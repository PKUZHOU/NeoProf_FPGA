// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
qzo1/ofihRE8xQuaPrNDT+7uxK6tOzMADFmkQeM+n2zd+ARTDoOdDYEa4eYW
jT3vyzRu43jJ2LHJoTkFnfmhm4+H2++lkikWGvqPz0vgN36DhmcaB+CNkoq9
Ss0czlchvHEHUPcoO+tPDEdRS1wbtBPKHs2P1IynX1aFdaXJchF//6KfgHtN
bPk023HQEGGDf1ArBjU0vs4Y8v4fl5czdfRO3/AxISNMBvfr5po6ncoA/Y5I
L7l4nc3oSPwomEeJy7/ryp/sBOphtNqMpaYKhsbLitJEqGnsyOgZeun0KvJs
asg689YFHiegmcIfStHxTORG5oMX/cu9Y61URK0oog==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Uj7CxatsM1/nYtFuKV3FxcySxSaAZnFchAoiKWAPAmzx2ekyqwzi67v/bc42
tlchOVgaagVwP7Pf1Ks9xL2LBpPmyNoedi0SRC9nHnq/8j5UDKkQPHEuHfqR
zpd3mvzqP9Io/y9s+AXWxLGA96FyDmpqU2gYbpL3XXpiZSvwth3t1SsbN303
bhlC3Pd5WgKijnPIV4lZit3E2polhLOMMWutTK6b6hgJ8QRyZW/PlSI6EykE
UXDct33hlP4SI8rkQTqlaQJhH6kCFaBba2PWWCyW9/uca4AAPv5b/c0KIkhr
EebLyyavusfGEhFGrew8Wef2kEB52Zr2KHzlOqNs4A==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
OBfz39MCB5cUkawoS9TXNiwtLK6S79s9HrndI4P6QjdZTU28BY7FC07FjrSD
Tgug681p+8oKU4gOEidJmejQcm3OUnUXdXD8EguZs5lRkvHQWawrvANlyEsl
akvuUHOtYGrZPJQbvjc57P4Oe0ASY71IwAvpLqzZl8gV1ZJYQGMQwpEvlsD9
8DiH3RFFkSDhqPnrGYiUd3ZQlAUQEtVq0O8M0dnKYJceoFKc19nAR8ylqf+g
wiz3c+a3gujzFb7ZMWtxneeIwtXTEuaxSLIWJb96nr+Qt2S4iM60JAL43e2B
47ywNASJPeFHi0fRjJMkSoUo83umwPfoKyl3EtNHzQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
lOqhIC9JjXZwIvarPKb6WJBHtDvhr6qGyKAqCBXdDsZtTjBrMohy4OxSVnGX
YWfRFQ7ZGrlZ+uc1/79hu6i9aBqjbH61DSzTgkx9fcu7iQsehlQnlSvWSr+m
fVa/plBtM6hg/7ALTucggryQDBGj1oBn1niz8FIIProvw8RVu+Y=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
oW2IBBjb7wBIUrHKdMhVDyeK3R8nTFWpSlN7eG3LVSC8daIiwQ8ONLGhVjNS
j8PeWoJ6OS+vzHOs8N6chomALTCNeV2cRjJnTlZSFZtBwf+iETcrhiEllDpn
TT7b2TbcRMMV6rxo9Fa5YY6NPsMcYJjExN8HN1b44yVtdJolczg5TdDBLDxC
yTyItNmQ/NwdLfQHIRC1/4b1PIffmrQNvecokE6HspBGvaE+r2kUynUvEuu/
1VrE+j/U049eF38tFjRaLhRBpvW0pXGgLhnciPZTyGV0BMq22j+jSL/vp8V6
jcQkmzqA/Uy667cYQpfyUMs4RHbSEkeJasA+jvXy/vL30/C7VgyEh0mT5Nez
aVdQ6b0xRegPiwxEARgVQdKCoUooFP9uVYeEZyArhaoOcSgBdjKKnHjpoJqe
aNJFqVFjMBZ0rDZR75ZDkqacw6MbIaYdG17CbNePWTGE0jMwQ3c14FWTue7+
BC3mVTgV5YxzEFflDiniiesGWfm1FbBr


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
OjSgeCYNYjMGLpk0SRdlbNODADIkYbtM/Udrjvw0r89CYR3eLFu4/BmHvq+M
36UUsgCjf6eYDN8tKmG3KsUPLZ+7NDukEqMWSQiNqHYKUcGEIi+lCGJaeWxU
lpjm9dF962MbNmjMkm/kTlHiZLBklbz7cYQms+7AiQTISK7mQZQ=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Q5jEAZF4Gh7J/5Mv1/EsQJBUHoyLLntlkMr3pPkKRcOk0x0nsYtVLKWJ2Mh0
/+Lu1A6/62kdFZoRvFu+XmKvE29nSFzViNnBGKQ4aGbceeqaNVQJQ/fjo7aU
WQ2Rmw3KGraRSBFJi6rnaahgskX8xqamby/7pglgrhx66dIaXiM=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 194128)
`pragma protect data_block
wDwaqvdZhqHi4/JiJCAdA2PkRjikDPuzaDITKkptdPtSYlP745k15tl/I+Hf
DLqNefYMMOfRqXXOS/beRxaqnH2bFqI95WBoQHvfVEhjr5Zz8mmABUJaTcXk
HIj+M5TZVjzhTu5pqJcXmfTkwWt3F4QP7Pk8626KqAHoUg6UQAuDFT5jOvPO
Pzn/g2LgUg9FhRz1p7QCrioFPWdKJc/82YVl86lGB+azqof8JkCaww985kQv
bakK8fjjYJGL2Tzbrh37MIKp3l1aNe4plv1AF3tyDAJE0rnH5caDgssPBcna
LhmzYbmgwo7o+luXeHLDMMY1v5QHIxwsTV8kEyp9xF0i5FS31vs5hoafIR6m
eR9+oltfDVF9JvBETQSVUcCiD3Px5RLE0dGTIyYuEbi03y18pY6Hz9M+4QCf
5EJMnI/RiKIjfW9DE07ISOMmhbzXeHOK2BVxGakrwd5cMFTDmp3YALBhW4Du
V2aKR3bkC3GI4yj0ZK5j68/PZ8P43U56HgccMQURIxInVukYCZYaeLoAKHeD
2y3kQ6Ct5urDOZyvyFAcwAMLkdp6AJDxfEnEaunU0RtBm1nRZLyhqOKYftd3
CFJ5KPv6oDzo+Y4a3Xp+RcD2pZnuKr2iITbsip6JG+W4Lhb23EzSNwmIwAh+
omrLwcoIih7MV27XdvHmwDncpEXGh2av/pd2ovkrlAOIvVFeRfBVs/Up8ybE
4wlAfVEim3EPnha2WXOip0fCJ2tFYFx7J2BpF+69IsdHGcHYlE+ItFpiVbC8
xOx47lIftjD5b5q5VHbFQxMDQNS4k42y3dg38A1rjyNkkgjJBy2k3UtsMMjb
+hLwD2kWcO2u/zkRkGxSNMixQuqFlaUaHIXXb3yUlpfbWdAsUdlCpOXXlI/w
cfXf2C09TY1rJ0FlQowXCVv24kMPVhgRd2TEZ5sv9q5GOocA/xaqQ+at1JKM
32vEKtK9b0yFKAQlVo9L0CfWQiLz2ZPGVSYaWJY0vK5lymZTiEsMWNQgOPpa
hQRkRJkJhwxxpcTJ/hQwGwsBEr7bMpMilq36mRX841njDJeUohM7KAZUzZOZ
zqjbhJHaoDYbV/iMK+87on2gnCmI5JzxnA5dfX9pIuzhRtwJ8cleg+ctDQa7
kvXlVZ3IzJ4U7r7LbXtOPX3hOpFjUyHcoK8erme+jI+lHK5uBin+IXQyF0tK
WZU8ctDJvu1KwTXy1rygjSwhx/8zFazTu4uSPqoiFmZmGPkgCXJqHto2mwY7
QO0rBbIAMD9R0qEYcVQGMU1dKLP2qV/vxZzLAL26trX7p2Uzk3UfnJcaICRn
IVzrY3lskppv5m0wr6p0LvMltJ+rd9d4dJIsWaspoc2kArAhZGSkh3wQsaJ/
oi+Wj0DKBqXyNc++cOjLGiTDWLfju1bPUTU3rZXjITa0ORhGMLB3l4epCjdA
QXK4i//dm7bn3NdBxmrLVbim4+n9L+Nh54PZ/P3UeaaKkYH3dQjG9Vr7KDz+
+kTL3Q1BHs2GTZ8nptXdSh9NTgnEerFBXkZ+IGS+LYPm7UvsRMw2uJIO55/K
EgCrYYnH6pQKRKHqhv03oUSNtrhmUW4nNKK3QTlQrXJwP4h73TyQZALr0IdF
e+JH1ntFzcDX/BMb/wzFjC3tE1I4/E+hIflg++sN077I0Csh9azzM3MsQnXa
poa/Xzcpky77gDxR4FN+45UlJfamQkYYlXnIO3H6GQF85B9qqNu7O6lPT3EG
Lir55YzyQLd1vuq2eFqD54lckVPGEV+Xwiy3eCiPFg7zFvL88qDjau00n23n
ZykaHZ9ANZOCiwWCkGLCJyXUQmrYwbcB+CGv3Aq1+Y0qDtn28tMze68a5x02
0Xb+fLukktDLV0SlXVMOeF1uWKyZrgYUaq3ZlnS4IGlwap+76nerpYBT4wAc
Xfj6c7zczI7VqE5R9WHaZbTHNvAAvnPRjv4eRwe5lpxlFmf6UOhhFYJz01wX
nzX2uOaYLyx7FVGDLvuOZP7ggNqrjxXkeTDLlWUXApbGz4Q64sYmJi6my/u3
qYn3Zmlxu9gOt5FZp41/vozOP41LQduEYJ9vO8Ju6lNbyBIT5p2fReVWZz/r
vagO4pjt0JMr6OBW/B8IIvXK/lXWZxxUV7wpn8VhDXzUt/VNPEg0KC2Susmf
zkTl9BgD3KFDorGiyOqOLfkcTXxg4MbLlJO8hE/LdXgaPj3/exKpARVm9iyV
ORneoaZqOcoo9gMyWRd9H/uR3DMKE9YJ9GBopouMaUglLr7e/ZFcGSIlSyLo
vWsWlh2En0sZb2AoQPuCDmgeG8DZX+ryJBPCUBE1dWWMHSQ5371A7/9CWW0i
7LV4rSBVUC1udyZQnj3FKrwIxcnowZmtjjMdDZZq6LPc4tXZMvG7CNgqLoIP
uwe93lqbF8ZHKDrAdHbudFxSULKCOWeOn1nvJGcbefuE3gED66gLUVt46j9L
PJ2itgY+c1A/QHxP/iEUsNcQjR2QpP0x4jY5pJ2QbXunj1H6eab1PjMM0Elq
AqhjiGySxWymw3qGZT7Dz0oIQe7ATsi3joctVIWzwCu8QXrkTSfShjfKToVF
D1rZSYleyltV4u4Edabg3P5m/lD2mcIQRS+wyI5mGZUMS2wmfaR5kqKKbWQa
zBTAsMfdrxUdqaTWQcM+8QbiFd2aFYZ+4Xe3HH3sCO9K3Rc25buAqfYfGUjH
RRE/WjSfQYfzzXBTaKa6YD1kUO8sICVnAQ+ya8+LnCtEducNpITYh6MqPQJm
HS+GwLsasSVGT636gT+Z4nxBGwUhFBrxBlzrfqz7sJLyaUkFzxuDWVsO7X+2
yaDBTCPv1OomcRE5dyBr55V7QhdBTTtCQMOVtWl+yZZhd8yyGC4JhH5oGiQw
8v7jn8gT+WjjNlwGKEweRQP9urYTNdIXlaBU7L95WXhK806N8H+M/63rQj5E
DkaiRKTT5oJbu3Huke2iDTZ7Mmv9hm8gWit/P44UgebgPDqM5fxcKVzl+3nu
aOhT6CKz4klvpgtyUBwCWk7P+yHx/eZZhtitVibZBPmLOtShPqddnahizk5n
a2WHlwpp6F3KwNDQFkN6zQCEEECe4bMky1+PNddDRnlsq47gv+30Eqc3+CI3
/o9bDPVDfxPc53voZ2XSV+9zvkPJZKgVfZw11dgg/DzjtVRAai5b8+L6ex5E
RokoezkKTSCZFxPCBlMwhBP/26B8AQ/Y9ZkZTCU/qb39huaUygA+oPBtks5D
Kh7sRKdLdsDJJRQBbc4l0WgWFVFrMftyzOWLd22w27o0cB7hQxhBfxc/DpPI
gtJKGPz3MZzFh3/LlcO5djGyCcwSxGw4jfbd54cJgTy3Ui8RkAQDuHUofSOR
lAks+UwDVlNwv25MUQQJ6FbTqDPFi2PsNBHTChcK9vsYkoOexcTedMz3U2tL
L6Le1gZHNfBLtxLYPGE3ejON06aPjDvb95czyS2FrUOV0l/RbTY5yWLpkOJq
DSzPc6hEBaUtvyvENbbXtu67xvPjwVgYVancRg/d2AAsbq3EZuufxS9z8cVf
FA56tm5EuR3AsYQJTRupez39yDa7EgAkpcICgfAJvYzNmlqKTqLnevg4N0/K
pWbxfwpwFAELs0ZUgFTmHs73o0yaeWjQHK56QghclOWpWl51qL111lyeBOxd
nFOZ5m163vBbWHrF9IwCGVqf5QiW8xHik+NQefK8QVUkY9H9mWFbynhyS5fT
hiFaMuPMjwiNpO2gCbD1GSa09ukBxBqhRg7LjTry4HrKkA4Gk0Y8+sMlpWzg
mJamqxH5GY5dm5ElK7EKvnfqvCKP/co64JMrFV292X9q+sN7BD+NDsEejMnY
GWVEeHF27UXFcn7G4kkzKzeCJXdYRJ2PAwbDeoNrKsuUakCwtxFhtL9fjZ3P
Mn514E8ffm6daTGXPS9PT3rVgAM7SDwaxwOXWQPD2rhAI06nwTLteMNXbC1A
SY09n+0GngtenrOTrvSMmAp2Iinnq79FsQf0bpfPNaNZRcEBK5WgYMjPJnA9
skSFYDMeQKlOKwPTDTb0m9xdos+TPrCCCBxTLQuiHJu9Alwd3cpBUUeChEKI
IvV7F4G0Yi2/lM2NniRJQBuh5QRr/yNUwfnWJZlDRNL6XTGCsoFbtasQDMx+
d+1Lr49SxYe9UiQkIuq2jxFUKQlI6CEgi8RLShSsUvgVmwz/47FIdCWGg0iv
CupUYK5bODvTg5Yo90Su+IXoenBPaPDqghlEIpAGdQy/jCOfKDfipqH8c88b
+6noUMNCEm0NnQhU2R8N3AO3wo6Fg82oEiH2qePCUDM5nvgewIWn+Pd/XBAD
iz9XUdKU7GyRPoGE3+glUm3A3tBxgt/n0IDhp+BYakDstUjq5hJI77sBhaBZ
OP7iJtSWGKUQxZ5kdHYNuUAdydISz2+eMIEGaPtYqY1egtV/NdOngEvPcdAx
Z98BnCRBbXSp46RVgbOPVUnz83d0F4yMrx+LgBwbJfnwUA/zc7YCffzWdP0E
SyCuKOU6eZGx/NFISch3Qv3GYrtelJOpPYp0Tpw8tC+m/cWUWJy9dZqX3kR/
L+YJgt4jVyFUR7dk68M+S12r5zQt6WS8VRptXM03xQ440kasixyz/3xAi5PF
x2hBfmD0aEbiTgnY37432aT8WLR4VYYokHWO4FgD4/iAFsv8qJhkOeLoHdan
J2DPQRBCq8b/TZ3mVp6jetWBIBf9etiXejW26h7XOZc9g/4wukVSxNo3E5VE
hoRyTfFOy71lkmBMp8crNzrr2J4lM2oBCIJ2M763tpb21lJrp8rQAHMvJunR
ON3LZoBr93PfhnLLTS1SIKntuP62gjrqbyMVLrsox1fVHuL/FXfD1vpFkgb6
LSV+1JzFH9RxU2jdCWe+93wfiMNJ6vd0yWTJGQntcbgTie0w/SGic3DdeJEO
LXg4t9bNMXT/jpHo39cBZW5on798Fr0ekD12xQ0+QBWFeu36AOhLLUQzjvPp
X42b3nsG3SEX6XvDRRi0KsdIMdCJ0SkPCTNPr66lGo0ZyvTZ3JT5Vt9q8TzJ
221YcUnl9p1qy+uJ+YUoA6qqMSGsfAz3vuHr6Vnpk4ylJCXdWOOPSvV5F2Lq
visPBS1ycUOWE/SKyZXgekHDxoh+ZJQ/C4QlMibvy5EkSbksIdKbojPwDlez
Xb0ZpnB8AUWM+9Zbh2+itIPVL+yX+wpa085bgWcoVKLbMM3Fk0HZ+tbb3kSQ
rCWYs3ljIgjMpjCP6MBrMyx4osENPFUiFo+r2rnPBToDjUp5OJkHw4WPOeky
oaX5Dk1vuJtzQnoUQspCGuNN8lOXmu4K1PYyZOxy5G3P8A7a0a/H5LzaMMo4
krTeT1HlUDMqxNATr5IWhFWzK1LH65S63YuxnqlHTZY3gkHYrOorRGe9Kwp/
T52L1VPtkGQhn5BQurDt8lmSzTY6QqTaLncwL6o547jhDPaUFkFzqENlmQ/w
jN7Wdcd2Cyor+wuc60/VeA53sN4sb6+KdiCqvtbGUYRuZiudynhiVAZB6bLW
ETd4yEixspL6r/fE+Hd905uvrrdMbxqTiv6u9FrMU0ELXXgw69V9lxTcivml
v4sack+7S/918mlRnpedaoWbsWRZ7RDUwv4VgIVY6qdPHIsUb5Bco3Zjnq08
w4Qge0bCZOl+x1e8wIpRxSDGEnas4eMj5GaZhtJQ8NbBEvs84caiKV0ruy3O
VpD80NLpeb7h1jrThAX1AtewkP4jihXvJpOZfco631V1OCQIgu45KDktDGeD
09lkM4G2o88yspQhUBBxq/SRHPCuveCT5wrOSRNztj1PDIUhR/DqRyKERr2W
ekyYDtpfrbqMgOHMLoCrBuk9eL7+pngkP++soVDeDgBpQRJw0D9GNkW6hIqa
K/nERx/WUd7QumLhLHNRebvgZIa6PGJk8vI3x6POTRVjYVNmveltLAV+Aj9z
9mrZZhBv5OUwR09eSFGDAPeuK2QN/5/AMUzwhUCK+LM0WgYol26wh8ePkaTP
7/0uEE48lQMhGjg88wQ1iQm716GN2dQ7ihg9s4+dRCV8MjtNnf6BXE44ZG9U
ZWaOwscvI4iEhA1BbZcfPtPQcjqX2j6IBifAtwfSS/3DqFYpSPdYNfG1e/+j
wxcREkuTIKtlNSJ+N8RkYHPzFPvjFOQPS9BPfUjeqeKgD0UrN5bCbbHm59fi
xTjc3JfLRC8cT8AXfJA162TU8eIcnGpFDHvIMCOpKbeTsEKO3Ef7p7BUqHtU
LBL8P2F0ks3yRAcKAuiZfOQpJhZCfimrObVceL9nucFSULVmgUdsQ91wa+Mp
kfBIxUB7AnXbJJcZhjWODQUG0A1vNv6AyQyVxPW0azRHK7RNtIAeP6EQrq2h
craxWeR5XYSTZzxfRUf3qn52s2sAEco0s5i1MpFKVlcEqBOqhEX4A4nZPaVG
CBXEBkAelFpQ1WSBpUeVscQquADhOHxp86MG1trvnlEw/aoGm52ZQvheJGVZ
H5c3pVSvROr8EFe0YYeIOadi3BsLk4Y+BwejqSqmBFnQCNzD6L8h0nLja2Tv
g0TV6tfoxNaHmiPRuTYK0b7XJxF9FAdZyCIdCR6LQPMJgVCY0bmvXdxXT40j
7IKxs/2b96VM8J7M3SiGq4Vb02F3oRjBHXdSTd/gV4rLDfYRUfISCiheLVmx
vE8eHayN+J4iX47UJAMah78CdWXn6811ce0+itYrgcVRueweesPkUWiKNVIB
1XeOwjISZx73BjMKmqRhWFpX7skfM2GlbdHLvBc2/MTCgN/3FFprWTRl94Zl
Jb6Lz2Lm4HFeagSam+aJcq5yVJfdrmDVEe+lY1KAaJ9BO/ETzqOGJ7bP7Fu1
OODA4DVusGzlYAvMw8flZaG1sgMh7vNTZIS+9MBuUGz8c8mmBtkUFeKYukGq
j+Qn1cEl9W0cR9s7m3Qdq0dKPCI4wBHGMLjc90NfgXyd8josfGyrrVgF2QXN
GiRIFioTdcejhY9fZbClOrh7Sx867j8Q+ss/fhuotukR+Ma+p4z7gRtghBoi
zgsvpxxBZDRPLevDyNAfa1eqdpL2JH/3yepg6G4gP6ZdHL65+HMup690tgoO
eftU4R3f6lwm76nPwr6azKgaSSKNAhphLGmuO/5VuxL+Li+KZifU58eKTp7x
8fu2E7jP7sm1CMNLsqF5ivAQrIimV1+rOFQmoAQoA9PIu54kYKe5GgXS1xgS
5cMf0XM8+TxItgEEbtardshPORJYvbNe64/iRKx1Q++OG5tfhyRUYcZ/3Ay7
nnWfnsJ8n6cOu5vSEqInSve4KlWOQvi5YGz9en2HArVrPmoGkK+ReQ9AgL6R
hrDHUiw5oLPjusV37awgy66Pz3fRFazL9e7nwi7p0AbpP/dUq30ll175Wow5
DB7rr0N5UR1m+bCkGUZokK4aBf1aJ6PdBIxG6BeCQOtk5fnS3VUL9zqH08YJ
Ie0MYxy32bMIALDBYyTG7nn6pJnZWFa5+CBAsMnar5m4pQAxLtFipzsnmYnh
YefQuZvokDmrl18YDqdPLRisztuCCpr8vy5l3AtQmI+qdRX7e/9eZhE3QeBS
JqMlK91oAkCip6vFwg9geMVJltRyhJoUq3kfFizGriB0jSs+Z6toiFaGGc+E
u0SD+Q+8w8plWvpOOxdQvh5CeBmuLXYaWrhAJEvivYB52XyN8QJxBvtnfrDs
74jGkIU7N5U9Ak9+Qje+MpAV/tB1UuuzYzQ3fa4jq/8DobFIcG5yk5oy+ryW
tmDU8xuJj4zwp3kH7ti7JMe2LNBLwtDyvsh07bWlIfRHzw98FYwY5akArXsI
wBbDV+MJpEFX7h4r6D9DYJWGuHDRVp9swfaEHkDainXKU40HAjmmXrdpppPZ
x59ImrDU9KzmfFoLnI4LxtIP5eel2vHWgaOIZPkOp7DOBDFAjoHzI2BxH4bm
1YwySd9VhZoFjy81XJVfC7sBW9jKR1Hp7JBmiBJqbV4tG1R+/O6Rsbd54Fed
EqB0kGmt9PlyJ9y1F3S/c4hgmpR9Ov95N4uS/tvW4QyCLChWvPovbpOJZ79J
iHdHokSUL4yBSISNILsL7ocDl7H2dkWcfIBP9oc4F7iflx5R6AmlMXCkPu3X
lva5P4svIt4UZIwhHZeSkS0mHn1RzDGxv2YUikKH4pWBTYNR6iFDVfO2jk51
F7IZYhCJhPg910WtR4L1MBb8u6sc/ehhAHYBzilOEY9NN5+ySJ9tqs4ksiIJ
4SoettG5c7YBY00EhFv35M+srpwOfJg9g3Gf/8XASB/AAXdDhZwFtC0qvBNz
M2P3XsNolwvRaRtdwsxFFo+i7df0CC4qcXJEqjdOzIR+4S6HaJ70teDoP07s
AN0T4OXWsH1QIg7xvSDMEFrAxQeQILSgiN43iWvaYgFo6AQeurGNHICpnp3E
oBzcJqHm8yY3Tz4WEibnQlCqmlJe7Gh+XiDvdyYXe2n2fO13FEt8DwWDippn
O0WpWBwOXYZp/StxXK21Hjo5xH7SglR7Y6B7lecY8ngVeytDFdFzqoBzfA0H
pCFNvIQTTsWKPOydd1qjFWxck8fdzsxMwsFba5lKhup6YzUzYwpd/aPZRMxZ
6Ua3qLyPVcu+GC4mzfd+9aXEPxlJHspPZJhxkSL/9qI2bBjGWAJWe70nR0wo
laqIN8ByQn3CGxrVp0oKT2KfwHnGD+DtHMmvmfnxjMz5NWtllzc146yl8l+a
7/rB5P5r0lnYTI/9WVkF+KahEXcjvqzlrtH7ca5QtIJlKBuIQ/7Y631aPCeV
9ITuXo5l388nhQGzUTXwMo3KuCkHs6BERxxN9VBV6TJnbjMZlcf2qoRDI5dT
DOa8+o1IZs+ZWIQ5AALYcdpSGi6WHkCp14+3/Fz2Gk3aq/6UCNXwFfFvy3Y0
uair3ADY+9h9deRKmfvM1fx4yGkHRT9OMUDRVO507MB3ykOJGF3hltyMk3tT
iivnOhj/M7Ve4AwWvC1bH9969VhqlO5LAGcGhUsTbR1ICedLGsnSbgfUCKWG
hSNLHchEFNLYEqQYqNU9QOyYfc9xxj5DCzBXjSnFbostCWLBjV21XbsbYm8d
TkX4O+tmd0TdrNvsz1znftzc2uQ/0cxn0lMbtw2yg9XnM0OLgJXgo+gf8ust
8liv6U+hTLYYRQjStKJY8Uzc9mdZzG9qIwtZOg1TG9UPr1VFUa/WAVNMcdYH
N2sbj1110EcHM343jLNdgVci86oV0rL74gw6dDng7KKPVrIr4gYT/B07IC8p
nclbfAfap2rPonvpz1IYolWJmPjErBO3ZLEeZUhmMF7BU4ub/nYybz6gPSDp
HeFmb7lvSqUJoZpzk8mJG1BzuQv6+AVEXUKGh+4lpNXRsQW/XuPTbVuHLwoa
N11MpuWnBB6B/B6LmT284wn/LBPW2y0QW2GblQeiXhVZSXJpYQPRJioJv2/l
OoyLpS5r50oZAcMvDzost32VLVhmClQGQDuCND+ghPCCiv0pXc31QWEvYhpN
6Wp77LYdclPwrep5fWPDV+hPoRVZlZPPyxqk4TbgUUPftykCXLMB/3QIa35t
0x9+l9RuWreOFZoXiasOcwVyzWsK+Q/31cKgCkJhwMVLcBJeUDxp4JL0HLWJ
LMstHcfdN8J91D/1wa0vtv3WZ1v+xnYQI8ybewYJmaiGJTw9kzEfErtkoqx8
9yehjsCW88YVxTJa0cH9tYdeoqYiDqtjfRFKinXII5HhCiniSsR4CUSOOWO3
WXu4P8jC5WbJcH89ht8MYTcJ3XE8xc2I1kYSaumHYLW8dFJAtXeLy/ykhapd
fDaevD4YSMprUpwop4uAphMc1fIOMK4TJLVwDGXGwdk4AtYIjAQE+ovrPvXJ
wHibVyVt9dpa/Isx6akqmkkUNzP2ijYBQWwcllFKrpSjVrkR+A+6pfxC4wTK
+t2OtQjdGVXfFWEzjvAihLa4ogeYDowNL2+zzjS2z98lOk9/ebkgYLZNHujU
yWs7KsrY4dQP90R9vMynNRDtimJfcXAILoWi50x9Vu0FLkbnUZOxoBOW2SUM
2I7gz6NdkRvaKF8HMsJQGOiyuTJXnE0CdXhd5JURS2TGcKUPcOmjkks6n52D
Mt5UBj0+LJcRCpopayslzAyie0FV+K4UI2sIl6DGmHTf4A4qwXiAA8tzc9iC
SdO43ija2zY0LHV1tWcYwO7fN4GIvhxfjElvuCdSMu11vlJMHYtk+7grGMgf
iOdyx7kd4RsPsofbZLI8jsZA4Z7DyTXKZLFKS8CcNZc7Fb3OKK6ho1XMfKly
H86vK8+a3zaGFP673iH88lZB9YxxEkqJFJ8sdXXnDsPmOpGonitDuw1ozQyn
BkhEWQ9wHvStTmXo5Z4HQTKmCJEGr2+gBEh/W39a+h0Ov3HBLboHeL9dc/UP
G6wQ+Kd/QiUTw5ghh870OM/IEeUueUXgzBMN5MA1djOVmXpsWEh8yV+vapNl
W0fUIGdAQgQztSpWTQFe2LP6PasteRGOCxY74adhxk2nFvvAEg2B9e0wTvNq
TKn4J8JYX4DPX5GwXrJVyrrD1zfUhlg4DqpgHRdJOtWM9oskMhxjYyAFEW5N
VXqSugn0Vd+Jkvn+nvH4cQSx/WmBZ/+0LzIk+GdozuqyqGJul9c7cDeae6Ux
I3hVL46DyVY1G590MTdWxWG8X4zLFGTXbLXXXoKey/4OGptPoorthgbsFByg
gosn0SolivLX5MsiyLKlw7Cnt9XFN6/pSs4azbadKAbLSYUYyIDhDNuxH6p9
hoWywacolGGO4WlFU7IJJez1MUBTL/JiFHtE64EYmhUHkKXkKn6IToNs9CAK
M/fKTwmZ7eRhyI2wwGME0FSs1kFOGkZWJxXZdMkAMeOJliZ6RUOs0lKPEtKX
lm59Pv35hMXCST21uYi3YP0/bQA8iFBlxtiHB/Jsgv2ETCQ6BXHn7Oi6vPa4
H0VwHN+q6lrgeog4oeehlWS54ncpJ7+E7zLDreQFirlEA+fZiRJbW4VsG3z/
f5QDgi2lOUMoGcvIGs0PwriLjHUknb5DwjezATeuXoUKSE4dmYZL/PevlGST
q7pyk8oDkXY1frh0K633gzhWNdjfYuCAnqraRQ+3jjdaPwo+lcNzkbjiEQAl
ybE2LBm/UzWyRIRsW2+pva/Fu5xHmavCZwYQ+kDcKKvtMo2qMiiSllis+mk3
tdGasaOpASuPGALaItvP7xhpied4N7AWlyyWqptHR2Hu+amsVp538hDAFrXF
mKZIEBrPBNsPZgunnsJJhN6zCpU7BC46nQrXzFdQcyK/xy6l1wsjieptA6am
AcWvpclZcixQNlLa5ADjT+SeNZzyoH4GDjh9u1byRIVlMFLKfNs0UkV3xuvz
2FxCaiPUGys4uklL/HHPKzD36m1Bzj9BPJvAHTQMwJD5Erq/mlQfiJiaVjwX
Y20Y42kkHOpwS7qt9o/az5GypyGrBAmuF+M5pYFISFDFW03wDbofSAvqjxxl
nDjPuXwlfJgzs4y0BPa+z5DxteODPDV/oFilLEM6b4ytRnn98TWymLmAog7P
Ip9AvffWS4Tvz1tWX7xqwg2BTVdjedMyJgt0gHkB0w7NsYz+uYpaLm1ghlg5
fLETx2LxiX+1PtAEq9XZJ3PokFcAty/TuqoHqs0O+eUM03omSx94xi2Ofc98
ZSR2tOc5BFg9wT5Mhx4NoTxwTQ8JXKBFj2R0JLysmZA6ksCrPIGbVPUcKLer
4G1JTmUCRuCaDCVGXEcQS+okmx/zMyO0n7upmitxTd4nr26T4IIowkpNXbD7
D8iEIdzVpiXgiuNps1uUJlpon76QUE/phFSLBL2C83Zc4iEMoOUdEK35h3Ff
onmdKA+jPaevormyxx9nEeIU2CiWBOLyA9jeVuHGIGzjIwW8KoQSvDRChgu5
kTBabH626H4EQGuyPDkd5k35GS2d7YBP7lQFhjAUyA3RkZrnYpQTxcGcnsxb
29XUW/p/EtW/nQJiYmZaMDXxGKDhNPEAjxYDrTyX9XQXbCtSt0CmeriuzF9e
ZfTILGhyZTC0HdssvtQnN82oWTarmuNT3XUrkxqO6+YBdHk9beCJ4lfQCgls
uj8MsKtErFN9f+gSYpG7DZLJSrkwek5KFSs1+XdsDj6lq3g0HZlDHhn9A046
iBiAHuF32u/7v9xBzaChYH+lU2oCAph+fsnpRbjgFFirx0e4CcQRFxaXcdlf
oh9yuWL4ogvZlz7Fs6q99pSk/+2w4qRmuKYaepFt4wGMyFzBVwoX1JRiVO67
DJbMGob3c9BAh4m+a3gse5UB0dDGx247YhxCXwV5z1WIPfZpMAV4bJLCfpBo
J0oQbZfLm+QXvwvAYoeiYGzWzrCq4K22ltKw8y+cOaXYBwS6xNBSTG0kZ9ZS
H5xCDLnkrwADZyfLDc6JQ/hvlwSHN3b0muPBHGfsmLxOYPcFmoRwTmgQzvo0
mlPfDJk1GT2auTmEcrtmEJn0rePv2J2Cjjy0iZ5Y7sLvUI+KfDhw0fTuu22l
n0o2ctXZLL+ZvYkJ3/HGxZlAPBr3DnaAtW8fPpPQH+4nRhLic6f97HRzqqTt
H63pCUYtaIAHV8Odcx4vLLwcDKquh0Zuw1FBUM3jlcq7HlpUwkTJ4gVOsS53
sGHFDj+IUoPE8RMWvZXEPSqHQr6dyfrmZxZJIzhUKoFMBNpQBVvdSKh/7wpP
jvoc37hhdjqSK42prL7nlD1Puz78Z1xcskHkdlAdd9BuCKQwkILx0XUarA05
qJws5seGMT3CtuyMkCGDohIy6CT8HmzL4Bn62y+dB4DLKoq+23LihBWEoRdy
Z5irE9CwR2LIJcJTFynIgfywg8VX3k4GZV6ffnR5V90PLm1OAcsqmXokFDrZ
+hMs5QRCZwjXjPfCUtau94vyuWul4io/ur8gZBtUaUNj3vmiYlkbQoVRHF02
sHFez3hA4HXRduVRcWPAGG2Q7h5AfpBXyt6Eo3y6iSiHQnOYvrEXTZNp6TzU
rCLiNSnuwKg1sp/1t9n9zFrCe6XABlUDGD/nwNyJW9HnxIRjKbuPWJYCbrdL
wBaReB6tLGqofmzXCWmY5/4u7ldrpm/HvTt7ViEc9rpqU+sLAJRnOnDYLQaX
6PakDavyi58hljYmCh3erPKY+fPHpdx1jfzIQJohF3I2EhoOAIH6Zbebcs0I
L9Nr5lT+czhPWOxX4y8jtw0EE1Vct1FadkmTmXuHbcEv2QtSmQqUerxB4OOY
XswbE3RN0fZO1cumYa1CZCnraQeRjdc4NGfnapZ0Qmnv+RX49AqgbgTWOJ3I
Yvu775DdrXLbur4gBkKZ/jPJcWn81HP/0npTb/cKRBbP9FfYZYqjwFhliBAx
RUYoZ/KCXbGTz1kJmZslUOBaOam3JmOFwkR9BHj6Xlpu28zvHrdlR5DPPn+2
Bc+LVYOSQDXNkgiRMeWA6nnrQkC1QTtr7Q3HXYnsmqL1U2zCAS+JEXeIRwO7
e48i1q5yAmJD1DN+rPeDB2PYMHL1G59mknfZEHokjpDxg7ptuG0YpvTX9LSa
ezl4ZpKLon+2p7A4o6Tnm1EktVgiEABddtzh2F/+4JS4KfmQZLUghAsAkE8Q
pK33R+ozmwfldTNJQzFhzYnS0EWz4dTQD9Msc15CcSPQbyDv/e4Fbd3CZMf2
7+wvEPgumyqeYWKzAdIsiK9wEiXEShYI39ammfTBxp0lUYsG1VTfBtOlF4S3
sx4pYKz9p/dLWPwo/zhuaWMj82bPxz5s/k1bo53T3pvbZbdXvhmvElLK/ifY
mnCNaHlnFIMzz8Toid7JvSYlQb8BKHrZlcys0Uc2Q52ZR2p99Qa/ElqB4yFN
nyfB+F7EuEumSZva45uJUtYf6p3H8Jst+mW7HnbKog8tGKuaa1hKrP0HJ8oZ
vkqzZqCfea5VMK67usuWcDZerfW1xNKOa4z3KpbolofI9Zl+CPdv33zRw6G5
ITePktq+EwtejLS7ocRFrmorK0AGRCLdRQIcGD5VmXAxUw7lqi/x4iaTBI7x
VBCQshDT5tRJ0uuGmiJsJqbp58+K91jDIIGBANPHw2KeOwt4nSOh5cJOTVUU
1D98Y+CJLgVFkR+KP3E1tHjF7tDj5ZegTsYyGvj98InUmXQdi/OfqbXReEJ1
AJB0+QT8k2zPbQl9BBKH4SDbDE/dTZF36zyygNwX+4H/yvfJsu5tY0E5TzFW
avN8D3El1puG/Pxa+FnkwRZTjc2ydVo6SgqwvYKWt5lj7+jecAlnBbhtr8AG
PyvcfEkK0PAINJ8W6CjopELC42kvDueHw3e6Hl2UUqByFQBZvgNykIHoG1RZ
1NHBgFPc4aCGGS19/Jhx8wA5W0HXq1GMBq/gIpucNsWyE1NsGPCyAnH+xAcx
3e9azhY9ZwngF152+TrRiQt+f91xfnXPiZaAV3U2VJ1HUxPOLTlSI/G24rOh
DAIJb4Nj2OpK6eikIt9CXMETYK2fUp7omPV7n9XFZwXxJWYorQGiYTDt6hDK
dS6buqZJQ5bkF0cznvA1r1FVVW2HmiOmwqbGbFlWEkuXHHj4fgG9I26LcHa5
RcqMgnMx97gbyuCSeQ9E6f+cCm8XNSETG1A486NVPkVnuIvv/frPukjo0PR2
xgou+flfOi/Q0Go0tPfyweSdxVFtypOvAVVsipNeBWxsVexgIrawwoAKHAGe
pE3pD3Y3VkrHniXB0DrOodgAqz/UoVXuokMwGlmQ+R3Wj4JBLJOj30RBUD3F
JdYwRXhKE6XDrj4/j74G9LLIVWCf1xHhSFrcU07KQVB4c9t1F4hjOPa85D9X
+iBA+c7lkGnjxzx4SwNr8OGEH0SBuYx+QiyK+i1HmyfaIh4QD5ZwRnpbVdYz
Y3IcdfCn4EuOpzLJtGSxZpS1Ed/Ff/GC/XIWFpl8qjs8h9wh3vCI+X0GHgF7
FaZWcnmLzwlnNQm+2JBJKkp5zk7NEygAWgLuQvBjO69jxlhj9HqG5kwWOJOu
B0cHVXZCI+mwBgDq3ObDV6QTIKk3dvHoZmG/U2amNJf/orNY2LWQB6HyhSYt
rhwQIvtoFxP+kfodbBUVCzRI4zt0sOjyLhMkTMuuffAJ+u+ObzOIIMd/phvo
raLKRvwXjHMy1dZxvX+90fvr6dhl2+qC8wX7VO1PeNKGS0qGEt7YRZBAex2A
o+TTLp1/Yyh+6wMQIGKGagl+xjbNlP/fLuFq3T6W+hg+zdLbxlnCyzatblPl
Lf9RBJf6CFrstnixx3jYaZy9P65UXUwzB5y2/QisXQEwt3lSx3hIF/aZEwWC
dAjCv3yq298QXHNUPIp8zA55TYo3cpU+EWtAOIZ9LezTzS/xbX/H60Dk07+k
axOQpyxn3NRDwKrRGZFq6dbPDs2bP02f44Lk+j3P8IqIh5fzMlTylNcjpPff
f3AkY/x7p9GV7b8Nbds4kcxnp8PmH5qYP+RD4AfEvlpT6K7gThvxaI1gortG
cSO+8iSDfG6W9B8MP2OUSqjkTOW9nvr/T7sYnCjcE6RE1kYxYTEJD4NC7zv7
XdaCI3CK5HfEcvlWOpUTqbVZlGLknLgAWety6x/tB/GKdHtW3Ul/gYnsIQUz
Qgia1iwmQBfM8PqC604s1wweZsEWa5mJcR7qgxV30HAE/tI+MJkgRA339eDM
jSJETpgNmtRAUAeFQKj8muGaTplOK+q5H6zZfwmITvKLC8l1cKzewMEJXtoy
3EDqPog5pp0tuAf4n+UGzcFrEtdbS9eSSrNKCLxA3AuIEAXKHRGoHNzjjsIm
GjRSyVK88+K9+tUQHgGEP06G+ekyqebw9HPp+FARRNn0mpiscL1r0IoMO96Q
bfOKe7UQaFtjtLd/eSxgji54gD9xqpXrgAt42hrGYVNIMlC6KuSjaNNtGOxi
mJqVySQOfBEwPuw6M+mR3yRvsQud0e2RLBsS4V8sqiWP4+qQZ4RVBBjIiCNm
ujHyVroSAUY8gXvvpqDLovIhM7/t2iFURbMFRoFRA7By34YyzocpE6BbQTgm
QzZ/B5CPvo9yyxsvjtOH0UiarVlduslHyv1mYwRhKMQmC5tfl2JjhSSUqEGD
Bm7mtZ1LEosnwn4AskOaZQBOLy4crL2sDWCw4qDEXv4Zr28CIw01lKVTKaKt
cAl0EtT5TZPQNfDbQv+T/jFMbMLL7N/oPDjLKqtFFOObcOVdR6cqbmeae6ok
deetK7YHVMnufmijzd5nfYekstq3ZSWCI38jX8cvYGyVnzcQAkD+XusOLW0J
WWoaqYrhsqX/sdY6Ec9bhxZhTAryxqWigZk1K0jtkPeaQoxGgYASjyKS9Q4f
RQicui/GriYE9GdYCg45EZbyyaTB5wrDhtgRJv29bD/9zcAvtvRwi/8Nr+lj
De8eQxiKpQWL5cGWZT5qkhev0Bt5SqVeQ+CMtD640WK1NNZumy0W5le/a1bk
yPn9RXLDdsDO8bXu386RukCkac+Mv8N161zCRwXHIK3bdepk9Qb8jmTlatIl
eJ31xhfy75DEccovQj2toFvJIBW+2ICsdEjHBlMYoxGvnSnl4BUZ5A/bola8
Cq1PxtdJTxuFtNPNbfnq0BGPljZTONJ9S8EoGFo9nldHQBSxdd4EsLsDhl0V
td/8K1kFuNt8si1QM01eMoXeAYTnT3IW6p7w0H9vXvFmhYneDSN2Dm1pGwnp
5y6lsj2B1QNtLySFdBDQ8DglWOwBjgrao+LIh9TNGQGgu7W9qhitPs6YIDPR
c/n6U9Zj9yiiKSUREC632/hHR3sVXTPFw8Tyyg2REsYB2/1Y2RdADv41CXba
WrpfyMVIbMlihTrBEYb3b8iiws3nhRBDzsVsJsUORhBcFFL4PuqOSKWjL/L+
5liYOB4MHqXbBk2lxnHCzH2Pt/reFxHjAWkQPfhxsY2jf6BT5wsHXaHMt9ks
B+7CI/J3Qg+J4umYKLsgCGr3WZPBddjU+m0VUBrf1N04D59Pp2KZtzXBp9we
RIihjW0ZT4+JTimARAiHO1wHihDI1XGoq3m+LmO5CvVW28CnlfhrEucsxduO
HX5B9RsPK/v+HxRzNM2ZesXSUKtH9kUcWPub745OcWSQbABiI6XoZLW5VSoD
HgX7zJ3SGleHgjY84rXZGkSekO1NtsfYik7Ah6J21faIdz/7HkfPkRdfYxaq
Kio35gvhIKd7Xg3nqG0PsYv9iGnoVxJaqrV6jltThh48ku5nnOakhFkuZK0S
VJi/hLxRlKWMF7Zkl2Ey2QcMIME9WUAGiBS1Qprv3HKSL8lmynEHzAT03lfW
8+0clmmYsjgkd5tHtBI4gasgMC48LkRv/4hFH2M1EGJz3ieN1C0v3RTg9NOy
qscL4mMXBq6eHLdUBH2pUjm/5gmRlUmr79chsI3/WJ5c/QnU9nU9dO4XrOXq
39mBX95rnwVMiejSU5qc8UJ+bc0X6Y/3iefpkuX/Con40EDr4ynriGCpKDJH
8uEDUpycmjeW5xaM3yHUOywdIaXpajO8hgoabKbPQDKuhZUB2oOWz6cgFLJX
DX3XsS5chtr8bIXW92LAL8x/mkZXcJKrNJF4LPpYoO4q8WuMWEbAv9ov1TdQ
n8Sa5r6MQ3j/7VCikB9veDKdjY0kuA1NetrZs8a1F2C4t0xxHm419+zmbJd+
UL03FBSuazbtNqKmwLyNeGsokfl1wn2CtdygBuBCx7VPhxviY+E1wILTZcxD
niUXYVk1SU3/OWKDkYO0cOVAp6IqV87G7N6wG+MA4H0QMXMbZJ2AxDzZJ/NB
e4znT4XtRSJgGJlwgunENYC1xPEuHmnFE6eQGnsoUC54R0zFpCChuLdOpNie
qFiGtRcUCbSPY+3g52iDoYfta0V6osdkDDslwje1qkKtKKpmGQdUaAvDqLUy
UTrQXoRrkDaSYi+iyHlKYaDAGF1Z+4A+nsfVabVKPOWJG0iNQBD/q9vK5qAI
hvohijELZXeE6ARzgUKxsvxT4KuWHgQOLyejOXRCCyiWqEniMzSUoP0/Jqsu
VzYRivur14XgAtI8r4CIFbjI6qYHma6Yr7Bqvd3VFJMK6TVxBfsdPIjkNXbJ
8yjOArBbNApHd6kgL6dzWd+ZAJSI7a2YW5AdEpDT9pvJm9fKcscD14llJwIA
/K1MEtkqH4GLiVvxR3NN9csbDSoJNjwyD8kOHObSVpA9evEGpI5H8bE75pWF
YUNzmQpWWB3i/PtYqxs1CkhJpFNygmOAh3eEDGed9KVj4DiFaMiboyeHaaoo
Te56yXFYbgvhl6fDhyYpfI3MblP6Uodk3vcsfokmMAuDJ8UBT8PObYh+yhjU
W+/kzAM4Hh70wRmFK9sdhopK9x80LAMlvwC1yV/DqvFza7yBHFS5Ancd0/Ry
OmkUeE5BC83D0vg0rQz+CFoiaCnoHauCrqDMqqN4k5o/0Op7GwCxEY099G0C
1VQpLEbuV3wFP0NhpTqStFPukcmKka28SHxCUzPrl2I4nI94w5wZTM/yO656
D1ECdDqsVId/lWsKbS6o47YCcF3OguacdX/nD05ysoYd3FZ2kerrYfoN9ALH
XGskRmCKud9sPAiF+wzDp4iapdcPLHAYy6BHAMqNq0EIuCLFTNnVlyDK8cmY
ONX9DhMksDNH/e9GVv00UgcR8J1d/OaC8W1iHs9xO9CMoGxVa4Hy7b6pRSNQ
2XpX6TVEvvc1dbq2PQNi9YZumb5Y/b2zrXQjQMo2Fn92s9BmS3ZikV6/pL8s
F9s92I1bN3J7ZLpJZeBdzkxo7vY5SzoEDWnEEIzcWGrFyNBp/Fxnz0Sj0KYR
HYPf1FrJb3zm5HHwuwZ3rzOTws0jjz1l4OiNFgdYbIIydFyh8854NI2YByhN
2NE7e0+JtRQaauSf10Bqh6o/yZWtaJaF58OvhvTLZFF5DS0JjJ3ln/54FzhZ
0ufrBoyjv/Ki0XUfj+bTlwFmlkId8Dqk2lw8diechxOh02EJcBTOvGDxMIJi
Vwi+6gfg2kL963Umck2KdXZ1t7OgaPMEtZrljFXVSAYAwWAf92xHH8VUVRGx
pIHIkeRqWaXAYJX23tvdvGKVt3qGftm8cCoNvP18D0gLN+YMtaGFXl5SjWYE
SYfL9tuj35Wd6uLzPAHa1vt9YCv4My78DHR125zQGjB7/QQtWbuHMbcIu8py
zDCkXBgoO2Y/f1qk2kjBTn9ppfjwZHjEfKEgiHamtjCZmwYoK3zfpfVfDORY
KzOGACKwu763lPWtLDemUA5qJKlKEY+0U40WcVpuikQ/9i/0ED5lSnmbFfAg
ZZ5NGIq6Dv9xaDuGiwtcm7TePIh924ZH/ap5cUt0LCeHIJS2FhP6bNo8ddny
jPS1JMyR0dQZWnX1iK8PmLIjDVAxDVUzIoqieOiEKfCjM1u9ANkppCNMJFhe
ScKN25KwRHacT93ziJGwYZcrdXeO87eo9Krh/lfQn4k1yd/K8xqgcsHF7OnH
zUwbBwQYCMmgb6Xo9tC/Wu2wuCsu1WW5LjTaxcnTdBT37nhix8EYpkXLdyUL
QU5l9ZsS7oAz8aRVdAYwPMSuYkh8wwieiERtM8o+LklfRNMtKDW9vypN/vCB
Mhg/GCzN6yXO7/5tIZnaFI0N9R4tUpTPrIfWMjGkk/s91hN1KKmP1PxOkXUD
1vnK9LFU0i5muYpJKww9HhQd6nFyDzin25NX4mjnPwKiSYOXb0zssBcGZJKj
CzZQz8m2pYyamBy9uRKoydCoDsqz3y8jI7+PuSOk3Wa4KvkposWlZzDh7SLf
oJLsUW7C+RqGZAkINlIqRjguO8/qIcV7uRkjSvE5fCMHysw6Ll/WpdejaVpR
AWKWvVHox4xSYo3zPZni2pADaqtae1Q4Ufflh4uGJwJoiyRdFqWLH4ujqW34
Vn6d3Pr+gtblhbGlgHlBwI7gU1SZ5e3iECJF5Wclc/H2Ir8E585Z8Mzmp/xH
nRAIDDhdbQulNQmtfGQyv9vkiiM3kYtXOwTnRWfGuR1grV6ge7CyfSVzqNqy
kcf+eaaQLZQDmGCgl05SpykOPMYyG+u7eshH/9Z7pR1D5cn/BHLzSfdSoQRa
AHNuUXJ3oJpBaI2+tT+QcaRGDdv8/vMj5u5eboTIlfZiGSxG7Bkr97vaNFBL
UhgL57LiN4mQlnYWGG5b6siwHj4Jxiqxa6Ef68U64jQyp8D7UY1QT5fjDqXV
oRAfuCu1idTflYzNUBnAbfv3AywcIRWE8cDJO64BbVpXqCo7z0srushNOoJY
A7XgdJOu0EXgcn0ccbP6RKYu9TEl0X0MKe6ZxZeHFCYXwWZ0SEufTHVHYYF7
KIIU6fJw3wkpMzFSR7mzFFfzwuP/rbdOQrhO3i+crI6nttqkpdSHnMVbBFs9
OnWnKyA5NUgUEMiCBXo5V9CT61Nt/iXRzaM0FeROV9fYB/cNPqXb4VBftQGK
3/lanIm+4iXQONuywcnHbuBCn23K+qkQtmROTiJ0BXa6t66DxsMLO/mLC1HF
aMrJR+1rrrCqEdmR8Edoye7Xhdlt61iFauKSunMDjjTK22uH4QPjJRSpTG1D
mjhQCnKmXm44+ITrQfmSI3ts6p9cGcnq2h1cJ2KzF/2iUOQIJZ6MewylMTaZ
KMLuYY7be+U8lmHCVOZXE6xHHzbfgfAPrS2GxSMsw0torFLNKkl54vlESFfN
plKXhAlRVfiluwfQT+sxdt2rdJ9eAvhBhm4zvEtLzjwS95xOFEjnJLigJUb9
OKWDtbZE8/hrPYmTCvUrX22EzGtwntFF3duVWHIM8SXoTj+ttCRRFCwn/YSL
srorBFfi5cUx7XdvzdeFtA+gtfGdOx8oLFHHblxH81U/k8w6Doo5CcdxrRVS
YtUkil2L6w0ovRGRCclCVtF6kSArh5pMyZO/sG6rkTM9yCn1dtsy7+oxG9lE
cUaPkSPK3EqkTp6P3W0LhhTrA+kVWKZq5BP0V5j+4c597duMNz5bEjNDQMB5
6tR56YC3DQVjhzwRl3U+fFsCAdp7vQRyZ/G6CyoeAOhJRYs6HvVHb3ad5dO3
I3vfSEoga+mBCIZYEBZEcTG6mmGK29ouEQFxDNCQymZ4Lijvil2WOM2/b2bz
y7Uq6AJSezSp932Y7kqZg42PAhkMnLRCmcTJ/OT4iyn1ZUSbUrFJq0BvSXbd
AP15DSYeKAzmL/jubqnF2OBiswu5uHsiOUXlKyh8ZzurscVV+BAe3B1egEBX
/JOVnD6dbGnHh+lDsnhUDL4Cr89sDek0KeWbOrPp56sG/N+kJR7pjSRkobep
alNQpbO+m/gEWfqsP7cMNK5JIiF+jV4gYAu9DhxCT9IaFCetEsTYtmzhxnW3
tCqccd2WMqWMigzkceEbMUpDVbsVMt+01KGgXiYKhts1vGkkmD5E4kqU5NUa
LHWflWO2AQEpefmaVYkzIV4rIAX2qmbVyEQ4L91cbk81oGqVR91fvpNnWXfi
QX2wQU7ycUzvO8/VE8HVjQjuQx6HIBjmw0geGF60+Cs3woDP1TWNM+iPFaRR
VLvc62gVTgv2I/TJuVS6az/lORxqVjIO5rwbk8cythFUIQGq+Asa6XC77tAn
wN5myckj44YPandVkv9DvII2Nma4wN2bRl/D6LLrWG9gKU7knLgNcmru18+j
0Q1HOWk1XLU5zIYwX4+4d6SrxBhoeZv/RdQg0GBItfunYGU+MU9elfOHZgF4
K8CeigbOu/ESlq0lj1MZ7Zci1DOGxvJ7avUPMV/V9wKLykyDuruZL5GA7ISs
6vMxMhcm6CyIf/4cNbxs3hZ3bnh86riHVzoHjwHhof/vWf2U/LL/eM2mzFAD
lvHOIev6RKKNHAxTyecPFE977n3FD20EiSKR16hfkWV9bd1upeHi/GYN69SY
Ylvw4SabzohBLmabMsiyInUs1otY3I6hFbS3OFXkKYV/nqn5lSksQUCAUzsq
x/jNGBUgjasqKpw/UWpKIjtNYs0GDiksiPj3VZphPzujIMz8XcuTMmOjO7Xq
DdD9OAiQzdLxkVlbGrQMHq0fRaoKiDlh97dib7VwWylmBbRWaWnX4wnlyC/K
gx/3qTZy+Q8ngfqDjWrIndLJJ0dguGwKv5zKSfCw7gBzycVmKzm/X5LnootG
lUJ8fAyQLo0nOcg7G9YaTr1ue7oinlWq9XGqDwIbEQEB7Qik1s98+bxkoig4
CBF2uJg5ltO/Jpsy5tzwMrCoKn62PcvXs+C+6ScSnuX7wQhkaQoYBDhYtpSa
doV+dTDO8i0+SBVhCTFpzwmzEAXWQGnhWuW9b/Gd4KQqi61Scy2xG18hCp1+
dKdKsCl526paZbLE4/94VZqH87UbBZeTynPo7m7Y2papaAm9EblvC2UBdrpv
X/GDH6ZA479lgmVRJpsKJms1IY/XOlsSmFw22Ki7++ZAQ+EoVYUhUxlqtlbB
HynEB3Klr4opnPpjcksxBzz6n1NPZwasc+++9gzqd7ipxGpD4SZTw3/UjjRA
9N7L9w7nbqlepP/rue/sWwZ/wcmGYqfYDJlftFp4r8QQ1eBb+0nTBdhKCCXL
Y6Vqqy3l9sI5o1EEisY6ksQ9IpA/4XzBucDHo8iFw5X1fYbynR/vIesqT/8F
zmdgJgfcAnisRl/z2uB5FEggaeNCWkVLy2fzbYpEywwdsmzHj3fC8hq6mXT6
zWYSIkcsjOt9odp9JrTFSAmt0upvgx3BnV1zGRmkr2/9zApG5tpznoHtzo1d
FPyjdj7Yn5kOqd+3vhWjgtpXE2moH7zMuHgcBVXjvF4nc5ad7liW2SrM9Vep
8xzVo9+iQIQ+d3xb5tZjSQkL0a6PDZ9lcPzQqaOpMZTGbBw64/vuJmTjTlq2
t92KaF9sRQK2x87PcRQYk5yKhxYtqpOyTM1ohcdusJ9XZshCMrHXNepqc9yH
ZhEHmrt0xBCvV8Fwartv3lTsBnSBX/MNFI1MqxF9KTghHFlVLaHkRlw6FWe+
+Q8u3dfEWHgh7TVdM3jZNWxgzpWOT6diQ4iG3E2HBJfqg7m3zqLjOT6jyt3O
U6pyKy/WLvcEaTS0HA7NLcvhThGETho6/nEIoVjajfsGOwCqR5/0Zdmr/Npj
GT3ZUtNeLXyQZUeJUFjpv3M+Jw7g3JgU1+ur+vVvCwOzcHS9vaz3k7zlmZrT
dYqJPMG65r7ZBwzMHsSNyZM6PbjEsUxcGQEMp1UzIZM3DROWFpxolZ2gweKF
5BDA/MYNaENlpHQnyp33I0tM1ulXEelZxKe4u6nGB7V13V4kGlSpbFMICMtZ
Yp17iiReyFiFESatWSoHufAOCpYZQ10Me9qfb+mILl+qziUr3zwpbwaOowQj
UnwpRp/nO8ou8nviNbX23Z76YN4JfKOcs/PHLglFe1dZr/ls4jMTqQetVCo+
stlKl8DEY4RQ95V/1w7RrFoPh44BtSdUgVpEUuHLZ5Ow+3usaYic2LgQhFLY
qLsmizN15ljBbGBoQj+NhbjitDN5uxYyzC+dAM5T75G2XwMBGjkvvV5DeI7Z
U1kzDxj4KTUooru7lG5amikM8nVjL/tmPiEo47uV6cHYKtur3vW0uhVNur91
Qn1dTr/tbrzczGasJbuJVLbgvDP6qYnDofEIN6PftxgPOqDEqMpciaJFHP5j
e+aO6JbA7MC0ytDFDr83Q77ecs3VRcyAvCRJR1StMe+/k4ex+0S+TrbXVnHV
XcVjKSHwn+FEpSPkqksuN/ShsKf1f/aaoBmV0ViEVoQiTYMVLy9Vr7b/T2M2
7UJqNa2yejdSJlNRyR2UwMFyYLaYEdoV8Rlk+9KIWFLUc0TkEQJIZvIiUctZ
ow0Mer5/ZdFpXXSzsk/4rF6NDe+RjpVJBpbaHA1VQPQjo7/t0zo72rQEb6h+
MBe+OqPzsygWQU1hzFO8ZNSELShkVSLTJwYVx/Ylxx+WvbZje8L8YlEYkxzv
hqff7K7shGkWuJSC92xvS1GTNqthfH8yys58VtR2dXc3XFnJoCFMT/c5LkOx
hOG0WjiGGxk6hr98MsQXUQ6jMvgV/Fni64xbxDiAA0sUJEwJ20NHiQOYESZO
pFIuyOXP7xnGuBQkrFrVl0pgZqYJHYjGRmH2QXK7yyRCOo6QeobqxrdeIUBe
L4QBiDxEXs6xYnQoYP6SWRRsZJbGACxTWaHxL6EpdfsD4WFdHD56mCo+6rZ9
zKIMKlW5MC2nHXYrR3iiQEuEjUprdCzkSoe2qiSy/2DP4XE7MaIsZs8ypgKA
GROZ9w1lWR2hb9Te2fpHv8T/gyGKoJELQgbTUREIGOZTejU84OF9yIRv2Hl2
/1J0tYAPeswOanzvx9G2MXk9m7FcXhaKLz6elP7fiDbWI+SLivDG49ARQu/I
I9rUecofJ5Bvcw8jMAqF3dCJbtICaD50nB45xBWRG3sGMf2k2v0bqHpewZsV
ZM+nZ0G4WAGGZwpecahIRqizDFHIJ2AH4JtR30HJb82w2B4Rgq6u6GX4YnzM
mZ52dyVHAHru7GrG8Pg6t3mgGzBSOwC4NJoqW8b0WMVAviGrEZv4YZZZ3uxh
C7oIPBB7N3qUTwYBIajUZL7YyAnBm2s30ST3mH5+2EPGX3x3+u0kEkb3H8z9
0ZkCvQzK0/Qg2dTkUNJc1SsdWpmfzVdqEJFhkPRy7Q6RRdakmHb/GfjFW2A4
5fADpqO4Gp6evBOoh4RALMSnpNUbFTXxEuTe++qsRNxc6/WPgaHxZBp1uZTB
ouAT/LrCLz1SlNJBi10Kj6+FUccb/0s1sHKKG8fv2CIx45IDv6FNgtWC05Vz
FDC4+0+MeUcIFkQ2r4jOuK0oF5omyh4Lyc0iGztiNFo4C2nvxQIiXyR1QqgM
XAtnDEeeolZoUOsDcWWKcp7gmhSm5ecnM/zo1/2CGtaLPdndNryFN9wOsm9m
pTkBGhMEMgnxEXPT9TA1wTOYwPddA3uhL8N5EjyVuzxVTw3kDgcUzGdkfkE8
5poXjgbW3xCOCjVpa9fahy3ApnWVUZXhaST+Y91msEj5DGdKK2vqd2P9gSdy
lDOx5nHwsE85cXOuc0RJBW7R4iHMB37zIR8N5yQOqV012oCpJVuhHxc5TjCG
Vz/0YMLYCo/z2oyQlane3ULoUX4r5o9tlZgkJFp9R/uH23AzLC2QEGNqNPat
8YMk9M6fouIu2xtW0pccdnmRt94u51G52P8dGlHpyxJitcxtfGhAuVVyaEOG
rJ00yAr2/A/tirhGGrCh4z9XJ9C1avjkN4vWw3RRYU5wWWYzM83R+5QwOaPW
FsEPfHAbYx+rGMVOl6hWUNXV3hP8si8SHitbXn1NswTLL0w11wQmXtE9v7cq
OBrAbHT8Fohyvrf7j7Q3pHTMPj3REoJCslbqPfvKIq7e4K532EPQd8H0goBD
dVE0qL0GDDhvifOQyh9OaFsyKD0rYSKm52fVyIo3Uo5VPSO62Tio8oSG6c/2
/raYemVJVSit14ca7jZq20xAhbjcdSi36YwTQzotsuC6LP5zB3It+pbnZUQj
oDJGHYhjfZEMmoY5TIpwzFCipXH1mNJNYnLFOrFy+7retCVyBVx3EWVxQA4x
4yt7BBG0jmq1HS1GBcL+HS+pOtW0uxOM6+HmI4i3pmRfaaDl4Xgicp9gm9yX
uSamT+yxKbzVLc3rluY4FE9g2JYiHLrXpmoIr1dJOU+FNCc+KLZS7MOtDgeL
zrC1xW5Su4km+NFQmNx90dM9PeaoFvogd5aSu3UHBecy2mrIgam5hVPErmeZ
QP8ONoSf1cVBoFr3K5anQ6UlgCNtViwWCHnWChymByARS3xzVY4J7lM5xrDR
K7gt6IQaLEd9kKTicqgLullNh7rirPfU36t0ByjrY4C2CghpSLnLKuYI2Snd
CQK50P6l3CVq8GYjJ/u0+PBXnKMr1xsgM9H77rL71+eTia669KVod/NZ/4Rn
OsxM7tnHvxBHJySZftwM832ND9K14kglRCiqkOn7RIiX3Aw8dSTdFM1G011Z
+LhEmtyEWaHSYnplSUM8QJe1tRlERl+Y5n8r+h2AAqvU/rXuuT31ZARtmENN
fR4nQ0ox1xmJtt06yszf2UYQTu868CeBN98qH1fya6bCNSPGTAdawJWSLwqd
Zw0q9HE8twHseMm8VC4L6p01cDzfA6RFn4/6ox2XKGG5Gh18BsChVYdPipSn
vifFPKhunl8juBlM87COa1Gel3MQie5wfNEajRcg98u089yT/XEKAfImKGI8
w50FfrCXu84L1el6tTTLAc94qh6T6vxc0JZsqC5FebGNLA8WfYIk6e/iNj8h
21IdsZBFIY93+28jXSichJaM0CC0dfham+qzg/F0uupQKNkU5+O1IWwPXVph
uEPEq2xrT1N2AKDnxDj5nOocIru0j10Wmt2WYulFOTWGrv+kk54/j4104Lla
QFd+iBkmYGYT19rSJQZPhmNk193UHuc/DW6OLy+qfA4YvGyn6H0UHXVY/adM
y3x+ZpUy8QaC5vEfVJ1echFOyQAXiFUY/CsPNqsQZhMIAyZM1/uWcb0Js+Mk
P783W6i+X0s+hU6yYWYFN+f1GjFal6FSwOvWosc2sOZsUzP/zRsm1/0EukSx
RGrTVps9I4rEUQ6wJ5KCQO+d4NkO7Ty2+RyEo03AizBP+sfkWg4HGhEWVyMy
sTz6fXCyFrlijTfQZdl4zUvpnaQZ1qGEhTmK975u5Q7N3lfcy0zG0Nvn0nZk
i4JfMDjq5aCD2roY/FMibvbx2Ym7mLyeDJzJ2lgFI4xgBzSLZuyfUahMetXF
/E5/Bn8TgrvpuHxvjyfwRb6bMc0ykwjz0PYLH2g2YUApnPyU2FzSae29D98J
FgXObV5mOjjnhXu2VmGJkMKfoOgBjsoPRtpY6RXdWlYAAJYaedRWKWJ1FmyB
lx42ZmR1Cob2e1LmCLlLvQM4S4J27HNZVS643DjfGTgxIBS6e08MqwRxK2s9
zhUBcjiMAf/tPqTLP+Rvs/hV9XHjDZu7N3XikCfL3Z3YM79EghGeS1k8lbFb
UvgBN61yUJBcR6NDfB8kzxFQLUyiEs1DsmBxUJCCbpYFSwDbsCcUGv3DzfMv
q7eo2i80gz1CpMLjYpm05wYDK6aRqaNlTNLbSEohNJ9NE/nT7DteC7yHolXf
oBxWMBr64vy1qvVuFMD78EljY5vhGdqwoyhn3SJo6CPZ1Z103uyQdb0MhDgY
ExQ3JyGDhTmeGAKZzD0ipqi9RijfF2KoVRTHd0pPZx/0CuwW9r2Kb0ObCI9M
yy9r+r6YSzQpj1FCPfteyxb/9lt29EBXijF8CvUVXGy/QWcuLwiBJBna/3Te
dwEeR9ZC1cbkRf3hyJ0xE0Tlu9hYGc/bxtu1xpYxIy82sBxBcaCL1hKtTwx7
aijXdDC5lnuv//QUtgEEFGsoYYdEqr3t4a+BhSTsS7T35u3ktd0ep7AMKhVg
E9g9Y9x0s3FVyZ0A+88IacwzwoulAGmMeQKdZSOuObQ0v76jyr6OzWZb3vFF
iirqA3lTfETIY9z2Khe+99AosKgLLY1vH/aDY3xMT7Bkp+GgOb9nSx3c91Qd
JBI8mvPgmcn+F9d23V1mcnChMQQYwgYpDlEUGjfhg2jDaqLnzmPYJnw4ufue
OIXEXgVnVZXsEcLdFa57YBay910VCjNYq1stIqTnJozU7OnAj1al1o4ir2Ln
2o0jtqU0Sr2yR5/+TOJElgi+0pqfdMZDIrFU84uBgR69NYhJBssPTeja8p5k
0LxBSn8ikFMIT8y6LXGV7rQiZ7OdulC+nobeo1v3T5W0aB2CguBRTpf0vCyE
ePeU+aYl7mvAWgqDkj/OQPETsjeAVRHe+fdTCukmXCWOxAZ1bGHsaRxEIo4Y
3DSrI3kmKamiAHjAdKxNy3hgGzatMzNZyMFuNEaGCv2fKFDrByMVe/92sOZe
Nrk0zoYUAmfugLSCJAzQxlDB7pmKyPEuhiyPX+UyfL/7QrLuZB0IcAPTiyrh
jn11VAxFeytr/4AiXHzyxhssGCfrfaHpmudX7NFkpinMx4PrA9+zOzSV+CFT
C9SjWrdLhJFMtAt/RaQO+6qddtXKPeTplz/sZ5BQV0TsYHEzbNg2lnVjXVOq
yo/GH3fMWPliHl5Y3Nzmwg6ZXE72bR5ySbUGktKWFBu31L3GU1iwBPgSB8X/
AFDMnPi3ECeI0TcYR2jsgDAkqv8rs0/wxC4H8N1M/66vJzrW0+qkubtgJ0I9
hyFvgoD3w07M8DUrkARedH8g5f1tNazdEq0PFkhx0HiyMub53RA8NN8CDYRA
JAGlqkLuV0iv8rP3dkwJ3xlnRTyen/qdCj1zYh5dGlYog+fhwUg0KKcK5Lo7
w2tE7NlrGGNOesdKp98wz4wEeVP3yYuh3Uy8U7IvzVBTXpt/H03++H/oMH20
TMqoagtmoXZybAMciDuD0fgONe11EWNTGBhgUYMUQu5KfAbN/Y506/3mKXIQ
62/QF2i/sfEwQCRtHX+YFTW+cPfskUvoGs2zqbLh0HflLgznyVlPunewEiQd
vvOD6oe2UILOPuhOQ58xrdwWMdz4lPGfpCiLlRqlj0pqrO/u99cQDevk58Ch
UXKab92gdOIiWuBCfa62wUInaz3P9M1wCf6NbQHh0ktlqKGdBTcWqaIrM7jH
e6jpF6tsx4A5OwS15Afym3MTcBgc+Nh/KAtYC/POar6LrM5ikIdJf6ncKue3
DvqLaLU8rvhLXNcAZ2C8ER97fhLSEIO9GSJjGMagjXZXS7jndLDZMr7troM8
cGCAfcamWPL+++NoZl+Fg++VXPm9ewP5xctyu9EAiXhv42PKNeyO1E+uUGOV
sTLRhB6BmNbYPZTBarmwklrUpKen+Rd40fvavu4Mg1P8YEQJIopgyz0tNfXM
ACRc2WldJTRa0nsdIL0PPUB1/AFJihxnuVAG3MB0NTvQANmJ3x1o9BLF8GSv
TrSo1ZoWdSMZB7Ak11itlQMnbMJ2ptEEK/F696ysK474OCoo7hAcaK6D8oQc
jRFRY8hoB5lApMP2WP4fXy4WED9eZ9oflRVKlJ9tVL6q7z9q9Y9YTSgxhnMX
3ji24nR1hlQB6TGMD8Y3p27jr9h5QFVZnEIbnufqD0xr5M55FuEVBTBBSo5b
0ub0s8At/76RdQI1aOtRkhGk7XtsIn4RCj8xGGs64SszOJ6ciOR6JFNdJc3E
cVjf4pC5a7fyQBlOUlEwlHsruh3NCq5FmE8Z6Ca9f04mPRteUjeRVNe2Nv5F
ZQTrfz9ljXqvCgWs39Ep8LlzUx5KV5kdnENC6y7Nkpl9OO3hgNv7pDY0I5mP
jx6gthAEZiB/oA+0NPayPvgBDl2bT1oQsjrEa9AoArSX83orZsTK3GDi0PtI
QpC4Mvfl8JzFEoLJ9dWRzw729cUL+1f3Jkql/He/fa1cF7vDREpBZ8cAAwOz
hQNJMFfe8/o6bV2LqK13MPTGpZFslrGG2IvPCkIgyDS7X4cACD3n8mU3DdTC
YsVSo3hg2eidcpQ6tYoeA4DSt92c1kcuY72eoea8700QxURuULldTD1/t94k
UUnJaDfrpRupjepisGkCR8kfppMs68dGmV0pGB5PWMf/+Fb57chADnxJZ9Tx
wd9cFgZyQA+9SCjzn3gX5xHjzW23mRhGxqcshcBEfhrFLezmeFMpBQ7wNKxV
ITzar08NA2rtG/JnmHbLFwD1YfLy4gjEO21/k5paDSAcWpkPF2ynlZ8VGZuI
3cDmOFr89WtHKMGYqQx1ugu/8P6qlPa/RJCBvexJN3O/z/1rJ4ioVh7zpYM1
g50lSsyAm0yU/zifBMLp+7svLyu9zTGmmbFL/wfHC0yv0KmNt3qusDObRIBi
BYESpt9lSJQuNiXzxVPuS/+DdHh4z435sgr6Kp+3+oI4WBaAzm1ph275CTIQ
+2+omyBMpteExQT9fHHiCrw6qO4JJDbupA77Jj9ZXtI0yGMkJvP5DYH4Qr8/
RLnYjpbZk/bM0E3fbOz4SWpBg0ppO+VH8GYLxB9lRDa3bhkdDwPVzgVp6Qop
13WtLeoQNu5GuYEUb5CNhMlQmE7qtqvvloyqaSjezfwR0DGAjY2z/KFwrYhJ
RCEM6/yuWmL515IRFZvVTGv9dO3SaRHahmLXVRKCzefHLZnYnXEi7YdV/7aq
EWSQLqCSZN5okV5rnOWXSM1e10LVGlvOV7uccuoAmFfsp2NSYTgjcEvKJSWT
Ys3q3qu8ED5W3OFJvscjhzPkwrIKK3xlG+at2B71WYzM63iqnbRw2d5xcG3y
5V60JsHLfYG721HrT4fgQA2FX+ubbvwGmQdGqpvBJjvZ7UE0TpVzroHzcAuf
DfD6m6u3yE6vOFmWoiI3mk9sI9JjEttU0gXmyhhjyBsTquslutVxcOG6i9LR
nZlXDiZwv5VEyy/en13Jyjj+xvB4x3Mm/LyCV+UqW5pevehssedGzp2DpuAa
XV6Rztpx3QzrAzkig3YMgoEYpK/MlXlKQs4681vkpgUOc7pJm53KMm/PgCEp
mOzkZRPyw4AVzOVqRMlRjFu3HjiDt4LSSY47kbQyqkxNGBFJfHz/VFlqDpxm
6VzdIgcel29jkRtuTZbgn7S9VuTFVkLyIZQ/0GFIeMatm5Rf9wQTtzOpTRdq
oAUwo4eNz36dt/aufkL1GZa5ikHSHo3jYaRfCDCGTWkL0+f7ICSL0y5URkSA
kWR3lieaUHpJG50JEftV31blTDy9mz1l13EH6PkaU3Ja6fnSGLuOSIOmaobt
jgPjRCWDc701njxMS4bHQaArlNNIVkobMiaID1c6Jet5dtFBrr/XU/j3pezL
tpd0tolhlYEawj8fAL2D3kY8aSeHCAJklHFW5nkyWHuVAwnqdM64Hk2WIH6f
WfYhGuINCmWGhU+oWC9o1iswLuxdI1AUrtB2fQd30bRphEL9rWvy2jfQMoF2
/RW7YxxHvSb/AsgC1K0akSraUZmymUIQSxP0Doi1Q5w6nRdlAnvrf9DosGpU
dbLuFCzI/KcA3+fUbfrw964I6o9CUegWQHUORqSu6i9w/S1VNfPQH6CNm8w7
F4nSuX86mSKuzat8JCJuFUBbaj9F4fr3i9AFcDUoSqdh4+2dDrtv+yLsH5bd
KJqoEjdA7z+hvznQFaP3lzVYMWqvasW8RkS9wCarWEymEWghdel6SgpWB76d
ikuEKhb46SGIwTzrSehjTaFv+qmSJ/zLILPnjKt/WtTEmsxp5uq31NpMJr4e
kWbNJ3A4qRAdO1F/UCZXBNJlujBnbC/7e3oRqz0oS0yMPnngMsioGnIDug6+
11yzLAUC2y/noZYnMtIg/aEf9GTVc8T9PmbdYyMQVAd8Vh0KJkwmWDA2o4u5
j7lspwxp9uLGsJY84Hw3xTihSz4NZMeSFPvjZXSxp9COzQ1pclwP/acYzuSU
LwGfPXoYZmpiKe+b+iTXpvzfXi94fezJBNszuMcD91dgsq1NxSuPwZXtFUs9
i4MP58LYtBO825rmiXeDTZfjivOG01RqyqiouF9YvDEJE5zthBAHQr8D6eh+
AGhaZ7F+RtJHFRQBm1IMzBAw4avUCna/EvYLiFbLs0QM7N3ju8bMYDmlyPNx
kDEz/xOyDC5z0yq7T1z9XwCrOTyhwNw8KWLr+hvz7//VpRgG8iA642jbROed
wPiy2avFAS9RBHHBaSf/2AT0P5WScQcjWuPPBNtuTNoLyhLdu2TNj5orhdL7
apfPzKqiJViNQeuSaUq9XGm3cYn8QWXH13blkzSTv56xQrPmMyIfQfl1oJnO
zEkffiNKLJorBp+DJVJKLsUHtjElMBDPMM7rp+t2rE+u2YKU1YsTFLTPN7IE
07Me/roRccYBj9D4tqnHZ6jWQdevjFd+Cn3lELcgKWr2sE3YK1kV+mz2yrgl
aQ4eDVokrYJRXGqXYXaZlTZhGkNOw0baR+TvyTv855ou9HeeHIaFBv4OoQlQ
q5JQ/Tl7Hc25g9By8G1o9nQRtbZVpcwTIWQdgzgOSW0vqbuKNG1+Ywy8XwSZ
roNI5Z7PbbLjnfFNDuiBN5zW+aK/0ycIsHE4uWhJZrjomz6fvo8cyswsbFQb
8Mtnc+IJZVsJLBcZZybLrDt9k55z5uODGI2tIJQNjFPTHaE4xwK7O9tcogB5
NxNllXbLljtRAi6aQZsZG0nCoxUKrVKi5ylfs5fWan7fU4F2pMpbfODKWkTm
bE0M1NJx0czgPDV5nzEbI59RKSxufnktLdTAPmk1csra0YwyI80jxd9Sfwcj
5oxUDPqSiBIe1DA6qJy2f0bhuaKtmaXsCLe1lL7kapeCwGiKQWHg/lvtHiCu
mftuRYmvIhC4hC80dbV8wz8Qq/XAelETrUoNDXfFqpz6hiyl4Z54ym/me+VN
MxsuI9G+wzmjcFcW3mnotVVkk9bBC0N2MbyZFfW8F0bBUzBwvuDl5g1Ge0gD
+AtWsp+CVR0u9hFDIgQKPmr+dULHSiu2Ru3XojUG6xg6g6UOkxUpsxxxX4eP
jHYVaxwmQlCyFbEqcFrsnd+psIwZ2EzePxct/nZF51Jauy8TcpT7LD3O0py0
KzZG6CopVQq/PjpXJP+EurGFwwLev3g9UUahWSdi9InZ5ifXp7GMmsuAqvqg
Jcf0hJDK4qITCnEHt/iNZyLfj7hvX81mxEfPZOT5phuC7VhA3kA8GsDwJu2y
Ic5X/TcQrVB4myxoL7aEMg5VDpkcmfznmBWdLJIbRDcvveX3vCQN5/03WgaI
t/erl6hJyyDsgcue0N+bcQugROy1oDDvytidi5IZ7Hzm5J927Y0IUeTGj45V
pgiy0FPKxqe8pMJfbWcutoQTFucHcfCbP1xOF+7sV4XfHG5gJiKmGidPsUeK
Lgvs1v5Y/r05NP9jZsr9lbNHH6TYa4879xYtRIduGJm9bjqCVaGX74cN+RIs
O1ZtBbaj1bwntwXzv8EzaQIkfyftuccaYi8Pi+STDZegUtvGmD1G6+sEh7nw
6NgHCkQomY4Y6Plcbr9cI8qmp6kLcOQssvc7CehDV39tEjrTku+Zda+r5RcM
7oNs9Zf8taKXrDwuov6+h5K0sxjUh66eIdDlm5nsz7bTAwpYRiB8Y0xf1+hl
y3xwSm3sZXFvrHD4BxQsPVWFywskjwmJh78YWsdBxhlHN3r3z2+W3sbpk5Pf
MFGMu6uyoodaPROSXJbacYeTCHxR6NlZDp1zVGYVXPoewitABypSVc5yybwN
y3/kdTYU01LcJQNfFD/n76DPxuLGdXctkJa+EVeCgTf7rXusVTiN1yMMILLk
itTfI0Co6a69Ix8dCI8QeQk4fAYfBaZSUrJTcYW2npem/Az+LHdz6ZfLzkCq
YMulB98X1tNj4Cnehc/8PlOyA0HzIawsTgod6BnPXlP3sraICagfVsX/skX9
k0pvvUbH6j73K8jCMSM+pAeqqxAi/WATddPu1xOOQX42DTsGskamVoyIPhzL
XzW1PGTm850bESF7ACxaRWvHSjH/NxXSxnued9hwxDne+YaJZKtxkX2JXSZ+
AHlS0CqL645afaIOqKPo+4svq2+wwvp2VxbT3IZCWwaV0DPvaMU+zVKZqZBG
s4+3uvDzoWL0Be0Sfa56dX/zbisZrtAbWCTHpS6yAjjmkAOdCqL/YcXPDSLF
vqxwFdtCz0yw0P3Ot5s92okGOOHjK0ZfBN/7xoLfhoyFKh/7xFFqJdQ/ZRMV
Mn4a/MK68DlnwUrJcHjeL/DFllNqnS1EYApUQA8A0U063etYH7YV6QBor/oH
eCRvRlxM9LepF0gVgAVerkb6N6lsseh0fQCSg5OLiu8nlj64ag2kd+VKQXzK
z3DydH9Z4PTnQ0nmsJJkUO8qIs9y79nTzIHoDD4BvYigWT6elw2jLbkLTwvh
tOJp//egC/US7js0NJHLMdwG2T1Giu0VrsVvPIrZrIDP156LdzCPoir8ndtC
eMmNklpjp+DhjnF/GNPiMPkf6LzRobMIopkrwDOfqdu4QxwYs6a/XBhzXPo4
wB1j5xATdB9bcQpm/5GH7nXYCNyXqYNHe6d6LPD2t89jOsxw0MV7OGA9XvN1
zdHaY8cF6m8VrJ6NpPA6k11CjU6gY/TOAteBZPE1S96QIpvZhAevC0oLsic7
/JlI0mMRiiRArVdxFDbDwH1UH66wtVFO21daDF7hWd0XbuSDsUOtpNVJXCWX
ewlEmexbElQCmQ3M/H0OetCSy8vMpcMpm3hZARBFc4ItPPA5edBSc4vdi/Fs
6mLtosHbdwHbvxtZMbOHl1imWFgfTxhJ9eOMDJtDHMLhZAnKtBMFKhegXTJE
YYlWZRbRGc8VHqha5o9Rl4ZG1B2MoPQ8ISExUsWZ2V8KYQkNbuiJUvZURDXh
BvJJVtoxvEFikbQvT0CVQvEQCqxRt25vV+NU0RfFnqoQJQLUPSGo2h8k7UHF
S6AUcvEHi6Aqwv+dzUM5AKHWILgqkP1IMdktiu5trR0iIncrOK6YmIeZSzux
BDXJ/qwDKLGREErPyYkOD1PEhR+2JR6KXtufUDGFHbeI/p2sH+YQDcNAgeLD
okci72tEhpkuvva/CpBp4JmWv7Nnj8lyppJ6SbFW7nerML8ZPFP7Cq+/0vzp
wISGixL8UG2dCuWYwcJyldHRiEupxK/F+kfhaLgWw0wVyXqDfD9aIeyWjKa2
4IWmnG6CHp+HSHRZBt/3gEu6p/KhCpSVGoaNfx0fW6pZ2w4B/jal1vO3tlJr
ZzcTgKssfGx/zyrzdBnwo1gXNKxHKjkfj89Nh606nwdTmyuWDDKP5y4opAEO
q2TVM5Yqh3Qz+BiGWIBkOL+wfvXAZu98ygfMVq6QDi0r63ApYyMDSOVp7Hq7
doUYBt0dFKuQQhr2+Kk5D1SmTUBcEMcCIxDgOa7Q4ckdlyY/TQoPiW5AUogG
lONPh5axw7Vhxsh2lthLmMuSGTDVk+TQrCLJCMYzI0thJcJio5XA0F9H9C7+
WqOklN1g5bYtWcBU1fpNjC4NvpyEX47/jE8xsRlTMY3AJ0Rxd2FArgit3I0b
1Q3tN+EcPIR6uFTv973sbA3j9EZmRp76LptwoEs9pJnoh2Z3+FTAXooo0bLy
laUtxVcVzdK4yQyoXFQ6/4wxSNpYRvl45MOHNViMiOhJu6s6ALfX3rFgGz1f
Sb5p266zhwNW5jQ8ZLjYYeqLMzTMN8QeUKJW9Y29rZ+cQxGlMi7lrTCqiUiD
2BqyQ3llbSHSNCXn8G9e/minurCPg2DNDeAFP2VKANqXe4i7WlJgv8LyR1NW
q28kSCWYgsio0PShlpecsC++8yTS8ZhHNZ5UqZr7J/3/wXZdQQ8EGI9EaTfS
ohKLUuu4+eK1T/RPfmx00rgA1F0kiMfikPhPLdbv0gAIxJKspPdvbKUR7MUq
jMZ/2C2+zxi2uLZ/MOdS4A3zPH/TjGnFkrn205+g5CmSztHSW73jV78a+PSg
fG4nT+gcKlaVBnVGjtLYXJvEk+9lI7PGeMZK1D3ekYzu94ux3WqY6pjyBrdN
8yd1ReboqVzynD+rnwJY1+V8p9+wEfcNIfTtsWrxu/ihvTZCZsqBCAlRkVv7
enKJ/4KN1ySw/isLfCfnc1GvwgbA1+W2+3MAe+4gDzt/Qsig+pg8lRpkddr9
/Aq7F8LPCjHI+seCZm3p60idCYcuNyKCiVSMRtw+xi05tekhx5YhmwdvPjD1
mmr8aAtjbDJda4+98luOgaEgFTnKqyxsx/mxggROzhzVAlUfEGWF42ExcPYA
UZRE24IqRzSGhCJEuVcEgQjuSLpAuyWWxuYUEzNnNFkZ7qb/8LK1/xOYa5Ie
iZQFLzk9ZOQP53ebdj1CiCgdjMsBmbCxD9/K/t88NJsnFFvXAGiZ4KUOqk4u
wJa9UDjUQZaX12c3NiuAP9GIpOlRQ98XZivVTZpHjkyh71ltuZ3QWEVwqnIJ
uBDIeY5Sn5RDP0iJYG/oznbi2ZAmkXQyLY614D6c7kL6oxzJo0xhHjyr8h28
Zl85nQZCWiQw3sV1b+ewLmUNBsyW1r9tywIFJG257YCHvcKtRBLtgAx0Aqxj
0lXZsu7p4k1ryY8I0OHQcwVGT0okZzjcdSh1OIEu+P0ZqXuSDAYMbC4YAOkQ
yLMyjwJqaRq28eVvzEae216UxzmEOHxwSOwGj/sY32cXBbCCmo4quezDDX4f
jo0tKEfAaEGdpml4vbBGkmyFg9UYE16UlwClFd0iMFQIH2/rn2H9T03zY1vU
rM2AAVPXC32xl1NqtFu6TvOcyrjDHnpslr3NZZHukIIZraSiWIAhIp9AOKKs
zBhGFHreiAl7hoFdRFd8Un7FzG87X3H55MGLc8hyj1SPhC68dP2GJnDYL5NH
HOorC4TJBn5zPBEpPpI1G2E2n8uMh8gfTnufs+w5632IAYC0K1KY40c85CU4
kqr8/RjwlKcnWx3agzoeghvA/raNqUW6GFGaj733hmErz88ejKQY6sqh78f8
2qQX5eVvHFKi+Hmp9oBDRZeJl4yN5nrG1HYEJ/pbgkoKqSKEtQLMJ0jDlSxf
onJ3DXvhHqujCeYhuuhMVuZfLpzM967oJYvgWXbw7l8BV1dHl8RYTi9FaT1S
MnQreAr5VISNrlqgVlN0by45W1Ki9FHN+n0ACN9lGlVFM1PMdXb9g4etZEW8
jHUdXlPJEhArFTUI2ilLS+vmeBduK5PvJGweE6QhFs4YnCcBES5xvmV2N9G/
2d6U7lDuFJj3mZj6lOzRv1yQgvnoXNKKo1OlLxWlfgBC23V2SFZp2WsVMsSx
JPi7innebThROfan65ahwM8vgT7Sk4aXeSKLfNcqA6w8LTpM0LYpseldnMnA
UYrjrpJiVOXJ2ZvegXIkgjmiznx5fEOVVzUr8RX8nCwNsNZAEgGR/Br5K1zg
4zWhCmERAOnunhNruFy+t+tC+f1OFSYkRF/KaIoxiNb0z4F+gWA0Xn6tcfo8
mzFLmsfi1Y1AZaktzpfkbK0eVaYGxCCfHu4xxfcCjT/zCVMq7afZlkl0dUUt
cFrytzx/K77B5SVrIYgvT40v8n/JLWTkCcLQgPXyFiB25rq2yEeh0qzzqGpt
yT4bJ8+bHIF5Lfk/g6612pNmRgvJNs5HlQQTOl9WFi7VgNRxB5YpyUvbmWvF
5qBu7xbx3MxjCFCzfSFks189GWcibgITub81mmRA/9bDvMGpC5osmf7WDVq7
mj9anJdU5CpxzzeXz9brsPswve9KciykgrF47OnlP5XzrqiEHT2ILuZbVItx
hAYwsNkChsQFSFSnOWr3ofrKN8gYWIFFMawjeriqZ54RSkxCLYmvri5y9k4z
BR8ZYlMK1EtrlmpzBnrlV4zy/m9z0LwcMizYnKxXyfSrjnOjBk5a/0yXe3bJ
L61bEqZXjuW6kYOL21+Ye64MmlBG4MO6oN5ByKce0ZTbcFcssmPYk+TjeCOd
L4LKSIc9eT5rbd7sLVLWnqdFz2Xg22zpn4kKhQtXxGaRXWFmBHmrfbeMPSla
tv+c0KVqIGJh7jotFSLJu+FPXkUyyX3Y/6pHvV/wCqENBhyQeve2XVpvt9kQ
DjYTMbJ7tAWUrXrEX5NBgSYaHJAXXQIG0CnldyWGd8ELkHMrggLwpC5U7glO
fv+KwINw5BspxT6T6zGHPnrFBYxGQCwvmZPl8c5ba5LZ9FNxW1eUmDnuJ3u3
d4UrL7QdnET7HS3iAuOk6XG/UWOeH6p8uiXk+FHcR5O8WjeBHtRscWSBGbSt
UHcq25qV9YQGiqmMTN9ckmmBYXSSewAhFnOPHTN4kMGAIiYxsHLJU1YNaquT
SGIWkROiZWcw6suI5Us3czxfReV6qmxABjeWLax+ZOb4fVWQXQUyMCj/xZkB
9MI9n6vQh5X49q3B0k1QefcxKbk59GRxgNdfrVjt44qLjZcjgaU/WoXtztp7
wkVeT/AEIUzQ4QTYVEgRbhCAN1RAsa1KqjD0jAYfMcFIcY7Vi9hT0C7Yqd7X
gQRmD2Xcar/M7zPBrG++9+00bD5XmzHKiwohoQTcSPxB8dGxqjFRyp4jZVYz
PWuPf4+T8Z6ZlpOXog4ZPQnEa7GuSn2ysxQtcQ6h9p9Pk9eAydfrNQNI7V9L
z5j+f/uMP6/2f7eo7P5dXUDPAWIcbpGdtMfHk6D7Bmmh8RVNx7ZhZ1gBhgtu
4IzKps0MOtlEhQD1qiqX9GNVOE3z8IsS5w7Z0Q1iQ9hl0xuwrH6vPre9IWyB
U5BdMuifVdKTJkhqRI8KsM5LQh9bdW+ORgk0e8811u4eYALPaujRWOh/iwRv
TpphaEafXxw6YYLyZ4Ilq4DGFwkJban5kwqygprIbrJN2j+glbDAb3lYbwra
N1qA3eqxBE5EThTX3s3RKvMlsYG2NWi4stPuTL6bPL1wYoph12N5Bujo4pde
pXKBbGKz4nEjdk0BrOdE/q2e2oWx5WFCVt+OVl7bPwRH6nTJniS/Ivd4iF5K
kPcYVV52FFGkDmlrRdOazxBEfdDv6I+GXlx5GWvVDP2RfZhbLWxP9bRlyRzd
uwrkmRv65TclkAv8bM1z5HII7W0LVnlZ/P5Nxd6TUq3TJE33lB2ZiSiZ6YEu
m7pQG6GkdSr53NzDa9OLLqQayvcNEs25DDOe8a7/6sXJsQBumXU3Z3M56Cx0
qIL+DSC7QrPHj0i4ffhAizzLxrlBy5klB9xyZBSuSCECoEaC1tGpLEX2Rvl2
6LACaOZjjF+q2zMwvGBXWzeU78HR4YGtW0khd34h/wFguf7An6VkzAPLWxjp
sBiV3tyAXc8YzvGixohNYQui+fyu+4O2aWegRrJGaRCPCn1FB7gUFaIWzLwf
tw95ovRgIyMJYX8f60PE4nZqSD3iLLudI/T/GKWtme67+Pbu8C1hSJThFU0Z
I4pQFa0HJa0nnX8GQ14+t0xpYckFaLBDh5m2s/6k2+fj9B4hlCUfPhoINGun
YH+Ae5hmHaBZuRx6Ojydd2oQb9pT+B+KoAt51Cj5Ru807ySj2js5E2nYcJjk
/uyfwaN33vENZk0eySGa4dQG35puyylGEYAuyr3Z8YVaobIA21PeuStsWXrW
YSttMIW75fm1foiRvVC+7MBiT2H8mjnWHsaNQjWa1BwgWcfY7zMGUroefMmA
+MXsYHg3xAqv+cUJGaueynJ/i0DS9zvr0mZ+72I1jaq9qf6c7MVNiXlvPrIC
ohhW+Vzd7YvQPfTe+q6zhSk7wmOoIlT+zqD41EZntm8TqPDOsN58JEKnjm9V
LLSaBjkOJlKqGHhO4OKfJK9JdRYa5ZKysnw6mPZlK6d5u8HhkreWakVdRG7a
OG3tCqCY7WrfLpLbXUP3g/fDbmfKGRLztduJaA5lsY6THCnh9pE0rTnalTNA
SNM2S365dB9vU+P9gzYW7y3jDXUuGSgey7dZogl79zl4D8RjhJxMMw0b92GF
zFlnTML1OVH/9JOY9sK8fPs0arZesI8GZJDhDvcrGTS7sjGN+BbTfFwgzniJ
AcX63oyHza9N5fpp7iI9xI46YaaPp6jFII1OPhRMOReyZ4TCYHr2AuoxpGXp
PbBMg11TnvnAgAXe6AenBuVWOeFv5DgUUZ79PZ0oqySl3Nau4xQR2CtUdvIe
qBVRJaTnKjXkHm6JnevD+/WXlMavIFL5biN6S11nX4P+5baBSpPkfvASkLWW
LaoUqwJ2jyBC8cxEeMUQPXcxFeouwowK1/xkEe2tFMxnUzd7XpCWqj2WwgRt
Je1QluKNcyFyS/kkaLxBilaWqz6Hur8XlO4UvA/npYgcKogtNvG6/TVbn+m4
OBa/EnRuThrv+qfz6zepWy0JDhioDeCJoSDGzwUKpUEQg7/pzVxNdZAeIC4o
RPpGrvNBGySUA1oyovq+qCgFo05Xfp+qQHZIJMKE8MvDaSBhdCTWKZTeQJTR
/OmijdJ8qR3YngMSXMFDH3RQXcSVHZjTW/Xw7y1PWN5R3My1Wl0UzHI1HqWo
FsDHu4LtB3R91Wp380aDj82cSwa9kjlpBJdJOKzQ1LCBDwX7lH1RoaiLAJ/V
4/DhMMfTnQSEEvIOkgCpvPxdVsAmNTQgQ1j8bVEh+SVUtLCObl3kiZn0CHFA
BLNhwpTsy0XREeFbRWoeb+1Az0eaMsTDmrCZMtLgDYCnFDWPyCy1KEaDmPKn
J47TxOUJRq+GEKDyRj44W/+v9hPwKvxMtHleZ8lm83jiehwK22yAoscJZQmt
bkFRJlk4kWTNFrIOrMpQFtle3XrY+t/DFC4EAnag6jCvUXyIvEf/amGT3TEd
Vc3DMcoiX7dou0wh+v/x5bbUM8cclfmyXbqneLPs4CLIk3fjRd8Y8tVWVApR
qkIAM+JuG5A96jMIlt7nrUx7jBnh+62XuH07TJsyr36+lDdsKfAm4+XN+aOO
VsF1xZgK60OY+QACYfFWNf8vAxPPNkXct0BHHS88lfSWTqXLpXpCi9Wtk0dI
Q/VWEki+X75tf+RlCB1AZIBnBM+sZQnXgBSMpnkQL7Kul+rvLtTEW12kKnnn
ZOqIdC6eQs7PbV4odgfLgncXn+JUi0UTod/lvjjRMrgZvIrJCgscq5P3R7aH
5I6cFn4mudrZCH8vFfzZiMyu8jiNO2ecg8MqQo7GmrAJTzWlHTVteLny8d5G
CUku/eJOEZGYJ/lglm+ucjRQLkn+wjsKVhz8OT0jPbKWyngAnKNvlpWm/t7a
LsWvcHlF/A/Mf4yYzpn4kTyo/CcJIGpGunJMs4eOcnPBhvVJ7fXQkXT7B5SH
AGy1f+NUPc8nxNQUiBoa0N+zuQ7ba99+w7paJO4GKNrwJv8AmVjclb32pcRX
Uc/6Bi66pUNB+uXozjPgtnjRmHWORJWBzB6mqvSHmWwdaTRiG5Y57Dne/+dY
XC3fY6uOMFc4l9WVuMpVg4znLj/u09cVftKE2vV0Jq6hc5jN0VBXI9pK99EC
L97er+I/lr/6Uv6GEEqZxLtBraLZE/mY6W4/VwzoErtKe3eki49GkzRAkwFb
dsiX2Zsv2LgUIZeT6gUf8uio0RlgIYahYZXQDgqqo79RdGBFV/Lmnj3dE17U
nWauo5FezNfOYWrhXzQutsguXFErejsItB6OBNJiO19PTht2kEd6oy2qFJp7
5syI7pSA/BZfw/DGZQ+hJj6tB7gC7PIcDbxkP3joSKrV6wJh4oCRr5QlZBXs
fFvtSMJ1KlCnlqJ5623oyMNkABr78oGYrnaGXoh+zggKsX67C8IZxDEyNNbi
iW22y0UWxdQLSsZBj5HytTVxuTVRysh08ePpxcPe+ZJz3DV6CGx322lbGx9j
K39oW6PH7kf0Ytrmr+f3ieR3xQ6D44i8cOGlMz0i25K/4/iWoc7gY61PFZPE
MvuS49Ct6NANJ+fKwr008JNhqDs7E5ZfcQyCky0NzbWxVjIH0kkcuTED2wxP
3QuX9HuZwGNc1W2LLhyt8p76knBI5XvESBMO4jDVP1d4A+u2MtGwl7HiVkAh
FybIm39pUNBRxqYLfLRzWqJ3EtDopqDuwMubcy/NS6oWCbnxU6uu3osCkvJ0
xBOTikTuaALcSWshHIlD1ROy+R3wzxloQdsP5uRP+FOUK3ng+4qUEW/H0WVs
OCBdh4W/Umd6dJYK87dPQ+zhrnLubcbwCv6NEoy0Fyw6A8KsfDU/2j/35diW
9OS+dK2imekXUbbn4I04bYKBLsd4lOUGQ52y0LVEuVLM/MvA90WLkHBcUtRY
1AoFcnl+wSyUjShTMJNqH2uRfYvd1B75IgfIeno8xXQWML2o0mtzxN2T0UE/
l+jo9PIo0m9pg8ExwS2N6bjLWXtMKmzquwq268cQMiwoRslALvbQm/HRBRUq
nDxBiFXT3GfUZxvQKAYXBVEHxMb7xnRtV5NBECHCx3WsbImD31qALMFbrKhR
/tOnvt7fhYsEeOCdPfbSGNlfNHa0BO9NjexnsSQnfHWF6hEF5M0Q4u1PwMtg
YqeuYrt8zkpvpiiKIZpvfRNQ6YjqUSXNZZA4YYiPahdWF+pSSk89Y1Skt/iT
mRgbU6UezlPlvAu1O01XjO4Pci5EnLSC93hN/5fPUZ+v1JTSInAjJgoe7f0U
ksSCku7RvBLWIUl5V87ajBa55VFX3d2SiGMlsHhjBoR3SEJpCIh4P5yeWOfa
ELMmB0ph9GPhNOsapaPBp7SEpDzgfrB7yMIqBgXzhfAq377aKUD7wlGt1x2h
o1q64V67oTXdCJ5cHixyIeScJliBNDwUiGQN+VO0Xs/c8Z8tXlQ7przJAYvV
48MNJ+VeR53tz0V1y7Xxr+aQwhqI61V240rQDVQc45rsHvX4n6YM1uJr5Lse
H6/R4AfGVPQkbsZ0h5z/OQO0OfsyrvEuSjfXKANHqIwwQddE9xzS8843j9Fy
lqrtx2cd5MtFWpxhUVxQ56aIP0bUx2itW40n5tTyk9f9AtJRXS0zdHJ1zSxe
lz4fACTx+seY43KRSuWQp5BfxeLEdbxsCu1aokmqBDkJ6KpMR7puvrMxpfzW
oq4rHR+v4hAadAursKFZTqwjRj8N/1CZNpepdrwXIFB1TyqEXMbiMf4lmrhZ
+vZF+jrR/BIVl66cVZ5Gw5rQPEEVHm6GoxzMpR/ShpmUE2S66j0X+cMaIv6/
BB1NtvmvuFBlcJKr8NpUd3Dwl9yI8aMGXUvKD45R7RYS4xk0kxQn1zWHudmj
Vs74AMb//tzJ0zHzB5eIEmracsHSbRWhvQ6vfLC64gOBFX0Jb5FpevoAVWuO
fjdpE7WIDi9Fem5lkICuKlLt1LJtPwgBXSWgFrzvWsx8Yk243BVw7MJZ9CBI
phDD0QcSXDERyXMbbYXkiUTU1bPmH+tslN30Z6zSHRV9asAcyIKV7tv+//FM
Nt5xHE3e3YoWycAuKIWbQgUsolBUQhfGL1a57FJB/ZaCrJ0EsfX5EOIk06Bs
ecpWNAf92GODXCuI5UHL23O6VthMMcDd2z6r93oi2d4GGXUfiI9YBd1XtEFw
ca7C0k3Zla8t8tdmOHRUJP16WvjO2Nt3g6xCw02evsTBjCqLaN7yZnkHcVpU
sk7/klY2jV7i9f/dOTOaK8leoZyOkcDmsqdw45ipVLfZnmXzgPfrXcUx7IXr
AykJaIwFOaE2iw6+zWUXPbibqTaagA5Xk0Weja2hYT02nC8tzL9wMAO98ExZ
k60c9ZTDW+LoCEJpQTK3DdwZPWr6A6J7ujIHG5pHKRa8s3FiYY5Xec1lx9Y0
Ym7AawdyrEC0kntatuUOL71wriw6u/fKmlY+UeF/DoVdw2HiDRi1jqaXqDu9
OXsCpaZwvfVqDupRRbaZ75rKE7FE79sCcxWKZR9fuf16tgQKv+/TQ79QwsWk
1DOzpENFEkT5SFL3sR01OpxXKExkPzI5fRvxZsCSR+4utrz95lIqW272DzF+
+Zp2gU6K4pOo5n71UlBEUZhn9rFaxwnr7SPjjIr+omWMeZVnSSTa+6nAdets
ZP5XwHxEcQwxSeMHTatsv5SWsH3cmMpILmeNLWKpI6wNWdUgX7eUS7ycyaEX
vc/MA9mNbAZcpmQ4lN4K4+cYL0LliF2J7dx6HVH7f5kb4fARFFBzjk9gEtF+
BsD5ff+FoGybs5DesVP3BIUqP9prKoTVQhd8dXHAhwIOWw/fXPZQ9uolZrqy
kv40DhCuTzRZ4IZO8tIlxH7/3juBeI8kVLt/MsDQrzDc8wcDNN1ifvGUHFUv
/QOxE48NVl5ZYCTxQFgQudM0Y+Lh0ZusWHb508EsmeVj5Mhd+G8qEkECgUVd
qsFWiL8Z60eq4D/+t+R1PliKqBGt4O/QywJzbpSO3Mu7aFCyXqKy/e8n8qy7
bqq12M7fNXDtqDwJYj/Y9pBtc5LdAzi3EzG3C2pALj3AdY/BFWzrG+TInhN8
fwtQm4G/VK9bXoMfIfm3MyhZCuJstb/CalZQoJmpXTaNslOKjMc86FJYUrv6
2DtzxGCQGcO1T8pCAaTQdWO9q4pKSy/LotYRMx5D/og97r6cpeFDv7BoJJoU
LlrK1PVBFGejq7qhlbK6+lmR8i9t3EU9SvnwjuLO5IyYtb/VhMWou40v64Ds
W+eNTCFh5/lu+9ThrI6R6rBwqSnYCc6s4rRJ1xsZdcLOuaJTfc02Qt0jKmDl
6wtGoXHrI+HBe9u9S4nB3RPrhzqiigljIce/mePd8xh0N1sgmA/D6YIMDmiB
80v5m76towyzHeaOi4zEFkHjeLAM8CTXy4BNhcM4FwbYTscL7DuOLhUpWoNQ
pt/wzTYUm1nozzIDHHn6ePV5AbDyrWRsVZ1a65QkWPvNI0ed2GG3F1UodE7k
lq569xcajQiw5bB1td03YLATxg+chkqJK1AUEbZt5sO6nugPBKy5xvC0uGSe
lspzAGw6RmQfJHS2f8sDHjQ3VZrUTHZorwxTG1l0r6X3MtlzwyiqFJi7Agtm
CRrRxjRmRrPavT44GNwpGw5oPSDP/ohSqCosEGceLSg+rr0e3T3bp14vkK87
WXmTpU/WvcH/ViE2KkvwlApFsdl/jfTYIZXiU23zTTQpl7R26X0JAVh5DaOl
j+tsjvYIgLsavtOsklTwvkUSjeHMEeam4XSwcvpEXKm8l6wCiiA8XIwkHRnu
cPOYbmgnuMfV7328cXvU30/birilMjhtZsYc7dkp1GdxTbhu35JW5YmmwlsZ
LeL1S9ehya6lYyrg9p1+Nn/YtAMWr0IyaNMwZM784wb00R8wogXgyehKysuC
njv6CopnrCtyss97nptGoQsM3n8C87In3ZFe8OPEhjHSLC0cOMlpVJFLkZw/
wc/+my6+lmm1Y3wUM9olgEE8YxVD53VSYaw9DwZOjiHvcyAt/p7AGd9+Qjg6
D0VMw5Orl2LMyIFyiEjo5eQPzp4DWB8JX3Wrslr2pjeJoKXm6iosNOjcpk76
1yAdqz4aZpBBRMdv9GcxvOczHD8Ivhnq9QaRCS+4qSgS9JmtAylOVnSmeMyd
oEvkWX2N+gD+7jJ4ssI6zyjLw6Uc/UNLwsAwHIcU455JXftFe0nZUtLbs6Km
CzmkO6i0MHt0hK6dQH9Pl9mC0q43AScI2wbHtGVx+KkGg17WYawuyCQe+W6/
sVyuhbkAwpq7yp01SZ6/Jo60k3yOw4mw6cumUX8V1RKD8ARfwkCaaAZ5Y0DT
whhSwNYARSKuHMaSJ9yFGEbufFNWETc9/ekL6X/E8j6pmeN3kOzMQTfjOSQT
BdEj5JPhvJW9M+WUDo0H6rGFIV8msumzmHNwSwip6KEk18kRoWMhpbSufduX
y8jY4yq3YP00k0RMmE0eJ0oqVJlfr+OS+byce6iO1mzzaWZFZgVQ3J/Bke+s
8jQZaXALNEP2FAIC5AFDjw3FAp6NmpCV6xyGneJNth0rN0J/GYOM7l+sJun0
fwZuG7UJGIqRCknEZu64pNYFNiGbn5p4L+z/QRRZrKyZq9ZPl3E2hKHANA/a
bV/9X8bRjeDmgon5DdhJ+h0nSSRp0+PVFydXi1pKceGH+7vHoKqeKGI8B6pJ
rtZtn5iEf1wq0VzOrJSY9cOKHFQLD2YRC2ZttU+d7LjXI3AZuOHb/bJmystB
cU13xqmOpM/P6RWoUi2aZXztGNivja6v9S6vIbIdCi3hKHhnyPKAncko25q5
stwvkOLR/c1MbMinVfMD5Z908GUItDa7UmCx+Ryx9rhyGwnJveZpS1UMbXOP
1QpczVDKVRG0PkrvHJ4qr2yTWFRR4eMa1YFKUP6cdsbgNjOtMn2ymSNp1y11
+iLK2F6Pu8eDhJS4Oqq84vC9Ai4OYV4frlYY2Du5B3UC70Pfd/Exuc/2uD+9
YLxNBTgIaaEyrN9nBIfqmSrLSs0/aipZ5kXTbaFxIfLxKVKPfHmJTe3RpB2U
cRiW4BtSFz7rsKAgYp4U+KZQPUi4MO15YCWknU5BQ56eSD66Cnc+rjzAClQ8
282VmKOZFYhNs9opyf2BFjq8SuwJRgTtiugi9ucbb55MrNYAizJdz3pXRlOe
3xsAmV6tbjFX3mtKKF56S/pnd7bVfaJ6qRe9nTgdGWm0OwSbeEf/dVDrBl5+
HmGWeoIm2m2/7z8oeQOfxgN9QiUIyGkuwycqtvr5SMCOG2qjKCe5O8w03kJ2
7ks8iTtk6QmQewqRcpVtq3Y2QFpkce2LvLUQnLaFIH2NBQMtIZrWihB/sRLO
yx4cxUHQ2nIe5RhJnOXkZP+GonskSG9CwawyMalWXqHANprkQx/zx1ILrEJM
ynC1HwGmx00gwBK2OWHRzj/vNWpo9K/gjtWpmszJPm5voMSgvghmzmni5bdl
KISgvVm8+DwL94IA8cnR0ja5oaOJJHoUkkdE+e3NVKl15UVdFge/ie9r2KQv
F04cgZBc+kl6aNiX3aarL2pkUN6OX8jtlX2ZfeQdXcTPLIYIoQjJ/VQarV2q
TfrpLLcaHHq+MCaXKuuKxeQC/23VpVg57oAh5TAmjGVZqo4bK+CsHF/YM9c6
QrjcNeot75mGj+UCy00fMoNTuD99UiEire4kQmUt/CagLqArgqomFhDLgyUC
wW5Yz+Ft6teJJKlD1TlStPz0srxiDe25wmhoES4LwcDKXeQNvM7WkHmZnJVZ
lx2E3Z17bH63TtO8XDly7pCJ1B6oZYVdQLF4YP+qcgmZDCuuhvIXaF4U/o9F
dJhI0QTVvM4SSQZw5mG0GS6P5Kj9LzL/o8XgTVM6mPGQ8mPtf9jKuj5LXuEH
7f9oRO5pZecUQq4lAErtN1E0BWqCgfR4kdmigTQJRKlwephRbG+hgW0prvYZ
4ntdo7i3rTYRGz36TuhG4qTS1GboVae6EyMRjrSQjmphIDfb8Ui60Zcy+NG5
W8LfKUeiz65TR7Cvio+qd4o8nR/1Di3FT3PHg3fhJAwlBkE7rF3trCVOhVPM
97WyX38DdI1sK+TrIu9Lf/P3qln3d/kYScQjvtwYPmb8kMZRBcleSy1pcR0s
zE0x7zmn6B9vjF5w8AJHHLUvewRwH/gJcbMGmRy1tq8ptqvcLGldVmGJKDnw
IsrqPTI+v2wQCs1YfoTPBdftuQNToz6gFfjuFwnHz7+ffpuoSA80BenJD+I7
SjqJrLgpfDFcCd77MdiUDkRnjYgS3BdsUqBVOxfByehVn4ES8388dpK9HZZk
K4D986YZYkl3QVz96+/79H85JDXZcm9a+m+Z2yxkX7WO4nFGoj3a93FxDF0Z
u7FhHpbuKRSPvT60h+TH1l+/fLj4BhVht3QamaKvZ5pvczuJoc23oCFLHLed
3Twi9KFOxKBhPIGzeSwR/A2LvXbVZcET6COxUqhSPeJ+fQ4G1tpF1HOkVjsK
N2O7/jRG7HOXgo+owrOs+j/OOqE5VFgm3Z7/AKo0ZYzshiKOkYPYJN6MxTea
0lh3NNMN0uh9cdxMbWvw/S3SUsfzvDkakiUHjWoYe3LoTtbdLMYOCepSb96E
dnEYg58Tolc5TC+RV952U9MSIryMlDcpa5chUUANQBXfjOCyfaB06r/dEfyh
/BR2Gn/MTE8mDD/JAFZ95V6bIL7H7lgbm8AEC80MTyPMAevJSysbkMHG/wJV
SHuz/CoOLn2vU7l4fY2OpnFA09U4pyY2XZG56qzzftBRrJPY9nMVejsgawWd
scforXqm2sAX0CfMBisXaMmgxyEYJ/c+qlEmwgUjspl2cmRSuuaggCH0xGBH
19KKTm/aeZ+6DkcNY08k2Y+jOL8XLfttkEF/JYigCRqlUZWdbtJNm6L/Xsly
RMStpySS62EpNGcS/yopKeFEbrKmwukQC1v2yQL/5SfF9m42wXO49CsQCbQg
4jIDe9tPttw4k9jpsxw5iZrLtP9j8BBel3EECsgbdrOAMe0l2vlEvE8CnBkc
OBCI7YRy6Ik29+7oaYBwsFM095B0wYLKlF36nzlpFq9QSJ/fR+mJi+sC+DeZ
6BPJBrbbxM3kEX3+L/Hi2oFsig9M0zA1qCx1VMt0Bm9l8FJPd8B41Wyg4ZnE
F/hFoknJvJ0qG77QZb79tSQsGn4FUyfJ7Hir9XAJ93slTx8KPawmG5uRMc+D
tZo/EK7TNqbN1GfpmAVnM3LAW8NYCIHBfT87Ih1F8hBhq+ZXQO9sqsG1K6tB
1o4S07Tlk5n5Q9SFCIw6xJMDi5waeGS0COogYRwxANrljGH0H1l87/qmpCge
8r5PelbOnvkXv9ntJLwV0QepEjlCjUbVR5OgUZhkW2NMYMchvI/T2evIgf/9
s/NK5yjXzHq6b0H0u/Tkd9b99c9h+6M31PBiGKkrXWhqVdIhBcQmIRWf1BrO
y3XyvhcwK7GIpv+/icRDUNZKkvYTXs1WwV2LvOVh3mnLsaQUTvrdPOmOo30M
J+Nx3ZlLDNKfb2XRODdHKxG13zfasOliz8RLr7JJG8uOgZ1Rf5QnfJkjHU/U
/vUKO+WAtkvWAchNu8mX7Km23hkXxyq1DgvpjBiyiQ5CjiMUMhm23KhRo9eM
APaJ0mcT99iYKO7qjMmUfaHfsBLo1XUt3Rti2Snby1EaOERuo2kTKr2N21Ul
v0h+P8JY2B3UMdo+QFymcnoxDPXCrmIts7/DHCF02JNwOxNvBg7d3rVPmRS8
9W9A0vmvqz5wr3VPSFqGvJ/enqtNirok/PEC+KCB/xwMcst7E5smhlRGXGAP
/0JXjIIaYZ0FOrSuIcY7S1KPHIsqnXuxGGUULHYx3DCk8e7L9tqS8vo3p2AV
Xp2i71WRbjHyLb7b30pciC+OBZ4Ud8QV1ltZ8/uhsZh5/6zoET3pwm/v+7lH
szoLa9f1y+P3IWRHsr6FJl+ZJBCU6X60ollludxQOR25YKNYNNJ4cYTFsECq
Qvt/K1OOQc3wlGaT64Pso6TpWMXfbOJNeAsWTsCqVl0ozuKWEwc5jPC3QvK2
Vq4J/DpZl6X1GLN4lXbRFj0A2joHQ5yNr60UfiUFn/IJvTZbgIkfBYjWXBCu
wJ16Li7hx1XlV1jUR99qtwCjkNV4LNV/m0SpK+5y38ul6dg51iE4fKpv8p6H
gvHkeaFIikBd9Rs8W6xE8aGImF7Vkq08FaLYrSE+HQ5VpZsytdH9/Irvcvad
JtqOT+GPtQeTpSeK4MhgU8lm+T42qNK/SaTvVtAU0TdrGlPgPpEjKe9byHA0
N//lbrPkHRBoi1NcOfHW8vSg+GQU1rcKUhL05S0tDPsLARJyxk9nagR9i33e
vKtVQHes0fnjvlQ1u3CgFU5CsWyCYfg0DapVw0m8qvtBNUadFVOkwTvUjcIa
zjsxttl6Q+isQPl7Drv1q7A/Tz1SjkVV0XK/VIYG/1Bksu3VfD9cKiTjRZ2a
WBrYLnmSxUeopZxs9yGVqct2OLq7EW5dBdkurxawXZ6xFSU30H4I1fN4zR17
fXeiUJdeA64Hgn9RBuVOdBlNUfBJAH0+MrhIAKepaG3sqkKKkcUhsoVjqUtv
sBtIPYQK65HFXddhUhZxhVM56L20rwWBmpnrksfJoYCtrv7GuoEIs475SP5q
5kzw6Pa2WsYkvqz/9OP52lX0VkSeKVM13FrEUjw5LZBeUMRzuUAP5EgsHrEI
PHfEMgF1bJiLD5Kxnm7pyy+gzHtRtn8o+whWws6pLUP0KYfsbY71Lm1nsqca
kZtVODo+MXfyTCXnrfGfCn6X9JLGNsQVwCYZb7yJ7u2uDnnJTPSo/MhgercN
pXrvzrFDd8vykFeVfU4C0IOkZfXQO2PDKJ/XBgsXFSeQ7WR6jqyaf8h3X4qz
SiRdte0ql9C1N14c62O1heHq2aHsf2VP47GrGCwquQqazO/1R0g5ViY1wc8i
d66Rg8S/TLuaQH/GkKNC7SukDsUeocojltio+MG8LxqbE4yeGx5eu5/taJlx
937Z0FSDkHdmwKFHLzTCLORhdlC5aTW3M7BzkMwDTLbFpBipHxJZEiGqm+zL
i7fR7nX7wzD/x/7l3Z7vm0822WPLxExJwkojplLGIKowD1cq4XMvGdNQek7f
/t9Ed0YtNKni8CcYe0xr5q7+dlrY0UOd8kJgVhnAtWrbq63hhNiX86dX/6lc
E3yks4ttM8Mh6D37/8p4Rby9aufUkbkFXLiNpVw7lL0KlWCSU4kh5HUOJ3kb
YwrZ80ajdNoOG5dI68kPtWyKTt4e3Ho8wmeasSXcLfVynqtbaYKCJpTBqO3W
DsDCCsi0p3jzkTDdDHXlYTa/wAsAp0oZK00zGKiqmXwtZVF6+nCg9u5vzT+r
NKlHHm6Uq/9EWWrhkXuZnD8DWnhJtZ4O4SSxLQakidfeV67yQmDeKZNGzyZz
ATALYLD2QU3EcJtS4kdoVy7Vg8JbUfIz06CqLqdaEg/I7uuvJbISvWVcfEMe
mkl+BFsYvVYg5NmYTxustvgToVRzCOawhnysvBYhpvK6fsWJaQOb3sL1QNTT
c/jIF18A1/2oUq+9FdRKoQGyxhbSFuY13CGOXRs/O4zR+CLiD8HKz3VXVZ4p
t2KMzU+QmZXQ0YRGa6X1SLEyg9+9wdsg9bcsNo1tZQHyWD3TEEOoAc65dyPD
a46CZp3lK2uUYaGrLBu6vZ/OC15usnFAyllwKHWZkgOmefuthT6i6f4CGKJ9
CpNCZNm3quLtqKrvOpwoh/2XDL9fbZxgw/0lSpwYuJMDo/Y3rpnYAefCTLO0
nrvHupt9M+3sN1syCOhZ+f7xbhYQBI8Vp0fUegEPRN7oIWvWXGrWrcUd3lDU
tIhv+AV9pSQ6Mt4fb+hzfsZ+k8cuUw0vXVpLI9WJXKOs7T6TS9e8K0Hbit8O
tLUFaYuLmVneGMSMSFUjPBAJX4IaGnD2Zg791aJvGNHnos59KXlcItchGAGT
K0awD4xXYNg8Vocis35oYtv9EID++pHiCSEHCptMSL/feKDxVKfr4R9DF+Sr
+VdpxeTWof+Ry7t0ZMWYt7FchC2HBzKcX1DcIZ4s8RCeGo1lBbHEAY6Ez4pX
32IVLIEzKW2aU4IJK+A3Gm05CR+biPloP7H6aOat3TrZ4BwJ9wfptCSjeWgD
CahQsPCV39soKAr+JDPUlqAFD3EqppeDZjm9+GPhA2p4LfgpY0aqdVaBFZkp
NsZRpfpUsPiWKrBO8G6CnJ0t8SjMLTtRZ8ISulJ2eYJIqO7wZl7bPP5IXmDX
ytE00eT4ZVjwmqfo9wWsX44WJ3CexJZjjHYB9nhCJjoDmCMajnWKUzYAjVwK
ysWeLMp1KfBO2XM7MnsDnNQ0Z6yX6SpHRCKTEdOmSv6zH4Oi2gRKF5rNrdqt
TT2SAJ8sPH2o5jPVsZ6tjfcmxkhqSpZValEngGZM6aXbXmZNdCoLoWsjBaJ/
JE1gF9AsnxCJUNo8UstkRhF08qCGkdy3DkCq9eGb4VX0dAWQHR85Dz7O6I5h
8QBaVdmpbh7Jry2aFq4t2SdXUYBmgUpRzwGNLVR7kbEIdmxi1GeyoJ4ZjjXy
BTgrq0CsfWR540md0A0N0KU6U5QYGJVPHvlpauIZ923yQ9qYWjU1d0NdvBmu
snKrtYuNB4jo+QXa2j0n5i0KJyC8IdIf9x1wz/vMSr7LtVHb797R+gHT5ZoJ
NJ5bDW1Za+IrGqFLONDDpwirpAIHduJjBh0naY+WQE1WQycZkn7XFgvQYkr9
PssmxgT8RJ3YHP+XA5eCr2ChzETKJx0P3MFiJanKSdNzKAVCtfteunXmTT3m
XnHRdNNEl2xa1Q2hWV+iQpBj0wBApDF3NSgOLOlC2gzGrAQlB1Jl6/lJzgfx
eY7OUhvVJRK9JhHOuU5DxUmF6nb5TMQxZbqHTjDV2jC3l7P4bPM/7ZcL7hPl
2J0ZGeUlZlj2Def0OlyJcPcxUyGg51htBbEfjQY+lbv+rkZBxDVmqrMkhHEG
o0VTH4u3IJC0lphDcrLf2sjsTE0aNsbObK2GtoA7i/C4h/+Cb/SofNMi+HXx
QEjzm0UoHqKYAhTa0L8emt0qd2qpayG2WrqAti88/yZmGEjGFDfG3ljvY5dK
kgeuhpTr4YEuYl7S/hAqQYBGr5B7aNW6gygIyzNKWac+uA1sAc/AG1IZK5MO
gTMAAOsJCpO9koykCkOL3q+hBcx7mi8xKT3encRDDh0Z07ixAWuuiJ25Qw1z
tDQgT4uwer28Rq2VInWb6oW0WpD1or2DmVvt8dm+qGQ6MJF4gAFmIQ1g8xPi
nLx2yNqPO8cWirt+/CDoWaLmxWBrog2SpzkGwDuUfPJ9eI29M1AlkS8SpvWh
So+LdA6NCuDntpXZocQ/bHwaiFFi2SiFaUUGRZTIxMKHO9DnP2Vjbpd8L5yf
x74DCsE/LYxUDEddeTMigLqkXJuX5/0W448pwqKjq7/gmw2VgTu/4ey4Uiwq
3Tn7sJHNxQPFvfcALQY8YufAE/M9lVLUz7HxOivwXbIMXH1Hdf/4Bc+inQWF
VvMX9E/wrZJrXi/mCDXdnpqM/6AeZVHohijlKKK1puZBRHL1NxH2L12g+/zt
5VVGRFj7FOKOCfSUguRJ1KI+tuHWUo5PVgxCVgOAv9UDVAUnuV35s0h5CFWa
laDKLgoP4pYORG4FdQpNFEQWoh3ogTYaJqUpt9AP97qwD2qCJJAuqxTiUnw8
oE8sn1aSQAcaj+H8hS5ZHlXZJWYNgxP0K3+vxhlsSDjOlEfLEY6ukcdI+hFa
h8p2Vh3a+J8HxRoYegMqMQX9FW+YMCyIkwlzjFtvOLn1GUn7mGCHAL4KQqyV
38C1D8L+avOYlyJVKTrWfF3cLAGZ5bosjmsjdpyYJda3a0l6l0AYfpeFLEdp
q663H6TAjfaR5UwoNhK4DRHphhEMouRcXdgunoI2Yg5RZ4mHnDhdZsi7J104
5Wsfz7feiEzzIDhg2p9cgeyRR5Hwi/xPuuYMWllkIzggI/CdU+GuGn51dx+J
R3sE39D9SLQlT1duJBgNKw0Tce7mjTwM0Jq3Os1RP0M6wBWzNZ/lvbWTPgcE
4wmtg3xAc51OuWUH4Vg4HIV3qZM3anRwH/Z63pRhXPd/mr/tSypUkp/XDmow
HQVnZRx/Wur7+8ROM/txeZ4Ri/J5pckJ6bCwhlfJZjtWgNFhqlCBXte9FYCB
fC43Plh6uSkI7J3/8VmqAF+Df3ekfG1goxmvfZ36DGAcbj+1U9v3I6gUW/pg
rFcm/Zs4f7QJCvybX+KUhw3yaf0AgpuS/jCAoV5+D/q0E1vUvLSac+ILy8uz
m7Qa1cneFDLeWcUu/6xqNlr0kIgMyBkoAaLm+RnR38Nk2Bd6POOkLeVXOJB7
pGlp/XNGGmFh+n+oM+hdFqrl1am+izKvk70mcgWHIEE3Vz5rbqDHKpsgeCFa
UVzhVKE7L2/BMgoR4R5oOfQt7OGHYOtX6vUFRZTnPjT+2X/eYRybugXTzupA
QdiCKchiSmQ14fGVSwAbMzANz1odkiBhJr92x0W2BGkA3Mb6Npfe5pSVLgZc
oNf4kvOlQsjTf7o1MtXOUZiB40QKwx9bcFRlWD+XdOjfCbVlxwOdXivws3kN
I2wjqHnoHj91jcRIAqtMmHBi3+d8S/sYWY1tnOCLPh+12m4+2lyps2/I2yVU
Gp07aaRu27M6xJCg0WDvG70/EICIJ1NoorA7wH7xhCfe0r4sfK37W7DeQPvr
P9en01veoDf1KZ/Hq7obEJnf99lJT7xKPlW5UJJzXUYjReiTVHsCYQRYXJ/6
PoOgSAjUnrKMm++dNZw3kXZ51lWhUax0MH7/dqvWK3THKfLYjAOfZlNIpFvC
88smPmq+l8Uokzapkme5ofRsG4sSiyB2IyhhcIQd83qJAA/xWFchGEOnE1lc
CxG+AT/0PO5bjNh2GIbB72zMzeE44CjwDmnlLCjD0NJ9o/0qj5/IQCKhXAKS
b0IiTtznD0cIqRpeaZKYEL2A/wuq0LKHwB2DvsnjTZp7ucAOUMy7K5wbHC8K
d6X80kadUSsxVUmA7/K7CWyDxw4di3G1FthrC5x/gP92ADRXcmGihkV98hq6
uMNTlTIvJXOy7nXW67S3gTGj5FRcl1w0VWW6sAzOv6KnFD0SL3Goj8Y6y+dD
BWbKbffCvj8zuQNt7d18e0gFdtQXMtcUKR4sYeASEtp81N20KFv/m2Dr0Q0F
Li1aqEYdjhWDVpBlVujYWAGf1RiYX+HnQx8In0ZLG90d88urz0PSHPW/T4D5
PdoCON6VVqtuCrGbmVRbXtGYP0ulGqMAoJpjjzZTz6B70EI6wK0H2AMZWmes
uca7m6zhEBog1c4sapdcSui/6TFPNT6N3bTYFktiPaUnfSzdP8Q6XltJCcWc
msF/dN2eCunC/yNsHbI4/AJ3J+LZASPF3TPZbFRh2crYaMteQrUs5NjvkuPl
+H7lT7ZJfFdFHGCxsHMCJC6kifamTe2cRBCg9JvSz+2q3mN7+N6o6EGGCihf
9o3zci/ins5wI5ir0S9UkO18t071zWHO3PIiFcLbz/GWT6Pc8tFSLRDuTRPN
ojyBQ04Nak64uC8J0u/G6r4c8bI2Qe6WiXTdJK+I3OLZPN9AUqYsVpCcCo9i
346XVPaGfq6SukRwisQysJemt1xS/d/EH1DuZWMOy2HxAt6mucNAAft+ZdfY
8sEHLhda7APQnExEc9CGTn6z4ZYBFvaWhD3wbS6ZNLK7QLLffKBebPdSEDjM
hacOQBuuqDNgZFEKQuxn2J+SWAHYhSD2Obc2vtIGbpw3ysSOLlXEfgO8XLiS
D1mhAqufXUHtRjI8ouUQr9mJzPOYbhS0dOnrpz61mvW9u81UhEBxuOTzWjTh
iAdddlPl2ItJDRSYRqTn+QCIEExcyK1S1KGE3FsyBjBh8vRS6pdP9bxaKrIm
LktEUxo07GUXRfGxCO1QWOEek9GN5y47isTxdne2RQZldb414nbYXqxnKcDn
3QGC36ksTYDVCmkUB55vYcGlMC73uC4dIe/PD7xHciNoNBeKJTlSmEz/grvw
WFcY1dTSQQeH0npVgk+ppWKntc1JGWUwkkQpZgnmsmA25RspnS9uSsEVlgTT
j0aHNrgezgDk9hw2TCTIzZpbfrA5zCjTDKQvgR007B8or7wj63KlqbZ5LLJ8
H9nkaKbgzES5k1IM1/YFUCd2AegqK/W/6MDYhSGu7mHk8UUi43rWNTo/RfnA
ZmQYbzQJh+QlbR0QvUGHne9HMCBD/C53MG2+I88wU7iFfG36m4zDP/NIQPwl
2ArtUEq6qCujBDrXq79CJB2FP4zJmPm81/nG67zUlj9S7YDM0YATn6/Iwigy
2kzRjbW4uT4fDkhUGqao6Y4RUmiA6veMr/85gWE7yySv3z0jvBVwGlhxeShO
fA67j2t8LOcd+yOpDMq7lMTEIMvAVbgwm9HT+Sf1BmwTx/HREgzFl14nRAf6
QrO3kdPP18h2EDJejIKEQzTPYgOnt+/+iQIRjmpsdbQ6X1nqggDt+M+b5Ysf
v162i/GgQlkVJVznjOti0jyGKWaQUm75i2SR9TEwcAKpJV1MZEi/9pJwG6/d
cYr4yHR1LSn/6g9OimjVNYj7KQfxxhKXKLHVMpeS7dmyheHx8Ml29S1DTcbd
HCPHi6Q3H3SrZCmwq/y9leWpxJ7PzRYFaRcjcRr9NQ9eDn0m2ScZO1bjXkY8
oWXb5JXAeZpgSP9Ykr/yMPMvad9Q2ymUvASCIPE5bdQNqdIafrrFSXIuHTvJ
udZAbQBuOYm2C6q8fCJp4EFT04CHRmMjJez7g1y8HNQz8kHQVOA1tFWQZ426
ggsyurzcfdS4lVe72ZDEw/SAqEvH8ohBZf7Q8hJOk+XIiNjUu1+Tmnmxlfcm
/O9Di5ZNZPC7tDyVyNXYci6eTClMaoLkTTeCS5Cj5SNVwVE7ZGqxf33HSQtN
buc4YxFX1HTOsNinSvJEcbpinAwKx+FqOLIrzxVLWOde5T4fZMHzkN7eiZ0z
/Pq4pRiClWnPGWugoKXysb/qmUUibVHAhLzWNNneI8HGUTdW8/S48e/UPM1B
Efb0MbTjC/K3s5H/JVQZ3pfKMG/9fs+Xe8WG9dcrC+RU8vjH2vcb3M5Xzcxq
JmEFtlTzHlTFPt7JEF9njOHSGC1gcrexEB5n6ERKZN6OjQERtp5xbYLsALRZ
tru99ZN8ho8vvjNG2DsGPoX+kzepnOfnAY/ggcE6liliK918rRMOrWWrpzM7
wS01vgE50G3H7tIQCnfMgIOOikjaWMtU/CE1NlLhlaAa74Qq9TXtFHK0JdBu
asLHdcpTMi7XUNLdaQl4GBsikJin8uKkkcw5SYzHGC0kKClXyv0HKlG31rVS
QRNaa2a0cPsZg77VcJJyCwtulAzT/LKJ+xuuTBmPCjnnfyICUnxAdcLEWWzt
W8uXMyHon3IiP6GCODMe2SSsF4wO3pfTkvNjrk5boe3bJ5nDFIoEp8NKziz9
HvB9WQqW8cWYkBVF3ZbW17/UEz9SqFAvOoMOftQTxg0RA2K1uPPsOpw9w78H
vQxt42IWHHI8PwwkgsVmhBLM3uBRSBuOZy2OJnkgzOFwh+TGUk758anK9Blb
ccnhfJBGpNMDBFIwtoy3W8m8YFVgma62l2uQWuQXaFLKgJbUO10xmo/of6IM
PS4mSbJgMN3rDdkBX2yovYzIM50M/ulAmWCZVohxaUf7MOtQQVcjAurhFci3
1UudtOi9T3uirtpZe+VbrbyC9mwXmsDfWUTvkA3i6LQ4PU1N2LusZm+1FN8f
/YSiAsdmsheKKMsQFQQsyULlbGfzaULOBwL7GoE1zFYMUMncnR1DkiLTOr+n
EqlRM4TZqV5BmOnApMKHFJk7E3GYj/CBBPCvn8oner1cdYjYKR37Ai1byU4r
MJg12RT6pucpWGoUr6Cxxv3jIznOLhHwXGjRvOWGBKe+IphWRrzfgz0bzXik
GNKEDsNHxgBGmyhHTtF1kohNtGyiNWIeW5Jsom1q/SKkxtVo43DMnKVaokI5
GVgZSVPlxwsJ1Hl+SzuQEo+xTa66Be7kGVv/ZI7qiQGGY0mR1sl0xjZZh1Kx
QNKqrcGSknx4QiKEos2j8k2HaxKSTqwdZszUfCeJlhXBezwjr8js9X7zrFB6
NC6BJ3iPNgeHLDq0WXjYIefX/bjOLhWizKtp1eaRpj6LSKJeEOL84wzA6nbt
+PSGhEOWZSxmzzXU0bbpcrWwNRBZ3ZM0uWAI7y8q52cL/jS35lDFWeJVIDJn
ZDCMMFRxLydyPqBmrWLzAmOOoEBtPU+FNQitpvGRlgE2Rh+rSjOtYjqvNTId
c9P2Eu0n6WSv0KXdwE+QZ+jZe6Rwj5wI/6PNjimIWcFzGwvJ7WwzoZT6QLK4
kxKic3wlzW+tby1yAu55JOXphkIn4pOKaonA5fpWQo+7dyOfX3tBR5VgSEDr
iZWEjXwG02ksq0bRoEklp77dF8M2PBpNAUgYiJcgY8e2B/RPYHNOXTM9yNvI
3CSBl33V/7KOEtfJk0GGxphE5AxuXBdoLzf3uGQC4zYZMvqkqp0xPNCM9x7e
/c4O8ORAOao0hIQSE7GcEjJzrKpkBSpBE9mtfuo+mTIub9NCoZK2ZAWDvKH+
/FYeu/wGCDFhQpJDqeiAF1WmItXPljH8qOd2YLFPSq7D2XXBdXZKM4/rquop
egk0nE+xWAFu598cC8ImSaGfPJngFg0ZQLKqvVRbyjKpbEhUdzeQdslv+N0m
O0eHpQ36bCf343/hRlSe3zwpHrl7La03rBnscqEW74Aopx+9ucASj2Hf4dki
fkEwLgFQ3F8Ydu4ZiO2/gKYECSjYjA14tKDJHYoBB9l13BJxbudOOusnRufm
mW3ljreGk3QTowBHFxcvsZZv8dcVFQGg4HdgSIlG2rOQAkvc5TtK95KQOvnj
oYR026nWSFciRsVpRwjkpWkUR0bxqghyn0/uzfkv8okw1jV1klzU/o+WgI6V
RuN/2D/ivXo9gclZ4sop5b9yia1rWwG8CERipvCEoem7pyC2zPxjU8HdALV+
I3VbHFWrjWSaC/jOggFt4ivPKn7scURTt4o3xpxRn9aVRp0G2kQOe/jDuooB
RBCfSWLyne+Vy3ogse5i7MR3pP2NZLEIOgZnGfh0/TN4Ta8tiM4pHQotVcKi
npxWz1Bexkc7kWNfgXq3aHXsgAf97WkLeLRUpbPqqYGjMrYoKZ8G2pV099MS
s/0pFmaUjjnmiqL7pW1mHw67sGtF8nB1DZkt0DxUKIJhcFHuYl8BoBkiI+rf
omg4r40HynR72lLJXPVJx8JmQDWRhMf7WIsXcTNKyYWgthfT9wYETA0ccLcL
qOZGJrtQQqJ7b5RY2YuykSV/wKSN1fhdYDkqMhvVF6WTNHOQd1sVCAAsDwp1
7u/ZRgWk4nZTw/FTiyZVP/OcJmSc3jE9BHr82BexQ16GG+BWr0nhxogCkbgn
AFZWBu47R7hHYMcoZK8/hLhiDb/eq8by3Wbn2C0sOEk5NU3OFwgHawPk/lHf
2W+6CV085VfnKoIpkBUdc6D+pzJyq7ZiBgOMUWQ57kGaTH3z8CzF720JbpMY
7vdDPbPe7kv6ALcL48rlO53N7qEp90w8R+AjAfSOOgWnxU9HZIbMxpE+Vsls
NY/43tZhVzrAhEYbEi7Y3y9DQT4gx3eT8fixV5DufUmfgXT8SL18rknp0r9n
1kMOwoRdXoQO4Nj2s6b1RynvEWoZPJ4XwnDN7cJzYJNhz8TVAihW0DD8Vcfp
NaXgplHK7YaWrYUNu8D2G5lwlnX68oPVYpztNDIUXyaSXc0CSh2CbwXq4022
/g7FVTpHrqZfy5/wkBElIVt3qI3Vbv6k/FjWdcfcj+PYmO/q53wRJ1v7p2dC
E8dmKyoLano84hrJoqtlKE7UemxsOh6C3a9U2vjkJYq+28j+NK2YOOVyVoIT
UHUb150MI9C+5z8iwGH8Kl04NlTkoYOx4jiCEP2Fjc8+rzpUnUyCdluwHdPR
dk+HIYMdAwQlnOP4VlGR6deanlf2U39OSyegRo9lChtVkjbNr0tNLMZ7JQCd
9lNvGmlDEVWQQFfQkv5bHk3GQexdOkh0QUqd9WWSge5xwzmL0Ns9WUu+tmu5
i0VlSDb8/ngCIe10cquE8LgfA1LJZRpd/KQUX45LHy5oVMSTerosRJu/RVQn
IF27WxeW/64WpeNEcFryHY5zx2OHCewnWULonQ3aH82fXVqjpCwZfX/34vnj
TRsX+KsfUypnE1YQhzpwHB9LyNLyy4/Efna8fEIGjOSvt8uN9kaqVciRVFwD
rcIvTkSFK986f3VAgzL81f1ifPysBWeCug7lPwn7aTJ9nVVKdughB+yOCTYe
JItMXLCEyJ5VGeLO3xMWAeMHSXXHTLcfHAxI7ULoMAN4wbiit5Vp1ewts8GS
FZVHTXqLEJ39jkNVHLhvCWOC2CLPr9+tDa86lUhuNLiq7rqvK9QkvI6IaaI3
DE69Sm/IZ+M3rgjnog2FMufLV28216ZoEqJdoPSjVTOh0RN+oCfh+VBbExyA
1UvJJpvwEx4f0WfgAjjkXTQWQUvsgJu9XBhYejx9EHkixQ5uV3UFYkjaWINx
vf8n7UFXITCPYjGQDDeqHhk+W+YK7IVQow2HzxcMs9ZDrSmAmvdlyF2UPga5
cNSS5zR97kl7UR3QYRmcR1bsa2Le+FgQgVPz3yUXIJ56Xbt2qzi8AhGvKs4m
xHylyC9Jc47LkFzAB+YCu+HDvwUgjBylMVXItzPazFmZU+kwOmuzBZRGKXUW
ZE4p88X+w0lgFOcqReeXhD5tYb0n1NLtnfyLR027MDPcplJ0kttbz30+9oqI
xvXcmFKHNjqH1SA0goalGwJh7PoCPrS7mZL6mdKNzzSDRh3BTwdmIWz0gTHn
9ptX8RGE8DZJlGVJ2biOPuqVAkN0mKOrD+7Aa1j3c364DF1GrqrbMfqImMnC
s8cmp819TvJg/vpCl6i6Fiwip+QDfpIYFPc2hJ71+JyzJ/qppTk4tPNp6X9v
LZ5ZwptfNk+GRmIZzbeyVDyLCh//qNBMXY5x3PRmqgE3WCYcvLgBTCxb04A6
SEJrv+uU6Q6BPBBew0rzuV1zX4etsO6DkK8iVx7JDLchT2aQXYC7e0ZFr61A
cMt6cgTRHnu6idCwUFtqlQ/D35yWDN0fuBMyrqk+suqd0T7STtqy3RcBPg44
FZuASd3xoVWnS0PASfbRtBLEg3URqACp1CZ6Y5sona0vfhBAYLfFfRlLbiym
t9gEgPszelGp+3YO8EGyUc4N/YumLrlKLdTV0Pz1pH8nTW9+zKiiHw1NO7c7
+da4Ii3H4yufu61w9cpyZWjJEAjYfkn7uZ/0uSVEE4557Z2M6XW6XWO70ynz
xTnk8u0Wk6ZGljb8HNYtohsKKBjq4jjauyqrgzOoL+pmroVI42nUexqVADNY
EH+KT6SI+dg6zoOkklQ5pN3fjEhNcygzEWKoIKhAAnErjLfx6XplA4Dh/tLO
BpEpu8B8me+Ay5HQQvzZGoyMzGT2ScMEKGTKOizIYhbcZBDrlVHQ3WmeT7Ix
ME4Z2EYlDmnOVTXqQyfB8twPDd16fr/zqVdYQmUTubfMtE0sBu7EDDDRNe3Q
dVN081g6HbzzwU2msA8mI3pjyUt6q4xgK7NPRkltHCiM0VlA0rhFezurvoKW
0SAmRchmyIYzo6+0op2NTWKJJ9RPTZyKfvYm1sK+h5SvtiJbuxJ0T+MgQ6bo
qFD1+mE2p6863AiAsbeSYlGAqiZWW2VSCQ6uviCYWDWrq95gU14eLVG0YmNA
lebkhCrDQK6XuXFAAOJES4NWTHd0yLJJia80KsrCHv1qrKETrhZzWO+hcFNc
Wlx7dxbZxZKoe51BXtUx6oM6wvoDSgqHgc4dvy9c/Q8xBnXWvYznli/VfUNZ
KVcjJpPcOy7qGYWNfHCdozkYMoxazc0ht18w2w1lBk/omP3xpiGSrUiRIMO/
2z5EcWAqvYznCDUVpoU3EOuPkP7mMQCz4OXiKFCCA/VIHrhSy9+DJADO71zg
vsxGaslqptDRLsddJr0RI5C66nbe+jmUoHVn37MEvd1ilrlflxK7O/N9+x+7
Hv8+TvVRpMbY1pcQt+fWfSIiyBwwT6eucVQZGbFzyCsbiFQ/JRMR4yPdWGx/
ogw7tTsmGeUyORC88/IwC0qipk9Ny6LMFCat2JrjiCiDi/3NLn/MHxZLYxIx
/YAtsO+Kb2VA9KTFqK/JwjR5ArJ2pByoRpjUICR0niC1WnZZAZQ36cjDIkNb
+kr/nCMMr+US7SO3f3XpnG3iARZr/a6lCnDis09coxpOEEGyYjS8c0fBz2z2
D0UHjGV8eGunlOmWquEBU3OB1RdL6F92rZmG0F9fLc4SNpgRPhv3UOkZWZlG
f2I14C9tXqvsGdUM2cqxMnsrUeD2TSS3TTMgejXpmLSRydyb50i2H8P5c800
YTftcG9624ADIzi0YnSHwm5KzeTfdzclm/siZWBYLooTynX4V3MZ2dwjkkg4
PBtWXoa6/ipjCGFO7sZ4DjyhoKY0yeShqrr8jeGLIHOg+HTgs+lCxWbesMxW
gTTXJRr0qoBjKK3kVLLN5L/4WPKLRTVzo+S3JTkf1yszXL5SfQFwmNFamJ4T
nVNHQMTICbFQyW0Lnel29pVcVly9OBGpFb4NtySDIUzWLqdpk9qDzJZIXptA
xlQ80sUbPIjXwPrnf44tI9Ok4YPPzYXSmhR+g0nAseYzd3WVoBpNPjYvePbs
owlOMAwLUsz76Z9YVZD5ALhNruONWuguh8H+DysgE3ChR0V6CkgfDVJjtwg1
0sqh1bLiwOVekWe671bImYD7oYMsMJKFoW6mcB5V+FZyUDzDlhAqgtJtHDv+
tTyeYqeN2FH6lCQCcJpxFy73fBrf+tsHM9w+2m6b3Dv4FqrYot7PqwRml95A
xm6gZvxuB1pEto3GkJgqmwLDm2XYUALEgHN+HS6SYiEh19rCQdcdguP/PxMF
YiWeCIis2kSpj4sQXIjpkwl6oq1gkQIRcEjrHYyJt/VeE5e6rXBBgvrh03PI
DGcB9VMqWG9WA1CJ9nkGcW6onCi2V2WS0in8C8qhZlfF4LHC50BDS1EEScCM
Y9oVcATpS76qN/sIkySNaSBIgMdkaOHhcF9YohFKU/4CY30iatVq+L3UyWhI
qDhDRHREtD3o7sTK9AjVJuW/x/baIr05bv9f0AwJ3yerbeCa0QA9mGjuO22t
fNM8Bj+3etjyzCLd8OOEAdvD806oO8d0qtE/Y/G+vNHXVUVfJgn9k0OnSfQ6
e44KCazgXoVm2a4lp/wpL/azWcrswsmucw9E7vo6YfQvT7Q+aGI4ewYx0w0v
d8cr9tn3cFyC8Qd3vas106H159fGaJTU5Ees1D7P+qqVQE7fO5vQlAAZsTD2
kAkvuat0cFjMtFm5aK6hPdc3qgBD1BVXjzMSbTPpwkd5+d55ii7s3tmL1lZ2
2bfc4tr/TWWHuLoitxvgGktSolgJNuIL3p54kdHYSlC5WKj/9E/EYQGjfhkG
YhoSnmE6hbfqQOtd9nTCfrYJShsP8pVaUFw1fQ7iRMyQYlxKeOtMh7Fj0of7
b9uYqG7n5wN3EHbtZ2Vn7tQm4+ckyA4dxYKmkApDPvBCKOaxmMN4Gk3oqAzd
fm712GnTxrtIO2ElDNSgqhhUC2mx8C0CxYY72LqaVMhcqgtODvUEGVK2JPCK
O5rbPQ3StDV9oF8W1wQvCfaQZBVkDldhBiuvDfIYkr6E89N0BLQqw3YLK3BQ
J+cLI3vCG10R2A+eKulKChnVoy0jgW5uI6+HPFNo3l5REz46N+lW0PmKXYZA
WUjfiCIVx2I4GruxEg7EQeOj0hllZM55CTwuzvyqmcR31DL/lSKIxvQO6dP7
cGTPD9CLOBMuOmmAHv01Efdkp0lQtVdfcAXM+Z/nzDSKQjCPluy48amL2IHg
tageZoOEvo9OLbB+/48xzhg5iu3NP8ap1zhepkXyktfN7CBHT01H3TweffqI
JrzLYDrqKfecH3zyxZJnkxK+XUunx68L2LDFzes7lX04qFjeL2Kyy4bXXOoK
uT/bRxkLA57hnnNTbF+NqSj9xi8dheC5W+LSxuYUm2dKWPgRs4PhYYLuNbZw
qlQHDDoEk0ElKEVNOMyMWbRfEWJpRt8axUW7c6DcvU+3oELLrfX+5Ug18o8f
guxj6bt6JYcKXud/xK1FwhjZ1FbM+KYplxS3tcdnVsOmrJGiQHMZe0pjkkpN
lANYLUfsXE9HdW5Ex/Zryg8eX09RbiyKMUOE6gybd57xCN5nkHYpDlD7CL3l
5Rb3EI+x8GxEsOJ7ctblsFgxYEQU0moQWuBRQ9hntUr7Qj4cois0MIpDy1Pi
SqkMmoZkk1Z7LrqjfHPE+nOmTwOzXFnZ/+QNXBXKFzeqp7PVpEVBV/SgJemj
rgAntBW9J6Nt5N3A1zM6+JjDQOQfVDM87gX1AcbFFG2HzNBOj3cxnnJ2CgtS
gqfenubZIBB/P5KZtNNlQ12JOTgW+KZz8WheH9ND83TNNFRt0d/oGx27EFC6
LR2z5fXUz1yEkMjn/UV6jKqRuIGi3svYZa6626eL+kvSLI5W7rXak3bjjJo3
yMVtv/GZ0uOYFLMzaT2fUAddJUDbFj2OCyJ5q+WfZRwC58/tam11phaVUHHB
ZGEhFjfAdXlL2a5mpD6BfW6aZUcGL6qvVWnc++fGna9VYXzPHr/3Pth2KOVq
wYase7e8x1rlObTiLpKOu9Ul/q8M3hfSRUV4Rs6AbL30fkxwMejuy9qy02nc
yJqXu3k+lkYLyxyF+3zv12zGsRRYuZMf8fsdWsWeO6BU1kPmjCTNoSJ0l41y
Sb38gQMDbabt4Dw7enVxzdfTD/nr+ZBSuzXQUPv5I0ua+3zek+PVbbMsFP41
ST19heH3+HjXoqNlKB8h69OcS2xgDKzXeShI4yGGJJemnf8LYMdVlThFa1uK
SHu/JSCi2x/qEsLVwX1ZEIj5vCYCTKN8rvp1TRUgEMDQ952LVQk5tYA3WwWX
/+oTuBFvrpEuNl9EoRMxMbB74z2G9ZldTMHn+2EcdQo3E1/Jw9CqzBg51yE6
Z7vV6Yao3+4YoPIuB7iaxBOsClSKvRBlaVxN20djNzNUp/n384xhQ8wPe0jf
FO+vJPTCTVsNevNM50n+SajhAxRhZULmcKRG1HruSDtFampjmKFodxSlc+GE
eIZJIyCEjuosIyKFisbGglwQym1B8wfCSPmoDBNlVGmGHSJkSXbwlOQ8m612
CsyftrGRNTJyM7bz+48ci/f0Tnx0MuZb0oawMy6tptRyrVBJYE+fCY21gCjw
e4QCGPTxz2PAjL8C/NAuHY5V2crw/s3pWS6uWzvxCCMZUtADtqcdZa5uqFD2
1w4sJ++STptY1Cz/UpJDxxlz+AOuFKMoDNB0eB2/t2Uj1v71+gYi8Efs1SLS
drW6/0sgJ71ERjdaSbb1zNTegzYW5RX265NBxybxhMR1Dj7QwJltRrKjlra9
xYVGxE0TM5RJRtLOuNJ7VMtTQkC+TjoxwGA2DJ4mQVsoByZQcqehUNLGzZDh
XNJISUnAFluH7tkmEBKrYiSWG6gA9jmQN+unAg85oyV2XjsAGlxxO0TMK32K
whBcdO/aCJ6Y09WFM9wBCSsyHSMllx4i06hFjDOw/584WN37uFsWn/jRdqTJ
DpBYTHfMYwR3NSA2gli3PWKHZgdi5AjJK8ks06uvL2Cabrbs3f2GaEIszk9H
0II1CxRyBCsGK3TB57PVa+KfeeS1aaHabhajJ7pZ6qCQQt01cljSjkTF/Xaj
K4DyC6B9A7DqsPqix57Z59vLoFkjTyCwDVrx3bpJ6CmhT4nDsHXH4GZANHgh
+BjhwRlauMhG1+xJErLqEcvW+KqI+1UEyIXpYcuolmWgHjoX5DpX5OcZChBc
figOWmUmT7tG6Zl4RlXfwC4LyHtPW5m8UFPNhXQDXhIXI0rXcEv41jTwpL+T
nBnNP++/jLmNXNR93o/e2Pb7aWBiNBjfedjgSozRY3c9Fcex0Wlt3AqJza0l
LKEY5UM3nw7S3XKgBUhWe3UaPTDljaiC7zth3cvGYaE4d5M4C25HKT6cPehq
dE0tjjMiSJroxnGnyAbkztfpwNVhHVZQJZASDX/xeh4eABVe8KX2CoTBvPkw
shyA7A3KTRqzvv0FEgd/L0pugSOGEiFPC3FHtfQJR73BFVM/D8JihIv+WGjA
xYFrG3J4oXaz2LE7TUmBa7vUbynsNSWs7PQzU/ogT/RGo91Gd9TjvSm2x4Rq
8+lmfgabyCXBfbL3AaAXlMmt6hHFzbNX5ZfkOt8I0IyqVBRrty8el3qVg1P3
fFBvIDDr81wrHJ6IuN0VbrHvooZgtb9GopgteG9nnMKmKpXSl7KtfmFsWJtn
tVS+UUlzxLrmAjse37K81R/QuUD86IHxp8wvmn9AMvoVovY3VrU2Xgo1gozZ
npngIbzmTDyJh2hQfLgtg2GRbacgMf/sz6LAi8jk1NVcz9AMSEKdmZyUkKLF
q3C7VQIPmUHtKaFqzgEiU6FxAQd2rjN2/k94Wan9VzVSEu2bVxYFGpYkqFYa
nJh7xYwPebbm2xlvFN0DbnSsxm511uoi48W4iJUsTXhfio20l4hPeKk11fFp
zs1jxfboAVxbLtR6Zgv2xiKUfrs15Jj6u/c+20Fsk7nBwhOxq3CfgTtKmp3N
ZZNx4gvY9rOEoieQb5XVM884gO8Er2zJ1hSFkoBJolJx3dBjgSduOlxxVP1u
Pg0eRG1ihAph379R/u/s467ONdNmg8mQFh5JpbX6+MIqiSx+/OE7VhdQ7e44
NLCF6Dc7RgZtteUJGAwcPZqOJMUEbbVZHdIhg/E5LAQyZEgaZv9ITatczRi4
27mwdGORo5F5pJC8aoqtAC8P/kh/MMMfnBCIT2c33tZPF2ooh/YitqbTm2Gg
mYRhIMUa0LFSZpwgGSWSbwuRMT/8nWw0UPOdyn06I23DYasKH0F9OAxwExeN
NuU6LqMKQnOLsu5KQxIE2zCJNjXIrSLWJqGVMIwi/TtASuIcka/d2RyPFFdk
Qkyku7U9DysQFudk6E3QUOex7aYksPjZmErkkzNX617UNjtoxreeoKwXAjaT
OIDnFbOPJ/43ZV6mt7rRVjzw327iOrclhyHLsGyQl4xzs+hN4te/H7y/wrg/
uu3Nb6+sp58NXf/jinRsRg9tEgg7joAjj0IByZBehPAZzfsYZ5tX1ivY2i2B
gGKgMTmUG7HoSz60AkvplqVl85tsjOVK1Z6svIOuUSJ+OrsOrPN5QSvFr/6v
fyORHobUSMzRrF0AqK+Yn5vq2CaMW3Pe90FTeQATitgU26CsPABTsUVcZ+ra
+0VVfp52b1W11rI6/XgEm+L+4hEbrHJIi4McsdqXk7UfithL7T+aKsl/G1Wx
L0WERC81Er4y24HpJNJdIE9KAg7yWbfS7xjHKEGAGimiDJxuqiJHCe5m/BMA
gJh+8eK2Lxa19gaybcPK32TA6jRolJFd5Beae6GTROb6uPsI6fce2oGzgO/J
VkIhM7MgvyYg4UZ3Hn77Z7OmTdVpGlgqouSL5f6LVwmUbBBO7KJjT/Hi5U9Z
5na2tGElmpBlNZynJjfq3mysyGWPY2TfTpTTLE8I04ktj09brVEIK2qkHNd6
Sw1CDOgBZAxUrBARySdN0rHAi7+TG6Cj5Mz5xD4Hz2LrmNlUjzgbNqvidjyf
WbaozFyqgc9gk0kQHivvizn4gTRHKRq3fs63eRXivjgGxtgWktohcDy1UMsA
/eyFFQEL0M6k9O7w8U6A0sSgjnHfwAifTlHjiRX3NfzGkwo9xEz9Z0JWxTHY
dIP4FpdBdOtHDxW2RuxAfYeyEF2GmBuCL/2gs5OA7dn4wkU1DszhA+Gifqzn
ZgEntaM6lj3N+3RSLw539xG70BuuUhOTBH2UD0NCBtM0jDeOId+YQL77NQ5F
1z1bmJH+51N9IcRcjLQuwRkfWFFFt3QQDrmyGW+ASKBMSLxYCZy3wygZ0fJb
oEZqQbsIZyyqnwAUc9eLcGeR/DyWhmJQCQVrqUkOEX6J9rfV2VBBGhxlDyJn
gOyzRh1Pg5b200Z9JoVFCrFl0ItMw1wm9vceAI/OBwy9+vbLBPyU7M1JK3FQ
kjUxVxQlWf1rOaFB3DR1NzbkULClIaecXJhPAiHxgrFMnWvsHkE7nELMqNBf
PsiYxxZFbpXR4JmRDkVNtHtKUUjDa4flUS2Kk7T0+9ZIk0nuFRjKNeHNx4WE
NA5e0ftNBmFiAxmk5XmesKqY3/co4rFq6S21f4Rc/FgP8LZFFJG0VOHr4Bvf
Tu2UFGEJd40QYCQH5rl72m3TAuGHKK1zVPPTHqdWtswJr6gc+doJ+G7GeCwh
89P+YglPISHNpzb/ohGF34WVCO87cnr/pbtrz9sUgXvBGhPnet+TGLZPOklt
6H/2vGSTUiJsVxiMoMYGN2RekE18vlnijS6n2JUKxYgjgmjWPK2X1ZWxSh+q
UCTaOICGCqQ1j2EXrhu9GqZP6CpU+DcP6z+efTHiXBG/ei5sy47qdcErFYJf
FCpf6V3w09aGINrzvvpewFhFniRRsyS/LJifHKH+zGXaK+SdbjCpLVtF7pX6
I174xDxNfE/Yp18R0ZPX9vFJhJ75rvv5LT4/npRy1KsvO0cB+Etco5hyODB5
6tX/CGiZ6wwcVz8nJFnjZZPa19fnVTd0EE3pcHx2R6M0t2dAZ9Lc3OsZTzO/
usiUChFP2sa7Bu/wf33nAlKty+SpA5g6v+5E2gsEeO6/g4pxD5wYrp6GFXPt
8C1ttlWYFmlY/sSCM1eidtwCMjl61dO71q32keHSEF4AuMsyc/IIKy5uTmXJ
A5Nuu+tkES0Yrt2aukpylKDJb0kEyN6KtLhjh9r2hwOKOVsKidsfJ3lx7fGk
nViGTbNiy8s+8YwGrXmWXAQDisS5rSdQ18uxQTsO6TbZM575ZzOl2h9Ly+Yt
kgRetZFZFWrL7E0NPD0ocUrPooGJ8f67ozOSoVQtbbsPxAXvtHLq9j/E/wfs
iLPc4UYhBpgnm7FF7KHRMywEeZAWEzLTC2QM6BopjFrTwbSyHw7pDeMw9/ub
aK29EVTVMk88MvGUD7xFb5IV5uwVH2MIhTgx3J067DaUcN/gy5xPJVToD4/u
DirBvC+LWOGFll1npJLQvCghu1ek87VnOXlCTE75ENNVN/kA+H1EP52pPcN/
i2Sdv2O9MihGCRT4njsrhAxmTLyZrQyC8RzxM1TpjJfAOAqaQy3nPBp5caK+
UNNdsPj3k+kFm/gohbhShZWZs3eJuvMySpY3EHVMKWon896PiCc1KjwDSB3E
lW/HD1X6W1gbOZfWfFhfsh0/A1acle0PXO+Bp1KVda1u9LeJRrh424j/f46r
Re5O6xkmwjfMepsix/pMpI+rRPFX+E3E615KcE6EpPMhOZd7JJKLa9gOn4Fp
s+3o72ngMTXzpTqKZhmi4P34DCJ69eX5vt9+jzPpbqoq3fqT9HoNiE7q+jB7
RjtLIFLHzeSkKQ6T2s51CrV1Zyv462ObI3HdX5yBIpAKzt2dSP1bTkDIPu1i
6HpF8hi8Hca7yll+p52xf1b8/8RpXBZ8P9/ipT3adVWsqD/JguyoGSCJW5Uh
+G212Qx1UsVe3QFBmoOo8Xx0g/1I+rQI4qj+foi4okVToWWzeluO9I5AZefo
P27YOPzXE78GFKkj0mgVJ0g4dmVy+u1X9nUH0tNjy827wQsXA654srGlKLQP
GiJZXjDxMgtrJdi79b2+kCD2kaHIaJ7QA7AtE8g3Zft/sVIpHr/H5tnmrJYG
u9YOaVlA9ISSGKk1b2BBbx91F6AQS2fejRTvxQd9JhLZgJI7U/huPwVaEBVr
mgTrGkCvu2orSoE31E+37VW63cxtFXoxkg2CGFLrYIyTGzDP8yKsAAjERoql
lM6M9IFglqgzjfBevEOKUKIz3/S7EI7jZelGM3IdKmW9bH9s4uSixeGCpblw
LrUcAWbR6llu0vKglBE7tBAMys0p34iFJsdoY2gd6lAc9/d8iW9hsBv8ZTyl
EZpXFexRMYyC4L+RjgwrSFlxYGAvhc282tpZtbYD6Byms9fopXBMn1Q/7tL2
BpnbXH8f5fA+sUjUttmaGp0yjKjRPQTG1pycEc+PucIPCywmDxh87wxwZy9I
vyfyZdIwcLCRyAEoAmv7jTQt5bcDqkecvl7up1AAlwIAE0NGUmwr8ybchIiL
MxwFI5bh9k9NXG5K7IGbCPKCWAvsJmhJZtxKZNYU7hc4l5anzyRgJoopQDHh
EqeutE1o+b6ffYoXls7gNLXE0p45bCnUEEX2nGks+gMC8JcKoRqrP6bcnrfq
ZF/vrqYKoY/Hp8XneVRoHefaUskihV8KvcCcujf899K7bZc0o1hRuBPChMOQ
9OgCurEev07Y2vB1x+NCKsp44Nc/MOfk+Rf7yXK/r8G9H+BLSmpR629vJrOq
JeCsYZlTvMN+FmFsuJukXlkiftuKJqvyOfPgY6YKEwQjwN3sNKPJAqe13lIn
g+t3ACnrhBtTcFCSLZZ6tdTv0ma8tC9NMy42iGG4XuHcS+rcSr0xFbw47xGW
y+PdbPINHTCHbFalvErNafyl6OrnnWdx/HiXG619uaQ5f1Vc85wUYsebNvgU
70/k2/hd+4NgrPh3Fbj9lgM5IfYVpBJT/zyeBCIubYXv0pqYdzNXYN3oD06Q
fdh68pQL6h7UomquiFoUSuweIBy182lzXwZ7mzVJShPYaa/vHk8hZFjOQDER
X/4G+adHlPZiWSVdrGeT29IIBlb8q4tiaOmWcchwzAOODAY20QAnaSTRlDsa
5M+82XpQHYNzXt15HXYHT8EvPGxdj96So1Y8x3J1EnI1P/edwIEtciw1hRrU
jzclnUEMKSQcU+MA+EtYQLc/ojSxLFTOWrkehpPBvtvqtxbl5Rhm52Yrddv6
/3jsDF4KKE0WK3yLUTps74k4blkHdnkmsi1pab1nDNjYDlkdFJqWroqKYTw9
VAyLuto4Or3sFzUCZTOGbAWwFFZwfEwuBkiq89+FpiDk42wu4JTTFdvkhvDZ
ZZLaJEAD1JooSIRcbp8k8T2SSP8R9N09msHd/xyJMPaqwQnKQbgsai9RQ4qy
u6ggihhfIfLsd74Kc0eBHLsxFI4uIHP9JvhftMLyDhPxHKpiQSs7NEhShMjT
Nyw0GuyxFl6ppAlXFiywgW09v7h3y1u1VHSAuK8XqGpfvvpbzmyPuK7JWfDf
VDkyqtVG7bp5RjdTBokSB7pYM23I5BJCHkO9hPdImmdPPzRVj0HQJoUlJz9H
yLgeUkmGPhObios4uYqGxAW/ERl9WIkhhi9DDbm677kQRQYt1USdAJIS09TB
pnzSa06iy3CRScDwC/bUHwG775XJ84Mjsv2L0GxPy5e4uzbYSQrGcZfMFsYm
MMN1VEYkgunch7KqmXo87uT2hGrSudLB/8CecWLUQQsU4Aj0QzDs8clxfKsQ
zXEtSbqctYNUPjLgJGr7qAOOJXNKyi37dx54RlzTIFohr4qUpArrWDtG2rRE
6JV/wCp9k8iZqAzJgl8raU8DKjB1Haq3O0pDF9k/Hr+AsNjPmq5tlVeluWMo
A+4HFivHxgHZmIcH0ZGtyh24oFHEvGgc8Hy+IeaDqHO2OoHQF1NbYMtM+Lz1
gHpHCcO+/53AQaO/ny/eZGkKn/xMYTcPykbgZr+1gKArIjpT9WeFL3702Mho
ZuOdVPRyjsFrio22UptZ6MXmAf+FemrPUrGnGmTDMfzVfQTZ8ZT6RRVPOO9x
JJE4U/kdRmPGsVz/ODnMoUf6lx+lxIvKKY0AuHRgwJrVAzay1D7bWzCO3ifq
RQE8XQzFikTd940oUqKSPeJjRegMFfddcgpHw42ASm5ecR4HlS09g+ZqqK2D
lis5WYQb/ODmw6e1ozu0OyiRcmhJTdo2DugZ941uv4rKvSptL5W0GU61Ckc4
Sk4xRhyJQDlapU5lNuezaSdDruW313Xn3xM3V83hVlmIlSoIYsJAJbJXPyvI
5y4KubRDMaLLUWy3GnRmGh/nVMo930sCNDlNKU2Fg2B5NONeH+3gOxtHoHEn
G1JcjBrC0IPe7KSJ62OCOUxGFpCJekfDXyzQSBnHJaXJLPEXuLHne08K/ug1
7r13z9IWpMSTTjbAymAb6IGJ49nMIstb1bIhK4iikacvRD4aAa7CBiyu782+
0M3RqriEUq27jYIHlGkxse+u/Tr/onoqQu7011NHMQu2bcJ5pHWdGcbyIGwI
QLsxkHUnVvdayKpTy7Bqr0eLN5p79jxXjpzANojG4pStC5/UAV1+w+ZnHI6y
1R0qXH1WOjUXNrtgOw9yRqiwxeJL7op8y3RNSUvfeeAwWOGGtSuM58IoRCau
adHPp3wHhPQQhmf8PEcUt+g1nuTDDKfhtBA0u9iOpJ9EbWa0wf6b8RErxa/T
WXk89hf5eAlFXSPGqJ5GqJXEnLT7iRd+muiuG9byhjWHeq/8ESKiPRs2zMAX
r8PvuDprFVqBEui4QnvR1KhQoFOHbVGbsnpASNLWy/EkMgQCYcK2hH4sIW7g
ZeUPIeoxpk0MvSdbLwCiTiS4z1oKFBBcyjnvgt0xhYfk30pC/zvzRGS0sub7
EwkN5XNTIGAQ65w3GH7ZD/HYr4Sygjp+Wfbg9d/P+xjbUjc9RCKAgCzwPhz1
E8jVCWNLrE63b507XxRSyN4Oicn2ImJh9A7Wjlzw7O0U7MnK4MzaIxjAevsO
S+Uu3KgCGrrWe0YbY4yLqLLloxCxX3rDe6+cHNWVbGfeRutI8Ubmp9lD4oLm
meVr1SytoEr+WQmFWJTA5bLHnMomwnEmpQeDBX3E4AuwHmQmrkyryCGzrUPS
yk9XaQxq04naHqDZk0jfB+uzjm2cO4gXiIbW/2n6sCrkKazT7AYJA6AaQ87+
kabMpNVaURSb5K0qGQOOcru1S4Dvr0ivq+xNv3DGFJNjyhKoHMKBdjkZDW+m
vefO4jlsnX9I22/sHm/5tviyLbgRA0Tm7DQl+NKrgbpIFfVq8knrPgaDuYpI
tB/HWM8eKdnkJAOSsaSbINnZCOuWIljoJPwq7Er67k4/OpsWIRmVqQ4oN/fU
JKiZZaRU2jrl+Jgd+eCnpJsF6EZE7eK6FVpPWSBM1gP5RyY+XtQlDM1zlO/a
3hndalmrhrBczdYZyM1igquPl/mIzJnOFVIH9JnRi7I8kjrHlqowMDAcUtm1
1Mp1jv8Xhn7BsU8ApQfg+vIGcR979kPzkHexmJUabyuz9ld3RaYyREo9lzDi
qfmVGQTpphTnX5B7/nWecFiB3q/dQVcHoLV89mwVeObb+b7Pp8EtdvTwKwwe
L9D0x+37NqfpXPHQp1VriBX0jpT3J8dPBsbWiqwrhC4WIq0hNqznsLF6mk4U
Z8eRKstkXVRpkxLRvKm2VyVHWwszjKYUMZBgJZPWDEiGreGk2sezqkFq4DKr
KOpL5monrrbXCOqYMmhTNLIpQALeCoMjJuHoCqDQMvdAd5q8Aj2Cb8LtOEsk
DDy/VZGpioh4xBSZ4zFJ9I94CA+yGRwWY0KOokpmhukAZsUpHpthmAHvp0Oy
/giohdQHwGcg6YUgntX7bwQQi3eFiU0tyapWyWIezXdqoG5PFEN+ddjjVl+a
SMWg5LLlNYbgfgvN7dvs//MCKO0v+h+7hq/iAeC+Q9awl/aAsO+fBRRW30XY
Svp5HB1RWj7AhXiJO/IHyCcOlwQwzCVbGtLarMrNxkf6HgpoFttrWB83X5K6
CEfr9ezgotTpYlANxP+kmZ1wZZl3vb2pKmbLDJNB5aHVK+tZpp8hfhHInZWf
O5zxiQiizJk/tBzNR0bqSkLAvJuFCSEH3q5ARy6P7orZn0DPPZUBzhal1qlQ
13YMVMY+4OvYT7SIsQOWkAltHOt0kXWSD5imWI+ZJcDk9cVXroJT7h+shZjC
Vm6LjaumG9dYwXLx39ePmxafL8WNBM3YUw/1605+RnzLqZHc9cfaWutC7Ne7
5X13WP5Wthuz+NjaNiEDRrmxj8Hxz+6qCRZK/0YEze3YrRHWVDjnsE0kox1z
8Kh5agDUyaw4zCUBJ0nVQFjCVLjNSVT6axyg/uihKyyKSyehAYgQOknqG1ce
EkOhHMAdYWxWriNOa9ttFxPdxLLOdd1DDFPON4jV6tpoOCtZ2BkGfvyeAjfZ
KMQIMAe3/zOzAEOKj2qRzijKM/8+HImUaguHmEb1bKzabHQZG9be+i+5hByl
PkIplQZw3KwqVzR9XzV6Um7MagTB2tiG5eUEvoRWK7bYrgkcjnpmBXo2B19b
rOB0/8GfE3qAx+5a7MKi8IHxmmFMkCZjr/9VX8ze3fW4mUIa441e5YkA8m8K
a0i4eJHQ4mlw6jrm8qMUwSTPZvBE5+nOXSIS04U2f6GDjmj1ORGQwP79S6Bc
oKBu6FDWebzvNVDo39tS6k8vRj+t3TT2s4I+5PZMuzxA3FUhLxsZdTV8KvTx
MNUH95LUBjFqCJ4+ocKjTh7rnhTH8V9bGmbSC6MzS56F+yI0A5qxOXoXBrfb
9bZpIzsO/Bx0Oeen3hMehzfqgJjz931/ivI7gENCRmvyY8ejCs3iQBVmn7tb
O6p4S94KkVD5t22XIsOZZMyDpFPXhnhPK6L1KyOhSpIioA/T31t0AHkiQ/d2
ahYRFO8Garv6Ez2Yb/brcoYkEwOdtM2LvKBMwLclC0PpOHR314HCUkDEzu+F
+KWLbRxgQt5PqIh5rZJWMMunWvnLPuFhjGz1vFtiP71sU4LRnCugcb1UYUro
psBFMNFxvsIpkr6WL7tT30taiSu2hDzO9bDFnBM+zFr2urgGbYp+baEc7uBI
+kft+gaZOFXGS+yTgbtCk6jouqCY2NWyfvDLg+pvCuo61269c8LFQMZZXxNF
XvzR/yGrzM4BI9urJKYOx9T7DOjQoB/gDGcYUuubWMHwcdSeBJMJXOISvWuA
7Rki8bebtPkopMvR2Q2N/2qWgA5vh4QCFQOB7DxMYKGn9s9Hwm5A1mLLwqnt
bOK+qH9NY8Bb2XbUFAUjvYyaTys+UAL5tel3v52KBXd5Kb/8p2RixarTzIJL
FIdz8Sj3KxwwnEdmG2UDfVeQq+vrv2ybFjACkMhFlqk41QScIK0nC/rCPAtc
KK2eDYjzHX/kN0k2i0/oS/qG6649mGOMCtstBHjFROIfZb9dtt8jb4kt18A1
GhEHeJ2lCKtN4TzwPesIYzv+11BeyXKAwSVMl9J+TK8j71W7hsFfxvgCI6Se
2U76hhtVzeXSeBcfGOV+dToUCZIPEVQSwHE5uRxG8EXSFq7UuxDo8wuyyBOY
WQrwdjpK3LJMauDm85yk/8eoNQ9nYpV5R/mwA+ZGzv0mH8q9+z0eMCTWt6OO
ucVcmdAucX5b91DG7pbv10iVcId8C6G6hGmYpa00m+UBrYFhc6ZbUMKOZ+uu
mPKq13pxaafyR+jFYYxTzM3l8B0onSpMY9D3oUPcrNbhjq1/5RfAVWSWyjfr
hzRuKnjcuBYb/0l7RM5XRLkx7U2pk8SKeM+ifX1IqbH/hBm7Nc3lHQPGe44n
7rt1HXV+5mpPdqoZK7w3fR6HQ1PZQKuK4aanYp9u8Vjt0pu/39Y15ZwCO99b
M57gHFs00JPqpIeEjp1JOdlJ3RNS6mMsT5Mzt9DlYo3NKllotm/U0IIY9TK1
3Nt1behRc842lYPV7BR0xvYVmDrHdpC8HkivOFBUUcrLyZGBVRVkAFE/MDZ0
/ASnKjKBA//qkyFiI6ezYO4+dQs9gt+ZHAFtGAv7PmwWYLVoODIbcsBW3fBP
nKHYXTdKRSIJQVVDjXlG4pyXMAKywM/GPsBGea6BZtnEIAQDjxV7AQeCpzwg
l+dSp8CZVKU1VMbOI/cem1ONGRIiNJZixfrPDr3p+5fy1/i0/WGPNUl4wqS2
fPXZcIJGsHr597z4FkCMgbaoojeerWx6zvWbegMkdpuJlIRi6pknIVDSHTb/
RjvaYtWj6ul7ZQFg4dKCt921DtlgItARQmj7zjGNYj5ZBW6rSlyvAo0YhUOO
RjpW0AaxP4+CYI+aUn/k5FgmuyJI7F8aq8rYzbtIW9MLrgm9rsTkeJJfguBv
5hTXmXorMVGzXtZ3KDE3okW8SkJKcUOcDqC+om3/F8bb8PkFL+e326fxqRf0
z2KKK8sYT695x/u7z1v90lpPjsRWoE6xc5swPDSqEPQ3IsjZgSjh2g6NqaEH
fuXh7vy2AHrj8LN2ka2UNeyHq0yg13tiO6zpNb+q9VQA6FMLqRs2MQDSN2Hx
FnityPfobnsdDPhVTB6gkk3a0MNn2E+5LBO+irATYx7Gvrgo+v5I1HVCc4Ut
7ooTeo3ppkly33oxw6I5scCVFpL7HBA+vcTX5cuBnm4itOfCr2MJ5jLzJasq
wvE5GNAWcaWpfpFoyEvrqkI72drc1pruH6DNUZasqaFEkEabtY/eQj+2IHtY
y2DQ0+Fd7Cuy2qNRa/JMdZh15J9oiJKhOExAk1GhVx5DjDpaccb8wSNCkpe7
PHSUOvKRLct2vFaozAlX44pp+QQ2ITDjRmIpe9rwjaNweyyCMEfa95uAakV7
VJzlmuwJ0RrwedO0y5KwBXNhrIStmxLErkI37vZG/DCBr7Q2WcYJpYKpKsa4
SQTXlAFkW2o2Fqbs8w8EKCHMw/Q+i71AhEEDLLbqQlnJaLt5gAK7lESTDLlN
DlQMNuHn42dYE3SLtQPPuVT4b0+AMM6fOH4OtGdtS0OKrW2ITZUxsp1mEh9m
ZkjR4gNfwF1ooekVVZp7PrKFP1nGlK+M5qwVUdBjyAo4mVwY0lSqiHAAxI1+
xIdUyrlvyboGW6e8rj5ma2F1pOSTjfZPJLNdlWv1zIhIlyc5HQgWJo0c0t9P
10HaWcTP0+Xqv+xLFfpdvbgISQO19S+gf5ksLGsxnz33KLcCX7WSF+dWSqzQ
qQECnNOqYzSayBzTP5JQoMRGI4Vx/kSYhW8myfUH0/sI3kNc+I6jq6bcSArO
c+Z6IXr0fMlfl+hmvU7Bg9yylL25oBvVgTO+ybYxUTdB/FIiiIYsS2MmNtH4
6vUOTyRVGELH0Be8NqgZ2Px9lDdzKs3JZFOj284I3KjgqHv4/Z0qrsXxiDPO
FPTDr7MBoR6Wa61JnOOmO1Usf2MDzUryDnuYlXr7SfwQqIBB+8X19Y2GLz6r
KIEYzMmXAOwV4MTWHx4dkd6grplEQx8d5hrUum/ZujHiX8YplYqR6086lcMz
bLg/Ity4Ife6drNkEL0KEg6v3Ko+inv2edVT3qnQyJ1nDt24EZ5H1n43b6Oe
x5oi6lF5x0p75FmHB9XCnGUQE4Vqhq36h/mOa63H2TfR7j3AAC6ybHkTpoNK
3GM3/h/6BsK3LOpzy9uoCD3kjg3LOdSV2YLZXbwJyRITc8xGBz94Fyc7AMKi
bd9leKFEhgdbcaJpMX0t2d+le8QCFS95FCJ0ZanL7L661MF1s5E45vscmBxQ
B5TLdJZOrTNI2xHbVDCSZNXkfQB/rUcwdR9F6nN0yZjcI19DiocihPRjYe+0
jv+eW78MTq3212B51KfQN4/sS+CuJ5J9Zl2gnLldoSjdgSGNiaKSScHvezyO
p1m8zf/MgtzNX/c/2Rqtn4bthHLLGmG2znDynuWfvHVf6UHlplOv/5XQ0hDt
rN5J0/aKNngbVKxrRMbXxgCHr1eD++22/VuBLQ0azEf82GI2yfuD/wDujN8C
RXeRA+DiGlAXrpDIkqW1qMbvOlHXb4LrqcfMniNc0mNsWBtFEhLNFRhrXXoJ
M77QcZzm3WVO/r4UV+WEDf0Bq+aYJ+GEZ1X6SHvGukcEUpfHlUtAFQZyk/0C
qvG9P4hKz/7pTC7mb9SXwiivDmhgHdlUXyU4K7YRy3d8d7Cr9sd1eiANdHd+
HuRRNAq91SOnP8msGm09IBfo4WvsdUvWhaxETfdIk7OedISKLfJO7JMLX/F3
Ws2+PnQ6uZLqc0cCrB9tdQf+EqRgsOLZOwF7JsBuOxE/tnjSNm+IuxuJMop9
Nq8+OxeCDmDkJpFbtDRqC6qB+KTnwiXaSXG5grNanThzxTYkkary9V0uRZ5n
rAO6ZRf04crT1sctOzOLKkwm7SJfD9QekOVhWy5e36jllcddRBA4buG/WXx7
PaJWDsZXWCr7wa2YxEXmBmbUBrWHVswlcGlEpViyzCVu4fyVulELEVpNIEcJ
hOyKIW6U9Pkds75/7K77aCtbHIx5Mk9AivJfet5CX6HZw432zZOt1qNRj5nh
ahmDqUKm7BTPg252lq+lZdjqrT5Agyxmx7WTwLx4fBQKGk0eHt06BlzJGIam
CYyG6JiKjvC78zFwgzGZ4yrDIP/UT/XUB9lqoIO3NyLENjeOgnVT3qqfVy0w
cxuGMvPsP6T4sFR8WCKnTnje8WHcRShtY6wAk40q/t8dl05LwbpRo+hCibW1
pzy0/jO0iDajKor/4LFKrPs7Nb2teUGf0F3UeyWvLkQwl1iJr4yd9WmzyQkw
DBpOUJHLSWDLZmHJVKUsb6CHz+s4Wazt3cAFUQz0JB1gq50S+CrISTq1CdN/
XVy2WYk02M1bpw0lcAQyc4cVfLlif82+Y6+pkWspYVNbBXfwAImpcVfURJL9
boQ3LGpzQR8Oo6gNXgyA7nUDBVRpjBWVf35DZ5ndIBto4bwxfjjmWB72v+Kl
KN770LjppxQ438X91YkNjVMalwRd1faSCU6Z9+lSXd7w6UU8HiQu/GWUw7qq
DPGViuKArOUF4I9u/rpMYzAsAQEPWA68oaJkslZTTyEIjclXLjbQsNtMaIh0
QSynRBf9J9TRBtu59P0IzzeOUsRYzvMBELxWn9WCuhhU4eOmaEcISpCbIzHh
ZYHeYAl6hYNm8Dc5DxKbhn9lg+YemD6e74YuQA5H+ytCgzgMHnCF4KyTlbRI
T/4ngIvk1GUlK3mPG+k031jfNloET7H7Kj/+Y8t9MfwWn3Wyc1qCnl7WxDsN
EGTIA/9bVQPjq4OZwR5VCd07R8tetOMZLCSoXTdujiAhK05NOsKCdO20dIgj
3RPgHRhHzBUU3Gw0Ue47Fd/wBfl9rLHGALmd+SDsCqpxdY4ZzV8X4eKdQAYl
RGffHDKAN3FiTqtP1avzeRD4DSUdsGPE6ZuyHRXfLE5Kbb5E1fpsPGmj9aND
KzK7jLeg8dEznpoEfrggnyo6IsgfHFi90fvhiTfwt3v+4pVVEARxJUEYJQir
x/mJMEhwXiWqb0YyEC/apyFhxB72o8mNV2C8w5cUWFGEFAR0zTfMroy3F1Bv
97RVYCsvLlglxD0v3WmdqyYP3PAyPwug0Hq03r8+VxIXtDeFnGBtxmW/i6rc
bTTaG3yqnXjTH6Fpw0Hojq7RFslGRfwapNv8eYNLKtamGUppchwfDK5GdRLa
sCsJO8iV7wLlq+fr/lxD8/xIuTFe4XHguLh2MAT8g1oAcstl2e8lTkOkNy7w
yictviNU5+kr0bVBnEybH2NzbdXt3d7USczvh2aWXbu222ZFqNh98TJVPDMv
nkVboO2RYnKx4TEg8BcbKu1wUL4qHywsaJLTO9jeW9mo3j35WHcxIf3qFOD9
epTvNhcLRo94rWw4QEEzpO90oP+TPdjpgcWJLMRdokXz4YUNiIUgBCVJn7Pf
PHfhDHPyYbNRQVOak9xrX0szFs+RdAMQ3eTw5hh2b8VWOQ2FYy11x3JUSm3k
/W5Q6dOlyIVLWEKsD70eZdL+m62m7rw0gANoXJt17NTvAiqndAdm4eQZ9T11
Iv9wiMZrzntD7JP5n8TjSBJNqH8ZdBo3mCl3hccH9Uvc+ZtcxQIsjOaYJQAO
eiz2aQEagcN1PpVzcB4i5yYZheq90bKxQRg+5Yl3g85d6GWVb+wcTqtGix99
jLdAgflKQMYDg0O5vIjEF/8YPwW+TEht0Q7MtIAEssIcSTx639qoHph7erDZ
MvX9rphym/J5V6IWXX1SaIW2//2x6u4VJk3Y6kMfl3EFIzUIMBK27LFvRnLw
ORj84zaPLzPkXtWAh444gOauWUS3ldhyfghcX/8y6mRBeo4Nzr4ASKzP58Qt
xrpesBUvp8+KieVNGPVDZ+RS4jRy7prKcydChokKHKyDVPtckZED1l34QD89
h6u0Ig6zregmQQ/2I90xNR+0Do+LfuOb2xCUFRC0rjF6XcYBqG9tVgS4fTz+
pCEpY/h0fqLbeGZOqYPrI/B216k97WY7bWGO7WTz5kntEleR5oU4ML4k4rj/
fptg6cPaYMVc/xrFvsNhdogqRxddMoq2aT9tsYYfxB5XXmChpRO0AWlmZCaE
q/C00x77D+Ilza8hRnpvvPryrJQ+zj125rfLsnIIgz6XAKrN7qMoPQ1JCa4p
WA9oVbkgvXvwCQz+m4/5FpJOK96xMazeLyh5J2u5jAU/Q+P+XX7d0leMSJ/E
Li8H0wk81dOM6Wb4TIaYZhwnafA9BXQbuflx8gG8kekBfmIlamBdzhfyVK5E
iwTN9q1XJtusThWawFk5umkPv7awsoyL52n8gajzPuKyNzmx0DjKCTggKc6L
c10Giz/eBzY38ECUIJYhLKuPEaZQJhTZq/jk7IG7TLmSnCXXUK6wzxE11/BG
EtSoQJpbkiD5TLcxylNwihRGakF/C7PehKgrF4feYQ4gZ8zXM9TCpJw0Zn3o
xhJDOnb13DKOZ9Yf/0xOQbj/uEzW/onDCcqeFP+BQm1Uso+u7jldW79xJrXE
wHVi0oOvTpleXVy82s2aaIzHrscV/rXTkMpdlRTQZbBS17LyldbTn/q0kPYd
Cm/LOD9basmAX4/PxGBgXZkyGxyCYo281xWImG0VkBMnXnq+A126poo3SI2s
SmUMRrJ4crR3XnQ0JPbabO76JKToOee1C4xEQ9ZFMXBAGl5jql3oHOM62rKq
jCgcA8SZzxPshu1DCXJc8VefnUCpb0yc9X4bVMgGZ0BkrREVDiccBSRan8x8
PEdffyqdcaK79Zub2OjXpcymTa1w3FufvqriGdvC5CI5/jUqBcgITJYmeeJd
hQl5WLK2IfDvSjTh68V/v0ioD0FIJHk8VWV/KxBvaeiQLf1Rh3AjYdW9GJ9v
xlwQqsGRBr9s6t7b2iftVxvXSnayI2dCyo7qbleHrJ2c8HdMDEfbDuatVF/r
GbreRm6+Lnv86W565LJrcsfthOzYPwrJyZ0ciwAFm5LSkjLtwvCi8dzVA356
nkXf6JlI1kWet+g9M8MkOIDM80Oq3h20+Vh7l7GRE5DelN6C2UPwf7/+C6EU
tbfs8kLWfdnrvvZlBnexSPll/BmZyIJfq7Uv+9y7tPxE61MBHgtqW88yvQZ8
8IAnHLfaQ/XWbqE1Hg5t7qHCnxSyqA7F5C2FuPHcewGRz+H5n5g6p3tB+ULj
nw3YCXEMzu4jMpuBfHQm5+PcOnOyzJ9t8KNuBj4tahfe1vPzEoLsokvNpo3y
c5AGCfNiBopzhO8ApXKqOKfzwEXkbke7SaenoISKU/fJQ5geg+RH1kMtQhFO
Z6LMEiUsLzDomS9XGnb01Il9D5lGvRzr3HUkxxlEdC6bh3u0/A+9t8heK+tR
35bcPpNs4ruI0R/vjHfGjbrTWxCyfFfFf0aqVGlaEX1ZlHYHrxnPojO+N/te
C/PBdKrNDjX0WP+Ir9IO3AeucTWn2EWP79+B4X0XpCX7xzCRB6ZbgYLS6Rq2
lprUH8e5DJSbWVnGHV/dqI9HEHRVEB9gcOUNeLZa2zgZHwPd6xh+NYNmVjZo
6tvXfQOtNTe0PYZvdvqd4EzOicTuBFuxyfYNSzlHpQIOW7AyTHPGt9valUZl
m5PGzXVdbeZu+rhAC9kQdogj5iIjgT0XC3ds0XYduTMef+FD4QzxLdHy2rLm
xU2zNnyWM37VaoNXTVqOGT+/SWmjZBP2bnNLhYPl5zpaYBf14fdZ/rCEJ//6
ab7uzg1uiUcn/FvDbUT9+Ufq9XjsTSRIk6Gq0uX+UMvH6+qD3fPODriXlaMw
MqGynW4EW56nloQterJNlSlhed/mxkttin7qgQ9l8Npbn31dQAjVuKkYls/4
FTh8QKk+1qEn6xvlvqr+Cvge9r4TscsoqQvORJNeXySPSnIVP6lIGvpBtsLR
I3WI8Og8b7c0+Qx8fCpuOyDrI8CIKTNbjPrY750gfSuKzI4KvXu52UPEKNPv
KCPqy4lxXeZ3eQpnFFB0wf4RE/uQYg3dHWsSPEEoCZSZrFujzup4ysi0ffu1
quYlDaRgo/eG4k6ADhyBmzQXLgagWFUd51F9l4qNGaPUOEUGMOnsDToANtJ2
CewGzahSJtAWYDvkrAbteYT5hk1RvUWNVZ0mAx7zLUVuEOjqrtvLf16SavPj
q/ZtWwTQimRkAAelcUL95/xysPRs1GClSF32+owBYHHO8h7QqAlTuS4dme+Y
XLeh8oHlWCO2bAMzQOWiEPfcbPyvDAslLp/mugsPDqpWHKgsAX6xm8D2jZyO
Z/AxUI1Zu9McMlWRMn6gH8xgCNNi/vsWChd+ARLYm8TTL0MKNa/a3WJthXRf
oMBkZXaRotXtl+uktxRfCew3xx6MNA1YAtF4QQwHHQLRiuj0DmC1M7I0LTPF
w/3xVpt8nXJhduQt/gjAjCzi6Z3/vyVz5hAEmWOX+eSpLJJ3JPGFqmKcmuHE
3lDGvzJi1SG7VDK+gVsBiAnWOcrzgM8bbEic+1Gu4wmEA8M4y41yHkYjgJ8L
sfC+iiiDY7MBsxYoF8/mrLkKbCVsukTvnhbFWbJb5/2CngASUEnJKm0FXjgv
jG9V3JTEibgFsgP9GO0fVkmzYhguFHIwO5unQvUYyyLCpLSPdF+k7vPZoY6d
eXYXe0vsMYcbSwMj0M13TkzmGf9pEVSB3IK45bZRrBdFFx8TILB9+gEgezrV
YPI+OZenuF8kVUfOgzNkdEII0cKMIbYctVzYZo8Kq/HzVKxc0MaD1WqWRkeZ
SEaJvtrMxpRtJH0mnTawjZCvniCQoGvzwn6CKcuK2V/nJAJUJLpGM3LcPyPF
22HGgJYPIm7uW2gIrSlVK7odcesBIH0u+bLJnYmMpdLfB+GXqq7UcUTsFwSo
PhcMqjow/f2i7t4MNfHL1EFXPVLJVri/Vj9pQ56ZUaeZbfwgXO8qH4bRjGFr
PAsmPPNrF4ZVf1zAIwmeztNOaLlncgasgRLF97o7PT2JPB1thhSN6GYfoyWT
V/p2CwcdAHOKWdAZu8jmFYaz7xhS72rlj/gqc46hJuBHBV1fDl8GPpkKBRxc
M/gZkMXbO6F7/C+fVm0nff8cqNNkW/ucqo8EBIPut4vLtxgUBP807OpD//FR
7f0di1GhN84a8jFvj/tfUc19zCXxaD5WNVDFDx6W19wGeOL+s6Bjtf/91ihN
pqskWpaMdQJaH2GGdkua20d6wUPq1/ze1/7WMMU0/FAdoK7SHv43ejGqxkIR
QU21eqfz8FOolF2t691/KLrIsG50sEufaZG9lijsmq1yR/Q1E/Vd832Dg07l
Tbxp4a9eKG/87rWPANl+NIBUIoMJVlC3GLz6ovmyy+V+UTqNhr8f6XgFkLZ7
dYObOC4OtN/eb4RJoQL7JXOi7ungkD83s0NN6/OdJ4Lzm4QDLq96N5keKnGU
k5I30N+pxC3K8c2iBh+OBYttzz4QZ2ZpRSKfxtgDz7mVmzWZt+r28/AnwkP9
VYULNF8v3u5WZgNF2vdcfA8d9kBrYm02Wy5CzbgqfsdVKilrIANTlO+8CY0+
UhodvBX6O+DF6kn6PfYavrFqiYE6ZXUAS7mi/Wohxe433IcosGKORFI8+Ojv
p39N/6yGdzSmulTgpk3DjpjzaJmb9JUYjH1coQNfvDtyLUhiRwshaEFRWjLq
Uje9ERGUH/j7nj6h5xlMKzR6+Ta7xMeunQ4uSN4X6JSxR4f2AFUCIfEaqjHo
B5KIGYS6vuO7vQ6M8qCtD0JQcgU2n0euxB60vfxQSGMWcKPlil/ZVRT+JunR
vNPq6eV7PRiaBReHJVALs54aTqt3VrlzRonKhiTfWTTXwChMbsrGJvGAReML
NNlYaV4TJ1eB+tc268ULkI2W/LHmy9KIHHzkIgkk2RLpdOwtI51n6ncJtP2w
Wr2RG/ltqY34K5l+xIZSc61FrTa/fmZwZA6LKKoYbQt8J8r+jFcTOR3UWPDI
Akl0d5wNMRM1C6etzgfOJYO7oKja434JfxaU6EyQZgQW3Gla7+emCQYdvc8n
A4Rp9RNtrO3TtMJGVsHu8nikH/9vcp6HECE5fPSnuyvvDUIgqvdEjM8oYWik
f2KI2mkeMSBJeZdRi/pEqWvmiIRMmRS73TPCD3lAwvlA4DQCCNa4UBzhnOVX
GM/ErUjRLDI2CHOdGYIIMXMc6NH6Va8djSV6R/PRylYOT5tB2CRhJcdvgou/
fuFPALJPGNfWsUgmJuHRwwdKbpY4X53mNVmkJ88NXSI9eWlPFMq6pHANywyc
a92FEZQP71MosCoQUAYlyKHPocO1QuPrGWCqIAiH0181lRWu6wV45t0F/0Pu
nnRdaHMrPKMxobaHigWlKRqTTwxL4udXrAa7ScK6hyd6yZCGnV9GCrQsCHbA
jToRtXOQZxodXJoAQHvio8h6lKhVFHCWSJMO+Os8v4WI6e5kUCOb8YL966rn
fjz3anyUZYHWBHbksd2tdMoRT2KSbwIYa2Dj7hkVcL02+cy9D9uKoRyTxwl6
LOJedzhiWa3BzjMwu5BxxqqjH6XeEpgkTjqiiqHbNgQOhUbf9hpkO9UwuPEl
KLcs/gwXq12vbOR8h1omHmMZL3az6YLJJNnbS5ksYS3v0H2zW/8QHob2dkyY
swn1DK5+wgYV/zAFxdFKhJlAFFFGN2legOJbiZhA63Io1gzpCSSYSYAppj7v
23+1i8L59Me2klTt5I/LxkzyZ+9D6r0NdqQFJ7yZRPgIVRrEcNDPcUeXpcZf
k+FZ66EyMzuY/EVHb/NZ9H6eGWgef6HVK5zvE36fQzfc6S6PSFTk+GKbyXtY
AFXu9o67L+OVJkZUT+5lgtmm7zAxSQ6PTozUxcWclaLGxLs/ViDyWCbHdqka
bNuPibHraLhErM8DZqTf1gI5CJV4W8g1I6a3UnaigwSfWkfdKbNOuG5Grxyi
qCpe42SFUKi2FxnO9IL1M38Vtuu2EovFJbzoIVLCi/Zvtx0Qq5/59+ccn15Y
RvFSOQsQPMRz65braReZKBDpJDzkiWinLQCaS6etu1BuV4KBqJ9HEVgqDL+T
MPMw7z3bOe6lKW4NKb666eqy+5eZ7p1+gJ7Na/82bJQeae/DXJDwLT9wSkB7
I11yksCMcvz0LKIbKYCobwxs2dgbUh6b/0eRLBkyuMSiukWcJJ6ucEOn9ZeD
nyqu5L7X7p9WxYWmyU0AqTGBvzjUcZbVM8sFSu6bA9D57PB7H1K37nfcwOh6
+ZawnKws04WQQU9CfC76bgsy2u+5SjbMxTVBPutSTjNzUM3DEjsoHBcYGBP7
Adokgk6tG1bOftkWN9Jecaj3Tc3QX+MT1McSBMo3lydh1rp02pp/BhisLJgX
rVgLfcBuicn4qZwhvCPrHMDqArYNw4AXXnh4RJjMnCFrtAEBl63BPqu8FA2n
/OWjasa9RHzc0UIAzH4YTJhm9ls2u0FCz1VLaW14h1rBVBzcv3+8ychsPhV7
EqH+J/eyD0AxdGejC3996rT5iyeAnK8HaqFUQq23YzzlWVsd5MqmcZsfxUZW
XvPFrujctUt4hWgWI9cTeyoetFHYUqd8oBYIJ5cIR/rARaa2yTuYJTfdzwBF
j92FEqbWOLnLNFIVQUeVeuFnd2wFmrE4VCXyzUkKeKbBqWra5x2qMVJ54kJr
1/zp51jYEdMIwotyZxWzU97dw7w1VL5gvLqQdoXj08pc7LM7t2NYYQH+7o++
/HGyOw0h9HoGCZm0AqEmIJvQa1YNz1MQc2gxzuDF+D6W+8WrJHu0260DQNaR
jGVXouFI7Da606cByjI5FzR2qUTO+YWFNhCWM2iQZmw2pY36lCqatAbzHopv
F3IzJX/pJvBVEJXTTxjsvfckBLF0d2Jmm2FAvg1NOBRGaBzpGCiss/gjN4RF
VTY/zBQtvG3Q8R8syrZ+mVBxiGLSeXdbFIjTNKV4lCQX5dLIx1N12PxHFW38
xAsZ+fUJiiZBsq3IwGqaDABYL4J91xeJxdmmMNXOf3vpdVnRpuK+2mPXDy16
6CCLWGbg0rNEQKtBTVYR83l8JNsBBQ3om18uBUd+omkNzQZN5Yr1NjGOfTti
eCZ3NhvfTG3oxgON7aTLP3y7l4Z+wqLEGKay7L2MDQ+98xLp9a4ETKIij4mU
W48DWDOupbBBId+B6LlcoBe28aE18N58tbXBIv8Kr7+Y8KIcXWz9Qv2lU3Om
LsiB9lCtllnnilGxhPEiQNz4/bpwJAxzDbrXjZKJaaWYV1Dgaw751rPr1ubq
JQdKUIYKhUjC+r6YbpcgH2AGx8padz+qDSEr/8vQEoElpVQP8LUGCkJMZiJ9
5/zdHX+Az/vb83iWDPTS1HgGe+CF8OXUNI2ZE5WYOtXy2/1q13zXteaYGBbh
eOnryYPhX3RQHt1TTaEuWl+QXG45FK1pFSqWjf6dsEcTBPH9QiE3q9SSw1eq
F759iySRVdW/1nWfsjKDXgp6RITY8nut21pxVZrO1P46uH7WoJC3sMdJt91x
jm1+tBhQvHZNlpsYOb8JoW5r2mU+B0JS6Vpvh5Ii3zU0I7ysF1R7bP7dSM4G
tBuyyLMYmWNxziVWJyLkv4aBWu+QeG/RfEb5C2ef/0OsOaU3+Vu+2cXlrLon
9fiSdngaXgtrSE4ALX2hn21Hg2UikDhgsTjtvuQMUyAVMvCyqyS2D4Xyt6LJ
zhLV13ATG6w+1TQNI/ajP3CllGN8wEs9BB/6oFR/iPNCkkTGb2KOJHFYj41M
1f+TTBmOvwIAHJDYkjrhECT7l45a4BR8uv4X9C2EvYp3lKjj62EJsBrF2pgX
9NXQiHBoTidSvWmWZkokWO4pjVlrVYalQu6D88wxGjYnCEP51M576pigQcGF
E2v8//NlR77RvO/op49mFteCmO6lmTh03M0OAaEBxDYeyiZhBwgF1oek3hyb
OdMQRJuVJZ8Nq+VG0VSJoAfEbKOWa7pqpHPWYkVpucTJpbb63z5nbx1KkO4F
qzgEGPVTFWmIV8JTlcdbj9U/o66XqytrNYPyRcKqPRPV6VthQnWvrYnHdYvK
0WAhcIRiopJmGtPv8otZD+EHQh53C5HEtIO3wlugzJ4JOcfteGtxhryIkPVb
FrwBCN5HkfKrKHNied6wSwU2C1eAeIcMwFNukj21950QHwr+MOf7orhVjhfF
1GjQtTo+sw48xeSn96z3irTeIRZ2tN4fFGaHLhe6notTiNecwuIMaoQHPsRI
fyKySdPjmS2NdMadUEl+Eyqxi3mgMEuM0zjudEEsXxze6Ew+MdJuH/Hi7V4T
kgXoVH71dX/Sb24KLrS+GpMfGLozQyYh7n6yJuLd9SURh+WjyXTq3PxHARxD
tn08xT+48uaWoD+wxW6VEo2xQ2UNCUvZdpAcrK+/fJ8kncarRaXbunZlrSuK
ifNNR7cDP3vdePlSb/+Z7ygwVBhC1EC3yAvE5NVjcOJsZfWI//piSCofV1hw
qWdFt1tYEhFmClx6Hco9fMGTDk1hfNKcKYvTJn1IiulIRKtLLxqk9Lxcupyi
Yr1oQ1QXXTOG0azdQxoYk7pDsSKl+k43g4Dy12OLBFQ+aLKdz3eFB5n1rNgA
DWcD1DEn4OawptA8lt5qLyKYqiwWlsdGnElVsKk9/IH/vgo6Zr1rLX7A0yYp
iOwJ9KdPtH5YH+RJGngQiau8N0PAbpkEZ4Oi5ar5kH96dFYyiIq47CwCm7Q9
D8+Qdumbh1hPAlmayXXnuWTHTiotmYXVPHsvbhleNlWeWKAzrvFquLHIyv2l
ayF2MTj6xtZegi8OF9j5+6086Y8VrXGnI6gcYOJs68p5ErBc4bTTfQaIpOpR
zOX/gG68kWMc0H4IwDXaPFXwePJPg+KAaqGyNj1o87JQkPagXlfKCBHG37dk
okqgdB87+ZcDw5HUZq6meU5NsL+YK12fwre8NdXwD2Ao0ChTshjru/xpEOrM
JZQ40Kkx3tLSXjLxO/f00553ZoCforG7IWZaqruohfAObeQm7TTNdFQn3zC7
7n6g4nI/FLdhAqQtbrK198VlBLs6QnDMkeM4l9aWB3cuq83hKQECqB98LhAN
4wHN4kMGj8SWdaN8XD+k5K7ZSHr12a7ZBFCtrlLED3s7FmqbMyDTxGN6RjKB
juYgUg3M/cRECHejoFERPaXxcpMu5bxTMSTGPAaIhJB/RCeCri3hOBcA6fpc
u8HMEfScdcUXrwRdm33YGKOUDzB/8WpxcdXwvyim5fW9YdzDAtP5bdJ/oY7w
gfQHDlEtDcsump9Rf4T4JrOmk9/p6Zaf6zi7cX2cETHVw836p8BtQnazvGQf
+3+7GuRiVHf8+R4z45L0Ra0pTDM6pVtkxdh5KrRgMqieYckMz6qc4zQRCi72
LDDvZTQeQJw42mBNV/PvGtuUpU0/ZAu08uqVRnajyzEbKol7BKkMbDUNctyF
sqUuj7H+jtG4NHLCuVzeBmc5BYYTCPyuMBzxXV3LvLl729J5KuzG5Xb1QsDK
o0UDGpTuHqirt42t4F9dYCGxHsNot/bLJ9iljBOQel0SS7e2hMFAwKHo7nXz
bOrTEZmAD+l1iaWTaDH+6T7Na+8qPv7YbBaqgDttw66Pf3A2KXsNhhUsTpzm
kCYNP8bqVjAW2mPs5MfC7s96oQ0OW/eJq0+L7xj3sw/5zIPnVZqbaEjdoOM2
2nEUn6Q39/hJXq4XRX4JVaapti8VO6aXXMc8ZM3+mxuyiFzNW1UzDmCizXwt
kRGfKgRINmJR979hQ7iQTVzvkmdhl7rKGadTkIUlq879ys2xkpLDqTxt7Cq5
PUxePkOR6RV9cswPulau8BpkeksdA08TSg23zWeKtOTG0JX/vLVTJlIsp4cI
vZuwWkmqXvbkzdu/aD1W8aIfku3bbEwGqVs/XfI/Z0IXzGPc3KIz8QI+nz5q
m+X5WxmziroImOexY2shX4ljVtrv1aP9BCUWaLtUkXAbiP4HtzKL/z24CJRM
ain3nMA4l5QbH2wwG5uN9GOct1h0xRYBK3apZsehoGIdoHybiQmj8FoI/FMl
NXSKPTzzjP9FdmPlh0eFjZnaLoagJ16Lp/5Vo61oOyzZxN6uGtyFs4ulJX6Z
x9lA/QfruftNIZd8QHVCHAznSu5sRK37811EBEQOaMcCaocDo6gcbNPr3AXY
+Xb+BSc3QjLCMfh5GqM71SKlbc1wP2+2ZXP2j0owALnHcdm557CBmoAP3OKB
fpc+WRcTVl/MBghGyKL0M+L/cGxQdihoiokoNwHQMqgqyfntJli+RtNmz0Lt
0XM/I//jS7dLEIu64OtV9Pl3X1rWEP/VgkxdlsH9Ajq2/U/FtGZMpgWYaT58
0dTsrysWiIttQ4BHFDp8pQaY93yR/ba11HpruuT2tVE8p9On/sC4CzinSFqm
6F2wDAuzeNz7W1QCBpUykQ/NBIK4Fa6MM66qV2oKf5mu8aOEQ3HNC28tnGxg
/klsC3dZ9wQP7A1gcW1YlFkUVVg+RbGePxecLtV6Ls2u4H2MajuxPoUBJ6kU
97dTFZ5+oZdK0730N7cHo3wQe7Llfay0s0KaReU8T3MWHUXukdW03kzZYnJ8
uzhSXg8XMe+L5rGSVZ5KkDp6S4yC9FlUk17+qbVp1A44D8bsIYkSfybGp7P9
RAg7lIvxUkAtnwCh228hVeAQpNfAc11rQ3SpzpjumNloycNtCovhsdUajT9n
aiFw3nQKJT1fYZye/fKAheC7VzEHmQIIkOn1Uc7dV8jXGEqbMH4GyM6biGDU
1q28R2K57mr6SXKWoTEd1tScThNPzRryomF2DmBxTkiG0rcSMa2ix08uL4+H
d3ZHOW67ykL4vP2BoiRKaudQvL2zHaBx6rPWOPNh34hg75tlhvgc9zcDIDWF
2Y9QWERbuOJHn7HMIwJur3puQkpV3agM9ZeeGbvDR2lh96ciq1jf/XOzjtGh
bdC3DPGwfMlaGfpZeEsswl5VlgTgJshsADn5guJUltvxW5uzrnTvgcKptZRm
0loglifK57EZsGIIK9ZhIsgADk7JTadp3knYXhMIEcnPW/1zFVG6xlSlHYvi
abM+7nPpU61adFD6xT+m+JokZG7a5KCkj6REWAfuT4TQZzgdml2QHqfl0DWt
Ua2AT8n2aU0nIhVD2eVVx7zmwkGM3790gPP25g9SE6iOgJG8fRMzaFFP/DbW
nvBxFF2TiVzhC78YaotZv8sX9qTq/MrO1hO12QsxTI3l/Ax4eYK0NX7IiYaa
7rRQeNa2voc96f7hCLqBWzdP2gAkiM/VK1SJPEw34wSGUc/UzEDXPnO/HEGh
SQVsuRrRuoev84i+RQbDfTg+SzuaB0URCEyv6+SITzUuEYxX/d7o2i/RM94E
/fCl5vn+kfxyWrhpK9O8YisJHzhLUTXPKjOQlUZmBR0mfyzxohrJ/9TTDL5h
yFaVZOOArSEbDXkk2T6eVtXKJW37L+vqa4L3dSJ8QQ0/tRj9pRFe45TqmumK
e9e1L3d+XRMAGVuuTYD3nlbo6d2/X3tDsTXJM+kWBit0PHJuxPzXo5ZG3Vit
LAKZyct2/9aWchA1RoWEskjOpfWvBdo8Y7ZwGZ/244dsorpHyv4ltPPkgRB4
sLFYOmsrEur8wuSdyQS3RzfVNYzLAgKgxNbfoCIRkU7kING0IWd+cRsVA9dM
9UvzcHIdE1JvynwV3iPi+MwZ92sOScv4i2jLWpY4FurxkgfKt9dGSTtzWMbx
BbFdC0nePHMMo3VIYqLQLSoIRg17f5X4m0bVP5K8muIbFVwrllor54I+cntS
Jg776kWVXPU2CpEPlb89+e/CoAwUmQy/uUfO1BjyONglWOW7GTDnRmM99fWS
EuDFnuz9Ld3c6e5zB478n2hI6quTcH+tFmF2L1BorfPeQsPCt6LS8ywjto9L
/1nWliCilNjx31Ecn08b8O/AIYrxx8vU9dtsCFgqknhf5JY9D9nDXh/WqDLj
qz5CrQvIoaosaMwaWgsX5v84NkZ/YR/TrYfizxSBkv8cCqDkMEb2usovYfx9
7kXkyS8bBj5zdhm8KDEH+6KpHoGeODTD0g6YL67ybRsv/0MOlBddOGeLeu3Y
LwxqgrIdEBbfw0c8mHzEZJbkZ2qpcZDhT63WyNQt4yReR9WTPTR2c1gIT/W2
hWCevWZWBJ3WgSQaoLjCQ2JqksafNGM8VWBBGDyYDgz0MRYXa1JtL3iwFw7y
sjaUS8hoaxr7uXgVerLjAHqXD/PqnY9Cx3BJ3tGXFVQOnqLHt5+yOIbzler0
xlr8hsDD1GJxX+DyoKf41wDtx0WZ9T3uZMWtx8fGhZDZbnYkV4818MDUMVs3
Xh1uPBSDl5KxAm2O2+GTcElITgg+HIM9RVglojiIeh0slvzkOGDM3BdplRWs
5nMJmNwlMJOjtSuONAfr/QDRsuW2DPBzaze4sf14n28KpjyVsICOm9UGBjHR
b5/t4zob6RdWT7oKzwf1nuTpYuiTir6u+35KJZgW+S0ych2ZJ9OBn/sXh2WC
iNO+TNoErs1wDBu5Kglb0az0K2BCS+RvMjg5V+EPkqv5q894cPvlTnum1q2q
QCHdd4mRxAvFQ/pJIXcRmccxMsbvgygMOJ0ytdN/OR4W2yCMOw95MH5bFdOS
YUGeDjY8esoOKEpi4Da16XyRUbxxjDTY48kGjdzT8dp6N6o6eQTvDRH1LDcN
LAceNcEQ13XeUxfe2pTXL06RUj2v513dBHCIhR/SgRdpgCX+nqiHoaP8Bgk5
iZdCXqnB4K2Ccu27ujNC/jNh/lnrvCvYUgGyvG9svB5JjTb7OYzWlO/7U08a
U19P6wWpdsootVRygrg6uJcRBk55H3/NMQo+v7fHdXWcubUfFLxnO6IPYbTU
JT8u5UXsHjsp67KpOPqkafKUdQ3o2vPmRuylaMeedmEnfUwK8r7wNq4d6CLz
w73vFiVSZ2g7Tp434SyRo2gN8wPib3z8ciGnaiRyeNgwMDu4gcXR4OIrY5bw
Ubdljw6uRxCxevTr4ksaMZ4t0Q5M4kQcMcq2FoLomtn1lb1JNl6Em3ErYNO0
N7tHnvfWcjo5x+Kt2dYFpqCa8cxIfONPvcdvPNmo2IHQuqi53Dm/FTJQ9YFc
RJ3+edVWqllAjJpFIdiqHfOWbQhnKftFTURUUuzkMmGCm/jekW6vIn2DoMrU
xJMwsh70FCzxaYOOrx1dBnjZvusxOgKp0i+hM48s7jy9pchvHUwad9Lg3Oog
5AuUiJlq6i1LKfUj2z3NnOxGKvdesCufSNpqYvPz890E9Xr6a9835BIrfiwo
3C0KLf2I+OUF+CqfHjvFRehGmHiNFv9nVtcM2ZznKVVu0BxvNfBiSJk4LDxq
lyGp7ienwPHC/Byjl3b+7iA2Nv2j3FCTmL6TILEf3w8ftYM8KCh+olnc++M9
C9kXeKmvcqvBiFtDG/LGlOhiDS9XTfgYaiHHFiBalz6RGntEs38SraXNIyUX
Qu6o9QNPqPLST7vsb5Xgxjs2FyFm2j3AUMreV2zhKdxcgLdvnk5n7kiCdtrV
/C+Bimmq0xXWC9VVuY2uleHgzb/1gyWLEzfsp8/e4jSTRL3OCMT2yAUbWCDc
gmMLIM3cwapN52f76f9pu88UETa08R7SJzeugApvu+0tWeQ61czKS5vmqy4O
NFawdzjTSwDa0OGb19u+0iP++uno7j/i+t/z26HsysjATV4RHI4YdXLjQQg5
uRXayvCMEi3OcyT0Ouo0T7VG+8Zcvp7ZPoqAEvQXjqN4A0tdgKXe31RTYPkQ
jNz6baIXL+t8q2Zn7LBW3mao3ZBSszk83KzqTVY20hbmsLhl6yPtzlt6Gm5p
Bb7Nr1/3QLHeQHGuDxevjTCNXj6hGbZvCFIAn+X1wqJGEOppv8rYD5GwrTim
Qo+71Ao+r1ZM5I2n+6VodsyCyImhKSW1Ld8XjtVXqy1CotCINNW6euhSP00T
YG8sihBiuraYr/Jp01J31+OilRdXqr6AZNeJOHYlRHc/djr73UvDm+8GSZqL
pEds7tvyoE6t1A//J479Hb6Yh/ZCfRe0840vTRp46mIJOXMrmrGJdS/pvT9M
Cl2NIeQnL6vWmV8wIDv8kDx8fyXljuYoPVNMvLYZLOeRv2TlXRjMsz48JPgS
hvZ0OiMK9AIkCvV8Dxt+8rKWQCJes2YKfjUhzMUlE7gn8e4WIc4SO9WLDYCb
s//wf0kwMhagr2Gg3AiEJYFcn43rx2dm6qln2FJHHq43gyvyT6M+P41e2U2F
e6UWKISWyUQOrQHt7NAkr//ainpWg8scBGJE1I8iifr/UPaqPfmvjj9r+B8R
T6bnyEWXcDZ/43HMRBUO5HFiEDhN04UnVR9l1BAoAtSSl4uX/1iOveki3kYV
C4sgtlGU2IXH7DswBl1r8sCu6Abxt4LultqdMFkIhpQWIJLDhYizIdCApsYL
qNzUd/qLSxtaXi6Rr2HkmFqAC3gXSkNTRRbgxYSAE9F63zgNgqRitHnOJihj
xJo0ItuXVTDTdtTOH50rN/y7/js5YMSaERBVzAj4HjmX0SWGxXWUm/g3EcuW
FFN3ftTavWNNQufit+DcPWkR8qMZ2UtTOQFya8Z8Anb4w9Lz3E08Vli0eD3O
ArSpAvghTPZB7e1wCOK4FHzQ3tGDiZfUFX0gr2YEiNPrNyQe4i4nvWXnramO
08OCAToaLfQH1NWZEueJtWCB8U7zS1gQ7rHuDSAkg6e/dVwUwTT+4EJs5m+9
P64Xu8+mSfSFZ5aqCsYl/9htsFdI+YD9t2CSbK3p4ixMp0mn30OodYQ8uJfa
XohYWT21rIW5HDieohQGQCl6Y6+I4IGIjQeUA/0qgCHAF1yziBh8TiIQA95y
dBdW1Lz0OWNylHe/K5QyV4spnaw3ta/aP+MSL4Ie/s1vWal4S5aBZm35H74Z
z0kVoI4O3b168yRwi9eRqRQH/FuBQLPe2N4pMgjhV2UcqSpKxNQuGOUtN+Hf
naeuT98U7dtKaWes1APRqIT+V9ksN/EldhzKrWIZnhZD6Gd38tB3UeZfnCLA
7716RTsyKpnKvhCCYVMcP8NEYaaRZXOyMAWRSO3YXDgHiBm27ESl6u96oKG6
xygzbmEvFCMBbqb+u6xwJPGlQArh+3zpmYo8S8w9LMeSz1ycNsX05doAWrOO
oSanvzRx1etD9y6wOwXDtIZsi++YoKqNd/eoPm0VlI9BRzG1HCwCLIYtjn7F
pMwJHbsX3JiEGwHUW3bfVd/ldK2FSnUjaZXFGkeGfc83ky1Qo94dSa4rAzMo
pB/436Zu3bz7OGPheBCkNF5DsVMab3+sKD82R2VhjfEfzTPdPAqv8apCQ3Rz
MdwMui7HUH+7rkzvRR+UoiwJzXA8mpOfy+/V60dvWzYytOLQwbA93U42gEvr
jB7T+r0cD0KYrw+yYIJbSEP8+3D35WZ1owuCtzrYyx1sAPrp7JD9oSKz4TQZ
thS5pC7RWdOPiPEggk3rof+IDeTSBokZQu3ZzvupdmiFI3YkaPeLMEm0OAbM
o7JYfni09I69udn9pn8GuBMzk0ubxX61JqLblB9bVqnIhF/DoiDPhWby2zYr
RtudrCcIlkGVH/MLTWvalG1fWXXxo0mUWODRTgcF8hjyLQUC6lZtkYrZ/z0B
B5AegK1+6SJWTK9KUyVSI+vAjG0o2n3adULENGV+Dg5sMPjYxbMAFINBj1h5
/J8BiI9lzqLOf9C30WBxhxR8piyANNEvPaF+9a0S8MAApKt7pidt/+ygpyT/
nt1yHUV1meEgaqQb0G3w8++3XwiC3Lxwt4iEL5LafIqDtfANNVZQywivb+bw
TiCK25bv5YsjzPVuwqeTg3YGfBz/0ywKTVDkoLtijt9CE6/RE74ovPdMIl6G
QiED9pKHjEJXh7IdrAfcvRH4O4TfWKprZq45wQ0O6vB1Blwbt+cGGDG6V/Ux
eN9AUhJ6N35VL4tY8XihwOThQqL3pH34HHFtskl6gqjE9HIcWQ+Tq3lSzerI
3HqR0Hd0uSI453iL6iTTsDMVV75o6h1ZISrUEgYqy2vzWF4G3ztB0wWfzibB
kSDqFczsYeAtD9g0RCABS3GwWX6FwbZg2O9MJksaMXROJBAyA9bI36r2ytoV
hHxOR2DWeqFZgHYREzhuese4fR9nnRdBjLTn4qROGNDErheeeyNfYRD/k9Ax
EUXJ0dje+MUI6vKlOrAinCZ7VgLy+ZeNfOS9yk7TtSpnr6QVfVgyu4x5LPi7
rDOp7sXeb/SCb/5eV2td6UjA85ygqcdYTQmvZ8qpvZlC0/p2YlDMckVt4MRu
Y4NmoiXzeUZ9r4WOL/NEfzVrJLtjAKS3C3ZcxVhZgtIsGooXF6ylRA9f1rRL
Tjcw02bc7/q/RjDUJUs4Inc9kmk76ivllnv4LZfgqlMi4PlBZAzRhS+Kwi96
xXewlXMLMU0sYRaCUEFbDo9/3bG0bUyA8X6dvkM/TsloX4M4oNc4QCWLBTXP
Ytuu8IIoORWpKgaqWqaFH1yVC3UmLQholati3LFn9+DEYfJ+fXOVNCjikNk4
Nk5nRzxQ4WUss+cmBxHUKm2S137U/87ltTLiXrIFNRUBGFH82CzjVvE3Xz89
qeV6PTBar24Q2hGrMzumc/BiG5y5G6exbsTPzmsfu/7xeQji5sULDKgsYGQI
i0SAhk1xJW8RTwhFDgvo1u92VNxsCvUi1oCL8nxiAGvwmCnWzpHfBEk5aDVo
wSAh1It/Dl+oeASgHuv396NM+ntPKrUtxCU6WdiDx++xHYGDQoXs4g5tIVDG
ijX3l0u/l77/P9Q8Lgb2nqy/v1YIu1MvtPQtxakQkYFpvh06SAIuWc4V5xMn
Ew7Xl1Hsf8cDq9cqfIwPI1wIDc4cRAZgqU+eLV5RlC5EloxAHKczzKJQs8LQ
OFKt7OlVDWvAqoK2qOxWEFP+uKtjAOC5lGCDysGf4H+52dSbAHfEAX+ft0wA
39duJoX+WnO1gLBve9JgrZdGs0/pzvDg5km4fX6gDy+e0GWOTePqlDZbKIqV
d9/UGIZ7a/q125jxMHZIZlAjLvE8cnQp7c7wGnFAnyqxlk8edjDnjrHNxvrP
cLzwhoKB+ZnTo9fYap6IQuJCFQtGIY4cMnnynXmQ3W730jMHy13vsUtYuMjH
0DXf9EWLjnjCwGxIGEzBNj16UkW36+1VtFfhNOHonC8rJWWGsmqhvRMLcyCU
sMNshuhO7sEYjAbR86wzQWCZN2dh+lHxMOyxPYb5cP2BaHkysdu+KFAHrRsi
xr81dQRr458jDTeIxLZ6bjYfwSMhNbl0CeDVrLzMUCtt9rsVkiB0d10Egbpe
WOth1wfpmeLpOejX0DvhVV3CPrLnOuMoFQlvJGt+psvvobwg/sTpo047VDDx
rF3ZPlNtlzl0SStNhBxCK9ehFbN3m5GRP706IgG3BqgHR5KSADpN6sS4xNwZ
xawyuRY6b4ChLRLfDGuwp48JCmgvSxpgQ3ZsmjQl1DJrrvD+bus+e2b0wEWF
XY5HThdym5fZWufkyC4DpXGTJQDL66AqV/Z59PtYGL9WYOsJkzcSIS1G5Mc5
z3Hsr4/U9LEjPnHes37FmYQRcBKE/c4aNEPlE0+ZNBH3wWA6n74RBHxgL3ZT
TW2BHvWNpB48ii2s5KgMq4oSZvkvg2Zp34wLFYk3tFPvVJyRaJvXOc3NygaC
WevdSmL0TA+FS6+plB72QlbrYHXEK1FyavxL70ShTdI/Rdn9FXYO4ehhV0kP
61heM+PBcBAYRWtyk8IbzhTo//fkTnoXy7A5P+iQM7bxsLjSfztTSn1Rt0Y2
X0oBs0F+180XEp6/R/I+QaEoPTaH6AApMNO78YPvEtP48ZhiHT8Z6EySM377
0kIOME0jchN4baVqimR2ICCNFBU2ghHiVL9RmM2uNd1oCDWdumR9vJiVwndq
oduWA6NI9Kpqbowu3lNJj5KGBhdmJ+pOqzHp1tYuMKgHGzjET4umqAfNsFSv
5w7SeNQg5LGLep5tRaM3sgjd6jTbre9029iSf+DNYwwXyvQBRCHgEgLvC+If
s6SjBA3Ux356re7uFspSPclT7Nbvr3yZlIB5fI8WYcwvMvpS7NdHkPUjcjDX
9NZ3JdaG3D0mzbOxGVkYUzNPucGk/kaUsdXYXKZLfrEJToNzb8oHsepUQSmU
W9wAuZHgWqkjBV6vmtWuUvLU0i8qloqzgZrIcAszxhbkNXmCv3+qrUbonNYO
VgUF/fIm5Kyip4WIW6sA5Pf32Lma5AK/lXEGYMJYNxBoqkRk2Pyufw17oam1
/VDTTXA/eM2WKvPstH0B/wKf9P0zcXdN86rItFaKb8FsiFzuxKlIfgoeKY/4
X0OqA0RXaEbxkYpYkZBALKaLcdhBA0WZcEJcHDx6Gv9abb0SFmxXDPR77vUu
zvGIZi1CVkeFPj4FM8pgqAkMhM2g6b3TLsPUTTDHgvHvhEKpjbz/lPXTMiEl
P1oDkuE2n0bim9JtKF6Pm8SgK4R8QvuFkwsbqPRbwxWUpY7GYaDy2vyN50BJ
LI1ekVRrF7Y1iICl4N5snH7syZTzWStZhOBvuYFFxOtNcgXO7K5IZFhkWA3m
eZmmVp+LqI8rsIeVa5UYkTjjlHkdF6+o10k5UnnCGXkhxMoIql6P0/Eo8bte
wtwJplIlyPlaedIgvmUn5TXAFPX9SnTXVuSUd7gxLqEaFh30TV2CNM497Cq6
FRgUahaCqodzFJCHKAdVU6Oa9OmyLP7RD4SB+yYYoRHu4jmM/Z3/SeHTZBNT
8tJtkEVQaHKSjQtTVmSe7WbsrF+c6P418RW8aJQhytmNxUVPmEdP4509WhVO
rU2l8uWij+o+B817tVZSllNc1bghVBNDF9p9PC1/+uEDMbgRhIGhK4lYFzel
Y/UsA131o2eROTYvo4Q3j6Lly5ostgyMbee1CpJiX1pcXYHdOQX/vaQMSH7I
gRDELQhydzhbm2+LKiMVBJGkbj93xe11T1Afq3oz4wwp7N4hKcczHZpKeo75
uksIBgJ/zM00yTraB28iMCuzlr7y/7amvK6RmqFG42RaHFpZwkACVyq2XMlC
Guk0VFIdp4HcybBFp70isZLhM8L+ziyAE0WKTtGUrIvcWcVXGF8ppiEOZvxJ
K5MARNQfORwLMnoPXDq3XO4D58ozXetIXswnHQ1d3E+pMvXb6Zqd2ZmxSr2o
gC2FgqrJjuLKlPb7ZYGy1tYAXLUTdEaARdS+Gq10+IvMqbHIvDqDZb9bftUx
Lp27M7kJPpgnUd6HwGAsP4UPxE9euzB4dCLw9IAlcdyxzgUOjSBnZlNumWca
wxyzSZiSzfiusdQTFGRZ/GWh9dQdJwmfP+sNpXON9r/jx6MPXAo0AYxS/NOh
Z5eWi0tl5JKEIsQiHQoJsVbaSd+iWXOl1Gr4h+0ZVgYZG/XszyOEzkiideA4
lmr5+QIy1KbppnoU2gs80HYrYt8dMLEy3Zg2uFmKmcMOPGoNImJljGLnidqQ
I9EXHIzl21q4URERG2E4Nihao8r4uJ1PqIYYPb+18smCy6RMSXBXMpXV/0+1
kpXgj5T13zpvKGo12cDKP1XdeTGuBLbyAC81ohoDzKaR/3q//54aNzdnEO9q
7TE0oBhzquZtaPTi3rnSrDS2H5p9QuLxhgAG8qfUF0ZlqaddRzrCKQwyD00l
eNe/HQYFUzuTIylL6TbwVGBjxlFWut6VX0zxvzotwxgO+t8a527paLphOw+F
SAfGDtuDdBfAQI+8t+UIeGcFQG1bwHpywCXqP0PyjspBy9EF4Jo27BuuLbmI
bJ1MtA4GU5xs8MbqwDC+2jPW1oGKsbgQz2ekAPJ073cuhwtQKCHX9Bm3rQh0
kTAHw8z8zgEXGTjFopUr0NH1iScZFjxntCt26TRDHLt0OSsDthkU7GlbFK8W
rGNxRccza+kMQG/j9Dee861JYZ8wuZGUMUzFPwIBHchH3/23E76fBHneLlde
n9zK6r8xeAsZdUqH1XzoFXCtKMGMJh/YtRqftRQSmfh9gU61VfbyN7zmWHRi
kWzhMo8WrrzJsUCoXWnJ9ncjH6y+cftOGs7mvlofHnBrqHyzhr9FXZGFESoL
/d7EcMWryKCvhS9f3F3PNU5lH3xIdqixh18prJPE+NIaY4YpAHV3ugYc1fxZ
QW5AB4sYZ32+XV/9WgaTC3WjnprjQnsR5wgeL+8jmKIrbJPQykzYElkhyDSb
s3bqBkjxg3CmK/nKzRMjPKai5h/K4g9OyDr5t4HiKiuA+QXgqiJj8HqbJ7/g
qyVGvLBfKLpxMbXeiXj9ecwV9bfCU1dDcsvJg/TzeT6L+l+GlFpUDDVAOCYb
OJaNYdbqRCgpmzwWBdlGqyn6mfu3h+3/9SCcLCpruMUXY/hSs2t+TevkgfD0
Clpygd9epFlBzKejXKbIPVSj65RZnFI+JM9Fl6m9d8Om2seKMO7Yah2vEGRP
KR2rS91zfcK4Z6JmRx/Yvu5+fQFipR8SOrpSTCPKIpTxCvQzP0jh3W0veIO1
E9oGtsFm52U3iLaYfcbAurOsW6CjCJ2RdKH5f12Lrmrnjhtdlj6DNyVeeMx5
HxjnndXPS0RSIGevUObd3KpLD16dfGZ0bqbe+X7Nq7WwWmvi327HB5GCWvRr
3CXCwirGtlXOblKQzRYKuK+oFMsqgLXXFEOTQC+jFYw81cHTsYazgfbkWW6Y
JDPOhiDa5ZyXu4/wuEJ/0MC2DVmkNDzVjj/SXKheL18YR3eLOykXw9AqwE7V
xOz9e8keZAi6xqJIV0ml5k9PmFmc050aBRXWpTBEIOealV7mAwCQqV8+OolQ
0feUWe6DRGkw8H1qnovwa7wNT3DqtwpzC99B1rePY557fWMPNlv/W3OeViQv
cbOPQ7BARG3nqtvOxqaV+jOKLu5Az1iEbTaG/13iEDQwfm4dL1QEjgw1Co72
/2cvB9s/OXStMqqnHYq9VTW0hrrumFN19jYmkBaAWN9z7reE46fBUVu7T+y2
YtAbHo8JAbtqIwdeEU8Ff5m3ZCb/yjPDqzcHpjtmJVURddObhOubGFreziXF
WO1VJTYUB2uGAvT/fxIvZqSulzQPMWqihuvkfMu/jhsQ25g0/D6V9ELgHvhK
RSEhE32eD2icSbUKQzROzFbmnl23HsTIzfBhTyVE4TpOj+6S26L2LsGiJ7V/
KhoiW49PoDOakZKa6deMMZb0MIjNy5zwgZfEe0VXtNdm3evrp3EgjKcxbco0
PnqGaZ2rL3PnwtvjxP2rsOn13aW7lyk/5UDUEuWjSg7xxvtJunErWxM8Aym3
+o2tXb5Xmeo4gL57DfWlRoGmIo8rVmnadLMN8CRj36TLBMMEsZnKZ3Fu0mbJ
zDXJnAz6wqH91ArVJ9QCyewoqT+nD9yRPm4m5PiOYsCtksVc55RPCJhJfA8r
N0L9ch6o+UtpFtZdPFkjj/tt/Yw31eTtAaxURdZLrjS3YSz7+pzCGYK4B9dC
/KyM3c+yo4EMSTPuPH3oA8g65vJcFEuLXZ9YB8t1bi7lc6MVBwD8km6eyZ8+
WNTdtSQFv4rcsI9Kaq/SAoxWou5ercjh9wgV1X1XibIGOQDfctRmYXVV3Pn7
f2sGlkwTx6qiBKWbXvYKbh8ElXWxcMFS8WmQ2aisFtSYO4KB//1ofuWBfpJV
BdZsFv8EztXkimqRI+IMCMh4yYEKK/oUSKOCvo9xQqrRpTps64hNzzhSa6yK
ZAUvDoCnD40vKzCE0EnVxY71bt9d9kNHGBvUqsNI3+SwyE1b506W+ogg5jJI
oKGZ3rrlFZUHYw22cwJITvpGTJ3QKRqY08h38tJ8K1D+hWPKOy0q5ZF/tOVU
jolKWnae19upVEmtmvERySIxesDlwwmdoVh6XsqmjO+/Nhp1Tgtf5iWyU3BU
Zi0/PVetRkeaMZ0bnaueqCIajEf6QU1z62hT8X4ZOPcUCLSu95TDCXwjufGK
Jj6/oglYqI6/veqb+UTowIYnemAbwMWk1kjxOiDcsQoU2vta4MWhhyzVYrWE
5gup136zKI/ZAkSkuJDgIuZUsywTYD3G1wdk9nyb5ZGPN+9x8qa1G9EhiBSr
RyfioSayJUJVK4im57UbfJRk9HibTw9NtzLcuWpoHFRBoN5rcLsxr+h+vz/T
aUEnBEXQ8na0O2rvsSkqUybw1YcNQnoZkFwWt+PmoHE2nYrhfpINCqhJaRyv
tXjmQEdGUVxp7Klfd6fGgDwVje7SUN9lVyxSXXqAzx6uc9O4aQ0hkGXFQVwE
w9j12T5Y3aEH9j0pZQHKTbJZyRqHXM6Omxpoci2aSMOlZmTHuhA33pgX+YnQ
ZRliTkQpq6FX0VfylUFhF4gRW0egdks2+qpDsadz9JjEP5fEVVLDMHt5YiSc
+ocOFul8IWYb6aIkZ9uGO4+U8kYTs10F+BfhA+u6W/iTFv2B0LsdGnoUevEB
7lam+HweQ9EcWSOkJJkFHTX5U7T3SrWR1qmIHhWX9wyaPC0GsGuOavsdSzG6
6kzRr8O2b2+VRW4yT9zCchO7SYGaRAI8t0gBEE4TX9gWEwQxK0tPeqAHE9rx
Qt/R6fsCKFf/LFox4hVp+kEfJWQQluUgYE1PSA8WsDnlratOoC3D/RibWDDM
f7zuv4uJY+2qvPmLlfOUALvxg9/3f0wu+TV8kgh838Pc+M94O0G3xZHGlkoo
OyLID8xhPPTv6/CvRLE93ojcYahQqNjtW9+tktnoLsnAZGNbUMJRtxbpDbMT
guXjgOsgBJVIDiJb1GJB8KeTwyz9QZGC3+A2vXClNOFBgjBypOgkkzDCy2OO
LimA7xcMO9MvDRuL/FR3AV/X3yOQ9aX/MqLEA0wNLnMQLXmrL8tSG+pyKZ3Z
ny124IqEcGa+Q/KhNelyrDCTXG5yTPO85wqn3JLasVfrqbdh6EVjzaufnnDn
YYZ/kLKtWEIzg5AI+S8xtHIAeOP8oih+kmAk0sSxdgzkh8+Evr1AUlLooNBb
HAn0AxhweeU+P3H3ejA9/IhairAYT80sWU2G282yUJ+G/3OQdbeBgS46jhMA
9nxPfB2fJvohldUj1TUn5Q7BHUTq1Ht/3TvTDq0csDjTs0aWdpkwx2TjJ9C/
CaC9i1d8jlKBJsJZXCVaMV3adx3u1T+1PEJsfP5Tj0DKZPg99UJv407XtRda
l6vBrbPYToo6NUsU5G+d+rubOljW/wUDnJNa5vJxG6ESHkv3tMCW7I4jcmQ7
0IOZ/KKFOJvRbVH4QdwQCzsmCfKfiGeMZN8xKLwrclTWNyS1v0OHjsPVueC5
EiKriEzRqwYwKFRVzQlW9G/touvaQq7c5H6AvRvzfaO4IahYh8Am2YmVyEv4
4Yfv32NTGswRlcFb1GjLuXMZTZifE+fskVKRHGrAJheCuDqihj5FKw58wvlm
mGtuOGkHLLZJjMYXWUwukGv6xdd+bh4pNMyi0GBgTIsd/OKWx/UBmlq8TTzx
1ku8CIpV/mRpa0uMAJPa0b50xbiPL+hhX6xhQexjHyZvkN7AP4Z41JNPx7wu
gZHr1m1pGrbxcw9Tl16mdoh63+r3HertR3D8dxZjbRg0VN1hR6TKE0RGLNoQ
wOFbmIWjWD8ah4kZxAsXSicNA633P9dgiSNmgy/SwjwoWgjB7uvfa4SVlUz7
0fN/3a+tyWL6S2qoKZQRVNZPQoHO48AiOU2XAIlaZPqTswfTUoXkq6vXqbFw
6yY5TTIlfJNrjXWlHLqu6a9aCqbqd8YOJm8bSOfLciGTmHiMF2y6fRyoOtEj
s+NxW6egN305RKHfa8kIelSsJiVedzlkMlg2kPCGjkTGX/ts/qdrllkHQSTt
/XP2FlwqcboxuhyqoxlZ2duVVXlmskjlOjoZGK7dzYILrvdR99u1+tn6bSu/
Qm5V1jqTb/e7TUaZ6TdtA0UDYKRpQci9NibVQLQ5LKYHrPoCt1bYA5GBy+Lh
P0BUUBqph/uZmmA8quB9bzquXpAe8R+4tjuiv5JAeKfPG35FtOAcBxDE47Vy
j+HpSwP/9OSnx9UH4Som+9XKX0KYUzm1RI3IGciR9OFN87bjIz2Tf6QRo48r
65A3l0urKTza1/F/a6I0ofkeBvMfC5/YO83323jlAPCwOgq1b6j5vo7cV/qy
0iYQoBbv0MOAGDsj57CQswpkDuq0ttg8x7Ps4U44/29iUej34nVu6nJigZdQ
k0VCjliKc5KH4kJdsauGNqmfK3+hHvSK6R4TyuWyiBNr1xDJEHXR9kuFgIGY
fc+KKxBonXg6XnBJJENV++UjRQzJpfRXGwv02KoyP0Jj005eLEr5D38L2CGR
RPKsEjopzUYjlx5HFVwCNYgPv4B1Bt+HNgWEfO46qlToDrnlK8E5W8BpQ0Wc
ajqyXUcMRTmMyf4MfCq7DoOhqQhSAnaZZnYLAiW5k1w5Cg10lJIbXSdCRbP8
Vhci3s3a255/7UhjUx0cV4fBBc5ArKhJ4ekCsgqb/bWi9Lt2anHUlAK13EaH
uqiPks4inF+/hvRyCPri7pKRgqMBy34XZK+pSuFWGTX81d9/iq9IPfY4Pphf
iN6/1lg3hYXYaS4mGMEy+XBwHJ6CvrkFQMCDr5SAMhs+oPcNv+BbQvwn2Wrz
KK2ACMlIzWrjy8PCfUm7M1T0Nq5SfqrsKxqMxHW8if1wATJ+h3aBkTPtYMtk
CI1wVVYO4a6lrTKx06dChFPecherx4WdBCXwHasLrAU9vonorrDG4GRt+tVR
Bbn0HPe1cE1dAgiqKF7uscULoGONf7N6iTqP+5dxsm0RpPcGq5gOT82EErA5
ZnNurvHhxok378Bnwr6aVw4fIq1bJ2JvysPFRJTnh9f+iuXIrSCHFwQbYvIi
BuNid84Clgtuh93/RBzK1aQo2p8rKzWD9PEg236Kqx0y3qVdU9tpWTEWJ+gT
RiB0Q4oMh/P5CYm+FL2L56zw1xnoUIN7zWJSPaawnRDcOjq+BsEy9mzfoFVc
Gy9/GdKGeazUEiRMe1LRdXK7Hkg5GZkG5MTJSrGWDr3yL8s7/2nOgk2vFTao
NCPjcLpVCSqC+4EztaRkn5s8MpbYNwkXUf8cnobPSWzung4dkf2J2VKreCCt
xJl0QtwB68DP6oaIsBYlwytVlLyz4rrvw57DrRAaU6S6zs5TEzz7mOKq9Pqb
JzechtsKoNPOA3SEebRiWvaFn6YVYfVzENLFF8ttzSe/xmbUlQzSdLZFedrI
tDdd4iJHxvF1EFU2dseJSgoqbkrwmL9YpLTG3Ap2O41oovC33N0Oxuv+cqaV
Ke/bwBr4xkEzGw1k7tyEBNvCDx+m5q9/Ec2JIAsPM4p02nzbPicjLeqbU5O4
i9LyBJbfBNSUGQgsr6ClBARapZS5pMT0wWD2NEYVjNmeycBVEVIEVT8XoBLQ
0Hkt6rcN5vNMxzNJ9zBxto7ay3qHk7849acEL83mH/xraT1LLNBNXpu0Ta1C
F7YWG3YJaWsZ/ST4Ukbs7t2xq4xUH3A8iKMWrzeBfxOiNZxdZGr1T5wArxnr
P1eintOmyow4DFrzhCZrkpuU4EDdZwz92T3ctybYg8QaXz/oTgYVHF6UeFux
OI3KWauamlh2CT9dwhF7PkKb3jS++UBoT/tXl7KjC+XJ/YCwo7fDFzzbEpyA
whUvuwdljB6vN/7Qv2M+u5crzYwdtGQr/iXIiuUPevLOzFBKkZbK4lII6P8F
Dw3Lxko1e+EWJ+GSNE2+Jq7TPnrz3d9txKDCj3xXVh59Op2rexnuQZvGmfve
DlZBMt85thIgd2/VOhSyUDTd8lGvXwmPowro338utykvHcjkDZ4+tBWMn0XL
nQQxdqEMisxxwaA5wAjNvwHPf7OZbtuu10BW4quVfmTu0z3NT8V31uKXvnxv
uALen6cZak0eiy4DFY+0OWBY4ZWnDQ0E/0EbyVMPaozWDd+v0wvdmmL1giZ/
co0b5j4zy181RCc46abeWi5kyeOez6gm7YpA5rAP6FPGrEXRAiBSp1jNJGQ7
t68jMSkErQ6tBnmMRmt+ZpRfPi3zC0Rt3kQIQskdNDVd8ggyzaHA02qvL/vw
BmIRFSLho71zSF4M3H646WShFy/DEXYLPhBpQ9CZxDRLjZ/mzxsO9x0EA6IT
Iwfs3Jr5xtw6QklLXclQ9Zu3z5eN8GbPxQfuO5uJomt87PgA2Tjq34FJaqbL
t7xE/vyfffRuO+hPSy4N09xavjvPlubH/XeODgHBWqzCkowIYsddkjj1RDGf
P4M/bKMkx4cOoZ3YP021lHhACp+H7NG87/oLfc16xdQfQWPSUheflppg2IAG
ZrkOWqI7n2nLAAgch2Rc3mwpEAM4M9Gf8jOK/TWgKFsoaFL70/88uU8TGULV
cY5abAp2AWUZrBKBjTHubps1Ycn01xc0WFPmi934GFoJrcjZnLpKxepNEVbp
qa+/a+qL+UN/sgAdzr7miKQpQOtp/GbO6ISZBuIOJDtnB6+MCeSoXQDcg0uD
S3T+kwNhsTXne7KK7hN/Z44Ckw/ZUFJEAzyZj+FYJKUpi3hbYhTEwm1QbwI4
WZBeK/hJJr1+MIhU8MLSQwMMa5u7Q0JYLLDUKy4mP7lYE/gkmJTU0JgGt55b
9ObZ3XR6E33WmLf/TYS/lC+5aIZw81OYHX4nVqqzOdm3VM6uuJtu/Fg3hrKI
VNdyhZDqNvXxvgWUXTgMeH7Hl7vtfrRgVPi5HnU3+JjX/HBqH/8h+MuaA/Oh
1N2pbL0hXTTNoHsPJYwC/NginpREBDPPg+IIKJksjRiXHAFAbFMTmXkLbIVj
J0734CxdYScZSb5lvXuaAikFsswOYzQ9OlSQLKS/lnKMq3kgyPIz1NcSvjQI
VdswEGcO0MY1JuaC5Wk5Ji9anzXOyWB/A+IunW8eiN7W6DfJ1kFHaTk9i9kk
s/uyrh0jryLxORbu30MzVs666KgdO+PC99HIKAc5cDN3v7smGSRYc3fOyH6R
gEy8ziriWaEyAemwbT6ny18M/atZ2B7s787misXUbILCf9Xptgw59FciaZYe
+nvZTxgTElhN8XQUuhPJX1H/YrCeFlDt6JtavpmaoHhQK/EPF2yBuSrMX+5B
f1WD/eKatIOJ4rX+iRGDplSa5tWKSVwJhUtBNALX29pdTYobhBlmL3MKqPmU
nlWEc2d/qZAlnVecNNPRw5ME3jecEdtBaP4qxHHhKUvU6+8WNL2AegMOmY87
KtOF15946JolbDpJdxTyYDpg1TFkDbGrk1OgmaV9kqE4FN1ZlxoKD7Jpnr75
hdD0ddOPfT6WcANvrLIkDxvtj0WPQSA4t3zRTuaaHTZdMBl8G/zpXJjfRdRH
IYD3IKPIdIm/UjtbDOySqZhPqIRoTrfnKanLq5wCl3GiaYiIaQbhnisSyoKR
8iHbXIcj1zrVSE2nc8nalbumak2x98F2rHMt6jXH0lHuE5CGuVxm8T3NY3dQ
ysS3oEwtwHVEWdia0pCwWVQ/kepPO7j6ACKgZ2iK+FNyaybPGbP6C8hzhtpV
3FjsOs4mSunEZV/DmCihB7TbFU0cQbHAQHu9YU9Hlrq+uBIZ5zd/XZ5mZrMG
OXJy/XPgOLFQQuOyKgybK4QVL1N6pQkLAOuQC34LrFgpARk+sA647if/tAs8
+271GMk2m8J8dj01kWSFEQDpbGjiinumExwoDkWsG7mnpwJfH6vD1jHa/Eth
CpH1fA8X0qTct9Uzvh7pC5crn4d/L+DHG1eVxR3CNns7fph6ngnw1VQiNxi3
HjM8tYpQIWb74xKbKVzkbOoFiaGRH8WkwkILBp7BA4IW0N/SaDjFl0WH7+L8
2n9/U95IO0CI/ate/NmE3XFqzKuD8TOn+UZKdCeMN+hO0rfNXBWdjTfds742
nnVNaa4wE2sg8TZAwnx5W4E+iXFdtKHRNcqIgVyRq6uzJMcXdluFplC/LUVr
rxfLgugDGeYXhCRKe69dQDqysfJlPJo67FXL8HGqYORHXJEpO/vmmwtf6ZE/
En8rTtbK+FrIxWokbPOSffoXJRYDHMXJrmqZvFLVIWVhkNRHw2NRaksfXgZL
oTZzmyNtHxltYbJptColbuXq2t09dppaWCDTNCzYb+eh0MONiVXHHpwdgS/q
g7cviUKRRXqXtxhvge1Hi/IJ0trrvoQ88U14lQNrPsidF9kDfUGlzlHKBBve
X6ptqkeeNr9xmCEU82HJ9sle85jPBPIqwzKbVfCwC4cSmISNY/1mPnoqUcAE
W6/bxKw8FMfI674Tr5G3ugvkrsV+6raMEVILHu9yJzYOWNYpk6tCik6suRb9
XsyZLRSDxDXxOifs2uSI77G6wW9qfMvlbp9hW7ZRg/uP/fvEJeAZzRr7RQLn
dlE3K0mr3D9d9MZpFZqvuYD3R0A/btcdJOz/LKvm8tPLiAwlbOpHR3ozgnXt
JWHZmDY00g9+LnQe/bnDxpr7ujqX/v347tMQ6br9g1smtuKejVSh715j5zGN
063uiYPQ4I9wSvgAXoThXzBfcE+Z7yxkTrrRVpqDNV1mJpYg3SmcVRM/h0XA
uTZyAhQvO6u96r64AA5hTM3nCIByYYccFJHaGag1FyNYAdEoeYtmscnhKXPJ
YJnbGunCuDPawYHqaFachuUkEp7SiaWfH+evTmlHQDDJwIT9u8gETNtlMv8h
Vu0ZCj1CLygthonMzC9sfaXBlAahKC+6Qjt5e7DuyLcjMltwAyGPotDQGRWS
JfvQkGjUlTwasFzA49iuphctH6uaBo5iuHIFKK7p6QzafbaXcQYLFk5KqNz9
tVoer0bRHpEF780jX8rm63vLGBS1PXTORhdVtGYpTgvEivdMI1osIuzd1ZBE
QZfuyeUHxUn8O7YyTrMCzYyfxJVVfqK/5NBktbviYFJbBjTwEATskIscWlnM
0X6J9BAqGOtBt+WdO5jLgwGlLB2iKbmGUpesr2pvP9vqD8RnaeC+W8N8rXfd
ZPGG0tiO17VHaNEJdRtDT+406DlSGtr545r4J0GEacEw4T81RhLqBMGFEvLT
6xdZyb5mxUUT2kponMmcYD/Vja1wnr5Di6/3DssM8yDU23/vvbh5OG5sq4h+
mRfbF7xVqJQT7uzcOKcHf4NW1iCdHu9SqYr1NSnYqWobnyDe3/gFd1kDPLcc
Ggetz76tMU4OPiMzUCYfxm/NPmo3qx5mJ/Ar7Hp7gUm+k3lsYnHuJteq+r+2
EfpBnVundkQbGv0pw9OalKk7ISFCiOCWDZVIK75GvensJJ2cDs051kKmGctK
IJcgH4iSRRe9RzLe3XHJ3sSf/JO9BCwS2g94NHqOqxRnyj/QT4zEA3f/qi5i
ux576G6nHY2W+yTSjphNtOTrqv073Qa4dceV6dDT8SOM2Sf95GjZOuszpUVV
VeFaqqw5nrZ+YlGHLFggfjA9gQdFRDLHPZux90Ps9sLZiP2KjsH04M46Egil
Vhud1MjTdNHf3e4qNRjDve6ECj/Lo2rdxML2V84Bh6z4F+cxWRFUuxJvfdhS
uThkK2DqtONkPahQ9GEhbxXC0KztX03RN6IPCJJNlbiY+wG8YUhK6TeYrtrF
vNObeOF7RzyF8pmP62dLuhuzo1+pEX8ujs13ZYaJfGuk1vkarxxEzs0x5C2f
r2X9mbvqc2P46fjhRLRlKH9FPqChVoaQdQ5J7KWHrNTrNaARjVP+OhEKZmB6
tD3QR4tkhWOVHWjHpI/c+wrJ3R255aKk+1h/OLwKnD8aECut6elH2w3fJV8s
evYg6H0szgLCbDwFifRIxDXv5rF53GhrsWaEeyndB0h8hQ4rhZUUhjN+PiBy
TyGmqXtWBPs7Y5AinHhRR4V3Me5Uccnl3erZxQ7Bfttwwxc4bz3OYnq3U1H3
Sh22m/+DMa+dzhfSrL7TjrejQTEoEyVPVQIIjAag4IU0rzGkJGUuDdH9AjDH
RT4WpXwxKsZvv6apEi57lEQyxgwIZc4lwe/Sz5Hm4K/872sEMl9IRKGbLxSQ
csr5dRgaDzmQ9O6zGxvNCAPwbTwmgxhi6t95Rw2CPqN+izDKj93iJMw8ISfV
YixghDfw0dg5vc7493xYt+R59OxpY/OLnZKzmEORedO/FdOR7Bw2/VpZ0evt
9+5wMGRq2DkDDbR6mpv/kvYWFAIo4U+QWVHgTxf67JDBmQw72Y4+SBH406CY
3fYjtfRF8JcWhJ8TJdWXvKHHagHsT0FrfKMD1wbbzYtGlhUAFRKHGuMIl+Cw
DCmvVwCbNFfcgD5+fxKCEpIYd32cM0dbz09WUedigb77jAaPjfBrnFlhcJJ3
UWEb/VaPq5vS6BMIYM1zXGcPwwxf44KOabGYSKtjPCge7mfLBgzAbg+jAQv8
1i1v39IV0UFNE2Z70TURrqXtuDaPlTUwrpFcM6pVezY+HiNWtaFGCzKQKHUR
dIa36ASfL7v8ACIYM8HwY9je0dk2e53X/5JXucxwD147BQQ5WeHD3AC1v7wM
SeLSd6zD4u2rBFrZR/gloHdueniBUJ4IpcAHhDHK4EydtNuMx27/3HgMtqE3
J2R+BCyNImGwNXemG0H/hoARYNtRT+OlT4xQ94zhGEan+r5cAuQuKJeeyM/s
rYtyd35APebMqmlJge424L/Cdi+svxbuJ7AEYHazMXJgboo6oGSvsYaHlPjN
rasJCQHhqrfYeOCmEr/mgZKj4nnwARp1zn3iOa/L9fVJ6YjR7KAegWab7Xu+
MhgGaZg4jP4ttPe8oSe3V4x7WiHzVM1e/9AX78L39K3mvCcMyIYcHQhmLDo+
XpVKWkpTfjFt1QEapdKKZz/LG/F2Kjs++VxvpgbD7zJh3eZEf4191sWUKt/z
MIJ0KoUcQ5c8lNktfRA/iZT1Gd/i3duEOn6rYEd/ULjUMnM1VY6sUJo5jBIM
nM9ucGW4QDPdrbJUe1sneTW3PzWzInuHoGwPk69+Q3rNP51KBJFL+5KnWJGC
TGx68OyBkhQlY4ONK2OnhIdxCH/ixFtaHq7ukw425ehyor/QQLwsFM/SxLRY
Tt5A7dgxYn8wpBKvlqVQuwpVoSZ19iOkzG0X1RN75zHjg5Czko/ICSrteMhv
5dS+c3nUadf45GoS9Pd2z9T1um9ciyPPHbcfM4xAydFTL2BLdnj/3OxlWRZu
35/hMxuwTXFR4qJ4vxxD3G2afTGutEmQ+FK46DmZ14iuOAHfWYF+EnsFQQuh
TaWt4U+tJcaxjqCFTqOhnGR7aSqt260G0j0zAcs+XdDN1nunSeebU2Fjyp0f
Z4xxEcY88IkAqdRHq7YrkkoQ77I0cFUZXZEbEDwwUMjb8H1Qo72WexoQ+Ruj
JTNKc/6AdAh+rF3E7MOmXHweVityP/tlsZJaZBNG0J6hmJYYqWsb5QYzj5wj
6F/kelaQW+yFtgRzcIFcGsQs3Qp1TPDwdVHMJJ1xqpWmilR/O2ls5cdstMxd
JJokk4Hiyzi3TsNAOMWiTFYOLgTFlIeNOc8/+5HQIDtSgd9AaA/mATL12RSH
5KdjscuMftE5+zpAAhljzGDO4rbCazkD+MNWLlEhsuSBhWnKP89L/+tigUog
6twFJUT4PbOKl1onrOrj8QSo9D9QwOEh1JrVsyteEG61ohZuXxf5JK/Kfvfz
Ot70En0vpUM/LwnxCVw8K3FuKSh3Y+TtmUMlx4QZFFVLF5uiugtS4XJRHhqC
Z0BYOB/nY/myWEWOF+VOJoHt6L2LYaELp8E/+LsAnXy788mkSdxdDDpoyThk
J0swjYouJYvazAW7y7AGIEt4MCNCE+eXGVo1Imu5lmYR67leU8z/+diWZw60
laTAJ2wR87VIMamGA7IicwDXMTLiWjfZgSiWXvVy+ac87m1yiLbFhtmgchJv
aJ5JofB+tiORI96F3Ci7+0sD//eGa+hYZxZ/QdfuxSlvlykp+H8cEoJLe3Na
scWOwj/x2kbM/HmWD9w9rbNW2LkvkI9ZgPEHtQ7AhsbzEXKtAKAzXtF5Actj
9JX1A9nLJvVh63cuEJHsPBHnl56SBw6bJB5hb8MeqEg1bKjFEzvMQ/JfTw9o
Az0E/MJ4cMSonHZE3+xmL5/XBGjmtIU0NSMazwOaah0w1fwocs0BiJunE1x+
VMwR0He4xxMKW9DqHKqn1FruOBerVtZjVLc9ASveO8iBCoBfnQRnpunEnTtC
KrRB8+kyxG0vzYprNfZtm9EP3briq1eoKIEqYGQ0JYmRTrbUXOF4zq8ZHXLe
vUkVkOs83Salg6AcfqvC7eBRG5gLfNFfTruiKy20HE8U1dCyvqS0HBdCARyO
TzOkBuojZBGHlpEVSoztQyINQOFGL4+joGK2u/Vof2G770803PUx8aUy0oRp
vGYJWP5KOxu/FbRWEfSd/xa46YeeAOji3ClSd6Vk2kqUUiykswB1X3y+ZkmA
hvVe+nCIrcrbcM5jajD3WvIKQAYcW72TLOBPRInRel4ajRNkjOIsEVDXMSMn
MRoJ6aO9gVieKD+ACA+Hbbd+55tbKtsQij/pCNjg5/bo853LtqZq6c0pVS5M
6af98Gt+5R9ExUlglnqT7G8qa1QqB7GG3bAf9ARjhoz0vWp5BJasFXoUL2ds
x7rlSwFu2nBTFuHob81VkyohuQa8xEW41OfDH201q/vrw86uzL494qHWKo+f
92MKaYV/ntp+AvjbB7ZDehw/25tNv48C7v2mhe1qsxC7UiNuG8AbE28WCrJg
7ivdH6sjbioDu9g2+VRNvQUxBRHOpJsXo4YHbLmVQJHfJmY5o36Z3cHWfOJI
G4/byKmG7kYwGmr/5/Fq0o1dcUrtpw4VbAgQl9+5E0hSozOl3O4cMfeOXRXw
1emN0dUouXeoOKJEQBzYhlhHvs2twYEJ7hcyVMCI/E1866l/ybHZyCsdtZ32
W2ijha4bCUu3oVnCw59K3Z7PXZzxk5Zle8O4e7LrGhJpTZdA6W9APTUXUFNd
9ADtjRo1cbWeZ/IBaiNb4JaBi3d8V2Gf+FIG07kQ/RyXJE63CGSBM2YNEVPl
I4O++ebASJvsT4kCrlEI2ELoo4lvIjcWhFkIJpKHGpa6SMal/rL3W3jvaIth
1mxO8UAR4HOPLu+MJ7fHVXpVkUkBn++gDQrE0uDr6Yy9ovUyD1Fe3bZaY+cr
TZ+/zPCN1d4AMNr+n7ljnViXOVLqMK5ah5NtqfTrM+7wLQen5XHpfgXYaY0m
G4czKgE8VUFJ4bhqnbXbJI4xfxtfNKsFl3/EyHk2yySuh4uM+K7EoT0UfGwM
A/j0IEkXAzU/svINQ8deQ+t0EXoi587GINLABMqFJoIPqCbmfuwg78K92M02
IxaHH22Oe63uPsINEvi2/0m5Ct/l77JdTUY3rkFxbS1cBJADW6hjJIL4RVOy
3mTaG6yhYm8Otu2G1yPH4clN5wyhan4K7333Mbxzjjfrj6pvrw9e6yi7jCyQ
C/TpazRlZRDWwWT2JrKUwInTU33BlolWMsC91fhsMRzSCcuUd3kALDLdpYX5
IuKpQtJ9cLP8j8sdflM/dSodfyUfChAUjlMePysKvYSFsjuEiN80D516fwqM
c06n7l6bqteQ+HMAb+EQHnCCvO+kSo4rbPnq99D3dpYVRY0NcljkYnwbucEi
iF0kY4/NIoFs4Q33vx8TA0Ee/Rkz6Y6/IfvCet7LhBdkf15AVbq89LQylQXI
jKvPp3jwPAX08RxFSmQ0ArMUExQlwXnn60uafwHWqF2TFJn95WcQ+MdE+yMJ
UPtPJeC4OZa2G8UPCu4zwQfwvuFpZRk1gKAhUcKcvQsTQHci4xqnAPr9II6G
ETrOkQtNuImFOCIWKC43dvBMa5w5anfMnG5Rmq4z0ZMpWKEiPJNNlrWHe9uM
XtAUzJMGSC9/Sk1+e0OO34FpbstOw+JY1J+eDNYl3Aw/RbiPXYawOUP7t5Bn
HVam2NaGyaFaKiV19Nk6kYSM/kvtzAbMev+q4Fq6LpU8jYjx+tb8f/DF/nb4
ic/MRiOeDbcW5Y7bJzxRRuowjJb2HhcczKZJDKQ7gJnnZi2LYAsGgerjYYOo
tal7XaCxVYsuVqHDfzITsyRayYfoLvTwJX0W59ROtDNsvTb4sAW1AX4KQyR+
u2LapyT+k+6MSRrkrCtL0siLIZWpaZHiRJXaiDm/2onXD5LE81aG9YzDmm6e
ZdnC6vhQroXN5gAC6PhmMc8zI+TTBHgFj+/5quI7Q2B5/rQw8gMQYITB4TDy
m7tgF/NLe+PGg9Eml3/jtV1ZZJBYXMchz7AMwqnryGas0WiqEAfchCeWZ5uy
ZHpzgSCOX1TRJo2isCdBrGRbeyl/ZidPZ+WgPzyhAxtsv+ejc09+TA/OOai8
cSJcGWKPc/Sctebv8iB9UUKgBDtJAkhO/GWt4rmvw+zvEvLNRQ395yHL9NZL
sr/FkWCwA0p9ydvDedvY83TgxmfUOJGNTAXIEtkj9XaZdJBOlkV0sGwJICN7
kQ3Zd4UMEcFGDNIqxT3sWXdABp9FmOHqUVgvAtmJr98AJsX7rbi8tFNAGlgk
7Ic36Qp/vZj/0B7ydpdpPrCfBZ79N1Ao/LHC8aeQ+/1Xar1CQ1hQ8NHZmJJO
TXyCLAsF6/oT48WcpTgqfi1gRDYexkb69oPJRF8t/SwE7WPFR3S8wAj1tH7N
5cHLdiGvui+EBETwaKYr5regbV77UYdGbmtbKc3O/HJSC+kG5rVEN+sJ3Y6r
Voa8MbwfsdeFqjyrS1eeix3JU1Iy9N81pwDbPhBokwBLytxQEc9UHUIVqRoH
E9xu5431BAevr8CJ6+VTW9vnswupbkgNnVGBsNNAtPFlgNza/OSpnQflXPTS
RIq24Y1kFaR6v8rxfrq+pAQXVgn+tm2RLucfonpcc9SYvPfUafjBxYAfIyvu
BXee45XUy8sk1GR+D/Csm3LbdeHr1HU7s+pCHNIg/ldjI3CDTFclDVOYiKXC
IBdbwo2IHnjBTUAk21UQ+FwUE2LEFpBcRXr4naoE1a7bQT7DtgvDAJTLZRwp
52IhMsfDCCgUveEmc3hP8KvBuHur8XqDxF56BO4s1NDmklOB8LvmVNfXt3j0
GJix0A4cp5gJbA4YQH+fZxVL8jk3T6QQdUd/HixHFGIQz9kGOETXk8giIi/X
NyUQ2uLQ8LVnskbPhvXooCkEQI/G10KNuY7V5c/fFG2Bmg/u0N5ePtabENZo
lRClhd/tEqOSNNurgUcdIDiSSQnFAInx2CKTOkIQC6o0rDPdRm6mXNo7MDIs
yt372CjGkOAzUv65dsOtPHZ/haQXBTPQ9RiYcTlbbh0SGQffEk6dBUEsHWgY
MrBGlP0spXFkPHYjIkvR9KPAoILdBftzHUmwL0AXP35RuBW8X0zoPtM2Nssp
vBomqV76qDhscIYt3cOoAf7oBOtCOlxIqgzLdSaiRwb9oofuxYH3Jwc51YOK
hNG3pJAYU7HhxljhBbmIwBSHvVuYskf0+Ul5+jq/PHc+Cc2RHqN2TLRvOcuO
nx94DMbo+nA53P1g4xMEj5pHgzbQVOdGEEJVXaS4a0J5TG2ewjR9iXUJuw2R
Q7PyYIHFxxS3IZkmOBuA3OVBsRfr869PZv0QPrCdpgyi5bBJnXN8s4ygkhWt
N3j7PE8lL0P4a99SzMUea10mx8ooT73NjtVynKMXHCWOfh0mRxyE3MRpR5fr
iCiUhmyS+/wODzmP3D08OMSFKO5uc2fxR0T6JxY9TSPv3/WEBPtOp9YH3tQn
efJ1eGBJqoxQN2zgIaA5frapRJIgsSbnF6OuWP/qdmcdNlcmSXRP041qm2+e
y/0ikeTuZjuocOo+7FqPaZTugx9ohw0d2vWhqN5EqUmnTQwmp9e0q4Wfdawo
I9nTaeuwlkwoXmv6XZmRdOhElvwXiWHSvRoIibPhCd3ZfoTvL7CaRxxv+N+l
cRpkT+HPIs61d4iJCdQ7OpFnbMG61zGZHULUeBhBOE5DuxeeeejTy5cRMNkp
+azUEZr/Tuw/PAuRYZunMXZODQF3IahDFbok10JmpZ2cy/hZemZ8rr8rLo0+
tE6yv2x1uah8fXpOhYJ/cWc7XtvFbnDsCqli0NkxlleouyjsqiwD3v0a9wF2
Wh7fQua3HmEfFtYJNgYzbZlWVIPFXtdRTwdqtdO1JB3zMUPf+XdWyA0UVq7f
duKinsPpdk7ItoRylmrP4RTvPep09MFNqIRhRwAAL5fthibpkHRXY9ysTvu0
tkcoYVzI9jzkfGF9xp1gHGm/VpfnDwecYkS+7V5bE4z9Q/pxmabeOcPK1QoN
ox8eD7cs6uipKsuZ7WvaZAE8v2zaMvkrN13CqgHkt3VUdYgZAtZe49zUGNPP
xrK3/svjqn18RSMiY1fAhRbPeQH7hwjYGXl1jSTjuOqEcHSdozdeYnGvgbmE
pEjuaDH0QD7n7lAwXSTe3CNkBIdJYte/WHrWR05f4Hp2lPrJS2uFcWkxwgKT
uyM+V+CWTDozMBdKQCWmfyBYBfSjnRJk2Hngu8V3Tzd0yovjVL4eANROC9JD
IXDmvQkQAKCGd+erO6BEovj8NV3l9ttI+W5m+Lb7Kie+xkdtAVIqUtUT8RFD
JHzuBL4Y5LW6iDgaUsDLwfH0hgbsZ1Q0Lr9cQ+JM6Yc37n2OCkzPhYJJU98M
VzfS7xT5R7E7yneSqXAx3XoXQVvEIqdebf6H7uOFapctdT2iGVfOSFcOyi82
riojEqFFAmHptMNiZb6dx3PpJaGc3+NHq0//T+8E2EKPbPHE/U/GrlVl+D8K
prA7xESiS1UKyPW4kOaDu889iLbOaxHkvWYB/xqd3zz/NySSegLa+0y03FaK
vOyRPW6EZlvGtwl9amrj7Gyw0ZoaiiTPWqNT1Y24c2HeVGh90MqJTFzBqho3
xEhmdsyWNGdflExnaFB16550r5F8YqazquJxSHl03DCNih0v9ZDQDZ7489+0
0RBrNxuu/ieHFUq429uc6QeXxkBzs4ql6j9ZD7G5IrtjrIP2pzzF3BlOez5F
2jFVd2TU8ohW2fsp4CZJZB4JqMFzi/RPk8eNNyGYNUOqAZ8f+VZBjgfYr/OU
NE18L0dvySxuHB+TMJl2IzUnSpyejrYdj0QmvAT/H8yKQyf28R/MnZlAfm3C
PZYAj/3wCUxyefnn8KrL0h44CNhH/FBziXHjm+LKIaCWrYfV1mRSMTL7K/K1
9WgpDOOwnc3+1CO91caD8tY7+xBaXaHB/O9i7U9oELI5OMnnQ4ahmsocLraA
Wv3JtFdb3njX2jUDE1HBNWAbuy82AJJkpMlRSN55oY9HIKeuvfrRv0/snWKM
nvFzt7XUiq0K2B/KboE76sOTv449TSWdvHhWEcCDiCghI7XkI6QzZtMngaS3
lx4TusQE8NH9xIXVD6cywyp/DsY8ktKl9NSbb5oxkDH9FyhMIOjwGOqYdN3r
cd2uIuhjnd0R02zA0gfc9v/piVTTUYR0ep9J1VsBskpf7uVLThFOO1+evtgX
MJ1jSzU66KLR/hQ85qdPnuPCB01KjHaJVWM29642fqcXfWkC403Q8UgPKlFw
K/mt8zZGUDWyvvP0NvG185TjtzoSdArv27PFde5hhfFHTvnwOc2T+26vvW9a
XKwdxtT0bb/RiBTgDkmc8qcb8Ch+j2COFoq7v7sIy0oEwQW1rxE48yavREFg
19S5kkNe0Xdj2bMtcdSyKETnk/8wzzfs+6XLNeE3qXH7MvAyJjklyGG01IWN
r1yj4I8jqW1pUWAbHM/kcsUaT9uC3Vzj27E9ZRFyu79j/ciTsDWp5+C6O7xp
PR6SVjFczw/NLmJRL62y27TF3V/Gqibn90xMuuWNEnEYZCmP5emabR4shi+7
mI+t3CvVz9QbmCjG2NhiaCrtYRiNDxRUFtI42PFJWD8Z3PUPlYOfvNsPN6hH
kZtGm0O6gvt9w+MdNSfcIDFNCjQn22HBsmgEpX+8LeTvM8slyG6nawkmgTmn
HUVHM6gULZ9YLHxvEiX9akm2Tj8TuNaGCH+GAekmKR+3HHfbkVwmQWyItuET
+32jwU4QY/Q6u3tRgnvbGg4Hk5Inx5TvF4XtxxXZ8i8xo6I6+1rsp0lArZnj
CCmMs8XszjIz7HMSWd7dlNObkFKJy+KU8x3RwvHmw4p4KPTjIZ/n19etKH2A
3QJJkSWyJ2hVqVtEUoYuNCTCL7dXgB+Wi1C0Ea/8r+gbcmaLUt4POyfxnym3
GzcGwX4eAdTXXb4eAYFtbwipbQ475B4gge7S9RduADPnWsJClPfdRD4wvNtR
DgfmYwPcjhGEjypcfYfo+imS+kZZ0lwDvoQiQ9j+9SIVma7WQ2dbiQ7+kwow
zARd2Qrc9bxvap9VsEMMSbu7znV60Hz7xbfJQVur9jjprL7D4gokexiGE1lJ
jCmiQtLwLWtag6sl/Nsp9vSf5FXcNx8JDtay47W8UYiEr/cmvGqRKFWj55Al
/iCOF9JiXjU6EGSqkLNxu5B0m7jryoWZ1bPcTjxfsgaDozJEoK9PuqhGvsNN
C+cSmU1/fn8qC2EHj5QuKAmRuu13txuTbPGPFuRkUwx8HZ9rUQHG9WsSixRb
iyzws1yr9ibobL4tVGH4BMpVsQzPyq0hhXFBULRZxf1EXDqVuEZjuvUFyMLj
7mB7QmFPeTG2TPKPl72l+7NHcsARSgFLLw3CnIgdZwhqpFK8W9wfiRy06JFG
UL4Ce+/LGSRQQuyh97kHyiiVSNrMRq4J1F5//Zby+N6HBTsGOCVK78bxvELp
SegZxVY+1lXUq3FfkYvKTKaqSxl9VxwLcllwmcqZVSVboCr3W+ybIS5H3ziv
/DgRTkySIb2xCknwsI5NcC9Owa11O843uh1yMr1mpG36TIBfU8p6T3PpEb/M
iK/WSVX9SVmjTBYrAwJSb0aiDVegbKqObUhH34XiKNPyDgAa5eAnJKx/LCaZ
CbK1eEisthqu9MqNM/7R0w4QADm5zoxLFprgExOWKA/H23K/pMQ1FCu4oInf
8YNizuQlyVRw1xQGE0d6ITvc1ra2+oibEmNeT+9zOQ4QYkXEGzEyB0LOUyHD
xCr7Wb9e7QUBg+BtAEhuWLpQfrAWmzgbxbW3TkyCksnoztwCr66MZVYGCQFQ
PeuQUQ3mq8lh690csKq9rjkF0e8nRNSTI3aFK4YeZvFBSOCjb2x+A3JJj3li
ZP+79n0zwu63/RVdbMKtY1zhzKgSDxZlcvrmMNJHLi/SplE6s4Hdyppcy8cc
2X10poj6MN0pkbhGjIZOf1ysfExEzfvmD1Vmg3s8hC6M1XKJykDcJI0+HNVW
XFI5AJxo0/XOjCOunU+vNuxBbcCC9WNmQXgwC1S9jsmm/L+QQczmjeoF5kWw
1LVLYeUmtZirzVeO7TdB0nOtJkGk2bDX50WuUJD0X/G3Kz6eAUUuMWuLvsMg
tgiaqWV8k3MgRJkDZvLi+Nk2ph8xq2SxfBOUTBBd0Fdm0PsMHmsVXR2rAGJl
oH9cIeUfrPl9jHKdztakzc8ZkJRSyOto1uvY+YmM0EFM3r7ZPgUVA1CNIVxo
vnSh2i2BHO3cqhLk1HAJrnx+It448QDbxxqGUqebh3Cnh0pMfpliH71sp0+z
/QyVNxMTYx01Xrqwg9psq8lfGuVqI/hRls5A1hiIWk2Q+5rDQPOs0DzrAvsL
hBuJkOryGvhjeZqs/K8Po/8PGImwb//1DFJdUB5lRaMGao29moPchQ9iSJy0
iM8sEl3U7XtY5g3rbAl/CKpJQPtFo5XFB/3eJjiwjYZxkN34ZmGFZaXE36wC
wenKDdcd/pMqJZq796VLznh0rBgt+zxd3YQKUwJqTJpXE07f6P9CzLKikVLl
fCUNXl5zpEnZHZHuSQRAd8xESVPXf2O81wjHIkiziebqJW2mmHOkfQK6L3ss
o1bfsG6hqRPAZWfY/hE1XhUuPUZWLlUDr7hvRPVl48TCVf32M02xdgwc1MK1
T3X//ddML79LO208J50yNzAAfDQ4ke+Y+WbM8GtEtSgFb6ffvEbigvue7/bm
vdhbHcS77HhLp7WEbHpLHIAMSiS2GRj49KavLPwvt4EKbFUmUDiKEPhUjsJ2
OZMxOFmDqCsETTacuAY6cxU8L9Un3VcB8SbSlDtWoP9Zxj/FG3hZd4O4Y/Yo
dDWBq3Bb/BpCP5mKVdTCuZgxShqfr4zOuFwp8AQZQF9mSnKz4UgLCzMDnFUN
tumz0qsdgUeWQVEANidiIE5cxGYcjO21+NvPsN7xWafr5Iz8u3wgiaDDsSPU
zZ9/jh4hjhMa5829MGj8DYMd/xXjcPasPDT5Q5WSW1ppXENxuUYltykT1hG8
F6951RgB9nhz8tjGOOJCGd2mWEES6ZdqaeS7vYm2e8cdg35CV5K+GPh/uW20
AAbRzcP0CVm6acGUC23bYKDNliebQNCBmqvakAX+a5ZWY4WO8EyJrd9MEX/D
PKcQeCAnNNFVdqiFjDm57GrkpjXUKJir5CcKt2WRkG3HlWtJVcdGbAlaEg4v
lXJD4q40xA8bduVypTNgyhNjx3h1mTBSLnO9zQz6qcMrE3JxyOxf3n7Hp5g7
slsH6luWN8p6eEayz4o7mu+VZ4LkyMJsJlfl8nG5+7CUwKir8+lBIokCBBCo
uY9ldpyYdbnIwwisTqCvTUw9w+zgjWNyfl+4vEV3msIPRb1d3vXZaSAkwB54
EdvivbjTbsVAoKj3y/mkbP6+n8enlr6NUVK5aySRfdb6hmCvlbmz6l2qWDtv
mfme2BPaLCrpSl1qR/hGnHx5iJydBAQe9MgoUnUpeoj+8FXI0WbngcHb827s
w9uCPLVxvFP8cmUGZjJLylUP3i86cN476VHXeeu1emqgP2EiXATSCbk0dJLf
RNw+EFlxpLyEk2hLErOeODVYWoV5EqlEeyBAzHBRZzQRDwPM187gzC6iUTLo
F7qtSqkx5qMYUmJzSlywOjBhjFOoPQF4VzU9oV8/Ij3/C8ZCucR4U8Eivnq2
ORNYA/WWz+4gW5NZgNKaoiKyVGYLQwpNp0yjrjOhGwySHjaCRkIDZhtGCh2f
Nk+t75J4oAFeQJM0GtOVRmqqsoTWyAZvDb+64iIN9rEFU7c/WhHpxvhAI3xF
mYbstWagoowKNObRZdd0H0dY32N5/8fb26XQ2YEUe2s30TtgLnzIRtU+72//
SEWd2YDqYvGA20w5eZiQSoYc6mKBn5RuyjTzCnCKmPHggTdgAzzWmsqk4zCC
Mt7Sx5GSo0zConGPWOxBsm/og/0VQDIoc+6i5gYdEQYHw1O+20ODl53QxbdE
FrIBWJOyTHjj7HDt3LMRlcxm6LdrOSsMaHtY8oPaiLrE/LhEdTNzgYFXlaZV
Q2ZexLvMq23IJMDgnNT4awXCA5ECusFUZ3YOGGCQ8M2Kx6hSRUyYDH8/fKlH
0nuuQv7sePXVpY14XSuVku7GhXIGc7LjRMrY7uLm6XVQzAmnMg9C+LKrCVsk
p6nSF42hQkhofTRYavGoa9GzBLeNUKTP0m+GqJsF29nAoDw2Zq6GczknmsO8
18qXmhWx4SoYUQwohKCjfJtRCpnt2JCAQ3GXWBHusX9tYyjV5cTHm7LgrPAw
IFZ8r2HNaukrRxBNaSLvwGaPX2aZrDWa4eJbrzFycf7Uu3esJYpsySeogHVH
fGFO9v7RCKjyBlq+OLB3aBw5/GJ49fil32qbeUSoPEMvPcVlTfTW5JA81SAG
+8u05SMhBrndyAa3bJUyqmHDdt6EjjjjrPKgkTyrdNxNXEdU/yJyejmBxGRR
m5vNxzr4tseOTsPZ4NrauSN608av4Baq1tLBlHjlPGuabfiw2HBiAMVVZwHj
BsAInCJaIKV8M1vDgeJsYLbKyKANd6uzt2cno5Kp9zS3m9N2TU7NBxLLNk3D
/fJRJR+Uxd143Ifp+QkvSM81z2zePiBbffJF/00yEcgjOhRl/uoScz615xl4
jUkxPA1tkvqV9iFpyJJT3t/TQTCMcr/4eqJRDrXbPVV+1Dh4L9iacS+P5qeK
bQRVHrbmEYNsv78WYap25xP9rYP+omBVij7eTNUbQYQbveqp5V+ttqdQpfUh
5J2fpNESc0+ylQfijGxYqnHpe6MPs0fHTtrNGvWkXpJUKNPpBtUm62idd0Y/
taxm44ccfWv/xw/J+OYfc7e1nBgx3tKWvZ6DnQRtl0iugsw5Jw2S5k/qC1Eo
neGVa3Otg6BbHv5tHiro6x74qBLi6yTsLnfQcShumJksRNViOOJv6LFwFimR
90LBAyvN3kqgU7tBDLBdEhvdPsqLG/f5lTaqjdH9GlLfY5fA78lgudVOrcMA
IOJmcaJh5K8Fz9fcRhi7VN2rhYW+cx++QAt5eFjaL7J+d5XYXb1bBP/w++KE
IzWMtLSeFR0n20H2kJjTVp3vInJ19kLoGpatB48SjbZRGxh+BPJFVdsk4gmH
H3CHvx7C8dcuuuNou9yNxC3Pmhd90qjBdE2r8iMVVcVC4LrBIhSUssoWV7Qk
kDcyDXuCI9GqPFBbfqVIS08SXxf8BbhHc0G1nWeTkRtnR2v3qk27bJpppcJp
4c9xzHzbQtYG6BOGF5y5NHJVGFsCunFk8aWndMK+hzI/qXibl+DTPie4L7f8
yJLCMxDWOvmfC3jr57wBz+/Os1nC6Mx9u73G0fJAEZYF6sZpiDdxh50RpYgn
Ddp+vxBghZ2bPRk7teVkDDpUsUEFrwQ1PTInw6FMuZAdjrOrC927wN39GHAT
B9ataubpzaxLjV8DG+ZkOYsxUJlDRBz8mT2t2d/mFkTDS0wxVGqUBknW+MCn
54enY8okUWJFSIGX1921klDrY0HHldZYOvxHqxXWtHe93UzD3PqH9c1fKGoU
ZdLB+TjIaVlN+e31Z9iEmHSUKPo3ImhvwQikvz6qk7JdWJZx1vz2kE2b/IVQ
Yrvv1cCJcjc0hafQvavRb8HHDv5rROZaYWjf7sDhW/gTHq4MSHAAXp70HvAM
3dZlXFNYtTrTCYAZe+CVaiF+TDjzKtUIsX/2c9IPFYSEAPs3iqNJaP9Wu9h+
En0RgpQYQvhDEMSr1+k0kcAooRUC5vD4RM3cAzoI42FlgOonagBgdMRhRxrK
NhqqKxHp4Oum0HCKTfMKX58gGmTHoqtBtJeHFMj0ga1mhNnnqCr/mbYQ63hh
J+SRGjNloMDaVc/9TC+tjPWiPmOjPLF1g54wpptBUBzCxXF7i05hotwGuII0
n9XOmWdyT81Y/84NNZSd9Dmt/Rgn2WyLNqkL1FSLngPitByk5BHdsWJwsGTk
UvBlKE5bpuF5NHa7q7iWntBdW1Wyx77k38/uhBLrPmOii3wwZDFfbO4ayeAO
31xf9G318eGhNW0P8sMnE98l36PUvsrxlKsgxCPTTW/9yeBPEdJw/7td7wOC
C7PtqrTKH7AjN4RkGhkxehtsBljkKysj+JOqpxnBmd416eSUoP0YZiMwVRce
Wy9BFnE0OR6GBPs149PFekKT3egtnWgTvEw3RsSL2qlFWz6HduGas6AgrsXI
glOySb4JzYhzEe9mfBgn6AeI09dBcqub2SLiK3LD3EGIoyHvAImc9qVQqtbZ
hbgo7S6h7Sz1Nb3jkrooExmXXGOQs+7iIzZTFvuYLeV79OBOcu0EglcJqCOk
D0tevAtTVdyqPa2/PuGhBoDCWLQaCEoVeae6dtMwtHOmhTFcLvFsNU3bErtV
icT+j4ZLUPqulKUcrKKkzI71RgWTuB18gOJI64jH+i13cmKPgYO+VZ7G2Qvc
kXgjGtfQVkf5lXCsCzxj6z52PF9mYNG0NlqizdXiKww+74C3Q9+URVzMH2Tp
iel3u+CRLoUMT47dSVXwiA5nCYG1gm+1CRJopJKsGZa3X8e90EuNbnGNRGX5
1qWOKsrIC51l4V5pEz9/c52SEbLs2uLlJgVxJadrJBl5WQ0MR4WHRLPcwN3P
3Mp4wCgeMZs4CIGdSTn5596HeOTM5JuhOZh7c8wNDN/dq3oM303qnZLloIG5
6wwk1AoR/uAimcpriZ2pz6O/xd2F3YcBp4yo9exPi94Cs0M4HWgcUk3L7+No
t66wsIlL0IE1idADcUpfha64dhX2vrVLAqIO6qMgk82vAjGXlOjdIo79YABh
MfDo5jqhmexJ7iyt9eN33KGHiP6IegT9v4ojF4ssPCekuxjZZyiTe7A3CILG
IAoDEHKp4yMT9pyy5w4omqPcNbSpEQBCPRwgZ7Jkd5iwUnsDrL7+QLwVL+tF
nUGwMKhiPvrSeJNgCQbL8UHojLKuzr1Tf5ndzDiKcO6OzBirGmzsJ0MRfsIg
vVsQAcGiHqa9hr86DREu0LMysKNzGVT4OvcXn7s1jtuuZLkl+FYzYPvM+XS8
moKMRuk1c7tktRwou3fTZJrOEkNmfw56XhYKCzKfvimUUJ7ZxFAw4p3TeUwB
57MsExiHVBRDPHqRn5dWgUaFD0dVLL+iTGWZMqiL9oENo7zhydOJE5wmE7Jz
Ar9yjWhAw6UiKB9Du7JEfUCw7flOEj5eYBxxGRVWRsvWdFIURWOnnWTdGXKY
+ou6U3Uq59x0U+TeWcJxR8ubzJ7YTxpoNmoMiEMD7vWLxWSr08u9f6DB9GvZ
jiNEQpa7j9u8rj0K90MXRTJfu0YoLa/NX3fdWfcJda0dUelEZLZmFpbTIX4Y
xe6nyRY/rzL153wXJ6hRQ53p2xGel4Xv4fv9DXtuEotyC2LM0KfMR0GYDiUQ
o45+PNcDnSxLOhzd5r0TXy5/I1rUp8BtRNZJC6VnxxkGk7N5wU0AdoPK2ILT
+Bsx96uDn0QFqcOmteMoAX9cx2GhOa+sizvru/m6ASJgEZh6OOcl6mR501DN
nfaUkco7Uo1WLhpbijFphovBFjwSwKGZh+85QxxNJ2Zx9Zwctk1V7eQqFgYy
QvQdCOQBQ6x9Px123TKpkpkiUOqB91DdNv7s6OwrF5CIpkk9Lamr1WkGklH2
jOpa6E2wtQ6+6vjLjqaFnVVHL8PpsDP/YzbCTEJoy0jjbkcoTEEE4b2JbVNb
sx0DFRq+lMef4ajFFeaxmMCDxKJtQKXhE5rTJ/XZjFN504n2A4eJp9Lfg6CQ
28C58ihnog9IMb6FODdnzGZsFfMeRMpK6Xg90mVcTMNsSOh4H0NHYis50DTt
M1Rs3LAxdHHPSK29GmCAy9xeuOGUKK6ZIlmZe0VtLX74VI7xZjKJf+I30Ed0
QS6OzuIk77llo4+RC7LhscR9lzz70CSVnfw97QtfcTCqTuNv9GLG0Ij9R50T
pDNKXKov2p2HJzIBGFIvKdPpvksunGQUIy9gt50hA0+IZYX6QNVe7KsFuE+k
v4UkgpBcTsaV1jhXD67drVv7PrOkNX90mbSU0dSftz2dASnf5gmv1AvY4/h9
Tcb4wGyeVbO/O50lJJdFGxtXoNDnSP8YdLLgALlfL1J19c8LndsKwNuzENXj
DDM5SCQ1tnWkNWbzd8+k2cRs+07AXf3GY5RZVLzUobV3K5ABvrq0NuzlXn52
a3z79PFDLO3da49OjE/MS2GmloJaidWwatlBVwu30YtbzAC77BwUFvV+bAB/
G1q0IoGqMOYDSND7QqBJkSYDb+u6mL9KOljQgxaFmnhRHKcpQNVCCWRLyuXx
bT0HkCuDhHjYR1nlFYpL3gPNSplpe8VZFhEFYIzQ+Z2XLQKpvnJ5BkbNu3K2
DAFI+2uJYB9cl1P66PLCJesG5HJQHRTzjSie2O2VPtli3dLGB27Z6d8Qup/o
ifUejjB/BEptdYUU1+IjVdS2KPzycUoBpoOWVTp6+7aSNM07B2SkuTeC3EhY
Cd4/vbWnMl9G2wdIzzkPp5pJ/Xr7CXshMrp3BbTFSCV8FmXBUV453QQVdJXI
bEzGE4yZFGHiPyTRx+sVyVeFZgjTR3fBw0P0dOMoLXCbdWVGavYz4+8BCP1q
SMzofeH5cWFePnS5+iMvh73bjWRks5xC7OcqG/9XKd8zMYHkcIsbLC0xaXOU
hKirR6tNkV01C6ZXhHlnUYGWDsy39RcMG2K4+khvM6sbKfKevgY/QnHs6yd0
RljxbsZNPOG6PbbG7V/kXbmeQvRQmnCnhQcQuYeCySXYajL2oz1tFJ4zbLSk
tSUbQp6aVJVlKh5jiRo2eBlaLN4aLnb+dZkn7n6j4FmFw4Qrl3iXYhIosa1Y
iZjzsrJGqjpo6HoSy4DwPb7twXduK12saii3nOZ8hjqEDyhOW9w/DC1JwrCV
1zSOLsK9q5Ry8zyVbFRHXzBmmMnvy6QvdIxfoCPLCxyWbQbJlcn7igni6odA
TS/Jxo9qDIMHfuf+wjeuXNw67q4aEI7+HLSkcma6S9Z3PDS9Ho80i9Su5ruQ
cNWciTPDpOT5v6WW/cCybE8aEHXyTq7qXYtHwWEKS/3lPFxfetNiXYp+s8Il
bSTn6l4AiQtNj0pQmeA5DHipdljzlcDhNKDNAuwN2bWQRG45i5qIkz2xvLtD
RPaN6RbELSAQrkeFz1LGNscKyCd4p/tfCrLMwW2bK5PY4HjdGGZI5JpNybKA
Bt7I7Izc8HqRXg19YKw7Zcr4kmMgxHvqJzcMi33r00CIgQiZGuRKwlpMVLZM
3S/ZZvBItSnJ6pv2h34SKt4iShm7IBYKnuLUf4lCUaCUZnFY+f6piRdv+Jaz
gBS+kwn1L6y9BRRgRhcV92J6jXnf9QTC733EwZLmmrolIeOykmIgXS+SZtyW
Teg3AVITMHCS9QhCQQRf9cfiEewpjHvKVPti/WZ8MRbd4TZb+ekUczw3aSt1
IjNbh2TjwmOEFHzDsGoi9W1OtCmPHMBqdqQzI2ASmKEgAtQuVh2uI1Nbgwfk
DAZW+IBLT6JKnhF+a5t1MTjHEQncLkH7pq2Hh1X+hHAvirzlf93eIdyneVm0
uvzyQrovinCI+rADxFANTxex9T51SAGapQRrdlfaBACdy5l9A0Q5ari6tKfw
Uo94S9mrtqn6hvDg1vLJxzE5Gag7DI1vj+ooBq212X2xkjhbXkYD3q9ikqEQ
vnmUVv36RD75NDaW2fhgNbRBDR8hgDPtWBdMTlcv/FnYgH69lFkJeK7V5lCW
MlHI6zhBuhYgSNjKjtW4DGThntJO4ToViNx10oYXqABNE4nTGH57pwZP4l0e
ClKyASl5OM22jrRkTdOIKqoKTK1zA/cANG9eSd/Y9LK/gN+qjDJz+2iTQxvF
7eLcgfthor2hvq73i+WT5ZQo8XiMqFEx/F44F7xJTUs1IVf4g6Y33qHlh2YV
wNeTvDni9x5PLyeas10qlY/J+VZly0/D7+lG6TCzDEEtpV4VfAZZBHgjsHi4
+QRW14UzhEmPNQS/7bwsw87qPeIuSch8BIzzjdf9ZEPIkEad+76Npib+Q6PJ
+HjxUgxwXUZlbwqTqmGw8CuoFuMCLBLPwBjLf0AAs+ehv4C/kdXDV9d5t7p1
tsFIDY5sg0m5OUBF3PwJgI6QpWCUW1Fi3FCvqmimYSsv3Qc+MmneR9Opuqbg
Ch9qAgS8O+ZCM+lrCq4Gqn+vAkJjH8gdaMfJETOEGp3t5KE2Gn8GYhu+/F1L
dOXFd85WLf/x4nKheNvWeUnMbwBpbRRTEt7j2mEK83+sAZEj6w/qA2uXpjsM
tICC92UTXnAHSuDr79e3l8byS3eHSMUnnd6xJDh583TCbEw/AM4DLqgHfQnv
wihxfQDC1s49RylCDFDXsjTl1ghR0vnLC8x/CK+QsM2rFYeMGmg/26OhgW6J
EDnXX8mBKbgL1SxyRbmSDUgmkVtUg54IodwDpf6L4QKVyjqf0vW2+W5ZmDr9
P02tjavrN7oDu71uQQ5+ZOjeWCDJuexQSgNG7grAlaqWIiN+6siYBu/MyYJ0
wZj3VCUnzizYx61z9PrN/S9ZEwbLMlZRL3iMcQ7/8wCAP0Oup4FQe+maBh5o
PjsfEAXd6tjBFD6IO5NtWL+/PPN2tk3FgcOE+a1w8tEvbNiL/jPQsD4+TW9x
pWtkkLDWs12I6OZEFqHgRbKqjSUVgAnIUm50o15BhOKh7rxoqHCNtAEaYhd/
7LJGzKFjCJsWG36GE5B8EfYjbSbwSUkSki2zZtays/PxFjjZHDiEI6wPj/bP
Y/yJXEbQIEEkyIDj7uhvHlg1ZPQnHuGVCQ6fpetIi5AuViOKZn9T6d92UQVD
Z5ewVWMhHLF6czLIuf2x9ZwsAFLCBbi4jXHKLntycnddeUfll7PBc2tRODCp
vjiOraP9dUX44MlW9vR/wtnX1ndrVgjFBDONBvp5XUO9IZghYTPO8//nrj/u
6nfvpqm5cIT9kytZE+/KSG2X1FMyH3ZySzpkMaDheU2t4zwKzCrE8BysDcba
8R1JG5hc/tho17IDKZScTn2RPDe48QijMKzNiWdRUNR+SxNiUbNo/pJOqT7+
xnDrHuS3ruSC6I83zJu20qkXV7YEM9Qv6uD2VOmaZxnH7thoEMv02em8xXn4
WqDoa/Y3yPECcCJLdOK0O1WsOI5XYHClsZhTd53CX015txyMmR2qjybRjJE5
l91yGnnvToLoZLKN3xNpLSJK9ZgTPzVN5POE/CKNt02AM8dPSS2tgi3xGt7g
ghP1/c0krXG7vfh67S8IFT/oz1gjUC8HOv1DDQmyCEdK9GNSkfmnPuuuecoh
m+em82RtJjLZDDviqebFL1C+14naD8WJTFzNfwwJzHJRVIW3xH3y9pobveas
mgeQI11bplmDAL6Sbe/vwfmvtajxMJPdaNDXSgy5rbegKqqJTFzMA2Yg0uuN
ft3Tw1ZuXGa1fZpuJQ/VZjXsYdTVlI0W8PI/AKwm29UWEiASE59d3gfOQaq6
/LJkbjuZucGgVpVCOd+oxE9YJ9InOV8X3100L6J1iMC7IV7paziuf2AsWCYF
ADv730Qg3+1/1yNVrTHlj4VfbuhrRrCLnbtcyKCkKrJ5nxQZLUEEW+Bx0i26
e0nZpF+OvzstMXbgs9TBiA822HFJ8iT2+WmlNkIFH2LzcDwqwfzBGdcXh9gp
uFJFoiPUwBYxlEpBFpnEcGl8fMionV5A9qlG50pgVQvJ4aSf6TeUm6guVmEZ
57DYT2sX3fAZmPhpPp15RGU5kYu7GzR7Jp7kZg0hHBraKRVU0IhNasEbauW1
n+RV04FKkOzS2xP1dkdTtLUftixCuQK6gS/3qXVyz8ccMjnK7qFJbWDdBXhJ
NvM7d+gKx63MmoP967ye7wWxQInNOsuudlorMgwSLcMsad0pDsK0C8zcSlqf
RoC6Xdmh1j4xtBLbGO7KMayAImnMSXz4d3FQ6h//ePZ4Jv5FQMKxyq+fD6Qh
l/CcmmCRp7YGWmMV9qXq1yRhTvEvYkVm+QaifhNw+n8KhqCpvd0f+E/gC38w
In+RR2xsn2ZII6HQiKu+wk8JO8TAmQWz7Jkh0Gwoy0vWHLsf9X51amDoq3rG
j/imdK5eRXF3l0AD6fFVU288hGxB/koaxigeDbvRnM8pwnoSHhqgLOo4tSHx
FUQnx25tGPcqE7QBr0aO/YowVwEyFSGATlNNXaR4V2oX3z2k8R+wC/MRTX7L
o5X16YAzkc/nGBELcsi+pgH6bs61YLmAoex680ALieONUK6wSuk+VFwTuils
Z9ooRjavxuYcjOBKxYOfhELoEysq5Fpy6p/HLCXHk1I6Kn81FVqUdHN6hz3X
GDJW/CcP7VqHK43zBhUXY9A3ZbWsrZGlAooyZJsI/Ht071CN5c8g/cWcbIYX
l41bzs+5RD9irUDunDyKMDOKEkVzbLVp48mcq7cQjN6D7V2i4JPZyEoLb0VJ
19pHaRw8cwYgodkluZpK3ggGXX+LZw8R0jQgc4+yZ+KCDGYwmX1TvIv12Cp/
ymB1gp0Lg8Wp0rNj3LrBTRllmJBmom+oD13D0JRz/6V8Skw6F6iGokv1bF7u
wuFn5qui6yS17hhvi2s9ZUkv2w7CJV31YLejnwMLuZATgi4E78qk70TiGYWQ
yXq8PqpHz8t+cQ/RAItTjkZH3Ab52XezmNiz55EDuMcO1/HpwQAuJggaLZK1
C+VwtpggqNoab+8EgFKyZJRc6NJsIrqTmrIIAEro2VrTQPdE8HvKP7GLZIs8
uouAwBEP7sUMn9p/2sAKeEw2SQDln1cbiXLsWC4xxEyy4YPnyD7A9TFBpyjS
p+supf6grCTW7wuRkdYFY1vcjPin+MwpnfMTER6enKQxFbU3JLV7Y286pqN9
9svxcvkftIX9Iwax63il1VKrSimE0ZIPJ4UaWZL7GPKb42PNesxCUpRslhVc
L2lVAyxa6ArVF4kJkh+jz3XReJN8fTvjZX3cXh1NceqQ6m/zKj5KckDR7Y3U
upplJIG1J+DalxhzWKmQm0Q4PavYFAtZYjNcZHsBG+9yPyY8jsYt+IlabB33
SrdUhG3Yg1wSTlXmFDQxOUVU4pMOsFlslY45jZoBtm+puNuNKt7dw2AaDytr
lMTeURgt/VwFTKZny0yhIuhBx4rGwHuKP3/f25dsE3dxBIt3saVmmQ8b6Yxo
q1hlkuS1FCF4XZYrD0ZeGQN56nac5XYU/gdp8OuI6agxOSYw+jIggSPYXefz
EBHrBkVNzYP4iEaIHC3qFoGm6Yf4PynIhoY+HjqmvJRaAm/rrrCUM17TZJkT
eJ8IAUqdZrN83ld1+ZJRk6MHJg+mPbV1WsUBOafV2lRz48A2uK/R3ofS1d1R
AnMkAH5Jn2riTFEBSHNvdfFz//v0L6zIwF7hrYClrzT3wxW/sEvegGri/sPs
C5La+jMjldP9RdOMaS8gIDywcG18toEQpPXflrod9LfZDqN/9YIl1pyXITJY
MmTanwfvTOMev+qmvT2apoAGVgMaLMRKv81EPim2jCnQkKFy8pksfX4/rxyq
Z4qB1zBj0HbtKpBVpUOkv8lSjB7RqLwbpyaqYfT//koNrt/t4f0yskRLj3Gt
e4YICmzuKR2vr1bImu4DBCOOLcRHnpY5HKqCaRR4Bbd5jozktVdtQCV6e/v7
cEKbtZVTnk3Dfo2zSoZOHFB9Kw5TFBp1xkCYsIHscvLIuAa5H6oid+5qrwmo
iQBAY3kdH4WJFz1PCtbkvIl4BrQcd+nVNt+4FFGdaFRJM1GhoQQ0HDTdapQo
pkV8s5FPby4RkOoTk5VCSGxOdFtYIwBLKmbro/rGXXFgH+Oi5T395PNGUa9k
/dwkZKPx6+Ywkd08605vM5LDycz+A9lXU+Jvd8o4PKo/GScx13+INh+vtyyS
R19BaTPlQWJJXE7QPUHxTrjECznQLAfjI9C40WPDw1clcIOX5qVqzroGmQbs
CzyMC2uzYCV9vAVUlPnabc1IB+35wuhA4pjyqqCC0WVnAylRFeNeOJa/oiMS
Lev9ms0BcJmlyBWWoc1D26v6LH8faeI6A0M7cCKD3OX5rT0UGHsd7jIZZHdG
tm/3miq7aKudX2k/SQQsn3bhaziWhHjaoNc/f1/AjRlZx2eP6QHLtgbFVBQ0
O5TIeduo4kyfudfEcoTJh4ive7CseRTzJoTVcC7b9gJcFCyMIRmWrqd5M9xa
JJNcw0ENbxk02edE2Fcm5bSv1C13souHCgXLi/DqP7ZAoVNXmR9KvpdYaF8G
kL8dL+Brwk+xB7wn1c9CHAUF00Ld+tDGRCnjmwuEARJ8k1WfU2+xlFWwh0h2
VQpOdUTRuayHJDCCApF3UAqUKbfNjQfcLGgDfPdGXLNp/0r5RPAktvNbRJ7d
h4+RoQEh/wQi8lZhzrYub6o+lQYzEBlCTvqcO280k2pn0FhZcopNFiZ/bouq
WmJqooWdvua2q2vjc/zhzyeUrtOGw7Ul+Xbjwlmrvm/aBxQ24gs/5kulAQdn
WKnhZXbicC8EEAEtCJH+h3pGiARjTK2zaW7/5jHeEUE8L/geGQehXojrGSQX
j+saUmtaqIHUbpR25AvDDJ+4OHofjHzUuGZlr22HCWVhcZEEKb9Ubv4lLrIw
nVRT349lecRZIFgQw+DtCWXB8RVmyjvSoDTMjK8qPvnldSDV8nyCT3RmEkFg
hSi98U1bK8wvKUNy7BTuKhohsZgjVblYWiuADQoBgMoYxtcdAYDtSI4zCwB+
4QQXD1CZcaQPcIpHlVr9Au6K3wb0faEm17k28O1yIJQPqmTcMFr2mphHS5ts
kYbrJnzzKEmfCr/Byj48gWNYTpZS/w9k44j0+puKvUwT/WQnNzqH5KL9oo15
Z0I1+Wp8thghwP3qUDbcXXHdOiQIRYOVloLAn6ysAUf5O0uxQSWa1CXvI/sh
egEfbKGah8HxlitYrrYD6KgT2GqvP7CBiC6xQjDkt1F5r91oPHzAgokhK5N0
/PCJzNz9JWpiWKo7piaQ8pgTU4uosJsAUfJkkBg4n+Xxbr9ZLmVquT4hzm0U
F4KMWHBOfq3o8AjNThZywxMmMug522emti41edpoMMxRgmOa6YPHB2fIXhNd
cFlCtp7KTCa+lT4FNH0PAyZLkd0eBamSQF4JNGfIR457VVXyfotWPs2aRp9Y
A4+t2hIcjZQ+wBxx11a1+BYovdw2eFr0t3Wgw/hGDsbkJLGpAKR+0cFtzIcL
QyI8tw7KVO3+lmAnGs9pRnYZVKLtxZohFyO9wMeXxVBDlolbLBVBYK1YehyR
cXh5eSLAbojG1BF/B4rll79Uj3BEe12kwV2DCqMfHFE5NIk3G75c2hLrCH01
Xw4W4Pce+htDWw6k2vPDaIcMiFiqVXgTHGcEj+gVpTHF3axRhy0SMwc0lQW+
y0gjN7YhOTmAaPjqImU8t62BBZ1y5KMcLtYIFGCGPFuVoHSteKwZdjfniGm3
XH+DcD7gsNkzEetEMFUdbnCgdy7JSoFK7eCPDQGteVuaUl1jlm9omYArYfzT
1j/rN5h76zeZQDX9cH/T7LEHQawrs4eJWKU25/WMnD+GiIM7wNexESl4T3Jb
upv4j/wIz2tZtDcXeibmOZm6PpqdOoQGwdcHV5WTF195ajssLjrzHGL88I7F
0KXHEXYdFB2mPiifXk1NoRpKWVzPtpT0mX7x6iOKLygZKufO7e/Ih/1ddXCm
Ix0I+CBFJOS8Ofg9SNTgSwIfiDMwlbxoBb3zcBr3319GctmbDVOCXNkL6xDG
5DGI0pRKuLsIR3V2o3U0ue16CS/Jtaib4oDH8RN3NRhIdgZr8BQfqFhGxmvv
cD7t1W3Xr2XHe0simd4S8IoTJWIPdH3KfRzm+b+1OJBAaaD35wmzRCQruiOi
aT6v/+z5Hpv5rq6cqggrOXhZs1B7jlxGi1wtpUAc0MB3qyN9YTbnYM1mWLdb
LuQylgtX6qQ34h8QO0Q+T2jfLo1D28IL6czNF9DMbEif3n7RTJ3tJEgE5MBQ
tN8KBBXqQTwU6pqpr521t6o6Q38y6fTcIKHyFchxhlY11DPZQOvayvOgjC4e
/JMyYjE5iSGcUuvH+omtCVgCIvOMJl4VB+cKkd+AVKsmtXdo35Q4bnlNg+CG
snbTffybGv4F0HMLPKhyuHKFJjaXomC9HVj+yoD4MsS+6r9n7/xl5TIg7iWL
l1InWDv8L+TeN6Vcvl9AvYbOjwukOckvvB9Bz2B8Xb15GhXp0Klk2RyrVKlU
fMa609maa0mv2gbZzK99R5Dz5g07ecYARRBsDqwEKQl2q4uvXrLRBTKguPWv
bj0gEUTcU+MmxxKmUfAYSnXuu05r33MKkRCqOsEwVqLpf8v94dV8YwcR47vL
FVhoI98dP9FvqR+gjqYUhH8xsrfcViizrX/VXzhUiHFXT3V+qz/Kg7rJ+haL
aefzcY4Pg98hnz4QTUMgQF5wGUHdH8h5XxFD82o/3E0uEjZ4vc+Vi7qeqCwK
1kpWJhLBx7zaERzb77bL9N759hcdw5vAlSQ3L5FW2nMTLHUuwOnY/uJ+o0Ud
QjKCTJFOw+OTaFLBLTv4o9DFzzQ8mN3LM5nLQwLrDZUA4vb8Me77CsgCj4Rt
tB0GnHXXq/Evky+tGpPjkh/po+oYICe9SEO8UmdGjlvF2Uw583v3zgYjnBjc
Yr7IXE6ohEFtve67UyRCj5/tdhnsQrAhoXdcRc7Y3bnyp5Vic5+khymf9UTo
+jO78vjAPgC2kj2kiM3ZxM4iOrytWIMnfG1wvEaEpa20K3S0fDtBmPNG8fnB
YOsL7b5antLDcxxS1htwWHOzx7fiLyL8v82h/NL5Jd3wsrJdDaTmaGz7SF7u
cWl2jsiLIIye6c3QNqarUewhyC1+Sp10+N3X446GUH7AtMZ0MoNrZRZHYcEm
WMsqehhYrZJyJy8UyAfCW33Qp/WITN2x4Ha291KqviXJYIKAV2P+wqDj2Dj9
p/0GCdRfk2z0DlDjj8XWZ2ECG1l4txB1koMIqEmWjeXtrMqmk83iKu7zRWzL
vFlLW9RfwW/3CUcmRtJkwHgWEj00dmirxQ9pl2Kc45zvGr8cRnbFQx3Bg0x2
ytk+UxyYXmjO2lof4A05pXPy9j5vbm0ZZpOb+rETBt1D0gM0jDloHaYhns2t
vkaOekOWfB3qyvBYHyk4zO3gspguPG+Ccui+ySVmmEj3v7OsqkWFsNCQ5wQ5
HYxw8tBamvetCoR3F7en5SqBMJl1Oe+s9FjssUFGi1ab3b0/LirNg7rN7t2r
W0kpnA4mP/ejLsCjlmsIuktALi+RxXXddb58J4b9rR7wYNyeY4yFagDKmBp7
QGL65EaFvfiDthCQuYsdFNMlzCE9x14cWN9i7ngahWXtAGgHFemvRio8mfwX
KjFZmgPet325sCLJB6/k3OlM1NouwBmmliSKf8Jp9pX9wvmAfg1da2i8crGT
wXxqgwPS+rpN8pO5l2tAqjsosGGpvRIIZ7esbbVdSSQ3HZaY7ZAllrnc5Ytw
yicpE6fBtWRdIAalRJ/gInDCEV1+IACospqjcZPJFJcl18FsWtsAKjQM0TSm
eTQ3561EL/18QuM6w41J8mVhKxKb/Y5LMuFRBqj5QhLTBeSuFyddk6+Dm5NX
Vo2L6F+/qE4X0dopBAon0l2rXxHV6wfT0daMSf9rjIGJUIGEO26KSZD4Cp9E
cRDjnTOP8fe4KoHSwpvjaoLW0oXtv0KjWC13mjecmYxmgzkU/WpKLsZTdwGI
XHjZ2hsEIGTgUdoJ9KieBXThLyze6VixR4KscZIOgoMVkNtPCfNCiiBlZYFs
aU+OocAziFN49MiBGjj/foqkkuX4pGEPeHrAT+wXJZaVsIXrmqjnQwSosZ6P
w94lST/fkd9exfPwv2BFekBBW4r33swkvVlEdntX+c0GU8MkcUHC5s6EkoCh
glGlA9oTUdOIkE7+LVyj+mRS1zBCGNd7ULpMLnxi5gG5bCGBX3Ai86tAcTTO
zbEZ24sXxieuJ0/xNcLLr5zpOd4CfdIevOv+G6iP4bbTcHAh6JM/hOIGKMD6
icBvOpAF+06eXk6zzedBYH27QciZ6klbccwGXkCUDrhTdRpbd/MV1RcbHdZD
eGEVOIdfjPRxUD/if+k5plzSb/ltUrnZl8Qeb0TWCIaRXER00Sclmggz9YzG
0lRxmf/yUlZGN7PDgytXq9kN5Kf+URQ6HhWl5d3LjYLT1Z4c3s8dhRr3xVby
7UU3TIo7diNllIKQS2Ii8kPCq/UiMtHLo3FRstC8BVg24JV6j4KdyedvwVDV
WrZMIry977Xjn1mfadadOB+Ji4c9VOBZRP5uMtUga6nrQuRZ62fqN0PNaZrA
m4edIhyLqJAYYGhkcKQU3SHvgl4fq8ZlRTTwf6ICf7/EAa7nfD0T8A5gno+I
T/IuLmNyLvrIvHW6sIi9dFBeB/DhzoBM65sFF82ybfREa8Qn5cg4ctCDLLwN
PRzqFOgj+DSY2mMoMC3h+V4+q+RuBhdgMNfycU4qc3oL7X/JUehqQshtvFFT
COzgsCZBE/qXxk+FosjetR1jxZ59yEXd5HKMXSCk/WqceEISlIDx72RhiKhN
bQSQaoCoSiZmDGdA7K6fO9GfhGjjemqbrZzqt8XKVOFlhJucGrgTxjOw0+sK
VhKpZtOGsjZo20P/LDGNYFkHeXHehAH1cP9ehBfsw2NcMQFYkAfdGaWziQBN
4Hs/hQ/eavQT8lstKh7SgOlHyINzNUG7lFokqcAVjYOo6qmNTZkbUDlPzqIX
m4viEiWFNilPdi3rkRgNbiihmUh8dbGmfdARQBura5IXh0Zh2tRc+QwsFIvG
EPLdoSJNbtKJfVmat8kUUBmrNCg0gmZz5pz0UCxt1QLVYGa3e24eWdKWjPhC
f6+HIkvhPP5FmIuCspqvfPF7xBC8Zv/fP1u315tDs1kUK81tTefp+Xg3XMF0
Y+omGWlzLaa0/XtrFRc3SL3V3QrXFcLIRQj5zxQclXvS9D8QTs4i0trxvJXk
XY42jmFjLfYBQi5IXCbNCWcUrflbf4A2+DH9jQtT+xFOfl+SN2ZBXyqQxbn0
2AD/EwOfnpkq4RZSYdLFzr1chNq8qZj4Qy9jFNSZOiuZW63OTvBwifZymHUM
6He/GereYKK1b2Pm/56sH/6CoHFM2CvMPFDlX8cLtun8t0NaRbCbby/0Zotp
EiBNGMjWtRcTZY15S4tEXPZ2+7b5j3aYu350RqqL2OJKiBuruMdJzi2Zvisi
SyBjJbos/+cReWe7w5LVjs+YmTsbP916RMRZRmH+KWjDavjg1iGmxVwO1rff
3JUlpbowr2EFWscLAsjfg0rTTpzftDBqwt0TBop486lLPksOJA5jCcn1guJH
uUQ6rQanohvIXaGdLB/YP8csroCrfKpv2RqiZ1+Ow4ZlAPaeGighQ2gc7XWR
xe6YWsuWoJisGnCiEEWtzjCNi84tbQilm9UNfV5batDsMQeu3gqZn3/pLsMa
edRAOxQLaNYv6ThiOXLENKxy6qZzckjlILEydwYHFIZ20y9v6OeIiOCbG7Ox
cNI+qbRKdlWz/ft9Oxo6czBo4jjEN8oOxtwIU3Fe8a12uF9EDO6VLjbe8vvC
CIlt/P1iI3oUSBmECJ+yfM+7eE7YQQOcs4LP0un5m3Xw0QJ46W2f6McHYWp9
Wgy2ePVZMky4Q60vK+yEbAfZAbIZbOcpsYNac7OnYqol9+4kc6YWX8nph/Ss
wYeT+nf06YisxDwQguU52SgEpITOsgt9Xw1BP/zb3UUEkzBMRg7rF70q7bc4
CzUbCzWuDZGKkTY2dnolhO1jgxzRcq13ggQi+GDA0KEEeNZY/VyZHM0O14tJ
z1LumWKHvuR1N91r3nD1I4NyoZiD9TkCD6IXspZeX+2rzr9hezx+FuEAsjZF
QdJpK4TKGWX5W6RxdKVOcKGyXWOOJ02asYzk4UmR8FOcSAtt6RcyN31mQKGs
rDMrFECFf8+jDNiZ0ZXB6zVZxXZ13nMcUlRgYalEzxlsRen83VnsOMLS9x7Y
MRff/+TRXruTIo2NEFVondM7uaSk12hVSYlNplKGOhYO/OtAFZvLOkq6RWRw
Rr4UaE6UtaW2U8Pwi/Q+vJdXAtAPB5iabyCX/G45FeEj+09QIVzjcKtLB0u3
rjk+GDB9cvhjbfbDyzASt296BvYUKwBfQg7o/M7X/MwBgqYlQ7wJirYaKQde
vQuVnNPfLTl3yjEm66NdV6TBSzlNm4eNHo32JiCx0fUVMNeMX+qhFtksrjc7
UlRQ+/qlll1SO9j0eMejByQUyQJM9roU++wSCa7qLMas1VKvVxDa5BN+/TBm
9Ra4jcWd3d1mm2xIFpewzatOWFg46381UCDy6aT45VuX54xrzHa7guoVfsyF
xjopb71Ej6A5T7RFG/gRg11HwRrISvGwJ9rhXQ15z8Tsp6F2qmKsZPYAllY+
dC3Ycq0EZZQg6xYCg8cer50XdYPHUCOC9cZRfwXOwJnCMtF7ESs0uKE6Ql+o
AfxNGhNomjyUrEUM5c+91kwEbIQ3ivT9Xzp52vyNhMTPNEXFC1din+326x2T
CFYQ9/mkJhsYg3oQY3xaXwlGdi5DsnSbjoN2Gs1Fr19NcjojRJ7bTBN7mIWx
p702Z7d8N2sVPj0f2DLpRRI1ThF5bBdyO5QuTNrAJzKT9vx2ea34mkWCyzlP
M9Z3Ig2bRi7smkYcv9ciLo+MF4oRQD92ZqzgHJ8fgxsSX1TAlWDx1/jhCgeq
Lr3B59po8cJqSozQZu4c6QH4Zo7rvAQt6G1UENWTfHUxeCZnsfX4BhXpSPIQ
4GD3iDLRBUAQIfLTBwRdBY7X6lCyDIHFDNtne/Nbf3sRcBvEdMxI5nQKaOtz
tGvidh5ZkIwD1VlRpnYv1eetd3GIN/Fnk0oQo4H6kydQEE/PRuEfA25my2Xh
5eYFfFA/X0mxe3E9J9BOwKDjLJFQXcL1MrfUdnOAjVrHxJ+tKK8A/RkHx1Ab
VQ9dXgxXGRcv/NvOn7+Uxx1TOU1OtQ1bH1hMvUCbQMscYx+U3a6P0mN25Zw0
hpIK86kh711xsPYPwBBDLdbA354s1y6+sQOlYkwNyCaL7ihrDsTpadQn1qho
M0OITRpjQVMvC7mzsFbbSmdXeN/Qde/u14F+lkKzFc0qeNFh4ihzSMaDB/z1
gmoCj03pkqH+JHwFQcUf78TSJmjpKa5dLIPX6aVbyCgZgRRKrn6TRxBWAUgi
1PGenUFhuDI0RlJhaK3gdV5YdlNOTyrfWe78xg4uXnXRbxtv+66yxUAQhuQM
NlGaRx8suUfURqn1h71bGQudKgvwDH1Qi4itJeSYJMjPGYcEjtJY1BtbU6Wp
o8ArS/B4EykDesszrqydtibnQPyeDHE4fPKw76yh+q1tJ5UjAi66eJ1iDdeB
PNkPk7udrBdokN0KBBoAKBJH8mzpg8FQiNrJ0dYn9DrPfX5CIj9ed4QCiU8p
ivWfPtJYhnt4CKe0zBQkyGBstVcFFs3keeMWiHmHnVweCQdCxgG1Ds5sLvVL
QNzyUTRQ9g6AftNPYplt6IT1XkPYxmkFP10XmzoQkW58uzILBCJTJBlOZCJK
dVsgmIg5X7MDqhQY210K8nrz6Q+8wa06UHnt00l5VPRPVF3/5+am87efQXpG
wpIcy1ecsEmpBwjhg/Z0OLCR8l7NgLr43xh9G1uHZDAwjvpE0JapArfcPBA/
gYtU+MOzObQOajNqXjZw9RCoWwym5S2pO0svJtnACcSiE0t3256M6TtW71Hw
zFAKgmzoOb9EZMA/0gJcnv7jSMR+QvUaThPfOMbtDgjkL9e0a37ZW4Yhs9XF
6DZmIXoMSYmS/lJLACaBUvnRHfP/xr1wQ2/XtfsuwMEzk95R430F1i714hf9
LawwOO2EkFm26PuL1x21psVV9gzszlKOEfXAU5pqEH43PEnkm3IxW2iIYZKm
ypQulQq6rRj021+xJ3BMeAsoIsyoHHxXmUq7NeMvx/1TN90cJKu+S4bVzrUW
L2pCb1MUQPYxERIs/0DccBxUBVN0kzsx0/9qyq43rCtAaBxZ0CUIl6m3QeWw
MnCdCQV4ZhI38sldExYC5nq9yDOqzrjErsC8klOzPyXxOjHJ2iuah4letceG
wRqEyjGqPz4NfOeh61L2tRuP4cd/1U4MIHtgHC7PzjSSwDBDybv7372H2jdA
AZIzff9b9X59Wiw/Av9dfXYKfgZZjVDpi3dL99NdujABDjWCAFoEkVA1/VOS
1RvVpdAIISS/0o7/gYqoWPe26aCjstMKJu0XqJX3FyF+VhrmoImClcRHpt9v
hLdGsUA073ao3h570v9FUipDAVOdCxDL/buZZlGwOAhlh7VcDcGFSK27iPHL
w96Fq1VORNvsQHsGAFeqMJNeU7bqphTMJC5a2CbB2rva1vtkKNcG68uvZJzX
SjouscvGA3ql93RyDepvkW/o4hVo8IOVZVSYO6Ii0I+Yv7q7W1qbF0APhhgV
Lw/Hvuj1Se9tIzZENBaeOq2M2guLpcDH1Kik8WylN8jnNQTZ1nmmaDvQzDaq
+aYKdM+RDLrGMVqUWKyVXVQgDYLskQotWNZjGFS4+Sn4qlvgyPvcfKzW/ig/
ebUWVkos8KLMgRCjKTSlLqq5H4AHDknvJTtEniUn345Ia9oMcqLOZSGzRmm6
o1sYeD1PUxCy13XZBIxQlkIYHyoXDUDkyGA+bgU3eNJUFAp6iwH4wohnIDNM
Lrw65J/eXDpMrDNX2daJ7/7o4bGZe4XDKv1pjHU/oawCcDrjg1UTwGJYyN+k
sKN4rHkiyOJfXt3T+B4x0rGkkobbdZmlS9jlUANZWP7xyHh6nFtd64tJsxhZ
Tw18V/e5PUwgi4uX1zFiNN/FzF4vxaOIAkwWZn1C65MdRiLMmq+CAS3fYkDm
8TeHkuZrKKBDfRCv3u5a/wx1YFh9tvID/vWOPoUdPFcUo2lCH5H3vkMekMN/
b8xQoVLcPzeBaH4KFKdQZNdyECHE3pQx4+md/aVHqAPN0YFVc45HenkS2HZi
1/FDavOQPe6nnOQtkz8wYVPJErEaDav/5yc7qwjaVRPb+t+hA5qU4AMCIRkh
l+/a5fXTIocv2I09Ljk4rUxrevIIRkQY9fDNklUZccemMjV5BwtrPSPCChGA
+H7s15lGTfamvQiEbbda0vHokfYJbBDAsE8eLTmsAGszW0AMkQdHoc4R15l2
8oU5427wDiCZLKeXmxp+mzn1A0r/AAvCCaYoNDMfU1tkzfkPx10Unft/xnUo
Uu3Ga+/XEy9qvlSlGOEGhe6svPNFzieW+gj4w5t7aci3/7wbzqfsDYQ/McFT
CX5PmkJsRBsBAN76ObmN7I8AzKNkX1TYFObKAWacZdyS4cDHcfbj9g1ZlYyJ
xdEp1ttFlh6y3arFt4qzvdDCm0CO9cOjbXig6LTPP29k7OseansQ8hCnhkZz
YQkYirddu7doGuVA9HkNFEPNKmR/NcWEJkEP0APGbzad43Svxu86VASpMBvh
7DJSAiMMjLfmLeu0kl+CaKFA5H8UGVh7mG4DJh02JzYvpMrvbiQXawYtUX71
PThcijzXEq2xR1QMuq+dd8ajafV4qR5pNu1XoW+QHF+gJF9ZDH+YIEj4nmla
4nznRvDuyvk0CdHtEWcUo6QYIPyHH/18OMNSwe3BSfLMEGzkPy0sIPC56WNS
vUL/LcBuZnPTDa7xIMdGyuDvtZVmkWwtoqzw8F2G3IHN4027YS4xHmJav/nb
se1K7uLsJtYSPVWLmhvvnZDEk4Vwq2pjEF17O1/1G5ESLH+YnblSLYG8b2Tn
bqbpFLNDIHok//nSJFnhXp6yj7nftfnYW8X8TARhCScn08ro5f6mPw7jQpiL
zIfVDcgo/srVdblXVW6IYVo4EdapaflneHiD/twFDCmWbYs0OkiyBj9Ej91n
Wwj/35FaoV4KFfLJTn6G759qjSw6qHcjY0/dw3wWQEti4zfIQVcIHXUIqoAl
iC+eeh0in5kHYBT6lXPUa1Mq5Qf4grkXBfdrb3SQ2ptVSr0SIB96EXoaPbya
s2iBgJTr9h6+hw7T5J2Y/2s4mXfqJZ3OPw1Z3Lt/ZQYk85gXJQNJpRMTxbU9
gS9FudG7CzkW8GhZuP3gCq40bALJ2j2dBEvvARq9m0ptRtljG7Ho5QMCHsib
Ejj48xyANfPxscLWIFloJfSeqHZu58O8x9SRnGsvRCdVZdzHAWGDEik0NIpj
KrZCTUe5qvG2585tUeYcFV7MN4jltFUOoYfushiPBToDYjSQgDopVr0MzZmE
Ja3/danOB5mhzUMCjb+rDMZN8SawGV2mc2cqO2KucTGoIdFYj1IXC4CNN+MN
0vf+0SyT2juYXc9lFn/6e7rTxSTy6vMPfLQEyL33ZcG/pJXtlgfv+aKp+Ztf
GvdfHMO/0YutwoS1OvGjCc/zH7wbARIlDDOpS6XBIi2Gwn9ol5CWi9D87lmQ
hZ1eteju3ruaewWp4NX811AOKM9MyNawvatqhpTTAdbuNFYksSvgKoc9L4NO
xtNUmQ5WgWKl4aWuav1IK5Sm7ESrWnmsNLr+CEI9DU0uJtOGOLV+5AunTgpX
KMOTD+wj5IvOdJewMvKCPCGYQRAQk8QYHL+Ak6zFPCMyv6G+o75xhnWcYJaO
HrAKF3LSTCM9TXOXA7/vR2yGhD16Xwm66CN6mermZwtJgg32k8W85+waNPav
3/trsmO3eRq6DfoGgntD3bCqbf0pDcWtmYQ6N9+6yW4Iq18zVWVRnLk/4hC8
NxZv+MvprMBf5d8ELFyhcv9GS9oN59wKPj1UPhZNNRcI5vIkB1KZLg/NLp5s
yZ1Q5efURRzOycSMcUoq5JgnWTUtp9/zbTgM/mj5t7LArssEyr1ovTgvfntH
gob40cjj9JnXliBOX7yedmVH9kHGT2anmgFu4NIz0a/Y2UCRSK2sLHFta/gT
AH1Wt1JOyeXWw2cr1D/e07PIpQOZbP5Xs5wdgDWn9Qom+dKVbUfZLOEzQFXq
Qtb6E+hUJH7ojq1P5PJwQw2WMohoAYhJpN4wlta1tzFQIZ8XqiulvTzlRw9O
ZHNVS0GZddLhM7N5XDGElGNG9vREXIbwLQ+B4q3mux+FMY8ge2wzWgROhvSB
gd6DmAp8MCQhnGtcsTjbW+a/7MwXHqtyOZvDCz3Rkj46qjjBlyAKRT4bsGwa
eNZlJtX50hq6iJYGj9C0njvQlAU53sWqteDxugCLO6JhzDg6I6CFk9d8Y5vB
ZFxa5PhllT6ON3pIA9sGZQqc/Amte6dQVEN+L51Ucwv3rZd2pKaG0BrBNpZy
aqaiz4d+GnHdBY4uEKTzXTWHaXGxkTDgU28Ia/TFqk1cMKK5Eiohw1ym982L
U2zzVGpNiFhaWWgYI1v3EPlEux5W1/jvRHJOxmcETJre57vs0mN+7Xj7LLYY
O50xR3chNZXPcwm0IUD1m7gA7GQDPG1XKxFC/i/T7dzrYbKvVSMhIZmaIoDV
Tv8XXAS+KzA43C9bHb97rMmP8iK0D0FXClK9e3H3Y/Py6cHwceX9+MrLUcXS
L6js8xcXsv4BFiDMSsoF3j8kvjktwqbDmpGrLW4ZpA6rMP0rPX3WR1v+IZZh
MFCYnV+ERUxnEZuzeOKM/XtmYgSZKTAT3wJe8GU7KuCyR2EHUZQnos+9gC3z
8cbd3re1x9MUOnqg5ZR6oiibNUpwFcdJAfc/qIyqmKgSFOTB3T8pj+J3FaFQ
3W5mXJ7PtO8qzNlQhgThBPeHmKdjVI0Q51Y5Cltp0kMjFI2un/dMvPNn0vC9
cL+xvZob7tl3Pju0NU/5QzYqoY9a7MvnPadLuBPOSUkEk3jKQLRj1ZFl8Lit
yzyryT0p8Msmtbs5irL9t/wnEjq6X1/cXDiwpCpuvDnMa267YM9BmTLo1NrQ
zk5JRrof+f7mqF9u8wxCYD8HFaPt2TM0px/JfEzKHReH9qLcFt/AreffkqwN
UoelkotdRkCqgDd8Fg5jFmrMTOSmT0kc+n6URQ4psXpRVXl/khrxPZnUzwi2
oAxgWNhYemBgyIOTZ49abT0DYGgVdUYaCl7DINtCKkSCfFCo7wY8f0+5UGeE
VBIhw3wqpaPuMvXk9unVdoYq6pZemw24htaeOOG3BT7eiEQpccIbg/Kt2LAe
QOPwtHDuncROh8y+0ePMhiKrNot/J+7gtPpKC0w68rwHuxq/D/0stJxF+BG8
tMWRy50hqWQ6CuAuN9bOOK2yfofRJkJKlPo9x3tbSXcVvkqgzNPvlTuPbtQl
2FoUOI0X0mir0ZFa5vix2ktYGbJUeUhKRVsFCws/07gxqorMwdSA7N0PDLaJ
QNmRgz7CmdKnovu8j14VCp+Gk/7daF/oVJpf82u576aPmKC12jaGPBnnvkrc
aq4wk4iMGhE4sqaZbbuPtZsFtURukyxgLOIOfsLWsAykR6l03nqvJ5sKMtwt
R3heqtiMAanRwFOzRWYHtj2IukpId/Qr3jgkEdPAaHpuiz77yTJufvY1MHoa
hLoLCPimx5iumz9PLoWkz8tRSqP/hfJLhuuQaIEFif18Xi9oKdMo/TaIdFz8
BTjGgE0OO9MTS+YtVWnF6gos/dfhu9sxz0Fkqcs/xzUN1LKqRdR28SUZ0QFE
f6tV9qQhk0WBlEHYMoCADZGENCKxonHbYkCyhANB6cxwzVRdhE+LF70xbGB5
IBjQyqmbJsUpUAqSqP3XSebydAEZYq6GBHwSf26ANpqw1spilUB6XjmgXVBD
gOrAwZabRFwObmGIdE0VCjjA/W8wbpir46o+clg1bxT8BBbj2r4kh8VHB5Ke
4NNBB1T5GXQV+enjDrwepv7BQaOxUbNIMYVTHusAX7k8gXNd4M+ecUKwGJmf
eplN7j9H7I8J3xZXCSSnfREUFS1z5PfVPuCwa09wrMV7f58LEbdWsJBhDoqM
SHx/uyI0Yz1OAoJAU84JcJD1ry5LNN2qcgg6FxWac39wBkHuPKMIra2J2gLw
7+0SGwxlxbl7brqdP2i87q5WcQifEd+yFq0ewbv/hfZVWZZYMlB7b8bo5pLF
NpcMf5oWXejbjMxonfDjXlXAtBJ9dIu2z2zOQS0lOEavQaiaDxEIlFUPKKVp
yQ/KyHWopyw0t1Z91DKl1zLU9a92lmkr52RmOkzdRFtD1+xFi3DbF3a1rWyN
xIyRNRq/yDnPK6vg1pV8L5X89NmpmOhAGA1dFmO91UQWdTFHGdGRu3tpvSp2
N/3ZsnVMnheocX2GRjxpcK5b6XWSL7O00K4wuv5xW7d1XaY8DZqxZBw7MH5S
3ruLH7L6PrPxUm0FJgIzl0I9UGmfY2urgHnaVuz8b2jLgaQBJYhE4kXEmCBW
R5XVgXooEaRUEaDu2xrUw5L8yKSjXwMgn+mVIlf4Fii9nEEGBfYzPzXj+SIj
z2b9tV1mtwbcen0Nk8UlXY6FvNznojEZLu8XC8RmgEJoA7VV9OP+Av+37ngB
Vlt4e4Z8xipFlAJIm9Q3o/wh9cPO0+7eEIDdl9w5OaPFoXBHH0QLxeE3pGab
2KfHA2I1pLweAqMcUJ255dfp8VuZwVOHvy1/KyO7QKDTwn22sQHoT+FmcRZP
KhfAtX3NyH4wX3AMboQWkXW1cH2/OsGSBxYlR9dVu1xOmoCeYLChKKImIVXY
0Famb2387ke2ZTejpWGlXXAoHvUfPsiinqVDTrVEUR+Gh1SKD/QKRgqnAc6B
F3NT4BY8fOEFXAP6/PHGu2/cVP4Fcc2s6xnVxHR/K1nXoNE98o51xCP8jIyV
ozT9zCjZTiDygyr0NiOGSypDyGkhyfM+VS/bNWsCofzG8h3VD7XZl1M0CKzn
O1GngAp661dihM+GDWyURiTWhCnSG4bQHNxTvb9b4ctoykG0QT52U3ZMgIOB
Jf4ruA7b/dVVn9oqbOdhvy4iSR3YcMexPdDjRtb/9DX5KrE/b0Rx0erJwkqp
Ok/6j5dq9zI3Q11YBj5BL2UnvnBnFNvoUUbhUROLi4FIyf9BoEjUju8wjj//
CJQUQ1OdrNX4TezG4KLQbvTtMX5xHloa4UutyZ8PgV72gYsJZzVpPvIeub3L
p/HOVHPjwQKTlU+9p0AQjaFelwnAOvCzxnS8af4ORl81/WmbJ4F/lGwKC0Sh
6EUobnVQ4ta7ZznHUIeTe91HAo3QEJVYbBIC7d/atnB5+jjQQq7HVAsR9M5y
Ogp9ngxrE3HMbE/h++BrOyDyjBKjAYvrgpgU+SsTjdW+3EV1oBF75uCuVR3X
Xi/tJ+35RiFxM6Qs8UlW4SQIO/OTylhE2VW39MU6a0DkM8gjB2vm9W0hkstj
rodRFMxSi/3HwaU6lTQmQkWC7sNiW6D3QbjAimK0Oq/6ETBa4JRshqUQz/to
XmfrHEbpOi2fFt0zgh8ppjHc2XcGUq4CqBu7graif0ELuV8+gMVFw9fe/6wc
WhwsdNhws6BzPElKDeVkHfZn5at6ATGrTPRiU8o6Btr5RKNfsKUuEu6ilY1m
w7xkl8M43vv0J5ipu0fdHQSLD2xPVy9gyC+7SGGuTg54ehDucsRPIjffxuc5
roaKl/EmgXfM7Q8ykW8C47mbnlCfeadGYFRCMEPuPG6bl72JeVefCXsSnbHq
5KaZUXPHEg7EaW7KKXD1DIcoxV8wfJt8B8onBpsq7cuzM/BqazjvM4s55pBi
v5TO4FsxGDAaNMya/3GyU35a2HVH7KS93Xg4SwWtpHlWEQOjTmGCRZEoIUyq
Z82AQEBzrr2lBjU3zh7wj1CDphpSrMnAyt6hhW9cAsduNt+nWtgTbgF44exc
Ow5u+b+hwmiPWNpxW0ci4FK/0LIoXuPoLVEyrl/sfBaEZ9v5Yhe3zRjtRN/s
F4zJH63MDWydhbfzx1p58ZZkRtewLxXYt8F4MhVNnmvKEAEKN9QeOq7J/lVi
WI/Cwse7Jr72ecKg3ft5pJ3Wql84ZdJW40GDgrPdG3Yra2WkFyvMqcg6BOQx
W66DWmPDfYk4XhBDuqdTJ+GEAAPw33JSmy/j7yjCrVYioGmVv6H+FcXeLZwA
Ql39qqRSe25iOTgbH75jyFeMpO/LzE+aSoJSW0vQb5VF6Qei+0ih2BB6i1Ex
jBqFVx7tk0LYuDZd0pjAGAFHTvoFormH/uHMaimDnZkSCpnNG9JaxfUGYgmI
3w+6qJyy4AFbrburPPym4loi9pXh/TdmF0ri56FJ3zq92dJGt1xwqCutDbHL
QUGMPPOb/lQfJ9te7Q84K88GV9rhC01lF25AybJzdtvTIoTs6IJUbMaiLhQw
0vcOUDohix1CND2znmNMK7bkGG/qCQjpy4m5kXw6ZoH3PkPzBnHuyODAAYzu
45I09FUsMnsUtgdDvEKDpqA2e0O8I4K410baJS3GDsyIa6b8pX5sP2Pbby0K
IKe27MRn3Lek4Zr5rZf6GyyYG2/UT7Pl2F/j19zjyJKWVLjopxfUnjCKeR1z
UtM98kruvWYTeKyJzSOeNNrc9bUphYejEaVSlY5mkpaoKU77V5g1Lk9dTPkC
KxQ66NnLjmUE159rzOLXjJVIGYf/dZt8PJNbzRNKWIuvDIINUrHhiaZ3DLIS
KRMxekyNLD3N4+CbXJbIW7UA1E8LjoXbcWQIMSjSzMvx+dDZD5IJiID2XR15
UADeWokwvnVPe7N2yuvuV6WOpgrST5zfj9Mf5urMxkTjLMHoAVJVO5+fDQM3
OkgWR/b+i8vpCl6l4nCAtq8vTaxBI2karsfVDzavBoZLubvZc2dvqJTv6m6K
Wqd5xzmT1Cg7GrEEFZTaR/8Ch7mR+hNZ8NmZLe/4d2BhgEmhgJE5SP7WgxkP
TNz2bC4ILhs76ZvhoDNggrMFA9kqglV0ul/Qce6djyfSagHqbmaO8QZ5xZN+
TAqFd4I5veWg0TuLftlmSl9aeM14bjaleSkr8XWpsmhJjhcPkCDMWAwr8Kyp
SUVze74H+uB4oEry+r9guzWnVGlahYrQHHm4ciJc4HNWNkwTbBSKkbYXP2is
BOSip5Wu4ZjjmCmITKUTMAaRLbQPTZIZn2a7tKz5rX9YHUqD/XLSt8zfbmWK
WKzKydM51hkyxYljMFCFRup9Qk+Ldcq+Rpzwg/Tqg/Ba0A3o22lZcPw36X+o
Air1sIpZHTlfCAJP8zHirVJdllCTMgLYqKDF33/0c4vagQibiDR+qA2i6O9a
D7Tm27b9YkgBnLYwtSnq8S313Dv9IGl9I6vZuMr+Mqhm4eNqPdtCznP2YW/E
IAAWGANAXpWFL6zdnPIV4BAHuUglnS42Vo9ywkC5olzIv7FHkA9N1+0owULK
ft3wD0pwRwDrIRAObpa67PyKGqgj0uRJh5Rr52i5nf+TXsbz9VclwS23C9gp
NOpt8WJc90MGrtdYMmEse9RFXP9Z0qvZnlAcNbSjXf7RVAsPtcFoqYkeYuEa
n+1+VIhn881ZnIHgBvDi0J5mz3LpJ8TUZHJ6iDcEEahw94Wffu2V5paX/al1
0fdUcowjfCjIjidO4z032VyFtOW62PrK0AWZ1WHv2YPeUFvm7SkR1b9WCFU/
b4QohRHIPbAWctvEkoRHXB+cXIpePxvclc1HaLxQaNZW89kMK5N/bbCmwOlf
QYA9vwIm434krOMq61IV6VQhcw30N5dY7G0v3q3vcRsp0bUeV5DoBWdSOZ35
E0N8zG7usLLzkV2t32GR0PgyQeXMB9cV0Syavb+lanQqK2Lgmiqr8oWLzSON
ZjcRxgPwu52X7Mwd2zpVr2Czc1yt0dN2Trpv6J5SzgWCAwXG6wdg5Qr8L+sk
7nGZNsn5eQwNyF7CqD8ie8LatyeqyTNX7RG+qLBI1vshNubUd7ZGLcd29//n
VntT2DGQ3ZyvJjvmkeI5VakwVGjCaWrwG1t6jtKWZTJVHfNmrFIdZWKrjzqA
C0UHGqrNb0ir8zRshHBX8QH78psr++X4elJH6TP/GMgynvQvO2wW99QDjGHX
TAHs9qrXG5USq2eoqvMLJOTObl9HZGnPIgQi+wjk6n9zRHGrdU/4LnnaBxKC
1mOi9ZJEXnlT1M1FQ1xNbeRnhr5ogCy5AVfJW7l9WWWU9KH/75yag/oHx9e2
b68EeVHdvlRzj/WBBR1UeaoEhnx5v6rQ7qUcpddQPST7brq2jOfhusX9AOzX
NYpt/Z0CpOkmn/bunmVNjK4t1KO23WDZUIrDKSW+MhIKGVKbh2jsKxuDJADs
BUCF+phCoDHBzqCR0oIAVFNvHLZy0NjFB7xrvmZXfJd1EX4+xIAkJ8H1AIaY
YnUh+AOzhTjb2ncPlYLkcFmjxtbS03IicXp5RpJW2WA9j1A7SZKpYGBXA6zn
z8aCAZ6QB/G/DOvg6LfaDXx7hFiExiFFhF+jSgzYG2ZxH4WqwZXL0CQNZSgA
wW7KRhDCctzVoblp1YdFxVQfKVC+pvyfadomdsVlJ4QXecGyyZgInS+7GD6w
+u//NSj9HMp0DA+yX5s9pTRKs9eHFx8GSUxg5d479Cur4gC9xWZfofpk2Hf2
fZi3wzb41Z6ocnyN2n/9adplk1ATqeIdkZ1YpSg7k5+/feRkJ0sKV7ZCWDAB
jY1NXiPZ1zsc9n3C4v0hxorPGFPMJVR4dPsFQKki8n+K8RLzKvrKVJPVy3Gg
kFvPMzycfVhzRPb3Sumje8n69QjgkolW4vt20zyEVWT6VhjLzapbeAWNkFpF
roNXvzW6S4D8io8MJe2ZaqEgcYckmAaf2GtjyuZtKsfAgcw1rOhBzUYfwpkB
1UR+VmlNgozlMiSJuauUe8DPAyZaMtdqZBwL+HmVzxYATKtEtX4E7lUKd34e
VdOA8KAPwlVwrMyLcc2AFwiPhLwFpHQdnGnLa+/lHm/zd+alV/AKnXkbYNSP
/Te213lape/eTODifP3t6hyLrfFZQJWHoJW13uQRZ8vWnQUTpcZpeZaBz8dj
ac1AGWr/bDuxryLNppzYgn1UjnDGVsP3W09RVDcvMO6zvxAzCUOInGggks5F
v301YmApfsZmCZ3bZfPZz6j51Y2i+o7XVcqNyXKAKMgAapUSS8Umc9YGCY04
ldqQFK0Wy11jgA++3alQVN2jJkK15lnGKSbk9BQZBipMscHvbykHTH97hFwD
nh84tJaG3bxESi3VK19gbfkr3iSdcf0Q+NXrKRtWW3oJW0vKeIJ7Kn6zRYlJ
IDO0qSCd75bPuVf4uZGiIIVU1hEZIqkiAP+dMGDIVdGdU6Ob6Da9l9KZIv06
yLh4Nl/c6T2mpUdsozGqOfzv860NIgzQSXh3SQni1foxohe0f+p1VODihKYk
XRwd+CflmMGD+3FYjnrzCryY+Kiizh6SNq91DJXkB4lo1WlglOT1x7kCtpWC
8WKTwt9O7iTRkPrPp1453EyC4S3oTjddi6hhdz/sdoqI4SFdIrBTWgmnxVuM
bfM7zi8iwWTZ42bI3oaC9t1ZQL80KUWrcdfvZD/vn2d1Fn40byuf8kUL3WQ3
E2Ioxde8hovFDxS7zT00vM7IdcTKmDrUisSXiXpkWqnhXcRM8E+5Tu2ktW49
1cEt4iwHjCNX1bOxRkngHl9HizQHpLsmSc0ihRCwvyrIEaZ07md+qantgwn9
FZK8xlwXZGTJ0U/ThfqBwoSpVFghrM1VAAoWRBVVPM3EsFGuArVi1a/VnK7Z
Dxxy4315pknYhfamZQFDFQnS74u/fK0QcasaOnj/W+Z1O5fnar7Kj1YBU4Rx
k7tSgHExwy/pLsFl/ZM8mQTASjt65TfcBF8nxxCbqZvzWRKm4CUZ5h8zF4Oy
6tiLi4E7Mq5lE655or4fGXLleFlZOn/2vwT9sfmTys3QK6AZVSt2gw99LsEl
vCzugmeYr1N9cvIH0rk+6h1qRBXnzCJFjgEqHROjmgL3/CkNskzIPeouZweF
lWv2n7jIit4z8CUIA1OuE94/eZlfcMIQGAb+L8uUuRXFI52M5c1sYYr4pKux
rl/m4flojD6zbVcbsGGUVL/y762QlF66+mvAeJYpYFSO8XjsIAkhToDrowR9
Lbi7SUTeJoxo+zjgBd9wrlUIUGHA8uXvm8p5jvc5xhdatiK03wKf/CqzvSpx
qNnr9+/xVXTbSkUNzLQD8mwbI1l8YBp6FBX/oZcj61LQQrKT5qCQhykTrmui
mIMvEpNcScnvIwy9rPJS17qXq3zr4WtOknKmZGUflzK8fKmVkkzftoYIcsmA
oW93XDohKzJ8CfRVFND4UGkdFlvPcijkSHZT1sBCvuFToVy0S6+j/pYQQJ1V
OBE7AjKARaowYjnF2n0xpwh9L4ynzcRbY8+s6kypvs0gMf+GDOhNDIhsS/s4
IzQoEFsJDuL+eDk6EaJDEP3Pp4mVqZzRY+GmzbfBcCW14u/cB9e4MZ4I20Ec
8QYfP9ocwBFGkYfY1vb+EgjeSnpxBXVNrZorH1PPCIpAdtGNxy+1e0JJ+cWx
Hlg4jDan28wLCVHfJJNKTng87buwq8iaQGsUTLCjdG2NIrFNVzQ0iQ1Sdkcw
vldeFtBsSpkSdm1tZPkql+Qm2pkhl/YhUxjHw42ozMuypsZPP6/m5BeeQj7p
zKQh4GXHYp1+2cjWSBaKAYBxOiYZSaiiZQ8y1XiQkVAGT8VkIIoS+JfQ9m2T
O/jJbeqBZfwY90Eln7aC4RmymDBsWl3VpK4PRFp/Eael7TcmogMl8Ww8x6H7
pv4xJIYiA4fCRMPB44QKSNYDnxkZHrvD9fY5EkNcd4V+KmOQ1v6x+7+EYjWU
l0zyVuIprr/YN8YrFnq2M41nHLM9Um//+C1plGzDtwyLoqIhG2/pEl6bQl6a
cW+CmpjuCbTv7EhXmbozJI/VDSeellkFxaooaSCjQz6BpMItNTZJJdoOPKWd
aaiV/nIVj1EYwA76OW5uvDp3GLjwmkp/XH9/O3OmP8GY0uTBm9nGvKRqTXFi
j3r5rIbOgLtxYF2U5N/qkLbX/NT5jtPC8x8hi7JhnPf978iTBBMWDpU421mo
LEjskbdYiUw6rL6FBG9pvTHVUvI2LRtGzlkW4b9h/l72HVmTcVasBY/Hp+lw
g/K6A808Ybf+ggdS9nIsous8T1v0CXkPylu4IYWNw3UsYFQWNNj+msU9Wi8F
MbixjmsGRiyzosTs+8/SNdHDQsV5fxyaODD6HWOapAGGgmM2rLEVoa+ZehT2
mkXIR2O9TdAA1JcPUZwrmMw/KVZSPQVnqFIfOM7yL/TXAAImu1XAFAxwkT+N
G5EoGd9g2628FRfnM9TEo+ISo/1zTh6cbbr/m2pu2rzobysyA9zWs6hyCxHk
t8SCOY2/YXx5lJ4KzjEh2vZbcn5U2lHhQsn88B1ZcdYyv6op7Oe26uAcekD5
Muh02Y50jYr2P2IER/pnpBZJxo5LN+abmxhrHMo/H2x1q1tPOHVjU7KQYCl2
IFZPe2rsnImijT9gtfXuS4DhpmIk8inyHtHzRSf3mYzQWTPHyjn5EWO8NKy5
xT9YboeLQlmMHmZ/d+ZCj+CQyO7aepcVCOUvjj7hBrWhuVveIX5gDNy+6w0Z
73qErIbCVW7rLiquKNDROC5MOcKnDGM/gNPhZKVx4LcwAkoISJVGAWPwjIas
3rO7ZZuIpNx8Tdioj0eQXZDRsNrpQgctMiw/gBWwtYq5vKO69Y7O1U/WNq8y
VkLwtX6vTxPjjndwybNlPXgz4DifQkftVUgbKZUNmCdY/YfrXHu+dXxQZthT
cpQSPB5YVKqLdi4tk/YKtFC3yQL+03DXXfn0b9XJcfy9K4YIXEdHvBVLT61q
dpNECWcNa5TAvc5wNGKRwrCDd5n0btLf9yWyD+FqD2YbOOVh1KQ0CmLhsOmS
iJFJL/ATPVZaztWkLFpJ5rdSqlHYpIzOpT9e28E5IDP5LkdKYhb7Ijdqzhfd
PI3qD2TwKYWFgPvCT2AAq0WxQCAVRgpjcv4Dty3NbpDgpexVSZv18GGLunr7
9A/ZN7bMnGwG2vutKy2TsW2gLn2UHpV9ewjB7v6QQ/bN8wO+2EOkyQHVKWlU
CImYcMivW5AK/aK1C4e48/jgcbbSoh3FgMvArap/MlFxM413lTTUsGpi32+J
ad88z4gW9gSR9te8RTQvwdDogkUMl1nB7SVaeFtLrEPhwx4xar5aYWRsNElE
JnWgJuh2/Fscg49i8YIcda8pMB38zu4TBAu9/+9Pd86EQt0WmUVMH6s0X99q
a1ebHniZtG6PWvU5x6Hulnv4GoyTX599kWRdfqsbpeOOtr2ul5lvUi7c5Sjx
xJZP6TPnX5O59+wyzQaBuhfdNCPGiDaWw8Q5tw5BM3DGGalkApP+sy2kcsUQ
RtDAZn0g0tbc06QDPCdmT2BQ3N31AqWMm2bUYEHBWBAz1EiLBjOPrrXBALVd
21+emtmucEkvXqnVUA1HC4RjC8DPHrZrjfvSvB+XumQnaqVpXjvYQLKgIg+f
QBMuDF1N0QyVL6NPqevq+TTo94gPbisZx/nrJHIKnqHjV7KNdlyFL8m2CVUl
A9N1r5Ij/+Ytrmz6B2nphjnQz0YOkvJGqWV3ba778xax6VCqxMdBdLkwN8cJ
rhy/3PvJgPHoGOe1WxG3cOetatmlfeOQIYDqPotAsBIUGSR5vDk7TPAmH60F
rpGl0cLG+HDtitzUyco1IUmrpsAWKKUMMA3EdkDw6UM17/mMSklx5jMNmHWk
+hEbAS+MT0oUq7gTwx0Nzgu0mSVqoTJUpJQkB68QW58Q3P08ucnGXwOo3KKx
y1YIQgquKma/yyHFmTjM5w1Wxd2BYZlWX5CAV7cv8y3nIPlCu8HVrvqW5GZe
I8YP2crL6HXdyM0kQjVmBOFLrC83URN31+BeQr8i1DUxfjHMpz1LScd6Nuu2
NuLezRuz6NXvk7i55kwQCCH9yas7K41akdpIUNauxVG1it0FVlFEWyoQFZzA
7bWN1nYxsxwiCxd8W1n/9tOCQi8nCqY8TOPKuTld9VGh1//wj65ot1pLu1rI
ZXGvKBVBnV+TtOK2qlf4alQ19JuVBFH25YQSPPLKgILlbpQsldkG22z9hUBT
et1ldIyrEFHoZJ6qajQEapydIx/yWG6ew/OEdCIv6lAvMaLoIJjf3PZhspda
2gvn8wuegrAZg7Hfa79JN+e+7E1pF8I8L6jKj6bJWrjGWl+6edlxoXaCFLqO
miQIJp1HSO0rCd61AZPSkFPHOWL5jmQIXuyvo7TxjFJqMh9Uu9IHIicaL8+n
Zf9DgbPfnyWtb7u5rxfIH+IMkHwlLIRZ25F3ltwdinTsbn7dIz7jHZ6KBfnJ
4Y+2VK1u5OubKuTgPHIlra4Y+f/itDU759QyXZYEOs9EKcLC7peRM04B0sda
CpUzKhrFjrlvYyXI8TY7wXVyDreE8ZiHks4RLPaHEJtZQTdge29Nz5rr++PU
4M1Ho9bt6YN/pJVpjK0sxB4P+3oLX3C3BkJoou1uyK0+xBLpp+axHz1/sPAB
zpmUx7Cg3mdz2QAqLWqZ5qGpjDoRsmre+brO0NU1E2NbRR8TrpAnyawD/7/0
xlVoNHNey445KXQdTbk+mpC3MROjjhaDM/olYCSiefXpDdBr6GtfSGpXutVJ
k2ob091VDEPc4n7hBQDst1p5GrGWSpFf+QKgulP7ItW6PFHmFlOSUvcfNuL3
l+NkKQVSjdeSZ13ruYjlCkC/xcb85e6AbKDSZKhlwioDSLJfKmOObEvXQeLv
ViLisyqz2tC0NOFKZR5sDj31cWLsjrZTJ/xjEms9ieCUBlfuCDA1BesUF9O8
MoyVsIedb6G8sBk30eBtm867ntyRg30txonTxsf1djNv5/fNp0h6BPTZ2NBl
G20DrmRKhqC6ZAXOykP83MSROOLQFthWzLTi9jQ2yXS4BK1AT5x9Wmz/Gg1u
Vpv/nL5kX5dHNfwnkyeiicsyDWmD+T4BPMJN4WX3N7yxeLoRZe1HZwEq0/Fm
dFTn+YXNaAP0CCg5fWBXYddoUaULXQAQpbPlgH3OykOljFQwl/hAN6CEo0Kv
H5uInCSu4+6c2Yl6DPAHy4eFqzMfcah5u9m0+de9B3f6HZR2+0Q+5sZlisQ/
k1zy97E3+thvM/cfhR82HcGE3sLtVLchKgrPwpb1mnGLGVoeSa6ZsjJmexgM
Aej7Yzpf6SljoRRNWielpaXhIYdc7kBn+FmLrf/QaCnWgnR+8BhOflnk+zmf
Xs6ndoYB2xPgq6xyaCxEHU4Wl0CCdS6IFKgr78g9HZcxm6qfY16NLYmO1B1t
Qyjlybg/vaQ24rg3tz7MCWZerfhOZLgHNUyX8OM1GgycCM+yMkHHkArWaVQT
bV+PV/75OpzvoV9Yl7Gxvz1yXBesYZ9PICzXcfpphu2vTKfxDuZGYvtYCe/r
ROp2i9souvPqqV53DcQosSILUU1034A0biDzqOwV9lhsRypKMzddcbVhPrVK
+fRXAfwdvcn3AUSOQGC4uq1SwC3UqG+hHyXE4cYfQvVTdb+sIB2oI/EMUHbs
FhNI4JawWN5fjJG2uo1f+ihsUNcCV1kpi5shvqel1zBdO5iKTX06KxQ8nVxT
rkEn8bSX1nmViyF+QCxZRKh5QLi9Osy5s0buXKdJgeM4kdHbkjbRLOUX31yQ
VuSSbvQlXYZ02Mh4Z74f764of59wjtao5/eZHf1eo/47U/CIfcu8jwCZZASx
nEN1R+iYnoHWWonreg+9uvoA5j4NggI9cU2DtKytAdO/d5MLoPVV84DRws3H
jbD69QuusMWoQkSdRRrCM/qK23ySvfIW6MnnscnoeXjusu8yoOIvKCxE60VR
ypPJDST+cG/61t/Kl4rXhbeG+gzduEVR+4mRiupZ0DTVbXywc60cxcA2xtVe
aRLyXLsLDUOtGJyW3l2jRgHWC3JeEgESabNcYVOSt8FcEdKYNr4wsOkoojKf
ibAtCtG9IddCMs64HaP1Ay8c5hyjl6ZqNK0HP6063alCF8lEwjof7mF9C6Md
dezLVHL7n0hfZ9aIYP3jS8ZoQHbchWZw7Rc9iZ3DEnGzV2kUGc56JOHX1qv9
ZuMiP/l4s/bD98pFibSyxwK5lOFGMn6Dr05Il9ZGUneuNXo2TJgRBVm00LrF
NfI5GOvwIXqha27iZLHQvxReapcpY/7d4LPyIJuFFMybYH2zG+TFPrNS47lT
o1gvt/oIut4pSs2X2fh87U6S/nBa3ah6ph9xj+Zy1P/1AclcD9cbq8G2VHgt
Yeo3L/f/VQYh5MIRSNffdt6nUMktLq9aUGhLIjtpzt/r0rDhRlCmDYBTQhym
3jMah0uOeTimYUuJL/ue7EMK54TmyVyAOgXzW5I/r2MTbpHKFppXWz1nVwNX
qGDwFXYvAqLxw/jTs2GrdLaTeOEBgAAoG8BSEaF5tGYPL5n75P4JoO2TzrzU
QKANkymOTo60TSFmajSZa9+MQtwQypPTPrd6snMqKMb/daOC5yakq5i1+Uqy
0z0GvNxrGMltnZj1/JJXlXxwhVM13iQc11yPbqfb59qnFEpTzLx2fQoHsyNa
l56Z5kCqslPvPqr7nw+TTz5jeu79cioSekMkILSAWHt4Y8fm6AVA4iy/cNw7
lbD4pxUdJDEbDJp2dDJunlaWEJhuWpbSexc/y5Rb5QotCSrAAmsl2PQRB/Xg
ExxHRaBj/CFf0GDkZYLl3sEMUK0IUuDN7luSz3iVM9nzhna7FfoVqHPQIpdC
oom6c4asqoeixapaaXfzpQf/lSx6MQ222oNrQ34L+Ntgx50TkxNkj2bOZY/7
mwCdRyNCTXJESyBm+1qSrpF28e4zR1tEvTwPR423GTKar1xA3QWXpOmXqyjH
fUyZQO7wy6+Atbx5gGPMMi9/RA10CVhV+E7IS63cYjDw0eLTCVRllHUk9WOG
bbALgmbWW2T46ZMO3Gsj/1q5HHb6hiG5OHGQFScjUmFp0FTHmygjgYAa9xWB
Kssc+fWzJ9ZR9Qs+30OP1ZWhaldW4z/r5ybMJeajWCkKtGoOhOIDYWKSBGTi
Q3RWne1nPzK6MO46LyTbGfpGccNRIuDEi1nhCa8FzfglomlHPX1xiu0l7eij
T5abaGuT7JZXj9Le+CbpEb1i/HGsyobINfIm9GxhlvsHFmQLAVTmLBYpRNMf
V+/xaAWA0vsT03mQrkJ60atVwEu/vdyILvj5hm/+0lsSNFDYHihWE0Y5hrjj
YTeRayuekRRsbP9QppsJYxNNWnq9724bPB9ZDSt7vx0myZHfbeC2wh5t0ss4
zaBDxHbPp7Bbbgfg+cDzrAk70qYb84s7PhWlfLEIxI8Gz1qaXhTLOwaJpKdp
gvZNrlNrutCABPYXCp4czt/yLGGz9VYgVw3OOEebDhdYs7X+AFmaIyMdmcnZ
/ZLhTSoD8YzRcBrER7TDbOVOIxMWGfUJIiHFmuI/kkdolDLuTOnKb53+mboj
iSMZljEsMzMBR/+WaK7447sI4hllLE5ck24ObC4mmbfvNJR5sXwdjNJH4lO6
45rITm9uOil6x9ZYZOp5885hERJLI3iWe+tFI9vaSXu7UcogUrNyCRfS+bQR
VJtd67T90RX4A7eQgxLPD7v80Gg7L+pnxGR5Zk3rPATe92WnSWUOlqqUMiFu
chX5VWvNWCPXU21G5I6KAV+EF2mTYGRkl09U5b/1Nu+h2Y+O6n9nug8oqpae
4sfN1uZYm8H3s3sl4RVdx/dD0vuFrGG7RAVydfZkH+TocUBBTTWhNYSJERjH
BPSB7TWEqBQXQXkoLlu1ZqyN11k0T5F37U5Joy9PYwSwGdd7qxUJUkTVwlSo
SkBWWjSF6UzVtMS0fMoWVI0b0uYVIWfDpwnsbAdt7YAeLECQzcg+vSMpirjk
bCrTf71/awhqyI1aMgYcTbesnG3fioB4TGnaTx4CPgAPQo46V+ZhGzC1SU6D
zQ0IxNWLW4Jt9/aTHAM1CRG+qBEQygat1I5pHh6bXJmVFVWpZn2MRuWlzr2q
XAbKWFIPutBOGDiVf8Kmga+mBgtCRCJdTayavGXXMcNq3fEFRYloq7n0jOTx
JetbQHCWY3QYYnVIkI8u0Fs4AGPyj+t4nBL/MIP7xdhXAETfkd3Igox7dvyp
I75AC8RVN7rTwjU9lVdkR24b6x8GAbaEVXPDgs9hmjOFuhQT7zjTplP7xfHr
OukOlD2Q2IHtnNmm1ZMZXosNx6g5+rn9v7qPUBzNTw0/uwsZOiL+wPAqJufH
XpQQmbFEYl4/8f02mF31xDCzsynT0bDAlekN7XzXop9x1rBQbE+fpbH/SobU
q4aipXi2eqrXvAjSKKsNSUtE4PvbSXEN8cBUyLeShRaPBjKSjUDw0RGZdtxu
dD6mlpu9Gmhr9iJmMyZQf4IR635qfBAzOLVRrPYI52bx/O5QjgoKWhJzQCcY
ekynykgxxbAogRxfPNWrH1THJrUX4xfru4ZFI8ecITtgeD4rBWOTs3083RFt
i9aF8dXUgNnCln0ZRvjWO5eQKDMZZwUbsREMzWKCasUxcAsOZaB/SL0VWY0k
qksgl8k94GTIPpa1XYLvq0wTDTxGXP342VPrtyIuJgFSn2kF59/zdFGxeRGO
8pT22gbb5TcCFDJmWosbJVNPhcktYRnqbD7Yu0urNRHP1vsm/jLasbZMmybL
cmPC9hxG3FInu3JWBdnT8k4AWBzV/XBp3WmxIrFDx9a8ZaBbUfVfC2VHR6ro
S9q2rXEdrM5rGNgCvW6v3TOQbqnPBFfdkh7J9zK4+Z0FsNeVd0x+PqPZc5OX
kMSvNuMgwW1GC3Ed/DioKPRWsvyoK20IPQ0Tb4hXs0IHDyag4V2wVZD7hK9d
6R3wub9uwfMTyTsPbFYill6X5HME2RPzGrg8ZgXRvQnyyghhOxuCuNXm79vq
+a8FFxKIGFcJk6SYbNU+f80ROhunFki74/z1N8eQu8QAkePmKPx/WtlxLrs6
9MGi+5nrKI4RfTwT5jycIs2K1cJ8HjLay3liBK2FPVKZuRIAJaDg46OJZ/1j
AdRs9fLppsed1mXk0/9BFXaJmhdvfWN5rw/04I8BzvJUFYq6+5/KxURf/ZmZ
YsYVCeEXJ70Uvy3NFIhCvpYNTcQDcPqxriKTJznTRr2EoJaQuzLMnABX+cSy
EP3MNSKCrTERX4LX11OnOSXDNKHGsi4RFitS3XX/LNUSqOifBlW3Z/PsiLgh
GWl8nC/quDXdJjg6PxTpOsrnuIGCBwQsJPx9kwtRwaVT3n2t6Y71jlQmJohY
+3ZY7qEe6d46ZteO79hRDCP9GHGE8jesszGTeG7dsrmovsqMRNH4VSRckri7
HV1YkuQN7+63WG1qZxCECZ5G5iPMHmvzjQQOPqKUtImCyijK3BHkdEZIj6/n
RdrGlWn3FQ/gGwMdPeC3ZzgyfZ0c9v1oY/byDWoKaTnHzIYlg2zdfQ4pGSQH
vnl8EDp/Lbg1LVQpDtgKdvJt8XrXDQ+yUn0e4FcscH5effV1XRkCY2pTZCWo
vCkJ07vp/PTRUzN9zt0Skuvs1dbyfsg/BCvrd4S2oU977esrp/rkTGImX573
4GR3Irr5YDRJw4AGJhhwHPva0gpnKRbkdkLUcPk/jMom3f7T5dbQPJkYkwbV
fs7lzPLe1APrlnK1auvEeL9/Epr4mW/LPJoWNWE1FvcMfibvEZA035dKTQnS
R98KpUilRW21rrCvta+OR9yRWjNbHIujQR1xXbGX6Q8s+zwod1ryFToJhw9i
s5cxlhRT2iD9kPzDFtW9QNQ+9hfTDSV6Ko882dIW0o51+AQAwtqETseCCrnn
/Vxqij8wGKcVgrReogQ8mE3hRaLY4A0LC5BhGx/A19h3j4NeIwRXTOX1lTG6
F1gUVFI7H4Xbss21+39Y7sMa5AVEZPZMkZ9dCFS73xTdYl41vb/NapXDBMca
v/wfPmPLHmkIyaKerZPxH3BZx14Ca1qeH6FGbsLQ9xRHk2K4uM1pAVCSqX09
KXAcIJH/tO+d8GVRCIFXRG/zSU1L67S7IhT8n50wbruC0lbGpxFniSaL64Fs
y5TM5b8PICppTGKPcw1OVpD7gxdE30om5ZsSb/5wrdFjDTs9sfi27+QFNFba
8J3dkjL/asv+M+twkyC4X6EMverVcF9e6/5yScriLF26s+tNcA5JSVmXoATC
GDEpVpfI4I351JKcWcZD/6Tjm0orVdLyUpXPUQlx+VNUI0k8sf+o0hIW/Lcs
9r25bX5OduCk4J02VzHc/CrAZpc5xFxehG0myHZxmQIzz+hdHIRscrIrc86F
heCqy0FyK5y4I9OFolLbT4vnPUc5eK7AUkozH+1CTD2Gg/kt5pYa55ygmsLn
pykL6jiNeiWYDNF/R+wnf7yCgdJByvmZkhUXq5RJQhwjq2HM/1LuKEfMB9EZ
W2tE3DTfdIZXx5h4MQyUGMybx3G2L4jRbzBReybGZ3RoA0aAgLPvRyaiW4ik
yBqd0JTRZ+zuNkzqQgIw9TTrVGndvIPiGhSVPLqNJWALM8WhUsX8CWfYoDNJ
YrENsiQsHRQc0x7cUEviIKrXVdzsQWMv/CSvg+rJ4pOg/eedlwn3NS0nkFtG
TdBN1QVXFRLfDdS26ME3Kh9CYb2acnDu6oI6F4zkkw0EBufr40fHDXB/Om4q
WMILl7JZiwSBC0V0LXT/wflCF355sO7g6BkREiqGM9FT5mC6swYjOHkQvT/7
I+P9O8uMZYaQl6fbV6Y557OsHvPGPb99qVJrMnP+CZHEYKo8/4xjCQc+Jam+
HD7eZTm0DhvBk44Rv4lFX9pNwfARJ9bj7BJEwIxkfCDlyMQhaWwo9AW6vH6H
SUFwDEXlc2JrbnhlsTc55hq34HOM8xzRfGN4EiQWtbyoJ841XPG/LsRhVb0a
RufcLtT4dxTXDarZVN/BIwfpXZk1qc5awxyhxOmcT1J+9sHd9TL1AubMkp5u
4PZCyeVEqBUAFRP1A4ogwHaKOD+lpaHT+5iWX0aKgZuTc2U9OecLRL1EKRQ8
rijoSu+daawHGXUNG2XjPgn9ZDN4xPmiH01QPl0BQNU2tHLjZ3ZaHeWJ9N75
Sqt2Xc7Jbcq6cP1GQtsbvWXQG9JHsFwRk6tRnhiSA3XmsaXwwihOXo3xLtd6
EBEJJDKhlWvMInnnjzkduBJDEL6ZHPTVa5F0rblxaO4YHg2fOzBI+okXmZxY
YH6O2IwaX/RAVn3xwXDqGsBe9P0hiNw5istwFdVWHje8YKjELy0xCNomkrI2
uZKW6RP/QKcjRTFaXN4eML7YRR4HiUVqZZtIsSdxb6QaCWA0NouSPBXdiXoc
+WoZ5h3oLboiRiG9l3EftCC2WJ/pwS/VyFyx1KH/7TzrdwecJFmNXT0l56l9
bA8aL/o8Bd72DAHD7uqZjKsrCe7dTOIzHu0REnkod8RHG7ZeLX60BdCA0QFu
R3rb5JUeNO1BHwgoFXd5AcMEvmiDdJtNH67aNJZBYqOdzScVUoil+kYM8587
rcMnf2+/nsxVERBmhOXeHcQz9Fbe/9TMzfb+MAgzzvw2O+zcBN8MV5PiXWCO
UNh1ckS/3pTwPp4R0ia04hC8Kaq3fEyAN1sfmxgPEI3GF2lLxU9qrAgSF0PL
mvtnJAeRjQP5HhkERkwRrmsyUxOa7ee3b7O+TLtVk700HDAD4S96GoDp/DtL
dLlF3FOkbopCQMMBANhc8Cqxipf+IgGIw2fOvQGkc/MdsTNTYOsIf0fr2yES
FQRJM775OuMSnoIhDmQx3DMgI/JklJI5qWrm4I03onNFmqaiTK1FRHAosCx9
EP/lEI3w84aYP9AkUf8LiY7asd1w8sCBy13of6fgSoChr1V/LlJEms6WMS8N
jkQbAld5F1fvwpv/99RDqad+8inv6gM+EzuQd/07XiX7l7+COUX9q54NkUrk
fVPB5CM/xptH5kq4J5H9a4l6EZYhsVG+KpRrLTtAmUOisYzhd0LMd9AkMGL0
8dZ7GXdD8IdCnroDdvGsY386t8qAPrcim/XVqA/EonkaunhvJ8NqzT2FUA0l
DwLyFiN35CeuqaOaHB6tdFJhjMsIqOULritmCRLwJePfMD495uGQ40GCppLR
/KJjQ4s+RyaIm0mseuK4PfthUAXHBtvyHTzo/9h1OBrmbaOfJ08w2JPWtnQP
9v7QnkQ8nSg1MXCploX78fu2apzjT/t2t22nxYoWFXshj5JYU/yG93QHinW9
FZ7BkZpYaFHQhgMRVHTDQrAwU8cju+ywaS4LjnwA9zSg9CILvX+e0srh1zm4
DGDJH4cZka73e97jd16qLKaPmNY1CpWF68NpZZNsKohupyUEfKrIEwnngFBL
RXVYpCdC9T/WOqTP3fziQDG2nUPAnUeSO9W5EOhSQx4CwTLA/TWfkAdD/cWE
mRaHOFCYGnTJgrYYZ8WrUBn1mElSTD4Y0ojD6M4gk5yvpnucshu0QQJarDQf
Z5mCURl8qGuslyawxpL4U8xy5ZN96pwO5GiFzqh2GLFQMQqe5qY9oVVPYhI5
sO2iG8yTQX2SW/VOLkpj+iwvmcXTtuOfnxHLuU5Y3J20jW2PVlmLBk+ZunAV
G9zHmowA6nH+JKMT/nXVC58+QqrnnlNrL2V69lTtfXBcB4g6cSrJ9IPOPv+m
EOzV2DRhD6DMeNE87N4HGeMgiiwbScQXqxPYuJHmCtAwSIGW0kMSUGLcjhmB
E/9vLMlFHC6ET4BIJJHbj4jcL8ePpfUujhZ3PUuqsnuXAwAM13ubV436hNhx
IOo8reeToJvQUBsWLF0kByNQOJlQR7yZgdbYK127/q88xxtqBF7EaWWJMBth
854WoajLZ34DYee4ZqzjCVtqavFPgnp0uvcmsOpF0NqNRwrV+o6jawMOq7tR
woSK3KDSU+sn2CJ4uEqtI/MN286L3A2fZhlbf+njIBmOBIOahqg+EaPZ091M
AgSVlzoa4sH0tYkb9cQ/FCC5td6sgBSIcXKgpYEYOguOM5hzhHoa/7e92tHu
peTpXKVNYTKRRtMbMd201klcilRUYU7j9glLI40nE8HI0X14pTTzK0XK+dnp
aSg7lVzxTjhx9b6kQHh9d0DCtHjxtNfEXuu8JRn+mDckLa3Yi5ammgXFijh9
BU/XFz62knI7WWbzgGKVCuR63YuLoXAKMz0su6zI1m0CLB+06ElI9oU6oje/
Xs3qFXm2NncKEbu571maMKtM58JHX3OoENoDdOiKyRdp0DrtPKgSyImhdq3p
br/W7Eg5UhVLEaMrnFgMeSjDHFWXiGN1aHk32JutAqSiPPa4kFhbCcrfH0qa
pxPpF/du6x6k/c0XIj/+hhsoJHLr3f17ZP91NJARifsZSABqtusYSD7Z0GJT
+JH3yVPbZLHaSZNVGacRmSWY52YFaHm23rJiSvY4K+w+jNnhXAc0gtWYrhY8
w2NJq5YwhsFXKPMBNUYFfz0M3/JLRERFCP1eUXOQQ17b2xoAoJD7kWsDx2Dp
45ImYLhoAB3szXKCmFc2PvPX0TTBI1Pi4VEprRsc3CM28ELv+MuPdvuSE2Kc
9OR5VyaKtVWt3lx5MHMQVrVAI2u0WRtssYZosTdO+cTkgpnvo9xQjNl1qo/e
nzaHnK0fLjiRTDEpiytS1fRO+gn6YSDaH/rp+LCpNr7ZaNfJ/saCAJi4mPr6
FjP7dr4lCnBkoVkHO+CCHbCV9ebwKOWFh44zD+dZ/jk8fRqq4XSaLNI4YS/d
AOODWOWKJ/J771/wkNqcjh4HPclPrgz7OA1DKv3PUGgsRZdB2V1VDwdiFClg
oOmyFpSc8ifF6RGjKYWxBBK37c4YWJta59O4bVelpHv0uFqgGVlUzxGGstZi
BVjQQ4Du6cGFd2ZiOhLsmSbS58a3jI8KzCZNbFENHURiYAvQpG68SF8q3oo5
Cms/61Pyn0pzg3w2s2aqR0rbEznESt/FhOREpEoRaS+ywSAqlt6sNfOTHQJx
gmwvCR5+7JxqsQQ6gyD9KF5QtLPgKW4xXYxl59bo2vtsgixsAB9Y4Cpa0BMo
W9sVV87jueBwXtK/Usd+UFgk8PDQ3KoC0XbFR/tCNus1rVSZMR98ctFDhmYw
a+tFVItr9Wj+4wpDWyPnprOR8/O/UOz7CmRZ+GLFbzG+Mc0v3/NInqduQ6d3
Q+1/sc05Idz9izDQ47EBGBRXQanNIHhNGGVUBPpEgb/VkEpiZuIqSPIgFVKV
46NqABjQSxZp52chFSA/oZLVPqww8WeWEjW5IuzlWoXdwX1MEcfihxYLjjlD
6PK43eZdmMtJzVYp+vtkRUYpCTa/JnTOgZ4rgULGb8zW6z83XfnRaUjvsivj
W1pd3m2ADQUv2mMQGfEbo9G5Bc/pZerb3Li2SVoYTxy79HuzMtlKhoUXpAS9
wc3Hd+fgAs6vF4BCG8zTFDVAsaXil6hVHRxK6bNENVbobqjijmGs7H3xpL4W
KSUujJmU8QrmrkfQyjyu1YmuL4pS7oJtamjGRzWu85zhcNEBsDPEgHOq9IMz
s+EZAMhJPmeH32/x3DXIoA2DnXiQhCO3h3pCSLzJiYvM6VJHqiy7KB/P8Hzh
Ui1jv74twLnlZ3vraowEICiHSsUWA3mA/aWjZmkt8nmnY8kJmUrdyRUvx98u
dQvDnPCO3CyW8S4eQAasIdTq6LPuvH+dWRUDqyY20N03gin8V2fWlLudUQfV
g4wvd+UL03K4udsqxEK+G2nblNx6f1G3DlHu9mucn85WmI/k6oBkVHMQ6zAd
Qwvf+s6v2IeYRq1oyAe0VgwX3EF3+PtaIS9OHNJciYORExnBeaxJZKI6SONj
mcPzZWe+VsA4sXHMx1ZCxGP6xpakahYfnooogBimdC0RwHNncGBJ/FkC5Nhj
5G4NeoaYsSKHR39Qjftih6HoYCAYxxszZgrOwDS1Rxse+ofq+BvclZIiBYmw
RUqcSvb9S9KT8dEsKUJumg66yrzi3jLWhOfglUGfih5HogWiYCnUW/GZjM0t
7jHwFooqUqC+XZOvBq9aiAGkHuS2P7IVbVdU6wdnFA0hEf48CyRp8NCvK7As
uqHvHdx2K+MUG363eKwhL+UgTKRDDq/RfSGzWHNd5XU5J6YyaMcv+xTBqKHU
Yj4ozS3ljSs0ANlE4R5/TsGXqtEt79t6n0Itf1sSSzB64cqiiRrLchLYHTux
x2BYVe/XVn8BlnGeQzr5bwlGjL2pJqi/yO/wWqWPV26R2yUXxy+5asuXOkNG
BkVMNaVToiDjVXB/ZAhiWzTh4DqqkVcn4S8Gs6UEXC6jpew4hEpU5vrrFHn4
B2KbFYMm5ZJuNxhr4aPDvvgWOL6X/xCTyt+kcbdwwr3bm2gzb5Wh/efNuY7u
9iT4+4cv0dyomO58x1mD+pmk151mIbVwwY6D3PWNo5zZ3F5S27r9PGxNOjK7
+JNo+KuEyFQErZ7YMpiEBhkUcnrT0cccOXKMG4iQNvqeI4lNn81i2fMbZ8UG
ShtyVRs3QU73R6D3G35auf9DI2KFXO8ja/y+tLu5kGWQ7mzBYTw/BajMHlO3
WPOLGaQRShGaLYAUOHtj3o199+vhZn4ipbsJnAQNg5VaWYW0GbGkoiE9vumf
HSoTuSkGziQRRS5taLAJB+gq6bR0y3ZtHbVG9P85cqMOTImhqfU8AxC786aV
rxPmCMIdrwVR0sftWavebbix8sMmtsfQdBdLEs42DUc46urcs45pw4TFlCTi
XcOZTnIvAmXq87KZufmzVgEueYXQpyboOACl5v2OpHmH4DLClnlGj1RAb9HK
k9VTNGx1JBDWNX7ikC+T3+8APj16ne5pQGrUhTmdPTnCzSpwahjIlc1dBrHG
KfbRgx77M84H8FbMHGvRPaIcR3VvOe5XMjqTHz2z7/fTVv3319rFZ6ykQ9Gl
XHhgPsGwSyrQzmbCKUiW/FzvzZg2VxyeQWjFi04u0TE5JHQTA7Sigsd2iw62
mpXGp1he/4oUTgBMxNrHcLariWFTaXSkJXnh3VMhHg/P2P9daJnpq7E89p0a
ngqBPlm8oSod1OWp9hM6rMdV/c09KjZr5GgDkGAAB0i8vJDmoqIQNsuhpXj/
W5K6j8V8s9Y4kl3axwUjLvJ41hxuVYMvduv4N0t5WrrpG4G8PgB74tfdm7yS
8AGqIaO5eduTjxuzwDUSrKFivoSfLFVC5o7x0DYwZ0MMJLKpUOVvkd0LA/Ma
HYA1VOa9HbdLhz3rL6oeZh25YS2tY2SPgKSe2uWxIHHcsBAdvYkQYLEgthAn
OROzxLWyIaTWfICQFiSmpA1dmbua0qRh95L95d0ncYTIVYz6cHbSiweREZiI
p5Lq1kyju4KgI0KvdLTdtHFEEVScoFBbCSXGUOI/d0R/r7eFFHstHHBtLhCw
3KB9BCNhOKyCmc8c1Ry3TNPo2aXY0KEqJmHqfN1x8BigYhusrbdikYTPFhFI
9rRN+AKWCEBoQnT9JGY3Oe/aOy6dO+IcgN7pwj0RlYCHR0CukcHshAJS0qgr
m2UWeC5okss01jPm5P4FkYuVP1vyALpmL2EKPRpiK4A4mW8XgGrlCVAXpWBa
t8t8QGMf1yT1xfv6L1xoArG3P7jmh/vO/QIB/TYqMBocphq7cUt10UVia0mF
hVEfw+CG7U1yZ5PzVXcbR06dP91QKA1s6G6rZ6mrD4WMv/1A7zBC1+9B648Q
ULSStTSYt8x+BvPss6ueSg96QwQHIlpNUtNbon38hwbnO65hsNWH3O+B6n75
zvN3rcFGKfZa4X1ptFHF5qiqhhCBgqDRWAR4XPZcAAxza6rSnYm2tR1+d7sQ
Nw9nuwujDBv0zJi/UejHz6VANmQyGbx0uyibGnE1Nj4J0HUqLjGcsLdkODvu
Z+h2/fUcGp7Q5WWJ7AvdWftUFhBX3Jx+ylHkY2BMXZoywGuDc0RjzCHDLY3t
qDqE+9OVU/tEH1TEwVhIqqBZucG4s+qCr+AL/EDMq6pfyjEx6JkMB+qprFRk
HESwQHLAYJ/MyY1rWGw2S2OZDUT8cNvfG8i2E7dMcdwWuZh1BcJqn6XCrFsm
m2GKKuEPBmuTlp0BUATm4oKqfiZvrl8lMSJBpFrPD9TTeErA3RAUsbwYXKy/
AyZTUQH6f4VFzyZW5fDOcURdCdlRw3R30wSFbWcaExhhYovfP6hVZtpPkMNv
GiE0ahWzROdfVq4OOx8sSe3ZlWXBTGo9AiYpCkscyQWAzpy27/7Tcbwfll+2
mIi6eFJbfVparIMGo6TigM6gVXoQ6L8+Hav2zLomAyxzqXhnwjBfsICtDOtU
BDkWYXFPpKEByZd+PCuQl4MXID51LvYGrDv4r9zXpu7Gu7gxPpfJYfOFvdm2
2EDp6LnRQ7+5pPebCkOwoJwpOREyFIac0GZMTqgiw482X8c+ZRV80m1KdFwi
qzMJuwaI7MikVgnwfxgbgwbMHMLGHRaX77otXfMkJtAHP5FLrSpwp+RjmviN
jAVUihQEigNQxdgEqjco5E4ZzUjNmBYsPYJ7AtyH9x9hvdZv6wGB6IfBxixP
r110As6hjOFVkaepY8c/OAnctgGkTlmMEBQqqUt6gLCk9Fb+w0ojz00P7Ul+
yKgD6IGwZbM9vhDmSqGw5WxQord7O+g0tFFHt/ZQeBYmawzmCkVrHJquvIcu
xN/baT3zxxn02+7K9ZDRyl0//mQQtMlL/VDA6o+tntLlSsbpwucLl+NCZ1A8
RWgM2QKMr2WNI6/41AuA0zIsl2oGobOGyUY3ezPucJgCzm8NEF4djTt9KpEE
JZN+df6VOIlUnstW4FzLjr94e9vCkiZcyfBIX4DtlRDgRE7QIiO9CYYITehM
pEznim4z9y9A5qu+73791YeocxX+zc3jvlOaF3oitLJS6bAlmlFy/rzvK5p2
zF4hmz6k9qV4BfxERdnmfADkplTt4AKJa9rZg2BrvoeLf1cKhkTQaTSZHpXW
RnijL3xB35GlFrjNQiaTSBeI1n3Fc7M5o4uHB4FR244ZLBQcXzDI9l4zrq9x
0pFopojsrRpgQJmG3SP9n85EhcxPeTsZL6r6Na7k463wHj/T0PU0/z0pWaru
5i2BimvQZpZcmMQ5s3X5YgaBfczj+UAp+oYP45NvGmfhgvhy6+FShGc5nKEO
AxVwgBdRFXz/IpYRl2urHUDtNpB9d8lkx0fndbDVXyj09IKLOdsSeKIsovte
1JKOuqocluKKAwJNJRLu97SI6cG4ddFqNUcTs+Hg95eKohgBJoqFbb78yZf0
ACahDgIztGU1cOWib3Jd1sEnzq5pjQguitlzqTSqNHBrGyVyHjzOhsstAv5x
nBqHOJcxmXY9HBUrIk71WlTBnXbvmYtavKRwU+DAYiOkFaII3sFK8ZunInIm
qOU500etuBgeZX+ThkPxjoygtTU21VLeic7Y0ktKPcuYpgLhQtk1eXJXQO6/
HG9r+vtEO64UvwEK67nBdBxRNeHkzllxV5DvI0jP55gAi//iZ43MsAEoUEI+
DcOnZfo3qeQRgBYYBnp+jMFhfdwVY04byCMONZ3Nh5KaLmFh0FBonWYUwMPf
CIlRtxHt6iuAEBRrWVy1zsvFo0bteeXJr5BElLyztM5PHgXk1I+hxwfuH2rZ
DUB6XjhYIbNj+7D6Vl6Zx3EzA40h1E8HnHMOvjKaUyew45RxIXs/tL0MNITs
aGBz40zHg+gx0+MdIGnmfcskbXBBvfZPYIZrNP0196vocthFNZuBmzbE3vOS
pGs+itowA4Uuur8S6UrALjhNzo3UK/ECD1AXkbE0XGgTtgv6n0q116Bvq4Ik
pByqDkJPrpccMmms0PON6Qm0V4HHDkokkvxiSII2JBJJXATjY2g85bBmGUts
s+g6BUV/fvGqFKmxW17lGOxH7IHtaAT3cAU4Ru1a8pHPdjI2QijsG80B3wJS
GhVLrrK4bXp0fygKlaDeCh6h92rlLOujTQ8tFI3P6r/r8d9+UVkwKoyUcmGH
j3V8BY0CKURtPMxVuKpXe7GC9kI5PxPopllkoXFjJ2V+xgh8Tme8GwOPB3y1
RytrnmNhDBTp+MP5wGTRcCEJO4oaQgUTZYtAgFQ/5Po63YoULtC3vSYC05EZ
seX8h3Tz1Oi/TnpnSB1iXlnfO0yy0UQYhGYM4/lycbPbvTQMlJijqRgTv3C7
jtv6wH6NZ/aT3Q0gKGzQ3UjpHVAqXFCD8L51ux7h7dCKCXmws5MWcj+hCDOw
JDqXmoY1grYhwDut9Dy6xnuD1r3pbaYPBSv0J8OOog/Co3jr5g5EEL7BrWP2
QNDJ0S8N6L4JHtes/yqxbWd6bFVf9m7DWyyDOQX/z2K4XvCXBK7tT4me7Gfb
3FRnuiggyA/NDmPfVM5n3/89BcOMS8pKVkLCLyCzckE2D5l8DWc+M4p/+S0H
YI2/8wmpT4HawKAR6+D2AqH+mWMntog3bMIu8pokXvSErJj9TPuNcelvy6Tl
l6mkrv4Ve0LpSkNOjgKCT/UK4+ifsIjatltpe4/mREv3KAl20E+/xFbOatYX
ga5WS1lphw3NLQ46VZcYI7aOiLcZgtZyCWv3rPupsQrp2klbSjk2tXI8fUNT
GDtNDTqQ8VRliTSna7asBZUYu1AXWCbMXXV1T50VI82O1QQh56D5AWqBcwFO
SaorSqirGyVwPcB+QZ7Xz8Sd2Dj2sOkDcF+Dk3fDF5ujbnVytaqAjfhdEx/s
vzz8mI1Rvx/gS+/kUtQ+KFR5qO0Q4malrpKyGPeatl9bp1PpkdtulyZLMfgf
RYQBZfp2AttPbvz64ISZUcFctwHWCs4Aykz8KjsGSoXYbadDEhhRKdyDPRmP
mjLD03/66g+XaIus+oDf/X1PsfzL4TIofdJhEyESvU5f7puu0dShyjQBGO0Q
xsVJyYHIZiqItIcfqGYuXX/g94GAd4yJvVY05M0ryS+es9ijKiLb8FK6mXq5
cRXLsD3rX8Q22LWJw0wqUYgm4yUZDJoNWWGzxhosCKfj3/pbjSby82/A9a77
jpLhKj52mVefqh5ATCNd4F/807J82F8QYoG7LVVMi38W3vqGaf2P1Uj+8bpX
bxDn2ucszoI3uAsWi/tXHtE4XlhM65jYrFzapnYazXGsQHjikFkEnK4tmalV
i6F1uAfHSS+v5Ktza9UP4FUc/XtsTjSGhHKMtuNaZUkTodSek0NjpkCN6WuJ
5ROaPr4Vk0qXI2R+tMLOvYdN384csdz1D4GKhrSRWujXXT9LIAuNxSxxTvJy
C8l9DDAhAAZ6z5XTgie87SWV9vagX630sv5CY/jsOIwkfRsIyUJRWxxKgblB
sH4WrAFpj6xgf6YWpLRlRKBWnkLzdFnq8D/USV4RxEaR/dZxdCMsf92wZ7B8
F9hKWFo1NwgHtinV8iruzyKss3geiKFVmbbtkGEpEwYL3Wqrdd9LF65yE5YK
Er7j4MHJZKeH/aUnfzddBZ0iRf9W7vo5Rc9D/SmUlW1FQJAa27M/J78X7rHY
WrYE5Qht5wXRhG1gvnD8WAhhbkl5q6m0CM2Lqg1Yhk4HHAztuVmINO5cTEeQ
t5whGM19dkMktFInwabzzj8Oc+uZpXq0SaVvAyunabaRTT2BkluZpym9fkTH
H9Igs5muRJtdAp3ySCrCf957GHL3uZWSXXwaOsiHFmI5U9Fopxhne130uo2T
LI2hvDM9ySn041ztwtMzT/WANCalyOeT95OnoJ7JzP/PiueMrMlmhiwwhEVd
FeCPfZd4PPyOi97cK/1k0cmKrgtP/62dfGumI8CIP9DlSXPEf8G6A1WOtNoN
cDrdrCRSaN8Tma7pZmeHYeQ8q54/BOrseQcR9h7zACjMB7w4HzIG1hu8U0Gk
23s/zTolSCEiiH9qH1aST5Cnbys+RBaWwLGEg9Z8Y/QgZ0vRUHM0dIzsRxZ1
3X49K5JbdAqcS230LizSFe122eJpZzoH3o5BVY51SK+C7Lgf4z+qsDVqxL4C
r170OECQPItN7bOBbymD6y+AnXA1hd/dGbRe7Ow2L0tSLMk9wSAYf09oeUyv
0ySDq/a+NGQDEMBd3j9UcSxw7ds1lvswXGVYxNZThHukAxeUoAtGie+l2n+4
q+6VXAJPNHwXMaxj8zV1GVBbttgpxAH+Smy1oICXUvsOPXJ2iAjhj/XEJqCJ
lXUlwgGzqrKuKTnbO7fQ51pubGIGF4unKqtrRbSHmgscqbO2dFsptTOQDgLa
5YCX+OidqPwFnWhspR6v64QQhmJd9shDFNe2SgBcji+v59LAQqgdrmNOB7ke
KNJFaahon05eQ8WEM1rt8w+J0OlvHCBjJ/zQpSlaK+nrafziKbPf21ltJf6x
ll6IJu3R22VVoxO/nfgK/xiCGL3jT2/BVA6F5Gi6GkmmtZLpr2rK+2Iw0qmS
0+8ehewvruU7RzgJFaGjsbrxDqzzwCHn6BKRQSgqEazRrFMAqHunVh3MCdC0
ZPbBK3pGlhwOv8/QTv27UJXt7tyaZLnxJJju5f71WKFsS2QLaDo+5bmo6CfG
niZURvzOhzGoI9nlP49qUFGyT6UTBkS0q0RgFuIekUK6ruHGeAPADJgvo5XD
NyuZMk9+Mfhw5vC01gEkIzUNXOvmux/ML5ugqfBXcHG1tVbbtZKdQEVX0q6w
BC4rjS40c7d7uvePHetcYiE+E9UVgI4d6fQj2NuiMNBhkkL3cmcuwczUn7vo
hi2digOKQSkc2uOIYegTaNa53+PYnPGmQemL7ImArzPew1GgVE+HWcazdN6y
N6TAjFie+2lH9eRprr1myvnVJu++HxHcVtFFvOGF2tcor6RNgEAM1vzo0J0M
5iJQP12VDYXuHFrc8Ck9huIb4c2NulLuhEmAwrXvr9sgXJSUrknib1jaAfgG
uGe/odpTubLEu6BlxJfq//06h7BU8c44U9FpyXQ1muclQsQcwlzWAEjUpC1Z
0fMbk7A2jTt/wpH/fACtojsrVpMHN+vWdgDem3o/yIK4nEpDtMwmQaOuvzh6
uxzGw08NpehidSvu1gqdcDS//s2eH0NEbfq7TZ9RWrcRVxNCQaJQEIaq2ELX
JU3Ohs6ENjRlA62rOIpm+Vv5bCjpIyh5e/tx7DumbTgGwH/lsD2zypIjxNH8
6WSrkKd7tliMdDKitV1qg2biKKKS5olmM03bcLSZ3KX+f4NSUYfMHm4I8Zgd
vCx+9WAgeCNw/fH1S4jawqk8a0fUAneX6Kq7x5utmaEpih0OHpcjG8xcKY/q
NhcwvHPUatwH1zX7bc+EEokLdld712QHSVp6P2vwBOQwCGcq3+g+X3dH77wb
ykZNgYln5k6SS7T2f4rscwC76DmbzfQ/oMxXoY6MvuuUYGfHXL8geFIfohLO
F7Blbk9S8gYqliaQ9fbR1lYYNeV2AkAWNw76Uy4yWWwqmZkDjgQZLYQtLpbN
yT2Embx3hVrjnfj4AdwLsVjr5aWpVT2e+t10cL8ePSXDqcFga8TavwbM57nT
c5eL5H/FToLl5F/99DnX3Ztz5oM4vv5yNTEGPIk2FqIOnvsiUOlFHK9JDMBz
vE56Ak+KTMDpyHMajNPSkGs8g54jUkgWdR+bgaKKJFG+K4SuZ6MZSkCvchzs
+6drp+dnoUoQoCZneRdHxbgvxzHp8s7oAr1SeW34c89Ue7N0AhTUsaoIH4jT
H9RT9n6axU/2PDNS4KVhderV4XiWOy/mc7uueXdYE2sd8pdUopI6Kn2W/r6R
901VjMsY9kTC37xS3db87Leq5E3zbQui9WZTsmCj01erEx5Jr6pehHNMYsFk
baWhnsqI7s6tZSk6e98x3zYOI28tgPyP7nmvC1PJ7rVso/CnF6yGoruiFdLW
FyEC4Cm62PE673nWwELuk1xGME3m8rxUhA6foqeh5zksj88/rA97bIXTx0W/
d3gkVUyCxyVRce0CJhXg7Gg2rOrF2aebxj2NtMP4Xpojb1XoM/7Zu189WMNu
b/iK7l4+Hmop2yEUDGFVndVrXLsryQOi7DLj4yWeheyN1qX4/yaU8er+fadG
LyX2TG8VOd7IopJTgU97Kqs0tKSYoHXdMVkDXtGBpM8UVQtXas97o2AT40Mz
YNWddgzVCc/2XGg3MmD2v8hT4THKDhSxKa+ydggQg/SGLNGPd7DRvl2Dt7aa
G9g6KKw2iKhd+cDFvt1yPxob0gYsiGfdZoGBAPIByCJt5nWrJh5u7J17iEgG
UTLsQZDK+gCyJkiVxvj60xD1oe7ZkKFiBTThizkGpZE8fNeJVxiWMGr5iWHO
g4rEaAOkqDOTpopu5CXx7/NjjDkoZXrb2hTkaof7HMXRVJUql1i+B4N9XvDN
P+nlCMs+qn1QTztz1mKNWkYXwrMY6jSbzjnzDMSyILmp2E5TK+rgdGCbGsxe
4Nlq+7p4pbZ6XRuhkmCp477998kX58Xpqr63pS1O5BCS683rq4JkolKY0CkM
gkUHMpJLejV2v19X9/GIgtLM5jNv5FDle/6nVSYW/i8iad+W5Nz2ecw4OZOr
v8NdAlF0mL8XjL7HhyqELgVyqiShgboIgXnaF6A/j4jR/cjyUDY0F8IwEYjH
WqJ+XotnJJtsFm2dWfV0ozF3fsBVuCssw7vi0VyCEELKn6oG8pjxVBxzv89C
AHprm8ZU3+j5ZFawgpk/dkkYWe1JrvOJmZFhrKpH9s1yegFeBERA1AwMDN+w
cAJM3ObONcoaVZyZbgIGrcxNA7ypOfW7Uoz+3fqZc3AsNRMAp74A8WcHKDhD
ahEx6xg7Jl0L+fK7U3BQFkI7IlOzJw9hhFI7igPtVM7EUuQekjsBlq4jPq/X
iAZNgiwtyuCpEuEnqWdUHK1NCFslT/EQwm/KzXI+0STFI7bPmf1KuDhmp6Be
zgmHkaahLcnB82FdLhHj1H+YlnlvMnGcQLXrBLTD+vFEVNW5k8N9udpbS23F
lHGjYnqtOB/PjMwiEyMOWZ6QFlOH5T2J1oFwdwEyT8VE2DTidlVIMmwzdwtg
qSHRRLLhxzo3ezr/l+GtnAtbZMYbhAszLFjx594hS2IG7Dragk1HmbTCr/1D
ag1pK+FgwsRLw6dqwHej0p40VCr9EzbJpU333n8rOPMfS6txtuY02LuIwOJn
pvONyZGuqoJzb41oOqTqx/D5YP+3N4gaWLJz9FcH4+xYMUnYeTqyEG/9KD35
6TYwLeqBprswewwOjHTRoL7YPmb9swfYP9Yif37ICDHXFpwaVenDH1BazZrt
7qOnaUJPA9kR8ToGDwPXCwxgv4tRge1CMzehtQN+oQVkcAuwfRtNDllY6SaC
KXxw+uWH6ZkxE2vPQSTqewbOFyNKJC3LFtO8mNWlzmEAuT+4sbyjySZyKdde
yEjQVvIBfGqvQtxcu8iU4+Zs1EBnHZKp4yo+SN/VPkCBfnwP7V6I2pBZaZrZ
No90UvLrpJyIvewWd2Ic9mr7stTtdf3Sa4QwgzIyL+MJ31ySd2XNP2XJYNuM
5waYOmDGGR6HdsbLnwgRGHnN4g3xYO4k38nRWg6sXDpL2ClYkl2750Waz9PH
CUZNGpeUH6A6yzkQM7j34qASMX8gjipAGC3J+MSpQQYUi7HaAMbloGWnG7NJ
s0azooRebvKTWG1HiX1ci3dkCL/w1nfhHBTimY1QNSAcJ4c3/BgI18sh5SNX
TCsE36rBZd/detnXNk6H2q5rxAMwQZSLilXB0GkKjh1wsVhwgVrQyw8ynH9t
qHJkRMtFxuU8a3MGivrHtZ/XSyUYqf5dNmbJ2kb9EBej4yaxe5D76I7T9xT1
LItAKkfLoWuNtHSL0p11kR58b03pYxdCRWmw+xcDDFgnsY63vLlEAEwpaMjs
XaXZNR35vwsij5CG0oPfI8rslbsZoU1NAtU+SNq5CPxkDASGET9vrdm8A0RO
QIRmA41EoY+A+1cPHdTJFMzdkfSXKvE/9iJYFZ0iJGDQg5CWS5ko3llAJwjz
wiyq7wVhMrFZdwgqk/sqjJl7KxGt9kyTd0sV5PTn4Y9yApuu0zay9/xX7jzg
7Dh8Xcaeaouo2b83NQ+qq2R6BYKRnUMe01N4d+5LcX4rP/lUk1AtxAGUUVV0
nGIGRLCoSQ/wmrAj0Bb4S0DP87qihdICWwD+BR+YGHvmudGX9CspR2RjaYDC
Xa89GctiU+jNoxGR2/+00/gnPmpvZk6VRl/eNJ7mCOWozPLhKxWk7LF0x5oy
r+O8Hmxoio/4N2TyOkT32lQHyebObVWAK2WOOrUu0kbc5R6TFgdO+iedQUlq
O663iVcqr1hqijEZDlMmqpvvTso6QmRDxS5nEDrOmeNsbhsVV+3+5b+LEZxj
cNYjLixI0Uype8/zwC5T8EQ3IoEkUVKbcIfMYCwY3c8uERZRa2RIstYfkXil
w4L73HKfcMU/zWRESz8yPGuMz5jdMicut58e4KQRlf+UTzhFpipgbi5Xg3Dl
3r7CaVlTToIfgz7YrNR2zalRg8Gdr63A6lHXKS69M1cYYEiQuN+Tbuc19WMh
tsd5guMIziu7ckWQXj49iEkMG3gDOLI21olXXMK1SXppqt/56hAK7UHv7d4c
QyKOzzcNlTkDVAD7Z9AAslBoCs6iRD7D0zwT1r3M5D5a65pafhoDV8Tofi9u
7ON/khh77eD2bEG0DRD3OsM55TzCKvSTZby5kJh5M1eM+9+RIhDfiRH9H9hA
hD8tUgwgamScbGB+GCH9kyBsh6T90i6gKkJxMu7ju+dGI2/5K8ZEP2znlAt1
y+GQkPdmHTeP5MpfvnMljeZzeCrA3F6rHt5ui8lfxoyR8+lu9QDDMIiqbRqz
GDwG5sfbq20f1ZFMMTIyqzrsj9lNeLOqepJ4+KPv48yAj3Q8UGI3xYPRrIH/
zI80WgVgbDk5VMKUo/1AHlgqHpFkP1S4LL+jXgYChZ+hhrxO3aJDF1gGVB8x
oP2IBnL/aC47UswC/ACkLtrm6E9zIv52NSI8/+p9etKSZXqNG634g3DvboN3
7RG4ikEkKtBz41bsZzVjNimgoGjZcCUbpD27whbmJ9bBvmlDYfNTPB1spOj+
lwtSvI8L7/Dx1Lyph1W2zRVRqz/qztjsjFFfO0IKHnZH/Bpf21hygzTbdKhB
DeIeF9HQMugReRRRH67poUNFT0EhRz41JK9RisaeI9fE+69yx8VAU4RzXi2K
5ahsMMBVFo4vXkwDwaGa7p1rKkQSh5eScbp8zslZrwNGWcDqTc+x38guSHwP
gtDphT+00kTObOAyZ793uaHfpASuSoOPHeETmwY4XA15mq2r41bLwWOvMeUq
//HvAh9/lfUAQZGf3RLgc1s1FymJz5TOYB+zU7aT9lAT9Q71dFh/3Ih7vhXP
Gv1AVXbdNo5guRJ05N+RNfc1F9OGSvGw5lUohByavDA9OE8wDqpzK0LMZjmC
N19lGRCt0oFIP6iXLoRHxjrh/c6yPPuNF4IspDb1xipf+BIDYHC8n5qiN56B
PJdLXuEY2kGXX43bU0Z/Rpuo+4H9n3u9LUJNpoZrtG48lEzr+VOUtLyk49oW
/HrJgPcY5OV4K26hGMtSoyj3j/K1jILnTuVTUC486yW1zvTy4s6Spcu1gogs
iQLVVwsNxldP9jqnMJsqcCfTTSkVGLSnwkITExTeyjvfT6xAbSKyxFSVNSfe
brZaqTtnxEij+Hr+pfXNvRGKWKl+/ZlFEw384uBH5QDR5w1FSaSdfg0AXUMl
jDkfjQgOgX2ZSDN9G2so2asj1NgbRrK2aXlxqohTSv9uJ67WOB1kG66gAnxI
5TCAMrdeY19PZWUAosrkEOBWF37t6cV2CSlnCC9dCX9qJW76yDA1kpRMtPOG
jEOXNIj85YbZh3K9bGsI5OQCkark2stkaSKxucf2dQaHM57mLFLyNAvxKP2L
+waRgap7b4s/TaYYl5wGC0dM5S+N9IGxx6qx1D7+DEaidXRvEN8DRqORlGzy
l91yWCdr9rEfi1r40ceVuVxc0tFlKHMSUICVkeGKjUzfLA8GM9U20h4qzmXz
/+jDm0BEGkvIoqE+QitZT/PEaYe2APDYLUya/k7ausGm/Gv0Rr8hj9uZgTR8
3sFUhvxIrx1RZ6gpYz0VrwXWV8V6lrPF6oL0wW+GDy+xqIUZXSphF55QbxJX
I+AXinf4Izwi5xmBWQx7dNLAGm8wZp5KnQSlIwLoKn9idfOYFIAlotXUm9Yu
AGUsxm9XLmxtCmqRgthKU8p/gjs9y9toX1CGE9/hR0+3kr2bImmsBXRUaWpA
ihFYKMGiHwOSdpUBb+XMurJO+gumc8a3bh4ldlBvltimBwO/AbYxMDAWdkL5
A6NqVh389EmrjczhcLU2Rsn7yIvQuv0W2qx3ItIcmb7b3b4hra/n0WfA59uX
sd+tXhLnktMkWWJNLUA8x+h5/rKqLjJgXAlVN8hWhodt8PBPKUSeyz2xKZTI
evE2PDkYj5KJFPal15hNkFgQjB2QM9Ot35S3riOu6Fvo16dUjLfTdMY1EnoT
RHgbOWAkOK4itxKCOKDbnh3lRyxLvuWsIExdT5qqHcgBSMUpi+WLDNMbYMB+
aFF0HmEVehW5GOhxDK+fGGHnPcSfVz8BoRkdYrg6n3QGczwuLYILWM82+vRZ
uXEtUhUbjgiR4O0+jdm5IyC0S7LSzDh0+SzlTAXig1c2tZ/UCs5DVzWvZjSY
lBAX2t3rBw3JePgTV0LYjxCDoppvETvVEKXSiCS1zaDVhowoxJWT9SOmTvQ/
QSa1t6p6j2+a4nwWCimge6+HVTQydToRrJGCA7KW55bUEIGQ4v3qx0DG2WHQ
zjCcGKtUnYaMXO9MoaM6AqaKtiZF2qxhVPzaSsn+vkBej/0u/QLg7G10Bqxw
nB0WPJRzIz8lApT6SVwB2YbkXdT/a7LvhX0AbltzpyI5aNvD27uA+6QZo/FP
VYJJ14JPer4zyIiFeNkMDYAzoMUxDOZDfXAhQYD0c82VqHSQWj76nYWXfYTZ
TArFtkOCGviVsU0H52rweQGYNi4ZYOmPrcc8teB9Q7DdUgy2yQ7ZOcp8Rd9L
aIjPPIvKNTrK1eotSvvgUH1HS85vznECPVfXrWwpyv8nPQGLH9iRIsKCKvGF
xfEvJ/rf4c1+cO90itzQfZ5PdydkzVAyOf6mzojuN9MmJc6IF+J84XssWFPJ
gzmYUsC8BOa/AizcMoaPZyQLchgn7PB6sN84CxdtibETwCIUVDwYV8bgwzac
IihvVU8XMMzwOrWtAh+qvLVx+D+hYEKxl7zzzVE72rdtvnnVBmfG0ekZMZf2
rsO7MatO+oB85xnj9NIhxIp3RXCjWkUn+ZCpApLsoL9W1e6dbPRW+yZrFMtx
d5YiFEysYNB2Al6oOJhf4g3LBHPIt9O3AI3GiaWBNLROW3U6tno89b2W3IPM
Cm3A9+v0v+FUUu97eS9lPylNYyoF19iWopsFUorY7bzBzQ67MMzz0V/Jqe8t
Q5y475NvHabntpVeOBOiXlebmBHhE9JZsRu46Pl4KachSeM4oB3CvPTIkCfl
MvN8KfCI9wcXgUUwrbTNGUWTRs6UnuuyuS+T0M4qMQcsRKdQ8RkxWEZfAcX6
PnGcbdzlgsxdwg22LvGiqAlQKZBIm44i5WV0tcuZ5oe8RYXAy4yzGB/uhTHZ
LftCFrbaeDUd2xBNUd1+0rwDY3ydzP9WJmKwIZtrALDjGhTzVHr7Dx+a7aE2
uNvYF7UmJWlltSzzn8HtXKteo1kFitXZFUCgT/vRsQiZTWV7K/31+oeFt2hF
csNL7Oa99FXKERPiU1twCWRixZMkMfzSNZxaGLNB8BJbApBQNc5FCZdQUakf
Zw2fn7mfJ2YyJl0oN/+//mlB47BnkjQX8zOAd8zQ/B9IixeP+yyuE+ji3qv8
yibR7h5QVbWhZJm41dGNTA+NG0uEIbvjq08Fn8xXkh8FI50OjH7fQB0r0W4z
93ISqEZVoO5+ic3tH107e+28JpZl9s+fq+rmRGbdbLwS89/Hm2b5RQddIXqe
VuiKFSpaaeMC0RPVgvob+kPLKf/Q7VoiGXDkyszbdV9teLyjC8b7UlJOKDi9
XIZcgRpenvXbsAwfAHbAWUhT1zPo2o3NZKbxDJvb/qRSscr6ucNtV4di6D90
sHwu6gpw+gpRCWcQ4XDqhN1qUGvaoB7OaZYaO4zV0i8bE2DioPG9kDqxX+MB
uFdT0KEEF0TnkbKTNNulg3L6h8S8bTU5Buy/Aj44ot4PYkzbS7FzSu3LlCGz
41B+tAYcgvtLeSYmJ1/CK0y24gVKDrL/ONaho1Kgt5fWzJ45G38VpQ48zJ2L
TniyLeO8SLT7FYHkQYf0RwfNNGLhcO+aPfQ5Iil422ZpqZTkLj3TeXqCoYEF
wK5PqbsIpOouoPwUYpJUs2BkCf6JYQ2uZvKxBjENr8DGFhuhMjN+4m/aqHDQ
JY3B7i6cnGY+Sdhu1upnHi9bEP0nYtW9t/2MTkAbbNBws6tLQ46IRpQi4rdR
esAuZ9d0HZjPTCKE77aE8Lb9rLMtO8O9W4eMX7Lyr9vXNs6xPrp1ZYemFKUc
uuj+zvzlZemsFNfFiTEjeVsjlGfYutYwY3liY4nu8/ShITNgOMVJjFgL8dRb
6uGx8DcxPGdrKVl7/jgHjUhhd6qYRYSlXyh1QWw6W523eroZvMDe4E8mPiTh
ouQfVnJf703CN8UQB/5mgC37OTD80t7u2UShppvO1PaljVNZUbNdI8nkwb6a
gjHZkuvxF2mkKidqWzSVNTonCRLYiJgxQ2jGeBA5iWDFLE69plhDv+t7yJuB
mw1qSkzH1Tc23VDlcIqL6d7sqs15XsZKCYUrJ4Hu4BxR10eh7rAlqMBs2hb6
HlxKadwtqQciutG8rJpzK5wFKCSKLH1Lkj6SmgFxrcbJibHGVHAPsUYPQelh
6W7lqsZptjyaoknal9QkHeiT1EoMMtnULFe2NrIbEC424D7JNjt978n2NtS2
xWwOSFXe6Bsh7nOYFJJeP2Ya+yEl5Vk+xDyiP/ShU5tx3HucI2mWbtq9CyUt
wT7stYv3fmv3zzZBAQtnGL87ON31Z797HlcE+L3M8HgeKTv0ts6PCm/Ajp2R
hPy9wNBQDEfsJ/Z889HNYM2MY8/TdtpZOD7UXxJi32dEG+PuJvMBvm9W70G7
U8PsFkkXp8aKasMxEnjkt/7MA1kSkmLrQNlkHWGT36dUeYVfDAbdqYIONHkw
2EyfhWxHTcoOKa0QxD+PWU6nuM/uwVMcEyXn/1j8mK2USU1b7Qb7fyFrrmKa
6+iGiQZCXaV9P2sWRER+oaEN6xV5C008kMf8IjRaYTiiQ442UoPm76Ibzm+k
V1YfVXmC5D5oMrLF3x6/XnK6bj5wNCmzI+n1zDxosnYpRBYmBrajrzkD6kyp
083xsx4yfJmtT7fkGYehwI5S2LOwuTKrkgGxsjhaD/9CTGk1dC2Vl52YKzb8
erP1bzkHFmW+TwpjbcCjTiJEDgwRQC3gf9edMGbNRcFQJBIv+HU7k1tYFKHB
kMWpMl7YhdyxH1HDaZgIByihe7fOudB1sq8K/Yv7bpYAwjy2LmkMoB4kgUU8
QfRpTJ06VoNimo3teFHddH4r6yeVBt5ASDXWdjdJr7cQ2h50hL9pE6t7m4Ix
cC8h/BHwBwpgXeybvVnVR8xipa/kQbRP9gc1DsELTPRGg83OIKaaeVOHDbNd
R45BOuuZQpEk0FM0PCDZyo6ekhXRDydgQY138NoG9KN+4FW6rqkbwPs8GUUk
1SVSHNLCg8DBtw6DpetLsiZ54br8iVyYwnZeWmrU5AKCx5tQ7IHIkLBn/UB7
sFlDkzpJfw+W/QjfUDiPOlBcRRJ6gCbFVCS+2444iOX9MgcMRShb7Qp5xcYp
U8Wlb9j4myISlzfb/lA/8wW2LfpkShBz6V7Na8FznIYy6b7v3Fq6WDIQvHcJ
Jch4sCImSb73/JHDA/mT+6Kt45NOD+CHGwYSlvtHVRMEMUgQQvJV9r3LMi3U
ZH51U/l5Bg64VOyxhfzuB3CjpMHSHGZ2dGwukK2cNwkOIBAimkHACxlPkkOv
7EdQiKdsjbAvFutEbq29WnMBZZ2K5PMx/25NEBuuk2VjDI1u1cJM/YZxbssG
3jbaHhw7GGle2zYOzRaHsa2y2ni8C0dWHqT1vjxFIY9qnevSl4N8kyUADdUX
eJGfJFR0+BXwTQLQ6LbQjMovgFsW9WEyVzzriz++h2jC0BkkOyxp+FaVKdJi
6mdCfbm2KKA10dHwWFaNKuqfc2UPwk38ufzwN/3WcYon0bxDHGHh2L46kxMP
reiYiG8puhV1IcnZUF5LMXgm6oIaellkHSta7kqIRi+1GGzfnM40EIAlH0xp
ogKjCtqvpQcUK3dQU+GqSyib7OZxxBSQ9OdwCplwF8qhtBejue28rAOHU5o1
V+Kk5VjbMh75Tvv7sSuMMsPys/4O86qNGZImn2jocN4JIqDIvI/wDmhUquRG
bxi23kf0peGJGM/QkbhLuhUtIv9KMBzk+KUjUJ+O2eG1w5a1j4Kiy8+babt1
8sEr7KWMoTxDE65cG9Whc3C0NJ2InLp8T/8rhV0ac2fIaThERmqSZFQu6ec9
9yp2EfDiOXRjTQC68f++3kjj9g18JAiiTuwIdmDuJE/tJ+LRXhMrwgh7Gvvg
0h7haOjkcsXbvQLn98xJu7fIgiZyhXt91SLvOFHEnyJQmkazBjTOCI1ERnEk
jcf0jmtc/35m3aDNNQ9e8al9HYPm6dfErybQTTaxPEqWiXNLoWY4kcXIoIy0
umTaEp/mZtm92slj0ZraXD1xKqwJhq3M6EvjjjnF/eTcmKG7zteTlqtWWiKJ
zxD33XtMLo7nQkAIoF4am5jDb8i9eYFT7d6t5hvmEA/3eGt1E+/kNuvcPmOH
NUL1EHh/DhSRt1WTUS4VE8thlFmzFLcTH4YwR+nkGouV+k3GR4erYjmlsji0
P4d0O1bvlunlwjq5nkQ90OswkRxjjIxFXoEjBIGrDFjb0mZaer2F1Nu+OO6H
AqHKWoboUKFV7CQcucuETlmehoawvyTvkEWBQ+31nspIWr8hEk2AcfH+VN5O
lS4jvpn5Gscd5ciygwwKp8nqx5tW+addn0QdXDmXyXxOcAjKUajFVGZ3A8jm
nPFTJ0PQMURZRUYHirLCd1Nh21bWPzHMFaF+mxxEcMrVIPFqTnknOeZaOdtZ
1OjR0Gv/lZzDJxu2DPEiw8Iq9NwanghAXv78L5RGc+m6lu0JeflHIejmoUYA
y/ejJxJF4+Nl4NluY8KPUq/GyvuyUrrc4q7NBC4bObi4QAZP6LAdkTtMk2aq
QP/uit1sULRQV7akkOcmA/k7QDBqCauVrMCojdxFGDjLCDRFWWJsfs913GzU
PgjNCKkm9JaNfe1IX6O0EjaispDy5kKK8/CDpSzmY5FTL0/+UiRPAK2lGgRK
/QmJxHv9dmWiH7lHFFLMLkh8yp1UBHM8aLtoDD0Yl3+6iaasEIk5HtsLRdi2
3nTtwbY+LvlPM8Xsu+ZvKnp+Db483y8ZTP59488dB/Q2dIOpSlVBTlXhjgBX
475m9q6mk/xZRKbpyZjPfNP0biLdvMws8kVLg/R9ocyrKzpCWzx3ANXThWOn
5hgrckYdrK51OviDSE3kq7VugYQx08sLd5FaaGaPVh4sb8jpAzHtuVLmPL63
ysG63qepqUQ3KitQjcevaB05Ldo9F6lE42chBoEIbnxbJOcHB/gzzgRQr7Mv
iM2R059LxQOHcg8zQwnCrqKCLsgJHQMP1FSySDKPKd2NabapPrABiMjdVwlZ
IcFSYTpdGEdNVhWDWqIRYpAeM8tEFrSkjGLIc5RjG5mFic+hclYEc+TjLV9b
IefeFEw6l7JfJLQxsLlDN2qsJTmIFwMfcU2wN/2jM5ijb5zzHvBkbzszJ9lK
/xgLlmeDh9FJuwoE+zCsEthlt2XOqRcsbNlq2/Es+MZ+R712jFoc8zVA7DmX
MtrRPFdSLXl5RP67lboAON7gsSA5PKpj9drwZK2s4keJgZtNl96yW+5DGyE/
DedPavJ1wtfpmGINziP5VUEj7SXqSE2gtfRIICpdAAda1knfkFnzsLCyjQgm
gykxjOg3qmuYFHHvQE7DcQS3z/TPjPkKpJotZ7ShhnCnWDt9t+2NpnEGYWql
6KUCA5DmSjV3Ix/NSvHhSmPrJFpykN05o4F+PxW+G4kOljZ6IlWne4o18GOq
Jt65oCmP58GjZE6F6LbHB/j2ILga+FN6p/6NTMybbbEIJieTzBM3XfSiQApt
FKN25RrOGqfeY1anFK+cldqQpWWexA91rrgCPA+nAbbAPfiKzyqLHswiDSfP
r8aKnia9m69HwNqIzbo0ZElE6FFDG2ZtXBpOO7KM5+uhR5ZDKmqOq/S+KHnz
Y6iU539ihVdJZ9f0pahGkVWOOeD/hbzV2ymQiCiJJtsGlx3kZXjEFtOy/mmV
52Wc2xrHUDrCbqpgIiidoiuEXdhklDk0ZaiafF163f2UAw06wEE/GFDEeCmm
Yz99Oz2QY7n+iAgTlQWuBS+sQA1tAmFT4WCQFcbb+dVHk4cleRTKN5ASstRD
RD9qQ8i1hKrxwKCJgokzHKwEp+V7g2knaJjSEChD5B1PT0t7S9Hlzaflkd3C
HqeZjYKvLB+iIM3wTXxZa/Tn+cS2P79yEJ0ueSt/CApzwXvuvL93ioXL+JJl
mqktYGCLaP6vuSj9Ux6H9ss5980eU4q+FeWeTvSJJTc77KJ8gsA1/IOb28eV
98/s60D6OSn5J+UmqdL/+gEgHzSTx1kr1NLRRtgHbz4yk5jrSvTLpOzB0u84
b+tgrTDHpJnr8Ra8gEE3WV5KbWEfi3jT5tBtp12SAThSlCRvIlbgSGzD+KML
2G806Q5BYbtvQThCdD3VQGjsNq05K/8t7SW3uA+BkGSZc4FZ1fa6mN2gsiFH
YFFeXTEcLmOoX4O07VeaCMYFERDbhXaZDUnxQ7PM209dQzmtuV5xUZQsrX9q
EtYS+7c4i3C0QvwlVHxVjAYmMQn32Ob00RWzOQ2POnR2JNpsSay2WxIb2tkY
fNEPqETu6px4kt+qxvJoc/oKbEgfFqf+JgKvv+ivrUCorXx5DpZhgR0XAONa
1w8s0bAclzIcuhpd5AS7NRh9+4shNhaxYwQG4MZ/W+gDgAlvewfLZaYL/8J9
9PAYVaY4WoA1TXgX+Rk1tSQb7VZb1QjBE/BE50Lqe9RZktc/2wL7Eg8ZW0Yr
1EgkCDjjhlem3Vuw1Z/ZUfVss6d/myarEoEPGxMqe21ZsKE5ap96r0H1+6BF
JxCvpESCnNlVM4A2D9R+wd5sUSDlNyq71XR3TbjLV5iR5Y1dnORd8RApaTIC
6W98eXA/MZ97k8xxQKlKR5HOwtHX4y/psV1ZQBQTQVglZ161b3ueCYxZbT97
LiH7Pi8DhKLVah2hiUEQBGLKHYSz0aNzK1inM9VXeFPJEnS6N5kcgOfKuZoV
oQ/Dk6U7M8T7oFn5JV0BJZh0cgMUgmOWFKV8Bd7kXwRL+OsIkRI1DFILPuC2
EaYnodg1gMntEzK22Dki2nk7WdzN9GkTO6QhKJ8wUOBFQhgObqUzUsB93SZe
NyNFSaszi9wtllApZMTuLSI9q/wNtbiw0E2xNrsK9fdBOxqJEZJJawgfGCd5
6dY5iOjNbFN8Ds6/Z/6mKpzVHkD/qg/vCAX1tY/l7pcHaDaRJtJQGvf4mp1X
eih3xPG4BWfnQxWy3uDBGlRUNf+LDRLZqfNbz+zOqOsDn9X1844u/x08nOJy
/iXseBaCJJbpKrAT4laM5w27uYxFXRLEY29wKNZMG25f0QTx3sNEn5zVDb6S
pJUxRMCdWTCtn8VKzYFUUaGVA2hjebZ9tsHxEcXdw1/q6lppCG6QWSke0+r0
t33TqRF+boZlAgbq4M7NPdLR3ksd/FmmM9wJLLMdI71HVlcw/haT17i0ZJwD
li7kfEubOnhMeQLOpPJvhW3lJXg3Fure2X9u34WE4XOuDQVdWKWCocEBlw6Q
D46CCUKGfhNsn/U7/jRK0YHck+IhlRxm0435qcEBFrbSKUZTJojl9CvRSomt
6PgWxJxQeGrIQtMWqumf0TeusCEJAmvoFTDjx7wrg36zSeIo58IZ0h2boumK
VmJwGQpU+7SQyC+VDC68+HP77L664HnW/WA4ehKMsyAb7yQIfuP9gYinZev7
dXYQExAFTAFG1zJ7AMLYk5g7IQXzrQWN1IIa1ZUE2ZUEBGgnHTHZFVxoAoCH
GPTBeW6IIgv3UmcZW4P9B/UFcEya15v2fdpBY1Kb+CVYZiKn1QW6+tRfAkqY
3lr09rA6CyyxcjPH/oTw8rxngevCJF7TBKqgc9IaeQvLNbF/1Ae+Du/b1EZP
5py9MN/v2WsaV6q3VaFTt4izVUYyCKkUXKqgrXJPvhrG5dlvZb6Zs72/g1er
55/qGeSKtpIt49Kp6voqtIXAgrd1oGk0VY3ZL3C2ZuGYldPes/dlDbgkA9Z5
x7yNtEXitZK9MtDNjdhPic0A5vJ0cVNaMdFqcTsF54icxpUMINA5tIGbSj0x
KN2UJAcoarRQq7gON4MxSZETqYavllSxGy4ti+GYTKpT2+1DyUvt1TFXocHo
NYnlwHuwLZZbnPHlFcdfZFwdZpMlp4pRe/1XkBmYGYbQzr1IAaZC9CFDELMj
SzNYGoICHKZELvvSTBv00wpJwE1/wBb4FLIOCyhtaTVypmHyba8oNKK7uPme
F5dI1VEnpAYgp13MUbVSi4Rt8m2rPd9V84x36n/Xop2SJO3o87wXnkds6dfS
W/bQdVEyQLvjiA6NySIQuxiEnUYU7EcIz4ve+/5zPy5iIzkrVaq2crwOFsTl
egneFZeF1mWNTREjXK1Y6Rr/FcvHunItfmHFFbBiebvbxk9ZNuJBsseLO1xI
WQhO5wL5uwowwDrYPMVidwMYU9ut4CcQomHV3Rz/jr5BLCYaMVXH90NstwWC
0xS91NmYpKwBZXp4lsaVsgUIsgAvQE7jG/LQc4JWCKsKMbeWYDS71im2OFZT
+yMU+TW7Y1x1zKE3ZEK408ReyGbPZHQYAmBhyRZlTjVTuIRzkD8z+d5kXzCV
XYE8R8ZbhcnFrcURi5tS7PRB+CKSJsXBIVlsXu8iVOaVcR5kMRPepLoi0j/F
EbHS2sIh+zH5mibk8E4JPlbwcNdiw0ePeqDGQpihJX8lMI/Leuj28HVpomcs
2vVEs9h8mjBCQBiDyKUhR8zi9Mbb92m5ueQxEX1gDr4RgooIhEqOTzUqHuP7
RX0pOTWyjoOiFMkTX+bTzSh0lJqVxb7ZgjwtEHahAoy0XHo2Q5XwRhyYQXeM
vSFvfY2h+v+f5A9WpQzWNOw7CLh5fnkzSVAs0TN5i4NB88IpW9bztRQ9/kg2
H8Ux5bD25Bm4MPOESTxaHpg/4/TYT4OPyLrN01wpsiBWvCgCQvvSu20lMlFH
nCfxQZT57NnSf+DTBDzi5wZJyMnk/zvFOKlH84Q1FxjYAFlIdHFqckqnQDSU
XDDsrKk6hwJ3AUtCYpGxZsBHVTLCp4MOeA7bP7W8NB9qbhwV4G72UCYr/tte
KxnPKfwJUqnDyjdnwK1suZFOpQUKHc7hnQXK8EoIvWEYMlU50RN5yBSdAuih
Do40ftfyuDGhBedNsmGVSmRiwnirdxVRRgX5qOs+nx04qtozjhujM42FAm4R
IRQn2OExD5jjwH+fysQEuDq3FxlQVL33nnvkrI4IZKaYEBDuQm3F2xh2oHBp
BxvsdPDo5tfHNnEe53nolmXhpiwRLm8/+3SOXadHaMzhUempiWBvkM0fg+UA
NUCeAzqPCGY9YOt9qnip664cU+8TL2d1nw0V+9/lZTzsRlpXeCQGAJJlwC0g
62z2MhI2DP8smkCLaMPlgtZS1i09nsdeJZGdNb1Teq59/jTPBZBL1DQjvoh6
rOFA6hpmfaKG/Q48ClJaZAeXgvKxZfIvvLM58QB4xl4QNPPK6vRpYCTjidD6
mHrzeLY0DRJf161xWld7XJdtxWwSp/8nMOAhrLhYeWuaRt7FKL/WcjKq/fTo
4LF6JpjTB/5Ow5ZT1ROX3UzS+I2Fzf3GxY3H7ei5Fwmqpsn0WPfi7wkWBxkO
Ehi2WXUkEI0aPC+aotdltBDCoLynqR8nlBdBTFsFywSO5YeyVSDCWzpuP4NO
lQ9E5s8TNghBG8Pj8gvNYqRaG/liCbRIQ6e3Qj8bv4ZqfQhzXFAIK03JdH8x
Cd8eXs7gKUBH+5B9fEC4+msem8+4fMPuZdsJgCEVSguutd7toxsA11lvWdGm
a7DlDUAkA/vpVrwALMub0Ej/IDYee3/gSdDDpJFcMe+NcBi6Y9Gze0F5nfC/
+Eso+rZvoCNUbEEfZvHE2ezoX+gWxJ7Mu0cPW4s4nwuN+nc98ly1LJVTZjBJ
fF8b1DlTapQi7P3MMXdw07oTNjGOiz5y/uI7ZFjn0qQQ5Ek7MaYz7Gaz/UOb
ZFvSysprVg4wWROKbeHMH0DVJ55Uf61qr93guYnSxGLbKUEBrBAadg92ICBQ
6nsyavdY9uH6pqhTi65tFRobCOql3Tw6UBW1pZR/M2UXXBjWIjsLlY/B2Jmh
pgtUzHpohMA/j6Q/FYmnCvnPIIQhp7lX0YiwRinfcObrbjPvlWhVj3siu/iw
lupeU93P2anTILlT6qQvSZd55ibmswe36K/c93eJLijvqIgZJKqSrFsrroxK
GPWGQIEb14vS8NCAt6IsqKkm+ODMUJ5zoHXJlAlz4srakuo5DJz2ml+YBeJQ
bwS48juRmXES4fvRC2zZplcE+CaH5Hm7mVDcEnlvc7w6LydAuflgEcXDDRhC
21z8JMxAQGrbljVL0D6egl2irdbnvZDxcwPp7W6YD3dJMGGRzbFeviZiyQf0
ZhvTZDp/AIq14atusrWWjhTtAgeHFalsXnuZ3XkAx+kY14u9HbRtZhgYesBC
yzo/HfNmhV1r51TImK7wJrc2t4A6O/gCn73mvRCfPUjEWSK6Gu7c+X9EALqo
/h3lFxMrsiZIyj121VTeI64fz+zl2QFvdOq1I6/7uuUHNVKwAbp0QThfo/16
8BIfrn2EhZYz3181CwIVft5FJKv6xCZiP/oH8INAn5jtULhkMCYdrrK59Mk9
T2EpB08R34jYON6gQv1hu+GIJI9pkp8anS6/mm0OpJhnhetasn9esEVTSOAs
PJc4Yq0m+roUDHppBXTnRZCcdUiS98J5B28DN9yaRify027xfiG2E05O3jAq
GSAgfD9Te3tnzAwVR6FoWwoMGoN8DLatBuCd7otV3L2Rmxuvhg5Vkah/OSrD
BqW6Tj0Y9zEw9BZqW7lEuaeJHl4up2kf+Q4bYjxHzGyb7FxkoZqaeTlY59lO
psq2KDACtuIyCA/xo3RAvkidG+l/ePtVetNKNSxUnjh6nrIoQdBJtPhy6B0R
/str7LRHQbQF4cxKwsYsXosaT++prAtxr8qbyiYFOrpUpQ96HJYxJnk7jfSv
lWe6uBZEy8pSgBprrCaN8f4YJqSB5/oahz/ObN9MG7qhDN45DeAjno0FlumW
OXUkOAlB6kmVn+mrRTq3HXsEtp4jRj4FTBzx5kqsEG7BDHKmvP2ysfTYqld0
NqFW1RK5Wtaatyk0w326LY8dniLWKefmtVZaqxrwYkL9Y/RwxdG8B6bPlpX6
V5JZDh3LjcRjIxVXHXDtRb1wxXDKE0jiDEFgBofAYzdAMdwdq/A6totigijJ
/+NBsrpDwoQ195g17JTlGCIeEGj/BkXE/oaqEC1WXwCIa8pzEMtB78W5p4rB
uA7hEG+eCq6onN18F+/XvJK3L6Q6qjy/mZog0fr9L1iuamNZ7KTHDEH703vs
d5iGBy3K6MlgCS1+uiDmBQy5xKKi6cZdEG/eXial8rw11J635JvIYFt2v6nK
aJicddCxRgYlBsw1cfsWaS8HhDGDC2lu85jCr9xgTbKy8RLENK1Uw2WRQ9Ed
g8UaZFVtNnqfHvZLq0JO1uBJP+rGKx7qJfqil2ip9770T8G+Pfr38vrmtI+E
FXhRn/PhTrHBMBjfHwgxbxyKVu26Bhw7nRxObiUiKE9dtGsCfymcr3HEhWH9
+PExy7oAjBB992i5wxGKXzvFbOKGVPOY3qiYZxD1Pp+aIi3b0N0xaCEraYRn
Eue3RvWbevDvEoeMO1gYh25DclPmSsK6IsPBPRZ30oKUekYKCNOukgSyGSSG
w9NOdcWavpE5IuD94JinGPdDXw7Newq2GkvPo/nXDR+4XZgAPaZIp9RNqxX5
KWjA5sKYiYEjOeWNy1w/hN7fA7UcG7eHLeHL56HQCNSXk92e2kx4vzDHtSIG
e7n/gfLZNGzKBq1SqZ1evOu9+wybnhTmGFc/5szxVn+qtlC36Y6OtkgP2Tyt
j4/EfEg9VkiGYC4/t8f4D4JNZyh4XGFTqoYhOLxVbl0B1cFCorY3V1t2mGrl
gBznIfGCFIv0rIr/1zf1O4k6A413sP1E0xkfEE8T02pY6NtYEIy3fv7n9Oak
1OURoTDOLX2tE5kHJE7I7ZFzkFTCD453YF3GF90B3kJhWM0PNJUlCPimonvx
R+6YPkda13sJiSUyaaBuO7gQVkWczULtqdLuOL6BuQigMzCYE7dR/nd6Mtzp
1jYty+bHziwchwkSSCYtrRW278YX/n60QguTfZDdLpuhJb/6oY4XqwYU1fKm
9RMrsmomEo7ZgSTSVtqcB6V9qWPPYTvvhI6WIuX7WPbtEWFmnQgXLdHm9iKE
/LDciKT4AcOdFB0q/VO4o+nuDxXl3U3mmNjmuqF1S7zpUEAfeAmlVgb8bAbX
0mKKj9Pm3wXVtzqjvbd7ovi4TQklrpCYpjV1Z3VuxdWnUIKraqCxuKmJkUPB
jViIXae0hnnFK7vW6+s0a2Lq5K0SnQyJy+E44icJWkHaU7I2fYfMfVoNSadh
WWUYtdu6q2mWYNcR0/mv/SfqEx9jRc6bxfAMRQs+jZsZlXqry2u/IurPdnu5
1SqcTacLeFugqsghqrg82tv4rJaGyzSmaKgwv9PJSUEh8bUV/8aiPBCVHRDM
RhqsvMGY3TKSCatyXciHzJp9cTCm0yB69oIcRRxJgs1N9xLHBXpLAVGHDuHS
TyFnAQYUfs7THUxYOyPGCZEczrzGa7B6/8DzhiWooOQItND4bU9KKg6Iq/7K
uoVuQnyJZ8w6QATIQQ2NAYRLq0jm4H4hPUKvNhfFd2sohyHQdXqm23r5TsHS
YjJ4riraubOohgZuyrguf+OsTrX4RYHB3G35IsBeQHdm4B/FJhQAPm2+U7EX
XZHczhYUXlsJJAgewO0sKjT9qu05C0m+5XtUWv2EzyPVyq7mkW1eN2F4QBgA
ntvCDzTwTPuhMrdXWTDDhvZhA7bGwBxFcIRU2fiIb0pELGoZEwLioVIK7FnA
2x+d7HVLCjOg9PWbx7VdtMmCgkzvkRyTupvrDZQNMxyGZHphyvzKI+eCi/fv
b+pZHG/q1Dqma9xkCiNXY7RkmCcVc4Fp9pFcY+AtEaBjIjx/lKXYt3RdR0BO
2jboQ4bcoQuGhoGMN4mZ9j6Ky12wTlCXE1d5aanzRt2qlf+cYsT6b6yqSggi
7LtgWb4r2RkkN2SrdIhdNWe6TUTX4RTykFX3NHq7Z+t5P1VK9myKM8ClC74l
zQdGHqIHc10oFNeqc6MF4wEmeZVsb5RziIYGj8rpQbx5W0E5Ly5bX0IfBYQb
P1UzG0vyR37Tujw10WZcgnjiXNROHSpGUHaTlFCKnjpKRQenvqahLGQb0rFi
Xt4c6YGei3ig0n8UMvHr9iuO4fTnLcalBM45mK2A5g5F2/uR3YbRBEEpqpU1
SLX4u0FrHj3HK9gMiNqOFaL2j1cOPGlWNCCr3OCPWjzkrhyCPxlPm61r/aBc
kxXLmQu2zNqhn9nwki0z+qCXJEJDoX4mON9eRuHRjiGoNJLucIenYzsJjCMN
rmRF1Hpm8Wmz5o15rwpLIyEgngjiI7v/URH5FdyG147GHv3m7txXKPODGKSi
iLwTK6cM6xvqMkcUt+4XAIYIFDfNpo0TB/v0nqa167ccPnNNMAcRLNuxMQSm
AKgPLNoTsdJ7IVywor7yURvIzpWsPgTaOhC0yt5znUBTav2r/F+hG0lymXXb
x7X0TqMbnjU94XhQ1v3qNUBDGsb6u66BIWT86D2LUl8x+f6jKivt/WwWw4iZ
mor/7rI/vflFacdu8t4PTNdIy7N/3iPqrBufEp8j5PQGAQmZQbw6s3R5yNsP
er+Q2Y+NDg/8vKqRdwboWUHO42t7FwDGyqHxbuXG+Spmkm1HzIII14eim9cd
ylviXTrGxKLJoLX/pE/XD3QKWXCNKxmGBMVLjEuWxwxwNhDjvoTIPcI46pSv
goJaqCDJBzZ8Lst7Y1HAHTInky/flH1/jzH9hl07iPxV5EJnti3eUX1hgcxp
+3k1aEhFhdK88O/NjfbPRenOyYsAI2giVmPCVwQ1U3gI2M61ksIfCilUUzoc
x6WMhOGkC7xnY7P0Uz/Sdz886EF6KGFrNtCpspeuysFwX3L9CUM4BJjd3L93
hsMeeayfjs+JwBZL6iFJGmnsNsb4EVCwX1ysmmgcM2hT28E/0ad8pEe9ojiw
0sBuDPdfStUrcUCQVPBmetmIdUsctx8+lieofKPLuzKFm9dvasTTa+H+0tEA
lPOdSb4iVkzPfSw0lh7S2tMg5N61IZxt85kICINZ4ZIl7C112ExaaB/cE6V1
Eo/J8LCuA5Ay5Xqul7dO+zT3Vg0/vzz1DIze+OjtwiJzV6uPbG3dx44kAdw1
LANNIS5rTZamqi5hf5spxi1hCOLdb0kbdLhWom2jbUWoRiMkn8uoG/n/7EDi
GiM+2WUujrTWbdblBFfq6jkMC4M3mT2Z+7LZ6b7MC65g2/zMcoRAzM7CBWVa
tLBREqHtM0wW4PNYdrsliUa11Lg+7oBYYy83hYRcJgOniwPdeq/r5+MZqBa7
Nu0q4GCHHuaC6CbH/SviNcwdaCqZQT+LC7/Pk7AFN+r9Ttj3VdfX3NUFF8PS
a773+IgnfiJVomA4MMwiKCFEyUR4lQoeAGmF4DDDxW9+Nw2jLThgaTCQhh72
9Bt53HrV4pONVgpdrV6Os84+Vs152krlrOsy2asRdoA60bPWMzizGxfxT+LP
mzq+7K915vjAcJa7mSpfGFyzBhtV91HlhBqcHktH0c1oFxY2azecheuo50em
B6ZUWL2wcXJMGqE6d/nXfcIrzW1OK3VBJd3Qgc2zkWwzE9LYM5UcxAmIDsyh
i32whrfQuHvKm5PEaMHuxSICdK+KTegWILkxSvbCNOS09ucVKa1tzgqNsFCm
NXNQSOCtsmDvT4ZrWmR935mjk+DfvsnP/sPM/YH8WL062FE1lh7Cj9GDA6NV
plGt1G7BQA/vwbNAqmW7PM7AnofB7lyctRSd7HGml34PR3iyI3uGO+w5t4+w
0dZE92Mb0exEkAHWk7KhNUcz6NcXUxcghYlEAfsd7MX+hNQdwLlzsQUgS2ev
azheUpM596IojQ3P+k/Gg3AcQ0o9F/MxzkTmi5w5XfLpMBxeRe3hrU7Ah6Ra
kvGgEJu9t0Xafpf6QNRYuTBqKHJ/aYBrqveEfdOE50PhT2yPOJdwHXhQ20LE
VGMgYsse3ZgAUaLpptftZBxsS+WZtsTalCGjyhD/1ncIzmVBV7vrtHeD86/V
J4ByWsYR7LpPFz+o65dtUQhh5KwYC50+o7yRHz/tDBj+XVTM6Wp8MR9mJ88z
oRsn/1BWqc0u/45nXbOEhJBw1T6waR51zEi+YdCPJSVjiEFCkV8fxYuKIBWD
SuQ42msFVzlAz2xB6q631l9TFNjA1PAsmz+h14KuXe25dV+WyOYOyTTsjbpi
SD+KXgeCX8RJTURbxbNyDUYI39K7gTmh3vJ+SjrcryVsui8NDe9BwdE0Xooh
mhzFC+ojhi6aGbw5kmUIND2N/eCfadw72TT9x5Ka4zWg5O8qyDoxHgd/OtmO
IYmxyJgFSZfNPybUmkYEbXsAKePh+Is2XTI95aB4kCJeSMt/oplgDo0FleG2
e38UntMdYPR1u5vEm0SHy3Nrd3csB2YjlbFbv6CCsSr+vowlCdjGu6KY3zw+
Xv0WTe6t50rjLGlqlVhMi2aPy/osVcFHUxQth6oV43cS9sw4pRjsxHN7S5NY
syAIB64kkPjn5przD4CQ6mw/tg5wYL5mj0HAaUzetP2dAhCyLFQywLTpwiHq
89WrnwgigFUDFUQXNIcHlXk50qPNUmifeb9uGS9DtkWBx8FpZI3HvxERTPcD
ReiINVfq4/8OEg25Bhp9PERMGOT8U+lF5goRtTN2WZTU68t6oEVegnil14RO
CFqJNmei3F3BaJwTHdn6TFaQLbSId3+8f4VyaITRAp5xZQKH+JTc3U/jE24C
Sw8qf6nxYbS4xUnIUYQElQ22tBR51Rd5FqpzTnUgw7vy8T4M643PUabWT3XM
+uXC7M3TGrUSgzjdV7vCu/3lE5VX/WkspCxW8jFK2JKwddNoKX0H2uJdBfS6
+EG4hezbxpulmPuBeOKURLRj/ogKziJgogxXi0r1ro2cUjJqG/RE7S9fij/M
plcMQEhUmEvBKHVRt179KqyQoVipwAM11NoiXaOSg23qgRwp/Js5gTfUgpFT
d9z/m4uBXxNxxtjTkXlh0iWOQdQC+RxU1EFX/awXqwrCfoZOOhQwGOtli4Vh
v2/ssFISG8b5XS8WzGjpA+/Mye8uqvL4U74nx+vzT6FY9S8XPlFvENKI4MB/
Xm+i6lNwj7btID8XAQY1iy/crrKEyD01IT5HIM1DGzPnWkabodSQavj7UQMO
tNdGDWGHjAAyeyEvndtFEuWvhyZkQRCRnDt7w/WRm9PxXKrLcaKsZlxAoBX3
5su1CunFeBDA7fMoARvSGcf6HVtV9EXVfzfGdgLLx4RI9TyMfbH53ynQ4wMT
sV65Ek6Kj06hdopTOmuNDc9fIKK+d/CcPEkubJSSaZy/kKEpMsVg+oGmg6nU
oOZaZmHJHj3She3amk17ZgIjntLgoc8HMfZk29eVEaY/apW0AQGGNfZRKFEQ
sdPcNuhQEzibq7FOn9HAGmnJzrnLUpcs4iOEQDa5KTUNoEbasp7zUnXL7cNf
0Rk40bgSpfuALJcIb0GcFX8KCfT+VwlfPtD/sp1qv/1ouX+lW57/IjoFjBIp
T51YiowOmN+jpEbjC0d6ywTDGZOHjdg4RUL6wGLH/yJgUSiczST4sTQyZ3NZ
Dzpqsm/H9OkEjpdyNweB7A3Qr1FNIrtscjtp+nSwz8y9kKPue4PVC5a5n7H/
SMCMVcWGCpSY0Agx2pqlRDcYtJv2+DIvVnYvCa9NW5ry5pxZ1tem8WoY451F
66HiQ/HTu9sAtQ+lIXb8wGJ47Gwjxuoeb1mO1w4byM6vUy7BsuQXO2KZwve2
GKIeGmPkM3qIMEJRAxwD0RK19ij7vN6FweRT0us3auSz4OYKaNLNUgF/8Thn
V0jiG1pFoJLUWu/NkUka//AV3faT2r5EylbgWRNQNaKKWO0zEqyS1/eEcwST
BrM/KmhjRwhzO7QSaxv6pPmm2lIv5bKMLx7LAmYy/6KK4a0RBINDmOBk59cx
4OhiCWQ4RhJOLMmVlZccAnxLFs9AP9QWZZuPlzlQc/c8cc9U1cR2j9iiMdFO
KE2Cg24bDBawlWQIKQFF9zYjW7XCZbii03QgdBEv+/+gy8UNw/r1yeVmtIc2
DspX8/XaQPM9+4Ugps+9vbohQP4qshEdRuQ1MY/N5jviMfNKceNbDOgMQAYM
jekhL8IXacPUpsG6nX6OwfcwF3POMYErokmJMn2KQqcqIK8LIXp1jLmcXPfS
FhBqzpbRvYMLBQD/0Sbk+gO7O0ZZlYSMjwieQ0OwoY5MFGtIO66CJC1xRwC9
FiYAXseBLPrd9M6VCd8nWHCaYq6Xhb3irIZvoL04IKCp3JAxIB6bxuTjQXGO
AVmOo93p1FbGwTYAaJfLEhvve5osMe8FOXK8N05Q57OFMhIGLUprJlMzHEK5
LYPoZHhkYeVdrgkcF5x2ylPA7NRmRiXhc2MKMtYtro3DM20nqTbupq1Ske5V
Yawhqqd1DHKGKnFpdwH6n+5WMgURMkm4p2L4G4LCi/gu+eqpgCxfEdOOo0pA
lKR5TNAFw3FCCGKiCTf66IiLFgBTNIR5u+F7QNDFwYjJlKYl5Jm4BsSRvyiT
Ek//gAbD8P1Ty0eEXOCtZgv1BhUdik8Se1bDsExtK/zhZJW1PkNaiQZm5GS9
voWPm4smZ3LBJZSNbOBxAzUHzbVQ2c8E2azWxeKGZrj4nmsEyK0KEx5cF390
Wt0wBy4zQGv8Y34YUh/Fyz3Y3mbNI00BW93h6iG2OEf6aI9bNRwxD5PfZkra
YuW0LvREjiEcWTN6btDq7TjOJShEPApORxNoQBVLs+Inm48b/CG4Nts+TJXB
ByqvDCDHWw9MP0E3EWXCTgROLziLEhzxXzJ6S2NwQ78SOBYs3VEwM+QPWRBJ
kfcCaVpP3JmnYa4wb5w7z1KSiGmaYhLljlkUqRk/J7pS4dlsjNO8xkpT1BOM
yFDEl1Ybjz8W9d7g/rk6RFb6q8AxXMSrO5STscTPT14gJhpWxeHvUPHutgiJ
W9WESF/TTcZwV07i4AZo9gKvZLPaIl3BuwqE503Lw8z2seYNUmYABU/lcUBQ
acwXGPqmDvjNCO3Ivh+lLvDJVBwpK8RX+j3EKUdr4Rmlf/0vOgCmxjZ8YBe5
X0c/2lNktN3IQg5CLM3PwA0KnVFCtEb7nl9FGL7ey4dBvy/LCG55NIgMdICm
9CwKvtGDVNDY8QOwgW8g50RexjMVNcTd7iCp1lQpXZYLQdVO1W++MKp2XoiO
3MNRHmHwORYqRb8h2BSs9lwHSM0+V195dAeRKRcn6gXOU3KzQ8edbeYWKshB
w0joiFfQOAsx6PZLYICiP4zneVBOhXroJaC8e4zZphVq0/WS5sk1PSr49Wft
A4RUtUvuKwGzFAGBWKXD5LnakVRWwMmsV6tgLh6Qo+VoLSGAbPmSlFaj7YHc
nNsDn/mf5eJI8S5rEl6sTqYhuHm1zTj/Dxq53Kt2axZulimUpuLtVzhZl/ZA
Igq5SfWqiyv06EIIDRCxznhM7JQTyG4MY/39nui4SodcCnnsdRIVP8vq+y69
UJcxFC6dFlr48qbohiYrVC76jpXgFfRISi9F2Havre8y7qnuy77dQz2/Qpx4
uPEVW09Weya6+k/iuod55H09Vo18tXCWI1hP+BzLrkpSs/s9oap3c5cS3Oq1
u9KTuov6ZsPPb25i7Wb74JfDhLt6mj6GmhmwQbvPB4zMekT2S3QVQx94cnAH
2AifeuXApJD8lWRQqhg8x6HywA0l2vYfUBaZNAR5WON9em5ZvCocS+uRy3Uk
EzKKBG99f2q4kP4Nd3fhJOeO4Hf1CK/LLubI4pc0jBYeR48bQSRYugOqWF9i
O4QD3aa43MGSjaOkTq/wfyjekDJTGBwcEe4p97myVtTxUJovK2k+eQogJ75l
+miO9by2pMHapaRmw8hEDpc2joilOMUVQPCg+COqehbuUjhIcRGyrNq3YOMf
CRr60h+r094XT79eXVMKNrmY7wng3/ZTIofhE8Q62BroNC5a1AIxZzCr8wcA
GtISwrEL9SM2dZCdyNJ5IkskbchuXztFCEmqNezEsXJGcrY4GNr8obX59SCK
sBA5sEbbkGcSOvcSSMozGmrPZCAVVTB7rqfjVxHKpjjxo2ujnTAZVEqCJARY
1PQR+VsFLvivo2ENjPWeSN5nfCFSjN8rMG6SWIBEM/smylqbbcO6xntJSw78
5b93HFmPpdPHkM1AEzXbXfjiZ9qauG/hhQq1osWvjc+4+cfLQoAvedQtJOkX
3JTPa8Hzz6z7OckDtVFtbnv1VKycWzVAcZrE2UX1O3suiNx/4hGXxOqAmnEz
ZBw1XR+OP9wZpsYClfOkp7FTGV3JmRIeqkqmKbdsRpXOWb4mGscDUut76SFy
SB8P1Gjgmri4pw8TW9SrdyAQ9QavITfa37yZhBIbRwOWAWFbKZI5yUm3Xg9b
xbRCYFNGDVXAc7rSZFyCNMW+DbJKoTO+H1dr7JQvex3duyd3I+u9zKhZrmyP
zweSVh964kxOnviB5yrJrb6S0gQ3bTsw+R7DWugCHIM7m5fHJCCehdL8OI8k
DC8BhArcv6bP52QRCeWaPZd5ox4zyaf0sEms8enwr8cofLGiqNezG3DVV8o6
7GpVHzy5k5j//eTb/uxch3cL45mp7maoxxWN3HFjv2ZfzEKSGKIE/v6S6WLD
dzs+1dJX4qSOLa237mWxWMEWBelEZBFjefxWOcuxRTwLPHBN4H16t0vfutzn
bQFvv7cwoyMTW6hyyQy4Ciwit/OSw0xgXyJsFBMdpDC5raeukAkO2irRWJBF
ETP1DBWZMKQ10OonEZ/tlavi4hvyXRwi/EhNShnlumwM0gx4AYlpky1Ik1xX
ZHsfcaI/GxUFyen3s0eYfd0Fu+RKXjCjnGhMdyNGLZL+rvABFT4JbAdCBf0d
9yNxf4RAQR3Pp04Mrxdv9gxXobJOgLuhSpYg4maVG9iZmvIxtkGjVRSvjNII
+Y/J7sAIP8uJi89nAUNmsmLimEjBonv+5eq5GM53IitVR9JBsSKiT4akyB7/
UvvfN4ntY59YxShUaOcoJ1jvpDC/ZitKFTc93d64DIFYNfkeuVlp4ShdmqiG
jUsvw7ekgVsebR40lLwxjaoFsmO4TbnuvjD3ghwrydSR28HeE2flX4zM+ZPt
l31x7fCgpJzCL8NIWZFI87hlh4thXKIXWfqs8hiYcGKSw0cFvMdPYyOEi9Sb
ETqXbukHlisXXrERE0XOJr6SMcVuPnroB5n5PfxPzBxTnABRsnzSTyVaG0ck
KmpSROSXdlEdZB4xAzVLnpqsJLAg3cSlRSPamTp8vMWDkGMV1n7wDK1rWCvi
ddaMj24uPfot+CNqiA88XuAofD6jcuInL60WqpvkwORSKge7wKDRBwYRLAdN
ItX74izv1pNDVE34rZ8AyD/F5uOPlOqqC8ncSJB2qciYfFO4Rv3yTlQ6Zt6k
lAZq34Jx9YOzZhW1IdrTW2EfQuWSupp5pfAbb39EDvWd8vYey7MC0hWpacem
/yoih0XyYfxnt5km0J2n26Poce9t4X1aiX/Mvan1FwcuLvA9dpRlHR77d45q
mZVpVaI50GqIRZi5R4p5D3jSKNAe4hTYeZOrQOUw4zQeAgKNnTDL1wx5Kx98
PhNE+tW4SUUyT2kaIB9INDgS/UwV+RJnBR5j5k81oDYSDCbTBjUtCWofCQVV
bGdeaZMzf5//tGPPh1y+3fNdxm/+lb6rk+tdnLZFHz6BHL9gt9gOd1Dh2rKk
CthlYGataZyN2cuoXOi5KIkIktUTJPtxKF7pneMpfxpTw50uUb53SkkA4X1J
tPTLa+FIqN17UBR3gbhBKaUI8p+sZbzBrcHNFEE3QwmxN27YNESPX6f4J+g9
psjrYh6UmoHmIeCzl6XwB2w9MJBJs0oA183cuENHfsumQEEym4IhakDvjwyY
nbLu/LytaviSZ7LxK/5hpJcY0f69JbspMRzDbAtpT15yYez0LKBF3SJchbBN
jenPM2IIxele/uWGbvsencf8O1a6RDYckfpxTQGUeyMhwXfigyRLD6F8yHU5
OSmUIvyQZOuJDvwAMvq3lwml/sUnJ5Bdiq9duQzQjqNbLPef9/3ZqMQWaeiO
9unGJ/jSz1GsHhsMegUzMpe2Fm38GgLhcGNVT3ColnCNsPJ7kj1D9SSX5SJx
Sn0m+mxQIU79ieu8tV6StJLv+Vl7A8MNIxEsiDx6dklOtrLacAQNMQLnCy7B
tHDxIva5NwlYGOdGS7n6U8rh6MFV8kx9U6qiscI2nAC1eUQBD3EOTS1WOsOy
joHW7ai/taskFIFNb37ulFlA849hwEjb0EXmWFCAzF6tR9CROHnQvfxDfEnO
xB+LQu/B+aONtAg/jk+3mvci5xOVp9ljS74ugLU2JCynzTMUVUTj/PKpa8B1
RUG0d3nG+x6Mh9pLEZPLKPsBrLizKx0Fob7pr/ZNWQIfu8l/gpQSU9Hmzlz4
3XOZBrsOiTE01VRE+b0SxA5/pjuZow1DsqYeTaAxudIHKEBTSpzq5BY4jVLI
aJTC7sBXSxqqP/jeByYGxK25SoiR/HHLYO8jh+Hz9NBDa32yEzE2hih4A2ZC
Wby3LUdMmrHarvRwYxgcrgKfoVyxpfGWKNlagkLCibpKKZJYyLIcCCnKXuUi
ozCEN1t9QZ0b/lbAtKg7rckXEpKe2Arrjtcf/iG0WIYmagMVzLWqZ+3w5JTa
yIzF8XhWXG++YVjJjTMPZ83qbrzrfNt29Mkf5Ir8/lvXVJQ1jYkYcQxeRHaM
5FInn03f7DLjUu8DUOBDRhTa2Y2Jtz+H9Of5qelJONzjY5jW05qt2I0rqlMB
Og9+AB8J+PGErOepiv7XGu/yJqlyqCPAWUQGmUGIBlzrKm9P5ToZxfbmTnmo
hYssDVEdgMPfVru8/yh/JpBbphraHGvzpoy9LjG6j2+gzhOx2lBVi4sfRj+/
ttC7nn4ukuDOKx/UL2PJ5EUk5+5aBFRViMXE0TYMkNS4jWjPy+yrynVu64bp
mxr8VczddRcBVleg+q/kF8S4F5sPDvjgEnjfS+3taZTIIPYBc3y239diMjUk
q4r1GHp+d+9Fxc5pxOGz4UH1tx91Hs1LVd+rDeTKMA3UBj5KlC2GSZRWsWAQ
9Roay9G3yu4Cn8Ic48NonqX6RKxjf2Kn9TZFf5kyBwKoYTBsbW9GNzG5nZab
hH2BvQsXUB3ncV3QuGDi+QjYxiKTLSOOWzUugPr7jX1o78X799zBLpLyzS2j
iLOOvAoaeiZ8Evv2QjA91N92oGPcigWpbRY2ZbxeXc9VIs8HHiw345Hs1xoP
wIRZ0J+xme+oDIbvnUG2kncaC6QgDvXDrkTBuY6blBC5nTp7Dh476PeZI07y
K+wRJ8CDkyXJlJ0hFfwM5dzBM7kcMMRFTCGKaLbnbEhyMCDxvnpnF35Tm1hp
0ZWdfCuBwMCddwpN9CwzVXX+axrGD4rNSDYi/IknUfu2ox82aE6+mwLOmgST
dOZD1OifcMiQUnklWwyHBTd45MzPbiuPi93WeGXvE9tF7S89Y0nUYh+rOz0t
WlKJeQw/7oGAQU/7B/4PWn5Ko7EKucC4vUCxTxdpcBPVQnuxqlgVFaDFYavZ
oTbEYib4uEFGARO56i5y29wK1XMEG01o4fNwf+aqyyVWlqwQexsl5jkZwpbY
uh2nh8XG5T350OfbhWwpvzAweAC6A27i1jGmtszFS7Bw+PXj9BM4yH2E/Iem
PJuF9WcGCXnRgUxX/YOHns3WQKg9ZPHCjki7O+bfpcwteek93STNRVSoagAY
4auNod6n+c2u9xn9lWmT44UdoMfPwI0j1GBiOn71Fnz3WKGrVPbJgX6eZJ/r
8Np78sfnpkBIBHGaOxN8r3FA+xY6vmSq2Zn2kxP7QfGVuz901ZDwd/G3dg9U
bQaYluwz3biWsdgHRVnxcLSbutNcdvHq99TnLCw4ISwACGOgebyO4ECt7NmM
FoTixxWN+atqe9txcd62Nj/Fw7NY7+YkQsr4p/8TXL52JgMPcpeE9GGKpn5t
xO3Yi+QtTa5cpf+dj4T2QfPyiPkZi6WRqxF2uEhlFzFcdXhcOYNa708iUjgO
4BkpxG/8sPOBvVCetz6wz0JCK+YXyP2rSyrS+Y0YdIURXz6mU64cJDOOLEPU
ad4/GIBZqn7GLjkGt/AgzFAX9DoR7b8Xn9nB2mSkjDdb83Cv56AHCDXzPuXc
HB6UxmBglDHsbvnGY0/UEofi7mn+GrxHFMYJpSFVoubvL0lL6yVidQzyrKUH
vl9j0wK9ZclzJadFZoM+n35ZKXFjljwcXQRuWnAUswr4aNtmb4G3niQZPXkb
3gYk+QtxNx+Kz04AkVrTZw93KdUNft436/D9ljgPPqY8QbnmHvqbACeu6exn
JPFZ0iFzNzhHR2F0I81eircsu3creGwnalMCsrJpszZIr7ivAiRllCXXm0lU
S2/5zzP5jcqW5ME21VTY/28VHlKpKRcYhfB3NNDZ/ZJ3IcQMk7xkjpYYSCWp
A2dGsu21yt0oBFxeEvvgokGEVpCKe0/QeT+anHkHHiL165sLkk8PANSGxi8B
RPp6btzvi3bJV+KR1mgspXHM865oLJIWTY9GqRga1IiAm5NXtyHznlN44aZ+
cdL27AoCD6+ZjMrqdeVkgt6Rh0mjHJ2yVyzcwDhXAiMDooN+t+NZguvjS5N0
k7HYeoCvBSdC54WXZiYUYxgS7gPxWJnS+PANPhWUuctAfVUUY2UuAFa5GGlI
IlFsBMMoLepDyaHVh0+HqltRj2BFizWQ+vvV8/tcArlrdvBRoB3+GqELQQQG
Q2oWhsfmZ7+RMYQ54bSGzqEKubLrGhv7j0ID1/SpvDMcSp+Vm1xMUyqE0L6H
1yK0m3h4oZ2XlPORQqcEBlunejJ7M3r/KyreqmeoXOyPk0TAVWeZJg2BMMt9
8LybDOL7XcumXjORlAqp5ZM1ef67EKCLJ4EheEJ9JVZZsK0eAha2NwODwKNn
4LveydKNbp9uFuA5ngOYh91xy6gE8xux54QgHBJ3OoodbTnYrCk/XcrBA8VX
jywUU8VDsqWIJwfDwrzngxdsD/STVZa+a2j0A3oSx3sPfhaUhdQ2/OvK7HVe
v7gvrcpXuzrF7yb2WcwTvNG4dViZ9rTa1pJnUxfEYlYscVkGY3meFpQlzC5j
wVGMJqUr7Ut1vKvEv6Yd16aOT20tkS7HH13WLx+iqizqAf+r8EAOUbaZc8oL
Qx/jwwHXnzbLm9kztneCRv8sK1XEa2DPdE7CHXzuEtkOP38tqrgVPF3oQ3/N
kf3Tf8cDq5iQO03YX8nBFz5wHpiP7atwBSKpPVn4ZGsMoerZgEdibRVet6Vk
278lX9Ka67lvTLm/59Lp8C5/xEUGiILvHgGaLBuDDIfCwesjUBrRCx+x9GMi
IvBmeJxSlSQ1Q8dS5GOsjuAoAVYMaz74ifXea7KK373sIqpnMQMjnHObcF7N
KKlm/qnXPzpVuV34mEAOFOj/2P8e2jgH59O2YGg7sAivEnM3SndR0DPOInhT
1YmzLFalcvuup+6JmxeVspz5wi3aewa7SC7XWD0J7Cf9m75psgpmFbfUT+64
QKsYzipb7CiMRHN78o8D2IxIpfUk139UZFNpic5WRl2v/uabpAwxnqPc2JE1
GpQNd1/Zy6rjBKIG2Ov++B5vSkB/QL6hbkC8qlYDcBXLc59jnnqZHm54xx/R
wPQ2/Vb1BxvX1vhSTYKiSb4VPXAqNIe+eAo0VYoXR57otrR4HcIpYfUM2rmQ
UBMi6FMefpSWIOhz0JRhsnV7KsNYU5fLQlTpXs1OViANI4Y185HHxi0ybda1
fcObykNDnFnEVf0oCXQgCch9litOj462InVmzaPASd/D7j+H9Mm0BvwZVOuy
Hl2dnpBHyohjagrul86/8lRQw8HERtZ9mGRRTS6Jg+oiY8xi0pG+3g8Kfecc
SpLMXx0DpB/2iihmdV9f/JQ7Lf0u5SwDCVG8qEPzX/F/WLi0Vbnps+NHptjF
0BzL75Dmh59bsg4Rgax0luNSST9q6Gkc/iZsGkifaDYhYp3n7JQNKixol93+
sTSPBl57w1tDfcCeZCoyfD63jzVWixGffekr55C+FV3A9lb18nkipKRu2Z6z
4CHkD2bK/RYyAVFSU6OVpEK0IU5b/W4a2eOEf4LVuueNKwMwn7b29yt8fqWY
yhl5zy9mFQijgS/nU1+e9Kv5MmfS7up+ShkFpHWJbr03ViRR2ZXhMS9M4kOa
dvUJmVr1XT/OawpOQSISnBcA0gzRyTq6fWQjwrtnv5vYeVe574lJoLIjaRw4
YBjPRWX5SIl2/iRoPFIBqHvPfHSugPZJv7yd2VeSB2+yT9a7q6EkFjDoF1Bh
RQOKRdS4OnPhUhirSe4r4T9fnylgpP/s1zgg2+Ro3+Yx7tF6Nm5sy1UyrLQP
m0njREVMiRZgi+xpztN+GPZM29I8lIZlXJlYYTgDg6GQR/ZSDUDL+LHnSDES
7YRMvvq8MrMqpj2EZivPuyK78QU8joiienpsFc3rwSD1/1A4IVhybeAsLWRG
lVTET6xcPQbSKpwV3PMF//WSdB8V3llIx0zcmGWDCcMQZBDeEy/BE2UIdm0F
NquOJj8wplfon11E6l/RAxYxgvY9WO9Z8/I1i+IDtwZEoPSiXVxVNGU5IbPi
Xf5X7k2At0fW3eCZQda3Wus37TSPnOvSziyNll3FfSrMVK1csS3Me+nj4Jj4
oq6VF+XPLhFa41ojaJ6Uo52HiFfsbF4nMze+dObm4Rt9LUQ6LZAW6LY5juKB
Gqd834Tk7ohczzla9XyCllOy4vwcIR76o2jTArWbCEGqxOPlg30jXz5MJVxv
Sy33y5KKQ/bYpDPxQZ7ZMdLNEL3OgjpSfFTAvkJCTdJl209I+TAyIznCM2oG
AZL8sr5sEdMs3nnC/YWxv4S1SWSv93FBKW5wF0CqfGOoNtJ/qLjWDZIipLZ0
rA8irRIUd0ftRxZSGqJqllT91bhDqJORTw5JML7jllLg/8jhITp0PDKD5b0s
gd5tB/VdHalQb1ZzPSrJr5tECneIuTkL3TnJT/A4E3M/P4Jjyn/quPXilaEo
EV0apirPt0JSHXE2j+0p5sHd1usS+qlmgLKk8N6SARzwl9qJ0XdiI157F+ph
yC8CBzYyhs3jx6vwkWD/BVVDgAmlZX1OzkKjd2DOV9le3HhdbhST1OZGPu/O
l6EVeaJnekPkeq8U2Q1EZjAA7zvLFIH3heavgtYCqIyaQqOy7Kvs1GBQWPFG
d3WzsM/RTwgN0QsRjJCb1jQKsRkI5X7H58+KFPunErwu10J8rlILMeiq4WZd
qcyjpJVpWIC2dTMd+fk0scgZvppBMUZ7CxBagJvrJK3T82pLkvUOU+3nsb49
1XSF4MYpqt9oGOnUttp2ZeWh5qk+0+L0Pz7RHDoUeRegXk2mStFcVEP/PurY
5y1l/CbAxhgkKZjQlvIo2lgyZZElswIvaYbgad0uNiKoZtvd1e7h4HxE1nDf
jwSydgg+2fBFmtDbEZuLE8bNZwgdudaFOMN9ULI1OHLfRyXrMUPZh5rSfFey
DUu7JhAHv2EbAi4wYUqarxbwbaar5iKdcrCNtnV3awq2LvTOG4yTL7eCg+G1
ehrPR1yGAnq4+XURBMf94ytH1vtGgqsXUBTqaosS/SegqqadwpkYc+/e0Fq5
62U6Jc74YDexa3euy2DJI+YqTFm4AxN2tRfaX5zR1NwZfLDET6PtJCeScl+g
CMbnyreT86NGNac1zjYaXX8DWbL7Edsq5GI51hdsxz8N5G7dTvA2hOjZhhw2
ymN3YZqZCgnjs8c7J/Gr0t/SACMbWzAv7h8bzBYHiK9u6Ywxdglvl2kZaAkZ
x31BAMyq2pi71Xx7jobGyIEJ14O8+AbPL34xys4jHElgTaDizhIOI3EnwjWS
cZm2xax8sUleH79R5LR1xb/NMxyc2l+FE7be9GnnjSXy198XT0R0BbXbOKfU
O+RFAM+9Xg0XYF8Kp6NpzY1UK6OGaWLsOvsL3pd/tcJBqDMd10iAEqvN6jpD
rEZTIvCTsgvrifuS2+qDToc4bBtoxEp0r8H7UY0AqcCT5xF5oYRvIMTz8cob
TzVImIFxygm7Mf4jUGbZvFmOe5QeixtXIEPELbyQSXr3Y6nS1qXXk9Th+k4/
Vu8FxYjJVbnkrjwFGJZbCPp0hv1rdKSRJP0p9S5WskOGJgZfQyfc9+HheNJd
TL3U+Hoh93lk9qP171XHuNSo5hbboc+XjGqzLKaaz+DLCKnOYb+Q/ZortDAt
K8FldyhBknv8Jb4VLprM66tIqJTnFl1wS8kNS7w+k62G6SLMR9+M0U94/Nzo
RPrFClrZbGrq6S7icIW/OKaMsgHD+lNSq9raPynFjjcETrIDsX4QT71jAPFW
YEscN8oAVDqJ53hrhW1KDCDBLSRuVT9VtLu98Q0+AAeadmpr2zwIN+Uv9isp
RdrD1qy0ILades8ZdFFrsV1T2NOdIpAEBJ5rV9ZrDY53dtD8LGm5r4A9+tVB
B6QRemawVr18SMoA6misNRTkeeJ4GZt4rZonh20ItGCuyWmFxAoZDG96I/xN
yV/X1F6dK2GnJes+3cpE2tUaUqZCbne7rNw+z36LM2BhzV/lKW9jNcOur2Zx
K1Z186HmD1p1nwMRbriCemlDgfwaqQLL7jhdK5WWnyHqPY+coeoeilPdCXqa
hbdehwpsvPwbuSBZc2wzx/QjFaWqpJO7jDv9L41fKweBuM/1o+weIFZGJFlS
8ktgl61r6qzjJinx2wSTtsviOZZWBqJR2mpAI7dCi9kZuotKPVG9nLWCn8On
Mja3wptRSCsZmD0cjSV3rCY7zaGMVT6Q1ObW4C1J9cSXoi6Sth7MWwNgL0yJ
ru8IHi6yTwKNKOGTFAkPavoBXKZes1OZ5sWgQFODH9qL44R60zEzW1Y/FUZ6
jf8lBZT2GToDmmhknD+eKjxye8ojBg9R2GeQRC705qzMv3phqA0S0KwI4YeX
f7d3kavq9RNgB4uYgzUr7mSM6Ce1b64fUoJYpCScahQwjQPooXhUftl0d2XJ
jfNhlyU7YGpNfHODVB04SxTqK4h02vYoeHFCcApO2h4vDnBgcC3stTvGCBjS
nZU8KxjQlHK4og5v38aaue4bTfIDzZcnWxKTDr57jlxXWNpTKlQ/l7iMYRYf
MsiUMmkvQeA4AN+kicx1SF7GKiwLz4QkB7j1aEeJ3YiMeqH5cDw1UK+CIEly
GHlGKHeH66FtjQHBfw+UveWwP0OMGQN1nJOZ1tGkA34xGBljNglCB+3XjWAe
h+VdGXA49B9poOPz1LWbX7AvwcyP2rvoClIS1AkWyL59dYIiXdRdaeSOD6cj
StikE8gsk/vya4IgnoCCxULxcJhbDsaw6P3N2I1QOfuoL1781ycJ+DsUpsc5
7uy03/SpHU2qYo7HRIl2MPEpojgAAVmI5e5XnSYMT2Haa6wH6V6xp6DAnP6X
a9Ba1nwYLhtD41Whw4QfAhnzeCLzRiwtITcFfFSWK94C9EcG9rL1ekBB6oiS
cy4xT/cdXbb/7t9wo7N3SAT1/DrLE0XGdVz9Lx8E32DbhhwjwBsXEG17z7Ct
SgcuEt6lsEbS3btCkJCgqfkVLajDSH+d7Ujvf6fIEJzyf/mEXICxcIcMW1bX
oGZ8Fv1skPrI0Te/veX0tC5Oe0Wv6RI79AEAlSJFHKOvbYLvFR25XTmPYjVv
GeljNk+vYoINFxQY3IvypbWWIHJY0h4R4KNg8IsrRui/SHYXVV3XldQeFkbJ
D0SZVWKuD5CuIS7jqp6yp5ntySiM/8pV82ziY3HoEPqGFtAdQXqIDmCSy96C
pIyv7DNYhxTwJiaqgKmU6sCcMajL6082RxSHMATVDaInMDeU9fe/k8DajMtw
oc97LmrnoRNfJllscp2RgOldjJnQ0/LjoQs8yUcng2fCT+zZb4FPFty4XYoe
JJk09jF4moYxcVmWuu75xih+wg6YG9iM3yo1J8rg6obOXTvxtBwU26M/OOAn
ZZI2rsvLI0yRnH8jY8KHnSQxKCZSASUC1SeuP/w+8wuMmHYbdUHpBshRS94z
DqzQEz7APlMNqNuCGBpcVote99y9OCW7n1ORtSfCJ/lut3hFmaDOy8VPYJ4s
avJ9HogkC8AA4thvhAcC9PNd6kv0s+FUL8RtpUc6vkcN2c9flEjlUvaLb6a/
WOTVBY932RM3gZlH9YOUWFRMWaTi2ADVWHqiRcEgnGH0ngLZlIGQD2V//p87
Uec1fHgTnkagwjglNPw7oTdBV1Okd3IAnIbbwDm1ti3+Vm8YDyYCtuAXE99T
QKfi+nFWGgYSeE7/2BX5K2bdS2Ysv96C4m2iqLGKx4qZEri1ogMx9hmPqdg9
gmM/51ygSjzvluy0MpR0gRB0qk8DJojpcVOhZQhbuH9reco+32Wv4SsGr51Q
6Y8TOfFWgNXjpnjtQAg2wADvMbc1dl/s4bVTtw4tJlVACwjrkhKcWoeQd50J
WAzTsONaFhBWqegaRCxZgQr4H9UBVBhyJclNc89PgsZQMmn9n/HYKjm37FR8
SoG0uIPa8fJuIGoPM+QnTbXFmGpaGRQMXsTKg7CDZceNHnzDBPtQL55Jsswe
2ajDDPHsk9/nuhHvlwcYJgnx3bvfIINVs5UDyAGxY4CtDlu2N7bX68JI5pDG
8JGTUKHu65w50fA2qKeq78nEsfI8FV0IdyKhAeHItygxF2D9nSsMOVX0xqm/
HeXR2IUl05+ITLEIOWyiiKHjd1toVEx2ux6xyMPWVkKeWVRjWSzOp7SLLqVK
GO3DYZN+1LNJFFdjSUITLtkhAzOwavKUD74/As/gEk+G0qtyel6rAJGArvay
YL9GRcV5Rr0EMFb+mJPWPxib1mJ9FU94/krZpUa1sWyRS0F/GWIeceJjeRFL
Doy6tJ6OBqKkq7kc3z0R5TwSsZ1ALTQDdYpyrWoO7gvps3RlraUXGRph5HMI
7b8TIsV4bW1fnJFe26CxGidbbNz6t0iBRuq53Z/2FYIdnlIQSW6M0Idsj6mn
7nl3Wydl1+nI3T/dZj5cPbAPCxjjTXI9hzvt0zZSKsymLoshOfKA7vWnxTxe
xU6cvySjS85bbQqCcwn8l4VRqi0F+PgyFiDiWPyMe441Bc7+BO1LdOFMS9Hv
TYuXScUbwu7apI6/AhkjonObdRRUxrChJHf20iWKm28/Sck4vHNN2zsnjFl8
sMPSRnSgXICa3qfN1WPCOC5LF4OTPtQEUKOQNh9pM5UocJRrRNjtqqjdroF/
Si5rnB4noyCxJc1gHF1ArTCSbJAENSy6aTw2ovsBUrP0q1ovvsiq2hFpjSop
tW3nkICQcR3lKmV0uRUDmXzImayEonIT21QA6Jj+Vyp8gVGyyTv7TRyr8Pn7
YWImDJ5r+u5IOB/IBIJts7i/lYf3tXTPqdI15X4H26jmeHuEwyz/rS0unB6d
Qg+cKnm5FBYDG84FfuD7ru/sXTCTTpaWZJFysuy8EiuYTnjmWZ5uzvjBvKgw
to7gj6UpkCPshbfFtK/BRaSA1u17Z6MFg+64po4QAa/Q1gb1bla9ivGsRiDH
9Jz8AF9UxEI6qlfv0vL+n1cogY9GQUU4n/lnupAMBXZGPpw3lLbSx7CU67JC
BCNMfjJTFGn9kjoPFe3NFAdzG7+vvtq7JttAhXan0cNri01ALdGyZE0FtybQ
GJWBl9UDhLG65ccKJUDQ36qGThalUQfpZ8L2CdN3/jtPBgBslmuFFTvnH8tp
wmgO3zKdOE3UiQ7/boUEV47MNG3kQZDJo/FbnhJ2GDYiZCada/pGbr8m+4+O
xwCgUYsdEx5suYZL14B/3cywhsR0aVGdfgmOSjSy6Hg/E+EylJ06kD5kUOSj
JedPCy26/P/BFU9FLppv/NMuRS2v3gzBcjKyEXsYh0cFRdovtdtBhvgiMwNc
iygx0iv9jQmQLnz0keXMYxXPDUoG3p9jntHOPLRJ3YcT4wCvF1qKzhg7VoLK
mOeh4StzB9wmoTug/cfeTyBvsOaIUO5ha703D413kwFLMTtWLiqpudondpN/
WxCD5YUqNAungFal7GibEJoyX+wZ1w8FvV9so5tkmuK7n7+G8XO1D5NJOf+e
dyTMVzRizFUnOzIHlM5nxVmma9wXkAvxxfpXNOYeaTm43XFVyJH4RPgLF2HL
UMOrNo88TtPhuN0UgtZ0W11Tq3LeGVpHoFWDf8xLL3RANJIsiJGwvNGTpThq
ScVhMhrRZi8slOuM5PvkNj6OPi0MlMXSFkRR5MWYI7/G7bwLXnDOr556B4hk
lHKh5/2rzq26JKlkIqP96QwjG1z5KiPXMKYXSD/zw1/uJIK6Wz7v0qIT+VeU
OD+PMlAgdRhKiDd9yBmOFVIaFJTmf61TTp1TJtjV6Vpx5USX9mxLne3a4sdY
MUq1hKkeWphTkXidbNLKTu91smLcjbC2GlNGuyK3iEUY8CriaGn+BajDIEIE
VH6Fg9JFCbyWs0s3iZ9lvCHVkUdIAbwmAKwOSUTgkvoC2cUbTO03SciFY+JN
eS+LFrI4G2/BfzgUNgJ9aJ15I5hABNukJq+z4yKVj+Aw8SbP6zEV4/xEuIAh
tSN77iS4hX/G5gzD0cOrIkhB/d3oAjSm6rXXdYD6RfGNRIYmIf+9UisODcu9
bmO/o2wj8jsTREsYWqFn1upK9YpFvwH/KmcGwT3EcIzOcclsanrNxhpt9nVB
ENRQtELDusKZXCD2GtQB599CyobXoS0FXtd5OOreVzv/5e0wo2p1kFfpPgEp
Eyux3ZnFYyo3GzaR5VlFLwldDUCzEs/fQkxws0gqMIk1JFNUdFoMzbwe7Ac+
tZnVdSw3Irf7KydSAF6WFYkl7/gEkDSlkZvIc/eKeapDSeoUnxyZkMGqqDoO
ZGgnY3e0lLsfJB6yqzVoYoEU+jDTGjOnoXd/+MX4D9rmwM5/+CwwkW3T3zH+
zlHxl6RsP8fqIKVE//JtmEmsLW7PC6fqOyBZtJ6i3KAGC4wFsObsMvubffpu
SHtCt+XsV7QZKYB5riF63F69i61wV2U7fV6+Xhpkkv9irDgaBi96Jz1MOx7U
SIcpoDg1skQX+BEEyHHbnzcXmQRnq6XXkKoljlO3Fx/Ood3GNmPCyarKr03w
H2heUkKk4MPX6dM27ewwtI5raITNyb0yw/9hXhe4UPfb6EXYmyTcfPjtgHL5
uKtdn7Is0PtDrbqGwm5T+9Y1u8i3acdmxZgD9GVVyLbUcQWeZ5SQPpBF4Xem
wZgrjQxYYAYFenrCOxKi7vIM5jEftk/8VHdsbGi3Jp9dtGjHnsk7bxG7/ayL
pt1HsoxQh+ySZ3aZM2WNGdUSF5WEMIKvHRBRZPFroM+YUmi94W4j6OTbOTl1
dIjZkvAR0W6yLgf9JEfPZJHiqlTt4j2b8cqzF3h4yBrMUtWDRbhm+rDle9jY
huiAKbnUcH+WME9uVIjO8cKLdQ3ZABo2uRRbjRidZ+12Qa2h6btXoetICvQ7
XOrcf6UG0Jr+nErdEqgKaPOXUrlEq1t3ZuU2L6x+pgjcB62dVVme2omNNt0c
75tZ4Cpgrv5avJamufoVpMg+OhoGM5RNqUzzrhgi98z6goHsnLsEk0TextR5
n654D0RBOUFXNav0PlSIJ1h4u1l7c8XAKwZrUEGsrEppi1fq0cxYt+1LjK8/
urVipCVHeBW/l/FIY/Hw8w0/iS6wKMX5r9pcho8UioHVepFKz6mV9rWeXijZ
cHqT2duyHeuRTwsmQqHmVl0nRPDkO4VVeP0Gvs9IWXnYu+lALIlvFChtve2U
+RCbha950vskLD8m46Dkvirt8+w2xAqByk8Cx9iV5C4kP/xkInuZVG1/HBmh
LAa/Gf8o4P+u6bPoPvowvuA6B8uJMt0kPyzWSEwVoS01Mw4ULWynOd0DUoal
9CLZvXrnlDTghTbrnQFIWjfYt3aO3sr8jt5zT4lvCkJUYNQmyTQxMYhYPWlt
1cQ1Gu5+bW2yAFKCmdg5ahnFZ/fTou5HxEBaN52gx5blafxjY1fpp9zvmK3S
A63HeGXbob2F6CHRqmlEtlgkHg0Ptdvm9zFHoMHH5BVkI7TM0iwN+SDqFSaS
6gE4/25E8VTYnzVlX/Ywg3vAa79f9b823WfUR2131/yEVLAdmnHubyLCljJC
ilax0sZeEBCWZNp18cZmP0RbTG7f27arnXfwb09D1zZhUZT5ZxIAx+tltjnl
iCCypRCtguAFf7sVvqIHoz0Ts4KxF5mg3pttbKZJt13uSfcZN5Rmk+mZ5iCZ
Q5KLDVoCH21PU935KZ0yxGT/jnY04i+bzFgbyLRx5Gn975/lXmwXPgJRHlu9
dZEp4cnCrYLSj4hqe2Eik7oy/QzU6GJivRgzRf2YNU9CXkbkV+5BRJd/ipsF
wk/ouzbYVNjT5C8FQCHP5tGbfmTHifuMSGooN+2PI5BzhNwSlpUrMFNpHlm9
9rZ2kw5hRdE1cTG93zLCrUYlVzopvfX4QHR7mj5SVWhdGkGq0CSGumRClHYV
6KSDj14zZ93bQtXR7Yy2C/579HeMfjO7ZQ3bryzN2pp/mlIktcJsZEw52H4k
QRBUq4VF/tjayVfE3CgropfisHlQO6AW6kvTmJjPoZtCHVzX82ggJaBlNueX
XhO4uqKBH5JcH+KWwVQ1XGb6B3jRpkoJuMLkrjK+zwluGpOvafjjJEHIQxvu
l3RMPHYION9LxJvcQxXbb6acdpAZqWHuUKE7sDNu0ZLiEvZt/R5imulFkpjk
fWDJztBeRZPMaCsX/rP2mHgLYdcXlVIj91KVek/nsMOcARa+9dQw5UJVd7xA
MKHH7r53WWjGosVymjQmPmIbwew1IPG6IpEhOklQQx+lYq6ZPUwHhtG2OrFN
ok/VgzODJJBn0Lx/UgtxOazR3Uy8msHOVi8x+T4pT6EwysaScJUM1RNrpJbe
iraC92H4q3W4qbAEowSUcDYMEhzEgJ4/LyvQ+iy9TN3U2o5IgGqrp03POKt0
VnDk72klZ+X38LSAYfEeIbQ8HnKS9t2dfZ26O8C9P4R5+UJpcAQdNM8b3t+F
15s+bkeB2m52JTbW+0FZBHxWzrHTJ4+SUkrUIANAuwFdZQN3Ro5rSWkK+oef
edeTYLwOtfeFc6KjJ3yJkcjfwYX8KLZ7lvENLt+igaryL11wAI7AUMNnFVR+
JnFg6qmwcUMqQzjvtR8wqL94KcwnEfbmJchYbpvSDq4ADgGQ57W6kkZxvtYC
mxMoyp6Sk1BxBK9GXiUZjhKx0YR6CiD5xO9JRMDOrV4xLkNN7eBqsAEYwQe1
wWEde+7UetkpzrcASVf6NG//siqc92pTntaF8gZNBNzfD/NlKGcDe3vf7GjN
mCmsAYV0bdAhUH9DS9U/RSO7svzTAHAekeZERP9QOuysDdDVGZ/JyAQ4HDnU
zYeazbxl2nlCP0pbcHp2Z1LBvxi1MsyKCJtoOfL7EH0XlWPzI/KgiebnsVLG
Cp1grahEQ2vHtX/0kLPUtvhLpyudl4oVRQGYO2jDp38p8p85ydHhutmvjFFm
sLylmn/9LX8gyEtOQ8fdtwb+gHx7zhHkA9moFeUd0ACGEXaL7xMvIfdBsogV
oAWLG6icMBGT1YsnffK14vtR5YIZx3blI8kAUfHaTZJh22EhCUMbH4ToMLwb
9F+niRf2/byPoKjY+MDInvBxS8lvQXNqE6GxL0KodPK7UaiaUCBoD4JgRZp5
3SVaIzm2cGTyKbZLgWt/cIRioOIUR4tX/3ItCkvfcACs/YkdzQUSQPUVALHG
G1W+JpeXCG5nZkL+NKlYmm/uOLpVMcraiDLTsnvYbTpb0Wc1bBnbp2wu72EV
BurQ92Zi9dkmiemGLw8QNKaDGHo4xC8wOdEgLlFtkYe/tYDkkSWTTNFNLNK3
9PqmnZoY0c5MGI8oUnRpNhvZbBgk5Xxqh69JvZaRzLvKI19bBqSfK2KkK78N
BVuQlWi8sEMjVkQR2lNDZPJC7fuz7pLqUmzo94EF0C8CqzBJcg26qB7FMeDo
CIVQpG4rGXq3tqiNrHV+NksPL+f5ZX1G0xyVYjQ6hE+VWv5GoN0Tpw94ozkE
3X5HIUMvnXLey+lczHo1fLwpYmLWXHEIML/+oMR/sE5f/rK96Z49D/HMhONe
i7bjIhUGshYRRrnreTpdH50UncRcn+rT7b9Ed3hO7XDCs3m5OaWV9xTVTI4q
WtKK+qTHA+GdB7yMPhkMXYx0vg8vMPM8Fum+LOIJsmmGYB6IjOmmMmyUo9Nc
B9I3U8YnjjfS6y9oo5ezee7Acp6XMDqFKyhBnM2t5bMKUX3vDVILr4USaFgy
ZeadsidNc1KLohqsqBO9jWGvHz6hcEB4FAv4sE6AJRe7wqtK9djh9JSHGsBH
1ul+i5tpf42GoTg/zGa7YLTaagNSfojzD4tHUdE/+DgxSzsThLIHAS7AWH1q
5sTdm84w2s8Rotc18e4WhL5sGCvXJ8yKToxAQFk7FJ39eujyYvFAWyQBkQIy
EHtqZ9I1zyV0Ro6KQFxGmDwH127hUBPR+xXCZvkYNzfldXPHVKz0WhtjbQDV
ok6sfa+Z8TZTsQZPR6mNVzkJFui7xki56yW+tEdWoNoaKxRsL/qt38rP1aWi
INCBWt1IIG3VL5Hqx2fWRKbR7J6KmYOJU+GBlhDrQMvONj1+XNrkVA7IWbyy
AvhvxEjoRxhzZ1j8sfUo03xbqWbtLtz8Fo76EOx39z5yKQAL7cvozYlbQSjm
p5inUGnV2zPzeiOMePQgw6UQ7MKri5Ju81X56489VYqIhNNokzlF8IekTp3R
xBZ/TUVWS1t7ti7QlSRxDbFthbPu7MDcbFyeXoqxkD0M3cE4rhVX/oJjSywr
FdHdPgVJGW6uI/v0q3ANiHOKjKgff0PSmpKg94j6TCIzDA66BCQBnn7+fmJQ
nmFBrpkc7at9/8+AI89hI1iiElEVZfxFhhJDUfyniF1a85l8RNIHc4fxWwlC
+zKBbjLBGFzPLtnlMiz0YvYkPFSpRWt5WpzTH+XAEBqliave4509SqdG/njc
fUIKsp60sfGqXnJ93d5C1xiT+OxQQVNnAToeWNYlARASu+tP0NXqUHoXE5tT
ukhu6QOKrmPdpvVvnaVV6Vvu0mF9MJhJkWdeCUh1UMD8PIwUJBghwyHRRkEz
Q8193IenIGX5PpKMEwh6gHWGK+toCfiut1Vte91mo9HEdt2sMbQeoqgUWu11
qZxAk6gP8Zea4ZRq3vYjcYBv+Kewm3IsLGy9UDhzO4jCxTqAMZyi5SKl8H02
0JLwMpsvzL5nwRLAJs3Oa78gg1XDcsW++p203bhzHKTAAQPin6jRRpXUq+xr
rx1o/XxQgPHpOXSlzNkRrj29LFQM4tC3Xvib/f/Fo4FYZGRTgIu5nWMKmMCP
W7XtpDJOzqUmthh9opXKL0yR6RqrtKBu/YyWF90CbxjWV86veL9qId1A7Mxu
6QeTPDcHQ4hTyHlo0PTGTLMNG870aLiH0vffs3bJNw98No8uNr4C6+tFdI6j
YUsM0ZUNzaLt29aoTyoi2XCGMmgzFlPHvrcDL01g1GRDphm1/lF4HZslXzmT
qAQbN5PtG2hV4Lp+mQ6oMxap4Jv5uwNuG3phc+Q12hCmERyemmhs2hCygeX4
a8bduProqrkgg8hQoqZbpw0Ape7KHJtp7IlBDRBXcYjgGhAPWkjS3Pbv+Seh
vuSrlCiMh8ooHZ+8LVwQpMTkQlTUUPh/QPRtpmJMsRuZq+RmP1is/8rJSztm
CpGn1xLQpUVBo3REkOD/El9Cfkdd6w/yMoBg+xNlEau0IqF3Eqj0KhzduUff
hYaUb4VYGhPw1vp8EMO3/I/IH6tbOvnoEdgQjLFDkdNIOZg+n6l1t5o+wyRa
UUJNKTJdziHVaJPMyYlsKN6/PIcn+B/CiUY6Z2zs52zbRGEZOWwTg8xfwRBh
64NQPn0rIdbxmtX7+stjOVfCm/+yYIz3Litfz4MVfjQEsqsYRivsYIs6ozkf
JQRiwYSj1+MN1riTWA73E4vwaWTnJ5F4iu34N4o6PBuKKdrPnQnWKMIohvi7
X6MB0ZHes3/5o1NZzDSM33zUa7mglk3KD09d4p/cbIajMkiu8YUC8EquvQC8
T6c0RbqeHRlSedatYT2vVqk1SemDMbOG4OhVPT5GjEVJAyPUDQXTMkGFspD6
yohDE/oYhfd2uoXm745b+Xd28b6mjpLHwj3Jv7YsZEO79holPcFnjbYBN6ok
pOBi5Ti4c4k4zYsg2KZe5FBpHN5GHcXUwozcp+T5RdxyoevdodFQHY2kdbuX
f857JXVgb5RHbz+MekbgRqHQLTy1kbrfvuBDTEE7N7TPLcg5widToSXk0X9/
JWV7xoLloNHxOac5QPAlLaNgAVBHk+3jO1hHVcGrFOy6ILn/4Se5FIXluvbn
J8blbiPrujGklxVXKU+Tf//Sw9CbLOjW9UdYWjBznGhsQOGrx2hfFLwlghWr
rEWECRw7niAqhb6lOWvbLRITew2vTtxXIhc/MigZwYertpdXnprkT5LO8IKf
kmxKAmtPpLQVetTy+pgWgI/kvf5TtV7P/SZ+JHXZ0qZQTCcd78RNfTF6JmLW
kjaMmGiEx0lLN1KHx9gvZ35j6OxKtH0t67gaZoNgTJQCaCuQT56H5eBgNzc5
4J8uza12LSEv6OH3dFunP2PHyMBmgLNyuXltE15cftL5aHteJ8gZAqW3uhzO
s/JM4fkLt2645160COiulP2tr6xjqHgqirc+8Wmp/BvgnY0XIX5gnHLmTAo3
GFqyLjLeHAYsa+ERyklx78c6JPiGXIMaIyHjkmhYt56uF/gu/mOPMhXay309
9jfUyM5UBg2o990kHLtxTcaPlzRtlMjxvE5EBmGbMvH2R9FBfEF4VhyTDX1r
jep7bBqxw5jXEY8mdn93hYpQRBjUMw6X8NHRsjWAS6Str9wRZ2P+POeF0rB7
iICI7vTyv/7aOHdW89r7BVM/qoZGdtKsi3QagyznZfnaXi4s5Otu0ntTij3h
dhhkTALAzKOeRfQl6wp3ztFjANgy7PqokLiwtiE5Tz/KEqSdrLzLJqmD/7AC
xcKbkBGJygDiq1fjEi7N+xz5nlPFOUgdKIjcERiTQd2dPrK1/pZkcMEKkH6f
mMRqXneJZT4T0M6EkM3coHa0j+c+9flS23K9lTvz4EWbSMYOqy2VL1vhvCTH
Zru993/4JgZEcHw6+TQNCjaXaib1hOQW756F5kBbu2A1RGgAji8B2u6ISGO0
Qn7DjzaG6GWVpzpzrMC5vtgMiWa8rYRfLLsYh9bCMqdf2bEXSr7pWrnljYui
YKRiN0JKyAXgQ87CmXfRG6mJ1kO8XjSG2flqv5ZD1QGiMyOq1XM1o2KrtTLI
0JNWc/M+6sjt6kBA8sRe2Oy5RZn1PO29WUov1cGAVE9I7h4wXzcReP7SkDNQ
PZqWV2upmAe+/PcdQNATOtCsV8UorvAP+HoaXKc9S03Jlzn/y3K9fsA7oLAM
FOAJz0nNqERk4YgpjycfbnClb1YZQsshchz2CTOxBosGm4Nc5cGDtXJ4yt9q
B6p3KdP+LO2M313zoPHK+VwvqELU64uZzhXZwjAYRoNRegyKyDIzSYMF4u6m
hj4CKyCq986JpCzlbrzTAQDj5wczhR1CHegzlVsnR9Ndrrth2VanH5jgUeyy
iUV07LKKHFQk2kdCWeXvTM9iKdaxtMmbF4aqI33+sSp1whIKdc0b0UU3WPu3
rML/hrmtV9izcPAixpmfC7qJEAsDRNn4txH6ZepN6K+HiGffLvoGBYJ+UjLM
3Bk18nm/Os6avpHtgFxt1GoFkj9RIQN+0ZGzkYn3wGWqcBVSd4F8k3jPeDo/
RcRCHiLflIhqosz0VNsgN0M6yQiC+6jMXRROXDOg74gBoPyXInT4RbRSyZTg
isgziU1Z/EzhpBlUw/JsB6CDlCXdqu/F0mD6REb7WTFdeLq612+0TaAQ8R1I
Xl3poXv+SDSp1opLUI7PWQpo3g+EVuh0SMFeuptWKAvxQrsMh6UcUwDf3XCr
WwmCWqTl489xLS2OfSZBRov3joBN+XPbW2i0YKTnx7zsypxigY8gIJsOXQnq
91Hk/7pr1XPIrfZPSKWTFKsgzuluwjOovnSxkjiYa/kFe7rm5C8e9SWg4Y+f
nUc8VF20YVZi4N7QFMjJI+ehrzxDxPdVJTVpdDd7SQURsPGUe2BDYQEbTtvG
EJjHU2T0ae+vZZKFxE2EHk2x223T3cvlMGEhJWrGz5VWOrfU6Hn/FiK/1shd
SMy248dDk//eoYO+UxbJaaaB6u1K/RK701UCRLeFsR8pWgsX4s8l6Y8Sz59l
wq6z4YRtozdajtDez51j+T9A3QA8ovEpvRr17qSjnicHvI/1rdI4r5xCfqhx
gYLv67gnnRKLI21o+Zi47o/pl5uNBVX7+ebbOtQ6pgdYt01DKnsmcEB8MsAd
2ORNtEiRFnhuNR2VkEwWAGuDva84hzYecltzJ5Ki0knxz7R6qJ3YsVEh+UNh
j0IUu2j5pRYPwVPLw6hr9CWF9bZ00wfiflMq6TGIt59dHUUhuuoaDTfpT5d4
MWARVUVOKo35dLD8+sbTtu3X/TyaXuK5cPyF1QIGxeLwLO5YJ4ZAE8KEgMKI
VJ0By0QElG+xr3mbNY9PPsJhWEQp+a1reX04ar1LHdqI1WanYvwjsHg6TIvX
5xzXbTm9vcXG4NScWTQpLJX/3ZsI/Q5UumtT0bYIlEdTQJbEerAaH9saZdq3
YQEsSSYgsR839C6FUaryyXP400Bk9Ei5geu809R6I0nJm5hvGBhPz/6OTUDz
tk5RLkvBdRuMHd0QMKckuYHHK861dusOH+cI8OtN7OpuOjClhPqNSy11GCOX
KXZtTbVWzasSflSwUeZ7et9HTQpPHBSG6dYOerLwEiJvaVPFiA30YjBC8ZD8
P2LwnBhlhulpSmfWxp6P9z7tzmfweDUxgCQpppImAGLw4iw8kFOKhB9HB6P4
B/TIWs6BfDnV0OJiZ08s41jMuqBqNAlHEy+ABCJFd9w+gaWMA0BGdhSchtym
76Hsec6r7d1DeqGx5+0KjzfqJXBcCtuHpYPKzVamV2Er8Uip31on4tJYVCl9
oXnxuPjjZJdb3/O9AZjZmAAIbg/oOaZoJ5OYLpCy0HDrT3rmwSH0jRUgqzMx
UWVbmlf2ti2bRsEVag/Sgx3siMNx1SGxfiiOk/vtfJa43bJNrNu6r3opjtKT
OuQ924msHvUTK2epw2HEdQD+z9TsgOi8HwY+h2X5O7QkHTgc5T7bJLMAWLV4
zPjFecAq0ZhRrNd1P/oRTVpTPqsvzbKGZPzP4wElS+99fUlBWqxSJkbwgf5o
W4oU6uwDRqSB09kE+BQ4Iph0p61ov7FcxlnVF6qrl9iXf3M3w+WItyv8yepU
hfHO+6YgE6tdDlgJrvYkcivwiHj9bgh04QRaskNsqWUoy8k2jfPYy9lI0CfO
9On7z3/jyW90c7sMXK5PhsNGWDbCpuM4hMjlSAMCVuxRDl2vaZWnqq5A6HEF
hMZLe0C20QE5LSk+ZtkrksqkIkxYOmFQu3YNUsVoCGLaR0lTTv5ZvGYhm7iX
gT8f0Wv3j0zccbk2JpSn3Bn6DuL+vx+fyOpdxRnG2nxv1dVwDE1iZl3ca/gd
xNd6j58ka5o2cxp4Q9dCasnSHpgweHiLpQRU3d2hvQ+BXbgYwSosxSQX/mHN
RSMK9869HdUBspUJEd2on6h85fOecgBRaqdVQt9HjR9lqmEUbENehaQXbYuA
pk/YIyNkZ1trsg8xNyjbg+zfPXv0yyUzH2BHf8TJrzKWvlgfM5N5/P+sibFU
UU8j/Lz3xT5bHuasfG8tTNNawgWd4UN0QVA/VY7SLF941QE+KTfQ4Uhtmad1
+NxxeoTplAxPu3QtPedSIEK7a/D7FzOlZevVsGIugJbdtHp9a01SCWKibCL3
FFCopLUSlWnAxDj/aRWNyeTBtzcwqKGujlCY/ulAvyjLji5p00BaFsqi6XKg
Br661lJljOAiv+m0swTnLt/5NPz9itfZwG8qMCpKlzur2vbZTm5m3z0aA0LX
zlUTR4KS1Sn3tCfX3dHG4SIckDZY1v21y4EhGZK9ef0gZplv0BXABvo98DNv
UX8GraivD1BQYXxZXnyfqVO1HHmJfb92M8IODyr2VYz5XvR4IaXmLLBi8ZMP
Pm0UegqsBS7SGFNmX68vI29rZltOlPJYNyDL7GYSo+94Brb1bUsOvKuDwRRM
yTu+mRwdTZkaTasqkxZu0e3o9f0oPxKbXV8tZs0Vne0BAKzG2kviiqXZvP5E
fhoixg+IG2REznZ290QxjflDls9ueB4gKuf72oZZo+5wq07A+mbXFDCkGqS0
g53r1eLVN2hUflk0EgFFu2AE0rU8a45vrHoeJWoWOGbc0Ob7aTDDhTFtxwxn
65vC0yeGlYmbxs+D3P+Ly+YMf6HrpchAGoc2BAL+jHBrRxUZqVzxPaayznmQ
g9eQ+GaMGYNC/IO7n3OzmuRVJUYkcuh2MYjsxXCDEYT35scCFBXYXKZ4koxe
b5zgrT2dyrN/gdClOje4fv+xpFcpeZLnWgNU9TXfMD4mU4js7mN3P5PK9Zxk
P5G385ue4qylTTs/TNpPyjtksTOtbeaBUdutyPyBqRbfQ8ABhNAuHO6QKYfn
jd0Uv4gCQVB9nvfa2TfFDLahZbC0nRIu4MbUOwIeKzNcO0T5rkH5G31frlf1
u4jgSrD19OY3eo1tV0f2HoOay1KGHR5gBAbZ+WANlteSaWmZkZ9zBtm5JZKz
kljZIvDtkND5fDIUGUAfXGAmhODhJDR39SxdiFbVJc3b1ZK0/62WUVxL+Fs4
iXr2IMwJ/kIsEZhG0MTSwNSH4LxIe7pGWgtzgUMowSx6M8gI/uyLssF0Fky1
kNje/uMxlIsZmc7hC5/c11eEUkxma0mmETh13BzG6CmqIHICZ1sC+wtDDhFz
mrlzJDLTzpoLl5CF0c/SJOjiVD0b5a44xb4mmAAt9bfEgjimJGhs7d9NiH1T
5fow+QoXDqVk33EUw/0iZlh7bVx5nTVv0zgjeXNTkbO2c6QwaTeCH1ybPTqe
sYOgtxDDroL5wEjMzJ0ahiGzaHGypse+Y5MKD6hXOTpIBH0qttQBfvW0dIuw
bm8jbTbUXszAUtsfDHEdGtE8zuHB9/8/dNSOKStmwRnQ23Ncn9jlKG49PAsz
poc3bOXP68wd0vIKqXUxk+KlU3dQ+ObVSqFv1EAHZaKrRmJO5i08dyXO2nF8
RTQG1Tt+gxFLBf3yHaf4bKo9MAuv5Cfdna8wPqN4GozPs+O/yympwy2TQ2x+
pwM3EZfSV2Ybzc5k9mRCKyu1XgOrpfVEMwkSj2sLjGBxrsN4IULv5Jbl+Fxf
00fUZB1nBtQvTY8aJ+D1cu3l2x8C7WzJu4CrJnmwSLil4ZGe79f5nHJS/uvg
8zTF1+hzmy0/mJbxNBDGJ2uC3bWIBj4l51Uq/UkWzptUivs6AxD66E5/5SPj
2YIYKS/+A9tySBd9BVBoZS2eRH+DWP3et4oGo6pBv+GfrR3syYaoM9+uB5lC
+p8pIkRbaFMXmsZu9Qow7+q4zHGWZzj3Pndlc8DrEXkF/ze100qVe8IvqLcU
IIJzCara12x32O22W561L8amlAnRYzFCx9h9RBK6x2oYZnXUMLFwkSGcSpm7
NP9XNcgFtA3deL6lzS2QL3aQEck8/Jrjyd+HjQ05TLMFV52ViKQDOD0RQHaC
gjOgOuWElUrUEyFeOR9GnVanxB7C7DZwz68S0EYPWJ/UwQYRKKddHKjZ8JkN
CMfc5vMIGUxTCblnJ4z0AIQ00I/+xU8ZYqwlbpetJe9JuSTd/sZpe9NgnqH4
YEPE4Q2zaCJYke5hU1NSTnKXPHoLpa9vMyHQG+BGGLUGd/cBAwBHQ+sviSKx
JUTWg02fnJuNABEaN0xGoVzfrHys11AcUmTv44KxI7/5OvA1uRNC449EzJ0U
hq6XL5lj1VKFsnin3mhPakzEobMk+rPLDpyLZauXEZbbUy0y4XpfsEQdgOdi
14QRrLvIeRlcMAWKRwdVGJ4C4aj7mTetDppbd2NjNTLmrhxwIPjbi0vqxGeR
tClblDfprGc30gqvRdWvvPFtWsbAuaMMqHUzYqGRHlRjy2ld4ldSCfkCdjJu
PFud8WUaP14neCnw7sWjh2vd24XDte8XRyH3onjpHiFvzW12axmAHHiiLSVf
KhzjuQZ1Oi07ZxYEHyxqsOhUK8pZ8ro4vsz+h+duWqrWVHv+g8s9rVn5UP7k
fn8uor2Ea94YLhFmAYvudv5hWhyqKKecYNxA7H1QAdTmu9lly2wM49TUSbfH
gEUxDCukcoSVOAbzn+wR+iGYg/YB9qiDpFGCgbX9HPdUfDViECp50UW+4ETF
qCvu74WzJS5bZU6z1U5u5nWZuLBhbBs6Un0MSnXB3kRJq/f4oxJ/XNKax/7v
W50tgirWvZRiI3vv6KoV3tc0OMktqNB7vhrMarmvJPH8nn0tFKUIQK9Yt7FR
HFvyX9zcUgpO9MSC7S4YWPN7m0gRnBmubgL5H9HbNx2Xazudb0jVH3+Tu0Ik
AIqhVeUZr4NdDqEjyl4hwrAySXzcVYvS3Dz51iAKta2nI1fCZxZRq5Gq6RV8
td2VfTsz+Frw2gLbN9wmlyRyrQQLBKOMOehEaEB4wh2oRwrSP10u551VmV6E
IuyyMiJhIjA7QslUr/iH8MU08ghW/S4lOyD9ym/2r1s3delhHUeus2UlhCPG
oj8VUGznSrbr9ViWNdkNmdrCeQHEprgqQBTymiTtTB9J9DJ1YWGAuoVyOg7h
Z+zDlcFRKM+9eqSXXEMjql9yIqFnH1ti+6sEBW0dk+eVXl4O4ETACk1PL25V
+wy/EYUXdh9XY5V7FjAsnohGbWAdrnDDtQwfyw5DAuh6eaij09IsroZV2fyJ
+wnS+UG+3JzokzmGsGMytXxMDvQ8ylw7HGCMzK1UwBL3hwBwSUaCiGBhLHBR
oEGUCw/jLESFqGE1CxDLbMCzbSnvEQkrw5lcE6WlyQP0qjSEPdbUGfATQmua
hjSqFPQYGdAal0FegJ733G8c45VnuCrITC+9VxVdG4p4vAuBUJDHfu/ajIWf
7B0BzMRLTapoMvaICzCY4G2S/UQHl8PutbK9ModI8BoNmBr9RrM6SfOYRdNO
y3HfnOOEBexv16QEc4ren8HZIoKpxHwTgEs3ITSpL1d1TuoA7QMmr69eJ2KS
hbdgxT0s1gaxP6flxuMXb/b46sMoKWOxz0rdb043XYM+5vXW4/QscIn3qmLW
E9RlwatK0Ae5fxJKLwmDGCIC/Wwf5UhnqReimKeoP1fgx6kRytZSXJc3tZPR
Ny3qX7Mo6lpIVo9h55dfEPTLTsC1Uj6SmyBSdq5NHh8kAMsjEFS0PEayDPc0
D4R6rtpP+sU0cDEqT1UgSHo0OD9fA2dOw0gzFFXQJoxfcVYZZE/zQ1aLvD1n
H1StT5yeUdREpAL/91vzS+Fd4wc1WTG41P1k0u90Iht9Xgc+weTNma7pAfgI
F+GzcsShGpySpaYJX8s/yvKbCJknA7V2E3AMGrAGM742xIoL4Ih6+dMZicnD
q7mPNQ8eOmeFZftGifJm/zlI0VWvcBm9XR2DTR+VVaxp7A/R2yfDd6IwrZBM
9ynvc9X8WotPw6soVlpjGbgGWHpoBcYxbtqZmuuaqqitrGdOU4nhOGpEeYRy
wYvJ2OVh6z5QQ/3UTlV95+hkpXBWwfJpPcqVaoP1P7eSUoIpYJ/b4cLcgTjk
PMVimb9HTsrehiGDt/nOnYa5DCGPT1YVqTAULSyVwrFJrZkicleqk7kMK/xS
B+uLuDhjhJjaXG/O7n2tGM4+bC79odz9KX+0zn9PbGgNgK9fafRzAhuAseCC
AZCbl5UjQO5kSnXV7CbVM140fnEaUzvD+9EyOJr4J2PSV4G7P6Lnj9i1R8kZ
Qrx0BSHPYkl5HWMW001jBCH6LGKCRW99Aj4tIV9wPRkyZ68SKgaNwCe/4+YC
G0HHzeawvqEGNXzNCPXaS/bqlfJE8NSkRVHEtizYJcLyAzpWqRaM6esm/zpH
grvrBLmbfmoZurZIGdddCcSTW8S4pedk9af7kQtWcq3elLcq/0HGexsaApu0
L5QH8P3oh5R/S7Cll/lwHrZnIddmPnzz2Xzoipw8qT8gLf84h1/a5UrPxvo4
Ewc2tzBooeV+yomJq4qi0L0sy43Sr2XdkXO7o1n4d6utMEkPairOXxTze1QA
3XyqK7lWe9PKGjMX1usfjbpD1SVTA5awbujnynQTp+LBxGA7ZJRPAxcLWVwf
lKnOT6ddQKQBVzM8beSy6oRXfWREdABsEkKXo9wV1p2fynp9YBZ2KYKWWtpg
Qj80e7JFotpywJQaEwLvSJJG8UWqmCU/nM8D2eBmEM31Cj6lMU8VG0SFGHLt
Knb/DfMyv5LPYt2lip4qp1a0cMcH0Z3Ny1kSDmPGmcylMMApDSK7Vygkqecf
7SG9IspdiHKmle4syN7MlagbM5F1FpqonfIAWrU5BHMbPi+czANyllYji2A+
7HEcVu90SO37xtO50XxsC3ca+HjcGttLmNHNQPW7+SRwPgzI4TixlhPrSrg8
5Ge00iMHoyjaA7+a9Bfp3unpVQUgUl2HyvrKDSGmpataL9H2zqBu99pEQYrN
73JmBptgBq8tPluSBg26Mka29AbCgSHM+0gRA9McH24cMfjjhbbvjucDwTFx
IEizatGP6S75ETuHlIrTUAV0cTN0agfjoLCor/FoZisu0MTEV36XSs76Qb1S
g0389SqDD4AF5dT7SA7cvycQKQjL1eMlgpa+pIuvwCW4SvUAg3Rk4cl45rSi
dKuNsrP65N3PnMRBt5HcPoPgO45/z8J0yOiOmyAYrq1PU7wuavnDS7GCo4N2
sv9XXLpxKSRpJhDJvBVRgLmaiV8U/oGtlrEiQ6b7nZl62/GLurBPYd63XBQA
J3+Cs32L75u4fxLaFqmx5X2PPDT49VD2ka1jnej6fAD4pUoqQdQrPhfNH3j0
MkNZIZkF8XbBKw5IvN8bKU3W2UwlDAxUQNOGwz1YZh2I2unpiZJG2THhb1ui
mtb2m1UQs0cCEZqrs6bMi1abBt6MYdeIzwmkCBRGoO0E/vYd3876zBtTOLyq
kdedPaRl+jjrbFZakuGUKilZM0K3g/BSLl4/4AQZNWhqzv1ULNo4+Srr8OTn
K+z9bssc91eWHfV7jGzIVY9kQIbrW+cgDRvNbcBV5NUwDmwmByqvvQ36it9D
ZiCeipJHfVBR3uyl3KSsuT7hjaGduRLIOCln1+tmysK1pXCdVFrwwrthD9cR
K4Xx81CKKVOJ8o2FpMQx9gCx+uhIklOG/R3sk4fQiheHmijEmzjAb4nFuki3
y9V+JmpwqkQYGIKgkMVOw9EZ6RMAcaimgbqCjPpoZ0dKHtZKkGOnbfmUyJLd
BoZwzKNMovtIDJjTJqbgNG9fGVKOWIsxQ+bFta6VyXV8zHM7wiz5ceVgJv4N
4vZ3u13ei/DauMDn9mlaDE4nSCD626FgTqkzrEX63RB9mQzG6AqEGLETp30x
993ayMaCY+WuUk2MIM4QhDONFADSeQ8XZIpUWSIa/poAwFRGlf0aBsxanCZ3
vYL/BL/R/F/BcNlpbhzRNG4D51SqrxLAm4hLfmPKQ1DgHP9/jrf2bmQ4gTbm
xRPdFM52eG/sOjYTM3k7L3xuExpwAsPzNM0bcpz5xqCSLm6dZPDzbJ1vAdqb
m6QSedhNlthLn8GUwRR4O1CaKEA+IAmdzR7abZ39c1OQIstCH56fBwHWW8H0
ofEDz+wyPtVXfD7nR1VfLAEENwFO/9mPRPViiM5zYeIeAvoa3sIJqS0CbBL2
1k1k+hAYDoDaKEX5kjCuZ2nhanCQY6U0ThXsyXfQ7oaQUjYw3/uG71aPWfa8
i+KIRbbzer84vC6++e0OXmuPwOk//NQJQNFDRH/y3nze8WEjMiYzqOjBJ4Ua
+2Qo9RftYsKrFYbJlsfGv1w3atzzLKTl64/wPJ5U5+4i6ub3U6y17NKQ7b1y
Ku91adCKr0ljlkFYm5nv+mxjqoUlwvZHvdKte4+vqVWvc5KNKlYAlflhwR/w
hq+RgedjbRbQRLbWSr5KWsjRkMBqxklvnW76E3HtWVNEk8FxdfpoYVtd0rJe
a3RUq7H+fQzpl6JHfS0hCZ8lEiscpghNMomnoU9PgkjMLY0IBx146iGkHeoR
rqOho9GBGROVfm8xP6a5wQ9bN0IR+mfxS+6yCvO2hd0NvuUS4DA988QRgXAX
uJ+Y56DrLMPvVEbz/zgZcVAdfd6uXr3u5G/KqCfaELoeperFSnVQbN5WH2Cg
yMHHbPGKyIOY8pt3hRyetktUYgCVpv53GQOTNL79ZddqjLxG9oB4+nZzjDSO
R7tXbK7RYSmy4KxHgTbLtnLSid5aByTmTgZqn19RWZ0K+vf0QIwBPuXPr6q5
ME6i6kfVcmpQq56Oe8cwc3xcEDfdHzrMP+wmtfXS6R8JiVMZlZveGnLX6Tc5
q3yJIq/4KQH11P+nGzhygxW3tCiqT67ioeoiokLLQGtYJPMv8dHAGGwfDWpL
K22Ycnup4KfRpA87RZ/nFJw+OCFF6aCOp1XeTLSvwyDxSX7DAcEcwG+CBjUV
3d7IytYu9M9biHxrk2BDHT3JEbd+xxG+vPNOp4N1JCDyYoICU9hVVfAlT729
TuclrolJy3pFKKNTh6ywvXvlHHd3WO4xOVXsdyH2XWcloQU+Dnukz+IioZTr
BepgtnwlEJaC9kTL7fVIv0CcV+HauaW1ggSLO66Kv7O3Crly/5kHvJHReK49
D/YPS9NNZNd/G/oEXOVC0DU5zlTXH/cE5OstZYxNA3XRf+OQcOPWXvXSUC4f
PJOMm6tolI7JNbhcaC+MU3gV8z8JdSA5qbPsROl0i2XY9uXInsbbpN+e+MUl
fsEIMXXDYAH4nag4dO7ifbwC0jitXPFrR0tWp7fnEy5/anSTLynhCsoPP8Sv
4UQE9oiPC2VDKx1F27b+vQCHxXXSX4cLY2dcwBsLPfhpeQh4ajcoqW26zI6h
ap+oyuZ0G/cvSzPRYfOXWgaoTgLeaZYAWU6g7em0rz+t9/W3qtFlw54hh6Xf
7keNlH6p8+DtTomLiHgtkGcJ1Xt163Ihq82CJ+kLwoqlS0+OUlo9nzwxghok
EuAa/J+Pah8sR9My/1QrD7/81MNdg2l8zWjmEhZXMUkUX8dNKO4l/A09sztv
bofPzDsvMHETqiNQz0dtL30qwDoQauQgnwqg7PgOpc8fmBejFkiUoJNMvurk
CkPLcd9Re/1p0qpC1nnvc2R41ydYiL2ROD5NYeX8c+mFPbQQ7cVZpPO1Uagg
VdEKCMLxE2aoxdFJz9R+CTmhLXCdLZE1CJpr7vbbqhrNqjCW6QT4NqS8azBe
q3VvLR+BGbx9YimPRlOx8onlWlJtXIbnrFBvatc3jNQmrCuifjOaOJ0JV0hs
UJoMZcHFrKm6ADIrZH+WOwMJXO/3uwSf3w0BUfeAb4o6el+2ZPshlD034rlT
a3f96hNBXHWNFN5iS2G8J/WhNlcdvJz1JiJw3kncRkw5ViXtDwJ49iywi0By
a6MrYT2aY5H4B1a8rl52RAxck+hrYqO6H/gqo7vsljB4UxsbyC+P8PV81Nzl
TZz0G9Lb/FfJ6uXdqEO3fph/y0Q+wUkC3Y7MGfrwa0+D6AkkAtfY2sC/+vqz
WAnuiwRa/Vm22XH5iBvOUT8em+qjljtbL3aokBC4hHiszgxFu9x61kSOmtl6
o5R3qx2TRkZ+dVz0wULdSXMtqyca7kL4nS/2GLcMC3SCZ4skoFrHfAlP1nfZ
m84U2U+WaxTrB9E9HCMQnBl+kxCHXSzPuZyygHWxI+hydt9Z4q3y58jbjT/Y
5JRtFdVnRc78a7rLAcZbYOVSEJvrvghmoYeKWY+87gTrqs23kaz+n2wAyHBE
5S9Q5deeAQGLp4yd7ZkzV3Nr0LwM8XUYZD61PX602OLN60qBvdCsbHSsKlEh
KU+GdKz1RpL+t6vnO7uzUD8Nfs84GcSv7oCpFvVeOaFIPMBL2CzHYxY7ccDA
BLu7aUa6v09+jN61OxNDl3eNu/jG1PfM551x9DnJso322tx3vfhD2B6ZYbpT
ryBxzIRO7q6LhSCVVgRO2fG7FK4BdrDII2Jj0vK1sJFGpPBpFJ3v06IKe5ws
24iPokwdS+sTByCgW98FiGWaP4zXtERhxyl8W7+Lo6lMPtVZp7IcdPFpDkk2
zWAnIu/ZZ1sGv3qDnvz+p3pZgU4lCGTfZlLJPFEC+LgI9VPHhuYE7O7p63uy
LD1I+Ccr71Bjs9ZSaFOuK2IDML+mqXbmeoVBQ9xC85EvSTBJAcyoARFmVqtN
TsggCdfqQ25IyphztD6ds+pcr66Rl+WZWXeqUjOx2GAFscU8P6GexXbsPirQ
irMzPRNFWQP9TZVaj4vX4Q7sGomTQO2G6/3jZApoLKZxwuph7lJP5LTOkzN/
5iiO71BxxjhYR7TNHZSVi20zS7t3asr1OmHLst8wBGNXhnK4XqlN+HDLV7AS
yF+jC9VDP+6YTINHSgCcTtfSyi4rhhmTYqcX20/uZ7LjgrGDchdo0gkFRyPX
qm0rS1ApOnnCwmWc5+nvIvuMzh/25p2XchWgD1hxa/Kjx8lGI3Qg1o+K07zM
nWgfWhPhg4jBb0jLTtYVDhRMQShEVgfW5ONlbNE5/aVhDF4Oj8eMSNAkkp3f
ggtbv/J1nxqUnvMQUaXmuiPOOXJQJXIMEsIFlz1LWH6ycbLWETFJmO0BksCE
ctM5D2C2KyYlv8kfY2m4wePzPTrdVoUrt9oqX50WQY4Se2AGuZCYLvwnubyG
00qiSiKe6X34lgPqtwwY7dDsYMjR3DqTfDKeGcJD0R9fp5WWS7L5SjQKq+ix
McZ68xIFfKr8VA37dFciQK+J/dIpAlUo1nT7dBacxY1cTaIh0B4r/aVajho/
g2EJvotCtJbGXKHFc6+jT2vnHV2M0VyuCpqEK+MBYZE0CnAO9+XAaaIYZxMh
HRclLEFIfII2D5yClsdVGcnEU4B9enB22+4+8YVU6/ljmSIleTfjk/FVwodr
p3qMVqP8AWRxIZyYw3xTXyBroKQB4so9ovYG6sILVGTqB98xlP58QRa29oB7
s4JUUMe4Zo2eiK0AjUOWsJuUnUdcAtwYmZD/dh9AG0j51o1F72C+XC34OIYF
Vt1UDarKih554HhupSO2XyEW/ZJmdOqACp/eeAmzYEoHYCHesEyTy0p+9gor
ng/CpiBW6JB1tbCZ/HAK8AQq7xGUeSqy4q0IEcwDIS13gYm8ppqmWNT4RI78
8t75YkEuS7/JZseg5Ps8ekjtCP6TEuCBSLryz0d9TgK1xnpub5bxvTjR3Jk0
IXrYRVyv1AIBShxogVPw73aIKQ+e0D/HJSAOMkKnsMRxzqmbJpNcJJBVj5on
AvFpIsI8/TfO1DiPzyc5HAXSokArnr8O+NDUmUC31Id5RegzoVTHoeRI5scz
qq162vB3ZHRrlEuLzOK969GgTBhvj3mC/TH3WH3vB6KgNPDAUaU9PM1nIC6I
WnIzAUSEIuAfu8BUAHWMTu9JTMXOjdK1w2dKqDTG8sfoSL6FtxNktZDqym1m
YalMxTKztDdB2DFJMsnE3utzhLIOymSBT5E4HnWc05H1vYgkMZueiOXl121p
SZlzbUVvlpmyuRiVGau8NolcrrYTiGnC3WyDKaHOrcthoOMtrGim9Jq2xagt
5ZCdubhD6kOcIqYCDRKrljrV7vrhFLfmicIPnfaf0G+RDuaAkU2fiBVIxsUH
LdxAfvT0u909ZmPpmiZfxMmQKI9Wf1icBeBHcRynjWsq8bV032dna38vfToY
s8+32dwHKNCbhqhSkXblYEMItTdebDzOPPbzR7ojlslo4/ApXnMYaYUno6AE
vWE3/H1cXJHQWBg0ELWw/xGZJF5V1O/TfMjCc5pKkmslr3uNWqEMlagraqth
uRExfps8ui4eMW0bAANFGHEHU35Sw61O3imfwzgjm6WqlZEIW4TwJqqhZNRK
d/Ikvetocrsc0mJGd3gFpCk+So2fT8ui1NH0OHoqw7qXHXrG7nsqp4WOvZrF
Da8JUoAyLrLoMMh5FiS2xx+ycXWxVUNTaS8CdEaix0lvukdfC2JGtBA8gTp3
ut445llUEC+VX6H1AUR5MEsK+4JfhVnj7Vys2CDbmJz6pUeWzPckJwuw4MVY
Ik7XmWZ1MK6CbcAufl7K0NGdDza0YTSIdc/KQgpRyBQ+zmHY5aFNfXbUuJ55
CugVvbwDxQSpGlHqIGEHjYnbvVRR+TaiYQy73NLHAOIC5ikLSM56piJtj/P+
Kx3JUoDZk6oIkqdSQD/bHcKNwoGsw3F+7K+RfRZPSgOPCjD4yek+o8XetlNi
6MlmKrjxl2fRLxbCKiDaVJtxB8BropG/bE0p8EZQssNTW4iC41KimpXtp382
I73ORPWZJmchorQ4pO02Vk2hTvy5PnljXaRQf42ZirqQtd+xaetU1CwU4/xi
QyXjr9Zr0XmOsT5sJsdYkXOGsxDtzkbKM2L9jr12WibcIIXh9LH58WC6YqEN
rWv663CWZVurgEX+TCafVZotaKVtjI23TLuHknXAX8DbNg/COIK55sDKx/pI
cSN865H6wO/4HYMz2JwIr1bXiz43IIxA7FkktpP+qMEaEqDEH7nplgLiSJ1K
VQQ9TfMeATYas55Mz962FhuznegjwDCddrJDaUqxFpV5Fyz8RIp38irBC8bP
3/f2BTkoQ8rSLAquOy+605jazrRlq/Ql5BAsZT+Ce6Znzhayw9EXIqDWJLmu
PKehlWW4VHfwX7RNuJM5ImM8O2eAx3sSsOjdwqKUo9ji11nHJF9nfFK/Ctzs
mdnJdnlv9Xd/aLbvYPKKohy58xywSVO70elrccV6A6nRZpI+/gu2nfAX6YdW
qF9FVfIVCHK1rDLCE4ILA8z3QOnDsL7zWKJTCd1A8vv6nn9jQBJU86+FbySK
dFR97AX+ykTE1XxpOORBA4/Lcf0dsSbs5DVJHq8UPWM2KJ7UfzIdoxa+01Ps
mqoul/TDP+zgdo8wPDpt0iJY3+1JWcSFoTAjD9yPCujvHn/C/YPljPqaM3im
aBEhtKsVOak/Sn3DIn81HFjrYr7e59kI5QG2hwMsefmJpJUMk5+E8CW/7stJ
S6jwLRtOeWg6/n36/NQ1jfblE4DB/b/GExI4s4mkxVqQhb1G/64wdOwauO7R
gzfOg3FLVSUiayf2lf4EIdSA6g95nqlgzgBqkGsvZioJn8lvSPCrH6X2plNZ
Tyl2qTqUd3sqUX4Aw/h+5xCgy1AcK6zaa9wqoAHmzJYcCr9QIPLilbaUjcCD
WtpSzrQurEvTibIZcTNdABXXuic+gxchAM5+ORlBbE4zIP82z/baW8NNpqQ3
rymaGEuvgICJeg1hnOT4cA10aOxJHcO4eRCAaZisnuxFckE2NHcY5U9i+6vs
aLdVoQ9cIdyvK3gT+LGC7BHq24mtu8e8v/SxBhRCHAKMyBjZigGyGOFNOplT
jBmZS2ZbhcPmqEhfo2Vwq/NItU/CzTHjF2vvHNJrLzKANWABYxTmwsIl5pw7
JplLOxh9xgDLHqIG8zJmlCP6cgW2HsjHly18MybqT/yvd4XA98sR07EQ8ePW
vNVuiOLHtJlXLBUrJ1++BjrPkuCecbm9wg0iypM1QLW06K+uDrJx/4BcKo4f
WFXSpvj2cZxFl3NlHYd4GHHEjJ5OuSgoQR2Pq7K4Kgd6/3yEnZGKTjKr9pIq
JGsAlqCgx4RwTBhPQ3iZPcJIQkPZtgFntpi5nkXQHbhuud9YwicKlIsMjfLP
gsdlhYvzUCCTI7VBjrLZeFmrwCG1FxCLQaDwT0op/bMEbqnpWGaA7mpEPSp7
z2YXXylX40qD6RgZSXMQTmXZ8+wZkwbnrqrb8BS3VRwK6nMQarAXL2eVZLUY
rU7lRBbxTcY2Ux0nGfczkP4iUR8X87Ter7N/hacGhCe9tRZ4FQxOM2LxuGxp
O+Q2Nc5RkTYMOnbUFuBecCckN+raLR2C+38FESQ8P2aRzMqDQroY4IbbAENd
dsFhx+ngkki1w3Ds+frTiXPR1OiGiyIVvnLq77W2gGGV3KVt92PP0xJPnmw+
/6e+dk4cJxaxV7a4vKKgnTdVLARXXiPdQsIrqcrGR0seBEx7nP/gEQsciUjy
M2kW/8dtLqOIdgzebteqfbqjiZoEQYUMXAxV+7do9GdE8HTG2nvqsPPM1gOB
0GkUgzbZ6yX1BihL7jqDYFovLmFh+71Ic2A00YTl0B+KoNY6FdM3pTPZByfq
h/0rfYWLLHthKA1p9TdhD7HkrsTon8DolUnT+pX+tEKXMsM35NPR2WZbCJ5v
Ozce8Riv5qzLsIBmHc03UrZ1EgkjTxRf3kGH3R+t6jabO3KxLvjTp74+Jc7K
Vq0MzjIpfO+BmbqG5bNRHUgBYgwH8MbT76v/QUQoZJBzOoBN+VwXcM+LoyVt
D0SHyXCbSywBvODNVW0/cPVH6Xg3t8AT80EBgK4VuiMmLeAaIzJBDPLrexH8
/x8r9vzuhieudp6iJp7afwLIsojrwqx6N8FohiD7EXuo8b1Fv0d8NfRUxEAy
Dzmmj06bLEPFuDaTt1vBEenim7yTnVIp7vsyw8+KgdxECn8ke+XrLn0dSx07
ukqhWIbnPOHPjOq1Nsm+y3SN4fn2QNlGAWqgOHnMTUqwaTE3d8knO90mm3Gx
9g2ObgGethld3mT/FDFrrcn7pFybjX9Vjq8dmFkTFK/KwweOY8EX6cJvKMa4
R4zTKr57Kx+AJwsdRD8PRnsJsjldsAyzP9AaTogHPFfZbROLVD0wMaNqRRx3
T4aFRnW5mYsFAvSrraMa9pnNvZURqqQ78/t8Ur//8pFGWGEmORE4FBUPNNLR
5CLBStPWx+D1oY30bjVSn4pIcVfGwLhyn0e/fgoQae2bp6oHwunNyI4sD8hR
ok9f0uPVgk6w6eerWR7/X6CMwS16qPDTt2hoQUa7ty+SfbCbAQXRBfK3FydN
0D5L6JaqZFNPjMGEWunPEeJfznLfzmX54O4mXotjZQOrkAM3BJdRcDRHoaZ1
ttVrfx84N8EGLn+4IWQT2rVLexnCms1CE9YO45ZJB08IZ4xAtRXVxpAhBj+O
KxgdDWOg6CFs2Ue9P/vv3a50W1dq3XR8GJ+W0zsyS3kIFk3vr6JYUpgiPKwe
QSQd1G1j0P0v0Kq903dGcYv1UfE0F1Sc8ghDNPbD6t3AgH1wYcbsZS0VLrz8
fStejORxLiYsAYk7sCdSBG0EV9r6FYvMNfZ9o0/H+6UzuGdsA5GmFF1De2Ck
H/CYdVkir1gJV3wrUQ3sTyfrLYbfKBqnjfu0F05JcmJDb4jWDKzMBIHW/Oo5
nsd007fgHDD2e8K2GMf1naLbW9fJmXWFPZ/M5qt9IXQJOHyV76w1VCjyNovh
bFKoeuh3i/jxH/KiXh5qAoh2vLMqqSxefbH710HAoVvFqyzwMTjVnRcxfs5V
On6J2qxrwtBzIs3UxEVnZAeS3h0JGUrx2OEDeeNRyabyiGUSVHEDBQ0La6YF
eIhAuoyhKjPEtYgwY5XupOZ9tzjT80/h/exrtrtqEs6skwUqe9odXlhtMqBh
s4OTcbawLF2ruPWTaBvw3invDFJ+JYCKRAe+9Mi1cvqN6aYGdDQPwzfOtB9A
rwhACEfcpdXaJcggCkCun+R6mXwJPvqLpE1Zt5417So4Z7zdOteZkHMbtrpg
Nt9hunX8D4DTTNVBS2JjxZ6gnilkirj1rlmWnvLIZT5iQQZ0VtZe3UOcTJy3
2m4LGF+2P/2lHMHQzHOCjmscXUo7+ztEaGgcOvXPuSC1XCxFKtPPu5eAkmSK
vC008tcqzdZoFbc2nI8pZucXUwdwgJdE+UtlQfIhMBgwp39d+yGZADf19k4u
z8SsSdV76aMup2h4STr4SsL5CMq/h8xcUoekK1yIxw0/REaBBmzjoK7IvZC7
V3L2xSEKatmnvUux1PFeDIcOyZ5RU3noXH/pVH8Y4k/6xPi+VrRR9mnmU0fc
2yA0X7+F7m/mkljm0R5u/1STj0dMRiDTokerLDAiIyz82f+1Xcww1jJlUbQD
fEBfGS6u9rOEOBbTqfN5ULbO4oc2U1jzAflvzmpVD3PPekM+dDPXAyjHUrIN
8TioBfXyHW2ZnQKvNzPgJaxL5j6DznkBbHnHygvRvbUETtHHJkMV5JeCKobQ
D+p59Rdi+aNESnOGHPBPcioXKm2viIMU6POXswnwARELZ4nktWzlOipHQCy3
WdP/1o+ditRI8VrxrEcY7GlI/2g1w9/JB/+NDLwstQkhFXrgUagAXZOb+FkS
8p56q3RRdu7NYwDlrxd4yV9kiFHLLdZ2ZFpbH24LeT9aRQzjXz6PRPhw7SLd
JfCkQAZDmBiXf3eKHzjRwFj4keKKIWN5liIpD6aic57/U+SWUE+zNtGaTUxS
3aEB0Gxa6eEwrTF8hAQ3s/G2RcZJ5XBN/kOQqzF46kdbYM3c99pI5qWXtvTJ
6v0iYdLddkCd3V/MeiNLmeQ3YMT0BYfXerXj2H41JwyaHhM/aO16wQwhhqWW
8bzrtuFmNOV0MVD8OIsmw3OImcVx2HDIJM6AMNN1vOcf+KhCriTbwFfJzodp
iopD7swVEH2WwaPUsfhX/79uWNRtPSxSLCC5f5jubylocPha8Hcr3c/RSgFX
VgSPpqGTz5imLbPrm8yh5D2a8GVtualCtHXRWAR9OxKDl9/sQnWvRFdZJyzz
O+Nfs3gUzfP2xOYr+aOX1YT8yG1yjU0K74l8VSnxbGY6zXQNiFDJbilOM99B
saOh6o2be9b8mvtciW1jRdL6brt1soyUINXqpWGQrTxFowB9Eu9MLmX/oBrC
R7L66dYwRgFZ5yd3lYDQcQ4hunDwlkod2R/u4ov23V9ITTu5/EqY0+DRTWrb
HmsAawY193RIo5Zo5D5zTDWBwYLopmUEGrTeGXKK6Z1HlF9TDLuDb5ZhqyKU
JkVUPAsSwSOS5lqPg+DAPW0YGCprZlTUiu3ZQHPudza2Acw2npcooIkZDbHy
5x0PzFzfE4fLbPykbezbYoDMOGliMUO9wmizhw3ESEsuaSUpAyNdpmycxG3C
7xq2w8Sn5eqktUvFeOmcfchFGAD4bv+GuL/pTFqVqcpiIgAHFNPJ4WGT1bOu
tzJ5sVYP/yMUMbYMVzGKqO++ynAXeoHR7N+mdu2tvnET/vq4thOf3rcCKttA
9PF8bDujh7K9aNhbz7WAP4JH5r+gEWMpbS1d8sHXutIWpHfOp6Mlce4qccmv
Xf+EisvwWtiSIHssLkgE1hnnuLt9xQTb0oXRueqKIF1qr7N6D0FaVkZw9WJo
DkQgqzVKfEvbUevPw+uKj/0RQpkBgCXpEjzn7DSuQg59eWKMjyYXrUcs8D1W
MC4QBb3jCME+IsX+PF00IpNlJcv83UTPS0uV+OkXtdG9kKGhW3qZwZvAC7Ep
TAi4Yyn8ExtoBunxDQtfoyFvtT+Xqe8GpiKvg1dwB19PLn7R0w4x0MsnzE9d
lGPrunF86zZoLJsBHNFIaG084c05akWykAAYB04Q+icQlg7Nw5He21zMza2r
BVUIX8JC74NkULtL5hRYZNVZC4EZXNIsnxPcVUlDJ7d2mcpkcPajFjVGXUd4
FN/q5YlFpt00vOHD32lYynQtGZRbMkIQ4xQLXAXCCben29f8T0bvCksXnD4N
JmBQLqS8M9xt0FbYimms+s8jtKQVawKfRwYlHEteoGLa/jxQj/97yzDpRybw
S4wpHa7V0TI5aOv0bgkbpqydIBfwWdWSNapEf0QdYn16JXZr1PX84m7+FoaH
BWRSCJQcxYsmgVGl+yAPi6p6DRWdIXyEBiJal2FFf7pP3XuvPaaPg//omJLv
w6UWo2nQXCgTPlzRwt434i12dvVYYdZOkocRBLzSoPPPEzeiHeVVBgba9Di+
VQqzLwfSEvxdVNpc1N7hXAODPLTTkLL2YODGzsxFlVrF51C4SARJJ6VY8JHi
DA1UNkCCSYjTyqhpWND/9tzydQjRGdaKOQ3hL5wI/TIyd42lijl88tZImLxh
XiiWSlfnxoCH/ysBegNshWXWSXxtpQzoPiC8gvP2HGAR+h6qSL8784cFCP1+
SpnHFWr9b9lKDnHVhCqODexTENaSjZTrGD2/PZXqFyTJ1uIv+YH36mQeUREC
z8rNF/ZZvXKVnS/n9+/tLP/qZc2sfDEZr199Np40nLH+VSqtlhoENPD+sywl
bmMBFMK5/R7cf8mNb0p+U9fYa+edxjzDXYwcR6rcvml1rAgeK7rdV9zD1bNR
LnudLorkdrp4QajgqO2RAcyyjT6h9VrMHwy7GYH95sjE948YB13NcOAi+5aI
W+d1L6/awTH5EQXYcu5pMYgS+75jolpp/o9Lxr9+vvTAFGueAl0K22TWvpMB
75Nu92+wbR3m62OekEGTWoWXHysGs73pu2cfENVYSQTJDOMJ5Mg46bZxLysC
k6phNH/VHNk2Hh/jFe7ErCPjMFyvvdzpiDbZAwN/Blo0Gous2gsfJIm1CDZv
uq0zJ6/WCl+QI6ZxD3nOnVa2Dr6TYDVcTCCY61zvJtALaqosh+2X9Zvxcy5d
Xxkef/8YmiIZlh+cruaXLLTdNP2v35z0gya2v/HWOdsgC022K+Duu5znhB5B
1XoEs5kJxFQTS97/BfsLblFrZJik53i0XiuPCq9EUCyxGtm09drZlkg7VM2s
EJl5c78RyyyHEOUGUUD8T/QUAa/8TaOhLzuyA1KIjlGXtIvcjLrE2katehwo
yhtt/RxuOz/5Rf668vPyysODadeM09CyFsmWaMvJJjIP+f1FZOjkP+sukkg1
lyqEWKRI2AvjAckdTkaP8Xyx7QDLO24ILRxI0ocsVl0M6Zvn7alFTBxhYX4p
OJ99Em02vO2IJ1jAAKJFXcxgCqEJaubmOLI1NwB97LsNtdRaZ39fOLk5DzVP
Wgqo8tPE9UuY+FAMU2ez10yfmbv80jBv2d3RZtHO0njDTsuRbkTtJNT/4kW6
An+IrI+YsWteZD6xXo78wAFV8WwtACXIIO/5+KlHHRIsSlM3TLhIj4VAbRSf
rrNtLCkTCOFdPJ2T0G4glnUmrtxiALOiMCoas1Uft3XSnPFTSQibxh+56Pi3
yYcrldVczCyGle7f5JTZ3cl5Gcrb+xQbafwGCm927JIgKq6q50iT1MNVMnaT
EpW7qAR3yZJt30dZNy/fiPn63P6bXDR/bLd12Cz8ONAy37rSYx+yfbTqeCr6
H6Gjg6l2Ih39AXbxL158EnEPK7rpiX7Lgm0rrgNv61EqHUox1PV4IU9NYvql
SC4ifT4Op8OgK2BuULGmge/+MFcUw0uZ8YNbF3Zc2Yj2KSN3l2uF8nqHhwYC
7w0dWzQbEq92cpA0hUf7a+Y0GnL2VOjkeOOE/OhR07E/4CCu9HTaJ/2zc435
1Rbyonm834dM/vekF5x0W/DBKCHLSTymwj01Q3o6DKCTDr+05awYkv6SYxV2
B3Ksfl1CMBE8fuNDeewPYURpg1hjWNo6hCUNPvLnmT9aHAIxtuWpFdjPGNQ6
2S6GBISlDoGncdEIZyMFRPiO0DtYTl3QiVW13/8EVJACz7MXoazna8N+SeH/
65E9r66IkXFoGH/YPjeP4Wz6fpltwhRyzDV7+8QGu2xv9vPSwrzH3YQee4WT
rD3HZA276zVpArJCA0zfZGOSVd8rzmbdl6kG77LPdcILGfByc3ubE04x5HH2
lDESfdxCeEKZj30OGkw8ZeYiw300VaeYk2vD3IbR/9N/krZ021mF/HJkTQIg
x6hrSSYs7UTbDGBcuR1gakMLFXgTrOwYiT+pnx2wuzqp/1+oD7T3Czh/eu13
c2UdiQ3duISeRsbuAXH9els56nI4DUP7IMEVm10ufpOZ7aXLtTFuEBvKlG8c
RtD0vHgHAcSYZb2UcnZiy/9uwqxv5YLcjXfPJKjeUs3YsUhN8gfTF3yDuhds
kuRlujs8Gf7iKVuuErLVQdqRjME7XgyTQtX+Ff2O62I6nilCNR/P8LzFW4P/
xthcV3FZzToaT2reV7ljQND+dvnex57Hd18jnW1X8khxrBSAsfmVHTugbq+Y
NUHpf0v1GIMOmC3CFvFK5Lo5beBMK7L9T6DABanu4n2itF115ZJitJ1egTwX
0AIqOCAShF0d7ORci7OirwM98gez/Nyq22YciAdQxbwc6PGUK030N1uwPLaE
hdgXgO9sCoQHoTtVpp4JRU1Bk6JEjjB/6Vqkg52uawcbOppn71q3u5IVmXIH
7cdm9IUZhQnXjvnBpSoppBvV7X7xIWj9vL/kW7i1uz5U65ECyXVcesCw1J5R
x0+N5fas71XfNI/8oLd563XnGzCcMKqdOWTREWKj51R7sOXaL7jt9qvmwq7U
5lZwyen8VKhwnhwIiSMcCjfTEBBS0Rr4qa70BMSGVoRvx8HXCm+S2yU3bJuf
N0XbTZQHOpb4yKxPS+Hrwlrlf+TLgpU/BTGZGS+e/AbeKnL+eO4lsqjGkMk0
jNk3syEbPV7CeIh2hffpd9N0BIXw7mgGkTw15I+38ijZtr/ClLUqXtdc/neK
AOR3zIMdTGXZonhgBOgIpvyrjIuh1vDSFip0H7J4z9B435mUnI3Bow8vJE/j
ELtMobS+h11xiwVlEqlOjbMqTVl3oIYcWp0YcOL0SDz1HZN5bLg8Ojg0C9vr
tZ1133dQEsRcOpIri6W/jFxB6//I+t39NAp63DbZ+lku334mZw7AiEQAud9T
eOZxuX87UYg9mBBvPMXcmtD8kRu2qDuEmsZGz/f6+PBHYh+u8R8XrPL02w93
wG65uI38bRKs59SKxqgk3yHlio9bB7mYc1XjZMkvW2Lb/PjthGuIGIs0kPHw
kfvmDugzCPB35T0RfynjoaAXH+5tlu9xqfQtsIF1LGNub5/i6cbleoelVINc
ERCWFiJ+ggSMG6xTeP7Pec6qPErswGSopCl0pKpDheXfiyhFJwGd/8pSorOc
xmWSPvs9iVFfI1pK3O13h7qLuV0P4/NL/fea9WaNlSt51a76mWBXzV5d1vwi
2nlXEhCs3cIRRpOO6mAm/Wzp+IpJ10y9ZfGxJeuF64NeYJm6n3ivv+Owy2GB
+yb6dAUSLedOU609zAlwPTEFMWQTm6wgmYCtxJyj96I3lFjnn2vs8xdIK8ez
gfAeYGKt4D/u50G9kkxpxx0Ywa4phBnQhholO+tkg6PiNx57gXnup+yGxvUR
QqyV1c/mBEJJpjHjyUMx6acxQBH5CIILZDw2uOTWV8XkDfRRTio+rCisqJZa
JZIB45nzrdvFGIvpGcjg8YvH3ID6slRa0MOAWWIRKysJYTHyeieoOx9uYVtK
NPNbZCeK6aW+TVy15TpxOMM72HuMrFII3cgK6yeZUy9c6QqDTpdw2BIEd/CZ
vNChMRmrP/T+YmJj+3TH1F4ezjnF7GLvseWmMfC78LSWM4JGZQOiofNlK31Y
9rdbItv1klNRkLIQC5bcBRf/iPSgvSl4Xw1O91BDOZ52FUPHFe8EubZSJ0y0
sCScgafclWZAPiUbI0Vns0f48+/ofOKNuywMIvmCJ1T86JlZ5GiUSnU56u58
1xJDh4z6IuFJGuI2u4VE/u83K2dQoZxHhfhNmzy2KExiOJsaoAngPfNJfOTw
JPNwblqXCSBhivThEIGhmC+XZvDkBqQOfhtQVwY0jiAaUcKhrIyttD9+RIW7
6sZ7MNKBVTR4RLJfLgHo8hftyIbv594Wju22Hn/hgrIeX1Hh6THBueItT5Jb
YxVNy3vIvy2jR0U7gWJwZb845IM8wZ1qU0ALaDId5vLpIEYn7+ZsA6lhLqUv
hpWx/H3DtRS3HxXBiG81+zMmBUwGF5/W1kcRcdgrSb3z516N1lDRwd3sDQ1d
4QXssIhzSi5mo5FhQfpigYk6oR3rWfY/rDwa8c4dZSjbEgAGQFXQgOGIEYDQ
htsDddcR/WY/SWWs3GNcEpasXDw8iSWx+S4MewNv8nzQISsSxl317LJ0sK8F
koTLad2AJwWw+d7+6zIvjtE1mTg6ILohRnsVdEM7UzsBa6/0ls3VZqj1OsoJ
Jk+jihZEutLr0xE67IBUqGjV2bFSmwgSXvKc1ksGnqqip/skBNxU7QE44ggD
OTMO8jgPTrGaHFTDm+9yCEfgR+dBWn7FO+s7F02UcIi9jpGOCNxoRsSqGG63
e2OYNV6T3HbN2CPr8bpMoi/Il7d8oBKhc75A/ctC3Mk/nzStGVUB3nz1bpwI
oBhCZ3WZH1DhuqJtVdYuSH5Pgh/tcFcZ/38wG0Ltyy/iJqlWentaoaHcj8B3
o5jJNkktVwBFX5KpFplaKtuOTWRoe0j3ll7P5F4ngXQpy/P6mFe1YhyZIWdu
wL0SFOshc3/CM0OnbUNA15q0pzMNPV9dI/kB7/2B4YT2h+Vc4uAkZwHB95HI
tpjJvrXDv9qLOeRhs55GdXkMar9jab0ytX0tUrWwcPJmrB2MCt9oQNLoI0Wa
JGtCbhGomp8rq18GUICFs8AZeKnzbAZS/VP7ak5kB1GrgL141G6ewlMJnfyn
l+BfdvI3vs1it4yQ+VajMvGeYACtlEUjhL8IUYLKKBz2jvrEcsC7SEg5WCsC
AeZJVmvLNPYFtRg4O2SsvHAhP6YMdx4wA3w21MUnb2jIBqbTcWItmt0aKl4c
GvCvMNukmMYTTmJNEMA/KLTlrlm7qiUTeRtRQ4S8LmrqLoZv+p2nRhacAckc
5hV9T93J80qinLj5HJ4kaAnKASKxx2yyFee9L1njQUBLzapARhwX6ju/drZt
UzksTORre1J+bKZSVuM1rm+G3U4l6tAIcTe6t8VvC3x2ex8aIAF1LxA1PQL4
aqpmueKFKKIR6YZrrZxTx4JsCLxLZbv1dkoscrXlldzRgnJLIdlR9VMLxtZP
yKPFCad+fIATyJgLTtxIJGM7gpfbt6GO2XOo/z9gJVBXRpulPD+2CKXwgJr5
+ThYIzQBHedsJS0QHee7G1sYWkTq9CIrfiErHEVXXpdL6tNECwmL22VCOrAm
xpIAEoPi0wS3U5hwtS8zft3GB+IvtyQlCa+2W9+YrKm8BKJ1fB6YQDPVc8ZB
/q7yxWbjgbVcxa99BkXr7+gu2poxhlXmmKbEUK4Ra0r61SNN/ohOWlTIXImj
4DMAGKkCFil2e2DohHg7uXT07yWa68hKNURoEaOAQEzfA2krjABxDFDjqkWe
x/b631GaZ32ab8gHPUyMPlb6s1gIH3sK+C/vE4d78XxFfvImR1c86aOhoCdi
axhoGYnw4UjnjlzQpi/jF0fuRoHnia6SolWayiyDUrK7HfMZbv4TPUGORsSX
HO+C8NKHH3USDxonRMwkdCu50Yx/sdVh3e+GhehFiOfiYZYzLHrVKNI0ssvF
X7EjRQqzfVQnKokd41NlbnOrUcLAVLPzAG+6XN4RLs7KuV4z4WJVts0Vj0QC
d8CWwkkuLxU4CFCo+FS2NbW+Eujz+YqbSfSHTSc87Cim4YEg1seeWNaWRbl0
qcK4wwQRVY/pAUqCgJChBrmzpNfBT22FKLP+cy+ST7okME2o6Ewbj2niknXC
9iwaKsn4hnq7PB+Qj8UhSfqYeM9+ZFs4AJgmQ41N+28UQrh9dsihRjPDSTcW
2zkSCP1dW/OUz7wT5F/eiR6WOu/epCsEgh69HsGLJoQW8n9O1a534zvSJdtX
cyUhEQ8URkaMeXa3v1MQi3yhXLKtXMdMwioFDJZAjYfRlcnhGB8MPrL7Mgwg
gvMfEnvKrNipOVFWJ7vD2lASKYTBCixpWgpOu1RsCVN5SN1BDBl6G1KwA3HZ
cI/QBCB3OmubDjGwRrf/FHdwSxxNfq7uzurgkkZbftCYmYwOHo76+o1xSUKM
9p+NVvWXIitRJhWG67MWtTJTVlkyPYSjh6jS9lSa5Amor64GpzaQLAR1LYK7
KqbwP2nl/+2CeTk24S+RwahGsMloejM2W9Y+v62Uye/8zfOGiSLxYGKIAHGB
JDlOwTgqNsMzUoMbacf3cCFhx+c3W++3s0p66LxU9eLuO8sEO9l1fAA4yjjC
fvoWcRZPSosAFPeBRPpvCU9WiMQpprgD95ayLuWfohlBTGRcOK13gxBznX2n
unu33CZGOLr2E8qvMvyFpZsFZD1llqaN8USwEMMS1drAxahwvxRPpHzzJ2ak
4PQAmW5oATfTx0I5AhHPXP8IeLkKZuFnPx4vsCVCdNKLHn9L/BGAO7Ok/SDx
d3wopSHcq6bJMdVo92xaVeI3k6kgJdJxTSH/w6QZl+iPw8IC+nBOvvcB0D7/
bTu1jOX8xOUdUbCPrFRpVpzY3OS997GMtg8F9ZjAEmwd8yEff8m2G3fj8+jS
O+3CxsmlKIW8Kg1DACLBhGDzExi0iaQ+c327NEz3THooi4ZWTNWu37aFVmhq
l21rQMn4RDZRQrao8Mt59lZ9LFk8dXdkv6fISJlEcsxq3cE5hz4QEMojjesY
gql49VMD3D2ZQWhtGXneqZk62swJFDYLEGMC6VKwd8LfVgbfQhzANwZtQuKW
CpTCgX3djWmJLBe+KMyJmFAP7lxfvHigtTh1GG/cEcan7oTkS8EF0t/axUQr
p4Rd4m5vrcKfGEP5lwmeK2GpSRe3zJOzhA4nI0H4hKp0A6PgcxRje0nvPX0F
Wkgz/bghUmacS+HgiruUFCIDfp2Jv4jKROv+FrpH2vpdUmMdBsG3oumuEfWt
wiKQwbUqfswGiW45ncDeIbh4EjGAtH/JARKWImRa48eZJJC6c15Sx3iaSe7F
/G8gvC1UzV9Zo6PfGzTZfkdvrJ8kWxF36vwwox1MxVQjHG4ft5rVhjiul2xZ
HbHiRrNAa+zyhCCaqxnNxmGZY3JzLibgK2Tiq8jq6rOXEyqlnp8CnL48EUat
hQYj1Q3BvK9tmOl0eKHNFuMz1YujNiAyOQB/28+tvKDBuO6iXNnhvtud6lOn
rNSuMKICofev6h8p03YNcLaXFyjt+J6rPMeAq/WtDFB+DeNWfw0Dn9yGyMvV
72VdeGn+Ice4w7sQdF4jfXMQOLosoF8YZYdsUxZXnhNb1nqCs/ZNRmSt8OFR
wXv4xA4yry5ulB1rDXEc61ZyqPy2xEyBANapmtBNzH5k8sc7VNFQiUjEgx5f
XEa6NViee7I2UTpgsRFxYp/T0kBr8iejIgdWEm+TD+WKroAYkeHAx9I65dEs
Ewy/oRKPenHRobYdXx1OKljC119aOpu3ooUdZgWMkiiSqX04x0r3oDTBw8Di
Kvlo5lK1XhQkmMfpRqvCWd2oW8GBaWbKuDt+Bv/u2zS17HB3RqE6fHk+9owy
0HIj5s+QIxb2z1Zy01pB9QSKX7uT8x/FjOJSyZwWL5BpeLl3ciKlZjQbL8wE
caFMjgGz9X5PU5uSlQ6Q2HVKuCe8IVS6EQLYm1kBY1klaKWGt3t+z4SH60HZ
kGfqoGQ3lPdpuxyS+4DJ1VLw4AWyy5LODAgr1r6BlKNa5467tdOGBOBj03ie
2kVh3p971M4bhnCSVL4gjE4Y781apRjBDl/FdMp15cqAnmUEAvOUtCWIo1Gr
Ov5VCkVykM98NGP/93Ka/KSlLLwBMRu9rBiGD50+CSMtX+BJ0V6rar4s4t2C
xw3OiRaSxe1X0xbdNIWUAA7z3lacAGB2cuXkaS7V453oYT8N0UG3MOVZGGqU
oxf8d7eRdUdHc2dqfj1gP4dhxWfNHYsyEfj2otl9AyU3RHAoZGz7wHmJZFBi
fhvSMatoqWnYcblBHl6lnwW6kzkJdkZl0Sc6QFX7uiI66MW3QcdRVJjUud1N
Oftbp+KxqoaMytdzbydfo1KV8ugd3PS6llOZAF8QuJ9OE7BekCzN4Rhs5pme
cZ/PVI5Lb+YbIkQilrA2nNPK+9NigckoYGcAzIHVcneXrHumT/xPns1haojv
k2Y+sOrtPdkLkCdwAU9n5N1hd0ZfRVm61DifsHE3sLZpzHBiKStrtEsnhuVy
NmU8JMtGAQYmFoakKX+KQ+XViXANrrrDyePVdRsVIMHxctXivwZcih5FXaVE
lb4lcdVCzjr/w/CtrAG2PCCrQFXs4gyX/nv9OdztXnH4++Y6LsB3vghqddG5
pYgaEaPgkz4wWvcah86K4VdHlqHKfKJbUdh7QMatPjBgc3cm8ddmSGjhFDW6
dIQno9v+vM1AP8fAf0fjByqCVr1cgIEIZgeCvCHMxF1asuC5oF8u8pTm+mEL
/ptMzOhhLoYa9KZOdN7Dc3hJlBf5jfzb01O3AYdS3LPIcRj0zEmZ2elMZ7tf
+EwAZPbRkBSsumfedkbP2V2h/KshOMyKRjIPrnQ6HW4/G5bOuQ9RLli9rocd
2ajKuf2OP8Uk0QRfpUvt5SvrGR9DpbQc1mbxev9UcKaHG0qwBZ3iyKEa43en
bWNPUOlHBeLoYyISi6WLywtC/w+p9vCQwHkaSJ3r9RGUjpJJ6bBrEhXUSBvY
zRVyinI6lLxONiRYArVY/RYwoF9krvgTN5Sxx6NIYCs5luebOTDw6IDFXrS+
GKSnYKXoPAwy10hGoWqCeEa9lFgWCfaZB6V/wHpyCqhByYrnhYxMzWZ+GKGZ
DJmT8Lo+hbg+OFd3+qG8Q+5RPiB7Qz1wzZpk3rwovMM6cv3e8dtHG+bLPg05
jlUGRqI53lHOKEuF4IStjF3Vipuf+1uJ/LVcNoKsDD2oihwrv+V4q7AJtmFd
oQ7shs/2SGKzr3AV1mfAuksSmGqeC4eD8cmPTrcqGsX838g+c9qswBNB+V1F
0VwvXgADpRlysm1/4XN8h0fjm0PxqjeHslCBOeMKL+imhp0OwnRyc2vPQ/Mw
g44SALGc4P7eaSsdOn5UGgqb2AvQDXQ2Pk5TQuRUtQ6JuYM+VHogOpVThnLs
wq5z/qdbPCHOnP44oeEltZ+7j7cc9w5u4egFXfY72Ns61ZZVtatxBVySLmUP
3ocBcxtV7XkOzQhO9PZaJOP6UXqTaQla0QpQ5BhIzZWfffkUj8JuVy4x51Q4
Lyqs8zib5V/EdfMjLxC8toWaQgE9cMyguJtFu5JQQPqoQRK5vk8xfVHZaX88
16gYeW9HxJByR8K6Sp/g0MCUgglB5EeKc79HTKefSJtUjepM5yV317RzRQ4S
kseyYftELawD6r6X8zYGNjiYWMc/oeTCECuW5thF0t2zm0mHuZDWTu4W22vv
V7Xyd/rT5ifQ1WZyvXCUN1i47Z76IncVvm7PxZtKfCg/3ZnDhypnK3QavTm+
RxPcEY6/D6Di9YUFWi/O4eDNDEZ7trW4zJuDZcB8wKqvdhgeuwSU+cE73Q/i
16Pumm4S+g+wRJ2B30Pe5lY/KqTICi+dEkyidS8kkkYAWzke5VgeLhTnDCla
3mVz3MMkLlogtR75/goly37PvRA3z3yBqW/cPde4Wq+IL/fHBl4ZvTgMVikT
Dd2jfiS2du3zlo+aVUyCtykvPo4c8gyRO8Sl/P53/Eym9v9RWJmNOxwdyuOt
Pt4cBeUrh7KgbUufX3Wbxz5rIHwVl+WTB7y/08+IFPdymBiFIrBV260OMNq1
ARCLt7ENGr4ZP4ZFPQEgSEex76582Aitn52huf+phFP7oqOq4eAKQU+wafIS
F9/FndvhVktVaqmef4fdh0FZd+Ah2xu/LZm0Kxj/fdlYr2zJjjjrn3FT/5OW
z+mDEnhlp92MLkY5Jps0qc0luqFK5ZAvzKqVmbxKpB9OIXIO9uIJhtKoywBJ
qU+Dpn/qKe+BmT1k80FRhqNhpemdKQiKwPYTvKHKdjarxaWZfixH5FkeGvDc
4M4p3lLZA47/iq4ovvLbGgRUw98mjAR+3MtoBFUdq/TDqSwp9VaOsbxQx/dw
0C9bsQEzmYo8QVel1ncVfqBH55bry5FdBh7bL2mMgYjG+Or4cdC+P+QJjH72
T38DDIwYWCIycZLy25c4aKCOnlTNrY/KJAwe/y1DDy9Pod1GSM3ezFfr42Xs
i8gZkf2sB7PbIbyis2poF/yjw5WORfxuUZ8gnK9jX8uCU3dQlRG4iQQKnvxd
eSk5owUCistpZvZOM9Ll5hek0WhdFI7lsL6YN4ebP3bhrQrK/5reP0AuEGaM
3HLciu25SRoJBnKN0wg6dWqvNXpcc31ScbpZMV/HjkCU911+d2PetqOOYqfr
6n7uiajLRfTo0D/PC4W+4G9FFfYkwBnfqzhGwkm8uWpudpcEL/L09zl66rd5
zK0MWddV9jPBALV24OGpmGn3ejqlxAakGMT5FMBav/d5FwJulrqp69+jKQtf
YcPsCE0mkbZsBfUhTJDx4r9iaMUXy4njgrHYk7g6TPu1w+nEBA1xOgKE0x2r
I0NgamHZl3UYuHbsuDqnOszShqVm6FpFK3o2+KoDLz27UL4vV6TmjYhtvx87
H10MQr9mwLTzS4MD066mNwjj5STVNqm3urmErs5KNwIUnlH8n5sDsRQo37kE
EeaL7Qw07G6tVel7krekPKO2yljJ3nCkSaLkK8Yz4i3LAH61hlwaQuTXunEV
k3/nvDZGnyWIGwxDbIec87civfvbNYDudnOAV6PHgBqDTfovC8L3d91wYcHC
Viw/t7KvuF7qMT2ZBcH/tjPGQZSMydbjD0mj1T7WU6qPlPuOw6W5jvv/Ozen
Wsf7tktUBfq7QGy+7xG39POs9kxFQuGbM4Q2S/LX3w5GCawJwf3CeorqpiQl
09t0BIYW4hHR+rveGDMhl4tyzd2IFhBWovGoESKwZgoVrbhs0w5iFUembJsr
ldnxTKG2BUNdD1I220B0g6hhA0vAVMDxchvP8hWAqpb2FOvxZDiGvujQTFPH
RnAgRmvT96XdNSDpmAxCJaLgWw1W2V8Bt1Om0Vu2dmIcs9rJaFta3+et2111
cVEVn7areAkVftqFTjqYw38PgTbZqRaJUGpSQRpQlFT+hstilE6OVJwtJtvs
GkdIcxmv1Q3m9oX+z4wQ22x4bq0D9V3gE7RcavFPreyCEqhNq3svUTrqd/3X
sA6EqS/m73UXO5/+vsPQfEFM/NVAJw6Q3OEpBgxcJi4ptlYe5ydahn4EdQEL
vIDq0drJE2WirG10h/eFqccMLttK5kpQbM2cv4cgN+Pu8avlY786BPIZPmSi
pa4lf5btrtrLxhTbQMxvFhUDzUjtvkp+z0WQ6JFzA0CQEmNpYQw5ySDIZvak
fz92rKfrBFW9fIsPs85iY9lnNSUUXHXWgBqBYfOM1veQigTMo0OvnLc4DwIf
RJxwYagXIdRlZOgfLFM0S94qpDs/0PB7fntJNrGbc6KJI6+oXHtOR+InAYd/
uuwOUpafQ61K3bNv6PzRX8Tw+giNJmAAtyKY6HqBBqMMbeQeGFeK+cXdpk+R
ixzHQ2tHBA3h9AcRKociAHzqrNWhHr5pHZyWVS+CmqtnyXgcVytCrc9b+6vF
qDDCbu0boIsEJNSnGhQYqS9v4aOrwPRtNpbyCgOJk4qK3H2sRmiMyGZpTP5z
RfCVE+jmGFivxZE3MLg0gCyczKlWKfsGFNU+VVEWfXSpphntPKbPPkA9fBSP
JNp4GkexOwB5f4XqBYED52bi9g9dAeIsMvTaK9rn3UoeI1PQ6eEKAKUTRLwQ
zMdQQPP72K+ncX4XwrYeQJw1vK5KorzeHjZxCwlxvWgWPVJyu2LazBdTVpev
JyqqzdCBnUnWjLUbt5K5plh95cJqS6L3/oqDmubyNbom5L1c0tfozl8aMrci
I7oNpU3BWjpNVsAGnjNCcYem0215Y65IDUyZjDhnIU6/IdDB1DL8MqSxstT8
XWP1XXjh0f1EC6cnWJuYj+Y7Dz92/w0+2DYeCEfCFWumUW53jmQITgz4CSsj
vu2BUHloUx8/CZU6jOm6scyki83jB5kG2txGuIQV0wDm8Q319MCQpWGzGeJQ
UwJMCRueo8KzjuB10sYk1lSVgj7gDUrZ1KXQcz1N34vY60tNygIL8g/OjG98
bPEQNfU6d19Dnm6AtwobHo+05LS/WFaZqqTXnGuxTKr98+IXLb3Wx5s9od0/
K5EcmoSzDtLxYdbiU5bnwCSbP2SfJMoBrSLOL5Ckbx0JBCO79HFQhttCedMM
sKHbmusI9gsRfHNnb1IYdE8eSFg4BFpoy6xXO6cY8pJaNombnOZAAPj2F5HU
8fzPxcIEBLojh1WPGRtlDtSSZ+uWEZkK2b+f6OgktRUHjAeeI3CAIJIZPbZB
Aor9z3fkcDUgRUq0v5Cbi7XBoe9lMyYs4HkC4+HKvSmrO8ylMZG5ReocH49t
DYh2onl4ccRIIrN1feBJ+GWM7kGVoICiiMA60QC1deVcOkAV9lZgJ/F04lpz
RpiDWvE5YrC1GYRFCf1m0W7TVJlcAQ75uWkF8Z3C2SLrULdZeYCtVPoQWMg3
PtfRUlepKgKXg10Db+S7lmwVlSrqr4r9nfoOPhYKSjXuEBsgk70oXsJ3flI+
nzOE7WlfWuv+1l+QpHeq2cvDZigkK7w2KI5exD8fzROfAiL3lr9r1f1e+BN5
ITtHJ247dswE0Z1yHPxBxMaOIFOL1aSdylkrJntjdLyTHFZNLEpgfKkuRhRW
IN6C3V0U6d2DMIdLkl7R12mB0g8p67EdU3sgZ33fYA5td5qRS8oOHq3Zqhpk
KeW6q9XpE7NSvWPNd4JthctHWoYxNjj0maQ1d6gXchSNcTI3d5ADZA3810/G
YfAtTJDs9D+XFnrQJDwJgUHlyGikHUhBKm6aM5yjiRJ62ChrXnQawnCquPgB
JWQCg2wR5nz+Kx3sD4X3e/OteOFWYe6Kd0VZgTstcmCb9xgkICoabGNQNfm4
fuLqUfkPZoec8eXfQAnOwzjg9qaeK8SISUgkvYeddGp69pAIpdJ3WdXPx20F
wAQkNt71fOu7ior990Hu2SU40f5xfPXqzlo0PgdKT00J/qnfEZmMHo63fwp0
7xWJB4j0xyw9le869tW+cEcZtOb6rPz2k2d38XUmo9aAeUTJoX+4hv/OQ9t8
oiCWqDwVV/l+vVxsVE44Ej8KfS3ecXeSNO+bHtDA7uCIZTv3NIdMOEcQn730
0PE6dm25pBp5MeOwT2XFP16toahIgJelapf3HJEBWefhE102e/cY3QP26xCJ
dKqgNONeSah/7EAtlw6/+00oYsq05qXiM7Vp2nSwHv7IfI+A76TgOz6/IyD5
RhRuIgradanA6fQvIfzXwjbcQ/FVr+wmeyxXNe2HTXA5jCtcXOlvYbTlvWAH
k+qvbGRapdJJfcVDuEF00N7nqzDAtABXYHrppdoHJ1GnAKW1A2sNnPSd7rus
ihSUBArAA8Gr8+hv1LHSmhpakBbY8LmbvOdIdu5rJO6vvQhRiHA0eiHlNAXn
hw3vIqoJE8N9ZeyT1ylh17yjvjH7laxDVicAW+K42fnwH+CWQXjF97X4HREO
mJPtYi+R0exfVtmxR0zX28XI3lLhsmtWr1Pb+Qyw76qfsiznqP8AvieT/knM
qOv0WR2kyUGyc0UnFpPheNQ1UmTX7WY4NCXGF7AxbvgjtYqzXn+hf2WQX5lx
GitOsl88kKTysPjoXmzp1c6LMalRXmyRoJYOMkxrO1bWjmSVWwkAmnjcZtQ1
TH6R62B+TF20OA3vWtz8THz0RevzgQ2JDuf7hyjQzfev9BAiYKHANgWT6jJW
ZuKuRZI5Wbswugnq27fOdcCpRHkWvRMccC6obFTZkUHtEBTbbPTjTQD6kNAO
twBweWQHL5W2QekTbAMmPyQkuOg+ndvvqM4Ucnl4Mx1YZZ4942o/U3GwEH3V
Jggl+ScswZ0/fbFe0wffJA+WufqWeZ7WCEZ46wmOOebqet2lMpVIC+BiD/gX
lvGC8rXE6pSyXAXwfmITfIloztEjeTZCd1RmPXo1Vs2Wr61tHwCtFcT6l84E
6NXkW4tnHDEpSbtQJUo5CMxtOOTB7Ic6EpwqeseYDYd73Ld9P1ahtFcfcENZ
acXo9Lii+qZaJCf9w6X+pfg9Kp/MVJbgNpWlpgGUdPu8SPGaYfohil+wgPZR
ccsobY80kOyBNfIwtP5IYth8Xndi0sZkocWYe7i+5Kfqf8bn0RjtHz1dO/WU
6JkXObbONgHFYS/gkVj0YMsCvxFbcQGxzY3CeniDd2iyPnqGL2BEfub101o7
MYAA8GIBPKv6zHb7hGIvIdBpQg+dSMTstYdl0//Bsn8djjNIifG2tVaA4MfI
ZvDIMmD1TMFrjTzogijyK5yXB72WFMMyDcHlO3Q+AnqQLNyVrxLf22vXGq+M
6gFTL6AF7UW71jKiha2U3yJb0Uqf4OORie3Ia1Yxw7/Lul1Vh0HwWfkivw0F
0SKOdRm1gaTcXay7qEOIXiFJkJNGMxAdclPA3roQdOxsQmSUgd1t++Qid6kt
kFC2ntkpyA9/WjZ2e/j2DdWIj6jL9/IXcmRZ4tQ0caUYkG4G3xr03m1WoQr9
xC0ywZcFPkKs5TxbROAlKNJHJNxTZPP5ZR5Mmti0Sl4AQjc2Gjkp5x4ITwQE
EOYZTjJGCdnA0zYeDsw0VEJcVYxMhd3VvJ0RSQ6dU872Y/AivG1GjiXDzAiV
VhLASALgVzRUSpuOiTZ5V/CGMB1o6ayGhuuV9gEDSLi0x1nDJ4NssKgYPN55
IqTZbrZUFlzEp+NAjzUGdMBYQ9D2DKcwwX7yZu9shnVPHkgBAjRsviMTVu1t
Fph3uGzgi7i5+OmXyi7LGCpM/JHp5zZQyfOgXCL+yJ3tUGlicTL8jROxxMM1
8vrmK6adx9fmxzuBu2VdFXEMPvU73SwtgeV7uXyg/LPLKOK882tHHqpm8jLC
oZF07A3f67eeBe9owf4mQEPtj9AohoGn1Uj4/mZseFwOyE8fHcWrdnMAbalo
b5bG4uQnBxudsbia+dRDXvMsgPE2ZiJWe4aefoKhzYtF3LF209Lx5FScvXXS
ofv2fR5eX2r+A0dU+4zgvOrxRBV2z0SsnLymeW7lBhv+AvA+UjR7ShZZeS09
LNW13pV/3vp3Ph8A6JWxTLbnuEQsx2/jLkbL63treOOlDK/V2Z6hHx3Swx9b
HqTLUJLa96NquafoVr9zOvYMAlfJxSn9bqnq41Gb2gD7L8hw4iI+Kd22QAuk
j2Jl0YKjHAoILOJvMQwfhp0dKVCSqN5eq/a6UbcL8vUWZ2ZtICaviA0dldtk
CgSARtSmQpuvxOm8HmphMSEiGVciEQGPO81T42HtDl8A/Pq1Pujzh/DuNzNO
lcPMEAQVh1/aW+Pl0MWKMz1FUepD91iOt+etkw7SqhckAplGwi95EhMyNrtw
tYmPDFXCOgb93TMOTUHgPirldTdegJkYGwbOZZHILP3pRO9m0BcpjdZCQoOT
xDKYCA3QzlMlDRWV+A8sxuBvPHQ9SQHaWuYh097hdo/CBrr/f3S+c//B9KmT
Fj7B44A0yJpdk9GbH/OLMml40IMan22Qikpm8/fvXmVo3FeVM11zVHrziufJ
iRL0oBBSOHzjS4kMoWIevrZZl6Xf5fz0vDM4mMtR9OdyCPqRI3QhUrpRVDkt
4zZEE3gIxYPiC4GyvcEuZQgfXnV35mPlLJtDh3rBSZNCWdGPzsl+Iy20bLvC
dZqRH3LRFnybsmp10SYBJyQlJZwKSNgwshnwld1vTirFXDSVubAtdopHZDiL
Us08DEt2u5nmWHiR0b2kMo0GdTMmQP56KR//TZYRH1qwtFrfiiZnI6QPjWM/
2fiH/iIRQCz2H6sL+MplJ4AGGmmbJLgPls0tc3tUuTQiiLjipFMXlIdnw5bo
fkF4casQV1iguvbhnf7lTxq/mVLzDsV71FhVUlPFw3fG8AQquwod+gzIPE7+
ei4SLFpV4uzTnNDwXgaBgpJANSOrsOWRe8xXkOtt6BVrAAcmzI7m5verhDx+
UVbvEoida6IMMZ3SOosKe9hNaw9AbSDwD0jxYdVhwxB2PCB7r4eqLFHBZK/n
WO369dhdPEiLH50TJ69IFM4b+K+woq5rbG25ypmLFXjCdmIU4XqIB5l/crMY
qnkw50fWUC1fsMZ3DfsHwEvxeGZ4cLqA+AWPBiTfJgkUe79CKw1vdK2kHi05
62kjq8OnQw4oOAfUx446pVxG1pAwqu23mzG/ii0gAtCwOOzwReiR9J/9WO+1
EWW9UNxDzI7/8ElKlG1miY9HURvtEDhWybse3ybIF7+zbBXlnA2jQKT8GchX
nFxQJzKTqno2YI++1U9O9vyN4wnTHagtouVRwwR7ZiOMPRaAc354EXPX3mP2
EsbbqFKvF1UwxTvpFUdecwfGc+6NyizumMZ163hoIyDpazpEarQibeLGexJI
pLDZmjeP0EBCPRLUFq1MsZC/9Fo52FI+hDJU3ErfqvYiMni1FIiYZMTEjjFu
mVXMHYh3km4RbKx7mX8X4p/IP1NWsbgqwfl6wZAuzy1eKpYM4wh7vIWvkeId
YZyMNUsp+1rG6aR9zvT7ta1dl9nTmZf3zuVew5kzUd2zB2K6nNN17EjJDMqF
B1iMb8nqqtcdJFCjd0yCzy6Rbpm7G5sSbxx2Oz81gZU8kRBS3ZhTGLHOILJw
L4tawtJv/E6D7Kc31Ti04ZpcEp9d23YYt3nJOOYjCs77Aj4Wfj9Wa5OF5Tti
d0udYMqQ9JNuUqUMeOMtF2JEC8+K11gxJguCkONSzjHGGm3IEWEfF5Y5f2B0
L1M+H7MnKuRin++f+pffOO/Dhm6nLsYiVVLsLm3u+neNt6oqVaDvQmoTFHY0
vH0LDQu/NqSVQvfXuhBfBUCxmGRgAa8lfrTLnGly/ZbS6UcDLoN2A5Hd/lqs
oqANxMw0y1A1unxRCFbXd/QX+0ybmeHKAq70ZStrt/ALtUz/LgfHKRkFNQx0
xo9qcGko3vz+SqfS0rv5ceU8XKxGGympTXZQ/8WZfkKNliKR+hitf4//wV2m
0xGZ6Q9EKJeqZh3i0s5sSmHCx+BbDQS1J35rleayQQv7KQopUwf7QrXTeBiW
58/FnR+ILMVCuWzJwppUZF/NnIWFHzzom9qusY0BfW0Mq5SoskVYMIXb0ygM
VrVIC8lJLN5+u2FmIzEHvWtMs4JTTsF4eeWcp0fPggQofxrgMLVzGOQ8Mrct
TUZ4M1ulxD9nEnuBdHwwjIFU2GqgIirVsbD9y4dlzs/Qmza2NSajkpCBDDFa
+SjQGlOSVd9VYQBkE3nS33sSd8Ec+adckmYNYK/mDEKss2H3OJzZYFsCwpA5
w6vPppRmSnIwAyg0C126LGTSmdd6wAJUVFRByQD/kRf23Kt5P3hes9mP8poi
EcwrLYw2cTE0AF6uBDxHDX+KgPKfNUxc1AaIFaZUzSoGEMyMSAh07gp53sd4
bB/WSzCS60W6NMrN8hu8cT5wK7cX7kr6TlQlIfLd7oKXQx/e8LEJzp7QT5/1
uWd/QmP1nbjbO4ZcYkJzuZiC2aSGV0S6sCDN7/joGLPEsiRyXVYPYdw9yzEE
/J4cAkoB+Sew3azirRhx41KEt8liQralMw7PiGWvm1vAdXhfdVGWmip93+c1
vR0T3c7uhayqJyifLrnXV5tTIXLJVz4gbk096q/MkAAX5MBgi0arpspePaB6
YYN12BCey8+tBDIVuj+o5+7E/cJu4FL52neavcwxSd0McShKuRyUalVuEPrH
KgKwqZ+EYmD7d3//dj/b1utuDrMXrujCMz6Ij8qXjoS8RclKJaynZm6fwvzg
F/arXs82K/TiUU8Eim+trqfWIbTXjI87jlOOEa4DOGw/jq7JgEEk9vbbeL5K
3YBsLBFeNXE2oF1fou07sZeTYGfJGO2q0byI3+0YIx0rWK8S7k4xg19szBQs
IrgagbrWFEOmenQzO5nMqc9XgPkMRx0LEuCFxFbddp0ziufCOKFXYa4DdcwZ
M4wuZDgLNLm5nMZuaDwbYqB2mxFQP7DdiwRBoxV5qGFecLj20bOf4a9xA2I2
8gWhiYldKpgfI1LSm+idAALDuz3dImrOMc1e50e+FPJYnAyY6hOqinQkM8uY
NLRyn+uVIF3JEVAFRZEpWOoeZ+lKRAt2uio21UGBz6J8Lubtx2uLn8ScMHL7
6jIa5F7D7OwFt8ZxK4SHj9DhvJN7E8tBD5hB7QRZmxKniir+gMicgQQHNakV
cxoi2yaViXs6KlghW3dqnGu4nZtsSlyI+ZYICM6Dq5IHx9+6JqLv4Tx0CIig
PBkIsX7xRHFo1R3Qf2gGITHmpc2RrHpwmi0A/So2XhRzxetOXVzp3aUAa55d
jXKWvcHPOCx5ieap7iGjRtkFwYWqScurtbEslxsjTRJBOctEuCXAONRspEIX
e6OaQNs5cJF85NG2CoJV53XGmq+rf9ePQTsFJM6J3A3BKOUQXASHjnWeLF6Z
H67WSF4M+VOEsts05qR1M81F6mm/1O2ue5iSUen8cMj3hv0OIKB5GpMpYbqX
O6b+kOFMWJLsZfL5LD7EnvsW9sW6Hu/JnnCPWN5DIWHhNZ9xI+TEzj/gAyFf
KyPgPq8iYmzzIfqul1dMqc0ZQfSeCgBRJXOeYd31Fld9lc3Rwjd7OvIEIO+F
1lgAnKZJI4gckybdZhy8DZyY6Y0d+ZD49JH0tKcJmLE+5MIH786DK32NPcCQ
vWrwsvKbgzF1ya2hI/2OyhFR6JoJvIWEWy6Dwjdok54ZHGCJ9iiMhGWQ5EhD
wa0Q10V5DAgr7qiNI2MMwfgYvrsvdiPogIgJuGed5y6FAL44ksTuKkoUPx51
AexCzy+KbFPUfpnSfSdywB0wmi2T9gGS+YYx05p6QPqkIkF0cSeCskNakdH/
1nIvsKDklegflKsD+mqe9Rs+BO6zpHAeeMc+KUPLl87MKxsgJU6coCLBmbV8
ajJ1hBPuXHlW4xWJv8hzB0v/XnKY1q6d45EkV0es0Ok2VKXqPk9B2xF6ZBUb
851Nt2yxbiaJy9cwC2/SuvPZ8VsQiI3O3FMPml6skM5sSafACSp+nPGsV548
9Yl8cpdG4CzmzE8be+lyvilRdEw5scWIa2TBrxDzUq5ifoi3yWmxZeKJ+AKN
9T2YZ8lrSeCiua4ih+UAtRgVPYBXvaaXpqkiNR1uNX7bvf6WZqdd9u1KR7rT
6Nj4Git4tbt8YR469VCBCKV/i1HwaTuBYD3Ldg+zHQK+xiVnCTnTGsW2VENm
zQ3ac60emc5Vs9JyKnfxZ3+4vwdeskhAwAXOkYn9F20DzdvPhxT0ouhzVUs4
RgnK/BXz+rA4uWMgM/q3ao449KBCRMUfG622P9l87pBHyxchKporRkd1Jify
fqKnWn4M/PfXyo/b2LHi0ctrSL0yr6v0HQYNsuw2Op0QW9g66U6VIzbu1zgW
Tmrhz7xOO0j0D8Mced5b8TvVmkgzpmxh/jz4T7MuATVGIYj4tKx4MgWEvfsX
1E84YRxh/Mm1EpLhH7UF8wkcWuDREmXsGeTkwnFHyJ5l2XsdFUdA4qNXPP3Y
22JRuAUI+u09BI5E6U5vf0frv/cfCa2Qm4W6HSqN6Qu3gfXT9B0wjmsBHCQx
cvx8uyBH8uSDNyCRWymA7ZxAdny8oQe9p3Y0h1LbX0m27zFEDMpPn7EZSimW
OJVse/jSffQOHGs3oN46D3LuFDsgG540lTqg9xEnQ9Qbwc6VDVqf9075QJ6H
KtPukmomTcGIAEIhf9Y1XqO5vQrTR8CMOC8BzuVHllKd+B8b6fEdkBmUPchF
u4MUrM4tTj4TguUS0Ks2FqyllgeVFnOJJ28+GRLz1xGWQC3y2rooDEM7EhQp
YD/i1AjDsS0Rms9NPYYlkd7065j4iCGSCFW13rlaoBSTx3cRhbJWvuUDVPPW
4WrBaPkcC5TuohWkmSTWbHdmEQdTpbKtUI2kP8C1yLoBDlv0if6UFf3QDsff
v693lRpHLuoPwY99kUJOAUDhBXDSErrQPCoeqk12ChSQDcpUDmnKT0E+WFHj
+Wa4M5Pc3fhdjkP92wq/JKhepFLlwoxJMR8fjAgQ1EiFS0qccbxjeMRHpC+5
XwNOyB0HoAq++4NenrBK1IqzXTWgupuEQj80Wk0ks0KnhZQ8ynX1ZmVArjJi
aZNrJUCsCbs3SEKZixptXTvIXegbRDbd80uBBV4/0E8ahCx6uK1TH9cMt5jh
1ai2EuhewPjfxMl+m6Zin9ElbtFkBV59/hZhFy0pq+eP6ijObRANr0cXglt3
JnD5GQ+bOHnjH18aQG6A7GgicQmkNjXDj8Y/Iltm7LmoTzhKJVlXMzkX5ylc
2u7VPMk4l54gjgw2WZJsm1w+qspYWWURGFxKpF0KmwdZZmXwEQxCzBjVFePN
uuEqBhmgEM+FTOWFEwMNsiiTMijen2NObggTCVwU1tmncB8GhH7H6SeQPcsh
CpEwZnk8BrkLXAJYovYyHgJXFDjrJ029bXEjAx63IT65eZl8Sw3/7ePPicAn
0INhlLGOWs7JfJX7io+IVrF9CVfueH7o3xqp9sZg4s4X8Uz/6zACMMb8ib9e
hV3Vf1+vs79fxIv3xQnLTpF1JVIBoelQ4N70wGHzl9bZIiKdCXdCFVgP2zDP
wZ8M4g/MUqo1p9D7UuSlxRWpsyTqqi1j4On4r5SERLHKfRVG1XCGPJY9UlqX
jj8MXPPm4fyIpQyA7DJ9sztnSREH5gm7qUbm7tXeMu+Wj8LsfGbJA5ihHp4y
dh58EOsl5CsFPeGacYKAuE+Vw29OuV0iFMCv/Q3zn2C/IPDD+bQQkJ2fPLui
eGlAmGtNzgrJ05XXl826mi2ajs1IsfpD20Z7kiVMnglBLGVbw3Rv4bmEEJlV
ogaDy7UgEJycMqsrr/vemt2eLxf2f+skhFLflnGSPm6NJLzIwM9YY+Pgfliy
/tjASgzpvtUg5IyWPoQZrAsmhuay2d5ETE174TvRaQtYj1Z1p6O+P/vsKVFY
NUVvK0XfrTvLNRu/4BcEY89WHETy/BcBPGadMs0Gd/NsjJgWqN3Eyu7qAvC6
WA5hz88klmGFbG8guNjyT/56qtTTEnFZbYReRqIw1vUIYypsfepEsz1MfbXQ
IDvUch5gW2ru2mPlY+4idiZE2071zWwvUH7cl643tQ/iR6UV5h9H24BTJjrH
TSv0PIJmIgS8bB/g7Yzt4CDyFpTeYV8R8RBOsDouOUwLMcHmk+f3rSGZ7Jts
p62o6URB+bYR3NFOZNkVe4eI86YYdsjszLds8HYkhxuYM2NgNOd0pHdCsGPG
AkZSqyykwrWD5YdFBSzDQjQ+6VYwM3mXCtwQz66Z3Zrux7Hzu3PXaRLk6PVn
GCy5kD4Bl9uBvrsy0p8E/ZXTmkrpqqhvEGmpuZi51kNzFmw4g1sb3CKcYWe4
UOT4zwuaxV9p2fBPIx/FWuSOXiCJUrrctb56DwHV/psUjr4z1Qrg72Cvd4gF
qYEwWl6cigR73nheXwvdeYcm8NE/Kapz6FxGHCclsg1mOIsxDCU+SE60ymof
KtMtG2/9Zr9ozeYdxWjM05BtE6ZBrwmIVrLmb0D47UMjgWRKiZGUXsuVuw6s
XHHJ07yUVEfZLUINWJFQN3WqJYNOBiAKraFe1R35YLCAQ2cIqjH5N7+7ZmSA
iVnrAyVmA4e5Izt6YbmZ529Mj54YefnFAawrIqAzsSsY5w+X/9Lik9RueyLc
ZM8URwJvsvDNgk/dtELMbiWoii54L3m3NTdFeNUrxyJdQe8wZisCpQMNX0Jt
xHH0w5eHTQxguC20D6MNpzdDrJiQqVbSKXxLsPo1RgRtVEqc0dgF4mNCl/oO
VOM8JcmgenmgPpmLo/X0EeKiLk+VZbG+5oQ/EZvzoYXSrInqlEWRJAeCZs8m
o9e0CmXoI6QivKTdLOapx9Ujec+CaQK8jBnRDJmNttRtZpEyoaWzv1tpaYQo
jghsi8YfR9v64uA08cBsar/2gWCbNkfl+zaJ49vHD09R5YP2y133JrJqzqL2
dWk2FTalD7pcbBrXJyZhXOFV3rG4rzXhBfn3B3OsR+VknIIrkx9OLyXj9IUr
M5TSUh+/baZnlZhqseeXN0Q3UAxM/A67bwPMvFIEzI/KnJMgOdlnBuag32Sk
PCF7+qkMDSBiJVFv5gfrwTFWMMwx9IN3rRTYfw3hIZx1eoTsS954DYIhCXAK
+eSNZgJVd+Psy2acoo4kIwAE64Tnf1CRJm9My1bpXgCvERZ4dbv1D3MkqHmF
wYk56pWrSGteeo7cDJpU2Aszx34mbs43FR0o4RpTQPwIPqf0P7xejTrm0OPm
ViZLNKzv3aBqn0/ti2lFVb41VluCQMGAMKFp0Tfh+UNAokbkUWb1k34lZxl7
fgmmNv2OL/Msm4JQ1qHXASzN8xlVnEnDeBI3ukI9FffmwroKT+K58Czg8k9F
vvLXogzaiuX9V1UScYFpAk6VQ9FGTZ4Z91NElg+a7t5IaTDqK02/teeEwxdd
fvzns3jc/7sRA7Pm+NDbtQxuQYSkKPs895hH9SEnQl9MmgGLiorVhW7ZNtIO
1MooELqyvv92TMyqK9MAT1eh3U3C2p4z57pPfO5u9JP2g/dG1Ds9PXL65XbJ
jiilL7prhXcfISz8iSAwq6OvME0iecmc9aBKWGm/wzXtcV/xS+BV8NGfXtMP
bAL9KZI+JmEZ1aHpVe2mouU4W1UvhVMkntBwGisbX9Ia4kxvw3SgYz0jy+Ne
W+5D60Z26Wo7A9RE9Xcr7tTKz/+OX3UWna0WbTiS7EGQS8yHcNQs7YbXfxs/
I7ytUBogXVHdO8pVKX/SeFAC4pZ8AeNOD+T31mYgR8fJ87W+3rIRLCC+3SeU
AkkQjsY7Mae+2HsS0xaU7XobpGdbq06ZFjB5191dmJLTDbUXK48mb+65VEcC
UfacpI5PNYAaxybEP1vYGOYeuYkNvoX1RCHutkiFz6s3coU192xkdTmui3mY
MLTs+0SfWlXArtnUR/WEazoI0OH+HX5lRSnJRLlGBK0biN6VWXnoO/qaBpFf
WRTKqJmpy8lfsklX+r/EgrKbKygS1kbJD7j66PHVdG9oMHePRvaPd85OeSIZ
TXeRI7sfTFRFzMGbi4Kwwbqz6w0p9BjL2diKubOknGhC503ajU06R6ZXo6xw
O6gn5jIct2mu2AUHvNpwqatbI1vNhhDLWpjkoMxTOhv6aOrV4jPgxgU02Hjr
dpaNkvcVPxm+BV27di/TMT1/rjykt4qHwtWqVxK4RCjaqNcqJ5GJ/lfvE9xD
KMs65rqjrWVaTjSVXST5RcsP4B4mF5yZJgankkqE5Lpv+woi7b3djrGS0wg8
r86HGcOL9JtxoruEnQ9P0Xojq2icvM7N80mHDLTI/iFu/dJ68sdQLdqj9JVh
49WHOQiFqbF94EELtm4EOmHJFQN9zCrZw9x1ywEyfPRhKr0cayDcS+72jvW1
bVjTHCt53t5AJt0OEw9GNc1Hz0iDcioe4av4MjcIE6T+47EmNcquoq6RUQU3
sZRa8XlhZAiH7f4KefJYrEeRf/WTNAp8B/o18KA3UYWjJQ3hx3AjngrymYUg
QZwTPH5s2I9C+jHMkhaMdvDHfHB4vFOlWP8XhjJXG1fj3DfHCiEFq5UZVXIQ
jRGE+EfEWX7Tzk3zoarx8+pjq6XVmil/1PxMn0FsyTLzAfb+L36jXa/JFDlD
ZqMmgMdrNG0Syzp1pBLs9nIrLEGVkfwHEl8AwTNr2C0uyXbSmqY+heM4J71z
n0AxDOQCzm99htgeZL27iCxT/445I81mI6Xy23zc+G7qupYhyJAx8gUIugr/
g+n3JjPQDnjdV9oCrw6/GJJteQwFB4X+Qk0ZEezDy8p85ZunXWZglsox4U+x
BiSWFVn5RqaHXclkXuDaNSNzXXnb1qR8hHQxzFoZIrocHbHRktPUyX/C/pr3
rh3bM0zjMcTg+9RZ0PBcOcugHGWhWGVleZodFJgNiPAzub47TiSra9GFGacZ
maGUcsR1KVmNNM2hA9JP8S5hTBjNMfHK1jHf6Q7yy55pkpKrZNcBWccvDlZ+
pl5mgOGB+xKqkH6qmCwuUQ/0koirsw3GYmxA9goJR6kCaQwj+2+pG5nP9fAd
AR3vQ/jHFztDFowClDipRi5UQqKiDBMTqydlvvNQ8ySRUpsUv/DJpTk/AMMb
qGe3vX76GEM0htL7N7bFvu6A9L5g0II8ZrLm77CfSizZ7wkLD/NCpeJwZWI8
NDgR/w/UiVsNz5VfdfO8yotkq/ueKtsUsMPDGAV7yOpbJX3RJG8YqfRFIneQ
niqhA9C1Jd+o+gYOjaV6p4z2gN2sgdnGCf0n7+FbruidJsoOF4QyGp2y+oM+
i+wuyJbYjn9hLHAACGr3dfGWH7NI5q0Mkw22KJgGrzLS/Oavr50sQM463XfT
mnHRJexEZbyCLj+MO2uIXvzoqsoLXfsnLtt+eF0ohoK1Z3m38M0jRK497PXQ
hJGFHprrHu/GJqLk7FDvKQ1qB9DZ2Ss+O7UmIVnpKiqK0xa0hyIG+alYW9sU
DxFGOc0mUsZaorNwsUMgFjCTb4e7kb64smYTyLWdwyKRfCma9t3GhDyUfwdh
doibpaKtY6tOL72wBybCBsI7eidy5RmUfQWs8E0gztfkTEKurxdpzzQWQLvZ
u0Y3jpE/xJIZrLMVT9oWJ86H4F2fT8nwFdvI3nXcjVAxFiEdk0Dk+oCUIqft
mEkcQ+l5wTiEHJL74L14DP3QwwBpprR6N3JA1aQ7aFpHW3A+9o8NclrZlOlr
K7g/oh2OtDqZC2uC55IoxspiHVJvIbiwri/oFvVGziID1Asc2iaZDEMcceEe
4WfSsyjMiQLMmbHVgKwOSMDzTw7Qo86Iw3ug2gq+x7hU5IqIwwjgM2Fzy/HO
C5+NuJ8ygAANsW7w0nuQZ7+KRbVEIzZT0+yrbKnWN6l/VcnaCG+SB0LjOhs3
CUqDfV9pcUH43yMiJz29qKwLofTMG8WKNP1wWea18kJ7sdE8OqoDZeCuK097
WEogsxqdc8FwLsfMMTpNZaJEOdc2V5PY4L+c9/cXeBDz76XZ5hWhMLrvjJSP
TTylNzBc5nYe7pvfvnHbllvNBJWF6SCdrD9+hUw69ojR/tjLYejlFDpb0RKV
m6VluePL2GSL3nmqbIyzMW0iBOlX6SEwkji/gddvQtY1ToXmJQ2Q4mzynBpn
g4ExpnV7nh7dtTbxv/COEIhQS4iX3bTZOoT4F633TOPy0o7Nj6V37r6P5OLX
Zlchnfky993qvhr4RPu2NaOHOWrG1GRlycuO4NYJ8GAXwi0VKsq3byoP+WpO
CzSB7CynkofDXCAY4k/Tf9qeCdqSAdYWIA0r+oMoAbkdm4XqyWP0eBndFnRz
Cq+Dff9xNQJLzbhkBPzIjp264EotF/rK4nFD+TW4D8WjLdxoTzGJqEFDvkob
52p0YqGH7go1G/MG0bf+/aCk2SM+VfZi4Q0tqW+UdGpkF6NMBsmKtgv5T6E+
pjjStygP9lOTV6UkS0mYLAkudyEUd0Ai1CdTb/UQwqGqqrOS+jbSiJpTp6SD
niNZmz/6AoCU8gn1ZJvrXbbOVv8BbaSxAXLgl4/9Xx32y6eF6iXKdJD5L6bR
R2PDZJuihfejBDCmefFIWTM2dxhEqnnhavbjjNciOwa24aSPiMZepE4jnGT2
cMpSvViOhv64H8pYry35LKAPGudZYIhz7lycKz4S1eCoL7bblDAA2UrfPmuL
6YfRGHo2++UV7i3dMMYHKQUPcdWWU255TyuBS9EBlzNz9RQNyWyg7V7JrHEa
U+SsIdKdXBVJwuPnI1dTmSMV5NKpwhTwNLlRpzvUfdseQamRzeTCXLXyUI6I
NMxieakRBvHTJk+THo5jo1NmSWUkAYiYnDChGDw1BtLIdizxhsSftE/bBzu0
ScksL6uj+5bKmsPwxK6HOOeUE5NSRTC9CAP6M3qBh1F6QfHQ2zpSt5132tlu
XW+5//IJF1blpVltHan8AXV9UdggvbbJ0cAQLSMjyeCUrz2oi2eARRzLcPnw
dLqzeLRWOuiLAt5wNAikLs8+2VevebVdJcCEvmb8mf7wSYj90vd1NAxOt4Ro
mpyE6uXaTCDH50Vx9KDrJAUcnxwiJ37rG6BJzAMTv4V9UzDaQyKILPVW0olX
IGNG9JdATVWMiUcDkBQsxrtVQrjec6AkDRLIhMsoyBlTISFKXLb3RcyXGdea
UBxxc8StN1eIPaUm5LrEpL96CSFDZHwXMS3ziNHPsrRy9AIGYS1nX8QTzbl0
DnAzKHs4KM1AhA6Hk5jmO8rL8SfNysz2z/KDeXMQgmRtoXaeC8k/Sfu4lBOe
N7C6L/TtqwuQXS9XdMKoAKetYr+RRzKCW0fwLQfrLcjqyI+O+gSWaVjrZKdJ
3UH9VjnPj42/kUnueA/KV7e13QQntmPHU3i5IC2WD9EJDRUgKE+q/P7jF0Za
HRtJ6DPoye4B1XEBidYq3LfH7WEfd41MNtdgLK0CuDAq9aA3o2kjEPiWA4SJ
QSlu1A1yBCGvuSE/7BlBV9rHT4853xLJ5GmXxf+BXkD14j7ruji5piMN//vj
w0V7hPBZfNSsNvNM5Uba3mc9YIW/ziYQTyvM0pv40+M1eQQG4L9hYc7uhZeE
4we88HRwGk17bw0xDaFEI0b3PCcaTF/DoCHZMt2Q+lLYOHTQsPz7IKGrKNXs
CHRKiAhWETYiMzW6Z/DE+vXgljxWB4opHdqAHhLzaecZ/hj5UaOEC8wt5VY9
IlOaSrG4us4R0FJqItj7kFVs00DXQv//jDbwoHcMdJ5f0Dcy0rZAYs3BJvtZ
G3QTkovQ4a+LlgfadoJGKxMXSnZayYJ0oo7N//osZA8qergZ24HdogwKQR7D
In7DzGP0g0LF+T5w91+OkZroh307VvNfXEmu5bw2Gzht3qwUZa8x9KelZJ/T
wZ0xrwN3WO3daU7sF5oq47D4lua7+1H+m0y/w4m3Z4is8Q9Gu1hqcH8lYHPV
2ZTGqJN1f2kieNgbEfQugJ+NMOnmVDo2b06rJAZ5bFC0fRPJ42TYijNyEfU3
5YZAsg6vULVPvVG4jGWB/sOxCPYwt8Du16YRiDKWDnUPpkb3MM+XPdKr9VGi
7t+I9v9ZuIujfPVg/isTtDpTU+5Q0xcOFvrTrKxQHl6ZvhG9ITkuLZR3ggiY
WAFS5lX5biojd2E1T7I+AmtHXyMSoBMPGSCWicRz3MJtlnogmBiBrC5IyoR9
oGP9tt0zvcxydZ54dD3LEKdWha26axR5Y7DrCXC8lcSLok805GvmLwLif2qP
KoJhSypspnjtDIb1D2M0bTeaKIpQuLVAgUHUpYaTz9VRcHu9LLwm72bUgZTQ
LhOwSCjuJ8lf58Cb1m2w6W80OMh1fEQckVJCIged7ZIL1NaPr3quo26+26am
wgUhNHvJE2A8vaC2zYjuikVndiiG/UkdXm4nBnyNhkXieTfVEOXsnAoyZhdO
xbiYqm0sTNhX91R9WNTSY00y65l5AqsEk+jWmlWqQb730jaoYahh4SGtdHf7
Ack7nljMtN1Cyhgjr4HItOp6nEaPAWzGRzMziu6/12zLHHeJ6uMibPDxqg==

`pragma protect end_protected
