// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
BtTmWp1GdVl0XVb84LE2Riy4MITXyzLVwWFIJDMcVTbnAt1KTcbTq4aXoQyD
kB5n6V2E9MmaLwjJkSbRe1LefAIXIGJQX3s7iRY/eJNcaG6APP+ECRfYn/xw
kfjWurUhMf2HdcCT3TTgt11JmOCobm9NXpM2XWT2UWp4mMKkCArx9ssSkCV3
Tos2MtUraf41vHp1/XrthQAIe6IbSwJ3WSGzFG+Hx88xV1VIKGTytlcHdqKp
SZNplPtIsyAGhb86z0lXmHzKOuNwMUT2sd8xKIQOsoIgXbYHkLiyeaovywuu
9ndugscS8v/GYS9MWm2ZhpAHpq7XVSblaNW31zM8vw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
p/hFSD6z+FYlUj80UmPYd7g/vPPqzhmF9GTqGMAHeQmvqX2gPIGab88dGlfA
Zo8OtIBfQFu/wiJoYxmZAUCJgXPNJoliPH+H39MXp7Rh98/i+9OGOg3/xM6N
Yn1hBKjBUGV8Ktaqfv0r2rXEv5Jlpdqx6ck6DMdPfpCtavv/iA2/yhgxE4XB
G1UqlunOWEdJFI29pXsc9Jy7sbk28lofne7pBljCbhtUQwbaTVJH8zPFlnx7
fX+Xn8SL1Y+qHGMYN4Af2nQZjj1VTk3HxJHYG9YM0IHHA63Uv3p+4JpInPD5
T+L/sHOw/GZAGbKN26LcVkcUay2mzT6LHQ/R3ZIcGA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Y5oPGQTW2jmr/oB7zFkTDA9udNxzraMn4cc/M8724VKKxUxxecKYBFMgsFmK
QHb3DBmOj8yH3MfLyP4u5Qpba0AS5rELWW1V//Dsfq03UrZ5PCI5V3jLamxY
AGR9ESAjgai8++CKxgd/WilYg+BNQXSYMmwqL7sh61wfHJJYB1YHbbg9AQ8A
OflVw6nWhb9ViDbPcsUMMIHv2YO6toz6gN64clNXeluSvYZU5AmkL/FH0ItP
nXk2QJBlmjmbetYaCJnUboCjLopby5bt0IGHFgPRoPpHVdH9fHSInS09NUm9
N6ZLgtCdkEcqPGD6Y81pNVjIlbTbCIVnMfEXfZ3ECg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
B1uRsm4Ibu8epsYn8pB4Mjq4aHqsRdZxmUhYd6KaV0t2dgEWOeokA0rMGzsM
7OEWUBe1BunN/iohfg5H/OAJiqddPhuX53CDPEIe64NQOZH8Sa9k5LrqaMSH
b+KY3ggk21Zk+s29DfxPgOxE2baj66HRj71kUNiJJMm2Tw3UYoc=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
PdXkyW+JCColoDYg6r4Ni97hMaC9ScUWrSDzjwznhBEW/LjJkrIDdsue6mPK
KnzIGSYEKokGx02iW/AcSBWKTOI7OH02mMLcMR4U6lGMu0BtGXSl31ARb/T6
Aebj2eJM6VaRS9k7cQwIxQb1BEdLV3XKI0E1bJ1kIsutT0QMgI0tharYS9+c
xXjdf+llGsu93Ut6z2JOdE98Ds5l553aAAYh3Ru7NnxcqT48BGW5LwOHBSH1
+ZTVdd0zRVYvdnuB9L/tAseMjT1H4mFpPZbHv7IlQRbvgVq6/ftfNkbPj+I3
0TYH9u39U3I/1cAaC4ubNAbzFxvRnV8vWMVh4MW7ca3KAhJhTxvnpasewNB9
vpkKCiDDa8KpweQeW+y7z0GdCAjRgZ6DODY/vOMnTyGws8RJgfIlNLF1hrJ3
NsuFX93wO1vu1ukV2PogZXd/rl8bThTJIJLVTY1EjjVIy+D3lkuHg8mZ9/a0
HJ6iei3Jsm0X3lbHKNyNGgfVFQKuCTAX


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
mAcS6XJNPInQEC9ILOu3cnOz+gwcomllFhsocnk3PeBfY2jSVMJKGwLvRdwx
T/LACQMLQecbobdjq1ya+BRnyq0CGX0L5sfUpTCjTu5xgP4we1XkjFq0itdp
XcdUcDWEJIahlgek6Et8TzjymOhus0s5+ydXjdoUL+RoIiL7VNk=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
goDrHpc01j5UpvQEbmvjUPCFj24KEY2BQVlLAlnG+7nLeI/iuAEwkqVCOCR6
1cIuo7YQxofhim6LgB9/qjC4fLRsUOzAiZRs3GmmIEHRntn1TR2KmweVKfvx
z1dw65aYRTN/iXjqCE+zNKzN5WBgTXLEdKywiuQKqEa31wP6cNw=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 13072)
`pragma protect data_block
JlQKslA7H1RTbuuaEvAE/wjFSIdYBfDB42rZRVnuxhOX+psTs0ngnKLD0BNn
OZvkAh8g7uIDfoG/7j50U/Xjkyv62RqWRMknHNl3R1qC5ux8Ff3trZTz/7Ob
jlGKtbGA6BO9WvzHGyGXOFnf4+KwiknUMbLGVIjJEkBEeVU0/20Q8BC52Fku
iGqWAluaHYcNRAYP/xcLnSAis504A9tPJmZ2vAT6YMVJUeNQLXt5w4V6h8Dp
W4nuqD9twFkiAciLDJfxAOAnvAYg1cU2kRoZQ1JHJMHqSzi+wlkMrIvy7NwI
kqRPDVA3d2V7+DL/j8SLOHXZ1P7QB8Ywb3dg2Y7KN8CuynV7TTt5kxYI24I9
S6rE6GDkERudWzbZM9hsZy62sy22P6/1/ULrna13xPMb87Jhm1GoVcz5kLaY
lxSwz8vm9gqSV97jYxjJOrdl+7KJ77MpaSrANEQ4hZUo4HV5dN2B54FijeyU
B3bJ1R+CcetJ/Hpdp7CFnMdOMEXFoPzBlYr/bWteddxWqKfH3BAiV9FCYkQG
T5uaEMptPqEkcX2vBNFZkKTuF9zNYo3mPaORJIpebSRlnZAEhdtdfxbFWG6D
TvxOFlJSLfHfjbs5IYuvN63FZlVSbGQzZwsvlOkOwWcj5bu5AuxyxkwXdcri
byx3l40npREiEYFmcLWh0qHMgiFWWf4iyox15Nq6IQ/pzTOM2GgZta5i30ze
UNLb+P2DTsCT2b2HWoPOWeMdaqP+U04hc+qq2AbZmSJ85B/uz12P9fXRBarK
VU1Pzo3Gy2oWHdpTpUzfgjSgv0P7o52SZZcYWZ2kcPz7XLfEp5s8iek4MaQ1
C4g6x4Gw1qrFL6I9ITeBwDfAdkejTXmvjUBEjzSof7FkWB/xwHQgTC0Qdotp
LKmbv9rEEiO1s8SZJnLBVUm+3ruBUZ+2DRy7at1m4DSgoQb39LsxcgAWDu4t
pNwapsBbXaEZhBiQUnqI0T6p5SaWzzLYHfgZ/3Nxtp/SCV/EUD0vnvbT3ESi
yK1SwbRMkShw+2NerKQDAgc/PMR7ht0VbkP9mi8PqWBJAuUFhw4TyJ1btjVN
B3UK76np/+CCK736Du5Kw9k4+bfzG7TKcSMegJAXxnvesd3QguPW8nENCD3c
wQ+YGRRuAg6HN4mnscIH4uicYfNJVbCYZvsfEkozy3Muj3S1WzNcg58gOuf+
9dCzbNVnSBif1UCHcqcb4wPGOxsO7kJqxvEoH1oDx4af5pQ5vNbZr0+m71Ei
TMTwvRsW++ijpuMHuoOKziBWxnVvNOsazBSdWZLHzRxxEd3zcWI/WoNcsgoj
eXpE6ipqtCxtG9RYhCh02cFonEOT7EK1pag1m/XyFIhBRE54QR0s5FSUJ1Kz
6m0/2tLe5avLIm4qnjxfCu5UTMLGQv7ABKD6Pr1L/ypftOGdtlERsFPfsZwq
04zFm2AwJCW3fB1/djrNFJkxLnvA2ez7KIZS+VaFaq/ydaDlgbaUaX+mlbj8
mYqOoNXfSk8p7J+d40s0bfzCMwV6sfJ1BEfHNfSk33Ry3kvr0m5URiTnHvkv
TVO3teKm7sVbj40XLMupM+DqXcTaP3YLRbZqBMlZN2G336BnxD/ei9LwKFL7
R3QuWbCo4YiwD6elN6twDW83szKBrauhZtCPx0O9Tb/Ht6vg7u80rOtFRMnN
rX4h+yBSnRSDQOkom8whdoP7MdYPSI/EGapB2KlkaeazwD1Q7Z3bKF0yIPUT
sWPFpehaX7/pTg8mxgBMabxw2sAPLUj+jrIF8edPtepPVOJiwIf9yhI/6DsW
6Ddy3XKhbHPQPi8j66N2V/JnTsqzvgoTaZCedmsqyh7Nn0pcvB5+grEKj6Iz
jXAkpPJSknmv1a+5kvhptrAA7atB+8VnipG0hORei7SEiOZIiShQ8Qw3lYfG
I1ujkbof4R9RMbrSohioNbRzMt3GPD7/i6Z9MwsKEfNzu0FVYKQnP06/mxgL
t5Vbkolr+d6UoFqIq3zEXEpYsfAYyxUG88uSrPDUKnn36jQ4gx5e+EQvcZft
lLN+cdA9R63r3Gd/woalY/G0fRodoP5IEQuE+W0rzruXtgLu84JEwLF1lVrI
L6JQ8wK6SXOkoORmOV30xv/Il00QNXFylLs+x7ROH9Lw2p6ptPhSz9ImkztL
dyDn+vVDEkKbgCo+y05276DT7aQ1snQAM9mBApvzMa6u0z/wklorWRuhqAeD
6ATsqBOB3FkGtQHEByDmv6kv5powUHwgcwX7dE+qFqeyaXGrUa6Gv/toIqm2
eY4wJt1B8UdCj1eUuF2RSN5p2guYhX7FZncBNLpqw2up9unvEhN7xObp87d+
9pb17Ud3sIfsySeRGu+ZSv+qhIyjuPWMgx609HfbppJUv0KXtD1T3t/G+49L
9zJZY36ohN88tnzmvIY5vlRqZAkOPTD5njbM8j5mVkA86g5+gb7WD8+NrdID
aVgTY8PbZWK9R7JrdIY2rTPBMaJKLB9DsMd0EI4akpOpZFarSsZwoLciCDwc
ebWDB4+kkMvbNZAavTd5+yCmmEqBIxS83zIcF5SoucLFzFzVxylV5CErhdXU
3QJgGxNQIbc3+MIuQRO3p/dbQgE+bJSUFL+OlbMwD/d8fPnw4HLVhmzTd/E1
v/9KJvM0fN0nyaE1r0PJqH5owcE8r1Qi1z82wW24ydeP+2xWTfzBYXSHz9hR
nPKohgn6DLGzAJai3ACzj1z7Rv4xCg4G7YMS94Fb352e+KtpUrf2XwbItws4
Kz130YUoASQ5xr5RgYGvkkMKSjfBczAP7UU3+5Q7z0KPXFoYXUmEXb7seFLE
xygfB31VtbDJ2sqdlW5/XeZnyP1crREECtWBYVMdcOTLEUCJwyjcwyA3MMpW
yooydS42Rq3xwoqKtlOHmzg8pAYaopQyw13uGBYrsO1eo2TFgH3Jquwr7cqN
aeJLdgcNqXb4FUq4J94tOKkftr/HHScFn4wAsGZ+ZmgsG/zHHbvmJpbytqD2
ZALT8mNnOvLlb2ytmmhiNmebEoc5Ueam6nM8eYMcw3ycYp6SIokjdjYyPjPQ
tEbBvfTAPRrBzyowS97l16ko388OKI878hWs5CL8xprl98Zvq1D7lszAY+ew
+kT2u9k9L6zgptQXUYV/VKwPLVJIFa/l+Cuy7MyAj9P9TXIXzr9nXP38OOUu
ByYKKVsFylumO8yaFJgN3XKCghFSbuujXf9lEjqwN2hp2DSfuGQ+xqQv2H11
K3Wcg68X7vTmLPkwD13WmRsa7uxjn2/gSI5KivZlyCEh30NhKLDw65xzl2AI
2tNV+toa04qTqrJaKu7PVWAlEzZhW6tajt8Vhk/8B5vF/F3Ju+vkG4WkcLs2
dySRd6aCikTFiKHmCffhuzU14mateLYtncHhCmcZG49zjkoB2M6UBsR25KX2
AC+jFInR6zP18ZFokxOy0IVO/w97z4fug9udDUKgK/QhPRJEq7eqeYxchH0r
zX5FDps6EEja9szVGvVIK95A3xMNDgmimLsBqRJ+aqjN9v+BWxODK6UxjK9y
BWOjE04HIKbcu186bk+pi0jYeW0wNq1Iyt2qBF6177Y1df5GHLCuC51vKQNw
eA+dKOvzb9B+9RCGFiRQvK0P3tsyD/a2MOEe4DIKkHjoM5IpjOTS+MrgYYPZ
t+ZH5PGVhaG0007YZuTTvGC+y7Wk88JH8JC4D0oXqJhvHiUiTlDtV0jgJF+2
inhTNnVvpc64eDnwYkFpFPMt1uYFW4waSK+z7DENqi16oSXmrNx59+BwUXon
mzQJVW5UYbj+daiPmEnDdIZVUT05UzZsxJkrJ8R8GOS0oNHm8Xb7oCofnbOP
jnU4NcZE4qumjeMk3q46/lzllSi61V1dj0mBTvUFWFACNvjxLYkomX5evaN9
UIc+gDP/JmsnXQ0F72hox95+dslkcNGuxReO83AADoqDnXsgZhKGXfNt/eL3
2bN4zwEvK6pc/gxdATZSVraSMa2nx6mv0lweJ4vKAHCfIWLmMye3ZW+sZhCG
OY+wPNvzMhmjxII4c9ov1OyVmfD7RMCcNvqP3vWjBi/hQF8JVxDX5/zOW1Uk
aUmv58TtxYf8DST8HeMgX1OE1ACimk6XE4vnMxYmvXoSkacTfbyxAAYo6NRY
EBmhBUBJfgHxZRevwdzy2XmafJVcozeUMEfiHSYtLwA4MztsSUxAu9dqIs+e
X5ekC8lN+GHRyNEG86qkbOIxAvavRWLahRmX1DA36HVTdE0pLW4kiO62YEa7
9FyP6bEC+PazCUReNtDHxMEuFKUOiYJ3pOjzQla0rdXl5VjyUTbOqXh8Tb/y
7N+q1cvajOqeK3oSS9vTaJUCCN9IwKXvHkBtoyjB+WG6O0ZZBdQRC9Lr98+5
O1gSmCDooKp3RyWwGgwYu7t5YkT1nZDiSQffILGKSrZ+XytAHbBJ4YpoiR9g
MfAyERbjVhU5juZn578b6xX4KXsn29BHdO1vWVY9ymrYiQHE7hW/AqJYQGG9
rNy6gAjNHEjh6WyoVjQzhMd2NJYB6xa/lRcRQuXm+/hjZKhIqiU1HD6bG6Gl
dQ9NBFuWXpVAfyr0zky0NAEyg9Ll1NcTsxcTlP1SmllnVUCmKBNA0Y2+IOJo
S/XDgIFQ+i4VO9Bh/QS26YkSqFY07U/o4+JIqqE4TBykm9l6mwVVXCtUO0jM
KyatvQOWXx/ms3XGkXXRmGlVQ77Vh73jEKRXPrg4LPuq+oYNhmicfwNbLsIq
0WbQn+q1PCc7OArbw3Jv8A/KbWZN0J52nu06I9V8kfx83bJmgBXzzKsSN0Br
APddI/CbmcWPFPS8F9qop1DPsmXVSd7qkRb5tlCf6OZatjotZf7s5UyjtE23
XVTFdCMuDoOWWCFRLP1CwfGAvdihLIhECBNBjsFOT+HD2wkwnW+eCfxNnV94
khuLm39NoXS7w+epPZ6ZltJHY82EkXbscpTNuURcx8BBg6/vg4LKs5aM2MoQ
B1AxyzroZmr9FzKIe6rthQDdieoOTs+PCweJio8QwkxFTFZ3cgEcFdKd66od
ZwhZiT6mRC5nEbLvYl98Jql+cjn43ZCI3UDO9k/jaoJI/FHVM+GX05uXzv4I
gnUNw0Xsp2tywT//ct6fJ7JxUgtyhIyxo4Kbed65wPYbHVn8ARXH8l9QixX6
MAsu4EwdvKyBgebyD7yZf//+2A5M9V0Ib7FTM+ppJ7HzdwFFd/sHx5cExZlw
zZV1+A+xPHV9LiX+B/ll5l4V1teLFulYuMjMh3N6d1Mftzu8AzAZAn7z4RYh
ZmzbU3PEcelWZFIDqJCeqCcHR26icUZ0xVyDVA/TAmy8WCnv4e1Pi4vCpSxR
Ll5/rV5lbkcE+18bYTovrpiaVLV8tOePi3iVYQwfYYEnX5l5VFfCxm9HuoVf
BzO0G8Hfu9RDwfavP7y3OZdrWAjBtMZCYzxs5cFy+V1ZLrKXGuP9rodtVYCH
1ER+SDxnnoeDgJshmI/1qV9nlJMoXyGviVsQR7EWpLXw6uUNW7YZdzmmeFWR
8toOmhVyMDFw19Xgu25H4U2cI3KXGChxBEHqWEw0PipYQmtC2RwyZ2pczs2m
MJh51briHiVbHZhXZAsJX7iaO5CeqkSzXuaKOyDRd6DntGjj6e+gr/hLvhRz
eVDdW7XLEGBOBBtn2d7tuOC9mCn+jQNIS97/bt5lQjhP698613tgh+EbjCD0
dem7wVpYVBx/Jv+TtMSi2WbYG4iFDefp2ZTgFwuA61aWblhuXiYVpwQUoUBA
cSsI2fGeQXEY9ci/Z84cj5xarUV7JFmTwzLQheSMf20QBbUrLS1+KRKyD7zw
k7s7ww6pq3O4WBD564iMlx1jmoD5VULIBCtkAKmx26eZkY+JW+ngy641sq0h
J1obHpd6Yl12FvyqzQ4boOUHKAlN6lB0jAbM9eRd3dX2O0tktpuPSmDobneH
1kneqmFKZk+6qBR9oXUsm/YBg2gc2gS9COW5pMvQxniDeuK9KdNcHmw8AbWU
6Ytuq2Kkl+py1N37+bChU9pri7IM2UP7MN5PGLU/gAKaGWUFTYnvVE8vwdjc
FedWUASPnu9bjdhna5yPUke3Y0v21PUg2bYWvzS6l61UMb3eHH7DTTpAxZfd
ERA0T8NVIQmfNkrtutqArusjzRiSNrk/9EnmJqsnI1taA95vgXM7u8lsv+dV
9K14gHt5DGZYdrx9BxUZ0KnJpmljG9rkBIPqyCfX+f+UaQAlMf0FrCZMgjtv
S1xoi2L/o3ChUkDNfniXU9fcBG6UAqwU9jflhqxVHNpFlVO2RAURX1iKrWLx
AalgIkbbn4XMR/vV5LmDEtU+O+KWkYVL8wmPgDpRMOpJEeFFdPXRcsvIdAWT
7j4y2eyJge8bX3rlj3dP3g6kF5rrs1/uWbJxEVU2S4hWT/yRX4jUQrCyA1Jz
Anqep2cdP43FqhUALwz6qp1EPDt3NV3gzFgxAE9vcF2qJkjXg7tsr8GI9alH
Uq8/eTFR50GsMMCLjb4sLcAlqOaZWG6+PvMfZc5lby+QD33dH43w76thGMEB
T7MAwYFe5YsfV30NJGobWqt0Je+u8OKqTqikyZeX3L8NdrxymKHvFwD29/uE
zpdVA9jzg0hjb34TlCXpUE70h7OvdlRkKX5hUO0Qreli8kbdZAnTg+BY8Vt1
T61AMUuWFiDadGYmMMxi8CBwBgK/vPLbrbxs5TVDZQQpijFwR839phQfz7KO
3mNtMaEhuC91Ppljw8qSIZlc9WLchtHCLtYAiH67V/mFTI/v+Qn5e8brH3ms
x6hT7Uc1AwVxaBRmk78PxuYssktOgJegR39XhlKa3difkiZhXjFtIMgOlTYS
jSdjMk5ENHzFUQb1wY2COdgnWPvMLqjWz2/+MBbCW9Z56C7cO3mUEZaMSqW6
D13mQxoc6e3sThZej6c/Acgt9ehrgIRGeUwmRVD2q8AsRf6XhWdlQ8fENbAm
5G8TGrCD50MCHLNGpo0mky5PxUVLaQhfza0bX2z40y+jK/RFC+Cel0OnXebg
OebM8PQUFfUD5jfqfS8eh229rXXNoQtYlfH2Gb1OCHZSwx8j0GpM5C+tsQBd
yN8Q0e77A4JMw+IlJpzw0JRXREXbpnzf/Yd6QD3+pgvnm9vHZNTUvqiExa7X
WSrLGN5VKaDi3RSu9O1wf7iyImpKVj7XJx3466ftKbKLihhZyTfM+qVy5DnJ
mcdhjDriytEKYT1cwidUDIi2BQq1je2yf8p2Ezue/tPJreSlpdyH3AkUUyAx
N912I84kFkRJ+kVf1KhmkINtWQGxzYEyxMTEiMYAAVbCMrvCh8fluBarXsW4
/qrArr1jNBnBtq9ihgLhz+wRG9lcyFjGcSm8KqdOZ8j+4BL30DYSi6seDokL
rzkcEXxKGBes+jjEMCxFa3NRtAeuKEGTq8ZHN4V69NwEBpjOvjyW07B7Vx7H
uSGgsMIPwH6Qi7fMrxchDW3eaAlmndip1F67C9FpnL2HjLq8fKGWmfU230Sn
ziTm7wQb7o2O2yROKNzi/ojrfNCy50n2uNq8eM4ES2oZUsT5yFvaJiCsltNA
7lrzfeLc7348kFp0fcBQ9riZ5yJVMQTcFrETSSXleaDh9ZNrw6Wt64LKeH/W
19kFGKOYprvPG96kcy2/yt140HKbKZ7MFTdR4eqc3YM1EMNmMlg7LAxxwtcx
b/pgBmTNyrscqF7QbrHGskxkcU6psEHAH1PSucG+I06gzgprWLA1SlZzGwnF
1OF3J8aKiBVrNcaIvFST3G+KvWTlE0Bb9NrHGE6SdNeDv/LvEqTr2TWr7up6
/+KfHKHIWOdaIJwlwijbaC/rSFIF1IwSyg4/NBAQeyBKM4kgc+/hQWcGJg+I
e7cxKHBuKoSCzEY2QHJ0aBYkbMZIXxvbJyN5wb5FOdemBTLCMgjNDwZhGIiT
9VFZsisthqEFz0zSWeHDGadXgX/i85l9I6UIel4Zl6566hphezZWEEgznMRv
kjwjlHFG/CTZaq1/P1/tx2j1mGN5dM7ANA9kQbyVef0uHoiKrVfyMJG366XM
wsbrhIW93quRgegTOlSKYr7jpvZXE9+mTzGeogL70oa8J8Jx3Wzgy17may2t
G+OpJOJudPXMUCj/R6QBFelVL2ond+qpTnV7JZSzOAwyfZpJXTv/FvScXji2
rA5d/61S0h/LYNLqC9qg0w6CWj4XcVaqrOccoD4eNP49CmtRR0WKCbICQP+t
4o25yjlW3fJHTePgtek9gBRDNm5e8/4i3GBW0n45eidIZ1GsKllzZp0ZzaU5
Gdxmrni3c+C3NwuQ1leFXeB9uT8CY6yILlD8rzU56Oe7/iNhhNLdMJIHmU19
0AnX6aHXKNEnQqP41kzKL7C6fGGbQkPYzmyqLCdBISiYXMfA+CAUsF5hx6cv
h4A02SFRuupYRpuUQna51O2qyhCFAtCUWAX3bHh6HYu+0QJHDUbqqKlBi+ez
86lTrn4WcAfCucmcsBZQKdj2AEbzIdOcZBbrlrx/XmPplxmtTx6fKi7bCsY3
N5d8F/YOZe8lV35ib8fcKwmBTpngtZ6hMXr1JUnKCKqmh+KqxSyMt+7GW6iY
6APAVO5pJz3uSwy8qQJTTwMmuuObdDANYQ0NTQeMv3LImglJ8lSF9gIsYrRt
wVd4Lpinp2ke6aGvFbL5P+hdPndIGXnezVqbm2HknziN2kS8ms+8UyCTyYTr
sYHdWC3L3D2++J0lA6BY1BOfrPzRCumTCLgX2xLBTozf3jNirWGkr3AS5qmb
85TKp5rJS598wp1fA/PsqwfB1AnWplEvac2s4MgIx92c0QSDIGZbjYkLVWA1
Ef3UhLlkCaIk6LJEAz6Lo4iFBXduClxghLGFsOmTgMJgts742FH5HcK16J8V
UXHINS0olcwbwzVp9DJFY1B1CHhsUxvrErBVYE6x5iLe8O0MUR9rWRcxCPQu
m+HNpwBWMUM7unX5JD6YYpsAwJgpQ1PkgVwAkRvZPJqEaU0kBFzoNskU+FE4
Qon22IiS0KE94dNo0KZgUPT9RHa+rfmYBv9W4BK29BjVH7dOhlg6gWx18KsD
tMChebzq+bIOC1dA9YcfZhHgj4hBniqvyKM/AoeCyP9P2Qv8uX7XRbia1AVu
T2L27p3rXclYHdMd/8bCFrD4aOGUkBRompIqU6cJdpY2AQK5hH1K99iFx6fd
00ZUy+UemJlwGrXDc3z/DzuPLsY84HVHDDxtbO1Vq8r0TG91QWq+etWEzW/6
Noy3mNPPYN7sAzgewtHLxBcgd59R79qS+BDKwDJcws8SPQuvjTlPZV+u+AgI
ajdIJVkuAhWFv1ue3iqeUxHVbCrhDrSEtRh5brPx9wB7yY3hT5b6iFE4X7EH
uI+1bgrqhxfNSzLkUEDFprCs90b5UnBTaxDprgzYCLQQP7lEGPpQluzE+VDO
9DSRgTRQuFs0G8QaJGoZGqEiZnUSpQs6On+ASmju9u5SKbwQFEY27Y0tSrMR
V8VUZIzEpPSoQmbPd2vgODZUpmB2LAq5mD5fDFIWEMNPxd2Ijq1YXJ6lbpvR
bS0ZhvVy65oVA/tIxzqqgzXYHd3Q/z77gbsR/2V01SZ5z6X1kUX1n4htLsL4
I6Vg+I4RAWuNSC+NNRhja8NuDAG+ayF10yo8fY0jls6IBxv6RCYD+gjiRIrp
HZC8IFE+L0vdZyNXe8oaxwDHrY3QrX9XBYBBaMWbuNPPozXLxdb1qDqYtHA5
YmQIzPud1r8eX1iM65efv47+FQCH8MG6jkmQ1SpUvHKKYXLL7GjcuoBVqcXS
v2akwYTGqK+SSisQW3lc553uoGBLYc/5pNWXwZTDLtL29/A7qM5wAz9nqvoD
zYqxVOxvYJGou62ADm8JvJ/jNzDO4/aNoGD7pWjN7eqSu0nSsIQUwusgsyWR
WIumbyHcdrLWpyOgfCPOjQhBXpScgzWyCIZyAguh4caiK28WQvKvAsg7tQp7
zH3+TRUjywB4AV3X1OyWCW32SVao7qsSG8uCzLhKIVRQ5N4b/ufncgykYWe7
PiICj9Ca56aLSKUCW1CuxSagJ7eqIqflmEamwe8VqQ292JcnTp44SWtSLRI0
I7u7o1cYUSYJLmCbmlDy35PeHdTe96ZsVh+acL58ck7ZRnqDE9zXhUi7xs07
lqhBCFyJ9jp5zFqzWioQ0K4ZMfIA5In595iKzLPbwEQqVe8fgIzMMGVQwesc
jJJ4eAp59o0NVTiTDRNY6t6mPJ3dVUG8dtLmqSx6wzgHJemD+0p+Sj+NMugZ
Ew9qLLh+9h1IDHVa+/c/JvMmlEuR/iRbImoz+ht7NraQH/Hydrux1kjNkmoT
pBK6YwuqL+FTKOy7UgcZ61K2AsTycDiDQG+GLFE2r02DK/rwKP2vaVPBAFVl
m1zfLB1E7cw+MK774WXS+olL1GMIApCwngMhsnXTYOw/rFLUVlkK2KkzJK/y
y+OKUdx7LRRvXAdNT1umLOprHe8Uy8ZhmKKjfixY2/q0HC1yLUX4IiKm3ujL
Fgmrdk+kz+06qebW13hgCPmW453g3DE9oeE2Jas5x9tr6qXqW0OCJW1jydos
QeTS6xspPMMxxC54KpzAyRc53bEY7IlIgJSRu/aZKS7WSDTUERu+f/qLSQGa
J34TlJE3TKZhNScVcq/gRN0bt18llk5bnw6EaKcYPncAXvtRoXTFdyx9TZmq
VuFjaoKuDQOxNYjBSpx+xfpICV6VgpwfnFn79Xl9p20vEMxYuanBHOn0afcq
aIFo0I9y/J4CnGTMGN1Mmu3fECXvkICI4QebUw7VzQfSaLSZACqBmweCkrXG
jlNxu6oc/GhpGN+KhskMvWtUcCPznIRF1RWjpJRgf09EYuARVu8ZqOPm+3cY
BuQ7MBYYsW632hLRZSTEf8RfHyCftHE2ITaJWniFnZM7aVbnHiNiD6sC+a4u
do0x+vEOCDHVkdIztaH+O+tYKDY5621lwEqoJW5gvomw3tzAacvTC7PxpDYh
cENmgXsZe6vpOSL2k8YvEt1WULqFDqIXnbZ6xPZHolJ8dIJFABb8nq4lvzE2
ouuf8kEtAItNN/CszUhuqtytkFE4N3OEqfdAqktMnwGS1sR93XzQ4uO78eWR
60FRlZL+vjIV3cAp4+uRn2pBgVMqOr/KzRpX19UqoEo6XVaoiftEuNSoIr7y
rg0PzxBT6RulqU1Nl+TUy1ETo1t1ELpMJ4dBKMykBQwaTpfEEwrO0GWQnICz
XxfeThPOVPWueb7PW5lAZ7HmN3YFZLI0gxJZEWAsRx8y6AB9CXUw2B0DdGGD
/mwAjT5GPt5svGeBWVYjgFdQToI3PvBLg+S1HOEyv1e19L0nAz8AnKRtFOFK
nVrjuQYdxCvCZ6yas4yklzssIOfEk5hFOiuk6mdmHOl2hYFfsUFC6ctYWwi7
3oQSoH6cVRXQ8pT5cCTx4A4rLxVTDR3BtyE1t78otRHAbafRmeY5GvVKro1d
1kC2U1xkvjuGIlsIaRA0eWqTQgCNxMLFMU8lV6devBfHDCFxd81u1O4eClD6
3c0VTRq3QLkMurDArKMI2Ag0yDx3lbMBROUkJiNi1/J4Tu8HDbAIblEjPp3d
KONITW9wEM8Py4i0DOQZy8iTa2gUpbGFXqc2n9XE3KK5z3jSGUz3DD0ZJefx
/T7EfPX8uwgEbsdH0VVnDidbg3DlfhQsRuBpAMqGEs3pjRssKX1gYkMbTJlr
sXQb6am3AJ9X7p5a12ivZDiqmRlJTffM8Fqn2mAv9+9vgysyIC/PDpD+HKEv
CVHzVOVKWpFVUgZ/4iQnOEX0PY4QbE/DjjiFx/aDecmbRRbcvVov7FR0icvK
pGG8VsXyrfANizgpcvBnU5A6Yc0K4EzAoN3ZZuUa3EuGIp0akYLKbPHgbF8j
+XIogypMwQ7+JveVPxs6UCyVYwhEu0PySx+zVCRE9PI22dLnq2C/DrLg2V6d
0KhXX6KG/Z2cv5fkDENJNQR78PsxL2rHBGCU7w+fG1cGZqof9LqhLXaOfkqR
DMdeL/qDkZvn1uDP3rECuJErojjAAYQEcgkUWvzjGB7VrK/eZM1a5kfiKfE+
ock20D+CFHlXIVQ+Sg3s1Ex2uqsyQVu5nb7oYXesEUgwStuAFJfHS8rPPXpH
cRgY91GEbdMzOOmk7jrvBXNHCImR9u5B/jFh0hgrM7tSoMlb1pvaKnYKABW3
qI7Cn+Lk121LmvjfwFycCyTw5o8WPjZbctnrPvVnQAWOPqS03MWNJcTlO67e
4gXgqvWOKgbrNPjc+/8W5/EjUgOZU2TVbgLrzcFGORR3qsuupzMpLCHdySJi
nTMq7wKm+mSWJbdaW1HY4MIeWGP6gEMTsOV/kIJyVtcO3JiH1U8g5QtyXQ8h
k+smfUeqY98GMXLJvn1gvHhButduvEnQkIXQd/aSdYq8PEoTEkiZ6wS5kJ/K
ZhnTNZYhQL90i+gdF0NJ1gao3k4H+fIzzzQWzwkQbRaw/uuoCAq+eyuRSGR6
0udz2aQ25vtfd/KNwG/dJ7Zsj1wxXWMbf2dqYtE8zQ6jvl5QK/ZTfeSU8qsf
Xkhmx3JI2KA71Y7fzdamBROEit6i83AeOkJEma5EwjGsIx7PsQCWPkB5Q4Oq
7EorB5/rzjxCtZZ2Inl8w85WgIhoiZ+tvEVhUN+T+DowW/VMBTp/gtCo0/y9
ZosP0Vs+LyNefMegH/dowr9fBkgzUqjlOhkqYrPav4ticVcb7Nm0aNnjYOtQ
KWvjo71oMxyRk8d/v6gehuyyoa0p8IrmaapWKvTd9i4fWUouXg/i9fk9uq4/
QwVfSqXFX1xNcb9wm2MhRTUMCew1hUPhJmZPfR3QHa8UYbmKxUmyvtnAUaam
oapMofbZZjHqPW5R/Rnqkm0HPPbpTgp7aM3Hjnf8hRolf/LfvWoFpFtdT3wn
Jc1hFJgOY2yCSjPdvUx61MyuNnIa0qqkLZQVokWXlt+LbF8S4JZEoONSqAQD
LRzAfHkeRbJ0tI2TqoxCI69EYMHKRF1Oc9y1Mt/RQnVwpMS+5kUy+j3OY4A8
d03Pbfa0XF+RFwxfH5CSdyIcQotauw1ueF6Z9EYrZ1nqClS+eE0pI8Jv0ERc
jgPxiz8cL6sywI9yLT8JiG3No+1zOhbL7FxVY5vT/qv/GObAcr6hhlctLXnz
4tmSloHVvHSekKr76FvxOE6g/MN2ksqQt7nWvzWLFn2LvN4cg7xy2fx98FnV
2B+kXU4dOWNrPlyQzU3+6x98DBVCjkpzwxZgYEAXiwgBbiCm947jJml+jqm2
RGG+ezyCBSqDJS5JceYVNaBbswK0GQkweO6ekpSAHOQyQY0/wbHDCpfKxeUR
XSz4bzlJie8KsHkUahpOOfSHEeK5klxBoYmjhfaOb508sPcDCqSfnJrL+Idm
z0nAzPBHuBlJaM8JHi4IlgvOnt2pHDtBDKfUO+v/E7qsD/FYixM5uOUuDET+
a16W/G1qEB+XyjCdE0WBwW11nhyKRaRJ2+BT7dJy9/2TyBQSIghs++mJRsvd
KaVsNfSBYJuD+QVmzATRrLHOijbuSFy1shrYO/W6Q5d0EeDaOK3WSwai4trf
+TZ2N8rEW4KVR4m+GN6e8hE+YiMRAJNFttd51Vvjsj9BqQuXgjcdjlp4yux5
NAMPbyz56ln0HlkLZL7Iw20RyvaHJFUKTMSE+MSomxy1bsAeVeBn2tMmcdgW
6BoA3COmiHkTvOaC/aIuvTf+JqvFyByuSfYnR2p/NuyMklvAWHXcmGEKxxTw
H6I4+4odaq7RRZPlGJ+mpXzuXifrYKYGLI9gjXpvGoA0KIAZhTlMIao457Ab
UFxe0SUawF14QPjynaApBLTROqq4k38fIB3q8dbMJc8c0Zu8N+YCs2PGJhzc
knYUAzE8HUoxhncWAZk0fnF8g7n2tLLzKLs/ToSaCyvTNJxIyGOMUP38roTh
b6UnaSuDcakN5KQCvFhXqkcbtQoNczSkdizNB+cVqbts9JnqLwW3GbLeNV8O
1s9k4wh80txsuJBbSfOQUSdKmJFnq1i/ssZDsbuJgkNBI5L5TfObhRahwlPm
6bcuiBHYNW7IdD2tnM9PhT+Rr4gUGkVaVJdMdtz87waZr6v71j9nJ6QczSqe
ZQQxlFO2kc7TC4FOdd5gTgbMJICW/U2cmZuF2hNDUy6vUBybgFiC2uSQHu4f
L0KLM/PJpHqgIug4EhbrqRRJpecXtFVG8xPQKWLkhibb2T2EC2NTT5dNs5Uv
rxIAEKLndGJ9K7KL5KJ+nw3iPlD42wmmIwy2BAFgaBR3oqdzirHiV9tk0/Jh
D+PsxaH58q18m2/hBMu7RkoCjWSKgnlMHcPiYlv8wTo2E/fVheHJea+LwepS
Gof5lwQm2klRRsDn8Hh8Jsi78yALj1GzCFK0Ms5HXOtjyfEiA9iza3+jwWE9
26JEAMKdiOT5NJQuKaxbQTdHd5Hv+5U5KiJpEbWcniM8hfW92hYtAUWqJ6cj
SK2DyE2PD9qEevcl5ECP53uBUMXxxsXijnwcpKIxK36ZgE5i04dfkT/580LF
d8DMH6QKbd7zIOM54aW+/nxacGeng/FYNo1X06T+VwLUp3lstVXmsksCvcQo
n2XdELej3nWOaYjUWy7eNehQ3Zayz4BmV/KDdKGQg45K3rxT35YN3duhwdjG
Mjl/NpVva0Os5F9dZlwNdhbbL7Av2Qf/C8uHsvAb0VUlnSDiqRoTfhNUuHgX
x/l0LYUD6AVIwQbJ2grwoy9RsgxSieKgrJSt0lhDUlzram21IDICI5PoYTHm
OL+ztRbaS1e1PCcn37uzGjCkKb6NTa7g/V46A91Wa45Jca4b7RGjB5MFxjxw
tRxbYPrI0GHmdIK5Jrg22cSr2k6X/7ShR7ayh9/TUyGZP6ePa263tjZLzl7L
N5Ii0HWfQV63xcDu9b12bOG6izKxT2Ntq8CCZOLXSeU5uBvbNsYjz9VsJm45
1de0SYClqaD5o+W5HHsUsCzjcAVgn8MS98BVkBYB7H8EaTRfjMim2hWnd79L
S8NhDeG6qQkpFV0GQ1kHcJMD7kWx3x7nhcHyo0k5W8anJksfZTEXz2gitGyH
jYExvjmh0C9TwPiXAJx3dfOWueFC0Hre4AcBip63NKRTyhX+o0PfwRTUR7+Y
ae++riPxgWNgD83ndl1XgIx3+aE0VW0EXuYlAVEPRkv2mMgEV45X/fgPRj9B
b1uZKlK+m8uhLip5t+qqLuXNYhNuhQAwlSeKIKSpphdXFUGCbatg6zo5Oazu
RmxJnTQVlmUddwnR2ohCRc8rlYlaal990VXQ05ByhGD1lpOujZrt3UsRFxGg
/2hYKmL9gYhHTrXZ+M6rcxe4av+OqDqJJebNx3jBjG+ntRTM1IQob+pBeX08
5YUH4sZzBgnG2i+g/+kM6/ZmDZc7yoTfrW0++8hyn7it3u8FHVSKxWxhFDwP
Mh8JsEIUWheN0iHLK7UShAoRa9YAqp6n/ddaReJPiRhfp+KkQWARy9r7F+CW
DwQ3q08Th8swCT3skHIx9kLIOsNJIut7PtpoytA84uQdoEAbyzPlhKem+And
4H2ryPrbdQaeIiMH/LeErlL+y7LKQOyk6uwwD9LhdlR2NRV5QZTPpI3xuzw8
0V8tUAGn14qUNJJojYXCCYS6FsxcLLWsrgr+0IBiVWyY2yTD8UuhpVDnoO4P
erRLu9WEyofgM8ElX9RKy58U1qX1JeJF8gA3rCZ03AOQ+CPROxS53ku+T38M
NAjz34EPFxxJwdRUtk2QZMM9RlMC9XIHsRuTgcANxbukOinfZgPffFQRPBgl
jI5tTjVcWG7KDJWZOf9iixk8OAYM6qhtZlvePdktV9TYv7jgFSqnqXYVty66
jHSIUoUSxmjRmXXxBZKKo1rzE4ugB36oCyQPawxY3ltIoAul0VjtDqrBznnx
xfkr30k1b7xuUk/I6U42d+ZkDcJQivpsDLFuP7i5YkecIH0baQ21PymvoO3k
gEdTRBmhOgxyzClkjvIwPY9asLb7jm7Qglv1LVtHkNgC0ECfl62uoDCGD1S5
LCrXQMt3USNiJW4kU0T+thKAqqB+v497bmyhfJe8OzP00XlOewIZWcZDzBBh
U2qwuKz/r09RPtHzvTa9DSZVL1i/FNkHcJ6C3CTvtDLzLPXviMrut723yJOX
/0CyW0rWdI6hKJRR/c6E4Rw5wLRDBlSF1OUhNBnjdrCcSb/CpvO4iSm+XFLv
cRnUNUCdIiQqdzf2V/Fus1v6CleeqE7IQmZ9/lvq5jccYBA88qY66AmFhxDY
fAr/UVKjc0IQH6ZlI/yL2OOOBzp5U6ttsozs8lBhcKsaf+0jEYQ4MF8hlihu
BzuHPolQs9IeN9W6yCTygOpFrtfGhf0VWM55bzh3uSye6Hzge6lckr+35dPc
0eDgIP8wgdZ1Sky/l7hZeiUcQju/+NEZ7S16t8chGO4y9YKuu+VpUQLeaZQS
nyKg87PcO/N5HM1tKLkcgQMtfqCo6tY1yYA8EqfxXY97N3rQlfkwoenIvSO7
mSpAwpFkJDAJ/trPYMht0O6+G8psALzCkrVVeLlcj3F0q5j0PAojbw41ICvi
EPwdvWzUH1Gq4XDB8LTWb0/vJxcxEj93NX6IXou9ulMZ/NJEo1r9hsyLSZwK
+4Bzcct81rob8G2y5IhB+mM5m0XkW0T5tCX9mR3JNgvcbG9zrsxZAMpfDLd1
RSVyO6upOMGpA+aBZinMu6y6r7uTewKIq3lkl0HuaBbk8w2cijS+HRIFLcJE
k0hubvE3v0e0erIj7CjKbJLtIpwHLbBBE/E25riKYGbdpA4/9WMg37Ks2lZV
WarTglIj9JX71QOOr4IbYB48Zu7xv+719CJZBxrAM4QORlkWc17tGnGoVAzx
jZAQXHzywdJ8RdOsxMn3EpbBTnD7kBgFxwbfDC0prYEFCnsAGr3Gu2VI8JMV
uiI5pGMmy3OrMlMIBKA6XRhHnQlfUOfb7mj0DKSG5BLsepzTKFsWXCxfpdjk
q4TXwWarCjJa5Tx8PRTohdUF32Q5ckO8C1CXFS8KyMo+Cr/btoyFGYHGWAf/
vmnU9+1E3Z5RdZDIVgJBbxbi/OsI/EndfCpj+73KCrLcRaK7teMu3HL+RLlL
lT9Q2T+Cy78rspZaLiRzorik/k/yP6pmXmgCQ18kxzglroGRhNhe7E6ch7qu
OEiZdEzIhsVhY8X4TyutaelSiN/kS+QqJDRRVM+jtfOfxveOXi+mC+3IWrPe
npom9bQy6sy+ZHVnvkDVLTCHWcwkQN3Hl7Zn/vsUlNY+tgikBLu3ubbuy//Y
dL9MqlQjdSH4dsY9ITzB721f9FW8QlLUgygLd0TwfB44TzH/5AQhOkR88dWw
7sSzbicQQnAlZQJxf8UUTU325SIgz/2Yqo7/d7cAbrG/kj4Vjx9p8eeZg4Cm
O+7kJY6ILD6zFCQfzlP23sLlO7FqQQ==

`pragma protect end_protected
