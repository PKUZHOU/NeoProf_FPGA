// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
a918YayEnTjNUj1SDAJySHumwjaK7zZ6xPm8eVjkO5dXlobeZgesi1Y/7pQGFUzkd2hPO0tnbIBo
QG3koc1rl8Z+xlEvCW40L95YWuJznk0SUJWSA3+qYaBDXzbWJW1nSMftTYeKNSYheW/UnpcxMLag
5DWMUHe0kxxbi4vVhmReXb0DdswvI5wTJmqj1+6aXEvm+KJUindtR4AVyrsj2xrB9ptRZyW9o83L
TM87WG3VYB0BFtyNNiLW9GmxH6sj8dOxQPerv1BNYO83/asOqANVQ998k1t9N66aonFaoCy/Ku9h
yIlsHqrIWkQUnU3lpPFmH6IpEqV9w+FiDbXK7g==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 59792)
lGxWP0DYKpvGUWBcxZDps0dTUxrFEYHQx5cZD2PAEpyqibemyRNqeoJ8TBV+NMs03yKaQQePfWbz
2MRYj7hbKEiaxbvI+34ixJQqFrNN5Ct33R0pn38rxwbObbAK4yKXfoLhckLt7ds/p88XIc9FSUzh
PfChFk/FxUDZTOnBaxWTuRMfVRu5/WLWTwIXr8R7Hf0o114p732XKe5WRc2lRqS+bQk8IKqbgdmK
lKOj5/2sno+1Pezx31Gj1fimtCTIVpEy7FnEWEiRd+5vKJV59DdGAvBD9mILpiJmOS3PTwf2DQ6R
Hyz3R9/y+27Qznzk5i7JgAlUFR1PUzyFU4WC0gfhpjOGjD4lYHIzT8nFEozLiwvNwhfcdaseTtYU
jWAn5RDqh0HZ9M+lESs+rkpZ09/nNW9lR5s/UIirrU2NwNpsQ1yOAUYMuJPZQN2fiq8eDXM/Se/V
FYoer/Zw5jh0tCgFYPiUEcsV9aoOxXEu6wt2xBoMNcYvu1867yqiFmLXmSHavROMR/j2s/PvTK4x
6TvFgBNGaL7zrFoloS2PuTl0xo2x56wyD3qrtjJamm+jwC8zRSV8vwc4ssk1wjsP+zdrXkW171V0
1ODKr5AMeSYrOC88un4pa5GgH0izMTSSMciQucDjPsCCc4HfCF25ozzK21pa/UeT6vMqZtoaIA4b
zcr2eCcALzU8hx7VFAZqyp87HZ79hpDVopUorK8BZcZ993+f0g9FCGYal/O/B1UISVK0TOjDGWkZ
LYohDxSodDyjmQgQOe18TUOVSbogboJrSlft8W/uoWGGkqccMA+vVbJducLxW0k2BIpU/zQNAqHN
pFmRiZlgomU/23PlMZ59E+GJ3Agl+BuNYjHqxECvXOay81LQhaKBafU4+BJsJE84AsgEcE/NP/fM
x7WqufISnvytfVN7LpM7I1prChmV0MBB1G40M06gaQtBd+jC/Bf+msE0wWymvif5Apd0alj2msv/
0tuHa7W2/oF95vp705F6yEkq2j1CBk8U23S3/xIW8SQvV1qnQYqwp3IdgViv0dGaV2qkSTRNceuM
+wbSB+R0F5I7HzeEYLJp4IhTJ8vjUza/mwmUGdU+p3L/DjEYIYmcSa8PH60FQT4mmq0ghF1IWKqc
ujn4aJb0+Hu0yj/MhtD0cA1/kZ52FxSXibkk4CHTZE6Cv9ZaUZ89Fy6CzTXJ/ZM9o9jAK4rgnXZN
HXc0qL43t4JYx28vr/IpjFVznL6ISRqCXBv9MVI+BibqMlS+OQZf4GVVflmPd04Vs7zuisnFkuGF
niVHMUGPswT6uzrzbJLF12UmN2fV7HZEZ4cTFsWxJJP7X2GAHBYLlFB7x3bnbaIDwy2tnfvdYgPm
Fu8DJjrBpALKVbOFLWYh6CMLvIRCe6Cn13euSyCw1VTCpNtkphexPV1m6yb2THjUuwIYnRNCpMKU
KvnSYGbtHeLWIitBRn26EfwRG83iioWP/5JGTaWS/VTsWzjN3ajA3vn8vlaE8fSi8prV8ubMgpEx
fo1JBvoHEJUxnh2S9+0QBUr2IgObUyqXVhPawc3zkvEnnQsHwsbm2GLO2Fet9vXRJneOIx/35FoM
MJPy6A6Ac8BuUbqXrwKFEIrePoLki1JzG+drD8HuS5rcMz6walQWv4O/mKLfahPDTdqyzQK/BQ0R
6DEOLuuv7tN8S5IZ5IGHMH9ht8OBMxzGyFAjkDb1q8Ecd0vd5KeOW4R9EnRYxsH5WtME+A/zEI+9
bXnrqvANlHhU/ZsTm3WzW0QG0KCf1rKmjqZ4w67zbwP+Wc2YT0tmT9hXiqMWqEpX/kRLLNh68O3I
SUu2tZDBLAD3kXe0veJLW4CVF3JP94u6mDXM468SscnJCS9w+eTKZTppzi1YTu4GPWn9kGXh1Mzw
s3UWW0D5eGftvFkCnlYVq4pIYHFs3+tE1+CQr80Jg1ePrqjAF9+A7jtkg08O1l87GX76M6oXQA3M
As3sIwQhYWGFkcctFUxN49vXxiND8BaZ40NDexTWp/gAeMv5uv/syUBgvoET+lx1jpvnDBE08LcU
f7k/iByo94B+iu3R5H7YAzK4y54Mwu/3T7zb06keK/i37P9kvWW4th36tHsDKmlmrVSxoeAEP7o1
Z5xOdmh3y6WpvW9hAEYa6gxA7Rr2TOcNP2FwH1gTpZm7F1JV1K0C9jJ5Fcf6w5F0pQiiZrcEMUz1
fCCgUxF3Ipr4ov+cshM+w7YgwjsX5mP1I2g2fQaXwr5mWFLHLQ4zqqiz7uZLmWAQcD1WLtZdODyc
AM935Ef6st15DDdHbenJ1ASfRBYU7OsYMqTOPA9H+K0TEuEItmGofGCDzo8q3PBq26wJaxDvnru8
VpsEIa1nvUF6UMHfhiIClh1FHZcMRGx4XDqoazYA1cBi4xAdkvS2ZwMBWlbprJG1P/dDxTRPKUU+
zRSnMgpo49RTQAxhIxvl9FBGVe8SQ8MVh0VMpxS6jw9d5sG7tWhZnKyo8Pp0xpy2c1Ser1oxn3eu
MBJ88nuSMD2NII6947BKuYwAyamCD+tmH+SaKeZ0np4yrQhJgzeHEpLLIhurCT13R7PVKsoikVTD
BoimfixgcInGunrzXCMiPZ2Whuc2XkDin0WvtPwDvcO9z9Usv8oxnWLjfaZp/J+930hq66TB+Qs7
tQOj+818yyrHgpO8kLgQJ70Cv6wkIMbSS9bPT5mNcuniCugWpGUn7zqoqrRZh3qx1ejRj1XbQnIj
MT3ReRbX8yigVvdw347zeLITELyXiN+J1BtjbT8/SfEMTYu622c/3Hs4XQ7x/cHcGb1vjOGdR1t7
DNG2TlusDUh0J0WItuSAk1nUr9GNxymMG9pdKk2HwIEOUzP+k9RKefxYYwl8y5FetRAWuvFb34jc
rTbR52LWSJqpH+esm6CtDE9tczEOpvEn3ueO8OHoEMScBMyJb8fuC2P1XVDlOhnZGz7MGJ58x2dK
tGtLgwwgE14/ejCjGOMkJm/2XiEe3qnKCCb0azvTyiZZcZGuLppYA9jRhVwyhjHp+CvAci4V6I+C
a9/SPDEnaRuMgyFeSqZsG0ab5hSn9NOj30WI2AHyqliDQAUTYwXBd3Oe4IB5eBvmAihsxlBioxIx
wgUarIMIR5YVkYYfxzLoXajSjkGPfu50f64jPeFDwLvqZ5yOgUp6I+j22o/zpBUIjjokKjjeeiGI
JMqABq+XslKFi2rZInnLmcGzfpbvdYy12ozm57daIzGyT7I3ESuZmIRhRiJe3LBNSOwp6IhGEHBD
VVgPWukLQf4/NLYmrK6Ditr0Hh1mkXET4ePKqV4ds7zhFHJ1gsGFDeX1k+2TLH25RBng++Mx7q2j
kIlvBqF+ROD7U2bM5t6uFOQRYEStd8Yt88RND+hwzqpt0LsC7CxAsjp3UL9EC+9L5KlVO3hOa7U3
mFMJG9dR2ZquFkxz32g6vV+FPosucsR7/LF572vuiQs8M8tkrvMaw9b58Ip7qoyq5odE4j5t2US7
IiTVIwekDaspiWxgcm5p2AbYQcil3it9tpW84XsjNdnpw9rDlnX0naPbOEtj6fxJwQyf2B51CPVL
JOp/8LtdYVn6dif+SGsvWXT2IS6n/zNhznZax7tZfuC5NVUDmbacFRO1WjPecMksBi8qiga/52Sx
M+E/JFrsprMOBimn95H0hbypfbL9D99KyQLdc7T4sJ2rkKdeI5+9/+ebl8/tK3XgHZAgZyPrMNyg
TGSt+PM51RrSsvzjIeiSbxZA+HpJLPirDNYJ1tkjlIwiOVRKx70wEkA5a+F8+WbsLrbtXdegBTXW
QcVdJcC4txLGDOrl3DvkUh2uR3saAyU81jb3ra12m9nvslcafxXNiDmHLVcv29n5zYjz8VPcOj2B
LDs/PbwX8XEzhtTc6YmA/GRh3klcjB8t93IExdAja4zfW0vYNe2lPBBno4aMsMzrqK81v0aNLiva
xtXFrGk4Kd4yHb0Pd8mnWPDdumZl4C9xUanTX/sV+3avJoBQHXscP4Z9mTgKi5jy7Z4NVVvM329b
YwgORGCmDxv4GurpwURbiTS2SEhvZsMtmMcsBkbaJsZsad6cGMvAd1nJaXJzY5B7zMiDqPNh/aW4
CYsce6Tqte62Gs9qLvXzV+Gp8GUHqj3XlDSwrK/zXmf7jFoGZu6oQ2B7IwBzkp9pkWRZQ2h60k+m
zAsc2KASeRdJ9z1Afpa15dKvMpuDG13PScO/W9h1f9PjAL5emXYd7x/+ma47z3p96K6GJjPU2Oza
1vCD+PJydCsFq5EAw+AHc1g0WZTQAp1H/m/sA2l3YYcHneTXH4IMNVRFCgZKK7VpIDzoXk0NRP6J
KyHbztL+w+ZZ+ub2Jyw69diEC3XdZSlqsDpLqUnp3yZWOfCy0lyZFsxYuDxmhOeiN77iaWDIpvgF
a2hy5uVk7sVEtbTcu0oMAKi9gHoUvadYK0c5yCz9SVnBR2iQC4BVveWfLHAmpAfM7m43rcrb7ufK
XBK5CuZJt0trRKXGsWVWs+ZY2ppl5CRKCvlNFbB7yjzx/h3J9NmNuWhWgxoVryA8AIU4x+BDRh4N
sNnp0yiC458gVfDuzSDKHLOZdn98IccvDJo8j95ptWDGRnJBdf5Wmn9A5R+SvuIWkj5Jo2Flvobb
1fl4J7VjWWDHN84HyBxc0GhdpoHvvi5xGRJdCPZpYg7ejSHb7wJHAHZBhFL/4VVyRu9uAJ7nZiuO
fHo1jnjf8rAYB4yQxaLtfduPxahfydE6ZJszAUVxt47cbfl7g1d6syTNcp0STXwuCSQffQ3K5q9Z
D7DIw5MOsJnTQdtwQNkmB4O2cPsoP+NtOk+EztB8jMCgsdCovkdzy8neKbAqecIFh/tN0K0jjBi0
Z+1SC1VvLjWkmF/rECjpnORM7xI26QpTQV7lPEZh35cqqhZZJA/IvNbXZP6B9VMaAAsO6Jv/+Y7E
7CfAwr+ApnI9LTR7NZFZQBPoxjPD+RpTjhvL6gc3N6x9DeUuxpnMVVHw7k8qu1nT+qXaKaZukxrA
alJnMg5jLDY7oqRJax1AzClBYaI7PhglcO6DW8oKXbJ//nPCveGmP4XpeUrnuYg1TcbAFmRKyoKZ
fOLlwGUeGc4zH93c6168zC1aL85aqoEMeHibrnZRmbN1EmXKC3fIOTUSHgjqp6AaCG3HT0J73O9b
CBmoD5rIJKNnp5fAmEafkfwfQojuLFr6BK8CP6lbRIgsYi5pR7eZwdU1KurfACtg0e3mlS0BlQIr
LSIbnR8kMQlSk23KTi7i8sTW4sDan9v7AekApc3Wh16uPDgLJnmGfJWVRFEJXoSp/2gE+VVYKW3O
I6eu4GZoh6o6bUsqUxy20dZIrbAjunM0RI+JClubtyEswq2ssQGYHRARUockdNJ17xzCLzJmcAz7
I9uNGN9u4+/hQEfvIsHSC8VhQxKvtszsSMgwzYe7+pTK/TmnuJ/6NuogHsZVpP8fFXpa81lewsCc
BWeu2/j23QhUdRIr6b5Ca8YtcD1YxKb/RJZHjf20NlaRtIka1fX3C8FPd1r29o8JNPvjh0u2cmvT
Bshr34MUs1NBDVw+dvAwEJVYp2HC5Cnt3npWj1uNRE0izzFqTCo7qIPCNtw4UJiTKTrxph92rGv4
oiXHG49RIR/3v1QV+AMZ1zTbR8d7Vab1JNPG53YF+4gBdaDzbdP8QDSPxhOR2tSQOWmU3urJFVpj
xQyVjUJNBQ9mxzUEo8QIkrWg0pyZyMS99q239QK7IyUUsxv2N+ZkUuZmosuRpI3HRLeGCxtpOmnM
ikpWKgwgo81BM6+NQmKBabXWptSwTyOcpIsovfNGY/+36lIR6ULQz9zUaY429RyRWCBOgsqpMzOM
HGTjL5VqgBaE9/coQ90ZMcFCOfibypc/XGhxgVDdq9PjaCVE4Mpk9PWGWRVQKyDLB+L7IbRXOqZb
pyIQkC0RQNJupN2/7T3aqlERaRKEqVI2Jgkv8FTieq3uCJ08RDhBxVIAEv0Zv6UMme2tMVKjOHEq
FqSc8EmqJEJTuXxirY5gBQj5/r6BHto9Ahi857ha9e8foeNYq34JdNbB/9vLbc8kNcFh1znwAJx8
eckLGQ9CU0tvsH3J92uzEAUe+mPEfpteOjNUSSq1zvtEMzZKcg1XgGTZ7OuMZfrTJaJ4vmRkc2os
sBXI9qngrWyV5UVFhdlaEt6DVAc9CASye1koHmphsPR3XlzevGeGU5KDSSZAs0ADpw+0xisRVWwE
XvU/FeCnphzCUzWPk13U8uRcRmZv2G9nxBqbImwq91Ib7Vbw/bxBGUeS95yHTQmdsklQyIFHEJ3J
5+7KdwNaBSMkgU4xoKDsfV98EAnlmhJKAiCQDosmetzBUVIKzqxvGf1tx76a0of/NVNtkvDrMDfh
v3sYyTeNmb5XyP6wqM/syRNHMzqxnHtx8hmEfKL3fAJuR2ZuHXag+Qt0bv0xgUUwTM//oD9O5mgf
h5VvqsYBWdX8NkOSmhuX11wAp8LEfPll8PcpFlZxzkyVj4vhCJUJMSa18Ru3KRYpMFIcJXUPilix
wtlYb9yk3LA6mp6C4MMYbfPTWh8+d/MkEoxdDW6mIfk8qf1u6bL4He1WPJDGfPGZuztqjsnsgxZa
EaouhgbdN45B8ojKMv+CR5j1VWFwF+qrDMOoRQJRMRvO4rmP0b+RUigDzJ51zemvBVx+sgSTwk4q
dgr6R/rxbQkK9xaEXvpx8d1ma/BM2XgJKVyJl9j8R8XjSTOhvRmEDWUS+jMGBoxdj57BNhNWrP9Q
ud00iWIBPXv/+lxYWjlwruQFg29uXYI3yD01xwVEkmknV1GppDMzawgIADk6hmE9V4YQO6T0svum
8kDU7dkq6eu/2wIdwvIn3Ok/yPN+Ybxs6yKuREh5Mq+A8tUdmrkCTjB6M6IfPZ4jdYFBTbRr11h7
LyIbkeECfmH9HJdGS9CHVaI0h/9tg2naCAhBvrJaQLr5/7RNhjOLpFO1I6Q9Jdi4Q7ZAF4V08rV9
OOFiA37F5JtSd2rLEZ/EKoZgXBYvZL19R+vk+Zd/N+uh95FPsva0wIETRIwKeqOU2lMTeK7u69mS
DWJbCHROCPckS8OTYn8gdtz7cw/lNunUy4/SiU/yW1975g91kdPwR3e7dXaGtYx5LnL+ZARYK0lY
oNT9k4w/vayIfoI5f45eMpGvU67CMbkH93XFkaQ8rRJZvHjafcUMbsTaOkdraiRRvDCbJZyXmGhc
IjTpA7EM3suGqs5xsxzCWULl768botBES8vKgGMBwItbPigBCIfzfiiZYSfZcDnm4aOnBY4iQiKB
sGDlhXrIcawMpnd4m5+2N7maI+BffcAuEmTUqALBfFuYV4fj9LOjRdwdKcd61pSUZkUd+J1514vM
KW19up0yqPjpQ7m/+y1w65j5pFCYSIFFL2lHnBcgkoBC1+P8g6SKoJGKvomuIk5veaPqQiFtjXhi
YMrBrxKgtiVOSg/jUsf6Rvo3HwgDx887RiY2G01rsr0+eboH7g6252G4kar3VbxnrP2HqOyMCbsr
89AHY0aJ3wFyZqz7qam/FSSymE9iEmoXqqDSokJLDJ9WIDCbGXw0TGrY6eTbNWMwLUvKGvjqcCmO
BLmMmXbFpBkBSLirb0l/vH9GRHopt3Kn/sUA8tCYKNn+/H5fVg2lFZOxHi4wiwfKksO8R+bYDDpW
c3vJcPtXp/IEXoxPJGe9uZ8uHjC2j9TEELER/wBi9Ut2Yuev+NEUyBhz0imuQsVjiESWHFCqEKGU
OFUo6SQyN6asoWw3aVgNLdlndG5pF0hHXRc522FRBuSTdI4zIyCC1AnaoKrl2d2w6/RLTAYYVOIW
ii5O5f5Zbn5PaTLTwOkxF5pQJBW8mUjavyMvL6NCxBXmQVhHuHi2LxGdRUTdpDf8dTE6BQ3/iQxa
fIkuZumVp9jj95aImqM6Kx5CxOew8B828Rrs8Uu1t9nB4re8q+iIsT3XDmmj0+CgE0eg7aq0RNoZ
PmJ+JwYbrTiBuAmt2jRur7gN6luGW8UVIkVXJBdKg/qu4U2H8T5djbouv5CRopGlTg9CIvDkdwpO
71QthO44Xzo4gXFl9WI+T4unGUkuHdBxiOTUy33xZJJHaJ61yN38OAbT0DVO7BBxnMq8gy3H1R5g
Gu9CxNRkZoEpJm5ByGYtJ9aO1Mf7dgp36Mafw1TH0qCuSQoDwmAQuRDrs95JSgJ0svi24vT8Lpgk
8Mo9Rs0utEjmy1Sc059dPV10K3Uf4Vo0IdLbBqag0NnoSK5ySQMtO154h0+U2epq+ED6O+VAv0Kd
f6loSybPF8nsEU6KZstaWpDegqw1xNgcoegTZBcTRkqdsL59Tw99MBs30eWAVbCBUYkvP6fj8MX8
y2WN+qLKD1eOymmt94Ly3KHXpi0yQbUrEfuYrZFAePudQjlT+6lM3+Fv4MxXDuXPsFrGYUjP3V5c
qx4LWB6AZHX82Glpmp8C0mtj5OCKNf0fC1rjBhdKrXp/QkxsSwwmdLADnXYXGdkE2gWRD2CV+Cwt
/6xlg4gjS+mgO+ILXG+xM3XZ5fDzyLYft7q0m/PYPA066qO9S/9qRU2i8n1CvurUeCGgB0Do1Ucy
HQfTOK2r8lrnhTSbcIYLI/4IOpOMv/LsGVP34RNdgI4QEBHmsIsZrNRS0treSwU3MLwQTebgWAla
PCfiXemEky7+LIgcOUcyn21BoMhrT8MbSFiYmEGHt9s25BwOOXPD+lnbmfr/PcmefSJ3SMTr/hjZ
UaLoko4jfbotek+A5aC0vNadJX3eYKHZjy8qB+CenyHZ+SDpt5cqfHphpnjX66HL8CcM+z5KTlIh
Grp+u8TMstjz7plb2qUvNMuTHUoheiAbQu0KnDrgBjxP32g4Gf8EhxCCkxPJbrR8gEAlVEIqlCop
y7nAI5WKtSzWWhzLHjUXz1KqmLHuz0M9qcYX9Tz3Hg4Z6BkUgm1GrbT7fBHP+a5HMh8SHV8faips
y9IBYvUXklF1A2E6gu+wSDCGhT+COIXS5/sI/cDUfHkGQjJH25GgUVxryjP6MCq6B6MWchOpqDWb
LRFHcnt9iZsS2oq8Kk/W1e/nk9P3Ie3x2p2I9TZYotPXtII0X0hE2JBWMH92/GTxa+CrwFbbvikf
5wDdKifmBkHgZKwpIL4rVyGwD4S4X4qd1oEnraqoOKjPYIqOzxbfDsuqWo5XrHdQWt+ezrGt8V1k
ago6zMSfY/2SCbbqt4FyRNRXmS+loh3FCXvxQQgaB339AcdmeosvnEUrcTICBhMRI3tPs/Qxs0vY
tAjvkbzUp4MwLQWgUL4cvGTpf/EkhXTPXIZFva+4UMaacAdpTdtMzA0kgqUh9iXTUuOCZTJCuL1O
vc0AVmZtjcL1pDq4Gq8QGyX09XvlQT2xnZwD8TkUF3U5u7MbUTLsFLIBhhkvzV3ewCTnwzlfXyBl
IoCbCXruVnA8RAtKN8ziphFjKZOCydHuKARcn1y+Qh5/hY60kuqTwCJyGipupGE5KsLg4sWtfpvL
PjNACQPJhj7EmNxU/OOyg7Be/07rEwb2HijvxuIyNtwaEiqJUuSUSFG6LX1+880VNobBnUAVQs7B
DS8rk1g5f92KA0LWTYTy+pPLyIgEGPE+GtV5j3oG4EmIN55pL9WvWH49pwOowwnc2jHfh6NUQY65
vGXrIlyjN0zpOGsQvBvb7+ERgc/MEhjR2qOM2cBXkhJ7AWbcwuvPfO6SsjFxcrWSAJZ5y9J6NdIH
ZAwFBxQviK4ohZ+hGeHnWlr6pdSiAgnrBn/Lpdrd1bbBOAga2G2maMSbKdYCjwt/5E0J1f/W7nWE
4/6q7tofr2kVJrbSQTi/NgEVTPS+3HkCMxIAG2MeZml8MWyavhdTvNihcqeaFJlJJ454NVsWHUWx
gYqhnRvrczPTR5BE02HghFjULMx1+mYE/Tr1OpVCNhhWW4tw7PFU1YHE6TsqJIC/IX9Owm3SLwCo
uLxuk9OtkH2o++bZJIgvTjSl3mMsh6yZgnnNILu62aAWy8qPun/lPDsax2h/RAyIuBRuncn6ud30
wYyt7h/NuSHiLaM2lbiN55CN4ZI+k9/OGdKvgK18SOSqr/7zShsGJ9bY+ov0x33VUHso7NWlnRLV
8TfA52Fp+NMKGR3F3VV1k1enhE+CJCNWbwjhqoUNEPX1AgLRM122fc0hy0GsrGQd90oaYpkyg/ih
/tYDKt6PEy6I5NM6/ivHQAACVoBEVQDyLxQ13y4G3n+EfL9gbr3Fxcwdz5yd/OkxmmaIJrRm5t22
8ts7F4NJAqQcHE/4iza2+Bw89BRvlVi2Ag0ARunzmn40hQb25b+PFDhWy8a7EbVbvhpegrPIW/tA
JL2Ck+MWCeOwgHRB3KzTz7u9fJ3BF1Z6r1FY2gVXPYu7Ee+GWQbXGPllE5EbcS9pkswepiKfx38e
3lg9B2z3UCgkSDaRnseHvb6uKbO/f/7I1e60+ft6pG1tpa6aR5M/F6C7VWeG64vR28leI2Gjfs0/
YIFpevYeiOuSpTufg0Xr/IY1K+QeM8iw4H51PIu9ASBNET9VlmU2vunGPzx2eDehQyaeBx6UAaZ1
jKc5BU9mICcxt8nlUAzDZkFbZAyaRpA/zudK8RDEFYc/yu94S1unaa4BI2thjxqgZEZ2Qil42BxE
kf5u8LuqGDURsYJvaMeHh/Vv5hgFNfKv62hdgLOLcJCYrY+3vxw1dRmK9K6g34bokQiFRMggxYC6
Q8L4o3fwoHPdUjvnm0sXZPP5oYVij92n1VUlabN/TAdyB5abW0hgZVhZPgNmvek9ojqtYO2NYzpP
wWMMRpci8nxXbJ/tDSU8L6JLna3IJEgpKxNhxQRyzDeehTALFRV6vLKr7Ded1RxqAgJcdjXwUXtV
+snKC1WC8EhEWcX32ub6Izgydw8X0syZAQZWaOJEUIvGw4E/UvODVqyWO4UoaCBiEFWpKrRG3sZl
pp4yEzxYdr7ZDcLCaNTjVK0Ng5OxHHx9O+mEVNjE+QPJWOTm18oJSdq1S3cweynSG9hKoNtjJec6
YdvmE/AXYOau6KAu38Gkl6gZI5+F5DZQyqoSD2i1GXc1WNE4aAHoMpOZ0p0uw6w7dxC2siHn02Cb
CZ75aUA7rs9BlIBufvrhWPC5UXCD4aRTi9UjhsIwhZPFYBCOc7t17NZXXlgzsiOWvS19MR6zjTv1
RT180b7un1vfzoyA4xV+Mx9RhqmNbBwcLkSzwz0aU/t8Wt+9Xxq/tDTdWmZtffdRXrVOqjN7aeAm
OttTgfvD5YuYwi7rDN93i3utfhgbhQNMr44LXJLKCzhZ/uELBNW0fKy+XyH/12LLvMIVqjoikq+5
+3+7uEBpm1PNVzOj4p1iR4HcdRUT1vQlf7trwA50wIWgFZTZKjKCcqdnXVfJDyvNYjj6/6wORl60
vdrK7a5wDkGpTk/nW9hKyIoygyfQr227ZBom6bg+g/xYN41wWApv15fgzoEm0BGwkVMsABcEy/0G
nGC4/jA9Q4Hg4EsCRLWmg8lZw5/Y/Ppn2KHQQN0ybfW7AIhYfhlbSkMvn4X0Sj+oMOrqe80eHIxe
QiBDHp0SkKPF+qHy8n9MUrmTwfYNC6Sfki4n6zHTdUtF9VTrL+5l2SEMu03KslZX9uZlIEVPgBSl
uooIyuFN7pb0CgfCLb5+JDQQ542ntUgDStbSJvZbRQKZrLRJCr2MStob+vml56HKO3OpkjDUo0sV
en1lgpXnGXDmqQKaq46jAy8B5WKXIrU02x49DCyj/0p3PWZp+vyZ69CzLz0dZZMrsnx1qGmAL4gh
4G4UWsNn55Fie+NNL6vtVnmpx5cCtBcUsTNFtqOVHkXM4WjNd10Sl29aWPz3MzWgOJK+pDVk6EwE
/kfFvYKN/NbiztT9illL9T0LjyMZZv4Srrc19Yai5/iEI2E0qQlsQW76PpyOpqbuU/sWwTw4x5K5
fhtPqV0Vdtx1RYLP+8rpvppURSsBGbLYqdIGpBhWqMZS2WHsx2eQVzltSet+iX0DH4mwOV8YR4fX
59lI6GhgstRHMb0EqxdzDf1jn7oqUGaWIqkTmzkwykyR6YDbmb17zTQY3Esg1EbAvXxlNitrxlaK
qMDwmkhmeTHTglRt5GGDyH3CpQd87Z9C00vXFOFiAahBX/0f4vqkCn/vpTMTQOKc3ykkF2o9Qfyp
Ee5V0vbKAKxlHYUHEsiX1DIqq0OAMpt1K97ZFKrhf36CdOqjadYw98tJp0eYewB6LpquC9zBqMZL
3WODhD6Zc47OBcznK/fNexfKqOws7I/JD79vUGo4oeegGJDMl+VzFo7/XfioXTIyLw+ztQ3xnyOb
Kjrrw4tRw4qDY2F3PuE6qq3Z8K9ouzl8d73Y050sRRx6Lr7oPXzL4+VAoQLPKhgjnFlI8UYOlMpa
lWEt2qnfhyQqkHvZ/s9Qu5A+7L3+0AHs9J1ItR3kN8rzXcPUIeOZv91bz53YQxTnP6wg1OILjEXs
9JolVN8eDEyzRJTnUPj4hvwpEm1rUdtY51qOivLeyvBfvhozi2m/Lc031aOg0Rxvbn4kh9DJC5Ms
b2wsyWDGfwXeaxO0bucwc2qTPOhmlbuUVOIPBGYjXoagRrFxE0kt8JBvW2R9MzvEF8Sit+T1uvD4
M8V2+Gogz4hyu+SYVO9qQvlYl8cFeskJ6e2j2GcTHd/aKDdzM5z24n2ffD6bCd0wz0xd4U7euaOK
6rZ0NFyLM9ZH8Cj4O7/N3iqLUKun3+B8sq2/Af5P0yMJ29osgEGyViywQM8sC1JbirH7UjUDvUbW
tkgklLXV4iHyueEa6aD9KGwd15QhmgdhA7pejDqxFriPocz7dj1WIojX4ES5r48yDQFoE3GUL14l
k300XwQrOhXcv1QkxtQgPV2KsYRek4F4Amwnwzd3x271neW1NavDB7nRkMDc0H2ZZjos6ThvbbM/
mfSuMM7hyvTHEzz0DSyTnEIoc4XTLUOPMu83ofDAluLNbWjmluZL9IbjigyiP0lSD77LtHhji3L0
O0BOgz6sN+Bo98RV11aoOgTbFIi11TKH5tZ57RQzXTLkxLp4fVIMmHxtJ2rs61kGvn5ODznEDSzv
qRqYZr19MmycZHG529MYBFbfnA6xPpLQWn1TGwGVcg7rJf/41gA+YHhVI9Uy9rTV5eWmUeb03Ukl
WQm1DfEGwbau4leFaeo8qb0J0cu+z+P7+CmvWut6TxY5upzCY0ph3l8ZW42hvKf24xECfqTtmzzE
Yv/69K8wzd9Cjy9oIFI3ICnmfzWoqq2g/IUMlQItUERisNlPBTYQOGnlNeuysyEGsAqVdqSAg9ua
XkEaiFtOM/aW/CVHkAwu7D4GpKLnymvsFCcSaRy3AxGJCDXCiGRqrm5bBOde4hb3/IjaeIhWYavd
AlHOIPSSJkFpu2REwmu2PqiQWUroOZZa8/m41rmaLB+A1Trfag6/GS8FKJFHEQfMacAq2QnWkFlm
EZXPMIYx3YEH2YFounEGplW4/Du+m+fypT8w5mt8irb7Wddu0X8Tr6M9Fi8i2bYIWiKoW0S2JQVF
YehyUtwsWGcS03YEamFB/PGx04FWaU0GKvSt+1xDIfSt0oh52RQibzz87nNvDqzumQbsSC49Cfdo
5rjLM+8mQdJc8BxY2yfOJKVM/gu9U1hqNQUBjFVlWveon+aJVNz64vpIdualx6ytyLt7POTjFgNV
3kg/vd42z5W4/mAopV0p3KnLrFQQgZW785fCb/JbnKJ14FHxD/Jpy9kD8t9m9YbiNzWIOWFUoeJF
4GbYiHZ6GNwtBkJ5mElOQOUZA9IGDAXpeAmu5rUReqcOVUya257hFCQOX/5IxbOeGJ+wYdQx7+tL
x9IQ+I2icxzW0zokos91zBL7bh6iPEAf9UURvswr6IEZt/efWqzkLqAFGVGHEN2lmUV0IkFJP6Mg
f/dAzdDCzxoVk/u0W8/Fm9tb61Z3qO3nFqKvIuNLL86zq4Q9APGNh0uGNCQwzqkQBJBTqGM/2o8a
eVLaOviseOBqVfd4CUqxcU2EGmfSFwzRVinCMAEli7cVqds6OKyrAXY9dVbuKg6yvKCeyRVQcpLp
Thh+RfIIXht1rdcx1amdT0tc8h5MJsEXfV9cQb2DYen9X+/qnYU8FN+LLrhEWfppE527DYPcK2QS
X/tn810aL4Kj+zBxA1QOmV0LyPMmBK8LXGgZ9ZP41d0rsIyTbHqy9ZRGWS9dA+GMkc4U9wdCKMuq
5DpcBrBfHmBISqXre+y3Gj/gyT80/NQ+GM267R7ibnhDY5WuDZFF3/veLJwlICfGwTPEIjI2un4a
DfkT3qEFRWtxrmKVlXXIdNqE3kl9+3DcxHWuoIxjwDdgivf9nxbR1peZJZWs5z6WJsVJ0z2BkGaB
rmx3dZh5CQq/jo++6cO50iIz0zmqb97Cj7Y9eJUoeqN9u912ysr+tH1baTyrsequ9lWQxe4y0cPy
SPpyDtT3iU20smUmEnNtE8Iexw9Ddc/Nq66qr74D8RpXg1Jofvs/y/sJ4g/i35ESgI8PFruM+/k3
CVSeHFWSeypxpJIHcEnnUV0aegwNdpT8YiO8hNIr6JFhOJi730shrrvnSCiFcEDo2SEpHcPymkoX
lj6yUv80xSOgIfJm8CDZHEqqBIkha/43me+NDmJPfXmlqUzQcbHyV4oRc4NoqDYUmK9q85Zaikdm
A0fjIy6nekUVdrR8M95NQftzi+cbzIOy2otbhOd4SdOWHDleBzUFWjTN+s7xiYBNPIb5WiDqiCD2
NTm0xOyEr7BbvHUrtNiJYngbJQsMa66CYx8EKpf+QZTbiGboARD4N7gvnfYE11Loznb5JmgX9k2B
bOmlrPTXo8VZgncsoQi4g86uQUfx7pAce0JwAWGLSgxrqzZr61PjrwepT/TG6uRCeUfO+t789PzX
Fr0MMOEeL2hTtxqXIJOfYeApGY8Aw1Zg1augqZcO6pROFBo6urRpjp2SXnU26evScjej4Jsk+rCB
QQGSWAio6uODuXGe8qMP6TiojPvtfCn0pnY9cFLSSGpwWCdxxAczOiKKwJmSlB+BjGevA9FkocoH
QA1QzKWYQFvgG24ePplXFcVovQtBu4kCYTlRAt4TTEx3QAGnQYx/c9P/viC7sBr5byes8nc0IEDK
MbLuH5LWYOw0eougvhlsKCrbsBj70e+jJRzZXjrf0ku/aqYkcctrov8x4duMJiXLD+S1VZpbTvtp
QdNMiF7/um5JFaKabZ0rG/hJiDXe6MsmGxuPto0PDvenbIoSUNfEc9wFbBpaWYSANNNWLtl6dQqo
ALjRmhnQ2ovxSA8Iacieg8FvvN3mdHS9Gm7uK5a/bmVZ5Y5C3Z0+EGs51rN8zyTuvSopoQGl84Xa
rYvVZy8BjIGQWzOlAXakHl5zBOd60sVvmssPdumCNXq/JUESiPvuELxnRRIsQ4/vNxS1bILJp871
Npa89LAUZuCnxsHo6cEPYOwQ08AMXJI/ym3PB7SZ54WyzkV6gsW5RkqC4cTqd7gEv6K2WNGbtYtH
kf6Wbeg31Zey6ex5pIk840su6VxWiZEuSMtx03rffi1sQIl3cUDhx4nvCFnOsh8+ODODLPdWJR2c
NxanOTHJJueIFa5ioVHRH0AAo5KKPdWSrUCm0EDGit0+2lRgzkuoZPc1CMyvHw7+kxylcGP3ffKc
lfdRL8q/IxozNZ3vHO65tljFGud0wG38wq1R+/OtrJ+GaICd7sUsf6ts8rptTT9H55gOzdTDLPZq
wOtK8HZVIphyOGjZt1yO0U/6l1hEVSfkYYzIDv0Lh+EC3HKvV1ek2ulym1INW1raWJgIutxPVFpG
7xRcIQn53lup5PCAHHKYP9+VENhfEarPtv+gIylcoPlHlEz/2e+A+UZlFABQctpYZ5Ro0t/C7CBh
Lq/YXhA8oRXxLxOeDvHgK49uKv2vCJjDpVpX8Z1GbLU4CCgE4B4NtuAOb+9s3yaGnJL09ZVqvT0p
0O91+pAH0ixLGVST+f5cCUQOBLrE1vSncqoR1SOVYk4W4spGIqQwPRuFEaRlsQyiHBdFJNv0VkyP
zVIwyThsplURtaVGelqfZHJdm2lhlkyps5f/8+d7pGyCkoakkoZec6pNveIi6fAGL0YhjCRPXXVX
3zCX56iX24n4mNA/R4AksCHYKimJ70PYcuMe29Grqbh/2tvRhPMGC7Re1fU6GjLb4g4fBf2jMxps
1opdnTAtwwHF6RyziRYRN9GKnj3iZjV6Zf5H1jxfPqUyBHjkymYlEkIjlS+A5FwmVfhxI4Jx9wh7
x9f6oEPk8VlqyO2NUxV/rw4jSQFdpOqCXx5nc6KkPUiEASs17jgK6mOU8OIspE9EvhI7y2+LBM89
GACSRu5bx0PbJkKqhAUU742m8SRbAOa/x9FZiI2UMs0c8ugGf3EtlEUhqKboERxDAEXCCZbiya0R
Gpxuja1NSn4Q9Fv/b6MB2mB/PeutYwzM4DDmzaHAKzNSP6/qWJu1AmiaZT/2v3n0ZWcFLRNA1k/s
sGQGdsSb+T6KWNLk1CtcZPsvzA++VHcQ0f5OkFJGH4QNdF3bRE2VXqe3cD/+L2qsl+U+6UDM0X8m
vMx/vIZqt7mmqHRsb3dX97/r9FdiYeydukookbMBceuAjdWtiWq22tGtusm4XedAfkje+msK4uFL
Wi+Z9tbmU4K2THpCpjoZe7h7yuzViOjMTuWWFE3J//GTfSqRqxmjkY0kwWZiMt/JkyiziK9dpkMV
gZY+cBl9SHP483eVrTT08wRkSJgLCAg6j3g2D/Ev4PHLmHDQwmyFZGIxLO4Vomchf7goFI1M7FeM
PiAsU+MSa8GXmCCttC4kLdL2wr/TCD4gcyoHwRBLMpjccmN1OFi68leDOtpSs5TvGTCCFUz69kiU
Ahe5xOPGJDGSqyl5URxHFmtP34YkMImxVT3CvozjtexdjoxUWlIUBfuKQzMQmEDAJSaQ2QzrMT9j
Gs5najr1H0/RfCwtxm1A4dnCq+8rT483ad/H96ZoySoMQ0xilYlw+9HXnBUvwXWHwBQ8gkLah3QE
SOSrvM8S6swbaSYoVL2R0pNoRe6vc7NSc7VkVvk0R56uh3yblYUU1iNFgNQh9yBOMAYb3jLBOpFp
rCF2+VldBObySa7CZGziyWs7cNdAsXQehF8P9H5vbVT741E24qDHEn0A/XT+sXGihT+13PBWreiz
KExSOliCc9aXwZdY13WMtKKvau642IAPtqoaOTTQHw0yAr9NpoKO6Ld1uiMCI+awaJdZxaMiBKdY
ZnROKyX4mOZk2/jfscJ68TubaDDJQP8uMSYRtoeTbbI6Zl2NvzBBcXhTlkpP0gNQj3ljCfpSKC5k
iQDrs7PomeXmIiBg47wUDEqFpCPkkQNK11NKM4uJIzcomQh0NpIkpILZvR4aI/MGsldfFExYqC6m
RsY6JIjyknIryAArVTVk060L/WTjoSCziUia7SrH1vVzPivXz8PU/mkQbtwN8Sg7SY79AHq9A5lF
RMWNnkvDA3wKvVdhFlSwcxVdOgnG0aoygiDjl9/w1V/xRRAmVMmNia+4XtSUWR8x9s96MhVt1mmr
qQqL7wvAPwzFTeJJmfBSsChOmPbSlYVpsVEBeq/CJ7n3o8/4NczlLmAMMdNnI9cj6yyiUYw02x3i
8r5jqbzFwJzYiRNgbRi+ZFi6GQ7z2I3xnB5zVt+J+0jsuumYHAq2Cn4Uh8bp66ogGzzJRhf0e/hN
z2l7+sD7zVyjJfBj8YUL3EsU/EQQsb1HBy1aQOUbiuK7s3P7oxEY9vrF1xjfF3qFNru75q/qZSZQ
Irs8ZajyrJ9hCTZa66V5xxiHx5JwYg/wUk3xTMkdie6x9LHa7IXi/f4a8CWyNJeM1pE5UhJXq6ty
7cD/HNab6WMSZEwqi2x7WRQMcYsjZzVxbrMAnb+kvdNheXu1D8WySw4Zn7Jv96g1epUAYSgqkd1G
AyiRIMe53fu4EmlEzWMK1G8fG5EkYIncIaFubwEjDuQvb5qefI821s6zIjHQJEBnF2rXkmcs80Tj
jiw5x2Y1Uv6ITKirGjX3g4foLWMuShVDCqTqUObXdO991wzBjzHDliZxMipG3XtsBJQWEWWE3oOs
2C6xdixMlKT9OF79HStKAiBO9AAaZnmquNzIS70aNt2UXyyXbztu7nTHUte4NmfPnRy53d2WlpQ6
FMOGMvYvzu8ZBbdDQcCqQp4qgN7YncRcuqAXNu3A0Wwymi4MIVEKgfVm9ndsPCxgK9K7quzujafd
NjcHgDIzU+g4jGe1djNr2Tft6/jNg0XfQLcTwn8YW+qJWMzf2Xqwc7iBH7yvGTdgThFy29EHF6ar
XQ3JunwNdcTLi9X4tmzUCCYFCk5jGpy9SHVbBwM0ur2iUQ2nlmOoBS3AHs91VrE9xFjhcyJQoPhK
Fb9IL/em3C5GdzkmLz2AyDXfklElBI/PGCf3c8gkRd7LYtyKxDu3/Hc3Pn/gl06tY3f+ssnMzNoK
nCx1D6vwfq/YzfHwDnby+dfvcptPAV12UnqM/fxTToYFE8hA+/LPcnwpFyGBUY+4jBV5xtw+ENCX
nayfolNkc/PWU/EIfQSNyrdWGpnrYy7oXqOXRHvNgTGP2s3HB87CNol0i4159tO28IyitYzP43Cq
/3Y7O2KXx6pGYg2m7B/QQtv9HTm69Lg7zQvB5WOpA9IUjlFOML3vc6yh7rrd9aeNDEK8UU/kChW0
44kVQ1oUVks5euGys01iFB0XFgO3Wct6TPaI5AHLkoC0oAeRnjFClgmgrdtbZNVbt6pIDKNPgM0Y
dvcbARX+173zSMQFICwxU59jlSyRcsKF/kqml+74+xhzAgH6OSAUWkrJ1M6mTLHpg4+rF8UGH9h1
SUu+7z3cecLarhZ91oZO7iyfTow4n1oR3EHzb9p52khWr4uGolIXARdlOoRMoQinCdea7RhghQr7
cj3Nr9jCjD+28vhFZNaWoBiX3YvsRd7f67qnRK+y22nctKNofvZzSfMUG3J626T3JstTTjjh/jpN
LdfcKeTgj7v+1GTrVypeZpfZ9LfYBtKJIBw1NMpIqC5Mpgsfc1LAYmpvmihB/aEvjhRzDE6jIaCH
S/0NvCY+inPjIYQW0C3EkFC4Qq2dDoJypouY0wAbNxpkoxrpbTpJV6bDc2IQNAqg6vHQA7dX51c4
+i+KDXB+1+ceL+Owf2mKGcwiwg4aVDXceuGOQj/k4ALlEPD6qDiqDtwCICtfyt9+e5B0o1Vw8KiM
i8LQBpJJlb1z1jButGG8N5x6t2pscwdFgJ309vxvEbqITLJLdRaKaVwcaMDN3RZL9gUoDk0Qrqxq
I4bnDLIwx9KUWXy2aUlg0r8vm9IOT7yyennIm26Pwl9KG53/fKPzbJw7jIYNEIKuirEZDqyF2HZe
+QaZZa1tT5lYDlhrPlPTdW73y7y6/H6JyetwMDLPrIRB4MV6a0TBTo0NJdeRf/7umVVAi2nNBG5M
MzwtVXYifNzuCO9VFtDht+i6u+3Mv2pEgYgjaKtBx6tBDX3iM71layeoSDplNid7z/LWsWrL1Wh4
lcT4hfXFTPJP0xV1g+j3OksukRAHc6pQKryUyTendELK26LTgjXyF11Ooflv67wTxAUcBTLDGBH7
DSpSekLu6w8m6FMarbxVKSFKZ4CIN8LQFMqeHEKrO1Q+y803qPutochB61TZdPZn2mkuRszIuVad
tJOp81tzgKQtJxnn2UmmQmG+WxTmIY7YoM4vy2bBUUy0nseAtydp2camXCPRsHig8pcal6Bmr9In
q7pCq4lps3SLXEidEDGtbjoV2Vu/iRTt0AI6DA/1MJJpnifRA7JBTMlkchwez1YtWak6wCcpdso7
ylL91RkoMG1jm1JZWpJRXofClibwm1suwzGLNW3KzRJyMLOMFLIxMqvI1rCFDw3RyMeBfJGgd5i7
HhDT0gwgmuqud1C2ZTS6y6ifwtcZGrV7rvhLQACDhq1UloWNc6zdKC8I/jQwgCn98KFY4i2//H7v
cpZTte6gLUNGQgeu9ftTRN2WtMmrKDwE0FAge92GmYarLFnKDMLfW4ueMIVnXFKKWgi+vmElCbY4
s3iVxtRvzAZM4XZVUvOfT7M1Q0iGsBPC+eRMHDQle6a75sb7xrtnW6BcuFCtJEDu62SFi5nQZd8A
jcY+wmUSJtbyyrMQfpOiJlte4fIpGcdMry9YXOJPISz0uo2vEcq5dZRUoaaZvkt2Peq8nexkQe+6
jbeW9iNhTjEKBn8lY/QTmB6a9pJ1oRsgmZsybnc9+Gk38mbJ1DIF4qCtJzn49FRqGse7evuSi2sW
Qe4gu0Lp1GgYM2W/mF6bk4g3EAmbNTVU1e+xDE/zDpCyRHGYPlM00HWZbvlyIGsFHmw9gxcuK5sQ
7IJal0GKG9hyyrQGG9RLHS7S+t3KQN7DTd2wx7B7kja9a9ZMHO7c89vbxOBxmNXFGyqX/u0bEM9K
v7jQBHGHOTLFBjmEoRr/1c0lFsYSdpRe2jVDbzZpggxKVDh0zrPkdDNFNp9Ro6TDWEtI7cf4npPH
WcjCXQ+UNWZqdK3Ua26TosYntcQpdKWZx8z/WaRPaBAPz8YNtYXu4MtislCLkI3CdboxA8Xq1IqU
sLtvebBjuZH4mhiFeuoHlTuBXsgIFXi23l7SJmeH77K9j8lev8zLMmgk+ZvV5wa2p4xF0H4iyBbD
+NvBlFCQLYkPvICCH/gOF9cL0ZkWApH6StsHO0WNVUKpkVT9yzcbNO0YXqFhykGE1mWnimtXvmLp
dHrx8s6nuSPvZ7KA6mBu54OQrlQ1+buRksjQvIIMz4KVank4r/zcfDkVN35OLEcYGxrFIdnAOPOJ
RZPfaCPRwVwMTtb95pykBX1yZVaeCoYSv88i0cNIuKLYBBt+DfDI4jwgS93+jHNYsMdVJc1hjErl
oOeoHtiZ9bdyPONgy0AmdKygsymYPmOCGrwEOcN2BcZ9I0+y45tDROpTAwav1ztzfp2eiCDhx1bd
JxAq4NaWL5F4nZAcgNY/zMIQbhvNO+QruE7NsrBoxTCIL9gDTx/OG4Hkh6i+bEaVlkbZmT2P9V+q
58KLdpTDwc0j8QaZapQCoMmUB35bUdfP9+sz19RaFs37eeNAYX6SPS9GxaMiHoLUCAWaWtCkzkGb
kmu/dPlMS7G7zvvUWkXRtIMpodi+GrxX+CBRdxcMtfBThk38SqttpRXFW1JEc89LNxAJAbGAdy7m
tCUu/0b6guvaV+7f/IqA/1KOLPZ35KXgI6x9P9gnjQrulpPn+IwTHCURw9YAo2RbJP2dR+8CRXeu
i/d+cI4M9vJ3tFuZSqTvBnEWPOHUT4AItMiUypjJjkpN2zZKSvmyj5ho10CONzaQlvUF2gXH3nhF
SMs00/JUMWU3am1G5SheNSfJrrfhSnpFJ7pyPsN8yGHmktNdWQqUqCX4MV8IYB4ocBNG4ZpQZkKn
xq2fAasHkZrno+jzdE8YMXqBhYAfxDNy1zTYRoOh/AsvnsMIjAE7awhxbl6sn7ynFF1XPCpmM5zu
uC72ExAP3LbWbcyhi36H12HcpvBtHHgEbmJewWE9EFBBx1QDLbszUgNM/NunsSVtZi+KHQxVynVQ
HjhODxpGT2WkVOa8kUcgGEavly0FYtrl1dcQs1ZVw5uQmd4SAV823ctkKp9LwSrcMZGMQWgjmdzz
EAxxHOVboEP8C9YLXq9Fu9a5xaYkorFkNQzP+O3ZS/27+rKQJEv5Ml3uyVoc7MEuPor0VxR3S5z0
C/66ZLfiahU7yX+rgTIlrq2faOiVlTHsXRW3mmLWLM0OlxhCB89PcGGTUmVm2eVOBnO+LmyqOpGI
mP38ku3LogB8wQgQz6Yrn3sze58c4tGP4wlq/Xs3DOgxprmGdyMok7h511QlR3HeB5aZzabLdeBD
C2DJXieHDx+5wkw5itwT4TDQI1S1vq/CU07yvr3zHGgEDfdP1zXWR2PoHEdXWGp96xKYbPsTzzWL
WFBgqXvzPSFfybjF/M00jjQGn7veu7wjaffUGsKJJ/XQDt0KINArN99zc4zV9772slaJTbR0go2T
ZKjfkJT+ss1HX+454KC6na7qkZ9ik9l61FR+bprCeycLVa85KTDeeOHHMlmoEUYAJMaSAssB/WxQ
wQpm2Gx4pi8MrNhfhhaDZNoGupPDR6m2PIh23lsgU/xqtpbgfj5xPSIqV2LQ6IlXAwTwPe4EzwO6
nvgaOlH1bBcyeDwFmLSj/rE0wFte1lk+MwvjuTAd+8q8Tc172odLceWMGFLeYx2lV6Xc7J0Md0jl
lS7n3d4i6j6rOso7C74abN/RTBvoh6JZpgAVkqS3qN0IP+OMkszC+0mMS+mMDTWw2zeiICdLyKrR
ANIV22rR4T/dkw8+ORm/POuVeigQW788VoWryuLLDzjyIQNSZEQ88k0/oKS+DVuFfsKf+s+XyQCT
pqyQl5XWRZKnt7ERZ/ZYHVtwVx5GVVuWTZzuxgeoGfqfNzZXpC6PLkoGe13dNgNP5/oRG6Cy4SOC
G3XshXsTJBiWXFhFY4LOsO7xjOEgT8HncOkGjG/EYyW0jK3nfB1M4/HiOzds5ercTHE9YM0l8mn1
l4RMQ7jLJAthLghlhmApI+lFjfzN1MQNfkDLs55qnGpOba4ArbsZb7L1LLDJUDzkc/mTdlaOAEoQ
8XnYYwSh1+qpf8BlG4LDjBA3Sz/JukpQoXq+imhxp/LWOL/8oOmE/Int2D1X/6EL0Fp8lHrQ9oPj
cxfv6d0X7SvXJtZuK+wAVMUYcq+viNxRanRHzTdzIikt8rEHqnEqMoNL6xdvpkSeExCgPzxSn33O
CL485smUEDrTM1rEsDtNPDWIOiIKfdWsmG3oVeYAxDnaM6niwDVXHbLRKtXlKNDLjnSJvuvtM8XI
1dTHn6Vm50qA5qodNumvKr6KBCzZi65wpyyotWVVUHNSpjIjkIO199EBYQUl/t4KW2HWqAd8E/q6
FiRagrYKbcrwfBXqXTZcOlsAhIeJYYBzZaadq8Yi7Xd9xYiBVdkeas1IKbmuimG9K2lDBorbz+BC
Ihku9E6b4h6NzMjVj32dSwJn0iJEaWNlqii1Y6PKwJVunK34MfrVWX7y+kIb1mogqldexskjDJIt
diaE3IgNVFVYSaE+qzX61I9uzK60mk9JITs7P/FRr/KzbY8weCmupVU3CRtkVd6NP/N+SqP0+vPb
KAxSdThOoMvDT74h+jJ4tjb4f/S0IwYINaIzqtuAvYovYRLKghGRiIBxxiVuJmUyG9jkHAn5Hj+Z
irjEUfnGeKIvg8ad+AgSClhufe4Zg7Wa/tg5P8OhGYcGpGpLrF+pOPzTuI9fm5KCmJabN27UXrxG
o25Xa4dfoYwjq6gg0pig5Utcqu1zB+vOI4xpLTKYFiTJEwPVXZ6vzEgRsAgOH2yv9lBbKGs0Ne7w
Rfy8qxhS4uKQSTjUHpele9WIJsuX23gAPCNRsXMDuYZo/oAQ+7NUl5lmQRjjsr5vpPAYI4W4HsaZ
lbcqdEIVFRFMeRJRZ2Da4XKThvh/BB2v2ffqFvHJn2om6jjjs1dUR1rU6nOAO3VPoobr1Xm9kFup
eHVUkti4INmrwyca6xkxET0ehF9IQu3iey30IdWYz6kRfUDPIvkGNu8/549kxFt5tEHJD6vlHBKs
NtYJYzOf90QpmMNyDOxn5ppl8cVaST2sbwY+0UxJvBTO30pXut2L3LSnL4j92ZZcH2FEtiE3zyX1
xjs5tZEpnyrsrQUGWdi2ld4FYaPRrAu1wEk/OELcTOicUkC1iwdgIjp9WWJHUuoEdQaFT/hdutFI
RQe1Acw7LgmUPkqmVyhQ176lX1I09lCK90UvaFDMCjEYscCoMcth58jzHcl4DaDoIalcQ+m21N3H
YUtfHJN6SL8i6GBtncvUT0DeJUMBxjiW6FN4nmw+rd/gCeAJIpCCDYwQQu4V3An2fzVznzI08FB0
IXjsuz03/5/lJmI+cZ2GwJtV73wDm85jS/MXWUSfpmIxSjQHjWn0h6mDVlywA7DnDjU5YI1xMjMO
CELD6UzBjPoY6gHSwEs2lAqjsDrr1MCnL8npr2/B1ObP8iHfxWUj7wOeMhUY71iIu5EUOgLTRMrb
OjXFPmQM4XsuMXdg84GsB+VtSkWEndoAJ+f/X9FU4c1NsoJcL7VrC+M5NhSREDA/3Gh1vW5m9g0d
/R90vbOmqwn6tQhDUxX85dS0yLn1gMyWHdOMUiNJJKBoEScAQQiysP2WSxkjXdmHjPa4iQ4IjNKx
9y0PUnNNruNbD6lOotgp1wUqT/HoeWoujg06Inb9kzrihXrOi7Q5EcYWDswRE3oqL85Ca34/5rTP
4c8rocetqs8VbfppHpNXo3d31YwHBmJGMDqa0FOjyc8k1rHS8G0HmnrC/7Q9VN+C/1ls96tSJsge
ulXdAZ3wHzOhLkD/ZU03DVkyjMDOvXMGPbulT6wyAF53xscBDyNw2UpPcIpNeKLjnmm4I7ctU6hi
uz/Wv3fr4RPbjWMzjck7fNyQyrFLSEenuT2kD/Q/hbGbNUwhgRJ7Y6gDnfvF5Vsg4utPff7RSdDL
b8wMHXuy3hnRyLK37kR923/rWPB9+HAKkIh+D+gPodDWV0BLBJSf+2H1hfBkP+1sM8pKm+s0IpgQ
biyyAouBQQlOhnAikaYViSwLaAsatYVTFlQwcc63UR4P2HTGEP3/iAzsOJxZEPbPVE5GcTXMNe+n
1iaH+ZAJY6A/GfGfDiyl5U8KYpw/ly13AKD+ez19zjRQ2N8tBA17ekbNDj9YhFexhJ6hZJcnKoN7
QBpWilLvZ5GF692SUDwOfDlMFLMmKoVJrhk0lZZX7YAnQjaRCfSMATaA1MhO59p+K+M1oHfcWz0t
0RfYEolxX8C6lYl7QgPpKVADfBr8bvW3p7aFTrJR8+ymvq4xVJoGAv4c3CNsn80N7ZgCcDzGjEKX
mXPKFggLYnTLUv7CZ9H2hi5kFA/NgJ/rp5QCGZixam54uE5zXkpDL44aQPa6S3NpCPuE5XnTmiUR
8IQPDVLyXM+q7UiZG0xuMY9rJqgNFPy6SVE8TF+m8yCY9iD5ajz541uNprYo1f17Uj8g7PMEjV8m
C9FTHK3OL8MP0VLgQfGJuvmAxsz8jqNUB8B2Do/WSg8eBAcmAEh8kAtCbqxFhOC39mqnINoHfbud
ivTbgqM+ti2acBNkR9GwPVuArDVuViuE5nHg4dIwXJ7Hc+/U6LL9n0KkMYGFCAcn+/FYM4qdf20W
Unu2iozjs8maX+MmeVslfJmw/f+rdrd4ZoaJQ9fVPDYKFgPNMRGkCS0NFWAtyMh8zSqGK27uBr/j
C8o9civsXKJIgRbaOgTSNQ/TqohD5q0LNe9Erm20c9eHAQQBvbQgmXkSb5X4pp6kCJ45nYWxKHAq
vnlTsPD8mKLRjzl3bh2jAxcaMoUTNktgtRqkyMXsCBhvcphHTlVcMh/I/5pB5ebqpbc6Anc2ODhL
uF8bzMNsvonKAgJ0q6u7xOiV7LpODuvIUVO310BmKKDXo/h+t63HOR+8XiQqLWyYituVeqPyHmj6
P88OsH/pKjGbHxcJ63BmuwPja1JtYBwjitOJpAyg3Z+g2tigw1Gi5ISS9H8SiykAxjMUyPbToqph
+xosLlg+tM01GIIwm3Mq2e3Qq/SBvVuE1SlSYlBYd4jyNBg+eR0aokbeDZ8FaR9Em1jHS2LVHfdh
0pCXXVggHYL6dXoHpzxWbGS6MdJdXEQCsnzhPOBFxtD1+EkmlKrQ+jPvTClqilIVlYZ3Sjgz4HMW
pFe4Wzinsw5E9yd6Z9mXf8DvprqGUORJiCzaTAbpA1ufvDhJRN9NM+ou9j2WGRXimijIkZ6UIZmH
sjyFQX7zLG7m7TsTB06Je6m/BvAUa7RCmqK+a0veQBrOZAGARZlr8p4f+4F0ZnEBg4pXLUoiRphM
CbiK+1gjq4FHLGNvcPOTN+ZXkUgeTL8OB14+9/hatJQCnmF57cLGo93ch7vnSI41DrPsoZ0Thsot
x9dcqqYIy8GnkW4Y/XgCbv5ZbYRlTR+YQl+C78E32Aljpl4i/KFYbWD9dlJddKd+HUZeaxvNnvx9
B2EMsaAKMq88gemyDhfG70QImWQFjWgbI+iHNgJNlPd8cHf65DWgBTEdKgASCahiR58HRyWXUEMP
vBrS+jdlEmxIzJA5kDlWiNL8YU3lfNsjysbzLlPVNXeonlkmPLqCwTINUQnkKS/FoKf6E8xj+MYw
9xu8FR8m4AYsrV2o06VMQbb1qdMmnxzVxFVO1/20fHlpqlvMCYEaFcubdvtH6+r2YTS18XCB34BI
zj4ZLNfwdF0OtMAAiQ8GnKbBwlZMiszmkc6ba5KAFodYKMyHvrf8ROWxprqxGLsatAJuBi3yPoLc
gZmb3qeBpFDuKhEkfBa/o5r7EE1s3XxrWHGZLGhwppd4STghTjtQ8UC3FJMxEx4f+UX8Z0q4hRWS
+eIRD6hGeZSwIql4X4Y/WPcvqm0w+mdYYUSFqPqvPpJ/wsO92fwBQP841Gk4TjzB7f2vruySziUK
WQMwLNA6zcNJDRc+SkplBXXfertxpStpzPf9P04A8il0QrwZLrVaHnEP9NZy0V81kNblp6iG3kkp
xs3yw+uGn+T/iCCwngO5Em+szNxy5ssvrlyNMKHsAHqC1nC0mV8pnQR55J48L4yoltdYiAUlHjuH
3RlxRqJ2jazhgShYrnnoYZuHE59p0jr61BjBC0ds8058dzHTwvA7taALFJtrEPS/XNk1VS3Ld7M+
yG62x/SBZsTn00/LSBFmBmVB5xC94QCrXj/HtV3iw4/5T1dnb/UbVXjBGrxhA11yrey875Cz8HZb
FuzO9vqVAdKel6m+NXZO02Rn2ThKPHR2gW6FAPMxjL0w9RTSGNat1XS9m2oLGuCEpI6S00/tO8/G
EeRWeik79ZfOiCTn474edrZne80gSBpZdL7QiONoWzl4CzMpagegEVMyCMMv8y0v/haQoDw3agDv
3Y0RP8bcMpUWnYiH1cHmyHRD3pVtHwYJ0m25Gk/q13W1qQHEmXysAIoTPYvCSGdwShnDS+DvWDEi
hWxJD4pAZBp/7nY/nrGvZJ7ff1WYRGExHfrmObJJTacoxTxhnBx3wVO9mlnWM0gEC1KIc6fhXEVG
j78mdSLSuydxcV4STNsAOClHoOfJBiS6l8KgkwHYbicJIXGFtYFrFK3azgXSl4btuPX5bezJtHS+
8yFKf3qjHgZmtjqdUODBcVKY1inToUhpzcNOL+VSHSD0erjrbf4Wb6oD9mdXJD8uY8AUAKK1qY4U
SJ7Gdgsc3tm2+a1M26NtKlT/5eYVU2ffl+gmyqpv8W4mbURfCN25PpA7t4isIosSfHzDRitPSmtv
V4mcJFc/N7RbNXFWYUykOq0sPr4eju8qrWbZj4P5xqWfpjSyuKPKVtLUYucN0N4BTbj06eTKooik
gkvYZ76rLsTHn+C3MZxtJ8B6T6nb92cp5H+tlk2ytUHvR3XRAG4WL7CArIqYYAsMwmXDLzG8e68o
znswKTSpJaZq6XEvLofFsZvrnBj0ae/qyuehzVrbQ6gnoPYVBirfdKnS8hWh2kKV8wbbii096yO6
6d6ocQvmaOq5RMNRYbS4nnPVNQSwrt0jwXeijZvoNIvKf4LbLeEU++1021Otw5q6i+9ptyL/9hCz
xvp1Ye4aJ5whRRBYoGgZ4XB4ylsHHaLOrxNq8RcGJJJc0maHj8yBNNRZlAByboLjQRhXlA+1PRaF
6E0Y7ajXRIxRvVdJhoB7dj8yULmLw49vjqryOP1pXPuhJXnGEaY9s8LIGtd6E9Z+HeU4bN52bz7h
bLpBzg8DTbxHUZAWsWNjfNJaY+VbuBOpFNvHakRV9nDi9xYkhXXMl5MAafmOUFQKF9hq7FjDut/2
syioHQQSJ945RVhbOOEuvORKmZboFts4IJtr60eNRcFs9egGHuiBC+PQllbu+/RCXYQxKmZlLsNJ
HUe4ATlvjj6n6jAn1TrZAxHBHjjvw8PYH96rdUXMDalbgi0wpvDMKT0to//9trAX0FH+QarxqQO7
Qiu3AbiJYjBRz5PPrzEOSW/E7K4g1sgZg1PVKWtW5qOF8QwSuQOurMeFxbg4O5xgsmUKGIB4zrqR
3pqms6qF4Iknm9V7ZygcXm1z4ORj96vknICdx9Fr8nX6x6hq+VSffRCaYWLmXOU6QNoclOysM/N6
fImCEpzEFUDJT1jfISsKW8mpLMVswZdgEVjituOkTvrBseQL/yvKiqsbCY7DnHpRAdg6I+1iNtut
5MlYFjIFroaWWcbNQjTgYaXKoMXN6LT7XQVCbG0V75xP23KK0/rkzASV0rAEbN2XZItkFGtGcPfl
ezB1ABzqOWiXPYEQtI8vf9NBQP1mNpXq927ToGpygAsIDZ1KUOnNcD5KDkqZYNWLbQSWNV039Ij6
Ejvd8v4lfevanJuBsf4X5lrTaTuOS7vhp+CKgwcDdwrokKMFaBK1GwcWIl7TokiKXqJgIIBQ5x5+
pWEzeFJGpHuHzPAyQRB++rNySCPzAVEoCKwpTR1ydev5+6fe4T7jJ6zR0ce9FjNXt4as6RMbKk0v
K0xYh6Orj4GAT5mzUuUFyPYPPUDTitYCkOMX8LWylSmx0YVepIaEVr+XUZyKw2s7zQxXxAsQ5xnR
l0QTZi0nz8unzxTFkpVTVwA+3oGkng9GOTwwOeF6sFAt0CRAa170SJ5SX+5LI74k9ImOcmQy9B0W
fsAKLWk+nXOeIgUjSzYWAKW/Jw4leTjyS/vD3GC1OJkViZBzOP7mJ9ucxMwGVUbUM2sWNAJ9ij+h
lWZspls1Rp8NUv1QojzYhOUYVsDKFYZL7kKfOqgkRYb0qcSadlqbgN7Lu72ohpGSSyStwTxsdy1f
/nwzyZTTB7/JO8XIxQ1+3rR7+IAbyAXxC7AIZ6VkRd2SL2WUnRZx/tFxlV/6wTPxFjzKhfmzdLPg
OONn7uSxwnKEkztSVChP8WohK2L08QPxfM7uSAwqwZqWILFVj5ZjHKm6lMx4ZZKlQBP+VE6zE/Va
EM7VQnc25jM4gBFIiEvEI2Ui+H3p8cyMpm9GJU1I1idW/6hZEJegyPLCj6ZmhDHYOohlS/mF1C6U
CajbVlcKYZQUMkp4UFfeuMf9KQtgaR8nZx1uYlqe9sth5Z9G70W4hVuHgmtvVDz6lUUdtJ86kF1l
nng1v2dSB7dDjXzEK5TgRXWZGTlcDFyh760mwx/W6fns9PCvCbOlzAtbYoaPD6q+5+oyANzVhWlY
ZZjNoTI5CaljIlK9VwQn3HiHoZiUVMvS/mlGl/kk2KyVHRS7KiorBV0zKFw84hivSNWKjVcU5mdP
vstmIxxjfZqdH7FDMBtgsWDzwEeflEEuXBcbAdPBsbDBIrLzTx/X+YMWmU+gvq/+ifrj3DRgaKSz
i7enTB/iSzoN7ZBhP6Ghao0824umEuPsGRycjFXBHJRtKHTOR9T/h1Tg3xORKdNA6sGl0xxplhu/
uc5wwycuCTc46yttWb3gfbKSf+haRwIs0/jRS7XntugS8hwpauIX5V6BnOi+SnmgFCLgfE9bz0Mi
NlpaVFNtmucYOeEOUUS2abQic+Ur1rhbRFoChOa64DvgdWqDZrYM15G0Es8lhiepu4qXQywQUz0i
eQDz/gMaIXBhSWChXjOWfNRWpJoUsqRq66urz0oqt2HG1uOylXd7nOWQwOxKsGKkhsuwzb5+TC+h
i4ktGQU8Ua+BGVmR7K6JXWMiBWIKcgXJdU0pp8zu+ZmLiqbPvVCvGcQQT13NAyMA29yhJMvoU9OR
hoXT+SgPue3luN5srVe8CFxu9qK9dv33+/VZBjrmcg70Qq2Dq/M959WhbNu1DizT20Vwx/fxBp/S
b9gkpWLHc6+7SHLtG0honvs0orChA7DJfRuorY4naIhs+WYbcA/3M2PJcE13sqOY78Txm/MSg6fp
ZRHphTT6YyTN8rz8SeB4YAgK3HSaFAjKPgCsxDOX0XDs7wRHpbqVKLZZB0b4zooskvPYIoy7FvON
gH3Bik42a5h8+e9nzF6BCDAuiEv1u5laR/ysUgI9BLAHCJ6qxFjVn0WuyNsjt84y9psYGH84ZooR
5Ll6WKk1q0gnKAnUDsn8PxD1v3TPPuQ5RDOSEMrew1vmD3Ryi7KxpBYT4Z2wgPDXI/zaaGbu2foT
bGGgQUqM80MnLQxl8Zu1zO30rsVh6qq7vyX89FUleseRCSvplnkQWqiZN5luXdnMvxnWauNMwV8U
zQWXegbnLOjmr3FH68zybBD/9Dr8IH4Wa29LNMMugLcCQXwp7ZhodewmyvlB8aeHMgARaKzPRjAs
hV3pdnQ24pyGgY0d6zC6W3m4Rd47el7ogLwe8A2joHvW7tILHaGaMDiFp2ILNS90TnOoArDtNtTF
h9Q236+iIv9eBmXUDMdV/pyzyQ/yPQI1fXj5ORIPI7/66ArXqS1ddgUtGWf5haYK0sGCP0jONI6L
391wnv9NNSG0PbRU/MwvD0APerZQffhYxnq0hjqLuqh7ANFhWz91q0gaSfH2kQDzGUbjFz/3SWUA
O2Eqleekp4fQj+eUpAsrWUtobnz2HCB+/IlYS5dSIZ0AybckL9p31aKD8bT25v5ngNoHZQveWIta
gKCExj6AxSa3+ug78MIiRc1DvEYnakonM/SwhDmxznCnZCTwsSiinZ61r73Z8h9u6e5Bz7s9C05O
N0vNz1wxvyaINPuV35S9Bu8UQiD+ByoW4kk/sr2TPVTZPGW0oMw0cdui5OV3TjQDZnGYkcD73Erf
dZGxrHVYvnWh+10UEr49FZA9qriCQc8FVn5icFAt/C0B8DMb7iSp+wZdptyltm48khzrBPusmMAr
dmzQ3KVKWPPE/jH1SAv6VUu1qyvPaQW8qgVJx7n1WIdM8MWcnUCCPRYvz4gEnFQqI5sJqXippuXg
3tMW480GHZrsACv4KjA/tvqqjO36UUl93GMNKpAvU2V7ci9KpfMrp8Cj+0Vg+cK9AheUUKKgybZ/
oA6FSuSdV6rDWhZ0Yk92l5tnEMzlHLY9B+du6yzMkQfip3taYYLTmmQZGHqKPfEFtqXmKd/fS3me
9aNJYRItbAq+MLx61C2qT+F8EDmeBg9XbxeanB2Cs9rimmn+5YXR6nc4zieCuU4BeVOavad2TpYO
O+0B6hWcLj7hl2Dpx/pgVo1O9NmBwpMpPvBDjgCJx9/x6lFuF37YeANLR0bzt0N7Ag5hZ+6ymrXT
7VXAQCvCYS2zir5GhjkzGwkH3UCrMjvEGGxGWUuigPKLtOHhWtcBKt6rfMxYjwlIUbDikqKQH4Vo
hDlv6CbXeLmDdF6TPZ2cbPMAIieG1I5c3gcH2h5098ajwR/s11qBV+ZMHsE8+kHdtvhVkUNWuioP
Ezz3P933/WlJiBqD78Sj57MSkfufAs6qX9Q72HeKdlOn8FWUdprtHJQDAeAb3Gqym9hL1aOuK280
fuUBdEFib90UdcpZSoTW405N7DOn+H4f8plWPSpF0swkDAUJRI4HPcg5kYABxKlBinGODC1CkyOs
5pXMYAVga5iKH9iLINoCIpBdapw3QQMr0n+1TdOF2H8NhIozT6UKbeVmCdGMtzD9RfDcURj+LHFR
EtMJLAJwRAokbRBzA8gWkAy4mZyjBy6d1fWENZvKA7q3hmxFcaiLkQC+92PHTAZcdAkN5y+8ER19
cpbi7pp6SbtjW2WVNNG6wykptQVgATDtUjKJ0j5QnCJxtwPZQazIxLs/7Qfqs2tHa9N8IstufwXg
mIgNAobboH0tAoduKFQYqUf//0b7LmNbL/BqeReGPb6i9NCh2/ecku1bR8Ggt8S3Lo1z4JxwKeE8
u3N17uT5ThO9V00Ae4ZD8gyoj0P0YBT639fDUCmnxl+8eX7GN9ai6Q91F8L9lzOPNAHxEMQUzDMr
dCfjXV3EDpP02zIbI3tqWBAfa7gEtlljf7otbrylkl+TgT1vEkXsU84AUVs5gf7WPJL9IoF0Qtxe
gjFjRJC6j9qwb7SjUt0+ScKW8fX+NvpyBJMl7nThQjXvSOgDv1kV0IoEFEOdzpwAVK34iYJeBJph
qEPE/98LsmHgPcnRG4huSK2V7LUzDUSs19UTopwbOoyflTp2oETkM4frbEMLzP2hzPqv3XwyMGBq
XIEi5mYTY+9ylHAMe1JJOoFGTItXa51O5ryS6mAlZ1iVlnl9jZgD0sHo9uVHDvr6vcnIqLhVaMZ4
yNrbmtnh6wnjthtdw/lQyAhz1qLNynlNJrhKz/2LqYXiFes9jloGyexYntgjt5bjSp610r3bVI6F
XGth2VqVpaq1hmvj/Bdpbf17zdxgQ6Zx8wlmD7CqZD/gUYGjbnsG9idM0idy1MZOaEFrqc1dJnpM
gOz7oRlI7qFCYXh9lyU2ZBAzvjA+Ti2tIQ4hBUo7KeqybTxIELFMknOzkWhcuNjxoaeTxyD7P/9b
4T4jl2GV9ks/PjNNOcCuEpc6ymuOX5LnzgyO6YgYskOW5ulvURWqY1eZFVEjA8qQom4cIPlypGkp
WG4qLpJcZOvdrUyO3YlqNFa4fXi/Blc/n2c1sw6ontZLBdd3Ygql7sdD7qrUrBhzrypwsuN9TnmK
wdFStWHt6mNG3HpqJitCTBz4244OHm+kux4XvOZOf4/c0ncrYqXFFjb+t1GCvTWvZKWlnlaUFXdT
QfopE7LibDf9qh0/yeCdYdHxU7PYMOp83ZIqXkMhFDAWgRtVhU4XeBNJfIgqVsjAIOAzbaJ5/L8l
nHL6ciasa+vN3gxtWFF6IxLpB8oYu50KsCRhfeOpzO3ghg9DTJBX8P1gMa2lCM7OYdZ0pUX5YSJT
zVhvqTSpIG9b4QQ2EdVH6aoslE1iqhIzE0Rb0vuvRukB29dQmIAVwZsNjEQOK2MZTpRk+F4Mzv1Z
OTlCuPD/OMUI2yNYEzfPggxzqznPkGuMI8PrPsjdUxrktbdRaiuzANqAn7lPCwwQphzb6iA8WJeP
tRtIXAJj4c3HFLRE+2OZkRVwYRnkWxJL6vqyqUn8URSAHPA81zgyepFMhaPh+KqCSZDz2OwxjfSV
KKL9YAMsnlJfwZa1W+Vig7f+O4lKYZBEr6XKmw63tMI833YMjZPBOY4oCqApt641mvBJ8tRs81WG
cPAAQRdPTSR7ou+PXkqTuh9VbzVrdLoaJqk8VxfHEKd8z3Rk9Lsd3nAvA/I9vRqcHfildfVFfNFC
yER/UUJCz2EfTJcjra8kF2MwPW2yJ/Xu10S+tyM9WwhytUqkcTg8pIv+me0HKWMmIQoH0RJgK6qh
B8vN/rk7Q7yZPL3+ykt4n8Kj0ltTl/d7k9hx3gQloxgBEK5kshITAU2YzSv6UiLBbMtnRL54mhhQ
lTZcJtYOj4ZKrjRAITC88bWpHMk+EPd4nwkwlBI7fbV8bIarvidRmnOCOcqetcm0gIhsW3FkDnrf
4dNye/OdROJG2aJTj/k+LQMyK1la1JX5FwyF0GooUxFcw7EOHCsSxJvyIdsAwqGfWObIo+ipWe4I
4dGdWDx1PVHlonGlMRxMV4tbABBqr/fLcs4TrbE+L4UJtjA8cxsSR1mLA3omxVGkDW1ndBj8ib+f
/faEEnfbGmI6KuJyHWSQqCjAcHKLSG+MVuLUUG8bhhs0C8vlP7xOPxRL+e78jpE3fqEIesFuYNw0
DbK85fHwJVzXmWPUVQGervgW99pdsdVdOqgWvL02BQEOkhyChS9mbq5y192o/vPF77zGIMs7j7Cz
gyKLAiVKvwcZwXMSOxDeanZIB7sdp27dmXYwE2XUPZKtt9IKecfV4RRuN/N7juiJp0vtnAwajYt/
/gWEd7YdZiGKRckcXkF28TqqYb7gSnY8eCc4W54TjmeHKgJsKxvvOMCE8nzx/vVkSZi8UjSEXDG5
34eCSkxivSO/ynDZYqk63e92oORoCagZfqXdGKzsjqBSWQ50hkcG4ZA2DO3NRhWv5VEf2RsCwP/F
gmf0H1W9eLv5SQms47qPNGNe6fyptpMG5bLOoJHN8mUz6Bw60lvIu0YUWl/6dmETkzZnnfA9LC0E
RVcskWY6A5OF34jAFb8y5rmIA3pHr51y3Ui9VwnPWkqq2S4Fa1QbntotX2yxb+kAczvS/RjkG0AR
TOQkZ0+w58KLWNuTyOqH9CFU083v/u0DRobyUEktbdqGDS1JjLJ8+EmSPqtG322ygngWf1CZtB3H
Hb6qw6ROyO8JG8f6S37YIM5FG05MmRvmJhdK+t09vMZAzZGITiBtmD7A6iwwYI3tJni9EuGSSald
WcjEOzpgD0MbSC74ahqXADlkYGNj1mcF63WUC+g1QHqdBBIrlCnvVIRdRjtHqRQUzarEPS9mjWRk
6j5FFb14HgRGp3upTl/z69Gd+xhYfctzgnmGe+VqFbjZwieBYooIc1qN4VB/mtHeGRzXEgqxr9Wv
ftJipOgsSJEuYM+/TClq+emTq1K8sYuwIVCRTUJd5pgoTtodI2aD1wCeiv4YGYyBfyM98MS2u18r
qf0Ai+w5WSHzZIVosR9nqRCRsscdCz1SfpeJe+e5S/AC6cs32u+1z5Ot/WAgs9hoXiSsl3L1rfha
PLkXXUSqGtL8n2JotbsBkRycX3bvyATPaDYu+vNrONol7VekTxjQXMD9zxqF7L4mGQ8xB1JqdlQv
8PM95tsqdsbQ0d7C/TG8CyzYqS6NzSlR/M0zgqvZz5wAEDGOOHG7vLHo0iyvwfElJ27dAtcJpUj+
Urq241RYkgxU8ztoEXHcMlwoj6OgAyIYL8vycs3uoXcfEqvY01KgIoiQ2EuKJxPgARYTX1XHVb2b
38w4IdyggdvSCUYuIxurfRgYZmJIz+A7Q7FitVRxYwTbQCqyPT/00gJnj+cXjB7DRamwNeMgK9HW
PjUxVDbmX0fYzmfEPYA6nWv2pMsidx67jg3ES97cVV4kAy8cYSkmQcczGtqY0HkQYqq/bEsfqG0m
HkM24k7c3DzvWj+sEs2Dsg67uNHY3a5//sWf7ppZ5SQAwiyfyDicPePvricNran7hrjO8evU6FOH
zRD+T4bjxKIgaxVDuxJn6MJu+hTec9j4gwg6e0Nd5qjCPng+hdNIrYHPej3iHaWzcWCdLpDORDVW
NIyMiY9WGJf4ku3EULoU1PkRT6TdyOAwsoR8dhyRALEl/TMNBnwt4YzkAAhvUhZnzZrQs/EoIFuK
DlAv0krEonHKc3r+cRKmC2+MvC5yLMH8IN+rct+hXSyQhPOFfPoAY2laQd8QuHfkh3dJxPqbnlNQ
sjCO85On+DRGdrOOWdHgxV8e92jWL1ZpSzfZHKNORo2YNuaxZjIbKFnM3CJuu/wQCa6O85O4AGdD
8pC5W7XWy2slPi2usI8C+yq0CylzrYIj5usQoa4pPFfLmVYkmqSLKO7bdXFUnEwe9NKqszHqspql
vQekzxmq6M8WqkzWBZlhZdXK4fzQqa2wikGBYZYnlMxdc/PeJSqdhqcIf/TI3JHE0RXbOJdqnRAH
u8E3HYIJzV0+ch7yX/HC6MTCwCSKQSjKvr+hyTxcarAeODTr0ipdJ5bt62tdrovMmUS6FkkM9YJh
qa5eDftKbOPfX4xZdJBXb/Xm4hObXiOh58EqBrFMbh5E2D3LrVmTEIxOAKaEgUPzzWLo7Gukhzkk
2SbYgumgD9APotTLx+M+H5AEimY8XQwTgp282c3KACuWwEYCc5ILKhNtMGAO/pz/6rk5EbsXo8xM
BsLYsAO2ITpDv9TE6lb/ULGAZVQ6MD7UdUXSi1M71VNWoNx4LQA+1Cegej+ELTWuu9xz2RPAkb/5
UXpVTSDlheQU83TTiucbf0lSbHpdLDnvWzOS7tqEwbJDtlgHTsT0OB+LUxdQKNtwdNocUFq2ncK/
qmyFq9LHx2VTW7MaPww1rMTWaaGcLGhthBlVBVl21OPX2Vypwph1JVrzMh3TdR05PuXQjUlsDbZh
hG2zUuWlLI/sEFSUUsPElkV6ziutAl4q4q+uJYQs379NMLILsWap0aHCaELnVeEE10eWpmOnyOBE
LYwzw0nVA3Jm93sS6XbVaPrxlTkZ1m7rHAtLdQZ5icD7CY1l5q6D+GMoWJKkWzZHFy4pknSYhCjw
f/lWT1UtU5s6AR4Gmz9oSgFR8xH/YQYFU08Oqhpo6mkYtZErZRxg2p4/CfjoJLaxtyXnU86rEK5t
HQb/aIcl/TumYZqDKWAmrEvlCkjICzdLvyhMWg8ICPrZVNIOIlhDJ9+t/14yRIzxmBTJz+PlmLjd
V3fEilxu3b19XNat6Nr5c2g7DTPhyf5JBWmKKmdppyqvMCQtP/KTa+2ak642ijfQNcNe976RAzCW
q4W1wKQT04AW5MMO3N/yEuUArz7lQpMkt6oqx2Ta9mkG22ef+i24SVHDLfBb+aapF0hHiLi7KWC1
ef1hyc/I7L/JWHT1WrsLf6dr8jDmES1mpf9+LbPSkeVGOHb/+DqA0yckQDPIy1sa8ABsbnx2/WQN
jO1A0FDfw5d0iRpRI+udpP6zNhhHWeb+RW0jSmyWraeUAPzMPyUasf/EWcWw/WZVHdKps6ev7u2w
/u8AypJp3GSXPulQefiF7fLnrR5GhbiPRTR5eDad+0Lukr79caSXuQCwTirSS9ylv5L4FTj5Zam+
JwIJSP3dzsMk9KA+GVmuJSN3cr6Y9Y7cCWg1h4MGokbfm+5CV0sPcXEEFSh0mZ5Tf39gyJeD5jWY
Dm9KneIlwuzrXU+Ox3XttYJ7InT1ENSRciRKPAk8Vb9zN1fP9YpwWFgjuFzFLZfJj9c0AK+DtOP3
UAnUB+GUqNjv702/APmOoXJ4dbVhxh6rQB2MrEA+DDTxbOUAxmAqq3CS88YdTavF/28vCiqHQmDq
2QomqOwIIGJXAGXVpdVCvdaF1MKNYRgNZ1PhPtwDZAUPh7tNGlzDEe6O3P4o3fNeOy7AcNbSjV7z
dIiLJX+REbJviPFAkVO441Mk7cAm/CqB2fcGqkmzrgGRzofowYJIv6B6lUFV2a8poFDXiYrirj8M
dSIlWfgqPW4o9L2zM1i07u/ocGuOSuNOsu6Vt2Dyr17SGs4DK0MDlKni2S8Z58VxooaZPX2YuEvr
XvRIXF7mQa0KtarClO9vbptw3herwfmoHkx2WW5x5rHvlYScyAI8eNRJCPN5K9MyNAe0Yk2DHUqs
57nzjDvn7HwSky/XV0LLsfWjOVBvXY4iG41+6s4pUp9eblwOwagkVb0ZLuOJN184QWBa0Bbn6w9n
3s49CEGFZA/LdGqj+gYBaYmffvcyWEfPYihrqD22+SeRRcMvTz+Gy2GdhPtAXpDT6SV0X85YZeS3
e277I92Agyy5YSQnXIt7rLUdWruTM2IVkmDJKAhCJjzBovwJ6MXIeQPc/sGOufsx+VjtmC0GY1DH
L1R6PWX9VmJI5vofMkAacH3+B0k21vPWoMeTGGzl2Tn+mM0mBfwIItvtjTWMikO2PfN97j8NDaxd
l/XcE1k3rcc7g0uMfGuR1CVPfImmDqiPbE7DDx4yOsMlqqGO+bO+VcMstTf7LZHisElmv/XZke8b
Ec/o6Ip+Hn/NTUnK1ksqjP/44s0Rut4B6qD/2q4/42fcq1LAMXTqzPGJNJ//w/v1N0P2d5gCUCbd
OWS+hfmHhzijhNohRsSuiRN1RCMBboZXNc/YB6o5uT7LOoNWDlHVN0ZiuWEksBc/8gwluuVyEmjM
yzTvr8NgWdRwlApSjMKLBBuK9NvRoB0LZtc7Os/ZpnSvMtwDPmcmOriMRoZ3pCdOZ8/iaSnz75jZ
0coeUA6No4kHcxg6Jxeh6Hl7PUTyoeOxKJxoV1XZp3wQXv+q70ODgty88tU14jBw9hXN629bAzn2
TQpCS5/3WUtqr6s/NeF3gJ2TdDE+Ax+kvGZGaiyS6GVMwu790c6Ul08JPcyY7aoQZGwg/iZJ4JId
QclFtNTxW6F1pbnK5CsUPt6+l0zTRM2YDHXxSCuPWt38S2W9gdbK+waP7MhCc4EtMgoBWm2iOlBT
VzerFMHlTf8FyBpGCtNQB1DAngpNuHV4vHqsch4AR5NvxJHUhOnxObWZZZ0EUsc1g3MjLqv+0N0u
s7UID7TsQmVkr1Ir0hCXVXoSMfepQvXWvU4V4ejQNuJbSic92A0wij10gY1bhVAS/4SGjiVUFxsR
oCvV2Qro+DNbNMAUChZB1orQdH7amh9eXHOpcJQXD4l8GaNQCJDNpK2eHzjk7zSmfSBjV9LsGiqJ
r/03PZu4O3h44ugywQGvy4Y2I01n/wJJo4Tl2/Sahf/YG2R003XXeiSr/8kVX7Jo5tf0D4qYIp/U
hyRAfyPeSrvFtQ3gE//VPSleIwRnqzDdTuo4Gux8UZWEvnrIcdMkh36ZsE3jVpQg3UBGSs1+v2pB
rs6NEsm4jTO+xwxCgUlMpc7b6EtqrcE+tR2LyEBy2+zu4An0w0vRjTROFNEN4mwS9Hit7huujIgW
WM+x4TEUD+UdtNbeMDSVEeH6ACwGCNfzVLK0j0GB8dtNdQXlsBvQmP8fcTkjSu6l2A9mb7OxOYAv
I/bF26R2skSKpd8j1r1R2TA5MutQjvgLa9Mf1kivUuu44DwSDEU0OIjtmWvd+Mql7n82FFRalD8S
mbSRN4WdYXmRUvVsW1mSoCN33x1jG/2Cf9NUOEdZbOq373hF2eC9efho6a4BpfAB827z/sXyoXuR
ZiPhwoHtjiNK+Hys1y+h5iflxl3YGMeFBDUsb79TeiTnM1dfzovBHmM6EJCqvXysn33E+SLt++30
appU8teeMg3yROxEYPaafKNoHzYSSyZ9zHi6qhjtqEt9u/YKGg7w3FSN+0c7qiT0NJVnr7bX0XEJ
1FbFBlpE1nT0BhZpmMwoJkZQhqlrZILsRmzoZjtTLnhfwMPnTgWIuzeP83JcwF/ZbX24rEl3BWkP
As90p811Nz5GXucDgvnxuUnd3Qdr0tw1AjOqpSw8/5NE/MY9ED8CdhOC+LcC79Hq0rVgjZenB6+C
mu6RQRv21EowHn0WJ/JVPg8IE5kBlhJESCtAAmr2z39sgEaOAAdPNvyzDySc+iQTi9s9F/4g9Fxt
OowW34DfreD9EIswygd3jjHzhSqTS+dl1o9RkP3DnliFmB7HG0OD7RVI61oeGc9YvCyrbWEN9uaB
WMbBWKyOZSarRdbx82sKU38NJsORh5Lg4bTay2jPvKtHxGpi2YvewHmJ2Dv3B/uTzShbAeDmnSsN
EOQEZqH25eRrMU3WnldQ2+jXuQOtiWPRisiNm7GPrTnRE7mPrpBqWqzpXMTE8A4GpvFyyh7/Q+Ln
dm9fCXXDdpE8/2mIJbEDP7SNRU0AW/IVzpfGClt/h0XTup20OyBQ36mkyJV7bwlTCMTdRWNynXWa
ar349TZayKAxJt2dO7YfnCY2lZ0ct7Z4lUuBiwO6c9NzNKD6S0v0W9y28Wv67XPoi0Tawc1ye6f/
mI+sSA5nHjFl1Wb1iHuQ9J/0y9fyD/nOoCCRpHEE5KuUPrhPNC+6ub44b6ph4szGN9+Ck/5DBOnX
fWN1pYFY+2WTB6EKRjTxyHyQ+RgmDm6T6rgCPloQbaPERZYlzcR8eG4Yjxjr8HJD2ovDR7TCIqQr
578650RLCQBPWL2ryjenp3PvdfRgKQvWCLxQi+5H80JnoH7bYe/WEFeV4jVoa3d0LXOzCbCjLzIY
+/MazuZ/DvnCF8/UwHzWrOX4gk3VbUjWyInA0O0PnO9LwDS0k5ysc3v/lgqOxzingxAwPSt1j/4+
0wYgForUMqHGYGvGvPWKHtuVoETPSrxbvX/Cp7q+SlWOTXpmon/lZ8G1hs89TFZUN1/XVgOab5aH
FbvZ61Va7sfuBaIW9pBHzp6G8eyAM3xWm9yo6GUBtclE41sHMHqhQz89EI6GkMRq3JSh56XD/5xe
rW8ZKahov8/IWy89UoiYniAKIz6QTijYDclRKPr0G0JsVg8vnOqcZRErfxgBIEIs1hK7sXBquupP
u7g11LEcsHrkI99LJNWfQJo4/ta2bOWSPsg+TIS7V58iRs317OGDS4jpl3Hr4iZuRHlAtsuheDza
3Lgn2WUKGFHy/hbiRf2ioejaIzemMq6DUITN+uM7AdEUaB1og9ks4Be+1QtMK2TauTyBDfqaKbDy
pU6bD/MBUNmnMlLnoowmcb/xAnWzc+29dR/brrQ6lUBsBfZRjKLaKZUUtP+GFlyNFpBPWMFB+jPJ
KD9FY8q3Lfq0WMjOB4Lz7pkmzLcIJiCn304IeVCLQsTSN2VY7iZcDcdI9KBjASerDsDD5B5I4p4i
QxyLCbGpLjKs1rtOMPGkPmg94nJ1cBHg5svwmwa4rEGe2AZhtccJ75wdh7S7dsd0Ms1FHIIjZEHS
0Hikf9Wiz1Hd0ZoWDX6xmlWYTo/YW5tLDNJDli1nZGum0lj0ugbEqI5FQCIOsuE8a3MfK5Qb5HNJ
NTkR+X1YegiLjYJ+orKqdLCItdC94o7OADUEg4YtmRdsmOzbYQViJ9JRn+/PeJc1sc8FAhM3dpH+
ibADQZ+iEU3gXVk0RyvnJH1VMZxbybXx1KTa7ROnBYObwMX233mi42KEcoT6vK3RCdEeQyGOnYbU
w2Eoz86dxeaEE6FkexEz9IfZae7c21prX8Ig52SuSvlMyRcpXwwU/sQET43BNl5bLEKq7QfDFgX5
xLiXKFSuFue1h2n++f8mAjHFBHn3uMXqTktw+wxshFDhClTSRrKkY689gOAMbqNyQCpEpVkuvgVo
wGSGdeCS7yc3ftPoolfXYtJ81z5jbUzG/c8083WDlFB7d00/G7OU+spEkH+G7g7wXPlJmKhJX9QK
eNRYA8GRdmlZ4/WWNbnreno6T+l9vv8vzABTQsaMcXI8UJ3bDKTwduar8ug8GhB9ldQk0QjEOQlf
Jr8+kffgDZFDiU2CRoxUWbQs6ybqR382BbiRisZM80tb95qYuyugXx1KoHfwrGncLeGl9ne6J98Z
9nErLUJMQlty9fuCfdaod+AiO0XX03EAqanbb104DIPWN7c+dgeP+xpFInFZiRJFt6Eo4EeQrC68
UrujAwmUJGuy6uu2NEq2DgGlTOrs1R5lZEPWgxqtdRYPtYTFJT/1G4slyGRRgdBmFnouE5S0a964
thM/3F/JR8WeyIRf1bTHZbkK4rhp2BG0OEDh2SjXSCQ9cXrmNtLVHHvwOoBuCMWi3vfoMXy2UOdE
9vPTAVxd4/FyNpke0+prnoSazHGxz8k0WeFUttQHJPCJXszOQgFRW+DOn/IFlh3RyjikLsgcV3ky
cIUnpSsdkOfU+LOgejtfy5YSYnumnqGLUjTlKnO7NgiqzX0h8mVIZ8xVNKSlxftqE9zPQBKtC9An
hcR3hfyLHO79IetlLJob1gBhY5QH8cclp6uKzKIl8TbbabQre2KFVPVfZmt5L+39K2lVXKWJ+824
5zobgWJYAVA1JMX+fFiKmzsbim+XHtzY59IdCu0cMM5R84hglgMjyrefTlw7TIvoL3l2b1Z66+Gn
SlfERjZcQddAJ3DMTKfA2+QlxmD/uvACSkGYYlw70xEOJ1+QcvhespEqRJ34CfPZLY5pLrwI3wPh
qudl5DDuZHehMKDNJoZnm5CZ+y+3SFMuY+l/bgpb5vhO7pkUohT0RdQcr8zO326CpaZsmHfVY0R6
iQyH43vat+FUrOe1oSDEWM50KH4A0o52AT8I20SDBvGGb9GgYOMuJkGRYpca0F7NsAZkA5MAzGVH
FR30otCLSn6p5yN1e3m65wkwNQXB60GNYXw4z2S5Bls2eBmWjPSVgv81ZMx0P9ySnk8FICbhUnyJ
TSL/MZfNsGwdtKj5TDXEWLDbZWiqsIGpqzGAffFHE2PFIFHdabQeAlOy7UAZ3hpqYXrUk6T8+ue8
Tx3zhs9+M7hhirTCFjwuj2MunXU1YZ3CD/jKirU2cbxiX6A04V+Un+hnR/cnFYd6y1ZQpbKnPtJF
kKPS6m/pfLBWz25Vb6CY4bGHORkmYUwit8NPgZSIDXY/KHYPrZUVaeV+lhtAJwrZRD3RmLVR9Rxo
ThfRIvsKxEjrnF8DdBDTdjXFyCGR5VFOZw+RRL1DpQJepw6FUYcltX7YGqk00pUiHTszLOLLhCxR
2gxJWRhV7UR8Np190oQBFyXaB06DuWXnNyQvmqcd/awe5ynQcxmeFBDKsM9qdJLhCns23K1hK0x3
TQWHgwoH3iwFGMKJKa7/MqSdUUkF+yZTfN/1KoAQKtg6/I0dwF6nUmoyPMcIpwKLjhbXYLFJfzwT
4Ph1YumRNbmc2RtvCWJxy/UkJQ+6480PM/m2pHVs360pHd86sFeXPccl+9PErLQgie/iffvCeLGn
ktJaWOtkldvoWQPjQb/NN4jhjvPzBHtsM6RJp5CauYN9RNbdq9u6qUEMytGfVQOCv2j+d8Lj9Lm5
SDw+J67hlIVUT3dailqzLbNo4MLJlFhPp0igaboH5AJzQwSD87NELcE+WD5neUz+KVKl2kjE6rVo
qa6Dxi4uA88Vwm9l7McoKI2aJTs9+02Wk3hKglkz6+qxNyPFyOowq4Xqs938gEzAUkoBlPI/lELr
WPQMPL+6hDS2efRr8Rmv2ggdlqJ4kuz9MELoFKrTXA+pRFcyTu+SxEoOCj+n7U6VK5egZlLc+iqX
wyJMKOB5idDtS+IrCpBYOMaIs8cjgTBvKGe4zV7GjY0ShT94AFkZLAjV7+QmC1YuMEvfcr0QN7RK
ULFDmX8aIQ0vEDkieofjUM3J6WfkhkJ1Y1jKgUlMQlYvVreU2J+7IsMYYybjG3k2HtyJq8RlmbGk
MEkGo0H3W9PGLEXFlrHzWbgE4MhQLI+W3gNv5L/0em48R6QdEkcNGoQYq3hnbccciQZm9Mhw6iTa
Dk+RojdT3TDa9I9js8dY90CoUgo8WhDg9bkNiMsu/oWoGDmdJsE7rl7p+aA7cB+cJB5OOm4itxBr
KRdFclhssH34nc48FcJH0MG9FlPwWga5pLeiT3lSG1bdfDrscpEsXYTNqcLgSzN3bMFkPgkfHFYM
gL3e3TYlOeKAeCAT7XzPWl/41a/aDu6yqfihWAtR3C42z/WywZGXhqT/Gxxgn/1aoOII6F0RD32b
yQDf1aeK/LMaiCf6+hqCu8MMbIZVqrW6Pq/nTaUf65S8pUyWWBC6jJb9JFrozBK/ScMY0mmO5/Bv
eS4GUS8T5YLLwcJNTUdfXrhv02RJa1fAj9D9zjNWnj82Kn06Gr6POW1gevyRQV5xd9qKiv+TH4tp
QI6MLlsux2dkQBqh6ro199cL2f/q4GbTLDFVl470i3eeHOd+PEv4FTs5yTUzVsqSKx7x6e0fSn+P
yIk4PN8YH/LWbUxMqSgRYDK+sRx18nX8//AZ6aJ0Nr1WNVIDUdnirDVakBTBM4P1VGun8tyNbwQ/
hQj7bsUG8HMdrYS3timTR28WOX4OzuO6Rs09EnwlBRVECvWKgE0+NHm9pJcRfsHB/LMagJe+Wk18
PNixSHBaZhJ/B/xrEgxFunNlxfcJ7SPskWv4JkNwUK72PmKJnY0KJ2EBXKwkzxu00kyhE6B1DEyy
xj0vAQGQwM48AMfO9o0TdDzWgWdKXiOyvPiSQyHeQBEVJVh0+6Dqf9Aoz3UskQ1iMQ0e6udIsUrg
/YdoMc/NB7baq4YLFfVXThXOtVatyAIVoyUsT2CXo//fVQbbpUVqha3tPKvbDDsDujczy1ONB0pI
TNVkZbX9nchbSPyQmR/vZAPgxadRF4qHpH5tUqULHUqK1xWbGeeI6IuqjEBIJCL1PpRgXhaFUO8j
jiv1Lev0Xe2DCkwuj0BA8ah44Cj6x4eCT9dfMJv4weDs+n2nrUb9Ef9z2Ow+X8Z4V3jTG7iHaxz/
OMATld+ESv9rg25WSmEut7J83CEVNMcHjDe93wGfnPLej9pmQ+kV2Q1Yi3FmVONYJNeJAQUiUMtW
oLNjLwKO+H0BJKlPe069rM8xHauq6FZWgPwrv5HspO4Z5Hz+3AE5d4ghcfNFUGyAnOdPgJdlaQ8g
JKsmG3Cmp5IcYgtZIREQ0brqejn9tZrBNuSW7uGiUHXIVIaoBUyLbVl9vb8/B+glsPOOq6eGMTKc
zN0/fFGJY9NgzNTOYTWCHJBxCYVPNcKWp8TuRORQEE/XTt9uhW90aPRwvn6rbIQNq35whdDQYKma
2vyryqCb1AziQyB+NS4GhFRA5Yv7Ye48wzRQvs/gvqr87qdlbTZdXF5y7AKwKB4Ty4VHdTzZ4tK0
mXoEGaeLt2bjh+hMfO10rSUNXTC7XJ16prsHzWopkS1jSWPJ5VCilYK2Yx9WHIvSEyHzZJcrD4pW
kHoq+jj0312WTj8eYiw6RQgwzvq1GSBa7T65kukRvTBC+/Z8xMNSwSw0CtAtCPTecTgHAEvGXZFn
8O9pJglzRotP+iIhCk2YtGnqFYQyeRiHxgAU/2ExpMfJPVWTsNx8Wwmejhayi+OGnwSSjlDwliRj
EkbMETqyPKJrhfka+QwO2PdX4VfousdGmM1XhSHVAgzb/MLoQv+s2kecL3y3IuHDKg5EEJOvVDC3
mUgdvaNAn4R8Q/DvHpoxqfHbLZ72ZqhPGQmybdjPKJIQO5Mcsv/y0ui9lY8jnJKs2RttBozqsZ2E
XBJFU2BrYs7wQHicnUHny6WzSQSp/N61Z2LCQEtx9q/co0g2HB5XmoOH90F5q28B9HmQao7/wqhQ
JFzeQ/PmD3o9EEU8lswWmEimo3UGagWgxZcuV+8v/ipcMIxoNE7kJrfC8nclOLUpKoAXdkr/ud2G
XKoiHt/Z4aIYLoItEdd7pwaTd5UVR/nvdpRXM8N9cxhOHVpWam1BNml62HB8PqR05IwwpzLsa3dx
6Ku0n7OJG1ktnNQx5uZ9iw4PQxZk+YeD9KOUE3rJOP9mVXTRhU7tPB7BJv/GEhlLPmVhuZ72PId1
nVtZ904Ld63/As5OfcSFV0w45Jgzd6KyToP3+7qTO+rHuXWagQzUWS3L21J/pDVL6i/QqvfJSE06
2Y+EOL+U5P64oWNDg0a+V6Si2Q7pO85pzAglWNU+am5Ow7hq2hsA23eP06QBbZvTEya8m2APgdEL
Bearicz8jRHTJ2gUcLmMwo6ZaJX+2GeIOo9AzjP/H6MCV2HIsTz2VaUqWi5ti01DmhFi1I7obfFh
YUXrQIaCPSi3VlenDn8Q2RrbbHvf3Dy2EoeTO3g18SPeQb956dDCATphSCqWM7R7RyP4ZF3UCcnX
3UJXGF/aqkdPMlRD/e+EQY5hGmDL/tvM/a+fNlwz7CW7IBaApf/vHdmsLC0OpPReBo6PFrQE7aK0
DxIll0YAOIyJIR+2j9mep8cHwJ+YSiri+Xo1tq4Jpjx54NgrqxwVf3t7JyTIdHNsCQejdXBfhW2e
dnOIw6dU0s4VJYrulUwROo8cjLAnenAxNwAZ18cu1SMDsqcUzpdp1f6ono2rZcUUML5vqQbNfaWx
rV4c+Zoznk9Cu2OPH/lX5MfF5FIic/FBXRTc+yYC/aYqRUf7ixBVtmb0YIdQvq6H/3PrwDQaOiJR
3jwxUON6Lwh+NTMgwgh+kfqEjP2Q4iRbs1dzLNYw0CbWXRSUaI+xJ5iVb/XPXVS2/96wKLp6hSdS
/gfyBaYQ1XU2aLoQJ9N/nxvNJNOgNN32hE56432+Ewh8QX1OXrAcVRuRNmBUPAZKnDGWyJ1ddOea
X+sP5EFSrrpnTyfAurdU0T+FKkLCPj1hLt/u3rWhLtFSiknYCC1eeFi3GIgpATo8+fCgHKqKEhYP
3Ykwgcjp4mvfm0Lj19Z1SFQW629FRTipu4MkcD0aqSOFoIr8wtp1mEzD9NvutpsH31W+qSC/wLSv
57BxI3QNuIQo+WAsxRomLBqApgM0Mrt4eW8b/s3qtfHitquVL4+AWpWLvhw8+AbQDLVLW3k6wy3h
d0v0e39lV1xZAkcgeRHc17QCf0gIqoqC0CTgOqNOfGTZ9JTsTa6FL2YSm2yts8lY+SeFGfLyOpVw
0ck6PsLbicWJX0E97XsfMnSvExA8HO43gklpHW/RIt/UWJrLsJpcUIR8Zx/rOqWb00RaupZPYacD
NgiAO8HZJ7jrs7qf8E4pqzbWRD2WbAH33fMOum8yjDI77xXpUsn6FQ8iMvzw5O5L+0oJW+mH56lW
5PYzgqo2ipj1LLcgUJj+q0Oc70y4ng8U++1Gkf9xvpdUdf2nnvlilYhhGWIITgPicD4YBYyYYOaI
6k7untrRqADXj9zYt/FAV9n6dsSE425jfQs8M2anEFMpJlaWK4OHjNtWXL4a8JudQUujtSbOevtK
h8fNH1bz1H0HTlrCVj/pXMetEZTY45/Avwqa7pDTm38y2dNW6m3jloCL0oyQCJEVSV00u5uRNKGB
UXI+WN+sFtbdlVr3x8BOnPQz+vWtBFGUO/KB5G90RDgvmIw8oSC5p0rcIrGwsrPe47vilyPBnGkJ
dVbKcMpmjYw0gdNu7hy8duPKkwDTuvpySMjso0Vcb0zF7j6glgSei2zE5M9i9AkVdse/XULNnWCs
y7T0d2dMBgv+6jFzFxIS5TIbLHeF1hJxXi1xFoL7nWViAAEq0nbP0kleAnbsKLIjrbFtpju+2792
+QL6wkHM/Pm+XqKx22jREVWXRZ7uEWucBKGNbhqp/mxPE/BEzCF3Ic3SfF0MA+S3hPjpdOhmS0xK
4YxMaNg+SV+71zLcxhADU2CP0H0XFb39U3UXg5ec+5YpFUZTGYLLP0YfY9ka1x8qesWdSlS8DQba
8X+cAaeKPQccwdLmhJItXrzmDKQKSLf3eV2gvkEQkmTBFXW0heXIZ6uOpfNOfYsHxie9Ykvoguu/
nXK8I3eokdSKvNzHEd2stydJfIyX1D40EYip+lUAkiz0mCW0qFPA5BcLwL+swafmNkAnwjHFWXkG
x7HZehrYPVRmmg64jkOrOUUYE/7AglujQ4NBR7KXx7p0IkuIc6bhkQbHPOC23DJYTjrCmDWyny4H
jz3QWKfDoo7EZnFWIxfgz6nv0Zo1bjr0EdKMe20AqgBvjZFTQ7zUCWYPHFGndcBmqImrKzKx0WeQ
gW1tA8rr+yXJt0zlD7X60h+0cNIcmeqU4TLmL5tmfN2iVOvxzqYHAo2RXkC6G4Nbb7kTX3QYwesI
zN0/sELNgbVmhG+oBXxM2zuOUQfd0jNQ0gEbeOmoMfNPaDZ2D8I/43nDlGofN+xV7Vxj1HJwylSP
kKMA/JKSNDlJFj35YiMVIq2HOpR4oQ5Pi8ndtXiMhiZfoNXSjDp1xeaD88IqNIe7++hUJ6Q3GgwK
kmGfoZ8blMWDDzVUC6Hk+6RrpQzTTp2nT28qAOTGmhlwAiuPeGb+DIZKcpVRYRf9aubJXctenK2e
Srv674jXJDBjRyoz66TucqupiD5kczGlYonydQL5/0C5LDDWSpeOL9lkbBTtI/jPuPX+7zMD/k2+
y1vz+NHhYQSrHqvjhebKMPtmIXujkqmIZnNxHEV+eE1dibF90JSgYVUF/lnqtvuzTMeLdT7BWKgj
ofl5vpKXTyRMLZRJNYM6lh22z6GPk9d0IDFfvtgfuk9Gew8rINfEYBIGSyG4kC2dlqDX0akFkwCP
WYXH8OvgQNhnZiO6OCIT5rWJco2KgGMgM1BRV+MkyMMt6gG0loLV0F4kjp4vHqoeXNgezh9X6Vth
fpqi2Dqf4ZYRWDy2fpfWR4Zdsv5SLlVBV9laeXE+nQJWju7Yu+HXPtMESoh5ep63GVS9Zl7BwExP
Fz1MHZhXPWBjtAi4pmPLnd1WbHU3MEqEscn/SAX21eWx2VSy4eZRijY2eDtSWTAGnKWdJAtU16ID
q274aX4krFEPluxnv7qgJp13a2uB1Ci279tD5q74WKESOxXdwCXn+FZdLMyG9x66icSsP+dwmhQV
9GuQeh8RFLMwCiGqLyvUCgjuIoD5mF7poHOx7WRwaHdGjuPmDwydOwoDFpy2klwive1vnFeF3Z/v
zHcPui4dJeemdpzSDyG/mSIGjoLyHYoC675GxAjyKK7WXWxj++rW7RvHAPKsMm1do4uOZeSs+MAb
IIVtniM03+n3O/+VJpGKavlYv/s3dC0WJpUDwZRz/O588puKbuWq3gzST7o9O6+ENwMj1LmAcf4r
5YuBIPQDiPygtFHCG4YLusu3K41glUCVs6RQkHf468P2hg6fu3RXSBkdGjpLLNvZ3sVhYcZXszpp
4PEta5YeKcYguC8v9j6efqVFYAIkZ+Ez+nXWpTQWGHbV3Kjc7OUPds3qlcoaaphdwI5wvPbxKhBi
gDSs1EmHGSpskwqMXRMgPrpPYEa/iAq12iEUdau0m0o8jaH9kQXzpvVb+tKrWNDhpQeQ/f3WrtRn
OL2F3tYWgty+Z2F/LFxG0OfsAjPCZIoM9TFf1MES9zZ9st0oA/aOv3SxQZcMwOQNScKd1+m6R40T
X10Nk3KFrzLPfhd56b7kB/pSYzyTZSVASuCgOHZah4isEx+lnMDFQNL9ipSK7KQ0M5bhMVbMVvwO
H+NfbSRjqa67lGFHn61icPjuNmLYTz8kbDOedZdIjcVAkc8hO7hYp70FPbCg05MG1J2T0VsQS9kp
8/jN0Xti93kBEqpd6HgPwL32SYGkOKg2ifsgn2d4wRjUJ0+S7U9yY4IaI1dcJuVRxUXZsxcPmJ6z
Nv7Yra9FFdEoc98Quy34DXoeh12iS3ovjLJTaoKAM5jdfocvTxjbwERPfdKik+EqXSzRZpMffl81
ZXEDuuk5YDuVTrmUlpqA9ngjSpS1um1Qfpys5CI8yZ9Exp6/XLS4XeNZjPOJnWgLomggUcsViVnx
NiGDMXlwMlpmeKVm4aOeZB6BIlq8Jq7SRr1kKIRVDWJf0fDJCwJghxfwwcp9GFs41jAVlM2fh2Bn
VzDwTMZ5lxanEQ3T+l0DbjscRfTr6dBNHJgU1q2HnrL9d7n9TCwlXfbeZUNiWcd98KIK4yp8t1ra
43oWG0zlYyvnsIpnCPi75+eQEkDxglTWPq99fVrdBqEDJ1dSNNYtxjAfX1Hk3tiYpjENzbeJb6cY
pey68RzZqUO+J22/brYv7jPXESLmLDjLUp3BD3lGUaV0DfBnPeen0JG64D907DIihDZQKPcr5mH5
UyFFZtBj+UseW+6lQVMEiX5XDORvb5fQMtkd32nohIjndd0uFED4GGXuopscDKoqGq7al+Zmv70O
D+ukd6SNeKNcoLBPyZIwzsHtB28b/+8Pnb6t7vwPYzsWNhsVqvPz0P1FxoJ+Palqyyim/LfOtD/R
X+Ye5a7K6QGWfw9T5HwcF4RrCssccjWjuFMdE2p15yfR0tKNwPTGhNd8aH7XTlLQKk6euQ5xpVIp
I7l3ShfoT4XKPdXRDAsXENaRnl6qwkHHDp4cN+G/Y1MIO/iTdTsm+vLgJ8UHG5YQ5ughwjtlzlyO
wQz0bXrpg8ieDzJtQ8U3hErhdK3N3Zw6txnDZR9wzvX0jw4/KLYWkN2zd2ftfPNaQBqxZ/D8Jnge
CtF322aOBwKh2KEBLeNC0Iiw62YN7wIviCk+6t/EgMjz+ardBjif7m4S7J5PhU/RsNgu/x5FHCom
E5bamJ2t0e8Z7YUqj5Mi7ud+Kb6pSUJZ/bKihQJX559BhKtC+nMlL26t+a1FmY1PKftF1yKKq/E1
xwPgmXx3s7G3HP7K9WnaSfqXqQJT5tbu65bFZHwJ5k92SH7OrdmFbIjdvnT7T7P8pg8JN9NaNdFn
B4GNRMpv31rC0xiKCaPjsorOElDmfb8DAFe++8nRWGB3Rew1cMYJqbLsElcfm3zOGu5rc/ibE3lf
ioxDivsLL8xa83MUj3WYwnPpDOEZl/vo0p13Gz8r4qxKYUv0Z2dG6frDWmhi0BaqtW15bqXId2bU
1urxD2jLppE/YtfTWA2QQ5ub8tWhVLVRKxB2CFBJuSQtT9MdMkkc4kGXzoy7W7mhnc163f/o68mr
z1G4pQiuE04NJhMc+BaWHqG278fqw2i0cJEkTWmR0yA6md82hf0WY+BXlc0eLW5kaWih9KEsSxaZ
suCMlkN8obhO5H4nMbS1Qh7zXRkXmJuMD7zfhzIcf+JHaXwjjaSpN9eqNAKgV5DKi79/Gvj0dugt
acl22rE4JhmmuXNbLV8Km4Bxtb2AWxnOdN3uozZHRm5Dm9mNRHamB334lyviu3/XRxthCdnlz8HF
x0wWvqRlNTlFP18wEftHnUsrV+TbWIwXip14xEmouybI1jg+OS3W2IhVncA3D0b2SGWnSSQO1qfm
Ea9x1LHw2MA+ZEQQhR1PY+L52TCeLnAY/uTZEQlxzowLnBAX5+aHPfx53rxSLv+oTuHHBh9TJh1j
R0C0acGGT6aybApkiZC30r/oTRnGZZVAd4rulXAfPkUpJG/KDcsuNt/8VFhozr4MgcCvNQDFVAAA
L2gQ+l7w75+iLBy5sUdN7bsC9wNlGKTck7eHXaqO8TZUgW8Y3/99cDXnc3KsiH5PZ9SLEk+4XBoo
wbEnAzbguZTZM4F3U1dPgJMR7O+0tLNGTM7OMqFWtx94x+hEf2K8p7BBF+F9qY/V0isSnWUb+uok
pfDWuOvgetjW6Uv3V9aE1mqE2k2ghjjvE84t0KHwj9eSMkY9GfNozeL02rz3ylcXea7eCcoxwHaT
CyyBD0iN/bPVPeypGx037CPIDPKMb+dMNp27Oypxllw/vut0jjZZPmnpmS6Ve32c10YfaKOwRBha
vTsk+H4nQjk1qMkOJ5DA1sNCYd6Wc9PaBkVFjbhZxpqfX6vLTYi2Ouyy6wuawEQxrovackkDAAkr
C1+9Ow5135ICJCF7zYMygp+5cqKvN4NnipEDruAEkjTlHnbChAIw5AcaEwN5xl1CaO0AGRWYmPsq
5XEGuNuN8+7wBghWdOJJgvQwYAUh02b3GE3+PbME/L1R9hwcVjbsk/uzB7Ttc3Cj5aRAADvoDKX4
ju1QJYsl9mFKhFxZyXJXNrvy1UFEjve/+SJ3cRRiz2u8WZAVMRf7noEaZ/uWpeZW9yUf0f+rQ6YY
jt/a6VfMMxI+etmW7uS6vgA5oy1WP2/Wn8e2KGdqazzf539YtdnN1R122+Hxf+sM3vFrHnlhnGou
50IqRjvDw6HsYVnJQL4/QJseUQK8RKyMWeIwKlBXIkpALtom6y6XizVkT4ODVyrmpNHMbuy/Kjn8
Jpm5xRtvtWnW+HEigh8FNUXQ2NsoCf7jcpNQvGfUdDYcjIJuXO8qxltugGD+EMgQTb68aMFemThg
PDw7lsJBYfQDGjW5mfil05M5KjAn6FUAmtLYvXvF//8rkPdJOdw6kjyvYTjcee394vnN6COhAQdN
HxE6WZ8utNGHrYf0H1OhHX79F+mRlS/V+43wesnsgJeBjKY6/V+0sRTNug2oaVtnDUt2NNZ5ukm7
X7uwIbnpcUATQ+r/rB/6JYmVlhD1+kSJoSi73SalIHxh9lQ4nRZo0nblPZiL83CIokkbuq5XVZXs
RqeYrnwzpUreVtE6RSF5jXE5XPecK3Q4H9QfWQu1E2+A7b0m7sFFLHlIRUQ4Oagrw2pmLhHcuSJ7
A3Q7uNhaJgKIhw+h7tDSkScHkrC5f88J6pbFDHLmb4jnVP2XhaDrAOnCTWuXAMVhXDVOWefWuQ+k
b7w8PKf4DHS0l6R0y4RE5fE28s2OcoveBw0JGfQ69O/cc9ioT03likAAaU4/XGss9lWqqxa++TuQ
WrZ9RhQAYEwRneFT+Gv2x2OVk7bm0oIAuONlY5BQhDcE+IKFMXg02Dbxjyf97bjgw71t9E3MhoHq
sqsMJ0RzVD76kmBerb7GdwwsAbkldZSAYwpFejFwchBv9BbtFCGDuxH85S5IgQuheEuLWkWLhDi0
8tMdPODrz6FgeoRvrVQohOco9gne4ByfbqAyn+S49ucyaog4ED5ahDoVG3uBsoxWvnTJ9BjdorVN
dTTcVcGIBzLPk4vtvEMwLBvenro4KMQ/kzoZqpfVe3Lh0yrPr8GBFDeVb5z9RPcWbmSKqjcPeVno
w4YxxtcBmD3huqaFs2jMtZ8mgLs8aKRsg/HpZjLNG1IeW/kBKAemT+EaltJXyvqP3103iZ78r4zo
ROhUZWVlaTuMx1dSx3xNGG02V8FltKBrOGPCyhz72AaJadHIlHaT/Ni6HL6ebszE/1xuQXQQ1VCU
OhceWtY0UnjdpgXuJtXefuaBYXJHVdzu035cNVzqbI0XypnSO4Lg4PeGE1F6qqPHXdEU13WXTp9r
dDIaPJyHr/n+YufuXa65V4aCIY+0g2oQH4uHVCaNmPLPNO8uz6rhzyIaWh3i99Mh6IUWMQOfIpZF
6w4C4SezxNdfYzyJNHdTLSWBCHtor9+6J9Q7C0pN7KyKw9jBLtxaYMhbXLGRoDytXy8d06bjwwQ7
Un1Y4shv1SX2AXbSzxIZKsQwEsqaNqvY37eEdo5LWBpWTFnitgD4qr2AF82C6qlfmxv26l+5W0ea
bL0CkYPbPLNDVfngZUXUVgdxmVBN7y8npUrJCXlBOkLXowASG12TUHvVcwlxd6fTaFUnw3NbnMOS
7o8oUxbVayqbw4aFskfm9ldH47sgWIMkSe4B+1x0sKh2y3+3MH39VCCmV72Lm2p1+uC8oXoE+bFM
5JnL5289/Q1BupCtOMUi+uueiCNjlQL7KnhU1gpcYiLpzVTHxMD0EI/9fSgVSlrzO5p90AJ3hH5Z
w2EJWeh0DeGmOI3QXRmsIUmEry5B9RVDUCYltTR0PZbYnWBBrHVCoOkyNbH96I8fp0DTodMLboBO
Eghax/ugdUTxRUMji8KUK8ykaTz/CtCbEGDbpf/pXQCTmuoPxQlM8OCNcFIyacZ+RMNvg4s1baIR
Eq1M3dhLMBqRj5R7XB8p7zdQegHoenBlIUdgWGWIcPQsDKef2i00xc9ihVanfb3t3zDpGvKna/XY
wbqmf66PG3PWf/kfNJAjdVgvR8fA6s6FUmpkwdYfBGIHEfPIg0HQ9HSGr5w4AH28IJX0o3cfhWGx
SNPc/mzHhos3P0mlaCzwEx0lcqRORtKYV3FI39gMuqKk4Lf5l1/onJf2GUtDuZgHmjiR80TdCe+E
7bVX092GypRDJixAFUJup271ycnGPFCCynyVDk1UCl9DTiTXUyih2Mei25uvfTk5eODUs1h9VUt4
jp/ZCBAyPAgyIJtb5KC8+BWPUk90fdgjhm4tX+2yLbXcFSNHlzwEBxa3oM7IPytPzdmYzGg215mL
BS6V2CzCluJe3o5jWx9gUf2fHgmrfwS/Kq5WpfweCw7+2CqKD+hO+pw5ZM1kHmdUnYLHrejBnlip
+OxsQRYKTu9CTTAdRpAihlueArcTCjzATxag/z8H+pUUO85ZylBBK8ovzsARpLIyK11BaL7ty/Ai
/fk4HosLT/isFBZ7+ti9YnEuHK4kxdA5gVGGL++VW0lxHYgPSCnMc51kcm9eF5NRmCQZ56biLi3J
QT0RGKpLbVcJe34JBpeArgO8WW54s6bqy6DYKI7NSqUE7Ow84Kh/RaMwH+DZV/dalapP0r71W9qJ
rUiEyrI48Om7v5q4gH7AkCDSwiuP1ezXEASRXWFsaYgJFlqDuDzv7RSQudfGovkhAzi04pqkGsm2
toaPtwnaD20agCIk8QRK1Awh54JdfDY2GBXNVSMLxM5bilzHZ9kfh6PR3sVDJFsN06G2QIqSL26X
Q6ALqH7X9r5DDzIncccuavDOltajIDpmV9zL9biCXX5ECfQ8kpmsHctNXsGhreWyIy+rTxKuDMD/
vrLa20SIZtlCFZLtIdvgELOeeBAeGoYcwEULnKglcJ2WRRNUjlFB1apzHTH6CaHnJZ2S0xVKdGNs
NlHEhsHe22lMOTu0DtvffgK4RL/GqcNrRnLDujCLSFjLX8I7qsukFyK+C56yxHQZn8YQvmcUqUft
1LZHUi0Hq+WNHibe5h5ObT0JvMwvEfyp6gSmRTSmju3ub96rKKpcaOj4Etgw313eFS5oHasNTx7i
a9NCHr7MRf9v8BBKKHKOoj1X/ysQxXmAOmOhNq5zC7yDVhyKjgN5klSTvFXhhqu5hGrd/dcOdKJV
7qS9kv7913w+YuDyz4ia5pRsZAnB8k4h9zivUFJrtF30I2QMOEh/IZ77tTKSKaDaOH0vrnQcCxvq
mI0HqbtCA3IJR9Q6ev+pmPkHaeE4uEfHOn/pdVQFVCCB9zJSJPTbZ1XkcFZ0+KuahH2vq4gY3ykW
ClyRrBh5cxMVXCmJ5FH5m5A3F4vJTASi4FNBcAb9rSVrlGy2PRPsvhP7+7cKroLQNd9/2QTdvs5E
rhH4HbhBIo5/8cVH8Xw2FaixWnArjcCEIoFFTb0PMSY9FKiLCbUw89ntWIrTkAPXoZo73wiy1S4I
ejODVmOi5Xsrqm7gx9zr1oqERdfkZe34z2v23WlcaWVH8h1/2fY8asb3acV91cyabbFlAFfQWibb
o5Qz3P2VlyJj+quZiozjMFcF91kYcUBBx2ACOiV0HTGa7qx48LcvoUY/ifYV12AtT2OiLb1LZsCk
gJyl5NP8GUErSVIVSMHRbLVFdqIJ4n+1vy8ScA1QQSjAMZAuXPqoCvZ56EsXvBQX0Pw8H6UlWRVf
m26UqQbaaVh7bDY/3c7z1r95LEca7vlt1zDuqpzhtwY49+72R1n+hFdUDJu/s2xQuaDP5WngnNhE
N3NB2TEfqcAbjqdhvAOjMUNyLQX2LotnT/Pflg3/gHAwEL3oBVwux2sZ5bQFRmvBg78joNvmvCQ7
0mBywy4150sVq1D7Gnm5zqT1XeIH+Dm6iwObObILdfs+Rtjgd/g+2ZvN/nDT+ghJPeuGLBUb4XsD
H04PU1J5eUp65cX8zWAA+cEDOBYqEVGorbpMnqrsBF5ZPg9MHGNTmrBE7PhavW7B5J6o//TFsrT6
sGTi+KXAB4eWYY6v5dBuhxK2znpD6Kt2ZAXklHWn64rIlL6Zwv5irD6Ja8Q3ADu25PJPcoJbAx1p
+Jv7DPZFtC8ig75vu7VbCIcngZ6OGK9iJEJuh0kiwRovPxJaroM9upLvTGp4J+VYe44m1DcgUJHH
FZOE2QlxwhlLYeRgmHMc5JjcmuSAhhWJ2Aa0TY2h/2NdL2F4Uf5o2It/0gJ13QUSpDwBzxEi/zOn
JziWk+45HsWBdHdM3HkvC4nKbUTIWrE6w54cDkqxzv3hzSqi6m78Pl3LLb7oQZ3Hng5phgDE4k4P
EK+BSX8hx61vS0LOyNuSwm8PRotRaoUTckU8aLwvQRe/9oXZhte3HiLP43f8PPvTfdUBYC+Mpet0
iut421s+369t549lI8aGhfUnOSQL5Q+CsCLKs67dr7w2t+yav3Y9/f1E6XSpW5K5kQrwOaQKhKaF
DxJDee8mwgxV2SeNmiqpvcWsygDCCV0CUeML13JOvHRwYMYCy7cjf5sqTpjDmKaDa9snPWSiZuzu
Y7oQLE6u1OIxulPMfl/kR1daL54whXCRjBX7tVxU0yKopqcKKnizCa/vfJRMEMT+vCcB4qKwfSlc
k4ppsN9jRHiia64QebbxcdZM8SvRHzQdOsqY5tbQkxIWYUypDzVaVdnRGz0iVSxKsIw1+uXiGjON
ag66Lat+fRHIxj0PxJI1kHxZJPjSWWKQQ5d6Vvekv4qrYYrzY0M2RQxU6pLSgxB60hM0liR52P1G
IUiXKwBghq2J+vUBdv63V8zq/QUv06ErzvuqR71NJOQ/FaVyy4S69DyG41/6bVZoTJ4zwQKwMgpN
mD0p5tXQwOA4Ru1S0A9MtVa/RjDQZXuaCLAqDl5KDUTdlz4WSzlukDsts98HX5svkMnOJa3z72p0
gg0577oHr672jNk9sOPLMFWFX3qG92Sgkj/iFQaF4SiYkQ1LYmPIAKr1V6/h9j++rW4IE4h3p4oz
Jd/k9F56hXLiqGwkgZL3ZsJPCvamQGLhui7G3sW22BJ62hCkHnqlzjEahKQblG6jupxMDoLFSG/+
8uG6nFN8JRNOhAr6u9Eedgh5BYdkv4Bq0hmHYhOQ4szANiCyqkQddg7kd0caLhFfovjHCi29WGCM
nWcJVbx7VX9zgYb3ZdifrZ7XnVfs0azopeCzXlP+k08RKZFweJ37quwG4QLIxFaGg3rhi44XjM+V
TKTCt00Y+qqN/NSgVtCZuAS56y+rXbfdd5bV4eHdfqHzia072LDLrBGh2qSjZ235+C/Gk3GkY/Uk
P2DR+Gqh6+ZmaZYN1mNYKh9q+ZhuiairlWrTV3Ub+XgzhuS+x0xQs1Q30N0po6SNtwQpwDUs7Egv
peQ6MKALkNf6nDXqOOfea64kq6Nr3pt3ZVARILk9U1UnyOKh0DmQAs3KA2G38Hvxau8iNZ5QMeqK
hzxG0td1AwPj0EDEc0zMD2QvHXpttECD0WdPrmAfp3pxI8fBk4T+rJ+oqrH13Qal4cE/6RTwIEDi
sieiT/6QTt78zAGKQFZnC2p4zG+0Th7s7kKVjthSs5XpQnsxnr61RCjE5dOMBRC/VkacDyMrtUpZ
wx5la4qPgt9njgHuIz7334whKVq10BdIta44QaelYVvzMAedgnrGM3qOG8YiY6pwdbEwzc8FHB4c
rP3Sl+rOE9dlTOT4TvHjU/q8KX/eg1G0fsu30/cg1hTOTiogM9OGstH4f0V4V6/7z8f/t0MEMs2y
ZVwS+WVThxrVpA+2lNpdaTt23F4Hq/XHe+nWAG8Y5xwRD0Ofa9d0JsCnRTwPjrKxJm/ngvc71HPm
WHcD1C5lFSC5zY8/47ADSBgDgSg8gn8pEpjG3BaD91nt1ySYku1dBboCxDxv0W1JQfu/zA4fttYO
Bdo7kWQv65TauznhbU3MOeV8CJbAHYYBsgrj1g1sAOGrAsU2NXV1Ur3Wnrw1tGFXOd74WoPYslZD
pd/cgRT7HDYl+1xyifejW0dZC1NQyiNM7i5kqxSQ8vDjowvSBfdOaojxPsIKZHKO3SLywUINpMPN
ywg7Q7gpKureachRic44Q1eMHjHyk4qHLCAuJvQOIOABcZYNkpePVoMPOLIGNBLGudzGjM0b6afU
95YdVAk6B/+5i32/YrMAy8qMQnYdjOpFnHDN2QmF3r7tnXSkWxCP+4km0RTzaPtLLoKxwsERmam7
PZS2MqoM/9c1LMJ9AMJPi0XMwC/5fJoLsViYWyrt9jIph4813SL93Y8kYi0yAVo/PCt7W2Qf8CiP
iaEre4uYU6b4djpK84UQCEL1xiUNcpWA+p3ZiQ2SM4jAL54kaa2K0gwlHPmtKMz28JHNzEARfPKk
7LXC3BzM6Mteoaa9LQH2HrL/CeY87YTGPE1l8hAJqOYQ0eybKtAVnO7Elb8BEz986LZLY9V2gMHa
eIeRTKyjvj1dc3tU2uEadzhvpFGnse33nncFNwm9avmzQHVdEDIbhqPB4RDw6eW9SUQnXNz6oJg+
FNtfwyoKeJTHvwlLFRMMZZLZ3+1suMjQOR+C9Z+cbA25Da8pjZfZgwJcfowRhVBkmCWqTXCDgGqW
RFDDCshv74vyXRdhhmHkojbI1PbUMLCIxuzpebCMI+0pgeJZYBT/w5+9ysS7N0GN+YP/mEPEJrx5
YS8VsEyx3z+cbYUyoc23YDQCqXL77iBdzvogNN2sw113GgG+JKELaRtK50z2PfyPqkzNyT9bcTrk
Sh0T2QVCugvjeuK1rKzYREIXxFcLfx61WBhJIR1zuQTCdwWndRr4TH9AZllW26Qp2KvfrUHLpleh
xsXX7DIY4hnFw9aILfTZtH7jVntasM9gdOBDVcqeHgzEPEQ25dJLXXCQY0H+cXIUaN8oKg8LTkkI
XfODQpHYEAqwe4JiSXys7mJiZuKu5W+1znKpCD/RGm/BdZPL95haa1zPy9G6ir3Z8g4OlU6hOWx7
dXgTNZho3+aXG5vwnjyzTlp82XUCeZOT8TgO5ilmLplxH0SUyGrwKU4wr/N2NMSh/82f/wS9ltCh
sg0pnqtSu+ihCcKys3qcbP6aEJkxTYYdpsk3wOLWRT6YwvSfiJs0pH5ExPOM9KpUnuS7a7BaKUHL
zc5IKWslMcOBKv/HaStOs45jw5W2IMXPR3cJ7WZNjlX88+o+koPlM6cUKcr1QtwSaUZA71u1Il6Z
q2smelfu1vn1IImdi5Qt6esZ2nlhbubUv/05hzV4L5hCLnS7cdtKqt8Df2SmSpNdKLPviwphJf6h
qfLPOl/aOGpGZWUSsCKUIFgk7hdcl0qbtVe9Hs7ZAzHhRNhJZ9luma1S3lcMxDbF8pk0gl8RcTeT
ybKBydEtqJJZdqGSWHwM85KtB2ihCNk7TsoXi6igkaexg2mSL6Z6uCDSzaH/3vcgdC6z5xCQ5HT0
XoDevtWIFjoDRsJOATBbzSNolZaTrkhwLce0dJWHgro6lDIuNkqFAdcaN36ntvwZx45iWci7MqXH
R/YLhrAs3c7cNfJOWzjzwCwZisxrZ/35wz6YLhMlc/eOKfU1m7rVQKAVB3dWsX07g8ZU5/idZoPg
DTsAs8nhNJC5ZMS1yftT29F03ZUrZwLp50piTOUOVPZmwiZUZEdu4gZNhTiND/UcnZP7G5IFXYE1
DkBVrdANUne3krls3fiig1O4aJ+aS+ge898SXMjcyyi2wMa5JOOnBcxv7+cSzoNHtoCEhh91RgD9
lziwfjG9TpoMoYaBVtSNERhncAz9aXijlem7F+DPJXlJD8/z0gzzzRCStAdmrmHam8kX/QzXn3lk
AEXlv1SuLGHfjzreO/Q50IefAjPnHPN1vAptGBY+j+Gh4TE7kCsH5P1gJEMvG9CSxRXstijFL0Xl
rBG5Ru1QMP0Aox7AJcDPWB+xNlGRiUSJ/hbpW1e/fm52q3ijiktNXhrR2Zyss2PyQIttF0YUJNt6
i0lsvTBWilvGaihq0wXvRajBenVWwat1jRBDUgyJiolCsZZLafy2J583osLBSeFzoGrplzjkLE+P
KQ7bGiJrsoscjrisx+lrQHOEbm82im3D2o2EelzOXoNzvmobtwFZtkt1qLmNAfU929TZA7o7c5w6
yH4bnFIEJcHuABCSSfbj4vylTROXI6sou8cPHNx36nl3kCCzE1zxYezsnYQ5mar+rgIMrmHl5ADr
fB4leAOBQnLaR5AuL3WycQKUyZTduNq0tj746btjXMLT1wnVXx3lHf2poc9z/81fe9Nh67jylcGP
kd86481xe/IRb1m3EoC7QFA9zUZRKW/e3EpgD8syrQxspo0o+S9jYHTV0dKOBNk85re4hvPzSg9W
l8QWouwcafbcWFHVF81HKzHV4TM9XWVdtRLpzHKRLJcO35vmOcihunAwJKqee2BT19tT1IjOmb1t
XbTZCEqHnHMGRTYyN6PGqoPPSE1QPMYJdPui3t/wVMsX/JxzNNzIqWWIG+lcevmePCzYfl7lbQi5
GEw8sPEKRBYe4EIhIqLbrx5PlHrLzG30GYW/j2Tpglw6/6/AqU1sPTB8/UPm7GvnJCQVGYASDSN9
NtmAn+7WZSMz29j+vsUqXdC4hsZSKPgjpUHQNYXO488GVgEkBD4WtYo2VmW8eEQ8j7VYeN5aGHw+
QYu8i3q3fTq4KUZy7bDw+nbtpwVF9mNyk9vLacsKE45m0MygTJziYCXRyNKGj1xfWl1fX7r9vI/Y
QnJnUxrXNwCZ28ZA6JVrf79T3wCUfNENkhpLKF0wup6ZEMtE2MX0VPYi/SbsqV3GOM9TUg8UhbBa
lbXVm/A5HRevllxhJAIARlXoelBHITvMhBE8JGqXzhTrd3q7j9j/M0UeJIY/YVe+RquIJ+FSA7RB
3ZVMHe4uq7poS0A1YM8IF6WqSqaf72/mukBeXnmvnqlqA0S0pUmuWwUDYQIuR+0/aGr/I4476sSd
L/jlGLt7hTP4SwWUSPlBIW9gN42lGmwT/fEgVQsAaHCQNm17vXyPKEjv44FfZMighXixEM0wLFht
BQ/wc7e2g2FXdz47p3wD44yixN99GNadXLoYHBJtOdPd9PwhvB5zOOcDAwG33cq/rohNMjLwR5VA
1neZgu1RRrPsGYhtmbR72JqO0Cf8oBgHrk7CCxv7XkJtdOXyn3UY8hwggdWDKHY0Mj46iA+e6bit
KGQIGO1Z5zoSkf6Kd3n0vkBMqdsgJWooGkqNaB2gRzVQxwi7bZW7QZpCFIGzP+lfR2RGvNtwVyRa
3ViqONvRZr92f7qjEhJ7fx4z5xcC5iIcBXmBAVw1QJqrAUJsdu+ttQmshetYh0yyUSZwrWcXmpD6
1dncnL7Dg9G64zj5ov6ZVcqUUCIW1VJ+08mzhYejBjW9EEu/fk70v+88ZmD6nH6N8A/r440XCik8
8U6RXB4nO2HDvfXHiGh+F06blYxDSfS4VLiFl5RJiwloW988/bM6cBpMWaSqnaM5qXXuUdaactGK
7fhab/Rmhwfe7Cx8itHXPeafA70Av6Ko56XPrfteCKzbpWe1BDahFgKWt4j9ZNwjTPlssSXcdVCl
XwJ2/58jb5RYUhVNJlcmKtfSG0KSXPkc+MIQKc38i4ztme5m0a+txIyL4xGWlUOjM3MWLi8SunQ7
z1pMLQajhqh8oQHVZiueqaWoxElaAwy77nPCVsDv1mw2Zb8i4dyfWsd4To0EEOKK1BQc7oyB9uYU
l/pvD1/JvX9O1yXx2ba0tjtPcq7JxCuN+3602u+R1YiJ4WeT3ddeflCLbw4aGFEIPyBbw+j8v9gU
NBg4P12GxaJE9iTNNcjGO8HsWLxsioK5d98UDI4i5ERAXxOrb+K9O2JMJBpesKuAzxT9IDFb036N
qtKBZQwNl85PDmEIqndVM7bXZqHKlYMLuXdr6hli3xy2zQf6N07g4ukxb6XE6eHM9AJcdtNtnDMK
ORkym2W55DDU4CJWC9cx6lwUQsDWXcyRxKaykZZlw4HUZ/pAa8yfC9t7xtXlj0I3g3FF/LRcbSP2
QierrVDRc/NkXhmZSNdl1tDhVsUiVzW6oUszHrf8CNxeveX/EByzKI5AqPeOK7aTG5Tg486gTs8h
J8B05s7HDdY/1CkcXZr9HJLAHsrGjSS4CS9E7Q77Srh/rythKNg+n16Av1bI7/7oD+eHjuPRnXJR
018DW43CtLHWtIJgpUw/5WLno1gqNZfys7AWIWBCDQg2fMluQo4glo6NV7Y60/kDIjwHIu1HrqSC
cvEB0CL1il47q6Y6YjTorpots9lUUBseoDe+8rWkcWDrV5gKiZi8YXCb6cmklj0YH1HAn6uGp18A
rhcFvsbVirWukCs4ruG64iy9Tyj7bNrXE+ldzKrvPLjoIqH454KxgHhqaD0ayTrceZKTXdIMaHs7
Brid7eBzdQmE0wh76sE+AjBveWnTt36MYBaV+jZT6d+jXkRgfdPlkSw1LOSoNz5ctINEs8JN9pQN
BKbfZ30WaW5p/IKDCkgnmfYyTFeKjoXoIdWQaojJp8wgfHnuHemY+sbIC+fsSS4QuBpUFpxflEj0
5LbZ++6tfvACo66IqhPLoXVIZ8+6Mf7uhRMa+Al4pT3xCF+c882fpdoo7k4W5NoELVL26jpjvq02
stvr0x3eWNf9+k5JWafhuLjyX81ffSR1VfRHcJ5KQK19yG/eGnvJlTZg/OYi9jy5bduLXSpXuX2y
XrQTyPuUtYeXLux5lauNCGd+GoZgbEO3L1gVWhH8ObEbDlWMfI6/UuwuncX/mWu3TVFGsaq2WJWu
I1a5CMpR3QA56q9eUZbK/YG+OULfAB2sdK6dXBKI2aaEOqHkXezVoZLtr0YTnVWqGCXq97sppelc
Nv5arUncNS7scHN0G557yA4GuWZ70pVTb5JX2N8zik95Z7Sv7kfUuPZUled24BQxvWuqumtQ5oxC
5h/DAO6cniwFFmATZRr8dOfzdWbc84xRsKXE6QiylA1gDTJ98cdeZiBdbAskAOb+YKEcA1EHtYuL
s01efKwildDGJec5efbK65d5jYyCxrvSHDfJFzgX93QDI4FDnHmQvg0EeQ337J62qiVQXvaXrkjt
qDg5RDHJ+K/hP5PqTme0YauLZdq3eXZ7qPLFkTnSiVXBOH99f86HMENZqITW/kNg4bN6zdUrb8m5
Nwje9Tpl3tXm9WBn6pmo6FS/dpYR4ZJaIPsHq5ibg+/rEuCJfqqzj+zWISY35MABr0Q2qODrGJNq
+sheWXvPQLxPlqJQStjnbxwtqGnKVAGMbfRg2J6JrDVGiRX/Y2FIQW4ldo4UGeWArbxAKkq9pB9D
Tz8InnSDPO+TghHTwg5a0P5Q1cOw2jdD+aimuQInypLP3ocpoBzU4+gZu9eamGo5qZD8QVQK6LlD
zgQUOUs/Re0kqbjz2AmDpkOC+TzlZRj7rxSn5PC254bEkwXyTon3nKsCnSiizyrEO7Q8gxcj5win
9wfdhpWGGaSJa2Vi5K5Cq/u/CF26sNsENw8q5FnBONdf6CE8nooAlZj38WKI05J039g6HaolV8rt
olBwkq85/kba2cFdcoEVWHAxvXW8JLYpBye1tcvNp9Y40cV9GNiEB9KzpjSu/8FGkJt8eZNikPzO
t/Y4qTUhtUijqXp+v55NLHi2bUn5/0vQ2Rf/JjAz5UUBSYzt2vEl604U22XvC/rtRPoOyub1z5r2
2lX3zOOrEyh7XhwtuZh4u5Qh+jYbPVFQneWh5LlgbF7YODFCjxJnhZ3d7SVdffiokXmpNfYSnaz6
z6VSgex4bjcky5LGzOs1KNKLzafn+ICiFx88zuAp948X11Mo5DVdj7Zc1yT5Wmjne4eiiTkLYeXP
A5NuWRyXLawXJ6MbCnfz3ApTT3LI4kEG7qDsTL4lIsZAw4BYBIwllIRAMmWEcCeC75hYHp0SB4zo
MqJsbKmMdkq09c41KH0T7emwTbVkVs0ovhlaDvETBnMPj01DRngXvH37I7ryzmqqtExXNbldGngW
JiwSOiz7G+pP50Wa/DtQWA5iOTxbu8FyiPwz1qEkPlWueU6N1utyDufBe1lPl4I7I54BoFu4QPXj
WGKFdrlWOebEgFeMc1bVk/1FKFlC8jHofQe/FmU1KWhFGCHL4SkZReS3k1jyBwBo1q6e2xLv5PEl
RTkDgk2rI85jSh7QcKIviv8gQhJhSaO4JTLG9oS3/6BBMpcB+4DmffqOxSICE+CVKfi7ik7vMjoT
9u7ThLHN7/wCFZpzjvaypTZL90NdWy8EFEd5gXrAmWorKq/WHUkmz70+J6pFRukLhdXo3BNfp9yi
BFg5o1YZyTdia0zIfooTv2D7lvMfc/yBDudnG4ffoFGpoc7FRVMAGSURkXbR0HT6Jt+UDNllX+Tu
8iPBRup33iwUiISIF+13ZI3wjG1ULmgT93xMeixpxvTgWYVXKjIHw98rqoHMbhgTl3ymEiAcPf6l
QHGd0aEsGLV2YtZC7urrRMl1fQvTzvKqWrgJbhP0cPfM16yp2kphwlYtOY8c7YcB1Sy68lIKgEQP
+oCWn3Zc/GTj+riSqX0z/IrRJlop9WlqFoMLl4X3C8L4zfc2E0Czjsv5s//cCf43RFneenTleI7v
oAP3MtKQsBgGGzR5M0HBWGD/CaGtIKwW4rz3cEg8tzDniKgVMFkhcIcncz92KDEy47+9S3Th3/uX
Rjq3+ZrHZvC8ZJnAtmVxBSpt4EjpbPCZ5EXjyD7GSV9FKI4cu2e89PbQwAtfEfzvHZW975Yfc1GF
BKfbKyfnu52IoWMb+XFKmaSBUcKiKv6hGpZtA65Ul4osCCirGzE1k2kYfixdaMzRHdvr8j0DNZuO
DHfPMlal8mm7Q+j8CWItSxRzM3ayxOkneIK3N59qgEE4YSEq1VOkm+Kuqr28iHs43YdCSgrFU5jw
181/MO0RDREv7GH4NBb2qpWC70sDtGK67B2bH0ldVqZNWjcW9RTxQ8ULGiAzPLL8IvrAfH1k6KOJ
2uudi/XvXriKwNbV+0T5s3VUOTB5hbLcCuPGDutkiuctJd+HrJiUrvoj3yBxjtQToeTO0mY4+a++
wsFjpNgwhi+gMtTRlRWhULINBDDEIrOJ4Y5AdLYFsyVIKAKq3JYoREQbLzUt3F0AuPqx0C28A+c/
VBNmuqIfscnQWWj3NP+laRlMst0EsFPvW9j9BW7QwxfTkgoCQj0oJcXPziTGSD8cxouOKeyLph9K
nZVspu1WKmczHxEnYw/01ZHTGY0mLQeGpu54mHE3TcNDbWuzHX73aWcnW6neXRdZ4P80mcGRHaRt
NXcmAW4Ktfs01ewLww3uuLiwQ+lQ3EnWSQJfbOIdoI1PjDeCz2yEVs7KZXdWEjew0mTp/UpwV3vR
Xx22UwvNDov7cpEQW91xkHLQs7oEHRrQYa6QsFwMUdcj6yy54J2IjL1rPfsPM2/RZbqRQdpYmn9x
eT+OnCe7eNgsPW8f1lcI6wOzwZsQzHb9kd+wVLawHnY19Cvs52Xkwjv6oDTv0IMlFxHKRXhWUgc6
M58rC+VTy2vOS8OydvfDMvVRL1KRKNvRhPrz7Wo855QZS1E0wM9nvWiEkA4zFckluP72OOo23InX
2P9x6/gf1kaygWCfEOYqbs6SqJ/Kgr8ti47sAu0LyPhAp/2cWEh6wrufTHOTTJNl6uu9G209CNtR
0eTkkMk5XCJH9Uq3R/KG6rYwRUkPY6bLdt6ak/h5Kk68ZyzL6ShCcjwYaYga66wifYtUvubk9iKg
hbcnYj5jx9fLMCWGittcbbelmQwbk0D7fFTFV+8zIFvNDGHwGch2JK8WkgFOYm4vQDT9sLbJG4Ze
gLoFL5sTESEm0w9JI3OS0HsnNjfL+8eLWNnKNMteSQ4Bgv7j0HwhtFDPbfnGpa4mtt1v7SXqv8Vh
PYP/Yu8oTjXCw5uzQMhIM5Hy24/OFXY4pk7b340XNned5J49DMnWtcMUwtwwz0/PRhOxe/k7aids
CZa1dWnEVg2dvqRSaXRfhs3CLbbOKUv3WMMlDYdRqdapxhBo2dTYYyoKVbr40gAnbgICLUdEX7Wi
npMckGxIE857/tNboDPIjIw03mjRYmv9dxw2QyEiNr8RlOP2+LAI9vykNVqwc8rAUG6i/hkrAWcs
MkI8cDF13dgFoWZLJsQ3t8g/DvK/glAy0eZfA/tmaxPlMgUVwzi+uJX8IF9mLzzlcRcuuccR9flB
dsefXOWlwKZ22fb2aWJNnampk41QktgS5umYWwBwckwVtnRZy1hHFX1Tu41euhNw/T5mLbWHjn33
/Qa587Fr1T2qc3igln1i4l0tuTEFIM7tR5swB7Z2sT/x4u6jbnWU9YKLOzGZ8CKPpzQqS6QfR8fn
LP9UyNRYorjPmCrNoYAzebyUH6TTJG/8hOfSo5KdoFUQLkWmyUc+A6BRA912B5RcePFVvQeHE38B
ba8odBo7WrwLCGQen8RQHixaM5AhmvrPNfEjGF+vBVXbW6EH506c9cCFCjHlasUnjUYE882/TNuH
uwxJGH10sbU+1uTMPEJozUgaC49AQRRRYGJhSeSu4Yl6XM+Nvh/GJo5TLYbo78buWnmBlGLPFx7e
V/LMcD3io/WJ2QUB7mFV+00WUrW44WRPiReZC3uiPiqZdSwuLzDMxE9PXvJPq6Vel6fHvt7h0ENU
y/vcG87yhXw018tte1363wr2wbXl6KneYD2/GJW7QMO/n2hH5buGS3E6dVOEVB1NOsbqZ/I4SIId
Sn1TwoZAh/JVEPnT8wcKGJ0nVpJugc5vTKQC9QXbJ+y/QSRn4Aor1fyOHyEtCebokaP1tchwc3dQ
X4HR/nu27aao/iSQ2wmI4rYQN7UK/rt+XxxM5o5t+xB8TjWNXJaY7oDxEQKgp47Oe+KgALxhi7PQ
6ajvmWxfDTTl2NfvLxdN75hUROAQFDiLOiZc3gcf6uW7DmHUUWTOtI8L3LLrQd5wDKhySy0i9dep
mw7q/rV8NgeyJQ3OhfCLKx4UVTV3IPDZ0MYZI2c9bfbykpalb35gk6Nc6UfzCOaheJGnWECAguTV
IdP2sVHte7PCS6ixtaBDGoxZ0c8IzDOCw3lrCvJaHzrzjM25O95WGYkMkkR+L090NUNKLH0zgv8T
hVQ4tt/HslpCAMPD5Xvwu1/mpZvHz4LThfN9njTmFiLo8fodKGwfeEJ2fLPtGsbryVwoDf7EZ/Oq
b63cMmWkwGVzOMg3d/D6JMavyvYfKAWIwKlkZKAY+u0cOXNGFcuOgEyod4PsOFYyExFZEb4jzeEs
E4D0uRk/c5VTSriqRGMgGGQn7i2zrwNrbg+HVRblBw5X+CKVbrtK/z4jR2G5stmtcyqZb/+35Ao2
F180iqXb3R5dKbKH69pnEWeI/3iLDxk7EKCkdP/7dR1k9HkGeAzfIFVoSbNXlnDZTAmsPxEG0Edb
bIuuuOpCNqo9bHP3qbM8lLrpyGYFsXnTJh9SQrSUKMdRxoMTpd65CBbGIDTyI9cVYR7v3KZdNdX1
rqywvW1YyNsAd5Pkx2bYkMWvqh6w/0MIUu8alWGKEdsLJe1jPRRef2rTCB/73KBnBFDijLQR/Iq5
eQSwZqWf6bWKOUM1K2HAPOV69LfjKDJJVX+9d8FGv7122QLC2Ukyzi5itl0wGmoU3TtxfbYz5Jm1
DqGDifX/flQRWM+G4aEA8izZAdd3e0+9CUq/3BffvcS/iR26HKNiJU6ToxLYiV96XNKrItuBrLQ6
xmx7YAp/tykmUbWAAcvn0gW3XtyMAz1M4J/qYdKPtQJ/Cf/f/ubpvuE0rRSgFmwierd+2KGUfo7p
mEMjw25XlqHa/hbZX/kguYi/x1MXbWVMuiuyLt0LH9VVE26q0mJvO3f1T0Evy10j9nDFTB2cagIw
NlUE293C11JN3Jdl6curABBYjorLD8RB3LNCy7bLhy6lgnEolcPjzPYZ0+S+s+o17rPoUH9IOEco
VhGUuPDXj2+MmbQwFnQzT/bM+TCbkD1rtrLTbR0WwVsKhFYyHY5n2p+BaXBRjRPKvnjugykSEW/U
/YVepELESh9QTGvkuZqb7auA6H/LVsgT8hujIBRcK7MgWNRjqJuZRDYKGR3d8aQ7ms93uT6IeC4Z
qm14Xq0wpkrGGRGjGxZGnAEtSbnsGhEplmYjs5XW8pSxtcwD84rtpb9lvabnMFnSkXLlk5jfJr8L
XBEizR5/nnvEUeMix52OotV5F98uFfdV9NEgWV353oI84Xoy2OpJV6CscpggO4hZ4074evKVfjEC
qtGKMyIdWxVDv3ZEiIq4rvZl0H46oHh7bFPuVQ7+XhU3ccKRVnNVW3m6lodqWqMusFF9MQApJjvV
BTcQp/o5HysX60PJiIHW6SPHk6GDkBsKVQYqdaQ1xzV+iBAABqwEA3kfUIUMnaPy/VDev4ncrbnU
Q/DzRnDLPBRH8oi0PIoImkPfY+PV3BLTD7oK8/MAHjq5NGsucPF00i6gxEK/dc0oesh5Z7A3iqp6
Um2iyY6Wqwec2EEytwrjo/fTp5YfqHRqBeMT63UlNPXIc0bHr42KLpJa/JZCRipDKrD586flKc1E
7z2vs4iDej7bPXL1VpZmMPchMj1amAV2NotJ2MDCC4qq0a2ViMW8w8T7yZ7OIGVbqL3uMcskhIv1
kLuP24yp52YmEDtVtW929miVXjGfegOZ/lV4D4cEraXRUsYjzAS8O7tZpttYFPtlTX89MaaaCh48
53adQr3/GG1LWYTXzEoaZos8kkmKQxbUFbzgrOskzbewLgUk/NTmFHu09ChyJwjx6A3bVYZceP9E
TLeoUoHFituC3hMTI2HoGJbiap2bZnOpWxcUi0eCPqRr6HGiYrD9w8JGi4yIVyiMabVaHabOuKVJ
3KCRTRP1nH6lM9UUIH6NQ8hsep/rA6JhAGVnXrBVJX7sm2CMajOugyi8VkgVI84jJn2xcksQUety
MC7RFyDYTMkdRjFn6iUOBFEmYZ1OLwOFCtJyy3OS3AHj3ow1caP4vsgW/Gz6p44iG4ONZVoCdSTT
CeKxFDpZXYcXdYhPYV0DvmNN8M9hWdmNiSZtRvFQPHO8P2yuCvukXqc6LTMRyN9ZYfgU59RlAy4d
UjbkxPaJofJ1a+f8tWt0dsXSXJjEst2k55qYcvILd2HJgd+EyZrABt63yGu59gqQQiauJ+1EZHtq
LUDoSSjGjJSYXsfWQL8I7yknAlxmoy6RQy9JRVJE59Nkqeu1WVDQSoNq2YcESYmqv9GrGRXUSNa0
pLmXYsuFTzCl9ipMe8ArLRM+kZ85y1IjLfvYVSOn9CdZaORxCjsfIiyT/HyPjjJTR1Joqrchmhob
piBeMfQ1oE92xEpRyuqR3QLmyaRfoKswQvMkU/qtw51mC6Efk/4QJUF2mrJ1U2a6NsYRVd69iokV
5Asb1GwyS1DET1ZpnfseetBY4KcigUyBg5K7mVrTbtZb/LzroS/VlZYkjCPbcT0lgr68W2WoCiDy
R8mNfKC/ZY0PDxnILaWZ07VQSnR1emUCDpb91TcnUIeqlxvE9YWrkQpwfHYGy+O5XXN6tSt77l5z
yQJqX15PQeBa7GkctD1kTx8G1iODY0RxRAeqXwHZUbXkiu6N2/dYeo5zEbZCH5DT4SduvsvQ7H2E
7UZ0Aw0R4rDhwaNW6SxR/2+aK13cg5BBsA4z/BX3ZodH86yQnjOe8NFxnTFyvoixhNt2sLdMcvlI
BEpwV2KOLxjvsCU1F0JxqCsGjfCWcfiDjInarV6SwjNj6jEp1hapZp4qUweJa7MxH8UCx2tsWy9S
D9v03DyiuIbgtgGItbMXAKGG4wLv2zLLrmzPI328KPDhDA5wa9FoM67STAb8f/1v+luIX81Hng/j
qxYb9AYROm/VTJhvjIJcuWoFnOFuaWGdh3AZbtGigvBUgFg+xMRuq135IlkiIhyfV/YL/k0UoKRk
KbWViof8vtMcYmpDlWOFuXiGkc8ppJxf4oju8rcYq+MO9zPpfRjGDYnsmGjS0pNbtgiARhTNiXZu
ygEnfDIwS/w+rmDbZ0+yhCqqi53HOW0GwnUp1pEdV3pnLVYOT+bhmFkhyCFaMvMGRthi+TkqiLNX
R4hqmop8MDgEjnk8zwRYKS7cRJ8ix8TwMpHknxmKCmsR9u6kAml4bVqha+YuUuL3ZFPDLh2tPLbb
g0cBM1KmLHiIa/pmvtOxYwPUh7jmNLGonWY20z8dZ0l8L3ZtDZOmJoL5aJm6lw6du+7ie2oZ3SNn
ZGudAXUu5BoSB3tzEtyezvnu/XSKLrvesT/StUDEsrpMP9NldTetcS3MLrgqKMRhXtKuPlvZ+xTf
w7p+r3DW9PBlmCvS47W4UlzdWN13Ef16tb9sWkIXjoTikE0jEUGvMHSqHJsnWi7pEmW70GyEZNoa
MMjZDdXlbPny4kRwGEYnq7110/4q/uWiPFHlXqzQO3f3x0V+X3D4SvhQfCXllI93ZHb3bED7knyA
7oP8wHCTISgifuMa/bnEmqja1m8l3fuImd4N8GZd8kkaqUZkBFgjF5+byHvaKpFqMrDxXzE2qzPa
Orkq1yzvpSggpXiJ0q2Dm7tyrVHkegcJ3Qln2sR24ltMuZzLwFy3993ZUtNct6jQzrGJCGOgS+ib
fnbQwjytHs0fo1Aj84E6OcWHIdiFwPCQ2Eq5S/JZ4rlWdk9wpRsEWpOZ/1xdjd4OVyge/K8SeOqa
rJ8dXp+SlBtcPgRGd4o6aeED56MUmUI3ayFQo3oFHiz3jKP8iwWKoXVlOzD5qIBJRpXgHHDtQRj0
WIaJoV9kz/pArJjx6mmY8ooCHe11sboA1k1RrzgAG7SffGln3am/2/LrO9P5/pJhq2AHRxW5aua5
YXp4+VQPb4O4ysYlhq6nHW7jKS4k1Q/xli8DEoMVsucOF9aXkDzEetjWcrCIkro+Bq9iOuvjuicc
yByRd3P200Pc6zq4p46YNnX1Zo9CG4bQ/FOY1qovaKzoWBzqdx8PiKo1w5UGs86tCn+dWTAC/wmJ
NOkPuZuk5gGnbqbR12wHxU4l2p+d7LXvodz83pTiCX5IJTpK1EkebjvXBatHxWYfXiOZUZ+7D0QC
wckL2stZ2dw1aP9znRP7RBV4eMXO0svD/eMae1+1IKLHrMSy7maQxt16xmOEBF7c5Z4eg1bxzwIJ
aNHvq8wqY2CVgk8W9UeR44xpznzuCR1MSSqrVLZBi9N+tY5S/IZvI2iDdOZVgRYj2Ka0q9HI+9+J
Y54Z3rBQL8JzYePSvAAvbe2PVb6Oor+itot4X9Yl4q1lV6NhM30R1LavRlS0vujPdHudIyTd04Fb
8dtuxB84xe3E3c5SI6HgcGFTr7ZGvKykux9m2yqvhUk6O2XvEJEWJhQtsUZ1C7kMbfRhkYwLFFR2
qstp/m4+Gvmdw6J9AtzV9kZnOp0z3F5Z0ceewYNBnc4VKol9JcFnDFnFcauEJnB5QS7O5CozUp9A
hMcW0LjTYCgfciuDukEcJ91iu69R8o/GkjrDe/97XgiXMlascRraqP5Sauiwj0LBhXVt33Hwbm1Y
y3fUYSV+coYFpL0b27ZBowPTevw/mv68eGSSsqL+e61MactchIpEjNJS9VXmqcVppiNidLdybUVt
YdmwX4AU4lX4NxgARARDiZAXBzcEt8yNvYBPA2Rd9ohJEcWeNc6DGwXpw3sl5sgdHDqc9lAEvEL4
2R2HM5D1R9V805UgGC5fTlptaVDWRIs1cyjN3SYGMBxDuFKfLr3t5SyKkFcHZdb5RW+ycrRgtwUg
8uryN+yFWk7oQvVrhchf/btr464dWaVDMFcFu6Kw61uhnlAPAaqfnqf6kIbM/tYYiWkb62LaQe45
bM8aRwJCrz3UCobF/JWiO2QRBwLRtqp2BC/GfALSImsic8JSKs7z04AjEmlaYTMX0YqwvFtMA1+k
XzW8ibHkaAq3PZO0BYezx6CdSpFe3+fAaJ4fqzc8x3xhJ5tx7ieta4AmL8FzEUQk3TR0y7RlxVPD
klNe8FhGgPrKJuuRC0p59al3bfpHfsCyzTPM83THbuNlXTax+b0iZStoHcsrOrpc6GSazqU+ttEy
LX44HjL1cR1VeXTxIdwH3rxsIEQtNdvSy5ITeqHhzof34h7mcIQm7blMs4P0QVgK9XuenxkjvtYU
6lcdPjozQfG8XLtA7jqIScH+NDpfvVDvER3ty6x84I9dbNyDhctHtRqoGV0HccrkkLPUKA0SsEcY
Y2s3SlLhWOScc9PwkYmSDMQtiJNgCZg5q3gdYhCazyb6vdkeAFO6ZCS19jcKeiYHkrNKqPa/Nufy
loUEHusIC8brDAcJC0z8J838/JTnaMy6cWO8h4n1XcBpeQkf9DsOpHXD+x+fTU5O7X+4shUKs3ZV
e7wtJMJhkXLpG7Iby6CLHAJtjTXMDNJaB+DM4/59GnymyZvQGeRclXof+OkbSBTqiwkf31C9/Xld
ENfMV9Pw5eFI+aw4CvGBmwtzFElDUGJDfIvfQplRuLig3NLrQR/nOMoK11OxriScA0TVgNtS50Xa
UXRIZZYzZjXMdwXYpkDgIAT07GC0VuiHJLl86FOKxopthkS20yhoIh3F1elOZfLU31UpEnrCW8I6
0TKdJKVkfLuKqnY3yqmbbynd2QkLmRMSwKTXvpiDrdxXq6d8KOcb8Gez9KhARN12NNya3XeeCEVP
msQp2UuaqA2aW7neM1M+5sBZgt430JqCv7aaWePaMbX1YTxAQiTZGVRIYgN1bqRXQwukKNxlI6Y5
1bFS634w+2YUAfpWQGM38WekGYkP9lqu7zTbI6msUSmHi87oUtgYwCUINywNXs7THA2Oz/tSsu6X
37W0dm2GMALEWHGutb/gKdfzE2kDCW0NQ5i9awXLi+UuC22wt2rVt1m9xeNxYj4vqGHzphM9Y9T6
AtbJdg/lfFUFcrcsEdM5lKGEp5oSvGvkmZtTHGeTCiDDEwhTa2YR43ufUp4wetJipMWhBN4ciNax
Ww4n/FA96JmhElRK/pmEdJEMuvLfKdVICn0RpTydm+AkVd8ge/XSwCqH8qmiO8Cp6tTLGaFo04xs
mD5rZ2E2gKDKJSf5gXJxaVV1LdSs7HwKq1lwfu+0/rvJOeY09gnUXRcS0b5zBNxilVyOORRC5Ujj
tLnCirpr/5KtKYBY3Bg2AOdNu2TNPKai83J3Myt5OtVK9ar1bcqJ6g9W/hB9PYK4u8/n9I2fgZRC
sRoJp6JwCqaptyadAeK4k02gsjeS+UONnu2O/swzZZ8gjW7ZRFWspOv+7VSYX6sNupD6YsU986tn
ZP5wbXaDWDmWB8ENpTyxa8jRkqn3hL4lNfWRCs44aNt0rhy2BamcgfAc+wP5WlMNBA75oWOQLD/v
Db6lh1v0TrEpYikTXoxNqx1N/bVuckzMa4uqgTKRphBE+wxnRy4oE0lYKfpmQwtb+0GJMF0Oa/Bg
/9g/TNskXmSPnpUovMku89uWb7oNEQkACpzLjqg/50fcSnBnCqQUxOzXolA8gUVjnBn0xyjjZHoK
I3LetdttlrgYFjYnUWCiHEG6gnSPg59K6KxY3DuWtXEOdt+KDuua/iL4EIlTSl+x20oKkNB4VP5L
DV6SxG8p4xuPcOeVzIIgSO25P7WDxYTNZzPYdB4zH7U5vgjV/lQ68pt0/vqsJmkdd2JTBm0P26C1
W7Ke/47iiMbPofvE/DlSnfB2CDack33oPd2pd/zexLYBsgl67ixFh7yT1HIskMD8kGBDzW5v8MFq
RXVoxJpbaYAcauBH7axoqiFeEvvJuDjNh0NqXqDd4c9yW0uxHMQ/Vwwx+I3BEBvnJvz69IYR4ulX
RTx+0m3v6+U/Ipj3fJWF36shlM29ZzDnxv+rcvoQpsMi8H1dEwMaB3jnGcsz+VQtA1LFC4KZfPVU
wmJ2+gQn6/eoc2FTkIhG4ZQiSvbRfPFGkDeA3RAZn7RAPV42U/euLZ8p/ChA5khi9OiZqtTNRBdd
38PIIvrk536GO6zLp9TbhABbJoJ81a+wGRx2XIve4XenmIrELWyyLQ1vHJZZVySa588jaeU3pMWY
2v4qZf1N1xPGYsEJw4VENi3/hO4QkY6JfspWXfZIjn6jlVxDjgIoq5EFcD8y9+dG95bolg1amusE
3/QXhmklMsih5/I/iKPXVZOu3zo5cZT33MhIyjNgFbRLj1taWYSSgFvpnXEamb4CWOloXrmqidr2
garhvWRfe5aGlHj1Pjow4zJZTWKzhXjTTdAapRKsXsoa7Jh2yHW7dKdaE+lD+4umTOh0pRax43eW
PHBI8UMqepojuBUzAwMPyalB1WhuW4i0zsVQf/f9Jw+j84Y1CamyqbxLsxi8pTLX+kI88YDiFlCg
x4PdIz194WXOFEmoZiIP2JdomM9sDgFtr5hp6gBW9oJqiiV+v5FKImCAQ+ygjhi4o2anOrjb6O+M
xIN/lx3ijNhtBSZVPa4b3d6O6DcBaX9owFU7Q8fz8nKWB8YS1m3NRQel/9rClfjOQjsOtU8nAOud
YHHAdDMaFJfzSYyo6KxChijpajF0FvdcYHQFGzNTtWq7oICTuwYt0VqmlbeUxnZDkDwI1+24oX5J
7OSjp/bI7Dc/0Oygha8waWfT6skYOxWM0qxUOecMQaWAebRn6oKfkCjJ6cq50gIFD5eGn+K3yNF9
G5lYPE2D1mtc8BtfK+aYwRroZ0aK0wpBsoFDsjvraabneqdCGfcTjcZyYs3XW2lv/Xb7HvooRGne
h2Qupy2WMaf2Ch/aVyZfHYhO2riAHo0jtENGg9kmQGYDifsSmNBqdjfkI0JxvDi3febTChZiDdOw
qsjv4aSBpP5G40h/NROCOs/b07m61mw3zdQnFTt4MJunCMMgGgBCI5NfODuFbl/jOomsIvw5vwvP
ilnwSwv/yI8bG8KkjgF2NLE59MJz8RgXtcWvgavkI74+xXsAG61ClH76tTlz41u+yztcJJrJ/hLk
n0sdIFx2RCH4UfBDhvodEk6eCQmqVH77Hfkurr371tZXLQgEXyje2KAgercNuqdyVykkSfM8D3Vo
rXgxwi+5LtFwYx1OVK5Z+JxEVkrdGcBYrFVoyK8S9pTRM5aLm150+T2TjOAaIfuOT0X5fXivQRZT
HCQh0d8YFt3WoTPcsClnqlLdIqb85L9IaEzggrGSqvKnarX7q78znfl8/kKUcIvYFPpQ91jOg6Sw
4vRTSaH4mEHGZCOTUbSAih4Hc3CcF+WyWoZLYXxWBPhTKtsoOP4vd86URl3JVhoW5Uzz211r9i6d
+Z+QoarnihIIxmJ6v0sAEWrUQXu8rE1oAL7oMMStXiTyyj1XXynbjZD8O8cvMjqbnIjEcEV8MuSZ
OaybypL5vsrVdfeetgzdB7XzlwMqf/kQ+LYRuCPacbKwjwuyHoEZh4qJiLqc27Q0/t/XHGZIOU2r
h2bG00BhpFaJSAe1fTnfAk6R5cWfR0XIk8sdFVZAqDOGdQwIANSzkinW8bHDrz6EB7lOcNLkdGRQ
a7yiRZ7lb5ZUNzq0e39hdklrnCSAOZ3heqK85b+1FdUdjwzdprsAeM02rZ4JodrrS4wFGCopSGMv
OXJrXaBwI0wAMPMG26/3YzhTpyLMHPxsoTdzpo3U0STT3LibGqMg5hfgAtgo7nRAx4HaIeqmkYjA
HDyTkKdSFhIFHLLGOK+fECOqegveBQ/WSwRyNhG0zoi2N7XlTPoSieriELXfdqiDBuxH/99Qg4Md
Ug1mYSaTTzTUpU7YW1pil/a0fTP2enKr0NR0eWi7OGbYEd9ogpUVX7Eqf6qW+EFYkRxxuQ2AHFv0
k62lq8RykGq6uSN9rU+oAdjKoIvHzEJDdHuUN1vi4mwxb86VmpCuIoV4keNJkhSnbq5QAx+bnUVj
p5vUixu/JAg55q9mgpbvEYS5hGoprtz/T2Znu2+NkBEXds8y7XgQzmHYAAAFFA/uvWkFDptuYBEa
oc6Cwv9Y6oj2OsqrBNWUilEATZVLNNyqcydBfY+5I6/ATJFkQoSs+to58bu/jg/d06xYyeykIUJg
CAStGF3aFv71fTEcj+1NQ2CBAF0DZh3YcK6pCvxSlMi35aoYPY0yk4EJ6B/8ZjGiB8buiUoODpHa
8/D5X1ddlFqYkzpg7ql5jtu1r5gNmmnf5glWdOCJRNvT2ohggWCKXVR8AhhZfXdb9fF9dKg4IDM8
P2q/Osrz6n+PsuiVQoHAixioeCKeNOvrahlhovhproYQis56mr7JvG30F46mcyIpKbMzgEzM88g6
ixBARWCRzrAM2dCi6nBoUqPy5p/xY/iOo0//iCP9/mJZyd6dc5pLDnrdVyYTOV4e4vYZmO8z0ugA
3u6tJjEiuhX85twonlcy+Vn1zcBBjTfwidnzMiuOeD1lsFPEU6XydS+Xq1T7U6ssafTCHTE0xNYo
2gcN3Y7FywfslSNag7IlY/1UQWyuu0nlKFE/0Ug3L8FMxd7v4GM0X8sUBgRDs05BJ54kusiT0dMg
BkWBdP2fA1b2LLWtQvMlIq4l4qy5R2a429b4oVoxc5aRUZIGoJf4tfYKn0Em2epRwm997X3kVpYR
4iygaMoRjuJOsIWjxxoqIOE/AeiFBm2ppBPzekzlInrDIY1Jcaq/d/WDquCHhSAe7XZJS4goyGA2
durAzj64iAeJxBTz8F1A3jucdoErjedoHqW7eJC1/7/8ukxEv2lRv+Nd64YNVCifgjQjjW6Omc7p
4KsI/ldcen21Sgm3oqQn+kgTtMVeIk5WXsJaLIYH0cfR+e5z4kGIRHzJEnAFAcFpkqfJvdfy7DDs
UwEdXDJqTofNmBPeejMRcFsL0tcGLRwniKYJ5YgCLqV/CLQB+4O2dUicW6pROSyaPx1KSjzvMXLM
rLNvjNa8it/8lctgLWoS94oJAkD3zfFsjuAMOvRPXM5w9Qmj1Q8M8d7W1UNRcuvJYUEHoghPN8Wh
7ULmJDvchAshJqD8Upoi1c6/UuA5AyO2AMQZ0GKan28mwqco1PsFabrvP/gWBQzw26Sr2CtOqzBo
0+f9SYGffdNPeMCHoEe1d605fQOYXofWtkS/ruLYDS1SuZrE0aeuugRInjuDMIj8ebkvYBaC9m+q
grVmYrrgj5rqNOpziIKCll09CrNMUB2h8SyfajHyI8QKlK/apfi4TJtw6hmN/Mr1M/yJosnG5Nmd
AdP5hScLstCl5naAUfOUj8wgqzuRkfYQrVOZS7K7H1XZ5oOyVE5weO5JJDZc8V5CTv0GmmY9hUWx
xxgIprPRGpoKc46isYdIyMpLPxtb0U/Ftj58rU8kCyL9UK0ZQUJ0MmNCsTOe650j14m6hTPEqKRU
+dzfyv4fzu8F1oeQmFDK657ta0AHl2Qh1cbQJRRP0hi+dtP19s+CQHO/GFUMcrpYaEojH6oCO+N7
JIfpFSZZtwzZ+Z1g88GSjCEBe9z4mcdonkdCFU7Y5FK8zXdw145sYoxo25eS2mF/Z1wsjcDnejkh
YnBoZGxBYRMin3DxKkojPdYXXv98x1NDABEB1crWp7pqgDd1nfJSXyKz0Px2UH6jEOmqP/1N6vuH
VFK0Pj+R5olNs/yBFSDmJnSAQnFDwtxO4NrE2isGrHjif1WbfYzmknT4pzYy8wRLOavrcbLVC4V3
nv00jRKqqegmNjc6P1sFb8V/LtUerdDrRb0SYTWERI74Z4pyn7hOfFMGJNx8TrRZuSd+s4PMxQpG
mSSV+Jgm1EWr1F4xjVhL5DeuEA7ofxVaPOIXlqQ9TV2TwokvhRVhKtiX5K1M1WZuYJo3BAQsEFwc
FJ9exbSkvHk1xje/y3tQFceVUkXAHU7j11E1ufg0dP1orFOy0Zw1RSHHQ8NvPlUPFK2V2NNNS/eK
Tzz+dU8gJ3uu4WI5zYL7GfJE67oX5Q6zylS/jL8x5/81q2Momcs3NE6shyKWMIUDzoHjFL7f0PWV
x6XJPN9MDExAiSt4yEbQI7Mo9Jhg07K+ZkUh57s0TVr/row+AOGUzBhkDqIus/Bv8AW/tMg55aby
tDOan1QF6Lhom0uq82a2Thzyoe+e3DYdvoiRZRyOOba+eaNYVA66GHmy7fSERMMwFyPCZNAqDYJw
TdPZpbbRPL6k58C2I8F1BzrdZMuuRAkNxcqOAOaV3sj1ZfKaIPNUVZ9dS8rEs3FA5bP4czq3qUVK
EMOcjbyFNXLxKf+OSdjC6+V69Y4HG/MIwrrBqA8lAxWntWFNFloiYHsdQwxMVjXZx2OKaGadfTDU
WMdP1h6w8olOyNTTzODP55awiNANZcDf/9mq19CHFWFlftY/8U5GqjhmOrbLKl4M9CqGFap267Ln
vPVMjzBMzgV05rlAwX3hNlQpVL0H3J9ZglnJA8dtDRxRPAcPxDpzuWzEsqbwaKSMiD4/i5X7l1gk
pXfxYGcwXBXQ7/RV8LOa1KEg9oAim5JZEdZFOV78XmAfdaf/sP55U+AvOAesxTf70WZ2JPUu80p7
ZVZbhXPaKRawA3qW2Cn6QMSU2Wv3XLn0yHIcV5wDQf+7u96AdVLMSoP/T+ZXnUN9A3st9H/4oC2h
2keFg4ebHDPrhVIMMpMY6Or6vurC4YCRRP9IfIWOThaQxOj2oRgejUWOrU3qMK0L5AyLb17CqVfb
0Q9pt8dWR+fgkdOtEneiKG+cYez9CVbvIxGTvIaUzIeHHWA5WY5sL5C+aD5OJJgjkep5iLWD3xWG
8z2yu0lqPjERFCeCClSWqqox5+CVb3AHQjh8EIS0w9qZolgOxZ2u1Ol8DDHNzOLtYueuEU6FUJ31
Fk68mYQMWkGxD7LUjNNVMrZQIR1qHQ2cMoVsxHwZCjewCU9Ws+ldaS0nldB43U6fZ3yBSQc9DrKj
mwXBPwBIPl/+tNHFoa1jEA81dw4IIANQX8JI/rAJld9q6NUIuQ7M4LLyNT9YirXduW0OGNrLadHq
aX6Seqzohys7zq/KTbSZFl6xC8H1OHkl8Yg7aguvFLl2VxxEdQ/iXYBTNE/lgHIl+p+B3bNLoZzi
X8s+ISdwJ5BmCgd5JPIyCSbfOZAlAUGY68n5J+hDsex+6q5sZscUbCefb2rAr0vNgJ1WJ0Xz2oMy
na1c+lwARM48nY586kcMDWGWOedYXhrMKagL7ncadMLT80D6eyFd2BtA2owO56Mx6Ya7C1uLFY8w
l0BX3IF9YPHZGEBPGOPy9mL8C002IxKaAQJoTym/TS1jmdU30eqz8IRL8wSx4z2yratNgJVFADlx
WhuAfq7U8Jw9fL7LOkQ5f/clM9opKqNX00QyrZIUTuroq0hVSXdry9gp2pHLcEXZZW5DAkHU/MA0
zP5iBLuZlyqxwpd40tcak5Q4t8rzR+EmrlpgtGyhL6bGod++snpu71Ieo7mVK7OOab8r0suwjGBT
vdLi/kU3xcIgz6NTy7eRsdiOGWQYv6ShiPc9PnpXR9n+wiYl92AUfxla1vAy+p0b9gOY1Av7GzGO
vP0AgI2HWLuqLYVOEpmQz1GKA8+K/Kq7rt8CCm7+Fc8FAYl0xnSFhdioT00xrgswe+xczrD1PAnS
DlhpFvBAkiq9/pJ92kvIPiHVF2BUjyV6PAAzdomy8p9/s2G9WTbds+R3snwmF95zR/h+p4qNylZM
PnpcyQO7NiJHX3Tm0iqz2tbRYM2OszGxN5/SVMW3h7Wa4IoNCryaGM5c9PfyYbd8GZ1bsmehJ8Gw
8ahGNx2HC3aZvl2FH/LNtGNQuFpDTnedbdMSoRDhq2jRN0ePN0WBCQf+qAPNHqlpIKNptjDQSGKb
ZWR9DsM8HZfgHK4uY+AqWJc7gJgCLluO0mI49pu4qMwuX01pThJbUFCDrphdmZPKnem9Y04tPiDU
SGSYjZS1FqxJDpXop4+3+/bl5PBQwtcB2saN+gbwQhXKudT1eM2Yww+cJWQk8y5nSuIkuHF7Mes2
6wVeyxrA5Y+BtCtHEMXK1BpMllOUbiMyyyR/CTQBvj1VM9Z/MPWnp8sWO49+IA3wJQLPruao/0Hg
Zu/qXuhu5E6Woq8amHBQXhYLwSVE0QyLcnv+emnm8pPjn6yDTfcWRRbx5zAxUTQqEmnpg58Wa1op
BZAb+m1Aup1BcK9hiDxpuFyOoaAFnBiIYKWAPOM9kt+CfP8g5xYHdkecUxfI9TpF/aFJCdXwoxCn
cz6ThkGAMinTeY9qaGSyp4D8GTASgeALjghi4kC0+W9Cps7OFLiT3uIq60WY4C69k+odC7sy/sdP
qNKTInK9CKviMSaUg4piCxEImd7tRGEoQdDy7VCrDNfjPneF6X/UvKSzgzYq/+QByFfYHwr5amQ5
Gn8UJ2GV3KLkSfaJu9+R8MOvGz3t/qTljrBueZB1jwgQuPF5o7VkrDSF0r+dkikqp94TmSmoQqho
7r+dnNb4BriIWnk9mnQupUsa/6qXC8IOvE/qnLwuFdMUFTgoNM8ioC0pT9FlDPcAvNGzfzRqNp0w
Veou79C+PbPqgVeabU08AQidMt/cmxMCjlNkm14yMIq7ncgmtBsZKnvpnFMOg6jCP1fTqOFTvN9N
jvEvMScVsNq8ACMQanu5B5xiplGlduxeG0T6nSn0pT4vdl3PhchCQ4Pmm6J5ffBlXKaMjUtwgU4K
Q1L43Hn6VrJdcc9vCi17ID+1jUndih06h0LRwR1LMJFMnXW7lzvqzTDsbfCbqtOaSPv2h9ilMgR6
hKk3JYVFuDkkuPTKxrTbExZJbqRds5lsNEhZQ/vdoTb9Xrko/+p1KkP9f9K4g8AJNm/42fkyHti7
7eyC7knvbOo2mDV+MfdJmZFTVcqbgV0dToARE+jWgm6YWwTg2LWyXC/dJZ0QCTSeL1KYt3qNijWK
ILQI1zDwVHz+mypPblWl1hJ1+YVCIjb4kpIUp4dKYV7RSeumOmuo0/J37KFa+Z/ILXvrO7f0yn0=
`pragma protect end_protected
