// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
vOBM5IekGGr9K12WY8NWeGbB65IGcJ5oL6LqEHK6J5YVarjyngLnVIx+kh0WQzq8
SEZr6RGRG0jaf7jc+z0MhYQC/cnZVoF3dQ4yk1Nnip5VVZC3r2UiydVnAcoYlSTD
VtyQHuZl6MnaGaHfFPqdDTIfEvKKMBEFktXYtbEYBhv6KO1SZRYNSA==
//pragma protect end_key_block
//pragma protect digest_block
k5C74WwFSg0tJ5OcXnHvyqoqrZM=
//pragma protect end_digest_block
//pragma protect data_block
G+pM1M5ApGrsBwiIUYpcik9550l8gZ0AEDyQh3PUybZuwajaDLN5/GCTIj1rxV4J
AnIJaMq2952SmhnGKzqzo7e2B0Yrhgw6UDBsPBwE/sOJmKps1VsFZU87NOX8otpa
PwYO1oHuYY/ykGBTQP1UzWPcyGLtOzF+KPZYKcrmOgciZyv8IRDAXGXu8JhAevWb
NJdag/RzZgrUKa11gvFVQQf97jWVOdepLDJ0HqDW6BZfB8ciBRAj/JCsjPhzcB78
6YtVU1aDxg80kVII9qIr/gzvfVQgUFknXJtZ53oGOnCTjk6xVVgDWRuLnEabw8TJ
ItNNlvzXMextaPnKD6y/o9ORKRxR9C/boeZEiH8KTyXtYLDetC2nSwKmiH3RPl9d
i9s94PoExAj7U0XmwwV+bJ+EF+bKGjd46kYY4xJ53P9OxHFasx8eKJPV0kKmosPs
lT0SgYky69CFKuJRdm54xLkveYl9++dKEXOv/vra/MmYeoQYPH55SG+uvW1/AJp3
Hih/PTefWdiqLzLjbk4XZDB4VKaVYFikEVjTXDapJww6EmESIVaJShqzwzQwCDsO
xWZJxBmiA4nC0gzhMKzDvqXl6mJ5QD/u+r1+YSdNMAc+KBAVsYujQDyQPGRADTbf
fB3u2TVKyY/opkG8++C/0Vo2yczDXwbo1IlyjyQuQqkpswBkzehzi9JNqIYYCdX+
PXkYtNV3kauLM32DTeZxtZXrqTAeHSQB658RAjIJas8s8ArreyjOQwMITlE6S1RT
huYJCVgzEhqNot8FOpDqezJx02jReqezDjGbv7iC5LuA43OCOd5ZjWVJnbc9XZxa
38Uc0QRhG9OfWiu/+OIWDWf8hvLPv7Cd7ymc/HRtxjoLApYik+NF9E31dyzsYi/N
J+65ssW1G8dHmjCZaBOFU0HbKYXOwHbEO2ZSaNP4nrPc+MiT+mCezDPfNw8eDrRG
spWbDOJOLFVdlaP99ruh7q9JPtCq1hoVCRz5piHWHcrOvSz+JoZJZxaPnZRi9w9k
pIi7qvw0hV1n4x9WnlnVloGVxP1dS293GbaDj3GyYHYtnmx8z0lLQ/IKSxvsVatC
ceih7jRNaEBzOOkzYXmokt5AgejKTqSMNCWQPUDS33lNwURrRaMOtJbeDR/QvcBn
kGjvGAx1KkCf/nP5B9zN+q2HTpyqqB9faGfm5vrg4XMVYnwP2TdVlCoNZ1sfrulC
U6cq0pP7OMTOPYs36AmJyCM1qwS+Yi3hXWKEfXeayZOwWXnTkmx3OmX/S77ZIUR7
ZAOX4nsVJpVpugkF0v0OIL84Yfj9vlmPpl0Eul6QPmuEh65n4QEojpsCsmKY51Qo
O+47ZN9k6GME0q0V89+v+eea1BVdgkLCCOqqO2vgpzEhGJ1zJ28eB0JYWYMMmT46
5wDiN6HzVJ7REnzAI9QMdtetdR1TqNSWCl7XnXwsZCOGft9KRdnnU/vIMy1NMzGP
Eho0HxjWkTUTVzFMUEz9Dw00KuEdBq5nBBEm93TCfRhCQM1gpN4YmtZtl4uDVLK3
jRrhYPioRw4UqwYlbgrlYmCIZ00sV8v4gyDNtSPtXcrhHh3mehY+7KlNe4sqY7JZ
6lmop55bkaxMfO6ZaJuWy16R77LD0mVFDzu18mTp1n5TX37qMi0I5qLYtoHVj7Fd
N5msJB4q6H3wadaTTcLPJEvx4CusLlRApgVrfjhgCi7YyFvztB+kLF18Igig1+qQ
Dbp1gas/QhHyXmowvymj9Q/xwE4TSQw8a4bNTpwkM03/KA38B7DntFiTSKC+gmlj
jWWTjEqFUeCXFmKTtBbna7yp4fc53pYVjz9G7iimTOn3kYXcOFjrOnWne3tU82iy
gZ84Vyg4Tf3iWbXz543d3P8DDzo7KhrgWtZQM1U9bDvUIBfCwWHRtkGJXCfvAZAA
xcuygQN9dTpxsujAPh4oDuU5EPkhGkNIy6lxr6XFULqP0jBg3H29xs2EmLuZ5NZe
bTWjDhLsGClQFs7XhGUaT5gSvhEa7kwomDqk2u9D3DAnQ8h4fxq0rYBAcxDCVxAc
frkjn7xi34GtpFz2goGSF/pd3mJd2EiRiicSC6refoIzA5UHgzsuQUUlF/fmtX6j
qRE7IkhHncvPrJOLBU6wO2jr5422USXlXaVzVsAYbsVZ/Ah5RTmyA02q9FujrmYa
QFycHUS08RHMiQJ4ZNnnoL2JF6U53YZ3BIcTjUh8UXKLNxLngM/PmXdS/SsXKU4E
oIpMPsxZP+tmnWOHKD1m27g497OVTYeiTUJ/rcTk70S7v16i0RKCQF3sLHHQkctT
t6MryUeZjQFRZZ84+dTd8fiRQH2Sj8eeNuTdOTdGkSTzoR3Jlhu1oXX7S74BmgGF
ueTfyyO7+dD/Gyud73REEUpZxioWVhr25gchc6VsMeYXDiLYBuw6irTFKEKJSySo
eqauCBib2RBCoXlEYe9XKNkeGD3ZTxIvgPxXa3RxxgUc3b5XJF5YTJzL97Kz4yu9
2i956/xNGhnpKPTKxXMjHKef0a3SPMdH1zw6MygLCLD79dIy7cufdpy8z6AMpkyf
1BUoYAa1DhIH2mc6lRZoY7izmGIzjhcJMVu5Xtg6sBiDbjthhPIvLpEwCm+0gH2Y
LT1YGNY9HaCutHufXbGnBD73IsbhQnEYy5+nzZC3atOuqiWgiJsWgQ+meKQuydeo
6gLkUTh6ICJDRih9p4Da3IQ38U6NR4Rp8pY2+cTHfI0mqxYf/YdEfoXfV4RjiIqZ
LKESbXoKyDHW4Tu/xKZbh0fZEdnpXdCaI3cXZaPnBydcAwdU9s+qqPmvC3M/4jRA
Rg0h8dexHmcERht35u/SLRWB8dBuI5HIXCLldc/M2tYeMoUX7tb9QTmSBbkudkBv
DqGocplKmRdTZ/2cyYdiUQ0Jnq8JECLISifVAXvJ9OBnaMro4wHVhQtAE6wD3u0A
aAyYFTfv/X4N7PKy+A7vM3pWi1gE2ld/D7wmaC3YCqSfVVO1AlQdl7DwFukNErrU
z8Dg73lNuEPzyibeh/fmy8y/ONYBemoFMy8PCV16OVZylQV8nFwo7VEoh07UE2ja
ZCZMODVU1DxWfhSA5lchsQZFV/sI9CFVD1wK7m1TLOjMfpQcKxXgtwoUjs7nbYvf
ZG3V09Y+vEhXJFTqbqn7CTwcUhMWCYbODMnJpbXP9XKbkdV8jCFIhxJjFfkWC58v
qrd8LqnCApryghoB8HM8282VqUMGf8+qzu048worLIpJc3pWV3BKzvPG8WCMywyQ
wH3CS/GuzbqrjK+NqlJlAsQ3Zx/O2PyQTFYJvoHG2h+X5MLayea+yCgf9PRcRBPu
AJWToBoTeq94ESVSGf38eWfJM9hQ85fYQshMM4gvu9/Ssgtj0qt9uR+mE+Fzbv5p
qTFMKDkLdtsTytXIw0nTzLEN23eqqWEt84BCO/NkgCWocCpejVlUVxb8Mq6w7ve6
Z+9vF1qOS8ZDAuP9aEisBwk+zomTPzitA1G2Bc6iNtZ71IE4lftzUsJymboUIEDX
RawtEkX2ycli3GlskPpUZ0Qv6xKobbD8stBVAe4Lwvj3b4ChvaSkgBVi3gibPL+7
nTbs95cMMgQmlwNd2WUExbFHV8W/vh104S0vgVA//aLE1e72mbrtZdKVtPcDYeR0
jf5peXu3uMQ0WOhTTDgHnTbNQzJ2lxvns0X5UubYiqz25LB8gHnl0FeimEMWiB7W
l7SsX2HPB28CPhGi7UA/QJ0awcATAx8MqFLXLjheq3T44JFVcy6ArrWkdFX9ORGk
3cABCTYSZY0Chgx2/yq2Pm/egu1l++v+dEdgKkdEs/F/SgXc1GuSGZPTBAloN4/G
GapV/X4mTUygDgWuBid8Cnlpt7H+39Rw+1ArPLOZya3xhsJcDmPdB/yY+Q8ncuJO
gvQwKJnjPLGo0M1eyO8rzAvNcw8QS/thvUpUwuTv+NxhOxufHAfR2QX1+dPFnmZr
bU5Ivw1LASSJUP/3zfE1iN5C9BcyGac50td1W4aY80kEMG5BOnfYzC66CCFiSc1x
kZA75dhrcFJ6hqGV3kL2xFj6QD+ypUt2EIGolBbLgxuY6OY1oJ4lTABLYHKMlclI
oZi0maR+S1Rrelgf7Vm/xbwL3NlWKBT33ksAFUPOrIdcQq/hdkET099hU7S9s1Qs
k20egAbHGPdxzFs6W2LApqylTiHkNtxZpk3B3Pgh0oGU4Ud1WtYaiUJTJ3gkHyU2
IyzfBl8UPP49ZEI2yWz5Gl+cr/6u6VY2Kzdft7Nl+/FuS3lfVufrjPmyvKsMMJla
+Ac9X1sHZqFT84HcGzLKM6/DdZtFdoiW1WNZAuT9zoBCnRS1kTw3Hai23b9hQ9Pi
VBT1IhqlzN29ZknsNSFQWe5Id3cuYniftBpIV4YWiaiFShl6rQwmnVu7eFLjJe8A
4ZzYXMh4MC4lBg+FkxsprqZAC/+nxVV6fdbSFmwhOj8y1QET7BKYYIrnm2Y6nGnO
v1MVPr07gCEXu8z2MSsbOjmorHP/skkuF1RF02/nqX3nZZRiWZ1ajMJlG3xYOkPv
yVicg56louWCntBBqDuHAjcMmhFPzn9FYRdXPWwQQQN1t/TimDoieTIpnyWGl7XN
XLTCEGCC+xtyOju+/ErC1BzaKsmcKdroIQ4gjx6jhanBqvI7K/QtSmY++FqHrzC1
DGPMikYPsApKKVhn9fc8P+XixhNGRzEZIVVtD8OkzS0TEMRnvb/A/vAWPmBxT1tt
LWP1W2Z2Od4RqN5iE/oJ6TN9GHR8GwJFlrCwcMeL8yEJAixW95PAQs4mVGTy4tP/
3wewRN71mQFAtOhPokCLAGDpaqxLIPEtLzXD+Lp1K1islVlKwYej4buLL21++wuO
i8AFH5SoYoLfXvsqp0MHrWQvzuQmyMgd9tMAC6V6kEToJZflKzJmrDFU9CrFPUIl
aOkOV+gItMlKKBEdzV1NNXbUXo8qWpI59vVnGD7wqrGBTv/Pc4Xd9FSjMKM9MFXY
5iyxU58wNEW1IeaOn9tasterKKNdiX/VQ+2X+jhcy4Dl6EdnJkZs4dnkF79WHzzT
hyE2mKJ5qhN7dLUVPjZqzDxvfaI7Yp3Xlxw8oMoWOUSH1yJLuQRg/RRyILXRJuur
EeNwqwAXHsPBMsn8UUdhHaYC7BG/kDHa7zJ9FGQ5PhZD73fXmiJ7drXChni4YSTM
3bR3ube99+mvTqJOavaA7b8KD7y+8si1heYM+flFPUSJX/GC59gq938Xe+hcEHGl
tpXJsgeZ65eIzKZXFfpuZy+1Ebs3zKsNaXqfPWZqEAhbCtEJWtNd1Uy6iNVjRSbi
mExOKaGRXM/0fDDG0aHOfcSu2pEIHC8eESXQtHOYRZfbLk7bxJmU9ZxuOZyVWdKz
Y38jCIFMzOZ4OEqTa5q2jSPzt30FnmO1RQPuCO3lz6vWsdvpYdU0CS0n+0+5r9ra
GIGmp8OXJJ4LyydZlOg7/GEjpO5Mx83RbqL70yeKP6yEgrEzw60/1EAKrfzupS5g
QS6jZilCA0/QUC0th7/LpA3BmwbxpmjMPYI/2dLxc3M+fiet49MCj3aZQIZgnQu8
7quG4ZlUq5G1b5Y+KL4EbRULR+Bfe9CFjM9fAxm6sh+gXnhU8Hp1QIlxKJzaU92r
iWjEUZGbAE/hfEgXYqwGZUfAFjrMC47nnzFOSfcmFezDYitDIQTiYO+1nPiAcgar
CoeC8oLG4smDjt4XtJXMa9mJT8AVmwBmcA708GLSqOKsdG1bcv6Vu8gv8O/P3aF+
KWbkBwgDLTl5gq9RDseN8eyAme0QwYFco03rtAUct/GdIEoqWMJqah0j7V/yTqYw
tvqM4KkHWM++RqK6SOS87PfT1Jv2pdrh9v0pBZOLFmPe7E8xN3se5KkDitCDVByV
H82zj+5AYy3aWiB/Jo9G1WsMd8guDt0quZ7TUxL/FoM/8+1LnC2Dz/pfKmoqIK1u
Dr6pTn61vsFWqoIsJu7QP5KUFqfRALzpIpSBSUvvA3DPYFrey6IXmo1CFkkG0Gkg
9dS6i8wzTbkQjGTr6Caajp0U645DLhbKGwolJL4BY0CHKm7zZ7Mc8YZjbtZ6Aesf
tb+zMsyNsqV/ysBRbqzWM9qyRGWj02NIocJSuyXCiDJ7B6Jch/4UtPUYcdPKnTcw
itxUyQXlwuy2yJScO9WI6g0XcO77Wqeu6picfBJNiTpK+Y8VloboJwQ8J54XjBMx
i/L4MkhC3ZS3wORUa9qfkFn2uxaSkNT1qa93+fjP670K+iNyVvOYGYw/I9nMCspX
FLeQDgFEfk1OLvzFGZVHHYaUc8AuKF/XdcPP+Jh11EYsrFEVqN1OVdad27LGZcy5
zI0oobyhDdskTc1ws8rw3GtV/bJn0TQ6ZahwZbt2C5Fs4KgBwaMHXbFf56QwhVOH
bgTBo2uFHdSP50HIcM3nxg2dG1Co5Rfd1hXap9FqBPZtJnG/2RhbkjKFFokaoIz1
tZiwPQpq3bMllYOXibButLG/p8Ls0Klm5BoWZSk1wytOCdfrDe8ng8bWftJO0DL7
2fS38v/yzJDAsBOdm0E7oA0Dw5dkHp8R2ebfNIg3LK8flH3JcHbvGzSTsmvmNp5j
j/ZdgSOd2oBZ0jNqubdApb22LxNIkVDrY5GX+p4R6ksz2UqU4FmFIGTWM+WjvadD
jR2kKrra5DIFfF6H+XPI08ebIHwLQFNhCaD0KWRzpGhvjzIfe/a7AUXzgczPcu1W
XI4TEebzQjtN1Pe1DNOAby9gkGDv6O9Z6dmY+/uStASFZTneQv4IKA1XwDrnFL2x
m0bbZ85Qwt1ZoTI6+7usnUdh9ytx9GMhfR1bz7O6+seOTp9dScAGbOg07uVsBo77
RubpSjm/QnzBU0eSMKjqwoxZ2bTfEJgrMy+9xK028rHyQ9FjZoX9lHkHZ+AX5GhZ
6rb3gqrjvO5ErehKR7jZ8wi7y678QOdqMf4dPRaEAXLdeHzAnyO6Nzhcq8aMXrcY
oQne5XJ1zY4d/SXfSihSvvrPUJPqOw6yyNFgRwUTOxmZGZLxKk/CPA4zZeV6JT7t
sqLjCazP1uHQvf4JWq5PbfOHWbwAoYkvq6QxqQZjBNWdfpeOQQzzXyQu4QhoKW1Z
YrCAgZ0AOJ3PKwvBtLDJQ9sjEHFFTCDIJ96+Ld3BC4cz+mg8rOX8Zmpu+V2EASFk
+CHcxNxFPch+qI3mo2IotCht2hkipFIUzlLheLUIQ5QA0UkQ/qvySqe8WWx1DdiL
pCBQygl0zNDsZ0srXIxRIEbYybXIQ7RhfIdGCXWxwg/aEBhz2trfLaOyT6uasHDr
hTElKL11YZ2lQm7IhRsGlg7xGRmYLUMByLfiEKFz0YVby8xYYXp201AEqytv0w9l
LwvZLhapgE7AsRVc9jPruy+dTntslj0eo6pcV75q+7zkJ4YI/Q/fmXpXFzej3TnK
hxHbN8/hyGVKweFTneCD4cpabt3HJ6JIPYibZkyhrP3yrBjGvVD8FrkJDxBga9BE
fdCkv0ga8VLDdoMHA9G4gsIKiym9hP55fvHgfkZs1kvnx14blHhinKtKhqmF+N0G
gtp+DtNxEEl2mIBxWOcHnfkkKyXG84Kg6ejZmMWXo0lxmWaEGKls7gNYfHnnXdyX
1n8SW0pge1BqWaWzLzbUDGKTiLH7taY1UeJ3IYjnoFn7sSlAsthrisTCrXdxXbEi
UM7zsnkBxvKI+wuhjfHK13B3PBuMrGvVc2q7rz+Ols5J/XZZRf4Yog93t1SuY8nP
8nx7NIwMPmjirJ6NJh3mRloWy1WP023FtNuh8mt6rGGLPWb06QIaVflUsNhpA2+Y
+nwpC3MZF3rx5PqbQRfv4TcYwPksFnOlKlDPvQS9/3oSggove2gYBUnsH4sBMIa+
HTRWSm4wx+QHUK7hBw0T9IVMEZVVJ0+eV6l5icd6T7fMvtfDqv4Itb7Wc8l1AC+q
hca/8Pw9xZIfbO0TCEsHYiwingSX08wSdvW+6a0ovj0RWt4fLzwlClTUFNuq96FS
tQ3DDgXZpkuqyxh16yaWz+j3yNMjWS0wQoWf4BsNGUPi+dZIb/NH0OcasxG/0QqA
N9C7wFRpYSrg4GrcbmqGXpMUyKPUYyqDJ3Rx6/qJj5lRguX+mSmQo14HUQpGmchV
hGLzZPLFgHf/PDcreAn9PvKWDXu1Uhq/oZ8//8aI7FNFjDxd18rfcavonnNhjzU4
fEB+XCPGb12wPNH9synyb/CSzQiY5ot3Rr0mf84JG0zJjWsNVSuhjwr+fiSjTjIA
X8nLC9qTnuehtWa+E5Tmd3w5FiPN1h2YllayL/PLKZC3zgh4yPW+KiRm74CVm8yn
Udhf2ksow5DXVjbtnYfpWvbHp8H+5wFxJu4b5y9fjje/gnc5TUHD11umpXH7tArj
cJr+ai0XEJFQX71cAzVO+SsKmT+HBL5K1QbT1ZC74r7eZunXaPWqpO4/MkpeJMA9
SS+4kl5f93Qy1na6/SCg6DOwEBWHeeXdR6UT3pdgJpwcdQ75BGARMYEJ8gSpmBq5
E+xzKqCAPxN+wff0kHWAiW176O/OxjmjZTsNrEGcSSItUfaScIdLyQ5sqL0Bf/nL
YGVQVegC7pRHW1BE6JIfbPFCzGkgFA4wsXAxpo05lIPW6sAMdLadWwU81ky1RWey
IkLBxJmBnacIE9NE3JzeefuHmYDY37hUKESQzV62E5pwZ7OtMkbigDPj6rfF4SLL
fqFs02qx/9IysgDIozkMwNjyhlg6TztSWwdBAosnOyxp0b88UwAHig8hB7a7esPd
1ROsKTyEJ01OfSPfP2m++aRXclIgq96fR9WvDbAUuKtx3MqVND4RweaUC8uZURRM
KwrVLvT+cH1FFcxJQfTqPaGiAhwPA9nZHwY8TP648o8yfZUo7Tsc74OUamxWSxfY
rpHz9UG/azK5LynSotuCE+Vcqt9TSiRHV7Z1f/LOO+10+ZTVFa/7oTxFUXvizz76
Wn1WuwI8IJ1oqqltsRl6/R8KMR5fUOrEHVVtn9wS2YeCAuLSNL0dMid+Tqvflrwq
ogHYICYDuwRP4qcPezC1Gi/sWWuuo19jjl+3mftPwdt7XYBxwdqazYpu34hb1g+V
0mCm+FxzN/yNxiPcZE6q6ok+/2ZZWgd5U24rbxypyU2D//Lzr4FZlZzKWUOag51i
hN+bE7tsqZ9WuorahD0ouNADgAdn987hT15CTqOAE6Cbhad4IXpqzw2ZLQbpVkAd
StmvDKMUwwOTHTqPNuZnHKWnjsvq/FybEFhMzQStFBNLFBu9PvGi2akDgys3UBTb
jDYpKMZ0PdW8JvS4RrhlBd8Wnor22rragAIRJxKBmtayS5NnNL5Qyo48l5HnRvKD
2xi6uUeZXDcbH3AICYTfa1xCdXz6COPPANmWnfb5c6qoFTOjMrMj2arcywxGdxgg
Kkxpn5aloVo78evR8Z1k/fsFqJhWIXP/Vx8/5Rg7fsZtpYJDStQY7bnAReso6zQN
oMWUvuGO7WhEJ0BJwpCTyGIalt/+Sk8gDJsq1Djc4BusJWMviA0sAlWPWxovADhR
JKbMCm/jlsZqsfd/sbDa1oJD9YxqicFj4nrBnMba/5hHCb/3o4b7LJMtACnQ+dsf
l7wtkGZCsgm2zTudi9gAeizqOMFGWtd7D76KEFA3j8WxPJYVDSyeT9dDaZMZRAZo
5PfpSb3iOEc85Nva6KD9XPDM2vrqtfDvUZv7HFjJE23T2nkgvgXhlKOWKbsuGREd
HI5lDEjSfa4cJgdbbMqWJyuShRTJnxs5Ym8DHDY3VSWQn2FyQVzfR0KFNJjtQBb0
dOaqPG0NP/NX33rJmj3eH2EyDbiapp9GgHANbwvy4boPX3V4Vnyq5DArFwABN0nP
S5EW0RJrvB1R3usJcVE89AEVMc65heyosyplFXz1J7SnDAi2LuGg7xz1/lQ70aRX
yOabcFn/PH0ZjXk5rdQh/G3VK+hQTi+MqvLwueN0JNdkGTCD3vAsfznBToy1nU/N
EgEiBqQ7fM6Pk0AgGWUM0uK8lK9N5KyVdzkl8L9ojuTbwab+wpkjV0CtNfKZX5z4
26UMZfeOSDsyJ0ZnbJnHdjUp3Hdw4SJyxNj1H9arv78SF4dnEcYsWMAPSYT91Atp
lhAuDHPU4y0hpaK7ksJBLQa/CQBBwTInE0XKTaAS+Ed5+0Zscpl46PHH8PZLgXuP
oBYh4Xv9RXfC2VSk8Vpk8d0BkSd0BT8RFrGg25qn7oHtrj5FFQ6nFV72ZOE8OJPc
h8hmeILvjX4EMMjYmyDt9aRpksMjWenHZKboY7dONWU1Fm3+CYCQ+suIpU+nO8bS
2cmft8wlcEk8qowakPQjxbwDhNs+po52EdThlrFwtz9ZVyuqMAgm4K8iMXANTg+r
hXtHGvmfJn1nap7FB2m01VipcwO72D4kQaAQ1AkKt4Yaq6EhF9LakjPI+lEwiagb
ZpFScAQ5druboa1cJTDdu6Cz9gYNs36b53yVVrV52fZHXpjUasG92wsapCRxjue4
1xS7QwrkLiXSRKn14V05kXelDs2KWDTGNNfvdo3N0UMkQkLLcfwbRKX8q0CVHo5U
d6DFnXFJYqZcSn3TLBPzieVfzMvW4j68fpnZI5nA52BCowq94Yj0FWk7seb/c3zw
55hruNZBTAM3qGEk9+SFeeQw4qV2uQktDAN34cH/lIjKEmBl/KQM1//+cjlZAlst
ilpkN8Jbp60FvHe3AJoh3ayH9o+5QkLw86d9ATfqEglkpkI9ngenqCbNbtkSq7rT
YAtQvS0pzJyoM5tLFO8HX6ey6P6XpiDqWrGikgXIIGyFzvkKbI2grELFUIrQU385
kpdRums4D8ngFxAHD32xHMVbxsTLqeWLDGgYb4DbZHTUh6v2QEouv7Nwx/EIu//c
t0HRzxJOlVQ2QSHeXskjxM8ghIVBj5NBDcnyHuOgT5M4CXbTACGu6jHhIlFYoSjV
d49LK6hxMSB7bvqHAd911ymtnOyHcuZpEQJpzrjsPzpxKXNX2YGxQMoUk2dy8DeP
REioY4dU+jzRxsWbVd2ycDLxnONc/CFe/lJVOgqxAzX9IHlM5i8pipnie/TSJbdN
3Cn7WJOQaDLUc4WjQzkAGhhbmgtVeJGlNmtReqgBy1BEaVq9ciMS95XkplRoxvpF
k4cSQMTeAGa1nrGpqUx8b2CR3ZyIVVuOAm86QdWZs1CkRe5Eas/z9KrYi5Qdbs7a
OSBNIBeJGmMq5baTPFY0w78qTEnF9nmYxaakjubul1Rty+ZdlQRQ9A5CCUZyAfvW
tt/fSYyM0s6DbUJUsun/r6RJQpJrVmSt0D3gMMoiaR/SpMtPx0ZeK0eGJr2T/GTS
OdHP8wZWXLj7C7zmEUWhewLXUVSHNqzoy7+rOkZPNzIObZuGNWtthOj6dozkm6KM
pUpRbYn0VxfJJ0++x/HWZhzuumI+wygBDvfxZWLxTjnkxEbd15ze1rxxGaB+j5wz
X/pVljp3S7Zw7C7uDcOn1e1LyJv8nHZu46A29wOo7wJRRxPrOAEMHnQocZM8/BCy
5CQCgSSoDfSToHXN69dYXmtQ7wmfLW/r6niPTV5YxEHhFlveCHWw0hQh69/afDQp
CpUxojTCpDKJXDuB/+QlCNKS37kIdpnTqXffbBY/IBB65TjiQLnfBkljdfpu+0/O

//pragma protect end_data_block
//pragma protect digest_block
Iin7ykZtdEafSu4hzyv96hOOn1E=
//pragma protect end_digest_block
//pragma protect end_protected
