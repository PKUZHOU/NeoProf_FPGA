// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
PaG/Bvefwj4t1EduJWqVnEb3LI8Ys4p9wv85to/3mApSPCwVc6/0wDCKbwU7qh1X
Dx3Z2sLr55CyzPRGN2tgX7aKV8mZjzbj08IoBVOOKzafX3N3JnyKJx3VPIlo7REg
8QlnlZekLptZwti8QhAgxcOCHwGqOXh3navIuUuwNY4=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 23552 )
`pragma protect data_block
ZZ5PnU4c6Yk/UlfKttpKtEBhrJe5uWkPRBjkwhB5xeTJp+Utv7u2tglxdKltAkrg
Mwx0sfqUe8jochoLF2mhI6l67qXsbNJ0KkJ/czVyc+Q5MOAOpRS7Fxj4p6/0J7cj
E4vl3mGaX3jx/DogMID7P92sNa7b7JK+6hiU/b0LsEOrLEWwmO31gUb3S2ZqZjQ1
1rTzAr6WF4Mjkcr7zkRF6XTtXKSxkZj8p+m0ivg1FtwLaYkuNxC5/gBzDutQ5wIx
a8a07l+jGkv+zeyX+2N47onVdHqaWSyl2CZxQWfxfsVJbq4hWWgXiIm54gEiLLap
VBfdhxhh4JbPGdUD0sFUatzm1+av0TDmCJWM67GkvvAnnVPPULgi/lcB1n6+6whz
xWy+3rbHB1E+l/nAjI1LLMJiF37k3LNDtAq22XjlKtPI3gWjYtc3VrM+jvy3YhD/
y2s6Q5lVV4uTId0m/n322HlvtYr5tv24BuktgCLBKuMXGMsInJZUlDXLZIEG/I5t
PcMDjXOb8xpXeC7S76YJCfhAt1jbBaHtYsLluHrc+S0bBS+JWqYVuNHlWG4NiOrk
wA4UCkgOCibZ6atC1dGB1V7/ovorNuOQHakZx9kM5K6kqNb07lQY66j7PyIVGKGa
veGSbDFZ+wEh3zhk2CK3mDSUmv0h3woqhginInDrGpo/7ghPCBbdNrPhLjlCsrhd
RW2jPmWEq+KE9Kg+LWSSfmWn/nHFskf011LCENH5UGHmx3XWGpG9EZrvPGclBGtD
deJK+PJlNXiZg8nkI8cxO3wr4zNE6lgeOU54NuRXZe4LbsaLTb2sNvhDU9rAQM9v
eV8osk8Wsj7bafNOxZPDvrhzEyIL1t0rW6NcdynMSBhU0fGtmKRpXYipvQHI1oxL
YyPP/KmUqxd6kb16K1q7o5IVxOzUGNN68H63DYNv5PiVbkzeHfKETgZKw+ph4UCZ
rTmddvk8qSq+K9e91E/JfNLxTlnCFnNEOAk6cVPpBtMad1ZIQ2e/1Xg2hKqnNu5P
lVEviU0N2C3USWqxcp+2K3eqN7dQf1aFXOJGS8bXLCbXVGpnCeHUQqCLTF+jsBRT
H8Al3lMEmW0HbBfn/N8NNglsbsAANhFs8EgP9oRB2vKeo3oYSM5lBmH5O3veqxf0
inZdSMfuIICb1fy1JFfjW9G+VHGEYRn+8GRVQuFL8Z7T9rRBb824xcVoh0I4GrOL
UqxIkmUzV7pNiVNESFThXyEHFhSOAaqwV7chNzhyrKaH69e1pDToluI9NOSIVcuO
scsCs7W7+dDfrIKY7HvKlRUWqCz4djVstrGweYygBhI9uID56ZrnK9XtO0ld529J
q64cStTPE8lmXh9iG+zxHFcIAZZgauDPQfia0OeHKCBzsINq6f/UDxcslAoOTPaB
NUevdazba/EKGtzfSiX3xW5U2abHXt8mXDhoZj+Viblni1c4Vmvj4dgBfvMWDmZ2
HRJJ7vy3x8nXZYSs33VsYA008sTWylPj8hIFL1NK4AC0xQbCbFy4eWTF8IIzs9RI
theHE6vkBGRlvQvQ74tOdeApQoZRFfO+9n0JucP3MIiL1AJP6/a/A39c2RU1T585
LS9KwbkXlshxbr6kWx7WfwHsBCGIoGo47FdMU2tPquBn1LFkgsrlCuq55OvyBb4w
7NA4tl/ePR2tZHvJ2zQYXlq2C80Goeppn6uySU/+emv7pd7mZvgai6mjaimkmo/R
e7mDLBmPtPxLNKY4QYF1C6n/riEUWINWHYp4pxuz8Bf/gdZ7fCTT9FF/pEEqi+/w
JsyvTg+cveV+RHmd1YDR6/LS5iiB1lPsfGIcYUsQAORDFdRz3HnCl5YA0woreOYx
UGBZmsQxIJOu7hefpTG+XUls6n58KxkmHDKsWRF8rkpyyFQvsX+g6bRJSswb+Jh1
ndUbAo2Kp77z2O2KJ7TCG++N1Zm4q7f2GYfPRt+xSAw5JIhCnh9FyBxHW/T9OqtF
kHjPmVXGmN1jdPCE5NgWDt4gntX2S5RzofMX1n/s7h4uGMFWWwj+UZGtbIPhbnwy
77Z829GgawB/Py1CAVQUpoMyzcr1A0+RADZsWNQvivxdojUg3m5P2/d1J7fU4oQL
RD4VOVkDXN0ZU/gErGlXhFcSD4GJ/gstCziIRVXE7U+KytecheGB7PgVDEcH4as5
BnbQhNFukRqKkoi4x1HxUpzmCXPcGScnKF+L4hp7ZCBhkN0yxoKGbiPykaYaF6FE
fxlEjPKr8n1ImM2AkNGMKBThiLB9sOb/4SilSEZl7LMWYiJHf1FRFa4QgEZWOmA+
zRTBVtHFLRvA4DPvmcBiZ3grA8eDvwEn+zYiL65njcmvBiBouUdlS3Ex3UKc3GrN
09MMN2fBdpIj9ZesVvDW/u3Jj3+pJitB+nmw75NMLn+GMIh/zcCbk+i9m3+Z66hX
U35t7EHmXINwku3dqP+D91rpYGov1kSSWYi9L6cUySlKTN9kcLEZEYrqcAnIH3qR
Tnu0kBWyK6syFbEuBzqLHW1uu/K4t5zu2EPUmP7FBsIctSbvRilwMbCjp+BU1fhv
5CUPHYWBH5LRgbrDFJrfQ042Rjxy01Yz3mQWt2NN5yLtoFCEpGxvD3AfOrb3E4pj
MVPEKbHNRuT4Ai3QncqPdzeLYVXbpzvbaALGkwunYYPOWUd9drdMhK4hdaqo23Lj
PB9P6Hwjgegh3rt/WjBcxgM05d8A5HOMfbcGndT9r3VT0qC8moMP1wAtYWOstFSi
adOtJvnTjwQuRJ9joovBd+MgQzI8lujJjyS+UMDvZ7Y9eJiw/MOWZC2E+EaN4wIa
X75HAHWhpDeWVKM2oR4q19CIIeIVMMKzeZ7KCSFp84DmAcpylk2NyF25ym/A846P
XBMIYT28BfsKlackEJ81xciG1pxzhuBB8vjVBT0xQkhPZI3RmYKCtjVb1DVIKLwz
DbvFB1gdkE3TkiOqkO4IHlXAeDgepe/CEXlBNJMHA1hwF174usvC9fPzUq0tyAEr
KE12pVrrcIm5PxIhUunS8hoAwDhX3VI/IwxwqcZPtHRdVYItDSkp2WXF7H1JChFw
Cudc6zRbhA2b+pyz6DYJ5/G8s0UQpJocmGXcJbujL93VMQa3UxOjeA3Uwt8xsZhy
DNBqnusLdXUH0Zkl6kPTuhyksKw0jkN5MhNUo4iTYM+gPT08ROwqxQ5BJJ4KerhJ
0QBzB8aJ1V7QAy510Gk8dtVGieKEcnhs2UOOmMca/jPUSbOUR/l/viyRCGi1EIP2
X171doyK51cig2zcTBHJNfZs+N9cNo38apHO0UyHcWGHCsqKvYLSITgt/4Cfysec
MflHHr5ZOGvbijv/cz3XJRqPajFZLShgv+xRXFdVa70RK080njttyYLw/Rhi7/ca
l64dVJC00Etlkei8aM6p8CX+zzY/VAAfDiQYuwgbwzEG+yZI/gqYTPBUMM/gcpY/
Fp9wsnZY4JjHvwOlwclVwWPcTTDw5LitAh8qp4jSDrZ6/zukDyDHmJnQ9fyOtK0R
ewGtKbfn3u+GE+2PDkBeUlycdatjcEkX+Pg7Q2RUYhxR93glb16goBjGB4v0hFeb
+JtUf/L9MCxtkA0+FsftMuEQMkWOboo/OWF9jIX1Vyj/MT/lmcVtkaIoxig21QMx
HvsDeBZpeidMAAny6rCvEcAJ/Yg55blToaKd2TjqJUcjEjPuJAM9J+RG6eZp4QEA
fcor/vj44LcXij2nwoxulj4PVs8Wv1LBTTMVNp8ZWzTYOte6Elfts5lg4O1naykU
da4cz2oRD8VbbCjCf8bo1M1f8meOCt7KOtMUEUSC5ogb08BCoA52UNEKcx4IZLKG
xE1z/BWq+R+6onZs+/osDIRD4mUIIfOV6ALEErQc8pbiO1zWcKyCn82ZgNqb3iXO
Ktgf54LHu4gnZmrqlpAbb8SKBSJz+AuGFncnmtDrRiquS6UiVLpls5uZEb9s3QIv
rvkbgXroKFCpiamQMsp//aeh5s+FA0hxB5ngtLF4gIIEHaZ5m1KKSZLu6U2gq0iC
AF2XfgJKQPhUCvxfzoASH/+8nAbl8IxggIeqFLjsPxdMQGgSQIZc81RKZ/6wxccX
RrlrxNplzvdP8e9PQUCpS4Uogs69uNtgkbaXJ+qsYXbO0jAYKDD0SgwjnFrcDeMx
/mNBvetdE8V9DohwHCQJQMrg4YRXCZUEahonblG3UVivb2rWyJIdmNmBCsjfuorz
G0XCjRQfPIQhMEAXNewaSFoUn2UGNolaFYhh3TWU7tlXBDqc6Onp6depnQoW9pdk
72ErKxUROFfelUE+5r6VdHiPZOhgiQcMfHRkDDPhqltmKJOof9++GSuR/4YyTzAp
R2OwcVhQnVmu61qPXKghVV7hbFl4dt3F6djfuRff+IPR7zhaBhBWP+Y0pm7kunkD
3w+eefocGinoTy7chwd0Tnvw72yQoWi6kHvAWWaRp9WJpwQ5p03v0YDtwExLhbro
unMdzupy6KCOwjrVCGnPYEeOrN/3hsBrH3Ws7SCIx5Z2whszBnhDbRV4Jwkv/cYz
7slaQaDhIeWFErtAQ7iUs+LLD0JEBGe635AtmseYSrrPX86+sBj89SXlwT4PwJxJ
QXO4b63fZ1U6JIwLScrCX24tJbm7RUtmAD1O8LZHfQjba2fBez3rIpilfpv/PA1c
aGnnzfMeSB8OuNhIUCI0tfhXNDTdu8r7T2YO1Y/5wpe1nKJLrbX3IWKc5sfTSWZt
dr1hip0qEqUmTdTvIHKXj5mCicZ7iCmXK84A2yQN7MMded3/DE5WlLv3FUkivyRN
AzN2vPGvGDtPV5iaXhOUbY1d09PV9vL+8YfBaTxKliGF3O8u0xCm7qkq+71yfbS2
JrVDzJXIPY4c/UiewdyEI4C1H6CTgkMKb4K5zqVib0UalzD7F+ll2qE+/wrkiJZc
h7F3RwitvFOxfduqUccfA8oE1vQzTOfEBRJhb7gvEZ9NS9255ZkW5a53372O1Qyd
ya8gaAj5YJCkL0v29GeX15Pbiqo4H2LOkQBhJZJyTzEE/yOTDDlWTxlOrTKeRvEa
gTvxJ/fYwQRPjeV0apx6eJ4oWvGonIFhWtbA5EQZRV3xyfnPb7E+wndq6RfEiMWp
VKuiggpdOk17+/cGCcyFwPhHCRP+zrp9EVJOYDLDe3jJ2qEeUCi6KGDtueTG8lUj
GNLb2YlkU/yXzpGVUdCvHEIbeilBHJoQs2Gw+2m2uUxN4wnP4Q24rBwsMNfU6MMQ
y2hft1fyBIen3Z8pDmqzK1ljSaOIJ8b8FAEudVsPaLW7d6n/kOGdL6XTg6e1Li3p
J/HajnirRUHkhpoINXN5YjSPLIzHs2MBvyUKzzgo7+qqWs3jC8sUjSz+WHEo2tn7
Gedn6/clkdCyLB7xMtZj9AaYvS6rR8bt8zfN9yyJg8fK3CCSy6jHu82S8EkYbagu
VpBEkP/sVwBu45ewRa8J8jd8eFzenaMwy8K3O2DSnJ3Xg8nxVrIiP6QTafxEB+Lp
KGemKX0psaYg+pxyC4xuUlP/Re0OlrwhcbwZJe/xJVbsRQcoJdj78VIeqHmhJ6ZG
u1pPlXQGzAewHhfIBitrNCtH2kOa511BfPBIkQzGCJVN3rudojUV+f8GQ6vSBcCJ
37QxY45eWa37vunQNOSiEiqKabU0NVUO93lBWB7Q5MoZdrQOTlyi8dVgAGEmoZJv
XPIPj4Ndixba30M8FahILYQZb4OCYdPRC6cztD+sgEJ8T/AJUX6/GvmUdxRE9oQS
RcRGDQvBECjXEMK8I61yein2TNF6WpDLxEm6WiD+DSO+HUOR65+o3jv0hcn9TaVf
s8kX5f/2R3S3pOazm1c8yAXkU5EsPDEZlaefSPWy9Ilp76R+u54n9bVgNw8qZ28W
pUD5zXrouxNzSqKrf5xkIK7/DBcg3XY83K0jvM81lQ4gf7Gftft3UtlrBm0CfYCJ
iTWmfDPZ0daJwMCYp/Ky2jxRg7BhvHc1E8eKxBYM7ZbxxFm/c/rhTCIjq0nZG137
pWUjJgxuprUoCvZ1YszowFWx/9VCgl48tp9C5yiePTm9iVEUfwNxIKFKGbNIF93+
Lk+QlrNW3viAjQPPJfvfscrcf1TDOqPbh6JPtxaetPshFCTeynljf8tGh9KGC5Z6
IBOyDPeDva4RJ4bzBDNBpRQYhkfkqdqYkmWCmKzpnadKTc8zJU7QrxuGlOsiX/gW
OX266qjwDHTB0ZOWGkB9AKtSvTHCmit9raQPPbPrnfo6bsrnHSvycAb1iEipDmCG
zwQxLOM9Rf3vuBQr1jA8pmdv1TjdPoLjQEbR45kesWOf1ZMVHhd9mDcXQcIwoFNH
FbFSX0kIptYc6sRvIIAGEsrhSDSl3DKe2DpcdMkDQIRgZbZtCSBWyqQT0TlUXQOb
/FVn5Nrj05nkeL7szd72CzjlK4dWNY4nUCWGk9u4l6FEDNkjGorTncQQTJTK6oUK
nDcpgHR880u4x7i7b6NRl85+4Y7VkwbapMW9uoGuOkPXPxWdMj+2tJohLvm/kSV1
o489zbs6hTmyBnWrlHiMMGnobJ3jPDCtClTY+sc5h7mX75i6AcAP0MwzITSuxqEv
XY1+ZdSAuBbXn4DCQ6xIzjX0ZOUaJcvUnjeN5h+XdAAffQrrKowZyN+2Yy57oMWO
7idN7pMPZojQXx0VhvVn6bhagJwWGPZHV0RACWRuZpMGSBOWKLHisEyRFGO8coPC
wEbzexNMM6LDUNQHazOI++n9wRvRNw4EIRpZB4kLGI59XWtMm7vDB2Ncu8auzh1O
o48HxkN6ZbrNf6FVB3QbljqyQV8zrC8M2a3EgeRC6WfScJ8uPzDZwa/+EcqB6CnF
IbKLlewZ4IGo3EqJY5ixjSNHdPsDjIlPbET/ZP9hIsGtqwo7FVJAyx1dXi3GSvA9
3bW4B1cqkMVEXCQkAzlbAeveqjdBrZgjMSRGoJd+7y3kDw8vqP/P9rTi1W5QpCKi
OLziFEnVeoVVaxBi6Q1AQTVpaImB3h9w0TMiCUR9IkriJOACpkkuMsszZFD28+sX
If4MtdAeeuSfi50Cqfz3wVvNokEcbBAzagPNSZHK51yFaOk76hD6rsb+8uTWIgzr
GKPHpbiEJ+6+JIbJFzk5zqh1JVmi868cQ3JFyBrDsXTZvwFzr1ygpihJpITVbkBP
KgZW0D402N8YALKvNFa16YdPX+RPtyMEzNNco6sTiN4UTgsvLpW0A7AFvK/zFmXp
4fOhRel8wHssHE9GC/nySQ9Ps3b1mjByYPw54nuC1W1XuZrJGVcv60Ekdiqq7xJU
mN3Nxo2JIsRXPyI4cNKjTWqLagm61RulWy1v/lHNby7Cvvev0WbfpY+STmFZYMNJ
j1laxhDAWKNxxN9gqCKufDfVfigkoUklyZ/mEed7Y/KS4wj8sWlI4fdTHtMcJLBw
8UMhN443LHy4i28zjxsVkBXzKwr9sIvZ9arkXWJhcE+QDAfSm+EGCADBiJQ213ux
I56+dVUsb7RGkO9+wXn0q2jZ3G3NHFE0vUmMrJ8fYgNjtQZtdy5W6QYTcTPfx90A
KztoEgPLjO0BlF/bVBZuXTLNVDKJLvDnA+yVaQSaF8nxngau+zyoS8Aq6sFw+DxR
hexJra1eKsjdTyIXq/Em4vrvKUqKemLXa5zihw21CKaA84/1AmDx77elWabQYeNp
eh983oYqLAdrVRHoOyv6GoUZDs71+c8zp0HLJF9ZCpomhYNkpkt9XT7u31QN9LyJ
uRRZTBAJ1mKwenrNl8xVw2QhlSEXpXXVan6oX7MMabYU90uktknaPH8IRpbhYBJN
sdDN37ApOa6qLqEN1XOD2F7RsHSB5SYMGrEbgQ/MjwU5qEM/oXBQAynYx4N/a6ca
NecG5Bm0T8whGUz2D3dkXx9zjtuC+xsRKP4Nh9YmQ3J32BYsJ4+yY4QB3uBR7vVv
uJ94sgUtbTlDFUNArtnMyZ5KGZleKfAr3xaVpTVQ8t+MQTU2jf+cP+alUOryTe1A
ziFKkigtW79IedEzcRU7CiQXPucjBE/scPnqxA5aGUNUBtsDLw9x1CEElzBo1cLs
CrE9umWGQ0FYApvorqpUkouG0v4koo0sKwdHVyMCi6TMMSarUCa8grV2CFBF2Ff+
psZG9OET2Ii4ZO+SA4Sq8749jqyXNaz9EGbH0hxTOsZEOgf8zoHOOq5/q5J5g+mV
YKxAmCStDygvOSVY1REl9IwvmzNgtHkjiph61GNRmwqyxRl+SjmY3hXgZjFDKiZJ
ZCRQhGjLgpvSsQmQY887H7AKXOO82j3Od5QuzDXi7cRu14x0kjgKk6aduG5JvS4S
fAqdBkr+LjzGF5m+Ih4fD0PWFQnnqxRJTRcQkqWNtn1wDoLdNwq946qY4djqqQed
2TyleE6L4WdWcKgquW0XXbXQydRaL3A4fsCLqGrSiu80vvzYzJ6nmteeUImzEuKM
oQ6+q0TrL65Qu6T1O+fhf4O9q4bJDKOqyuWCIrsvlBO2DYde0hNrYle8nxf7FFD0
WIqk15kX33Npc9RbXkYZaJHX3gDDx9mJLfo/U6tCnt2mFyVkHyjaSXy14eKmqce7
OsqhI4/v/llDqbuhFq8nkVQrS5ay8K/A2+ZV+gHS4C96LGqKk8G+DQ4F0GjQ6NfG
PuoerZtootXMmliaS1ZG5N7/hTKNF1AC4dTa4Hh+WGq6GVuBMlXV2c90EUIytV8B
CsA3e0UhoCZz4Vf+BkfPPXubya/+VOHUUWLq4jKKup2ft11BYiHa6h2EXwVnM7xG
uabTG46BGzLL66AKkIb2Oj2zZPVPl8FCpg/cbIHpk2SP+uAHY68puRtzG27tk8Q+
Vuzt3wav2IMQjAgRt+tiediwusukl1ui8ZVmtMklHBX8bwzn7uHOfTU02ErFtUtn
esjOkox42hyJpNXdSxPG09kqHe2cQVIJZEmQ/bTTgHyA02y5cs+vDIHs1XkI+l2j
tCXNRL3CKt9eTOTgU03UAbaksAZCGSv5SCRPTFe8qZvqsxcwwtgIhW+xgiok9SW3
VUb+1HA98oYa4EkplcqKgyONHq9OcvhVXGk4eHJrZR00lZUEVlD+6YjYXSf+v60Z
OJ2UKrXXrMkCVj0sHADhvTeBrxBkA2CTQUBML8+roxk46eRcVZek/xuk+e9VTJEM
MzoeLfSisDl3CsP+EaL0wTbH+RW4HrZKtE9Rz+yLWjuoPUDC3TgjbEvW/LyrXGr6
dwRZTY7gGOBg7aHDTgtR/pYQJsbvr3hLQ/ROEasdQPyJ5mlSxvRysATHZok32vK5
M5RbX5WpfPTlU92/1Sw7Pm63xWOVu1glEdDIPFhiiFWEuRhqDbMpTD7GRJOPc34i
BiPwZabfBbVq9RBJ8UT6X/gdk7RffNPYSJPA2isYQOMJWLlIwl4We0Oej+HFSv7d
w1x6U1U6EiHU5FaC86MIJahJKxO8cu9JYnNCc0VsNSSTgnMtpo+2sEjrHlNfVQGy
v2JXONsqTtLayuGh3IlBqaBUDliwomlzjncpbJejwxTUAL44UC+88+8pphcYe629
SndvOztvtUVhJ0wwgSSFughwKw7QHwL1LOoldVDIkNTWTeBysEGxloxCs0RfSLwQ
yaMTfqoVUbUSKJuNR3Z2c9bo3sWRLb48Sxi63ofgyy0p1bEmjrREz8PuQcSf3s5r
Ptkn5v8dcWobU0Rqhp0VldmKK+xl8M9Wwlrzs3W1Ed7I97Jjfqu9+uS7joybJ0lQ
SV99qDVwJeKihk5br0SBwMyiTBY2JPHf+XvjWbRAMI2bc27rxlEbUzCbWlFpc6Af
jOnCbRBaKuMx1nFhehm5iJjj6Y5ezGRzIjGp4TAhWYlfKqjrbd8VNKXvDj8b52kM
cc6/704WW63dT/tzpzZAT6oklEgttSWqVGkHBZxReI+iYhgmvD6I+Kv/GlrgIG7X
DMakf0ZmyMgiZGVARq4Ywv5cUpwATUtpxXbXRpCvY4Otga8I5bZ6LNAKIYfDG0px
vp80TkFRbJQpaYWseWXF1S30Xp9RFrodFaTzhffAsGSB0LzOKPwzXEOTK4Nz5SGl
90X745ME0L+m9g/H9kIVFgMWmdgVFq2U0lVYPL6ix6bwZbk2I4SgpUqIQQCdO7ww
yVL0iCm9F3k7E6y0Dj/VjfBbAkoPoqo2z4jqEA1F2NkVE5WKzOOxGbnEcE6u7Ljv
Jf5nJiWVTkkgSHMt9yl3vLYri8dqmZve6veO+UxnQfsEvUPS3uG6SGkHv0VraAKb
uZohfJnIXsXdI4IWENxzhGWDzbkr7XZa4k8xCkK8Hqk+pVCbalVthITRQmqlFvvG
YsXg5S8j9+znQq1hKwE9sEgc6kOsuVMo9TXyVmWhOFgTW2JchWsQD+iB/mhdWPDZ
JVntCtdh9V6p2iBjEIVhBd7c1VNP/Icc2tdsSqvg6Ejlb3vzSIWz0EosWTrQLmN3
GMMdBJ5xRxmYHHjkLi/CDUBQRTZA2VLnfXlSp+KQD2ntYWGIFHFU+LXUVkC2c0Ap
52NlCJwg4qWA6wWkPWZeuZtDfy+LJC1cXNEhh7WwDuToPJU9gQc6pkTuc0XfMrbg
jUEOh9uRdJlDe7rHm/ZXfSwyDAYl50IeB/1/WX0pMboYbjeambIizdnM5FE+oTmE
1zG4sqqeG0US9AZKQy7mVdhfuHaHS6ekDiMLTV3KLJYiP2WlbT0ChFzmrQB7E8zf
lg1iV9HzUSG4UvO69pcrUuQj9/Q53YrOd5389A2Swg+sUwfanFNXzHNz9LUaj46z
UTukGYfD4BORJ53vctSFS/vPowJgS5NZpfiozN/p0N1hI00cefrvbQ16Cm1OhtWY
m0paOUsa/GC8LNYbtsH/cPoC3rFp2j+ayAq5/YkmMM5HcOH/l+5dqt+WcgfRvIqr
j/4tfuqTvg8frm8DZKwjajqBx0c2hFtraBXWGv9nOtfeWzz30u53Rh+vUNNHmUNN
s+gbqf5M+riIP3LTrXD39u0h6vCG5SCQy8EYnxIjXfQLkyMjGyLlcaq7H2Q6JRQN
dWJ3h8evQlTy6/wKVGyYrpLf2+d6sR70zbvdh2w2jiLX08kWO3223wYLHHMwlMhn
lgmvi4SggeYzSKB9bJYQUFuXn+wDVuHiR4E8+Z0xuN+rlworcCmaGVFk5vvmmVIu
4kDBOmq+4HNpRyIjbz83vf/3y69xtyDZHRE9mP4MS2fMa73y0SBQSOMaBH4L3qx+
l75wp/9jmDZxe2Tax2U9SFx/Nlj/haHCNeHS7QwVuKtTr+YTWJkvUef4U8eLlcGs
zQfoSCTKE2pNs2UqVQcfKK39j0FueYZuvHBHWx4kmukiVolBuLcqPLa7zN0Kd3Xd
dJjHSCnt5D8ipIHMHQM31N8Mv/zp6YrPyEJcd9GQ4HoJKGnE8Dkea6uiS1Ga33cG
+FkIPGAxpF1qpBTb8r4X7xzV39r6Z3ePgQaH/MzqwysOtbbP5z8mtQPs3gdVz4DG
jCqef2ex1iWt8lgjzhMVjCZklQwVvqD07s9Z3OJMfnWOk6nduAGz/DvAHH9ndmPG
PTFWDSpMu7iSW4pzxCtI7PCr6dQucxjI+TLVxhQ2SYTZ7x6UaiU/EWELrfi7KD1w
kcyb1UQEDND8riTJw2i0kTYpGd7E98SQlPoYxvAviibQ3+UU3ImYXHKPQHM/5pZI
ATbWDQjzngg9iCXA1mFET+hGwHWmLLxNOlDRQUA8bAa/jIai6B2EW3AJIu2uw0jN
v+q1s+vGiJfdvdmZUdnBKg5ZtaTLOeEsEx8gNOm9NYQk+hpvyTGp66aHbxcYj8X6
g2AEsXAork0wNHwxt4rPZeSzdv1W6+FEc8ImuGAt3NPIirv9m5C73YJ9gsXkbn8k
MFfij1DkiGQdujB2lBJEKYgKuyKmhe0tB2mJTCHSqIuQ/L2QJHHVGPQGquzov0kR
6Eio9ySeH9iwGi0oaVLdz+VUcFIxd2iUnGYR6A/BWmMbd+9qq8Bem7di4YUkc2dH
IQcCXv9lhxyNt8Cea4vj2E4n1I0cfPmqwnTgSY7JtLeuoVtEvf00yhMX/DkFxx9Y
wM4OToRyfkD5Ry2eghLZA5qm+7bnyGOG2FYIVHHPI/ULZPBQF0D85QmBDi3iRbBR
rAg/DkxTA/+AQGpGRKcBSCTFDDfWuvYFuerTqevUXAOtxaQVt9UndPmsd+BdmCpZ
IcoQ6qnk+1rEssHxSRr4pX+YxokOWPFHX0z1Rxw5HHQFnvdQqL2LpPgEzo7u1Awl
pz35Tddl1fjgEl8Znebi/tBoTrkyKJ10ErIka6fZpBmMy3Asaga1sFFPIdawFdZI
wYvIq8Q2qif1nlCBF9hmNB9UYIxChQe/2mAkajc6VXdtjbQElMmc/Rml1kvNFZ7q
/SMVZvwjVWo1P6weVO2V/w2TeO14IdQSCYFcSbBzEiFmcoQCzLpqZIF7WABrO3R0
tgE19kH0RzSE9GEpuJtIZK5Ohk1bMNGBCNyzk1LmnAOwsHENWQpD9+uaeObp3eIE
G1wEcM8QSWSnk5MOKY1mq4PoKw7X0xjcGNpGOJo2S+5g7hiAcuPsBAw6Wl94cxmZ
YbrT1c4P/FBVkNNi5CRs6ivCn7i5DJcm55GojIY2ABet0oDrFvwQCQ11PaaN8Xxx
x+EH2DyKhWdEy3GIy+GB5u4v9x2bxbejVNn9+Qs56ud6YWUUJXL+Lx+efuNv6k4D
dEJCK2Fimwu5TEia0eRQs9OGu1Aqjbh4IvQrd778csqHrV0o204G/PRCf3YL71lD
u9911S9bGivSm0szfQQj3oHi8aYAxtfQxemzR5UrZOxsYRpPachYj5cY7SB2fLXy
0XCPDZX05ayH9+Qzi1OBsU0G9FjUbgmjhbXwonK8UpAIqu16uRsc7NZR+0ZHG/xm
0NdR7EMfuMR5WWhqsgttKbB1BDr7tIWNxDjlVZuFOV1PoJEOdJeE4Hg45zICKp5Q
g4vL4bTaZg62ji71D88J4dtf/y/5WlChJMse1VqN/7CWw13gQVnf5pq4y82+ur0J
l+9mnOMUelX8Dj1jyCcmaNIMRY9lDuBuUd1o9fcApmDK/VHnos2vbjlxJlPWvw5I
skATS2ja/FYjMevKixjMOgu9vqQ1OujZemtZKOa1q/+eKlhtWlMfA5JECwqkJj94
yun8uQhl1EAIqYf2casXoWo6JpGT0HnHxL0w+GHhFj7iQhZYegPSDapLK0vvDHuo
4RD2+tLoVISw6E3qX+GcrTG38AFE5maNeFneOvzF8eteDTgxwKzcKgqDjWyiutX5
VBhVZLgImk5XT9wWxiUqMVa/W8UNfzCbxwhhAVhqsw6cJLLJmXrWzunQtt1bbUwU
7u11NurgCbTlNkmcpw5U2TIf6n8/W0ut4WStjGEoIVUZ3kfqZHVhW+y3LK2qm754
yyl8rXKqLFBJDUUWkcj5G3rPZxXfbJS5JsoYA9frcr6mh/nq87RXplcV2XSmx/OV
hFZa3hY8w11RvVj9TNYAPCzD4vMpS6e8B1xurzz1R66sY428hjkO65FohoC8wmhp
RdFnoF2eyRMrRU4l5V2UIfST3MTufq6wRiyMTQY5GeC1f3laN9Eg1WXR3Fv2nirF
KlSOdGXh45MJpbal8PgAtda23LQtpTJm0iyUOGGm2cHBhtZEbS1qADUjqhjqoQyN
kE3sGEFSQNHqV3kcqMQvcThB2YixeOqdehiafhcbjUvzOyVLbPpZlEQ831tmf6VJ
5dknPaBHY3/eCrnZ4t4aF+9TneF+mggnwO8VliYWMAQFs38DWjbMIkmNofOV9RnT
soejYSz/qS4SA73/l35qxYNj0ZrSizsRDktzRbBHwORkhnivJjYRD24JJR1LjndY
t3vParjoApMcCiA7OwIA5d/fUuVy28zerDGc+qJfumXzglPOIX2n0DAbpXlXbMcY
4qvIAuzo3mY30xDSGMfgt7cfguZHoBfoLwN9c8kHc6M4AcK/NyuWKimqAEdd8lBC
uZG9CjyTSiR2BDclk2Y68pk8+g90TSwXKCbMN9rMsfi96XkkD06iEgMETVzChO9Q
zfy2JVZbvnd/Mzm7U0THEEkD7Yow4b+HdoS+WJtYR8w24UBtyBVqvmecy+u2E4A1
ljsoWbIe7qYAf+a54oyqVxQfZGmM1cDUhHp3x31K8bcis6KjeYdyYRIJJ8ufnm/b
p9dZy3VcSgyebLhArZv5ibvw1DT7UdP0bdg+/ofiWrkSRQnguubg8RKLH6p7/zxy
6zWZvwXTKg1i93quS1tIJLfhWj053Qj5WzydnTQWn5qTOm5HsHlEpMErKx4qN81a
mp/7fxhhzE1kCbUCrUlmWVJ/7ju5cNZCPNptqZ/5uE9aUkWGyN/tViyHRzP9AVKE
ux8XaqP5aFIT2DN+LpCD5x38EL0E7rvk6nWEwmlk2qeGoZuESiLt0zUfblMB3e0d
c9QY/IZlgPseu19y1/HHopKkWotOnxeCday6OKL3ICiLeEihVDIWUHDXu7kUwBt+
A4HhUOvOO+zZbdwOkk3rwj3vvg40dWHBCaoedCLbrDp9FR21PmNXOKuVZy55dcUF
dbIBZ+9Mu5TzyeEtLahW1OfidArBUSrDvNtDIMEgMdh8WLyCZ/k9aDYX3rfvgITf
yZMdTpOcvhKzjqwrcmGbTAjJfAHPUlEWFNMqQnRxc1SvgjSniDNzjoKv729vIf29
z/jhZ+hO4u4LXfbSiYlwkf9bWTVZVBzoryRmTFjCc6HQGDdTO2tH3JrxFb+2/dXk
gS7x8yKuV19AdoRhsIPGKuS6i3VpITbbDlT8MUKXM6eJgkmWrtmOkfSBiDXUwBG2
PBtGVGFYmSBvVPUpQcbuw2DoOYkWf99lJAMrPp1PgcR/0hSuDjCRdwS2YuqGoYGa
jdmFW1OyzIlqAqaqt1hvhtvqQefdv3IYgJt7u+ooH+htOxjbMjEeBReb5yd1wwFH
mXIdKSbBmnCwlussmB2dMBhlxXlHhGCAvO7To3q4QYCs7ASUJebIe1pIjId7mySc
KnGtYVN3SAsN/Ct44vL2RZYIKZE5eJpLEZUPMtam/DwMTdl9vEaJUdPcsjgI8hX6
UjUahfKtRwz2CfHptEVDKWQDAhTNm5Za0QAUluGiElJ5A6vxgWQDvSZThasgebZA
DJMVHlodGnO8T8A+Z76ZmucbqTa6CtInJmmgxOj7awWZ5FGr4atsu+RlQ7bTYUno
0dcg1Jp4Ki1t5e1FqEnz+nubN5mQzuvrijIH1iGt2iKVVh5WVM7wOoY9iMhksMAr
uf8uB9YZmX92EzXbbbnq/hVH+5Ke0qjbf9Ld4xhwtifMxufmj4MD9bVa2oyOjDv8
8Qren9CWIFwTHUti+MTN7oK5kHXiTj6/3JT5er5KbRCeqegnsPZbRDBhOlZ+h/1H
7DD8i8fF/G5aVo8KlniqiR1JeZ5pyazzzysI+aiTuLt9ny2N0hFw1ISigIHxxjYw
QjakiPEkYeH1nj1woz77Qbd51l6z9I9p8nMguO22/Nts8Rafmng/UJGyPmBZ0iHo
KLrCSfhy54PMdoMNIc1ZbEwE80G6eFgBXViACcUj/Z81bFndxN66ItCXyK3KahKb
brSaG/rxfZSCMa47o24fvJoEXNju+bU8cXPfpSpeEmKTAf+PT0mePL133n3dinpB
9P04QXTrjgXYPwmz+XIOsc2hOP5dWf/T3k87ZsEsa52Lt5pMRk6zbrzhmzcONhdl
ZyixUbVF6lFFXYvnMeqJvGyycT3gAV2/3PvDeb1ur5LgtO3wvAqhspRz2NsbyqVF
YChYwJu/J3XfT3CjToZ76tBKz3TVglQi8pFT+B2n0EQuaIFZ+dJWDhlwNiWd6dNp
EKE52QkAyCKWfsvIwTVcDm1Qj0JfqLN127mo4K4g7BRrJBrDaFFXKFUKlk+T2Z8m
bHBx0FfQufKSgJgSwc2d30GPkrIWHn8qtArxguRDprptjY4/IAkMTxWPLfPE5B1s
2yPanbmbuFWZyr5xmJP5chKG9q8IQAeTSavKNrqGZsScwo6Hw/ewXWJYO1By57EJ
9D7n29vTWqZflkzYCY/c3oLGnwKI/Cds9mWHLYqlvwO5eI19Dz1AB5ERiIITsviW
UGV6kuyg28wAwwZJATaE4geCHjqsZyuFxcYijZWLDtZHlqMRbVsFTQJvR0J2MKLy
U/6JqVfhFzum44x+TtNLCibp9Im5ZxUp2eGU6nDjjxjR3QTM9NcgGOrSpFWrp1Iv
jW89JpJ8djBcniTtHBNd4rRHy1n8XOLgcKt5DCXO5eUuLz+77koYoXk6p1iyuNla
QxmqsY2b9uRqbEIopEHaXaj2/wHxKz0aZYNGDzJ8m18c50QGuZlRNaUGlMlP21tN
UboTfNAfqBxJaUkVtJZoOVk54LB5GzuEgRTvXADUjGwBnXC/DL6zPmUr3qHRJgvz
Q8re8rRlJftEqoHUdDPjtZo+ONfQtbRNNfc+XYl28CzbD7eBT5Rh3viWGnAVhuzj
H8gRucGu/MafbEnRDNynygjkCRZldE9HzvI4Vt+O54L25siaUkwFy/yEGqtyquNS
fHT4GVUhCGrRHEiHQD8oURCpCbpO3WAieahtSzTLDVPO5p0rQE/CGp2RJ9F6ncMZ
7lGSat9ybneQhTw3YiJ2AdE2o3ggxzlNV9xUsL1yn0nnSXgTbsphKwap6fn8jlRl
Nvs8EPsrI1E5dAq4y1FW4cGBs2yPTDUDjHjXP9e51gDoXqdIEaVjua6EXWc00lv6
O26J3B2rKqtqFW1U6Bve2kixQkJ74Z9Pwqk+DF/WS6pdwQuaObRbQjKNOzEgpKze
74zffiUzH2so4Rf53QcoOgoAJieu3p/m6j/PmI/k2XSKhR92hf3xLBvJKcvIzK1L
LyKwsv7a2k6baoIS2xENtBjDuCpyImeJTlbPq//94nuQ5+HWGI5z+tcy/OBuuEGT
BKYer54B5MVIAuGGGv/6Xk7desajMUhyN2qWY1/L4/Ul/g5RGIhI+LJ0VK1uOXPu
jZwT4lJi6U7AXQBc9sGsqh1cKa/pyqlWUfOY8zUZSKryEPAPs/8eALzUBqqQEwc3
jnBh5udohIMer2Q3IYjQHk9Fp7XzLjrf+YO/1klSH4goOzztnp8CSUyUvEC3M32l
VtiJdwWvJx7ywB7xcu0pp+Xx1T208q2FNH2Q0qjGlQp6LhsxdG8gTd6D7xGwNb1W
FcLuaq0yTH4RnWIDlp4QIHnrps5tEao40W56EfS5BHuVUeQ/FHA9mpYo2tHN1oqa
Rvss1Ea7S+X9A5XAL4gX+RdbQqsQ0CIlk85xHK/4sXHBJG2fFDHWubHETQjoiAEK
Pxsdq4/f/eB7ZhS3G5BzQf7y7GOgvGmILT+W1AvSVL2CHckW7NZnAkOCqjIF6Z5/
q7aP1OrWUoIbNzz0flp1K1fN4jxyybTZlbeAr2+ZZciAtXVolBogDm+Y83EdKZOB
9j443Pr3QiCiPvzUC7PobNXhJZtqVKNFA1MaB0cAwG2qyuBtkWiIJKyte4um1ilm
XnX4N55myJTsDLhgiozNwgvBje/9HZVhyQqyIVeeNF9iHDvBrWre+xaDiwcEAOm4
69yTaJt2WlvmjgYOHBYjY9mEtOKFBUmEnDJlde8T4Gwkzajad+fkSFUQ+h8JyeVj
44HpWTQl1R4fvgik0B3YOuNuie4cs6DAEh/VG35B9Tdq7UDoCpXMYKfdI/C6h0pG
0UlswgWQ5sc2qvqwtTCujf3rApakS8cj2ZdS+mkQNf6KCu8BjgN5owLrbfacRFa1
I0SqbVkRh2yH51VVBZKZeqfL11kUOApjBglvok/5SpRA5qZn19B2DuQdTiMXvVKH
QFVkTb7boIVKWgqlrQOB9XcAyLYVxqQJImg6c2WIFV6NmyOcT6QlqOOBCtuPrL8G
8hR59jHosiB/Viup9cUqyd7R2n1Q9FW5O0Jl4DO/8LedCXQLkUaczFvDefE4PAtr
DKJ62ZwvIPCjuWIvklSVPferx40lJvHVvgdOxKq6BtN5fYV3SgVRzmpuDjipfkvl
BetLKJe1FuQJYB6rwFYVCWc9jVn0/1w6eRdpilvRcmVnV/+hdtSuHAk1UP0TFcYd
qVjP2H2lj/dufdu2mcXdWz853QSgUux4P/zim+JYDJZ3brqeUx+d90VZBBPAJm17
jwCRDNLNK6nmaQL7D3iEdBf0eFmDapoKh/V1WQNVWY+hXx5fSCmIywwU3gvgMM17
SB1VIIZZXRCh8r7WVM6MXkvnjgdn6H3Qf24VdrvrmR6WU9vYYyZP74S4xiPlL5V1
GI2pxSridldsgGCtpmIU1kWLyfXXEyh8y9c2/HxXZ7UOUPcsImjWRh766kv0kB/b
x/NLuJeTae+48xsqXQEruH4jxzswlBhn0+2YIwASj0CPt88vqZ/HDjBp8wD6to/6
Uv4Pp1gbL2E1oHxadgbDV0RNy+XjvYrr+U1ltpNcGGgrmY3/9k8ZP28EiGGuGzZl
oU+fSj+U8HGYY21Wx+B+DoCxF3uRxHGMH+TlwG19AowBBQiEQ9HzCXa83YodK/du
AMv+dAV9j9K22qFyJtVF7M45OVsxWzgXw0szm8Qwvg2ic/mDhLDUDxpST5x0hlBM
FdlR51BsDdrwvXhR8k7T1cC2eyCZN/rSzLPy0AmxbX3q6jg35yUk/+cHAdKFTqLI
rQFW4z/+ZDlUjmXITSBKLmZ4n/GtwTBfdZMAGmRa66Ogk5mv+yAvdIg+OWsv1BoF
V7+Ljd3Wn5boofQnaTDZx1LQAZ5GVP0IAM5It7QRRGdbxyVs1f63Bgo7P9ypZ2sD
7v+nf9aOnTZWFYO+riBHZfXnwGuhbUpEzkTCFk5JIx99r7ydsJueidSsf1UtaNE0
1mnd4e4OEeCHR6cpdEw/0v35q1ZnWFXFXSdBAWjC7hI51OL/jP9LQBtVfyyiGOgG
eTIAyt2oCd+QGCwRHHPpneUwQSfPc+LnfgskFPXcVeLYXq1ghJmLTbaKH+XMu+GL
wF61LMVmtPj/+4qWdqJeXqJvYXndr/YpGjfIeFNwNSqUrk9eq7l4DOx5lXQIPOg1
W2iL/T62sJTYgclHk1bCxKAKodF07Rsd6v52Mru3W0YRpPH1kqTN0SIp6LJtonIj
CxODEyNG7XMaayZdwYsqgIUgfMnQ7IC4Cg902ToIqKriaLgpfkHgJEhSGEBIEPak
bneJznNuNqFLVYW7vxMeCOwVgTMP2sVG/KSHNK/4jmze7SR9FdeqZShsf4ZZINkk
bgl1Hbz2dvAF43seXRWFAZ5JT2YbrpVzTsfRdx4B6iJJWdeAvpd9uZSBX7JOX55l
PrwKvn46UBAfMi6DN178c+1u1tIAY6kLGfGV8nNq5zPdqBgyPvWvZOLOSTH8zay5
E1aaSHG+2gWElLU9a5KA0Fr4CdaHMdnkah0w57m5fjcPhfIpvcIA77zZHY+lNo3i
2eS4PvQbqWorU1Yv3+DO8DrLWrPCxU+zFzg2rvfvE7WVP02uGOD2ckMb3kYgX/bv
Rz0+pwov3cOEyeYdnCIEl9iboC2r0DqxPvLRxHJdr5AdNPipTxzt/LJYRq0AHL3w
+FB4tcL7Ys8eE1zndT03RYptsuEPm/fcX681gk7MzAQm7h+egB07r5Ddt+rCMBV2
4RlJvY4ba31gaRdTRFD+qo6GeXkp/ki5AI3FDUI9vZNM5TAnxepMwappKEk1+2NH
FkZ9Fd/FoXDEazq0BRMnLR4iSC4EmSaUkapoC7shktgl+9nM8wWbI9/LHzzrjB5S
kT/ZIEHh3RwfPtUT2cVYWYjXQSgpY5qFEw9YDWmmXJAwRJWLJ7jyr6mN33MW4tzi
zRvnWs1gcqdBmYwdC8TUnBSx7QKh3DL+c5OoypTWE2Bmv14lZJdPszvKZnaSc8eC
zg4MqJOyfPDYRg1VHxMroZWmxY1tlJ4JunCTaghQJMx6MTg4HI+H2XlDA9oztKIr
ciXnM5V7NAQ2wLlZ+NFd/HAZOWUnA9WI+44f0CHYQsavtCBCKs7y58vi/zYjGwGB
YMmsRfXF+fgTaEAf7b1+/JeqBMY703amvD8Ths1FtzcUsxoHh8GGjt3fBCSiW1wq
lS9EPd+rmaKCsoENaLbbxCoUvpLZ2XreFa1AqVODzzK+jcK0p35tg8GeZsJ73n2C
/KAylQZCvX33L52vOhhmTMghuR8i7BDEqkqcrdcITyRQmEKEzYfkQevWUFlYmQOr
onp3ebX1X+hwRlswgyOmANpHfeKocUnDifVrVT4Pndn07BfNc9XKZFIxsVhJysKL
ZEmbLpBMFPKDyM/+p7zv9O9s8TVUdVQsEitVr3RG0wQu+chaxpyhUYjKfeTETJfJ
DPR8WkHB3GOSKiawZbY+20gWNIMpLxXzgqMGUfrysQeY4tJQJVijeoe5p9OPPVpo
Zu4e104LUDuG9oEkItVouu74UzP1AXg0E2u4DqEY/TORAwRanqDerLCLfI4q0DI0
dnKfasD0A1y6RZgmi57DKB/o7YFf6iewoNK/BfVybajfm5LmRLWz5pXn/R0FKQQO
IU5jpIRQZzn0BoTBp3u4mMAWAJsRyzoyOfza31h3ptP1nJcbyW4pwDOwlxb8P9xT
ZWGlTAZecIPxKBiBv19bQBanYWN0a3L2Y1k9JGHgoOrLl62YiAU56J7VpXUXar28
ZvtdMC/EYBbRFsjGSvoIwC1fRprpJrd0k5KaCQTdvTNPr8jI80xHPknZdSXb/7/z
28a7ct64N39yFRLxRL3e6dWN1LIqV6jeqKuid55+a4IyQZVd5ZaMlQ1KgL2NV8Nw
hTumQyE2GGvrQO3iNxDiBpqOcgYgh62++09ZrkcKpBueckMgY4K8bOWg0LCk7IvH
cxKt8TCsa/IKvYlpWX+Jom6rXBIzcnkwhfXcnKRZPXp8ZUew274u7gAdPthmBEBc
m1q6YjczyzkBf13r+NA2GPwACSIb9RwC+scPa06xIvspVW9Oi7BIOy7/kkL+kECO
+EtczCKTnlzOnxddr4HH1o3N87fK8uu/U0ZyUfIn7932mh7W6pHMINTBikjT5jtp
FKwFZk8a0AvlcAX2Wu+G4oroOJoZ86WU/PKnf9Eex6iCkWMFP27qhCcLwbG3tPsr
BpnG64hKzpVwU2VlztnIz0C74cOJzY0cdXLsav5w2d78BD1dwk2Mi9SaYBn6MVHk
R5OpKuO+LXDZ5OIbGsMoewVohCSJKZuqN83Sqh0KTnDizUbyob9EjYILVqIGV8YW
4T2zwkmiIyN9IupJLBEFWsepvzRKYTwgjnN4nIOgLH6FTvV0NMwY6v5kqPwv5uZE
j4xIgtzCKk0rYU6tYloXCfZDrD5q7IcMMyk+ROLgzjNmt4i0MMzixEvUrPg7gz3v
2p106w5mKu08noEONp72XirQTYQuLhJH2hGFCE3j7OWHmJP4rX527He2fwDPETZY
D0Px0+pVE4g0t8JGxJhXOkrzkNJ7O2HJCp/StvaO34upvt7BuwpmqtzhYSPaMUDx
rqx73BouVV3lpvjbE5i97hF19xoLo30MSd+yLk5wPn3AVwSvJ/vSIfyX71PohV4l
HreJJKQX4nl1gaot4n/YbgBVg9hLThaqg2gutbelmhk4I3Wo9fYPnqBQBsmAbK1d
ohOmTQGTm0Bue6fsfxgTu6SBadAoFUgALJkzyYmSy55dQpUCfcXpGY1vyuWn+EEQ
tpRSG9idVB6aeKDufbuKNqdM742wIfjYN7VrT1AcMAEUTKXwATCIGYzaMr4hRFZw
q4L0amiv39ZXkhK0AHpsXLnnJVb3S1uY+eJzn1RFcNhVZRYKcwGvG/Bp8rhGpIbi
pPD2rZceRC3GwNTwWve/U1/J9sHK6CgWiIF9hhQapgVfhVl2HOcNyzwBnSY6Uthq
X3OBGcfZsBtfSTFXDQQI/bgiiqIE109B5mF76DzMG2WhBsGJmmKAKAxMMjdIdoqI
lcaLBXnu6Ekw2rOrWukCrJcea0ThP94GjPle33aZYmHVgSb2VQQlXu36PNfuu2cq
w0KQAi7FNHiGoPt92wq2BGuksajCW7I0K7cRoynN5l8fwajBVP2O7E0CGg2V1Qoy
Yu/frwkCie76z8tySGMpe9dTIMZD0cF9MgCOuY6SiyI0gfc1awWyDTHmZz9OhCAu
lq0twtfOT4Q4DgTL1+avG+fHimM4QwoBSQ4uxPNb0cW1J93iRABDawgqVcbk4s8D
AwNwX2mLkN8cMB8zbcg8JArjyxfU4IISipMpmgrF5IOqJmqcPRbZDsz4q1aPoBMr
Z8sgQpD8ZsaU+LELOXIeGOx9gdpelzaU+Kejoqs4Y9O5/w1KP2zK+dT+N48+Cv3p
wbI0jbxYb+2zldBejoqT/HHhFbszq98YAGn3kE6fl14iTxVZJrpW/w1jj9rKL96E
OZL+Kv4vvVm9Jtj4MWHROeuv/7zoYEwM0UbzjDHM2Y78VgH69fhhGj4fMtPMyRyJ
hZ2j1/mLXMgRG+94EwpNuv8AsOuJfnjm+Jo/rJg82+fcK7Vq7jYnxdtu5aowRJpf
NNrHZthSscxVpo3fTqZdcAr4Sfoh1fb/1iEokbJ5DRVEhE73/S8dct30vVIXtsTQ
273OxKA47+a6khdDR9lQfgE8mVZPlMbTsRmttl6XreAYNvKF+hST/cbRTtbLRwv+
puA0SFO9y6yMWr+EearMUG7Ar2rSazB69tFWoMIZ6Gu4kaAmvAjgQPP0JnEFtfX+
yA0zeS+CVfAhx17tJBG1k5cbrThT66piNqyBa7YIT+D2BmT/S8L6IB4JSj08kQSL
zmucoiX4hnFaYMn1Fz+jrI0HB2hV16LE7VRFuiE5yZBp978JOWK8cDbalHuSnPUY
saje/iOcaoGXRUpt4agRmzCMDg+e7vNnmZxFTm6Me5vyiMPovelDICx9tyAzC/w/
G6h5ZENR2HShdlhKCK3RmBbjmzL2GWRujpFrQlDRa4GuPD6IkjHSoZHwkymkQdgz
amJZFTDfSliTduCchqAy8uZuWYlGwqNHK4H0TZxYAfoGf7DBx/2bxbTB7U2DRPJr
Se9pOvOfjq3OrP7UkdYH/ZmcWV1utPesWPkR9e7hKN3dgULdjfRAOs9FheQyu6P3
C8fDWhvtymvJ/R2mLmZeBBoC2QlVNwMFCT27wMvNOBlZPvEvttA0KIjFE0TP0T51
pwOE/JJnC6pVyJyguZXySibfZg6pf9qirCaRYoU7oN8FPKNvuoNM/hRlTb6S026Y
lOh+cnwU37rr5edX0PyMVIPDqjr6EVxGDINpQpVZw8knmglFXn2mQmd4Q1VzX8kD
aIRcYqTzjmg2M/o3sGSyVDSBosJUPRVftAncxhKOTItXsxsZgjNjrpX71CgR6+D2
NlXN4wzIcVFEwVTPQX/rwPm1VhYB7UkxTI+hLMUVOHU3xeRI+hTgpUU0UQHtTS1S
qV52g0nbj98iQkDbxv69tHW229osJ3KnW7KwU2mVN+uTxM0fwmuVREO70EKq3jE9
2TRthZ6J9sik+bLPB+5Fn+MyZaheoyJgppEB7jo9YdhD1yKRBEWTo++xQWqIWYNV
eqtogKxakkHaTXIQJcLlfXLCrNBBPCKC8u8rxplVuBoHDklOuIhNKq49xR8H4Pci
r9vX6DO3lum06v2OvhR8yQ1b+uSXuGZqtVNOephZ5NXrHhLrOYKsmbKrZ6vJ6ACp
8xTMFD+dbFS42NydAgQSrU/u0oLALtYset1w3TNdGIDpI+s0fEeGPGYPbVl7Bj1F
zmH8d9178TVZ3wvkTG767ZVjFcOM7OW8RxvuJQcFPPxaSQDaLXoCF7kmT36kNCFt
3mA++WIEfmpXbaxi9G0up9vct66GvzkxqUyXKcEOTujTYUjbMmTGzwFngGQvRJJh
8X3QByVz09j4R2cYYtoPm31OE7iSNIh2sU9gKUN6RVf8gcJ+7+5ozqyRRSMiDsHs
HNivXPEz3W6xDB8ON4oxs9LFlCXxYPNp593K1ac6IcplnhssQBAfo4+z5RY9mv7S
Y4JsUk7DWC2KupF5phW98MvziNEGWEo62g8GRWGsE7wATwsW86x0wIBAtSm2n03i
U6QYV8fzJxXii9cEXDuEnn6cKNZMJ7sHs5dq6i0UMiNBMmIyYjpES4pmkKuf6ndT
H0TykfEnppomrwJqGdiibNiG/9SNqjtg2ynQJjVaW+CXPRKSDWO1vja9eiWIUZqU
phnmMIdWV/vg0LHakZ7wfQa4eeFp/18jE3jbj2ZS8JIY6RsLWLCvvOHd1loQHtn0
I1g0hiRJgpw5mzRkEA/eT0WERUxNtAK9/1TcwDk8//0zz32Wllp5NZBVzBeY0PnU
R7OGgZPBj2vkwzYyzwCdfKkneI2ZXnIZb5/d9jWGSb/+H10MgRh5MJXMC/njVn4h
ZQWrDtPFz2ZPKwEulcBX7F+JCHpj8X0znJLi+ImJJ+NVyskCltypZCH9VKPBNZYF
Q1fuOP+b6TlOxvfLmgjw7BtrJ+nhEKaICrS4zYRLVztIbu3A4YZTg1lvAqO0oell
5VMx0eh+x61ZMw0IaBY54UlBuh9HbiF1bDwf89huIRMJY5cLZvSDKjEHd8ctaE1Z
GMxt1T0xG6VpuzDH5e6/oaO/UxPrGSljVBKF/idGdn2wHzT01FldCmxOrRhjk9/d
akvNdZqOW7ddZiG0MXm6DmzqOZgBZi/J512oFVtmYD9FNE7lkskLv+IWPQu4Mj7b
M0rtxfVvO2kMqPRlP5MrIkbArbX+EULCj7jU5rkTZg7Ko5oSZDep6Ea3FJ7Nw53x
IBmvL3bCsY011/mD7Z2J/sWrXWA11cDb43vzR0vMhLFNK/vSHBlkQICIbCurna4e
Y/fFhtUdux37TH4ql6OyXUYOnQabTn3t/6WymnudP1UpjqEvYUKGxTsbYpTpBVKK
h8vgpsHTvtywKwkQisQHXLHislHgli5I5JtRun9FlPu6xVHiLhOTQUw75lPs7BOs
WVqXkxkL4d3VAlp+d4+WC2YojPDiAeBnqiU9froU9aKd1+DLzkcDFeJY8Y1SLBJJ
5SkUnkm+kkWbLt4Aftt45SyuFA5mViTpa++CBHJYf2w+Zqgj1R9787x5+q8nT2+V
mGkVObZSAJfDQtCWP9kpNEDaXpVqeueqGRldHUUyj/0V/+N6giMGDHxKQIs2A+fg
yB4ZgwkAQ4HMWO0U9UYLVlbrNwUVhY6r4WcvYvVAT+VIRfA20zbj9OZv4PCYszYJ
Sz2V7PuV4IX+//WkSjOyejvEg439A29ydcic/uR1vp48vdpXkNQaaIuuGjfLFyqm
p75ulYSLS8J6P4YiCpHdMq2z6he3Ig3wa0/GyLW3HbzE3TzJd1ScF0OKWCFTPbZw
vJcZzxTwZ/tnSEJNgOyLuEpJtdiquCSxfCZlbhkm5qDuVaNJ69lAsvtTS7BHluPB
03CdChlYItuQErMm48qp/bajocmEpHzg70xeCpk9rZ+8wstVwtwAxhlxkgpPyFxK
+nMVrFq5iNpw85bK/gxRQEabiIdvJYjUe8bUMQ+CDvgaED+zm+t3ZuFhNAbGJK6g
4/jija/5fYs8Ic1Xr6K/Aw5CvTyrbiNYPv+DcrGGUtZ4EcsT0r5HI6ln79rcAIQf
ytk5v/z48MxZGqJK04aWlzroZlvl4ZohczHjMgiiTEXWWGEY/MlyL6uKhlS7IGxU
Cd48DRF3qzKye5eNSULy/elWx4PWyWow3tmqqScWlz1hljlMDsnAtcM2YQh9R8o2
N8GwUWfpEtE42JnMDibUYk7tnLkS825fgctCnsrsSsOLng89gL6VR6FkeNVeooEr
KFEi5ZyjsxQWpA0aLsswuq1IKWD+SoiRyQPOAM/o10NMFEBi5N6xqTrZzAfuX0Pj
Ah9JogJ92hNCSUngULL/dJF7whond4tyxEV5caAPUZajXyedJmY1+BNNztu3VQYS
zwwShFsmzIgpHrMpSzEwJdme322LYU4SEEHfKQ0eOLsm9vMM+D3uHfifnglQlRo8
OIRuX9OHN1ZFp4AwJEieJR8HDPEdmD8sBsMbmlbJ7WtMFYriwODRr9JAd982OVs9
sjdSyc6+qTozyrVlCM14G/ikwAxih37gwNZeFi5HQ6MRptouxwcqIIH1I0oogOBx
mui7S0bizw/Mndm8s9oO3aCPC0NhXkKyGw61+BY18EVjNHTBLcX/ZkiBZ5cIZOt9
JxYEba+8rzvmxodaj7beXvedQc+fzFxWzfUU7XsYR+k2MS7FeaYxO/YpTx2nDZPj
HwuHu1OdB6GY8qyP9Q8n0aGcDY+HZh6zOEK6WGjZHYs4bzB3KKBH8km4QevRwfHA
6y2l93eS6emn0HdmDuZ7LAUBqr1mVlawUKgAIzQgsD0NGMBoQ1cYdWMDZWaFF7lf
8rhRQfer0JL+JxVj8UewxRi53TlhRL/DN1cgkcjQqP7hCyt0RSg/28OU/46CNyL0
9qe2iTmhMrEtM2Kup994ZQy1Vt7yxDcSfk2go0pbS0vP/OibiqIhSEIZISda0ajV
G4Yy9x3GQ3vnVPo18tcbSeD4jkpV85AVzdcWSALOTfYwJnprBDqtr/gCu0TKG7zp
1ikA2ayJl4M72sIXVusuCg9K53F9uHDQzONkAlhD0PwkSTior8xtTx5zqlDQ+88A
6x07SApMpij4/PHM5JO/gJeVISPDnEH79xFPvL+29CTLes6PnVrMduD8f9CJ0vMy
XvNfZM/FxOl89VDKwA63GpSXnzBDdaH29WkiIcXfnQZgaeC0sL5WbRUo57ttKSi0
ooj62gs/5FZ153E+Cgb3xRmKPgzhxp6sUjH8LgBqvv7yqEG7ErIM6JWYGxKC0ELR
oobm6mzlSaJj4V8wxd3OKhmWQYkTBTf7HLJJidUwCWKQnwZ/1IqtTM/nJB96Lvbk
zSXgasK4ST4wJ6s9AAtsfKbOLGmTNtsO+FCYe/OKrULj+VBEYLteCkQlDh4ScOiQ
aZisj2KG28cVhMm2JNWmjXS8Q4qvS0dfX/OrULQuOyPe82nrd6TfLs7SkysQmBw1
KIDWZQGWJf8DRbScAtxn7xetC0ahAUAYq3gPzTq0tCrbBoZqw8yVmwXptx+3YFkc
U+fCy5yWYmUNBBjinTSKcGmlUcyVs3JUruMfFR/ky3UGDHcR2+hEIceew4WC5GPX
EQsPMBWUZkfbJxnPOvbPK6SFBwWqF9jX0rqYt8iwFJ+ijIfjbamSdVKXxW+DgcTm
18urNbMrENP7iQGKU5BeF+YwxtnDIYgR8U+/lmWbK2hXuwaAvt+foepW2SzKm244
Vj9rskz422+PfZr5wWQCZKB7XChBm6TlUMv/G5/DUxsJUkg7R2ClwoiatF5rCMje
G3tsApwAwY3Z/sCLPiFJqI8iFFSEsbSnkdf8Au+nNl6rh1AHbkmCCqi2Uy7w4jTV
W5rGsfDsxcxX4tKRyoHMyvpA9sP7z1KNh+T4odPoSopBRm/GbJKf7DjYN/DLOQVP
NJ2/KVpmbnpt94FNBfxHNnhbPd2TrP/DLNRiWJtvRDH50N2fxn4MwR/iiAQkfri0
GP4QjCIebI1wvuu461Fn66dBUblDKzoVR/i0p75edZl4NE6EpNj2jn72AwBX/XE2
wC1PmF7diVaLcHnGJwcRWyqwqqgqiXhbbGNHsTMv3PWYNIxsfrAHuR835ogNhFic
XgDdDt7ktXYd1c5JgrXGiT7jLGjhVmZNxiFd6QtKmcSLuacURkigA39hiHtZrKhe
+bynNjGKPd9to+DXqVLCUNEmIH1b4FigDYAsu/P5Wo2ual3D8k+eGot4yr3zddrd
j7Y8LG73rKRUoFFYWd9aQpFL+MXQ6XG12k9LJFa2P6/VNLgpxUC2iu3xt/3zpL4+
vPcz4g5BVwJY8p+71Xwkz1y9u53GVUkha/TWkkLraFQ/YjbV98O6lvtbNIaKAYVp
VAzNeX85ipIGfrsPzMXoS5klqSsjZVQJ4Seto1ezhmwKMOLtOvkhTW1uyDqybOjb
x0cdpOD2tSdxImXJ09LXssL8tVegrCD/c/q6Kh+bwq4JvzPj+VLRZX+JmloiiZCA
c/u1ogshpjQFX4zo78vv4tHEUrkd6k0wMJl49WujdGG7/dq6k0KL1WMxqP0xnwaz
Z2OL5Xbmf8GL4JPGOk0Cn2bqmwjZmKVC4xuzRMC23w8XBjbqWPntJiQKilK3vQoq
w9czjKgpVCDquyJcTda9ol82CzBNApYfgMorPD1DCg0pmexPdp+rmXg+f/uWvL08
rpURuwSOX7O0rOm9MxTWJP5axX6CSRQ1xMdDpigCjyxIqL12pPCI4O4nzQlXJ/x6
5psn2qxy6KLTp5gG9FcA8bklUqx0ZHxQ/hvJdILVoFtE2/a7Lzi9d0Zd+vl3A2rk
xrooIZwIYRE47k9F+m3cB700FB5aCwOseUNQ7jPX3SyitHqOIAkPgCUMTGX00Lg5
T8rCVbFIdGXRQqqHiZ+a9tiUT4Sl0rlEBoxaaTpK2AN1Es3AJPmEdOvCodkfgEab
y94BJZfRAtRCNdF3Ze6jH6ZT1mLRTRGynEmw1ula5u7wClqt3WUVGPj1T/RNd+Na
Lb4Ba4gQnQZrzmvlkCXgScCsaj7NwLwdiplcb9jZR3IbY4AmX4TrTwG1TvomZtmv
5cT5luA65LtNWZF3BmHHNzB5Mr+DG+vO7x9Xg/hPlOiIb69+33ghVQWbvQzKUWv0
6YE7HLdIjbajz8eNZlNbqA4im3QBS3Q/xwMW7vrRCX8xmV18xH7czqjUzAZE4sSS
Ntdo2aaKWOfHKcvkOUjDWpNltSAExnk/LaAcs8w0NTwLKGivFB+zo6oiVcoJznZC
WYhZATHWLyPo8KpUGPIqGzpkDH5KRPbsCUgHkdr3iNL/HMgii9rI40UwvB81H1mr
RdJG1wM+7zkQnG4j+BNHT1yCkISYKh9XEEqUCy1llflTJbeT0vPbdNfkVcXB/oRm
43uJNTXM0oXeWEpsfwuw85LWK73MoQQLuk5E7NcJp14fuaSJS0XBQFy3Cx2bZIrR
d+mBnDT4nD6n5xhtNyaCr69VAWZJphr+yCGbEMnhZ+N/RUjlzuZ30VV0zkbp0Ysr
k2n9kFwanRSXrGnJUpvqYVPrkM8o+/yZ3P0UnjO59FQd/WMsY9prMFCHXOvMph1M
D933tZlGShwwES1mqTdflhZGb9r3IuQWvTCKkdCdUShJ/GUX+IDilZ7PwcqDg8m+
7sRUEtGx6QzLOtwhPj4d7Iz90Jv80c9DC68KVHGe9RnfV6Xs6oozVHA1waBx12vE
YbjuwAM3U95EF/4bAQqzm/v181KWB/fVyvNoc9hLstsEux2LagSAIZaU73lcj+0D
/g/vK2dkrj+eXWmG7EKGKzD0JlgiO2+6uo7MNriX6m8/jKWZTXeMgx0dn2TS6ZfE
9hpw0qRONtDCrwcCFUzP/xzfe5Ku/zS3M27MjmTfXtCAeOYQWAnDnrhumrIe/322
mwy/xIiqmpZ2Arb6TdCMyB0Z5zMsvj+59i109qmr7/B+0LelzVm/l2ANKCur6zWS
jIY7MBCUUptEgrDyJAdhKmiHDTyjnV2gKBaEGUxeFI+7rV36DDpJrEy+zB+ZL5mf
G4YHJHXzXpnFOfy0LlTtKK8pMF2vG00zrgtsJRIT2EYFjOCv8nhd9YL7rRJaNs38
TA8KbpG8Pf7EFUAs2F242SiVU6BtNjXpTuGEvkceDSI5SD28xKEtNlrARdJiaadC
oAoDIuDGVYPS976SGBCUluApmnkgGsZqxaOw067s7V0cMfYBB1pxX1h7H1anuvZE
XrWjur1NH1l02frDi5LidudSiLEEKc5X5N1GSqR4ewA8iPl9FdBOMI1X0R3EfYQP
ziZlCcqneJl/DKcCLVDcUNjXghbq1AikeYFO8ktkWHMoWfRAj1SnG2A2C3GJVD2H
W6IVSB7OtQ9ErTfvbu2QUJqh4c/OhufzuHvk38QIK9gE0EF4D4VyA7G0fjNaCNXw
d4ba9jgiC93r+6WuZka06fqcOcwrTkThie6yHLc04OGw3pgbKRHmMZVl1NvATZO6
J4jE/zPqV3PCSC+vqGlKQvIg/lv27N0Q9mk/TymVYUHMn4AxXY/QeKgCSDNipegR
o6n3hgXzDqtBe5WOvV9Q0No7OsTx7VcK1JVAkFDqTCad8xM06vrn92cngJIIaTn/
CnzrX4aGt1ltDWdRNpvHMguJckBP6ME32vKAzEwc85nT9HVo97VaPWCQmM53mvpB
LzXKpRXWNPV+tknvY1gQJcvwgzZ4dNjd0RWV0f4oAi/KMVlHlsCJEgH0Uwxt3V5T
uiTe8ExTYdbTZxTs5sjK/gSsnsHAfRbW1O2wsRqw59045taY9MPWS8QkpmMg3q+0
sjm91V8EYRlMiuJAhemK1ytZulidIbfT05arUe9kqCtFXCyjfjzTDurKbLhKsG0l
Rc0PaTeYML6gCYwE2Yj4xW4MH8Ps9LYd6k42EU/wy6mu4bTY2PnZs5eblUjy7FMy
nTrsGcawfE7apPJDFiKZrjOkzzDTKaJc1F5F6W//nxyYQsWK/4POT2ZBmtWDBE1m
FOzTvPYm59XouTUEufWGHXkV1Ov44RAKyez240NE3rXnQU2K5Ttj0Z+b5uJCyAhJ
2FHXbev42LET/yKeFWH7aByfuvW7U6CbFLMXOD64mkH9mVF/Py6ICdnNcgDXYjop
8fnkI4HoNDaYBTa32Dszg/V5kbCCRpSfHQ/fJig4J7cfq8o0KFXsWTjUlw/2imZB
1i6Thqome0nOkC1cLihumC7ZLXGQV94vDRDz5ug67iBeCYxk0xx1h3YBq0ahpdOZ
BVWEZiQUlrDmQJMZL8NbtpZWxEfjG14PLI78LcC3LWEx7cODseKJ/0k/15QJkI1H
/CO1R7TMAFxRjgTSnYuS3tcCeUVjTiMZxLXJ7AiYj3C7ENiJZUAt0yrSKZpschc1
DYk6ilQQuQ0SfptBee+XUShAqTZhqoYXU4fAMTSEIJjom8AGGraBLhOqIlEkaYcS
FlwLVWgCxHDlFP9SMvX8+BXtuiIcZeYjpgjpXVouK1Hcqt4CMetY0xQU3uZRV2KI
B/zpv4q+ftqiVWVD+YWqd/jZW5TSoijMpjZyu+yHJOVifp4Ef0hpg6vwx8dJMR7U
kGPyrT7SI5isJ0vwiPlJv5sltHCLTiSZm3lIvuG96anvOJCJMctemB545AUGvcBF
F7Z/A+b+vsJVHPVd17E6xEl+iHWL7DMH4I7r5SnjBiZSdlqZmlYe4eJ7aUWL+v92
y/slhrDl4eLGyXc2ruaicfyy1ph/Rd0QZZSKZkI/IAfHmEVYAuj/Jlk3IqdFqYZg
sSF3epCD5i+WQHf+vtE29GbFuR4R1jFHWusj2U3f1ZzoJQpWlkKrPrSFjohwsnOM
aVudBa1tPJpKWwqEiNxYWfNN/srDDEnxvP/h8MZtuagnN7W+5M0b8TehYaduFrbA
Wb0D1cAaEPG5kvWcsVSAT+VNuZwiX2H5P9jqOKBU6uM=

`pragma protect end_protected
