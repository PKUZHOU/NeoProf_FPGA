// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
dhBHdvdPIDYrr5KN2y4QA+3EZYhe66YAemGmrZAy+TCI/ccBuhgQWTAR6nja
To/sNVlrzAm4PIJHBQwEKJf+qgMrrlFBnxxvZTeWxvJ4c5vgrpU5u6YigrF7
UFrRRiFv0xDZYb6mSsmf/4quN/KcBvMJvUy1DwjoGiWQUWYNh5x0sbDKZV7E
ltlrnyaoPQta/z0GSSFwYpi98UCWkwpCHPZoR2EzxQFOUSB8+qBPm3f8qNu9
cxr6AbcLENMiqXhMpGN3ZJoKhoV+JMslNii8Fzc+OUqlWABjSD5vjZqNMqIz
IqZTL/8a5FXtfuktzeXSzlHZBd3plQEomBWlEtLViA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
GATdSn/6B5YNsAQq22uZG93WsF0jgwv7jkfvLvAcXq6ko2rf32EJqWEDkWQU
GQIzPe1TzwLl0ALqfCParbBB88CgW9USoePKSL/EngZtuU0V1QvO62Rn9x2B
ObbSunTNZsg8p4UniX+kggBoFaWruFs0dSXwDvG7fTTuhI+psGp04hL8XhG4
XxPf3iFXXc0CWWI7cQUx+hSjf1qRvvAGj/AcWlTP1oNYHRNI+FmQPgKiZ7vR
LJuClOidGtNmC+TRNFUmpwhK1CvoSyWiK9KaHHI9A81/6hhUcoLp3VKPbXmp
/kBjDNQCLb0KQHRMZJlaHDZY1U34q/ylLbtYMQwNwQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
aGrIpXWsfl/LWpVwHMueM17zgT2NnrEqlrGoB9UIsOcJaVF8iyhmLAKKfYli
Aw8C5QvS61rFWp5jZzrn1sRDTwlYuyznxgxuFe3/6rqvErhEgBByS8IFYx0a
pk+IL8vS/jj7ZmngrOZS3EwYG/lsYd1NjX+GBAx0RYcDkhN9+KnaSFGh2/W+
igBfHdxYyAg/buchlonBYwM0wANFHgpYIT5NxP6/Bc5jEm9wEAQm5+QXgj6O
raa0bPaNeZNG2qdfGDyrSSxxmBU8Hu+7QAuyZScj4iuNRvg0gm8YRMH+EFZU
YLifEDnc6lO9MSFBQNGBR/gOhtzrgNDkj7JKdE5ePw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
JMT1yB6AtKmyqeIDfRXTwe8Kxydtrfq3AyFj7nvetYKkHHGfOatN9TEh9w9U
s6K7ipwYJfCG9ChaMf3OlCHMCiSPzSYX6h3LkUTec/QenEvfl+w7XOI7kE5n
lhbH4QA/+6n7ldgPQEwJnlwuDf9SzoNMYqwyxxQknH9RKd/Hgks=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
e4p7+wc8aEgs7Xv4aynZ1SauGQqQeGkAc6biNUG9V1E825xWKcXAZHMt6cJ9
o+JYnEf5ZGjj3dZXv9pGvgs4DduLnFKdSmIYm0w11GgeHgUuyWUmbNh/3wqN
Sh4W0VHwtiacCE61OQWkLrcC7dSy3wclNMq4MLicSongFzVZSqfUPhERuuKf
q8vPozuFBaTGLrh+zLb2Tx9g7YsF6xCyGJVjuLFiuj8fHPKwsieNaCQsSDRZ
8YKvKfwE8T5TYHAsHJByqVUvcC2BCfXGOmgDAkUovrmvKd9FlNmnT/e9GqB7
aaQTntKOu1jBqye2VJn2O/IOk+phHgF/kA0czg/6LEVm3HM98ejb9Mt1OEU4
OeeJlwspkrjxsPIruIc18LFzLLnO3ambXMnk2IzIZv7zh1BDQsoYTNdCEyeY
m7QOSw9Ql7QbIBJS33Ip3CVm3XcWx7vhM9nCBY/c7iACjveDVEjOXtILyz1h
dT7lr8oXjdDZ+VN0/yAFNxrgb9uj8nM8


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
drgbP3DjrGDRYbKTS5W8H5eTNUXUBLCVxU6XdWY0n1VkeWVeYiFzjavrVUIx
KvvHhbNCKSH2l4JDyFY8RQyLcOIvVYTHZZnBT87haV6Cc4f01jdjb7DO/ypy
8uVQo3+XJfa+ObywKi76PMPrW2aS1XCfrZbltqPymLybrR/UIgE=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
UpHBsGBj2KLPBc3SYAOwrEUdCg1OKZQLM6EK5vETlMEK6ZA5Sn+IAPnhhjQY
fNKwJzvgKn5lvgNJnYWKJrWg1b1syDAdI1HbDoWlfdWFDOky7GOtyBfm2o2W
WBZ+ca975T/aypI5CAqCnF8IjfkbS4gXXw2AtpcyTMYf3h+a5MY=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 17440)
`pragma protect data_block
1ZpF/+isUayRUYksX7ASsVqCTRTjIE4WMm++XhgaMLBLZDWmG2wm+RFlhpdp
DnRnHcRK+ULqUCVg/uP7FcR0J3aoYCNutWI9nWJ5Qihc3Zz7WPxsy/ghLBQ/
l+HBw/iY/KKKFD5JFR8QIDYJiNa+w6yQQPCHT8NGWW3yyGNh+cG5qKYbK2QB
kVFsQC8MImHO1zcDuC2HG1emKgeRKLyr9xUmy1WlvMvkvRiNl3WyGq5WE8Dj
xYhGaBhUGbK83fQxbsiDAv8VqkzKvwhfWkSfJELt+qdoAdl1yjBtBkEneTS6
cTgJPWWT+wAMMJoHbOFFsZEf+qW+Kyy+b1Gb/5ppxvhuGN29ajhgUq5KkNwi
OtMYoehzCn13o6I2so0Ckusc0u9rGrBojJ0KnRv+3TCGT9UM+Gz51ZDRgUcI
9DkXnD4C9hWKV62Ox64qU26uSSxvBSY4/yLCBAJQ1WrpFXtlA+ZlSWT/qI3v
6EjmKZ4HyKnTU6X9ZM0VfFBj+g/dQNOuaQuwqGDuA6+vxE28BX52NE4gggcX
yUHRAMZJ+UQNhqxyNkPtJtbnQFEWrsRLNUldW1CgK28hmZjijFUeDdEZTwd0
8AH89XorREHO7kHCKbZg38RFhzB/5gY+776wR9/NxSXLOyVhdWsnqoEotn/0
/xsONivRXE7qowY6SU3TZ2io7sWb21iacrjlImnXiVWsoZuOS3HZF9LhLSB+
iE+l38E87/mkGPc9meb4TYJUzg4rUumNb37R77FOgRQh6pSexBTts75i39aV
IaoonMlT/0WrXaJbHjfSJV7Dr56G7mh6F8bDdgbb0YFKgv21W1GZWSffM4PV
8jjlfkqIDAmTVGxbZmWo20vWvLup9uFWSNTg2VzB+OqE7HdE7gKyOYLfo9Rx
qRi63xcl6m8wvwcz8uy6l++JD8deMQ8NG9k7uKzN0UBrR5Bsav7Oh5qFZcJ+
V8E/9NIrK1oynozawE4C/lWJ35R6auX3g2sL5f18UBnK0g1XL9fd4L53o24Q
jIxwXsYlfwPAtqpoePzjbVE+Hgyyu7Q+RxOWxmKvWx35OvWQVgXKpx3TZa4R
TeJZY453YOt9K/HfQMicIVXF72auD/7o7WnqbOfSZ7Tu7XQoiWppiRjj8s5D
Gtml5jz4bM/aQgWPvjlu/2XcmfncfGaZBBAvURUOTo3NVy8qJe4rB1Nf8yMq
1ullq0EX1bVGeJtSXSPy11FTRf/L+XvrZM+n4laUMNIVamnMZzwGjCApzFex
f+zqeUwa6zZRdR5+7DfxgrqWZ2wEpBQ+sDk8BdAwFh9Fs0dJmpPdUkh5K535
I2jidt5zVupQHZmnDWLjZdyjZ49voNDrm6IOVRg4ip7EnbcCF+WfeMyoOwCH
2vRP99n1bZyW1Y5OsvYkSZfgxsvfX4b43mFcy3FOr7koI7BFiHCtlnbBd6Hz
nyAPIZtsvl6WqR24t9sYwpDxwTGzYMSeo0agpAARNUv86kaNIRtyMyxLAEJa
WlyQ/wXzapVywjWL43XLIOyzrKyfZ2ba7A6akD6gZu5rKS3lFaKOjIE+y/b2
/bvgCOMeyzTuNU9qhcbbkCCGM+zLz7Kj54wLKFFUwcdgunpBdvsr68/weLe0
VFeTGyZK0Ex1VH2UsJILHpPqVahGQNExkjZdoTWDa+CMffo1ykpWOLvGbyhC
vaxw9pKh1mva9qztaYwrh+8udfH8fpdmgvMi3FL3IvsHlrmQMkmzH1cabSPK
mhGn5G0HClnj/DtI6zZqtkSQo0neCat2gYixYQimljZn8U2UZFkl1lzNc6v/
5sOavLwonoFdVLzARi4iDoJbP2yOOwFQea6aZoaRCzqU6MoHocNdtDrTIYGd
bJJSzbp1NPcI3GEH/lJPt+wDteBFM3XoxcsfQ19FKbSlMtPkOjOBFutRa79x
b5y5wOfdWyCgOT90tjH+tkD54fwrHPa93fZ4zL4kYry4DgsYXxI6TJuWvUAT
5xtdmCwWyJEJ/BAZT4fU1PPetXlc+8dOIiXjUO1ByhPuxM6TXhxMt2GcFoPp
0dexZgfyYYoQp39wleEqfcRFK0h9aHSTbT94p6opLC3YI3eXlaKCrTrviWe+
U7aXYmp+QZsH2OuyUgOhj5D1HY4IPsuhqMIHoznh0EGmf7cxuQUblP8YV/61
ENPMWJPsysm5DAAzTPXqseNOtZy6z2KAvq18UIszy/262jH5DjP2vxkXBTSe
TanL/xY+V9f0FiS9kxBFH6fVuQS4hLyxPXWEH0tzB69G1Ftn2X0a9tw43maI
5UTqyHBugMqCM0VBBv+Wiczv1qKMdlkRKm/zpq58mpwuTpRa4CD/8CQGJ5Nf
jySyoDGQbwmhWbGqxPwinr5c0aWQkJBoFBI+mf6ywYOJAilqrr1oa7h3q0kM
ESAK5X8NfFM42FgXTwKwu6C6n+F2/ae//w8vlWFwDHq37f2+3zbWG0vTMKR5
CQtqajqWo62/H6G2BTh/Q7aCISHrVjVq5W1CSCRo9qaIDRUH6793qWAPy92w
k9Vp4llg0IPEP1ZDOaK49jBfTcfUYLzFT4upagy3xo3TrrsHJW9VhFXkxmGq
ri0k+C+RDprqhm6dtcrCfHLGlHcjkEghfPxixhBT1hQs7rOKtrIyahRGVjPJ
caMnT2CWjXaS1ewO2KvY54T7Fo9lzWOhHzMs78pCS3ezRzu/454ufQ6qkcJA
Mpq216+sNTDQpp2AlF5qQKU7JltnZPtxm8ntZLadGYkrF8kTCSTqMmwibhG8
IeK3Vo12R24CfP9G0pZrUiowms/wXaTHQNXVSvV3UpDqXyvh0ObqUlnpA6zR
MJADgJV8OczyHlR7roYAzm3ra1dRdDIj0N7UDgMkFK2gJ0uHYAk17024U/vl
1SqXrn7ZZpqB156FkmHjNUgZ+nZyeIvT2sx+XWWG03CMqpFl4Xvg9EihOwr0
JRCGwCmy4e+bT4MMeBqaGqEt9mJGhOnYOAexwpJv3He7VBPsZrzwkfG0sJu2
RpvPre4rW7GL12ynzIowM3sEd+4JubwjXAc/SFV+k0un+6gyBO4kIgYC9Dab
ZWEHqc9+47gV+ejaQH6WVoqfm8l2I8FpfPpyTuIsl5wviYo61x+BWONRL6kZ
/6qXtVRAtKurHTKvK/r+jbRjKHkNVINtkx9O+xs/qpzZTgRDmioNUl7KEkGH
HsvuIwWskUb9UQW7BBXguWvLQP7U3CgA/ssVLi5JwSlD7vzakpBGrriv2fUR
BP0T65Aqu/QL1lCLbRVB94cMXtTJJsVn5WuEXaykyQEVCSzDuKgcD3meUOOU
5iiue4Px9VLUXznXaLVs69r+h6rycsQ8RQ934RLUE0aaaTzDNREgyl6CjIdg
lSe037jtXRGo2ygu1r8UlcOHvL1c6D9PrgSZhkoCHuX2ivFvxozwau762XWR
CYdESxxv2KsHTGYQ0FE9k4VA7j6NCgLp9J90BepwCcybV8Cm/CxcVbEjIMJk
w3hnvc5bQPdaU/dV3Pp8yfNso2uB2VbbSG9JEuLt2qBdoOjrhHTWizyOkgdU
5dSgVVAzyflf3skQNTtuoxpcwBj29Jnb5zeP4kze94rxzcZU7MV/MfkD0NyH
S6rci+RypHJWox/bvDzNy1d2xqMrElnWaDYvoHwP5Z5rf855DlkyAc7S5ydG
tJvN13iYqU+HK0qS66C6gXL4zCfUY3JRkBMuMo+mOKFonWZXdULboh1a6uF9
BHYnxEkpB4cXKYok9Wr+SaOj3BoUPZREYv29mAX/X3U4wfSlRE30htybLZCh
bqgD1br44FhnhQYoUq36c+dEkRLLPR4WiSi13x8IkXGpPBO9usBacvPoSty5
pGsBXpg0Jd/dm3cHg9cmdzBCpBk9WjKRCEGRkzMBFUsC2cIM9PZAtZ+aawWd
4gb+p4jfHBnEOlOVLgzao+tOtchkJbb5PGzcNni2kTByME1yFStC74lSDuCH
ULTKsUSpXxHQJ3A92oIaWmt5HCGUfHiXk0HabmyoMZCn+DYTM9yOt5Hvzo1w
6zDGXx/MHBqW/fTvUX4hjhqNamyG7dlq6ElcOTj6bxUD2pyypjrIjbSZ3tAv
dy6DeaynWN8DPuV+rQ6qmTtChjoNin8iGMDooqyrcZskLYpp0Ay5SyatgBBy
Fw5hlCGtSHwxrHOsI06S3jaYWK8cOmb04jdIP++w8RVYGbkJlezIuP58DjL/
KUbE+9baP3SwcF4xUmnfK0JDhbCqY8XveMN175vU1lezwx4oC4nOYKW6v2kt
wsA3qiwBR9FSJ3d5kbDeJkWY+GQ6aeCyigx6J9hV3ULMyymwL06lfNJgeDnw
jSgstkHZlVDP5CkuWEg1f/6de2UR4bk4aiTC6cL87HE64JyAB4sJbXZWgVFb
8409ayf4ZTszpNdVCVP8d02yjWifAtrFB6GfcijkOtee57jr6fjjdiapEJQH
4c984NXfvPi1jGObUwdRXdCXiF6A0u8Ds0sGR1ou6JLWWW0SJdlCJW67xVfg
1OLkhJHzGHhqFR3L3lFahBpuTdkOdnzOIdMgFBAPJj0qMBf1kixAPS4uBFDm
CXjKTmY2uboZWiPHOg1NfOUyc44mu63DRuWVScUvPkOob2dGOacxP2YY1M2o
VK18ZQHMfymewVBC20m8PI3u1LfAoFHrmfsvfSJpgfQghetIJfbaI5lPdgcK
AyOKbREgpMOL17wWEc9zT85mjQFDRdBjMuA66mSYTHV3LRe4WFNKn8W+3axI
YRuoKpv4FhEq2Rb6dv3M1sY2d/gYTKVQFR8dqwc+/Go8ykuEKBc0fcOLDYDQ
VhpYrNME+EZbGCw7iEiIv+W5MCEQqhO0KOfCFNvLJT7YBUong48t+XK6Xzyl
/Lw2RauocI6HdeTGAKHIr3+rU2LUk9FmlBIVhRiZSQIkOSWChjx9LSssDsNp
Bef1cewTBuGlCOGEomTPrWRySdRG32dt5x5II2NSyNurwBsWW8mJ5InS1emC
ncyukeiYfrbs6NParZGZjGnJjGMaY8g27bxjsM0Ihkm2oupVnKGLTksz3iGY
X6xxJUsyizKE+uD3sofrqjr+1FxMQ0GGxDm2NyQraTh+pOy5ahU9pAeZPrU1
bHK58SW3yzggWcu/Vq+33OXsJJe60t3NmB50KNF+lZHpUuX/TIcCjF0o6uVz
+2n0DN4yiQGkhhvOjFI1t/5aMtJGzw08yuti6dMfYD7QUL0WhmCsUVHBjHr0
7tNWQK3RW1o+0XMI8CTEWvz6M47l9P3xrGYgCUZAXUVKdK0hbSGat92mufOU
yqPjU+1fko7uRf9EWiXvlY5W+ekooZ9P9FqMBS1xy3pCbHgCBNLuxsTtUdxt
ZY0bpaemGpK3P7jQ0+sbdtGG0YL8Mb6rs4kCUxvl7f1MICyzJIOSGVfYZErt
0kX101fdtLOP9v7E70iJuMXmw4unqWPXLmqVuBgUyGDBAbcvCuTTbYRBYqRH
qDVayGwZShacrQoiSjCvmmOHF6U4C6hyl1GIkY+X2uGns2rHlqKoFs9B10xD
+PfLuxPadbnRKlEzA6n4w5GjPGlWu0aVrrfzhVNNAaecs/B8NQNoVSO56qQZ
1GB3AFKiPf5r+bPnaaQ4A7PwOEZ9jXvlJGCkujNf6ealHvd8w1P4GtZrKia+
39Z9RkDthLi0ICoEvqLI9YxY/3WXcVqskioM8BSMu9GWeujTzHx+odpFL+Ng
hP8Q0de98ifGT82ZF10ylZjpLbWJ3Cigblu6aOoZmGf9p1GWEc9XjMhjQBLB
L9yPqTNvzTLSCBnG+yDe8y6MCVPWjsx0oNYxMHSpmA9YbwcTeLFvPjo0TK3e
0jkV7cCPSqHMfI0RKCh0fQYJzVAUfT/MCNB05KZZ0jpYeD5MvipEee0cSJd6
6jukttcYl4rjPtGVtzIsAwoMkbfSI5TiDrKPKHTA4RRI0znwcCK8JpH2ubFq
81v6eA8O0g0H7KU+qKC5vXLEZ5f97ZQ/4QF7Dekxo8bpIJt4zvY7ESIyxbAD
JBA5/TvgjM6k5YkXRAJg1xqJHvJVerAoXS3AxlsiLFqrqC322DfFm/hg98Cr
U7Uk7urVAC5tBHVr5KGRlT/5ILTytmhyKpVrX1nZdK5pWeU4/5Q4g9EwnZnH
qeWKIgczqtZkSaRtiXO8KL+SIFqVTk1IfcRXO7I6HmwF33rntgcHThnWFBvS
C0FFRSSTw5GYhuxNAOIv9Up+uSnH4RP0lGoJIw9N0+lCwnBdUIeUzaSXM/p6
PTgD3wCOpn+gRZob7XAeKkWNf2D/tIFITkP1vIlcxVFa/bamB+4aBpINxp4d
O6ZPVwXpUNngsIqKgHjqllIMoF3PZMfrkjDmWd8o1himdP2VdkwLhx2R8SPN
tCxwhBnDCxzpAHWhsxyrmAjOLLycdikdJeoGyw2Z9SImU6tNg1kS5U9WJGCm
p/WKRbNTNJcjiLlGmVEoBtQLzcvVjC4OD07IRRuocfr+tFwjTE/mGvZhdT96
oIVayRPiu8BTh9a/g4uFbgVrPfYTBgXbe26F2giI3oBcSmPGwBAsFQHzF8Uz
kPStCf7Ut1GlK/wxZbQltx93dxFdeMo6nYME2wmyimjUTP1nmX77HzxYNATP
9zKKsyqyJB+lE4kSjLYTFU59mkiOd3WRUbRgh7eb5QheGP/kg2SgQSJLjQy3
IoV7ICznOZGrgpLtJCb6J/e9P2I4vMKEFqMKf+/4+qSS2TAFX0aEIhTOfQ4t
4LF3yMJYj+t3I3/b1am6k7e6dhfKVbrgcMrXK7uIzYVeQNthbtbvzeo1G4lg
eKFGgtIk3VAUoMB8mCxvDpRYkcKYKsUf9Eg3XJDg4noon8k9vh/vkUSpaZwL
H65gqEv07rvDZFgsokavNqvfxeHp1OtM5NKZFLTjS/3tL57pfqZ3aLVRqH/q
qW0FkGq9mPDWAJhrGpuaBaYSvRaFTRl8YhdTSjD82ahJ4/7Z4czwKIOxOFxv
/9JVuvL87JAJNkhb/K0eBTu31URc53WpNV89j3qMYBLDT0BCzgzZ9SKJetbq
fP0DS3EjyBUFgUJuBUAoorqB4J/0Vgy/lWqPBo+cvsmVDSilWxnJsjtKiRyb
tVI9cYT99488LH5wtiE2tMssZOqX5Ph7NtphrKdPR7ALgm8xs4NXi7QTH+0S
I2K0hDS8Wsw9ytP1PvYvF2tvqP91L8ftrOBdcaCvt19zxpHh5SuQJCdRFxpU
Q1m4CU0JZSqQFu4jUrx/44UwRQhxsqRs0IetKI5d+c4gCRxbQzTUiJpEBr1x
mL6T1ZbC+u36SD6vogJK+Aea6u1tKp6+6wxXg3ewgMgPI83R+0tUDV7Ay/Hu
xZGNENNPU3W/xtvD4jVbf5ZHrrK1wK7Pjft8XHftdJKCKdeE5O79oZeNFJus
IARs9mi8QXW8NencL3N96bWclSSet8Mgsx4ybqDiu0Tx8c+uUfImXmRXgck/
6RX6RKGR5mJgtbrRAEX67qne5Yq3NHlrzRiyr14GFYXZUM3fBqPMfS/ttQQA
B/8nb49BJ8UW9iU71iRgk+nrabTS7mqBTAQ+TwGn2ryfuCPNLZCckO/d30sB
i7RBXX7WbucvB1iwT9oRGZBRCgzNeCxRPDJPuHckcE9qwEPM3k69zt3Sn1DF
bCLf3BpfB+ciDEyicRCrSDvn3WYzubeUOppXgV0xmYV27kDeYaeAZhpMqnN1
F1hzY/42sDzPXD6NJvNlQPAsY7dhCA2ir23fy7h/ve/ewfGI5vqMRZAJeMob
A7Sb/G2xFXR1nLtK687Ja63TG4zcHwhf2567hwrvN9BDgJ0xUAtcNdHR+nc+
N/rjNzKRmzw7XYUQWcMXyQ7AlRUluI0IDzpgshhNIDR9fcpldhZa4dpIzL3V
h8soZypRKURHyi1hw44KcVumAkILt+4Ae25B6fpkwB64+c9nglUQ0WWO5rwn
eYR55ogDEvccZlCoSJQHHolpPYWdxQwtMQ7gkp5aJrujGgynRObBdUcz0l/J
KPEXK8GzW+gaHZxmiru/wWResKPoM7KX4zRWTPkKdkHenF0VIDmcStbwrMLp
FL0O4xnfCjuOXx8TkjxgHhE367vn/hFzfhxcIN1DGnzr8WoFM2uQiwavvHzk
eSJcN6eBI3M/7DSNe+cPrqutezDD3G0cn8rZ4F7MRr8i8nx9VPPOsWFymudY
kBHcXGxCbsYlK91sA+NGPikTLce3/ruBxyU8+Mqkv/Rs6/sPqBTLzUmLCC8e
x6ooMij+g01Q7Cln12WrV4wja5c2x2cLnTl6oK5gx+efA4j5O8IVG0/B/ie6
fH8fw54890SyQ3vEd8YaivR4mKTRcQlmJnaLRGe/d46SB8ltbLISMfa7BSzo
InrGIbC2VgQOdQEkHnvDhOlksKze+rnl5ExG3NZYKNQimy++IwlpJAYYHlgc
6NcX+APJsll1hnwg56P1esH5ISAts4cQp7t4M/hBxuqw9OCA+DiguIz8iKGo
v8gLZZnorJzuGtQZdaC7eVPVM6HVbh5nRHi2pcbPuVzOekZ4cwQvk0KvMOb+
ctKcjXMZgvKoZeZdkACzLa2Nn6Y5ze4js1w7wRNFyVSn8DZClxq6x+GD1+zj
LnwD0I8ZDhKqzGTAipwxh26fNAeg0MgP9ZbqK6qTgOCNBPvnxiaGQ3ghZ/FR
q0hxMr1tmExHTC198bFfqoOGFFu09PQeta/pA+mSgFJjhEcgpL/DjX5x+EOX
SiGyxOZECiS62aPQS5ux9K5OVQLmngsZRP5WYtY5jVds8DeO7dBs3zktBhhJ
X2vdWVooQO2oCUMuziXwOij+PqTNwTglQ8lsJnI1sghj1FwQiX32AtvHTb2r
+fP6Oxb38/4V5JtUJF6zN0wgjUAe1KlXcaP5DUdA49j6HFj7G5eRk6I/PlmY
hwmcRDDK9uHi6qjLWidzdOjBSN5bwccNH2O3DQ22vt1H/q/OuMw6SaoSlczR
s6Tm0nQBkxsSzBpWUmqMfnZ8y43pCFKnXYQHeQ/Cc1fP7MXsreRnN8Txiusm
k3Jn2E3rd+d+L7liYcTVbYWFOdis23pFuehcxK+7Y2/SMLN6wyJYefV7JD+5
qCHF8S31DVVi2IdHy7VTUtn+RibL7JUttz+XO8a1NwFvjOqD46lrEVm/ZhZo
JakCifjtYHlrPOTvO6Snkx/vhrDJE8OpWq+bvJ3G8+AreKnLL72tjC4j54H2
5fKUwhpHg2UIrn8gnN3YluklZb8OSVvc35YZrmtMkFU9oXQQhrAKSTfvbSZk
sZCXkU8HnvCrPSrG4UC41dfGrtoXJ+Xg3JLiX3IEhHjm4wCfYf8/50HJFFZb
V4YG43+qEvi68RNQN7+rAumSGGFvaJqkJMD1/9OIBzUMmeed4pBHMl4JL1An
rSQmqQ9rB98ENjZa7SLIheVHxjC1mxt/3XwUxeYCupvlW6juG4NvfZDyo4sj
XPrnE00BWkTTj3WcLRBSVRF0BSu0lR51HJaokuQShO5BoF3LzI8znlsLb8H4
5/PqaKajbMtqSTwMju0j/zmXcW9J5k6Ih0q1VupcQtGqFTl/IGfqHWsh0myj
vDBvych6heJRPlMdFMhlrhm0u6mbjZNvNIRkyb7uaq+jJ3FQuu9bzv7LrvTc
wLhrLDjGKUdbRUvyHN9mrtOlgTMTQV8KBmPcjUimm/0gaHRTP5OTS+76BlXm
B10CXVsYLvr1gQ8KzKVtLA/R2cXjQS4NSuo4SrhgcG5D0G3Ib7KjOhc/9Gfo
hBJiUP8arIPXqFQWsPX9OugudrZGSdY1lDBIMLyjcKijODMcvJst+uLOsCt8
ooWHPqLgXb/10gflpkGdJYpafyDwx5YPYlN2dn0G9X1Pay0B+x+RdlrCenAv
KWH2FLq8cgrldkjawLfQGlMznvF+WnEdz+wFIQl9Kk3T623o1poWdsNawLbp
1DAvi32OW32iOdS/q2sFcTvsDNUmjqRMG/s17DN/+qTR0ePB3970S1XVAZJy
XezH3FrYuPTHkHenLqIVeCdHGzNjCgh9nJyYw/NzP1cejBKWp+Fwd0KPp1v1
jBfD+TNmN+vsqmMS1hhWqFULX79ylgCBa4lKZv60QrF89BRqsA7bWi+VGZvR
JuMGgMDihO5oUFdK4Y/T3LDtZ4t97BK6aHffcjvfEQOl7a2W7vx8ssgq48hj
FUtet5bDeClQ8+KQJPV+52Ogg9ZuzZZRb1a3HzRdjT/pVl9bhRqitkItcJPQ
ZIQMrfyFCeOwZtfyKdAGx2dRt7i0WNxTKuJ5jk1c3YstVWa/6o2DprbYujdt
c22d36T0r0e1L39UNYFvFnF2LU8FevCPBV6klx89idPX2IKTjCRL+Se5+qMU
zvlWAgMqGODoxE3H8A13qQT4m2vtZ57KeiyTIsQnzYB5tDqQ0zfTSCaPQEE1
LfLcVcLEc6nUl1Otcl3R+YH3grzeZ0VlNKsZqe2KCgQdMoVxSkiMM67xxELf
hHYBZU5jdqur0t9lcVB4WeWRn5n23lyui8XO5LsY4CZBo4kc/V5PXQ/lgfmB
vXRWIi4kVBJn2YG5My4XPZoEEzGLkgOGA1VdN9W4rTDWraz23TAzlXf9oK2A
6PYBqIdchRkJ+3jRlfNCXk0IwAj/kt+e74SZzCD1sbNCs1kkDvh+Gj26WsiC
/hRB5CbK5NM2h7FrzfwU7Uo2KWg+pDfM16UyV1HwQPUyikoPkOfaWIrkCHH6
1rJxk1Xaan7Wd26jVpZHsomaTItwqL6e4t8+ZzJe9F0HuhSPLt9PRfLOck1p
DzHEXZHBlJQQcsK4Xu/YUKJaBhcIHTdGQnbazjwJYfInLsBvSwd2ZWJqnu/Q
Hlcg+C4y9sqesXTNFdOwhoZW7/w6j7wG4aDZZwgMdINZXaiDDX6rubz4QLvo
3l1c/a7LXIGKe+BoJ/OSv/T1/3VsxBSVGuFtU/BYzJp+550bXFsW6ZmDa31b
B1r8ndCIVqTYvjw9rpxmKHgAJVbuqWfg8AFEsQVmuap+lD2gnuqdH73uPIem
7xqR/T60NIknAUnojRgaw4YKOKk1u/T6JZRIugdPNQY0WTdlrTQKR+GG/eMr
rFVMjgRqW2fVDSUVRVesw5MeElXVlPQGKk2pOxEIRmaZxV5f4etV6bH2gyGT
V7pnGk3y7aj0JvK9MvXaCytVbWKFoZQg7YK3mphdnP0x61zHffJE5gHNskiZ
mY+h47JupvG6NzyziqvS1g5919QH7M5CB5bm3gmn3DRxHPDULjvc8ACFG9Ca
alGEcH1OCW6oOZ0Ol+5sUDKdY2ww4K2MRF4qas1XLOPSLIhPnhM8enEPodQo
k5MMFW/M+G5lFTg58Vjn0VY84KNbG8GaKmW0cTHqe3+mNCefPxb0Nb272D94
1guzXWDkn7xFt1hmGTR1WEGDY75XrxsP0xQrsvDE5oF1v02e+BV6NQ3XN93n
UOdsilTBD1k2SiW7C4Az04te5tEnFvYW/dMixwOnMyprquT64ArhAaqrWA47
V/jl3gPs0vaRkyZe+Ep29bOrskWfeV7VcaXp3oFfDipA9vQZ6zMqu8OKcBBM
aSnuZ3MUGxPG+0JbOaxhm9LEtRyd7D7os/LdojaFrsQpQFjwB6fdlO2bb67W
l75D3M9MrpxIZhGmVHOJVwCXG5SQzYN7/hASXblA+xx1yfOPCIb0flny5bf4
6dH3G0M13O790OhN4MTQCVuZyvXNATQ1r2gDHmBIECusPr1UENw61oyIFl6a
dvRG7Mw//W/itk2oUH0Q/FLEeGNC/9Qrn6UH95+t0PWbZwMZrO3HPA6/FzTo
gQiupY4stleK7l0ZbpPNGbI3Nr540ISpXju4O7ZKB7wpcI77xvjIdi8zcSbX
vC4Tk3T5woyznWwmROW61lKgRLSCkCnWeYJmTJHJiMS2tFxfwsHr0l8TLnVt
Fyr2kcXj7Ad7qeonCVZs0e+qa5ce4ex7dhDCWOSeN87MvxMvYIeXyhyn5AYI
S2NIgG6XtnbGl7sgo9NS13EzdqTKJzH76JQ6tYmaNXePLQHWXr6DX7L3vmt8
hi8szs1F1krTnN/TauIu+3UCsgpW6zwpYsaLEIv7OcTOlv36K288GiUky7dA
EU6oU356YZeooCc2LQW++1Mpq/QnA4lH7B+ftNvT8nuQYvKshwAWLxL+A9ei
D5h+pn7S31GQAuQq+P6k9l4U6rxh/GcEf3gnJ0LrNvlih9F7peRl+ilcY8Cc
T9S9PzrobItYe+jn7dOnLdTZl2kTbIIzENXWZYcLJGEkaQzVbkG9UophIOtW
VoAQm5OLUKF2m5wm7eJD9fKWTWdlWkxLn856juFoy47iqhDkFNw+xn4oWhl9
gMC1ttC12fDCdcb3VBsTyHSI2j2MMF9Fa6LbLT1JqpCTMwCqnnzLBOevkvPU
1wVagQm+9bVWSApDSjtL3dcA2BKJiQAPPDLgMFciz7gOtIwfPUMxIuM/KtvF
oMhHxf5hlv/FdxAY4BEiWdTmAuKM7Q2g5kdTLRmUKa1/PK2Nf/xyIW6hsAIF
2UIbpyTRxKKpzj48ZIlJPhncBzWt5LS0O0NQQQSw5Hx15gJ4f1UazI+X60Vm
el+fWCkpr3UIG6kyWQPjzS1OPvvOvXEHGqsz9Cn+M5OHaBWyNYFNJlu2m9Mv
BQsaRFRScT8Z6OhJpH+Z7CigXjkpMKrRk3maMY4zyz3i/TuQYbPtmQdh7lKx
ksfY3dv+rrYBDg9cvG7tFr5HXMhO6h9IU+P7qtzYl5dlqlY3K5Fk18BNGWp9
1uZrPttHRUbu3VSTK99UUFA1lgOSxLMlIPRFXmX5l9ukvE7liJZlTZnLhp+a
8Ufyuv1Axek9hEIWeqnb37TRQnq3CdicDbzeyMMbVEsnRLR6kXw3cpM3mAnD
H/Y/l6TZ6I/6nvTqUcGB5CQTEKUZQlCli5b2AJfs4OkxZMwySZDr/VVLGumn
NI0h3JKbs6EQUx7LyMEykMmXYYG1/uutdlYmdv6PMPP+F88wApRmE8lNz76R
JmQ7C4ePZJbakfzMhvtjkbuV4PF7wEazkPYbmiMauxT7KhsMKiRvZAXEvyfM
htpQ1qx03UOqrNtzsRSnyIonPntVvC0lDOqahtCnylaoIG/zkDULN1QnP6Wp
HXKvGWxKPXkmdN2UH+X7awF8yJXhNUIQjv0ssvinCNxxrSIXfDj4N9axWtTR
4kGSt2JrV5HZFV1FYAqHE+7edzUuFTZ/m7vyDmDLWpCtc9x9ig8M11zY4iR/
WHYPBOr/XYy8OaDwg3UjzRaCUCczA4pfqh6fdgKI2PMhhKhHioJ597ldNoTl
SqZlvok7TE8Q3ryImn+tAyVmCM4+kbLKqLjf8pSFNh18M3yYI32ND1kyGMfF
tn2qH+p31mIw+VgldeVLhlaOx4MhuPnFBLaXh3rImoQ0rAn8xQzrOPihgxni
OAMV00ZaHd/rM2Yx+yYX/HzF6J64Z24d+GNr6xvGiUawGQbG4vdhUF9jEAy6
LlunHZnKT7S5QDgBFEEh0ZCj9uXhCyDztWCENTfkJQqxUcjwv9r0Hc0ym6vQ
q03263CdCkSUXr/VpPoQldDy09p+qXW+Ul4lW0zFUCsQCmxWma/WcEYEEI9Y
NHX1SQxuM2fshAQXx6r+8DES+GsbsPzHATBfbTiscO+R73q+v/98jywajfcz
rKkafJQY900susQW+pVK9orAAk7+vjsYC8AqOJ4gPCXdcQiTRAD7QPBb/l5O
Rfg+eIpFpp351GT2bnGTLDvnK/Af56Kkh7QNFoE4vYFvJSzxCwElaa7KZX9M
PVMu+8IBX9y8HfrvBzwSCMNldKFELnzEevWisKa0yYSOkbdf075Jfg6NoFOa
uSOAmsHmVXOXGCTOTnE6+aXxs3ikeTcHvUY5kJ/nQD2mnG+IWYY8xy1O9Nas
RRyd6rNJsSOelhzXMFO6n8XQFH/uJlM0xgz/+Vx7K/9xPDZt2ecBFkxnohGF
dm0Pp0268P98ORBqKzBS8Kwwgvk1fPLPrOFj92kSFn8ufLHszWjKXTUndP9h
bof0kZNKLCYuIacc+ARqWsj00HQ5Iva4id816FLyy44cWNeR76j8ATM2hMa2
HylLl2uYJAQHKrZAQMXU2jmcjgTAo0zEeLZC16A5QJrSf81qliqAoGIir4ii
q0box+v253siWAS9FUx6zaIHq+Jgw4kZ18+MWRyOl2A3UAT1V1Qp5whe26Yx
5GycEyBmXGTJ0KhShueXKOvYA7eYZM2gxJTfGEs27UKBp75EsllDcdde2n02
j7VnnCnn2txCcZj0rgJKdbEJQ0H1AU8Brt7QnyhPAhg6DO53MzkVXeBrUjk1
8HskiMbmCIrtTbHv7AQ3NocnnzBrcLxUycNR5ivYT1NyiRNTQluVVbDo04d2
It4931fAV/lD8YMvK7vYMNZQScV5BVUW2ZbI4465eMEL/DigqCU7N6Kz+Uif
vQ/cRCPsww4tzB7NqEEyokLucw6p5DIY26EVKSg3DVAcL2u8GGux23GfKWS6
mePas014VNlwiYrdA5R5H14dcExpMWQtr3selddSXIzloiGuLjcdsmwsw3l6
XmB/vLFaBC43KyLXANkcitd07rdnHDAQCZrkulxEvUCLsozIRzt0RfON/Z8v
Tyw/5p3rxJ5Ki9FncG8QGHOMRpZCVc5Zu0pbj3lQfsknKwigL9k+rgNMq8UF
ERESFKDim3At258abiTuSOLuTr3WEDaB/Q9U2z236PyG/mt8kKOroN4aPZ5M
YbsHDoMEhmQwyfXwqIjXfB7ZAIaDbm6pfD0UhDosQikZdwMkF6ic3vQeTWK1
mBbGTwLieo55IH6ufZr+AWOQEmIosrIWV+bKOdbdZ6ke3w97WT/4LU4Yhmhb
oGZiI1q6QD66MqU1HtEzv2hnSaZvCsof1zrxpuhRDde531aIrGjYti3KXIva
HjvECp2cxrEbumGbjpX7AojidJXRcQ9D80d/+FxYh9b1fPYzCCSj+BDLiTey
odiIEtMWCcOepeezEeVMRMaGZjCjqI5QaWmfaKlqZxE/xP5dA9RXoxfsM54E
nLkU0W0raxbttUXQK8PlfjI8fGVM3mm3Cg2nejMPoIqJb1a79mm9Ns6FiT1A
E6ozACUjWNfWlCcRRvMgybeCSLojNYi1MFECx2+sOe2hSrUBW85jylAylGlR
aLxwP453syFpnp+MkvhLiM+BC9QlsFbtQvDyMrO0wz9E9r0jJmcH40i5jbi6
kM6shTdig0KorE0SNk0+QdhsxmVyuBpvs8o9zv4XEZyVPLNFz7SsM8jDS+8p
l9rSr5VF32qt/ySMPKBVuuahgOuRt5+xoGB/UVGIHLzdi32Chx+t/ypeU8qc
WnqDlcRzcjcfQv3TQRSr2uqxxssyjyj+6Gma690t/It9qlSPTNXr6JHvVjZi
E4BRFfyI9G0kFQcajJ1w6S7UVSirZqazXa0g76WtsmAjWttG7nGA32MjsfIk
6fSIyy8TuesaF3bBqAfoCUU6LjYKhVlo2tIEOk+XNigJoMVReWzjE1uUHFlR
Rt8NZCLvCq1r1GSMvTgkRPqulSfJrG8UPeEcTPtuAOEmoeTV4Pmc6yHO98rD
gHfI8rS6WX+M8Nue/GpWJFTuXelLGbXSiga5o9ew3JqSJNeDEKfvhSNaNkQG
vibhvXoWQHYmBM7kk98++FhzLGMgCE9zlRx7CMMTDmHqTdHojwIUNLU9mAOj
0L4zCaIBSSc/OHhzknVTOG4olbVYmAChLfIC7Cr/oFlnO9Ewe5GhpKc4osR9
E1CC/bwil58rzqsEKhlkkg3PYAquazQ+IOHZuP0GhZlsEqfMgcMv4KL0ymQh
gxcdKQO8p68AdWSL7BM7Dc28J3zdy3AN4+Jj7+FaikU40dPkW0MjAr7c4WMv
duAKGY0YDlsapCT9Hw9pzEFfKYytMMerkUdi/UWgd7+zY5cTfl/Po84CtpIC
C/or26J6e/UAhsFwzwn60Zw7JG+bOwAaQoOKoWDAwIEyTgqPMo1kGXMJw47U
Co6UI9dbkxZGBiCwoV+G3dsOzURKKrMP9PkYfW+IZPg5yPEgz/gHTe57pamv
qwum2ICCAnagkgdqXxrGObEm87BH3kYJryoUddZE0oetF1cI6qOq8N/0rtUH
RFFWiMWYCrjsedGqvJhzKcpXa8qy754mxptjo8CcAVNR6k5wTjMyR3COkuvt
OWgv+wd0AkDdDvEaRDxTFRsWlenMF73KsJwab1fvWSzkNTnG5I3wGzutRSr9
2NitcfSkdSXx/JLXQWSs5mF9PmxXSaHZk9aWZ1723WbzZqS5BsgRuH+tG4kW
IYR8c7zb6lH3sVSRCSFO8Y+HYwGdFc0XAfC8fm0xtRq2IMyW3TPI5/6zkjs2
Ah+7ha/z3hUpHOGD3biRSXj/vqHAUMd4M99bMDjm0Ki411ZIJQtXDvfJMgWL
sx/kWQeHR96AKlo5pd4vdo/6x1WtRTHl4XbmKnaVWTeLavftgYVpZE64pzGf
8WxUNKRCdKGAXAJtnux3DYuTEm7SuM1k/5GpCCZk7SdnaloYsGxqSp1WwZ98
xltDCTYkNpZiimcwnjmQl7q+xZJw1yC6RqZl2yivN0oOhTCWTqXAiiXQmzdg
CXDJ6PwV4ZSLdRIXjMhlw3XlHdyDhoU0mVc/M2ru5RyHvmO08D6n88nJBUGz
pCF7M612rbtVCxWU3kfgs8CS+/PCUBg8LaBq1tFKGsICDu9iG/2I1f3cVC3x
7SA/qs1nzurDCQ6rIs06n5iwoDixbr7/+an6RxFTefqfFij+uhX1eOhF2H/I
fnkoVurBekR5Am6QQ43+fwbiL2H0JtsaEugyV7bNfVNriocDugbQFcOoCXZt
KbDx+ZOKlUGR0bKzKlnlCWopoa+OwgpRGnErDRpBVtBm6J0RPXMa/dWtBEhF
Qn6AGIbDuJVAOJDx5r6QzQ9Ne41A5Ovz0EBxpmIym7VN5CeUAklWxSXXfwdJ
hzYkO9EmvaBumZo1k9TYWKkTdDgjpg5YKLIRLSlTO3Yev/M6w2yb5iLIJDoP
C0RYO7aKsoVKtM8OuPnh5y4PwjYmkLR6G3AC//EsLLYrC5bRUXauEEnjM1Ua
Fd8Zi+wvzyrm6lSy47UNoMVxqakBtm6gaWeUzTNkjxBhP+9ZjGbz+taJ4x9A
18cxUIqbVegsN5akcEg2N/puyuPF5N7w6UlkX+I9853o/gXu5qUwNKAI0BV3
P+JD77DVWdpuYiKJ/Jl0TERPPH9G47I+OzB6GLdBkTpODlqQyXdYr/3ZiVMD
MtDXMsyNuPIbmTWgt4A9fn1U5xZEHDb1PltqVhzmBUOkc3M76T2yjyDMP0Rx
B6AnBxNIubnqtTbx7AEULKopDNFvOzSvaNlFxjmR9ZQtuhry7UYi4VdqXnah
abvpuIhwOS/iy1oZSqf48+Rr7/1ZjMlseZ5r0R2F/6qiHlUh6Es6XERb4xZ1
ezn/b/PkPmG7P7sROcSGuwuui5lubW9xEPBuAt0dPVkLEFp0KuzOSo8IRItw
+0Zt5q7gOOnqIxSOVbbRBPiowEBEytyAJrymCJZLNKLdovi8XaGPg/Q8kU6r
LfQqP0PXxUFGI1AvomsZ1HQTKxZPImtVW+jUf3EyI/pjqsRlgEGAI04ykoJd
hAUNDtik7ucIF7X5m8eU12m3PjNphfB6QPO85ArJA8yNyaMN2lkRbYOG2xwV
vpNr63gseVae01NxiTkGmdEmXE/XxvgACh5G6IPbMD3F20sE39JBHbOSsSv/
498qCeE+UKx/x2x/qrz8fp7NdDPPU+9Y1u8yCsqvKDF6N57q7bEjouyPUFqO
sCjIOO8+p1b8+0w/yb+LKd8W0i602D05px747bbvZBLf4ywbf+0IoHDZ5Z8u
XAxY9HIlUAy6VTseR1YWJ5kOCS98yUsYyuvMezX+5D9PEndo7F1iYJpFI3os
TGel5dNmXYcQPeMNRAeJkzctJddc52xta49MgyMud9qwmC2NblIr08IZmhMp
oj522jJ5siLHegtkRMxwadWoJfJpzX1m8Mu9Xn7EBm5m3wR/RB8LvyTksEOe
ZI749A4c0VzAu+ZS3KMTS981FBOq22MAHKIH6ut/g2aSYKYpRkLvB5F6+OWE
ovgJnpIyJVOVSN0ZNMH1PfC0znDrCh7LAxOOStLT7oWda9paxNmic8ULKuOg
aX9Y09gmL7EtCE+f3m+OwdmnS3QN8C6TXMUBvLkWJAiMVESqzYHBEjYKRFaW
tTvpty94azzuGmXC3+GQiVhHVlNNxOfikV0WoEeOhKcgc81B3zefsyNxJLKl
pYeEBo5OmcdLIVWT6hRj4M7RHr870sGvVyNO5kIoqyRFrk8bL8ba0M3Ff4KC
22D+BZo+ka80RzowvRi6KXc+yJ5n9Ah2MXaeCqO8SV0YS4jsX6gZEP9eo+c/
+Nm4DV601CpL+3zwxnVIw90diRlzRWsRBWVkCVfCkDBsUbdYuX7AQvP2MSZK
Q7+87TlUQxR8CV8dBCeZnv2HI6CjTJglCKbXbXAv5tjrqEKbQLI1vA9THyUm
Lr+ymLXqxGT6X4bFHcqXUrW+RzCjx5pxXb4t3h96ERgN/Crqt7AhQKb6IC7t
s6D4pLhltbjUjOP7HhWXUbKI/ZXXBTCiH/Pucos1lYm3QF+UfdV/+t9hfntG
63UuJE5nAjl6ajoaGrRVsmvnrTqkViZjCGf5ZHsIXclBiFAm/bATlpU+5Nbc
2m4QGhhP0B4jnWmIRLhwSO50yXrspvth0og7dfuyrMFZox3kZ0c7kkll4z8K
pw+NeyxDaB8k+/L94CI3i8t4e3YU4BhQ1hLyIkzvCx5bDmlA7IAr0cueZyeE
naA4s4FV1N2cByTNkyKpEmKfpAv6Alpw/uybisDQwvnmzyBJS0IiHHUEe7Al
WEGDqb712SSl+WehctSZO5UpRMhy6cD2gDVONCdSwe9iyPCAxqGjmQqJnLni
nrQQTWLOmw2DYTFzP6k+uLkaSxNnKRabACPyq5qzIQMezHF4WUlQqtLq67LM
WAZteSKe+xURfj6HaHjKuAW6dbmidfHYG9TOI/Kib2bub9x5r1BvF3ln1TaD
AZ1xOj21R8oL5/FA9FVdYirGQ3P4ADUUV+8XWiVNL41T/Bf/fVoFFTuZbmX6
JXAlTRbYvuR0kcO6XMs9oECZ2UY6VcD3oW0LFmkV7mvs33t4MYOufPi30+mv
X+dFCSKJK+47tmrVGqH8Sp+N/hJKuomh8S+/FBK3asfF+SezUwWXnfVVydcp
T2O6iFM6RlfdVuvLHfh8mv0si+NGLpBws4pyKkeuXnvJTvLKB7sXjZjxv6VB
bYOpY2hCKLt9S72HSz1M5ECl8I7nirqKozK87ZfceheLVc1SNLBqvgF0BBAu
HWOJGCSngrrjbVTpdHDuHvgMljOAOIIUejlYVx02L9R8Rit/BjSVxmdIAaeN
Fi1EVeR/4vtwAwKBWxIBR5hnxNmQQ2b5YJFTK1qOgWIi5wLCEC/nHfx/CdMo
/nBJvxxNGnvVVdGRHhi+9JofemA9H+m/8IyyzOEmhnsdEhOrJP+HNo9EknMM
G0FB9Ztt4kL0ptsU25W5XczV6yUBvzCQzhsOXsXZ0DL0hkpmLcFJCHnoHo05
ZBrlU+WGqctIc+7StZsDlXFSwTcqHI3EJQpzFR+G66U+6ud1CHu0CnIv7T9y
MJqocD/dpEEF2e1XbA80L8cBtu4zzcdY6j9jVpe53Zl2ELvTJVNRnFcT84UD
bNAfFcqJsTCGTy8VCy7d0NDKxVxbYPB7O9TG0ZOtSo4ZTWZlBzj2lyfQ8ZEL
IXzf167wjLg4o29N2TmEEyFKkjJz0fdHYACw+dFwonYtUIcWacCXseCvz7dg
6suDV90GSeuB8FAyFfXdT3WG8k7JBLvoJ9AeTZDlMWNR8X6U3D4wxFriOqD0
q4jcDnYIVh75lauTIOlkNflc7y1mfx8WeYNS1RnkO9VS9JO8O/BsCdOL/Ac6
/SC54TWiwe9CZYOKtTESuPiMNTZM57YXCRYJq+elbNZrIB4eSOFFL2knxA6R
Q23ehu+tU1tZpJffOEHn0s8GIKX9QFsNRxGp+Auau01FE41uCNs2uG//PVHb
aHoKoVMpBicAjk2OBx3HsX0BpZo5NitSSNM5/ruoBp9NELT+C8mxW6to5Br1
CGYAHhZSMOHVoAAM2+nCvN5UHOokJU36h8hH0NkQSMTveWLzZ17EZYxDMNB/
o3awcEet5a2J/j9JRGzq5QsbsDnb8tS9OJIn82GTijuYqWnCOmv63Jvo71AC
yeM4FFbTTXZH4vo0NV/kLZC45tcKsH6A4OBvsb9J7w+3ejFMK6/VITSGxmLi
uQt9+jryB78xlm8H+8CMehypIEmDrI8LXzOJ2h0nti5BQ9TU7S4awNYYo/IO
eJRHTpOsN+dnUtHqh74hW+5/6A266G3p3A5OExIEC/TDJXZsC+3w0zCKmz73
aCSqkHdApnd6SbiLCAqe+TL48pV+wEXx/S3dSsJvvJnuF17DD9Op2Jx4JQZD
HBjhaPxlnIq2QHEJ/9gU9yfH7uLM7FCga67HjHDiiycK+FKWxPlolNjrMUoK
8Ges7Pl8dtIFt/KnyK94rLjRPnGrxNVNqZgkbtQEm63/TE0MehIC+QtDqKZ0
DN/Jskp7WRk+mtsOrceD/M6iW2+oqrXRKHZMqswYyAxeGB8GkcrmotrGz0l2
ecnWBT4NHN01c2Gla/Lf0apmRC/wzxhKG8Mr1Osb58oYhwZ/yEwF995BbIgG
rMxT1Q+sfF5SvsR+zVqEpdNBZ4iXLPDoUO7vdVn+cGy9sLJW8P3t2BTh5+Sd
QgjPxPAbfr/8C0cFi81qzFsA0YUiognIEvt6/581tOr2/yye+oS1ysXSHxx9
NdzbrrDltJJf8RucaCX+aveA7QIQ85mJO5c+UanE+rxGb3vjYkopA7Ewk0OX
6wK+b+9KJzPyWseQouwp1CIS2/m88x4xjZkYD9vlT6msqIoWR6YamPwsBCh5
lGodTt/ml7S+PDy47Cc77JG183Q/4aXY0bmVjOx2BjG/Crcc/760e5rB68li
iK0L6B9mefGfxQ/Nfu48/DSqK/zKPNlmW6mcKWtdI4WVHw93zAafv44/b7ey
M8Vucd5Hb7gcPjKMR07Ok1ZoNbk4uI3OBqd5FMtwMNPeU3hYP3+DD7qi9lQa
ZqcVGfU8nLjPLvEokQmK/Z0fhY2W8kdCYui1kNAd+m2v+j/T0g9EKCkL4HcX
7BDqy/6tsurMjjwugibJEh4IsPWNI1KmFmzTVNwvv/8wdN/atMKumBmVIBoG
42hPR+7wVh11EeucGKR1DRd6sUeAkM2+Hr0hS4P5XlCK7TQ4aj0fD+U5Imva
14LIukT7+9g8BWD2YWhHFgLhOMwY3HORS6Dd0CaeEdH/Kyr0TYgxvftB2ufO
zBvVNsgWwJjcM4skdCRHaINBACu7s2C9UmLUlOtp0yFM5o4kDPU8Yjl8gpMO
dYIduX3pMXzmJ21/fliBuc7FXkzDLwmG9oYSm10eX/ecQ3I2fShoiwK19kKU
cHbDQsOBRARtdVXj76L9G4blRaTXrbkNlPrABiLEZOoWEl1UpQRoialmlOd4
y6qIO+bFAb09KZRloBTX7DuOuh9nq/y3aXmwChBb8jp9WTUUnrT5NOBxILm/
Z4m1PGwFyGVpATV6lUjjsJ4vLc5uWILb2zIDe04hEeNV5H5C2cmMfyNZflYM
g9H0PDsY1hywY6pHUOs/OWkcXRsSW/N9keeSikS0pVJi28IBZ5qJFbVLaDhy
z9VCzkM1v6GhobabHyZYopuZeQEdxrVNpeDZJ8AKC2dHz4tFxX6s8R94qf4J
uwtwngwpjWEmpQlcILCMJ/0APw8XQQqow4SDDPbfFHKZ1J2WV2ro/1nGkIOG
RP5paZd+qXkxJ/BsjjjzH993ctzRCwTi+GXui/G8qYPkfmkujQHLVAemhJ9L
fM/Fhek1CQG7Z1CCcpzcY5tfbjquEg8xwKeLWBqkmTd3DcjW9x5ZEmXdu7YJ
qXtTEksvypINIJT8Ke7asCjsAmvWNGHk+Usw3Y53gEEcw9xaT0UBkGPK5gog
CU9qybWuYu0HA/ok4EhHzkqQ8s+S7lGGxyV0+Gj14tlQdTHYfHIaTtqcXrfK
/Krz3hi4YcFRl5GdkY4Am17nn1ZrwFrLY08gp0xlIbRzrWMyhZZ6TsB97lN4
cBBZDv8p35r0AphnDE0bMmtvIQ1k1RhnLT2KtFXPPOY+1sPqPxN1Y2IXtrtf
bJJ77Jbzkwl+sdYUKNUpE57fJlF9+hHlmkGES/yJ/T5+BRY3+xphmYmRFmqW
tq+1o4SWVApEY+/DrQBidy18kKK1JLss3kBgXm+wVc2OhZzLU0k9Tlcm07DG
99xOnIQrCetODM8d2PvUoZFKvHOGUXUqdpfTxMwwJxaTehru8U9ARUzKJEqy
oYQMhe+ww193V5YkvvEbufJAn2UzYKbgSNMalct1y0Hm+LQ7b7utuN/KTANH
rjtErkOwfHe3IPMot1cpFuym+bKQprk/O5J1FlTxTEUHHH5bAm7VtuO3xKfF
zsfa9tYOp1nL1PKuJ4oz3Zi2MmnVuWFUjAwQgyqSGflRyQBe+2kNsowNTrJC
U2wUIKIJo8XE7anjjb2eg2t1MmaZsjBdi4THnidWN36WTWhic6YSTzXKRqbW
VK0cdOzm8FWwASf9Nqu4skMQkFL/TtgLIBpSkM3O4MN+jfZ7wAcYNFaD1aND
gAP7UpcZgAfGuGzKV7JVSXcmduR0immZo+reBjUiIx6KuRDV9wJRFAujnSJH
zk/EkcDP9h+Gs9kK3p0HTB2TdkdXONIw8UTky0Hw+mPVCMuOVIUgnQYkcqfl
OG4tK0+AYJ2q3Sq3T9B1JX9a1Yi7peFS18jb5Di9iR4EMmLeiqnx1jGRhzWS
IVIABLDlSgtg4p0dBgsukOD4kFsaS/LEhzmXKZ6T4KfLEYEo5ISAPrhfps5A
jYfmpkZ5q6h+PWCpVF48S0i55zR790JCmkGFWij3wTK1N5ooX46vWyEAW2IG
kEROT+KevL2PXigCkw1yLvtcxad2SV/k5p3FJfbAx5u8pcrUDs1SB9qABCzG
hNYUuohgVvqbr8q0dc4RYbbph+F7VPJJ/00nnRGZ4f7BJcCdWDK+M0k1OBuA
iU7HC44wIn1zNGNSsdt1xLkUYpot+fi9o13vqb15yfhyvDZZ3kRBLcwM3xKl
7fzWRqA856uuPOgj49HAODQVy+orZdlMpmaLUOSRpTBN6MaIq+DuYgzOD8wz
IuHGFjlkL/KAHDD+4C3iI2pgWw/r9Fxf3A==

`pragma protect end_protected
