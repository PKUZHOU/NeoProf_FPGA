// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
EpOaP1i8Yx1c7wY0ncMYFq5iJ7PqtSvGwJZY0VVQto7gHmmoCzLnD4g3G+3K
a9kHqO8EngK2T8R+H3nL0ICBj4rmYmm0npHS4gS8hKehJ5pZ7niH12v9TRY5
qiac5lRo8D5VKEuW71mpUJ+RoPJlWA2pn6SM18zl8IPo9NE2pfIsQ9La8tQv
i2V/XjHH6AtQP6NsqjwVCMGO4wxM+pEnee3u1Etyz2+uolSpxqTXTuDdRD7M
P0N/VUjCTjE1xJPASWUA43tnEUK0sqHgB8JhAe3E9mS6Yaisgfyzu07g3e32
ZXeyZbPOONWnLY367ACvRvhyoUHJg5fjgigDKn6+hw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
cK28QUdG49NECZXgb6+hkrt568RoIp7nXxxWvkhMX7suDx1qSP5rnmyTKj7T
v/8fPyFY5TVaRD5Vr6eyWT4Qo3RbKs7VaiO0hwdUKm0F+TomyMAo4ZNTJhNU
h5rUirTLxJytXJfJDGQlOM0RbMmPj3U41k+brU/PqQK/l04TOxEVryfcQ9V6
T6Pa/zPCYq+qw8Sb4i4jwK7j7nOa0np9xUPqdPk/Zjy7f+1AwcjBahm4hKNI
R0VfM2YBoF2X/fEaEQiCf6Fm11jbNApTbIhprdCP8qNv7+yKQFscEeUnKVHH
dSNgnAL/jNwtw034Tjjo43KITuR2dUW5ABzL93IUFQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
QC/iyi75TTsDGPKeuTO0kEx5f7ouZmzejpbHv6Wy/9hbJPN4nKa7yieuYXAA
9kPNJzgxhY4tfQW4xr/IcUZi5x5LM+J4lc39yP93niJK5WCAcylphJQMlKV5
kDFPdcooiwFLY1RvPYeeFhCYjkeXXdqA2jMekg4m4RDmnJHGfCgzN1TrGHYC
mw3Y2cz7qc8r8kfwAlCEUcNUnFeFz43O68tq12iT33B+VZBri2Oj7gF2+YxO
Cgwjw6r8EgDNiM0vDFQp2kvruZSA03kKh1YIyvYsudUR6CSIMFBgjGzrfoBN
QiMwZw6VVlAxQfi5o2AqN6iBY/6sqzpsNAUklOhiEA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
BAdP8sfNmUeQ1l0g7+CrHAwxOZ/WjxF1m13kPdqMNK54+SkUVhM7XoBfJdDz
ijj6/fo4t4bu7EUCbi0FRPV83WzgSVW7Gb0SmXMmAYngxg1GGegI86UoTK6g
3RTu/ls5HYIdHXoWgNUpegApyTk8wyil4KAgsp7P5N3LOaA7QJQ=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
hi4RwiWaEaALTKqSDaOZPN8ttAYNY1MoWdnugrGxMN5Zp3ToSen7Ncq/ZDNj
aD19TB1e2FaNQvth6Mvs7CxYHS9Z9oxbsPi5j5vUEOQXJve2dzj/TVVkYCDG
jfr+WVtumEkerMvwyrwIjW8b/wdnISpfsBpILc2HDTiGXb8k7wDS94uzImiX
ArnweLgKX53tvUOD1DxBNFKfG5irlTo4TfTKsjIb+SJT4iVlGqhg9NWMOkOc
VI5nOLozr8plRHnys6hE2J1sgtVaf+XEu6khpEbG04Uq7uCuzW2la6CwAKR3
bTgJSCfFWOvL0qiKEYAWsitXishKNA73L5BEgz4XTNwTvV7noGPHWtQOv5CG
3v6w0muRgxfaBWhLjQ50PplAArhbMwUGRQ0K05WGa9GpRCIsn6/3zZhvIEAj
8Begwt6Uy935CeAEa9Lv2Zr4GIJsriWutVVhxKSfjSES3RHvPdvn8QxIV8TA
LzCyI+04qDoJthXO2F7cZLRieWxFmY6e


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
adzw4RxoIyxJZuy+CdQZwbiH/2mVTcPmeBHCLSO0yzoQeR/2ZorKeceThITK
oHGjmKr3uxFpqxucZeEn9yNMloObhTY4zaNu5frai1+jU5UUH8QkGzg5eeBt
vUkAVxpG+73b0oDXQzfqzCB7bv7AVJgsOmHW2OZbSL5MEeVSB3Q=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
cM721wjVjkE6Y4JtuluHfGikRP6CTWJ9TX6m436qC1AR0YnS9h5ZJgEznhwB
f22rRxubVXT0U+C7u0C05AriYLewSm+aqx+kaL1tg4e3tjJ2gbANI9WFgM2J
hPtNchiJqhX46u7nn7+BYOhYE3rvulC63l69nJC7f5DKB7u+F/Q=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 3296)
`pragma protect data_block
SsJqmwRXDcQfZqOU8GG05yXBdRG+pZNWICiScXu40IndkscsEnPLwkj+BUyr
5B7NRIuPtXJ4EQe3drJIMDSna8oh1UUTqk84GYm5z28F3me0tIsoKaESHfe3
VyBC1zFYZsQDumzUORvJfxKkabrZpOVGlrt9EYtVmM0EmbVQ/bFDGVEi8+JD
YKJnT864jUcgIEjMHJWpSp6yUrvgRXsoNHEcAYGA/Pcwtk4ZlKmEGuisOClF
8BJXzB0IINhEANpPPRbMicSWfjpelcUD11sjycYp9sHzM/y9/Ht6zIj7J9AO
m75rA2N1jNuob7jSVWloU43ndTmT06ZCiUYuwLq8S0HnjerFeXSFkNc23bX6
v2+Ftbf69UI4nDHJVXdN8zed5mmkZV5BVZoNiuvzJDbsD1PbG+x6Wt6jbV74
hMej+oLTq+HuiW07P15FeSHTI+13dSAZmSlLkSer6R3Obn79OvHEBTB0fNyl
PPdrSdQ0ZuFAzqgUggNXxa04CtAV02POqJvf8H9NM3yu6WhuQaNxPE5Q7m/r
hEK0CQtKZardBSYf0zeMIgbfJf083GmljEMUkirNkDwOChr+w54Hjk8fk9Un
JPghdt16VVb5knPfEdXUvVMesFcVMx+rw/4DOKuAK/VGt3xoEU0Y1NzeDn5v
9AcKMHRrYaczIuYObpKR+Vrsb+E6UGwjSjA+pNWnerI1EhIhfa2i+6GlOwMl
0krU8qvRIf423LoswRRANYb2lREEFSolpIC62rpv406J/5LEJvHDcxo1yZEj
TBwuEnk2aEOoIf7amAFTDU2kMzTleEwqlSavMWzk+BPzG0p3w+MxU1P52qgQ
uM17eYrzXt2a+daTVKs2SpM4JE9SQ8rMX8Qa+FopBPF63YRfJCm8Wdto0aF7
yPD4A4P6pvjWQds3Do6a/3MIBQmBfu0Z6G+npNybuzENctYa4wDbsOzbXYbe
EkayAl6TXQ9vfbQY8BpT0HQt0bnUo5YiCvQ1NkYJQdl3eScc0sVwncYc+U7A
tAPgtz11eaGNxdqG1eIpu1JnTqK2NnMnJqb8kjzeKmpU5E7yJOC4EPBYfN0a
/qZIkWJslr98GB+TCOfS3BgCk93qmoltf1IkmNz78IbeAiFIqcJq2UkDUZGy
KwOBi0MIgh9vNKOAw4OGqYl5GHUd1lNdqhawRPKN3jBzejojmQ/tU6ZRJNgL
zD6YiQKndujGfDBrwJMaveQz1zJTQ/ilUpL28qq9MFOkntUpW2O0C2llRKGF
Vm88bxAecqnAKrWvAz0lk9nAqsTdRotMvVcPni6y0hYfEOWMdEmIiE5DVIsA
ei+HILSknK+aAohZgoaCT+sqaHLWgtcMj2k2ZuZ08eU5JYNgm2elKSkiUDUo
Yx33hjFnzZEkvkaRXm+QdMKSoiwDFxZCFo8FMB33pkkLGE8bjyUhhAIGxxwN
wQivYN6y3C7UJSSyvYf6r0832iOihmG0CS4NC2HYWOzapTqtzH4R67ZNnxak
Jk30RBQv/evty4ffWwuxGW3FHHmj0g9lb8RPTHlI9Z1OttgzxVbsxnfgE/Rc
ucRX1QTTBshAFZre+NBM9NO1sj8nZIunGUoujcxl9yP8GZ6aptYj0pX1agQw
CVUkPv/RAcf/ThDcuk39qhP3fMUyLp7tLRHG+x/d68mwImygBHKTsrBrX81j
QfSMfA4T+1P2ZVSdJvui8t7/KYNzWi0DNuEzE+XByR/3QSW5seMXmB2gzd+p
gThKHoevNfTv2A2RJ5OUbs2P6kCethdq9YEzNBUAHXVNqaLCAA4VG17b/qmv
h+K9RtkczqJbFt7eyNlO+x2AHS4AvHxYF7K9Uq9sxtaauvmk0xWhqVsQ3QIm
qaTZOG/+ZnIbYZH2hR6VYaEMPD6IyN20cPVXotT535pmQmY3ijnY7kinf2x0
bAYHPVnkxoFiXGHbVpLjgrEI/zlldnupKpTey3kVhIMBzewtFUL79bINwwaV
t4Liqak1Aw3tiZPQ7xW5atiBP7gHIYZh+X5v0BezIX21H9fZz0IHdKgP+JCL
d4y1C1+6/np5g4tZWzor2ZhESWob15WzhFK6Mv7jcforVjt7nBN3tyUNhkiB
vpXrZl2nH/Euw0im2N3XJI9jWsdXgPcWHan1R8idLDq1cznr0sHNWTze+RKA
9KaLamAYfzVN1cZWYigP5pH0qlcJ2OB8tvws22DT7aU39oM7wyx3Z0IkBoz9
qTXswzOYirSjnjJMaL7yzVCz6uPOfFJyK0fDBch9spi+aInm3W655iidocfl
CvHhK7azLNQ+u5/rn9b4wpjOLCXvCCp5X2LKDp50ThMsrZRRG7GoTBfxlcEY
wq1c2RhtqIkpFuv3Y2sWp5ml2eM9+DOvlMAkRuurha45utgIaqnFJCCMA8MZ
C/WZ4MgW7ro/nCowRvnUGPCNIYlKHCk3/ouixm5RsUyigz/PPJ0gYHgPe7CM
ehlw1En7hO80DeKbrbHoJErLUulpBUvr0p65fPShHpn3pOTvaHRxtsBUlmD2
ijJ5nXRznBuF3wyMbsSSQGzmJkuYuufKmdOgdJ4JbHqVWV1Fyer5HHaxINFt
Af1EDp+aT0mD9nCLHe9a4OcOoE87b+7unvCCi94HcsmhF4KXO1hXi6r3PaFd
0qD6nlPy37/b/CIPl0U2IJ7isUVJ3vbIVht5mA71IGFfAZQStLVYEWZeWtuN
Dn3W6YQJXZly+Xe3GsokeURNQgojpWScdNw8Rf10GfIwKtbwcZayIajOxTIh
u6NptpDKpnsM0jD1JMmw8SDP/hwsBXFjDVq9rKIv1QwgUOjJG085hMV4y7Qi
bHhJFR55wyd2YCy439IqGtXzXx1Abuz5W8v1U6EHi8Xwrw0JKFS3TjXYr4o3
nnzgijgzYb8/55UmJRuaBkxsHWSyLFepLZVAL5QydpAokS0UV2r3L0HnNFv0
7NjflZg31NIzE7NGv9jBFf42WcMVWifK12x9Ysf9J5jnZaXyGL0nQVhi5xXe
7Ga3hrN9QyZyXd7C+vA/kBu/oDbjbzsGUsjrhs1A81nmonxMHhET6TwDdD5P
UApdXR0HKYxYXZIrEvTsotHKfsbn1KzgM7yIEo1b1jbXTwI8o2yrCcaf2OLx
U/erA0yXIxmk8jZAATkFTb3vparC2604NZZARDgyDyFg86XoEhk1FN3xwaXQ
tjV1vyr8poCdaHMzt9x4IttLoh9pI55N02rUuOlFmmod+8mqARbyvPI7H9MU
8dMXmPqVG1UeLKyg1j7e4NSr5P+uZyxdENdqiydHw/22okjobmpHiy38f0T5
9STxJyPlHpARyYftGC5iSrYLYFzW+snJAXV/K69yQQE/t5aceJdijaE9w6qM
HKGcEE3qaTvS7b1n03VwrUCFJRcTovLeMhGDG59hUbF+8ssxgzwex5nSc7uE
fmObpMzjayPxuFv7wyWUSX6vpEuBmONX1WJr5d+RhVN560LZtup96VT3wQ5z
LEnMsi3DYFk1q75l2fRpi+4dsiwBjMNsZiAr431ImvdtGx8yds3CUN6f+uZ8
f/O7STkVKeUnmSZjfnAYXDg9023ELfWZbMSJ03ec1LCVLjnUPJ2Rse+E+RSo
Im40VDe5xsI3e3YOqvgkOl85yhqYn7Wkl3EtAaFENow6sN57dChgOCsxje7R
njipsK0f7GbI8mdQrXUS+gcLeOnKPLEhhrAAAQwjl/MPGIe4CatfJO9dN6JC
YYF/oCm8W6pvpImFZ3xuvkXYeMxUe3AUc/wZCSfRzY/+yZVQwXxvVt5v2nuz
kajLBqzCmoJTbxFNBRqY4Zv0h6rs8EgBdSew9hkagxPq2S8bBW9wRpA+dnF1
IFGf9dgj+5rVLaavym0d2tcivCcELnREljd6j560KkIiDmG62coGZ+8oiJL/
Fi0RupcvheY9kKXQLK2r1vHqY/0mjyk5ZqqOXBL6CLi8gGd+/JCsFaFYnLFk
XHGgZA6f7U8HQZbfEz9OtLYa3zsi+SypYT7Sn3kKHZTb2VN0ShMJuAAHp0wb
kMSN6uHKfp5mscoDX4zwfPAffsdVgQ1P9u56gBSBR5d4HsSZjSafcis2Cxb3
oKnAiwWMvf0qsoMkGEZ79F2T2g7GCfTz6XOESRXrb1mBhpbcHVWt4ap95QI9
PnZWcHbozVKXWGnLXmTupwpLGDRI4JJeq5i2ChnmzYTjyaicwFtxfj8ByDRX
i1shDatiq3vA/vVcH8h3N/u3jWUe/isO17i2iJFxwyt896u3NqRtLFBW6t8S
LZbpoZ6tF3mwY/pIIkprPyVV+H/tEgGKLbV2k/Bov6KVFstGZ7gZ3OqjCEJF
1A3hsGeE975kqRK+dJa9INWHlK3xEceJaq5VEGZoAsnKCxVd4OzRK8VfXVHm
8eQ47uEq9wPAdQc=

`pragma protect end_protected
