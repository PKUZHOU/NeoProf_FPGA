// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
vudVNOVCxpkUEwWQeIwR+EDAv5bZ04aMxRUtDDQRp1TEZrntB0tb6sgX75eGGlE5
3prEXnE+7p+GlJ6SI0w3q4keLIV3J1CuxddXDcjGyOHu0Asj65jsbYPGlsfIKfk/
e2L3wFqeFPWKcUK43eWF8Vb52WWTQ6YlYDPfTyY1EcpYO6Ai56GFeQ==
//pragma protect end_key_block
//pragma protect digest_block
E4Gyg2YixgLeNJJZULxG3HftWaA=
//pragma protect end_digest_block
//pragma protect data_block
lrH3vgTcNR5AnkB8526YZVc8EXusNcE7DZt5/3WQDcJ2TnCAN5LjdTbtOYTbnz2w
N7FBI3CjWiCNFH6otnGAsntwpqYBfBmJY6HcJ6f/T4eyesYDtRphCrTLU52nazWN
CLiau8r8z8lVEd+uHY45vNjgpp2XkpkyFUY8KiW42Sa811zXHOLiMj5cYsoq4vHn
MppErsm5awSC5dV20BEM9eGnHuP8JGsFfqrNemYYIWv3KFBqMq6o01yZ6zFWdFXH
O7Y+PQY54pkTvjcAJT8b38d68/LqySCeIRkFkyXUviCvmAWVa4wW7t0PYpOpWhad
FfYMuroidEWsVwuV3H4gGj7RomzHXcl6nM6Jh0QGt2V1Oh8dfU9Gf3J/DEgEQHSP
vrkg5+EfynKa67gis04/kYCp5lthaWmJXla5cKnn64e8HJ/dzQAu56csC7jMPcuq
hfHJNiJstWEABWm94CcD+rg2sTlXVCy8Jht63IfFnBiyrH4FHhXdHUGYSx2/N+nS
UrNLwx8WLnSFBtPUKp0I0xVLdGERln6ixrj9zP9dmU7w/HFO84/vsSwepnzLT5YY
/l4H37Eh10dCHNf58lx3Kw4P8+YC04pMBMpaF0lZ4AYp6dR7459lGTaHi08Bd/rh
opMdp16GqVw0m5VncVAzIR7YhCIZsK6mOcOT3TbFb3HUxFPqKeNQ4pxlja98C329
xLLLbKDyezvSgjgCbgk/fwV7rjoEx+dPq7v5rg/cBJ5ZceEBMp9TMh7ZBU3I9AvS
mPC2WbxneOA15O/FPC4tLDI7wubPLKadMHvphbob8ht/i07T0SXF2XNPkA9rQLb0
Wo/7TkM70Sut9anSJkpmRHb3CAzgioQxdAmYpKraA9k3U/3aENoaAdsjdHftqlOX
zuFSGLX7vi89Hu8Asaq+i/TVhq0InRrpEZV1nTz60+a9kZ5JLOpRDMnPxMmn9uUw
H4EgQT6RwALj+wRw55/Y4/3cPP7cpIr84I60ZomuYDN/+oTqaCRO3GAFwglQjhZu
YTqfZRrYKoYlNsX4NrmO0LdnXaBFpyfIZI+6VGXnZBNK4qERhotLAfQ4XfG474Tc
znIXmwF00si6oVdJWliXjD3cLGn6GKRHmLcDa8hbUdA/fDPET9RbymYcApTlNCXf
7mTCscECXZUaaYuiL/6MFAxozLWh3XQ4v1Md0Rr/EC6miTlX/NQ/qZOxD8Abxcz4
i7KNTL0VBiR0SIw6wpHW+j3u1RIrI+W1u0Ar185k/gstynaPuRSOmrBQisgiqzy2
8wzhY8Qxu21ImZpCO/ags7Un8pgAaBWChxsvteBb9SpnmAqFwkTSoy6OYlmMOn24
nno5uzJ6XqNLIvgmFXLolxqrzfOuAQFCOSnIXTVEpJGBBoc+Gg1tZmmLyaozMIuT
kz5B/IQ7XBKYfYAFJ9jsmtBYjOWOp2LG356PQlAPGLbzfOZliiOCbTqrhUG9sA92
d9P/mPkIZ4b8n1hQnTvwmqSZFLz4//1B9yjJDbkRu6EUYJvBBPeHPmoeV/qHelI3
9NaC8TVOZCNHzanMR41AdGCBWQhFPJP8DfDernAL3mLgSYHdjjPRjqwnqFFnZKf5
woEHLwjYT65ABKGPCFoaNZW4PvhhVa+jpEIf2XuhPHe+Oh9u2m6iOMomTDf5N8SY
9Lt53NVLe+hC0ywfajUJTeTscUJTGVZqB/TYfMbKB3FW8L1b2sJihttXn6b9LVfQ
XoDw0fA8t++hzQ1D5jYrrmy0dVWsj+6zniIM1KPKNadz6QnZ4HhqU9Azls1kcWtE
w815NVvBHtiZgktNHCA1oCQdu03591XJVma08dDzNdtx6Inrzbbtv6DzeRcofgba
W30abOZC5fbmMb32eUQQT+HFJsLmLhU/xlTVmS6c18CSYCnoWB/zoTFwGMjiGQ7Q
dMzLSE05aJk3+R5RZDC8yfx1fzxnvqX5aaDmqmDm1uWl+DV6+H/334/X2iAh3/Uj
yJiONBxtsCWGMKtTCkT74sY66IJByC2Le/tuLhMfSqb8y+Mn1YGsmaSrA62Y1aoO
0q9/ILNrqHTP7Lh3ari2MhkwiVUES6uCnQuzIESB015ZixbyvIzXlCqIiGQI8RjP
FKVmZPALo/5pacxXwSp8z/4jZqcsPm2HNL+tkli+3M+d6Q5P5bFxSx36BRv0kj5Y
H7VIC6dZaP4+gYmfcUlFbo67NxFIiFadQvCeo07LcUa56CExW8D7U4yOeaGW9hoL
Ko/DnpwqjKuzXAZk4mNtre9ESRwgx+olWUmX0HKUZfQyPB0K95IIB1E907vnpbQP
QjtKZQq0yEEgjBJOaY2mw5H8opGTNcXAwtnuhRR4VcclDtprEbDvgPRbbkgdnbYM
QJVA1GAcoSh/xTg2sA9I6QRFi1eULRS/EK17jXXRaH7PVqFcXzC60JIiORK4t4mK
0ybn43Dd8RspRmEhaHqk6zBpSdMarHO8G7AUr/7pBcA1v8oJH48jTglkMcNPaxyH
SnNhPwhxhYdQDMALNBirRIisF7sCAWfFbQ44+SWBJaRN0Bv5f/zots9IwuIipKR1
Rfl+yTbgUY/L9E+tKBeSzYhd0w/kOGYI3wkX6g8UYpQfsaugILhDXY7bleT5GsJP
vmwL5VayMrgZ/s4m5mj/1mpaXvrVz8p7nweI4EMviD0yOPuxCd2x835kLbr/lLCL
+hRZ3vpH0wx0kJ0tYLHQcG0G2/ewo25Ia2W5QkM09yi5MFU+v69WYUpj3OInqEYw
+6U7eoTfbdPk+Xs77qy4V8/ZtJKnpIz3qEBqsEw4H6pRcnFaqGpGskFfpITdk/d6
fizsX6K8uEdMO1z0VPMjQ+qjqfmVsfcJSRxM1cGdADlF9AtTFbCXiuB73FG6R7cU
nVkQ8DBAnhwLyzHo5sZCBOtiaY0IhZWJlq9XA41G0XP29H+wE2JV3uHj4FjpaQgn
WGcLGUn6maRY7cXWwIMTIJFsaQkKvmNF4reuk6dsRyoocANJ/des03dnVZ+9Vn5R
wL76YWxO/DpIU1RR+MjXce/LE1GkfB7kDySis+BPybcTGrw6c920XT+8wEdmEPcW
DYMQvG/A/8cjx+G44gJua6BRO21NhIDxWRBrSWm8QdJq7/04s/Ro5gWhj+WTwNmA
woCQq3DtumwbBeA6ktdNz8R1ICVM321ExY1rMBExvhtYbxKHvJ23v1KBEVdmfr2V
oStnguVjXm9kwiz2KKLnzyNjVjYrw2n7fKEuqVYvfmWMTZhQHFmAkFio4b2t1o3o
FJXxczXsxSowGo9t0ayUxrUcbgcRmbq9EKZqBJD/Botl67hnPY8j7503dhzuyYZM
CklHC3PyUhs07LmDFuayIcbzdXPvUno9cjPdUY7cFPVFANRW2eNiytTIgTX+5KXv
H1s69sP8EaYFiNwJ8J1zDlStQuT6ci0hVsQuaJY90xhwHynr4v/sQZG8cK9G7od3
dJE5uhXH6SgKpgn+//8kHS4QDo+KqwCtK+NbXioyWDFCAC5HH35LIduGOvXQWGpH
JZkHq9xkvU6d6BM6begtuY+j6qVfOnd72y94CHRQ/bpLQYjd7YgWMTXykB7uhtAx
s+27m6Kr00bPwKoLkTLv+4wfiXS+Au1QUGuSnjpOFO6ymE5/PoPHylRi+x7MZ2j6
QdOxO5Wbdei2pl6Ptx8HrYCF4gqveZyA+r9qpZNps60cn/Nz3QEyK+5FI5anmvqc
7V+OdDo6axd/u6NJ28eYGTHDXXDEp0jFbJQPd8rL1BXVpU895nExIl33yCdqo5sq
24LTCJmzmb4J76L5RvpSuylQ38Ym9ynwaSNHlHsArVaG/aaDUM8026SBcmoXN1JL
WKt9JVU/80HLK0maP1KjqoK5LV+r9CEJkDmK3J+4j6/1rKHCAHhafreEnTN0yKuQ
wBzwgZYlR2xp3KOVNUkglWDITe3GOH7nMNkuwUp1HgfxUXcZipG15C5myIMuYv37
p5WahE074qEEfj10vyaTq8e6eTscqSMstgHMmSOaO5jZ9yn4hus1HGyeOkY8bJhx
7yWXrIOepA68rQXrM/60JhZ3h8inyi1ZAYQkhqjbZz1g8ymfAX3k2YCpBZ5Pylxp
OvAD/6DOW4Z0BB+RhJHbIsSkn7wNgsrrz/whDzEctvLgJEZhAGhmgYTXu7bChX8t
9IR4ap2Uro9bLPSC9DBbbGq+g/IR7NMMLZSPMh0ny9y2DwHXQXlGefo+tGSfTrDY
RuIlmEwfJs9CsjHfRxjiaHqOjdYs/NUTWDooRU9/+0zlrEZyPvWJ2t31/47q1cuP
H5yKKegHdw9ZEvuwnflAQO736GGBnUrrbYmA3BdVdBNvm5hQdsQIcB5YeXDRgRx4
RmZS8xu+SbhgnhiYEn7fdBfSM2bA2pxotqwtxBdiucxdvYDcu/hs2Tafeefg41HB
P0OOU9BNGRVa060tpZ+wna0I+PgNODJb9GtRiso+Cb7GgkS6U1n05Cz5Q8Tv2TvL
aRi4+efxoY+RMP39GzbOuWBrxUf/tpSAZWaj1N4XVZb7Hg/wLMilxUkduPRKgGAM
LnCddtaJhSJw5hzIerHu0kPOOSoowTPjN3tN/iR5Whw8j0xIdVeUXcFkzfIDsD/L
oN7SF3jtJJbGJY86a5SzY0gVtLv6AsyJukkApUDwZPJJmCA5q14JAkvYGLGqw/VJ
iJrWrJ9jQsRtFK6GADdgDrZ5faSfdoLLJv75IBl0J2TSnCsABFENAoOnvL6XZMmV
aCmkEzOvh74FI7Ga4vvwYI8805AYcnj5xKxU4EPQpmUEII41cAmIwrEEI6hpRmHb
G1Nv/bL//W63f15hRBgKxhFcwMAI4mKU7RI16kp0xsWpbSVqN7oTSZZ4UA3sIyt+
bSz2nG2/xf8rqmRovaTz+EISY0o0N/nmqrn27vt1YGn0x7y36g+n5oXru74z1wD/
PYPuFvPHQxC9Th2cBTKCCo/yqxBMW2+E+LNhiQZGoudPzfs+tVjCvkPW/Gb9DnIQ
zTRAEHG/92zdhXYDv3YkMvP6ohjoYcC3cZJKJ27td6TItVLsDCOlJRbyPnUhoEZt
U8KSGvhMLw6clMJW60ME+i+IUc2rgBbizYOkAKA6HYr3R0OdlKtj4HMMOLZ7Kab4
sk2K43JG4lfkmcFKNvw4Y6kPMSf4nuXcGAFy75V0xvmAG938CPChIXCxvrXhk7jq
HjvIXghebABTnV7Bs1Ak22UiOXo2IqVpp18OTuLYnsvT1q0VyMbujZPlpdDOhHuz
5SC0JZSSnoCyZZeoGGlXbc1Jb47u4F8VQUMse1ep+zE9ZsAyZXhpfNskMxPssrX6
JRCe9EgCJ5unDEoCDzCfpLsiTwEvaadkdnXMeBUzuk6+3xvZGL/n08hfNIlRfnnM
96K/Tu74eCJVV5GGsKaTIVqNGAz0syxy+Wh2tllbiPB74VSkX/N4kCcW4xI37kaa
O4xSYFlsTskcDbrAjjGBJC+BEORkURiUXRkncTvP1YsYTzjkLWiluZ3BbfKYFa+C
NE/0XLF6d48wyIzFT/05qXJJV6QCyTv/SthqPlK/XmFexJ1yszIj4eiMcxZGYoSl
WARI3LwbbgMfCCqndPI8O3kR6d+VwCNvArlMOWnP6U/UV4fMmXN1NfzRlup4PtvX
SY8Xhlaz/ruvaeiuCqRaKaXPp5FYS3UA0FINdhKOW41IFIwQU0NgagdnbvYDDj4b
2HH+JqMfcK3XlEdhG9msyQBVmDw3INFlfR+SR4rdjejtecHogESq7K3I7fMIdC2I
k6Iy++pavRecD3b1r8wyKwoBcUqQEFQHNg9jBzcnBtQfWWObDYp1stKCWDsv6NPF
Nj/Me7qakGIFjOTCwI7pCPMYtmK8cYbI85WvY7K5CASFizpGdASZlisZBiBBZnmZ
K8xQDhDqCACm6qmBPKgxv3LYIEq4k37XyDLAtMq0QecIdLbpBsrPYAYXUAALUyXV
zdzVtNdo0u2530A+2mAfrcUZC1B6aU16vgAtvCNO2Bbjdp/FnLrmHZaqlKqiazNp
B/8w9avVVg2kCKSnpN6Nyu85suLNtXnFjh+3mscyqAvMmCTww3a+V8iHwI7idKyJ
8D1TT+DnoK0YmvMVPqpjj/xtlmEIZs5FWSSjo4BswpoUqyHdISmIxlRo4Ri8Ey7d
PBLJluPGIYBjYtRhT6XgxptI5qaQnjjzJY1jqyUVb+YILjcBMcHKkNs+t7dUIKwx
MKKPbjvYCjnkGAn0QjaIqlAXKRsm2Oc+akmeav1VBK1MZY2xdDuRGbfp/+W2a/Ob
S64ZoLkVSTAhDzysY6uX/kBxmptDbqJc5C9V/CiODz+tZaOXIfzhtU5cOB2yOs0D
6Qssra4n+15D7s48Sao8tflniizgSCpXv06dCB3Aied1pT5UT6VQYxFBFMdezI7E
4YVCrlKOzrrBN7urFGjicbeawVdUoQPFSlGtH4yAZB2e2qHJcR389EtemSnvw55c
r3WElpdmEqCCajtOGPT7gd1Ez57ncUCBzjErYbtEJ96hR6yZf3nF5QqSg00GMOzY
IXtZUTOIaJ06i+YoooqpR28sBa3rybNZy3Zgy+N4O4ATabsg8lUiwCNBEJdBAy5u
zQLxYoh9DuSmxnP9FsG7jnuo74pTbB7TfcmDtaslj0ogeJ2u9bc++c4ZgsKZIanP
8Kx5WXPDQK6JJlaWNf86127dSkZJdJ3M8COps9elCK3oCIqH1iSKYsJVNF7MbfJB
ApajZm3t9PhjHIhnQScTCUm7M40LDBO0sjZEhraFypZMW3+x3sizmXAHQ/nzlHIA
oSh2hVye1OgrP1qEvkQGZbJzsFC34FtV24gXl0njlT9zukDrmJ+zFVfaDPIl7nB9
iEzv0JfkD15Vd4N1svDAQ+Rs9p8wpfMq4k7WF8mFLtiUsUUOFFtE6rdVTTfSi95r
od0Kfp+gIBYSy9RGt6H00SgXNhMmr53jVxXcEpBqCMchkRJn06YRkMkKzUFPkWAM
G74AKnhi2jaUrtQh24S+xrhVm+Oy10vZ+x+6hE3KXSFmpZgQSGDGpGwVdEWHzJVU
hIsdW4C721CaPKOuqQwPAWR+FRTikLS6hjnXwbOzFsOz+0CzTf8xiTWQbGX0JZod
XdiHb85YXX0iigME50fPGT9BPOOoL6Epj2RZyWkB+W4jVm+uK1PoPnPZ11zRV3vk
eEO73QjKEBJFm47kwxCCo/7z4a2w9xJrj2Wf2+/+3skg4TemkVp0e4yvLRuLni1v
MTNykN14+ySTCpXATssr50CZ9/7ZTGxmHWhqfmi570mmDsN7lDRjaQGW7Km1wbSq
FoBQMaWQPuDBOI3nbUpiwmkJbRJDIyitqdtt8CvnmUHbW6MY2qsksJx1kjtaaudU
uivoyD5tRggeZmnDST/kBb4jLqaw1SVGKccRr94N/9+mruf7ZI7YLWPSyMKGmrXL
p6A7KZV4SuDr5p37mP53YMfpx7DEmFPxtk/Z4KulF8ONferK8xxIvubIeWPybEVa
/csjxWevSfh5o4GduypSllfEVC43k9RXAAQ4P4bc3/66bDBmzTbpSbSFaDsPAr8h
JRjT342uDKtOSDk0ZnZpke+d5DeW0LYGynHC8rmSWMYFhhkLsqagmZo/HEjOn0Xt
uFZU2/imEjd755DtmiSoAAS00kFAZX221wsOldDsbWI7SvPatpW5ELrZp4PkHCyy
fmD8l4PUXlOH6/ldPewxXhVxQIQ0Zy+KE6QWlmxoZTW/fFTJYgTYvSm3p+4355AH
1SFwWKtq6VwQ796xSjBA7mm3Rt4buc2YkEPcabnhwsxM+8Gur4NYpnjmAqztvxA7
a3SXlYPtBvcJ6qZ9ZvesT/dez9Zrm9Csz22vIr8yLd0wgvgFeJeVxZxB7BblNnze
XYd4WulVXCjhJR7f+BSE+r7f0cMGLLQYzYUf0vO/bFJ234RzWkwUo5j/NMmWgzV0
L3EIVyj8G7XJB8z9UHGqAUAEPfIxIMfK0tTq9PBh5MEEGTsehhEXK4yPi+c+H8Ri
b/Sqr6SYOmw00LCQnd49UtSaznIbBfSxlhEh5/mGzspPqdDRwFeQkT72ECUK20Pv
lgg/P4P96TkXUjgD6CzrA4lrYlfIhhM7OdX5obP5SdVm+FwRMw/p/F76rIz3snWM
PzI0YeRAUR3hGlH3GYDz831tfHmOI9+qmWuvAy9oOykHn+CuSoJf719LoyDUjgR9
85lorf8+4vNEsqsC5YVdbhNWbW56Gpgjd5cBh2IJJTZnAP0q2J3AzakbZIcJcLHR
07wqVeokJHRwsp/qUMrFxkpmwOdPBVo76ipVmwUtd3lFz9sdgVGBW29i9H/Q62nW
/vMM3zKAH4+1kFh8rsfNnrxCQ3QszL1N9iQqf3SsLe/E5nwZSnMPCW/1NpK2cwDA
/5BxlwXzqiYG06Iqly55Lgf8hQUeM6klkfmknCK0/B7UK1NisdgXuiEagxqaAD75
U7qkV6kmgGruSEm5tUL44OAyCswoKNYrXGD1oBcpvrp/yP+g30Vj78emxBSItH56
/yxVJjGhcbSGBT6yUvIvRzZdABv2uKK47RLiHzYj38GDY1L1PBPvdCsPHk6nE/c+
HxXOvJovUec24Ds/JkZvIWAoXfuJojNsScbLNc4w14CMW53PiRycPRMUEBLc4nO5
EHFg9mTFYGqjEYe6HEhkNtuY8gHmNiFPoVuJqU7xnt+g/YnhtYUDDeI6a551cKpH
3PY/cxkTj7yknl7lhRxD5CzzdcEEnrxu7a2TGOtXIWqNsXorOAGgVn6EO8GfjRBt
yP/T5yPd7CHH36uJCI9qYV8/h38Am8OdUU8QzW+a0ehwiOSfMDG0yTbhBXOBG486
oGIyYSZv8Y70QITs0X2b03RxJg2gXnkf1gF4NyPEdhj72c2gC2nhSxyl6fTgeFuV
wmGE3mdGwmura9JWp66FbYt1u4MhqEUymllu8n/xeyaAEJ1Emrk7qNisBUAgrKFF
/Dl0U9Bq3iSwbADswAxbQOP6ug5EjzlxKL9xzW7Azngf7sfr5HAyysDYZaoAUsA7
/lqjJB42mes4prnb/oN7zjf3yO0g2LCLX2bTUfCNl8dgdcl7l2GKNR7oVS1gm7gW
BCJrJxJJmPcizSd9UB4FsEzJH0L/I3xzYG77I2XPvErKxhUyfYV5yKb8adju2OiJ
bWpwouCcNtkNayKLmfD9rXkY7oEgE1ZlOlB/9BviQtDhdcPaeM5eUR8fi2zf5tzQ
ului67T2Tpb6KuHEttUUlXLVl9eQ8W+EHw0SfNJ8ikod0TPtH6LeS7GtjmgG6jLx
PlY4YkG7lrNqXXEhD7bCeEPXj19hhS8a56fIj58Spt8WHpR+0L0NXPune5Ek5Twa
Xnq5dkccJOh82reR/fU8zDmJQdB4aZAXfmU2tfF9tryRtaFmPOdT1VD1WccYxMWB
m8O82eNjof8Jxd8zH6VKS4+kjO6Phgd9/gOxzyfQRa3iKTgml+i7rJdBwbUAbfSE
XbAbm6vJa8t1dQNfwmeKyzvV3v1FHQ6nDeqpR2QM1/RewJY/sDhVtXWCRm4boMal
yv8/MvEDfYX9Ac4pS4Iq7rcxtpf9dPlVoFJ+QBMU12x3IbxbMD00D/sWZeB0aRYX
0nULNZ33crwCEnVXPU3hZSUYx5Z9ctT526Jtd/Y4Mv6hDlENhMFtAYuscDpvqjRR
lDi5e4dhpQOXMoc8YfKPDjnUyAOlxvI7eztgPYLU4niUd3kZ0WXJZxzLqnFliAjH
g1wZlDEur0WeBPt70FMWJlSZ95aDh1ATvz3YAW79J80vVUU2Ij4pi1Rd6nFK6nXr
XdqclGAUbsrt7fBfP+StIEzisOAVNl8neQmbQ3kV0PLkwEML+WtH2UXMuZHYJrWu
3iXiRwsj0yNp5GadQpdPAmtXkTiXn0t8cJyN9EbYtuJQxDDq4IdNwEIsbnwkcx8V
n2ecRBvvEtmQW+WhPCHDyFf++2foFqHeTKKALg5jB6kPM5XeYmpomblv2Qo38muC
4IVod+JmT8YRxtGV7lplhikMUEGtC65vZ9OL5e3+gU28J0i27lsApqeOeUpL1Zqr
GWT4tIWP0YDu02D3jsEhd7OWSqAbgKu6Xup+0oX3IktZIihCnjxGEPnXGv1NXQI6
LN8C5+bPDaquBRgQjeZDFEf/9/t2A3tG96fZzCKAcpCToDmyNs28oQ/5kjp78ARA
URCfbpAdGDCkdWV8y/ufCM2m4gn7be2DfwiX7NUFRlYVvnbS/H9/s7rnDobBwC/f
q288zHJ5fdujd/NJXwdSB4tUBX3IkhgaBwUEdmqJlYET1swnpEUJSRtR8JfE0cp3
zrDThzS0bkSfjHMjHW9ILd2riRNDG643j+R1zZ9BrhxPxpaJTOLxk4jACoOPr03r
z7Aw3VE/h7I7rlwM9o+G1CKNGaCjv/AUblsjP9rzuLg7gwSr3Yft8LYBaAJMb3ss
FEkL+nvBXKLCA73FyjcWE5bDwJ69qoNjzsWKACLTpgkKx4ngWGRRumNrgb5j5GZy
bxbqIiANIdDCDqaoL14MPOnOXlIUOz6srde+lm801uDN4sl0FF+wlOzRYnQN6NAS
XujP3y3rjl1atFeJcBxoeYSSdGvk74zZ1KDpNtA6UkwNec1URdVy8oR8cNeZSg+u
BmvQ49o6JoBoICiVdtnn5D1fpn9S4bV57qKV/HjK0hb9PGjCf8eAwD0FxEs+2idf
FbnIWNRPDYt+2Hv86TQmSEs4QQ/vaFiPvomojmrW+stafjY9imsnu9Kg1iPdeqvn
thLZHR+nOjTEUyyLcS/CHWttEun8xUjneHvDxfgbZU5AT8NMvdoA0LKzkQV06pK6
X7lEjQC9/95rRNT0cCxsa/VhFvD4Am2C3aXL5ICi+co+yp0VYrmutODxyk4Cb5iH
FdvXNWqxKpZiqa6oSKNxzvrArHyL/YQQ3qXQFBl4Ovk3HUf+bilYlIb/AKI2+hkG
byUaLy2Np1q58A9Xo9ZlTELZEMPI7AEvgdh3ysVs29DH1pFd7s9WENuyqczKPpNk
ciQn+3XQ5K6m6IUMotXqnhlw2L3rnxKa55uv1A0ogX1D4hRUHczVsR9IS8aMqMLo
/mHE9ElHInwyLPANmN7obM9rV0BXLZOOVxPwnnTopup3Z03uGhLWOWnD+f6a5t2P
n974qdsunxhJYiBNToWqs/DbbMNm87AC9JlktUQVHTTQrsVJeJ4xnWrhml4uz5+8
vrzBsSyoS8mrQcFWI0KWM+McSFSfrzqxe6vfhuJY4K+0jfvvnHL5LKWS69QBXypY
JnPFXzVSqlSvZ2leQpcoPEC2zDMOZlqONgJ5UM8DrT9/LbL7xX0OW2b1oYJ2DNWF
somYjSQcetXt3BHq1eEayYDX4Ap7J0O6N2lbgBgs8Iz56tkzmy5dvWoQMTPR1N0H
uM/KUkWSCAmNt6bfIos7aeqe/Su8fPm5g8nAmItEsNL6zuuFnfjMiQ0umpA37yei
RfuIkhwpv/Z9aZ7boX3Rip5nZtXdzmYQUDsDjxyzRBNRm6XGey6C7UJG6gtmQO7W
62Ptb3tXvHxFYhsqK19wsAECnreYaSWEmxYuXSiIep2QcZy5O+a+rrqZuZtxcqnK
/UJZt9/hSNAWbtv2n8daDnacy/enmfw5hEJqb3Am1Mxie/RuIY3kP3t+7UHSm8lx
65jNdfi2SWzmg5iSp0Npxa7Ai0E5pEn7ewjHU72rCQHZIIjMfA4WJ+8EuPlcupz9
cj4trLVKqG/OE1BFsnYXKu4WBip0AsN/mbv4Q6qQ6u3HPeRk2vTh4pIDsiXDetTR
U3J0j6AE8PRz+Ra394/Obzq9dHH/EI+iOU+6EbOlfNOUBFakzyPGhdym9ahlJ1kC
E2yNK8/tKB0eDeG7ZIbothkjjx43HqFIMQy1iMYXG5ruml+YD7DVOAZ12cnhsuSF
ms5NAFwU4PbKxeh8fr6cDVWOxZzX0cliH6rlX2Rw3TL66rY754V2ML5nwMGjknCA
0LhZUU+N3znyd2IKd/SoLgzu4NL0QCYsAyf3+jxBQYw5yTVVo0QiOpKWGmvt6S5K
9/eM19xsnhu5KUulPbNgpQgp9P84MTuyc/RI0GbomEgstzPo/aUS3WKFAEWRolw8
+JTYyxUTUx+zbY5IpmtplBGmrVg8fNHuGJCXcp7d9+nVAu1YyVTk1gLysdTzAUll
Njhn9Milr2oQPe3MARMS56TYpAy+aayPVUPs9ZkNCQUX2XrL4S9Jr88q3ydIL+hT
HaN1/e2t+DZmxNFP5II0bhcQmK3ur33JNGDvYdnHPxiT7aoeaJZvPGNQ1woJMUJG
sEXBxLJueUkES0j6JBqk4/Lb1Qed5+8GF98ZYgZRznjdpYdV/AsvslZWcOPSurVL
Gk9c2aFDuu4FSHFnWFWWQjM3KM56txyy9VzvyUlUV+InIU4EwX/1z8Tr0aytJux4
WP4zoi7lq9zfvcyyAdBBU3H3cwGRgwHbpx5ExOEazqlN5bhvCWeN7W0ymutMj7eM
iUL/5nY2hIcKHh1XLPHsFpb2jv90ME5qyQNiCQxRh2Tfp1gmDz4wU+OoWVYQYdkc
h/0sJ+D1/smKZcXhkgI5zN18sYXHl9IgKdAP6YPmX0NX59OvU7gKli4U89NF98fr
PNhv70Ok3tuhNf+RhnxJBly3bzqsiRbsutRIPawflbl3VVm1H6ZhnhqgNEZcYa9x
0ZOvdKWTJpCDmod+zIrqFsW30hUPCpm+IlYj2X8FSkssWK66k3p5mVSeMT6PoIjh
MaoWhUkvjkK3nRDSUT9ssBNtR0F8p6+PYCWHFdBCy05LPNyMowyt+FRc0P5ASS77
ZSwzazfq0LBgvchAtwloOBOs+DdvMJfjBqgJsxtMeqyLXhNg6ENOHi2YXxy31Q/j
O4Nrv2hGOiL2KYbt2WSG5UkUcCvNzQNnDZluy995w9Z1/t63wVRu5KNV0b5+kMWr
lv+SxjXmKw+8/q6Yr1gw/DTLo4lRkxgrvcxxaUIWvoNRAulgjd6cyPtI7FdTSRe9
N0A6J/NI6BFnmqZWNgrSxkLUPJGwtYZsNB51NQLzeDP+MHoT1w4MK9jowaSpITuw
WFW/e2EjOBxJeCgHL6FtgsanpN5kx5FJWb/sp6DoZOEGAKyfs4ogRySTHwJVMMSX
8sW4qdBq274kFc88bwG46HLDmdIG7IfZF2YSyIJYkZpNpNX08B22wpJDOnF/pkaA
FGwIpMPpngqJkGuEkA2RfxjTy8aSKIzy9YhP4cIdkj6RKspnhIR2MgyC0GEoVgK9
Sid9Cf+ZB0AdNphGaEWftUDmO/5yZ/4METg46XMnScYaCQ1J+0nU/os2DZC3UgAn
luJB0ICyTI/08xf/4V3pBdlvqAQ8Nc/YGiz1hx5PHoNGm68mXEQImkc9gWPa8Rua
V2Khd7IemNcRfU3LT6ssMRVjtoHIUoY3CWAc97H1i0wdQoPEy2InbReP7kQmY5NB
VwaPyeJ2lyryIFLPzAHDoRcjhnbkFbbOUDS1DkmbPi4542+9mGpMqIuCsP+ZIVAy
VeNLpM88KNJOyF7272/GfoutdRmtY/QMENo7z3MsjPnK/qWAzqMPMO8fYrPiKJ6j
o3oUyZrcWsA01g+GBpn7AVckCr+qTuJqwPM3gMFSGtHr/YSE1fsFtv6tRNL0gPiC
PPW+InBT/l1zfxK7uV3NSiMv9g5YJcr+OF29jckj20L5IUlmw9C6IChRod6yYdaV
ev1vbhl58e8bDE5ToRtj8gj3E5J++3VJxN1LhfJG07iCG8c/hKhSf4jdy1Fulo9y
lrg4OLKKVCGvu13qMajBvabe6qM6hTvRqdtgm+wG7ZDikDgf6nFqLHoWnHBKCYxx
JVnZBJxrd7UmZTd00tRm+6A2ciMK+31vwmrJWBhEi/hmJtIC7BPausA4E1xunbum
hOaY6ovbhQ6FD8VmgzCTpgIwVavT/+i972CpLZGl2Fyixi+Ign4GaZqZ8ejjFvRy
oacbHHAEboflacn5lx5cO4mcqMc0BXV+Cq/P53VBsG1lf+2+pKSGuEndmj+TGWiu
CqAJt1syP9aIa2Ui1cYC8bCUJxTxLgc9NzND7giBifA27YN6S+5VHEBdriMSc6he
Gpln+1jRcloKeCVkep+QRrlXF6lMF7iCrEqJM0O9FdaA1QuhF7o4jfBZck4HYnol
u/NVeGtNqFRydkadxu8IS9VQxQGqwR8f3NyHxl5D0/TR46zTxde6WKOcWuEnJsnf
amWKw3DFPAZbytJ3T5x6H7iO2VGYTwsGVrkxP7qAHChcnazpE3Digc57an8bYGoV
mjR+Ly/sUi8ObUXzNi5DaEtx7NtqSQJK9OIt8FAG6V55KBuzLbIjUVJNKvh2dSTb
JrmFwOH4tKI4oeJeawMef6Mt9xm1xrgcvsPP15R459INCPOioYAUtidTlyanEOZ0
f5Szv9HK1kVu9floUonjI4jVomPIkPM34kGzUZ/skz8FtBKMQwQEOkIsxYjXS73H
oK4ynG2/03wqKtHj4VV4yZ7WmB8hW1XbsPolLKIeXIPHtsna/2qP2+Ino+R8UUZi
Cox6mmkXoAHWGEXzzJH8iU/f29QVhQpeFTB7GbLuRR2uMwpRvd7ukKmsviHqOiv5
AYqiZy/KiEUX6zwa5FHoWsuzOiYrQIUrETlJFzoRPQJl1fDmwWfTS0yOJVrhmoO/
ccFvLkZhRuKM+Mv4tGWEAzT1EQWveT4L33pn6umOdtQWSu2ap35/UbdtoujX1dJr
s3h//IzmZNocY/AIclF/Ypj8u32H9xin28YA104srpyfgvgrGxm9LZnv9OdG3A5e
b5Z6Ie11dgHTR1Sg/+WtctnF7v7b/wSIYgg57pvmBaXDFu9F5lkANahkM9+NklA6
AScyG9+r3bptH4vOABJOTVbQ4OO/SMWKCmol1g5hqM+UZ4CLXFySEhkdQvZkxwH4
AnOSJTkoW44jPaotvpssS2haD0wqMo+rzqmuY75X9mFCPln0f/XXkW2Sa+chyrvq
xzcp0W+TBEAHX9fwwl3FJFJbWt7sU2fGEF1k1mZeyc5ARfpgQHcZWQv91X7s3jnP
L1SQtVKQL0ubvaRWJ2AOVvW2g8OdueGZ7/c7oMhG0LhnLqma4EFhY5KflV10JS6s
8GeI+Pg1TIwvfXnwdABzXf3tCuyMJCqaZsMXy3npN8wxaz8EaXaCvrNcXjP3Bf/i
AlwMIfPQ+6tSGuLWoB7WdbpIf3OlBcQfsOtzug4wgHtrDykmzjidr48baVFiiIOc
ocaC+VGg+h8GCfrN9PdQhFQwDmyQfYpyDAW5UOK4U+AXPjcszhXndDi9DM32Rv4R
AvpLREkemWSsGeomJY0HzGO86qVsQxj3+KvZr5ZBpoOUjySnlu/aC/eeYsvqDSAB
wNaHp49DhsgRi7OtlQJrG3PxSdP7ZkiEYFua0THA6/DLCH3rUdRGTxGMz0zBCuOJ
QbDoSRHqi8W1N6KA92ft7VXX8NpkdqDxAfSIsRrhVC7UkoBneGR3Dr+PdDxRTPIC
sSuv+L9fXFkThWMuEIQevOX902J5/MCE/N2joEGEZu7OB8UE/OIrIBn7LrDFrPNb
GOzJR6HFN0X8h+XxbqvMJPI9eIVibT8pWY3AlLiDDGzRZk4zq3lPRlVA8W7dzO8R
3ej4bhnXbFTA2j1JirP8kos0KA5QbO0f/qv8714Ovk7ziqJ0maJ9ng9mNj8WGeu8
sP+C0he7csCs5LVdC1pxvI6ASllo5kWTAFwmVupyVSG8ziVnIDuDXexKeZIKVWnh
YkQoq2lPaiH9uP6ilbhL8SdfFotwYZPELPO2s+bi00jrbxxzXCUnQi2jLCtiGmt9
EBmRopJ3x0fZcspJbkMUU+xTGJTq0+8kQ7u1ZZig4PTDF1VmTlBMSmZ4cPWmV8rL
V8mdhEBJ/mIRshI8ge9dgIB8kXfwNWh/NTyAMWs20CqKWvljfimXq3F/hn2UlKz2
DXhOI+qf6wSmCzZT5MnhOHLqJ4rcB+b2udRJO2fiBLwIRVG0Krbt1wNyger897e0
WEEigwaV5yPeKjZqVKfLzt3N8avXVC1QO5MKmxbBNl6EBUJ/m8THpcg35p694d7b
Zz7Kd/xrbjFpW0PAqzHwlKcf94wJZsY8yZh9F0q3cmAMycgF+eJ8L+5dzSBbaLbs
tAi3UbkffVpEz6P3w+wRim7BmD8TMoDou6cNXsd9F7XOz2NtJjISA7GrTpIAxgWf
R2i+UsLc6LahCTpvzVJjcQO85oBnOHMBgEjEO/WUVhN/0CY62HHc1pYQ4chLohGr
i9ZsVhALtHiReSo8QcD5BhNeVvASLnynzKP3RFphoZiqz78SlYtayUTamnsMQ4ii
c82+letfpmfFZaID4pjqsiqgZ7u9RuMKWFjeh868iXnBbxE9uF+y5qw6QOuoi3ft
XjgIOlzpFAU3bu6JozvZUSj0Uqn8xXRZBN5IpIQkP9QMCVf+CsQ2a92zdDFy7gFg
WOWAQVSfLDmZdQ0ENOPbJMQ1+EyKlSYy6BVy3kToGrzuDy3hVIW59d6BtjL4cDMm
8igA6gzXTp+yvhq1kcl+NCjTaw1KdvwI/M1qeQG5p846gm1POSgKDZ0Xwrtd78S8
t1e5yZbqS0zUV0E9orTi6bAiqB73R4jJEKkAoA0tZs0zJ81F/Dzd4vewYoVKKzm9
skbrqzmwy5HaoXhxwoTrrdtG3pB9+uwCqz5DAsxcv2Ys0857/TtQwiq/C03BggM7
FZvsN1nc36LPhatWVz8eiDu9miKYWccuXxUuTjSFJEou3Vux+3rTpoFI0nXxP6zZ
DL/HmirPNfKKsfyOpi8lESMpoJnDCZJ6USnCnbm/9Z9A2YODsLussYjrOF2Mcp3r
6iXtw+bplYUZPkxmwX1xvnXNOjsQB3f71A2fJzjRm4uaYrHcDkFFgVBIr566Nf3k
15l8USnj7O2T5ssrpOh0MaXCA4uAPwJbWy1GJCK8DEpeyEv929zxI5s5G9JJPjWn
ZGmhJBK9f0heJdqdBXpAmZ5GwGcPISwJUTYsCxDK+vRzQhuD/shvP0ytWpnTaX8E
6kAPNFg49M90kqd5s8EUuaKPINd02j0VSWUBh5O2mHIlqxvFmHp2ihuIA0osCZF2
R/hJqn9frya54oCEv+MSvOi/6nF10vuY/DxV6sKC3AFvmjHmX5CSA+ERbYDTLthC
DOzZqNfLOKc8Gn6+mL463Had2xH8i2VOGPXSAZIUctK3kTyJL6B58+7aOTFD+Zeo
jZ6HKiFHNzFHiysHIovgFtM0xxZ5AIheS7piI/OCGaSEhcOfWI9rL93c86G1kJZw
cO8TcStUsIdosOOexT8hG5b2e1UUbn4uS8EeAAM6u+zL1vum78L4FlIXi5hpNa6T
f03DAvrmq1E1boDVbUVppWgr0TYaQ+Bpia28eIWF3qmrXH1vD8tWKw28yntH0U4I
wRZpeYzNe0yIYsU5l+d+VpzQMLyTIg7LERfBPknP3rOYFiUCExCAW97kxlMna8yK
rmZqrYzy1xlk2sCmM4x9BLpiOBcrWz6hXaOhHvrYLVnfoF8ZWyx1vDWnqs73jJHg
oVzFSgiltun6PjK69b8geCPpHXpLOtHIBkYBGk0Co0jGsMhxXXcKKEnSBjOUmKg6
ncA8gvq961hV278Q8/dps65tjGNBGQyXOCTHQJNCwCsOSIsBGlwTuoP7M88Eb09t
1xwtv0qEQy+LKnSY44XbEL6EXhZOpn0q/jd3fQdADQPRfA7K/1caB5sDKr0JB/+f
EJqwRGhs18a0pjarnPalrPSqCtRasQifBTYXKnt860GA12HPMhhjyWyPHnS7MqFi
XJMT8lpj0Cficmz/dT5oZNKHQjGpS+x1ztu8ra7MLY50vYvRIyS6yB/IIs0BNs9p
hF/LT9kG9IGuMrMpHGdm+5bjsNPWQ1UqfW9P6U5P4KKTw1b4Zj9NHf8/ffZsk5AB
McwTYw/5peKRrPyEGlyir686pgrMZRrDyXVFXyQ5w68JU2iAthGsrgdnJczwMuDo
FG9O9iOUwhV01AQlq2GpvOAC9XuGsivMMdRApDI4Jkxi9ISEL11liT+PXBK8eXby
iCkIebmyD93MgZrYWZZeAzExDFIatLlVs0rsAKat6o82/a+mbfhqutmcsZOvae91
Xe7QKtuZqKs6Oi2eddjrRvW7ZKKdUG1QKsAWHuQYQlTMDCuF/SyKfM0y2L0gjiWU
zk7EjDbmB1hs6zdNjLo6tDf9N/0lQKYuYtP9nHnTItDbSwzUCf+oaZxvsh3GGXoD
be5wSGDqAbHIDtdcfhyD8f0HxRkNISiGR1wFLBH5MCLhtlTTqfg+aZATJHl69iXC
PomJWeExEJFjfC5X+YKHjMp7OPtrXIr1JVepoxqznJv4PuRhCF+rTx0wr0vg3Gvg
S+HJyfxnZPxGk9C+b2q/r3qV52xN9peRuZSJbyriYApVJSnVum+kPzt/oPujDEX5
8zcFMxEPBdo1SEgjd9Y8xbuHIz+Zvq5KjL7JjP5sF2ULemHLPfKPFhTOS42FUuze
+BQhnar/Qa1ZVEx5L9NK+HWIGfwvkaOBrAwCTxfIjRj7VwfrdkQxzfdmYAXGGFKl
miIjrkhTN8UL5OXZnrSS0Ry+SpkG6F3uq4Jm8pkWxTYrBMqpnq5Ci7Vl6YRk8ppP
uQVwjO0w2ilcOw7x8ilY1ShYF4YNGhtvlcElafPfYUCegTrbda1B5SELdpKNfGQT
/BZjo346da4wgrQ5oUE9M0arnVsVFKoj8wgiKKh2nzgXhpcjiuQbkPuKrrXcEcMY
od9PpRCP60lV0TkdJZccrM/7luZaNOq65DQnH2jPDfK38g/A2Ev5cJ2x1FIIMY+f
FMpfCHulMmMh2j2nS2tWctFSHUEjNrbLQz4JeVTKFwJYtfT/pdmE1PbcF7+YxWQu
iwKF6SD0Y0ZYcvbXHhiGFgt2VGIOnh5HfeEHFhclZz/VMa5yM3Ctps1qHvJ+XnA+
Ohj+XlTHFrEFFxMJn9aVQsuqhnYSF3kMv/QvlzolGtbzPbuiPPPR9swm99oNER6j
L6iAY9R3YRXbflH6g6ezG/igR3FaCcMCAfC1BJCujopZ1YT+4Xb+b1KDjvr5lh5S
0FGEhMd4R8AKfCDi2BD/mm02rcF33XTL5Z7k61adnRQRlolB8xhIcbr8D96rRbvs
maBG4lJS2eUyeBbHoPvnTsmIeVwGKNyYtszf01GwiYH1/+P9zBzzu52VGh0nMhJi
kV9anPZmZ5F4QyTYAgs7EPS8JHtw6a/OPgen+r+X7t1KHvP3jduyTxqLN68PtAzN
uYDh6San7vWwUzc9QZLm+JMI9UnGajCciUgzforPCfLo3Mak1cUK4FSH8Vun9wZM
pFOLeqXgZfrEPFDldDqJiTpoLEUnheABq4Z3I3xLxfOh+lmeb7uOwBJkhajsNQ8l
pbnZCFObrC+VQYSy7wm1HfwcQk/ITgzN2iA+EaJFo7C6AhalWanfiY/DaPJboM/S
26f0foKeNAiFm39BVguZCdLhw1/BJCNDC4YoveVQ1eqbGYAbiUJ2kZn37Y3OvrIy
G3dgUSy9BRidO7Iz7WtQDmJ3wBetBJANS33JsmsKN+qqZt7+tK2D7TQ5am/UfZ9m
5DlfuB0+vBEk1dzyQjsSDO8jEWb5kUYXH53Xkx48Vu9J1ykhH//tFOYdWq30hloD
d16/0rcU/DjJzuoggZw8SZlbvKWx2cWufJG+JbIY/xwR2LMKUDHpXEU/fGdy1rm9
TYFknHxZlkBIzmoJKLLuvkMRpCgWt0bslQkUZbA9DvA7YmPUw+p4+/x/h0Qyruyl
rMs8RSIj2/NGiWKCJ+YY7hi4QnNAvj4d5+30UtycvYs00K3u7H0ZeUjOFSVt7bzw
eO98aCoLpxwoYeLn6OptQTdifxRYmv07TNqkPo6gU/6r1xfiO9pkwqwu9rRrR8Pc
N+rIYOPheGm0yPxLVyZcj1CLhjEFUmDCYzTsiFY8vwRMkUQd/2kVPg+24dv+DAZ8
/oXCPTN/YT1QfWKpVaApbq4Fp5EMHc4+5b2zJZ/tXC161ghCVFEueSeFs5O8dvSo
EQzT3L2ZpAbisgTyGpqTF1HaNO2iW6YoSVHHRJI10rsTt6mCuayuGJHj+XB7ZtLv
ho1gNM2WxInw4vAkI4159VxkJgozRvZBqa7YJdalTTF+btk8htsPPvTUC8RUe3yr
dGj+Suv+5mvO55KAfJqmNrqBUBmCETgvRsVYuAophWTZn0m8Iie4FWLVxmKvNjod
sSM8VnE1migvJmmQUrXR4NE80aJh0vjOuAOCdHSnLkzXIbH3/NUtRMufZnpQiZRn
OdU+VykdzBzA1IEl6wpw2LzWl6tglfx+IYpMux/Yh4P3yDVbYnegLnSGb+95nZOK
2J9GBECgZnUDWPg/Qu1OBPKdNRblypN2xxpkfsVk4EP7u+fF4+WHfLhv8AcT9gMH
btFJVGZXRb54Kjpiz4y8vmtQjo2usQkSsk2Z9cX4zl1D8GC6DBQJxP5snHlhISSz
NGeTOPjMXCCtjozoScy1FcWrDX+hUU9ap+yX32iQ3wTSWNz2kZzFRfNkCsbM8nJ2
Zh/aYCKqphKOUHDDDMREqlATCB1zdeyotMOEuweTzUjiP9DOlGTwumn4syhW9lbL
Ivhm21XxgHSjGfpjRbWYPT/e8gY7LNUnGSb+tpYkSlWkrASbcQnWPVK22sBKoKFy
XVsnPpE+eUqebrGlcwpHTX7z3bYTanWUgPBoMcfvlBH5FpGjse9MtnIg3XZUJLAF
bAi3TrroaXYi+7S5JseTMZf/Kdk8cnCIYn74Quu+X3LPRIKFidVvzcJ2+7gFJSdA
cc964IEyO59nJYSV/0NDi/eVje99/asq856Jr4MnYAU3+k2elBbATifH3rHD1KtM
B6GfvZJCUzqWJCY+cWU3huzsl5hIQR9JMqYLKHGFzyUnC7e+arROA6Lh86T5Laii
PGGlBdC6me+Mn9d7hRw1gxbTNQIn/hWxvqaF2Xl2t0/EU5NyoYukIzIMKMnpY+qI
n00OaVxWS1a9a53SCT/E7mj1yheGdEqnIoSmiALbNnLTNBn4+N2DZqAsZVTZiQBK
c99XPWDMZ50ZJP6XaNqiWoAUoYIzj4jdi8w0grghYod5Lm4G1yxes09rpfgLA4//
xokrJQfqh2m8V7En+Xlv7p/zdCJqwnwRXS/7gyHK80RSf0S+7SJ8PvzMJfMjQcKr
0e1/DdH9qSNz571j3ddww4ShsXAIpvtg9xFAdGS0ESUbSTuLT10hhB8ntRqXMQq1
VmLCV/y8NpVF2MVrCtCT4+m7FS0H1buDw3hrYJvEvDvc4LAeJTL6G/1YqU8L4ysy
L0lNjU6ldgkJX/IYQETlseTibaUMgBhVzt2oImFA2ynuYlUDen6havHR00ME6YoZ
fT7FcCsxDk78UMgMgo0vvDeGn6xhcs5cQ6eWmwIreEkz0Ic77W6rWJhe3mg9xgAQ
f9fqREO76v6H+ASrxVkTUT1NYU6EmQrfppwXFhF0z8iugqz8aMYoZ5skOckwPyNA
q9VG0mnOY9QvBvlIxAGZ2USxenxnfYdoi1SmTghy8NK6bhb/5HgQ0tOvFVQ1SGvF
NojGAs6qXXu1/d+2FNmi7mfFBO3McF+k4TKHO/Byg2P4c4Ls0uERfwOdit1D9f3u
rvXaVIIENvWC6ZRF6TAQ2xgtmMNLazFfT0qfve2RD3Xv/pZRU/cE/H5wPYSRqR81
9G+thkynQWCtGxtBTWPry1BF0h9FSd6TtgF+lgjq3wqNN7sdGCAmgH/kHvR9Cm1g
ZOrwgDbUbt9glSnWBscMtrgxnwxbWvARf5mO3sfYTFgmpAaahQ4Qo7r2WlXTwJJu
42VDhIo7reEdGMLpjzJ0mReHBfuIXTZThzz+ioPuJWHD6XseEe3S9BpByenK612J
PmrDS2qbN9CU5E0tVnl/LQVfNSEH6kzkSprsJ7aut527EI3cZtxcKjOkbVu0JMBS
cUKQSLzUxh0lqcS9+gCsZqbOZPk8lp2lSF/I2jP4iujAySSAlR37DOsFlE7e1U+l
ujGyc9ncqnqsM+saL+DZD+McQbBjTesS7oIdKW/cZp5bSgPwEzgGzNjt4dcVzPvo
3RN18joscPMqqNKWrys4aceu0TCo1yCIpXpjGrjzL1qqdpM9z5wLn97FqBBsUf37
G9/dDsa9rJ/tg8C/s/DwFc7QGDQCioSOBqz8INb6HsKZyGIoDqLGw29NJSFD2DNf
Nx0rE3tyN7AhLbfHjWAEAj7/PpLHPoyAeTPx1uys46J5ceg6wOGoWNGG/+uJDsWW
e0ifId+Wm/1Zv1pWe7Tp+njygBCJ57RQOSMn/4OMny0JTR2YTwWpr7VhE0uIuPkJ
PTgKTy4KgIYdr0FC5ibSGK2RIO6fiiZvQUZMx4pOLKNznUPshaLXYMFBRk2Bh7K3
FqpI9h5VLRQOqLYfG+X3R6glKqY5PQ3RCViIHrrMdJLSDYmzL2kR706rX9Zd2FoR
V0xO4adkEPObY15ieUWYxr7KNF1o6V7MbyBZECB4oh1h30a8R5WZt176iVtL9frz
b0f73hdtWO84RC+K0444TtirWFKtyucde1ev9XLo45Ay2Tt1FfebZt8xopbCmq87
reJWwYrJ0FIkpsTec2I3MzIAPSNf7TNFaUbPfG4EqJG5WRSLDmhYpjcY+p2Kfamf
IdOA6fzUSU2ocErWmT6IkPFrmPme79kZoUo7Hj6NHRNjTvx7JDJemKmSxc770OIn
DOp7N5N5Hcznz+V7AyE7V7cMKwmIv+Y+y6fxGLct7J03e3UpUpYqbcvzOVz1hu9V
pMWNovG1BuIJ5x3L3xh4CwBXqL//oOmIFO3kJNRolgQ9EUjLgpSKe0NLU6W68W1x
nQWSZwQcYBaI9NDQzUSv0oB2kypl5LOrkaT6pl3LHk4ooFWE6gnEVo3ldxnzego6
RsME7YArWnnI/pTndYthIxg6TuCsyA18WzVbiAyb2xkNCCMXsjHxWq+U7lOEZV2N
7GKcUpfC5wPi/Z2a2Nq4osHzNpxV6S07XjpIe8g+bKJIgOysREZS9gwVK3jWZYNO
yy87RsnRzIoV7vj2cQgjOzV7jRa0WL0I0uCKtWIiZ1UNhFAz6FoswLpo+gVk213m
zmGJoCo2+c+Ogj+0FXMy9BmCnMzBfM/SsJnL//UGVYfY4Yz4hAxlcodfqTzS+IEP
Os7+cetO2RT4aFRMn1Xa8wupsp6w7Ke5h28h9bfv+UNvOzQk1fSmALKv5VtnVqdx
jZDmPwZVzgUIc5KHwSZgPjU6v+pZL83kMoJ7x0VtFR03WjTVbM1m4qQVegONsneO
VxzGjCzOI9jyhgzRHptPnOL2YRkIq0MRt3H1Q+3v/uKpg0SXSRUKw8bGeVOmm5Zf
3CivewLNaSnRM0WMesGAmASkiI5nMEVIpbPH1ehltdyAgt/8NeWxeTj+VqH3CBT9
V94RR213ptQj4WNY7KGLwCHWYKW78oWE12Yzw+u+ZTBqs45ofiIGR0BHWBBdk99N
VSyItlTEdRuPh9OUCUaVkX4fUzNU8X7Y/yXM4ZxI9mSJIjalNeF7pqGF+YgQZmb0
7maemU2kniMF5WeVqPk9gvsJNBKPTaDkw0gLJDANa6Pi22rCok9+nOGeGsnU8pho
3zQSG7Q1vr36WTsiXHX6ThH9rz7dgr+h3N4bM6Jf19U9Gf4Aw2bAWaf+dwSALUk5
dTCeE4HJm8LAwO5/3XXQeAi3kNiRnyG/EIT12EPo/Qfva4rxCS0UsZd98/TXha8w
cCZffO36R562I7kSGoJV8m/b08RjLIsCyMJgRN4neo4ZWS5eYR4AEVgwHMvGo0rY
HSDZS5iS+ofNjmnaamTfye5OS7za5SQ/P5zCrRbIv6QoJlG8WndmpPH74lLEeL0s
1mFQP7WVctpsq7teUooaMtimz2AiXXCPVwNWjvI2zermshQHAOxBQpb8P4PLcGWc
qCJY5AtgiNEj6aTYdly5HcAD14lMD2jdMizfuNzDvzCXmilponjV4L3n10+GXUTL
uDRaAeF4FwrfgZzEeYMzTKDsaE/8WicevWB87v4NG2ku048r2/kjJX8mivfWu0sE
NqBRGEkwJwe1/gl4377Hz8ewizL/SYR1846GtmOSTRi6kdnQeROOxgEX3Iwggy7v
+GSlr+4+2ivjNuPXa5M2uIFNAifSDsEIaaD37tl7nPOk30gbNX53uaPRDSz/7VUx
skcnryO6CKVr7RTuICaFLl8FgqhCchljWhSh7dWsUWNG0HO+UFwbCX4EBx31blkK
KuHU48Fms4mHFdVNnL/XBUQgErM1VcJ5Ati+Q/Rbd0/l0o8fwCJNYm0SMeq/HSze
terCFDWIbesYgTMXKjuvOEvZkyl7YYID282vIdyW766YZNfUxuywtkbgLIbcSA8m
1LnX3ZweNEP1qIp0DKXdS8ICqU+feNZZEa8+IRG4Flb7lYjv2X+ibOlvTml5dtHc
5ctG+iA/hn7lvVIzkDg4NFLFhzfl0PEAU/7d98hg5iVvZHMhrRh+qpkI542e0hrM
vyYGDcwiJRBeEvj64o3tjljslVmboG2YZZ9X/z/C90RvNxLsTwDMuDrW5oFyrqWx
+I07OsgZvf/HeiFb6PMTpD8ytrw2aO8i6Jvx8HAcREQ7R8SXbbm/sVw0rrpFnXld
+15xLv76apODRts/pLKiHSOTFla8kq0A0ZFsf/tYCT36vV2y1s9S3u77bYjzCbbh
ZJmd4j3L7E3YoOvsg5dE+YJaM7xN01EYu3CVm5O/ClT3mf0YXguCj+DxJ5CWMkZu
LDNO6PdyEvPY9fFf8vpu6asDaPY69TrliEYwdaBIl7lzm7GxTwfSOi0vAZKPH8Jf
Vs0Wa1w7eFTaguEs1ROmFG9RkkzHXh6bc5gO1vYG+Oof/7pOO+Voi5nC4REtFw8A
zj+csT0tIo2MV4m31Te1/4eMQ5kbljambh8kDTJvE9a6xWXxF65BrQ6s3jz0NW7E
3vghRfS8gHDOF/9gSJFmALByhz1PE8yGHjiNxswWyn9OW+ouk2y8pxfp+sWFjoBq
cjS4N+gHOZ74Q7uCdwH1WMEWIOctbdReK67J0NPm7Ukn40WHcZl1BqcrVeZ0qNh8
9Z/anw+W9x3LfN9hVciMp6d0UjFV7UrLvuRKJ9FdHk8a9F0YLNmhte4rEcQNJ2qi
h4xEc1kihcbEeBBKrW3LMykDTvKGlRoo8+x7GMftPxMUcNCgmtOdUi89JS+8TBE2
0Nt7PD14LS3ZRM1oLZS7PLz/EcUjdHS7zvxjaVEozUEBJnMvXjrRNpQF8P+X8dT8
xmrWxHae6FxAOTZZk3spNW0NDvTbLU9yCKovXUl1uqj+QBXAijJocVzPTdp2j47r
cDkC6RFZSRIJMA1O7ofg74sQ0ZR7U8DUthqdcp9mpDqR/923vaLNxG2aBhAJZ6Ok
IRE1VBTxXtbeYzjKsRBK7D6EszV3PP3T0N7TzrM6yLWlYTqikb2oDLJNO+sCURwk
ELZPx7XQkv0jaKib7FA0xLO8f+pCAHraNzp5L4Kx+TE6n5dxuuAskigCZ032abE6
30A3Twe66yMQEFxch/w1v/71U8pjU/ijYbUJ61CTFHxFeaRXIufO6MMcCx1OsQMS
1YorHIPMlXHvTpx2oALdoXSa7xGZXHSw1/EbeB8wrZ+oxObDbxWNwS92pW5bLHIU
M6X0irlOjRCrTNMbl594fesssixwPDfOyN1lhu1WfGJKiFmNolzt42XXeDDcN1qD
2swN0nHfUNCB91ILh8FdWoc0rfiPnuoaN6IERG0ifaR7uvQqKa8tOAu17BOFELOJ
qHx3yU+BC+9iUq8zoxRMtbWgw8jFIUn9vtbcgV+vOo+/lVr9aaEfuPCe/OkEO7pL
a8ProSOd3YlYf/VGW1k2jsvhVJMG49F2UL8AQ2p5jqHE9JrJ56RFljD9KpgMywrY
jg391AAkeGZkOIEzwqD3Nj67JMLCTgaRCgb1sPBqsn8Ea+sDJW8CRqsPGaPv6GgX
/hJwvdtXyVEEpt2A4/imNL7C2ZM4A+BHClfuHbpO45r3RY87tVIOilCPVpqRpquS
0pWWWkEWBxreDEXzjMnKgMpone+GoKmIXLzDlPfVPniJ9Gy2OOvKCRSoVyLhiG6L
gBFoSsoM36HpyNZkWCa4q9OMWAPCK6xEojQnWYY5UFDn8dZjYrkatOHTOaO2AW5F
kI+xDqAGXys55f5x3SmTxZHRlZdDgyEBznCtUsdjz61TVnttPIfKSYU2TPErIlHF
Vts/koocUNQND5GvIki1Skv4RW3PH1KhsrniCPMDMnfLqgE+RDAfHueuDFePAn1H
w3x69p19i1UIyL3Pj4Yma/eq3g5z2gw6hKhf6bz/r3YgGmFR6pUioguKecSD2wN2
C0dLtq6X8l/pRqbfT3hSR4xU9nfbLqXzhF0Gbbq7mf8uqHvi8gNptHdDxcLkyjsR
eSLnDLXWYugnMR1/rfxhcPtDLTiH9FJhHVhv2E3T0hCyFGIze6MXYrnYAq3+qRNI
cRMB6rLyl8+3ZZT4DPjRl42FGNKQ2J7a8I2HBFyfst5lRt4zgP2NRlK737EBkSII
U5UMXKVwnGKl+Ac5idBzj/yfHTEiY2m9dw783RliB5aszAm32csmd8/ary+Wv9ON
LNCbaNQEsfeAXZuma4cuDsaPyn2ouT//gLDjFBAk+MXvO/oe2inZQHrJbJwa5Hdz
q3BI13BXlfzgCJQnHbgSuzciYTnmc/ivSuj+HCvb0DOvt6Rtjrrp3T3htQ26CQeT
S4uRvjmQCBkV4rPP45e8/mN1YANVkgXXwsIyApVIEHBZ8loPht3KX5rqKpq3pViK
ROVQK9GZaMEVRpbhv9dpXjWmHxfokVfvIHjMUdxlYJ40ZyG8sZ2z1opLpJHFM+R/
97bz5/i2aXcBgA3CDGNtpNt0GvGsD+BVp+xepDmsbIrEORZADEwmoN3x+1sg3ZSu
kYMFpc0xJchYJ62xKCOU4YNJNQZnoke6J9Bv3T3ZPhA=
//pragma protect end_data_block
//pragma protect digest_block
ktXhy2xDeRSKDk78S3HSrAs9b2E=
//pragma protect end_digest_block
//pragma protect end_protected
