// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
XqwBKBGq5L0TjaCgXBefAOvIE2+9P1WS1Nk813fPgQy5VpVC2WAI0lZ9dRlL
QMTOFUidDVdgz8ODfMYoJcqovdxDlQnLDuKk2M4EAuGRfaOpBHBfG4HHQjXA
FagkA228VyywVIa4DDeNJy9KCIc4Lw6SUskzOCIDrwxwMZrMw42jGo7BqURL
xiMMqY52JRAu6A77tXMa5fy7yELQOQ5pB0gScspw8rmFt8peikDbgUocqyrd
oBJm9V9imGQiSJAdLm02M50FVzNB8DgMJkQ3L6iebsNt5nAEmW03ZjzfW/le
QZwMZayNDEHT1moVOdEBNyyIKaRjTt0GS0NQiwjqbA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
VqrDlIpdXXCvKYS0UtsNHVrRRkPs5HpIkID5I8WDlufujsja2chVe52qngQJ
YYee/kAJ38WfxigVSkHdzsYPZO1r8fYO46LaACiFRNIK16kqKcJe6DCvuPaz
7blgaai0/rRV3ZrYypU8EgCWuuF10Rd/ZPUjWpdRKQ37jzEG308IWkY4HU07
zdKasVTy/XGmWUNeUqpgkOF0mIPoEC+b3oIsQCf9VizsQohLZwNKuUOyWsFe
mJXOTudSrrzkT0RzdwTGttGiIwfImvxn4KV+zrlVRZkEEe001kpgekZbZxDv
kYQmeci5eA+7j+l/MOhP9PqjaJ1waWzKV//YKBIKzQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
XGZLS2AEsOgLEKZyCMfI3KNvIi2QuR5JUsVJi9Y2BmgPoMGe7RNIQL2OCiWC
AxKg1c2cqAS/ql9Y9kV1AXSJp5smZ4hRFdAIvZd69B7TN453XzkoaFj4ODRy
tO9yY/ccxcK/Unb03BLkhsKjhBuR7F/zZm7+i3UJ56/c8PWGsrwqj13AhDTl
9KFvMPcdguFNmU9ZIwwPAb6J8tVJ3Wj1CXvhdif8+ZXoSttTdNnsoj1Vhi8w
LpSjivnTVVDiGatsUgp8OMxtzdTJN5UHdJX6DsdsY4gvY6jZjfMzkkImXsgW
pZ2bFs5gznHKtHo9x3hcD3nupWI/1UpgOJ1z8IWL6Q==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
kHgg5BB0yWByP1OJWy/48DSuaEujmaHJFkrEPd4r+lCS0n9Pids+nrBGvgNO
kkTWYJ8+QWiHFF4D6OHqgSkt1Y4riZQER7W0cDmmkXkiySJrT9IriPSKapKt
vxfG2mEWw6sz5hLIGhDN0FqNE9/3lDo9cfcrePxVIPdlO5y+geg=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
aq4BxB+3AD1oRZfwZUtQINsMgg/X47MEMh2KkG6ZBHs0uim/i/PoZ4nO18sy
1Fm9hGUuO2xyz0gwxoNq5OdrVFesrlalCmJWxofgmKkmgtEnScx434B5ocKy
dBFOScknm4f+mvpNdykVkWCp0WiHluuQOZasxFdEz1lQrvkZoDm8jB6nXUXb
BQH3XhU972rhUTl4boa/ItJZbKdoVbxNlfqTkmxUYiZrwmldvI1BVxP7/O+q
Q0HZgHJ4QHom076Sqhsk16z6PTACzANttdV7HztRgRMfSLUsUCgSQ4FS5XoA
UoSoDvDU9yeNpED6dWPvOTcyVGHcL2+IGHskB8GPYTMGS0VKziu+UYI+I235
LtizrVyb3ZbqNPsdqHyUTaFjJlNB3o/NDgMUji+sjsdpIUH406yAv0OJSefV
8stAGo9bOcMQrprI/S/EltbFRgbYoW/WdWbevU4+YUHPA8CsQTXnCvcnXkGj
15tPkY5VdnaqB0ZbYrTHKT440mALCmV9


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
snYpevRchvqfSX/facCEqLrEyqrY8qSBN5/27b9KaW9l6iaDm2tRvrv9R/nD
pMzl4MtO3GyUTWLp1bt4NCHfyqFHTv3ffuRrxTB7KDMt8HGDtSmthgXydSDh
MCQF8yNY5bI2ILabRNh3Hrwfc1uhgoPBTfpkzdaeH+d299qTUNc=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
G9ejC22H9yhsF1Rg1gFg9jX5BT4uOqiY+QnBvOIeNRoFJCK7R79FJPvF049T
E9fe84A9/QDPgSLy/jxYAkYHF0YaNVifuGKgFFmkJrCbUA5s9mCd4+4EwUVv
pMcq28E9m9v23v8KMXUgGQCW5hRgxqWFrKcCUhN3Rsa50cCsasU=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 2464)
`pragma protect data_block
3zBaPLjgj4U9FJvBsZmroPRjsFBb+aVTlSCRSQcXlr73AYbn5EomAV0B5jwO
xk0CX7V379f5RKDXE06raLJW4bEw+oyYhExYK+MTqC9zTC/ZDtuTJyLio+vI
fhBGvVyAUMxdS8Y7NyeE3GyyErZFocMd4y1pQhpmrzgEO5v6FkY61v8cDcEB
W94drBBPyXRlureT2GCHy6CAdXrHb8hnQIuy3wLqaeQbrMDMON+zcIvcP0QE
SeU/twbCN61cc9OaFDOvyhojftYKpuh/pAWyVczqaJz6B6QoisSCqHNJ3Phl
s1cCdEFy0RxiVrd+ypnV6ELj3bwxaZnnzysD8l/VwO1XnNXDlusqt0DRiPDC
1bWoYzH3+TSwIQnVuqrLX0FmcQIPKB7/UkiRVpBsHtWspMnuiPNNYYMpmZFS
Ipo9Ch2CoEvGes/75gAeZQLa/lyxFMQFa40GJs+44kuxuR9wAYCzIbo+K5xN
7F9eCwb59NS0HWtHXJFKGelptNekvFI+Y9zKdFh+UCXdQjLtcjkAjaVrNl41
1xqVK/8jGD9VUzm7CivAW4OFYau05ERarkt+Ib4oR0Itivz3IYfHvYNrhv1P
WRmhu73TwV2hNTuT7JXTrgnLgQBM5oNZ865eCdkzhRogdcvCbjTOlZdg7ynp
FTGvCjrlei6cXF+vt6hcSs2k0udKSB1BydMb2Lg6zi4L5ErjuNPcioXE4YMu
CrArkFgjWbt4F+/8xRxpJMRWyLmKOCEQggPnAdAMi9JF7n/Bz1yExqWhZ7O1
0UOo9YCqkaq3cKoPFoqIs3VFQcLj2vfRZhpZdGO2oqkDrpIkYgqnXJkTunky
zp52nMernyFANBaUwoQmQ0yCLiXwaco+JgkkVUbvqTpJuFmU2WjQ7SREK/Lp
XBZLt+8KbVvOchEjUB7HEE+FE4KscKR27c9/W0bw6y15Gki7dlLN1U7549Bz
Cr1fkARcMwkaq3UL38khg8iEM5aZAkrztXk2hfgcXKIpuHfqWTfCbO7alN9k
1AWFo+00C3hL4Pk5JFSBSJv3H4D2lo2046Nn10rLzpCjffMlToI8PFAzZOyA
Ffx7NpGvXV3Dl4mjRUSu2D/c2xlq/42+XlsXueyXydzXTRoa/nVSQixs9eqD
yCL+Mxo1WQxBdRWZtw9DwxHpnpzO7Zg7RKoJACtbJU+zBhL+7hsBNPwHU4CI
DMKGueXz6GuhrMpJNYtvI9fDSFVnTxXBRFxdE4hESTg91H91Nd2qt761xqsV
o0E/2EBAjVihuDGwGmbC+GU12lpPzk15u6BNzcmABfp8tdBO7A4a03qnfukK
nBRJSegObcVi1UjF94YP+xGJsF5MnZde6vazm8UYvaL4qVWRCLmkRIzbp6TF
Q4wUD0qmhfhr/XZWa0SYs4tA8Kaq/EU+RTKWPR4bQQxYlE2JOIyujhcte678
ysC0/FhR5iu/OytqjfO7e0wEtfsNe96VrBTRnjOR3ECLVn0Cgnwg1KKdBICL
r7er/1USuz0XjvHU+hl9FeJXXf8cBQ1aZsK3if3ykE/D9JV0hnVh7+hsIiFn
BNkWFNyiPJrvpWUIAYKaXq1Xbd2ffFxy+7arq57Lb7atQx48sFVwoXmVleKd
4gBZKE9kveFqll06TKnVfSMFuvzfYOGPiurX6HYOzkgI6yV18XhgW5V8DDMu
zWo1l1IAmvT0PckHUPNVCo99Il6mrV3zIFDaYhgNpZyje8FNKnJeWxNfEzEk
7U+qUlCcz6V3/iNuCwijUOAq8nHJ9ylCPxSjEG9cPrHNOHwyG6G+DG+xMTfz
hXa/mHJ1RDQZPBiLDiGaathCUMuTMWQMRsp810zMJikwZKIc2pt3z0lMZEcP
StSms6ntrZyZIWxObrds0GPMFj8kHmN4sX1GKmPY6Yw+mcr374K9v5aIDHRM
3HBNG9hL/BcumX6MOnzponyKZBTkD20+CrH2smTBmFwJoK6SqOVc9GkiWlNf
L27ktx9L3UCaMAw3S09a61Arj9iXWon8www2tnlHszgYSSKrfvIN6J9sbv0+
1uS66eTf3nnwLj+po6PR4AlSEPpAcngk/EeGHG2YOw91+xOI+kXyy9fI7NB0
ry+ciouWTrs3NrNAFe4VAxnlcued1LKeos8nwqUfRWaDK5LBOUS/ejS7j+R9
87ojk7ncy3KxLxDfqZ2fJV7LSUcMxGc8szXsdSLEcuwg+tKr1/Gom2/+PU8M
RPdyDy+KBlCuE9NwhXgqgNzB20jelsY39WfY/jcO/wTMfpK3mb6/ZnBuS3g5
Btz3vnnbDMkOIlSSUbnpMFcWEQQu5w1Q/zphR1xMo62TDHx4aTVb5KmnMOqE
w5JASR7UBuSat71brR64EMSi5+T1Ib24Z0H6E7oI9zDbBUNOKbRhGnjEFY+5
MSJjF2KWzvYHAIXne3YnOkVrPdCflp0NrHiHNclPIN1q6PPFTo5tiE8MYLQy
uMzZMZfKAeJMNuaOP8lUlCRlP/134t1xvXbtcl8z0mdBUj4Nvu/YArSceA3Y
eQLG8EfMOPk59c7nEoU9P/NfSU+JGXx7+LHzBBtiT/xPWgLieRSezRVi9BM4
CwyJxnewo0evi2anU8LPPke5c0wlOPOleRrdnACUXhViesxoN7luAen7RAFw
tK+6X7lIOPE4ECHEpCxQDO2mWzea1dp53yi8hW+r7zWyJLVjKUX+Ni1+n7vs
/FF4cx5qMwfzEOSV72FOXf+WJcTniW73GLmS2lSHZrZ2xOGghQ9jHxyGLOWq
kMN2RoGEeP/NKUDGPh37U4Na1iyToNc5GBOxy1+SpsTtP6J8jxujke3KMeMi
XSEPvZMiXk2RgMlP+Kc0Fl/wfWCkixlIrMTyc4JugcdUcUYMdQ9WKDSzuxN5
2iuF3oNlT/MWHg0j8++9Zxk6nQexq8ECE7L38rDqyAGs1H+KZAGP5UjQSWux
yEe9/9MY/MVYjh9RP+LKOuPiwl03IHbuEtOAI+X74P1X1loerv3gSguDPXVX
W3ZseQlk2UtJ8aowMuEr5swR77cEng5SVH2crrXx56CgStq2Q/DyHTBrWttE
pnDSB4g0UrNBXc/gpTujVb95t4afySixoOQDnkSU+gkIuxrLWTOntP1HLSZB
Uz8YB3zERoyfC+Sv9wKM2nLkrjwBRitSS0FeyveJUl7RNdnm5gPvwXv99Bb6
D/azhpr08JvIFg/6TL4GV/ejfuF7qg2P6twLEP1EFTtljEHJW1GDJFVpvzZT
rdNabtTAQBszB5PdI+Z2kwX6S0bRC43+Y+IokuOfcydmWQ==

`pragma protect end_protected
