// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
FykovdGkxkews0evWIk7MFljjamAkIy8jaTMIrvEnjLQxa9z5R4x81kC8MFIJfII
9QtTzl/uxTIPe7GUs+6z4lPEnA7stLAMfV+mhZ9aA1qOH2gMgvq72TcRxJkOZdRQ
tP86DEUjRE8So6KvmV90D3ne1Aeo6HS0XIzlE01GgkL8/g+l3Dn2Ig==
//pragma protect end_key_block
//pragma protect digest_block
67z0VFgVF7a584bNTRLuzl/taLI=
//pragma protect end_digest_block
//pragma protect data_block
qjScV6Y4KW+ChnAKgjHquarF80WTbzU0IaxxzfYaKl2sqNAkcXpKOvj5SfloTkDn
DUwPc8PlnMChC0jd7Uu9Ht98TNs78GjJvKm8vR5rjeZHhMpDjSf51CihWlrqe7kq
6ZBYcZNQ/p8EMITSGmjjtmBRsOL5/KTr7cSq3RAXceQPNAHJbuciaXk+dYmhbR4z
FrxXKYeiIG1S0OQjNnyD6aO+DGBmzSMY/Dt0DvV0UyJphbWKGM5zEqjbKEljLEjs
6QkEubPvyP6SJsm5P2rjTVXmJBzAUOnhvL9vOIfigXnsA1AA1/k+UUSilQE+bMTi
Alc4GdwS8vVK5+r/dvItxvvyjZRsUsrNBxstZ1RvLGdjwnM0eFwd01dwln3TZtOe
2cUTh7qGqfy6HIqHEVNhdI9jk3pLX0c0SybAzJCSVUiPfhUMEI7mb9OzFJwBAndY
UM8ZrUEI+n7+o+PSaPYv9PUykb7BLixbHgVyd+I7/siavNK3citLHIMea46PLmsc
Lv1x8KwzgNJnGi0Z+wKxnbqXUvthGpJYiZffLNomcEuqM5al5yIWWFUzoyCa39GR
q5foVhGK//8iD+QtkglUqP1Iassy+s0YtC0VsG8oDS2i33dY/IbGxVpAONfk+2Sv
SZjijbv72SIJAYjROGkhIZiIoE4rspFMCEBVPfSrkDLbCPHlxULKLFyusNfPPSH1
mpWxGxuY961XKVlQD0aFclPx8oN9r/HUW1F0d4p7j+z1ownIt9GkIQV69OrIX4/u
W1uMrRqYWx3TjwKdjZ3525eY7d1N+Isgm5/+Yole/x8hMDFz8n7PYOMF3VoGlBfK
L7vHQnkcr8Wbp4j9J71x8lo+Xxx7WRbkje6U1a5Vf8Ug5D42o8ywY1ZRjHSPoNYl
gpgLLKZDfd7DKCjaLUlsO9YRq46x1jfdOMYZs1WdsghHgi3x+OL40CzgXaIW8zSI
BSwRfEtMwRSO9Ll7r+VQIfePPy00qP0NW8mVr78y2ldusb3t/18FBR498mn7wIxN
OrJIJXRIyuiFZmmObBTFR2qTLAXMUkaFg2ndYTylj8TtoqvUTJCiIRlU2OiVH9ES
PrlTIUjp4XP63Sr6yxvpoUGHhntV++MY/TYrWAm6wN3pobMlx5Mn5TO9j+wHOtmB
xOvJgsGAPZVJmS6TuaBtqCn6lEe2JAbK3lRbbMsEYTPgBAR8+QHtVl8YL9M7LA2X
w7/bdYK8P2aCtaM84jxPVQaoSMGUqV55FxdLWTzCPVOjD8+w2N9l0z9MIsqgpltZ
V4J87qu8QKM2AdVsePR7h+dQc4IkNqJfIXIga/hj9GGcdnAshccuQaeUhAwuMqhL
mbKqTXrqjfjv3pA5R7qF2HGxNmRnb3C9IapWE+DwZ2AcA8yc0P3AKahNanoinDUm
17xWFuLXXlVLorhj47wQQcH1Fc23FvAIVKgBDJh0HXdKpq83vj6Jf0QPGE4uKdll
cUHvvS/rE2ielXyaItaT8UCA2ljn2NFe8nboxLZOarZ+aFzoeDa6MObLRSkA3OFu
TCIgBVB+PT1BRwO2cfqyNIQXyGHqwbxtB63pJBXWHEJ+IZy6HkiKvJnFtkq6LtOK
2ojseuXMSNMHpiPbgorbU3QKH5WyIl3936rNZ25C4kEEqfIHUa9m7WojluCe1wpK
vh4vAF8/rzMx+ZLq0OUHzqnZsAEcAsloxYRRDNtGyg3DWrK4toDF5RI4SvGcFA66
1ixko9t/FWuhKG3TOUdiqnHANkagQZfpRYTPK8tUmAvvJrBhpKTe0Bnt9AEDfXOJ
+WrLx2wEykS7olbD6ElWLqC20/kvdrS+mwXcsiIoDHRO2bRQpuvSeuSv8xxU/+Oc
z0CDN8zu5FkIKnNWAPCfLL0z9ayIXI24rUESF2iu8x5wHO35X6B21PB3bQVMlrhC
kBsNQ8iEQ1KYv7cRMpe0HWWD5u67FKVi5gyA4hP4PopktUMnZCrbiABnO8uZYl0F
MtuIfmrtseksKJ1EcUt6atW8csXgwsthrxuxaqBBuEiAkdI2QjOzVflQOR5FXwmy
DvAfV7w9oukbkQdoYqw66rRpzd7WoXZ5PsuwcN9c4iHUpr6FByv/G0AWKLBS7KeK
gduVnvLeWP/BXFypQWgYPwFM1baQqwWXXRvwVJy+Kh6UX2pKzCY13rxGzpU3XGP7
Y6JVi9qiq1V1HdqLwS/6ck1n4wilWLcL8fDgnfzbqO18pU2mvTrQBkG6czcoidjS
ftXwzLQ2HmLAlFamuoIIDvQqEESObmYzrtpvaNtnypVwZaIoT5AJ0VMMnjk4F2rY
rtXNwBwuP7q2rylgriHuxhzY4FfeU5m6SsrCLacMjblEKXWH7gz/H2qUdUcYr6zz
+xP151mEFK/1y+KLxfOV2J49tsmMr3+iz1HaMdHwwCB1GEkvcFRJZMLB+6xgMmTb
MqM/Uc5azjAaftnIDVP1LXym1iQ32D7VgJ5v+n8rZ2WjJj4olrDSczSKEmSxXC71
U56MUgujN/wqrOMTnxiawD6IInOWdN2OkHfw8LO9GYlMReFAGTKlgwtLIrTuG9FU
2GTnl+EOgVfTFH96a0k3qdUvK3sdf58B/L1w56sOMijH7QQ0ObBOQoXhguNhSw25
+gil6RDL3z/SNhvKlXlSrNUs5wkaBygPQnwWuKE2unvOluvl7a7oHiRAwx1zU+pW
B0QyLuLTAhTXTzb1Z6fnunibYhAHC2yskYtFcIr1GffHlNLeoRdv2BG+/AlJ+TWa
HWt3xoCDG+9naplXCfW3Eq/aJ9VuxY8lQqQ8dhCJ0mtIbW0XaTPMnrEby91TRPkg
1OTueQlne42pa6VIQ1q79sZ8WLRjoqO6rUpJDlMWm7r592YH0HUXKNXDbmXRR6kk
l6P7wF2Y4pxaJUJNyKKFlQK9wlZVmscPQ39UThNOoYyKmYJUzPbPHvP8Kx4dSRaZ
RJ8r9J8FwC4f6MNIOgzJKzV3o9ZbKu52josXyMe0bDMdu53IjxAXPOjzNhvW/jpM
TUTm21LCraYhaAuYVb10LrO5M8blOU+pr0FXtgNe6h+Vv+HL2gNGC9/9GvPFqnPN
8pzey38BZxQ3WafR3QIBL9HXtMWblD+63v3BwbLnx+La3Cg8716wTeFTPDv7rPk/
R/zRTtSV0IGMG//zhwgr99he2I4s5fKZlWWB49MAA/pRwvHepvWNujkMVYElD424
/IhyOS3lzkBJCewa8dvuPdqBrTHknFgTh+gIzT5U0WjphJbJYC0kSNm+DN5/ZbP8
1sR0/1N58mJ0uIBq+RC4ZlCZHyl8MPcvRAwR2zptvy7Ied+hocK6yLzc1/MH+vQu
x49QkSVa/GzjcHKoDdPiibKiclm6nRDJNFLiDQVw6JBPbF6VLi+lBIrSc0KynUqI
FDfih6d3ZJPIeNB/CRrrwar7GnFVkDRFW4ro6hkZswU28X2iPY3B0Dwbr98nDIir
ZmnTkE/sBqv/mtZTSJ5Q4ASeXmQcCatzmMlq6LfT6yDE4H80eWKc+jA2X2yLhc9J
dRJjPgf+jJteMu1tiGSzeIDoRFnhmINFRV/tcwu+7XT96qENmF7uIuTA3kM9h/U+
eK98RnAiVxyOZEo/0B6pThRGH7GxmPTj5yBrFFX+6fhQpBQD8dsldMMs3w2/UEW+
pCnfG6XvSUzP9hXV2oOasxdvkLSonqS8EhwVgBzYHqOj5jDRmLzq2uEtMHheu02F
/qxsnW8D1wxH+k6tXCNZHW5h8Pz+LfHS9/2Ji7vtCnTemkG/bgngd2YpOBjxaYFH
x4yH49zL/kHAmNvse0YOONuxF5bWSLje3jXyGujvaXRIQ7sKRSL4g/Q81oPI/E5l
nhup/z0XevomOQX4CMZiKvARmjs6/h2r2j92XXEGNw9U26IlMg0XujW6qmIGijY0
qR743dA26wnkgEvnVEU1p5tsQcJx2LyXHcnizkFFbwYqYxXTujlpREvgD06PniWv
x2uQzaMw8+PvRah1Q4PnhDrA/1oFNDt+lgNd/7FCR9W160gEl0rIfzkhye3+g5cw
iYFspkFGn1oGmz7fef34eXiRcd+EVMacuYNrRYGTCNZ9zVQLe9EsxDRAT30zLZgN
VgfZ22e+pyBVTOfLPDnPdeo5+pqibYDMtP+BOF7MUpTF58RcZgmhl8fzuTpzx49S
MhnNS+MVIeL0eStryns4Hr3Ib61LrszfbSQoMtRn1EaaNXyvU1snZtdoA2IMqB4R
MD9TEqAkJNkDWFhMqp3E09xr34YY4JVMt/+9rHslkK0bBOuKGoqcAiw7PBZDvA8M
MCkScfYpZehM3jjZZ8cVPxaCaiaj9NI/wMoVUhTADM1bXo9gcChxm+B7KNRMyKGp
AiFW7I7aHwLTcZT2lWjmVGt5aiDhFoDirYAbR399FoFWbtmo5sfJ3YL1I7Bbvd3+
AC65AmSMQz6QlN3745S8q2AWVvXa4GpWsARSilltZiwGh+1aBIMgHpfZlAWpXllq
lOze7GWc/u0lgD+malCbWoxSZbb6OO+aFd18TugaaAq9o+6t8aUxLXG1mCwhHatM
coGAevChwYtGB0QoaerKWOLAOq40epaqOkBlscFfBzhQN7tTAeTj3ilmc2sP+8V2
8Yvrs2uBV5XXCbSKd5HfKyQ/XHa6KNe4QJiYhn3Lq/R/P6dlYp1Tbuyo3lLVBwNH
63CuJFvYnsUm78FyZUuhgbGW7rv6OBFQozvSdlO1sdQyf566hf/flGugOtZr7SSO
YL/JN/FbaFw9aypw7IsXndaDndh53JWpG9HnIgo6g4mJi3OYJ2FJ7WxEtDQcovfs
YkxlFjI8s7vcVi1UesQTiq+/tf24Do81hux9mlWMjjjkEknA0/3vBmAhh+RraD3E
GiXkQLjE3TIOMbNmJS44VdHd7xjKqWoqRoEcFhaQdhPnTh1MeZJZQBUNs+OOgLae
JJrhTGBA38Urti7Az0FhOfHWRe1o74Dz1os6UR6KHm2ScEYi8vU6unQ/VkrlMmOr
BZycTQ1iU1u4MguZkysWKcMEIJwmThBuClpVkdmPanzD6hpdZZb/nbOFOVQzVPSh
xUVr/ZIO0jhzKKCd/LWOrruqR0TWeSOvxeL0NWLLdkjLsKMIhr19OGc8ADtIdKbH
ibdtz0uluU+KF3wNGUrjtLyG76sbvZ1jO57l5W9Mr/tlXL3JOd7mlN550AoJgBjC
EFjppiYSJY1ISYwbnPxsQqcB/95YAnKjKFZO/eeEpRWONidoaetywx2lHiag0KJJ
V0lKiu2igY8EAKMdqAN0BR78/Rn6AVCN0l5TB6YZxIB9+cdqEkscRlcjXiWBw16o
wJi2WcbC6YnY6HZ0eZ4psn7HjZDlUzA9d//SjtRnUHWPECOPKiC2C+h/EzI5g+V6
SRtz2HFypthGaIAQmJRRfjO/QrkoUq+00ugJ314q4rVz3qR9yozrOb80RKhz69KO
d0Z+lQIoK9/g/kh7OZB3yCZzlkci+6EJaSzN8v8/qBJs3h005e1z8bU0IT2fiUHE
7djfpLbs//cG1v/jxdMGeJiD5CM6SihoBFzBCas0HVELjYcEokfm4MLu6oW8pXDg
8UvnsITPgHt8UTVKvu8R2pOLw0GeC1sKX6PXqPCXM+gcNERQ7SBSjeY5K3j0AUMR
KWcB5FM4JTrx06eefUimKMQZ0j/ngzbDnUMb/aiRpq4L453eUR7nN8lqd17mzhDe
HzR3QM0VtXduJJDx2gAD50B7eU1tdbZjVuhtxhwSqslX+TdceuPXJwZwNHNVJepB
fUKilWxCNz0p9Z0HEp/u63mXkXR1sUds+SX/qUK2Nvr4KyJe6iQILQQQ9YS+I2nr
0A+wsRGkoxA8ZP354tpDXVt5ZrYJtIcKygK1a7ARUnhl2y+T40qpyuz0lLsNnv0G
ocQ1E/YXflvQfjcuBlzuntW5uZPuW2AeSajgLW4ATvKPVseG8EzfQ/QPaEDvTBIT
sAQX7f3KOXtM3UI6CB8bmcD5T3myUKPcK67MiRZh/PMcrJgqt8+OMmXGLvgiyiJL
R/JmNUvY+JQCn7ZvE6q/DIbRb5EueNgYE8lCX0q9/vDlTjCFdvleEAMLvMsmYoYW
bC1vOb3syk2s65fd2fwlchpccBbYbe/NYXCYHcWEkrQWPYvqIfC4H+Qpe9TWheHQ
EVC43p6DAexj6qHXdJgSezGsqDc2/Usrm2qn4uyK652QZd+1S3NFYwBfP7hc0mgA
NDi7iyYGTQrFVGcQK3sxZBFWT/YnHMdci5RIuExrO9dWC3FbMNDLWZxQfzo2w4l4
S7dSaEQIafRKW0KBLLyCGQPESztFys/8Ez7BFyXzb9uBtj6HJuwqUcCH9E2jd/o2
e5tzVfdD3hnflFo4hI3EpNyiv0j87ap7PSgDYlzkvofF+G2Ma2/ZCo4PJvk6eaUZ
7F5D+EhexZ026c4W7+25IMsQBfKGnLCxgFvYTGE2nziQNTDDTxBngxnjmVFEvFex
l/J1K5wsJHbl30GhvVu6LHB7dfX+HVcmi+2nYr86uz6UP42OCEwq/C1f7ephTDDx
wEYWzx+b8vP2HRJrcGqUp2hNFKgbeNMlfI8M8xLwbRujLPx0PsA1G/rp3O9iSyZy
bDNww+QXIbiIdQ0R930KSATWsxFAb8GhIh6X1vdIB7MrZ2zQpvOMBp76t6oibGzN
/3d/vOfc6Uu6XBdK2i0zTrSDeXyrFRmty9xE7QPgzpQLCfkbsxV7eF4QSuVAS9wC
Zq3k+gJLy2TTbaJo+G1THKt3yfAdajQ5nLdUrT4NHkEUyMTFVMSZraQcTgerbMkH
fd2MWdV59jEgBqIsHSRz6v/2tLo/vBDnDhU+RGEoHoCYiPJWfuP58o0wKVMxB6T7
T8YjFJQ4NkMBsEm437qHhsVY2ChGGE4frbPejXfXKf6Trc3WmLVq1kfUKjS8lyQW
4DWUEUBpZQF0JzkPUnKuS9aQvuw1X5NY2Ql6H+LDm7cOHHnS5/Vkyxyt+7itneYw
uqj/DL8JzjPitjqS3cvL+eTOeTi1wLXfyv0ibvWipnuNc61rms+CeFfj0RzNbm6o
r8NzdoDwhmZ4XFz8kPSDduJIwL8PSDQm8V51GDxHFHEZ70rJI5LQB2hqTpIQZG0v
5ZzNyX7eHyJtlge1l8iIqFjscz2KQPRabvrPHjmhkUuC8ouqadb2DoXhgjIpQVHx
P5SpUg3uBC3vyi2H4OKH7UMKWL3rqJV5Qa9lXqjuyctAZrd400HpAMNyXQtfx99F
puoru1EC+Wu/MyM9JpxY5OWywS6oP412kW+7r5waeYZVrNcyAL/IlUteGhjQjO4E
0+ESK4TkOM9egobQRiKhllJ8N+FaSikWoEK4/6cD1rezhJq3Tct3IXRmHyc13rbZ
SlCell+UD6ibTyeL6AlWiE8bm+rjajzkX239J4L0GhL3jVtpSGdBo/0wi5WAdJiR
zSBR3srEjBXXGgxw051ddO4HEh02VXYPi3KjXtL7/8vamgRH/PA5TjRyqn8vEWtS
FyRWZ2uAAJl85Ejd8usLgJtaUx/FDftzxLEmAiijlrJrmy7+fxXPHd11OBC3+Yce
9wqducY/2dssmpUx2x+/R2j1D0vWR9kwUF1ayqdZvg2DzdrDHEk/QquMU2mkoOqx
OCxwBvfn4o98YOc9TePokHHAutWxwROs+FcEbDUMVI7JkKyCkhE0XbXM6+j6PawL
nQ99Hkl8I+wVLP+Uer5ysLtsQj2/D9a1AoB4ALPrMeTP4o8//tAw+v9gE5Qzx530
j2d78WTJkTDRHv7qMDOfUh2MQQ3v5t60C4DcizBV381Nq5xhICOT0UNPyqCTMKlJ
LzNUSFDZlJkXglwWDJ5WsFd5aU4gJLKEzPo0muZFXKDdpSn6mIXbbn8Y3IQ0B1Zl
epEN7I7nLp7MTB4nDdSvxT62Ox9+3eUaJYiznCr98YZJNcJNSaZcQ8l1OJbdivCa
P1Em7RuPbCmO8WHSLBuRk89UVtrTSW9+uCFHyugNjxb2IvJgaSSpfKzbkQCejz4n
RvLSeqzAXhrQSvpyL//g7l8sGPhgMlYJT1DcU0Geh2M/kAEMOQeLRFk57ewMo+A1
mpRAO07drZOpSsdnGHxs4fwE9Vwog78t+aU6YG8LJ6f8lMHEhYlAG/6F2nTVLAS6
HxaH2C4X+uBi7/5FZzHUD5pV8rcZmvY6eqDuwilNVIwczFrxexkIQOd8zwsL2xuV
JRqR5hRAFq5MHxNdY94s4nxAYNK5CPJqFfpyWLUgZynMg8jom4OQPEWLFsrJqa8v
dwRNH/FeBW8XuQ5AX8UISIvSnEKF7dwYl2+gu8NpEsgjIN7RhnPPKmxEJrUBv8Ly
zLR8e0bsSPPraceByBxB7umzIqENCbNS2bZIIWRwxBoGNZIcDBEyCi3UZvGjJOHi
+41ZfT8qRONn2XCBgpU6I5X12E6IhLM/Ijv2xM+g0NbebKkzoLYzVDIjPopC/B7R
cKEcTx+fe//n0b3UhxDi2CaRiJinF8/8ewCi16kt+Vx3MpuxGF/7UQJmchauHjUI
AkyvaHaQKsrOgFNJXmEYho7hz9O9gTogOWF+wplwZx5zpspB+4DrnlmiMyWFYjP5
1zwy0XeL+VC49bKNg1aBX7bfSyvSPSjhWT74sUBVFQK1TVvpQBiMBzASuABsYnB7
tqqzQne189X8mC+dZGuSN+KFbBKVa83PH3SOrxC6VfuriE1ju2OnmWjEmTPu+OA7
j28VkBXbXQgBUoMpSeUWKinZCrPugaiP+yosCrjjgy2cDMiphy6+WEtIwep2Yc4K
+NXdl3Bq/dXc9jbek/DfNHWmQuhRfEzKeMuzcDzB6RnpVld6dqqdC8thjzks1GTK
Y3Fp4/LzsZld+4pQTeCsX6on0i201SI/jrApLG+pta0CvkAMUVpejNvmZPvmcE7S
1EvKnZi9SfJzBvdZaWIIzPxcyvQqWT4HlkBx7AZJOAqndzk2J9LJi1/ZKVr5uNZX
uYdyF4SRUvIIa1KnaFKpsVJ9Tw73gWCpce6zfrJyHQiwX6D3gxyN+0ceRszvJCnP
OJziyA7/vGFb3bMtst7+UkuwzxiDIlMwrBd0dKtP75fCL/U50n8bdDUijUmmeoDl
oS7xQqjS1Un0JqiKDzday8KE74lv+lYW8bo+rTrHDDWv42npGNZWYcg/Topqw/++
Vl3FphnJ0xNrkN+8yAm3JI8Uu7XloGLID6MxO/h6UeYzFxiT9KV7kjP+/n3vqidR
wPe5B5aSYwZCLtFdChBpM4ApDrDKyjgi5pVdDkAO8pBfVhPefI1Tz6S9eB3XF2fd
jNYhC5qdQqrWI2DoW230dQnh+sfCXTRFYZEy08EZ6phFlAzUomw0sKbrXn/FWQMH
ZB3oX6x75IYggh7oUSnfmLxklrtWyYaRoueDY/kV49rhWGq+tK7VRSg5cpSD+B/6
7CEExn+tO4YT/61emV8AMeYiPqqNmNlcdHfOJQqIe8aBgpJlQs/Et+VH6PHKoi+X
YI/lePuceHrrezgqG2SQrlSUOdHGtfLztyq3rOU/v0U0H9iJwtsfOIm01merhT8E
aaIF2lRaoxBC1CvnB19O9J2bhpu4YHEL52Grb7L8VR4bCziN0BQzaFj2OdaRF/8f
A2lE6jYw9ZdhWGFiW5nIx+lkQLfmWL0qA6gQIMD+l+J0muSaPP7lZnIusRh/jVJ1
HVj3FvATU7x2aOsZKZddocO25390Xnyb3WsZEnQyBVkq8AinhGJ6rXSIXWprl9X2
1JM30AU+6ltBm6pUPoSJWllx938rOeIS8amnn16ya0cINcpWRIwZIeNKxV0s7Gd2
rC1xGq1kymRmi34zwAvC4BawqysfZLWgMVA/9orqWRKL5B9BAGQhqngGJzXFXBgl
1C20a1uPrcRBMTg+wo2g/Kmu3mrx6KeShouA8X6pEzmrxo3TWjwjoABObANwXkJV
awF2VvdkfAQ7Fdresqi3lUpR+QWLV7VWNNkP1Cn1ylZbZHX2+M2emRNvXSoFEY3g
fXm5q0Qao6xIN2SJEFevTZGKH0TFyrV0iU+lRMROoP5mdw37P7PEkSkOOR0OGzWY
CeGNXAsqtHNRe6GtSRumXKnSAC2ksoVEC3Omz5ZdDlT4nHOTTKI+ejfTYwxXJYtX
mTSxUNEe7Dozm2VJAKgF+NAtvw44DEpM+nGnbhxGLZs1z7QJR84sDtwQcrVZHeVg
dvTTy86z3O6LOI6V5f2md7HycXZkgUurhN9jfCPPT8Jgv5P4B91N/VQkF7KZulEY
UHsqmUaQn+S1zz9isqhIRDuv4/j5+Ykd430Tm1ul+fsgQDCi/qFq+T+o8xybrZZ1
7Otxpq6lgdjeEXHg2onh9AYwevcekohxE+GrVsb+Lz4wBStCa87xmu4X5mJpqEew
KydtzYSytvw8yoou3u1HXMMhg/dMDCSACNb59mk7Mx8lBGEam6UXLUUwS8XWrxVq
4jk9b53bUYKHfAuyT7gQJTkf3GA7VTuB+yE8z5X+EbgUpYcSR++59n7z5X8qfIWU
JL/6vIaziup8YdZ61jFRloCHnpm6zL++Ck4IbVBjxQkXskazVPUU+JoXRSTF4w27
bEih1T4N8e5CZPdmM/0Ot1XEdytDVag6K4E2dVj1vZP1N0Syb4JewS5aAdp3oidF
lLXtRTlTR/c4NmDOfbKvv9J6ClPxjjxq0spG97Nwn9WApfBXQ+DjVFfxatjo8VbJ
K/e7/29TC6QIazLIXJkYwpnCbZnVd+Z6prki+cFZRj4AGupqzYW0wA7GGo94v4LU
ZCqwRgcD0Q6aFceo0i4P9CiHxpBjJFjKZoCEN5O9/cZdWCj9T1kUWCPk06vTJ5RA
OG3UmWbN6QuO544DiGRtu4YAqSW6rDfFLJUU+dX+tFvJFTt639fHJEziad13nwbF
V4alqPkUjAEFJBUCP99iG83rOCcWmCawLjJMwFRjL8OqgeS32MWu3rFIP0vnKStc
ZpNbHBqXdEipjPgR7MXYJ/ybwmzIfQi7vp8BZOJoq8zgJCVBpUdP5JGjFjWF0Pe4
I2pcpIZCv4Ixojqqqx/0RmNe9+sI1RxSosL4lOjxnjdMqQqe93hxJMo3DedJ/vbx
HCXsRq4+CqS0+U81gETpiz0L3PlTRXrFMFP6mOhcSRPQdv/k7sKoyKDz4HeSujUx
Ga3aRfz2yLYt06SorL1p8d/FptIHE5c1v7wmGwcdy3zjJFwoP08a8B67jBuroXCH
nL1xrg7BoRtjlhLkiUrJ+L0dxGGHOWTchwvmdtJdJ5lRYK6vV2dSdm6xx96tbUpz
oPAGIz45tUEKstzIrbQJDW8/fp4NqbLBhoRtYq0NzrB5i1++mmiuVIomXeM9F7HZ
h8GhwERfg4Ev3QZkqa+s4ymkAvsxmI4WMH3YpPWQbwfdDn0T0dIbUU1A49K4Lx0L
NCFNNiMxEIad13J8e4K9W13bSAQuFLLWhcV6N153wwVCc3iYOvZ++uADAMGB+q37
JDTPMikxcgJqsmLVoruxo7W08yTEI/iOe+dbQAmZ8AK9biNlT9fgKBaXoqdADekf
kiBUlQkHPmUSJ2H/y+e3UNgxdNyc1aMPmu8dkU5FX30dRwGzCX0lhTWySQo/8m/k
x0rmWfdpBBE3t2JiKKg8MhRz7Imf6/Vmjd1+pI0GCZovZzRPTgP+3zbt8NcITgbe
20D1JEw7W9Nxy4jZvbrEsI/2crenwYPnblNz7Ge9RW+xayfE3ooNer2bfgT6SsZe
iIPaAwXRCBAPaWaOmqBxLxSgBMSKQy4graoM8h73mTA1AyCHErf7unhRddn+fAx8
k/XpNtHCwzdO2cCPHf/bx4G3OjMDv815CM6RdV0gIvgQEiHqFlrmBSmq/VUbKf8U
Dr+ZsWiLMNFkfqzSoljJKckwqhD9rYMq345GLsubPIkdhatP7AX34TcOeL0Vhwm5
pYuffdFnwVjqEOACf3uxye9/1Q323onJ/eEcOsipEwxub64UeHRrP07F4WOegG1V
r9fLTMLxszCmV5t0eKvafxngC/BKnrjX4y4DFWRvIwbkL4J0kBolESgu6+FTexSr
1eJ/UbWpta5zx7I0jgceVJ6guBDhvjId+MKoobYJ7E4QDZv4pUYIQ0zNH9S+dAGi
lXgTvvQGv3VH4zjUGWC0jcHkd/tjSuHQ1fZxZ3bGDKinH93NDPrhNoPrEJEfG5sT
bmKHvVcSO9ewz5JaeiMWs3D3dB+TJxho3kpoFF0L8X/xRJISGKU3YzvBRx5Sq5qb
bQbK896/gMy2gFYtrP9xvpv+T7khdaJ/JWpF04IHjX0mXawYEdaUTC6cqeIA3dD6
7epZlAEJVQq1Nqn7nmp3SmCAr2iWmoWZGEU1P/d6E6w+0KRMzpY8RU8apj+p9Yy7
u5c8wPdqfJAaWFOgiANSE/LQxJ0Md1S5/60OPuC3iJjf6JbMVH7hLvjhzp1JGbFQ
Wpwp078g3DsxOvBlSNhVNiiWZPdMynllMUvphe92HCBvA+k2HRm3lYQMkMCGdn6v
un8NXtCLaChbPJbkS72WuAZyjjDnIsfTZiUIKnreLt0tmT6SpaYS+g5O6tSwX0fR
gnh4lA0f/XnP54uYUAagZyqoXkOFJfGAkz70Gb2oXLjpNA8GiZ7Nnme6lT1/TuYk
6gN2URZ88z9c80fxKtajSAdAeBs07d6vX0H2tuDCrtnDNXe8cecQZ/TSRma7g8wz
+j7oqKEYkDhLPowE1w0d9LTcaPnlZhj5zhL42KphYhsbUxXaKpBttdOO+uV7h6wk
IF8JFfAsWrlxoFxYtvQlu2s53XzuyEbJ7hPTPMigd5NE3qR03PTP/4ZQ3B4Wdyjr
DSxYo7H+mw4OpiplxXK/edB/w/h6f6DZgSn76ewHIThJR4kZJ5D6pMaLl1d/NkXz
AHQbAddc+z4vYM3WyX+tubdOjzieX6yB/WDRfzlRyVZv/rcAhwicH7U6FaeDPTMy
oihMd3J764yphtjMDcDocEF2b5qDV6AuHEbpiHRYL5U35TJAF+AQwG3RTmMCOX6t
tyFFY13i71dCJmZNbaOhpw==
//pragma protect end_data_block
//pragma protect digest_block
jW2Zb9hzqlvMvTHv6peSy0UfpnQ=
//pragma protect end_digest_block
//pragma protect end_protected
