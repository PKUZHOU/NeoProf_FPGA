// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
jVxSF+cHUZ5P2wOkjmMo/Fu6SBLp46kYoQjfHM7SEXTDnfZDteRLbDZSJ0hEV3O3
qR/wyT4Te8MyMdhwCgmBc3GcBxLiXgCJqy/YMIRp798zG3Ea363oViDnFgSkYXoI
jJn88UJ1VLEx4tMnFNzo2MjJ+x14X1EIL4p5G1tXSAWtnk4Z6KjXOQ==
//pragma protect end_key_block
//pragma protect digest_block
KhTVxaVhQ8Ez+saRAzx/iphpLOI=
//pragma protect end_digest_block
//pragma protect data_block
FUA8ngCvp2ZijKjeowb9VvX3rprOiRBktFVZaVBRePOMq/tMGp3tufgkqi9MANJc
F9SyOXp23Vbs4jizA/J8v0SO/pZXlSWlkuvo+blD1Qq2Rd2bt3QVlPAM8+CIaCaz
YVvbQAJSTnJV/JYbPFfqpXH4AAlXQXqWvbofRD2F+2LzIvflV6ztz2VR1aiuYYLY
VuqqjB3NdAPVBzNFssxsOq9js6qhmvXHV91d6YiJd2n6osxR5OSlI+WloczB2oGF
bFcoitHVFlAXpJ1bg50Wab1dycmnnxdN1o8G3wfsUSNdVWuISy2H6aLJLbBLYqVl
YOgR1xS+qMtDJyLVYlmDcPqK3aEhKKBlzh6eT9fifNWOljWjbtlMLMOSy5Yge5oE
vGyhp7hMIiifb4wC7OL4mJOUA3S4knDtM1TDL06Bpnah82kP1iO6G0TAZQYJIwE5
xgsI8L3J/elMNkU1L1PL1vKeI3okqFG9FHOaAucudayWFN6mW1eEdWNvxSy6Mt1u
Ca9hUZuDACkeCS0ZBPfhCTqrUIKCfd/s8HhpF2Oi9pCYjO/kUflmOrJTT4Wr9B4P
zt8iyH7NassNCZoR3s2DChWLZTGSLEAouWGvAOKLgf8toxzRZRjQceQWOSomC9XA
kkugaGHFZiqduasoCl1S0KjG0hqLaMbqyMq12BCs5dKqYcw47eW4Ei9zVMP9zH82
bTG9co4NFDEfrSBE31/+s0uLh0yBqAe68PkVlQzUQYuzy51uxF/zV1QzXq/1Js3e
LaGe7cVZlwdY8/AtOOYUBPzNPgYs8SUH9mjC2qhHjq7tJk+6zdgQ1AweU+dSxFTv
LCpuCOPC3rMOVpPWce96SvTTifsMwpzf5QlbZW9oGdHEV2HV3fOSnmVdvnyoG34q
91HuVu6iB2em5bGCjMcp4il6MWMNoWlSU8zktEKUC6ixaLf7AJo/PtK1UUcf1VXm
8V++TTzvAKK+UcjvGSNn3bRkdvCzf1fe6Konq1pOB50k4CmmLShsHK7YAsgrKh41
6icNdTAUhw4B1KeO/Dkuk1eYCnraFWsAgsgsY3xpQQWQ7nljzElJFtTm/A/+mkjB
MLJUiezv0SUjyK+r7IvBYMZtrzZdQWAHo9X9hvpIGEQc8uDsl7HsjSoSZjcHVNlj
IteOPrZq+69DGCQEnfzAWbK7Ull1Q/l4YhCw/i8lpV/9PK0yVvfxEeUamps7qtGE
bkXUbGQVAFL793LPPH3vWpfg7FD1+e1AkGTwVXMZvN0tdCqGW/dyX1APoZSiPFVf
S7Sb17qFHwyC8Zpt2SVmLDZleqGxsBzHDUD7XS3V3PT3X8htgpw6IjaQl+Qt/7pi
lD12pmIY2cFsxhYAQECf3yQCho3Z7ZH9z3HnxGDnkOvOx4mNCTvluWpMZHYosMWc
tg/+ERPduiIqjJNOcmCIjG8QL+I7qKxr4wBtgsakpcBPe53NPSvL3BOTUL3IzjB1
DTujwwae3AXYBTCfQpbwrkGRTliblitblETZiVs9PIC5PVxIo1Rw4EREcssEIxLA
vnwh+dQhUyRMmxWEVt70Zd0tU2/7XVzWhGxE39jCeaNAzXTywMqTOeOwTSmJ07Eg
9jW54GDYFW4X88bOU8BlBwOOJONN14gl1hMUN1AHzIgPO5r37Iv2sZdXVJsMsypm
ljKWEuXtv90W7X5WDz71Gz6TwRuymo49wwOxURjVfAENU1FUTiFazTJ11eIxej+z
8VNSBsR171fw1ifqPxTZhVCUZzdudpX8fwuZdpAupK9sKlrDaT6Kej6ffA/TtfVP
0HR/AeiMTYl2seM+K9preopxDc9B60lEbQx4ovOLrVDPMA4MF/lm5C94FGExrDJb
2Ftn2aWGUUyUKjEntnhyZ9EiMBHi2MdgzPaVEiNwlVLdsQoJeF+ZHEF1YNK6WIFK
Pl6/pt2QmdCU0Y4RPGDUa22BKatcJmGxUKu8qoMw+bwiXaV9PPDSWOPaKqGWt97a
nYg9WCq28Ui3evp3/x1MMfPy1ekIOnl9DRsvTul+svsGmDyIsYJZIXnoWPT1UjDw
3ojzW7g6559ceQG6ptAv2CQRtmjZvsSxFP3QLpm7AveD9QiFfcj7DPd5gnfjQHaF
j/homBmzrpsrS8ABNdSjX448yPqUczi4g0WJ+y3Bd5HNGN2hUM9oSfV4tlvmHIn8
U+LqQoIDbLdqdIjFlKUc4N9TSCAmnoQQwYxLl/EQKBDE43alRuqfIiqv8GME3j+Y
nckB+bde1Ys6IUz93KF+EHJ0K3vVYVT0NE3qoRDPd9Qe2nDavtK7R4jCr/HG+TNt
f1abRCjJMVKtgvaIfJsR76H361Pl4L1gjRiB6p/xccGhSgxSgnuEsp1+BmoLHTJj
7kGg/eI/B4cVEUCtwPavfmgX3T7ikkHyGv8FDHId+xvvkU0VkDCjze+cdcr9senI
yM9xwAO4fueyE7eW3KTOj40fPCx+zwuIZ2wqmsOET1TKMDMpu/IXFMrYKVgLPbS7
O3naV5RRls2L5GZMPY62BadIgtToshL6WQ2Gvf+y4Kmdycp+RT40VnKBP8mIc2oy
iH5QeW7eTJgsvUGLuo2mxucKuZrIBY8yhgb/+Rus6clFrWoAgznqi49VrLcdprvM
9vt3Al19nlixVd3xn+8Nf1MV9ewty+77YbbPyqjk6gI6eYO95cLuAWny7cUJVM5W
Gu8uWBE5BCKaD+sQfbpCwvntM8TE9GjOsBayetbA/kgWSRTU8B1TyiUG+Iog9m+x
vBEVcldEEmdq1n4xLMOk16deOODNkaLkszGRLNFLu8OfzgY706mACo9w6O9esIpy
olnGDTtSqJ9aR8GE9e42JddkM2ke8Y0Cqy7zV0ba/QmC/hp3iGDyvG8bK22447V2
uqrMG5pLUopir1mLgG/sSu8XK3r1pc82UmfvdBQQR1SEQ8Km0S1OEbBop7R+VrD4
jNr11y9q5EjIO9gaNUXwqH+PotRTeraY4BbpAxP+4OSOJn7qTHvtl/bwCTAXUuVO
a05umkBE3oROnu5/OPgJedi4C6+7qV+Q0KNw1EvXo8sZdNI0hSNdR5QSHfQT3NPu
yjA3zRQU3UxDlz9AOxfhfQ88v7DpJ5jqbHM9fZNmsuT3dpQ1Yz3IfW1/J0R+LPKD
0a2QoN6fJp7YBo+Hwgg+QaTCRMmmQmmgQ1Wtslerysp/ljzNxqv5U6YclXQqOhhO
p9beDds7N5dSxP7pcatxx5Orz2WH0Eg5SOYN1nD1I+5+fKavsiE0vLAJdMY+EU0x
bVSQM8s1aF+ZNiCuuWGg/RNwBmrS/DcdRqGzbO/NYUgZmj4hyl1tu2+hR3OlD1KM
6T0o1mAEiP5uIR0VU0NHNtcCyeASWxWlhYQASGdh5RAJQ+KzrKtZL5tkhtOdX58S
MSJ+lK970hPNQYthu5yitBM6XMJ6Avk10+rpnHsdHzWudkOZiZ6K1+D0ktGp7uwi
0Eq6TEFV4/dP2mdwSSu/binPbGYFAyMf0BAlj5SQ/qbKSXym2FuypmcDS/lluEpz
sOuCzPESOYc4/t0zi7SFj+klXbBItRou3UxKRaCBRGm/D9LJFQh10cKbhR9R3yCH
rSgK4eX0k/0tF/B4pLiKqy/tCMXl6m7SM3ijrHRrmvLyjRB48tgI8uSKtvpcim/T
Y/IRrPkIv9ROLCBpv9yEYZdrUJofCT+39PpQpF5yWwe/yp22Qzv5OB5TMJfGfOMZ
sPzmT5jzIOSPp/FlbKPLQZs0P+C8luNJHcDdagJjVxkbLbME8DwMZkHCdY0gD0Lh
dc8gkFGCKjvU21A9onAArYtuq/9hgYqLBXvUIwTiJBlplvtVnxYYxljR8agiPpDb
uGtGkzjydXhgG9Z2d0R9juAH5JqPpfEeXfYwW07SOHc0fUJXelx+3q6dpgQpwHSa
3elBp3uhLoN6WluLE2jqbqvuArDptxMKtMu8oAuQbdDVGMC30Pa+ulsjIsTdvuw5
gn4Juqis7Nqxoe23FmpIYGMEZiMiiX9MVaFjdLRZYfMU9C5xmtwW88JXLhb9Wiuw
B8kcLJCL3AUK4/Bt8ZmoxRy+52tkJSKFi+UTi1SbjnT4KdR+0SWh0iXElpITGLzi
bcHiChLWrXBQby3WVsTHAM8EGpmDXKJaUd0gR74vOR81M8m8BgLCJ4q5NfVlRPUR
EyZSCATNEazdBTaPsLmnAgVhZ1+p0utF/MjvbexdaGiWQ/CtQomVBkQQMklVJjxK
PlJMPqBNhZLPPCKq+tu7jn0nBt1IIpbkQdOQxZfyqyEWOavuEuj5Tl3iTQ0Mrv8O
UBmzL4vKuI5a8E6NZP2bKR0stbpGs/VAZbcxUaSVWLRIamiJjXuYQGMOkP8jM3xq
afoVjXnmy8mhc4l6siYTcvrRWaLfnrNjaTUh6gj0Bd6wEC7M7hj03T67t+mada7X
pC0pudfhG4mMJsljF2xJ1KzgK5ryt5FLhs4RRZje3u0qRf5VkeJ1ysgEjagpT8Cm
eRq+8onLaIF4esR45HatcHbPMnp43ayc2QxC7JNQP/xHaL2+V85cOSG2j5vYd9i5
qtdD0A7PigRQKxlhjNjXDhL8gun7MSDhd76ZwbaOyhMhqeHZRDwNytTwF+awRWEC
GKD/vcPjVToiWlXql0bgJhb4Hf8NGuhG2fCgA7K196UaiGRtmHZdND84NJOujO0J
I8PKCXsTUZokCNW7XQKvYvcGX1wpHuFFXKmIKiUo1KaTnGAzBuNQSo2ssvIYmaAd
CH5b4ovtPhjae2UZjILT8Fp8srS+oQeHv5UkKT3lboIQQuD3hhz2IDwebmZZlesB
L5wStBF3YXgbUT6Msxm1ZHiaWo/1F5Ut1iyNKhGwKVH3V5UN2ApM3xUIFiTwfoiH
3kQrpBsSUOKiY7BS23xpMy7/3zwbaEdlTnv6EyacLfp1EhJ9K4+82eSTqIqXo0rU
p/uqjF/C5ELrElJ5Lfd90w984qqZgg5czWxXhDsulYuw+GCOYAV+p2/NG9Me2kEJ
OrZit0UGhB9RIi7eNDUy4Frd8ZD5qzdYnc0/eikfIPflxOY2in56orCJXxCtIDia
YLgVXdRzPXaiwVDqJIKWUcW6ENwq+xFuwasG4YuyrA4fNyt/MNTwOS60PVeh0pAp
901GNNouCRFMVHCbOUVVZlzd3QAEvAyYs/1vGR9p6xav4JWk//C9ux9lVvBQx6a0
rsJpgUHiFfzF+ncx1NT4RITlMc5Sg1XS/ZMLcCupx5XfssQEmE8MaobKxOe5fVvd
8wcKkTSORYNa6mA7SJF179mKRrXueYHAbgMfVF0EAVwn7vDuYokqvdSfFjs7D8QG
dTSp9u7vtPrE1+Gqj5Y3N8WH+XUeiM3E6JMZktQOyD2As6B/w2XHQ3XEHu0z1DYo
rJA8Pvt4PzWaYdsxkyko4wQXNrLhTh90/LQZPiMV0nQz+FZhzqPqwXR7dt8BUh/E
/oasEB7DKv/voHe36M4mMrqlWGVD6ZCRQONGBWVIftN5s6wJtU5lP2k/XGcJJGsR
sbLQN+36a0QJ/mMeFYYruMGY2mz+y73AWidVsXXlunrQkF+a/OPnK55JSBT1vmH9
GTMyaKUx+A0rX5vP4TjO5Wh3tejgd+gaZrkTJ+wxEL8AO+B7hnT/0tDSOaUeC2Lu
Y8EtpDLaCpfdyy5L/fl9/3gukh/JEWKlRVBmEhpIcHeEio7wMIEKk+rT9ygK2fds
A9kxPI638wQOEe66oNtcdYGWPQkMh8Lq0VsctWCASQz5pZ1zVbdlICjYm++J3SX6
DB6NMRD5cIvLP+sg4/vDMc4tpecJKvPnlwRNA3uzCZF2YvdJp5XP4kxqFpH7ICt5
WqH+DR2PjUyw+1Hc7O3KW7cYo20EaRnkHhYRSBNa7kxcsJGgSVTfmFapDS8I7pzs
kg4kRAtZ72ouvRyZkG+SwnRpkTHvJPPXR5R5O+u2nWeVSUDAQ7tPS+w1+Pc5nX0G
BaDsvMRynw8A0IBZWfXyVVIfKN1vY6GACa5MKK6+bAd+hyyvTd8ebOHZZ0fSGTIC
WN8DEkDs3ABL4bYrT+0ivdh1OQ89VJHPr+iMG92cm31vefjH5qrIndIu0819PpjD
AgWXyVDfUoRpbVul3KaNjuWD6vx5KEPtM/CIINXPOaEc3gsWg48bIzZ6e1+HYNcG
uyKs89Z1SQm9yc0D6wwEhTKmh1hYdJTJ+Ti1N4iiALja4iFFqQ5pCRdrJOVql001
rhMwxFRzxwNRtl5GwjUyc/FbqqrVyhpOQGVMR2H62esq6CWA3vxBgOZ17ILjEHDR
aTiUxYukgTdLsiinO/BhyzZqdmtClSvN8C7TFk7UaauaQ/d5gwXoY61cPEWITjUr
q5MwStFNQKTaEZEIuCWQKXxXkRwr1mmespCr5v5tzDhXwFdvKdAuXR8AGhkxwGYz
m3rr+T+fjKs4brq6yXvHQVoNidYMRGvnldiNSzXMVH61dTYWXvEUXFyLJgkghvZ3
SJYQf7Y+Y2Jhd7acwDgPlGmdmkOg/SvrANIpwbTQirzzv1/xaLo99cmpaLsm72LF
6v2oXODuMPLdWMaL8yShYwlRDJO9H4rbv2UNjI8oAvKeZJBAloOqMHaVClu8uKx9
BjI0NZlaQsHwdSmMBRkeiHClMJVEPSIEH7O6KwUxFZ4Ux2keE5420+B5BJ8FLGUD
laPe6//6Q1oatNP7/RiSZpfu1uUlZwB/spUaYxTPgDVSc3WgHs+f2eslX+oVPSoD
RWJrherbxzHjqBdJxXWYw6M9n/zYzXbzhbgsVjKD8YVbf4UGqmqgtjpZHQXZqoGn
zvqI9s2W152G+L2vB2+ihH1Ey7rU2jOx7b8Sm1fWbhfgx2JiZ8Q3nzB86QQk5YWH
3+u5jln//BvHEmKJcEnTrmN4YzKIYxSobMww6FbgaSYq9QFhRZi5DbTZJ+5EgMOn
d4idfWCyQHAWz+ekTuRJSe4XJoIYaoxXp3se/bqNSYO3O3r8mmYywDZyvfVM+Q1a
EsoUWBvy3NzxXoi9XE2Ps9643yReZMkYy91KeweMqCGOqxNvjK+NsfcWq2JGN1Sw
QevA92XhS/ucl6fvlw/phNBvvfdbZOsH4tQWQzoZirsAa4WbX4JpAJf5uLFtmiEB
tudD2TB4zahwNazNlc9ZKJMraW/nlE9uEpp9GuIi08EL4vUFfdnPJfJANOuNGE4X
i7k8gxuHCuHEKoCwYa9CHUJXcnISqf7kjobS4c0wjSq5BM1053EGqVZL0F29lV1o
IUrleJPwE0Khu3zjEOWKm4ovX7yCJLUYm9DRsuv8yRA0OWxQMsrTHfU5iYCYixqs
JCYC7eJmoPARrdM3lL+hs7PM+aHo/eNlIU6BysvtDbMgg5u2IMnzzrBOa0eonPIY
EYp2fzsG89SoWOQu6btu9zA3ZdA99euWG3iDBZHeGRq+NfHo5iB39RQDUeh94g+A
+40zqcya5DoRgPQuoDWKufJPec/tktoRbfx+NEYl5GZQ8jJG5nmKXiYrMmrc2GxS
lqU3hM3WgioCcpKYfiE32WsKUpA7sq2OQieoW2dLENd+uttUNPHiz6J3MIsbMpDY
P+p+O03lT1yceLT5IC8lmPd6Gr0GjqnUZBuow8k/i8DC2KzIBqESHBLFywQ3lE7N
Jq/RB4UCsrTh7Vc/PlepbB3b+BFWm7T0OLmda3qgRhVfkmUIzfOLmfd7TwmMFJLK
IcNIpaRwVAUC1jD1qthcbkKJPR2sg4y+T+x0hS+9w1NCI2XVXOsOiiB1yPC+Dm5X
SrP8q0cSb4Ugbh1Mg9UbHyFvAUm5pEo6Azo4tr4ARPH36TLZESh8dXfNRaU3cPL3
ltPip8uv5KJE2vE1QuAu/O8UxG44oTvpwGHYe5RRueXFMFs/i7THebbA8qXhZr/F
4WM9SjQ0x2st9oR3i/En+RGHTeCRjOcmM9404UkeJxAMVYrwTFQ0KbzfWvLBIOy+
oHoY2xuCYtpfmAqVFhPmtrTYS4up+Q6n+8YfMLHT91spbno8SQihK0Za+ZLJYUlW
GOE8u8q7H1mVwOF+JPM/F4mniGIP7Qst/OKW7WLGxo8dPvzjGv6j9bbRqAF+2eFd
L78OTESEN2k2+sp1Vzhe/NQRsNej/WkNLqgM6+uL2ts7P6hSLfGgt0RBk+oJPAAs
r0iMVan+OcBlg6tKOrbPPfJbcGSdY2ayJiZVf7N/SEJyYbQt9/8wwqWl3EF6ImWY
lJR1SKoJ80vdI8rLJNdgePA7OponbZOO6zH8sKewxGZ/ogLfZWY3EKtWMDlmxNTF
FobVqBcAX1zAu7g0GHqu2DYrJQQa1dKegdV72vkYwmSKXKqcjx2OkHJuJ1hERM0w
cqRPjwZL8RuDBpFGghIrwZ4fZ0h/f3ebkTtrDKfwX4T9Jn+nmQhADvyaH1ZSJUNI
8C0N356crMwY+Tna9WB8omYlQzzAopOX8Ez3bNaP6ZGEmGbftKI92G3dKLAc/633
A4uxN3hx6W87hwIo6PWN7CMqTkImwbR/lp2+TNOey/EV8xtz0/URR1hqvPpTquoM
i706jHdxBPwqkdPdLs7pkIaU3gSeEDjvMB0cLnXAxq1Z+9GaEg+So/bw8vkXbPf6
Fwwx+2uHoiswgOXdL4/7mjmBH256d8aWNsk2wYo9hzziLibfbDW3euQnZSsxqptt
XoZY8eFCFAOC/Q/iJmh/6pv/ZY4A/QfmttY8qBfNe7o8tOdaM26tIKc9D+oPNiAm
X1KTngQtX1N9Jd2tNektlqznscHNxS2Xijkrn0Qu2h9z0vAba5zHXRXCbTe9p/ar
pKjS0F7u/XH69gZpuLy/l+fbwbm6SAkxnV2PNq/EEivMVJBsVdWsmvBzn5TO8txD
bLH2lj/I21+C1sAdHG19hapJMm3WF3ngjXkBLqmGttr2ftlJM/LNtUiDjTceNf/4
1kahCZwBxSiXeQaufaiCJlW+weSQHM1wvwwiFuwC4mt1vjbSv6rSO/lA2/XL1vh3
mNMDrr+7YA8JEa9CaXSR71b3r70I+VibeOdX0cvprxYwKxD2OM2MOGsBw7GY3KwL
3jw0iPLmscL+AGD3otMGcDlKdZQ95vP4juTolkrxsSqjCgeNgSBEV+5VausO0get
+mnN5X/a8mP7GKJxuEVLHzv0bn9gYUrpM7mcmd/7sWzTv6UPEB4uieBG0LdjV3ef
oza7KTHsxJdpV0RmOFuiocOSSRNaZv7oLVYRdKI4Au2h/qARIX9nl7EUK2CYwRwk
LaYnPEra3j1Ki8wW3ZxlM+Fp1NS3FLsjvMweVkLovWsH2MAhvwLtALvprrvexWlE
w6vplgqBmGXP8UruqtMkiz6dL22kyEUDdKrkqHTi3UXzDPgcBPOOxuk+fOnd0ZVH
CFhFSoEMX1VLxRLvYhlkXTJ3zxw09z3xIIZn2OTVgyGhze0da438ooJRVZTRH8It
BHJeY0s+bsOTjEZEiZOKXKIGm6edPzF7KURj5PK85fV1QP3khyeF7Ki/6i5orphe
K2BWH+N3ZsVsVTEDSA7tZdhCGrthrwW3cRC1hUXg5aaCKDWhP1+Q9ERGSzZOwqat
O9puTqPqif/Qkyb40JKjOUXmvNDdk9vOVA0o1+6aqg/L64pUG+LWldpZnOuB5tzl
Sg84YoNJ5qF4ZEnAMztQPcwoExn5ZgeTM+xrrFP51Y31PxxCk/AgXiyb7gvYhIJ7
qNJh+RydPCcXmDeUawTSytXqvYRN0HNlHfNUXs4GafX1pSa28qLz6tPc0bTaua4y
v7Hrrr7E3R/ej4jumvk9xDY/EnuZMs+PPL6294gq0HSHmm5vy2pinIwRU/hI/x8s
n/Gaej6C0l9/vq0QRCdYW14P3CYqX7UctKkLkaNZtPDB3gCSJrxAM5DNtIEFAcr/
NwX5GnBPXZ3QvxRMKUEd33puFRl6jyotIrs/uFv4a4dZLg3zFCZT8K5GFSArJIjY
UzEnzrm65Tl10dDYFXaCxCGHbBdAo9EpQNU8RO3YTfXuP0mxQ9cqI4mAM8+kzk3t
y6b9EDhOQ3FyEaIIKD97pgNr7DtpzWqGsmtRNdK06Llfm6koqb1OA7GJ2f29Dcw7
sfcd37zyHfZtzskHhOntJyb9hjBLpMc64190B9lJuxkIPQGXMtqLKYNPRKu11cG9
AP9KBMSH7zMIZJwHeYRTk4e+R91ITYaYo9s3lohNUD5jOuzaGcElnlHasIyqu7la
b4JASZw+hlSiHcPJ6H2gHHmoXbsxLEUoVOnJZy3sjbyV2sNuiEuczafS3KwCZsIE
NSykVvor17tzgHLTM49abfJv+FVTSe97xNkKUtsB2JgFbgxuz4OjZtDfOvLzWx9X
qPbTcVJiLVuZ71Q8ihav8j9lYjDn1Er5WJBaJF375RmLcil5r00cNBG7zRh8VAES
Mb2CCSK1xrTwV2LFiCWdSdYmovKmSMwTUvj7TELt15YI2wrSdfgmDM6pnt8v9Y8h
lHtikHMkwxIS8Us/wBVuDXuGn5qqVA+2z7fbk5EvVxUk1ttRwdYDBJD98twzRxfv
TaKk/RC4dOpA9rwL4CRBD2Pnp/vKfx0es24oOfBwPkIptU0aa89OSKImZaKufp8a
1W80vzlxT4/wg1Pg2LwkpCyRtwukGQYfaveEeskbT0jzcAMgGWBknvDEBoM3HavP
YFTBGmRWkZXu19GT+vVOC2T0bZcVBscSVbQNvc6Qi+UEQ44rFcOo1we34DkOF6QM
nTIRH/di5JCswn/tXFqeHNNi2U5NA1dNEKCPzensSrkkEio61ZqtFEQijE7hES93
V1EqA6MfWPNp2ajpTfdf0cZoYwDAE616QMgV81QMXKhSCvNUhQjLjwTJ6Gr571hp
fb/MZauTqr8U9ox4A3MS1kRgdq7L2LV6thHF/pj/FA9uYnNM8R4I/XRRXwAd2CUi
1IWg9wR2xrEgOpvOKXK7nXg8oWb5RNcmV8NjQ9n9LzQ0HEyIH5aHHqP2+vTdx9CS
+Sdy0fi8ID8PvpE7x4UDKwJwmQawU1f1/A5iRytvgVE8IuukBUJDlM1BsL0QBp4k
hofbWvqcF/o47vQ4McjF2j+H1FLMcgWQ5Q8y/laBO6iB/ilgVbeqPxrXPHcGTxz4
fnhi0JgZfl5LwdSI+FHduorK2jHdV0Rl4DRKgcFpIVZiVYGaDGnsJbmhXghsVWnU
IEwf/Uv8FrvBg17WDDt9gLY8FZB6vwXLxEN03aNzdduiREqmZR3u7KxjoQ1OnUPk
/RXLEuI48WTy1exm2+nZy6Wm7L6Mb6qk5ZT/GcASggTZ++BtJrFN2DFug1qopUwc
AGEU4rlQJsfHLnoq1oEiS6AGqkgBJdbcpPGEVsez11WGrb986HUhwPzdRG+k21xZ
KwnaUIqJn4ocFE4+b1tFBfJKwcgPHBlGAnf9IoPASIYkErQVwi+HapGgOUjUfNER
x6SZZGk+pDMACggex7mQn4+LWKNzXEPTsYescVHjTB6DfGHE3Mbn3lZQ0iRF+SrM
CCeAQ1VtSvZ+aDEywsB3MIe7M7ouzDKxbNt0SK9/+F6evrmHYm2L0Xev8fTWcuzJ
/nNL+TX0r83i102hvgB5+UobYQ3mT6n1rbYoQMSsYx/fx5yKW5ByQEifrq0FhT5/
TjV/tYPsXno0wwE+q7FzX3q41a1L/JY7nfAZ8+Zwobhr8/w9RzifwoJeTwtpBKBl
dQErNQytNRX2jLBHFiLlG7IcreLCu6OP3UxapwOWCISyzllW849Wsgok/aB3Fuii
xob12FvSbtSIjQ5JylZzTaR+JfVkD/U5+5FYSBGbY0lUhE0nCj7bunZ31Ht22UH9
dpJs9iu/C1aJqbWj21x9QoUmoXexdzBFbXHtDyWNodoY1Zq3uMmHI5eQJQiV2v+y
6FlVeoXuezMGiC86ul+ZUKEyoEqWTIV7vprSQUwNQ4+YTo7/kb0gPKHstGRedlGu
Q3j3nho56XfdXjfWRM2GJNFpmQycxy+EK5eKb1BdXyZMJCU2tsngUZt8JUygQW1y
RKOHng5QgJzhx2hENfYZv5EPnxrwFqc3rMPZO381Mj8INJQouvZdDFDGsXYPpLFR
3MLqjljqxeFkjYn9C6NtQaCJWhpa3D7Zae9QV9OnEJwx7E7E/S/AxL8O5CI9Krog
KrjnaN14mjghZxe6MCI0psiVVu08CqlPww4MUOFES+tR8jj4nLap3TeCz3kV3CdA
HzoBcqzb7B6guoNI/RXZ+3bua9eO87+YJiX4O/5wfXqsqjKQVgyCVwBePOpwX0Ad
LiLVuzR8Bsw4vb6UBGZEp1i43dU+lSisyA9xa05mvuMefSthgOixxc3pJQLMlaSl
LcAWgrG2c2PoTUlHhoOWtRGKYYrAqdYGG5amu0X2DE5VvexHXScrWxBpxeq9h2LJ
ZkY7v4es9tByTKyNJiUqeWeQvA7gIkEap/e8OP3UEtKruWrZ0VtED2Vl8ir9xtla
XCCoKNNlWwnGtDpahPzUZpZXfjKu9RwmINnUjXNcwkcBC6c+rh2jpC8Oafc759rH
IkG9ZxmfaYw/JXto6glWcvk0RFq2pKHGliBsk+fF9nZZwzpSm2FWkikBdYMdUb3p
xbmjzfMWeE6npl3oiABvxDLd9ZvdHDNSz+7eiFocBEKxnRhSSLFw8q6ckN+2wWsj
J/kXN/5RBKXZbSJuvg065l27oNoEcn15Qqu5pBHZ1h7P0Q5YhPs4tgxsXv5oiZ5c
98zquZG7CSCVCWE4q4Bq9MkM3npvetMAwiJLu3N1SNLbC9XqgbZcYskA+Ue1RzRB
ZfQCqELgchU/yd89eI9ySy/EKL1oLSP3dku4Bu7o0m1l3HGaI6ZhNmEyh/YT7Su3
TgDRS5M5szy1q0mEtXcN4V6nll41z7SLAtEg/4VU79eW1KHmhch534HzoMsDZ7ds
1HbqyhJKcNVtRPVwJa2pQc7+ZzJ6356XehmK8N8rYCgu9Mjyc91WPhMoBNC9IBZE
kmnBswgQHRtcuiqbCtrBcXlcdQZiPSeNAIMWFN747Rd8YlQaQ8dPLoScuTL9SfgI
r+o48j0Lf5SytZ0n4aOZvTVc/Daealn9cAGVixSTQgl1gFhbz4Z6HzqShxyZz1LJ
YvTc8hkmt+hz9/c0BzW+gfSgZmXcAgUlU58p5ygd2niwW014pL8LL4opcwJcIEwu
tQ8dGTuLI6s/3i8jSmxskmcQRo3/Tfj1lFV4lqyIzPOqRH1TSangA62rlDvaP9s3
D0JV5Aht6ZPRGMDCanM2/glgrdBQnUgg6J2dULzOAd/eYBGn+5VCWDdEviHnEPVz
MlTE9hv+YqRxwlpNDG+3Rl4lvL8Rs5wBK4gOgQtx2gT/1BFtaZhNqfOwB2LVmu5F
U7l2QHM6L7mVClWYvZgNh1hNjpyHrAUGlABH786tUvoC8amQLkSKL38rau+syCfr
0iIBYKd55DqgcCn2HUOByU7b+BZdQ0skHakQ+o8VkHHQMWi8VIPtpdFEiKGD8JMh
i9TNQ9PovTlerlbQZNCQg9LEpnUigZ/lRn1u8+RaTB7zLicG1pfFmy9yjx6SYxR9
+VOqy7IA0ctKDXUZBdoTAKSZwMkFy2p/9zhfcaVdQOhwBacg8UwJbl7RNMYzf5tI
SbJN2P+6i2Ddhf0y84K3u7QrsnzsJlOeRyxMjYaBNUT+KGT1hcFm913p26bJ74N7
cNazl7A5yN3LY2KASCyiOzH20Vap/3ei8ntWd2han0NXRWpDGuuTsv8ChlLYcYoL
y0GUk86HA/9JKhgj38ZJ9285au9AzyfZVa0KlbELUNahtIXuDBjLLweWsJreexGy
RE0SLV1TY+8tXem+XrWMTk3zGOW6nGMreSbonLGeo6Jqu9yySqCDaDkScYj8t+aw
Bt0YzXOyIYsgxQHBZoUgWsCXi3OHaB/VUxbWQrTjhpKvOQPA7IC9xk8T6mxSFRkw
tgSy3L7S12L2PQHlcIxncQ9dNpfK7C5/mxFATSGbr27RUmR+dZ6zP+twXNrf1Wor
GOQn1FycPz1nLPJvMiUfnb/JP1Blb08xQ223/R6/jzjdqwpPE9b3HzwscnGtKol2
hYJGIKggMLnve/2eI9ZS+ZVuIyjoDuqkjN1NEp94Rop6kqcDMLuGSDAA4W4EJrVI

//pragma protect end_data_block
//pragma protect digest_block
FqvJ6Llm54h+V0U/r245q7eNE+o=
//pragma protect end_digest_block
//pragma protect end_protected
