// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
j6MeXe1UUbvy0XBr2K5IDrDtckvhaqXC92iA31UgBKVUCHC0aDXvDyb16XP4LCiL
foJlbQWBybBqFDnm1j9CKvTmpRU4RJn5EcyHCjIBcM1MLyDRp5Z4/N1fmHxwjkv1
ObtxsNL76JwXK8L52OyirOAYJMtFASlqmfEna5GR5xk=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 4624 )
`pragma protect data_block
BEEWjqA6B3BjECsTx3BJNib5/z5LDD+fXMTZl4qJn5L1Dmh1tGsn25WEsIIO/RR2
Bjh7K9Fn5rR6FkIDZ5zBidCz1NsjevHXQx0EpU0aT6UEfeX05mVWUEZ6zOJh5TJ+
17NwfzxTpw52WvOauQiVxb1+3Rc88HkvazTC+IlYjDa+SirJ+cx4la7ZwUs+NDhN
8WGTzsOe9eAMo3zSDbJAyrSdAKzl6TgNKJmyN5ZgRQUy9Cm2cSWa+mMsrCpk4XPZ
ZD62Z82wPW7N7pO3vHTdr8LBmCglrwQ47OrKu5K7oEIhaBlW8c8B/tTHoH2e0ZoJ
we3LbBtXlFNLWjvGob0RsOtLcfJEg8ow9QP7+yEvLvhUnkiaUj1amMOwG4tkx54E
kLRDwtOBC/Im/yG28fHxIvbd5vJHvDOZjrkyN+4UpvN6F0qfsb97BbpZFdzgxIhS
/exWDJloT6Eokj8TcJTMjr/Tp0UD4hT++xkEzY2lCSqI1394c1hJJS/QO5UvX8eQ
RqxEykl0wos+MguQOVp6rhQC2qDchAbaMx/1xmXGjmy7K4ZVdU+oBXFAP9v+Yrgy
82UbSTEsUCs6R+RupoSR1PypPC/ECKtnfAQs388dterFvzNlVjUzPkKenatS9LcJ
g6exK8PGWvvBlk9fTKWLUjXJtHRw1ZHQVGXL294j8+TwsMevVMVkcs2zPrEovoWI
8/9vbRNDw6g8QpVC+QA2iuwfCh31cIcjVjv0j3yOJqLBj4HG66PZc5ApAZy0iDZ7
Sx813ezbsAMS+4kQMmkGRZuRBCBRBPM3kg3R58CB90fMiThfq4dMPZe8yYiTXpPp
2OunGjqBTUfevdROUakkitXLdXrtVGXe+9p6+FPuPJVPGF3XnD7Cyr4Jr9SNqzWj
rjSgYStgh5KA9kiMAzKza6r0ItL79ApEw58wZJJ6RRMYQikTVbxEg3tivX8YwVKW
vwxO74YRwj8uzXoRY+pdNi464MdRV63T9mUyzWYewENHirMt7vttLxgZKTOzYGsj
WEC/8SsKKFDQo4tcroNvIxVY8zWBlChsd13JZnMvUMrx3OmKi/4AVGxI5GpdN8xq
uEXz9+bcW6oQ13ht+LhL2/BLURhDI5P6fNmALYdzLS7v2xKBCPLPMmyqYyAOb5DT
mn81NxHsEEDbnPkoGy+GEOPSn86vsOov8LcSjIO4WFkNG5uBxuHpxC5Stzs7WQto
3g+d3uBshNo0PPDIXbzpWNNBerTvkm/vII6ieMDv2/UNCtYK4KwvixzCB/x9uCpn
3gDEHUQ3Dp6h2+jLve87p4uoymghldEVVJX07SYNidVnAXqOxP3soh5d4nujUnH6
IEKrL2n6W213Wn4oQ+dNrRYGmw71yDqO5/Xsk2BGX27VJLjvDK5vrZMctyto+zhO
brAtkKkLPQgzqCYOaJkaJaewe4KRAAzlJJTJ7WlqqwgXfCIwE+GBDuFUm2LClbXl
ne8dosmfx9rsS1nbgq7wPyJQHc4IDu5nyChVWZgK8Llv5CtDHXkMdf5BCkSp2W4M
/ewzvl9rCAC98KzYVzPIg0sITv4nure/r7QS6Gyi3c/d6HW7gipLPwlQBvQWiHLf
cSmwMvdBkzfFCm+lCxPSx8KdA6kEfJGDBSgRjD9htOgUn6OqMgdI62V5acN2Jxuf
6Mw/659qe4cWMv0cgtVrrvsg6DwyGOMHORRfOXC5PkTN1JdSA9Vg6T+G9D0ExaWZ
RqE12UNK3E2la8pNh44cnSJzTQSqq+XXPDgw0Q1JaIdsheKx/jCbY2YXXdo7c6a5
8dTcCJUdPBlSZMhs/OieJ7FUz/t4tisbwJ425DJb4TknZM227bg+DRZCO6Xjivae
laTgaTD4MyHRrkLpeqHcSPeIlR5aZ4BeMYEgXQVQla+0bzYz5eTlupGQ9UKFXxKj
tgw3ZYY0n1SsS7VwMPGWK7GY8BfDsljHdRGZLo3+2vMW/aHvXQUxPgPZPbTQrVhJ
uNogtWY2AGRwLuSKMQ/3e+UF/Q3MSIDsyCM/jqU7PU7U4aajS6rB0AJOX3mNoZ4u
WWUeY/ME3dNbTkoJdYDIvGbcGJTA+dXb0uIM4vkENclVG019Wk9C28FRB9tbpzQs
uoKPUJCDMrGcz4aR2tpbxvd6bO+0t+Y87Dkw+au9AUORi3kA4XK9PJ2p8c4VUcxV
eng5WNkP1Bbk0k4rJ6AL7IoZNzmkNGtWeZP+E6nprc4VnlppsbdQUN4id8eenwnm
oaxd56giBy/YqUR8yFLl3/KJA0FjJJV6FzvuDr98kFza0VgiPzUTefTDgF2YvOBO
ZdjuizXRTvYcMAcnLmGLGA461IC8En8Aqbm488/+DBH+5DKjdABCNBowAIb/v+Q2
RmJd69YQysuBh3nTWGpyX/OyQ0xA9vG87oXbX0CGjQFmBo5y9ZvCnNKI5s6KuRCU
rOwPM8oEcOlwnJv41bsLaoTFVcFRyehN+e7TdGFO/HweXg8yMLnkCJOTPyjsEZT9
slLbIkCU4+Kc7RbufMAceSPI39avbExXiVYLtx2Nj5oX+qoMVcR7bPJipIyw6xy8
yRcbF80zb1MPIgDQwGIYOkma13uPomnA7exlcjFgdzX0yMFVbzsVWBXl9BPuJpZP
plxhv7yCVXryP2RKnCR1Z1k4nx72lKmugqyxqH6QTfSDa6FnIZKu0cXrAljxBgXK
gmX+lkK7hgceASFJOS3ywR3SxUPWUYIQaHj0c4rUoapHjSIO5LCt3n7DXTWNOYDE
YW9dMzlkWtaaqTd6rNL4RiMx6zo079Vp0+jadKWcIhz1wOuiLa/8wfc9Y5C4UkUv
CyL4UJPEBEf21iXiOaIj3XQCqfB+IbAHGNlHciuaTL5rHxCbH6rlcyupU3BW+GRs
jBNch3LJZk6m7cn0wcm6EqC951esp3Ub1muRtNLpybbx7PWMijGLVlKJp6A538OU
5GVweZZrG+7VYQB4TRWstz7ukKrMV0uwf9dNLcJYAKJp5v96Vuj+nQz53hxNpC36
m9IGjxNfHL8pMb+vLKaeakTgzUwDWcMPa5DgyVFfSwwEMEf9Yqsyc9Cag1XIHCWY
ojhWfWA/CesBF7vzI1oKMx4Mn9odcswv/j4fjvWglv5PI5xORpZWxFgJ7ERwTYrv
XKVg4DWRcCOuZHN1up7+6UHrRZzMZpC1JWjMZPJDBPQo06gwsJNvnCGRroA2NmBy
WEWKFW9f1M2yTi+3uXdYbZu4KADCCLhSGBAEq9CTl/rkZTMR9SL8MFrFkWeQycUA
kgQHAYPgn8Ea+HyEP82KETfY5WEWif4XT+t+blelgjNV/Z5ODKfUjnh9hEx0PUgH
u0yLFgBpnSs041b2E7wc3KfoSe7NQTnzaaEFURT4Wof5U2RGuqsckuJ3o57faUYm
k5qnSwJfNrYbbaOvIzHsp0ywkgVAqIIjTDO4cNvZJj68cUBqLGDWoQzpPPaFyH7b
RNiRohLbYwt4S+ARVFdVOqX0fXRVYRdUQEgc89lMDxRwDv46YPlMNndaFBFhtbQS
kuYaheC8EQSqCwi57nj4gGQZDwug6x3Q1cYRxzjtn7IuuP9UYJrjFgK+x7gwVXY8
F3pZAhKVej8CndxsNrIZf2oj1bO3PubmYpXljVs48uE8WF9Xt0ue9GVzn5r/MV9s
9Qw2OMKsXq4W93TLMtkzl5P8UCLUX0E2bsyXfGa/geexgTPcsuUNsYQ2Ta0VCoG3
7Os7/5EKfjE5mS+2RIJI5e9vHZ5OJiXSzRb0a+VEbj9MOP+4KNPoCIcJPjSmW7oh
WPrf5VIFPkT7H3VwMEebj9T1u0O+5GQTqkp3HNW7IXcLvVRzmPrQ1iR/mO52B3ES
ZxayucGqYXf2743ABMPPnnenVBu6KV1mdWuHe+hVJCNt5AhLYpKJlEfSECbzsq+3
HatWy/vQ4TUia3Po4KQmIDaeEfUgzPtmF7bCMaHoqAaAFCM11LJVkPN+r4eb6+Lt
lnqYk2d91Z7ror6wOPJTNzrlWRZVv7i2wj4bQvEteOHoPEugoPLXHedZfuKV/c93
VJuxd7zdLL8k5SAuPj1SwbueC3/x/uhLvh+DArBY9Mx00ASfqXDUvoAM4AkE13Mb
+M9r+wCYSJ8O2ICTvhnqQuim553VkxSV74pOWMzy12P8UQUR/EHsuQp2PpJ11Szm
E6POiMz9aiN0UCewuRWIlqZqjwrLj2D8bpMaawfpYuWXpXlkIe+1knermPFA7ItZ
pYrZGGfMyXP2Fd5LwKNTzgqN1rLs3mtX+GboO08+a9UeAIVr/O03gkEj9EV2C+e7
eCbueG/KAPzLXExCpI3SNFL4FJDzn7tBf1PBJ1TM3JBhH1Y8c91qSRfeY5j2hwEJ
zngd87Vu5FiF2BBuyqRkYGDbMOuziwZCaFz+yMTyzacuiFDoIiomYVRGorZEtIcA
R/DqkEfcSDawxSJGrDQedsn7P0cpkUvtOv6cWj5+6aNgVOG3agcgI7BQmue+8hcH
EoGfKY84wbQgjb/xN78JU0u3VjMOhgGNYMtqZ/eOWvxiD+fHGRhvSNCckGFEKuHj
r1xHKNoqlqwARO5f2mr4sK/d+53NA03nDT4pU66bgL/GaYcxVUU+PVBSr62L+JRy
MQJh1d53kPlYXr4pkpwyW3dfxC8CTsbuUahgMNbGx2U1wlxQ0XkHDnYW+DPCK1OX
Sx05OOKl1DGIpU91sz59FxQZ4nfZ/wFx+yp9Ne+AHaGLE0TNArgQ+d30idi+Br7J
TxHcs7k+dljyBT3+eMj8oIktcQ73h4b4EmC4CKtSw5SJ00izvUVHydiay9N/Jh7b
929fEALI/+deuhIplKuD0nGTP8ytINcc9PT0Q5dzBAbEs5dzWNmZG4FA9BOhMN6W
ckRr0zGfBJiUsL1JLzMXmVq8kMaxUv9pcLhqeLiEygHM8NHVHhrlk7ee5d+stQBx
idstfNn/N9cG0TBndrac0Ial1LcUopsqWKmEfDlcDIAJzR8plmgzpQ5UShRJ2ALs
gX1Ij7ZWurxFqFegpcASHm/aiT0HJ3Q2BdE4vB0YHsgbVfyMlEHgPtFDpiM8A8HO
0yq2q5gF4m/cDgiNKHWfauB33Fx2DRKZmTOhnfyPR6TsQmxUUWHHBl9ineIs5wiH
WRj/HASi8e7KIUQqB0R3YzCc0AWfigfhHW8Y/ZEaIk+Y+UBx7axOisGiLKR7fC6L
HXrf03EtWqu2QNS/QmYEJMgEyiyiOIpGAeuqqBTerqYJIEeuFbDggNz76YtuP+ze
47csYPhTQGdmrwhRT2GjNCNXejbs7S5kAK4fJc/E/NWrQARycHmfJEVuCUMSXToj
/qqFLYVB6L2gahnvsc38Rgs8HPWMflYJJhaxAScSIA5O9fZg9DTJEaPN7LDBr4Zi
jeTU5Pd87DrwkRJ293qeE2zNaC2wwDwOcQ8gcE3tkhFtIua+8R8oxx0tvloq2t50
P+99fJzrdNhMNas26tDk6zmKzWr1y5B74Y6J9mtGdzU6BExABGgYsT05/f2G9nXj
2qzPGneh/azofbqQOrUrypE/ls6CAEAupvzD3xXTEEtGDJpi4uHSbnxGo6QsuzaW
mkpKG1bscrhNTKXezIJuTrgB7gQZyR/ZrBXZ8/4s+labgiCX1MwJUAt29Zaha237
zopaV7Ud8e0cNzpIDPocrdTpP3bCX3DTb0sJl3FoyZ4bNQZK92ccSCwXNUi9IOGF
Mkis8qxbOWVIq7FL8t3GPvb1jA2f1o4EWUqQoHWU2L3Fson0PTk5D3GFFyI+/O+T
9kKtHfR9r7zqKOf+lZJ2jIIWD1+NuhQnfduVflijbmCuASmrFr/H1pdFdLAZtTUr
tDjniwuHLiH6FSWkPH74zHk01OsJDOIOaGZzL5kTFcv6ojzrEuHEZ96NJ4V+QnKW
8EgSLzHRPzM5gkHDWcXttFMuQXHOJb/R9fREdd10mlHvyjf4CMrTqsir3NQANJGd
PsUtCp3dStmdOrYS8TWDacv3dgZl4ulQHoM46ijPyZBTFl6xo/EWVbx1FpbMe8I3
ZeQFYFYQAKhbp2CQFQUkiLWf2SQtVPNSc2goe5x4X2z0ocMgBxHVtMoOCg8yoleB
DjR8+Fn4xBSuRu5BFQmg7ZKAz4Z8m+RjVXc9A1q6fOeb97o3w1AaCg6oQN2UMrAA
I9CT4dbsbYSxEpjfr6ClHg==

`pragma protect end_protected
