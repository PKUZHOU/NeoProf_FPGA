// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
QeLRB9goLjAI7t5X5pbXAHBz0PYlSoBIdPgh4FTHuvT7AuQXyTU63sfzCO/J3Ahe
lHAucGiOtF6UpyrUOiFWPt17qKWdMLQWrqAWT5Kaprn7xzlrgO2fm4SwymPUUuQP
8pIAk+xKgm4UezhZuVdBnS8R0wgx0gdoZZXh3kTBteA=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 9536 )
`pragma protect data_block
tiNz5f6tQMzPTQPqu3VX8aKhzixEcJdOU63m4PIj8tpNErvZtgll0Dl4GrBuC+w5
bSCU1CWX6qNxkTM0bnXKwdomhdTb2Qse6x/V4QcoQk+hveYhCBtSnRDJ3W1wMX+r
iyEaeIQAzt06SEb8O1hfYCAHO8Wy6kGfTJfGabSbdLhxQ2g54fHIzx739Aop01RS
nctfexeNbBibRv3m2EvZ8flJXnFwdD6CmqGJS+kF9Pe8wAOEhnu2UmyiXL16kIH3
E14TysUBu9oE69072WH4yaHrRql7J3ZybTSL6TbbMy73BjJdoIklfWx4H+gaFYjo
D7xRBvyQgfUOahPtkH4DsUe+uu47bWQ3GuIO1vpe3o2Xk8Za1GMPfe1zn9IedtWr
gpKrXHbNAmB567NFD4mLAD1ygYFecNhl86mBT3cocZqcWVwlQk1Fixekgkc8YWrI
FnN6M13i2PiRywtgacP8ICSNXuUDcJ6BxCH1cWsQbF4PfxDGUyUUNXCEzXKv2xf0
iyugKKqFDZb/FoSCoj9vJxxBUrq9rHXSwLP63c2+V/Nt6/kPxmdkBHv4rQ5NEADp
VcNoNrNz+shbniT2bcT4h7SCKmxb717BBL4kfUq6UItQFanX7vLCq0eLreTEiJ+S
jjH5jk68lpadIykeVb8dOC1oPHKVhElaunMnj4eM7w73kMiBbOcD5XTmZRt59oFU
EHIPT1Fd1xDH46ui9UDs6ho57TZgpvrbfjmxy9opC/nO0Wu038l7UX5lbiOFFBQS
SzRn08MGqSThhGp3Hqf5qzIxGKi+pEO4KT9ukuJ7FZyp+inrHZD7z6gd/cjuw6nh
4H+mBJWlu2wqEd1/HISnxh/XO+vdKXgBMD1GzGasKEluSXdmhMi0XU6e890RyLLG
esixbEdG8Ns4ibWrBIRFC3P5IU56FZBc51IhJyt17KlkKwfn8SHvi1tDkS9H6+SJ
PUaLGAiaHsSv4l2VfAc5Tk28woX+lbe5nXi8PzjJ7dpqeVJVqI4WaRgn2jKXE00e
uHlxXrQ860GbZJwHjoW+AREhVHb+0S/gtWjUMFBZgVMMka8aMzxI1zPrB4+7SPdV
EMWhCHjmeGv8OMyErzwKdY2wJKxxELk7ooMOTVVba5SiAAjw632uCDiirUe4NMC1
F4b1EGs/TH5qnsB/Zw45FS5MRq08YnaqhzP4NFrhowu7DkjVYwofcT8PC6P3+Hc+
o7jqFdbIUz+iRQREW+MqxT1C9vG4zmwp0ewQpJhN/k6uilQMB7GpeH3ZI3Gn8NfE
DmMt5iE/ZXJGxoAQOyD2/AlYRkyrEsPmopD8CCvS1Nsg8hF2+rKNqRO6g3pWI8ka
YonA4kiNSNPCeu2kPi1G9169FUaMwXb2gDoxuao4E43XN4XEF1rgG70DgaZPFhrB
0Nf68xepHxA9mELUT4r3xTPqnZWyra8ogKlFn5cQ6fBhd9+KhBfAEaP5MGzoIONq
P6A91qxa7aquZ17nA72hHNGN8n2h9SEwkdtJnzGk+gl5W5NGQjQhUHl9f81N60iW
epdoyDM0qkoz5/fLoTIYPy/MJbFv1Dchyg8KqT/paRk4L49i2FfIOPQz9LLEBEaM
uSUJQoWDy5muy8LBaY58rHK00gmC29EkGbJTltSh370OMddMltiUojTdtGihlFao
XhetDp6Fk6V2FtC/J4DU6QZnUfwWazYKL4MokhoOXrNRnUfRec9c4LD5/GNd+7BP
sCjnm9/zVAaUhHSbw7l6QElrFjjzOP1WZMNv7jFJl67wZboOusVxK5Mh7Jptm7Mc
FNBAZ6Nrdm178Vb8T3JErrTh1G4EuqEq990EbJ7TDcEj/weYuaNXMdCtHQyXcvhb
abqxZCUS6JODgm9ywjirIdq0bQT2Y7Hyo263SSU5hMx+oToMeoU+uYDi6eQLROf1
DTmIsteFDxNZSSS8c6HqddBg09ffhOvngqj/IaIgsXXEj/lj/P/ghNWun/BoSwnz
f8HT86wp1oyX1ZVCrvHhfPsJCbf3HeoE920zFx6pFJ2iRVIVnh38yn8liWlU6o5t
Q/Lt3S5z+ODo+SIQTsGKsbUfZB05ECptohyyEBHE0qRX/t6bj6ds4j25CKjBG1vI
3ySTr1WnrB1okvpDJEbU8r7+lHDKDSXR8l1UoUmpD3eV6XEzEtdGA8elmFsh2YW/
BGA+77terU3bYUxGdDAnRh2okzVN7D9MR/3Qh4WOupnf73r58RLZhmEGcIQm2b3+
2L3a89IZueGKjxNxZzsJedO3Vbct95aarvqhpudQXS+YxkHMvO5PDsnPxTgKAwjR
u/HLkL3u/3ahNXyd1xuwwqqFUsf+JNL47kRhuTapRX+mElipp9iq7tT0SsjI+I1C
w6o+1Xi/j3FmgayoVnvl0sBWsE1UqRubtk3/jmSSVmd23TVJDWdY6EPUa4bL3Wdh
12gxQvkjFjN8VxAsbwrnojePbFWJzOlyEFWqtXFVYnBmdyXdH2rsPQJw27M2jQ4p
AObd3z4zHm4mVnKEqGzXT7g5/fW86qaQTZS7d4fdTSomA+lBSUnYjFT49bK8FMk0
AjgIenqIJ/fufPkQ5U+9/LvmNv+H+nHIIerDQV6VPk9iGfNYY6MynbNdJgYeb8+z
tLUwuOWxQhqHzFRTuVPGkV9GRklo44YinEY2fYc54reJmUf3l4Eg4KL4FxgMqfGt
jlidXwz5S51G5wlZvmOCPmsDfTysdrwDida87NT0L6Dx+84/grcBrW5KU5Dvqnmz
5y8XpGhHhb/8NLhbd6T+kYn3mvPFt521vSHJ7J3GG9f0SG/XPfWtXA2y7etvvPqh
0bjah5bUV6n1678FPCsRFmAWg1JXpUNRAtyLctvYz5HinIP7Ka1qdVOjQ3MO1Qzm
hWhfCyZecDTXkMT9GLJxOMHnP/oDg31DsrZbCUsC00oJzA5sO7JdLdHBkhCplNoh
aruiN7yU5lbeuXvteqDKaiERwykDrrgpNeIET6znkJ9o4ZVPlENf7AK8To3fiabQ
uaDl0L5h1JaCoPovAB/IR7MpaHSQ6mns3AXLLpxMW5yDdZtvBj/1yjnrDesGkfHo
TT4npcu4dpmnAirPCxTJdKOVwBMpTfLM4iy6niJ9snaTzHwgBQ4k48zOfL6MFxJ/
12i6//9fo9lGIFA2KO6uISo2KnzHf1d68YbBVhYQsrN/rJHxg108nkw9Lr09X9qd
L1Anhfp5JNGGJExamlSnZHh7cyWQ9GUWr3yqgdS3R1LcgHoQXFQJetqyMIUJpbhz
0lILnXtu+nfHMuCcmBAs5qIEU1exPUsXaTvM2/Q3Gu/wWW3iENH9Zyy3y9QKaNtt
xW69vTFslTVymD8gYFn3v80i+Mi4NgUmC6Sau+GZiu/fye2Y++e55cIGW35uJxJf
penj31gdUD6olo+ZaY1opk+uJbarb2663xGomuR4i0/yIBiD/dqGx8iAiVgAhmoo
TF6XQeumYbq/o4z7+WhJH8lbBmMCXPEHhM8aZLS+qs0Z63u9yTt0/g9F8JyeI6kQ
zG7/sk2iFmqTvs78EIq1bIT6AOyyK5fKNJWIQn8APYjCTihyIrJ7YOEQkI5dmpqS
puKX1m/AUwjTd4IvEZyP+omejmqkbQGQtoWvZMxV/peIQDa8TlcE8cbe/iCPJg3U
vu6r2Uy9gP6XN4HYDidjwMUncgwsOZma00twcVKyU41aLUsSDijTaXAUpA5O+KTq
GCTDkHLx+gqdG8Sz4JH14DqR08EfDj8H8GxZq9bPL6gYrzt3UojHGFXAcb3urFhc
VUxMrEDa/7hv1TCmV01UFd8l4hyMgDNdH7aprZt6viQADaCWrbn69WXl49C5PJp+
bhVlwMtbpkFZz2lyJ+1arUrfM0C8wSPK9nie4EOvAxZDfPVrzawzyJLO9pIDvpYP
JSHpWHRjxwdvBY5sbIPxWN99unVjug5TsQzcBDgenjgeYPIY//B8ShfhSE0bRNWh
JR2cNAtRuTjvdP6XQC446TRnXBOyQoKPFxoQTc5jlc2M7wg3A3VGw3B5L2t8XjNS
JX3zMijFC8K6nelcWJsQMoL07i5JL8+S9YOSFXwioTegEo9DmlO+uxYXwt4I6O8o
I3y23EZ72GK5W4rDivNHgyj9TrzhbvwFBci1IhZ2VM7zKn+Mg813CvzUUKlu/U58
QWv3AU5YQYKRAr73bKDlY2wLXH//e8Pl2/9m1TJ85IE/G119yK5pI/tN/x4GEahh
1nJlAG05R0WWQ+FG+lPej3Xq+67mmBITcFYQyPGwu/9Ho6XrFaw/vqh8r3VwyI9m
VSyY56DT2IHVwqEBCdh80MDlxdYngEd8/qLbtqI6QOOKhvllM+xxyEv3LNEAHiqP
zCVTgN97ePAFek5cIjnre304Q3PAr+v6CcN2TxPC+wJJdN0BIelcDzGO+rMCum2Z
5nESV5ad5OqkMTQPVWETWzvUtHzY01OnwyfJjVtFNQDKsZA0fcdz9UKD69CpHVvg
sbnXSr46JuhWw1hh7AEXWuxn5/kRlN5GOisD5TbH9ypcoSHSkKnu2cErH7QrHdQ8
rKJ6Q55Lan2WOBWCl1GujmrSXi8jAgq8ilJ6uqhec9kyOWpFwVICeUGzQ3bLSBwu
GZsVrH/Qj6KLW7rgsTQgC+zCEoQogjBjvHwk0OBTzDzX4N+baOtQpx36NkZvh7zR
tL/EEOJ9/ukwV7enIIBG2fvkCFI3Yuky6z9mYp2l3DLEO34myKH7iuuX2jyBiww3
RdF/sFwPKGvcZRkaGw9xOYuZ3Mx2whH31Wq8mSQCq4nH4zgIVRIaTjQ0wprqqVFG
kZIRhvTy4W5j5BwvgYXyw8b3xwtA+l+t5USmStAztiK55QC24lZ6W/PuB7cRDogx
oOHeWWsnDbbqod9ERpkkEB840qZ2nzeUuRbLaWcNrSoGg/LMxOOUYnyqtkkInAd9
PAjoUxCQ2sQiz28Kt29QY1fBI9/S8P/8OY+OIMDCgiMCuPqzgKRHwK53BPVwgeuB
BQ9FrUyQCZJkcGnG/UE/EO/kXuxIYT9YwbAypPyd0eQjIP0O+OosCTHtRzO0kJA5
wrxhMs9uDQbmgBah7XoTJFxchR5qh8aTjhSNvmDtTfamAdX0hUxnibuQPsNyPvjD
WSmyK/eog8Fg7GU2sSPzxYtNfgII1mqRJV1Yr8KnsAcZK6y6cPegHIAgw9pyxzCC
rqWBBwSsR6IsYdp8+E9xXudIp7EHYyPIcUF4aE7IBZfiF7jeouvFSYJpUgoqKu0n
BGGtbuIhANHVIN8cWsfyLA7B+gHNM5cDmQeLQ40wjhzKfpNtx9V+DZMzCNwzQo2j
TC0XNlfr03XPLltJzh+KLEVqtPpHh/3B3O7aa08Q/rkpV7h3fGGLa/kgoFygMb/n
C1rlmCtyplphYBjClXN8QtR6HWwKUSYNaK6FWko/Q0j7tadK5kdszwYagdCblrl5
HZoCQC+NFe2U8Xzp0xeX6yUOzIVwsXPrhrKoF6wTFZ9g6reH2v98OCUOJDDQ28Si
a5rhRiH6n+kMagqDqTQ3QfdXPIt09S6qUybOp//O2dvDbUlW738RXIcOO5dZe0Lo
tH+znqIwzhYhy3fSFD2uL7T850qxG+Q2u5oDfWo4qKJn9d9B8vAik8pPgPV5e+3D
hXlWxj6K2I0vSCdkwRHL39utsDCpBeg4DiD7FZ5sA5DjU0/TO/z/WxUkp8BEoymB
tC9G4wG4JJC/1HLd1P4jeyd/tkzC7bQ0PCcYw57Y0Lj5ykAIUiGoop7CgkoxR77p
SJiYJo5ljTlvA86jH5UAIRwkWQe5PdVztRJS5mV5T/f3+YcbpPClBQJzPw3x/NIJ
fqTG5V8M5mPFqKeY1i8KEkziSeYTvOBRX5nvo2EYawmMEHvxxxWwm2KXg4P/Ka4N
GqlUfjLfrLHeHRZzX/dPcbwB7Js+LspJAfWVWU+MFjXGSdgqHeAWsrAgJM3//6gF
HYHblx0hL3I3HUSC/CO+vuKBug+PT30+UPea3bPlCh53B+6mXs1yIH3GK6u1UDD/
x00jbNZXtkuco+Lz15hzpuNOOWakj4toYntCXSR0s1xwhY/a1LDxJqVYT3RJOWjZ
dGzk3WvYX7fmkkGP0dsaaqqhhC3YPTguE5ZIPuFE+r22A3e1ggcNWlSxY0zxDmfz
poH7v3yU2ry9QBMTuqeI1A652YnesYI7Aq4EE//oq0sdqGyysA4BOU9jcG1QA/7l
rqpf3popSgGkUvMLg7UN0GGL3Z//im3GdrA8FKSbzcW70nKc0PGL6/kuMRV5mevv
0XwsPIvFhMpKwAPHSE7zbZepDA3fOGhg83TBK4q7Jqs3FHIt6E7RKqMbptYjSZJw
AuuqhsdC01PRNGhfG+9Knm8BX+2e6PhN1cDGvkjTfxZNw3TBWPlMhuO1CaQeEyKB
LLP8kgPqDejPOfTW4YvD9izQ4jljSv9wXg9gWg3EngoGqzaBcM5ueNzJdFQl2UAn
N25JJUZ/DaMQlPL7KZUzOSlPRyquJNCWmg7OR0RZhc7H3P+nvNKuFWlx1N/qGS1w
7MZfBYzT+sauBhOX6t6Lr8Muii/Tf48YmSM93OwxPIz6RHeS7w2bS0Vo3tH6POVC
pyyUdFhTD1x1I2eCEDD1wAPd83f0jYpL1P2R0WE9NDTHOuEU6n+rsAxKhfcwyn0/
ETcSv0SgKM3bYT+sXfub/tMh6+BeZu6+CeCV7adAnzoBFMlIlWramxbamd6eSrOm
63dRZtdurqiyn6p9GrKIYJyJOmztrFkLfida8ck6hPxGUM9AzCErEtLO51aHiRc+
87+/XYcT2vG7VzjpFXv5v4pO7YBff8VuxvIT7Vq/Z5gf7pl3LF+1osmp+JhcBjYY
SSv3QNvrWOVsrT6mOPNT1kclfc7kcrDI+JJzTIsaHlrolK5JwPPw+deiW0+xbq+6
3zzsXtmxeTE8mhnS29W0xwceS675JIt1yxvMKPct7ClI/wVmiwR7a/AutANF85kN
se8y25RFd5XkrRjWAnLSdowPAv0U3HL+ZIGJCvz0q0it/o1dlqlntPu3YsmCj0E3
wExriMN4jIpAD7o3Q9rf6KEIRZw1/f4vfOkxO7X4HSe7iU6yRqi9zy+wLEUkeJWS
/y+0gg7U20Rq3gzBUxg5Dti3m6qdre3Hu0Flr32empfjn2I7WeKy5Bt6kOxx1sw+
XDHY1eC5niVu/gi55co0s3US9hmBWbPnvunUPJbYLo4k293TKCdGMRx14UjaAnf4
eexf3KxkebxuRUE7OiN3i4E51QoqAKVWDAsn2F3/6eDIJsrKCRXLuwcOyuht6D/E
G3W2S0io2gg3QYN+Gv8su4TB/rDZy7ESdohy4zeYTNAPUxhDTxoYxMXN/SqPQMOa
R8gRkH5edRAzxqpob/crlfWOJmY1phvBpgZPJUnsx5kpwCAOoxwjyvp+kj+yqKq+
LBk0bne1zRTYHVT7lN9ilytnEknFBXdlxHJuZuyzAEcR/Q+yED99TuNBCZf+Om6L
lePXa5L9J8ZipfRQkIeGrHy5cv6jGy/sCcJdPXI1yN/5ms764SkoSAESxTcq9fVV
w/oL8Hoer0M8fGVJ4K9MnE6yR2BlqfGjQHq64tPlYMB75Jl8vFEQkOkI/YG1Ygd5
pr36LI8xmQJRmegOMeoHa6ckkc1uu6hARDu3GJininpHTJUeyuDp6pxo9wXx7ayH
B0EnWtpQXXlswiHFmfiezXf6WGseUWyxQlHuUU79DlW0ky8thTUjjSE8Ms0RDpei
5nA0kVrThtGEobFKALNv7CrKexUq42961qP4mDrdtQ6POB/N9/rXt5VrY0OQRTbX
iQrYPriSLLd64GGrutTswxrKIm25Zi7pbYp9xiX06nbbXiKdwuNXwwUkWSjDjEBF
A9IO+u7lKrpkWVnF2wyHCi2aWO+NoEkngntyuRk8zeZm00INU+iTk7qKNSCJT4bu
8CyGW/EHRFzkxsKf82TLRDNi1KFP9PDyOg5lfF6ZxZoIk6EWy5hF8zdiQoRxGAMY
n0RBT/xs0z1Bj3d4mzENkRWOmHl//wpSXBXpLpJ8HRuFsv7ZwpfeBTqT4abGC5e1
4dn4SCBhXZknZ93W8w1aUajP9AJZdfASAOyb6KjypuMWkUekoi8oDJyQ3CIJJuTA
BwuOA/u1GMaO0Fj8iBH5dMX/WCEuqhEgHk0JTShDbbF6d7yYEqTNQAIrhbkm+IzM
JDeupnaDd0nI++cDyef2YWlFVIxitSjyR3Q4DZv3b8wGlzxqhG9+UGg22rYtqC3A
kS7U2wyPo5DdWWikSPMT5V1Udu9VIDZ47ZR7dhNTLA/E4O2b/OqofUjZXj1dnM8Z
vZXTTvF+f5iEarjei8TsdHsftpeXkoSZrr6lQ4KM2U4VruuVydIgGfEOjIOyhJD+
26lnW6q2UK2blPVIP+wug5B1xTDY9ovwGCMhoNLzse3tba6p1tPEZjejMcNT9ES3
R7ie7mKTVuojnfjKfE6p5jSPd9UB/C8jKrfPuf4a8HWtdEAsae66nyyjlHJ5wyZc
uQi5/47Ive0X+pISiFptpLYldyZGFTbK1x/ZSfKQS6bs1ZNQDkF6y3X+EKIVMdD6
LoAwozrVe49vhdBstXffraNz4Zg6uV6VYsYyTJ6pfrZZCCDnWNVMiEEjuLDn0QI7
jWf5BHvJCsS3Mn+n4xqoH30OSoG3Ny00EhWCllrnWXxDf3mLMhSaGJVIzyK9SdZY
8n1UKkZ60xLcVCeCGQuxtyepR+dgtnqBGOoWoMpHucYjMgSfe/krAf6SwfHx+6ai
Uc67fKpFtCjcRJVERnI+M4F0OZjakZDm/p2HAFrC0L8xqbufEIrKjNieANbp23vd
gzv2yveo4huy3wErnEkn1stIH1btJsmWTXS0idF+U1V9W0BhpkKUPy1pO0pMFiOZ
aSfyBBSoGSOjrGOPPKtfI/twcKGiB4yrJs8k9CB0dQ1QPTrIiD5ItXe/C2TuNYZY
1NnsNXHSqktPyq/d5a9ulQsQuYYNFA3Q+mCa5NEDS/TRJ4KKDFosWH6wjb8h2qVj
CoWN/qm4Iq+qelBSAcbGqVVkVWlf86rHeN3Fh5vKC1JAOIz1ce/7F0LOiejysLuS
utJmeKbW+2dLCFRCo4mZNMZJ8A6BzflOQx+e6AlmcHzqB5sQSN9GGOsVvaQjeqyV
cIbxjW2Op6X2qyrZ3XEE1/Yc35HE5eZ45VAgzRyG8h1ZP4zzqJfAPNBrVXDQfXu2
rjU25250ucX+RZLKESgmqKAi4m1HM4846Luaj5oMQWe4/qa1jbnhYFrK6Y097xEQ
ItRKpnzKtUsv2KZ9mB5UvXdKTk3yhsFQdrHubXcPlb/gr0PTthCPIeGHyhISyWrk
RynjwRMGYzCRMl74ax6uQtghI8UdxNetDkf8Pc6//z4JY9M/sruD/+xvzX/2Q1g3
E2+/MBZ2ZRRdQYNcGbQ24XkLHj7pPFA6sNNrfbihYTzJpCrmvjuQhFXdF+K4KaVc
G3BiBQ/mtqzDeTYP/oldOB1URoqiSEr/2GtMVuX4Li4Ev5S7+tBlX6+OHz2WQSh0
VmH2aqNPR+saUXVHOjdzDqGYNv5ZclSlBtQW1zd7/OcmkZH7JelQ7X+LNKkgT0FM
yLn8R+KnQLYuuDL1eadlsP7Q2VBQLxG2ewXgeebNPJgXGfdgCkFqgR1M8q89yar6
jmJ8CrOnyul9Pl7ntQMBybPTe6X1RgEEq8rNxIcDduQ7chy7dj8G/Q2G3T0sshAo
ZOJqAup5sPICNE/49KYj+NM3Dpb+xZcvKBO1aRZLh5F0IdJ+qr5qCgxWJI6yC78Y
efcRI8ZbsoYG5II56ZPaaHoYEo8CVq+6wksypdr58JaacauR34ej1T70NkQYOwtR
CpIeJEdGVrPNaIZ+S6BYY33rWa36+dFFfzRBHmWrMgY1r8oI2LZDtVsAylzMGzXs
rOgA6JRn7K6sVUVd2/nJVSK/U98RWH5c5OiUQtBlUrn0jIbXny/P49mtbhLeavy7
NG3NBu7+y12uKN0h96tByyU3N3imqHnGA9Xwnkr3yK9JLXYSKMPvMoXrXQYrKnXR
R9ApLlTo6imuwilo/DiL5AWTVBkqp9dg6wh3de7NJ2Q44xJ/VhdTTDbj6FQjFtVd
Thc5mLkdKLrpvcfwbEqbSx5AhZ5JTb1pIA0hXEuF0yHSgkgXHYcl045V6+5vOC7P
EHrGXmwhxRRExnO8hPp0lh4v1BkNA9oU9SzIEKHuu0sQy83zNYGJAvH4SNkx2pMk
LWParkAaiGdMlMSM3m5cWLUGwTIlkmQ70ViPO1to+Me/lyF04wVUkJGCwM21dwp7
cxmsf0JN7EggNgKTNyHCrxix+sjOO/ERTIzDYWhuv5PQ3irlICUHLFfrRP4+uMXx
L76C6LoUZWeUwiLI8/qPanBBr6XeD4n8Gd90tM1qI8iKnI2mDrzrhI6L9ub8smrX
Ksh6WfZUhLCeE8w9ud49H7OeXtIaCzy8yY1J7RDziNAhkJRnLrDMPiineQHJVCAB
BOg8BdifGW+YuY53Z5pFQqGIJILDidHyRKnBVG1YO5k5ngRGcaRZzRsUx6sNrS/9
5cpHQluKmYXvCdMgDv7b5Ps6wx8XFTnWCUcm1PPBKOevXf7AtpyoMf+2psVqRuqA
6Jw9XI0RQWEzmwwqj+svy3h3DZ+3lLGQ1kVMUnvKyNaDVN89VfxWT/IyYDnuUL0O
3uodvULPNGxjqlTTEXxFNqi95N1Cufl40DX7NMqA1BoNtDq3KUCfq2e6iElO44U+
Gf1Sqg0d5UY0hQsE20PGUuQ3w6ltuEpR6217uDzOtVAO/Ir5KwmdYs0VmA6pTzbi
Fn3yV/YeM/k/Nz2ikdyJbPqO/fdKM4Ds4QZHIPfOaxTjhhUWZPRmltKhtQduodQY
ZzZ10WswrIBlUeXNLYRqP5+e429SEoP7LthI8x3FqszxT+W4BQd8yKH6+a8NLNI5
a8D2kQjhRuuY3/fYtC2dukcBX/rdzVEHq6ngd4qP44tQ9ENEt6F2afKgG/+8MDvb
2xepOHL83RUgY6n8JvDLprwDTU8ovXuEgURU+FV6N2xzyuUW9cBSb2hI9rMpesZ3
vM7W/4A840tCmQQIpVRiib1zmQk1MWsQO8Dsie933C081dwz2QcFsz48/ZEXVvCb
wAh8gplu8W1hgTh3WzJGzkNqGBjUdZPVAp6Sk+280QsjbW2EBDx8P3PqT5fEPM49
zcdlaoib4mtRmhHhuj0BeWXRWcfk1s99LBDGvDEvrOXrm4EMfbVLbc9eLXQOrgqc
cQ0CXr5pszI+/exWYfpIRSCodOevzxsiEd1F3ucc5WiNrUbEYczLRzYy8byWdLAp
4P9lxbfhTPptcjdHdWLaV9Vn3QmFwO/kVfu8eLddXz/vMM7AWO9URvP25Xek7wIm
S63H9pjG/x4Cz9JmzxK3udmvpZjYKdSKvf93aojVIjMCqa6CBwjng9Wzvs9Hye+n
DvKoS7suZ2eRcfeT0pknskSXozxDPtMbhBvAKjr0z89+O6E0rxp89YZNTesffDyp
GjWlFHefs94099EFOGjRTPoXQ98GCwhYelrxdYaae0wtaJItmLSsus4Ug2qBYPSC
grwbUPMCMo/ZqoMTa/A6kyFW5u5/0Y24/upxlvsIcPHu8KT699Jgzu9hO2QdxJe6
rfE136Hv42Eqg4DKG2wmoXcRgPGiEL6HhrMwIE/EOL3l60tR4Kryb6h68Cd+sruh
FfNQY3bSQfLOcVReRhpCKeBBjeCe8rdtorz/ykmSay/dIwDq8HTGgHmBzz/BYCZ9
g3THy5zQJ0yLV1oCEX8gj1kLgHa/YFGjRkoe7zMd4mdNOG83n/dixvqymGstQSMS
1gY6P/szuH/jJzL1VIXbFEc5Wymb750cXwTz2ab2EhDBxmLSFOCBjyVmvaI9FTEz
tDTktRr5dyZrP9KQfZozpztnh46b1tbk8dd9NHwiBatcUd3kxtcMFVc316Mb2356
1OrA9hGzWrtISKVn4xf5QVIdbuWCiCH+xmg+G/pHQbmjNZgSgxqnFMmkB9MstNdU
dS4LiiEC44634O78Y5jqnloid56mdIplrcoNtPNNTtF7P4IbLAmnfVqHguHKjLLc
gRS4986Z3uSuzczn2ZHuOdB6QPjxhgd/bPQVXsv9Wau2B8qCK81sAW3WZxItMIMR
qcfQTbha66VMsHgDIBY7dQLl3LijvOUITZSPjw+p1HA5xrMm5DDQ0xHnjVHmG2nE
bpRkaYRgFDIrGgpZSLRLJMyZmF2Tr9TDFG1hCReyIRN52WkSQi1NWHCrCRJiA3Kl
VGcdNgs63vahjqpfSylUuH7aOKk0EM6s7Ozf7arBprmHzUW2/t0t0THdWbwPZCEM
JVi4ybZKcTUL5P9pNS3fccWkRUJsLiEMEIiIKLlOZyk3pS8K/UBs6tdaBfVRuahq
EWGdI/HofUNo549jx0OKM2UzWYdYQVuujjketfit3c+7ZWetOP0nbHCUL/AdDzmP
b73lKsWT1F91fQ800HiSyFYWk9adn7BH6xZ8h5PuAq7pc4DULNswP4UmVg1UghGD
iOef1DRT6jNCK5MYA073sD1lthSMlDmtu4UwMZtFuS7Awb2g9W+nrEsJLiI1gPKE
Z9GgX0fojJxz9qw5rXOyj9nKwrLofoRa7Z0OS03dmoq+RtmRIsp0dOkU4eFda8OO
cf+sYUA3FgiBQEbG3sL3XhZlK4PVmo3dp7uHMPJhlOI=

`pragma protect end_protected
