// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
o/z30+an1aVYGly6mfX+cWCPCnOMqKSzGvPWbFQnzpEmEtQ9Zg90EDr9YDpepiD2
N5vHl8tUmKtF0ODy3UuMFjaRIgqTMOJuUOB0Ors/331OF1GJaBHEq77ukZMQJZy/
he078mOw/tgUC6tg2zKfluxP6+mspSM5bsuu8BYgqXhLZtbQTCOkKA==
//pragma protect end_key_block
//pragma protect digest_block
BQ9SE3frkm7fCqI+vf8a/DsjXVc=
//pragma protect end_digest_block
//pragma protect data_block
ILcjhNKBJM6v7H6PZ3aHsWICMYfgJAqyBPzguWu3W8fGuEj/5QBONv0WGrHyE2qa
JCeE8ljGRny9UO/EYxri1eQvTOIcABfgtKtlM00hCGsVL+ahrboL+wWkfj7vbplc
HBIkLu7NDYATTCYUx7Fzo8coQOxGJV4SWl50IZmSGVWidqj7G7oZbGI2S7hHfnUT
0ma0eHva6iJPNT3ELEdTzy39E2/8gzxp0nmWMn10IgLA/wDwMTLxMOSqrsvpELow
UzSTNG6/Tggwbb+nW4C5FoG8FIR/SySvgRsKGaLMColBuSahJTl+gB7ppOCMGXU0
H/yiPgoMcFZWA+hi/Y16c35sNyu3NJZ/1upIbtiM6BsunQTAtvVVoIRf2Q72anV+
4szOrOko4/sYj4KnxliT3Fjy0oLDZvemecrB94/3oIpRkR37US/m5uK39K5xtJg+
FLry5PfPnVdWdaZ2B7Ef0JIPZ2VD0sd+7SCDYamYqiE6DRnyEmjA2Dgna+mRdzWd
Ccz+a0ligVtRRjrZiifTLiclkAw9yHDtwk577Fxq4ZdfaIr+KuIJSpS4ERKxf3gH
j3mLiu4lfVN8dgw7U7FFyuAN51qDGidCeHfoso+9kgXsrXr4GfFW6tExh3zoIZcT
XaksbstRJZOpg654ecXIuB/TD/9AWrL3v9BepUSwI7gbg+toQ56OIrm4Ph45+Y8A
IXGpS5LV9Q9on/k80FscfQTIQx4fgovkk2nPbKi7Oymc9roTOrwiv3bqR1fr6Zpc
rhz0DtELiqAlyn5SCpJuLoD//pGa/ttxYU9r5K+xIA/GvAcx59sh05/cnpW7XT6u
Fh1iTT4cEV+jy7jzZo3EJZ5RI7nyESoJYM6m6e6gq6JolFkJjaGEu1uMozWpdHRB
+2MMs9M68yh1gy3r9vhUkDGQuwvTZROjeFGn4IHXXQUTLxBkxvmGcRjHXDQGYjmc
aQR535lV+nKPYdmrrfDckrwX0NYSZjH2vEIRIjxThH+BGpqjTybex5bHOTUIhB9t
XEa81/AJbEnA8bn+i+5xymUGIA7XJW76F5qk3nwwUWGFHOl1qSm0WHtAZ18QjY6I
zfvr1WNQ3whHCAfKvuJMdmNpJylUR5XOIac1Lavz3JAyKxqCdqUMdxJaGFEHb2aN
osZpZwF2e6drAE0tQGs8mq9bG6nhUlf1PXlwW3Jy4CeMFY6Ub6qowdS3CMB07DP2
lDdsvkh4BLrhpX5/84+137sN/UhuS7dOhudjw4myixjr18lOBLEZnHsfKTAYtvSu
dqhMjAFW43GmPOaacrtqFLkuU2ubwtneYxEt4zvcIDVvma5QjUR6uo9mM1IcHHv8
abWR13KOZ7oMKCQFaS8ZKW4tKA9KVcsU0YVVraKOIybbZGUNpLC1PMC91iWg6NgC
vRS4mm5NhH0UvodnOxGhD2Ww7+I7JbKhHR+fdo4iNTe4xoGvsUV9DjZe9qgSWId3
LJWfS60EhwwHuF8PHHvjcp0kelkjZ/KYyZBk/G5SW1nKSVJTrMPiWVWPVm4kCR6v
aVOB/dexa7g79EvFT4Yi6K2lsnCYadlRCW/o5OPRZKWAc3ldRANnf0mPjwBjrmaX
qJnhmLnb0VDCdFnz0E7b1xSlO64pdGoRVAhLsc8QCwpui+KY6rl/+DnoAaWhiUaR
mNtZdCs1MHfMgPhVGkwigd6R0Gd8JxPDgkKIJO2DF8C7+/BEzOFpFDqB9dnyBZ9m
VDq1HeA744d96/BsD9KBUZsi3EJ+KA/XtHd19iTyXmFwrmXt47dONh9DX7Ywu7z3
ZyB9988Qjwymndl7tSEE2PhEOq40kJBTzh7ZT5qTHmCdwTQhUjS4uAiYh/+X4hyv
Vk/Hb4NZ5dcfVDKdAK/SqGX9ab9cCPK3wMcwz5HzxG82T0dVJOJ1Xg1Q49ngEaNa
XO2FMBNqrI5SYqwx2VoWTGKAsSCN+1CXARAzBoOuy+fD2HrxxICt/xvx1RBOj9wE
7+NHi+R/flTbcksD+rEEok4rB7GWmmsezXXn8ezWnljP/9qp7EMPw0+IkyDXxHeM
8bMmaeiO1b1EW5YkS/0IK8/FdtGVvezbqy7NdUcszDhP2/cRaLxOz4PnRAMXXZR6
QhotyaGOTW7YlsJl4YQ5B5tSFwxqfAkQJtvf4K5WGMi5SbkASPrJ6ply57ht0UDm
g6Dyt3QGZuTN2O2GaJ6N8srl34NEVYW+9XFIDSQqJF5IvVdPSjcWMwZ0ruETHk2A
Kc8w+W9IXXkxCRHBqLXANwUBAYzv5pCGADCnSDxUnmNOuh/xmz9kCrAz3hIAqEvU
v+uNJyPt24/sRytiwONLJBF7MxuRCg2ENCloRASgV9+52g9JLPUUAW2ROKZtdTtT
kXZ/Vyz7Xz6evQlBexJlQ6O8ofZi0VgWF51fHt0ZZ4b+nSWPRCuhcFURDq15ep07
lkeZeIJC+YxwBukh4jv9YDjJ93TZZXMCr+FxSiZ5yM1pbpn0li6ijsa3ZsOv5Rqq
HeTU5MgsuDnVr03efQhRxSpFWCIn7O4JvpgCH+BH43T1V9hwIw5EfhKPjqrbe9Wg
cDangPxiuxsBmiNpVLoKzULdvejYVV9rKbXpEU6ETBiuambND6U0209SKuvCubR1
tRJOcJrbyInh6eEsxUhX2exJqUVu+bJFwq4937xozIGuR2ozF+1a9x5KX9ENb5Bl
6+cKqXTtdn2dKVRo2V0Cfkl/g19689vCxV13KfDQGodhzeajdTWCgNSruUhC3Wxz
XAF5Tj2wavWwSB8uutoRjqxSVLyqPAIVZzsWIYpAkXkelj8kaLxtNRP+CJG/uQl3
ARFTiSf/sBa4Rsyl/kk8EvIoxe3alMVqf5JC2k201EvG8k1mKMATircKNmpCvGPp
tucWj6TQmPLpzGB2Ww2PAB/HAEY5O0v1TMcOlhxqXbavxzTbmrhDCJZHUVlwlmMZ
fXm8qZXvGomiXkANgG9e7mbkcVD/svwfQm6Nv4BvVfTqqMRm2Oqhy+2M9uGLWluN
BnmutnFX6VMqDub3Uyt3bJXTQ6Q71YZNDO+3t1nKWEg1j09yYtK/T1ds1FOg4Bw3
tJX52LRucs3Oq1QzQIjX1gBB0cos1xAsNHh7K//HEvu7WUdnCTmGCUSdBBuuXjg3
ld1lx7zEv2hVpw++hnLxgk1ZAEkCUAWBXBS2TuPJX+FvFPwD+DRNkgomjtrLpuTX
PG93O0msnY6ThKCaVyiGCvs3AJXvoJZpjYai7WFd+AGnIuFsU63ZsXm9KVcffvNg
5aT/rNlwfrxZ33CbDBYw5o4pPRKeahMowdnurHq8fokWSbb4+SrSyo8Uhf1kaTkT
1BZTSkXl4ecMoCw50O+405HzjvEf4dzKBYOVL3CgyADvSShUqcegS4Hv4bqAmZjD
MsqxcYUgW4GNjjBKdorZkGueaqB31ITk2/OxUVzZjnFUEEJpMqCtEXcmkrocczQp
vXxg+hGKCPscp9nqwtA2IBr58XgUrautmNLepLCLo77Dmw0X41Ond0wcFCFpyuD1
X5v/Nm/OERrSUyVn5GypZ/Pdq84qG8FnNf0H1rzNGbRWPiH+hY1MfdOKhDliopXY
XcGEcw0PBc3429Qq8eatqQL833vNsyA8+9T0UbQXvv5bocLhLlUmZeXrNsVDExFY
maGDI/tShTbhNM7Oa8yw47fJSlHzT7N+bTB3arUaAYsJtnuJed503QFEE7dJucgo
a9ktwLhX3FuKEtqdbnMUEBhRO8SnI0Nha+9YxBX9qLjspEWS2YkmY5PygrPyvnv+
JWHmifEeiFJAAZTPAVgJKQXhmoQO8Zqm3PUcp85G2H4EiC5Cc/H9dTiWQ35tskkH
Ovp2kxNNBhaQ13IisyDRHgr14M3qXG8RpiVKN4S9U7U0rGnC0ubPX/Ti0nb18IX3
PTsgv/JSwnPZy8QVGr9Kcuozszf++mtVOYT3XmNqfdv5kWAh/Cc3PJR7C8oqueEF
Ya1SAT1NNMF2mOb0NEP70cHrJ09ahQ3UJ9E7NuUbtGGzezfQMGKaHLHLisS/np9o
lpypY8fPoc3b18fQeGR5DfqSgx9qcCfVnzDq6hhLfhnezDUMypytMpdHp0S2gUSP
Z+Uq4LQY09JVxKDfu17UAJw5uNM5fYWZSku/vI5UWveH9URWMdu97BHVFFsUPFRN
yRrGDaWMn2vIk+IUS93qmBXHAwBqg938Gih+p2DshpN/79lFnHOZk+lUOQX3WL+Q
wke8+6XR3G3xmbk97COYakGK57ZprLvU2H+O13TzYfvEA4tBYQ3GwPLuKJsEOGjV
NdDwL6e6y7038jv9WjQhJvu5inWjxzr1fdSiZ2yZ8Ph/d1QgCyWlDWO+lTuorSsH
EyJ21RUw4zGIq06yCQvUFYrRhf/PNwtn0DSEKyHDtJsh+3oDWy448x23igb/Pkjl
S85ejdBJpdatOyDVxUK21tTncY/WYi/5AkJqzFpFnaGiWGuUHxIU+M7CeSCTsFvU
jRZHKh4QFE9QmIor3lDPQRgZzTSAqJ/F77smbACGkhAtktTfqJssvtl1DwD6cvEB
l3s+bO7FCG1tiR4zffhG+9/BsJvM4ijYAxhXBrqHRWIZv4ZtqLVxI96yDlb1kt7k
g8tqW//OM2/Z4/Eqx54Gyxco+IqWiEC9gulm4CathjRlM1CgYUIs1VtB045+t6jC
qu8+75OcP47KJjxV0hoa8Mk4Y8tet8OKQQgzfbBMhRMV2SJ/qy31WVC2PmFRqZIE
4MPAmYrNOyCmsB49K4XO5nAc3cmxefIHMwFB23CKWvOUNjRC1uAi8K0LHJnKJFA2
oEmcjgDgEzris9FCRUi7/2F77qoOT8ME2e4215gEljX/HCdT3mNfPjGdSzUsWNPw
plfpL6ojzozNM0f+P/jIuZ5IYJeuqJ0Mz9zvnNyhOr9bZbGpMIPL/JNn5AQIxM88
DCPgOpbbFQtKfgMwsTe3paOYQv5wYnC4xrOCQE0ReGy90U1xcDPs0S5vkJlD4+Eo
hA389TIvdQVI26wEKDAQl+gU1hP6qCKDWs69TIEvElk0FmQyxW5j/Kc0acvOgDRh
amCVqyVxO8dd/Fu8+UE/lj0rRcecwEscc+uPhkUePn0wVoZ7dUBroPt/eeuTfytY
G2eAhaEVIJ33I1XZ2Et0sHRIbh6H+QffM/ySw4+ltAdzKHQ5sEo35NucEsZN+r69
/o/PK77oZUlAg+xjBD6M1ohNj+VEAD/EeXcxX/TDlVh/32jRxgpKoxuzGl2W4oUk
vbd5VEObqjmOnCqtHU9Bn7We2vPh/R6WFCO3N2sdzFfB/RfN/sRdPd/P/nvYwFGM
0+6M0tJLkbbP4HyTAPP8OXetQXKJ6CbOnd0YeE8pQB7bSTHH7hXCgQUlkArs4iR5
GvFsJnI+dp6oPLqhlOvTYZNIq/39JWMt0yTcN9Lj6+TsbiRdlGBbskxSzOt34oU2
4m8a+Rg0ZfPs8bB1M0UbNOqD1qNi6Iul5qD5q3/7x7MhnquVX7dT8jdgUmTTZ7A6
JAleAXg/7zQuch8OIgOAPLThbAMys2jImWpYkNH6WfGziE+4FxVna1aZtFWL2dlx
YDS91PGOT1hjBQPi1G9MilfMs0Jo6+JG+9B2F+hlr/2MAWjPcHIgNjaNSc7vKG6V
6ooI1yANHPcf9VZDFHGixl5i0R9CR7gWVbEs/0yjHquHZJbHg4KgxrYO5ZQQjK+2
Ti2nofgVTRaHajuM5hCP+2lLq2ulzWwYTrtWQgpNWeb2oQgXSoZWh2IkoYdIm4yF
dFgisdNFYggvKA/qaAUq0eLrpg0AZJDnWOwhKgpTEVpNLmwqEvVSYhKqkitFE7gy
T+6/u79e8FBIizeX7GI2J/NUd7ndserUYD9eFyo8vMOKk4WtJ35JUdB4zXPgrAIN
xzQGQh54FfKu/sJm6EpCpCATrxTWasDqdiUgFZHjTO0Ek1nfYSdQBLCGeO1KHbQz
W7zScQrsLFDQz8JdDTxbeU0pmr/C7QTyeWzgwPRHC6B7po3wRUb3ya9cikDE9GEJ
Bx7eDPSS3L/EKkq8acmtvbQBk+yd7a4+OwJsj4mGuSPdqSvrM3ZQJ0Yo4jpEgJ6r
8Tlu/Fxcqby7pb7mlVBaEjsqmT5NNMTRi4H1JQ3e65P5obiVJxbhdZmisUYw3cEx
tChLiMvM+7tftopDbjz6Q6lFImp6mW9qTycq2Xyq4dtO3+W2eXigHrrBEJknMjYV
i3ykxIyTKxi1YsLL9qMBZGFIaPgcdL4kBe/Xt6HW2SP803J4uJoYWBy5KxvX275F
dzBLFTe+6XoeeGXwWtE+bDXf9x73moMhUMW1SZvJnogKi8gnYIb6CnvT0uqwjltg
X8sPkH2pfGp4jZUy699U8ImF4/Lz4vomQassEq7tfEAo5LqTc8ptxjWw//+MyJJx
qGnpYS8lCHOoYoJhn1fbcmwR04N7kY9jefIqgJHlEDugHN6rTNOgiJFUPF9+Xx66
yKjlxdSn0oUHukFSr1YsZDJ5YRWVIslPd7NxeuUwR1l3+HYg/LqYi9VGmHEkpVNS
RcVn42PIQqctrTn+PbKUn4DXze/LtPnUfD6EBb0HLNuH+hW7ezUZVh3hMd/TiCDb
YIiXzpRPaiOieWvHI7R+G82tffVemm8n9AlMZ0S3pvEfbeq3mjI0gb8jhzHocPi9
noYvgaJIbpyBLCPsoVROhWxuzJoBozyspt9RRx8MwH/mEY6Rj+jfUyBTDubWfP3N
fDvH8WhNglVRSM9xdKIJrpS29aMVS/Tgjynw1+ERG/Q/O2KZ+i3LVSe4Q2IOKZNP
SvrjCn4lo0gr3jlE8xsshmarIYkUFI0djCytMmFIms8rR2tVfn9wGSldJ8fOBnhQ
iDIPWa+rx6Q5a1WM1jjxIRiVwlX1KYtWbxQ8ACPbimiQPVvXuZQf58Z5uM2y7wPF
o2VUZTCeUflHEOJNeDUScG46//2Tc4ea0fliRgUR8vG3JhXBqCBSiHCQ74Km08y+
EaLqQtwtjYEcv5p2HmazzjQLr5Dx//0BcQLO0HDpfH3z0uapg1O7tIidn+43gTJl
3YwK7YNuMUDJcBn8j7X1NTbM9QcVpCWDaz9VdAvZuc88rZLD8Rb41gsDWObQuTlY
VtNiIU+UTZdxWXSxRt7Mo/dxCYW0pJ9dLHKQrRi3a9vxe4NJ/4h6y9dlgy54lLbN
HDtwVjnJMD4ysu3AOP71bOa0bkJCRv4zxRDXjJAyycIRed2Ftobq3VXfbD3//ozI
J7h63mgWP8YdsbkBJ5q2XHI65KsqahvXUquicu0basD73R8vwuhpA2yb7D173/4+
ZjaFfff2MTvNlPYzP8Z9n2zMZwEMRYfuOjlpzRilvhfFpzJrdNZOBmoFSjieDGyz
PHKp+WZEX2aM6X/pDzzo35+mRwA/6OW7NzfoeGMnvvmDXeJub1+nCVl3q+WmrzRa
gP6f66tTQ3OYNjezOdAG8PBa8Q20i0s2azu/e8A+lPsZ4cRdfx/bELyYDOfFrgrU
QQXv+uJYsINdFG2cTFA2fPfGVoczXR3fQnS3o2IaevtSy5073HTXWgQQbgpbhuCA
wL1vz0lIIzHO87S7s1UnSRGD8i3cU13zu8kNGg5/ES+vKPDklIul7Wgp1u70CEz+
3+tHxRUDF0dkh5WKuxtxqaynRSD0VipoT/gN/zpivMHu3vvLQnyZIlVb4TvvRHf6
8eHTDg/wGtfZ8WzIC8JV16WTJ3AApMij9jyoOpD/RgVXWWhQ2yiMfsj158zUUxOW
gAFeY8pqWwVVvp3HMiNsz4Rhd5HQhPpI59CWGYzsMrz1qKXwAKy+mjydM0Rpkrzk
Iz4SXgWmEsU+W+PwGzqcx9UEqlt2skTe5sYwQoVqQOZDsUuf7mJzQ7NM54KQQKjY
D4Pn/7KqSYKqLPPv9DYrZTA8g40fAqSYF5xtrPU90Um5ygx3+0T4V2Cqsvqq5AlX
nGvO4DOxyEQXtwJq2IatjcWQxdLh4AVi1tVQJmtRK9zrMAZwL8tD33Ts8kgWuIsT
2Que/Au6mgxDJieYJC+a14AXakecukkfApub4wwy/zQ2CVLAbgyKqwMLA3n8R6Ex
JWQD5eAQV3nODtmDC4PFQU3iBQud/HMhf02VUGjwaizsjehG5qP8OFIdG+EWeECl
NPCzPfaNQMJTFU9+ADv+J6fjvcasSoGSM/fpCt81ECVBGshvGWgztAJbXnH8Z4Nx
5WKemyepizFugUtk2PEN1Z8bN4uuiTUXzPdmVtU1E9PomndWpsnbmqKyBBvOPlnZ
dvHwzPN5IDsx1WPiIbHTCY7WTc9uuosc4CRkSUuZLg+u1PRX19mpYZ8C/8TueL72
/JdcWjn+vcPvG452yViKeui0OYaHZPMyI0I3Gtd16dUDjkJ277zec2qDL2UvVFsW
/cOMBN4/a9l5LzRvIUwrziosCgAuL6A/Dq2Y4rQDTouXU7eHENvYZQCODjxyZ5uS
AV0YZIWgVB98hTP+YyP2DbXqi9hdZ7CqmtmUejcQ0mHS4gYWGdo3f19ACZ8Cu3/M
ECG5ogK+8QgTrj9Duj/axx+XDyESI6dF1K7/tZVdPercXmmuqw7wtX4YE/itxIo8
PiJGvBzCovaUbdGWGiZEjIoTMGcYRQiYDDtNn1Ernw+9gWY5aD1ZbupecZLFQxVA
dIuzkLZJNLaTM93cYOOaagAGqaAfU+HxNiwJrNBnjKHdNFk6K+qVe8OI43qIi66c
oFcxoIq1cH/6yoXoT8FLSuPLjFuCmbFatYXoKhJjL5SEwr4KdNuR3NVuYyP4KR3/
Igjm/KF6Q90E1ToQPDPW4kjS0AbTwqaIKDANi0PT9lPDz9peotKwJ2T/DgXC2KMo
HVhk2A2YMxbNyiHTxW1qHVypnXOe/NGC7zu9K64ExOFn3ufx4mE35U8Kom72NaqK
C9kbNGOlzWCJKEnkmyy0yU/n/h9paWADx9cTgpIu7o8Dj+UFnz341yERfuBWoq9Z
jSqYBkSgWhVsw/5fE8GtL7eWczIUt69AIyj5yXSAAoVaKVuYq2rW0H5tpXyJ+bLd
vj7VbJQe+w1jqt6z44hJQLfbhnC0aJKSN4IYQDBqBefTrvquFL2G5Jqm5F7q3hs9
uOy/YYzSdsH8zgYuFhLCckQt5+jjeweFr9Weuns7uYvTbCsxeqvpkP+iAgmyKsmp
L4xG2Udvtfi2wSl0Z74jFgLeuzWL07XlOsZwHbDtMrhaYMxgogDkL2OPt3gLf9E/
G5QuhdxVNMEEtUxmWSrvdnl6UzWiiht5EKiAARyFHDZguPKAAdF+pWUYtm3pNpci
8KqKChcWOJKx1IksIyvqm5WI0o2a3oY+O5eCPJ+uCbukNBiM/DqcrEZZUtjTvmh8
f58b0Plz8ugBWz5/i16XPW7suF4LV7LeqAarmYfXRhaqVAj+/CSC2xhnKmYUpy40
yOYma4uOEA6tLhRW5eu3hqqblL6Oexxg852vT21JIRs0RM/rrLe9KAhzvbhMJx1q
ZnsPs/+LM3qOz9Efof+h5b9dtyHWKTzWarWe7gylhHIXwJBBdpnQW/mU360BvSG6
MFl+xP0b7+KsU7zRSYzhuYKujukuqTvci9plJks1BowvM5xERVOKPMq2rsIWFjTN
2D+CsIOLmeIY1n70gakr1+ZaXuNs+dk3tGNxrDuSMSId0+6vWJliP72Uf7+41Mym
g+tbyBnDcF7EuAZVJrUN+hgkp5ktQoEspm17ON/OTtQHo+e84zowaODNAAmgOoUi
6TQpyY7MIA0Y1af3l8nGvC7lVgifItqgNYtmHvbdLrV+ffM78m9IzXqX+zTJ/jHI
dc/3y46t4gL92Xi8blzgSeVY4+iv2niN+avuVV9hcgRE56ebmKR7h1TpTuhRGZ3A
WJhAuWbqARFqwd6W2WUoKy++Sq4Qlwrh+FDZevsnylIB67XahKJ+w8GybqG5j67I
yzxlHlMvxZ1Iqj9De8TLKjSZHXsDr9dAY2KKxD7jQawvzlDyD7nvF4mfJPLa6u6n
CdeEpUj6uhUsaCXTvRD5VS7q0kT3zNIJfkWoG7ejtPd5T0VThwUzUZgQfHRBzEN7
/ivIrexaPXb3VDMkJ9gAV1hbes7GHsaOWXhCJXx5Yrg11TEP87XAxnz62rg2JZ2B
rAFzXEDA5nO1A2JDF0LTTJ4EndBzBquphirpbbYyzgf57LwIF+UmPvYhgHSSUSJA
+vx2QJogOwDUY1WuNYurbB/ujoNY6u/DtS4Q3wNoKu82mlO72jNJ+MXxWyrY9ggV
xXUBE3xtBHITCG/NAZfuCpgWJNg3IReE4z3YdSU1Bxvl4jhNTgblSazerZ2shV4A
m5TObweAKYi2k8HevrB1NakME9EUhcAcog43nStBkSkYeTye9zPkTR6F6OTeSOWb
XgbN5BVBHPsoM5WsbSxKAzP8vOXG5OAokYhJG1nzCLr2AJL1aEiKthhbBs/2/yQw
LvDfTOTAXJGyPSMRC6oBkOTYMlvkmMgECywONEX+ngR6onrU830tNFhG7hoewlJq
RhqAh3z6f5tlUOFlcS+r1Uuxwe9kSnAatUQKjzqxEIzbng8xonfNOJa9sfGndA/L
a+3QF92JiR5SxU60AuQpbEQwModDK72B6qmPYM3xq9ks7p6fgxIFG/Eyk6zff6fV
K8boSxyjnr4/Qn1fRDXch7CSvpUaiA0XofN962UH4qNRgMNMsQZF4+9/aa5ZyYkZ
jc7o0F96QrKTni8fvQPG2d9w2Vs0dqCEacgE8uGaItBcBJMN3QP2ZCpyUAbh8MZA
/0a68zO57Y03STY/LH3SHYt5yStegjH66/ZhmT6zeIiLM3/k9BevqoMcNFE79cOK
UzyVx5fFxWty4EddY7UbdyqUS6u0w9TgQ/sPxI1owRl1KSQOSKzmRsNUG7qVZFHc
iapDCnOhEzVyx7N4B9YDsHeoof5TeSgfw6YdQi0r+76tLlVHM0Ewb+y7A+6AGgks
zwfaKIA5W0ynL9g4tCV7vICjgsyZ8cX5OslTwWAMVLDhARFfS4q2CeFKH3qXOrmB
8HIA74Hy/4cN2NZTU/TWcBfkeryD7EoxPcvv6mroLVHqwPtBsjOSomZF/1hVgTY5
6aRruHmBRfJyxNCmXo3QGROVz2svKSrKfC6UvjuS1fweubiZnf0N9aodIQ4mf9gz
edv/i7mDtr6K56N5ghgghH2QeKOGAzRPLySLnZsrxzLGc2embSF74oeGO/kzHfuA
UnpQlhcC7lTiSqk4rwIxOu94J/SToXyYfBXgsOAW30qY5myezZPs4blH8hcPbDEU
qnerF4u+xVaE7WJi+mMgkJBThN9CgDl780XKeI/71wGJOwFao+fOmhrigXsuZMik
8oXkQ/1LOj/AyTlD80KhTndKFdWVipaxwbYMwxN3EH6taj4VZJuiAlYOVqwWKe3l
fVreMikMGC2nLCGvQd7z+nqmQvURZJ/n2/bwSvnPTquLDe5BvIx1aJDcqussHX1g
84RQcuolFT1FzqNmaerzPON92/ygNI7F9hl+PyEl14TzhE6JP0F/y4BbtOQOfbt/
UAIbU3V3tGGTQ1uF3/6WwmvCM4KlQrYjxCea6RPBiGLTFTsq2wUtw5yeyWOG0HLT
3hsuxX3rcv7TktUcdZiH3jRqJSp7miZcgiGFkSCvr3JWttCUMRYiMBhmMH0LwNp+
VcKZ+S2PiD859c9HwXlMUZHfEtzHeni5aHX47xfCd8yxBlunx6Vvho1KLw1wkZ2I
jp7Xja3cEH30YrCVTDo94LQbz59CD3iUassGpIv4k5CtS66oLJ5Do7vAgZzFIfCq
r51eiZ521aU/q8KRo319+XKacRFzDzKeLy7U2dIuaG7Y8r0ed2D7qm7upk0ofTBT
Yu+oZn3yxC9iVS1EHOXAGxJz1Kd4rIxzK+W2v8pKI6ZIfiq7o2aqZBomhtP/gUki
NDiWpWbth1FwymXukxvh7yrZ97K/WM0sOtP4kOySgyaAFTBIBDcxELrtUtN3axIo
7nfyyaihb59/ItWjS+NUKWmTH6xD1/L0ggoHfhqx0c/2Km2yN6DtJYPT4dcjUqAK
ank8RQbgjebIHgUti7lQBWoycid9um/JUsaDKl0bDcvbD3oZD0+/8HbUvUgpRSTB
1QTmanZQxt7gPbWilDUAATlq1m+IN9GzmYWkgrCYLRP+aP5//z6DitH6We9rw+6H
LvzDxMoRMB4epOx9mEwoqbRHkS8S2EvH6Hk5Un1bZRbJ/g3mZLHPWo55U8uxSRM0
q6nMeNzYJ11njWZPeMeh/DevZmZMI0G8HceqJh/paDSDn9CrhYxjaFO1d8Rh+x/2
bT4BX+L+ytbvq4OlXNCulElbSso7JLcQznBU3OMV/skMt8tBCCsxhToJgl0GqNVH
s5rzvIFuKfUqqM+ZnMKkVUgqRS5fofiQ4KIWaaW9lAqwH+voCjO8BhgZW4uUrLVK
+jnKf/vmyNv2fwGNn449rdF+QNeuYPAynZKY3eDbvwqJLk6FFboAEMXf7Aq18XAE
pNOOEXI6ZiD1FLCyFNmP6c/TOB5x164ACNRBaCCuXJRRnxgSrfoW8oX55+xfHqKM
iAChT0quC35UDBmhyzSWjbB3qyElJEoj2+Wp2QwySHRXieIOCU6xao1wrGNFvabk
B3vYcE5jLH5rWS6yn8nT1BjuGXvFqp9xaGN3avAjkaiF+eqNOAD1t+uNtdtqSrXW
WXu3XYl9MDtk6+0CnbZcnMV/1Dnbw1CZaz1q0yiz6/F8A8HBSelhjvYlY5HqQ6HN
j3s/mjcB5PxkapfwZnMEZ4kYid4/VIecG3jP1WbGiib15BUwN4aCa4XjP/j0tWtv
/VRHlwYrmpOpxpfhoWNKzgW0UOJR0w4Mmnep6v3PreBuhuD5eCyhrnoyuRDJ173q
Yn6z6a4o/KVlmDMJqg9tzzYNNTyfdb8EW0oupQ/5FFOxDEVamoWjqcLDIwdLe3KI
2QkiKw0bJXdOk7Q3S4/pJqsVkCNmWH4Cl7MBsPNFWiMnvSFHEQuXlE7MPXxTaZGo
6U+ai3B+MAfSXa2fDhGjrFUc8y9Ok4970CF/ViXLTLGT3q3KvG5tUYpY20dPpql4
H31iUT1AdkL+hUyvbUk+rofHdg1mHooK9KetO81AdRgwnWtMjYd7jFYg6JJFpBqv
GV223xM/hZiPvw8Rgs7mqhcKG430o4t9GBdvCrPYqeU+X8DK8ZIxGMTWFfvp7WJ1
EH9mciDWBgzwsRfwgUsN8yq0ez+wVGiByxlUyn8o/HEYIAmmn0PFxBrCW+JEdH31
9S2YOzxiw5BrWYdDL25N2V0PI7fwGtAu6PNy4ZZ0KOOcgChuBGTxzjO1m2mn6ZYM
1UJldVnd2i108sdpHrmKVH+uUAYhGJVQoWyUZX1600Qj/yBJd+tNB2NoF/VKXJ8N
Rqjy5mv800LdwoI3oRLzhOakEpvAHn2L+wx5HA7N2hMF2VveiezOdDNlsgi10vcj
Yz2FqvZwSTcWvSo0Wuvii8YuKRx657twdFq2HhkcVhQ/OV/IaFk7hNPWb/xZX8/4
xc8I4rlstiFYbGKTHWFhR+c3gj/D/SQzGXN2eXvwhRE13ikm/TX4Pld13d8cOKO5
6kvoXU9Mna7fJn1QUyd1hiMOYDf792TG2W2vZ25RSYfhTpos9UvpFekLF5Baewvc
AXm+ni7qO0U7KnZFB0yxKlsUxvrQY0MMT+8gpKZQ6jiZlNBXxIZ+l+ONvsNTyswC
1dLR3lMKRKTSXzLIJsaZsjOLhMb8mrzQy4D3BOPN5BJM/tzGYXsL3XmVNlKP5CVo
t1NQdkeBq89qMg5mcV3ppEqBrZMStHFVQig3iWgWmovUKkkQ6kCEkSSL1XRGJ8Ko
1OptogmwREFgscpwwUnDX4S2hcBeRDNoQWOOp7yPfPR8g3CSx+5JIarXnzW2DRk0
Tl/RHzt4TYGHDftha3WTbYgV1wOyKVuagDe6R3awPE0xEUTbZ20um2KxMrSYgeLT
CQWFkkABvi6kbggAVsMXiKGmU0FhYp+iye3X42pHqJdDbenxqeYis/wbEAos10zi
hCcYhoQTQQgjOWPgFjkilsW+dM7ipTwWGsPjl0UjH4wM7CT7yh1HdlMvI3xeEbcf
F/TwU/wVu6TSE4OsiaauHPhGi0LRfAVhoXwvjHboZYkOIPEjeQyDIdf1p7YYwi/g
+zHYYwA/t90ZdweRdKLcGmBmUuCE/xNXkvfkdD9aImI1WuBssq3EPMBYpoa8RNxv
333f0Zknu+Cn9VBA315DBAhT7+897PU6BcPkpT0PIh+vO5W3F9uacVN2LzJUb2xr
f24IUrCbUu/9F1nN6s1w1QozWZ/YBvD6iTyTFTcZy8CrYRW8X9lb5AQr4g04x5rM
9NEHL6CBeSvsgGnqIS9r9ixINdCQ6ouF8UUkXteOtfC2vnJPst0BGGiIYeHupTSZ
3Xe4TfmHH1AoBr6fyNQFJedkx0BU+oQKU41hXXKQB1XiJLkwua44E3OK3DCM3e+M
YxPY2VrGTMjyTrDopntAazYuLdhON17TH3mtN9eYV8JXMuSIeoTbT1tgO2oZtOa4
NHV7gqSnXnEIVM6ZViqJFWGOZwwVFcKILWW2pOd0LXEE1D4EzJBms+AfSOFzMOmF
pdgAn16XMM+td6bGs02axWlqI+WbuEVs3hpMIkE2HsV3Ye24kv/zj7iis4UFN3jl
5zZdInxLMOXRSe/T9jN9UBTaTsYgRXHgE1Gt0uYz1zyPaUO85il9zCaXeK5tWsNl
k+qQg3MnQzjzBnf7mRlfJE8wbabSYIZDEJe2ToHE6Hp1Wg9blh2Vp4ORhnnC0zM5
nOh/2GLSIBhvGBH4G4tWNwm4yXdFezsdVy4F9cfsBOYrryOniJvLiAw0R9wnejiE
kmrffKyoAIAYdkIMAYc7EIREYcxS1GxQMd9znv5bYxx/9jVdAs4QmNmxxtEV1x+J
RbCWgzuLSK/iYlbee5kuoDODaVumHzQa9Ez6DnoKhLTFis4OlnYjcY7GFsgJrhSe
5zH0q2U+m2j5DMVizXE1YYP5EsasH6EUBQIq7xdRXLywXnT1HAzbfYcaKU55ujpz
03V4QGXAPX21QRVhpGsV7hvz+bgDYLifn2gq2wdTiuPnew8JUfD3oyCfVF96XgoK
L5eFvZR7lpr2ptpcA67v90/viY237Xp/tWDNDskUPMAO2T9Vwn7Iz43gY2Iwjo83
06vquwsb2iGw3RjPQmATQWBU70nJSUOeObA9J9xV365tKHv0jxj2vQyRRK4JUuFY
TFr2DTnHQn72yS9QY8yVhINfngNkHu3olwiXIiHaQlKg9NnD1agDfh8on3jiushV
AydlUC98hVoSWqIMLpLGw3FXL3jG9PoNh6mKCl4YfPJ9kwS1Pd4yZXW1ZpMIorsX
+H4nZBWXMGu69CrRJvUaMgJE+Q0P1G5ENc3KM4JGQA6fl4aeTYeTiW/v+v5lJFOC
2KZO+//RhK7gpC15rKZz02N5p2Q3D0hg9DaGuQ+dhNjKUuR0CcMKgZHNqKeTmkd6
aPTq/WRvGK5Vt4SXd6LVA1MLjkQPjGWGWDr3j6ioC7QQ0ZpGRL48XWvvRh/tA3k4
2uDsKsCM+UN+qTILdx39p/aIz97BKJXxITp79xcRLUzOZLfXj1Qlh9X6VGroMxq0
yBgTEfs+FjkpbtximeVSTsps4EBfLE2O9BAefN5uX/d4BCE7J5FpBgvFK82NLNp9
dDATTTERd8izBcDiWbRDCWoF5kfOQnc0+uxuR/zGfrTHh+6mCWaIzObYen3HqSy/
Rpjgz2nljCtdIXgTHDMOLSINod2OIoxqvxwH0qVEouNtxMVFP92+d5arX5Xglh8y
kkR5j2q1pekGOs25CtAER5ihV29IKJNrkjGa7gZb6b4GpYxi3ZL/YniSt69ccdXa
5KHu5/EpRR4rjGgOnW34Jdk1bTplNVFmLB5X36r8/h+gRkEDq0LYXJctH3hQTqBX
yusCUST0X/0hJIDOKnWotRA/12HMezMQXjGZrts82M+PXfVIqn4W6Qzc1ai5Jk+t
QqsUj1joZCGNARRDTyxRP5n60hIXPJ0LCRU6L5xfiUtQwVKTG8SMZ161HWpy6w9Q
QXpIQBKx/HyqpdyvZnKPtGwRDTsmns0W88HjECDxg4diVLEBlu8plyafAEQYilQT
0Siix5/oHB+8LIhLmPIdnHU6+xmIjQTl6TXvtcmOmxZWBkb0QsYLqHCYCZgUlvNc
ZjGCTgYmcwezfi4P4ps3qrqlke3btVnyzgrFiegKwkpOK8aPXqHS6eiJL/EgsSl/
YwL2oDTPeEfMbmkZqclSHQ6H5l7RPbKfuM+dXXK3Bbql2dvG+ZuoB+xHtoQl5rSO
blA0SMD2tonLnfwiE1LGMIzaNUigK6CGRslY7SsdtrLYgbdZ4m+PkwBhWmSplvyR
trse2V6+JPMixXMeNkJXORmkuRcR+7NB2qHyPjqaGk2dcCB2J01jNG9HgrfvFsKf
O12+Mbt3pXs7XH1nQxhZVGnZZoqzPpTBcu7yMJE1ZNvn5wBY9q/8ScwgaBKr9/v1
79iYpzk10IPhhWW4KFglQ/Qr110fty5YIM08isWRxQ8j3TYwpy9yH342YN5vKzJi
2GCysKEDR4dYUX0Lz20T0gre2sOrNMM7Dmi7JPMzdSHBkTLtMwd/HibG+MZKVpmk
muplwx9AyxJj35oay6e6D0oxdYz/lz/EH5FvUCuZ4L+wZn+CQWOZmOjyop951teO
1Pb01Rb154Cv5ql2D75RSbmPcWn7p8RowINTYDrLXagBIyOpYgVWCLCx0kLwaRqC
KP80QaBQXHmDKu5wV1Whpsufp9l82Qduh31SFawbsJLMtrx9VPgKie6ka2vRzgsO
QX9WMez+p5GQrqTixR7Qwso0XCYTcJwxR61U7sM+jqqVyi80H1ROyIHBA7QOZQKy
amV9orbsu2YNiUpjXiMqIpUQDaFe+6CTRquHfrZVlG9B456h/Lwg9Fdvq2VrGSQ7
+dooSti2J1Oi93sYTmH45Ltxib1FUgKWvH8ZaHdt2ND/M+rO90FtDZpwhNf+nzfz
AOOfTbOCb2PVsJ8V1VhUhmgghktnR32E28yj0k2u6tMvR0i9P5j2wy1guTwRcL2M
X5R0z49vuy+oEel3racLxcc4/xRukSQj5V9opfs6r3DxxBvF0/U2itwMI7wlr018
R/G2jaT16+GSxyCZ1+dr1I7W7EgCnNMcn/ChWDgNb51ATX7PFESVabfPnUdJ0kq7
2qYCM8QRT/ZJbQVNkGQOEoI0iE5VAx4Efgoji2NbKHlCvVA6gqdPpHVBC3s8gkXc
ZF4KtsHJeoQiKZKkCDSULO4KAZirHb4q7UocXJkz9I2CSPc28PWqih54fCbkLfXi
CDL9cLpbBZieR5aQhXq04BlSYy6Uv8r11Ujj4P/fKK8+pOjFste3fcMK+dW4cSt9
i04HJZ7CHSMiCqLoLu+JDxlo0tr/Hr4R+ssIJ/GtnU86KkGa+rwQIM1GId2Pxq47
DSbnFjhR5Oeaens6zVeFYsR/ImPt8bGrFwiFQYOXnH7fcpI1MLR1cgZzi+54mKyb
l3in8ImyFEQG3jszZ9rs9zlmlWfm/oGsO/YHcc7M2xNu02yuxOoOefmflsIg4RBK
HjqkPQRcLhCDokWHanwd5nJhNKL5NaHpJZUpFBJT0AaZJrs4JyM1sjFnY3Dmi7m6
g2hbwelvIlX9i3xRM7w8m8M5/Fn9zxUWVTkdB0vXq5RWjDdLqJ9vabKYrQwpwTgS
TG+HRE+SZbiLKAA20CiKfmNhXKztOxUDuk+mZqF1FWKc3n/4wszxNCojbFJLnT69
OxVLMCucYYYJeeU++uzLYps5gUbBkir1DIpIQTkbYPk3xjx/DswiX+YQR4Ic9NgC
xZ1tGBFObeemwxsTrou45/IX+RxhZaANOYDUP3dJ7Kn4ur+SlCneKzEL69w9RZ4x
ujgkRwsvi/6Uw//2weGDaDZGbyjaM+Ad7HFV1hwGz6KRdcff9L8LT/NJtJWBfUsT
QxPY7ps9VSpNQfCuIgYwtcrGBPs88Psqn4cZ+WMFimrpuIcTu6bRzqknFBDUh503
2A+zNPspYt5mTg/TAsyPldaDpkwZ+0/Yg44j7/RYm3gQRseYqIePWR1lhbCIzz+t
iNV6aiI/83kEyCbNXE/j2djhCZkaDQQUjRvfdVg0hruvJuYkbMX51NOncXTz57PG
40lXPJ0cJUz4Id5gdHZ0NWcdES5h/oMYrQopEF/ZGedyovQSSL0xjEUsOf/Dr/E8
yLSvheDpDYx3WubxObMA9XN3r8yTIot7iepagmx/ASh9UZj5vTDKxTDFFUi2RJvg
ynyhHzwey3KbmNjCJODNP8OnVvF+oRIMrTVhUaLTZs3bCzclKzxdwojVj4pUc+BQ
jvZWirZViSYdutyDUDTRBMj3FI+5NEyJ8VsGiEvtFbDYgpNyje/H+XpQISUMbpV5
Q3AgEcWNrVdl9yMhGjOwnjHaeBWg3OPBXTL3Wk73/l+hnIOAy6t8iPG4hhd3n68p
z1jtI0u+fdlAgZaZVP6CT7Y1Zw8OVcicUu4q7doOZZoPUplzMbu7vRdiNZYmIWH1
+Fems63BDGedKDbojzyT+sKQBlAO0QpO6XaAz/DTnsAt5Z7/QCpNXQB/RZf3KeUu
qt+9dAv/yCMhhg3vxgByDZN31p+f2iOTo/4Op20SXioOnwdbYZXszFq8x0Osdlzn
zY97+ZUMGt4h6vVg2R/XqRjp/5Vai7d/nNwHIwcFbDPVsIxZYWlnUfN8v9VP+Zpi
ylppzDkHOfpRetTdDgeO4ti3JJ1igBSFkd/Yo/vmZWDGt+zUbgcCuozgnGq2AVDU
CnXDiIpJPnUou+Ex3ozQ19Jua4FbohPUMRQFSKWt4ULby/PtUNdBuDSImjq6pVLy
aY18meVHtdAXvUremNMPuzE9Uw1iI6SS+ePnNwv/GgZ7ikSg9ntm2WA/vqR/R6Ry
nW3FS03NNWpgC+f7ZWMDxZ6i6Pfj+dQ1zGLZHibWRsa6fDlFhTcZJ8LMrnR4J/vJ
urKPSrTQ88f0dEYflp2Rr1aVsE95uNiVzvbx2T71aB7TgSCPKntx7zecR/fL1Q1g
5IQVVbcPXrXaOjF6daYicItlROJH2OD5dfDl+6oAAXzy/PtS6ePX1JICg1AhfS94
U3K5I3TSYZuG3Hus5IzBFHm2uWoZQVyEEFUERiJfOCmOWwBJYMQm4/BtKVwCtyP8
IUu3B+cLSBeGWMi9aKnDpwKx9gkJAVkAV927nmuXGMF5IHYKEXuDhidRELG31ZDC
TN54ApUC0gtRjFrn3z1xcY/AM3jOHZ8jrkOUHwZ9Jfo3sW1pZX1/eQgEFy2WPO0G
TUtO/985O9m/i+9Yv07QuVJSJ/N943AjtLDPffKZioY1bGjHgqfp/muPzdzD6f4R
0D/lB/aW86sUW7uBt3+c+LhxnQ9W+ehLXJE9ddGW0KnjCyFdR5gU+u2q59vzzWVh
nCySlpThvCTwbIiPA25z5AgodvQ8vZQTtFWZNYsDXt2OrXquXbZeDHwgAAkRvmPQ
Awpm00EaIhUToYbQjziQb/lHrugDpK7etXbFAG62AQSCMUrWKJgYHBoomDVOr4m9
J3huhb8ZQVDoy1HuKrXaaRstpJoJagET/M5DntCi5nrTbISWvoEPwawSSKjFF1vy
GGuSBXhJUElWfhME4mrT2QaCeuhjbCXh84e84+NblZJSixtM/2lYkX2Kpv6XiTGp
49jAoJHUqBXLKAhtCmJhnU9sADNAiVQyBMyfDwWfXVvBcmA582hYqBB3SMRj2+02
B16IcK/ClZcGv8w8BHSfpGrpXRpXJ9cjShMw3QRmZV35AQOmmalNWHTAwDKbJUXg
tTsgwPmWSM0NFejLh15bOlSuSwvzYIaPRzuOt4aE0GsrW3LXXRNaRl+rD/MrOlgB
PVRrNWeOpAgi5UQ/4NmQuCWfhDEwMexE4yzIqvRGQJ8J76LCKRJovg0YTTB2SORp
SfPeZcNP059U1tv1T9qF/xIbjl0Iouu8Qp/RtPdZoyIT3qBnCGgo8vnfuFnyUYrt
QTlOw3u1aJdqZiizOk4jKCIz0PQORozAxXvktLnOou1MtYG3QRhaR3t3+URiT4ui
VapYVEnBWIKp26ws1leYpg+Qpu3nHildK9/QpH7u0N5IfXwU32jLxXK4dkalFlUt
8h2/iUdMxnU9jh0RaeuYBiX8oSz5FSEEkExn8Xt/lbgcIcbKOqrVlvqqTlV8THsO
1iGuLeVjmjA5XpTO8cShnnJuYWJfQJ2LKYSH9DbZy21U8SGOi8dCkB7EtWOErsE+
ojGnBbsnHg8YJyQw2yBmyC7evBX/o4rQBR/oiCnSvk+Co1ZbK5E5HxCNP+XCUVgi
DjT0QYquFvhlEXD/Uv5qCZNr/AOuDy1H5jmjAoen1CfEopFEOG0KGlGZPa4ymr7w
+smeSCoBPqjThJMB9FgPJQcpXm3Ke9v5mX97LqGA82hJ3r4BisSLxMSOSsEeGSX3
r0bI2R93FKhoGY/3ZxTOyK28nXYl/sjc591nBGws9gqreiE/y5YjkfTZ3Lhevv2Q
mrIQc3DrR6QLL7d/AVC8hu4EP9R0tYaKYzkAyTmtWKuoMtCgmiLNOK8RIiaa+ciQ
hAmWXb1i4bLDnhkWSDnbqQL64WS2Aiv/S3SiYjUjsUn/Uf3iJr410Hx0Jf3BG3Zy
E0zH3mf3NwaMkExU0FQbfKFiQ6ajwPAv6Tjb9pT3883d2I0rpWO9g+5mEuduDVmH
7SmNjeJmkO6Rx6GpiZ5jmihPgpbT5tToIwSYJy/sJV/fzUtCCrclAzI0R9N1CAVD
WZnZJzlDJGF7zf1BiX/knc1DFIvxjDr/BAcY5g+nVS5tiWKHQw9Jtt4rMRYX0vqh
DLfXZQfD4ucLJdtGPXjlhFB2boDZGeUMFilkvdBBalSiuTWOaHGOfPKKc1PDSBgp
IHK8/0CZf0l9U/YZNnFrDOE9utVyhBWsqJMC1ZLn4LHCWXxDgLx8Kfva1HabiuhY
qD0971pZepxnDOn2mqbZaiN74gAGeE+tNEvX/JSnjOMeXjzE6Yt+gn9IIhz5NtGK
V5ZjhQ+1IYKvFJNPneSnXw5aud011DGbFOb61V3pRsFmEm3frLmf5gSMFOe/FLBV
Y7a19nLhBNyWMgYc5qem/PkR+JRB1ikhv9U0jTYdUMcgmO+Pn2sCW3K42LvQYGZR
xW1o7DK6pF9xujUK3USE3n/p2m3ZDedK8fsM9TcnqXBF2Ji2GxgjS2BaOGhNyelQ
PYcfIOJynr84hQxy2zZyvdpMrFrgjP00+BWFFTogT0bkvCNbhF2ghlZRNTGSS2Im
rY2Y4ZD6ez/E1g3f4uqWrIefOEUuLZYG2ssEYqACoiPj+9D3/aBqTgBdclPBJbAa
6ShfeXDdf97eIPk329poJLgDXpRwZ3sRKlpS3qjZ+vi49OxSopsRzaydDnm+b5V2
LRA19LWmeV+L58pE4V066+exMpIRjOLzGmWelZKYkcwBjSloT1cHhO3DrPYSRBow
DFfmNycIqUv9m3ldHS+xTsuYzBnabvbGuqz+tEyHycT5+CqrCwj+nrrrl2l61m5O
gL789zBhOis2oRb6EeX/7XHHOW8hDf/Ue8iWHeb5r0R9gc61Mbv/jPulQ3f4wsIo
U5lOgi1lMJiG9qvn0u5c30U4b4P0T1xK0Hquw9a0fQMsKrvY1O0m4AyXbfMXIHXA
cUAHfRSJ0zDH7loOZRyNCX8o+TlR5A09ML7xWIsCJ+RljvE7Td4Hrs+q1z7m/nZg
grYA9qCnZx2XA6WZ4brxkeDKufs08fqL+B6sXE01kEuK28sDOm59/uqhOxNeI9KJ
It8AbuVwUyvG3xzYJ3uiKf4OxwBrlNLgWhzF3BhKUa5hn9w8XJIDMlzohsREyVWh
VguammCNpVjF9XwU+i1e74TD6AIVYh4lyFEVstR1re839/SVWg0IR8ASvYrG+kfC
DvbwT07JFidcpDM/VFf/ME37zvmft7zDLAyemIlKrmjQ3uMyrshaskLhECOKzo/i
4cBU/Lo57N4Ke6tUPxzol88yxE8YRm7hx3njtpBud1suraNOKHIm0bnbTd1mjIh2
Cl9M6ZYKHxOxeXzhBD7wvuvIS9l96y7V1Zv8Nb8Cf9/qPAaCXVAu4zCWpUqKRqNn
Yi/ShvcUEbVGYJrxBjbUEyWSvbYzWq1N2uA/BOXXwLiT9wEeoKUQISq9z3vOduQS
yMfcvzFxr/dVrbUicgyjFTqyolRjoF00O/tRT+2ng8wewW6fmO6MJ7Hg4IlVbLP1
4dEKL+6B4QtlVleTha5/QbutANpZJUd2EZZtP8GLrKGzMoNb1BQHkvKEo2h9ACpH
cASewWs/1Xg8YBOJ1qQNmJXrahD/zSC6/34w4gBYJ/iZMa2zKU6HBawZxpaqHusl
sT/GDmufJrxhxclapIk4m6V4GO7DKCepXYI2f6o/oUbVHDLmFrsk/iDxvThIOFMt
qYyVXoG9Z30eeRdl31obf9Vkg2P4fvbMcrTN+LltYJaorIogBzDOPLQN9dFERy7Z
slHVM0h3Yvsjo0YN4N3xE9shA7jkLOBcTLUDC/fpcMZAJNEew686R6svTEi5llz/
x/ko3Tqxllwjw7zNzQifBwDnr4jMM9akg9GPBFiQdFEj3e3kPAOUV5XxIdDGT34V
qG2oNhwk6sD/tEYujYHm2AMvkRKJRw95gIypUADhM+qGmDk8zqJbQygUvabG1Zpq
VJfyS+Q4KsL+y9cd0zGzvZUejF6+lyHwFUrGH23yrBLSnbr6Lut3YJufDa7c90tk
L0rvrxwWMQrtnjyZtcOC4NKX4IGJuJMUpi02ONsWSjrckuzD3RJhlcpuMF0lRiUN
EmesN477q6mdaWXFDpveJO1wqdgHa1OKRP8rG0mCoMCWGSm/vu568zzF8Kaq/rYX
hhQs1p+dODSBm/tLKXmK8hwkhgiKDzRExpOnKepbszkLXUCN/IbAim3MqwIqqO8x
1VQqu8RG7gOJZKNEFESMAq7xmga+qcc9hsf+9P7QN8dXDWlc3/XQ7s+XIGkrRPUT
CrY0oD/xLNBfJt/KPizuvWPHNswbZ2bh0xc7vBW83BNO157tcMyah8L0Mph5e6cV
zeQUk44p1RQSBZ1VQ8q4h1ZgbKGuSvqkLvOeaKxufYHSTf3ESW5sKqhe4nYyUyL8
HrxFerdDEtLdHxhO4GwD0X9LZuIStTpFB7dUl2fXGmJHk0IiCKYiwafzKOxP+E4S
Zg486CkG1A7X4p/Z2fyccWmNb5H/Rz+XD4mmZL51miNvFGcw4Iw74bFZMLTF7MIx
7tRiPZEgHrdFNuiIo+49JNxoBpXhXJTBqBjDIjdvejNyRSxWgq5Kpbgc+cWYBBQd
wkfw2ytv+/NbKA5lItGIOypkrNCnuuLrhxarqKlm+MqVCgIZMDoYS4roPUlz65c3
c+a1BtOQ/tVEcI5QBxl7y9e98Fc7rtBtzfEciDCl+XY0pwMU3vdR1sV2g7f0DGyJ
W741xIEqEdk3GvCAUioEx3wTmEERBIRaN+qHTboUV3S12ITLxrRbRe7RBCNUEi5T
8Il+ICX8V6QtSNuVrXDXWBaOuPfxOtc6kBQto2aDQRU5J3IzxF4raLkspzEmGvpB
zX5tSizC0e53OjJl4WUJXQjlAcKYjmA5rq9HCqdEyQK4WnZQJ0hcvhz8e3yyFVLv
t8BPfHDdtakIJEMhMYYORcy+Hbmc7lyhqPVx3rf3YnvPkDOqjSCSPboBvrJqUaKr
nv/GNUB26WTrOGBPjZUfKMrud6iSW4NWjrRo4x82IK52T+v8Jf85seOAwwGcfKZn
hye3tzZlQ6xnZ78StK4ryAQ4fiN3UwPlIk9h3aBEeRVYttYUuYQo3AIlwI02kojR
2Vk4ddqnlRkKX3YIMQXjOaTU94VA6AHF4cM15KJNcV0fXeN+ArGtzVMSN5Thu7tN
u/9fGu0CtH1bOHKr0Nc3PPmXHUX40dOrnWz9tcJiKbGQ1m0aNR/539eh8sotslMA
C0gOokIRi6gTlrQ/cHEvdeAMwfuB+mFrP+9qWFYJ1Ogd1uwqunV9BCNJJBCl3fUG
dR+Ll6mDDWF1pK4sFCAyUQjHeX5P3+fVXjxWQtX3Zg8Jgk6Rr3fVsH9y3O+H2vBq
W5O8Nui8HO36KUYEuLK2N40mxn+BjFO0Ld+MmQVt2Y5uvl37I9EUPmeflycaakmU
5Xr8yYyXD/2d9aZFj5fF9+jE4+U3kQXlAl9K72tKJmhkSfLs0sg4F1LHaHzBQcD0
T4DpD7zrYR7Fb2dhowJ7ZylpZLDAJhd6RZt+5oVDfIZ40j48uRmhwHdO+6ZWdYiI
ZOTlWYBOBlxybFoKX7wc/z88sd4vg1xBaR2CIzRuNhIXueBAtl1cuvhX2qHUu/Bv
RYGToXyXsR3LZre+qHwkdUw2S80HCyQ753fbXrabSd19bJeKfxpd19h5jiNEpcZ3
uiHL2OeL3iQJ7NhO1YqkRHi700qU33qfiic6A9vXEYKaJGk7dPQVB1GH34V22OLN
pSlZr1DDEC7fjdd0biR+6quhUBpXTvK10IMROopRDUYXrZ+mpvmqOlejdbWGedCE
fNPsNDS8pPotucJD61vaqFGialAT7V+9xMSS1hJb96VSk+v2mflAtygpMFvYHhML
AzDweJ7BNTs4MlFKR25F8Albe4zywv9LjjdjfIKL+hFv3Rsja1NSczgag7Rvi0zP
5tKGxu6CGda82swruj+rWEFBBGOen8azxrnXIuNso8TUsZ6NyQon5V/sbR6FOwFL
6oDoVH5Vjbaawz91QkT+ozv+t70/xBkhBu+JPMbdcuUL5bI7wcUFJUOHKA+E0x7i
1CelPrs/ve4/6FTaDHwQuWiyyKKyR7CtLUgwiNXV15FO4nmZzMHsBNsx9abWcoj6
N6k1TOE1K+tm/JSoJsxiJ5Yb1LMbC8G3Xmgwj+y98IKFjrVyjns9nZo/q2WnDvrc
Qa5D/sJ9JL1OWjWs6HOmVGt5tJf74GCH86TeU/jG38bsfpKM7Re7lllcGfADSy41
PzyOEl5GIl/vPIBApF3jS9kPpl6zk3tzagRsIMBhKp9bahQy+IZXp3PGDjLyDo7O
4rJ0tLdBz2OYbSSsSgs/U8OiQw/BY4hQi8Abo4t61GkJcSHhbyc6PHMVPpt4OJ6m
81R9JfL2wiQmh7tfWFzBryqxTDkvGi9HaOTKbjYQGggpZ2qjyInE279Tz9OOF6Vt
RWi8Dx3bq5m9sKr4Uy08+e+kvirPfIVXNM3YqvX5hTP5a3M40OGtr2HfVWODK+tl
v3fC1xmWnjQPGgzZCbdH+uSRx1Fu2CEflkZtCO6suZt4JTLFbk8iWotSY4kr9mb5
MybQsqCtYe9fHkU3mdZrwrwW8Zg1+tH/Wlvp/7AstyUpQjzig5wTQmhLrlo3MsPz
gtYelqmBt00cOS6IVtMVRyiH2T/96eElEmMNUAlWrgBL5sie0JgnnZhvJ8HNMMP6
PPNSno3+qp0Uttc8UAAJrR9zSmQqdX1XT3+Xoc+15eDbNbeMkACaMtYkj0NdasKH
foPxn3cv6QdfKyWxpd3wsxskW/gnwhP7AZWLF0hSZ4WatGUhvXPuXRi4DhkWL4bo
U6KKXYYcaxkjp6O1ik/AtQuTDsi+b5oE+qYPMqAnXrEbrynISXIpfnPMFY5/0NNF
FS2Ek4zpjoEuSLwyCC+HdiiBaQ8GOCKzpWN4r+O7HkMln4IXb1UZYT3+q8Z4EwMj
cvUMJsaEND3YcNsy1xRPWHhsyu36GuGhlvolpWQX3kJBk0Pt33HsUtmdqqkGLASS
fcrfhP+WoE2damjfAkdJKapLN9JmBDRgmfQQcvfTapwncJI7Bo9wi+mHjOOkf/W9
LxW77tKGQlriakcLF7K+w2cCkrX0gbOZgm8TgYKc8G8B6KrqD+5jP/UtXD/1uLyp
h6rKyrf89QjscbWGAp4IlkALTWdk6z8CxscCC8ZYxtV6Ye9jnzTIQHCtgl6DK1KP
0pFrunY+7F/aXto93HHhF71DYQWZHIY5vm8oROYqvqHwapOJUqM2TGNnllz2vrmG
ypXIMee65bHQFObThKgrivPT0/tq/6x4RSL3a3c/g4CWVoeEeugW7nNw5tOAVBJq
1vIvpLG+u5CQr7VFQ6jogGuoilvfrhlSj67hHW2u6mnROBAgXpjIh2c8yZYmnK2p
4kKvqdrmRFAVSnhfc1+DwSCVgHwr78kb7wB9l5ahkF3RHrO2njkbaevoCjK1ZFa7
1G+6/0x7HbYOq83rPJvr1+GcNQwRzYuJFivLqKZBS6z4c/DUHgCHEYKSVOmU5WI0
QV10wLh3rlCPRevf11vPACHCAuo7mckYcIpOI/nwF0qEQfljJCpwB1Jw9hVHtFlC
KVBsseypYkZsfOcZdhca3OcGA9lmxWdfrbbeA4G5jtmfZ4AhDEvrxLQheNE9N21Z
U5GoYPBmSde4DGekOHps9N9Rqa1zVGfKogTQT2Dq1Sm07hw5+gjobAimaDZ9RcZZ
TCmWVsPnuUyucEBbEzKQsXmVtqhPwl+hGT0CkUg9tK4uPNNuw6+/E+TP2iIbCOlj
Njp1S0YCaHTmBScTydqEqPpuP0DoSVvNaTPgmtd75ku3CCtjCXYEx1mFVPDKu/vV
MxQxsxWPTtDoI2bDkuV30bcLqkLip94VEyVl0uXQKopd+qMYMeNuC6B0mJmN2yoL
ErZbmOT0RZYPnZAU7fOqGCKXVg+I53H12OcFdqslEwkAydfqxKQd0EWIW5HOcWbq
Z6dzb0W+7cXK32FWJbzDrjXexWgNQHhh2ZJvObOLKIV2+8ZURZK7M6DHe+ArHEAM
IXt9D5Zf04xBK/40lO/npwDQtv7mt+sog7NLDgICvitIbLmd2rHw8aqHM94vPRav
Mgwi69dJ8Ve5swPMkTfcmcROEa042g7+6WxHtuY7Wr7iuAKq9m+4E4bZco3oqq8j
vP3aaYhey9N7KnnTppDnApMaqtUWirzF1Wv7fOMVbhxuS21QK8q/Xz1qP4cL619l
QE10yW/b/bWsiq6AUVifxyL4L+d3+7dySTeQughTGIdNPMSBDKFRzJ4ibLCSBSbG
F4pHlQvQqsDIKW2XGCdyBYmkMjXjX3s6SzYk4nG2JvTfEzbYM+xjiZP+qac3FUQy
FrYUrQc0xiU8sTcdT7JwH1KnzfFJDRfws6DCZlU6r4uAywSkvS4Rsi4oSTtMwrnH
b/O9WvfZspq6FH1fIa7XGQ6AWEueJzT0oIhNFIgx5Ee96uMLVrimypNHce/so1Nl
L8AVY3RD/jfl9b8PbZLJIh2zHSgSUpspE6M0upgowzlNIEYu7mrH6BTLRj1hFIPb
Z/7lw1kByPbMHq6VPBY+lq9PjaBDHBk9VqL8zvAIuYOhtWi5V5d2Jvy+Z7ZS1N0f
DEOA3uSLOeYsnWl8X7Fu2S43kU+yFp3XNOwTGT1pSq66uknryJgN4Vjd5wcgoPsk
jfjs/ZFCLM8c5eEFXrbeMlW//9VR3BZEY2MG12HUVIDwg9NRYtYhlYaPGb2YoHxC
jJua6sYkZ07UTqs1DMOXy7wr8c8M8vM0q7E9Ao0Ykor+HgpzapgZQlm78DcOFXnS
ysCBi4SSDGEvJ5zs3T4ZA6k5jTmFGiAFPJ0A9j0ZF/xhZzPNwgsT2KdxYAzsrC5i
mehJ0GGO1uc5P3FoCIe/4RxtKIIqIq83n7Zc8AmxwFxKBRU9AwFF1EaHDMeCZh24
p6+ibHe3Pro+vf0alv0numaBcQWa6j565r7TMtfjmmIMN5NwW6tXc5cQr/zGOI+m
NAWOQ2uU5hqnH6bctl8BfAnUe/RL3qy9MaC97RcyaK/vnFic5zjbeQczekOTzRb7
mLANnDlbpOR77KUTD9qYg3cOVS6BhEtQSXSdg0FkCHHw3V2sMKgCEDsgDUv6UI9N
U22QRpyanCMZua6nmXvJNnwbIFhqI3z2MbkE8dpCXip2j/0sdmKC3IUyfXVcceIi
6WA7pJaR4iSLEsyz3v7550xyJwvm1MG0upys1U3AdNxeWa5DHedpRvXG1TW42p47
bHNbRDNhrKj5M5cU2mTR7/9Q+pRuejmQBFIqzHtIMxKQk4g2l5qoaOexO3HFyhRr
eFcJa/Mx6Yqt2J2C36rm5mzJDnhmQWjdghtmJP4iApW1oULVUIOiI1uRz68jV0vY
4rpgzZMxKV6c31HYu9OoOf9fCSSSIXDi7s0edvc8vGRaJ0gAylKT2LwzlQ0PYkem
kgLHTuecooWwNr/QtlPNlFsBP354kfyQZdIIqZZQH81S3GsJM4hMcLb+BpdW6Q5r
UfW7xz/RROUnNl9CCE/lZj5DuJY3YmykwErvwTBBHKfqPnbHdLo0z1nF6PxOMnzJ
uXnyF9AwKufFzC7RbT6h85zYqRQXDNxrcBNiEGTBgCIM5j+AuGEWrGyWy267W9y1
kms/0jpa6rFVFTTkgiaKuW+eNHnQ+KE63VKqLNJeC4Okso0kesHtikKy43JKpoMO
eFQ9QR2A8U3N2f2r1/+mNU6yE93mHTJ5LIxapqwYDim+y3rAjT6rKH3vVgiVo3kI
9nkCFw3GaGxOVOCfLGaRTXxW90uOTb+2HTyDK+zdhbBAm2ivc5rYu145UR+U56rq
cdmjZKbILsYb70gXvxCtpYt66hWeHnvKuJgWiNYfDBsXJXDcmfbAvVuQUycSGqNd
9NcxW/TAU+R74nGNNluQwBY/GiM00mc44t9jS2GXIspVvX+h6VcI0trPMKmxbofD
MPtSf/hJRe/c1rL+qS1qrCqk/n4rM5RAEqqMAh+31Ak84PB4r4MR1y3Zqp6Utk2+
JrQU5xb6hwMqx1z/jAYrSTfhsoXNzaNmBSuAxgEiVppurkeA51h+iyaB3Zq1/Tw2
anR/wwrzz9R5H02cbLfeUxZAZ//gHjjoUV0KLDpUweH7+mp7y6R0qqdnksDTwa3W
z3HD70GbYqzgBkdgjdtDb1DrWjXJCnNHXXQdY+U0f01BEK0V577Sckht2X6EGDWw
jRr3VWSBEQEkB5Ijo0NBJePkzibNaanKRYIJ91t9Zr+Wqk+fHIx4aaNXzZTQMNXE
zcxrEl8uV0C4LHz3WvED3GoeS1iZBVNk88j76eJBDbEsXllAt4FiJRw9ZhC4K2b4
NpzBFPTXZNUvvuCA4e1ku2LDfv6SluX38B876CgpL3l9IpqH6UuhaJL1pN0wfS/Q
ZI8JvNg95kTDodVLn0o0nWEaOFJy82wIQhd7qr1OkbPzGugwsfev1acQMzhepTjr
Zk1F3OL4NvB+ll7TblAKnJNuqY4/Ci1vt2cJ4D2eLnAtsm7vVqgY3OhbLYXLLtYh
6dITQ9Jag837Q+JdM7pO3Au3ZiQNnXfXgkRmw6z6F3TMxNLLoSB5ys5IuoB4lorv
rKmgU07Jjg+/gOX35VQa/xi0KQDmDRiZJayudb4jDh7jMwdIIMEq5p2/ulQvH1Zn
zr+WXa2y4tEE7a6Op86HvBBcKihMwSGWHcD2VNPyQOpIvrivoEKItdNZr0EaErcL
A6cW61Db6D/V5BA0kZYQQ44w6ZvCWXm5VF1v1MhCZNeOdiWSpsDGv4PRSgAzv1k6
4b+uCOdXhgeR1DBf6/+zFLNP6ZyM0LVROrePpo2JrPX1WDOWv4GK82P8w99WJtiw
U8vAmPkJszCsm20OfI9f/LJQQPMNpasD1kP2pKZnXlMP8o1tA6/6qi6IJBvedRUw
a8cCRyUIodjMjUhpCsevwvTmLXtvjKaZU+pYa1rH8CINi/pVQq8/lVQ1saXZo8PP
gdtP4o7SeOIxWfzxCUpFHcb8Re5NapFUrIQjq/uKy0iS4QzfTWsrjUCr1Jw6vFUt
MndBcnqgmKVPHPuhf4piK8icY1NfiwP+adeLb4cFcIsTrCf7iaKnP+fBIP++FSyf
p8atpcSp8OYxtz6Vj3D80cP1c+Hoq3XlMbOC5tPugmuG8w4Yv4fhCDYkj0/uoYLI
iSt/nA8k16bgqjLAdPzVnsdbvBhCcMm4xI2IvSZJVAEpn6iMSQq3NPRiS9UrjONU
IKKrQbbQBMd59xQEfcOORosMnu8vj0sLeUlE7S6o7Pl07s6Mgu6iu3tW2ex8mwIN
iXnkuVYvD8m2P6EWtylISlygv/BfFDqFmv4UapzJZ/pzh7LEpO2O5zCZOSMNTEs3
/kvoChgPvliRfhr9fJjvdJiH4OGrMwImZA7HD4M9vYYSniH6KwgSCQmrpfYkhfq8
8IrTmWUhNdqjpM2o8SSYA6mEx39FiCJo/VFNUswhiVMYkVLvhiF4RDBDhDBAgbHH
dVvaUqzOlPtXsXhqyHIBsknDU0xiClwzZIZdjJYDKmOHxGrx/ar7xd05sap7bkyU
CwsG/uBfiPaPRJjHP45LZtHbw/W5ZzjOBw/th+DVI/Sb4dcv9HfTxbU3LDRjp3ee
P/lVAKBOaUF+Y38/RVf6y7YihCUaMVgHf6b7FD98CGqwR491fDe44YHaGPd++M8k
NRFvQ1BX9gtNbKepCUbO1ZOp1AxpmB2QXnkZgHC5zvSJBn2wxF/r48IvPS5rZyGS
XhgaLhnPcNU/ylViV6wqZp0DKJfVMUeMwmKE/yN7Mh/8bD/Wzbppa56eLitMvj4N
/j8hdHgzOB070B9XMd5ORRdMA59jUXuBjcELswibz4esZlwiKv2cyirt+rQyofnA
NMKExAuQP9iEIhbP1D6qdjhcj+9H8B54VbqtWSpRWA3q9qbN1oXYc8J2wP2ab3Fw
z5LWHYFsYt7FATHZHUuPQ4Q/HWRXZ8YDHMwpvbWfvCo+mWComHWNNvczua9rSqRH
dxPQK/0OBLGET26RJ5UGQOTUDP0LeiB8mhG/hpfQNsY9084HEjiFfPH/5mr5AXmn
878iMEi+U164ArNftFmOcHqcZkoTA9wSakmaRzXLaJ694aebY72AyDXag5yubUtp
mVQeId/+a5YxGoAMXatnpUqPF+ISJ04SxpMc++nt2gCIBvZvMH87ndGH0I7zcNvf
8zstsnRNslyeoCWPsVDYq1F6vXFZMYmvfx3dlAo7bAqIn/bCo/6W0yFE0prqmFKy
HcxiOB8t11baRsFt5J/nytIqjFh1CDCXmqDQF0+IVlWCxYZg0uQcVPX7iYWhLoJ6
ksBHvRA/pCo64KPFzkV6s2uF8pzMZ10issSzaH+tLAPujAq+i8wzbYHG41I+vG+L
1cR8TRgZ7D23x76Jp2+nFb3bG9dy/+8HpprgpJUnleksXx1TnNpRLmIVkcFJfbB4
7B9K++p8fHfOxSA5F5vX02J5Lxl0v+KRmaB+tRUgtKYDUzy9nnz0rj3hNwgXcOFD
EMxbnsPDuuMYjflYd5NCQOZLCEyqeevSbhXmUlyZzTcmV9NTjfPkgYBR7EXo+kYg
7/qNo5qWjK+G1g36jgwun4lCWX0fsFzhc/k/+oODzQtBln7s31KPRlzbmFCyXjT3
yn8b4Q6HSbYS1WD1E9wgMuErga1WZnQStmq5Kjm/BPURBwz+pkS6y6bBfpWPzUyD
0rJ1xTsg2oC8jf/Oer/y+mYOTZf+z4Dm9ag4pUBmHe4YZxyCADKqyfkAqzVJVGDe
FInphKnfPtqC3bVN78JWUyeh3QNNP11wFdzH0Z3aYj/sSlpGTVbFVGDdvCqEbVjk
amD6xxiQpqj+zhbJIZVlVSi9A2zWFNJgTr4M2jBziZGQ+xQfYXYVxTkGApPm809e
h/sADJ9M5ab/VK+XkyYbtQJlmGZMPYGUCdCU2QRVZFWFqRf+U+k059VmLGytJ2np
/TXpohFiaCcFoIzU23C6gAxYn9brI5bgJkUByDaqO7vi9XZVh+uZZYTbto8itZvz
xNYON1RoA0DoCl+o7zt2ek31f3kcFFC29Cj7m9MXrjwdqqOLL8vkMsWrK5f7Z0iJ
enMFtNr91EuBmI1tH/BTVEo/JSrr7yZ7MGP4yTaiVZrLpnS8KHsYmmD4O6mmlyd9
ecXlv2uIUaJ/r3E0+LG0URIVXHol8NReBNixgyeuXL+DigwWariDWVXRGwvjHNn7
39uPHvjcvQAbX+9vmXoEuSSkwtOBz5T6kJ1Fn6GYuvhjk12HpBrIkbW2MzFL4444
T/HGqJ1DylpQ6pVIPoypP4rL/MayTW+R3EPq1AGH05ArYOmU3NS6z70OIASHGfcv
QY4B8C07exHZXIh5R1Yg+mplEqBh5VNWwgSAHU+Ht4nBxKYVOMpPH4QMRGzukBde
QEE46o1BFF44K9YXRmgc22OtPIFi2rPKmYjtgAh9izM7/bSZ0ZsVPzq/nTtFniMC
lqm9mxgQLxGBkmqVWKqUQh7QABU79BiDQXnMgiVyqBWYF++EFHsLU1F9H0DIC2uX
Lz6f+jKcf9TptvgNgfWb3R1xHs0+QJd8Ag93vbVpHCvMgJ3V8oGQ8bw/OPNpWx8s
LtQfNvUmUNkBCo9HUnoKUIvQoNKJOJaVkxr1WTr1abcVMTABehiocwt/2lVgASOq
iNXKEHd8WjZyxQfbfh0nDGifb1xeJyJD/zilFEpW8i/26UKOpflGgyuLDKZoVSgC
cOceuwxGpRt4kmIo1UOwg/HJOYK5mhsJfj8lq4jLQf7HItk9C+xV4senE4D3NFkk
M2ZWidXaD3+j3C2G0ZUi6SgKkc4hknmdSH6i4CpfnT9BbBGrq5mX3om1luKiTGfQ
oI8amWFBmnw6SVqgv7RhKp5mgXlZ7VA2dAuBZjk1T28gDv6LraHVW02aJtl2EppZ
oLocxX2GOrzM25F5q+e87lDoK92p3gYC+Dz5whXxWxyjk9prS8NnSgoZ7iENA+Hy
e40I8zfD/F+hXGv8It2Qptd2j+6A2KJMNy3ucUMwg/w4w6lpWQax4R3wNHaoaz5m
7RpBkVz2mjbKQv7q2aRC1/813qqeDI9zwr+Crac38AreLuoo2pzYOsGciE+HUe7B
nssMYaqpkR3kbagKo+vNWS4Pm2/pgoPyOWR+yjjlq3oqgyH7FHRnTPVnTfdKNkzR
5bRyGS583nNUmX1aesheLDDeAs5f++/yjQ2mq0eYBo2XlfbJLNTnySWkNwYvrA+4
UJ+LYQB6wJjfxMgO4lsSmAm967URuYCzKILqmwaiTzxR8XkLniDP9Z4dsN2voyFK
DYsoBVUrB4uKsCVfGAK1zTvN8y9fGVJ0cTjAyGMQ95Tl61696IpXJePfxD7Tyk6u
3CRSt/adkwdjwYnq/NYXa2gQ2hxmKUkQnxngA48Wo4gvDWc9tXY3npWhYS2tuhSS
+tmXzOKkcvDw138c22sx+tCPV6ZBgPysTBXEpC2OChSP01xyBlS+N51wziJIOqlA
jM4nmPKzfU/0XUmpIgQUMh9QWzE7a475taiuM2NA8yDNVrb0/Qwxq6jvEWtnes9s
lfJ5l5yW245NthVyujTt/8z+nwhpPG0HyC62CWscmmduMFUZZyK1W+CiO11MfpjL
eID3Y0YOcOcQrD66u1+0tZ7wRRlSGe33DLPFAP9AzMXF1UHymhfCmcw6FhouOR8o
wr2Ea7/aD+BNOIti4r5hEc+i4U76EMWdM8wWIO6sbrnixZ1QkJzf9mFzYY4dhlEi
pOgBkZhsNFq0zUddVk+onv8RgilgaARg0OQv7UFt3O1ApsjBTySzNHD+Zwct/7GY
2YcMDIpu2UuELvAmtC5duZAsaigWkNcE+gycnvSRxvObVfKxc6i3OcZe9OQ0+SCy
1uJuGbWsAUYmG2mVasYFCthI4LNV/SJz1U7bBBQ6thETBrPKq25juMSjZ+ODDlD6
Y39cTmtS4qrorR8RuKRAFKUTwwunIofsSh4+EGZZRvSZWovSA89qSzIiOoweY15+
cry4sXjhAS4QJXgRCfbiMypDiiBNOpjKU7KH3E2w42TX4MqvPapRm5Ax9yeaMzNF
3hmSAYD4K/Elx10DJ/CaE9Pj1xpKA4u+sWcIHrBY9ACiZOKJz6jWZqYk5Xdyt1cA
0ZHjEFyB9A74q/di9z+YxcsbIQFoK6PON5sb3R9YRTzytrhkBEk5hWaYKCAL4fOi
C2QaflfX0o1YF098PRUk70GbUnbskWQFd7/OzKs0Eriw/PrpN8+bw2p1KbtCTMbm
aVTKDKRniiTqd/chIrG2/Prz0V1Wv02pEhtiE7mEwHkRtl3099I//yRjLS/SH+HU
SAlydFl9bWfbcENdFRAhulSzMoQlbI5q+o1FgvXebmH4eTJ9TCrruIcd9u1RiVql
Y1vLISn6wvlGMzCYIaHatw9Ox/dnm94u97G8hZY0RWQNEEomCx63PDb3RGHaOGUE
lUMxJ2Zi6EKrUSAdxMEa0yVmzwNPeww6l87ExMnogQjOx7E20XRnQhsJhH31L6wS
L8pN61gMclKvo/kOsi3LUK5NdCCjvq73e/EVjZHeUMgSImdAOIBK1gieLylrnvoc
qm9fc9yUZ3KQz0ic3twr0Eb0cZVDn+MufLDBcP6jAmdVVUW2J1LoblyJiuZ6i2qM
Dm271tk1IlwkTD2h87hsCvnwJfiK0rgRzmKEWp76CEVjGR/+5klf7ojuVFRbbPZg
IPuVdnLneUFVLymvTDuPqc7wuym+UMdvWcKEMD8UPVl9pJhJuqdlwDu6+T2344xm
hb1sGCrsEBzzBDmCaA3gGYfZFnHeGNAZXJ8T/+fwM+k4fUZ4YVJCmC7jlKF0Q7cL
nlB3K03FE576NwJiMS9M2HvsNB2IVWHziMdCTGDjtWSwN4/qr7QmT75jYJAVLWio
nfX12hwB972nrUPGjRIptU6iAS9KP0/YINDcj2WZRaPuhI8Cq2C0y3se63zeFvVS
A5WixhmEb3672Dfi5AD6l4xZi/JrI/KcFs0NHBEf6G2U/KaeBRr89nutbffcZZzi
Liw07DWa/HL+R96geKagOCnupvg8c4KCGyOODn/bYJRu/rf8mTcXNTbYTGCY4rMc
KJKW9zcm3mzWUQPy4irDFW3UbPtbIbQPU1oDpwJbne2FAEfM7GYvM++cl1nScOJJ
nDJuADcig8DQRzE81UGXJf2ym1sLOcEBlB8axHIsbWBmH7fH6qWAyfbOXhs3TtmT
5wuGjtxbemQjSKcePfNiRHLzIWM2Sv9l3YetolqTm+roV4ZICrooVjomC/sZLm8n
2gSs1aA6P24L85BXtzTZaBCvg3+mZjCrbxKVKSJuB6Tb2sfodrhf95lWnryufPtx
3xzI3Kf20ogwvYiP65JwkxoaPVZ0YF3YhNzGjpz+vRc3+k86HGlBjCn30dYvuGnP
ITyLayV/dK3pvp0YwySFZY+rPgREO5IfMPkXNZso1NCZAYtHKGpSPHtcerbTOZLj
J7OiVj8Q4Dc8LMLrheSl+DKi0RDbRLE/ATK4vPt0+joFQP9lac2ZvO23nwzggHnc
N0tlhjmzUzN4bRHXl1S+GGVVykLuhiOxV25WPqwwp42K2BiZn/AVGovFE9giMC6r
cMe8zkfl6tyFWOHCetf5hRXH1ggDW+LAjp0gZ2+Y6C7NtzSN0mvTm3kE4/QKPcKk
4GocdvTeKJoOAPfFEpctUV9EwQTWsaKCAR+AIlRd3hxEmUJLonLMEVJAo0vq5VhI
Er5LhMMwX79Nvwe3unc0YXKjYunE5VDrY4PP15YygmhHVVVhtJ0tCM5qaixOpksA
0keUs/ZfN4Z0chK7LG4XMy093VvKQICd/dgALbpCIOlghBNV4xGuPT7H2tTG5FNS
PF30/BFv/Gtl5SP3l4Fk8jvCMNeyxMAwwXEmZJDMsFM8tFheVcLoeZrosu2CMApi
1FbRtXPxw8+zNS6lN3bzNMI2h3znnyf0Rj/lSA1b17JwH3bwymtY8t09xE/3WfdS
c7N0BQuMqcwHj15puRhIKCTkgZjVcc3jpoMuAJvqaRG7Ufayv3d4J6Fb2AksvHlN
jpxxSPNtLIfswfLjJ7xOQzXOiZns4T9ozWiOKZS6GV1sN2zce9swEtK9Q2sspm89
soNjwac59gb6RGLRrD81LVbP+FwiZRkzA1iGmOUxjf1qctP7jjBc4HpzNSQJhaHD
h9JKBC03bQoZDiBotoPOZ39HMCLqEl+LOicyRchnibw/t7DWNcANgOK9tclDpODe
1POFAscIkpdy8yhKU/FtDjnDepxC7P5scF4k2GKDSg5rsobQEQ9jKFToGEt4b+mB
/6459v5UbiJWmNUHxiVPBhpr6T2C+jrlSEFXqinL3tStICQf/qgUllZsKRtmulVQ
7KmBQzI9Anh9RJEPTdUAcbfaQAGDKAkS6dGBgqrJEcjzftwAx613AYlv7i1CwRl8
NTM9W3S2bcp4mJh6Adv9UGkNZoohJ7hZQDH8lvWo/n0MLF42JWEB5q0eXXCqLgjX
hX4HjGTUh5ivxaWu1b5TrRn6JLreCl1U5F7sohtQmCU7sv+E+hTQz1G2fz8TafLM
ce83hzTzt2eUDvq99SrCmSHZYs+IwudJRUY/mKtQFKykqMXotZjfAuAXE0meF4ZF
UdqSh7SO0lt6Dnq6E4m/o2lzmxwO0PUtjqcZ5a/lC0ANFDQT0DpM/tXG6D03xpHU
MA56NafZXVQacPWJVB+SJwSTg7J0iTu3Zz58oul7NOWgLCFzV0JDM4e8ZfE2MQHk
d1plDMSLeBndSOTaDOcNh2CEXe2BaqYyVgHt54V2sT6c9tQIGudwR/dD0xotMYkC
7awqYx2dGgW7qDaK8P72NIEKpys7s6cO2urL41hnWDOVQ+kx6H2W/jyDiR4hOjGy
GC//nwf1856nsFiyqyHsOnvLYBLutdc30K4fOYAd54vJMpAhnXmaDbqQue0Vsq57
WAx+ObmsKAeqlfuEPN47MVLEl2ghnxe8M9SgaaJX/jpf7iDktRh/HTnnlTuxTF+j
DLd0m1u4arvVFBtXYKkeF9HQZkRWdmr0G/jSXPNz9cvwHM6v7XKrL7inx8FswyrI
i1ghmX1nvK1gPyg6yJlTucdapPb5fcMJzXi1U/+p3++mghTo98aTt4mDkadwcbsc
46jlQhhghLm1T8S3IdD+x76aqszmrRsYCrZ13hu5LtPn/XmUJmzFAEzjfzK6ZedN
2rymfdTviLsEhTmo7rZ2Shx3BPpqXzwajjsVNBu4ClCw9vYNz7WMDiDmzXaiz5RG
1o2qbUeMDovh/q2aPK6CD53xE69JCcKgLN7kKAnWnCDyXZy3t9kl5l7zNcWTYZhD
MRRenR24OSDuxeMQdxxKJejOtQhZbNNZsjYUe+IIJJKf9sEnONL16AEmpWbXtnz7
Z5nCjocuaFMuMgvfi5iLC8rffkLhfqN15upw7I0lh+8eQPrk5glLI+6NBHe7wmVS
8wUtL2ap8i6pL0bFmETx312kfDlSh+uf5AjVyq8/x9sacGkTNx/hMVFxVZleh6V2
Im1SNivtH1V5pThZnqA5ylQ2FU3W2nTsyrgga62kKeiFENW3visWXBKqJHJO7y+I
HpHfdmeWBEg2PG0sJmkYBMTpY1rlkNcy41pjc/zr5Bq5XwwUroaa96nfW1VAunrC
uaUE/xaJP6h/WFnzAjJBlGd7ns+LcY36eD5Mj2pwKA3rkuT3CDvnBUmQ9qBnUX5z
Gta4Q5X5sDo36Fj/dEpmDZaTRc832nnK9UfAQ3Qy2O21Q+/RxH6sFlyxs0y/14Q7
OknoBwWEsMpK/pJyJoIfvLeDq9n66ru6yFNH2Ukj2w6GwnV/4Xl8OSPAivKCAjqG
mN8fwO/5ZexVGl9hDTeSaDBLBm0K+mBL/IJrxQmK69uQWqgwp6MwbO8F4recj/2O
iFf2+m6NCRkwR1qKXbK+yYSRghwZC0YKz1zyEmMdAjRkEQe89/+TXCslVaugkTzy
JzUeQZKQdUjQHdwsT1VwYeVD9h0RZ2eVv0O6/dFyMwv7Tmq1uhOtem0tKnspg5ME
4YTOGqIn+hHsJUTJGbaq5H1dmhEodtCEvAW9HkYEnLJ+EChNQI1jTwevJ1IJE9x8
98hsfFYw16ZzQDzsb25oHcO+HyhIZiaXhIEL17odQZG6k94qLZK93KFcBYdYf1J2
goMHWPLdBC5/qUxHcPuphtHNwgEmEIbp8Ou4vs3aOD+paXTgRAw+ckLB2LnQXtwe
+me409ombKt4AU1IPJdqCEuqQuimWphO7pqOtueEeOUkGWJLE+bJAfmTLD8JAJY5
H31ZeMzbQV7ZjwbqSOAczNjHnpQg0aBHhxqcsruhaWlA8qib0BsIm9ENJHOAsUPQ
R0fBRfgay1cTP8eSbnBGLuWcSO+cbstPukDsA0g0zTUl7R2cjDdipPUTtZ9APHyi
xKCPxuq+bQHfa6JaSmM01SyHM0KrXB1Bo3OeX/HDtx70gQNigYR795ksyK7uuGyM
TIw4i4g7L8WSHPM4QZ+p0ZEITswj9yK78G1ciLU0RgGapkprjntnJkIf4wSLQfzl
C09XARh2szDP8bz8Glq8JK+MRGrlHfLHIqlzFuHlwoxtjGTBj1dcqmTrU03m/ZEb
f+3nFNlV+ET9oyZgCaMDOE6+RUE/0x13eJw8/9G1vfSYCC2AnOyxLrRcMl25aU4z
9uDQOhtqgkFSBGLeSxy3Z8bSYXDwOdGZ1fVJ2PEHLCZjS7SmWIXcM5qkcnzLbdIG
yz4VW6eQua/+zwtnycB8iQWRdcKs9fae05W+kmEqaQl2dq3i1/mRB0vHUrMfUUj8
KwQS4TM6PsBzQwuZeibVJa8St5IctiuNSSO07P/WbSX1HR+4heM87/DutSUtJ7Ln
1qx0/+gFAHvAz74nx3iiRusA4iG4GBZv1KX3JnSuZ50cBVpYSwSDvMpEctWFL4cF
2GbR7cPfemv3wo2TXX10KhKcmBFizokl507Z7g7cUCdNozgk9e/2A1qD8iBuas/3
ZFEEe3MPuMTPvTJThgcorVkLkliMw5rHDdYkV+KIfrCVUY/XhSZBV6ibI5rHaKLa
G5wFHrxeP8CRkHTCR1sAIUdBdXVLqAr8+vKo1FixlSiCASM9JKLaBGYu/D52yg+G
I5In/dgHA+oRtgkGBQUIzGXYIwybii+X1kc1KN2ZyyUOHiBKM8pv2Lwxam2Fn7OL
gjSC3Y+si8YbR6XCgsmI1UmDqlnZ0VxzjJAh3V8a1T4nA5o3K0pgMdXocrAQldlm
XTY8re0npsbM18fyleq/O6OH3VUTWz6e09I031tTaMJn9mj89+fZrzS7CoJVRlig
j74w9CopBPQ2XMsKlfqs5irji/jXEq7XyoTHuNOfrBOyOalCaH8p7Zri75h5LgtK
mN3Rabj2qo5dE1osrzB2jGHnMl9YSVnArtSa3DbucNTZxdTp4cE2rwY/7oByqzD/
Fn5rHd+JEKW2E6Wdi3LcZQqYgSA0zBejDxVr8FOlo2woDNYkS8NUuJ74Vb44lWbY
veAc9idDLobR+pwHuQ3lNjyqqz078+DiHgTfhQSZvqKUhn/scC7IjNmypfX8wlvR
mU3WXv3GPvXH7MhNHU6LzcMisKoUcPuGYwL51iHoS9uUQa+EjSobQmPQREVieR09
kbLxcch4AIHTib9IK6nm5Q==
//pragma protect end_data_block
//pragma protect digest_block
rOIOgpjOpSQNkMGFm6w2pxsdvlU=
//pragma protect end_digest_block
//pragma protect end_protected
