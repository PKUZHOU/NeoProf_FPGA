// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
iW6kmMWouiARWc727OIbY4ZjAQZtik5mH1yUs1xAiZa18g/Q0mctDtcHslIkpTmA
MUpMjO+tD1McLoRFchlHCJUlewEf2ibeKQd8Ns0PtRHKYVmGg5xtq2i0g+2iE0Zx
XGqFn+hJMz+fMx+DPwcLurKBpHsqsJLVnVBveFR6CsI=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 28640 )
`pragma protect data_block
2wQXC/u+lZOXnnjeB5Y0o7579knS5a3mcRUe89bstxuaEy7Xr6CesXDzA04F6y0a
jRbYDHZJw2B3YHOHdUXcnc+99k12y20x7LwIntBjeYd2G40hE8WH/1JWHnTiskcA
1GVR72EeB2uZlpy8Dk6lWLkPfzneIJj+ej573bKPmw/mvYekBe2L8yWxW+LwZkOl
61Eucb+/QuIkR/N3+Ys0W0bAyjIz10ORf6Kz9Ozg+FtI44tg8jgv4BPp16mtWVAW
PXnstzQWhehQntKpGa1gBxucr2a2e4BC3GqWkLksalKoL87FS4nmD6PaH2ja7hzU
lH7ZB2d0z9OFpDLpsEnj5KEXxVSJFr/LzvFMERTZMNXlX8aEVG/FEXLR+6zsZQVj
EDnQXcEXChw9QJpUI094zTZaAMjTwEUIhKgVQBJkNh0uyd8EVpxQGzFo0T48+nqC
mTLuZHSGDw0Bos0EDN/b8vpNwY9IB1l9NKcuNuZxSy3rOXoBU4/xpjVfpAUZ7lDu
XHmvxJle3LX/KgQGY0CR/Ek1YsdHxNr9mW94CsjMw1KlXtp7UeLU+dWCPCInGxhy
+gX5bEc8VGZzLB9cQfR7ZuhfYJf9RTtFJ8QYfnasARMAuCSr5viobLCvUE7MVcmQ
Vu8zcFYcLhTT8G7WWLxjgce6dISo+nUcrJ+Sqoa9aVxXh0Qk0K2Njz98/WSa81T6
fz8zQsDegKV/REdVn372UHEgKKUJdenmpZRWJrELUw9S1/e7gYDaMT+8rU6Ndqsa
RqI1qa7KRFkq1UeU9+ckhkI9jh+GclCEq6XMWi1MLTsKjPpkaE2O4A8KuZTRWZUF
V7MiaJm8o5C/iF6jdJys440EFNPndsH2O7eNQCwNTiSx4lvNqKCnR71qhUOU8/Nf
WTkbr3b0mvGKuqUj+/9BjfWdbZm1wsuTT5WNRzh6AYfwCYgfluoYsrKcwovNe7Q6
EiHe/jsCuPPru4wS9iFCljU68x0o2DlMYaNTswqWyW2pd+7o9KGZiJR4FTjhHnd1
yhRe8moRkIdFazUty+M76X0vafZsZlKDkrEdD1QVOJrav+SCEuAyR6yYIdQH9P0o
divBMEdemQd82XCSG0iypSVYpwFTZgP9cQZKY5nfBA3QJ5cdokTpkPfIfNv3qr8k
Cwbgg7L2C+z9OrDRvh/2HFZ24A7zj9ReSh7Uk6n2U1SlysbDIPunAaYS591WPVUJ
cmdl18YfLJ5qGmKRxbYFELSGAxqOMUzEGptsgqLxaR1dIMAtdobX7Bp9gIRMwK3a
L1Wx2PonnbcWwhF8eCqlba63Hv/d54UwY+1SvC9GNczbuUEomifLf5Eax8aW6YVH
DC5GF8xrJHi29NXia03DIFCRWHru1xp2+nSR7c9HqZtZbwHOS0NLQQpv4RzNE/D7
FJqb0o2LJ2cgAcz2zyEc+inLVseEbwvZxQzbfEjt4Z1dD5lDioTlxJPQ968EqxES
H/F2dLnQO/iz08S4iWqLPYmZa/PZIgiHNWnw26NdF9JQ6LDTlvSw4D5sagQXexRT
ADTCbeFKaKbPuLfm2eNBjerr7my0OoxXoutOxMw/o8cv/SO4iXoDCB1fr9JsvILA
jah+kaFEHocuIUXVTe2rzp/nm1M1MVWC4qqhg7cgxkkbMA/h0SFmK80TH6hqWkmE
f57MJYJ/s365gIUoLgR/gcfvgesp4TJnDpc5bkCerkkpCn/yL1XqkfzcYbUxv3YL
btXR+17uyRqcosGM9Ag9wkhw93FbmsIEt1pWtiDYTGe745ziSyIAQcOFBoAuHor+
Ge9GIWbDl8FCZOg92mk5+EB0pfDJfU4hlJdoCCUWkVtQ+y0qxxGoYUyq5LceXRaQ
Wu4caTrMie+gw2StlE1L+Ie1aRthZCroQ+PTS+flSLBIYl8tEGshLhXmV4g8dhD4
bIRvL/sz3np+s4Kw/qoAtycJ/t5VFHZCllZBs3xoXoXUf2ArPctty4C1GsUdVvsi
LtKkC+MvdZPhxgWSfKWZ174S/qJW8e5FWoG9Xjm9icHzWePK7SCGNhLEakivpKcB
qJmOqq1fW5RXCu5kLYd6v93dtfGSoRH6WlBxTY91OZEIaQS0DaLN3se4mMhXG8Ko
9qCvI7u0KaHvi3XVy97FKafr5d3PbrgMlPqpk45c8WIyoj9KsCYgZKG/zbyO4fCa
TnuMkqkX+VxOkrVSREfu9x9sd6LQt6BLAQR/rOlVB9WdDDyOI3EmGF3UNjfbObXO
auEIO7XSOAh5L69SHCGsX41L53tqb7aogFP+4V+eRIoHSlYnO2C1tmfmJhH/jsR1
nBYMiZcXIMJhEK61d/Uk+k1hv6d9HMCeDvzFjMjdOHepufUxnoX2lzfT5K4SnMrp
4qZo4Im4lLlzZLI014oYGEXqyLCoUva8yKHilvKo6ci+r5/WSPdV131Gg853EM1z
fcB5MjoBf3A2Uo55GM0lv0jMYPCBZvoy+7pNzvaYJKQrRFe0SIZLGwT4HaKVP1sa
Y2ItGFh5XP9tSSsMxahUevPvYl8WYhLpZ4gwd3AYa5ksbsKoDLH8UoGEGnmJirtT
58NLnzkXyvQi5lehfwJb+jhgwaSf+u/h8AMqYW4QXz/lUPqPvcXnxKD03vhytTeA
UAghCN25AD9woAZep+9+k9X4vpTkHcLcdyNScwC+mv6IuwAtX+H4MdV7x0wofey8
+nVAaO7qQD925BPqAJs3OiPVbVv0LxM7iXcEOpfcx+biCXZm/WNRQBtffycLF/k7
uZKpuedA/lUS97kqxRAXY0HBrNAb3+KNgBH8YkBSmO7H0p7AN+oEY8lqMRsLXXEy
ga/TfMIn2q+B/QClRpeh8V/1om/dTHVjTY8etDw/DTI7EBdTbsmLNeQkkMp3enWe
Qyat2ekj/IdPnLb33TgXpZuSWjYdHKXuxdwABjJWnGQmn7dd65t+ci/3MPpiK2IA
SgNyhoFbjlVqI4nKBqYC5/9tHmtbFDNWo9uzJ3ElnjErWJ6FDepZY2+/22ouClUJ
ygD3pVJU99PeUdHWjBWC8PV//1rhDjUdl/6e/cHLYQcpTk3ZdlAxprnNi+Iell3r
P/IBjtGcfjUehwNImC9hvpLkuSCZ4MQ9nFyDUD7Xhiweqs9JWqs4KG+7Nmm7tirh
RqmpAk+otCCf6EgBDCmHnfpeM+LdDzyHb1kqVHhl+lIYSjn9ylvOPG6jc0HmP9Pq
JYt0e/Na0oSta4/pt505CuF6lDiD8IGUPCFfll97K+ZYGEb2skaa383rlXuUQ1JH
nJfuveUfE9c0FuFmvrZYPOaaoXBPbI7uoo1SvHPZj5mUp7T7fgLXPlnTH2ihCnR+
G6i8ItuRnFds8b2WJYyTls3UvdWx4I3jePDKYeldGlh7sU+XXsz4J0fetVoqpAWx
4RVWwC/Ms08JBrX26pAVclqS36pzJBSgr4X6phNOcqwqypu0/vNiBOaVJlp5jqXf
wDynjXD95c3fx3pajsYPNx1XUC+Gh0IOD9uSspCaJoTMCW4mgEIxLKJW+P25edYz
Cqg5yaB/lx175txTqN9AD/5TlKiOw/e+7ljKoKrrNnxSEa4eUNeuAs4JDeOs8H/Q
hMle+X1r2VvDeYDRZgveVAXXEFytMX+5L/G+tnvwE06hGLGdvPOkZxz2Wb65Aa4B
BP6mvUn5vdBS5CvlwZPItNUaLUkpIGkx4qc1XaghxIbi7v9w+ezx6g03H+gCupvC
Dpxv2xhy6iH+S8EI9clmebdxh8AXwgrChVEWzjqic1rTzDFICm/vKwqXqTASdvgn
C1WPvap2gz6S46ltbMmBF/+SUlgDGdEBbmznA6mBn3Cd8jw4hih2tyqihLg2HfYB
TEaz+81Hk1/4u7BaokA93jsgCie1zGh2n5K5wZyA6GYWHOw9dMRdKNqPPLzblX/G
MlIqmHwqLsKAEM2wN7DpvO4GuMQ4PCyAtPAwtmSnwhSSoo5/ZRIQFs+UU0FjVnpI
X/QBMjGXpfXY3bnI+aHMZXkzCbTMq5olHnUOhgQDELCUMRV3WrlR1CiLVy8QOUYP
BDs8W2e5UMK1pEeqqh2s+4p8Vw+EcncnNIjLFbQMgzwQsY1WW1y+eIIKulAbX63Z
l3M1Nm76f3dI4KKyxfruxfs1ZMJM/X+A5Hb8wdnFicaCe8L1VxZEekOEVo07yDo5
WSlUfWTnse0qy7rITHVbWUDVaGCFAf1vWJkn2uyrDEmMHiWfz+j3QuZQCM4XZpgy
+EvDGYWL7dGlx9ACLDJlvaqcYnOouuM3q1842lz8QobQEPuy8M1OSptyKQdzqG4O
4K5cANM4BaqMPVBuesUaxXckZ0CCsrCrMXDq5Ohmc1n/2jGdBFpmxIzbbakR8QwC
FhACzMYeeBSuY7fIR0stxwg5BiymebO40e6uvxtUsdx2o6r7JgPJ0e3Oz3ZwQICi
LOdmmBIXXQV3l7FZNWp7F3y0/NmQGKQE2IOImpUSGRxP3LLYrKVuxLvziAImIHVe
LhOyp/BCClhniIoHUvD5sLM2CCaqwTH/T6O71RMollXHEBgtjzGElY2t/wWy17JM
FXGxqWtjybWOGfgKCh1e+wkNd8+JHBR/004fKNr0KcBYAI/vf44yk5LSUjxjFrKn
ycjAwf5vJEEHwaf9qN5/hQEZ1EfInVWxS+oLFOyib803zyyPHpKM0i7ebpfBVZYC
A7Ex/8tyaGnn7pyntOzsH/mhKQicCfHIXadzfrFx/hb3qI7az3AqXYPAxGm8bQN9
OQPWb56IOw2Z0QVEE/Rf+zGeZbAnUd/dtuYP13Y0WatoopQt6e4neRtfF2Q2/5X0
oYLPlgRKw2DshwLSk+SQGU8xuC6QSRGKJSe90wd64zTAdJlRhDPrbILnBXESD2cH
7qnj5PlWBslu78c8tRhyQFQ6zx1/hCYRfRbVCO6605iTtsUknbfKk2RprZr8/SMq
oeJgAr2t9/ZPM2CBpb4Bsm7ghljECup2DG2jEr/bAdqz0GhVNei2DAfmQR/8sqKF
kFE/KZZZnyxScwoVQ8hj62EtyCW46JwF2rUcBdAEPtagRx3xuJyguyli4VM+vtW1
Iw3TRPUfOwfCdjpepD7G7OgbrbsSHmW9vt+yP5e36PMjG/4rg5MNdGtISlNJtc7T
8N87BWwnlJU3V21PS8PbRQyv+5CeCRz0Sub+OgnWxMGj0StLKtGjUJIZwm45iW4z
YTlzdGRDKIKS6ZmRRIVq9LMyNgzZ9f/WN3yKrZsgw9vSI0sBkrZ3r6s/pSxKT7Bw
QvkQ4n4kz/fqTC9wPz+LmTPrsbT1saaRQJ00mf0euRNFdBYwbRGXhrDdYVt1l4pA
ccls+hXMVJt2eAo0QFrprTsTHkpkPRK49lYgWYv/2BDF1M4DSSHXJZtHVldifFp1
XMzAfuKsPHvSzSDJrdrvjaT3///yZqpmLbGhgW/uOu39+9Ynp9w+zFg1XX1/iO4m
6rIMBntekcW+JoLAzPLOdTqOMtQOK8k7rx7yV3cso82bMeGllx12qcQIFherC2cR
EPprWa8lsZDMjej7J6IBFRvBLO2mFFjcWl4dlVNIoCB3KJngvAOFMMLDPOopu/dJ
WnWnfHz3Ux0R46PqHUjiJrEOwV9kPB3C2mFZaDZYH/36H+hQMpdYvYHCIqIFGBer
7S7OH1Hf+qPuz5SLQiR2ohWpTOIjVfaCl/IhuZ3hKaiyQ9O8VNOKtLyI0VCHkdld
+C2CCeZ0NDrZKnG7aJHq0oIqr+Ym7+bdoGAwZSrIS2fq7uQX7nbsuvOnqt/fwLBT
Wwo2wiOh0YLhNOcUiORnPrOoppx/2t/t5SIsB7r01+j3RYd1F8tG4TZ9OzWdpIZa
UQYzDdhkmkTn8mxvPBcEIEZ//HnZ14brZBEQ5+B2G4qDo7FBztpQe0vjefrAN/xf
5dfeu7rD5r1pz4ifOI2Hlg63xdcKFcRYGsppl3PpjKUBJNLYZrhJHtkDvFWvSUfm
WzmisF6YQmF7dIA3XR316cMyTLcBg62iE2iqr+12vfyK0VbC6MRjr3Jy/bcpkCKK
nkpcihJpIrYqtr+U5t+rPmarTxOop6e367/eApdwc9ZjG/Plp2NS2+L2lMxh/vck
SFhOnoLk59AfSquyTPs51Oq238gdh5NrzjjDh83MSleIkPTdnpPjOoKwvu0zNH1r
dXj9GsLQbHfsr+2MR6A8KQ61k9wIpB7Ut3p7rLX1z8FrH6ptL67Deqn1PP/EARoy
y2wSKsPKvOd/GtVtBVg1cKGT+BPjOrjRpmqwMMVabWVdKvZUnMd5Om2jhk+oYr2s
n6E5aafz19V96ZvyjxyGWiWIFQeirK+v3alkwJJZSFe/6xeg4zFnEflpoe8f9YLS
veVbyyLxgoW8M5W46f17rAQE6vouvTjtIaDLXhF7LXgVa4PCg6O7tWqeq1s6m/CC
YJeVD6IkPkW/80N2P3iV0+YHGA8ej44tfoKOdHIvmBm/NmAgPe47KN5FDuq7rB/a
7AZY/Q0S9IeK+E5D+u6GP2MT5f9y5WcAmcohtv9CdxHaaoukJn4r1eCGuEUs0e7o
QA3rYdjDNNNluejDTao50WyGB0CFGqBlD0CG/J0PuKLRAr7fTh13crFHfSwg2l1r
4Bv6Vz7jv+gt/qrgiPk00iWn96N9kedeWQYYbKnoCQMdHCHm3no0d/8UfdUtQFs/
gytxLTyw35XsWlejCPvGPYOE5WHWoYeZgD7USlv5gkXs8m1seIgbU+WBHakpcMCs
sfx/qbKdrcv+s8Lu1bt9BOPt4pH1yzXRlDS3toVDmtl5+KAKQJZFefOX7wLJuShv
+AtuWbrtgjS7Cmv8CFFXkYO17JWTV7C1JOsZhH3g59BYSxP59NTFjjXnvXivXX+6
dE/VSgx0bD7pnhPOGcN/0klAItSpy4IUEhKEb3FFsC81X0Ywz11KZv+nZf5GygZb
sb9I6XtyhqI+qwEXAO2wMYrH61tMUJZsoPhWPNXxs15MxdfzLiN3/s7CVEerrdt+
UnLcMGMxwMmqMIBY5SCl5xLm/glkotz3YnOWdg1WVGepmm13V/XXWjFfgmF2n/FU
eaZKH0QB0JQb8/xAgv7ySqsW4P1zbEbkfYzdfsIRYFlLevQ97hgeXhOeK7zK3pla
ovGwlL9YcMRciqZ1B9OoI/HxGZ0EVfFK+v96xjFU7zNuJ0EWFf7HsAAD5r+kbUdS
HzCNWMiw6B91cdQKilX5TBBq/auhycIDLwNqHOK5aZFroHq1ln258TXkrUOatBDN
j5sInyznpHiG6eZ3dGDsk0gQOuojx9c6Ta2hqGoQjkg81ML93aNE7Wyq/78Kmflf
l5DV/GdTb+rOm7NUrm0eV3wUpsOqjeeMTfI+zN9p7eYgh3YjmqEuDjVgQLRC1BNc
D8CqbrDjVQS4nKLQKUWTuJR0WyC+zL85lkrQTy5Wvin4GWQiwsds5J8beh1ChFqH
xZqvTGEu0Hgc0SsPJcmJJ20zUhCz1DBQuDouXA+y+5Ka6klGMaUkrAEwI29vLmNY
YGyqeaMq82kkSCOwxPwjRW7BjiY1nUQTSuYuJFa+KkIqG8D5VAMDhdAvR1Fsilob
plHxTWbh0XMaT7Q1Jh/XMU4qGmkcBvsP7NHMqdkp92cXh36JAzs7mCAjuddM4GJ7
jRzsNXHT6l+lzCy4iGwnijt6vyC1qgTsGyYhRU8md7+JOyY/jaT8o+iaRzlhvAEP
HBLpk2yC1gRCU8gHZ3IMdoV7bHKgwh1lzHIlzHvdMLHO8AV7XjADYJeLvUFE2z7v
H8FgBSw31Tu7RpkBdzUldJiORisy0VO1urapeTMihhpdZW/luUJGW2RSPnhUpZi/
wKLZi7jtDNuthQ58DoHjqVSbQPLwWtgszEf2km3Nl2sI1bVMEcgJmT0z3Av9kgxK
36EP6n303UqX9q0qVOxE9r0KadlTfYhQPrRSboRNK7dE5Yq3ZtL0aUMmJmwJXEM6
Ql23TYL8KMgjvjnJRZJlzg8HzZFwPwofDxXoD5jnuZlROu60ntjKEbOGp7yRqe7u
fX9ohBBoyaLndqivNCe2aeYa9s1Q4mxg8TS/RgLU060D3MbR5+j6rO2nphOUveHE
bAbDaA2BlrREHe2o7ioU7/bLYiXsduXwUpAPMqrIrzgh/6aLs2kz546B8khWWAnM
wi5rKqHRXhZw3Bwf2ag6LU4dxOYzkzYiKq7UzA14BXwlxtT8IyD5mm3vZaL6naZ5
52gQ5A/EsnpN6gHbi2GzUqxylewb51DC4MCqT5Afy/ZlLcKkAEqHZM70cNfVgKuj
eWbkvvpL4XEgn3GObh2Tt2loewCMYRdyvHmvSTYRd77kC6eGsMaXZ46furxAQX71
MMF2K2OcJ0shP1W0B5e8kQaRvdaj/OnQMUGi5MYVwjFe7ilFNuv7SOl6DI1LX1kS
RFDHiNbwYyt1NnrRP46YK4QFxuZPUxie9OTFue4vww6s0kS5ydMmQbgqdxWFZYHb
ukNlK+WbBaqrjsEW5F51IGxs17m1fr6FOMc5FGBU6P6t7KlG5Hl0DWyzYKOFaGqw
HJGw0IvNKZmduoXiDQRZxM0zpawLIm2xG4ZgLXxcd+v8s/D+rHUP8b3eMwgvksM/
hX1a9FT03ag8eppA5sOv8OXwNtecnB7ODiDiIyVl3hY5ZCksWFO21A5lytAhape0
ubCkbGnNQak0KWPBG8ie92scIYJaTLfyTEhbOZvYW2raKSy7Gs0YO09MBZsdm09c
1kgvaUuACC7yG1aN/TA5ukge2Cdc+7oGa599fkiGdD+CQv+g4Glop4Vtbubd7lff
ZYb71nC+cGoM+20RHfFSVRY7t01wma3ZDzl83zhHMjc6tapftUINeburY7PidUNV
ZzvWZSGXZ38pocJSdtlNJGBvn3vOFqTQK3M+GW+AzKG9PpKF/6KnWiXu98YIl9Af
KXErCanFobvZSUxL8uaJTOMwcsppOn/Opo8DqmDPIEeQK8ncyQxQNIF6MZBnzyLN
5XWO4G15ivR/KIuI3Y1nz2rHRAh9g89JgqPsSiKGdMOMvjBbyrpGx3ogITED1xqQ
kxi1WZK4MxRO9ZWkvKoeLAFELAaFwxZRSV9Cv/Yw6tlG2VXJUqYrdp6kCmJLkqsf
a2L50j6PU6qksdi0NtTTMh95CuITAlrf+WctMZUqYLmsSJXrH7EX8YQUqyE64z3f
XRwSeMbFFuAySxViosTpYkz+i6NmrVuYx4BDa5LjwPqwnsTzLFHC4aA4kCCoEkDL
D3iCtG4Ir5rxDiZxkGvdDO+f+o+KqgfRo0zBHoO7Z8VS0GmFhpMakBSoFBXhtz6f
RcLPXlu7VSpZeHZk+UIvuLKMYRQosGUaY90FWlq3yAHA3AMENl3VFGT7H9xsaois
WIZ4rSSJNx27m9r671bVS6L5j1Kz+4dsfrqCbpFIXKAMkZzSYjOEN4OV0yKr/YUc
pBtVmsKGwmzFMjKvb2HbL8FX5G2ujvsu7DkN4Xhl/eBnIng/dKHshFZO4l19HmlE
m+Lee0qBXmM2GtTwKTJQqbp/zm5EslIVrPnGWv8R5LBLH2B8tzyJ/SaeGnim0M8h
oqFHakD9eoD2VfOcJkg0AgsyzQZogm000PMVuj647qBEwzENvh7Qfa67e/iKEHdW
KZ7vQxkCRRKN9R85UAwuRrOYNa+Z5uvMP2K2a1UnvmKgQbv5V3M6X0EP1YkmlU1Q
o6jCiHjMDNynH+jJjHTBAv7qAefTUwKRoxW3y7gz/Bqf5FXobDB7ndDPUIxO8lG+
2BCkGas51Bvg4yUBjBSXawti1zL3/MEEgQUpvG2UU5pRf8XHqdEGwkC2YJim7fae
loK4yvxlcKAK3g5x21OZIenUupHgquLKMcNXJ9WgqmUuy2QJP8yunSyO7Lwf6NZL
JC6ScZ7zeP7k5OkPpaTQ3WxbFDgJjKtG/j5Lk97PAEgh6br5S/HQac0EFTKIb1X+
081wjoHRPKDOphZVlOWaCp5Yu0zbt53TpbBq8Y5zG+Erz72NaBqT/OsEZx3eRhR2
g3I5ybFXdeZYyRwfJ1VfqHweBab/xxBsVnJWQJa30GgPlF26QPZOQZCxou501Llp
+IaVZv5poogztBYviLkQAuR1XZ3wRCaa8Hr36W/arqXSyn2XTM4RpnY0MdYuu1Kc
NtTB+gUhL52T+a/YMXkgWQ7Qq/2AnrN4rHgk9RzmKv8Sr61qN5mWPv4FVMSYpLIy
gnY+MUqKTVLDeUpziuBgfVOVTTpGtaUV4QTCfr/0HruIpXF8vW6qOzs9yo/EuRp8
0g09ZivX+63JJAvwiSfrZoZjFr51ox1eqA0kU/fUeBgJya8KOEhRRZuGALKXZUiw
m1JnUQd4RLbSkcQulN0aP8BKkaGG4sBCEtQuUJjEDrXqYxcXFdAxPb8JE3XrfvZ9
Af0ZK67P1ENF2BLTqrxHCEqbOChd6AY+KfFUCKQRB5PQm6x2T0To8LWIbiyRsJA0
Iqszso4nH7wylxSY+somwPtxIXTNnrsEO08d9KlxkBRYvMO+7HCEssHSgps7FHly
E5wTG8F5Ro6lHx3hvJCMAKNKrel8cP/umePARncqT3jmetG6FJcoH8jZ8Log75qv
5wV56fNXuE+fXiM0sGXiY11hb5+bHRPy8/jpzj/DnBbyiF/Lpi/NCjwNSQYTlKDC
hIbgwOZIaGjYkAmLi0vaZE7t9yRXEMI5MN1WVw8lHY9MpTwmdD4mbBaj4sn5T2Mx
f62azIgrWxke+719DgOtDzOsZ+13llPCHzQkVV3JE7nNXT+IFTLuwE9e95rUidII
BJXvx0NmxW2K56e2aGvYhJYpydsqHY2KQyCIpcEzcOJukvh7wAtCCCyJ/kG75C1N
bpAiJn9XNCOM6U72CxaFkUsLbNX+11f8TOLRsKrDN3S9JgVj5xOosewCmLoNCoK1
mbQmmXGzI6nbhGoG7uosIODltKXXBqY9MtunOPDI2A9MwrTDUAZu62ZBRpEmbcjh
2XFik3jvbnorwID0aMJ1V4YAC+zpHFGdJLDbc1+a2GBOFj1njYEXcgSbjWlSrXJe
Z7/MUSKTxAbg6Zy7qSsyvtaeV075fuTdHOwAvo1cVqxLkmmRUHCW5zqoOuWL8/Uz
vhgL2G7GogOgz7HmyQJ2FvlHvGryHSFGdTU4SWQlz3rQtEdKxVyI8S1HjIlIKCqR
wshRfSiLP+aQa9gvn7Rh2WQHXOlx5EpfRqtFbfSM4oKwvA87ltjHPIpv70OUx/1/
iDIubZ23pbLHQ1cpyxSC487jmF6fgnpslhVqG4Ot/miI4KFh+XhwsFmSgVjy/meH
9zD1kdU5zxlbtHJuNlQLayKRV9WJeP0/rvDwAX9m0GUdVcdBF9lRZglCcT97KP4c
BbBJKz8wOe7achnKWKFd4SosZf7N285jqdMRedoAd4i4CAES4E9CaeCPYsr0b+FG
bCw8yzZZnKOkN8XCB4Tm04JavzfTMItWBoAUFBPuYi5Li3sjpp3rZAzwgc7ceup1
OvNuEmVvwcSSCQSiQDoOc6uqzKsFg02oDJfn30699BToue6PI1xunN/BGVVrOV/r
NoP5uoq+vrhPD4DTiIU2DtGcwmIRGfOSDALGNSbUMIZPsaU3f2Pv0ZAKLuPI0z/k
CAcJMRdujH1vGEs7GG3PGfo62lmY+n4Gg1aZuRxPyH4dM7tSlrdP31eJxR5hjqlP
wnvjtVvvwTkEA8+OJSKvN2EpbXA2XL1h4zBEZ2K+Fkb3Eukp5cF1sXtIlh4l+Ltt
l0HgC/eC14npdjFA2HB7Hvgf+4ShgrjMVSFJ6IotbELjRSZFGxNv6zpojXrLpiSA
QeiwieKLEtaqdWEV/z6OK/NkGO1y1gaVROvtUQJPHLP3ZTkZAVtcqv8xBBj/AFtx
BGFf2pG1X+ZMRqoekjfwiVvYYO/bgj15qC9N57gARVXRaUapXRsBFfqNzL1kepSh
PMuB+iOKl6rPJs6G1CAdHg5V0sVm0pxn+EToURimqzEZq0NmqfDGhbQDQOD8NsaS
l0WnlzWYFr8Jxx2YQrgvnRVhSgyguks4ufYZ6nPiF4jLDMMM3WDF1Yy4WVPrK78c
aU3mhpCN1NOBuKL5bIvGDXqnJkBti1ID/LrcvhFZoeelYUIQ7TYZNNSU8t6KIcBg
VxDh+qUpIhdFXGXer2TI5RgEkIoWK2SDuAQyNKrGrS0RSX1gKph1c/7qObm4JX5j
oH8SlYRhv2YoRkS1H44CA+/SL9OxfrDvNQ3ks4gei7BnJPpubfyZOMnibQcUIMUf
wiCEsUPxuN/8xDfTxY+JxzuUPejB9BSw9iWyPeArfHgYIGubXrkXfHoqcCu/IH5s
bpCe/bPXUS21GoHjVhuFxrYyl7T2INMvV2IInAUF1qihQdBKVMApSUJEnaXaxrAq
mL4FOM6LifxXvxfIfJHbKvRsiNN/vM1JTANZIKRGu1cmekL5tvqJOxajVgyZmUlV
0pK22lKjDF1JTcx8FLxcrdKRW+yQnkhILEU+RQYHBA3KyXENvxa+/rnI5bolgtwM
JT4BH6l47Nw2t8QGxISPMmkDBOVv2VRNOMkg3ZGj3fzhFGEx/XvVR0Y8yffu4P3t
LA/fhyo5HdMvlu8KbULnSXqNk6JDRzjl6Zspz8yKs+sRab3dQGi70HLfM0TwgZye
am0gLlQcpF7Av/u+3jD26P5GcVRZYkynhl2tzJV2zhvt/sLYDV+2fNLSdaTMzVky
9knhVk/YvhJ4vbeW9pXCl3pJ4P8Fsbd1yTzuqIPDQTl7BT5NTaysikXd9hFQOj6u
C1Whlazv7QnkSOzdyLlBliNSO2x6pxhd5agjFd/aBwQtqIG0xa1fpTnGxmQU9DKv
cOIHIV9KO6GYPRrpRKAmsoMZIfmtVfCrX89wpTHZaFQn2gxHiLJg9KWR5YuSa7Ff
i+7rqC6h4Uoqx2vCZPS3tQ92E9mQBcAfxKzT8wGvdB7uk55tv6ZQFsfdRkI37iZH
9O02u/WJhpjH547ohljlqyyYkOWzWGh63ibzP9lYUe0JzgNnvM+LHgQdSBWoNM3a
3Vawso3Yx3xxd00EmVQCFi2YrXzlw1PUv2yDE6Uo/oHPVZ7HDbv6R8Ew0kyC88AB
lzyGwE19izd75h6cIx4FrGiAxZH9EXhpaJExJhO+YsFk5APw+kOQ0EJweapUDAJO
kw6tpyB9blPKRjqFfagV4CureTLGxvzayVn2zmUDh+fQVBfvFyl37Chg1luNOyJN
gNpu22Vnd3MhNr7uMojdkK8YM7aewd0NwkZhOlge+bX6UOEtDIqvXHr3dLtEV31s
CWMGHoIspmTSgeISqEV1V5lS+bZR7jP6aKGfzx8Y6dNE7FOHRU4nV/fPr1vyW64O
lXCWT4LVaDE5vPiaV8sD521B6N/hHEn8WqFho/dliyg9DqNvSpHbsba/E6cCOqgf
+IY1Ght+cWCKqk6LcD5hbTNYMK9IeMoACn6ukMSHv9y53GyCVKmZ56oG4eQjlcmg
If/b/RsxW1UVg6E7zUltfUku9wdVQrGXerKaTiaa0/pyBHn/O1lnihCqdwABwKMF
mYiI3TXVCA635jXkXTXitHNJ9xVLbhmE2hbvrQPmp4rMJBDwu5c+l/0GZEZbdcQO
qUhtfCWUUQ4JOYuK685z9cDr9T/mTCLUdXe6g9fWv+4j90+3e+pq7TVGlWUi7y0v
R7cATdkeLOLJwlW2WREhhfmnL69n/WLMHlTZG9yjjs++D+lrkqE2IotNh8B9hBbz
EZmKLa6cmCiao/+g3VyoNamBjPYEnqLwMEONnYIYz8vlIJBtuWY6MLI+xSMhu8ME
7UqoDcKxOCubrVY/TOXVx32jiKOHxqhlaxSQdbE+tjrz8ueZRk8RdeQ8JSdpGu05
aD0kFDLJcxCa7Kz6CwJEdWHg/ZPgsEPY64LPFvgclWNzum5DdMk1uZF82UiV2zhZ
Xmlpw2R5sFkajdYNklwM61hoagaKDL35+O2dd3jK4CpP5Z6o98cpI699rzkJRiG0
1PPf2lBdVdG4PG/edXX1MCe9OrwFexGTXJiQpLfZKrqXyOYInNtLEn4Phy71ebNV
gkM7RV9+oBEqdKhJKbnrPvXkqnJAZaJpHcAQPzRmTePykNK5nzHMtJIyW101NyC/
8CMJ44uJJBd+2++VAaLZOoj4mDEm+JbokhU6zqpPcVCm6UHAs+nkohuzTWrc13kP
jwvceJu4+sfDFDyFM5Yh/O4dCTrFBbhyuUa+h8nS92WWXNl1Gh0iZS9h62kf0LEL
Nq71krxiiE4OEHYTNK7J8ticmocW5887QPCAW8CaTtrnkNPXZ5+3dNxrN7f95DrN
M48bbyKoL4JU1R3ysnrMkhigKl5EYutbNYUW8gNSpJBaPsJQplzmMONVDrJ+kJIa
NCdzqiJgxequim88amQ/I46tyxmvHlbbjzMRbzTGZwen6sb9V/H+0TfMBnmBLsYf
3kqNn1qNP+Sg/BIRwbNEZSWGTSgotobGHkCTaizR25vmIzGjSDYhqxpsbQ/QLiOE
oplcBoAR3YJT8idH75fmYwVJAczAzQ5Ft8oLQ0vOrme95AyBitYCD1d7BbR9WyiR
59YHzo/TEUGKhaeYcvq7ZoAWiey1b0I/0FUjpHzBRaSTxe67nrZpkFAG7n0T8Xtb
iojjpxnJBVitSlKZM7MT2F6pailAk1Dp3GY1JcdZmPE6lZoCXkQbZSi4z3mZFdkY
PZjyHGajrRDh4xnTxrkHfMsRidxMZ/q/39hn5hKu9ycP14FqZMq15QS/BI+H4QqR
+ZLUbthlaGKc0rFDOJV8ORd+XD+1SKMMRmPSmYEgXybCAA5J5hbPlWZTZ7shPtdB
Vk1g56Dke4UNCSc7L7SGV3xH1FjrJ8tRXuz6aux6eXB27/QcoFmvGtNSIbVwdvFs
jpUbRQmGZKB7IPJ+Ke/yOXfrI2HtrkIsjdJqqFTInAxGpoMQ5JSvJxIzaJn0mwxy
8pSCS/wp7nyctbU3WcPHDMvhpKtmv+7pflW2joa47aMHqWxTsMVWSNoaalKdzO5c
15UGZvuApSK0zyMaTEOxCwxxwqC8ulI+uu6ZcMiF3gqpjB7gWHRNKJ2PGoo+Xrij
krV2svFm3TwBOB4vuPgtoW6wS7YW0tSQ+VbdUpaeNIO+IN/p7cL94zdwwJe6QxLB
h5D18xqt5TrfiLOR9GNo3SyxShvKsC6TY8/2YIMv/sTi2KOnLYfk3AP0aO9qRHqt
ZCdg7W76BGsqawixnEHGo4TliheeJYHNTR8RnOzLoE5URlUdAjthODmogMEpLLkz
2T40p1o7RTmcM1ACkBEDuF5EiNMEVlZ/BXGyX0sEyb+8zQLUEgx88xQVJJPMYADr
38zBVXhZGO4fPd0i/HRsFtIR69cTpwEGXDxJ3lvWxk1zB+R7PFSVD3dbHtMXFfQF
kTKhaKOHKZuLEMKk+x2xBNfzR1wZzMEjO4wGtppOJmea3R9tKmEJA//7jrRUKNQa
fJCEbdfZdaqbVcm2yfmf5uW0inZ4EcozSbiXP/CW/eoL6XDNDg23hz+dstcJ9ZFz
TgQuUsmkJ4SdDvXITf8jATgXYuM2OLEhu7+uQ01tMOj0RUK8qAaUPbVmn3Pe8Y1Q
ihtV5GSJQ1HDceO53lyse7yrLfeZtUSaGOzck8W7zSbP3d/E+x8J4a87gKO/VMcm
vpizLpQAeSrmsoaHeJj5JyqSda46rw+IoCbfQbePLe/2Lfqzlq7oHUtDePyByvza
HilAlcS/tW04EQ6YgYzfJ8YoyOXNHV/X4ToLFhvxSI1HZboBsP9XHpunun50uDDp
Xj2qCU3IV1mtmVRf+/6KSA0yK9fTmDeDXvwf45zBMkkZShLX+NHFZX7Np6pTBf78
Zq+GjCJY/u1uA/Z1hflWiqcF62HB+pZugZFmfxJQfmUfs4dacvDTsYIN72fxQXWe
2wePhLpDCZjoFDIHHXx6dpKegUjZl4U2SifjZei+ISClkEtyX9iU45W++Yp5++Ag
BgVR4wvgJKkjjOvbpa402fyTunCNZQ2vjJNQ+py3QSi6Tkk6ewrjI6qAxM+LXogf
t+SdK+CmYPtpHKohE9VO2aUFdQs6U2zqSvCQ/jqXkohNDt08CW+aOraRMm1VzkO4
fL/C5OXxAKzX+NF9Y7Q1tFHcShfd4j3MTIUe8f7gSUOho/d8kwjEoM5LY/DniT8v
3gXn0yKeDMblVv3zfv+mbMicEwOGjZWWCCVW2ZUhCi057iWqkG6UMIFulCLmeIdD
agflGK1Zs3QMJ6RrdBmL3MeIfjFLPIGklPOmCVoDf24SigZVKtw+rrdSZNhlGMJ2
+JiQ6X27j8shIrTRLMW3e7stmtuCEFJ73R8p3CYFI670IGJorQdASHa5lk34JR3W
ZgtFI4lk8LxOYODDfAuP9T4XmTfPc6brg4ZOozWI4QIc10IN7T9FYh6agAZkKsLT
MjdBaZwmTtmTQxnx1iO4nX5CIvKNI6URyImz5+b/svpS5nRI++4giLsH8uqvrQ7i
otMZ/iezSCoGUpoJA9JLQbH/1J1DkFNkCP5M/iPP5HEE2eWIdThVHRGgTz6nqyLW
sWYxUbSTwoXmT7z/C+WkuFp/P+X+ioTMpC/vNBxIAI+VpcUq4YzLCVyI7vtOIUnx
vAbMjWERJx3VaRfNIJVdEmFSY4EYgKOmwdjGQRrOmC8oPNqlFWsUQj6krI8OMEI3
njaq1ILt1WGOy6N68oixXwzw5uUGlNGis9AdIeFgZYyRqqxwGIe7UBUxCTRJgx7b
2uWu8N53lLIIT66/AgKyYrQq6FbxR1hp5LPKJzQa+2q3UVC3dfrlGPc3seafKtO4
O50CLIuHQDlHEYG8byv+rVl2RlGyDxROmfYzyTL7TJBOo6F1QOLUciZuvfFUT7Sr
BL1DgLgCpz+n7E43AXB1C3DeTZQYS65ghcRTm5IW9+nme2aw7XlLumwweYId22NV
ZEz9Ivuq1JYKo6aOmLlryoBNnB4l/Jzn2wHm0i9HIoXzED//a0/REdCdefvttgxS
A1jSkSRylY/sFHfRg5ulIzOaYqat+swfXv8242EuyV4B5wtc4Gbpzm53qlCwfgL+
nv4Dp2DlHZKirgIRASryPWDqUBvZW4iVIM4K2KcCKQ2Gcu/GlvA47HkT7W7sJAS0
DaxS5ai0DUJgSzUyGbyaGMw7M/J41D8WWZS6LYlJuD5j9/Sec4N9QoB6Luzdp6gX
11rSgAvBLmbrm7WbMn/yIK9q7kEs2u1UIjIgmgKNOMEVZAlKtZXnLws04/pnZ8i4
NmBQMtDpGtmJXHYZq8RFZt8cuM/PvITdbNazFRfD6UYvBABn9/jEsrFUNkDIe77V
HvuhXwzrKiKFe9zsYsN7MY38kqzSj4uH1NpEAywO1+mXDriKcE8IaHkP4qJsmt8V
wHGFiF0PwiBilveNUBwuFn5osJCy1FrHG2NbdmZ8ySZtIZKgxMMbguBc2VcA8K+s
EZqjhipPugzpn8YBAtKvkA24a/Xo89yyWuZ0i92YoF/EYIi2L5jFF2ny8S9JkAoQ
N6bXE0C000tF0OAYxifFj7+DgLTXUGE5ej9SoRR+HRg8w0a2f7HvKYUmB97qF3tH
7O1mfyf/25EIUvdzWqL1zmikldy4go8Ae8J5ltPduy/P/bV6b+X1uzlfjNXcrbQw
BF9h3izGdJ1WtWM2vTF3/3JNz3lgrOR+SQqGZoaeyI20t7ZQCeoNR+wEFGYNT6zR
ywTbit5RP3OC0lp5b1QiJJotah1QTwObkJfYS/NyuUXwoX6+oSfzZKsJihbvykmT
MXRPcXHfEovRqPux89pd50KSVzCtKo8cvVgamZ/Sd0E0DPF+sRtpW1sY1lhbXW5e
LvYW/ASD+gBI/gCLgmB95rrZbMvZnXIK7a+SXNpfuQ4/VpJ7ncKbJCOAVHGXADYu
6LYnF1SrF/u1zhoAbPg7LY0Vv1e4gkKilHuOqnSOm3zHf3RBH24zmfbkjGlcG3IM
BDH/eX9d+ZDe9vNRsTLiuoe2AfVmP9EhnXnMadXN8NdMx9yOBE0Tqi1vFUMCIPj2
q5kCrhxtXwq/jH0MAEJGH5NcUod6HSngDdbe+2sgat4qo4gINyxaqoETU6+UC47O
AaVEVUrm/x8rlUVxgnsDKTp+XTP7jSl4495A1h+GhletcsNWB7OgdmtUXu2jH6Mw
ZO8vbfSInKHrCw8JnyGcfg7UwwMIEbyUm/wvPdacaToZyV7v15rMHrUssZRpfO/O
Iz0C/P/Jn9u+NgGWNtftysJyj+ElLRHQkqmFc3qxWPMZUj6c8VoobmZjaY3Bo80q
fcup5YpqTeHB4dhoH04WWL1Pe8FaMoOflpqKrZWFG5gSRgbb8K7b6d/laqhtYtuF
zZE1+wobsGtmV+NCfqtsMaPNmVr0jUV6JUtqD/eVfkA7ZTydLF5jckQXXiOZkKiO
82g6CoRsvcw+x5dWS+hz4aBmJMIQZeFDtVbR9ChDPNlENeJa24X8v5qkIZBlAZs0
D4qQszEGc2Wln/llRRFgcIW9IrRTaj13ax+nqUzjCiDa9lQn41axfoMjNGAd/Q3N
JngHGFuTAKzrq/NatHmpT2kMj7TcePcd0qd4YieyyQ0ZJCLKT2idDcVSfMCdHFwG
24gIdXog7wzZVJQY2V9o1/2vJ24PJunovpIQm0cGldzBV52YtkwAhhQHGAsEY9fR
9j2i6peTWGyWJcygG64H0WmL3XOTbAeynn0/7iCW+baTEg3usV/UInY5QrSKDrrB
80h01YD6nPkxW1XqzcZXbQGPbmuVdJDsuCORiVJPzDkyVVWLEhEtTOBYBtHtIpMV
iIW8019eVulFDKVMpX+ZhH+XUbWKhvjzuTmKkigkEZ1ZioHOmfiZMzZRSAGQenG1
LjEOQDhAccJCE9XeyvV3kk5z5MF2cOTaw4flrNbnktqxEuLbg7yjy9TPY21mrNYs
ecKu+zWmMDK1sbv4dpzZ7J/QzKANMMzBJA0YdxeIGBGi3QaKlbRbuqRp4oTPhuxX
JlN6WX5eALAYPsj1pdDUp/EAFKX1Nymx2g0Iu3VDK8XVKlCZdFs5rAsybpBWTW8l
UPHe7o1Er4mLHNuMGegkz0HvgdtkxiwPrjXeIJwia4OPp8f31tBzH1KkrpCYKrEF
G1ny/wWL7bcHfkA/0LC9i7BPF9ijfQUjPsr0+8OSJEbtfKTGtbpeIabNN7yUjmum
0TFOsI7eVE8oEeL7PkY93j6c8MpbbLK1yUMYeaC5lXZ+mEu21zaIk30gU2fk2h3r
eZ9YzTtNjr5nyuxltlPYDOen3P1U2KLsIMMe/uSZgb38Wr8wlsnVMPMV8PskWpaZ
YhAO/ZoZgu666rU0Ap8A3x+/GKHOuh5pQpinl2f6arc34zII4oNRCMaO6Fz+mufN
b//J8D3CojyuLJy2M2YwRzLpjfrgxSm+JrbCfLnez6KhF3iUNxdhBGFoIDwtfwo+
TPbqZi4lLEjgHRU0Dd+uheUIX86d8ReumQZjSiC3oRHn4hTruJm/K+vwSpTX3N0I
Fker9CPAnOIxA9XMInMgSqiDlesV6XAWl9EvAuTjf9+daXk4JwAKN/GlhQHHe51A
5IC7s9zL55BIR2mfvYTMMt/pIAVk38VuaJgzoGrBv5rT0rq+UjBcLT41nUUA8MfV
jwbnQpBOPpf2uLaE1nAD6LDwvwKcBa+hp6i6D64VVOjB+PIjYHnOO0zJiYDBKjc0
wjJpYIdg0nckrRc5lkkHm3Cc5aoInkG5iYkos5ywHeoEJUVTb/PrDnyIudG5hM7e
91sMGekGbe8CaR34wYPFtPDAyjPDb6tC+c25v/bCsRantSs5qLkAhU2uCqXE5ca9
ANAXx5jZYBeTWvoMXI5xsZokZ6XAHCMAtM8FygPftkwE6GS33mhWzd676b8ulUxo
tSUkbVuksngHoC4P4UPuUouixmQjLg+rZp3M65+WDHH+bZMYPT5B29EP2O3MwD13
eoD9GzPbCLRCrShPupJCgbKbMOKKSrSCyYZMTxHMtcY7Xu7V04W74OItWjOxNg1X
MDEbez2SU92+KqqykB5rP2cEQe0dwixfTek2vj+F5ol25vDpxQblpFFvmRjg0FCf
t6pmvJKgtn6yw4itvm/7UTIBlAk/asSzedaDr16Ql5eR6o/CkZQK89P4v0uJZi3k
whODq4ti171u5OMUpB3TFWRxX+I4BKLaAdW1B1kvYuJ3m+ou58NaNByB4/KDvlsm
5o2hsSjqx0v55wbPEmrNDfIm2z1gO+jdjmtnpIqGwlV8fQLa1YwpqgQfrMiB6idj
YfJl4/ifc8V+BKXnw9POgwW0+Ct+ixGqPsC3xJrrxFmzT/vlm+sIwnlD9VcI9o0+
5bxYt9dr+VKqAAniAqkRPIFQLgz+9MppiKlwHeS0hI/DPUMJKIixgdoHJMvhkf0K
nrqvdYb9gEu2P70l7lUh/I3CEtcO5me5faBbBd7nSPNAIXU5tmfRQVS8dlAxjT4I
LFP3+wpEvcqpy/nxYLOuHDrDpiN5FlPkB7ILTUXZAeGIuE+t9pea+jer/Bh9u2DV
a8rJhij0BFw1iYssLbBVJe05WBQo59x1zQxXWzrS8PtvkZQsg/58tZsHWr+PkoUC
gFPZcc8y5UtcE0cveP/zzdv0sVOdUdsuYAm+ni1FLHAiZqN8Pi0VNCykWq50BTRZ
vasIONh2b3NBt77St0Y6GgVqUGuGrwtg4+LUpnSFV9g93K2+QzV+0sa0roxiponv
qpLrYL45LBx6RLQkr0uiGdabR5QjIO4gp8QVBuggM4VhTAkCbE1YKYQAzJWwfoTP
4i806IKptOCLOwjWHo0/PniBsUbrhDcINEETxWJxgrt4QG+behjINCLYHEXrsZh6
RQiA/O1I+tsSK4KyrRddeqizXtEQ7OXH9BHXmrCeLiJY7jo9rswzGIEf7fv3d+J5
vNXH9p3Nr8wuQsMKvMhjhIMbNA3LF7/99fPJor7yuYhnAbPdYyJXiPHK6fYbZSW4
NuwVtzxLiDi1raLxw+n+uj4BXSxoQjA1JxDn1b2+6L3vb8n/N+Drvq4sVFHk0WVk
pPJtzXDj7lCCoUooufaAPDzvyCGTIYSHyomt/w6gRjsJnchMiZDy1zsScLNgBwqS
5G17mX2dBbgVobhQk90Lb2n08NcL7n+tz/MRXFOrI97saBlu+hZo2ft1bTHe10FK
AYCDdsKeacANhCL4fj6u1UeDjQDIqwTzhQ+i8fE0GNU7Yk/8SwJcABz51a86kRuL
DDcy9I4xKulqn6q6g+3sLsHmUO0VxrIbN4aYBuSZrtBHjy2R7/CEcvEw71fw7xIy
vetmFJx2iU00lUR4Nq8vBA2H9Rp+Ua4eTIjHv6uCL+JNJpy7qdqfSYDq/7s8jgot
bBgFzzW8mRGytUmkJtYDm3DKcLvPFXxS8eTjWHZuX0W/au9SGEUTetz2iMM+VV2w
jVwkkljW9KQrqCLJiFSBwar75fFg9cHzhbkTsVfkhdSnfzsnandndfCg/KBs88IA
omv7SMsL3ZI6As4xMFAc9sWkhQDKRThTw34TqH+eDyJ/+qOxK2GAVAwYSJrdG/Cp
rF5AWw2s/ZbviRYiffr40sw2OP/p0iTDxS1mlSrb5zsB6YS23jQ8PmvoOB+3BIvz
OnoklGRhTm+/9gE9lJgcPUDxs6xGSMHRdUbY0zYT8+RyWz2PBN7VNHMWFa+bVpAj
aveFPtsP8tc8VCQhtrP+b+hJzNIJvso2H1gLeQYD6Ycws8CXA08F0MmKZUOUiPTU
Yd5W6iOZZ8eVE4lQhUyY5snNwAWyxGbO3MFieWTDtlwQxgSpwZpzALRfI9mmHzfY
NS13PmrzhbuSSxDC/xdxKKOztRxAsRqBf0Exi4f69UMpV2Q66ki7MbdPREkphOpQ
dXfT9PgsNdLEsSIkaiLbwOayv7KL1zVir+IQuJDqJ7xmeCAlfdLa/RsPRy3aCXX9
1GZmTmjxc7WupToskG5JzD2XNnjWzSHbOBd6ebTNzdel22LWbf3oomkHPZpWns0U
N4Foz8/2Umalm9iu6Bl1UUzDc1O5yOWD1NHG4h1HP9vIJiyVANrJphUD1rHENbqc
FQQCMOEff5ukDgMm0upAqIaCaMGZVRJeL460dO1Ssn7dQjgWsbA4oSvCJWwJ49nE
UJiPf/TPM6dpXVRSoimKQM7nIMbVMa5jgUk+tHBlju530VWztbFju2bkNPjDBx6o
fieF3WUshOWqt7ltK1Iy2DztDBQk32j2C6DgxpkRSVIc6qoIdiOGwP56417Hw5qF
6L99XjAeRD0V8y0qS/2nIYT1hGu76LQO2f8aH7zXIZnLzMhD8UXTBzEOExZt9UST
1URxp9SVgg5sF0HstfprhIeStJWfq2qbr97wUXCzyBYhE24ZKU4gNmr0JUzzDkch
B8NiZF1zODSbjTO4+3buihotemF1Ej/gpFvwaGaNxqKmRIupm7dantxQvu0oFlNl
M3z9vFXCZZu5SBUn9GUAMsHNkyT/XECBauVHhy1Kt1mpAcuYcGYsbhauXjJ6YhYf
4bV+qfcuryKgaQRRqaSGjD3c2jJIKNloZXEYzjbtdhQlSpdm4Bpacp7cpMy600IE
R7rqbvH8CTwEgcBufKNUk0MqYFL8BmRScdnwiXnWBO6dc/OGVRt/bOZ+YPAyCTsM
HCQJeXmPkFC2wrYnHZ+YylyKr7BxmZlY4Dmev72LhAaJEyuUD1ohJ9K4Pg0hL8ds
IZxpY/TkhgU812sPfI5P9Q+WDH9M8sL7UBlmU3KFhQr64d3F3IA233HhnxFWkrA2
TwdObdvCUkVQqiGgMwsEQ8Rx12AuCp4YxoKlHL9ad16HGVsFdFzrNbgpXXqhKVjF
4uwDnY0qjeznYvSZ7MJOR9PSmxItLklCFSiQxvIrmbVD1FXzl+Tw7PMrGy8wkd2v
Iaibvj/1W2Bd6HqvjMLmRVWq6nXP5cfTujvt83BY1YBr/0zQtAeWnA7szg7FOe9A
mALG86UONiRBTo/LKHx42x6xHraoq+FYMYX+CHVXhOjVxFc8StF61eNLN6IcLQc2
FSe9nGu8G9rKpoAm0EqJ8FgQPxsICuni1ik4caltRBbsZD/kqp+Fmp3jz/BooIXI
gDeUm/ZmpItGzI/qCThyZ9jrbagHualANGHJ/SoeiF+OKfRCxR+ROZdObJC0yy2T
fB3Wtp1OHBrWVUh5+pWnX0t+ejDWsqTGkW70LsRPfEieMZkbfVZjvHIJ2Yt2MG42
+L1tp4YwolFly7NAm6O7ScGUA/fTYH5kEDrRXNqqAdLYuLu05OWfEjx+6hTgqnsD
+A3WiZuGUf1LHjQdyj/Dx23pTV259Z1U12AaHje4XSgB4rcdilS4x/p1PsQePbxK
cZO7eGSePqS+M9f8PUtvNP6v5Q7Ak1NC/zYUXGbCw5lpjF11VOLp42B3S+LI2cNb
hwCPtky+N1S4HCu7yUN8CRKfeyVI8G7MUOZ8lqXUufIAstWITQwK4LVb9slIxp0/
Da7xaaTpe1/FjOjwaoEEnMeu8ch3609/EhG1LGZVWrNzIlaxT8FaO5CSN5mVRmtu
NUMNLOLT0kY2IuBgJD2CeisvZ+GgGanpH9n64+d6DZQ9Tog2byXvekXPmqiti/5o
UwX7HnBl7O6zLFzlUEST9OpRpw50/581v4Nl+b2fSqXLfOsrIpfgdFPDgglHf8oe
KQ3s4rzkbktIRXYRzvjZY2zmuo+/mcCEd7btjhCOjLl3y/zqp4PchU+UkT/pEpmo
UMCTL+eOznioGj8ZSNVKqJerAGDCUgfsaWI7vyFQeTGpDFXBNAuNyS3jBSyfZVx4
T/cZoHpHnEnxGSyVx0qCzZlGVA6eXH5X2nb5DDMWsoCy/uv6/kQGj7TET4r07b/i
FbiJZ7FlAkQ4Beqb/fMdytT62K7CBSt+5xlGlbjV0MvOfX36jW35CTsiT+40BCOI
cFzEtS6t/uiL6vvc9DUL1Ig09eg1/ss07RiBoEXyL+ouUR5pgi/VVGsgfJ4yhdjm
CW1hZ/QAyfK964XLjJBIrUl/ALe7jw7kGj9lDgUgYbpaL5nkd8zhyFTZ2FXznMjP
L8F2E2D7njDAvdKxfcY7OWNXQ668AaS4b0+SuSojxIj5cZHWxYJu/0LMWlQeNKSd
uyXt0FYPoT1Eimi1svJzkGDdIeePRWkuHJgPoaxj0QhZCXdoxfnn4yFIDqrTqHVC
kVpXubkMW6aNuippH2d77szpSYUF/DwwiX4VnhCdoK8BRgX7s9Juw26YimkISJj0
jNEidzCdNNOsoAoPm4kj68foi6ckyLQUrn/MSoZRl6b+gJLfzjY7ONp/W1L18yIM
2+P6G3px+Q5iXKYIrHlKHKCxVTJJMBppXBHgio70JyUIbJeFSz/biHpP5bKFjnzk
tHrztRlMGt5NHJ8y/6QVLngoqgTpnGRuTRZW8/wD5VhzlmAPA+rFTYTcDj51rpPm
Uizj2n6V2RzNficucgtwHFfc46hnFdbl086VUXQZx5RHwOPcnqbuWxRd8/+10PCu
wATJgZr84OStakBLXayGsXLfmmwBc58VBfJObXT4VSafIKypFeyI2Y1LZOIfh/Vo
n3Uyve0Ndr+w6nr6duKdgZgP94mqI47bYtjULR7qKkJ3lNSKy53eNnjcSpvw0Sog
BWzDJBQ3hExDPyoMhV86X8rhWUo2vDg80BeAdNNzDy0ecqKUIqvIsCTxgveMlPO7
EYznSDSDbIjEvG7PCylxvZGQeLqaiS0J2k772N/CRuf4nru5PLqPtd5TeDCKbluo
8TGwBj8XmDfDfSRh6HhtoKB8eFOxOaue3o7s8NNV36RpKOnh+SZ6dH2zYCya3FOE
BnR/byxMbWjN+AU7VLSKO8/NUorijCQs/F2wCapJorRdDTeyx1uIc3iCJW6u8/sl
slF4d62XV08jP7jon/xk0S+InqvQRiJMJHzrXJnktYib6VhVohvGaWt9uQEFs0JR
U2Fgz8zNqYs6OiU2obdLzBq4ZYwDN+RI/vGL5ptGu6sZP0xc/F8kn5LMSqFVSJxU
iHIsTARTSIIUjHCPRGA9CMLQOiamUuKFQCjsaayS2f0+IVY8Feh/O6ejhVWMg8IP
kJeUyW44QZlVCZvEH+cY0235rlwb5X2Y6ZzrDxohvZnmiYgoNvDpnLbG8eBYILiM
m9sRrBPXcpQai8j6VJ4wrPhmGU0tn0H1ZybUFlUgZkuzrMrDLgLpdDyL5cuk3dZM
j+NsdHVhZe9ybmNLrP6Ynv4Q1q/KQEDWb9md5olq0ZmPv53VE8fTR86OqjlFk2Oo
7gRdxc2OjFiUuuIi6mbqM0FWgsq9kK7B+B10Uo97BoiqCdqaQE5UU0xT8KHEExTv
/7R+y2vWu/STcYbZjgeHbK4HiAlNidpKBKv3+fhdGRuL+mT2lrmK47P3XL6Kc/Zw
90axvvpM/m6ddQ7FLAXeaqMmTsHsfA3TIgHUe/3SPT6FLscyxj1uxbifSta7OEwU
zySDfyhldxZLGM774KGbpfZm9bE0HSry5fmgi8Srbgz4tETrqzh0yUa7vQQ1QJZM
xgu617XbuRvAkYIs9ArRzhoTLRyvxrzsPqywrQccFHlDNWMlCGI4OpnFl2pay6my
5KBMIoldnmmNQqExk57nRVTCdRFk7+bmqd5AlTlpEMUohdAXlZlfu80t+xOpK9HB
ZprJ/nFCIoVl40wqRmzLBXGmsiZ3OES9wtLKeGzLR4SvYTuYFjvi/HSZlMp/rN/I
9Q4BC6rIf749G3EhvynauwS0EufZCkAsKSwugZgeXRFSU6Qo9Z10b5vtEH3YSpkD
dOxKFskvWzp4qHa8m69JRkAU6DAKNvRwaAxhyWBqNNkq0UmVlpzbNguGraJV7KKU
Fzfqg6t093tLujObWetRhxwZXNhscFdIsh6VtV5HW8ChXcwTOJTzuEmqMaTN+DHf
GiG5T1Z8K4sHJzKk4/j9aV5jTY0j4l6LWXiDonjjhfeKSIp1zBxlEmiiqJ6CyrZ1
Mqvc9j4lU0MPyu+KBPR24z+5IB4HSZKtzyK5nbCx4AdDp0cmwAJQ/XL8jw5wMyJt
dy9AHxMAdK3aROBmpUkrzn3OfS7T0v+WuGOl3JVeShLsJ+8d7hjBvGKogpOktrAi
LfKl8b2+b7a24d+YLNp7z4xrOpmaJoFsfxgfr1sGquo2nkNNT77661mpWVi5D9Ph
v4+9OfLBh+zqu8QoXEs9nbp3b3gRuxGOBAD2nnSCFInWKhjzQpNB2NbXu5kZpVw4
rlIBFx9uwy5UaBP7xbDW5SiXdN01Pdof4ReU8LuNuAO9QBxR5YAXp+bVtJTFpv6R
mVwj0vDtf+zRv+FYRh/WZa0bTdtQPVLSVEi1bHIS8NLOs5PG2mnajBTCX4i6WQeP
CxJ1bClPosUZYLQ6eQ6IaNFWiiReu+DBYm0Q5R+NHcMb/nmNgYrF1h02JSjnLOXl
//6c7fNfW/YdoOVVClfSZtfJS4XQSgHGoRU7xMNzLiyawPXwilTiJ4M+iqWYi4TY
aa8A4Y+Scv3uQbqtyXweFa1n3Fec1hruIU2IAUbkn+laPdUa9wBT28nIIezmM/qo
FCgL9LPPOQGDZOxEPLzQ0cXRnYLyxQubE9+NB7GBZRNKLRMad3nYlM+H++DVcYDY
5J1D4yj9B1jus6RfLeTrjekk6FTXp/DRw3uWCmVAzlH9Xo158oyiXPit3Dh4IE/h
GDE3Oel/K2DolD51tSNUUWY0oLa7EtW7hrsfeCfGjhuY6LhmVgKECudbKbJz8apm
FPwALaR4irUid6TcnFOf/33w/SsEplJ9xsjI/m4kTyje61qcJOFfjifCGEAZGbIx
OTfjBFBFM+u26srpyUMv3noAX1dgZk1GupwItzAoYgF9D5EVxPrLqrrLuH/Dpz46
F8Zp8h2+xQnlUdYnr/O34+nCK9NemCYjLkdlYEuVxjkRTaKjEfpZDfmZMUZA4Wp7
vML4VlfwG5MvN+ttyk19Je/SrTvn0G/Y2tZ325ZwvYA9eJUpMFQrwDgQ3EyvUE3k
232IQ3Ow6+sfbYOPeRDVkkEO2n8kSGstt2aEhsw1gv0nbTwT4Dg2491E3Xi1209e
jXauxGJDW4su+98LohyMT/Y9yj5AgJugPM/8hzU+cMf/zz/lyjgGCJITrQyT7Gja
yNKqVC5ZsVGzTbv3GewJyAq21RbnR6vLbN5u5mger2yi73lP3KpwYMhxHtDvhXd2
DzZQ7Mpt0rwnFmFVQFaVfeIOZ3jqERd+Plsbniy0HxUjuJYmGuFK9OV2yGX2OucP
E81YMfPUYNjLnGW27ig8ecypJcRgsbmSE/zq13CK7AGBaPRnsrEKq56R5/+UV0JQ
ptdRCTCcVZamsWW9M69ru3zNPAKfsqzG4cROFyUtVpXrMrrVugTtakPJ7VOSf4gW
lXH5oKYQ2i/MOk8YAC7R8+seecHWk6cBn8fKKgX7zpOb1jq3kRsrTloEOXsg7zrA
6gXfu2lpb4C/x3Slu2RZi+hKpqgqvUD/VJUweX6dR/YDV9+HbS2d2l1PVtl7agI9
mEo9djqiiZHYl+OmBJta0nB6Naaki1LvhXRH4JzDRllUJJMzGVajZ4/fM9E9YLHQ
sZPs/CkcDEbPatqt/DlovnlkYG4oXTeq16l7YaOPEkiZ9pldOjzn8IZ47kTCRj6B
aEzNjCjvNZKVZYBLeJjNs8GjreYJg+ymmR9t/5NxVj+4sPrtcZ9xh/JnIqaYrG3C
eP/FXCdPD06VQj/yTPffO6GA62zoSu9xLOgBVWAFSooyjCchCfFxETt+OKJ3rbEb
gxOq4V8kAaJ00TZ75g4YNzC0K3tcRnPLO1Kc/5NbhIxm/gMM2ooJ1unjwPAUUBqv
dsn0UF8rB+0GqWRkkPGo0GFv0ZVqE9HaX0/VNpG5jBDxD1ZWi+0RCY0rBL+rxa++
u6BAnffL2inQ/dGwFU60QTrrJsnnwH3Jl97a32RjirttvNa8+mNj6NpcUe9cn9Kh
NGVDf8YcQ54F2ib+FHWuWBVf9zVQixKO4JS60YHGZlxCSrxDYRVs3hcuqRzo7m9m
jRIwTV8XugJUwJ6PIZIfcizjR9EpGaxdYrsXQi1WzBuYTsoKsw/6Tzr4wP3Ud8Kv
B2oDkMzKvqySFFTtvkhHoiDo1X+q1UzbF2GoYP8cUbBzTlyFvq5IVOIM/pIC0UfP
F2JfUkVbLw6hVLgbLdhPwF6HiItF/0znPIJT+PQPrXh0VLTfHAGiOyQPRbe31l9R
Twp4e0y73gu0948pRw3XFl2Ihi3ZdlmDKN8T2lFjj5MprGhppaBPLrm4uqN3pk6U
jlyN8AbemodCs+Z0SxVXIxi5Fif1R826DlcWSymdvmHS+wr6fa/A6gFsfQrKGBDS
jkGYHKry0JSOIApgDAGjChnjk6yI/LzwLzuWwc1+bipaHQD04JHp7RPAHGblKZpO
9lgMTHjnhrMm/yCDqpqaM3qa2cbbU5n893AnfoUNiYsIYyue9Vu7Z5e1XaFQTs6m
/OZEGAr1InJBVELlb6rnaw+FBnCLuZnzKuOxXB1yVpaDHt1n62OjXV9Q5A4yQhuI
0xLlraOPbPSCLsgtQblIVqr/Zu1pU6f9utwdF5jp8prkyzddxkF2/etqQaBnkqZ6
+JJk6toIXsdTs8revzgqwdIbbEVaY+Xv0S1RhfT3685DeOV3N1y83JouHg9QFdyK
suYoho2E0WYM3+Scjy5ryYvuJHylLYBL/Qc0j3LR0U9SXdvGUz4FylfPnVBT5vd5
L4EQVEfjlb0PWtC+PGL6x+hMvWHyZwRXwvPd2NPvCiKWO2XbCTMjbV2fLB8R6+/w
k2bNNrLpzes5iNyM0qHSwfrDlagEzfGZZNGke/NjyX4e36ZsIwx3jrugvzIhYF6s
LqpnyllUOlSVTikn4r+8WEmJBGTaqrTd7jR9DqYT5exGJCPHYUJjcudzm6Iq1LS8
dJ3/xPN/V5ZrZvFSpSsmExB7HfXyKsURg5zq14Q4faZgO+CX9caf+1aTaoaGgY7U
jaDAnkTmiQjzPtrLMlr6xH5awqIJ3w9uwaxaiqbReCXqovmar71gVW/85GiYNPmB
tacOIZ/W1Dew20HtJ0ExqLGtLklBWqprS6Y2Ep1POMsDGFww2aKWiVs3tKIH8KKr
OfwXloOV9HTwJ+qfmn2Ubgig/sE7leJrFTTYIVm6vdHM9jkSAddqnV+B2as+XVcy
e1mseArhCPpcWvtepDNBaFJhVG2gd4KkhkAvDNZ7YqqMKguhLUUAJ9wCJy4OkHaI
FmF1mo/9uxnwxOpHBkS4IAYSkJ/HCW8Bct3SEli0bgNL5JUGfv88meheC+ewaPGr
JinKItqrsdWWdujoezID3dJuhQtTUEHxoDGvq7k9zqfPZHaCRH+Ov3zp/WIKZYli
X7H80z1TR1haOEskhyiHFoecozUifV/gfVu6nhtYIBWYKkUkQYNGplC95OJw9I/M
XTyjXHpfKuhDFumtTxwwwB6lehYTdrFTmeuqoj81fQ6wSVAMzf4yjybHN9gupn6g
JFEiry6RVAdHf+kfMxAWgjhkIy3bQzh/a2s39+i5a4yLzoSUdG4YhWrVTKP5EDdJ
2Hjt4y0DOJTJxscXnUsjG93D+/Tt8X18g0ej+W8+wDJcf/piWLIlZAkZOlm46NV4
PzQHOvYRDDlOpDNMs6jZFtbqR9E42b4MvtfcbAJ5lUoOmOdnmyw+VN7G6O1AtIqw
LoiiIu4TQuxCe4zpex0d6ZruuO9EmlImgItNFW9Ih4hBECUchwwGEHbWI7XuoeXy
ptLMqVAJljW8dfVn8sAPor3NmWyPlyF7VTR6HdbMa7nyWALHGNgp4FJOUW/t3C27
XQGopEpnarA6sagEicg60TsQVVC93sqbW5csxm8Vrx9yKeTtIhRq9wRhn4tLQ2TJ
ZfOxA3Zb2NlkHstCktdib//YMcLOWkiZooz3NFe3lZmNZvxzu21vgAmAulA6umPM
nh9EmTFnOQztGkti2X44mtXOP1WIdyDXGbVyMRnEWIwMfOfQx/QRRGLPVLfGHOk8
Mw/vBOWwLBdC9gigspbhJbevu6Kgz+ASauuO5UCs6xnRsBKF8e4MojPpELXTRCoA
pK2To3dgWzI+94mqXDLZ+badofJ0BT1dZVMbc3qdoBRGe08T0C08HVVpuMZuxhCS
dRgJDRu/UrALhszVRB5CntEW2ktXzqcGZjLn3ArNTq+q3PsNL+kwT+W+JuayjCsP
CriDC07bdohllS1bfUraOWKEwhM4GiZ9vlj6iBZYeyV5+T+PXCZ1xH6No99WIQGV
lehtB5xdaPimI08nAD26F9lwtDaawJuzddQLj3frnrrDGaZf7C1Y6RypGGWQfXjx
ePxrBIzPte05tmAQ2Xl04ddXHfsVyrMn9pZ9a+gPu1L6all1jd5DTlLKzLZHehYV
GlPVIaGcnCx9VzgcxcmlA36w1W9hZ+soyxWc2auymPYMZOVZAwNUUSa+N48d+Gif
WZlvrdYrM5D7DSTWH4dRwsnofVIXT8iBohpcrJYROy1wFcnxLGiOna8LSJeUwQg9
2MBLAfgK0HExEIct1jN3eOwFbwz7ysjNXchpF5Ex1KpV2Xdc0uXSYHh6ePi8IX0q
vonzLLu+1WFzZ2iWNlmFRHfxGTf524fFsM652AQWeCmlmvp/kEPzRgKxAE7jEYR/
6/9qJloXHVDjtp9llLua+HKsbxDBPlHjyIya3TjnWrgW2nhqZVU2CetwclRdaGGQ
Rz/InymY/Bw2dMpEcPjI4p1SowENWjcZY6J6X70FSfPkrW8iwBIROHZaslbRXI4T
EcTVmU6APwpLPDjueRB4+MNS/XhVrRhH3jqPzmmKL+6DNLB71k5BLbxUiPvUV2/c
uRZRCEAZiAJJf/gc+caDFjOzXsFVMjm/sBM5/f1R8wvNWY83KzV+7fc0g9aJYjOm
kJuKo+C/3qQhRfZovka5z8tSx4IpuAPpZpFnb87+W76wdwXcnNyExJR/pjB7ZJJ/
1DVSIrBKFOudmaSZQthdFJHT2fjzRjPqF5II7m1ObS/O0If8z9ulJh5cCz3lwhcw
cgnTcWI+FJihSO6Lj5RGXNPeQjniNMjDaorCWaoWIZGrZlXL/lcEKkRvaVJ0ogiw
s8McQvl5bR+QvDE6PvWZLX1MIFvHQQcyhoMnhHcE0KpALdZV7OVvwCZzuq8FnZBP
A1P0I52imGUQS3xDS/LykuElMfQ6mQX8hE558rQlcL9B4CbQgYRgH9zPLXTlvmBU
/oReDyvp6c7OMprTsXsfnFoFD4OWbzilC5Xt1eopEHfnH6etKOT3u0pW2ddrSvEH
YzJfgjy/90hCLRdVbC5oIw0rhueWw3uy+KzHuVCal/KgZWZeir1fF8w0Ac7S3ahu
+NTqMDhfxpDvf+Mnz/s6TTyywpCDE0U/PomU465LS2bR63ee2NLM92UtrBov2Izz
cea3NTRZeBAhOopZJFvphlkx/MXh+V3d3+2Q00YWzCxKsg6nRgZ0e8thp8Bz8NH/
LWvWbEj2NXE/Nbof/qxiDthn+tvQX/y6bxP3o+RIj33eNZUtU0i4JTKLwQ2cBgRx
K3wFelyNexoRYTVoq0ysrg4lFHdJQ6qkBhifwP6oPcmkLaQW/addLOSokKPuf5db
8+OfekbVxClTij6Y4xn29fMAvjfRrYsv1lR1DPReEyNr7qFk5EjIvZ81XvjdVpRb
9S0tOh/K0OtNWwuaSFjupj+oMocbJOYy0NVgy/pl3McJdOhNBjYLmo4+2S5TE58F
BvrceCApXXEcolIxXPsQwRmCrLdXpx5iVSRtxoKR7+6+FEkUDnuFuLir8BCVP3ts
lYjFY1w5Fy8ni2qsTkyV1rgo0/zYgYopHBvVFjFqNvyz8MYKiAY042VQCQmr49Y+
zOPOLGS5i/eMEb/4L1w+5I/l7vWfCaXeUoOUzKSDNshO14LQ0iTJDn0/evOiZadI
mHzK+ZXbakMwhxTbTWKlDDpzZxOMzbisDwlQg3vvH3y+rBSUqoJLoupnFeAP889D
4PfH2pfdGGBxDu1chTb0+VvQauAncJTAmEEV9y6Mo/kkLNgVcasoIAB5qtoFrthX
PXNh/ZXhXDh7GQYKko6Y2K5Dkx4WUO9uKWlV9a2g2dl94JG0VA+QcCYb/fS0Ep1z
pYNyb9mFOWGpTJDg6XMjmUT18jcT1m8I/4AFpjij3dLVvV5nZliBS9Sq/YrK6y+Z
d3d6RHNPuO7QTg3dM9fwP+FZMqSXZHgw5if8c79XTbRRGn2TAqpJCxju95dcF7Dw
Sz7v/F6LlVZcQxUZxQNPen7RYpZFloydK0ph98Ix94oXxFtgYSvJqqxlReMgGG9h
e+BaK+v8Q5ac6tDlbCTHBUhMhMkGgUWwkxokqxqDZecdOBh43O1NxncCqUoxspYJ
8iOtO2x1hq7BgWhEFyl266K0aQzvi06+Yk3jiNK9jrio87fXbsvOhdeYcgJLseGZ
cV98h6/pTwB5W+BuXEEjXdg3l67tkq/h73jzZbHQUdbpHGwPaE90OYIhpoxlEFOw
+9DyPehv41p/xMP3tlzMkJd6WzgIlfZzUsYoPKCcKaoerRqM4+kNuCx3B2nWwMHe
D8Tq4RS8LO3zJpAWPZZV9vpGwAxAnOYa/2QRg800kjLJ+1vWrkIYuiV+1K/F0j6/
yOA/kRaD5Rmtd041+e15reax75Om3uLifWoJ9wd7sY5IM6W89muNRNYON4CF2zNf
RFypfEECLXHqPlst1nj11T8Lp0M8WLHs7Y0XcvYa03Y8sNO4zm/WAjmQXM94d1Ez
HYrzd/TH0Wrj7rVtlcGi0GiXROXELNYZRwoDgmJsIQpJRgSnfdc0C8McSTDq8S7T
W/b4aNDDv0n++JICUdhbeRvCDqe6U6zGwf4O2VUQZ/9THZ4oeAoi3q8z69QJcpQu
PmWhbgSXGJDqSewO/p9aWLjpcX1nszsFhqWAefO36i5WUtF39n9ia8Q6VH6bS8/K
VIhFuYJIVO6NYG0g3QRneQ9PWcl4u4BU3Py0jViv6bSCaC6mVKc2QdUOFCHtVCv4
lRyjecqXhmUKoyyyD34D3iXXAt3cb4qKl9gw/54XDZRUtItQg/TT0vk2O4WWmTWn
+zMUB150rWAMPo6Sb69q4LKisjj+WXgNyX9phqByOItXQqw0NMJ5/FcN7mSXx2h4
D7BroG+CSjVqFNZ0TL0b1cKStZapTMmDHhMva2XBswu1xs08VmDcIfY5SsP9siiw
1P0NWCcwy62phJEutPHKz55RqK+tueDhxOxuvrOJg2OPk+4wyIcQMPWfLQmcAaLm
juYR/0zwbernwPQoa0eKISAzYDTq0thzfb+Gfp3piw4c8l8s5d2XBPCK9KxQAcde
UlnmerwDwqjcrgnA6F2eFJ1iLuucYS85loy01wOU1rS1E+n4KKHQhac36m5GhK3r
8RxnQk0f2uzP89kJxOLdjKV8Ii4+166iJycDR6NAKqIikUtM6YFqTFVFFuoqH4dG
OYopuhgp75N1zi2aA4q4hfOHRVK3GGHzirEl63aH46ItUBoC8mqtHGMpuk6Bbj3V
0gOrJnryLfszpxNE8xIvT5StaIavcdbvRS5DLmM8KRKxN8oYdQBx0JslOqwnNaQo
iB6Dnrby/c6Kgax4Vg3BzDPc6Ryhe362vBHBB+BdnYjzG/ByW3c2UJlWgk5JE3ty
5Cn6XH3KiYZ864oxDIXI2wnEtDU29Wrb/N2ma0xrHCeE517HNpIV0jzBQFBMgDz+
Az8MTxtrR4OFqu8zMY/qOfa1NsRSkwzZDL1hCS0x02lUjsQLR6xQS/v7AkNEoJcF
sZy99eIlzRjM3DDP4aiPqhKJSlkKjjxRypDEYYAwGTQpNccM2fHE73T+dSYyBKOW
tBQr9ky4YAPeZhrTAzpeesRB4Nn4pXvkRe2IkgN/8baNjPb8gO6fTAgz23EmGmfB
YN8EKkGdXua1lTzqndqPmC1n5Ctc/VfLtQuXMsthYAImKwyeCkzD3URIMpZFaFP0
5u07SxiJKlk8pfgjKzqkE/McSxsodeRH7UT1JKOiCVS2GrQp58mrFYfiPmpoXSp+
OWinwQohc6UC00tMd4So2ByQsdeQeKk1uu9sN2varRNpb3EESOqMPIhz0eQj7ykk
bxEygR9SMsai+ODR9EldhX5sawYI6liSrHvVk5xwh82g9FE1RrHku/EVqgf+BkJY
8r9SanxcfikNpr1wANSpv7xmVUjdvI1ePo5hqYb1PBezHfUld/mVDsLPmlW1XSN0
fC9r2A9RQMW2M00ErxPiUmZ628iddcshHhGZnkomUp+Q0ybEh5rGZ2UcKF1Gjt76
uKaSAAhgdo5oNWyNh2p6LPzRGMopSD+3WTreNkhkqlnV6xtsZAPscYluEJbu9lqC
S/0iaCLA7rxSh7D1jCgTXCe179WVo4+o7rgdihFfq266qii3zpCgMU7rRm2vfatx
42xYiDwgJYPR0PaihoYGrY4Scbczj3iiK4CGi+7Xs9kL3/faG2RkP7AGm7/YvRDm
nm5JMoETZcmyOi5nmCd/SY8t0c/LQ6DbF6yJniSxc6CBPa/6y2mxiar459uUu4UO
YSKkpKJpUuGtxhv2tqnAv+v/3vu4s7NnCs63+Fff1hwUrTxIv0CG2bcra6xcW6WN
dgvM4jmpVNns2QN1/BSSLYTlNG57y3y85PafUkYtEPeudnr+yckYMTsNtQWtQkS6
sRVxZTnPIzYjxDahz74EBe+rMYWA++Z6H5r0r7J1cK7u00GvJlpVwuVU7BsbPd7i
YM2mOS3J39mf99n2FVhV6Dq1mJAMWakDoDsoZrYfXr66O/lmWwuqScwObBW2Zt2E
aT8XBQp02bJPog4THyP8v1CVgAyqIO5pSyrbWEdFCxQ7aE/WLylk1oDNFFUr2Vny
Ic3IvXhmLOslN2XseEJFn3Ih9NpRqjpY5iW0uGmNhqrJl1iWpI6xAW9B6gCB3NJy
Dlv3tNJHW0yCaB77eaL1QRDWs9JHsI2Lzrd0XVOz7ZtwYlG5YNxA7lc8Qha+6p7x
IrZpKxKt/9lK8BBnOPVHVt/o4eC37hYwqhcJmWXSHHbSG5O3roR/WixQPefqOcKp
Dyq2COV6JfbE6j6+7nmxlXzg+vgf3UC6fPGNWTfbBgfY6BVciXu3h2DgX6kvCe56
xcZDxQmRFG8Dqooe3OLI19yjEh9/5qAtyDEKKGYJy2GhY+joi050mwRKUuwxhHip
VdB8vX6tK9MToU4lBM9xFY+bgGL4nNTLbipU8aPP+JQFFlUJtJKppRdj/hwsdRAP
PiWIyUSNlmNB3ZXYNLRJY0i/cAtit6vZhCfQ0Sq6GyrKuadJxZGZuyKGwFr50SOw
O+fm6k3z+f8gDgeNk0K95ObLOVT4lRgqZfnf9owuGvlAQvxdApHQFU5g9w7eQzNe
TVQbp7TvjVMFvL1A8YCysZzyHxAxGey51TIwpFs4WpvtFIjv3eF21TIfU1ylGmu8
mVjccwEUnBuTZKJcdUTo7Ssr85muPOG5D9yXUtrKPoPCMDgOnNPBzqi1+NW/2MyJ
Oh9a+bFZkdQ6kyeUhxj0FRuk9OS8KQGVzaiTKfu7MLl5/o17GwbIZijZ05Edd+4t
wsH6wymf/R9bATfvrRT7d1stPgHjWHiTMeFke1cRolHJLrjb0ujkF1a3K41F+uBH
4Mkq9EEiNfIawyKyfAZMa81tL54XkPHVjcIqyFPjIxl+WoeBUiaFNsQf1PXr07AX
mhE0MxTdinPYz2ECXgB0ccUO3R4mtUbeNICoomSfSnuC8vjmkq8mox5JlqU0BiNU
cebxl9Eng70buLe+b7ANt9GeLvQUw5NdldG+sp6ArgBsievKlb4dEFQr7Z6c1P5s
0xRwVkRdgmzdj56vX76mArkEQ99CgCP3r8HETZm52++xZffiZJVa2++zs6DVgYWk
U+WsOMxpH7oErrxt8oc3J5aQn2pp+gP1o1PorOxqEhxAr9RlQn1B9g7L3AWGsbgO
f4arPmNaDdELE/IWs28KKVivwAvNK7XGBefWnOn07ZyuFg7i7wVm7aiLs7cCF9oT
lLxGovnvCwTx7VG0XKecTKQ1mco6U/Dq2eAWYC/WGP+AbbJXVasEvt3kqOI5HPiP
7gpOlPZcnNzn2THxA1UqTWlErwnZfEWeDh30ksbK5H2Dg8+cvy91BhossyENru9+
t1gSk/sjqFmu2879ybRqjXSx4VY2m4N/lDOz+wMwA3I0g71yjLlTg/HOl0WbXOGt
F5PfeyEqthSK81oVAmrMeYWGlQS9VeEFCTdh+wE1tf5vPLavQJY4W5AQZK7rlDLi
vmLuRgQ8KdxkKANi9cRaR5yA+yZKelAYx1EurZZtGJSS2yAbT4S3/+i1XXt093bR
YH6K0wFTzBd1GXRP/CmeK6yLWAJRNh0aTMep2HaVyP+u6yn/399HSeCyxyWPh5Dc
DLP0mZ+Pf9BvnL634geWd8twSETAoQxA4ghC2EQdRWcKjG7nfSGHihiZoX752OYL
B0dGj2ayzZBtJ2J8QH/wQzW7TKfGIIthH8MWehYRoyB6V84wiKFrE8G/XNiZQlau
NCABBX/AWDZjr1RDjK93dJTnYHtCP5F2aVejNct9eefo3Vc7r3bkOyZsfZ3II3Az
+jC5OFcg9Mlc+wks43rIo9ox/cQ8+ik5p05Ee6hnVOHFIHk/I+DeGOK+60MQi3yn
smyGJIsx1WHoeWPDgD+zrhBx7C7oTHRQjsjfsC0VVWyhn1qdtPgz6Mn8Vz6K+hV9
69Jex7cNWfIMWzlP1XbAI+sI00KP+nPzfO8KKF094sbBDs7+uFpKvSYCQxiKvSqr
6ii+FjXIysfd0+jiDKYws5LgI0JdyE1mTvoVe7U0skVNSLPu4RW4ICdGjvf+AB/X
JXb8Uz3e4cnd7aAh/ksBzKbhoK/r1gWexoKunehwGs7xZ1yy5IdwJVKyam+WeK7/
CLRwTOH5w849IxDd9IzuoPTFeM/lWpMd74AHkCm+SDNUawfgf80i5Z/Ito4SK+VL
gAJ5/iO0KH2prIpMELi9W2g2puq8ORY+8mxVfO0h3MC5BK/InHJaES0BVnfvntYm
0WzEfX5RUjFxNdalyZcK99CHlVpCRmufBPs8MplB12ieRLzPVEG+HsV45deJ/lCW
BQjJ96kCFml9ddV1KNq4As8upup2XMTc3keCopchqi6L0hNEpXEhNtIA9uQ6vIcH
exFGGETOAsndwAXEbiPH5UzSBzpuxVFWO9Es63itwKDs/Ie63CKg12+LLx5+DUo+
TsbUb03rrna/j+PVvduHQ9bs1bT1sMaGWT/rZKNIPOo7CR4r87e/HUkHSuHWUGtr
giyBGuUs3515rD8e0+HBzZB7YdS4yF+BZqLb4rJJy7Bg2WuaX5h/E2z0LLfZZwEv
3PboD+q6P6VHP0pYZ32GuwMkHSrjZXB+CtJaqrDQrVSjURjwa2izL0S3IDlRJJ/A
9ZJAjLxo0wSf/XEwkU59QoNXSUzAkdVRCoIDA7STZnpuzSclsXY7BMnqOXX/L9/O
9kZpkNvwTSR2+ed3/5NjzMbixE/LD7OtiNi+pH/3z6AMbs8jAg89RZs2KniNa1n7
aCO+0QvTy2bmRAog8Ksfjip5VnKprq9XjfTvLcrwYs5M32guJP87z8Gp3mvXnULR
PVxBkf2ey1WibMZIyOVPEguPw0P1kH5q8jY1LsKGJ/WSSpttBBvX/vVRCxZWLAJx
16NYgWJdvKgtuTg0l779ZTqLLNghHD/NXgETrPmhyn38SX+OWl4hWF1Stnp2W72S
eLU/YJ2jgI8QOs0T+XKGTPji1xlCBwa5gBd8Bip/kKYwyq4E4/KexThTZE0XUCmB
09brZmwD4wmCtGFxeIT9j6YRlXZou+TL5g35yOpKOKUoWUKLA81l+6lEzpXhg8tm
7zEjLTwmSv7iA+n+EYTz/UkPohQOx7phMkUYppav2tnK+J5n+Fz5E+hggFJG5cEP
0P/+ZOeeyI/VSzUmaWjuuGCiKzMK1BY4irstx7NLQdYPBOroqXa1JcHr58urbXn2
pQ/fqvydAdOBXDErVrZtWEayriRaUPTYAV3Nzu8FrFGGBSceaZz5LESHzU/40EO7
RxT4q9QaDaGMRzIoKWXkKMu8KMeIZQkpVOLknXp613eWRPwRrtKVh9uykZR3KDtA
aturxJ2thuUALDc/bkRqGwPmjcgfFI8SMQkTGv4dqNV7/k/QErmk9Y/NANy5VRqv
6+VF34aQDMM9Re4TyIbJ5IisjxW9thbudADF0mNue8w=

`pragma protect end_protected
