`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
BRN1H3nvUJ3wVE+KJ1giaoEeJau8FmqegtM0pO02FBd/znweZpSmO7B9hyEmN2re
SaOjjDU8WukG3Z5xnn/SqEGtjHt0jpRNNjIUD4E2GxTtXWPBdEUKKYVXzMz+ekwc
IS+J7bEu5ii0fnQVsDapMxCrCwZTAHi/8+elBPBCUpA=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 3200), data_block
lBU6Nve5xTI5YU92CgWhaUgslTy8Ldduuhk/FKYwnBROVzrtkadd0dktEr6UcJlb
aSJNIajkccb0YuVVKMdrriQXLHH7qpCmiDJoDQzeyuA4uLdZnpNCcqjxqxz9YzPJ
ET78Hv620x5y5SvgrKkBmvfcwjJjWdtg4EHBPUjRyFTFlGKwKD1OCTPoFN+3Jnte
535cuaiB8mDVs8BowGcCjjTstx5lvHZQMIXhhQ1HIF6GP8GfLxKU0lxUqwDH4n0D
6RPfyYBpHLGS0YB71Jwi90ywtZIkQ176wJiOe92n8Fkth4HC9DYTaUldWv2yZdsw
Y3Nf0sbC0NY6iHQs325/lP8sEt6P3G13wJxS/XYFl+gLOIg4nN3GTjDVbHhilLZF
PIyREtXzTSyOuY3YlwnfZ7ha0AAeYKXDokLRIDJd/qeBVachJjlI5EW8QhMdVSAK
qyVdCRnxCtU8IOcqvN3lqy0asX++G8Va2yCEIpzlnmOQjVE8cPESiledlSdLacGa
KY5m55GfjpafYjQgLJNTU7m12zBZlPb/SpLLraAY0EzK8C7RtEuXjAQGvElclqL7
p7AGKxv8BAvm7A3Oi/DAIQA+yE3h3OU2h7ltlLw4rxDAbucw4OXlrfnUQHtBTvBZ
z86Q+Lhdi1pi++BVcUPrimkeLZ3zWmhK3iRoL+b3cYOoyX2W0wUYrMX+MXAFdJtP
lPEgFMKZbfrhnRXtuVV1q2AnWeLIWDX2ahyOliSECct39vTVukh7iDW/O6TmGRdH
454z2P/uKFNZ9uXn8UkEEndOV7lTdEPcOiRl31f++TxXUYxxIHQ2eeHsCPyGtbnY
f86xAFlVNZ6pL2aO/qHRVwbZwVZDBkOuPNkVk6diBfBswDC0dyuftWQ6OE1HQzVN
FaahJV4VDB1KDnGaM6WIy/lSE7AmGdRC01/u9oSXdrB1AJTHqJrKDpMH5nEVo6iU
zprEH2fqQN1BmBDrtg2XuZ7gt2crOKbczNBKRcCOXQKvaSa91SHb16qXjorVtIRX
JVhUSq8khLm5vU2Xn53col7YUeCPY4P5BjdycOgLMS1ClqbxKc3ELOE/xyXlqzdU
Zh/Vr1Ybwh9L6kNXVA2k1WDTc090xo+ckNWg1XgfLYdZ40UvkS9mPxBvXRywXPuE
wRBQcS5qHJWkLdtfmwdMjWYtwsiJv450QojL03LUnNw1+b3tp5faIKGIbfOTX5Iw
Clytfnz+1yUvmtk768yKE5x00myoTV0uPg+Vq/vOBBiaRuWKU/MruLRqMoV5XjKi
DcpegGcMtXwWtdyXO2yvN9e2A6clSQLthYbIcxlR8Ft5kM6R+2FEOd8O+wyBfxhx
gBa577Azlk+9HNAYYFlew8bLcVu6tRLwYuF8h114tNeYef9p5U4J+y1fNfKfh2eg
kiiKDDk6QA4fEtxcNVrXBLoITIA2fGHs1h5ls7qI2VZrNlF3f6VPw+J/VHQXBooQ
EsCLu+UZIiVJEqZ+5DYOinfNnXdSJnqIl1Dnh1flJa7SjimnfZfW9IkYmbTiq4w7
3QVLC7vSkZqiDlcrj97fsX7vNgpGBCp0iBV2ZXV1tiMHgV9TT1Kdz6cZ8+JOWHZ2
SAf38brzeI6FBK/wZvq73kGAsm7QI72Y+LnINsCTofI654opMvSRkkrbV1blPgz3
7Wy+8HiTmAyUAUzvBBFrQMqRA/WeUcryEuc+cPJJIAX60aNzcL1/3LaubwPTD1dX
ZI/Gkp2I3qFMhBw5g8Pdj6j1jtwvH0JXdpsUJ2JQn72DXYBPnX4Lz4ZMXsoZpRdn
UydVHV8dxik1V0G43n1XZGuJsZrzdOr+BpE4cOUVde6sxPHv+xjjGrlOk9E/J/fN
dLh6kaLZGbKWLKxbrA1Zh3j/6FQtswft+cUmenqM1Ga/heJmLwoztpPxzD7LGnrL
MUoUYoIwlawJaUoQiYZq+ORQmF+s5uyXxI2OxSZh9Yl1iNWqcvsgnOBGF3X1RxDk
W9+VLx3wRYoRkSIz1pUtslHoGlZPK0/yGE9j62DDBhmiZOdsNWqkO6IOB9Ta8u9F
I01mq94y0Lhn0CgcFS3v4nm0/NziEAsHtzjnVq0c4OYCPmr2vWB8jn0S+0yDWZc8
xsgY62CpYiUQCkqm+U+Ete7lPyGiPE5FmssgXiSMikai7DxR1iEGGrU3xfUZQTHV
/zSWlDJ3unWIMd5kIoLCPooSNo0sshF+b8U2/Gy9svX22d90cCBzZfzMA0mMOM+r
2WwdkIMo8ro3RwStq7kruPVNylnhvZVujsY/ZGbujag6KCbjC7GL+cpZl/pcVQRq
2BC+OlNNFRVMTFPdhHptv/30f9TyPiJqL0jF/GzPNGqB+tgJbPhqBGHHLryfI1Wm
KpQtFiU875dUxnVx2uRyLXE4XhwpPLzBhG6A+rdcTgZwMjw9YLBQMEqT0IXMs5MJ
FXmjHuFYtTrmWtCuUc3OJN8UajhIjtQ21GNNU9CLVFcXYFmwR6auY3GfPz1VM22V
/AcslMjf+w0YRQRBFoVZXrbBwJM3eQjCfpvDeSNCSyAvx5SdRLv3nbc+jvVZpGR9
Nrx9dlqmUUYcUrPYPYjuCSb7w8l+NbJbRfI2clIgFV8bxvcQPr4bNlj/LdGQTSXG
DjK1lstppBFY6iggQs0MFB9UWysc6rVszDAioqh+7m0oI6aoEJAXCFWxlioEuMOT
9v/PZ2JLbghh+2YydMUKmtZSytGKAodTeBZ53MH+kQdjy0HHHEPwUi6xLQkjQKx+
Mx/ag888pBrmvUExSuETnYfj35xZIK24ILpV5Is3xlbJiFpeJDZ3mxhDCbupUMDB
vn4AiVptGscfVZsese341c2Z9wJGkIQutJmy8UVzhtK9+RL8HU4gNJnDm4XycrIo
FPJuFJiFaOWVwJwynGlYtJ7o4zVwJQ7JJk0oiVhPg7fVXEQj3YKFgOqZ6hbzFR1J
vtgJ0eN2SlzzPJdhtz35XlcWC0CHSRxQYkNukd/VmJ1X4To5NZVX7As2FQPTYbrd
1YeRCAfS9mjs4H+2iWwgt3uG1X2QioMRGRzdIDEwYhCvs4VlLDQehbGaWA3AwNlv
VJjiSNW+tqjVmhPzeiJcJnVXe6gleKUGz7e9gEaQVh4fxWShPE2BKdWllG/S8VHX
NWVpSNKDrHw6eVCT6xbt0HM9c0oJVOTxojEY6ZToYMBoJEjSbtRkdq6Fgq/okRAh
WYAea8+tdMfrlnmjAl8pE/l/sgAwdL0L8LDOh1YncDf/Obumlb8KAWZoa6iogbHm
yvYUZ9m2iwGfUreDuwuvmukDtiH8m7kb+ro4MQq+ABQxLyk0D0fdsG7L2+b7KzMX
BT0nt/J4NjoqSwMwMepkq81yDli5+J4BVUaZS6rRSwNY9osPl5NtNZ7xiO53PKBG
mYCOGRFnPqrkzMd9dnvUTpCbx4Oqm7hqJ+fzS6LSm0RDYAD0d6YlpSeKEWKkpEkL
Xq/Wd9kHol4dVEYC63FVcynSi+FBtmBLqlSSS/qsT5/US0SyXY/QM9LNwMqhHwfh
DEPvrd73jtXL9j333xkDDc0yzp3i9fFWnI8MWzP+vuhXQmytgBqZ+8TQGn7gaS/p
BxrMNl9byamytfsBuKpEXlq63Ngz3rVu2pJ8ddIFuosnr0a/U5MXCJqT8SNVTjTU
RipG633btdhZvZ5LV3timw+ojqZ7cH2x8+jjTlhhj5msW/vZ+Tia+dzD4Hd3bcuB
N8uBWMe71PPSdljdnvgwOjq5DWU4uvWWpvpF52K0dX+upXRno+WEraNlDrmuzzr1
D0Jfa0J6UuH/XmUXEoMuZFqXNjefhsBaMUSaCOv+VgMA+UY0PmcAhjqKEKlT5Rd4
oz6I2sp+sv2sn2RemXsyPicJ9GELi2Hen3lLR5+i+2tVM7aAjBvSp4pMrGjFD3du
9uN2uGkadt43ehfO2bpyCUbzb2iiK9bHS59s//XScmSQa6tyfCqKiI9YtCRGbUEt
2AieUCIfoB4Xft1NxFhN8d4rTFXWXDT3pchvqV2R0ty1I+n8gvCooc4v4ZuNnbd4
NzJzU+gOuQwQb5BSdQcWcdK609vgZw0V41VI7EvuW0Wp1Uco/pAkc7BPPUvmGk/U
Ykiv0xFPEhIleTGlB4Wdeu8qkZEZkllHrqia5kCGImg1S7OQfe3hg73mpM/1uiAQ
HsA4Zf4cJqTJcxltqngj+/NpMpiTHM/af0v2qPaAvuw7Sa50jemsus8N+pQIvWSM
vkhAt3QuGMTfr5E8Ylzk94h4c2eO4JssV8NQ1fmqWw4=
`pragma protect end_protected
