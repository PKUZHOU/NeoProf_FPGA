// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
HNbzdsuSTxYEG6UzAVZxSi4IYy1HwhZTX3kDdrPZX0vgwiviFd6YB/4+bCV/iP6Z
uyZ+dcijDYsbnrn76FkaYNBo6tZKCxQNdOEdrqy/0+2i6QMfLrtuRWgnjE1vzVde
vuTaDoXWjZErYvv8rvSFSFGGMwIipUaaRKQn10yK9hZzepXbnkIKWw==
//pragma protect end_key_block
//pragma protect digest_block
OvhKNGiAx5BONP9FOVVJ2RcMPNs=
//pragma protect end_digest_block
//pragma protect data_block
lLzOfdOOvwP0t2++7pnz5cuA2NCt9St7Bv2vAXRZm4EUHF74eLjWjDpIPzH4R4Sb
gaFAdQJJeCdak5G3DuvPPHNqHgOr4rwXbwXvlO3Sl+e2CpxahF+j8+fPGR8rg7WJ
xkC6KLFBXVFAe8haLlU2BfnFUKk7k/9BKkhu1FvN+XjQWtAOsO2KrNaQUZJ3gNWI
Y/Fx9r86W+yumPb7drklWJm2B/sLZ/jOQ34sFyEkPZ0CKM0NavFqgMJvBRZv4DZq
KQ29IRcW5KXWvubqt6D8dlhDnNU3vJq+ONhkyfW4tf0S1VRs2AKVzJECyP7elSKz
PWxX7iOnjY3O3+ptPTT02vv48c4JhHMTX3+dg0cJ2QZU+oqgThJS1bi2ODT4K16x
SJOipKa0osR6QkGE2Gdy2HYiLw/jcFjh+yZX+gnnP9Tfk76Zns/W0mUc81hz2Ll4
N+EHlZl6sNGstJkGNDUL++3VX/9hS0Le/40KaR4GtNzQPf4l1eSYWDykL6z8gnQ7
etW1+81Awxa35X1MZe0ACVE7PsUHr3w/oI+SYy9hErfjrLVCmDrnUVV5wNuuloiB
mXgWhYkiNXPKnlZ+1kEsOL8Z7KB7zywQQ20Q61L54IYThSHf1ZwuSHq4JTjFB+wR
YSwgKAid8EAGndZhrJPRxzo0MoHuh62p0NF2w+nMNs83NXIbAzPWNXsclTKTyZZi
EGvB9Pt6CqiigNCsSNLqw1IL5KXCgYm+2BOCiRv5MdC2wDRBXm3bLNGeyeJe32fw
SGeRsPJxh1GyjBc7ALtPfCgdZcercjabcMGzxEvVJ2+lobzeWO5+KJrpebctfMbN
T3VHnho9ZD670Th4nuHngU4QLvICOTpa7m8vwMXmgeiev5tDFT5EoLU1A678GCK2
WnBjqynnv0UfqYXVR5olywaaLad3yCo99dSKcMp6yxycVczuWDZ0VDTnjtvJ3jta
0vSrslYrj+NeL1wXmcRvQj7TM0sWaCcHAX1U9MaO/d3cesj6gm7hApCZfu6DV6/s
eEuj7Y2Uo5sOXF99/Sa7slrcgj1Ns49wHOvwFFPva/PHP793LkYd0y6uWERF+PYa
OiIgGrLmwOf8N/729koD5+BQcGsGIrXzha8ZORfTVfjCcd428cJS9xmUm9a3coIQ
2CIBcKK5e9YfRebVM3vw2qDwTzAiQnxlck6hbed6iCkebZVTHCQr3AEqor1QQbw8
NvU2fh4vbzv/WBwUuOFbEmsasdy3PXnW2+Bt6rmjlxSMr5/eO8rM6R816/cR5jZ6
WmPgWheIvyqYlH4SuuqztA7EcJ2f3hXeMuHDIsAgBajk+08n89nreWB1SkCH6hf7
YEUhq061Th7AiXDZf038qQzVTXrM4cIoDUpGGpF13JIYm/BEo69KHfjkQfWvKwUH
LxNU1hKY6FbrckMAVSZMZw+mCKccBPbWU5i14AcL4ATVy2kJ06t1zxuB8P9WzNjY
AAu4OBs7AUU3WklCf+j6ZbN934oeARFykMROQ4U5PhlGlrn+kSRjAZWVVncqz1XF
L8nZajsb6AvjmyoKTqKlsii0DQEBHJRt+BB8s7Y9RQnmbSBhmx4HQO9DptCPtq7u
ZeMnYM0T6FX71JCEta1wgYijL9tozwJ/EUWpxw1zGT2KJ28yYAuwKe3Q3UIZ8zLq
H2mxDUEIN3Fv2olCTLK2Xv9DStgD9xqPP3SutKyM9VEa7wr1ZpbZTPe6qt3sdZt9
U+zMVM5RpThA/ATnxSiysV5jkx1bzcfc3KAVDnVZkgRRhhhDvJrWibmDs6VTLsK8
KXuplkAMHKfChItWsUnM74tANBy3K4F1FpcHVx+gXJ71Y2GJCSxl6kaqab32hnyn
CaOcJgLcbC3LxzzaRTAzJHlXNffaOtm3WnPvmKW7yo11YuHbGr2lPvEgODSAFyIT
aPqrCEIFkiEutmedkT7hJRXXLOd2dLgFnbWGmdnE0DgK1riFJA82SKFdPPtjoEvK
0BzibDMOadcEK9gyQgEHGYSjuAn/HY0l0s04yfd3RNsCbztEaQoFjAsi5QluaAz5
DXYe5EdXIIYPmZML8rHSXIbG4OPEJr6e43v7VEUgPaXbtWUitOQi7SPmlJ985Zrr
JvJAcb4ho+ccRIBbJY88ge6FPsc2lAiWvyQybUqJdDa+7D6/lv0bXDGE1mn8GFyZ
eYlS4e51U5ImPn+jnMQrlVDJ7QGngkk0AjlsLkxQ5T/vMG8JdCmg6V4VzZqByBgT
RM/zEVVhUD9UMQ/HUPkdLl2lKTnq/Nwh1ySZRKld1cuo8ZY+5JP22ZgJPgv+/m2R
KMznzPivmTxAk06zAKE5LKEbYje5GqI8FQZZ2ZjA/NadSViEyU3FRhGTqApej1k2
pbQqmE9lLA+iGgWFR8xFKKWJ9hQeMiWtEjSxKDFEAActsNpNhehEpgljdwKbK2Li
dPzAC81F8mHMs5X/htm++mBfPZTs28830ft81SW3oaHHDn8pOdybllyjy8+dKN60
nhScbZ7oMmaTPuoGvthhOrBP5gG9CctnJHwJVoZFaHZg1rUpjpiJF5CggJsxfLZO
YvzekJ9WeLMM++3M8LjJ+AzR3paLFj5WArlcovtMy21jlKcH6OWYYZGqXSOoFvvP
5CRQcNp2tz6cPSY6YlSrKdzQJLDA54dEi47ZNRY99b35IxPMw9puY1h8vcP0Z4iN
q0kXqZRT4ZJIN7L8lbA5YjXmZXWFJ8XGk86gqRc/RDmmETVL29At/5ycjHPqbfVu
0J3yvES+chZ/Rm01y384njjCUARaG95nmqgte5kR6juwfQsdPzNEgM+5vD8qlNoz
xkYP3LBG9rxKXCX3eQxcK1szIzFGSNnaUxNpUidcXyUKSfVGXyim//FMIxwb4dVf
Qx8rX824CKhX3wBotvCtnO4QIOH2pMG796116OcPkK86TxkAlrizsRgNrDXdMxR+
FFsChNn/U1CKXZG9Oxbqy9jOlHrikYlrw+mWd3biGDCygSJzlVC0fYg8q5U1lwZ9
bVa29gfjcBP0eUOx8Pjk9RfAuG/Q7qhM/nCI5Whpuq39SfWGU2OtLw5/e30WnRTf
dIc48d9A+i6yT9sEzS/9/aHNbj7R4L2Q/IEAC1zeeDxWDw+LRswf2+eYysm8dQor
JU+ZSLycmbGjfiG0CHWUCX58wyv1lqGbfv55CsPFgiB5Zf+D5zA0lJR+oET9rHVe
QrCIMi29gIAHnxRg2Fo1XI44Rf1uT4UWtihDIUUvhMqYK0hEdzyGO2zvsq7t96ec
cR6NqrRMET7LiD6fNYKKXzMUMdCtt5cXBta2H1v9feF1jvVkXTP5EQozE9Dc+8JA
7tZam+DmKotoMW+wfpmbAuq2V0o4ZBi/CMRHfcfaBzo7gKOijPuYvHbDWzMzgXJe
g9VToopne4oXx8owWpK3VpJ0h6rLF8iER+WNdZ8vkLEO8bpCysrPegioDSXl1mrm
eBSb90MKUk2wdONGqBk768TnYpepIXOtvP9jDo5aNikzrBZPjnWqoaYmLgKDLTxj
gWRIIRtsyTJfXdmV8B1gWAgVtfaGhNIIO9d54+W57YVdjkJRIiIyAaJL95Yv0Vap
AG7/DaRcXjolSv2rAjKqWl1r3mJ8ZitYMbO2c2g+XgeXWKS1Sg6hKBvgKHyY99Kf
jDHORypIzr3OFn80vBmWEAmbMQTCLbYDv/Rlq39Ug16xyJx56SIMxB+od4m53keq
gMWY3G0Q6HoXyGJsttJTICQAtiGqgK94ovN8ulZxSMYGVkKu0DyINDPFkohpCxAF
+k3tTGiPhAFfBQtK9AhkMviUAVcI/uCBJydDuv/kc5PH4oDPs15zGzG0nAahEQaa
t+QZQorxOdnZjnKQLwCcD4R4p0U6pRoRq8VXLvXSjJmQV4MuNcuZebiuGz9HowDP
mOu0EZNrY78j4Uix8fi2iCmywQ5NAMfTs9o6GrwxHO8Z7lMrT0LPu5lonenb+OqJ
Ye6kVhe1esm98VrfGo9zOXu7/NHxSnFMbKD8yv0q5NikEjsJZgzCNeTBdRWgv9iz
IYKdt1e5z4Efo8Q8b3M06ocmqO1Ifgqb88k9LzfysGjue3tCGaRWl/vTyJjeZ9Oz
9Vennnl3MuERrKgUueHRlNDuEMWR6uYtaS+6OBoOXvjnmNcIwbNpdFTwi7NjHqHV
DHo0u7pvcMQCeY+3eUACkLoHJLuBAZpcmU8ry4Jnc9rbvp7VRz3zsZpEdxcIS/E1
Bend0sMqkPWi6XBTX2T4TxKfQMDbq/jnuwlI19CdEJQ4E4oj/jV6vgktHJHuzadT
zrsVjfPsjkUhdU1AYeFh9gQ+7HqSLM9mVVnJKoYhc15vQaRFncPaY4j+zMTkhbu5
tnw3xZ+VBxJ14s+S2+44BYc89BZ3An+0J/zODs7JrCZsjbQdnb42p5cwro3IiJUt
JHSEao/v+EbOsJzCfcMZJZnq63K0C9kEOuZG3FNzVXxH17Ar3qxZbmlL/2RVGhRO
D81HfU+O4xMU0N0ZCVSwZw82yodXwViY4/saW/vyEHeQcqe76mt+dqO2j5tgXvY0
llCLOhnzZ7/XbvFuY0cohdX4XBZQpwN1MfBfRlyQJtNFLgUXW8fNaQBIBqyvLorP
EgR8y2Jy3L7gX9SSmpicklzXAikRM49eUd3uscfrwUzw08ACLytqDmim+FHeC2uu
aICKWvHjqWXVqavG46vZg8jOh0RfKs94XKyS43uFp/ng3SpsSxGBtuLDsMGa3FO/
bl22f/zfJmO9Xl3Q7jQpAx/SjyW76IoONE7No1gE6z7vJn0V17n4F8Wjr10YBG2r
XwHe5zyQAjq54/Dog3OHR89Zsuxm1idIsO4MmKJXZb9Qy7CsKfhL1T49bt+SwEYi
Yk9QYiBaEL9k/0Wwoj6CViwXdflvg+D16FS/I5A48XfISF8hxM468wAmGmGWy27/
5nGh6D04lnMzFlhT5hTxKm+SIsoLEIXyjwYWM22UugBhnzVJvrLUVHNSdT1UBh/Q
5Xr4TMympuFRJZjBStoB+tZalKYiXqL1A1t+XwIjMSDZ7CLIyZK4Fz7q1Gk85roK
/p64HNWJYdouv/BX4uMOkqbAE5LdBrrlWn20yYfHOVMVKQcpVdPZQBQ3RAoFtWVb
+awacdEewGrGQstziYYS/cFHog7EpiDNNYOd5aV2BrRikKhAG8hhUaxXtd/8hz+K
B6vsilibVw4EvHDGGCiS8lrfmp/a9DtgxSmPD8gK5imqdkkk+Kq7Cyg/hbrZ2Pnv
l4Dj7K1IiE5VzqrQsi/cwWw3sBfS/JirOSLLXgjuwtZzuuXIoH2nZaYR9gvlT+r4
ndTS48vcIGpDKYY2UCNwDRvhs9qbfJ24i+/xnislIuJqc1HH4S0qdKgpUhNPBa1/
G9pVA/WLRT6gdRY/PsVTyHFoNk/DrBcD12kC5OS/sXFhaOqbVZcL1LJL95jO8ES9
4VIhhX2CFOCQZzjH0Uce9sQrXZBWmXbY0W7QrEc6a77dcR19TqBeSWJIq3prxOOH
tOCQnVvqjCAmBEbCMtOLPjia/NqE55J4RGWwxwZjwK2XsZgej6IQkiZpiDNbD9eh
h7JcxUPfAFfQWXvDB0kywCcDfGr74gnUBsvQ7DgYrvpq7mNla3FGcx8yn4k1ByTL
5ErI28oLL0RiJ5fVPJ2iiimtKHnttwhII8OED9FX/W/4U8nwW6kzUqeYVz/tjzYH
JXfg5b79mxqGaP4mFpBrt0IfegSHc6DbZ7Ak+PBnL5BQAYw1TqFzch/u1L8Kpr9F
mU5jMX/moA5QdcwqdregQjC8f13u27cR1L5kdy/8MCcMBQuTDrK5gqsEvIdPdlT1
jL8pvp9QoYhWSVHCa6hKEsUdWsgFjZjR+4WOnM0anTcQ6IL5ulIz5V+xOmgx6DBy
nGyl4iS+bYFCE0o1ahc75NBvoR5Eqpyxt4yfK0/26FYs3FzmfRywRmsSC/LVVTjn
G5VP5lFaHhsSLZ3l03LYxGVFSIcAawnh0QD0ivldq4SNWSNRo1Y1roEAvKFirPBS
QYdmwf1V3aD7/RRuFISu8tJmb+a3F6TPEWMN5wFfPo2BE7161wgZzV/bcTj/oAmq
YYp40IqkZCnfesuy5UTeJrx2G2FW3yp48q0AHb+GGi819VfLPx9KjJ7xykuCGWMg
rqZF2bAWlav2XIb2VRf0WRWeevEYdhzfgyHgVMUvU/KF62Ih0IiIaQUJHXHL800H
3hVYiXsE3Ychj8HgIS6yWgof/XQXIqMVkxqoHHk15MlcPsGTtzrnK27sk6bFfUoT
alnzky0aBDh1elUY6MsJ3N5nI/5fEGHpE/BmLAOKJOu3mewVSr+4UepqiP2x0PET
lDbbC39NGaUTbrVww2xRHL541Oktpo3rgDdhF3sDm6i0/ABEx7pW/JJVKF8HnSil
B+wxEW+JfALV56/FDzFUJKzBSVRbr9IUlcuWWkapswiKSbgVZdca2T/l41GR3mJG
1gCS5QW85ITeqtDT9qQRzCAYr9DYarmBwt+hhGoOXh6BzFttNYNEMs0W++fE96KN
TGRQ9C5STk2w2NiMUU6nj2m0GrPjct1fSLt7to1mCy56DDUqhbL0Iny+6aPpTP3C
y4cGIHqwNL08Rca1JDvq+vjJMo+Q8nnd8RHw27LZQHVkHsqZf5jVa3XsgIiHNC6f
r6HqHR0SYvXmntK4vUNff1iLqEwSlMSoG1Nls0i7ZPRk4l8PsM296zvUxDvB8LIM
RGu4nG7JgCcJ52yUroNnsFRy9bPLsvKg64M9i5aa8g9PZpi5Cv9LWzm9QAKuHX9M
znZSm4OVnJtbOlFjFMXSIigzdY5OPjvq7jq2UlfwUV8HESwmroA/fJ+CL3aBP7ST
nU66ImGukMxrdOL5yPOQoqatJopXGj6jBkonQcwnwlvlNjygV76zscpaPi92LQdF
vwisWYGT16SuNlHgCF30qwmJmQ+1Dt+MHFPvKUWJCbWMc/IVBogTybJStZ7sOahF
5JbEYz4qAqCkU7oazrqY9lRHc+aQ+Lsd3ka26uDQrUN6z8pWaidO2cj1/iAfh+yx
66qI2d06NuViXErHUVkESHUjil+Xa+28RU+1CUl8NnqIoUfmiUFanBRivDIEyj58
F6zYuJTUgJxA0Z/pTl7x+KUEVoa/zIacYfgiwBfb6j6MuIQfsSH30nAvYvaIMQU+
GnfY6AQ5HMfzEK/ZgOedbpSS8RERV8GkaFBzqG20NvSSym8ZqsoGBrjaev+U4hk5
nkUXp3jxGk/+jccPGm8AQ7Xqt8YroMs7GLqKHFlBIYLA/slm87VNEcGGLyVUKTa2
T1qI2qZqpWxK7JtYBEybbtgeGx6UFGIb+f4w2Jc7EWAR+S1hW5iWvAV0AIAnyPU0
P41lW6nYpSoYMkUdTaL8iPRSEpTl2M+s7PIePE8BUbeJOFhR7YoKZmdqzDWiKvwW
Bvp2Ow/82NvfFrDWWbjHlkORFMkjRmI3fgV+i9Ba8lARFgI9PIeaccwS5/cI/E3f
PBP9ZSMiAxn6AzGxp4O4NXbl2X/zRnjgLYnthwhlxravDHmkZpGNtxcteyjDBTdO
ER/uVlZgR9D/bKW1N63BtCztwykBj74CoO+y/C0Aj0wJQsk82Zu1Y5ZYFvbX06+l
UXrdRnOVoX/Uxh8qLNqa3OT2UTojXeiCdMLCMSEXFeat+av2ycyfLs3o2Hr/nX++
+tpFjGSJ38ZgpXxMMuel6bhNQrBLI8e2nqlRFv7Ur7xePa81Jj4eZ9wwB1ybg9LK
gTtz/cV7IRkA7JXmfnD88VPJXPjSBm8d85Et96WvOljjMO3YGfDCN5hIEvF+lAlH
vx8pc2LF9qG6s2tfq7b5BBW3SRT/XKxDJZfq0gsuWNrtHkgYqr5uaQ4TD/jFvy0z
+1aYcjZAcQspKEqZLYvhVEv757krAuQ0Gl8dqG63dQRPZqbG/5kDAC6id9MupxHQ
aVevuTgxlrF8zqzSLfRwtqcSrO60gwDL/HsEntDAIo9HB8qwHr6RkfTEg8q4/9WL
gd7ctNuJa7AlUXeVNoPDEP0ELrXgJgwTXzHep40HIEq71nmdCkquJEZTA4RxJe4r
AGpyh0e5hMbU6x+XDiYRC7+Q+RtzURb77tp/z8ErY5YR6K2WDC3q4z+FbFlNe+Vx
F2FxYLppP7guBpSjK7KE7CGao87p5NNYSwshfGkjA4wS1bHW/FRnIwIJ2mkYEywl
UNabWoCqKAmbO616WEH1pLWu/g2zPB6fwnxH6s49euA4azdZpm2EwT4NQZl02TfN
EJprfpv5HwlOXbvna4/YoX3HnFN6to5aDx/AD+UwNfZvbQnnXPd+iRKjJwNdW5kI
9Vnj8BhFdGaPfIqV9Mkttzlf34RYYusnqU2Pb7X02jdM/pF2P5GTRYQTu49RXYPW
lUbP8P84NFe+jydFeozi40xLf1R7gnlI/Cx16CBCsADX9KkAYP4kNZYnNEE9tfEP
0PxM8tvdD7+zugLlnTmV1Xr0I6DBsiQXUzc/uAbBLxO0zN1G36MLuFW0tkAaFHXT
A+cQpMplWDNFR7DArMyZXW7ykrkUVFUkxp9BTsZpyp5zVqZTecx6BfV0V+m0kfzI
JyMrGvn0rUnU0pyz+7UvNpo5Xwj7/fuydDXXLiRsM/EIpnJR8GWR+UF9/RtKUsd6
Jh60T7ZrOg84czqL/Yt3MmuWBULAQlJhCDmY4qUKVoRoapAv+zeX05rM/wkj/KTU
eo0xPA1DSuufsmOjpN7TTOe5hrPsDeqa6F53E88ybse5pIXS/Xl1SwCVHj8Re6Vk
P+R/BC/4CdaIgeSDijGTqq/CUrEKwQ5Ss6bZYGnQaemyCgLs4WRE6tVnj2RTXA5Z
8C98KaCehVk793fRUkbUglsPdqcJYeG1KHvG1Ya4pLUky3LXBdCNyvWqPKLbN7/O
yDQrsUphrwS0dTYZSEml1qLc4zrKPYiEg4SDh0SjmFQapF8npD/UqIXn9HWUGllL
4SXKDwFQBEwqdQilh7BXIumCH1ZcUdpRu5zaG+37oq1Vs4mA19+AbuRJ6dXpOU1Q
HaZlR/9dH0kjTzAIiLc2tOQGghC+E4BeMgp/aCliBLae3sUcuuYG/V7OivZTBt7o
wgkHYsK0lV/WzF2DtTF5a9J4Yaufh7jj8TOsNh0jxIktxR6smtx0eZmKshrQTU1i
nwkRK870kUh/Y+Zmj56n9eacNGxAwNFDNckPWg3uMNThIsE7rR05wq1xh4Xfw5td
6FlUM9QG2RQeUphYv6LpwiqsbL+1dRGi8PvPUNuB0kBx5mLjNe8+GxHV0iz6SsUq
/cit3CrobbENAmB9prP00QNjZVmUAQUiYTVDhnO5zINJ+n+B1c7PRuuw6GfRqFHg
hP1PZqDtwWtNa4uNrRw8CBOMOPZrCS3BOhZTjyRuXpOi2gqkCJps/l0ZyZMU4JMw
XYEjhm1HVYikdALLWknBZ6rMsfHVEMV4stAvMpRN0q9AEeZjhay9DmR3GDVJQI7z
TPiDt4pXKP6mdeOJefQhxBHOWthzLUc9YAnxePWB3Y31c7B3WaFgFnnAC15QaCyC
7EvKVwQX4bUUwYdAdA4pUggoOxLhauDrMugA79xLOlCtIkUH9rUqxTfeVkQIuKuj
cTLHBHdqq/urNmpQH4i+MR688rf/hEbDvaUosgAx00JuoBKBZJT/8jNOFB4Y1eVT
1C1xi7ED+ohWL51siLbl24dmwX2rZ0PTpL9dXLepzXQGoET3ItsKxPl03XsNNfkB
ydo5KoJ9QohFH1nYU4/LXc4F5rnOIMmZoIaT8598YbCKPtSGimCBgQERL6/+ba2V
rL48gpiFtTBrgWFDSSLaW+23rgJtKA1Kc996eJqfC0rAkUenAh8PPzWmFKOXzXoE
c5ewo7IHom0L07TV2sOj5Oo9GfrVESQDOTZhl5VKmhV2SKv3l8jIToCPLVtP1Lj+
FG0aw0MHBniRXw3/Eoj8FAW3TNVaz1WnerIhmoYLh005+W5l0rPVECVmO2H9pBBt
jub/6yXBjUn08O2YXikLeRyT9N+kjVoT+HVTYOS0DZSu5pz6idsDeQ1N3KAwIawB
u0oqFBe59nb3N226Ylcghk5aOKltKBN4XpXXIsD1e1zEbqwWUCNp021lE+u86V8w
p4NwC2SOOzoNHVFGAAS8CKk/PyECmbZxYm4d9soF3nAqRHhNdefdEcKJGHlXRInC
Du8nCeoDYgaU/5MB1m4ZtyfYI8aKyV4RgU/ICtprUZiMLwVKHVnnt5ldSNC+0I1T
u9XnNq5VaCyDdmjwb/3mtn2RJBa6q18H4gDLJRJhQs+K4Nsq0IZHVOZ3paWFcs2F
qslvRv8TRGk6hdhmIwl7vGmFoduAJpE0RC8kdTPZ18ukVwXI/YN2+WBZiDfhXb8P
1/hUWrpRKhHwbGHOq7/P8UAddWGdKmZ9n/5+aXevZP+2eCc3+wCD4PqFG/B8sLVy
Y7Gc5CSoUW1MPzv/+FokhAGWlyMByGs4hyHxM5HR6eg+7bFqM1oebJmQmhCvCcHS
o7yY/v8Oxr9FqLu6fKTU8PDTTnSeBkzNZbDvze02SnBeoH1u2Z+SFqwx8gsXaWcI
V6VzfTOTBoifKxZoUvzBN2sX5eC/Qi4hhgYye3Tw2mrsprNWoYSfIDrMLjuUdnIY
PEK+vzRmU5bPTwayta+3Jntu3gQ8y2xsxvvafLNkYtf32zC6jlRsVU99yqQv3t4Z
7Rpwx2wi24TYHqJv+rZdj4h5MhwO73OBryJwhw/MjN8gBqtOADecTHeLzWIXuENG
IZrsU0vbv0GW63/7Ub4wkh6IJHz8qlvoAfUyv5UQrUYlb6dXUVKjx1CtFAIIBFgf
9lhq/R5u1vedIjFXz8sCneFAqbi2pek0kKQrexGJdq03C04E0zbExgaRLKX9G3z/
ueEO0fk86ZJl3tVNLFLg7nnsNagEYjYuIDNZrZmvLdtU5kc2ZcZybq4haYHXjJHm
3o0Vy3v0TlsiFQ5sXRKZV3qgb6CHOu9KqnAqazVGbqTkwq53X+JnDJcGfCedV7/0
2iDaskO4MdO++p5wV2Ol0YAo6381zr39HlPoHZGaI3Ip2wcrGRaoSjUxmVpzvIFK
9nj0xY3QgcZ0+Duae/LU7whGTXmw7QvBaghbDD73JuZiP9FzDY71MO5kG5U7Dftz
zk0GXzGPiPuMkHahraxPHviIH+sZznD6H9+njzaGSpDdXG4wMXW1YGX1+2s9Lbav
lR8C8OUMG4ybeFaGL+QnQx7zmn95iHpKFrM9thGErqgiUjG+X+6R1KzRHm0+1sI9
dx9YFV3jUSo8nEntz3y7EpXOdgdl9I/8qZqc/o2mctR26TqmMcfQO9Ic+nXyCkCa
kAqf7k1bMNXAwmFTMMsf4Tm5BnHyff+/0fzuLsizYSjwKrpbyE+g1J/U6C45qDFs
lTSVdzrF8dxxySTxGuxBn2Ia5D5qJ+T2vyQHVidKuY8haroYl3b36IygEoZM9bTm
oMJcRaJepxGRYXZL3KkKkaqYHC0TeQ3u/9Ms3l4UBe+z/GTF83YeBPszBto1fp58
uIiBr2YxU56yM1pHqwmKG9n9gdX3JLEwCloLQkQNmi648apoZ9W+MaTGOIyuT747
nuF9N2JDOa+vwHTaNZ9WICEHjAuJINSA4fmgfafD8OK7hnJzuLHi5RH7SkJmaqkX
g2u8tYNMrG9US6z9TiakotxY6vqLMGFZPKEitQQOrPVca8lqkdXMsYOVZPVXIS+o
Tq5wY2ebW1rG1gSoP3cCJ5rPTSiIkG5bA5xFatL6TzVXLhi81VVsDkpQcJOtt1rI
5RDNXpud1Yl9YNpSUVhdCx8f6Bf9wVo6TaUpENYkvGgTp2+ZNruK38/VfzrNuysn

//pragma protect end_data_block
//pragma protect digest_block
G0e6nuWhcOTnX9lOgftmlqXbuGY=
//pragma protect end_digest_block
//pragma protect end_protected
