// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
yivGC56pmJtJqsna7SMgPVaTi0ZjOC2c3DRcxqZq2ChkWjSE/FwqBW5LF/8g
Hk1J2sIYaIXQt5JKGsEVy19tIwDgLRk5GwTm2QmpM3o2leHQm5UlPfcMhxwq
WkUr3wrYpaU7YGqWkQXCcJL4ke64O3ofLhO7XhI+EFQwQEuiY5yylCH2V6jv
h8udV066SHBPY2JlLPRLMiq5unyADESRAcv2GELx88ynGHeshfGv7skQGKfO
ybORrU6UMyuvafvoT/c4yy3613a4+eHOoLzuM5xwP4s2Pyny/6UHkAKpmorr
t/Sx4BLFugmKbmRP9FTJ4hCrcIRoROt4bKljDmjxOg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
UWKEplboidjgKZSVj7os5EAGRxsxsKCwfPma8jsDdYStuqjNgqFFX+ahiHoN
0MGyzq29qMGwr+0L85tkR6qMI7dYKf7hcM674yL7zUUfphK/aW75neZ1FH1e
ZXGYar2C4ccNUwKgtBLyrn5UFP1tsLYU6mVx8GpwrIx3Xy7yy6pKgOycVbd7
uETVv+ZuMsB264CYwnz5RhEcPG4d+o0bfnLUwpkx/3cc9JnrszRpTfqyhdPu
b+VjKTEYeOhmhKDh4HVBR3Ty5V30sGn6/VtaBerCrih+lojU90H5dIOBwg9A
f/jD0P9PKNTEZGSJdAwPCZvt2en4R//EWjjZHu4QKw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Tfjs66TEnD/zkwMTdT8Gfx46wBl4aOk/GuOP0q/Al1Hh5LyTL4r91CDr+N4b
ZuABCiOC/WLIIReYeC+Xi7nn+CZ6GLapRXWFBqw/Evq0APodQQi0rifNXsTH
zQtN5JLZivvGaXImc08c8Ca3eAzd0RkXxY8GAukylZY+PEikAm8OU1Gsuywn
vSk3wbH65jYSjnJaYUWQz1zzk9lSqmX6fKHLA2l6I8t9S81+PQUO+se/5k8L
dM2iZmR15I3zd85p+xKZMeE7125PFEA0oSvssz5odNXPGvoMtjjnjIULk7FP
GRixvYySRYM4jzfcUtD5z3jnLFaB0To/Ak/Nfzllvg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
MYYcZi98/9g/DmXiQsP1TQzdkjeZusKyHSebbSk+T1owuJjvidcHWOzBzYDQ
BUGOgQYKFIlUyzOl3C28KBty5/NAvi6V8knm2kzEUQcrZLcz0tfi079gimNI
QgYeSDLDGoaeuwKBVw8MUnX8eyrRH6IlCvcSpPWFfDtvIDt6AVI=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
eyzhVBVdj+UWNiaRFXMZ6KfxsuBqCyUgLP/eMDUNXVA9TUK8aTdPs97OJze1
81OWDePBz6pm0+hKBYqQkOV3OEjnVp5zm9ZIrUM5xoJ8LD/U5lHLADEMxQts
45mQVZjcK+jvoN8V0u/3dLtWUrMlvcFoRl+2uAikRLpR6eIFEWS6sTi+Esh+
idYhhRr71Yk7nd538g8Fv1M5FuGoLICHbH7HqcCathFn5rtZ6lfaEKrSg35B
yDtzJaEcxgIJnF4LGxP66IVIx0IpIImCKa3mEo2/nK3a0Auek+A32EhqMEGw
Bu0ISWFwYOUxcVcSpBO9SRdqikgnUtPeYFxN7nUy+uDf+n75vj7HcENMnLpx
/DV14SwzsDlwBWCUEITeNyOIb9b+0LGBGSqMsKFgEYKRdRXe7GGGa89cZVya
vrf+p+1Mw7v/QyYITe1R9+l41Q+/O/4emIugjobali2++2bdY6vaTsPdu219
KOnWC3/el0JG1/byuszBYR/KEVE6ld2X


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
UW7RZGSGM5WK7Os/ZtzeZVeLZVUzO+N385HA7ARpOzy1uADlyLO11Ued2vUp
RtOb79xJPRPKJouWkHnF0FbrDJQl6V3qJiZVosOG08ztqwNpWGhXct0Wjcp0
5WixsqPz5WOJJWWug/AS5oweaBOX0TcCmf9ngyUJ6OGcE1Vj5BY=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
XiNiZFzOJsZ+N7iAM2c4eVRLgIf+HSOaKor9Im8ixm2AZtAIn9B9vA3lmZ5o
ZA4iNyYS+7vn8Tq3ea+ntc8ZQAY+PHvNXL8aR70Fd6smb16U+K48bOXknEtI
kKcd7Sb0INzc78DGwGDERXLk8MCTE2GPgYJp5ngWXmvJj7wuTKU=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 8272)
`pragma protect data_block
HTc3daRzEYgPzUf8Nq9dEWDce6jsrKh45e5sgecjpSx/90gVUBA3IJ//Vv02
TOxyTes3BYeOO29W2xJ7pgBvW2OxGdYzmgg/oEvvVEJ4QQWm+YTRvlWdFU21
lQYNK8captsiZ1w8WkvKAaTWUiTYOJjTIZm/WECxeSiG31+LiZ5pPzTrx5m0
qCw1Kknfchy1bmuNBS6UId4/DabQbJ9fDgw9UXtj8UdQKeIsxEMTWKgNDELD
p4YlSCak5gK+tPAMRy0Rzy2vka1DGjEpFGGdZCIaAlYG4DC9CQyY3DW+Ih5R
Hfb1TgDrUwp58uUBW7EBxllIYcMBxuOIEXXQELL84maVO1y9DhhmRTOmOfvq
Oi8H+XieRkP6XeM3G7NTb9jV/D7pSACpCGL9n0pl6Uqpn1Xhn4Vj0UIxaBh3
73p+SlvSo9oeFq+aFHW6G5iPOA2HBJaqjzikUf2s6jbdLmV2h55pMm6QDzSX
CYoyj4xZgJ9HHX9esT/OvIzROCHRO0ceNQM3zetaSqtsFkU6huqmLnDHQ8Dn
MG4FPI+PzifTSs56KsmxzptmIHDQTu29vVLQ56yycVRsZXa/luYuRcutvYFv
Kpu90V0jSuc7xLpKEi3+n9z1RhHG17RWo80KxNraOaSJWdSP7gMzh09jbH8I
9AoX0FUKaQmBSa8DaZ+BGrKgOoXKqlu9YTtvZ9uXBxa+FqPbNB2jq3Qc0Eru
pRQN23PnzYDdVqrSzQMM4JjZdRf9seKRMBOR5HQYMZrVP7x2RG10fvpVE7QB
7TDXS576CthJtVz2QYO9SKZ6CSmwF8Jvi5oicvecOw/U1SDlb1sncaiSCXhJ
yhg0ezR2lbAcejCeP8t2OWMpBA8wmS5HvcW2zC8QFb7wqovbiAT1BHqKTNL2
sM/Hn3vJQ/d3zKSPBxriBTo5DjcugFJ8Tkp82McVTzUr7rqyCIbJ81TO9z6B
E6su20XHQeRmP9Jzy3LECfpq+BN+6cNG0zTarvtwTQIlKqEc6Y7aB36qCD1i
Uyo640xEXAX2aQCWlFfZEC0h7sfzMO4TZOj52mKTlklMt2N/qlU4ZrtSxBaO
ETP4dwHinRzrzv64IBFudSQx22z670ml/eguzH0S8sH4AiZ0eyB+ZOWJ/ERA
3GACYOEDQiAueXeeFZRbgwyYWxjge1M+N3i1/8lBMSWNr+gF9EabAE6GWds2
ETOGMHeioGiN9vDeIc6nSiKQD7ydgMosqWcbMQ7HK/bSBiiYbvvGSXw8mvSP
nTO5gKfG7pKMfDXFrda2jAzfBY7F5LNkXyzJLV65BXBj8u+MByXS836rLnky
hhUzRgOjqPLetG8YzA4xoBz3ew8lB9HYmpHoT/QJrT5MKAVcpuAXPncT6MOH
serbvLC/Jq80R6ZeH7GEJG4BUXiRHCOmlnXv51cVNzv5606KTzcr7/fNqkeT
rZan8c3eUdy4MBGy0C1EpPL1GPI/6KHf9A7JGr4dArvKCpg7pJOs6Wkzns/U
uc7DSCInsRoTsDfn/NKezrfdQkNmC7Jx+w0DocrkEdiPeK8FcYGtQPOkZm/s
j8dHw9mVdoLf37XPIZ0S1kwsu4ZPcG1K/dy64wXOxNX1ov3e4C3kXc7oCPk6
VLXT/BHK131eSI0lafecUxkXRzRLAgKcf5NfJgElUV65ojKV7mQBg2Qil4Zh
UPNntgSG4ak7ZwsTTtAQjZM6+hZqPQu+weIbxGTgmA4XSInjK9j8t8PcvuSM
KfbcFNl9+ywPRqor6/JRoq9FjF8lhV4lMYg9+YFDMRXokUZIsOuqDaAApHTv
9cSrSJoLrD9peN0ZAW/hCLDDAwUX+1ybEifPMZRDU9jFG8/oYzsKJeTZ0B+e
FjjJ/3do03iDm7JKitD+FE/GOJliRPP8f2DCzpSUigMzfAx7mypKZNNBHPl4
p/cCl0nzizHCGFZ43yyXdl8qyXuOMd4ido42ojZ+H7tf40Z8G+lum35RgDLz
/CSqGpAfO3duPySO4Vnspcwh6dto2EeIr6vQG4DfOOkeyXhOUdrji50qYE8J
fB3rhQ1AGAcsJ3jC6uImt6IAtyVZW0OqVAou1xMhzZ2+ZGK3TKgDrKrUOrQr
21DgoiWLS11CttnxPIg+1kCB48xKzdmF8zRU9RlQ9T0xWo0jv2+KM1yJNlOZ
w/a4liRgkUAytHu2bZjGFkfRL/052GXE3INLRtLQ+jGNhBKdPizDJROao5K7
W0ted4Lb9HgljE72XSMmEoOAYb53HsonZD41oCAkcv5wSC8iC5IwcE04c+xR
+FfkzG0X9FGhOmrnilC8CkTMp5caMlxukTtxK71X9OlXSCqQUS6iSwjDuLvs
Qa5QxbwfrENymfZQtn1ez+wfBTB7C6SphDLXZAvcr2kbiKyjIO37POAUIFhD
SXUJL6RL7fMPJe0Nzv/iUz0+Be7bR7LVWhcZ1gb4goSGd4ziACxvTGwyohwx
pB19Q553KOo6FKOFMEA+gR2bPOcwgMlMgy3h8Le650+j9Vy1yJ8mL0Y0oFBV
Ng3GLYfpnblW+f+9nCA8DUTdSR0TqCEl2L0Zfmf1sudxUaswNpcJ0rawEuoS
XTV2LY11bLOaQEyRPeGYUp+y46D+l9c9qFodVxgH6IecCxXpTnqj+3+G6Jlp
NuxJZlM+Jx/lcHXVI0A0Cwg2Qq5ip4EjZLNhT919gT3QSNFGsqCC9W0xWSQb
NE2Q/ExaN1fm1ICx20kJacUbLjT03J/yWSrM+PLSKBL00cEXvk54IfN75TbQ
/qMK9YwjsKGdwmqE2LunK5oD34Q2NX13/QwmVm+9uRxuIBl3ZROAP8G3v4Lw
q1UoVwgt65Nv8P0BBvOlWSbpJaGWSJp4rdb6unJh1wb8vuf3Pvqwg0NfI6mx
yibw68ComEpKM0KdzsjvoCBaleGfYBlDItl83g/WhYb/AV9Cp1sgdy+JM+zB
A1oothx9kGzS+MP7zLrN5a18b0K94x4KL+2qZKgFNbWme5v9XHLzaJ23sYO9
2CEDWSv/MWDB7rgYR9Yesx6dMv47/GrvlXT4Oz+eBPhCmLKR8Bbt7JY6edKW
46VUfNuxt77Mc5qIjLatlbkm/zp0Cbrq3J/H/x7Zka8kvpv/e2L13aH9z0Le
KUTC48vZx51HVQe3Dh2BKq1xhDdELfsD+2n3+5kXfaYqo2ebXxHNnTV/5vgI
Lcnk8I+XTdJeGI2Oi9TucujLEKhEH+8KJqhlw7g+B0+lTkUuFmU/DKsWqsUM
n0mzDMqf7wcD8kw13nRP/Uo4nav4uXE34axY8Es9yQ5JgJqMMitg3dTtjjbl
FYBxWYHF3K796W7T9vg3MR55UB90EYxuQNpYHg3iMMzBe9B67kUA3ItBVfU7
Vn87C/6KJV7b7KB6IyJrUYizpcRtkTa/yhKJbz79SFAQtrICzIIZLJ6AwLgJ
ukGrarkVtm6MngPoatjCbQx19UdO3mO9g6toaT/h+W0BygEUBCB1RQWkodpl
lSV8NDf8NuCPhRUZ7S/hX1qtKGt+of9eArG2Hin+p9EqYm63r3U1h25BchbM
sNJEhFKOBp6inXaC11tx447b8DAgvp7EQZNbV1M86oKWlZz+Kxr1SDwLNYr9
FjOp1r9osTcKUzEu692I+rvbIw0ksueK9t8fbIGo5mN4VLUxhSVsQYTFdUMo
KK1rixqAS/h2RN5gTKIJvmBdqq0G6c5Em6eWUnyfUG/v/AW+wPWOlmje5dd4
H8HKL+AEc8tAb7w6zpBG6F8msHVefKFDCaIGKGAFmMacLJEafOI4AKY1wOpi
IK3NNOgtF1SVKMybUCRGd48egQQ+5gFfp7/87ut/FWUSdxXHheGSl50A45xq
tU7wd+anEbTJj5K/EuYPrugzCDgLXD8NBa2VXAYBeiMqMqrL5WxP6AkFX/GP
ZJHCYoMXL8i+MJagWuUVVBrrQHi1iUqBdTVa075Bc5J0p8bv18A40c9tv/Ny
MAbQoCj1u5LrXKCwzGMbWYKDOr5A7JGpCKHK3bqw3MpTe2fxeEuy/yVwzTXA
Ly3iX5YhwGLS5zaT/a53VkiCcYoPutl+n/c7meitq9wmu6sxnbbNTGTKWbgE
3FjpRhSI04mpL+R5XoXEyvBdY34WPJSpWhB8n+nWlpxNGsVaYhUxDi8gZUjR
kLiI7eiABsAJbqyNdMoqmcdkSN3PDYKwsnCOmfW6EEMEIBeyrz6DDtDNrmAy
wSRBgvO2Ux+82+9jYPKskn9yiXHRKqfe60AddsOH6AE6FGwiACkoVVVh6J+K
J4/eyy9xYq4o0B7sAintpKkB2Z64ZXK5Dn0f+prEPGR/VOnKV3QULuuEHErI
d828zUpewNlY4zy9Mkujs65cHZ8v/2ALABtWPOwhI59pMhm1J8WDCzBNkyKd
Uy18VM5kP9kf5PaSU/TOYX7ngkJV/aw7mqWmT6YXyuJPt3CROcbw0AQAsjmw
VQEoC87P3iL9ZxWXErqo8nfpCnAqPZN5gC2yOwha9YOOgovi4maekHxJuy1e
FCCuLy8NTaIwKnsOT8b1wiqMdC6ImjHfr1L+8BN+qCSuOcNXlg94RUChlOxW
sx+GMY89QrxPS8c/jg0EKcz8KgMltc8tXvkRa3OYi6/O75ENkLGggfQ9L+z5
QPmuft4/JuXkzOnQy/97Dvtsr7l+F195iEY60yEQ2uxxGEDrguy0Xcm3DwgU
OUIF9U9OObCt8mt/bVMp6gxSm6t0HWoXbrSJI2Qv8CXGBKrRa0K1ykwTIpm2
QYBVBL2L/Mlwf6rTFtc6SZ5qo1V4DKQlJDGbCjeHI/MvTtspOngznxy0ZaOd
fwX5S/bKLshR3ISao2POm6jeCNBId6fKjBhOmbtiybol73XN5pfXZz9zp62e
Vmu8qolILAsqoyjEYq5Kb6qoGgWqPO9+KSd8WMS4VHrKy5OV4qzW2+3ceumV
Iplw1P6joV1pYwGnYxh8gdGMPbrfcr2JGyEunLOglp3fBqkS6yz9OPuCZuMr
UNFYDgYwJySO2YOOEZGUEIC39SeiHH6USz/V9oAgH1uFHCeNeRIGxEbfWDxI
oTT7XhKUR9tJjo0O4VmeC04pYqIVEDtY5OuNhUuf9RQBOd66tTIJLXYVbjkA
KwaXLOYGjLysXgNx8fRIv+so78/8J/Rxl/isw3kAKYBFkXS9wqsVOY0JhYIH
v5D39dFO0zJCY9JXXVw11ZDx1NH3hdp3MFma8gPLoYRmpYT0rc6xfFD7/P5N
DEvQ2ymkA9JfxxYK2YDN4S1SymgdWRiAAJAE0eqPc19zl1TZqoyWJjvddkNE
7TQvyAyo8E8a1X67hz7YAO+SkKBY+6qimMCtkwz+w4JN6tSxNjr1gbDrH6Zs
FjpG9O29qq69h7Id0UOT6EDlzdfcUZ7IgBumnfUhREOHP3hZW27kNQ+B6UyL
SW/Aw0QJCazRIlTIppDv7XRhn0tIISS5ZnwWKrxYyoNJ3FHLzXvfClskT3f7
cr+SjcXLr9zMdDS7FqKHRmGgUEjQO+CLO653BIUjuHuJHBYGBXA5gI+rtjci
sN+WQUbPvV4qWFfjnfiAFA003rJAN3YJnmtnvRPyiheUjsQwo3TG/HgIIUis
eStHJE0CG8NlvVTxmpUD0tDPxlE5QVLxO5oBA15IFGtQO+xj9TS6s9D63meW
edDqH3riV23KPQpRDQHOAGSSds/LDlkeZERTqda+PZcVvVRRaLnprMqYkTv2
yul1mSDv6/9xvpuXqGBllVzSeWb+2FNqLA1rnq7rfM2TU9LJ49OWziAR7dfE
+3L9EU15Bd7XraTrDLXj4Q06o44v/jSFkW8SMuJ6qW8RjV4ArCIigI6wn+dp
PuSumMoYisYl1+hILMuGa7zoR0ivrafuNfjHVQpgg7Ec9RkCTIU6cyXolqAP
qozUZnXNqljh7TLqiv5jxdpfIVjPbltRY/Nuabu2MfMBubnD/NkADYQZVpm3
UFMUSMQm8XF2RHLATrda8zKLQejiw5l9ZgrJdX1EZ98rbt+x7t/NWbDqVbQ5
dQZQmJy5ByJPhH2pKfxRnyVYPEmusgk4DOh9KRW/J1hUepO5joFGrxy32pUe
ka4FkQ4J3hrsOZYbR7UMpFtODH+QWiJZtvzozuw9apZ7oogi6EnYWjJ1hb8I
r3X+jhOj5/JdYhAA/l8bX4B/odWGgBQjdvQUi3tIIAXDFrvuaFlVIbBC/vto
4qT6MkhivxZp16LDD5XWuDjoXkq+GxPiGGZAWa/tgkKCcChSlZe1ZKunja2O
mjb7jfng76GepIfjOO/Gn/k/mZEwReBn/Hdd6U+IF5krhHKpIU2Te1alQsEE
8WSYSaDFJKcpaO7Jfo8yj6COhtuFqdFJyJCI0Hl+kNXpHeg7jZFnJqGgtsw1
T+ifI9Bk/LWmTu2DP4x6IxnTrH2Hc8+hLkdBJxT2PUXEGzh6qi3FppQQnuok
6sOGA+NdY+XvYQLtu+G3JH4Kdti/QKQHiHz1RNjdhcztif3IO1n4vte1TpoB
IgrK+dsItx39+k6ClRN9FXPgOUMUYtTAHsao2XLEKpnAu5Sh8nmLwVwBQ72F
+XdCyBj3WoRGc9iQdTjP0AazmupB3uYGQh2C2oGlHXxc59Se7NEQR9aZKG6k
FSh1B6/hNack7+Ce7wwXey3s+/ioDAcsNvQZE5i+Ou/+tI6cTOHiUX8aRmW0
TPZdWpZpNwbqEonmTQqbJpfQbIgJGGUGPo4NNJvYauvWOhoclT2mIhHLoEbJ
yhEeD0N9ZOxPAbS0Vuk3DQrS+0fF22c1rrcW/y8vr/P6JiWfD2zigQt4S1TB
wZrseQcG1W4OgUbNjyiqXbUquqTWIXxbxjza1+e7Ja90KA6yk6ASbBHFNfWC
SSSQKutSDBBAwj2nwzAKLImVsGxDUNKhLEM+uwME4F3NPzp9AKe1tV4dx7bO
ZtydheQGZ+tl4/sPHF92o5iZdzMEz8WrO8HAC+AbB88EqFK9WHWNf8KsD44u
zojkLoqnMmkQiIRmFwmxzpsIPA5Sij2MSyf9UyZHRZBlIHsdRfbTpXuCx0rQ
FOXYM6i4+VotvFwh1DXdEGUj2qPeYOX078Nl6HFpzmelJKoDI/ffk+F1Mxj5
NtU7dVDkT1ecTr8dFGuqQWRcq0KBusESKaQSA3P6HwNm3GRH2fYlrZCcLipM
I4x4hAbqsuiz/rrYIE8bJFRNrC0JUCphMEraNEJluDQTbSfBjMrxqGXb7lx4
pfNrQlwbZbA/aO5IY7k4hiCNuuGiAWmtPeyCGq/r+qYB0ykm+4EZWrwKoUpO
XfP5t4aHyi552OfFYWUQsgfJgH8E1/tSSJ/fpUYqEJtrjEv+SKhsMaI9Y7y0
8tQiTMAJoXdYEpoqss42FMPxGEYg/67uEnsfFDzLCxZBl6MR7y1f5fJJf+lU
0t8++3p5MAKSmprQmZVN0E9H1svGmJ5dSOI3wn8SAYBQzLgW6N3N0dKMsedM
OsNwEj0S7o6ATI68fHQyeCCuta/NdKU7liol4CBwaEyBEMh1fRiDRSh3sjA0
deG0nPl/nxRnnFE6nbAWz+npT/iEAW2yMNirkvWN2NeZI78ittqo5lQY6biy
ZwOLrfASBFwukkCFYsj6QUNwFk1JNOt2pfjf/g9W1RB0oYe9Au7KwlhHzCDe
iWI48Lu2TNbjLQepc0sQ4Z6ffQjeggm0kYgM6n4UXIyrN2BBzcYnL1CowBFV
d73QIN6ltrsSqhFOUt4r8FPkrqw4TvE0Z5pDhDImD8rdNLEgXu8txoMOuX0J
Ur+F/V+WjrqwZNIfLC1Qrzur1htzWCup9AdZ95EdHwn/nCeLcqMLAkKq7n2n
UicpnGDc15qWECvqxsawGt3k4nL7EcmIE2D6ZI5FcpGjfQh3mUXs0aTq+cEZ
ZPbQcmNAocopdkS0Z2j9U5m8H1/gyvpjJrCf08fxQ8Q6AJGq+1sSy9FIxb7K
yJ+LdX+fjb6IbAaqG3t4nmcbBP7H4EeRsRtdyuZak7zJeAAeWkXblNBOjEWC
sT2x65Zfxk+SJNVWTrLV48LM05L6XpiysafoYdg9IRByykD6JONLWXIyVgph
A89wv9rSdWe6WuAHa489jGDGbUbu5RkyQBNsET6hoHOlsKBv9oE1dS+ZOzd7
fEulYXwzICVKX8Fd8dWvv7ojtQOTji4wS6mAK1PXdfI3E26zP19W5vbTSNxq
uHliotUnwPgEnWoevOUyzmrRhiYpceAb1hPHStqn0e2VdO7WlPMvpr7tdfKZ
T9NA2HnmGJ8onhz5b6sCg0aD0bNQjqD7iErKfApH77n8jxXrfkHFUFDAaTxh
rTlIPZTM4ov0XrAHhyQsxWYup3qtxfugSvbVLUOxHsyuFiaQcshhG2HddIDH
S7a4eE9zzjbnjM8ZoRftRd6mODBZAvV0gr5fMj46n+mAloFMZ67tAMMO/7Sk
a6E27T5eOol0KUciITVKCrvKt9elabcADHtLr3pTu4Pkvz3+ny9O1LshLiSE
Qu/Bohg78U9R2XBeN42N35bKgvo4/+LCE2rDkCVAOTxr77ZnsJ/yRd1dwleS
brtZM+Lgz74dNzPeWD+UCBXcuVrU+wWx99VPw7I5BimEFs+9XGWwdGfuUc8z
vku5S6mF4JDc8d70bfq3tAlusvWE1QOhL5f3iAHPZMsuaufY0++gV9CWpHZa
1N6QW0BR+gGpXi6LoMdj5Q4EhHeW8UgMCHODnHI8Yc7e2CwjxKa0Lw/eJwyK
e/Bh2QLwFFawFsRr2HAkj7PDabjQIIhCABl4+9PgRQ2vbM326pzn+X42r6Pv
agLptgk/lxaqZu3rEDz4HZL3cZe2krHu9bPbB55jfr6Ctk5RGFRJVl8WZK7b
sWMESlNfwneBcwbe7oNOb+Imv6q7uR6GntDoXPasO6j8tcJ9ehWEDTq6Zehf
o1mcKEiPTobI9Iosg/Im4t92AOoOLClr+RJ5J/TU3FrXEtx+jd0kO4FNX4bD
nqgVMnTTmO3IL362vxjLpAaaQcw/31qv6VXxzr9yy74uogY14YClv/YgDJhB
T7qsyInTUIiwOBMjaxisO4FcU8KR5hZfZPVBJFpEnS/oKTKFo5nfwOeT/CbN
jvS7bEencq5Qk45t8LEiQqpOzdWzwNd8Qhw95XmsK8g0HHDG4cP+yPxma9UN
ZOkD3Q1Irq46eILQElU1nsBgi0PSYInJ41v1ayqTzA91yX5AS8oUO6nbD/Li
LdN0Ht7HlRl5ExEb9aZDQzH0c7J4IZrk8frI3aTU08+WzNG2vhjF7Q6pHfdW
oQI9zmCxOJVAKdZuowAI9j6brGwpZulLgjE2x+i93CWs1DXSshCHPuTyBRyy
tQLM2dcMXKZZVdvxJJZs+nVSt0qes+pw/gjLDLtuRVQIaQhArpmL/EvyhiNS
cVVOPR7lAzKYojBiLUQpBx44UccDdw9DuIK1RDg0xzV2ZFTe3Uh1h/bGsCUg
+XILe18MTzlDgMvAWv+8KyCA3ipxAnqgn6AW32iGZCmPC8L2nO3NhIdt3F2D
euPojqOosBFgZGgACMTl7MrcfMBNeiWymXlzdwkwDJKClDdnkdrNn8fzyL7Q
FD69FZuBgDEb+T7aBlHf+kQeScij2CYF8h6Si2hc7zyB14pljW9K9uRfB2w/
UWa32V1L4Kv11NOKa5hTnlkXXYLTixfUbuzXpjAAkNc2hHeVRbLZnatm+s9Z
HReHLG1cJuYSLwKEPXtKLZGdqNU9wLLnMKq4FDqZM4BWFZCU9N/jKefupu/R
NNr7HtfAPKAcKnh7J4yGjtV/AUa2ioDGq2bnFtGrltO2qiPOmJ8R5671f7rg
L1erqK+tawslBKVoP0+X/eWX1oZHhlaLzeWKNEgv7qimhd+SifCB5+jkKZvm
aKrnIqotZhv5DjFveXczD4DN+kCWUONuZURxak5AlYCqXOZib2tGfvElucJd
LknrsP4fHffSOGIIk/0CiPEhW3FAWxlUuNK0F5WvZcDhPaFdQzT6GuLgRjJ2
BcXScazOB5YsA2CcvjZ37H0wXAyf642EXMvpQFkIC6onjv/pvTzRCUSQgwcE
Z4BDa4BGkoB6hAj2IEXxXWSRlN4K6FPU+MHep/bAFQiiODdBeml5rwN+COwE
XkJU+2t/4WlKWghITJLocav5AbGCR0P/bYk+6sNm27JgCcOTain47/d6f50E
wugLsCRhgRtopcfuRCUn8/wRvLkKm319HGI838943+DR8ApWEghMu1WyVCBe
VD737B13y6JC8nFzmFJhOLnh+PrOmFxVkXPWVA9TuKLmgFMNyze+5+Y6xikq
VtIaJwtvu+echskz98mM5JMDG2JGl2J61BP/9j5WghQ/0P03/HcQy3ezF39l
wJNUMEz/lnUwdARhkkX59ljQOS5/6SPRJClVnqUzcvnsxPJBUdNFY8HRM91f
hhEqzPtDRoxKetbPwlwkRntdUtXPqA7fCDl3v8CLsYQkebzbC5mOR0Wxb7k+
ojwGDQhdT4dxKTihrKCwD/Wc3Ohrvez+5rEtnbhjbJUqxNxzKskXVhZPyX0h
Mge1Skc/3pddntreuh8qJbGvn3lVco1n7HC+UsDs6gOGSrEo8wQ2909gwlbB
091NId1wXcadwL6x/ckzYasks9QQO8I0uwLMF5Rywd02GnBPSh38z94pLHT/
iaQXkJtpvZJnTrsfIuaACXTDJZS/DAN9vpimb4EGezWPuxfcrjsO06DIhDDy
e5PkDtINvi7NrjVLZ6Zm2iVluxLlQ4DBfUjo8XViDSK2/morhKlqY8bvyWWz
+T1MuYG1lDHr0R7qtmUq6GJ6ISgaVPerD7BwHBwCDa82tLXXa5JE7bsLN4uD
+/2wrg5NDivCTfwnz1Syoi6lU+rHzZotVy/DHQpHJaI4Z/OuAG3w2DImwGKh
TdZFMU+VWuRw0MuxY43FSCV2D/AIR19+Z8ct5OkvC00QyqB+PzY7xmncX8No
nctBxypV64spKYksQTMKyvaxked2x4QgoA+JJLZ8dB8cNSBj2uOkNWob3OBl
UcBf7VCc3o7b/X+TWWl7lecks+llaGqhyt3xv58N4e8sCmOLMw==

`pragma protect end_protected
