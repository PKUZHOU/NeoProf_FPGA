// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
am2Coy07Us6lvAU1RIko4uudO8Qfqc6igTruXMI8imn3GuclI3eq0YJiA0Cb9onT
qYAtZ/mE0P75CKEpiijsv00sNK2uetWyh4G3WJqCzkjAoSzlNsjJfLjkMzaNtHaE
YKIDaZjfQVxdotpoXWaTgNYWKx1ds1WLFtqi7CTG2eI=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 8544 )
`pragma protect data_block
fn5VIRWla6Q67cek3yLdbDW7COHalsCsM7TsYXWZnB+nNu9W9an6K6fVggvC+2SA
+Tlj5e1xXdXN7ur3Sigt+vBkI9WmQ7417p/JuqhsPJJCMgaXWgMJl5v0IyC/rqOf
PQDwXEq8sfHUjgNl72wBR9QHrDYnGxQ5Q22qba/Y6XZHYV9OkFKFfJalOAGhWhry
qsDH1VTKn7TD9S8zTuQ/c+SE1onTvOVHxfQHKDBuEe5HieZovk4BgBSHPAIoVf97
DuUqG7yGol0s/MkZ2aLAXDnkxuiCzAGaJ1QtISurGJFzB0ohQHuSRFYhAScGTxmJ
rLfJ0UkNwI89m1dw8KQR9YFqpDPM4wHpjnEb21snd/HBg0+6wuEwt3paDMRboclD
zmrxQ43ra+yDebUUVJGU1iaMbUks7DjE259uBpFvoNTzV6EFRnTPuuNlUh4ObliJ
jO7ju9t4z4iulzurWl/fJstIfR4BqCSr/PNRJj6R5mlk4Y2O9gdomqM2BGcA6hfF
/uOUbe76M0HgULrM/E5M1TDhABHNdMrHyaStVsYTCDW4gJT8ZsrQn0NQD8CUpSLY
nZG0uOQZd5Om2bju0ul/8H2Mrvw5s+V+I9Lwdaj7X+p0gVYCXPzPEMoPJgZ2PmCh
EpkAPOuMExmdy0qpN12ZOoqkSclf2ylxE2xAwGuLjyELd7km7eg0Hz3jQ8C0PwV8
zz3yDQWVoa79aU9i0xMS4AaHhDgjtGV0j/2OfNaC4aa/ib2DOsR3NkrY9SqfO7OF
dr3c+JIdFRQb24LVVMDoE8eCUpjsaOTHds8A/pJjy9OXKeg1Ciw/GF72fTEuCYQv
ScWTKV1bbGnI5RdDhkr+fvxCSphbAExC087GuFK+iN0jklPv2pPwE9HspQ00+k1E
zPtaqxgXddOyE3x4/KgxCQQXlWk1VM+J4u+q728+FpQOtIAjTQwPMgSuP25KHGLn
LU1EdDFYzhZ9dvSGYtYpOJxJY5N52Zui/NMai6nCAAm0Hz+yqWj9KSn8T6hLPKQ3
18wp5u0CWIwmsB8R1d8lxNKGlZE9ez3J6pv+uBFOxjOxC4eZdQwenyUzPPThDUdc
Wk/4wlpHLEX73rUWgRWeiDhwBoP5aLW23Z913as2+cJj/ISpsHGhhMAAStRdvoG6
M5g5Zwdce6lOLFoHiBcIVKL6j+M+IyqCHzi+TeTw8Rw1nrqqRDJVk6GU/uoxiSwt
MOvqi/LIvD3C8Tf4zzpvyF3+rIZT2u6vwTxbU3HSFFFikDlYeUmNXCf1fW+XFm83
YF5TceCCoVKhIEU4VZdIvx6uNeebuU41uOFTtEQ9tS9ozyD2CV5TbuU6gPSBx/Gm
enPo9muASz6dHzzZ4dNIUXsAKJVJZ7XM7XmZIh0kKTlJC8svF4tEALhcuheAgo13
YEhbhpDdEoi0PTbF2mB+pob47VILPMUflSMW8fbcLaa8i5g9aeP52ZjmU1XDwrzo
CC2R14j+lmM1040EmywXUBlJ0gzZop8z+6FGUU46zJeUVKWU17UtbhNQz6spQN3i
metTZ2WEWDB7gIBUY5dyJRVyqDN1wZdGbH2wtedVB1KYpgr3h6QJSx8RwDTp1/pm
NnKXgGbvgMLLjGCglVtDmzKyN9iXMvztHvJIP3xqNDPb4efGC7X1n+FQjP2NGrwe
4jmTclcDoxWYEkY1yk7VhpPkt5c9CuP825f5+Fs2u6tSy7IdDA2c9BHVsZBMPc8X
QUp3ZekzcjtostuR6NH0b/QFI8TlTiQaQWyQIqGvgbAqo5yGvS41AikwyJsLBiyK
R+bz2lIZ50LxypNI0Km6o2+um88sHkO7UD+u2BK1KLrsDqYZJ+3YlHYxHXoPf/Pz
hhY0cAmtII12CNNYh2Vfsh+7tXv/t5n3+aFNJad4488XTv1gZ2DXqb+LLEp4QHBg
qV7VnxzP5a+gX6JxQZegwn27rzErUUqNu7UAdhBfFKKxHuaMCMJ8PfXkIklA5OaK
kh+Ub5ij7NBPbmwMsOInlGUoipO5wtcyh6O3W+ATw0dmnIZSZab46jwIylhvKckZ
Uq29xyl5IxVdv+fvKl93VznCtW+YzjZIKwJSLmKriB8sxd50K2yAR+sxwwhwqSEg
VESDaxYU/VswPZmQMr0+rw1PP4Ig9AwTJJrO3g4AYeHDwpvMuQlQlQoK7yNFFOcT
byABsPtxvu0fRrdgPC/F9K0+94NZmL264kKEhxqxdv4NzxT4OHDOq9Sk1IZEnj0a
iSSmQSJK2tHcJ325UVM0FcSaGWBO9qgKURk6uP524JIxjcXNItH/Ui5ecELgV1c8
3nEi/9uSqyLdd/Uv70jYbumV0GI18K8ZVpwLbkaORVyR6C1c6+l41hxNMrVN9yBI
qRY1SwOFQ9Fq4e3N8PDeuy5lxo9vXDAKSrESNY4QbFhR4PFmI3c+61DQIod02urN
qFIOyuIZ+O4Xd1zON4ljxWwM+0zGksmAn7K0tN6TpsBeBs1FGlVfH5Cmw9ygjyKz
LBDqPpwgoWF4Kvj8GSLjOLI6G6U0PY/iS8Fbjs+bVaXNkPEmo/nsBQQ5Q2x4OtSG
KvPGfbcDcPbVWhHkzaaKSQ0RKqONIlBtnGB9syZXoRRK5XN0BheE+Gd6RLQzFum3
n6Yxe0G9AmjL23s/R59brT0Ujy072/mMbzK+rJjfIautmTwKUFrm29raWQR0wqxG
QTB4DRrZ9KZ4xllyoe1oeyi7PNXfQu7QolSdADZBw/Ke9IG1L/s4y2Ly6rQAmSax
5KRXB7/WRDyWJWorZjXTzKcmTutrQLr/dPAauX1rWd3XHHvXfd1R8sWqZ0Ht8nAa
EHF2/Cie+ilcdX2rbmfmZfltz3msCMZgP7856zeRw+OVQid1QxLecAfez46NfPN2
2bN3nOyQftI6nAVkaWZmsqa4iL3g8uPcsqMdWMT7cDKeBdUfTJTpM9ye2PBY4WUH
q+SUeaUTWfBDeF50jZ2p6xnZf+mnxRIrzkLS8bX2eFrU63csnh1gCdrc0ag9fYxE
DvEiVftWnU9dbjTDElxWoMptRnNaEpexsbH8uY+c8+V2EeCOTn27qJNsfPKy0MXc
XmYxNKRghDKLL08G1a+kQoRLazoUbdMQeXsiY1z7XHtaei4LTxgVDe9vTdmS+m9f
IQcDDXeNUDymDvXdxBMYYBKhfo/6DvzQuI/gGqislJW0kcYazykj/DTEuEjdKqVv
CGz568EolaLToHi8Ph6AdfHIxfdPEPN5khgT1dVWVHu5OvdD6yM4JThjAAjtLAkH
h51XyDWYXkCe0g+tjzhBk6vlTiJa6he5ZsC1Co7Xddei4M6OJA2BlaSBVsXICTcJ
N0CDD9KWGYvbdNxAdQk5zLNnWVdsOYo25+l9buskNZQalluIRz7slbqDfXT/YVrC
/uAt8kUPQwxoAEZKdgU+QZyTBN6fSNQE2ZhBuDjtRpEtEIB0E/ge0yiv5Cw1eXV2
zdC8vlc0lMGQalU+A9SXYNu98cwGvoOE3j2lfVX952p/WoY6XOTh0DJfLpExgVER
cN+jnI33S8jTo9ne5UxApUjY4KYsXBLVMg3RyLVaB6u61HKEX4fvjn9LGZaS7LiK
pgRRM/NFFkrqZD5M8ivrJDFouaonoXsNIr6kLr0jXyz916gTFPRT4K65t3oEcfRq
EYK+gmygNvSfBuN0AjjsKuh2MRL/9LzVee4YduRT1iemnqzeNmFXlq0DLOAjyKVL
y4aHjiqyA6oQpPZY2laBMiykHF6SYP2i6Aeuve81TzfYM7sU/PpV28dyUV9Qj5+W
C0gMRikfzKVQELo4+LlxHEiGIRmTnwWOaaOw5eqahii3FyFEU0sezCRfQJd+bM4t
FWxZMqSR08v8cQA7QknSUALuZw8IzEL1q/r3iXxDgqyViGp2H2+7ZM48JBfUxzXg
xhWGHtSwRZIa8TC79+bwXBGOAW1inx7F3OOYQoa6jd7pcaFJuK6PP9ZMdZ7Yif0u
SuI9+7iOtvm3hATyy2sdHDA3rappHRTERQUus4E1vdFa+ciA0UDKXH+lr+fMcMAl
J7GXuJ23jpL39lbjF1n3MPyoa3ZzjkFzUHXahqWJHxWGUV7D735Pp7zvIPRvphzD
9Dy1JeqUrp7C72LxusUx3Fe4cbIunYNfSTjymO4tOIYB78xAFMysAHMIzh/SUxoy
/M8kR5882bM/eB/r823M6auQWkb2hw/YXYoUY6FAJ5m+jUFrrNhqH8q2onuyqyFY
+4Q7MHC/mhRzr0Dn6NYb7VX4Ei64/uRpcgO8pZqZtPKca92x8EWb3y4XEnooKW8X
zTQCvgkZ0zF1UbVp9plL3RGWO6YDtxKJcGaXCPjXrzCybcNig9QpsQW79m2/9afE
lXX8ujQD4OpoE1qCy2JGTr1xVvqr4VZB8LOcvRZqlINLjHOx1FqEienHXHRaWApa
mOqdxsvXxcRxL/YaYpOeMfw+Wy7ApuFTAK5tpJMOHCVjgHN+U+b0n3VnGiEDe9lm
v5n25MCtXssZ69mKKulsv/m4kKn1jzT4AOB0ob3Fc7FTcbYqtdUNpIXZP7iWW3CS
1RaaebWgnKJpLbGcSLPXpXz3aCBkPNAWwt3JTZGaWFJ2/fP8sH+p8Sq3G/5sAxMR
/Ou/eh6QgNCGHVu78+qZ67nGpk5Ch4AlQ1Jx15UC5gxDbLz0/0K8nPac4otjf2dN
ySmif+qMh3+N+3Cv1B1uxLQ/s/PGmaYcKyeu1SZn9xGqtC1Z78NtYoDg578Rubro
3/BmoL9H4cVpHF3yfBDAwwyu7m7cuHPuBt86nDbDuak4paNfkYXIUH5FvT3ScyGT
UDIUwQSGuonddAKnJotLQYX4eOqpZonplovWaH6QUENFyEFVOnPvlF8dbKnuV9Zf
wgLzlC9psvqjRrLpKCf8AZ2Z6w+nHB1CUIc8S0+vEpNrmVqiWr4kvbKaT2fLsJ0A
mn6yN0627tU1SiafEZVnCwaRfnFRH/QN4Y1y25mFIh/CfZnSl9kEedlSy2jcrYOi
Msn+GxMOaER61y9jWHnprf1IIVCTjfb5fblPgd016owG7I2Dz/481lYHVcP0RdQi
3r69lIwzAHZ2fBr8ztyucyS8vSYQbtgkGP577bmeGuK5keDXINzU1QFkqnlAhyAX
FzlZkKmMVu0w16eL6QQGTU34v0oELCEofgej3URORF7s0+GfNo4HOLx8+wxmNKYG
yFWQgY3YxhgiWZz0XfjllGkpfieGqCQIYd0FhHfzo8R4AMQXy6zN7Md57S//jely
zm729pRE6DT9d2GEyLYLNQCgUk/PX2Cgk82zEFVMQ+vuV0rWvFD1XLnCIcXUOI5X
Tlv2LemtNyG1j+3IivIPi4w5KrxDiR4yYcEhGBqkXZGl6ESbbQyKyaq12E4wKrKl
Zq95B8OZ15pK5w0ryjE5Kv+CM7Fa2arqkl/fAGgdZBVc3XNM4g11PhxBgMeo3HAh
ng0X3MkTjM5Gl3AyT57qOmcdScoYz++5V3sP2TqSV+A2qEfZyp6dkTaI5HZf2cep
cT/KbIggsIZgLI053jP0Ly41V+TmwEGV2BuYHKQW93iR8+Yrxmlhibp0iwSIxXyu
xebnRdV15eX+Xr6+yNRBRPAdUMTSJHslQWh7f/2MmWStztL4t2MMUJjvlU/eRLAM
HqR+8QwnZ2fDBA5B8LkTq8CPXLI4rnsQzFy2E/TZzlFHqb6D3dKqDD8G923jHvAr
DXt0thqxFLYaf+Q1Ry1NCU6snHNJnDvkmYLR/ZDHxPK4ERtgUtKdPPB0LQUSi/z2
niDOkyHrHjiOhklfoTNQqxb/dUfGRnYOG3dcUxyuiVyPVd4CI6QUEAJrnOkvmhS7
un/tsmmhMxzXWBZOTD2ZOThov+Yxlts5q2bZ7V9gmLaVqrbH5xNylcdoE1lSXi7e
x6JNlgyb0qypwRJcnbDVdUMRZvYx/yuYjSjO9ePF4fnbijqb515fadwuWX7YslXQ
vZLqQLeLoY7iyek+7ZjnOZbqXlY27NTE0He4DP/TOLxe+7Jln8oGsMRpEytGWDjl
L6qImWsE0vfBYWlRVkvkhnv5YBVpXxLhVyAPsDfJI3CB3GJS1O212IiwHuzMr4vb
yK5wSlX29wqbvdDeybfnjn6dW0qykbYmGdWMRENei6TVTfI0hI3GNflWYbszcRl1
MOGdEFprAs7Bm7y2nPIkwPI0oxLj0Sje/9v9ftR1INsWUgNyVAsni8gXWeox+JAY
zrLgPIzKKRpXPNGao5DS+bRyRxHXYs4mCtmQwOfOeO2LeAl8e4ApqG9OZhdTNLhf
wJyRfp6XIGNoW8STR6ZootESOf2BpdwW5G/4pUsDl4x6WgamPJJK2jysbz8yIfmY
d334u7yynODi2byxVqJqZIqkum+0DK2xMiq0vPlD/F/bL7V+QXPu6JFvZOIniCq0
4akxn+azt9m1C7dEEw+GAJEUk16lDCtcYmACnrnH7GO3ADttP4f1Fxyhzg6JN1qV
k9ef0Ok9Mg4nUUsLX5Htkmj3UYC8g0LiUdWUT+d6AHCcPTjGmkiUNxATzNLia0S+
xcSRo+hS7649JSGX21vftOeFMLUsd/0PlZJEIrcmPrhwZhuXYM20sLJRGTWkAGAY
l/p0/QILXZG8TFSMp10XJOByQvmYhutJCrj1hLlEZSStdstM4Ib7wuosQPl8E8o4
5JnP9ISif8lc7Cy75nj0CsqpDbor0OlL+wgRDgyneIAZQIR2/5Cj7CPLtG6HC94L
zBe1OUHYx/LzUVpwr5pntArzEWuiyR1LeJzL+7a7yu8PvJKfYakfq+H3S8Q5d/Os
NBEdSHuCzvG9//cc+DqWU8Ifej42KXDzVrwlKQaSzoaaqcIAnl2wz8Z/Od4rfGYZ
MwnX5Ym+8PfoGI+Xg3IXmsALOqOgUZHM3ONh/1plrtc2ITvp5Ilm8ueIQbQ2r2bO
bKYCijrL3qRfxurDnpX4Bkv0SaGGhA42Ut+S537eJV/3Kb0ArGswLGzf0cKkuqzL
ipC9IfVAWlilhTYhC9GyuNwj31rrFj6OIg2PtHfMWmrok3XGTeL/VPaZxzMBmnOJ
CTpcCmITwDa5jPuRkMUsoDpjQ8Ns1AUwFv7ZFgDLgC7xDzUwveheToIErOiRKGCq
dHK4PExJf05HD0GrJMIWhHu50+eOw0DaVmQ/ReTvnSRKsayGBsi49PQqF2md8VDm
Ls8bp0a/br/tJC7AxVH+Rf19YnTAiWLWkIxfdTkDCMDJv+e9GbV4O6LW4JSdsnKJ
79Sn3ZsxX3rQV0AC5duQl5CHzIBdVrx5kl3H/p4Z5WuAdn5B9uKN57/hd1W1o2H/
5FpID/qKBnN9QjO319F7chPTdWLaMFgsJV+Q3EgQAfOJbI+PtmWp5TFkvAcDZ/MR
ec4yLHYvCi/VRckzy/mDd5odNiE5bIFYDc6UjWT8999x9v2I9RXRDmOw577iHmIa
tGpAd9tuiDEqsZ3oHkWh8w3BvmgPczA8Taqlexyelji6KAy+Azhi8UY2XciXxIRd
DU3LKQiKH0VzmOK4hJhqsjuvAT7tQXd0S17mrwbLOS8eaYwYazz/4Xu8DhtA6ZVo
ATwC6Lsh5rNcn2wH1Ef0SKhpMTZEeqIkCeI3lGWvnDo1l116GrjkVRwaHBrWd0QQ
iMBW+NADhKFk3og8G9EqI3fnlj0X+TRQPtqXeZsk5IUeWzrQHADnCrOZyFuVowvT
qZ86wTgfD4zkGsMUxk7Uu7/I9zV9fQd1fbltXRK6VYTnpe+Eh15GXNMPKe7YlGXv
LYevqmG2oPIEhd8ybYyGs6HxdNvHhmTP3g7V7jTk3uPRztox8jEuo+Oz80/AsMbN
/P4GfEh+6y+GRXku+Q9DA3ngqdE5lTI2fEa7vsES+lmrJeqhOvDXjY7MhrZbcqbD
eLl0qu7YXGQ3HDQ1qlRnVqHMrN7C5XlZTFdwo0C6ZxSx2K6If7kgjQII2ofRiRfi
RqOpDqkVmDiieaHOQmJ/vWVQ7Yay02PDvtu+HZTNlk30d82yxPpbXV1nQwDG0zYe
BD4jmng2F6fUKAxSCF51XDtLqDHL90x+0VCtdI57CHvKPTFFqcx/RGOMVU3nl6+L
9fFWd4Eza4P9bld0BkZBgZvSYYzfsvjaarkIVufrafKeLbMhsYMuAXEyemrv3D+d
xspW7ZB+UWW/QCMfRJUNRl7509oul6aW/JPAtDiNjR9v7Z8SZrruXh67XHylkdV+
LEGQy6YsPSTXnJEOjH2r5Wd7k2FmJI2Zc1yH8cr6yyF1s+dBBN2aUELAq4S3gQSh
IzpgLx42cc00zJ803La2xQyQ7engLPPFMatchlMhEy/S4vY7UFhFBD9xWJnOc53n
Svn+xKThHLxzWBWblAH9TUPJjUTJ8Rc6osGaNWMtclibjxpR2ct0+60iIHOg35EL
2lK9gW6u0qjmiheMEN+C0XQ3PBlNDoIJS3dCRpiviIa/cdN10jQSKOXzrAT0biIs
anKWIXoRSsvTc2lWX/yqK0lHt18RJF2T40r35UMsq8SpEHOf1YSBdjrckGbAtYCQ
CJMqmROB6p/vrP+qIfqGZjaBnnXmDrMzzY/AYgeW0ijgm2U0k9MVbaP2eN+HoaGJ
CRDUXfCEZcpEKwXzKMMwzL/4IsD5VD1LQwe9kJl2Cqmtu67EHoUszhJli/Mh/8N1
Zwm5RE1QIahACKh6vxOirvX7FEOD16uarWBCUP9GOwVKjQGqWx41tnsRCqUujipX
ExdEFCad+y5ojRpewzTkOQ12WrIphPQCfIvAQk66oavBCTk1S+oIpLE5F30lN3y+
ngyLHj58LyGnzDiYK5U+jHKJ7ie7OsKJ1DPIzi9fh7+Gu0+NQ4emWUazs3evf4tn
TBSN8UNVDbJpEOdXuzZj5HEsO1lYGWjFTuGzkVg3XO/+TsSRSif6wg1kk1ql/eIv
EUn803opWAI/ckv2YLZMD7S2iKzqcg4Pm6DiURo24ApGYNIgAYtQjVA3sFf5bl3N
Y14diJEIy6S0xFt67te1v3YHYxBL2Mmu0W7SWikpFfgvOZ1MfhBlsyCkIGynPA/2
5Sv7jFTLACJhur1QMsMJ78wt0XVNHNWNCbe3qJyaul9HZ9K47kC2BoEgJER57aHt
2+vd7sbKVVdaUULNSLwFEmNhpGnfukI6Tw9Qd161iynKhPi3rWNppoWXFQR1xnKR
PhGHVR0fqWndj/WLpQ+FOfg3eDPTpUasQKqaqiYo4lEpZtoHyjYdy15oxckJTKVj
Q/GsAudQe/rqBizEUJhaCkWt6RcRP68VVSV2aNmpJ+1+bIQd6T6VxbU7YAicvsSC
66QLUdZsO38KPi1F8XDGXG8KG9lPZuzgr7ywkaZ64uAzGjGttOLxi6fA+qh1FPtp
TK140+QPtFQ903MylDB3PAuZ3G2AP8nW191emds1MbTkQgF24J9j6IfV4/FKCLuZ
BqNLepobhm31FLrNjxgAXIMYcQnXcKKnd3tApZo8FkOfn67G2jRAEGZRT/esOCHn
BY2+tlfyFxysyPQ0HMnnZxVyqTgymBFO33gS9+Ru9vGckL1FHIaO1XXS65dFs1HX
e5Gx4Agj/EASbRXCb3KwmFKThPz68MIv9V5Q+IPaRWM60iMiaAEh9DWvfoyYe/h8
6KkX99RmIs/s3gIMEabf3iwmNHLSsj1Hry22nqDMYl8ezeOz9h5LLeLghxTYhWbz
d6u7uz32PcMgPWw+7iZYkyy0mvPl3262JDTa5MGDnsmnv1rru5Vjf08RKE1YSQzA
EtJSQ6eaUEDkBFlPjZtHSMhqe41cdWVgUpb+aO/vguFEaZoHVo19VTDlashYW+jf
8k0JTNPjYXB5pW+NsxCt6ZmHhWyBO52nkRvd7p5Yb1vUZK+qD8G8fiFLK4uXuu81
EwMnUa//iZdxRNMXB48Jt1n9ukxrPsQi7otnlEslmdO+R3XX6OF1G/uXIGSIssdv
kBAKuQaD0qeTXRhE0G2XjthFsBFe/fwmeDQkHiSPkvzZ1Hb+yPdMzwUMMRQTK313
VZOPI3heV9JgmBg6eRt/57QyshMJYgE8ohAQiqF54GEkK7NnmykslV6n9G/5qvOg
UahQIu6Yfx+4tTjldi8InLaATB4pvx7dqFV4kYdy6zy0ULyLjJqqluPTXXxgLF3Y
cOog3JHinSsDqUwNhmqVsnmlScZRiQ61sTXkpo2LnX8EkUlJ99XQ7zwE4aX20U2S
u6CyKUHPEUNjNM85zC6yuXOxLu4sPuviA+UuDg2LLRTtTgtwdkPtOWaSwAYQ57zM
mnMA/8+L/RbYkQwO2EaSW8yAKm8R0SKAnXDCXJ9gdYmyMgGxgjMrPlym0HGWx+/9
pM9YjJfqhY2JFa4FxRk2MLWNSQKsi6OqR+ZfvABOEqLg9AnGgOM6GrnWgg/sdW9D
Y4vesvdx9QZ8cHZheG3f0sLlQt1KXID6khb1j+KgHD0iCCWYrs4Yj8wN8mMw74Cg
KVDGcT7FDXFM490wmOIYNX8YvWjOkB+iO87tZdqhbbt++3EdFlDRZrDZaSmCVYCh
unu0yXn315fPslph2XIwSXSltVl9p7YBhZlz6byO5LHvXwm4llCH+7FPa5MrNIvp
fWdNt+0LSWv2CH9BS9CI3ejkXooD4Sh9z9MdYPrWaDg59rqJOzB3JN20q9KAaAT1
3pb7m6bd2McPXPugE89Nh2lq4aCLWpoluyrFDbceH3gZlAYnwKFe8E3jZvwOgBae
bdEX/e2+vaBXUdMLZOfVbsdYnRtVHHzay+5fy8HXSzajIVLtW7N6RTzBWXz1lDWl
cDSX4Oq3ZwqbSsV2BC6uPOc0FafKiLe92SOSaz8KvzEF87QJyuyEH/gWpWROYhJO
3U61Yl4dVkq+Lkbc/qA5QQyN0Q4gVt+mY3OZzd2vXqa1zcYQfOS7QfdFVPuN9NpH
Jd69IRDqxdvWFw7PS6ucnFbe/eLzG0MbMNxlQsFxfu2+Bv6fOT3XjKU7HXKgz/uA
H6q3DXeSIVxOLG7iRaulJ3VA2p5QWjbZU7Sy42fe3IjNQ0ICnoXpk9SwWn1/XyFd
V4M/iPYK1d35xkbDK86lRxib4qT56NG+rlgzZ4qmB/vRoF7DJazQ+7xQzmiA8sl8
Y7fHSQDTbgPuexj+2Cy1kfqh3NjdR8p6hHSQW5UqS+eq5n23DjM1UPfCmfsidA8a
Si3+HslMMdsfVziKJHCVWzTk6lUUyFBDK+1urFiXn+y6d1HkYC36OgGgVbkXVH0G
/S2UX9pw8hyzWe+ofzKGrzQNRyhE0ZkGe0BZ8bx2NT3GILR5Dvpg//ZrPUOOYJ0Q
9X9ZmDNqulcvqQBziIZDeDRAoyaAARaanOxOUMjkax9y+ZtuMtlqSY82VdvMJGNl
muqqzWyg6kydBKvo1TWfvGEE5eScZpZfn6QNEadPSD3NSIdl1tlfvIiQmy9ygJ5J

`pragma protect end_protected
