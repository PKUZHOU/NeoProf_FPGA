// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
AVV7H5IVR6fmPcN4Lxb0tsX8RxaTlhlxLlbbKgcJpa6XcX569IcBeZ5cvYcb
tv3Wvi5h2cLRDXjPq/hyKQbgUXVO/ePXL//cyyrQwwtkxD3MwWvFemCVAsNv
sAHZwKJDtzKS9hyt56hP96udzQvRkOzy2v6IB5hosqv8ocMt79pkC2/e3+KC
1y9NxS7dVQf8y1GZsE5tqV9VXGPuw//cn1oxWSRPkwn9Up+bM+n+1Cbs6gDh
abjgUm7uJVxJYNf5r+hjGKHONKoAXCqmreFwwRsJqalf1lNWWtvhjUcWbQaR
AucSQyDOYhofJ9Df/tpx3aHQkVsQWdfXi9ZPmfgiwA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
i0Yjb+BQxlv1QtsuIw+n/adl54xbeDLsNmI6O69sDijQlJmqyUjgQl8lb1H5
JSkgStTzFkdRFfeaB5dYa4HWaWEOYQ5VaA977n4ira4zQtEYaIEw4HDb8xvu
fO2u5FqiffMbsJGWcIOBmj+3VgeLMgpqvbNL3Hp75GseQzylfI090FctWRtO
S5jBiEbrXA4bOt181DQS3469LOuTBB7VNNFwJ+EQThSqU10HsmPZn0/otLd8
OD1WizHTmnFPvmor5l58T/Tut7WMfJClu2q2cxoidyTM1oVYUB9PQ/dCKjbW
BofnC8hIiXl+1lFJ3FR0k20P1kVchN1rMnZQYExkkw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
pwQz0JQzTu/WIAtDFyIcv2G8AMfVdRJf2bFKXSw+9IrH7wMvQlAAeEgNnkx/
J9uqBTOOJnoK9uhxBIH5xPh1rwK5GQ/hDQX+S+i4NvI7dKA1GbK8O8Bv9tSz
Dr4Be730O3T7uTmh5qMQPE3WPw1PMgkowhz6rfa+wRAJKyeyOeuit8aQp3/R
/TjX0+cVh7zHtBG6DjsCExCkaZEXCQKACLAyvwubRQsQwkdx8CcHeJMrqfQH
lVhJMIqXgiKS7z6sak79qbzq0tZEYqc6OR8c80Iz3HYRuN9jixCYYL+/XjBq
qL+yrOu5g3M/7ZoQ15Rn4rz+SqA+/g9K+Q9ubrG26w==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
dna2z6i8xbOOeQLPsx48Xx9TUgIZRzrroO/MrpIKd4jNFnRKnXPTwdKS6F6y
wGnAl59BxW4G3nC5QjJex2keQG/eZ4VCZGKFmQtobXc9rqGdXUG070G1WX5e
3agL/flZfckvJm7pdCw7LB9xrxJBboopkDrTY4TF3ys5G8369qE=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
YTgorO8TS971VeiNN9jOsK7eGqEPndxIET/wN75MIO/x8qiy3DIAjNOojFea
Zwt9fPH5Yt+YzUWB+JzdvUC3iW2lWTm/SMHjvLpuaagxaUny2V8edHy80eDq
LqFUUK5JK25hyeCf+MMdeQLdlbANKIlzrvKuw5MIHx2S/cQ+TKn10V848m/j
1pHxy0PIICBw4anuTF9AW2/xtCipUWV/xj0OebOvuSBMwYmJSh7JJjAT/3pP
PtoUKqmTe38ohmJ5nMAir8vsQBKIEhZAlrokjZeBh/0vEIqI3496TIdsjjEa
12GSoQFV35ek/iHc1U9ZWNAG4vF/ndcVW8LK+aKDE2xuhxMwbSy63RXxnnGW
WQ2URVmK7z7JGCmE1PmOMYthm22KTyeiW86pV16Ql2kHZcMT7cqT/7nSTfQD
HX4/Y161hNIZnLNpD2ftplzSpfV9z2Gpd4wlBajAICjmu7bwIxPDTwC7wRaB
2NFWME+fzjFEaG7OPKjhaTJhqr9EubBM


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
CUNSH3KjzxIiPgkxuzT3T080/Mg9R9NZqC777Q2ROXG7yIzqbvXJkkJcrccp
Jaizl5l/Mug3FPyeoUNh2ghqaGcS4dZJFJ1/dayzSxGdWyT1duq5KsE2Zvc3
XxVO6iOaHfmqti47kxEZWk8MrS33vp/ZbKax6nlzl8s0PsPGKKA=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
a2vNF6wqAp/+GxqLlSOTxnrImSkv0+MimOfFdnB4f1MywpPV17+HRmAczvQJ
T5sFKmZbOouW+FsQkCQa/LMnWdcxQCzxrmHQDBUkpXI+xAAfXUu4a0FHbrDJ
HHlqeeShf+lvkWioS0Gkb4Qc5Oplu1cEv3P14VF0NPUCoHoVpEY=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 16880)
`pragma protect data_block
x8/G26mewGyXaSyMtJWPDnvfwxP0xVsQa1wCk7DNf+GYda7Vyz/mSi8LheQW
L8V5yTvMGk4fxXju8YP8MVZeo6TdF8OrPqp6I8unkMZ+/z/lhf2B1WTdsij8
b0Ctw6iqShdeJyEMYHnd0Q84qTfXgPyDkg6qN/rcAfO83UpgkXOEURzQnxb8
+xziMPh/WoRpWpU4Dter/bUbtVrvlInT8eoq1s9nMBhQBnfGrf8xj0qW0NSb
YRWC9MapCvtilMrCppGig+SNe0FfQZ+o/CgGNoRTQzVFveLSDEDcR6DKk4dW
F9r8rJq9rl1nchwoaWxIbJbKkmggo71RIuZz2gNmgkGc4U61hAtI3G04q5F4
3HHmxSo0s9+FyV/vc+HwQmqgHT36fPUNSwzHbDDtK//yL6E7HoznNxhpNoDk
2AqSGBA6FfgQtlF2VYqLBwQflolZr54yzyuubaiaQzx0jFgd5EotZ1PcB/zA
lRoc1FE8BLBoWo4sBnnQBnfAVbxI1Mf4+VmZKozj9SblJQ84IE3iopvaZf2p
VEyJBDVomT/dC8RaRzpxdHEkYAUbbZGNx9pPfBsV19LvHIG9SmsB3OecR94P
isKcT8hL1Np20ec1TTzD2AjcBnZ+ib/jHJmgg6LTdQpMZn3psAgc47kFdkhS
t1/bBqKSYzOaAxRF0Vm5Ryh1ot86EN7RkeCK1h+9eV6Uwmjj1b2rCsHZ4T/n
3fEZLbAjmXaTljqKI4JWTgcR3ksSUKUfIU8Ji8TDbfGnqjM8DtSBfvN+JGyJ
Vi/CJFS/3yL0ZoszSdJUhw/4CuVRItS9gaEjQEgZsaB7iDTRnv5jC5OJy0ZX
gzc93JLAGAvTA7grgpqHOewJ35tDXdMrLic+r3dPF+WkZn2DFEyFFonos6jp
CIkZVzRxxyksappJLMhnXhz+2xAlb/+/KIjeWOKS5MFJ4E7U6yujwNTmHAMX
fxQCiok8bxq7YeM+OzMFOcLh51FaXBqXhiGvWPxjjOdX914ZHXSZXNLspUKl
NaXa4+c50IlIP/y/SsChoNQFCAWN8XweK2WDmPkze7wRdBalB97kRLdzYYZF
ErjMmJj/Erqrx+QTMzkviA+sNxfEMVn4rY0N+jYTcVtwNvI+2Dd3VHV3K6fI
TAfiPO5IOX+R2tBVECisBK3FAnP5l6OZ6zRLuz8Cjf27rzFzbeoXy/f0jtCD
4GeX7iVl/rOakLTcLFVvuXtfB5JSE+PD/MS9ALpOhwVDA1AJd7TVcyR29gP0
jBJ3tS/ikMS26KnAwQDjkkjwJwRMPGd/LfmHlCskI8YKqctHEIEPTo9YIqb0
bFEOUnB8qftNsQOP4qnslkBv83aIiqT8/7YrOIAOztTTBPtnTN9jRT6BVCCz
uQjaJT9egV3SzvxQOpZnGOs3pQT/DCOJ5BvuAC29ob90tCRj3LDtM7wjaibV
EvRfWcaAaN5OWUV0dS+k0iIW+5v5c8bQDBTuZzGUrUuIM/I0cv0FeaLwM5/B
67X1TgenHgmPKTzjUwJtYkyVfBUKcFw/QUR20D2Kyy/6z/TRuGLEUP35aJ1/
uu302+ILj7Ks/2mCV16d7majCPg+co9Wxxkm4xHmv9ZnyMJ0Cjt3WMU465EX
epmc0o1Q3O63fb11qYgYobPJiixH1WAVVRUljDJphg/dIeztZ4x2R2Fli07x
YchieYRgzDQ6y59Ss6J6eeYGaq/9JrufRgVvBI1dJfLmvJohHjZTtR5nQJ0s
uYJy86nEFMesHXfnJ6pF4ZLzh0/yAPzJqt5q2qkbEplJIywHxrLaMwhvO1Zl
zuOMRDYeC/58qOluanrgXyIcIvfvIzpUDQFrHNpzNz1KnIRtxbnYRIQ6tDqU
ZlpXybwW88iJ0J9g3B/UfZixuGYeN2vSw3C9ANrHWHZgGzcJFxTL+BQLANdM
LpK3AylggMqpdZWqg69zrSDiVVsqwl34pt6MKRndWSBpQ+/LYRH6vm7mGVT1
EQbtdf//Z/Iy6Al3kM2qwLftZbRKDQ/SBWe9g0HsLzrI6uPrR8MpN9lQGCaT
g0/gWGba3w9Af7fcwqHB7sRFZq2PZCWgKzh8xzPoaTc7VoqD7yOe72DKPr5l
rQRMF7C5A4XZpCRU/TwPGHxE6tEGMcATzRJCzd7y7WbD4CcYiTN0gLezjRm0
0gOCsUGZmkB+a7SL3yU8OcTTRCOdSeuWX/QTHhIXz5JGbzPjS33NVBO9HkUg
HJYH/1tKoIfavQEyDQ+DOjMvomMbe5SaZVcGZS5xoNJVon1jxTFPTn0xkqdQ
XJEmu98z/MKiRQ2PaEW3KhWRd0NQduCWa+Jb9wU4Wc5ZjW62P5Vskhqg0LoW
YLF2rinYGv9R1RM4sIym6p821IuoehQeByrkQGGmYa8JAQJBKfJRWehbPIFM
IOxbIpCZfyoqClsqMtlcA0zhxOE0AdhxCI90MMalLu52BhwxgMzSsPODJEwj
Xik6ZPrGDKI5op/QL7Kdmi6ovXftE485Glv5ctIauRRg+qX2ch2e6AE1MMEO
vx8Zvl/bEmgxk3Kp4obGrrgYBqS62Yy4iA7diq85BGf7xJ8LpekFGKBENihQ
xfV/R1QDIWHvn56p1U4TPAWv275gxVwzdI6HijpBUhYq3a3eJtY36eziScCe
/ZyLSpJ66OluekQydHK6hrFPvb6KQtwhg4Iy/tzPJ3NMkSoLVs+dUwp6LLXn
DzFC4UIL/ue4IEKMRJ6DPElHfN80pGcxCWJrMAIGmV0cr14kKDdBmk6Ctwcq
IwrjaOJknN/KsCU3/Np6oRIQWiFKjT1bPuhHd+XxBG6PTo7V7CPePiIaT4X6
vnwyVyli2gcW6wOi3QhDF4+W9o89Hs8AAX9Bh7DJLZNXOjrrXISCbYAr97h4
/jpZ47sHjleY2BCwhyD4FYftpkCNoUlsvwt79dSywjiz4G1sQFCGuQaWQYvJ
qM/SlSTh9arvaL1jGfB8bV/ShM7nOrNhqp0oqY1CNWtN5l+/pPmGuG52txzo
GB5u633HynVWF1hE21o69/l7ZSXnnWJHlZxK7P23j01Hylb+W+bAOUUJqdwC
QhO9ieRTxwJXM8PPBEClb4qLGe0RQ2U5SS7q78YabpTEbqIiPgAMICVac3yr
3YGCIUm2jOE5n5gnuCVgBWkj3k/9EuU3lusk9qUrNxWVaXgB5IfQd31r2oVO
Ll6tWKv3TKQH7CW2++BGpFAgoU5362MVgcCoPaeYCIaQMl81YNxB7WbAD1iS
aQN8W5mis3JzPpLwAnQ4kx0oeEAOIqxr22dCBpKU05qVVh//Cb6oMJKz0RUg
mlDkkSD+dgr+06YdES9DKdlbVq7sLOKDcDxeLIFhsXTN0epHAGkbRsy22jrr
N+sZitaeAkyiNiG1Kif7fAsV5N/LLYtkXHlTyfIczq7NXgIpcV5+ACTwfMAF
itEZGGbGK48vPkGfi+a1l6rEQQq7EU5qgOFVlG5BsMLJhgA2ZgpHT4lDcP0q
g/rmhVanbyfIfRYUSTrP+qllxGXk1M25tagstwJBgPOb5LjPu/ma7iU4ZnWk
BEXDg6Ae9BpyWFx3OYE8Fecla/nIZKZXgNqzJUjThXIRLf0IOfNfPfLBAZ0z
SypHqjzRsVTH2GThu+41s17rGvfuW3gmnWcR7ZNNM++RxMgQ+bGpJ2HTqshM
AZkbDEjDJQA8O+FIpKC/CbpyCmPVBEnkH2lUhJawBoE+LCgoOKIjsaJicN3A
BuCLrSwKRHBDZU/xWIg+vjifYyexSKNxMGFlYReLQqt+VNWZ4bQKLCUMqGW7
g6TkXl68qdgswKWBYFx4z4u9R2pLBRZxUrHv5B9mkOhsTeMr7BMaKFdOrqav
CmE0ELM1e6Soq1sNEzfts/fUfY71/ZRYByWw1IP9081fT/hnY9RJaMeUFRdL
F89TcFBpGAA0dtJB0oUFGMBDmNX/utwNL1phmvYDTi+I/gotGyq+4T11Teiz
b9qWGIfMr2wWOTxNsP5qFvwTecVbTJHcPX8y9ZnejARrIjBxsIf3VYT2V9hQ
2Vfq/yOf+2yW6+10LTgpdftrG8nK1a7x0MhesO4Mrl3E4VtfdSa8zHYVvRic
USfzxh4kZAyykKEeTHye87wijgzEEWvx3ah+7fgrNWpfKDu2udD3qEFagJVU
YEV2A07jIgC/K39OSvqIlaq7QoqbxQJN5qc0NGbB1n0UXtZyJr2hYDnz8mU+
gwyYyltqMHmftni5ko73C904F10L9iFoQoe+9pqQw3D9RBRbPoOKrvLC1Sgy
kNUJQxuKwm+mUaovA49OV8SPrjqby6ioS+eGF8R3HZoGJwXMJ7hAe2nWfbCA
K4AE9WqQcrBPadrRTmSgm1fHTEFaemzVVC55btp+WecDphoKOve8+MnoCfWJ
gCVe0yyw/Bx6wIxYvVdHmBVCmbwtGO40njF7OLg/h7i56YaHFZ/Mb1ivTzC0
THMw/L3zKIREVNohIcV84BBgDUVlV6ItAE8mVLZ+Ys4EyAiFIpU8f5XIeziT
xvnFGAhkFdrxg6ul3bQBOcdvGrLw0LmvQPGwJYECzseRJRY0iH5GcY/yeZYw
cNy3AlXE9geJusWFBR/QTWiNyF6OfDh9bha+lbpJPBUIEyoGXQu1hRf3jfF4
/cq/5Nm0Rt5UVC9sa4mwitbYZUKVtxIh6BxFtCJ936eRn+qZ1K8uHWkJci3Y
A03aTgkayuq08rZ1bIVOBiVzDey3kITR5ZfBGpHNUwt9/eOmb2/xxy8ZGRwT
Ll6E3gYoyI6pLW5dyMkiL2l2JQcUfgdR334zizInjqg/Dpc/dWlTgANPPO+x
DoDMP/x8WGZHi1X68ZeeNYNKyZjVJuszLynb05nyDtxmmmKX+4sF/bri9loh
JVXLww6pGJAd+hIaRyRcW5vvh1MkJOYwTM+oPRumJbzcZ3XrHCkG3dCM8TzI
9XiFEgs7xnv2bybqjM7fRKrA7LhpslDq+u2E1M7e0zHT2Vw5cV++WPHGL/dR
WV85Dr56GlchabLxzeq2IvRIj4pWG0KY/JCDMZaO6qVmfxM4Ofumlun/SEn/
UWzVvYL9g/Ns4jH6pPmGrjS8kywlhvBo45UzvTJr7TVdRPf9GWWxZGNVRJwL
1SPEf1vbQuEppzhohqOqVHj/SUS/mXWZAeW7/PsLTTEl0qZVR2aidaOs42nB
xVQsz1FNwVfTZDBFfiWdUyfWiY0byRJ8p2uSz2x/6bifDGkUPF6UeBCKi+va
6OMt3kgUtFAKq7TQrPY5bwNv+/ui/okuYy6pBAydTsAf14ngwcO/+8aH1tZn
Ae8zuuW1IA0Xk+x6uEgyK+AX1ih1TiD25Koah1LHCw0WcHLhFph2acFP72sG
qCxxU3qxblntRoag/DFMCKog6dOBm2RIbOeZkLCyyE87TsHYBuSdTOrLb8GI
k7XLz42qIqwdDlcBSbFuAqs+cwupwzfPq29OkY/hgKiZ7Azu7aat62d0HTff
4DFkHL+WdOd3ZKKc5lnt20wHiT0N24JjlKOFBWs+hSzUVCJN9HMXOvACXKVe
aNwqcJ7XfEObUIsr4RtKVGQpm/B6j1rLNxVxfiYNAFs8H0PNEOiLJV8vT6jW
v7fP0REcE2pZVcDkRnS3wHow3z/0KGUXUvrTv+4a/YEX6+hTX15/Q/rrEP0l
MHjSrusPDmh4ObHMFSXo5b033QVUgN5c2Lu0AToZZo1ivhRbuX2LSrt0CK8r
X8W8qknqFx1wgrlWy3ruf6MIkYuVGzDgOQR7o1q3tkEYp6hnEmUng2iNCTuS
X20vwFXG+I/Es5G9SdzlH7299HDaciNxEGX8f5cnYfOGypbq/scU11LcVJCE
0MN7XY8WeJEw6qmpal0yJnewpFU7YSzO7NENBayHt/MIaJOpCrq47ce2M57R
MRNun82awASo2Y8sPd+ENAs3pcW9ZT2PdGsA2kn7XwoM/r/9Lgghot8YO9qp
jO9FKVyaUZpgoxczmshoRQq20nSjLC3CSh/mU1FW23qJfA+BN/MIzLbNtkGv
rCJedgcAgdKxcr6ofQ1btuFjD9BMbba+hvH31vLSloDkgtzYwirXdbFayRuf
65dEIH1rplE0A3DuW/gqmHHk8u9i7vn6Ttla5WMJmWts/dMkvx/MwynJcnbR
Er141QMm3FEPRrtMshDdaP3tb16H/CWc9omcAQuyFeEWUUwDEQA+OvwwpeYg
seubm0cz2nYkDGis7/QBLBhe3aWFEBM0IBdKgCYNc4iTRUcISR2C4FF6sF3J
VG7PEuVOjeJR9b68Zl9YO2ezYcBUiE6RdZAr7vKrfX9kWp7bXnG66PBbSmvg
uLV5HH7845gQawO6HMjx9bwiwhdJyYjh/QtgTsc4q6XXmueSnBicHDC9ZsoS
F0c6z19JkC5xxPxtwz1ymNlaQKRmz6HSa16rsEiaEYGl1wBvLw3ZOgd79nQq
uiOW02V2jjmasjmUgeqWBn1HVY8KrxVkOxuDA+VqXWsAUmYbp8za4uYGJLvk
Ng7RdSv9Qhgd/kHnehg8kElwkf59M1MSXa3qQk7z3qiXjGqLD0l5yGcPDibt
37166Jhqi7uTjsm1VoFTlIe6PiPqjzXPyL0KqmWJZMHcq+Jd9lyPe3Trj+IA
Kn7/omrA1z7mrLsdWUJbYpeQECbvUuj9M3nPJTMsMZe92zK8ab8DlO69qban
8hH06iszFyMnHsJfWxh5cIoPsFRwZrk/cAxiEqJL9sP8AbV5RvIuaBIgDShY
9OA9VVH0dVFt+QDy0fL4xC5qj0P8QVFPWtiAxOU4DjNIQQmJS6fhsvzEl9Oc
5T0sA0XuQO1P3ZM4m+qmbPg1lu/MhKlRwkIzFoUnxhiukPpkLtKRBOfo/LMB
kSkhSnwOTInyRmL3VoZtSVFYC3lAnkSqVX7jIvKmS1BHt4sCXr8pg3X8trnk
UuJQd8z7QsSx5doypv6s3ZOTKAz/0oLvDdb9fIPzQtS7UeMrDKOvZV6Uf3Z5
vb7kIdnwvsc5h4ieNvOREllgz+hhaMvW9zS+MSEdRplukl5UlaOZWLEKUmnO
3Rtn7VYLono6lt5sEl75rW7+apeHTu/tAYaeq+kc7mfoorZVqBuCeSu6E0p0
EbNuEXiCSB2obcw31fOlewpaMx91hIikN1ybHZfE6CTBK66vL3tVX1O8K8oP
3Urqx1Q3R354ixMvZdbVCtBeJuhjRbIA2t0jTD5hixdadGVCo8IODT8mQyrw
tDAFhGty/DGNsOZrnJrY58LrTWIedI2fojb3yU46ALyrF9gQjjaBolpClT0R
v582MLMoZIaVsj0XvTMqNESjlFU7YJDD4VuZ6PVtNKTb4VXMyv96Ng5iSkZg
jPHic0lfUQ5HCWouWCW/xU6Zcvlbe/GneHW6eTc2YDalti394qzq4Vg+uB3/
D5nkA5F3Y0shT7LYy3ISV3nfjnrFxWRt7oHdvxL+WVzsSIb1tlbSAPy3USN7
7sz9/o5VN3smt6qI8kAfQs1r8XH4LKxLh42c6rSBL4xf7N956YA9GPqufNTb
BUJp0AOcP4CuwynErY2sC9KdbyaBCwNhdol5xiKXwNRZk2AFQrhx7CZyQfOL
qHi9oeIaC5d9CLMDJDtnG3IFhgqNKgAQ+4Pa3Z/66iMOhe0sLzRUgTZxrxro
V9kx1OXsDlzZ/+ca2nv8Vb44UFGU+zqsFciW5lgGunzvCkF3ICYz3gUFtFKI
plbUftTS5kBKmRTLxRc1S/pjQeyYG+B1dBl0s3LhF2J7BQ24KstqnfWsgGm/
x1uLFp4Hf2hKTUFalCeDmIM9w42Ln18uaH4E4DL/t7Q06EJXIbfcdr0xvl3a
0u0skrUEVi4UTxROOUaQy1Mq7Rh8JZbictPswmVwg1q4Gkq4n32jaktp0rVp
BNrVnsBxqmmZAD7c6JF3qBImMxcN0Kg3Hai9AoKeut52SkwRVJNnR+yb7LXA
meAuSHCAIJpunJAwH+ZzI7T5rOEo7CO0AAwv9CfkCkYKIhGAzS1VNdxC2RNy
Z/cd5w/UhwXCQ4/8nlyUMg9R4AGrA7ESKulM9BwL6Bw6tHRpfBVvtfikb0cs
PSWAeA3jnJkUlu4C2QvmTO9Uw/4GBPyS7kbTJyudDboBDceaRyvsnH0BM+/q
EDxC7NmgRH07nhZWC+WqD/TmNTsxtIcyx9fDM0L49aGCUmqfc5LNVYJ7UuCQ
MdxFUugvJDbHPmnABmGw+oRgcNLlpiPsRyk8xJFlxYAZlgPlchDADy2jms50
s3jFwzFCnWEjREme2KHWG8r7CO03vnzu2VX5rRzJLpRLTax3HY9WsBptIfpK
+pln4npUYZfGlw9yiHyre3WIjpLgiNf4DJo6guP0yljKeo78qjIzPxrbr097
IrC7z6eXT4SGOhO5Cl/hJBrXkf2OYSL10MRJwe2hmyYXx6cA7VhgLdJih8di
myzScVQ9b4DDVimQQW68ViM/bnsIvHhXcekLn+0a3Ig+UO3OnJshUCgIKaMT
G0Hfb6MfVYlJoXK8c9C+ejnO4m9mk1JrYs4OhbOChoTL8Zqk6NS0X1lc/XLy
Jp878u2CitwP44IvPO5hurbxuj5l9m9eUkRqDyMLT0r5NSSo0TIaY120u2tQ
yymAyCizHgSGIsKJgAE3AOaLan0e5injfYe/UQA9Usdo5ibk6VQqdxTV/Y1A
BqnINfXr6ocV77kBcBcVxpSkuWT/86lwn8V7cS0o3yYS2Y037z4vjvtteud0
lDUu14woXydEaTHX5YWUCY/GmiS4l3B/CyUuhjS/P6JQrm79KID5MOwlLec6
6/KoYyjHk8PTexLBZQKchB14pWG8jFRJ9C7zOLzzU07qWPViLgmQTvgqrsSU
HKeOcr4CA3+x9PPWI7xqK7AqbthKI0VyvmmME8BiVUX6jT7mYlpaKFxqNaLD
QYVl2UNHjWk9p4ux4wdX/jjSS1/WiXbpRoCPHcgKAPY63QGdvxJPGDFrwRLy
OjRoLmDU4e1XZYRVbEIqzosnsL2rLYy6tPfl1G9lHzi5bkMaJDgVfOfa2AUR
lsGQ6LBgjWTvaLFICXFM6yHd1Bnd1hCseJXu7Wq4j4pG09xANNqok0JPaZqY
1XMlJRrnBPaltKqS3AXKknneFF3FTKTCIGnaMzpdE2mofK6ChX9PrcoMT6j6
9aU/K5VH2wIMSEQluGgxHlGgT/3ErZr7TIn1wMpvVj5llEAq32yvVOievH9q
7gzoukzZPz5AQLBY2KN/sPJbjYORrUqmKOhDKPP+wSP8cYrCTJGjG/qK9Lqj
QbPFOvoIZyABbOHWAXhNSvuk7/06c31tBL55Y6agDOzEmalxpfYEp/S/1r0H
VklkSUwwN/0JJVlzIzs3QQKXhIOQF19+Ax+voeb5puMJsnC3V9hnC0TXfqvz
A0jivT6e2IZsWcTeiYdWQ/Ed82dWMJ0sqglbWrAQucJizsKVDAQSVsUYBTpB
nlSlqyiC0BP4EcE/BStQFQ10x5u8vLxZeeipMUVfTmqGl17/OG2f2cTrhKXB
XKBko4iGnEURUBOgLwKt/UoVODV9pUiRfhyU2z6V6wdFzqC3M3Y6cDK1Y6VV
th1AggxFds+82BWqfazIlHtbrNb3ReLFDWan3hoEwYZLdB5AyJZ8XQ5s7N3O
GguSTp72hjtzkS+KzziFmz2yCyTrm/hwAns/h8/WPqJDYOpZEdbU3i11wDnn
IDve39dQPoAEKDG9FqBKLgjKr3tPPE3aAGo6xBe9LevlEZyVScbiUMiQYam+
WnytNbIJsbRba+DQS6PZol56FLku9rodoLwYOZZm98113569v1T26X/8kWA0
bk/LXL3cHSGAuE2KV31Bl7kCGfUnBu43BNiD2HzkUZ2O/ABHalcAo4i7GDsY
aLIw2pKLvPqK/v4edG5B5HEl768ykbpjOkIt4dQCZ9cU0Duj/0KwCx6g4/qK
p2SWMuwc2fKuKC5/UPmcvDT0Cav18j1DGr8IdrORLkTd99TVxNZtfTb+pZOf
55H7IXHC7boB78C9RtA+5v35mCALooxDcHJAVFOArsIoBgZ+UpNinR7RW7UO
+IfNHpY1Thk18gsBN1pPrtImQRh2OhFDxIwxrQRhh+5tvSIOJCB4d5ce+imb
DKH6D5WEyHQGRzGkFthmHXrx/otuQgvMFeezdHYI/avI7e+GsBiQT5U55Cw9
SwR/kpPnbdfgkTPw355Ya8NVL/xYHNFmi/ofSJF5U69BGLphI7kOw2hghuCH
vuLZPQ4cYLtkMsUNVL/a0tw4HCuywaLjvHxULdxH87JzBIlzyAvPKoh4+wxD
z1sNaspP7mFt0E1a5M6nKdNNR8cpKWc7l00vtSytYO6iavdze1oGPGdprSmA
6N5skslEqXwCIJGKnrw0QSUhNnwAcNWRvEDkZDyrjILaBGJRpwqmg/J5BCKC
XK3Vuny7ttIImT3YlTrSJQQk/BWKSHLFPmbpsrTWfnTQq5yD0y/G2blB1QK8
P5bNYKtqzqvtIYsMSbsm/iKxPaFwUSDHF9uwlO3q8x6fy7of+hESdSaO82kx
CXDlaISJloSrzsYMzkTLoE5EIgagBNFa5WuSq8BPu+6uc40vRLwYXuJUb4+x
yPhkX9pee/QAOmX0JlHJ5rS1OErdzG+tTGHAcCDUFEu+HZjdn4LNEavBCwRg
4z9Xm3NbBOS42vW9W+1GznuYa3s+/5lixfJBeKXXGdfiazICEDNcH7Q7hffD
BO6YDbBwrM53pQJO0gMOUhjeLY0yZ916wWw3PahoSg+fT3y1Wna//dJml9tH
dXUEyyD51wfQUb2HKKbVgnrShGJ0ffWtUV9RlReWfZts2eh0hFUpNiMD/oWO
V9X22WgLZChZbRg8+82pOg9A9lOt20yNwW1V9XYCb9JgEJYqyYO2ipRqSeDk
mTgV2tK8k+4darLUFNsGAMfJMVrXqEBlsVm0K6V3hQdzFSE92YsrgPbxOpGI
nJRWjBd8Ca+3u7PrTG0Ybh3oW7PlneE0sDlnvJAk3R4urpdCs8648iIuQXhw
nTfJigeh389WJZmdJkHj+YtwwdthIyQb8adMihdN7R1GEnoypd3YuTr6B6kC
4pL/nl+8hirXRto4MasHoFqzShRO72fUtVnF+pUp3OlU3zzbvj5jaaNloGCR
lXr6k+4Ba6AsY7CXOh9YEo2argg+d5A646s9TUkCj+nuc7B6atY1pqI24nM9
X1UYvlSdtTo/JUAeoMHw0yuA5PGGi6yvx45OhJGu4oOY2SWP23IVb7K/834V
Fd54Vb1XKVaUbhqT8XG7Mpe/Xk1oQ32aaLgtU352lMCAIinCr+eHfOBCYaLk
bhgLAHpV6/68wqY9FeA2aCLOpR1DQtwcmF6R0dtxaxrUFaxeXOjKwH206Lkh
6hYXaTmhySi5y0xiOtbF6h+Dap1cTE+y2o0gUDZ54YzhNeHuBQnYzEm+0wWJ
YyI/lEtBb6hSshi6YKRlOEZB1Vi3W0CG0B47V5IMJRU3EKi2sm7EmLAoILKA
XysY5aIL8V1W6P+OI5nT8WnzqES+6l1uER5Q/Ir3kJil/2zVv3CNRS7I+FK2
jzwk1WgVrNfD3ykCfikGAD6ILYhX6P0wg/p1rR3D3Eo6CegBW4f0274OMXL/
Mdo4Y+0qXFZzFZoXTl5gSPXACRHdKGmtOpAP2LJT/6flxfaDkcylF1m8vL9K
MwpeifumwlKP2SkHHtkA+/qOE4HHukm5xydHObcFJ+3B9qcdxIm6FvznKWQR
aPAVkGE6JfcEm/JkbzLvpsnlPHkZ7Zpf6gaoRQrovqs3q63uGD4amicTsUfo
yKipG43Z6Pnnp1kOQ2pFJ5zQ3FCXalXAUSGz4r/AwkX/R9HDDERmfNzNeMOJ
1q4xu5nV6zY4F8sokxrIXUaJS7tqR6aUGBEJzs9yThSWXrUm9htGMfyUgqBC
TaSE0ilolbYEj6xXPFF7JkC7x2HtMEDQ1sw/+oep/v1BjiXH8PCZa6o+1G8a
qIDDELRE20NB68zNlbcY3yiJXV21H/8GjLfVM90Z+TKigK8Azl8BHLMiWk/f
Z8t6+crpIXsvR2BjS4y4V4HLN90G+lEXftbgbzlwpKGhbTfg1w5XWp/161jk
/nEkObEy5pgEm0pZin0i4/mgM3ee3HCXHFZQqiZIUSJJjFyFUXnNawY2Hcnf
hbYHpac0L7GFro/nOANlrSOjVK+tbH0qkOhqCWGRmA1cxCBqvp75bWX3zqNP
HM8JYq1zgDZkTSar9rEDO3+wGrZC7vZZfjJtfg+ACjphPHNgLCnBujCWPTjX
WelHNNWl5+3r76Gu42C+z04utk4bqE65S7TvogQRKISY+I0va4OsTdFBldDy
g3WAnrFhPUyey/U01S92fmjrLSIVp1kt16FuCL/Vdkv2HzNH2q7hNywc2PPZ
s2qxDji/W0KcHLIV5EgZmUe8fOFemGtNN8PH8h07jQoEsJyCLKv/jqlTMy+P
Z/Alj3NRzlGZNlb705AFgc6mntywasDGRz5cJr4EQC9PKJ5tHRy8oNTh+yKm
AtgbTETt/SYpWPkkieTGDn5HaQCkv/cexpY9nm4OSxGZHkQO66ZZZg0vTBPK
iK/4t9hVINYkfGiRtyKr7hbdKFnNHDve9yLRwZfx0kPtB8CAO8bPhrn1Uc9S
pNPWiprUrvirrdBBOJu6ku0jCNW4eRHB9K2TwZtoxsx2dUG1CeGSsSdmHQyU
IhR5pZijgzXNqjfJC6Mj7PGXozwI6LUhc9NVj1Nze/WLbsmYSW59AdpZQb7I
BBtlHHOCbAwiECGb4l+KNydVfYhBuHbzl+X7OdB00zo1LEFiYtq4yKhy/WP/
/KoIS89zA/SN/1u4I63MP9e0KZQjbNNz6175BnJqPqvlPmFU9VBPn5OmiNLh
GzqgSnws9RAf11dme6yVNphs1UMewaMg9PXA+1o7t0DMZyuiEDG7UZCnvUIP
7Lemstn8tmpbEFLbY+DvcLbn079AfUK8v+VaJcR8y7NV6qvaSMr93YVzgsOE
GRmSOPt/sVxjTCqAaqdONj/JFq3iVJ+VQM+vo83pRY2DtuPH9TlYwMaTiluI
SCVejPU2GIh5OVEz/6AcW19V9tmQ9nGd6iTDGpArYu7JNco7QZ+Y8tuuXiag
Iuc6UXjmxaVOPPRi4xpe+/cCGF/uS9uWYgG/66K5oh+ZMJO6DeoyR/Eig6CJ
bEplde53o78sfXGA/uTV6zkDDtDaILS/LQTBhlh7hHiXjIimX2uTn9bETP1C
a9JMnpLglsu/Lf9TtLYipjJaCaiuMW8vfGz1+8xGgvaDZLO4zAR1Oy1tulL5
mBo7XDY2dBOMi8EDp4bc7V3evLY58LSXrYLMkBKdeOBGGTWDREzu1dDTyC34
WQwDkEA4FVzoaaz8E6ezz1KbhVAHJQx74scU/FLalOFp9eAUtF5nCvkgCDI0
v45TGTGsHB4hEY24ysf/tkkyxdTF5CPpOAJpZrQEXfGkF+rDDgX+3oAUGyys
UqfROP6Zm3t+tuXh3roZVlU5QyG8w4SNXQ2S4zvWfR0OZXnmjL5xaV7WD9ZJ
Rz9+ZE+I4wefw/l3bi69MvkpbyiMND6zLmsNhm35kQsG1T3DzHLKACN5ND7Z
LlBYXPC6KrKD5sexx/TbHmv94o8/GfrezwZc+7MWYRETmPdcUcSQekF1VurP
OSagbE7+AUDzc0ihLZc6YvBIU/9epYM9ZgLjGTRutYGd3eWH1MI5OJxwpNGY
Jv4XtNo7vcBXPQLPcYssH1FWMIqUv0FY881x4xoGqgkh/ym95GMjnUKhZmDY
UFYFe2a/g+en3EV4Qjqm7msWuLp7kD2FQy9jsKr5kjGhCK4k3welaseNSyUq
kBRlYpZI4bV3pjhcdi65oaM0b9nuQT2eV1FIRYzAFHGmqdYCix91P8GxZRk/
klRnSRsSDChaPbrTeXbHywu+i43PpntS+rMbNtFQXy1pXYJ3UqM8ijLRt99D
v8M7DrRb+iHhe5DFTMBZx6f917vrXsgFM0ppmFZDNHUCXid+gjxMhywSKirc
rNTywJTt5yZIYWmlo7nrsIjC+ty4P8yPphIsszYdl330HDgPFHJ5U2Sfjkii
Q5+SCJ9CEH/GQUHgX2zXPHTRM6yNPo107TzHoFcLqHqV5x2NgPKFbEkHyh67
ldfOyLD5u5M3HMZ0q/tbTkfaGzC6d9+9FEMbhQJnK9kgae2cD3aO5NqeMTnQ
1ecUe+LgvUv5PtfnQHak8KGCdjRsysUm4TGnrVt1KyMEYiUSHtOkvZr1NYcF
FJnYgcDdhOpT/SiNRIv07Wgz9k9TgzXKLI3AqLcRLp7Qq4JlSl6oyHdD9LiA
7f/UOI0RrD4fd6df2/6gEVZwqRF0CzPvmOOWceBdVKgtJkl395Mtk35uQ3uO
yOW44QJ/SX1cNsQrwSe+TRJewhDAtWW1ZqSEaP+xLXMjGCTPe2oC/NCFxJAA
2dKd8rwu5J/QvfPKKgR4GqDZtRpl4r33qYXmHi8G+ys/SVkVrdTAyWbrlwDi
WReO8bn78KOQshWoTMwf72H6ssKNlWOJqRahqzyoowfhliiU5KP0zWPX98G1
iSLXStuncpbwnPLXG5ifsQF6vP5Kn2loKNtRSu9R9QyQL2G0vM5/R0ddf9Wb
+0+MADirJt0u1uQNiP1j4tGuEVjFoXTejjUY5FgT15R26D2B8m5MjWoV9OQc
YbG5AoTroGAHnamriwe//R92EZwKNMDG0jOToZ0CsjNITsgRTkmQWNMz8loT
JsMqOFG7ZA5A7UFtxvUiP0iJN+J9odovZ2BXLh53PN7Nxe5qd02zNBhbHvqJ
rRSvNJVauQf0qV28PYlRqefXTKhVnvSYoVqSJP64uSzgzNsCf6u78TSM7cRg
N7Rhuf/xdOhJdYNuR6T32ByCE4oR77/enu1pzQ5qPioFy3ypa1Qz56AcxPFG
v+VrU5GXWaaPWRx0A1ttl+UHewP8WcV++bV2eXWrPQqnCYRH2iNVVBxKmCf5
fsqF4qpCMgkMMpoko8o211M5LqFhsW/Z7cyW1JxxQ7FcpiaN7SzatwiFqgJ/
xhZy2GlVDQE0JmSZrpMvsXscFMyVs5PTdztUENwfiHAH1h3kCxEzgeXjhGuW
HhUiRqlh4LSwSx/iKtItbHmL7dsPQP6xsUodtrlIsOj7C7j5MuPnhn1P9xmc
e47g8RBOmH7SZfd8dAXIHaHo00SBMtvtzsjoUfZFe0FDu3SyPhR+SwZq/4Ph
ja6twxyL8bwnVds3jTfiKKDbGKmrBjfmCrcOd9b/ua1+2DGyp5ViaCDJQCBe
a27srlOupdSit8QPCaK03X+XbUPBz7amk4uU7POuQmKIOiyU5CSZzcazKeSs
dojFTshsZI7NlsoPXI7p7qVFv+msn27s4VP6xIteO2YPRIiOyICe3sYZ0HQu
bh0nrH+WTvnKARgvtlcQFnI1iTL+NY2s7DRwztTqHpJY4c+UL2QEAmOAXNZp
Rz2PJtACRlW9Zamf34EYr7uIt8g5LTEyfW9PC27W7jQfKkJq6tuaQDEW9rLD
+i/Te+4FR3u75hkC/sEyLzEHu1v9rcK3gkZ5X1Q5qvjcBgS/onmgzPRL0tRu
Ba5vVFR0B2kZGBgrkiy3V7Wyt41uLIuxG77RjVz0lio8q/xRL6MZP2SGq8kG
atfIg5AmlB7B5BbRH0EDghjKZzxpcbpg8KVSluu3bACaL63XySXOXsaUg/fx
3xfngDv8lwiYGeFyOUqtFrw4EiqfNaH6bU6FcpzWIhYh13m2QX39jdk93AnT
PwxTqAaszb8tru8A8F5i5vyyV7OaAKqzfPwLzG08mmLjPR7GpPw8AIFkxmY1
xVKdnvKzonZhjMhI+stMhOYbqZrVr2N6H3tMclLGdH2NxvT3Lgdez9Z/nGqd
9WqXwEUGJ/iempb6LGNPPacUh+Co/+uSNfkX1iX1nS0YMga4zVS+gAMmw1i6
z+vDB2jBqpJnVOcivZiU7lMJjoAlVgrLE9QTpqr9KbDjbTZWyAtS3pbI8ZU8
mnK/piXqrzpYdov7RIgxbxG53tuVfQv/tykhyLFlKqQsPw0DxgERVTeKLcm2
kMTeKTgwvw/3b5mUOYC/zOLZdrvCI2s4EjHaJKLfxk7P8Dxb+sA4prj6K8v1
MFYo7K7FWFQ38hTXN5ZqsZouxul0l6z2+sxvINgTPttoRSq5xK+vw+A1f/L7
LDHEGyGO2U5i7UOiEwal0OCXhvx70J/jV8yCN4wdb8rTbJyRR0JizIQHZ6G6
WE5VPjJpJWYSAenghEDtIOLuRv1ffvLwjXap70U7sLkU4EV992P88iB/25Bt
dHqNkh0MkbDNepDA0f9YWKZYquAL9dN0/nbjvv/EKrC4mGMAoUgqs5l3lpSg
C3Xy0+LUwyzFBCK6+RN4of3YH+wUC46kvimh9260WqMNOda8L4zZde/Qtr+9
arzW3QJL8iVXDYjvYcN8iUNoNm1xfy78mcTCB4cHTvC4SPh8FW55EWl6JU0s
v5FtejzhhTWHNPnNMSu/wW68qgQIAWC0r96GwcIkuWtputIIrVDTyd724fqZ
M6yVKQ8zX0thsTTdDQfyGmjJWvz2Mi9p5ikYf0IEKZTHBTtgAQjFoJzzBwyW
P+6dSbpFxFYYhkS4M6xnsHGrFWzpz0B1qHwhMW321GCQgqrFWeDdx7Xg5H9J
O8cP4qTty/rKs9lgbcvbY0F6ggRXZMB1Br2P257QDyLGX2pMCIjSEPjTlgC2
dWsnWyH9EiXdTaWV3GRD34tVmTuBpBAhpUyXHEjU1rR+lYnkQ3dYdePHrvZ9
Q9AzBl9B7E+uTEMk368JNcWGzi6qyfZR5Vets7oTFSgElpTZ7CIp+PMSxli/
uLIPDkf2EHbgf4SS6/ky2n4yWYMhuoSvk3Zf69M+FqF9YMMdUVzSxq58hent
ncG8d4Z0u64ZUipeDqZl7o2mJfeoBje+FO02v6AbvySH1fM804tuZSFXI44J
4cvH0oGEblmAFqeOAK9BiS8lE8wMomCrh1LyileaRN7RkP72tOTIVFr6qcBu
yx2y4uUynbV6PapZAIpvqGGdyoug4YrPPB40+aoYI6MeXJyirbmCw2C2ZRXL
Ye/Ry4jL8G4g4eV2a6i49omLFXfZMLiFDhQZHv2IBc2cSdo+AaEZLVAKabPI
HBEBCeEWciWReBP9/sjys/ugfC80ZLbKJCz+718/Uc1oX+tjg/W1SoLbooT3
07D969Sas0PQTyrHFolBq6SMT7Fz0Chm5OEIX542fwFAY6Uz1mWeTdC4B5EM
Mw32WCwCT3lyw0oFf6K0zOPEBcvIE8ZyLYXCx9w1WaPlPncmdxPU9DdGDla9
VTB0gJpdBWILncqN0NzkMAH+3tpg+isVk97M/qQ43BELluAvgv1pWa420oy8
zBCtXM6Tr/TauTsQuZJ87YJPNuONqRjOZdqHz8inv+UjkVSb014qjzEk/upQ
LlmHnEuRCKTtc/N8lfPYx8qkwEKZ5gQpWASjBcxCzzYk3EMF4lxzrz8knaev
K/Fxvzbz+URfTYKj51/bE7oVefkrJbpJwL5oSXdTDfbeY/96id/2GeZ4le9t
LlAKF6Cz+0mXJaVuWpsu9GrkzPOLl/Z+x2JJrH1dbYscpbBTRsUOyrMDvUU6
FWMBfmytYxSzZNUHny3ePxQNgZsqXFS2CFbfIRWm/MDeRqSblr45apjGkMOo
yiFHf6pMoR8RS7To2Oq60zv6y7/vSjO6S+rAbGwZacflTwglKq6u2bmba9eU
s+C9UWfOZYzALTi1c9L9QqCIsb4LnV/7lrVaw1hIJkydZ/srbj0pY8WNVxaS
HKdvcWoFpUIjDVuJRl4BjUr+ZhsCYoH0eoyzlPMTvZ371rI1YV/ApzkoOfk/
HDh3QdjUw5GWN3D8tD71zFkfAgPif4FQC5a4fk70jjulIatta6GncRb70LHU
ACciuwBCeqtubaqJSphAsWI6IucEE6AOWf9jTja8MoH76A+TAkyMkxQ2NNuh
nemMx7nHi24p7iFsUu8MOF6LTXQWfx4Pl9MI4CBDYGsUdaktqIdRZ+Ovdvnr
X3rrxsGCEleB0RhlWNRVE62nod9vTfOrt7xeDjwk23m6a+b0qDWjNjIqOMal
m6zCGWlDheA5Ls708CBuPxbgcesO3Z91x14V0s1rnF8mxjXuIT30nywSirjp
/bSq/OEbcmZnb+wORLO84VX91v2PrLJQUCn+0UL9K+Lxs2rq4ciApQ75ydvC
Mmlxeij1zuDyIPmTCcKnGC42uIzGkdvYleMyNjbbMUVcwjTMt41qH7s1USgE
XQBl63ilLr19OJAitv1TNsTjChmv/U6TubPR/UqRbPwevc1oxNZwIlegsYvx
dYimYhcbBwaxTwk4tMzugUvp8U714qgyye0pobzxFdAPvD8ZzJdjctLFMYI0
ALPem/wOIzWsexTa+GOWI+Ww67RY9mkGK3TdH2mKemi8vMjdG9ZwI2++wxIS
V43dcHGpPs17Y0nZKyje2HYhsVaYYZ0CLIA0cGGQkQ+OzgAWhURrOCnwPKE5
1yuQ7Ct+hT0yRscSYiWr2J/KH8sBu0hVMFcT0XdVaAXil5KZ+p7GlkfyaMqu
njGgP8HmHzWu6c6BfXyb8oLVfRfFre0mkFXBAlcA79lqGbD82iyX+X+gQnKY
fheD4hP8YQpkBZ74PKTatgWsgFSwIOn2WF/qqXjdbVD/D4LB0mn9CVaL+U8E
GxXtvsWqVNZ5EpSTYXufLcskngF6ROpBIcoKQWUEfA4v9VLoVMDqtGB265CG
02j0ujaHsQyE97M/VWPQyeFdzM6ta47cEo8SOtZxjlC8tA+ZJm2DsgdHfIto
+eBPaZSG0QSQ0DEHOS6G6tlBAi7g8hR9/F3bREytS0VGbokBAGYjNbt6XyCU
UqG4f6PT/qzGiRPZNfzCRcOkpc+z+0QNfLU8KZ5xk9ItIa65cu8NN/gNCeDj
/7LwhRZojoWAgzwQBKvk8hijYFA6jNP1gx8SWIhPQPIeeH7NOyxNYxHJVrpo
ItBjsulOgJQB2tXxypBj+WfrPHOPoa7o5bwgzaCZeEYJ6v8ByVuW9B/l1sP9
+Wxcach78x3Fpm5iEOpNMvGfig6I+PsHOiHxKc6HOk6hZTZDJoK6n1LhmXvy
pMMqTGtlveBKPB+XOPehm6TDke6uME088LeKz+KUgdlllvBBSdl9OfLrM1Sn
TcPsV6Paw8HdCJkjNdhfvV8gvnETt0OYV9SDmiPrqdOr55NVAIrnnzr9ID69
1G9im8+sFQaz/v9kINrwVUd3l4dmheD/Kk/0+qLI6NOH+1LQgq+ECOy0Q7Vb
twIEe0JtEQLkfsj0T3x0UoaTP2LPkw5geu2pnPeIYeKyWC7MCJuommOYFew5
+GE9KhsekYB6gLRdvQIdo47wVahLrUovaT2OKEhQtkY8BGSIeO1HVfM4lwBJ
IDpGLhxjKUyHcaoio/Q6/xjsADdCYs7hTj3QTymnFnMgB4EMeoUni21YV+sD
K36I0EdqPqAYEviRg/7x+9j6+kURX6Mu2Ve4HjwrubuWDHlPbE2Am3lsyLh8
LBPJzr4CgAr/JRWBJ/HMkIwvSYQgCbnaLAu0hAQvufhx7woKj5iW7B7LFtRS
I92VWO7VmXnvgNMUi6mZIrNiIr0cdoAnOZWExB2jdyRsRCGegesQeR2ZKTRS
cReQt0BdzcLw6saRa0IqQtzkKgSu/DZ9WuBidACX5s5u4DJvlqZjnm/hhNe9
qzMop3OlBb9BHuLiiHhiAn1uVxN0qSnzfvYwUIDnWdfxVzCu9AUtHvMYJXPe
xKxrBfaeq9U9kmsA/vb+PWmOF6/nJ2aRe1ITRJvstREmMLQIW59+4PkmnBQc
wi2XtyZmvjBmi5c31c4ssAzqebh6jg2cKWkVTB3eyYMlsAxGfsV6Jj/edJG8
e/21imOW+fsgYLisTI57ssLfsi3ZxA0wKKg7n9GeVwkQSh5EVjUZoFl/DEmt
/ust7K+/CKh/d1LU7epckdY9s2TIicGX8wf5wybY8E0E28LxwNrxN7o7yOLb
fayH6HwFwt5/DSHw6I05Kge2Tw8ZMH4iB66ZWK4KjLzVUzTmn/rFqR7bde8q
1DddX1pCFmiGtJjEUNBfoMq9bTR9x/f+OGPxsjS+GbNLMMId3dxO0RTzAUIi
LsA8oIlUQdkvToBK5IcTytkGVD35zeYuiqdJzT6kKQCYPjSSbbeRzx+xYHf8
80muBtsiGkmIdEXMhqkKXar6G0hONEFPzblES2vx4bn83JYtLmA7N2Xx3hUM
dn+TulMUoLyFtyP6YFi+B01xx8sg0N57VMGlXsTzWX/tIvdBhbmtv7tMVtqZ
IICP9Jz0B1mUZwU7wuLhjaH9cZc2BcUIhUJD3SmB6MxJks+/lSwMVg9rITZZ
ds6t7BOtrvv/HD3ivv+KtH8734t76iGqIRoONN+TLQC/TqkIfk2F/oMzhUYN
p63o7KFHIMxVFbxT+APCngHLjUtQN5lKqRn+nezxyEr/UOuLE3NV1rEQ+bX8
KeUoilNun0/vkg5rngS06tVa/7OdsQcdYV80ZYLdNQMpUK4iXNsQ/+kVX/Oe
BeWC/8zW9fa16FmU6PeITLPI9VFJ8q75Xh0vwlhNVL3V6yLs7Cb4tjlDdgZu
GhoewJAtzMuy69aPR2r2FMvvFfrXBExnYjzIh+2CCh4S9D/lv9nyjSe7aNNy
tsKc4/CQk/2glXz38j3ayZ32sRoE61N34tNsOz2c/bpjPFYV7uo8pu/h5vbK
2nJHtonniY+ayxVyFdIOvC1fBT9vNxELTLY6yyQ5mJy063gOrV1Fj5jJ8olV
sDz5cHiFOUkpUj9Ze0w9n9fqB7F7iH8Qlt0q2NIj42MkJALXMHcrMnymCUAH
T4PWMS/10vhHabyZLJy8iiLFLL+AhfQzd4cSqymwDhV958CbkKjnDTHtpjY/
XnZKM3zpn8M4qW7cTvlLFBYIFMpfLWPHNusFnwnrKfAwcQteLDYQ7LSUCFDZ
NHtVn7RmzbftI/f3Z729lBCMnbZ5tMX1eR7pJUCL4bk7xDSEwmG91awUuBp2
QztHn6kFzZKWD9UZ3CZe8LtgKaBzPRAtoq7qksIM2XURBAJlSkyVTrVmymmR
MhR9F9QJZCNKHrDUahZioc2G+xxjtqeuzLFdv3FaqbiseIM/suNXc4713gQH
9hQQdVUwrbF6zk7pz3NE00kk5tbfebrUR9yEF2h31GTfFzCvyIiPmIkIxyta
3bHJdgkq4bpJXVBoj2RXejwPBdSTdOxRyTOewQvoEWcjNEpNj0gFSBPmLIzX
JdYSKkz7mgu6qDg4fgym5X/ufoUp1ydJ2dxZucTV9xockSzCk64G417l5QUV
1QiKyubyVAfkGNWdjamLRlG8dQ35ibTsWbY4Yz9i0AWc68Oa+YPpdRf4+k12
l2JK5Z365xSEGGTwK/PmJ3W/WznDPuwEJTibRXLc2PGYEEstDIBIBeD0e00Q
neo4J3BZVIefvbc0g2MMx3UsjNVSqjT3wh3n7UrgEvpkWBFHvcgBDVey1RHM
R4sb264hy5wCY9m16Ro76OUYsIe4agMDibRo1FNAmh1j8pNcWBd7AgyW7Xl8
9wBrgBBVFdrtoAs/3gCk1MxBbN+7KTjU/03TXhxOug6y6VAPjNxLJDIPxXJ3
KrInEcwwfNaMu8DhkuTy6d64edDns69hbfs+hXwMZXkAWbaTscqK2levyVvK
uPMy3ZJRNMLQ8/CCVmVDRVbFPipFeBJFFq4aEOs6ljDwnQTRMpZssp3VcOLE
cZ2DAvnTqLHtM5ZWQpbNel2U/u7ugHTyU5BRXtz8yLn70f72myyqJ1qbCvO/
+z4SrGAZjt8Jb1oFPEZez2QseavGqYDmIFy/GSSjvd1uC2GUqBawvNi+f/aZ
u250jcO1ur4CvXp0NcKI2+fJ+EuUOVasDHaZvKW0Lgqnteyn7LzKyJ/6AxZC
kv3ulYf8KTBKzwAoqqP9RhwjA+Mt30FQIb8ZcFaD4jL1iE8qOxQLZAqieUf8
IGDhRHJKGdAAUbT3pt0618pWgMk0yBB9Pdl5jSr2sAwF04XVMMJBJDdhAULh
dn2ig7SW4IvgM/3S23yteS6Lf4tTLfzNdPBuTOs6s0ymF2/aZ3lfNeXQEWgi
dMmpHP3AI933Jv+UrzwmzFbVYRAhaQGaGL1oU/fE8aRx0fuEr2MeYl6gv7pg
Gt83HHowTZMiAF3BkmbiJgjaFjghwPbMnrNX49qa2wJG7i/lS08SzXs7Abur
p3sCjKPRuziBzLzSBuuTGO0bVHScRPdz6BahbYqgBO7EVGnwS8orJ3VwukuC
HMyGh1rHNlGHBMFQPe/rvJKoTx+u6efHlCrYXTJVKt3kv/Q2Rt7oq2m7AX6C
n676gMufeNFq9d9wjQAtteJiPhvS9G3o9w3IS7Onk1C66RywUbgnKGKOD/XJ
U22EYFTUofnXNIRZJncz1hIq9JVGx3abb37HERiI3lsCOGRF9woXwqx5LxAb
9qiPE6W87p2VWr//Le9ZsW7NuvO+GeLQ9crbsbmGztleuyz+M/gFvjG9cFed
4v5eAC8=

`pragma protect end_protected
