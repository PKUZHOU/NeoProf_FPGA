// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Jto+C/r1gxz5rA7vvuH7eouYpSy0PQ+bZR0KN0iRzXCcPXO1sazuSoz1ycKS
X3CZDUxxha2NWcgO5L52nKmQNUmLDOcesHokWu7cBvD+zajqRLheQ+vpw9jJ
1ZJ9kr84wqIeaZKDTEZt4tkFpoeKM0HKp2WIWXdpmec1YNrldzB+Iwv65BRH
Tjb5fa6d//JNHuxOuSxy3kLlE78qMocbOR81oPm5RNruAWWE/OZ2MhYaVpGA
sBFt9KuqF5hWWyu0ipSn+npYSZe0xBqdtvAdRe49bKg1MCEOi3JAJviJ9wkk
ze1awcEUX68Nk2WWJ8L3ZBDzVZ9uMTn0/1egaE3AyQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
TEzWXArKIh1WCmcejr7MLEUxqo9R+cxPg6eUSxEIEidpxktvtS/HEuhDYSpL
qSMepsh55x8cwh9Jf0Lq2ujNyu2ND8U8bg4lDSKzSyBTYDte8AFCoQNuJqGu
ZGZW74Z5h8k2jqHQ9nbP8sBnQVZoCg/QVrWLpHHrVnDvM81BCPMdecOpg/RQ
Ooqv6eeFoC741slyov4/brua7B1rR0jjgMa8FEqGZQkkFNKLMFxu73bw5C+7
Zw7MxqskE/g1c+ts+v6BN978qNrePHOPSMifl6VT66Zv9HXZjOwRbake4jrW
WLtby4Jl8fK8BidWIsUNXTzTXD6g2zHvKKFg2G8M+A==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
hIHKWent8k/OUUgmTSRXq7k/vtX0iz9P8Wgp9E7rpRNLkZ7yT8459cGRuO9v
4yoQL+lJ7EQoEZlb35sJ1lMaBobYwAXj5YCgJjbOZwCrn4e72s8MS44oQmjR
1sTtTLpflG47h22fbA549TeRPGLiEwlPpioz0PbfbiTkWEEdyHq9189tZUcn
cZhwIZDZ5Y2dwAgCiLADZ/dZNST/voja5KG/Wmd6zSRObWBgyL+W1iceL7TC
0TRP42armE9kAR7ZsuzKxLh5xBrzUYgCUGiiHyGAma9jZd0yYaCukeRd0Dzj
Q4cR0PzrylZ+KxzXj4I+69aVIW6okUq7y60zgftR8A==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Fmn8y8l1Ahi3jIFw6qZYU7iCNoHsOszPEnLcfHC768uK0h7w0X1/UD2zwYO0
9doy3msuK2EM/7GINoC0Jc+Y/lKw2YySTpxdtM7YHUN8dHlKZnQLVLJ1TcEN
KUUz5nBnVtAPo1Wc9s8HSzN6OFCHsS05asBc7LN8ZwBZ52oRQXg=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
tMjm2/I7mRER1Rt0KrVnaVcP9ygypss0G7X118pYezf11nHpbO4VXAZfFpXC
Hwd7ahNzV44ZegOnSrRnV/i8DHfWhd1uhIES3wWuCMrNJhTxvVuzvdHmr2Ov
uqtSOWSWDdfvoUmqzWKj3ZUY1qRwJlkHSyjdX17QTTANsVcYDUVhqVCNNrVh
ijMXk4twZMsAYBKxF7mICXO0iUMaDrGmnLsmN/lAOZ5GVxq3wvoTE2eArr9w
9R/gPPnkBzA+U7C+43422fCOxYfpUTg3C/cRy7/W6J58qZjpLkJqs8uOsJNT
P+D/N5AKBZknUe3Ht1b1XPsg7WFCmn7fOk7C+8uiG5o6vsa0lhuvPc/37hzf
C1AscnT4LBuu1UZjUCAxWxvVS+VuACI006KJpq1s52aEFAR4C9HQVqoAJnQq
T5lDdpp1oVKCMoTQSSnBKgLru4mzTdIpyBtbECnhs0SInWMJ6fZS2k3CAMgV
sy91T4EiyH3WSrBSKaiKFvq7LfWSL36g


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
IA7wtlz30zLeH8CLspGCtLJyUYD2avy8B7KmL361ZzkYTOsGe/vQ0UuPp8gB
0Sy6wkQQjFdBpNaQOukHkisytt/IPzLKV95m8RYNjASaORC6nOIt/7o0b3jo
jfJa5K1L3J53JYMHXyOVnb8QKNRNO0Qa2+oi52F8U7cCqKdPNxo=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
L0wzAGVMc3O39fYr2Wytl7Fy2dm3EnBxHHr2O88Se/gq1lx4pUzDG0zKixU5
2vS751GPp9IuK6nFhVTGMOqZgz5aJXmbuUeWSMU78y2UZUFXbBb3ef1V7bSe
REFhd3UBIeZeC8kfeCqbqaIDzZP7VyxIZlk4bORRE62MjEpQ5tw=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 3952)
`pragma protect data_block
BaevXNQnvDB5+2gu8DPcY0xsA4iqrYc5jn9cFFrg0Tt50t1dz3UHPcDDeeib
k12YxKH6yhuuND8r6cOPd0pT43ePxfzUxYYMWZtS9IpXCSAYlmex8iB1g8YQ
F19DBxECAdTf9KckmIhXEr19J6/E4oj4hCEIhidZ5BP2eJej8rTkpiwVDxXW
DiKyADz8JFI++TkxP+i7ClO/E30/bw9aTam7iS/qLqi4/V9oC405UZ6olomV
rvmzYfjP3YtteWsCJsbXcQTQeF2JhW3hcN63hDZud1ug8J65SePxO/bf75Cn
F6d7kyq4oDHiiORcpThdkaLRrj+DvlS8OVIgEvEmlCqpnDXj3DbzR0s+EDUN
n8lHaoIsSXAjTcz33jSPMhcgXulMGXBLlUDtuJRhS/ULzMiPnxq88PWv6c/i
Ztzem7ACh89x7sBIvUZCGtOEc1Ae3xLhU24KQ8Aj0kX6bUEhBoeFlIZwuUjp
ov8lhacAwiE09rlVh5rfdTi2WlKY1QnG4OEyV58aIqXEHl7sbQAtVyTANdQs
CJYDZ30/5+2O1rniQ+ARh39qnBwWWLhr80UeQdkWHihKGwV8QLzR/NeDqmGs
vz1Lj9E4dIIJKsB4qYkUFqx90PTX4q+r8npIvxaQCCl6miXgMBuAhHNst1Fh
goPmgW8qgSJm2VtbyB0GXtH/cPHyERglyUFA4MD27eMoxSPBvaICp6PQFVsY
QbEI0VUVMDKkJEobOYK86YVQWkZKxFBTU31+7XNM6bUp6YeAzgH0NVYPCFT/
+PShYRnONjrzuxauFbUqxNQ+0M6bGjXkWG5QViEDZQ07yt6qkD3fj3cAh6LN
DDTEvz+WMcXA0jC3f5g91rONb5lYHcOQ5x/3eCX+5V8eAaTakrtJbUPrHX5H
Bcrb4MlWBBkg1L2D5Ig9zCo4TNJ0ro48WVjpnXqmWb8tV9UPoHWqxzFkzXt9
xS3ZH43ppv3qEaPFsEW2pJ/StwNfblPTE/YcdQ1W+MWLkcm2kw9V/hFWhb0z
lXrfQkfnHaqhhtQCvsWYucPDcIHU0Jt0tv8Bw6UEbEtrTkjiL3sNQdfSQnSP
jY7Onzemd89Mr3fPYowKrnqE7duqeDhgx5JES0wtZxNr1PyfHAXuC/oE0yR4
ih6YTyJ2rCtFiPSG668hj71K427+CMohO8CqYFA316T9zKUrtlC7dr1PJrQl
RdqrY3VHYYguWvtr6Hq3LjO0OGt3IJwclxY5aL+l/efnHFRxjadhf0ITFsRg
mnkjFZpdUP2u7gfgBR/dA9Uo2/tSxWvAT0OYszFfualt05kqpLdmER9RB1ZQ
d7GxnwWLbyDFPN3mWX0BWwN8y53r2jEHEl5Wlu20IY80CWqzcsS/giXamRsr
B0uYJnR3OkDKXbRv9lrwTGNN0TwcWOvYzyYJmDrZ/WOlk6YbTeVIvbXiYnt1
lZlLRtgC3yO2l9y93/BpRjJAJu2UJcNzeob+6UxWXJvqLf0Icxv5SwYykQY4
U6uPhxY4gqqUQSPRtLCCC0UGxkhLEyHyIxB4MrHOY7CxrYd5eWDK3GTSMx5L
R8oclgG0tukbhtTHbcO4VpYJ9Xc/jM+i6gmOkTQq/4KJixP5bDLg5en70Tb+
puYDigErGhudb22P3uYteFVVYfcgX343LaJ5n1ddNp3HAlYMSfjVVvzOwWrB
aMi1q8jySX6PZP8FRKyi8P9gptIDdx4ch+2X7Wy73/HZ1A445M68QQCatWfJ
WLPvZGMjecQ9BId2JPr5fN5vYLPNsZHIelTE3FU6gZrB4jxQCkvtqsaG7ejY
1XULacJtZm3jWCQXqfQsM3qBGmDws1/mfV0Ic9rfSp8S435DC/ODnCGEukEN
glpqLIOqq41fnmvLpS5TAoZyBE8q+raX6TAUbSxehR2PwOwUq5tqRrvtTn+i
pBvTVgq2GUbuRK2lUHTxt7KQwIc1FvR20zZz9oXxifenBxwozRPzNrOulDG/
EG9vuoXrBt7oCscNHC/0hSFg2e4KazR1/vx2m9UX8sE3uBq6gf4rz/s7mkfJ
xnh4v13DCckZFOp+QvAENTsq8Jktf4zfE3StM07DQ14PMzq/kTysU5wHCnuk
wSpx3R+d0L07fd3wnYSdRt3UQipmhBw2fwWGyH/fujlanazDxlh62qxGyx+h
w6WMZVUPV5u8DhkFx1RN/r1Jd608B3AJ2Ck/5f1nJKirWPdnz+jjmfXmZH3b
W8Emfv2wAAZAt7TalgbCu38DgDZc8hEM0vouxiV+sPKYGDkhzVWKLDbFvT56
wcGzf4zCM5VisLx6RI7QSZzG9iFwwcUZZCAbXgbHc2Y1YT6wQxZO+5vtSPoo
7X3wbaioMZgpvEC9sbphQSRjFz0yFerDI7kE/hBNW5cVeceg4ajcWJ8bAV7o
7NXg6f28nz+5JsTz4rtAcI9IbWFssdMIeBrabCk5iCQNVYMTCxj3pImVnK6M
C1WYAONhlKJGlOBozUrYpvEz0XbvJUFXWlP2A3zATWk7oOXJ1ywcUcqKOILG
1u0grzDF73xyEOxY/lXOA+88JmzyyJj0IqVnrwH/Zy1pTjo4Nl3ykPvCzQ9T
+VubBcc0B2kcTnQ3duztYuyBSgZjQvEka5m+4CqhdCCU3FLh6D+Cf75u6fbD
167CUp62W44RWuM302KErnU25JMdUH2aZKROgdl69RfddgvjSzB30fsODJ2z
EsX5vkn3slGlvX2be1PtaFTZSsuKZRLQJRxPPqEvnSrQOieeCmqcxiL98ssT
unsbrBM/12FAD3m5qW+X7e/wCLz8BLzJqGd1Xv8+ip3oqX4anYQMG13WFuTV
J7mVYmqsiifJeBV/BpGFEFEC1GB1DZEAmZ5sE7ViKjTPxJOLdjc+zhVbf7vk
3ramkby+Q+Yqvjb4BJWJGDVaYDgiPsBq7dLZtI0SrKo2zytKezODJGjvI9LP
e783lR7Jtm/bLG4hLcNMDr5xc/Ywww+v8qTqIU60qvoByyg2TSFmX2CfC8G1
Ad2q8kHbJL2KCmq8/Sacqk6JDbvI44VTsnT9xYZkNz/T42vgTdR3Y8+jwBeu
ifdSOQAAPGiFvHe2Ms0JGK4w1UDgsY9uL86dMVT5lzejRX7nAzKxd8JPuBX/
+gJ46e7AptjlLUStvhQXRR8gSbNgeGQ6EyQ+aKq8Bia/gq5PySthBwd35OBJ
Zdh/MdZdfzf8G5+fcEwfaIEDGIsfeem9XwS5nsB3SH/EKqGhmOlgk26saUce
AiK8g2sNce9c47eT0WzG8Dm6w56w4IKEQ2zXZemO30kJzYwQOslZzFQ5SUr9
wf7HHqgEtftZF2TzZAVL4KK93MSgqVndUQTjVAi/STk4ytcEOzQ7gPUOUyZJ
ljhP7V0DZcsB2ZVrrMtricWWBfFugOh8tgYMQeRjCtkTAc+XDEkLVQq4t+8M
y9bMraNdDcPrijfjsYnVJc3VZQSvXSbEPD640Yrop6XWnBGJjvschm7kuivq
qSPzH+JMbY9mTN5LLS0/MRsxuD6gRQEXppczLBwluXhHSiK02CUcmnroLY78
M9arVhsb3QkQsix3vooRYI5VMTNUhbaVz9sxfC9qguwihSKVK8SODFmpwcc3
8wAXAvm/E6N0/laZThNXQcMzWnEjVumWuzm+7wO97lnDMvIliI6PJpmhSNBD
Yi6aYT/EeRJbJ6IUWuHSsRjOHFVDwfBad3NP2StTE8pnCQ6dn9YgKKdHeUYd
lTbML6ZG6+mBLUsGCb6pqtjKBbRYew4oSp5F6bm/fNNFN3pJCnoIITO8Uy5O
7zlAEGWNOLLoenq8o3GdXZqvPPwWgY9QQQ9JRm7xOcQo87gcbBAiXAjGBY4L
wF5PQrJ2u8N0tpZX//DAAREkx30npe1NaSLBcuFEsGJWAOVLcAF4GjQ3tnFO
v8TGtp+MCcgCq12RTKWaZNNPR7bfygrDXZnGI3KxQxe+dQHpERL/nMmG6toh
xnvttTGDSU9Jsi6vaK6GqAC7q+3GuPfB7rJYg5LSGNw3+PF9FfM02DLiqH6P
/YJBubmivXyisMQ6qnZpATTVtMjwYjbXWm3hvW1+bknOmTPxEBmbEd9qTE0W
QcUI0ya8hRV0s6OPe96ic+laCR012QLLGkkYlqZVyjvtCvqEje4+P0A89lfS
cVSwixROTA+fFKVhUy+pgU3yG0WHMukaUBCNJQov6yQoqLphEabZjId6++zP
vSP1LQGA6lNRb0iT8N9Qb44BQHqChmTVUtrDnCEgeDjg7x4quoHf2KvIYqsb
4WWPJUx9hxHFdNvCX/rPbIsASiQ48Ri1ZAbNPZEbQv6sfJmrnWp/kjlLFrMZ
5iPHg7UR7AWpTo6CM4vDUSvbqLeDu5+4hDfToRVr1SB+xT6u4wHwB6/AwPK2
QJoh8AqoiYiiTnlslWiBW+2yLOxiqCtiv3gwMTGDIuncXkxwl55Ht3vwDKCL
ZwnBdtxMq92Q7wI5fvu4z0mCfd/kBSRKU4CGQvVtDIdtczEXH7Hkfbb+CZp5
6Qs8l2ZQI188KyGAMa6eCAfRKsLEcOWiNFKm+FhSa2GYHL6zs7Sz0na7B/sG
Zh4HkUh3De2XORmG0aCVIYL5AEwD+0RTdv5VbrO4ohMgjrV/dhapJqjoMJ+U
LTfnggzIyBi17PoDyPYNRjlkwmxNMmuVW22ikvh0mR/8D5RjtrzHLawOmMFi
RKGqNNdFPmiCTRzIWUvStagsjxfY95ESTCiA2g+imPeYsJeeJGEeHEVjRh0/
8/XYgkBRAW2DMLYakdRxxs+w5HbXso1GvqlTMV4GTkIgr5OdOG1YWxwxR4eD
33WP/5Cnx4zwztqyfS4wkPFZCOgVvr+lXhF5HTLeWNCu+xHA+PB8lny71l5f
5NFTDqWAi0iC3eKSeSYRbck6m1HZt4i0X5SGJHtrasNQLcht0p8ph9f6AM5H
Ez0MKjVz3Zcdd+nPcVGVVQR8OhHmpFBtfchWj+jDEp9C09qFTBrMupoxRPOS
a1cMEafKXcGNZ7DrhwdLBlpNQQQBRmqoogghJlgTVqQmhRALP0bQO6hBstIP
2C+fM6I+I064BdvZLX3Z8SDZuFvMEy8yki42W/ORDqNWNOn+B/YVYLDM2jf1
JH5IvaJU5qbH38V3daANFwl+KzGFuPH6mNH7mepNpiI/MG5bZ2NTH+oe6fJE
20pYG71nec/p2lMxmAabcuF/qWCFJ60pW3LDMV6G4o41vL92KG2yC3WsiWAh
HAx3Bp/v8div1y6t3XzdCq8pNA9ErZpTRwQXvIg/Utyh4YYmJQ==

`pragma protect end_protected
