`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
rngEClwSJKQgPM+Ij78/2nywZzom5Y+LsBY4acp+V8wnDEhcIQIJTvvxHarvVVvY
AejtFaEAbLTna5q/tIqhFTJmye5Ghg3h0lXP55i42tKjsuOfP3TCaMW7SDwp4Eby
BMR2iIaNiU662TA3hdURAkBgZBBgNQmKS1NFqWWxkoc=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 22816), data_block
wj8iYVR4VZ334vR94NGHoccoCU7O4E+pl5ILbMrCNovqOItcPO6IC9/LXh0kklZg
dqKbKpaCGTJgKq6ytJKgDr8y9UNW5y1iSU1ZG99KCoHH8OiEholwRQu6azWJMGIa
bR0CYBhnOM8nwW9cTEEebW7qtKFzQEQvkK/9I7Yppo0Y7y62gDDxe+7J+R1x2xer
okazVCQ8+lDNVcXpr7RVrAAUVSApWGp+ARVhyQh4GUVa+clWR3NraPZVUzgYvssv
tfIBM63hpw8KioKxXEsXSy5Flf6tDd9+vG2NILaL8D8eMpoAQBZLKM6mL+GPmjVM
qkHZAXk/dus23FqfdnpKYUF3nQEgzKgTAM9rq6s/ddyBs/xDd/HRJK3FrTK1BTPf
oqt3J1JKincT86NWTGX6BPcfHUYWjDag1H+hprV+JxzhZ30nz79W0UWXRFRIQFzA
ulWkCdYP0PftcgNX3Nqsol6zMixCd7hIfuH1jN0OHsBWz2/rh6RpmoK5UHzPNlmw
4wCbW9iV3hVFotIFF/aIYxRatc0P9EPix+0aiLgZ3Vb+j12zDcGJk/3o2jS7lZ3M
KX8b+nCN3PCtJVJj2Hh3tVhl3TK2EkJHnIhx5rvuYhyJinF9Ql8F/JTgr49wr0U1
ckgJdS/Xe7P/H9BjGSdKiIF/NzypRsH8ayG7nIdNOtQt/4aymBtEgT6YQUkNsj8Q
rC5VBhrmsmQz2Zks0omygRL197+u1bq+P5VnHQQBM/GR1dQFqJGCzmO2kdEOo1Qd
ysMERHvjcjyyYzeG47cN5qIHARjUWdQt5rfpj7DfWtcNQFlToj6HLU6qxwMhpnEb
eSNeW1OTIXFgGk3gFsNZe1b4smn6EVxENbvmsQyJwB38BFLMYMIv5wba6iv6b1/F
FHrOIYYYtLGk3WFSa42agru6yLxxuVKYD9ssEH+cRsOFhWUrChfC6oqbZXo1XO5c
fMkyivZah66mhXzJplx5q9QXAQ0ago+RRWAKca059xV9CjKB597GgHgTtpfmQAuJ
ekE3alDN01hAq98Rh30gJg9/qn0/zGo1QgzDYUpiLcWa9w/hzF2xvmSRSUTPhrhN
h5+z+K1IcvHFSLm7r7Q+ICeBdGjcyO/wt+nR5grazeDY6nxHSFOzwvbkXR+nfFjx
Ht/9YnYlbzk4ZZqDCZFV371oEfh4F+JtculRw4NsdnVZtve0Tm2ZTLQyQskl7UJZ
FNiTnsFasT7xGOmXwfa9l0clMpvoLX5IEYRh8HBQA8bicIeySQ8yy6nxhEViPNZW
Jv6Mc1uUXhe86g4udG0N54YeVeO67sL2l/XM+YnggzO7phW1BWZn/ex9hV+wB0kO
7Gu5DmsM2pEpGMvs6zS2i1hp7gKJON6OirVZm0xw4s9IfczrhuK0KfQXOfMabp97
jlMaX7/kQAHV54obIMIhxhJxXWUVIhY0EeJ2c6UUBWSbMkofudZirKMePu/9KkRK
CxA7RikyaYFu20DiiaYZdf1Cyw7j6TStWH6fIrC7C023xR2/qIQyx2OdVFX9xRrN
5v1ES27hovoeqLu8hK6mAsuUTuWU2s/AfE2Ii/ieIOm4AbryV5t29NFBo6+gGWLg
gJnN7jKCWNBxkSQe+pt/KQddbloh45uQX/vZPNDE+FndqeMElE3f0GgRcNpvfKJ6
/SMQIPPZHgbLkZYYhxL4uz9xH08CB/a7Yaj82ZUvGEYgMuY+G5dBxNtcVZK2+hTx
rZNTtnh74qoRVywF3fcnKcligvTKqnvZ/+sda9cDfluCsA3L8ikIrMoVvcFaTPlZ
HFPIUYHiQReD7QxoGqLAiDQpMO20k1qOU1WghgGgV869WAEhukQvBZdzZ3AqXFwD
TQG11AAw8847ms1E0o9pvznlj670wOjrU7rlz+sjYmdHdlUPyIr/DLlIyMzgCmOr
k6ByR+3KCUYytBtdBPSv7g1JcMir8m5ZY4battl8KMLbLBP5Qoa/5VkJCRx6ngcW
uG2PQ+ODP/mydUJ3TKCqx9w3kgQYr8OOqViMNd8E4u3PT1B0ja7+y8gFbSo2+F4R
t+Y2JMpcDguAandxFlXF6fbjaH6296KqANR0fQPMOakBKSIG1GogZml/Rv6EYfIa
cqRsV3bqQsnmndnq1d6djsEr3e+lez8onQMepVQ7rfhB/2zTJx9Hr+G3KjeX2bUs
d4yOOKmpdq5vz755HQNun+Ii3nTcrcwQEpBD6mMbeDMAymvTtn0ZVpmFPMEDyAsC
4KQmQnmRv+z0kcQ3shXnmEK9Cp5LQRLzFnPK10M3lMjfax0HhZRq4HNil51XKj0I
RgpXidJ8VIHEJmFk32pdE6w/fdo0LiqvsUoIwxpi5xjOdBKMMZaKiczNE5qazMeE
6gaNcCFjER5m0MSFb14Gy4HEs2oudJVjumxgnIWRawE/b+UYCNl1PKLAbzuwRcAI
C31LsTxNexSWCP0bC9qHeoM55MwRTxKD24dukWoNDmFinsJ9WLN4+jwA2O3ehCjy
j1PRd8Qvcb6kyxxiUrVAH8cE3PBUQR/XTzpGxgtZF1J12FQq+dt0gZpQiFqcyR1+
j8ND+II//SMGijZBY8ppn111UtwIkuZCAITDv0s6UgcXsAicQ7pKiWXJSrL784zn
v3inkqatXXfkiMEvQUkS/CHGRup1ZQCFl3rPq+8fhfTTXAvcdAWH6cSIQBXs1Zcy
1N4su0GDmRPuj6EPuNkrEsSC4rC5RxZrftzcVPFIlVRB1D86i5bVClWewvLHyDY4
hT0IWHh7Q/U9NqxsMmDYXGhcydHN2XU/juZ57CPOrO1LsulLXFnq6uVQR8KWu++j
AIUHepP/k+1xOkQuoMpok7Zyqi+rAHkhIWFn+bKzgDQvEExvWlAKnTsjySu7jfVk
83ABZz/vA9fEfyW1y3dNX4MYC10yNp/Sfqurpw9PDm7YbZIR+HkBIR8oyevq9LYp
X9IpR4NKNx+WqxECkJPrL0UCCCerkUDqwjrY9WXbyE3fIChvItdJljiFsCPvXQ2c
Ma9J/gavVafFqU0y9+WF4kG6L2wcXm/aX2K7+FVmLkj6DAdl0OIajNiepO2vYLKU
3DdttkArVl2WbDQPdhXfE5GS4WPqRcNfBgj36pluuMk8bkZMRWLmSZUK7c3qniOu
e30Gr2ywxDPkg7Ndd2d5SwEuKgfbbNjkwu9ykvjlGpD3J3UglHKA8DnGmrMdlSQ6
h37YG5YHO/H35Vi5TZT0BiV8O2xADM2tjPyyfU1qH3hAybOER/ARpaGuuE92ru0s
eb9GXqSLzm4XCzMWaYxw/bO7+kGKt2hadmZhFHl9hcjOf/Qfh3brcRCn62jRlt97
GTspAi7STE8NiCUpTT1zF3zlrV/z+LzfTdZGgKug1OdNqWbvJYJYPaPAjRnHkuFD
tUxbkHgYafDezjh6PuCCjfIcbY3J2HRk9bYCLqx6Y61gHpY6pB8wbDaiTUrli54Y
ZgonP+KsZQAASwtn4Z5omfN6wxqlsv4WIg05iCMiFlu7tHzrHx2Comb3siwd78RK
HJ6zZGt/fuLci43LNYdIjfQjSVibupGc4oj7xr5vwfv2OUjhxDMvJCVDfWn15Z9Q
SSKz5fuuawfoTVOAa8B2wDwyQDbXaLwM06a2RbptMd1lMh2B8io2NrlGXY1OYvWj
RxK+fbZSHTxxTkbAPi651OykIXCsLUzEo0TM1cAi8V1QGv3yK2HNtLEeowDh+6l/
SeHB1rPuY8lt57bOmsr8xPbNHGM5jFnl9oMAVna8QdQnVEhUmO0cSHVkkKdHJxZd
wATGFllPJKoIXyspBCYYdf3LZvMDTvZroXgdwiMwGIpu2VuBk4hEXe3RiCmFGVIV
7xAQ8i4+jeH0BU8tmRHWV8Et9iDlb9dxTdigB/75BYL8lZsw18CCS92uQquPDpDq
ei0v8vmAkYK8T8cRYP6X9hBgr5Ttf9oL0fdTP6PhHx3IGA5a1+qaBv5VxqN0QLUk
/25/qVjblk051trkUzrtD0bTsCVraCUc5XuUpmgXATuqYHcrxJ/FozokNMx9XFQf
yQlPTCOCBLVPkr+aBB9zPlZRcpI+RrvAD7n79z1b81YOMPFd3WvFgAEGsSWf8OJU
YkHhG4zNzBImsZmJVS7BQ6VoeQr/FM9H41oAE9PZCspGLzuMEvZtarEZV/hGULPQ
/OWKiSbBvlz/tM2VAzAt32odPtCAQyUOXD2Jt2Kk9ey8Vn4ozH2SvyH+i0CMqj5X
e5eXgLuL4XPSyhU/kGuAVyrDjnDYDUeDK7PPJOK8VsJl48LPIW4BjWZvj5uTuarB
XtCD5etDWZ/bABov5Qsc5KUIxqcmh2OTVE/xiJ2aVHJWu72vBD1HnsSSPWrFQfG9
yRPxwXqfS9gNCvaCswR3mxIODMpo6zCYutP5hSu27ju2dYdEYkM4ioEP5WiX+tGC
Ogtv2DnyV358mLLG6W+7sVQE1SqN9jwCbR9RCZw8s/fXjx4P/i1SFjackWxWIcyr
Y5cphYR04XyA+VoaAeJ0VgAuJZEH9gIidmZoqBp2J2FcOWX36RN+YglewvsVUK5U
iOfVj1LGWyZpPb3hMWOkLr2OzkchiNBGQuBqtRItMV9GEI26Fohj3PHBdIujU0Hx
LFwi97ssx7HBMndxxqFHyp8C/K4vcY7j5Ke4JWc0J/5xGY2jCljNgvyy7PL7hVXr
hUNDhuSMB6qwAHigjLNKgeQX9hHzYdEd1z8OGFKtgUiw1yvcP6a4HToXJYky+8VA
oRIMXZnfUYvmEUNorzHZddgfLx4bpL1pSau41ewOEz9F/5HMKlvOQKx32mzmAiEm
VC3gqBt+IgerPKuGQ7K7ECPTOD8nruaj3x9ohzrf/rkyHy89Senbe4QWIFGDNdom
gTgr2+FFxp0mRx5DonhgHgXKj5xGW9pjqjdF+RJ2/rVdxzCpotdUMST5wyDL+jnR
byl/IYzm5R8otSL6Zr6+JNy49l7l5khRSg/R31fZO/G3axm+X9uMYhUOtmZKd6RT
nOY9rLz9SQKDf47oyrFSUT7xqDW0hcQQKh2yhQZnXm48fVWZ7XmVnMrgRyWUYsCQ
3ZFkkczoHLTB61nEBj/pHb44/mOX84U6xKuzVhPNf2pxZFxpb5MSDanXM9qXFYkb
S3NbfDBCItrW9krfdp2Os2yntBj7qQs7+h7PJIFYmDIHkdO2JG1QMvFZLoS0ExCS
qIv3r6wYf+6IhUnQgdJp+skK6OJYfFNNIK2JMP00DJzSHNUkdcD/qFDwx9lS+eTK
nRQ1O+dFUOFACfwKNsKQz/VU/KcsbQ6CAlsCdjOMKLDyzxguIuOZrLe2LfbqPo9g
iSMk3hTpJPgGVowbQJaejWcpdikaFPJ2c3PMW4tKVZwRQyubYTD7Gd0B+Qa4lvuZ
MMCK7JeD5IlfLHvKwwXSunmEDfqkNDHV+WXEOUUCONz//PR9ICXEWuRgda6qaB4q
IyijeW8ldFWZJzlP/7hPVg0TZq1RfQr0w5Lo85kU2npTG+FJhMhJaFDrhyyFzEfp
yRTI/DsxL1kOn21AMGDJXN5G1ShQETTlLX8YHrYve96vaRBO2OIHUaHFqpBjlAiQ
slHeQfI338q9PkfCIPIWL4KIco8MO0PjQTeVTDh3vz7sFDbmy0P9l5EOlCmmaX/S
ExoAiezcM5piSdpKgu/mejR3VpnHiGWLp4AMJIC/7er+zjs3tccH6ceVRfJENw3e
6ZZ6P2lOaS3/Cd7wzsipdUcGUcK8FrNPOgIEfvXRQOBNnFdqx4CiSB/yungbnVpZ
wRSxV43DIuvZns33kTy/kFrSKikAKnSCZu101uwodkanHptgD1LXFRWdZm1pIKx2
40JcgaWGOA13jbWs1lbImOmG+w3u+XcSYFLBFLXITnyHM3JPSOcOJLyXRTJmVnA/
NkkQEMHqCajarDwsLjQ7VeNz2hLYfaV7+CCWbTA+3wA50/6yWjeAw5IqV0mR3sVG
8STfrQUVmTiMAoOfIv8fxM92vp1+ud4oWN9k7hoyi8IEdpcjL2aL0OAES2XcF+mv
cu3fDbc61w98nXHTpLjm9h+7E2ulJbM7yGGt83zvdLctFa7F2lhWX6zo9Q9hfPWj
JNf/EGjM57uXifdvPk/KUqOHiClXqUPB9r5MrfZySUumOspbwLz8YVzg4zmvIc+/
WgAvdHp3lryeCDxMMGQ3YCmQxXO8Wzh4l0VD0VaZL02duP1tcc9rWcjh1kNDiYrz
xYAJjUyGXsc8jpJRoMP8KA14cCCfbve9Y21XURDnMKje663iRXh1l9VCcStjabc6
gVj8vpzYn6JYhyENp9dPIo08QiqCO0STYw1FWpMJn5EnTrTL3H3wQ7uTfnxCAiNC
gjsHfjAraMfCfBgtS208iKIvSON+/08TQ7HriLXUfC1Pd+Caslk1ECHLY5ZglI+4
su1vk1Wpe1aJ0hmdCi597V3LcbcqGsfaiq4yClmFnvVNEqcosf9Z+W0DAHFC9QSd
ZPep/yUazKsATrP+HxO62nl/rXIS2WBdYcXq+uZWO9y71GIVNDvLFyp4enGBcQpc
rtDvxUWA0sP1j51PSHQFk5HEzUjOX7RJH3EnYEC0GB6Sqva1i0Oe185A7Mnj1Lcn
s7JrqwZ7Xdka9m7l3v5KA8Z8HLhakOgu37PxQ2zRGA79k2Xgw6p5xtNywM7xV6MM
Eh+zXjLmIf9bA8RcBp2vL2EN3rBgJBs4fcVxuzUoUpO+diW/K583aYqnrJMNF3h2
bVMov3VEpgmbs6ENqQ75NfVLDOjzJJi8CZMnxD8NBqXgolugmlkoJC2JkRZuME+T
rv5whe9SXLU/UhePvZp2zcp9Y5KOZosGtYYzeUZL/HW2ER3pujhBulHqAm80TZcv
BkftHvxLRJIeAGSb4HCAiCi0SHA/SXJ5zjARFqRwIY2V2wUdt8lvPfcKr651WCng
XbXdIIVm2En4IU2E6sh8y2T1jmtMu3p85JAHrOOXvWSL781YFtb6rvLtnbfsk33A
TPRvtvRym0OrLkWoIyoFaKEIJPClbI2xCI+GGb/fF3+xCTYDa9P9mA/odb6R8c7c
TIApyRo32c5dfADDiQv9YGZCf7r+pJjgLwP4eJ5On50NWAsb51VB4DOtCQHvCp9c
fUJIM2E2imWzOFuvwVeCp/hIWuYWFNOLVUYmxcJ6Jx6Q3fuBu5KTH1BNV4HExhiT
EinRRILp9jxz59Gs7chSItJJnuDrCWwom8OK6jbzRQjW5ZqvJAJHQ+jIG7W/qJQF
BHMoXqETpk9NABOrYuZtinceoJTd9XTvdwPD7SgJngqgZuJkdAQYFC9VJhA+9nt7
5j9pbpRpcPj3hapo/hahHpJ3V87PrFulkVASHRQyy012Fc6gjOmGBkni1NI/MOgG
zFgvmbaPjSskz80yHqxDXQS8XF5Ti4cmT2CTnZiYmKYLIy8LDmKBJ3OAxgwnx2Rd
UNLkUNZZpvdfisVCzhWigadmQZpY8W+wlIlPejQ3CfEx6P9KtyIlnV8F5soCU2tl
1JxJaYk+Blz0lRIT3EYs9/h5nm8fiZzeFajjWCLwGouqDYT3g54KsKsotK9EtYUG
zC+Ibv4VE+0sQ/Ug3WuLV6PGl5dZXbD8akiHunu2hzfbofaq6meZCuCXSLHvyc/d
tE/JP+GSroSI+RlFBR99Q+kk4F3IfCl9WF11d/GEl/rCErpdvbITKRfLdrLQMFy2
bo2fD7pis+HSES5uwg5wZ+5DzPceamAfV9vYuVnxXdlwRn8tlic+LWidDYfFnByF
xzEaU1a1ujvsd2Nc2ag/9+3LHJvOjoU0j3n7sCqOPV0l6HkrQKZ/SOrFmvExTC/I
gA1zq1NYYJPhnueJvypLczq3MC4gSd86ZuaiNG71III0pqwMX3aTdO/9+BLQS3Vd
O6z3FaXNyoBhD384KzOk6UilXVK+gtGKljIvg3B2VMFij81P7C8mVO0tmyaKxgws
e3p2Tr+aKBFvVUdG/1zb/cyOaVgA8zaSr0fQatOde3EPOlYcSDeFkPb+OBxWFSOh
PGSeE9q/XqLdcjoGhurU5t5gLKVL9A0pkBTr5YxQNuaYbdp6GymEV8YWmzHD/7Bk
X3ZbhirLJVkt4F/2YH2JNqv9M3D/ZkJ7QT7oLQ/w199Sk1uoQnGKdiptRd9uXjQz
7FuuPxgpZ/U0ziXzldOWn4rBt034tICkw8x53QcU3X4D4PT6hQ6A6cxiVLaj//so
RcvWdqheXsdTxqAdRDoKq5z5QTefUPdUwLWUdkOaomAzRm37rDBgBpZft5rNuoVm
WiP1mgvvgXv8mc68NEMqbEks1PqTcb7LC+D9x1m6+k7yzOEtswHh67Bw1KjEaZuZ
828MElHMjaD20li8adIrpAeJPRvcawQYnOoYvN1c8xovSI2YQMRIqpQ6+m64qpjp
5NA7Rg4x/KclhtCI/v4K/8b5Ps6Vmj9BiCRonqkQ2D5rXEDkgYreA4T4RBmwuNn4
OgQBgpBbHKMt0Rr2zMrQ8IdvBA8y059WvyS2OczStSgyHbc95qKtDa6nnrzJwgtd
UK2t3fACD5clmgDRewoEwF1fGDjP5sTvmw+KcxqyQ0uwVJ0UD/xyX3HtucqVFHWc
1aHzK+u0l3WnLcl6hdpIclFFH6HzDjCCTgo8zUIyoleVtciJDW8rVMBO20lq7MC/
R5o9xqdDIo4aRnnDkJ7hCb2Of4Uk46MaC0vxBrJvcHol3qyGnKuDomt5jTS1VNXP
6YdxiWjzaGGv0ckGuHW8F7/oy8E0Y/rsqNMYSKs6yazw/F+SldmqdVRfhTwzUefe
0olc4x8t68Pv1NbGd1bjfoGQuJMbitFZ9cSdv+gZ2YtfFdif3tRDvjRVBumfLwK8
DHE7KGLNA7tc7nWMIf8T0Rd4k0Xp/NhIjJkahYlMwTyfozUZsJu7MmZ75n3s7Kmk
AftzRS0EZOHPXCdDI5InYuaBMSVbMkz75MroX2vzJZRLD5RDFz4brnYat8EGfv/I
IWuC5VVDYgvYYToSg+Nqgwn0XobQRtX3slnY5z/ZGI+QUDBf4h9xqv5FDjGTWCtM
49Tp5Pfe8t8MfJERuwJftGYJ1bav7EQqG2Y09OAhU4O+JS3n9z895Rz1Vo3puA9N
SPwJoLMb2QysCDqCMDhb1xmiWhuXSEptX5yS5/cv7UYNxuMQ5H0q29WJd7VXnnJY
mJ63DBnaNS772hyauzCScG9l0Kt+WqaF+60YEayVBuEZZydqHwfi2cAHnCWL9Dd3
yaFjNFER8ZtuI0OOXeb2q9aDx68q13eQwet/RbnY7sLa7rc4WsL6/efd6PT01G6a
UYwHg8z3ZWkWDjyKgBn5WvahiZ+D20ZikxcPBcN9J8Ibw42sxcbvY4Yf81QSzsOg
2sRwqkpuuHwC/+e4IyWSxqoUUpcwtMWZm3oV8Up9mgWcDwl5O4uEXYCRYWtwDj0B
Dqys2n9O06FeINkzQdMpy5yXd6Q0KFXOtRxYn91qbMP/jpx3JCXoLzwCEzmD11dZ
SafYAdICr8REiQHWB7y5tWjD53jxosC2LRT03DaWsZCoWBxtmeAJZNoxcAyr5xDM
btO6A+jF2ijZlMvKtBsUF8bo/tZsBMG2T7bBPZu1YNxTRU2ueUo/6GFJeRmgBgm2
rrau50mI/xFMJB4OewIVqCEhnmhJxFYm6ijcF7N7ZiBomcEOPXikHDLCwtz3omGv
Oehy7q1FJbTh96LvEgoTPvrNCUjPRShiyUOs3KYhdXJNSjr7SVgWzawISSSnWJem
5PwNpPQG71/0ZpZ/Bxmu6mBJXJlgLxXVUD037/mrkXa0JURKYRKJyuT+hUopNSeY
nxhtOuerkwKKuooNLl26DgfuHHxntj4GnmgroHEDMND0bTOe6uHY3UDSz8e8iwDf
emDKL/QWxe/7DGlJH8fAk7IlY7EL5VcG2k0sK1d4Gy6Bh4B933vCiYXfFLy1a2dU
TTZmdkIRGissUBPs0uSeiZTiooF2WKiKjfOIk4hTmcvySFoMX2VM6ghUInqgf8c7
n2mm6PNj4q1yOBnH+vhfLW+SCZ4+riEmTrJ3b80IeV9K7f2qoH4JB0/3zbRQa5mN
KiOxPsSlQVgLuk/1P9yLOKm6tATOJtre65fh3acmH/PkyLq+CJhEw7vXobTJPn0l
Et9wydLR2UA9MfxHGK/mg/J2e+1DPGKefvpCRshRSwCbLkGqTjvRNz9lEJDgSapa
2vmtwwtM0pK119VmFjqIQFPs13geRDMYyqoTpENWoq9Vl2IpvwDeMI/1uF+SAc3F
cTane7cfhcVkhLd4Iwua9fcz9nhPTVVk1DMb9Q3YBTLM9Oa2FsAaWZXNXdKN+kgS
MpvkI++y4vCJ11gXnPjAaPd3ZEqAd4wqzvSGwGrwYVoo8e2hSnC+Fx++SgR7m7rU
WIpoi8zGSyiFuosTSqRvjEKPkVaUcA8+6AUuVbtxLt1MZ7HCbm8KvObp61RQeRmH
gy1hqInpwc0AG7log9QUqdgQcqng9JzIL27TUkov04TWBBamrvOqfMQB4KOOmmb7
FCMKv6YLlNwyyZ6d9694jXPmTb4nz+bAYVcP6TFs0ed0TE/IhxKIEwEzRth2gS3q
lzVonOou+tk1REBdapmybhT1bWhQylhadmunsqrQRHOI5czEWzUc4rNkLInCjtnt
0ZU0S4UxamdtgPzQeLRCP5cAXuRoAaz5z74Y96estG1v9/jmh8aFDT+glSW2M/cy
/Wyo8skgv+eJZb/KfsO/kUtRfz2PA89wBusEgQ8sszX/YB3MzkYWFEXuFpKsjGPN
5pyJqqHsIfX1attalkZHn6Lea/QqH4pfPnUhYS32QPR6fnSaUhCLPMVjmm1mnErZ
QBcY4yDyIomHCaOKF9Km3XZ4yHQdzglmKBR5ujly4dhBvvrSVkXt8HpnXH7folLH
tVEc3YmPYNDujI5VUQwCRyNUSFGs22D7Gciw1hqmFZHZv/5PQrf7bpsVg9VqQhp5
Dq1kgmYTixSlORgBD0vXt+upw6wGyfZXhtzAxBFN3UiY+5Jmxar3qWeaeaiiBFcl
RcQEZFrQW03md5XiGOIbSFZ/rxuwyHmq+Rt+JjMWPReHzeZ0jbc6LtjP+QjlgIcv
yNF+E4CVwbgk40SV96QEvox78v51TyCnDHLQkI+vdQiDCV+hiL/B1t3bWKhrvt6i
HUC8avkbm1ab7QCoG1I/YbIAhiaV6NiJhjR354UXrjLb4XzSWwPueteRQimEmepy
Y91F3Jf6KV9zYdqt/pZanPqK4XJZ2EDbF2rtYey+QRMiOxfuTFpFglj0AwO1ioWl
UJziOF6tsjYWyGAvwuHziUgJ8CDpdxAxrxDePDIr7g5iTRa/asqkpoNYa9kTSDCJ
AFOydi8JD4tXdWMTkq/EgjfLEG0h1KSdUv65d2XH7eutYE+QRd4qAh/HKWqpmpud
xg6UYaW9hSuKg8hBeS49ZXY6E8SsRRGJp3WnyEwyYxrvYhk46dTfB59T2OOPmMyh
Qfn9kDA5ZCafV5N+nYxk3ezuenCYwCKrwhTjykkYvo+Qs0cc0G/h9tZnjJoJErae
WAEOHy1nU6yi+IwIIunue6ItLdKUD76Dvj/BYR5dS8DKgMMH2ESNZwgYsI+dl4a3
Hb1Em3Uf430trWAkhYCZ/9sn8akIe/caTyDJxctvueGe8yI1EZ8dlkbOlOeIKoz6
GOnZFs6YVG29ry0HFXg5PLzek2HrTgIjXm0JKbdCdxNJ9zs3sYfeO0t4iyptPGrP
d77//SxJKWuNQwzlE93tvMGW+q64lbYrIhnWz1x4mRb9rfBXuP68Ayx2frzhBgzo
zh1bFuvA/L/Qq6DJjb5E/JeFkHpBeYKHVPYgMCGpsHoeeQlVKVP0wHtxBGVKnVRb
eLh02+h4bVD/KIjHo0aHXy1p66XftQqE2eNscQAyO4pZHE8/Dl6TXcP/j5+PTMSi
X2FErQ9Vmn/pz+W4NC7FpfNXDAajXmKkEKf1V/qlRWhAszPr/G/ZgVnkkLiEPU/j
N2knM1dl9I8yTX/piFCjvdhBbZGN0fbEG3OWLEX9lSkzEm8tIgZjaMui5fM4nDAz
8SCxApHZdMlPtcS9+9FSczntkBQSxOsv9CaGkpgdBkcDZKv0S41YziXgpdubZ3QE
nd/xTtIyGIgrOd96JM/VvxpLL2D9lRWB+tVxnxjFyfOmej84fYKinrR3EfVNk212
HXYVg8aaxEmXBz6sdReGasKc1+T8hKDxpvLyyyi1g7+SIUzsUR4QvKGpyhPizbQD
7n98HZpVEMtYrOXjHHSKoT56JX8tYY+IYB28+tyNQLC5VFt8PZEbAYpOFet67ZIW
fVwj4ab5rbBznWfFxjNzXyVsZVuHMZZYelPgBBdavdL0GVOicgknmm1WD0VoOkOJ
J5HclvVQRJN4GNaGKqG2GpeskFjgjWaDcNrfwPSmvCOEl5IgB804WfSBoypcrk72
zZkuVKVLkVbypg8ak5MuVLEFkThjLYtrAYrJyZqC9HcixPTCdWhVP9KPyuN2ewAa
FraiI1tTa/T0BT56pCuDKfgSQWLdjemShtArQjsoW+IJXAS8GSh1aUFLacyzhLw6
Iz1uRHH8aprBF5vy0Ep+f8NZHl88YOeeQ6FvEjeQBwB8mcYEIDDJi11q3hEjw93A
0RuSZsyV4tj/BfoeKY8EtXhfrGp/De72QOYVAT6rUPAapD3cz9B6FY7I7GSRa8sE
tHyDOqU6LOVXh/qcUVxko/TDJnY1vdImz3fNsEhGqjHLIv6sdOD2TMXKdIL/q2YG
WDUKtImHgF5ijc/Bybhmhc7uPEx2oxCGRPvHl4da9r4/a026/SFcMdE74bcDh2va
60QS/pep/yox64vYvExchUhyLhDeCzkzuVXvCAsmplBCutls0kGD3tBR5h2up7K+
+Od/Vrxb+VEgTmJ1C2eVaK8kG1ObK4wMeLpihXeidhkzo3GvC7V6ZLh/1TrBuJqR
JCSYpB0sEZdRDyf6mZO31zdCC2Fm8erKO02g+TFaDTnGqZ6ESn+UsCnNekpkTdp2
Jpzn4aCmsrZZMWC0j993HD6cH3ZxMpKJyFvgjfTnIPgo4zRwLNvGcqyXLjBKs4GI
mVJXuNp4ajMZHX694xgfeSGhHqs7MgXXrFAr6iVmrhGXuxMaMXMKatxhGTuZJhdu
bS4QsRfT+KYJssFXrV8H5ayIylB/dT8pEcdsiJsEN/5areG8RlqnkR3ZBcbRJWy/
dtZ8QXyqrmw7FwMg4zzVMAKJDGl3Jq7rT7zxaSBVEdJaaBRpZckG+PaVs6KM5VN3
zRjHdD44nDOUNmcSKYCsKnJ0ym93sgyTapmFfxTbd3J0ag/VryGmeS0lwl4//3pn
XPyTwnhsX5OdWJBReKMaRnOwbJX/E4NIaoQQ6kEjwsyRw9bngdASpyxPYarc4wXA
hfxE3jqzXndc5CSsAtwgXkb73G8vYRLU2IrmQuF6t+EA85fuxrrzdClGtzT+wVtA
0XDPaoUVKO21IOwXFrDE+jopkQ6PfN0S0dqDRtsT2/Y4YU+2ysVKWwYzYDGo73cc
x+SrT03ItIKoFjjGSmVxASZF4wrKKJgWrBgP+FdgT16bIR+q2qHnm9QaSszmr6yb
5uKMulp0ZT9GEkNGSoU6YsIrXWWgZJcq0hSr2DwuuEqPmCvlJ6CoalT/pTdeFb/j
MTeOqBfj8fyA+VrOD+URmgficCgvY7HvyAVyia6TACuQMFszTf1awlpL3ENdeSMI
XeOOdoRjYhRlNmSbOqdTTo53GevQsR+n73ymskVawLy4/PkXv2QoPUobNOoBGrTX
2etUQT+whDBKbYcK9rKqgTx8I57sU7P557/+ne3le2VPo5fmEqSkgJrESaSW58cx
wbFs/M4Ii6TVzGj0IwRbQVeO0XeEh2VmWXBB57GjP3uwjR80/jKg25hJyLLReSyH
WxLJhfvHgxkK0B9U0l0byOhQN4EywDGfDPbyzHzcnGOa9WRArpk8EuLk76mnKSOw
TNg2/5FCmfgFQtVJah5KB/ZzKLAc9B2/AN7nDW5caPpaMkCpCmcfbXEeUDtJdKuZ
us8ZLTYbO6pEecbTGgPvWMYJk84lO2tx9Gl4VfiGhMo7jNSCcu/hqCALCG3yl9OM
KxOEqNKf9TR92jGw7cB0Dwy02+TxknolnZmkFr5WW/Lm7qNa3dDbpXtnYoF0bfXH
NaxPzGjWldXGTvS3VuJiApPyBW88sWi3Xwqe+IjyYQq16ZLA6PJVB7ccfY3QqltZ
22F3Hx+X0HhEO8C3/cOl5adDWiIYZVoCoOn1PJMxaLH4+wdjJrT/pPFupSm4QuiU
Wm/4rOHh0J2ivP0pFMojVN5SJjjpF7vimTcUQCm52PaDvJybl04hBZ7uKjuJYir+
6Zc013FLg+pOwlpvYzptJe+QrsfSiKLs/1CN8MDpfQuilNZe4uQwgMTNqjh2/ADv
JujKmOxG/HfCr1O3a6dyJDHBLfCAK6Wj1gBAxVB2HWAeiQlmx5/fGfmLVxghZBu2
Xy9ZdnQ/MNHaHSRJwOd19HW4nDT6p9k2j97mj5RbLjiqR6NoI0Sr82PN+MdS8Aen
kiJXIWDr1FKLw4Wx8rVGDK0rnEP9TMNHVnhTJ5mAGBUoqDRmjccmVn6Hl9s5ymgY
sJ3Gmf7Fcty2C0FQxxht1gvzSuecjwLrMTxITEmlJcyOECpZawRmAdO+hRP5hKfB
Bx9sW76NhrlcUSjXCGU6WJnhaXgB/oygRz4mimJ0jNx5QjmKq+1L58ITzwc+y67D
Sv4SpG0e0CVUe33L5qbJ1VtqFG6He3+bqqFljxKgH0aP2tgMlQq5X4d8K+OR9Z0c
xeOmrgk0fbokTNout4lzdAp5MZrlq02zhASpNRxTkpP8jiolZIPPEMU2gRuiU6so
NnKolj1SvV4mcROiHBGFB2RkbFEzdF6a0TQ9Gn8HvlX1wTSq3SBpUbVRCwxKuhiW
xAvvstGaOBYuMZSw+FaqAkZwfi8YFsqJy64v12hbcXoqnRZyDIDDL++Krt8Irpy4
fLu35kzxa/b52b57LJU4Re8ZprhbvgwtZYiSN0FJIXq/lnlD5tifrC+Ihhky6N2H
adDi1NKyK3Q2t0sm5KOiLainkzOBioNOM2re0yle988hynUTD1wHRv8pFl2RXItK
pnRFLgEaPguy2x0N8mpz0cVkZJDLcIjZwBN7iKUoJFnt3YG0/n5rc2nq3DL5nkgE
IzYsDqbws42HtMqpgm+lXoiBwV+TULFWY92bjLQg+v5s+GJrrDpu1/iR+nx0zvNb
tqLAjXJZG2DAd3CONTqsQPXkEQfwCVjgtOU7TEMlSMFcDH3D2/pycP0VmBfyZ3oh
mIdzExO5q9XaKjY03i51J2rV6WqrXxFDGFbGY0eb14gGdGnY8PiVOTXL5JV21v09
EIMcrEGDBlTJHnmHQtUGfhioPAg8u4i1FT3n45djYThhqEI4OqaurofntmpNqI6O
YEN97f1UQIloq9Q4nLeHVnQafU27oEJbGwNgMCLFkX8aznXsKcNIOvKeL3UX3XWA
vHsMBa7dqaoufqs4CiOEmwOw6oeAbFro8w5nC5tmVsxJCyR0CNnn9Wewb3W3yqvS
DR0rakQ3ztwav83X7LLzqPQemz1pClocudntpOUIhJ01j6ke3n/i6T/pLz1Midnc
giI8/S0G9WdH++Zl4XjKcqUmA/XES1H1GACUuVwpfLe7zRqrr8luvvnYEaMwJueJ
QgErxH3I3/UtMlQlPPoOTZAMtC5M8381HI49yxpbDzkY3qB0Tam6upwVLUqPyI5I
cYYHnsUaVzr+IKOtqgs6c6qsgCbn0ggI/lhO06SF/8nDl55+fidX+EqJnriIYLuT
kZJDfmDe6JtatOH8+pzRZq6OEvispByt2Q6wfLvfd7H0YPUt7OWLFzcVPxJi4pxN
gjNVyuTcdZ2EI0zoUqpwxmEQBITXHzAQCiyYKW7ZWoxirLXe1YIJ8hvvqJIcWjWH
5iu13CXDFfyVu8QFWwlCG8ShmjYdyxkQpIccK2kUE8MQtkwax/VKZu4drlqBdh2+
nmMfjQEnNOnCcKQH/Amb/KqAE0SBz0B9uFJZdp371lZUq8FrsXpdwpamJyca29bE
iHzf2a8cKY+9+nHlNrR3F91zyuDwSN04D0OkxPdF8QY6DuaMa+UWW+sQKuSPhf77
4oInjEzjhhaF6CKk69iizL3o1a7Zjz7zFd+Yi2u320Sx6P/0hAON6Yvw5UfYJv6a
6Dp8bts80Nx8tbhXVT2C+Xxcy+glAZqEanays8eTguZixpk1gyrDslCuRXjLg7DH
P4oibBnUl+P3KKKjHpsLeIodIkNLIOVNDoEJM43yGJkKSu6hefsJXirLxl80qucU
pApM7gHtUXdS62yh6iGggLNk4tSdPz1FSESQMEyJzf1+eFn0XssPZY5MwXF6A7DO
Z1VtSY9rUmwTAzcsje8SXc8p2qAHbPtm7GD8/2fU/7NaAiCXRUzPvOurr/CCi4+n
ysujIEaXjSgimhi+vSEN4auiRYUGJLJPgwpFwUSpIeDdxi3Jr2ZpL6jWwrVvo/dP
2Sg7RfRCXPKas4jCIacaQND7JK++kXq2YFPgw0gFOnbLUleL44/ZUDvavZlI8AMq
7Ppv5YiHBv+Ukqjbh6JADb4gR+qk4Dw+Zm3HqbUlarw+YEvjtWLqwciU6AnEithP
rOqjOQV/D1OiiiuqXbHE6QfBp0mRmfQN+s6CQCr+H7eobhVzggSRKFFahS/go9lt
wWzkENxZBHb1j9SowiwjS3SpSX0bV3gZE82od66BIVCiHrkiS5QvFIjiO877/4lU
UKaPY/jekiCufXeP83y7IWXDdvaqfwkhPlTxFvs/WAu70/ZL0ZUtZ5eFwe6RFrtI
O+OZ8yh2MO9QixRXRb7mARFKjoNN/ObWPXhVHrjOKtLiHwqUqXXvuBNJdYiBeVru
3HL/92dS/Vy6KOm8UITR4oMLSAu/cZg/Qjl114CHWoI1FzllMBNpgPYD1WFX74A9
/6b6nu8JpKMJG40v6PS7SPqU9IetgtpMlgzPthb3RvqIEwhDXZQ7YZi9PIU/F7Y9
enes/eGlX1jd+F84d9rcar+WYmdTce1F+MiWxUu0r8OSptw6hME5JC7QE8goHNkM
tH+xhw2qmHn6+CgGIVO9o8HDuCIcZ+JlQHHKGtC9sHDlc0DquiPASVwVi6nVXWa0
CDbcjMbnUmGrmErWhOPkItxdNAO8oyv4y53hemiD4/Q5IRUEv9SULJlf3u+Lc8Cx
/W7wgn8Bv8ctCRhoueaOmqOeS1z2Z+pgNKP9vXSj3r+0tDB4h8p6hF3vGobKFRLz
7ASItVrnI0sVpO3Cbu4XXZ9J2fgoseHVg8egMsptMZLgt2rU7OO3g/MNJrv1gK9C
8dYgCvmcby1kdobVp2CYHskoWZO5RGzqG85hqp67n1fPYbnw4pETJBHlZa4cbKvd
srnPlZq4XU2MgUan+6NvaisZuvd+SaZ3tYEvAfD5FD83mFtMH3u89jYSzMO2W4h2
VlnquTCHJj+PFxmsHhy6hKng3P8AumWMFRA9mkeS0UkP+wI/3V/0EwvP8ou7WiOm
R5gRq4McnTUdRh+hQJzsEg+veBaFN1L75zMdeUwUIOt9pUkG1Czbrv7Qkhe5aFZ2
iy8p7CKGTk08ez8kICmSJuiN5VXEW9+ROAiqaqpS460h2pobg1lwuqLNafaUfeOL
+x4c0uS6SpqPklBIMedGahreu4daK+7KER+NV1EFzMrAbtkmPX0g/TFBQ7uK3Jnu
cpqPsN3YLiy8nt8Mz2/lwo134HD1dQJMTbO6VIK1i5LUE4siYnZoz0QAGiExfaT5
yje7jQQ0Y9+6LbEaZACI2cdvGYKUgsKuvcFYTkMP+4oyd4ZR7Lq7XL52+9eTZqJf
KGfqOjyPWTJQQnwLAHdUUGXaPTo7O8FKjoPQso82KVKvmX49Zx9nX4HeQns4Hu47
TYUiZQQL2jz2WlCzxep58JGOzEDE9IuDl4A79dsAycRm9j/3rjreYwvFmvVIlvpW
JSf0Hgsj0JzLx/2Md5fKshkssFgthhdPyaUhXmQSongZulbUM3/w3Dn3re055tjp
W+bDrJM51H2dhC0OJY7AJl3DP2KiMBvhk5JRFVIrATzK9FGteNShzW27ub/P15p0
OcWmGzxAr1e0Z5cTodFFKQn1jnkNePZQheLtOH4Xn8VEPaUK4mhVS/VmGHmwHo4J
PVxszU5/9wcAFngWHU/yJDwEjvlvUt3R5J64LQlrAne2U3lMhwrKFAeehhjbdxMu
jrMyZ6OuPiZB7Jx4Tfk3k5eqtVfObZBPoWWfCAFSTriHIqbMzwJwOXW9j8GJJapb
07o4bAgUtlZ92D5qLgu3tkx7V/wIvnHvPF7LNGHxfuN2QHDXV5nEMSQpVJ47Xk6g
+J9BDBQ3tmM7Wzd+swjuQPMPpAfORrfLBoA1yoLC8mbEbqAVKoXQcjwasSX8u0ay
7CdTpvdxuNHXYs251W1Dj3Kc8f8F8nAgzR80eE04UBeFz82xLd+kv42TUGFdYI1J
dVCN2hsHzS1cu4XouH7Yis8Az7vAzB3cil0DB9UEUPVv/p7LBdeID3dIlqXivfr6
NF+btv1mefLa3qZOiN4+QhSWOMw+1FEqe1CFFNT9ILqY0SmOvsjoaSWiY8i+Ce/q
TQwnHkxFKROCm1QiSAzW6QfSQ8SitptytcDgAJfVqBPM7OSUvt1go61BCvGfG5t4
WUTi7LFQng5SzSgRq+GFLRma5rvwBCiBuIk2UQ81bZxCPhSg71wrWG6ATzgv328q
ejY7r8RMpXaz0BaFn5GoiUX+dqIHtQSKqayeiEf/Q6MvC7AnTUNAO3hnqhS/Zm6P
wo3B0F3ath2MKnWuP0shred0699AVgRxpzdsTvllm1U3kCr24NfZsH1v0VAdVl3C
MVOWYyqxmLRUk1kdDEQ/njyUxKXekBQzmG/yokUnwjiK4URSDhcriK67VjQxk2gl
ygTt+KwuKgaRq7YC4+TNeZi/VCd+oaTCVydygHzqL0E8icrSIhQH3y3O0W0zGZax
CMYZnAWXrOl8DsGfvxJaigg+eFrC23HD+xP696Wr83iZsmL41e22OPI9xL4vws47
zjbjKDnROZGaIlaUFs3CgUkkB2Oo11up78AWTPxfJSG0F5bWAwgFXKhxhIBhU14k
0kIUSz8XQ3k4lLc/Y96e5V9cuxBx8xISLSpL8Z9mUbPEzHLcTp8odwoOPKpJK2M4
lgnE14ah9/04Lypv2Qil+OUYryhabEy+0V4dKt2Ive1kdjuPCgymof0CNXZ6+jcF
FhcJm7bwijIKS9AWvU7IkqnRtGzjpzPOgpPB88NXneo6UfqXslprQ2ryQBrZeqLo
irIihlRvPvqXXpYirO9dsq4c//ycJzU5K7rwvlF6d8vBRc0uzRTO61hw2eNtklJO
4x57ytTP9be84/Hl3EHYcDGs1MTv4f8K5log6+AYcaO4oLO37BTzNwq4+uhuB/R0
J57XfKb6IxATw1V0t42ZUHuRjHN8dv8ONFjpssZKdsoiVL4I8NCKehy3rGwrIJli
cc6apQiSc3cDybdwU62xKsgI9+Vgb4rUY5q7ziSsYDyoFV2gtkEJSwmGYu66rk5l
FqHU9ICdYy3kh5yUCpS8A9zpDqoG8Mh5hKagVeJVCFv+vnKahCfg2t7bo1aVjHl9
noe/43045fPSgqJx0wiWnShJal08Gd4VQI4IEplMzOCZfhsIXlikMnvs+l9Zt2OW
DqPLMFebCL5iYhtSJZWDMtQMcWEN9AbrZdFz2YPTqSEaLyo89x9u4dUiUu8X/XLp
Mtksb/5vP4OEuvq0976Fj4L/bI8EAYjXpKKzX9fCA1pxcMw97viMUVl7tmdCV9+P
Ws0t/JqwcVDa1T81clm+hDX/EgwJHwpJ7YXSJ/Y4Dc3ZjbzuKlsIe48Klccgk/rF
p0jL5RAO+7d32wggwhO4j7xiyIZG/08LQFVmajNMg6UwX/+EUplkSg2uNCx+UW8+
dG7RaWRONixHBR4OjUJUMKkMHu4OXjyC77rhFOrjDwGyasMDBt1kf14Al93pSeEN
DFrSstxt8840U//4fladtdDR1A/2C8Dlt0kh8Ivy4QB1Ok9ZjOzbRPaGyl5CEARi
KksR/2O5JbrxF2jyzmzZqcdMjFTx7ieCWMbMPqqoynylAXCF1jMaoziWCcTmuQiZ
w6/OULQQU3vh+bBJ4zD8Scs00Yrnn0lUN/XQQVc8TICBADnWxqgiScrVYPWDZmyF
7PRE3NRK/z1aw9t6Sl8Woh9gIcqp6qftQenm7uqBcVOWisqdamxxEKixLAia1TxB
fIMbCrp3OWmQADfm3Q6rIPMIjZApt3Kv7UB+k0qgQZd8Q4ITfvJwK9H5q7aJf0m7
JKI04zYYQ7PSDR/wixXjI0jTkfqtKC0E0F3mxj7IV/KE3YO/OZsLfv8bv6ahhnXI
53WFVJv69hjvJE2AiIUKcKp0ekKdh3+7I5Sre0tucNtag1C1j3IR8NezyohdjyDI
B+158hYjvDGdju+q/XcyJFh709HHlKl9E4eVj3e1vhj0a8qcSWnqHLFNxaVH4ZfB
A6goGhwv1sq2UmWETmY6XMv+IXadoSFKEuKzsIt3ns+sieFahPvkMoEQS/yf/I8q
4ptgBnW20j3unek+1lAvHrHZocfvuptipzfRXPJy8j6OUx/4925DrxHS909blcpy
dLKNSF19lKXUfN0iZ+2tp+6vPtG9+e91SFjvT+4XZmVLitcbTCimu46nVWWWDPUu
4NF/geQOqu5i0WOagvsajdZZ8W8/cf3QIzZ9YOHypon4HxmV1WvCF1msjectJDrH
ZLVqUhLkEhZZ/lcn5GuqR8z3yuOQVuihCD+Ukv964b2qWTI/lFts0A19OAe1NS7S
1ZB8m0gXi2Mf8K/PVldU+7aRTaJkVCYDqwotNMoFtK+Or0jPFfvy3sjbYNsp9OML
qWRJYbOjTycwlsMJ51UTlu88UR6Ayh2PDI2FhDBQja5tdCUNUXp+yZ0AHZHQSNbc
jJuq5LS4mJJI+unexK8G+KQpPwXHToaKjrYz0NdeYu4+eJnhuFBsbfkUgR6d5COC
mMtIRvKNxx7E6i9TqXGApcPzmVngWyMw6IK03SMsRUQThM4kvKzfJG/x3QwbMb7n
80bH6SSGWoNL8K7UvR0gcJc9XX2cQfYkQNZAk0jnKuKABP8tjJSmnmMBqLnIRxmd
e9Kc+wiDFrucugREZEKdNADn1uWyNNSLTFKWMY0FgFMvgh9BIYbww01RbEZfB0Us
NbW5pK1LjokrrOWPSrb8jqQcIinq0bRCDCUEd3HMAeKNHrtIqwUjrdAsrtVfWYau
icAW4GeUxyrPP0+mw5ZTzQzohEGV0ZYM/O6/jaJdSfXImb0FgbTJhzLgHwjh7DV6
tDpPYViGf/hL9eSkueDmZrzzplN78dnDR55r+7JOy1cRbP8wwhgWKAaC8LtsouCV
jXOeL0ZR7Z6afWWwX6xL+h6U+HPrFc1IfdtCNERKobDzCrbe/7SKSJ/Dntcvqih8
GUGETn9dNgz5YWV0TTxu4gXRn/r5hhLbhXqWGL9iMaiYACpBDjJQLdY7A4c9JBV2
7yYW3Tl5Nnu151bAmcFcQWZMG9JnQCXUWUFXWHxESuWckS7pKME29am+inwhX9Rx
KCv/Pr6c50zyY5vo5Mc0Tt16sgdSKfdHda/O/0dBZwUtqldB6yMmgan8nE5UCtzk
GziD+KBfL2RtHbNKwnuuG3yAjpgx9tzMIKB93GkTVKSoLNtMTRykm5LnoEczGwIT
w6ArG+rZ7NOOqNYOiw9e+PfiQU0AXZ43jOlFfdrS0ZUm1z1TxE8bQ91OGfR6ds+a
Gz7QqRgCk9FYJdCypalpPoVdbtCILpjUXVayd33TzjAdWAwXdX3JkgvdsWByQREZ
oT7zJOxZGwlrp7leoSq0MGWG2u/HqStDN0Yu1jCn2Pftlk3k2g/gMvndxHYwn8yo
JlpAVGW3vwGNxEd2+fexTHVridEG/UFPDvy6QU/1KO0QZVirWG//sgRdz8VytP/R
bSEeDKFEPWW3Q1VXH7Ur0gdlbTnzz4eiYsL8es5VtIMiyRMOgG4snjvQ5a36nxxg
Rj2MpsSlbz4hrhSAHbYBUeiSIaXUUFuiL/zd7Znle9OzvsGh5pc4FctPJUo4SPui
IbjEUsDvPSYNLJQAtKXep7MOz9wPK0TDoCmNZmj7Q9qr74eNosz7CPijHAfeoIGO
8TQkxjcFfp1S+wH7w68+fg41uozdXE6qF9DbNDmZXc/EArbKS/m01a1NTYrXSATl
D8qq5ycg18/WLSUo5EFM+WWxlFV0LIxES2tYZ0b4JDCFEsBuf2vd1VyNinOScRLd
ZgLP4YiSi6kWgDDYTNfReURBPTzuBVPfSzg/A5nvYgtzCd1adAipM7Qi8tbVhF/z
DotbD4uEn+9IOGq+Wr9jniVuZCzaVnGesKg6m0XvJr5gksvE2p19icJdF2CitWK0
hV958cKSepd1jKCR4N6S94d96EgwTuKRgHX5fFVhcyCpzE5s7JSKpstPX2wfwCwk
9M+cllvXZqmhBcMWBCg4AdtZ2a5KHlnrOPGVYal7zM/A/V9kyrS8zvGVgpCFdeW3
tvTyDadwOXFbBarNDBS9ryQ6KJGMu5OHorvCjHnSEbNjG2Ov2AYTINPRM8W5iA5k
YNIu9EkEugr+9Or+XaEacEncesbIs81ovmQlcZnxfS1pm7lU4AADz07B7NBiIXxB
hG+GdjGJ5GriHOYttTzAfGtwOsquE37tG30Hcupl4SJpU2zmV8hPEGSnaH+B9aXa
qhFzI1PiPs2g3yDnW9N7HUUDSIV9RdDldOQPTIszb+uK9Avl7MtXIZpraXZ3X4ff
/EuTz9LnR1B+kHVBUPDgF/d3S+sn/s1yr8tEkoAF7tjORb436gvqX653Dd1EP5Fm
ps5dic9PFWYljW/PfYJIq8GXAbct5keGpw4amCSFcaF8JEQbMOUEGBjoXvghsMIi
n5RMkkkTrAeD+Y8eZnJ52D8ymAG3TzdxoJAMN4jiJviniyXAcNQGrlnyi/SJjQB+
6wdQyLv+7CwWOw+roaJWRaJ1Fv4ri32jWjkk64B6MNWrcgRYZjII2BmncNgPvUnG
7v5428SdOv70qc8dZz1LFp0VMvMHseSAos+ZiISuRSrEJIlAQU9ygnfO1c8mg+9U
qysQTNxGgg/tCa7/i6hU00Ovk4XZRgaoxJo6rAJqTy5Wub/aIIFF1pDEICiiGaf5
23fMuX0pQoPSmB/3+NMfTAcQ8B+BKYjfmOq6Zt+BbyscOEKJ9J/sjERaKlEXTGs0
qX2vmtCep92iMjZgNchvKEVo8cY+stZOHDuHkw/zCLfNuoOtjHEs33Y+uikSduri
Frt+A54kmWP7S/gOm8ZA4/kSeIB3vnaSS2yq2LL1IYkLhxhOasiL4QiG7dMN+MYq
bfiqwpk5twGqIYG1zPpUpZWbd9nR25safrjF8PAbmyBrkfWzmIcNI+b2lpJvnUHd
Qgunpp95NG6qV5krEFlEteVbgMXtHA/RFf568l3PO7DZWTXXxGyiR5yyKB72X/mN
xmz2M4lxbLPfnwTknZFOfd5hBdDFc2ADQY3XZkaxEEK2Mx5Or3AdqIYCvHqjjbPR
fnEQIuVzaE7Dfe+y9lW+gfwjGAS5vZzO4NCarr36TlnaEHlI41XqHuUVIgtH3jzX
4Nz/G4bA3pcUGc4GEc7QygaENsxRIVKw8v2UXwQlW+Zou1fcZd8/7WmooGopvCoK
+FwEKnjT+PZzewZR/HBnXIPeUTiWfYBAk0JkGehglUZP6q89flnvsf11G/qWOeWr
bAUCttPcreJZZ8ML4fgd/Y/UJhdXnUtv3AXb/l7uxoWiu3l6GLSZ1GFfPWmiNMSA
gnEOb4FqVDW2KN3UgFXqhPmFAxWwNk1b0+Wuhg0iUcRZ5e0A5fMD+b9lSuhro7gY
0XUGurzFugeTaJm9z5ayoMmS7p9/kp3lxDbgBVnjtQXCp0mvrxR2Y3C6B9Disj41
hQt4thUvK2AkwdmeDnDCbVdmh7xsUF4dgc1HJyKcodrJv9SZCtI3o7zjP2WJ6Omx
+dNhHaEaoEf66LTg7FPSwpUwFXgSKGJ99NmQwpiGYO9ef8V5oHK8GXi0p77ln6+s
tzk4oTTm19uYbizldlnGKjgNqj3YrVHBrzZyeNlx6gQJLrzL/Wc0j0atxeN1oQrW
xKZOpOep7xPNiwmpxcBVm4BMphDegdKP+tKNFRbiOu5jG0cbJ20kpdcW8oFbjLKs
3OoCj6TxiTxDeitboqiqAXsl3rq9JBxROx45dMN3njFuAv3h8tnm+cTyahfVhAmn
JX4PwRanLannxAC/4DtBjbGWT3pDtzThbvpRjoEjePRBDdAytVgfyQ2P3Q/dmqGC
su7rM7443Zr+zl/n1gE5dR1jEuyE1whamWuUS7skMf5GgU1F0yO4RUNfQk7ULBJS
s9G8FpV+B4L9o9PxSQ/KTgFhN39U36mPVb9J/SVN8Pm/SMFZLieYcNrwHZrZbDSr
tizf70imFKNDFfuiqt5hu1wE0VBSCzkJCCjZdD5nwvPPbR0fg5kbNbZnll+9FKue
favEkDYRfwGy1x2i3otaCjRjAbDaKmYceG1iP/6eMbeG0OI2LGjhF64q7d7edzT6
JjpbqgnlJN97CkTnPL8hoWRY5qTlrxDHzZN4dIRFMngnn8oOk+x+HvQwjMjfqzLU
0/XJPZqJr4Tx03r5b4RXkI6jdZ5wmNT4qPO+SexiICBfW8WIx+5cQM/O4mRLzEDF
sXhTc7no1CQ65rH2Md5LMgUeXViEAkxWywVrHmRX8cCndvCHerxG5kAfceISIaJu
g64UijKVXurHQKfvR7gIZeH7XHbhphPfqBjgmBDwF61nRFuOQDzDp6PGZkVo/Qij
xw9uQPLBgJteKWH1elh5On6FIaecRI04/ywGLDnnr7F78TLCYxPxPXBL4ciij9Ri
Z6UdUpJpA5IRH8kJ1je1SUcmBleN+2YO84iKPPBcbtqb6JMShJd7lGxUjvIqFUnV
L17RSi3g3tMw+dVwrAAlIM3hGR9KKegsBYAiCTeUKF8cWdex6dTT1nZjHoCK3y/n
FaNBerqJZu0lbfNIsJMtSOz8PIp3OT/65gnHDEqpoev4FM+yaEkgZNK0w/AZa8OL
Qjr7gfGB4qKThS6zjX/co3zGsBhxAVNaO99kEF8tsrrmA4HWkfzoOzf58g2xERA5
BYaeShSdupTZFvOP6sFrtzBBrhMhcEQOQ4ZKzgmQD5BLDZavmFGGChdCIaOv3Kgo
Cfs3AXo3aeeqARDU5gP2bWu3DUkzTI5yc0SkCWckNE07nLWeX5YFRbM4MbVZaTN/
wvKmiXsWMvbqNf/gY35ItHRKBGQfh0giZ1IMZ8L12zW95fYt282ItheykIJqPPsY
NbJ/1eREEDenn1CPHv7XE99Kv04gSypgGBwV3tkPYLxDX4vNkSaFScc97Y+kI/S6
lpi/WqmEJtrZcj9e/ObI4JeGjWwqKcdMjC7fQGC0OvrJ/DXPo7QN5kacuZoXOiM+
5sR9Jq5+wX+vRQK88JmsYqR59b7UesGMPuKXzFGacY9KfaOdMOFkuAAMvg5MPZaH
lZntY9RQa/kzRanCRlikQDtbTyc9HPC8qjpN1TopPOCQODmwJ9BfCvXnQ0kpcidZ
oEZhEKA4TxnY76W48hPsKRuo1/FzjA8/b9vS0qp4agudr6c7kkC2bDttyXJM/Bjv
dNvXDrMdpIxKedcruydsch9L0FAWLlvdrcbfVe7aFzz1lDn6JJVWTKfpm2i9AOKL
0SeIzV1g7UFBVD53Jke7eQuNuHO5ckfieRjrXV3Eg1GgwL+u6BslHJwhOqDGFsJl
xu1E7xb8e1PbIySBjHjJuXL1sTpxND3tfh3b4Xu2RQI4MzDjcdmCBmdzpDvNkP/l
I4JsWbm60QhKoJAhSdgDABwDIyNw15Qan/q4CZrFd0LJ37EH3Vk3CaNPrpe963Ym
kUxiymCkSkd5Arbljf7Zwu18zIwt9Obv1m5tkdEGmKRLBPU1iWdaEaZlofLfPOIG
rB3YXkwgVw9tQsHxRPShUJjPKs2LxezbLa92AW1+QNkvrxzWcUEwLPQMPTk7mbQ0
McYiVekWPjQv2YWi/PX6pnoNKpkAoGhJeCiQ1HvUP63lZaLKC3og6azvms997Z9A
PGjfeQ1SUXfJgGE1c031U+KBSqu9kUIo5TGUvajW1HZgli/iGgEKCP565iV8CGbp
BkkYWyMb/jpKBPV/1ARKMHFoGfTu4vuEDyajk9JNKsHUBh+IUa5ScVTcIrkrCx0q
T2VUY9ro+ODb7r9lKIhjtteDveB1NHWCMrg4ITxXXbsOM5sTv8eMSDIUBw0ocO92
Ssci+di4SGU+9sLdePx+D6ZF9y5F5dYLmKdeBXwGvxbfohYhPLQJsGLWgmPo0tqj
EWjFSgOLpX27coFUHStK7D+Y5mhOOZcmSYuJpvAcI0qTaUa3FA5ehWFpR4N23uNB
fP5RUk4/oTCRK+B/yh4G1uZB2p2YwUr4juSGHhaEE3nlOCTkW4YoUtLShgLHvW4U
DhlFDkENU7aOrTVIbMGhLtKzDypnDxNXIM3DCdKjvjmZ5lPPONz0/wQ7xD76X0Wi
Rqlr2v4+5Ihh7a3WfZdod6258uLVV6fDS+Th5FhFHKERlJcsTZ3a8+9v3WjOP7Sr
kzxJQA9/PsknHo2l12PuB8hjyofIu6/B43AGHfKOr79Aw/2JQ6CTnDqihp2wVHxk
WxoSQkqC5umEd2rTbg9bp22fvqTZM2mqX12RhEfP0nn7rRe4js7GbtmNHTTblcVU
KMTyTDdMnS2rEQlfPeGzro6+Dcq4Nq4N8lOH4B9ReV3aMsJDSM8SVMRTUydE3CV2
s3/kVgQZdOqtitF8pxKesP3x3FRh1MsOarlnVatrgXsdU3OLV8QY7n9MNyWmp3Ku
2Tf2Ob9cMiHU1a07RSSSEzwNuz0e6eH93lZbvuowQ2D1YJoeBkQ3cof1FA1rdE1T
0vOmCddhegUDCehIcTQ7PXBUkb6Cv1hu0mAqa4g7lUCTEAsLLaG+1ZnTrNU66lsw
NZtsrD1mcB8OjD6DyCGCwvh4RQqInq2ujjHL3KlWMHaDxxZz5E0wItqRFbAceNAy
3bm+ZFvwV1UGK3vy7xiiy/Rid3K0MSuFMgCUXbCCwCSHLs4/WS1rThHWmhFxUOci
4RLufPASLidVYB1xpKusLzuIkqZ43bEYSTq+BAGjpp2L5/EzyhaB3Z9BLe/PSYlh
Lt4dDAoC4kwVPd2KGkazAaO+mBYF16wGVYusewcxap0YNKgBzskIJVs9T623X1tH
zwgUi0p/42QjCfL7Am/S1S0wYAAMqP3IYgUErfjfKi1rfdkKimyF20sEt2tLVMNF
H0eGUOino/n1nhZ9wDyT+1tP8tNL158IkrRwvPECxLVl9AjAXJUulDSbB6f2u07J
nSRkBdd09I2JqFnf7YO2BDOAX5hNxkNI2Gy/FZ77mDKntk54YN+5/CGm9E/sJEG8
GeYN7bdmadRHv+DTqz0ZCVkVon7D+pQ4oBGOB09/q4CqiU4jtxDj8cLUNdAXaA19
pZENyYPiHXFmFj3uF8Lkl0eH3mvif1ra/xKMXF91NxtCK4C2YYqWOyh4M843q/Rx
4uFd8a+lHd9k25P8KPg4Ht6sfgWNLJyf88F+qE7SeRdrXR0G0E/alL7l6V7fGsj4
g6muHTXnc4r+fkk4AUnhYc9ecltle7xJiw/97moMS19JKqSbq069lYrb1Ci5IiuB
aAiHnF3mXxWGAJY1ru3KvS3Qe0OvNdvT09UJVR4WQOCz6PzAUrzkKYVD01wj+i3V
dpRUA6iJkhmuMKrroIvF+kJAJV11MyZUw/iLgw0YH/NE0SuqBs7x2kr63wq6RFvb
q2MXi7P3Iq/NK3dbr/g/VxrmUJUU9LeIEMvnaLTpv3zmWBwBaywcrQGDOc/FPbtt
biPtXCLPXkhknkVVQ7BGOiDiGsVYKbw4P65ludVCIr2g34ZqZRhjP6tLltEvDPt9
qhhC08XrlCdkWda8MpDl+2HGAIn02knqZbmssMk+qR/YYggJlY6C16QxAuz9t3Gg
mapVoR6fUfEP9IHuET/ZoEU+yzh7kZTdMXsKpCxyo7j/rKCRWiXPNPKPz8KD3ndm
9Ec2zhtMiA2i6aAIMn26mrIlfRxkqRNY1ZQxtntCbBfA9wY9rwRJMfBujjUE3PQh
jfnRM01fPUmbv4qPHlsonbXg/5i+2BY4hlJkuRjAmtCAFVwRKb5R6mDYahDNZdsU
wUYWbzqpNrCmvB2mayP15MZeQLUnd4YiMoDUATZVHsvJMCVcXuF09K92ifk3pBzE
n4bdT6A1gcQLAwIZBj7ufPge25jmThZAIVTn84awDsid3luX2Rec/MkFcOGO8i8j
/czvt9OcRQgXELW1MLz9zhy03UgUYsFkmTlJ16vPI5ueMZOe0Bi6GUlqfW5HbX9k
ccWLVN8mKjOhbLDomzY/otWxaVS47jbtpvZ+8NvKinJCkKW9ZfY4EE/vgtgde3V5
cWAsxbQhsGGSlVPaSmUaRNavPovatzOIfFjE6v9D5Om+mlgFAc9/Nppp8SxJpGqT
QyRPNd1sSG34J3B93OaOggy5MpAY87Px/HgBgWtXcSgEpRAkJEcQl0kycwo+x9dm
OhGjOCt10KWu3QinNrPB3CvR7I6OU6O+b0JcilV2mWAGjsZAn3j9oygopEMNaSua
MVixQOWbxT4gndEWJj4e9jsKqRV6G0/0hmxeygLNEI9Upta0kwP15BHQz6Cb8Zl0
EtcH/Esm0UuIvoe5XJ4IfK5Bf/O7PUDCi0O22GpBMugFIh7ikkh9+PKBx7Pn5F+L
1EHXsN6LijSa25PnW7XYOix6P8AiYGtl2CLnHVgYHyYCJOxRi0SAHriCI8hgwNPq
LC6STqO2bPSygM8o2tY5brPiWJIlipngM9ggJLlR4+lMyFV2MGuYmzQN88QCN/zb
bWU5g9itGZsJaHQhWJKCyeoQkOINy9CMNzBuIR2YVMq92y8gy03u9V/oE3r7uuS6
L61BERNi54N0UcIjfpKthDfYyjkdt3bI5EJ1ZbmoimGymPMsTt214DxmfzU02X7z
meDwIfZeTN9B24fpEIHJj6tRg8MNg+08kJ8s4bdTvBCGxqCa9fiEZGTyADGXcKid
qmuR5mC4FcZhnTpZNYKE16jfzIb8VDSUdMSd+weAT8XQm2E2K0+hzj9mx4BxRDPR
bzNNaS1DyjOM/tyxJKPRnOlD6wf4zsj4PZcixIdW9z5ZhtsJfySLrj0hHX53g2n0
NzXyGfaIeM6B+GWIZiYBYVH2zyEgYabw9jt19iVBrp1sRCof0XIwKHIGAio4xODT
6e9jqD+EDktM/gK/0G2uUplbI+QQuu86+xGsEj9AjZwecSmf1/woa2Z36w0ECujZ
8fgm4vGfAPcc2QLMUANtHU/gL3BbTglAmclV90PWT2QdynGheWk3nAN+Q2ppkJQd
HIhY6v8A3P/NyNzncDwAa/nOMgt5l/XwVkoZkv50FQ4OauEdlL5tzJADeXXPWkJt
rgIu3n4cdLtVqeCcMSLLKP15fVv2pmLpiZk42iyUtWBUD8apHAAbqSiS16NUtaIJ
0EDnwFdAblQ1ZMxnHDrhfcBzG9c189+WFQmV/XB1Bu6I2LyJDGwaNJvch5eK1ouI
gSu2prFcswoXGBJvYArIKUFJDjpVcYTexqLqImKkR1MQ1atXjOkS3p9bIlX8MzeS
XAvMplhi3ljAwHLZrGriiICZthST567eOsGQS5SLe4m6QswxIBb39hv0xkDE+kZ8
ssu+I+/6tAgy5ZVPfTInA3zLxyee7HKYc+qWq+/LoFxGWSp1CwCc4gWK89DRyVeF
/a6DRbTPdECRIYuQ1L1+m0N+pmGIALuUAgqjVtsEwl9R6ka737Dy3rZkQlUrK0/c
mUKGabRB/HUA+SOh4w3G2G4f+u/nyIa3lJ7EEwz5j/Ej+sWyjOd697nZzaFboKTQ
oiqSGjok9k16FN3w7D5lLuRBPR/ijSk8I4K0l1l3VoJG9X+aLBCznK4ZknlBGURF
nQLL+q43uiVgMa0hI6caXBvUf/9yIaG7IjGRfbtuCTbp1LtEzfgmtFTX/BYsA0Ty
88oNuK1ypdMKbFRA2NpdtWID1uo/eIDE+Nn0Os1UC8JBFTKKouna8RfTPLk070Ov
nYbhyRPiPK0Y3iqkAmn+oEItPi9a+Z7TTi3dnuF6HcHowaYaRnj0wgDndnzRjdOy
y2lIVem38CHzPJeqecBbvWe2+ruVV3+Xihyotvpx2BzNT797ziXNQHADdvCHmMKE
A7xOAFb5eBIswUODJDKsbKhbRBbZM0ulmJ1AD8MDmi8azasI8RRrkT3o69kkBu9X
yMuCQAN2OWEF6BHbolQpDQ==
`pragma protect end_protected
