// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Gz538IIUGGBaalwcmdjTS0CDTvHAMmJfT57qFv+oVf/lSfCvA1CH0I7fJzik
YLNEC8Rht9S43xbdGI+gMyVdZ6UvCjchxJ0S7gpMUnszpquhmjdK5K/QFIk5
rKJrRJjWy+bmiqxETLgoN1Bg7BfVClM8va33r2sbpzDXGsFcUFb9ivLUL6R7
DR3TXrpv8sSrsam2WHu73gyu9BWKc3e4gNY2kwz4jR2VulZzckiYpxrtQFyE
7LjGkOz1FIqZHZk1TkkW4Xj3AVAwxrac6FKfAcluIN351YH1RLKD1goccNnv
/xdgTp92Wjdj+lRrZTE73Y4zTxR8ikUdEpr2X7HXwQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
okBebZyPZrmGEuKOKbeSlNq9hs2MavffIx9sOnnZNxdh3mK6/Vt56O3MJexv
yIXkbRwLUD9EDpcoDdPhwb3U38VUyRbEpbgYMlV1rdfKuXio60l0A/DKzSr2
rCsUSOWOiuZtyYf5YxqmmbrrYnhFc5bLjJqVbS3HQ1O/6gEnhivGELGtaPMY
vs5mwuGY3RT8iWFM+YovyH39Uz+EuyGxZL6cG4MLib2klVEtMf12/7TW2QBI
TA32GTr6YBFKRbCEJR16uje4U3SpAs2fvHvEkNsWkxZduBMgyIo40ok2KMJG
8jm4OWN5lZUCrm25VqUyNSjeahtHii+7FTWog8qDOA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
WEfkqhVX2w/mkQomNBSAKjbv1MxjaNhYK2Dkj9tOF6ZChcKaNaOQXDhjXdUN
0OZu6b4wyYoC65vrk6yBpwXdLUk8lr2rDxdyr8gKTvQeVvPrjeyCr8W5aY6N
BJF9iNo8pxykHTZR2SWMWSViWtx8KQEVG95ic/zdFEMVuRVDBLtmOFQ5oQhq
NERizIyK5mp5T9B/KE1svFrvFOf6otfbhOggGCZ8fjjd1vH1v0F3cyM0eh8u
H/UBUv3jXJ4h4NBkRD/gaY/rZRkLYAx5XH8PegwvS0s3x6LGZ53sG6j/519H
DLBF8/IzXzgsUfKGd/MULCsfWWyC6ymuKumKoh9Ubg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
jj4ViWVQIMaSgy5MRXOI2u+vKiWjKxjPmyM/CKSFDrRt7zgYi7V0nMjLI1Py
SGLuWKqcbzX1N1+QwEiQchfJgFT8BNod0Hv7le46QGmp3KLxrUBsYTpmp0Er
mi+hYqMpEJjfH6slYOCsy3n6E6srZ8RuvQn7wlI6uQvGy/3fLK4=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
MC135Adkl2VC1R4f+7lxS6AfdLsKWMt8+UXHlHF8wbODIpuEzGKrGKMQiJmM
GFStF2fpYHTc8WEimxU0B1zexkws2mBxsdg/fERr1p4wbgkGfYU+NGxIujoE
yNpFktW7D2qvpokOvwx60gJOLUSfry916/b2S9WaujqEa2enAZlxIlKNRk+C
nQHqxPbVOlNJoI4GxlCPW9kukEZW2cmaLk8jepRS3uPmbuYQKkqZpB1l479I
2KlvBPXMff306K88/RFJ4M0rnCkT030RAGaqAfZtq8CwY7ru88ig75V35LKF
AaIth6pC0vBbvFAZSYO3fgEOhjPE7NAq1ekKRuzkkmaJ3/JBBgO1QU/E9Rwk
XKtLfQbEdV/Ipoc5udJhNNG+Jv48tkNjq4pVp4Ik5KKPmBlD2PcJlQDaPyZI
SvuSZb9mtFK44cWKGmitt1xcn6NNHfEX94VzrKzcJdj6EWtZ70YeO6Xr94Cj
YJlbIyn9GYLWHgRlbbMToi5qifx6U83U


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
bBiigXnRiAHAulJvvfrBgMIpbhqIPe4wVJYbo2VJX42CFEbQ0pqFhAYKbeTz
rEULjP8vKRufPXyaaICFK1aXrpDQFDfVuVzI+Kf0z7JqrXo3LQrfZsmNSxr6
PqorPmf8as9nMbd2PYZvIfQz7L27MFJYC/+CVtyP6+FK15S6Jfg=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Y04Qqdrqj8ZOnAfppyq4A4QbpWiNU9qBmK79c5fCl7zkB9VN6Ww1p7B+AqmJ
6j5EB0gjzmyR5P55bT42WGshx5vZZodqBW3YDwDaxUZDmR6qE3Gf1sHGzIH2
VJoIqmNjVaetdFkl2etj/R8jrk+8hcbYh5uXuV5SHrpWHEmXnsw=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 9808)
`pragma protect data_block
r6/8pkVjWjOxSGDlhN0pxTEdKCpM5zaua+3drufwt7AMCZ5jZFQNynLK7Wyy
ChrB+KD4tQ6x4MaggKHONcqNXNLUvhnRKHhGP0+Yj+tYzaCGrbGzPn6D7MWt
638JxI7szj+G0fKRYoBM3GuT+1BAXYyobFHY+y3AZo03l9gOXRgNNL+RlsUq
UxeQ++baJCR0GRvbgqyoKJG6vIYC+Z/xHWBt8/m/rZPS78P0Of67OHItdjaX
hjtucdJ/KGeLpjiSSYJIFQKgc3T4WDVGuEg+2VXk0XizM33AdMPAAnd/ikrb
FUEdgVIuY2vriXdYQcJSXv001LEQ52zgHb3d5F+X7XT/HAABdsE1Qs5dWVpI
tYHyOPxCrLnruATploCWe4mMtO7zAzcezBnMQ1fQ6OBVF63Um/EH7YHfmG4q
kz97+0nomMdL3irAzP9JlLmHIuTIFxiLegADpauNu+bE5X5iPM8B322R23S7
OFnmDBMw7GI9QnI8fUt8EbxtuI3JNyjMrhbhdj/6iJVkGsDxbagmRluWO/uL
Fo5VoPkRQd24DckawODT4vs1f5F2GHcz/xaIKCiSWv/1/AE5fkp1bT87loov
1nowm77Y7zZEs0gU80JsitlKpWavO1SMO7pq9auSXCW8A9dMH2FvKsryjnEs
dWZ/THIH0z4Ij1AYD1yGlIHF0bfsML+xwk4fLuURTRvl0VDOT0G/52JLqKjQ
bf+Y5NcNKYDtDfUGvwddj/XO3Zo4TlURlmYebl7T+341Wyy5FPJG+Ht/HWY2
nHqDo/g1cSvJtoL5+Q0BjBJu68zAcrszyYjr3gK6nYfrbFfQ5oXD4IWVEC1T
3XSK6V4nLIZ7JFczD+/VNUipYRjVXoYgTBqF+qYbUwL6prTJH6xPZqOM1wZG
a/SqWIxmWziKXlFseMo4inaBj1DHHphE3RZxuO/KTdRFzbUdMp4FD4C/jgBK
7iU5p2FOaJzJFAOG/cdXis9eSQhtXakQoR3jSFtZaxNTj+LmDuPJDLpZbUca
DtxuKSfNYYka5+LONzOHHRTaDC+E5cjzVIJfFtbCxgRtW56PRzCScQEurrj/
bXF06nQ0/0SoK2VzhxWLKTVxC4MKDXZ0DwjZGTxALZiLe8UwtvfkBPqXPcZ/
vJklCU+2rjE9lFlWdI0RUC1nN39/dywSbMb1uEOufg6B7lE1hBE1GShrNmOc
lB21d65JcKaNbUeZYZAPET0BVIvHXqNTBeY/FtdzAWtQ1HpchNQSTyIZ/e1V
W0F+OvOoo51VpEVoVg/0AoElXF9NiIt5rbq1IVGqD5k1bDf4b7pQ2UDiyXo2
pl5/QZHdHPLkqJ38BQKbYTCetYn60MO5NkAYUnbSHAs25ibS07CiclJRiCB8
dL2Z1/IObvNTDBPDrJguJRU/YvrxYjv69EjnesyQxq0vztH1BNkPqvxGxBDW
ZlTr1tLhtJO9wUpX8vXbxX4YghXSkLuSDmYzVjVuVV9f5nm8U3w0xY2xNM4k
gPLSbdq5eyXXtf3o9yB1qACIgrKOMuo4i3nhgUYfbirKqvg93NuSH1KIsPFX
xz42l8PFHA72GyS96D4e28+C+skUTn3dV8zkrJF6Y6JtsfySadRjFvuXMh+O
FC8RC6nX9GqoX3xGIr64+1FsWSQv6dF6be6FfDPXu0sY5Obi6AePzEzFAYEW
Z1ykgxb6dATDmdUDGvb8HynbNPG6XlaKbqoT17Cn+MqTa4r46Ibl+TJU7Hty
TqjR2kjjl+opIS3cKb8qtW12HXhezLX71wapg4Q7g68ESXoDTu46dWjPGsNR
0wLXxKZ7aRMT7PNei4MI8G4zkbvMGi+HAayyI9tF7c5MBTq7Li0KSo6f3P3L
KZesZqDKT1ZIQRoId+uS9+iX7pgalLV6++AaREn/IBnmtQ3sx0ISdi/arZy3
Ajl9lbN4THH2YPv9CDZr5qqo/3QEu6huS9nXbnSTUYIq8RhRxyI5lNfkUyZo
GgouiL73v4TCv63OoyPtmh3wq0YhKlx1MrdOOSFyq8iroi9emVeEoiStxd0z
GmL2K/dO2gdC9vQKxuckAP/K2PVLurL99/ZA8NNJc54S9E5ys5O4URmF8nuD
P7sTg7j5mXbv8dQ93xPe/2CbMNe2e0zmZOcECOVXaXIwf/BQGiWXVmdBtAdd
dwhn7jYOjHreGusEdiKmR0rgI20RM2Fb3LnDDrA7b/2uZaPfYMr09cTvGAli
DU8BqkZDElCAG6vhggRG41hPUPTY91wUIDdZaSJUqTnFdnWsttkY/gpYv/4f
OkyFV1Zo0N+/FYTGFscqknwiovWWa5FqciC/7Li0iRN4ToDyM+/nMh3D02k9
Gth0QmUUQLosSflyHa9D7GTRUmB6SK/xOd4VHFuLQ1AXXRd4gTEtznR+KWEx
EmMjVMGHCdMR1LQjd6JPVltapjM3NZi0FabqmTo9MCADEoHGPyJx9Ktiug+l
TTKdD5yy3LrNN0Bc7HH7IT1EAItTgpDKbgRIkNeMY5Jk9MsOLSxZGmJI8Yp0
xqJ/PANRXWkseW0czRXveF9/COfJCPax2nqtazZQDTY989P7hESRRrSJOhpk
OlWhCSs1tCcK973BiHjG5pquxb+xvtdFjfqqLnKLMw2X5QCp+ZebaWXTfb+i
LP1UvGR7QR2HPnTjHY23LltFXH33BABwSBUNkOuqrHqhn6clZ3DKCHSXxuke
FTZfxcW6bNS3FiJqtGiQV0mvJLJIi0P7iic5knlodnI/ozSqrqOQOBvlg3hR
LR8thZj0sck1DxKP6jkW/EYwEhRUHIcPfMu8qsL7BiPKcs66N0jtJmaqEcU4
t0m8jB8Gs5jono4IGMMThl9qCyF+eexEaPgB9Rd6n9cE8Wh7dWbUUCLs1fM5
1tv7UCF95A7b1+Gxg6WFWGjO1WYyIH4yNlptAgRbN5CwVgf9p1wpc2tVp4y1
4F+86RnN8RbMHjzjwavyFtjq68+Jbaf/u7a/55KiPWFeIk/O9TLMsDFfEwnX
T4Ect+oGtnF+qkyD1hclCFNlsrPNX2IfxUqiYzfY+/Mbsb+zglutsJWsoT5x
eZyIQjn8whtELTsRV0905oPpCqnFOIo1140k9uHeoXRuuX8Hcbocy+holN8z
QGKuQzdxHJszXgbpnFoqDTsiCe4QtGnaIx07kJqu8LhfM9OL/AFkFoEsZO7i
76mMqlqAiv7GNqKP68fuCpmiIECWBl3MlPed+ySF21QedL7eEMBu+9Mj8fhG
pSHlmKjewYSjpc7nOVpYOnKwoEtQJypWETLc+DoDtNAr6OjK5vNEJFGaFk5X
UYqU+7j6PQq4it5jLDDqaKoJ3ExXZ0lmSBJbBbBR1gcMsHLddGJuT607prdB
Fs4izCnBI1qrahBIUTgYwlBVTE75JmEEljMkxTavE5nB9z0ObjLC3QjxIxsV
CgZ9sIcmXv7FbvABDhrQNZJKXq7CY+2nQPTallxrxvWp/d6JHCDWvPPUaeSH
lwylDYKh+kWAfP456SFxBlb6yQtyV+hCTk/91weqCPmwVFkUHlleyEGNCklG
FLbVCmRU9cLqUnCvREk0+mVsT0ILUpVgWqcDIefveLw4K5+Gnejk0rVJ412i
17oNwzDz3GcUbMbGbkoBI5wDYWdKF6LydBmCXtm17tHXIc0OLDBtxcy30zl4
fVg/l078O28IOganD/T/dtQghgywElIgR9JKWWRSXN0cVHWeWqy9frBFPaVi
NlwpciqRUNqlirU3a5R66/JMK0pDGPMBmysdZn2zpPzjluezGS6uVR61E5tB
+PTnaSv4r9rkf25MeJiwYrZvOeGNeYggC9FsMwoiNOzfa9eBWj6TXsPheMIc
uWk03HpZs5rX8vWRrt1WgGP0JFxqZAYYFOjFWpjRpe6XHhEBtQ3q7Ppa2pvf
dF9uY2VJwNODbb8cLyO30hZQE9iWD1IgLIsSvYg0zCtMSApUWUCa85qiyi7u
19b41aNs5S0di3RGvqKg536wloUyWdmUpyrADve7R8PHhlw4WHHqXz4/YMJK
QTr4wjBC9xPfUQEUxXCfg9PPcph2OksN311LIW4Gh0SlfgaOU20u+MR3JqCP
xbThoICnbz3Ht8OgOjGCqr26QfAbIrE8Z2w2t0Cu9FwEwTTvxliWsh+9tlTo
DqsLss0CbkvirX3dxHugahwx4qT6zqp89hMUhJDz9hiag4KqJXyOEi972ixf
Qm148ZvuUij4FwG4zOs56qp7nxlLKYWb7dfTph9yW0MFTL1Gmh9aM9wzVTQr
1okTU2YlYJOMxA3rfBk9pkckAFR0sseiuvXzMK63cvs46trNlcF3egAyX/WH
O0d8V50vryz+MDEZWlEVEnWXY0iW9dNpe8ndqtqqmSNEDlJFZCz8Sv7P1CDK
Lr8HjIh77gjoyXqwZzrSgtekJ8S5C8s+jVHaAbRHV8quKEyfDGt7/35esoYv
caSBq+NKGs+Y2Vlvf1nhmK1kuUIDB9x5y3hmWodJB7p4GoxaYXtuXXb+eMFR
SWzkwhvQCK4XfXfE4sLtdvzmcXbYc/5x3j1zT7p9+g90eZ78zeUGrDdju7UW
qV7jogQ8vC1pBrpXz4zf61XFRFRXaFPZ1zHGvvwm6D6/BhxcfVsSzOTti8Xg
gOHlHUV8VRXj6irh9DWJ/OaQCvtG2VM3+B228ConEc0hTQppSgvvx9g+FTAM
u6TaZ9hYCFF0tHP+xWauJYCPewbVfEYG5DNxHxRDtu7GoSU8KccDzWcBssCT
veGiFRSxHhM3hixyfRr9axINvQVX5GWD6GdQD8cW6i5GA9h83rZf3E+0tvzp
nnbDaq7G+TV65AuxqkN6wxo5ptboOUcGBH9UQyTJWSlXnlpVKlovQKd+RKvH
tieujjL4LXMEn6YzGht8fhla8XJTEV8lw9W7KoaVkzb+Boho9eKKbJAVLErV
xj14JYL5RYrKM8ldR08+iPIs0yIqXlIDWvq2TKnaKygf8Z5Igfdsv5O+Eswc
yMAH9TcOSIggVEtW/myqXhNeX0SYv2lyzseeCOaUH5KNv6fp50lJVf/Pyvh1
MlJtIZtJfl67yBzPIxgrDoCZZbcYmdUIUvI0w8nEgJxxkedsZrdsdoB/Zg/Z
/ex/97Bc5IhoV/icvEZIk+ZmHYxLHWpeksOkCoaOx1DEomqMyRhIQoY8pGWG
eH+XnOFFjpqbKtJ12uDwmAJ6h8xxacfHKO+BO5tzIuc5we0aDjmsknDVrZu5
jQ8RzER4aGuRYyRPvSQZHAugE4Or9G0m7c6XdCPP0TB4hZqhMe8esb33Pa7h
HpB7/IQeaYkg1rZnMZiVdF/iUdZqNqcddrEqtGnvOMi6aXMLtIo0WJpn9H/Q
2y0BflqjUhYFDJwHque82Wr31kDDFB1U5j32kQMFC8KRNPIL9JA6FuhiLyQo
pnkpPrKEkmwo10OipB29Hl8QLgAKyyAXIlFstC29bu/4a1fOLgYJ77HY4w9D
Gxp9EZpZqbf2w83lubJEuvo+quD2Bg0N7omvrB8tHgwG3nNJIny/HYa9HVbX
Vq6j7h7jzRYAQrHfMdg9fK72vzS7aRhiDlJtAI3gV/X/4/D1oo+wUXkImid7
mnWOqp1EeQXzYpU1ZBQZ7pMRPJeo1ULO53Tzvwy0GL/UjKOQ7KqeTVLrOBul
j9a16qlf/riU6+Jta0aHu+GTjGL9CRu+y16DmHRocWt25qHTMYLeZ3CrQwZq
GvXOshJ2KmED3kl6esEjikUx6yryB0DJeatdhNpmSJMgpfQVq00rRhrP8d5u
9GsUPQg+Ft2jhjJ8cITIa5wdtNOg0y6VUN/Gmy4od5rri5WO6O6/TmE4DtCJ
cZZk33zKKYdj2bTkJq1m3vOAObKeDoKMegtjkj68wizdXHJztXDFMevZ434l
FgD67K5psGssDCkfoZWC75aL92gCr5o8XnQkChrqZz2LAEFjmOaagxi/FXO4
+9yEpRUc/QbVrAN8g/5vT0P4fuCrYsSeDi6KeEj1uE23tsjAv5wc2o3LqtQA
f/HdATYlzECrj+WbTbK6PW/i/beBqNONNtbS0qTZmL5Cwj45nCANg4pN4bcD
TX9q3ZN+0CUjKMvyBVzpLPVgN4FCg5gMvitIyDgk+uEhw/x139JbF6Hhxczw
3jawamm1XhtBgRJ0579SOx9nliGZFP9UHQv122SagjlBK0vRhSQVK6gExcZm
d4g4Cf+xG2kqLCly1c6XqnDY3MLcvG9oXmlbqAmjHC2LHkChyZ55kI3boqWn
mK/cbjM4m02q7lRyFD1T10LyJsCwtlmQyDOETZSZ4q7DLso//QIqs44YWw3n
VDf4XeJdk9y+8wfRK484CypZEnyVocwUEwMDpLhQrAhkSQRn2ZX2yNPEsi8k
M3E5LUHBo3uGTxomM2DccRFq5Es1vTGrr/NrygYzSzbNV1bDpOFYbGIXD8ma
jcqEcQNgCp4kENuPM1Bf6GU2kQZlmm43EQkV0RF1o+pOgwT4kHoW9SgI2xEn
WRzJLpGl22+uztw33DkspJL7ANIj992ImfXETkWAAeqYVLHkJ/lUvJLFJlSE
83Ro5tQy496K0Qgo2LuFxRMncn2PaAlP/Gm2ifG+ONAGs6edLzpqHpgwr9Hz
VzxBSKIKUd+thtOFXBHlh3tNt2GrUl9cE+rpBIKXJqTTb9/v7O2KvCb6hP4L
BeJJ7BV68qX0es484Z0UGlrSfCOkI2xzniCPnR4DMlxVbVdmvsAmeb02KMCE
WLz7Zj5zegmS3b1tOj9BDkwzcs5tcEBv30BoZAn6CWu+hI0pfjKHLeLGgRPr
cDU6NM/Zqr9/1hUtRJL8JI2V3ar7ay5Q/bmTwObMynvhFBjEwqs9007tld4g
c5ScL1O5v6UPAwNQe8AlZb1dyZdZPoN8xA4MfSagMMjCWdPJKmfyojCGmXNp
W76Yr4RyoklNRLib1Jo74SOuEjDBRAMmM9Mqa4dG6goBiy03jAjcW/MNmbky
kgr3z2IFLLBAZ+F1xJSZyQwvCywDPeyqD4YRPPeaL0hcMck7gRBP0TQO0ldv
pz96rbY9ct3cbb5pIivk80OiyUjc/XqXXw+f6xPH9aFXK9h/yUI4oOE+u8cs
Cg4t4QeI6+aRu2AxmToGtlbHctML3lig4Hq9SCnNu9TfMsnu1FN1QWu/zcQn
aD1pvvTszPDSFwU0fABDychhzmC41U8+lIN8qBGz9gWPO7rk0m20L24/LFrU
1thX8hYqko+y14SDiyn/twKJvTPgAHs45ZHl6eQP/OiEhLUp12diIqpK6uyS
3KlRkSoQxGzmn6WN3Oa4I7A22JAv8mFOi0dp1JPSEqrnZn6hx/igQPD9Hzx3
IaOYc55082W788AQ2l+/J49ptw8xCrRP1U+OtjS2hBi+wp0OBZIFVh+8bMg1
10KulJNGOUNbzNqMHqnMXGi3BQCjgV2YlseC/0o3Sqp5E0GJZ7QWGVveCnhU
Mo0HP6jS848mFyKyT+eqKwUSCdjLT792xoueySpAc2zoriqcYyNU4C+T/cyb
bwEF9By2cvl+C5JKk/4dUUD/LGpI7254QkBmuC1V2hmerHm9MAFztt+027Eq
QuC4AMlr5Pn9LNt2fw/i6fHBSw5Wdg0aZf7xImUjJYfDVTvHj5jlIQLATkr2
wSgcf+9eGGK9CSJ6c3j52mxHqe5RzWlWByZlnFnh34YU0Mv1h+QvYiWxuEqu
QjJqKtBaRlNYrXWmHYUF+mxbKptla5lta65EOipsGCSYMc0urslJzp8cSHle
I+zAefmonyFIKjP79WpBNwM5TYbQZkuMikk98+Gdrxfmov04AIyfkolMB2H3
wIFjZ7p5XCCnQQwN6FPHp+mGS/zlw93fGgvA8+rIzxqKsnSgC1uFrKSelcys
v/OybYKX3PKziAnGiJBfpCeYMndR8RJ4AVr8mdXmCzlqaUY5wtEjeBbnNx4c
oovdpMJ7+cHjqd/DoLiqgxOk4mnPrQuowJvRHhPJeJYG0XwWiMah2e12Xd7z
sDohp+6YxLL+oW4r/XiRF2FOuCIre3WZUimZ4rvqUgYKYrM8/iJN0ZGwGrFZ
Kjahn3sbFIaC9yL6LgtCU6GQlzPxHfknp+Ya710JV0pp//LFSFMNaZNkvMiz
mhA+xdTavlPjA3o1aIFFYOZfbhjKVaUnWAA4XbH1bqkDawQOH5mUSPNAVex5
2omQNWk7BwdVJfEc1Pgosxu4wnWdjDP1GJwSSUtNrmr4HOz5Awh9QksuSB7G
v/hsX2wXxpOir+V40L/rBVfXx44WVkphCwtqwMVE62q81PW+XzpNoJHuzwo8
oPWJ6zR6J7GwW6dvrrlLzJq4HjmOet/9dOknOlCOXRdbmCsy7ewzx/u/kasp
M4S281Y0LYabwLoybLsOfpI/xI6tPYpot/cYLaBXKr0PjuBZtOoYpFkd5fpC
Z+OzkD7NZ74q3I3WyAOmz/ClMgNaIEbC62eIfhWdYVHdnOfxFHcgzYYcTwAI
OFE3qcOj1i6iaE1Z2NSBYGUFaJPRp5K2EFH/8VNnGCAZ/XxJUS0L1ylzzqFP
2lRPTYR0zNNGodv0uIfrOHYuBwU8hkqrvCYvPfrqQ6HXyIYRDs4vV5e45lct
1TiuJSc9/N/xGexoozSG48Yp0ueNhh/FSnUZdnwUbPqXmqXEWJg20B1UC5Pl
SkYIWgRg5Xld3nOeHJ/1a7ytwLd3lxSm/Q9lEIPMhyL4oLk4JYP//9KsxK1b
74/cyxKaIHL/lzdDPfKD5u1f8JQnsg0H4aZMIf/m6p1yyz9lDWW4z04sopgv
7ME9AWQumm7GSgn1MTsNJ4/iEw2zvf5f1XrZjVYaf/iesp8OW05b7ZOnc9MR
eOqBCFho+UL+awwLjMZwidOT9wGHfOr94qivQ1pStN4VIgDE4733od/gSeA/
D+Jrh2AJJK8KRoYcoT6Gvq07VhOAoXvfZ/0mIX+0+XOYx0nXrkcJQ0chMIv3
X2xURdcSdLA28eQvtUP56156pl0hnT8IbO1ikJAs9w3rubB1uW0yKYGFuwpy
YVh7PieKYG28euMYqugFz5qzHdOT8+H9FjozcGz9tLVC5FmHmTbdpYNo7eo7
0jr905lTop5edoYQ/ZWx6CZQ4PxFZIzcRA1EedyJInxaw2bzNVBb68WgA1EV
XDT5uHAkmlk14DlO0BhomjljdzqPMHz6megLm0gOkRpgbR2TBTuCHCnNVERz
eoyCosVUMaYKUzSa9F4StGHdX7LWBZsEKLqg/uWArulbH6ajQLHieh6NNmHS
/wEub4BBlSo2mOhbnN/cVVwHGpx/pryEqlXcCQ8kSjggx5zRP5b7xgAyWdVJ
YIg4vF5YzdrNSs7CiSICgSCKZ/c/5FyyviXa0S6GmV4OKkG4dZIyWsKsOK46
kIvbf/sVA0LaBP2p88zWWtBxqzQvNgTtfCsZa8TklPNHUB/O3afbiylwmKfM
u6hUoQODUjUkSy4vWYEo2fjxRM1Q2Tn5PFg1njX1BNveLBuBn1+2rqun05N4
S/tUlxgwtN7uDcdd7wnteC04KCnWaMWmJuiSZ+aAycqucVsa0Iw8w6CyTzI6
OOguCo0bKA/Xchs3Wudim6tyTASPWJPc0PhC5LKvLK43+EPklDGr0iISsI87
csET0s3J7nUi2+qBFFMtJdQhEtI+2Xo0JRNDPGUNSDae42i44s2aI4UhmnDb
qmwWZLGf99u9gXZdtVDJCCTGoOEQoa3ouHIc15k78BAWoDJUfXR7jySkTct0
DFOIOM+3vid7b8d4ysel0spHxw8ftKHcidCIe2XZU5ldBEgd/I6fdqy/HCOO
qxeN5BVoZ5NWid9wEmMYMxVW/X0riBbX5vdb/OLx1Uf4QLHtAQz9FWMfBVJ5
YATWypxWiHcRem7bMhkqG3At7x7+itSAvIpk8V8yq9bueanOxrXqnKHhYvBp
ZDPRuKqXPu1NvnUmHGWXFrgRKCy/exKvqzIiDg2Dgn5YJNTIJNohk+ofKZbf
W2PgZhN3IQ0ENMlOqE6lUzDIYLT4Z8Bq6TFqqtfMIbv0AcLY5DPhf0Ez3CjW
vh6m7Zk9nlpe53hW7kZiyelv9UKk9aeJFsRjE9r0Oy7jg1KbYuNH7cPWI9cg
qhbl+UkPBAekHWUkzagdvKkX6wVCsVdhDTevJa/7c8dGQzI323l8+W7fppsS
uS1N0U4hAwEPZaf8X7JzLNWNjSxPnS0M5PATOy41eRTU0gQlhZ9CxHPT92Fg
Q/9c4XkKi60GpQwoOh+ItcQONCfjR21ULpQXjEsFRcrX0Jpk5EMLqHmQz/YI
POyHyJEjiYRXtCuZ8jvVaiO68EDtHvOk3QEvDk9H1s4GHJRa8e2NErxKdiBM
FGOQdzxj6VCbDC5D8fjYyhVURVU/ZPrOGwQyJsHPuu/rmj2nPZSC2nn7/7z5
eJKbVF4naSdF+9TAnpo78v8AXI4dkglWUe80PJ4e+Lj6yGJ8aouY+nn0B0M2
O/Y4hom3vv8ns4++gIO1dA0c1W0aehIORQ+w7gH3PoqZMUWdkhVtccu8Loxb
TH1Ic73dzJBo7RchsNBAL3bdpU3X254Es14uOnAl1jVNnVNrV7Qr1+b+UKQ1
JrMu1qmXTWNj+HU0J9A/0UkMzpZAD5ex8k1FrovtAwMGscblSWWrw0tKi+fd
d+Zi+Y0NBCODUygqLUWVJYhS0vK7oMi3JTz+UmWTyMT3gfzqdQ1fR+FZvuWR
tZDTFu2qbepNr7c+KioSKkblpvhQpDUqRYtLZkxoJS5NXU+Gq8/ciyJkHwTW
VTuXOSwRWwlLpGHicUmY6m+Or4Tyaj79NmcclkNa2G0xQCn35uJ1ipx/wZay
+fJS5jOtdMvpBZ0xQEZHQlpCUls9aZvvkNj3z517YpiB0OXIblx0sstSXWCu
rPImpHUUn9WnFt+O36CmpXQnhYQEfysGG0ei5SyVPfqhH1ZLo9+wPSwgfisY
BBVQuA/OxGSeOWaLFEHPV1gNnRCrVle092yVHoRfoOE4fgy1NXAwvnxD/TPx
9WfcfmPECtG3lQVKp8keS67xtuW45PORMaPujIBHIA/V9XNooC5rmMSUo67Q
O8ffD1bD09wxSxJ5xlY9J2m/M40kKG2nMt6197hyYXBL9txobpA+yyUa2bxt
a2NWbSqCUW4PTSvbJtV5pC/MtyfM6P8BwzJGqt3IyDH8vrLLvVcwHHYMVfPl
PcNlJdG3y38dvgXT2M4t/FtzmRWP0jjl8EslYc8WPSRWhhbjYheSp5Zfkuaa
A67qW53Vwkz6OXltrFyzxDWi0ekYIxrUvM5iXFCRnzoFty9ynZ/luYRGy/zs
1Hex1z17sbJw6m9PV7Le+tRzK6EuinomOpRNbQ9o6q3EbOXlWz/8OuYeBqo/
d7ypYc+XIzgryIwJeX3+EKV0EgBr8pgqyC3qkw8W6mq/SP0kIfC/nZEGiX5f
3YGAL0lMyZh7e8n/IT9Oq1kQEU3llJeohbfSKrXwP7qI2Eq8MpaHvfr+ppC0
W925qFreywsCHEZG3pJWeg4gGvfXjwRpLTDdsIA8b4iZIMEH4R2O1I8E/UAx
8dTDJOMgBAvfu711e55aWHB14auc6sk28xqwxsyg4iRId9Prm5gPyYMMvxxL
1AcXTqixvX3OV8dxKduV2rP+JMTj7+hDLfqAXEKwpB5yrTnaGBXOk8jNd2iu
dclZ6LIuSR0ZllyWz+Fb7e482NTNUXeLyv1CRl8hlZzHv6rjo4kkEAJ12kDC
i+dvkwfrFleBM2AMzUGguerl1JFC1m6atwNl+Nq5fCF5JQWAAj0fkaMqfgLc
z7PifPTsUtwvlcE+CfNIY8I+hKURAbfIqe6rvquTQbs0QTqgEXm7cvtqxUdl
wEMsRe3OUe33LP0uMo/2sQ9GeCqnVWlWgMadgkc5zLZvlp2bV6FvgLVme3xF
f3wQk6YYri97DbCpBJro0sXNE4/9ElxONx4QJkC0u2IUzxVjjJrC4RWdpjOK
TqxwAlT86y1HnPZx3pSOz90/5tGjI4cmA3OZOMIwmDOYwIGXZjzmJoeuPu9t
3aCtp7M5hFLCvC4tqsKLPueBetixJyHYGlsXr8YTZ/bsmxRl7D0cTEmF+rM+
jnN0DvwZSOZFCZNJ3QsGfklWWYcG7U7j4pMocvxlE2r+7qUud4UdGrIu4PLO
lba1RPKB3pQVDAkEz/n6fvEBV3qhxqsOjxGlFhzObriYYCJlz2IGBbFf1U/r
dAGH9UQOUNxEnKcv3lU/B0fzV4YsP/0KAOrUUSTm9DnwaQLDjL3r7FRdHB1c
AMggrkOorKP7BJTCzq7Cb0GYlHuSlAUByZQJkwPFp0R+1XJMTq7qfQkfk0i3
1fvtFtvQM+6cDXvQVpQkT9pLJkl9M9qliQfPDUmjraFufB8K+ZrqWTZZTozg
3dUAJpJCCzZ5Ec+CDgO3jVnTPonnHkTFAkhtqBeFVIXycQMI2Ma5m4Z9BeBA
b5BTNLduF8FqzQxRquoTafxdygOJvgKjKCvwhwEbGSKyLG6//UCRxog2h8tf
CwfBkrDJgc6Eym7HMRBL6im+bQkYyCNFBNiR5XQN0ovbGt0eY8nHyv3AeZSa
OdfnPFIc7p05jyCQG5BzcehBTR8JtvCtjkxbixf6ByOTjvCO7qZi1IyPifEA
vPKKqDjeOBYdvcaSzNxUNYtC/jusndNejYU/1WoSkJCqXbgFc0QY0NfV6O6N
kIwwCXV4NEsw8vQY9fBfLKM5wSe6/KlqUprjDFw5LiEQSI/iVun4jf2BKw9t
+T4tAshauNVsLecfeivWC5WzsxroeureBp0HafhbBf2rcEH6dROWPelFEWAa
UkjQ7eFPPOVI+G0XLRMvytch7OU21OZ9luUEAI6313eWMhEmtBt0C6BeuSuI
nIQb0SoT2h/6I7XbwnHcf3/e5HW8f54KfXDRt8b2j22lhb/7AfGxN7itmUEX
rsu/IPPsm4OMNtG9Av1BbmVGDt5wloV2VNBnARyitG0XL6810vRC4OBk4bhL
rKeB8P15Pn/YMzXz9ZNZPLQlSisN1+d0+juJyTHCmcyFerUISZX4lX6h3No+
EYIn6+vopwgL76X/ik1LvyGZfONwbymmhfKV+YZSxcF/edxI9zrh4E6DkQ==

`pragma protect end_protected
