// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
WaTyS5/nJxQJV6ae0zdu8KKRe+szLhOahgaNiP0TWHCYkzJrZ0KP1EnZ1Go+ffSn
9aCyc6P1elK01Wh/K6WyXmuAlIU1mN9zTgrKv4Rs26tYShNGej3fxOqr9B7T+HTA
YO3GaIGcxpMeukVhpCghb/AQ8a8hDQxI/EOorH3A5gk=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 10848 )
`pragma protect data_block
N34JUMIsC68N+37BBd4WDtLDn5Q11JyEsQziPcc86Fiqro+s8Dlpi79FoRrX4lIa
knrBp3w7l6KDLQpyfoOlKPGJ4R3fw5DZV1tY/RClHB5LZHFNYGu0O8y5pC1vqpfA
NBarrFM3LmAJF9FZwoNKyl+QXKb+SQ0nQRLCkGtgUy05PWTHwjr10oONk4ApYRXq
Heetbw2Oiuuur6eOmP+8TFTT8TNmQT8lP1zpcDjA+Tgpq0v8ZkUAaJO/OrzdGhp6
s8vU6xlS7rK+GtCSvbB9Ir5EyUpKguWCRTlD9M9EM2IraSj5pKK3EKLqli6nsddz
kfviHg9j8xx3WYAyJhNKAj2L9DPOOKJFWGSJ/sMH8GXsVrcCeTR5BZH/tLhLoeJ6
ArMalLmiH5UjK6IuUOzQnF7I7vBZ1j8vkfYdggPIxBlJPB8K9SYvIAIeDJ2v0J6Z
1LL3onWwDkOckLnM5INtIrllNENePwbTRmlUrN8fnuHWr3SEumtv3NAHfL4UdcMG
i1OWRrJnbIQLf73mayRmo/w+699vqR5yvwTiZJnU5fJfFUz8RkGwd2ZVXJcw7fpi
CHI4/BUvxmfJB/FXiM4k29wcZJ4Ntd8ule4Gt/0hgZSkTonir9ypiLY3y4oHkXU+
4N5g3PeJI181I5ysnK43JjW2e+YfPnBhuginy2vZSHMSUhhBeMFWYJt8UmWq8fJI
+W4HLy3sGH8IGjC3kFv1L01Wndu/PMAoOAydAEEGK9W+ba8RDSiRvAfjHuDeS7Wm
yxANZ1x17Y/3d/KTzdkxDF2VShUEAuoJzLXVrXoHsVCa2j9sGZXDxvG00aTbR5rt
r7dIhh+wSZwYuY1XC+eT7a/pAKEGFJl+78yBhnxmY7fAf04oFkSO9IlPFX0DrHIV
ZAXJC05Mhuq/6wqSpQ9IHdaYTpG72XhF+mJyVIex1C4KjHkwphdM7A7S5+AhiJ0p
PJJpmGdTDF7UbhLSlvVRaDTROs6+2urKgzetmU0sEjX5JVzhXudWkQg0u0x6Nwz4
ELU7qQeerU3mUqYS1ODUtCdaoOLnua4wKF+nD5cZZiq3GEsIczHBlp+7cpkLI4eh
9Rl/RSSg/VV1dH5tWWnbJuJ3koFwvDt0ON1Ql28pN1tVwHf3mMrEaQilZcp7fY/0
0mRF02q3O4h4FIlWlb1641rLV7VyLWF/BdkEfAv21ux9/Cum0BfXCEieblTMqYI7
uP0P4Orene7wP3DE6YWekV9RT0t9wsg/tPyyaIcL8+ldFZyDBuUo2eijJkCKg1eg
f0SOx2RdkaSsJom/kDe2DhAPn0m8WVPQ10OOCVSUIW6PxsF+UCWeaZJJOTKTD1qc
oFyVVRDmLbwAZ+iHGuKQ3ev4gYZXF/m+p3/qPsbp6xCqrIfV972IRF54vbKCnzbd
E0Emu6deU7OL2L83N2QRGx+7quYByuWheVTRxsqDCeYnpu48ibljBPQT5PCkvtpF
1zUSDFqDUZvpzGvTwZ2nkvx/05bnh/nNT4VZmbdYV2s0m5Kswb7vcIN/SiBkmbKp
dQFUeWAk95v/nlHKn2DyoPham8G6IwYYnRfu6jeA0lv2KsfUJFvnX3OcvQSDf8Rn
46Zo2S7EDvwz9oTJLiocePsGAHRWHj65WsBWZ3HUPZzp4OFjeDUjQ9HHQbjozx7g
ngc21TmdD1LuLeUMOgy9VJjUAmymjC8y9j7C8E1+fFsESVpwUHPB1rYz21Cp2McU
PIt0TJEqnOQf+xRSWRuSvbHEWTKWt3cN+ldNm94JnCF/9Y4Fk1sEsag/E1qSta/D
KWV3GFYYxSP4X/W22yRdB5rx4DYOodF20ooeN2GeNFvCRnhl5zsiQLavURfQwdJ3
4exGvgMI8XiovXH5RipFL+jx0oE34M3a0VD+VDe1nobiapy/iqII2QAjd7hF42fx
8Z/RbdQ0mTAwn8mg9lLC89L6kV0O0avbq4syzGAzxL/OEA4epZn9NjbqVa8dpKtb
XnXDvZlpD9YBq5wucyz0xzvSI993fZCtTAp/7zEUAZ71emzYgu4ShWGsmG/Bb2gd
GeY6gVji6rNA811KW19zRcEhJ0AA/KrCqCffd30ZUDWScy7oW6Vd8CGIqoFWsQlR
P1VFV5FUnBXMVj03G1i2wn3qxsFUVzOgEh6m8TjTOo/M4hbfOe6Ul2EpRM5TJig6
3KfIh1lops+XJhR9iI6CZP3GXKowGd2VLsy7uLlTJY6M/xvQVp5s+yn64KXuHiZ9
UE6P4RYNthcuT5JiR+urPYVqlRNUBpfm3NTBJo4z3ZiKcIiReZD1gTdNYGSBKcb8
vJpO61AQqPYGJJZBaUhu9hQetvOzXd4dzbHQW8woQArMqa8QGDvnNxU7NqJyc2Lz
I3xx0ZAhUYwFFdILTyatEOoUzqhM7LTWtn7mIGJlSog9hSrXW+feuU9zYAV7sQ13
/of3wCnDstqSlboMpEBdOqheDp3/iXeJbB81Z8WkkFNx4QAijpsiHQc0lNgY0QOq
J/78X5xOhOnbizt2rDDMCCutJlpe6oRqJTFxX7jMSZYpw9H3odDO53nUmv1ZYgsa
G+xuxs+4Whk0Fh4mJtL5xi6Fo1X4zqsn+v3jh9Y5ZOrOMSI0nVZjTkOEHdQJ2/Ue
95eQrew+009pcfsqPmFNGvtndOf8pUQH3PGUJ9+Ziy3pnoqrD7oAGF6qYrHjK0T7
Nix259q5E6TOeS0+f0UgU2GifQr5TVWejFc053g2S+4G+f7TNXU5kqM29kBnrYeB
NUVL2HybLox1MHpCFQUN81+uzymPgrzlr3JW2rvI+hMqPi3syXLb/Hrj9suIK0qz
Ecva5zioQtvRwPpQh+ZxSu0e+CRfvHDXw61kU1yxT+w1XblDc+3gxDs64QTAPb3i
9o3+NYEdHvXU+4t2pcH6YuY4GPU3VhLMXiZOnOveAW7qDncsSWTCB23ywavoaClz
JTLFa881WEK/Ga+yIn4zhDSgx6ecTX42GHNRax8dNWC6HCiO9u+mEykAMquSbrSq
R5JmBtiRE8eMz3eI7hpYU8jIqtK+kskYOAXXxjnLwdCurspWo2/CEvvS685pcu5H
eI9b1uWQnZzn7My7V82uM1U73Uc847mqJmGUB2rRuSwxFgLtBkVoKEXSUVeqK+Ah
v56lNeOtg2LkkA8uX4JoV1mtqm8PXum+ZX9iCA/O5AWZYPrVWV7hlZ7yA7CLdf+q
wcW7vIsspq/rJYwhp0rnugiuVo4DdH9SLIeU9Dt4lzkkqp0+RUqmdIUhM+65cX/c
UwS7uE7PbEW/1IoON2xIEnKNSE5HiHv91I3ljLgopBxwoxCiiEwrQY39N2cMfvv9
10iBdVJzOXZFBQ+RnrLRxe0qPVdupvyZpFK2efCzVoT//qpeo8dfO60bYVu+pBvR
XSwQAalmM2zmqgHZiNkvjDpiJYkgpXJEOetVkpNZF133iTAuVTG9z3dGPpc1n4mm
Bcj3c4QEJZDmwdngk8wM0tQVqQNnZfEKDGD5wnPYfNFv/cGfdTuXN8sCKczsFE6k
9Lr9Cg7sHb6jNVIFDgvBHv4jwWV3K/gSHqSBLi9L5Am+gVQsN9X6iotT1SzGJCE4
0ET99SrKMA59Feb98iYdCKzHM1cVqenKfZfuNrlml+uyVBwhvaHY9p1hMJaDdQWJ
1jdVaUoMvKdKpdKtoaRHj4JsBZ7Al0DUxv1eplsiSAcd2udGSa7WLCQx500u2qp2
FkdYiPDIYwboF0Dul9L6DnlpWnY3eqtTmigS0jJMX6VukTkkGZKDrxEy2q579nET
58WBsH3zXHHypgNtdcZZ9FQwN4elNm+imKqimpGbwUJhH6k/949qq2NHFPQP7SKN
j6NlLLO8wEPLGmzXPZz9EML3pUjIFahzji0mK1qZqKsfj+gO6wnSTgvOpl9+FamI
iJ7eKqMPlmnuA3VnlEn/835v0TWtqj6PAdBnInDC3T6AIU6WBuNlbl8csA8Li6Q3
3bF5vLM4+kgXR3rS8LLlcva/Kp5Ubfmyv2gX7alPO91Fi/Hb+kYWV12PBX3OzRl2
o6q7+ULsvfslE4uf2EaMWQiefYRj1TpczE+j+GCs7gt2Tm6o+w4Lpdft1zF7lnrT
cNCgTI1ZWll+OD1IS0P0ox6V8NjQQDcsBz9MmgJpdX9laTorZmCw8LF6viL+xQc3
NXHeVvokfbwlZer6x7QCUHw0ImTLtZ6xo++DJHj5LMyqAO2rd84ejolGa/6wTZNg
hGYV4nJuX8A/jfpJUmO5m+yVVgk1HSmaoyxMEDUuxqs5ArLFjU/Weo2jI9ipmjTZ
H9GyTJSCNfB9b1fQ164NCAuV+xaxjXrQruNglO5gHQFdlla5MKyf2OEP7/AriQZz
sv4jEnZ8VODNxzowPTQqNz1qn+I3EHabg30iB2ods6WKlb3O4uySX3fCKtVDZeZz
8RBS0SNraTnBMj7alPxrcH4F7CYqy0TgeQ9Abt/oTZKW8I0i0Va7umU+gDRJWwS+
SZQe5BXDco151g4MFblSO02Slzor28oeG2QhqQOgKArFNnha6uV7aIKmXo50jb1Y
I8fcWDrHjqfhsS7blRtehLgX9cY/w0uke7cT0fzoYLMSMFqkHVeoKpsw7EE8Jx2A
tGp6BOSitGb5/sojLDYg+oHM3gXUlxOxuQ8R9JwU9f1FjYD34yZwQHDc7+qMQKnQ
zUno8u2a9MInfId0S3lYw1rtqTlIxylBZSaSsrgiR3LkgPdlO0fmYyhv2VYwNJLR
v1OFbaaMs1hJxpeLkFdNWkagNAHeb0a7g518J89isfw9EA7LzcC5QtX+WRFMGOvd
Cy63e0VmaDgbWNaiI8qbodJzrz5jXOHb+PLWYa/HWNhg4Oqkl6Hu2T+x7MvNnGct
O813AUHEick9v+vwmbq2JQyFQ9zPX3MJlO4u81uhqpatCxClBvDU8LLGnT3kte4T
7rT7D+/q+rC99PM8dL5zYrh8q+1fhLw0wOCyY2il7dTUEENTzhul/6i+8MabO6gW
gX/J4AbrIuRMvYkW/XT7ISKFjtc7AhYNthQvOSmCXP9Pdp56kdEAOtw/BSmp8g7V
SJy86XUojSae+dR26Bxc7uhDPBn/WNg+Jt6Jij192pRF+gRcZbhZGMS2ehLYfbSp
K7BeXW7HRWrR4PJ+x1j/9ZXhjYIno28H+IUBgxxREtNjNEiD7Kq9RZFnDtWFJHXG
8GxbnmpuINbvdbIkAPRMv2FyAj8J+wFjQdPSlvdO3Angihd7Th+NQeqPg+f6emoK
FM2JX7+tveJQxwDBhAqnZOp3klofLsZrZ3TVwniuApB5IxbsZP2Hacs2AS71Fulr
ws0qIBIL4PCzowAbwigjHZB+6jSp+nZJT7DOmZ48Lqmx6e2iOozuTd9Gvce2E79B
Q9aJRJtQBkzkA8JeBnZINM8aVaFmPyY/o17iw7jid4fBJkb55rMukm94XJfzSKEH
H88eyhilROEUPmuyhCvexe6WzvUx0TH5HcfAnDt5ltO9sT0GL28dbTSDfcpWcysg
6OD2GjTj1wm2KA/AWmkloFDq65AmtnR35l6imMoPjcXlZ/cngETNFM2EhqKxrCt3
ceBc90mldUpVPi5P2z4oM5twwdkwE6mak9AEYkOzTIjx/tOQaNpB2jL7gS8ECVLq
ykowjAgvD+GoNOe4++QVY7HC3/O6q832sXPyiefxu7QoCOuQKAQt9iLze303UFyT
CjUWSw6Ii1hdBgohClaJe62tyyNWoajGT7o8PVsN1TKy2UcEWUvocIoit9DpS5vT
oziqeQ0cOpvR0Gb+dX5YIupgiCODnXF5qMHLpD5MMAEqtZ7dhl4hyin5Mcfb7mVU
fQxZhRn8eKDCFRR0+TmdV+m6LUM24znLVGzrAnDtMkhCxFUndhmw9IQX6yP1d80d
qdhCBkoXBXwU/ZBHkTVp6Vu85TeUtBK/0UqFl5frugKKgFwWNYmjtpWgOpt2ZWBv
85yN1ett3SuU5ZWVgqneHqPgeU76OiD3freq+ZdCijM/V/ItW60SkKnwXpPur5FQ
fP3juXZBDqPYcA0GAx/c3k2sciTzWDO4HU2G2qzJFEHVqGhktx/b9P20PY3944ob
w2etb3ykrRsnBMIEXcxynQ1l4slrxfOLNQhvTVg9OI7I0ec81TSnWrtbGuTqbKPB
yisDkjSpH4KEF74fLP2AaMTuJ0hFS9qLrV6AtHM5oo6QsCtYW9kWFgw0sKRExSI+
Bp9IRtBAxh8uoWejqpKcDD2I4TzkFrzTc1ojWBbYstT/SgHdW+F3Fkyr2rPi528r
xdlXsC/Dw6iPCd2azOuoy/QbGJXYMbnt6GJ7z+Bygri9+zSQRSqmYN4YjZTflxNh
knC5DI1iE4Dk/ZdWhTWtj3ZPv9BkHJbstQIWqTUQARxiTvQW05XNrfFroIIa2yGQ
MlE+wtUl1ldxyIQFeuwtdDqE4Nm9n2qQ5FthfnhincUOQjTu4ZeZi5F0uXo/s6ny
SSEbod3qSsAOpeeD/jGMe3Cf7HGBypOy+mxfgeh+a0fo4/T/zlrqLG2OTHj02U6C
Crvyfyp6xWpKVuBf8x04CmWVxKmn/XR3N3ACnuNdll2YrjjeTC4xdAbBG/yvTCRz
lwV2T+rxSj0b6JDh+21IafxG4X/njMGLb/kEb9pnj/vClWFwMhyzOXGkjotZh/dv
y5Fp2gg8yudKyj9XW/11lB2ubp8Q/s+ck1QEOwMOTpwU8WrVlpQAh6xNZXPXEsEM
VO/lFVGtOYrSds334hI1BSP0ppdIQP5qzfoOLQaMIZ8OGPv/9I0aC0ERs6OoJmSW
rDVpEBh8AeCAXqMkdL0MSpk34/dYMw9XMe3jBu/dC0m8gdSqIxqQWRQ/5jWCrWwm
YvsTUW9xqR8NWHKIUoCrw6EcRUO2gyW76cEAxekI2S5LkdxdH7aphR4mI3VgMX1e
mfiXxgrBoFbkcq8b52aU1FoZvi6rPa8SYKNsZJfQLcMnEjK0fapeLqpZY0RLfMTS
L51IS7PADacS0Dw/0frrqUHo4x9Zk8YkQ8fCbcoTHRmK5qodKHzGRswYGigYOgKo
LSQvp9uDrtNXAykes9oQJnxEn8OnpIqW5ZSCOnHUSHY2nFFKkF2kxxl1BfhANzUa
Zuil3wtALtAd+J511EFi/2olTygz5NQuDT1SOSnSWh4mh/UDcHp1XgTuKDwOul0V
cutB+oLuiSF598UiL/w1KLpXhJGDAxqasXNd5tmBNGfOT9DRbq9gkrYQEs8ql9vJ
F62Bjx9JLlwxzArVGAwXiowLjFYfVbnpsv2n+V3JLxDQsLK9usv5e5jd4hnFcdOa
NEitc21lu2yHtefSJNInC4hCo+Jrxd6tTy47SUHxV0pwL6izSR2TtM8rQrdy+nky
QtYEHZbNsv8aGu8L+v82ob5wSLhGwK6BkTernWIDwodV/Mb4w/iE/U0RUYYWAfNx
nWxPNe1pckI87oStlM/F8b3ue2FOpPfVh7z81zgqRVVB/6rgeSWVEUKcxou5hdeq
plIgp2HvD1erx5AYLZao9c2ykusRUyJf5mZrXdxAG8NSNEK6SZS08YmMYypPDr8l
rvVixTU4vmomU0Rl3hD8dfqCE1LgKoaEqYRH5nW4GtXObWOQPIPB01esmb46kUXh
7TftzVqkHabNmA+oPbqp6JE6oSQeXpMo1q23v5LDUC62th/9rmDVs2ygmfgZTbtK
sij1ia7rRciM6eOdS/30g7Le/xK0Bpdmmydhw2GpXGLo/epWfnjFtnyiQ4sZ+zox
x5NrEJZ2flgCZzxtRfblGx498hXI5assOUREoyKYusfjUNQwLJOU+gHkifPUGDKz
MTc1bSprQIeD+RT67EWu/B4NIBM7jzMBCxP7u/42GocgXa3zp7NmALcARJCiOmFO
gOxsmQxc2DCnvrEUkQ0FCxJuRc66ZVyf5UaRdLc65rVjU3tSH7sMYmvVpiql1pgD
O2LiYTQ4JerkrekjHBTah0Qh++PkD6RPe8m0AKKPCSWeLY/lPEc+zA13EzDgTTSB
VggZS3WrhpGmJRv0eB934HCUSHyg2VtZy51OwWfMxZBI/owCEgua7LrPV9fNhlmC
7AGc1AG/C7CdFNgbv2evedHBh1o339PzhmEGflxwd9IvU/K0gJGsu6vCa/eogIZu
G0Ihsju/QSwubw5DMpT6gzDqi4N/OASjVNrFxyrbBRgkfXqNrBtZLzlRUwiwDcVy
KBTY3w1JOy/tpWEd0GqpNAbl8edlrG+CcFyvjtIVF8318Q3CXjI61jijs8MsnvQB
AoPhva7zLL2rgO3f5GgFCslTBtCgoci/rfaijHIRWuLdVY4NEn90N3vPpqRUh6s4
4NUEoS18EJo/1UKcLnfBF7Lmyjab0uzwyt0gRdPcBECnpM4d021pArZpmU1lZSVo
EeA2MnXfvkfkQlpo/lIUQFmxq2X+hVPXVtavOrAs7HvKlLtW1yYgsJ4audTkayDP
U4ASx2jZjUGGbG7RzX9BshlgJymO5Tl8DiibaioCp+261HBA+kselsrv8FQtMuhm
q0fiz3RNssVqTPVd6t98zvlTZJ/0Qr/rXj6WS/wcyU+yyuH3INxLIByl1AsRumOa
R7k27lx5odQqWOLlHHdZIeqLrPLR2RmYz4eibLxZTBNB2UM0MJNEaiZ6U27ulRyf
0AhHBaBusLdb9JSD2h0WQzIDmbx0KF3ByZ/nzwQ/1CRYIdh2MX7BtrhyBOTq17Th
aUx3uEYk7rv1GxGl/SrEfGF9VaGoSzw6MAzJwl3KWS1i54sai++DhohM9KccpL/h
QfAGCOdSw7k5BXWIYtYbHD0QWqXuy5JYlNx6Feys32bfGwfySgKfcoY5fwDFtOE7
VVWqcJuSQhmdkDgVStF9+P0RP0ipfjD03Onlv1Kaq7l9F0Am4ZNI08vsRaMfpaIK
QrgHbwnTtvMdnrXb/D5ArfxlPiAQatYRtDq3DkITrKLv77FEbXcuioABIxxVTrlz
Wshqa4MfB61UKZ9r1MOAHC4Z/tcIQaCDV0Bp8fPuNOxSKzqMelIpTxiLYv1X84Sb
0yyH1pkjJjlelFN1Djt/GA7BDQcBztQrX8+dY+EKkhqrwC7KB9aBOxX1GHSUF+h7
Lix9zsC8bqL3RbUOMA3vyuE7GvjEXgIQSYIPq5jSKGy+T67amxPCfOnOCXcUXm3p
hsixkpIT2beBm4wmEEgh84NzayNvJv0FP8U2APxrOrpsxci6SJrPrmluPOb42i+q
kwvh9xLmi9GRlc9rSjx0r+gF8bP5yZv0wBwhCf6FEadEerege6UXSmCeluq/OyOG
TOGrihhTF1UAo7StrXGVhD+C0OjWrL/V5EeVWpFrC9cpL6gIomN0j//u13GOhzdy
hftrJv4RnM7V9VRx3d8GoD6fP1wsVqo3IXb2XDhFTSVXW0VK+5jyGILtZQI1Cj3D
Kl1zOXe4w2B4LRPjkt6G+Guv6iZSc+n/HCFiRD1P+TLPgRsWT+rbJ8ooKxOG9Yb1
IVebzFPN+VZJnoOYaCYe641w5re8vI6Z2gjDBMs/7ynjEnCZ3CjTW3FbBb+shuD6
gZOBFyP6QWUATna6+yFKvBA7JciUKuP9bQ1BrIefs4WLX0jI6REKXcAbpjlSqwgc
msekdA9LYNrw7uJwES0reqMrQjrjwXPP/LhjvGz4X7K4Rvri2Uq3JcX1SwmJGnSa
OyfEK/aoGjH2Afx6V7SY4IVCJaN4lFFAL24PVe1h1r8o56LL/71iyKB6FaeJnkEO
xqYK4amowcGH0qPc+iOfAIQb8bedaUnCnfsvgHbOR66shwM1UUoKDVHT0H7VMw5P
2/fnSoEq3FVXmlv7BlINBAihS24DXNLZDpv5F4ad+McQVd0fShd92yMi0IpBCGoS
5V4uReA3F4OIBclLF4rzpb6q22xiUOHzKUvqKDQnP7QJ24+kTKYuaK2dfpKNHM+L
BsI2wJOzkJlq8IHF7yTxdyoRC242Ow5K6hKIXTIVrK8G0FSv9iHenfXWzrvnPJXs
WLMomxhuB/oIsACDACwQI0R7nMrLedk2aByyPpk7Cu7xJKVEhe+SXIdH+3EDLDY5
hjPO9rE7ua6qe8uIiUyMJl2qXwURnwKQ6NTUNWQfgTAdBdJ9ct7AJntiqU8VPT5t
c6IiDNuecw1SfTSzwfDPT4bLf7m4Ao9iojP5NpCachLbOSDbswDAXxjItwjWDriL
rfBu3YMUWTaHLv5tg41A9rPu4ovAI1DuhgzfuKkY/qrybPsuTQAEyrOzWiqIhnso
LN7B+ThNavEYyWV/6hGjfC9EKvSBvZKBedkG1lIvU9y/yzBWlpz51/IsQ7IWgD9M
QwPxK9d50XPbw4vmarVebm4uBlmcOJ7BNjO3pAQp1lyjp/Shjrj9rqGi5i549bmx
ilKlDKuSpp2giURAgIN5yXDpgdIPuPrbAGzeExUZkLtf3QUqRMHzx4JCqb2AJ22l
nHmTITobIkraMhUH+LkKY756tZhitXHdBZMtMCXSlMj60VgIxxH5j2EYIL2zBCfy
eqxzqv0MHYWgox6OmnEekjkvfqY5g0neySpr4ga4Kw2TIGULSEkWh5XEyhht04Ir
HqQbSMpJMJluRJUYlYYD9utkqCrcIXSpzLsmVLnx1fAjc7P/y+El+QnKZQhxlnAO
ldsmcTp8iYOK/aUZYXXrCm32/OZ8uS8gdBOP0ZVtBUBGHd/ZUr2zxmakV1D4CMJx
pnTNyQV52UsEyXWBrTwdrUf2hbJfdOrsF4rJQyq6JKufzl4FS8AdyXz1mr0M8Xb+
CHMs1gupgvfCFpKwu12O4dIO0NLoFGCItP0fMMkGhkS5zlXdxhFCILnRW6+yGjRN
Qk4OkS+Fw4ymjkTkyG3GBD2oy3H4AUhLMumwErRu0N/7oG+ZwtN2Gc2IyuzLhVI5
0zYt+GD1d7w00kjDF20yhggYa2k/BPbRVH+1o/ppKqnPmebF7Z1gQM5XosAV9m8Z
bROETgQd3ud0YB07s1k5flB/4v3GnWBnYnsAKuPrxrRU1mOsoXmBZndufNUmi3Tq
rSDkLIYVMuZuVJd4rbOU5bg/UynK/oiXO3QYcOLx+csgE8M3l+nWKS01cfSbpLsI
e2+L3gNhK5HSYqy8m3JwcajiCg8wm3H20ePLzMeVJZbw440+9f9eL1rWeEnGlapa
JO5Ko2NIfCjM6v37P3gHqgFolFoPBqpqnPBL/7hlvTyIiyJGB8u4CYajybbUuSoJ
hnadZNoc66Ds2F0BPZeOegAX22fu/RLVjVjN7Paxro4SJlJmujsw+H1EBsAZx9No
iCn/NMPGSAeUhtmALJMEIWXPrHaodtMfEQBqUK33SFLCUikY9ldD6rWPLMFv8fDA
PQbs/RQRfDoeZ1cDjei3ZR8WOkEYfQBqS5ZYkzsdkO1eyc1Zu+40SSxJCOQiq/5W
dlPBCZh5A20Quu8ziSfjK8WadDtlC9N5Cq5kuKN4EW4TMv85umzmHFvniQzfyb0/
/FwuGjFv1adk4+GTqYrT1uWuugnvs+2nQ0iM70RC7wS/wJBM9E0TpDXjiyZTluRm
qXgpLnBATzwWYGm6aujLA7mlNjLcLZlD4VsJfpYjAAOgenu2Yez49CAX+5WXZEuE
zBjI0+4cNVJ3yHMpQBkLmXvR4rIBo5+MDJ1gjfT5YjQanMHdsKb04PYocJTUcNbg
iPPW4oF24HXpGVsP+mKY3ec6N1D+woduwo0F8rP+arMszK3Ozje94YnK2yotEsI+
d+8qIxk1DdE446I18CWMnrj5RcKq1tTc87kMRwA3DJy5F1nNgHiWwZShU7A+/bol
pWWxl/VC38FCBD2cEAdYMd7+9Q5k3JvE7TcmXE5BmnTyQ89M06HrWwT/r1Q9SK8+
QESt3umta0v0iEvHkzLElVdgi3kKcnEA0TK3gvs3UAFS7gAt03C64Ezt/WY9B+54
ztuRSPR6k9F6kgllgun9qHNWHkXzAfIzELjGgzSXMZwdT6SionEjTxdcA0K1V1bi
A9s27cKJzIONIMoYDYwfthf4GJslx5WUFeI7+GvlJ61I9uxLaXuQJSeoKLZaaRP2
ZwR9P9EV2BKjZ66jZQGy29jRXhOA4LjrL1yr4nEfGVSKA7m9TzAm4CeDaQk0woci
0f+OvJ+WnY+JhJdsgU9qND2BuyXuuVyo9/989z40hvxWCv1Sp4Ce8KsATFOUcgCm
NiAyJRMONhxF++G8t+a5uv0KvTmCl0OA52O1FVWO3hfoucVIXNbeRDSW1mbhEdiC
bwwIiVEHEbemX1HlMr/kVXExbPSqcK9AOe2hBGKeaX3Czq7l4Al4sk1xZjF8CsfC
H8qRYj8PHP3WCE6TjvvisWaHpku3uVDeRzYkeL9ao01p3DKu1QJaStCZxgDcQ5MM
Ydsa+yh/EX9ziBQFpncf9wS7xyluU3k5VZlx7oxg0Qis3SlGjbRwfeLalF3e+4YM
RgARMPyaJYsazVGqg1xkoYrnCX9Gjssug1tL0REH4xOH9/bnEb6eBe6DJNMUzE8Q
UJlxpdkHy2SF5sKn0aFzwTJSCdtFMcEVzHhz+GfbxekfwGd2ZnbJ313Gbp8iTL2l
h93BcRnGYvQMLIWusxDRoULTCPzpxOXiwPUExJfixqU43P5hy8Yt22uKjYe6Lf98
JdJA6SIY4NqVQoBJ4zcWPtq9BPfCp8H1hUexkd9PVR+Uj9d4hVFVO4F4lwUZ/K9s
hA810AcX/z2/L2P8MVpfmD8ueO+uZ37rH/+J9ruYt+YMMUTxy+OsIAw8aJZH3ock
vCH9OlSMJDlUNZLChtsUzvWS8HucTv1aAoAV30bQIVSZ3qNkFDsribI+sH1JBu5+
Vou9iQ0vYMGKAl9CxdgcIPPdNQGiFj5aQIkTPdLbHMn+65O4vkiMI0RvxC5hDEsC
OIFcOOPwtxlLSN+OmNykwMfzHB3YZrFdHxbA1+fW7jjRzhZ/LVcTiSqdzFDRZzoq
g3iHOCArj9JQs0FEMmjH9u4Z7L/wyUmESh6DG0JEQljgXfCFIQNTWas8WK5+KD92
7y13uKKry6WRG31BXoPzapC1PhsjnKP9wxmVdZHo0BqAdSEiaERN5PN398Ylq3e7
ULlf/rreBtcNJX11ar/YJebxl3Dyptn/uCJbwEvKmrG5cJ798CysFJunGooYd/e5
LKrsOgqbqoR7kosgST6Nyi6QuJX2Pp681QiDHQzEg2Rr1YDoXhKfdLjeG6HShFgd
psJG5GdlAbnoVjCklC+yclxT8QZRn/jidlJj/N7jJmTJhJS9agnhw0/ZwUXfHlcf
jnXmhztjsKuQUXEUWXu3uWOQLteI36QreHl5qS5sCzwRay5PR/6wfU/pzeiyVlAe
VIfF4vmIzOW8MjwPcvWH7yMkroR0V3wPpWEShty7PDM35bItqGgOhajFLihZbhcl
DWYitMGgq6qpb7in8EuBwKlWunDlKKtF1V/1+5L88CUuCeL0naFPuu13yur2iKFa
WlIV508S7Acg7hAdEbXJxmxCYx+IqQvZ1u5v8bayhrjJlWlAFstm7MzPUW4M4OaY
L6OQYFudvERn4y2OIeW6mndlM6BmLR4EKQ8EW7jlO3khBE8e8e0zKG4ApFR7zTCr
FL4xuQ8mgiUFE7UfyAb9kxQiISfniE0dLieKx5lk1kdTtgg3HcbR7uHcyjCEvh1x
Hcl5IrspgdT5sLdXdGAkYpu3CRjBtegYVGJdgXpke8PuFhkbbRq55Hg9Gz4mUf2b
6x+5MLivv1sMNfP73A0El5eahScm5GIgZ4B+43fu8yqW1oCngVkeD2vsMIaNQ4vt
3MPPK1h2bfMsmRGeftnd8cEVZaGkZTUzDxuolJI27WRG5q3mjoKPv4Lgeh/jDQme
8ppVl3M7zCDTSONYYE/JRCjHimtrGYUTTzoGDAz7DkifX6n8jVd2wCHgHnuuw9tO
dozd3iyYpsrQSUHWcgyMz9K8Tap69dwA78GkSCDnxVBx4PKiI/2jANCLH6fZqoVz
6kitXPC9M7S7588RrfSi0rs5yRJ72bWJ9zcsn34jUvkXji+Li/ZEQoSVYxRYwrBu
eVJmZuvju32wsF9lSrXELQl+MyZCOuGam6Web0FI+OwG8eM7aP20vt/pObMbJQo1
lezRGr0CNk3nIrT+9uuSu1NJGHDvJQaCv0U873/JuY6j0I4XQHHZOFfTsB+oHeOD
Yg+1Gbz42brKGD5tfqGDcO/Bbdd61VdpkK7NBMHafq9dcEkLffqir0z1wqkH/wIg
YMWNKf+Q2/yTOJ7XED69Jh+H1j3ax2WsKSDa/KRIzK4HWi1cMddM6CAWmXQjY7za
dirgDuxvonPzfgkgAaj25fVQK6cdk0+Zs6rL3MP4qcZI6eA6KrmZzpvYNd3U/7sH
IOxW9JhIWuVD+lat42L8Y7hik33SGxY9PGbNloA5hOqSyjKNGSD8ztwv5CqJgshJ
PngDVCn2rRDbOG68rYL4Zd1BM58TVKYNYPhCnt7SaWrJK9cDN+DJmn6KQlGRzlL8

`pragma protect end_protected
