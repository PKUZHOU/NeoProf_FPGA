// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
FsyzNZyl+PeIEWONlbHH7Za/co1UsCXMiIarcNKvniQ3Et6hjUWMIAdFEE4QXKum
SNYDhzqj6L0i/AQAMkh6MiNzC7cKf8dHYw06qt6T0fidiRycWBkQTdrTOc9aEoha
TaCVQnSMEqhWO+ugPUfjBDX+8nMsRJD6C5Rz4wJgGNc=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 5312 )
`pragma protect data_block
m5NrY+oaviMjEMom2zs6p7Uyw843qeuKlK2JsJQD/SRx1lFEgmKFyLi0gFZ+/09j
E+1iBbSyX/iaSJUCprLzbtugIV7GQMC/zYtCJrKMZS8IyjU2LXtJiSHBNXpU0hXg
3L1PAUQAkfhuG2kIuPqBTzSJCDuKjhFL7Kb2GMd66rPDgecMF/1SYtMdQ5y6KCjf
3a70KjlTWDMrui5J3X08pNaSD9JgPS8YBS/Oho9X7TD1C9+shHiLMRL8Pt8E4SP+
2CuUltFq87lELh4BtSmoBblB+hMeyY6kVc/IPG9j5kbKQiKvOiF3+1GNxH1sHpp/
ZNmUDvLfk4sTaCqNNJT7kHCpOCfXo7xI8uytNct0FfDCwHNS8Ay8QttoB+9YLx7S
5olYqMv45QC8DiALvrmZO4BH/3Bd/yivHMjszp1zsWYOJLzT5ChWaYGuwcQLdB0A
YS2nRg8sRi3YpUDehfzvggnTHIUWoRpZj1rTmwkt5DoCxvP3qBo+7UrFJxrBOixc
fbghKMFasjMvUIa4pmtyQvdAmHTC34eFkwDlkoCmesJ8jgMdkEIoD6GFQWatVLgS
ubClxQCObE+/r7OoERNXJsFGnu14ARebNno3GxAqpw/Qw+JCA4IMd5KrxZfcmr6N
VvsF6pPOd+NbgEXYd5VXPM12MnhraVfdhQ9/Olua+xdr2l6fT9nvMOgUWXLYm0sx
QBaS5xYi3lsFdvY0ji/d4C3Nv2IRR9FCOHBFXdpG/XzHRX7JVF5VAqVwHKqb/moa
Z1+V+0DbxdGheu5DUfH/x0jodd1YjULcDCmj0hiox02rGX+dS470UmIl6rIuAPje
SvmQ7K+hSy8pEgUz2dIucwaNJWvZ315JJRIwdIctKczgtEow68Y3XzEE0rtTKau+
W/+pKv6axcxilh7RwEB0ghzTL6Iz+CjbHSOjrImK1kUWb7yUoCzMu7/RtAh+XLGg
uxwhYUXe+dKB+hMktOwXHt2wo77q/l7SLaR02Npl1NigQD7te2E3uNge06bZdPrB
49/dEki7A+r4Vgdst2pDyNvtUcWtOkeWSJ4lE+YV/PLIj95eABs0h7VKRXU0mdPg
ViH4YA3jQQj5/2intGIRDEjZ4ae76FbMOCqVO4+r/OP1b/PoTGgD3bagNECE3lMt
nyUtEHPp0jXyxiNw2NCYQ9VqqPMh8H86saJagWIAbNpaWKZiw+kRnWcyghDDE0ga
qIsJ+qNjYLBZMPNwMpU+qmPXYFYQlbCyPzpS7UHy86mYls2738unSWYzK2z+OdtL
XXY+HT6Y9kHmBWG8rpvqnk/um60rGPuYncbmYdoc2W69HneFqDu4hy93EPdUf6XS
F/sGa1JXFliYdGNFHoN+MwzgUSdhmV1PPOpGnoJcRurcgBnkAB0bmqLBdlaYAi/A
qpi3YKOSC5xkBiQIsoniQ4GYAtHODWtVyu6KmO0+IJEaX8slQVaRE3LeKty30jrE
RtJQW7QPmcjRet/4JoCJjlzDQSSP4OUfa//e1khfRe0iKs/CcmNlDFMeuJwnyCQT
/p9pPsEyh7ouplrEmxF5Zwr2fChWJYVSrVBt94hV92xblpbE/83Ugj2f1gQxAB9A
WRIag4bFRjEZ5q4UTs/1wzS54ckkw7UegTV5WQzcA8Lsm2gEBAf8eDw3Qw9p2w57
wmuqiFSRmuZEeuHNMvQclwQsvuJIoEbjfRu73HwYdoAb9bnKUotCXW8Q+nNiK5Rm
qMKhdyev0wPIeQMW9LIYfnMY07xeKFJC23rwYmBU2G48ooteLd2kIzTpfCbERXk0
ybAgx+oKnksCqnRR9SwgV4xfgppVxEQS0/q7GEnMKNtAzcgU0m61Zb41/Mburpyj
YEWsBrelXvAVgBCi9j4dk+gMmsu4CVzFL7bw59CBqnSR2aCwp7ClbaiAYYGzdCgo
x5xWjSRYHXqxUPsF7JJk0grz4QfxFivFCWY+F1LWW5FIdsRJ6MYGZwbPWPHrcc1v
tYE8iMR+r7oP6TelkpLFXE8tF6E8uytSpny0wCE1h3q8LIHdUct2IoCiPYfbIC1U
qEWA6bsn4ikhpV6U1S/SgYj2ksOU3FsZH6C9de715LA6/JBRjfA3G85mOzYgeU0s
9bo61miomc2L2rOluBaqjwnr8onyxOgWKCCAM57+N5IcShnqcX809HvG4+t+INXh
/JWfct/0CPTVpMn4oTjINYaai0JRyoKrVpJEZzTdtKOCpj6Bc9E67/OcSPOoKK6h
gTvolf4QHA27m0OtD38xSKANzBErAejhsQxpBf6Mq63O2l1xk/6RKAo6MeJat2oU
MZyNvbd5aKtJ7rnSLJvb+IqF9XNTmWc22kqngM3qOW8+PrI7HvCjmyJooshXPAt/
hU0IcoXKIXAmz5UEVkoc5dnV+sZm4aG3DrgEJdkO5OhuJP39NPSrdwUm+00hALdA
ImhBZhGl3WmuMLmpWbNxP9JZcl+PGlbDmbjeCeBHpkmDvpr4jow47t1/HeoCEqTH
1asBDqM7PUnAct/B9MCWdgQn94HDhnj6BfspjBg03joNP2PnJlkCwbvVY6QdMTyp
uKYVZ54h/OmT/REgEjPCbRfAZPDpl9Gs47du0iyGTyhFJ2oOpfzze0oDpVzRZJvi
U0YDpfiROB/EIgwgGepA1IZqKqLFm5X1eH1aSQ5/3hp5kmDGcHH+9DUs5/Mp1dF+
NYfuxiUO+LHgm3eOlHRE3YhZuQ9El/objr1JgrBgmHCFmzxMU3iXQ6ACigJI23Z7
ZKArK0eQu1s8DiXOxAx7/JpvUYQyMi5a/TUF5WYLS79anqQt1Iz0TzQoAgEuaFOc
1qmwRBQQgk8+xF976hU3+YbXAkXsmdXXwIftEkefGGVKHBb/buCe8c5CuYx10khZ
7GAGbt9tJHhlsbPPJkN104Zar8mgHzPOA8llThQPpIlr6Djt4CO6qcRGkTsZfiHn
pB1viiIbI128kLeG/GtEgHSrN0QuusXcSpfTevGZp9L22kbfTHLIYu2LgLEvFfN1
92sgTbiewTBljZn/VbV4Ee1PPNrGtgarxSbTYHskNkJPQI/Buz93zLE4VSkT5j4y
ymsyUxzSvVDQIGVW3NRepFdnu3HOWEJxDv8p4/Mzk62eL/4Ffaypv6kgOd1izNIS
Ds0w3lP2/YTerUFmuTDyS3agjaAt15b0jAzko/cd3qfkYhm+QCpefLQ8M4cts1tH
5ssCPbCaXHT9HZOu1X3Z6oFi1ccIRU1aAq3Vp7wwzqoeFd9eYX2T9sti1Z/TX3EV
oBEzXZQrOM6HKuM+YsdfeTp/LNx/hF9n8hNW0cqKsWM5DNfhiPhT5H+P1CVDJ38a
HS7fDEYtm/3DK9d3734JRaV+/j09yoLf0IPd6M7HciS6C+lkhZDF+3SOp3TH31Ma
yxQ9g2yMJLeC5fwAlDSTZ/01Is+1exKeSTgN0a3rpybZSjMdPLCIj6mWoQfDBMqc
0JVc29NhihAaPNUYyhBhT3nEXN697sdHnnpqt4afzNt+uvOtNjtUiqYUGJ1ex10t
n5dfiWgh6BgPkAdsav01gHimJ+YJMfamYQucjzdhFpvX2Q+Ohw/exVlI1n2s8kpz
2LK8wVj2hxz3LgXYSu2e6nTs94ElZYITi/s9vYQ6fSxt5n7EuEGNg2hVqRLMXCSQ
plJqzxAj/pgtobDhwl9MeUwLqEZg5d+VL+wOrn1BmHs2XdF8YtituW4FnfW1YZOZ
8wE0LTMBLPP2OPCZCAvEwQ4caEM/b8A+LQMP4JtB7JczgbXqFMPsupKisKVcLGv7
inWRaSB1Udgqip4AuAq91wqWggl5UaZpgWbEF1gpH44oy0e0Wm9gO7xujlNjU+DF
A7ROVSrgp9lUZQ6UsdHmEtDwPXD4n9l9aDz/Xyq4qvq16r2U1N/T4klBASsOcv82
nC0hOJAGXMn3K38RvL2nGfvH0uuMxtRxp5lwFy1zdPTcqVhV7Wt89RQjw9aauo6a
Bs1YNLvMUQSAYo/eHhwNnDxuf5oXs97iVV5mYwSV3nQo19hcILYVWbzr75RnniBj
RfQijuWG/3Inhi9v/JPvq5VO+2lYZykiRvXzOiXfRv+DO6v8cRCQQOKU0P/xYaok
kyxz+DcRRMATNtYqCY80nrBFYaLehi+vZmxqqngDzN2W7A6LLvI56MF7g0qqWybu
1f672m/8HqlQhh2yxoouEU0XrlddQWym4zgM86G7VOwRD7BeyZdWtnSiOc60ysWn
j0AyHIpDcrkANe5jlYtlH2RJX4k6Dlfj9KeUrgZhvOc5k2oh8+4hJW0g9VLIAj2M
2E3XTORr0gi06ZITaEAoKrQM4Ds+bEVglPFb4JV0MmWkMAKiorvT/NAtLkGnC2Aj
ERkjIF0BTE83uPQjV6D3eJl7KjunG2mRTocXSYjdrNzb+CLLdX59hxGE175bAqej
kIONEd7pCMm7DtQz8CGlk6M3GOYXWGOh4/QjKMwthx3k7O7mylhajXBetQhfTXkF
4pkZW9/FpeJedQBho+Y9qBP3IXa/vky68bbX+U4QZRe24xA/P5V0lnuwDh39dsEc
5IpVijc06jHBTmUyXQgeqK5ZbnJl6h7eekCisKweZCU/p0R0u87zIq71LHgpRPgu
/io0NLhc6fqmyEZe01b1fpN+qGOPNTc2NDntgx41BuSO2umtPU6bOiyMr5iMkL5w
rnU4kUodEKmOfqlzCr9lpxl/pFJBnungt37Xq9PTbdfF9+ci4DiEZQX7/lx2PGr2
cxVmwAlTLWGdTJlEfZKlNMYN5fxLxo8dXerFthCi8dt11o83mdwD7cDNpj+O0ihw
xqP8rfj6G8NJuCwA8s6HPY+5lrq5mmKSW6BWdr2I2crtpyF9VugM7LPAUUu4VWZr
cB40jADwCTa3pDxhbWoMvt9qpxmvzc3zNY7WjqifX2SfikFrg5hqvvSjlOoxkbwL
mqm1pXIUPeBgp6pKwKhLTL22S5z2NkHEGJv2pwA2nUmGPC/oykVw1Bhb93qQIvuM
RrrudbYHrUCCrWjBFeMNlqqhd5EXZKAiE8LTBXoL46NDVjNHB6IhD0yE/z7xTYRc
bhkcaNkpD1oQEcwEQtY9rtLW+XEQ9rIHnHSfJpHsPpfahgBOwIpsisEMV+RrTa74
jiktGpAl71bORSkBB/HtyQDZzEYcXn78q9qQvZAuQmkKApm5YXkYGwgK9RANYbgE
6/CncB8N9r4VCWcIJYk2ZhXV5aMnPhiJRCAWsfioEeOBAMgSg2crrhcO1RwaYB42
oJGTfYW2CdSD+mfBZiAWjRVOmygwgYNaRWEKyyMQRqKXELnZRZhh3lsEC1DONU90
O2yzuhXjP6qG4I8lzsTyCaAUgZl5qr1MYiQBeKRLkp9/Lm7qgaFirxnKo/muMA2R
Dh416UggPutrL6GMFtGk+ZQ26lLWGOm9cqOHcEvb/LW6nkyTGM93QgOkgPZPAjFj
KtcmltD81NbBODVOp41X4azYPbqPnndvnarxItDYrAbXJoca0XWW+DwLB7aNExiy
jln0ou/wfLi+iY29WgDqjlc9rUF/qbTcVpbJeoO75NH/TXQjhQ/y5xnuTrsugLgL
uSepwy9bCIB9kDFiEU7m5/q1Fhb9V94i9hmmjEVnFFcAQioTV3qkNoOS+LMjMTXc
vcjuoBLF2OYPtYTIJ2T2+HnbduZRlNITGkONcXXPZ7+XszgLeidKTNEjbTR0YnBa
g56V4XjBEPoEXHUT4k8CyPJ07h4zY0PC/YQ4KevKWNLIakQ6ifnlCgfasFbL12ex
y47dk/aX/uQcLQV8U6TmFGXQjetDMfCefk4lBdEH188K+Coq/luYsVH8b+jcTa/D
K2QtgMPNR+WTGn58qONxfM/hoP1NmdSyw10PctclWuPra5fcZFuFyzS/NkHvSOMB
uhETkHgNebvSR6kDql+z+jk8ZfuzainhdNMyvokhoLKEDW0C+WOJH78RIxP3ODCF
p7MezP+0ZkijbSGctsjLHfs1IuaID9IUcXNgduNIfHM4zHf1hnwg+QILrZEyatoY
vRVoBSKYTimwp8MvjqJQwtaTmjewbwXhVpoZV1DzD1yTwUJaJlyxy0X1LvXAn0Ho
Z6RwgeKZBbIdWSYHh0hbT52iqZfMGP8gHnuzDlCIneUfQLMrx7m5eyLJX7JSC2Wf
wpdWDsn6dpREZhoEiyh9qx1Hqt9rxTQmi8b3jNCqDQpRknzJt/gSimd1+2NctEp0
9ChHm2jWpnbP6Zgp1o8K4GzqakL5Zzqbu8jW1Mcd4VyXN63XVI/wr2L1Bde63DKP
8wJeIXAOu+mtG9DTBbmfwsKStkMH0CVXewRfK2mak0mPueemhLSJ+atuz99u+DYx
GWuJjGzfLxj+DgkMDhsA4yPmjwIK+4/8dkjBEeJSfzig3dtUtl7rDMCj80iSqBN4
t+f2tfNdk4ThStxoFEoVoMm4EKzinA3TV1msu5KRehZnBKvY9hgK/yU0amjpTp5M
58VXKZILWH7As1pCKUEdzxQjnYwTiu6XHgfnpAhopNyA2d9Ay9sFvakWTqpPdcBR
BZXTkqlQuF6sX89OUyzfhsa8zb+qWicpBdeQGkBT07VMPCTwg1+M/TDaJlMq7QOL
9JO1YzNLXDYzejid8SvskOoP7MBRceEdDS29+QJgrFWr0wVbYl9inU+VpfJjB3to
HHfvY15qbF+LKVwDgapbWswLwphRgpQ76KBeTea4clvGvCJxNJyBcUgfjQsXnpEr
wC9RjWhdfybGjTd3eZkx5FueyRQRLG1G3WLk0UuenjsZ5gRRBKAKYTVhcBVOR5QI
yC3cprQyZl2+LLLf+KdQGEUUDIfWvWNFa2GPGATd9gK0ztURVQA755zzYc46IX5Q
qRLXbFpDtu9cUo7dEsDh+l6SarSJMfBSkzEypKDH4iHOk4f96xHJRCfghbWt1UQp
A/hQfP3l79ZI+apiT9lqh2VlSr1V2JLApjauEA59yzNrfbamO0H42WI9HuKq9M9o
G+QPwKtVpV79KxI98GssESDPWilZdc3ClMwwndAApsaRLaEFn8SoDnrO4xIm/vTa
Y62cmW7/qY/PauQPoejlHJTlrsUH2Ph0YwXxAzg/Dp8=

`pragma protect end_protected
