// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
w42dnzpxC8jwig8RqR3zoylgRtzjPXG0TutLJfwQDZ0s7g/Ub3CV0kKbXqqXlyFS
IkbqJ50JEJMOfWRa1yYHLfE0sEJIXjsaGz6VnzQO6aZNOKn/sF0qy3Swln5cfcF9
ezDbL1cHNeu6KGK8M5NXG2z2T3sm6Ug4v59NXAZUMoHsJy+5ZZ5OzQ==
//pragma protect end_key_block
//pragma protect digest_block
lT04ti0VTmcpljstQklihHsF4DY=
//pragma protect end_digest_block
//pragma protect data_block
V0Cf6oFuCfO6MZXIKDj63R1DxoFYRptqlae9HuRz0yUzeOhCnKwD0ZgQ5ddAia6h
jywsWfXLxQGQpGcaOAmbdgRoRzBw66KPj3623byp+snrxZ4y09EoQjhPDPfVOeeH
StNSQvu5ZbGkVAtR8HfR+IbS3aozlAEBRlQiJbm1XpMkk8ykzzEdC07dezpfrKit
ATv2k66y6KnYwA6V6B/lDcuLnDCqjM++34mRpYkrpYw8ESyyax4b+aSOhpwHEEHG
09k3QhxXfkU6lPE21p55k5VaI7mN5x/bPC3ehft3ui4RPTM0aGRxM9yy8zrXAE6M
Y5qs0h826cCghg+X/EL++5Me1/aT5fYefKfVwvX9zYw45vSkAq86MPMacgaeKr5/
P39HX1mEer/sX+4fdVKAWciF9aPv4trCeusSIEtT/Q6iBqwm/8kkbsekb/NtqlDY
wxRoGj0NkPXFmFN64PvzAIZbuWoIADjinqSd2UwBtSsxJ3s3tM7da0ldoT3nG+Gc
sygu6SNAx5Myr7mNQRPSkr2KMTQKZTzqDyoiBT9jCLETCkj/hLyfkbKErXBdE5kr
m2rQCcv74iEodHy515b/wAzKOyDMalHXzRiVjEtFI8UC4xlvIMhy02EaKzaBsraM
pyVU24x3jsJ8X4N8/ztHesggvMzYuX0qaQZvO2FDXrRG9UuWyP58+XFpflbwTk7/
H3LSRd/zAOlttmajZfLn9Bfn8F32D1Ki91rzj5OMsIXsG9+3uD7M/ujKndIkSj/p
gQPlU5pBKhQe7iWNUNRPFQy7ivSW3ZfiwVTZPuIXWyIgpXYldkwXu7PdvaLSa6R+
AqjpbI2kfjKlQNHFsxb+k6ZZVilFkBjLsIX6iV7a40ULhIkDFW96A48b6sAm/ux8
inJ1lv0IJwwJ8U32enrK7Kc4OAqr+lAV1lhebvPR7WxrbYuhx15gI+mkOhJ70gX0
kCol1DQmrxKKNXl1kmO820XJvdITnbKpcVsl3fmy402uwEjKNRNLhT04ZH2Nr1r+
/qSMvPBzeATECBuwlHNEM3PbU6sA/tNgdCUFg5q6Y8cbX7Z9bI5zJMm1bPnH9ey+
QXo92WGWcmt2Eje0oagaEPI5FnSWLJil96GUljkMmxpmyDYKixVH02UcLISuQiGu
+VeRQwTCWNd9sHzHMnHcDF2mXfyGlCcl0vC3Q1WSrya/jMkaoN83QPDgRQn693FH
5ZvZ9KhfCC+nGe/o3adAMhJykVR2d61LGtlJrOnhSZjhvT6HXa6vb1ldhqsdccaJ
T+Ul4WlabSvKHjlCpEOCdTtWFP55fCc+n/0PU7Y0PzPRtjY2P3frV9icUhUgjIIC
e+cKKHYJBgpqTw6KRzwANMQEHe5D8hLo6wFP1dh1DFDT5YkWxDbEnVy6aPHJ5RyF
+hYVlizTRgJSFLF7z6pqFwZcBszT8XpGQcxeZS+n3HVDG+WBJNW2p/hZzHM7WVvY
x6VozHmbmHyON84tS0hDsF4bYz+4H0iAfNLnMiEjyzFBPyHc7RxLyEGzAkvq1Bit
zQnnpkYvKvApl23GeXiYhbQBmmS+TUPjHrPGZiNNIlTxwcfcpv2uaPQIWovU8DnO
q9DQQVjB8YtvONQj0cKx2sjCeiyxH6ZE1BsYmqKk0NpHB+tz5xeh1RtEsoHWaUX0
/nvGAbBZUjPFb5f2xpPpsUrauNLEyaYGefMczn6OU2vEpI4W6xUPq1uzA+w+iUCT
1YEQ5wSMewh0jPEAALVdvU0MCbeYgSbhqF+R2E/kYqIfXKJfSKbvvf2sxWC4Jtf9
+hTTb245++O2FYxjrppRHTpFLCmosdCyTkZSDH897AS3dcY7QghT2TsbMbuV9G0A
a89dTh9TL/AzATJLHcusuwkUR2TYOB7adYpZMuUWxN/rTN9ycdbVblUb1mx2Rk93
dstlPC7CAvfBLU2cCnBd4IBB373ocoD5rjYwaVqg07w9vSm0mH5qbzGbnBPalHAu
w859LbvpbVb4aaQRI2EO79W1XnuiWaxf89DpU56r8+5tH0jfNum/GGtuzUw0ICZT
I3COmehxWdrnvgsFhIMfJI/3anBvgkAUuAg6I3CExu8ESRCJyjOwG9P1Tp0dnwSm
e28EXPSKxSxpld32BOX4GZKkjFxrxE6B6RXShAIA8nLXugd857F5sIXb68fq3GoE
ERGL1/rqlLO3B819iVseKpXabORAtCe7J9dx2iyeFs36bfHGDIwlaZcLryRJG2Eh
vSFoOx5RHx5XwylTNLzobiL874WWWCs5J4bKk/QQgTL+CvShtWvJbkRzAi9mREhx
hoUntSWWjRFvI2IdFBqfrsv+LiGO2emaHQz8puDZMIOVtY/kTzQve4n8YEoktKMG
Y5mgqew+PGszwFErta851a3nhUISUaa+61prFSO+9wiSY6nc63Q/k+o6p8zDWgCn
Jd7M5TqoYJrJ/VunbvCb1X26mipb6Javf11jjK7Af3v4a3H8AEAgsJu+Oy29sdUr
SWFrZ0wa0LOR0jVnQzEmMOs066YMXB6AKTA8vaLMfHaBHtDanMlRLaoPbN3voH07
NnFZM+/xg+UK8KFxV/iFCxU6dGJszpjWrCUrCPeRuWHkDNGC2Fv4lJlihyjlnz2v
tF2LFTmGBLit7bxtSHdKOIqZVKqLn2Uqduo1zymm8QLWwQFQX3p8aEiOwSHXLcNf
gxscjK0I/m9TiPOf/t5pd9r9zz/K5GVRSpUbGVJ6sUwGpZparbekmbZJlPcIIxXm
TLMAjBq8mPD0wRF60Jb3900BaHuKtbCVaEbIW+8LrpvewpgFUd3aa0FPWmIRBpBl
8nCC346+4Tu4/pAwE5rhg/WSJU+9eSxzNYwsQ1u+ecLMu1ebrziUEjSS7wbuTu/O
2Vd6TL0pz36FXbqeet5bc4f8R5mtAjrxK4Ddx4VRzdeMbNZI/RboGAfNyRYZ7oTK
GBt6zo+Bk/5dEDOyBljmJmoM2EBJt+U5CQ3s46FH0lZmQBRpuwRc9EfKBQRJ9gwF
hwZrzpecu2RdMJp0h14bejMyvBLw6w8RliAJwPkwQVSb12X5FYr+Jmi+yrJakkc7
ZOINY84ju+qIhKrORA23j56QNmnNxDnpV8RA0DoLigDKDa29cHbBvjvus79sx53M
hCzPYyTWJWNcYCWdzaYcUVo+Sc6OLeGQfKwiWKsJ1cV6etlGLgK7R8g/MlAfOauL
PAyNXwIq+bXCIzwXnF3nMsVEsPtml17FPqwV2toRfBO7RxVEjphM2d/DdIX2G78T
r27giokFeg8C1F4/a+o63V8D17gp/yklOt9Dr3f7xeEZKmSiMXMFK5cBbwEubLRp
i4fdQrMq9oDQeAUUaGT8wuEnyFRRpfb33snRhcyTK64OAYMdlzUxsSWN7UQU2wXn
uDziQKgAEdPgrvjC+5UglT949dBWTvo1iIl7v1aZlO7AvNobYZFEtDKU3+Oak6jd
ZTnXgXGOGvmfOgBp+jrSK6A5RiFj5GzLOVZfECqWWgTVxMpmyw6F763wchmeqU5x
xmAV03MrEQya6s2wRM+96dMeuAIMInLXLPxPQvMbNRmnSUmjEYw2sKhAmBdAwlod
R3yaaer47MkE9B1mXmumxv4Uj1RUIgQsumLHUKSyAQ1r2PvxMUwh6XqJRL14fT1t
LuVjEriCtpiLapDI27cAmkV1Xtpe8BKMvSZWe4MAk9/uJKG3v0Qm0dnfbU7I51vp
k1UOum3z2UNpJHrjp+ne5eoeU6B1YH3baZkOba0uMNBIxyW19GFci24zEMmc/++5
caQEsqRjgOIJ2YFF+S7tA22ISVsvRJ13ti4ddZ5v9a4DtWPjkZ8kyblVLg2wGSJS
wTHm2KqfuWkEpSAq5CGqxo98+77E8Le9OMVmYBlLnJ0jmGBXvO71Z+TxPWbgzBPC
Cf/bVXKEXdgxyE73NjA83lgudfwg7SWhxjK58qYt5hN435m1lz9lFf3AtK99xJoT
CzfUWctCvG7cEw8IY+AMgMm5OAXuJxTG+yDotwryRrwvsXRqirIzcBBh4NJyuPur
+3PXzMfiUGD52nnM4MDzYyKusWUXmHh47NIFjfXfdqSeQBZRnsYSpeLkNkRHMS0L
Ci2E2NsFyDHffhg6sMlnXFLR4C3sPD3Dcf0YYqhKI4pmQ+VZ1Ke014t9rrKN256J
wmTGwSIfMe+o2qMr15suNBlmhq8bidjZ3McmU4EQ4Mv2r5louhKxuLdObjjMaiBa
MrslvnBAA3trLyDsc+VGL9ny8iT7rUYDBQQrM/KIUT3/fvL/7AvNA5BI9DqBq7IH
msTF/oTh97VheQ6MRvsJAv6MA0ffVkNOqjaGWladz/CcsRzJ5ENcMIHfDJ9N5OaX
m1wRA/30RtYlqRUaOXP5EodUS0xZvbsAea3AhN6MmsulK1y/CWEs8NZvfV/9W0RC
zSezc9QE+QVXwcbNSHZqnkeLzhS8qFuoqPI5RjujRXgIGJYSpp7MKibtgYVo9zll
z7JfL7n654IkdRtppT11gTzGO4lyxprJS01e87LSiI0AOg+mD8KcUz1+4KEYJLXD
o8tzkOpHwnZTUU8o3oJkFIkPeP5xH86tRpoH5YJdDKVkW9pOzvpXD7bNWeOHbFO5
OAW6S+JMY0imJ5WsoABKOw3eGWLkCfJduLgGqR/99DQr2qpycnnwST/USaTrni3A
5cNjW5vUMwMnG4S6XIH2NzPoUh+7WI1ovunY7L4T97YL7Y9GEl8viuN+PpndwD3t
qvj1ut504A3aTBJ8as88LO0kla2ZTnpTFP83K8NuM5ex/O/qTZJ1aaD3fE92CQOI
U0FVXmXLsV5Dx/wYZs3QrisCsecUfi3eQHYUjbf6F3KgrKIOAcalig0G9IpIlxSa
JIn7R62MMfdtQpFK+ctHhejHu+sKaVoUR7y6giE4ozj+WbFR/usMx+nz9q7kogPk
e7DrdrFkRboz5WbpFc7RG7Jjt8pq5z1/F6FsvBK3erjV0AQBXrjv7Hu50hUfbSPo
aG/qTyi6jKJZWxqeA0cVHZ7w18eugl5qsEd4tNwu90pWK6o7///xeJskysrf6t9I
/46eYtBvu8IZpYvRqzM//F5vg7KZPzjXB43NdSi0tjbvu4+UnphAYb/uCqF3YQ1l
YUUszfCMXzS5Sx41MmIwG/+1YIlEC0fM5aziccpspUUK7npdMgS9/LObdVYoyFPR
82bHWplELS5OO5m6rzBQSmgZpuqPfGJpr4ixBn94YbitA7dFIdtc5in64QQqFUjX
jw3vMUcZ/bujjEccIxeKItfeqQSDdGnpTiQnJ2cUxS9eQh64jeuGf+2ryOlWZ/Xt
YtoYeFg7K0y2wwQhcS28dHqgm7L1wucxSns6j8BNs4gEK2P+06HLmcojeX+q+dQh
8fmQ4qJmbi6FHktjyJ1Vj6jJlsyX/HF8V/MggD7+o9jnkZj40LqZUWuEGiAOOCjy
x77AxRcPodm37iGDa1GyDCOBDKlMlj3zO/KE3mt/edQlEKc16OtSJoApN9DRmzHF
2Qy1YrtGOKDz00dNUE036q4lTz7iEDkipYAweUtgw1uy8W/W6g9gxZ0csS7LyE9c
adRuHAtgIysAYOGWDaXi1N/KKV1p67zVWxcDl9wMxTyCIpNzOTGdcIGcO8qGGZ8n
EkdkV2yNa+IANHXb6w8z8cE0Y8p1/n7YsDD/rAIAWMRsAmDPwZxvaxplTF7s7f6y
SXsadEdDhsf4RbwjxYmdwZKYr/DQQxuMn2yFLW/owSPbAJzmF4k8FfcTxyjx+H5z
ApYvXESqY3YVjyNP0TLOgZNqGcwG2L7hvZc3ain7sR/WqO4lXJSqjZ9VeWTE3fja
Y0gbssGnqgw9o7cUkOVCuvUh0XTr4jIrPeDuahAOFXQAAISXWhH/2mulQ4+kHvcB
ptBvkOKEPEjwAheYpCYfwvMgXsA8PBsJCk06afVZlm5Xx0CYWtErWiAB49sZuWDN
m0XMWmZPYnaMCjQ/AYkTc21EnNdOoM0WwlD3iW2RPltkZ1EJGQeLBEFSdUASRoFt
xi/PpGBfu8ZhlmPp87yuMeXtkOuWxYgn+XdpO+PruS6o5hu3nSGBqoqXkYmu8/X6
9gMI8ONBN9pjMUqM43H3ZzwYniie34H77Pvl6uVaf22UF3TFCl1rgQad0FGz/7kh
d6C+sEqBqVIGOhfqdnAWurxVt4ftjjK4dhZ+EgFVJDqj5OSar4M2nRYBUUeH1LjL
27HpJLSZn6JF0LBFmeMBdIDo/xBz3hcwZp4DaIhYXvigASgBUatC0cxTPJkuvkm7
03oWR+1ct6ygFCTCse8EXkjatrdRihdlNzJg1CJHR/9hictOV+qa5krxHD59Fqmt
i/6L0qod1rSzLr50ggSHFOHG0pH1p9HBO1FLcKhq2mYswo7FrT549yNOzggA0A6a
NvOKYggi+8//iUtF7Wf4E23Bwh2vVss1I1RLoVHYQDGOrEivYP95/pvwHC/HdiTb
Kf0yeygQ6NmKSKZHl8XX1SI1xoiGwmzhB7ewS6uzMxJboTIWU0KpFVRE/YeJLvfO
sh/R7u5MTr77uKtnVgfRBgXdSY+VBADGXfwfzO6XnJz35W3/+fMLsQw8z0rRE5vq
z8eu+VtvAVqFg2N8V3u6WaaVDt3pcCMy1D95ULoBXovVsXOP1Y2nCpPwUuKwsmSi
Kw8IH7R6rkOlgiCUmENjGDay4QjNMUJVwKAyNkVbH/ZaNH7nFCQanVAtY0fiwRAj
CH+nZAUpJ9tIT1sefZeuiiUf+gFkFU4c8DKGPTzxQPlOizJBiLLtfiF3+4C1O8RX
R8LIzhxJEKgJmX5VgM+d3o1S6M0i7SzhxlgIrkdJhUNts1Uvqo4iZLKPm+08baV6
OSXIa4vl/J9CSaUA9hCdOWoZqMgmKBu4t8FmCdzJ9GFujelYpSORbkwKt7wO1KYV
OkFAzotD8Juv7ViBTxeVLo+yhvrnPalg6R/Pqu1Qki0yYCfGivJVv/GHrO3GNKC9
nVg8RK6phn/viBH3H4K7syqAHV5XcERDiipPpK3NMGx7AyLpnMluLHF3kbm5BEGS
/NXotDGxngaduqcLirZmMM8cwJGQ5K5BFrWbNLcK6w/Nvi1TBSAkOBB87oxdT+ne
R/sOpBGtiMIkER4GKuFl1wuoEsdk040XrOy9/19PcoABspDUoViSKjVIbbgHBSqF
ZJ6cXYrW6ipUJH875HE/tbRT2Q4YcSZA97Epu5PegSNdO1s/u6QDkviBbwz3Kb+y
PBL+WYyR/SgadlCusBEza5tyLZq6K+Pibw5DdZnaRigPBmELRgJ1YAwvsChmugAi
z82i/3H8jymbZckHbUNalieujB5DEyu2HQ310Hmkcnsy15dAOxZ+VUGS1z6kyG23
kkLRA17eTy7/g3zjqO/9OY7QiRRHr8kpyMdL1FlBZM33D/Ly96NqIaJmtYYAubqH
NURpSU2ONv4o5ZSrnljx3fIQoq8YSNN1Mkrzadfw3Q4jjXJD/tadKrhpJq860ucO
BgAramyCjM2oH9zvo/FQ6M32yv6ds+vOcuJ+IxDmsrXTFvwDe6EPkOEZhMmxMG00
Ne8b7jc7RgMyoeMfmG29zaolkjWTtUpNTZ+a2/u4Zdtz46Gh/3jwtQzJzOTURDic
O97A9FjOsPsiAgF3AjhbiodQP6jiJNcLa6o3JOA7aITiCu4Zb4X/4yHTn7Mi9Bqr
pYvDuwQCO8B5cAywv0oTKpgX6p502Gv+gBcx0EN8qgqwGnYQtAq1HIA3M92+olxS
cfNLJOsMLguAelb1QB6mwyNZv14lQxwUeIpIc+Rw78drq0/3y8P1cdKp0mpCgTSy
Pa5XoDhz6R5apyNsHO3ZKO3fHQLBtBoyFpgk7jgbui05nKqYzz0Ae0+yRmQC94k2
0IRsJPjoy36jWPghlG1wlIPNtutgq3jP99pV/qbKgkXfvdlLZa8Y+NryXLbZlKs2
bgWxwGE7CSc9HT4Fvn9lxuSz31HkPuO+lF3+/atq85mR0lHIzzaGfQ3PBnLy7Wvd
52HocqZRzdqX6U0f/YVBhCyracAFPaSoUrfQK8Iw7EbamdJQE26I9GJcKf6S4rcp
cucB2ufelhCmo0jdnhLTcpQW3F0irlCYs1LYQWAd+Xs4/yfHlYJp+Xi7Yt3nARCT
hWlSJc7ZJhM8+ldP3TrxrMxsgSxwMNrc0Q0S7hkSslF0e5l+hErsLvwtrm9OruGo
dKkA+R8lv5oo0SJB3Xv7quorT7ik/SdOBoUIwb4De6A0ZwJ0gXeYUDWVtLPBMSEQ
uCQ0orLswakimzQRmybaKVtNbWI8DBusN/XM7UuO3R7QnyHl7JUa8Cr2/vy9LQeS
I+CsHWrmWlvugPHIyp4hjgizOCsK7agXy8QBu8Iktn5HqX2/Gn+04AzI431bxr/F
2F9TTLXbdIEz3G91+cyWVO6J5VAVd5pPTNLDQ1vrp6OOWP/B5mhILs8I8W+Hky5y
wlWtTwSOwqRnD6G133gVImrtzEvJ2bB6RBv5fzCM9uNXbpGllcFFJpPMNR+JZIj8
eFOPMvfILxcKa5vKyrTexdJOMSxjVbqRuan0vd+kfHWr1Xr7jqYkK+wyM17tRXFH
s+o+KmVxhC7rnyFZBCoA1jRZY+hLhUKKwYJJlHqQzVEhWuxVwmkxVv3RYIFzC4Al
pKXx0B5G7OGvjxecoSJu5gJB43maFlcs3BMaRU8wgQ4N8qXwTEHs3CF2e8MQoa6T
Oc2NGPKmY3blolCeIa/dlP6GhGHGf3zKxSoj+kDuBRfl7PP2ud4/ooNo7kdh5nrI
hruRO7V6MG36+bJ3pDc20nBXfiakIVp92KrBFiT+/tDgEKSBnxmRWJ3cVTHHjjW7
UukbuuSFWzqxfbnGiMeuD1xv+RqYowh/cqn7fu05PYbOKOzE9zO0p9G9uDYh/1u0
RZBYxPIVlSCNOHYNmzn1MjrTCLYINlvUbTn6Ntntw+wytRStboXc7MqobRTR3uBi
0qckRxGT6d3Jibn4+a0EwBslizg25W6f6dVRY+bU09dJXqx6l2jcAbiTOyEQ2jL8
lWMG2JS7cLpsm1gSmQsQRZLW5k0JypdQiTSMjBXtrrg3znorQC2eI4VsDMntjWX3
A0VlAk2WhCODwxsDpq8SnS49NiBlG3AIufcYSS1LOrtOxkqsMBhfGEKZ4+D+CX8h
FZmJWBlbO5BnnACN+lS9aaKubU/tEz1j5bVZxgF+rY9GK1qzCLC1tCHuaC7pkmR+
Y+3ukn9igen8xzjl2Q1vT7QQATN4VVOYmsMsErP4e52IhjHPkDtibNGguytRJLqD
yb7dbw52ZeazvXpwn4VpexNvDMeLTCoKBsVh/nZLbQ1wm0VGTyJcUoLtLMA9x+uQ
GJPj0T/jiBUZnLmTtrnxnmL3wlBy0FETvGbF/rw2IXrRcjUbQ64dYAQ4YxgOG1gm
j2rQ9ukMiQ4J2DBry6jSxOtT6+owDIdJdaToPpUMto+5ilwvqcTQ6gf5yQSyZlO/
ZN5cbka9hAJClmM9OzAZUhf/5+W4JeVyz8wD1sHsH16981MfvTqfhzh5TC+txhXB
x0bQ9GVn+HpC4PYAnY87WjT7iTB9/Ah1hzOjaseWQa6dAAOx2GvfwXT+ak4WTJXj
8jI/sSUgaqrk/SVhm+JF8fmpiKK4cuPU3rDcaz7z6aD2l9IPfPWHLJReB3ZhhU6a
eb9s48u5dV38pO15AKW7m9YuIiG2Nyxo8fXz2zmvDZWsIGEOTW+rxVuH/5U6vqVs
oquM6T0CR0bb8SnHlcTHnnJG2BfrSUSMTLOcSLEYfithwhZOqLylxf06VfoK0ct8
/e09aQovRMm3XIALwQ24F8wVGaRUAYUSk6JvHw1lL359iqNlwM0XXxLhL14i80Ar
GkDmC5RzPK7++0V9sdy5/Xc/tsR7ktgOi8JgmanqDA1fTxhgsjLzDz0EhsHySy6V
ZLLenD5BdkwI0gD7AiqW4nUH9EA2KTBGqf2okFqLFBBAjimFdqesrnddGFNGx106
9DEJ0Ei07rHg2bcKm/uwxpUzOFW61HGi9Uc9sSsYG6uH1XeHChwAdkYqNgw7orD5
oc2VlCPeIB/SACOPdkDxDFDhtlXgPnipjzICt/GHT52de+6bVQCwvgmRIUhAd9dZ
JSbPyfxnhemQxYelFZWo0cwJMSk9zBVbEo35AEe5QCrpyov9jgV4edrWJRHlTVow
A1a1LasO4ihXcBsQQ58N5HBvfa0Fz24dFz/xjuFif2Qc36EQJ1ZdZqTQABY/nrnu
8ZGcyrMUxUqVc+T9zUowI4j6rDgDLTAjFKGhg1+9DBWPDr7V5YO2IrT4drNfVKi3
5zHhZnqiUdH4kCla7gWeEGrMPERqZYC227NdzUqdvK67uVGMAqDT+dC9fnRhoY1I
dXNYhEyiUskRVw+JsnGe45aevHHUqjZog6bMXnmOvd6zyGKiDo/AMwvmef3/2KCE
Weji6EQqOpN4t5ETKHjvEtZlaRLeN20FUCg/xJSMh+sOKS8swCqNy+u9doHwRRGM
RuTqRAD0NDY7IcBlII1ZiHsDXXDgIyoktSdB3AaH9ofMNkYeMEG5AH4J8Xsn0Yxq
dz6IO9+TjkBaWApCrcEAL69bZFj7Tqjw06My6HYUQmP+L3GWCMEBj65UqLPFO+2w
q/tdzGKhBxc3Dm6yRiQ4UwgddvKZZEX/ErMrR7TxrlRZ8Uqmw+sMQJvNc3qCBcfW
DUV9a/SyT4rFSWpxw4gEAY/c/ofvVVHeHvVIeF3t4nle5rmmNFCjSxRJl/hNIeSg
zQIzyywT22ZTZUs0lhJsH3QRlPFTeWXiKT+VuZS0uye89Qnrp2TbZzC0C418dAbD
ZWHC12944wUUDa5gpJ3iC80Cgbxo/uehko0oQPAu2EL4cvcJfn+sAXWqOwcJgNtP
8GzyhhRX2KAGMbEijTCGVIxf/+8BqaNTYB6U8b16fjiFDzQb1/XGQ24GKNdJa5Sp
fBH2Q2RYdP1DrV/eNT2Dzk+ijCAkZS+d6zsXmDN39dHAVyODks4eCDPTe5bwxDMz
Q4aDfi1xvi2Cr15nMXTqEI/ZI5/DnhXddG5pOSgEvLWWtlzdjexpSzv+ss1tm15l
/bM5rSe27kvrh4RXvUa3XxKmYmEftQhk8wScVl0yyglB+gNy2E0LXxY/Vv8Of4Ln
aRsYwynKEdieepiBut/xIeELbXcSS68ExYdAEXdHzKlYv4SwQ9C/7svYOIavANSJ
58UPCamzhmokBWrKd62fEKWyl8DLakCINTf5c46C3i9d4GYqsS7/v61Qjks/P9SQ
cYnJFYvQyX3p9mju2askJJX57e+JLbstgR1hmel+6CURunZjP6c7D7Ghm9iNJWMR
Ave79V+ie8Ux4CC6hmkm9PX+ysmza6c6Tp+zXF4yHFNP8+H2Qbd8swtDcbL5c3nQ
vVWyCsD+0LzZkh4syQEl3Kq6sgHC64/vtb6CjAARdmqCxT30yS14exn36W2pMGq7
8VoZVv4vt9V4Hj/hzteMLF+DVw8Nb7UYZG7xEKuKCLC8N/SHfpSzaEH0NJaUK7MC
UXgHV33eNhhJ79uaha2G3vPFil1GjgfXKnu2RomWHfU2HWDpz0d2NLFToqjKbhkC
zq0Z6N20QstRze1J5Mn9+aztKoeC20tmCjGVaEipldbV7/7pUQFr6ajDwGUouo9N
PngyMg3OxDJ6o1o3lVZkFaipkEx/n67vWiFnE/mvLh6iYPYMHRY680JUqWq7UnLP
79Ek6VKgKdwcPLHlvuw87C6yKtBB4gWBy4pUaD2OlIeICYbKf264UTvM9E2AAGPB
C0D6K6r08Rirl8lLITvnnKhfFERDERP6pdiQqx6zgDFZ74PMHraz13o4GJ3fpcP1
pUeJ0mGNC1VM0DoCSmnFcnnzI2TMx+80i9clJeVP6CqS5+E2GRc+glf7GhRgKzk8
d4mBiG1+rJD/cxjp6WUo2MYTg/fxjSZf234nAIj+mQAOqqaVNA78UIdod1gyn9yz
XcSmr/bXt2gA46pqB7RB3Myrp4qm+4gq+mPHDsS8oddXsg04V4vsbhep+Fbp+yHx
SL3wx7841iVmuu8bAHNQ9E03tFkwlSz49vv2K0zMbn+iEaGXq/nKvEkcYouPR9Gp
3mj/BZ5XjsMZoYjIiTO+ZySbqNbcv58N9UTgZvKxIRSDIvCVlXmtQEIsvt8FipTg
tNbxYyhau9jiGkNI0tpnPubazaEeXVwDgZ3Znw3oalREytsCEPyhFgKYR4KlqdL9
cnUAo0u8vGLhgSmzBvQfCyusrC4roDAx04PnNIBpKpPRAnzfFtUODhz3/pjQGE0o
5jGUPWwiRy2E0MeFStljLKX7LWC4hEXLht7P/omkKcY5QPcYG0vd2Ee3wUdutxQ3
q19VlcOCuaX5AiCm8VSukvGKTKvyd4ACn+OjBhxoKwsffh01U13oNN6C/6O1A1fD
Dy6llCEqwcbibGIogHRu6+MH5kqLL+YOHtMzRYM5w/d9jNvg+8274cgwh7S/M4gM
OHMkqakIYBFIK4uZIMq2GNg0JpTqIMgTM0iasUImYYkCSWNv7GhrVmNptH874GrE
liiqW0Lj7d86jH+T4FRn9ho/bd4kN/p+zsGuhl/tpO1yqUAz4KBGDgdi9c9vWzqp
P67H/LEXjWKIEz7R3WMfwLVRwRwgwtpLbeqgPnZDQsSBppJaci1b1VL22LnR9psG
gAyW+T9mq0z8BWpeRhClYzZ1kCfH7CnoC20+SR/5PQESPm3YLy3WhqGzwytZDUNu
FRLuuuQmuuQFqIjeumzg0YgnWrJ8Xr9J1DOzjL+4ANm54D7+UDxUSzlVdVO6w3hA
hNDDStkcIJoOgCjBOo3skQBabCgq9JgGoWZ1+i63Ff/m902LHdotUfXf71V1KEQ6
P8JAh9U9zLBK+4LL1OqPndaOgXUHKipRonBjkGwiDR8NipfPDFRHe3yvDaKYUPFM
PL+EJT5N2MIQK32p8nkYIT+mv1KLpeEeH3SQj9kn2UDsiAJNcxIyuVFXZDM5E+3k
n0Yn5VjI1Iifi1JZ4Sj7aRHx0RnBSSVU24PlTwMxjTq+opVRr1GVztcpW9SvNmhE
gmJQjKaTkcS+j1bPYUYmxtKhwQTeERiaZaoT+b+tUMsa7tlNehMTNbN+Z2eDbJaS
/0lCPzeAV7W5TAWjkJ+FWG0r9F6XQHeuDbfZncfAXMfhQohhjcchWfuHlRdkDGgs
zmhXIB6IuoevZaW3qLIjYv2zSd/bHLBD5+4BSbhgO2AoiVNO2nwIvaZ040bTQGwu
Tk0rZjeKkfNg/bGy6Uy5AV/UKCq1wPsv5d3KfNV+4i8QFIXfKtaF2XPzpLnMq4Sr
MxGRxH5/LIwlN1HuetpmNETt1IRmdse5MFZd0ju2KFfHthc2Uzm6pVlxRTvkadOq
skygOAzHZjNrPmCcAqbAfu/gVrt67iSuVg/2t060KnfQ534VmxlN3k1PYUvEdw5e
45Ms65Zs4NF5xdm7cJ5juuyNvcROaTvAy+xX/prq76fpvLnYZaA3Y8jVnx8VyIL4
oO6T3jV/MqpXQhbxG6XUgqvJWkKX9pumf/huQo9p/4kvlFLPAHlDszQkXNfOCSCi
71/+2bramEnqMfyZpoqGeCktKexZyvQBk/XPqf6Shp6/6ZBHpiNysBgR5jWGUi67
9nE8OtFbB6f4mqBqs0I8NmvKlt0OUSCtckk2V+N4XbJP4OnortDfI1pQ17wsvoSb
uJP26OrVd19+w0cIwFZjSqD52j+GkyMJG3+l+85WgHvUsY31Glb12LkaPQTICrb8
wXMXAF2UMs0t/fF85Jpdd9+9qat2VMr5Ar63rgV1+IwjnN7siTglJHsf/XVaGsJw
E5jBKmXV3MShWe5/N4daa2GXX3HNoc3/pm7zukF0VmP4zw8y5PwDGF6zs8r4+ghq
78LL9zedBIkiZh6mbEokykKJXctMCqs+q4PAfaplNjGfisnHUihcErL9oS1wsoGs
ofYpfKeqJJyjhLLbD3sZvlY8v6cZaSijCoob7L0fz+SKoWTNJ/sCgStOsqkRfXMv
fwJC9Mgw4QNZxyanyIZddYjIrujHR6Dznkex4NUAi6hpq1rbQHgKM0myWMb6OYO9
+v/6nVhqwNKBHhAQMVt0g8g4Mw9kmXsCjRqoZIityB9DjUDnCXaKHdv9UqGOtJG2
01qZO817e+10FYGiYxFny23kJgpU+nFlStCCYr4uw4hFNQkI2qYwSIOuvnDPwjAl
9RgeTX3nueGafu3PJw2nJL3mhRjn3PHbN9Ukvl+g0k6HTVx1BQE85/KyUP+wr/zf
rV9DhGSw0OsxF48uVh9fxLeZ37193SooTYjO0ANfi/VypI2KZh3IvqXVtORI5JxP
So22mgIuRVYcpvsOwk2Xx2mL891L8OPsKWEGa7hRz6196qUTVKcgzgiH68+6ngkh
XA7OnPUNbYfq7znenEAEQgSFYu71zdHIlKZidii6VpyHPACBOrOd7KQEQxU5ZjDp
FrhKAxzflI4UrLPuwfZBV0jNTeU4p1eCl4a/tAuolOjgrjlPArpvtoDENvR/X5A8
TIE8PQ/PHZPex2WhtEjPXWCVGv2OaraDNGGP5LNPPJ30V+DvtccXquLidLwpnM3q
i1sxCcMS1kBnih1vYcX8vsLnGmd38EJSyrc9NNstDcI2vxETo4iFHc+bWZ1ZP/NJ
pwGmyO7I3TaMQAVRczly+teS27B+5zOnskL4OdJETxzU09Wui/PiUrDw8tfCtKAA
S4QOtEUw4COo6BHSgzPy/YvANNIJZkwqmDuAg5rmD9W7xRWLURS0hvbS+SKvh7Qm
/Zn5H0/+lmHdFWZ2Re5Y7xdzuzTRPsuUiqLOCQknkjUPw/Lw7VOa2BxN4R/ts06C
oOBQsZL2j8edZ0vkqiMaHzgtN2S81knmwYgMgErDlgVT8M828xtxqOGWEhPFiXMt
iJbJvQrJnm6PWIGN5uKDvJn1TbfLXTgB9hLM+y31zs6WEGZGdIOJPGLHYkDtvCQ+
5RqRY2uqke04oHpW+PiYV7b0A6CuRsSu+zobpLZbHlfDn9p4/93VgL93HDiuR7UZ
gPCIOX58W5PZrcQ2zf+NWR3MWt5u/VR25Cc+ISYgBA3Xl19Z5VyPeMXdDX9mjCdG
m8PEbep9JsGTDZYlxq8Z7suJ1DLM4EyJFm8AWvncou4sJiD4TmNEB2pPm0RrH8wO
6YpusEapVKugNPlexvfsxzNST0o7tHVqDhwP4KZbSHKcGAT6zp3kn7QtGX4LoCey
livmYfqqkMWGhzCLegd0LC9kC6WB8fevBSfvPBpdbx7FTCZkbTjh9vVvsIwN8hOO
hn9J/BC8grdjURuRd1gALb1LugEhUpDzMjFPM6GSFw4lP2g6HNDsoSfzymCmWPPv
EFDC1JkxUUUUACXkyjo6fvbwW08v9WGnMJrUu6Tp8cx2PAposJ/Qthn8dzgEVCT3
ZN84Ufzl1wrZ2ST2Hve3ZvBR9xJ4Kyn7+/pzLiTx4JtzSqw7UvaiqZ5HQqVxFisk
irqIr1PMCYe/pdg4ci3yuAAlQKfCojDSHkrZS5vq19+11rMFX+/xf9iHbAbOb9at
jtJMm9viNpl1Jfr3KYSDjHv5aC4+FDqA+2nYfARGFo032yj0RrPZHbqPyyJ/VeCw
izA1vHunbuo0wie3I6YDxF2TQqhmFGJmq1y3Y0ZYx9Uh3PW72y/YpG5nfUhm4IVk
40JsGMHSm6BriGvvIK1oeuCTqfSajGFZ+GHGlbcvhVaSfETk9ZYlkb+/nGdnGjXZ
lhhdqDa0sAmYKm8lDoBzd2yZqcMRVXQ/JVdHDE5hWb6/E+xfr5JX+BdnBbqokBd3
XC0jihYTvOxEHBuMgRRXonbGL7uu0pfwNBUwRfSB6EKnjXZwE+DNQOktx4TLETER
4x4nhGy1k6gVaRRsWm9S8tvHxJf+kspscnj3HRjsEnAufGJ5cKKhz5X9jyNmAEZ+
0UbRL7deYNPkyvyVUrsn+yQQGbErIQT/uBqsIYFnIS06UsD3a9FCsISYRTMp/juh
vfy082UW03rmUQ5/aGH73/d5srnL3um/KVm8mqemxVR3KSnkosZMz/NZY5L2TC4n
FaGRfogK9UkeFf5Ko4+Vu4qksyxK+xJ8WV6hE0rcqZOZrqsW8eSYt4OU/SAUJiLm
153qKKIpl1YkgQvCaYAwLk4HMgIGzWrRSjTKx0J/gF7I8g7qzBS3kYYQVwM4Ohof
wOBiSGrBYDXdmfpEMs0ya+9hKTm0PFDyy8vKPbiz8kLEAeaudyy0MGi120hBQ0xl
b2ePiqlJ2efMqFTgphFCvKIEB2oXdND8zHAz5tNKu4/eEUKOp1aXSD0BQ7BbBbvC
wMehy1CoO8Sck6Jva/P1IDeaS/tTsFMb93DcoSOKcYvJL0bNOlkrU8J5od+J77jn
itynFZTy0532GVc/AjxjI8PGZ9fL/2JM2X7VwUUlYWOaSRmBaF+oU/hf/qB/x0bI
+nVvPO7vrNGUVnnsmy4HdFah1WNQ8aw1pXT/w2nFBDZ2wdH3AokQdR6NZ5ipFO/k
aUQa0PW9l+xJRLTXWuvtUYRBW27oGGLGB/qJCbBzRvnscSl5CLNEtJKQ5vnqSs69
28IvG5eh4KcNpt1xrIAfIvAsYGolBkGoaDch3x4nU2yoCjthOM94s8GTAVzxbpH8
QAbaNPOmFA/flM+Inf0h1eUYDysltS+Lz9/EmqNaKfcCRSxjfSIckkvfkIkV4UhY
KAaPrHtgfJELW3OgM83Vev+Bkqa6TkvV1Hl1tsCMy2Xe4P3mv099GspXNyfDuw+2
im3JNprvmryeKC8ceEWQxVkgg9vsk8DfNBI1b4yS25vgZNas9qx6C1o0YHnn1yvq
N5MXkTs2N/GLCcB7AzrJFyfog+2HiRCyjAYSU+TakCIqkA0AQGg1/bu678gKAHZ7
36mb8Rl7AM9rKlCQ0BlhpZ7ltNNPswgB1HL5jtxQrjh8r373wdkER+KZMVD9JU44
ZSWg3CIZoNaveUM5z1kfJ+qi6eqhaxgUXos29PHluDYKlb9Bn050TlLCe9ZhZJ2u
O1hlbCJjrQo1vrzq9yQbtqvdlWwvCnYYhFpHcqjQuozVUMwWI3ZzTT3Ue/L4PFwC
4fY6s1iEP1lls443JBjuEBeeZ9g16E7fEIsOEKSvzt6IpykBns0lyKnPU6xLWWYf
iCs31XbW6zeF6dBk7m6iXsmU999CWKUmcCBTTwKeHUsl7lFAeYLm8LS89pgCuV70
PUPx/NCrFyAqejiREy3MM9O1l3Hcsd1iKTqjKGciD2N5kG/kXW2Johpe4/NEhaiO
/IBdsn7wZF8IZxoj+FsFx7MLpBQqUmAC92i2TAqO2Y3xXOX7pWer0cZTDH8Pl1Cw
K4bOR5S2qGKlDO7ldgqRgyJUTTVy4Umuy9nDqBeL7nJwdRwQo2N9+bcJoPW/c0tF
fYw1yTXd3oToIiQKTmTtfTTcWJhscPJYJtiEga2u4V962bMAHAvDVPU4nWjlMk4t
6R3O+7dxXY5IehqIJJU8Oowa+gBJfYSscFYHXFeUcATbxJWtwUED3gnweOhdJp/0
XfysTZWcVUZyF3kOrMx9Kwm+14dCrovcBp0Ff46oIP583qkf2OuXAFkNdA16nFUa
J97MPW8D6fCLIeFnyryG5P3qNxJP8JQXmCBJ3ee0fU931hNLVkp7HVDLUAaw52HI
xQJKP/KPpDJjJ3ORrPy9/aANGrUtfHrfAb1paC0pqpHgD0HX8jXJtERLIo65XkYX
FGMePUKWEu6tUngnceqEGsfkJwyxyFPsZoF67GrrJpTZ2tio+nru7QYlCW09TJHL
lT41n5vPRVsTrFSW/gw4QfZ5Wh5Oi4X216N+5C95boOmDTE+vdDFybwZOwJaEk03
ExSSwLOHMBcUylWbXGhDCHY/BpyF6EKz8LQWYJB2grJUwxyyNUe+aUH7pM8BEqog
esL1dTTvUqTuCTQlShu0CJFsn/2/wg9RU0Xu8JnE+MgQHMtZRpkBKiT4eMqXTl7h
1P6u81mRvyXpmiz3g1XD4mTYmukuRZ9SXHLksWMkem7FPupDRhlVowo3tzfeizdQ
CuAtmUjtuef6xO/tILyePAsnnF+T+U/0MYrqWNtHJIywU9MPjmRF5zkF9LpbFONJ
FNeISwoQ4WKfBfwp5My35Iioo52Sl8Qj6tSKZngPQybYoNc4XIeZqAitg14m4aFx
4RlYh7InmPjN90SmKVtE//3eUEkHXbTiy0mpUr0ZaeYnwek/A73+DHMvXk13absD
0SHPPsdcWURAIG8kvEZ7EC61isLDM6Z2DoxYZr4F2iky4gbZJsraa5t3mHn4IlWv
q7Tdmt3EQ/5Cxk2KFQq40ItJ8K2oM0mZTZvMBb9Sh0/2BXH/2TSrUn2AuYKf0oKy
siu3wE9PR5k1X28VkmPp1XSTx31KnUGLSmUzk6Fi6A7j09BAdnXXUX1+qCgZbcZj
a+HL2IrTxKa+zSOnN4UGQ47F7SJhuAcaxf+z+Ij0HGQL/VoHputm0ClHWmAuP1Nk
0hkhicEU4DU3vYbthTaqVitpsGYFcyhlNPVgP/fuihYGKREtJst/aRueFuqL5ITx
wvvV4iJcAT0Dqrshu+XQ+aQdvr7R3o+y7WP7/4+mDCT/3puKmckaUCEMOd2471RM
wJzM6StD2I80BlhmxC6zQ7JFMaryD/P4oXlUdB3rHtz8wpz12NO4mXrHftQ3FYDH
dnML+Jv5n73ZItgElqf9SzRgPAf2d2RvhFaHuhx/u5VnfgXh4h9wQ7ABGZncFwPQ
sptnxbeaOXs0W7/R/ExYXPL1KjhordnlWZlz7mIfZbRtgCRBcEg+Arr68MI+BBiD
PV3OVuThD7VenEtpEArzIGqspg6CXwZM2qEK4FchUFMS2F+g5XFcGzjSM7hdpYsv
49mMQPTvIopteS0UI2q4eO8GG+AJF9Fjyt7kbNg39W1J41hn85Scv6W9fB44rXYW
XcgW1Gr28iGF6nv0xNj0cS8QvPoo2vf2nAqGIDopOCtcPyOtwZJjma1SKsIz/+Ns
mwsABAeg4yubXcFz+RhalZZKdoTF4sCE3m8+bAistFCOz/5mZAnYWPFWu9ZCbF9X
iLhtaf/HLRgBn7h8JU4AHoU3EdDimd4zUxTvyV2aToCPsbBu3RNt0yb/UfPeu1eR
2uEuioi60umcVBMKgex5K96WSIUHmbUZwu47Mq7fzqmbO7VxCCE1YRvavqigw4OT
6Bxek6yxdaEwx8kLxY2u0e+j0D8Gas4gaj8KGgMSq0ph9vtq9TvwrV+CBcGGeWQ6
01cafTtAxSQ6wsRDZ5gsCLWnMXJWM4THC6RH7Px1/MzL/9G33+MSQvBfBPIfOazw
5zCOKEMOnTLbO2MsoFWSh6mW5Jp4oKXv40Vfzje6qlIO21+8nhSYyWWTfgMrUTi3
pY4a39y+2G/zh/+mLYnlDcn3ZZGHmOIlZbxJRJCyX8g2znLvijoo5ZYUYr3dM5mB
n4x8TxEtGdJM8EfwjQKs7DX+7rth+DT/KnjU1rVjRAcPsuCYTHyhYLBSlvlQKKaG
t+lWtJr7FzV4LDHyjrAvMN1vmheaIzGOnvjpkN4m+oaaDpOhIjguiXNlQWegfuxc
iXiOaKsxrmdPtMmfiTBbc2j3RzJWZG0oeHsol2sdu1WW+NLsfcG1Es/Yee6e7AaT
Nl1M0ZKZipuw5QeDgLtOdCQGbvauJa3jzlrQjdnM4KXrF4RV9ExJZqehtOkJssl1
O+4IJkAjon92PDvR/PoFpz4Lz76Wi5432TElH8UfbPKm8F2nk+DBQj0KmRdHCUfj
JwkNRwbNbStlLvT/yLEecuvrnVswoddd2l/rhfELp2Nz3j2Ub8ZLFly9AJlhAl2n
FqSMzb7P34yLe3M43i1gXE1Ss8Je871xKzEbP9WQRqfayuhGdZJNNEgDWORtYTfW
7a8ja3AcRj3kvX30fNgEFHxXxkhJIqm5ddW1071e22Wv2aDW215N8K4aIxuvC95y
7Ddo4ogbPYTvX72P0HNNCsFdwIKmep9rBMsxp3y3TVvdGL9iujonMsiCPRY7ISx1
JW7toZBI1MkmgvS0frJadifUGAf3EdZ/Fdk9QOXrx0fK2GqIjGc50CQuPVWZqvUf
E7VIeGbJMbmjJRLGIAs/5c4Z9vgOfwtp3+/3jNQW7DsRdtK3vJRYjBZJqTXMQ3Br
CvE+eaCHQOESVvIdyGVDrYjerpNWJy7c3ljAwjTo1p61YZnfq8/wP1DnbuP4LEHG
K+TqkHrCH2s6v5reFaB1KpYoIZvNtSkeFfIULrg/FrdiQ+DEzUAxOVtNr5eX8zOU
Y6eeyrm1wHQY4HR3ZS1Y9gyeO/APyvGsXJHCaiFW1oYQJtc+7CVJKQnbIx/rzZOr
lcdq/rUgeFXULm2j27ybeiMEEK9y1o17lNtd9bw1+2qFivOvDSZa84pnteI0IaKs
kxZhnVmOp84UCsIRYg+wfT42IZ7Mxabms0rQ6hpu/w6lWhdNsJUhYBXtTfOOXbyE
mSDUxsRDdYkl3oqqVpxLXUDu0thn3Fhz5MUVsIrx903WbQzAkwUiPGcvjID/2Pe/
cwm5VAHXFdC5QWBCUqZ6jaAYDm3RgDYPco09M4x2nPL2T101ZWGmcoAKkMfD6Tiu
qDYTgKuh75GF9N7zlQqPUfbdIa7oNHScfUelMSvlJ3NYXG1vqBm+0L+SKT485is3
RMG+v15sGeytBLnDaD58Lk4qHCCsnIHWsYP5hzDmA2l+NDRDVttyelGpVuci5Cik
P0Z/A1GwZHaVa+yVPjDR7GtopErvRw3yvp0d7ZIpymg5Qa6phqIszt+ic7yDO+yK
wJSVSos1b81xTBHnSorovO5oPgpQvg14nup2ETqU66px7B6k/3Xhm0YyXnj5z7Ne
XM+C/vlWMV2v5GVQuHp6KXkR7EfTp5V8C/kqM37krf2oCWoTIMW66sdDICgmZsfj
gL1VkKeWUIJr/YdzNpZAm7zNn/CxQ8GTE7vmY2SPcVQmgnmHwDVwEftD1zPWVeXc
j6lV0Kw/63BcIHQyt6367KKQOvaQvWocZ1ruFTEhkPz7pmpxMT0OOg1yfkBv84Ya
Eaw/XQZn5ImWiPrZmZstTRk5VHUUTOHWNaldl7bdiq5GmOmcLump8CcSgXwzlToN
guOscmTri9uJ86ZJPFdvSGv43PjEDGVeAl6rkHdR7OCCGtWXAzRrRno/0v819+af
dz5iot7q5YJxCCZGtwkz9akDJIYxz03vPjFN61RXuswil0RIjcqMi7dZ2HEH63ar
F5B3Y3jVgSo2Cghh7qY0zWdsrGsMoYvGmN5c4zPUFvXS8qyhQrf7YZ5Djl39iDQO
Xenm5zxOCdFW1rORqYzmytckhSbSosSIjNiJQqQs1Rb9EDjf7RVrLR1ywgqSKQ7d
J5iRfJtQJv5UQL4ozS03iyAphxnB5KP4fqrd5QVfxFGpqgDFpWyyWBxANrbpVeEi
m1As8J//T3uX8sVZ2yXfaFpDuFanAeTnFWl3H4lc2fc3HzBcfSFcV04ipiDfPcqd
HLO1RrFVS3JXbPH7BwUqF5Usb1PQdHv9wP65XzusrBPjA2hXgjQ5OLXb88Z+1nPm
u+Aj7er506VLMWzhPzqq+6LljqHcVl7FxwBmy6+fslTAX5IkHXrYs/TFPPNoKgab
tB+JOiQV3fcOV/wOTNwaKkzWQVctXDWMb5P+0e8uW1wJZebWm09XZlJ/dsd6krVN
A06N7dRTWd2vtJSof7R7L4TImDHT9PlP0ykqSSxXFS/S5ayTTWYnL9XqXlMvchSL
+OwTsH+y5fwLihqOvJV6dC5ZOB8wqoic0cCdJE2CEpUXpfRfi2HtHHAtj7p13snT
Xg6JorBeAxZDrnUxaduy5Zgw5gAjLSE7Xed75F/f/oycz7j5t/kkpoa2OxkIj+dl
BPBtpaPPef/whdL+Y7NJddmzbim8P32Dacpc5pQm0e3Og7mAa7levdBvtIEGCMHM
poBKnWhZjuv3M2U+pbJBw82ErCpHFx0r2ZliMc8Lunwfjj4TJjtwO3wWNoMQhi6d
sZXKTj88kndKPhejAR6hhy6DpknURzqwPedczRgExqN9xJtZPoeGSPJSDwvFnD00
2tHH2xvcjTnTbS+FOZT5RqrGLEfRzWp3CALH71HkOVMPeeASojY3jU7WfMyLWegi
7bCyCTcrkgCyepc6Vu9rNh+UvCNN5pWbA4r0HVaKU7nDGiuqPhG1QQO+4Yd82Hk0
cT7ndp/1x61f9IaQyMuqGUWpdmAEoUNE4jtEJ4g/YsqWLhKQzJ33+YWYXXadzLA/
K9ezglTgs1TwH0a3GL3Z7DxhO5rRWaHgSaXLj9nNE+fZz+ddccJoOT6+KMdws+76
fJiLHZWk8EtJi48CQfJG5DoAdSUBSca+PQBGBHcKoWgjsNlTiobRE4ox17Z20Crk
9LGN5zn0dI130pNt5qZ8U75Wne6jFmxu9So8/USIvDpfHqjFsRY/hJDZT2pIqCgU
/QIWR5vEI/+Sc9Too7HRQlUap/0L+qduXCKo/f0EGz+/D2cr5wd/ioro5GKsI3dO
YYdFoKGHgl1hCEf69lHLbjZd9Oadt39NhszkO3RvIRIBVMsf+UGaGR55+Tieh1Q9
+6Junp0HylbD14ki8pg+/L5n9cUnqplc5K4da4RddvvEl7Q8d7HdbUoB20Ra05Tr
GOi49dY3zaLHbLs4ATAWgjOgR3/qz8Gjk+YpkxutVeNnA28a41DhZknyfzhULr+q
/cLQqkSqgr/w8wmUsSKF23oaq407FoMUxx4GVNmsYpPja3eyDAnpMxBLkp3IAZso
uGwewW6gam0bhdOWr0wbz4pOM/QzFIQIDOJwsUTlI+zOdg+o+R/43rMTAvGpgvZ7
CejZ3mMpY+Oa55LETrcZiU7OF+aL21r6tjC0PXRGSE6z1nsNgsAeTexPVAduy7qb
vSbqcY0Qq6NoInxhkzoR/xWCO8z2uCU2mK650mt445/8DAq4fuK/21MHF25zTjP8
TDr2bFhoIZVVLs7j5cSnpFNCiglioGUjjr8DN5iGsYQSVrSOSW4J1RueAKqx9w4p
LV7giSGPw9J57aAl2jgvUl/tOan17b9lbegob5C2xajzJndWPhj7MBoit7PuI00k
otx+HSsUEwpMI4TEJRHEghNKW4frhb1VRKNTOV9T+4xafzmI1HYeyJ/qZs/37cZO
peKa/rgFy0PmGQ/OvMblq/bb2OPjw/N04U9mFqAxJGC4neEcA/rbGzxfYHm7zsRJ
LZwYSbmfnjxm6A0VjJvK5Vufo/xTKFE2nhi7+tqy0KwhlhJoOZJCmw3loVBWqhPB
KsYiaZxl+pwEDItTpEZk2MVsyU6W0lQ0AYBuk5vHPoPsqVXsQZIcWyht0ZBQzw59
jFKdt+g4/+poVOPWw5VFNsvXao/qaO65jvxkwbAiR3+SSzq4kZpmoADzXN7PK9V0
KTRCVfEaEmimQSI3KKKLiX8Os5w7VleU2yY5nzoANvSA7lJmqNEWNirqRqDWZonY
Y/RIQcoNGi6sigCkIlPZLVuMwgou0tJk1v3ProX3h1w6RzFICYFMn5K8EiYZFCZB
stiTyn45F1GEkVIobgQTuvEHS7HuxzNmoIaOe7P2M8kPPtGbe1FGAaqWIbN8EkUY
kZQle74fIqXg/7PoEIsz+CpHod1CeDFvnEGCpiqCqAsicQ0BECNzCVLIb/MZRI7p
/p4DBHC1APeKKgRjejGCWFlsFuQxk+3aPK+65TWbLkwN0oP7c04LsWFWJaOS9hyo
h/2qaPlu3oqUX9y22X3rjDgGNF0nTF1G792NQMxestbgQiS0qwAtMA2Oqwuchqtg
U01QqC+SP7HHTa0E+LKQSfAoJcnSSHFIQhVm9eDgvVodEWARHLoffhKM3+qqJpSX
GVOvCdJfv6uuddy/msR9XkIo9Gx+2gk2gBUZN5mVAgOP6AR17TjPI9MURiSR5D3u
j9jVLB8Mhzpb3UVfucrVWjhewgmDKenUEJPeIcwYV5s3Sj9WWkvbTrX2RkjnhDnq
yvjhAofhzp/mcom8vjZ5/7cEEWWfTLCeXZ/JmGXEu5FFYCehJnftN8JDb3da0YBm
uU06iwHQPwtQT1wHYAm7q3AOESro5Ow7bIIImwQRdhu/LeljNowVvVfotY++MN4/
iVBNXtEpfhp/cYeiAm0tBJnkh+1rBurQnVnpthdDgkrLnAu8XLUAq2Tth8HuzlVJ
rj++qPRMWYHOEO2JNB02tIMjoZC1Iwo11W3rPoAcDPigptJbqV5iq8Pbf2wTJXpK
A3SFiS51y1kvvWlAFyzVR/6TWyAaxFArj34u3FuOttAUi81Z2tyBaN0XHWOcpS9D
3oVIzJZ93wUEXjacRoBYPPBSl/KcOTLeZDJUAM9yrSecOTfZmqKme/JuZobnkOWl
pFvYMOVT/7AyHw3IcsexQaEVO52vfQh3sB2SRWvciEHi0IbnyyIDGr7l4Wh/OgO+
zyj8VIHPInOi461Mgx/yOmoM1l/5fqs3sFhrw3m6wnLJJs0u3CQ+OaP388QdTvny
hVYlteMwteY8geUE280mx7aWQ4aTzPV1uUS0NaEP1Gj0XwHASYrIB+3EzhXldPGG
Gkk0r3nxHoP6aeDGmcc4iaHkpMX9gpmJH+PjYt+nX0tEUirWDZ1ScMvJuPgdQLe6
x/KILI+25Av2cXsGYKyeE4wC/s/gglNHaKzZ3zS3w8zOP2d6G744NnZwh+kscTr4
WM5eOY+Q7LMjVoYafkuPnxICC8UeNKEqK03azdZlOPT+k4R69JuY7dICcG8wKIhp
2ppfJRo0hwA8A7awE90L+hkKsmNIIRLfbHNRD0e1CIVzjAu9hBEHyT5PYtRAXXcp
FqDhP9uCEA92P8HmioKjkV0m6KhDhnDdT3v7PfV8AYAxi0BRecvwti0zJdhsW30p
9jfht6jc/N7zsTlp9/Z38tKMkfkwK+C7dNEAcsDSAUpseYosR7+UC/PB0wa1JNCZ
dvp5rEwfBglfo1dkT09sEldWcudH10exNkb/JMVmRJ2uGYEdvZTLqkBxnhI566oi
LxNGp2gKWhZTnuI0cC1+u07/14JgIU2+fmZayYIMkoHxnA876AcDTG3b5uSllcRd
zaiQwwglT21gqifnehd48E4GtrMFGTKhH/2e8JvvpLzSGpINftvoejWtaztxZRSY
TM8qmemgIUA9bV8ptA3pvnLWvjpDPK0izjk15pSbO+Qs2ibJ1j2BJMYrPtBB423W
t3qNUyHfnBMdleZuEzU+ZwqRdAXbODFzvIprAlOmUz5381K/QD9HXl0sCZWqMX3B
HHuvUjE216vaidUmsGHkm8N3Xdwc9sd3xbzX6D5SbMqknD1CyYhyWi4JDRvPOWZ7
Br3CGXKn0KEGRjW4vr5DJvrvQaTTVrzkR7q+eMEic8ERyQbcsQHS4AYQm6e8tNqx
k6nZzn81RvrPodJgM5T5ClBJatag46M4IYBiu8kaKI6CjUGcQ3mCamw83G+fcilC
zCwIQDuNjCdUXQkDpGhXQiYDgwc74pp4F95hH1pNJAIwPnKNBnUV0SKinLgv8ZUA
P+hGzax9vBNrDNx/oMOfoTCY+SRjrLnmvPTGQ6uQZwMUFyhz9SL7F0SgHjTvHekp
eHmQt9Qbo+bfSOIqwmtO/66QvzxPjqly7+MOFMgD8qz77e/l0rPbSO2Y4WqeV+8G
vsEf3LVVKqo0y6tNla3MCC9eC8ydeX1JCrhxPZJjTcJFVUIaRdAnyMlmGDJbiQe9
ZcR5GXGfoK0qYl+Lv1Sv8HW7a+U3uX5Zh1fBF57U+8dw40Yxav5Kkck7fdF/5BRU
BvGUZXdRy0M1G1DMP4vbIN4mye201+MEDfmsgQH70EF5rs1PBeRglduKWS9EWDNH
Fs0xRJf/92+Db58kIyVCCgM0Jbiq1pkJchwb9TYO1pDY89kmdtv7laejnNcEgZnh
YKrhsIo02338k9GFt4InqU4PO1ikQDEmXps2Nhxw+5xC8hUmagIAjg56O4dA+KHT
6a7fsI0qbkuAKFQE4mq6iVQyMH39UAeai6QcLy/jf3EXXj+z34SbFlcLlGpBHqRa
QBl9Q+KC4ddFMZTlqm4iFvRVSTki7M9kxjdFHZVEjl+ZGjt9a5YIM/owacbG6mlB
clAlyx79x/p/lOOv7XMg0USOfjiRZq76iMB1+uF6JBXt3+Be//rJX+mNwrFoj+yJ
U2UWNlK9bSpJ8vEk345jk+O3zdd7WI0MDpZ6MSaJZmiyMz7MmaiSQfLrNjLR1tGI
xKXpMKXc8pLu1RVEQRJGsHS0xVbWIVWPljtMoKGnsuHOiGhIkusmX8j/rWTk33Un
vqclU4NkwDpbaT6pmbKGkbf8FyM9VcF+HPqF1a1Vk/y/309wHKQb+JkFACfWbhQy
bEL+LcrAmcAL5+47qMorHeN2PKP47KKUAbhVNyoAsB8W7y9sO4yZ4jxf6EmcAaT8
SFsV1KMOr/1KDl7prF2VTAPfKr5X9sVgD9M66CiUhINFV1kF+b54n92bcbz0kVV5
1eaPDU/vGTTGSLFM2+KC7ojTGz/qGMkZ0WvVHowGb6CDb0zfX5rxXsgUzyP14ES8
sFpR7xHT15mQkbOLNYiYo9Y+0AcU5yIJ6Vka8hRZ/Sv+ISL8y1r67km3crnz9mAm
aeWBIjPeVBYkh32KaNjSgqdOwlj4vIFaGlw5ILUPbqRG7IMrK66e/r7LJrpb2NeC
hVHauLO2uPcDKf35ghj8KzABKbd4cq5AoWFII3GghGRNUKWFMgpmd4oEWgQsjzxU
iOUTGL9WEpE+kxlL3vI/O0Dyo4IocfPxOMZuiw7/nRxCd9z1R+wy7GSHuxcqq+VB
/j9JUvkaUgHxNY6LRBxo5Fo0NTu59W41twxKPweyh4QDh16DTtNuoJFQFr8ikeJx
WYmSmFZIwEE9hSma/YMQMXsLaEJdjiPgYulFDGg2jDFKIHSbRyCCHw/QYccwkD99
to+k10CHiEdnMGvlgBRmyqDJpvjpidhagsDtfX9MtrbU8cFFMSfiBhgz+D06Hgt/
2bEVvQQZFDH3OwBMqlWNYAJpdPBTxivfD3Rnq/F9DO1eiCAcPZ/H5cs6kJl+cwYe
MB5UU7h41wadcZkDtrXjIhV/gotw8wOyWnnSyzDwxoVvXdR1AmZeSut9Sxf+o9uM
OUVf6mcveZlmhBoxhU0/3YTlwP2T+UFb3uxtN8GQRRgHmybML4IOqtMWbYhWZ1JG
hlaQyfBV0N0Dh9dh+FFlW2rzYcHbF8RYal/BVapmK4mrCu2WIZPZbHJ0WbJW4qcS
LqY278/liEA3+UhI4T5PzrkRxufMElFnlVGpWfGUqdXLtd73TfIZzpF0DXCw5TKr
tvKim60LHQ6hG5x44KLyj+BQ0yC1HA04X8R2A2WHk6iH7xmO9gVcPwqNo7ZbnABE
rSNGuuyvDdm2FyzHO73m/Utxn0OYFSjO9SZ6N1k7+ja5t9yk83vxZTu36pRKQbMg
CxTBlgx8JVtD0qfTxz8k7tQ6zsvV+qJvxRKZlh6klmT92lT1c0+w7ayEyTXrhuB1
rq2c3I3enS32jU+nWfLtpOVOpx6LxdHvM9WkcJm8c+xnAM93mX1csiZSRqXOLoWq
TepLwVpSTQ6ePh3rhvnoZ9a80Ag//cUdwGEOaFtklTibOkw+Ak7lDd98+2DwY2ym
CQavZCZasNwS6awSlrquXCYlUfA88Gv7IpAjpGRkGrCTAK860TN+8+cHXcSQbZ3N
RufPW/RpduBL+zpvqP4N/FVqBMO8OegU0dDirljgOF+R4zK+mEUtBigxnbqUm3lr
bN46LKDREdiQuvRnAhIS8dNsjKAlGy9bItoXKtg+aHE12kTBGbaO6JrApp9Uh+hk
VX4QfzwaxLz5xkCeHNpL7wNCDYGTV88La4X8JL78Jn3zC3kpvAkFcgNxNQOomHac
YWT6YpUbJOexISE0VDA9GHUww6wIsU0Yu0GZ0GLixxeadVUA4AC69ES/eNJNqQyk
XEZDy/Er+ypEMtrFUEcxNLPQgF/42NgiyREwNIQiwvP8LyIqeEToPgb22qIn/IwV
GFO3TRmwXYJQ1DCEMD9xV7o2ybhFNecFbxIRTY8GKsAj1MmpE6aJPUwJYqsegTii
bc/ztZECkRlu33KMlDSSi2EhjV/8Jjju06jkciDaAwKOv/9/byIQ2kbkGCGNKq4h
Jg3SX8/Z5p7jVC1E5g3/Nu/a9CVHE6B39iAo6AF/swOA708CwYYf007JOAZXDkAn
+qITGtAchFq7VyfgdCewayHxwnE+7mpL67Z2MRFb3mtqGZRxrirdL5Q4szGCAvdB
f7R2OFcJrWmkig1uXfegUYu80qWHaF2oSO7T/ZHXsyv2JaMOwtd3/VKogGQSHJbw
0L29JWh0Lr++ysVH2t6EYmT/mYM3PhPrtkWOXgFe0qPJJ1S5Cy3fwRcCeti/TWvY
e3ofmRZ1bHIzs4ryq2Smg/M1xEUkRPHqbK6FvOdajbPBDYHNXQ4u+PwHg32K+hIq
pY3pGIoHxPoK6HVyMS/xafYXogj8vQkj6hPHR3xJYse7iUTR3x2WCkVqbheigvO6
dwxdOG+FB3W4eOcdscFVED2M5L1gVCnqiNxC2SHUtRk0gHYhbLRz7dbjhBFsNsD+
bEmz/bSj8zygJrru4bL/XKINs/kucMXKgvzbq25nGx2tdiCIwN+0EdLsqXXQXJJM
S6rc9I1yBghvFqYRZLJpghJDPKyoGjm/Sr6q6fne0ujW4U6kjkPZLP9QTfajCsDl
ldUqBOV0FkbrTuYjW2Qv8Nj7x4fgWChbpwRZC26JN5mkMdqP3E6TUFZrmt452ypJ
Bu8grZGKUpbAchKJQ/ITcYuIRWKNnw1gu+diO0MYwtSAgd/6FCR6Iom65dyKH2X+
hYlEWLUkZp8fpLcXciLw1mWMe1Aio3WXw/223car5p436oHlD66VDFs7jXbehPSG
JTmvJ8ZRIP78WLHy1f5jAnE/7k1CIG1Y6QMbJmmtkOw9bo/RsTOcHerUUrP525mR
y+8OsAC+7xEMJWwIO66S2Px+QwQ38LnzI/dByB4C2hOdiQ6az/RBdqeTQ7uxAmgY
XexJz2EyiVc62qx4kjN77/Zl4XlWkiLxNxkFN4W8vvQbvyNnHYPYDXoxaclsMHVc
ui4HZKQhs1DtjMKhgjrvohdj5VVdr74QhTtULs6f4V6OEOdLFmvmqPCAY2UFhenY
3a694t/imClOVatJKZ+AJm6XVu/N99xB3Tzd+pqc0b2vWIKT96lztqBkPIVpbJks
TFaWe/hzHp+hzAGxLImfcgCNHcQYLSUSyyZ6tEgP4HUvB2PBNr3Rvu8/+5vLO4m7
Oup9PMAbYKiBLdK28YnRGI3z/AUFJeT6ast+Tx9WkvTmdjHslluOUlzkcXjhr6kb
oFbMAHU+YJ7mmRvW7tdPEje8SVpZQ2+yUGsGE8rOp0QRDy5ulMSJ6LdETKaz3nOc
Ya2svs1zf7lWXcn4lhAVRMHIjopdks+nykJBaorSO3sakWOb6ZPZngyPy0WD5vbk
v4nYGocQPMs8ajDnukiezRsgNT75DrQ437r9bG1mJMNseE8axQGkpUXLQ7U2OhzZ
b9gPjXX+nk03osfLcXbro5mCUo6y6o9VY9KXOUEuOffI2cLzp+XmMs5bOMZxGKLV
LrfF3s5uQM2vDzLKFvApu+gZv3zcQeVNmeHD+o4Q8qroposYjHmftmOo42yJwiy8
Pxrz/NzUxxSFza7Y4W32s46/XTiEYfuTiXAkHV7VTmunD70HFOFs+PPK1rpQDxfy
EFHM9BzehgRpAr5k0bmN1CMLoHpikckRcsFy+/vzuLvLQJ+TxpewZfemt8r6UZku
U9P3ryq3Vp7X/orBcYgfmDKV7qFS+hgibVq+b4VCqrvd5Lp0BuHnDj8ZVmFwofXk
tZOOS9kc/s9KobZ5ddZN01683mp8JOtTn9YVumFStA4Litc1jmHyDubSevBzaSws
haQ5G0zgEf2OY39R7emRXz10zuBFqabu2lgC53JcHWLJpVrkAWXx+dOwAEaNbc70
a66sUrNeMqBXWP/9xdeCP1ENZrGiVs0dUjGVOE3nR2Wn0VP5hMGhBueB4xGB12yT
ZhbEW/+LEnrHba7P6/whDSCHTaBthBK6a7/gC3nixaBnRlfCwMy3PdvRmkV+xWbg
FVnd504c3pXkXtcrJj7ALAb0P+T2ovkKAj0ImDY/LkV9fR4NDoROl9BDdt/kuO6U
mHNXhKytIMzPogblMwDWiwksNatw+92mTOrtSC93b7tZ7L18afvf5Vo4Oi8Do/I2
3LFy15AhEDWlOo4WnKLYvi3+65SrEoKtjow1s9q4KgKRyAQiC+eyp+kfJ/KXh453
5n9dXeClZ/AAz8lLTlUX3vlCHizeJU/hmp+6oPyP8pdD5zJor28/stchbdIyjgWD
No2Ddf4H87fZnVnvKRGKOmyMGen5X8FZJpnnJsHQGrxwru8HmtKF8p01U472gn5n
DPVBcILxfRdt3WqX1loS6ewqaKg5pd7R1jnGHxJcQ3Ho+JUvFFiON4LsM5RY6iSF
OBTPg3TQPwBEJ1XVPS6oM/51eevylg+zQaeP1cSTsPbwddAr/PSPScQsBkbDAm1O
fS9mKwSSLi4sQTNhgSGXGyiR9P3tlwsWs0ApHUMB4yACXV6SkUfE4AaJJsyDk6sm
HxYOkpO+5+kiD2aNypYBZulCwviJACrZ4mKjrfOSs7fotwM3aTDYHVRztKQEdtck
ZsppRSB1ZigGe2NL4U8jMMt/mVAl0y/dxgAmbL8/lTvRdq/VdEg4H3l7IMZ6C6xG
Egc7NP+TCRDLWrY6zIOzMY+oMa22uRZVE9Kjcnxkcm4HctYXYY9wsZvWKPRAoOV6
cQGdXLO9mkO/wFygVd/f4Fl5E4Ncz9oncnos8rQLMunT1MzdhjgFEZYvCyEjvk/Z
UOGI/awtRxDCyuoaPb0MpsF2y4iUiHE0xFYHF9j/JKPEMUngnyOmisaU1HMo+24Y
0bEzoKb2X/dRSpXZcXyNd40i/4kwn/Ij0vDtXn9vgImfRpkmwKI0l2WVK/gDO7PG
xJ54d/7AYOyERvfp/k+D1Bv8clAgsRH6R4QIWkQkz2UekLsdqyzN69mypmHBtcWP
5y4XYJmcrQQnCw9gWVu9cnWn/V0GoOwmS6Xn5OROHNNon49+/UstWs+jXspc8QzM
Oxx9kJCnXnJQOV3VTPgptMWwPmAAli9krFW/AZeS5N0AFkjJddz8JPNsS0v1aX7E
vXJ7r2V3OdMrsVks3fEpreBJ2NHdYSwuPKffFCJAQy1ro4DLH39u8oaTF8sD1PWb
k1bFbDfLCmv1Ro6R/twKskwvGF/EchoCEJqYbbmytS+Urz9CnGeX8+kvB1LbeQfX
UYbFsbcFaMhgH3Kmq11HSSg4urPBP8VboksKCC7Oim/tiWxWPqkpxsLO09h7CSOa
2Bu/hbcvHL95G8N2KNVXGt5NEjuqwcRWAwAWssbxPswWZ4FFnj1UiNwZYeZzBizc
V34XkooPYhZ/n7lexT2qI5uJ3j2JaP+HtFMRU4WDwrps0I3o8FTj4nA3ClnRSpyD
bes+mckGm3taAsmpLe4Dd8XYoB/+ePMcx4j4ynbTqvaMV9ArDG5plEnbLY+09zTC
t/yNAzNoJ799vowT5ixRWxZa/QObBz/iD4Gtb/ZApfcRXvZHzsAUWF9FLsOu//Ev
enlaZr3KPoS9aSp4c0gLTsHWuyFkPmgDKzwLBN+fddAVZnE5xDeisYHlNmLsCpeh
NGwBVzDrV61ImAoFuJFoNsGEa/F9Gfm5KUvN0BZXvsNtNw6gJYCz4k41GOr9xVqd
5aj8iUVFGWRLnj0SLNBLRSxMii+Z2oQc23zcowo8ZePKYHLSuNujaoluAV/v3qe6
f90+aqG8V9yQZ9HBcv9OC4VG0eZcf14I3wZiDH+dcTm8xxzDZRO/2o7S73wwxT51
tIoQpI4pxtha4SDPp02qHhCH0V3lOsanOf81cElDjm8ndEzN/q00J9THEcFgHPSX
6SUeeBcmIEh/e9pv2HjdVmOB/EohECbDphF8CCffwY1wXUfx79r9WlQ7+x+KgU8g
akXPtVzLgtW1w6QwfRDA5V4RocmqGDOdMJFEuyRDtnyjhh5GxmAD+4UGPTObUKXp
YXs5kVwTczIYtm5D8E6z4Udq69ukTLGxO+io0NX3trlzcDhKqa+g9oB1XUrg6MaO
wa3af52Z9puDomdpOobnVeV3xFVhCfkRvzZAVCqvS350yB/XgWqW0Vlt5hPXnFKo
95wzr5D9OPsKofDYGZp+1a8382QUacGhDQU12cKGkW0tSGcVPZ0FdA/o1kfounpo
Vk9hOl0cX48J/VaETOdi5sjvZtbKniKJ4346yS7FEF88LJZOw2mDHafxkG1GWJxV
+YtiveYBROwbO2uSi3mAK/XPy0lzN9zBHS5E6l6utTIEephKjM3a1aDjVEp8e1gY
VRoKRdl+pRofDeLYpo5OV7B6rEkUYltBuOCQrpccBN2bxnXhQPtwa4Tqnzu0N85t
HXkOQ1M43TO2np6wPaOV9X90vzsfhYiCXQVvegOiyueRTsZMKys7JvZLw5BGO1KC
J/R8P9u1XkRIyUdInqgbaj56FKO4yBeXY9RdvvAuGRC1vlAP6qWizXbSNVc7mEUS
VVdxioItdZJSC8OogDi3wbS76BiiiIU6TfY0jmcfrmeuA4hWp8VZOoc9XWkByueF
jRs4s7+RVdYD/M/OZUaTDDzeno3tEEIo8UT308WS1d184ju7TY3VMgb09t8l1fjz
Sp+f68IClDpVU1SrwHJqJbZ+Bqap3TXeylNP5n6T9FIKX/wqNELJhlG9aSqW3fVt
Qd9viRkZww6zqxJx9kwB/hXjkHvpKpw/xu+JdNnyKFAVtghtwf3/X49fFMRt2Htq
gICp/qpjR7ieukgzt7rshFXcWynnDnFxyFY6LMD6KZJhL8HKuBIR7uDCRMbI+rjo
9Fbdy1QctRzZJBouI1nE9q/nxAKCDqwlZ6q2FeHM6GqX7daz/zoxmlLOEjz6z72j
GwxI66TzyD+jv7nMT+K+Q4lwGyOzTHw6mUJekVG23VMBtScS8vs2On8ucuP268fS
3hQwvvHIgQRsm6uhFCWBY4eDuFEqgu6VMvXLDBeoAMZo9JkZDUyj8iq9iZP9PfGj
5KQmUoVQQ7J0UtdfKfwi+ahQvUaoel+jW8g+YpUGZv2W3jSAHrNZbX0CNSpt1/q2
Jxcp3DrN/oaC2U7vqkmhLwokiS6qkEYLng6Tzb3eIu8/pUVCYBjKMzduRU57u8X4
Ym3Cig6zg5inoepmUcBdG6Y1Ax3dx7eB0od2ma13ciYYFq82RJBlhuALmnIUriVN
hC5i4FA+ThyUOqseU7ebjucQG771yos7KuvUeP+UXeBLgOB8dMtSxgU1j6eurMy0
q9iFklxo+whzHuDtEYHG4VudCs4IJf+7njlor9u8+T7HaKsPysEAok829jSWs3X3
bx38EYUL+qK+aq3pYAN35D/iVsl6r/bWEUkp7JCYLqaeuT+Ihv/Zs2GSfvXadaIT
XStmoMXx2trCGcyYf7xEu7R2xLIKjx9/2AbAL2B6AtNm3D3Jqj0c2/WtUBZGdVal
UpuOJqerRXZYJufgrkzVAuStfG5FiV/gFLT4/26uUcY0tX4BBMShSL0SSESU9kah
hls5nGcF2GkWc+Ys/nK76tzjG1Jp9+fKLIbhxKMdoJSkOrGtZwWbxjNzN7n8JJfD
B2I1eF4VnV9SJZM8vJni0lMP2LtvZ45ggxz/mLHtJR+Zs5bBfsa31hTMoRGXYDho
WicUNV0VVyalEVrPqpCGVsJsW0nH1rLAL852X0Ik/5s+vHuMfJw+nzctmy/1J3Xr
hAiY8ng8cvuJc0GGtmdSpv8mTJJk111ZtaLlPhvY8WmE7qOuJX7tMAOeSmLaEt5M
aV5MtTuiB5mHx3i9/j8k4E7eTw3uDhxgnVDEc0H9S6rPNTyKhd/m3+Q/WH/hlhEX
6x0WmeGbm7J8KXvYh8gqxUGc+3u3+y4JYFKedtu+XaiePhlIcBZLIdMSCRwgc5Lu
zZXnjUdygFuK0RnTRpK1RxlUa60SNxHx1/r4XKQvqP28VCW62prCyK28WSQILpIa
1HgpBXdHttS4FBg/y41SJRmtvIgRwGXBoEvRV+gr0a5geSpuff+SmsfQ2MqOg9qh
uGdpoz1HikBKkMzAvhdHwKe6+N98zAcHHh6sbEhldRY0rgxtgNArDdzsLSlzH09X
WgtgzhZzr8EOwWrX7r/GrYaA26Eqe8HHlwXZdlRQ2ke+QaYMaUTqvC2RQjuzq2u5
1O8HbgJSDYTRECtPolOe4pQs+PtpAtkiuCwz8MvwXLsRDiKXQrRYZFzNSSW3Jbjb
9SsnOofXUfUAOwE1q9XLj1zO5GBUul+/FxtCIv8QCexBNNeVMQGB+KtjCM53tqLw
iJsmz0YSsJgoAzlJJx9os9+/tpZ2B3/cH+SABAMctUhx0qd0E+Lg4Nn1xLwRZ4FE
d6QEtlDvrfX8slULqEGIdDXgcn05GJciWhBEbDOU56h8d4pJBUhgc4UJv5YfTbFH
JarTb4Th+fSuGTaX48S7N+qtXO+BuVjtMlMoL4ht0rODoQJS2U+X0etyJIBLqbcg
QJ8eLRPyBNU1B+9YpHT2dYbQn1bKKK9IJS9U6ehYyOvzFf9Ta5zJSgzbJg24m/cg
pR0TJE8PAqnKZF9Kq3MMP+Etryrh99PTwY+8uyZbhhpFIBW2g/dsjScT1j8ilqQ6
yydJpSxS4KIhAhdMBYPEZA+x3SZF+NhoZbh0D1Hem7vDPUnpkXJMFflyzUpzF/Gu
HQG1MUklYJwRln9GLQoLwN8TlTKdlPI1KuhpXsWk7U/KiA709V0Hd3Rj7allfJhH
s57i+VBYjA6YXDh3pwcV/J19lEIixW3awncBlZeS82nfkePGb1aG3I46sGkj8NMa
FvNt7NCFoC0k91MRE8D1vpv9FMxW+IE34E670r3gS8v9Fy8w2CNRPJOH0Ulggyx+
0/GwKZ08IMkLesUdlgcu7HCugq9AN9vfBRuieI5kXH37KMLxfMB2LVkxEwcmH9Lv
7ZVJ0ID7nVIPbVXuhMc0Y+aN0kWxfDth4mWs9uhDddJwcPIlOFXljbCBo0rmpiSw
BlgwiW6nOeLN9EVNbUgMKuWXZB8ufGdCiPyOku6n5PmX4ksYc+TjmvQPOgCDWTRw
gQygi+tA0nEc/A9afinB80edxuaSINwPkuZNlT+YykyeDR07/5Qsp5isaKdzYL8K
RSv11fYaYPKzs4VPCaFjwVjNOdvY9w5osyweT68GD3lVSj7YMwN6zCioldFo5jSE
+lz1VtDk/J92lCsoiv8MHQpuVXDEslKt2kZyD2g3CvAtce6yEr5PFO2TL+ywdiPP
BcbS8f8RTgnE1QM70kaGmdnMh8cDbDBvLIuKQN3tcNX4ztnQUdGVCFzhobxn9USN
m9ashu/B0oVwELA2UphOlvVQuFyMW9Xt3Fgfnvux0zCv6h5+r38jDYuvIYUQHi3Y
y+KGwdN1Eo7u9Cnd+6ikj6gxEKahH1kwGDAzr9OhAcvx4wrCH+dKHhAs43iEv152
Sc1i61kT6Ap3t2nUpHwGs9CXPZ36vOiROpNmA5B9N+QxXVGJDp4fhPp026l8DAGo
OkpOo5aitCVXVAYiB1lMLFjtKMBfi9bO9sNz+7qYs7S/+46fWQFeu1SDCmIJLVkS
MTXFcP2EDCPjQRBB3NRDmcD5QtiZTukeavw4wDhHMeLPwLhgfkaXRaIzOHy5qS1X
jb3svvEzLjPFPPxMA7bQVLJGLw7H5X3nvW+5T6HyQh5PYPFg/jW0fF/xCk0UprJo
XxjzkgdKfPuhEYcWl4B55BzTW6kCDGjxxjDuLGUEzoNqQuj5yb9W3A/upIPyOWcm
AjTbScqOFG/1Fly57hNdMOfL09/T2O2oH2idz6W/FCBGcxS446EsLgjK17eu93SM
22GwRpwxIKvHYnECPfmm+7/AWrR2vFJt+xHkYHp7CwrYWMoaeOlYJ8CaruRT9rbn
OQbyJtuEHBgpyfFVn28NGCUPwuHS2AsxGfHFhau2SiUX9iaFBtY7YsTiqtcPW92r
JOPgjBsseuDbfOM514K4xwBY3Laxochps4hnDS55D+vau8yGEXXV5xoSQ+/GK305
ZuiRlVTPwOdbShK2/EGkVhjVi06/3oSIxCyUDmVbKi6w9j4WnPeWSoP7P57yRI35
cKh/msmZ6F71VEK6KudG4OPskLvLGzNb1AgcmWSavfz+26Nm1i/7CXdAyWggztbQ
EU6n3K+bpRqD/HP5b22IHwuxFKs2bHhByW6GDWC9xHwC7r1wWmRvD2MtCmsZQQlr
tdqEgmFnB+hkF5oViWMgJOrgUcnb29hM2uAyIJ8N6ED62Vhxf3k0gcftbGMTQK+B
UBjTTO/OVlD67c7t6jM9NkZlZ/18gAo8htaAX8EquCuBTqBmlVWHsXBn6WP8fD45
C07tqKQzaG7X67YPNaeBFkXpqouC+2aSxyiaWCh2KfibNON3eff41PmOGKxoKNqQ
YS0jMAkltVdLZbjAN+TRVH6Nd0MUOsGIMJ7AsVwwwJ6V3lRe5I9ZQ3PUio5D0Mvo
u4JJffwXakrBgqzE96f413yWTqdfGNMvGAPbARXGD2g+nRyt7j77v2CsBvTEI6Ug
GkKTbRZCDLDscM68LckdXuTff0QbaX7by4awDAI8mOOKk5wImTI6zHlz1SNkzJ0k
zfpy5MVIzDtmqagalClz/+gy2rY6TALtMDiIUI62sCzhy1/yhXgSOSXIj9c4qJkr
Uj5/B4etZ2xXeIkiHZ9e0j7F4skmUzIvQHJep9js9Z/8tdPnGMlOZeDwXSuBKOa/
mcp5v49aDibrtHdrzBYtfPay/4Gm31zzlBwlrGyNMH5vFUe0y1ECX7XboLYHsyLu
igVQ+JyVpUv4w5rE/f37SOwg9ARQuTbo1WsRqLXbmyo4EyjIFv4YEoGyPUH4MMYd
nYUNgaZNM8kwesbIhOs8mIXsS0CPhRc/Wi4Tdy4I7oHNgyk/IEkFeE1X6cJgXNvk
SriIIQbLTNEW4Hi2kJChTPC22QZ0ZB6Nqwzzi8H2z2oYCH5ljqFr79ld/U7RCgXJ
aDd3TEbhXKydTTyFDZm5aeJzZ4I97Y0Z4WRJkjhN34gOS5qJIRTFwbIlKeAOG5uF
kos6pGjYu8ilBUcwaQA4nFXdZn/9R33c0THm6LfuwBjqhj5825MOX2bslytULT6n
D4hMRLVUNDpc0z4da2A72gfxQtYNkgjN4/mTaC9vtSLgrlxw5CeIGFak0yYAV2ob
Up8R0uFOVjxRNbgp4E+h87KNeF7/xRIbdprwwHNeqt7FL8uG0Gtr6jmjUF90Kyul
jNRJdB3GXlQsh9ey1bfx2MKVMiQKBnCXqtdhwYJiR5WleUaUFQFOYOxS/xtapXaM
4TvVrGY+AHgQEYKqXdNpEjGG6Py8t6fJYceG02x/ewevwWWljHeanp/qfr0/r+uk
rgjJC6WpgeNtj303/jGiJViUIMvXIDnCj1jmcQxPSP7LngYJxMSlIwtUf9fZrvIS
rdK0fpmSGeH1fVptZMXeT9OlqJL5RV8rm29KgSzGqcnpyFr0ie43qbgaI/a5BK1F
ZYII12uX12FBacXEbunB+VgXJkWsB7C2Mm8YryMiKsQHmoltJKUmB8ouabT9xOg0
iJvpmnz6oRIDfu2qp5RxbFnStbqMlQfoHt3hNRDnf/2pF3Vfy4z1/csbw0S9+xjr
sZYmZhygYFYuUvYu/GWWOiB6dg6wo8n9NKgGFgR3JDTJzPQRxCJkZpJ1YEsq8kOo
Ivb1NIWEJZPlK9BMKQ1m1XDMWe8Q+smiL8j7OETM9PHUf+dkTUzR9pKxZzCEzyZX
32umgfJsAApmooBJvRhOY+oxbO+jBqCKjm4XuxpP+Ld/h0O4jMMdGJWcmNf1pSWs
8lGK+/Ys93pgnsqnH16WBw71GB6QuI1AeYtyu1RiEkdieEea/CLALInQA9/HJ51E
ezJXzZLcaAsS1ZAqmtwWafGdHvbThp2ZXvhJYeOgjUGKwSblsNijTwgQeFNT6uwV
BVlBkAbxAl+FDQeFrwssw20VdNRUYsQMPSEhV1YPWRSbgpTMbhX8gbMFSupV6wjc
NkYDB8gKkBglSsTBH4zR2+qizvE9c5uWCYGi0LldW+5pyMayuyd+eYnTG/e8IbzK
1n/sX0ITZKQWyAm6o/MUnLTkrYyMNkrjOzobImyJ/OUBNmnhH2FJzaVBIzwSzqxG
Lf4CCdSjBo40fbbt9FRBZzH81nkxZdOUeA63uUSGKVd53qlO+rRObqlWyo5OTWU+
PC3TtbT6aQiy0ya1U6ET+Gc9Fb1DJxjeCyXnBXtZPPClaOCh0tZqILJJqwb1B1OI
Z0ghUSPMy/l3d3Wi81fK6jFbARBmxmkbl+cbgla8cdD8D/Og40gdIPbcljroJrkn
IXPop2UZBptBsrhbmavd43QDhqxnW9IBoEtogpoPi9sRtoIiSd0HpDJeSb4tXFJl
5cXvS5cICdT7Y5aT4et/0b7ppXbIzum9iSsFtwEjqgrX+4vrJrjL98riYSS6elM/
T2cEsn1w2p2qjO5tzdF7h8qbZSBs3j9VY1aIzs/wDAlp1ycSt6QQsIPuB/sYM8Ap
SlPfP6ncF+dJ+VoQCwJlx7OkF7ZX7S7nzI9AKdtoI3oopYrMu58KXmNPESbIOpdW
ceethRSb6SQv289G5kOJOTw4aX3WwDDomf7FKvwM02hSIOxVXw0lOhdcy8Ox5xSv
k5SSUxcUqZ1AIY4ZFP4Hnb0eqzM5rD+TKWPubZjnC4pjXoXv8SM4fWNwi3CBVFCU
4HTRGgVHS3wfrDNAS2lsb8hjo7E6R9M1bcxqAINV9mG9HO0Q9e1Sz9lvXs4uFK+R
bmzb0TI7wvFmEKizmMloiIItXTc3IfxH+RRoo65rESGzXNTtB3GJu2ds9YaqKFiA
x1HQq6AUcMbWjAgt3ILsXjSN4xyzq1wZjL7NjX/zcTfI35hblPD2kBzsITXFk9uY
8/qos8gSniLfL/Zcy95W8i/L6X0NwjV9ruAiZ6wxuzzme2oCdRcZW1QCxd4GyZz4
F9L+ajh6zuPK2Yc9WjCnYixbV+fiFok0WvowjuF7lPy/X1MNlz4Hc1olrVE7p3zV
+fWcnu4pPi98ciyw49nbIdT35P2ZZKnB9RVodfsEu0f0dtf4aiauVDFGiilBwgWp
o2Z1IyrMNL+/bTXcHMWdsP5xnGC+XgE7xYNh4TOCFxURkhcKHtCq+8ZSRw9mwuwL
APSMOT8vojOWZkjW2LHMEACk8/vQA0ZGqi/eLVzGbEMwqir2l3qRXWFmMdDqQBAO
X667ubClSuPofvfxqHW1ql6198Slc1vt3O6OdxvaBjXNXkeHKDpLp2AzNT+gmQeU
KcRLuPstjt00KUJ2ewnNCn5E+LJui6d24W+L6CqbxeiH7vDY9mX+BXZS+DuLUtCe
g1TSy/kcY2w/mNkEPq1C65+zi55+ThFph+nQthD+4o9jWeshKD1gyb3TW0sA43MO
wHPjNA9LqiFZJ9kUwj83I46M5l5OIV+a5g+wCS5XvOvRRLtYoEdrIozZ905CYsvK
q1+VM3Oz1psfWib1WBnueh3Ob/IaoBdp7iQvfKeWthIlmvY6S9hRSHM/sJDU3v8b
KFxz/FGU0+5Cqu4dj6QoZ4TIXmFEWNhqI3MgiSgs4+vfkbbyrIAQQgJDSA8My0DS
Z+USiM42eZXEVuiwc+hoXb3xIK3zBOasy3OA+5voQ7YkrGJCX/8b8IUi/5IVjnke
pVkXhG0OiJj0LDXULUAmYLHyVjtcaeQ7iqcCP/krYnhDYsEBm42ic3tFJRti7Jsv
eRQ5kF/B4RAtPfIke43QLVmtvHYBtNVq/1RrRwNaIO1qPeH2ympJjU6gZPUJWrQd
vTgGl02AzvwkAt7gJZ9i4lfgnm4+WoebN1BE1dGQhc6hPhM3pBWCqgGNXKfp+IdG
3TuPTaVK6W+aMYelexoyM5UUj8NXe/qtriqtcAUdItgDxlFPAgsO4VOlGSAAlYXM
x9CzLbrubklKksMfJJcRhlaePA4MCMQj5QAxqhtgofLEwCjJsNnBlLyvHtASz3BY
xWwpL0vdmK2T7wLSvINgJzHXbAg9IVcB5yQiX1t72AVqSasINMt69Chnq3HC0iWi
SIjleUfbi+Mrbog+JEf6V+D5lX/zmwRZlowHM5L1D0HZkhc6eG0FsrEKQ9Gtoe3v
MrlrWNAuQd0qIQl2+z2Zv3fTgDv5nrIBgvHMOh8WGGqUJGfMFlyAt//bxoy0YNbk
w3STZLm1wKfEFTdjKWlsZJ+otz3lxi/Qoc+kVNHKcAgarlYMO//OA/djZxhm10vW
75oHVy9+W/5CQCAoveRA7LUJt/ToS8cBH6uVig7GwstCwk/NCl7hMXITOtX/tD33
DgA4QO8FIjNMZJDzBtrqRnmP1sNMYppCfn/DfAugJA7WzV3a8ugWUxCj9OrnaWDT
i2bOhSx8NcANpVUXBz/+TXB1u12KpiPuexJHwghIk8j9NmpbThY1Gi514XY7zz5D
l0FSWgKhTi2z5NmSyTUcUaFrNYzAfJbhmEjrGzazVaNtAgGGz4FZXVF+vSRnKMGQ
aJUvuWFgO6BaO1lBAvPq1V4SzvvBAYCsv78ZNjE0PZ9bLspyjSnS7o7LF+Ky/kO/
YxQKLWR0z5FM9K0y+Hdxn4USJOCr5CWWWOKwFrckR7FXe0Ez/xeBtgthH/1pK7bc
Q3MQnzjHArX/I1zRS+t3R8+mvkdQA11FdUlHkS2XdrXnb00HxKvnmJ6K+nLJWhti
5llklpBbCrtPu+PUmZ5a/fw/oNMtwznL7LddS4TKmB7++jOzrDIAdKHfK80+LqX1
uJyZrG/nWljP1C6PIRY0Jb5HmYza+NqIs3Mmds1mqSo8f/k9M4p4FXmVe+LjZLU5
+tRqPgQXkv+LVhrfiAgR+rNvxg2KEfDutKruT2va4RnCf53U55fL0sQsSPQt4q5J
WW7XVM9f0XhhM/wiBVXwENE4CAtJ9sCkPVyQkyyeVMTegegv0biDuKJYpgaErAvA
rfwQG1Mi65fYSMa5+LzS7nHuTc6uCo8mM1asxCZkl9DN+mEqQDBWLOJxo+XpmXmE
9HpL94Z1WKBWsyRtyeSlPM/Y2m3jWya+uILvYgUYDg14wlQGHW4lyvWrAgKVhisY
fCrZ0EAZ3SPg7HAO1UyXVJTPM+6TM8vNMYOpH1X346u2zxKfA/ngCsVB3fcvPzbO
07QjxMO8oOqsOGQIH6dcDiKfbMjwCcLEYNz+/Jid+BCNWz8HmaXbx7GmH4rRfjJh
XYvbQ8dZ74vuIxpFgm+5yki/Uf0Yo1A0s3FVBruzyPUIO5HrnW0Lo0aGoI+rw1jp
PyTHwX/ooOhxxtwuQvmLeSLMiJMchdOZm5D+frxrBUIFYhAj/uzlF2zzYHdefQoJ
dd7QCKqUiXPWxFak/AokVUfdYPxRSVdkUMS9FY1vgPjGBGbIABcRKGPZS6yOxe8C
vG70Re8j1nI54geSTP9E2MoKcrnsdMthjrUsZDyUFeWHle9FtxXbcFXbtVIyCCcS
buzc2aSsbj7W5tTtCeppJLY/OTkXVpDvQXGZMyjstPS1XXOjXy3EsFro/5XfWNig
tURxMxJbd/exGnhOznEWXzE8q6imeFc0zM/PDgFNe0hXXPhAuyWuEQ4eUB8KarP/
8vPS2VeGoxFtFpLDevHI57XFE6+35KKy8ieJ/arIeAy89wM/IGhWRp7NdsQbmN7U
9ivxbECmQiZDVNX7RgmVzfE2OTIUktztrYTA2p7iWktPU4yQnDzWlNSmeqPmZNc1
4YcCBGQVEAwir3qCwTGT+p/DTxHLl+js9JWm2DI9LSSydky2oLFxY7UmkCNwQIXi
bce2WMu9yWHY9rnvPhgmHIaZ9hy4x4MUV78Ye1YrpjIZA0Nf4beoEs7KLURSLU+B
bAzSCiSR7q5ztNn95dygGV2LwEjZZGixBVrLsIqmZR3BT4q/zouYXBKu7bnHKj2I
JqW/1miOX2/owWTt4iV5JWqTb6yYQQroRCW3Tnujk01/BbMlIYI68YIqnqoRlAx9
WNEXJoY0ymspvK0FtS+Rkj6NUBwNpaewPlTVrueMRE16xzpsj1fVgcpHlE3/1QYI
HL66qA12rDH0FJZla4ExJpFrHzbcrLMG2v/CpaXcEMzFNEixquhJKDQW1/LAvztp
1JiGZ9JTSR2OZT6RH5mGPYAGKNgR0q0T6Swm3aLrzWK2k98UeHcecw6DId9rqJQD
WssmyX6gXR5DR+aiTZrK7j5KQqjCrJOYmWxYeQvrOHU+iY4dqSiAyz1BpiUlSXhk
tGv8HZCT6DY5T9efIh3Te/KFLxqMR13ia3F0JjbB0CbP/1XDV8B2WwziMKkEKUDh
SAD0WElzNAfIU5jMnQ0a0LPBcZNL23HXyzHSk7fwClH/oezFX2ophPj45Pz/9+JC
W4Asvn/yXlEeDCUMVl21xuvoJDlTFyCNi0wPVTRzF6/IVhH30USdtSyjj9q07bNL
oIT3/TidO+DwQgKTqcTO0aBcZ3uEZo8rIJ91zRU7QEjRt1BMQ1oW7SPNv9u30cbG
NVMjVrHUzsxo51PEa7hTb0YufvkSS7ys7KwG5ogVDWAvbrbgyBDDvUkhgdvQreJS
WAZ2Id1OvMeeIwwwdzv60ViEfyHnfMpLvop+xAC1J0M2LeVpqjTG/KWOFzNwttWu
o4gfpqU4AQkII5rVlfN/sfNRsY7tOkA/3kSSd6b8WewbXJsNnYWx3UjqDvirXc6C
GB2jMga85S3/ELF1Elfk4Ackrzke14Unh1kC0NIydNbH0A7gOVs9cKjSj+kVy3WE
W8+OHSXTCtYDX39tzZoc2y11rsycHrYyOkp9anz+S3ocHMxZ4rptv0Qupf0brQnJ
95BeixFsqXmaxQ/9SIjM10zV+WxKznSi21CbcSs8+o+OOaJ+07JVxKjD6+rjBtVw
jurVNGXcYk333nZJOWrUNqU0RBmqA9D7vsUiw0577ybQpOFc++iFiC1aJyc53dkB
U0JyfpYxjyoG5wXPjMWDgJrbTJyNrE3X0mFDek8hM+RU4z6Sfb3X3R+J+UVcpGc3
wOEJhV/bTIwxyS8Sn0TORzbfPiuyDpHg2NATIuLX54JsICQkCp8HwYWTK1k3UQN3
WBI6DtiZADzm7a4c0Dy8t/aKcLOEd6p2SoknLqNcp6lVbZRshYXKv4k596cxJIow
/pu2N5NzB4RiU1+bYoG4jKyJOvHUhMwmazZoJj7ub4Mj4FcZFk4jhkIDGW1MHYD8
KBwYZ6EBs689VWiMa8p/P9gvrxSDxaEnZDPSsz5tvdwpQSY7uK6AfeAO1U1EZnoL
GdDyYlvaAlt6OK71Nbpu2FZeSiyk8+a0i6rL2JY9Mc8Cfiv5Znbv+bP6zXLFyqaN
XSuEfc5ANQJIOgzPwiZz/KP+AeQMLcLXT0MxtsPWNRrxyUZE9Nhdbg7RPtL3Zn6B
AKxYKgJQZ+SK7piBEu/78SDPWpLe7yl7GlABSUBP7nXNWEDEKhKFlj4RDNjQ/7WZ
DVrMBOdn1ycnZwkfrO+aY+0hL1MZSSukHIn9keGLAN3lHg++l/Oexb7Mr11fICbN
yM8Clrl0+tXMUcIrd6+udLvKzdArh3EWAtMkfqHVHlPfg8S/5e5TNfAO5lRDXG+w
K2hcvL1JGtm5LV0PBi2o+JxdyKa/+EN+z917ycoPE/Fn9CdGOueLrgYZjdfm5DBk
6wlTLQtlTeCI0Wmzfr04a0o7n/8GacI+HrrxY9noO/Lvfj3iQrQW9XJaS+F8dYfQ
MWYj4JWZ3S/QaLxWs7q3o1GnRDx9KTx9WmYhyIEumj3xs+0f1nQtuH//laj8vZzu
G0e/kZQW32wjXzD/JAKkIwjE1Wjxtt3txPtPeXNQzaTro3Mxvf5yuvHnjnxgUkF7
xKHy7LHbLMjRn5GOPQsJNw1DlDWJIn+7Dq4ZWPW18rh8r3VNfgb3Bgd+9HWpY5Ei
pXC0OfETFIkgYNRe3TRdPfkWTKERZFq5NApDj3BCTJ4la8rfGTR7VlFORKyzgWR6
eYdQessoHBiPXLoD8RrnJp4ZpoLmtk/gRe4aD08eyRSh506XZiOwY9JccXd76AwW
LxMQEer/1o/vvMYThe7NZjrxHwbxta99pmW5VXt50b4MhTm1/qTXxpBqOnlEuk/v
BVIdbCF3mX/jhstDGHtTg8G/SrjUoI8jr6rq18v9E2f8fPyoLYMhUhn8+6IK0DIY
3A1L1NVioeun51dd0emrCh41lGXILa8VxtCubrwK/PyfUfcTazyunPKmdytg+IU9
Rk7nHmWcsyjkjlzLnhxjDytPek8Z8g1xuyXnTS7dhNR1f2Zqn9f9yaGTwh2coK6Y
MKXABOdnoaphyAmSsNkgYBNMY3daUWkRB8FurF6bw3Pmh9AbDyPXJBWXk7pYqW1G
rV6X3Pc5Ij5ocaUYA33KsOEha67iltdSqkbO/7bBNm8lRorbl+5vVqzz8u1hy7qA
AnL0oLuOtN0eM6iB00X1oZo0jIMZoL5mkEuDllpKEaSPASa85R5d1vr6Nxm2sl/Q
ceKzap6tHLz2nPn6ZCjVCdTRhDgw11NTtNaCra6Khatjy99l4IcUbfqzI23J+Z50
YUrkM3uKojCZoAL6EpKIwD1iraTAWscUy3dVUXIFbYEGm+EBHhqGZUzi+TTq3AM0
n7VIlDpVWsYw+qYY766updonbSddXwRV4RLA/cMCVNxc/N6Wi3xL9cjOwxOU543z
9N5S0St7CV1UPna2CwobH5n1uooT5RXTZLOX9ITiZiNuoPZ82yO8nPReCZbFGbwq
AQNSj4zZkPNyk+AHFOFnK0weNiDVTJvsi7I97ocWqHzJjridaF3Jx/UzbkGgR+BS
juk6k7xZXj4BbdOuj4IDRGS3hnZVj3voBuvgmUVy8Q+MTNOmSNkwwNb61jiHZC2E
Jcfa9quPtY8i96QCh4TBhqLQscpw5XLuR1MeMtDxp79NhFlXT0dK1lRdhKVUaUjb
CAPZmd5jsG3G1+jiQ2bW5o/grJsxXDOo44P94QN/mDTgTYwkxYxOQkU9qO/E1+BJ
LZupYoJWoMHsHR8vHdY9C+fGh7TSl+ydEdKpPYs59ZNJV7UsRToebuU2lKY14tUS
cm+imML/Xpy/NKfp6uPuofQznJLqL2j1Xd2I0q7jgf0WhJlHc0VUxEEgDq/7phPZ
uKh6BdbZO8VdVZ0060R5g4Lo53kMqajozTab+PW1MzixV3xpAje65/n0kniv0QG3
GZl1n2+sis1nQJyw91GTnheob2aXdv8YVfDUcGmng6JJhaXYX8qr8kGUhKhn/s+b
g+pj9vOQhTILU04U1TfxrKaTzE7IwZsiiAwubXni09rAPL6VjqKmdz4K28QX10IX
xz6JQKqz61R7HmlgfzfHvSSKkrJ+QrD5DcBarH/aZE3C3bjqlKE0C2MXKa5e/csi
CqeVwKyX0WvfVJI2pMv0AcNZYjhgQpjZj+5y7ENdgOZHi6mvluqpMYqwTUgYoFgN
fk+6hKIp+f6AGe7CZ91zgfMIShDgJGlzq6GUUHCJ1u/Y4tXy9lDnUTxYZyBnLKdh
oqUOxxNMlPdOUco00Znhl9aQi+5J83dcUr5Nrtq4wwFa+EdKN5UtqzWBkIqWJVAH
1eIkpa7hHOlFwTdMo3wgVfvn515SjfQULZwLOd6Z40CmJOTHFEUxI1NO2WL8zVL3
oVkx68k6o1zVIwjgnU7VejX84XBcvsXBF5Ux/IIp6hii9JxLIYT8PW1GsVpzSDm9
3ARrBL2HDiUMtO0ZaB8BUYKjOKfKsfeNH2QV6UtojonqXePoQEsWWOLUChndogYJ
aQ0ivB8AGZ0ZzyH5ZGSgJTuEv6XlCzi2VE2TZDlF4wQa3lmhMAhLgG5aOEVc0kYb
8HFvEKmt4DSIIcXkSTWMQla13vOnKX4Drsc/vYLoZwGollrhpvUV50pC/gVc7M7g
FxRmpXrZcsHPhrwyAIrZwcvNmm/rJOsfj5PJiCcRsTdGbyFyazShzl+iMhh7713c
/CBE7LYYnl//WVvXvGSJUlPb9IMV1g90SEezjqxewWDpl7tpF4B/giSJbsoaWYmh
Da16giYy3MmZiQXl9ojOReLpUV8EdX/Y0j7g6qzZ/1hl8YoUReepqhv58VvKBw5g
AMMxPsTr78T0Sq8oYYKsRgJD7Q2QGtjR2pJMNLbsd1KFhaYKVFw0NwjadKDfEPU8
PHUSR8+TA6/SsQvLieD2ZuOnWtqcJO8/yFGt/fSFzgHyMiVZHpkzaZMvJjHIQ6cN
X9bh49mtFuoDt0viYKSvEet21BTSqWt+X4iQTN4OnGHTl+rR/VNdQc+H3YlCYes8
hHaljFsiBTmcQ13Y634i/58vKih50hvH0eukuY4FAR1eIVQ75W2r9zoRyk65QlN6
sZwURFc10SxaRng31gzzXk96raHDLTvbjtLtGsaxCkYZb7+r94OqpwGbWAiH4f8B
qhcVrmfjasnSMTlb5MPrQ/xiflYGExGDwYEB588GgsJJGO1CdtEDPF3lqzQr01Uj
MQGR7uExHuYcIVS38ITW0g/mX88pD2NBWkSlyvhnCphES97P2iZh24gc6wHac2zj
xu5AujCvXMDQl7I43tcCWXhd1mx1bunJQXcFn6k0uaiLZwZf+WPpsG6qwUzXFjc7
KBISiRhN+o5Jo67SjC2BS3fSWuIIVNRm8/ZPLX/coypqIeEOu4xLSqIZHCkbwN7Q
0vfK+aaDZi2wlJ8nOPLR4Fb6BtW2V/dS+j+Npb5n2GH8Z8jwj7u42CwwmUcDM6bs
vOw7PyHILEi9z7crAEBKV1tfEoPCBkOXBa5vPMuYo7O/xBZWKpS2O58zJTtNuSyr
8QpzrRIxvYn3YShE/32e77e5jnBQN9/dB6Gj7E5egVbrGSKqnOpp5PiNJ5dPJi7e
CNYIr5dHVi1Bm7Bjt2qs6lzcu7amUc9hfxVrYJdppYq8GHlhWr8Oy2Jihw8/krXI
TMPgL9pbM40O1GGp6oKxVnlE3YWBJjTJVVCQ/LKsfknq3XI+kNkF6ZB372ExB/0T
FauT+Scu4XAqOICxFbs7kWnmMYXuUR6aTE5lzvqVGCdQqKtJlKOC9McbxCQBUcSq
KAVxJAwI2F5a8EqkQBMX7OLJgKO0aKHFZXJGoC16SAt4aH6N8tVkQD03upFrJPad
78D8KoRpmjI85gOFwaBOqaxwjY+IWjTj0sq0rhBCNIQvqUzcNKIIApUAz/WX3GCs
n4myxiLxZNBwXPCU8S0GnRL8GSwQeLSwoeSMVdxR7eIuePDYlQdtJjxrxMtxcP0c
4dByeStLVb05jOQjt+UMjoRU9MdTBmgLjnhWIqxOA76SdMdoLcnHobCo6xTYla/x
357Gg/PWKU9pq/Z74LS6g3ad3m2ta02fojxxHl8w3veul24Il874iL+LBHdDfCao
qTvSkoPTZEZG13JE96fOC+ht46zvp4EhdFaymUN18zwENEASNrItbLBmcZJn9JM+
ztjbj26i9dXQM4lqxkdcYc/mABF+SdmRCkm3nAedCT6gwPyt4XWnGimuKgXmjavf
OPjpTk1cxez9rCtokZymMaMpuDTDuEmbZg9ocwCtrzfTl3ONe8kuPmFqpwmjbQk4
bG3V9DyicgCIJa0hXE2k7u98lwNfo99mdzlFIo4Zoc98am4Fng0Fmhioq1DIPO9A
tX4Yhzo9lbqfZtVnXCr9cVA53PR9HZHUfc1b4qpcZ1tVJ2g5P1xTtF/stB2ISQn2
SPFJAApSSB1G4HwGJKI/neceYo5wLg7Risdo6eFFmdseqMeN1CRdVQm5pNgpec1R
hEFmZEi9QNEJK2rqlZME4LPrd1gzvRpGbNFiv/MLv4MHJXp5dKaiN1lJ4TILGOuM
g5o3KOVLZsO5fNZukNdpet0QuzMd+3kncw15z87S/QNMGRjDfq3ETemuvWPPTX6u
yAgCTh2Q/O2LEj5leFvfwYc5tVzZjNj4/KlTHb/uw9xtPIMvyVNlYH7i5StAJB75
se1Bd7wPCdfY/Zuu+FF4AshUFtSfUJe3PkCQcRq4Sopedb2M8lfoZBU8hgDT+wD8
rOCxutcKYXK31YH4Uxjq3pPOnkhYtdwke/l0eKyJMpJP+QbMfcRfmDDth/UwZ+/j
Q/6H3A6TKMDNsDdiSehK4Tjwc09cDZ0Fp3ZL62fkqP7PWBmjmSnw9B82bqvdOYrS
U9NxSy0FT58J1uN0FWiLT+xcCCpYz2qgI/dhw0axGIpEDclL9LDm2xXWOj4viDfv
gE4ECSJ+KLrmcKxBAmY75i6A8o2k4Uis/i1ZxFVXaBVDLd2nH5YJK0/aH3oi+3V8
6XlIeQ8Wdkh3+512sq5b3ML6AuJl/Y2CIcuFQ4QeR71LA4yQ22s1p1fZY5FiBstS
qKDzA6Uq+TlL5+cBMiqLg/17rnrH0GJjNLQqDdHxF72wIqJvLxCvvhf1lQnx1j2C
Af2knFKf5V+ks0uTbWpI4kV/rwsiPb194zTlqSdRpmBY+OgQPOaxtKKamyW/8iE7
wqGnAu+XbimZ8tmOGRzyyygu6p/zebNTRFTU5hv3WUz3JbmvY5Atprb5Wv7feMET
g+dCfj3ZjcvzJzNqXKqlVe2h1qf5mpE8OhrQTT34DaNDKj77SsVIjdZrv7y5bMhB
LxVMNAh4+z8aZmlX983EzVX1UrASxMujNDxAhUzA6Lg8xJgUK55I8chzGsC6xA6q
69PXTCu0AghinDaXrt2H6/7JRh9YhG3pKKywC+98dbpzMuYFzyPg8xdXplVW2nMo
UXIvotLz6DBa5+XpZZ7G/X1VNpKp8FRezmiGOQ3+xYkW/lPZ6p3I1k3fAn4/t5C6
VjW8VZXYX7UAHTWxAtTUuxdBfpPIbtGybKDpNF+50iNTN8NS3LoZ9d4jPF3NG5mT
I9EULDYdGFwOoAHWEwgUXGnOQR4ozHHO/mkMWejxZF3/iYHP6OFXjfwUHzJnJR/w
z4DaPX4SLI0bJVsNZcc0iWw6aERDRBsixkInbASj0v83bPBqbmNgJkM4IZXFU4ML
fT8ljePkQ13nIBI8NhX6muLKQVhdhnTbk/AdHbshS8jHshQia/4vUYkaS2YV70Tj
QSk34u5Ge8cQGz8ymKwz+BVwnFGBD6tHi6q5fPhVHjtHH7cH1U803gJQ3vJ6Up9n
NJPdjUHkqvZus+0JZ3TRRDdLetTTjH+6pmks09e6QJt3NN/QELQ1CtJN/YuatKyn
OPWMdKGz4iIYU49O8DqXPEwFUtK+F8LMvvU19Ji+xJYJLcx/zF8Q6IgIZqkvSQuo
5TPD+jTK3wRM9WUvPOS0bM5/Ny+XKG8bIZUBoSz4C7pqyBBBXIArnGZv3y2XhZS6
11UskwDHojXEaW+5Lyq4C8RrjBaJzPx44F0b9iWCBcm+MUpF2TAoexxzeD9exa1Q
Hl6u+pJGDqdbieUldfqy9WQ9Eq9DBZisXokUzAec3k+ohYrET/bjGWW3gmEbdv5C
QZBr9p3uPGOCelDre6akMnPtWWEsqPS1jc0k5f6HJW1BwNvSwUPfYyA0IPCmgtxH
ZkwlVITIPQU7m5CuG02fToZtaXbHEVKerx+9HvUY03AJZA2BfUlyUSwVqovaBD9l
UqBBGDC79/0Azd2eQ2436APc3qjZvv00uqnKvNxi/ENWcxpCobZq/EJ/D+EhQUtY
BL4szC06nxlkBX9bNR4yq3ZEs2YpPeNK0kuU4lteERnvrrI4o/2dEXXSsoK1owcJ
NUOMfBCGZnfvsRKGFTZMnu6DhpdmNe0JwnmcIYv+D8qI30/pGaGq3Kr0AwiwX39b
PfEK8IBV+xmb+YQIzz+DjE8xc3SH/SjvLVjw4XRQaVVEG0SAra1uc4dwHJIBjU9l
cHX/LeN5IzxL+w4KnX/AAefMe7iMnxRlPbgNnvcIq51BIdOQ8CHPb5j57M6op++z
O72iGYGcj9gd4NBRc36J1USoBCWBvzrm7JpxrqeUpHEcu/WOd9US68DalkuaISvS
2byQMHPdLsVRSHYJA6bG49aaoj1xOqsxpK1iGiS8GJ2Qgm7PFV4jo/ZxU7eqwvtv
hQNbpm4pzO1b/XmVad5Hjcv6E2mbzARqDNP4COw9ZWFYSiG5YmcXAvh7FCfVWXc7
Rm/8NPR+82Ky919G+nJBEoH0b1tlNL2Uc1yDPALSiV5k3ktkG1CezGHfvZhawAAI
QATS32eoWLrEoj1yuzfTw5m1/j1qmmWaX4J2j2DnNRlCA8tjKoCRLZmXiRZ4jd7r
ZY/Y7xfkcaJ87DeD2x6IMqYSh4sIWQPt2HzFzWCEgrJwJSKDohgNqHed1LXgtTuK
SnZ1ZmwBNNQDYNH2pWUS2s4DQVt2uSks43ON4q1FEd/WA4OYvl7TrzoD0A5Rekc3
V9Wu7JaVys4YyHsrFAgCvf0n6Wy5O0LVYLjDMlYj615wskRVHikJaAGLQep2nPz9
f4NiZv1GqvZ9erTCDmIQIWQuyTvRAz6Rf8y6Z1QurLZM6qbRkxa0Iw8SZQMxiUvp
bXRwu/EJKg148sSBY/bRSQTld+E4DbVj9Ot1v83d53CwQwjkFhPwZ4EPT9Wa0J1X
i9XLvl5ntJ1bMYdKddC9muFsuU12Oo7iFjg4Xs/xw8i115mLtiUZT+fmQRxINBo0
xk1SFVTKtVPFFLPeHY0nh0cvf6uizDFYOQk6JtXEQzLy7WV7pDxIIea/JMb9Iz7P
WwsGynIARt8P51FBJP4c8Y9z5HSiZ6v/aGirkQaaF+iMF9zRaycYPeasw+QJfQ//
tPnD7pT4qfcnsPcrd47icriCHk/rb3P9EmWrh1zLO1JqUGwOj5JEUz0/t9wIa83Q
DQ1JUX5p0w7zbreM6d7L73LMsYQmEzAnNZdGTT9wPjMmKYffvgJz1SeenZupKPnu
y3iAtjcrCFx6OnLiI1eAu2lT7hs8Z5jY54Xlb72FtIr6TcFXkQif6UM41RmXyr5h
rE9tB5qrlVB0MZo4gv2DqtIKLJFMKMcP3PuByyZkyx5rRUvWlrHboj2NCUphlq9C
K3SwIHWZ4AsXMIUysVa/PkEI3dCgwmupDasF/g8CEGQaUL6hYsVYZf0temgUNIu/
DGMl1LLOufCBdmmaBKMY456ig131jkC44QvSKqQhXAWGPTpQy95fuBRlV4smdE8W
Gp843M64ubyN9pl+L5PB+9HZ0fnH+Rt+KDDX5StMRuhr/blbFPIv/2d8dRoOstDE
upv3LWFavTcQk50miu2Y0R7ltf0R8sPZuxf2WzBo3hWTKSFU/d89hwqFxlgd7D1E
KNrlAh+0PZE7bDAoT5vEbx3BmDL2Bmp4FDdHvLmbM8x3GSHKMmkK2iiEkuLa1AWS
mIHN9RfrVBk7B2WkQLalXddd7QuMPSamXj9ueNgYyLHazcl7hsGxcZtF+plo7oLs
oqcCgAzt6fo5MuATD9Uh0vIAsIbzd/z7+wHMpZkfb4QDZYCYlOkpRWGvsTxProSE
4hFXEU8LeqlN5rG4YMWVBj9k8SXoylG6Cp2ru/8sZKs93R3HC8OQfybi09C2MSpH
GT0kyu/8Nz1OAF8TKlRlpoWyiQ/VxIYmdNebh2uOwc0J9QxLZ8wzqg9yLRBbaxGH
PZI2hP9oMI9JabNJ56RoT7vDeUdz1Ra0ILyuvwnAjnLOlHbiMCtEZedtdSyIm3ru
lFXnryEUKcNlPvQNEPleUmDphjioNzadYAQxpzuK4Cy+Yz9UstsoaRVOFxIVWMhC
UzDPJsSBMO1cw4cxr6EcXYaH6So+U3OuQ42YDj/aOTfui/L45XP1Y/An91M+d9FA
WLej6y/z9KBd3fJUFVLexjk7aH/1Nhh2XOz/vPMy+Fbu1KHbkEwL+oHrt4yHKHFb
N2BFLWyiRBaLa0YW+7Yah1Q2NGvuCUR8zyOYvl4wCFcj3noUJoqvBAdFV5xRlY7m
6mrOF6h6JiCn7L/HG/A2ApR5lhiQ89LthAA26zDrHDQumXsTpCcENMLHFxgPlzi7
Ky8DORL4Y4ftwrevmzDXViLNe5TKkZidusCcpmEH0+3SpOGKOihmNfSFpfWxYQZ5
uuGAC0ORi6ntCwwrcTtFqcsulN2SkPQntH3sNFlueskavwgIBjxhw1RgG5byrGvR
fuFEVUhjzRz8nTBw4HXjAzXpiKJvrT87Q2iWeKm09fX4rnS3qiGDondpgieJGCu5
NmE9H2kMUmpL+XL4+e6k8oyPV3NXkxw5dueXya8MiR+Y/+ujcuK7M55JRRiGhq/T
bHXTC4GeZElc7ch2FaFmffB0k6p5S51wN8cSyaQ/RpKi+uvRa8tu2x/WrhG/9oqG
TNGkuwW66fxIu5qiXSTCorEf+as+CMaIweisZRA0dppGHXB6q6bfQJCnHJaxPymB
D7N0n/kmbAwPoFi+A5Pp+A375ilj/+7QxSsmBfn0Q8qusH3SUfQyLNedWsTchVpn
VMXD228ZAYp46tkWkO9B0JgRsXZNJtOmDk3boekSbUjxfJby6SDn/Msg03W1NQ+B
YsnEiJNLFIQ78mVaybD/d468Z0EHORhb6t9ZSSB3880JOee0o2J2DeqLn2BRjtdN
mYNuzhhKoB07Rmot/9AkLw7sIG8SrZ8soSAfawnQ2o8XeEmx2ANj7Cu0CpQ5NBTS
eBsu/ascuMiVk1qyOSQaG0mg0YVki0I9LGmBjvRt1WEcqxLqXSh0KRLTcetPDxzu
6Qv5BjwZtsh/KhyOX0evJ9bww/yxLvUDQ3cb4Vz9st1lRVicdOfOM2OEmfSq15j0
o8WYR5aPFg6h3+awKcqp7aIvMcssQeZEj6TGM1dLhZaCswuNaDnkoWzvYHi6aTKM
KKx52PWQ8JonCUvy2IN+5dzJa8GuzGOVO27K5UspEARABsaq8ljzNy4bMmlePpj6
Gz0AqTmgZn51xCjaFiOeV4cAvpjCBnI0vT9O1lrF3PSzO38VUWqXNHYa+eGPSm5c
L+1KEReWXf+pJom2/MaU8FyIDh1hz6SerJmhNCFDN2GhXvUjB6U189kSz6oc/FGR
Tvnrbu/iSRglrNF/VE8vx4BTawW0zP3XtJVQXjVraETd4rYq2mHQqSSo1GbeNXOk
EulSP/v/zbzLsVkkg2DxBUM0U63yRPRodhaCzfDABy/T8X7+gpoggdVUGc5rThXs
zOGW+ZUzi0Tm2+JKpm+aJ7yi0rKXwb15foWdfWqgOqr09iTxogDWJNBMe7DEfqOH
lA6v4LSyCZqTulB1JQ7Opq4SDoCwp9oY1MIDCKQGIACYUBu18+oH07dbi9vehc1r
ZNkOni9rblz0lIEWVeJ57Fn0DWbrcs2QiHReYqfu8q8+AxRl77UXcJj/xurAn+rM
9ottCmWM/QsqFFYnfrXKYVfDOs2drNnMF+nbuqHJTdKxV/Zf1t2S+RBt/3kHL+lG
NDsss9rJFPQ2qzyV9GrC4PgIr9tl9w7uBqkukIU2WK9H9bsKBSwsOfX0cpUW9TzR
jbiYxGT+djxtRS2zGH3vo0SJ3p/78SpPVJriQZ66dS81iMlC3ucoTehnTUKAXlqc
KqAvHOONbY1lIUCFbzPrrQAkFElZk6xJ2V6RIC/HixtZP25hzKeur0S6UrRr3VdK
AuBfPE7mAw9m63BHzpeVejxgBYw1CJARtGzsL71bmid//PQsF5797IIPYFMqbm1o
c3jZYzd0l5L05YoQvMm5hhUUZ8axoxGVKNRSWdNyBtUT4cmq+A0i6OoV+mKyjNfA
LTlOif7jQSQNmesuj9m+AwPeufV+1zfSl2UQb/mhC2r81ZiyM+QnWFI9yB8Yd4r/
csEQddnBeryhjwrM8PVCa47hT2Iem7iXAufcmdUHkOOUjA7/hJekC+evn5x3s7BJ
/ME86xzcTpGpVw/WeGflbTnBaKxtDfQxcjatX0/WuTRqsQ3leSWwfE7dmqEFdeXF
5g0JVrDwgNLXw1oxEwZ+dgpolBn12OlIgrc7379g5iSZBuKIX6yD+oJAiU44F8C7
mz3yIwX8FnlXj2V5v6YkWge/JGwbmugB0kZGodkZ8OEtdkab7IRjPFYLAIGu9gXO
v+DSFBFy+cEIdxamRnuGkLF3p44n7PMLjHanESQuze/7GDa50gjxf6Sl27kSF+Ez
nEfJPSOC7aS++D/dEj6KL95dSlCX/9rmaRMEwYO9J8iJ9LNpfl3dVUo0Zy1dm+CL
HiaZAP7ge62JOJif+Hc9vgIXupG92y9GOHt3Ao3stq97c42gVAomcqawHNbvEQMl
hDKhkhPZHU+MnSiNitkUJYYkA9+rB98hhxBzwWfW8XD0eIzRM4BUItY7SuuZR0RE
JfMXFGu96VAMctGZk5A8QrM/W8nv0PQRlCPVGayetLPIjVYihU0JX6C/Sye5dL+M
hNbZx0ar7IwCVTNZ9WOqf76DsY1/12eCyNxcciRxsipIW92pqikZs2eWFDZBC5EV
wBg0OgnB431AkVUnq81CgaeXdL4JNrdmJBKYxitK58OqxFikSA1jta4hyTh/IRaO
bpVIT7SExKawuq3UftsndR1LI9XyghXLbKdsrhBUr0idrAWyS9/LIHZdOiHgNkex
PyZgAl18X4GRwnKovneg8E0aDCCd0LXK6XWl4cV+srFyXuSpuLsOv/AMtfpnd0tE
WVOgTBIfU6PU0wN0vCg7/IKp46TSamYODRt6edWpHNCCsPTrnOp8/7MOwxMLM8BH
GvJ+V5xOwHU1krD662gbKWu0QuTSolDbUHoDGSwaxaQDqaS4VcCmYmyuihGbqCzf
+s9kYERiPHeLReimgwhyFsFnj4dxzFPl5C5tDKRufQNtgvkHSsaCpfZu3f8ze7BU
3I5ISRXCKAdzYaVE+pUuwxeT/G7UlWH28a55EDeUjNdHiuv6yrvIRj933yXDtRJy
pSOuKhVP9wOIcL2cf4yF92xZtMWECra4c/a9rjnwRHYmjEmLPvE78JrOKt3rgzD1
R53nywG8ViN/0OdrgXpom4Kbvtvv8FEspOmpPd/ZraSwHKa8ev5Yk7H6D0bTjXV/
hX9PVLrYY9vgelaL3PiJVrUHVjazFgrleEcZkBb/pQR842/4kWoHGXM+A+knmhwf
7Dc2TSrCfKuc8oAyG2FoWNQStl4YCi8v/28AX7gtfmEk28WGjr/zSl1Vc6QFIeKr
boh5fjRc/OuGED1UPTVJWG+ps8+YLy+ozq56bVh7+kjSxZALl/1tOgibJt2eRBoE
nxTYLOLWySX3+IXMlN3jC8HKDd6aH7mXO/n4cM5Za2X0p5nXLTEopdmyjA9VP5v8
LXvn8okgC2c7YlKMgmbZojQGiFOWmDJUbtjsC9yaEKIIlkVLhQACLW5cDzqRD6E6
TqT8c+ADT1sKDA0U7rlms0VFLzikKum3C4F7u/ucziPjYgYZ7cfq7fwDU5h5GHsw
YJxOVlrGW1oZHTVli5XvW4TlHY3e5QiFzYG0TFKcLYnMahH/z5nrgC+rn0SWCEDX
nX36lzIxEBRR66/L6s/yrLjffhsh0pNuyqPcU0jhfgT0ScadW4vDI8yvf0jLf6Ql
t6vXPzXeJTCEkcTRN8yAnGPQKADa7Nn9cTY+k62cx+5e25JmcCETKextzZh/Jo4S
b5jsB8xcBlabJNMmZldgrtK/A1funf1nG+2hDl89iDMqNUOjCz+VLlhyOaLqPkb8
f6Xr0IcSB5OKjFvObKGcgVuxvOasw147N//1mkTEyNHIA3x4CvWU2EmfZmZNPILF
vUbFI6pd/IV8jZBGqiUDNPL+8kwFocwYY+bmibgjj3HwJqUfy4Pg9b1ZasbW/Fzy
gQsptvut6jFAKnI/85zgCIr2KgxxG1LYUDLqnbZamzo0Ulzv24n+bvow5hcV1mJt
Dkr0Mc9EHd84YI7W5PJKUJmwfNC+zhPOEP9I1d3Vih+n4RmTAYSdxA2h4NZDrlFi
ZbwIL4JpO4wyKIGh0rGTgl+hSz+6AO4j8SSnQoDpfsuAkV/SXbRY4bivqtIvIiSq
apttDz2svRE4XVUlEDosAuQ2E/8J/eWid3hS9D/jeFmOzkntuXHfNNCgZzuqif2S
cswmj34MkZ8JZhxPTN6yF0y93TYVxSl6yRcYhV50JMRlux0j7EkDwuvuTmj0Bt7W
BgJnaRYJdt2p2K+OeowOJX3nE1X8Y+r2gAqxOCSP7REQJ1l3Otd7v6MMb4QVVlBw
+l5tDuOfkNKpn7g6jzXB2KOZ3a0DVe0IvuzGXQJ18FnFSsY3nyrlFbneylLsE/mH
Pt4zsac2nle5oqTsDdLP+dftBFwbBAlgMCzp1vNu/Hite1kt3mDxi2nvFNzlslOG
7G4gl+ygsjqE6bcDVFSn0HgyiPjsP0J6CeEBWSu2IlZ8wO0jhpG2IYslBXifC3j0
TmR2rWUDX8qgE5c0ZTHMM24oYrIjY3QmALEqSxlPVaa41x0PvdejnLaG9PhoMS05
T+Y8skbUEhzyXBzjv1htqwzO7/m7Pe8ABe8X5N9yzY55SZF+tFXBmGO/+Xw9yE/R
hQyg9WSOgx28jUvgZw4nWgZ27g+Nt+CoIqUPFvmhoOB82jEzTFvoxG3xFHtQ8yC5
+g5Uwn5jxRF/Xya4vDDUH+pg4Fo5zVU9QZU/4JtokyFMkTDzILOl00U+32/6k4e2
pq2AWVis1C4uF6MqmW6vYWp5bDq7obiXZSH8g3/NikIeW+Q/L9xhsO1gZT/Ol3fV
ZjIsvgSsn6hHqaOghVUmky37JmTJ58BEzAuWStSBQ6tR23n5AsTI9uBdhMfFN1G6
zk8liPGw4RPyh6rYAJn09KVd93/C7ElTAEOTGjrp0vQvLHEWnxS+/4x+xXABHEth
r8W3v5i2Q2Ul0xwGK85He9v8Zx6taeYKCGWmc0k7Z4iTMDDooToCVsV5Z1yk3TQK
6a+sprHgkQJd8MRt3hb6kmOf5QuvPE8auF9j24JUDaoRArkKmjfKKmUAivEbLDr0
8TylNENGA1sigQVYAy8IsjS/ErswtJnk5NvAoKffWeyErRX11nrG9hZhVwQ7cjwk
EqE1/7cBKrHxB4qHC45TlqBOUPD4bq//HYJlw6HeTdm9XxVKNL1ZM4DR1+atGRYf
RdILMVzt0FASpZ+RKEfI5adLAzaod+QNrQW0odTEcbc1c3TiqirmmPoIiKZ4zvbY
E8Js9b0u8allE2wG73xfeeGQLmT64jH0hx3v6/UB88KNvXs3Oy5JNFdn61/9vUqy
p3+Tdl/IxaALKAPDot/iiv/MQByoQNFiNpTfpr6KWRiuJ7Z+jiLQqdUhUvYjHYFR
yGM777yXNwsqmWkJunJW9O9iZ0lPBPSPkeJFjXDzPBfs5dFPqUK5r150xo0c2hj5
x0dnKPsVnKw6IPdedLYvboQXVYZCGXI091xtyKqK/QfVh9gET9U4jFrnWOb6OE5b
ysezZ8KEw+qQHbArNa/mYfu1D3EmVImU9ljSpIdsaCvw5KJq2zdOvMYEm1rOveFc
8/FdahxhbYK17AAl+dDfPzXcT1zquRUfvAgjM8vfGVKSwdGUzwfvWUE2LtC4UtFB
PdqhP+la31qJDQr082ypYYJBCu4lzKlT11PCCQkSFnPQ5/X3ceEMk+e+R5rDM1L9
GfnExriPT+kfqoHl1jPlBmdaeBAsM72M++id0bzaBy4barI6AcOM1S9DNptCCXEW
WwD24gPozJ5asf8ElWUOmnPq0ulFeCO5swt3C5fx1faW1xg9BbuelOuEJUIO/b/N
olDp1NPFWp4eoT7L1ZoafF1eEFeqTTe9UgUskFkXtm9QSWDyKeVB9lkquI+7zPpz
FELMHtW+p9pxgvdPZ55PhvyNOgHEMVfsidCcr/ausULBuc4ly0GxagvDW1Pmn2XF
wFyJAsB6K5y7PkNQ8G5czGJxEpTaaFVhgprdxa0+DrA/nu8Wi+TYYZH3ELTJe3zR
oOZxlXdPnOeFwou4qgW2X5wL+jT3nXGU57flGSxHWNPpykAq5VVD1Mwx/J5FMdPL
linc772vig9zajFArue1u4fqsxJ3E25wB/JHf9es9VyVxO/MOG0lGVLD7zqHO598
TCDX9tCykPyk+aPO//WcEBVyYzvFNbPnD/ZH5aAIB0ewN0IYi6ThjUmB8sdkRz0A
mTEfry6zUMO4mJzHpOG5U8rMOMlKaiogFvaKkOgAKER8hQGH0jKjC9+8jJBaNkHW
epzxurSV89L1c6/YafYe+qhj+XQAEju3MQ8bE7liNBzKsL+xC0VAXd16BQAtYgTQ
Gps5CC8JWL7GStOTbrTw867x/uFDO0GaXSv7dfETdcCtjGm2wJfEBjolAr0BVaQX
UhVdYJkUBLdHfu2fvL7XU2oI4U4/+bJDbgd+LNuIQU+7kGhlHlhWYTsjv+WtXHaW
4r6PCJyCyBB5QVcW+s1i1qtL483vBtduEw95UVSTOE9bBfX1YYaPugI8QUGfFPJy
V8pSZ5UQh2YcocRwu/8kHDKVxw8sfzPToGdOn9b+tW0rp7R0WRweDTgbuN0U4jJ8
h00nchG7qBgljUXIJ0e6rsbuHAK5/cXxKr056j774Xk9YKgWFsFZ6+fDZArUvMMM
RO6VYlF7AaZFViJ71O48mgJ4N07yPoOBqrCBXl+WleewE+K1Werd6/oNT3Rzr1uR
+X89Wj+upZjYQucQ55srnV/OyGlRoazmRnL+9/8bqWYe4VNcA9wqbheP5mJ3zKVS
ni5UxGwk8N2ynzx0QkH5LOzt3ryHn1Oe4sCFAeSkB0sYr2f+U0TC9jXMaiDNwskx
pJAqfZmv7o3tLK9XsJovBSbFYzaYRAgFgLdLoDDorGvbURlQ8BehOWTUlnlwFAKI
Ajq8TFjLtX6v5ehmZ3dg/lbSpHUJQ0YwOFfO7cF+7P4MNC0o+p6ounOfUdn0Dxdx
+B8g6/BN2K3itRPNV8u63QQij2KY0BtdZ5ji9g1vLVIwzIAjvZOYZ0hdH/JVH8+9
Q1CdsBP3+ayoWZKb42lh5egnW5s1b5fErcIckeBVeacRWX7jza2S+SzMDtZe9GU0
woC/Cc0FIn3jnWM4iT61eZ13twNapcTog7FvqQshdF2h3PaGjAommW+2zqkoDy8j
pLcsKCIHJkWh4CJ0nB4nwGn6L1ksi/RzKGWUxJbJXlQQvX3sRLiLwc/1ExtBzcE+
jaA/5au3zhvTsKts+3vZqOQjXA/Ao3yeZ8EUcA8DoGPEmm/bV9SGPL7QPoKht+c+
2Po5pYDa2eB7UZUfPvNojS6O2l+IwqVXsMb0XQ9XmEJGNytfzR091Azpsb9yXznr
KLPm6ui5A6vREKoPSDRCnmQ5vDIQDyGnDpgzGPBsE2456Lga2/PDqAkatd6lRGgn
O21hEOMuk5mx03yzTZ9XKW9HBaZE+wX9qFn3XKkOZTkCVaUPE4uoc0bQivoHKAaR
D8RgR67Aajzf0tGH/N1mXsdFl0R8Jntq8uXrIV6U8nv8sYNppmklmaJCPp5QVK3Y
ZvwN9aX3SRsWasqUmh/4WAGUlPQ4es4oPmAGeoH7HunOv8tTzJnpFgrlzpB6AUNu
KIp18wTAJRdzaJ17KUUp+oXnGxCZp/c2H2i/0LaS9N1uimsomq986qn2b/NFdgfF
rTp5mw8Zh3mOQZT/Mmh3b4dhJVErRC2/yVKEhbQyhXPUQyihWbR9N3McrONFbEOe
JmvtZ+JdpoO14lw69aGTrTKMfhqRxM2rCmsIrn9g4mHO0GqaurllRxVQFhtNOzGF
52rcrqF36SWPEkIegqit8yyu/r2E28zfnOppDC//rV1QRyJ9pqNihX/XlkUT6D37
aB20aSUJbIbqiu5nGjcWoLw8X+H5N9kDZTz6F0t4/1mwM/cozyO1oO2psblOfM2K
IYqmH7DMgw/fo0A4BHnwIvo7TRKiW0RaIFvU/7kp6nqau7W/SpS1y7jN2j0NEckq
TFJKiWxTb4Q0FOheHOjuplfwBWRIqVm6ig8Hm3D3PwRGUakz9ENQ+o8auHf65nhU
nQje3Ipz41mld/F6nkp87W0mgscSRt1y9Oc96UiPEzNPux9wbXU877lSYG8QTwJZ
VA30bLKQeEOx68Mg0X3JE7zioHQ+9fWTP1mhcnogAScJNou0V71sBJREWSVKb0PD
4i9ZhALav6jjAdGVfbW1gg==
//pragma protect end_data_block
//pragma protect digest_block
NkYSys2JWZnM8YgFwyE9HRUcFXo=
//pragma protect end_digest_block
//pragma protect end_protected
