// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
mzETyGGXcjFMNDBbs0nMnoDPA47pC94p2GwAbsTXjTnor5E05votL3WwdeIPPo6s
uv3j/ns8E+g50VGwUDJXjJyojpHW7Pe4joc/RNnitdWCpt5LFTzRNjs9NvrfgBqe
p3tc0MOrn4BmFQ4quD+/QCTo+ZOmiZqQuSusQfzzDGNId6aURBFtGQ==
//pragma protect end_key_block
//pragma protect digest_block
jCm44IHHaj5atQzCBwo+89J+l+U=
//pragma protect end_digest_block
//pragma protect data_block
K0i6yBPc/2qGLP5cHmNOswWstB3h/dfGiMWbyFt/DUXKaoMUOZnUr5bQqFGlqqRv
bjfWFXdzBqpyFSa/SMUVNM2uV8/lBHlN81hp08c7GFgLs4EjPFqX8ELWlhJibfwG
QvdIrz9h+3iodgzTBWtP77KkHFRmxDijYmv8Zqn6G4+zgZQ0QTujTQRwHK+yIXSd
9F5LuBggJeR6ctJ9ct5LpW3ZTqYXP9oHGPIBWP0PiM6DF+pZ575O/EoQu13W6ze/
IAV5V7yMtsw6GxGZsVy+rWdPkIIdC3o6BuDixuf4CMTHeIXnR3iRWzi+aP/C7Eaa
C39ef+cnZNeujG+AkQWLUM2DQI4CY6t7OaTAEW2WoZgZiVoAxUssBjqt+NksGo+D
exOpx9zJRN/jj/RsD+6arSt8TCqpOeBf0P6v6vTWOS5aebs7X2LYUnd9Zo5w4Otn
MSiUcvYPhxDzcpR43f19KKQsy6RweTQKEc8sE0qEZlGaipHM7zLRMaeezFboDZAe
soCh/Cz2ZCBQD5np0aG0xYFm21Vr/bvaKY/6guyKrTqY9RoYnazx+UpeMA3HsSkE
TzuUvaaBJX82r0Gt7t1hwQzYQwkiHpOUJe7Xgl6QzDfhb82K44t9XqcKUed2gqMa
pLKFw9cOdC3H0ZwZx84B89CBwt96texAsXxorR6EW1dgkvq/IuCjBXzorBEaySIN
biRtZmphyE9v2X7fzqttHVXr1lPinmHmKvHML+qLlRyIy0ytkQsHgvxemfafAtGV
dbnWyvTKwi8ija0QOQ+mrrlP2c77cIYuPvd8woeZTmrHIoqMjP0An5r2Q03X2OqJ
jdtACScCThPR8S7RmCTagVK8AVd3F25W6rg8xBAwqBMZaDe1vEQga7gt0siVfusI
JM72fE4Ic0aBqrBengpW1BZYRqB5H5Os8FNA+K043QHDC4uTYNIyw3aV/XTZUpLJ
iz/ROiEXXlE2DYsVYt1ceUzrC/h+JPHyOW0US1UGk8FJGQwUbPU5n/VTO8xF458n
Y32g4neXTLdce2akg0A2Nuj9GfZvfN/HnVVQ+Z4vIShq8Q4b9EaUdHVKxpGQaIrG
KTo3kYlctSv40EaNffQemHaQksnM3o9sOm91WWpKd7Ku3kE8MRFATqNkIVZwgw2r
mTEWP0BFy7bbex3iP5XK3AUcDzxK2rC6kzvKvEpggxRnPqIf8FXl9ymCinodg9RE
c9cEvkhawoAq/TAHdZwKDFnk89otu2NRfB9ltt1+QFa32wG+MIcMLEER1djpgpUF
W1VftRrWwzD0gYcq3P7HK9sKlr0tr6nZs+LiYbRuyk+zzaEnczMsNqaav8Jgt0vI
O3FaFBAwlFwsbNFoEF7CxMcXd9jlT0DSbwG/y535hGsGDJFTDKywepA/FvD8gXHV
V9i6S2aM/rj27MAhT4a/pnCcWT6cEHwuU9NSDVA13rz+YHB6zNfjhKMHD/TnHhlB
ZDhgiKU2212tHbKaSR+aEb6Om7hfuhYSDOfzA7iTMRV3g6e/8lQK3xj2rFjemBQc
fG3om1TNlGGruE8kQODnS+U5kdeX2v8rq/8oYP5PEGlcwmGhvTreph4usmPzhi3g
m8Iq8pmJ9i+kGE3BiEseXLdEm60kD2Ea/Wah1nTSevKDsyCcy7Mu3JBil+3wEjm/
s5i5z1UgOaJS74JrY4zRb6AmSDdb4Z/FKqyGB8NEwReXryoRhLbSlMM4a47MVVaZ
31TAprXeq7ZlX55D5Q+KnocIvIsb2r9AZu9pztIsQKOvP3YSSH/iTiIiU5Pdg+a0
8saVQLuvp7TX9W8JFzRoqmOyNkd2cb100ylaMmheFh3uhe1tRORlTbCIvec+LE1x
GzuxOFTUSf5yoT8usx/MVK6ng+kfOyrVS9UN8Zbhp0r3YQCoFsQq9atsqT591PBa
W1CK8vB8iXqjl/k2a1EIn1jI5Oc0lpIiBncobec5Ca5gEIialLzr7lXvBMxFwfpV
2JsuSPCOAVlTVGUskfctsTS7nvxXLVdFgZrKrEgyb84/SkNhr6+xyApyqWZ4popK
/y4TaX0VGI//QDIiV+EAEkbGZdEBNoTDgX+9VdCop/it9oHJev0IZB+548A43RY2
ees1qWbO5AYylO0ojAzqOUlUNyioAnc98bjKgjWRYhWabvGpHPUhiFVpbEzEMmOr
lSQ3oFPPq6WUTQtWGHVTBGFbgAtCCfk/K6Y3to76O/Bq7nunWOjZFwiDyCbDHpP+
PuAneQxbKNwtrNEMBtas8r2zcecSTGqSbdZreJ+ubuEGdtDwMmEa3T8hrmDLQVmw
I/Yp1GKHLWnGPNRBkqdXYHviKgiyeVXLMRLI0gekFw96A7taHDnxpdxzEIklR4BX
qTpnIz1KLIHEodiFZo5/kgHAEBzwouRSdnMjkz4Tr6N1j59S9JBuNCClvTcUKqTu
ggdu36Z6l7/lMu87nxc1nBwjH+P6qMbCffEwdbilOoGHDfr67d+DVbmvC9Tswxmv
SSEqmzK2u8TOyxRpa6+pdM/QmU1DAvz7nQsCzUqtFFy0FuWLCCTupBGEVAri9G4c
fmESHpNvO557YDbwgq4cpBdeUVZDDlvEjA/een7FXgvonX9rysZd26eEJfD5Q7I4
1jR4NxyncCpEsc4kSL+dnkCYjlwDlQhaS306Lk1TfEquC2/V/p7lJIjocve47AP3
fvBACWfnpFPwiETHhBaO1FXcFL2aMkKQDt/bM0jWl/BxA0p1WEESU+6vZYByfqTx
HAM+FkJYm0+kZgE2292L2fSN9KjFhHEn1StKbCdA729MeJxD3WukbSIlfLUweNIK
tKea4TE85bxFD9ahcCJeRPksBSir7tM+jIXBDE7dYLUI3eQUytm6gwDIJodu8awo
rQzHRb5YvvbXihosms66NrAgBFL+McNnDbFwRbxtQk7wVAkS1bi9915+NqXhZwm+
zKB2uYzKgIE/dx2ajldSRyaVaeeeVlYgeZmoUy+N2VLIRqYsVEQzrzsGVYiZrlWA
xDM9HhUEC/o1sRfQOggpTn0GaZ4I6FEJ4kFqbSgdKJtsfW7tMrdgjhSLP5PHriDs
W07TvqdCtMbqUWkgGV26NsVcvXDjZyWq5GFlCbdQVWv6YFTuKiJDxVBfCc8ClFXe
vyzoQFMunDI5RbZvzB7WeLWuqp0x4W9DtbfuFVrwULyqkkAxZ6+tSfXIcc2BfldU
kilAFnm2jI6Ciw4wBW3UzJa8d1pR4nOP2si7X8Jy5RsCTHXYWybOH1hSArWW2NHD
g+bK7mvNrZLKSBNDqSjmg2dDivmRfLTmcKhYJ2njlzT3XNNi6ZgbazVrtPYjgVkI
6eQXSJa2QT41chanufgu0UrrB+HorlzvkniFPHlqddDOF2eoHhRgqAZEdb51COyV
RSuTQXY6xjjualkFNBLR0gdKI8LoLdxivvCt9ZWSoi4o3slD6xtIoclsa8Qi5DJK
ifsXvqmOIKNuoNL0n0yFGwERd1Zu89/7WM0OFSRcDiGg05Bmju70ss8bECay4pfN
WlLm0Puk4wmH1hHzSnlAhdYVxqn0cPAw3pd2joa3Hvoje+QqwKTF0RyIjLxZTyJ9
LK7djrCq2KcpM1kYSC4a+w0VO5a4PRDgYz1C44v8du0S6LH1m1gFdtnbPiCH09I6
RPIv9xDMGS7fzMffzdBRnBeFYfltthClmZtapXI56hIWWxbGk9NP6Y262b+PUSHe
TDRqt2gKfJi4mjhc5FeMJ+BDkSMETUK8OrNCmo3Cs4aOESPgouwXQGI6Gyz2gZ1y
63A21fyKg0vhw00EEZ/nPtMDQGyQxQpg3rcBNqGd3UH8wM5uBsjuhxmfAErXhWUC
oR0dNT5/Ktoy2/byyH6Mb5S8yufsXA0icnAUlrcZKhVpkSiaroo/+MYzdFYc9aEQ
CwJqamdyipJi6pReYxn/lhfF1vnbcea9AltFQiaMhXkdfDd0SigJItw3WdWR7rGS
0tYDMdig8H1ajHUogh/G+kKQ9yGfftle1ls/fFA7MsaNZfZkf3bKVUoPbNq3iJBY
XGpR/aV1w7vC6P6Cyy30QNwgCpnbfDrdfGkWqAmcjObz8vlutzcutGPL/Y2KCmN0
pu2XC4VFKa+x5h2RJk8KkisTYon2sk0zrcUWyNvT4lNQwNq/nkIA1vppIVvT12Mf
i+jsKf7AETptRzxJS/yDRfW22bvlX3XJ4NxDhpkRwx+kohZLs/62kiY14uog0HpO
Jf4RAXRlMRQIu5T8IO7lzhv7cNexQEKDjZsuUuutqbqOq7PJ36pV1On7HIspp5H4
ZFDlPGmMSPEvrByZX4shTRfyOkuLwNAsbeteE5CL0nslD1lVabORrYDmMk79d4Py
JkwjfN3AU3qBrz4wV+y4N4dBU3fo8UZkdEdepK8SXbgsFooLVe9hv+DzELR0Bc+p
JYKTICnWOtGzAjLonl7sdFHJ4VQjsmVHOY0SQg0z90ufEmSSlE5mgCMNkZi2LPZM
de0eM3KC8V58t0+yJOulFbOOs1QuyCeKeFvJI0ICI1scfogPR0klKmb6edZ3nM5Z
mjxr9sCW1LS1tHwG50Q6CPOqzNqYxyS7P0DiJe+gv2qJuqGUhQQe9X0g3xpl64vj
03rsHiFsP+8u744g/b37VkWU83MOONbP8kzTg73dNCaUUUVJg2S66SfLo/p0t6Cs
TiEHA3FVEYKbKrkoHOkKIARBj3Etg2RtqDEminr/GzC63IXWM02F/CH61U3oZq0p
3qSsiu6Ru3e+PBsf21hq6FCrqguqB2Z5CAbaflDgHtjBl6dvfaH3MilLALt3jure
O/BXlykbu76rOjECLd7BAStdim3oSwECYUskeaQRcvAQC9jh4wpw6PctVVkpBrGN
wwnY7MNJD5i1XYbxxK6eaBdGHwDRd8DtQNQyVZV/U1/9nstGp77nHRFNort+jhNN
ecaxWfrt5RImaplGHifxAIS+FxixhYwKCM14xbo+UPtcoUlR2ouqHmDc0b956w9x
txdMmles/5+4kxjXBg21qSWL4zSopLXLhoUFn6jHt30BwIzVHkVs24xnZNIsPcqu
W/KoBIUmYvAu7hTQ3VI+ZQHH5ScBuveJuJAk7f3hYcvNdIgQsi1XC75bJN1bRzk5
+UVOFbr1iPXZgrvWYPALYzvI8jH6zdTow+sbd5E4VbFuuWrMVYDFG5XzZF+Jl1ck
IcaaeMqGH4PCCiUwLLvTKU1Kyk3+qhPBKjv+5GcYExQguRHmHc7lFAW/Y8YQZTEN
iHwvbL1yIdXjS442tSongWL1KJiPC439KGRaxNT6N+HECULXT1n+YS+CmKq/Ukhg
D3+bvLowqtkbXKUqedVdpLddLh8jo538yavCE2ZXxA/BnXoOZEle+UeN9S+ZQ3nb
nzQrInyK5V3e4J2OXDJwcF6fCcDXw9iTqSV1PX42rCaVtZgpSJp73Or4WKSvxnFW
K7MKKxiVuKxf/7dGQruWBcfmVG+7cK9jg34BpuHP2N50XeUmEKI/28bVT70aVHar
GEWYKs0GoZMSr6coJjyYExSaJsRC64Hu9fa+d/VoBOsv8Jxsg7H5zpgcCiQmckGu
XNJ4Nki13D1aQ07a0Q6HsbCAcDNF3qnzpKw0nJNlM3S0zGdAZ4Wqs6ENXeMCB6nQ
mI0fR/HEE5B6X1aRqA42qkn6JclU0NPD/kxif6wcUJo0xJNyQga2Dhmads8lIn2f
TFdbLXdrEIGbadEUM5N1ItiZN4fEClUdA6gEsYUQNx+UAYwydL/sF5lBDvRk4VZD
FdnjYSI6YMom0CUpmHpALUFq7R1RbyThhUeg4gu4tIz22tL8QB2NT/wNb4H2SkWN
9Y+ALaTx7iVWDyaQh0LKne/SaM1Gss2Hhqq4X5+afHzgLbJDFcFi2CrC9Gwuqabe
2H+99UY5+dnRxaCUeoVnHUExFSpjr5jvSVbcwCafFUR4amwb6j6lMIpdBSpMvRpX
cnJqIeOm/lkrcSHsT26GzGoQRVwls5j1Tgt3sm4VV+E2Hn++/L8ozTtdIOV0FM2a
V0M2jrIQEv3WNdRRNdC+BCDoR5+8LdbkAxp4SribsdLD0pDXaFwc02HZOCyd7v4o
ArBCkPikOT6S8aaxGyyq1b51RVsG+R02BtSubv+PVOpo9tRAAsOYAH1bvb8S4zbE
zplra+TVyLRGmMtLf0nFPpEVOIub4PWSP+EraGvtFMJQQ3YEXDcsGOAMIjz3Tp95
TEkQcokc9ISBKEXFTTzG76rrf93QoquCLTZPfWJLhHqW7Tn0GbdrLdYLJaX7A981
69UVcrQoxXPcZdnCdCQsY2aAxpzL91EcFXiIqJxichSjhtc9YDuAZNKIYOWsULLn
ThSmJDFJdzaCyR9RENfpmsJEcvBdWm1LhYowxHUKDE7vj8d2wm1wyGQhx+uXblE+
Eevt8omAxd2+OIg7yfKymxfMzxKLQs655l2fqOPuA9VJJpu1+Y2B5RALnNW59GXi
E1TCrLHclPbcdiKS1qT/YPsXg0Ue4bipsrqEUcrUTW2dxULcjCXTsdglBJhByCky
HNQXeEN8iUN3O0Q/V6zdv/ur5V2yunUQo9lGtdcliLNYnztig3JaYB0pc49RrGaq
UAqX4/qB6nCpzoDdbh5GQHjCld7/iW2wsjX5Vn1LjXhTeJoon+fm1HY19ZsEg09T
GVO86WBdD2ki++dpJBKZJ5c/9VnXE4aF252AINqb+g6u2+ZpLaIsFlURpsXcveOq
UUtSoQtdOEoGCpYHpkgatmLg/Z8SXNQWG7vGHgF1mdW3DoYuUVgZmzXqH+Ow7UMa
kcCKw3wQkbYeNXP0d4JqgXQtaKqyUx/hs49n4yDDnCVmo8sh0reHB6PFZs98i8lE
0BwdokBwj5PscUfzmVzb6X/hM51o/1Mx/ITD0AHw+ph8KcSPvXWt1lCca99JVvIO
ZYmZ/yRUIilQCFBYwWNYICScTsynBgVLjepFtKzjjqRNWgOD/IX2qn/VlmBK+nF2
qryx6/hv6OrQRlgbXUsd12RNOIzSMdfbwzjgBOXJbIDmzqFoxzrB+OE3xW7X4kTy
foOPmvW8OvlR/Nf9bn49gL0YXaBnTImR3J3q6ydRmVbYs+sv+CK735c5eQn9a8Mp
uJYHpFsg2ep5+zsVfA5ed57JjDImx8Qr4f5/8sXfyT1nTf8/h4Wk1DK3PEDYBijh
6yd5BmzN/54+63bVDHqrmeQAL31dX72ihfojIJ+nln9HvtPK2ODvM2eiMWkiRZLh
oO8Ca3oKokN7hoGi2u0K5iTCm3BdZFKyyzEtr/a4yp+p16lLgR9bw4DigAX8tAmM
rP04xTYCXSKNcsGGS4vRrMrX2RTe8Y4M9Yijh4uOqkgGLcE3R9vSw7mMN4s1yJh9
1BeyPuMdJ+Mzrup4hJrNWjxYvSkyUFu7KsM67eoXctxqe2TgCggTPKbQizlyG/IB
BLMcEzoGGRrXpMH2nZxSz1DlTLZTerymVx8ArMNUZZj0tcbEswk7BqDV4J+3M3cc
Rzoj2m02N925IN8o7JWVgNPNsqeXcjzLYoH6GKcU8lY+qWcwirwswZn9zZ25pesH
IHjB9vSQKd4Fo+sIXxFhuVquuxE7tbhnLfLOo3GmK4XoX37GURodALkv2ejgIEKB
cj29Anzje4J0KIwISu9K8Ni4eBuipieBnOEnCRg1R6cf7zvZdU96i/TerrylZQPv
+/yzcYwBvvcKGLhyWab1/XvmVmImbf7muFdaTa3KV/LiJ52GqlqI0VkWGsT98RfA
lB+WCg/ZZKCQ79cI7YuBYYCCWYm0DPFx08zNfcbxLhjcDMZoSlVJWswG5TWYfkic
xtqxooA1XZCVzLQHNytxMXdxf88R7Y3dCPkBvq3ITFxPYewfr6N+Pj6MvceE4EhN
eS6E+Vzu0fsavLefm53KyNXTyKktlMJ7W2kUqM0xaCUZSAZY7VCByDZ9zd0HudAm
rwUjtu9eGe+DdSP5d3DiW7MWhjCMylqURcBaRTE5daYuwatU97FGZ0TE15sHejR2
D6Y4LUSGwglZ+hhhbZgqeRGPI+rdCjnyg3P+6C4KyJoT4VOI61q9zJuhQ/+pjwVo
hAL6FqtxyH6y4Ae2gxm/hEpdiwoaTSCIqRoWN0QjPNsQGi0sMpSBSUr1tzC+G+eD
izddTtlhjhE7yUYA5649U/mWKZ1RuWU5D76OQo+hzfxhlhtElb/DdApMeYGWkJ3k
Z6garDHdNJNuwResc3Dp9ifDTmHeRN8iWKcMtgEfr4QPmB2gjqakWh2GOw4H4y1J
pAd4AVPa5DA6wnC/Sb/h7fDna6Zg8Fo6xYKijxp0k1XifbRGyNGCACz/SEYo3M0p
S5eMcWGTiVhfQIVJxZ7GKc0p81Ln/RYjYnCWgp8Zg2vYF44/OfgkPcyRxKJOQE3g
hZdxp5FJiMvMVIMtb3lN96T60plE32zRrOHmlM9aRbbx+hSRJzXXV6O9JFSQyHpk
oEFmmvNa9+2eNrPWjKvJMCmMeIrFV8pG1sNpZRCTXgSTYQZIgnw8KBaFao1YxGdw
D44mTuIaioA3ZOlSCLB71oDYpWsx1Tr8DvhyJEcPI5YxdkukXyWAIs8mwtFTkPTN
nssqjnGQbMftOhz6O9mXXtTMxXvXmCBp0hVWP+ZLzF4cMs2Q/nc6n+hpHf9CF8AN
quY7rj1Fq4J372VKxuZiAAjd9Ih7XuNsoBBaqOQqqhigpQPCxr31JYx6CBS+G9av
fdHIEEO3SEQ9SoWcumRJ/bg7nqIi+rzHe06ltX+Saf7Y/ifi9mUmcPygeHq4zmHU
4q16VwTVit81FHEEBUTvuv6mR4t7l2izj4GVllI9+BXEyIbUQxjREfW8S0dkgfYM
ibltowqGTdNkLTL/C0Wq4vy4gKDyRsByXpaPrEL3adncixbWjgQJYrmANSHXWJcc
sDhplAXRgnmTZITHhFolQLiUrhAbPy1vN6nqMMTkS5QJ19NmKFMFTp4oip1xShbu
e4MR0Pwnes2rPCOpU70KmelhugOYccP3PAiHnE9xd3Q7rfIseHpabhHLSOYGbeUR
X1kim7MeOiEItfHK5YMZar4pmpmUdUslx9PfWbRp32TNa+iEQ9+Tlb4Yr8XwTMxR
RqyIAXCeLGdETuDYGB9+mIXz+c4MV15HRs5NlNBMVqD/489JZh5t1OzsUSaiWedp
DBo8iGE4kIqZA7PzNH5eab9DECB5KQo0FfL0qHwBTzTMo7T4pImSMblvrGVYcnki
qZt71Fpdi4xDkQbWgsy3BeHqPHGlDLThFhgDz1mJts02ybi5O6KjeC6YzUNKeGRk
0c2f/8Omnme23WvYh6vjOk8SM2uqqFSy0sJU0nWVJ0LgT2JGqKTeOayt+9J/xyfh
sHcsINo2XyrKH5WjLQ2OyNZzZCqWjfdv8jl9EvwwwOwpP9TBRFZ7fcpFK8u5mVpl
OQhEJITsc216y15AzdYxEvtTS5lVn7e5B/36gYuEeQW9mrCmy/LZSEnUTSl61WTf
es1YSmvSE+JJJfGjMjh7DOfh5urPf5bWK6Ctjp+zYuIanX8rvoMH+JKrcY0Tnt8f
z/YZ/uVfEREP9MHfBKEvNRalLVYiJAOxNW3m61dmRWHTa7rJiofDLKiliUUOZy1f
FxN8tu4B97TEWsm0bj2iKRYogSXASMiaReLUYGvirUwiWVMG03g+YODEWvw9O6VN
iXwjWjNL2J3q58g+E286sN2GhER1afs+4UWKXTvivWTvUl+u/AX0hMYRv/RaCd7k
YWI5eusRFgq8bDuKsobIj8k5eY3IueTomnxDqa5tMZTjEef9hwQmhTPhpqwpenY9
LMen7Uxny52+AcvT7OBKvGFM80yUQdA0pijn4C4LSE1+FeS/K2ZGv2jP3DFe39H0
5MPD8Lsb8fvjxENVV4uFAJ4ZctxFlvBUahdKginRvjfu543W/6w/kQi0cp+IkGnC
+zbJ0m9efY27me4/Ex6tXt6nzgpvs8MTQrbKVFCbJOssE1NX43Ggf3ZdXE3DLiNk
vbqyWe61eTME3PbcuqljuHhecRLgNHyIaEpJkLWRtkAv25uBJpRlqiVkaqTq+1vB
RBQc041o+iEJB3hpQ5w24gBlBtTdjJb8GIc7CCXs8x85iZZXxyg7EBmc2fCfVhF1
pkamqlMn5T2VolDhNWclcePyGU8khZD1Y6KsgEoEn7j3dF9UmvZf/xqRfirAOE1c
oNP9R1BPszMXgDVT1nWElbFXSaJ4nQb8OESitGPDyUHXC6Dzz4FV3qWHCdsgYNpB
3bVXEt0Ny7/XJsPnYXXGDTu+B6zIcCvGNdeP/WagxgoEylvi9jq+p1lgWqFCUNOI
7KnyINCrrzj1Zhzx7bMMd0Yw7+rdNxL8pwusgAiKdRk2UgfxnUN2pIylmXRvkt0D
1DwqSfQFCESQMxMTs2Mz2VKIDbm5mEo7dPlQHJ6V2GgCwLR/p7fuDNL+IcMIAfGD
7Bnh+KkI8AAanrM7UWlIOtxbTk1E28b+WXrwrRE6+Ttp8fwcucwhEO7mB/gsFNrK
mUBvlGiP+oGuKOg7Ni7+JoVOFqm9bbPPbrbz5v8COVMT9RfI0cVQ+Qbx4vMg2LpU
YAkwDNP0bo7eh2Ad8CD7JMk604nPvf2fLq5nLPnIoaJxTTFG9K4kU4n9zMQapT8n
YwdyWDuvfGKnHduyCtF9AJBy+nKkk1VtqJLZA/Rl6pwqcC/mN1QXuCz0mzZnNvFE
J9LOcKvKonr/hG+PqfRoEsJbQDteCZdmltRmsnpC6ubFx1TMAbLXpNBZcUFFpa27
G6+TbvXFD/CtuFc7J0umAWzvyrp/jQL6tpoc9Tf0JlKbOEy9ujKj8yR9xvxbFf7c
MGDI3BmYRFm4zyeu0NGFUKl39BHhM7wU51aOOuYpX3bCsmxSoEjnBVczQ0efHHdY
ZTUlnjjn5kxnXA5zcuuyDZCAg3kz9y6EPthewdU4fXau88GA38nv0+rfYPIKG0MZ
NBYWp7o4b/y5gUMFEx3howvFPRmCKVgqgYCH6IWRao8R1OyqaIC+RGKIVJl8yXkH
CT3gS4Wd7Gx4I5kbDrfJl/RS2PtbpXgnmXSbifqwabaTKq5fUKYLTNh9LcT4YVRX
lpus1wkKZhSz6181bqe/DNfwylTM0BJ21kHlh26+rbhhPfffDYA8NvPHCk/VDTMQ
StTVP5r2QIRixbRsIiNbdHjNzjkD5JtIVH2pO+yV9yLUcgoGpzmIDeXT+HtMTzgr
oy8K3ADgDlamfznxpmqjzQ3ONCW/aIWjco5NU46NeoLNh8+UUK6+rkXDZLpEENoe
B2R2H8HnrQ8gU0YxQ7HXQCdMt0FBB3r8wxgpPyfkl38U/Grshc3FV5xKvphkKziY
pwTImIzhIGuWBrjG+hShigGyEOpDkVu5ux7dxxfP2ya/rHjL4RrZwPpZMvu8DutP
6mUIph8uoVOxaomd/5RbCk66xsgkmfYDdQbOzyY0wOpaoKqJGzkuCTFYPS6d79du
dkMl4Fw0nbyZYamIfMjnrTR8fNd6ahdIkLt75i2/SxvLqFO9UfEHYnkC5vm3FGa/
DQts60pVi1yfuLPe577m9npBuS6rAg5W8+7ZIJNzlq0jNYKLMu4cq5hn9w0m7qoh
6vPBfhG5ANmSm+sqXELRbGoe+Lzz3Gf7SPrynW6FZsUzETXzEgFuXEkzAQh1LRBI

//pragma protect end_data_block
//pragma protect digest_block
BV9oqwKtmNRg5vOF3LYrAU6IKSU=
//pragma protect end_digest_block
//pragma protect end_protected
