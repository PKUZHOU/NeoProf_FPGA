// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
NPouWsiErTaLqtGSVWUZaBgvp+kr9FzPkCaAuiktuo6gvVyqNeKzzIej7gIw
cq12W6b653VIQqORwQk4EKu+GF0kqAnT98CeIEGciSSO0Oe9uz+LDVVDFKgp
GOuHeyDAqY5XydMmUgYuxXVKZwSQPG1aGSus8IGKJLOvcQCON8pht0i3NKpD
yDWpiiKf2NToGKYu9zYjFX5vRlRX9j4mw30aGvvGrFlb//ylOJMDtSSRzFK0
6opl5RaSVeP+W/CYTibcg/awze83q4kqlzDeIgyW9gNGLBDnFYyqR6N33F0R
o2X7YhjugsG6PvaJz3dUNvZpIlCJsvN37HIer0+GeQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
U3XTBmPgM9HfOSNEONm8+TaFpjUH4QbGE12WkpalntkuYDZ1tzx5EXGYYdYS
zf2j7UCin+C6FpGOWkEIKuK/0vQxPtPOelBNGP8XbMOYsxN5h5WHiAnM+eeD
1wTFeyhsb/xkxzAXDLbcZ3CoCm5FoRNWuNYA/RLBmIDBiDevST54V8q5VycN
nbHfN2aJUsFBWN4wwPbjRsrTNTW+E5/3Ts3Wg5qUI4pSslmevikxZhSxUlYP
U8HoCiB4iMveUktIeMLv03DkKB2LCDZ/T1AmZzdbyx9My1kxZOG64c39sszE
Wjbne87hYdUtZkK5ohAxkL2qTCb3UydSRYDbAgiDiA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
MJN8dnovZ8TwiGHOfvANjyaUe997Bfm6OSu8bUPY6AUn2WV4RR5hDFd/VzdK
GqPTt8Nb89k6fqKriXC5bLXJ4wC99rFZXIl568ov2Eks6ooCx4mSjeteGjxI
CMmWYfihnCtAG1jntGiNKSO6DpUWFb7MhJESkvnjehjQfZVLLzCPIORa7pan
c20hknBrl+xXF5XhUWeh/8liFSgMxn7LTepHuWlkYw3RXQthK3GuZsJHwtgr
1DRlN/EHZz7P3d2TOKptHHMPy69+n4Hf2+N5ZnzQ/89aQQxn+o7qUCDXYeFN
+0cP0X2hF8dHEswcgoRidyOrVX86iSJOYg0lA332Ug==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
SVnjxdaWWQNYtfGatzwXgCyA9hJ4WOa6ujzq9/rLEBPtlpUCGfWzU+T749rB
5hBgobU2Z5nJHhln5D+BmPx9wzRCCDCP68TXl6LcV6PT8lB7BtCqcB5DG+Rd
IZgWBFQlCjSr7cHFqGII8YfiayWdnDmBLFpfMwCUK25MB6PoUI4=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
NHm4neI2xwxIlCb+cFEwXb00otQFEKfta8soGy4aO7V6XQEl2IerJzAXabM7
d81roeRoBQviXOCAn5O7nmHpeNWVAi3qp/g2Q5Dy6OPxPkLwiJCwSTuujCOQ
89XXt7XC1LiYelX8hcxGjMA5G/0UrQyenkeRGAniC8kbDbtOU7A728V7NgkP
g2Tkn34QmZIW2qJeJ0o3KexN7pKrMcPk0qAGzy5ZUIucyHQ+nbWcMpcxj9GB
sTguEVfyg2DCKLRQjH8ObLSc7Y0dcDXYBn8cS/1U2cBPVPSMICYDZyCjc9Ps
Tpcf02acouimRyCeZYtqJD7wIthMPB2rwxq2ofOqhLPAQCNklAKRVwNO4bZp
Ox+UB4oYn1LiSqVVifUXUvx7a2eakcJsDGfjqZoAVmPvWgnFNOQSz2ASJuUB
7JLgkSs5QaigFKCBJ1r52ZAKAuzMLifbLfyRGvsAtmYnZw17pj3r0pVXECmE
EhmDOar80Ana5cXNGsbXxfmFlESYlEI+


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
kmGNsELZ25vPJdPNzBzSJd5ElHeUS53QQh3Q+LdkrrSQS1dTjIArfDx973/K
ovbcrwetdPqwaD7574f1Xt0E8oOPSNqBMjj7E2EwOLLb5VHOGRXrG2V6NunL
UDA63e3OPhqTCQhcRbJkf04zK1R8N7UTecIHj3Nv7luk3ko6h7A=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
jwbCV1NiMVDAESpYccvZGg2IVxdB0e6Jr7A/ihnEk6JoJSoi+PQnlvx8aOq3
9YrDQUGwnADkBZznQLhqfobysassFmP4eTg2Mt3S1nCbc6bI7k4HYtpnDPlI
BV8tfmxqJ3IKATJzF4iW30wa/V4NZxyv+NWx9I6hZljraTM5sUU=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 176544)
`pragma protect data_block
W5PBcGgyhpch5xHoTVG4w2Dy7gRWYiYYH8ZUdKMzAFKNJd4kcRWu16l5M302
v5X1ROAZD9vuDyuWhaOxPM93+KpnWEons+5qPvCZD36dtBVGZ0v/TSWT2rtF
V5tswP0n81+I7VYsNW4vDZkaDIVtBzi1fG9LBmlBOpID+rEmjwLISWXrBDPu
ptm73DMNkyHhVCa5pqjIFIWLMBJo5yhNqou7O4t0wkXerbYeZV/B8fjRzR27
Sv4qzf812xbbT5qm8kcHo2CUJEFIY3nJfkJNu8Yn/Gs5N5+TQ9+RLAqQSvRC
KT5bk/tJVfJ99eBsxrlu10i0Wc18eAZt2vz7x5oNzVWWMzQma4fJuZAX6TgC
jA8ODVRMV3UQA78D2r4eCgkOi1E/qxzZaL131mzoxXJhXM4ECxn2Sa1neBeQ
EwCbgbKtLyEeD9vnylnviLP8kPWwFTbOUJW4hR7muEbxil0TJF/uoF1PZfpU
bqwQKusg2hitnReYR65VIo2AZpOosSc0muQetp/+Qcb6Xg9ATDaDHrc6R519
Z7fvQjeIODwHqLD926JMT6Wey0lV32CkLF5Ls8Wwka3FMWQLyYnKGpGRi3hR
NhKCrZvUcyByp9v7K/c/ShPcAMIuKlxoyEpF5W9wp0KBoH0zDUkhIOcbOy2s
TGCT8LiApYky1hov5Dy4Iyr2xs1cErkr9YK+mwla0HRiT4kCMnVV1iVK7Jtz
/rc/leM6dKWBvvdxKpDLPeDAgaLLgMBWaVS9JN6yLXQWfhXLrYADYbmmi+bk
PANiTkaxG865oJj92Dqp2Is3XY0etXSLSPyDjQZbIblBLDKivQpzBp3cDrfB
ASGtoVEQ0SzzZtN8SsVqdo4zQ7yFrkGhTGM39lgFNeds7GA6OvHk8WeBiQoN
f8FjI57exTTmzNZ0S7Hme/ZyuZ9usjVej/99LJjnqBWcjIqodXwsd8/d94bf
qPpXHTQDPT1Om4/qNekPyc2FKxiqberqCksqFKqaq9Nj0NMDN7WrIECI9Cgo
5/Fljr4yqFmlWsSuRKqaSQ06vGIu3RAK0TqCIhxPe5MImoMY1H0VVcumzbrf
Hyashv9OVJrIq3nVhMzHvRHDIRDUAkqlRX7zwT8G5xF1F0pLuHmEFiJgL4Ue
fexIbyUiiXNCjGk1hJnbtE+68JW8J+d/gxXEhDHgOMU14QsNXov0ZBKjU/EH
XOMuvh3+KZq8RiniYKmEjL5B+PZVt9Idiw8FYbM6miLxRCrmVqMif3/0u3WN
sMQ131/ks6ZUCnmdzZikTbjSOhyZNh3B+mHym5wtRW8J3uuhD1inOeGrtZTc
ea5sNcjP//2JTib1RavNEyaN4NnTIeK60drNQBaq8yLFUm8Lt47EP97q6Gbk
YJNfKJ3IkMahUuX43FiAvPdAIvTopbU4xa1665hZU6vfD9/KNuoagjg/PEVR
dcQpCkv755hBx6hWgpDXT7xI9YPel2vhEAeqx01+OtpWqfbQ9Fw3bmXdsAF6
KuOmJkVzc1S4VeYod1E25CwimJFHiYsogpiig3u7cFF61qw+V5PIRq9AqQ41
+qK4YoPSGiVPh0KYjMoxR19uikncrnTwg5E3sqaUblIVsNozodszQ31UQqcM
6Td5UbBBXOPY99m0l2K3Y4OtJlDiAl47soO+EdRp5kPpB+V9L1jrpuShMTrH
F1ejBZr0r3E09+LmTmvCg9zAyMRo+ph1AIfySDT8xWF8eThCYYpFqpiTNQ4V
koYlDo1rEQSk/2QSgrOhlynCK6SOeKhHzIFLCNHykEwzYXA2DTOPqZMWkC4q
o5cz5Pb6XcoQ0CfqyjxlyFZHB7W4sanVMHKWgdm56he7Xipsv0+1PV1jd89D
frUt9Y/nChR8y70xBfW4pI7+HAJ1lSmcHeTWFQLbWNHJ6gI4cGvXITM6L5jE
waMdi63c5rOO/az8jtmh6XTWOpcVIP0HU94GyNp8TpNrW0p0A4AIb2I5c3kN
tt0rdL0KWMPoH20CnFY5DJA+uD8vM8Ebe79Cghn83GVqgWBmUKNt8wGhf8Qs
ML5qpNnl+3N3/QLaSPhLgY75swKtkgw9ZZfglqD0lexciAqxrfAsoGS3aVMH
MkJ6qWi/H0aibT/uNVZ9EvNv1gGR/CqSkEh3XdpqKQuZzhvSBHNip9+u7PXl
sOCkCeJg1gZqFQHq8hYiJDYcRAHHdpGK0QG9vYfGoxCNt08CIlK8J9RcMCf+
IhrGXQkJzaA+gkPVjydIFQCRo8z4N/TY8g51npBptAcZoOlE3oKKIqp9NVoV
X/do2IoDNKP+ZrIxVE4LYTmqUdOt0GDH7yk0JODFWLbDQYhQ2BgKQ+rnLXNe
5p6t7YF3kw8REWOUt12NPwgYrRC6yZ9AKiUiQneU+A3qYufPde4cHODjtK35
LmEZnF3DiL6exHUV5wkni83nMaoanzDu13Q/3ofrmM6fb10AcSs7QA0bZzqy
lpNtA4hP8z4Bib7edNbMDc+XxnJNuRM30BKz946dZ8q41vkJCMplnPwwijO7
+IqyXpt3kSsVIp7gnrVj5T90EGuwgF7GGa2fFTT2PNsg46rv5rMUk/LXTc8X
lbPoyZya0ECiyBvqh0M0LWroblDpHmOKYKgtIpcj9zHduYfhVt89kAa8rSkE
XLFQ1BsWYd35KgHrwDRiF329Rm5bYV7gsGx6qcRRItOxL/3inMbpOtQ9eHfe
793Nws8dTeutE93/+lX6DdGrj7AInXqlow3+zxnkmL0RD+XSNecmWGENBr6b
+4cUTM1DpkGkeFoH14CGhA4w/aG8KBkTERfjTSygeN5L9d/+2+FNx45kduBV
HG+pPUAd3FS5wEfeWr3NPyUw0GPdMEZO0TCIPacXIHHLzpeUs8zEZvSSJbZ1
AaouBqWB4WD/EO5Gb6VXWkWQLk9FyL1AOlwWAyi6JAm2y2k+I3L1Y2XCSoAC
w+p9p4/pCJeqUJ3cYk3Frl4YxUVUsOtL+RpP5w1DWNILHxM3GlxnPCmTQK3v
i/27isN3BItk0AQVj7rbnjW1xI64FReLye0DlcnqIu+c/5NQnx6F/e3CvI0J
8S2LPf5/4sHo/au2Jth+MV/UT0L0Yq/pshsGvZhCZEJylLocm23jfPVqXwCh
F6XAcd6acZSyv++WRV1622VWgywbGVKwGziCi/NwR7B6/wWCMNjBTbTA7nBM
AxIlyLeTlj1ecCIa9ostm+lQPhHWhSKWvsM3mYtZAevAH5mvSh7uuMbm9yJV
DXMjcetegRj+Ck9ojQ1YBlsFedNqfWVh4MB/Q7XYn3FdWsCiN6+/Dcd0vNnD
OJRbWjHbCU88SZR5bO+KAHMCNhnI/EfdLwt+hzwbusRoSD8BDb43C4tengAd
8ETT5hq8T+r7lHG3zgNjH578ohzybsHO1GK9mbqRpkOmiYtp+cs+qJiiBATl
hwpb89D9yhWsjjmzX819UFHjkofaTCxs3+edTyqhUZpmZI6b+aFs6KhEKYfM
u8GaZT6H5rilL8+Fxrrmf0fph08Q3pEBWAB15m2AWagSfY0uHjFgpC4Sm8sX
Zg4OgTfRmEQyzEEo0XFf27TYurA2uDU1TqC7uZXT+Vy+n6DUkXaxUxQv+cPs
lKVPrXxQ2yUp31IPUOGlJ0DYtoNiknAjDEckeLOWCvMccV7SPe1ubgCqpoxc
/+GB8xEJC4ZmdkrO1+d9JbLMSERRdB3wJcyR3mam3lwEsjnXT3hU5P1qvQiG
TK48ocHhX7lgWnbP1iVl0+aHxw8rJcQbULF1aIPcZH1j1IOlnL4Au5lrVcC8
sf7mGqp4BlL95YBNJbx0DDKdPZAYaLLRSNfS4pS4bxAnIlKd5vlqmHuOnDzI
WGxcJCeZ6e5wyFobIHvhp5dEDnFz60d5r9tY21WoQ/UAX4XR+G2+4YaWAEYW
9WKs10NIDpXZRr86BX+vZ2TBfWuFDvzSwB3SrU6xpD9Oy1F1zxFpIG7Eed/J
rd4TwJWv3FcgzLDznzIsrqaCsnmMkQpDRWdSbXsLARxHRtASJgAl7livVr4M
xhHMMk4tYLDPSLLVVsFdDdM/hX2ivUbyILuPLPmCfS9w/6Z6sLaOQfiRjQmo
bigxVy4/lGxkwIwlSnPTDQf3RMmaQsboTeWLQ28ZODGiE0rE7srweKHVnkPv
yLGqaCwkCjGTYrLJCzVg4q+B8szD+J+u5U5IOKBBDPmYSyWCJJ3tfTBLdI/c
FzBPwbw6mBmsYCbnyyqlIrgjsoKiYW3rRzciqVQn9AXoQ6aceL32ViT+P/IZ
uJuw0wSoR9+Ce/QEunQHfGOpQ1VgPBgXEdYCnOkF+UkzfKl9UVj1x6amtqVq
qVJ+oeM5aaBQ9ked0qtbFsuuGJ71nPKGI4aJwXggJEYtbGL0akr0HcDupjm3
/ssLiiisLCQ06ei8dJINmQSKOa8hlCoKztmpw33lV08W4225DgV+M1npVTA/
Ih78UuMooXQ61TEAKttASEv6z83oqqJ9+XiOcRBaSlQrhBpvCVKHRmEYI7b1
H66Gf9i1ZRDtD3qIsWrmT4XubxpKDRFiR7r07+9fCDLeTWQNZI54X3XYSHNH
OSLoJEHDyAYD7g84k7bBjoHXY8Yj1EdHdguc81gP+aT9GrFzQJT3+PoqKEc0
PpGq8uGUWzGR9UnXb8CCTEbgoX/6+CHEVcrgXraFq781jn4lBQR1pW1Ivxon
DZwnHSJm+getsb+I9R1IjLNBL+pQ17I+9b5e1rxuTun29O1UQ9EEa4di7Yip
v9y20xDhEyNy286/6GUTQUMTQOxtFgPhbxBcXudqCgL+CcCs2fwurK+7SjE4
XkWI0LwQUA24L1k4+ZAWuazt1h1bIPOxuWE7Ur8c0MAEjgBX8PtZdkVn7duP
DNz3WyzV7qUckzpE58pCUZRtBveZDfWzPv528oVR+nMVGBgwjIvym45gyNJB
t3QL8JchXgX3QRIkWsE8NGpC1ZrstjHgYGXuzeLom8WdUNgOQ8GiLTyLSJjO
b5Y6jFF0wIzX3jx3eZ9nCPKglhLxiUgBuzLqerMIxwuq3fF1bhvaxwA9eXUc
tnIFguuhk5KgE+ROMd0WEDcTait48/mZ0dgTNEBlfLrARRDtmQ77g/pbxEjn
ciyr5zJQEVpVLwJcHHqNQc4wOwjc8Vl0EjB73RlZiNjgEvXUkfeGtvhHHqpd
O5mlkYXMGrRj82aHOG1KSIN09n/T8rYOt0+/C/ilaDOdi8s/EB/D85g2vU69
HUnp9qg5ZmJ9pHHCUmtdTWxQ3G4X5Svi+CbfoWAXrYXuznHRU4sGs3LmNlO6
/wc9T9hi8yd37LrrNsINcXkxxAkPSRh6cHz9FyTJgatOT/aCoNBjdB/efH1u
aqqgLs1bEUyeMxKmXtNjoG0jnyrtJAarT8XX8EYMy9Qwz6CtuSUFbE+AOtaj
B4+IiUqf9uMVkAtVNb66hIHK5ElZfRUpLqidpz0jtlLYARjlGFPVTkR2ddlS
NaXTuLD0xTT6wZ9B/Fac2oyX9S0zWvW4H5zz8Z3vN4yIOLBWdtgmH5I0/li6
kT/8wbao1iaMJcWx7iLmKPOHb+C9zqWb62LCoPLEMe0xuhuhhWz/saSmM7Ca
H5JR6BIRBFOBjD9yhCobIOGAWqfvOFZ2FKXtYMcqWfX/s3UYluAQH7oIZEO7
6sG1TP+ZpkstoZJUrrNBFalsHFb9y+cjxP6zvzL1tNlIPqwti1AeWhoCTiA/
KkumaewldGAexSVZ7VkTvCTT0hfyNMjXHULP6pSHGyGwvTf2Eg8HZZSHIT4q
gx+PJJRLdzVk8yE8zv9T8miYmJAM4V2zm3Zkg1V8qFFx+OgvpJrttuSMXf7o
6fSfrpVtH/wI1Ohs+o5RNCh0mKW31VTm4hB/D74WHS/FVLTrBwcw/tIxKO3k
5TtMjBrf4XwhLivdxEcWz3tvcCI+XlVXyDDGN7ER49bONuE5Q99fFAxHlmOW
cqoZDeDD+kHW05B8DImG3AQvMsQnJI/szkM0Dv0RYgGHmOGuTbez9Fzrhcsi
xKpLonQVHaeA1RwGZ3aDXRsb2jVwLg6yytJbV4zuIS6WHNLr4pUUK52lV1wF
hd0VOUM/4gzO2YbOAxTHxf501xu5LO8BVTgljErQ07/4cVnvMFk7F5ebaSJe
EecuOpHwbyhVBEjtxsBwaS7tlM22qQiHvo7vz3iChiMkMEqJZlvPJ9EPtgfI
e+Opyq/l30Pvi+Msgde1Wv5s+meNY8kPsHUBGQMo92vFVA0i3UFZ1/WDkwj3
QjaeMdoeV5FK59caJeJza4fA4Y5V+S7wTcdZNBSiU27WOhrx52lEPO/e3FwM
7zkVrX1JVefkOCiyDJLd6afjGKcGnLnAwRrRA+hqdTnsx9p0MGHyWJ3Q5n+z
FCjaKz4jaANLQlDYdtEghW3GuEoVefJ2eK0CZAaRXeHhO+F7Tvmnh/UQRhki
LK1F821uFhCM4YrzPRQhl8jWzgE02lpKhcy1MHYpIU4/rlNezgOIKrST8/Mb
1oa9CqpY1sqz5E6T2D9DN+TJ9KRmCYeKtEF521w1Gw853pNqfzZ2zuKV1hHQ
DoMuEwIyny5is24Kfv/ymTSYqWWcGgwnzyJbiWUMsGz3exQuxUF22Rh0cPE9
MT3VuA2/FfjF2ClQ053Y8hwbSmXB4y8t5nt9m9zi4g3xanUh5G7Z3QAcDJWb
jGRgS1sN8hpnZHTcLzadebDbpqMBjtl9jWJ5w5dP8Yar3qa6k2UsRGGInTcE
mvw5ai7B7PJVKHlR7spuwJo4BRd3efuz1iQFT0zYHo7tyU90EMiKCvjghY35
j6fpqBEerL+RX0OO9sDKGgRCGG8eu6OE4YLtbD7DmQVhCimGa5mVzfeJGZNR
Al7HZ3yxsY5gpHvjb/YhfE1hObpEYs97zbjg2DRS6C/sgzx4TFD3cDeuh2Bl
Sza/iyqIvwQkfdccX/0kpXggHBHhlxcdI5gg0UD8g7Ln/55IzBD9SvkQnq39
PyTevf+eahj8bb7kBEdP0zdQUJuskNXmtUHi7EpE84p/LDL7mmZZ4cT9xmDa
JMmQ7BXFbHJw/JuyGjS7bb/fxiFwk8uN4ffq2k0YtL2xTqEVowMsrTE1qGBO
0FXjDjo5rZNabz0nRGuJSXHSck98UigWTUObHpwNOEVkPge8u06htXzCTqit
75ZX79Eub9Y5XDRBc5pbKF9lfHrN2ZtoGJkGMRGXYkfl1dqvnMRzwmbkpFnO
Uud515osJpJo6s1Jxi3ejXNsV8RGdaYV+klkARvA7pbN9cxmPuLZjfAFsdvA
XcJ++g6TD6jLStTgOkdfPXx9eGU6FCDTWcmucyn4Oh4avuYDgeZyu3868xWK
RSmG9HNw1Hacihqa4ESkY+SyEBO2h7ScSL37BLRllsA2gc1Ouoko27N+gX5R
tBJ8+X8srw8ziVyPimuYrb/q8cq3SX8DOmtHf5CslJ9NiGvkIag/OZM1n14V
XH42EVFFmW3hMIzNeaLfsOH/DRNrMIeHFLhxbPDn9G6XqEEVWEm1VxVLWqmN
a3hM4v2UzOHy+lQJW0+viueke5Z1FV0WPkhx2B9g7FfN737JlQL87hBg65B+
FLSNXXKMgoVMWif68JOwMBi53rRHw5cG/h8PtUJ3u87lCPwRn8Gw8/2G5uWa
b2zmj2OJa6MlI4eO0BEvRKkWUi3fOUvT5dm9/Pirg979iBMx5zTr9xEbd3VT
rwCrsboQp+Jv3JqPQjwCN5y0aEcENU3Fm5N6dvURx1ezliswiXKuBnI6U6Kn
lQu/Hp9+JtHwxk2RPls9pqW1hMRDqS42VBo/te49JxODhPZJAXT848+vounc
oTYzRe67kvu5ctziJ2vK+Au2IHm9s3RJRkf/cirt99We7184/mdywi9K8lTO
ZrEOGfGWGJw3EuqckfDaGJSSUd6g6ROQAyTz62rx0bEXx0x/pOO1a1g5Ih04
c24FktXPFIGOD5LFss/dcR2gKaW4E8gC9R94MvgL6PUWRP2GaOUKMGIXaNxC
N2hQL/50IsNFUW50pY5liGLncR+4jz6fSTQDEo65XC/vnLRGB1I5PEQ4s3UV
zkHaxEVln7jOx6n3sPRM5iB0rzxAjngZU+IlA1xnMIYJMacwWWaTDH/7XsEg
a/flfXDgXyfZUIz97A4XvYIQRVZY4mXW9QrK7H5oSxZVq7TjBeHvq7xw1wop
Vpb77emULnsc3W2af/KYFgsreD07kT01ZuCLoCOEXsjwhBcpsgxGNx70/ZX8
bBivWNc8yWiTygXMfGar0vHVFIKID5TxEhPu0RyITQ5+Ni7j0QGKwEoltrto
efL1qBLQ6dO8+SXUHn6N336dDZwd52X2Qd+pgwFynG00/6GYjIeflVSs+LZN
x3QJqtlTen5V+XQH0DHDKjc13yTMgPi5DVVLduNJNcjG0bMWvoEma0pYGjXE
Z2+YwqBBNp3TLbmSeQjfaIIlsFWQy9f+7HwxYNVHAjHDe9hom+PZS/VHKD1L
Ft1nxPGviSR03RCUOhYqVFThtNmZR02ihKu5hrcVSanY9wcZwpT6DfqOnWhh
EA6pFBQ+vG0toi1AbyMsseB3spUtsALnt5/RJcdXTwo3a+7Hej0ko4xRIsyi
1quwanyK26xcQgOjF2pypjPbbgVjloae8N/jhfU7+KM7yFa1LEvDsHY50Mqp
vsiCPIZQia2hCpJ5S/pbmK0suGNMt7o+xp/a97qJH7krR+0Bihy8s6vBkyWo
RGJVyoeW3MDG2Q8axnWRyjYnnPafs+y/V0UaQYHvNLzFRnK+Yz0ooA5uL6Qj
U6Mv/nEW0hH+/ukQMi7B1GF2Y0Aq/i97fjRm9F90xgaMlRjhJlqFLDMIYeXb
COXVbJZU1fB5Nw0OD86cf/KbyOqa8wFBWoGWRFBIj1hbpRnZKmyp5i1s55wK
nPBgs7xJsHgE6yr7HjwIU7U5pTHDWRnF403+FM6UJpFrq5X+VsqhlDffEYqN
YvxXh6y/79W21ZvxWdljxc6MUktRpHjA3ZcnVzBsrYWS/s+oA7c3JbWAsMfn
Dsp7CbLkXrESXNv/GQ/i9cp3G4B7Rmdb2j0ah2TsGqbWNUgZDoUa/msTFwcL
TaUM+ADrEl67Hi4SN//uMqtX/fJexdpyHWPZrYVML0IKq4voiurpsA6eG5Qs
AA5+ukDmu8/mbkXf4/A7R2bKvftJ2grVfVFfHW5uuBMrgugOiV1Z7WMR1bNu
MPja+mPfZqzBt116zacwCKsYb0AqeWBw77TxZBXGMUwNqGS3MMIhPAYlfQZ/
2ytBryHVQAj0jyuzJ78D1MC0A/GWNQaMG/wdtDFROzDZw7nDeRSyoz2d8Urz
SA+TG/j3Op3PaFpPsExzjcwD5msC/i0PqtqB7HOAZRQ9RdWZqsB9h0+d0zAV
P/eJXGSeXiSijq0CEGb6JvRAvJG+7eD2Ii6ERUJrHqqJmd+dYnRIXsSKwBzS
jLyHA0UgoVjAIoO3Wm0SjAzQAKtU7u39h6SQQsGK1lbXTIaBU/LFv99+VmHC
8yST96nadQLPN+jNLQpNqdl/dHJmuJO8thJDDfMG4g7GwM1kgLlyKegtXLKs
bu8hSXi0/w2/k1bs/BDTPAqegWJL0V6hA5AF9byzumlhM35K9Eb/x+UtdF9X
F1xIoAt/oGU+omNZTMQyK7qmCYRhP4VD5QF6eycSaM4/7wIgT2L4Ipd+ELXm
8ZDOU3pBGgZClr9XfKupz4aY/4wYT3s5wvOKKyqI4tSX4Yzzdl66yx/YGCTg
pP18amwLIaTDWKJGLAUfX5Aq99IhTDl51kQAYi3m3RTiQORuU+MM0fVyHrRt
vR4XmdJf2btOENbpObuNdG8vCQYgpFEfPyEXBIMuRNVF7m1+H6NRti2+dGvs
xe98A7T7L6gL7EjV0Lo62jUHFK3pBUO7UQl8j0n9ju/hxI2wlXNQVkPWXm5z
0tSMWzR1LrRxdiZHJX6DAZKs/eRycV+HCtKYCzOMrHtUhSitJlHfcr+gGytt
pSr4WYKngW0OZN2nGmkqrAWutCwlY1ylIYJxU3mNxjgaIkPDk4W5+Y4CBKKY
ukhSn9nrMcxDb4Jbhyo3q4f4MAu30txz6O1vhjpdKryxiB3cmxWAkNV0rqob
fv8u+RgtTu9nonUzD11iWHgB+xtQV//j+qlIqYdbwXGdNlCbz4qWTMC0HMdZ
tPvVRTfagBJ7LO1kCitviA1y6M5N9IQuvU25+FKUFHta2b2aJ7updydbr4e/
1lli2xtS9SjeY4yLS5wEdpRmLcmG3YsY7dSyHoEzr9+kt1k6079WOBbU/u8y
YrofI2PfDjlObai7/FiA6X4Z+35Gr4alzVqGVkG7HGCPcS2wIVKsWBARj7y8
ldV/MwaG8VpSFFHNsnKxaSvkXw4kceZgNVROIBGUNn+tz2zG7a1IeBRi7Xbp
uHBJ3U3hwl7mymeR19HFnzz+LspUCJNY/ytQ6+jMopDJC+OhV22U/Bj+/d0i
qzj1HoTIkrQlTLV38qJXwTbakkQcqi4DGhlw1YhGQUDyuqNH0N2yxte5U1bL
Yspv3HPweSH0rc49z5iBJB0hQizYh3anSbSldrV3y3FIDmBu8CivkVfbWL4U
Q2O4J3oE28Px55NTt4GOrHXiiJW7+phlH9ZRYuqYjBoEDKb6aPMNdq3fRDcl
shl6nltlNWmLKaxv6GL9NFWz2OH1z8QnMHRpLhOOaU8v8E2dTKEQVjkEX/MV
LbL/wx+0YL7JG44ttO9PeTQQRcE47qnEM7Zh0K+bgkkdgK5nO/IJ7gmeYG+w
i7KLULB+J89fCv6h5WoUgMA4LkYPADopxH1a5CnIneSrBsK772aJXTyKPA10
YAlgHdM1A2JG6bG6gPP/nN5guMM3F6IOGT0+Z7dOEMSO1sDRzdrKRyL4H5tx
2KAxwimeP3PycsOZZ1mKmrNpsLLrKrmZkcDTrY3VgFoHnqrcTe9NI0wKOavk
mm0SLePu3IbR7QwWqLUmNKjo/sBXqbUZwj7IYnmcLue43XsCVUdKyZuONMoW
VyXwlHZI4OUvSFB/oHj01RgCvSiO+hmM+oCYzhACi/SbBF9G8lFhW9jS2beh
rUrDQqyZ7lRefv3DS/i70ToYl2m9P5UDO6vKsruujd6sURED+pXyM9dJiNhR
yjrMwu871TxRXtRVmpAW8yOzIOjhlokzsLvz7xhkiOjg8Nzfqp1ZMCrJurvo
KdL0Hakf9D00n+VaerN6bLPMQbgtquWNQv4X01Ef0wE5GWfroskLE+v5je/F
+a3+vZDGaMQyntHZjdZWzIFMxkagUA95SwNNvdh28KfX8kZ6GgKCULQq2bt2
cCBk7323bQgGCskHrspZflYhCTI1Bi01cHVV68nnHLr402PgL5hVwQpYppZY
2n98KUx1tFLIpT6nVZpKqdMDMhs2yyZAaUwx4BFIITRd332N61xffYJjtVt8
We1HCWtT7Vt8dtKGbDN3I/P3yiTBBybGt8dMlHB2S0tbqyElonl/VMJBNR4y
Y5i3LXpjQ8Sz9yR6kcy8+n1UhxozkdIGnsPW9rX7r0nzNLc1t06YQsJu0GMi
W3yKnj6aiBmd14+pLYw++Yogu2Sd9svlIRHBnVu0J/QVz6Eqf9xm1pJTntEv
3w5UBk7GNJ1c+wX1gx4GqzK5fQadeAtZ5xyCIqo5TTfP996cS0jsgzbwvT68
3Xp6rQGlMhAWsrldZ1u4CmT8fIpz4mMX2Ax71NxDG3649EvZi9JNAL10Zp6N
zQXSEwLcaTeCrXTdf7c3A2OU626sCX4XzKLPP9X/ghGkVUqGH4fVS5BLkLo+
PxWMP63VvBOoaHUWNyd4jJNAr9DXaXniBihd/6Fj0IwxqupQAqRjlZiMOs/q
uHhl2Xib+2eSaVgcLw3uqyBraR+j3mSzKKdGe/fFaOoiytYHTjE8ObjgZrob
Nc/9nbyKfzjFh5eGaXLwib5z7Gm0envgk0Wm6OMRGheW3iCQlJ2JDpmb6lcc
d+CZoxkDtKjF+pNx9zNnfJXy0T+fSG5QwyFV8Qadp3BMB/M04DW4mOwXdv0p
m37XRA3rSsKBX7j6ijSnihRQuYs9NnctipcPJ+eZ7iwYD5HQEl6428FbgOVN
64DMuxRmy0k0CGsGiSPFMhqKE/UA350wHnTZKtZwACp8pfI4e95pHyzr2Y30
Rgwku2bjdSPJBA4Ak89Rlv124vaeDztfTIeZdNckN+n6jvmW+jL9kPohyaDl
PQ0JHWWaqF9P4VAmyjCKG4scCAL58QOgi5/aPxhX3rbRdf3kAM4n+MZyUKYL
U35liQPks5+vUWPkYuUnut2LB0T9EPVdk75sR9I1LG04zDyXyQodk95Mfxhz
c5GlSXC6J62o5bKoQcE8flt4uhRKvO6GPK6/2QyQqaNOigIWl2w9JydVg2P4
GZJWY5tAyV9wSD0XgEB+i1hEmDKGAkLaUfykyJVJIfdIdp5s4VGAo1I6DIuF
2vH2mOVth2DA7pTfxD1mew8ni48Ov89lWKABKx4m8RPwDiHfjnzJ4fX/90ti
OfVpHrEcp4s0fZUvDCVN0//j9QZlSMPYbc/V93Y+aZ2eAAPOldjPhqM35HDB
vhNXr8C36OKG2s/h3VT4auf4BTEgrIi2jdXuGJ5obmdoRKMSz2+xcUQWFbW4
XWheQEnSlTfTLEM/v5bTjnLUi9JNUJ0a12m90TuyQsP3kHk+y64VJ4ztz+Ld
IgsFfmjYurMIiGZnP9+DV1dKpgcTt50zmHp5+l0CotICFK6v+GoSyQipOCdj
1u0DgiNJ/PD/tquiWgi6MgNPDntP5HSMr4t37ONlTxTu+03d4yWVHW+XJ8pP
4pdnpb5qhJ25WXWUfIQWPNWuc1CTu5EulokKPSxQoRuNg1uEL0Nt9GY7qVUo
L9dk9MXDztx+kxzjIf2tRv4M8ItOAf8Zc4+oqojqKgEIjXH+axf2e0qCSj5n
5DkDJo+k00kEfFtDQlRPOLi8WJr1aujYnexoRdLzhpUXp52Z5u/d1tQr6Doq
DIo7wOrnynvSSAe02QzC5nuXscsXimGfTOFeeLXbsf1zgiYQv9cvztpc3zpO
qhUPc+jtJdFUgWca1lBSztdpqG7Bfthb0krIuhEzvzyD6IkEMa0KQc+9ZvD9
FM3na//IbXgAjXdFQnQEt90fNvNrNzaryqtwthH8nOxv8zyWq/JRhuHu0ASe
49uvuUr74rohfEYca666gVshAlzEe+V6pJG1hzgHd8kLoJHNMqqWMKAUnXnL
KxMy1T3iyxp5aaPAhx6hR2N80EXD+Al5V6oFNvgZE6AjPw8BxzcKNrcqZM8F
Jbe6e2Z38x8YspW4ywN2ElFc+nFdWeimNXbbNTIM2HOS9usNTSC3vLukXK0N
CvaQYdOyEgrMCyp8xlF5hkVPnJkw8kQzNCgjwD2zBjznTdXy9OEBXLWKlhch
JE4GKipb5F3jjRiMn2s03z6wW/r4plzr41ceRCvUwJsQ2rGP3qjdWCx1rRzn
lLskYBTpQp1kqqxRP2TKj8s35hcTwjIwV2K/guF68QalhR/Mww1T8icYyGb6
UE7kyIUzTE84Bmfjduilx8Yx3+no6B3Cn32OGS/UZ9IgjSoWMscItCT8A5Wc
NZTHGCbcWXRSiajNIF58V3PlRUXG02jbzgCyjOTBLawVZ1ZvDuGQ5h6yE7A2
l3RTanE36W0qNwZWeKQQVGte4BJ6qaEGo2cIx6o4odIqJIhdJQFPSIF3yRIL
2WkevWsVTvcXIOFL1I5i1sFpjBC3LTx+x/lO8A7RHOS0oravAwsG5/8H/uoM
3I9yAyiJ+JXQ8Jb0paRryoz+3kOC6X8YFCDgbswJkyggKrRQpFdWwIrdTcvW
riEAoIKFdliEG7ijW6jvarwGxMkOlgpzbsXVIr6yBBRZk0nud62zT+SD6q5E
zozyZbWKHbooGAOHeOEQdiweexLJ1lZG1vBk/s+XoD99apeKtJN/vLmhcH/e
s0L4iFgEqRHd+8IUrlx74NU6Q3Y+zOdgMXwm+/bLT55RKrgjXtXvTCLclYC4
C3/MyNjSrDCUXMrZ9aDvJMjrV6CI4DSTOVoBGHhL1r9dn6qqNbN4b7ZTMnDK
hikp9wNetSx3tnslj/nQFi6OthHXs5OfgCi5RmOx5/rkpiMrr/Ua1+7xs8wP
sM5xmaYElkr4yvXwFerp+ftxrNq5pByY59qvoB/DP1I2wHsVAGX5HLtC6D/t
3sIxU7aFsqqMMn9ocn47nb00oN3Hd4nymmFXuSfXqwOqV+r8sfwveVqi/W0B
g1Uqp6DYW4hLNAE8AjMlY8kdPgGUscizRGrW+pVtL8WJakQQLvHRXZNRdAcn
zBK/KrIBWNJtaJhDh3MTF+MlngS/jzAfqYrELdboRAx6qTZFD1Zs/eU4re7g
wH38WfOkW9mVJw9I9F9sX4TQ0i3uimfr1Hq1IuIedgYBjnPI7EX3laOn/Hdg
tZLl1Y+VeIPTu3SkF05Vqup1RWWqZ2auzHwDWTgzWMTjn3pzl2cv+q8UZNjI
cjaurIG9GAdHU1ujd/1UGGP5JuSunvCmy79MipbIOu0K8JLImZuZBaaJd9LN
xH+Z5fB4qDmO/Tu+CHm6LNs3ilOHmQBrJUoy4ZY2epx+dJIWVNYLZ7LjNdIV
7Fk/5B9wm3ceDQqPte/CsAEdWJDK3fR1MPEceD+uyg3esL+VaW4qyA4v2G+M
ZFqAbQlreWTx9YJHTXTu3SYnlh7VE7KHAaMXeQMqQ2bNd4iQ1qtXKl8x6gFM
/JoQ2JX28bsX5W1wX9X4IlwSpK3pxTo535gumWdW/9eWu8u4SvxJLQmum4wW
T0th1lgQPHaBPQPDKLsw7KXRQLus1UWrENqzWqQ54k2pLn2hwAcdwbBAjmeg
yfDrr/C3AAAebyltWLhuoPFBUApxKss/UGovbrl2NFz/9vJtcme4QvPXPKlu
behllGyO9okbuIMKnfCv0bXKmPBwhJW7TtVtbWVFgugpnj3JibFQoGGzP315
1zMJsotNNpZyEONC8zHkbS7vWH7KbBA77sVRzDdXoGyCiaal2xVycSQaqqzK
2w/rrOwBd6PaRF1qqa7q6sDxhCjsWpPyp71uKTxtaueppWMk/IZWYuwyf2b3
uSa8UO5S0Lcvsp75trYOtBVdHr3N6qxgjbv1hnwMh+59ioJMl8ifpu4pIeHZ
VVc+CFR86lkuWrX62Nql0vDuZLsNi5Ssj6nqFVRlPQht8gJJHy/mDJzFi5bo
4U0Nfo4foLXZpSZkGiSVc0nePHom4Zuf/9lhwnIirf1TUX2bJH4RDy2YrKc2
dhjsG08y/1rbfy/dEzPrD2XviIYQK8rJunpkKSyyu1TtzqGqeTlYYALU137X
YBYEr5Qxw6L+Tus3KEitrTFGbl8ahJhalxJshA7iN/IA0Z+QPQmCfv1asjCu
0m9nqCxWB/1GLWwQH36bF5vC5/28+qbcA1dE5dAVJyzVA+2J6jjaG0AC8uN4
x0ybqvTVv/oob8N05hiqevOpbmVyVj2prp12Kg6Hg+1Pw7U6W3E+ZAmPeekR
3yQYOV5Z+dCTm6QnkjczmMPJy2+gv9UXvqDvmtiLYXa6f8fhfkSdrHNsDRBq
mMd35djWxw1Gv4Zwcvuo0fnOEdzA+Bp8NxjXORZgbIdbnXdrpsei2XNvveON
ZWChCzXbLVPa6eR2gr93WF9PnyoY6FbwxbZ+/JmXe0+2v4CARqksl1JiqTAH
MfWukZqdH3g7LZFmNxQT3r6ysSCW8me69ZGk0vmOf0zGWF4lmfXHOV3EFdV3
1Ogt0M26aMHuw8Hk9dbFsH9a3Srbl3mFJKpyoy3LqQPGOsvvJbuFocLq1AcZ
vFdiy130JI9NCVyQbXUC4Sp4SZCxDaJ15az5y9FfP5ZfxVSV8vEDD47JZ8Xd
uZd8Yh5QlpCBt+AXrpgbMvMXRQwmdtNJE3E2C2v+MryfWxy3FbQTrle1o/lx
MheNSnk81TQoUusWFkv5rdV+5RvGzR/UNElXNsVqZtQmWlVTKE9ZE2VB6x3V
VkKt8JWFx1e1AKNYLo/yKX/1bcFlimvB/qKgkTZi2XtrDRTgjhFRlndDuaXD
yX8QbdkDC0394SWtrDvgCjanBzsjTRH7rW3DwfXU97sMcb3U+Pm0Pp75FIzz
ybMUvKtbgndUZC+qmhJo25eojU03tuktYc2iZipZ9jkdLn7LA0t90PhyC+BH
rGTM8DHL151TjWz3pYj+rJVXDm9+ZO5aO1xip8T6YEHTz/HHbLrUkCImhyT0
Yri9/PNhTpw434tBFvw9NIbop+rpbUFxIlkLql6KvPEcHokGO0mYgez0JDRD
flrYt/T197ezJcOGlv2Ncq9OuBycs5m+msdWH3vCbcv+ckzSSpfVWUG6t7Yt
M7T757FnRWBsnQD7DyEdfVKs8OK5t5q9IMRCZa7GM/AHy4WpdR+2lv7OLsmf
zRTF8FoMWENB22x+tIuDcqeNk8SrBUwerxpc55t7+p2E/iTlirpog9NMX7vz
5oS9VElh2eUX2lmWO0ZfCJh9h6qntU+P3sjVahK2R2SEkUVylyFWCMjlotus
WAx3xvZFpDQQ8l/YrGnxATSHFdZA1hv//6zDD6cNyALirI2+1HfVZPuZeZVg
ltxroC6Rt3CexbrZYWoUpK8NP1NSpMHm6aVZGk2aOjXdxQRHf3emNtzg2zSa
rIuG/U5wLxa2TODgrRN39/PBWIbztuZzLpWext9gWW8LDnYltgs4w3e+8Z7e
gyQgqVFz8EZTZB6kYacrxsoBlFGPmW5PfIASncsCPMqrgqXDkVKHfQV4eNHQ
jwOVIrs3qQgsdzGkiPOs7iXWTF8e65T1pMcBptGlT+FRcFkPi7CPn3oKZGwL
cFcNMD3p7btX4n9Lnu+ancc1rrnhGE46Pd6EB6zeDpUX4r6gBpTHnXIsZC5O
3xt9Cwtv5akCdfZpcDfqeyYctvPIXcIoXWCR1k+aeMTjwtX9uUF/ARZUwfeh
Oc0XlpMbEeJehPavbYUS/giQ46YQkY6NMTpf3MCWqlQ3E9bExJ8fefYDo0HH
G8qHgoVGtgmAzdlvzHyuCD/PKh0lrzEO/7YID0iylaUZrM95FPcU/XuGI+8y
UNbJTyfUwxRx6aBJs0fvyRQWWxllEY50YoDa9e2jEtXXdHeECHbHuEVMJzVT
IoEcR83vH30TiAgXr/sjcRspzwf8csQH/sKZ0QfyJSFgbX8Te3dEevcrsUn5
uDEYMoPUBrYujPmqFswvlRasQ/HsIbZb+gnUgzeNSiwGu+GsrSK4QSqlnyDb
wx7ptapurp82Vn0L0eOUUP37v5CWFwdn3OeABlsxm5DWr8WsMRZsa7xMu3ck
v2fPoy/klp5MPDWOm1X5Pv2Mxmh3dNh+4k29CuxOe/1h+2BVJlfJikzfqPPt
kTpSo2XODTyeQbd/6XfWft2dM+wvow6O82Jl93zRTdb2B+GG6vIDpvFgfXdB
yMqjzJNDUulwTipKH4URwJNyM4PdeQDZTeOU8FHi2qEWfdkpcRR5YAQwdrro
89ClvlWIUXA4+2YDQApGCiUBHcFzoKP/4JDj0zrdCZxm9t45aUQ7Ym5HaMJx
HI+rbMf8y0gMEwaTN/2uRQIr8Qn+CxFO/pf8b5ADqSS4sQKwpzVEG4DJFwPE
8Oys0kFDQ60Iobw3y2QPKx4ihm2+oNvjzlllxqPEnesCWbPl4mWmNYaMgDv2
at5l9dJQ3d9heKBpUKuHy8+7duI5GHHmbRNNKoSdjPQwJ9S4eVj4aIjDP39S
mvoh2Qe0B2aRszcrvQfDfkTrVTKER/17/Hi1UCdYgMs9oESW5rdqrmNfdU9y
84NpLyaRx4e9C7LZB37yCDMpHExSIuG9AB5gp6lrl0M6tAlLQ1sXC7N5qNFF
Gf5dkadm1CpniCGPz+gbHYgRf97zoRi+76U5/dUs9PeihTpDvNqyuIgEmtQl
sFX57PXJ2m+tShxHWg3agMJSPeIp+YQYoqIrwpAKhhc/bGj0UFH/PdchY77x
utsKbzly5C79zq9jTMI4FKbPc50yI+vOrRJX09EoFiHPvv+bq/wWWOcjxa9p
DbGg06rNS2XiMGSL5ppuqr8POC+zyThq1p0Ezz9h/htU/Rufk2djaupjMSTA
ycEUOHKCXxjQAAMRACOa5+DhDnP3SECavtdl6WO5pUDUHoueXsPNPcpkqoKf
TUTOxEOTLAOfXKYcl39LjJ3ZtswcqoUJwd/noJekZNu+q7LVMB3gnLsVOFiQ
vCWHg1LwmAgHpcYQGAiYQneNsxxxi8SbwOC0TYzjR3fNko2XG4v4WwDUzVqz
g5EckaJwoXSXYDM0+SK7FIlMqR2jb2W9ZF3mlZHdERAHUJA4Dnd9++G6jPK6
9tLmzGqD5vtka3PtGP+kr1EiySKgSVY7+/U+ILS3BtJrQA6ErF0zuOW4wLI9
tqOZk/glZsK+o21GG93BsPKAAjHV+jcScjJYSFfOknA4212jEbrvMI8CEkTZ
Xa+0pYXNN4zFZV111UYLff1sp5F7Amrq4nWO1rA9Vsvio5TWo2SSdeCqCYKG
6oyqIF4MFvu6h87QaECbYDHYPphlk7l5KnorJ0AmrX3Ti6gkABrwJMXd8pTe
Ba8Wfh5smCgIapr37jQKnmh3DM5hEtTw7Rq5I0omexi90PbVKGvkNeak7JuY
fGHan0EUI7pbk1UGowzrFR6wcFY+I2lRY0GWDEudBHQ/1cvYuJxW6OCbQCIs
ZZeOCJXj90dTb8NDRORedfka01xXImN2kx/WqGnnO+zLg/JDGCcrd1SPifzh
uIW3JfSJ/OWfwAJlU/D0daHjBWbO9IzpAJIUru9LVgs/bRcFVVY0/jzSL7Jp
PuSU2qhP1O7/yBiVH7yzNta5aLK0yNkN5zlN1IjFb5l5LRfZ8/gV/YzzpVOB
ecf7hb2qyR5DYDFox3Fi1yulySnhoLCNFAFV4y2frYYok4xc3bOCDTVLdmIb
sNxcj3gZlhK6YcVW/L08/InSHGrxpUXbJ5Xd/Z9dVNzX6z0kDTexc8p9q4km
Jf6HU3QOtKP7pRE1KWHFHpiAV7XL0FvppBf6QY7ecm2gaggF6wEsr889LYX7
yAfoOOuRFi15B+uuR6hznEENn2DlRFCHqq1BCU7YOzHPWjJxV4bf2GbDMe6/
54rjXhfJCFW4UncSgP4YGQ86ZoNuqeWms8jJaKD1Q+NZ33iBz8pOeZr8xPNw
gZ201x5Rtp52hs3iB6PirMCVeOvqocq0Gd2V4rzgRAU9/FekAyOMgeIu4jh6
14A6205lJ5b7RkWIjoVFjjUbhorRmbN6wkQt2DYeA2TOAAFfolTd5UP5VylH
YvT6Y33KcTxJJ1/t56vIeOu0wdBlYrT2Y8kDuC3/baF9X2DiSRAnQ8I3hM/c
1z6kxGT1KD51yNN9MLOgg14zgJSXyu3XpyWTwPdC3ldL7hLvPAJnEWXj1Qis
nEbJECA4RLYlQYcmOJsKuTonxlctcUK9FTq1qLVB2m1B1ACllc80t0LZBuCh
7pj0nu2RJ3mkb59FSFxmn6SXCMxm1GjH8d6j8rxNUkpleoAWIwk6+FANaxsu
P005x2OOYfNsLwgWK5YSnv018kb1sAO85v1hk/s+7RkwymU7YSUiE8uFi6Yi
GfWhkYgV7FH4hZVSHJA6VYCUobk54t/u2VhDYSrGJPxNu4hI8RAx2M1Y+Jys
VFzos3XM8Obd0xQXsCnpdi/V4QMk+zAYRUW0SpHLvIF3kZYU4/GZF0wkNa/G
CT58DdcHvsDRF8opLxyR0WkywWFTLAgkc/5gb0UBm2fZC5qBJvXTsGzrRrtQ
n4/xRwfHnhU2ywzKiiQbGFmSJNSb/eiHIy7Gm4M/UrrlcFEO3c5TF3WxkBZl
wOwECTjrEW4VSjBBSagKAj24iby38yFzP13lM6GjD28cVOc3KJPNxbZa+6i2
3F5Xj9Wa9g57kfiIdApVAnZckySQQMixJyy/uV7mwkRt3lNlM92RXWOCz7FD
fCcRfP3ETov0aMKN73TNsxoAuHUEymWrnPKamByIaNIaio/nu7KovHoGzCBg
MqV22ZEjVA0l/ehaxQ7VtZ/BkYLhUTVvXG5sJp32CmgNs9ZFnGtW/hfDRLn9
14/4e5Xc0KUUz8G9kdKZ61AF5N4A7rLX37WYoh8J6E4tMNzc8dgno6fGsKdx
5atIF4i29qL/XByU7KAoIon/GVNWwht2EueRfMfLzqcgKihZasUR2qR0/0Ay
j73bRZme2A2TZrbZfP6xXrejiko7sfSdXPimaFKLNAthBh0q0ANAZJZILGzU
acs87I3HYT2b9tZ0MtpLQE8qn2VD4/BKdIitSheGDsJiJDy8zgoINp9saKGV
tWihkzRIl+uhMyV8hkSNY8XHyYAbRO5wq+VazhccfHHBKXeC9epML+X8qLme
mVVm5wIULlKcIzR9Zdb46y3Hf6dqLq1qeBReRQ7jq3/edPvbGVNl6Q/gFchm
7AD0et0/7/ZvtOwtjn4ESAHywtjyZOAar1SEt0mHk/B16jn2wNH7C7IKDFAC
4RSI8jsnL5Z8gX9PQgA6FMI+MiTQLUp5d/RHluUvI+Bv9btDntqyiG2Nt6Ne
bHbisNQKNndsrNbVNZvdi3g4al0PWrkkHSAL9fEooilw8O208zP36vsvWnEb
xwr+29DW+dqGTYVfvEALNMCPmcGJoRp3/kNj5pnIPJzaZNfuI1gFtN3Bx8l7
MIgSe+Ji8HBlMT3rDdZTAEQC5erEvWtFKumfVls6uZMnVmsE7GaxXU5GK9jr
mOiccneCNXJYdFFlky5+HdhqXujtztGssW+1NQEk8rdRlVaJllOfJ+kIFU87
iQEL2d2YrxSI+DMlWJYNvTI8HNGWXBWbfc5jhjV2nqDCuslkKNv2OHNpHjNj
YBApwqeOLQzwo+52Ihues4Di6w+gBDBneCN+iTTDBkzD9vHnAgQNYhJGtBFs
Px7i2wKVeXeHwiiCQ7MKlJtzEZUkvJruH+61+rgtfBspHP8bYf5bMIArZt0o
G/sb/iTyW2SsixVr9/iLDwP4KZGHcYlzP9lXpBD2u6vu63uBB1fJS786QIce
yjYX6UZoKObBIjFEr95x5Kdeef8oy3IEjXN+RQn5ajNc4QzlNEQwe76+IyTX
qgbmBr+M1LYzs7g3LBKcgYL0rwPg+3nEHUNxJGH2NwS1TfUT3ZEQAVeHlBVn
UNn/fEs0iPv3KuX4RHnRGocV2/sHAAcQVAM+OEWKNHbM3TkPrehF3SoeZGLf
fmW6oDupb8VrzJClYLn5jCX3YTwRyjtrvEFApZKI6hO1+0VObJMBM0XLlwjZ
oP87m2KXMEtRsQQazU9XZ5PTILKtlr/eP6Ri0/sPrSBFuAp2WHmAoTNJkdpe
y9OjS+Bl9EBYSRi0iYCLuYjvuATIKsKt0Rnxe4TejZgaI2l5k3hbG/ksK98L
uTAe9A98p/QOPcRZf/yW8a5f/lBgMnTGu1bnEOLPxJYWI/uLefKbtpWHUW5L
PlSiTXFJ3pELh0/z/+D4e37rSGNkEHwLsdeLdJUpRcpOGYmISPh2tGC2PR+2
LJ7TwbTbTJLKfeyqawj4fyfKzvMukV84U3CHQJoGREB/8U4NTUEUTBgZpkQR
v3dTKlS1owf3xvuVzQ8Wn8QcoX/6Z/0aNxzRpp3vVdJM6wvEIoo5CZhXbyL9
vKW2CJUKYqAUlaeiPOeoQ9NvCamywop8daenzwdUPuA704IliW8clA/NcZKj
F8K1vyndOOWaJbbtJgOyU1GKRhg+gIxH/NIoJxU5GIC+wdQPYDAaDGsl5v7w
Ft2sMhgO4dcP+aypc7eA6lU4zNBKgPLhAUrhDDwuwTxvGC/A9LPUpkYCmuCA
cjkzCR7EYCjTcjCu+XlBr5K4gUwGueG6DuZeLpOZuzi4zygQjbdFWN+UGmxt
kYeazYx+4rxzSWGz85MupmmTtT47r4p0nOPVZPPA9dtTYoGN8hwcXDWCYcKU
wrvPLklgl0OX6EUBR2A+fOKnV8Juqe5Kk9+meUrxYgfT7mOaAjbsTJhWNUZ8
1U0ubEz/pNu4kY6GxDH14Df+ocG9WYlZDbHEUKkQnJVCRtHMU8exbSCtw0Ji
jhtTSLqp2O0Dq4TWfPVjcAJaFO4+CvXjNRkLvRz5R0mcvAoToRr6Y2/qF6c+
JkJ+iAfposYuFiKmsuK2/1eEx/XzF1CY/t97VYooBnxQV9paPsZT3z0ykeCn
tcUs8I1ISirlml2WN/Le9xWGVUWN3TyPYf+ZRWIHtnpGLrMXt5F3X6v1V3/E
PclhW/1nS0GZlxvs6bcfHYC5+kDoEHYruCIOhIVIdDWgDUl3EyhKxqgOJKjh
+BepRdiRgLeDxQ5HOEb6XestUjEwZFuNiK0wxGCfyhXcQhD4cn/KAmb3K3/O
Ld3j7DQdiq7aYN192d940hfrXhyr2CFiRLQTXFkT85NhAauLzS1k2ZJBs8Bg
PId7mTqx95cnWQCV7g4iGhNaiqftaA1hQJOeUlfVAwkiUt9bfScMoyMliT0I
IZBvG41bVgEKebwTEc7Xw7+HkE3vE7ENkusKM23pKcjHW8ADqBceGbUJopVq
lu0Uk3R9YElh1TSdl6gkUvWlOvL0HIAgQXajtCL0vaNonJVxqeIbv/l0//Dn
lJwoSUnGNHePqofHKDj8p5j35gTz8Xhx02fsdFXZRg6q4KC2o11WA9YpBJ7c
51Ib67MHxJaP5Y2oPBEXrzvH5EdHh6IbhiSdY3OOVV1g3TLJeEt6AP2P51sL
5vp7Dt7THtebjSojEtm9q6nm4xfQeooYBfH9g3DJY7jJMhmgWkCX0ngO1nNB
XOvSmrm+E9Ckn/mKqEJZDyKNFLB7Cm9wMwzH09sCAlyPbkU+Zb3RD1FbmrH+
l1476G3cvQ4s0+SYwx3fKhUK79Noe1Z9Cp6dMrp2/KdgMdo0ls0uCT135kXd
d5kiZEj7qEmFev0X8+lGtBwC/IcV6ZF505a1j80mYLjOS1r8bXXmJ17zEe/o
SCfvwu61an+qbz0qmgyQCo7bQXEhleUD6kmLtJLTsZ3Kg1RfzvMWzeXFSfaa
P/ubKWP4yHJwU3zwXOsCU0nSt4s8MJL++jqSUzK+9HbOnhQvl8u3BwQPmaqk
vWcaUezpiimoEmNNJ2HQe8avqAEBu7L8CnxU9S6rxo7FDJL/B2pSjzrIqhVW
wXt3QsnuKfyWX17Kn/8TrDEsf90xdkTMqEG6Guiunn9szJ7dqdUl9tfYcnoU
XdcdXYoVx6lMd7XW/ij3aGYrWscw8Uh1sobhRMzyVB+OU+bfGrMt4fT8miNn
J1NKgOko3hy0iDQBA3KVQKaeUyC8eXFAIItskKtX4dwYyNtY4GP0/DTlKgSp
+qdXxCT6ZF2MMSbJ2GiIUpnHDjOueFZ4t6Hap8VySRNw4ly+i34uXeg2NUa0
MnWo2TF+aXipgdt/tC/H1Fk8s5ToWLRCY93DzGJjYIXY91fbrX9B7zql4qJb
dLZvf4S5NXT1szv5Gg9z/m9quchORb9/uUu5ZvlMBGED3DYI/02lcFmIdF6o
YcHMjHGN0V68WJck+DO2sOUPhzpsIpkLaZ3WvYAd7h874CfrO4Dyn6YJlYo5
RtbyGJTBuGXZ0dzQRwmpTe3Nhj1D7Je8C3MzvrBinNh308rl0xoWyVcjXdMg
Gc36UoPqKDdtX35+M9kor5RLZA4ueDlYtBzqtQ5HeHA5LwMEeCkFV76A5vjQ
vIkclWdOS7kwoOVtCXWosZRlNA/sik0Lld1d3nCg+rL/Vow25tBGwC5Zwfuq
annw+5lu4McfXCBfnDGboT2+XmK+7jv+OSHI1mowxLm606WkEHTQMqyPpQZl
jargWWS5Xqb29dzom5VFRZCYzzSBzW8Q5U1zwNEOsMycvlLjhTf/iRcktdnL
HeiiZLwjAvLumqhuQrhk5yopvC4KnFujyn90oGHr7+sijQUqlqAoFS4PMOTu
N0jTNMmaf/7dvNMORGfXAXKrbbjdryntGu39X8Djx5XZEc2GBW0sA/Ndi9R6
x9K+CvbpAMEG8QWWDV8rFemLZ8I8/Jodjpu8WpyIp9UwyvUo0if72S4xYg1n
Fd3/y+I2wOoO9V8czo80b2RljUS7GhBHqCkm8mSyZYJaoLyhWWyrxlEWpnRE
G+j7p1zC5cpcJBhCSPL3lXBNkUhdBPn4YA9O4u7eHKEoVDhJiyx8E3w8d7gw
nbm1zxry+0hxwj2aVylck9rVBYz/AwHVzaBiNKi2H2eUODxgxGwt9BEkVcT8
9ohUQoZiXbF5GAk8kuzfFQMCT1a4S5CCgiEVZCKBCu7BKddb+ZDbAScJTikq
wefL4GXuPjlVY+/ZGWCaaCXiWhAKy9sq0/vDjSK21pkVguy36AaQGlNVLenI
m/bKeVZG6DzzT4Gl0PlnCLapHuM4ov9wo1wYDUw6gbgRSGmhq6NFd216R3ud
B7DJH4/h2MD/hJ3tvRxluht953ak5wvDZ/MaXHXMhdWFzsNOT5yo0sP6hIGC
3LL1W8g9uveMOdCL+RT7XA2zQGPvegE/VFJzjxU436VnjaqhhTAsxbSyT21h
UH1j7Glj+SV7G59CTND4gp3Z5DaHDGyq0exvNatH9SXSAcYpOTHESWiQnN7Y
CpCQaa+TUK0/t+TGoaB2Pk6WzrKWSRfq3lwCESxWwc72AXihuyNe+PAk0R/j
Wy+AorE32Jn/VBkxMU2axniXZOFHoT78j7LSjjGFNfz0mYPr2o693iYPTvxr
7zV4sl/PEtIGaOJ6OEr7qYrNWujUqe/g9t69fCsS0oOAFUIdpEcgUpZBubpR
VuUttmN3d60bU+7o3iCXeRVyFtYjkV7QoVIlKeI+nFEp5iH86/OyHc5qxwsi
Ea7PbB9aK8n+e55aGbio9tR4sJvLzlWPPxd7Yjs6acwY/HWbvFnQ24RpMC5D
Cee577JaWz1Ors5Y9nbxeJBjU22GEh3fpDMRYVxuWx+7ki3NG4CPLrGbvQrs
ZZ4Zgu6/q2zs0xntf6YBLU2zsnYZkQnelrmsKRCyO/lGa+8a5lqPNSDyQK0X
nC54lQwlLCCyaYqk4HxVyrHwbO/4HBH1LLQj9AcKNkJ+CxsACx+2HW2d4Rm0
D0EKM/KzbzQAMNz6e2Vnnh0e85fWdyobgXE1rWZcguimtjFYeb0lQbtSZCfm
5D/9l0jqLPr5HMdiqDCD4tr0l0tlwbnKRi5PKMqrCQzEQmVlMpodwZu9pmVi
OL9B29lRclIA7rvURmjmCfPk+GzMQd71jxIcnEor5t03Nimfmz0hiS12zLrL
3WISEAKpqsBjKLFP2tbAneXJWGIc98UpouOYs8O6o1ZPc8iuiG/AsdvxnauO
o2Y7SXj0icCNKmJuX9kK6rBPrSjy7u96OzOiAUMPD5RAZuLs9VZZdIgaXkQM
m0NWpfmIfsnCC+4KcQ3u8JzxcOcJAYl6V6fOGpBzZAbA/iRVrtKkvYKSxcPH
Xg11gdH60KKAmLiAV6kxS2Vb+a0twtqCl+Y4uqKsG70sMRBQ/EZivWSb4myZ
r+tUs4fixMRWq/yk4yPkF3j+KEkPCe9zyhjtGLoLDQkzu9Si8VUU7MeonIFr
DUJGypaUz7LcqtBNjVzoLYEqHJFAgKjEvrGOhrJhiwYiEH1Vs8LX3LuyoAqq
crg4/moclRsZAgvdZJQxiyFMinn80BAeRU8xXh6sSbBFm7p2tRyVOJA8D1RJ
NKmLGtPlQIzVc0oKDLvKi/YyWYiDpzV2ETodNpheWPsjY/mfKQmU2MarFhQd
cnibX1Vqlm+RnHXWNbIXyZqMrV6DKsGeo5xdYh5I4tfgaoYLu7QFhe0Cq9xh
72BJrPaGOzbwfaBtcLN48Hu1w3rKcvD1b8VP6RV265Vo2K+xPufxBmw8F+ny
Tx3FNskDLMf/V6ZgM9XnSWgatFvuA8LNl6mud/N7QMLx89FphYl/PPPoVKnw
roA/Ib8YhGcmoHfT5RJ3E1wf9IQiuOIdHM5vv3YXET/fF615U+xgueWtKW2U
/AcaFdz0VPSo5s9t+wB4+qtrkmhnAa3O8NoMfQ/QWUiQk7e3W0kf77rFX20c
iWe2R1/PE3zHi0UAq+hCZNZWZkan/qFeCeHzNHWozu1h9/w3UdUELC7lAK3i
SGQT01+ER0KmB1jJRSO5ZAyrRQnHy82SH5q1jXHERlWCJ//PW3Y1CxpudR1u
fLSN9QuGrJ/STVDw8KLq2PY8LXnmvU0oC3gQBTb2VHt/t21XaG0NTi196hcA
Ogx88IVmhpurfh9jVUIBzIQ6//tFcEMEgVsiwubLEKjK61/vdSpRUzhq/7V1
e7o+zn5L47CFMtNacVVZFpk/s/AURSP/9ojeqzXjSmoKL7sL1IUpSW45JPL/
9yXrsftpUJD+39csZ8TPhrPVLOC9JGys/6idESlw6loxNwNmuQZds8Z8o2/1
KdPWbmdj5YfSJPeOTpFSoTbkZqHQmgkLUQU+YDbMKCMqsjFjZXzhBt68HqTB
ACPba+VNK2UR9pYBTV7OKoOh9VLVVbQu421KsslctBnzs2COhvlLbBpaBHpn
e6xkW499VMBfdvs/qUJoRfQgyoRVbXgpBuXLIUgPxaV5OwEDZv4piH0iEjnN
PAU4uVxrsOnwaZX+9YDImO0WjWzqIOjH0kZ3WTR0wh8m4s7JHaRRnBWMMTK3
p8/CBlbV3u2yXyd+kn02qB2hSjdUMfB94CDmJofjBbJmcU7EPLlS20sIu6tK
dFuadfBTdyauu4zDZWFfolV/4DKcmfF2Tyn32zR4QVwmjAB+Qaey6bHoGi4W
Ge5ltQtqrXmZiJ5uKgGOSqxXFkb6CheKC3ybEsOgrHRJYgRZ3LIVLwQWoNKh
HJfmH7gLVMnchxFODEpQrL4A8ApV+fYatwzcILBCikbHTKTClY3CRQjlbsU0
cD7OushXD+HtNsozOE+OpQ3lyZu+e9ycQJ8SGxNDQdpT23jHTL5c7+y1cXjU
sN3D0bGYFYTIWQK1gt851rAH73o185DzLHt67EoIQ/IQIQBFf9oBdm1OQvYT
a5Em4UXuH8vrIs3PwnpEWN/7H1TRdNpo4Hr7b4GGVzrpch+xaQrcjVrqieDZ
n7XbWr2Sk8Spaq2yUrZKhMu75GcDPJFJttvOF7gKMms1P+LWfovx06TotfFq
NjMPlTofYCd+J1RYTeX6KvxMEWe7lAVrbsAigz6yjSJCsc2au0lNMuPqvbm5
It3STEC8yqdke9D1dqJvUIuH3Qc3CRVv3lf9fhrouNOXwDg0VqisSydJb1EG
s3pRCWvRUvIlBm4tHF2j5yzSqrWtrheBV4I1hdyGejAVx/aIYIhO7jycth01
9FLwbtWiscsiOPi2qQE8ml1gjeQT0EFbQWGWlJfhrBpl8JH3bgX+VKKa7U+Q
eLfCy/29OPovNOBWzEwBq6f6kt0XyOFaAN1RdRN/1ClmNY5pCMXKloq1HJiA
2800/SxkgL0ShHUFhq+YPWEl7OpQP9v6PYy4YOD1/ci4fQbshkhInRntCiYl
5DmTvBWkEeIJcxVqPqFUEnAI4A6c0DhNLfpO/x6wqn0B2zddOTeQd3Yo+Y42
9sMhTgythCq5b7uAXU0beQcAs8UqcITxjaOIZAvQ7wGv33lkcxOQUNge4Toa
Z2I+lNgeL6FZI35XCXu3DbW1B9QwtU/se0djvrDL/+9OKlQMq78dY4fS0uR9
Cs1Xp3ANbHGfp4CrgRn4srQ+FGvosbn/huoUFEazUkL7d5saBBA/r9ynWDqn
dErTYUXNrlAFlnIVDDpzb1x8GRrJtszF1i0DYzuYDf6wsdsy5mHYogP2HoUN
Y4vK2nU5e8zRjbJPnw7/tnA7uEzUpXOWJ6QwFYocqRAcqG/uBd+sbs0TygqN
84CysdvyTtwsYkc9r3D0qoaDj9yQQwzLLK06/IDd8OXTJ57XkJNpcDBBorzE
rWi2XB4u+ibBnDoZu2cRWHhBGmouJnPEUm/ntpWYKvrtMz1NQ0V29zvBK5mr
ngoczydgKd9oUkqFXjNJAClBAiO70KIUIK+CENf7aM+iEAB4lfVNlbs5TODj
ttlONdX66/W8OIvrFxdSEJ0XV7rWRYC2snVO3dQuepymRHx/FZ4tR+EIrMRA
7mouGIGxBBp3sgT6rBb8IabObx4AhQUwSBhTO+qwfSgw7mYLOsKllggzCQ8S
nQXCWcugJJIirNO6+csT4C0ptS0u2Vu29oIqMf4TjU70DrSjlV3+hHYSho3C
YkwztJktgn0266T8DYMXyDQfFdK+uUdnUFx7+wWnrSudS+gYt1kzG5jEFyUL
7js9Log8tG+H6dmrWXF0vKYlmbwf3UFCP7SPR1PyTNp9ds7rge2/MSnEmxkn
REWXJ7IGIwbJumVu2dhrOTwGJwX6KoV0A83IMqHY6NjGPPz6D+vOXDI0wy0+
tfk/nIOc415DxmsPez/4fYrNkQICkV6cgj0BOnXuS9Lew55gE6iyKAE2oAni
KE7HQZPGaAZNXwgcW8DqXcU4ryzJ2QPZautthS0uv7muT9QEdsFtT0+ZBFvq
lhU+qXVbmT5bHTxQTQj21D8LBh/NLXiF5FCwhWrtUgtPFbeeAfaipgehP3pc
fws3lfW9mhfo9FxtTK312oVqOR8NakvN9WOK6Q1WNNGxVXvgfFS3uoQdxm4j
3L5VkI6oHuQk09TgYMVn3u/isAQAMYzU66pVYkTlbeWwBVdlkLynRE8DePwq
7jGm9H+XyDVPi+oCGrx1nm+Z4en/YPenDb0Qk8b/+iMI0BTU3gUejuAK8l6c
bcCDAyOiUl0e/8Xlme1E19I27yCW/dfIQe81x5LeA/kUMqIGn0LTsZ6msuj9
KKHVcuBc5uU5B7UGaskQjoNdQg0DigF1rsfRNsO1ZSjUBHzwk7xgxEQgIYOR
nHHQfw8wrZ8opCZqHR3JBFSqr2cRMaMFhborJIcYo/XGEpbvDR1sX54Puuc1
VMUQoHAt4hhur/ii2UdM3XIpchdOma3Bry5Fn2V60J/HeVV7Rg8+l1LQZlWb
RyCHSHn2GOadvkQyeDm5do/YHQmks3KAJUsBPlOzV9L59xiBDPqev1AiEvMg
4VSqPF91czDIUrFewKPmcyWHJlbEz6YR7NyXHAEnfJQvRSD85KBlpi+ds6Lx
41LkOOUrET85EVo/KmXWXVTJyHdAqozHvdp+JM6OGr45m/wWvmQWG23f7s0r
CDGhkJeXk2qI6JpHQg3EXwMNzSGyybraO9sQFOX11K4tDOAWjR9wjyk7aEho
q9Wx/tCFmu3Dp/TSRRh9Xh3XUw1MfvE6LBrYAkm/ATmTlM7QWmAeXKP3uA39
wfMEd8h1m9mLPGXtMU27U+VxUCZaoFk4h5PEYLigYZEEk32goLeiPGuE5zXb
7Ua6LGLBP6i/6PCQmo/VhjbOnxO9H5s/YvJNJL2Bu2bLravD9V4Yrscp0RaN
irvqQelb6VxdJ7jefQnqOyUNGzeXC8qpAD8AwIq4Opxp9T6hRs8Pn/dj+7cb
9bZnF2/Ux3o5zMC5rzkhVtkD3q7Bc1LOzGrw/5PE/0dX52gswBktkHfiWjEB
yKWyy1QJ0O7qJa/GJ3IKTecDb3CwabKFxeyg/2dKveAUM/r0yjeRBJ3x0Uty
x9wJgLQ6Fsh30xWNUCLKs9p9CZOUWwwoP3REHVZGdxHO21dAJ24kJ/P7F6RH
u5JVeB/Pjm9V0ArmYzcbc4e6yvnFXarjwx5H74Q0YBYmGCsiBKFxej/mvEQz
T4G4mI4TnfMkPKBC/gE16Kn3kUxt8sJKXIKe+OdeGngaFIXZfnegf4ptEa/h
nkSPiqASY5pcnfBIpzoSk+1u1mjwrKNDyHyXQ0s1q8Zlibszzyipt69NA4Dy
XyYK/McQLqtntjnyP6A7iJaX1H1Y4GYJJLojM9RzX4Re8TKe4ILRkYHzdHrX
9XCt/3ZZhJc0JM4Q5n7s+6W3UNebSsazelLJ9VptrQm7qF1G/YXWgA3WIkkU
sqwfTvRqM9OpgmRNFKTg0TP3yo1oiItt1kmcIg5rPiN1LfgQQsfxqZVuYtbG
TbEiuha12C+1/nDLKSM+zmLNI0YGVp9ZnUVv787nAu1R91aV6ibfP5LB08h4
EfQ8+Xsubu0/S6VJu7umXf9K2V9hgHPg8PAa/YkxYkeUJF/mFgXtEDM43fSB
1hcuywU2lpKFZ4NyMXUuC2H0B5Jx6A8dN5Q61qghzPKUZoX8xiti2tvTey+s
LV0vDbziGWNSoBVoJgK1GyvWQPeiWlsaNyJZmcvjR+ZdrJ85ZEKQBVgyszii
RPhn1eFotJki/1qugJVKUMGRN3BRuh/SYoPa46iirt7m2FTiQFbZdl95cgH/
3tCW1NvGiwd5IRE/60ePK5wTk596JH1x4Aw9DAU4+DOm3CLQbAx+YinKFE0+
pREfQq9Tv7ObJjlFJHi+z82LDyL7ExsbWT1XmH+wl+o7K0kKRpPsqU+qVjkj
8gQ5pWWmF9jgsV4vUdSsem65+xW8vhXdJxr3dEvgbz5AaUVmvtQRhub/EYLg
IheZvI3FBdWVKzYtK8qvXfWdVXg66kkZ3gq+c8gEhaqKIz9p8WkEQAN1ipo9
HU2+bfYsaVElkP5Z6WW9SJuv2zPJFZjsDkQIz+YRGPBq/vIf2QAEP3OKGT/T
vog9/u/mT5qJLN+aL5joDLThhpnC5C8s65ha8Pv6W9CXCJVqASfCaWhLQyKr
K33qrpNboDSWRUgogwRcRO8FD6aq2TZN/3BJiywE/gCGFD9aTj27mXGM5vgd
Q3YmZLB04yoD9ZgKLmXuT7TcaU34ZmIWsEgdiywcnUqjZFAH7VCime4LFpgx
EIg4K3kITIkK5Vr51yanEujE9b2TxXZgH+pMIYpHWtGCc/N+p6EzIFPzv4Av
8GubFcXTdZjeH8xa0F31fY1egBHN1ax1Vw+fl9wNmSEVzoVehiuaQ5aFTy97
w2GDxiMYqB5nPhBuBc57kWADiJEaI7zRQlOI2unxocY82oSs3IwIvojkdijD
Pg6hmv4XWVxLuK3Yht95KTEkz71ybEtge5uRKpw+LhH0cFXiStAzaCfepzmr
wEfYEYL4VmM9h1xXPlZ21V/lnIzlKiLGVDJVQDSZ7rtZnRc3gOYCjzhWq+p7
h6bLaLHixbMPrE3PcyC+IJ6tfOSwD4SRleAiqf+xO1dtsM8DxVohifyYIJOm
MwkP+jUV7NRGOg38aYb649dD+vGPMnfzaphcog4f3GWEhkJF0XxRMPV/HE2x
Y6THuKwazLelDPxe1QU2VaMx4dZCIBY4BqMl6etOjRiS+DGBCXdt0/+DeNo3
3PPM3h7PPiD34lsWkNIZrvQU0hjxtzlwCy/6r+9xYcgwWF1KU18Ppz8Tp0/R
CM1Byf8NX5TuE80pQKdtCdeuIXCG354qnTQAZrjRVBGzlEO4W0NmuJWRf95t
w1z4yFZfOx7S7AWFCcQOqLqc51bwrU5B36cit4Pu0YFnX8+PTPOe7wIfoynF
nryMKIjFMrS47yDHeIDv8k0SwzUkIlLxVulESTgz0VUx4sJEzwtJMuhaNhM1
PWVpE1t0PVTeDSLo408YhGicAAVpqfMX1y0onEcTuOcc0fJ8ou196WLYyPmR
v3izviABYZsGD4dXwvqjTjZ6uTEuxiR22OWXDg02c/SzmoNF3DSk4nmYQsm3
dvAYqZkNl2nOp+h4Qn5Yh0Chi/0eE0cK4KbbmD6x3qr2W09ky3OFqDrJM9Uq
pBlSpC42OWSj1L0/fh0GXrl//d/lTsApgTO0K/Tmkucf0fF+tRzJdDgUqMFC
oMFzTPWhmX83AiBAp5Mh++eFVL9+7MoP444W9XksS99cGhoDtLCxWWusBF/D
gohe5oBdxBW6oPSiVJdpqc6e265IZ+TXLPAzj8pYfN9fkPSoHUNg7XyMfa4b
G+xgw+p6eU+v0KS9nTwIdRVMx/6rBgQ11a3e6kDcI0dBheM6hB11EyHxxd0N
byQULVBZcj6UrhrdWMX73HJXsN/SxcJ9WxOV4/coQqJN4Uu7viuL4nPcvGyM
oVqKauM4jcmDuPzO5Hq5XPr8X2xYKxQBuuafm1c0Nq3BPUrDeQtrNbDyGyqu
2krpZ1C5l2ghChGX/mWDHINDgyw42jbSbwphY3q70A2v/Osai5ZbxIs+ATz8
Kv63K2ojx5Uaenq0wD2iUWYxriu3edo6GWANja/H9Q7k96TjsnDTwQeWncNT
AxHZMHnJvd74ApYpgIhYGIw8cVkhLLtWiHiFiwMbzfx3BXdrhb9UWv/yj9lg
S4SKOCBKRpdGfDtj2kAQXPOLln8rpdRzNgPQ2UztiEARK7LSKhKLdB7PhTy/
u5m5gQuYi21hoFh9BJ4GtpYJbu5mtg3dA8Ln0CYvrL5wSZUh7XMTJveqnaM9
GlKGLFxB83awNth5isMOpsVZMNdMntBBaZvybDp2iOgqn+GZUg51/xYUcZ62
obsXkwy7fCKvgNSPWtUL0kv245MmcXKbTrOemh1VDEy54f6yVReatbuDxcQv
zKAN4dP2YTk6Uekq2ZtpEiOdYR9S8/ARVz0WAcJqr70I1bQM2ABizhYvKNcA
5qN3k1NL+VwqTjb3C/itNWHyEVN4/uBwKSgbXNna54wYLYVWFCqGtU8Bju+q
afieE5e8O5G1+Pp1WYojvK2Z8vFEtjZi3dpo4QCLP/iOz32aJz7jrtlNxv99
u57wxwx2BHGCoAcsNzyC7aw1etNHauKjsdqSHtwWSLcWVkS91plQy81GbOGh
4t1r/X9cbwgHRN8Viu6KO+Gi/w+9t1o//IqqXvN6jRC3hkeHhrWiKlyqzDSV
MQsIYsgklFXWAskal87OmJQfOHD7Vzw4wg1OTtMJ/k1ATzAQoteawaeKOSMK
aFtRkKAUv1tS7WXDGe1SnaC7EO2fWT1I+OZXYkbp4f9Cef9SJVeK2e8kUhsd
c9xYMt3d8tsXWNIjTbOG810wxzAO7vDqp1mEehQnlF/hxixeKWMJLFv2Viq2
uz0QKpzsGpcXEw1Z34SChjn/ma7Ep1JdKzdM2caERUxV3+odlxTkFerjZlzn
nRxHg19mduLPsS3AfvXCmsGS+YL9VCmmC21ywKXFLFfP+4ja3poFLFOM4SU3
SzDxlfqn3XzKnOI9D0SfJloHGjAZyGNEYbTxP9V2l1LOeT2YkUWc5InFhfH9
SCGTLEC1yLhw3bfJLLkRGg9pYqUHqba32BfT2p99XkcILooQovhTRqCQm5kc
eNszhNAU4I8x6WPvAYhU0ThvG15x1jD/zw5ifmX0ofDxjL1tA+XQeRgDEfaR
aGYa2KBPpSFxyDrD+xJaC58GuNsVniiWWVKJX6S32/H5AQZkkx/orxfqMeKV
VMEgCkXSpVkUm8g0BU+cBHADnYAHwXNb8BUDKwC12doBD66A1JyD3M9evjjG
Dfg9CfhE21ecIWhOaJuZ+XUGHWM/kJxzJmaOw+3UsO1sioW/zBPslCS5YJOA
NafwEK9NCfb7At7EI9/uWGrZvr+rPi+0REfs9BLWEAjQ7zYWcux0erD/UR8g
txyNsWVohwQntPseUWKTiwVyTApAHEe1SF60QzXxYmgGmGnb6lULEdrSemLz
WSKTLuMzkeZpsHzTz9GGOofe/4w6pETjzcGL+DlEUowEbWx9TT9x6DhOOe5C
QryoAEqdoRLblSSJ2nd9meE1O9KFt9rO8slZI2exwvfz345OrZi7Xok8r1cS
gxF1wZqZJm0zPpo3hkKTkvK/mkWY2XjLwOCgdv9M6xY8Y7KU/WhDT2d0cUq9
a6xl4Ie4XxvbGkxkhXXm2vucfMPVX1qTF4UQLzhqxelS/4J4USlCYNWdvnas
layJEJVJvzg/+lXD+JGwxS8nMksmTcYyzQKMCCZ+8gwyYZMfKSNiiPcY55gc
JfnnCKcS7ne2Ux/dLKUnIC7lRkRI6CdhAYm6b8eSbfR25p3KGHwE2fKnOCso
qHPtnlOy9K9h/VnmRKn6ldcUdvLXBLeS4rBypevCnWV+A8j7P0l1AzDWqTyT
MeqDd70CFQ/JJkGkEHX84o3ihAe7KEVS5XaHx8w5PVUSTSeLQfia0oWSZt9n
/YWqJA5TMGTN0OUPOeFkBp6Ss3zGdZm2+4vwTG7a5Ste1NULJVh3Y2O84kBr
trGs+CFbPgOB5+lyufTTxuLi8Hj4WIyDfIWRrwf9Zbr4A96FqFngDrLJDqfM
0Vy9Om4ZqOx4A68JqGIHdwF862Ead4wIqwIJyNqqxohpM1Tb2nL/YjY7WPq0
AAddKV24z9KR1gqPEoQSw63SPyTMkpJci3GRw1oGZPfbC8LjQXob+1I5bh6j
whsExWtVRGdRKKqlCgzaHkkVjtVpy6LcgN16q1XGC2S49Ib2tZMgUVmeCN9L
XLFsfmGYG+1JW6A98vefhCa2GTUBR76YSQiT7Qll0cp5zpZ0qDnr6zL2OX+5
ehhikSbIu8Wv8CP6cBoY740n+P7wNh5Isf2LDvcxHEzSzKm6e7mui1/OUrLQ
rvjn8aGkD9M2HG/061S2p4WZszDv8Xk396l8xIetJg6MqSKKKzS4Qw4omD4x
DCgn5iOiIHGypfUC+xmsQkFAvdcZEMF/iny0unIonQpVzC+SXesjhtbQ2vuI
oSYT9y14ulIvPGUmHq6NG2MgDITetrcr4WmXSqfguuRRGHa6wCZu8m6+Np+k
vboS0MEuzcgjc8rSvQNgGfdMjYb/Ee8KEMRQl/gu1dKPr1F7bMOXPR0YIec1
JSjO84IHclsYndIfEq01n2dN5Nb7dB9hjW9VDayFxL0kqmQGiNhbQ1Cjt5Y6
mna1/orpcR8n9cmvt3Co9Z8R9rR1TM2Sdvq8CvSQLl38ygOIEJWTJRRF7z22
nNxWxoWEStmsUg9OQ53L9qMT9nr9gJrIhNhceZb1JkEdL6UdgNhOQ0w0Qxbb
06+/5/khT4IjYZhO1lQICIxXqR9MtIHaE1s1Aqxm3OO7QzjvV8HItvYyzgM9
KlCliwosRjHCRDcr1yhUMW2DlfRDekk5XErGv1tfA6PEzl1wne6ZHMKj375Y
BRkZFXFzD7MBrfT3xuk6fVo4nbs9e/u+KIJIlFc28Z6BueYrmMY9DkHJtAue
OVyLorgKEL4b3F2ZJVH8Jisxezvmonzo+U+a+2odYdnc3WSmTfhDCu78w/RU
kq00vE2J013+SOEJPCxiO2R0CiyezP67JqCdO/++ey9a7sfPLvZLUegp0x3R
/oBEKbo3GbvunkPGQB229HvHD0vuFmdsk/JH0AyuNXz8BWYz4ukHilx4tsVt
ZVYX5qWLK1roRmQH/nxx5uhim9opI1SUZ7n9HT4uD1RSog3i6blF6UlRsuUg
FrasURJuaNlg8zjq6Wt0/FkpbEofSEiaMB/UfEl3ZQCJ+PXzt0Z1kKN9kxk9
ffrssWaSyzU3cWNsmL/qkLB9EY/RIXod7/3qHLEjQA+I2xllhUcfGXP3UiCZ
cS5tnAPKQg7iYL/r1FoZpI0jP03ebD2BqsqZ2c/rq+6pxzH2VX+YT5JJWu1k
xfA84qu2d7QEq3OgD0TJvwqNUsTQAyufQPEsBu1vOJ0FLQB1L/JC2MRrdqAz
HMjRTFtnGJpRGJb4VS1ETsXE8+n9faJQ+n3tyADbaJHqqz6WyuSLbI534yXF
vktmT7iVzLjh+SplC4TD6wawlM0y18xQ94ZzTqDlkGp/v/AgnIlggs/ak+eQ
1iWZixDnDqgfdLlvaH2fk9GlK3g6PJ7UMJtNPqoKwyqkCpBRl0/6KipNQ6rZ
gNzhVxCrBCurxcrR9tRSsDSlqomUL7kLBPgJ94GtdxYR798FsL6kN2vHXq+B
yEhMxggvAoQujdCZZO5feZyDtinTSzAyUkTBK8W2rSqHRLWM3C2HtKX/XbwP
Y+FeyMw/n3uNbBgcPrpYBoecf3Uk/bIDN5VTQdrdR/LMn6Mg3YWUrJOzsKOq
K9lI7yXc+2KkuTdvi/8cENVVcwwyjiz8MMVT0sfZF++deRJoayprGDguYTh2
CAc6aOvkpliSIMbCFdKN69dg9qd7ztTCZUZLJ8o4fm9YtzqD0TqeyUqP3lES
O0q/46ay6K+QT4uDVbwb576hBzhdmfX4VP8rlBmHPFkjxiQVL9WzMgvUMLgF
ZJJFSqBFuZ5mM6H5PlqCwnzPIP9wC+pfsU7cu9mg/jiKMjcur4dY+M7NhmJm
Gp6BqR/kzgfoJNU//U+dY7EpWl/A88L077faipkWXKbpuIY6qcKOuI2cRN40
Xu0ySvb+rJ4NljuTxuw99OwaZWuVNRtnTLZKTcxtZp8zfjrYvzWoGsJJSt4o
0AiJ6+3PETW1WyU+iIxYKaD56DaRNS73Rqa+vOZWGFxxiW0xQxjy7cNR/zrB
pjXLZtSz2UJ12iBAO76yMqjTzoy24C1pvOUhjalzGNe3WqprP29galWNUHix
eW1oWx8fkoAxwgRH/gOxqmOdKczgZyLze85aakHGmt+z+L9+Q2iBKWNNnWOu
DNBvnOOiB1Msxe/zfIs/1zN0a8NziSZEA+9z8dQyJOaJSvNkBxWroIAuWGbm
itmHLsL+FBlHg5OUpukhpGT1VjOOaB0i/mF5xXJfZiQxKL7TXL6hvmPHq+in
45ZVuhkRZRdauAFT4GNFa7AbeuoFORc5ECP5J4UKIujC2SDZvoSHvt06RFwL
IJDR9Dcc6LeXoY6x1UEwMP90SNlXwNEh0xeA7wWZnDdncjrqoAH07xZWFDnc
HomnFRT8M+qndAopXaT3MCGZvS+T3l1/0vsoAShnDiUvU9MbjYIKk/z5hBPT
E3W+r+i1uX2ciU82b9gYNRIsCqhDCJqO6IxfTjPdFrMDffJjsWCgaMnRWAfp
YH/AbDcAR1umE/DNvjMH2z+nLivnCOVvFs/FSfrisQHjVEMtTFsq4q4UnXOe
sZ0TvdiKLuezxj+gx673mVvf2U1mYXd5QbiUXUG/wjoRZNbgMDR+LQbtn4e+
NixkyNAd6y3trAqlyCkdSkHyvZ4xo7e8iVl1f5fOuKT0XVmN8csbeMXTbccd
/9OEdwKQlngvZmY59iUJ3kRK9+5W9/oFfjZmVloFo0hQjC9PNqnMuSUsaO0F
Hoqok2abvGL0nbpJTNM1cGIctMiWAWL0gnqoxPi19c+Pn5JvszklkKWxzcTB
qjUHmYjiIpts3J3XLqmIWeMOTzMQ6YxSnbiA2WyrlkKI/N61a38BrHNr4bAI
fqWlawiqur5Hz5pn7Gg9mtKaEQFGgKZ+oH0aABNmGh7w8wX8Hg+dt7bEvm4S
uoPQKwlcRbUuqZW0dRL0w+gOYS9hwqKxTJk6cvkWgp2vr2aUFRwk2icdUd4x
fLigCuN/Wuy3UbDTV2I6g68vTeqop8x+7PKex0nudnbtbZIfjKCdlGHF+owG
39jO8RvftSc0cjyil9jbUqVxgGBV0wECXHf28mPMA7xyZfBNtxZFnxjPy7+8
4e8G8liDNiyptEjCybpNfa9fTZ3FgeavcP3o9kGorRnY3qjcD/UXqPG//wiV
YvrgmpXfoDteAuAfgGkHYnNhIW1UQ+Aeto6hyS0B2omsk7xrhWuDKOt7wLui
84UAEje8I5m+ErLiw60zqiVzfqlcAJwcqD8oBYC4gcRCKqO8rtvzm6Q0idgK
DGvjMstMkL5g8NAcS5mZn8NSDskOKS6mo1IU9bvs6G9ojffZGsZjzQxN55dE
GOgg6rFzUIyzmuT7XGJbV623KIF42sZ08B53Uyo4B+e1cqQtUUmOoujcr+s2
ex0vcFHDMJR+ptZ2K+WvGzMUMh7KZMtsswb9YY0R3a4tFwDqV5ylkNvi4qy5
XSEI+4hC6Madutx7jnyjOyN3d8WtEy0HYdnNKUY+3uYfurF+YqCq4fZT7wte
nxRPh7/QSdMinXJKMPN5LGVvFbGouC7X4JrBQbSdF7low8Koz9LOtLUJYSIk
/RCpbE9nla2v+PorBEEZHzUKVFkQOEmXz92w/qt1d2tmQubbQ8xNcQSyjJAF
1DwA+u/YvGfeq+Wti+X5845Ba6LBzET+V6+UJqSm91mCVc6+0TJjReAHpih1
dbcP1ZGDHKxu9crtR6mZ8qsVs256FfVQVW7E9GuAH4CIUoqEaGr0odZ4WtIG
POLVF0gU0yi3Gz962bKRSIAGf5OEP5aq/4iHNuYC/f0HlC/gWm6juLkTLyuB
tjGevc8M3Z8hlO35WDhjbKcWphzAnni+eO31PJh5wWVZeseNhvN34ZL6vsv4
l0gtTKM9EAVJphHfpIpfOEqxjFsDVd1tauri7eTeqhRUu7Vd1wHVqZ7FTFun
W7bBaKdIZGlsAXiulP5csZR5jrje/Wm+xoTcvBmu+70mvMTbZyGg3mJkHf1S
2/UO87DkE2bXQjDSQrVjb/u1wmh4Vw5EjHW59Q3/V9CNzrz0Wy5cCICiYhTB
mJ0At56UtQCEPX7jCHF8JHuN9fTkTTVcHnPEQeSxCcdZ50TPN8jmMgVLlTBS
6atYpKxRPZ2Ob9l8sSmXGPG0HsZPYFTwLRuS/ZCH9yKmSWpomWMj9HMAdray
YVa0fN03SASBVnIXYJB5/0FWwvtKLWWpJv/xFvXcL28kgw5D6dWnanmmfbsW
ytYLTb/9Gia42CGS/Th4M1gxnHowjKugYtqfRQYgV0HniiUJ8l/A5GBFPl5U
9ScBEQA06thv/45hA4AO2YBtbpy9js5jiKa8nwPv+4eU1Gzc2GuSgBky0RdW
QfjV3x6WqBBnzU3km4ZYst2D8DU9lqrSoonG5jog2X1cTBZEKk/KucoApjkY
AEuqqZDRRLU2sezkTEK7SrnnCPYmYJVZBnSFFpQQU4QorXsmdL66IbIXoUCt
boE7YLAXMN+QmRNcNyp/ack1QrwneA6H5Zkq757o1r1gv1wmsi3vosnbxzzu
Tf4XDHMmWcGuJgsS6cgiVpCKEM32lWiJaTuIDe0OHQ2aGT7KWuXRwu3VC+SM
9PsoJMVtThjUmNDRNKcPcf7GNx/N3IHyn8Nd2Vqrhb3z72jSL1VIYYldzH5e
qt5n6fLXcfY6Rc3xDhNQQOyBGZC94v6uUnQdHNPSz6+jRtrKFkfzqpsT2htm
8VlfHbzEn63+BVtiWaOQHOubSn0AMwQqq5F/bPnPTc8PznhjRAQ6t32Z5TAI
eRE9nDbwyZj0M+tKjuYw1lGyaDMoyYsowokR6f7gGx8ljA/3k2xf+GHWYWYh
kvvm5VEIkqzoTMc/zqIdQcEbMrQSyoxm+zCC4j5ByTTU3titqYngscRVzwvL
cuQ0kPcI566t3E1kC6t/EWWOyVMDbFFcBSteT3SM5WOoVuJ0MVf3PdjV2uJB
WaqKBcvZG3sjrcJCIxQltBmgzfEPnYIcFS7L+9AKYrmu49zSR/Z4eHWTpJlJ
KLSyt1bPntmHQUtN33gQuyVS6hLiXr310fYnpAW9NpcdSrtnU/89ZpocM6lp
vZ4esddyv+j2SS3Lq1tD0MopoSYTJBZcdqh/M6kJwS9fgxmk2JU1P2JMqUtH
kSsPrseoHv9pNfhZZSUnoQrf90Q/1K0nGRYV/Jk2YdD+eYuxdec0oYuBOX24
PPNWsRb1QADJwuAR1sSMHy39KalM5VqS6wO+Err7VpYE/nX8XM8yAInnmJh4
CwJnAZ0YVGqYW+t3x2CmYGF5sji30rUgfs+WVJvdzMUuLgYTTCgFHxs/3iE6
LjQlh+StjXqzIDtKhFW0pgtFGT+QLqOMSF4wci4COxheb0KbYX/ZVLpF2q9r
LA4JJiM2PNs5RHGMDhmAxDBo/XJ5tzjGdxSkyJSPr9vUXL3IwrhIl3ovpcgo
YXRhpEZO8whymTcKqO9vJof9ONm5T2fyh8KRR1UkSf9BPW+knSFcbT/vH/T8
xpFxr0Sukc0972sCLmn9mHmv6pi69ls4acR43XnaEV/UxI41dklbKY7Ynvs2
fjG3angAVftCUhGzmxF59RBpoBeuiIULxIawQAfeXwqtwg2ERezfBXmgrK5T
5tS9+CokAyDy/svddTsGkGo0t0R++V6Ddr3zWMwf7i2DotDXk9t73mtesdXe
6i9S6PstwpEY0Rzta4h4qYKTiOdTKQoTpQ0pn22mh1+itmgzHueT4Xy2crOQ
nXpkn7kJa3846TnsAXxCe3jMoGHlRDS8yK/absa5nhSkppp75AnUXxozLu98
KxXh4n0dQHBHjw8GqVus462QVS6UPFiG1prZZQApGzib8UscED86mDIoAC+k
QwFKxKmQp00gar4VBVjSYj67c8l+YtM3VmDy3dWjc36J9yxSgYpnHuFeNZvk
NJbAVYteuhjgdCAAOQtc6yUyHvGB57xnOzT47Dbd8jR6XKzhMDGTf86Q6hWS
wkdWauh+4pwSWURK7ZAbggnLarUSKqV5b6qBobf4aK/1gsjXHK5ieYcuwQ3O
fqXlQNJ1+qqARU8bklCb0OdFV0WE3cxewuKxZpnE3JW5g2j7nR5BC9YJTtph
M19rgoNgEAnOky4y0X0Tia2GsLOl8wCNIkFOyqdvYV1Y0yjDGf2x+x0IHa1K
h3Ory5WYOpFp1GcDcsmqzuCAcusgCVzNQT6F8RSmTKJyJ+kndB/uzXkFMeZQ
AKknp/2aLn8VTvAiTmDzlqjQL657cMlcfyLZsY1fKV/Z6V5lflabvChWJnUR
R9PdfIE192oncgKlWhCI40qUiCezYK+EDw65o7ethaBuTobwopMP/VLqEUVn
JN6U4ISexCtG7xlL2tzHv6SFYc395vG26FgKh/1RBcZ40quIPhpezJMzY7Gi
ql1pZ968tmUGjJkZZ6sgtQ4N8j/ZoeqXUj5aXtdueT05KSJvhIQu6jcy51JK
RJBU+XhoC1dhYbkSW0azI4CGlVDRcNV3oJQkMRI4D1USY4DQeEebgpwktbE/
JTOi2LciiFXsKfYQw/fsIVrV4cn6WL3y5ylslJtQdAvLpHHcMdwZck+l98WB
fpcIuup0HhYs5vsVoeTalj81WvB3F43Liy/nv20JhzBvNY/1OtRmmGdxuvTU
aHmXu444S8l6nNpV9yil9T7OAsr8d6+QlR/CfZohlLXRD9OrktnZyRa5x4uh
u9cB8aS9cPCd5f3/3QJxi0LIKJsfFB05HVXm5Wgr2JKDVwRVJA0HiCp9BK2m
v5vke94+c5nZ8pDtbReMLa4b5LPo04gpcwK7pe8wmp2V1BHtHEJLwwhvglMc
lNeDcMTMoHJgBQth6xMkozCxNBllmpT6MUCEu1J5X4MZOdlJU9srUAf1nBWq
iSHWyVtoMpVULe/WCv3sESD1KJJP1K6zp8hcJM9eoKpBtx9fWCMvXpH3VkfF
VdwaldDPhRM7Bf+LqfAl7wOZq7RI5MAIjpMDdoKFSdgl7OkZyjHhDvuH5MKC
OEyCgxA1UEw4awx0nR1hUYeKFgWi1ZqPIaXjpJYGBHyas467+fC6bziNrrbo
wqQbEO66+Tq/AGdoOcaDCMuBG9G1fMSPkfcTAtJXELvqNWTF+U8JWXfz/jK1
ikgknTKY2hw1xD8/KNJIkn8FXKoFBXcOyLcM1aTrvCReavmdGEnHSUnLMovf
egI9qMq5wGU7ZiHHe5CVaNrgt7tueayzHTlk0Ax9/+2rDYltiKivuA+8M1QB
Wr0hGcW/0E7SOEelWLIIVVaDFOFQODrWUFtTn9CMtF6ww7Kg2lXkAldFw+EM
boomeudMUU4rclZWJC7JMPNyBcphT2GUFiKH662I+OaBoKxCL8+gZi8PCshP
wltYA1QXf3pNgtvjNg00tBbMYoENPGmWE7GTQCK/1Irew2PuR+IWaua/akX/
jIXEGlAuGtbCXM6w6Dmp9Oq7uU2Lh6dH2v63nBOdIrADj7sqjSxCC6EJL9Ns
PeNa40PH8sBnrtjDT32u+djgVBriFapRoGQQyUqBmJoYipTEn/AC5y6N8Ico
LcMFdQKSatddUAjWWnpgdqUEzL9EJGEaSJK5QHp6hscG0GSqogPhf+un3XAB
RJWnQyEI9cxR9Ymwf4o8tNwnNZoXIwok5A8lEb+RX2O+GY0X1HixUo+lDnyT
WaWKxMapz0TgJFDMHXUjwhbIlOxjCl/478RPO/X5VNABMSlX9/OAn+ymEtup
XCsC8wMx0R7x9gfuN8odNQtAI/Be7WKipNulpuzhAWkrNlVl+YTIg7C/J08v
MnLPbeaHBSZl57ikrDfby6emOB53pJiJ7JK1tNp8d3vDTe0OVo7fHk0VipgP
mQhz5GBVRu3QgSdJPS0UzoYOl4ToIg/VUPTXpo0RFAckuVOZi+VUpUSExfNG
gFJ3UwF/KGd2IfwChroyEeXyUGbeRscbTeUaaVMmzZCfVpmV8QlEX7rH1MZb
0m2C1Dwb/6TvElUmv+OZWxZK1HHpvoAvbJn76dneWwbP4QAeeaFOvDwPgxQ8
pDgBcfgWF8LFsibwFUPoNNiHvCo0pqbg8HNsVURsBHubZC585s0Sekn0ilNC
l/WLb31Lm0H2vzAVBlfG+0APl+HC63qXcjXW+oSnEPPvDfR8jT8ZHbteqKe8
X5gwZcP3BI8ydfrjI+kPZys8VJOoFSfZY3637NKSHS0Quv77VzJKR9LfvtK1
0XG7fUV+AViM+xbbAhnHSJrMPJ5LOoob8JSdK8jtSLzkq6/TpV7twFO29ZSB
xntNCWup/KQhfMeU01/bMgtd4M1Jx7k6+UkH+hKde/0e8ZFu4yC4eH8oRjrn
N3+uvKNhK081Qhmjv788Us99GWxY0GZlvQQRt5uenFjHJA1mrK3QPgn8IyVu
5NDo9gmKg7DzafkOcYYxF8XvCZ2gAoHpyQapK3gvyjFeXBY1g6O7rIO/Zyqz
Ib9k1LimWBCmhCWCAWWQnBcZ9bXntZIvErUNfAOTDMjt/zQPx/HN6A6hj8I6
fCLPdTOaNViI+/ZnweAgyVXFkT3l4tHSnEmyErW3TjtCozzcLScyQG+UP/Jd
CHG7CmduIkb2CRLTRzQZPO13GJHjEaDT3qhD0cL9CKDCG12kTHjkkcNliRpH
oeLthSXZqegohmxfj/JkMNsTzVC8PRZ+PitDpCY+jIhnPWpY+HH2vcdr3eU/
hhGZHx+CTEaZkfV25O5AugStLgTPP1es4ig9J0Pnfw6xAavc8n4ARpKiYYtX
PWEYF1DBcJPdG9JRcJ4CBOa5zdNBMM4rtkXLek0hJ0RFVSPG3Mx7dVJxv6kb
HwU9ClX7sdCcY1sSQ8RNEO/OE6ERa0F4M0QyOQ7D+7ZFAiRod7HvhfCl14yZ
BCQrADYtiwNMtImCWFbzcA++rkJRDAOiDTL0C1suk6JAfFajl/4pdUn/sl10
BGtHg+kak1tRrUa7fz07h1cZJfAYFp4v3+KNIp7FKO/VHBqWqjhHif/BIowv
LIJROO1uodInbDsfzhe3KUTtez5QWPVQ9+jODSPqU7NV3qQq/y5N6mRi5fWk
WgUoMLgtPveNBGl4LvGXoOuIHImklyWob0j95AGOBsrC7MvCkL3yifc2gfWi
pBVj9VZZYFL5mf2uwDTFRO57tMgh/afk1n1wPyUViH9rSGCfCTZEIdEib6Ih
SkuQcSoLloza7W/vUMuCuCBk2Rw+UWEuPtWlO4YJtwZRidO2cGWxTqEtonnv
5NW1GgdhBDTREcPDL5wTL7z2BLUGfYiZebuPhLTM8A/vW4x+7yqYj9UoZ6hh
mhp+OqoGNsPxr2jIgSqBjwFWgSpJ8h5gkVFBMBxeFx7V/VKPzkIjXwb4HMEM
FfEnWRdOkrIw1ZkRwic28rH4Vrz3XD4qurCH8IhIu9TbH6W7vS4jvsMsO+1z
m2D/htulfYXIZL560KxJtLrKccBXxHE2aZaxOupnGdg7BmLL1sjKX4D8n+6h
elpPdoHFOGgp3y60CgsFMM5SCUG7Aoi/AAyP+HpXWFsNzBPsht/qx/nlcAbD
5NxuR1M6UQ8TP6dTp1dLr/IKoS36ChFM2qfoLnLW9Cmzna76MYT60mnK5c/k
6C/GC5al7K4w9BZ3o0miepxRS3bWEbAzxTbJxl2PSfJuTMjNX/MXJ6rdT+ma
kCxPE+EdXJffnWsmfL5pDSEJ2gB9njTZM+aui5YlQSmy+AgkCn6y/j8pHRdY
kinAxCuCPbnr1UxXxj4/7SadjXTKf43wYYAoPDBSCZCM5w14BBXAT4/Z2r+B
pb/nRAtFukRHHZxPp2ui2jmwRIPUI7NBN4+A8wfEB7+XvezdOBNIcByk87fN
Ww9sRcyGmBg3p7kzVpRuIdLBDo6biZjfRgt8GwtI5BQN5GmAxPbXUhYDPzKg
7mavMVehxWHrIEO5On7mixQEVAIZXtGdcBENLHTB7HzTcsWOJcXuE5ZQKgwP
ADeXpO9/02MhivARX+cqXYvS445LKr95LtX2mtvwjuy3EJ1qbabPMz49Q8XW
cItEtMVewG0m0rY726zf9J7JWhl7SANyOs2sCwIc51YKu6MAPGnRVsr4pk39
Accx3Zs2pCgSK44FHMzA9UoMPmHWqSVtownkwMzfbPVoV9bWIwivDbJjACBx
G1LrG3NdDTv1QElASqkn/Pm2E05mBk6PkLr26EDA5R3+EsHu4B6R4euxelNe
ZB7G9Bj9NkYdCi4lvOA+3td+AIQ0SBfpFzCyDNx6hdTQb06b8bKiWWRzrp7P
sh24s8M+kQSYWKMEQJgVeIrHcTeYk41F4ynKX9on1SQ2VC/wzJu0JnDASlhi
QCLfssjU6kQbendiMcubLNqXmoelan8Zn27MlOMRjU2gEZeqqWghnHUCgUsM
BjK+jOoT5YZvi6OEdNaocMJq5ZjVPkUlPyxTU/2CrrgBOSmsb1Pn2d1TU/xw
txeVdkv+N6Fgg1MdCrQGzXEowns4y5A0s8SM5uhgVTJQk+Zlb+SNY/UtTzXQ
EdMljyB/e/Xno1C5vQ+rDLS9VTuT1Z38rKmwWRm8Hy4V6h0tJXEF8XkXDbX1
W9VpE5R07kPDx4N9qsjxIzdpzl2HFuU+U8m4isHHu/R01PotqCPTIANPQ8oH
7CdN2PuZdN+Fz0hxlzt9VJy9sqnhIVWLea5NM2LkXMw/F0t4HtNlyIgpdO9O
5EIbFk9UGxB77o4LdTdNrEzzXIAa4p/IXDx63dsT2bQ6PixJVBUWXRePCkLc
VJjZcdziE8uEMJjYP+DAYVTmXZWtu9v64l2D+GzdV28Zsh3XbUhUPu4SnGXX
oQsbiGFifZ53+Du8WiLEpMktf4+T7vbYvGTMPEq0AqZQvzlfLQJqBpXegPJA
kAGbk3K674XFHBvXxNU4Qon8pc2yJXYk96Ym9Awxl5fko7cJhxQiYQSZ9yVN
pcBYoTzK3NyPwpnlggeR6rgTJOkgVCouE+ORxrEYFKpCImYW26HYYPGahXEo
hwLyrGyMyQ2HcTpqF6FjBrcn9FLLv8YYLCLu7RLLjrhmUeNe8gaCRsfP5xAb
CoBq0hqoYYmXEIt4ZC3XLXca4xl21A7bEmKLfXGOfoGaVi7sFCoB42o2FefC
CO8zDjB4tbqvHp1oyr6JrG8XwMELs4SygVx8g9R+PwSmhf3kVLxkSKFvrJPB
EATynXV3pugnwRF1wtJyU0evYGiA/VkrFWyz8wGC65Ax2KUxHMiByD8ce03o
EOA+L+wYL/MRkVAYz77PyI2RsIL9QJtTS5IG7PjrnBYfnJbFxtluTXaekU6A
YD7mi6GxQvyhS3Lki+7kxzO8jfIgxPpXTimqyoOnZnQwOQqW4j6ssd6ayDx/
5Y8/sS3lZUqiIAWmx3bINXoxRksOBl1Y+z7XP2HFn0aahW6Eak8sl9WNC5wb
bkzR6qkPcBTcgxzdpWjGyUEULygA7qYfcs7cUlcqzuKY4Fb4tDxCBAiGiGgg
8t0KoZsPY8btS9fwfWScPKBKow+LQrnF5Wn9k2Oe0TEL/Kd+t4vO9WMkzavC
Xmt5dRGslNW9VLO+/I2yBo2vycmlXuVqa/bdnrm87elhwSTJfbPXcn9LrNtO
Rq8FsEkYt2wnFH1mioOB4Sif+HK69Bg8dNsaSEIDRwwGXcYqN2HShG3jCK8T
+V1qcvABpRP5g4B1CCe8SSlxuy9aEDObn0WdQQdqKsuxUxnhxtmGKCWrS83V
hhcEQln+NiyTpiVorjl3rRmG4v42kyoCtB0/U6Qs9q8VCSREvSlg0yB22dI/
fAFryeUE018VgW/nHMiHB1TKXDnELUv+gr0CZRl+MRP4mIKRRupB8ywOX4Hn
EPs9/cpX9IKVZZXw4JRH1w0Mq0ozQdKrV5ByhddN0Y3tW3uJ3z4NCEk7EhMv
Nw1kNDp26EByWde+upwZqNX9IIs/Sq+YavZhGxVzP64UkbhcepbqwYkTVAC8
rR1NF388gJmb4K7tng1dEh5rJyK9NH1JTwN1xpQVOi+bYk6rd/UCcRmPjbPl
4B8E6GICMpwwooOGt6jHNRXkeRPnqlFAD4huB2d39cuLufqznAU8Cg9WQbBE
YAkDogavE4D7oWYbiC951mWKouuKZ8qg7mobabC1vBScaJNzhA/4X3PsfBQK
WIS8LPrAZZZzSymYr3G+u+dwVPRA4OPz2qiX2YOtzhjd2DRxcGALkZOoitsf
XtPq3bljDdNnbgo6fGRtvFZYfGh6H/2eatE87t/7ZfUU5UNNyHJT1Dg2IAm5
FBOPhVAiVqCqARjaDKBe6IEsYMs/Tdyzw/D9aZef28wC0VuX3gQOfcq/KvxG
rZRVAFk+Va8EU3+L1dSoxHnzkr/me1zezAgBdypgEb0AFypuV+e0C1IPtG2Y
nrP5KJpmFtu+C2wMtdmPkZh8QfOzc4RTM34R3dXKaSgO/csJak02OH6psu2r
bUG3hUplE3IWq+L94qqQ/1MVKBnGtY/EvqCGVN2DZSy5A0l3gBaoGkjTWTBk
jY1Q4Q60O8quHUvkdZ+F+oYqakuJ02P44ue8+4U/C+Revg3ngQHHhvY+NS1V
4pxOgw3DM7M6AbD8T6uVAAUVwGHZlufVye+xiMKoe5MlO76lYhQKw8cI3of5
iBxmwbGpomxJxNNjdTUMnwpDAxfbfbr9PjGiw98dGDiFqdMZz7NtyKryhj3e
LHWcar5Mcs7+jNLDLXim1npJAaimuA5LNyJVvQ4Yt9RzhztT3WFPqytH34Fw
HWj/eUzBxDEnpIxlyT1zeRX5CiMhjBZPN1xADcsk+yqkOFkFv5Qh4dDAI/UM
89EcPp6UynTNRXayz0LBLLpdnsBZVJTFrOhlxDxbUaSK0iawkI+MD+M+BM/x
WX/B32EiWKeSoUdEEUgWD/BGHCuM4UBzcjptuQgJWwBuoD6B8us1DfxQtbyd
hsje3YrOnGuQbcrI9JLhymd2GMVYihA4LbT0IYcM1+PDMQb0AxvnWS4n9iHk
ljJNwV7EdbjnlMnRso+pkyBj65Ri129f5nTNZ7glvFWmoLhsvXdWVrjxMVND
1T2S8HqEQoj0L/0yt/1sEEkgtb+C3e4GT82CJB/Hmv7y8cid4wgB//7PVspM
Gzz1J7CNa4QNQDBPcBxVbpnPnl2FOsVEQK7CxOEVyA0wrgii/89DKi+QlgVP
PUiZmk101YTlo+h/SRA3EBtuTIlTr/JogYvoQU7BP9mzRCTeQG8/UXBtAjlc
WKtgM5L4FaXsZcSd+lr+kQddiYXXlrgfR1PDjvW+bM/BMeB6YHcif6PODP7H
LgBT3tbMMlPOm6JmwAPpZGfutyAVa7cOKyCskmWHxHYXeOXroSPJE0Q/auiq
dBt3rkIN92JW4zwN4ZFa2b+tANL9D2jSDREbOW2CXZU9WU5GbTlDETHx1ovg
cHEnh+FPWSMdl3IjiS8uujbso010+S3QQzcFz8uukF9bCEmZrD8XFcqIdhz3
8CND1XoL0x9Bv9Elpg/OvcBghLQ5Z0nr9q80dFYkjwQqUVRwjU6mrNZPwjX+
YsXt9KfiYZyohnLey7C/27eoyqKVcPYQGUx1wSUnsLFryIqtmkSr+zaD9NJg
zsbLezwozLdCcOdTOECRSaXHp4lCAKUdbE65AeVWx5MQCkpYvr5zY3cftRr2
QQw/pnuIWwoIUZQYTQisyM4Utjqhnbsw7ZdbPwAgclJFxcQHP1O16ALrQo6e
ZTMKr1LHlipJcDMZJNAMYgSO0AH1VfzF9OgoXfRd0npKW5azdUXa5uzVtgZZ
zpUO0yYtpKO32837YRZhWSFl61yyjNx0ZUQazGIW3Lq3TLubtRunKKygNNgf
6Ne8UWofK81jVn87WlEwq451LEDLJXzMY5RNLj1MmXRBxxmwr8pqMCT2+mGs
VLpR2bCP3cqwLURefwBLJo891BkdvkFfyKGTcaxGpcV6BIxuJVdfe6SFZIco
hgT1dV7FM5dsl46S4LQuMjm+hZR0gH3Fna8g/lFwJlnpckmrueHK1/Ca/gh7
O+TZmec5mYya6et3AHHCD4hZBH5BaONqBz/cyjb5eeX+47sAvZ3Lo538ovbw
DR/VuFt6uRIVjBFyx2syvBj1RJJtJVFBsSKQ0P7r6KA7vm7laLJ8TGumZNB5
IOlONTXbw3Z+14m0rJlQIROgtOv3ZJoJPc/gdJPCVhDIBrBzIMR73E9XBdx5
NeSSf4Q/gQJVqG8M7CRVJgaid35ybbTPQiIRJUYQWr52oFge9g6/isDeCf8p
XS3sGKaf7B3t4ok+gK73xatygGtuPZcLxE3LP4/Biofh6/H7KbB8AhPE/a5F
41pHm1LwWYd9wtQeSShg7Gwh5S3XCqvdKnDcdSpDhGOWi7MrVcvVFqhMMPRH
RqAI/Q6hJuFRoVEz+tCynuOsvAVxQmAeKSxOKXq1tsHzUWVBqR8xFWkySoc3
6i/0k30jX8ezn/c5sNyOVGKZiWyMzczxvGNP8S2AOV1Z6Xk92hYN0g54zWKi
cxicrViQMkCIG6TmyO5uOK179/3sC58DZvByd0NDaDZkFbIVMo8/bxdS7lmE
xszPgdU0xER14X0tojSrxCkFFnUgsLdvJNTKh9FIBZYGaLLwDSK4xNP0K7T7
Pe9gRGM2wOuma67GbOYVUg0/1HCIp+vEhL4v27UGrDjB5rKnWqtBYlAqhbm9
uLgYYVUQXVeXA+hlBODNJNWCDOaJU3mHkT4PKbEvYUJxU6tqxX4wbz7jN2qc
6rUMYVmUaGHtDwd665nX+G267FxV9rL7EOJfBVAcV+DqCDzOdL3+hm1oMavL
UhzSctP3Yf0q7kCLCkAsV+U6MXQ/iI/FC3cS9DF1SkLb7ASwWW0gJDyqKl64
Bp2XvsNJkXbnAaQvKl66x1OLyC6ZEzFzEt6YNm9YhWdfPt7GqRBpNy5z5/LJ
/V9b4Ejo43IXAx2SLQthHqH5ekodyM3jrbPLAl4pF5H7RiAAtw1xf3qtOt5E
b8OOPay+DzExMsKP4ZBAwJTRaoVXcyvu3JzFlDV5GrzpEDxy7LurXdV6Qsbe
W5AMwtyLUi7tSGcMxp1rAwS/w3lI2GcEimtLG+Dh9/mNFaMHQVJ4yNfAc9K9
WWoo1WG2Qljxw87zgpN7G8BBMQixOXryhOeloX7Wpj4Zm+vJ55fLDTx/+XAJ
whYveRvGVwwP6qjnjHaNuzqFqtq8itVyGHcN+8+O9/YTQjoBAc4Y2UD7w1aa
MHsDkycZcCV3bzXJkuouJJYPWvOfSH0t6yCdvQQ62++tLAe/kGqkt2HyBq4H
ojEnhYnJXTVyuL3vMxluzEz4ICDRA8fjzX5sL+yJ8//Zdy6PP8lXsW0GoFFm
jA4EDD89Av9uK6eMneUrNFvU3Ng4DR/DPR6D6zwTeSkF5AXXSrB84OaIhf9e
af8wB37vOHPudLAskcvMUJa/f2sK+y2qyTtG4pkOjCpoiNrYH96TXUziPTiy
cxZrTq+im5J4bLdRD5Wqex3CFSFz+nq0LsWFUCW0ue7wEDOTFMY27mJcVB2p
PYyN7I+xefbYIgAqRx70wsFBmPf+M4FzL4raCGy+E1tgWU+Gjqgjxup3kaV1
b5KRq5qSmoNU1XPouq+OsXJqXF/yAWUR3DGPZfwZEKzTztOqQLVJ8myebIif
v4Dy1yu29GF4O170P3woaeULp3Iqt7wk6a5gQHhBltDSRf3ZRqyqwnDxZd5u
JRTYlRs5V1pIoHcnI6bA68N7ZjmT+y6r7H8dmhz/cqT22+6TvTDSWeLAetfO
x3wLgBLZ28JWKZNMvSlz4milGtd5Q4R5Ji3k9BnU4Drfj9K9kSmtEB/dFiUt
6db594Rlm9T+eVuEofNSZfFL5GdukfHz6C5ZSZxE1508J+PYmJBTIxEj6Fwv
1nVq3iGmDkQ5CChTuWmSiQLOkKGsuCGtqqj5oCykmb+pH3p7QhsHIKw8nLIb
akmMeu+rju2Tdg5kyfpYF84NojRMRxd4kjbe2yGDNNmaVh0ft9wtzE9cSK4t
YHvxV7RDzqwo9bMxAgDOvUgkU0Jvpgjg88be3jcSUF3mVH9Mi2W9V07rLAeH
4HTta1BMaLA9/toLkeVMXs1mbvIBFlHEhRRgXD/BATMGJdFJSZzGULW7DOXv
nPL9Y2FdjbZrAsOP5/1Tzzid2klDL/j7xC2LvZ56XIAvN/xEk4fmqTTey9Jr
ApawZ3yuJvjMjqEX7oVK9aCb1bZMUpNhSKH06F3jfSDLArTuoEUbW0EpPdD0
P1F+hS+zAbU1wrlEucJHRK7hTT6JcC80rdlkeNFabylpAf0UuldfN1irBODB
o/wFvXoYu3DuVVhk7zBGmJFIvmnE9YxE/oQtfM5IYAEWPDTn8X8N2j/POTdV
8eY2XEY89xVGVysKV+cMpw+rARV+vzmJ86yEpbjzCa+G0r/duuZpSoHILpj/
IrcsdxZkG5QXwXvrMS0o2050zgxqUgtiaQ+CJT8jUB8yAXxfjswgSeeZ2ysm
MdY1mn1rjJsMRAMPHtM1gHnzZBRHe7kgeNjGsHL8R14hFBWNEmYR0HEE9Pfa
F8lxcHN5gT8PhztSouTy19ZBWAKVktzSOPiNLmZni+N4oS/APstxRkcg13vv
8us3IyJHPzcKcxy5t+hgDo06Fwytxz+xnC9Pe9utVECnTty/M6yNWc9qm3nH
JqB9YUkrniEf+br0GpbNMk4h/D7mkBDI0s2Avi60jK236Bf8g+UjQsRNXpU6
SjYrAM7xuqRai0vwzBaTCipGLdiJHFjmAsZf3532dGEY7dEeY+jaRX/IVfPA
pa4wJqVvyHug61weirQeiCzkIgrOTMtaG1Zp9p6cRlJ+X37ZCkjClHuMwz+3
Xvz/tXBeSC5GTzg00V2lY2MLg3L+sESvaqCuf3xgT3PzyhcJ8Kze2H0H0ojH
NGmwT/Ie1dT1pcIpSSYf1O7DK65VTs6sevltfZPvtWC/An7b3kfQLszUSYIR
bbQ0ajOZvIG46cgKlnHfudfcDEZsyQf2AfK7IwcK7QqkZ2VugZDjMiSE58zM
caQeQO13YXgQ8GKiKxtEfX//Fwa8+4pEH5J9L0yqqFXVm2kzz8tKGARlWdt7
sNxjvEQngRDjI1I2G8zDMBGmJeu1GPxvOQoYr5YQ9dfAYXU/IlkCdBi6O6S7
XEXSPm/mQQNm4hc/InleZU/fgzMyRc083nq3X+tZCSo0/J90SjNykA/DOvTp
62DasuEPOL0tOxqYxZEZdOPyDpGUn9MUEZh3Z2/aw/BMstlNdMKMGfO9egCQ
AWLz2Na03R2T2CxYLsyy4EYlPw7KSHQhLgk98Goh4QSsWRUXFf9hbfAoqF5F
K3CzyjrDeWYqllhdxiIUN8b7oS08V53n0SlgAHPE4vKKb4/8QsPg14lwt8Ma
cn5YN9vodHodAdbV6WeRACkhs4FaoynrUPZulNuf9FTeBoXsh3is/8ZGbTrO
fesZOvy9e3JHZ0J3v9qzdYu3mVgQIedGF//Hvs4M+VhhxxcntmSYos0Tzg83
Vc92+N4KEgTKpGWrneP5f0sXIChePtlN0HKJsQUSiMTn4fBrQrZLZBkJ1qjD
U6x0mFuZDCLTh+IhUxmEySho/F8HkNbz8uc7QRHi3P1vch17yR1asyptT5vm
4XTJXAAXoZBR9vKVGLZV83k5uDuiKv/ocoR4U/KjxTEM8OsFU7W9yslXBPbe
Xyj8nTxNdlG1cZ2vAWwN98YYBh9ihepWQ90sUVgIn2d7piMR+kyp3x/Ztqq3
+B5daL77W8mkaZVIL90tUF6tQ+9Lm7ZuZN9yyaKvjRmFtFw61+vSNX9RPGdZ
dtwqWqtywPA383DRgPDGfrnNBacxZvxyNeLfkxZISDqXo1N9kPMOgbANEsXR
/JV1ryfPJVG4ykBrmwKm/y0xgVSMGuHMdQpHmgNjYW1AHpsgZ7dIdvDR6GFO
GhnrAT000yu1ejau7l7BCbSLkJ8rnwLxz9gUKLlskBtuyJ8aKHCsk6c+2x4a
uDsyUKewmb2NNEIhbWQoRzt8fGhgoRtBBdnJNQRCnBpLCUhr/ApVYyovTt5U
7eg1BhwG6jUI1ivkHoHcT8V+7jnxwIId8udbbAJDc8mcwGvS8JBKuEHGB7I0
uTvPd1Zm72EUOISMOz0pG8HAoEK5S5g/ww3Av8DcntL57vrFBs+u4PJcmvV3
jErVhHiqzN1YaliHcsovWVsZfUlvfJWvInqb3wlmmlq6lhdyc7tSsm1fClc5
5YETkUA4ttfJzl9OjacpyBPuOo+C6luWOodQCGRjLzrc42JEtc8DFSichm+3
9tKl/YmLluNyqpFUuEZCuH/uiIy7nFL+IugHBDLKqEtQV+j7WTDwxAOdQOt7
iqwLXWKjnf13qVVfp9Cz4KzPQ8T+AnJ7ffXu9MGia9YFBmePsleTCnqeeEdd
i8AbEtfRx2CIukVJ5dG2sy3wsqumNMFUVSZdpYegPj3nnlNQ6rgygeYFG9Wh
M0Fi7+lrVgDzcqFAenwQPTRmHrBlONEl97Y38okBfRK3VHC8cTwPLxTi4Wei
IdRxCeLOU5teiGXcjw0auXCDNpBHyTKEthb2Te4EkfCQ+8ocBYM1dHlvghL6
qRm4t1bXEuR1UNbQ9+4/O6lyrAF8Z4Hv809it04yfAXZkOXuIyADawBhMbFv
QPjTuyfkYvDPZUfOxpRqPHZ0PsVQMbCn+8BcY/HHs9tA8FjQmS+6memOesy4
4VJGoe0OoTLRqki1xU4hq5w/VkArb5pww+rlW8aamTigKAnQ0BIVakr0T9ZJ
Ayv5LOebFwhhrSf3v8TlA12bfeb95bHnGlICtO+kS77LsgumkgYacRrO+FiJ
0wTEoJEJVYYcTSqCs18l6zljLFsvhSY3Kn9+JXXpYs3EyGQT5SgmTnz+Rprb
U/7g+6fzSqD8unMQ2fYIowiP1WNessJdXRroW5S8nq54lhvi6l3jNXshhHBF
0O3Bg4pzoTEw83XUG3AWfcCBR3exHGiS37qeZM1ggJi23EWQ2ml2dywBO300
NugkJIr7I84sgWzsW9tVRYUdyrDO/g3np44ZCrza+nCeqwReAlaug4Km2M5n
TEidCDuZCx75+ABnE8enSE4T12c/0/I3KReEtu1ao4EFWD1f8M8Gc0gbSkWi
DxWaW0l1r4thWgM28wxzFL+tL0EjzYpADGanCsh03eA+Jatde5U6CgMSL26e
Y5F6hORMEoWMXrFMveuhOiYENIs7tCWswcZWlZO9jyk2PWjj0Ro5DwchR0Fp
ATMp1YpD5wtkHjSue0R/2n2xOV/tZe6DSc0ar4oouHWaP5GGQIGfzeOsLTPi
pdiGZzOjgrR9U0CwrYcqS2QGTleb2lTPNT4fAFEg2iZH6uhhzOvzwp6/RnVO
1Bh0A2MCkhlhL/+WMPgO67a5A/ooxii2kXnh9fBhHzOfCfo1QgtEbhkFwRlx
7ab3wVTP3h7udk0tr4HhRAlh036vEqLpi4qIdtqAC/8tF5wNiCPSl2Ef9UUF
c4bhGpza1fZVETjpLUbZD3xxKXS6karzUdN91KdpfbhCrB5/LruEp3m6DIhU
QyKvt5cs/vsJxhWjvWCVi3YLFOBhGI3ZEqEiYdjX205pivP0GepP9m6MvOyJ
JlBKPfKpL0wXzOF5LHGdypRLK9x7sJqiqC8Omo4/FD0f81rJxujLX703nxq0
Sw1bShy3oqfx4zEnPNEW3pa9ghW1Hc8Ungp6K4Wrw+byWSRCc6lX7HdOhz9R
iyWXWqQ52/EfQ/RSHWgzOgCO1m7xQsHd0CQlR1dDZHxYMo6VRNFIMw1CkXT+
ZtTQADT8+kw83xvcb9bdYPS9dQcwC19WreK5aU5P4jkap8AOttqzQ3e/I1pI
2s4MZ6z3QH6KOjpwHrtgsNcJxaYPe2X/GW6Zsyv+gR2zu+qdwi45jZ0GFjuH
oR7E9ZsQU2HaaoqXx7M1GW0pzoKFOaZAhDKee5geCOWCS+FhW2V7EcRKvCmV
QiYzZ/+zrOSsuzMmL5eXX0vQxRL7TvkvPLj/Qhl4okE4g3o4c7lH0JY0ISGt
utppHFMaK7otMjKs52cH6ECH2NcTR/jEZIY71oGhGQx5KVd/W+GTIH+vHQbs
0A0DS+NPZKyJLvKcD9IKAVxQJkdaI5oqho4M0lGvUXQTyTrhsVCp7697taF7
clLa985stZq146J8qPCYIoaX2NCXiHXAc5PaDVF83l1/eIJqkkbe+pfZr/4N
KnqVzkfDxxXBkuuihIf+J4fVFi80pXXJV8gc+FdntU/G5LQpuKmpwOu08rXZ
CORbm6vohwUsiLI3ygG3twEW6yVdonxr8BXAghOrfArh5qbDPeJtgWGJNBzX
w4O7HW+iWLlBiNt/NxwgagGHCsNML91dKUWnsRffljRu9KgcZjmcr2EgOXt1
X6et8I6xCqoMuvwUcBQUJU4k+iZ3A7HpjDmUKYvvTWkxM3uMPJXCSobMMUOF
begKdiaHWQp1iVj1slqgPvVNZh+DvnEZS60zOwDyvkArFp0BIdHA6p4V8u28
iDanW9cNdxsfOi7br8jfIO7/L0LygyJozxnsnnoQa3pR10VHwm/8ktJr/PZ3
qbm6kIta3Ard+nUJqNkqlqQnGDrzq5jk5PM4uljgbOnK9xKYlolrDXAacI5s
A5Bjq1jT+cl0vRmbo684jDX2EyFHhx+CZ5PxFQQEYqyj5uqg4RqMQ9ec52xu
knKHe2SEVGQydkh2QHTWtkRMolk/tUxafdsBibZ8tOMalnAy7KZt2gZHbgMC
cbbTf8cY5WCFOujABFD7SWF6pm97OOn2ZakMv+2oL4KB49nL31usDOAuFKhH
fBGGpaRnDfiQeTtWTQFBYuqSxYJl7MfNI6fWHTLfyG9y6FJxt1b7/hH04Bcx
S4dz52qnC+1g4RshgSZBPefA0MyciNa2dD8eSX+LWaWsRmNysKDXwJ/O+URq
jin/KmVb4jwyr0/I+TT7dlYIcDX++4+jPNx80zAIlEJ/+HbzygAzKuaz9cmL
fM+8NHd3X3iLBIIUnclRcWF9lmyFp26g3qaKLLtPKgm9mCLo2lQW2m1EE+E2
6c1Amu2KvvuyBhrt87AM0u1ga0kpq1gfSIlSI9iLKvliSFS1z5k+7HjdG1th
JMA/KTlU5NkPZ9YKZx93x7Bc/GQgHehRTQDz133KHG1ISi+ao+DRxHarifCr
bzj86ebrbowb6FONN+nAMZN/hYH8DlG7zsIbnVwE8LKQusSCHd4bI9i2FDFp
PKjzoBhVs4Wkb4VxnvxA1y+McQimIY258aXmEppk6cdGYSadeu61bghHuhSj
BXouMCSxA8RGP4SJHVbHAoKiQniyk6/pB6TJV1m0PyiYDw/KGyKztNg7GJ34
MmCEsiqctneW1iUvK/6GMyfXlFgsP0cGPBAgzrKFuh9ThrAzWapL1AZl/5UI
Y7zNa6cjZq9pGLTWmhyUSoV8nwkpYLI9ZGvJTXl7+GEevKuVCXFpmKXfvqEA
JWLD+y9idy9ce98ftLCIbG6ME0BEsOZn+rDWVOsKc1wezgvJbbHwwCPrjZ+z
uwQDlIS/fuVZ/5VznbzxZKUmAB6etSg4lfWBjWjkHG1EW/Q8TMq7Aj66wih7
Ypw7FV63WV1cZNfHMaUcraNe0WWatOYmRSGq9+byJXDuPJDuQVps8QgOYPl4
OGVoY2TyuyiSBP7xZG7LIqOCrjFsFGMOuza9/NlasUFoldh3bSRwSG2upXcU
PQyq2iNA1e7WYPr5MauSa0QEE4GWtFK0GcrfoYjhW1UUGU9FG7dWSI2HB1il
RBEzMVh8zOFHurgtBVBq8Pz1u7RHv/9+AvgmpewA2sCoJK1ciJj9QAcCQEc9
+bSvsvH/UipqDtfeDggypEYAqL2vvsexNthHOGstgUCuOlTR8Q5lsAKiyv1q
e1JdIA7kJwS6sZ618wPEMT6rsWhCTn+quxTJD3KItT/DpPmfREKHSK0PJ7fc
zToQ2gU/djRyqpPEaTWJpggAC3yV24pALfuj7aAod66FJ2Dtgg7NtNPpBOx4
kuyBdHSczriNL6RsC8lq1mYAGkZjqbqEZODmJLBfk1qwCUeSMneUIN4CKqOE
EerifWyEbgmpgaFpXOH8EASj5KcxRSGFUQBXtTZdlJm8WWHRVTrYOzhkSTyC
tNrdrdepVjwOCdpaghC4BD7sn3SKvk791d81iV96kYOuxjgBYu4jzxge6dSL
0pLz4ggiVaQlCukrpcioowFiXXbSbXCJfQwDasePliQvxOVLJjOeuOS5TBnn
vt0YUzOeIeNsUv6nHtTNPsNYXS7LFEUJkro9q6i6c+uqVvgB+opAFms5MYQg
cHSKTghQMlDJV3ABoefWLE5js63ok6xwYseAuCJys2j+rqcTut7/cE3rFoON
OEpGr/FDmLmL98yuzmpZ4Wh1d66SFRt7Wp7WYd0FUeKEw8JUGTjmPpbvOWAf
YgFebwNP5B4Yfcm2pvB1iLRkzG3M6wCVhCqZGLFDj00KWDIUh9vhtpeh8b3E
KuMYQk4/9/Aj2bhZOnW6+XXap1xok8r4O5KUwaRCPoqXFBEt5VOxA3tyf9WH
e8OP2VXwJe8V8BUQCYnm2/aYsmBiz7GCmWsWiblMibDmQ02KEgcQEeRWedjw
hC7T7TBYIJhGwOZIgoeceRjcH+kPsPJbzYNPwZdlCRb1mpNo5BKYYPESw6Dv
TCf9JLJd4nQLAeFl0HoALYW2aEcg5V4KmojhKd/p//r4Dw27sRktFd8t7B/P
6dwkx30Wn3x+Ulg83Jwbs3MpB8EMsd38y5nK4uTHzQJai+JoYDda8trnKRi4
q4tRy6VmuGLfLRejsl5nG8XLnX7Mey3hRfAnW8nNL/y9z5GzygRbA0Ts6qX6
CocN5Ds+ZJbrHCPkghjkhoMrXq3Z0lZRGzKRiIgvrHSqws6qein2b8KpvjJL
EGsfYHQaL1nNRfA+rsxMPyTIxrD1uoxVkorFO7bbj3VPJAtWuOmOh3pizYOU
9SmraXc+QQMD5xeGZmwvqwV1dvXAwVLkYDH1LoVY/GeVAeHLLle0YrMqPHdC
p33SaW+3xg6Fc797oeWqiezbQHjdLEQ4iYu236TtNSWJ+Jl4/z8hDmT3aCie
XKrCj+FXQnUZ7GYtARNUVwdVTPPd39awy6HIGJUBdH7xWCcdK6oCwH2+eQ2e
Whoe0cubarjJmA5SiJVHFeDiDvvjEoRGIjxHZIi1QS3eA7NVcPJSAjeG27zk
ATj/xOoI/sRKe6r4UklCV0UyrUq5hsDIM004PlMnr6VVq1tF9UkTHeH19TrX
iNwvqWih8Q8r0z6t43SrUjgSX+sZ0SkXyveYJrMy1uj6rAlK5jg66H0lQTjQ
ITlkvxr0niBCoozR+lFNTpD3jZT3sofbfLZj9Q8DttvHeEKdpGmIRVBgrNSG
AZDvwBlKyu/PrA/itzfKmbPC0nPYdxNXAu0NLHesdT/a3NngcFDafyVh9dt7
mGuKBuDvYlRrXFmf4qDpILn8eeVTHmoeShAtRMYwj6PBaW+wdRHHOhPXIwvj
ig/BqCXlwKuOl56JtJUdwKwmlMAz9w0hcJf3f7kQKBsCda2sbuMLXSNAoyQE
EdILl1/OEfNFLyde+wIIT/Zx5JHTkKrM+dkJeiLmaoO/3kaCttGAgXYlY0At
0sO+fOf3AXQiTEGlCRFtrdQfr2Tay97Ggzu11V1O89F16cF1Te9MZr6PBgvx
meOEnCsahEyXu7rMQEYTwPnUpfUklQEnQJ05SDZfzaAL1T4WtzhFEXlzeLKU
tfxzlBQakG7bKOFP5Y2vbkXWM7iyHOalYNV7AJfwyM37+ycDd2xvO8xH8pck
mhcfwX/WI2BIkugQE5tKPPSnBgLnmoCKbbPmR8NO44hI49o56wSzl5eSNhB1
pTghq6QvsNTTFIhtHuTggab4Oeowk2WP/xfw6HgjBTDr3k1PLm+yBkmGWQt0
lOCVWsVqdd3tJY+NN3uA6UQCsmeAIX2Z4oHoUTb288bBnGNpHAvaBNAFQbid
tiapYmqft/ddavlOIt4/2xdQo2nrVlcyQZQa+6HTDagqzflZVVqbQwgU5Nzv
ypPIBJ+9y9Kquz3rGtwirm5gkuAD5T+GVz1ApLqdZ9yDEQOGVkzopeUugtp3
aZF/ufz/ZbgBCd8vfB7WRb13dpzCvY1HgH7CBv7ZNFe/ipXn4i/RqF6mHglE
QQ0NyruAiQn4lrh9DowS3foR/LYSH8oA//d4erk7RkPMCngRnqFK5/QE7jwD
5UtYjplxMvT5dvqartXbDiGL2JZbK2crn1ksOV3Gh/vSnMu2mpY6cXNOBqnr
kpoG73xw8VWrpcGkoYOkMRbNm3WDSdxAogQyq5wC/gfk8MrdT7jOZYidXnGr
+ABxZYnktJEYzFJpEE2UMv8oKBHwRd5ukqrKYQFS6EtIo85l0W3WIzS+/EWG
OLfMm5thgCGj9MTh8o6XCeZ9QK6zwGqxoL9SFn6rTzDiZ9iwgLkhHeKLe3xA
t6+P9Dpd1tipj2ABm0DF8If3hhxuZtrbrt0UiYp90bMdV36zGI93C1MGLVj0
YWR3UCM7AWNtNn6kYtUlhPclOD5BEBFAVJWa5oRf3uCNPctvgYIWlliMQWIF
lEAdg/JVKtt9tfZxZtGQmR5XQmei+lvQF0xxu2sWH5IMFObCA2gNttKvi7Wj
eH3yCkUwj0BaH2tAJ5HIWJbLnH416kp6Soivy2WzeZXdHWY96+ZAenGjFVRU
wMjOkLplCy1CpPFmtg181tDHpJYCvCDjAkUGoQ4aKZW5iiXl6E9RHXzV/ERu
0q5TKn8QKwWFJZosk4hH2whzTYAq04L5XJhDL2sr1yiAY299gmcA8uT3JUtN
6kQ4ySnI2tlPKM7AQFHYh/7MapD48vnWgWDiKn40rHFsptT0+VUke7Jxcd4a
0hkoYktc67Oc5COmK+XhMSrDEil4Ynpd4TLRPP1ACcHtJUDqExKXSzRaSnEo
oGrgSh+ZQ6mubCc1JKtm95Ie8SF3uH0r5hZvsD0rG2Rv+KpHAUN5/PDv1lCU
B5nNWbik9XconFCv+Py68/PdPmCtZ5e1BBVYCCN5JaPeq5vRSlhh7LlfaAek
NJLTleFv6yWRkd4x8pMdB4aQimkR5gydKOLw4beDgjXBDdisWUwg0hF6y149
eOGSSMjwE01Iw02KnymC9KmVgBYTMMeL4sSsU0BiY4EkrEL3gO7dnKw5J5j2
QWJW7Jg+it/j9hWiclfTpxeU7zBhGfBupuRkrAr4TV+d7IH3WQ97rpsECUxH
bcR9BiiXyy9gRCN1r6pQv7dKeQuIDcgoJSDAcX2++a1Raqj0GTGWA/wlk8YT
SI5XiF9wm9V4UyUwNCleqFIErVXnDgEzKcoBZgUrXLQlWp4kCxj2MpBd4wWe
igpAc9Bk10ZI4YvBTtmtUZGpQ3Jq0Va0cj2KkIyvxtmJkOlSrmrwgldRXzdF
vh2jrZUWjqXWISaFv++hHvTO1v4n8cn56uDdidGZaaDP+yTVlEpeFqk23Fgp
879CsQXLAKI3BtzYvyLbo1R4K0MKbRieubzpqsUqsbcQjCHJgezVL0HY6zz2
mTseDfDQZH08zDysQLPpXhV2dLAPYnI7uoa0h39P8Hll2tgBgR/Llzz/LrLS
OiNhSz4imkzxSEolSHF12lwMmTIwl9p1W6kfreCuzgEjMEkIXtye7dK3vjYu
DJcDZzXYwA7tTAixTluu5hBnej6rCt0euNv1m2sryiCp3AefpRdAlPLJdJ0W
tT3ACCMssC27Uqn/spAs/OJMDb+kr4wU+SskgOBVLbmrna1RAvDTLdPJ5zyC
fiA1VJUoc1abjgMgRt50XEkL4tZ+Rk+U/kvCGwqeemq8phxKCYJDBXxW/xMy
PlhGb7tzw2vRrVsw4ZYbI/3NLuosMoV/tkDNAf+16H3tbgQ/KLDJiWi7ijRt
fezYlc8gtZGOTwFpO9mDzdPwOwpmRr6y4++Z8xmSbFh/uR0F96KxvmrGXTDl
m61/T0OOTg2Ajo0UyyAHrmYjPICr9X5nK4T/18FvhWA3mhGLBzsUjOIrCx39
hRyaW3ZnmCQdRmXGxy2s5/E8yla5jxcO3UJCe7TqTKQAyVUM3osNzeQkeJ9u
yH4Aaj2TJhxDllfSe4rjl3P4p1rWIMhuGeJWEUH5iWPdNqCHZq1iogJ1Hfn5
i0cy+DKIMTdHo4kIezvgoSBzIhDkW+qW7eDTZRHNa77eCDFAc5EvK/3A3lJu
hZiFeToMruBlGnamKqpyq43UKm4k+V9f6MYfCTMBo614ONpoalqhdq0qBfNS
xFMlObwFOg23qtfnOKr/U/aZnWau+nJIwWXFkTZcLLOTApEnrmcReA0kKAqs
Vp+0Wh34rjp00XLf/09JMyJaNmgCwmsv+Jk6sc2EgF99BKqEnzgiW8M89uEp
tEN/3oSsMrXyh00THub1rABYA6n/bJjyTSc4qUtZDWdniFzVMGFqvFfIIyKC
ONs78vSzW8QkxkxRwlzU5qL+2SPtmbP0RMfG+d9rSRjKXVhqQ7rLUOotpWdY
S0UTsYdWV5hE52QgPtZzNe6m3k2Vkr+kRNVQlC4SrwBN+l7m4v+HX6O2uFT+
SFoentk84FKmGjqUUoR+8/q37UcJ3U8VloIlxGO2/rjrtlrc9mnA4tA4Lzjb
1yLf7FQPTao2sXzz+p5zzHRyM6H2yCeolEs2JBMBqM6EiwI73Sz/ePab0NwD
gwCHl2PSsWjE7mhVp3IBFb7PLZd6Bt2XMK6Gqi58PRpfdzHxcJSKQeS08Fs4
Qp9c6MnebzAeh+YlUZEUCRa+nauT/iLFkqJTD6lksciWyYBN99hGZkJ8z/58
8GRpJGgYtm/+G5Hc26y150cVAZQAPkY2KK6xfX11MhFsuSXuJrCMk0cF/8PY
dVwXpIxAbBzOJYwjDRoQGul9EBmLj+E5AjTWY9xx9GN6pnsHLvLPzLnYNEvH
RZVlsNEGf+ehBhjggM8X2wVJvASKR2j3y9AnhlP+PlR1QST6BhOFymKT8PMM
cQ4YaTbsbh7lWkgPWrARjl5ZRimJb2Fgj9V0BUdU+8wN72q12CF8SP/PvU9w
jQaRqi98uLgMIQtssONh+LzFng6Thv3dkYtotuykaOW9lEI6KrLd0Wz50qU+
tz/vVMjPh/8iTn18llEPi7AK9Dmw0IvkVo2Zqh5fE8+FQzc2D6Yor45R2yfe
NylwjrzMXjb61oykg1KcDcaKXk1AK9FDIw1UbFRNFeCi9GwGadqMa0ZFgyky
DJel6rj+BIX5STx6HHdaCjxFQsZ2C4RDHvZx9eHJdZ8xCPxt00w0u7YSaxRJ
7Xlf9WauFBtTP2TNIVccM6m5k4fAii98/L8PcFnU1TgAgrtAFRoAnhKvX7va
lsj/Wz0Nz2GZ8GAV1Y9+OfacSGGJ2YgacnVN1argCF9tywDFlZ8s/bveqdNL
t6GIwVzfCF3nNzbCEy792EPwrAt/Prla8wgqFNR+Rdd+sbDkB5tjy23G1B3V
R2FAOZuY8rVb6HOz1bBX9rYj4pBL2lYfxl4zKScnqs/CKHrPxDL6LXRFG1pA
0ZuumZyqm4Ybl2wgW+LRYkV6LRte6mtFXcnoh4ktkbBPvf+9aWz2NKUd+eol
W8KrrtMEFcK/cTQulYzNSxOHKOzrU7q/5adxI+VbvMa37jrvySG/ABJAC6j9
DPBLsm2hkecAquS5PE5/L3C5mPBexOEY+xO0XOMM2x8Q9JhyBh7T+lFHNbu6
gARcafmVVB9eswIq5bVn8HNiz5JupNPYbL6Sr2NaDkr5+oKB5DqqOIUj8zBY
BxvamUAfvPnRI1vtO4dQUU7JRofAJWOQFk9EBvXWAW4swCZSmnpU4mrzHqy8
276c7wOYEKL4IzdArs4xJL9S48IKNUaxCdJA1IZ/le8uHAWy7+zB6bDXyMKn
zbClHT1joH/33mJrFdzTcooGPc7uzdUWNhOW49ctGIyCZGFC+piROYj5Au+F
koLbW2JBTvO9okwSHZTUDm5uPWV0RmUlkiJJFF3rJ9lP297DTxlXXf+pJDlW
lpFE5Q16LNIz+YvCCRynT2Vufu3HxR8Hzobd3bRpPg8pDYdztI7hUeh9RrCh
tAUN+gVhJ3ZhZgrw9DxocA2GR73+qenkR1dCrhvWJ5aLfq4m3L5u+SPVtso/
i2kLrNnWb94vlL72PrEVOY+GgdyUBNvSjMM1YRyYEHgaMg4e8Sd4bLYKVYIh
fHLFftQBvjM+ippUcTmXaJMFWTgygcjzOS2G6Tu3GWbGNE3fuZPRgFAXdGZn
jro3eJrH0cRFfeqPyNOpzREViMlPCCj9wgtFeTxyF77t3oExXRY/mXbeYpNv
6t+nX2t/ejZOz9o4rxtjF2FK/n+K48ACMP5cA/SLxvb8IARj6Ag1ixoRM2QR
Vq/QGcR3jHmPNFr13HJR/MywgRcLButbz56fYJ4nWG1HKkhI4qCDoS8ivkOj
h4X8cbLgJDuHU1Nep9p77lUWLiVPifczaB15uGHy36UQ75e0Ui4gSOBAhaQS
lyeTrt/MguNFTDcAN+F5Q1nmn1ZrxLJ3sYq5b9XLAVKm2AfFZwO7I5s39EJI
uNETd+Jbmd5uO4/UN0WX2QIGN4PrNWMUensiAL0FHQ/V8MC2eJAG8OQWvWr3
yqxTn++wHQuCoihksq8aK1iyJScQmNIKjZKLb4lvAtcgCJd8Nyc4hC4Ofte4
eR3GNOpv68Yw9xZmeP5Dg8YvA7hOa8IIjbY4tEHNC1J2+BOa+brhGoQLVHEH
5jrPP6iyst8uQTVZH/h5ZXjabbb4G18eVdyXKgL0x+v0qxTNFf/uRNJVtLDs
kcZUAEwLHYg5n/Bk9+DlsZ9RatG9u7vKQ/f2vV2o7Nn7dnSC2KDpGXfGTC7O
IMG/s68rRjsQglBTJrIPF9y8a7s/6107L6j8DW5KZ2BMhBC0aD8pqFlMEgzm
VE5s5yQ3b7nC8Tf3orSC/DuLhTDrbKr9OqCG4zN0wZlchPMU36m2enmsy/WY
y7/wAYCcLIFVH+G8cpk8y0BiIn0Ww/aNd7VuxsEXBxPyyzBzMfjP2N++K1y+
HFxsqlKJw895f3yjfdtD9kOd3TTFedyikAM5yahQbkyOa8ma6xBKZ3oCTB8t
bkXWgp0kh07FSk1yUqPL0kwL+DX/tSd3/3wNo1dD0DHYchxRNvResbM6E4al
tEkUk/Q3p0Jk2wkVT8U+hgkDUToX/9Ej/Thp24oB/7rM+2qapo0ci3LOQKTB
91BJwbZBWpwXI4Dj4LuwzTIsrqtMcYUX0Z8vbLgBqatC4iHqMRfPwBipte7V
HYfGS7p4ITq6RPYNZPpJbHH22GqEZRD2RCI9VmpUpiGL4Smzk2fgC48pOeQl
AawMFnqg6Eo4P2ILOKaXa6oj7nyZjhiqNj+0jsWKUU5vgK/Oe7kaUjtTlVzm
p/e+nirDiK7FcInJW74Dp/t+uKmtsQwm7El9KK6I91l+H7iJp+uzyq0mACmh
1iBhbKAEjsxyE0lA6tDiDsLjUNy72D0C7OMQLFFyI8QLj8Q06uoaHt8KgnVo
Hmqkhl/nx6Zp767vPpmvfrkZRPNJUPBuQ4Azm8T1D4YCx29hYrknClOI0r7U
7xzVjuQi/ENl3UJaITkqr9RLEeUAMVBVT/hSgbvTrcHA+F5cX6jXCjeGIiUq
v9YnmxqUxRrmqGxCMmG/A3Z7nqySRcga/SHFMTbIqwauNrNOLO5mIj3Hs5b+
sqUJiHfNJt7Ck9tr/RWheggynj54V3FK3wD2Cj/0jc/sIGNsLPRPOYL8cKT2
n3OIbycYxf2X5rl6DU77I1BXmWCUp4SYSGyx0dfAERu3v1XOLFCV/TPaql+b
lihH3733XgFWF86U/cA6aHtyW3w/phBP7B2Ncvj1wwYXANle3Z6YUUY6rfVH
p/CagR4f3XiUsL+BZZQWjy3cBqnvJYS6H5ARkprd2Z2dLthyKLGQsDc+UTJK
MRFmgabovKmmbiQ0E1gMEA3EOv3WlCXYem1+hyLoy7W5K1XdWX7Q3noafFFT
ewhfaqBVYccMjzA8maWBPqiqOFnOE9RoJzIfKmX4D/zn9+n5iUo10vrl8yHi
uxz+Wg6dvB8Mm5FpqwswKXX4jL7XAzNE0YadDN24ACKj2Tm0LxHQqrfRxwal
zrUzq9Bf64gv0byJrsfnGRNPGSMbFS0ILPSeFLGi+2O/wYFSl9B7jqUJ1DcQ
XIiTeXtxUe3qFI/G824lcOqE6ro3JPL0v9mWtkdzxVTHg0BEqpRABqguUV0m
fdgoxwplyDEYvUUkjZ+jqZTSBT0wAi7fiBCBaFBeYc5flqoZYV9eSLincL+P
7kkSrM17Wx/l8NeUD5TMDnKdZA/dvVjy44wFLIrpYBqLFeYD78gq3a48sZQx
0puTgy/KkwUW8b205Zk7RWui9PoqB0p+BCa215U1F4s8G9VG1NuzmEZ75X7W
q4DhWPKKLpAQ4dT1vbLbMGEiJRREaQsYBtC2LJ+ywSTNevMkyvumub88KW4i
+wt7Y1x9eFfD83AjggLn+PVbfEnSMauIJ2izqLxYQphSdJGjjjPpYApt8iKq
v8KRw4WXcieN3LBeCk0TUynGeM658cQMEoivOYtwHV9Vm4XS7+BatEZmjax7
uQXL03PUSBknuO7eS28Ejf9TjhN6YCEsfi7nKcVcHsL0+n/6eR1vOm5BmM+B
IlEbdLWnGN3Xh7XRqK/FyczLvEqaSgeSG0iMg8BEfI9hjGlg2S0GyGFiNI7g
NibF4lCAQK3p7RkHihMk0eFcs1G9MYn7V2XSdsbGbIslo3V8o5nwRLe1CpKb
LbF3AxgCYoD22ONiVNPMCAVblHj4gJtI2kV54bYl+h2u1YTlKjilWO08yjF8
QlQttMtu1ZvVgepkmpK3d1ju6oPvMCRAAdj4WxJjOWxDH2YW9obpYXZe7U8U
0jwWAHHSagmsX5PHNQkcOnN5sEmsy2FAySCkTYzhwVdvurGiaDNxTD+ENCNu
KgMWxG+TzcjWRRr4rGUZGbGR7JS1SFCxtOeFCHOluN+4J1jSOyRhXbhznzsG
OVb3TPZRIpQBS1zJ6l1ehNS/CKpi+03xRR5NjFYzD+L5ttm9B3OorXAM/ZWi
+CVCd8UJDCCjPnyA5iav6s/ETa6pXyKtaorSBsNPjm7hB+bcfoNzH09h8xyF
mgFBxYEWoRtYa6vc2ljLdEX7O06gmHJ2rE51aPuMEjEBHwRxH8DhEEh3f7zF
UhVLlbpDLXrsCIz9S5a5RcoNHCaWC5PodUUB+F4LpCHqWLLBV1IVpPoRgqAH
2xlP9f5Ouh9Fu1QS41LOpwm5pQq0OHDwfd9XDrRKDwLMzmibIBFpoaDveFHB
hZ9VFiubdBQKDpNxFfN+trLmrDpLU41KtdYavyyQTckPj8+CceJLzd7vuOGM
JCKUkAo9T2N0uoTJ1y0JkbARM57NUIKtJQrUr+Rze/pxcx2MtkL9sTFc14F8
MW+mdzrqxKaavAmG2QikYujFHSHcLEsvxnKLqZPhD6TZ9NVXbaqhKf5BnNrs
K5L+rPPUFmVZ/x60pe+Wre6Hw2DuDQoZnOXI5M/GUKjaVpdVoRcuZDeZXunT
Jd2iS94gFv2OUDLJ2BwmXdaOrUCwLn0xoUXWTwnc7J3IJerucvgJnD2u9cBw
URHhSEyjyW/qjW+AqS3IPOllzg2gMtG0o7BT+UoXRRtr+AYJ7R34plR2GE4m
25T6xyoY7UBA/YdMeuxk2xZhxAoDXAah1s973HcKKfcN2N8kBXYqT/jS+pHU
lNZd1NOR20qSS2H+4J9FDdNrd9HJPOVNYr7qBjk4sxr7uf8wVkr7RcihuzMq
lkoHTnd5aXuWNL+CGoasrL/a0OM81FF4MFHACWqH9opKGMCF7qQVCr99gK59
9i1gPprBZ/UTpTBlNJ/X4INCFr5siDOzLchXUI0lnric+sAH8wtZtAHFe4Wy
DjW2dHTHK3X/2wI/IZIWPZxYadxidYpC0r40/QUN4lz6amzTTu3/tGILQ9BA
TY+uSioKZDNMWZC87melWD8GGNLEiZ/5p0ujA9WNdxRVcDokuMEoBMN02BHy
jKb12pxNRWDlSSVYB9vssGJ3OfcXzJir9ed3d7zFEQA7K6COi+2qiivXgUrt
G/VPB3XsMbVgkpgOhxvJJBturFJKZEOi3P+6G+C2rkSrs/y8cms7DLmfdXq9
KO8i/NaF58j/1JpVuSFgYVZRT7SWUnN3Zh9aghy5zk65bfYeKTXXY762Xfco
hyXRypzWk22/Z4Novvq5UOYPTgnQE4OW2HUGhJH+QMCl3aCgf4GJk9MICp3j
c8BxsOPNvyeeReUXV4VslPRYrB1kM8k+K07GhSltQMiwmyABXFHXzye7S/nC
kZpowijVmIG0+mJPN+vkMKj4HvDOlqx3z3PyQHCsWDFDqxzph1jb8yh3nx//
Yd20L9Vhg9Ajpk7fkcie2jLpDQaE6ecpM21ys8TWXCA4PDhtBlLY8SOXWhCa
GPWKXurHEFWXdVpP6wXU75Li1nwi1CyFRzo1TeQWWDxoGp8+eW4peuLcfsww
ZdoQpUQifYKVLthM295Y0Gq37REw2mv5vxHu1O699KFy9jPydY/IiAlCjpM+
sngY9eGljRWMQY7GXvJsEwMyQbnEBIh7kSjygxohyw8cZ6WCYuiVBwccNwpU
WWdJqfSGErEcN13cyVy6JOcpSeQfyKJWxcfURT5iiJP0fSmpqtFUMF8raCPb
XxztjJU6PVJBtZ1N5u3NdFZRJbeSoXdX97CJ1FW6fWLWmPmR8uSBdofBPPUs
xo/uDNSzDWFNtaPgrLkgnNxabBcNP92wDiGkLelxPrHUeSKAifUVGj51K6rA
pVWFGj6vFN3GHPlK3UXS/3MZJZnO7mmZ7ESd4nClMfqhhdUTEyBh5bE90Vgy
1ct4a8jyeiex2DjBzijikmTc2yzjQsUHCynf+SJA8D8MuQKryhhP9YTnK8co
dUDShr6qrSfy4j1QX2FxwpUuG9u4q/fQPNy12sqOFXPdY+9b80C+X9ioMbNh
XYQIiA/0vjpznxRQmo3jDht1CqY5A3AtDjyHEC4lWVTP9rLR57hcJnDAEMpQ
jLgS/p7c+BsWbiQe1xnujAZ3vYAQh9mESq8YShtTc2DX2KcMfCRzIuO8LaCu
/Pbuhxkkm74NaahVHAQBWsWq28V4e7lkRHWdPQHZOpn54PyzRUxfSi7jPvWj
UUtRk0NYR5mK8P4kOJTkTYI7nYzY2YtZQuR7y5pm0GR5Rzp25YXGWwnEIIfg
lYbp8qPlnfU+TJbb5V1vsaVIjbhMXx/ALZubnrwrUmXBY5VN3KQsRxze5Mq6
OcPs22350t/O5pENqq6fzganRcM6W2KKIoTqy8zBpCJQ4wc3xI0Wq+oFdsV4
vTDgdjpdyn50EkaCjVkbAX2ohPzbav1s7iek0or6IjDW5yMjGuayXF+Gtdze
3FCoxqTibott9KAk+DJ6MEOqLGsy+/IgAa8siKD1ojWe6yenjVBmRLhrRHMa
CLgl++PkCQtAjfob9Tl91EcokVUCnPhSBnNpoQjBmNRR7QAMgHcxmI0WEqb5
JNGcvTVqD2Y1m2oP59vmHCAeuYe9waOtuF5kqvppOzrVnBhj9AnfnL+7aNgz
nU6FyfSskvEd0cLBYFQ4lyTmtbF5Ff0OUbgCwtndZ6A/RosJ2rdyRCJELnfK
8swDHk9mPoXf0EqN3jE5DZ+jW3anRCeNwUk7auMSzeKmJ4NokUTVy0yzLYl9
SU4e6ajpaWzStogDdVIJkS4cBUvCNYNvjrU1mzbG+GA2oQJEPop5TLHGhZoE
7kSnIAxsvdyGSlEDvXHHIYbGeHi2NAfdFzFMSxZUeff9bkePuow7HlQ77VX/
zavffgbj/Sy3RzaDburblaDdteLsLF6Z4ddRw0TXCMiAtTLoxkP+Q5MZukDB
5xwOOqxSyFgyry2sOfEIuWDenA1fZIioxseNK1Y12iK4bGOReytPz+D2miYV
I3wf9q9qxXFbM74FNZBgfxIopbUnBHwkvF/pHsL6qcRzvUwS5cp3smiJZgUF
r0Edoazl1E+EblgqpzBdMFLUK3XIsQNLi+AKvLephfbF0Uu1bL4Z1oceWghv
qNruHkZwpSWI286zjckxo4kofSd1baGJxs39jNKuIyCz6nwjmcFM/qDPthsZ
zNPU3CRWlAzVYRMqKTWK1ZmRqoVgqYGXtGm9hyBNWTA1r69erWDl2nfL2e3j
FvCeyrOZnnoSrrOHYZNkF68q0K9sEXtaqcJpZfTGa5H8EM349VK7VC5OtLET
HhYa16yUyBqA0xbtAD92J3MM9xHGcW1pgj3KgufzARVUbMOt/r684ldbuwAG
qIqrcKkRWI3wMMyUnUUD3Cp+DsxmPCLeGwS3Rp/yQQZWBKgIO4qIcEFG8ug/
t+zL1hzdqKnPX9HqTiA7hQ1lCrV34d6TwaIjr9j52pmP37G7hsv0yhJjKbNy
j/SYgS7Eh02DJuo9xobsG4EZ54R2ESDGfFq1i8nJYiWv4b7h8HUMEHOvqJQx
NJaz6UpdrsRSjXkFd3ERmIbzYssq4OFkxTCKSHUYuhEeybWjNvK16FY+wqvk
h3osK6XtZcuF5BIC4090Jcd2XPJR3+4VL49SLVZLr/DFxs9vzj9zYcRcdCiW
ftPLukIbAti9L/ppT7e6LX/qC6MiFAIkeq4zF1gYeIYnWwA6ffFfKPc9ZIy9
wg6UXOcaEbwBw63XLPjfz5Chg7VI3NR3Ki+OOXBWtITRBb7adHgeTG9ABx4X
z6mro7sWrW/RSwEt+beIKe4eCfbamZahsJUqCh+JIn+rCJpH8wt9Imfw7Dww
BZ7+ZWkdZeC8hzf5Z3MzlIjwqeXHkXzFvBGvryMELandZzQOQQdGxfFxIbVg
aULBsf0u4H9rqK8+8fJd5FbH7Tzzcquf9tnvS4+H26JlKIYiE0BwoYlVddnT
cD8nCYa2agyokkBPGsA5hBfvnlxh8Rmnajwbnywmzn9Gf4a+jOpndwvYQZp0
NpmerEHYp6qy0Me5sR7i1ZKvHjDAL7aeprdWh2MiuWcY1kELQgqfhGqj+LSF
t724u0snWTnETr3LbQO8bE2tCWeU+GIHuoumiRXTDSZIeooV5L5hwpPeTTBu
hKPUceePrVNpMSpifb2WUfabuYJpII1+AUkej85xCFsv/oSakr/Tn4ZhLwbs
y18HUhWhFRRJ8u0NCB7ADeMnTZERf4MomdiKEVnirvMQZNt4h/szi8Qakfl9
Yp+YW774hjbu1sMN0GtxJY1LQ/r7DhPpLGa7JMiW95kIn1c31H2uUTLJcxlv
KzJpjbKbzbGFbtZysfHewrMCrvMb5pE6TLUBfAU7iaVBJnGhETBMnUrHlGo5
Ertn2W0QY6BTQgY02q3HWIVbNWWGudN80a8ua67hkBuiY+xpfaY2g4mc5bKG
ppByKY9oejJfljSli6YRIavWaUvcOJmGfjEZ8YrV8YoB48CwBy4Oca2G83jE
hOBzMT2kD3kvOeTfQGRREG3hEnS8Uv0gmFDdF7uNUz6fzapXMYU8M5FOZ3+Q
/oOoD7jZMcfrEbjPZlXjc6Yd5AOJo2X5oW+ZqHgV+0hK0RVm+u1O6q9YX2Fw
s6Lk7jPng4jmGuttdvIFPxnOZX5SJQ1WVJ4YPiaNIcBvHudiRu7mXHpzwPO5
MCN6IQZFGLcqdL4Yh+8JenctLDm+sdnMKkLpIcKCAGFXYGUbBv5utNhsjmEQ
JMeKsRhNRzbiKS0v3q8x/boE8JE4MI0/oFHbC06IqtuLq2H6KFi6J7ljHurM
cFe/xJHY/c63VdP2zr/3IL/NKyMREmOztpW77UZN8rdyKvGxt3sbr68ZAq+m
8UCs/GgiLlGrmgfv+lXRVBzZ7U2poO8h9dz2y42IDEug1l7a523+MjT9zc/X
/LezaJ7ECVfXupHsiU16Cdo8v7ZNvWFUL/VW9+OYrOLQYxN+6Ljloo0ax5Zr
lqFi6TniuIapEQsPoxIgt5YPNYduO1bdZ6Eqx+IKDKfbuwLm7w/vJ1pjSUUN
k+Q1zPbHd4BNFLwBr5KdpjRkECP/GE+RyMsPKkQkpsJHOMzkKEzzUSrfUylw
sX20fEQ5lix7B7SLRbso+NIFo4g49jtAPdOPm1hjap6kfhhMXo007Tm1BDh2
jfD+hLf3m+5L1WaSqF3Kr9U7fGfDmwupGPbrNDIWTWI71IWmL1wKU25+3Esv
/FUxvXNKpDTBvw1WzPW7NJYTByPSwVXEz858fR0VX5+JgifudOys2CGsC1hr
FZgXNqgr3VVyVJDlty8NEjRUeYDRHLRSaR5BbVtlRKC9NVorQFMcmL5e3Zla
5iqu3gGrxYrwPjObjyZhACrDMkbCkl4OeLNns4OBVlx9vUj+5DPxa1UBO72C
hTAN+jbM1kiCDqjimh3nCDW82+viFCT6rftx8CeqH0r8UhdqNK/bkKftQqyt
jP3lO0RnHIRuf2gs4eVQK0kxlWgfenRtBHSpdLTHdROObqpgNqQQo+QxlTOH
c8vr7XHYDEWi7lNlmngN9M1qiNYLTxmbx6PwqkIZ+NE2CWlFKg10iWx2jZDo
vEd2R0P4AdkzShA26FNMs3UneM8jT8+cB8MwsH80Z2vXslqBmKeh0vaUxF64
i+wL+ffPzhsZ/pc9Xf2TTvFVxL0OmSQkG8s+ByN8oaPMwmAkFJLoDKf1MAH7
L4CvtZkzXl82incAcm4PcsjW9PWPf2mFtQchWW7A+QW8+Nwbmz9/nrDoIWfe
u270yH8PseEuAAQUBkhAWVekfU4u/tKBsRGSJVSx1/Cqa1h0lxA7t0TZbYkt
5jJvYElfFo42jvWMOegPAJQ4uQEEJ8KFRA1gScXI8MphMKfy0j/IcyrVE+8h
eSy+WtfIQS2Tiy/gE5Yym+3MFOJzUGRqSbtg2Vf6dgfO0IUvSQObOyuUnR02
gcmDr1usQs0iSfVn50gqnNn9NKIzqEuTMEVutuFYgJRESRoShDFFGvcGw42x
XpCMgBwlHmqK8pEmA30JeCgDuTJVtfHdVk2T9QdAKsCLV1fwMFvcLJ8lbzKu
UoL5JeeQLnRj5SIdPtGbH+T7FtYHHoYzGCGoNYWcc8woWCqE7gZswvqaHoPZ
8edlRwoEYmA/7vS6zqWueuYr5UPhAuY8TmGUypfKxe45x5DP49QeqIj0jgsH
OrDCRwz12JshKle+CB2MPHit05hZuReu5kYE+JVxMXcdTpyk40huNsYvZ7Ia
TsDr6xeo2L/8xR9vp4PfI5Dl67KCxrJFMXTM1nDRkOtExvEtSui4ECbGYeEi
1sQsdNfqRcGO8XA8fVD3TAwsemWX2HTQp78loyciWdZ1iT47zeS6Ig6w4zVc
R5Suv68Ky+hpGYM29Xfn/O0HdzkddinWSuxy/pJoYLGIk/6YoJIctdC5iB1G
Ziwv105fRVFMyobbkDctw931o4JHXiFSmpm5gaJCjb9PZLKiQgtKOmUasavG
AHb7wYs3lem7Rtj23HT9k98GRkycK9PcI5wihA+Zt3ZYSU96yH+jfXa0vgtp
+V/Af1d+tBOEQ0aElJY+aOjiQXbzIjX8iWJXFk73VFvlJdjjqMtLmts4yV9q
iy4FGjr4ak9u6JykxlOnEow3KSvk/FC73kEriojibOvxDLdkPC6L6PQiV4Ha
Rl5BmL/KztArtQ8WiVmPPRav8l100SoXN/MbE+/MR+rf1TCwn9H18zY5ID+4
BQNSdDSvPpawBA13Bh/Rp7XPTwlc1mwZHy6VlS619ECahqU9v2hPHoJHn3gu
CTt4D5MN6M6aRtgUjdFINVoX3CNX05Ygi3gT1YChNHMa/ypsO2iuRqfHO/iD
yZ/5KqEYjwExQLX/awnID7jEMJoeYNPA4P6VNa4OnWy1n1cu8E6ybuhHfvvD
vH5th/xne7NnCAvqcxiEctkNAUyotL2mBK/a2+y1W64zmdYYCigKKbxRmZyG
9S8sHn4oUKuTepRMcTLrQHmn6fTRqkmMJFnkTuATgfBwKo1JkM97AMsF8D/X
SCJOfRxGSZcPoS68yulEDTlM0FMzwl28AX8fuTsYV6DnxcyW1rdRsyAaEbAW
pE/N6dVt0yNx3+xVPFDrWTR3qEmF9i8J/XeXhuWJTr+vNk50e3iPw2RkxWc2
+1rx2KPIQwd/oTZ0+uN08GQOt4NppSLoRuG5R1OzVNoBjN1nK/fU4KRfAV/F
D33bCcSy/0CIAj+qrAZpdNNQDrw8hovbkaK4DifH9PXpOyrbrJwjkxPTf8ah
Pc6LnQ5Pf4I3aFha1NndczKYqil6snHgTmj0xYiRRcngeWOzKGs5l1wjeAaZ
9xf6IvTaj/ZK/tbn10KHVJcvNA/syTFY70o1+JPWyG2PuaLz2G2EWJbRKoop
4QtlZaCEXXK6Uw72wicrhXZiOJhVB2gJ3iM+OTZ6Wvq2iRNI+o83nL/vQ8PS
qR1mC/+LZhn/y+svFPwrKYkR/Dxx84zpjQfccrYRS0PBzhzi9qd8sx60v9SD
dbrcOKQzCPTp+ItSqV36JE8gLqIAVg9hedxOphHNpEq8gGutMqzaaX7qfJgf
9fdcYNr+opEO/ySQyBq2/IMyy3H3H/6sbCraocD/lCqXNeU/Q1iOQNmbOP7O
/BxcJXuA/RnLNCcJmGAEDEunJ9roQyirvUzLCvhuEkMWRScbky3ErhxxZsPx
8+R/KF6So5GP5TdZCWx345b0ZZWJW1ZRr3o5rw9lCdX00tvHrYrBUrpQg3nQ
4S70RHOBx0sksYgVjPXZyU3cezNoOhP7P91jkqDYjOtL20y4X5Zw5plMjZ5M
Tkafsv9BXq75jluDAN/dny8O1Q8uxl44CB5TFU8J04UIKZr5/yZS6mYsFQ4Z
3qYJjqNheMaTRhECQDzyfIYzGVVI1MTQemhtHlf8VIOlr7x77N0kEQs81zd4
LWL+mZpO3Cdl8WXnKi/WmMRE+yJ7iVeCZ9OPuLeMUspF1o4rcw/kk3xB4R+T
L26BExMOmWqPxaTXBpdOLXrODZa2aJSHbw3AQqqYEBuhg2R1oiyCeyDHK8Kh
T0W4kv2Lppnu8digP7Pfza9iN8hxV19sdp5QM/NsJxUocZVkrZiweSWbsdoM
szfNheM9h8wXm+xit60iWmA/u0XvtgZshy9ezOxDfB94jgc3EvUyVbg3PSsi
Y1pnfv+/DW0v/C0O4UOrbai27Z0N/jTndM90Rn77XMSeNl0GLyf6zc9HFGCV
ysWwCUvp7amEvrni05qM5Wzj8f4pxHCJ+C1WskH17NN4aYmRObZM2i3qMW+a
T/EG5vDX8+fXbkl8Q2cSBOvC/FIS/Q3TPk6TuglBYfrNha0tSU9c6el/BqYh
tV38IuxfUz6fLsSpcr2Jw+v+c3CppYfxrccSqAavTAo1gQXchdN5reqTYJeL
ewnpSYfzXtzUEZpgQdn1XGy3nRxEvH8nn1tc/gkiYSsOC2niFuMLiHSawI7h
ub1npRH7ViqxH4OHwbSC77lfp1sdgGcf/+sBMgN6YFJAXB7s0Uy8dutw2SeG
iQSRCKVG9m0kg8/vzCA07BVXRBhf/AnVklJ0GXYTJUruHsVpZ5Bv5KdpI9HM
AagpzpySm3lVzMQN9ra+pd/qqL2XOaUNh+JAMETl1bpJvC+HmbrWYAM/gpVN
mw5cgyrPO+fSYlAGI0Q05Ig/epT4XI+nEbBwQ5Mr7i1rP+NgRRTiPZGzbpR5
oX2fpmkmlYbabzs2FLoQkZp6U7UE3NI/6y34UVeYV6MXtNnkie6VS9WQvSQK
rIF96iyVosiZ0qPb7iM1bMlq1/VHiAnbZmNE4QIOw4+ZGHCmjNkf7AbT0d0Y
MpB0Be+FMOEzYP03YmWBqgF0gz8xYTRnrD+Gp/BrKoXPuSDZHUJjXLpWFiLN
JYjxgkFy0r9bS25hGqC+kil337fCbGfqG0yGDqE6xQnG6APAiXISB6OloQo0
9gcZkV5TpR38Nrf8B1poen9W/VhNWZwj5NdMTcoMPubFkusY5bdEaebKWxXS
vkioAdabuRdg53yMTYRra3l8Qf4zg3ijztbnwOJUQNF276ZDzgHtUtXbIT4k
g9QZ4DzQiq8L61JqQiNq+c2j5H7J0ZTOZTA5JTj7DVOmRaJyPQ3nVKfTa/j+
V/BTM+P1sulymV6NSZt5J53lHuAUdg/4qw5htIvE1TiVrHBAI+TTAmvs7pFj
aaLbWaVoFclyWy9J65BYVFDSwfyz81Oc5OUU8AW5nzkcxfcwFfLd15fWBAm7
fQdOKb625vaALtU+8zq58JRDkrip/++uzKdFwBBzmrsa1Xb3eE/Q8ulnk05/
gzuDGMsuJbhSsKaqQj9NpNP4EFAWKClhShsmbWLiaRkM+LS/hsZWxJ6sq9n6
/coWmJeqo+/lDLExaMHE7Ei8SbxormMBTXuEfiKsDoc/0l/elGqZrRHL/lmi
GDBNz6xaBpse9xidWEG5/67JcivoE3LzlWsu4jXfysZroLctmoojXQdvWbym
tNRg4Nc7OIMUx1M9BQwxTurMLxXzqbQfy5dvLUTCVuAD+fjn9B2vkRtr9zhb
8IeqZWH/oHb4bWWGJEdgNR1KUZCKsAE/DfvWSIt2FITPS6T2A5/U3FgreZLf
iBKqpUQE49tcmcNTUUneZdwJakGCZgJ0Jjk+n2OHTRgUpqJ49gdYBoRGUuYl
qtmxkt1rMLBwsmKjzR7ugru5XJxGNd5O1V0nSz2nKmWGOkAYsf3IiH1q8yLZ
J/lG4zhox3a4Qj2KKtChZtVftV2z/cLj/K8OB0DLvSM5yFegcL7Osyokkc/n
ce5vUwn9g8faVGUPDK653eUOvSukdAgx/nW5mFMLtQE9592GVJUBo4ZlLcyL
TKCXv7IGZSBw6rS4MLAKCTYkbi4b8h0K4Al7bQgkgvjSCF8zhwWsAQ50C42r
9SFXUhKf3PXOjvwnNjsuLorswAbRbWypY/yi5N7+Gqiu+IS9vij9VG2r3Klq
wakLx+wU5WMkS9UoRtYSnDEQJH+y2jaRFmwTv+VP/l2ueRd7Tb6hn5yLY2mf
ZNfTVw8XJFT3OHsh5Lqsyg9Ki/pIe4thVUvvfi2/iImligKADOiVTZYXCm3V
ZNjNLX6snMh6jXwBOH/03ZIXFeINhTGNeZ7zum09aCg+f/XiH3nVBlLcc9xT
Jgbpvs5NYYyKDAzABv0vDy1hdBQIzcPzX0yFqzkhl8bt7HHqRiA5cTwEwge2
wd4r/v9pP714FP5rtGY6xTlCW1IDfdY+OaKUzXkZwfmbGvlUc98/ZgAhyX4K
RUpNvQUuJqmtinL4f7Y3lQ9BE92Il+14wZIGG1eGRnFJcxH6GHyzD5BgJaL1
/vcu9aSIYUiw5T6gryMzin162721Hpap8L/xhMDPpFA5E9NnB0y/4UrZPcI4
ODlN+jzEsr+TiuwOvGXOioPiLlCM8KIkq98YH8Zf1yZpeX3qmPLVKHdnA3z7
MyZf4XIjFTrN6peS1m7HbsWBTtDVVxcI1un2wknoJgB/UQWCUOs8EqnTJH43
PppmGehru2+fkJZUWeLUp3O2C06SnRDwmV3iJWK7E3/uOMwB2yJ+0hKxPdqk
Wfov1Naw5a8uAHqoWJYmUzh7DMkdE5ImhNzQy2uwXbbErhNQO9MYhBq2/elD
vWtXJUpvuCSLYWe4MUFlOrfRj1qGAOe977tDSsLm4dP/MGTjwicMgbjgjB+d
M77dyb/kV55JpgkaAXtgfOL8vaTbmuwknZiQQNakCTMO2zU7nMYUd5/+355D
DFqOQnW+nFVhAMd4gRo4XpsNnSlSL1WLaAkE20uPv2zW2LJO3xVR5IqzXT+R
ncoJ5L9qd7qhfrwdN/EZlBVY6dimv+tIOziyuDqZ3g9kGqHtiSowFN1gO8fu
12s0f8d2tgJk2UdlU6Z3QFrRAV31trTT1ibqDAJOY+juIgRZNEsnRNHeTXHP
Y8Se8lCzeU2M5WmccNJpRmnouIXjuVz5mu7DipVisQYVnYKNeN880W1z/dtz
5ryJ6jzCc/BcOHsnYAKmiUcFxKXAd9elbVDe4VcvSFsnFTpWOIGM7JeqZt93
hopKRUJeC1+S3J5tDtehAbVGO894tmLDDKIqhLBgLHUAlOOFgyOdvte2HndZ
XowD3utwezXN1PRXK0ELWI/pL+jQi0MXNav87kxghBEEYQPiuREc2nQ0K08p
e+gYZ4xOtUxtu8d1I7tHNchegAsIBEDJQeKd1NCdLOcSspyitdLYAZcMkeDl
MetlCnmFevhFupWeJqaBSdYZt2eKkchDWq88Gm8O0nNrGxtKLiRPc/1kfzEG
hJ1/rYlCzgdwPQ9dhBg+dTP3tY70yINeLF+kP7LyluWCdwD3GM2LaTyblFyC
pm9eWR+GZI9F9IJqgirPQDxoS1q8xM/hQrez/bLXNBtY2Iat/2x5f+IkHLio
HkgPv/gSNaf/CKG5cF+GDsq1MagouOX8IumWUTwa9SEm191s1S4rYFtjjEd4
JCCbd5RwRa+pG5NXIaMhdupzUJxnNdyg67ueS+IieUvuOwfj2fGrzT1NxgUc
v2fsh82vdGrHaiKDZOM8AxGefUqDgfu0u6okm/qPAAPqgAjGOo4Rsuy6f4ZR
WiOUpGCHH0DdJKAON1yvpYFwzBvVcBeTZ4tci4VFjrG7ZE82+q6VLy5QNOcY
bekLBhQ79LvL/xTmG+SH+2dOcq9A4xtZ3M62pC1hNHMzL0wWV1wCp5g+8D8V
ZHgnYAz17Dxd3hRirunWhQ5jNkxeWwPi2ck3ZI9PflgT6v/UbwVfvTC5H1Xv
sH6/8O5W092FCnClgtlt0I36mpl5mv2/I836o/k7llpcEynznqnOoqSF6nhS
xwY69VjFwm8FQB1QB0HVmacw45m78rk8RtiZQ02BiPtn/AaE40wypuvHn7dF
aDn2Hx61QreoO7zbOWby8uVe9NOyMB9TuGxL0vGtK07tY1HMdiJRc7WulJyR
DLCJg9SVKp7lVjYqKnI9huprS6t5upsK/cFDOWBQtINpCa7iShCK/VklwDtF
JTP29GGk29V3qR7uUyOIpvovDbbSlOMZBvv/ihAYLI+3DMSkyquJ7b44BPZa
Y/pbujmiwool2WT5EDZIPzhiYOgF3wCBo2CJNYohdqERh7vTSnliR5XCKF+o
/TPGOW6errw4xvQPV99M+bod8Q8UbeaVB2D2Xyp2+Z800pr1mxyz0bCkwMY7
3gXUbgtMv4qsrvVI2v9sDmjhV0I5TdMoU1l7TW5VYOt5VjC4Of5dslM1fLK2
kaMB+JozQ+2Lu+wnkJnYZ4vMyumiX/ogDJPbqvihh6ip/wZtRIbbdCF0EDmJ
rINbdxzfJyCW7VR7GU81x3gnWvwe1y6ikEG2sIPrmttlLw7DDWiiQsBMDRgA
zOSaLNxIMxpcVokvOUb7v0apmzUjPx9W2pIGxcmyi+rsGF5kdefHMwv5Q3Nq
JvPmAKm426Uy1p0aYsg6ma5Gms+5mJQpN9xI4Dac9ZGn8bOOjnRvDVxN6fK1
KEWV1Kw/41DJ/I6nJq2QN7FaCfAXDQ0JHa7AgtufSWdnW0qCkHasrJ39nriG
cALxpF5mtEYksDryUmd/Q3lbfPajxYRA1T6ooCcp7u38qszC+NmK/Or47Gyk
tt8kMLHG5yX9iby8SdR7fV6gYIBPu4AG9ASgqValqrZI2GM63Km/YveKAtza
sCjfKurg2wYNR+iAE5YbiEpw7ls1GWMtGQOwvK9mCOReyc60iB7kAWbmw+YD
PABIjZdjAqRCEd15nAr8LEjFNkX5s0bUTcAXibVST350GiL4y1tgXT1D5IoU
0EymAJhJXO8A5+m8tYq1N/r3y8m2y5eS5O2RHVySeJS9s4hCimqpIZSa2W+E
qxjj17VUcgVRcM+2e9lbT+GJeleL9bpiNZjH/kqK3bi/mKWcnxTm/9UIqLyq
O+rQfr0e0CNuvvY24mKiw87iQak/AnYhmdNg6u4vsu+cLnvoma9ANtFQkzwS
Hi+CdOH9dR0tXZp+yyQQsN7KLcpO4lSDsi0K6fRv4bQGOuspyMAaOdpIjD0Q
v6l8jveKWttk0c8iuq1dy+0E6sRCzKl65c5/L+KOlh111R5m5XzwLaeyVw7D
RLcyE9P6ThrAfMkyLXm4TQoYEvNuyoT3m99wFggdKwCLOwyvBAw1pEOIsE0B
cWzUNC/WMjq7t7/Jz4zv0jCEYE6LpFMq40hpYAEO4v+Y6f41Bx1pAc9LKpT+
lwfNcB3bd58eT1mePs4erMSDc1Ll/KLGq/UCleRyw5oWh3VDImJHPuTb4CYb
m0+MS5r1w0N8aRV9linzTneDdxeT0dNcFtGKnQDioHRud7dcHhZgdQUfYAw8
6gc+jrL5r4LVzB0MO9pSxb3vKDrrtiiyNADbTw1Um9ywax3sZRsN6VvVVg3u
hzjQPp48nNXNUfMVjdSTBUKrfIy2xmsANC+8hqGihAboyis9w3tkYTji4+ne
Wghh68sXJ3KlFK7Gp8h23Cix7mFjsN5a5qSEV0708oTc3tfqy531Wt31nYeV
UP1LT3tnUHJTre6q1xzwyhea93kw7UkTvzauNb8OniE61YIceqJfaFG3fG05
zGlNI1jRExlxCM1TBKlIINl9biIIJ41W9iHVwyX/rGzfHCfQN3nV2VAlPZfl
PZ4EeaJGAxUP4OAX4SziYPbG3lwpUzT1n8eneH4ncA6EeoKlnvmszjK/QVYn
AARJ35gqmOxIRKy5A1oFynBovlrzETYHsX/aQ37pQ5ljvhLj/yaRnFOaI3Af
C09fRmu3LyT+Y0CxyOUrHkR+SXnAyLgt65ZnMRrWQRA+DRgCA58uMVpFT6nu
Mhavx+K4cdyX1EHCTflgM3+gNJ8iq1Cg4RKc/0j64U/PDND96B0rlGusvGkO
4TnW7mLlK2TZ0LpZHIFN+80uhMCyJRfpTVTuC0+9/NrJTf5Gu3XtZkcgTP8/
m4lcbIkKZZMC/MWjvhh3eMc1dQduNWHOaVQN7yKMrpxi/LXE8VOdTiurGmIk
tJ1XlrhWie8w4eZiHWdnp2z8roV1O8szdfZJa8qqDSnUFH9qiNmjcKeOpAP4
8P4aehElwomVYwPsVbMWhMYiw4CakqA2xR1JxvMLbBdjIQzeL501v9FLtysL
VcqBIEEQPPXHEu1Vg3Y3MPQ3SYL1PD9Hi/LTt3FXJ/ieeQCXy/X3GIDc2gIu
beP7EVHkce26+6qlwUx5yrc7uGJXBE1aIWKhe7yfCJ2TUhaKyUhzWn4nZlfJ
L9PPZ389vrPe5PmZPMMxwHKBwQ+75+PwPeIKx7YWb0mjnrsbTukhvBtGEzYP
jUrcbOsb8xhs0Dt1V63+CTUDx1xziOSxtfYKQOZAriVGhpAG0MihcB8oOmfu
hCYw84tjfkVgSiH52k9gQu8HfmVhRwvVtWxTG8OU6akG5D5lnc/hTI/w8gmb
/0mQ8+Q1pUMZmkWkPjSwH8Uac8F5uVBN9wFUVBcsM6kzGxaYynqLeQFmuu5X
IGTlBa5G4UG5q9+Uwy51fiVhFZUdI/65zeDtHUyBD9MZ8ZlBpD8vOuwjnfmy
hZOF9kdCIRFOZeryZ2AzOr46ZuxFjcVckXal7qWtcLxGFhpZJIClU4+v8olq
I7QLt4Li98dzTLVfgRuL/5qWq48JQRXHGL8q3x6lB5lcvTAkIcoVPqWEvDib
+wAqmVFJEYEWk/zqT5lJaqfLxtLsVSfqT/do83j7dDjn+rwI9yP0J3Ig8nsf
m81IWft6uCt0FveyQ5y5Cn85LwyU9u2hymMx1ODfs1qobhn7E5HnNWE5eHim
mHs9qRJ5a8a5kgldX1Z0jukxluB1QQMeeBE8o0wNG1ghWyrrSgLRQDQu9CXl
0lAf8aZ1nE1nJmEtCkmaEm7Be66eJ/l010NEKE9DUBTIqlJOLtmkN+Srm0Xs
nRthNABemhuckHPrFlCywjh9dzgpScj32h0C6+Fyk8u8jFBVo114MaL0xlPV
PjtC2po+5lOd09NMAhDcDmM6zOJfcrXthpnyfxDJQBiI9eLy72qGjatD2vnQ
n0Rzp+szX4+OkSvZw4SFgpon6qBag56bP0vmzx1A31nOm9LzzlMDoDejb13j
WxbScvedHXy5eATa5SAzVryr8TxWVVlZJc43EAq1CAFQJzph9LcvrzbshOEB
6c7/1+//7iGH0dUHx+TXZbGefG5C5+FHqO4OUfPfFpeM2yH3SRN1g0XXsnXY
8thc0LGhfdnCHFC5PpZoUEBqQ+VDxVAFDOUGdZ5A5rF+Wvl8ZKL2RBoTUL4p
n1aeq1mpBEsyaNTq87dfmY4giSNwNC2ejm+3EzZ9VEVXz/oieVzV6Leg1uE0
cUJ36Y6FYdwsogUI3riz1aHFTWcZis/ssACE6o+XFmh4KP8cGlOPhrznIQs2
BR2/Xm44A32X4iVDWSfK10WjpGD4XnO9V5RMplZf3J40uVIwQBys+TgYUwyV
KB5Y+tOHxS4qFGELi4kk13Sp+EHv2fq7352flYOSllhTyo79KnpkNnVFalJn
+bnI0x8y8v3dAV+qJLADVSp6SZfw3UbOrw5BoHt7gmW9yfcC/bHRA+0NCuCo
X3u5ypDMEglJ/S36Yj/NNzl1NaumNce0Qyi5MwU7mKiBxG7/KNcAEqJ+DU06
4nfqm1I7Hgx5HDHJbfvil7hQA7T70N0PUq1ChzpS0Prv28WZy0f2GCghFbfU
M9WmO0zR1b87ZKvW9RpCH163mU9m0w9xJjeNo1Ri903Cu2rrWJjicmi4hd8u
ubQvwsJGcCS655EviHqlDjDA6FqT9pDcAa3Er8y0u0w0JncvR2r6Sd1s+9wc
hgYlqB/EJam1w6vS/6z1TFQUvljxN2P47cZrP/V0MDamWf1L1YnunuOCLtnY
g3CHdB2IjKGmhBsDfkql0FqR0hsCgNh72rmp9nfZliF5z1z7AvMHZmULo7EY
YNdKpkykEu2siB3pHjtO5JINmBmggeUEsB/MyV4KCzjeb8OlZrvVi+VtO3UD
UMeeFZMvSMsiotAuNnvIohkSPYWjoePQHPKCEH6tx7mQo52O6guvLXXRJlKj
mbuVaxSqsa3DC5k+fneeZbJTpcdAm8eUsy7aGoNTVN10nRMv9QuhDce1yg/Q
eMQw/YmRUjmmFh3ESIlb4OpN7UzxpA+BNigA48YJVPRoyx8NcphtzQ2xg4WD
20FMdiCJwXcMJPAQiMJodf+aK8AHk00zlbxSdGkAo6bAiHd56WyHdX8Hsr8v
p1mdIVt8mWJXUmYHCnK9a2mqgNc9eYsIo3fgOnx3OCNVElTVdvFatMR12kmd
bvL31Xy/9TZZjvFbx/Ia5Q8na23UkI7VUAFM5yhxXnIXTTWT9ozwzEaTZVMX
bQlbjGf9joP+rUJ0iIbnkG/qGF1woIXMBn4C3TCdf+0lr1fBc8NrH0cT7FOY
5pezaWe7YFROGQHxWOiD0mjR6EGQ+6FpWQnFCrlKZoHoa9iJxyzn8rvPbbPv
PgnmMQX9C6PKRJOlEOftcEMrBvZTjsdsrl5wO6bu2XrCRBi0dOAzASHD6wNi
ZBFR0tMFo9+rEHx+tuqzkV/+KvvTUvp/g8QEz9TtDuiEHdmA/Pb468BkUBiy
HmOURt7pqYVKlXYJ8xZkCzn9SRn2E2CgBeqC4xTD51EKrVz22aKnsghzF2u1
lOxpK+FL3oduuYZjDSQc8fN8wCSV+T/UmB5PBh3K3GAi1T6ub1wxCIWVWXA+
6JTHwogIpbEErh+XX/M2q908Vd8c9KNSs98vRIVdm6C2mKhF3uyVAPf1HKtw
g8Up3kona7ZzUD6y0hBjKRnv4JCH28XXr/O2AFi2CxGpFLud3pjgGS+iOD2W
DAJtst4YrLPlkHh2cP/pYHgEPtEC/yfZddNKFt9czyZzIy1PVdJfZph51QKC
PVsghui83uQ1ppMQaOdXcb++lmhZXEYUK0VfJ7ErZNLE2fWLoOfZefG4HINO
sIpm9gdwI+lJoaBGDDRX1N0nSHDjFUl+ETPtWn9HdVGB2xyLG63Dui2d+Kpl
gEbI8OFx6uaFMn/H2gptBCNVVEOYcmSA5PHNlgcAD2KVmJLjWNawhrBe4Kjz
NHu58egLIXIWH8b4oyTxKNCbSyMK3IV85o0nWrivH4PXK2bRbnlfn5es7oVI
TwjS1NbEdbqPUAYHTsA1/0bAd4pqVgOlQKCwkU3kK1YAIjHBQOeHvzZW2iOt
7/jypfIdARVlHKpynJP/av4a/8l1rKufM/bc3Qzl90cP0TNNVFRS7eMDhn09
iRu+WsfGf/XeKzug2BTaQo4RWGGevmeNUvDxVgSDtnKlAzj8c2y6Q6h5wJvr
oacIwb1RvRfXT4Ij4P5o75XTzT6dkM8Wwb8fgS1U65HKeYLU6jJ3Qky/CSaz
NxHMgnGI47zGlACnHClo67mX1n2WRJQ/3OYNkTn1nTJUwC6iOrnjqhld/HOH
QDiY4aJixE6J1QRLXtCpikbbWT6mc0CVh5SmsAo+gXTl6nq7AltU+96pXk61
Aku5QHWuVd+kouI1ZsdTvh03Dc2RvPXz8CrT4nOxg8j/aaSOJie8fnicjVZo
dE/7Z2fIfeV/IZXMYXeW0fx6chvMyw/hm46YiHpxFs3jJf9LZIGnqPv+Epd1
JlhAiBituJnoT+DSHK0WIB/rET890vuYguU/DtHqLTgi7/qjjT05jgzniHGQ
/ehbVQJIMpenxckrrbyVhnhqz72kxeCMHehXCDaaPqicDmUil8nvDApfH7ho
mF0sYp2GedqIAi3fkk8G4xgw/dhWrpanhE+EZkAqHrRBKF/4q9m4Y9+tBf3P
VanIavlZz1QevyhiOuKQ9DGwpwrMSC6C7SefrtQ9L/o0IEEIIUhw1SuAd8w7
JP2zgIektmgNF5M37Foe1WB3x+NVeBRyCvSfQPiRQtPfR/gKDyKRizMxuKOE
q1/ND/ovAS1scG+6ruhJCIoOLj5fSPkZ52RvL9BLgPTN1I4t/eVXimOYXmfS
JgxOPy7ct7VKcf26qyBF6DcsMjYp0TxBbYHio9wg5q9XBAnJ3eAzyDxgvNjG
c1wPX9xOglr+lXaHB+u2EMhpO8udR2TpXXgK+6RQC3qHunVQqZTfkR7URJzS
B+Cu5nyluXeGxVfhx9CTfauV5yoRWmyxIJCi69Rlx8j96x7P1d/XxDsTkhYV
M3I6xloyeJEZvOXCKT50KDZbFvap5LSHk96qyq0UhMwNaOODN1zyUX4InZfS
h8aIhS/kdzvZdTizvz3ldGv5jvpEed0Nsg5eSZgSp04ghoAL+ySqV/qygZYg
7yblo7JP+1jqg2Csw+85jMXv/dr0WS9VKIMdTiLUFPrCfH5qJ7jOlCb0zX/e
NMQGjZJcIhlUv59ww4lXSO10YzHshGkMDrFAQIqRYmbZbFcnG3oDAMto+2/o
obA/ypHj5PBFfuV+QSZhnmO5Di+bDitDAkh686sZ4gVBQOLOQKW5Twl3vEWa
yCCcsgXnYqqOVq4Pyk8bpjwQdaSWA1unW/DhvwI5gv8+X0M9hZQlkFyH6Og4
MHV7JPVsIhYcGZ6g4ZhMYo5X1mnkkXtIqNax5wu8Tacltu+Y7WcYV2MBuVxv
tmD524IyNqDs+H5+Z6L64Wepo0H6quvXfyfDj3ZJJiNtA2+Bbj11mddz98Ny
QM1sSjo/cnST+0QiLIfmVAPmGS419ksAkh1ItwqszD4QxaxxJxyRgG9lfZSY
vqYHKO0jP5ZsylOI+sWT64aforQNz9XG2N8g/Maj2jdBNRrCnJ3YyTSqpaOi
/k1w2Q71/NOoNJJLKbrSntwZ7+s+pmYjgaMIIS/l+XQ/EIfWkghrwtA+9Z7g
gP5iuN0G7OcwLTdM4f9RTYfLdqLhXGPR8nCN1tie8w4Fhau+hg66Oat19Azf
1scYuk8C1KuJLH56tkxRDn7TsnsGP00GKy7XnXIvi2Qt0rYfz/YdQItohPpe
mcaMQWtHKV19Veh+qwFwePRng7ZRk7I6azwVm0NkgJjDZMwNxg6tDL9dOtNm
9sDLjVPj6626sKJajs1myYEikixJbMUUUbSPTtwSAUE9UkQZ8Pz+3VP1LCYh
mwbUiRgcQ+mdxUXnM+6ADEUs0V8iobkYLORSzwa/7myHB9TpDiC3qlfKuGMA
VnwRKcRAFyJJV6sH2qvWfvGoOsRFK9aVEi0fb7o/3Ky0ACCN9NMFU6Y/aWlK
cFzR0ch8u1lqc+nm0gTusMf6n0DuevFYAMYFMXFwPmxkKPTO1rREiTRteewX
x7EQMKVylUS9oztIeO4ZEtcWTYlJfgvXygpjnz2u6nfQ4LZ2Ywym5wu/L9sc
TZVgnGg9/YLg9ZdosuUIMPHE2HBynLELHn7V24PxYGQfRR7SMj6NyrEeIHzc
bR2PBXo91nCYDN+I7gff741Gc1129S28iCccDN0whV/wj9bxn9F7mDPFUN3n
IxCgESaOLVkPFpMDB8pJDILzKgB/d/F3dU6o5RWd/IhVsPFzRQo0qpnD3Qgn
3tLoUT6qXjc4S4o18W4Fg08IkXw/04nGjjxtZsdO+Dz99VpHyfJIxX9wZJgV
7rgnQ1vLmxfAtSEGshTNOa5KIzLlNenjwzd7EtoPZN98UKw28qYVrm2E0+mZ
nnXRNIqEWO09aOMOcA3cpCia6sCIwTuTRoIle+0acYpIrSYM3otxCL4KkC4S
3amGnO/5Ern/DGPfv+zHRJS1XAeTxuAwVWGQ6FaJAJ3QgfjpOsOeCsltmjGd
ehvZYx60mat+/5/3lJInDdK7g5T0wvuny78wQd/6qJPJRVVp2iPUtFDG8Gcp
Ts1sbDx8cH4UaF5X3E6e1viaLMwBn6TZmu4l6+n5G/83LZXDM73W8gL6M1nW
D05U86j0e8BWomcJtXV5JtQFkzmpPuEIGI4NuS+H9Eo59bAvdeKKyJe2BuiN
yqmOqhSL2GiHcni3gZJ3sZ5ZReRm/eU5EIBRO6Y58Brx1yHqbERU4SCZOw7m
8GemtAX170/wRD3dulClv4Cs5V5di1hNRCq8inBouDgNWOiO/Uea7ZLj70zY
atlt5ylxqzkjw+1nIFkxBkKcI/aaL6upkREVM+Mz66HmCAi416dq2acJYwmv
a5GvthoKz9kvgat/1QLdaLZQtmDPVL+zwts0XmNqvAOR5SDZgQpq/4ZQ+gad
GEmQDENPgQUFmmCpyxkHxbERv9yY+47o84S4IE9K897jc/IZlQLivJBwkzFy
R/dXkwDYU5DVIv6HN/rNe/mH8HugweAuSQmL9xX8JBagbMCliVtBPFQfnIAB
pI6/bnFeNw6Q+ksHRVGyWiBquFiqZq3+ypeA1fhaN11a1gMGTdcz40YJd9KH
v5WiJRFZR+tFHk/+sWhEvcRwXlDVC7s0yzY9IrK95FMQ64WJZWZUAksfgoSE
neckwUmeyUWRNtFnZn3p4MUGCy0raurgi9R+rsMvBlpCvhd/x4oHNPFfDgax
CrVpMu6lBrKI6GniH2Adlrw3W/uucHsG7rGNtZXAFCYkC4dv7WDLJINYtBfS
iNlJPU8AiGA2MqkIrH/ov5SoePWn3Vrwn6nQuzjojMzuoIoP5iLOIKBh5VcW
0hxrKXTeDJolohaRcNaiObRBTwQEpjvnRXErrhYeYzNGjg+IlckPguxp/2Q5
HOG3qLoNrvqDZr+zFOaEoTiv3lxCzci6dSugawmPMgA9ZezIUHFRMqM4nBgU
TVSxMB563spARl92gqM9lFTgUiEPxzKjADo5r7KBExKbd93XB9bIS2IelQHY
K6Sfz76b5WnC2v3xZkuXrzSfOofxFn/bzZw+HK/4MrgGE2oExf+dHQBnWee4
k/v++39dsyJYrcfn84SuUofkZojwPUqkdpfgMxnHlQgVqjgKPfTJkp1g+xM7
Vjn58isEEr68Aae1ymJvy2n334m3F58SGrMsMQM5x6pLJIaeCT31BqbByken
BNl3sBJq8QMfL3ODBElopampcyxHO67A3cbdKZgoQVpeGSeLTaZM7xpVBj5b
OL/gUiJFYiD43NAy2luSMgQwExgdzYF1/q7FAQpS1c5kKwNQvOFgyARzGJZS
KBuvkTkMaS1V4zSHuZiVDBmUcrZXDWuI1+qip9n43v/gu1zw4JROKoPJDMYc
Ac2KFKETsPjl04M4KT3fJIW4Xqo2bLwY5PZim/Dl5hRT4GOx/g+uvxwvwjtn
ut/40KI3LpAwubAv8K/MH2PJv6ygJmumtTGbCovxn3C6sg/w/TX4RARJ+13e
7RE+6pBGA9icHnNxeImOBnZaPmONGIftaQFVxxxDE/3hNGAt4VKFv/uyPyAF
fmgajUCad75Ga1zW6wXIVXrWYs8aQTr68Cu5s2UD1VYuXcx3+tUGY3GFnWlp
NYOdMzR/dBU3lK89F8VbiyKq5WV0rcu27DOso6lFEMqzW172JVGThNXmyCDY
l/A5Us6VvJ+Nu2dyCYDRdSdmZ1Ije9ggo4QsrDKL23vJFwlQ2SinC65GXYzs
SO3g8v2l/fxFehS/q8TB0iJICGlYoDuTZvAkIFbwHRsohGJXzMFwY2JS03tm
cO5hwKpWDBs871xaMmOmPzzun9zVUPYWnJmunkZfUWLl3ZW/ShJwMbPnQ3bC
aHtImc5QACaqyUh+pcAGN8RYIQjk5m5v9fJP5MAI9/D/bqz57XLf3tw5QtVQ
Jql/hpuVHwYgB8Cj/68emM7vrsOZrqxLRbMx/vTD1ebRY9IZIV8tQtFKueID
Fxicsr4IhLBS6ZZJ7Ax58QRabgi2BVol2mxC3B6rrm04wwoVnA4+8WOnY0DR
34YYigyi6pDk/whaZ/exrqnraBgC2ZOVvix67P7OR4kjVYLQGpgMy5vt7fl1
PRm6QLPmjKSnkXDilHIPcOnDufQ0yZmqY03LYwPvBFLBmIxdD4eRRI64raCM
CA8yNZfyMzPp4y7HkoQZUDr1EGICKzQ+IEOpupjcAbqICtgM1SXwMV+IvXap
a7XItDsylMYAD4T2Oh3x2cursNO+L3otYWhoxXHUtQ8nbpyFyHvJhH2jRQTx
DbXOBUjNUiCXBOTrWbBR4Dm5txFCZ5LkBW//k0mkfoXckqT7PPuOgtjeq4hz
KQbAp78TcHT4cC0oWLQYIPLInB5KLa8fKhfshkH83/HJ9SEmA06nnSX90tZh
eBfBhl2RCNoRnrwApsXDyEHz5dQwYtNJI9VgZyIbxyQEG/VLED+0UAR1ubCv
KCzsmcDRVihPPVTOrXbLZD7QStSX4Ia0osnQV4gBRrKAUw4AdODhy9lmePR9
+aLiv9ijw66Qizxz1MC7VqFQiQepm5GKhlPvjtmbE1XMtoclHbdxgCcRIbJ8
c76QP0bXi/U3v59v7nKgrvlUDj9WNQekCmlx5EhxuT3NbNivJ6Drjpwvss+c
BnowOqWVDEStQfAHnIsoSqe2+AFTE4M5L0a4nEQcYkc6Bl0M88uK+RyKGAQD
c5U3KsDrd0WdYYKjOaLGW3QaY8wqOr3wuLDnpArpc+92A17seQX9G4a5H0iC
hve8FNXBjlmCzl3K1XhomcuTCmaDO8vP7M7rAiUxmTdDBtL1m3aO2HAyU/M0
ZsrtXumG+mrU/s8x3tP9GL/JbNDiZnzVtbk1Bx6mE979LHTCz8fPDsr4Rk8W
bTQblT+VoPf+ZyfurQRummvLNCpMMWzHbfA3wWgw9sIl3Ts0UjK68fKX2t/r
hP+s4BDN6v6VuRllYh0ytA+a50BAP2QOZzFTvsbnZkftqd10GvKaFSX1pQD+
vNFss7ELh1+mSJc309847WwRDtVjaDx1W+0RQA4jPYt3Bv1BRh5Q8W33vt1z
ZrMW1r18Ty8Ail9NYynWUHuJL7hFPBDYZkFZj7Dc/heGiErE97bqTdR86l1h
BhNeQUdDYf2g1hQWlGQ1+dSN4B6m7+LlKNRjyD/WjHhExkKS1JCw78XUeLrP
ncYGj5bX5PVItqvwg6F6oaNDq3u+YfAHTKB2hcYSfbAdX6ynu3qMaJ822jbz
SjmIC0l0Bo4KHDHnwE+UMo+26SguSTQK9oqzhxxN+AbzHxCYclbBL3O8DO9p
16EIj3mxF2vO9mhV14P0RCpxxl467ej01NtsfWKrdQwr8wcF3bw15m10pba3
9i7aKFwpF8K7gq8Y/zbHJnKtKrUArgaZ3OLrn7H2HaIm2RSGeuL0Qe4PKnP0
qR2ECZ5fqspIdDDv+P7aMi2Vjl06z9FtXBARoiPu0ph0z8itQ0jNQh1rxGht
V3MWCDs0HRkAtrPHwfU/TRLi3EV26Rp74BCbnwYWuzJ8viKU1Xu4H2pvKIFW
QAbdB4Lwa83Bom/C4Qlt0FKK6mlZUbHZ3QR/WXR0eFfQRNYb/2rctK+X91EN
/OvRSeSfYn81Pq5+S7S6WKpIppRP354P9DvrM/cp+c9yfnORru1T1tBl8qtY
kdjnUBzvl78oycdteCI1gAuMlS/1igBtFcUEUjcWcn4uams1basaGL6YgMg4
8oRFHin7w+HOFob1HlpcuvGjkmDpoElCVWF0QeXBZ2Lm6WbyoxUvKgs1EcuK
265AK/yn+rVVlXgwB0Yr3LFjXku9RirU8h1cieUPEZIi0Gf2JZgD1HuCUvwr
QNrtMqUGxJmJJwWtoRFgkOCV8o9lPIQBrFBbTArSSkoSo7Ii6SYSMnTOVeLl
iXGxO5BIBDtVNZsq+JrrJGEy2ii9N98O3PIRhqB6mKrjSOKxRYQOxuJ7iDgL
IIvRK4eTvsC3IaAN+ytBq7VoT70xitRjorN4FnN/pitBnJ/FrwMQ/QGv1qBL
rzGJ7HwzWo0D5brPKJq5fLmDuzFD2pnCoZOCFFr2yQgX6ZPKZqvftkrXSewv
IUcBh+JQ9dDB9bbW1EW5+BAb5Jig+oJYbCka3ae3ShHXP3N+x141gwv8YJ5V
p45heyASLnhnAjgE27UlJoTrxw4WSk0t9fM5J2Csb0ssOTIAnWj1lLcta3Ti
bE3did+xFKG2LLjPQXMwwi1JwkiS5g8dIR/BjM8Lhkeof9bUChQ75iGz3umA
ALMFIfbWjtWFLSGf77EyVrx4qW7mZODfw6GSGTRoOd4aWc+trVjJt8JMO5OJ
B9KvwdYJdO3r2BjFAGuQWueNekBuUKTPED7h1HQKSsRV9K/rrIFWmJZ3GDCZ
JcFYwKQMcDtrJ5ELNfgFGYeRWDJRDiBv2+eNXosH3AjdNs7T9P+O9KdTR7KM
Bz7C4ljlveM3fvMK5F3kI4M0gUs0jjjHWs/Oa3vLGs5irrDkOiku3yksxirC
O4JldEyLkLSKJUNdt9QVas9WkzpKtX+HDrlp8ra2KPYmi0jeOQeCPTjKT2qU
l8H6W09C8/Dz8CU9RvOgpj9Zcg24cO2xHh/138opcVyjeqLw2wTDh6G/h8dy
yTYL1CCHtjeFBSu1bJrvkoFM1wfmuK6vv+WA/0LXiogJbTM471EajOJkKdSL
T7pn4x14/BCl7MTeuUIJtEdtJWW+5jpHZyKZPVJRi5CGvQ+Zg1Sbozmgtfeo
lxs49sa9zyCH18ujUs64AZbcoGhlhWZOqk5WAHSMqNIN2BlSV7xfQE1qxS3U
TbmcqjBJOfib4YcTjkCaFMwjGILfP2csE9N63b4MakxxQk3yE9FseFz5aK++
g9qS5RBlYkOL1WemntwFjdlSPmW4mBDwdngErUXnL3xWjjpXu7qJubQn4rT/
Xc+umDOlJYiHFcOiv57r+WooWNcM352ybNE7Hf9UmOQhGHBZpWqmCC8SnpvT
C6ZZ8193wrQGOq4IRQEIa5a296mdakZhxrRiYQYeSYLUx5hMFollXdXmG50o
UvGDSQ5EbcoyaVsC/H2atHU5CheBsLfTFqn103vjzSyN6oIf7V90uaDsuFIP
9kMzhhVp0Y5onkN/h75PY3NG19VWfdofVlrrQprLwFpyCgMww4SHFAnRXv/F
uPACElLsDZ9WbtgezmWaXGc1S/ou5jrJb4jtx2FrhGTUNuksEs/H3hspFQhw
g3mH5dWKCd2hiQVfbDG0SqbxELjLeRGvSI6Iep46E/OXsEjtVJ1ccnaDPhdl
Z6yIFTaybcEzVy93JXkG8abOQG/jVcn0XkGRLAKBraBgSesI8OoeUpmdjlv1
/wOsLkFLr/OuQsMjfH7VEIRsuzGUPgkiPoq+AYi+7oLRREqllisK4XdiIuvj
yjHqJbUJr8dR719k46wUyOPmv6jCD2Dp6UFlF4Q0jT0Lz4XiNlMiZSLYy/G9
Yc9zz1LqpKjcQGiV6AtGoH8f0TaZqO6GJIrcUsPZvSh1SK9LBvQ3AAK27jBo
aniRV6JRriJdanFSEqij61fEIxkZ6/UjkIUc5O0fsoSDQzd6R3AUdCeRIFw9
anhNgorWo/mHxRybsbB7xK+4NwgyeG/a0cHhgu/kuaqZ7PsAugLhPKeXBY3z
VH5qnx9J3k12RgmIYr0ySiFnZjfPP8qDXYO+kCeccFZqHuRFKZPi0k1CzjuT
8VmXqy8R0T26GxPMr3lkX14Sx1kIFAIdOdqg4iCf5kqO84pePKeNglW5eO6e
nxd8KhWnRzBlh00hHxzgx6xNfWBUNnJffZyqnyr3hXBaMYKqZV2UOX4Qsdx3
csRDCFN3ubIaVvRz9d/N8SPw8kxcd5j7fRwSBGTR85wYo7TCZG5m69vGfafl
zlpreQxzVk+ZvZficfTVSGR4htbXjGRBCt2gybm4JQPKH2gPQrS8iTZtfZ4j
TMly380neYAqajjQTsz0aOzArCPgY1t/zWNa1dEKHK5lcsQ/R8LKY+XDX/43
YzcnUiPobOvvrgMS8Wiu6wlQNvtz5+0xOyXTzrwmqNTYH0YzTKlPT2ozYyr8
Tk57mnDN8VbclYVS1yWJMHCCBcdY6AsuNlgKRFzWf6YYlEhChAYwE4xzUxyD
kSzn+a43LODkzvXOikjsHnzTVYgumTWMHmtS988O5NcAXK8CykkvN6eMqNJh
ggjthzDZeFAKHV0zZa5FWTZznVYaiIPVdPCPdyLttcN4fo5MUMBCeI4LFBZB
z0chXy1UY1Im1roqml2QJzcbwfpckwsBfWGz5i3G6yUfFiF8yNDxHWBedBtQ
KxOThzL2giWGhnT4Wo0HxGJ4GPxR7p/GcWbh0JLTN1fMnZIW3K5fSIKcTAOq
EKLN3WxIIs/bx+ykJdoAIeme9r1Qc45WhQhvTSPDaDSb3k3VZ+HYi/C29C7V
Zh9dLfo7CG7FMwrhDgLtL524LQdOHeprdkQ0h7Q4AoDElGCZtt/gTglm9SI3
WH/aJlG4fKolRIAT9QzxyrusfKnpjGHKD6dGRWATfPb//gSgUG9lQX3Vpp9x
+Ys9eWST6f3B4aUNlcttGtVuE0s1p2+k7oVVk5FUBCYylOHgDYMKNk7sgFIh
5wzIQewbTYwFCUVE1HETBaVwkk1FZjhKexOqSKGT1dwKqeGinL8eHWKua6NX
xRV9VaEOq8pYSN+AXrSwUTfqHtinHLxmhRyhir/IbwyiJvnQ7tsKZ8f3K+Hx
q10oODMEUv81KWCcztcr4I4IW17mylNeuwj8MdqPeNZrpL/+8lZXjgIIzxRF
RpCWQ5/BMcvcPpCzvrfP22u6Tsg4jgdK1No/LL77HkQ1Hw7nHRgCazPKJ6Jg
GvHIaUy7ewoxkXe7tpaP5npJNQrggBCTM21tCKhSIfT2NWKZ3Rwd2LRPGAdR
ss/zqhz414Tg5dbDTzCk0ldILz3kCu2RbSBQnE0ywOtLeJLvqKQGiiRxTYu9
7B9iiqPzO+ovKtkLw07gRQt+n2BF7AWcfIWskVg2Tj7T5lM8izl2upkY5pRx
2tILWOLByBfEPwcVzr14uETOeGQW+6Sy8dnASfoATKr69rWrnbAT/Il09mmI
yFASxlAMR+namHwGz4y8AFblcU2NnhUM3JaKS/vaEzb7q4zybv1MY3LZqq4E
Q2Yd0o+lkoUx9kZCmUDyr2914TOqrxRjvBgk4tAeRfgIbK2Q0A+gAT97rvUg
vhi9gDr3B6XeH3wopDvcjdm22wgAQJXwHjTujorsxtGhRaKPl/hy/GWN8Fyn
c4owHbWWK/fXo8u9amO7ieiUJlFU039Np6LiI0L9Kgg0TarxEm5uFZQ+HxmP
E0msnIS30XPdBgAPjo1WhoGqVGjLxbCJW2hhpCiGv7cIjOKszoft/ghtBqWu
VZXISjc4z7wJf0xQu+KeFMcyA8CTdqc5z4PM5Gk3J5Oy5wFiHDIe229neEiS
aFgew9azg7iH8eSUhbtnL1ab/Vm0VFdBcShwNyQteOx0FLKG5X2zwTXlZYEw
9Us/IfEEVoukMk5vipgXp7Hhx3dVl0pmPdpRcpOowjLBjiddW/A5KhmMisjU
AUF9sqAiannF/3tJB344eEGuYM3lj43fYdXd01gMhJdfEGno8bomPjiwqq60
4Yk/hOc3gwcNvcVtSz5BBhG57uqqXhWL8vbQ9AuflN6Wmy2yQNgT6fAKWFOI
v+e4svPfemLXMcdZjGqiAwJc8hg4kVGpdIk9gemDN8yPW84GfQWk8ZiP610G
1jFgEU5uFp9kRzmCxRGKk2J6bTFPpdP8yY/FeYEVUvv3qCMvVqg6+WXOr+U0
LyQLOTz1Hg6hwU1W6/68X+yVtCBO0m6tRu6yHe8iKAASIKXbeH1peHfpEDV6
fGVlB3hTGNfsdRJ+fK6rK/q/RvNnSq3FLt3yt1hn5T1u7EogHtr8q94lzzN5
azaQGnD4Xxh8zg5JnaP62LWmKPTeyVFKjWaABNqq9qJguqDMYCZV6gRE9NZ8
9Kx1ZAqEIYRMW15q4Jtij5hYauDUM4yV1aYGtIBHx35nZVZ9atAYn+f5l15o
3eTuRjapP7wfZXVA7FAceKx6Q4SRzJR4UbyVvDis/gg+JkN8uRVP6QBMJHps
FD1V6W0ECxg1kIZPTajOx/qTgnXbF0TOCoMetm062WkkyhI6tNLTr2sb347u
cW4TyTiBBIgYdlRPdwBM2uXzLAqjsRMHySrol5ccS87zmVx7gFJRPJfp3/MK
TbLexVZzriP6Z3Gv6vHjW9ueJQ7XjUkhcqFJfWBMuIaFANsS2Wovp4lBRr65
uEJTxU9UraMrLitSwAwubhoezIGkab4JBLX1PGzaFQCkaggPqCB6N2sc6Koi
fG59pk4ZRyLUKz4gcXVf1n2Oq1xc3dCyb/ZH9wb7fw+RLFcOOx9fWsVPmQg7
ZKFXMuZoS5NYD4/pks3KsIz0ryiBOj37YvcSN+aFGJsldkqASXddw7e6MI0P
40pNXw8RmscvT2OAwfzWaW8Z+77BE8bH7MKxbmh2fmrK7l0YLY9pwodDIZae
2z6pOfaePf9K037P4FddE1LXa1D0TdkdvLdtg1hTqqwWLpHJ9YcUuU8BzfIz
Z9Y3QccNA13p0n6+zPpsCsdXmBrXig1PKoTKjsmvZsWbeAGRNHh+J/hCDvGJ
dgdoz1NLKGUMaYW7keT1urEq5yiiR3nYRsvbH2Ul5W6HNAhg2TWuFOePgz0A
aC3I5bXckiAp/CtbALpX2ZCCLkMvQWeUCrLFTCgSzJzNNC50X/ml5g0I4/56
xKsMjeUyMtUuO5n84aslv7uMSVS4L2ZRUOQ1uLkKZnom1fguVttarJw/bmHe
LXPpyfk1HmfXZU0FTqaMDnd7tgIYySv2EpptCzEfP7Xo2/oZmrxfXL/jOZLj
Bjl287VGYyyAY6D3lbXvDppR7bb6981xPUrKhjzB++7t/OVSTYE/BG93nGhm
E8eXy3MykRIvem+GHHamllLfwukbtaDkAvpqi/CkPzpzF38cx9ecciR2rxjk
vxQHSAlvlH01THLw7fcyzMdWzP2WfzL6DH9eI4Nhb1yyYYHBaMsZRcn5BENw
1ygXq+32s5o0kX+ORvVOCEw+ZLVw96E6E0LEojiXh7g+BHfOdCq4DNqbBUKl
5UEgu/f4fyQY4jeajSfB0HMMMZvBJM7BWBLDe7iJ/XnyZUr7aSR5LbSY2Bnr
SNP9NhvOtVs+HRjc9rJn1ADR5VTiOxlYgxrM9FPsU4ffcxLmULBPWppV6pAC
YhS3Acmb3kkB6kmoZMdL6FTwoooiQzt9y41x1j2b74MzqOaeOYmCqsxUAqmM
z5wWz4Svs7tQbUJca/3qY3b49vUrxCTmDkHURDQ3Ef1BuEeWU0oc4N3FaF8H
0Pl+5MgxQLNf1u7djiQ0HA3NVvuyPIOR527qj/vQhu0/ZjygjedtmonehP2J
R+TTymAd1sVC2x05wxBlFccQBtJ8vhOL8sVogw9/shJK29K7WUSlzcT9hwGy
39BHV96solmFvNZZVfSxjvRXlzcb1CPefNQ1FSVvFSgmyDm8bFmGiPSdddub
dbR4XIYxdEDJbirO7ao6Kamj1Lyu9lcUR3TULzMIVaFs8LvYMlUMFQD+j2pA
ImipSoKkb//a5ZY8cS8f6NIjo2Xze72i7YsLIoDYQt5rSDvG2+aDfzwt2ZKp
m5N+DXPgERscDN+zdzQg/6vsTw76+pMrPdzWshLQd8mPgnIO3kEtkDGssnUa
5HaNYoDImzDKFZfeg+EpnbOQ2rT7Ha5P3ICsxrXXiqRzZmEIjMMkis7vqRQS
nK15Ds9FQ3Fhh8VVkA2nvcwUuWssGihTZCK81+kCcl9C7qvbWGO2PR01gjDg
wosSJDwG9EpFkWkx68JzKHhN2oWFRSsTqRL2zewttdBvQmf8w1SNNn+Cy6IS
43+MjtS0w2d6Vm7525hwVJ5Y1NqW9zTAAtLBGHxJM+HOjE10GxdZm/5zqsMd
5yVaew93hQ0cZPDh1tLJ7qHMHF7kQLYIBSlbMKW7+Xk1jvxfd85SLwwolRnz
gvmAEp/LsyAepjrdwu9IDJ3FXk79v9tYeRxodmQGZTN1vGrPTeQ+AaXCq3pS
0DqkRXpfDalJd8tq3Tan6dhOkF8Ip0w6VJoCGVlQgrq6JAm9Rn91pUD+7QO/
WGRwYZm0yx7gtfyBIurEMQhZOEeJC8JYpurXJaMYQm/BJCLQ7DDAla2lhp06
TV+nu34aqoZduPFWFarfqVW035rtrBYxu4bHGLTOsnry2XC6Gg1TgvnuMLDS
amj0n2Ua05hc7y2K9ZlIwNPdojpOU0NJYIhUXHjy+cjt5/JW7/UcYUzWRLR2
OdZoPAZArBmozztQr1WlZomBviVXM7GHEejw44knU6I4koJaUwEtm3CbzZRx
mddYzg6qCSudxAZBsXyY0TcbrIctMRwqm6rngS7oxu11/xjUtqHRVrlQPPKv
2WqlYVvB3ePsnoH2JS4+4/R9hf7QyeMUlV1up3HsNpNg4O68Rg/bdhIaGhyM
wB0jzB1y2qrbuAH1TmalHEcI286PsU40SS+IYV7OO6HR2pz/sODe9V0RDhI6
unN+rEk302qm8EfyY7115jkS48ZIfcne2/u1RpPgeQPbL851veH714QuA8/m
eaoJd9s9r7rhtzEjAMaKo5CiJ+2ppmtK7iNTBLh9tny/uZsQXBnw3iv9eU83
EPA24A3GX4bQqxWPtxd+pLKhXu5qOC+kEsell2QNfkugVpJiEhyFQe/2uZNZ
cxvZGqxusHBUj+HSSkTG+VbeUyMLlHhTwdHeetQx+h4aoQSxKbi/Xefwia01
g3tjUKO2w65ZO3d7dRdfe5EAn3iw1MnuHThaw0y0JkVSYhFID+53dJJuNwjw
4LPQHTovI+8iOsaTEoE7vSgCk8taa5LKqEFNvKuh3+ENcmSqdojKjvbr+Wy5
o+/5ZHOoPYQGR3TWfNl4TgNAWZ9prdP0WgCtnkx+WgZK7Lt6/YPWpufbyx1o
3o6G+VXgM49887a7liyZ6Px83J1LyRHCAJyuJJWEQw/JdjMK2KQWROHp+Dno
a+gHdvTPUz0VV76H5IpztB8ZWtoTtLAi6P5ML6DlxR0e4HK0S2vSRTNkIjZB
7J/FfxTxsmSVZvyYFOF9B4f7lqMxhR/8mECOas1BjCrZyqQBfVI5CZ2fOIY+
oXeDeD9dpfSLtWIF+1jVw7it5RSEWjKEaMoLH/4pMPH7g3GGzFegMEJJWZmh
vl1RDTEJByGPbUr0fCukrSmQQxZ3GqaBgQXjSpTuNYOv7jM4iOdKpzNzYye9
O8Y6Opy2ZYcNQDUm+zjYwaJmP+Y3wlqt33e3CjFhoIQxbymHZTN3uBp8yDeo
NZtSsskal8kUFCYaffmR88VUzagAxiWXGVK22vIE6kHnxzkPfLieRoqaPkHl
wpdP3OIw0mpy1sjiyUx7HeMjH93SZjGv8R42FvqvFpvY1eCG/kmq0LY66+Vx
dWHN/OJ/fIgWLYDBMnBAzRk4vKOqPbFHT5cm15V0oLFTsKcW0nl9P0vQgKAq
WesZRb1OD6ILUsmOblgLpcGBNsqbZ/G/mMopfMQGwmnUmI9NXYo4L1YZXqy6
9MILUtbB7Yx9B8LY9oN82G1PQYob6rm4eetuG5z5xmsixbjPi3vatDYYIRTh
0ICDUkU3xRPw9+aqXVqADSw4ATVkj7Fms0nGGTyONXeHE49PH8ieRNRHu1G5
VmQqFnkMG2tJkGYjWtn1Jx/huSt4h22M/d/SR8Q0H/j4zh3858N8q3zQ8nVg
XT6MWgRLgrTaiCxFjK8unSgpNYd8yt9pmCpkazuB47ZUnDcZPeD/NlcbfBV7
amglIq1oYpdqMaA7tgelDXdjyFbECWLR/a0f4E3B7VuknprYuXLCd/jWjbqS
4WYOX2SWQdcMWRjHrWnR0Q8l7SpGi4cVgt0IXPLY5adyH6Iu0Iqfm+rC4IMk
z9f8ve/g1xe4KTMLnWoAc8P7LOnMcAEeYDFeAIpXCnQf78bJi27aFRFZ8mdS
kViqP3PQ20BcLQsXN/Y1l9LZwLVZKt+M6a8U0CTCruTi/JiHmqRMkXu3kdTH
FMqcPbOUca73s1mlg8Syr3pIRGBqUPbhAiewt3SWZZPBInA5BO3Rcg7a1Z4g
I5svSbKEQHg+pG+39/PothIKaxCucJf5yA7nOG3uAAWebnt9B6BIZgZIv04y
r95lJZhSNb5DpYmCsAHjrCmgxFkpjpKTS9IuK0eC5WMYtFdIonRKaC+RtxtS
fuReijxFQQh/UI2yBxxte4xWiZcmNq0oErxzuIqAFFqbu/8vdQGk+3Wai4ED
GD0NIlaVAb1qxrQVhCSHgRE3vPbHpzLLQnaG4QRYXGyeihx1HW94Ql0M7Std
W3hc/aBx0EYJCWNnp2CA744urZ4JS2tQQK60ecAELMTlioRBBUyOj3vXUkch
FoGv37F0xidQOInHNkyPCWV4gvEq7KmUv+zSRYIBB0ckJDIE3vNHKls+7T3v
w3TDGvZJE6SLLfU/xx+Yvpv4sWURtxzFjSKhDkXNNC1gqKTNArK3AclZAxkK
s5PUO4/t6ecaSg8v5B7vKozADs5kpx3d+YN0hbpNnuOz0EYf2taMMtAiIF3C
Vz2szJL81EnCE147xAykb6BsVeIlR6NcpbZCuvOB9bWo4p2frHPNgaIH+NMO
x9yA2T3qaSdyMtRZlt9wps7TADpaKuJDVEVgAPkIbzcXXWJ5B6u4UnKzmevC
97VDi4ivXTtClJidevlcpUZ7TC+l3fxkFE5KFMrFGjTdOwzrQIY6Pf249LiM
m9W8JPtd1THsu6Mm5HdICr+SbhHkMBvslx40e9kMvb4YDXNyDWafTb8MNdyw
0Cbq3NC2YjJmz9aeJ4Fa8QKLM/GT1cjY0cJAxOzcCT++sbg+eGt62hBOZtda
Jjjk5zxyoRnaaUIdJGfBqTO6sxawVyw0aHzCIYCCTSMBJxe9NYkK+RvtEME4
9Es5iLKNcRxzKgTZZ0qqMRFJG4hdlvVBkUjseAQRe3mXoKjf5rcbjij68OJp
IUjj3YDomZhDk5hfM/6L5oJjlnX5+5wK+GSHGL8ASaSkFJaAvIG0iNG5C/27
wvc+wv8AWne78eGobURGQp48xCB2RSlzpkT/aAIzC4F5MTQTeGTb6uC++lCu
fE9T4r4VexzOi0IU6PqBQorApD3CdVAAs/XdS2XZZ1sQfSTFozMZOu24tKYK
fFaTbQSp1RBX6Oi/23b/lIqaq8k1L9oY8XnUBHlaErRxiQLmL4mygptOLzC6
4EUcdU2W8puw0aAikGU+TXX+BXwscjHstid8NUwsf8gR9m6fm3Pwd/AEgOt7
BG/8ErIgvjPInn4OWvEyJZNpXwN2vyNXpMd3yYBFisj/wolKQFEhry9uhtZz
GZnI0aX0QPStql1MHsqY/Gpkz9iboW8Ko+QHEMC3PudExxtTMb5/q6PHCJ36
BCpIeIlwoc35B64x5dU9xVu2gQjKsYGloFUlg+xKd9fnlyx2lisUkzrapoMz
QD0ZST/HGRPdvzEiywLDIsHWl9ZJFlstqXo+au7b6wbRovXrTwv4p8SNZjcT
9MGHDKFl9k2zOtSC3UWzOghVHxbomZsAiKkSmcaLuRd31YYB4hs3QaSPrx5p
s0yhe5InxD66hqWPpAG9IfRL8jNXuL/G5flBdEzFcBHUvl17/RKaiG0v8UAK
7RqH/aF/dllPW+/jjlNVUqcFRXap0IYzg4AJD3AX2dKtWnCycc+vUCqSn1N7
Aw6fTLgQQ4f2krYNCD+Pw1JG9SD2mPUiTNhvD5p7VxZa5OV6c/wWgJPbl+iS
urqOW+cp+aUee9YZ1KqjsS0NvpvXAWc/z0pMFSxI7zXWRSUe0URFYTVfwXVz
PVImR+bDdmU04BvD1S+zL8fNSKTxItFKKDMVJ/9j+pkBN6kWzeg6sFY9BRUs
ZM0WHgaHQg9/GhfjaXTeCAbNf9u+AzGaEEK2lZUKRaU8EgPRnSIFhssMHpDc
H29JOkNcDR/ptaI1sMG60q9EV+3+6QkM1GWdcGKdIu3+jdpNxq0Gc1ZtEnj8
6N21rispKTRAd+sQmE3JN6XLQI5s2BR02bMMk7SfJmsAJBR2o0kgkosgRSGS
bqc843obuz97S4KapMyq7uVfUzlm9iNdnNRw2wGviKphR9sEb2d+R94qVMEE
RVpIz9xzYRdyuGiimCczmYXpLGqOp6TPHLUkcp75Ao9s4G5gKPSFznRzO3iA
1DfsbrT5T8v3+YLKFSXXh2N9yVQBZv1N5puqTutTE3SmuDrUECn6ZjgnAHKG
oJHZAKAlg/WAEuLdKuKSuCHNl6e2b8KI2LAntjG6hasLwwzijAQ1rlj0UTf8
D9KClKfEVbbOhxPD/8kJVVMSFah8p9buNwKOwgzSBlRxzqWkcSxIhOChhalx
XwAhhw1plTIyXSYWwFPLkU1URFqR6DU0O0dy3BTm0yBsH3YDOlVDrhiwZLVC
XEcbxbT/+4hqy1RgOFsT82E52iBKB7srVQmjLCQ/1FRU1KTmLrgCJukRHTmg
1kJkWffLfHx6shj3YRySERUwMyHL862CvuRrCO6nIo9rWoVFeQMJTFl1BhE+
Mi5FurN67mcVYkFxs+0Uy4o0pkR+RmVP0Kex8fMU5Mlqq5k3dAUlxCpV1XfU
jo9a+uy1V7bO1pmMuq0lqf82hapBvlq1mxO3UbKjTIzVK/g6DUeUDrgyo/Fh
q1Fd22bzsebD+POb4nR1SURZ75qLgA2OdzgxFUpI1ZnvsETbvY+72KD0he1+
bfSiSNB00dMY0AVxrIcc+6HJbucptZf9A8zvLDGgvGRBFhfCRPbH6InhgOVv
ZeQaP6gwweT7787kKZo3lxQXPqX1B40G+slkA6xRhNRlzi2JwmbVmMOLb2L8
Z1PaCHn5lNxEGYXXE4ffyTBMhtSiS3XRrQGsISX1SLUJ56eDKnzMhiWpJ4zf
ctX5STnGgy90nxioRHbAptgIeijse25p4cZKQT7BTCUR4XJ+jyQmSyhL8Ysv
LjR9ka4N6TzqSaSmptMeE2TZ7ENgPardlEkRFzUr4s8pNZ4dfDdSYXo3ufZ9
9bWLxk0kNRJv7Hu2ub0J3duKOKL3kVOJ34s3OnVTZAo9b/57sPIRWeKuRO/7
JD38999f59TuVwwvbZyeyaa3hh7PgBaMeMobpiDC6jculHIfftIfxAnHxWMN
WZfSyE90ZK10gr65TtaKpHHcQS88y3UYRjEpjTNQHSvop3Q7nAjsVDVkvcWo
uV8JLjbeDDaIxDU3x5TZdeuFGmmFj9ifOuoR0PrOv4Yy7mVOM5phbnzwYth3
2RgYL8ybgjdboITveCLmLlYZdj+rNTjTqjnXBfX0Q9alPSgSBCFFTKIv0Nzo
Rsu4OX+pInfHWxwlcjp+DoU0EW9MoV59RgSrT+jwdDBlcX0MqDWmyZLkOGiN
qlRc2Zf22zxasgA+OxzzvU+4YzFIFSGPC2QnOQG9MCiO+bU1t7kYGBSCMSs/
jRDg3WgG045kVbYbZWrmG7f+FSjssDJbs1cSNpM4JkTz7R2g1L+iheVeoGB8
jp448WOv9weARcLYEOk7l9l1rXgMmo3y2LB4PA/r+l5L8uU60YLE1RaYGdcj
2m98F6Wd6dRTv6PtenCaKo6g5Q6j9BFyQurJ4W3k472aim+776iB7LubenKc
CXyzA2/oHBNxw6Yp+9IlpVX2TQY6CboTlIopxYrsrvPT40R+bohKxmDyVRIP
M3pqvjDgj6xwHGbcLB8Iu5/Dy1aZ90hPmnd72UhdPhaqeRDhAuuQ+pVGRmwS
73VzgQOBodZHTT94h08ELziLm98UpE1YpOX0A6/1YnzDIiuoiD3TTepOpnO5
ZhcFv1oN/IhKj2aTSOmUzqOmpf2IqSPLA5cwfcmVOxteSSK1ONkoPKG90aDD
BsmNlovEE36be28ad6p19RPvhZiAL+ElCra+epAtmhnRrHu8kTenYYRYMK0+
/y7rF4hDG1N32edZpEWiCRiG4d8GjfrePiepTXu6OH66ekoEJ6KOF2lGcUJz
Yjm1moFize+zELhik2xz/K2Ra+Fqykvy3IclOOrcjFzaQZ3YBGdQDD/IdoZY
+c1byuHDH+CxKCt/zPFFx/XV8donA5sJ63zZmS1Zsz8al6TbMEwL+3lIwYaq
E+e8toScMIFKLx1351N++mzewIkxGD8R8Y/xBYJlCPmQseetPUhrJkPGTE0J
HTzkttIQQuwAmu4tKiMNUxqiKbI/AdLs5Aj0dDr2BSCg/4RKUn1/gM+K4BUw
449hnEM8Vvj5/DUK3+HwgLFK0OikTkrfdq+SIYz6NdWvkzLwQwVkNjD03gZU
OQJBRrd2FO8BQy5KPJK5KoSAimqh3kcIETNYJDjNaGywcx+awO2tmC1hsbAL
N9lVn3anBq7zPzHBqDcdBOxaKlxHZpuEdNl+5hfUoB0y3Nblv6XS6IYZhpKY
EuVWr4GMxoqVkaBdO4yF5q3MSe5xdUqq8qOOjE7OrdlWRavFTNkBWNHIEzUk
WDsDYW/cxV6A3DRuOBBoq2EnZxB+PECYUmB/+zYTtH2u3owUIFY6Z2XPQe2o
T2qUD3LMdKCK4deCSJMpi8cYBwCoC0JDJubknUt0aaV4u5eSye+tjgP2jEKo
gG+AScNgTfuwpwy7aE/BK94RAKAkFH4rqCvElxU56z8xV+dju6GGO0S5ADrv
lzIuJcKzmg8e94N4V6CHLD3bHOZY9Jg7nVAn1zy4hx7jqj8L/99kF6QIxF+G
+r42gsR5aRwnxG+ULUq7j2nNadr8nPS1/Cfgp5Ubtq3hv0HwAVA5B0sK3sXM
T6wrVsArSBWVpCVzgj6yGg+sJC6bLJy6AUrQhgj4wU+j5C/ST/soqzTIvR87
Rl9HdpmsVbNjFdFiEMe1R/N2aySUyB2Qb1pmUJZeBfW0JiNOZ3WrJpytNOpi
KY0WwHGihKkDoZsrmBhErClV9XEoc1rblqhLOwVfTdmYQb3Yq04SEdZrDJ18
YWH6lYXQ1VuQuTt2UQB2+vUrl0ld+8DHXs3nrbRse7dNJwb0wF5jzg++VAAH
ldgaolc+Yq76wsawOYfIMYbrJUFWeNePvDjhQ5gq3ymhydgTicJyZJeCbCaw
BStZ6ROXRVtxQYLC534c6GcUMP7ePMf/xL6sXO6Z0grtXWfWcq7FKRGVcXQY
5iY9ATa5+TUClf/fWTPheHT4zk8uya155oINq5p35BCUJKzKVwvSm8F2VAMy
2oy2DJGC4IB8/KI7aHSwM5bIT+xtwcAyOY8CZ4rmUJt0lJd6mX9lwn8GHIyH
syJjyRSK1kq0iwBAon671MRnN1FiNEID0ob7zzW0RF6hQYUcN5K/1Drm0riK
ZpFCRAcL3KtbfH4lbOSm+w+ZAc+o/86QKes+xp0YwRitR1m60FvodQQzSTPy
gN5KCg96HT4Ck56wKSo3ENQDKspYEzHF8/LZvWiU1VshEv6xFGzRDCLvZF1Y
2FntVIsEDVOlxvAyX4h6vI3BoPIhnsgdmBUpqvXBweJzYaKIAXfkRAhzXMUf
Qa0EheTiGPo96jaKJdn7Po0P2VPdAPi2poQ4NrBz0ObGI9EdRKU7E4t3cmTr
rTDBqprVEiebcZcKtr/Sl9m6TioSiHaVpc+vZxxpfdRD7tUTnnt8IGnL/u7G
yb9Sc3knB29V46ZVH4l/1bsbcQqNH9usKqh9hrfV9icP9UPh6P4hORXSBG6j
GLNHEYB7OT6kvS1aJSsUdCJP4cBzLgiT+Qn9KpcdbCO5NiJPV8DAyWhTpqLN
IKoEM1OFlTZMNx2DtF2xVuVbu+nGILwA+Z4b/Pn+qg+aIDhTowh6akaQStZ6
EzQYW8jPxTm0W81kOB/nrQ4w79IkEb7pR4FjSHlUA5bKPsKWY0xEozTD32Bs
0davXCcN1hX09SMRJcGsIa99hV4e/3aOWmS3lzd3tVfze4lfr05ZGhXp0mIM
VIc0120jKog9nMRO7hzlDUg4WZELnqUkMeZhxTBNZF4MycfAOcFbPw6ZE0H6
6Iy/6UvF1F0guUuaWZin69nNEijifkC4XGTW8CB8V4MXsG1UdA41wIzTCwMy
XZx+uExbFTg6oWdGq9FBVa8dQ6KUQvpcpaZr0FCyUcQ/ox+qtXKRCEz8RpGu
AoaEVPNwn7ecyvX/fXdZgVseJNyrB7Dr5wF6BXRpsSN66RAPb5CHEDhvJtyJ
g1LiHR2TtbJzy2EGG+NH9q+G2n6aVyLv5k4/b5SdWkkPwRRb5deR0R4MhZfQ
Qjjc2gNwYysaOnIuK1jUb++k4sCgRg1lUcNTzzSTVzt5b7KYLa90AKqI9ylW
i8fYFct63FBgSYJUI8WGakH12bfJWofyd+LcdFygJQ89h3REPpoT0qD+ljj+
HXDF3UdBlJRvLMPvDfVnKIOQbJMvCtqtjSKf3XonRIuZQQCI44h6YD/sFeQ3
ydr+uNviH9w+uzN68hyyRddYHFwhOXEP0uZt+Xu5a9HfiR58nUzzMHOBRaVg
tdJrf3QQ8N8fk5OOCcH6m4HqRNM2uNZsQlwVr+9CTRHcSNtSZOhNDpgIjlVi
zOm55gfyDzdaQtc4OeqEpdMAggyWjsl/7AdAPlxGH68FQKJLCXVcWgcfDrEQ
NKe2t6sNVbjEfnD05Fw7X1OnRkvUQqkHdGa1MziB/WYlUA4mA+fqy1Z55RtC
ycfWHS1JBOkm0QTfiCG7KYamFdg91Dt5oUuKTTc+N7DaeKUxAedcessy7W9d
gUOtwKOZ68jv3NdgXnQu1db0mdOMcUBbOREs/SNQ4oITJxleb9F0DJN1rm7E
NTjoOnIZ0z7RMiq+hyf47M7yu+6Wv02smQIIWJWT2z1XaQ2j3xJZDVKJjm1h
bb1pzxp6lXeraKD8JB5uEAqIRcGmaD1VDtdzwybXpftNmTJXpYuSpVccsS/L
XGeiXHzZJZfeLJcMjw7nnWSMb/ES09xKfu4A+n154sCqq6J06wFKuvUMr4G0
J9tP4nq8UQgMjxTBOHEGPvWvuJL6EIhSz4U0fYd8fG+QGwS8DHakINTc+XnS
5qmIFU8FSiGH53VLjL+KVY6WFz9TkntbZLUXyfopiBvtbEt5ohP+2MP0y1nt
tLhhRDIi0C76kYQeW7wUiLtIBXqSukp828BH28AZCbHE29A60gj5M0uoI6r9
NPMBQOWVSvW5lzmFd24Ak5eVXQU38lHBHt936wvEaoDSUTRo8eBYFroHFmF7
SkruklQ05tTdo4uY7sndjk2Hjdm4Efsxk3L3WThUlzKs9LjDm6v4V12VnoYx
yYaUfc7zFgvoDhOut351cYwy12yYaSJms4lGQ/HFuLK8KsdBJU3Qyq91/5d9
c609Q/FPMQCoQWAnR+SYEkGz8ydcv9nz4QvvthWkTwTTgGpKgK8EYFESiH3n
sEsJ3CRPE2iCGB/qN0VCm9BEZv6HivuMPfLXB6t2+QbfOKddkZ+/MWlsWjMK
1yq7r8qcHqGmTtwZLdvNyIODBh+lFM16HgjfylYW5zZfcjGb9mcHDn+zoUxx
2/xq90Lkc8GD6bPfApliEQUB+nlbqXHXEl6+khdr1ddr23Xu8q5NJylHX6fI
4fd4d580kwj/Hg2UV+i9hE3JVodMDcslqqRuaysIxBz86sRF4U3AGAsJYSbb
O51uO7gzXpJOZhetBIZ9PsGXgbMCcP7W2vU7lOyzh+E2oZx7X2eH96rqnzpN
+HqHpzKjI4zpPhgQ/8cHEiOGiuZN92+NNYH2BgHbN1ynqASfJgT/dYLAE+qN
nI/7nGeI/Y3Afm+6hYmM4twIw6g8m9JIYfkmr+uN4i3+G64NMkl2YCJEUdPb
8z3OP+sd7JrvJ5mXoENrhZ8pF+DZt4YRR8GeyhTHeMIC/3mS40zMI3Jem/q4
2WfZMF9ULrZxPFhYKCf0kmIvU+k9U1+Oku7UsukKbfxt6jDUepC1QxTWTNGL
TUSDVD+W5l4Y1ScGe2JvKSBzHCNjwnNuxA+LhN1f7psuNeNLXuKCaqaCH+41
gqHm1WdE/cpttHMZYA9forZBFStz8tvb0TCp/vwMthTuKlxQ5q7joyaKlaCj
RoPI/8V8raqVOIXewKYn3Zd5kQ1eRot7SmXpKo8ZVml3IyFQh1E+9ees44jv
yoMi4KfxWinMFw7UkO84WJwWHVcj3CUNKqrmkGXBlzzlDCc0qMWMmuPjUJio
sH+1N1WhBiEXXMDq9vkaldUSBop6Kb4kISratJIo6wGnF0lu9b2XCxW5t3oA
B03TTcFS3ebMhsburrFiDNcDTE9M4BGYZaionM3tZhM+eH5me9rGQXONQ0JI
ji3MEvivQNaGdITL6dTLgIeaOian/It637Q2kLqEl4y+88owzxTAiC3wTiQa
RFTeXn/IDM5nWQlVfDnDgiWepbgyuX5ujHiTvpIOj4SxoPQSFbyDlsY40H4n
oumyJZKloTbj4UUIg8sGnBNKsnwcKMlPqRiG4SDHUVi3jm8xEcgn0VHcOOYl
uhZqtZM0KGJjRjfW0IiA1RqA+bUB9N9nZB1wh0tJzyaRyksu3KcBttW8gC2+
yOWTSk+TDhTjtbrzQC8L5wFr3mZFayTAONCL81sFK6+vDNSfJ0x4iGROsSEw
1mO+bREqj1AXq5idoryGFBpb2B94+1fvPEbFeC2HrkxYk97035fpQ1+4/9Tq
2TePNqbLtt8QwfM8iR70yKv1hjZQJ4nmJfmWj8z+p+k9kanx/oFmN1qKZloO
dgppS0qqmb1KxBeeWlbm2o+/72HzDOHBjPMev0ttRdgVSnSjI2ILLVY3Kbn+
Nv9JiDJ9+ka4MIpESTboQwyORbD5ZKRY7MQoLhCWiiuWWB8f/wMHPg8M/Nl9
sN/jW+XvtNmn5YHcU0VzOsGYuKzCX6iJZ/cG9Q1vU0/++uydcaCgAUQqS8Ir
PV7gNR2ZV3usAiGmNLIWAHuQEE+M1GXipu77p/hayuqcIihgmbAWBUP/lGHy
amEalze1SqOZ3OuIaKWC1hkBZobjePVDIpto41oH1Rtq7F7JIPOel2sBnycN
ZmTOplZudEPSj9JZK0xMyV+vf4ZktERITYrfmxwlFr4pkTQpgZf75OQT8pTQ
yo6cTfS/qlMTd9V3tMLceLmLK6mEah5iHH5He9gPtDhNFIxmPsMPQesXzOsA
rjEnyCkamuOom3AAYpO4sFcnjE3kwTyfZaCU0lqBdzQ9DGs71WqWkCDpa9tR
hsYtoemPB8x/7FllTHg3TDmSndVPcBT/n4svN5NCVHz6NAwCDK8xWqabLF+g
6kfnd2TUtjMYxeOhSa9miYbSqIHzRofrlX7WsA9sYAscJUxV+KBp4S1w5VJw
xtx7Fp0sFQ8YwFkkea/qMx6wEJIDJtVE7ryclRxov1+bdQno0JPTFHZiwoay
7d4WJQ+5f7TU/pBoYPbU/EkRGTERfA5EWC/wd8Y3gOIkps1w/lsr8R1euHjK
LqQX5HG0TrNd0R/BrfABfnvtm74yvZoznNdNtOUYGRa7EKG8hPnvJmRDm5r7
vUuu/SKnOP+Z9/lltNzVsnlSAU4qGxj560kyAuaPmZBbTxEqo54Nk1xZTe/C
pmdNIjd1TfH20XHciLO69tYEvewTQTMhUrzygSW17jRqSAJ8E7saGpdd8KyH
tpHD2xzkoWUOwE2/DYzphSInAwoPG/Coi9kSTIPmfjykxT991lrQTxfBAWiU
3l2sKo7Xb1T1Svf0TX0WvCKieUFG2+8kn4eiUON2qPjhuBxtVGfyWrZcCFaa
jGfDs6Fqyevueab/ZVeVpiQ4hxVGevBLkhWpEZMamQvdJKkkFZMWYG0KFITQ
rqNXqozZ+YoMnh0+QErB9oHQrOK8uA3sVqEBTEDbvaOWMkJcVuXKeIRmxeIU
6XTf0oa7Qnu0B8ilzGLVqUt+XGyItQowyBUHiJdBzuf3AD2+i9vH07SyHaRS
0dsQ5sEvPvg2xUECEIeOHQzekfoy8HPH+2Y/ZEPN8dFKEtWuv/DZ6CsatvU7
Fs3i/piDwCkXOkerE5Je8SRzYBq4TUXFZZBzvjPT7rhbAOMYRwMI173zpumO
EfhOgZziQy4Yb1lgiNheppvRdxv9vcYy4ZElZssoxMlQ8OF76yVRwjaxKOzb
YoQffJZgtCBoptba6melLSx80T8eDzqb0KatY/u6ahOrqeWz0Aat8+iwbSzs
oVeW/y2V5XhtPkYMzEpAkCkdcUGtWcnQF+vL0l0bEKlxyHn08vnnbWjk/hed
ZIX1bikHfqYQqAhUwfQEOvvOU+2DXmYt4T+Ivgnarj/JFKqiiZofSkxplRmK
Slr0ng/OHRmRWdmoBZzWNomtdDx2MAk3R2plAknjOsnkCojbXOcj/2FMeQi+
IOM186QUq+WGg83f1uyi2gHevw+/AtsW/dEQJmAw3CACth7ytqdYbrlHUfcM
2oCJDPrqLS16EDMEJRUy8lZQ5ZirCtMCWfKvD8Khs1GAvF4TFUh4cxV2chGE
+Dx4vPaTXBbR1UTWdZhan1/aSzi2nHbC/h6qPdxPK+PYwuOCWJCaw96Bp4i2
hz3DF6DPkraWK56OwPxMv9y+RYzI8l/4+B4nUekHZdRsXFDf0EC62FNSiUMA
UkzO7H6mXtpmZd1dCWgJV5hAfqgrfHgpSwCVJ8nsl6h/eTmyjZnoMA+fLIbC
yvJlVbqDDsjeDrA79mBE8CU63A8dODZqIg1pH4LVlI/gsyAFxvPNsl0L4woH
tWfkjkyazIikFTbncB10MdaH6NFqz8nJ7a845t8DfmqkQpSmgce9nxbXEl3E
uNYVG1m68bnwNbVWAAHJye90akKxOSW7BrrP6hj0JfiYAidgUbnTzYwM5V0+
4s3KmRPYZF5gbzbXwpdA/93oOQwrx7Ant0Wwj9+jiO0m1omGbegnzgZVAUQC
TPbB1ye6wkBep/mfVhH/aRRbSFoqlfE/LbItKIVXUY0/vqmCyOkmHoS3LsrP
Au3WIUinlJQCSDBciZCle01BajiUM21lqg7DwJVanNkbxKgkLPyavmINjvZR
AMm5WwbiOKO71KfMD8bOkRkqCLTKvOb98fbQmFXyMZPnv7fSRuKxycRVtYUE
vBu+26hEOgqyPR4KVCQhKc1eSLyZU+thoD+nB5JZ0/EEzfnAmMiWlkTupok3
Cz6mnbeU2tvfUgPjfROrulbPbMDigmmjDMZb/VjZcg+zv3cMywduf610plfp
4OhFf4t8wkCQeXlxHDdy//VFRSGCgu5e3p+O8dkF1Iju4EtPxydThQbAUbM/
lotpDPl1tCFfh5udLm9laCL5FUpBetoSKopd11xQl+rs1Y/Jq/+C67seWpAM
GSV+4+aJywll4teURVbXhm3xPMHsRPBaBB8lgvKjvhUMjyddZbYxPw0MF35l
eQxuWFnAD04I6iL5cjmoemgsfiOUfSMx256mHANZdVHfyqsCNMjPH4Wxb+gT
ghQtDZmXG+Femc5GEyEr6EIV0wl/yWh4moN9gk5rLxuiiIvFz5ljtvExE+dz
5fsE2VESc+MYIYAVmH/QgMkuTzsMbcqmjqhYz1xpdXuPcsPNgU98wpRI8l4W
1Y73M4u1VI/lvDM6KSFYv34cxtg21tUuBA9dmqAMv37JXWLzoFrLA2BkXpY9
QXpbmX9/H95QgeyURUWpg8E+aNT68RmibnHg6Ocnmh1VKs1WQLW1DfEDmcoa
d93Yol0NHcnNqiqazD/aIeGLyf14pegeT35iPTUq95nqT5jnQMihVUHpR/mh
n0L4juEEOUM77GP7e1lpBtKyAjBf48yUmjbbJgfZN7TG/Gl6F9gT1py0LCSk
rZxIB6KQInWwQeY0M+zcwKrUibSl3PPlxYdQApXXaWl7WvxtuACviv3elfpH
RIs2h7m1sso4vnQ3T8ouVPvcIGSCLSoYNWRML5D+DoDCzeKUEoKvU01CA3Tz
G2In5kQfIlQSLfmnZYLDArW/TzDL6yIwlgwVXIrRlvDseYTV70c2FPmF9ajq
RcEXYGjGgXFHLL1aywH13XaBAxrXEAw4YEzWz0Djb4jCt40KnLmo626IRWQn
kRX0Vew+NMNN3E8YOa8ndq7zrFxw97dW47mDi88W9X7HWdbCgySKgMnVcge0
Fti6G5PWIaFMco5Xvhk4ksYeBzGCRMHBCeopIFZ08gKN9PkoSyERmNJJOHUH
4y21ZBha/5Fz+jJ2c0yNpodNZr1SoyEZaZeKw8CqPUJeLIuW+8fUtgn5QE/b
vw+2sO5amFQhR+n1qVndkiCYN0QhcErZZysR91SBNV5jCSW/ckKoOf98tXA7
SsaZSWEgEG58sMxnobJwVYjUrEQ/BIDmiwTtqrWEqGBGPWHt/pC5B4NRdgGt
hshaTNHserU+Q/WR30gbJOXLDofWkjE8334J0vbsjdpVQqiAYG5GduwgFfCF
bCFpOUZEzUl1MgFgRxB7DsqrLn1VA265bgAbCjP7kz7rxrib6oRLoH0ys4xl
M5pXt9eMC312cS/tMG6YJIq7vDd2aXRge5Zg7qmnmU+0Q47qiOL6sjZ6PStY
FixZdTCaN6rlDHE39QXSYHVAtTk/dIBZTi5hrrMgBCYGmw42eGtL/tbOhEC7
m1q08mbUmvT4TAorN8l2qwDwrXGbenfNVt5I9CsYKbITfy8gYeOwCVFY3UU7
Nj653Jys6a9W4mMJVGKPotKVyj6f8oc4fCZZD9KySitoOvH3DvC1lwxBU8bT
oUAxE9ar6c6SRhWy9Roe51tjW5t3qZ54wn3YeLeGCNUSD1+TQu01HRQY/754
dVN/ofZ/w+7y6CPQ2PU2EPJycO+2fc8OgZpobjKww13eYU2RvRM6OA9cmF27
U6Kkf0h45bb3jMJEXfufHOPFiHPf2peDxsLXkHjfmGnSa0BYxH18gc59gc/9
zY8TLiYNHzUYbVI/fIqbBnIKq/cd3gT9viRLL9kcqrwM/pVyXxdWxRyP/eCY
gwlvAYvDV2nTFPs/8L7AragDg4OBJxgth40qdzOEG+1vD9S8pwa6lW0T5RuK
iF5fmstBHRymKtwsPWT3aUiEEM48Uh0pbVi4mV4RGokCFERseChgo+sfCNyq
YJO5n1qsZOuoWbkQZ315MSQT7ASLvfRtdyauqTdWpOMFeRG8klLEGGdrYReY
mNYs1CbDCyyQgMls2fEDNO6pCzuUfU1kaSqKc74kBlt7eBUQyFD4KWVclJrH
6GEZjJKuQwRjaPag84R5Lmw/4J7vZMCmx7qNpM3HzfQWEeM7MDtgnKx1eavf
O8/QpGs87SEVgTZcjsnt4AVZbn8RZ0s0PYe+ldCKw32g/HsxUEIW4Iz8WN7e
p40/spGHp3+nAxTPsCWAZ3ywUXDyvuPzmYE3wsbEhgKsUYeIC21UbYfIBMsZ
Wo1k4x3lYZiHpwCWJALDyOP0YFQKx+dN0cZgT8IsUl+K4adlyAt60wuExQC9
qY/bsFvJM7dnDJQWZxmsg7yOX6Z5kF7uQW9orADob+QJAIkWsay7qQ1SH0vR
F/wnKH4MRpbHfQeJ8q1APm45HvOfuDTZfzMAgoo4p54IVKcL5jkFT5t6DceH
nctqD/vvgbtT/64eOgi42V8/NIjvV9BPxv32VjJZlwW7km4AW6bhCdK6WNCw
sgyVq2x9YPE1H5n7/AKZpzl8NjvVk1k45IcaxgYkRcXoGlzz6xMLB6FLCLuY
p7bF41gau4KdWy1bzc+vcWodqiDk5TyT/80PAyaXvVbf0aGk+kTYSvDtd7br
seID2vS4FGtTKcMy/2lfPPaAPNNF/i3uFlHUZ2uAIlncl+zNH9oLSP6QTQ1Q
98Sh1+Aziik5FsxOoiU1G4C263ZpmAxf08wz0O0BdaDsE/4YcYHv1BoNojok
Ubrli4smfBmRgQAbFcQpWV6zUmoh0xY48y+/xIxySo962hhW3ifB/7x2hCM9
dnRC1ii2MAkzjEjxQJKfxbxR/oKh3gKUftqGOlH79BdttPf1M0I67/UMPgs8
rRVgc4MaQ5rPRr2I2MnuM9f/EneiFptYlw34kVaUIDK37Wu06U8tzmXjzkNA
qnJZBys5poJOO2w8e5vzClJYegwGlCKfgMqw4Gz2dlJDAjC9Xl827w7UXGw+
P3C48NxSMamLdkJBj+o0wn5We7jkrqjomgoD8t+uwHyQhLuc/n+0x1WylJAc
eOA7D2L9y8SbiTU/MulLQYUAUta9MjkBjUFy+1fwAKKL+0vpaT89v0a4mA/I
iFE2evDnIGDgsklGie8coqzTJ7fkM00En7p1QGkyY6RyvfW05wNFCv0tY3mS
83knGSQ4/78Ybl6Sr2labCknAHfTKC2W+kNJtZfQDkvBYXDNGKqQpfgmwJBm
HvLI/loHa3g7DcfDCOO4lNmZr0TQDEtJiJ4+VcRi7Z+rCSgj2ZmzTXqKox9B
CfxKKM1MBiMfXFkW4rby+EMVk74NE8G93Fdh08FJQhE+yPFaqDKgN680ltgh
+jgJ9GvefozjteK0n/RUxZCyJ0Shou7G9Gja2/POxAlCtiAAoEYYJMDRi09t
Bw9YO+X7V8NyDGRHVu18nVn+fgO15UdsWYydOiAWtNCldD8K6/r68w6TcOBZ
S0K7AGzqyq4zad+BHqxsBJDXJlTRBtRdP1IMjEkgOJayCpQGpeic06gq1ay3
kXsXsI9njbwLIh7f4qUxCm2oXIGaAXH6bkhF0Olzgnedr0+l9mBPrpICBQd7
cTTafbwpvMYfklU9jV7u26MsmYC5TXSc+aoE4Btom5izJByB/qaJF3fXF8k0
T5LeCV7MXk6MQ/37oTwrvYkpBUlSCepeDwibV7pRZo1mS9E/61CLLBLzSQnK
OsH4nEUt/ZVk+TqR4V2EU7VK/0yMZH7B7GNtJDTdYEZROmzW8adVJtcnj11v
6VvlGZEmPXzSK7JMqsCQ6PcvGaGZl74+WjTSeA03SGJC6jYHRUFk9cW9Pi6Y
rsMyCxnJMIDygzS8DLIBcY9+11crqZX4WJYzoMiy+tSWfWzcXJ/TJTHF5UFX
tIRNXVKB77iOjDvlAf2RZrJ8P5ZALzjhBI2t6qmrHckZxWKD3WoU4HtxiPkx
MjUjv4Y2kH4DbBDFVH5fy3hWSgGmGONEISEDYeN2SHLpp4W+RwsALCtndbTu
PhIFNiqkvC3YsUmHmVDmybuHxPiDtlhKlCmrJ6UtAmjBEqGNbX5+Gjr//cE8
vNmdk4LkWuJEs6e/Gx2HxPE6wFdHd3fUF1Qfi/racPDuQToPrpA2TRuRuLsm
lcaCXAGPOmQPgtywSic73DzxLhjrziULimhP+6VG6t3YsoVUae6nL5ysPzhF
O3tMqhxUHMPL+LBVUMD3gg93aRe3bTg2MR7epmY+EUyfZ04JOui2XkXJ4axv
GZTmfHzjnQKoxo+O/7DJ3ivy6EwCpa+Y8/y65hw8DdaBmso6koiygqSHiSy7
WmPqizueXsvDpqpkIXA58m/nH96SJiJn+vm7aMLk2GNJdaArR56gV+VerxYX
QPrrev60sOKRRD79aKfEmzDw5C+5vs9BBewettj0wR8LJ/KIeiB5M/btbaVF
+jR3/deWj+T4QbP9w5jgaN1fxG8XHoVPIaCsCeVzEJtIK9PvruTVqPJlUPzD
meWcyCx2+ByirTmiMHbubkfHufo2sSqVCiQJ8K7cabIMp8Gn0w9lQfQiicsM
eRuyMAco5AvN90LXcvqNQWN6wEtU5Tvjf1RT46sw0ru5eks2TpsQWMbKR/hA
EAQZ9Kz2BvQgHtbI+XN5RzqAXt+uYvWC6ONtMWv1IWBUcLJPRmwUrv03fIt6
JppXOT98nqeZK/qwHVOuU4xFbxJAVPDzvxWRu7vUtHyGZDHVG9C2IMYrwna5
6+bvGTZAhXiuCpZ+lhG/IBrChbxPZM0Es0thJEsk1oZuiHKzPxhjkVXquLTK
91b3S0h2/IM27YdAS9xiH9tsEvKES0fldf6AljZ9Gl0sB5Qmmizin1L76N5O
6DRJEzKf8dhnZKjnHEF7ZE/rKdrKUczBrki6XV7TOEDDdneML5r1Ix0RhRnc
pHwmiBsCmoX9dVzr3p7RsfF5QyBSk2LRZ5rrWcdcD6EZe/azs8Pyjvue8Jnr
qViP/sC8J7aM6Gb0PlmjOxW0gVMJuWP68WsFq78muW1ZHOjoC0Ha3maJxlbH
YMfqhbMOeHBxslmTABxWDJMx9YtczIFCEKToEPdgQE26twaDCFCkOu0mWGN9
bBaemMtlXk1lRzPcw5O0IWEFMNj/mwfiAkmbQ8Eske4Bpzl9fk6A/eMiBsbO
R5d5hQK48nRcXA2To2Vo2XZeae2SqMMpF0CgHYw+QcXuMO+mTvSpL7fP11vM
oNj9YDL/SsTkyj/vZeadvhaYAATtwEmJ9c/gffKxFolyz0ctxgtQtFbzU0WV
8fKnvzv9dW5lZOw/jB71gJSCpRqOEiTnj8DwiCpIz9Eajrj6gKM4RPrsUWkl
FjT88H9Wp1Qt4QFXhCZLi9BZ2rOcqEFe3IZ/t2HTPUyykHrLBByvQruFRpkK
1x1VyqWPtduGBo+NfQ37Ti+cQslW8UvSU14/RcqLnQ1bPPevL2Ize3MKMTi1
p6Q6LnnWNoaiRHSOSwjntRHxBStiFCAafOBCxX5gty8LvwLU4aWzZD3EC0wY
NZF4DuaZTCbNTLEdBeRzSaH9IdXBxygjlsaJHNiamtRcunWJvT1pQwGhf1PC
EXwQRjsut+hzbbp0bMf3XjqVYJBsR33ap2L9837c0UmNHntmZz5OxPoVil7d
2K32LAAi1JLb91ra0kSErTgHcGnavLywyWGM+3Ud2Eb9VfMeSdC1+ekxIJ2Z
QaINNVVcTUyLWPRBNY3ojCkS8o6iUw31wxc3KH2+2CjKDx98jVnQF/k/6s2Y
Lm+wLdIAo+7GbUy5pvYJOykXOYMaIrbQchi09dLEkQ8wXZRdlqkK0Mk5FITn
9VAEDph6wB24L54ATOz5YqnHLl28I8locQONxVfoKfeOqjf9krr5r5ny9d5b
LPH+PyXTom8cuSwY9WhlErY5wRvRTzlpRPbvutcwRe6o9Vq7MfQh3s9A2XoG
ykSnTr0vcZ5vQ5KV0R7zAzPIhEppBw6nuQlwb+FoGcGRrZODGuMuiZ5T0D4R
T5878sM9kxkRfxN4qV2PNnFaKTiIvkYIF/uZzaZfbIJ6/jZMuYSGgtqe13ak
OhkHOB8aGaauYA2u9yYCesJFrdLeac0BbTSeQQvUUVSseTCUV3ENiF9pwPFq
S0sBnUF+UTY5+LNNR2Se2qtd4lhGCWmE1iSZjMoiKROzSETzsKH9sO1zGuRz
BzU++IbmE4uUdQuVboROp2NdpngCIS0uPMt3tXcmNBNhdbnNgua2L8IzoceK
DnnmUrEo/UZQTBqhEkm4HHfv73JOlTQlhtWXHYV+VHhAW/MJoBX+R8C2bflZ
wDZV4Y72BA0q1vOefj9fVkw9SUuw0udpEUEvDxXxKtDOA5rxRqVC12JK4Wt2
EatY0XMPBByYssmu6P5MccJXaGUWD7B3XNsAJqIXOAzcrTAh+Bcvg0g/4Sii
eFJy8DOd3hZXnSXMUgoZiBieXUb8cacLtki7iiOy3VcEXdJOvV8mx0CpAyUb
jEEkJ/Gp6xNvAhsFNIbWt8P2qbtzbgScWU015RY5trVyioursiWcZ9Sf3uXw
EL4td7jrMRPCaa1chZp1g0pizjm6CPj1W0id2uYRA8TqJzVf1UHZDwhnYt1x
I4ygbow4m1YcloAaBwevWCAf220CUX6u30p3fE9K9cPPdBR4ammhCTSsDPfU
9wTAvLuMz85MeRuW7xY1mYfvHpdcJbOk5HIHxaZTsPrim47li/a9BIBckoAt
Fp7pSnk71CigiT7eLAKfn+1dOcCM+EGiUNqXGcKrF+Grdfj2EJImEkWiIIon
ppwleroSEj/KZf6N9oXRZKqJOEGgERQ1gBU12gom6v1byqriNcmICzHLl6tK
1NI5FMROTchNGohBDxq5ZLhi9DO+HeEpUIowncF2nrzyGvVwhPQHcO12n+OX
SaLl+0/ps+6uZ30rIilINyXH9EfL5IUuMoWVDE9ZLYlbITT0AM4uS0sc0mmJ
0QB/QXyKu0zJA+3vM7GrTyu8YozZR/w64lq8rSJRIJTGaVQCRHl90YIIP56Z
UimRznnog/cbdzJw5+H3v+s/EK6Xcr6zmpOqB41kXSDYiRFvrMaYGuLNelir
OECGYN/AE83C0n+43OW9gTopJ5oHHVILKDAde6wta/ZkcdbPe0Nm2voY9zVm
+b1TRy4LcokKPCnepJdaoZZxLXdBtzLF7ZlstbgjbTl6djaTuWKWyf4H13QD
iLS2RP948v1ZcRKiqQ9e6VjN/n0dJ+0E8TO8/Ik8B/2d/o3w8vjI59hXmaxU
tVtOz9CSLNB9QCw9Aii3ecJWYkJQaWdtes5NQTvfdHGSrbBagY+AXXwPQSxz
XtPVLhsnVGo4ZPKgNe3wwR/uuB+ZxkUPxxCwtzl2jIi5MglorIXPerzged8b
gUTqkXoqJZfpjqXC0tAVHiKm+/I45BCfwG+ZWrqMFhllcjqzeS0rIU1W+U/d
8O5KCnq6GcP/E1an/dpOZEpGCwe2qpz3k0a9GNnGmWCFiYQcyFnntR9zZgY1
evcxNuE3xE05pRnMlBAuyXgtLSEgAO7f1J3D3AecVe4TDrjMuDF6c+AkFTHv
heY2dRxjz+Nn5tOVDo8keKmAu31b8Klm8PTVXrwrS+yqBHG5d8PhFRgbaqnD
Lfy5QHB1atgudnLouBq+YboJZF/Q2r2T0kuXW6oQEliAz+IM55aYBWDdVH2z
swAhdxKZu75uHtcJKGjLA9n7YtvYkRr3IvLnfreYZz7/98gHDLmiq7D/X5ll
t7VzQywspJcKUE1tDOnKwZzYr8n/aiiVUlq3W8GSbGEmik3ff7VgsMo7uISz
Xlxoygx1+D3JPFUcU1ANDsxZuzDGEOI0RhqMW0AFFtzRttmCrNgj93zqbsOE
71N+XLdHjNXzMTbO5vWR44MY1O4UVZyoTYeTSHlNSJt47qQr1rV+jiIVjKjx
mkmvTJAlJB+46qig3knhzkjrKVL3nMKn51Z3WzUuQxh5IVi/h+ff6tgAbdMP
/rin4xpLFpUCxZ6PTKx4oFlx+ANvReuTd8yMCkDsEMwkDeTRl57nSCGeDznD
ypnApcdilx1N2q0Uszkplp4xEH9OiKP5SFaUt4oR808f6WuepHcwpTo9Ibyw
rNyp/+5+W/JSCUEjmJ6o+YaiL7KRp6V1QnqYOfjMzUou3jUouT4OGDArtN/Y
akqu7TqhJkii8RBonLLs5HoxPi2dmc1sCEIhcr7vwJmYbHJz8kmNSOx6Igzr
kQML2hJCsmYIf7OQ31qnhA2yrK5hKRPKx+ib/xoQkdBLAZtWl6MbD9bRUJ/Q
Ql5qzOdZkzq4kbqtT+gud9sRKI3Fcd65qYedtqac1/pEwNrcJ7zi7COzvAvi
w6jJZa2SEpWiXyWAxgheR3AFA1SCJAoP/gWhoD5kf5LJs8gFg3UCcjD1IvzS
Ke6nW3e2T7OssLsluw4iLHyaIBsye9MDHnilkklV7+P840xvoQMxGW5OcBFX
kZQQgC6ecQU8K531nL/1E4T28XT/krQpdRQG+SgyVUKlFc2bS5edW8G8mWzD
IkBG9UNG38+Ul30YrfOh1vFulkMIBQw/D+810DQR4Yfz40sJbAOX+IhSp1rQ
4ThKTk+/NsBWUE5q6DMzaW4N7z1s7dKjnVN1OASM7Bz2ImUaaoR7H14Kyb/f
FSq64OjE+PLgta9vbi1BDpnv91Yn+fDCsKOm1XcnBS0N0IzqpRr55cPhL/UE
lKhoMn0DayzWGJ88ih8BZvwjdqbDtBrgR7iboVBciZMj9W9m/Wbgf9I3VdZ2
sRrcENqKTFDYJYyuxOKDBq8JBfaEbeaKq9H7uGVzeb/eeFqI6xwliOTar2MS
fLhK5QQR12P6P7pD9qnHoD7l+tIpLj0Yqymb8CW6h9lDkrdV6fMuC8drZrY0
K2YF4WzaKqzNP6FVWqCKquas5RT+GC2WH/opnXM6vp50/m/c8f2lanWrhABs
3Whi3K1uQArTOIYrs7pGHywYrOlUoSvpIO/N1rtvx1wortML8ncnq10hMNLF
npIDhWZ1iygIQVbd1pbOEQKtafyzRorqzQQCTuGIwtQrErNgfk/MxzxDCam5
lzSdqmKWW+5GW8FKBIaFJaN1Gd0mLhRhIICqaPwRAOiPINxYENHiAvADuH81
3Up2vA3btZIoKRovw3onKLxiNe2Uwnt5dB6FnPq0bTVGmfhNgnyJA6NANYci
p2F05QkUBs8ZEe0xfk/IXeUjUxsXUNjVydBPyEjR7bMd5poNtBOJPyPuMejN
S5TRrKBDcaatGEUTn73eU5BepfsBxG/Lf6blLitvGyTBtvV3Uf8Ob0Su9yyH
TqyiNSqP3U1LTxK14mdGeKXiethehxaZ6CNPT3WnU92W12K5ULu18KUD9d3x
5MiCiZfFQOrviST9xw9q0N7oX1e8n7a7oqR3SLT4+x309k9Xe+xAk3cwqHOK
hF/TuNsUl152IT0jPCKkcOEGE77Nx3kmexY1UcvTmDnOJuhX0wEhVVMK+XhR
b13tuDRE8EB7tUnlOcJW3FZADlmHunIheRT9U51fAgWjf5nuZf9H+krKXDyv
ODFf+NTpKyRTDVgd8+rLWiMTXlUff09uDNK2wFLz+SmQ+hSZWR92WQLxNn9+
RHMFg+05cq4miaaoVK5/TQXrUoxx8vt6O/ht/dDlQgPcHBQhYzi5ltVXU0d7
kNu5x/4WMsEhygdFBkwqlfqNlsSlCelw2UypirGb1QGR+JeO6eW1GXC+yqGZ
jNVQXg+ck5gifjZnYTo4T51Jpf4mlLc1lX9f0KEf/vy1Xgd1c+d4Au/0xfpz
8WWCvjd4K0lkowavZAwWafge9C0iWngI139OdTdWP3bnxy766QoHRbNRCItN
x7y60IZLVvIGUwpT/AV4rP6o1kEadYXpTCdb6onweXa7G4ymbt5H1eZY43zZ
4tnJWHc3wevemROLI04UMEqYScsohh+3faEPLJp6MXpgC+FR0gooh+CBH7lF
fkqrnpRZaON1UjYJiU0C9nmKJ39Y9aagPKTLt9lDz54Dqfid+xuy1ten3hOm
9xuEaQ4llEGqqrLDP9+Y9Ib0HAyDMUCxQx6NXH3We55UQ42jFAqRsMrSDR+T
88vJdXabdUnyUJEx0P0uFLhLWQCdFs/m3fhvJlO37XkyxHOYHIH7IJU1fwaT
3Md7gtYIQeFkUgqeM5uZGCk+027hTB8tc/F8LqZYj+kjaCA1WNQwJNIxJLFl
Yd9GzjXGsG7U+rWmjhPxr7cMRVvnMPPU/Fk4pZWoYXlhHBKRU2JjIXfqlp7O
LiMdglqRTFZBMbeqyl5k+EPs27TobmsvKdm1opxika4lMeFqUpfpU8MBtfGV
eKM5bPcRWBbfUA5CUzLabtS5hLorm5rbsP4TibRLdx4WmoJ2rpOd2aMC969R
UZBSz/E6b8q3+HKTwDWgfcrLxphxrPVpucIBrnYdkEzZE2LxUiOsa7b8usO7
/Xmqnlh3im4jJhaiXrCYQ6vocCZrFPpirQ0JaNzGs5yxzil9u5R0IDNtm+9d
TP4TclRvAuxIVTbOl3bd1kyeqv4Pbh2GD3Snvn6NqX1mP44HL6Bzx++Lhmym
hCMeeLeJsmA5nzPvEzIgkLaOnh5wUyzTBgjlWp1DYEtQyR1MqBMMnrzl4kHi
2RSIZUXY6yAFMEgGlvRx1Yozl90CP9VSdmO3/AjrsFV8g7dzzS8AerDJxQLj
OkUuxhE17Lf704bdvVx+6jkg9f4sgm+WP2F7TCUQgM4LAKwGi89aJKzaSvI4
0tZv7gcfTufJBOuOHMkzUFNI+uWb2CrmREaQk3pa+vcuUsNm7falopVwIGGs
cuNyqOS7VhNHVCly4ViG/7gLQLF+bgvptWH0VNXLphPOxXwMgTUhpqn2vlHH
8V6Sa08bIfEz8LpRzK8fscipJ+EozHeINLXF2yJaUWf4D94rOIbllDdobGaq
8OKfGDKoM176c74r+zRbWcB+f64CPnwCHfcy6OAO9CYSxJt+bQGt7SpxV0Qo
l1T/muwWd8guEzEaJMMl6tBJT7xdxSgLp2aLjGj0mYh9yPAJbxs5EaAC2bSy
QzR0jo3O6LWMOIDeWn01IoX4rqAw74yl9TnYcvRjyRfNA7JND/epOICipvKl
9+TmImfERZItbJxFVhjBZ19KafBgU6khLgkUQhQn7vYs3WmAedG5l4TlWnN7
k8B3AeWDVTZS5pY2extiADfa0jFxRfL5cI9UqUHLX86hkONTYtdhJJEt7qrq
XBksRi+4Dg8Yfz58kQBNxmZf7G6WZquT5myBMX82nbDJbiRjw4MiVlqRdYhu
u2nCfYuEVngCsRH1W23ccPgh39JjeE7Wr/XFvsPrZovRwUPYKp3p8V1MJrSy
WMdZ6Qbfp7Bl+TxU1kV2m+8wz1oHr6n52dPmvJ9yAAJaeZ3LQqwFje6BI2B3
/VFzi7b7e4S4+FukdylMuV1zGiJPg/bIq95FfMA7SkBQsl9K6nOtk/VXuC02
A8Xl93oKNOEairpGmQ922GDF7qF89QSY6xoGw/YD0ki3h8Ba116Wh6xOXPg+
l4A2YP00Kt6gGOBrUO7pCdO+mguaKQvfjyo+lE0v/76W40jxWSr8kcw75UiW
1SxXMbD0NTY1Dn7ceHguFK+nEPj8CsxbzFbs0zC733jo53VRiYl1RME1Jnu6
REQ8xR0CW9uOcefBTrpGACQFaqnVTQ5FHUt1e2Xny0rvkZcOVNo8dHSHO+lW
X+yE6YYCLfFWZimW6dzVpKLcUhPbjCNR3FU1FO22vBABiCqM0mn55dPKVxj6
j83Xo7Kn2K6VLgm1ev9+MEwh0Ceu+9jdkCirQn5H9mVEDTm32lUYHF3Xjmtz
XSfmpvf2UeI6kuWIGdr70hPCFRLahURzek2Mr1TXmbzxTRLrI+2oMCu2uNZ/
VU9RCxb2K8fyORZdAkq4wSQct76Nj8KPy5pAXn2Qun6GORzoLVILFZm+C2nn
MQDQjdGKAP13EkblHYk7OM7wpWTTXFmxG+So9GwwWOXG4z68Wug5smYBkbVn
BcPOy87wRI5VXBAqhoD6UiSEZqCwqydkBP6Mjxm2W4/TRGuiWjvaeqmmF9ae
MeEqQ2g2T6g8Y3LYiehR2U+avDTu7SJ+zQr4WRm588QH2tJSzQYtRTgMtf23
sGDct6jD1sgt8cbCWuFFU1BKhtZ1+SSyIahvrxSOCNVO1X33YR9vy6vk/3nV
hQg4dwfFvxcfaImJaSMcaLtAek1+RlGf/kEWOO8tVjRCB4lqjOKHgAm0YnRq
kCRbAc3X8oYf6PsBuL9IDKy+wzbhbepDLlljgx2PaheJRqaqsQNbTGQuQ2zJ
UnDuoA5yU9sDNSR7raPz0K6laul5VpaS0Qmo4ptwpJOwbyjNIxJNe+vbDHjB
Bg+dbv2+0s3U0kTxWeuKLCSCirJwm28dVbK0aa53XVUObeeAsdU11Qzpqjyd
fwbAHy2eYTPUXZj0+GCClVIh8IMF2EKn9jwDPy+p3+NzZtH8U4Mq/7zL4wWt
YMAp0GYn+2qDVuh51ykKdPBjOWbTIPcOYJFDU9Cr6Rarxq84hwZiZAbOH2Sh
k0LwevgmfS54rSlegnebZ8lT6yb6p2km1WCyVbSOoXUsjKxMpYGrhc/D63OA
pGANxFNdrDpDtAcMG6plJsOueLBY3QjgpTm/wYcIfg8j7IyGLg6AccrMEf59
ifZfIbLYrA57iKlx11up8zo9uK3Lm4GptQxI9zuvkn2XZeTOWbFUDIvW2EWH
Q6CuQBFYgPxo+SROvXNqRm0yq9207idXjQHQxEo9ckstm4P4mD4CgLOhDrHC
76tEIGYgUcLE1oGcPnrqPerRCXUN3/GX23y7YYGgFv1Ga88IcMpNFgpwdUMR
mOfUZsq8Z7URNoUQ1kgOA+MW6AQ5hKW05qqJPyEnBwwn3gDYGmudIdPPYmDh
w1/racYooocABHsCAQaymFx2otCd8W8Lf3yKxIswrTmOLOlBoYsK8mEAePDg
xRqrgFw2qZpNQLPGVvXvWYxOq97W1i9cgi0abiV3FlMmgSi0vBDvpRXRU3fm
dJ9al97xGKA3UTarUQkya8eraBX01bkzsAyjAoH0DtMtIc8lUFsfmp3cL9+J
tjfyCD0LjkKA6UasCoNGwF0NnYfYJi2i6qhok+suzRBmJhvg2tMK2Ga7OYSf
3Y9is201JBnJf7QeTwOwL7ftNh3KSC5idyfoQjhFKdqRXPNQxWPO8YnVWRJM
rRTxUmSYUcfF9rM6+SWwr5lMtOXelvrkAJ/MWEKhvkjaaxJOWtvHScmDdsWf
u2NJg0DUhjy/0c8vHO0XRU0jeyjHB1MVMblSVmXslkcqQ9L787sGbI218kMR
gPd9zN1R2f0N1Zr0MlX+54GrB/NiBig5MfhkAmy3GtpmJ3DM3NJPtKvk1k6c
V+Ve5Mumlpb6V0iCU1SAPWmT/xzLoFKmJhJyXP4r7vatnbpRJBBxhJVd0nHF
UPhsvJz/5a+3tEUKDbIhDjqhRv65Ts9zyRUGNftZjtN9zOguXwvg1X0+CYhs
jDhSXPc1nbAeGbIl10TTuW28Apwydye7nwGCWTB0XyRgR61s9fb61RZ/bzGI
rSgkfM0fGP+YOFsBV/RRIQHSbfRbue4y3GtZ/4+ysKueQFrXI88qh1398n1a
eqiW0jd6ALgoGKS89OHeiHfmOL41QWmf0M3qfF7/0OJeMdHtsUy1cyt2rsFN
HPouMoZtZgNT/onLq9NR/lrjTcdEN3av2FfeOd40vj7IhQKAxwOMgzqU8kqe
6fjwTsEiNH5UChQS7JNk3vxYfEgkDPw3ZqahcyeG2Q2r2wfLHpyXUhsxVg/g
32wsnLFdQ6miIaVsyrRgIDR8I9Oqz216El4MjAgoP7dGnNVLQJrqPWJiRFrc
rFAmqOPW2gAKqYBhasAQC5EyevpkA7gqwjaePHDShYXReAdwtHhIy73Se/bg
fsJ2PPgj5hP4+meqKRBy0AEh93Sy2hUYZdEEVHiM3T8WeHrA1M8jq7LKFeLL
fZUoB/kIVXy/54QzmHawDTw007jrD3aXBXvl7lHaUFkCRexuG54rudGi2hCf
KNwm7zrFW1CpMWd/HHG98Zes4SKyZgq5xehxcj5PD0tlnwkbnZGClKfrpRmP
RWQb2awRY0NygrvJ+y1FbpbAeZLhwM1xXMGgfzF6RMgk+mIUELdSk1Rw5CKK
p0/U1Evjjav9kVDHxRT/B2qpyctcFUzAeTwS1kLlOq15qyNhAuFz+kg4bVVY
d5WptyM4MW+RwQ+DCqcU87P8yOhsKKvGDJw5I8KnvMvmNUFzlcVGevG2Edt+
0Ezp0Mj9tSxOI2rlNq09vSQfQa03hQlp8yRdQvXS4CmBIMXJyEo0r53hakNK
0PM0Es2Kx2LbijWM/b1xlz8mVCpT4UE6oFF83vBPYgaoZbX7h4uN3PsD/BvO
SQxWFX1EH/bbDo9pVdf8RolgvEeF1V5NHEuu7fxhnVhdjDdW6Fug1mp0zd2U
qWv/toe0fulQvqVt9yXq135ab3LCOintIcvB9kJgWIuhak9V05/uq9R6+4ui
mKq1ye6+syq2vXOXW+nwKvi9HspCFpBHNxrHgN8uRWQIVcMs4klYaWe/Ct9U
Z5FCXxRdc+NToiOdKyd3i/NNp+heyGRhxXPASyIdWryM+Guhqe9fRz3vO6kS
/XVZpucIpqczYVQ0jrqHHQGbMZaWZcbBPk2IQuJ9WhO9l/u5n6L54gQn5ioO
NPeg9L/H47ir8w9dHwsZ3oF1r2M+4/EahQ5g9jMCAWreKpF2zJzL+sK12i8y
V6LBeL665a80i6VIGWXcaVCFgBXMur/ZYKKWmLeW789X7T3TJiacZIiHzPf3
jFGN4mOuM8NGYQRY69LPbwq7HFeJphDKvYbtaMleIaMbI0Ly4+RPxpBug8Mp
GYCxUGkk3LdhOg+UYUiUT0zibj3T4MLGJxlX6+/1V4XRHFl3Twz5a72RSKWp
uMg67FK2bN8ZUBxU7KEHeCYNpYS9eTJAoGhPNKvVz0RH+bjmlqPS5AVZ53LU
NcCYw/1gwuDDr9CN2ZLlKR4m5td9xIHkMKrV1v4pLWjZT4IMZ633h5zxkvU8
MAvw/f9R4LUuJhLwO+bA7nvxfiQB5xWEVfzxhzrj5T9cPmnP+QUWEXFt1euz
tpbk4fSk7LrCyGLG8PZQD3XJFqVHhEAoDoRe77id1htwls9u2x7UavvxGgzO
Aw9TPghbsOs1t+wM+W6ltif6LFXoiAP246x/unS8UN651nwhaR3OBbZw9N39
fODiOkcb2IVixdbOHpqpAvIRKrFMbwAnxu4k5agjaYQTwCBMwyZHvXH2NB59
gf9dRdmBzoPhOiccn4KUJwuVGCDKWzv1wNwxOWzFOhU/G9HIHbJfDuM0cASI
0xNDxsJfGI3b2j5HIONgMiUTZ/OCgJYMLqdxRx9RE8lwIuaraflnkF2MFgIA
l3MCrB/LbYksZRsAAfieVEngLCnCa6lvm+FKduzuTz32gNu6w+nxBVoptjL1
osIXN6VIodFqqc3FaByP99wUUdDscZW5ib/ychWoesRrcl17Tzdhxf0FQ4wc
3NFmWlD2qHzLKnUGu0lmk8pxIQmfqOU9Kerp9ZtR4Ao8lMpGy4X69u/oNXbq
P49Bqtode1vZBeybsoYhTDWQZ8z/l9t6LlUvS9BoTgV0S/QOyb7wuJvJ7KzD
vqdBwqvB4sljrZ6ikFTTnSRoY4expiG/0z/X7YcgAhF2bQGysNtu8sIQCgUM
T348jq85ARGVxaoRMAYjNngcTtvpO7HgwO3ajfSMejSJzkDsajV4mTn96+9q
ON1Cl0EhDeyabEPHWpWESABhaXVdmtFu1irhjqYabLeLpMmo9zjB0BhopvsS
ARd7EcgKvHiG23rnFzyEi+mHRW47fFepcQrFI0A+L8AUmsQZk8NS/lKOyO3R
quUUzQYOkWrrrWNip3a+w8ImX1UV/U3xFyNwKyhnVs0WPB3F9dzd6cOatSwt
TQPvSDUTzIIU/1kfpKW1QxvSRGcJtV7Ssr/OrXn7qN0mW5+snsU9zAFNOyI6
93ogiICkczFvrTXFHLEVhiEW8YohZ2JktH2HqogXAQzBS4hA8WqS2JyKFCLI
QibEArtZwP7uV6bvK4Le5nV/ovcmoPZzm+WiEb/HpJ55OBgxve+OxRXwyH7v
6EeuwTz2faKLNL0EfZ4AVhL8brfOHfwOMm8HN+JpOCwyKFFz0xDkGp4d66TC
v3ZWTujlrGsYBUWq4hESSXXPBqn3RvAhxS6S8/bw+s7GvTZVIGMRkIVyttrT
782ZwSlRp/89LU8Qe9PYkhbC+kJdpd9TdV2YUx0+2LtA+bGtsD76yiu9+1eO
8v8vs9qJzd9KxKFS9ZOpk5HmrYMxA2Hg1vfk7ePT/18vvpHmK68bgdVBArt9
RG+aePgajQ+IuF2HkbFnMFYgypki219j8NeENjs+JIs+vkIR8xfns1IN9Mp/
tbYB6gzNpYSzqLocPS/7vHvqzLN4BSgySd41eEkWknlDgBEgFRxCfef+JBgz
UpkZucmRNKciK2SwYtV/mfuNmiAqVH0vms1ihKDDdCWieV8B3MK6l3fntpKh
eRlBALLIelaNcAuJXUHqhAfKllQPTSbikJzNaPY15+fN8sXWfiCQu/AN6nRX
FRWpLFDw12snw5UKw42/PvToPZDzrsEm0gQbyRITJRGMKbbSJZ7mlPMaSh3a
i1rf6LMwO+15MU7A9r/WVDEfvj6fowGKyMdmITtHVGR1rc62XQuk1MJjy0tD
E4u3khyhMwKUOiyGK8OMgDiGCn2JgE+LB544rlmxMfQiFgEyrck3Neevm5yf
MzFy8jUw1HH7fa97A9IaOQXx/7Wjs5G4kODkG7qD9+AlztEyyPgkx8rtA+wg
dusBHtFQC2dmV6xOa91vEPGj1b3pD3MSiDrHn6h3qgIvworZLYAusSaDLb+y
Qc1TaNOFJxhUMMyvJqlaePenw1xxiYzlHE+NKNxbCVOnjWzQxgfuHtRQuSI+
zfuKcsCr8XfafgY2RCJjHeOx48cc645TVzbBmM6la151xewDYKei1xHla+Rm
cnrEFcl/5Mv6tHDnwE7VPu08I10PNbIUOrk5SpSMb/PBbxpcUScFkRyEsJOb
eT/bRQjVrOQ2O29IEMMvYb8GT6Go3bONnu3N7sXud3O+j+LvSpWEMKjTcEbR
PpQh9yvxAJvQiZIjE3y/BK1DrBtFZ5jwsyVVRUjR1ygSJec3HnYWIJqwxQt+
UBB6vpTjAqu5KVES3D/vhnX2xzcb0H9Dd8Xhxh+xrm7zS6b28juQ4e4NSWVE
RIzCjP4+sAooPpXpetqksXGwQuQOz9OYXFcBilW+kxVj7F4IuCdGNB8EmQho
8RNQ1WGmjTVbIyupL4GcTPqYDo7EM45JGGtJ9QqH0DBpO70K/W5/VhVoHEh+
9OPfzDMX7s0suVYphp74b8jASVveFQVe+YaEszDKcUsFKqEHvnCBJSGuQLtv
WUhfMuNae5xhy1Mm8vyx6h3gs/kK9cs9noNNnblG5fs1nAqDpthEHpVeNMHP
hJSks4PS1mxDO7D3K5AZskt16+EMM+K0XXpXw9ySO2cVzTaYfHxOJfBapYz+
8N7zrQJgDg+5iikwqwZN8D6ynRf4kxAk2rpGH/gghWylX0Hb3iEV6Bwvxw1V
j6WqwBercBpb+euyhRMJ6UsU8epqcDHhZExFKXXpSGr0QgxstMhaKI6JXDCR
so2w4wdJK50dri6cjRVY2COesoKpcoYoa3OVWaO7qut+IhdxVZwvPMzQu9DF
G8yPjN+/Ro+Vvv7slB4/rlOjrfS/g+pq6BmbAFM3Noi8FOh8fINnRSosMwX1
Qb2bS+m0lm32OOhpLzP/SBUWN1Zb99ey2iopzIvfEl+20uP2J2FFLhzysx9A
n0tzMVgVgmm2NXuMxGz7vp9QzjHxsL1Uvg104dFZoU3ShynbhVl0Iez2hOvT
vSNZHp7zpelSR2v922b2xbHXRgnlFL6EExWBiyw8rfmeGVqoGcM1HH4OZEeG
jrRHCGkuGqG2FF1HyNqIR4/Kqy+QePpC1+ZxudiCH/YQD/Uj1eKs3mdH7pOw
xOlb3XCMl3Oo2+pXcGvUZ56Ig4KfgzaSKw+lbz67BPh1DawDUDXGu5kl9wNt
Fyvca3n6gHmQ8u6gTKIkKEFavmn6CuQHZUHFqvlH3DQy4+qEAkt/5nH5fnmv
u7E+kGNb1yxRDbr+Nx49W+CtkjUPV/aiN6ng+RYrfs8Zys71/GeUXJGBaZY1
hjccuaubFHgDOyhs77hDTnZMzPafRJ+DDdCb/S700gaYuokzxfOcZpfn08Xx
Trt4V1393M62IVAPnAfVRGTjUGVgZWmhBscXjL45PYARWTxY3GXhfP0kar9b
hK5T6spQPJoCkp2d260NhlZdOV2zB45Yaw4Y6p2vx9MQvlx71aFwOJxVyTKY
dvMIWRFfent+k1a3WZRFNWNdbCsNy75yJ46NeDeN+8kAqLAxthBDSYDnMwUC
1z/F4RcYQv9yUwYTmCBNNB+rh9/u68hPAboat6H9YRMAUZE+yK/RWbGj0Ykz
smrDVHqjZjkkqsffZBdROairQUKyVwFe5ihx7nHNSJsiX7hwBfR6KGSMGD7q
8BFkuhaomJdo8Q5d+X7wqIBY3YCenlWmXuFgQaIBhTGNRY8RCz6cq43ZO/rL
UVR/XvnAdbLJKCzp1CnZHOn7IMD5bMatXWYWYmiIIYdxSG1xMDmiDSae/EbM
P2sZbOqU7bfx9g4+9JjLl+LvFRonlsxt640wvUbYnVlvMizAahBPyCS8THEi
2C3cLH3KWBH8bVh9Bd6c7UW+J2A0m1PZ2FNR+xuDPJtGKpHfg1JiMQ0Ky+XZ
AOq66PEJfqAmg0ftF29kikZiX7XWGaJXaEePnnG6kB6lKyx3LLwhz3hMpX1D
RW4eKfvgroaMCCTvfvb4pCcyXLpPUJw1/4Droa2u8QyBbqf1tex+y7PGTk7D
Qr4UiSogeXQYxvrL8AtoKzMfX1vaT5naS/FAYgMJIJWM3dza9HbopXIj3Xtb
8hPt6G2Pe2PScfcJWvYoZ+BwzjXmqRizIAmbnXgZJ/PMY7oEgW0a/KWzIdMG
XeeI9Y0OlGhvqZK8ZVYIyeHVSXg+Lc1leONNOA1qwA+05tWN/FD92Q5V7RzM
xL64IVGer+4PPV4VEUQCQ8OEWO3Usp+zpiaKX/0++BA/+Moog2ykeV58kf8C
MIjVS+FKDiB2n2MD56zcHAHOWk2atG3DsgIpcMJTILdhG9IQNGAsz2xMPbAv
PjDvyd4jSM8cb/t6+/a3zefC/GoeeSBq0oN4b4zZWECJyHvo7dWqM68rl68w
msprkHwPedR2aIDG/YpVs1Jm3EdDVi5cpCdKPsPcUWyGlxamz2JAe4f4T/cE
KnQeYAM8+m6/jhMKnfTKeFsdjr9GoSIJjMpgO5RMC2789oW+49K5wFy028Dp
ArLjRfROnppc76GZsGiIuv5fTqwZQWCopkGtJfcNf1luWU+eHJImvJQjBj6b
Ii2Lr2EDh41MuxKYV6UUKaEDs/KTycSRLsbCQFVmo87w3VVVnzWAKNixfepS
ncOIf0Kob0w1V4PnUqAYTaLrXdR+p1vboZAkTXtYzGhZWfdcDIhkxxttA37k
dFo8ybrc+aO+9L9NkEybu7X8HB4gZOKWdtYyi8gF7KFHg4+Z+vBOwaT/7JDG
j+fYpd6VknjXNpmMklcALHoXVyVVklEdjbpuOXtVquNz8nIL7JrUP+pW7c6O
JlKZrx5M/nwg3m3jORZ73DLdDK54XS4xjxWNDmELYXsMmRYkhfJeqai+/IBp
tGcnDYW3jrFcgx9a0MvOtGTt/Nnp7OuAsXNSCEvG+cztRcn4e9UfCjJZ/ebe
VQVmymZ7LOyX5+NjtMpWwgZCWD7b+Yazsdb7fPYTSQ5jC/vTHNqBRdG2ds1O
DGNmksqm9e5xZZoDShFIfDCx/9Ntqfr++lLEcfCX/6mNF1vOTmNgy75LtVmq
YyGdOre/G191KdTxxDd7ojf7dOv36ioVKntnqtMC2r+ml2IetrpkuqjU1f3y
3ixF9wDyekNT6nOw9uiDbV2GcIn2BKYwOrB20+NzGYAA9DRswMK8Amv25WKF
STIcuDIR+rB/JhIH6jfC+UmlmE2PhKE+C/Wy1UJz8SNDZjcyu/xoMI9LlC32
WD6670kbXuLCuNXKSpwt4SE/RHn+2A0hBE3XSIh85uKVRAxbt9P2faDDAUhY
REajwzPVsGX01XVA2W2qN6K306WkqlMS58R3P6xE/Dh578lLBcsLlyWdQ2od
nDNsoydgeZ2uYI64yRYT3RZcfxvnh0RqxA5wUhOBE/ATCKwFCHymk0tMgsvM
L666JWw583qmVTXhQ8E78DUEE8HPmaaOz34aVlByNCPank9un1GEt6KTUCYq
p4EsHzyaEqItZAjHMDOMmbcxp2h3VuulqA5Nyn+aflMPFDKcd5ZCRRgqutqI
4afLwdPDzubMmR8fQJUmtjQy0/nzhxK/2oRzjJD3Vx98+NO1VjBpLg6lmfTd
8eOvYlhEUvAer3PZYcWixU9qXyHfGeh5v7Wi8pfKxJrTcWUiSaV6SeAzhUkV
LADcljtnTR8EF3AZnludJ+mywYhvms7CaJdwdP+8VLmbu/qYSVKRQISsQWFu
8Crum6FiuKdJ9GOioihK04BHFoFDIlbiUZ9tazCK0+XMABX88XdpP9pFsRo+
uyndad1eX7iFReQzAs//oea44ZVmJnJAljkzI+Ly8ar6PaRVTek8DJ/MY03f
QkHtE0cdI4t6cTeCC4zYoCR1zTuoyLnV5vOags+YxsWsXFFcy6c4bPTI3hcQ
hJshuG3iQRc+5UwugSkjReBFS4W4CXLlTZf3CMsSJCAoAu4Vw6Cxv+XDNdTM
wGxWCu3WYQBxadT2NU+syp+gCqXYxA2Nqqa17cArZgfhmyePRR9GP7Uw2z1a
rZG0wYpm0SWSkEfANMd7MIerp/XY/Cp29PebikHW4665mHKTrVnIY3Gt/fCq
5Aph61pSEPUp0WyptYtIrgJeyUhNs+j7EP12CdLSh8k+JkV5+mP9fVuYOjWN
vxG002r1aAp14ENBC8WjCxvhq7cb3UY+0M6lLL2DXUCe8Qur79KLrOeqZYdy
ntU6635EWcl7Ydb2X5FCAArRcPy1byQW6GW/0nHLZ/Bhz3mtaCZl5MNvDc12
c82HuDjSMiTDLUsDECCCOToQhklGAHhWfBsDLv8D8qM33lIYvuTUuRQz2TVf
9QH6YHrVaPnFr2KeOhhtJB9fG2p99ksoxt07UGuSU71O21zAIB4fjGatALTz
v9rFZfHtDQpCAI3wXZRzfC2gwKrOyusNmxwv/2GKH41dKsLce5jwFaQhKWtd
6y0J0iLDqt86xADE+mis/Y3nFC7zT2/sn1x5A5TQOKOOh7697Tx1jRvbTFC5
43wFbXb0mfSuRr1RdLFcI7W6eQvaAyOZ1koTMguo8xn1nTbL4Kzi1V4xVVWe
88cnJsp31pX1XqlUJO7NiWnHDxPqJxcvQz6KztTtWFAuq+1A7o1I0dOKM+69
y72vGa25NOpZUr13kRiNTqaHe5H+ajvQ3gUq6TmYIVr3jSbohDZlI7wnmsYS
fixfiYtYOK41qfFkAICn7p8ZzPyyTDLLYQoAuqMB0p79XpzzlYC6Jsi3kM4f
nYbmhAIbJ+34VprFsdJwG2rKoRUQN065b9oCb8z0lTHvyF5mQf4M7tfcMOBq
6Ma2X5jOS92QxZS8HAb0fjtbyVx5J9Cn6dQ3DyklxBHTUKc75SFEXei/tRJ3
mjHqhT5MJE+PQhwvnlgZLeo9aPF2SrSRtCY6MFSRetCuJY5Oelhmrkc/2bKL
SAWp9Qh7aNepRhLn7CgKlLB+VUGojvRCZh4Aidfco5Ci0VwUDP3ShKZKBbxJ
wgngVgrNUVAHLl2e5zhHJQWxVRnSdL0Z3l6rJzTx7Up27NxRAPjQsoJ6h3VQ
B7tkDVPneU2QTxIaSViWpkXczxsSGVMNMM6F9joSNkAQQ8hL0m1MY3k5vsck
8VUq/cZ9QymXoHlL+TcLHFSeuLkCSA8jUG5C1BrV8q9qXpiYLgf43VQC6Rfz
eg/rfV0plTeKBjJW+oms+AfjIUrmBib+wq4nS64OYS/R4NgrnAsG6WaYjsUX
sKeHIqxKnPpBovMiqPu40ngk/SI9Bsmw2G+2LE/iMbbTuF8QcxX4U4x573dx
4oVqaNyk4bybw84mJbk9nxx8ITT2RNLb3XVn4mbJRph69kNU9FeofMaPBYKk
2ve4p+0mZ1IoERQISpMK/nSQpsAr1oFytQxkJwaPviDWmDvhdrGhkN9JM1EV
rrSaQwhE9KiooldCjZdcklHBX6AlxvIJuV5DM6WL6tDfmSHS0iVM0qRn+nLn
J9eHkyQiMeGXTWyrOWA+jnlCDivQItfNSrzNPkZ2jTxnmkUykHV23Re+4CEE
CjMvDLP6YSbhWIM31lC5C6c+zMDpxtrTDpRSWxcv7Z9u5HOXPXs6O3kfo2vr
K4ZK5MdQOCw6svI/reLt2HcCaZEtYeura2A6yLnHtBW0hj4BWSxNarChOd0r
STxKRtg5BhgbqCFEv8I/xGDCXq+6XGEjgDLP/Sg0OdGWh5FsewcbuA3vQkLS
TS+7qHdV1/ZKIR3t3xnEhs11W++KhM83GtTSHbC6Y3eDmr8bsS1QiJkTlCje
/Kuzu5fPY14s1Ojsh9uzmYmv9kH7aPGoyyleXRt6WHfaXlfIplGLCcPsPcOV
AW4o5ouDBSQPmOGC/KjEBkMl6Rm/8rBNsLu05EcvuyjWPTlKeqIOahGIqAcO
A98/C1zUEpfCwd5chUsiDpkT+WBTwXZc0xPwKiwKsDhz3JWPEIItJFCE4l6x
Dr3AgJGl60Wf5Cnf4VT08ayC+QtQb0AYXy16moBz4CeoFY1qHcyecslfMnSx
wFn/6ExGLn6Mi67/WRP5INR0ngdLN5k2T4AcrMvikotH5iPX/KMT9DNa56c4
eWBk5Nvl2b5xHHO3Levv98zI/JZkew3Wq1M8+qJkastUsNWtJzwZGAG7Fzjx
Bxj9KtazmD4OXCOy0VAHJKabEW7NaXb0KJXTpoq3rAZqU0npNzfaj/97UchN
gSblkj2nPsNVbq53V95Ls1thXOf0RNGscwma7y2ysLsahJ+mdIQol7BBzCMc
8KzuQQTOLfnyATvv8U+KzskkBFG+nC7A/hSgoKtcOoyBPPKfPI+Lc0ZdMNgt
EdzZRHc26WIqI21pSnwF6bB1ziqLmwfMhfgRndaiRLxTePjtET7LSS0fEDbg
shSZ9hYGRUQ0MUyY1D34dX3gOJQID9nfllOIGHWADJA2pZP4ctmatxLNAN+q
oSpc07GN70/tvGgsFUmLDBUawFhiZV/jZxDQwu8cYTjYVQvMZL/srqFbO1yi
wcB/cnhOMpVqBcTuEy/bmOIeNSkx/imxK0uPg7G8ASDomBeAnbPGdp9+21iK
8u56u3xX/hS0WWoJ19eeOutXimXQjzSNBi9nXQ6zhVGU4AAQv+Q0KWV/I4Vx
Plr/a1aoLtlc/kSxAEN0jQkhyZ4BkwiT/vXQ+WwOOocGnumewwTuFDsajrw+
MQ9zap0ofrgYrtuig/bB9KEpUotE2mJRL71QTmZrQ6//9SPsm15Vk8JtO9QA
dX3HpcLZBdxIajdX5EhTPkTKP7AuT4i9MtoY/NRuSqHJd5nhBcG2V8OZJUF4
zlW4q8J+cF/cgwHP0f/phfxYLYn/eAKdeeDsUyCs2s99xbRwPtAitWuzgeV0
8gT2hRuupCiTSVmckOi1FdTO+bBYKBCiiW+WtRjaKqkdrY3pw+cFfMY45MIn
ne8mAr9JgZxV1DGcz5W32c4wojbIQ4W/9B9wdAdecSWlg5rcebEjPY2Uyv4Z
3ZAk2yZr/cEW2GUkLNjKme3nFg4EaFqk/ZKpYXJ+mrj+hW/MFzpZEcoPX3Q8
8A/KZ/TywBBrDkZK6U+wRvWR5HKqDRy1KjZvTjAEbWyxLXxEq96TGlzqe5h/
OnSKfvg5nuHgK3NnOnn1WR6AlKi6Ntt9bOZu09/gVipQW84wHla73KgCwRlY
O41giga58HfhIq3SMvETz6wTtgD4X5ApG8WPKj6alMLT9mCeATUalHHfLvfH
3IlVuAUPAbH79uU1Yel1xMv9xkHaaIMC53AarlWAB1Gz2vmnISIqB5pQa/SJ
AJMCkkhPw/3fkdEMNAfteEXg/GjDPec+V/OEC72b3ATAEdwk/aUKBeTCGRbV
0kcfMDVSF5bxKssPmSeb0FJKmM/mUQ3B9GC3zfSHxRxmEnDpTDvnECEHl8Fv
MuHAWzTnqhbDikiSNEeR2QnbXRn5quymaA6CSJvzmyKkcr55Qswe0t9oPJW4
RjaRISA3KjGsDFU66ZLNgBxXvbyFV7hFZy7pOT9FyGmXCF1qNnxjR1zz4rez
FbxfEGe4KWk+zy/6HPd/kwovesxYVxxSUjjNU2EdCq5luovexvqVcGbugOnJ
Cd44RORW4E5CWEkHQFwoUR38MN30diBJjs/Ai5GFuxkXMe7NFj+FTXorStMr
RDyfPSyja7sWxLtqkkad+2GUUec9xbs3tEWUiom8T2IWrQ/MNVIKivD22OrH
kdYM1dadeuDZcUv/epXNDlFizzmyeAHIoT/9+/hd68C7h4fW10a6NxBPuVY6
c3ZllosV73BWuZpKKbkfqdpddt+3ufiusNU56geIOB2GZ3OA9jMAlhACMSrV
Vv5Ee5OJuizLfNhmcFVH/jS+SGuLm8cLYmOUIJjVKy1yFiYyW3/Hlk3EutHg
Er3unDUXUbLnrt2GX0QSxVnHdz3rdS3JAQLLdHJRVy3yztSx4Alu9eWz9coy
nUD8gNLtmuuqmHvmNauVp66v3xNm6MUC7R/c/0m6drPeRnht2OXyrIRxPRLw
/BR9wPMEQkCZf0Tf14gsfVA1WBbfjrnlDmSf1lwYhcSn7z4vd7T8EF8RMpXf
xmvfWpCjVk9W1WfZ14l7GhFuh+ya2GmfACQg7iM5RV8Rft5CG2m8ZXtfuufG
8w4sYKX+BWKZPyI7GXzHJ88cdyi2bVCpv+JQvUHsSgg+pviWA1l6SyyL9v2j
rng0ry2UZ3IyDyxPkISAfKtpr3qQhAXsvI/S0GmDx3Oji3tv+b/YWrNP006a
CE66YzDtTbjpDUK6WdogFDRTq83xhH04ZZTi97LAx0QjxLOPygRZ9EDHRjei
wjVOHe14vVAcX9irYGHzSnGzys93aF2ZFjTuh8SqbilNfU7lxSsUV+VdOy1x
S6HFJIArMtkb73USDV57nqowo9MrXfbAHOEDsy1IOFs3sV01N5vU+ioe2tWK
Zpq4YkMQriEKcjAmTrd47VsHRsve9XL9qnCE+sZFcgq9fewFbFtendNUhfz9
MBSbkM/XCmGwjpswVClqehoDXHtJjv7NiUXC3vebiAwNWLekOb5G6u+BXk13
9B+whgxx3eDwtN0KzBeCiOph7OmqVYEeRbtX7f10dWFvGWqdesEKlsZlcj2M
Qk7gmss6K0CsC/dj7uzLUWSpZhX3rBxc2IGWqOqO6VoQyTHHtNy8y1s/C+uq
XlPR5CQjgh13z4BB5LoczmfieF5YO+QKlCQtUp/y9NxI+dJ3FnHGS/HnesVM
XF5VIHk5hDIXmShbNb4eCs0Efc5lQDzm8sNx2NfPzPG7F5sVGgPgYpbWTNhj
CpwfjxT5go93e+jAnQVyjhslB5CDBVpnO9g0bPGvLs5DTOl88adyFBgfE2gn
VmuTBVJ9Huw1AZYZ62pyMAwj0fW9SRYTtUP6rE4feqw2tiljgKSTX3zFTHAW
gG8mKYT654smQLXqCFKKF2vluovVwGnCOcvs1Xlkjqg+ujfPWGCgXT6OUpPb
PdMIoTfzqFUp5jHCi+85pi18C6J32jxwK0EynCRnQMeGbqC1+gKlCjEKEou7
/CVAsaZhGvqXGfKIqMsg+5QA8dLm2UgO9WJR/GivNPeeOIri7ewMB+r1QNid
eHnwgG1C/lGkrpglR5ciUTNQRJHus/4SF8AtsMKpkLzUcw55/n/Gqd6anu41
vQy3PXjZRWakRf9rUEAc4IbeRy3JJlrNsvcqQG4SYHVkR/3kv6p9MHOTV3eN
TuQGlZLOjY3eFXCXN7f9Len/nBFPqR1PDKdWZpnR0+E7z6aYbDi8aswCmrAJ
gJhv6QtOf3eDw08xNT45sCzZ78r/KKbKAsIvGLOZX6sjNpojTgOpjtTth18r
hBE/pOAObb5xYcR+lIpCst4fe8oVyv2SPMNaG7BIEF+nd75ua8WGAfOBZ+v5
i50zxtvLJTS/9dgTbYacF8SOM14RDx8QL8gagNSScK4YQlUTX6wZsH/6zEPK
rfL/VaJubEu/xjOtGF3jwj8D0GobEvA9kXblQcTQvOJsk56E+l7WxtrmlDzl
kJCMAOGgZQ/wfaY/ESB251HKvfBCv/p7Nq2FQ6HcGmFvMXevwkb38t99LYX9
Ecgqm2XxsRWIah9R8UW2rgG/nRc1iEXCMspwvutlPUGwSPUlYLpgesN5urU2
3XjD8dH/CLwke/b37mg0qE91n+RrqoU/0Cnar9Kh75aZRjzR8/5HqHd4W+vA
eeUQ14o9gy20vhgEZyT6kMVJokx6bcXpsgyk3xqPSr+1yxpafhk3NxSYl7mp
DCcnN4qrBBQ5u4SPDuAM3NwxDsUW1CMdCJAdbGT5q/7yhrIC6buihxQBh6JC
Nzkfd/7pwQk+87Yxy/N/ViLV2ZcFVK5DVbDauFDKejIHlyflAlwfCg49EVa/
29rCX1MTZX8+5vIXiGtppWUrkbS7HBV4vFyBZkWvM0Q1yHgHza08sp+qi4ZN
IHbxDVrvQMks1YXnmmh4EF8t8H8SYLqZ1tJx4PSX1tkh5lElIPZPn+Sj5bQN
hqZYeqTI/f92+PbU5KbJ3fpw+kkKJGHXAlD2JvX730zJAzPjuiYaDZELHRhC
0nBZ3dQK8GKSiwVztdhh/ocAwHhDxNI5+jsnk0b2hDKzk8u9LLDCe94RLFzE
034iAtLP/AGEOJsjZRynUv8ltMHewqf/aXkg+Osq5VKRkvSQ95/OsZLcTEU/
VHTEaQNQ3r6RSas/1Ur3hI6sIUwj4AuPmNuB/DTvUt+VOcqXvRijEvjlx2bU
XBUyvc75ldi8b2DXGqwhRRZ2YcOg7VOQtwOk7Kgs6xYCTWDlD9/Klx9bS1H/
5IQUiV5hPm18NUFc/YSWfIOy08XFq8H0+WaDrCpDqv3nsOfgy5j1s0zeMzt5
D9FGcRVnYvUCRvBWpuDwQ6Yr7tn+LGC1c5LdLjh08PirY1wbs8FCNMlb6ElI
kGRWAnVN2O3vcf5dvzvPO19FpYhK2CkJatJh36q/tDyHcNSNw239cZVUl/xa
BRe7juUjD0tOSMaTDB3M8nj7sRzCTwS1M3alB22UqyMHd0KybSb+yRZOWQia
xgHu7TeH/u0E66sfyF6deb2R9S4I54PENsScZH9FUThoEON0wMSmHYGFIp1X
d26237XaNguB/cxgRqMWfphcSFVo51NKmRUGt6mstZdDOXE1gL7fIZBizpFI
Nh8Egqp6L8IQcW/VIG0sKfR7aQEgHQaxFqYFxqG/WllKjuYq8B3eyDemgv9K
ZDlYK7AUYfnwBBHDPl6yO1zBDr6GBrlysbjzqpR4xjwCWLtqemE7boGgmMXT
GjYDyheI0JNGzi3DRpaQyHoIntbSOaq8atqXPlXakQGBv8L+6vVWS/OcD/mH
887eOCceCFDca78rQr12kPUYzg4KnQ06r530xrHQWTQk2gL2xFbpJsZ8qQsm
QETlqOOTWnsMPjxLcn38z0bkvl4FcqfaqY4ZIy1N6gPZCoWcU1EUAcnYjC8t
18uR/h4NLRvlm+edt/0OzX6UQBlW6mHw28Cnklb/m7ezb2voPJGk6vO5tPqW
/FX7fniL/1FNkItafleKdyE3WNT7bOQHz0y2jThnB+HNDBuTkzSSnYpGUUsx
iZ3OcOFyP2HgOamR4VyHxcXYWZQZMYOMfa1AEdgGkckz8jhLnFgtXk4FnSV8
sM2jHgnpdOrff+QDxEt65hthUrx8u/oiqehZnc10qBU2JgvdFPaT3sroAS7/
gVVL008Lz86BJf8YTj/VWsK+l+jO+S/RnnRJy20rHUuPpwOvaO2urzImSTzT
GeI4FeRJNks3zO6ql9xWOgU5N+q4zP/+MA6NweNPngoqzfGqkw5D1ePFk5Rm
rSR/mSL1IkoXzliQhSATbGhunFqsXCFwnaGUNFuNrt0vJuO3MEs5NnqNBi5M
hp/Ar8a2fCUZpZY0XYXASM5FBRV9DpKxanaVRhWmP88SLG1Hx5ty8Ths1/Gr
o3C12A+e4Ji+6RFH6cyjASNQGT1aaPlWuK4QEbsekGY9WnR/PkIuHoketC/y
w2rPJ3TJGzaKyHleTJ1zl+nmhir7Z0t33RS0ijhDNC3TT7OZi3w9ptoP5ccp
UCjz8hfFxOGw8NVmptjl5i/S3whze9jXTbtlG1GDeuz4hQGc8NMtONlmYNnp
LbP06Kc4Hr8wuGQcl8sFAzjXnTDAKEH8k5qBD0QBr2BINZ8O4shKWT6I5m0Z
fzQCaZIuJJ2pOGg2czd6ogofyP3AM/1sorwXv29WsrH/VXNdW4Z4W8hkkwdv
iBnQ5FMCO8ds9nZG/WcjNszyVkFXTNUL1LXj//5CjnALDViJCGkksMznvpc/
u8ZkFc9yTrlUrUi4YevirgpgQ9LStySvSyKtjl+tcS0PYdrMV7UBybT25hoP
lr1oL2iqyvwZ3S7zZaK3nbZegYySzRYhLfpY4a31vHibFK5HOSZoukU8T6sn
bcMDUAqgv0hhaQUVSh58hXivigHU4FMzEdiZa4+x6079aizQW41fIt192WUF
6iSmYoPg3vxIMOj+yJoJ0FF1zDdVqEbfJ8tVDoi4Nsg45n0SnLzAR/7bhwCo
FnnydSMW9JW7rfO4CoFisbdpWm/mKppciKhyogQyMxi/+3WjvcuF2DHF13Pq
/+XJZv/XB5IeFX+FjgN/HYO361tQGqrgkCKLAHbUmijijC+DNZ0+PTN95owa
9NTFDzdOERPZ4qt8SQY3ajb7i4hk7b1lquGglgxjbWN1jvZeX+dNowMUSM1Z
kDJ7EX7ZhduR8jtgpGP0USuujLNxWK6m43bYN7IHrNlJ/g6paT67qT4ePcLH
oP5GUzh4JYsKEsfftE+MYcCxf67+48R2Fs64XPfvhV7xWqbOz3hdkecDJAWV
wDezIM+tCVeYu3mOdGH9M3c2hvLbuTeERtqXHqLeum1TjobJ3lyKC9aw1qVB
X9zw71eIqc9zuyeoMzwu8VXs8+E+3qXexg837wsn2nS492FBWHaGXpNo7kxE
XPyGt7TGe3/LAPmwUODwri7sxRmaK9RL0/dGNchMxghe9b5UDhE3+R/woZSG
jyV3SFDlNZ3Q9qQ0JHeHSByrve85dVKfJ4bgKmE8xXgoVLF5i7PgLcmBG3tn
spLU9xyAdQLqPRPKb3t6veXNo+Hoyunntvz8I+0jlHm9frX8k6m6L4LBC0KL
1DWWY8LhvVvJoe3j+RYM46jpk9FCy2bxLsJttzCQFKI3jG62lQD+sspwjvk7
8AMqqRM8kYwJTOHHdslN2sOlVR1NDpDjtCJHmo+T9sfkzMo+sjoBcbxeZ1uQ
54S9d8g4464T45txryD4K8uz40yhZaj60WZyavD4DU+EQDPfCF0JRX77aGvz
8i9SiA7rN/guqG6RGEBkMZvbaL1fnQFwrFWMuhTeDjIq9ySl1haqY/dbcuiq
4NxhC7RKlZErnUCTcCEqqsCgkACEt6XY6UVP8Qp0+/1SNaNaCsNTSqFsTGq3
wq+v579jxzMbHfFSGog4J1Or83O6tuXwsGsSBY92cQ7IXUSKBqJuESS0sowR
VX+nen+cef6ugzqeGJQ1JZnsTNxHd1sPlieribNF0idEngvPNsi7HgbP5508
GsSsK4uD4scF9m9xs5TToga0Xk63E6mIzPtBa46Hza2nxZEH6VZoZIqRqSs9
2GEdo57YlGshzUCQUheb5OuCNrF5J6KsWYrGg+O4FFdEmi+B6FKkZuCAH+YK
9m+NG9NVckosvMoECvxECjJ2AC40qulEP8BPLfPO8VJIoILVTTpOBD8oh9YT
rjjaEF3y9LyLBhiDAwf/Z2vlsM1V+4i75RO0YOy6qcD/neKRi8rNZrnb1QHk
NgFPpkxBzu3wE+tN3CxIh0MxExzcBVn21+c5SqA4QLm2XylKCWMyIJLBap9n
8OVL4vco2Qrfwz1y+zW8PyEvBBDrAIXOICd+gEX5fdc+LkVik7K06EOCGyJd
dVakBrM3XEQrntWIwtECBblpU3xgswvluSP3Kl5rquvQmMaStcgvF4hUazE3
XiUEQoxNCqsa2ZqtFtXfDr1kD2GOSoxNHxhto3MyNagvjunefbUDUej+fSV4
hlmyTSjxDpRdrdtg/Ahs+HITPJMqTWGtP7rrz9Uk1QXBxFvzRBxontLapWHr
6328i6IBb4IsaPfC8vYDVZ0rPyNJvdtzwaHuI9BT9twtOucH/vYtu6y5yndY
BiGMIydqHk974/tZwDVeay6ualNY6DdqMaUhpwGOGxDgtQWnQYiQFVwORnNW
I8sTUrmJdNMYy83fZfrJycs8neiJNKtc8x9WcL1KFXAC8LYFzrLn/A30bBYU
weWLYhcl9m9JAN0u2EDQGDwYG0m2u4s0udPO5ukQDiN+Z2FI7ddGTQlX7GVz
30jOrrDtO+cnqmBbBuQbfA+7T+SM3fAo18voghRWbY2CWks3lToC8U6pY/gl
5fdLIOJ12ag64ZXkrFAtZl9CiwAAgb1FNqEjudkuH44j4Y+lly0Ir60v/i7I
VibZNVuZqIeSfqbvq89HC9uGUbyQPvEna7tNIza2+B160qHLu4oY4nMOAo/B
XBojx93VQoz5ZJa0p85WIJh2BUF1ELx8J5lNAAZAqxMNwqUXguhBIXlgmmoY
jIxBlVMY3Xy8CL2fbZz/CkAaD2/90cF3vH2AK9l3eaIouOPZsOznNRmkbCZx
jmuWqrnVAmZb4PT1GRpMLnb4MIf+LapDIPFlPvW3i6MUAHKq5ZAlg8Zh4j+y
wWi4kfWIcXRRXlkAQZ6CHdmK1tief8y0p+HdFFNC2uvAvVuITmYYS9XjERFh
dvEiEHKCMwUe/WvP7I83q9NcqdF9EtVmG+pwtDJPYMgD+of70F5e8p1JRz72
XFc3vdJBJYlHmnGYEAM39dZDRQewZQ2AQkTt25PmUTvSHZCjWb+0yQZ/v3mK
+J4Aecevwx9gx5ZAy5f5A48/CZx4CzjiDNhxFasGVZk3HLf1WmiKWH6Dz2yT
uK7KR9sysNng+Fk6BKkgCt0a7kzii85ebSAhLO1jc1A396dlyviG8jUiG7H9
7Ix7ukv7NDU1PHqaXtgqAuk1OyXO5de23TvNwVxYOJVr66WuJDMTWG39iWE1
4Ll5zn3OPf5Yj4Z9r7nG3BqknlElaBdwnDUBLXxduVzBEa159slaYBX6OF5t
AmdaPad0YytyuW8XvNgHGIceTHeymNZvu5mS+I3DhhKAZCrXW5/bExOdcpS6
BWTiZ6ykQ5FjNtt6eCy0lWfbqQlalRK8HXDKfIhC5O3cJoBTY9HK8F2JysPu
AmGTonvo1W5AJ7Lc1PkMXlDMeSc8rMRCNO/GSLvm8H5a93gPGjL2iTsB3BqN
R32iHb5dAMmYXFjNV5NnRjy7Ymp8XGWCxDcIex4+Pc8N3Qyq1k6OEkZtL0gk
rU+D8QFvRKTJ61+6Z1XmMa8DB0k2gnjkgR0MNdo8dLkc+BrPyMDUgnXnw9nq
M1pHzCHpboKFd1wBaE4toVg/QH9+9qzwBXHUybWsSjatDqJ/BvQN5Q/f+pPc
hYc7AMvAXHc/Okd66Awog8DKDiqXtioe4KxImXgt5PT7HtyIjhHbbnJOGNVz
LUnggqTADPloDXMuTaHsh+LoYR065ftU6h+PP2p2K4n5Dc6fxx3Bxc/6bJwC
s6hgVS4Mi0H3zlVSuLvn7e0nWsevBwTatxNFNEE9JTM9j3S2NRnqs/B7IYb5
mM7OBFNqwrpGb7X5WlLos84ufvuv16PidNfZjL02wlcxjZO/Yddf57NMGORh
BjJEsQFVhxCu6Py+tdw25IqaFfGVEvOyXgXLQRozVJrWQ4J8XZ29iFEOpu61
1pi8doGaNRw56yKJLEtLLu4UmZJcJyO5yAGn9AAe402btNnhKU/nvhDjDQtr
mtD+hkB5Y56DP6RVnqvWoUEQPeH70MNjoVSUrXMrpUajZQmSsHhohdf9ER2F
t7WUF0u5CkOZhn2iTQOzE+wKLR481wOxZYeBftoJmV0ubTt9jDKBzRSqGRDG
mGHV6QkeFSf3SKleNhkWbPBFULVsr5u6ZvtY5SS1tFls7MAbrujMpM5x/g93
mCUYRlvV1Exp1beWxs7PIawQaTUM2kJOOWGXb/6Pvp+c/WxJ/krXfycQ68fw
We2dFKaQsXGuyJP0SCCR2zEbHdCA7c7ItjIFtoufkULacS8bA0PNJyfVTn/w
pDAXWpB/FGFQUMZSt60lRMqqlf1mq8+iHJ80IcK1Rk8/vBSZMxktDf6QoIrv
TwajakjJPe366IqS4FiCmbenXQCaqaQF+TiL+53y/C5ULmmeMFaDN+zlPU/6
2vLZKpvIqf6981/9z7+CkCt5QF69CsNZPNRbj15hSJsv+wQ+6/8j2KfAEYhI
J+wpVtzj1WtiMq2w+GfW6EFP9k91Ri+x7dbSaR6QZWtf6Pxr/rvD4o9QuOQO
dwhtLI9t9vtl5fTxn+q8Lm/fgMXkwIl7MRQ+vVTOOgtWXFDae1PlL/AWAlxH
c8wF2dF5JDPf//k/8tS+xmKlNO8rRAhunbw1D4OWwGVUnLGECbpd6mLoDSPU
YOT99fGUiPJ04rsWIYfdmjQRFF6VMEGdHL+FsE+QhuOSTyvv5FoLR60jFuvS
pfMyAYLlDlp8uyHhYpT9Us8vuJMpyfacoPmRxGVrOWeWV4fD04YtEMq5UV9c
zxU6L3p5dvGLhrYgjpX6vy1ajFIEwDwcouN690cXrP+Qvd3tuIHHHBBySbwA
luj7P+u5s92Dhf/FmSHhjy9whZgJHmJujvwMAONOq+51O4WdO8OsQrwYOZMq
CyWaTOApOiV4+AKTeTSqSoZMehAGRtFvf33zq/x4tsub7r748mlSIgoYMRvC
G0uUg3CEHkOaxHP3eEJFgYgGNeOhutoQmSYIpIf/q2rzEJrTGI2Y5fs8eG++
zxE91j2IPAgbtZcvsq+Rlr7GPf8Beg7KhaZNBUl3w3nJ5kV3JWYnVOCPRMJO
1Ll2hGT5NHPC7dV2ZBSuA8KoZIJxmHPEOBLWmCEtR6nKU84eijd6lVWMp36P
03GHVea3D5FOgnpHFXaqAolUQRdz3hBIDKOGY0RHYQAQgOk6wFl7t9NvjOoh
tvVxBjMr+S0aidVY946nzqmSKG2rxU56hDPfaBNQDNIU05YLxJYopXCIKEcF
7zgoyhQoE7wPg6X0F4/Qhq5k71fXlwJIoMlHc1jq/1awmLq9YD0zXDJhSbMP
2krkmb/KKPWFgFoyjTjzrlKS8aJb/+HY9aaK6ME68o8HwgBzujvaCkxXTh9o
qPV6Kaf3VBqMmupRHo04EL3cs+mfkzBzRfEeQlkwnFV0yS2q4Co3JWUYwnmo
fEdfvyYbgoeU3OFh47BuFs7BYe1tLC2ClLiALDWy4m8hXRQGOiZ/DZ3d4j2c
/NQ7r75pyO5O6k/Zj9sgwhMhGVB3B9IOWq5BJgM7YbOx8FuRdYu5ypai1MmS
VDqyK3Hu4gsaxU4qmP6rgvm8hDhu11yGCY9/auSN5kNUxIBYII7DRkY0AyC3
RlTYXy12ijGQpTl7zt4LJI5DFwLxb30qth+YatEqWPhCoCrmGYMYFjUGEXt8
PmVtbNLlM+rcTpVKQiFmeGMMMnJVHtyBlVcuM+Kx4x+OfFT5Efg1qtjX9RFV
Vknak6cD0m3/BCOvTYyhOqhVdJW1ivWWadu7sQzbrkBeNx5m69HU8LD02Pvs
VcBAOGzsgMJTRQI6VA8+KidVCf1bAmsJG39rN5tX84cyJ/5Fbv1eWIWHIj7Q
6K91vDaVFjgy9qkAuT8JXW0nFFBLeI30x8QOkjyijNfYWrf5mY4ixn7hsnqQ
VQsS+pqAx1bn68D+zXxKU1FMa4IC5GLQohnEWcijojzomPG1Wo8b6TykzWr7
Ced/aRxTM03uOpbpf9sJ2VMgCLPqD7MX1dPLEaR5jZcBwYXHgc2Q90qiu9mh
+IHINW2+2k1qYtCWvs6xD5r/kRMVZ76Ux5b2oRLgq0p1EP6lK1Ld9zMGT9cL
zX9ojJJWirqavfgzZkE327JiXGNGatlTrdHfTKDWRtorbXKhrvBtsEHdJccB
SgzFADGw3H3D+jtr4t3YhN06wGg2+Ze/yEWuTZCbEkUUAw0I7sPkHjSRyGDP
wHQtWroNMcg2eTYVBIogUKmpVc6i2vrIPSdAcsWndtvZ8AbgtzlgxtOJrk+D
XUNSGkP200K1pMVVm9Cq0LypburjZ0QCLx74GvAm5vvbzcMon/PiIoCy7UVT
SU4qnx/Hh3l5zBaGbLeyUYtpVdfL5tLB+Y2k3BaoB0zNQRAAg5LZ1yaO0dlM
iD3GwCPP7/ISVnTZ1umpIO/8XIvTEfvBUYalqqa6oJcAHB5tQcYQNtz/ykv6
TMZdaDL2gkCpzO9+8ltPh7UhWeXthUNZOA5vXy1a9PekiE20h6rKPdW7SzpE
l8lvcZyqbIepEbyeGSoev4xNUrz+gQj7M6fVhyIL5TdR0MlDDgKdV8IS55/a
skvFCqTND1wXKY9m4eZZNvyUBySMUuX23xYEFPVse9VzI10zphToq34JUhZd
sVfuiGJupP35VoNceexCskY/CAs9ZAwk/XQOuIIs9u0zdgT3MAMMZVbgY4je
xiCbE/1mYNcF1dEKTcyW7l4zrkz2X3AzGnm82hHF2ElFdx5uf4AsZqJBThGp
KzJYMkQBBi3ttPH1kcVKCGsdXn29nnOGrvok9UZkXfDb8uuSQ0ROEfByd1Ub
pt3vTlSAdUvgAJBwGfPhxRPNqYcyfbYRjICcZEORmJp/QDheih+1RF9dLMG1
f9TDxugQT5aYxoZgQRhgw16aIhSgq9sVgUrpWT+qKYBdWtuZsouyIc1/OA0C
lbQy0Whl2JFBJ8yVWAwJBoPkdeKsI7Pf7xgBWlNjryoGaHMOQHS1KSWI4TQE
r4ZQw+uekT9ho9Fab40DpVhWpIKF82DGSKf3lnUXuOtDNgaifrkRTYTZYsuN
ArNfRy/ReRf6SlKGKihkkT50JiBR5SZwIN7MqFahJbXPiMdGV+wXGy2IiiFR
XgyzEbhJmB/D7NZKuxnlGhhz1cxRqcOrodTmMdpw3Iq3SoGHlcKh6sZu3yLI
weRUVAw5Zc1LK2w1YP/3/vNQi6e7piIoAfmAadZhzoW9x/10K/4LU5ZOfRp0
Uq3CgGDkWGCvZkpSAwmYvob1Pj+F87IDfT/FZQAQR1DEuBD5rDQ7Ep7aEyyb
J4GP8lv4GxLd2NcZBpY1g8Ft01FLEIZz7siOhifHNKuLxDijy3jx/KzttN9K
1wxWJwg0eSEIvtrsQvp1MtrLRMM2NT+E6ZjLYYM7qXT9J9l+jcjTauvio+F+
0G0mw23T+P73X7V495W0kRVVQIntMof2NFcxFY3Btx2XrHf/bd2TvMxdF0cg
tE/FbbFzUoX+zgdH8x+KlWfau25+m4dN8xWXPKcpxLlkPsn51pIfOP0cyjf4
H4O27dU1xKseIFdhEWto0ylqYjzIHTmyIMsFTpPO+8zCJAG15a4RvMRvOMaO
L5yMOUsCWZVN06vFihc2tH81CBLKbxgp6hn1J9AK5mcH6m3CJrKy3qZhJEey
UhNt4GE6eOAvnQ9UYKOGhuApsFso/Zn8cBPdseOHv6/rye+UXNMEGdZf2BUW
XjVwpEkmVfcikM17BS3dawEXW3cNzL1b5MWz5yjSFMZzloRpRUJzf/pEgmfT
cmI07cmP0h5qdBQdfgD4/7xDBVhp4zZAF38Jr55LwsHVC7CaEUjOn+5fdw02
F+Q4VTxMYOi03bXr0LLStFbcm6Goe+e/JN9ej3EB1XCyV9srSjHeL2aaA0L1
Rsenc+N9AvqMYTfahkg3dLxUISIZ3kBOGchBhlMgrwSqI5E2RX5Q7wrXqqKg
dz51av2oNCa5gNdbdCgZor89eeNbdbZ1e4bX6XFxpcohUJgGQbfOFIq5n/F3
0OOyYSzQY3AQKtcSTl9v7P83OP4yQBRFvB9d0wy9cqoM5LfZ6mP4dShPe0co
agR18tPG56N1rQToxakejDAdmheJ8nIDjxVRV+tKFQW8CowGrEH1TpCRjTIV
Iok4IODdCIwUPSi8PY8gzZBO7Im2LdQLU4dtv7NiFK3Cz7nvcWUOHoW8uSdH
+KY6sRz336xg/s4UpCqF+eBbYQdmrGsoFBV2E0g5jroTgE49HJYbVUpPGJO3
rYNWeBFbHSqEjIfM9MXCoc17pL6S3cwEYVzIDCL4jSnDLodX6ECjF7ndm6Hb
xJojKBPRuZC4TvpxSHG7zAknxrOvOytN3sox4BqghOS1hYHdyYwykxGFoqTn
GEBl8fZgV75pY+FMmdF6hxafAzXFrNkFDWYfcCIPxODKYDNa2zy2wHkkv5VR
yVvGG5XMW76y1YSx8RHc65EcoFlBRWznSw0y/7x5rHZU7oRr7MX4/HA/U0x4
8EHeO9KHiri8kZ1GV6umg+GwnqRoh0PSusbRC/copmEpvtE1l31npyKPpQOW
SiH70oIy5RpZ4zB49v0IJK631oNSgVjZQnHciR+XPnm+x5NSX90afRk9isvD
HXbdu7ijcnLJvl9fIAWoIg6+shXI/ZIMjk260A0lPzn6GhV+0UuHqJu5oV0o
S0mu1b/uoEbI4Ia83RMJ7X4Dvhk4t69WCQR+6dEnhYJz1g1eLXvHGh+OjwYk
8RoSYJUkjGi9c7pxGKHfnyX1QKbKX6nylZ1Tj7P3XTRaIiHKbUxdtW6keapb
Kf1vRe84lu+X8EtJf/JJ1OWLXfoscZ9b826xMOUDMQVa74FohMX/qoTDqGZM
7Uvg7WTDp6aqmVylYzKSn7DXPzz9EYGQbkmFcY8XKTwq2b9nAQOL5TN8uPrp
xFG8UHMtrC/H2YW3AMs/2tpXjvq5DvOb/pXFkZXWUH2/9z+nS68e/RkkG6ml
ZLIB7raA6VDFDE4cw7dDWj3mI4eK0XiVvmtmrZksxKdMtMlICi3z0twKCXUz
+6VlgOuzNUvMsVVOtfXx62acNmtt8u0mZvzw3tmjjgC9fZ6zGOXm5MMNI94D
j/YcyuWWH7hKTiS6l+/pbInk/SLlX1gq0YPvZC/ewYzl0cq+/CQy1ucTE3K6
SCKsnjyPGeah681zCpQoVQXRjZBYc5haFeG2qKH5Tu08USJ5pOTzFtbmB8Ua
9EGAzaoqwozJ05NcpdUrQcSWWJ5mGKikzctrYVxbEaRvwnlTV5kqcTvVkWq2
oQma2F2REQ6oa/TlF+Jtn7CDAcqdbTk8eciBywDWl2+C7mNNeOB3dwipFagq
BcCBnGOxl3DDmZHVieBARzOFrGAMlyV/eg3qeiKQRTAWg3eDFqbEBKDWZgSu
3bCV+hvzsgzeLAg6919dch6WoV5MhCUFJjnFuoIhmnlM0ipHBd/UWa1NoW6V
iAsl19PYhIptAqIGs1DR5RsQlw/UIxJ2h15C8FsR4UdXp1iGHTxks0e8sVxM
eqf70bCXFZ7l+doNiNJY7us3CbxIL+qGBbPjiWrLqckFTrMZF9lsahRZfdfU
4EElPUEFxzxKrFhhSt0C3gmW8G2IcoYRIXJ12uMXS9b/Bx4ZlHLXE5umQVkm
HCnao8XTyBcW+tF6izvq1zjAMnk7l6TFp/v2bsXKzYwI6NhbRHJq5meZLiUY
PrgtThpiyVfouMekZDExnI/3vWptYkL7CfCf6CWcb//u1wAiuwVutyskg12Z
GmkIvZ+bmGVLwwjlGzObfpA+pxOdPGuGmZu315pr9/4igepEs6ESBMIdkqzb
Zi+gFaM8X7iTEsFfpnyaHLz2Hgm9l++24aRYUWaZCa9toX3EY00v9qKg60fA
aX67hJfS8Ju7pRgSjtJL5gDyOhoDWslfYBTODa+rGAywAoMVXY2cB3UYzGmP
STkhb1Bc4HwbjQ9XfKEgZt0YWJ8VHm8ryqqXdOnvN8XQjScTY0U/kTPTdD5X
98624tgnUJaKb0S9fFOXN5Tg7doQceB0gD+w8KIO84w1uSHYcLRB0fh8lSMd
DKNf4qOaF14qnOyGJjSBx4nAzwjQjyU1Xcd8AQuC3ill0H+WDEPRzkyyYksd
0G5pt+mt/ccHUXSwKvgtfAvp/qw3fTZIF4A0dpcP21n+q4Wa9hFNUtHb90vj
fq2uDYFIsgd55n+ZsBH6r7+CMHQY0r1mrJEkqG/m63YaaB4Cqk5A/dys4nhu
NE4H7CJdDrU13hqFIqWiSNaQ/BUXSZ2edrm88CJjQTXgHKTvQdfvdpSHAxjo
zh8F5tac6i4d7e2KiI5hDzMR4MKvImlzRlCv6Fz22KGEhg/P+kXxpgo+MIaT
vc1dTG8V08DCTut13fOd7iIi4hlCJZ0NCnRmWIIdm1t2LC1MF9tZDKfok8YX
Xmc5rEXQ49Gw2jnCMCXWEqHKSLW0YrxRlZT17nRfabEckFG/cUj/zpfZ6qXM
zIAAz0bUV7eTkBwYIkmYLUm45N9vtFaf9dKTmiYTbgOlR8/ahyP1xwqB/A4E
Sl3nACKiu4/OdNzUStliQuKMMc63uPkzXpl2/WD6iuSzNVP1EJhzhSk4Cyq5
31eg5owahvBYywIT7IHD+L548jputq1AgFcXV185majdFHQ1l/7dpZo6kt7x
MrQN2etRQwQkJ/R8vPgLCJ9dnSoGTDrZ4rusPHvmgpXWXAvZ5Pf+N162NYev
G4UC/5/qmYP+MRGrJ6Vt6Ski8goOPHNakMIAAw+bxNr4kKAQDOhVizA2Ay+S
IV4z5Ax6zZdermBdRpHEv+KZuSXHgocTGisp6uxHjUuV+PnydQd4tJx75pgR
8JCAfoJRwWoK0kd8CB0MZgmRf2Gtl/Pvlr8um580qdwLDhuLK+3+wlqkDGow
gff+QoetsR/Dhq/3uvRWjImlzQoUlvB0bhH3/y3JaxT6sAZnHn/PMQkRraBO
l7y4U2MkGQbsNRF2ku6QV1cQLggTOUWJz2MxjB1Cnj9yUtAj2S6fLG/IBuo/
1Zo7hVXZuDGLMJ71BWOfYOkck/DhOUedG4ZYraTUJdkhl+xpRs/6YVRWrOVQ
5QjTGuVOXqt+Xk8ty3sod1f5g4t7KJqPmbV/dtUdqfoWezfzz7zyBRTSyF4T
COm5CU1XD24ebu+xejVWt1a+Nc66mBxrv5WMnmh8dJ4pp1U7bBQO/u/+QG8u
HmeLsmdpHDDhGI+YU6aH9dyJcOyO+lqbTgwj5GQyINqxjSkNrsFNnlsvqxat
atWITbHb+i4mFx4aYbvLOeiYr0YUUijfNRbxrR03Nvp9Hk5z2K/Rjg2z1wl8
Ufkow8jUTba17OzruF5AvlYyvPCgqnb1DJllT+qJ8//H8PXDzXD/w3T8c94T
YNh/Y5UNkJGMNWCCUtaj3WEXAumGS+v2C2pyJ/d4s6sIWbiK48XzL3CjhU3g
8sNqZkGiSElnqLjajUqo/qg6Ve1mxvRatO+94c3dV8qcCMJIHKyAoUwdyhsI
iJGPyxxcFAnmcbrtN5a1LBXcVuRnk3/7m2rdVwRVn3SRmH5zUUlRq458VKx/
HPwVeVcWMWAYE29oSrW55MwPzHuaXPGbXdCeigLYBbdf3Xys/ySGrt/JZtV5
WpoqVXWyD40h3ImlqNqKh6Se6RqP88PKfgCw7sFg/GV1v7MZRyOvCTTkzAfo
A+H7JzsAaq7UzpudFOafBzhqTHQFP0cIzdL5uK6FgWCAaVIIYvMsmM6pJWLb
PD4R1Zq99yK1cb99vsbAo4CqAr1/aYYam8v3xZjwPaz9TkxVTJ7YpG+XSJKT
V97rc+0kvnBLeNbTzN0jwac8IJCUyfmQJT/5Cfc2nQz9q9Vi2TwgoPwyhIig
y5QcEFWZ69Pmrnokrdvf9A9/qh+DcgUjixzxlgR4oiLRRhqMz+HqvZRh49zx
OhxZ/HckL5PwcDVNNQc8SxxnjyHFaL1dLseX+OVfAmEYR9ZlaVkJyd/MqhvJ
6Knr/Qfxr08kQboCyZL+IB6NTrLFs5rJZyFZK1PlmCsxib+ShWLUkT0P11Gk
IPRFhqsx/kbKTntRQmXPrwrjzCsiAUtUnTW3FkaZvfJLLjcHLkbvvn3Caq9Z
/yc5TlP/v9uaiLjAmt6vbRYfDhq32C8NKgmVevgvGXlCKjlq4Wxb3SGUyl+d
D24kF5/BZjHgsyJ1TktL390smkhnDmsAIsIZqCZTFLQLfYyuTfDB1QGPnQ98
J9w5Ybzaw0Vjq8/UiNK109Y99NBaIOhKfgVGyYbz8FbLVUJua19NYf/BeqhK
jBejLyBMtyPiK2OIQSUERsCxua0U1FhjyKmLQloDiFw7NMla6MgC3xu5Lfrm
Up1qTq+O4YWhdMVuJmvWIed1cJ66q0KEz0uxpJ5jMV/eAMhS1RzgdKiyJ3ON
0VEc/hO3t1IM5GmWv0+3E7Lutr4fo5iIsDXin2HE0KSzRSQ6DwmymX6aD5bU
hQgj8Dg+YLQYQXSivDPIHBINFr2V1tl97z0DHDEx3LZ4UIfRGasp08PfirqC
HMTSn4pgb4ig6zU45s+OyMafaKEKDP6nPubVzaiBD3afIkmhJPnycvQ2PNsm
WpoFZI8BAIQ8Z1OZldsgQVkf1KCGY3aYxT4L21G2s1EAIwykNg0bAeGQZX6J
L7om+R5cwvRcm4PdHXCOJc/kGDnm4t63KnvYy4cAN4mEdUxykwJs4wYECYZY
G/CUCZmHqIpDLgb5Y11Ts0ro9dC2KDDLpiKBbkp38SrqWazLmpHPaPepzsMi
pibBl/jNiBVcLCj+LfA4Yek2QpAwUwgjUlvcC4towwaK3RW2X1xEupe28WHg
vwXCcre0XMbLmiiYbuR54mEQnloCprGlH4gGt5bFPzl82bokE2LzsS5b8MeV
HQVNcESi251YSjMEmNhS2KYXMK/x7gqmz3yqEnAjnyBIyn0sGTXzZNz0ytbq
/qWtNJnVA81Sz4mf+cwejIU5SgpQ7aQXRv4fZM2yf4Ghc1pREist3U5KVtO2
p9QMPrBuCZcZiwXw+s7sFuMsosUkzl6dJePK/0cip3aX5Ju9BfJB3do1MrO4
vsC9KFkGFKHVUMUq1Bz9jbrNTOgfCqFxp4CrCfxDzV/5QC3jIdQow+jqzDkd
S4Q+A0VNp6iddEBV/nOYxfuEXZ2HEj0+hAgzABjDUlb+jdgm9bKqiTHVkYmh
SXI+MEu5h2fWdUC80axOyPlJVWnMBzHOpea1YCJBBZ/M8PBuS9YRA56vI6Sq
ZbH0Q9PtKSSvNNe2Pmu+AdykxF7g9BJ7sAk+Ko8NAVXw8hSmhytooFec2yB7
2SSCYUHYnYuY8c7gHSWD93ChTt/OK0O6dwArls8y7ZsO0jsnB72cIggIj1yH
Y3y4LMKYvGHwct+gUaaZ+Xnz8K/7u7hTnJZkSEH/OrHJTwGxwKTVdmOqNIvm
Itpy/v63o26pxQXJdInoaseRpjLPntMj+7LfLeSaxUNjTW8Ak+O2kXVVxPuB
WGpl/A+h1zxKbEeDwq4UHIPBkalMy2flBLqJWudXkYXmR3ghrOXD9Hp3ek7I
PFH9wEP8Hb82UFC+v//H8Xnuk/lZF7vohI7YUqe3L5+PmkNVXmjWMHSR/J/Q
YQ5QLOZ3kLZSsa7PChXJyFZz37gKcUyUqMsg8o+fd8xzd4qfy2EZHd0qx7F7
ztc0QRfCBpGogB3g4gspTXNl567R+1WKzBY5HwoMO4TpNw4eg61R7WNMhJOf
lz3by1npxxrvtp+qYu6k4xQP6M3QCBlkpKk6BcJABhvk1IV0OEr/PaxYvCrT
EPoTal0Jn0VJD3CXJHN3+lTWM6DGA5wXe0KIWuvWIlcHCUQZJXN8cwJMmAGT
dphZP51jo6xc2wmEL+w+u62VRVT7H6LMnmsxx9DBD+FMAHcn3zWKDhn9Uy4a
fjrTCdioMYSd2Ph8d3pYJ6aFhfQbpP3qZN4rg5gExzR2d1bFffeqSHUoQjfc
oWrtliC66tQkvry8bpWKV5fxILLSJ9z85Tu7r1B3cSLCcpa5LFnm79n1eyZA
ma26+ZvMa6n/Qg761gR1Dzs9DblSbJx3uhiBf8xcTFSmCBhg3YHoNwitml7k
ec/0magNngME6wmCiSGGAyb6YgNiKTGF0iJ+zuaTwEKEWz21DONlrlWnTe27
DQoqaLXtc71gVncDU4QX+IV8X9WNWS9RnaMqXPDFwJyXWItBEdwu7FKRIglz
E7gCaS9WyCfADMWDoI+194yTkERPeDKRvqdOT04PCB4nKLeK6AGWLRGEd/1W
dcW23FBhRUEiMREVc5R0Dv0bC0mk6E0jqnbDrdI9O6RQfbWbJ9Y/Qr8TucBF
ntoOT/kocwJexrg1qEWTGt2K+dv7P9yOWxfltvkCl/RbSV1in4M/eL9eHpHX
C435Xk+wFiEwKVVPdZPNqRkgiGmvLhmGPLkJV0ycFtf0LOTc9ZFelVJdwjME
c9YIQWeplWEQQUh9hM/+taPpco8AhIDAm11qtftZn+fZtKvDiGGy8ARHDE6r
teGu6wjIN/Jz3F065Ndnwm78wATVVhuMjM5zRIqzddQrq3cNXCBmaSclnONL
Oru62kSh7KInAohaV0kScvLh8b6G7cvqY3op51LBN6TshoCX7TWdmmS7yJrc
lMmvJUJ8GKCzIuxgwBYDTTuMem+WhRQnUGZM+rO5FPKLLEn28SMgvkFzsxfP
c8/nYorYFLbvlDEiVSHQyFXeT79y/pCHGh8yAOj+0p0F+XY/bsu69AQGodm8
fcmjySub3jCzZSDi1FMMytFq03rhxytbPiimGR3w8WhIURWBYml+MNKmG7/c
oHX/z6lz9UQYq+wQZ1VVfpC0Wo+pSsD+VkhYgKZ6zTCHMKmFRnSGUkfew1sz
WqJTuomNLvvjIBp2UVhqeoV6DyVfEa9uopWzU6XdTMcDLRLU2o1fccsWhnwR
qd5/M5h6EnFs4Nb/CRN6pSBsZw6TA1+QRqvo5QSEcZxlJ7N9yqv/FkfypR6r
89JeWKqCV95e9MikAkc3hGPoYodf79Dk8T3E6HyEpT68glIckeTFAVm6RWdm
/nVVRLTE1EQLVXF8QApKLhtoTwrmgaRvyxhyPPRPKq6ajyKn2G8SbDEnXA+A
k2l3UtEFi2baukwiSkDMnULdSTWyhbk+cVE+U1GNCkKgpasxHj2dGPQNzixF
1GWLeB5dZZ/lz5mvWvKL8aPFo8OLqHvREOHKlt8k3C6eH+fBuA3Mj/PtpGPH
K0lvTQsYFSt2GNNB/n/YJkcYn9AcHx0/cchujpjyn6Np9QYREnoGPejVRXkU
4xDvDisgd2uXvd5b+/Svi6NWUPkubgdw1gr/TdJ4hYfcqWhMtxzwgVDye8ec
G9v7157PDAaUnrFYq1WuzUHk0ZNneZwLkv52FbCJH+WSgzCc4w0g5ACclda/
0DQx+qaoa86IwF+Tgc+1NsTifPt8r1oDf4rNgbxYOG+bo/skShQybVxFbynG
qhN8Sz0NW3eLWElRm5Mu//4oINKYrp5bVM9CYapb2iREc9U5k2z/xJCo9nRp
QmXl7I99Lex8jasLOcb4gtJFCgxfiIwfFYtsQsMRXEbPVBWNbuByquXidJ1K
lkdImPp491YYx1yvOtihCxxo7sRmekS7F0rYTcUlzn2cidkqP1mvhTbo4Qf4
QqtVGFy5QGOXU1PDfMJQ5uMulMiKZePUEficMeu3/KruZlxFzmjaeVuv3HDL
TsKDo751g8Jv2P+rYJWhH7zNRmmm182XnUt1VAj0TcjjziRTQ9df2CuoYPMv
EVRzt05E/iy26pC3+KKN3FMuBWQbBJpOi3hDLAzoYNptvq7oYDqPM8VowKSQ
Vzamwo98n+CtTkCj5r1TI1pKQm+X4L4+EkMdyiWrin4iLvtcREFABiHLUlxA
TbqmZw0HLu5QJ8y+8oHYbVdcDXSIRKbHB3T3RCv8lsbSzXB/Gqw17Tcj6TQi
MASUb8op+K4fZIRMReDQ4UzLaAodTlEphq0vT2wQUYncjVwPd13+4UvUQXvE
2rhHGUPlwo3g+12sH7+kk/E6PCAqHLHtMKg4q3p1ISzJbdQSxvcQuyClIRuN
0JMwkRHTAWDi4E2lPmJb2DWfaPzVZQqcW3RBGxYCCdiMSeI3Zi8kQs+mp0SZ
Pbd5Vvuo2rG9gEZh4oEUMiY/Ee8mFDF9eXm2NufVb+ANpo4fIUPpgNCUnVAr
8Df/6B1JIYyDJkAZllJ7rUTMVUTNC00TMmBxp9g7tSZDDOiCzQDHsp27JP7T
gtXPQhsiJXcnUL/Ws9gYuob5MCOB4TflX9lEcIHpVYOWkUYhDKVRoRXMOL2Q
Z03tV9vUmxU5e9iybzTOKnnjVOQgazzHff7dU3PBTiWW0k6acZ74DuqgvqEr
C24k7ysHgLKVQhk/x1rdnhV8ih8T5XkabEMIJMb7tA+BJ4XNDWmMYz2i66qR
xSkYD1G6fFnvkN/66paAIRr3oF+NXkI2L6KwwaR+zqEwA+6nfdf6rZt7mTId
fdVmveXB0ij/OOWM8ktt6JRtT4V5JhEGXnqySRPt0q3b+OUlDSVChW2bXzjA
LwGRlGnSgVoh72fwUfaRs6OrUu3OVgOfI0pDfZUPsG6bDQwsW1g+a7Ru0zIr
68xCXGsFSaX/0BUvJ62HYvbKmlvAn8iOGTcB6PKsHXnfk+aGmfHLz5+Se+Dk
rq9lN85yv1R1QZChlAuXmDQKIuMawqRGkl+Ky7WLX6A0SU0UsldOqkSZmfjR
tbj+GxK362a2JxlxehEBsbaNQZypbg8AGlF2/1VD19e9Ct0MCLwfd9svidBN
mU1J/fsDkVbEbSKZk9Z6MYdY/ZgNLOgHusxRp5z+d54GKvTruG1IYW678OXT
ecyy5DDUGzp1bnTs1sn66xyrIplj0XLLXkrFXhiF4Buj+cvPqQjf3ugkH6l6
/RehFlUbmo7aFBKuNdtYos3v7bv38MpjLq1VQ17NDBp+Jv7JcR5sqYTn1dXG
4ZMM5JH69bFqCjtokFX+4ZwS5DPY2bBWVN+15cNdO6xqqWmaHaoDYd7tOnTk
AGD8/Qz1usg7oIRXhjir3SZFSX5FF7z7NLGHYm5OrdN1NMFurJT2+Ns5ShUp
l5Mu0BnPJUTsyTtejcU52wd4UIjS2BWfxM9f20a1wweh0aNEGVmTanJyfev4
gyZ8TV0Y6O0eRckT8FgLRXSLfZbXZ+2J5IgC47Uws1dCimQEjMUB3n0Sto17
fR4ejnS4Mqi5P+YmmS0OI951Z2Z7Nz9kPDczB67TriXqlvBEZCkDolEs1C/c
hQ3QMaUYIhZsg7hFevqtASjsgFRWod5rZ46SohfmpRCIALxD+j9ciimKaygO
L7d0xnZraP/J8omLaHEFBTiTv/e/JDkLtqqmISZILOrIBP57YD5TO1aG2fuc
8kHZ2C/CCH15i3rD4lUpt/wuUQPN4936RUCPd6mC5PBUj275xYY7CS8b/BXW
HN4nwOUQtVVpEvLhADwdYArw8GNcE7CnxOtzJDDXr1vTzuKJSm5hMKGFKjtt
65JUMjz34TZT/9XRFp+4FcIBsQdQGecz3l1IjWemZ8EzFbJOFQfWN+ong8i1
1+xNxeunE66s2hijqg3sudvnc8VpDJ8WwWWfdw/KxWiO4CjjxvUhfTX5X1Jh
98MhdHLngMc2SF+V1Sje6Bs2/sZXiHO1mXBGOUtCd3DWd+n0kllKYbKORRWM
sexBzxzH9MmmPDLpUWxmGadXeugA/+/ewyJn1SN70Z8uAzWQ5tMfq09l/Sa8
AV5nQwqsC0QTJYwLYu5NZIqR4WomZSucTOR1GVenG7W9H80+gLJf/tnhbbpk
QaE8NB/mdptueJlUtj6zDyeHjBoJZbOWYF0e/Snkz1yyfa9rGxE0O4bfCNSz
AwoAL2mnGt+0BGUsxBbtiUsj55t6grxoDrOHTtNKq7Z/gjy53He+/vBtkfrL
QddEc4d3uYHnFTcr75i0j3YIqiDe2Ov6Sb0q0zb499VQD0qDtUShkD9SI8qh
3A2tx9g471tD1HrW4kcuzrAtMS36euMLPc2SXXcvkGw8sXsR9wFn4If44f+I
11oRP0nr2ez/02Y1MS3KkRjo/vZNaPMS8884wTVUCumYPV/G8Cx7kLB4HKOM
L58fqKRkSj6taorSDl6flxs/wU6GH68iUOsoRdKnKm/y2aojX6juVj7HkuyA
hT4enLItXSlLI8kL8c5llRS43vHCPZxASJ5RcwBgheDNyotzNpxNUFUD8bJp
m19xrVrq10OHlyFWzwd7ZBpYugA3Poa/lElMrIqbYm1JzQEYeP6fjSHpV0dI
4+CBgsYXJn4mv+IirvYLq4qBXvAueNhGKJOkVmJk34dIvC3dcaVOP/q3hV1W
WTdnA11xXafnIVVwHBHd/dxU0+ccf8CF/tGX1AVFANQDT3uc2ba4ROllc7vG
xh+UppY/xo3WGbPIM0/EPjz2ZbBUJH7Ri2DnJHuBX12OVfjRq3D5cupDmGpC
VPTeDzuwx4X4hgAtyLq59vlMP1kca1dCsfm5ldrMkYs2zmc8Dsvig+5uj9E7
o7StIIMF9IV1Dk/SH+OjaV3RXYAqOEz955z7NR4LLm5w0kYCjwDbBvJioMN9
ax0D/6uCGLUDztvGQvSbtzOjUkEmSKUOTu11+i4S2/pbQsEdRhVZ+7HvsRUn
I7UUr5zx0Jm15aUQapNx4LZy2pL8dYxBlP6HTKRl8LlVf4P/zAjJNuQb1GOF
hdXFDLm4C9chMnng34LcGnWp6hz9IqDsN1QL9EiUaLu8mCrE+pRIT4OgA4OE
EGh6JfC4yX0PapZeaiGcZgPgkoFq7X2wzzReou9Ro6Wgw6020elfMXXmS9Jx
q2wwOaEDxBrsb2WL27X3fZm8Rx/60SuTVM5i3fpx27PyaZzeMgHgv7si/Ky3
f4tcOmSrV4JqGsPEtXI3oUtjx8wQqwHi50iw7wFsUkFabK9o3LjtN47gU0Oy
7kM+BriDUcTFhUqn5xq/xoW90ifZQv4Awjz45GF+2BljcpiL2x1klgE5zRrp
oHDhj3+ROw27tocKsn6ylpbM4isQTtwQqZUFeGL83HsYRoqGfIKPDioZqPsc
2AHzj3NEi8OW/uACqsfc3KNLl5KerNOUCCgRh7pmbsHplmzZoMMzoYztOM80
4DdQWrkdXuPw+McI1R0rDTljRHQ3hqEdC/tWY3zb4crRUlqzJvVE6YUktt6b
x3/bRYXS2mcs2Naj4+vcz7VYRz8gSoIJ8HlMR8wYW9ht7M4vKktMivxebWN/
LWQkLErLBYxaHjPa+bn4x6CrL3G27LDMQ4Lb4wwi+7Va2mIZ07a69/o0v9k7
yM0q+o1oHvTfUFVZHhGUnX0QdUYwfWFHpman354SLc38NwDXbsBRsGszIwHE
Ff1hObRhhxjn5eQCKC3+HIALEZl5kF/JWU0C84Wkp5B1iewf3k4aW2MS+maQ
rIzeDaWJo9kAptF96ymORVSe5h418qKK/jRau87d+FeHL8/757xrXi/ScRb5
f8OPJIGNYJp8WF8qKY7BC/CeI/ZUcQjTxZmEZOul89rLmFY7vFy0LHVWsN5J
zn+uUPnH0EDsGM9OvEdngmjITuEqQOcFrb6olTUb2jwKUnyLYirPqp6aY87C
wKBg2ZYxhQyZ8zkyaEOgG+xVL7URbasC0SgEhGTjb1PkZMIoB2jxz6sU7pdo
A/eQCxvd1NKoAkd/K8OoG4RgngOGvNBAcPbPw1T/A5AoDrPnZzzMzv/dqAsV
Ncbfe1lIK0ssiqoJuAU48MBt4lDJXS+r+s4R50DKuK7KLewD3o/JJit/xhC5
tvsZFss/LfiKJCxFF1TMTg6MPvGj55ht+Uws0mdWzLhMs8TGpHnwZUNMATAG
1TJIyrOatyb4hWW/yc8skaz1fXHWIj9GH0WrWqZP6jJJ13cIei9O0xBUl3BX
yByi3blESziORUsR1zTC93P4Ujlcbs/7PuifX+Sg3MEvifbEGVq46KNTuWzk
pDEYZ6NO7AR7EdUQo739tLoLDYbf4nPo1hInHAyjGNqHzTqQ6FLGmUOHFyal
Ajf6yonazqdz+4qHPQnYeDBOzZQMw4R4Nk2a59m07COS8SzNI7uiMZQf4HAX
aB9lBbhwF0lhijUoujGPhVNnp//bKFicO6UsnZR/ubLwFHjLSRcU/GxT5uOB
IWN1PzVOFAIlf2JG+fy1htgStrxXO9bEVCWZ4l0aQasNepaQaqX+o3WJMZKM
YUlQGR4Ng51MRToBeqdYGYR60MQgGsBB7iIfQR1ujd3tYczP5Uv8muYK38Hf
Xl9MRoJjiiMMSae3RQHOnjH47eI5jhjqUO6NlUsfIGHJbUUQ48+vm9eBB7SB
ZiZZwnoOX41C/VHpxWYSvHA9iDgQ8Q6z7vLxJQy0ig26HsTyVusNyYSPMBhV
nwDTN+VPyZMWmnh9YUwbtst75COsdA4VzocIpyh8VugEH86hG9utXoz0S4Xh
/zlWPleDJMI7uq17Fw/CsBgXJSxLgivQTqGWewG1awJHKv8NQ3QcXJEJjH40
F0Xuoa03mKfb3ZwBR4i3morkvwIOY/g1GdJK8XeycAOjFXecXTzoMv2kgwTd
aRq8tmYZfHr9SP7VhdR89dO7T68GAZ0iZYy7VeGJrZeNpuHZThC2ckqgXdZW
RSxjL/I0rHwi61p6OfTiJIb80DWDupSwsttZFvy+6u9gusb35p3M0EeCOgot
s1gse2ZdlPf8mYWxulTmCc06cpPezZBIzAGuueCdaisT2753D+88KyVZ2c57
vAKinXoMegQtL9KTbXFmLxea62OELNiuBVjzjdR+oPHiQpILBY6I67vaz7Ad
0JtLNli8OZv17w3W5qvN0Sxg4TfUSbKjWwHGbvve8DxqEHDwIpuukiNsD8gE
tAfZ3LpaMVRfK37foVSK+mnq6YEZsF4t2LOleB2Og71rdxvPY0yveC07x2q/
jA5ZuGA+QRjge3bsv/Agh/59kxwPfB5XrABC56HdjKfhKHbdRBdTuA/ZSEHJ
yxWEHPraS1SbwctSmtVWAiwhh9xokTlOD2ehO4c9fA1/M4QUUgSWIDiwZqrg
3WpFNHSDaadvxP8VXcA3nlT3VS39Qjr6nCOD5FuQXw+ShvcBfQlPrIZyzIvh
PkggcvPtg9uMoYxhlMQWJ9vorrBdnTDQgzp2T10zuLbR7SwHRNLsnLsf7Qjs
vsX1Usp9kuAW1a54H11EtErotwSsVz7Q52mRAxQCRIbSvQx5pkphGaE8rvmA
GbWLt2eSufVPgGUdNppNWWGC9/5X5jVUYOt1xenKa1+tzdbT7ylQNlpgaSuP
HI/AKXPJEi0xUI3slnWXC7daOLrUO7NOUoQtoOYvX8cXwHcoRmMszlCew+K2
jTCnDqIWXIjW744n8xABWHYBl/ejkKLfLS4Vf4VVFAGnUZThhXB5ExcnKnh4
TouTG9wi5dkqMCJpqUu/QZlakTcmQEhQV99gu69i4cClOTYtc54etOHcPC0o
YiPUfREP3mDgTNJOgfHbZOKcpQgkEYEd8abeJux/TFbXUj61bFe5DC7Kg8+5
owsscz7TOjN+0hk7bLjmB60tCo8ReI6sXYoffvuLnReIzdYl7HrYbOj7x3fP
Gth9xcoZEPK7cmlK6LwV4YLwZRGzXV8uReIcDu3eUKbi/VdrJ+CK4HIjhuwr
HtUhEBn6TA/ftXkH9XVA31yN7lPTwj7g5jkAoETmqOm1yhnNUuAiJF3nMpkL
6LSR5tPvzzPYoCfL5HK0zybkhDBO/5S1dn5/ZtoEUG3n0NXuAmKuLJzj3Na6
mqSGW8hH9i6p+Fiq8zD+MRJoftyQabdAdhXDH6I1IJX3z48oRETa1ImIVETL
PvR9rhz54ZJifhpbbjfMLHvB59EL/oVSZQQmtmIJeodW5UdvxkDqk8I2x3MM
5dY4t1rzzIeeyneVKgmn49A51LkKt2JUdKgFsSUH30N46cRcI9cUibTK3Ykf
xipp0sZafC8k8PJbsjcKrql2rXa7OE8GBVh4I3/p02Xoaj1mcIOxKLbLNTVg
2OUIOI5OwKF+KY+xJc7KXIGvMlIlh59PikJ2i3rasV0+WsV4zArQlfskshpk
Dyk1MtGK/URlWu1WVcy50YxY/zSXQH7JnmxE1sNEqTWbqiv1Ky4kCvnfxH8/
MczrCeLnIFNsKSzQ4TH91jLzZurqHMMI4JR4isrSmQcZST+DhmTwXCIBy0T0
U4PLj7pQtad89/zYDHrJC6X7QB2MI2TY0D6BVTIomWZ1utY2Szd9RN0w0EIl
0NLY4cG92RqR1lYdzzzbi3nNLq1Vd9ozwZzYcmisJKwurbzuUQFjMIA7YrGV
O4YU3sK535SPCue9sTvGE6Kz4LuiJdtAsicAQ6+VVGTkLAUYjcMuExBNKOy3
GRQVLfux8WwdEZDxUqd+vCa0AC96xvkEVebWNxV8Ge5u4HC4Iy+VpT9omnSD
aItAPaJp4T1e7U0iPxwm/XSS51crfaZcVbmybh6t38GZoh01z2kKf6f+BI2s
Qx0D9xh4eRRKD7ZnZuebVsHoIxlp/eAUDHwdnuRa6htSZvE7lX3ncdP8fMav
wogJVYCM5c5EBJ5a9/9+g2Rn2+rGoelbNpPo5R6eg3+/+mpRVSVBduceB099
VQkBvcLEmY55dNnQk9zqQABAz+DcKBA2FmwB9qrrmysdCV4Hx0aiMJKopjpq
bj8ILg0og6A3vDE9PqoInDpq/JT49o+g4XSogLZXqF+cx0IWfPHhHXD4RyNL
oaiMvPlMoQfZQ3qEwr3Ni0B9Se0CFYWGlMDuMsXKHTDqc8tIwdPjVfvO4o2f
05sc86UGQBjAdO9vsWO3ydxdhqL7wf+7nM2CGRDxbxqySJd5pfFSU/27B5D5
TOOsSeDaiDAqj3gL9d7LZInqhNs0fegZ+5Eyp/E17deCd4QevnbS9qjHxj3V
G9QDBMdr/VMWLBhp7AZ5xJRcQE7IR6viZChTlzDFOSZqr7+nr7gCHMaFbPHj
QiBLZ5b4Hfp1mFuo0l2ALaSry1372lFfBBwwTkNuzlETnG26aBCtifU7DfR5
KGRwcX8JQLN7fi0m9tr8NSLtEL44gjrx3CdWyzTj/4HcMFHfGO98ReEgLgJQ
KnWU4jwetwKOglEJxYhyB5uKTBSZsqRJKVzJcTJSY31EHcVmvWkOtjCOvdPY
dq19zo9JTNPRyBLEfgYNyqJqQgHoq4GghrtdQwcAuBZw7k916JDmndi8DYru
3G2lEOvxxpI+7yeM5pab5utDPvLLhUu7ovh7HQhQriqkHJnVMGPau9Dxa7Dd
576YFNqiOi4eKiULBcLqR96IrBFUxFrcphvwoHkaaLthLZhUY1z7S9NVFQPd
wOwWm4iDe5Ds9cukB5a4JFQs2pF39BXFpTOP3UVYILyQB5vXOfxkRf0jFVHq
sJp0d3ltD/Kv3qSXIMihx5bOF0/DGIuCyufs4KUBEilEJSkyIhHrDeqjR9Us
KeWDu52KT0c+FmHRmYY3EABgqJGe+p/FXBw40ivCYAUynsy40yRdSZOCzz7X
z+Zk2Og1egVP5W59ku87pnaNImQsgfFEDoeXw0SwZr7U8XmDyvnTPOIFZL/V
dIQiSem62Iws1qm9s83NmwI7IwEiL7IPScsNS+EvQoGoVmRYJbd25gvJzJ+4
VbhMuEeW2HSeR6fRhkhpQOEosODtEyeyoDpG7morm5PMKAhV0+4RisRu8ndq
8ukIfLbsC5oIN0+jnlmEjudG1sKmMQuuzm80OtmAFUSgf+YAVv/iFq35Ufsg
dhoaHBaV0doQ6s/gnMvVNMVZu+5WiHmWnU8YgPoMlG6n0BaeLOciveLhseSJ
MbxsOht0dGy9MTiQxhzOPtLTVnuYaKolskMTmXFEjeXkABedkWsnagDDDsBD
JhV+zpzU6rTiquBpMD71FyCwtxnbGbrts0qKzjPcf6TmUb2r3klo8h6XPub/
M2tty6k2xkMdEGzUjhGw8r2fojBdwrWJHNxwVGzhYIZ9GBKP5vzdX9dtJgaQ
olwVd9Sq9FkCn+u+boSG5dXo6lk5MxRLTPeFYuU0Dfj5luXfDdZN8/zZEmUj
37keyPvkgpCto93ztKcnGrobU03Bq8HqyQz0MyPqbAJJTodimDrIResxJK1i
1Se4UU3Ezz7jpHJzXpQHpdLlb5qjyMDeC3WrCNMaNfj0ohaQLm/dR8Lp1uCf
Idml0h77XYyjLZYbfTXh2hGeabFpWjvwUM2sdEr9AMRL5nymDi7DcsjVgCAY
EWS7zAr4aitzQhvBRZHEeLI/fnUB98tzNVlbivii8KVcMDbbWBNzVR6jjlpr
9LDpyLWGGMCJldiKHpdcvtYiX12QIUvL+AMssd75W2MwjkIb+DVnH/BXki1F
shQsCX61PniPywattuFV0hz0y8qdGWOaIX5zEfsDXWj3t3pCIS6HcDB7r5Rf
GvQDrUC09kpgexKDomGXjJhcgxcHSm3os3Xa6k9x3MicfTL8x/h/CJbHgKWo
x/+FkhpSsyOn0fbqm6318NOOvZzQ1yd+DQQ+wV6Z4LdR+pg2SZ67oMeNeVo5
rdZsB2ltgmur/fYUKzdxo2G2NHXOFgWcEroCkRcZnl9cr9Zeg9VM46Dx/1Y5
BP1aFybgQlie1F03LZN3FQ6rgOhwmNILqhSBUQ3FPuWWe6Gu1OK/3CdZiTyV
wUPdhGPdr0birQP7rkJcl+SdVFMZVlbN3C+aPo8oTYpB1mzIM8N+RR6Bhyf4
SnRLLpCoJVw35qjszmh57Q8VUwaknNqPmQFr5wEIZQyZO+kVVn3HlP0Tb1/Z
W/Yv9q9mYm4ghlciER7H3sgcVdLYpqT8Cwl2mtqIqxS9GOY/MwMY8OPwl/X9
y6KWP5+TxhzN7WijYekO9Y6Hj3HaqLYtsvVPqocxip1tLPqZBmZB8kLNpY3D
xXpyFufNBClwBxh6SDDX6glAIEDImiDw0/fbwoiPvJgJpyE2FfHuqw7jZcKt
d0ltOywjQtlECp1/8pkXMpxM4uBszNpvkh2FUbSpkH+3O4kYQXGANIqSINiw
Tp3Wc5b0u36yjhkz+e6ShocdMxJCzkUnvudZ2sQbaifVI86O7aUW6T3PdLWn
EHoZhITnye9kFjAwt17Pn1bTDwi2YT0W4ahg4QAHEOPaLZ7Q5LzXF4aQeK0X
VHsHo/KOnIxhIXG+F3mszgLEi6gQdVA1hjWknJmZiV6CQV59Y/inEjBote6s
KnfXICQnzGZXsy7EyvQ/5+S7Tsag9E0UHMgQKy0+MCaSjM0bz2bkyhJVKhMr
DfTqNFYDR1q00TSaxym8YT8Nn7uSx8rp6QctSp0Lj1q9O4JG5iKMkE/p8hgD
dSl30QqA9YFFbu6lDPOBSQxK7SWYUvTjt2vgp4gQt/py5iRHV3jhdVBjPuO2
qV3Fd7jHeKlEF53GYn3x2dfaG8WpdvWYWxaz7MfknH30jifIYPu8Smn39FGn
eTll1ujsg2PpL3wI3V6qku7LB4QNKvtPJzLad6bATR7V7GjOfX3Ym0ewWg00
ixnXU9Y+UH6AO3h29B8/lm9/ijfZsbfU4n3VGTLQjORE9mN7oaijj2Nb15SG
1y1iXNAHpHz46nuJv+SjGfCac8QCgB0Z+3ussesoZAMyZtLTHUt2F6pmz88Q
abDwLs9ho1BHlVYit01iMt0C+O8OQKyq70qSE94vqgb/HHsTf262QsTEldU+
36NWYMIBZMz/GGS81IMDzY4RmWevMelYER0V9Hzivp9HXWf3XgrU/CKA0xIz
aW/YUxXpkdVjlwmAnDSXsEMt3h0ZD/g+RNLIV+mtHnWWnOLObe1O0qZSC+G0
XvxmxXCklQxLnKZTCBNuMouuuvq8iAYJ/cu4NbSv6gOeK+dBUOlfDiQnFPVI
6lvrSAyn11pOePbU4+SheEXXBnWoeKvyIJF59Yl9wYavBB7K6HdzBxh7Yvq2
14tWgkTB7kpnQU/GXKFuhg5/vcZgjydqcIhPzwlWScEWzgDh3eqQkZAErufQ
waD6McJq5F4YDeKS5BrCUniXJFwGR4ujCD0JVptYgRmJTf2AAgMb5PUTDinB
oySZfVCXQPEojdYts8C1RJKhiL8VbgtDz3vVs/UEIdJ+saAFMWykb39BWlXn
seLB7Wwn+wtCwgR/BAWQZIR+QIVPRUpxWNKscNGU4iOfPwT/DcKsgjs/yhpG
CMw07yHCYM+RpsbvOn/m2LuTM+wrt2WE/gO3TU7EbeqLmvi0oaWIkjjrviu7
XIRKjCjekBH2vm9X4otlphX95ceIb9JT6H6BulVkpKzj5kOfSoUcTzaTEn3V
4+mmebrxBReRhDsFtr6KUR8uQnT1Iyyy91wS0+x6Tg/Bo7g5TR8EhmKmZV9b
eyRk1gQfk8h1NzCWXAaxRrvCDAPgVf+ESfZy47xNA/iWQ1YPQHpC8vUXw4nJ
cuL5Whrjm4ddKGKWRDpPMUspsacfI74NBFUBBaTh25mEoyGbY91trfWk2pT7
D6fQYWXeHz0S58hKDxjmLwfxJOwkCa+latMrjeT4dB6irNZh7HqICLCuKz1N
ifPRVjcJSSU4rsNfG7DCHOkt1amepw2ZMNMyaKxBYWdSFtCpNmjU2SLn7XC3
J0LAXLRgfaHlubMWvgxaij3nQZzB6sfxHh2TTN84u+vxxfe1NcIP4D2L65pf
I8AaD9LcSITxJpECug6p5/c5SHcxbtkZm7q5fe7InRbxx7hS2LTySYUeYLXQ
b35Lej2HOxvnao5/pPusXlodoIFQwI1dFA1Juadq392EEeTChekSUMLp4fpu
P95sEQ/U+i/sqms0y1tySdFQcs8Ip+tllQ2USCfotu43MbwXI85RiDa8yQ5b
F6XlAX1EVw1O7rVkiAKLDgg9VFIgXhXyjhqggdlRtkQQZXkXbVQTPEW129w+
puYXV/VMHslPx/L+c/OcRtEmOfK8K9fuOC30+KGCuE6U7TS50S5G4SLIBzSU
+gJhzE/OAMC6C4seQgYdQYjLf2wOr7G6lxvtNRpz7PANJvd8sE2dYWRJPy+x
vuPZ2krn7m0XxNDmjGYyzd9dH+edp0SU+4ckuWYEBpjOVBUGfbzONb5nd/ZZ
0fbF3t1I8nFLyQdAkPv6K+ftSWyTPg988eu0EHbt/jlq3bfv4qTupiTbUjwG
/NriEwDlSelkDPzGIS6F1sAoiKjfrAu1yaNeKtn8CcxEf0/CBLL4CxLtOwwI
YKTDaJFIcTWyEBskrVmfPxWnU32yyxfc+KuBAENQtl1nH/S9aK8psBxmdbVc
R4I/LujB87hNEzKs9MDiKawsqrXn4xITfb+faFhYnHzwMzSFsJII5X63v6k4
w2pPykXf1n+H/+iMjSpLKmteaZnLAPlB0QjPLOcpqh3WNvcSzPNa1FqYTGbY
fTBaPJ7LPnPK7sQ04740wjxBcF1hKQDi6Vmx+nqGDjL8u4DBPc3olocCqKS9
nA8PV/gxmkAq7qlHTvyEAC/8zotsEmpwOoL70j9PeKtDfi2Japwvvrsnz/0J
OmU0Sp+Rm76FrbmmzeTSPLEBE0LRzqG3I3tbv/N0WEw2CUHUIRBbkfJPvOv6
q90cw+9DfTNDSPiE10qTrCRQiVSuSLKhcDyxvxcd2s+SqklXQH2Qv6ru/zcr
pEPGwUMHfLSViubAD6o0WHOX/xXIGgFw6qVR6CVyaS9vpKizMTKwqRwEnX41
y6dYCJfZmsPSVuEwHW6V+tU5s8VHKOioBO6c9BOkbl36X4PxHTtnu+4IVkth
Ah7UCzrTqEl7V7yybU0U1jyUdqe65uYA4i0YproIHH3Lwce7CQosB2FunPdZ
CesoTt+rkQfoSSiuFl4PCbglhtbiwoAGsqYFTnz3B5UZu01AaY7b/9TEGOMz
ryVsCOQVtn15dAUru8jY9l/8h+eYibhERAhW+7mV5l2IxrkCxOvDOkQvcQGW
xORfrg3iLa4t+U3Gt9VLk+dNwGaycb1jLNMLs3hpo/ZTrYDkL/dJpAYHYJ/5
ryhIC5QDHozHSY8/fbOj9LopA/JfZUSEy9se9mrAPRLDOF319zID/4fL4NJA
ZJe5kSMB2kjiE3/iTFejuBWfYEBrPY0RsNcsBegBFEextc3Hq0cD6+yX/3zl
jGc123NhZVJj8vD92queXgv2AgGdbNZth6jJjCTm4VPQ8uc9iVkkUHhpEY30
rtFiwLF+/y8+qX5L+ILNLxyBsbI30qcagHsWatB2suyC0ocWcyC4h6OrUj3d
Y1xubUnhoM4qnnYOfJEbMFiQ1fZ8nvQtoT8+93AyYtrPYBinvahp69/ayYXS
bvb72G1hpEXCDOlv5ymzCdT4+QAh13OSM2dt3LsdPmrI0NmcYRPxXLFYMhYm
g1I1GNXPoi9sEtws4BwRcjMKyBmGeFkPVpu+RaTwYSL14utVl/9A52VHTnm9
t/PN+jJozk1HXfdOf+LBJxQJ58IUolX6QoS9D+EwFPz7nzQBVK/t/IbNQgjQ
53ve+8dl9w/FvQKleRdznMe5pDYwJA0PEbYWrud326IS7lN4pTyg0L/vMesw
PcdPRbPoDLs5lXjWb1S7z6STAUcxd2CzHOYwONpIhQyumi9TouH5lBZximXF
PQ+Cn9y5uo384+s/TZdDC5ozt7rQu74PjstBqMtfcQJImeOudIOPiXLds9+Q
d2auxyyfRmXPj139XexIZDzek6TRAkZHUhtbUwh1+9BVOuLFzPLPFM8Fln1D
G8O8P6UanFmR6IMeJs6sssrT77X1zEtEKYEAKIXgtJCHU8CbKznDN8LgtOJd
EUbpysOAtjjjOBHsS4SY4f66Fg7HWdaA6wg7hro3VYFktLPjNFKLSqV8gVOw
6FbSnrDF7Jln8xYjbYQ8eCJLKmHZgIRRb/XY9f4vZn4ABWO10ufX17+TefHq
ukjbPzSb6jHMRTXZubtG/XNzMOdTO3B8gfZanPjP7/ZkRpWpFOuGApu56IAu
SBCrUN1iz8VqKmy4nClZdqOislImhoQA29SzmhV1lgyqbxpYAKnkmfxKXGCB
bkEa5Y07S1L3ktjOZCpc3YDlFeKOp2SSC1fc5NBuqKtNmR3oiEkZarEXN5dJ
CXhLa1SqmQJE9zxwYFqkj7kt+Dgy7KqeR64uFxhbpeMq7+WiC/XBIgRHkm0c
PY71v1eVhAE2l2Ycv4Q/3gwcJWVBJzHYgi2lJCgRcaQrVNEnOLFvs8gVAKHm
QDmIHz7wmlZePWgIeitgYb7aMr1FnlkuYF/xIdTx7ot5Trgarw5y8R3JgCvd
wmJgM0OxA0BAKESBiXWSLUeB6S4m9LlNkmXcuJeI4XofbfUXLeJDwOGbBgG+
zGXTYDNURAfV+rLiIokqGWWNVrX/dXKVVSHEXyHx7tYn8AMuVfD5vn/l14KJ
4HlNiC7liNy22jLFkt/fDAv9P3ygsrCYU/xGz6dL2nds7RDxFM/5ThJYiW+i
JTMgltPxkUSfi4swip3cENV9M3uRKti9bdZud26O39+HWZe4bxTevjYbdwJ5
le0CVgW1UDarFr3mq6CFC0VamR7dt+hS9cr34eYncn/fTvnBxBppCvTyz3Mx
DNXaA72SKY9Kr6KaKx2zIvv1M/Zydz1/BTkqRsrmlGbeoQdOXBK1nfmHiqXz
FBKRLoO/ziMvdq+6e+oLpfd4J+xUJU7PNzj6WHOc6NdNxM9N0DJNc92amgww
irILaJAzGyW9eW69a4bR2a3OVe8TdzsEEQhx56LLALClEVdizRwIS7pEH/OT
q4bcfdijgGneNZvePI9xxduNrQhi8m4EZtDKxsB/rV5qcj/lPrvtAiKEhS1h
IPW6l4uRNBcwVkEoW/k+T2Bunmj6qQIuWaWoyp519MIq2AHq8RvRNLt3O0Lv
WwiJsft0NzudZkGAEOxJk1kWOi6p9xEtgvJVG47LjXEurDJVROPhm249aYwx
50GMdY/4yrUtxTIjYZ2kdGQQzabIeU1xIehNUE87/KsrImmyL8N2wVFpmv8v
B0V/SFOOMCJU303CHjyvC2xDLVdB2CE6L0x5V05BXZz0TGN3ZDt/o7EbcCqf
MlO/ny8L/7QDwc4W/ZIivXC0TMmBStjVDzRn5DqI4AtsGpHA5qOxGiHw2mmC
34mqYhhLIlgb5wUH7XHu9XKFdTYPmtIWwFM7SbgBOQNZ1lCj1pfRRKululOu
s7/HVhlU7hxzobkQHgcrDYUE7R0uZo3diMAoY1dPCfQl3gBryKmRaI6w5nRC
WnnpPPeGa8cw3JIFhXlTOUwNzzFRxKwFzzdPaVNfcLFVg/YAMN6DZAobRUJi
3wMXhtlTzuUG7oE3vZcwQXSvG0LC1evaK6JKudWX7eik4YODm20TSe12H+BL
O8dj5cP679R1Tx14vttfzbVT0GV4AZiTv9DGgPuAsdDNV3TK7SDH7o6nzZ9D
feBTTkTUB4zA489xEV/KLqtFr3LyDhoR+SFICEoh+6cI6S4H7yO752suTRhw
bU9kxUOAesDV3sFNIGTyOncQtFvpahLFgN+6AwF5tl8R2BnhCmDo2l4Qx2Ob
ZeVr4SWPbqmBUs8440vQa8OfMqu5YIyEoW5CzEovUEE1mII6Iw+gayBGNR9Y
yeTiOfTgQextXxGlYVsqEQHeCHsIpUb5UV9K4+miHDpvw+Dvd3LzjlkF7Q0w
mtHxEv/fHqgpNBr3GBuKbASDhgk6k8+3myVwG7to4gwyBIeY+eeh6l+awXQX
XCrBUQdQ0Zth4kA6iLL5Mss5FniqPJObbZtpfPMhvT2377eqEPgVzCEnUNlr
NNX0wnLjNVdo5kYCW5iA/kcwBX0ALta56bE5Z3lP//wAvAdP6EGjWAZhG6l1
Y0BeVJ4Zb5mXsITVewLn8RjahVQIJvaH7BPAzSEwO3ARTlZ9B+9vAv913Xqk
8xYqyMp8Q9GvenFtjORQi/ejAejCVXempqGr0NDEXP7r5E54EuMcxnSRpHEx
GDsc/4DxZdNHR2tm4xNmoUVA4qAp5uDDa2W/mZ/QKpncWKQ+l4L2Aevexm6D
Eh3f3QQaRuLiAjk4+68f7d8ysRyDbsR2oLa2jYXEj3TN7VbUgGkPl6whPycU
rFnWa2y/p8L17uw3oH4zKx2nbW5F6eS/yNs8i/9PGkvhO4PRNjaqZ9ClDsPX
EKWznNhL43HyJHjPff38YZNw+IIdrOhUupo811q7+7JOt5tn+m63Eo51rEeE
2rIa5SSKI4I0s4ONdVpV21sRxy6hhzKB0rvHGzfSfnRT3oBFx4DrF8IqZatS
3E4Z6KEuFMczVVUcAs+o0gXpqT6SjXe5BmKPPjWcpcqA4khhXFOo47HdYhb0
aQBjKThR62PRRAE35C01WrcFMG+1hGXGVPLfNR8HlLQ28aDFLJRz9Oh6iffv
ypJlXuZ85/TiCLihygd0AHFBt9DrCzn5f8xmlxWFtBjjQmFFACxNAjI64AGm
jLK7G2Ei0U7ZIOYhkytgLXEl8ttQl7mgIL70ltKypeG56rIkqv2t21IsKrs3
GA9Qfs/cttHwE2x9r4u7qrL7a8WVvi+REVNR2upNhJhouASX1B5dZbrXyNOV
wWcoefQxPtibhbLYEx2ulk3TQBiFI7DAPOux5YRG/TX9iYWyeb11bJ7cv813
ePQQQKECMCTcS8X5xxTpFHx7TS8GjwwxA3EW04mwXDML0KifSFrNe9drxFjZ
IAxUJlWABU6zCZfZINQiL2n1w9CGh+kZjRV9SecHkZZl6is/wEtaQpKnCfO+
qDZaEPdwrcXNPFFQMkPyk4iRV+OFjn3+nEpoM++6g/RTN18LkvzLDKBxcXL7
Mh8CsLgppViS5E+stAJHAtBl5HNRwSXgvm0hfzJVOXihTye7glqUSsISKeTQ
IAORVpR6UzVlMPrrAAxRR4LAku5Atx1RIYee/C8tND+9G/HqrlqZf96g7PGq
bYqNXjnRNjtB4JSUBEm9/WsfqCRaiCYyH+Z10jqcEtrk7+c8lhu7Yi62BVV+
IWtXsucr3wrZ9ZqN8q0/Zmi0y4h0RMJACZmJNAEBlkIWogzxCWqVLAelCDz7
kmCOV41/TsKYfKxaRP2OqWD7QstcFIk71Y7fpR0ejykA03uwplsxCzi+Vgf+
HbZwOi+nitBg8KDp7J40KYogrZxB/lXOezN2yC7v6FX71BYVCNYtpXAZdmrh
2jnALdvlF6TSHgMnY2ynEiDswXoAIb3s8Q1ZpH2VmI5lvJpVUUgIukYa039R
/nQNFp8QzOEHxCcnHxsO8bDNWNXHpm2OhuBe1ywish70tEoOCPi32wk1xp0c
Jb3UIdNWemqVg8lGLjB3epkjuFqtagh/EeyD5BROOVxovmfknqyaXMRll6UX
W1gUtJmiYYwVt2WTNpLS5zBrWPq2izHs3bDgGYapdVMpX4Bs423WQESmv481
/PAiawxVUnZE79bWzScIxeX67hRUaRJoSmVG8IBk32VUcM1AfSNvfAciZmYd
/zZ7AT8c9KXoAdEIFfZrGa3wpRs7/KmQo5Q7LloSc5iFUIYIcqRTv1KXk25H
MZ1jjZ19x8tbCSH6MZ4ungyZgq8mYtNPcvzZ9ZnNrMTylsPLVVLTZzVbtJYT
96k+MvkeUh5zsnIVLd2NgX2YBqFx+0pZyULmLz1WAB1A6x2aObjbqhe5NwYf
YHHdGUh2v0+i+YAfpqdBqTGlDTXFRoSn/xSi0twa4LxqXJjj0Auf7qs2CgUZ
SB4nCLUUUCu9JpQI1Ec0W9E2WY5ZEIsjNGpo9MRjnTEvOofRq2RRKibWZkvo
VxjdxWBgnZUNyRVTauGWTgr5qPC7G/CBUt4t2Tf+WTshPOAxFcCPn27NcDg/
NtAWPlkaeVZprWFxdKn6PYbRhiJDi74OxBtiI2l6pZC20IhZCsYxE+UWl80s
sl1PsUz4z6zrJYVa8+t4TyvJBM9cnAvJCWrYMDxJ6kgiRJXKyJe5RvyyZTv5
nvgd11yEEmdQIUzZty3nVgWs2aku5h4zUxGL3Sh5wmmmKccWq+39gvVXAQ/A
xIy9Nwg0b3awV4C+5EEH5+sdVPm6adEr+TT0PTNgTqAgZLPC6mMqbra4Gj93
JgaP4C4zP7mnBBggjpIlWKQY6ppQRFFgtXwig4+cBjXd8GlPw83Qtb8ZtsI9
SvDcTEThzhQJjJ9uU9oCsXe50oQvUvZm+txEm577Pc9X1pivTvzOavMOcHhr
p3JzvtTF7PXvnGsD2+OZo2hMgVoTs5Hfu4r+0fxIz/Weq+AQQTG+92bVY5v7
bqgluicWooDSC14M1dsrKiA+o0IKjh/iII1+fzkuO46jb2SA8d0eRwtLIeo0
lt62KOyzn80661iGRrLtm41ZsgemvgkYnotLdBMBIWKVvj/Yw2DFp0As4uTJ
fIUXPGmhJaOT+8U+YuIYD3IbTpgBF5CjO+Vj7yMhXM0yAnjYiTDGx7zJJF9J
ncCnXgbkkudguZ0blI1CkKiCltTUExB7SQ/KPO7wtdXCeX24pMcFvZDZL+XA
t7uvgna3+ATqKxQ+DZ05NF4Fpu5ocSHiEQqXWac/9YfRyauKM4LSQoJ5OFEP
hYYhYGuqsBabIma5olHiEMlyqOa6itNf9Cb+nJIw+7WFdDT+KMAgNNERh3ho
5QCHBOdE3bnNFsHP3v1zecAkhTGBFlyXlffyqb8OLHTp7MvUgcQr/szKv7z8
vp2A2N5MGYaZLlygqnjYrYFmGUstEdqOD8oUPJ96BZAnYR8rgz3h5HvCF/7x
S98uOCQN4rDOz7tXaMsfp2xbvNGbWRXpLKOyQ5G4zfRPiYbvpUXeS72yYrXQ
cvbqEZVwBM5b0qI2y2k6unLF8gUoHVy6/9DsP93rSUBhLcTnlUobjG3K49w/
ZJUAXsg7Xm8E2U/+tq38cRj/Ea/AKPxAuAiZFpV6Bw5vhXoacvGYXZNZUeXa
/JKT/7FU6mN//lUqXMt3irMM+z7GLZYADJrfpEuoxjpJIODr4sDF19vdJfeE
Sj1eaF9jutRyfyOuPHF3PywuemlXegiKGusIwyljaed0gYd+LPTRAqxNc5Dy
FyTZ+QfMunG91M50cdK6Zhd7rSUbGlB1rQOTrNts+CMApsqDokFujZ/4uGB2
M+wuDiH/LZJrHcYvqmxvuRq7Pu3l5lP1A1JiNyBby6wXWu+87HULyHveBnI6
ZsKw0mKMbkEKRr9cmSQWy5kEQRffn+tq5yY5ASbbVylZrdE5T0h5mipnvceG
BOkfuYvh+QUfWrIVLoiX5Dw0EtC1ABt1GidlYcDq/hWn4W4/znY+9oZtUuA+
MnDuKi/rADIwlCfOMPibX6T5+sGkeGjGLceXdt279JhadS+cy+n/GPGKR6IZ
KN7RNhYyUPWHg8aU7Wf/xgn8jEGCy29gt7em2XlJdFZZO0DYRjXjHYRmXB8L
2EoxyiTGv/LvTXwcmTCMb55/11RtYEb3NJPioVZz0Yk+oIoAIJO6w613fB1M
NHwmoCq5aTW08fwh/ldgfve8bqZ+/B5JpjMk3h0591vjx5Jw1hWNdHCFj3KN
7uBh4vlbJivI4u3XhO4yE2y/pdvHYtvuWZHTbzU7J9ElPamowFJCTReL9IVm
tCgshHluiGQzgmywgkDPokX/yYldZh4FK38NO7YpzC+iUyI0x/X5ACP6BriG
FcDQ99n+jjrQqE6aX5wDkIdns5ccSao2brrIimN8It45rkTCJnQKLldJgOEP
RXiSg12s8XvRcHCB93i91gCYe12G9MC8NvwD5lHI6KQEet+79ibzv1JUMIwG
DiCJ+LC2O42Sj7aJFV65JhG2ntYwxsnLrOF29Ikx6vpAu7C4CnUbBP1Q6s5T
/NJnM4ZgCK/dFzxonYNS4wt3lWhztKrnhiT0VO4B55K/eVfm2OoZ/HOV/a9t
2nCIlzEs4yP690SosiiadNRdzIJcxKMrXO0gLvr1niXXC/GhAqd9Bs76PnBj
u2pXHMdBkQp+qGA1jgHanCCsHqVVEys6cPv6JI5AhdAD85PDtC0HNT/TKMNN
/GjavTCnMTArqKRPI515/3TihKHLj0qAKfOhndw0tHnBWgKtcEbZQEGbFhSc
5yJcYOV2qxuWOgrcLFx4aVIIbDdTaQaRuRYwI2rSH0snMDGAxGGtfCVLkV+e
6z1r1zpm9JsgKzCL9xjiAe7tyjw81qq+ODuUcauc8f/4oqAxKwb/+9mOX4dr
NR7YDRXvQBvoaloGz4omnZKFCf2owek2xSVK0YYqZfVVHsOcr7xOaGLgAazi
8I6FNIqCDA0btpCzj3knSx5MQYiGe5yjZXPxy/fcVkNJvRoDBP8vptVh9PW8
gSZev575TqWqBw+z+pUSHnuaOyfaSKPWb8bYGhUxB4rX3BKFYmwieXABrLwQ
gn1oCfzNDAqTmn7ECNpzufEd3wwJ2azQMoEcYq4rQq3I8rJu21NS1lMVpu5H
kmF+073wpo9QyqVReNsLrj8OHae+Ikmzi1KA7Y8lnbLtvtcUqRDrupomN6J9
UYWxFt3hvqoTYIuqrOTlbRVNII30X3r8H/8Ekie3tCT11wrSA377qPGx7W3w
1M0Tf6Mw4mi/byuYfbBS/h+YVzbMGtI7wfeFnw9eH3X43s+JbeWCxobkD+mW
bdNRV8EazYq/JjJZcACu6PGLg4hfiPKUQkQv3ZD+KjUIU3Vs85PdGEDtKTTE
jjj0ktdzycRr/u5f3d6kQ1fXP7+F1gvFODSx02lBejsUSIKPFYusRVwhGuAB
LKp7s/la6hOy66i6CoeEXwvg2M2+mvOyGYjnu4ZeY//KB0+7qukV1G9Wcphb
bY4EdfRzix5tOgjc8ygoCsBXoK2DHfKa9TWQQDiX34lBzJEQFuZdfERJfzHv
BgpVLXXKgTzaBqqOAB+1YhJfItXYDMLBJ3Qk8f3gGMbUwoIWpgEnKq4KgUfE
2CRKqxNt2PITiuwT2lWsEstUsoa5XpP+/JVTXyFIevVA4yoMUm5Yfnzz+v8V
6I8fszra0ee9LBykiSoyHiTVY8+AHGcOdj0MWBDmztMuEA7wxDRLEeT31srr
2F7U16KAYOAVfcPAztbdCbMrrM8SYYxYFmghIIDgG2Jb4Jr21sUT4kxCwdML
A0RvMEdNr8Vm+zYYLU1f+arEo9WM98gIhIMbnUu/S06I6ebyohvQKpv/eEnl
8ZDVh7ITa7xiPV5Z4XxrbVX6HVpZz/dUcV6kBdxKPINybXBA0F09iUnH6txX
gy/SPrxejfwHbx184flXmBb7ByehPUBEk5bvBnqqRtltscVWqpZwJMwmsDkp
ybGDeT850tymDf60e4Atj1uAaRtVroa88hAxA96shy2B3TK+LoyLr5Fy44WR
wlGO1nlUdp8PIacviUpdOdqmvcDlDvMpKZlizt9noz5j9iTdkNTEbFIDaD9V
IGwWNmt5JbowdGnr63rTOl9r/pzlZQ91Yw3Fte2V3oimnvwtz7Z+++VEW5Wa
TSn0ie/702gytxaeTyIxauQ+RMdYuxgp02NAXEyyIGcoifPIFmDKs7oW1GPJ
+r+8utw3AIL0+euP+RzMRUawo2Fs5ONHr1PbIV8E3mKxbfmXc178UC7rnVUT
uaWe55vAaVlKAx+3BfaCjp9cbfcj1n/6+LPsK3HngCNlPp6OUHWFQqiA0Stw
N7LyvPJKsbTgs30XXog4YmGzO714uU2LPgEjU+gzQFBt907THOHekBDx7TEy
7JLyKFxTF9r6ANw7PnWqVBanACfGUYdw2UhiMbN90xE0Ui+tkurzDlwiFOig
G7ZF4drw7Cbd4hdBphPAVW46Xbg19OvltCVH5AES6CDy++vAC/ty+mzcNPKc
1VTJs+oLycHpUk8HfOvT7BoEghJ5+5D6Jv34lhRm6cxg7kK7Twdd/KtONRxk
Ea2H223fsNV6LDS6p/YF9W6cAKzx+BcV9qSc+qL6HT590mAhImH7jdkoMail
Mktq0+Tw4i5lny88Q2dzzrCfjtwp97erdxSGt0BeX/DvtBYg3yEZH/0609bD
JnLzjOMip0Zob3dx8xFT8Y9ddCiy2eCfMdnyApyN4fH+dD+ePm4Br9K6M7Tv
EmljToevJ9W4LpaDVyqJdvy5ux0LkCknli9LlPiackSa6bEN4baKOGazhBWn
GzmyKyXdo7zrbTpMfNlJ7O+4JAm8FA2+UWRSAras8hmuNIXwhnUNrdTRp/Yp
JeBkKAD6xbRgbR5nOjAWozaeNHFvWkXRPsE8Z9kUusfzI/9gSexL4V2mCM/C
2l92aWx3Y6QP/57V5BBcIGjE+S44dK1GHk/vutQvcClHKnJyB/uEN5rDWcEi
tVAELsr2M0HAgZVv1fVYQlOqvjDQZaaztzswUL/gLNmrvBtbWWchCl9dCprP
F+1ot6a8GUCrbsesUR0cB5Td+WRLkbjOGLuZj6XgHB6UAOO1kWCDRsqsv3px
BXBClXfIyKqfPovO0HAQcVmfKaHRDZWnYXH+guT1mJc1Vmk3aPJQbNVPFSUr
btmbjmyDcxCXhKSPlUksJ+LPyuM69AEcZS2YljlFTmDMZ4GlQsXB+bVo/CiE
5cfn2x9t1YNmxxK/SebVH1+CxtRvousLpBTqAuo+t0oP77juuAIqKzeK1KRb
djCDmGGwVNLOtXIo4zLP3NCruZIaOvBRiuB5A2c+FLxkcowsjKTQZzfSbGDh
5ZJWu9V+J9gWuVRMf7Cyx7Ehc1+5fEUGjRy8SGEZCMElOEv8QRz5TmwONih+
3ZAoMUSpagFK6L2GGKjDTm+PiOtm4a1CmXbKC66C22fibgUUyQslYXYc1c8M
J1wU65+0r1QoY2GL0XOf0uW1h60mMxxkMbDKHSd32vlytCofboTWO/7TfoN4
qhKPRXKGi5Cio5t4CfGQDBReANhZIrUfAk2AaRjOtW7s8pwi9v2qfSvBSae1
TtOQjx5IbLjUkP3V/4UqkmHJi2Hg4U1WLWe/f4j7/df6D3+MaK7Vd5ebdpmS
eMi6Cg0rwJateA03skB+0LM+ajtD+7Lf/Y6OOL2VYGWZOL9tZvDITA6nTva3
V/hoAxcJE5xhMCl2vnZfwo5ZRrqwyNRxW57ooWg5J1xqmkKqQfsHdjyt+hce
wtpNgLHNQNkk+xhOrxXyUY0UxhLchllq/i+e8YjlzAKtho3p3dsZl+o183Rg
fpIIkjgPCIW9fYsua6dAT6nuqfUEhS2vW8Wb8DSP2FkdsJBgYt2B3EzKV4Xz
1om3g5nkh+nSr7Dp+7yOgMDrUF8mg+8QyuqoKaxzWVv7sHsxWzCBfdlmqrBJ
e+uLZyXZdsnl0ZRrXl54FkgQtndi6s84G6YmZKavgISge0Fkyn6CzeR644hL
RzG4hP/1lWj3Dnhbee8Yc9pA5Et3BVdB4giJpbKiNFUFWcG8Tm0Uqj1E7UsR
4MvJGJnyPs0HyJwlnUJ9HALHVLdQIGGUGiYa8Orgla8vhciqO1TG8gxa1NCb
OuYKCMchKhCwKsZ2nObcTrWsqGC3zoXD5vti3OeBQMaH25/0w/v7xFjmhqBk
y/THPXtTtlemtDptCmjXWWgRPxNkPjEswFVF87xGyRQVwDagshi1HtsOHAEE
Gzug4FVhWBn1ypDvqxn1oAjDi71QA52KzhyCQ9KeiAPLKlICjkV565vXlMc6
lk5y2wZBTWsrkxX0l56u0LpSYtBSjf3kuBBLiiprx4jH49Yp1NSva6IC5uU3
aaijgutxmdo7aRLo7v4w7Jd1toGHOtxDRQk5q9Q9SCYybfKqK+9itSEpZ0a5
jyqeQ6CISHdhCFaOQC198ab/UdwxZGuGjHG6ovKaE9mCOUdYkb2aCvHfNjyS
e3pwhCxq/ZP056qA731CoMewf1+BGBOHaqBKIeKy3XOseFQQRhALeQyU+1Lx
jG4MQzPNo+nAm5o5Z05I+o5eiCOu0KzITrns8S+UBjxnfL+Psoj8X66NH0/o
LZFmtWcgLH8X1bVfuhyp43TkNWJTB4dAMA7PwkovA0nMC1OEkqPX35uRHDrf
kFdjo5Rh4LlvxDYrXYBv6sX4QZWHKg2beOKj0mWGzfBC9z+Ce37vG1lmv/TH
PvN+VDi54tG7XH7mS/4t2c7By5q3c+m4aPYiE+NvR+MMTrEKvev1xgK9GdT1
gbRws8deUyMQWA+UMBQA3jD42hw7IlYSEDGtczCEdUMXNXUDhg/7Jh+anU3V
y4BRdlNNak58UHxWld4xOxN1Gd6iPlFFyr2bu9N3nLpASt/AIm7bex/cLv1K
R7kP+s9GMVccT1UVVvBXqj3bQoROqqBvmS5SkUDrls3wQ1dXJ6MHdKG9RizN
5sj8p/6a2xlFqcmkl5Ej4iBPuIviJOhc73qrAFkRlB7FGmMoexJuJQONYhmn
xj5AyIycfib8mqYGxhf8NNJx5pccKruf8f8OGHOHRqRHFLFCTYe7467GEUhl
ew8d2kpO0Ae4AVLPtlR/flz+OONWzJ6boAMsN+TnOI3Dl8RVpLP0T3t/2yYz
j1/fbaN8zR177KUfDigG4F2JPgjKQ1e4sdk0Vbf9JuU9iSvuMCFz20PEewcl
m12sBcuC3zjaFtwAM0QPbHJVmuyxVTXayWMVoluaHk4CUSRkfJF2fzNzqI4/
ryFP0hYCDydf6KBKI93slEFL7n+P82qoTGM/WIkxDWDgnzbzUfTnuD4RAxfc
AI9s/VdH7I9vgXgEHoPaOTddyjM5YoIvOyyPvePP3BH5WDXIRGcqNGy8ob9j
RQMamPR/8cBq1tyZkElJhbdPGCmtQTITuM6gg1vrz8BR/GW4ITbnw5ZzzW9I
pmPRwPtZUgEgO5d3SRQAikY2i8idnhYxJFNVhFrQKqeUIWj3OY+rOM+jf6f9
tcyVIg5ktVb1pq8rhUlMtI0rN5qWTwL3pSR3ncC2FqKxrjx/0N6oVtwTkyZs
ch4hLVRuthNWF6J2snu3pfXmAAu8/mVo/7I7zoh91dXwXdpVewHH5wiuSypV
0K/3HwyqkAp/ccjpiteaVa6NVASe6w6tkDgnmA4NP04dvU4NirT21R6SKxtf
tXKclvMAnmcWiGHGytbDERvtljH5TPdS9ptDQrt3sAA9i0XvsT73DBprssGB
/rtqav6z8H51IDLnfsAJ3bsrh+0vqDuhIG5443RZ3T6E5l2S59uOhKkZ2F2S
lMaxEhF+x0wbMdLhjWamQdcuFq8LQpMpbkZ1FR+TmnjaJUrQLq0S6hoRrdMj
W8iZfanwx0ECccIco0lZBJo+j4Ree0x3YsUqdWkoU5ulR5CV7blrakMQXO99
Y/gY1VkE5DpDIIFFzHZAhA7MiB6+5xdCx2DE7zp5UH9lrslq/az0bX78HopX
PuP5scLXfI/ZzZLpzphAkfHqofYCcEFTU6tbMFrzpEzuZPfRpoUb0C+M3FeQ
cdj8ASUgtbMtKY5VemjlotR6OBamUV4FcjhNLuvmzt3ZctoZwh2q7cH1Tewj
5pUHEs0uTQiEOtSb8n5SnESZZQruGKX5ozKUT+VU/om09X6/Y8NfRaEBJSt/
K5Plmfi5LQMm9l6oGjlslSes+r5wnG1ysFTI77fZ/CDqrrV1GcwKE8Qq6JSm
iixbEUeAHvlmCHJpmFln949q69JzBY127LkohRD0bH/HHYST0K5V51rCHUPt
IOWcU+MOCVitCx7MSpTKrx2K6dPkkNIz0i+7OiM3AYCCpWmQkUejO74rjELC
ctQdqJ9ZXXN+dtKWxcT8dGinaGhPlZAjJCm4YPxToT1UVwxRqE4fZHFlHBiu
XRcxTxi2pCBOwhd/BREXoeB8nb9pRVuAS6Yqpwnk8fMD4GpcKLS4xyDwOXhA
KJ54r+GUM09Uk1HuH36yysqmYYyAVk9X/cMo2eq+ZnraiWyJH7lu4ed5t0e7
ODkSmHjFjYncDSlubcGU5CG2kGCurakGRxiR3vBCuizlpvRaEavy5PCVCzpr
RTj1KMhaVz6awSi458VzkprGcwHFfcez4Iqky4Um1RmMxoWif0TgqrNXsjYe
e6vwDxB860sKIFm9FaNnwTozLjED66+pHZCFudmPC5h/91GYWoOmHMjTUbSi
RkjNVDFCg6wduJp7GDs2QpS4ZZwpGSzFupz1MYkKzndNemNn0Rz2SdM7zlmv
y4EmM80ZUxxymWdoQEoDRB3zeiYLW/7rd4XvcH5IphwIijO2OyOSRRItJjb9
y5iTZiZy5ROReiStRlZkeZyorqhi7m/rHDaw0Sq+EiMIlBf0hEU5jHU/3WtZ
hKzIA9py4zc5NxKOEtRlJ1mJ9fDVWvmRQFgU+TcpK+QafLVKceGcFWPQWvYU
WSXGSToWq9cghGKYBstwiZZzjCdd7Mt4q75te625jLd4OKdMUCqblwp1ZWpg
Wokrfozxb8RPn88KHXTqmvvPEdIq/xZXa9UCjYzprOHlwY+OLPjvlX7rklnJ
W8yo0xGc5GXQORIdB9tiETrzofgwaEBwwzkPTqn42iE+ECwIfMCoaTUGiQ+8
YswsM41Y+H3V06HTmivNeg16gc7rX2k78AafqsNF/R8ZM2VTnXiO7JyopLVi
fWNWVucFPmNPE2rayrVk+BmOi79FZQwYyjrz0nCiqt/nb/zohU7U6/mmyFbW
QwrdG7qFH4WONQVGAGylV312Jd4TeSisvYBBta9ypo7Z/BWudzbQwyrom0yz
q32LhDW2zxcQ4KGqKvJT/V7r2EMrNHPF1Aaau5wqXflXIp7EpuC4OmWf61aX
JXIqe/ZTWRLSV4Mv3BG7A933bDsYGYCgWHu2dg9Vp3HTFAHozn4HuwfpAPT9
u5Mio99sZMHrTVrcE0E2QxnF3EwIa4oGLXtvjYqFYHPBHYIy8LsBs46WI5cq
u4C2am02sCReuFHockue7QqJaug+UofpFrQ+muhi5caC8lG4EF2WyXRMLtXT
U4bzrWRva9XvUDkeSgAPObSHpg4XWJNpcJiiEHUqQrq9PoQzUiOLTnkMVpKV
1F5ldHxg+BOSfAuUkKGnZEeTHruWpa6JGr2Mo8FNYq6J3I+bEXsK2owxLCKx
31msHAR89mydWfgyNjvJMlu153ioRh4ulOdY8tvZTdZhI9URBqcjRWsCwTqe
hm8y1pJEzVndoYyJ5StXZU7+1F7ZM9mtPdlkZ7Kv4PDMKQFil6zwWlc2DpNF
b01IG/K7nKr4byz1MXouIdkl+X84NKv2UVw3AJzWMT9ZVW6aO4oxwFlvGnMa
rX0WVCpoihquPzKAGNxwYVpj15L1u+LK28EkLk24PisfoOgujqvju15JtSX4
h6US6qiK2Q2T0ouMwTgn5g6wI9RZqZb4muiZvqqPgG4K6cXgodI3MVixmdoR
IIkmo4+aq8/s11xDl+vPqPJCSQGXJPoYGB8Q+sIzsWQ+D2QMAYJFqaE2bPUB
BZ7LXm8HJb4zzhcNKu2V4FF+AyBuK2OCjsaIFm/rWQQmesLcRJ6OGyDG0X8b
amcT2BdjpMOC7VkRp25PyHZ4R4V0iZfUOgOuxW/7r1qAzDCa0oPb1jMElfoC
+v9u4Ou32OzNQo1cSFFmgGpmbLCuH/neXYf8kzC7aA0yhzPj/Jxr8+TUnyIO
+TiVHt0nSwQHvY5A0c5yZ39ZAkkZ74Xt9enclzMVz8qecrkK7XK3kF3QKjyp
qY0NgbP7Gzr2kEt6cbXCQdJEn0MBXXe+8pWtoen8ZNv+YgljXnRSKa7lRVhz
aL6dr0gvYY/zGwbgmxSswxdw1U5XFXhU4yRxpVYOzWxnUSDKvhJWH5dB0MtP
GhuN/iMqm8x2q2tWHtN+dXROl5VZxqmNdrrFJVphcrAWycOxXXvpof92ef2u
AF9MxD2gAG1iFk/nJ8m9i41tJQxTtoVi9s6yZr0NdQM47ObLOoPPIdq6qItb
Jc3iRVAvaGquBogMDFMFf8cthUJ39D4nhmtHPcWWiAnHwyYuiFe0bI6CehsP
Sf0kZ4HDDqKdiE0sgjzdW0VVYXu3dmGGl6NEdu09kjFOdb1BMTBGm8PnY0hH
RUdVOtnnlpXlOn8CPWsi20ftHy4CzxH+3usdzUExjusJENJ4U7qkpS6cNcW3
c3Dm1is55rQtXyiOT4w9rchH6c70IPJT1HxELL/g82oDhWVh+KdQrTPRJ1CH
1AYWWwDWQ3/SASMEWbzliofwDWcD4UBjHeFHt/e5+RvcETs+SYuHKF6k65qG
3A/7ZGDc+CpVZiM01+Mv2kTEpk354v5zWhcEomXyeb2LHMho8vx0cC5AiBew
ucumqoTLyF9zuZX+fpZ8TE/+LvNDXikC/frGwsQu56DPsfIvAEdqK2FLNaTl
2nsaRFM52fAcEEMkrpH2gbDPpk6ClQEILv3zhRgXYiuWpBdPgcgc2qIsPg7y
TRZvrGidUx44D7Z26byDWXKGDh5Pgv7C10DSDIE8xJFnyoSU2o6rAWkToGNF
45NdF6gIRg+6FDv0CBMH/ekEXZNoSD8Lm+1jErde3ZCVCOWVv/Ydivwj5zmy
+KPX9lOhdQRbK/4D9alQdTzDt6YKpxZph0rOKUp0ApbVgORHRhFEpqm01mqS
xtsirpSow6UAtnPjaNdITCOjliksiA0dpuWyAF42v8soDWxWzUc2Wg2jGaPN
vUN2dYTIDSvacco/93l3FGBlSiBkAqfawsOL9AzH9yY2qlfgvDuVwG3UJ1xm
3Bc/h6VidztfyZxPm0sVCFihjFLEw76pkOgqrzr1npyBHVDyMQmKpVBONEDU
OPi5b2fTXi5g6Xi0NKJ4H3ZqJyj2XvI4J47aBF2VXHFI2WRoxmcF1Ie7lUhy
id4QnvPBg+ihTwhLvMWj33sPISuhrFHjWZeQvQpnGkP4uJp8zsMTT1DK3e8/
xEfrwNbKkbQIVAanFNMhPd7SfTuOZJmVLL1WTvXFErhQ3L2456cdIgS/Apiz
nB0phUxYGz+y65QyVrWC4SCDer7fDXfmOuv844GJy5yUoZOYXg28ICLzGH9I
OCeSUV4D5YORZZ8F0CXzQHt+QnE81IYU+gpS2gqmKj4hChTkXJqeF/UyOJXQ
bjoWTsMTfoCtoHXzVVU20MwviG7YEh+jPcqWRfutL+ABOK+fvrl3tbjbtLlE
vlC//N8ekMCvEdizv4lQ7tPMjuJH7j1QpGQ2xJbrkAgMEbHBRxT0LCP9PUO+
8xcwdO50NsT4iG8GS6n7hDn6MeZsCexCvrgE6L2PuERTlimZ14AixX2l0Vqu
ipCJtjMTkIWTVDyMtcM7EamgsfqLWNTlI1iAeRG0MAjE3x07hBxoqIZSeY7s
FkRBaVpX2dHF0c5/pskw8KDU9vXbuNaI7yn8PzoBV3G1zHvpkIEZeV+07EvU
CUsGgDAv/FxXuKmB0vakVAZ5hUuH4aQ8TESuAG2I6PzLh3GcGJCTql3iH531
yyWXtL29OZQJ7PD7Nsf+lo02yEHyyrSvn3QcGpPk65l6aoDGu0ujkyD0TG/s
HzQo/4b8pkEDr51APB1Ls56u7GxIJXVyZdtTuCRcjcfsLubyINDHgjoJPiDV
T0HmB7UL7CRUPYJNrF/qtdnkftcgAL7rszhQEP2SmlhxlmDgbxGv5dzqk3l2
CvUItqg6Qojlu3bonYxZdV7t3zgAJGIzORTwEioqXeqIzTcIhqauhqOw9R9D
PZaQTziwh1kOwXi/NWIo3Cf73bHVYlQMJSN9dTlFOB/e+rzMlZzNd7nNyBga
G6oBC6KSyBgQxZa6BEDTWlk/WcBuCegzkC9MxSAFkM2/eGY3SoHLZ8IbZpNn
WorBe2tFsMoRgt8Lw16ZgSiizMukcSF4oNTaBAPi0nYra19SWRIFwz3OxIOW
2qriUgXzH+TUkQBt010t+OLK6r1FSRlqyKP5iuo+gq+7/sBqT7JW0aik8NBF
A2ohc2VNAj3JB/KloyT7wU6gHlFOQ5OflMXN0GlYUqrpWHSkQL8xb3iv2wvD
L2tAa9SLTdfYbDGOZI4f3pRh6VzNJAxqMen3/S19bJnDDuMzdTjtAfUOeUUJ
q1Lis76pWyZo1FhckK0F5ahgdjTC6THHYgLBtZCHH1/EaHctoxkCO/29qcyE
cWmCiTzgYLr1FNAbMYc0g3eRf5CYk2bB2yeduaPzj7eFvlBJbtrxX8V8UgSp
QemGyd9I1M4Fd8DIlBv9YjRDJinElNo8PNzlEpshynL/bjAvUYHF6Xebb7SE
g/6SRI8WprTFdA+RQv+nyOR5/sPk8kvEQppM1WNl29ZzmkQfgGQV8JIuHWPQ
ovUx49J5Ne3eYEFYoIe+s2S04myAQ4mbuTq/EMJFHEX2bY6uyu1I9Fu6DMfx
6xZV6UvtsG0T2WAmwcf4hvHbUcyNCA0XyefT9+09gjWha1zJKAcZs+5nMKG0
J7NdJr9gRH05Q0UPTNZT8QsH5Fp/Y6lqrP4DReu5ArPdJCvjhLz/AmeYWJGq
nYi7/+fvhHzpV1pUW6C52347J9f3ErYwJgWs313lVfcgqgC/TPZ6d6pFrO/g
Fy3P6fukiVUzyD20MjeTBqEdw/b+Ua8pY/A4aIPkOIAKqeFmHDLDbU2Z9+we
PrecelFDHmBf3AtLHi+R+lh/3uvGQE7DusKblXKjkr74Cqz8H+bsG8tCVv9C
SR5+bvQV8HBbhkzxrLzYEy2kR1udeJjThhARs8EBMfDGNAEar6XEkfnJmG9l
AJ5eR6dcZIlD9rUylM6sdFt+bN9hpXnTIU68thXiIwYGlj4JGhSnyl6XTLw7
ymrzYAejT09w/84yvc0SdsIM9WH1aYuBatwJ1WhyohczP+i1XY7XlAun4m8B
zxCCC33itULxl4QEhQs6nxD1u7eOZOarUjAPRXRUHey1Ve5o7RyJ/FewdeY9
9M+xafOI177weFOUEFqhrXaH5jO2VTZnJN6goBcyTXOaJSTxkNhf2FFqfzlA
Yp6DaRLeini228GYpSw8yJEYjWTHV0P8RDkPRwiaMeMhn2JoBPz/u2e0cfbZ
dC8njbwZC+w4zvWRFvMLtI+heWXUSZo9lTeH16E8Tnw+7LTkeGxMsdRztXqV
IGUOAP2KwjIXUhMm9mpBwz3cqd/OWticOAWzlhquT3Be8h1wy7/raYkTVao2
IYMlSPb1KIvWAfNveKVTVXpTNKERJ/5UmiC8klXc0Fa9aeqmdUudOVyl5vRn
FxqX0uU0mHaqh46A09Qyb+Lg22o+RWLNOSLhEbAsb0MtzjIxAk1XyOZo8UwV
9w4tRfSlUsu/AMZv5hOzz8Wy4w6DNCN33WtTvpd/JIZtTH+ejCS0jdFEY+qj
HHz8X3Mow4EPNHcPIvENlgXjGXwJN418tOlX0aDZevSb1qr6UtduFh8xZb1V
0MT8NAUPKBv21LdTWGPEQKPgWy5c5YY4KYxyJ4AboO7AkmRgdS4RtU0uNgHZ
PXPflmJU4drNrsd884Q7VzZ4Pa/ZpnIonuh8thLXH1TMLvgGNP36COOC0hX6
E/ruVcSstanhdYGSJSgb6Wc067OzhrYh3HCUzp2HKIyOApTFNWQNZXJLkaAV
AxAp/NMZPgmX6hv9Bssw30kkhzXKHRxqa0cpfIyqndVesn3u1pPp5FTDqR4h
G9gDsSjD3V0c2C/n4PkZsVhEntlg0KH+lISVo5aR/mzv1S9NunBANjX5O701
AZMR9Mcc7w+basPNDiCqE641fhTM4M9LHalS3HhHLt5YqZtRORZsMP8Fypjh
tfA0cacz7gCW59XzMl0w1LE9LZXf2Xl/O4luk273QvaXzB5H2tACe9hshvbC
JhPuYro4VjzhT3FpPyniK2Iu0GlnGhjQ+ECEY6VJgZgvzpmK1XO4hUFiFrbc
dhZ+5Y1ieCUmMaEOZVJ5+hbYnVkYaMmpxI7lFwmYK2EJH6PBfgnOENXwtmVw
+eGO6WIMdqMUOs1Pmz1ez/ziGvwrhu5s98yV4o+BPti6nTO+ewVu8M1wxnTo
gQ55BCABxnqGokEAYGffLBK+3Y2aBrGHT9mmxQjD/Qt5VBoN8spemPArwINM
McyUnos3cBpDY5sMblOnCKoPUrz58tP0kKS+s4z2N+Gd2Xwc8QvNa7w0hIR9
Sdw1OpxcznS6jTTrucHMkrPU8VyXHoY82BqRzULfmG7vQ/L4PdKNK+WeSySH
uCbrAmrRwWfezLz1be8x1oLfGPpp1Slxo0kFEgz6wlDZTIIzL/cZdeBoA/NG
GCkITA1PlLYbVPWIi+QjbruXfA48OtoSrE04NY9Lz/sDRGDBTqGoy8grvvDN
QzK/0sRrbrgyLSRVAX+kekVAjza7hwIldlOBl20fA0qpttWECQYCjeoEWi6D
bbNAIzFBjP1GhB5hRqDqpDlZs/w/Nhh5p0dPAWps8rl3jnlobOA1REHwJrcA
98ytqNr7xL6ZT4FbX0UknWA4wc7UIlwLmo4lJLZKNfexMv8JK5k8w3vxp5fq
9LVix7yY7B6qSCqisaVW0sWCMRg0oiphM8XEp2bpTb0j9bZN7P2yV86tZHnT
b9dd8UUCwM27QeSQV9TJ2dbuXNwoPhGrM2oyJpgnPdYzJLdPfHxlWhX24//V
Q6vH0Ov3u3TrPahGsvjNiByM1oBzlTVj0iAHKuD1rbr9b5S5ZoAqM5lQv368
Ar8EV0SpfFDWB6/2vxYD8t7A4RRjrOZYbkZb4NUvqTvzkoV+3Urz+GNh65Mp
ldF4w56ZGnVBCGL/Ja8EZiIXcahO5ZIcMFlZ18P1cHWdv5J0FzJKd9tTq1Re
ygkOjqnJFrtaMmzPZ/aG1s9fu7PvKbgagL3yBZbj9TmyeWq0unhD6//jxpcU
va1PnwmjjCSey8L4gRMXLzIpvXGQ7Jk8OrQlGnJ5mJrF5xswyEO7Q25wJQ7s
ilvx8xEqPNDBcSeNh3NouB3BhaEcO3CxXddi/lXRHm726RsQUC7zvG9nnROv
h8t077hjaiobHztyNeqsF+VRMk5ExTMPUTmMsyUg1dUn11oGBFadcpvWCEKb
/hQROrEzKNzbtcVifQvG7Gx+fc0rVuAffAz6ybSqff/t7ZMICklCvBj4zz4S
nqpzDjuZTmeNiwFE2K6vshdaD6RzmNiM0DaNNptM5P58p/Szq1gav/i5bpMi
A6Lw+gnqM7kZh4tX4Ycae2iZWwPpNaWIn8G+z7s+gMNyVhoRPbaHCGJS9REB
VEJ61Zc0c65GBAusL7Yp6RqmNMWw22ieTTOn++iKP+WzVKsbVeApW4fpopDO
UGPCD6UuCv6oywicR5KrtSD9NkM+fpcvZSisbyUutptRwsYys74fMZVDT2+i
GfaG2WjJf4FpXV1AmQK+Bd9yKPp8eWZIppQNzfKfa5oH/JkAObJvoP5/KyQI
O2Ay8TkXnTI0SrGH4yGps31FSB25lnFPu/hKqenXrIE8OyeKCWLDbfAs9nf4
YO7PSEUDKv/KhX0yfqwOKNgcCGwc5LYogm8M2In6Xgt7bDpRDXtoKExjhnOT
oDq6ABa+D5vUCw6YRTgK+ny0sZt9bCXgF/8iq6NGJFsEqJQxonzbVz9WccUL
FuIh/7iUlKABW/ZDFE9LR1sDIHeZJhHsf+fVI8vqQ5uZU62aXYajKg+2ofmj
gbL32Lj6EDK+fuZtohA688v6XD4PuL6ldW5elYwuNtPm6tl4cSAlU0+Khr3d
vyQrSTqpmuM3PeyH1ng1CEQUXHikZVG6Zicubi3D3JH7+eXD/5e4IeKTIe2C
M2eqI7CxxNq7gRfdr7KMHhF/ityALB8JQ31XuXrwA4oTCcdIgG8TKWoewxOJ
7Dqf2hUnNZKLagpY4k4T0iT9FW+Sa0BUCiRIhX1daG/kzdxKCzrjWKufl2RH
hjPjCQdS52PC94HKEGqNpHQ5EcIiL3XTfr85f59j6z8SpCMBX49UPW0Es7BT
0/PPRxgbeeDzL9xnbmllM1Pj1zQ9M5t6X5NfeFiu+AwUNagwy6b4HTGKNu2Q
vGDR4vqzngighH8RLiO8HAZu3v9OxZT8TXuw9w6iYcLCGVkuufVOUnDQ7BxQ
rEWW66QLdsck1Uv6BguHpbJtKXpHHcgVTiN2bCzkZoNeRmMHqhH1xOs8o63C
xMqiom8pN5EOz8wwv2DHcjEXj0pYoNbO11WMSHB8eo4+nI1rK9z/il+e+8WM
3kD79U6pQWOYS9fyWPS069ZV5PPZsevwenmLKxHSC1aaZeFXd1YavWM6hIzC
aM7aqOMIiqUl+o4jEbddQDj51Ys38FDR+/yjnBcltfCM7C0M//rgBs4VPUgC
rJTWKVoGGQKsqorqdyBWX/KuQsPSbz5H4B+wqzsiQWpDRC1eUgU//YGWXqp7
pJy7cHcHfXBOU/YfHPgURYBHUxAV6YBzuGTe42xdED/4zXfHvdp8f0W4ceCd
zbE8bXNf7Rt9F2sykKm/1DdN6uBC3SeXL/h7MzcoMnNj6Pg1WhBhWg4/pOm+
qeV2vYVIe29PZGorWeJh34iL4Sc5jVnR8O2rP5MK+SV3+QGgiy3l5HzRpmNC
aJo1aJEHb0tv8V4OozIFVeXVweCjt3mJ/xkQ/QT2ysGJdVA+Cc/icAuTWNS0
JQ/J34+1nLFO4XmnujayRQKJ2pxfwLS6lHdrYpYXdSC7GJdH5C6kz3ac4kms
ox0DNsEOwgBOnotR/McBMI7MYg9eEI3HcAFxwU/tu7EjNAJv0MOlU0RACl1U
U3eAS7WlAAm/3FXZFyLzUvwjx8gtmbtfa2V7tuy9/r9oHCkLi/GMYigpz9aN
R2ZWeDjg5WiWuvAps7AAFkeK8Gl5J+7Q97DsvgRSe8mvNUgY1VaCLzVD6Wag
rwgJ21BVcQvGtWItkU8cnK+aY1LB3X/uVGOO84wtwRHdq4g97/x0uLUfNF27
tnnogEXNysdmy67n/MWxYtFKlScaxRt7BY2uB1WiEk9GzCMmxW6DOPEhBuaN
rNtFfwUw4Rd02gwYSLPkODnQtiP6RbB6OL1gQsFt2IVh2L5ocpgHKsuAIFxW
GF2JPr4+A+oA6+Onm4vOkH2pA9sArIh1nV6yT6hxS2agBNWUlOWBqeAuisPK
/OJmfXgl5tQ059I8FqfLYlMU+fWzMuT8g616wnao9LOmxwFUuOADEOSCAWpB
fs/XkySdkZtCWfH2xjxXb+rPelwcIvf8ZGHmKFEJQ0C1Cqw6aBSr3FOApBg5
PLw35Jq9wWvPCGWtkoe5BfIn0Eb31IjtP/CW+c4gaDzrUu4LpYdK2EZm8Qcg
6cpSIly/Kgdt4vNkxeknAq+nQomAsGoBZFs8yuQjS9gAYHq4dH9lo0CBmC6O
pjfn9Lc3R5mOzy/DLZjLbGOnKma3nRSWoJmQsjQ5NEWUu7A6vSSGO2tZwtPm
qHKHGSBjl9uKZEwEru8P0R2s7EXVs6TuJR2rnGvybp4S0KkNf6oq1Tq4HHGA
wLC3GA1HsqnT28MGqjg/78XsF2N9UX1dqfw+VsvA7cUX1TKwZYN+fxX1rCGN
F1PzRxYJJSvdJFkZcOZZ0Fi3LaT33OQuZ1O0BnzNgx5HwQtko1s4mevLPyZU
hfzTMSmOl3CW9CzHdi91Kw1JwYqPwq7uhJla+blvZDclJ3GRAYL7w6PSSWIU
WOfFiwf76rwzRZ8bWVTCmEcOJJY5sIBYlB3g3G7dnUhUMGvtsfWlqeMaZAK+
gfcvOMiAPLxNXQHGaUY97oHdoAbqBsXc/od3GBEN9M6tvxeK991jkFR5PnIw
QzZOMopNyEo+BiATJ+Cw+4+7GN2aA2Rim/ITfpu/n520G/rOsxtXQxNmzxSh
LY9kwLmW2kk/OASOLtUL1Mf1x6ZHHFqUMsUnwqxbT012DQ27JDJotrN6yQCN
9KBmEtL5zqcRiIwzuUb8jbGNPEs2cF38s8vTSrf6a+XKVO3sOZGXFCcxiaIs
mR3YDUFYdt49LAW9JOofvzySfYhcNHGVb4IpZvUCOMGL7Xy4t/HtO666mAb7
jp2FIgGFZG66iNRw6uaj+BRGDnZLkzECQqfWOMHv17vXf/Kwy193qkKyBxPH
fmBwJsR3P52E0CPWQIkrgE8oseKfRZBYq1L83GaFMVopPTsvryJu/Yh3WwIh
4D8OUxmuTwM4A056k1SGqTIH4KhvalHSrhbf3TIjC2KksA//qkaLw2ihoKfI
PuayX9jiO0aiuAg66AgzFrR3t7uFk4wwpiZiDPtPNU2ObU7/bnDyyu33Wz+e
aItgd9Eocy8vSQs6ltuiZUELDWaei3Qta7dh8yF7TE0YEXbGEGIiRI7ZFt16
OsGZVY5Zidd9XGOuDbBAXvkIr2XK0s/sh311n1MUc3TG4Apu5Br8VlCo2IOM
I4Zs3fnSA1vIlk85QvGtq7r5RecMZLIAHH+jOgc1cnAXX8sFV+NIk/FOMB+8
a4f54cChtB1H7kwNwkvb6NADN0LwfUBfA3cE4SkxpbkE2xDbHFURPRnMX6FB
S5oslNhz+6TglJSjKWOe+bDnWxuJJ1inaZg0RCUA1udBFc+MKdX1iLL461Pl
O9Opo/uRxwh68aEW3adnZLX3ZXDtAG8ZGOAChYq2JCmvtiD5FaPQrq0m05lL
U/sUGOJxg8XD8AzDcaait9rKfqi88A4ohwVVWTC8jo2BBJNzB88uO2YzMAhQ
kh5jmzybFAujKm7jOHERCZz9799GPh3qwD4ClucfJjLt4YlTYI+WHdxLcWX2
W2N/tZydxpFKx1wzVSl4kolyBcAuXmYaKHLqxU091+vC6NHPvlYAUFItrYBZ
SXN+XiZRWvZYjYc/RvHWZI5Ci6EH4VAmeb1B6GTw8r/YiX2Qxab5KZb/B10D
ZiAfML/qAjtS/Vb9rRmu8GF5wHDOrXUcwvO4LLIB4xHmD1MgOlhRuafsud9q
JVzPm6yShuR87KgOwBFH099DlXYZAlf9s9O04cwTuWHGta/wqAxMueNeMai2
bzTWJsOMSrSOtKeUYilkDguWGKNQosTUotQCUuY6GYVXLsxMxHWgzmuTEii5
6cLynelyaMLbtl/wSSrZGIXJiXA5U4ZQd93d7jHb3UfsPWZk4ER15fA8vEwY
BNBdCBqsKY4p/FoDXCMsFauerggWazFrmKDDF/lU+LbFXLdOIuVhmUyQYQHP
qD440d++KH1GjctusToRp1JvxfJDt2F2v3r+8DxuUqG1QKlp8/Pe7McxhD6Y
rYLO6qbTjbZ2nsdg5EehRY7XxYFdkEqACgJRihzYrlODKE+Fn7riLV1j0/YS
luOOXL6Cn9Se0aj6HabS1rKotgjczG7zLywvU0mQyjXjOtDi/sB8fuf7eF8N
zTfq6ug0RPhOCnxirloP9+ryLUtCMkoYE6/8h+QkAd0V6ukFdVbuP/ecVZPa
7ZZPe92eXxTMIdtmtHRYEe+CXFntsQ8LKszFY8sKd59N6nlmfzwDTo9l0UhW
GRCzocyVt1dSngtnMkoWT3ArkudwPeqA52K6rCF4ed35qPYlIH3ZRf1xFaYI
gXSl8cq3hPUpXbWTtuZdvr44n7G5ZzmO2K3vWgtR6NWAFyJIHp4qv6TsT/qI
Do0rjPl25mIQ2fE7oA9OSD8zdaucrvG4H+Hd46MoEU9WxpW+3VflXPUQw4Zi
BnbD8BTb4hXYBz/d09ww9Kt8ijw50BlBR+qPkHVuKtCQJ7WUS0Auyc/M52Or
5617VgrtD+kwgZYI3op/Xh7JELltwhEeRnuv19LoZ+am/wwcxtrGcPPdsGyq
4OSIWX1uJmEncF7eRiCsmK+WPQ4bF74te5Ty467iiXgw69vTEPVlwpCRjJR/
azVJGqkWCkASq5ET/gDruGrGOYDT/TfkvN93kkWWZxD5wHmRD16kNtwsv32X
For4waG1xeTgIWFUNXcExsWB2NrlHRloeYcwddawhQ+tFGP9QyPHJIfTiH8p
kvyiVCzzlFCPUWStjJIfoYBhDHWtDsIU+F0o/th+AdDPMTuK/Re522aobu3O
79BaKValzqbajSSNJvonHZ7LyR74oQfs7Li7PY5+snLUA6W5gmajjC/qklEQ
phitFxwORn5GiUTRF3EdEqynM3QYq5Ub9OpC65FTo+ZstrG/fddluUh9pmit
2WUMqTnCqRukMoi70xs3wKcwPhvFxQchLytIM6xdAY+/vnw0IxH0SmM1CQfo
BI2ZPD3zf5t/f6L7K4q+Suam7z0fePG1CWAkVchHtBotgmG/1t7U4DmrVD8I
e0J+Lq22Rdm5tyigSvDxxb+YQe0pBbdPhWO16A899cYCWyp5ka4OIHlhLxT+
JEktLO7fgHziAlQXy6DrjcZts58zzI7X4u5Zu0nZVocBfopgSfhhA5FvbkIA
D2dH84BdaIu8Y3L9vN7AQYXP2HGUZRenfW4JkDZmBd9I0+UgVn/sE0pddPT0
LRdN57QGXCwBgzdqw8OipSaVp9U2Ng3E7BibaXusCt3nWqBpsjks+IYsAYNS
RI3phyYlaMHDv7o5sEvbtVgfkMEAKn+59mbuYf8NdicHov1S4vK6SrLlQqza
ALXyKh+IajdzPcM03mXczU3yi/nJrzCVI5cRisxY0clDFjiXiSq76A6oDO8N
iehSqqt0tScQJcgniIRE2T8f7QN6xDJPBkoE6xiZAIuAiZxTmE0663CKccdq
l8f+d2Wr2upZDP0h+BVioizkA5mZQOJfILflnUXf0v2Ezr14hr5pg4OTMF/R
Dpgm6nJhEMG9DsLRhcXKKwmncYLexnR8rZ0gfmWSt661XHuDGvXPJtWPLzTf
zKYru/VFtdNz9BhxAp6lvz6CZetJhUa/ku3g+IyVvKrY/im6yz8duMCp6a2W
O+9PkrA95p5VhntPeyI2v0L4BamTLTQX6c973u3+GV1Y/KkAZWVoLRXbcpXU
EbszrvzX71WvKPx8Lc2wZwJ0SrQecDpbSIswWqAS7Q6gDcHE7mriJCKLsgw2
ibpqkWNkwvb3dk18l/QIaBXQca7ham2/U0uTIdRuMpet6AWsrftRbG2aTVzd
n3dA9K3ZqzMEhHiShVGyb9sDOwZjrSZ9O6eJu4bi5cM8L94OCWq64+g2ZQQ3
LWjmpEKrzvozq3rpKaVCcEPU1+UR8RBnvg5VzNFyukWps6EkOl+3XXoiJfgU
kQfR8IEOVx7EXHhj/TT0/j6PKAlim/9BmCwxqjjyn5tGZHSU8Cftmj+jSHhs
sUYzgehLwxXbBjDDj+6rqooiFGwRM6FHCAhx5MWMMvv0N2p/kRcHLjjRXGoC
ZNykLgJTpoGm2YziHHVE9Awl5Eb2tFW41uH/GCuFupQfS1rNSJZh7WWVDQZ2
SQcThDNMZk0QRJ8WON8U/YuW9UQTNhIJz7HiMs1SnV33uDWbaNe4V9Eau3hP
xI7YRbqEUXatPIhRU8WPOO8q58ioWLMAqMAm91FhyaijKsdu2jEXTuLGRNTC
uMjoWd5UqZp1q9e4+pNSY6wPrdkH+F5+hFDH42WSXVoCgYisRU82AB3fMvf2
Bls4O6m7UtJcgIJhiBSlDo0w2V6DSaI2/1RGlAvglOP4cIbKqAhRqE4fjjHp
FXpWH0LDC7Xl439Oz+mJ2S3KaPofN5ngGVsQl5kywDq9VnibkRIrsmPlwzL6
HNGF356QRBViN3VOQe9FHXhfWOrj8WO6TUKhFC5CdoyigQg5OGebSDzeH+kM
3WevRubJZFLGbMSWm5Fnv0ls/ggJvqCaJuhwTfU28rKFwOFnPYdMfoFCmiid
G3x7tz8qcLELQR6RHV3LBy679clUv3UGeWW16miVykXC98tjBRMWcJwMj0PA
47trLTBeTqshDVX7ybsWwXGQK+5wTFDJs2uW6cE8zCPibr7PToyvZGeTKULI
G3majgCHEz+2FJMGIsioY7GB9TAyHV/ymSwcQcR0Dw3Vwyk9aT4peyroxc/7
FKflWyHoqDjr531Gu65TTHOBSszwOe9h726pgDqiQem1JS5j+2vj2c50siMW
PtsPqZROh4tn2LlYHvyfwFQYISO99TkQfCboHkoYFjj7WZ+T5dvrKtCDvn6r
qUx1qct/LjWfzd5evzGpngJuirwXPMMdd7L6sbqN/RlbjMa841z0xktyLIZk
+mT53XkIEtY6WmFLqW7J94he7XPJWzdwtUNoN4zPH41gh64tWflnDD2c5aLu
5PR+v+4wEiLZk6uITMagsxvlAyF5uPX3nvwVTmcTJQ7O0ZKyC8/DjwhsaWd+
DFZSdRAPnV31hdUknzkeH3xSvt4mqFvF/y37O5pCUZaQg0r0m4R5195VyEL6
fidMwqgC1uSSVYwaDVeZyWFBYeVn6znUvVWxAdOZRSDlUbz0n1GoQzNI7WLU
67yFoyVNOEEHwFVZA95j/tbN9O+5Cy15Kq3zG0zFMH8lS0p5oR+4HLqA201w
yl5BVcu9lf8zlSBQwyfagZnwYaltIyuBlxWl4k6YUKwYHFjPcBzUFA+xFeNS
INN9J0zTpn7gJqPlUKwunDbWifGxB25bzYfyV6HGbjwtC3RbC/9Sx8/0jxQg
rzdCCoa5v7nmQc27Abs/dXfBwRqOli+tvObUIHLGB0ORfK1mt6pQuCBTXbA7
U1xsDSvzhRqsLtKMteuuyN1jSZloxvvVIXY462cxIGTvj8RflxJDwuP3KekB
P51YEv4xj1lKlFYVruAoFCf85/SoSrkzZZURocFaNDBpWr4D8N+tsVO72tF8
NQO4X/NI7istOBYti+CRZ0/a/ZeJfbeJADBxdAOONaMqmphwDvekBKwLCtJl
yC6ksw3amc5yBVV/AlKq4npkUw9VTGQErynSotm0U7B7LVe2iCb8/F4QiB8w
bO1mtFB2UdONhudh/UyLUmOg8kX9mac6I03lirr4ESItICZe9Tk0UPnaCKKw
eIhNEMZNcwmqLV479WhRDU/5F9BzzISLQnmdajMihC0nKZasusaTq6UlkaEh
8yt6AQ44tYqC4p/ZAlL460iYwgto7lQCpqLVXNBm812ax0fS+Mj3MzySJ0Qk
vtaasKthqN27HHknFxILjNC0S2QvlKEWAX4nk3v+72mK0lmlZp1x6VdwO2qm
QpApHvxhXoVbu66J66FbLX5+3P54Pl0DWA9wt0BXN4yZGtadlQ5y+duwFTfu
+TlnEu0Vi4OKC37WRyPHSavKSJf1SWz+VioNYfCzV5vdnlggVlKoTwV4LsL3
50hV4RBDe0bgATl/uT2yWro8cb8guKl5wM8HkbwcERho0rjCOYscYEgWn8iv
YvA5kZCNKGRlq41shdo8Nn3W2F3PCAkMec0fmQkNnRMBudxDanKEpnU2v5hV
lxVo0pwJmN8/Yfv9YFJIR8f2Jo+vcCVN+VxZ0c/oy6et1JzdvG3nSK6cah90
7yLcTp4/0ZVBhpDlUdaAiCmn3Gt+FbrZLx/dA7MtfRmXMwSHT2sL4pWZf6lD
cPj8/c6pZ/+GbSHhQR4YglgwK0xERmSmDB115Ov7u5umV+GkNO+dFSINgk5T
lOz23zjsNhUhiR7fvoK2hqoG4ZlzZEm0AiAz8xiWzrXn3Z6eQ9tSVpoTL7gm
RmJj7Jku8Y4bEcoELP747d7JoPI8F60OipJHdTTY7GpJXtjRgdrvnlJIe4MV
ztNbkoEQd+ZubLf+VAJf4U2OCPY1hREqvdSBXp+IgqjygKlvGNCUn0Rt7ikw
I1x8ThBq9AMvjfJUURBVBpvLnHo4+o0mgAyNcmwt7QNIzWc+BDWygGNBNkwT
WwCNdXZu2bdGPrCh3K7G4TBbwShthEz9mLRdbmrnSTKZIcmOr+s8aSKDmm6/
bvKkcp52rGbCW+ORNmdC8s7BbDIXhX1NtgHoBm4aiydjTG0T9aTaBxJA4dbl
Yr0xJNyXogi94DDoFa534HCSah2Pmt9vXydnXDgSt0Mw3UEQchc+kYydWy0i
kBY+xTG+1+EcWIBYDUm1ePtrrsllH72J27qkKG3go8a9dU8XY18wVzhLzeTn
+MFOUF4RwgqfRXbpFwq8a26Ex7AMzY47URnbKQwfNvkmfUOfjXmhgSjcKTFj
OlETWSDg59vbApNvWVh4tXoXf710Hp/UVIKi7kRNLKmeL9bm24SQcDOiXVta
GpaInGl1jPxeBwaXdsXsixY/dITgUvQNQDi36g/fdq3WHh4EsDKpCFG4EugF
5RJ5BMcLUoAcYQGc6iiM0xxf9YLpvZHIJN+1zqe0hoX3ri/yZU9PGYRUg2XQ
y45SL1AAyYd/L697RHR4AjFmQ1typx/KpuIhym+0DWnDJC7Q0ES5NvPHgkEH
fklKPCk/2oxBmP3ye8V+DmAyf5TguIViBYgcg476UAUPfq2g0kS5Ol9Ow1pD
M5mCb9qLq2ggeDonRyGKN6mkmqcRCRstBUIoUFnJ3hG2h04pXJFMKOkvdoG3
QZRzuD9MdrVYuWaotQlBEnfftwTbpqvPHzjCrNo+Cf2yC4OmsbIQ5TFTrzv8
M6OBFjiAY9ua11NnJsUJ1pEr9laBR9zE3W6664+Yxd+F4NWCYZXF7ZpvQS9I
EyZWKb1wWuv6aqAwyv3DlSz+6GdxBwDnMrW5dyf74t5/Kbr3lcf8UsiGkKsd
aoluzmsdP1CrGrPPIkeShJoRtzRvj6nm3PqrK26YCBIWhPdiK8IeewiLB+6v
3lZnoxS30m7e9dt5OuToF2bwts7+6hIUfsNuf6RG27ighj5xJN5Q5684wQhM
L4RPjTNYfZ3lyV3Rw9OR3neYIP8X0q34V7ha9G0TtjHY1WphlQhSYm24S8wA
OP3Hy2djm9g1rv/S+0GkUzUp5m4+NGBVGcw+efJ7Dk5sYx/p7Iw25kmTnUOo
DMvNn1+CoiCLPqCJXHqW3LsZiCZ5kCYKDvS4Sn3Gk39IeZzyYYsq6uMlo6e4
ZdGEnAR80hF3DFUfkxFUSIsxnSS4dF9mubeXczBUS76/myxzi5xWkm0nRq9H
EAGS/9ca3PZHTv9+nEZxm/Z1MMNWITQTlwNLtO2gXd8rlNnFv/sqbEx7yT+Z
gzp2TPpkbOZHrawT5M3SLbCnsZwsnVeu6R/tliftAwl0GEzF+aF4WS5gDR2A
6mSgQaZmojzXJ54aLST1GOTjFdUW0IKNAj/Wf+TQGuaKDo+edIPvIdIh6YEo
XL/keP59CxYv18ZST/JCckfEACKeUGjoR0x9JL3t4INQAbKXtCUGxlmh39Sd
/y9IX+w7n6lAsCSzjHEYdgKR4oZnuCWJghIasVh5m0mUij0i7GBA3wCisEhm
gAGNdAH1x++V8U7Li7XRV5THGPSI3DYmKR4FPHyM9qLlTIzEVdKzYka3kvph
NjTI6lB9HhRk0zM3AOVJWEOMZ+gZDKsgbKystonv4tCHFWkcIPAfRht3Zvxp
LwIhY/WbK9X77RRx/6kKeUmMwTRzkiQ8Bq1cUvONoKDQDYEURHzwFNha12I2
m6KQu4lQVI5A/Xh9zQIWh0Eqi1p+V/3rqdzQX5E3sM28JPOomNp+JaBnUvce
Z8LxPEEbXDcyglCYoo9YyTPq+dHYJhGxWv8MZbHlrsSMO7UytwHGPzMyMU4P
VyjxlTpOAOEFY8i054bUesMaKGQMHLvRyFaXVwwg/TjamjD3j1uBWDN0Rtw3
jczROFFqZZJ06V258njWEhCc9YYaaZPzeQub7TyekWKWsUYxvjYxanuXGdWz
0kAXD7An0ihQEazr+8zd0Muh3A1500C6kYETmD8VKZYoPeFy4q/3MWhidx8H
bw4XxSWZ0L/aGSnv27WvEvL+FuyDjqVx4D81zItcmPdUEtGz6byx1p3FRmE/
uA6aPiatpMJehbUQlaJ90pomiFaeApwSGCr105PqLNzxD8MVP4BjWuYRUpMu
GsTxsNjIy03kULRZxNc4EkApWpKDTwNjykGOSTqTdJlSTlvi1OW+TTW6oy3s
bU8xfkT3lFoQZ3FgPatG4waXjX1cLh/Ir2qkOtpMwKderM7GYcyxggCy2qkb
fkq4NY0G5Z7Pa4t68BRTk5oNX0sv71qr+YUNMeazyQ69wWLzn0kxGLTAIGJQ
keCe01DvN3AAoWXAnVP8P6dE2pnJko9TP3U9hohGbALvGLHIAu6Wb2U92Tht
/FP7LbChFQq4eEL3U93Zlw2HQ721zgJuwpIrRn20MWKqeY/SulSsVZA8eCHT
uKouiaUM6jhmHh7igkX2XOP4BxD0JB8XiLjV1carvBSBUqoXNn0HriNKosry
xmTHBxfHSFbHXWszhnZiV0khwZGmw667GPKJDfie58z02LYTR9Qo0Y0OiNw4
lNa2lF26zZ75b+03xChbO9ofiNFSsZniym9w/VRs8VpoPXFaD8vtfZN3rbHw
AgeEWs51Cfb6OB/zLyjq28UwFg8aebBmPWtPooV08ycuJCmwKc2SDkZJFXVY
Hx6BC3gn5e1smSI4qtlvXgX74FOeZm/6wt7zZW2bBPkyunSXWwzcSrBs19mJ
d4YDb1Y7mWL3JOaofNxnfSXBTy5RoV5+0ARF4PG94q5K8p88PB9ujuIO1+oO
YRRyVhSiNqkAtGUJfDrp/er3ygXqqB80i72Ro9+XqhnbacY2qLbq8AJYS7i+
RMfMkMfTWtRQUbB1qc8KMI/m+2nkXxetQbfq6aNw6CT9/66f8nz3Dsk21Hfh
gn3PUJRbx1K8MCk1/kYfaBFkJ9a/1FgOV3FIgTdJKSJXmz/YToKV8kpL16DP
0vjwXjxmPSVmo2TXWBUL4ZmyIBXewba8VdPvcT9lAk4cfEWI3igZ+oJbqKiK
atbKTjgTDbx6fexQhToFd2dU2cHRe+2EdokDH8z2GPPHqNDFH71KJRlmcesB
LdJhCuDYLs+rUHoGsTIuXCUoOHYWx2IxZRJidriYTLfUPJ7UpWBmKtFF5KlL
Gqnc2UpsRKn2j8c+H2ylr+7KIwIusf1Cv2tfMeavepJ7gF4Nag4SbYyVHaT6
zWrEqSA2a7JbVh1XiTfOrA8/kEEITJpEFSE0IUv9R2s5FJS1f2+M8AQ6wX0V
FOt9NFS3X00lf/dBI8eheStSG1aamx1Q2945TtPSVlcr8xnxqHpoRqvKIB0h
Aw+qA0R3R8DGk4Kyq8fFEySaNdcc/tJGeiqrgTmqzBduGW9rD/mKPI1OgI2+
aMkOZ5aJZsMYixZCkQUemnn9kbe5Jx6K59J7+0J0z5PeMhEUs8ysJfY0Cl66
2fOcVB0oEnjEtIMf6vZLgZ9WJAItQ+XhtFaK7KfZM8uw2oRHfMArleHReynN
MBF5mRS52hEwPXYbKNjelVwqWm/6Lv5Qpf3bM5FLxDT/LjrnzJ5ORnueNBf5
t1RTmV/1pFQmFuFJq0lR8VLk6VFx5dDxZIQpDi9LBbLrrHr/mo5MFt8CpNvB
uMCBjZ7NLs++hvOlukrmckZada9qtMX8mtLyvafYikn4HndYucWV9X+CrVHK
T7+5Jx3La3Wk85mogEDG953hVRt4KqXPLXITZHTvbAv5GtThbo71OauWAj2s
UE+SiMsYRqoKAuidx6USwePt3XZThg/7VIkSOXBI3+9QpdrzVF12I7/LOE6y
KvU7DUbiOD1sg1Fp28ZACARzX3SX9Q02fJ+6Yg22IMtNeKs6E+QBMUkWHx5K
chcipYMjX72nXZXiHGvTmvH3pNKPFXl67IlY6SLU4n/jkMp3K5hcD6WUIS3n
QqgPSLYpO9wyoa33DThbCgcIUC0BSk6Mjh2EsrTqSxyUSxiKPrqUa0x2xVpt
9B99LMtFY0PB+CizBsMSfuGGdLUcwi/DcHQNSM/j5Y30VXdVSo3s4RhFqnD9
AlUPhKQHeU8zGFTqnGH18J6fMaSncXUCcsDz30jCxybG17b8JAfdXRfI3xaL
J2+86g6dxykliv4/XM2SCGcnSjAB6uff2z1Pf35OMNNRjfY3J2fxQG/4rKvl
ARN5GeE68008QmcuGjpr1tvLvwxnZxoPBfzOE+Ag3B8UvtbDWwSHyeqK76Bi
DsrwUkRDr//i+acSi2/A3ulfZCNfXRTSbYMYylgEWU8qJ1pfMhTzVZ/77M76
lZNeb0Qyic/A5KJruBjLXzBmDFhYbgbY6mXYolPOf+BnOu4OlDs0Y0HzYe+N
a/YkIbu2hDnTcwIwKIjgbtZbdnvjhFyzR8N88tKUrLVXLY+5I9dQecA097u8
xjE4A8TKK9zPauhOx3O6WhULsAsxbCEOgBw4t4cXiEVOekRI41DTC1sTS/Ri
BNkkd8v7ySgihlgZfMGhxKg5OxU9yYJa5tDTb+4TYf7phejDGWGYWsjpfAM/
W2ZMI261oyIfanG0/4dJMWNxbPR/h5r0fSm9AUDJZKTy775B/ZrJ16P6hNlj
ftKJv33iNPnl0bilh/qfy9NC6dNSQp4KD3YD2pvvMek9/dK4cjxO/x/zoc+n
F50OIHlSuNl9nUbNpXohXu/ldSXxDy+JwAhEuQhYQqtDqUFuNDFOK21LHiBf
Eoj080IV6oJod6zAoJmHvTivkwDIIMIdORnvyGKuqJGXPAqbv/xPEaD+xcQ3
Axy1Gvj7fMoiNYdI+0lJT/bbNvnVRZBdvFSIr+GkE0RRsSVxXoMo0e8OYHUn
n2LwD2YQz7fCcN3rdOJJM5MCF7LbwG80j4C1U3FGkUZwv5bU9k764lCep+zK
H4xaZjk5u2MDf0Ysd55DAXy4HJJn1blc9O+UYle4sFe1H2vOrUIYSPcP8N6V
KBV0ObXfZ+bpGXOi2nhjXamtt080rZtukwjq2RdbBFwjvIgL/7tt4vIAHcYh
PUcjUKywQwLl4LiWMDFeYK8OFT6r6wxnMiIbXQZ3ZPrZmqhE9gnPkPXS/vD1
8XkgCj72C6qO4uJZhbGT8Cxaeaa/al1Y0BsQVsEQJC9nP29gyZjDhHvXSZei
XmVdbfKQdbGowgVFRYmiWhfSKWHNdlLsiCePlZ48ty/t/ct+b8nv/xQ7BzcJ
PFhLeYjJibw5QcjC799OTOAfIEhEwfSDsi9287A4QWo4EQEDF21XZ+Y8iLY/
+NpNhPOU42qVvVKKmF+kVBp05wAW5yCAV8gXim5J6LUBZV3fjacvgVTMSsXJ
GU0dGSsOZInEwJ3QkQhD2Ta6IFYJUEBj+qfoRcUSOBcU0D/nQzv6ttEiJS9f
adlGsCOskYYHCGXwetzIavvDzy3xH3xLiNkf6BpOpnueXhxn3Zcn1tHscbHp
pJMtAaT/cx3kv+Qk2gDT8ipQVcWN1TxKlzg7dfckz98Flnw97Wca0WEOWp7l
0s8xOSCnQzj8gXhfoXI8p/mtDJuz9fNkgVwbdrD3wg04F5CPT40N8+s5/Xbc
fuVfaeymFpsXun9w3plFJeyHM2iBRH8tC5ixmx01KISO/P5Q4QmDRl1PfGRP
ZxfQGPmjW2TGjnR1ZICzX39iWebdTzdHEWAgB5MgPd7LZfjDUIrz5LZXcVtV
lb89+F+qEuxP+TLPYrdz0PCOLGzp0iqFajpDwLdKa/2RI118ktHYfvW1pEb0
JvzRLee0rRKJY7KAmZxUAs4/1AbROHjFAGi/qWqJANMx2QPsLnpkiJMdm4Ss
dUwXWWgSEmssTorKSXew/hzjvtIuE5Pxwnq7xVUAMwkT2s5faCuJGHLbfhIZ
G5U35Aj3pZua3CFN0cZKJR3u43K6guGyg96cFf/+XORBFeYDNADUOH9Crae2
Ca/bPIKpvSfhXN6QJF5CnbvUBi5O/DKc2RITE6mlZhZqPUmoObl2IFXi8ifF
DBR6x6nAYzMqwF3s3OZ5VL2kr8GiGZy7TRNcm+Czpbby5gsUhbTFU/KSb6uy
XbCHN3ilH52GBNLsGtVMMvxiCZ9vtQOGdB+CxNHfuW74aAAPKU3TfkmpM4vE
QEaECb86hS0oX0Lb9brKkuBHRK0SLbxUTgC6WH1JUC0cfx8+VnAqUxogoahh
0oUkY7TsmS54eWSBDht7HGsrsdNu60zoE3wDAZ/tB66/hnNGnw2/PHEWxudk
9tTSnuo8nesY/Qeo44/anqXb3oSxG0V0EW2Mf+OyLpfKGqxNdXHzJpHFalKV
l7eGlCxo7r8/kj7gYKIupjllMiTb9bCepntuShxAwWK8kQU57wbNqVrNT6WS
tA79usXz54eOjANf+NCg1Tw1hX7QlyZg7KJZW4pJvwWgg0kx2vwUpQ3R+HFK
onMLvwM7a/FkVhsajn4O2cU8mzEtU4WHXZPOk7OEykHhxJuOrn9X3h9JdgXF
senUXNByxp5qRToSXiby+sI2kecSlvJ8F6ASUM3N1jx39OTu6KXtV1Q/w9fj
NKvgBqOhhCtI9GHEtf2/6+HASrWBAoCnVJ2FrqTFAUGuwhjYTcGc+/vQGtMN
MeLAFeGiQ6uT5XUlEHvVxBD4o56AtPOqilhjtaiUleaysrIL8L/15Rd5tPgT
gCh8/MmtgCu9Tg7Y0F8xIURzzGQXvdBuptukGUJ4r78zvq+b7dpvoZvOzNTf
ac7CnwRkMPGXXEDLfp1lxURYRTrIqHau2dLcfLWjqboy7ETrSLZTVS4m8Kvi
w96ZhMP8/KBubTXJ5xWNlyNlnILGFtJP/s3abvBBuapY4PADJsvSMfv7g5gs
1rCRn+NJyZu3ytHBrrd/clu8/AzMCFlO61YvV8D4qYQ5/cgsFCJv0UNLKjx1
JY8ZBIFcofGB+YTeglFbsHEWB/o6F8tbOMwJdPIQxu1RrOqK6oSy9i6toO2u
Y2GdwOdtWGDac9IS51KC6Avik5IoQr603XJ96uAiOR36tYIpItqS/Zq46yuZ
fxecUzul7lfDuB+L6ZzrdyCvS/vpywQHQrtCezYq47GaFH1PJCnrA79ckK7o
dAEIQnOIOgVPk+uf0Uf9/Mg9O+eXG6Y/E3EezgX4nRjM0tOTLh8Z6OPi6hdh
CEHg1cTsesN3zmaS9f4TyrkEytHAz93vozd6Jxd63z+WooI7Ffxeg83fh9kT
FUp+rhuSx7M2fmhHL+sEu5X+mi6hjuN8qACUNEKCXcjpbuhKmizp2z/1HEpX
eAB5/sJzLmwsNzIYnqikE6l+b2+SPS9eBdlzgR87EvpEigvdXJYYsOjZO6e1
8CjYiu/QWXkuVZnWdzOYWqsyKe0K74k3WFrgmsbWIRdyQMJIrj5AcpSJw4Kr
nqz8eJ6WzjQOkHxaSYRdeP1U1j/HY6MENuuAwhWtG/YVjuUo0W6ZLMmvr1x+
jYhqFJarmm7o7Np+Ow2MTkOclHlwjyMAYEiv5WlHfbzxYHRvJS0kEvZZEyYG
/k8NWsmhM7MykTyTiYRdiZzNSuma8sVtJl2pPBW5DngyIBx+GVkk4QgwRnSt
kxG6CdTgi2pmBceBWsX4AuVmpIvu4H5VmlZAboWe3CTfbbNu7zAFR/tvAOcX
PHfKpz1WskILq3eHxoW4RDYWX/8OY/+Rul63+hjhPC75z3DJ05jPwssc+tej
N190HlgMtKFo1WvFBY0bcKbD/Ed5nNkNkh5GHjYqCSJ+N3rprJU9ILqQTYkB
07IrZ/uEn3bPp5pBEqcO9ZicvAyy1VeqWVra4LcHw0m+jgxEcwkcY/KpgUW2
JLFUi/lWGC3bYcfDNI0oSR9wHC83krDFS6pkzRH8JxM4E7anqTKiCmYDiLeR
9DU0n8BK1KXk9czlomYpNzsrPLWeZ2JdH51P1KrDBzCHMCtJT/K2XAfvhthG
zC5oBJcp52rMvB2WJ6VvZcsNj7VksD4YYtgMesdKaMJ1zpZVgKaDNrixKV/w
4KSQjflyc9cDmS+q1b1IcwwVvKYzg8uRb7fCdHdBBbjgwn/NGKYvaCGnxQDL
tXO60VAYpDbCEOlOOyldwMhga1j17sQX71/RGJ+ggUEK6C4vhhSq0WIPwVxs
GrBT4EUhExJOEj37apD2fHAV+eeKi0phhbCHlcaPyNKb4490jyN7IdQZLjUa
1ADYoA/PXfEC9in4Es7TW6RRRiCZNBWemT7nKp+A9SazwA91U9qCJ1TkkLWl
ASIS4Vbhp2rniba+H0XXMXjMJIZ52/vDrkwlfrr3jaSK51B3rAOJ8Mg52h8H
p3UJJ1k4WMbaYw0xBCacwKmcxI0k+8Gi227yX+0qYpx6IQ3qTQ6NHMpocBJl
i5nT6Q5HdRtVd0KoTwY4uXmT399BVgs2/uzhH7UBrFMGeS8wrb0hQ0xjaH3e
FJrYURxePEre2WRHNQX9I/D5rWZV2qSuCaXSUfEl3OJJOT7tu4Xn/tZ68uPR
ZM5nxjlkXltPsRNvPtWA6SLzxjo+04Mxd5N77cRauxxjx8CpKvChrDGQAgt1
OhChPJMTCBvPwsCGxECCvkePGSfEcQN2BDuG8p8+upQldOxlPB0aYW94Tqw9
IcPvVYENGbZicHnwlLr5idAbVhEiJq/g3vnqRihLlOhvoyx3xp/6CNR5AXn9
CT9xKm/6C1F/OnkruzGw86jLia2Vx09ooo0G3xpJ3+eGmynKSqlKJRet0Cu+
KFYNW502BxVr6VgUN2Y3ldBZ8fwKLNOPlPHXTvn7ptAQd6zZSKWPhWuR9tZ2
pUDol49y+71yL1Mm0qMKKZEEzn/tiyZo7CwLz++4eHGoLbB7AKASl0l4fpcY
c6c8fjC1YJFmUIVdgEY1X7HgLvkD/f0RtFVI/nCgNyFHX5vStssBloZdg96K
IgIuYDmTjVVkLaNag22wAFPlv0Ot+KprV1IhSkoXtYdkSCq3dwZlPAsRKIy/
rmE0USGNPXpWlVo5wvnCQBBtbpNFV88a8resVWZ3zdi8LcI5qK/3gOdmr/ly
di7c+te17OXF+f25sdMr0uVC2I6goq/MOG/CaBqN8TjU5+NVeT+DFSBQ+6lE
5VSvx5tuQ9EZlUi9YS5PoCfv9CAlZNo1IvqrPbfnVvt34g4t7ibOzBIShvDx
IgoFJhY2EAlzTT3EoSD/wIIzJoHT9snRWH//3lRzye2rywuwxJm81OeZSrib
tlhagHKKZjj482hiHkzvFvHOC3IQXRqspiGEsh9uoeNQA+OkIIArJLb90hgx
/qTvdekHdFGR222FIcJAMysEfI8gPRPHrzPwREbfPMBIpiOOV/Tc4GMYR08u
PXvFVOLFe4MyHP/x2/HXbyesb3JHLl2x2APcL27ha6R8ykxDAq6UuMKxRX7n
E30w1sj0w2jBeu0sF8E6dV9VS38A9C+sgPRzpEAqb0eamyAfyxcaEmsYnT+N
0w3C4WKtyNHkba5mEVREqf2mZ5EatF7pDnfRDrODgzjgVVbbywi7qJ2XvIVi
59b6JokRBe8SfuyEnFpMC6ZGdji6wjBEUK0msjuxO/AIUOkX4+6ruXWEn+qZ
4JEoLtEOjyVRdv8Xhq2gYX46QiIT3zxTBaanhg3FeUe41bX6vN/EAYU9ERms
rECJ1MVkwadWe26pEPhklAyuUFDjhi43PS7n9jxmkrcnNGMpPfaDyzV09jBU
VzPHkU8iYXuxLgPN54KpwEZltC3HXVN6sV0Geas6YL5eFGZwgdEandZ3nfL5
5FmGJDnniBOH6SGD5EQZ/uc8tW9O08ziL2rw+e7dz+QGc6ZKIOcpiEqY01gd
h3NnXWX9N5OGidULbUfWPTnYOV5d45zsgoRUKBb1zI9hEEglHLnPZm4gIR+x
H3WMC/GhcibeQCk5ipxp3/X4lIX90kpn3fqDoSMOBMF1bjqq27H/BTOJ06h/
6mD3sthzSy2/6b2GtvMQC+Rp8Ghb0UAZrMM8UOPeG6RbIDK0TxhG6cMixUH0
u68k+WZZvYApiTX088HmsR0hllhDSfdcRBh30e7npzl3EjrGdWQbeYDPhlNv
2pLWPl5BpPs3GQiXGQoNNunm84obR/Qw3DUunUOvf2kKIJCr3oPG/0uLRT9q
HbBnjViX0nX89qYBt5uMVpH/Txm2lpjCRnvB+mDfMAH85J3kWlPJhzzQjafn
FNrXW3Tna4DuIorC2kmGqE5Lb5GyVmofryCarf/odrCEdC1LmpEEv+iBC+pW
IjjQa/1GhtGpAZYb6Al8N5Ki9Etc8Nt50iSQ97oVYaoUFgS43ojyqNSBHFIb
1f4+CQhJWFYzkcX42uJyPK/6vGhlz/vS0NWkxfNGA+k56iJO/elT25JkDYzz
5H/ksSOu6dkdB5uqHKULq8UFsOV10/p02xFQcc05Cvg58htBFYR7rlqsyMmi
jEmUju4bThRqw+VaFBWm3cY/Bd5DnT78eaNLwGXLuWdLHA1WyHctuyrdG5CD
bc9xPBnZKOjRj3vT060WmsDG1pq2Jvx+EDTYt2sUHWTowaD3+5KYEGALx7S3
h7NPBoU1mBl6KTRLsrXwFTYDJCM/R676WFeS7F+PF+bYzO/Pevqo1JwXwOLr
mWK+F3EYGbGsoD0jrUF+KBDCuQIT0qZOBHTuSAA3VNqDijQtT0oAGkhUIeot
LbaDB7sBIHFOG+g973AptovWvtD7b6C6Y60QSPXdh9T1XvM/6h6gwY8+1GGW
pSo4HzyiqsKdr7R1LuN/St6kntuBUjipiU9IrJB68oM0bnOeVB5ktsrpnwAs
OCjlVwy5sR1isNxXQCxndlE8q/I2tGpSJvR0nh6ujcFTxfBuOk0fJP/ckOgc
GQO3nQMU/ZBWLzMoj3osZFKXlsXASvm8pWOHk+FwxqBLGTNfNofEQOrHM0K7
PGfxLosSUwbKhelzpvyckq+t+1FUu+KCc3v97vAFhfLIYBFtyeMlNMHMuDEN
lcrV4N2XZSFDUjPdq+unOodEeF9xqhcszxghXCU7SkqnbMnh9JfB+MjoxM32
glZQFeLL59lo9yv1DK0imE+f5b1vBX/iE9wDa7up7UQ2zHVwMzSA92254KfW
4eo/QX4xgCJpIYXhEe7CeHzQV4OjjKEThud6nLFCeZNBBIdgo/7Er4r6tsMO
ZJQ1DgNH6zUoebHLJ5/IvC3mjbMnfJ6qf3ZJh8WEiBQwPQuKEoiogtnOkL9b
CrvmPWxxVUNSpyRaPlAQfIJysCXBDDkB4taEspBDefYjAE9+ksIE25xT+0sw
/qiOQqhOZ0FRIMc3U7R5sW+hrW5V1uB3g0WP1MOvP3o6xMf1ShD6muVVF39y
py7DERmIk9HT/XB1PaiAivmvkVZSrKEqYjhDuaYl4B9/i0mO1aRgvdtY44nL
ZNauBXZIfOFF7xrAMBgstF6rmcY1KVCq5FVI4Tpa6+AQwRpTmruwuzZjv0ju
/N+4rOutctdFKAo/BYHmjJYpCcvPhENZPonw6DdKe2h4Vowc1LSTd515pbCa
2f0YOquA6zqZE+Wr6gwF8HrDzUhS8V8F+xM83w64RSXqAWx2t2uyDx5zXqyb
hQjZenxzzWzyIYiXTM8u8oCuKMhOlQmW2i/+1RN0hk8wKJ+O4S79M1dnQWG1
/2CPKMKrqVX7EBbq3xNspGBeZMqCS3urL2S7UDmacL3yxBnt4r42cXeR/YI7
dGzufX6AA7UY79pzY9ejH3YdC0cu1svjhPvrOJVGeci8XshB+hvDQwK+cfyS
YQ4sJzuOcWqEys/7Te1BuBduVigQfeQQzWwXaDxguhTB0JtYtqNHCat7JoYD
zpoOcQL3bJ8HhXewLx7r/6mRyRDUiA47eP5EExX6HW/cniDlAz+J7JB2jBRM
CPaiIuTxRwSVxvsd3j19PobGiWiDjOGcvFSbwFwoX3jcojzBiHPpjIMlZl+6
MGJsLjOfjHK0aOe+L7eOHzLeZdSutejlVFwpV7e5YZObSmzNQWuVWRfwqg2b
iVf6SAGv+WooN42e2Eus4VsoVhig2X5mxBL3+5too+bEcf7YeCDCeYjmCpwB
bpE1T/vbQjVYvSPj6GgELaWurIrfB8c5lLqvKULNm+QnbqP2GqH4q/5PHZRo
d35NiNyBspGIH+RiAoX5RNt8HES+iWLJM2vTq6BHbEJoMAYTiyquYvVUJ0CF
3+9MnL+RlwU6SYFWqPuNvfQeQ1vsghvCo/w0/dI2p3UNjDbshRdIwQ+Hc0U3
yf9vHuuh7UfBVnD8dddz6cdHvuo8wwudHqIQIP1u05hhRrrgtUU4X38W5gLe
d/jn8TGJwjGIzxFvjgetL/mztNkaE6cRF0A4dBJ04I44rnwzntRp0XIjgk9r
jVDQHpzlB2nHft/Il8losLXokT5CSzVFHN2ubgcD1qbKOYRmxUMWHKwXkk1U
H2HrhD0c3AhXpnYgfqwAXetOmPS0PQtKXNT+V4slDHP8xo4SyvILkN9b5snj
+1gKkYE4hqN+XfeGllPX9AAbc+TiMahWA+ftSy/4bzw/LOUvsmbP+wtISjql
tZ8JuJI0dNWiZpdmg87efjGCKx6vVnhDzlvt4rDaxgVUU1WIIdVPW7I+mzOW
FYk8yyPAbOaKbFYkVYXzkQ4wtjqu1Tf1w4vfWvSSk6Jlxe5HXsrjj2Z4tG4M
287nx8sn24et3+fUyrafCG2+d7IMhpho7KK1v53D8jVTHTXYsjy23T+2v+lc
BG61u5Ubumr+J/gmsux3SVNErzG2MyLmDCEIOW2WUBjTctDF4TRB/l7j7E7l
zHqKB01Y95lxmFrIVdWW8YhJTf8cg6+a0iO3NlDoyBqZPn3wXfJYH2fsjj4B
tptKQ41c1Sh/klD6QMIwAyxwf3vm0MP8D3QmOTLL1E7IpXrGVeISLf6mRl2+
QBg6rifcjYxlEuZXBAcG+00qDeoBQ3sPqTEabTBG+D9ysK6r50AzcLh2gTHM
ZpSw3TJiNJwJp7ahorPDtPWfdPoAs/5VZn4vQtLID7bIlV+6qLLE8pomyLmg
3xoVG0Gs/arWlrQxFXFOHJ7QzZXXFi/lVXaSCVbEtNarjh63YsTJ/fXyDYnG
bNR7aktf10vBsXZ0g8RMrsV4YSH+a1mmP6LJ8kH/eYeI2XfrPorlr3QFKcRX
lfZEX0kgeTilLS8ReqNDE8rjP0Xy/YO7NAMCP1povqOgSirMFHZbVlBfGXCf
QzPulaG0vN+l56O4t7t776tChDDd6XbFRcbHwlDuMH2mM1LL4aE1caHclamy
ZpdVHHw9BVItOeCIOg77Upvrkrn54Jt7aDvOMKvEA5BnBsGTXFlcXkm/VihO
OW2+mvnWQ6AU52mXH4Al5YN1dyDjfhPNqHEfDAaepO8DoW+ZNlv7P08Q/FvV
GetCiQ0Hz2fVG5gVHIUwmlEdfwN4nntPqybX9uvWvo8/ZCIa5Xt8vNssR+tb
7HUBtiZ5g9B8epbBiN34F0F2Aqw2NumEUrBCcuzw/2VMh8IolWmzO7r3B4Ur
Kz6DpGcbGcIjtYxXb/4PWNidK5vDIK2sskvk12NnH6lCk9KVxNBwAOaKIb6p
j1l/F1PAYZvyEt7qfI5km4LcVPTUA+bwcZ8S+MzpvuZwU03ywSgodxD6GcB1
T2pb+p1tBl8ino5bPWPpdUXuO3nQhShZgauVuSCYK6EuddMCXZYemAmCXxVJ
5xtCaWeoRX3UuAGoXFLnWtISW5IAOdora4YH+s4S/pNEbwtxwpUedhqBdeBG
wo0Js2nSMPBsFRQEmNTA243EOfY73F3A5zdUUR823/gWw06wm9fS76VyELbT
UBE+OOLgw3+Lb/miqItVaSMD4IUXu/Z/PDUis3Oh+96guxJwLfpyfWFm+rpH
erhzqMxXYU36uAb3ICN4lJErFAFBOFXGfc80fjgtQC7xly8TBGCMJvgskZ3n
zzA1V2rxD0OxOtgXq9x6xVwwCJfsT34Hmf4GgSSFiDzDBH71zEP30lQbIhhe
+lmiaBSea5rhFGmpBAXQoPsztdCJfRI08lBtHSsV1KHsVGMjNgQmU1ST6thq
w0ZUkX654fuKuiA3a+AgsOUXa17E4yghVID/xmcN781bG+7rVZjzgXTnwP52
SNeH9P8y7zrY9ZT0lBnjsy2QSjl/j+SLiMTR4LB+j4qn5ScAXadS2zqFr51c
ReqKtUcPaRel27+zw9gVlY3DZT0BiRUJgUQAXgPU2ZcVq9wTuZf0lB8XTU9S
S4GJUyLNt/Xs63WZUSWBhdo4j8zssa78Qhc6sQ8DF76Sjt4ZZquG/nDvkZvP
E/PtFqVxBo0jZJDClh0OP7FosbmiPjb4UzbYItLP5EzFNW61vALJSn3bfGdz
JyLjsN2uOgLOCivS7mqtpZR1DFhnoaAJapBdPCAL6y+6PdGuCw52/fhZv5dB
c+iRiZcvJOQUrgVaMsXpfZmiSJVqGOgeBtp1QadArvL+Z+cwRVyE+NSca/Ug
V6sLiwPJCOEPTf0+xaI0TgS9I6Xn199ODVLcVbLH3DyTd6B0+t95uaLa9GN+
Npex8jPESc7V4W1g4nRuhr1bbd/zHLajsytr4OJJL4REJQAZpimVR2gnNamd
0oxroie7uUWHNPgKvO5n4HlmtoyJdM+zT4imUHbL9YA8Ye5p7aG3r4sW2q9T
TJ6Q4yEM+Og+9/WqwJBKwNXLlrDtOsqS+u3wco9CGskd6Z3eo5FDMxEYyv55
uVRa/A8lc0etZDfUlAZ8C7eiPeS00I/0dhISBU9Vq7btgi2ReygjGTSyzskE
uffJRQ6UuDRGQ8rITsaSAf3kpZyh5I1Jn/0kPAFCQLQ3q/a2PNmm1EKnjEeh
nUdMKLsj7D4EaiKhQbL9OTtM9N9xqz8cS2QiYEE4NTtrkF+EWSVzrhk1Bdt0
ZN3HEBxwLaH02fxMAwjghcnErf2i/7Px3lcRyRqK6/zKSd7tdCOTlNP5sS+N
uc/wfskgj3kCrBPZrM+D0UgV/0U7Tn/q4s8RHPPGCebdMM1XltBptQJlRF+l
lJLNJP2lH4xwucWYlE6u2Hl+4/C85F4/NivDAO/JPbqnoT7p7KND6g1sSpzL
Xzph4f6QRAE27WZAqhRABiYbTcbVRqEuTXFpOaLFBTVvUGQJ4bJ1Uk4z6OrY
ChnWKoq83+51ifRpvo8dwww1LO3xghIzpvSWyErQvQd6SvoGS+HvW5C4BDyq
f9/XWbCgEswxd57TSZqWfYDugRKNQmguhpFT1Rt4p9q1/to8yLPoOyrtds4z
GDmEgpsYUfYR8ff9r2hpAlWUkYqEYbtUpAPpDYUOxHStHfV/Hjl5gI8fOFSg
n9mzzHNz6SNR4yv0HgkO4nRZVyA0Ao36y9kpqakaoPz+H1fcTjIII2IsdxHl
NlQs+38GSzixo96wiJ4BlkMgJ2HBzAphRG5uP/n9h7TuKfbGLnc+XD42Xaib
arkRk3ctNB81nWsaemmz1QVlU90EOCPMLzJIUS+wMZp+lgamxV37zKHlVYmW
1kUHxNyruREklCxRB45i7tMz/Djpj0/STa7xoh2qolqZjtY3HlA6FYY98dYh
9WLD0yRAK+8PLi1Z5Tqho2l3EHJSJyO+IzKB74JRkuRi6QvkxtEah0RmntM9
xFdykySnYfpgxAsSM8sx721VRFOBHDaTD8qLMmGQHvgtv9rDH+OsogHp42PM
w4Q9xwx+2lxiotl3ZY3o9pXdaMojgygDnGWwmjqXM3RImmdBgPzk865HF6w3
d5Lr+A5pM1mA57t5bDTN+Ij+3ZPKvHgIoAvyj9F0kIDwatO5FUc5Q0spJogL
N0KplmyPy/0iQ3j9A3oD+NPHa8aF2ax1ESKPD8X4SB++15UrxnpSOtAFPHOo
0OvuqDpBQ+kwPd32l7RIe/M1F2rPRiGh7V9rrjRtf6/0QBwUQiGqZOrihbVD
3b8RPc7Ora3FtaYhG0K8nbykYLxM1YWx8TY8tDj8bxEViRdzX4CS/ieHSqxt
SdxvDj4uohzbW7bLGdicjMP2FPEfEkg44pRKJE0w1jfNq5aAG3XN6VGYQIC+
n7YzVnVlfMAiEOqimGENdaBsQDzTsMOxm2vU3FRLv3xZcYodnPwGH8MxasSP
gNBw76n9qnMBHeAlmCgd0+N03XxUDZxXakvGVeX4XVXBXg5EQSsfMSEpT6c2
Dr08XTU7trGxHg/5beV6KD+Pe7/6ygEhRWtf6/8DqYRORqP5zyhrmFuYkufi
QbJvI0pqaVIHMbLByQD+42NeytYPB//ddFxq4Dm9C1Z+9UYIduS1Yr6wb5hW
c+ezBra+ZxCZs8UcdMJb+Qfo1U5GC0f6WRM2SfmJ9mqu4UY4lRTQuU4xq9xH
/DtzWluiqELRutd98/ubX7GDtgkxW8V+dVjamtL4r+iAJMTRa+7EnFgwuuNm
kkfuLGUTIyJ6fvtr7XW6Im8wSOXdI/WiXa1rGZ69yTQI90umynlDV/mADMuz
PjtWRHGI0qJnjZIec/d3wDhgpj8RSIu0RVc+DSnTY1C8WQHJov+3CXK+0nW9
WtTm1TjWV+ab1N/aOs0ZcT/tAf8JAhpZz3aJBmVmcsxqZkxKxuO5KgSVSK5i
CvTkz01RBDY8zw5cIW6vBzLL9kyd/fvd3IMGhNJ6oAdev7taQaGZOw7GSlD3
6kT0igcNyiURHy+O08XNo6+R8DTq5H6FqJJpGgRWxS5Lv+vUWIZ5gdWaOAhu
zsqBgrBCnBmQbial+Gfxz4fyppDQixN87ISVTlYq7OKSP/YNb9AR/Sl+BcA8
2yWQMDID9tFRhwxRJTc2fCycB8XTQhYLJhoM/RLHG20UZ/tDjNVtrDYe1UJ5
qTSxajru2a4W7GqxcGpCg0JeMBUCRYovGo2QJPgcpa0/mDjXhSqX1VMyRDd6
ybh2yychMmv4TQWBv43UY/+vjLhVgaRPQInn2TKVEGSX4ekPAwvU/7SyFDu7
TQAngq8nB7VpzOXME9Wck7JgpMWKAiobXsg/qtzLYxPUqyuxUi1c35F9EcDH
0sk43Y3RVJOt2Sr6sbFzt0oS3TTTQmNRHVUMnV+XpUrA01ZvUMS26HHzm7Uv
dNTLhEUu4gQIrBYYNs+4aBhV9rqwbjZNo/rdcA/PXLakkfTfEKat32VVVDm4
wxyD1+WdwyAQ4FKhqpDjK2g3aEBjzaQul6XMe1s3130TZ9PgHI4ZF0PvGb93
u6fDUBGx7SnFj5dJF+lclCIk7FTK7d8IXW1CbDSeZmroov6K2QSea9YtgQzd
mHR2wwMQ4trV4LnKkUcBiIQb6ubh4fNVs+eOBmFwUbRH3EdMOLDAMGOXwz/r
iDu5f8ILTxGKk6rxltp4x/MPMkYhqM5GNHYO1+Xb1TM6FGYvngI+I6JcL6bT
NLCSRm0JA7mYt62RsAnKNYltDIWgXsYRfxbYBCPP0EL1UmZ5b4amWSHhH7+V
Vma3XzLHOJiiVPGDsEFSHAw/8nP6oAqJBj7SwEGoYC6g/xk8rcfNtc6v81ZM
ehwyLGKDbZNWiB7KZjhW9bi1vLk196GonJk6C9EaiZDl77tzuOIQ5IWZ+Q20
+trekS3qxVojKRc0FjlePGh2wF2IFCm0zSjQLPebQlmHIvwIbwCuJf8Rr32p
fApncBsy2MG5vOcRNw4qSVTWdLvBQgXEao77/Lq3lAaOmK5ZjdaYifz/Ohyh
KHURLxCIYjxyCSsmwxIU7/3f/168T5svQUdF5hAyFU3eJ5kP5hAqOv1dgMU5
LpnAER3nsMl5LS3aNoAKLbqw33ogn6U/rKUNs0kwe8DDEnMUgY9AWr+VHCcS
KTcM9D9IYYVyZPY5vb7Ur4uwgyEgH7nmdrJDSA/pqH/vQJydE6wPQzSK1QOB
FuwEtOYCNwHKveLHEeuVgihFbmLr5IaqQJXVi7dZrBSG6RIXMymxVJy8dPDa
Tj2J8hKazoMsc9NT84MtpqYJf2Iwd35m4r9HF2dhM4CWiIyn66N5UEB/+1OR
SB12xrA1wfRaJKJLSSn4A6/X51zhHVD+fIxvpUfiqC7uXSrabkq4miFM0yIx
yhB9zD/U+P/DEP2hEdXJk/zarAKqGZi+lE6iyW+Vsekatwnie33fhKCIUsGQ
nD2thxahP0SiG36ujlaGcDbSiAMlsQIksNj7yCnmpQ6Q8FgqLTzjTtRsd3ND
/bcg+UnGTfDaiPRlAc7jZhadpirCdVkHGH7ZeYOKwlex7w6z2dSZzmO/xRib
QLUMmg8Ff9Egk7pDR6OyVlR12/dcthNwTQ3v6LUFPy+j62Gi81u4bJJbelHu
uvLaqoMdoWT1gIMUjynGXAPXEXttD1KC1FdLffHuRbz4iGXEqI81FsKjfodo
v6eNSapDYkZ+MsN/uIucCVAh3UmKnLEiiomZIeClTS9bX78iCEambjqg0k//
Fsl+luTXNkK5Wq4yE3hHLpU6GOSWNPJQQFKni5sR7CeLweTW9iefOkj7nhIZ
dhbZ6j228Btwn/nk+r4mIvKCauhSDFk9UgvQuxs6jHFYJcb0lmFYZUv7AWiA
FL1LiJVcDAwM3cOaIEMWzRNrv+i82M0xbPe80NiWkdLTvDpFIW2YTDH4GNuG
miU2lZdDjuiyaax4ITui3IJr/PIhaZdSE0PxV8eI/3nDknh6KYReraPVvdKC
Yi6HGpkpcGEeTkFFgnZO6Iy3ISEmbT14loEMFT6DnX0wNQavOJKKmAXIR6N6
tBxV0XZeTtRT5ni9EOsojPuS1eTUek/DcGm52RFgiUUcBxHC1gCa+2uzrWMr
gDblCDGNz1M8b39Mn0C3JBRIxhjRL7U557A01QokcmiK4t65/7xtkxPuPCIS
E2NNbxuUeU2G3okwes8kYH9qWafQ5fbZ5jbpMZUYN1XTfP3LcifEHodsfCMQ
Zxjzsj4/KujXyA7aeTUwQXjogNJSmHTu0YzTnf3JSfA1dKyennpj4A53oQWB
9oZ8tbgke7LrPeKzsa0TvdICUq6GhbiDxuD+glA3+z1DMMjsOauwgjO24Q1F
/aPae/A2z76gu4bGMXZh//HlXZI803Efj4xHTTMgm2NJFiC+BafVjGbdtuKx
08TBJ5H7+CMP4sJu5lsU2eXSPTqM56E59gNCbD9J+A6CNplomF25TT7caaQH
mOWzEXyV0lyknkOiR75sAninF/ZBhgmVUuKgJ+yNyxtvVGMMYdTEt1RTmPxg
0YX+nP6ecABQGfrAQBHJKgMVDCRQ6Rg2A2qK3p2QQiGNCLCOKnWwyI6G6RhM
5xfFpBRSYRspe92fp0oQdpHxx9vfgBwlu37tAy2VAiZdHhYiRjpmw9tlZN2x
GmTI1xZhvrngyPr8xFdznrlngO3Ywe8pW+PRD6bCNNLviPjTXwWgUWPb8kij
hyGrpKmo+5VmSJSKyg/27TyoEZH/bQNUbY6YOKeCJQN25cCtad2Y4SRHwPqu
DmAZVr8pqOfOoz+ha4wHeH6a6CBZvYpHfN2ixHbdPkgh+cX1m0vaqDKKzDrt
pThSAXxUUCygFIJ7lknWFIYsJUdjwamf6vBzopxMNtT2pGFEse+djT7rY0Xz
Ni1BjB1F1HlYGacNrWvnIz6dPftiIxeb4ubzqRbleZRZaL/EFkrBxFy6i8aE
Xtsc6KWHU/Z8bQdglDgZwVPMQN/IBArQbhJzI9nP//mKhy6rLhDrx226dW6t
/KSnqnlzmfTuIGKdtZqWFV5X8KPlm1z6gQ0oa3KNmUjtz/GDLKga8oV7j458
vYPTeSfTBLmS8p+Bz9X4xDvP8u1WM4t8wofz5UkuN4YTgFz1MMk6Lsakh9X4
i6JU/RB8AdoiFkvbDWXTieJGnetWaGp8GadWPL5JChAo+bTsjopPSVQambyL
WX9DOvnyx0kEoUZXQOIsZrZFqOKUdhEzkrXonJlvLBBllP+hurZyT4bCUri1
nR5gIKhRPqmH+OMdogTCJqRs7nyffFukZmNzc36fofHFN13giWmuahWKfB1b
ix9ql+0HQQmt8KjpVTmq47UaDNSsH1ntVrZjnjWgpTcGS2dbotsml7XB18nJ
LL2/NMwEeiz756Kq0BELpkjUuczh9IMEuUpr7NvQOccUe4/+g8PhAVOn6QSB
5XTz6VxaEtq53I5EE8wSvtPGWjGVE+8b5yE+jeN0S9ZvLQ2NenPF1y6IJY+F
WJyS7fJAAdz1yBmZrOBJzHTjl5LBOsM/t23kT5ccLbUt/wlynrDFs5o/CCdO
5SvnT/BY+bZriXMTeY3oa88+M4gZYxEUgqp6PREuQ2MOwFTvZ2pJfwHwuRnH
mxJXAVp+f0EvAxc5+t7jnkLVbqBwFdJMGQbaH6reY9vdqbeg+xp7xXTrul82
4WDq6eDvVKfPVZv+HSGiMQsRA+ae9rbvztlYcWOwuomNlCabpjtgwjfuQW1M
eyYR5jqYWi3CWRPbRMd3+wpFY04JA2IOkno0VYYrKYldWx+o81YGNyAqlZHF
dkfyOOz8THAt+KH4k48NsQO3Mh8D7fwofJ8mslYz3FvzPgEjW2Ny89UMeESS
Id2KSsMMs5VC0gc00+nGXSsJiD8UEkeybwYKPQbE08XAX7ZyOOBxy4bSh2FJ
GWoVNO7EP7tr0fd5B/RES7w979gkc6zXNwoloPgCYL4OTNahfAscn6jVRx1f
p2GO0EC01kD85nq3TqSlYrI3RyXpuXNFtOJx85j68gETi8u0yJBIiYTa5cp+
68e4SRqIOATV/eBvSU8GOVeEugwLA/UHy8oO0H+3+ZIOOWLc8sMnVw8jJPhr
Wm4M2IHosQv1W07064lBCeZ8cuipZETVGAe0OobefJ+/yO/mrUwjWVQb09cJ
e6G1FJ5UaIutu7XN+8ZTOgrVfIxEhQMP6tx33bvuFSp4ref8BTOG6Zcgco6w
njgcBKsgrC3NZVgxYI2xHayZzofOUkKwKNOHknkO6RND5kXBzUWatnQmyO5q
AVjJ9rI24bc2WGkh0KPwa2LXTNsVh50ECQD49+uxTfSkjklOjLMqCD3nFvvX
NhgMiLk//Z8LaeLEeOoAJjwu4H5SXnbxZUSnRPKXNGtLExtY2fyofUZxMyTz
FlxNLjtvcaJAfMpgE6wrOa4BgnQmBDva9kaH/R9y1hXY62P4PtawEGTMhiWh
XDi0N/URy7oDaHzSb/G0Yc99QP3UckKOi8sEoLIqnYZ+qAYUmpk4/8ksj+FN
53rmgBv/+TZFIRPlD8TepNOUvPS2zJ3b4zl4UOBcvuP9dU8ou1xl/opy7lzK
a2yS//6VdYuMmnfr+OEXi7tTlnH3cJKyF4IHxU+ByFJnAII9KH/fBqcf3Eg6
pTQTZUgqxXUfz0TPVbOf+LH/t14TGUGCyCkeTOV0WEzFJarSk+JXHGrK6gay
eb7aPiJx70R27aIoP2GOh4y51ui8/bX22RNvEKXbRfZsP0JpzGsQANld8rm5
IDKk3BD/iDqH/0nea/W+u29agE1CDxA8XNpsl6u5xMeItagOpBIFfUyfmXcG
0spEE0gTONvanrIo7Eg6Ro1LoU9ewzTFsMRAOLnRV7CWy1faYXwdrmRklHKx
qLC7hIRJJvdDKs7d6dHt/3xwP1Uvz8PLRctm4/fiBac/Y9GyvYBP2HMUjqAb
AbCxUD3Q7i+Uc5zk3Epxav7dhufirtHFwqtIqqxrutgoVqZkN7hX72VhwnLc
GwwPLjgdTRQsWvD3JnPGR8oYousQ/6FZckvJ8aV9Cd6QhAVX77cSkiaPuMer
s0eDhkWu19KadRjmRGokfeLInoIILpjdATb7aIadWjcL6Bf3aN1yFQFjczIP
5NGSvE1ZxIXdnWCkjpvcnyNkONxYxq2ne/34wJh+25vNZVt9tFMFXCs+lImi
ti+UHylFyiGP5BRLPEQJ2hZ1cFFS3hhFsWYTEWQXYHaiUlNKQIPFLQeH6rvC
L5xjseXfBgeJGa3i67akOMwXWaoxf3Znytxy0gHDprbPHnX/NDq/lXPSTP5E
bPzmT0U+jHnQzYBy6snZFh46f2hMdJ8rjpK6n0uCgQgfiznqnA88eopFcWly
KJy+hz+pDSfKwtHDHYjIoivUYUNadXDnC1aCiJBmMXcQyGX31w1rHwO4PLC8
Mg5cKmitXL7kzlj6adDQuwDdZ1O4FRNFK+RWPRWOWV910EavvGJAIa2MHAUZ
qSafo+4wnAU5vN9TR2eGX8xWBDKPib2+XyZKHDSfYS33F5g6Pc4d5E0kub+u
T5+AvU7FDLUUJv/doUoTv5jTavtGlR6otH0d+yx/ecXytVxrNnoZxrcnnwz5
BtNusjm8gSxThlnTiyBGjY/xuVhLPj/SrAF6g1QzLFYdp5x9uMFgiHMahQ+k
as4R2I0ZySqqwCE6n91tbPB6nSAFgpjxBzMy0TzBfIhMCEpPoFPDZ9cs7NCF
liFHRxW/I4a85qn0v1WFFsDlwjUlI2+urgLrrnCYAtZdz/P5MAXlTaq4rQ/S
oDaiOGmJwn4YVc4xGu3k8eBlfj0OPGqa8ZEO7gNiSeX84jhkhjtbw9DxevZk
fBt32Tln4h6t3+4yY27kRydQPmfE+EGpcuZT/AiYWM2aSWC1lhd2UNwrlve4
DlARAvLxBXDJ/jnStqWOt3SOAM8wJHwu8kyuyXuQhKdcCoWeal6u+hAIu9vT
VHtE2iQcZZA4/Vm0tR5+h2PVrLjEJtMmF7m1WcGxzeDX9g4P5T4OYFZ7PcxG
F2uEJ/QqboFPx325VXxVfLzGWoG6oP4diw39Y2msbpwruErNUfRjBYldEI5R
fyyUcTFngk/ABqIGytMsIAdGQVxaArVX/1dFkE90C4ABo7GScxptFxgSXVfZ
yklHq54x2wUezaNsokBHiEnJYn+xrHd+I5eCCjVAFQmppYEk0uVJl6/BfuZ1
mXcHWjSmek/cUhqmEXSCMgBaE7BQ9OWuvxxM1ZBqT9RUOGlJ2QIqyP9WN1mm
wRnT9oB2G36l09epNBS35AL+wda8V0HNiMcnV15vThsIS/RoviS+f+EP9rh+
5Yl0L3vMMLpaYkfBBBkNca1k1t+OJLePnOHkZ1wH0HDDYL2Rova1NkwW7P4z
0KSWWRsemZYIoAIahMsXxwV+D3F4uh1nB6JifCflkUGKI3UxtfuTOhMd20X6
Q1Deqr0jHbOhYITeHUynyOGVYkHR4nNfrEryVPvLHq4RNqviWT/mMeC6DwyA
9txZowC9HXqSSsqq/Xp7BBpTidEEPlMNqzXnIuipbRhnBJEPcpI5ab6fET3c
brsNJSZgZud5sDUdv91YaDG/tJc7+UNudr/ocZjNqJJelw3y/79HmNeTcDdO
2R/3pOYxzzxdj9Qgzv9aI9pTtm8X/NLk3N3YFLCoF1Qb9kR+Rt7n5P1MzlwR
+q43cZZQRSwCbOYQ65kTzi+fwqdRabixho2hkrd7r0t5osN55m2tjO9VgXhP
svVDAbLvwn6CXNbdR+NdYaeJKUmL2+iZLwKegnfs7yLJfiQ4wirR+cjpaCha
UmbwF6BjepQdOk0kpGRJBdUUPQpLghmxPbUnPc/KOBXNE/Kn/9QLIzgyme0g
F1j2BTpMmPUa6pJrNRNA33FFHziWU4Vj7BCprPKg/YiyBcvfg4919IRv3T2b
play8cAGy0R0/ZfvlXU7MEqCcXlu+2wv5jVwEJBtic6T1I1N2qAPSEX3p5d2
mj/dK+cgQ0e2yp5sSi4Ts6j4R7T1ZstagVNjMcCwNhLvhQcQNq2Hlc2vWYVe
t4Op9LQFucZUs9KiapHgkOa68jeF36/blORUyOidgOstiXeD7HeolrxIA3az
Mwd6D6KZfwLx0PhGw66xgouqVyNRIOSFUjw0oZhXzJSJ9iUpQ2EsfFb6Tr8C
TiP+7BgOhiO2jnghtBuubhrJ3Hz7PezhUYux/lY5gKzd53QiYt36hB/M65yg
iy1hYl96gcJUerYkiY2UDJ84mWb758sDyZTzIefEBnu7QuY7xQOrZhqXSHfL
QuYBr631/+QTiPxE13hs3bXFDuWnp8aWjHUa25dTdwICEO9ZLH/9A2kzl7aH
N7tXTVB6VfaBzVH1bGke6l9n+m/547wnuSYIbfXgiyqluDTUgeMkqJ+/ElrH
66M+xrg0vKyvd6ylpw0ETfXs+v2KJeKPjHFAAMl0st+LR0jnVyYt3Z3rn+HE
j0PrYOFa6AZ9gaBvC87C9IH7gh3ZOv0mf1b/8YhFbQfsbkLL5q0Nve8IKZ5L
8i2JyGJpg1d7ciJX+VvHOKrI5/qid2hqwRMuQAx7lXaUqQChp8eTxWXTupB2
unEqVDcDayDgq8zpy0OVvAbiiJhHIWe1/rRtzywf8Qn5g9vHlssxdI7Slvx3
xlRuUOvUYl11xxxNki00XLiXcRAWpYhACOJ0Da9F7Ninfl+ikiL8kKiNLFLa
7K7lBF2Z6Dc/KckRS/UwPe+st+TVO2gFwxgvamgyJFkUjwzOenj9ZED+eg2U
C4CnkpwHjL9vLiTz7ypht/5IO+In95Ogf6RIjsSGP4qBgBm9T9RsUbI2iFL9
3jA3IP4jzSukaU0WKX7OxS7/hmyA5y2DGoWCQ0267nZcEWHJLpg3Bw4IBI10
mUwWEJKtnQDBcTw8QZ6St5/e58A1Nh1SxdckRIf8bLrEbdSm3EymybnnCBdA
Eo1CDkEL9L6rDZMFyBOx130WdO9Z8s3qe0nBMT2pk7k0Cn5j0ZMQZEkxM/TR
BEadLCfH8HeHFWpPXG50209f+m287kd1wmSPM0dxGS5kWwgvhCUuDwuDYsKo
qRJpIHgV1c2u2ZOlh8Pu6LApBiaFkx8tPgYJ/LaY1ydRQtNy0XFGHsKUm+1O
zihR9h9QQY4kSSmSZ49qJng2ggq/qjsITu14YKCpM/4Z4UGyqXAgsdn+WhG7
vlJfLLfCXF6+Ah/fugVuB3tCz0suzKsFretbFtvPbdCiHGvoWT22nclzvrCn
qwARHJf48T2//QctfQ/3xIVFK1zmaXc5LvBC4dYBasaQQ8fHNotTvGgoFHNu
tHpATDMXlNw080ee6CL6FQNpe06KDVG2E84iTr/JbPIDJQIvQIwkOeuziTXr
c3diaj2vrgOWFuOE5YVthhof1g9h5FZzS955Ow2v3BY4gSa11TcQ3Tx8Facu
XzaEMXfPtvQSJkv3wC8A8SJvAqO70J+Z2vNG2nJMvO/mN5XXgDQmmEXI6PaD
D1D0FOdPoKr714+6Wq8xAuJKUr8zV442RvLeIQ7mQ2hWSEFEP/COfctKwict
XCBJLtH1p+3h8NxBU95lmNWsXt213p6K1O6dwKEVuiQ/ybjkKgvuaKcp0TY6
KhePd58ZY0L70el+J7Y/PUW7BL8Ccq+oAIXMbI0urpHF1A5YlLloR2ce14oO
pS5+Up7q3vgDfKVp4xopEnT7BxIqrEMH0gIy5Wgxq0WBJveY00A3YjKwh0iZ
NVkmNV/UUi3TlOIBdjH1QEZO7VujNfmMH/kbtbY6eJIYdZtldIAT0J8+gwXy
7/XX0Y4cWoWJHdowrmC/b/oscxCmSarkpBL0U7O6wNDHO7tNpV1T109Aeysi
HE+b9RyJNFj7K6pyOA/Tr8wn/6zGE1YXuaJyKQuNwbrQYn/NpZv0Nchgb9x8
7lJz5yetI2eiW9f73q3KQibkVVDE0rb+wkQqV0yivVEn2yr4GFfeAv2QPnax
lMLvaEKwglvQNvu+lpkfJQON9/po0EsfQMyYtL43Iy02BCkMg9rQ1JEMMdJb
AL3QjQeJJFbm4CezHjLxblC0O3wD+i7druLWT71rS1SmEk8EHSzsEwsKRjpr
EOEZyvE4mNb1Ug9gZsuGHcGyEgBLlIzVP+4g0OEV/TlVaY50XMVJ24+9yEe0
BxGqS62JvE8E1IiMRDywpg+hdnzeprA/LLyWUfDAQZb2pY2D6B4Kg+Oy+Alg
y0Sk98FoRtn5qTiRhf7XNeFFtUX3aiYoSz++KNwvfWWCNZ2jQ6U7x0OTF3VA
QPBuS6G0kdCEvYlPo2kd5otGq1r5W5qqwoVSRYTeHnDbU0S47xogSuMyNmJK
yS4Lafq0Oa4BxzK0tc9oUpqsQVH9NrWTxotnN9S2S9bCE64CJwDq7wMYNa0e
CadSoks/vKpQScyF1sp0QKpx2XKtGqbOlnusIChVyZQ6l19r3FUaum+0T6HM
NX99kGpXjsvPESQZzkj6gfVqXSd54PesFv3ZompGbONJ5dIOEgcCDWJP2OrV
yn+qRTkfwHT2g8reBbcBA7iXL+CEru1sdcD71i5gE8TIxBx73oXwouQGcVQN
NLwdSj6mCfGyP8kqHQGxizWxtyD2eB1mamiSx4xvMHZ/NuMnBBUGrqwJKGTs
tg3ok+HeRuS0N6C8CmTzaEhSah80e1al6E3LT6cUCHXK7T95cNJ/Wu1eLfeK
yks4bMJ1LCpcybCDmlCPrTUJTSICaMb5TXkbanjhsT/H1+gErJMvRud40Oo/
U4H5m+75LnBzV9JyVufs0ROiM+1fdVlIyGuw5RtDK1mWO52JOQm/EeXXkJal
o8DGUBIvyL0wTr/Fv48X4EJC33/40LiAjFOMVFIsYJopZmCtDjt2MKLJ4wS1
iMGjWJ492I+MnetIQ8l6rXrhVsHVTSwnWeACIOuCT0ZD+HecafcnX62F5BH8
t4bpliU70CS5mj8oLKpBl+yI4wDBUVSXacaPAdTojLlDL5cAy7Rf71gSFMKq
Pvs7331e9U6iqVMK/p7rwqmC7ekASolfYopWW7Tu6tPMGT1nniM1XNUP4wCV
Mgby4A5vLvFY/OsrguK1bEgvPO4gXPJSElRFayZCN5u27zm0by68PSV58j0h
hi9wA+10ve6aiS0td7cl/rPt0HAsTLRGsvFOYNhbvuvtUbmq3sNfLmIjUCM8
m++ZflIvs4CtdsSYn5oEM347ZAprv/JQpF3vnQo2KtN2xDvwTkVS9pT5/oXp
bSjppm2Yx+EVjhHCk0w4bmZJABRhpCJCNSkSCcc4zG9m9xraEsT3BQKrxyZC
56GM/qHW52mDfPBWN3jjtTg2TtcjMpgTdPnTBNXGCBiQTMmuEXlf4xLnMdSW
x2db0iR7k89jzDiRy0QFwV+VO0hH8VKRFLX0Oqp4T7NqMqyItSnpCOc0VbCa
sGIbZ2VBfQdt7H4PsJaVSTGMlvvcpNvveR34skoCVEi6sjlqiop3jtFSibbq
TSmKAScpt9jzU/EzFcCKOQajn3+zurQrSDG+80CSJrhzAs8vkR2kB8VDqTQi
UVarWXxoEnYDElwtP1wr2lZB3oLP93bJ66Dh4K3UUUBJp6tjYNmh7EHqCw6s
v/1fK+JVAFui6blPy84BzSDQiZtpYov0q+XkvL+ixr/yLKrodXnmDneXcZDZ
AYSwxD0fvFCbwSA9GCyyxZZvVRJzKNE6cH2QMbdCGo+jy4xWuxQ9LCEcJv1F
jysfoYqE9tFLkfr0+NVy7ofMez7VARQioWxw0wtYJ3Lo1QYbuPNPTMILA6Yf
XxD8wBYExeQUIvhQu7P7kk7OYXuywLqYSckPuh4iyn6jagtdPQ9W6Uyc3ExB
/vXPzXYnLVBZEkX7sPa0tvYPKeZbqghOrZEJaDP5CoXl/gvTvmGIYPv+HNCH
8j/sdlPyYrzYEBCzIct0+VIPCgeEhUs30brbikODbHd8OmRJO6xnOtoTpf1e
fP7F7/1YJStVs8qyTX7YGpEgtfp7g+gUFQcJm85N8/e40aj5ZgEzHFTwnT42
ZYx+ET1kTvS9eaapOPz7j0hGheo0hjnqSPIpxY9vnAGtIgSDdMpcMsF+mllk
2j2Hydjjpk9Wn/3lfPAB3oUtiYivn5wtpjvRBD1NA8EdYkdZtQKzUE1L7ziN
61OoOcaDzPxxXPvcEBWJg3Vf5fUFZc4MJH2E/OWOSYGm+8vlAkdxsKutuzOR
PIC5bCxV2OxcaO6vjB6Oq92x4ssJfOvaiULu7lL7Sw71di5llvqVVVZw/4+I
0h1AHCBwTB4MyexxFGxyitmOvThwvSihiLTVLG9rOqK9VoRyyUt9wM4ThLif
bhY7lR8w6QiQ7GBspYwcm4WPzckZDG198+VKsyJSxjyqcRpER/tt8dvNEaO9
mQp0/dZDM4EwW1fXsrG/TK0bb4/FOozCgzvQQM0+iq5zRUwHMg6nf0GuqSvN
J3xqAz1J1LncBuVmXMOb5XjVzTApo5uhPBoP0dLAtEhi8moaptBhmcKLCGoK
z8CD3/oHwnvzWQoKcugUyCeiMvcJWE9El2qslX+SbTIsYKs3MTy+MpUbLOlv
Insd2IiOZRVKTY1o40ozTYMIda1E/o4eoO0Bs0kPsOn5qxbY8/RGpiBT+5tm
ereRTqv/FcLA7kxFZyEqiJWqxypseJuc/ZMcTvbQgpLbbjd6ftgpw0Zx9P+x
6kecg/nIjwCvOQPrXGshzj8CnrGKXRUfpsuy9uINoOr8yZgAT9lwtmjr0PQs
rVy48RhBIM1/vb/c1IfkE0EMFUMn5AT+iGZLpvzRs/uXLWiSYzh5GsBE8Frx
byNqcPsZG5sK4xJZPSC3v8UjfIsqfNGh4jzJELfOz9PWYrcUzBeBuuQjlNpm
g9w+or/QK+Xx7//wVCls8Xf6MkZVKjWoSpyihWLVqGcDr/HACCJ1thwHepKl
bEMJ4nTPn7i0IMZpClIsYhBAe2wH+IWwmTtH7ubcJXL7ajvn+UUcpczGL+SW
OQ/L9xTf2k7x5QCL1MHaBrZHSIx/OL9hbkJ+spFhbFeNW6SIYeESZWN3aqZW
WA5wT2Of13Vr+SDmSWFqCHFymPHxJD/5yVQ24pcRP+3GCBHigGU22VirT96M
jJsYs8rTZuqgLhiIV9VieoCuLvJy10bqTfUEKKWFL4m8OblLisNJQ2Q9WQZh
gVCIOaaQ2C2nd94BbwRIZC6Mm2cvKX3qrB+Grc7euamR8dpT7B/kQ/uU8rDh
1cBB3DHa8G8U91so0mMHsH5J2Ov8o44DVQBTaTGx3Ihi4IMOpG3hcPGrU4xo
FIZzvMh97cpYPjRw+OwRLp6+mH7hOjcbrty99d3iSoKw3IRGeuPiZKyNFHD6
9gzgoEeILCz0mQjmi1Uxw6fNzVoE0FxMpDfNqYMePvzgvTdl7XSXrvGNsgaI
UN8NASFxOpm9ZFr3Q2fcCSiMm52ACNK1LXoIlrAISUBR/cr5Ua0t0JDG3bWy
4eK80q2tD+NTXi3BBZCYLXNaD+Gnpr/NNxw7gbszqCbEg0HNp2afQc20gPQU
14DqMR02/CWcwS9cKWv3b7FWkw5Uq2yMpcbiKSiSoPJCp7kkrIBUBFyNnlJo
4QwYJXCCn9ImZesyb30aiNgMBcA0W1q8mBKeCu/4C4uFCVv3j7NKod2EHMYe
65lmxa/B47kj2vIy6LdFsca3bBXjudlmsh0W0GLg5J8u7sdDkl6cgCbb+7eb
L9b9/iQ2VGDicJFPNnvL3GSA7SIVPwH78pGZVCHKEiH1dRk2BzeuG6Oppco/
VwNjnz//WFig6oU0Dfu9lN1FsX6RCdwEksfPxpwo+QZ+FBv48yVrlyS3d+Vm
/nstnMO0AQVTUYDvM6X2OAYBD2XGhdSpw6F0hCWZ5KqLorMqR5Pf7mzSNTpL
56DuNExvEalcYgaAm4wCl+rVwxWSHWEx5tAmHhJibWCEu2F1VbvBqqd3TDQP
6n7iRAwAtiUEouyEj6EnmrJDC8xPB1nN8YTFa7fLpkDsdUhRX6v/auXlt++5
ia1vN2Ss5hu6acCqjJgRzilglyeDZO2gJXRPAMUIUpLHvrdnht54x+hB2F+E
qgL8CfeLi3+HDLkTcmUam1fO+e1fZCcgOEmyP/qVT8zV3CplY1NrE4vugSrQ
xF67SoGnGkoVqSzQXvhGJhBYRdEZN2Ar7senwdaRZanXuVccUNcV/EtueYHY
oE5/X/qoX5mppWMKHEie7AZZFGqVTIhtIzCSUAQ+wXu6WxvkZW9nU+RYcQve
8l1PI9M6+tShUGrstp02bms7fPhwQPw7FOy9E9h/M0o+XnVnRbqSStMWUDyr
yXc3b5ReU544t58PsOYqQtsEZ4M/YcTO1voaBiFI6ZQDozB/FcU6hfbRYcMo
Hx/7MKZGDqD4rp6SkzUdjHhcTZR+NLwWJJQBTs1QVkKp1wmAEj9MBzF2iPrI
3wpARoS/UTlm1HLTyIa6Rlyavzv68JQHy11GiSsY4RYZRjrfh8VL/kAS5Shr
XTUWHdXUku2nPCVyIRtRY5ZmYyDc0w9bM3IfzSseS4q0STz8LltjLCzYx+vj
lfFpebhNGb0z1DT3kfPWkjtdI7Gwz7eJznUAovutQNTpnYahlQAco0Z46Y5b
cvrm3a6c+UE7Cf3SR3/A1wMeg7/ulnDxyZGo9OsyAeumY1cGv4Kt4m5yx3RJ
cpfOrTkKvdqMdp1sBPXBKbX3UAFIrpWcPt5eKm8FtUuPKvwnVmL3m7okcg+X
wSNlAowdMh79wAGoGnkXaJ+sGwFgJwGtPjl+CG8IWJB8YUOOIQeMC5SoJRIh
0PF+IqOPWpp2k2OR8G8TmoSvEQFV7dWB/bNRpOjrUC8VX5ZsHXzDnhcXORlf
83mqsjGtHlK1ZE4ouYK54o2uk51XTo9Ie5bOYdDRkzsF1SNy30nvrM6pIX5c
Qj0jGi2KzdU36zkA74Ir/EnFGqHXvDd/h8ky26/3UnOZ1Re/3odHAiAej3PT
gdgvCznIqiQ0c9JZJgmjWsiJhj6qxJwiegOCp+adNnXaXCizTLcMJQE3ytip
RhJLPi9a2S4HbANNERepSryoq9Q4HBIQREefMo8hxUugQwwwfbX3oAyG/Qs9
CB5w9BMIsRRVVrdPpazwkDhg6/cWrQ8C/zc8QDIKmqdHR4j03HoMg2MyuA/n
ximOkQ+WCKWITCzg900Je1eYYPYEoo475Wy8IHgjmIoTj05wejSyGa/WGO4V
ciK+pNrfryrmzTvPr9dw3fexEQoZ1xM9/PciAp/ikUcBJcwgrhYkW1OEVOsp
lZRz3Zf1LuWxF9nZEzV/YpMp6ImjGr7VRwG39kGFSLFrBCEJyWrmZ/JGgfmT
8ruAWPdNSgE3hmXjWUMOAIBuUezIdKW1ILmv5LibIzDD9ONd6yftkzSJ+1xU
D417ZbsiRYJX1RDwCeWemv/weF292Zmt2XuDOXCfICQSP23apc+ubiGSngYR
lrZrZqrLTRinQ9fbl6PvT8zd9atsKWJ1u9KgGsJSfDtJJL6fnrLklpbqwKVm
qsdhjBs2Zxc56hGPfBqWZBuanfaMZjP/gj39wiW9EQrrbn+xfPTQ7IbuiCzp
D8YtxKjc9jE1anUfI7jEcuWVTpQKUbw2Ho/bvDwiFmeOAPimUBNcxPd8qioi
BiF+T1s/NErbnV13Adj/TipZ+KSRzg/HoU9jQVqatU+HG4P2H04QZLhV7L0j
qIuJx42bjaFzqzN0Ke/NgrW4ObrpWBmszF8pAKB2HNpQVQVPqhQksR7nE41r
8qkpjY/0wyIiVc1nnkxSZJPntERr3IP+ZrjEL1//CFPdhNyuEntx0wgUcvHB
xNVtTMqQLG2si4cqJqPGgvhp5aOsgrS9vbha9PNYWewTT7aSgEe8N394Yd7M
r+sfdfFDfRWHCTdi7S+cbQ0kpQo7mY2htB/oUBG4XDCs/6YogopNJQLmpb3B
EtFNx2RTIzYgbgHMdt0JDl8yaCGbgSOy6boS7AZojLNefZUmTXLeXdsQl5rI
bx4MHl22/zp12h81q0xUrac9mIuUip2p6+BDES4eZjVVakfBI2mge4i6jI/k
haebTEDU+GhCdTsBsGK6nasD/zpYBH/dlvlc7Wd/7eG3apVgfJH0RfZOcHxa
AbhBpShtwSxa4S5hh1N95rPxSedFGgESy0kJ/8G7f05YhDP4T/R37WkKvKCg
csmQb0uJX5PSbAiJ+zzgB9PkD0qyrD7ve9mLe6ar9+4SyhCkGhX9OhTdwnEt
mJT64O2Q6wmZsqz2v9UH8KlIbglKziraTnf1LDn6anKz66RYXcof3wjoSK6L
C1oqfPWkhv+6sH5cU29Udly0KEUwb/9uKrC8Mbc0xtaE/9BL8fYu+BYX+Ltf
tTIXFlF3LjPA+0Ywzd+DqOPzkEmEZgnxLxpJoAN98ne8DgSo9/UZ9k2M77E3
ixLsrnKO6Z5twSEuOciJ2ecTDISAMYg5FGKo7cYnYf2g4nqeLkkcIJ6YVxEK
rHF4gTpMKeVIqrwgf5Q8azTBNoU8hwMLaZuRxnCOUKyv2yO7DKeNjiUR4XVA
JiC1jup/MbLvp7NQftsblzY9Zx8nU10jX9zPTaHq7g326RATcZ0i4yVidafL
nz2gEY/iAounHi2GJ4zx2qFeD5UncVxKEvCIiB0sdjUKp63WUnKCpo8YhSpf
xhhRW54l4E8VxSfBBHD32a+/OjDGk2noqSTifJHDo0ndbaoWYH6zErG5GjUI
C/uhnfbz88TUmktagcHnuXCLrJ+vEwRskBKqK23ZiI7d2ujf4HB1BTy8T+QK
mQxRFsdGL+EjdPnezhhRretUHNF1ZbW1Il1kQ3Q5neDgfAW0X/PdTTICM0db
T+L0N7OkXQMkK288JbIE8X7KhEDzlRv0kTDWjTqthlCusrAI+l4SFHD3SoX0
OAbx05+RmDBg5eOogcvffw4mSQvT8MGel+28LXAL3W+w8YArq4t3BdlyFck2
GKJ7WpnKVoQ/+b8UJHNs3H+V/LmNez/X/KnRB35Wnh/JYFnCfuensK4cEmpV
ouVJ9h8m1dlacQ3lqjfSb+QmEmDS6tWoJB1yOgFWe7Th+kY1ns/gPOjj+1Fd
5ULqe7u4KclrKMOBvlQNWfoHVBg7bvLIkuRyQE+eqwjLjUnINPyFOFaclmWY
V3FcSrIHqiIY9euar9ICHC2kIFcCTvwy100p1xbKPXKq5zLTqSdfYnYcw5Ta
S3XjffzJQHZzOMgJPtBEMpBHtB3dDoRgg6M8bUY80RtNieKdmwI1NS8jlZaS
EkrY+BASW6ITm8wgX/W/iQzs2LWJ/Xo7oNxQCgoKXD6wGFwPNPB0Sf/R5y+S
Ics+ao3B3WR2E6FRq3+plFhaaTVtPSB+u38tIH1vvJbTOBz1LFuNvq0c0nTu
1Mc0WU+bsN7kvGh1VDfP9FHu9m/wDxYVrLNYdnlyRa35uX7ylwUUrBffWK02
kdfC+rByYLvbunasroUlF9ML+GYiL56YejXNTPZOrmFPOlwESr77slAKztzH
jdDBmEU/aJz8uN/dioe45rGCcup4aw0XWA6p1kanY59FutPgHyutkNVi+YB0
M2VvqSpDb2ddVrdKH3CzwXuQI2ctqpKPb9XfyaOkpIg/MqCuWjtxlkOz8wAN
MGGa1W4mG3kX5HKWXd27qauS0gszmY+prlYzA6KNqiyoCFVjytkIRiOVw172
/KHBgxngAlz/iNM/fYwUD6E2oVo29ihtSanVf6+pVYCVLKolhwP01CjT7DdP
VPMl332IeAMIO4BaDk1lhOWm/q6OuJKg77jM1j09YFyQCcQMnlzzR+0utXQ+
U3sAadWJxglODopfZzXdNxcUXa2Y8I7uR+kXfXcGOFFWdtKiaCVLeCD+JDzk
rlIHjgRlLOsxWgqFsW03At7wTIlFCwZ9DVlRzP4EMzCedhq+PH+GA7xZAcW9
rGIuC8/rTjwYvtKBBTSyW0AS2DNVPgAD4D+XMmdKKQMyumt2Y8v2wf9qJn2H
njPOAKBGABCqaWKjW8ZoY9sfvCDiBuADnJFTzAZBldt1VkDHFDCXg344v8ub
hAV43tt4hzonrvesNV+HTfQgU9+S7P8moUN6A1RinMQe3b+naKW/+drLrsKf
eF6Da8w6zLkUsLwpubcijUC+kJvfxVGXDfrjF6X6qpoGv0tLSAtqAictQMPW
ayj0MIkY1aVKwvETU9d0ii9SfdiIOXVCwHluwzg931wrb7sHmXxKny5FvKg7
gEVIkOCvr3kvEeCaRoq+ebh14XzHOH8tn7jbjW4MOaz9vbO6mq4zUnxzNLWz
PUNgRqal0QDC5SPERjf/WnTFEsYdLF2WO7Fw0Oplnfpz/EOwH2wbT2tqBq68
/1sL/QC6yuk0Dbr8zro6un253AKRL0ICv8SJQ+lCgcpvNepg4QUdYzgDUosc
BUcMRax3gCUe6cWmvPVlTH8xmC1shbQMR7Tjt5Fw+iHtsI6HOSbqTnNqzES8
/W+Vo57U2eTClY8AztQ2ue0ia4UOpP7mVm6Nl6R7iUR43OkyWHBMUlqpJXle
OewPP2NOS3yOSuz9yHrPAHMLnAa6qv05nz1rq/zJfdDtXun4ot+P+fF2a4eg
14gkGnf4WHvwMXl24BmVVVgajBNd32SjTLm5bOpbLGHfvTYCaQoYc1HX/iTy
lJSB3TNivH5yIu7PX3apR1Fd6uX8sRTUDpxvZCbFcNllhLjDn5R1/xV52S7X
Mdkt7Xq15CeU0I/9gWVCGBTFCl+bldcO1u0fqn3t2fXG1LFtLBVjIQpmU6fy
aRt4lVRVzBpt7vVKvo0hiZSnyG38IoT6O3B3tA2Qe2y2YQvB9J/FlSbeHpr6
fkJIIRM318JNfil5ITc9Em1WHqgpVmei3F2T4frl3N0KFpMS6h81v7JdCH8g
/6OcxxhnLcX2we8Nytispi9O/3WIpNtA1ffHy8gK+h21nrOVw3OggyJbnUaW
nwz5XYfu/WDG2eleIYPlJWuPfrvG3/7jNnbxGfsceBTbNdAR+tim8AMaDKOB
0F/tNI0jTi0Lns/IhX135iWbK4k3AGNee3pKKXR0yczd0wg8/EnlrtnLJwKx
IXxbLoSzeUJstCWM+Jibks0r98YPQFIQmzOAkXAeVgTpnohU/VBoUDlkZRjv
1n6ycyoAMuQL3+ec47PtHmBnVkPh8s+IK/h9JOsOQom2HEYcgT4hbmMpXRqK
vDEaeEsESqiANc36VB+qs4fJjuDYyGzBVPbhPpJI0I6Pj8psKVKeQq1dD/+1
u27kiQ/HXzf4lQHHoNaxnmDFAMiEg6u0R7caSrLcjFXzRBeGtNoWeouwBnDr
qRt+bmV1KTDwOLCmRW2gAkP37REuGmrTtchDujrdlI5TcyxORPj5RO6saF8B
pWT/665+6qkRQ51nZ3Kbm3GuHpYLD3pB+fvewZwrKY5X9Zi5FOZtQLsRd1Ko
+mbVipshzQioK240hv72t6Hq7j6ft8BkmFw9v1LHM6xxO153jr7OwliTksxu
po7CWBs1tXIzxI9Snf/zhRFE+CmAPk+/aLdQ11thoEmmKb92ueTrPaIA8M9g
s9dmOlX/NQcINddHNgHIxdtZL4lYxqP8Pq2uXCerA9HCQok/zG2eSoFOAoXt
4AULGcsukMKMQV9H2tzyfh01mCXq8rPjIz7XcnQFIxVvEeom5RD++k+zWn1p
1nzWio9Z25SJEGYV4tdz1RDm2hd7JlECpMmwQr/6KBuKZS60Ej+qPh+KuFWJ
LWFOS4eZz3ZQK7k0Oq8mNbVoVBeJjVXqtPQZUA79QjweKZNhsnHR4HFC7nEn
wWqRdXsh6FsUa++Hw7sBaFhME3htlhebYDoSegEjVf0Gkr/bs8l7OtiO8omQ
GRep7+C6CMNghCYK5aVI8WT1DAjSp29/V4mzimqvZ98mxHxYDrZbJ740CyLd
gWnT7XBYjuXPaQ8tDeVkagnE3NnO5bJTuDEr1tCkKP4PNFkDGcsP7vRX/Ojb
nxrCW8DkX5phlwCz+FlaAuxyjLS4khv1rCRxw1TgxH3t5gwO5iKNu+DjhC4m
TRIGOY9aaEyv1YLIV+wjjOrDZbFxA3v9rsh0NcyYK8KscKOKRD0pnzD9fJcY
DCV8IAvu/QIsxVJjHNpZ78Iw6hJalcB+Jj3oGa1sEr0WuAY3U7mkE3Y2RBHd
42YvH8FezFWV9RdczBQrIXbZfXmy9j/9B3iP2kV6jpkrMReMtX0RpXB2vNw8
SCoe/SjPW6c0SN3WPaG6I7B0haRjjkHz/dVaCSsgFP7gXxh2CVhl0vXKRqJf
fZxD17vTMdBGqcRIoF2x4r7RVMGbONDmVGrfdvCGscdJJ+BY9jhTXt06l21a
ShoLxlS0n7JEf2jJRlmBLMkeMEyJYuwuSmbIK61SpfQ2Jhp0fKFM6vl8qFbF
Tl82UtVe7LzDIVkcuYmVq/xUuwN9HhKWWnnzPr3rLplXNY02ey6nb29b3bmo
A4FEhsasEgpSkQ0phAiJXRW+dNJFx4zVt/qPaZIWPztTvFYinwbKheYfoO53
Z9MnI/avXtHbk8zi3lVBxbW+tmjFJ4nXflmb+5bi2k9m9E9tGdN0ylicZ/ms
PfqJi8Cmll1sL2Kp89G1xR665C8HGra2UxmD7XDWHrVY3ezuxtV56HSL9AUq
6ksofy7gjI1IscQhx6WEoZZk/a3Y9k5ctnXe5asg041GkaMUGiTSEDkawCiK
Zc3l4E24ZgB+lIhnApENUlFdDreS7uYYsCclYkDra/el0OYRHVsjMLPrZWco
v1FiK26ZlIOfUfgVYg0CjuE6bhy754EN23g8Gv4Sg9downQG2YZxSwyxOi2a
U2PCguGKyBRTjDGGDC+80QVSAjpHOVfI6GhRmqx/oVvngONzAGhYkso1FrQ7
r3EoGS+J6iG77ejlCizNe7jJxavMcKbTeOGItiwb0pxZuLlhEuRfeRrZ0DAW
9+1utxd3sPQZpAcYXaTxLyjUbC7yYBcQNuzXmUTMu1zPB9eqez6fdcx/K4te
0CDtUL041eC4VUGcV98yYq+pRXJwlVued7Vf0E3+QO4RoK9ENz+pE3RK5LCH
V1WpldiPs2V4u7LF3+XSanqXxN/kmX7SDmoHGEBdMGdPS+znbMc08ppapb8z
HiRGPt48qSXPDTwkD5lZ++zxSDANj5rHgSruHBLwm62YXY4cTEpJmEnLjRwX
p+sph0K2Uu9bnpb6bcxQIk01JpQJ1lmUDwdvpVd6CJwZ61fvy7XruGfc7HsJ
usJ0OzbSb1U+xmY9tdQDK+fBH57/aFZQpMJukemyIWi0V2r3pa6+UXdStFQP
ndbYeG6XjbFvJ7XpdzkfV7ro8BksgUiPaionXvaaZCLLFRyqhlri1IQfqCIe
dHd+9ntqJQNKshOu8TQOrvlc2jqIMyU0/Ue+FzOdjyqjJHLtwVhu4hdFz0c/
lY5kylCxDBvJvg9+/AQMINRCzpO2YN1orYZqSzqlP60QMMEYCZyrGzx7hpJB
4oqCnVMg4kwaFLlWOuX4Y/yG38dHelAChtLLMLp4MtzNgC/arpZF1Qh/cwqC
ubFsnFq/wghk+Lfqa9VhNTHfQUZ/u4mWFSQf9JtTWdX4JHOe+bc0b6II9Ekb
HiDl6IR1Q599GI9PUG201ppxOMVVUHRkYUGhFzkQms8AuScUY0GuVm6zn574
CsrrVlQwBMPLM9DO/YZDWDVyAb7fx1hmVtgSTSTEloMhVr+uvBN+QMNI1KOY
EoOuy6vU1ZlJqC7n5FP7B6iAyMmEtn0dmQXwyvPUMyGZYGB2UnxD3ZYEJh3+
6u9bB6HjKDtR8RbnKI4aAV+BXAWp9aXnBE298vOcMMvwNBYH3nIFDKllkLMD
MwOI7ybRe7dbZ/ESaXg/fhX6QVF54gcn5aEJKagup9GgI44IY7b1ZeYl/iO4
haD9y2rS+WsruxNreCimT6CnxDgVt5lD4WmzvOKjtAP8cihXQxrRjJFScssv
tEyWrv57bRKdYmVFVIMRCEOycdlnvotcvrgHvF5qp1jjlLuWfb0G/sfHXH6C
0znWrqKS0l0HDnybFo8ZOjNfbUZ0qXrN3g5e6N25UlgXjb8eFAqm1KwqrcH9
aJshjWYDDvtq5PwxePZTTfQ7QQODlLt32tohMcX1+gnWGsC8OzmhSEEmOfY4
nO5Ff3PqOo0wsyBkEHQG/OLru3c0R/2O2/XnhHxjhXhA4TD9WXnQatpSR01g
rfXxOzZ9cIs44QmjmD5cuKselV655Rrv9xkW7//jMQo9aQAlizD+PLH7A0fW
2osLhrpPUVqKfNxN5czeemk7ZIpPSlhBJ/8DtrPv2S01iyGI+ghk9GEDHlls
4cP8i0i79lWzvLtuet4OFTdsIoEz++EORgEIVlRLr1AuKxHwvEIHuR7nsjIJ
4AqxuM52hnRLi5pC7NZhx/8jOYRHjIaEURxANRPiAGPfCf3oiFQ2m8UI9zCV
4KfTLVAwvtHFiC4nXmB1WSfCUZ1CSKD1pDjEPrEnVEvfdnDOBIvEaOa+gIm1
WgPPxQZKqQmJuqX4oklZ9wy4LClILIFKzv8a7fGmgvxpKjQSlj/HI2hwpPEE
2wy/Mqq/TkHxVIJUALwaXoPujNhZxn+GhOMBEQsMVISDz8CGtQjgD3SK+4Ew
/fPVlZpQYvC1PcpkaqIp1mjSveIFW5RyQOnPhqOHokk122is/0GYkmReeyPS
6IHPF6311WehKj2Mh0NYfXaH26elY2UEjDzrLpZpeRzF/+0G5pnQcyC8KQi7
h1GXVkrhE6LpYs9Ojf0xkmvvqzjFYLHlnP/4r0zWrZJpJtUP7AJp3EDla+7E
FqcTNKgOne+XBdg1TbyZHTB7h80UBObGCuAac/78KWr3cufLCvTtSlYXQvWb
NhyOGkevx2NIpERyCU7IowwNzoWiinUMN6miiFkHS6HtK45t3dawRSheL7n/
caz4kU3Se+mkIC/qWfMPSLmMQ+D+JiawwGFZvGGuuixLJQRur9oOIyMTminM
SXx0y0PJ05LYaUARx/SdVb88SYpO+pTgGXW8W68YBQ01stmW3x5AEuGYLJdc
N5yyzdh+D2p7OKQxfJT6ToJi3GKeZ0JFwc2W1ynbHW14StsE8p9ThT5PB2zP
gDH5rhh6xAYy8gqh1Oh7vCOFjRcrjepcF6L88LELdKOGxtm0wudiooBkIMQn
7UItW66Rov4cPCI3CNHbKbSmzglzc/VUaki9WJRxIe5vsyT40hZ2oVcER6ds
DGRN6ELUQsO7JkvP/ZVt4tmsfNgGJBgn3ft6WrkCJKIoIcmuTpdSW49qQaiW
+kst471pAeUujUa3eAJQTBAcEA69DtsVZ9gAGy4Or1L+T502vp0s/fo/efBd
q3xFkCznozvdRPMoFcmUbbXsBtVJTOj3KQymwss7HLyRGW9frXnA+lhKyt4Q
1fx4hyPvWxT09T0M1i4ClPCIe0pt19DBk2jSMn0kw97omNGS5usA8PBc/4Ak
QI9TEI4NxgpnKuqVnhUc82D9mE9xs5wiGrcV1InutsfrSkb8ycADmkBZsHQj
1+2tL8Zril52j+OFVGqHt7rxN9FChXXXFPhd5dSY6u+Nco09vvLksXZfmPzI
1ToebsWwkpkUyjLXTtDjG9WgONExZlcW1A6/BWssd9/v5Q2jERQuxSRDYnQZ
rPOYaPLfkDJ53//CvY6QavkLeqYRZPq//P1QUSvGCXSgJr2+hbhtCM9NyvvX
uPpwZg+KCmFl4loSw30G7jnJleLIuKkPg7CIye1aOhZWcaLZfWJ5AelKXOw+
UGP3yrkVexxlqT0pqy5agiapkmk37XsQZWNdtT5aFoMQ6iBwFDOQzrlQcfQa
lQ7kSyQ0th/4ncrOsVmH7K/wfZXV0jyquuY1K5qRvh8bMbF/MYQcDQCUo3Sw
kl1bHYu1MBU1PC+qGUAVrhC6zw5Ma7HJJltP+CPhBu7gHVaMCNWJIK+BZfRH
5IkTaOK1GyjYEQXbo0JYkqdvFiTXPo4xu086drkWhkPqBjMt3ZxIbu0tZlBC
gau2+TekwknO6bNbZXgzQbfW0LcWe53MPzAgp8Nk+n76qrY9i81OzGO7bClz
35Keq3xCeXYOJmFBTtCs//3pdN1nnfFdsdRoFcajY/ys3I7/cAC9gxM4HVtg
IKmQpKNcXETOtnpuHfFpS2IqmTEcvRv/PAL0tDE/bZFZnNBMFkP4gdUPwsM6
SBTTgABR+K9FlgLE4Kx4cdo8Y5SZ0QHz8qe+pNx7PPlXs7J+edIDpdVe0cMH
FPmpn2lfscavAViwILU/AYtWNhR+FLXQli4ohYL0g0plc91aJ0A5VdXmeTVe
seR/CeKND0bXijBP8SlSuTx3bNYRuemvZ8/Lg2JVr6wLSwdpFKMuLe4HXALW
dWlQBkRFvY2bL6dkkGwG5Y0wCMbn543ICTTLsU8JV2xXwB+Pj6UQjV+UqwA9
QDYOlywLUnD4KBip8FCLRnue2+g4jrKrHMdOa/TKZbE5U/a0FGF4GZDS8mNJ
f5d6e5lhnoA3Jhp3sj+LQvaSyl4FeR6GLKQwmz5Ztf8U/EMnWoH9mR1MZSfd
or1Rk1p9bsXigMEibMwOQkgP4pU2voFt8/sfdv0aLJEtP0uEZinyeC9dD5fF
prxctZdD462qDGRG6mqmwUsIJDJC/j4fMF0QMGAi4ZgFxFXZh6cQZ0pBYaza
LMpTskgWn9gA6K7REVtD3wwR8wjU37AH0u4sLbQTbDvLwvUBKJ03SZLRl83e
1mdySTbES1Ydsa2/GyVbC+JOTWe+eCGp7YXRa8rPa02eAqjye4FQa6n+5FZb
agpHrzlVZQLHnHlQyOpymhoZjEGprGTrUPb8tZYYnTnL3WCLseGn9hsTOLQm
k6dstwX/bvdhgGk/pMkgIVGcXNnAqkDKbiihf8sqOlm4Ol4dvc8FfmV3mppb
aExvDOnv6hZ+iSM2zbcranEhWAyKxVzjEe5tsJ41TgOoOfqZahEvZ2aDw3ON
IO52/tieBLLO38eaHizJYj8FW4njgJrqytPlesVwTIp53IoPrl6ZgthEkaZe
sKAlZQBxkg7Xx4aZ9i3DlesGmxXiINhuH437P7CIOwx9qfVbl1Ud2X9xkwaS
qdubiyc5UQ9P/wzPJ1ukOHkPd4HFywZpZ8xtFVWHYNFbF56IJhthRHClVPom
bme+vcA4cAcmPD2w3KWHztIkKzEBfwa2PT2aLMurhhH5EIRlH3hpnkjfzqkt
Jaet4Ws0P7sl1IWUkWvYHuP+e1JodGkM88UkD9mNXUSfFbpax0/um/V15Y2F
cQq41TubHIKMXlrSJf8mXxQS5y9M/VYhIrp+oxG3o2vjK/SGwmsfX9Q0EL2+
IjFWf3tEOxuA/YN8qBvVfUrl1Sw9ckCBJZlHYmdFKxHA/iiumRGwZtTNyTuQ
ogce71ae0m6l4IGGk88DA3FT39rfPyBi76Y8YwYSBBlZBC0VsiIKxqnuIWtJ
BYZVhGPfNkv2QmlNIM554AU6cBOVCVaB2aJkMCqfZa3OgA1waiyhscVyca4N
P2ZgUqtaKVSPOOyEufLly5TczGCCvbfOuOYRuLButIdITaT/aEzPWXgwNY6a
nGwF9E2eTKp0Xb9h41wYxodWnFcIVbw31it2HFAYs5Zul3LGQ8x7Gf+3ekmD
g9dzNZgoGIPE6M2wC0bXPdlRdiETi7fqwx4+ygWYnbmHJD8FFksivaOYx3E2
zxqYO+jQxx3Ozm2CaR9eqYW/TVZd7ua4YZd2YvviWFufpGHjD9V46mSXvtz8
x+sywZPtNEcfhWjBl+3PquRxYt5oKctMz92taqHzkXc9a87RX735YqR1IA7M
3EqRin6QBBUqKSs2LSrdCMNFt2fR/m686lDUBfSpXAlTHIXwyZ0r6ho1Cb5P
5cvTMoZGaDv7kf0g5iQ/5wms8KU56ofzKN9YOLObRVuM531lfrwwaYGe6nwm
OefxojQ4BwJBeO8cndp2wEQZ1+EXap4O6K0acefs3gj53LiMavxio6BMralL
Dn9N3gr60CGoUdVwJEEWjZaFLQLFMJQmnimeryKRJqurU1zEh/ZhRASlRRxo
dMWxlMAOxBVh4+LocjIOWDANw+iFiTxa6raiZYnhoGdLdzb0q63r1rxjuDHg
zwoB1Keed72IJAflibjsqCE0CHijpYCWyu5PQipu8D1URUALFoCvvWz5md9t
NfxyCh9N2bJPIZZJ8W1fUucVfui/byfq+9nIdaV6CFe6m3bLkDiP8+WzyXUD
rdiKIIyxbnBni7kaIXFshUSB348cXK89U2HAszn95X+VrMGISNmtu/F1usyZ
7FmJT8/qDPFt3OCJYA3zaQK/flDpC9O0cXftZLOtn96iAFPB3c1EAyRtfw9d
7bu+INuJPOMV2ZIqSADND4r/NdgrxG/kasKA61QyNdExJ5tmvDwcrFgZ76Lh
vaHazwweR6tiEvS2DaEgO61n/t90dUY5lKLVDTmXfHvYiXmjMcY5bzywsTle
Hdba6iqBDYzw+oasZGt0+Y8vfIRL+TW41Yo0r76T3pORClb2d8t/tc1FkKBn
jLMrDb9U6hH4bmfzMPLdXpsW/q16bbUsKfFrpZfRv0ErjGBMvCVswZKd6tsq
wKR4wg/8/corzSnTdZ2D7dsXt/zqUcsNU6u0obg/DEbo6KF1yssQT+JJVM+w
xcPfCv/7hKo6olZpoEHbvcdPC9a89t3bN4iNknBksjCyzzyg13eXAgfgd0Uo
mALuHCjCJqjRMsIZ+5hL7JvnbQUGOyWODmk5k3mulzZMZCdAOXSC5PfAF56t
ggPZeiBnHc/bBeoXCduYxmn0wvzepaZcc6WoISvjmuLz6SRU3xXEL3AVE56S
/q079Q+d3mAlsiONB6SuSpBVeocqZTlznNk2UvzDETASvoeEgmpppFWgpprx
whEIdXmOCGfeeRlXoqHCV8ABylMaW7L7Am+CF08p5M+QjM6sxb9bkyBmJ5Dn
HM2A0vAWRavACZWhb76xK1Ljd7H1oOeJz1SwGJuPMyGFO6I9mzDVRczRSYhL
JWn9Opp3CmDtXWmGLHMGy9Vkz+9XFXk7SXF4zPdQXKsPP5fkhjvip5vvqODy
A9A5Sw1fLqzveWcQhzBkEDXomj0XJYFMka1MJO40CYJO/hjvuNqB1KXES8OR
EZBn6aFlRBsuZeW77tUdP24WlTeCoC10AE1SK7bdEQkhumdE6CTghhm6+DcX
VfIbdNf6PYp6KOEn4cHciQo9rs2YTZYF5NZwdVPQM9SY2UsB/C35nnKd4+OC
tNOenPrmKNv7/ehPGfI4jKoTA/d25U1ievnjxjBQwRFdohPpKPDWl+8nrIlr
zC4uRqMs18v8dnV1rs2hv572XZIynJej0NGSYS/4kjiM2x0gvw5JAzPjm+Mb
R+PKLaVlYAUugcxNanZi9i79qM3D6qox7sM4TfLT301ym2qZ01RNLQlaikoX
Be6jO9sCLw/aAd4EHI6bylgD6QOC6FbwQF70Mhwse5km+N6bwGZIFiWf5Xik
3L0ut9Zr7OxFXeOC5fK9UoIUfbOL7PPhc1FKf+iNk9YeLdBQ1guf3IUgIFgX
cxTWmR4MgOJh

`pragma protect end_protected
