`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
MuBxe7k5jQUiQLBqvTRyvVnUZScg6VdSanouDOSQGhebth26GslbKddfyCqqblW6
ie7OFIzM3XGhNx8MJh7QE9Y1dkEzkX4URFlsxI1Nn2eOXKL4lmTi765DBWFHh+ie
LjBT44zU5zwpZ5jxMpynw4vKHuLNDOt3iVIfOrksSLw=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 8848), data_block
YWtK+XhzLuo5CALZ6C6t4/vtUDTYYRn2ocDE7sNA4M4TTJvZ4n4lShhtdIPzZXti
kHwKZpGIlTBmNqglpDNdF4UVa8Ni62MIwYkJwFO3gV3N6fM4EKboVvF0DhgWI7qU
yAzCOLEl3Mb3gTR1ReW7W7g64O8YOeFOYoUMDIO8rMDAuoAIAZdKmDRdhBGcYdT3
B1E7g8oqw3j+BrdHpg6crdyddzL9R6iYHMoUsLQCFXinug2RBaKJDO3XVl1OWrd0
rib1jtup7Jv8hSyWcHfoU/5wsc3OuXTuGwTcGPwnXf02YyPiOWP7XV6J8R94Ok9c
NTCon4Wo0NQkvsuivN4ZLH0tq4wNZuqo7Bti3psvXrqzjMYf0+e4i1obJGZi2hYC
Zu+1pG7foE9tHkRn97F2RanVU/QiUmNnmCLq9RXN4mCRcdmsGt1/A6HwHQI9dNjV
tU11zhVogd+JjqDHWRPQ27OaUpLMiGZeSNACuRxb/k5L1npkpwD5syoJUaLlsNUH
A00NnQ/OXtgkMmDlRrepNiliLu9ii8xQHrstmdEi8xQ0lGKNB2arjblj5p+fzZXN
rPn7B7oVKqmWpYrKhkKlPm2rLHqgZaMNmGxvxX7JL6xDef8oKsiZytjXIPAMVSSA
2lV39LNc3Bel4ZMZwmjtWDaRW9ttdK/b0Z8t+dJ+w0umMI6RGmRq9d8lXEZ3FnQo
ZJFU4yjAg16NHi1fwguU4VFBlMD/yA7RNinsJfKJF3BbB9HTlev2NAwXPxmOugRr
og7SydztS2xoGfkV3gP7PT6dlLsU4zCSH9XL4Rus4f+h9QavTJW1rZZ8ZmYNSDNW
CjSykLAkpso6l9LzvEAy6cud/kuyiR6tdkcOwWlceK/XXz06k++3Rul3gZyCvrv+
aEirV30sjZxQYo2vH0Ui+OGctmP+iXMPELC3ineugv7onC+lwqImBy+TVWeOsyB4
M28CSMcj2l7t/UoTb9gwJ1eJMvENnKkXEKwnBuw/5FK/RAeKqaXxzNGK+MREj2wG
ADr94ZMhhXZhlsDjlyqlC/cXSfTTy+aQcuz4gsDNVdZtOyR+9uYz1r5Iw9EwOdN8
GpBYn92twUjKJOr3hFWaCZniA4WP7Fjv+T3mkt6dcs9FA4BygnMD6mYoXQLFOXDh
dV4YZ8bN1mXgaumsGbn0bdE4t2UEUMlYEK5sI6t48TYjuXVAmui8p5FIQgy+aL0a
0xmUUtykHPmMIogeCDN21mSPyIVVF0azormhMQzaGFonxBX9NrmnQDfmTgOVrZbl
I2eG36PCA+7YaWFbnjWabXdz49xt6G/xZHF2SrfzF5c0WyhfvYcw3po7I5h20xbi
dKDOTXV+pqIFW7LkGWOX2cFYeLv5ZjuCjPIbS6KEiAhDdvt8+YYyWMIa/eyPnuAG
hih+xHbzYBWP5BVK+CIs/lLDybi6NA2SP9aWF9hBa2Cl2Fy8Us6n6grrpJ6k7cZh
qK2bdLKWSVKjXCtYARF2yiZ+6m4dZJIwBPh7vkA1q9N9wMlykJlXIIpZSajjzjyI
PMMzBpKro9wHZ8qTS4Wvqeg5n5ginJ4UsJzGV1YQM0YG6r2jUz9KAh/3XeBAHOsP
Y2bXWVduaiA7KWvZHgRQhGBpPI7WjLxICkuuWfaYMVEmXAlZyFAS7uhg7kBlt+I4
+SSQ2BcmqdJ0fMyJLpRXrIdJPRzp6Mk3mQpvn05oLSvjIULhNiXvMhJKL4hIB1yF
mk+YV4yPjORRRSPgjCw2PcIagyH2HJm+l315zORQFZsfDmhegh6o2YA5feEkrtzE
73xEkORg2EvJacOlDKv2D9CO9mCq5Qmnvdhy7eQtA6oUstS8iwndOAKztZpfFjtN
oD9HuCHiFZboJwa49cGppSZcKf1z3+HNf3sxuJwxPDAylvjAYizcnzq5/RxOhqI4
t03FvHa0Cxmo8bEGW7bxAAfYkoTfmLZIEKShdrm7LGoTsagd7efXc6i9kz/egALB
//0uCsdO2XB/+4DLY1BSdJD6a//7q+yO+T6zdxH1TzdffFs92QC1XuDEQd5W3942
oXiNVzheLYkKuMHQTSsIpXMDICEGAgwCSgQMhrECWvFBSpEinZnHfmu1eGUyJueJ
MtUs06JYTwQEvD7AaDO7y/WTbanzZiUmgrZw4ugmL9Ew8HUxD2lZ/KgD5DjKPOQV
sCZJl7HlMmzUela1bWy0biI6ij3/VWDG2T1ER0zlgeQ1wFJj7tR/AQYD9bHUhilh
SWKGfH/c0c4w+VPLQxfdoRbqwWIxS2KjuBERIl4Tb8Y0BCNOZHZ8ereHSqZdA/QL
pyxokyyBp8VH78CMXYInBuKN0Iid3i+igERQXvLTAYjlIMlfZolJ/uhV4G79iq2/
rmdn/FAEeajFnY11Uyg3LYmRAeMoPk4RVMqKETJVtJNWhCXjLO2g6JLgtnKjEjwk
ND8eQ4teEbNEa/qe3tXisROdSWvNKgo4x/4Y0N6Y8yxNevwVoFg5lgfkC8uWSjIV
Eu5M/cv3ajJ1/FW8Yt5jiOIz3RoNOY94poKrL10iTwaKpqs4Ly4z4oXh9gxfgC4G
t7voCjndLebiihzTUkVbgbhBrVPBjlkLxSoIhR0tuRviNuTnfVuLMXHfSkaiQjQb
jKgjkU46I6XPhAqsM0TRe6AZq/EtNFLjbWTfLXuQC0XyzBgOiNHO/xdY4Q/hwapm
yMJsB+TiIx3+JjnnCuR/0L3CgjmSOg0mrxDg/9Tlj7T/i/4Z/uUKuNrf7Gcq1GL3
w5VEtH87oT0EED0myZTy3K31d0tqwdWONhzssnvwvv2Pyes0pdxrivoXwpbMTwmD
PJyFJm0P3N4yhITfe2FWieC9gvZqQWp/69hZ1V0C5rjwLoadrcJ5kVdjYiuBxzMi
TMNMvcF2vlE1K/lU3867CG7ZWvJiXktmWF0h7/FoeI2pyyGmk6XfL7R8aEHCP5vF
ZH1sQ7UaENegFEiefig5BZKVqZz6iiuQjF15TXqerbmFVPZX32TfomP1EFCGTVRe
CdbOEyA2ITlKs9ymqHfowauhdM01RcWiQocsSYz4xagOUpw/bDx+pGjkiMDnad/H
fd7XdhplmuSsvXP3WvALUD9FtggoAz6GbPfChaK1YG2QqIkVn5RM8Z9C9RUAQsrj
T3KVMQCRzk5tx/SXLNsyt0cJjjEDVb9H9dlTlnNG0V28NknbY6WihUScdv5LrXIu
Vei8jzPyGkpHSdAFIjXV2XXDdxC0vdTnVfStYQBP71MCpldn/bL22jJWAXPK2kjF
G5Bi+uM/RhIUD4FomUpp8kSJriOGwVuLNL4EOoMFx9tf1KYriG0nPMVag3IADaej
2SjN5YlXlwlrZdJs1jm7cj7VCGQn25OTYZCKNrcLjbeIzas4vxMFtVDS+0XJFXkc
IDGTsNccob99ogUbkfJfoqDXxSxcGWrydviA4elRYU0CYZDgI8GReyxtpP1N4tyI
KDDvZ2GFAtaWvR49nQMAfyh/mmgBVQktYouEO8yanVPzBs31geFQ+rHJv+BoRGU5
clSPI69I4TvgYRk/5I5L0WP5YTeh/IZF42FCdBbi8USOyj9Ohtv9W1FtqWEdJu0U
4N8f6O2mbvWwnrTzm46NTG3XiLbUCAfQwMVeEgoPlU/UZR23ePAATnupyhb2Euj4
XDX+YGwUu/BT8UWKiuYjVHeKCf/LJrLDZPzMpRyXrETckcs27ZKpkv1VVy8HXDT1
UjqoeUVmUOjX4cAet39jEb6tencP3xAJU6wLVp0dVpqlG5FRsCSQjJdFeMU66pVr
W8fr3RdsrsKAF/MAVFSUVDaeTsOPYXUgJhdeKQ6y2L1bipXNKH8eC0Fwszn7PkmH
CqasSjSbKkGGQtfkKzbLpwQKtGX5oFcvUQsiTwWGDdeLKCjuYOIOnbWNtZyCXzZk
6FpJFoyZr6PdEVHGA0GZpaHlsiRtKTvyte74Dhj4l6goMxEMDF6mA811PpNJ5bYb
uyk5C79zG9Q8nAMu0aT48l6PBZSzOPIZmbij5i+N30+rxf9heCg51Kc1AZi5gECQ
tuvvQTwhFymTSPcAgQpwE4izFTUi2iUOZGB2Ll70oHG3kyxFs7/KsSk6MlGE8NLm
KlcYfXF9CPJvxdwf3SQSI9VZNLagmPtTXBNFhTUctCpkMYPixcelVWRpCMU2TCeu
XeOWVNmcQGGZPJ18y6hENja9piY6O5wxOXzFeyG3hIa+jZPvRzyM3vlp0eT+gbg3
fWAK9BOIJIqMgn/ziegLCyEwrrwYHTHVHS/EVGfFHLzfiZRY7SzFgaN+zyMvo5S5
T0XyK23fmlUeAj5YFS8Bl5TiZ0GwY6FH7ZcVjyAi9nWYDzXsE7AJHI5GZgk2Hd9n
Hfwd82zttPWvos7lzbPiffaUAk6OhRHut2N3kgnC2HOUkJMRb5t85CBslbeM/KmV
TzaG3017ik+sDoP/lm1D+de3E0e+Bv9lb7DicBbvzssrKzhh7CzUSXQ0jDvp0G+n
PppXHwhWZEtNknbNrHT/PQeDT7DstUQ8oCg+bwcIXdJ/XsAHQFcZc3ftDxOij1LJ
Umgriv+lY5ue2ZRdjK2sIEsuGQNQuoOmPXzB7L5Aaqwrt1C0HoI8pVJQBXGhpCnm
qFu84eube/bLVjxyLA+o/zXtIS4B6kdOG0b6Gyg8gtnLuXqqykKuEHLeRtjsmbry
0i9ZGuBSHR6ASbOfL7bX1YWRWkkBUqPLi4yAQB+G7SEBCtxugs3Id+ClUV+ROwek
8cd74cVwIR1EGj0Uz2CUgOM6rQ2V4/zPzjc1Ubr+qQgN7Q/HS3jl0t9+4a/RI9Ye
R/10HU/mmdcexWZZIidLuZ2a1NjcFc/72Kyeg9MUJ5Ry4eYaFWgH2G6BkIWkAEGc
ojrP1nmarjRXAPirKc9WScG+SPnqsOEXg9zx8tYym1Ip1grL9zqLWc1eXxfioohU
SBg9ZAeWbzYUZSHOTzaJ/KepktQe16+ZQNxDpYwoqvlT1YS6LS+euabgZmdiyGUC
ibsM1URnQFlKisDWNHF/iX//hIxxpEwjGf1wHQHd4G9M0I/Fax2uOd68e7bM/OgJ
so75hdk4kpQJWORNdUaGLspyT2lqiMDx3y/HZ/AtKcjLJ1bsB0vuT/h5KWyiWFUC
ksrqLuvf8WEjBaI6dhTB2inR2m2V0muVoYzJqvWUtNX0pjgn23AvHbaOcLzV6/eP
zT4Ts2rFPEKhkd4A4P6bT3V6dxOK7fy+nW/ji3nRFQeUZ+zcSxmcJ3ijyjOL7JVx
DzABC5lH2zkqr7Nc7zlX5RWveTIZ5V7zT74faB//oGhkpyhnPQr5BLb46YI5EHdo
fSk5sxgP5Yk122FMMCNJ7IRbICVOwv6a4FAgkjkigRJ3fIAimmBDQqir3ksA7KZ8
WTPieou2UoeKhcc+67kTm6qXNIJkVGC8h4kmW4EAM/9LrZyXH3ZRUd1LzQOtkVsn
36IUJ6MkfIUiu2vnE2ua2+/JsoUeB+eQYpVhc3isZ5OYRCpeqoAcNB8HAmSx8cqH
O7xyzDl/ao91B16q/dvhU+yC1kUHE9Fq2I0nNK2lVIuvP9x5qLrxPDER4om9h0pQ
jhvC1ikzdIE6oZr6sdeMd4jxpy2fRgRhFpMTUimHE1R/zbr4m34lxYBPvTOVLCMV
z8J8klQpbWeYZ5pC67C8AkwbrnLr3KXYhf9HmbKk0hxtewUuHJ9kzNjDpVTbjYB6
OpKpMpdrw8EiRMnhgLfTtWDnXZW34v9lc3f9EcBWnVZa20FBloLJnXN4sQJDZPeX
1lJi3csxjXQAtmyVBn00SUHKOTAjWZVVj+Z8RFedrXiVXyhrlOV7JjoofWFUnKFC
dULtBIhpaolXB8dJnGE/M1YSDdVCqmt8/lE3MPPuE4+ToVhWwjdJuHeUAp7gxbBZ
AKz7OFdlM/8/MN7Ev6RddLZbmlEZek0RcljKqRMXbcm3CE1uEHX+izzAItIlNAI0
fXzGu5NeUQGx9p4tRlfsKJlIvt+We5Q3v8gxQLcHC8SMlqh9Y0wYqPeyUqPD/dqC
44mG55HnJ/q2PeZWHYUOJDJM3Z6GsX4A3olTxd5YZHINPxkmoYMyMh7dB9hgBVU3
AfuSd7LTlVWrGawDtu+J84stNQ2bVsCTXord8gSsc8H+Nuzz3z+iJJwDH4OvV9SJ
Kl60DV6MZLVUWGqD/Fs2wytGTZm+zIuT0r+4xYDp4eoFKCojsRn2cisDQJ30zLgd
UkKfnJbZrJRjLFL6EYS9gTSQNk3FzFqOoI5UNXeobc8X+ouuUEHpxPUD5dxL2a58
O6yEQ1ArOJ4dsnRr5L6oICyakXHeZ5LdQdUbeV7RbsoaZ1uqwUtWjTIjI+OOfhww
d26v+j/9FuVE9HCzuhZ6rs2NMFV7LEkArimZdvbAlRlhONaFsCkDetiY8v08XfRy
QGrJ0LMQ8qM6jclRCKDva8yW3dOmXlJdlBrDSZNw6ORw8+tnf7yhzWmKsQZ2eWdw
wlW7yKBD7KzP22ERW1hPayWxSNwpQWbaoJLuzlQsMtN7PahMSHIVXFxRT40dkwLN
J8cmH9xYo0Pi9F0uyyTc2H9WQMDQfHVTZUfdkLVgCJ8e61eQL3OqLB/bW9+ly5zm
IcvnOjPgruSqHtvROdXIfLBjB/a1sJGJWkKE2XeMr4OlyRilfdCntY0/ud9pAHzZ
/Ae4BVjhgaZqxzlody/g89wTQRpv70kg/LZyjl6v09EiFK0yHCSLR3Gp5pS+IK7Y
NKaaCuA6z/qCa3cO8dqyZqzzmTQY/yA1lccOGboAjdZgfEZbicAcV/GpEBEgFwa+
hD3tpzRQbTATB+e62+4lOR6yaxywChlPEkzX2FKwpLLmySI8TtcVE6jZiRpbFD6G
rjTzYXFLERDpr994vIDJExrhGgFsjpe4OsSLz7oTOEWej8eUaJKDoIXUumibjlGV
/TA2Opu3a2vJS3AnbJKNE6sRIxr9dSE7ALRZVjjy6TxudwyuQjgHXsCOVH8bL4l1
ymMlFWh0P1CzMSvBj3HXJXL8VvQMCDoCGGW5XZ19LaaoFjN7+yxvS3CXJP5KfRzf
lb9OU7XaFCq4l65+U3ncfNF2aV1p6eeUVOaOJ22H9x3VoB38KhQ3fxltI7cz4T9a
r1IKYRMtep0GDEWiKpD+9fXB7h9T4SPhk9NSmcpdAcEfrQTY5oyDe5yT5PrcrUkZ
dB5VYMpf9+xlZCyP3g1YNNeH5UK11T/XLb1i/7fcFDq0BjNpSYh7qGz9vBTbtg3F
zEW1q/Y7UsoayyLQpkR11fgRc9PFm38V5EJCh2jBMhos3OmatEjDvfhmt5HMgGUv
zdmBGNUGTp/oEZpcFs/uzab3sAWg1+EhlxtHgcDXKsa8mjBltucWadbOwFDpaufk
pfF4Nk9ihNeHNTZRQXDvcRFMblB7R6pS3NQxnPpw35SHVq5HkYHuky6uJm6MkpC3
AieWABurT/4aiewNXy6OR3IZ6hgNVsyJWBvLkEWOYF1nTBH2SdwH6UbkLEFmJvx0
RN3T2OoScXUHNkgEiejMfulh+0/0p+oRv+QF30Lfc07dsQ9zyM/haNh82jdpKgVu
iRPAkLwJmCfv436+UhWsOg0nyQCAjoYO10XPieWbcvKh5ZaF7kIhXc6Df1Gz8U+1
ZO1Oc/lbr+7ysWzq1BbVoPatwA8+uDfEmCJwSrXZtlWezPtZKe/azvYBf0fv5Yfy
cAPa+Pr4FO8/nBUkZsu/DKfHnNcanfZNP4CvEPwLifAo+ag4FIg8XBgWV+8TGbJH
3Hw2amtjsuO54ybl9fZ3NDAhMwxi35DmQSgpOhZeb/sohXAsJ2ewlsrlEM2Dpo6d
1+TVe/X9iT4Hgrl7C53yOs6DOTDC0QnhBUj/M9Jh7Xjqr5oMYuaBmlzAlzGgmiAy
MyaLnNpfjTx5dxsuSyCfx0+xxz3OgTT9XSxC+bNr64r9llxkkDKVUyTxuTpW91An
80kCFZ52GTYt5XxphME4H4a4QwwSBupZXbSZqMB+/DhZVHmKfsJmvv0c15ORC8Yf
BHSK8R/e0obKscuFwX3gEtb/C2TsSrcv5FW8nahqgqqPLyCSJs4TXoTjBSmUsSfX
Ut8yHevHL26Ny3wn0t/1P/mMEKBD9csSGJ2yHtXa3b6BGYquwMCKnntwh6D6/GGO
s3AUja/LDbWjn+ZeRHwy4b//VTGONxVD0iWfmQqLVMxtuLJ4jnef56zWwIghpAy+
4p/yXI3W/ap+vTwfllDK0xj20ymW+hwiGCf94/DCtwxvkfXIJgUVBjq2wnY8Wdno
0q/JcFaXdkKebL/q3DUj9v3knVdzv6ssVOZdwP7eKx942Dnw7g250Rnr1d73QAFl
tOjLaH9K45Rbc6kBqxsdPdYnixtJLk9sVMMnDiCkV1UIUJSgQXYvORTWMtyp4fF5
xxsn/bz2NWIIF2FsggozQzMyBgzbhhFuCVPXtMH5hHo7tBKRUZWNQoH+0FFCxfT0
Gj4JF8+UVkgDPfYmjhhHZZqlEmuQpM25sbk9247QEnEL8z7YV0IjStsPbAYmStQ8
EjuK3/eHS1F0zW1Qa71opvHQdN4nRD2ZgCAKSZypRZuJ7Be40gUe+BsjSh3LSu0h
90ZURtfKts+UWA3/FaUXrkvkc+fTbL4AWiMS9fGYSAdfpM/WV9r/SoLGVCD85khJ
OvgPdOtQCzl82HNlHn/lNSLJhK3TlpBP2JqxLhmuLitX3TLNwprvIAslbQT/6ZoW
HT9r3IE5BfbYTdfSptiHpCch4VS6yLqyANSPtdP+KIx5uvN73oPPXEX3hAOzGjiG
OmZzOGN/zthBOIPgte3T0PB1AXOoZGgQEOApH+T8n0q6qrzLYwf4nWsQbLPxLkR1
90/ez1r25sbaZ7HSyN/e1SszV+lO6EU9Heb2FY7u1Y3NdDMBGDWefBqaTSy+taPu
Olv5PeF3tl8+7cVbmXQycG08PU6MuuqsPn+KDlY8iL2hS1eD7RjqKDRP3Wu0AE3H
XG6QsmjBbcrC2qUoHVAxkhmBVy2nbIT+vvrxZK8xdk+8hIbhLxnVYeBAkxrGNsyY
dwYoprgw0Jawtj6e6zqpfRpHlPIh7jOoysNIp2fe+YesbymZ2/Rxrsu/WGr/t2b/
EYjcREunx4Qt2P18uqmJL8XSYgNzJq25O/7tBGHYqzXLYSR66jxVKPi0isfwntgR
DlOtqTz34Us1pEDBRkZXPSKSL8WZWvPFLtZ7Un8uaSGKlAchrL+mxUl5VLntY6nH
gK6Gf75ONcCPhoefyFBpC5o9+7aOjQvoyggAQGror/W3cBWk62J1WgJlG+joshWg
IM9wwyQBK+1smirN213s48YNTJQbnxKXmq0cfkgW5yfDolzrMU6itjTzfvWgRTQ+
Zvpy2fZ2HR+WVAvlB3dL0l8QAFv4dHrkElO+XKI2Rj7wLU9lZtPwAXuV4hOqfeAV
6jbLlTSv8joOC69GLjbn4k0DH+9mT0h8MIdj5kLNmcuLnjofagnmYOaWW+ZfkyPy
xoAAC1ncKuSd1oamMnyN3mTpY81x4TFd5K1sfUAIM4BP3wJBSt7JbfVwCQZoUqLH
Kjv+HUn+7ev7xuNnSOihbLx9bLT9j0j1XaI2CrYRUGTROSAadvR4z0hXR/Uc8bRW
Ckun+r36Ij3+fDuK2PFoXRsmUstCChBW5X0X5pmu+g+fzuH2CUQdcniniT4mvuQM
Qji4I8Rf9qgfpP6TLLomLuST9exjLrtkvyu6Ne/ZrIuggX9YmuD/xMWU2hfhaa/6
aV6A1xKAhCUZlmXnDThA6EwNM8VIZs5BOMaO2NmFqb7T3de8xTHz826CwIZJcEXO
0NREdKllPK8IsQMQIHtMqi8dgeN2emeLDY+rT9TXgSoXO4LyqnAAARyLyUciO1mi
5OigmZFOOJWkSHkBLpAEsuPvo6vv49L86GFIgvzfAM8vw8J11w/VtX9dZt4zjPz5
+UHGTiNFgpj4Rp4yPqAF5JGbPBtpBGz34NtE5UhoeZEuLWW0kcuoJFXeGUlJ0fJq
eXa5Jcbl+4jNK+8unyo+QXPobhTicasndzSRTVQsHgHZ2ka2ubNbPy6y01sqF11V
rRVlDMM7FLKDYZfH28JZNyy6m+IoOpeCXLQFFF146j5Wv7hW59vYAiAlHjZDic4Y
jOim+T3csK2yi/GvzaXxXdEaQyrO3vR74ZIMgN3tuNh6O1DFipWru0wi0nfmCr+X
J3ei4Dn47hLVUuMGr8NXPY7uwJaq5zYnhkojlAAOR6yh2PA8y1momUciMaY9fK5q
2rr+9PJF0MEtdjTcp3gYbWMLYOmYaAMt3f46I0vHsoOe2+hJ+02quO+b0VzPoX0n
FN85wmwaHY20fC+Lo60ybl6nBFy33Dg7LSLE86vlvQ3m4+ecx0RB413dxNgpxnLD
X3iWZhaNNk43Ur5mV3lJbseqt5xAxYk1/oIY3WNhoLg2Kd8yE871uwdNtTQKK7x4
3j8btKoOqin/G2dWNbbU7XAah41tuxAIRPtTBsOP6KWKgfE6sIX0C+Xk5enylr8P
iK2yJyIbzLzOtbay/RVSgNoNXiHyx5+RcgEVyiLJWmaqKbXD+yj3z20D6UWE4K+E
S/GNLqlzf3KjCmTFlkrIE/3ljV62FRVoT4gjNuaZNMIb64BMJTzPi4wtYDIez8lP
VweP4s9YmV4pKq/Hpdz/kWOwF1efYWg++MHck2/LGhhLt+RlqBNFFnt9LpCbUFL7
UeLtgsCz3OHT/l2J+cibQJbng9rh4EiizhKcPN2QSVrFC8glqZFH7tRoo29Pu1kC
ukwfFqChF05u0ueN8/F7koGzFZTPwPrkUIyTsAWT39ZNubsPlH5dg2gtcSXsY6+y
1kbaKPOObKDEkyYR1tiLVLIIACAHNlWJqe0XHS//kmzNNrwBS7UetN/1l6uQLsh6
x7lSMucs4FS4+iAwy0Rp2owRvFNrNj91m9AJdLTC7CHaopAOlmRbDScszkJ2QSpM
BO1TvEwwlxK7AC7vpvrgVke3RTGIkRNvnSJtD+064yDSg27MJ/O4qK/zQVvuzMLv
29YeKcMEclWEKIexuh7J24gZQxhVAyafIbIa/Y2xS18I8EBdIm8sqpWR6hziUAse
Jlgxmtw0T8QMiF//ejI1fUh83aUlG4hO6d0bcXGjBhMw6tdfR6noeGe1mWHmyMJy
Jj+rKhhIXv3kubwcWpkO2aGPZbdRUr0etseZire7Jj1q7fKKudxZZufeEO0jy3WF
134Q8CfCPBod+vf3MeeyzzeP0lvRaumu86LqzzPTBwem36k+mHiAGdZ7/IS4cfYc
jc7rMLmEWHIJdFKlpsgQ+GWf90awXHVCceHI7QALfAv+dqVJvGN2F6eNV1bBxWdp
aFE60uf1+ZKdTqqASM3FNJammXmnQu/5ngA61cSPy0frLpHXC+p0/jUP/5U6qJS4
qqSznMN6XnY3cvCxKFIeBJF1ZBtiW+lvk78hNAn68R9eJB/slXhIz9FiEJBSbFdh
nMShVP3zLjcS0OHUCitzcBfA6JcgaM69vc3GciDes8gqXK9S+8SVZ4oDeA2QmE85
b3tQX/EPn3xOAeNJ1sb6c0z3nFAgwyQ1Y25oK9/UaI8qPHZoY6Ugm1AG1vyiAe2j
nmFThvNk36TrSH0BAwHglKFwE0nfgRJyu9QVDbaTqIwsiy2HwLJq4dUwW+Hq189b
8tqVaN94wguJNQiTEkROElQm3qPTJFYCw96KMWjgGYBJ33pUOY951fns+XV9O2jW
7hhgxd/PTrpMX02Aycj5jGfy1JjYK5bEGIktRXydiNyueAjV1tKAKxWBkizaR0XC
8/S6v2H5udP/chUspscCww==
`pragma protect end_protected
