// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ZcQYC+pO+7Ym9rBxtpycRBZaQwn0YJAyEcUHVHYf7iMxmbWPimNOaZ/q6QJY
YIEg72EywwCB9FNsZd0avEpabg7rAkUfE1YFs2sJ3Cxfg84UJFhg1iLtg82L
vPkjb4HMiIpmPueMFg6IcL+KiFHBpSMu99D2p7sKTO5InankTv5ck0mbdyCM
Thj92kvwoYPQswWYFyOtl4tiBAYyCFIVaZLvS4FKRJtm+cw6oodB0OIsm3Vu
nbsLFr0G+vm65GjW+r6UHZ9BWu7fXENyRDNHh9nOrhZ055oIDgSOy8Vq3/Pp
LNIdCppLsuFLVHsXlTHl/FXEVPD/x2oXnduSDdOS/Q==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
hseQNWnx/bO92ZSXox966y0rUn7HaoRdGsO7P/J/acXMdT6QocBRfQrXAZ2F
CAVNfIdTJrRsLVlLqjFLpKOtX2TT+wFgGDfp0w/CKP2gm2mdogjfz2/zEUrg
KesNHs7XTrJ6NJlyrkssGJ+lwG9+b9fCpG02JNiKDOomVK4x1PXrMx4hzse1
Api8GGSgqDNx5w4YQNHWuJobaZtgVDzbQod7J2bxAwOkPusnoacvuvKExmWJ
LHqIFjYEbypu53DrxzzH4Ce7ALXKweFot0liREnZS8ni++s9CUTGBgpLsEA9
VkVFAp4kRZtcpLR7Girdcs2BbZWvLmYCegeRYDk64Q==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
AoeYEtHAZhQJhp+7IYGH8gqAYrveRet/Ov/+HRTDb9nVX9zn+gPLv8ohNhjf
ORGN+lGrFg174KbO7BcKlAQOcgfWdlFX6uFRvyL4kpUCuZmHR1LAYIvSMPNT
C/dLIiICDh4m1HnT2nAD+mwjOF0tphNJz1XL3NhIbs6Svwj7cIx49v71cTDi
cNX280jpvfkljPmbO+1jJKBFWleLzXx95NPL8bemNKVOkL5OZAPf66X5aJdq
B7x9hlm977Eia+PeAMFz7mZejuSxK9Q1lVPIwryjtcG2KXuVOgrA3AkRpxIZ
aSk0xtNRuCph0wCidyPGN9M2EHNJPlq82Uq938U3Zw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
MxGaszJrnBFlu4aWWPe2cFDDFlQfDMlNMWaK1yS2zzkb54ZxuKXpbATZEMHA
YcmpIPt99Z+RYmagTrzVk3TeGLn4rtyhVNyF9RQnFQgFi9ITUOrvQzuakS3X
7Qb/i+wEb3ePBmC9JwuuxniXdTpD31/agwx39WaSnwFKH8GytZs=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
DYbf8gXEO7pOxgbTyYknGFK8ubcpU0shOJB+e/qc69Kif/MM01oUgum5JkjV
zQ32yOK1KnL3wvs6P5we+j0Qj321okxZyW6lZIoCF6zzT2VfwiAsiJjVinLl
ekqZF95yIwPb/c24KrGX1c1M9s2bPztuY+aH2ZrRz9FZtqA0PbFry62nG7h+
JZ+1ltpMZAw36NipcWPEDkAhOLSwcjNV3opqUiyWvmMbteKagtZjMET5aQAO
eMbbUzDdogLFQfH8jv6vVujWNGjcTxCLjagvWZp5pzxEnehrgjl+XOS0lKjc
zn6FNh+f81I4mnPuFW44hncb/f81h0ohoGR8kuMIRxYoMHx3W5HhPT/AOCaJ
iLK63zadL22aaaH+VTqtwxY9reQpEnzb1XDnkeY5l/sEV9meH+lqm6s7eV7R
2XvDhx8j3axlQ0pfklgT/1yZSqgZyfysheTse4L+nvGHhanrhMlrKAK7a+Tx
TbhH5Vn+8DuBh8nEKIIUsTGhXyn5nWte


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
kvhhnHbf6NjCyVjks2kBbKmgbbNJqJ9OUyNgCfoNzbfDWvEU9BzVzy9ATdfZ
MfpldZFy4/OlR3R+fib4c0SifKxrZcxphcvVmOwTm2F/0eHHyfW6tktYhPaH
WsXj/DI37tPltk0YGXVrwfdgr72toul5mSEE/8GiCa46eQCs/cM=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
I1rnBVFbxUvHRbb0G5Rayuql+iCo5ySIPD5IIaKhNCwn5KRkOfuXvERVZ3vY
Yf1/UOS3al5TVSWS5/bjjqakVr0pB2Vg+B5ySmdTaI046qHy8JPcZ97B7kwK
FD+ybiZ1I0rcRTuDpMq9+TEfxvBiVmTp3XWLpzaEvmoS8S1YX84=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 8688)
`pragma protect data_block
z0k0Yls4E2zLnMDS5OVHVLwoUoZrgPILQqTwY5QMGUy9hjUyl4HVamP2dsrH
l8+odSI18gRRJcvQFFUH3IUI0Sk4qnXV+qNTu4f2FylgYC3Bkeh3iFnNjFlr
QDbH8r4H6AJYtnPjNX/ewwDBzT+hMwFT1z7Vs+KasNaH3IvToDBUm/qiHfE1
1kkFQKR0NXISvxld1w7cMwmO1vK9hg5oBdVoilj+rMheVE2Y1908az5RozEP
Oo4fh4rKJGTnl0Ija9pMCbhYfrqpOGPLsjIqZz6U/ffaxKqTrtF7FxG4fqKB
evL35Zwu8SajtCK3l/bD/v3b5GtNjK8IpOxg8RvHBo2NjBoFwb4QBmkuJeyC
E6bazFI8Rbt+I0akBmDUwXJesce4MLQZ0l1LALT43racxw+BNLhvzDrav7Pu
LfXvQKc1vIHVwvn+G1+yWtnX8anO1fZT263StqXa5cpAtSJG/JBXDzfQUqRy
ek9pzlYzXWQRzDXpJ3B24rCUgB9/HJbAxFobw5tAOXF19cIOauitAVvsMYkj
h4Hk8EFBCVksPWGkNx1rthIdP1w/jkfu+QgWNhWS1fmZ7NEm1iJcVYDQHt+C
XZiKDKo8q/Y7yfVPNijkE4OWdRDdZgtcpuc6kE4xbBgFCMGKG9t1l05/fDmv
4LZSxwqQbhJtbJWoRY22dwcJEhw0fx+SluvF/dhAbq9PPIa5VrSCR5fP6qR5
MJ0/RMM6nbDDN/fmUdp/nVNqQ9TbBQaIWwXIpAFgoBJKl8TvlPup87JpcMKU
ZyY5ht5Qjvw1bzSMjUZP6VtPSsuVmmAm6/rCM7SU9MvuqIdA6g+MWQq1iWLT
VUE6bD23m57NZsxgqHdNOEuhsm8iDhlWgOd+Ia586m6MBXn55f3VYJPiWWJM
NUZDb2sFByj2GIu/EsiP908t1Y+zI7hlADMwAvmplE2DovxB5PLEQMl5KbVM
1lJlZZwRdGnBzut4vO6SOsAtOjMR+3xrS/hbCY9v2Skmog18dZ1u2QwrcExE
L39NknoTeIO4ytEsg5n97X8PufXO5E0iGErNO+zptBlsiYf0bDFN+wD3dCAs
YOwXspL0Dv6Fd4OW5PXNV1WnOqejE4TJXJgBzVpprgTgIVyhr42cLkhkrHq+
h4Cr1fM/GkWeudHXK3V0JvJc6sjQARgNQgJwWLpT7lJFH+pvVz8LvyUts7Im
cFKg1q1hzSCMQkGuvcVg/IhlBBiK9o5bnMBJ169DQxCjxRZG7g4xf1f1iw74
xfwsNbi3WjeDo4khA4C6Ycm35Mgf/T0dKZezEtKl3GDVv2p+y5MIwwB1cvKo
bi4nGvsM+aJGWA/QSsLG2OoNjzrWN7l/3bggBU14WYGu9dbdvwe+K1vaxCNH
RJBeRkGP2mxER7EnwKT6QBoQ/NUsRq0mZI9knXth/moOw0Yx1SloAPDXrteI
UoC+DAM1oGXyZpILssqR1EGZJInc3iIbwPxJWmnEugO+7ckGq0VxaSnyr3IA
zu8VBmYCfDIyWzyAY+M3FaCZ3/aO7vCf+VNPovNKQ4AAOgdDSbhnhEWb98px
9MYLotFHvN2gaIQ6JV0cKeUFq6SioQuPsbK7Q1vdtQeU0FGcvyYinEz+Bu0g
hCZdUUG8ZLnhovJ5P9e1ix/TJHs0xx8l/Rw5fTC4JoZDPPzBHcpwx47ykIZc
svtobi+vPLEj5QHvXvT9A9OLjilrMCTsdTEhzOPX0Wjo3j4hoozd9aXSJ2Qo
HbcHwzFRXXCE0x3rulaifYxWsuaHyhBNkK4y5GzxJ/sRER7OdnZimLtlpu5i
TaJPegmcFxLSI2uVtx6JgNx6E88gMVEUZjhN91RlzwfqP/x9npxHlpHZgpn0
NMix0dkuX15J69o7Z4+wp5nuHFMn7McsbciQ7b1ck0SGIJFFvAXJ6YtcIn31
jvWEiUSev0XfNv5vDNQ9GUPDIn7QLyrSbuoKvvCMvrQLNFtpid9GFZ28m0Un
8Jqu8ukinUQmSG/9kIY6iY3ccAVM9zvSSRtfv5KbAp9H+HlVZaC8GMkJBGkR
ZyLPO8pCcPIDdnsZloI9xTgop6+wsBSI36UxtgHYzzlYhlftX96bC4ODlOcY
jRmb5337gnAyHZxEMqTss46CH4jvO4jiuMJnoWkoTuchsDGVISZ01rAzIH9u
4AiMplkLLpzm/arzpYe74fSSVviXslN8pR0iambqzmgJfRx+uIqziVm+9Jf0
t9vUkhWz2UqYzOqMvxP0yYd+TNmxQm7D5nkj2paFx4wce5v2rt0dTU4C7xCW
LiiGillQdW3WAIpsiYFXaZ25vwDJknzKoZjHcVqqDHMaTpqTXCL7cs0lWW33
HZM12AWUhnEaUi0kpXfTqFG/xQFaEkqQlQMOKmwUbNWXCBs2oUEM/jW4xzHr
5R7HcdDHWZ0MnnTIpB/0eg6l+RH8cruFn+CC7uvuJuXsjRgGGPd/oCabAzke
Y0ReheM/iErbiDU39Rp8sA8pCPpUGany3/taN3iDZ4HYWaQt3mFtDwYT8FLq
71OpKjkwvhI7aOrdbk4gca29wXVE67ZiU3vP6K7fYuC5VklJ+odZ3McctXd7
IpM3Ck8bKcdKoOifnw3zVI4BjJBPRTSWvTc7EwLwnbRP8/kOi0QT0DuMAGf4
DlPX5HZxvtZaep9stY5UIGaoMd4MnfTVZH3ywFX09nLN8N+5Gcuse93Usn6T
jtgaT5ufOOETfT2MMTk558bhpCtI9/Yy+06KS1F6TmQZcv7LQWNqemDusLFI
YZt0n5U5qr5kZ8VOduHETKly22J0IIgd2vfxWiahMpyX41N1nRBeT4Opn97+
cqv23raBzuN+chj3UrTqX/1hFcS9lDusokYlaX6X2z/SDPPIN77u9qEA+XG5
5lWiCh6URT68+fL5QlchYKGNZiVi/4wyqH3jhhl7GexUUHD6pWJE45COg6xo
6qutoxNTERxD08/0HCCw1TUDWdbPq1BxNgh393kJ/J3nK47Vmx7bIXOpVt6A
myu8CWvMgIzOZUspncIE8MFW4eGB/kmc7WQEy13qRXn3JWG55iQac/uizWeN
BwcrkFRPJbKQse+lDwk645eI2sbxgzSUodMDY9J/QNadQ2bH5eqQXTkk/ZI0
wARzRsIg+ESSLlMpCz6TSpSZnOu9HGamy9KpJJccK3+XXgpZZYfwiHLi+jWv
02Vh5BIzMPOS19yEKuQBPbtDkvxKXqsdgbMGwR7izEiH9McjcA6bMukmbQO+
PKvoyQY0s+zYYvMsGeMKEHL1eV/5Qjf9dKSHcPULZpC4bI0zrUKt68dTt8Sn
xwWy+uojQXApBYLoFvURHrcGYhYfGqIT40sQy65AoY4NmKzGGJZVZUa3g4Xi
7SVvMVXcWIITgUo+RIy6IWm/jDj2VKqrfvJ9uD3vP1FW+q1T1q8WBKlRke71
+EzefVqaeZ3M5XRZ7EwHf0B70mbtkzVmcjCLgLKEnR0xLnFpiWVfzU8aLxfq
ttdEMayeREjNb8b5gZehAhzBPe7sRTTIDLj4Dd8fuf/Qc8W2AA/Ysyb8BySH
8gkrHLt0NLZIiJf/Pkn1POFnJgW6QfGi6N/vQ3fieRrSj8OB50fjSB4fD1VA
L71A/lfKRknOD0GitzU/diuXeOSbngTWtpn8T54pFQvAar+dTUoZHGslnrEx
34wOSc1e2G/dHE0zb/IVu2Sv3DC2xmC0YThEOQ4bASic5MRFWetWLPQs2b2K
4tY+KXd642syacDSOrS8R8fYmRUTDFwy5VaQvBLB64PJzhkBMeTHATqc54uB
axr1vBWK+XUjpuj3/UfkhqPfj3fPYmQpULyILCWDsiwnNz+AbjsPJCEFbmg3
KJrudM3SSGyECSsBAlUgzVEoAtMMZk1h7CAa2uR60JgSSidJOQrwtVD8kgfj
qENILRl0YEvosm0CFaoYkXDRC1dat8eAF/rC9KGeu/ju1e7Fd63mQkic/3af
uxVbnR7os/RjliupVNt9mULaQzLCFOde8vI0ngTjO6/cs8SsM+w/4jMvlQq/
oUCmuBPPE+Ny3OZfVsrw+z62rOOUpT3JgSa/b1Y0yaoF2PVY7idFVSY2n/tE
ikDuQVT8RVVNqst++cfdNbp5iuBotbZKZbbeuA3Dmd2WFGq8S5ZPW1KKZb1i
pthVaeavHW5Ko3MNspRJpiU7K8qbuT7TrT2nK4Ua5srY+PT9PBbSTICRwGyM
FXK1Sd96sDGt4j1Ea3gpk9UmWyN33U7dJOn+zFMFaPLeMmMk55xAmZUwfTtE
3/XjWq6V86Q1nS0U93XHp25CNYwimYmFbi32c+n8zdl0quojZiZwLiQyCea3
XyWQbkMUstLcJV/NcpRv0wfp7JpoSqtLth0YwSzCi5IBcavQzp6Dd10R9vLg
h72BQ39gUEdLJx34tlRqiwaP5LfQ3ZuhbHMCQdcjpmLRgNpH9vIVCGjDNAiC
H+F8vplyejUBK3InPGfFtndKgNsM+tV33xLJfAcHWOXJFmrM9foQ6LCB/XQv
w/Rt+GU2o3r2SiG/cWnf2AW8UCcmOFhsDukoVpx2XCLPxcVuCEybdW63BrcX
+STIbdEPGOIGUN9EVKeWpmfbR6AaLseI927rB64WHRCjiG1aLuGG0hR5liR6
67p7UfiiZ0azp411yF0WnA0HvNXDjJN0wmm6khnFZzz7LPbxYHwe7vRDlfIY
pFz0HAlSXpSMcG2ZqJKT4Lgh2vVnFa5IziFM63GtRIlWFZVcvZSmOP+YU1FY
N5625yo6Gyt7oOhDBegxycvuZw7WNylbY8l/fPMWquWYSCzOPDzV0rp9cvxg
bTCmbOPiNreK3ZFUIe9WivDV8luCVWltH6v38bLZQamLRJM9Oowq3LivQA/r
r2jfuYo5J9Y503RiPL9lNs1jUMXTC18CeReMZsOTglkLdaaj5fk4lCgXs7r6
bv2VvOcuuzhGeaga1ZO94kO7ccjTsjjtUfWzZE1/8ItDDEsPXFjt3m9m9dtz
QJ9e5QsBGbCbdShIZeIYl0ei3jdAV7cNIhPloMQYndIv/7ZNnEd4a9CkxgCd
dweoWY8t61HbZR1cc/wlpH6/Uu+mRhRFmR0eVcsk0AGJjkYHiHXiWM48rwfh
kREY+y3Lk5L/wl6Shz+iDX5DJrY72C8lC1sLWTd4REiizeRyPUqUu0+MgyFX
FAyTmqJqKgWjnA7r1VRnubQYWe+LY8ymOFpC8MZ1qh1Um+RUnRb4IXtKmXRp
wnpPYsqDl7uvk19rY7T3dDXh4SRRwSmDAbKPUJ/lhIhI41Not7pbHOInCDHN
5x0TA8sbXv7JWm/Epvs00ffHhgwIllhVm4JUBKRvbbMBIb7WAeaN4N4uF5I7
m1lQY+iPnr7i5TgTen6W58lXfQ7jE++6uecyxDwuOHEgH9bAMyctoI8UeMtF
oHn45zW/1Xh91mslat5hAwJwmIOvyQYRsD/RgvcI83tXjj+868frkmNDAPGn
Wy4TsyIrkyUR/khfvtpwP1kHDByinlMotns1tL63rZrM9l9uESwhwDwODvp/
CEtA+vSw3m7kCKqAaq5EwDgfjVRR/1a5MJWJtSuWvVSryR8xUwNISSleAhfu
OgXHY5mhOsJDifrvIoW4LFZYYQ3hcIRzNN572D4K/EnSuZPocQC5wH6OOtwq
lPt/VMp30UojpRhhcqj0kke5SXbmh9+2fFa2QlUycO9ODos4JEbX2v38zNrX
PhaL5/1D5k5BfpKiv6bEMCqKCgrpNEJsXilDDuwQe4enJ3SQLjyGl3lpznLM
ARtn2ZtW0ZLg9xv5kualYBYN2VMPTHH9c15GoCfpWDMBTr7ETkHKgI3AeQXL
QVxJ6YeZoX/ieXmfdLgZkbnE6BlXiBwnUiJcXHc8ymfelehNQkNvTI0tEXKQ
DGV+PS0QncRo7bufVwOThn9j4GF7lCZzQCqpgNw/FrFCZK/jxbka1ZqFhx7n
upSLsc27T2vzkopuEdWW6eF6/FpUARQUvVWbcApab1oEnvRzwsz8UvP5PK3F
RCJfac479SGxrkwgGKIkf6dIJTBIM6zecx+EcFTHQLFupX8zrP+x1Y+R3RFl
MKi7vZrbu0RftFyeA5KslhI399V3x1BBQsZV1bWhFQRuAjoll8O+bZUuFyYB
N8LXO53X32APmSx38ObkjCLrVPxSwNAbyj5nZkeBwqXRm963KYHr7GItmrp8
ldclOm2L+nYGQaa1KEKPHexKShcQ/QhyA/d5EHpHwswgI1dEj+pkd1buUcU7
QoP2P3upEMfIgRI6Gt4UU1wm+Hcil9mwM4TtO577Fc2FjGJRhTdFTtnR7jTN
5ykqZFZbO8lmjbqSraBM09bShuX+oL+X/35u46GtRtLGA3yeG6lyC9nuZR3E
2HZKTMJA4WkUa5n/gBAhcZNHr2LLa8XUAJl6P/+mSCdWJdFSNmGvZLoOPDa8
Au7x5455T7LlpiXGK6v+Tf7DL2ld8UU1XThBKdDufkjLu1XCEg3J+gCyuvRL
oqXgAWNp+CTZPiujbOti91R2hoH89qCIybVFI0P2/rm+on6R6KqQfXfUFBKr
dc/9uAKmsNzdOO2C2S64AYyN9YSvTfcy9/+a4xCgAlDNzfEGiUc5aFPsTjTC
G3bAqi0/FDJRlnsrSWtZAvH/cdRRaFUHNM0ndQIFMjY93stvR9ssenjlvl1P
RmFYluKNL6Rc0fvf7DeEGm6qPZ4ldD6EQvpTCqg88rDSRaKr+/o8lXy0ufja
N2w5yYU3KJUMsru+x8g5h0ejD1i7boKEAvOExLIOvbnuguW8ADVsolJM/KFz
ip921eD8XQU2Si8AYJ1tfoBrQoKkAaOEfr/qJLXOJLNy9QdI+LAiJ+K9tjYV
2H3G1YOCt2inffG9qaZpU7uLPwxcKjwyr0gZJj9X+KPIrz3+C7cmDIaPvdn5
88yWqRSOPaeZuUaIWqJ4NT4KthlJV6ajxpQjGpzkECQt6uBQuuAYLScEWAF8
x2yAVCQAThWJ4mp5OgjSt2SkbDxPIoBJUPIeHKSmHcK+pGhmEnLODrwKcHN5
orVldomg5TsavxzRINFYnm1LdDg5YkXwkeHMNNOQVa8ajNjmcJMFmmiuCDYg
CFxqT3/q7fPhUFsG3IsPskVqIJwJxtTU4b0F3lz9fwzRdCmy2LjEtSzGgrpP
fJSf6rIrOqkgrTI8bbLUW11bTme36p16mYZ6aWe9VPohdsg6Av5aOVG8Xcjw
0KJRsTAY4TOVpH6T6FAGnt5efs5IJ0WgRZ7/TY9NuPyzglHTUUdFaIh2QaHs
0fRh2k9Tm4lsUcdgmqdyNssexdch+Gi5Q0fK/qNh+VBX0Tp8Uqvt1yeYx4bf
GhMbEPvOFhhvFON5thRx9Nsz38NWLvhn3dKXzUoYrWaQJzemFRYutIxkq3SP
C32IjX3yffKVCiiWFrUJx+8YNImh608b/XtjW0nVmjJ5CcsSh1KVnrfhSGCL
RE9VPIortstfENIbjRGkHtSh5yjX9VtgckaFpp8GtY18UkzVMFJR9LbnvB0/
F9tWcgZW0Ypr8UOz/lpXier+/yXoc7TcUYBxGo+D10EJdpRLvFv/SpYqVaiY
wDVOgrWHFR2pSS9JpeHMI7xmcMGezuv4e3j6ZsBstKmFQBtzvD6RIKoLFdNT
gmxFBhZLeCM4EG5JrLu0dOW3sCvKVtB/kqs+jC/nlth7cOc23oNsQe3zTc19
MTtXnhcbSB7VT7bbM8SfEsyannM/tOJh19pENddeJ/waJhNMeCs45hGYVI0+
0o3dAg3YPoY0AuxV6tl3oK74V4MvDURRui5F+88SdrBlq8s+Z9PRFUj1apZa
N8cpeaEQrz2siHHClqkVf5ySdR+Fri6zOJ9B6CRrnK+uWLCm8qnhZHB8Lyez
+wRrQIxj4308qAf7O47ieEcgtchPybdQjThfIz0CIsLfCI3RRhmYUvOXFyEj
3QbYjGl/SFyyEBHNxt2LoaDmK/b6w/NOlqyDTOhtRf/GRIM31MydYuDsMQq/
Wsdui2cPo/NZPj+53Jvk8PMCz2U0cMMM8J1yP/C0vHr7XRcTtbBJAoJw6GM9
pxpIU+WpdBStfTxdKW0P3rEiIrShHn9fGnPWjWm3TPS1I6TksHlIptwZYW1q
rNISuZOdANC8mXROi/suweeoer0OFB/dFbT/kfevK6r95Gi2ctoUq99dkmJw
lf1QosMRc+MIcC2m0hS8fCqKNjnU5zWistAYWvIkyvx1xAinfE9wXqDVhjJi
C74zCHSq3CVX5QyyQlAR9mMzDWtWdHHlv+O9A31h9VCJNfb/ZOkKbjOjBeYG
MmoZa/EiRgPhLdZNCHz/s288nT5KSwKAYv9JbFQmKti8wWYjs2VGK2iW2ZIE
ZotGt25eYjlOV2VeLwd1J7PkR7Fvru0YpIPM/b6XobhxctONTtVWAAfcnX1W
ehWlsaLtqGZlJ+X2zLT9KNR/LoxMD7LWiAKI5UEN5XdU9zOWHjyzXFmmBTmB
UG8GaPYaS3uPcW6qxe9WyW4USNo0j2+k7j7APqTWkfcIevnRNLi0JGhI2HYj
gDGtv2b1FPTZ60wMck9HdyoyL39HlffhSULCeiBNTk2NA1Bsb4tMB0l3WVRv
wbLTKpiNWaK4tOs3fYjuTYREkX4HsoMhgOB90g0bJgKl2mp0O61gxa2LhAiq
qTuC56rGoTOopkRQIPFLx/Kqs3DJbds67jOM6VRob7yZH4t4AIz0m0xY7Mut
iueo4lGeAgMxGvtJ4zQ1aoqNsFhn4f2ywGvCOpvWyfp2BN+B7xbg3oBamp2T
XW7R6Uv7IIJo+4oEmSpwNIZOtB9h0CKiQo4saq6pPyRgixAoZf+uDXD25Uy9
WU0fOGiFIRAvJHElvYZEHplnZdhvYk4SLoMFb7EseC8TtsZ3cj0Pz/m0WO56
Ir4LBh4Tz/pt8ZDDtAZaHPtdcxPHc+xybxA1GidN5q9Gew0dY+dKR1Xdsi2Q
SdOjT6P8yglksDmIUl1QKaw0uLLpUFRNinugWyfcZnkbX4cNAwhuhYM6uOOr
JjMJZnZaAxSfKtXmPR5us1+J/blh9eQ8k5wLELPataoYZRWEKGwItMFj3yYA
disX8bPo0Nxs1y+HN/yBsrvpY63GpQ0dJEl8aFjaE7+NG9BrEV5ehasIsiS/
R/fw/qtCQ3YhgkF4KtHDeRqWoee+L4YARXuNj8HqGsmYYVmy29Wg23Wcnbwv
2TfAtbyEKK0KR6CLusXbfbHyGaXHXQkmyRhvVgJKobUyfmvYRaG43iTJBn1p
kzsPgybVwqhU0jd6gKYBHZ0XlHUwsheD/MSofgVTtuIr+w7pVItR8IeOiXZm
MqzKzgAC52znYHPN2FjAU4pgu54hXdtYbvypI2FhQPJZpg671LlX5o15xgEJ
a6rLdvE0agBPQwRp9Zl5Ykx709ENi0o30j95MlfvO1DqjzRpUjGewdbzZmA4
97OUn3cDYMaFdeupfYZQtMTvgbK3ZHvnyrLKDjTGIAKNF7Of5ojolHtGHtL7
SPAMUHOKm0l46lp+iqtWgy4bJoN9i5ivCdjOGUZXTdCpSOH2nin7FVWnwJ8d
CuInPPF4D8YYiwSga2DPp2Ys8/qhFaC4a12PvhS2lHW5hF01TukfKVDKCYS0
ACc92pPPMGV83fBCKax88+zicoxmpLTBo0GcgYlta3UFT4/bHZu1qwaxYGBs
Uuei8kUk9MFlADrU5Bu/gPS9xkfapMO7gm5ydEO3TUlDEajmKVY85hESp7Bt
WVOJhniNSVtXJJG2f0yi68qphhIHgoh29+9mA7mdzJEKOJHVpbz44HjCKVfr
njH8KvroV1a6vRJLUbzMy5lZobdpqdwcmkApJ0/+UWd4oO5noBsmF0T/WLk/
IT9fzeDzoImwkg/N7NeOOlsMj6qVA7wLiMRY3rZnSNVrneZTssMu2xiBeXlT
UG6WtjfMUuTUdd6fIKmXaM5a/8csT+ZNfCTMHzd1W71QoO0QM/0xsemaPIaz
XVneL+mzidfxTWQK15fXMNU9e103Ut7f4k+gL4+I6E1GnTggqwQcl+titHEO
x5GkYusMDdGnTlqE3Zj0gAdx0lEXeSMaaFbiKJzzCQrotjNfYsNHKt+3lIVy
SdW5O8nankM5R5tYfJTA3UphFWY4ZwyoqsrwUd8Lks+6KMvW3qIvlROXV4ro
NyTIze7lMGaHX4RhlY/2kFQGY14o6FcycAtAaoWw5ruzss5mnmxDtG36wj8F
7znabMqAEXBOwFX1otOpXSiYd6JLcLAQ1fuxmslkYgmOSIJ9o6V7gFW2BCfe
mn2deyGKboTcc68svUApHHBO9gymdygXHAJu0HxvMQ9ByS6LOcTy42MJLrRi
q76m5pAYo0L7GRbnDQvGroIKsdjn7cLBSzywkBXn5c67l5YgCdNXdNq7EspP
2Ty6McpW+L+S+1sZIYkZD9gsVjUq+V2WPypXmI8rvhBTsEcZJQmDUMv1hgKJ
DMQMW9OqU3qbiXwMyInpW9TFZf6WstgytyHwOy+fty0qIvzmlkWgpAYt1mbs
oi3J6PI4ytaD6HWxftviaEEfplRxugq+YXmsX9MO4Gby22q5fFG2g2tuAbeE
L8ByfRGFLTCxosPYgx2Xkio5gVNhqkw26R7ZnYYPRkB3cEeS3xMmjDZbVoCA
Ln9k71ghwMM2SZvHcOhcyLjlIJiP8zZVExmvqds3Tn/5IVDv+S5AMe97ndJy
eq+06VcRIeLMDorV4bVcTuDMJoFArF5QzaPcBGSwtUAc2B4z27eKByV7gGY2
ePBcGB+7jjWgWfmLzJ1CvXCgBKMapwLt3pzeeageSUPe46IQtMcgtmYVfUNY
RXKiodSzwZA67Ga7/eRmZhOAYzenUSbgNvlxh++3BACzQATQJgdb923YzK6O
dgETCsrbvHb5rS3dhDXUCQUmpAgcs/407AKeb3nY6LQR3saZC2kY5s9AOfJC
H/OZLnzHfq7wezPkPUeWOUbLwWgNLn6en+yFicRtLMT6mBJBFyG/uNHgv4mF
cI2oKZF8khBtLRyZbA9BAdXc4sra3Zc7VrmmOmAHueXC1gwUfe0wDoJBAvQJ
Up4HKzeqWYSqJsnbYoXVyPjPgZBf8C4XyRpfko5X2WiWE4caqZf5a6AOyubO
RQaumfCYinKSP9PVZWu/XEVag594TQOed+j85KKgKRNopau/oPakygVeEus1
1hGOMXC4/vmSpJUlPDnGd/9w14R9D7s4w47DDb4gjJLNxGbvc+H525xNh5Wd
S3iMuAdUJN3w523T5mkxo0rQq7pBi63gj7xQmLypECJAfFvXmxSo0bl+XTnF
PAZ89Jw9xHa0rBXo8TSKf1XRzVkLe3MZgfY1JJaN7ZEnUzrVAV2eLwjsDpsr
EYIfSCa2IhBpsK3LhahqRFBRbIzL+s042GdMvHCNtd5t4NJ16PkQGFZbdJAs
RqRz+sS2AojwKxRNm3VG0fW0+0Mop9Y8efDrjvoNjynnsUVD9NDOUA+jycYw
/FUwA/FdEu40hmAL5/sAL6vIzTC1FLD42N48Gs3ylxcT8nrh/ix9Ul1xqX8W
8nOArUWgOIFLbqfnaZej/wwRRQSPthkKNdR+8gGN3L70hbA1DzO1Nh/jJc8u
9Zln

`pragma protect end_protected
