// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
d8rzLkPQMR6ih5qkBoSdw5gtu0B6iMNYBuE7SKCibJI2YgqctsuPMULhh5Jc24wG
g37reZcwmzI28spkWVy7nnbK0zYqBoCoQq71cKw7MWoN47IpuUhMPM+bqT813O2V
f+hnci/9xmGH83h6ihERWyO8ZVrIT340YZXMAOMf5uJ1XBDkxS47Ag==
//pragma protect end_key_block
//pragma protect digest_block
MLRWCcueo4U5w7HjJYM099/suWs=
//pragma protect end_digest_block
//pragma protect data_block
KKEc6/Qvs4HrXTS+nvsEnCMfHgWFutNg5DR8REUc3XkufeEpeJimKBMpakoeUvPH
VW3HeYe3XZV1Dw4+z00TKFsqYz/jDvmQB9x36LS2k3bViLFFzB25QLOHH1kFEgIe
gUkp9lpHUbdpZulJzzXDM1tYvKpOBqS8slvuMFq4DFKWsP2zy9rVd09TIJhMzeTs
ptdNcKpkBdM0fkCxfYlUMG3PkTIknV19TQ2jSlfANRm6iQKXZWKEctIkoAudW96h
DQioQL0C/41Wx1z3YvgMDMDW9HkL1giOIEdSWFT6elzXztsYKW+v7fNBl2i7heJv
0AzXVwQk+bzMoaJxx219+2Goo+TUG3ZMIRPLU/h5nyyTW9fiH5xBBrrMxN0gboXB
4nBtgMRk3JioVyj0jz3gFclDwzT45Zc1IZxqrHV+hAFA0qiACsb/6oCsLHdFPfwM
NaPnUUQAsEBmv3H4ZoXPU0bW/+LDVUZKskL6L/195nN2eCqm8AEcF7hzFeespFIz
XkJGx8+8d2uhIaVKr+kvzh065ChA5goA48mFJF0Sf82o5c3eKZJify8qzhOfsrvz
UbUdsHZfyXF9hYa6p+uGzUhZz/k/c1v4m1dPJ3y6eW9Ozo3+jGKrrLMOu8VBKEDn
t//48mYHDB/cQSU8VXJF3+glsU28z8tVWXKyx68Cg1K/IjsslB5PYOCz4p748d9D
sS2XuJm4TGR8lqCjF2ucOnb+iDft1gZ90jkGKZHnIovfZWjx7VEvdnE+WqOpbpwe
jpS4+to9q7V3dop3RVkPz9nsozu5059ue7aPpQlrVBwSdmbPg4IbM183K+T2klF/
JFeOFju/DeC7PnTqlgJY9Dc5XdVgCXNQ/DhUHT9UxclQmEhGnykpL5NXbQGb7dS1
NB4nYnPtZ3UJ7hiIrY70NdMpEKDNlUl7Lf+dXRkwA2HSqBDu2MeMDi/g6aLw8xP5
9hRl/R7VLVj6qRWGSKOBEjb0+Y6y84wLIqr/+6atjz9wOODfn5b226pi0AUmw+nI
un5s/wpCxbArZYZ3Olk4LR6lZbukpr4IflqSvNcHMWMdQewXspYWxcNJwGAMeio/
sywpQ8pV1fSkSYeXmUHre7zy9jAK1jKEzgjD0OZxx1FH4yIzEu/SL8xjSBnliMZV
AXV2KFN3tSIxVI8Fi39axdhdZ09YGBF7iti0q3ODHlVU86ZDd4fEWg0rNrse0z7Z
x4nQ18ubk2fQGdeUP4iVeaZ0ypScBQ1MuADUwHnrclFypdtLCu5lIU9jZwPtwsml
zVzXXKVOtSDtdNeQrhT9erIPiDi3apA1zf/R4IpD+METxttm5ux2nl3pS91aFOrW
I+mFEZ8R2K//OxwQSoga+p08NgL+j40Dx9qXfw0dSBRY5Z+9BrYNKqVmMg5i7v59
Am1LfJGbcPeNDCfgK9HX3SRZ6TAhhsbp0n2eZ4PwIUqEJTfhobcn99exS/qqMj/z
tju0nUkVu9nJG5O91LO+gaAthLqizU3ZnIfUa5w5DiVcxD6pkXYIgxhAz4RRsiU6
FEw78Xo5FK4ZrL+CZKWeWrZfVGSanDx26nIEUt2CmIusVImtgjxf9ThmrnUP4E1L
FjVEVjM1R77mPEvTMDFYYyVuLrJM1LLnoAbC8Gts8Xw1JA++PTCoUrL3lNXuJPTE
oRC+XdlMd14tERf/xk9RP0hI2kdXeymh4I5aYXeV/midITp9TypuFxrLb2Yd7zpE
oGeJI9YfsBXOFor/qKF/ajjV6GP4oTDvOHuaRNknSx89pm15AvY7QI3AdQWAVk5a
T0gyxIiJvU+bPHTe4b0YcougNvMtxM4xM1n2MhGIYRKtZxekEwxfmbuWGMM8BtrA
W/HHqeYtPuTHuu8SWsLuzEw2HLipKhPAj3Yn7myqwVvr0tx6VcuOUIQ4k7Rt8zBj
pPDcVnAc4rCkdQvYsRmkVFMW9bh83GQN/Dtf8nSBKy4/qV67JEpWj9jlCU5ZXyYU
SUHZks+LaygXkYzWXv/0xEnYLtRx6n7Ii1VF1NGIEzHYhF8UNpezH88MElzDKjUP
N87PsJjF2o0Lh7jnJzubLWhmqUsqpw9QLS47qK1b1SjqS2tbMBT55pncD8mTNNig
NRda4v3CbO9MiVIdo/1pQXqPpAayEDXSBzDPpv+ibjKa9zL3Qb1COdb5YCVB28ra
9+CE4vYjnuaeBVQNir4PxsBDBzhRr5cNZa0APtVGDs8N5cMb/+tkAa73DXpeVPJp
TT3ZGlUfRA1wtvTYiuRzW+hpV0LUz0VZ0iG7WDqfVKCD6kATIniz2Mo9UORJ+C09
Lwc1VB7zZjftjfIwwuTCjV5j0YB8LC30aSzNdnUmzkDCbWIXlhcTymeFRt2asLTu
Nx/sprOzg5O3gptJ5+63EedTM4WmwGzFuqTMWymlbrks6lvfGzh26Vb3pVZtvBAC
G7ltSut96zmV/5Sp7yAUPtWCgUD1/5sKJos7UjzyJWa2tNynUC8TMLdGif26BLbV
tkOwCx+BIiv8UGMr8DyLNJJmfFAKijIPbKBLyMmPFPgpICozav4BkYquQTojV+AG
K9ykCDwOFENg99e5/7Niyc7wKDaEwny+RPtFm/VG67t0zoij/ifd5Nmyo5/C7i1k
lYaW7MN9DqX0tNJQhU4GMzPRfwcxrwxQQY1DCHbloM98q5YBCfEGGrALA17rsPGO
3xZ9furSWEbHGuMdn2juLMiy4oQmKuAXluyOqhSTjzPT0yVsT3k1yfu4UCkYhu/h
EgMqlBNqq9IWtwUf17KkPWpjpd9qJe8o9OweoeSOPJnAL3jI9cRwOliTtyqn+r2c
IV/wLpKdDzd5/XloNiZLzKAm+YO/sv7ZryUg0vp5RaD+WbQjdJ+4Wq8e+n6rrP4k
S7jfl32tIuwikwLAK03maH1KyGF3s4jTR5sVKxVlFeL95qSr6yiSvREgBUZOf20I
q2z913Y/it7nKZRtGL1gts3meojFhq4CT5f0TflMY1dupdfJvTzeFjB9Q3gmGUEn
AD6AWzOZPOP0rN7buVKf07gOv2C9AYo4PEIT2NteXf10EcEKVArQvaSM9BIolwAj
Aum1+whlF/vqvLILm+YWTpxbvVMTOid3iu02crbax6JdM5Mn3JXX0DhnrZCuo4fU
eDcmS1KZbPj1QDydHNxZqAFVYxmC32I0xxK2SZqThKCjJWMiJt9lhdt+rDVY9FA8
JCVsB+9eTSxoZKPbOpTFL/LJY1cNdfyzi+72+MgNeODBkPp2MKY11I2kUUdEO2rA
aTKV34cXNV0pAUncgI49O64jN+QFNP0bpX52UpNiqj46m6RZkyQTOHDiHc8SZFkS
Z52wz5h4AExGNFy3m266+I2e20lt1MlRkILfW/M5JYkVZX25cK+JjVZ+544YosWD
wqwJG4kNUX6W6yei6c40sa9LMj0qUDVjc6l1dLrPtPU/9roH/70YWQMmaT7JpCEY
8zK9SSnea7JGZ+Gvm/8TqPTPkk6uoqouy2d7hqqJirnrBKymmeqrj80J8UAA1ybV
WahQp16qGLgVb1RiTKWAKutiDHBA5Rh4Sxw+ISEhztDnqMY9XXH8B28B1B9DRNdz
HgOGXk5C/aw7tKzEBCBGZtcYY0Ff9zo5pcu0SMS/PRMBJY2a4XUBVSXrxzdyFeo5
MoIdkpHUdtcbQAb2N9v3jkSXSlxHUCCg67Gh5lzPfyMNOX4czm2/OgJV3R/ENWk+
i50SJQfpvl5WgOrjaCzBL6t4gtJ6sCEcKcxSa+TDUfaeHRAYSfZe4iJpqLriTtXo
9gvXd4Lb514zPf91fX85XGKxYQcQ8pBhH08coSjmKlWAJdJLnh2Hcvqk0EKM+AqM
AdikLzRMt+RBEUPP130/lA6wTA81rWT8GMBj9f2IIW7zU5w1QivZBK9gza0NQLgG
5FCyeMcQ+1T3dLrjY6LvG4Lhrq3AoelPUTsKZ9LVX8nxkF8tjlmVsTdppkzMAXRQ
2SIU7XLEBj3S9RuzZGp6fw9fgZgvnTAGG9L0sPjwigSGn/Rdsp7CzEZau0Mwm6m9
M1HhM51WSuP9B7oQjsCaaiUljJwfxP8kY6104QXHPxswt5JPR68+eyFBmMD8RS9c
PW1oaeOuvFtq3LfXqICUu4VQHEMnz4Ttlpbg5U7VrOLcOhvrnXnShk7Rc6wWWAtj
bskMMgNBMzYA543QSt1Gdfp381Q3OTXdwPWhifeZieBrx0tWEGkxRbVRtxyEq4p3
8wN7z73V6yMhI3bJKv/8qvu9aUzPBXut/KfBxgwzHRHGLyiyFHH1vawePQpcYlh3
4mQEjJtm3h/WU4HaYmX+tekOkwnHZ4HRAsvOANCIjhOAKhbx/C2rEr65xVOAZd2R
v6AfkAwqhtJnjyf4MolrPjSPglD7U1KItE/8DuTcTxlfezn7DWLPtoY2nsE4ySCt
hgpAFGVUY2AjcJC2fJAFKmnuKjI1z4beUOC7MJEZTw4QecqEKailek699TNfkw4P
wjRja8avcnar+vxeIfze8XvK0H6rVFjghP+8pfzHYObkX84yNlayo1fGnO1fNDDO
TxAK5O0u+7McO+QW1lPG5ai+83seXvhNtiALq4Cp8Jqm/10ZZQ8M/csAc2c0yIsD
MrYKv7weh4PD7R6GT9wXpBWFGaa59usYZhX0lWJEhpJrRZuObDP5GiGlCvqSZ3zp
wEyoNyWKb2pTxlgUO6e1lvIy+0wz57h/L0GsdXxpnUthFd7CcXb+KK9GI3zPnTdc
ZlYB2FHbztmejriL88YgNRU77Jiv5Yj9n/hTFs0Al0CFet63M0zOjM/Zah0qFQNO
7hN8y+VMDWXZcCAVFZinGOpKCgfSiB/lS/OwhOBlX6pFnjvYR5KcflwlVEIT/lh2
+E8SaguJtidiJixpLqeITrSottXMyDRj3Od+yuCkgeWdESHWq6ptliOeUb+xtjkB
63OqtytPHTOjiNITMzRXVkn+wQXd2FcCbyY6pWnAm4Wf6DKGXqk6uhyFKnZlpxWx
ZCFGVHbjEMndr6ug9sy1wmGC1z6r7dcNilg/GgqBivJX4oWO0NNzyS5ud6YP9FuS
XhX1jjfwOE/If9IoALiHuzDNjPrqFuJziYdrT+A7KQwh3c8zZKR+SjFzODI35YSV
IStHG5kHVL3WERVaMH6yOTWNv+JsoMgT38avQHEhgPV/vGG/FkvhLmuqTdTr35PZ
dcb3An20DOsS8uGRh/3OwKBfB1uzAYd7oLCw3yykn88PCfw7IJ+lJ/2LrKEO6M3a
FNQiyUJy0H4QrJ0iEgwsJhIOYW7X9xvP49mG5XBZ1Zo/hMsPZ0uDYj5GolP1xND7
93bYvuU0uMBGvRWjYPxfYbel4bR0kL4ieU1duUw8RKp8IlTJ91JSZwsL5WkCstOW
IVjGTNjsoZJ1iDmari3YMzXqoldeGwmk/9iy3FSMDg/kGnpn80Pb1y1HMrvMvKbR
0/9uHZeM1Ddx0NtY+eaKykilxm+hRYPAnp0Jngww4lp7e1doZvO6mdec8f2tJ4n8
UVNhOnt5Jy7o/H+Jul0I5oYMDoX/a0ssPBPeq9nyK6f40UPXT1lTsXuG8ayo1QKs
YBQV39mJ9qFK0MXTBHgbqBUgzBmMO0aQMHVVLkQKnZCaVNzyjQ+PJjrpOW9r/3kY
z5W6Nx/vR0HWjWeU8cNUvEC2YMDQcVO4kdV9WtgqlEYYXyPcDDFkEunExQfsJuwT
4Z8a38aRh6bmWi+z3UYLoMG5gOKveKN+qSZjBY5KMx3OjcC/O3m5Us1w8p464i4X
KaXKn9eLOMfIhQHoCGDwvH78m84YbOwCUL4J5r1VefZt+taoJJWz/VEqXyq5kkmz
EULWQEMpInBqMiuLOgkv5a/7Wan5IOjU2V0LvtKMYaIc6FxI19wyKzOseGD16PJ9
7dA+QarhzPInH6WjHLUcFMTiw0q39CfZkQ+1kh/uUeQcTvsWEV3Koj/LWuLKLU05
jhp5IKdehHejP4lcypCLti8VXMIi9tn40083fxBHhqMs6DCOLxfcWVB/jX9yeliR
iNW48vlF9pLGV2fi4GUgjCZ0UbDgYm2ON+QzFGA/6KWQ7+54ZJfqFcYtiQJKh1Z0
yLu1/jBFYQyrFLWR9EcLgwGMxr6D+TgWUpqKNPJ//b2K0fQZkFfxjgXT05swOeq4
3hApJGwnx0auCI6w8xDFKrTqL3JAEoo2TTjwztwlBOYnh71GNyDk/KcrSWSfhowZ
pND2iUJnGjrnoWTiFEFLq7IPO2uJ7qq3Y8+aeqJbSao5HROUtgjciiKrv+C5jx7Y
/UsZp5XAQLDJGWQKtprSO5ESPna+zjrEWCd00/na3RRkg7NooK6BlYkEJ+KN9XVF
xaLqwbScNiqiQbqt7PvNehKwVclqvJNg+ZCJaoQelp3oB8Uuk0Zj0pX3djSeN1ws
D/UBVSHDd4fowZknq18pB6blZFpI8cU4DEfbKAQJoRQ=
//pragma protect end_data_block
//pragma protect digest_block
eFDWiJ0vlKV3ydEswz2HM2M43UM=
//pragma protect end_digest_block
//pragma protect end_protected
