// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
0nP5iTydmcPXiD1HS38uyylWGr2772C66Tv7Irvmt7RmjfEV8M66sRJArD4N
Iyb/v/egXk9SQqdjxCj+kq7kta49nmepXpnjC6L3lXc8OjBZgtXwbCxTdfWs
F6XlISFgeVMqDM3OiRfqjxSmC/kouCueuvSZFrYruXHWeKzCmVX8TTbVfveO
2/m/9WxGdn3hCCGTEj4iu7ryERM/Mswy8CFi+zpDpXO6JNBJUnDvgSThCYTY
yMLgcl+g4FaFVvDl+3PvlVHouL86a4G9rtJmWKHN6FWXldPzzSbnVmW7zslR
th6QIbKuDOIkPOqILejqVaMhzfBPDsKIFC1F3Ein7g==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
fZZLQnGKCWP77uyXTz7jwLn5J+WV8plcw1ZlipZnjgHjtPTp5tLiAjkofpzy
G24GRphY3l7UZig0lVBiRrWWcc9eH6T49a8q7wpUH3SNcAPK7dwFkqd3g3u1
gNwXe8AHKP4Mmbv1FxhjbGaPT5EZ6xhIarRcGdHxRd9yDFsaPHagFmRxVcMG
Gc56/3Xs8ZBsJ+JH594diG49v7/jEZE+LZ4gZ2jpzewaOGBxxo+R/68I/KfE
OVZjKRNejrTJE9g3j2YNL6ER6J+R65zGViwiWXZnYOXCvIVY8lfhsr2EMwwS
gnk2bA5Angv/GC2bnDuFuhehhY8uXR5BLQD01gamKA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
dgII8GZQ1XiS8R7ykbRG/lT0ySouTwrdPaojhvKE3vmPQdgIpENp1up8rkwy
SKN9RVLqv4PkT60hJC+KUnmtKVI708qJ/A0Na7mqZv2OiF0xL0Ajs88ZMhp/
twaOcJ8TUdh1WnCTAGSQEWpPNRKU+kK5tkN48KAWlzKOjbxongX4Q0zukleF
5ZrVh0vdDnj9Qvkrg3gTBbs4/bfKlm/qeJ3d/asZr9XNnJ4BkjodlfyQ7uZP
8hvqQrZ+mzoluDWEhf9DKCRQatC6FbjeC3/TEi0LpAebsksLBQF4a4DkLgSd
Q3wEkyApsCe5laMVgqQR0AYuKJzxsYO/nHDB8MOYuQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
kdPNiDDt+LJqGoi1yvhE837qORCklQDnXJL/V1a8mQ0N4o1vhiRwXsj3xRSX
7+Hk4HotoIqs6GqYV8BS3Re8p6dJ1Zc+/54vEtPmj9Bo6pLlmS0CpLWQeP4u
Ju9hlbcPAJI/Gyaf1GOFWIKgdLIfYV0GFfS786wwQ3rPxPImjfo=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
nQRA9nR7/2gyFSzNliF9+Awc+cKubqXJ8v5U9Z817I05Srx+LjtonbkhCHo2
gRXUmWs/iXJRvamJFLhKMbYZ+Q+L1RfRoRKXPshjUnVkULc/zoQR4jCoA0rL
JCMriox7mo16fjabp5U9tDJ0BGm2Qm3ULbVWn65Tft4iNk8pl4N3A96mhqTT
xLWziBB5vLxf40vpZkg03562A+w8b1KhA1R3k2B8Iji2LU/AKfeGvNCOdZlf
K9OTea/p4pQL2XA3rhH7pMSy1hSVrjeDkQvf8Pn7/K1jbMa7mjETCHvvciTD
pwO3toYSl1y5PA2ChGXWdWsm3rIGVM8QDxXbqeXzrgtPlKTed9mIbsYw97cv
MzjMCx1Rf9DFI0tyMbQZmwlZYJoUO6o7iGHqXz0cI/XbCGUlP1MIHCu0sl2N
0tOKZOmV3AQCidC5kJNDagm8/kBBEYB93U0o+e1kn/yhqHRmc+S1nixBq0S2
iloyyNKQkRll4FVJ9+Fljjx7ipzXzh1E


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
kmeIH2cZwmWrGdXwSSK39zFhP7fsBopmjI1JVyEl4r2PH+5+7jhYMcu1AKrE
rSggtWvtaLrjJr2QSCls1Z7d3KJpLxRhD6pdu/RMgn2fn7TuECNkV57Dms+C
Z5PYZdXTH92FQFd33lJt5EOk/S+wRQj+Z160if3cLGSXoneoSRo=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
qrJ+5ldIUrJa38ZCt9ywpp1O+RDJRirRv1Tl8iEGlqCEEdf3pFkQdNd1FTr/
WpMJdIICJ1KYYWHnDWRCXUKh+SsRejly3sZlzgobNyN/tEv2Il1SVfsHsikG
2VustXe5gD+yk26hCVlC1SRJ/yvcF/glvhy5/U0Ofo8khSmbrkQ=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 65472)
`pragma protect data_block
gnuru/2ip7/maeVwFF8L4FqOlPcyUtEu4itGAZu7kFRZ+S9OQWKyE4GTqXM+
zB37opFVhEEx4Tc/gxQFT36OOPdcLN1bWYlYZlbd9HrJ2PDqrNEI0LwSYmp9
P8jCjEoGaANwa7WwF1OgE5xhfWSp+6d6KGE+b4e8JQoQ3KfVjZf260y3tUjs
qftxRF0D/ehtWpG/C5+gOX8O4I8vpheLZj54e5SZmJa+9koPazPbu2TuX14V
dLPODyqXyWh8giDXUq90Fo5qtDqUMW+z4yWDz6uiBAez2nxG5vMwW61rzs2K
L3tzHIGcSggzHci5koL6RvK9tDB2wH4V4B4kJO7eYSHcoP+KFxLElU5RppM7
VmbM9Ue/XY4eUGQGFUQ1HbKVXzi7PJmE256RezmnxLsty22DZWPD+jyS6x3j
LjpxpwO+1oOnTV/n9sMvA8Aj8lR4nSnWvVg74kNp0CLBvSkEpNKI5BGxUJJK
Q/1zs9Sp1mMgf7YwFBf1OHZvrCsqOwBIpZMJnStNhsz4LwrWPXy1SGBwy+53
NIBRlQN81zMZvxP9CvFCipV+rn3nlewlF10KTNP9fVzyyriByz+l9a/50uOr
aOchhdIItuERqV9i5bxBNGl73NJaXjhsGBhDkCV1ulmdD6L8lTr2GVC8JzbU
6beJ+CqVqMstyLiEDZHwkOzEWKvuk2cZPzH5fXsYz98J1e+2pnIcPEgu2hkj
YfTzMYmdZyfYGDt2bA+PeObaZm6tzbwAKUskjQV/aOiLcFHq2KGroluhQsfd
RDGdqwLBidROm+jgnB6NnxyqdmZQrZO9zK+M8wAsic2R0FXmD3c3QOr4Atea
pIB/aY5uEayBFUtknBTNhl8cioG85pKyXhhBapMyhDh7Qqvs5jvC6tp695ls
pN5sIxX6WKODHz8tdicgkJqdQ2tvcVuco9Id+T5gncp3IXe7Ps7CuvbfGTOZ
T2Et5P+NE4wPXW25x9Gctp8gSnn48CfqGSkd8sMYMpKflD6S+dSC99VlVAse
z+JkVTxlCniv6OXGEx7jj882m1YdcevMVt4mdSXLB2gd+HBcaZyMtCP4n+Do
cQnsH4smpNLKFcUnYJLA8h3dlclSyhcW9K1jLe2A4d3OwL6yn/r0vBp3CusM
gH40rNc1BWyuAufa3qIsyzeQ82SLmVE3f9ahPzI5omxJOhge9kR/ENgcfToO
D6QnQueIm3/09v2NNmW20IELBj+xHZIMp08A/j9nR1TV5MDf97Sd5Ri5OcIh
lYK168aWqFcIb6w7So6G8jsWLodsV1pBPks6AxvHSxaCamAlg3DNn2R29tP1
+QaBbjpK5Fgj1vmFz/EVvL2LjJK63FH+t0nGZNzevDp/0FRq6ozY/qMfQhOW
VJonT1I4lFgrJAmAZII7EB66T2R9WYsLqbnDXK0VyJoMeAu/nT3nViiB/KBY
HFWhP4OyprE0tr21RmlleIeo+amAEJjLZMOYT10VHCy2gLSX7bjgMGeY3x+c
+61h+4inYQjV36DdjQgfsO+AgD4raVwtFeLNfj5SKB77wlz24+/FXdJBD9W4
R2IMSYoyytgMVA4CSW0mhdX4QHJmmscfgI/ckW94Jo62uJw8XL2CKyPGet33
fmL8vc6Op5MwmCtg0U9AyroCwejkEjbmSoEH43+hrjmNAJTooB8byHwbNoIC
2jovnPVEdcD7tA68NB9UaEvyctqfg3WwcKue45c+q8LsTaEnLTDFePlZS1oQ
+ooVl1FsLu9BGZ35hOOFk1NQ2/WVKgl5QD4EtkrTUTREy0HF2+nQPv2nz8tH
BLFGYHuiOvy1YYa8cfS4gxuaiDLFv8zdceQGzRXcz3Jqh0qvAXgclQd5lzML
v+4MGaadrGRReC911VJ3tNlStk/zfkFGjU72sn0HSeNLb1GUS7if6pwSaSnd
fzSoDQFGy55QyizROwqujWbmfM4kioGH6OQtX8yHPWMdZ1UfvNY1Q+cuvM5a
Ddg7n6feUPy/X69plRVL5qeyXz/EtNI7IxQAkXsgzJXAq8PfTakkGTZlrCcf
NYVWi5QrDL8y87Sg0fmT2lD6LBucxRjF3CWSxD0BV7QvT/Yawqx1ffR0mEgi
+y2WelyEN/rqzEhFkz9CZTfKCk2TqJdTadvVfz2g7h3R1TdUc7K8Af+spT43
dMUFXM7fi6J5ndRWGcgJCgstQAlfMnJGOw7Jzo9JEA82my5M88K81vgM4hxy
HP5WmOJL+oFkIVhbIjS6PkWZ339oqYwCokxj/d87bMczr4kRWd82/S3OujjC
8R3qP6NP9a/mfdXHRSXh+X5MRu3FSPXDF7FgunSpAyPxXMIY/sayvR1+iGch
WHuo7D5dVoyIVR3J+tOv6Kauy9/tB48bIhKYRJiQQriyJl1qpJLb8u9zolnC
6PbYshZc/CRpcWWSI3iMzqX9F/rCxcyQP6WIfGT3Wo8Mwdh7OWUUhhHBv3LT
u0oCx3i+rCzI8mq692r1OwUgsgW1DgtfAkroCIz/NmDFSFBw5IUP/7nhPXXr
RtE28rL1WjOK5IXNQ73enJ2WGdDYpi6dCPn6RsMoKU5ldkAK2BRTOMxmNEny
R6oZPIZk7s/5xUvHZPpYy4ejMJtQWKoVtjehfUB+VEum4GDnfglm3xkJ6XpK
SznxBJCtuIMgV/Q/5vqvdC6oUpumkTHUntVSN690dplafUnPx7UfLiqTXRym
fxr7hJcE7QY5OeUx7O0OQzbl7cpSaSzMz526OS5v9XnxXTRmG4InfxLXGoIZ
OE0FyZB9JMnoUDDw7NohGdaD6g9DOC2gOyhWXk/mZBNnmIm1ENTbMatyXDd7
3klNA+VIKRtIhE7pfrE29G9yP5zyb+/4x0+hFEtJWXamVFNdgkedFpQwEO30
3jdPeBAqQcrB2bOz5n1CS+osdhhsygS4Lv4Jq95dg8p5P1CA0N06irh3ux4t
J5+aUceiDslGF8/DyR1P6C9Q5p7AnK4uDzgp2ntMhivGOV7JlmWM06XtNwtg
qptxeMRjWUVfVRP7SjavDVBeeT9pfI1U8lDbnneTCx9T85GWBSBaVnPbKPNc
a6OfH9RmFHGu039xKC9lSiHPl02Ej/4CESnh3CqnLgiEbH4b7r86pX1aUzTP
Xo6kZJPp8xguBJW7F6BMZF+VhwbTx9HzCEc9lOUZbLIJfvbJ6IbIjH+i6ZDf
5walCvbvH531ilCAH/Aktq1bB3egvwemtdZHp1x0TkHHpOW113XJFlSzwSse
TbhQihWzWEoMDe8Y+Upyk2DJ1xh4aoL5WWlmkpSOUqn7VhI0mUVFNAcT3Arm
YPwbsBMdEhNk+rp75Uq8spYU6wtVTCbPlcsL8pRW9XzQIwRJpTXBhuqPpR/h
9PYfnX4vz427+zlLDYG8g62z1g7KFJggmLbZHsCocLuIDHSi0OM0vSvvvDMw
/TTyhjPi1PtiL3IucXrHcxWcU9PtUoc8aNf3Y29fxT4CNmxBYqSrAJz5Udb5
JZXUpwsgmoier/oRtLwtukFDiIcMP7R7Xxm6WiKtbrBlBgpjtSwwHTZ2vG/F
MgMRYppVxY496Pq2J9q7iZqvKrMgelDXUUYm96LUNobFiKjaSfWdSAISuXqD
DaHNGFmDJUGMcHi078vC7VoCU06DAcRQFO0LBQImsMO0q3un/xtQWPSyUQX9
TONvwHxg886EH827342zIDTUH86GIXZaqZEtl38TOapp37Vo0bsH3TZTWLHO
7P5kIwU9c+zYP/DeQKlepcFzwytdwW/FDoEQqKMvYlYXxVc0RuOKby6C0p83
Ioid2KiXgNtgRB5m44TzwOfkvRLybdskjtcygU817mU5nasRAaZtrKQ2fklF
536n127Q7Khl2mAd17RuBQw/ua3AOlRiPL6c3rQQ6IgGa3xB53RsWIJL/jKy
LvXu84AQLoKpEF+L5ayAmdZ/Mc5vVT6BEhiBWtQTBLXRj+rCsQ21XpJg/Bw2
WxqucERnDJTdH2ioaPDa/0VNKOX+yIZ3L23YG1jCOAFy9VC9Shpg3Kw9cpmC
wYgJD/npK8VDKYF5ArAoOWvB1sYoXodOrCPcqhhC8/9gibcHHWg/HZWHulmb
6Nk6VjVKCL2I3v+NWShzkETAqJ8UtukmbZhjy+A/+t/Af9DBHc/noyVdD142
WceqcYWioOGzibGHiZ8zICpuIkvB+kG5p+07HWFXBWhLQhREww/E+Liix5ds
bMgJX5kPvo0dQQqcvBLCL3F9i3+yL4rVo2b4eh33WDsYEQAvQhAE3B9y6ENC
ph3OV4GIdeaI4sw1JdnBH2bU8veSIiaw6S5lf6Yld4H3mCt9ccHAYS08G4Xu
I67YDAad3B3F5TNbhqBy9CjHKWimHEbgyU81SXeozcVwNmYgb1or9xbxMo6A
m3K3x+4r94r1g4ZBtmyUaVJjR27V2AWF3Jzw4JeQjLV6xq1UlFR3nluUwzqY
zZkKjnzMLvns1GMgQmex0HZMi13AnaQTnAgI3QDPtSmmJ0+aG3NXLHAcPolS
IgW/rrT0nO9NWi1pcrWSffSm0UWD8mn4ttt0rfTmhWArgT+GwmeKrSBHQlVr
le10xTpvou3WGItSmtaXqo/3KA06ayWfDHAlTjStbO9t3CKSdSrrDBoYc2Pt
AK5H2WlWM7kIm2b39pAo07nrc67/uED60Cwx3aC8wyW4dPqTKODJLikGnL+3
U1TEANt9lqpxJ+AHd1UCA4LK5+CedwpvapZZpEgsuVO9frSHCN5YOG+qU7VL
kM3tzo/yMjspETZqQIgnVJ+LQppnoHY+O6RJ2NSW5NZgkd8fBVmnihmszYwe
ALWI2qObnnRMZ4/3ijGzIE7sjOrcc2rOpFCLVHVk51K/m1EG/WNK8ZAHaJlV
V+nozahuW+dwTPn5MZzbmchGtLCk2Ru1Qccud+oWZMGogGq+5UJZ8HuSlXSg
Tgc+eLWrP0Q4YnAqgnsw/QO7mbtZh8UafEHVpliRXIU5qr7tst/jqkOI4mIZ
GUUMvwPNn6U/BuQyVJER7FKfNjuH9804dhnflmyoneMg5dGtEEwKxYciCCst
eYS0ouV65br9YXz8A05S0vdKN+5cM7g873IJ7tQCjPTXLU2u7DlKeVAXdREv
fTH2drqYdpY/RbpIyMvva/lcAmik1E4NgQny10mhYpYTRJ74xOcriaEtkasu
/WwZWBtuew0sFbl7Zhmifq1gS/y554XgyaYvuOdm2prduYLBtBdogcrbaJHu
EVoh3lHz4jywRWC8NgghuZGrEzYSvqVVI+pHYhTdb8MoGM6kznlHUO+JwEid
8OB+aSoU5US8ecF62wKNdO5eh519uaCxGkIL0mvgRGKu2kBCGYkmtCzoHWpm
5V/d5Hn9tJCMJFWFRPT3IjqFziVY6PDCVV7qaNsITxPWkHlPFEcNA67XcwlZ
oQ5TLoa6b2F699YI/TVBNev7saolCgrp+GUTB7D2zB2yfOTIQgpf33hspgMn
ZEUbNFqeN9nhT9E/CzuhQ4dzLQMPyDAsX9NZtTXreSafv5DS2ioJhccd/Oan
iAvN31CiFn6JsOLi1XX/EG3tXIs0epVIz9o6Ix0Up1Kyoh6mdXWlHyCD/B9S
qjgP06l2ou5Iftqysi+IPGKDmxncZVrILsS1K8Y4ZStj2YSNDq7TUnq3Sdmo
Qyj7EQfB1nKGj30xoF+pI3zBrRmI5BuhXj3PPH3lXoJ3F2NGk4ppXqHJTi3o
Fo1bZGac809XPbEjp3jaxLQWxFs2uLg3K6/3AJW3oBMWnzQ0YZ8DG98AXG7l
TjRbPvlkPB2eRoB6FeA+qV3kAz7zNE1LnNKJPvhnkV++XG2zOO0oLBfTVo/R
1oYollqC5dB5RvcV717cbyaKZM1EWupLDN5a/nz8RSAuOeZlvMLd0BkUPSba
lGwKALtAQvdK3wUE3+WfZnVcChPNJId9afKHNNyHD386hLZiOEXISBd45VrT
gegU1PINPRn12RLZn8RqxTEEr8hPfQRkBAOQlzsweqOlrq9Qu/wespfSma3w
ggS7yKW90+CioNd6pUlPxPvrlFQ8LTGcbE+IitdEr0NO1oiNgF6xeT4vBUba
RjnU3aPRkxDdHD30E/ZiA0UgHXSjoQCh39Y7YgkxxL3pMxBDKuOBj/Zs2bGM
xp63UXUf/o7+dOCDsB6LkS88d3McBt54igV8UJG+EITha15/RyyH2lczMcos
+iYgLfgrHLZsAybl/Dmq0Il0kXgtq3poYn17RqCU+jVsq7X0KzNRUY5L6WXI
AEQIQrBB1D68wNeE6f3v6Reir9hfj/zb17nJLiOXmLHtp6krd82X9bYiVszV
ebmcNUGPn1RyJt4td0Iw0sj3uig06SsLrrvBZ3XT5Q5NLCd+aDJePMBEYg7I
p2XwMZPyn4cvhtR2YP4B5nH0cDlPR7cavjbqcXzTdsuCoCWOl4S7JwvKFSkm
+vHoLNe8FtNfsTqovgZuMJG7bZdm65Kplfzyt5JuxmKpSNe7+B2zEnDW14RW
c1Z/JcXXRlvZfDhJue68i7mtE3LdE20UHLJuJxNgnLKXkBbQqISUyPyo1Dgw
2AX8JphYYLSJhAdYlW4MASdeDFBSQkPgFqMmFh/+KSjGa6/YasPStBbhLwaN
hJiICEkFEn87HfC3cgHzZDMr47ChDITv3+ugwnX6aF7Sxy+fuhyBNxT3FjpZ
xw+UUCAlIClaqfPytljfYoPBGnx49xb5F5FmuJVOd6G34SqmQAgxuD6ZtlEa
ReODR9T06vP+LlTRUci4Q3pDyNCV5X9hCoSEqt2ydQKu3XKNEL1NDJZ81DaH
7uvD+GVf3z+YGg5g1/J+0FOSaioLNGTK/iW0PHbNduZAMJg9jSfqXQg93zh/
+oHzp38Ih8H9lvYrVGowa19KHnEUCTZfsx7ccoHRv3ORz3eymIBhzSDRRUP0
dUBaxBhKsNLqts290n5pIZl2VbC5XzNC3iuW7Fi0efE5lU+7YI3pNgdSDPvv
O5o3hQK83PeEE+eWAKT2GBZCwZkUhivbKe5YUgB7AHYvKSDYvkFRb+71L6sq
bumqStTlph4TG3s+Et96JFSRjG7bQ4YxD/YIMt8TVlM5Y5fpEuczoqeKGjEG
MzqytaWoaF4qC2k/WbXdwoJ6JsUfCTA62GzhADbSAqjbIee5+g3xiSqpjVK6
8PPcNRRYbYDZcRFGZAji7u5J6dJnhmQydlNjB7R9XQaE5KIpNc0YTKP2swb6
QCTJZFw0pkc3YYdDLoDw/3mdZTbI7m3nuWH0dfnVFZf/Kobtu4blHbPLi30A
53SGHWAJAzCY3RDtdvpkH6WwTR1qmxmOqMG/1on78e0GNhw87MIQoYbvq+P7
gbkvzxMKSO6C1j7axAIlgRxZuOHpEUV+DMAl9gEi3UKUFDDRctCchBlq8hO9
HvicwA+3UwhHaAO5slLGCwMONhI7PLGyorkffaOoYdB8HyRbYlUQ6sBdoP++
egg/9nPAdbehLDquCNLjuwQlgHArEe8G+PJqxin3Wi/ho+Vcm6eiIc8QEGxH
TyfgjWPeHyB12/eYPdV8lKmF6Ar1/DVjHsvcRqt73y9ReiCQOXRpIczg4JD1
NChWj3TuosRZ6EW+KWGW0VWbAXt7rS1RfHMSSS+wSYoa1TXW+Ei13dUjdDVh
MlDvSH4QL7S/lhT1z+nMIQG6R7qt/PsA87k/S981S3xtDltjiwWZI8wpqJyB
L0aq6Ol7pg1Iw1s3U9oW2MaycBF1/55pepNq7lwN+SWxpCzMu2pN2ESwyMFU
OlWDGZeowBk48yyFY0a1hfrxLcNR/V2nNVrf+FIH9MjIyg/qG+ghWOmy924R
0x1PE4A/1aIiflNOc47fdrdNDLhRX4K2d+2VFaJTHIN6a+BzwINgQjtzqimO
AOyspLXrRVT3xuA2MMaktpf5wNBf1E2BxVGukO1ETJPgeDIm7U3829jajbiA
S5TSjrpJULqbr5+1n2rgtvMNAvELen+PaKGSqhijh/OLYeYgQV/Lb2ktchPA
YCSYtUtvuzq+wFPuo3ExZxcnTU7tu6tqev1Lt0xvyy/AYLDOk9coxY6nTFb8
Hm3g+B660HR/awNCipcPzV4nY6/CjI2nru0ptOEiLatSyawbVO+843hwR6B0
kTSeYyPc2CAU89aplxbBibbB86NdxxdHKTPYQs13tzBUiLHTBt7XYPZDrG+I
dwCAQnkipBfinxCqNV/uua1T7kuKAf7fCmMdTDgmKzsJVeTlKeFY4hpaum1g
Hs6J3fnW+F7oKvLaXWAtMKaJ2S1qtnwQjl4v5Jh7KLHIAV9jezxjPx/gV8L8
RVcY4cIuZDUNcki3V9tY/cmm8na0N80UfrGejlSuS4a7++rEuJukGhfeAPNo
k2Ngo74t6w1SeWbEIzQOakc108K804H22z30NqLUpnQXocAYXGQDs5wOXKQm
G3EM7U5j/AeAc5lmVN4j66HDMKq/yCw/TMGOu2uuKlHR3Y3Ru+R1IRtWF9xD
yVdzO2mgPa8fqEpbBVJqZ4YjdJZE4UUDgXPGsp8RFC58jRU78foFNiQi80vj
brD6kn31la24ECjlYPI7TcEqZ8Z5YrQVN4MT/nRejEpmLoLT6r3UG3IwiH5K
hGsIGK1jkVOeibC9RLvaOER6OdMru3lvey9ytY/tULok4syk9jFRPihqMnZR
lViuOAO4ToJt4jdlbNDrXZ3cbAJ0c6wWxBVc/i9S3rzwn80Nicjp+RgkpXWN
hf409NtgtOGinpr5gI5FQeWF8zUk5PJ/Nt+PYgLgnVXIKdwEVkCpsw7BQoUR
RcYP3EgJjdVS5lMKxktDIq2GX5MpW1eP1do7fe6sFokk/A6fJkOsaBH//LPc
93iWSD5pfM2qKH6dDI0+r4r4tNcBFELp8Y62LUjKgct8PMHYM0vZ/5/q3UEl
7ylv8X1/weS5QxWAqKy6IFbu+BuvVMISqx+qs7dYCN/zI6Ryr01F0pfxLRyv
Wtzt3PoWILLzlNWndZq7arQPNW9Nzk9LbY35RP4arl6HNmfKBKJ2xmywWvb9
voTShc09NuPAeLHAJSW/vb2lSHsFm7evgg2QO0iaMW1CMq/dx9A9g6RLuSze
qpL00LXCvVotZ5uWDwmap5H4WbA8pdYRgSEhi7tPoGQpaCugOFss6nWC8o0a
dVRsGYyomIGo6bIMbN9z6zM1cavymbgDUHFCu8jJPyCBhmfodEsaW0RLBa87
n4dPmYyyK3KvbzkAcNRVl3118Dn7K2oG0bTazC0uqCwH3ibXlKBdj4g1dPAO
qGtDbG0Xvi2BUAS4tWVXEBe9t6gG3YBCohdNmiawrqk4OZeNHB6DGzdONKZP
Is6+Mlbfx19+fE2aG6Vrah6QgTWAH2WhLzLmBK/C0zZDwxurtZSO0XAlzHor
ge+/sEkvN7Ofg0kxnnd7FgQfNNgukaxXAB13y4loMB328pduNfiwQgYpFzkD
GWdUryJYPs2rT6jm5CFLYjkI+1ZCQ4DujemLbElQFT4k4xnKqqeiObs+brqQ
8r3fraPN2R/4r1zOaKsMZwa80AI4BXA1OEh+ltEnizPtKQOpIfS/ygJYBGGs
eWs4zKq9PHImYvPXXMIFsOhx7fL3xhqMKI7KAwE9j8D/vw4E73l+LIJctYP4
D5XJIjqbbl4UIRzF/EfecRSW9oMLdC7H6Ba9hN9jo7InFLLCAhoILwfEEUoj
Z1ZUxEpzuzF8+h59oJHOgWN5vquuRvvM9N61TQOMVRbUYzLLzfUssc8Yasrh
3vCDIHBLrB5vg2CobiB6QuvyROTWhbmr/juN7bZ2C0GqgIEhYRTTa3as+zIi
tCegHt869h18kyOm5onYuG6R07Q0jA0OdBn51fuFfDz/dLUf8NEQn525ZFy2
TbA5e4awf2I65McohBTuVwrflfaI3l5joAmPclVzr40QN8EnTJ14RhzjUnm8
01B3OyudCyYxQDJc8uBEv19xbBQseHuaNtd7kn5JEDaaPXRQYjEExwkMMaOz
UbdutvKa81WgIfENp8hcXzC4LadaQzBlZjQv8pMSdCXIpnFnxo0joiIVMEcU
dOjczOyxO7/LEkG5WqenRH1fk8oNZ/8Cx/i0fIni/LEAi8CUYFg+69fTxj2S
jSGiEFxMKAgUYO/VWulmAJrmUq6K1W2gTvxK6OwrnMJnfU3R67AWPo1BygbO
2VUzPBZW0PANSEcKW71tGou+iufpucgJaTiRFIvh6GFzpJA6vou5kN5kFc6Y
7KgUZLkqlRV8IKknKnEVj+tIPJOOekmep9eL+w6HxXYrI3uC/liCeX46lKYk
4wBF366fl5N25XgnRaVQHe0W5BTZVT3glPV4ftrwMCS4S77bz0DO/xE7Iyj5
0Zy3m/Asom4e+4Glr/bAYQi3dLBt836HaVyhPkIA18lKBvufCo4pG2gikD+K
QWzF4Jatpk8UphoBoQzHXOjNV5paGNqMN7hqls1M0+m1Q9PScfLuS6K49wlz
hvQbiEL+9rMabC+jpVQ9bBsfL186/hTdOjEGu7JGUdLtAP/6k24Whn+qAUDI
kwxgIDw7A9ccgc3PuvW04wX34/rf/oVdCqYnGIRR9OJnjLmxMOZ8BzjcgdpP
7kLovnFSclXMU8lIrvdxdWBbrT2DvH7w2+jYmD/yETxdx0ZBGVmFrEPwJl2z
Blv436QllT2o+rVj1u3ExWld0VHJ1/xsKEdrpbTdJshS4ywTzg64Rq4fFPrd
YuyIK45/oiz0iHlFERQ7ykGKEoZ4LFEfZIk3uoNuN5wEHXoJ8fDSRsVAQGYv
1K9o027lNakxnxi/+jkgwno/fucFYzZ9gc4g2g+mrW5HLko0aV4YVcDqVNO3
dxn7WvmrxrQvQsHjLZhpZKIKXs98l6B6Ec56GxykSrVwmOXL7I7lOZMi1Fxq
9VOtbSBw8G/74JQnqL0M4QQizHa12CJ8HWNFUzyUvxMr2XstG2Ejw1uKfUQq
SILD8XVEto/2tgTFVidZThJTVvquTNkIem3wZyGoxjufwmcJToVbm+KRsCx0
nH4RXYO8bcU0rkG5p1nRd/WUhJBdV1v+4y+k2X3NWEiDETe+IIasSL6fB6EX
8K3/pjwvjY6d9wNqn1rh8oa0BlVyF5jKb3JdOODLFBQZqbY0meOsDjMnVb89
GkN2IuouXh1h29tdm4qgM0bIx2tb3R8bCyDuauUXR3HYYp9kyo0paiGBrG1i
CuydmBwpy5UOi/aJYGNNSM1vPtyFs6G4PLufItLwPCf2rc6BaruXh9U8gcn2
PDTkFYl2/mjhBAxTUzWRx8PVJY9yT0ysYi5Id9hGFbYQy5h/HS6ZZkCtAS/f
7/6TiXcEAVBaPVkiG4w97Ll0leWfHPzafZAkk7Fzh3f+PRPrevufscNF5p/m
IO3t7qtlZ/nSDT+IdWwLPRzPsj2WdPPLxnsx/cCDd0ICwm3vMdTMJ7fRzCJt
7GeLKyAEH7+Cc2meC0T4NZvSL5nAOIrJJsDH8OluR9nJm417TQFdhOBHp0Mn
nG2Yn/eUwfYfwsepHh+QGOznYAfad+pcobfqw2s7fgcFxCMg6IrA15U5l+c/
/00M7IEos+5kAkgFve4meMb7cP0TfTeg8Po2aAvdVkNI8GIW80rpwNApIDPg
xLgbXyykJttywkDl6P7tFS2KuNFPtlV3YSqYkwNf7KchfjAWtnrqxqXGDVxf
K1Zx7JFEmi+rzro1jbX+1qhiZy95WIfPTbd/J2h8GGqyP6rjkRb04fW7pH3H
iXdL1U1aJfB+uyldBA0ytdtfkGjlH0bPV37f2C803Ltf0/5+92QFIXoTgJaN
ZqBH466ug8Q8gLKyCdMwjkh6mftVewJ+fB4Lm9m/CFtOyILhdhSGbk6vxn3/
4EwzUFBUD8SIm5oU/ICeWVywnM0MWbTbju47ZNk0kOwTw4ffcRPI1nX5uCAs
qispKaCNC51LhWxEmkxvaUfSoS1iFqW6qTTb0coHUeh5GkPE5WV7KqyqCI3t
+yI5Xk+8LldTs56Nm8pM7451pCzXEunwrN9rNQGwnNmfe4Iu0bYtlVcDEeG4
fMmQWn7g6+yZ3X/crLdQfslq4fhhQ5H4RldaAEZUnjsZ0B+BntSBjp6tfnfn
XjHXzxK5Bw/XL9Go4A+xPtHR9dUnHFEAtF0IhowBdvseAiFL0Zv4XkTVVLGu
hriFDF1C5op/NMvk8X+/70QpyOyEbTfGVqrFFu2JKeta7i1TlJs1Hpfpm+XC
0AN6YaBUXegRYnJJw0u5nHvptCLpzL7VKj9qz/sFoOWtzyBvkQL6oYyonHrM
VGi+ewdMXTxVnGHsCAUWRoQuPN8shenIlyRcf4RkaOv7Comcez1vsS8JUH/V
4IKn3uWoGCMFFaQUGCkf2M5AvNbaS3AWI7G27bc+zUP3xQ7l06ZRaofBYy4g
M0qizmF+NVnsXFno2N7ntc0bEQ/lJvWQdKfTLzrjiGXPU1SNs+fzAROLYoFp
4HHFLEDH3jUZCdiquUUM3JUTkWsVgsT8xOejs82Ia0st+6ayU31k+xRdGb+W
nuw3JQ8WldpeuSD5NOV6cweepozlk2dy+E85QRi6CJrHrdvEy0VixvW1QgUc
3nQ7WNNHtwP5nkzHL+7wYb+MN9Oe82pT3Dh169oucJ8h+S/slRjXBGr8WrRZ
Pfd2E4D+DGSXW1FE8FRl7wEHGl4mBjEgsrHaOj5QZkm6uLXrh3+G2Ib7Ndfv
aWm2Emn61sAFjs+gK576EhlKTz+b7BHAoqyfjoBHX6Pn1E0grnnrHIU2KL17
1EskCnjgGpQvhiW2Vhhesp3sKf+p689yiEH75Ke/LEOmr6O+i7p5mrnZAjRO
moKil3iszF6xfP4lPbhVE5ORZUT2qsfzsWhfYx7Whe3peo+fVrX9ISdTHxZX
bprgAo1MTASMea1VTE8rzHJK1HnXVdlqtu1Bpk89/qGmcHxKzzx93XFuhiJd
/nrKGslCCe4efkT96D+L3FTaUDtuoBBpPIGA0n1fYMnfk7hAeGZ5bsIFdldE
X6XPSnl8Cz7viKce/zyONdpj3fciNvyTXbWkAxhfHViFstca7Hy7Ssk2qpeD
w9BaZCtumc9F/4KZyWejfFURpMQa2g1phTOmQBA69AzLSHHBhKKujvhESsxU
dAO5ngbNqIsePm3rZEdKjN88a8zLWivQ48tcMyhw04IvG6dQZZEPlRmNH2CA
2dwjgyYxnfIbBxBYsX4j2eAjVd3yRxw8u/F4zxnsVZdhbCEJg4JnWL8zC5Qq
sD3wadBdkewnZTTJ5XA7oNokUk+obwwoKM6/C24Wcnq3FimHfFux0EDhGGgl
4GH/oFn7P1miNJhui2fVrMKEzvuwdzFooQWO07JHRH63aawDdGvKwcgbgXbf
2maQOY6Tx8u4zHbjQm8JjhTKSiE0fSu51Cd9s2rRhqQnlktyIt+V/9c/YUhV
TPcKE7IAkE9P/kPEXGlMCV+p2drW3UUTNl228SzTrnwELjgbHHUUPE5kuDzF
0D+f0ipsz2nTVLsWI9iaH36amJwp92bvlzzvysdDB8IGssAlgi7WoqZX4FUz
Hbykk6+MlkU93iIjxGIk7pgm7+Ju/PRoF0jBucIXEwUOI/dw9ufsdKBMw7tW
YoMdDv3aFUi6RUnfcMXOJX+triLGkxPcNP2QS9sQ8sotKOg9tqvdUurb02Mq
SLo+hhNYncOxgn792VhB2/8HEsb10PQOOkSIzDr0jicLfhIFx7MlV+SKtDwc
RVGaCqFVczu6c3aCX25rNcdmy7PQz+eKUBfmx3E0i5eTpkCC0cIVmUjvL23L
J/6sFJ+Cw2YvEkoltn3MyGi5xXMetWxn7usqZj468cnlVn5D0xuuZlbvJdaD
SBX/3la4y6/4VPI+qnAYDDkCGxiCMbjrHZVCCbzhQsT1To6LYn67pEAnT1V0
mPLSkDvaYlbRcvf4hMJUOeTPMamiGW2sceBLfNlKHGRgw66/mlEYyaZA1/QD
/LJfgcBEQovQnYnr46qIlNiZ7Zp3lUHGjNUhecYUYYUYgOtcWfGnDV3vHSCF
Nt/+Gw3YrnVtAqxK+6347mGi2uPMA5BAZD999shC5xl+DYNhi2vpbeB+EqtZ
UcOvD7SmmjvkYrp2n46hRXLrEoN7c8gT00AHTXB9LG2Wvb4PvLhGVB6BZDjR
bGTEU3JlnBuIA+uyN5kcsRd72VvnA3zyn3yprKXfo2WW7/tQq114l4RL7yRa
bcCh2tuu9yno6byIo8MR+Ci5gpNI20MYu9CeWgAUzXbjH9bJJW+Yw7OYFpKw
HPSzymFLNatIzY/TODA0YgpxGW0GFbCUDnqJHv3qNLsijbe48CiESiYvq5WW
Da894ev2JbuhE2If6hRsVuF5RIhtLtJB406gtmxrqTkHyGtuQbx47Fdo2Jch
S1D5jLuCBhv0OUiDHR5VpiprnMKp3Cq0eMitaCdggZ4/iXeMLoEnM8fpBhwd
GI/aU3SKogX4VPH7IWROd3yKSQHGXlJqqEy8zaB0iUunyaRVpd8UbQXsuSz9
0OTtdzvIgDSoBJZi7Qur0S8Nmp39tSBCPgAYmyEU6OUX4SFhTJkGnaqRXTAV
A8m3vjThSXiJstxUFVbdSsxQehlvGHAcYW0Xu/jFxxRain0m6yuvgxt0hPpP
Gm7sxnKo64g68b7mWS5PlEN6rguIGl0qbvYTYbqehd0AIZOEun6PJJ8fCkrc
U/YdqlJiz0LqAopQri458DqSXAWObBzHf3ARJrjBUaODMf2gSFqFgPAlJzTm
dhm1UfBZNtfUuxQsBnXp46I309HFVwUTf6UwHxjm3SPWgZL32w0Hl0gVV0Ck
WQgdi8wrhs38B0kgeQJAllpenXR3DuTh2AxiF/n/RjjU7KaLQ3V3NLR5nizA
4SORv6aHpOq3pUxION3bB4sHwjQ1oKq0NXs1Q9CXsrTWZcPGTy/H9d0sCoOY
6Ak8s+XBYtshYjalWMRo91R3lKPBni7bVNAxZjUSKUVdGxeczMdmIM6s89yY
s6qOVxjY7hq+yq8ltHMvIY3/hdzTZCKH9l5p+9UelgUA2mxd/qjn7AV4Swau
RO5be3+44UIZLmIWnkUr8Rm/GECwTDiCK7y/2CPHi1jA5VqRPlIt9W4nNX7C
WYT6xKpjOYnWnl1As/tFJ1yqYEt4VhUmY1CM+EoP35gEFXzf1PbwWlnS2cqw
iD8avV2RVQezeowV/p7Kv5lbJByCtvZzQmGFiJKD41b2Y37lQybVl38huLfT
+hiG2hsnWIXp3QryjKOVO6kEFKVbNBQ0SfwhAgQJcMHZIoKr5zsWKx443dYp
Jk8PjSGgTamlNVLVWSwSU3JsHlgLn26gKREBDFPQiNvM2dyXT8tjI8WKSNt5
eCuESO5ZtsZ9vF1lGTeuqVhP7PWUmbIbowspxLeMnFtxnsqdeXxN5yvbElLl
BLmLriEw7TCP6Wfjg/0tT+DhBjrPrWhPRGCdBDXqLezNNdiVVsw6i/ejJH6T
CxAkyOq6yBSRDv4REwl5+2hZ+/z90lLsm8T5yiwusFGG0asRNzxwf087G+Le
sxs1xLPhukUwiQP9tgKhnDbRYLXGtAdEYQ3/5pYnHoGtRjxX0X8TAIWTEDXI
17OCGOVKL7rdk7di2bP9IZ+csCxAHLa++Jg0gzWDq9vyWx++EqPff1vvNHs8
Ew1we5MlWF8+ZIXq0ZbDllwS89xYTMTLRDTYRV8FgwAu8GLvgbcgAJhe9ePN
mSDyEr3dz6rvTXHUyxeHjHK3JlfXPxCZoVsPN4Hu4ys5i8WfvYvgQIeiXTUj
PAv+igUI8a1KY0e87qHmsV5AXCnArByXCCU48ikDaRokA6LGXs7fHwsvl6ly
7oLZcZ5hW5+IrRTyMThD0l9uzPqXPXxA2rpZQDSdSbO8yBI9e65x76NAGnVA
ZJtqfgH8And+6wod8/2Ott2CtKSFbK8bvOCx8nMA+ZqtwQSnGSFhZCysunNw
3mkEmLa+DB7DkMFoYgu7BCogQVP5EZQ24ooIHR9rPL/t7/1zXxtPgGKMD9Tv
k/DexQgNHt8aU1wTvzjIRiQYsKqC1xqgkqVUcyej9pmUBh3cD6lgs6SGbwK/
J6ZdbPNoeih390tf0c+PicSlX1yMDAg/D1XphVIRUc9ALwkb6rxQjzOCwK/z
nGfuZrXHOJY36Sgz1eF31gkYYaUE6ZTae3wzVbcZ0zOotr44ajf3R/jNy7Lr
4Qc5cV8jgcaRocwkDREzDLyBGZZaozJ2WvFpw8ljQ4vQxtg9+NzpVh4CVKvE
NAO7sCO+9rFfWswBjgHm7NSms4D4IFANkHds4hrSbevpHhlrcOe+eMnrH6NJ
w4u2G/Rv4uxGOd7eXKpZN45HFYWo8PeNcrzMsR9x/tjNUTDvPWGLmSaevdAz
mK2MnuxqTyWBOygxRoUEh7PV9kYe/prjd4LYDbi/A3cZSMAIWKMnR1saax4n
C9P14C13nVR/SKL9kGi7p+4jtemlh3TAMUDAIny27I/gEEqnfvsWr42I2SRM
7A77QW98kCUZCdZdF4OpbjZUgoPM5FiawlQCnGmHaZkhiBIN83thW1vSJT1D
0gM4lb/DYANxPRXpJo5G8TgmS7rkueG6lx51WJJcl/2LHvjCdbeXiqPGdUY6
05FErPltN0tlrvAoV39IjH13eziGjMM7A+x9eY2+Ea8fEalvHs1lla3Tg05d
pTOeqkx5+xm5U73gvlM088qSqw2Ebez2ec4Fv6cABHSbcJxvcVC01ysHnZrL
7i2tHiS92CC/q+VZSxeCCljAdiOTz2VAVKdc6Aue7WrBtrMw4Uq6eE42sQQM
n1dN/yjjKpkAfgW9RNEjMlGh/2SrH+Jx/qcyYZt2yJuo/bSDA90a3QEEd835
IlrA3Zep3JJk6N3tXqdk6fcN067lsAM9d3dOumFprxgTC4k0ifFwL56JDknA
dUfNeG9MgZRbs3JMiuqgaTPeMVYrGWQ/9CFKAGs4wic2PfqMzk0+1WR+uiws
4TPEsZP+psn907AQBN2Z7B+MRQTfQyRSLQKLgfeo/vbdUq9QhyaA6P2VePVV
5NIKt5aBu1SofZ2i8S0iMrCtGElwJaT5IVh1imWCowW0MXmGJ/FvgizteY2n
/U33hcRtGv4f/ANi35TtFy2AUKC/eVokHlzTQ5DrQ1PaAZQF3IWTE8Fj+Cfs
KjpgpI/SQYh0SMcPg1VMu0c5LHRaKVq6j1K7xtS2AvTpvVsLaEBO6cHOn+50
inq0EQ7h+COLpIgLail/UiEQVOxdX8OlkiLOtcl5lkYewqmgHbU7+X+nqsnw
cnDEsjM/FtFDYzS2NeHUc73k5VINq2z9WWJ0X7B2xTvhqGNqaSJkm8lCr4+K
Qd1GtZvRAaxk/izqNa/MEJ8CwsAdkxQOjG2YL/ZA5MLEpfzwhraflIy4kNBF
e6uJG2nrSzdUpRQMeVGs4RBdmSlcr5RGf9kfInGw5zMScqHLrjsxpcJEYZUJ
Ccl85rWJnxPbFJGMhzX6UEvnsK8/DttIFTp91pkb8gPFw+TXlQoNZHCpxctR
MapX/bR5dBHDpH6PWRIDQwOLUwjYTp/lKlepcal8ZxOIlKkJ4lTg4hR+JMsy
A6WeLi09+9e59SGMYNj4iD9UUN8ToutkL84vQm1A6z9zO62Ksi14Fx1fT/7r
WSz3IC0kqJ0ydBtd9xMpJyVQ2qx/ZfX2o3IW4vCeQAOt4NNGyI3n22qwL3SS
gbenqzsL1jE1H+qV2m4M8m40QfWCgaa/C7PezsRr2XSI18TuSTVTEm7qSCVo
VysHSkj6aBfJYXZsxtmHwgnR8rbAQbVQ6HppdvFm2seE8c8iTHzRiKTP7QdH
NXo9yHCyyxmEzy4y5fQnCptr2IaSWtFjelQdkXzNnfdcINNNgpPceGkSkbae
dvf4rok5X8s0iZF1qt0dywfkZEULmKXxpDCNNju7SFBf8RpNSuPohngLETeI
eNehddQPcrNOSzgaztJbPu6doyHld/EuBmfmC2ovgTi14TE/wiLxnbKmKy0g
4+l5mElYE/bk+JxgiTOz+ZhvdYeZrRePHPLjORVmf4MbPFwDaVpZbiJsXXQy
k5I5fd8s4qPAwgWFtVQ3zfFVf265XYXtcjoj9hnNuqlm7CwsTYoyl8uJgwS0
KoL0dcQjfpPsN6OSSjlNcnTI1RxacOs/8wyKu6aA04flQcc47E22ceDVkAR6
w6TEYk+1GgVrsM+ZhOTwJ7nscZXNup9fc+0PrnndUxHEhbfO9siWdOhW2Toz
1A0+Nk3OFsBvr6uMHaW6x3/WKWkkA4/rtl68Luqt+RZu2vlgNMYwSqUMFovv
LWx+Xb2iVPTEkdxz6toOHjGNn4qc03/ebwwM7bIlBIbjAX1kcvykNkdVHbKD
gyhaLHZgPE6vfcfAbJEeHsJEMAXlG/d6psJu+7vk53tHWUOmNAdLaEtLEL0w
XQXO7jN0gosn+/08lSnR8gIDOy1qAJBMNIDb3hKFCFIfpBSgDxdm8xq2VGOL
1K7X0YoKmnsKbOvTY0VvTnSioWi6ORDhBQCbhOYd0M9oOFAbbzOzdBK8mbav
Nv4LTNAAcEW7JrpRG56oxCoxqw0Y0XV3JTat4md7hq9QVhUJgEk32cBXeM3A
RB/y8ZUl7cJ2qQCr2Zmq6UEEPvDQEMSFHQZ0BNmXbj6+3/95hj0gC/++hBro
ps1WGn8nySB0NppKcPwJZpjVbcw0QvAvSFZDBv9YbQu0Rr0hG2aixnhMojLi
f+no72H1KCy/NQZKNnQntnS0mM/N7DO8JUzrx3B4USoHkNPPd1/pJmKksphV
1QiLQhxDo2DiCrkSLpljAfRhS0PCANC1t1clltGvBoGd+3BCvBPCahL10N+f
Jn8QyIfBR3fylxuJhiMo9txHMoBxRAMIRPyiSkcg18fdcXlXE4BJ0C6NvxZC
zlbT1Asf6MG1ocRXeyfS6IixWPM+2h78bTiMakdfgAoO5xbRc4DSiq7BMLNJ
XA2yRjTSc7ZkuKei5Jr2702LsPhH3wViz1RTf6oMVhgUo4x4L5o4Gkmt50Ej
Cpdcsuq4R1SwBAWf9YMv9gOHCBSTmKbiAScEeSDrI1pmTFFH0fQxUlYW4Q+S
1U3O4J4Sg6U6A4TPfYgvdwdzPYuXuO8D3SwCWpt4YG8bUdgnZMSIl12gj5oc
4W4zOPOuxP9+BY0zTr0UrhRSmK7ZtIxQS2ziiaMCp/lI+7LLeeVteagoAlp4
Zu3vzEKJXv5D7C7G3sj6HCVVXkYzl9hbbTTAJlqZi9l+Kjzb+P607sSqWtyb
cRA4KwVmbdcM/J4BpFErf2jbmLct+jz56a88YZXqIIhDR0snzY3+lkGZaxs0
QGpCIzXLKErga3373tsckxvUmN0J8v/aab/yurKIcvo7k+hAVXCk0TKk3Bf+
GCCgp4yYY99JRYoAV/U0Dn1OtEo1oyvyFX9EUhh6zZAN7kBNctLgRT7r7W65
Oc7oal6Lcufk28Hu3hi9POhka41xInGdJC51u+oyNIAgeHdPMnsdQscPUvyZ
WeRbcctuSqY+wfQQGqsWGeOee4LEB2G9Xs9H5Vi7Tqcgse8m+6znF8Qi6b2p
Wq94dVXldp08X8AbrxVNDBs2vCT4jDzrhYsN/psIb5cfTmyh35WCMlvmyh7O
0y7qJ45b62YC8BHkoFXeDOvP6dXsiGRF+47Zx2djC5+JhtVQw3AHgb+827j6
ALU32xFebsK1wk/9oeTt8wTyLZ6eENPdKI2ql7JIIJ++puGBXhqsBnuy5Yhn
1Hc7i+hkws1l21aejpm+aw9Eu9+o9lZOcOX0/um8Qu8IKNO4xhgfCbRLvki8
Vlb8VtBXlDm/hC+hZxg1gWgjb+FXQo5npLqktLg7oUkGlq8fxyoY2DBDXHju
XnJs8W7/Mf1EUoVRKivvOUZGHUz7g8FvdTCf4wCQvRx/uldW+CZBKcfUj5+6
v4OLpLIN1ErRNFiKDLtk2hkuXIfoEJl1xe4fzf/UB7IUKWh5G+QO2PcksleH
95oZMWVt/c1fXa9TkgyZ0L26SAUBPGpeH/RuQRnm6YYC2VDTYn/knUQjJsy2
zhv4veoF0lH20pAarq9axW1rx+xEY1eZq5dCTNhC0hrcr8RKmcnZhhi+rPN6
Mg4Qi8HHLoE+0tmF1rEML/CWe9+Jqi7rrqOB95UmkEeF6BU7Ltz6t13z/dXM
wxT2ElPB2lXgvHjmorlEGuIz2FP/MyRRl1poj4lX54ELbUc0u+9G/6pqPBuN
B9DLp6x/cbu/xTDz6nhRYBqVmRXTNNRjdo9iUmDA460EhfcN3dhtgpPrBOgH
xPIlnJU8kcfh1AtgEsmVdrDObUFxGVkOFa0oMIv7WkA2diMCTyxHLaybs//F
gSKmENKf/9sD+pjyFb/DN9xcqJE+QyAHs11IvHE4pwUNdfZHx4LjeVNs+6Be
+Y73H5ZSXGqGxQK8A+I2X1exSaurebKPp0GmqIWr3wdgWXhPVUtJ4jJ6fE79
pm9i5IzJx1RbWkO9FOnH2iSka8/7LSPPxAeyA0Tw5zsxvmxnY0VCaLsZAFDT
6nuTHKhZj4nta0mKKoMm9e7esp6uwm+eH8oFYDUd3whsnHgz41Df09mrlc9v
7pa0uy1YXQ2vcghExMUQHpEo28teUt8EMC/30A0jxFjGAyoH+TsPY4KVmjLQ
qcwQlTidrq0aPgQ07Jj6uS7JEXxN9WIKLRE3KGxqdR3orSsYjlqs17AMt7Bs
4wO/TJiXxvrPkfLjH9Jwz8ibbWY/K39N383sYkX7LyDlJVmTV1JFzyfffzLR
HOo8kmugjjry9eTRDhqu3XUA/2yGhHeIsb2jidc7197MB2N22FZA+FxuGiTb
4WhJ/6+bd8NfEV8cY2OMqEvHDiKdV3LG0y9PdisnT0rbAf6AsR+4M+tIy6Dv
L1Bh8w9fZW6AQLWlFRSuDFuPmROIhEHNhgVnphNXoj2Q6dZQiVm+EktU+09N
WaJ1KqJbJJwWiitGysk4gSJ3aHHbUmOfQFLrBYrKbYEjd1jU3iz8RtEDkStH
1qlhMasJIw0ww/JJ0KtR2ccJhPKBwupNucIquAQoQDuYI4KZW91o0wmbFsKW
fMysDvjWsz7rxmd7QQCYa2fTcS05G0hxGmOfcLeldDNhZmPxJp80jppY3PBU
GwRgnwZz315bkpffoM7asyJaW9+FyOKxaYI8YP6fBtv0xUwgps8/Sfa5y9y0
woT7kAShEAlOZTptY3uBgNOSxuOV/eBEZKzaaDkrGwinRZZU3fjq7QhgiGL4
xcBgOE5WwGp0eSGvF38eCS90m+x/+dhj9LWUtXCizuhrn8xlVh0355KOTo/Z
ECA0x/PyICzg7+yCwGMXs/afL5itL29OvFlZ00M5ESpjWamIXknvSqXonnXC
xGSm+Ui2CdTjMdGN4tQbPrO5MWBBpXP9f2mevpJSlsmjzpLwhg/QDFUIxlxO
Db5pTbj/m7rqlA19fgDPqef8c0wmcALh3Pdi9Qi4kEnr2pX1vTScVLFb9WHK
cZ58/42G8Hbo/QZHovP84EoSCmi+tPbr2pxiB+yvqLSr31BZJh9mXzXLEzWf
6HmHAZUH2/UsX2opR1atAwnZyF2uD9Y+UZXIwtML1lpMcG38syv4dqfrM0cA
AfjogTYRrgl9tp//b55Jtv/AGBxEK7WyPdikwhSUddM+vHJHJFfGtBEh8g85
nRuGpEt0xWt/nlSbu4X+AvQAAjOYxjH4CSCLRwVhVEQwSHB7wjIKmn6/iaxs
8KTLydstqkCdIyJ44/FFLNFYkUnVaERt/wp7fpwSfZVEaZpXkLuSVnBZpBMa
b9vOPyoF9OyCVyzmXryOJNlmAdkvcHAzEefgsHOL52iCBpdwPZAIThDS5Os8
VNZlfqCFVB3iGV88TeDP4llzYBuNLC9PtGUJbTF88kNE7PSXlRULDF4/j6rB
Wakq4dq312CmHQ0nsz8y/xEzn0PI+zqPobdf8Fi5LEsoibdv0shmPaCXduxL
HcTxG0gVfSb8M6jGdbPiZ0FTB89WehpyrTOyiDI/NmdT6HKX60ddNHqcoeg9
xnWa90b6UMlRWW8vHc+NHTruxQ0YfnXDWQU/39nyqEMv+YRfpDUNt18XKu7g
XZwZBKGVoFKInXri3hXKI7dCjVn5gmOsxQy7f1t1mPGMMq0PcURU31GG6Wk1
UmpzmRLnn/TO/Op9WY8fPawEUPeM9Sn8UCBRK7dvC3zoBHNQl6r3V39wNESj
nK01Lq1b/D/XOPmuktWWNIxcmQW5lOXKko4I4yznbStRZxXX/NyRBtHu6/Pp
7DQD7BSeulT4o05eQ5PkODlNF4HgS9qJzA43mEAJT3AfKqP7Z3PS4HMk0QrY
yu6Vl+m4mCTxdAeQE8wX2bzIktXWJlC4Im+eognuTwrGl7t8Dlp2f+f31XRl
urBq8k+YROjD/MoRhmm9QUihgXX8dx8T04CAJIf5qaF9IAVQHxRP+H/hXeOk
sI3vNlKn7hqYJeRFWuNyJZbRP3GX/Kg5M7lnriujRyDyBHWHa7l1OZkvHHdi
+OmHteMPTPXSpHeQDLDFI6k74QrhrLbteOMPq4/d/c+pvlbWG3vMYNjdGlAH
wMvYBuZfaMvbeY11pbVU+koiTD/v2acpyRs3ocQMUFkyO4IyL0gUWstfUql7
hKdM74LQC6uDR1QmtHTDwf51ey3dlD1AkamKjPpytdJfr6odw7kZMX1wA9ie
F/MJe7vDP2fakCaplEc+lP+24o7H4yluNXQrprpp/eOavl2O22Rh1Rrx7rDp
6j81qzmr+WTf2gy0WJUEpUH9QPtlD2FPfEOsVYfEfV6oarWvZYre/8WqVPRh
K5wQ38y011OOuU2/E0Zd5sH3rvBrm3lgWIbri/ha4hIU9KTA6X7kQQtlCG/D
IfhiC21EwpQARbC2rKnZZzet7lyGBakWKJT7m2P/c8wu9EcVuN63JniuKWQo
V6Q5J88MajpJ8eY8yheChpWFk6dEI+1fDvlwVFp9SglB+s68g8j4tn9LXKhw
T0gTMDldeOnRWRyUlsilBYeEKBgfM8M13O/W/7a5vbvYzcAM7PINAB4LxRzQ
q/w/VIfZYmgWDzli+oCWy9OX909LVHhQjwIuf5yN4Hmdznjljv8G5OYXyQOj
yg41xB/cW20xOE67W7bojzlICOYNE/2HM6OykrFV8KnTY9rqf0vQ56eiK9ZP
7yrHeFDhEem7pRgmIONTrlNDYjN9nwd3LhWq7jSLzwPr2Ch2Fc628jfciBeu
5e+7ZO0MYXGp8Iu128m/L4CMRjOsFFMjCYL8pVZ+9rbitfA+6V+odtz3BHhx
6RcyhKUtB9kB5K660rSmfca8WXOe6599qddlrlXQsNM/BNyg1W7uOWJatN9E
T6WqEnTkbnhAilGSZfP9xR/AiOZPMhb7JSmqKJqXghHuwNOjZkm0GE3zXHwW
laqIo0mViPVl0eNeYjGlDw3fsxVt9pL1FV93lQ5giFgzXC1oTM73sCQ37yIW
mZu5KWHPQUjDI/ssG+pT7D2yzGrm06SuihBoUD6/8BRLBEfIVNFEvYT4u3bm
h2renQS/A1jAR2b63E0YaVj/doQ+tJaeHnsUglHQ8scbx5UcqXFKW8VVka38
SeBPVRbih6MZ5qlzTiyEHBmrOCKPjaIRPBY2IkYV3reOj/WKKRVlP5bifCuL
dpGSB8INyqpKhCSDICAyutLddwPO8E8fv6fODZ3xGM7wu8KDduwlIuR/akWv
C1wbX7a7hf8PQdfNKWYK5IVOE5PHgimp7qaJjFC8gYbJGa7uIzsldK7hhjdU
8hY3OlH/5kJ0AS49xlpmB959ePdhLkUGaJoBsxzq063c3s+xZ4xGcLttXAGe
J8aAnC3VpiUrlG7lh3A508LDZcEb9NE2wfX+IMyNtpJISgxu7pqTUoE01cwp
zmfZ6pgbVM0BX1hbX6pIan+pjC4wzcOvypzc4tlF3gywqYxH8EYgNfNDasTE
PX5FA7vvIoH7wq8RSB1ovWW0rKlN2tE6vrNiNKhYPAUc35UhQDakStgYYDES
7pZUgQISZNOM5Mrasf1Wd1Fz8j0XMfsHLd9bXEwTePAM5L5pfYdL5z5WcvBb
sudJS6M12n1bUd2YA3Fn/9dsvZJyLIRO+8r62cJ+BYM9GpnkvRvpp5MR1dfQ
siuqYey/OUSzc6SzGw2rtBsOf092NxGkhZFBklGcOQYtdU7Nib9ObtKSU4kq
HP946q4qkL5oGXTESzLaQRVjPYusxTflh/H3eOfKePT14NXCRLuft8vldUkI
Sz7Pe5ptSY6hqXajaE9avHtpyKsAPNhxlOY539l0X/GgJgcwhz70aXlCNBFn
3XOVddSVl7JKq5ikvP0Id+j2Ec6G/hzlf2BwIJ0grF55oWFW/QlJjaZHYspo
opUoMQ7Foct6fWwkFJMS1xqRNJFOldLosbrmvuI7O67CeTnrMcyPB7ANlAiQ
IeOc8ITLDGj0aW1Zu6DJtU65xSs7i/KCfO5CvzDYjKKjCDcEB+z2EOaryW/G
f1vPv0750yP51VyQqShjMBouFe4auRIvsK2OOQHZVins1zjMpskpkmW+u2P2
HDwwQclobap0qc9ino0Vx9jpjeaZD+mPGDHEr/SGSnjOgPhhlLAf5Y/73FBj
r2zTyKQudC6dOnNy6yFyVhec8E6ZOYXJfJH+XBgfuUHxJ9XavxRRrn3UvtQe
kzR/flt765p9CgCdVmqRbrTS9e25jcwdtGnAundIEU+SAlrV8Fdqwx5tiVIg
QjHuMHIYT5CiQZaaOWUvmebv8VWKiA7Rc3HSZOHPrbkspUC89POcas2Z65Cf
kjYHNQdjoqZKKo3ftWGJTS4oQ1I2Hyrp/zEeYqZbIZa/oAR6huBrHeU2ilf/
M0DnQkHVy4ZRP3kfb4vH26jbT3I1drGFz/7ruZiG7AttbT8ISLRFGm1SeraY
H19uOIkvCkzwg7GEeszkYk3opuNK9yIm+8rmFCXOdg3Fm7zfnAXfQGs0gjDK
o2PQhqV9OH/YALTzY9ulkUeDOElh+t/gaSUsp5w6Zw7XR7XG3MYIgvD/X0SU
FxYjM4ZhgkmcjC3A8lVUxnrdbuSXpLhpGzShjbdQsQDcJxbjk7xeCpF7p038
320h7Kc8HIOSixGS6aco5fh9D0EoO+cdx1hfM0HDR7YLnfjnIJiMVvM8YvRu
90eTPhcCo4yTPG09U2BM6KK/TNSd8++uF9joQx3WwzUHTNp386y7Y5ZD3W3/
+GXewFrwQ4uC46qsuUau2MSb7mmqUZpD2V1M/E0UwztHNkQEt6nxGeeGxSZy
7JJD8DenikZnfWI4UqGamAIPadAF9rjzgKZ2BEmpITTcNC8tdXxuziuibqUZ
dGpVgPtvOmg1kU+TmwcVZyuIIgkIH2KGg2O4t/xgvB43weMrud+hpNjsunle
6ejvqGGEKn8Kh9qJP3dgaDx1cCDh4QeG6GfwDfQpNcntzatPeA/m0F0xt8e3
h8E9lUpXqngU5CXXvQqm/LEuqt6RadRTZg1p0+CQ4ph4tHx2PUDDTatQ2luU
WAFQud3kbBaKvotr5o+dRKNWVaPh04RYnFx/19R7zmlJpHZRjwLC4IHhYyOJ
goxi/mePs+hzKt8u6i+4xeJhJp6fUHFCE79f4gScN2Jsis7CEgB9fb2Z/1d4
LgVxC9LiKBVaWYtXqZp8u9A6KmTfPmShNQKzIPVPO2W49fbiI+LclNwX+cYc
vsb6bdrxnVbwUryVI2sZ959Uuv7j3ZGZM3vd5KZzXNNKqrx9e8YaKWOzLLNz
Am3wIcUYiCFU+lrA5tikTwAmjBJe70Swtgz89j7ngTo4S0n3beehHYjqA6xu
BgcSKOwHW7VV29u2H7pJJ9NVoQ6SbPbECY/oHsTQZWGKyappY+Ls5EJddAdT
wfUnaLwdICqRfmUYh8ZMX0TvxMeNGvB3ka8EAoT+8iY6gcRDaNNfiV9kpo9y
nI8SvuaQC9p8VoFsiCFbVctaosowbt93kxeeG0DT/gDlkYfgW0nb6GeXJC/p
0xAFfFNbwFULXu04YxPv9VycdD9QWD+qnnVfdHg99GWPuZrCECETT2xNvHpb
OGcsvZdIV7FrXGIeronTRiFF34Lvm3RG/wVmEnxKKxvwjh9nYgFqsKIBr/4M
ykEfBKxrDYicZd4HaOEpgX3DXcG+bRsmxQVrT8ncDhrrd2eCQr3fxw9cfE7I
Qrs7b35vPJk2afClrpek7OIaR0EORtIS9MWvUrwFzTDQ1P+92k9eRTID23UE
KjvmAu8+itwcv5rh3KV3YrUjzdFdj/ub1q6Lvx1PDZq8ZNiojEs0/xbwRvKY
eU8cGPYDqW96dnsqmwhOmo8VqtPSwYl4vOau/LCg45eamAbmVrQt5a3isIH8
mnYot2zBxUu+5BWh+BnWkHjqgzbS9Su1xoJ8m5foR8mxVu+kfS+kKRHfe664
kSI8tYf2T0P9iar9m4TzTkdGl52gA4cGTvw9nDEzGoYJD9e+eZVQm2E1f9xw
cvwr6lfI42mCyftTlDlbp684fu0kczzeTlg3LdfODmh2eTs4IkAHYPES9YMB
GQGQ/KFiyII94BsEDDGuvZjJ5Wo2siSZKFFZqq4tO5arP71Uvx2BDRIxIDzA
KBk6QDzxZDOKzTvVCV/J9+vmFuvJ/5ESVq1UqhsCQGOsnX57izEy3fiKxoO6
ry08gFjVlvag5iGa4+uE2c4Y2y/wgJuy/kULVhqMxEoGyviPdQ44qvHx0olv
lVYqnkdRBdtqptTM7Vl5cRWunUyAz83GShR/dK+rIVjk4/hMIu4qGwwyVLuN
t20vcE0NR0wu66kQlofOoravX2kBT21KPwFsA7F9fyxoF/O8Fi9tWdovk0Kd
HGm5kWMduNdMUc+qy303o6CP3e/GqQ9gLTJI4qOgaR4/1H+DUfCwr0G8RK40
xiKIzHhjpnqpGK0zuUZ7PGDMV1zk4wx3vXDeWDSDol8bx2Thnk28bHNXnNYf
R5DXs/36ysCjW6/sqwddFDRxyRkT8nOdeNfluEzN2GBVnc90EqSs+QWkvZ1/
vgxPwi0tyBOKfFHobcWo5mPWxtx3W91QrsNnrsn3oJkkVfpNtqobQBm9LpLD
PhvcdkQNzxJ+FcKGuuqWOMtdpdwWNtJ1N81qN8tBr+ZGU7NMU/cA4u7e63JU
0u40bt224jj31RHfiWpPI05nWXIp46tG6LqhnQSxn6Ht7Zzrpnfpnop2S7u9
MyD/2L1qi9YgsyMzaFmQ2TLnSZ3fvd/4MZ0YIofz9/lVTuprbwTEyuC10vxI
4KKE9bd+vbObBiTr9Gpe+gx5hhhvBygHKkRO1GpeoOVDkXrv5Ku6BgBRHukf
aiEA5JupixO9xr9aY4HnTzbrLlPu69zHTFbNGdCayaUpozeaZtIjJepqOF80
SqOA8fFkLgQAddiJZXP8OB/u1+BEJHY1TiWQ1bVG0VFGwDRJHvubhNA1eeF/
WwxW53eiQ23TjJIuWC4a8qYwEbJ0TceEFYiesCuJh7K/QHi3MNgrtDPV2Mvc
EKF4PzNmFfy4xks28RSF/7g6pAn86qMLAESJT+fLr6TaZczy9Emoo2ac/hpF
kH/jImeI/xEQ0/uDqPQ1GHZfzQvrZMRK9YIRU4Eud+PWk046lLciXrrZhUbG
9Gp+8oCNwLUeogp/v9Ih2klDBcsTojTfdO4ioB1k/vrLeMCNjqcb7AJIaoNq
pyExoLkCj3P38AzOnSqR2CkNjQ97vmDPWzxapqQ+fQTAHHZOuBQ7AKrz99HO
qfaUkTZVncf7zrjNsvonClaRfA8unVj7pwWd1UkrBqfgxu8hBGvXHs5MAVKV
p6d6qEsn/dkaLe2VIDjRN4kepD+y2PgWoSkEYQyM9m7Xjg4aQ87EJcV+dR9k
87nQOLiABNzOY4L726zw30xy7JNKkxORGOyH3etfIUSst7PrluHMXX4ki99S
M06+MpfCDIhhDrwZjHAhckufpRTbgyxNYBeQ0/rMBkZpg9R7cXRexxDc8Z/l
RjDXocTC63iN/CK8dHLByz4UUh33EnBUfQiCvAhrwbO1DrI+HXbfI/QkehmI
b/AxviGPcZF5JX84dwUeSZ5q7LjKqt3zKnoWnc6++uxo8t9gk1WmSEUJtoGD
w7PwAnRqsF8TaS2TiBvHysFSL0eca7HTuKYZJGmTHeYeFmATzRJ2XGsXubWn
np6YBDeNAnLu7qxk7rW81vZZRgS8CG0a4vWfcG3CHXuAmbogcf+VSF86o1f1
e+o7UB+ZLpchDXiIzjC9uSu1E2TM3dqR1/glTjNFYRdmXszOTQV6q+zfUl1N
UYbXzx1aS6YudTd/PWoB+sX1IugbiQcYFh2sGBbIVDYVPwNEXMZ1YDesDDc2
Y9KnC99Mc1Q82iRgp7Wrdl0vTuZ9vJh2Kjg/oNWjmT/b6uq/ocjbdDAHh5Sd
pQBaRiedjbF93hcxazGQPzwGS784gS91bv5mcLbQfUbGhpHnEUITw/tzi494
r1UTmFHQSiNWftyxAhZPw+zcFGmYid1G+aEyAcvkPMSAJDrzn4zfjT7+87Qx
X9cr8zqlPIyDDPKVVrJUCxP61/sSoqPgJs0Thv1nfnXe6Igo4HH8u0IA2Yji
V6DOlK0sTrvNZ7a4fJjPVmRfx1uLRBUjiI4pxp2+oyas7odXa02YWdP0fPS1
42CysqMVJDRvnyG0UzB2g9UakJ0FB3EuLNQiRlcxcTETXk1IpRvEAisBKkxw
DwVyUZGqt+tr2vIVRW3OIeO13FqpccNtc3e2iBWlCux/RRe37GQInVIdQjkY
3KmxFq25L/WD8ynsvXIUE0NJxvY7p4IGJUbjfcpQHh+2FNldoGmnwKu2jEZT
xLhgisy0HRwOq0VHcLPDqIBqH3pFNGms0a/D+i2zXP8gNvj6NhtMyqx8Z9yp
5Q3drUqrEL1eRcNHdPUqXXsf9AC0K5EpeK46WTYzzYa54mMFmPKK1m+qIQZy
94Lr/4JCkOOCxaOmBOr5ckSW7RT2MY5/W9xyV+iX8ELv6Av5R/Q1uZybCQuY
3mEQvH9A1A27ZMOnG5lYO29GXxJauUbxdsJuadSS7HLdfhhbiaoBXvQrdIng
0hKacqnzY8jixvlMr/7oVmeORmxgCx/EAco+BZ6l7BbxHjhObpS2mMCIiJDI
IqBt+WSejHcp+sEHS1W8xX/8YlK3NUDNvJugO7nCL2bRkgntx1m2Y9PfRkaM
RQkb4Rm/m76ebpiZ0DY4VKjMGd3QyXU7m2yhqobPQbOTBZYCBb1xGpM26p1H
1hzi41laENfnbUs46qaRe+tFJaNol5LrTuReGvJ3hxO5ZCik8aGcbktEEno5
Z3j138Amrv+MDLkfMhD4VPa3tJGB5cB3gbsAIZ/8QsE/nHslQ7sg8zn6Zb/l
NL5ifGgIJTJP98ydvUUrv9X/VXUBMHId5C8vzQel5CVvTdIW1Hh94Ftu4I/o
+fn8sWvtR+9pW7LmhMKJd4eYDVETxRGyRQnPDxPyLoV8DrX6312nfcnoJDmJ
+0IDEpA6ynzcQF+OtE6oQrw5N0o+7+k2WepoCPxzKPyDQN+kGHHQSXQdttx8
pVBnt0LIE7idYEHQdUdCRVwGnyvqzyL3mQZ/HTZDiiEktmrSqn3h3esyCwY4
EBE+0z7GDpKXLfRXPVvO8sjfUxSaRS4M4MSSAc7kUxvFW8nGVosI45Yyptpu
/9kJDe/zlI4g/ZdwT/f7bBlETVZh8pEbWBX9b9zSDEIEjw2tGsDxiG0XVk1m
JSXfVH9Bwd8yCu+QLuDs64XpQxNiSLqvEWglVlcXdYTBWyvBkGZK+mP/nyzF
0+1pEyVdJSbQ7kkIyMaOzx1oJMlBlT6b6sabsk/RrxQwwJA/pTQE8jjr1XnP
5J2eT3ERg/wy5V4ZAg5eMBI0RtAJQ84ns8+rxCBYOHncEBofdUG7EEnaFQMd
UL5XmMUl2tzSTzA2UWTYIomukV3+9ZQoVNk9hK25kg796H2iQYjjyyBpQoV6
oRO8bXOoggBZZ/TyRPwqZtRnGzPsESvlPE7H5scWRl/d7nFMpUI/t6ip8ivk
9HadFHgZeTUTJb+JtHKf2qeATAbjHmxiTwFHBRuprV8JHllbS2VAIOI8wXhu
R37N/tZpwLO5v6peX93qyy//SJCRIA9sJETBxQpPBDIWoj6rdII8+s8sxBn8
8KdeyCt++6cxEwi5xb6JE5b9trVHJYLXH7LHsXPeCV8GjXCMZBX3CGqAMsFl
qu5HPZtb6wpnk8xlxtmyt/eFWha+HHUTM5XMORiSYK8ZDyTz5iXamvINTVE/
nWWS9Dw0eMWfRkmti2Cw5kWqFf0HNlNuinx4L86vgoCjBUiUp7TFEIOA+k/X
qL+gbeWpRktRguSfVErfQrw0GacT/kkrSjOBHRklNPj00gpO/azvMkKe0whg
XawuQ5bpcpnZKl1N22RbetYFbvnO8Zj7MoD6ScU+MCSCAw2fFXm13XIt4qL3
lIKZdoSfpJ/bX0AZcxkoCNyXuQreirnh5nsGpUeduUsM+RqipvhV1t/3FVbg
a8XzlrwR/ZjaZF1JTbKr9h8UPW7WIumD44PUWnC4vQItnYaCGr9YHpllPYye
dHU3AQQu+Ojycg8IpVhcPihDlQ9xyw7c1/1cuYH2Te4hvQNY7AkCP26MmTZ2
ZdM7zXUx9V5ItBUpVZiJw9j63tGAYz65UT9RhbjKw2QqeW5zFBwKWHl6b3sC
PShURLcdEDaYGepooVvJbEwplE441h2lIAQTam4TQwwQAQFQJvy9uXcASlxg
xKaPRaa5JJE+nG+TOr3+kf5mvfY5aLoeYSFgT/LKjsAx8JPLR23aDMKz4rD8
7QJJDjik6GS5RpNoFndO7imnNxKtA9ce07qpK8mupJZ95hEzU2Ztau6gW//o
KCOWzAvXxcICOwlrkdBddVGCIApUzCoVfBU9Ls3p5BVGKvgntLcY5ZoVAPV7
8El5Ure58ZHXO00IlUVOrWHRip8FibrbNFoDUPyWtZGbu3hBQu87L79eD/1K
2nYzSiV8F/DrVbMloNd6GRDXvW19DIU93sgVHYtFutT9c2dBrOZlWHktH9vd
ArLE7M2nYBru6vyQKw10BueNRPPZDo3M4jgMgtX/BpcVUx5hWo1UrGWCeGS5
X5HdM7Ks7+T9UH2dXuokAn0AUK1WE5aOSPwdKChG3My5IX5qSLU2y7CL0x19
UCG0L7eXhZYWQvoolI54VP4D0DyYNeDkE9nIH8DQQ1q+gKJ6eviNl2z4ssgB
7p5slwvCTMiEW4VDOkOxSLXRKbjAXJ35S7CwcdypPGXNbRt8yY7HjQ7flpTz
Xk59fQUcfR/1Fj4r7DPxEF4haYVm4+HEmis3qeG8RRwhy6Zh5PNWZCp12bUq
Q1gR4W4+SR0loX/Z0YexvNQjq6CIK2FCfzgDSfJ12IG+LkhbmZ3r5Lizqx+t
5VR/6/MHGFccTX+X5h14L+p+vJmj/GWG3tl4XkqX0/tPgpfQgwrkgv+hRmW2
MmEseemkq348QnnNmp5JYing3ddsjdtObNJncjtb5ZNoNmsOO1HDpiEq6wiO
w9qYMEqGGH6xLTegF6VlJ75BbvvwXb1JJWkKl8YO9YkIV/EuLY/CBN9ViVT1
fBbQN+6AuI/tu0kAfoxSOSssBqrk9F2meoM3yUSG2HcGVASJGV8cxKjMFjVV
wn7Zioat5J94CrsUtJQRHb2lKsiavC9mSSQ5mHPVh9sOc9Uz47ZMvhGEKlPF
4bcs5Xjg5Upd46e+sUAApEmj5X12ihVDdTMGv2eP5Er/hCr2FVWrxWFCG1Cy
Rg5bxVjnSbS8wWjy7f128Or5/gdVO338Tb0QKfhCV5ol4vN219BXDmt50HH5
u5dCsb1U9ORov+Dn086unJ7achRgqUAf/QDe0Plc3Pi8G5Pm0MNEsRSvxOQg
x+wjwtsIv1dfXLObX6aTtQ7K5MnlboMTGPL3m4QbNIKrJKO3wV4F1OsUfH5r
kMyC155WWp8PU8TU7MLvFXX/ebhqpioTcdrLdBevqH2vvwd+oGRtn8J7tRRO
sZg3wTUOV7rKrdSlsQonqCxNEVRXymG11goCIPtDFtMIuR3vc4cgvUWnUFe7
TV5S795IZrmASaTGLbwEJU9YNs9xZdecbMJwnmaIy0jPBxWlqan8MGDKV36I
Z2gKGSwOsNSNSh2rk9QH6GwR+SSSNgbxpFDIkdGfZkrhPOMayHrJ8y+z3qkP
IKNwYWkcWZ4Ih0vlAJyh2m8wn0eXTlRn5AxibZOCU+NDH71RRvkW9mCdSPVY
sFU3+Dblum2JbQh2blesHZjxqvJfZeEYb0E+qRSVh32IGk2h0HnB0iAeqgCU
GbH+8mE4E/jkRCCU8jfwZlLXVf4DEecohN8Jc1bkmTX4xfo2huT3MdnJBX71
CtsXKWnJT03jLwWSrq5nbl6ih2R2lBKJz17ZGYa11ye94805t7g1IMvXWewF
fwbdtteSyVJ3A4JkYxUY15tHc9qRb0Cujb8QgPXDafONWRpWrFirShK1gnl+
88DgRGEBPwdwV0FOnyWLtpXbQPXzinGoqVfaeUeU5GEgmBZPxFOJ1lW6xFRS
kE4hMvGQSp+7QwjkCDYIOCBVzkI/7+jhpwTYOFVDiu5oi8pK44pO8BRHuOkn
XvtWsAo43QkkBxKFNJEEUYwbazXs10Q3DbApvF+Ys9PoKbq3aOpTQIov5KlY
tQ0Ckipia0TG1ALhKIqU5qReLdBVBjSEplmrZh30zvLwQI/cW5VqqPW4EfCq
txlP2j6LaQhJZR9d7IvukMvJ8M5oUuA9gM1NGSyCMEayWOB5GEqOkFj6WB7j
014/pvyNvPho5/8a86B5ENtTv7ret8g+cG/9olMzqPhBHv2/ToFLlIDalpFn
fRIyXFj2xA/mwDoBrS2HMLjJwb1OTrNOnSrYrnYIsd7CSrChDW5/vHXx7qaJ
SK6HMTnM9Z7MOL6sLatg+Vegu+8T4tslnOUAzvSZiRr28QCfwDa5NUvNzGfB
+Xnb3U9sPG3F21/9hMOCz5jsgLI48LxHorK3aI5GtQ4FNaQTZhNQdqTOHHMC
pHazqqVrp4mJ1RwrWKZGKB8v3vYouoxMcNz3lXNVwAWtX9iIq94h/L8XWAEH
+oZ+A7g20atIBl8C/EEAq1g3kppNDj/6CUHHPXK7TfyQ459r4lwhIaAWXsJj
rXzTjV7iDPt3gwpmPO1ah/rB3aOmx7wgCyZ02HSQJNpaslaLJMqp/6XmaqxN
NXOmu6k84KVPMOTLVZ3WPN0AEyPuw9OIwl0QJjdA/h63LPNjQS1Uw5rCy0tG
+Qruk1ZLoORFo736JqUoMUn7OXHsPsJDUCU2ZGXXKmwrW+BFGzSUS1hB6TV0
+jn8OLrWia3+kukuRn7c3i04XuQ3ND57UExjv+Vi4QyXBmeylhAAmd4uQhRv
n+Cn4au1/dhOTNa8vv5upcKCR0n/o+Dra7wfpD84fX3/OqR21g5YcVV72InU
qhb18fEdIXRpc57/3KsnpO5CkkDzaAj6gL+7xK23y4WGwl94naoSFKrDRitW
lDh308QOx/bhFtzJ8O7XDcCQeiI5NnHu2P/5fLipJXqLH0TFSz+O4w79B3M7
kqi19VlKYZQDBH4zwQQOj/J8QX6htsTrfvmh2QUWi3yEAUbbZ8iXV8RBQ1Fy
7Fz1MpnLfhDzXa6zg9N6frr+7/6d7VRo+DFcM/5II/qaaSWPFlpULkgrRsvF
bqJKES1uCGFn4LZbeYmWxiB73qMffIfqwuAYCON3BCo6rnunHKsZoaV2o8kv
t3OqJeLopUZTmBv0wH9U9b8AXYpu59wf/7wa9NJJXEbomUBmSEHqtIAxLBj2
lqkqSsZT6cBeODzTq2+ZlaYjTqVIUWWAb1tiYoMqveyUvyONY0qvDSd310od
Br9eDBzALV5NgrdV4btJbypkxRWB+NqErjM5qEVnzpwAgyCBurXUrRV16k+j
6Z9KR5ofCLMfXSHvwqfQam5HNPogMdUxtrO9HRyByCmwlkcH9h2v19rWO+SJ
vUqIsHBsKijg33qD7tTHl6DwoNeKxHvFBq9dgKtgDdEJ984/q7AAiO8q109C
E93i6fqxs1EHOmZpRuK5vTgHbhm9okDgAOx9xctJhe9ysCRhAKF2dKbm1JKl
rXxOwyRIU7mLa6bMOKN8hKOTllFnySvGC6yIZGKxIZIjtIlKmmBiMmUcvm5n
g5VGeA03pUHGWwUrjAi0Rf7m2t1sOUmti5hSYUOgjfp54U0CKPSN0+8BdxuK
HLp4LLtAuHQnuJY2RmS0WhJwG7Rej2t0pI1Rj0VRwAv8AUoouv9pbb1/IBuG
0izBeF6UoLTG55+JjGxsXj5/PGxcTox8LN3tcxEJ9d/fJnaVZCg6Lmc7tk6F
shfCOykFLGzkFlWJ0v9u+WinNWmc3i6rNPkFtFbMKLDWwla/p3Ud+glMa7R2
yHbdzVcA3MVXR/2h3BNQIF+jVePQY3c0mx0lOTBEqNU/mNq7SeipXVWjeDYa
5uXJvSxJV+9AT9W7/ITw5Vg38RuwTq5t3uN8kUY/AR1ErSvzbRMt3McXLrB6
uFMuwid6DUxYyeB7dLt/4bZjOY7VAYpWx9XVCHlXIdgR3FwgjNHlaowP5cO6
P1wpHMVH8wdSRhthZY22pJbnrrBfhdTqWEEoeD7rKKA7ynzjwjeidIqhuLRi
53zDvDjh9QSQGdGJqmHdge19wEq5NyJZysgXb5PABh0vo5a2rjB9YNNLCaIh
lEeHeo/48ST8rv4ur+arS+mID6RO8dvhXTvWmBEvF6LWuVdCtPKaoukB3TvE
SWPTS5OcLoY7H8s0LquaYz94//sgTv4/1puQt8qAPQY2OhGBSljApw9uXuOC
7fds0oUkUgFWhBDKdvpRnXHFmKUHEnuGZ6a50wAOPJdTCtF6p4YVHsVrRaKu
jyovJCtN1yWeDTB5h95xi6gnnBbfQqyvnj4GOfL6CJFRssomBakzRd2VAhY7
Ta7sy3NUQgMUzqmqHitCHR7UXKP2iYYt55fZL5rjYJdG/cSFJwKpgU+2BKGo
OM0PIwUoD2geSwHHp6+W+F/II8CkjiUZX2ONZEdOc8kRUEXbY8LHjhbQ94pl
IrOzLMu7cx/sGLjpXIvX3w/dTk4fpQEfUEOR1JHwpQcS4U/p19ZxuCbcoGoe
VT0ek7rQRyUDE/x7+KA5xFIDI66BTnA2+wop6rNjn9D413x4PIvR4AhfbvLw
HRANK2FUV7yYBA1uISN0A+riwWmpwQxzv0wqkVKmJGFQl5F+ZcCC8HXzlV1R
ld4BGphlMMbQUFf4e2CMhRUQ/jFJgARYuNgcsHDLd30FlOr7zLQzSByJw8DG
wXQYw7iCO3fGfF1bRfiJpc28h+vlzAKHkEWVqGICbqSspju3TZWWqgj3pQF5
6/1NcwuC577nQYvRtR2OGVPgNbAFidHMZk6OUgTsllVq68vu07CWet27sdnn
aWdq1u9gzooQFK2m4EZNKCcjcdJTKLeWkGXQaS/mz76XxAy2IUEXOXzmtdwF
ZeIUJcjduUgkq0MpLXn5UdfoNuThhPa0I+ZJrjMUsetcJwb9XIISZn7f9aTu
+BAfsKF1iKyVC71Xs3Mw6lCFLRySW4ymD5DvjrUbYYyJoZRBPwwtS43jMmN+
zGvNFvYl8GcsmmrI2Bvlyr0/eTv+fXmOMj8x0/ZP5moSPzS6+RwQQwHgQYJK
ij8aZlROgR7nZ2AA12k+TKc56WLNr3f1mtTHfQeA+ebDKEZsKYJnedZhrKz7
Q0VSAn9+LWNRXUojVG6VBgJxRrz1+vUNRqoFeqs7e28O+J+hT110SNW0GBmI
PSPzRgVbwbBciRGKx1Nlr7v5r4FyoSlI7nOTuTY8qZrp6BQdfq4NKxF4z3Lj
517ZLmWgkuS3IyqKuC81TB/ogIht96FDKql9/CFwKzRfGaw5ipqhwZqusEt+
2YRwhylFXSoM/8KVx5fZzpkNHGhuXUltCYUaowAmY0IPwrJbjUm57N9Nbjop
K4Cu8cIahNDKC4+oZmuIjUJMPgoOkYcZlSgxRLI+QPmJJ4+6Nti4Hts8sTtm
6WGfSp1xMepXEeiIkafzTWLixNyvbKMmO/XcWLJmW9zy+gbqFnbzFNMPSqJX
n7qVbS4j9iGz/ZcTpw6SNNuZTHJEb69Q2fpB/zWxM5g7KVTgloBUG5wRh7Lt
GiR4LJbaM4L+PGTz/LVnsK7p/YiVW5aChTgLOzgdIXQgf0LZ8YDEnHfdE7T1
yDxOKKqvBH5/WmF1LdWGSspjuImeAfnWLEcpw7YiI+2boqMLWL2/ZlRXq0Dj
cOLPPELTiUG2L9P37NDu/qX73bMJR4vpWOGHwE+YwV5KRHVqZjVaNsvaTf+X
4RJdefC7RovL9kPjIsOaFSmxHqxgOJRe5g8gD4nW6KskQctJwm0dkXzUOJu/
oE+5VXm3B7Nxxa+uE+bTDNvDuBgZ38PrSKefhs9BId8ykQWZHjXuXC3gxPLk
9YndA55nQXTCIvc/EXfTj3KdKXkyzqD1IZKCG3XKJbXmg9CKFAFmPgorHBwe
Fl/OLP4QlxusnIAVU64M6S/annTlEKXdL/yC4hoRawL0X1uNpXDgNwoezMYx
6TGeUo/yrGC1dLB3ZtGc69/hcYLj2mG8X5hNv951Ir7i7yaT0S26MfsYr3iO
6vZCZ47uwvmvoMg5L09joEMrU+s6F0DT6en8oBbgeb/xIW2Sg6rKq9T/lC92
2n8WsTL77OfiYWv4W5nk6bjDJuJvFRL3/dktpLsD+jFy2Rei2IqmFCIn/jXm
+wxpm+TTb1zPgndv7XYJOJOdnu+RLM111j/k1C6r4K2A+Xb0W9qcGOs6jsBg
NoAmURIIcVawVNBz0MWHk4StjIewQERHtlFOc58iIhTFRqlyqVa28/GnkC0R
9XPDK53rV8HCcNpwgIHxX64I/7uAy1vcxbrF9jbQLlNXspstJVU8L5UB4JiJ
O1hja01IVc33g8pvxz9zgdRQRDniKcK37wPytnqfSGMp/C0+M2QepgVVRPss
lbqQB5wUxtBfvVqLiDg2j8O88RekBVr3usYl+z2KzzGiM0DvEnQg16u0JswB
mg+kQm+D/iuVQS3SUEya3u5ve9ovaUobUHyPSj0idJDSityh0xehJG1JXxru
//Ge4qvSaWV/3q22W7aAjqMujJVjpkvB3QN0IH0eE1YnAA9nEBhzK6uddYxt
H3xcsE1ZkdoVicCfxS1Xcx4HphnMJReJe3u3v40aU/kCN06RvVA2QywDvFA1
wo1f2btTJ4w+KHIKqRlt35IDj1QIJdn02TQ2PT1EQboGvsZGowl4qTq1NmXv
eGkc7OmeyAjKA5/65/ejvjHABWyL7xr1Dt/d3QwsaqzyGkl632ystr5/gJPp
Vv+D4IAVxGxrE4LOSIJFLbvn+5hCYX14oFfBKy9nAofs8sgjOKmk8G7A02Ro
8d37G98a+GsWWAJ863G3VZ0TlBaQ0c/aBneGTjVWNH+kiIh9/CeswU6ZQ6dy
8jeIBuLU7/7YVfeT7FZe6fuf84WAJV6zUoYZME3tZO4cG/hiyP96ReDe7xS7
fGLjrVk07judk3x78LwKateK3DA9ZNi0xsEF3XDy2/+UmxeelZDg8BxuRKc9
XWbOe2npm551KFNjg4qZEWlqRv8gZq0F8GuxbhrHY/WOKjohBbQB1JrxGRcK
n9D9MCj93Pxjq8yH1ACD7b2f9u9gXskEvZRQYmgg9CsOlvNBmfJMgdIUPD0u
3Dr1xmfoDwxbPULADzHhP/jDLovaLYrRHNtXkKaYopR6Hyc/4IacuORYdyJ6
Bziv9KuGp07XIH52ceuHfSRDtjkVX8bZxUrgLY5IUauius7YLi1Q2WrGesER
zlDEcgyO43AkXXsB9auFMJa8tteNDlLFTt3Sa3VhZSX39A7zWlqActQr3Mv3
2ecpeWdm6491oWouf90winAlGQRK4m/kM41XUfHm1K/BT6dcnpDs7sAY4siM
dUeVOv81nEqTpu23hsGx2AYGsF3od4cnEswvw5/NKiNoQu12oExAfWNx2t/T
enAIFV1IkBy5+ueve4TL1HglR8Tjwm1Fjjkx+WcD7xniMDoV9/lckxz32wh1
wPYafwsMRfOwgsfOCYNegRQ8D4mWBtn4ktuwbxsID0Zk7ZHb6opp6RHUVluE
q6WtWiF+o23ILMZvBCuPdkCKG0Ez/Q7LTaTmuURGKxLgEWiw1qMCI5zcjTOl
2Zr8bJpZYdsCFIxeJvdWsw9i6Np399C/nOOEDOL6GMmwQgTTTZtqWJsSN/2r
8pqF9SMT8Mz3lib4gj1IZ0/YbROJcPoftoGpKjLXWyJcovgUMucm4j/l8xRt
lCLcXorY0Y/BdD96nJ9JKedNQpE2kLNpW1Q6tjqKvavhtnzpjW6nbB8QGAdv
UbVZZx0xRtu9LjhdM+tANi4ymmYz4LJe+2SIAEyD2SCpjJGvNYKv5PaXg9j4
UKbMb5NlQbUSeU1YkV2TeFOwGkNtQqy+oQrOQwzEMTwZjI3VdVSETdtLTn7U
A05NwcJXdZNHpwf7xgappvWFGBxX4TsdmIOqTKtqu7FsQy5GKQlnV6NdTX++
iqcFYm2+Toa2ayjkjp3R9u3lIgL4sLzkHnChkJCJ+SDfiA7n/LR451rXs3Dz
6UxrxR1YSTHYLTTjWjSqtsK1YfA02E2Zim3OHZL3LWnjtxxpKAqwCiPLaDgF
e0QOVqcVB5x8/fJwu122cFDk9s/UrDLVraP6mdyB69iiCrVODteBZhGozOw2
NbDiuoeTneyxNra2DlsD9zptHUsOscECyqyiyKymdpw1+vJg8uHqTIvEdR3B
tkwxUBuE+7JEkC/i+tbJQgf01Oan5Cb5O9T/lSJdxOttC9B+RHz2Xg7jsZ9Q
6JGBdA78gUK9oUe26yBcZFhXY5IRaOb7eT/ky6FxqgaG1cbV5cJWMxdvMoD0
fFdSjl4sGENCMCTLknDfy+yyZ2jpVk8mef1xiaSwmnPYIh9xsQ68va8IHt0F
LilSvor6yHJ45Op5LlQDA28WSMDwBzc9YehIqn9Z8WXcMYJrukAI5DPAhlxN
QvfWxlb5MVbNPslmAOQksAkLl6anNtTDri5g+jJcmgVxRD53hargFJbVmX6l
+qHfAJbHElmOHRiuZKGENJhW4vaLiGwIj5NWbws8BqeVT3O7CHFl0I/6bFmD
fnmn+uPmmdlunF3gf8ejBZ7DoqKDMryfs4L+7MeuOfhg0ToRbpbNab3OPMvp
A9JeYObw/Q6ZxSB205t1G3bQvgHZ6svq+zsLw7IFgbpcE1NfMASqb0DsH11H
kJ8ocJn0de3EUWjOonP1ZuRf3Q7TAeW9/y2rBOZrVtKNYm3t+5lR8Ko3NHBo
8kIES5vjxLIynWI7r+cKoo3p5IUYfZo4XKSgoPBcy3SpEZYLN6EjaYSe1Xeg
9PjG01WzEbDPlWVfJV8AXGWlwYMp7ySSlKZvErS+wiMJiSEvQtwdGvcl80Ru
yd9aagvv2i+Su9F4/kz3dWRL8mpR7m4mByK19Ew8Yj7iBP361CgOt6JWh47T
3XURWiEYLCMImnSz8dMZTXI+llXpXTAaT0/6OjW6pVzRI86JBGLsPg33Zf/F
bkXakiwlicbNnhph4BhCUOeXQHwPA9inB65RcHXYu1jS01wTeRHio8L9Atvh
5bGLqwJCQVpO7v4nxadZGWMJjzuEmuJRKb4AuflrdmyzlLt1QZVo2FsP9g4T
fzjcAJdh5Koow7gY780IuKFoSwxBabpopQqHlCHuuO6vQb/3k5mLCJOsxkqS
d3g/O6LLmUNEu3pmJSmaTHd0b4fVazdFepoAuyC43xuqMHjYc81tqJoUda/k
ZI9571Pk5PcyaDHFM0LcmFy+IXel13U2tkKvvHRSxwIlB6J9oUnuckF/FG71
Umq7oJzQ640znKW9qcUeFyvZJCViB4OPpmsCRaZdP4Qks+kFll1PSA+7CRp+
WAhCc2ch4Vr/gxXVFAccJsc+V3M4yizYlBxx1qQs7NpXIlgjBENX2S111Tym
uqarsWR66PiLKaWam4tH2nf/G5LELtijpd4SyABqw39fLqu1SKQRkWceoVI0
V67KLINT14u95AWTn1QsjJOPrPUwwQtllz/za7tNISv8hFTCaDc5QQr82B+X
/95Qtg6xNaPuP2rJyTgFJlzMkBcl5EbaAAzZlux0q9S/cTGFWw0/2oKrsaOa
blfuoj4MJFTXmZQ/LbAFNxx2KQgsi41BimZ14TaxCqIe/sCawiNA/TceFWf/
JJwbvidjhO+czIIoQyUJBlXrGL0h0HvMFnsO5XzSzl2US+3M4WJN7zUVSXPu
N3a3IV1DaUBh3w2kDe+31VHjoVPp2SuKyIXFpiyH6RIMvYL3D5StICjpIRko
eo9+82cLgNmwZDrEc2Bid9dWcVO+OgPkUBQIaiomZn67F894Gpb4sGqJc19R
cfGTwDgbmg12kfLZRMqDdx8x7M9DMobLySxt/FdngMBvKqG/uRsE8N7DmrCq
CJoniX3aTTYHHeG1xtTCXv5Pw/nAYpTzEwEO08Q5edLcSrnhy11bb+i7rXJ+
7n0D9q4shtEdlhXvFN5uWpjqzAnCL0AeiV+bGsd0LCVPID7B3PMFy+sNkmn1
ZTRk2i9l9Qzt/xr/7kWbpNyFzFm3KsGS/8atTpQE6wCQW1YWs04REGj8ZwP2
Yp24X5wZsYALPQ+y0wNmBam7YJOSo5t1+p7FSGyXW1Liext9xa/lcXxkuLlv
4JydptkEJfxmfCbVWFgzMa8JpM/cJu0ITjPDboUf6/FPyFopa/gKdYYm7xTe
1X6a0r13w9n5/2815ba4tPkXgTwkzjDpAIFFUiWWBIHh81uwSnfNzfFDAilr
AeqArBeaDRu446SJ6ZYrEuvkyTIUUoeY3O0i+aGo1PmgdBut2B+hZu10LMEB
7dNzoiBw/rKvj3Ae4pJP3CgnLQwTchWc1600cMK5/sGr8ESum4yT1QaDfafN
pp7ubu4jmFwkAHxiqzp7Mr3rdOlOiTduhMdx54j0Q/RZ3Xk49xhz3mY0blET
2nT0WzBLhhHWXH/0UCbxjfV2dTh/UeoP6whwRuHWYsTmpG8Zakm4YE7XghGV
TaoAI2irw9ayG9IiYdiluqhhjmtuaPL3QhL23gk7WNYV6mzjYVW1WNkqd2eh
OPAHJs01PzpfnNLE8rsepdz0YHH4DFYcl1TwZMlQ7u1h9OtjmL72QwXzWXWf
aSm4b5Z7Jm+pBD8g+INEWUWkGNHNO5SiYocr6KcikuiA6MdV9qh21n+AhhEB
c9vWW2nTmHAiijFDmwezPECj2520SwVFx7XGU678ipulMozajWjib+CKw0Ri
zO1YNdsfa9hwCnDHIR+lW2Q4cVlKLmzN9QxPkL7uKKMJfifwQVz/hess1uIV
CUXrZGGkIlETCeMzBORVZWd9VlvdqnIleAKN4nLhwRIvUchRnZ5za481KA2X
5zDmXn82AMmucEkqS30xJyCp5KpWvYguHKycL+u4dJbKBK37plHAMBX20SSr
R/HBoW+MmtYwEKdYrbk2pMzTcCw3Y2bKKqtZsozqfwdU6YKtZvHqNqp9YnJC
n6t0t6rkxGHPI1cFQzGNL97+phtqsZtQZIV2gDLwp6VvJRic/VnQuZpuguky
0llWGcf/8N1wBvk+Wt0YFLl6qS3PDZB14Gs9sKSGxZsFGC1akkcaKHOFacl3
2IvP+ikDmIDNJ7wbwqEolT+8qhOmv0yuDt21T6/Ahvsljse/wGpYtUTKBC9H
LdvQJETZmC0ZqAGFkr8nYktSLGE/qlrraqZwaFNAWfPInQgcUNlhj1F2QlPc
y8XWl4+f6bsPlwPu/qsc+3/AhYhsAMSEQvOK9yjo37RRTBGlU9vs+esSltfX
ZgA/QbwwR0Mt09UxTLi31qBC3kcEHsIYXANB459Et6sNTNi/KRaZ0vuVG0ZH
O7DE/4tx4O17yw58mzkfU3vJhCauVjvKGEEmMaEMRH7h1CNxB3gMVnibFNID
yFB5oakLcxfbdquzxX+WdtMrH1+50L1utAb5LsgMDjmUfpYEJNpW5UxrFSzY
BjJ8v5ZVhjENYK6WG3jlQZY1sXEjNczJUOGevZwngxQCVmsoWGMibEJHmS4E
dMitqhZcPjD9G9KWCZW0lnZLU9vLjrijkkrDP9Zr4S1kDcoib/I6mOjDj/wG
79wSWjedKTy8K2siAZ4GE2s194nVF0rj8HLeaX4xQIjewfsjeGoDOQ7fEWKS
wrvlJ4Gg9ZfcHRyx9JJt5Txx7iRavjpgLiVuL2cvjruhuyQFkMwMRk88fWPg
6uehsrLNx3x6eKUdF7U4HVFkCaNmz6H3WpwjqWCopoJMP0A2u7fV3kW5b+tW
u1lMK/O0rd4GjRQBdlK89I1XaPVIpnsvJRRwU1JYdaGRxKjbCzSC0VRtxc56
coWgG0I77D+B47yLMENuJ9uSlnYO6c3kcrtrh0Lx9XWRBUIq8OjcAveiKKid
SKFykvdAAWw2s+0JebXBixaf5kDe8tJMCzeketwibWqBSBsIVzjTb01PFY/1
KvV/j3rIQyEnNBqNRr6+dWqAvTtfgKC3saC3m8evr+4hQNjXv7HNWmomek3U
Cyq3OoMk8CYlJjJmrl5o8asunim6rUfOztO9eZSNu4OBQlELR1kSw0KGmFFu
I6NMpM2gXKBa9TKvuAJcOrjMsf84go+go5GwdZN2Kfc0M3wjuoZSWWA+Nu5+
b9a5kEq/HycZ7vAcvi5/jPhh4ZZtXGD2cKN3d+HC8WOoo7LmebyUucLDchg+
1pd2N1pcgXh9oAo+t6oPEUAQIx7so067EEwtEewb+InZjZX7BsHYIZvX6Pow
VQZLOtg4Er1+/wu8gwdx8gQeo5iblh4fc1/y64/cJ4HV3Yf5frW4R33HIkD7
rkdWSljyqu6FvNA8TvOsVP0r2y+IQtHveauLgiS/udERjCYEQ9OyYp52g+Zi
JMHbRbDShPDyGp3a0Pma1dsWL2n/BKY2VZGfxk6G78Vk1axzyq+9m5I0Y31a
FtUnsJ5tPG4cxFdKT9Ghi09uQDAD/dbWT122QFJMCwyU5pjCbo+7ns1eJgyh
vaCX4jbvZJsxr3TzmgCkKZk3fE0O2A50CAUaXGzB08zYIs5xV6/zZ2ANWtCX
ZnUVWqv/weeHoK77QFhCHu2YyPI0ItdwPCtBEozD2H1waMah46fCkEJFWJVi
FzW/HGOd50luoAlHryGhhyou00WNoz1YiGO8yvzNRAbbJd02XBrrOLHUmi5h
n+4paDV3g0EBOlXGWGIXVFqPzofyxI05ayYLgJkwbz58cD07ME50ZixjrCZn
jU3i8sLeCGcnZXA1QmRLhNqWmAB5fIkg7psoUND3voA9ZOtcoGKoFnolFXdl
C+o3yy+YSlsDK5yz08MCAJ1qL7wx9ai5KW5HehXDUtf8SrvbFJ8IV0iAvVoZ
NPI1A3vpLBg4uWxZ0Edt3eRTwN5Axjv4DWS2z6Dbitdk9Wlyd5RtreXfFzn+
f9EVfcKPKg24x5MS+djiyviDYcVUXJWVNAXaCInSSMU0Hn7w/SITpwvZJJse
uAteO9K9LHhm4/X7Yefj1mXb1Umai3NE2yQfv9v+Yrv8eQE9ju40jQcday0l
MHjVeGA9pFDMS8PmJlWAvlXX3LKzQlhrqNRnQwuggQvVz5XjGbjIOT3g5fYG
jAGYVFsHBoNzOp7bXllBXEjwcS/R/N3muf9vC4OxHI/utXNJcFwgVt0XMme+
rO8jY+UC1Y+eluZzJIFT8J9DYvgPPMztbHsAOr25/YduH+YbkfsL7KDQVoVH
lxwxY+9p0X58GgMj9J1rEs7f9PuX72g+mmIf+ynyQDbbHO1MdN1e/hTEodoH
4yqApn47xt1uoZZkYBuJ42hL/wH3ScCv8dBe9CXgFyOPfETEj9gI0jQkl+z+
W5Clbk8jUc5LeWYfIfSAHxNsvFEusuf6AVGqgJySprlRGwmW5/FvT0grG7oq
gMcSelgNmYaDeDMfI/TW9RWWEKRZjdE/yLqp8VxLjRdCty13zyNlOoOIfcr8
Imv7D+9fO54smHRdYjfkkZjI2KF4FHjrMt/v4COfmi36MySvhFMaKf5tdUY7
zFoHlPiB2pXxYw8AJ9D0l7/aSygm3jK0IddN0DbCidff1JH0S9Vw2dgm3L53
J2cjkGHJ2x7Cgy+ON8KgJCfNgcdg9WJ/bPZpOfd3Gi0R6GeIPRu8FH8S+Peo
THgwiYmtItVxy6VNEXLI79YiYprT78KOF0fcuYHya7WD9FpoQBANlzp85/+w
2y0a7NUcT2VjokxYi8/uB+Ycg7eRPejAwlFpf3/OdJT2ydUL7ZijMetJd6Og
l0NKsSfMMI8E0txsOnYIcgjOydUxbNDxqFCa5exVRIF+cisw9yY3vFFNSnaj
InGdTkemGcXImfWP4msfNp1nJDGZC/7uIxkjp174nIt1EbMyLkbUPw2z1VrA
dYOET0kuuwi0cJ9dyItbu7dglyhdvywZDS3L7DX/+/wXK1kK6YfHkuKYe0JH
proKA7Qq6od/jft+g95d98PHfBh7WODp0wvVL0BSySJnMVsJkRyVzDMNxXnH
zOmTJkF/J8VeBuSwmOJqTDXVe61bl7cgeJllMV/QKDJyfdnkrgCPezzqMvh8
4XacZxvqCWy5xwgsA36ptBUtgocw3ACAQ4CiqBR1wuf92K5nEJREjNSt7KVP
48X+Qy+JkSZ2Mu7fHG4x7jk659U+NRXla5UabO3e5XFo5pvUoVrwWHw9uUSF
0TJVsH3jXTfI2hVIIF3xTnt5U2+kudFrna9FH0vTJlLYB6lP/1hrcdeMa4sh
PELbmHp+8iEBaHYNm8y+/w/aGHjJOfELKpbm2+7268j41gdO8XMpayff2vCC
y7zS+iRCqgAdxjFnUmuqjLeWguTw9h9hxRkcZTNV9bO4/wVqr25AEC6sGrDJ
2XB/ai8nD661Drb7T66GEhmlMnYIhti6dvkrOgJ93tUmuekf1FSO8M6kusP1
yUY2SV5qfVq6kodmhrfUOkSYBVV24J8VuWSi94U+DpgnhS8q+9exzJb6crap
fzaqihRWNnXZIT7Rv7wI2oXfyTWL6yCq79xD1ryzeKNsuQJLk38hy+P8Eutr
FCF66OaVU4VhAWr2kP03hCe6PxEB/YMzhbb5zpr/GNaAm6L3fIi2OwjT5Pb6
PJhAL91ltjjgYnhFIYOWQXVKGWamY2leZL0/DFdR3MPT7DgiZlD2KlYvKKPE
dhPmvigQzo3Tcjl7ZjYA1sFDeu/6qlF7VTnHzRtMTfkeHM7qvvE7BdFiyMKN
hmb30ZwJcvVnLLixE4cibLPbcb9PUREwmfnwly+orvQjnyrOIv5V7DzvvX5y
MrQ+GHuQ0A423Cmaj9Po4i6AwHGI5g67TohB8mYdfr/TLKoHCbFyZwrF197J
5VFz3IdJnq8GtVkWfSzm7DriUPZC7j+nyCWNOttLt6mJJV+aRQFcj/G//RRc
iwCJ6/J2OhzNCOfvZn7wizp74hLEKsDHzfI8mAputGBY5Pt4fZBFFHo0nCYZ
zDzylYx/jNolpTq52nnVrNkL68z+w7znTW5VKu6ABEh6mgBzOXbpp8qBWRFG
+xChixl4kebq+jSQ/Ox6F0mbK6ZdaY+sdCdYcAxLzf0zGSJv+WODHM/KYzri
ZCEi6DYSemDbm10zHsgiQCSpoFB9/b/KMBOWTwpuDTKuI+pp7w9BA5/t3+/N
8EjnBODRLaIxBfISMM25//1+3cTY1zDbWCH8ZD5BuipXdXdxpWJq5gHGGfin
rR6lIUO9scGgQSrZyXpcfCMdoSM3WpUliQKjYby+QtO6WFJz1FY/gsjvL1Nl
PbLLT62sTP9LdE82HZKrVrkSOkC6SWOdDqVu94W2GLjI8MRKkOeZnt8/Dmrx
9I3rL5VXFtRNKVsU5rF/yy7s0HAy4xfw612sIwhoaW8t/k23YDAlTDUcB73G
tgwYaL9b+7TfmSFUzo8Ow8vpIQYGtfS/phgdRGMsO7lRDN29lTa3cwvgt2Zs
En24JgVQnk4fF/XvkIp+3VhX/WV1wGJM0iGlDe7BstZduWTkK2vTewGnT1Gc
c8FgivKvkeo2ppUooj5Zuf8/aVS+0TnruMw58Cpu+G4B5wb10Wkj5/xcnipJ
uU7sxzcbMjqFNdUGRmqeSmHlHAYUtvB5UFesKFnXXMcgDi1ukCkuI+30zud2
a4QAp2f4C0S04NgHDaAUFuYu67jJejduKgELMOoMK3OIIn9uCPntDdVuORgp
JQ2VfSDIWTI2PDKBT6bbWY/XGhh+zGPycJBSUiY1v/2+mxFsHT36TKQC5QbT
eDWYuwvD0sB1QgHP/BQTDcVneHfdxLaUwoeOFFQp//cvpDzbBP3uht2KIYf7
wy0XfeFIcFa75FMALrQapOMJjYmzWmIi2aHs9MgaNl6bdmtBuVbmUgJbimP8
EAmmsSE0gSWGtWSuPo5OQ9tj/O08QXuu5R9vjnCfCG6rV4KyNePVZ3KGEdpF
C8qWoYeJmHgte59tpHPxEp2lG6z04utK3/bBjT6q7jKdFNAJfxBlv5GQ34zP
2uLl1aM2QBJ36d2rI6ouJcL39iuwJfD8YywTfmkM2XvzngwJw/E6kk03cTgu
K3xcTXi0MOcEuCqMxq3Z0APyKXqj/UQzEYuyiQCxu2322spKVMcJcedonUMj
VGwuE3VDwvzn7R6kZucshpz4AnfI+xYzX4oesI+/OvE/Nla6lSIRig1D/xpH
NmjR8MRui+yMdxY2P+SA/S6iCkLUP5dLtxFdVtC1y4/zulipOvXneoWY/FoA
xJXCTU1uKMbOm9xU63tUwKWFr4nllhVHGRE3g6iOWGaFPl6u9OTmaKvxNlV6
gtEAnUYCDu12v+JYsGIzr0rTAiKWAZ+THKXmlHcg50Fqv+jNY076ryOWOIe0
NESDZ/LdenFpjkHlPhJnd4MbsnYCIeBBWE7aDUUJAq3BYGG1zX9yDBEc6OCE
ryTcyh1Km8Rz9fvvGx+4dVGXlNhjxV+vVk32PO34J/aaEDkRDk1B9V4270cB
IGx2Z1AucIMDhM1evzccyq5d/VeR4f3WJUVM5hAbCGf8z4iHsUPQB2EuEY7V
lULtgMrfePZEWSuQMAx3nLe0S59jjSOhVH0h7EcZrXOHEdrgDIkZsaGOkjOP
Ahw8wId6k4OOnrKjCEUvTu39YggNlMYYRnrnyr6RGDGQdg1YABkqDD835gxi
LcdabzbSCjtknZynokXXSVrX69tUohUVEdIS9k5MfgiZcBjR+k2SjsavACbb
XEkfoAV+G31CsyFzMWcBX7Mx2wAuH4L1PCRft26XCcu8dcQTQxLVOjLheDRO
Y4kgTL2h2ENWgNcqEeBC5VRDghUo3GJXOkECxBvlh7+eEkqdaFw4d8Wif3+q
+pXJrQ+K0z0BLB6/57pTLrlFDaGAY4eYx2cZeuF8/UG6/R4eexEWnetdk8+C
Jy/sDuaW30cE5mlIxWJyI07mq/bTV6waXK1S1MO2HglyDQpFXIUJ5Q7O1hiA
P46wAaKXqgFppqJXCkGjFAAwK8R5tD57OcHwjDxl/6oO6vTSs/BeQ8u7Hsww
3OtYiAfH8vrQ+mzGNcP5ndUtLkW7dzEUIQT5bukuNWF2agyd2/egGs0Wt8/K
DtlwYsboMDA59MFIeyoMSYW9psx/YRkyn+ic/NHklUBFM2rQIuerZdH5RgUK
LGA1h2rM922vG4ch/dROVJB+l8wMZxevicF8TF+WzKH/csfYTiK+zeyFxqdk
YouP7A+ZtIYtklNKUvpkNlbLx0eYsRCqMmRE6/+qyJSa2t/Zu5mxpxiBJ148
qV6Px5QLU8HInnUTa/IjQKpm1RUjA43lSO6WHbRQcx4BCXHQ7wXzaB4kLe2P
eJXiFCgKkfTlmOM0zOn75KLniSRAgRYsWx41C7eBZPJ6ZSe+n8eFCk2lxrHu
ef5ZoRMCPmYLuEU8NFbpaq1XN7pdqja6qSh5pGAaFxYSKtlE+zwn6Q/lXqUi
LWUdgZjzWnO/8274BMf1bRUdtQseQVdkQxqkIO39G7O2ZwKgFl8D5xlw8IOf
t8r9+FdIz2n6qzxyBvivXfnt96X8/Xis2n/Ifes+4Ii6iaj82gri75By5Vbs
xSjjKi93VR+dNLJDPthj8VEmWCMMKMlIEkUsVR5JlDOAaAgfk1W29Kho3Ifz
teayvuKWU6oHtkV40WsiMoPXzQh16UbDhEveSRf9ZpGjDUyK3xqHeRWmn8mx
KsM42KblCqYd+xNJxsuOfVwHjU5mI1WOF3xJFGlEYTSO7/LSxqOhnjIVp8Cm
Ws6EIc9LaJfD0EdQF7/SG1CnBzgcL7jRCgkfHcjD+CsLprQAWkX736N1FY4g
SZnprc1C1WhqjWw+NX7QFbMvsWFic1WCLwtjFEjibqBGR+2Q5IfXjdmFddi/
mN8IvQvmU7YRYgAdkbvxztP9UQERoxL7I81CJ/3u/G7VzPWjtFUkX0UoSoXR
oA5uATWwhbItTkfa3x9PekVYpcbdSsCFFNHgz1o1kwXFC+aNqncZPL1QmZKm
7P3+QycJ39wAcJISHrMYN3Y7r3w8mekbsepSVwxj4DC+yi9rhCcr9a1q2/hC
wVyTpJv+AGQvIrEdUp/wdJI/kxC1+yUXzL8YGkuaLrc2LbqY2HAC00ZB+y5T
MxyOV+dN5iSX8YcohXy6My9CI4doEtkudMbAXUxKkO82fw6RKVefMvuw2EvP
Przw0HF3893AI7GGUC6ZyxrAVGM+6KJhLRkMGOScKl7JB7cOtMglNOzpF9od
gwkV23jLEy4PpHnW0zlL6edqPYJxtY1up3OMw+0XjbiMUmwHl++g31brhoN9
eFk+OvQuwjx6abkEZma26+/GqidAOTgZ31BamcY5auJy4mq1sd6L2NWxyH8i
JYb+/KtGqPMVzkOh5WJDGP+L9uWJaYRQ+CeIKEJTKrdo8AeZ9l80Peoe8SYE
41bjtuWvRzKPvRINBXyCr/G5pClS/ZgMxUDLrie1fp4qghnmfCuLCn1z4Bo7
oq0gQdPQITUa20SYz2FhMYpelZJqSNyZY7iUvCEmxw6hlRHEp92sTeJuYiNI
8KZirZxaK5dCP7l3fDiX8i5v+cryaQnUA3jckRDwwz1nHaIPxw9JcOf37NN2
peC4Iq2Cx7i9xp7ucoaCIJW2DLliqphyvIBt3Qdqd7+SvTg2CAH7vNC3sLga
mKw/UvFaQ7ye1jxx4km6UeHO2DeOXz9kKNvsVIUz33xY7XmDit6YobAysPcg
hC0c+88/ph+blMHWLNwcGj/4o2mqcpVGHe5RNzAg6keLljCf87TBNFGhBlt2
7AR0CD1ew2IPFwHTpANIfHKxB32/ppjGMrlCF3KFViq/S1bFkQvUhi+DzGzs
SHha82MOgJvw2c4k3LbTqx+q6plh/zhf6Qgyiatf+8oxfsy46qNSg6ZVypyP
vacD4bvXycEgnDQRayeqZCZH1xQKkuvPvPFEefIPvouulxzP2ZMgdWub/Ksf
Syr0l11G9B7gsGcEvRSVt91jNA+aTFhW5kHIP4WkY3FcVmPzbHhEOoTXRk0r
JHbPuNo7RrUA/JuBMFIyeTuOyA9AIm1yJQoXkzPK5lyPzxF61/HM/S9rga3b
Q/Wi8uIFaXmSesJ+1hUAGq7SugD7LBbrwupkWv/l37PTEodJIrfhGp2Cqw/5
5xxlMWPxap4CGd04xyjkDQSIai0M9FY517pFXE81bjKYhGdvl3TanhXXXacp
9V5rfxDJEaCa8iJeBOigZ44zxgwPa1Iggnf+Mn5nwwxk2fMU1+1Bz3E1UOKl
WKX9+8rYeq8Q7TSlDKZuruMj00dYudGKm7+kcv79BGsydxZUKz7705aJGDs6
+BDP6xxjZ1IPq8wbsBmizwhz7qa0F3lErQ8K38AZ2/HXOMyGOjdjm1X3kYw5
dIybILY6VzL7Slzp0WlVdPBdVhpS4a3a+gmQyGHXhEvbTF97ZJyGHMU2hoIh
VBeS5SoA+/vD1RsNL3vBVUX9fSJMX1CquwLwtw82Rh7IN4uqRpjPbiba6ixr
noaRe8u5LrTgRoW5G8TI3I6W4Du4DbMZPFd3CNywPpO49p+Ai4HTskAabssF
TmYf0Dd8nzEuc1HHg5RRbembPH8ROs6aM8XnoKHwaLWzZmwS5DEwdyRzEDMJ
JTb33Mogtkt6gMf2WTrRnZWKRsBcEzfNxyQsiPPBdDNH74bF/Zvz41nmUt8J
J1eXYe2mnbVysS+9UNFXXCr6HZE998V3Zpa5BgesisVGVeWAGyJjqGWF3bz5
TfPjZDrJwOnXP5PjtbLjAniCdfIEtqHhpH9n1CIa7+Ox7ZBbdMV3vrh0UrBP
oH3czVrVjK0WRQJCECbPc5IAompusYG5LQo598bct4H+RxuotVHDSUXgati/
Zo5E13WBbsXtZCZlrnmpywty6LthHMZpxCbMal1Sz7FEPpkcSaEhK2S/9vBc
PRttsYxWO+cCgWw/rymUmLRfc6wWQgOrcUQvySTU/PQP/CBzdjzLpp4PTCs1
HnU2vnzylyAIyi7YFMJJ5Eb6O3FczMYRswH4Yd1Q+4qCG0jl6YGgFyK6qUHO
2L8xXtpJ3HJ0XYKu5CGlGRTsmqFUEBydupKKcYJ6sqcKb/ZePICphvJFKng3
VZl9zEX6fSTOAb1QLdmkSXv+VbSL4XU+TeqvUZxU6QlkwVRPUlFBlUQBJROn
dllYViMR2pAZCZHXaZ7pJtgg4Lz1PacPllwBr2VT3zWKEDRBvk7RAK47CA2x
KddqVPvL5Wv6ORJAF40kp8kZR9+FhgbdFpvzd2RKVEmVuluNr4qhwn2aYM+n
rhEs5NGwiStQ6ulkE3YoHwVdB8JO0ZdOtf7S/R/8pOTwkUW+yAeGv61/Gejj
yhSqxxkxyOSevmQXU5kyXArut9pcoIceT4s6hlJScP/3z+wHrvcm1FCa2LNT
lYpOyCyq2W/HJVuVOTFkkjx4O0vhfQPocm4A20ZAzdght0lMbPd3JKuKnDXI
5EitgSza0r7gcUaZ1RZH/bNWWQ7btgrmpcrLup6lv57aAGplQlnApAdnIOyN
HpX0e4a4HkOhqvsmiqBnC8qqwyyhdnL/20dXED2RUVurnp/zJ5oN06virl6N
kxMK/z8JHpw59H2ILkcyG5Ga8cSgUxVz2V6ki8NqJ26JskzNQeFFQ6/qqZUD
m01SjYmOLtXBJ4XkXYxta+2mkOy0mI6evSTtnPqdpQSoz0qH3tM6xJTdqM9G
Z3CF9CzjCbtdZwvqMsQQoW6idlrYB7/nOU6OLdOWhfvDHI8rN5dP1yTjcKQg
fIoM5bY+LTbdTdBRVYuR1x9N8cR+FWtsxWcJkXG7NxEc47lhEiKbG6Fomo6D
2+5zN5F+LoETQMGD1eAbiCk6MFwjleKKAihU2UEaNavU/wR3jR6CpAr7UA8W
f32+GaUm14IxhNmeNT+/aQnOOZRAm/Q7N3UEMr28laSaeDoAL02KLpLwyfvE
g2aEA/Lo3YwTulN3l1dOVetKexhcvQm1r7wZoPl7d1K8Ih5tKkFSPrvNGdXY
na5wyAFDziosCnmvjv8ZuI/ohxaikhOhUeU0g6KfGXSXVz4xmgIa0AbnRfvY
eUQ5gIsbv8YZ077qVHWkLrFeA9eZYLGflXy1E443R/aFCSGGiH2Nzx+eEW0s
CT0UECepzuuKuw33RyugxLSyjTLzSOINJVfI1GiY1SigjOnjxa8MQ2IShWBu
dCiD0AgVh+WaDrbHPMDXvuwlTxi4H3v0CBjniwz7rxds4Qeg9Y1KdLo2t+p+
JNwEBUFQFaLF7BFYjAa4bLnO9H5dco0tN7KgsDv8Zt1QjXxwDsrB5iDGG3Wf
hG6e5CedRhS2aU1S3637kVK8Q07AOmuud8uwPQYd8D0hg1O0+M0FidZSEaaG
60equSLCBopocCKL5fr1Qzd+k3uUMlDVPzjjbweldl04FcUMXVhil0bUbM9T
6qttNU45g2zB48bfZQiuKg35PFM0NV7bkYDEVKcMvdSz2+2ojeDo+XG4/KuS
UftT75FZw28moT8yLSw/55n/XWfQ6mwKyrYbw0difBRptv0DZNXl9DqsfHMU
6lXB1odU0ZciLMiMmMpAkLgRUKemYZBOgw6iQlSXkvVEOHWuw6OzDwf0tkLs
/V4mKnJQnMABXg7cxKhSuS3w1+OhzF02cmXkhuTvk//dKu3Xh16DjqIpKnEO
gCtPrbpHAbXKFb1n6zoeba7kTeUs9uEhGFo9LcLYhw2elZtFsfTjtXhdAANz
9oWIe3aIeYaspiqQbN/78K9MVPjjeHE5NmziwcYzhuEIrR5U5gh4PqYCMzIL
CGY7MDP4IuAJeP9JruX6tlm6B2MPOyaiZGBqUd+qK2rBzYXaw/H4pwSZL5+M
kjDhMHfLBF5U72BRrOiY+jm9mmSkT4IsO54w1XQhrxAw+opymQ37fsFK4wb2
aL1e2+Xd0/OKo/HUaltUk3T9om7JrTdCm1WJoy4bITEn5iHHLs3r6iEo1jl2
rKdGkHVE7EXrDY2V4zUbxc/Me6aurnO8fb7l8b6roAHs4f2qDZShjxCeI2hB
yVCt7eNocSvXDujRGAw6sifLGbgrOtsZBVubWabHRIYcD5yVu5x1oPxontrF
PCsxhy2z5TzQ6fhR0eRxsOL6cQ+ZbvIp7nOvsYGDWWwIT2ICeJw68LP2+ATL
4dRgDDKY5il8wq3Qz9yJ1zEQtFAZYJ3nc/A075osDpo5o71dbnw3czpiH1Zw
hjk5JHJgyNTnux1y5MSvtVua+dVrjeEKZxU6ngD7rXYgMurlMG4lqXr+2Va7
hX1kvHXUj8pkoyLGS5pr/itENSwfrp9Jc+0tMaWKrcp3flhNCQSXjL4jyjKc
o9gwfNTTZLLYMnNLRmQcuSygthwUxtjWgMvEpSH2ZKxMWt/3L8o2HHM5LQGw
tomBBsWve56g3yzHA8WjSco5/8NN0KQcLqcFduqi3HfCDxka2kl37y5XmljI
m6Saud5VidGo8Y8XAwgTloXB508wQj47RbgD1O/DQFczlGqJ5UMtpeZ3w85h
i9Gqk7iiRq8ABVzClaPUD1gAHSfHtQSLJfCCzw94+Ei5rliFyKLwfxxj5cq5
adkiPUisMQLGRDrOMGvRZ1PdlnnU6PWLNodt0pulz6n+uEYgVqOD6btfIfAH
DYBurafP5vezzpyd8wd+djAn+NTWDwJ9xW7mYg8v527ObLKFuNGUYb5t+ZCu
aJ90VPsxbJnZL2GJdEFLcNZcPi3fYUStW4qZrOaL0ZbtGUVrDJufoQyS68r0
ONejTT7QAjjruk9OMSgpqxVlloTry5ivdcRY8Oa5XJNZcdqC2XQKi3Bfn5bF
/SERMZtR9PJ1ZC4rRlMKgr/pdQhCizh2UF92Qhprs7TW+sNKYc1B75rZ3BSH
UO0ErkCHOyuvLDbzTvWnz1Buy9gCY7s5TXHwZEMijvCh3Mr5v9EVlXlw/TVJ
2xZUmA9okAdTK2KCTuyEfG7LyMPJVGHgcewFliPkNeThJnb2v8ihnLaRJXk5
6UGd9IRVpiZwcxeO1sAEWd1tomjLNjggw4tYAXD6MGBxWOfaAtnAeEQF/Qk3
slK8wGH2prg6jhjhBJXpNP4NHhoyW9TQvYYMnUjiDQs1FenihlxNhOumluJ6
FI+/hrxRYpg8qtsgbMaAY16lq2F0Z6vBiH2iHIas0IeLuKOgrPptdtCnrgOu
XrdJUrJVmdpWaIgQOI5x8Fm1Bp8kOcVcto0KKUWf9OYgMwl7y+AA1I8Ddkr9
30z49xB6QgNd2pzf33VMGmMNx/fB8FKWJQCRtIpGgD3XFhoE0TbSd2tZtZ80
jdnNu2dDnIDvnnjwy8HX3OQWU3T5M45dtRTqzeLKVl1WYxKrNTWQKUi80zuq
bO0JtIy/St8dtV087oq4FZdMAnyIgfe5f3FfYR7mfSgBR1CmakCkY8PItUxC
PiLSH4/HbZkfPy9Nnj1zbWIS0Kd63rXWFCe9F04cYxhO0ggUOdCTcEMlh6ID
TVUb1p7shCrjRAvnr96+IqL4MQz8HWAd/nCYO0sE5LW+rGmBTBuOWnPPmn6t
BYVXuSGcBqm5OgL0cnbBu7E3tLe6V8bI+BfXDsug49+sn0VR/0YivqoGX98L
IDWBa3Pi3n3Wnh40fYKvui5s/Vd67J0U4W61Kq4+s4JJEIV91hh14f31d54M
K+9lalWa5SiS9La4tljn1j738Mue+YObHCoQhOGQqVlc7ZjbXbjy4+k74cwD
15sKGGrE05M6hUD2AT6SHa2g10cxnC31AV4who3nfXXsu4dV17ADjJKPvF5Q
fptijJNCl0/orSlsB7EQju6hz9MUsKBV7eko65/VoYE7UlPayy8sdBpvhc3C
kUxLRCw0cDwTZURMcTxmHSotfkHeBZ3Fc2vZxHbwEv2A3QRtVdMiQZ2W8Eti
pxYuSE3TARuc8LoLNlgDhzX7IhB3HNZxJbF5HjSM60vqO+adLxuz4xaFz3Jv
NlP45Hhsc8IXYIsy/ulIYkSMEX/r8UHVGl2nX43Hkh4H2ugFne0t6n5bJwCo
s081d01TIrzwsQkQjwGG4RsjzmkTipWqJY34zudwCgm+LlXKaakBMzjQqmPo
GcWU/vYdKk+2yEE1MW1c5Py+swpT/m07/jn0Hc9kfSTwRvabohBbXFkUPJtp
/M3dmb56X9duNhj+Y6twf+pJd6BAr/ZvQPrOL5iQEgpyENtXtobeKrIg4b8f
ngebeYJo7zhkDHrLFVtWdzhAsDS1hKs9+EipKkc5ylCs++Fus7Ij5wBrbqVG
lTF/Ogbv/JfxBpydXUOlmdhf2BOU60HsD+qyT9Su03bV6woqA+LrlapJ8j1y
J6xItUgpUl4O2RnS/TgZiQFGemX6BKYMW7zYxCvMq8kEPdISIYlc7R4or5Mw
fvA0vQNj59dRifOT4uoZp47DIu3vYT56UwcqXFCNovARk1gcQPTsrJlpLCR0
6BT0KWeHvNBZR3Uu/LNSd0+p3O8LihVnDNVLp7i6ZIpbcvocTsWbb2k/qWWS
HlIYppCI5Y7kYln9puU0r5A5WxlhhN9bA4NYeBXcCeog1G2UHvFZWv7p+ENQ
qHAaCHUKB0wPNy98yb7efkR8CtflDJ+m6GZUj6KhHcCJu6kIBedLA2H9Vmvz
2/u3wE4B6xhg2Q833Bgg1JhOaDQP9Z1ULSmZT88mBy2mbBo/pOOoPRjkKsoG
MUfPBcwpdMrv/NqG6yD68Qm7h02y6w4tVhiWwddUzkm/2r6MNgK4gXp6nW8q
ULXWLx9+YH3V+dJJf0nuDFG+61M/CyRbm2vpNvPhiK+xJ1wS6ubxoUc2gSGS
wCrPCIYIVnwo74w/eMBPn5+RAdRc6Zrn9L0TLUG0RwP+OItc1dpQiENlDO9t
hcNxGo4GhYMAocLdBa/hPabc80jn6iNl8qjWGZM5qQ5RY3W8cX+EpPD55DDE
1tDxCiKfMNMHw3twkmb1oCiTqlZfzNkgde8SckLK4+DyzUcFjWN1x+5whnWG
dUJtFHp9nrlfChP7vPB09Gp5OVx1Zgj0+qphUgxgbyoOquL72XG+8YAn1BHC
xV6194c2cn94fpHY7sGuPe0BN0NHL3Gi9Qjw5hfBjbTiWovATSjoHewcX0r/
NqQgRK5v3KZOVObOxTJKzZG0EyGJfhgcRC58C7NW8KovfOB805wga8nebX0b
cChgQ5DEU1kMUReex0seMLH0ZjT62SwpN7zzvYJ9yD2DXakZRWNf2y01ll4p
KXJtAYzM8QOiNSvUSmj9h9ECb8FGe/XqfCi1bUqAsR55KP2nKPZa6LFyu8Ig
b8cQHK8g+2ysOVlx3xSQXgMJtMMT1CYCsf7Ahq64PhB8cUGw7FY4exIHTQaL
bgmnkLX9HvQU6tmy6FHz/nYTpGoV0g1qXgcfjZE48KxTIZsXVHG1nF5c7PHX
7yq/eAKbAJzzEsvaDyGrlElYhQDe/5xQIzKnjTMhA1kaQVWS0L/EC7psxbpG
QW9pmsLFVfWPdBP1SWAvJlfKr+AS+dIp36cckqG8PFqN3fx33QV/GU5pXDcc
GX4CWlS7VwMwGtJgf/6R2T0bg41KUMSVaKiiVwvCGwM2LQ0wv1pY2VKwsiK/
Sp/3EsCPDJOsJW0pwUCTEj9vT3E4EW8axyq76NPHZf/Zbsf6VRTLHPkg/Hz5
PQ9UL6BTiMX5n6GZHmWE6c/4AMrieDAf1RSAYvTiwAlp4pCwhHQi1oQq2Kns
sj70cVQBHtH8Rx1+PsGG61osp3yxvJKJlIIt71ohERUmqgYt7UnUzSn0jMq8
VXblavY9HUV2OOCYPKb7IBv7t98TP+aJfqSq7QA+D+hvt7ZUVZ5BfiKRbVlw
7rbIBvnmI5qmz1REHym4QuAWKcJlg/+1lKoTwcJcZzGEfO3ICXN96k7stQ+G
esOFh8CvEfR/j9yCB90Xk3ZGWia+mqmhEJWr3phW5+ksLQ23kUMElAucePkd
Go7Ot2ULiYrclShN/LZLvkw9Zt/qFPH3EKVrhwFDl0OT/l4UdVpn6D8zDxIk
wvr/DdzhU18Ag+wOhWARTV/wJD+TqoBZcB0TmGdIWy1fXamJVe0EckBVFREn
CU6OXGq5zJsrmEyAtqE8JarKZS4RMb0EB2doVSwA/xSuLN/R9H+9e/wMdn/B
B07aj/5j6cK/2bG+vijoSsUnzTE8974o6nAMQ4L4pKZrOieJ+dxMKSiiqZ1m
eeLIuV9yr0MKoN88GxnbSIM+0oyRT7UMbtmIF1UvdCqehYNnNpmAruaW8FJN
CkeppkhprhUx1g/mvpky0NRHgLwucYs7BQE2Wf6G+7+Yv2LrUJK7SCDmK+7I
dl/Zu7VkWvttip5+uwFQNCRqtRxH1Zb4fsQ/8Ptl4GATcaXPAtm7Y8EfND5W
n2aeiNP74w5a8RiYn418xZYztDBG2LRsOMDIQz3BGfAwr3iieiaV3NHufO7u
9aHd9ddkcfSpHnGyjFMGWPyGkIzja0lA8FM5y8HoBUnRfWIj5xncPVa5lvIN
Cv3FY+B/ueSzSPVMkKMwK6B4JC2WC2FGeJ84u+zzXGc9icPJ1tCRKMsRBf+X
4XLBxdtwfKb9bSjrz8oBO59Mgta6DgKpzxSflYL3UnVag5ozUoDBr67uGo5j
SxmdpP/F0/tuN2yP9Hdl45ZAVJj5CBCE6OPCeVyfsVBQOei7F1I6u8/gPKPI
mCRHdY8Tteri6e4uZr5PVeBCC5s7qzXJ+8ZEs35gf+fTEe1Zepi7wdxoquMQ
CRXtFscoFF1FXBIyI7Hg8/wxXx72lP8LghUy1WKKbcHYYdIbYwmUhA9fz4p8
bP9pF8rHMbFev+gIakSSsb/Ki210bK0hYG9oj+4lYcU8xq7ge+seZJg1jxbd
b7qT/3u3eoDCHIkpa/GaQLjgbRA8ZLfpLMZFDWYRhFN+ibYFXorh7454UqGu
4ZRyc3BnQT1PuLDGBB+DiASq0WnFPOm0pKu9ZY2p8UC9FV2xgo2Jk82Jm5Cy
C9fRWSp5ZT/4mAp5YGn2AljFEa3J+Ezb0jsTc6FcFEwbblYtCi41Lynp9ltz
F4/v3DuPlAZ5l5uTAdpsMySqNxFXOBuwc3aF/SjyMaj8/IJ6sasxyBbg2M7+
QWZVhXLkChl9Cc+JRwLJX4KQz9tjIJvIs9z1IZNDHRwcaQYF+G+PS8qjsEZm
AymVIUn6Y71rBe3yVVH6FFjCZUrMUyve20ZeIaEyZaIIkk2t75L5510wh78Z
oBpM5Mm/r1zAGReQ24wz9H1YJkAXsLheUiM3nL6rClY87IucUJxmTrRx6Lw+
8J3Jn3cfWGkE95GiOLmI1vlNMygUFYIZRvOOgVq3ST1tr6y7obgN1ZiQNJJm
ppfkwSPkGNN+3ycMF17RFBMDOUNAo90nA6mB3CnzjPhwCwjSEMyA22z85hpd
TATAQeahs663WP0C5XbSKrJ5firajsmsmnU7tDqyVXpDo21hKiNhzknC0E9H
uSYQPsKfG40g3Nn3wjAH+idw5ePSTkxczORZNcNgLRC78nJAZQlgWctkFG9E
yYjh6w7JK7otGiGlP7WjP6pW7KZsSQP3gDRJuiUmkt5TkXNVsXtcsW9gz1M9
jaKfoco3VRV3lPd+bwqxKBCJIQBowKSF7JMyvcUlFrFovdldf8mhvevcmFWl
soHlXX4YTD9iLZFyeBgSaayDLPQjhTQ4sAZU1/3kBfGF+dBPIbqsNFNaFgt7
4cfvWQF2LXP7HyzvNBavYjQ3sY+eHkgAMCS+HbP13Y4WxmKnhZ8KWgLSo3GA
QcO7sFeDuCwgWe6v4mirqujE3yhgQTNq5QVJWMfj30BAZ6mTmE9APumxJ5Mb
JBfOipsElhLysxqkqE/0i2kNVkvOqfMGUf4MC/ZAdleVnF+i6aKJ/AzHcbyf
X2ldMuh2a8LTOOh+G23BiyuNGhdxvuoGRbE6XleGxMb+WXFH2FwT8ipMoSgr
XPbcytbM10fcI001NoFpDOP02usRUl464RNcfFndWZgwLKLuoA2vTyuwoy95
WJoQgk8Ovh6gii+nCcwqLtgE0RTNMJ0iA4Wx8NY4kFo5W2w6xqO4RzDmUkDE
cKseGu4rIByfj/8m7PEkilEKMwZDHY5tIqc+LmSH5h+B2dmTYyEr7MLaufle
IWEtb16CbRpVMzxVnqBdyD0vHOLMMUHnKcMuCivTU5gzrXRTbSmRHLYLh3yT
cgH1K4dsguw7kQTNlJvPTC3kmNlrX7vJzT5S9/hPYz86vg0RkijzYhjZ6QmT
WTpvG/ZCfW3u/2C7NQSIU/p7Mr0X2//78iha0pzOiatq6FIOvWY6hvS3diNa
ySilbYaYbrCN3g2+GIlTlcxjndeYCr4WIFhxvL8Y/uDj/oPE+9DqRUJSg9IG
vlED7KJx99vm/cCNjXa5MK1KfeqB1CHOSjeFL/2Z9lg6JwqOv4RZUbqvm7Co
k4jGA6sfaxbMKv0EPYjhfBYGzE1alndL3GlTB8T0xPOuunReAe0biSpMYAaT
lYH03KHMggBX3sfJ0RUAUMr1/nhpFUaMy36uDeK7R8shGJrE7M8rbAcgnh3W
/IB6WjWqnicpTAcNOEvhAAX3HvRy2x6D0fVCTkxtvplOJNfuj3YRVBzKvhmS
1xjbPA87KdEco4StEGLVK7trMuubxqPA9tLD5IhnpP5w/vhxc/95ci+IZsZJ
28q1gvf0lDc9UQTg/7Ult+0CCucH9NaUG/2jiI3H5X/8C+V80Vafh2N3QG0o
bSs+JllNlO1xCgrLokaHzAbXuTSeyZaC16Kn2bxCizWY3bTWSzrzQmEwlNtP
7aSi9OJ1Gh4/u834LA3lum9YqhujQy7PTCGKEw8rl60Uguyp9/7fkPxaS1+0
MD7ghHBp4O3YZ65iFVslOSlyBZ4M2uHEUlFwBU955e6bCUIOqDeuMVEPeaR9
u9iQJ7prlQgqIpZ2lQd4Gl82DktEDSPpx5Ibe65IeumP9JByR96LKJwEpJ0j
hPMnL3hufGeqtcIvWTFof2bjNt7fozXemmmzlnwq6nAGpPTONyGGQXPMFEL3
GqAp6jlcblmefv6mJnrHqhwUvTlCwR8OYQz0dS5VXSRUtLCJB0sNVX044wux
Ad5TelNvkPVkx0M79vhmSnXrMjuSrycUPDwLOES1nmAonqqPHYtkw1umBYNf
STX1pWPDmy65Vq/Vy6ABonTxb4tNfb+XZk7gyYZ6cCOKnY/SO/s8iz/ussfH
1s5ctpwP3FhiPGdlw0JuT7CCqSvaf7VeMuYs9nJootFSa+fULcIUFvUNx9yj
KHkMzAb6C0tqtpfONwflkZCvjBk9yf84rTVkRQDs7mhhHaw3y3YhG3waOoSu
uGzXKBkZj0Qh3DR2BsmdSEeQdHwjn9f7T0deGCoDsHqksYJlqxcKQvX+BwmL
LpU+00SbCI8MaH6fY7a6OFp27HJNIsMQjf/ii/AdZt2gi66F9DylubmP1xLd
r7RAQE7arlPmDFwDWb8ZXyflMHFtYYhp1CEYf4Nux2RiD6pbn88YHtkjhm0R
qx4vfnKQ5LM7JXIApuoJJys4iW/dJ63QDQFYBs6pGhhOVRHHAo8jSA/Q2LDA
NqkV2xozdxHOk7jNT0boaXxbgF0vvCG1W8eyPyUsd/cvDm515WYzWTewYQPF
gHbpCyyiNWRbQ4SzI03LNJlP2AdNzcToGCyPBNz+XUHt3ekp1upu9KR8Skxs
6Hw/lth+rO6DMO7I4BFl1hcg0xVtemqSpc0oZlmbq8aewejILzMTcLYLE1EL
5wLCQodoSdnK8eWZLR13ItA5JktYj4PCpTykIvj9iu7iow3rkqS9H0TwHv2i
jq+Va5Ks4slHeBrzVP1e9HFWdYal5MziLjqYC9Tr2QJyuPv01DIWaNspf861
hsgNIRoFCaUjBKFqh1m4OHVW22jUAcGNjUML4FFvxf5QMTq3fJZdXbEyxWnC
HdD8OiR1jOh/NzQQCvMZI7gjR7g7VeBvmNr5HX7+DMIoA5WJf197OLiDZLb2
5p59CCmGETAHhyhrR/Y5HPqwSBHjGl16qDFn/AAtgZVkEmL2nNRebf2rmV44
ihXv7Igo1I1fpezEtNuManb/abi0MCQcWOgwNMjpoPimPdv4mCC8/unQiI50
otIShpwShnLFn4tvUBi51CVTrv/MQca3O5P8fo2B0aAjqu6/VVVxOCrUrPfu
OykM+f3tBK522Pln/EfmXec6W8Sx+soFD3lRYftrbzPUU7TSc0OK8Xv1OOH2
XMBZlVCI9uGNQNqpUsCdp3VCXJzmz6pkyv8Ayh8Xxx4np28vB74vWvPM8bNx
ylRWulvtdyZFJSmKoxFUgUDr/i7qchfhkkltzx8TwZEDcA0CdlZ4ZbBfPNho
HT9Jsxtv/mzBcEp0+9NeFyETtkF5CJugweTSAnFqHnzA3NxovyNoutupA+Wp
C98W1Wa30YlgVfkMKLp0O1UEE/K7sgkUanby9X9HRL7fSCKIzVP/Anj/W45a
l/NJGhOluT5mGyiKn77UB12x6DzIDY2/heDG/Iufa8fTujwELSv7BsN8ti85
wEMkQiBoVhEUjxaQtGUD4b/4ugrJtwLnsjZFSbqDIXf6+VrBhe6uvgZDHttJ
GkfAO6d7M6PlgPrCOOV0x/bBOy9vRzF79GcVx+l09N3w8sZotAP5CwWGVMc9
jt8RAooICgv+wLv/Z5++9tAccTGxyDhsBTUpA/cfLS7iEkHUHA1eq+Lzek+z
287iy/wIdkOAhDTN70eiwrQ/UvfDGuNF15Trd0RDN5b0E9OTHl6aB8psqIB4
qPmSVS/5kEfu9y2hCF943dxb1V7hbPZQH3whuMHWr8BJKLTpKOmcZgV9V04i
hcs8XEwhVRAPBj4QswVBDZQU7I9+AVHyDBc1XLbDdi538ziWK/kiYR9saRQd
I3AH1pGTp/Hsyd899U2cORBDb6W3e0fNU2iTebciVte+GMo4N5rJ18kca3YK
WA0r4MLCozD0Fh6gtaoBmBf7x0E8D5hbad6mrsKDOU+JbYN3htgie3r0pAni
JFVHrAg1oGWiZ1dItNz440AbSzy+oUBjz2SU8Yv1Fbwm3PXS3YD9ZPhsTwyT
N9MnofjXr6E5WYcrBHEWRKwWoOV8jpQ3HiVbpPXUyPAvCtHdVePJBIyouy7J
EjwKS5ROVY9dQgSW35WVTenTnysZFi+0/DtNn0H00VkuFXeyJQP/ViRrdieB
QQDrVG2uWFZpZhML90sR3tpCvBfc0klIuv037kJltbXlfh6ko2jzxxvdKciI
ZFi7UIlQ3gAyivKs42nFiDL9+jRX4B2P3n+Xv2gXQXT/zp5mFxYrHsL/H2d2
4QBEMs9uPwg2gcqjlH7Y9zH7XQUFpIh7j5DDsMwTsSuvoVo6i+5abovmyV1H
fCcdO/1NI0VQwPJX+LHRxHliq8t10qt7TfiH5dvLmTOmnZuSxJjNkLXFUCea
qamzojXE9u/cjWYyF4i6ClMI2JPiGznm5svdL7FRzPX5XltAv/YDUw03HbGY
Xx6paeB7Dg6HtYvzIKKOoxSl2sd+7OfQ5bWO6j9YclOzSlDXBQaOK9aqYVDM
1orhgQp2yg9VCYwcMIKKT1mV95QUvbOPPoXwpkw3CISMx9ziES0meZrv4l+c
aTUd1fGAkGvF2E/pPKMqe9ABH88T17opMZK444ooyfrCdnAL5guwnBKbsAbH
5jGLWHZjBrsMQ8wVhTxqd+ekJ61KdZs9uqZYofvAhJaX9eTkv7qmlI+sZyRG
gfdLwZUWpsWmU2bq6ILz7RvV1Xn0odE5P2DRVeXNvSht9RuNe8/m/M8isXP/
Mto3ZkJOW3itPFdm7drQJ9OounvUpyJ/5bqee+qEAkEgCwpSGxlMDVmBZbjS
VHZoQ9j6P/32LWAHrfPk13Yq4vGXJPFu/qzL7Hr++h/E3GElGbqnZ4+OxQqs
XQ80rSSHBo4AsxfS5zOyNYg7oCHaoUAzkBCD+rrNnDIld+7oT3NgVXUwXpSz
k8qPMG8e8fEwPcLMLUvsXmgUwWNBg/vSEprz3O8N1QAc3bgAzY8eWw310pDf
UfL/qy3lPhnHTbFSoUOOK9xCJTLLir/FhtoQpP4itftJUkpEEDlCxw5YIFkd
Bti/jvRIlnmPQUu3N7lvWfMp2YCUo+HzEj7KSc6BXi3PX+CHPSkABf29lAf6
x/f4hazSly8NWfXouE7s+S+vOfWaBa3kf7XSgUCPLxSM5ejVYmc/L7lwBdHD
XJ6/spkrfpliIecydLixpOk38WVCG7PaZcDiMV/cjL4vsDS/D7s4LWULEg2h
/Vvih1euFuXrTv21dr8C+qtg01SDHUyTNR2MnxhPo+AgFdnMbjxAeMvxGtHj
5aiMfdbI00wi8B8cOgXebzMSA52Uxw81jdklsFKtUqS/MMK/JgA6/OtqwUoi
6Ar/RVhrtfgDnQsI3YaB0wEY5LeGfpgYoURSGO+nQTehMDuZ18Km/+iynvmA
U6eQssPuiJC5QKHp4bwE9j8tWUcu2Tw880+IIowu0D1jPp3IUAWF2e0xuJem
Q2ZTOglLc9A3KkypeZ8IOg8xMsv6AzFB5Vj+WcjOT1kU3TQAL+yuJcJeAkfD
/xKYb2LREBmmL2Sz5CxJDzd4kVQ3JbAnvIwA7dMYUUuc/E+/Ja+Ihi6HJqsA
9l3pPcYbdSBMoGV/2F2HNYBlQv1eJA6HsLbnIYsbcNnsfLX7/xwxpTUzIFYK
Sk6zqCuTNxNVZrLtUyLoCrRjtkvOqhL4iuHDU5bB3TI1H+To1s5z2Az62XdN
45dAsMyKymTCr6FQz+CGayxyySP28EzEDpQMI7v9mZJltrqSaT/2Y/pkUJ54
2Iam/LhWn5FaTvHq2tHrVR/trR9x6UpZ74wKLFX+Xry/eGYWUWcM3WRgenjl
O/H0KeGVzHyB8ev6AWXBVdldZmA0BGy9dQHRUZ8qgTz+CtqWS2jL7aoxcBTj
bOvoJy5a1Wzw/1h19ZssF4Wh6uhnWkM3N87HY+yuFhwFUPmjGhlHZLecjaPL
Iw3T8l41xYQFTK3urRjcd0fsRJPb9+P6COXhWG8FYZWcKMuEFfpfmFz4OlNQ
qZ8KyWcVBspcX2txl+0CN1libkDhJqdFj2yAtX4JRSVEb4UKH5Lc8R5b4qgi
C1SJjA10AxlhE8/IjKWNLXQRqLitiinMgh7mavgghkLfBSKxcDftHV2H9ADL
v1O6i/xP9LXa17jebT9x9n6BA8v6AqHc7TeKkP9quUnd+ztqHcAM6v6AdNIg
MOivHD8BgxBGTM9qtLIoZ0SsREf0HY9pGY2aD2QyWgvYBnalIxrtRBoQd1zi
0Yv+qdpnB3nHwwg0BST0OqnbNQ9nKVm3hUz/XP14k7ovJvZO4jShQyirK6HH
a07ad5TDyc1hjTmdbECtzyaJF5Ul63BF/UurU/7emtMj5gGRDNxKxyXXBzgk
v/5DEFo7Bi6Lr70MuTLZqRyJjcEOmlfMXrzwL9hprYTwut+sf5+UOThd0gPK
mmOzpbK+2IccVpJTE3RfLzmCeMxZ3PGUMnzv1QZjKWjZsUigfgA6v6KSBNiu
ratbIqmzWxsSJPNpcYkAq7ju0Xx2irZaFafqwnrXh/A8YluJuxih3+2/OSTq
od3YTV+u0h80Nt5NFSv+3KcY/zKkxMgzos+QcAQ8XmmAnN0RXOOW8/6w04ql
9FhdrtzvOC5YiujZQOxBZ9c7scfIhZU1vpz3dpACe9tBhrtRftj6Z2ztVBbq
SB8fgwpPex0d+hhhJk2tNGAEn0pvCSuWp+5aoGPzfW/Y6ZtMTRJ09sET9Frp
j/acrosZXhmSoR1YAbs5eSueNwfC4oLFFmrgYBy79g/mvKSnlUcQjZTkK3yo
HG0651M4FQyZCzKIfK1QrpY5dFXLsVR0V70P/WGRIf9XgzdmXaNkiuJgepzh
bU20kReKw2O7tbrZe99VM6IaBQg9Zp2G2pIreKV3x27JjNknBBCL/8ZC0Dwa
576BxFPykSYKsFNNvv8QQdSSqu0/nBu4rO3POkL7s4+yOrwI+yIlQuSLwXJc
/ATjzOKx3p7KorabgZUcgANqDt0xprZyEekoEU0/ohIGzhZ+XCyPqiOHChKt
evDfJ8NLI5gg6uFiwqL1MSEBVODpwstgGWM4Q16fTMNwZkq1uG5uwkIC+FEW
MRaMVHr75ehWCQn4afT/NqMmsC2bi8f/XD9KNMUT2k8Zkww0750ErtsU+yh8
pdCZ41vOR1rD33bm+iu/k7HnafsFW3i71QKcweWUQt3VWZHYRuARv5dlqLXR
0LAIu43uZZUMyqO3XdiCpjz2t6e7dMmHwOjAEGnWS7nqRhM5Yl6w98Rav/+g
Q97OoFmJ8TQC1cd+wzEZ129bL3aFtXygQ2Y1XzI5OD2ExD4wx5+9CWte8lF0
0797D1CeVtxrFdtfopTOjnqnZ/pBfXLxzMLKnNu2AcpaKvBp1CYuRKZPI8UB
zBsgXChKxjTQP9h2GPg8Oqm5aMA0xhWD1BGsIdJZHRJ2UpC+9vDHfW8ptCKz
41sEmTscLYEkwVfhUGLERjdN4LV/jX2YuYxiHnAaQQ1o/IRC+aSxayNw2VIY
m/mTQrryNQch/8rvnxWTrZrqIs3eankJ/5louboBL1Nng2+sTPxJp55qrVzL
h7EoMk1FvsBPiN91YdR9yCx7H8zX2h4BwGFxfSO6sZ8pw7lHWWsQF7O7d0L1
ym4L9hJaoqsEoDLoZnFCzPYF5CjJEwOpEYfpJDJHFKDVP+qMR9ls63Tjq7i1
GwW6m2FKppx+os2BawBWBPITULAJPelNY5Tsr70ji5RORKij/mKUEPBGMJwF
+T3fIMj9nAjfXVNfdzwwCNRmHMVUnMbWyQCK5b9WlP1juYxU3yjE6f15lSE9
UyU37YV3cE0kJq9biM6Gm1M/RvEwQcgJJAW9XE4464ZNeM7CcQboESwh3gJn
E5wQ61q2bw/GdkSbTUPm4QXOFJ0C6zHx+XvALhiD/toVy87lFG+oF9jBObDh
MSU0FhDc2O/HA9VYkCvM6kCiEAhA6bdECllFI3XUb0FAWNrsGWPu2d7wMPSM
d7iEw/MkpG8lzbfZPWWY8/SE15Anb9xedLvLDeVHhA4AWZ0cwXkHQN2eidJ9
SjP8v+LbkhlZy0znZ1tF0Ll2mRe8sTleQC8QTBr7osgjr5luY85iki6PMwyF
TFrVceTJm1uidnxTwe83jDMgYlfjw2VxOYDMKQalmIld7nzpKF9G5lLFvN8n
ZPKJmJiBYcnNWrgTNO9DNRi7fJPV8zyV003vr19iN5GD4CShrJ1gR1Bs2/D6
y8ZBAo8DXN38qQbIf3IN4aTylg38eJjuprxRKc/GIVekD5Qiiq6VaAv1MGD4
y611/uMfuiRl3wv+os3YkwhxCyeKqYRgAopXPI4yBKOSvfzGoxaFvC1slvCs
e6DUoyowpFB0Mt1y1++Qh6bDJmRg0Z8SjIxYrHLoAmX5/NAPoSE9Kv3hH1bu
TcBhGjz5l6pZyOBSdlQVNfjQqMBGyE4865mg8zlb/5N+z8rFLr9boSb4DNwT
Tn87+jJPFob6gSYdB/UCv0ykmIBNH7yFXco4Birdl83la/v3hgzA9mptmjJL
XoiTS2CkGRK6ObbQ4gOdw+JXe+OEwnFRBGOj6B5Lg2UD7Wp1U6n6r064G1u+
Or5wojdZJByddlAqq7GcOCMBVcPAtDlSPZorsPdwWMCOM4xP9bILADF4BqNZ
1WOta3wQwRs8OEf5gxscVc1Ox9walPzCHYjRmSxrKdINbc79MZ3RfCU+ldc9
RZw03G0g3TtzNZLAFnrFNqyCNrpQGJ1vS50u2R7ns5M7Z5yAP6JT6A3AtzP+
8uQqVtcyXT30FVqyJILWZGHNAC6ZQMJczRIhwxqUiKBKJvm/4SxySrLVHRR4
8sl7ELjQqrkOwLT8sLy3tPdsVSid+3WLqDzsC7mrFWV2ZBVUnvnjY8Y07e65
e2/6Ht9lNpXLz5wuCkxX7sOZWbKWGFvTjzqcNywMu8S6jsAAcb/hJIUhoOT4
PDmuRDuKrXUAY7KqcQCKCMYMglFX2PfLy/DoJauVFVb4vjjexo9MFkvkGTP+
/Cqb6DbwD4Qeux2KjkYEhFk7M/2vdJaWDXKzlA2ELd0JuGD2C/6QEWVdJ4Gp
cGbyUPEv0X0Ei6EPR42c6r2wEuewJix1OFpl0+2SRhC/o8tcwHvS4z4e+Shu
7jT3vPVQYQxeq4ihc4gwxzXUeaEPCQ7HDounKGuM3jbo9eXVVEKmADAD9qeP
6/8sLqh7Ht5DNWZTQY6oRr9kaqtOrZZvJrhhqaVIcQQygotXrSsIxVu/S9Bh
4Ay7/73XaGy1iIBavJJYkA7FoC7sZlDGQ64xdbpqgKjOsPL4nO+c5cUiKhZW
lifwBlM/XMB9pT2TGSLhyY2gOxQ3WFylj7Y+797EG/PeNU1E1qpLat1rINAS
B4jQiE1Z89GoFvODAy2hyrU1ykJvk0sYcfN1GpPtEofWp+w3GkDDRZ8eAq8H
qVvV909C9idqUDfZjL9ZaMmkox/SDXb2DtxDo0QQ+MlASwD6iP7Q7/ccbpgb
sgQ6tQsi2ygZIrUS76sJSJXO0vMB5KxoD4DovNQwJSmupB9h3Bh4umKoXqFf
W43J2F6/f7d9Vw6g/qVwjmdJG0NkyQa7NsybT8otI5fWObMEl6v8MM/DxXVw
F4L7XgiOp9RGc9PO6iNMBDfpCfmdCqCVBG0NtMkoBxDItO5b0wr2+3OSkcfr
Z/4hFTmhRNLjVbCl1B4jd4Mpf2lYp7a/SjiBXliAAENq4JaAgSNwzlq9B2/9
Iv8SbQDG+VV5m38HpZSL8C0oKKDneBczhwY6UBo4mlpjTtdQw/ZbxS7k9VsL
xtWO46qtL51CJMc+I8IWrKivWzMY2Bc9i12SKkguIPdBvYT566BTnHDrcMD2
AEHOLV1tsErZZNHamBTtUGTgdHpRAjwVnS+oaLfPJaAsH+/qLW4R0ZvMnz4f
adAl7wzQU7LwtXSnwxm056K25OEObxGxDS8LVgSO+zcA4OmydQC9Na+PxYIE
SIPqJriISJGsM0WS1FLwqSCWgcGpbUFPvs+85WFl0YZno+5YmJ2/a1SiyD9q
Ry4XRc5k1z8UbkHJ/yGdA3xG0Re6/7cnntX0y2SWlJK2uFSwuhybp20hXCY0
U80SWCBnykS2dedzILSf5ohIa8lULU2iFmwcTb2m+ESb+fWQukoNOZtnZLFT
1qHOCnZLcA0g/5urYQlpOJVwZrNysiMCR1d+Yvmxxjaus6+CXcifLeTSqIla
+D5UHBgC+PGb5FevjP56VZferG+c+iLIQmmfUJI2HMGfhmORjmx3cKqbeIF0
1IFMQUP6GK0kCD+uyrqwDrbCxoncK//PFOlx4nYRhMKajGHQB7MExBNXCjXd
MXbPqrN8+n8DXOMMhuKdXqlX/gNPkp2BdOhETIFRbEi+baPByJm0am4hv3kE
mWqJ0lVzU2qQcn91svGlNLU9DCNTSXEqZzF2OqWG2ZHFuExFyiL8ktsYyLv1
Cfqp+xbbl1b1tueT1ODuwJuYydJTgF3Hf0KOQYIiN0oXxSQa2HRZiAB2S1mf
/JBy1tMg9SldUVPDMQWqC3ShqeeuAQGEKJEYWyFuuXNDRAh101OwAGL3r3+c
GHWx31tyPKkikBDn71HM8ASbJKCS6qsMPTvk/uuE2H4M83IgoVBawM4ynX6h
ohR9nB11qigKGEEmxa3N8hNgRh+3523nUzkvdzIXBLlSvwT89aY6VqWo/cnh
ajU7jfMEz/igslxpGzgBEMHYmPlAZ+IFY7WoEVqN5QdgqkwcgDRCdCGsI65Z
0VGitmNpIE+nosEfdtkq4uT0fuv5ogefCzR8eWl1JeXoaMMZxEpQRhBc2RNb
3RivYRG0WCCmxBpK/nOtN8s9qn+ihpi5QFAprO2DmPpGc5i494+zS00rscPy
z7v+fjemru8OceR7wC74FnFcBb95Tw0W3MlP75oRwuRzRB+MTi3lMQnNdbGf
sw8F8WuwJEUO/Cff5AyC/ouylfyX0WOKZBHKwu7n9oxxT1IesRxtZUfQuyy6
iahxnQXZRIEAZcBARu0E3Fs20sRHgpJin9vkNc14L5CTLIYMx6CczqCh9pM1
9NejRhCLP14IxJ1KlAJIsiClVcBU1wkgdDWEv2NLHUc2GvajGIixv6hraCO+
/Qq6A5hvxQ1V3JUFfhQxy7uybC5GjOEKyU43WOnjWs60B1IgMk+SViAhMfQ7
/hwxVLASfEpE1cphIXFPeT828Bv0qzm1YMMCjsrt8c7pqcAeGTkz+WvUsk0N
R0wsFxKlCGVNg4eFXFPdIkLZa/c9I/WzC73CiZNVb7LWYGsMjreEz8JWiHuD
f+36PH+aMFmJfnaOygGK90gjY4HYSQ7oJUxx0TTif7J0v+KqEPmIyelojQX6
/uooWT96MaOchpYUgvxcqj0usMCjk3FA7bIqraNrvxru/b3s4osM/ysIvejM
pf7ysjrNXVzEgDAlX4qQ/3u/g93y8haP/Fv91SIbHJ4ga4gQShTEPYvXYPFz
5pHdQN3TwHPgbLqDXMnoJUrjg9WzexmcrHbBTmBaAY2HZNnCCcb2+gAv+8bd
NN1uug/Rbnm8cL9NNrHl65FIPbtQb8Vueb35+s2MV2I5+Cw0ioKApfDG4LVl
LQZMr7GhckyzPadVbkFtjYfm1/V++61WUlqXA8hCszRf+GOUyEOdL7qjDEXt
p5YcbN35L3WcNke5zOjDlfMvreTG/0XllS+78LlkXeIGb/usSWaYKsuNtw+5
/C4svVkmINKc+TCTnHWLc2YPBwDF0fVYsdajeH/q2lv9zevyzW5n7gTiCUTT
a8fjhzkBcmQwrDUKllN5yjdCHeewXjoXUpDB1iUg2MZVc6i9Mp7OcKo7o/Vb
cKC60dg3qGLJXjS/3K5rVwa70es1DZPHoaOlYye1f8vngp8D7tICAzePLfN4
fej5IAI9LCT/1hny9QuYV4+BqRQscaNu+b41OvRYz46YJFfQvyT8Oa9tVlOw
p74dCPOl7M5tORZ++yKxEBTBGY/8qCuPd5U4NTZ41xfa3t1k46sE24WSipwo
nRfmA+RkTpyDdWpi2FmiXa9ljjdD5xOpkBB8vXkL/F5m9EsTqMpPd4ZqJF76
TMagUD3Pbl08Pr2rJQSQQhsBZmyDUuWQtWoSnjm4KaIqOGvi/FYwt/FvgcXz
9w+M7mNyFgnXQPyRuk8SQzTNzvfDSQ1xqmm20ClqqR2TinI+ZqrN/0rNzic4
ui6gFNyzMLq9nAxHMneGU/WeEufeZzpdC2p8LgNkjRxAQBbnLQeculH34o0c
bSxlo8l3t8VPsuVroePnV1XmvxYJjhgoY0oh1JyBrVAwoOUXkglvfSFjXvcM
9oyKihz5+zfizPT1p42RyR3FzBN2CnCba7IstQ2v0BqulJxOmeQ/deDZ1/W7
/5LbqrHacpN4hcOzMCgeSmzuPEYLRiFbw/iFbKs4BkPnSK1LJIIZgaOOsweC
1Q2/5WlbkC76wAhpt54YyrGdZOu03Me0Wu5d5MYgVS0uy4XmihqWPZkJuHdg
p3Po5h8wNvrFCAs/4M8QyPeYYbq5lLR1+H9VOaELPqqazo7r0q7akT9DlS5w
Kp21kp7KMlYIivHnWPINdVLwB92ymiBJQ7Gjr55gLUePrVDtzqlA0kQAH8Kx
slPLLwmxtdeXvREdAvheVsN9XadblIw0pv18ufnUAZtts+eGRtDYvsUPcmoK
K2vJi/bqVoQz1Mpr47plePBExhqj6/Sx5Ye7p3G+YCKpalTbAuhOKKzn4G0r
VGVUL8QuEUC6b6dDdx0eTjfDeffldGiU6HetYcaHCFkStHeAWtGOqhtUA21B
yHuX/QtjybZb2/fecbnoD3lDYDUC1gfTmuXXEf2SU1XWCQMd71zSwoIf7m2Y
zx8h5+5QlrXnoK3pPuutVuQZMmVcLbxfYVRIrN4x6FUR+/SdJMFK9JCyTui8
TVE28gbcdB/NvLoTiFVqrUaRpIVl/Xif8MKpScJ7F2XgsHHksM+I7Wt+Xbwq
Q3rSXUCk6xzaln6RdhZJcm7DJb1PRyDufHIl++viImFaVnmYC2cw79BDaJTX
gAU5Ecr8nJ8W5S+SxtkHhFhDHXmj0AVQ2ftqb5NSDdEMyhWKIVZJ2CkBOqA2
JYCCgxi3TD59nxHIfBF1ZABG/c7T+VwnoSuUcUTF/wEFOMLX0iMCQlXvHpN9
qJO2OuGwxH4or/w59TbO2UXA5PkwBSniWbBXGHxtFbITJTIIzbh98xKpvad9
cjxffF37E3uPnQhbnREMMYj3nPlb86UNI87y3W6fQ9ZlkcfdCZjLgLGK53Zg
CkaPLO+JeVyeqH0I+SlZJeNGaqZvMd0N74FkBv8JLhiqyIXwnW1SRrhj2jsf
sQgYWdsTdYKh/wpoj2x0vKoel+HRho84zCwoDSlsG7c63Ogz2m+DV3VHzFSo
SKSTxbXD/8Sf2s6IAqdmB76OdZu4Ew1GRDQozwDSY3IbWaITxf9fEbt323XU
nGAJT0CznVX/wiQuhWMi28i0I32/pNgWuX/C/53mLIl8Ib0/AAnuu6xYsD8V
FAkyJPjVPs38rmjXJkljESk6SyBdyg5MryjW9aJGYUgItPWWP8l18wfnu/jv
N7Z8F/c/6PAWWw72vsuiqtD4Smg+b0Mo9wYQwzvrx6jWrNI0hBY/aiDzRSgq
XmaYrYP3+TUkryOe2wBTYonfxx26C9mZwKd/Y4LQDRbc0Dc5cyehxOtjVzCM
8LML9I8sXfU6y3vd1d8BBhjssJvQD1T2Ti90oT/KJIBJFPPXDt2qIdOYsOl/
ojnmyBXDXGmEbDMYWwi16XlqRaGhFE/Caw+6HDcLxXGck/+rHzR6Z+GWVvmt
sfCNARf0/tjbahl+eWO3VRIM5kwu7iF0qt4BoJnUZgWJx/7oxcbfcAs8vQOZ
iphP/GIjSMUEz73vlAOEINcyHZ5rmD2YwzVrjgrfLE2+Q5ykR5mOLmkOBrxi
Cm7Rqv42SV2C2mWOKle+/GJQQPmH7Z1D+qJMXLnHT3gKM0cH2UFEz02jOTZ+
DdjmxKaH8ea2hrBax96YfD9MxoLYqjbrzTQehhIp4yEBOWXUVpWh6e5Y7m4v
NwE0FWYlJviBOXdLk6jz+AKlbUN5KSxckDWqQTIKnyYW+uZQlQ6oPTlrW2dD
oiJAtR6xAAXlO46dtT3LtyQU/ErUiYnpit7gVJcUBrk3im3rmmdhp9HDgZJk
YyYo+u5lCglSnmo8PaXUzQL4/gulFXnuRH8Bz+0pnHfKIJkskQjwm9ZMMI0s
FEKLJRDHhNXsW84UokC2XJ43DmFTCduOe3WeA3goMM4VRk1XYRN0+Ulb4wHJ
kHh1g6Gc6oOslg6ER4uvzM+my4QCS0rPQuF2Iv1GbNpryhij5wIMqnG+7u3O
kh4M/q5iuQS0u9Dr+IMsSq8dC0Umv/tVeZiNi2P3iCKqTBsVJm8qzTvV8SGH
MwqbbyJA0RPR2UzNu50BWmxvbP9PzXUQPwRyJfDeyyBDqUo05cBYK7gD0jNf
c3NpKzof72kpVk1uNb9hBRmtQO2b+/9C7q8ut1wtGB3NqcJ0GCTmCpaAe6Eh
2k05L5kjMGJao7tC7RssB98wb8pVy3Jk9N+wJwRYe3GQdq91+aVS9/WTKOG5
ZVTNZnLE9+7e3z8inMMPS+SLNNSrCTKHdBw3NfsryxAO6wY8SHQC+X/ljmlt
JwdIYADdRIdeoksNYaj475tOSib/pnjevqlMiZmHCFDMbKO3LIRrGob/KXJW
y+rXHzKm9laEJm7PPfylSsof/VDRV838LhGRU3u8l252C01Va2q+ap7Mh/tn
BJGZteMGrXjDiOoixm3yQXU1kmlYOyfnsPaLsFmvnYAR4k2FFsNc+V6fHrtS
DSmfP4teHJLe+4Ke1eRvBj1m+/Ml/hUKZPofxIcfppjuDPZCqiAR+B0qAs3k
D+ALZMjoxduI3qRo5ZcazABX0Hmq9VyNUxu6IQszcAIFQ0j7qWecSo7L/xJL
0yB1FqJVqPSxjXcCDxWtlR6KACPfOOZqhrmB2kpcfHHwbBV3HiH2NZEK+8Nc
97ac5wQcdIzJ6Dc2xf8wiqAD9R9f6h4BCCPXh4c0uA6wP7X8zv6Xi4QHPouh
aPaSOLup5x3mpsWealwxQ8kaVYSXUwyGjLYmkDDsToBBfwzIsb9RRjGB67zE
rKTN+eQit35+tZjlW+1/LYwtKg0safqSYDK4HGQRZqiDM/yYFCHQ/bSsADiD
kmvZoDxeJ98EsWWun/ZNdDgLNX9lamiysIIBXEn5PoErGj11og3I2HbNuVCf
JPgZqaf+Y5RpFQKxJ9lp6crTUTEgdqBUgzxvwR7B6+HH8MeWRVy09/cy3AXw
4jNrcL0EY1PE/99aFmnDXs2MKSuYSJRy0OJLPUkxJFCmugMDCOLLgMtjjppg
eoDRsgt38SyEAUPmta6Mfz5zP+7gqXV6jqmfcdyEL0oEYuPO6QCPUpMGBV3R
PqcDKOUvuLdzNArz1+xvUyfbPG3Fx782RECSyo4r60CrMI2Pum2GbCxRA3ez
g7aelkSGOxkHfRgjZGgKABypmrzdyA282G8kuaJ+UB3N/5W9bDAvtYXFpXYn
OAEo7ZuMPbTdncDiD86YBn5CK4O+BHN8NXCV2U2+s6Q72RTvVmNDHzQs0c3T
ki21B4Ria8gGKEqhTD6aAc/IANsJ3dSRjwCPUxcrWYyO68MDyX6yE3IgKhOc
cA1waJHI5a6v4k6WpvUB2PONrNF62IriCIVjAjtPpyxQonL5jKgFhPm7FO/A
+v50z9WJPtoQHX/7d49nIF5SuM2DSSWts6vPmw/hGdcK6TZr0Fk1GfWJeqJu
dUnKqsMGrNpv+5tpJwK/TJ4cz7CYKqPWNtvQTXM6d2nopdJ04e735uJZunI5
HZ3G8Q5txC/tnsJjuxvIdKc5KMNuVu1OxiU19ETBtjBpWjOxiuqqjuMf3DJE
aasJ2PCDxDIcGnUAWnEDVXnUnH1t2J4q8ih0syyevYtA/uAoLll4hrYKM6II
+uwArHEBCHFZtG/UHgibitbugzt7dKWLQgEoxxatIFARN4wSjcWLpDOXfc/H
keb+Ze3z957laiVueetBHr6W/tVt4h4pUlOd3q6aYWOIvuq6NPQSNg4Rs1yt
8Zp6+686vESzNRD6x069ay6JkMeJ0I/h0h+YAy0fZF/1XvUokgy0OVRfpwGT
mVbOTxtCM+XHaU5Gb9M9EYdyQXiaaSoy/zYti6KcqTYIp3axCM5WdRr3gxod
0QSrwuAgYYIx5Q/n8G0PPdbcXej/aDyWo8u1QGUEV/a4KXnLldTppRZveeTe
jGTB023EKnfIatNXUfFdOA7hJAOrq5qP6cF9uf6ifb8oefFteRyq2Ize1rMs
FSvjBzYsRKtjwocVKW5dX0h4bE0DsAkbQNT+NKZgfZkt8TsiFEyzzhXqX4m7
24zrmTjTXyHklOGecsasVb789RCuK71TTTyI0+UNiSPg/WLhYzS3Mk9I8Akr
PKP8f96tcIXyjluoan1+rJF/Kslt99gXr3kWI9USC3SKLA+cooyJKYbQY0fY
KKq7g0LYDV+Pw4nalcf92aYZVSEhI4sWAvHU+9b2Kty55iXByt3KrvZwOeFq
0DHvyUrc3b0vKUpO7UpBkcjMEfbmEUTbahDavQzy45//CpjGrn5WgATG6pwb
yq1AzvrnU1lGP4PH4CIz8fPYp6t5I2ypZImJae7g9pQXYSAK4PgioMpZGnh1
oy75DDoceuaK9olH6JQCW0U4LjHZEmzD/i3FIIP/DDBwu867cqi0yoDHRZw2
F9u9Yb/ElEjHIL2fnVJxUho0aJRfau1/AxIAjS1kI5X20mlQgGsSoi4e47hZ
s2StE0yQgpNuP8IYtHu/g8DGta6r7xunKSvFu0UHWfk71C/QMyhZklrja7b4
D5Dyle+ioLcFuUCOOZJ/r43xSkvF5kIIpS7Di+TYuYoK8Q3NBxUJ6TUU/rux
OPIlz7BsNM3hmpKyBfajDk10oJPHG9FDnEJUOrUeIkFHyuxm4tkDcD8+WpMT
Cw6GITWRSMmoTCvx7NjQS9j0DSB1lYtqR9HXv2tqVIsjYRq/nnBI5k4jpjdy
j6RHKq5NerIEv4tK5eyQvxiiImlubItf06iqAOgB+4wEH3EJxmA6FGnJbyfN
CFeH21fv+8nho6fASmbNL6StqRLlHjNsnkwXHWTV0AIhq76s3Vywt77ZGVki
y/0GrEdL8Jc6G7VxmQe//923YgrsBkmXapCNoVSsw24FwTC4+Z+FaJa6udEy
GmUUyQgoLmuoevW3Hoe5sIv8YguffO7/9wjdMMfnz5fRfqjyfNniqsAfC1U2
EJyaAISPOjaF0nw4lIfE4X4SVPYSB6Ill0H1+Utz7/w/h3885mEKFUpv+Q9+
ZjvPCMpAOb3O/nl+Z5s79EgsEsmnHgUv1sHKiYwwyl0VxmNQvzeISXwF2xP4
PP9jhHkTloZAlxZmHblyRiwEbkJf4eqoIpp6+J1FtGd9/fLrmzKVcq+E0FaM
fg6PWwJYiuuJQ+KIp1iAKDT5AwxWLT8Zqu5IPCIV9uVa+pb28dqhZvgRSA5X
v+NGX/CABb5jZCOIROr2oBGbHUE0Iad+4RG5c8T0uMu7le5leBg4ee9TYKdj
CpAfDbbg1hdcyt6khuc3u7n6arW1nXi6+AehsembE92AJ32+DuBjRZWwfgX0
NqyuOetfY/oJG6R/Cizm5l6cF+A4WRYnpa26lFbmq06lHSDLRHPHpf6pHkAq
wzDubQcHr7UoiYP/e4SKPAPrus6KsBnvMf2vL6raJJtd7yL2jPytBxIcISsk
J4m6OCGCeaeVxynHEtJG4H9/wDTn8JpAk3W+jPPFdgK/+yEs0xQ6Rtr4AuyD
SlGtXoFsLuFJXnoY3ZAKDkdBHenxxjSyZKaRvBe56RhKGlgK/Lt5UtlY17mX
RxXhMYZSMoCVJWwWE3Ha3SnsA+ckvUw9BeSxZjVvUc0nPMiMg+OHFKNwsTvl
RazeJ/jzfF1985vXvjFY04uzRe4zuhD7S5AxfnP3paNdYyqxWj3ZoRos7VNo
ym9UQKrtHd3v5/jR4Si2IHHexM79XYpa627YJXRZ9ko4B1yAKO169wJuo+8o
X+P6SAg17yg8bN76K2aKqykzLGLc3siE4HPiZOygOsweGOmfZ5iucux7b2h9
Rh9UPeUA5p7nehov6rAHMnAhUN3Cv04wyqqbFWQFzIreFijQQqxltLPGR+nL
50OrnVy0czQW5dHfSR9O9Vgpn6X7/sxs5L6bT66ypY8gthgMAF1IGfBMviX/
D4ExlZI0zJyIihOkCDTQhXEzr1o5o//ZHFEqLFXR2TAjOkIoSsYVkV8lhd9E
DTE6kyA2Ftx0YGJIQFNuoocVcdm6yTrkU6+EwdJ+thFyzNt905vNk85q/YIs
zHhehitGPf8A9+x314MzGYeNbUu2mZpkLW35IYdCtrZVknkOm7kbrV6lbWCm
W0U0/0wmnUd9ruheK3i8lPzE3R0PUAGBmyNvc264DjZyJ3o9w/GTKXf0JjeL
tofxbmaZCxn9kEapdcT+07kCXup75lZ8+exumZiB92nHL+yzHzu3FwOmZ3yX
LqE4XHwSLS86IxM9EnQHaZLZbAzlPjsDsjNDY25mEGJ7v+/MjeL2ulEwQmy+
tvVYjn7oUSG/xftO+uojUS60oy3rRT1GlcTfTaHGsv896ySXwNfCJ4iDh4Pf
3V7kO66y3ajwq2ADosjcujXoRfDzkF098kEr02heG1vYBTiR8sdXNQqiaXmt
Ybysi7RsaGRI3HU83on7U7raFDCUTqrC78v0tdAzyMXnn+tyAB7Wgo5qSIh0
lo9bTzeTbjvcUmzFLtzb9adbQoaTLahUhm1iMFNVuPF+WvqDXHWNor8BoaFB
XzdXTJB4x2dp3id9R1ntTuwzgvdwQBySTE31xy8/bB3qOkFcJ72x0MEo66a/
f8jiwlqkQ64mxRvkm7blWiBxe22U3pkEUhzwJ2qPHdyVl7LHpod13sTYN0GZ
6LYR0VzphKeaO6/msNphQWOfIDnf1EcKrrbJ0v++K9KJM/K/P6vLveBIGRT6
kw1YSqSKoNjE7PWla1Pdrf/JFxwjL+WTJnXLOIbTI9EsP5XjKIyaXOtPxGAg
xFZjS0H5+zinahKrwkR6FBxmIzDG7S7lSjNrHQpSK8VSVALamV/m7IznHTFV
JY1rKbMP43+XlJUBnJ9jLxR8L/ebNxOf80qblHvcAbtSk3CUg6YE8Fz07Ny5
xvJB9hvbmPDEKf6AfM5sO45ao5vSIaxacQ4cCVtNfGh0tWXiw0LA+1iJNXzn
UgdPoVWegx9gG5xCd6RDX131KzJ/xdWAeIPeT5LgQNkuZeWG+34quZWWp7pb
Loqy2MDC1Qi4Mj6DtT+bPhsqYS0S+WPUoyCvJrQc9g3+RhQBt3w6aQkl8VZi
ADpS05J4GDbtfBguC4L1n6H6Y+CAjJk1Bzz0+ZNIdkxmwQoJxU3XY7+IP5z4
ZRxf/mLwvGHtflyEu7+BxKadELEau6x6jmX5gbwHzRiS1ENV/LAH+4TqyiXC
MUGgeB3+Lz6GMN6j8THWoc6yoWWrN+QUscveuAju5Zp6uqBg3tDh5rXCCJFy
Ka8nG752n7iGhWL3pv3QIRzUMKU6qMNNbfnto+amNIBc+9r0qabSqGpnu11r
8NJtpJYmqf0NPNzvD9KVVGT3NDFe3bT/ogX60CFR4OAXLVz+fUW7FVPEo0w6
ixxoNp/BjKv4+Af5unlOPQBv60m7KX396XjFwQVbyQLu9G0cuJeANSjqp0b6
9YXKJwiG1Vt6HVz3XbufYhvE9NfMJ7+pun+7TeNa2m9ja+a6Uqm7UWjizsni
wKzWqdFDW+zrYWTc78MLnTIrGwq148+1o2HpcO5bciKqpV0/LFYonTjx4YY6
B2txSJz7MHybHUN187AUCQmiSgichFX96gRcXMBRsiVA6hXX44hEH32S7quj
65VSYpkNXOfWJNq3FR3I814IJ2PN6ijpdvS8bQlLme9VBhHSblzBhXW+wH67
DvGma1huuyEiqC53I4S+d8vMDlZ3QUH5PtTnsbcH2AmwvSpuF5kHiWKVccbt
p8GBCsE7wx5oUjSxU0uH5WXYdGICqJ6PP9t1sg2GN04daan/nazjkB5y1tjH
xCNXhQQiYB4MPpJvY3B5tPdQhVOsjFMgJ+uRVivpiMXLgFvjRpwfWiOrTHSN
PMJ1z8UwOX3f5odIQU+URY1D+WRCJrYHbO+o436/ValvgCvVZREfp2lGBKkB
jJC8ZuUI8QdyRcGQxV1HMczSboeieanePcicF3hn7Do0fAwbVzzl7m31S+Xp
e0dt//2xZ9rXgXn02gUav+5JPMlShL3S+COwqj98aZyiA3d2VDKIBX5+i3cV
g3xeiuqYDYntDn8cSM91rxHhuux0cjJTjwlxhvlBG53h0wpkV1zp5bWdULAZ
UPt83kOqyJ6+4S0yexS20DArow6UlgAiLePrywIH3yeb0LoLblnm7YWkiFPx
Vkq7VMWKIW0OZWWGDmcc2ljnt4HHz6WzD5di7RWy5MlCokrVCvuGoFSyr3Cy
oC6rq42TZYadG8jwsC8T7e76sVRB4AzEncpcV4KN1f3Q1UklbTKchxm6OEgZ
A9z1O/5HprX5cKciG1In6XyW7su32n+82jqrDA1oNVVhWU7u4tqz/c8H6TCq
qJbZ6LCxA2WtGq2baQgHDIfbx4v/+220lFf/Gvontq1+Ft6aEDiXIICoO7l6
evXdaPQprg++PJfUEiGL4+QriVH0ynQaMXb5rvaPiGzqwLGSkYtFs1zj+Nm3
osvhU/rxNMayt5v8PR6E600kGgg17ld1rooJ/LIArX723MoccHbHhpkB6UaQ
JnC4H1BOoQx+6uEBL3TSojy9bgMJAYKkGCGw9CYdXwZHwjP7WZMVz+SId3aG
eP9UAHNKC2Y3j6bVwbFlgQ16Y0YIwe2tdAfN6n3FgdxLXrKIDdl8oqOIi0M4
HJY9d3SI4hdD6XDh2cumBslLw8n2ZS6XyyDYdjs9M7Op+grZ5BvKAjmsR3se
/jRUKLQycjAZw+15CRW9H9LQtvG+cbDVP8xQubf12tuVSDakAknKGwmpuscq
oGQgnUTkVCDvMuyUtV6zqOQJNO7O0MK+tD1H9Mmh2LEWyEjPK1vZ+ahQnjtp
9LmBAZNgNWCZ6owKAHJeSsOtcdIZSLBsGHS6XaZXRIFShmKmgoQGB1ff8mZ8
H2/V5+efOPzHvPUAc4KhuP295zdB3s2qW+JMPeEnzsyjY6GqOiI+DZc0RWat
tgqjwbhxTbpDqaaD4t4UFAl0PQMRnfBdG7LowOthPNoHHVeBVi9B15FMP7uq
AE9TnnOJuou/aG64k6GGlcA9n6D3SFj2+ItKw59w77CFlb8KQt1faiBEdtbL
ZHJ+IQNcwVjoMqUtmTea3yUwMrpsbGenJ3adYO08mcz0GcWwpg34UdC5zItG
cTW8KzQGMXqLzBpiMV5ZYYtdKpBotWBoRDyIqSo4VFQSaibq1IvoHQVYyAtz
CaEY++cQDjVnMCwHkQR9DywvO0plNkxuaD+fHIjUFoWLdV+R9KPqCwvjsZAQ
4EiKztHqLdLUy6bpLUlUdgj7qysKpivCeE353Hw7Q0Wvp16QJfNBBThvuyAO
I+bnuy2pvEV5x73wT5RRTLIRnYY+M1yS56oT1FHoMI1b3jWUvZMAOfLWmWZy
BJTP2DqdrBeVA6dYxt8sHTKlNbZfx2ikMZjkRfTnURBir/GuSvaTA0IEd8Mn
uuDq5Y0SnxyIY4WduB8sRsBB9hYtUW09qlzksHNmAD4WRGkKFP9q+3Q07nCq
tyUYQmgP/lAqwByePUTxdeiS0mUR80SdnAQ/JkHPGsXTBVUhj9lICjIl78mJ
zWtkKAkXtVVjQUOwIMdh3Zs4bWOuNvWKne7xTHU4Oox9tDkd+j25j+kkUZQu
nyTmbXuo8Rq2hCKyzct0rbwRG0Ctu3r6h9U9UeMGfBU1j5/lX2EELC6ZrlfL
YwnpeHMoMT5cDINygyngECrQwfIsGqqNkvKSEAB39vFUpUZxfDkRpxgGgh3T
r1bZjVKdv4faurhYjkMBlZ5xHCWzz+8jYeJYkndkxw/blgsRBrelfwfubfkx
L+NQspronxwWX+/pOAp8umCkdzLMgs7vJj3IPJk2In/aoKfZSIOh8bj2DnAL
xQI6OTd6llwS9mnk1SONax/ibkiTDauigWZUtoKcaUyZJmwK0PlthJUr1KZ0
8ZOS34iDo1/I72AbJ0BWtvAepuc9dKpJyZoZYQH9GJ7n2zzfBT1Q2jWOSoNu
D038+NnTirjFZ4bRt2obQUvr0NfQuB4zQ8oNoV0bzalxCK3grV0T5UXGNI1y
wwPyspnpSrfMO76IBg+zR40Z34YI258NB3KimvntkQ2M7KaF8XoIBvEdk7MT
sodk/LDBbMlugML4BujXp0C/94sPl5SRhMnXUNptLirGz9/CfLiUJcaUs9Px
jd0/vhuE1by4OiZcIKPkoGjz2l0o3iUsDV2doa7zQkLLYoj/9eYvkR7+09kn
6rZEwkArY/Huius1CMYepsjYdpGAbyZouu0oUuAUl6YZHBubv2X6XLYAIn3J
5H91PROLDb/dxX0FM07in/L6HYe8KFHz+TMZgB8hCRGaAEa/1JXLg4xMgcfF
FnLVpsI933CSrhMGsFj8Ru9iQgYazk/fw2dV01pJ7zCb+JAJjtk+pJNqMRGl
j9WGlmXY4kiQ3vnjwBv4oTde12HGnmcsa7BTOg2JScaWA/1WIJaM3Y1GUnoe
mz0I/09ov/cZSYn7f4uIMWzk0Ih3HdCt6ZQTj3dvZRXnq7goXOhkx4ehBEI2
fQKiY7UPHXXU3W81yFBy6Vkp8n95fy/2qPXee68jTGqOLu6bFVw0LHI/oWaS
XG1hcsIRhqvRzLGcwxlaeG2iJMyGUsp6iyYUImyej0ySrhYQd/9HKC2PFmW2
FJnLOEpo4Qs9d9AOFUMw60VAYy2FOQoxai9DuLRjquOWhaGEii6it8ahDFBQ
EW4YEuvG3L8lwLaDNn0uQxFiuXpH3ayZuj7DWBZ6K1rsfR/cmsRu19cgmr+X
2j9lJmo5Z6GwSBQAgF5xwsimFg0JMO4FkKomsvHvlJgPu1c2TxlPJtXJ6nAw
fYMh6OOw14dBb+WU+QFzlbejzYQtcbHZSkMABqJ7f4rKXM2d8eT1fI4wZz3h
PNXOvhOn5Ypp083BeaO3S4VOrhbJAgIKZEY2HqVQ+idMYoiOrK/GNsPzCw6A
Y2YkyrhZQV2i5OoffDfLhc+/2ap1wJ8A+JToaMKZtpIS1zlD4wCnoVQgS+cQ
mJMWUpFu858DvV/OLJ0nLn+XWPFAaE6gqGCSOgO0Zag6eI9HJG+al408n7bU
U3an7lU7F2/xCSMNgurYW616bQTtAW/VQCy2h3siQOEolLfHIKrvWxWo9wNs
PpiTtUvT7o27AMC/zup7JzlAceBTGdZ73TTaiB6k13DAry/QvNa8NEuB7NK9
CXIl8WID4ATVQVWbpTriWD1EnaNrQu1PLdDAT0CPFDmj6k2QhtTp5vbW6Czl
3HFCWYxTQFZfa4gP+e72fxitCslzOgVB9pkwsw1R7dBG3C0YYXt3yBSPNMKY
ndhREvRPntZQnwxDPUp+Lw15trOA2oYjOLEfrRx11X4ZFuDonuoTdGSQdOa/
51of2zixUYwkbJ0RFGBDkcEPKFeLdWXealgYHjcZ2FEGSUtLuV4E3tuIfBZm
l21mJT5BsbyeZk7TsBZhWP9U4OrSGNTpvQhuvogU+IxGcvjqANXWaKepX41w
X8Wv6WBkZHztV3JCNcBb8SIr0CjNIxoDZtUUluLopw3a9CARNGN5yUKpUheQ
BTl6UEoN0HtPLz8ARWffAAGO3nQUy4RRtvMe3d3zwnOuI5SyTHNFnYKXMOLV
YhIy0VCBlzEh/1yuh3hVdlCGhTki+9CDKh02baY44YyFkKeEFTeqCtMLVd6Z
QC/jisHDl2NQL5kitAkMxgqGUzRIKj61XI7ddHeUXUzzYiXmIUyQhcvZdyTd
4XI73/pUmt6s4RbtOibWEpNynsNDDjnsNe3w6gaCsHbnw6cdUb5ubw5W+Oew
G4zdyghSgKStbM0yKK6M7zbOho+9K5fPlhLxSDllamGz0sl5yky7k6hK/Cx3
JEthcGc4B52JYxtUzocaTwWjgy5539mxszgrbE37j9rbeVapWSoD9W3OiXha
C8VWvZ2wNVQlVfa9+Pj6Li8nISnLLmj6cRP2WVZnInzG/XrwXQtIa6Klse9Q
RuxyHO1QAxc+QS6TRLQxtd8W7k3IBP+afqxRNAYFta2Lf4oZ+TtSIC5xpArR
UNAcS/pfL3MZfCrxZQBGrTgGl91p4wAoagDb0I2pZpafgQPi/l+YRG0LU3SZ
eQXkhB1S++a0Mc27ROYcKp3C9Hhwn+RqKuWhcatu30dmLP7os586olqlZeRC
NgF+uu9A0QRR3wryZ/n0rVwmnoifdGfGLTDTIg7sRj6/gNkI84OLliuLtrcQ
rPNV+zkNKM1KrVT/zWOAnM6HI4jKyx3mwaXLhgMH35hO0vJEDGiIF+J5I78+
yKv/BP3mKz4kT9kD3IH3E2HfScisX8N+d9+45X/tGUdYh5uXcLv9CxZ60YQ4
0ceJPI9BG/9+OT4+u65cXNdQ4ouyTW/9kkl1igPhAHvJaBMDtCRbWjjBlCyx
FCXgc7N1ePnDZwr/dPKndoI+OiSx/JEXOgeziCfmzQcButWk9gUttKxWkImI
lcPcLPvSBBcYIYjAM99c6Pk96KLbgcN2Ugko4hMoS3rl9dQITQcNcIo1mRnJ
gU0oOFK/gjSVIamS43nb9zQBS/NP+YBnwjXclBsRsOegzMX/j62jibpb7/ZJ
r9o6FHmoDkwwpwf8JgWhUzzD/7Tz8G8C2jnngX+Yyd7ZnnctH03fkcYgh8Xk
XDJwB0C8/6SKn5ftJPhMeUneHztBJAwFjdxLHKYeT6MiciZHuSXvqY7bBWaj
YHlsKS8nVUH5ZQlKvb8yHJF3ksWciFFAbHSaeQ/e0tkd1uRZUgDdJrLcf4fO
A1hTtyJjWTWn8dLk0c3e2ddj20bq8sbCKWS9PbTtaX1SGz3QHn4NKlBYLMpC
FMAX91h9XsCl+tU/qfKWkMuU2GRGLGd1Iez2NXUB0M8BgECUsmpFIVoo5YPB
iftFll+bqRU8v+8y8O5n7fjuEPLo4S1kUm50wry87V7dvTHtN1pf9nVpVrRc
NtMjvQdlzGxZ2ZojSC4fx9Om4lbpworYmLxXX+WNIl4Mkx2HPgHd+G1PRWb+
BdsNCplbBK53x/bCU330wpqOR9mQOteXYFxhAxCsnBt4jRiCVty+RuNVp4Jt
TKaCP54nuXeRW8v/OcSi4yE4lFErF/xYRpxQh5SRI0pfaTiDUK8XbOgO86mH
8+Yo1PpqQrDZVD3ugAEfwiCIg7maq7+uw4vNUUik29RWZFoF+UtuB2AZU4hL
lQpYNNK1Y+9h8rbMHMrkgcMU6+pmIv3wpo8Z6IUQHF1nsoIZGIYBb6RxyuHj
9xDMTJbNQfZYe785n3vpOd5A0bF6XXj/ccOLV/6DVdLRoqvJ5xdJMEZOvjW3
9MiLzeHWEFglM8hsXibjt+fzWkSzpqyGHtxCs88pyhDMJqL5VFy6FLJxkWr/
EZziu7qiV78qrducLzuPQ+efgzIkgoXbLmrY8oiqZrMQx0tLd8G6DuOTn82O
7CgvsdPaICjlxkZnKOm8J+6v67JOSizqPYCB6+c9UjdBzDQA2/KU5ZtGTUWn
gBA9BxkVhAMuACX1n+69/7LHJdcPw75AcwSwK3gFoV4EwCZapsv9MIsJwNl3
E1/zLS+tkWE1HhCJOHV7t+j7h6rcufu8pLHKQOrNQl+ICiMmeIIvHuxIAGi7
K9xosSfgY6aEZe0B4og0xp94LjwVa93etT8Xg7ZXK3GEcQny6RfgVGf39Knh
8PnbO+FkYJ/YQRj7/7rK9y0Bj0J9bpt+wmsuluddxBXmB3f9dRYGyao3HgLw
YOE/H2lzwy9wR/A2XWc9rRWAqfvt28TiiYee4Ws7QmEQdj0Jz2c6WkkaV+c5
aJaVq2lRV10cA+t59PglNYABrIqtcTPRKa+zO+lbIiAflVeBQYJkn6acedlV
B86HKyrgAg3uZzrEYoeiHMzpXzW1M0baF25iHvFbq2k9Zrf/V10vnJ/WaIXT
AR81Ifj3VhY9o7dd1zSxmqHw0X+RLy4IHCe0ACTkiixKFdLFaupAFGM32Txz
t0Zki1P8ywXNsdQ3+29dAVh7X8HSPEK9Mmqe3HXx54QCMoQ9hnSasPHlg1ib
YHJe15HXbu5DUz10yGE5u59ZKIDz8BaNt45h0i5VUKHr2/jLbZLQ4cG+6Ka6
6oelb5DGysGbyboJk9eQXW4GInmwFAnjbY4CB0NVroe7RrWFVUMU4imVOqhn
NftTjUXrdaq4hmiujK2eo8iapBin5gYxhiHYZv+QwTWJrCOsk+IG6VYSEqlb
0Z9YHBdbBFxBHqxJGEjAWUHN1Bdqvgwv31OGMEfetO4hoE448T8nKX0GmJdY
+3/O6o6nZQQIgzzvURuUGLYPLjhboiha2EIGeQO2KMfGxU3eZFa7ASWmrT/x
i/Mj5JMqrQ/47SnRafDIcyt2FIvcw2vLFTdCmBOupQGwYn7AC9eKDbJDiknk
5Hj3FJaZ5GVRlFTPsHGN5/E/Ij1+Tn7vNKvfOsEkIBxjiKGaXolMXporS4cQ
LK05fs0zCnayEqxry2s7cqTNZapFaX1VYPTxtIOnzQYJzd96Pj7WlgCsuDOQ
+bV+qaarMBJt9APkYSVD8tlQT/uLxl9gQ35akc3AwqELgxTnsVodalbxDE+m
g1v35rxr1cuxCNhZ/WiJry1sQIBstd2pu+3Mgoc8Zfp+8vijZPfidCUTYSc4
qVV7SLNJbeV+f+Ri7/zu1IGMxXNck2bo4DAQAIr/KUyVCbc+5ZCf5ocTuBcp
2P2tknUBxRtkb++GnRIq6VVCmJ2RiUSaLgi33q4dQChfOs5UOOVPviBAj/oh
7KdUIOBGkR2t+14d1vgigPuhNGEJTovICZae+RjwuPpebrfYYl5QkNBRuKoV
vk5LfU9M6lms+9sl9ewaO2RjT/VAaMs+nszbnNj7tmBc0kpEP/BhZWaBoUFO
ZnW0I/iRvJqkNYWTsF7dltP0/+QcHgjoH0Mp+o0+SwfANC2c25bdCp1adUB8
cmd9d3Za4cCt+gc4ywArBDZ4cIgnvffeHKAmRDg69rCl2cqf5VDCiOC0jBZy
Wl7cvqH7J0iT/eQmDkY+EsV8d1N1yGc1XpySNYO6MF1hrfXN+gWfOyQwQ6uD
n31l9A3w21e/HBWSL8mVK0TC9a3yqHlLiJUH5zWaLPqNyKt8wB0RGG+Y64tA
DxE2ipET1KXkoQoBlMBQRLJH9aTZqzSGKODjKl/9QUxeYlzgaOFEKemtrvlH
QrJPKItb9+VI4fnN1bJPDG1xgVmP258duernzT34QV5voOJ+9t9cqFApM5YI
g/xlRwwZDjnLKSMT9IHmUjvs8kQ+H7VzvLjQ0DtyiMP4mUwuazH17pmTSryQ
5OCSEJ/qyiG0iL7ZQPvvvgtpjdSZU2DfwuzPwvTX4BrP4FuubooaYCmJAoEQ
jTYRvEJJp1HKChb9XvJsXibjdhx9zFwG81kDmVzLLzokEckUNm21pd0pGgL0
GN7dxs/tEGyr0ykdOiNUQ0UsmF9AdBFpBYygDrUv6575wFZLIVfG6WmUCvYR
mEFxLaGGQS3WUTsjEeBH6a1dl5cn5YHtEDyIPsg47iHfgXDEC5fHXS+qpcLB
PzQTYJ8+j7GExJjeG+5h3B7FmrKUG+XBaRoAC6l0kotIkRL3RsQoYZ0eNKSE
ayn4w4m5Qa1i0o/ebeV+j9Aft6esBYMppz9xFtUSWRVZGRnaGJg7XYBDdVoX
kHeURTl6kZl1hOiXCNc3F2NdDyoVDCDr5i2z7ckxZbBhTzEwZA41vc1P5CUb
M8ySDvASZ9pUOTxg7BvRY3el93w9FcaoBzbDtMFo9g5Edu71AEXsEZc+Kcml
4g2ZDGhi8zWCSGUFhrzUHycWk2x8isFETPRV3O7ruF0zB94qHE+ZAuK9UWil
FLbqsz+MHhtsUU+ZHC+NfQ6SmvTqBzvpmQbP4b0QPimfu0ua4XOS9VoexeOD
WjjgwwdPVSLSkYFTVw2/eWFioQCi9iu+B7+zPnjh2oqR+W1TA7vVVCpooNj+
KIkFKB/be4cb74FSbOaGJa0G4sKSzxK+DpNOwHch9kLCEHHmAWKBEUbdOY70
/ps2JveCP1I4AAk50A1AzkbCVnR3KU4c463XbUWoqOk3Evg8RdcoLcerMVoB
tC4xdZN+bmzhWzUFRhKnAOAI3at6wEwtyGNC+ew84HZBbXZ4jnrEry4MsmNn
so4TwVKbUulV8RB+/bWJtvaFuXmwESRatuwqsJpo8bPWkOTcOZ0pauy0d+Nz
bipD1YGpoPwkYr8MSMrVKuX4cTyhv25w5pKJnxGwG9SLLrddiPNZJiWzgcG4
ILFvScsi6aKrv+vWr06uljHmc7UNIt807IuK007pzZd9cW6KrxUYVs/ckPNN
XnIQ9tDt43pOWyLrhHiwrKLtW67sgb3EmGF/KxWAxtCpmcyEMtycv9HQQdZ9
WxLM2yWo8Oa5ktLBUdmnS+9K8JFsw958ArK9HEoATpzdNNcLMjYsCMrJJvjG
exbYJ/dRy0qVVZsViax7xupqskymqJIqKlFxpBLGCWpwsIkFZ6Rp9sXAyfUH
FIiNQckGBnyTeBi8XYYnxRJTpHrFP8mMp+x2wuKKHdW8yMuYsxpBw59rtQoa
k9A5RBPdwpEAGHS2ZdoDS4c+gXoCxVYeleoTT4y8alox6t2e+u0q/yzGjz0y
DJaBVc8CTQhyxugZKZIUdWk1A3DlFQXP5zQ41M50+zFdSFK0t4zBvmR6dm3V
PlrZfTJJZFRhY4DzYSXLoWJh5jhXrgeKmrCwHS7tn7ik0/wjaAjPtkj2FTmN
HGlyOFahcbYCzL4cDSYzcaQCph53eRo97qUY60TvGYjqjq5WwaZ/wAgheAyc
wd3ZSgmfxFjzAXO5Nx0lNiE7BhfrZ14LoOzfdTb/C506CG7sJQ05HQhhs9Bv
qF6Q5ptNN6yZZC0YbbFH3lzsUBgK4keTQoJJWJkFwcoTC/s/SZvJKcPaxgvt
Y1K2RKJNFippJlMqhp6QWFirkFGneC/Rm8X7d2RLHO+lhGVMfmToqXdK3bcY
KR2PSCcW00XOfRAPVLSeq3/XkpnofUhFFZXrUrWF68kjBDeeK6epFEAeSgwa
M52Cc+ZYcuYqjRSA9DHeOp6PzRO0C6xwiEnA1QoO9IfJKj/m60PuSInhlzLY
wQhOHmbsGJeNiy/APEQq3DPZ/OG/aLkpSKBhcvEchBv+hLzy+Z02ha/JUCkP
U/bACSyAx3ZebmTRyWCYR3eyHRZnFnsDumm1Rhy8GPHbYibpKMjIleDqmdYF
vO+CF63E/d/Ka84Rq/XVcNs5agEH9/LipHtF3gGsea1We869SOpXdoil3+cC
xzK9F6yEtu4rtUoQK1yypX8Ux0Koq5bo0iHKTwaUkCZb+TMewk/Cv/O+uEV0
Tan2p2DBi8pW84OXKBKZEywunZVBBGBpOQqyHH15HeRt819hkPuEnUnVofed
qJWrxea6OKOt3fwNOsbX3z3PTUMth8sl4OFiP5eeKReSAM3OWXmPmc7ObFy5
CkvNsixQyn6cGCA3InLvYAta+kisfCJIzlijHxRzQ5Nh3xRGr4p2cxN/F4gQ
cAEKzvAoBZgN5CgSHsiKks17lIu7yOcFpPkKlZj/dk0vdDAfGm0shFdMIyAM
tb3A7BJ5b7Dws2xocm31C3L20bUo0taydP7ribzyOfotb+IwJ/cgYmUX

`pragma protect end_protected
