// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
otCuvlsUFnU4kLzx4QREk2dj6VHq6y4iiqi9XPzAgEG9SGMLrJy3XLgvzHSqnwUP
oItERh6ajVTAEEeZk6wt/Aedv4Z8d4nKQEdoatR6JWJ9ggh0yS3IYjr9XnVqknkX
dkbFIIY2NA8qDYrClRCIxy9T+EgaU58jCUtd+w69FNntbQ6Xcy73RQ==
//pragma protect end_key_block
//pragma protect digest_block
NrsFTgflzdXUzgrl4SYiWoItSW4=
//pragma protect end_digest_block
//pragma protect data_block
cI/apxKGCepS8wG3jB67X/z0QzJFJkxL7wHJVXV1Ti2RKvq1EO/GetbPtJvGr/sP
Lrncs5URN2KwaPyt5ntnFKw6d1Yhlc29PxONPOqERhoUE15zt2PPGI/N6WvL4bMp
gJvPZkEtPtiHUaF2NrTsp79kU4u1BSwk06DI1Zihf8+/f919T22L7BhDWzqBzwAJ
ghocd6MvxTQ+dxzpUv9J2OoM3b1/YbdeL6+yl5Qb6NdJHwPs5StQxJpUVjRIT68p
PRQLTXRKEYjuJCDakm9WA+LH67gZZ/b/X84/hHDtuclUcYpivM/A+cf3sx/SOtyq
oL6kzQZGB3xo8UGIAvHuNM4SSz/aTDOA7qk9tWvowbuJcbSXW4lQVqKQ58e2CqD3
2XYkkIYzDUiNMHlzfSaT7AQDzxzbrnCoNa3MbGwiDEqnQoWkXH9TUE/HyADy+GcA
4lzIgFOpJwIP894lEM9U3BUP/PHnpfMB/2SJtmvbBTjOYDIqYshez6LFiskLkVrU
k5205HrV2fGsU5wr+I+mhOt8cMAyiXzDQMaHSwpguC3M2sEE5EA8iCElTuOeeF0V
74WZSjbiwyg3G4gq6h1floOugtcLdhjUxjw/qS1QEQJY769EiaVeUcjyPWAj/CJ+
rjtdWDwp1cvejez5YeL0YbGkHnZKA05XMcVKyYJT40ldom3EE6/ZMG5R3MVeGFWV
jBz/yO5Fu9WpfuEvgLOQO3K8//U0/qwvpZGInNoLzdHwz15kY1D/+p5XTBKwUxFG
Fhch4SPp6jt/7FzPH0egSZgi/W/Tpqaw3H2Fg+UJhCLjAl1DSEeWdbn9ItxZMrJd
zEjXvJRtKxJH8qWcXrwK1n6PQVQRtvPBNdEGZBjYOPrmOPZQebIYL30BjRuhpZ7f
FybmYC+cQ7CyooLTSgi+udvGZny4Wo+pcRTFO2JHnhOLNYE+2987wd8xlb6fNPWA
TNkDdKdefUcRg+996UJPYT2mc/XC7ISVt49/x9ppEKfqoYoD3bwNsYu0x9pEEbrc
EldjIeoRtXp+cWOrDxtbm+GXDd9kT9NFPtoXthxqwFNe6JCtgP3ZeQHHCMFrcBNd
OHRHanMNp/OllLD+7apMo7h8l0Dov8tM5Yv3piOPhw5N8Ogxmxsw53tHq3bsLmbr
N0s014dHDWGmRfKJcoRT4zGyNmxEC++M1FzIQgqgYO+B4C1eA4FGhPjaKu/tGosp
Rwb7J9AtveNxawQkonnBF2txA/8rUpt9VLQOyLyDLrwoTV2tp9xC5y0JYPHJXUcv
Q586wF3mxw+g10DyYHMmLrZJUWzCbKceT3gtzqIWFCoTz3lDsB+42D19dE05sjsH
MaKY6Gm1G44Ag2LV3EkOI0he8dSkxcaLNTRoSg5ltR4z4MsDDi4SSL8WPN0cQJyF
Zp4nYjVGOEywNHAGGOfNA/lpxhg9ZORYsGwBPfWCdNysSAzMu1D5ZLoqxUC+jJAv
dCHHufx1ORlbK6S5PKwWTWDjEiqfy6AMPEn0Linwh00x6DPRHmKrB1Uslo6jeztI
r5LvWyOPMNyhaNny2QYv6e2GlftQqCFswJ9gmD22+swLrFqnnAnfMMx0pGo16U34
nwEKk2Y38dQE07LghkchuJ/rYolnpPudoJgefmH1blEsLPogLSxqBRzvquGFV9ur
qocHS2naw1TRQBkpwDPAFwd69WSYs51qVg/YUb4RwUMdZ0RjU7XYmybZ7Hh61heU
CSOud9hqXOTCVuzlCjp+fws30eOeFwNW2kYvfxudJ3Wg9/fz6ck51BQM+cdzyVUH
S/PgPtVo3GoA5G1eahTOq4ahmzrzZvHI5+iZTfU81MuqSDRLSLvgQDbjaJ9h8d1g
w935xrr7SZpVAmbCvQp5/qZ9ObVu8xX5rYmDuhkbdmoSp1UgcQaO5h0MBDqsD4eO
nykT+PdRm540DLklEgwpmMeZ24JqHdS/IW6O89L5SU/SI3UfPR0W7Brfj0pegwb5
hetXRCQgkqigmu4hr4kGy1TR4mf7DFxxqWniiNYtxM9oHYKYW/bapT/3EUWzuZEb
KZv/w5925vKYIWJ60k2cf4EFWAAPJ9sd3No0/VzDTuGPJRD28kzOsMP+4Gxfy6gr
lzRfgq4q9h5AkJv+EiA3cMTcWtB1Pac35ezrJm4BunF5EU3UfXh7y5AubxxHEDQj
ZgaHFP59aNoDexAn7XN4oxMvsk8MgYoEZXXJMhqe/mptqAbLA1yR4hGFthSOIkjZ
Gq2473SdLn3eISCkePNAJyVCdBRKdhL/IwMbH9CltjUdRWmiDYD/YbncStlxALB+
qhlslK9qFaIfWZB7PfG8riZc4TsLpX8WaqHtCf1vGZu9cxP5yHin6Fj6et+2j+wG
kdXw2uEX2AF/U+svYaX3G2GnYqX2F2ONTNPVj7FGUD/ybK3dL9Nm7VRG04WOv8Rg
aynWx+tSmzuO1yZHtY4WjlBXBR+rGrSyKNDueOWOieeqkROkFKALQ1HQhaaih4cV
3vfCLcCzO3NYxFCigFwl355wDXRyV5/Jaj91iuIeVmQB/v467M2ugEk2CwmUYubq
bkyPLPWe0ppgSFl/PhKv0ORV0O6ZSfuqrioYTTEN40YfXIn93PLdv0kjUs/aWdRy
SsGoVb5s2oLTGzinMOdiqqvwXHNgf5fXzzFyEIdmhBOjLvF8CMsHwod+35+nGjAJ
RSp+mlIf8B8rrXWM2HmY/iIlYp1Tx3b4YdXg9LI5H2SRN8iDZ9HXR+5C8gYu8h38
+2hBnt+e97yk5wQSqCUzCkKWj/UWvtk19i+Wv7tMdj4uuOliPlsu54m+iYb+kYpM
N727V19CzEZKNR+dcEDhvbGnvGG/DxIwu913eMxHVQzSMAnoQiD9NJmeecwaTKaA
IjGrqZx02AVLznR1nwylUhp3qe+60ydYztu2/osReZ7c+IrQhTCBL2Xb/hDKdjQc
X79TP5OGVZgpcguG3mHY+gUhLjnnDZx5JWVFGL8K/waxP3C4szm4lVf/H6GzNhiS
DNuAVKOOb+LVTCXX5J3N7x7Ip8jY/jGHziVrKyBxNl7/vjyJxNLMRiLEDhspFZAf
Fc0h4/0MxEOFD7k2CKwXCpJCLLfCZHxKF03iujef3plCQGSgh3kwwFnACMzceyU3
QC8lwUe9hhIvC08EsfyeT3GqK2KS1QGxNMyRq2GIkMyCvuGXu4vokEWJN61u6D7J
qlSObYOr5g94hvnqeC/wJy9s7zi81ql3opwPgmcE5qG3s5PxvWSkz2LXd13ZemqP
3/qkT/tmKkRiDoRey1+OKTFywmDxmuLE8PRNyyDBWfyjrjDp8xP1birwW9h1st9K
5zdkGBkz5oOemqSzhkT0Lz+F+4//wkawPqlW/+HuYQQ/U0jaSSNYekW4j5jluw/k
OpVwoR5hAe2fh8qV1QK1QsgAWU91RPIqM3RBl1yQ3RNZzIEW3zf19CAQwriyoNfg
22yIyR65UBFwav6DzzFQScrqy7ERAH/yro1OHtvcxfQytUziD3vsaFiRpD8bRZED
IL83Qr+xZKL+kUrnvH4xCEeqs4piqYq3TTVRpIIZMsxUaTBOOK/3yLM9bbNgksip
prOeYpVEfWtWc9IOlKTqg33R808jI6ZBiZporxNxHeoUeGKZSAWx/aCfXsVXVIUm
9bfoi8iLq2CDIQdStuabbBElNrFVud/hUtf1mBdbpjBw9W240gzwZ0mXanHZo6Nt
jeZYQpcOfeNJ/Yudav+bOeo24KBtyXKlFck02K2ZltY/tSA3JAO7fNL61D30yCRl
59eQ6q8wisfekE9Mc67dUJ2Zy4YvvSS3whX2qYMAGxP16RWIB8EO2SA8evNlOqjp
L9B5+DEe0fQpg7Rtp/ppUYNOg71/0JRxaZZs2ukwC62SZbGRtOM2cO4b67iNd341
/cgfWsLL4HfCklW3IjH2v+y4xoiz4OJb+jtFyuI8H3GrKKR7qS3UcHJqxCAbP+Qe
qEa9SxV3ppVU376dthJzk99D01jd2Dz4TFAalQIucqEPZqH+ezLgNjkL6ot0Fe/i
zWbj1yBNTF4wIxsUyHZYqIFgNSbpUEfCu/KR6Sy2cAcQpICxL3maTepAoPQWwSK2
uLbjlWLbW3j53Ds7mc8JYtAaCZrVEihPUosR/mwNDAN/LvaMfr6970AZYgTOyr/k
/VnE1oLZfs9PmZ2DGY14EGsghBjwwmKAi6J0PeZUq1peSDWIVCJaHyfl//6RBTte
vhrpJHnk+UAXkQirvSJAlIrdxoqml3scpchFGHJ5uj/RNvNahQKHLJzx1FXIZoDA
lIZVlWov7c2kAb4NlUzyyswtieDzYw4buGsF3HoiA79v5BYFA+wXZsEVAR0BN8y1
LyPE1TjGQl8AJzHIUacODB28V4rrXM67NgrG1FyYgD1uGdP4mf1iFM40hhkkExlG
zM5pt0u4oS21NGVXcReqQ5uMSK5h27wccPT4T775GHb1FhfUnW+3TbvjuB7HuZx7
h6VW38ggounhefU41HwX+ryM6pI/AKUwoV9+ATjKOP1pfD/fPUf/kij6aKstftR6
5++zMPZN1Wq4XI7mhw8O85oYWMRg2Org0p8+fJhBG5hcQIH/Sns5O3PCQekImYZz
Z6BBkZhCyCHCb3hrYY8HRsoE0a8sjSIJXPhAEwrqUQip8GPuEEWWrj+hdjB6eZCY
JstRmQYx57wLrO4r/4y6YrDaxc+78+IUgqfY/EEBxUAjxKwJ9csP5ptl5KMUxzmy
iRYXfbj8I7z3oQ1gSflatqEB0ECQ1sWIosrP1QKSIp9maRq6dSqcm7+E589soH8r
L35CA8KYZwbhTmbfOJSaqMXu3+UnIwkh5pV+1g2D13GekL1ndKPN0Q6Z79uD15xy
wJ9VCMAfVrkxj/sOLW4/NmqGJB64kNLNtlqvWP30ri6Hb8w/rqYykvO5CWg+ciuA
BB/mixBbgru6a4uHGij1p2jDpsdGw9gDxP7y34MY+4q63PXPd0T4+SuONo+adxZ8
oPo95Ll6T19suftXbxbaLQ0fMZkrHLB9SdFgqXX6B6G/x+xRWNrrhIJn3I36GRlC
hurtCCXpE5tdk2z3Zq6E7UPC0ZjE48EXl7Ve3TlslznmJAmbVqKobKQGLLQ/eXI/
R1MKQXVggLhVhyfZNiAvL4/7nGOgYWVbwlJAloBw5hfwR06TmZIWENGKpZHxH9Gc
MApRLHc/70eoL4hYWjDVAKuimTDjVGkIXHEEqBlaNfRpQpDZbOvflOh/NWfSKxzU
dNqIx0Lo7h1IFYQAFvsJCAyKyXrtWezxBtA5cz33FIioss2yG86/+PDrgd1OsWB2
OlI1CF03/2CB/e30AH6HuwqVymxzJFO0r+tTsE9tSuYGM05xwP3PmajKZW4FxPJd
VZTfAx5OjnQyrTle5rgUEUWdZaNBNhGGZ+oxFxNXCJdeDpZ2PEmsuBGfE6rgm4gI
0T0OoYO2kykK5Wm3RsJzSJ5S2lA8UD0IzSFgYXWnA4GFfdMbBp6YlJh50R028Ys6
8sCHj6NTg+JLVtWEBwKKsNu3odwIMiIqgc31BhsZs65ZIv7G+LbKVf4UVuw0c1z5
XfL0FjldJktec8VQ2YvrFxJOM/iSh5fmf5nX+WPzRa6yU3W2z3zEW92jAPSInTxD
RTZxaVCHSwQZgQu4QRiZ26l2li/qg2FPGhBUSRGxJIW2k1jqspxaKIOin3Zxs+0t
fJPmYUuOETVAP5Edp1lmMOWfYVVC2/uLr4wBSznIuv279smZL0IC2+hnJsTprHsx
HEoHZENG0mvt8Zy/SAkPxsvnqBwYWk5H0TPjVZbfd17XhEwbTggjnvJ7sIyZrSNz
WwjxDu4eIxVEdTfV16XgbGPKUahyBqeqo5D21jYHVCkwxnrqbwxXWCC9eSel/iLx
zAOT/cHZUkLOLpkmZaahJPXaqvOdbsOVXIiZlJAVE5bm4WIuWnq2tgCjOfy52GgZ
U5x/7hhbzqZNyF9HttkXqlie2toDr5+buUV8pm4wHawI0MiD6pC8di0oe8QKvyRy
+VM2A+A+KUiyW82gJq/8clLQlsLJk4Ilsc1J1EeT8A2Iucr5ByurCvlsxwlpcWXW
XnuZgKzQh6ax4bpKdpcQrnmNmfZFTq/g5rMBKpZoUp3jPG5bZmbu+cv03TM6/8yr
8O0KiWq6X5At4ak/iFuoLAKdfK0ZQgP3TdvyiTx98ODDz8KOqs2L3cYmLNnpcA8e
utUg0IIwv9+gkQcoLTsFkM5nTPQPtOdKfmS3dH1X8jXCoKKSOIZ3Bb+R/Cg5pY/G
DmLfJjhyi6WFDv22yqEUSHUC9LNqAy2Tglu5/i/KB4qywygsqHaqLEcIt6qD2jbP
ZuhKorZamy8JPLi/q5DCLNeuoRG3m5G9aL7mSRyzsT00WzLMLO/ij0Gyz9gWN80B
+72ahO9zlFmSVU3ZHPkrnqG+zlgwAusVXRZEa3KG1x/MuGtOWO8Va7YOrX/c4i/D
pDq6tpxbe1LyJB0PsVrmcTrLa9gqtxJRTieu8Iz+vjNMyu7zYAF8ZGL+Bj1uglya
pmBAy2hQ7QxhFxCiNBUfCeWB6hjATCePl6eCRnqbiCtYaNWhW+ZcSyfsbOZCaOL5
3Cjg/Sn5APBgddGTKDn1IShUWp2c2Ybp7TGEVRIkWYeMjE5ylXlF4062fyn0/t83
QVsgCwQgfFuRL1Do2BChrPJ0S/UldTrCQhc0tXFQPN0mnjVau3Ymy5fJ9aQH4g1E
8f2jyOPflHzaldoKK9IY546aqvfAFTkHUpNyvsLbUJysFLPTutvV4Oi/KxDJvDF0
hTn+QtwPnTlCxJNpiVj6slO2gYt9lHBALcmC+5UW5AokGtrD+tZ0zEQQincf+Ysr
O/ZefyCZvIkV7Y4Qd/Bbn5sftoQoS9hB65q4NQOt92Bmm1a1B9MTpH8K01Qbv1Bx
TzgHzQfvRhRjXsWYi/TbdjM0ukZDCyE9OohQa2ky6NWVSRJJfrJUkgqOmXttpi2u
1Ixnr/0mqu/PdbaWvfVHhr6ZYSlc+suLk7/c5WLqWqEsRTVIuI445x23UP+lVLmI
A388tFz0dH68JyUeDGKb3KDc+6iBBMwcoJ0/S8Ur3nwPpQzSmVvUXJGFk/kwsGcF
n6eQIWRQVpfL4FayvZbh6rjw/6YshN8X6Et1MG/kb8aU4+jAsSNmeUbJaey0PvDg
EUW0uL3Ioy9wMzpnXthbLgECQnmBdUy4T0KO8Jh1COpviC94ubRNeOpUzEsRgK6O
nBVodqLoRwujyYC23RFkY2p5Ud9yqhkF7Jq9+qKZc/1+sAn5Z7kD3C/kQ1IxubE7
hIAp2vhEDe+Fsk6P4fZ1om0WedmkybjKyOOnY5FjVwru7wweXL0evVrxfi/YnhNP
/L22kmzQLcY8JCpv/xb4l/cLSP5nWwQb4IDQfy7clzHNExyL7Q3mbuQTojSnqHTs
7Vq2yEwDwqhEnjSxhjfzJWagJffD31Uiqc/xh74jhor+NJrKycXIeWrQjGhuGOkt
ks/cPz7MPIIdPfCoYPl9EjBmwDrg5dkwaygXzAqdsmJi32eZDfm+9UN4NwzPcmb4
Uhd3+FocyHLoAkBm+W0Moz8ClpogpIGveqz8Ri7KghK2H6106Hf1eDMpS1mH3hn/
nO+32kCzI1IALTVCTEBJhOEoPWgDomVUqduCXRPADV9qj50jXvbgGg+pJB5OMaPD
ezga5FYGUeBGcdyI6T4vD2m5NH5UZrp30tDaduqegV7PIJsJDO/9UNNlPlHH8v92
CO/UtWx+qobboHs+ZBxfgBgBh/CKS7nKeK+yma4/NAJiV+DTxkeAJmklVT8U6tHJ
U+ESDpuYNLCGShsJw/23SheKgrqiKSQKleB8qVK+UN6TmyUaE/u5srB0r8HU2bO3
CICAhWUqU/0J1y6b/QIj1RGb6AvPRvEFdRGK/xHNGJ8DqA+b13f0sxHVuRxhxr89
8nMw6TfH9Aqiad9CDbBns1AAV8W5q2il+hzxRyUj61OUSYLSIiMLYUzvW2huF0DR
3nTqJ4kf4PiYaqXatKCbo044H48c4/QBmpUMevFvc11BSiNDN+oV7BHNLXpINVqj
in0iJDoETDWW+tTPKRDoNJ1Ybk9R7V+riiSs2ADHIII+/2HpDTiG2r1NMCParuhZ
JKzW5QWjLS7cFX/WlTlsU0MJbtgTeLl6e9PjRE6HSPZL5+xT9TAQ2DOHozwUmzqK
JHbVyVTg9dmVCi4JfO2l6KQyJDIOv7SN9aiZ/EzFA+9o73ItmMuUpSh9RQu+bgmj
TrgfqZ3eVOxOeIVvpiVXRmxasElP8N9gF67JdsJIPn76HexE9MrS8EKEZpaC1c/h
Bm201OooOxDZCvrJU4N7mm30y9BBcvoNOVKBYkRyA4aFfQFK7hBQ5xkTY+2+XtFw
UGBzGDykc3iZDp62Lpl/c5k2o4qtQgcsfJ+mQ1oEkeL6wRUWRrBb0IkSNKI+YvqG
xsL2LbIgQFy8SqpsWM2ReaXeVFOAJnTuCf5qwe+g5rX0La6ZoCRi//inhFbMK1t6
pZmNaBWNmXpWLSdAkRv3fzuz/omO62LgEIYrO134U1tBcPOQAulcuOkJhQS4e1Tr
RNjShwONx+iCzDxnKVvLNJY8vS4ilZ59Cd6Fy9J60Jdv7vOLPGVrI/2ib0+8dvAN
NHkVcvXCkfznBiq9OM8PAuEZtsJReiXfwC5/dbXE6u5ZN+wbhdEi8ey4BZWrR89c
CYAQO+D3xagRfxiHU3K7YO4CttXHQ1L06HPOs+JvjzWMpGHexNRBRO2sWjvjnkTU
gZKYK/iC7amo6599dlF9dJ8kOr2NJORZvog5Nkxs7Viu5SeQGUuy9dumT//hJeIu
v9koc/PDyDhSl1X4YL0+BHzsFpgV5d1jM1061YbwpdKKslPvBNXWBh3x7wYbXthC
lI7Kj9USeg76/GfjiYIdNbsmGM3LceEXHeX4zpwdC3PimDc6VbHWC8A3k79Du9zY
qU0Jd9rAmfw7LKSj1udAkdS8JTPunrpLEo5dxphMfrf/04eeImniGSAOah6IQ8pT
uonePADXNwMKbGWmLpU8eqOYqpvzb6ybb7bt65Rm08FclJ9Zuo8fNi3lmpiUVcbz
L5UIkMmYz6tpYYkWp9lf5pYYS8wJdTNgNlnPKmrblBgYArVTcv0J/b/nlVVGSWcz
d2GFVkHnzJyS2ZfajfdJ63BbCT/85uFp6kQW/JhecFjb30svBRXupDRY/59x5NoT
yeHEwxoqdf1q1vqYGBrw6Ag61EBcRI+Bp2XSysJWbEfK3tGcp8yBn+5yNXgaL+2R
xvTI0cSAvm6PtSxfOlO6lajq+NvnXh2jvzTnj0setMW1rcjh9J+sNO45g0ptToSt
xM2ewlTL1GfP1BSgnHBJzg+pE+CMV51SQdt8sRA4+GcjJzU49BAKZEuqibKUwFD7
9pkIWn0ga8G4VfzcGr+UQzp4UF1ajClPok7jL/54gL8rrXg6b1+x4MLTe0U0jPQY
xiK6N5XrscgS69LidODuJtHe2uI3mc8eJIh2JUMg1fQcpkY9FooRfM8AFmItWwI1
Buxu/QB2WjO7ykNPvTdZtFk56L36S2bHY0y29lAq3/oH7EgUJS4dUEl2Jzd7EIcy
VuNcKLhNXvbgOkbUFSsc3vgSBpzYMG3O6K5ImY8PvaKOeT0ln6tk5iZcJchpmZgR
Tf7AHslPUy1TFvVudCMOj0u04lYxr57mO8YuL8Vu4AkPt2APmt3hZiNVArMAvwvD
48QJoQec8VV0ediIJN7Ctm8+YXqLkmaG19DdqQiry9xIq7zg9I+AtakahBTNPPfV
ARfl+56Zmb3ETTWqmpxZ/Jb93BJAKJmuio7IQiXQCVSPzbVg6MCtUoNzU5pjFVC7
booRXTIHQgwz5zudx3RxPRdkPgQIp1AmFF4I2xHWnxcNshX18gmJ7v3RZtIe2Qb/
obJlWlRN6l1N67kKOVa2vaRHNoS3MMB7gfEABwlXI57o4Z6JGvpm3SV7hu5OecIr
22MzIyAlwdz1LnEddT4vPSgQDBv7uWDajSL7rkoZRfvcYyvvq8a3qOlL1N4Mgfjo
rWeHSwG1SsW3LlcS0JMzOu5UpmxQSvuQW1/s2e6aid/EMLoZdnx3VJ/tEyKAHOL/
ogNRK4emoeXv9t5ibinKtnvhnFrhLmYQO9w9wpfW0Zlfq+jxanAgbZZuWOqXmqcS
szmclTdq/iKPIaq65Gr0m4gPxC4sSst9RnR85QbPLbeCd5x50xHM5YJkvjRleuVz
E9KNPLm/n18XYFakCNj6NCEyZbKQ5R4NvacHbw+G9lLZpR6U3Zy1ziPg07cSejOE
TeGB3I8cAzuRjO+FVHs9zxAwAZ9QPZs7UDxfG2EV/avC0EcWBd/myVolJ+IYlWi9
VaAfEpl3tFfPkE553vQpQU3CZvm8cnXuuQA/FQ/yeXr4Ic/EyMRqz3LiaNbKJdKd
A5caMz/0HAWFGi6y2GrE1BZZOpBDh2EhM7a7RTCGGaomxW5U6dHIVxnawqJgGNxu
/vGfXSNlLU8AdHQ7TtB8O5aTkVPVzFaLbtooyXl+LJ676XtZuFGHudNbkpIx+vz2
B6gvZlHMmKw4P+T+sO5sbwEbhjXgd5CVVYYBA33+fP6FoT9uzmNHEHTu0yhMYL4h
mCCMh9Aye78rdj7Ad00v3ZGte+847pU8szMcKiGW1BZBKr9h6ueiejzYM6eH/0rZ
aMq/hiYFinaPOqBZ3zPNZ35NPK0wE+MKFO5iGB65o0NjFrxEOz2UjpvZShMfpBpL
q+X8LA9KVWOd+GKrJg3JFUHwhJpJzjZTfwqnmevaMTXUYG4ZbkFcosP/hcbuTVXo
JV2EiztEQ4OmButkySNoRFzfCWrrDXuzQm/HF4ANYIRUllumA0GoM6Wc6pmVFryq
tQTpGJnX76vnBqJG4J5h23e1C1oxPP95DXXqT/DXmsDFyqhmHWkXS2zTQfxTfy67
64gjSuqTZmHlwh6THQfcmOAWe5wkIOlo0TsHCY4qDptcF2fSLDllBC/BXUaQRvUR
LsNmfiRaM9KAaKkxLhQSZ7WLHbqZIT+6HDZnBVLrSIdIvuCsBS41MCOP5UreLSC/
kgAzxyV1HifsiEFgR5l3qLabhc0h4ws0OzmVmYLAopBPHUNMA0TQ5V0f8rFm1kEU
Z6PMSmOJoZUp9u/FYEZokjgK5/d7RdI4rVEmvXZGkuB/LNlTwnq/3PtToo2Ko7my
iN1rYJD7jcopPhC+h+R23pmgPiMWl5Mfzdhd22xIba73JbZ/0rH7/LkOEgbaPTHy
06XymUqTH7LVXhLfzVZfKDCtpKL1GqwUwACd2JPGCq8+pxWVGvTGNCsQhrHaEra1
UJP4/3I90McB1AnYtBbs10DVJfZZv28XVUzYPbFFsCWqJ+obJgqPsgfYlbmL4p/H
TzJGLJiP0cQ3KxY9ayzuKrH7SHthAVA4dmxesbFW1qEK/oHIgnzfJlIO+2IrJ8tl
ZZC92dKL3vMB2wM375e2v+Y+YkGFV2Qp5tO8oWqbm1dW/gZCrlM/JGisT1LsccKh
wSX9V2SxgqJURR2py6tMJ+0wiI3HXBLlP5WM7bcDhGlONIlfl1X+qQ+BzZLGMKVP
EW94n5d5Y+72Vmx4ag297c+zb+69Vvcs9cDQUARvLgkBc2tnJKbcIlvrT/FOF8bH
PEz3+ORX6bh2tEPLFBes9hDAJvILag+uQLnDaWllomWsXeSx+oXVQHa/RyTJNerM
oCxD5pk4SRAzanie/C2wPB4LowQ/dY5pXUPGf4I4MLKDQQ5S58hnbgXRbvCoF3SS
yErphNA0D98vC2BXG+phZy2mm8MZJrEUBTTFFyvNIgKZmxuCfnNN2Pp9XBGCPMbW
7qSEImKg/27oJ2cFBa2SuUfM651HYWkMKoy1Wzvxbis8n9m0zDKA8rITMORXEpAp
EDcd0jhd0f5Eap4ZZf3+XvOEWkL7uRd+lmS5JapWGy06T7Mk9fetXfF2MW9HfZ+j
DUVCrjXtbp6kySFvQjAm0j46JAyPnYSuRqgs1Jp6USwOPiVEJlbuGN37aZutt4Tc
Aovxdy0B7ifJ1/PXpnFBMrPpLj0X7SryKuFFZQcLuWQIv4O0qrTWvy3EQAheRdxl
t8ZaIQn1DYLa+sepfyckSRWvMn6+tvNtDdfTJ5W3H7qJt5+SfaDr7fACWUSOUgQC
cFm5Xbz531ocflK3sgjGp/gwz/R+4JCgxYFEL7sv5Sd5ELWW6d5kQKgQ64gbTTMZ
DUIb+CKMQ+/HYH8eHIDp8KbGew01o3akPi3YDwM33jZKz4JKsleXG3QAXk6wJFNQ
vqPxpMTsCmYNzH0DPb5F691NVemw7Yd//1M7qGuK/H+ovBcfiSYUr/JnlIU51aVy
H4GxSWQuR4piQ+IgsNk6OgCSA5Xtb2RYj4V8CXYsJ9lNoGXyiq1Nl6pSIu/kLyKt
duApA2HeMtOHz0S/64+BqnTzgV0MKyNpTUI7P2mX2T2T+4nDBeYN3+ekEXq0yq7h
/xWec5L+iMTvbxegoYnhg758vdmsTQFlqbwSWiWSw5OeV8SMMRzBMLM+NPc4+6M7
uqSwszxu2trQ5+Y1HOsuKBKWjy+iI4SZrzDC+NPfJzYrb/bMpdzU7SstQ5XXn0FY
d32gCYHDuOAn/w+HbTy5hMHdNw41J5YFVo1WRK4yL68LahMYwio42ZMsP0S5r3ee
37pS7qkNhk11+OSuuaCbo1oBTavtVdVE0irDUy34bl7551eVJoI71NRLhvlsu1FH
dl53P+c+P/rYRBhVTVDhQvjRoPuIdR59up5Ev1N4WIggy2Qag1nKl8hCO9FJ54nB
osWj1xYq1lJ4qQGJ5FMI60ZJ4av/xg13heLEUuzUAiiiW4fjvlDz1apxK7q/d67G
tviJ92SjCYt0GNDsGQkHydLkmF8xNa0xsj1GC17bF5FJ+iz1bu7kEG54YOxeGm0l
Qwykx/BdjcbdHP0CMdH1RuXOPL4oJ1tXb6iucABdErI8uKF09IfhCWPeeZEd4itP
1Sp3Y8JeflTaBgHYVPDDwbrhvSF5UU8japrH2owJp/OWFkWBRur7mjzI6Pxy+9/f
rLZcsZm0r1YUJZ97p28IOlcASebmW8Eh2eIG7a2G9Q/qBMQcnHNlNvsnYL2iqWP6
E1jEWt4Cn5QtAtLakwb9/CpT77iQpwjllIzTQQ/58S4GawQkOdWDgg+V1qtsHdp4
W5z0hoi6x6LZ4uUExn6yKskp+CNOUhFgZat4szC7Augt5K0P2fZjXK/5zxPWweb/
fKSAdxxMMbv0IYxOvS1Pgn0l+8K0AInoCsuRA0D2nq+uko+eCK3YVgNUgvNsQPj/
XanltIPlpJqBsl26pLv1iA5RUen0s+GFvg/QWggRCpCOrFSkI1Ch9vMFHLa8Vivy
S/HBPxfEZMtSbioKg4tIBIq9EOf5mMBs5RTIUjZ2d7CBUoiXuqZJK76i3ww1YEvU
NQGL8e7rGst/qYonYdJCQpENg+4e2EtNqcSjpo47l4N9Cl0gkMtscr9740gXJ5lf
V5XChvjPdy//t2AG+gOWcWTiZt7L2vffsV4b+zjslvb0W1wJBVvQ4mxhhe/FATt7
S0bdBo2gl1GDpz49MrNphKoDWlgXII5+lS1MidjzlZ8oSY8TyWfB5TSNqDRVcPvJ
L6rZ1a6HyZUk+8VVDdbpZ/NZMeXIGLSA0KDaLrmSZxOhF5iC+09WQ7jdxKMKLdug
uYq720HarNj8bTMc5GhbElZqAjsw+bSB6doFlMpQU5FDrbtbj3uRXGTHKSgv43V9
jljSyupbvM1NIu6FUj8Z4yZbA24ThqJ2SjzLSPINxQOQFEV14zU2SIBgv2KsB/xd
zd/OXgsoRecVNqo0meaQtqx7K659G8pRC8ycAnriwGf5+zHTf0sTG24v+s2J1Agn
cFD5+PD6Wx59kO1HQogoyD4QW4cnMSSlnppjyRj9Fsv1QETXaXICBFfEh0taMbfg
m12XPoIcAPCC5+k3UMQXKgd2X+aNYCHhePITsislUETTmanHjhC8Cx55u+Dr+tAb
0Vk7S4JZv6klhIyPlnoebYCl6d7ofo14J8ILSZU6XyaMM824DQTtB5eIu8eXYX1i
FcQuAsY4V7B3YD6G+Avfvt+KDp5RIWUW1VBgGq6aP5ix/JEKNvxVNBQwTFBhTnwe
fGeySadq0N3eNBEFe+53EEM6unIb5bqawAgQSPKSBsTwPo9xXnBm0/BnNjfcfzv6
6WwX5pSaB4DtBR0c77vD3r6o9HN2ROsmcDWlYIvZuNArjjTnUHNyfkZXKwPK16AD
K1JrzD6kF0JMf5rctVoR7UP+UJY4oFpEq+W29GziOo+v4Tr+Nl6DOXAcI9GuKMcg
MHNTflO6WGZ5hjEzKvlPh8BPKq6xeoDD9RJujyIa8WOhV0qURavGM9GGYBvPaOOw
9HmYFWhKAYIT4h4JpUTHPV/AyOuYx0ntWNbEZ9BWMEc8W3f2SA9/ir+9JtM6v9wo
csrfF3mC3Gi2/mZkFHke7CBM8uXqNhxmqfoNteA3339SO3BuLI6WogYAjJ5vvv4H
pDov9n64jr4bnW6eOtJiaWzfdSnQi/oLaiKf0KtreQi4yHkSD4VjrRdsbpJOjeu0
sXt68a6TRuYOFHemfOLYgwW6RGmf/tHVrvPKrg4qjMOLPYka5hSGD59+/6IMc/d6
3IjyD0r3jIdlZnsJtc4KapoPwP3LkCbepCUOeUX589W6LT0P7oyxJn+3mtPFOLi1
rEzoLmuELc/91ktW3MmzrUUWDAaLfq8o3CJxcZiagY961JnDBpV/l3wqmFOzP1IU
bZo4mYlSOmriucVUYhDcMc+mf8DyLLUrP0YKVsteaR+EiCt8ofNzgdltX5TR7h0Y
MpFrgR+C7A/m7ZXKCnrl5wypkq8WLrGFWsYHvRKzkMLe2vTnXNY0JbEA9yM0qDKr
AhwBuekwVqYPJsiJON/1cIUsttEWUdaVK0+p/OMVAQn/RXcSgZ64jyMN7XDGZbGX
miWB/CsOJIS/yGueyIGlIyrUpXKFoMXP+NDceCsDPUDOPp50opkWMV/7FNgp+6AY
ejWjDIL9R7m70Va3TEJ7/ijc+GhYA0q47183aiQRCXbcfmklpzbLG5qwYRvHaY+U
f1TjB2aKkcLjWcQtjRUHFb+uXN8brT6vMyxOAASX1vyS0/UPNqO1jmsD6+i0idoV
bcRf6sDGOAwNm9dDw02sqjHHcaQE7U7p6E+uICV7vUM31fifYum6uP60mIRgxoQp
pk+3VZhrFtWVkhDUebZG93PqW6LD+Rzwo/tHZCSOQBOSjz+FxPLQ1IkFlPfVUq92
mJ3t+OVcHynEnMZLrzq4St5YYUDDd7iymFio7SWcCg1IQoi+n86pdW0+ly/iULk8
gOSD/IaZSSAcEkPgK6h1DSTS077QtxTKv0Apa/fyvIRYXdJqAI+UVeNsqDkwLkD0
q5YetLSjfDiPMe1SjV7+VGFjNd5S7JkRHElauuu+b6x557XoJNkLcEA6Et1A3E08
P/btMawjBufKSvSf4nuVaRdOokrfMehugam+rtuJoU7HeSvLTFIafaubt0r4oPtj
HC71+FLP2B8pb5bDOl2QgCeyqFeztFM48LBwz+CZpXeIEymrleucaLwoSWdAxdEX
6ik5/6K5xisT2b15G/cuNVLtY/2c+c9xYtYR+Dz4ayGx95icRFWOz1A4EJIfy0q1
r8MWgkZQyK1YpclhmYGUbuMQBSfp3hbRrVESuZLerB6RgviyeadSlh6Ywu5qVYa0
Ww6nCHW21OtS+bfn+qS2PpXysn3FXoUj49ZBXezKmHD2PoXhdeYNwZNE5mh3V7HL
FMEvekl/xRcmgzPlZuBSDzF0ijT+pILM3al+wfG+Hpdp3DfJtU4JnaAG8A3Opz/V
ghHBXVdJrWOmtd2nezKljuJVw07/kcuMtCCQssgb6Unc7t6Vi20wO0Xckv2raAMx
PWUYlaGGeUi8Olj5Z1YDifn/qrtO8Ln3UZM19TPP51XPl5tagQrDBm1BuAPA5Dra
B+uvqN9k76K8keYA/U+bYmc9DijjyQM6bwVLF5P1OakKC4qyyKLrVW3s7zuxXL1e
09LAx5NGGFhMFyzSlgYNplicEuRZy4nh7+kAirXStG915TXT85uc1dWiAuIgpUH/
qjLZOTbyr5tXUj5+LzdJekeFozGvPaskSL4Vp74Vq8CFM3PsUZW1RBmVvKRgGpZY
AWDr7wiHyswauGzApgRHLtufKk3BVEejmeRUsl+0jHYbC4u/LtI6qBqE2pCEJpLg
rMvWF4h1VrQ08MfV4r5+qCfCHQBSpiDfjhythiks/ZWsLxC+f0cT1olue04bzEN5
AUGHYoOf1raLqvT7ry3ddyNyyc/YlmI/FMQnvZqFMmTrsRGgN/isca9T+Ch7ToSv
HuM8Sf3nwDorJFH5kXSTZgaJjxLl46zRvXo/SO5tKFZvgZqZqx7qPZUqv12+IVUt
73uGntzrztlTfvUr4EUKyxbEqImXjTEWgDcgTv7ACEzLWAq4el/rUCRBgSUjLY2p
Uj8fMnxJ7YXuhD4ToTeALbNrJiB6DjEhoxb10dgxz1oy4/XInyY5u41m4yYxvQgn
cCv3ZMTb9ZxWj+IQVqDW7AuiUkrS5n6Xln78WZ+FJleqHPNtJibb/xe13brOyjDx
vCgXkLGohzdnvts+IORdmC3O4vcGc6gKgYbGHadzCOhn7VdtiIOP7fsUtz4RJQrx
mMfHhuSo8dB3TJKKfF8bGPvahE7RensC1ehUEpOHI7UfNB9x1OtbmZLjKIthYda4
t9L21mUtohdnf61k2xFMaV0HYfAYJigeBC5xqI9VbLt/uZ9ShaKpHMbJGLcbyp3D
g1NCNZQxv5dLu1uJk799tSgR12PIKscyPYsyUvQqjoX124+d7ICW/Joyf4/O/WuF
mFJqpuP4IaAQljVGb/nK3qbRs6lLuw87TC2J4hcMGPkli0q9ESYqTrG8/J4QrGTp
zjK/vyQ8MwAQTZT4MjrWQ/Oa5w3FUaLa6m+AjVQTDIp+gCOosoM6sxcu506jz8wx
ZeLJhKcB90sLv4XZmJTLYKKg8pF9QAFrKAMHw8SF6meJsCkigFcgGx2q9CgXUi5i
PD1P3dCIYOAh0PhCXsVdorbKxLi5GrelYy7hEcPRDtwWsHOU/i4691o8hqClFVe8
zpyShtPnLWNNRCtrFTPaGc3CRXnwEW+7DsXEBIlp6z8XwZSpdMiHjesW06roGphh
v/sK8Q88SYlINHAUfXNqf+t1Sg5rOFerxqsjE1XqYCfQrrgni9Ds4/8GuJRiEHBo
PcNTyKt+b9eOqlymTiQVHkNI9GtAxWThMLyIxUP3NsxXky8lxtvrjDJ+eFbNFZGN
wYLlcMxpUFLJ/IN87ZgsVK0oCn5KROOicgrjUaOpACe9Jr9iLf1OxPv56JejA0L0
ZjbFrV7mVublgePUbfRcVUENBDHPgsoRLvOF1IypCylDYl1GBEwgnIxZk2lRrevZ
v2zz47pZkpW9SBqsxlKgENJfSreOx1RDcffeg6sSe99FPINbc9xphtEGLwwpNUNZ
/xU0mALac/qYwqsg90nsfHtgrW1Xq5aUwMeQrFGbcCEQsHPYOj7SFUMORFTRbUgL
32qbihWbkVsri6f3F0R1ZMyPRVlDT+rA8zctbZTFxXU0jLFPOPx0AWpnXdYRY7L6
Zg7eOxvAXPtLuI4FhpKuZltV3yQv8srx25qL0poWwobH7JTAWeGcKKhmn/oWPoBA
kI8M0eS3Hk9dw1Nb+8Q/3iR4YXuHN1191GlWCeP4EsdbxX9Sb0oxQcOjmBgBI/pY
znMk+Ub6231E/YhCG2zTygVP1JqnQKFuslN1pYUHP1I1YUFl4C2GubExOJyXIYJn
4pUZS/4YgpVrxJXKzX+/Kvug0ZguwNJYhtRLIEojNDYadsvJd3baay71k9EkC8u4
FkJFan5iYVUQGy8k0xIugcl9+jMIlkntbvKsN99LgK5zKmRtW6jbWm138AW+jlzD
J/rWywUU9qmt9neZMnKYPdKYa4FmrANgZkm7qixH+B32evQix2ivhHwLWMScPM52
Vee7wTWL+AriqBfFH21F3oSqiikStsYVUE7T1RENsEJXIwFKmD+xzzFh4oBER9eH
NhEtHUAInfAevfxGYyev6yUMbmLH6m+lhdWM/E325aTYj1VI75T7w/C0rDM/5JME
cGMXerKREIzMNZqyLqijuaGex7McUr7ydWHwjmUc71l7vVh1Ll+7FNEX/N+D6m6q
6xURD9j4A0dX3wp7bhWjzQUtITLIrJWvBxgs3epauZ83EC55fQiv8N7xRUqXoI/d
b5o4hRsLopPS2OQ3+YrwjSLKJAWPw7SlCX/iascMPNPPosayIUVOGbVfdc1bEdSU
juk3t+zGr218UwQk6eHMDruRpnLo5kFV3xBenGxiAa6elHukAReiiN5oFtI5PtxT
x9L1lRFxMu36XMTScCy0tMtBHNbVLl5K/u0DzWI1XDKK1H5R8RWKzxsIjKJgwU0c
gBxPMwYnByEo5c06tfEJ9LgI/9rjPH2TdgCV3u/q99IkaiBjREbOG//kfvjsF1nO
uNEIU2m6OMEoiYoFvroxG7ehbns0S3t3BqNF44aU3ZVRZg3R0fEQpps/nhOR7qtB
GmMZYpdEqQpqZsxpwJzx2YrdtfNp8RA6JTdtbZa0DVkL3wzYQ7wpl+NJAxFoNtWm
3tUSdy07mBBPp9yEto62jVaT/80NOERJTvXxyVA61+LA62+s54XG3XX0Q7/Way3h
s+6lQWlnE9U55YiXqkvm6VnC1XQNQjhyOdbMl1AD7gbSqbqzpqFnWk95756eL/+/
DW+2fnBwmmCJtDdZbe1rwqJg8zvSdSHYU8VRDMhIMJqIfuIY2WP98vP0GRaMs+Zv
BBkihqTqn335CuhbRs7BFeergi2hjlew23oFHd14IpWBmEGQIhmEYe7wDyMiUH3l
teEmoNcj17JoeY7gN0n/9a4I9gM/pFI9sdk4D6lkPLC7wZioUn2nWarSUl3/s+B4
nIbK2Qoi0Qi1uVnD9BQZa084ScXHCljx0blxrYI2TKvpNr7veJqtn4D9lJLHhxFY
tfoOZ5h007vRbB7Nb+41nh1deyTvdh5EtmTnvaJqJk+qv3y2JQS+aqsN/jhKD2yR
XH7CrZMTfyWmqmPmz2UV+JLcxt6hGAq4wIaxWuuRFKWOJToycU8xmznSyGIV3daw
7FL4T98R/pzNSJNnrbIjriM4rEil/2wZFHnxxwaPDtyRc2ha/WSKCPvvjcNdDZ5V
HWwtZmpeeHEWxK7vNLcNIHNJVyRjISeWcDl5xxJJ2A6PV7GL3IdNZGqmDgLQrjIs
4VAPNFkMA8ql+m/j5TlJQQtSD3g+Gpq6qLI5Qeeu+OKKD7vQFCzXhTAZwU045yGU
VEkxLEIHZwz1a27ugEs97V42XbnDxgNIdAAVYsonkEgAO91tPYbbJIwNpXwI1uuv
hbJhwBi4LR272mXlXJeLQm7OpakYAa6RZDyPUYHstREvVIoI9ZW3GT/Y80q1Qh+B
ctAr6dPBDHpYQJaR5HCIFAXGldxqbwbiBQ+SPLbKFjbAlbLpSUb0ftM2XGbWe2+s
h/Y1JHU2jpE9olZeb8L+xtZ1x1JLccLjl2QcjeF4ixQybH3XdZlQlv+IPzNNEGYR
Av8Rhgve9dDu1hozmzHeklUBMZVZ2Whf70WhAy6ueB4Fs+M6X9HvlLrrprlIjRmR
uc327bGNBNsBo78Qdanuyc6zuBHIoTqU3zh+b78D9HCt/576C0+vr4kaGUy9pwK+
gjgrWJzhEylDLQ788+s643whtVpvQK0Ojof2WUClmKO3TuSR+zlKf0TXhujT733Y
U4ZTVSGfkukzKJClxc/SMtOOsLpd5Iyx9TCp38f2YHMD6xLU66IeSFSVD0WztNbB
OK7gpsDZQrOOhwwAy+uWfP7TSb/Sj7skzvwTI7sIPin5i9CthM9xsszMQ6yk2ci3
SzHB+Xr/cPFkBkqAFWHVIp9pK8j06HozqLlZIXz4n8vp34+ALeXJ5di6wx24Hnco
seXWjYKp1J+7ldqAqxB7U4bVVf/YU4VF/NSkeMtriTx/aVoXek++D1mVhTtoAucO
cyJmaNZBAU3tuUV0pAyDdZSbP7zhzKPyNrfioor80nyPX4hBrF2GCGLh3y8LyL9Z
cWKmua0rW2v/mhiTllytzM3GpB3v45oUTlx9rQVTDlaNqoV/Ip5wUTZR98OBKsnP
49BUYn0U+ns+us97HHuZKICaNX2OAd/aXeC+gDa6TkrPGfvE30sR9hCDD0pDLolG
1FrF3NlSxdCRAu6SYtmTMZutAWlTPYie/maUQLjolNM8q0UWCfNcXvJZcGFEBWpD
nJk93hZcLTZySA7A+UWvU/87rNp7Db/ZQjbkGVvoDJKEwNDYT20LeB8bzd2Bmnra
bU1DC86unxOSB2SDrX5011EKV4TvMc5iid13ZuGfGoj8uKjp6mRp5yk6i+4e9jmZ
OPkJtIUU0uiMpkFL47QxJgRDrWm1u6TqnYtSLsKm4DopY57Jui2CWG/PWdJuL++M
LdDSFAjENx61o1gbGd762GYLYw6TcVCa3Ix6+WGQtnvvzUIiriMXK27Xa5bQC8x+
KzVSiUiOSMtXn8dgkna7dPXy80yS0i87MDsVcfHrIpoYzfjeAhA1w2CpunedmBN/
nEZlLDmu/7tkaEFGBhaL/aFQ37bOJuYoPNo3tv+OMdBPIyjQcFB1qJ0GdRLFZcj7
CNh3/bgbsmy+lAyLzV8u0frG8eoi8k6eC9ICMcQ2e5mBu/qUOKXhT0ANsMuv3F9T
3DsaY2TkSPaHVsqgW+E/pIJCyi5Gq/JvpFxQ7A7m6zSFWPgxMasJZ13vgY5PEq13
CIJ8AhDbXlmJgdmPNjk43QZqRLnssS7Ea2virVOwb2jOAdzY1dGkLf2dxGJEdCQB
Q/vrhcZZAnMoVMGKMRSJ4o+jpLhrlgkY4bQ1SyMK6h1AhSbHntdDeXxm1nV85pPM
E0T8kEQoa7/OYxxT5zmaXecpVZus5bf8vxN2jgxNEWOcIKwBnQeiKrCFlWgu0HoZ
W6oCl7tQobI+yurAQKfMX857Ym/N0dM90Ex31yUXmvMLAgc4bbZvaqfUaS6Uts6w
WjGzEogT2ODYiOVRGFP82KHXQF01SBhkojq/BhoeaAMIsnUshO5K4PWtYXM4a+S7
EO+GxotvhI5+cGGNu+X8X99Z1DY0p5q5pev3/Wgxe89sv4b3tWmm98GEEhbgoMC2
4wzqsTbmQNjSberhDRwGK+1Gh+2Rbrn8czLdpHRixalo2ilzvwpqyN8ev5z0Zj8A
kfwYQizeNw/nV8JSXkOx3IOmlMrUIQ+w6ArIJ7usLk2f+omC9lF6BklBSgEqEAT3
2bTvFH5689Xshcz8ixViy66lr2JgxKGmaZI0FrqOcPsFwPwJvq8ZOzEVS9NFXO3f
km+vfLF4cOpUkhD1PnqLudQRRLwtz+CPXRF4ZMtHuyI08ZWcRX8oZVoFkl+JI2FB
enKqowDcObfcWoZjXs5BZw1k1Zly3eg2YGyLSOAqz+f8YBerhg9Qml8ie9oDz2OD
s76ANwg4kZfJXqAHhhijlQjt+D4iEWuHZe2qpdyf5dLe3ydNyZSsF26xW7fu5LnO
E0zomTwne6+bC8NghD171AqjFja58Zlbq76fbsiZtXufkhpCcGe1o1wpvso/XF3R
i7FvHJB+05MmX3XfHu3SWZORXHR4x1eroS/aIqoYxekMoX5KIHJBuTS0l3kbs6kx
GdTgglhMCecHvbZpfKI6K4GpsLgzGwp2LK3ACNuw4HbErFyJBdJUM3RcR6skStLq
viGfn3Gxj1LG2mNua1wWOO5BOvpfvFAIkRmqIBuDRPIbYLQqgQTlSvbb+qn10ty3
EtiLV/iggvsfYAONp4IIejUCA+aeZweLk6uvEHeDYZs18okcQJPMg5Cm8PU9ldCn
TF08ZnUWM79RqbyoxtU36NJn3KJetPo4VmSmM2U7GjsXHzUfCk9B1Pp9+ZajXisT
i5ECp10Ubhc9RghMl/1+JcroL27wvkoO6at/cpiMDk4i0/1RW0X9JTvAcYaLomx0
bO8yWj/kPTNwp4ziPtGP+NlJWpAw36fcd/EUx3rTey9mrVcayjHH/sh9GNrFvFWa
bQ55mgTemYfp/z1PZs90Of+ygwcKXQG3cCgfNbCXWA7qfIj8CsxIcRpL6exybE0N
twE1CRN9RMpTCf9z4IhouiFgkLE/RJ3IXVQFxn7VyH2U1YeSEpcRgYyMBF/swOYP
1pdSLVBIKhyx/r1VoJeyP2u2QSa3/BNfb+P6JR0njC0EqndyLjKZAvLJ4LCwXdl1
6YX4a7o3rfju0xKb5TpXxrGXA1EFluwvSZTvOenlHDF2EFKY+9MRA3NzH6/dHAGW
mr/O3PFOfGg4KaJ8Ftbsf/5lJGyiQtoUfzwVInlShf77EMuq7QP7r5uQTpiopCun
L7fTOIxNdrq2RFGzoVezsgPThyGgf50K9qKEKEfhYlAbpdRIG9PKgF7OzyYnSNAr
paCO+arcYz9bg/YQaSANI9p0ohGPCDNcPW+BJfrTYB6sPhXYt4U+DcsWxVo+U8P+
tTAad2QQSyz5hUCqUh1R0RCRSw2cpNMHxQWsccIjtWpbERNxNpjs4U399xFUhzEA
mcWT9PSQqHjns7le/xGEmo1PaOwR5D3IGJkxX4o9kGE7pEXI300Cp7VFJrTWeT8r
b1iMLy7e2UZaSEfYmT0i8Sn7xbc22jZGm9O95hvM+f5y1dcFG0yxtCpTLhimRu0/
M5fIxm58TfuNVYUfQWhcO5Ig4ZHhKC+f+Y0prPqiEbWR4CIxlKUzelQUzKT8BrXg
Ue+JKhd3oaIZwddEnKH4zCewi3b/l6eBASbSgfBYHoSUeT/xoWTNcQjsTA9hzFzO
SFQW6wDohpIeu4F8vLrDXKywURFCmODC2Sc8K78VUH5trxWMIsXsTdCf78Ts6Dz4
SSUMP4UYpGhID/dFvOoIAb3rkhLNJy5KJhttxW5LT3WtPezM0MmIkbC6nhbAnvIy
cDysFrdXxFxRzlWKOtI1uBIuhJKYhEvfFtuUDltGEMFm/LF7nGCFTw2NB/06gHuv
p5LMxpOW84zugGGpE6HoI3mTqcVU0anZu/pWlvmwNZvub5kFwFor5DD4FCwng/LX
QjLZ3U7lq97Y6qbQIh9qUeYd7HNnPhW5Dt4IDZKPU6El+8jW7A+X/oiPMCDFSey8
LCBALb2MOq2Tzf7fOo8aB1LMJ/woBhsrZyYd7YeB1nktaiAuk9HIc7MxJ0S0qkik
DCMY+UKARKaV9yGVJELdj5kXgxCTQUHn/ObtZbl2dEsrdgSeJC/kX+fm8M5QcjN+
bfvkz5wEpYCEtZOlHRI7BRZHMFIWEsbegCER6JQjTSghUKchgaz274hrAIXIdYST
StG+/3WKxhCrbjOgOa++8HGo5TrwQJNL8qLpJechwzN3VE1/nrO6qRZVGR02/+um
Vr/C+9gMEsARMmOm3kfO+lh8Oy4ZSqzWd/ZM7FBCqO4Of+VdG7+4puErsWAAGo7/
VfuqHPDn9vyuMqpwzPZ9zWD8lejcx7YqnfQ+Sh/NH+0/zAZflUpF+CU5lTO8vRoh
JXIM9EYyGr0U1f0KWEnmFJDvV5xdPDBERKAyg6lUgps0I3vqQLKhYOFKj7QpINn/
JCaE7vXw8fXFWybGgRS3SlFvfoSByO4CWUjpudo+WLVi0mSCz4WIba5InJ3hg+WQ
EZqpkieRGNpddNYFs2Y+4Wkoh0IoWs+NH4vymGJq583Z83aJNMOS/xJlOCrBs9JS
sDLLnmpXYG72JxxFw9NqgwcLib6p32Rozpb2zZl0egIl0PkTI7mTM6+AkJoT8aS8
zGlCc1vzxJQhE+HaEdTAqSkgJwYzNdsaLRtxSPvLkeEGmTMA3zcST/IhKtgLDJdT
8uaXu0dk2n0WJRniMAafD+ONYAjfE/dLW4b20Xr2fDH/j9prVfIkl7ThqZ7t4DNm
1VlgslMiG+Zlq/RMfeFOSPq5OiuGPMxHuY9Mg1E61MWjvKgYRbTxKKhGojeypPTT
raKsbHN2O5dMl+XOr630XvoLC0pihTFdJf0Mbf5NTnYe4ecQPOuqzWQj4SIXO1ry
rsTBRPBCrAr/lOmiueh2u6i9CFR0IAmvg4RA3UnpNtH27MCKRRpinb//MX6UtDPV
PMbuSu59dSsCytofCRK4D8C1zl+zjfJWSnthPkQksUmRnX/pVk73iRraqJIuXZag
W7T4hX9T+B+RTICkufk4IJB0f9FieYYLufOZg75HRjhrBUPTBABPOsSMYVIJbp/G
OyKsaqZ4IhKsj7pWoB1J2dxHboWkLBAagy1g4uWWMNhY+QQdn/AdvEtVxZTiEXuY
KRHKgn8so7ALEJMFcmhm9xIpEpfDkKe6HucfC/jmXNgzxazvWraAfC2INxxThF8h
6guVtviF0gC3ifBhUXXVt6Qp2MDXSHfBhOQMbQZ5QYQumEP5Y1RyCi83kLGL4I3c
X1VT7gVV69XFoJnofcJf4cHD3iC9J9dqp3TBIY6dojOhdNBenryBOT16qdq+zfQN
ZyrS36Ez7ROw3wu9GWpjveLNit5u/a2v+03Mz0T+Ql4MI2163WBN7jjZIXrKTQ4j
24A1SQzYMpDLpywoTn3GOLM7lrGNCfdQdeW3wqVa/f7qE+UnFdmUglxzPd/BUauX
98ZRIBLKezH2hyWXaPBv/1Q24I8uWbCShvxmFotmufMw1B0dK8r9UVr/vS4QxSZY
C6ksIo+nwLY8Jh6LnH5dKGNLaPh0aehrzGsiw3xOFoXVPtNcSRlzAhi19USJZjdX
0RC3SP4hDldWNwCI6JVokWLJ49lhbw+H7x70iQ/o7FBrAQD1ocQatlBNLueuv4lu
qFkrx4INGm8MH3c+7flikRGqWqa6OuPW2cFPJSQmKFzckz4dCBsbILg4In03/OjP
bIiRjTeWW8++SPBH2E/wlVWkYQevoILGVmQlrWMY1ynUOz0BMj3bjyxt5NHUuKpF
zqe8hnbxWxKetYSDyGfcXlNLgPsQYBKMgU4M1mRY8n7h1TtxS0Ywf92S1pMy9e5f
qtYiV19HQmyocd8IApINaTel+5XF69XnbePP2O8BV64O0AucCkcM7M/QUMvJCEe8
P8iqWbLwALpnhzFEPMzqor13d3ZZjYOuWPeE/WTxyHXdZAOKkZAfdXjRH/Hzkx2v
3GlzvIjf+3vHgCMBhjD5lavpSgzpWdxGxaWhA3XJqvinE+oiD4ZarFE310c7llii
TtWlL2XJKRb4qEKSCnq+dERJ/B2YBDSujV5yDsFHJfGyTYsY92NPAKfS6fa+rmY3
qtoSQfCKiZWAdKNFSEPZQtUNP/YWLQ8c8gfdR1hINwjsT0iUgQ/t6bDT0VIWSvI/
VzK2/xLeDp9c989vlXMEHv4FSQn0wcYZ6wWdebRWdUYAcCcUqCzBmqWMH0npSqhp
nQm7uZgOeNQx6p9CUav2bT/ZBfh/CrPnfa98qrVEwoQC4+PqMhZX0ayCtiWDEBu8
EjWFCWrD6TqidrKSyijb3ocAGNDsdLt/Fu7UZMQChuutlGFYQhpOp8WoqfF4kGYD
FjbH6H9sMrArOfMa4RpaNrN9zo+WMRZFfWJ84okWYQ0H5s+zxwmX3+e1wRgJ1FEY
Eah4nvtFiRo9xM3L8Mfbb6uONuvi9Yd126QLvtC8xIhDkSuDWTp4zMlMS0f+0YlU
GVkBMXVS1vQ4Dsi0UjU6RvCThmfjXoHLdo98Z8d7FHGn42mN2IyXCE80w/+vjNic
jFJ/hJx1r7vYd5qLGJTuq3tLiwT3eKOv/qjXxXzN+HYmeYhJbYA2Kliviai2aw9d
WGWFEVV4nJOFRTemAa/MIUNjPGs+vrFLhUyWhY3bugh52sjJoDs3mBJAE8C9ei7x
5gUbxCEVxJCNQptxj0uUafC3t1/4F5uD7Z0PA8FWZLBAsTIOx14uYCyWZ+WjRpU7
wrku8KHy1rHRx8g1XGrEk8h4icgK+ySJgJ4bYyPbtFYHpMRrQ7B2/lEkSy2w4Hl0
vIfhLAGgCV6a9DL/0A9hRnm5gaN4RC6IZ2fWq4V9Yn95xWZb8Tw8iaVaxhnQMj+C
C+jHaFZNsDy00TKYRHMhKnff+TgmBLUZGCQsZnwf+ZSuaMO4CV7NpeqftmjffTCU
X7Dcu31vvz60Br1hgWxDbmWVq46OAzLuTP0MmBKql5nPNuLKVU/QfHBoP5gguMWS
DLLWiA8guz685yOfbsmWT93/LPGFaXPzdnGDbxbjUJ3HgbzEmcxBDrXnINEOl7DJ
/P5lz2FBclti4ZMFzOxGHa8OLpmT2sB6qTcjC1LNbdFLfTQSdwLdZzNSQiu32B4S
sm4+VXgjSZ6jYRteD9KOGbj3ac4jqNTw9Gx7yrkfs5p9OY1P5M1ngCbhkv+TiNdK
rHndITKf0hkml8os4M5OFkW49p4do6DrqX0+pGu5xPbJs4N/Cy3Lse3+0DTb/4Z+
bVlsX8ngqFsKOj5f4Tynn+5bV3CntTct3R/db27JFO3PXkzHgNIuktFqseoyh9BV
u8FXZdyGJIWcxClB00+rLvlPfqkPMYOc/9v9i1FdBvh45xYJVsMJ9Eyfd63v2DIg
4sGSs/UwjJ2r1tH9kyB/rrBw5hQ8iqGJg0Z10BOoBMXivI1OyjrEqVHW91SgH1iw
qCHyzY+jPl5X+ehF57h2YV2Xt/LGx07pOZgwld3bxUw2rlWibsT0AbDcuHMtJ6SG
zitv6GDZM5cQ2YX/puHYjjZIkPwVBc5ny47EwsCaATGctr7wivsYSkYXbWbzqE0h
LGm2jAql75+Gk/HgHX2e4q7RyU/K9+mm7ITVWtZcLKy/htwC647l7TrohWeSaZsg
X4r8+m6oETtb5Mlq/aqcqoavkVDd80+snNyZJ1LoYae+N9N3keWS8eXkcUo2G0fk
zh36LanbsGK6rf0NkUGDDO1cHNRWoZMez9rshak6dp+RAprbnxf78hlcjXMg/3UE
so7hJ0DyXVb3sMfhBDYOF4kM4/coxbLoCtqvB8qTFaB5bqNhOjtSVgsudiuymcVi
NpMyVXP+lYJ0ERL2AE4YcvY9ONrpakHC1ze4diAaqlB8xdfeE5Ur6zo2qz1XRXlD
Cu5ou4Kf7eJqaRwW1nzlp4EgCAh2sbWeErmDtAubJL2zmK0EyOx2pBRnrlpQjHka
0Yqsa0rBWlyJx2fq8DbaIChVaUd6aisCd1idfkUH10T5GdlkH0pLWBA9w7QgqCSa
9YkUwFm7XRCXLXY6Wf5/19dCjXmNpUUBqelHUqGBFvI3b99AZR0nvOTl8fvU9akd
E533fAYlU9XwipNb97ryF9Cf5pNkP9MGmDhu4DHbUVbeOrYMvyXMrFadHHgkBdxG
kFY48JPR+20Bubq8yfsb/07EQztvTFqg1857feQnNxtAhiiSuBXbR+IVtNdt4lk4
TbtkI1T68J+kaSgFmbKI5nBWzBjOapue9GJ9ELuyGxbTDzb+fDnbAraCoxXQrA9Z
79MSjKpHO11UXNRLQTZb193nAaE4O2hzjQtbGeJPRdlvM7o9rPGNsgFmYkERFsks
M05Tv2ltImvErEs+5AKQXF/+Dih57Ue/51CzxP5vyZshh0w5wH6TTGG+aUEb8SV3
jyZgmQSAXSN6EhpBV0aPdaBPU5sLJbELEyWYO+Or1dxMb7VtQU7fizda6LUq+yse
l347DSV0YcQYBTNQPcjUmb7uO7beqHe+sA5Wgi6G+nYxXS8t5ZudLXPhPImUqTAH
B55BRjmHOiKglNBWSeAaqPhap5a6G5iCTxbjTe/TAW2hh5W9uaHjl7oM+8joyLvN
kT7w9MoNpjYGjFTgBZXcKqS5gWqD1ONbLhguxbF079lTmnnxZisQsk2h+RwgcoZE
onG/51qSh59lPsM1xgK2em/6R1VjqmbvhJ0sUIZDSgSEfYiTya1HwBunQk7gi9wh
ASw4gbRTKafgDtVY6szT6BKFQt/OCheY4H/zxrDrCS/WOCkrMtE9iYqX0woNQHy0
eV2+dlb7RPpJKyi0Y4qO56gI2jhfc5NnWzpq0BXIdeasw0GW3JV6MgLDgPfZOEy6
NiEW4a/idrlFMJ59Nc695Z9CWJL5bR8ataZtFVXQdOmljcw4HQ0WHrOuEavNXUKC
eCB5fHjvHXFn4XeOLnKFkMSsftMuXDyeZSgL723iB31fwAY47l1+qx3m000KIt5k
oG39k0Li/2kXqU26GoeO8tGnWxvoOguD8kISbKx30sUwdfEp1DTV/IrR9732koCp
UPGH7nmnCwrPHtMbgp5qxtIfUUOMo++fsy1PGr9i5n4xRMeu1c65HuA9n0O2KhHa
N1GXQs0SXNiYyVuVCnyf1zkMWYZWobdnbOTEPlZadAvg6r4PHDr162NlxeHZvlPd
SzzCKQBcdIGnSz0xhjxtm0dYEgWEw0O1fl/2t8S2r5Cb2m6U+LBe7sXxqmQBQ9hZ
tNvMgOHFGbVbBcW7IojwyCm5RtQwlbR3nYHa1ZsfKBErnOlyY9DUK6y/Hcv3sjcs
UUF/pKgafbtf6Pcd2JP4Ewr3nD1/rrnyhE9+FmRrCQbbUx6L4PMbNd38Z1g9o1/r
sfQnFjz17pXGXfYC9ZRlA3M8Za+59S1hE/5bvN0mBd+CDNHOlLdBzbgpOQfrCZ1i
6yJeE3oBGYO7Hzhak5AhcYWgfhhVOqf7c/MpA4WWtwwO8T/uaHr2hwW3tdqpxIHs
86NBuE5UutWp5aOmu/5EfAjHhohcQCTz23yezra71XMrOJHpVb4RsyWf06IMiYNB
lrQ+jzuGffMn267ctzOoCoiMGTmPqMBUHvQhY3aBUpn9ngTCfiRVayxr/wCwSVgw
lRWBdGMirfzDlUrhi0aFdviYW2y/gpd71NT8FVQat+r2oiCvG1zXJyr2RtVH86iR
PDCHMkUtgM4UAID49IDHq4Q0dBdZCZSWqqE6fZmKzbVRbEFraOSPcN7/OpQ1g1HF
c6gCoHxQfdbn/9pfiG8Bblyy1yijNA+J5iZthvqkQsIFRnUgmkg8HQ7+An/3DeBz
U4qWwZxWy/KwQiauJ3D42u/o47nl6roiTpM3+Q5MqNJ2nQn7+fbJxji3BMc58R2F
aDKPGlMoCvFzqnAe9crVMTi8WtZvZ84usIVrLZewkSM8WhuyvBNTCJphP7T33ipi
lfdsdeTV+gjwRTABu2q/JUCIm4ZaEoZXd5T4pP4PJW2bLexkJM3zzRgpB1B+cxmb
ktaDzSbfhMgW9gAyGkRnzQz8692qvBqXqV9hKXx5Zjj8SuH2xk/Iz48ojqv0iS6l
pkNLXWc0F47SPb8xDx1elAU+uAmieob44CVvpOMkoF3M1+/ScYTHzP1XRHjnz5V8
QgjWx+Apq8pIAoN85s4wJbb0oyIUR46x/aEgXIAeu0j//2xbaSN8vjqarTsc18ZS
rm8aJ6BIFoKTnIzZQGtM+PtTAJfU4XppDxNzz8lLrFCTT+HXs530whyn/mnqwZIl
kJ80cLYHvAehKOKZ4yOFsFN49q6qL9Uyq0Nk4LQxXe4YwV5tzjfpQkJKsgFhEVsY
wfxN5KryuH8Ypuln3CRzBLNCjFvt2W4hVX5EPtSBEm17FrrVZ/asRuffdtiW1q66
qOYIeX5KMgzpmhN9fhtLPbVlJ3q/gRgU/fbYlSmyh3q1Rx2S3O8sByfNslDyeB3T
fLxSuCktYq96HT3EXrUeEzeMBKl2JF/f2Q2okRW1VZ2R0qeBXk8hJoogzFTSgWk5
v27EIGe+1a3OnNpsD/vEczUk8lH9L/LV0vfZ8SkpxO13Ib0ChAF963tVNxzgQpJh
aeP0H0HFWzEZgjO1hYBdR4BnCSAwuJWvf6oEZSnwW8ng/5VDyWaNRUI3aq297sUD
rfeOBFS4FaXEFZ8KS4rT7z6LR++zrKMwd1y0fEdhpm76PsLLg53UMEuN7C7hU6wr
5P/+eaS/MSeDt/Zxwzym2gDYLMWY8nbZa5KQ3WftJM23DplfM82BQL86UqkrGyQK
kE7gCzD8kbtPT26JCFu9N2HVX4u+w/Cw7l5gNj/epsEJ3l+PP9i8hU9tsNjbI6qB
hZFJacNpw08YYNI/i67N7KPzxocvYLHVv/s6CFoJ+BcpDzCeRNK2rhXotvuA34Vv
tNScO637vhQ48R9Hfa2g8C615c6HzuetBaWfsN1T9rzG9jkUkmQ8lnPLin4Gp7e1
EzuhCSzmoYKoaeE5OiLNSqEYfLeOGZF3Iy/RzBfLTayxcmIC8Dwm1sKS33ZWFlwy
ApGNKhMprlxEdn+Kww1cTDSMp7h4B7WeDAATDK5jW0UGv6LkmcLkmHr0aeb0LWlh
vMrYStucRES+prnbVdtXmeogAmp920hmoEhxNvMGfm2kzoP4zjklHIwefAIjIsPd
5mKqze0A/4mnQNt/E4HgSsZV19adjd19TurvB2FZndzXdKvI3B3W9BXSCMhQF9zm
jHM4wg66jHBRbI07C5V2ZMVAIVKkDazcJkyElnqShuSBjLwWidKAHHS+tFlonRRg
DN1p8a6Z4Vhf/er1ZGoamWCqlKYcYRls5KRlCtzu3HSoow4pabye3aoZfpMBeYN4
Lg8996m9DBvnBcSU/tBxvO1GbLDOiioXuEmgDWTG4fkY2e1RekfwW3JmWUuyK10A
jE1Rd24qkz179Oj+0MDdeEGc2nA2Z3NWd4imZXlJ7HxxY3/E/D1wN/Gls5oZJsEa
rbEWOgApJeELWNIMwyJt7uYFeq62oMkMHltZt4fK0W8pbXeraY9SzX2yRfELmRzo
PxugNQitwPV6oJ3mVhJQiDxsVmwbU2G0MNT2PTLMu5zww0Kx2alpBZwbGnqExnUk
maM+qzE+/nYj9zWpkTmyVjtTFVy1I0aCEGgGkR5Xo/9TFNfQtYE5tCsm869mL0uX
eGqruRYYTbDQnjfhPhjhZIHolZNWxG8/iOhV6zqAwRa7jR9es7GFo6mNrGlyZUhC
oeOWdsfgB9oP/xO8qDuU1zF93fSKKAvGqZL1mUApFLAjXjOakpjBhBIOaoUTQOHN
rQJe12ahV5ik+QOrZi3MGyhC34Y3rWUFhR5aqWnv5dqYGBnHJ5Yk8mwUr2uyZ2FH
5sAIXUZWD7WmfGf6ANJm3WmfwppRwI6BGX/yJ58wnC8sakfhNPJrVnwKfOez+upe
mscAdo/75HvJSUPp4rxLjZQ/HtFn8nN1rXHinPotsXHnkQoY8RAxJ8PKXjQXgjEP
cSFcRDj6dKNhHZa74+RJ6RRO1SHoyOFR6mCgMXPaZtSmCRH8MpFzTxozEXRmoWdp
lvj5aNEUWkhGnvj8TFEzVSqiiGr17PDb3tE8z43Jbv6qClbup0w9+VesDsiFXgyO
4G3lPQJpPf6vBZV9xnMPGeCe8Huq+NMhiAvL7tmZYnPAl8/kaUdSXvpkkgbaKY4L
pFsgVo2vZVhtTdBoqFdBdcsuQ7Z1xbXYLMaBc078nfV9tFS+XqgT8+21YhWZxKO/
65ox0Ydr/eG8AHMt5dls0EII5tDOmnZC2ah/eG/8tXO7WU5r5EjWWMagCwnCqpFu
V95/fax5O5Ex90NS6Q5xJNnbNL4EH56gvSKqgU+1Jk6Ve2xw99TNYc17FTCwl+Kt
ONr2a72nfLpVZFtIZCGrxEZuzjsuOQ6pCTtpQiJ0U88k/5jZlaiDgDFoy/33hw7y
jwPQ8nCPLdciz+o5NVeuQreVm3PFIco29Rg7L50I0uxtTQc82nLqgutjUOPcO/SO
M/nRKamBZ2u9fqw70lzA1fFoQ2jMtMYQOX1yNxJRwSLZ2T6vZKk/wsPYtQypDISr
7QMc3LT1Tg0lTvF6p4qak7HvoSSiw9L0JoosicpzepvO/0jipLmbgdzqvhsDEWEL
SVm9ERVyVDWd+e8fh2LiU4j/l+icv4NaBxATqXD6aGxgyZOppzt5eeSFx7RxZJKe
C7T3YoAx0j4qH8DWHtf46VBWHDWhKZBQjtEmCP/LvUipMXk3gCxySpovjppooE0X
YYkd9CHa6oFu8p8xZ2zvIJUQxf1p52EShuZB9iiF5N3KTTr8Od0ScMwNZ8Lki1Be
dy25ztC0DNm7hwFe4DHVwIY1OATbv47gJjYOPijTZsMny5/YCukPoKa/rpKrrO8x
jGCB92j/+ijdncgitESvA1lu5CZ+NSRbY7bm3fGbifr2rNPpqgFJ1O956i+VrZdh
XtKx9j0Z/ZKAb3+0yODI5V3aAiZJhUmtY5U8Sm4yKehcnNSD031MoTIiPuB45Lvu
nlXIOOoECh9hJ+DY5+FkIqxgGsjw3FvUqwspqHRevZ5dR6b3kFjKecApvMkbm30q
pVM4oEXkuqd25UhfBzz4pcaBNo1cA/sIjnJCRROLdmqNl9gu+f0Vvv4FhDmKYKxr
IDi5uMjsEHwHPC88ZPTy4iSk29C/yfyD/NZHya8e1jcooeqXkx5eSNrG977m58b7
okINsMMPlRAQuVCAqGpVZKT1FgKzi+GYwHyEuBOJaKdqGQsfrWy+qrRpk0P6T10A
oTbQRWkXWqwLgvm0IV6cnKiCMXcH//VYJ0dCsTpuAh/LBrbQi1zmmh38PkFL0Vqh
HhU2uPNSFQoguRDk6r3OaHIWYhC6Eitb62q7oMzB+eRDiszhFcCSzVL2s8nD65MH
pi9gKVULt/qXOg9WzVq5eImDSohtMgLDj79YwRj4N0rtJYdRxPnKBpeoFLgKG6c/
z5YVypoiB2RSietynRC1yrHEUkSxCJPakSZdyZbp97Rh61y/6BwTYqJKQ9liAdAn
v2qT4XE6IH+XaBA9AeOXpy3iQO8W4X14cu/n4kxQXBAasJPjDCfmoce0lBDAU8zT
svECqfVsRZxIk8PHRfqdyrT7da7Fk0GXcGCJARo95E7AgQjKOrRKw7n+J0j1r5DH
++UZv7c3h/pLU2NFn516KmPjTcS301LXU4jIrcsD26mol3Qct9h4Lqt0StpqELZj
ttMNByqW6jvUSuqswoBVBJ1Si8VFFnmWWWx4xupT1PKhY5sqffu44KnXrCZ0K6qV
01A/9q+9bXHaogsf51jZrrsWDRuHNw9ygnaUW9qWZyQolfzSnJhnJI46XHjQFtU/
mQHa1UnKcbyaphoE0BCwVlQ9NocdXbGA2xUd6X2QDZUcDQzN4mU+1eeo/NNRd8z6
BiEWjfK18Dvfbj39H161BNHt8pRzXfup14tpT9LKAjNH8tuSiusL0kyZaePc9Zqa
CUb67igCSCZQSxj9BLgzE7lc6u6KAg9GCeDA/7FKaKD7wPQ/VRXcCEFOPgOryUPp
+eu1dGAYsW6UL0wBGdJiphbnnimLAh4vMyH0e3mmFDacSQOjD5VRu7FnPUo96fom
DuywaRqwX0qU1JL4fnqWyOSadbwsKTXvYQW5NMaE/prTKQwpFnkOQj3nPEH721oZ
XOaJg/uBwl4tzt4kmdaeH4eECtMBhLtQiJe3iPzzCm9iOj0smOvAsIk1JNPM/J4O
XnrXWCCXzq0PbXbr6wUm08tvwORM5cmXtJZRy2jftQOYKYaGGXPCA3my2X2u2M2K
ufLbaQDb3LSMqkwVvwbHdPbH3u4RnQ5gQKVOM5t7WLi1eNbGC6FqJ4WuabI/0JEw
w5SX0W6zv2DEyfZlnvoULEQ+qFil7atcyPw+Lfqh3N2Jg8qKMH+T3swzR3gpb3eX
Q8wXrAyUbkMOAkDy3WqEWlUYU7lBYc8q8/sD0Q/wReJXBovLzsYhoC2bDoQ8xryn
JuOgDI7ItoTfCHkOMuoluzdt6zu9+JuWtZv6zd3BXzueNGqoauxoaSVunNroKQI+
Z0DK4tXWXRAXkJiJ8LCjxKIL1G/p6pMTvr0LRbygSurErIMgE+9gZ4FdCYTsI2Vc
luG7o9ekJS8hlB1vLZPn2/52jIGen307TJmXFfBjSzhvz+GivQhbhNEZfi81h0sX
oUOCi6Va2QMkUlhjcxSpZpjDspf2rluK/78z8t0qkhgJ6oEoaCI6dcb97He0dolV
cRlbyGDVGTjhJ+VgCk3EWJhbATyrBmzLkeHVlajamY6kQ/CHvwVSUi6wicQbn0Uy
NYYQ2R30O0ju2gTMecqw4lyxy4YEEhsRlSVk0IFGTsMhYjQP6IQOX6rVs4IEFE5+
n/goJQzcgTfmb6HtbhYB1mSFIhIfHbhNi/XiVXmO9FiIEt40y0u8Ygjg25hzc6Xc
D5tJWIbck+P/QkXG96qM0igHYxgJYXlc/eiEYfu3iAiRtSS1Ga9RAmquKNcL0dMV
a29Uh8eVlQd/n9z/J42AnCfKXbly0IKyzHHn+JXNS6gMhMrJ1KbGUsTAD2xgp+qP
qoDmGM6/LAOIfIGapxZKQ6DbsPK3ECoAEgSFKLdcdTt61hUNc4ktMZQME+FUjHoq
RoOVfoGW+qrLf6Fp/xqjdVpp3w+VWU/Itj9TrtZJvlYLF1BC3QNlu0sqTIVicG6t
ToNRSBaIAbg0A0zMweyjYlF+u1mnTwyDuc3iuID19dpbcu9yI2VZ9EBUjVkotr5T
OjugJSUUIyxHOoFJPWyLMPrx+CpKxpHSeVxbK42PgcnemW1RjBPBNeiCtoanM/EW
S7nA8tefcUMSAiOfPlWll4iC6F0kwjhgyfCkhAZUe0E=
//pragma protect end_data_block
//pragma protect digest_block
uxLzm22kwbdAyOn0Gy1yTBmoqGg=
//pragma protect end_digest_block
//pragma protect end_protected
