// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
HQN4sPPFI4q+afiblSGQfJSp84Yn21IB4K7c1Owd8P72P0+8teKcd4TUq69ykbHY
SSiCQLtPisbIRj41END6+VGhVfbpMWrhXLJTA1k3P6JoKOgT1X+jlI81tRVaL1+T
hVtTfDZmqsf3Oq0TSzWieBpFEUDFWgbtWKKxVthXYGE=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 5472 )
`pragma protect data_block
0eZ2oRjtv489tuzQdYm0ruvHsjCyqe7KFSWQsduqxng6r4HDYKJs0QqOmpJ3w0Z1
su73q9QSJAvh4xbtwbPxpt1DmNJBtQCE4dY/gS1IvOJ0boIgER0E30Xl3CEZ2QIb
Zh34P+Y7KxRGyxWeunrfx7GIvJdRGpqgvhLWbd3NJLLOJbesAUbfINItH5417Gfy
NwLVwBMK1l/LXAkqNQVVeCHG5XlfuPYRSvXz2mz3W7i9ClJPknU1TnUON1LVZ6Ev
Ae2HFZkRQGP7NHaqVP/f/dlu6cwShdIn5E88oFsDi7oIAUUwLuTWgBKevwxTGz5U
AOjE1yGWrhU3TqtGmWQnFRlPLvbyBOkrHcv5h41zFfvWdBqPGk+1igBuERn4Mcyz
pEOK6Ia/sdQQXEhCpJ1ZXsYlmEKTaC51/8T5UiKCDmv3VApCA9+dq9rW3mqq52nt
UVwzOuJvn0yyDBOJl7TmqflHtIvoY2pwuq+cpTlUvcjoAR2Uc036ct8CxSxN9W1k
E0R0TOn5/UUP33f1Xhwc8WvEqIScLZCa4VL4BtxjuP7MOGMpe6SCIhLuW8/mT0mu
xgK53gDX++1M4VfA34BPYSH7nlrA18PU9ZtvdIQzyeY8xH6E9T3cZ9UHf5vq/Q0C
Njh71YcQdSk725WL2BMrlDDmWCwMQeXwfC+GDSUc6Nb9i2uARcNjOhm/Qz4GcYDp
40KwYvbh791sCaISxomYcgkBt7Vnf0j6RTmZigzOXilR/vtCzhy5FK+J7mmw1VtF
PQSpvsLMNqZQ2qr4hwyzattgiG9Diajjcu3dpm99HXrb6MkEIBA6dIEDKhpFSkZ+
Qc7npMB9By7iS2um2x8yb+hnlZsi2LMbTtf1XOyAnx1ttKwphb0JRSZYAHIqVDCW
bwSrpwJMAjCQkl0SO9sQndcZZuSVGmDdYnyk6Hzfk/ojluYUcyzgys6LcrqvT2G4
DSyRHjy3SjAzstZg8Fl+MEWiilasJXsAv84bbUCyv43SD49oyibekA8cvTYGpzQP
oADQLk3KDyHS/ehbuKYqo4Rx6zu0kkuHaI2THZAgS88lpSmC0+Mf2vLQdtQ8rYZ2
05c78BmeDIDvRBFj+CCxcSdkBQ/oiwJzEWx3AXM7NlZvLvVoVrVaq7rARzsZVQmc
Cgmb3+Fmeiyxgez7SMXRA7FPYhahNBzQyYsl6jHB5JUSd813wLV8beXMG659aBre
3hrQz/JAefZVH0wryyoH8X0xDw/GiZg6Hx6uaY4WoM9gLxbzM4Mlwl9NtkZaPH1L
rhDBLFnau8SPLvdlTo0jb4rrO5im9Fch9CiSEQUt897woghGf7cOVOSgVjinXeg6
zysa+n0+OGVJl8SBgwyk0J23tOpPHxhwr94+TFugrQtim9zk0moqyj6bKbhfKrFw
9nWLQQvCv1hh06AAkQUQm/uAC7xpSMy5r74TT0Aqf4sOUA+bi5Z0BKdOFNOnYjCs
QG+HdfwWScWeUSPbSc/SK5xKLcJ7Lmu7o0Ioel+JJ5jKti86gKnwkCtUH+FT2TrF
KQIL3kvZk+s3MWsDGeBUHfpBV78eupOmrInThCwyiGwE23+yiI2bQGSgIroAasqm
g+x/O/mLJwG0bva5icFiya6LhavayBOV5nLyCSnvj+/hLGVx9iGSITnnKclbh2RC
A9jUYX8ZF7cxLDtG/H0iD0A5pZYwda0/aV3NFae+0PzC+VJa4Pr0JdP9P6hgkVJP
2a9r0pC2NacqJzEf5VbAks4/i2eHXphlUGVhqfo3xuef5XWwgBPFg2iNqLYVOoSH
ufhX8ZD5aevdv6j43sPe+2HGZjlxVvYCYExUXKQ+hsfse88GsS15lqPM8/7GMuv2
ADCnqHSGVfIf5fRdMpNpCdP7Wy+qu/lDcp/w7B50JL92h6x5Cgia97N1QQBvsxIp
cgddA39GzaUeQK6PFad/SY5F5E+755OpW9PkESfJl+0sqdVQn55XArsRvoXDArGo
FdSTku2fa6HHKVkcLLpaG0dEkTRGxP+k1NnQfoEC78oEpo0d2YmgKh5tL97jTVV2
LVZUTSZMSOo20mJZsqyxBDr7KuebtIUQL1Qe5yH0jH4wFzQj3dYThNCpE2Ee7zm6
285D7QOVI52suiu48GHGLVZ/QiolZOFM5zC4Ci5jkIlFfI2he5nPD2nT2lENj4Im
Ld79G4WA5fNg6sK4GKu4WFH9pzp2cKNfKjYZZXKFSAa4em1YmTQWIPpNE5zcA/aF
Q+AFlKrCH0gBtUBgkSnXXZPG4qTs+oLulJQnEOyVN6vrcrQUTmNjp7Zb2PM79lMz
ur88JwA/++nQfQyuAgsexgTtvJuhe+HdNRh66oGSYlF83JVwzcKCv6u7yBeFQA0s
B44PQwH1jL1GuR//kQHLxaq8FwUxxQdeGXeA7Wpv5ydJuf+J6K4Bla7c5zkv+7pE
JW449SDB76Ti1FJmIGy8MOXSXvyxxjJRq27TwNFzVRwynxIX7RqYguH58Z7CCDMY
hAtsyRIQvLJVYoP8PwJD+HbehQWC/jKQ+AUJrLFFmNMb0TuQ0HJWjud3hO+WbuNw
Q9ySRYcskbfbP0Y4EwTLywi3DsHNJjWRXuQ7f1FuExBqcF+bMF+xo5V6XzxUw7HT
0Bem+Uk3uYj0O/lg/oRixR86dgPTcJ7i2ZBm3a9m3pfx/TkQkgK4XxHKNKuRzJnR
8IkIOMZeDSfNDEVohsaBIyFMAelTIcfY0NeFLQYwl6nSOoasEJfjLXg5ucV3L6ns
NSnUK2XqNxLvAL8Ae6B7Rvvp3kuMc53HnvlKW630moejujn/w/lTAPlv3smWpVqM
oCRtRHi5qybfnrUU/wRT/W7VvqxVW8NR8klxMhhz+T/NoyCzdxEEwvZF/6J9ncPo
DNbuHp7sgCqej8yrtvtgnRg80X1QLJBUotcWYCKa4YNFNSh4xOQSqbg7zrPdDGYm
F1D52ZNILXsVktpM1oNFutBjx7hmOdlbZOgKvA3v9erqBoDcMVceuJXsU07y2aUj
KGB2Yc7pQxGJ33pUM6Q5d60FvlRWM6iM6UYnqgoznyQW8MBlxKnKkq6ajRaySh9k
/ZuaVyLl4hAoVNJOlbTe1SjzNey3d5VLfLeomBsZIVrfA5D0+C35gC5RpAeld3px
dqyTc02qro6KHoBzoldYgBTNoU4svxI+cbbHzxeV5TvfHfCmjGHbnmKbIDnhk0pe
gAGpYcMh4fCchM7ATgE66UvHJZMQEgniOkEuluRwxG75Wy2dNkgsmgRPL1FoWPl/
8Mi2Sxc9UN4AJD2cP6RfeWXDRnqtqOVreM9ezAEy+10zoiKRaXZfy/cnfpzqJVzm
MaT9CvcSRaBrVcqDhr2IKQBTn0mffws5dY1FS9iZOxdaUnzX6Hv/XqnugBchQx5N
0xQP5Q/j2OzurwJxdfFfOdr2CT8Y4uEOqoc9NL6JmuMEM2ZNtsY1k2NHBYkZaI3s
4/oPOTiLFtcoLNEqB0PVpJ2QnfxutMYyXadf2nNMYhcH9mCNqS1p42AkMHZxYR8c
8seh1hqml8XSV9i1TwgLyZ0sVzcY8OuP5yjt+28PP0I2uzi9DEh2bG9NhVtS5JwP
5HMCd0I8Rm/ykWOD+wN4vCVj5TJvXDVokwdgM86WDdHK55MkCgbOizjMDW9QvPvx
EFXWDTw4WYCWu8NuKgfPMNXj20VC2ytWyb3VO8pJqji9tA5q4zGQ6aD8etg1h5T0
+dCbLTqqocO7uq7ZoICw1qjDO5mtoM7NYd8YPiH07navf6OflC++In1ODQ0JRMak
Xdn4WQxgoc2vPjaLel692RFh+0aW03L0FCmkmA7xeJBpv8oQd93mrtWtiGuIubOg
Q6yoCms9TqT6scFfaA5xVdwlXhBFiwYfpHDCh9jr902tVQXrUWODXUMAtdU6fByL
QYzZAZXphXyHzvV520BH8CNYKEuolvk4HB5OSsQSEPhUdR2n0AMxB12oJmfAbcLP
RFUIp56CWm8oEPYcRgyphCUanTfCfZO8lBsxfY9xOsMLfP1SgeW+5tKsiKiVYZ2H
GgPN4+ZXetAi42rcFp6UL7FJHQSuvGXgJPdltxejSHyqd79HHAh7DDNPAmQRnCfi
LWMsSQQvjnt+9NaS9FeYZCGA0s/f+hJL5F3sgq10OYYmzH73ePGs45+jtqZZx+tu
NBx0hh8hGcNpBHXXUlQj6XNxA9BXN58kA4yz6vA3yb+6Espz8i7Jl58lUrmGD7TB
Ve8Z1jKxOB9lrQgbgBgkME0XoSMmdLzyLFKOCOVQ96axQzA2e0N2HqAsFpw+KgX+
gReq9RgG0y5S6pj5irO4CN3sCWFp885hlFKZtZU+R+2iXXSeBsaqrnI13JAWynXw
xNb/wwrspxy0mQwAK2dQDYi+gaHmL5oBIMEceLGLrXDsX89fUXdWO1sdjCE6akCy
6Rjp4C+OMCEkGDAZliOEwB0Rn8S0cXPwORXpYb1CQ6f83LKETKL4BJZ6OogV3J5D
rhQcJh46UPI1LsaJmaU1kbcmXhcfQ199qO15pq1XmNLLUulH2gLP8JGmeDS+vjDb
HinRZgRu1nuuV4UalB/+5+hMD7wdfckpHK2q4JJtUuKIJ1vNvGYmj8m5L5gNoIHG
Cyq3R0vQMfS2U8Om1wM73EXGdfaod+i36jCViOMCusWKUx40p14aPadnNUWBf+6l
FmEyVEE3wiZdsXGMOXU90qMjBKz0ynUJDS3P29RsBd3us3QjG1c1h2JvRdpARKZQ
vC6yu/mNgjKSIpckM6qFP7YmLgM9QcrJTO6RALl5+aLDEUpTb3rk/1no5G8exCjN
fMX8hz1qVXnLlACV2fryaMWh3iDXO1jciaZlzXjlFAMsKbZDn/rfkeYv+Mry7RiQ
HlFiS92lawkP16WrNrQRkg+MlXDPhGbXG0cgZ3K+muS4osdVb+0niiomS2D0CFi3
HWQEUvJcAxvtZg1rT9EtXFB/kYVHAyXQF8YGcOL2Z5RRdz48oQr8ZTxI+GQhcTA5
+DMi37Y2OUqEmevKtpcAsg7D5eosQIx2dJSlCWUvjSgSlBjoniIQ9LNyMEifVVW9
oF65nwXbUyL32bJsS2j78JAi2E3T8/1+k6EpM3yKQZ1tM99jWZ3TPbAKlYBQj3kO
WCCopdKpNDQlSB1ZF80lm+UBCEt/AjpKRcOUamSU0LJC9bTuYw80Kq1rUFP+1myG
cFE3HGcWWBHAvY9VFyZ2rOPNka8yM3k/k/154OZ6Fd0u9nE92Fr6O2aOnUbxixck
Y4/B8XNx3bV7ZhMWJWxVNTmsZT6dPzNyxe020B1NUzwEVsOJEsb2ZdZ/Cz8FCq9r
76lofCvC2aVE0yG9IjQe7MzMZ2EoqzR5zm2cd8le8y69YNmMOkwXIFszW4KkC3/v
MyVbcg72zCCt4a0rl2PjiU2C2Csdpk7Ou6cw1rmGtJLXZ0KQqffxcr0VhNjmBdv+
gPdCndwHJXPP+lqTb8QpXIqTNPC4JRKuIZVmxyyudyBdhMhsr2sdGaNcse1OUMKF
Q/vqVq7JQ3FFOgwYbGQdYGnw5q40qHEo+WcYOtSfrN0R4FqRilWNnhG4qj24m8Ok
C8A2nwreFAhA7TEpQC51HsfjTTh9UbBFU/ofL/IqCC10/MCYtzdAhbXKKu6D+oJq
/kfUr/eVVRHE/lHpfMRW8KqCyW+MT5DUJ9wTc2Cz4PhSv2FBxw/ZfSM/Q4vZY2F2
8+bTIfZo4Zc3og+tN65Qxst9++rm2h9+kTnQHeknssBoda3AZ4ZXMs8J0sxyB+74
P1IRIkeCG0LTSKK0gajpQGGWBe1eeZcggycVySjLuXVlRN5sfMRuNLcR2cWVWJ7J
WMRPyUeRUxfnLBe00/Dsk4G4uLNGeJxUq6drqpQIfBkQPod57ZE7RB3Zanvf66PJ
CPZygdmDMyb0dnd8Zc88SdQJIMW74lgs+mj+1pYQauoW179vec9TUHbg2e8XzUHe
9KmATtwQh7zeJRzBIhrTD4INkdwD4LdN08y0fm29eEYwiFObyOKl8FcjMpmFn9GY
Ryyo1Qu7+gNoqNM5mtfPgiL+OXoRmGOHnrg2ef3jnkwPIBOGq6N1jVUPdOMouJ/9
Mi17rskpLFR6CoyzB3OlcebMywnUd6UuStRufaWU9dvA8zWa/STz3Y3VIzBzv53v
Z0qvEbgLGPmBgh/iPlQYsHHpGhIFuwPS/rMZfXNrVHjPmKN0BGB1ojhlevkp5KOg
3qPlioTcstJhnFLhRexEJMWIt63VvKb3lMRPoDgjaHDJvOeqwGIWInxEbvMhqI1e
d+D8AqsjLe+KFFCOv6HIj0yavf4qT1UiXe/urjeFKSv1BbdGZv6vCku0nzgGiH27
xk6LgJQchDZCnruTcmmuTw1g3f8Bsco/yCuIYoS8YN6stfVb25hAAoB8y99X5rGM
OD5dkte5Dv1/ELdtdtCwQx2Orv6BV3GepEWHVjVOu7WSa0nVO1y1wySuGwQN8tux
mzTdNRURyWiQVGU67meBxtLV2Uj/suCSe6Y6cp/d+XLFoBZUrwVl3gEbEcQPQgrb
USqExF/rDY7wpkf8X9zsPoFOUyRvla3IzdA2R/+CQLYVc/bdWGCR9KyWmi4hwlcj
6ZbWG/Ifh1/Hkx5aOILT11MvtH3M5n6CVqhDthXMv1DshfED19D8psvi8YCe72lc
7lfO1BHcs4MKaQpjhcsMX/piGNfkVoLND5SzpdINhD9QGhpwzpcMJQXvu3jBUwee
GjSQmvSDOq3w0uW5WZ/ZQTLnK+GRPAIZKusZTsg0CVX7k86ouHSDwpGgEpaw5qWl
SZ7P0gSrZtXLplmD6xgOAi5QaY4u3/fTtzlXp4leaJYebUVDPpA5Y0Uhh5EiKwSf
BOofQYzMt5lA1cfcHWBzTrdD1UEhVFTWzkoIe154u+ehDBWlgnHml9LZG+mSUfRR
5m2nGFHCidO/sb6P3QmgnRNZvGImCNZWOLWM6qm4FZMj2RBq2yMJhoo8eUlwM7y+
mMc8h+xPm/d9wbypUZd3d2Rotona8oIPb6L7HpM3ySpEAZR4pfqF8WADUJxM7rB4
G40eeq5GcQBMypRz/Q2io5A7C1bIOxFmVLfelWqR9p20yqlaRP2LkwUTgNyVQ5tn
xUK8c2J1Ce0Y0+GzF5GMwDdva4ZWRpezkcQgFla4ey+Vk8lwLjE4vQiHhViiRGDV
jY8BU7R247RR0v2V1+YiiiLHWXmQOpfflUIiw1NGVpKgcDJ3pmlSc99/SnBm2jKj
X2pxrPCUwEZUibrxEtJ0SpuXsGm48DQxr5L3cOTaBBzq810gesYSSEmz5uX+1drX

`pragma protect end_protected
