// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
JKtLwieb269X+a7Chxq0gP7t8dA/c4Owqu4UysaaJYhuKDFvytoqiC8uvE4kEFv1
dVD+90L2IWQVdLXYaMZ5VroPbpTMN+N55hYKP4Mp3jLtorT8MDpUye+X4pUKleHC
usdIZZTRmLPKYAfW/gHiRDR3PkTfzv+qCR6KAizvyKU=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 6688 )
`pragma protect data_block
rru/m+UyvkPwG0gO2D81ihjye9RGd+OyFizREPkRRCWFDO/890GHrMmRWOk8lTco
E6y3X5LqNjyQ6c6yovlwT8CBWuOHaOlkSUOVigLxp2JINBeTggcdHtfpzQnNDJHJ
oav9Z/zxk9LtaCJQsDpWWsSrep7YULtUk+OO/XtzGmJLaeg50CL0n1ZwbYaljWgR
2OWYX85zuKmpvHSXr4YODxm1gajQSSutvC6LZWN6sWMDZxEcADvG2V2nlTA+sx3o
35cK/uxCvfvY0yAAMc4R5kDQ50DNCtRJQNOhc4zT6KX5mfObEFYqy3Dn4g4WM7EZ
Wp1BIwzSGOoYL+LBn48DSG7h2IlBw2kS2ate8v7978w8To4sxmLRSgURHC1zcbpE
3bgPwtC+FGm6vJvUgPteBbrBVsmJa5VDSq2oo+uKxvhBD2TJgFsvzAIliXsUpqKH
21mFGZDBKKPRYXOkqdHqDdAa5P8DTPgfj79mMh9f0nUQ0FY7tZhl3I4Brjh+Z7ap
ElTnFZUahPRdF2Or8vHi3A9s64JpwHuZ3xvLu0xEMjY//qrsOa7/JHUu34mnie/0
BR8q7WR8kElZFnTyRXrEzfmxDgrlDquHp3mK5GMQCXX1BZk+gakQa5uxo5UD3QJf
c4tLHcgNasAqwfi7+LDrUfXs99VykT+pKhUFEtGLfrPoQ9EA0gGfQFWwklbOJdg3
J1puUdWKWRaA+f0ad8wstXEFeCKlkiFKrmkx86C9glFxs63kAvXO6hZDydcjb3xq
BcCzoD1b8ZdgmvjIusbFGu9SImRPP4Ok6E6vmkkZVupDwAF6BFnSfwoBMf+23y2N
xeRdur+tMGRialT++BQeKHQ4uAG6cubKJiJqtKKhX1nGMJ79ertfdup+clN4W2BE
BkEri+DQG3Z9OZmaONo7puSefwajZwMa0ZF/g81YIk8ZR5LhLrZ90SylUqVIuuMp
jGc9Zhi6ICvd9ALwD5bfOEVt+dR6kenBcd/P1jK4NoWUEPDIunUwEyDCRJq56/66
hXip4F9G5vLvNYD4UNwscQxOe0rnAOOHN9nNWKW67CWZ7QX9+Ak0RPMzFOvIpvQw
Lb+jh2M05TzsFi3yepQNWCychozYdglIanR3d6eV+i3ILQIRjmzCcZFqJaa6mw34
ln6FCXCgQ0ZiKaYoWkIpYt5H4q1Ysptd0lp8clan/MwNiIDFqdWwfByGT0NVsxxm
ZnR8wsmM/RfPMCiC10DfNZT0DuHdwJIL0RBCFe2bNGs24T61ajSsXH12f7MkVWKe
iUZADajPqn/TUCuiagB43VQmEltnxmAT/vBCzdvUF23I4WlHHyES1CtO0wfpt/+d
3vGXXLQKyV4SSuYTkGFVrt+DubCbSfFqwK7wPYXWju39KY8d8zEpRlfvUIqbNLVH
1ruSaoRFwztjJfIfxryy1/RxybhO6RBmiUlAVcIVqYkgTURR7lTxEuI/NRNgBiF8
8NYHl0W8GJIuqqw96PPhwzHYzcW9+/64rJoQOxDS3Qlip1UsQ+AcTSWmK/jlOyPA
DhI37wd+Hr+oKyAWc4bwV/Qr/ZXxms5prAGN0obGTYPPUIoFk3ox/zQSgug1luwx
AQBiAaQjcSkSVXe2ySd7e6xn2JfQN/w1K3xltwcDlhuEEXcpLMbj6RcVj7m0C85O
pqWYzdqjrPjcVVlwqmwBW/rBfQNH17dMKM8blNCIeL1zntdugGToX7RvPeH+QmEN
Hfs8H5yKGeUvYQ8zsYEA23loHkgt03Ws4XzzqDsrXcfEuIbC7S78PmQby8llsmzf
3dzv5GSMTx+Sp0Cz8++HsBtg4Jw6cXbEO/7tsk+6E5CTONTDInjKGO7FCvKPw/Dr
+FqVE8xQC+QRp+v/00yebXL6CZLLNXjL33H28eeKqziEHmZ1IjjI2xE3mb7e6Ai+
+jFRZzixkyQ0fc0ixAyAVbSA7j8fRrStLDMj8qx4B0Ltd0vKNsUFTrd9sPYRp1DU
Lpocm76QboI1yF9HVJJPBi4x/Xm7EeYJmgOyp42p6CTSRqIVfDNM1ub7UsisooMZ
wdLVfSH6whYlfrBFkBhvm5/HwBVkM/8BDDAorIBwMiNy4Sc1REzN/NaljJgTADL0
8HvWmhGP3sjrGj8fpNgmxADU2Ch7XZFAlxGcSGrCeQMGAtUF0V/TWR48jjyD57EB
RoTPnPrU5fT9DiSDvJ8/vf97Wry3elm9cENa6SAnBPvNC+ki7C40YMTn0p7wrMxZ
yBb9F8C1C+u013T3l8XgzmZvwWr3XE/xccEcOUh0d8Y5c7yygAdPV86aIivHkJv6
dfvGlPvzV5Cjqye0qzNg9qQAPTayeCa5rJQ0os+rzn7KFpPVV8fnxmOhFC7M9Vuf
vX5carsEKm7e6fX7BwThJIU3eZyN8hUBCDyxXM2ZqHXbHDrRCjdMHCmItzoyrVBr
9RPVvbIqGyKa/FKWt4lMNHqO2b+oHMh5eZrbQ/7t6TEHHufRNagpbjTYANaZRPoM
49j16zqRaOLhvnFUY7fQ508L5i47KHAwiwRlEFQL5pXr5/dT7Y4rKJiHUluOsHvL
XlTb/Xoio3G45X012mBDVtoAWTAgW+5V8IG6mnxhGZECPZjTzCojz9CcwKk5qSZv
qYo/PDe7TzmUAnmi7V0ZfO0iun731n9yEHqMcblFv4kok9YlaBL4DOUVEo2Rx2/i
QVTc+Wpn6uta80GuQ4iqmLCRzqSVayblVS+gy1VtEdGO2ouctNHEyvJfyV05Ym2y
A4s9ZbGYdRbXL4es5yOZ7YkOuD1H5dwb/nHq6cIQgs2yAGkmX+SKOLHQynQZRZL4
tOUit5Xfg6tfjooCLYyFmXilxXpSJZv8aQDu8nUzU2gCLNV7sq5yNd0jZUnfRPg+
JhW/ftcaJ/jMn2VDlaI/SZLrYCLCkAdDcug9Az06vxJkXTOi1t9543oUOlgdpal6
pXg3fxhJl4t3QJZJzG++l2NgtOmofg9TNkJxiuJmm86ruSZ9vB86xH78rNFyH/OW
ruuzahVV3DxMomuO7iquijKGlUd17l8qWR2YhxCQxCjAkeiMC4WETo9NvdOGITwV
mWcC7J10o/1TS7KVDL2ItcQWHFbUeG6MHf3SVAYWvxfVnUTxHJTuZdcF0CbNpfpB
pJfUw/TAAT26XwPi1MMDeasgIgFr8F/FRLShsrFmNCiKaE/gN27pdG6DTLuaVSwh
Rfklpto/iMFfcJfQqkvuLadQiJ5KmsgveJL71zEPLxVoBKJ/GOgphivU7bc0AfS6
mFyhYepZz5hqPwWMXiay5rjAOUev1gHqPuZQ6ZfqmxJ7xlcU9/EwCpimC4x4Q5P6
+c2xCckmvw+uMJmW/GxILIdOpOcbmtEqP/RgSPJHEmVm2zmFdECwMLDjayFIvAT8
9eiDoPoSkHSVIYTxaxaWvhvE8Fpx0zoZ/RowFuvXmlwUQ//MvRB//fMYnpJQPlj6
R4CZVtaGNEd6ZhZR2ncxgHaLr5vvgDkVzAHPu4V6416WcAE36S8fLL6EJ+vcvQbv
OWRUMnomDtephNnwmlR2aZ0Ccdw1IwtxTvC3QeciEi9AabPmqXpjI8b5gIOfrHJo
xrcvD4kFj0zSxnbPA654vovxzEY7qiE9p2ort1c60JRZQEYAWsiDP3ptMKe7QBXA
SqHPtuHRbWRSgW8MVIkeXwiR9wGbEII0BQixeNeoNk9/NePF61BBwfoWDaYNFa3G
QqBn0A/0g4BTmDEo7sPhxB43txX9i0p9tH3aJv5Di1KKHDWxK5eErP8h/RXofXSZ
RqZHHIU4Lqrt2Qj2a44xHk+FXicNXQnVIlkRQExYQXQEYElAy2F3XI4ruqXwUyJO
5lpm5QsJeJ9xXxx97olatEvGy0Wibv6CD9tEPusdJUKc2uBYwadFwJ76OBZy1fpG
ULh/TPrjm79lLy89pURaZVSjTjxtHbw3/I6FmGltET9LF8WlN65eUwnqsgKHWyDd
t+cs7kIkDkNiHIGeu7iYWzT7ztXOAB+dmPEt68YjmtddQUrpVYtNS2fpmANF9IPS
kUyVnK1sntzdqVFDLaGEAOCx7PYt8T2gaoJE/KbEB8E5WyjZaTKBs1UIKYWoMMNw
DcR7ebMnwfLwcvc1ncyrEAhhlZ8ONVEx/fcxljIHVXPZzOWhQRqtYKEhtLHhboU5
AbIFqfDGLzUyGSu6RQj/aEy3dXf8Q9HTRtzkLr6Ege7NhzbZkQw5/dSq59rRzWUh
h66qCjmFXWGvZZZtsFqtn0iv+YoNYh89o7L2hEid6xlV5XTSHU4/YeB96geSGGiO
vWzMoL5A7gRBBPQqoJrCJoimqiOLoznvCYJZNmyr8TTqKWNHfUFZiFssx0OXvBK2
5ZCU7lyYfqjyHSpFBkXKhAWf0Z2bfo+KL4nfyWrPorRa0PJvDYpy5AnKoDILeq0D
PcnAtlaTvEyAa/WDREynUMRNm7KSU34mVQIwELk1rGdatmA067OV1MhUTrl9HVCC
GmrCbdC7zYk0SJhdJqnf5BGp419/9jfHHfI2cvv65BAnLUm3UfbtyOUZEzcroP1g
Kr6Aua6VcopAdtkMJmka7pcQRQhlxTZiSsYQArg4p8B9zSK8X2IpcgtKGrb6i6+I
jcC0zmzFI2yo6z7z+mhh5O/BMmYrvYkfWg9EXHc7rjGgD+GeWhAr/M7Xaa/+aVj4
/iiElZsamUedc/tMYP36lDNGYJ3nrydKQy0Cgpbvg/Q+mHOl1FFGBS7UpQH7IUDc
67bcrgKzpFVykLUHRuaC4jLPSw1UdQLWuzerLHpxOiFV3xyxwrOoHkzxPLRlP7Zi
llz5lsiaaRv1LLeTbjHgApbx5dZ7Lu4qdgG/s5P0FgWj6sa1kOa7RHl2BwHFWFYP
ljBdtqaUEFExDeAHgwr6oxKIxQ5cda4naHLm3wbM57oqNZHF7SW9ZU2oRlV2UL45
TojZahnn18NykuWndn/w7PqmTzkpK9JZOFKZEgicMD309H+qjpJ2XK2j64Gk65jk
bTC5Kmx++FiFrwzhL65PiBNYitEsJNRQ7CAYhiq7Q4va2Jr4BuK5DVqS4xNVEzTH
L2aBzySB3bmRYrUL+R50hXpYJtH1IEiOpM2393IBRj4bfFC/yr4zWH0Ed8BHx4Dg
si/M98XAsp8ApLo9RwyHC36mduzjLhrUfOfHsvnfQhr0I4OENCs7E/lDLtbNgjB7
o0s8YK9vxL7QhUYlmF7xXv75d0hACLy2AFRTDsi0Zwh9dsbcBeaHHuX2wAChZIm9
1+aphbgL7SVf/hvB7QmjrPJPfR+t711Q48hxQPLkizv6vioOuaV8J4WMOUaNcLlr
18N5SKUwP0Mq2srYMEz0Sf2PI5kG6fR2sNcis381nVAWDrush0hqlUUYFuC4BWFE
efCp+BO6m9h2VsYU4cirPClli87lAsPFp9yTbGGNQoa960pRQ++8TQhZBuHkUPza
YLOqPlR2tgO0kJZ9u2QP/Bd/SXo26BOVkvpRlQnC28IbRS368here8fxXl6ahifB
iQ6eYT9pwbyPMIhrKscYd1Ed+DOs4xcMJzLvgiZr4OxtktrkxvdukY9JNI7zHeZM
PXoyEX1MPwf1zU0HcJpMq7ojLDh0LXEJ/h5H3T5Ftr8A+lY6aiVvOfyoNJSauBtK
zCsWTBoHo7cg6bqRNYXaAT8ViUXRmIA+IjHV6+UvuKLPyH8sm4ITnqXZ/TK7X1PY
yKtqprCjkm8dabUCiFFrUJ+322RiMVIf6wSuR5WrWitAbaFOjOWcdDFVJXeItdhA
IPRC3dmSz3b9qJoryF/i5mZ3VdaF60jA3CI0R9p6WBDTcOGitYLbJWOxVKM/3yAi
0gxCaAPFnHRW5q6nXUJI9iORkus6qq8ncnFgG96U9K8c/An46raPeJV973+0VxL8
MeI8tPHmekzbFVzqk1989JxJsp0o9BXyaOxu9nT3ulfjL6Yeyi3UpBz9Yxqnor3A
bYdSwU4tlBqqUPyfjyMU0D+nrhqQCo4iAZ39ImGSI4n0+aKT9jJjb1To9fPa5B9J
XYIX+JpgE+3yyf6nC0lrgsrK6b0+A6/dXQC8DXRK7/dSwQ9wEKqOH6e6hCdWE4jh
e4cEdGuCpy8ASDkUgH64qfH1xdtMTL+vbfDlRHau2GP4+8M6uI1SDL8Afmk4PSNA
tHUnEtICe0mQS0+UyypZgvbC6/pnc1CI5miXAk4ToayUGYIAgXtbGeiFKi/uewAn
xXBJbd1vgtMPhk8SZbMHZbpFkaeE3bL+E8c+NqPOT/G28nNV+XfQw9w/fZGlCE3h
ZlyYRhc80KC2CJ5EgFQmxSs6CkCT5xJEUgGL5XFoiJNFz9RGWun0XQwpps15596k
P1lax+MIb8kba8Ba4Z3J3DTbuoPWH+Hkoa7SSZMzWhSe9Ct+/P6pnTjkpwUPl5yE
K+5h5VZrdI53wYYcjUC50BEeNPFjvH60JavTjzwWC4vBHFmeF2d11Y2CTsIBUKbx
/Mo/3A1As/PNqqy4dUIW0VlEQiY9rrBHF60IUlLDOAyt+kXQOrd/JjHtlJKKZE9e
mtGn2E3D1F7J4c+STibPse0XcmfMhXf1RAqkl0f9xE9Z9Rzl1bc0pOJ+gZqnqD4u
CRq5/sF0x2OA7lvXwtZpy35FLDugAUmf3b4O6SPLdmKMUOlYVcFI0nwzWHg+86L1
QWKxcGlLP89nstaSr6Tn0yGhY7VSISlLvC0TBRMRNZntj1GUabzzDVpFA8ClO1Lp
IhQXvKI1wILWLHRVl0Pgd2soHW56fy+3u/JX0yxlvtK77k6q1dQNnon1FUXz2vdD
Kd4F+I/LadAFMBb0kSiYcfFVOZghSSAncQOO815b1tdfUydZ7ujY1ILVutJLGvFj
wL0Q04fievM+z86MbowSYw2bjyg6s+qENLjXJqVAXwA3qtRyFPRPu8p+SXqsoSLm
QlAZOpzqXyjEAU4hbvn++skU4A3p2BPXUoWPhknVtl5q1otCZSkKDFFY9B8dTnvB
vnapKQPORZ4SZz8XVQ4hUzrhSPUVuPejvv7VJ2TqSrm8I2MvqzPj6L9ShH4eTckB
0y8IdZFOHv7EzgtIoo5PzI9reyvnPLM5jbzBBFHPiYbNWWK4tnlY5uckBFcPEyWW
V4RJgPGD4cX/RpH4sroim+SK3qGNlXuG89FA2CsR1j2FZpRGQvQlebPsOnsUi9mw
NH3nIklafT5jz3gsfohMQnO73by3YHQcgLtAkTCPWbySkZFKFyyM6MOUeTPiw1ar
5Jbi65LapFORE5BBaH7dTu5rtZSVg0ZJRQyJoKhBkmTQnLFmU94U0hUSiP9cQaTT
eQSpf79PA64yldxd6a3UAGXgBvqVJjz4iD0+ZEJJ8viw7dql9nUrMavstVCt3eho
vZ69z0dSPQ3G+/vaOReTB6F4NhJrsDz13QEHk2I8RYZc/phPV7S+/OJpg6OQuh0t
cf5BvA/Y9fmOIsGutTX4oLol9b66Nk1MZEJKpSAvC9FKerZ5XmEzVVhrPr+vylFW
jDOZPAtNCt5HuusyRQzIzhNnaH/cVOA+1nZXiz9UqL67xKkDPCxwrqpKh02FO0d9
myOvTFjyFDzZVnIlrO8RqCW55TFYlX3v/Rk6/avOwAXxtThdhtYeR7kM9rdKcOZh
RiAp5+D/PvW+BlEOaSHbHeeh7ljrC8334jVnmk0+MuDZYiZl5prWDLk0pcFeFGC7
Lf2g7/CtpDH+6hWIWdSgRptwkNHYTWPJstcOpJJYKIlKKrrxbmw1RVSu4l6GhMh/
BqAfu7Nn/f4owhEAaD4hPHgk0UxG4T4QVVTCOu2kdYAk1a9ED7pN9QUY1/r/FJ/f
uHWDGt5Ps8jJt4mFjgzczXGi7LjxIQZ62p+KOKwZTwnCc03fd9fgjRqbIk9TsqCD
HSmXitTqKvroS/OCRr/yVR3gUgAM8UMfOf8TvyXOoEEt5ojYSgNo24sP5Hqzyetk
w3gAAp8l9SdVZQ0UQQDARPH6puER4Y8BmV+MDIv+Bfx7LTeP6114z+HCWQCiTnHp
Q4xlwl/y+42jpeEKZGL2GYDi49TvdmkIq6N9Br4YIwGh+pHbYST1AN6I4t1k41km
lQyr7TlDhTejrVS8QuwcF9ripfPO4pHqsvA4n4sWC0EUWviV5q1is88Uq5a+B3TH
xsZ2UUbLRViEa1RvsDMc2M+C6BXEatt/udEj0puzNEPTwuO7RMSn7sEOCSceZyYQ
QG5fh1AO6ZC4UQweoKteQV+Q5MChbmLqFPol/Y39m8mNfLvRZWkpXrWiSex8uUHr
Aum88uJIYROv4I9MPurPKg37VgW1l+OwozkNj7VbnhJPmJirAu4j22CybUzz+ept
fhC9d4W9EsL0HwbYBodmAlKSy/Hzh6ph5kav8T4sh5C2EFG0HCWl6ySflVYoQDp+
az+3WOhJsIH/LlS8pXTjx7RknBVmjB3JIhFXHDKxzI7gJp25n9HWs6SxhU1hwQrt
VZZyrOQPylYFrWH7eipEpbtRTafBqxDILRFbDm9naaMkS0l7n1R/fLu5xadQonSI
sDvS1xgTu/DmX1N+i2K7ulRFXYFtHSlsA+8tP0f8QVhjmi4LujL3goT0wLD712Jf
bHCQ7dSaz7oxgN6scEw88ULntVwkvtc55Z0mHUffIoE1wtjbW5UDH1l56IHoPfzP
ecNjDOInfu2p1lpaU0WDhMJe8t3LBq8n/PFkkHJ6F1nqXpyQlQ0CXeVpM7WAoN5K
9e0FN2/PR9LDXHavSpe6Q+pZ7FuYBHul3vwRoaBG7uEbbAIxMGrRHqeoRATtxmIv
zR3CV+bF6g1cDZlv+4jM5lxmF0eEQspzjBzcgBpbqu/gyy+S1ZTOgISkQ2qokY+/
D011UI9MXltJBllV0Ze6g6I20MJV7FpoDqChmjiHlRfmV5UG4a6PEKN1+gqroAdB
xst0suwOAhBfT8EzgXOn5A==

`pragma protect end_protected
