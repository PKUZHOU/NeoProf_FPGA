// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
wrh97Gxl+ufBnRMrgNbzIXCp/0YaL9zyU07KnVjgzEexazdGZiuTzdP8BUPi
Om/kBeJudV45IWB2vYZITzsohcE7vwvhKDHbwpTH/uHuHRpMD33okUK6Vh8o
sKqUZbJF2y/aaQ7rSIjYzHdYKpv1hHdNbpR1xdhVuyG61cLF6nJgCOo9Lb3C
dVIbg76id8nUtrQ8dDpi5XAlUFQZ8BxSKF/0S2FZgGSbxGv/yIFcjkKhJZGA
Ov13t9X3thwcttXAAostK0/LG+YaATWvuAeJ0Eb5b8B9UsyGV23cRd1v6shn
xaoC0duBDB+oqZHPMDQG6h/Ew59aTlbhGc/JoIXohA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
qQzt6mpYyvMRa0wDfjfyd6xntnCYwcMUTJEehuABtfZ6VKIxEaStNw6dJX7X
l1wA9wEmRbmO5fjTS3JpcCYC7yn81eUxa5yn59kCvH1SAZuwxRNmykG96IjS
mAOS8/31ns0CcconSga01Qb5LREP4ZEvcdVuJKZwIpWWEzF2H/YC9awwUg1v
23XHFvGFFGgkTUCYzrVtPEunEZNEuBCEBxOsWNjV/7LBMSaw+teAZp1wEHf9
O0B2LJxFF1JDoGfY4OvASptkNbKfVQXT8yGinbiX/GMinuNdECH7G8gAzzoI
0B59VV8itZcdTulVa3pCwRquti7/5R+T2P1+7Xt1LQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
WpcF+Sauen7MATNPIWxi29qiRfEyg4RHfmqGLUOTk9/qSSw7Zr527po14ZnQ
6Ec2fM1mbwO0YwFU203dYob7CljHQUTG+WHxBeYxCJ52ZVNv15Mzy89qvy5P
zyKK/rfNNbI3jSwwn3aCHks0zOnhHpUQ5wFMIcjVStomcNzm3PqrDVSE0RTY
bLOocKQ0sBpgp+AgDTqXCwWJU1raKhi7bmSo9eJZSgxZUMneS3OCYiXyjoXk
dPC2DB+zTmEn4eFRmwGJreEfKLWSc6QKvgnLoTBc54mOxXVMwUT6IUeJa/4D
CLRgob5uitbww3RYfXI+CfSc7JWuS2fi5E6loTX60A==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
h3b4ayOA5EbKQ+933/E7XfqYDgi9YpON7fSukel+s1czuWJjP1n1OKRu0VlG
+77Vl7N/htmkw/DnZmdOyWafmoU3m5mk8CDOKYH1Pxb2DvThK367PvE7LYB9
3Sq6HwCkD3Y8sz3+OzrHwKIHvVOge9EPeFZZVrnmITCQT/Xmpew=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
gskC8qdZ6wzKA436ktAfOzSHA1ROn/KdIwE08Tvv8ab/WNOSCUTsnGsZ6SvF
2AyKMFYFqckq70ihR9t6wBhLRbKXtORBamblnlKEZgPoayGtrRng7F60iRzz
NuBGb5dgsAW2+dgU8GgObVQWP8YEEi84W13rv9UvDdns9B9/QQ21RWU8Tus9
BUYHoU5fX7tkpDU2jn0S+ZSWKpJvpT70uO4jR3DLB+A2wx/GJdKFn6x4pCpl
Y1voViWJGvd/OxVw6JMlVYQjWTkPRY4Npw9OhuMtNjsILqOaM1KPer3TLRj/
MbyQGTqrDELEQTSknY2Mxk4vHFghvIibLkvnd2IJmnfBc+qF55H7j8ZtomPO
VC1ZzkTgrsrhwvx+vIjiKy6chEVAXY6jTCqgaYApqOytR0mAtRsu8GLSHGdE
jq4OHhyNBr6p2izrkFzssoJEIjNVV03HYT9svCuAtZVhGi5+vW2UapXOKNJm
pJaN1xlbIkedQ9QTuRkqZZHJ6FYkz3Xc


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
WqDeWjcLNRZtNnYojbliJNAoEMiOTba7IhkYQ29NtIypU/ya2d3bjLDHly7+
2uOngr1hsVgcHeN1uP3MyvIJGJqKXhxD2O1Cm3tn18fdjRDDSLoaSnS+PFM6
RvKDsbQOgEFt5FQ/a+2ZBtgE/EOzuUulWZz1ItfBMxuJWRRKVWE=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Lc+Aq3m2+ehSRXysvD+WH5rHSAjNzLH2s6M1QleQ2OGxf2VY8sisHug4kyD1
7j25+xSMYV426OUE8waXcSco4xSL87mLf+uOXltIUgeBiSSCIq5GwUoj1+GX
nizKfX9eaa1kHlO31jqqzxupz4nai4uE97sVX8mHU7VGpq4r8r8=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 321680)
`pragma protect data_block
sUA3x73YkZQfTvw9mNIJjrzIRwXKWFtt+IpT7PaehrwVDJA3dUj3zphqlK8U
bGmh7zRe22wg8LtOoNxpBlufCvHsyycmCPdY7RFpnMDDgKCpeNkRxgOyq3BC
fyR0omTBDMN8d/HDZrVUp185tGgrl5nRRlZAYmFLICOGFu3ZKMQ/DZRwsPY7
vqNXwK+xBXVLki4fYk5qB6fyheD4oyjK5ZWUj33ih1yZCkdQLAsyo2mMH2+T
D2Rsh/hl6QlKEFXz5dzcNth58We0I2fXCVh+eUQE76xn/occzBEN3++CtAJr
J0366bHIzHwGX3MjHeIyklQh4IW+lztScxn7SmlsUriIpa4Mna8RBwcnY+SD
eQ1haKwlQqK26PLte4h42BbW2Fuk3jFW350/KSbr2qX/xngjZgH4xK1Yajhx
pGbH32iqK1YMBXRRrneJEVEJvXjVSi1nPl/mAHcl4ITUf63m3RjMAFbaZxYC
mAddF0Xih+xw9E8YsYP4IEIV94AYAudnF9s0GHXeH1soXLHS5t9SG+0FpsoI
vUDAqgkBZHVSb3xhyTSVfpI0wONLhBNWc9D0szx/NxW8lcoKXsqJUd6ejh5k
/QRD/Vwrhxpjun4u6PqNukpNyejKvK5ZlfsdLgBcw47liJyVy5TGbB2bdLfI
KHO/HuDkViEmmZYOHJ0KkX9ASqbjf4SlnDrJezP7InF4BtS7aGJ8hBu6k0fD
GdOnP36PISc/13Hy2beiVr/1Mcw87ItAjzOWwhZXhOb4XoeQ2FI6an7moto0
8pjbgr/EOL738PSKPrniICAV63+lOBHjDo9JxxrGFv9jQCU/2URmQRbvuJuX
SYoQhPtIOpVjnlkwkqMD65SgjwYKRxk7DGnx9ozjTHw7U/gYztW+A/BI4/hI
CxXirJNZZLopetHwI3nsM3/LzRfJqWoERmRiU0XgAj1MgYzTVyQMyCquPPxC
S1zqF0FT4Nyh8F1BtMD0NjDVfOHMGPmpk7sHz9gwdGIowaAGNnenZ0wklyON
DaHYU/I4fx7tHl4zJcDWvIuReBHrcEdX9eIRbpia9gKnxNkmsMIswStUzIrj
bhwFCz/eLdmBwdoRYN9Kud/DdP6dzyQqdNE+EsgxFgSr8t+XnGpPfNzvw+nc
acTp1pHa02HvZMCTC8a8qlpygm1Zp+SqQYi2YSdhMW6CoBalogTQLHJfMF6L
3welaDo7CmxmvNoztug+Fg0uc+3FfWVFyxr5GYWMrvt/d4MP3JswnNeSEP9E
rBLUI8N16V5oyFKg80+HvwZxPJYH8lJ+kteYstnfxa7qo0fWGCAQ99WPuqUv
OOhhHd9nCJQnuGztF/1+uYFNH2CZlOjmus6WYLEEMCm9x43nymLAmNr5qzIG
A+6Jsvh7E+KJ4a0UXz2A722sq6D5sns5GG7f5FnTUu/Vo76KeuM4Ace7VdIH
BFhIWK40CSBy0o8fPvucEVLox/B2gcnUuaQrFw3OBgVW40mLyiitZV5m6/51
RcxuMeMxBlK8R65oJ56yoZaQs0swadmM0bjC/KhSQFAbm/qaLhYwUj40XBDo
b32xv+RV2crxs1+vW1gsMvAg+uOtZ+tjepC5y7zPE+1kQS3x2D4EdUGdzS62
hWphEXInFMNOMXYnThdkTTbvjePBMNTLdATUY7qCaiHPHZBvm+zxyXuLwobX
LYDyqUW8QK6LZ4rxzqQz6bmZCnnEOAqOG+WsW6n8NB6wpeiwBW4LZRAyG0XA
DNVZtnQyCD2ogegPwh9m5Tt/aRj2geGcCGKXLE7QuA5JfYqQ33eFB5l6LFzm
aQC7mpUKexsg/sZ/W6QmPzmpHdQlnfVG1+i2pPmNvsbzI1qYOBdEVsmjDIDk
xaRkdfFcsNUcgAIhSytSG7ZaORToE7Rfg9MZt7vM4Ua/I7Re8THO/s09EQq/
dTOHLJl/C2VoKzokSE9hXSHgk1XQdSgEBlRoJRWGRL2wvUvYzGi6Hc4uXFb3
vzX9XS/aPT0UqatuOuOo7YnNOKkJzVAB0swFAxFdivi0HgxAH1LDFcU0nKc6
8kqVUHTPujWFqswzMr3nqPsv4KMHLYj9O7+yWii6ctGfU/qq3ywa11TRELmE
GGN8mIkkni7qHV2tX4O1Vpz3FccSIzszsf2nVQQEPzI6CkbXQPU/Vc6S8o9j
KcxQxrJEcwv8aJjh8TEbuPqw3NJ3gVzhaF+b7bin+xFtynbueNZOnmR/jnn7
bGrL6sL0iy6bwjnmdxH1UF6WQH3FVNGQJnNq76DsdjtuJcdF5ash/9x97CLx
agos+NbSeKtz7JE4YnStUoOrQMm+bYUADElNDXIz3gRf0qFhSaFbq5QNfA6L
ECu77WIChUZYjMw/8gzFzuntfFAYRgP9/+q3YYTc8C1dLldTwZfTkfO2LSHq
B2/x6EhsCngjKiWMKcEOcalYGhXkTawLZ391o5j03CI7q073VuKFUmTKuSEz
45Yyn6NDNE+uecQ9i8sOejIyWpOZz5MCguRbJFcDPUBmWoWea0OHxi+DOr0z
9xF8jb+irRGQjDJ/B1VVnCCD67Y4XaqEQ2atsnHB735i5+pUKESib9bOq02S
9o7kUeVAsQIu31syNFgyqRXI/6xJmGIQD1gXQsc1/2xkRozpg/a2IVjU87/z
imlam/png5WRN8sGJGamf3wB+71oOmUueRKuAgQdCoYW6cfeO+UjLPh32887
WR/2gz3QKGlsmi9xxVB6fnvQyHu43+N6CugTl0VqH4JghgJCz/xKNVoxAJR9
8JFsrcAd2nQq/NGI5Gfy1IL8R+yZEag9Uih4crhU/2lOyQNbgm/JAWvVZygV
zt6MolO1IFjYkmDAoICdKogBf7is1ok+c92QacMyUit1c9OxqaCvBzzB5mUI
DeVZqj46j6Wg4X18Rokwm/JIsCcA7dcRZRG/9EW9YOo3dEcjTRbTCovVxVUM
me+oyBReXOWcZRd+Bqt9S3IxduDgayeOeCcI8w//KaX3Rg4ljLMPXBK4jyrR
wfo4S9R1UWqXiNNU8Y397j1zXFGkD6rL9Yf2JAZmS5LKorRDOvueZlGgBBy8
yNmhROFxGNCVJjFhr44ZdR2ieG0locPo9kyo8t366GNAdxd/8cU+0sh11GKk
S9+o2MIJOdYg5v8dBtB+Rwb0w7EiOq8npqZavXoD085beMr+uEuZyFv+96/P
+NHDw48qtMTuWgAo0tRFCwOjfoAxOLNSNiiZ16xHS+jYnZjbaAFdQ+MhhcFb
zVz34jL5zTfgEnBSkpbrCMMnbTBt7Uy5VsfKDNukEGDyIfb2L3tQYbFYziIz
fzqydQxvMGoNwddTXCUJciWDp01k9d3i71DmWdNJzT4MiBaMXP2Znb2gZ037
dkF3oZsreWTxSt+plgLbwuvOsYQ1f2JaTMaok0tfzq23A7pjoS+rGhkROTdY
qIYclRF59M6jQywddY1HiVwyUDPpFMpejpS7mt18GPzCK70Df3unSb8CiMJq
dAgkCU8c+1R+LtLGveh6pbRamwAWP/gnPtERdRnUfT3fKDJhzHzKYJMonl0x
Ioa8+XL3wXaPlezLgIANSh5jMJOgytpDv1TNGe9n/Wux/XYnwwPQttN3kszH
bR0uR2Oxov9Ud3RsdvHQdW2+Qr4Ga2/v9IAXqadVchFlAcIttTCjgZ0HLaM7
lGiTv17vKQhqfoA/Xif30TwwUlhyg9QgNykQAUIZsJxPPtgXbg/RFe4W/ahd
GA0y47osmxUvcweydvLHk4CAVznt9CZhC8c/6ysbaPHhmmCy+X07IDH8akYe
Bxt1ezfFM/67e38jtj4CZcIm5vZkQFMsmL58vKN9NAmVfNQmMnnUbrCQYZpr
sdCRFjjPeqaCwCQEnQpR51P5OASCZ01slAI7QR5acHnHQgSrnaxoe1OhwF53
llLZ1QgJ2RdUjoVFULL5rM8KAXqXMXWKIZ8IkMGLLyBnIX0MJxU6m7rZDg33
jVFCb1HAq2mhCS+rgE9ITb9fjd+VFuik+Xjvj1ryR7VJFGT59qLWGAgGJglk
wab2mzW99cfwz5w+5dEcA70EWpwJDXAIoqLLad8NAwc11PSe5CNug1ubE1Sw
rnM65+e4tGrrPy7oLhJEvZoY8xsHIMRJeAu89qkyuVCrgO4gGPd1KYwF+z6i
blEIWr2GcJ8SyOMk1O2Xd6ec0sFhrfRrJtq8CZ2KUdu5Ut01SxNM4+5exH9d
l3NtqYYzHI82f67tNjvYRainr7Y4dlGgfDXal4ARPJW3tlE//gisyuc3h5rU
5qSHKu8aETaIp9gott1LyFUeYsSUXh5P1YWXgiAcOfqjUO71W2WSaYZTUyUO
V+vXSQmPJ+mS6VT+H9C8aAq0SL4eFZA1Juv6K6oFSPa0ZxXACPG0lyby3Avl
3SirixAAJ4WNz7Mm/SbWLos0SBKK35G/adsRDT7rwilj4PRvSYoscbgt37cF
wYeSnyK1SL140Izy1Dq7AA0QaIyFqE575SUmC9CzW9qcLBg0ao88BZAkJykh
+0icnoIlaYMUmYp/cMQF0HZY69NDpPu4KKoawMwfmUIueXsBjvRzSr7hPMVm
K04dvRDvWR1qTJctP5U0fCusF13n9BIYRna4z/oMSx52uIVuR3vD/kf9MucF
/iO2vZNbrvvjV/pzz58wTLtZc+wR4jQZpAk0okmVj6TxexiCoOjV/VOCsFn8
CONDujdp9E9x4Yi+RuMf2FXB6uZlk8/Ly1snnSlhjxsgjjR/Eof6/ulWbJsz
m7IfoRHG8hGSAxuX7LnukEnkSSu0FGdg+ctzBJcOzvYIvrIAxqfh1l39TnwW
ZSzg8NbMuoGtfBg942U2EfH6vzEFfgNxgAM+zgY5kbESd2X7FUFcv5n7l212
ipx2suuEU5Q6oRJYRuwyWRNSDUuqcfXwuiI4e51jKqVuRTXtjkam9CT1fKVx
dbQa//873wQI3Bhir2Gq4PiQ6i907Ma+wvHIlYghJavLOZLCr5FYIzPzvOHz
owHqVKqTcUtUYx4TXg9TTP+pqrD+QJ4l91RJt9lT0kjIqBItVEJixXIwV9aI
HmIoq3q9d28eyoWJ1l3czFvAEwX4DF8mpifBPZOgXf/58PRZmwu+lF/N8swC
8wzqEOt/lVMVscX/QNXoqrFoaBUwjoMgbXHj+zze6tfmuxrlXmkrBse5U6v4
GsLYV6sZhY4Lh1KcVKUWj0v6xig5sB0oFzQHslLtl9xNCKvGrLULmmtFBUck
osl3xcxQeIEN8DCZkTlwUiJy9AsiqxBBIPeTv7kMR/mJ3VYcw74wEk4DPI+G
i0bE9THmIR5ynd+HFvEYswyMt1KC7lkQltjiGQ4uMz060cdUQGFj1ApQFJ3G
P+Z+9LqV+IisS3dQZC1GOVNRKmbx9F1Q889I1+tqNPOnoUfA1JhzU4HiLJUD
5+9Y2ZD+ddxa07eMTpnAUD9BxCOi9k9Iuoj84hp7LzPY26CRb5eTBPPOY1gb
5fGA2GMK91BK/8/3wephcF1ShoS9otMk1G2Gix6dx0TMagnOYRyqn9hAAYVu
+ZfLSXC8D0d89J9fQv/qBQRyQlm5pDm8wbS4xI+Yf6vQF2u/ep9IVOvN+tpq
Le6O6ASUhOelbQm9yfNIsMpLp5JP4BIRJqvR2+rCUNN7yerS15YeTo8V5DXD
npfFXbwsWtmvVG7ICYJAN6OUgQ5yVaXM/8D86eXBwXTkGU31B8+eIuJKNnpT
lWyhQQiSoX39RJ9PaCDawXBQdQ+gQYJb56Wxgp7GDOeIRIH5aa3yoUoJL9AG
mUetUgI9XBL6s0afvh2FH2N8N0+QSrZeh15e8JNqI910gC+/e5+XZXgXomia
9w/HBwo5C8i3/9zx1VAdcYA3sF4k5kF1pFqwTSP1ELzNriUliwzZDT02SCJ7
IAKqo64akPiSMWz1cr45eyPgR/wK54eL1qpLoLzPbBZyIz8rsn0Ubewz4fJy
nkDeFjRBHPwyv3u2uiw/ouZh0arHFIbBpspLqf6AuWhGfvGsS9fb2/VspQGR
fCd3DR+JBNx5a4dtw8OLPq5DockjwPt/IzTmpK5akGBKOBpCGaRpnFzB5GUw
55eY/IVNy6MtAbWKCYtE+8oKxgOj96WsU4VSk8AoZSCqO676hef2BgzOSGeE
ZiGo+Cu9hbH5UO/vL/yTPFDjNFAAMjYiPrWm+pca2g9ifyzf9kSUwcCtZMXY
BkzCtRMYLvyKv+LkQQ2tXxHvXs4CbFeqcdDhqTNzfWkEGMufM8OnrKDFIVgm
z0QHjSqNxOzHQKAKZPxjhzf4BolIVnqTJyYBykGkZ+pP95lMeLpyjaeTAwen
Mg3eixu0YLI9Aez3fYms6VU90Ygz86DzhdDpU2eu6FflDkI1TsVxdPFuKKar
Lsk2ASlod/ijEbrlsNlHGcJ1RDQYo2UD5hHSgrXJexYDXYgadLzaallBzw1W
4STzL+MYJNEykgGz7qo8zL7ki7wHD/acPpTwrWHOjLwaVaJ/xtGBSr3DBJqu
xCe+J+mFXL8ePnoySDbfHwHtfS9gQoXYK0gI8uvw6hICmf/nrVFaWrroWile
jzlJIPShmMXMfc9FGw4B1dulNQFoOl/BRllGCBvcp9Tdjo/mgW9TDLmz4kTM
1b6lBan92aDPpkWY/qA+AfbdqWESqtlLwEER7CwKqztwqYhvdNnuD1rYOzMF
8+BFIxuDlduvI6LPaAMIRGjZX4bNHlhuMMvbynPDMJ6eROh7DHdw+uz6cfg7
r6koVuVSRIkffjVXLwsmSNjisWVBTSSp19Eql/sjyfdoRRCsAc9K/DNnCQSJ
t8NNwK5j5hlGAN9uERHWIiRFOUwQUUT9/24YXwPSJ5uTwDDSLbvtpxfWvdmh
oNMVOCGty6npJCLKCvcCNV3sizgbFQ4SDTclwN265vDW3pWebJLmU3EG2wCi
d8U2Jg7Diqdtt7p/LQgeNshG1OgQS5Jl3XyU6/CMNDnZxyyFD8g2/nDIPYBE
NyoYPBzi9egrbk/AaQQtoDJ62jnICkOlWfMvnhIB+IKIAynMUPrNSgfjMraJ
wdChY6sxRWfd25mA7JqJv8dGD6WkYucsMav/Pz2WHjN8rc/gU1W/JXs8UNZw
ldwI+Mb4gXbIxvDVEzyFtry1UheKOALhoGbzMOMDj/spt8EGlbiyRDJh+mrc
HDyi7xuz6vc3ZUXS+rqbnOgVPy6zusjcQOBwVAuFEaI+zd/CEqypNfxUp/4T
fH9c6h0LkGmU5OwnvYZhsVtFkpI0YzsSo4WHMrRrZg3Kpz65n+Shm5qcCHOK
qKXEPUJjT0vy6o/3adeI2Y+2g5B6edCR6x6W2HNAKjoReSYDGdTE+Qp6NlD+
dv/ttj6EaLrdPUOg5wrhlAyxIDI07cudSuj/v5nhAaL3FcQwQPX3j0K8R7fZ
8Q6kznT6HV1CwEraKfiJ96trZineeEO2NnU400JiqfIWT52TUZp5kQA9u9Hn
T4aA+PXxQMHmQQ3oZyl2Z/ocAGDAaISHc08UEa4By3NYKbt2NzaH0U2hr2fP
mxzi5iBONR6Jl92WWh70IMueJFCo21FyR6IpgoOO9JJldh/p6KKXiDKRUGFH
s2eXrzgd1TWVg5J0OZvbblp3dRXiuQYKhf2dEJwPbFa8at9e2aM9XbhBsxfP
cXqK5wCToAJgdbn+V7CssUqx9mYYYw2ZjMlz3Sb/CvdJMxfVbTKeO40F16VG
RrASagFlGhhRcLwghpSlPVvu1TIqbvRquPMNHY2jCd7R82rYOusF6AVoDMk4
E6WTJofmr6vQajo404qxOWpMUtCW/yd3q580e6mq5BfWZhVuKNpq4r4UumC4
MNjmEb5Bjd3/xq6ObrsWs+ArVVE4DQIc9BATREn8CmwppGAIMxRHpZO1R3W9
ZreMsWVxtliDSYxckDzGWPS9BRbOGhNMk6chZuz8UQE1LizZi+ZjOvKIHSxx
Wnzkd73/7fKNBLkoTBd4R1Z9/1j2UTKDo4rjN60AOjNS0dsAm1CBWY7jULDQ
U6V9fuQxB45UgrIUSpq5uNgmIqRdRMTg5I0bbwzAx7Gr0k1Cl7JbLL2fcKR4
9aMGzhSLynLPjeSWWU1gqZtq8VUebA/vn+Vvdzqi22i/69sQdv2rtlEDc0sC
WiYYGs7ONnKuEpyo/fs1mNVrseuUN2/F5pC+Gi5p8QdVeSa1Xq9H5V8Rj5bO
X147r+PSjXSbLF4DPkBh7qa5tn6X5YjE2njc5sLJzONSIBojnyHHvV63T5VG
4GtejsFeJhTyNwvMLsWBjC/Xur/8kyhOmIhj0BeAnW3pF3z3K6aqfs7h0sR4
avqbNqvXwXckAjJKWRy5nqE122ZVl5p9CohddXM5hkdvXouX1jCbDZJ2eK9m
QzuCmhOvxwmKCinNXqk2oiXt8MWGKO0ASAJE2qp8sZuq2Rx/wE68h+bN/OdR
73WpTSxjWw//UtKTqOVPbSpogMFzvO/jluR3pK5Q4Ma8RyrhKxJC/U6PvSyn
dUEmduigtfcugjPgBoagiST1Qy3nskc1ZB4z04uY8tiQjTNbN8Xw4m+f6qtf
Fmfc6WjajOtAuDo296Xzqfv/+Yk+dGoX5eXkCBA10UjXTiBbErU0uMfGCPZw
VSu4/TqZfeYPsLyF0fyHz6xHyZibgYxdERBnvYj2MmRCNbKsNthbCj9L1Y7d
++71dTjQXCSrFnXKAw7DQ69kmD/B03JlJ6ME80KyBcM08Mj0B4GUXV4fjfPh
DIkF337gWmxTKTC6zpY9RrodiMqbXVqo/iISRp/x5OYfo37sLqhH8gXSzA8y
yXCU6bIA9SnxHK8e84Uxgx5i+b1Oyf4CfLDckR6OZRpZeBLHgYwGbEiT96rh
eHgrIUqRFXyfeVAaXCeLnneGNPJERwGQTrFlx6q3vpO37OjuYbFVxT25JYqj
zzL7SvCWJQII+6vXKTOOI7juRmeEbh+RS+c5SPgfKRRWpSkS7vQP+Mh9j5j+
p39pjMKr1mAWsYQx+u/NuOCP0EPhSV2rem4Mce7SBECaxSHq3Tid1n3qHetB
bxgksMI1v0R9zkiGgveLOm1SaNDChb6XnM3Iut0bRP9wLT9xmhFUpzb5TR0r
qRc6WQEXt2mCGdEkARKcdI3OBAMD0SNZpcbg2dmZRadVW5vQQmzAEzlbg/mr
OQC2m3qyiQ5eKsU8P0gWjIkYeXjB30BCYhIzZuFj5bN2yKLwBzF6F8RKz3dH
dAEN289y1mjMNfqXnUcgrbttH/63VYUQuFtuBZAqnP5TxySiI2hbly6aVwQI
gHz5/cvCvBLrOXicz2FcrIXQ2tkew0d+GeBRpKeoTVIj8dJdXmos8OmUc9lA
bKgUSrrvx8fphPjoNX/UXVD+GRKhVdA8xOHkSDNvHyOSIV0aqn/3vgfALCif
/DKKCAzo3gVZPmLD6Row3h1Vl7lL2qBHvlWp9mUL7qKNpxgBScYA3LU3I7rh
AU7nsGimDlIVpOLWhxqYXv32/PXeQ7f7Xx4WtwnCi7rlBJefthgpTei6J/ER
UbNiwNgTXfyFR98nfzi+CGV2dplxY5hXgzACnzwP7tdlntwAfe/kMti4RzzP
jxgekpVhyagdW9jWtBew4K6Diut+fKtY0FXGhgZfCDRfMyzCQ71TFkHWdHfP
JuslTuMQCHwU9HYj4tH5HFsGhYdr5PFVjL6/ahRHlK44NN0+URXLqyjqoeK4
/YVxFEGxovRtcYE5Hu5ocYXeMvt4J3DTbmBWzldb+eFwv1M841/Ta4QiFxJb
w6rW05h/qdk0q7joFSayVJeGxv3xtlTeW7lf+ffFXIYIFgjHvIQTTp13oPKh
69XGQM/mlxmzJqZtY4/j1FtFA9UCIOfxKAcfBbsC8hkqwS1eZIKUyxJEhYtK
v1/6ta92Mya/+8zqwm9k70kMkfWa4TnBR5kZnnjrf+wp41FlqPJsU0iUiGxx
/3Tt94nFdF9KO56188Iz/hMxV0TCGMaE92nBWqMvLS8Oh2CYfeWOMeLXxsPY
8/9mbmj/QsoVLtMr8WAU7U2d+7kEnKwX5XyxSfzLcXkiVciSSiyUl1upsGIf
WNwo4F5yf+XKreRDFeyC6V6yDPCo8aDhc5fVPMz/KceIqD+KVLZYKiKRsn3y
i9QQEkW6sPNfYtJpJytS0p81jyoGa6daMvYnkn8VAwdeNZdJcPbnUwbYOGio
PG1iGCcMR6CObfQF6sgHynJMMy6vj9tdSu4LKd6yWUJp9VKH/9fgmlIaQOhY
/cl9ttgZl5dyT2SfgYylTLvCBEQQPZQtMhlLXEi87Wd7/saJSHdJEfF0Wx2k
UjBF0oTFlh4LAHQALmCVHX68to2XEHiaNw+llDR/BXiY6AltU85eJSuePMxT
A0XWG5u1stV5EwAO+AejOTwkxu0D3E/89r8z3aJAkQ3j6Rzcy++8iy9U0vgp
IAPO20IrwG/Z3gzc9F6nBZKG4u8P9rewsXXi0UKA5FUJxDBMIxs0j43rmMq9
QSXAL7QJP0hrQIcj3D5DrJqGJcdPqht4lk5uYD5MT4uTwCc3apxZZNQnHR9b
wdI4mIUMKn2WbXnr2+q0E4DQv/UmvsXyFW/U8YNaF3vJV0Y4agYRqrvYz8HI
bVWU5b6r0bwjXMUpusiBXnXqd3T2YQjHKIKdU5y2TFBDIjlDJPlW6iY+IS5W
SnUBQjXNgUbDTyC+Yry/oi7wMnXFu1jsXqnTBGOpZidrKsclrOjwJzXjKnQT
D8rYu9Wp8aKmbaE/08Qb0OEmEkM7yrK5Ui4VlaTgvL2GfUZte4YZe4+glPbU
sNMskNavYcY+XTV9aPelYWWP7rO8OAMI2Q/zz6ORipVDRNI+T67bBS5Ij+9u
9qk6mH7JGuw/8ywEbBWoW2fJrVHqiswuDvEuDEG/offQmJx+JZ7avqssg/RO
QoFiw1PFbGo9r4PwxhA0tDuPJUDmqG6D9BMjZyIn3HHRKFne/pFoGXzvbQti
8i+fzM6I4hciLu8LIKf3EGUbQ/OGOJylbzUWELYQsRPj97DSOAxhGWIQ/VyT
KnENvMeQiDkwJJkcTsiciDYyQ+A9OYXJxc7uZCkVytCCorMKJBfy76KPrvhK
AUY4vgPDMqO0i7nsf4ujPUzWW8oJK0ybcwCsCZsqMZ3B/mT7Eu+zYMBKpeWS
TBFAdqMqgqkJal4jNQxKaCT6RADC9A06p5fzM5Dv2QljhSHUwwAb0Ns8aV/o
f0jTaT9RhqZNAjghVLoKOc1s2zjyXxJFi6dv02V/YLnOA8BCR54AwGbs8i5/
5mCai3vljUBrlOd/w1MykmVcLOdiSevg8TDU6Wn1xXGjT89IoeY7boD/tGEr
YA+n+mWj7ONk0c79DC+H5VCEXc+kRXl6OltxCh/Helo3Slh60tQVXLTrNBvy
ZZsz81vY38jUlhLP9BqvvHyGJTQmeB/3rOGzSn20FUFT8Mel5Iw+8zpnrwJ7
QkeqfgJA4JA9kPtG4Foprnk4Z+ERDHLEume/eTpqJUn9JkmJr8PVUdCnCoAD
6WMwI0Ub5pktBRySiW0HnXBYNCx0SVgsMxpcsGZEOArt4D0cvJPPa8zygJAG
o3DGZdmvxb2ywvopIrGgz2ljAM31v27CYAru/w6zDVMFltn9E119DrlwNjnY
sBJXzlHJjyxmLlM2VJG9dxeRRc/SWJJsky+l1KPFRXikomnFgItnu7NPpG67
IrQ8phudvlIE6kWAXHHuBY8N2MpDDYAbg6/NspDCoUKTYBj6Y6pCBXMYESy7
Op7ao7HbotCVwgOMtvkJq0IW2jPaJ0QTPjE+E+4oRUErJ7ElfXdFsk3/XXC4
2529/8id882dB5mujEe8Fji7T26NhVB6A9Skz1E9V82E0xVx5EKLY8/yLgB1
b3StizSHMQYO9GDjPfQMwuDbp8irqV3ltLyjujgu46S2BiJalggNFmDqp5d5
FTHkjAs6x3ZD8Pw85KgnVI2XLqpm7QuECeBD44OV8tsB3wI1/yDnJfGXCfyI
QhEG8KfiqBukDCg1WnB3bDlk/PChOtxziSiWKI8bpDxmG71aNLlA6cLTIv69
DNb/Y5OvNW8VfOLJi3w3hsLNUMzNOjSNYdDnSoKi6viwjLAEBjHkRhDiz7Q3
Xtihz4MWmC+iiXbVEwDdkv7SQw0TAElWcYyEJIruMSdqf+yGn1w835xNh4g9
9Pj7yUZnyy7s5hYirMhIZ6e68/HDWzJZy+Rk/VMvemEXtrj9RJHvQsEEI7BV
uGY9/ITjf6d3n/tmWDP3u1PsOvS/CWqwTYROCk1ejXivlZsBUpoI9PvM+h5k
UtLQDQytz12F9VChd/o+KtXZWsF31eflxsT8MYViHzDC6gTKqltfi6H29Kz0
ZlIFDAX7KKjFSMa4VQuncVM6XA0g+BodMXYa+lNTiwviOGPeeLWWXi0RO7ak
MHv/ZZHsU/8r0ZNBfEfmRjHYnQmclZAqahfv/FifulL2OHnk0sCeOU7Pa5A2
XMGaKaKma42de6zFW4UrXG0ojU7YPM3WuaPrnr5W2euKG1lqoDGts0ao/tFx
VJ+Qf2SaZAzmfVtES18N8TYaMVBv5NS54uvRZFOzzqXRJ+FhDAnWJmRlzkgy
GrJKpfIM49la4KROFAnLZDKcn+WDp165SNQbZ8WgbyYJZ8fbwKRaXh2iMor4
LrC/dcMHpKq+cdA66XoZnISexCZC424WyFmQJBbAFFA6yHdztQPLYMbsl1r1
gZU4+P1lcTTmyCZkIaJjt6K8z+H8HKsiOQF9gOqe4xjudBLORRCIemBUrZwt
TKaZSERCRw5lNOzlWnpEeSkddKAMmCpUnH+02V05043AICM8VBYwtFeWkkKb
z7CC+qwoqr2+eIzj/GTZmYQqFONwneGa9Em5r7GZvCg3xQSEIjmml6JQw2gp
njYU7u0bdHlBiVWjcboz7LkKbz6kuKytdQl0wiHoAF9GXafA5GKWjtc3CD2U
v2k+Iqe8I7acB+FoIEkH4IiyAeFQsgP2ECkOdCq9Mitiy0Pc1FSMxMJbnQTG
lt59l4Wi96B5dv1W02CQTzLZeXo98ZgnGHR4ggI526QNmpkIbvj8O7lcUKCg
DVgsrtBVV0gUr7pjnkP7mNVVw6zdi/hAMK/kobitv5KRpMlBDvYYT/8YK+cF
DP0k0G7jjJw6Esp0x4IqeTwS29UYwZscNhllB3b2COS7Z7Tdzkd8DDwT810h
YlsDGOVOaHGuAh/yqqc4RfLRcC6eJOF+qiidMfRiL4DBF8bg0Fgp1BoRSDu2
U1DNcylJtXeD3rf9s30lGIiXlmD+cVzo7mVl9W3me5J6wENuDx7nMnBTCHaA
4SGzm1OX0BO0LGryzdZIbnzjEPF2ZZdAAhPm2WvWPJuNJkQ7z/cunZmippXU
CNCQKxgRDUaq+yOHsVeF2OffkCjftl8vEaTLwcA+IeP8GzZy2Wsu/ZB/6AKn
QH9yJzeQh61TkTz9iX+561K0xuUggwNPJ/oSkTvUnofR146G7eIXeGkdOZfx
ncKAqBKZkQUxCR2rYY5vuDzK/r0HrC4GADrn2X0v0Wo29I+jWrmdzReOeGPf
/sYmu33HKdjUyJFeZIR0t/tDrXjjn2Ls6PMFGXQ4SEuUKfzic7yxmWnHrvub
LtqnfBs+HTVvMGtoyYlnXYr4g6NLw5HKOIetjPfGdwci1r1ATOtvyBVq7p3c
9W118MCdQ1O0ZIdjtAOO6bRQby34Jb/oAaPvNW0TBc8YMdolsOVAGPnCIzLG
acOoPz6oBeJc4CAaifxTjnqH/r86YbKsN8b+BwCPdxO2z01vs7xL0BRPpNtK
4DkmDNJHdkgqAKrhKi3V5mRbY5sLnf/z5SujRYFbMY0q9lXEns43sEMYYc2C
buKZoqflMRX/aUKFceymCAkL0dLGZGoJ8dArc3pq4Y8JVWYkCa8f4F4e4lNW
8DliK6jmr37OGQFiqlhr3MhNzwgX/mjxc9L8GcGDBUgQ4w4QnvQbLDMsv3/x
/ZyfHEmjd+vIoh85/4mIj0F11ZSBhhDU6p4wOgN0m1v5VNX6JJ1EAy4vGWlO
JhYsEZ6epPpwe988snll+vGWycmtjC77ticzUyyi18lWd7J42abbIzRXSCFn
RN4yjtJB6LWzGSBW6XAhF3614u12YhgOFuG5xViYpfmHOqQctVajWwmd+fwD
oadXlxo5lvWDUdLpArRiz4NFnhQZK76MeM75EqEo9Qw8gtIc5UmO3A1/+o25
GUH8scwHAExJMRUg+VY0xnw/LXazr01udGA4jIkFfQnfStSNXMAZ8XpdSWxV
8ObYjiLtB/6a2BNnmKC/wXQr2lVz6P2UtNwX+lfi8ag7qWVeXh9EP/iKUL/r
FGp0SR7apuVhbVziq5r9stFwO+N4xdiuq9YhYfBFN3Y17jGKp7rj01i98ol/
Y068NgCFwxAsRcaGtOgDsJce6wD2+ngExteXmXWkWCXNNQMGw+kArUL5o2at
oUKLJqaBQc10yQessfSoStrMbOfNwlK6xZjUTBZRySfQdQhZFKuJm7cUigKo
mWodwydATDLCrSLOGVqUd5BjjK34E83imoCfDoSW0z2Nv4axeZYM7/csbs0o
OSzwUijScF1ZD0WcAYX4dFENZPZ/rz6sUtj2paFI94FzW4myRMNxJk3VniHs
1oGb4FIBFHJFqogTxruYwQ1qxNlTIORaE/8HEkN0Je4YWeqRSZOJxnv597yZ
KbBG6zYxotOsbzN2PXWuiFrUoUQz2MhZ6B7bedzQbJ+t8QVFNV2V+OHi+kFf
TJAk1fl/jeF4jo118ZMP38tWH/jWFssyJThUUePs79rU2ann6gpgKxxwxYaj
n9b3V2ksajEHthKdN2DIIz/6NBNdJLISL0QWsaYIt3qRyHBaOwAJfVpW533x
JxnY4bejxdpCGvd4MvjDkHS5Ht06EB34JaCo4VH/WlT+tNPjRTHENkRnx3dh
1UlrtT1nfzoVMk7y31OO5eARZcREq3W3x3zLDsIB7iPzl+QZajsuvC4pEP2l
ANh0Y1A9Fr7M6zMy+rfUDCMykDYP1RpTN+vhYxH2Ced8sKJ9R3wI4cDESAlN
zF3RlsrUKJq42GxEE6SomJdrR++zOs3LShNIDOUt8O7ZLUvWPnUyHaDhTiXF
nucqqZl4Kzw1ZWNE0qsE9mWb8NL5DVHZpizM9rYD1G29w/adeyMlZA45XRT8
MElno8FR51/RkS6kzwc1nQpeRcvRgJLk/dkgncCoGGwuIVChyFJNtoTK8Q0w
RO/UzS/3rJmbP+HhEYn0qcbu/ZjWOnnw2eLIAip0wOD7+Twu68ZzwcdNhScP
WjpnwMtF8GTN+Obn7HQcleH6ps642rsW20IyYNluVvm9RBWXGDvOm/Ngfnoq
3F4qtaVIub7IquWM1e2KNIT/eeZ4Z/AGHPbeurzwVp4xxo4BfIXVT5wlncAY
+M+gEnBKnnYpZJ/WjsPlL/o+wh94hiaTgAxbs67/AI1xpljRFi1lkj30lZhj
GQwFt4uJIWFl2nRGY/CMnUZJyBDzDa4P1xP/LuQ4u8ol2LF0ha275z/FI7OF
OkkmcPH2N4Dnwc5lnv4eiZ8ZJQzX3yZKK1wLXEesYO39NmkSRrvLy54mX72l
Tz5i8JZrTnMQKGq3dZiRTUtcgqStefJgtsAR1XSzioyhuZI/zzisEGQg0RUC
vkwYLTyJsmh0zYMC4ZDFBXaCenySKfYZGx4H3t393YEhXbvAVlb+Uk17Hb+S
vrjWSA0HdJYHwNicVOQM5nqD5Bjv9z0kwPRZH0601ekLsIk1qdc/lIkgTOzN
jLlxVnUPcUWYdMT4SVYtFEU3NUZ9BhZx99ML398IK/C8W+jHzMgWMZLuGyCJ
QUJwNf+4OJ7cgMTw1PvDdDz9WSW2aXhD/up55j8mHT+hHbEmHfN0gqYZcPa6
kEnSwauUqah1Od4/BF6sWCguBqGMeK6WLgNKFOYDQTjs9s0KX3McsquzRvvL
TW1iduTEXAzl3M9a79ySp4RwGXrRiALbsAKqQQCrO0zBnpMhPTMrrpPSJnR2
ZMv2G3T6TJr3B3+MDEDu2A5buz3yXUEACw0Wh1dsBr41H2ZmUUCTGIw5JbYm
mNJmiAieH5Zh2k7XSOosT92cyGqNKZX/vakO6eRoMYm8cMZlDz5qKbURIT1T
JjA64aOzecIy0ZDXlLjhdo7xA7rlE/9xDHthvapuy7TATnpiNNn7w85SAqrX
VinVuJ9lPaGTL5cpaNfa0wbPNdTlgciatBplferqyp30gUMb+l2kHkGoQVAw
pemLPlqvWXpc4+BhM/Ua5rYw926LteqAyosLxWxjTfcOkux+A86yNq7dcy1w
8FNWR6+gxljLF3iq0H81scv40gXQbFyFKpfagVMRoM+rlnZCrlMJDb0WVLRa
edk3tLg6ocVCyENaOgYD/fXtL9XgtZ/NmMo9dp3xssmBoDZZcYj1FgoX0nkL
t6AYdmlAkVIgoQj2wv2DikJaOT8845yi7wgOX9ENOSURMJckLmhOsoTNzkWd
M/mpIQUA1JxkE9tsqrB/8Nkv4Voqwovh8hpALj6GFL8DcwCG0YHzLQPvJYos
aKanXRbChoCBkMHv+ZqJj5a9aovbLolUvZ56K7pJd+WmSlifmbiL2iHtrxRH
spOgtNMZYBF/1lj+pPdyZAR2XHxtloaTFxcSjENk0HTgF+UY9GX++orZvfSR
5GRniXE9sti4hTVA2Hs4NtnX+FeHG5u28e0syOWXRxz9qGPsQJzj5JnrcTjA
gQ3hx8dsDnD0QmFYAV0nbdK88jmfyffQCXXnusNXDJ6JK64uFxaKMe/3oQLr
hg1E+3O0dG5vs6vQFhuh9h8QuKFriXZ74HnMexxoVfWea3sr7rD71EDrRNBy
/h/W5C9fICsPTXitmanvkX9JDe/E2HDuB3FJDwSmPBZTmRvqJBmGn6EjOqSC
m4LKDZONoqOUhzicDbVjiLFIAuiOfMOD6LyWT4Q3GYYRS2vwc4hFd7hoKfEe
vNLsTSKYMx9ze2gUJwWn+Yc26FvhSrHglJHxekxvHke89ninwIHmp2emSj6F
uTAn8FGkfIB/bP8NwI/5EP32ojdrHEZ80sVg7lLPyyjKjOQr0L7/kmIfz/O2
cPqdxmHwnn2P3tCAft2IX7uJ7U9qveAxnnS1j81Xdj7/Qz2KKL1GaQn8R8Kp
QrvLDPc8woPbNLM0y3qkfAkUzpMm3BIaA7liHdReL+veu194jP50SgKXGoKs
+95BEkz1IiqZlcori0eRPZ/tSXxVzkyXHKtWZpp2PdHJcO0j12AGSqnATrzW
pmyyup0Q1AyjlDLtTRJ0C1hbaJN9ATw1zk6j2fkNNWbgdW9Bm3eV7wqjRavP
bMotNHZTd/SarMRJAgYEMUCHnxcI6rIWqARQeov9Q+rx4eg9rOnQQOZpGk7o
LOgfJho2Dhir1E7ec2SO7dzPOgzMcX1aO8/8lW2JaVzeJ9V2ym2GsVO7ylHA
xYBK5u+RrS3Jvo49GulFfTpnF5EpkheGwdnjnp6msWLTrE1Z0jP13mTjY2w6
Dgba4tHbEpej6MiwgVjk52rZnFXKSd27MiZS7at+RNDOJ/dLWtTywsa+VsLp
VvvSwuPwBWzHxeajNBqE7/sGc+dGmKBE5j/r+aGhPISslkR40lPF0noSTipO
/IPHPzemaiLzji7FCyHO0AI1uZjTxofOJiWQ5Qvdfa9wR71KpI+lwHutyreF
c1U6pIqnTvmL04ugdq1BSfAs/yZ7RwpDi0v9O/yn43TrtVypXIj0WR5w1A9U
8VU/9x2JMBuff39WlZHpDBGMfw4LKQEnsQe6krobuVyWuBfJTmWZCzAq7ARv
zLeIe1oopBret8twFiTsmXJq6m0B3grOpE5bxUuJqBugUOwHLb4+sEQPxHxU
pbRLPyKLvOUq8TI/8eL7nJC9n5yObOC2FEMQpgApORqSEqkWQA0XxZ9UA91D
qV2MEnTJvsYwQiG7Hfx6R7pohMcGaIwFP3D3S4hTUWqFGTBo+Eb5mmNVORD5
RVSHIL3k/4YKgbZqD4QGx41WfEFLQCGIWc6v1tMgRg/nQObVOLJ2e83M7wkb
+czAm8xh9iD78bsxmmNzv1NAUbx5tNf9aNPN5aOlpqc8Uni415kOhuG6RSbh
ejv/iw9jnVY108X0g3P0MrkBvczUwzR2wqT7ONDsPSbklLajd0iAfaskx1T1
GkP6EYm7w87BEwutoHRusGRI5EvJEl6KBDg12JJPo06fGHlRNcnW4YgOf+v2
u8Wv7QDmu/bS86ANEjls++XNzvhIGFxCkiLomV+IzYrSKxDUJxL0L6uhbYWh
lCxw+saAdXIW3LE1BCh/wCF8Zvhf/rBIc+V9geed4RZfrocXrZVHVrLMj2pa
CZdGiNJmEMo0j0j+cy+GwR3TD5QBcpu6hK6VcE9RkG0cbwAX3K1q7cJPUW6/
jr8i2Q/rY20FjObmQVzuGR4AVarzH+wUCSR49czMQ3WROXOITdK2B37GiXuY
ds9dqlMfjhxQQNymnjevv24uXsCxGhG5vh3RIIqpWwG1zFMRgQgnNw8XBLS3
IXvOBCoFMjyH0lugQ4A00OoOGenGjp7cbTQCsjbspGMcvLfN+uX7nmXXKwek
o62+1sHp+r3ByFjCZ/nO7fwEvFhMdD5lgu75SrMX+rtOF/I6H6hTasPz2oWL
G9rIzXTriXhnL/T9Ldfkr90cHf3diZFMV0as9exl4Z5hT9NKKUZkOruKbGZN
8rCC4px2wkqYiuih4l6seqSu6GlBuVybmp07A8Qa2BCPVs5XAevqCmf5r9Pj
O2o/nOUdsUXfsRmNRDzCTemNBJHFT9TTJDkCLV3dWJjYdodJiKHcyofNggub
WLRMCA0IER/4ZODKl7loxW3JPfosQmSDxQx0hf4CPjfOSG2HTx3NlYSQeMwm
SmCgDi8vAq93eocJrpRb6Pe/PJWQVi5DzNmRcSEXxmHpIhSQ9q7jBQiKhiKj
fT1DwhXSrzLMv/8s8mf2QFAVMuFw0yWzSCbvOa7gCiRzFL0+qbVa1v6qz6vR
UWNvO8Bj2u924OjN7mCtdZqMa9DPjylZxy68dvhzcDoTaDhkmsvDOx4jFsiv
DzeFQr7WNCXZbbrWvvbcVmmIXXU0HshnA6a99E2DX3IzqcxQVL4fi21r3PmC
B2xr1rpTsSsutjukeZDBcISCNOaO8e2gxnfyx5wKm/gBy2o9mfwoACxWayrG
ecuo4HEgSK6m/ODuPyXe/RgWWpl98vP8GEeC4kjkfprEWiiR9MA7TUvjtP6K
uSrrptxFMiksQ4y107en9DYXp/eBy3KieNKL2oP14mwtclSJKu8BADNZxU9P
9libnPKW+HsuDb5nuBmfGLjA3vyKf07Ckf5KEPYesd5ie/ozdU5QRQ9K2oBI
lJS4BY3KcrMa2VTXxasRIaqKgmRxA1Rmroqp5VCANpOPjFfZN3RxOfBSTn3g
UAIMY+KxDesecxTKD8bUWmOD1fAftxVDFMRpxLpvhwEG5tPBqTMRn8dsh5Nj
ETZ5jo4kQZwPzSdzDY0+Z1Z1KidVkaT1E9eRsp02FXzxmvl8+CAAIvwuUMOG
n/7UV2EfcL/W0VzI4RRKGYgrGKUeXrVqkSsOZPMUFNrKGfspuS3zIQZ6Gdr1
+WhZGYJmeX1hSCYRBi6ZY5IsQcf2qGg93gE7jY+n3ht2QA8Fjdif4UxjIJZM
V2lYztX3ApfWDGMPVEp5lFEHaWiRFYGEbRe7aj6MyeqmmZeTJcsfD49QA4Jr
Lb1wjcVgNqZ8LWli9e0K+a/MrIFeBHkieVo2HyH4xa21d5eQdOhM3Yaen2ER
ZF+3bYOVN58moYyeXD8TOcHgBIT33cS4+juEsBqR1qaini2tF8SNpTR8S+Re
jEJfm/xJB81QLPJmbSqZoXSd7w0B/kCKeBLSvS+QAem52Te03BDCgD3nopKn
tMSKVldUH416oqZbAIqIH7RTgSTG7CVB05XSc17k2eGDH2gzmCV4VFyrGqA3
nxwEvtxjbfIBLkOOw4DLZXH8W/JNpwnp8apOnC6n5ISfEYNMJbahlHuVBF+4
2OA8q4I2Ud6o0KjBa8ETG+5eVUmZVkaH4c4PYm8kk8A9cTn/VcvEyu79Xw7S
SHWlb0Ff/Pvcqx8UPSn0XlpZq3ycxPyZYwyX0CMJ1kBa8FGQc37WAETXODMq
pMC5USmMYMlpOyQ/Z+sroNhtMpMiA/Le4VzwP9hxANfjgIycdfM89sgoTpTW
feM+GM0yyF2U6E02HEhA4JFQyytZchr/y8o5sEVD4oqvqFXBhq8NMZhSMVCO
jKQWeslromCZMLupKrbwQsbRuy72xhixNOsdM1bOd7AIvqf86ghljdS/41FW
gESV6h0GHrqX6cq3ODNEvl6zm/7WXYYN3Ap6x9avN14ssKdWXrr4jxtVuNBH
TNgYJ1xtfVVFqfvEPVkOPAC/xKDn6CbsuyRL4kQh+Qa28MFoHoWF2HmvZfu2
ODIDquNFJ80Phg051cwKSLolo0MxkQ/0HyRjf7FPuiBKATfkZcd0TSCVA/Xa
ysal79RQhQLpMBD8/L/V0g1mzrfpxbwH1BKQ7dvMDmF39MTldEJ8lwesSy8j
Av5n+zGqpVVdGm2M7uhscFY1gXXgrFKmpqMOTOD68l9qn2WZ6izniPSRVCtJ
0/DOamF49n+hQwgrpipiEAA7EEXHZ5VaLE10vapsMTmeX+3GlZyWWpSapi24
fMYdXGt2+rhG2/JqthV2rzpb3VrMuxaKeVHw8Oqfl9yU5O28w0DktMk9bP1H
ZB/w4GH7uXNyK//dtOcuPACWI3WNmxsqtOWM/843QAEXCibYeq6z68p69A1m
reeyM1yiMw2Hbjo9amfYokTsG78pTgN61B2OngwtPDA7awYAhQuwWpQ8N777
N0wxECEl0DlWJd3BosMPLhYcdfjQLOyTxR6/XGgO1pm/G1EexXsArfBbSQXV
zOz9tc9pUZNHQacN82MkPejjo0buYZr9RbuArSgjMUJlOI0c0oiAgsOEgxFg
R+H4ue8C+0yP04Kf+hE9/bc+rNKBL+UZEB74Jg1W3hg+WS0cLZwQdAJJO+Rg
RUEuEw2mAkqlf9zgUKvpejFuXW3vZX+V8kzYmd358C3z7nyoRzr6d2lGnu3I
vE0uvy41LgquX8VZo6Cbzgy0XJui18iNAPFtdWXehgT+KtJkdn6Y8UYsj054
FHLaztHHE5XBob+CYyK/jDgMGWrSqZw2PdoO9P8i3pdfoeSQvX6nb8zo1Kcg
lrEgmEEHTAltokvT/5ccu4+ZAEFygYHPRfhyMDYKAytvHegZjQOcll2Ytnkk
TrPxrRWrYJG1gyjIog7W9gZ5+PuRIoVSF66idJDTNMfOn6JuC9gGVXFOu8aW
WDOxAkD9AhtMte3fPhU7vf1PCPWxrO0runwBjbBnOzTk97+tpdLzdugcCguz
W7sVQpWJWCxPYnOOGvAgPXB5a2jMLnI/T8/XnDYvHHPoL6YG886hxPRxeTVx
20RD1eXY361uA8nx7l/necDrk2E9ZifADwEhbQrjvnKjHS26p9MVKTfTH992
W/vKgUEUyuv0CkHeyIjYKLahuHFtdw4nmXhtYDpj63zjaz9ITrhCz4tWUxoC
ijOVVTlfODeUSi2crchdgaQI0DFHgRecXXkytKS9gpYn6u7Z2svNshSHFaHT
NbFMZ4t24fbMsz4KNPrTM9hZ6Xkg3OwjDC6eRABbt9TeA7bIT58EiBsIluMx
CYK7GxA1f8FvkKWBUzSSQuL9YDXsERTLa7FGHQBDO9WuTTcNCYDPP+9GwUYW
iuWTquvTNu7D8EvxM7s+XLuATidduEdJ8ehLj+R0B/IDTzHKaXn1AcryofC5
XyLNuJgcyK8RDa3T0k6xewNJR/iYqWmouuKGAYpXXTXnXMg953CCq0bgafeo
4NT3nuCg9qTgMtxGJ1h2QTA61CmQioWYixQe/9B9dHxEjWdwd2u3UwhUTvVW
iKrCs7NeAvX+VHf+4lq+e2uZqUDNwnSeoZ77FTXcWdY7RsdwMZwl4qtdnPou
61TbBTpAY3VjV9gSLFtl9838iZSdAmCUC14CaPvJxvfMSZX5FdMDwi6lhlL7
lLt36BFx3NtYkmm1ZGSuly9D+2PSIUb125PiIpX7aW8StnXjMEazVJN3fucp
3SuwJHLzXScFdInO9j54LYTueKsf2t+YA9dSX4jz8+0KYyjfxIIbLCe4kubx
yPW+wacRGTA47V1GWtVTHiB9iHKG4lAy/WtiDjfzDZMPm/m+4byqMizl6O9u
rt2lwJgbupjfJ9x0EfYYph2oEuuT5JDV6CEzx4KxvkFWLNQEUvWWWUNOc0qb
dV0N1bWYonYfpBj8/1ojKXt7mA4LHOeyEV6e+4URiGpnQ9RxzbD13ew1x35p
LSjwGzuI9zv5wwkp0Ne+hNRA0s1bufiJwcxhuyWQ0gPRiExygLOw2T2E2/DG
d9FCZgu4zTnl9PBs+pzNv47N/iugNL7FBFaF/jHQGnuXlZcjSYU18zyxzDwL
JK/2SSin4uck5zMzgxBGamCds+emKa06hU5e/Il6qB6C+Q7JV/v9xAzJXiWE
zqjyIfX2Lop48/F32+HMgubpQjljbxB5M5J/vKRhU4Oq1FTdSriN8NRb7C/o
xpFsbM6dfSOw4mdwi3DnpcmPYHGgtH+VBTmw6XI2/5VJhD0BplTTRo5jiWsI
dripr/rIHcpbcYbZi+RYND7rq5gXbens1qWpsCsc3ImfQ4QWwinLlXJmDeLD
aC7Athu1Caw2hbaMZj+MMuEIE/LG0ElFOGtGEC6D0EUnhLs/RIlQxZIrMs03
Nt0luhScPR54w9o1iRRajqjNtPVnMirgMJv+3q/x5c+XsQWMZ3ePhbJMGhL8
x4QgZ7hD0KWOXyIZkPvPIrZ1cIEooNx/ozFqqvICu+gX9+2r0GCPJltbZHHN
Tp3rrs8cCWZUgvN+fju9MLvtTykBqCu7sHu4kO2jekljPdTBf+YK2YEZQZuS
vzV0AuincY864bVEnsZC7V3Hh1mlyBLNgsV8/mKOecJlkSKYREoJI2QnRZSa
F1baPcTbdSQkwFQuIwgHDFz0mHJRw78yzD4iPv2o14UXm1Dkq3+/fSkKx34y
j5NwTHDZi4B+AaF9UpmEiV20lRoydHyYRFK5uQ7f/ZaPYkZ9L26n9/BmmN/6
ZdcWBgvngvkKrLJVB83V2SIYZTcdsZ0LmU0QmgTanh8lBIAMVF7rzIDYuFwA
Qq15O1wivv4z4CvSnUL18g5zqo7Cq/JUil8zTYzoSWVtVKU0oPI+t8kGJ4J+
IofdJQCCug5bM1D14ItlWVmzLAzoLerjQWqqPkcfYtqGQ/fLMNXXeAqquvi3
TUoy9lryFjBJugoIZoAbVybvJQ7GaCO6+bVQd66AM/GfkAbvzW2oxkfm3Tit
FGCprK7y/G9Am2kXBBchzrFFghfbvh16cutkVugaGUrvXYkzRdu/U+u6VrY3
CXngKwhPccf6pY9acaOXyxu+yfXX5lceVVB43ZesQJ+WnRNIEtGAZVWbE9/G
FTfosEDoFHFTG9S+YjoPnGbc65Xk30FFC83itRAJcFS50dpPQLoyQQXSOLJQ
4ZPqs0pNMABiubT1/ngUo3ii3xs+Ea68tPHmlBpShh+v/aZcgt0re7cc3zo9
iOzDiSFdZ0LMxjgCoavPJfd+r0T9AcSfCaB4GSg+tKD7wK2RGYBw/xvnd55o
vngDBr93uagMm1SyDjcf+i/Z94WkwEGxOI5qfzzoF+pfpzX1qj7iEGOOmJvj
E5qxZ/2Y0xBkOyySPmRcU7QkDN+w5yePbRr3Jlo1ss5YaICXEacSF64Tniya
0gNwLI16zxH+A18/O1BkUu2GgUxMUiKrhBmoJLDIjcMa/TEdy51672V0hy7u
sIIpSWZP9js5XoIwCuhivmUKueScg2GGj8NANHeLKXrgMjVoCty9DLv96JZ8
u+GiWKFLpWEQR7G6CQzjxSjtdDxr/qP3gw/Gk0bOnJYwyX6EeZYHP+sLhUXH
ilIn7MZL8wN8+yK+mtFjRIcAPx7TZvUSHJHivQ/2N39a094+P+5lw4IAxeha
3n0KaFpT5LVdQ+XGpsYoDPYMZfLDlpSXGkfpLDC7ieSUMabUydOYmk7QX3ja
WZkHvLtWbsWLT4ZfFKd+yvH3+3LQIarXt+wvLY+14akffqeJQWGnzM51cJja
F9CdtdqZ+KxdlInsZJ3flYt3ecP8mdXwNZ7RBoTpCyJ9hxNKDzQOguEy0y6l
bamrJXgrps3uTnF8+HL0//v+p6hYR0wNi3jGqzCzMn0uhEVkXDGKXqDw5Qoz
PbdYUTkHkx/7hNiFdOQ+XAPqHjXt1YtiNhVMw41+SAxQU/IqwWbmn89GO1np
ziQuVKEJVd4xT7QWGhvNsYGX/ZCo/BmAdcthtB9KA6o9WU/BuMuiTfonnw7i
d9+SPfgcFiBrSADPpNaKqTgq1xCDdRljJr1WFxDimI/KnItRGxb/y25Iktmx
cqRiJ/Y8w1wNTs5eU/DRFcLQMZlXX+KXxkyi02JYelSjFdEf5kQfcPmUnZyc
N97F4/yvLR9OBtnnEfHSgku3r3HtXk8ed+iV2gSet25j3umRR+WF5cIrvx11
aTEz7sFzchA9lE3bd/bT5DvJshaXV3LG5FWI91UYzrcfvIiJW6qOv0k6c5ux
K9h0VHwLMh0QfvPcu+UYVuyurI2KqDnqCBTbvx3RTEmWaXkkgIGoi05say9C
LeE5//TT2JSHzKFKEmPcDmrSiPqY1ZdMaFAdYGQoYEcaXvbdZ4Q/sBm4B7YZ
gPUMpFtBwrqaosrH8MqpM6HN+301m2jRWo0kRvvLF3koTYAMXtM/d+dNYf80
gjcvxDs+wwTD140w3BcJHZwruq0cMwBIzP+/LBHrLCMALvTbRevVFeGhUO0H
vWTOs+ViaDM+P+sOztHRd9hENKe1HZlpJUVTnzD7U/TKjs+vc+LH4dlsZ7xf
PFiejR7P6GfwGBZ0o7a1TKUY0hWbHDo5TTRKETgGof0hLgNHdGP3uY8V9x7w
pECIXh7FAjZdGJIS7c7DpHTyzLdEJN4zqH9R7qxMrjPeryvpM5RFNAPdglID
FpyOy2O9xsbdy0s7yG21UUPNZMeR1Vet5zouaHFR6f+Vfbd9HABuuNjoH6uN
cHxgFlLLrlPpY5d7MZAjuL+NYkoKiBEQa+J79vNu5Q7gNwevBtkD2finRMWC
6UTzwi+Yk5Dr0BWbtjygtfU+7m2k+uZXwKZdCpdLJjpPgZkJTRX0sCPBNtyi
rV5La63ICkTmS8pyTVElvcFG4bNQnz53ZTq2Ki5nyb8ov9cuBNbW7VexcmY9
1x10EfzDT1mfUH8FzeGlFqBkSBXmIzTKsXcX5p+b7/f+A4vZNfrgSAd29KeR
wpUaG/C4vWsbhS/CYNmHZEYOd9lCwE+DOiPOd4q2OWru9MmIDdetH0pwkFVr
Y4vLC3lrqsFLvAz1lwGVecUMVDXO2S1AE+Tk4o9I14JTFjK37WADrYd+1XVc
4z9N0UPrxsPu85dGXduePEE7F45t3Yw4kfTeQoxSEtG/5k91mNDIL711uGrS
2GAYh7Q7gnVdYSsJglfSsvmaaT0jRffCLPO3A9UWM4L/2uY+Qy/LOLXfSdfU
9yC3aa2CsO9S/iC+cDe1FhayBZPrOGbeBMSF5K7rOfPyFmzZ6R6NS31+WBPn
wRk0+vSNV+fY5PXRkwAbDRUywHXibKzNXihiFP9k8yifrwnr9gT9A7Tuv4PO
K7VyktBNGOQDjvYV1lAg3W5wPOFd9LgRHByhz0SltnIq0Uho46QVolCSyXNe
hlIpQwpREbagWNGY3osKyhXQsHZ4LdBN0PLWvCfxivAdbJ2emyTiKlxPy3tW
nRnVlbHAua2XbZiqfR5MWqxFx97q4jj2lbPJ3SpjRG1n4K4+QR1oJcAuFcBm
daCzBF5ckuXLpSJzknngQlRrCI6lv8eMrdpZ+UHqVzVU21TdgLIhwyhcLE5l
XjO2ZttRYCYq29D/YW+riQ7KoIqMDkutRuZUblb98YksadzzzV47IqoVuvYh
Yb/3hJpbDKR7uyD5yIMMdOSeQpLmU6+MwbUcQ5H/CeptS3bPPXB7/8pb91rQ
Gl6RFPYPXBv8Zq2JnDorITOthEEAMYKTouGJ44xuAH/LkNBig9bEKaywfSHe
Cpm1C5DVPZ1GmPKt6Lvr0CgKGhBnv59Zh/NdUAqykT52Fzf8IWPuIrPENqgr
wiV3MFitPW4WQLsdLJQVRvlm8pVtR4hEcjkrpH2Hhv9JugUyiiID2Jkxq9ty
0jaBModYYWwKBuVvewqm3crwPrjExif1K1O1KWRmJFBYw82bFKO51mgahU+4
tR1qm4DYRN3KD1q8ShxCWWZI7ou6XmgHAh+WG4O9nfWZjJRWikVwrKZ1F025
oBYIce6q9zcMkwpIAD5D0C8MpRjxq+V81bAaDy8JKQEdP+95tjZZyKRYSHy5
BzDugWv8J8/4iTBVpnueqAGb/5cJVwRsqeXj2AHKLZonNt+r9/xezNPpoHMT
x0/W++CmoF5QMY5Y8yvB7vCknvYEwLT6hUW5UpWW2CrlQSrc0qJkdkDtrX0A
UJ6Zti7wfLxpdit4QgE6i3OT1lGLQZNSYoriIChMs7PYzia/xyDoO0/6vjO4
V3c5iCiNAEVR4JeBh2uMVV0fIPZ918oXJJttZHss79eE+RA4Rn6vMozsnyDG
ztbMvIgv0uc0CcLtkBdP81BidBSwVg8tElN4ETerJyPGymfr9KLdH3nPqg/N
7JGn+pkqZtsZjJW2Tg+xT1piQX7SMu4iPjdH7hcqggzMBHAdkbht+Vo/vBtZ
t8UAJL1QYUvxccfLN0fQVBJ2476g1BPX273pcGfJWJW7TBXcd2kFmwEWBkRE
2/2+FvzQcpl1RLvpSC2Qa5lLi/kVxnxFcNILyxp0FUPMdtaK1oEtF1PoQQJW
l13dUbTVs3QieWPw2Ke+VCm6Uyva0+wYCAdL9BHILskec1iaYADR739inOhW
0spctd2GBowPz/9Cjuc2Fi61HaLV9rHI2JUq2S8ZgKsrAsqMPfBPcnCzIr7M
NYZ40JfWXtxA3GyExLKZGT5i7noyR/fR/IRszAthOGEnadxI5LMfu/fHF7RF
9i33/mhTr2KZqJjvhu+tLVpmeOMZlxg5dFhD6KChE//BkImb7UR/krKdzV4H
VtwDuxmOKCQKmXwvO9oZ+RR0w21BcujEqiFW5Yy3ySbGLkDcna4mFwqsHDza
nk37grn4Gm9lLOd5y1WgSmEwydEcuzSfBQaB7QQY9EA6I2v+Fc7tssvZtm8I
vMyJd8SjmSmLQ8M1w8h89L+O20yirUD13aAZ4h659L0sRtPaGlVETQTlAFzn
bVEu9JKAfgMnaVT4p3ALNZ0cHMDodh7TFMLAX3yf7i+0M1usCHsTntzxSfWZ
Wa+wbRDwaHqvKDReKjta68SKu6TnumnY58/H2/N9MYxzuMZPCXyQ3IGvonQT
ng8ENjRDxiqpyNV6SWdt7wGOJSYGaUKIPEe1V1KH9dU7FfwEw5taim+93xwK
BwFsvdLLl6x0LNp8Uj96vp/WBfGPkLS8aSQnP3bJl+yNjvtz8+m3CLyHTY0j
mbgfetLu9QuiOfMrqUOZ3Axx5sseQEv+/HKuprIMVb+7mcIGB2mzKLWd2dmG
InhK08EdBm5LTtb9UAFyanOJ+pkYsry4luNZ3hbQsTG+td56UjAqJ+hRWdpd
/+spgjpdiDs1Jwr3ea7t3MRSM9tNS8uz7btqvaYT3gsYVYK3xt1AocfFdnGb
il0Gvy0TBpBtthkKr+JhOIWSepKylNQLqLOfLJ/VIGtobLZlPKXf8fFEcFRS
YgF5OMrbFy0YN9hvLVNK4xu8TmU8+nCKhNBgoezaSOT3IFDaOZQtYO+0tMNK
J19+h0NV4gOTFaNTU4z3pUhK9HtcieslLTR40XsXjssPU0vVXcIEd1HiDatR
sIBQ0nk3k14LZFSuQttWP71RrsglwKBtcXKnUdYBtjvnOK3fyOObn2gXAuRX
X6TD8Rnc04GNdoLdHiPJMy6pZBJ5msI0stnj6HbmH6lHEG6lo6j3qUQy9R6W
cpnhVhCD37wVSKCo0RdMadbDcpL7eiQBzG9npVSScmJWL8qgKFlPlb3QP4Km
58gL6qtHgNtr3/HOwZIvUwv42MRKT4Ma6ZSz4UnwzZgziZTjYuBLvRPpej7U
eetc5bYf3ncryr/4O4kDFVylUyC8LaCLxZTsN9lke4EL9SYNwj66ax2gJCkS
uAyAw4tWpSxqSib8qMkqHUrUZIJA7C7KGQxsjpaFu01bfBsWXppntX/kucaS
PD4p0o0oXIVs9DebaRRFjxtlavuHoBxArAHjGNe0DdrpZQZ87PNHZ0rkq5Gi
soX4TLG5TgdBrOj+nhaScFOHwxlDZe+jZxtiL9+c2VC0zIloZ5pOBmpPH9wF
RyFBVfGxWKD7wJfUfhcyupvtha0gRxLjGOsdiKJO9JS6127T2QI9GqMh7RQ+
kPqABV6tZHq3HHaSAXgwO/9q9MvlSSfQhpT5Q9rbh34KwYohbohVCmDbTlZq
j4GYTZdz6w2u/wOTht+iSz9noA/jJxorAXurxLnTu7jXODbMgIds5/BNAB+f
eQLEZ9QG5bTSzL54ordDfabDE+7mHgiHyNwSiDuPEU1x980DL7nzGOlfoNDg
gZnLwQDYW8ZxP6EGoX4/lL4ksMI35yR4ixTrPzTrESVtqqvmdgsXdDA6rI0B
xddWZAfTGvFwKC731iqAV/4QjYbWlYl3YvV2aJRFOiOBryNYQyvbHuf0wJVm
cW8ZwzJKVjRvLuqVMzu1crqIOa+Nq+5K9OvxbfREMhierrekgdwRz79jyoVS
rZg55fnureijzQnmZ38Re/26tj74vUgNfLpdaiq9ZaKFPYhZSN8RLBeofew/
zAgttuo4FRmUvaSiJWwg5SXz/5TS0jJyWTi4LgN8KC2p9W6ZEAypMOqyNyLq
FxCiaiq2BIZU7udLfkQQZkaRwGib8lgqRtn/SeM7Bq44R2RlGKgY81Qe+TFV
mfGm1myYv/e9wdoRI06bCBNJCPz37IKiynqP5saK7UsQh+CJMW3Nr4vdo9kS
eHXmryXOn8avRLncwFiyOvHXRy8+ePvlnZxSlRqSyqgQ8ATApe9EbwiHH+G2
vZHepKC62gL8MSgf4Tj8ay9BKrZJWfaxn1kTZOBGImLjmI086loqOHbpjjNm
5QHrHbk/QfnoxnvTU+O7Su6xF2epj4PLH3YoKiB/JuGMQ5jMpmJqr+txa3GN
E/0y1ng+yBdkdatcGEhDURnB3Ucd8/PuWudeQr1yPaPMK/fN61c5AGhclrcY
hUo3r1XKJemM8iFu7q00Rm/7Sem9/iH39JDBRnbjUJhv/jHHCuQmMeeVnysr
4XHYTv759Kx5s4ZRhk2W5n3GZRMPcy8HuyxcF6uYjYTXP2tb6ybruuy4GezD
gvIxM+mn3xPCtMl3rx5L2BfY5274pTlHoYc1+CuUug1fAO9mwlZjXEWuUzdH
bKJM9k9cGIQCBW1S6LoFTBBUZJy445YNbvAh+cjTqsdq+NVwd40ltsYFSm+0
hCVTpqGycxV8em2+vnrcji6WoZs4PlET/XCOGfZ+X0WxGXu1wBsxwINXVDfV
sLlYRiAjsF5FO3gAmiZjj90Ocjy7NL6pZLHf9WtfRIMMhMWCSwPpxGD7fToQ
7GZb364zyA7gRSgHw0XTsQAdLRAnU+Xo8+KH1F6qJb700+GJMN/sEjdfzOq0
5vmp7chRdHnAtc+rGpOGMscqsk5ndqK8Nb+2EyRKSFLX7pHXV74y0F5v0FaK
9rUdSwiTfXbTmMHH15OyqDRsx1x2/BXlDLGCP/0+Iuz/O/xIkJGZzlO8poNM
j20pqtP5SdjkBhYEGYMFg85CLypdSrxJm2vS+nyCBp6EqQbKUt5yYGIXFz4S
tUp2+74Qy+gThXX+sva6l9vE3KmkkxWJwsv04ZSi4ZnrX6GdntEJVaUS1uez
VvPA2dEPE+JDUgLP9ni7xsi9mnQmlpJkuV8Kqaakp5Xm9zQNs8M8o8pw11lX
W/7WfBesu5ph0wX8l7YzdiT1q1PNe+t1/Gbcmym3dOX6bekY451qd3tdN63H
6XrsOZmM3N7iUpB0ZhCZ9gmTl7rCdklyHZKEStKfmj1Ypjv27NxHh13hT2GH
tRk8EFp/q7PuT1CMBtbgGPFuoLmBnSF8ij/FC4DpLHNhDie+lEqiuLggVT4W
ba4eZE3tZv41/orTuMCfdPO/qaFVuTt+A0TeaGLG8+h7p+6UMbIv4qEDYh8T
K+ALqWKvMBOXtp/rZ7SytJbQcpwFLqamNd87Fcy6Q1u8TgczWz26axKDJV/P
sotNzd2L67MjSyVmDg5apfYrK+vhaRncBE7jKIm1yLRjwcS8z3tgtNQTNKn/
gav0rstksXeD0l2qEeez98sZeN2PYhxhQqI/PqCSUZf63x4MVffj0lMw+Bor
OPRfhLHWc5Sigv4ke/jrC7HfVNYJj0l9Dyt7XRJ1kG5phYEPIpzqQ5HQTIlG
n/dAWedu0asJP8U9Qlo4M+d51n3feJfwLRVLA4PpLq3jhaFQ0KQXgsRwa3C9
+t6SH173Lt31ySWibNuX1Ymiy57o6pczjLD+onjpcq+R+VPOOLPgxyn6Y74B
7G8UgDLVNP5RwrziRi+4UTNQffWav2kdM6vWH9aMl/THr3XBhyqODKHTEnM9
ktqwRSjnvZWhcOS10QHSBYD1x4ztpERrjF6WMJ08KopZ6JeLY4uIOuN9cMLv
8nHQEaW0H2zJ2sSWZeNrJ2ibuWKfHIMI+EMwZZmcLj9z5iGJde/9y4yv98GV
K3cXBvYVxJtzoSvYU3beieQDUmTB42FXitPi2Md6Mmrlm1QTOqC+lkOF1LHK
uk0vyb4tQjQdQ8t+NPvvN4IN92efA5IUyT79YqY4kKhIr46ThWNUEtT4DL5Y
K9NJejoT741F5iDavsIJHoD/EWNMHVc4+/RThSzNROJ5VUZt6XaMj5qSXm1v
C6nA1VqTotxvteEiR0Z9sfJxRStXZ7+brR9lDiZGBjp26o/lQAsBwa8MSMU4
TY1lTHXsyx5gl48WINcOqtNeMQhqZBJObQ587l5OVNxMBWjthTHXs+yhCVAe
lzs1yJdqCLxCdh+BWWnxUF7qhSF6JdfVIgFW5E4YJtG88/XB39RrzgR1yc8f
0tf3W+GnACC+pr9aaszbAI/+TVD9mpihKwK19bL1RBIws1/7XK0+tScWfSIv
GGGwV8n7CbQS1tPH+6Q4kBoqXgS0RVb4pt8y+Oni3+gvwKUOKYSgww6kdAeR
f/c+tHnJVzfbVlx1Su9aiVzutw9HMh2ri1IhC0OdWCh6glkPf3ee52eqj3HK
diraZdD9jb4nJaww1V2Mfaxmj5xvvhvfh/nC69lZLAgqyQ35iMC8XIXlQWoL
LbbY5aFODjQfuC7i3V7WRZnyuX1Z/kQ5FpFATeNALKsRhbiBiv6p8gOFXOQV
X5JDz/m9emX7fCEzXzeZ/sdW8eS4O7xMaBGTPg/FxW9nWLp1G9m0iXEZOx/I
u7LR6ahShEAdgQU063sWFfMSPsYPjhTQsiEunjepQEEW8XbLzRPawiKQKk1E
wRFuAHZbLvKp4bA05s3zmwiCtYHtpQOIeaoXz1aG2/VeRXSADAFYPLVBBHuC
5ujDvxOvFszXw4BkE+Zs0bcIojzRLJ4VFVIvlrjTkpbb7Ssg/ikPyT/lmo6T
1THx2WtzpcptjR0wJAUEn2e/cnVPUSS3eNKGa3wO0DoX3Gdp5PtgCWwwVyef
HjlHVNyKtWj0PZMUEiTgodQqSq4MSuK7YxXRTUfa8ccW+786gffkitEc43nx
YBaDF2HZ6FF9nYLb5r838HyaFdO+/rcx/KqVd1qagBhgqjQZ3Ix1TirQb3XP
7Mf9OTfqQlUCnfKbtNk4KjARrQ431ZSsUeYfbrtT/B+sS5iiMl/gzCvFmzrr
2YN5vp+0/TCpos+Qzz6xkwgGgBKipksLyqUo4MzNXR7bFSviMHZ25NTByjy8
VvlNmUOoX2Zv5zD2UOYKINICStujNErMGXx+sRkLL9km1QZPGjb62ydQ7mLk
gYjyAtmIcWd5btc5Qh4MBf9IOm4GOUh2RuKcUBC8Qa1jV014YuIMgtni/t+F
Fd5AfVVwq1YOM1iGTe+tetkrSMxfHmnmZLgKIeZWqqQoeKYMORQLjOBRLOKm
fgbQPp+fDdrValil2Zn1uRNSuIocxoFZqeKDMRKpot+6koSVT3dGXbZH4xLC
D1KPg7FSVBq5nw8NZ0Jez8G/8Gpf+e36qclPhwvdP5yfZ9JyB+MkM4qKzpg+
QrTpz5kHJxCsHSQJTZR1ytrrbH50eLazWEmWg8Rl5RM+OMN2Y0cB2PCgGHuH
JPMApcL8xWyupilLbI1VcP65JK9BQ8tBPyA9GdPOcYTX5MGPXmzH6hRfgWyX
1yloUgcLxvo/oxfjFrpIiJr7EZmxH+REnqexc5/NmzY1liJXJY+TnctEjLFS
dU+KYCnn6Cq28IQ1eOnY0pbiQpUtniaIdAHSrKePbpa36lUR9Vvmd/xL7H0i
K94gCuo+g3IgUtU1AefQqYCMiKQac1Sfxq/YONkJj/5o1n6snRcc22kquT7i
A7JlfY+uJ7Vibo5jCO+LBdOrosh7o/jBZIZ6gkKUlWiqMEwCxAetlOpYHtc4
kQ3p92VJmUC7Co92G9UIZFJ6Ab3Hg5bS02PsuL1sB5tIfSiD6WrfTUSBzq9V
TULw/dK9ln2cTC6AePV963Yuc8a9Y39gJxKRP7qxP42bBCg+8O73waErn7nT
wcABD1VZeakYz7OmomdJVD/ZFtKKreAMlde8Ndhr+szK19xd+FgXbcIxzP59
S0WzqXxvAYiwZSo5Nb2hzau4r8u8n+4b89USagE0/EiGZzxnXY6wfnBADflm
eZ+hAG/LTP4vbDa3518lWTiLxCRub7j+DfFha/celAt/0poHdYgpPxQwfqyh
OevcrCdQW/ZA6T3clMpW6GQySmynaQy0j2mRGYo0AGlD5A4ZGCAWI+qw/Vxs
VkC9ASJOnL/gaSCM7cI4XO9vgXejW7VyuvIB5v4UH1w3jEZTE7A8btjYMfh4
4ibWFvEFhJPBqnKV+sK+4vq6IDbjzd4bIWM/dhFWUOfWBPDwIZPuSoryxqhT
vkyPs6WZSWmqW0jonLd/lQwNWQqpareyv4s4sVuRIpXBWIBumtwAT+XP2w/6
1PI8DHjqhbWUqB6wMsAVIFdrZc0z8vJrbT47ou14DB+xLSW9vua+dnuBXSkW
wrcWJgDYPLjH7lIt1L0QTHVIDeLxg+pGmTMQQk9KmqTbr1vroy4Gz6te54Ai
luVOnyDvrmnE9nz+M0iA2tubW88NNFqzPVZ7itYHFPnLM2d+y65MnOTjfJcU
L1qMgV/Ny9B3iQ4Io3jZ8dYgDn0vu5XfA7gY524BG6n75jMnuY81NeXUlz7i
1K/9QCJdRtN+f37KS7bzeAyd/43N09Y+Rj+bTIzp06SGPntbxXuoRe73aq3V
L7D1FCxxFbbA57UtR9L5gAgyzXJCSyl1Hi1CLpywyJq9ZIBaBxCbFow/Udr/
Oq8BUGUxKjc924VhFeS5H5Tv3iJBMRM3R4wZB+3w4KtrS6asEwEBypTB3ayG
Brb/yrgUkAUu/SwavvrgIHG0GFjK3ULu0jcRsZiBt1k/+cmmelGuD6pM2cbu
bS+NetebwL5GSt4yLpOu9IWgbJz3yqLgMs+C+UrzX3XvhXDK5i+1SdbURlt5
vVWpQhSbvhgiAmDoGvuRVn6ngMwmt5CffVN6c5LvJ8aR/WRWuihlt9ZLCYhL
Ty65hgGumyFwfyJ/7cxGW60X1DCx7vM7KzWOhbUYra0EwO6Vl5xl2R/8a5G/
T7OA62YJY4V0DJCVyPSDpn66CL8yMxKO7TUSIxqXz5jSgwVVUox8+FBhVMLb
7ZKhZWkDEYiL2l5Ro16+yEkIEUQC2orQwk8xr+oVkVSIBcBfnSg2smPy7gNU
1UAsiEZ8VTaiq3pdAP/NIXbsqHECwzZQJq3O6jPiIPm28xlc7iaT/OhzNInh
ALmO0ogsytOQ74a6l99+Tz7eCcjYzJaPLqyJVg73njpmVwT8mheRi39RdZl5
sVTZgLBpiw8OIwUmgia3Ix4UDcyvHjdustS7RcBs+jZB5eBcj5rrFLVxdx4s
4HNYOCKdpJ9VszZQd6b0SjLcklAQbA4XuLE5bDhwHtHb5yFgotB/9NkNiKr6
lCMB/rznkSZfuDPASzceXRamz9sbeQQi9GXp81H3BnCKkNa+hmN6gOHF//zM
h3RWsTnX2KECeET/kBeKa7pgqyiG2nb878Ndznh2PPx1bOYB6/tk1ezxNcKY
6d2MHR5HXO4fkepGuAfjN3FtgWSYKFqV709WQHTvPgK7KMU/8PiuZwntVFbt
BQswNcStN34sGna60z2oXXCkooD4CnOhyUtBmNwsahhGJyrp7NQsyvFUZEeG
2buy9Me35SH6GRqeit1MPXbm5SqylIrXpmfbuRpurdjDaat1OAzyugbbBdiK
XG019Qr1kBY6zIYHBMr9k0oMblV6eyRp8hkRgHC8mxIKN4FRhYoqsaTBvA17
37OSCNOFY7Z5umPejf4Xlhx1b8NfTarQW/JiO3JH4LPsf/lX07JYWtgXp6Qo
n1SNZvFuCBAoPCHMqhLUebvVugqcnaNXA5VxU6mH7tuZAjV7KBuCmrTyZbq9
7QTXOyYDAaElJKwdNfYVOa1xsvMe0JsqpWtnbpkM5j8KOfkxE/bCBqcobjBn
FVgxsEyDUc2MqxlqOXnS9QIS2Q0JdTlTeThjZoy3rTgsaVTPfByWUxaSzPqx
eg/6dyMp/0iv5d+i0jPcasuHp+t5SfsTWpUVTH6LYE+T0dLH0XJWxosf9i/M
SFsl3k6Db9CVuEWvhbwROpWJCpmnAKtDsvDoCChy9QmDoPrJ8sj2XfdHLXUp
BhXyV3zkT9cqhu0ATRy4qOCVSs5vi8k4HzxLciA2ArL1Us5jewC+AsirtAsC
tbZFwR545eJhSXkqi114dLc30lkpf+sObvqoNoelroSlT0Dgt7tZTNKSWotE
yHFh+6yXbBEawqtPHJj2YL9JNnf5GRkYuAjyKuq6yiZD10tHd+3+MEIMtDXe
XhXlG4wQvNgGZTKTSHNrpMQnIjASqgUds7aH/qKORztH0x8pJ8F5AObnMHrK
zHDdocXAuWfgh+tRFwhk5WqtCBRVliWDn4JpqwXnG7rLkRtUbf0C8AqhB/Ms
LpYaqqufgXBNLNDijf/WwQdoSAmBHu20hBTu5NfkUtJlpCprtK+tp6Isr40O
7dB/wmERQzwWWYL3PNFHgjmlJuqGA4s3jFwAB57N+yfY71ZU3c/joyXgRSYa
m3Y4HJNblXLgSv/im9eiIe6XXsy/w+J25Ns1Yd8OM3Zz56BacEbOInRd+dro
Suj5zgdbbu6QLxYbxKas9JCISQOPAc7pO55MyCIalIXHZw2c60OD9fPsA4pC
/SWR6O0L8FtQ6YdEm1FXRe2YV5d/AkjvnkyRkXwPG5xa+vemVjpPx/V1i3JC
6Q4654mHfeinxCNZedeUqLmdztsFCYyxt7Pn4JhjdEZPYGAJhBhDmKg87l/N
zpo3qw6/W5ctxu4aoGg8wN0D9op3X8PxU5VMObGQ7lxx25J5syR8ni07/mp0
nuzKbw0aGeBZgFhrWABqcRTncfYmK0jp9Mqt4ouujWAZLJfbivFiR+lvHRdY
Ts+CNZMf2gHhmmM8pa26gFKCD7hiLQZONh3xEJj3XtB0R4DQCK4UmZjwluy8
2SDrfjbidK5m6YMvgS18TZ+Z+/vhUKB5dE8/V5BJ1CGRX3770s9vMa1DnnQc
WxqSwaY9mfnGRHihWdd0g1quWcZvgc8q7ObKDdbhOXoRNFIEXB41dJdiDnCo
+mzpNntgTMAT1ofa4ztYvB7UAMQ/uhNzM+8p2qB2FGDFoJE7vOCGq6C1d904
5BQKYPJXfRzAddwTGRLjfkZ2owQt1q3+EyDBv4oUpJyAQSM5LjLV464RBMLe
CnyvlcczXOtJTmrAVZrfpXMZgVp/xW26wrbpehby2wKrvKuitljwCxp7IeYZ
YeepnpWt+7RcEhJKy/bdxVkOQxPlHvwXvvZHKOtg+xrG3SzvrnzlE237QhTu
PMJKJdaij+7TcLMi4DrqZE7w3JTEtcjsqtmJBzkl2zqCCNJogxDTicoOq/tT
TIHXWECgt7aew40pXAVSp+mgxyqM3HDs5CI4S8WkA+//YWrMXvzELPziK8cO
QsFTJZT26dJ2uSVbCBFrJSKSSkSrQFBG+h0slTN/mdSRTsmFzoyp3WiOg2dD
NpP4kbDvVWwRHRy3QuNvvwr0YWaNcjXdwcRBl9zabT679Tf9liJkBbp9wpkE
1PccXKdTSVO+xtYw7fh679LBJUe5mUR/AXXbrCF0lnx6GhaK40oaTOkq7+PJ
XS6OK8sHSMiqbqmKfg1UaCaemw4idqJwZRkEyPi/5glxcn0fahDlXSCv0wU4
RrhMGrovesKY9c+TxT8M5O6tMtT6cVY0jCciEqxi+VEDIF4sfD0AsE/5Qrlf
FvL/F6PzMai8ct2h3eD+astrUmMjywv+79byE2mz0IMZS7JmVjr/Y27/6YJW
P1NkpX/G2aWNHxz+V9jU68w0iGODrkjkhwVt2+iKfb4UCWsNxXKwbWHsNJm/
iiRy4Cpdg28jJvHh04JcTAVBb13rGPXRbjjRPrk3DridZ63PLwWRb39r52wY
EI4jKFB8o8Ap2r8ShmmySxqNyJoTOUxYHTPGBdn5rLrNHv1MLddTigGNVCuE
lT1GFy8/58HaUMsGk0vdLQjnVu1yqxyfRGvqqm4jdLq+RGJ3lfvNvQLXv5Vf
uu+Gz1uzvVVaHvxsoNtSFy/1ClMec8H8xcODjO0uACaha9FNdWoedXoAdAjx
A5ILqz51v0Rldx8hIq+ZShmig3LTvFSl3RisMrtGRt86oLu9HUam6YfaC1D4
7D2E69S0OlzjatztPzcY5R7A6OPYmxP6ULDy+kC7sDEF8X97eXPfPPVvv4vY
PJApOytoomOHbF5eCW+tVAWkGW+NuR9n4CIFXE1Pqe9PkDdyu4xYSk/z17+w
EtsfZaw6S/R0ZN+4t41k6W+lXV/Tu1thM6fL0JEIUUm2enWn4lq3UEJukvGB
auLhogOZjONGUsHWthBwEziNmdUFT8bQNEPs1VlmETtCljG++skoouRhX+b4
n9eFAUUeGtYoWN0I+134zyA7W4lsc9lGjYLSL/58BgDpjpvzMuSiY84w3HAV
fSnTE3TRizJ9dNl082+JjS6Z4Bf98c/jIk36aCW1e/nI1aRPuRm/QGZ5qrLn
0cFB8Nr+4o+wIBuBTQSaX54doeDaF/IkXWUqXfGI0dXExtaCO6Wl58qov+c8
tiHOx9cRzjNkIhtnqYRNGB2/G6+VhjI15zmIDnaz7eKHUKCmUiJ5f+lpsnw6
9g4ryy3kcvfwtmH5pHUrsfvI7LW+ZpFatyc4GdjDC0Uv3mUEJ3tWtFdKbO/y
nHDKj5819Y/faTkEAROLZhHBhFeT8WgbENB0RylJD05xzTi8/rvH5I5Elz3I
9+Q/yGdwF9eCEvlmAciWrxL4d6KAZffbFCAgsiEo7pwCjJLzxbEqhoidhnnm
kgrWaW97NDzmzkZ49IOGqVPyGLcHdhqATcGDut/dCSjRgpc+D1wIjqXtaZRZ
yP4ZAmjJCjMIOPx8XQSfxKJ0zHL2JYxWw9bhxIwXCXdJOrEkSSG8ApQ6YOPn
niwUrLdbzKILO+P3/NINxW1uGapY8nTjpUQ0tAy+8oxnWIEug8ujg9EJoeNL
B5BvOQIDaW7Yy9zcKbqiaaXxwFgZkMhvA6YbusRfEwyViI3nzQjUc4wGPFbR
U+YOhpLoo6FJ5FDiFME0mjkRPKwDzhh3ogfOuXQoNHu04UYhGu+Kjnv0mOYG
dxJxIJQ+fYLbQfHE4TTiwyMGdBAcZpsPGVp5WH6UdaBjzIOno3nhvcknsm7S
vGIdVahRsseJzq1XIFmcN3WerhL7uGKcPBrGT3be/kLYxEpn6amkRNEnb3Xs
88E/6R6N1kMB0a/Cr6zreRhyLl5hshrRUI94IECPmwMcD2dJrHTPVW3AkQyC
YaPm1BEiyejbjSuLjxjHQPa60QL0+j0tgc2BQx8T55wyDowuzI6dXJWtk0wq
N+ZUfytMUQkRsSceXyOKj0lUo2Cfw/rkcunh2ABDfyAk7F+sHmMJeIB9n2Fc
5h4fzFYP9ohg3y38w3uF6br0AtiZqS2HYl9R5e4zYP2sIJ/ts4ICQjqo6H3L
NNBa/OOhze/LYUz2HeEp8MMq8uQy5j+Vtj3LrHzjyz1CpFHFRkwfcdfxQWWF
H5ixP+uoTmIA2CZ2NUQg/aDaWMQpGDcjEHfyWJoUZIrHHO1YZW/INTVQ/8KM
oYqT0sCxapChjxFMsXGPnqvR8ETv5Yg6vjXX6SAdpPBDexJktQJ2+1B82OvS
fBywoYGtc6IZRLUGn2Eje7r33Y69Zwi6W24NWwa+PtzJl554zQT47gWGRn8h
peHhTM2+BCkVw6nznaTtneuHKLobXP71SZzrtX416Iu5b/nt3xYw6Ws9sy4o
X7+g2Uea3pcqw8uBIORlgcenFIxwdCDyeq3f0TPkYTuFD9tTlAlWs3A8fWzs
yi0XMQdUZq6b66jOTygy65AnYbFNXVhqx8asFrubtfdKcWoP57zlfxC+4VuO
w1W8LzXIXUX0DvRTfhvzuYHrYmrNI6KRTT6rm/BuD2eLDfJqKPrsnbmTSxme
KvIu4ahpQW42/AEMe5TECeMFKIVfZIttlOHzk7YDeORl3M0/W1OFZa4Yl4J9
gzfpshKH75IpHoKc6x7XqW18te8Tl5VriYjOdCH6Jb8xcZl8utmNeUyLZM9/
ymztjnC1y/7WpSYJuSOgYCe7rebSRbRLQGJrusz8sc532jpRaKCAr7KV7mvS
uXTbyRHVa7SlUHJlyeDJtMJZBMzx/5JYhs0nAgIsV+bpySCbOk91Kd4QmwZj
/1Z0tKBUWIC8nt5DiJTzvl2whbkO20gxWaOCT/W+s/gYV9VhHIIsR0uOGLqK
dYcAFIYzFfDI1vXiuWhuO67/zkdyN5A6FOJtXRZSBXemeJOTkEOlCbkADShv
IS1UQ1nixW1nOqEu369l59C1GKBtjpUThZychbGxMIMy1mbnhk+ozjkQnXnl
PLOtZLO0EBjjGwk0hjMcwVVp6ALOZLDX/66IFFh198++jV8vS3/DZM4IDoxc
xbz+/Po5jbTnTkn7OVL3NCv3YGCJ8We6sDNGeJwQ9ATS4s8ihTopBXDAGtfr
+VekViz5y3h9had2zJh1z3Fzz3xPaUI5K8FkUKcYcHslJw7HPUr2zy+dL23g
UgCmAaQkXkebFVVrNcgRId5COHEyYZo3uP752KAIz8PC0KxGeoKLuTjvDLt6
k9Sf6p+wz8NQCCSw660QrxilbMHWkhZfExBa+u/rNldPkkQLuLUWfm+OxNwF
IM3BHz00PD3PTVcfJMyjLcKRTZWDKtYn6BnM12UF3OGXx2z1lonhEZA2n5cT
YQQUt/OFFCiU5TouZmb4cWBbCMf05qs/gt1A6pOqnIeP/yzbJNTtF4eqfP+r
gIIlJDfW7a8hqJbCfAampX+EV+4TgScwFfDafrtyeZsTlWg4/+utgxkRQhQN
hBKLnsg4LNMjnU5EDV2GTFLQE1m/fnHpJEZ151cEcETCzPDsCj3RUU8MPt7a
dwfRsXOZI99VbUnD8afy52/DhYnRheJyig0p8CH3Pm4Qrjq6ck9FvDy3ZAzo
lOUF0yuZWJw0HIlANoRsPTaAamcxMkIiURXfKJVf/ojyXtfdip2W3aPK6eCF
8KiuehdaVn3b/gwNTmSQZKrk/efBMpyg3ZDkQKfaZJDOsimYJXX77Sf8HIXx
kUTSeIYmsHBphqDSusXvPg1oMKbp2pktfdw+zZ/KtQ4ofkkep2hIhvuFVD2p
REIk1eOFTYN+EQ2mxPqBtsFOdWywFgm+JRSdV0hIE1ofzRV8qm7Y5K8+2xLK
Zrf8Mu2OcF7EBCBOH4C9gRXybkk0HtgWW2KNOxEBHBXOsIR6cgPppMwIzb8n
LAtuZpsQf3IaK2Zpi0caUibxYx+BAKsJfOakn2iJ4Jhgj0VIMPOgfpFHCUHG
loVJS9xZloMs+H9KawU9KQe9lqD+6RoXgMMIJc8H7z0ALd68dU2ywMxg6YD8
y0WP7YDn1lB9PJrlfkBO2CjWivWfh9w0zvTuBsiVWDJTClpiXpmV/O4xS5sS
hX/riaPfIqWa3jdKzHsHYQMKkLG2Ee/+LMNDRHKQ4iAv2DOASc8052bAZjjm
I5WLoAaZ8NJUmhzVUZUhL0RNFbpMCvHqfXPuQzCt+s75TnjrQrObtGmnb/a6
mNJMVDgbXjHx7Z7V5ujS3IgjTCEdwyx0N0POLn7jOrRPnEfDwtDQ0fgdBQNx
HKEhIfMXUgE6bt/ex7Dd8W9ZZcLb+VuDJ63qfglVdujH57zkrBWCWdUhsCeJ
KhBA28lslPnBpY/7B4FiKtyyX2M7IuJ0Fs8uJ8zPKoxW5sByTfBq2cSht7Lp
LUx4MkPuDuoX8/kD7gXhpE6NpxNdOkYyWvzR37yKeSFVpoB0ABJnveoBAu0R
6PpEvnfuaIWpwE7kbssKaq9Agq0Kea87iTZXZgJMd8KK2pjuQ9cnynenzjmM
ahXO2SMAhvlMpgwMzMr72ixv0r5BuaEJv3LKEW1ZNCZNh6eqs7NV4AQLpZnf
sQzu8742nRWkhugLSJDEdovX07mcaPgzu6NJt0tvJRXOrP2tvmUGvMENNdzF
tvioZnHWCU+ygBunu89WvLBfcSMDcpO2b65FxagCKoBuno9nwao5jaz+Htfx
mfIB2E0DJ1xxx4D1EDVlG8QG2R6YMMmeuGnzQGlaArNK/tM/xgfuNTdME9jQ
lDk1Oxyuz/AbhPgHUfZnvvvvnEM1Vh4u1Eh8q4wODWp0TW2p6KLpoCuJZbDn
WVlL2zLJeL4mcBbPcy+1gtkaW0bZf4El4PhhmGxTASqk7COFrBGF1AKHoywK
+Xjc1utyL4FBDXV1myXprZtmdsUx+LNowJaedAmOpWeVOK7limJ/NfKb6v83
tGNiLuhUtlN/kJotb+JdO3Bk78+Pi6oPaXKKd3tzHlNh2KNQTTMSdyhkUsXZ
Hmmcner+wQDL2Za6fFu3wTA6j8kZQt5wMm0cduWQShNXA2SreDqf0WwzdCUe
sLwT+TAlHyo4DJ5Q64OrLUpdTnCSj/yzBpsJSDS7pn9hRFwzSNJSExcn79iM
LxHi+eGfwj90vzhrydKPDiLmK+VwwNXW5ptNVqEPp0Kw9CJ7Vay0ln033y1I
gRJdYJrX7xAfqS5ZsYn9RkHK5DupTOgvsNoJnETMamuitaaYFhMBwxFD5xCV
xE/rTw2gAPXV3NSLOx25ZxBvwGSMKUE3mI4BovY0Bs7PFPRAguJQtgXNv3We
L0+YlBobZMCzXtfdZn3y7bemi7xNkZhh0JQZyK95lbUOAq3AcEs/6wyzStkc
UseMcRG0F9V5qpV3d7RezT3Btm9ys2e4Riyei9KDYvnh2NybbCY5US1F5jV+
LNMW8wWOMjIkN6zjJVG7UxUzu0QARGqwRfSSiu0oY1auqeqJXPUozFRCJmjR
qpf9ZbcHhYhQMv9PDiUapI0azsAr0zVfnEaUU4M1Oeh54MpThQefhsC+FH9m
YYm+6gL51bfu4X85BRtHXQ+sCWpMsdZraW5VGgvNsAtwvQcXIDEHnY7l8ren
4+xr0HnbYw5YfyFMid9Bsopx4HKG8ty7VxuQnZUxK386DWzdC5qZxGADVRha
WdP5fz9GsBwCbW8yISDQx7hjfmu3aVunFsp7hfZmnGE4NbT5yet/MZDTAOWP
du02wUN+56by5DuvOl94/YmM0lZDdhrV5npHpcCUCFHE7dzbTz4PtN/Iisw0
3K8XTwJs/BwUgQhbVsfBgtk96dhBxl72TSjZ4qjejXsQ9qdSq5wwz8lg2MRH
HZZPR0bFGVezTqWR6T7MeQYpxEavTPTA38ToPs/mpCGYxfosYbPEO3HOhK4N
Cl2W43jjQnm+MMHcn2q/uERXZoBlLEwP/hLUTMqnHlDq80OijCLZnd3aE2+v
iQZZW96jjJ8ecZPvmPL2F5wjA7wFenNblUCGHLCg8AU3sdHlQlHiQsBwKs1L
Dsc1PtM1aRvPkmgOE4HMRkfgc8AWCOXhKlwA1poFbueC9zdzfh4DPBEBaNeJ
RXqwlkOYts3Vof0UDTfPy5UqrvZ2QvmakNG5L1SiNqcOMiXZ072qRqI4rVOb
XCjdqZyJdjHE82XAq9NMvscOAsedDWylXpFxpZZCOoDW1KBmTNp6W+MeUw8R
QccUymh1wwUzSYMsPE+s0QuCvRhpAL2W8tSBRmU369XVEW6pZrfwFuu1c8qm
C3fPEGfheMhFU+y+uggxwU2lnTXXq56/Tm4cuYq5HCmzL/1Rozcd8E0CN+7R
8D2gEt3x1zTEy+c1UHc5Jd87tIEz36U5wQazflxCdiuft/GNBH9e/YOhcmO/
fCb0fOOm/HHXw3nNZc99wyvejBfZi+7AxOPBOWBS7zQz9PVh7adcJsBf8ZkX
ExVQXAYK62bk3jHWDId416Een5JnaHbKl72uu2zCwr1QXg4ICxX9XthSyAMS
T1zPBgnYGK3pLVhGtgmLHaDjGm60VrJeWBj4VXFzHrhmyyLTWmwSd0n60AgC
8TS5F/K8WnWpQouBjKdGNiKhXV+Wr2SeiiedXjKzo/3Z1s2MY6F2ge2fgS8y
p5Cn2iteqPPX2O5F+arpHerroeEPx10AD+uaADy5iR9qwv3Jk/QtLZfFUC2E
+XcBZlkFmfeKa47FsCY+tNKEk2BJpi+Sm7IuYGpT80w7MNI3GHGZnyJZRj3V
I/3GMG5MoC1B91u4uQdeRYAvxQxanqsby6q1asy/eXB+WlSPEweDiuvRqIwU
hhJjHf66exgvXm/g89cMg7XLeFW3l28wqKUSCsap1dmvpTUSkcSK94KPhRKa
Uzp1+K7XYAr6cGRAz26cdS7RgI7kLQyWUmDcGfRQ4Yxvlp4qfpRdeYO/1Lfe
mnCuCWkA/6vlD5pXtK3ND/jXabuBOdJcLFszmsWzD3KG4bHwSZpdudSwVLlS
7balwe+IFdVS5cFGk2x/NY+8mJeERdN/mtyKMVvM4b08oOQgW/w/TvWMcQK/
egKBNkdW0DgCPyk6piEh3eJ38us2h5H6MW92URJta6ayI1fWg1m6DV68axd/
sxNox1mC1r18GJV2PR/6MrC7T8zN73++0rELsaZpLoHj6/3KCgs7WlTS8GQX
hx7yjrkYTKz2GRDQh9/uUcaNkhee9/ivQpQhQ5gXw3soiJvIT88ayiXG2l/m
EmrxgTw5ZlMjw/rws7mi5VsTcMHIr4F2+ZVYbM226ONOxDvPXiO0K0ThADjx
bd34/xSqf3IIWqSyLEwrCdoRu71z3ajYBcVT3Tb6qhsbzbSR+1HMmlZ8Fbg9
T6R/F5yo1hC7zxcJuZt0QzhkErt2PIY01aYTtXJR3ieQiZasbLp2xogYaIw3
vH+tfjnNnx3YnSfQ5QSDqcXbuVLFjYROXf76oBDGYl7Pkyd4kz/EtHPekIuK
fFR51WFk3gJTzD4b9+0scdw/Szj8OL99QD+A/SGYGagRBP9Jhu/9NhP2bILE
+fXbzHylj9puTZkxFUChIDoUi87yySOwvHVTVuRT7bbiDtkPPtQaYOAVK1p/
pJdCPZ+cffehh0kHwViDy/YlHVKu6LWaj2TFAiM2+X9lFBsTuC+GSPHeQ0ey
JgNkJGCU8J9Q01IYVcQ+Lb/ts6dw3oFCMwHDHSaAWbKNx9ON93lRuuNA8WWk
dhqv2yNORepcjWskzBXQzE0XpuSrwfOoLJUDNPEBpHGcC3cl6lcYvHWt4TTj
2zGMh4UvCNoW7UYUr4cvM8hScpXDXTkr/masUu2K+dq75NJJUj4V+CanhfGw
7z8MZCPWoA1kXAvDV1VzcuTSJFY5ulZhSu2h0Zm9dhrvq5aXShoEzom1V1fY
inE2JJbHNTr70a0FTG0bxFTfN812foGYCSioUmlEne092jsg34v+D8bk5tAV
cx2krWUxIkYapkdPIBufmIFgVy7nds3KMrZozUiGwy7VIL1qLBLD4yqK+vWA
OZ8LdnP0mUc7titn0eSAbkrBSgsRzoKGa4yAExEnYzuThTwE4u2h/0VjqSSn
fWkSEuOqmizVouN3aLtYvfXjHVX93Kk5wXe7xZjM1IQIvLt5o2NSUHJcLDJY
oRv9HIz43cpSrTqzWFcV4Rg/K4qemFfOVc70P+SFrk8e1Nn6855YvgZhZkHg
EMtT+PfPK4h7O2B+r8fvAS+7O6r08AJxr5FEFoCQ8cUVj+T4ITpJLZhBJJMO
oCjmTqr/AL1GOVdzCwCtOsh3Kkwqq4yO4JQl0YHq1nFhw1KuzBG5GzLakLn+
p/rm/Y7azhRNKfZi7YOYZHx+2KqQLKC9hNIIzF8K88BYtSQUBtepVRlYQV4Y
31F2QKD1kcvS7nB1bFosGN0ZshbMmc2M4zG6IC2IB3NlQTdF7sJCJVH6BX5W
lpAoTh03iQtelx86FOrOJQhqnBJRAzZx7rTms8h5ArsqnxMeILyL2Wy6PwYn
Z8sRlS0FwMUkpw3vr0nl4N/9sLaL9Vei2VXbbpXYArER8pA2OGhCGvy4pXIQ
x+FLatbgTudkEoh+Z690DiOj/KfP/yFhLVEcr7ANCuoSTcmGeysYgg+ZMk+g
p4FJS394Z5n3WclEEjzHo9i3rJIw/I9VECiNJGB+djYk9/Xsopz2rNVOVR7g
umdO55GhLAi6KJVru8+lOFLwFi8xmQa+wY5G0tuIkA4U4ob0UWXTzxcSsXXz
+trzjMHmhyGyPo7W+7IAC7pQk+0F4jEx7crilhzj4WdAhlFPCHJIOoWy9qQm
QGZV3DyJjYTbnQNt3Txtrh/7CSj49LjbdOO8I9g3B95V35CedkHplIX8mE9C
ERmiByqWSPurSl9L+woMY9XLSUn+mMfa3cUr88yhmb9lfiojo715/24jBqeT
E9VxYcuXRd4jrek8RLYePwnyzKvnhHdekbkdqrVkRJg+8Oo02YCYd26Rwt2W
Il1UEaUaveyYfo2rS2d5uhxCJjJuz8q89q0V6+5zSjq9c9kP4X539uMwCqgu
/VC5EZVd+Zg1m1CsxuaqpAy3gAaHMmNbrCE0Dq6xPRuRT1P/LPE3n/NHrUuh
jd6FjEyILeFBM9MxL+tyIKFSMPTcha3r4C7US4EomoSKix2YC7SDwCpa3afa
S9oWfGyWg853AESX6xtK4cNx8NZCsFvQrUWU9WV1Jl93fb5yVn1nON6MG4wm
5Ss2NkEBbf0pEhlhC5p/fqRb1ncYc6W5tjCT0sYJu/upAqk+WeSABVG1k9w4
cr29NSQXuaJrY+6ASrhUToetbaSxQvxalvJ3qTHodrypKsDz8iK+KNTRYEHn
Qp1KqK9xRogtDTfWlzC/qZMgcrnv7A9fzb5A2spvD44I/qU617A9lTUNlWyF
5O5XQ78H8fjHXbpGJF+OeCAsUG0783SRMhJwqWL3+hK1xn9Fv/9kjOhQlU80
zbqs55iCfHtl0x0LmSHUjKDR6hRftAoD2F+/lRfjhbqFQY8yUDLYv4sgN+C8
yxVm+Z+j+hrnFKig+z2wHBCzKihOycTHu/X6cTGTFwZyNXDnqRAMiUalsLiI
BhfaejMVGYTq2Ke+VqLp2qk4BXTUiRUAI2NVGKhwN4C5Vn+vXwgBvz4s7O2a
csR8M06AnWPrNN819b9g8uU3/WsrfEYSbnVl8k9+11P5s09Aj8FzeSE5uX2D
aX4ccN62J4amcmifTex0cvK6E+EeqkFQSWzAOPurGdiaYHI2ZS7R70wRGbFY
bUoUO5pa+o8a+ScJ/0GW3tf4C70tsYTwUH49bZqUSICi2JgswpF9DML/DT1P
vZbA5HIf1wkuKj3704xw7v4cuWcEI/M/QqIiuMVkh881Y0Bg2mbu5cKyeUZZ
ewPplsCa04LFJIFTrb0silOTt300Z+3YyYZ0sz3voYAoNEHhuxALJnPCmRX1
ycN8zX1NQpYAesknoUf8ykS5o7hXnTlkxQ8shWjUqMllnIhnVVOO8/F2qI0t
tiusp1Slg5L2rVY8J0gFH7BTn7cwBIcjfn1LB4sentKT9SLXrjo+KMp5j9CF
Zp7D9oBWlA7Bddt1PdE27OeWtNFaJGv60wsDsSkq1wv7fxPPYUmZnaBqj1tF
tuZw9iybkmHJoWJ6IYMiHozRXJj5j3nvXjGvMJl0BKKZo8GKmybwQz8vfgMm
LKdk4TMWoO6tmvCWdNbk9UZ9XauP9YaVGPdZPTJt/M8Pi5gJDp65tEJw41FH
VV6cqE7iw48RJ+gEoAOcK68d2U3qi41+qAn4EgiQQEITt5QKxgsb9fpsH1nt
Zce9jc9ysX4Wa4rkn934T2gK8DQFB8PApWiq0b9h6n6IuzUTdgLesfjdD0Qj
M+0u4z1HxlcfhB+vsbP+jMMBDZL1dZWh0UkM2Ec07S5SKFciKM9CLmDY8bWt
2vKwvRJzOzSNeimFw7asFrllYkKyurXOhdzv/zqAhvA3rdLtDhTkHTd6QoYj
9CpWwbXSZzoufrYX/Qyyg1OgrbNlikmL0CLGsVNjKCL7A3r7MbBLRLI434Lm
LcfneZ9ihLNhKgp9f8cLD1zr+4PcIuy6xnaNvqgsZ1t9qap9KC2WFoS92zgf
8/rTzG0qNJZj6PHnJyAIGGgS2wMNw9Vc8YFEBQUsk/5sYR+FPKfZtB4JIrmW
l0vBSF6hpfKO0G7rXr+7WFjuwowQrO6Npv/t2MOk/OpsCg4mmKG01V6KzEYr
SzkkH2swvrV0o4XYWxPRAawdhM7mu5ZyqziYZY2GkmvfpwWxwFpCvVN4+55c
piZ/kuC2giEoKo8U/Ckyna+Ebi+EKVDRAGDbTpzBPaZSh3N2fXto2OFUNRl4
98T1QZmr3TFoowh+QFp1ZkFPT6HM7yRe+Bx+zjxdIzYQWNbJUMA6E02Yx1mg
bxaa3/VTySNpUI4SDpfhEAVrg5ndwRaFIMY4UhStIHkEDItttSrbSBP4q8/D
vi43UiUyeUB5lqeUGe+5Vm7DUj4jiCJwmFkhgfT/afUuR4pCd3hdzFhXbk+9
aJZqB5vksla/FiiiFXzxFxhwg+CzzsCfsvTHXd4qD9t7I68bRa6VUAx7rHTa
Has9jXUJT2adYIVnYtbTXYjNPn855X0u+J7Xtsxp7G94LTVQmiMkfwbC77V5
weW02e68kdMhZmJ4mdVkfIVLEsGx+P0bN3NO4ajEux5spcvYRRenea7NNevL
r8grXoeQBlaDMx2EyAo0X69IsXfTXDB/VPY5jB1T7xkWwWBpFIN7CXh+0iOk
ep5E2rKDaR67YrPXdMYqzV9zb0+MU6BiRY8Dm1vADUZsQ4Lk9MKEf9C7JWBy
Yj/YVKVXU5hOfjuf+ECf5UkxuzTMTHsN96t5HvWlmgDZSTgvua6pNxOhcDDy
t/Jz3ckRy6pUIEveot+K4c5BzMYyl5+LLJaroy6TiY+zuptA1xvwFRbRTUy3
XmqB02PfSO5UWXoB9SlQdgvEyN/2fqi146RYU6UwQ7n71mzdhyYgrJt82dYh
/Mg5EAkxCvI9zTcUh1ee0SxgscalWlujJPr0QEAynUL9QEkzP4/oLB9t65TH
f/gBS9x8cDlhC3Uf2g5HPsNYB/6Ak4/Ze8yo5mu7dYJ4DSt01i0u/K0JOq0x
KLkLrr8GdmOxUiK5ClU/mTiikGKlYv6yjB7UcdHRSLPwYTZ1xHR5J9+5roG2
jAKhz2CzVp2Jlv3z9tB3DIe1cZxmuNEGpStJYZdFxfEbtVtfvxQClarzNkJe
E06Ys67XsrFWp4vhsym7BHBIGC5SKdwAnqunSwtrG51P6/aL0cGBJzP1oN49
60TMZGxLFR401JBaSSro3XGHl37luDk9h0THhNOrP3odS7S8TXNg5G2kITOw
Trq/sjED1QtHUvT+Xd2MIlSzHY4k1XmbHBLHeOvQmK7O8uUkTwK7cz1kalEi
g+96uGsOyE0LtjSTy1I9h/woOcKRzrN6Gw5bU95SMCC9CQOhOFjvY06z4yo4
VbpvmKCyetsN71E9CXd6a2gZnTbVBhVDOm+1F2mqhuhgepRKqqkith0ruTAm
a2eoOYOSXgCLO334w2yd8eNsAjKl8OG0l1ymtCpCcyBBUZd+BCXdD9X/krP/
/K4hbbVadvnVUOsHJFzkdxoZhE+PqH58oL93uNmT9eECYZ7zcKIeJIn5b2A8
rLfoU6NEE/krJh+O64mP2qVHTw1vqSthIGWja7XYp5vB14ppUxjAHgu9Gh0f
3vUckL7Uq375mj3xscXTxMEAkCRxUEuyTC8dVxgt0t6G5WOOsKI91hL4/2Uk
eVPDcR3rwW1YkLpNI27tC3WdH2pbtoyFKAYomDu7qgs2NF976JuDsU/OaZBw
87IFudU/5GTc8aEYxXtR4fhAnfjXSmFKEDLHqK9sMBYfvIs1CaEdf0sSps+g
wcMyIapaJeKygzyqK0/G6DwcaPE/eDV3cuuQlers3TeHzDdcazLxqXgd+Ybw
1yMI82Sr52N/sQhmlikY9jiQxT519JeKqN9Q5LqpjyHNOUMTKK1lIojoFeQx
3UrxiwC0Yku2OlauZL3hXguqUCjH2wru3XqXPZAF9Sgj9QHpyabN9QU4jYsL
I3CiD6Be+/A2n2cOVOFZJdPrLR6Hk6bUAjKzHMZpPSaabxhTzOAKk93h/q1w
xh46LezS/mEQHWcg/pyde0+faf1WEovU5xcwmCKQv/VqPsE/dgU29/WpYp51
kkSVqKih+KmylFDmLAD6B/rge3ANiDwIugWJsBD8ErOXwOpHh5hxj4iDUZzG
rXqy8Kt/p9QwuLteqvfvRctXWjJF+8PV0HCYoQ2LydhJXcZXrOrW6YM0W6VT
BNc9juIrlqYGJt2bxLMvaA/M9BYYqVFhIYBNaTjl3O7yxzvJi/n0qtfzj+d7
D0CoblQ4kMRj1HpJlC1MZM/vr6lH2Ct4arqDSpANRxk4G9Iw0P3KPW/HTRbA
s6ZX3jjc8hsX7DMvjB3b6gU34KkXFqYxOc6fUf9FdRiiZRngb1Hb6yFUJpNq
MGr4zob2agp5ZShMan+S57VmDGK85ollpNCpTMQO7XpKBn/GiAlDgLtzKGqx
FufrbBjPtOPU7+QUJJ0uV8g1NDoQK3pOgLpBzgR2jvkNlgXsRh0625Y9JukN
sOxH4sAeWoFLNcqjrUhEGvnPHV7ZE8uXhtr+8PBPUos1s1oS9rmp/ATEly0U
3c8DpTPug/klEKjvCScsRI1iMKp0d3OoTYcKwC6lHNm+YqHV/38VfEcge26u
Ja0KuzJzYYxX12J4UXDwxgc+gK9uDcM3iKDra6Ki3FrSozqt+ptd0lAG/+ge
QqfVLYO2k6yHDwPweqDt8lznQf4V93VUGG+PbGDUtTQRa907Fy+qoYbM1rsX
mrcNonLlphXp+lXfkPvJBO1KS8tQduTMMYfPTAIznDgtCMn9dNVuR5pjBnaI
d4kqT9bgLAS2G+ls/DzCYzAucwNdulHDL6uVwHCs1Ve29zIVm32GtIPEVIgW
DjtmzebZ2ccgD3sPBSoFbeYgWRrDLPLs4ZGUQvBbPEF/uJ3Gsuk/qSUQsgAj
ZmHZf2NJU8fH0CLo1xiplkuj83/Dm+jIQP4qbW0g99EiaS1yBALU3wcu5AOK
N26eosu4X8po5Yvcwwd6izWOL0COd7EKQOR1RpOPZFlmY4KgO8ftayyiHfCH
iVilbvW1Luq+2lk8ePnv5dq/9u72Dhyzs3maaHtGGYMzFvmZzDh2Q1MfWZT/
Kr4FXH9EupEGtJTsYSW6zHrBnZu+ZGE2XNS9K3r+mARGSa7eF84RWT5kOhmA
IqX/lop0gTl+i8C15es7iFCyqbaQC+/aEoj7jpshowfmEtXqOX6V/HD4T1kS
PPxQabQK0CIFdzhFLqtJFyB4opgsxPPK7/CNnhNleUelyBznUAafeDUN4e+C
Jg1tvyEmLk6lhQRa1Q841LyNVpKSFPT46YllrY+X6BH7tCoGYoDo04oOQVFl
U2AzWKQc8tVOD8A52nNkyLVvIRCpDQYnwvgUOHXhtL3bqEXiMojkkzijWi48
D7FxRthLT6BLD6iDjEIJf6HzJWYY5IYSOCTP5QL/IG6NsOoxaQviE770kgup
E46ALBjT0VpbUXXcJG/YiSgbRZZV1mfrEJwOyXC0vAAyfhPhTALGAQU6YFDp
xO5S5jcx0jE02EguuysvpX0AeSGdcQ+mP8p0pUtL4+0cqHcuvMlhneiD6rGu
M1/ot67JjRkU5AiYM9t7szfPZulgRYbRIGSkY2V7CuHQH1Kk5R0ki2U0I83i
48ljw+DTQ22Rb1FCouV7KzIW09/kFVz1h67lcsiX7t0MkuyIEmf1pqbFbBRk
8D2hwltTHp31+Equ0fQ8Fu3OizsfoW+0ThF3lI2mIawm9kjJDChYRKf9wxNm
DFYFXqcIePBkV+CJeCskOZuuslgDtP5dTdgfg4fw9lI1NonrQkPsZREj/B/f
qHJA9MHQSlePv0q10KK0CRkns7QPpGqI4cXK8C5hQjW9QL/11OakAG2HJqIT
tvjUwUmgN05eZNrPMgLMNOIuh6wD1SwrooxEYff2hkq8SoYSD4Kj/5XsVP28
7ceiSk67mMMnxCw55eoA+vc3FO/Wr8sBCBRFj4oORXacw14H33CGYDS0vh48
ZeRdkc6V5DOG2nuLVzn9qOXipCoZjdKE7iD2qUeHoEt9HvgyJhsLnvjW1JTP
lmBPy6mWRu/fOWNoMz61pByIa6Gx0JReTVICmPClRNBfzMnYMAI2ekOJlV68
D8LYyYYy9DFTC03zGscG5cwu7POdrbCe7xvZaDZv43NF56hdOqTjd+hz5vWq
Ee0y9F7YKCIVnNHvoGfBFoaEUa7TL9yw2yIdwkBBMc7ONx0mm6GDlOcZYZps
d9ekCHhI2rn5oZOP0t9XeP5wq18ecIlZQrKoVyLWB1o3cYCupKpZy6VbvNSb
rjT79hx8Q62XLIOW2NrCgOs5WyLC+sjO9SGZo4Uyv7NP7TaFZqWFjEN70nJ0
Z/h++yZciTifZgK+ZHH37z+nbYOLMV7rWhwv8KCiHCECgvU0PM/62w/w25oK
rzRiq782vEVwgoz1WOwGR52q2mFkstKlES73gct0mQWS0/MYqwdUUmH3pjdM
y0HNrofvODDf8SyxZvRTHqnGSZ2aIqnoXeYwUGcqVkgd9Pc06ig/f8133Otu
CB5IMgJx8568Bh95BZyWqalj7MvOmehtbeRqwtaa3D9r+zhacDGmKiTxcwzv
tUWep7npZyZAbuE3w+NbWOy5A3HsO6tdX0fqFYlmMDADWt6kRXiHsvLTyCxV
HaihcrOJ8ix7S2I+72txvwGU3pP4aDDuD3e5pi3GvMEl95tuwbMEokxOO3zw
793K9u/sKOBdIpx4jA5Y1rRyx0FISeutLb/MurtLB14WAkRpJlAz7LXwrCDu
4/92p52yjC1Z8IkB3gfIyP3AT2oLcboH12Fo9ArSwOwmG5gQmVxKdebT6AQ/
HOG9URjfec81b5bwK4co7DpgpF0Fc6Jzdl6m8t/NgLNWNtbf810BpkWBvURF
2f2fi7MyKOPJdAM9AxVHfsk9LA9ft/oFCdlAKNdbhWuAZJ36u+kXdt0+xrMl
mNGHLDxrtc2tY0B65KPW2PASokKyKHxZ4FcPocaZ71ATQB9Tbn9HiUQgdZL6
EWNByvHo5IJZY2PuweC2WYh7nkUdTunubE3D3zJxHZKPs0awsrlte5qx/beJ
LdmS/aIlEL5HNvXcy92YqiSCoGykwJw9Ko+ji6ZvvcAjbJRP9SyrTS3XSmWa
zrIn70DbQcsdVELYxgDMs6qccIkJd7lPn3Owg8uFhAr1g90H3w3vrXE7HhdT
Bcd9z+TAxzDBBtxjTg/zPnKinGNjJrm4Y6G04ZkJR+WWtWVr05YKOYwgNjW1
O4xcyL/ayX1Sg2sdlpbhnISNH3paxjCj1busc47a2MpFuPAVEsTLmsjJFw1w
txoajVr05/kzXSZV53NneWM5JN7bu0TlAq33S1c66H2TL9bn9rQ5n7Y1T3ZU
y9cWRSPNOLAURvttEcF0YlIOqBKtr4cLxVvFtQPoJdiL+ItYtgeeGFMKVhN5
wWGfcLwXCr5RXp8WC3sEKgOhW8eAIwNa8yJxQg4ZmsRPjo5bGE7DW/jyjxbK
XenNXIaZ/ILvEibbQz3EH9kIKj06W8K23I/BhpfB5Pp7QDVhXZjTc2Y98ICB
8wSrjcEWhU9NNZfpE7qUOHTtAe20salp6IDEAfvpvjwozqnDGTorzNYCvDTC
Gz2l90/x+v2ecG1wJF3LGSVQy45MYRIyutCOT1b7uuqgqwBgpzMZrxhZTaUk
9ZUw3IMzOQnhL593VnmABxc9GJ4ZErkOUQ57IsLYRlQ5rtcIh/Pw1Ratg0Cw
KqYQFHLF5fVEnTdPrepb6CobkjTcKwmrK/emD0GI5/2ypFia21yNXGRE+HCB
ugJBBUYjnMNAp+q8PCMLqGBICs/2X/XRw2s31GD517rZ6ipDFHBEkHmBHdu7
+kBbVpYFtZDjdKhGw3UGJj4Nk3ayC7dv/GolopmgMlYXXpFl6mMn7jueHPbX
QLmCqQdaf1Z6GKZ1fsL6g7tmFRPhf8F/gNe1MmmNauoQirjGkGc1vYHXK7dh
xp6Fov17alqCrc7c02kq54351K+I08oJJbybnP5f/JbO+9zoAvMZ3mFiYc7z
cAiq5+1GDN4bz6O5b3XxQo+X5YDw84aXjZ7kVPrX8DO8a13aK3V/mxB1WIql
wZ1asOKJewjX7fYCq2ewX1PNivlyxIXxmZxATt/ELvwxh9A68AmkrwM0DrTM
g7+zvxtH8RA8WlUB69ZHhsnlE9qr5Q1yX1GEHbkj2AsnKX7+fFuFBpqjgOKq
QapxdvvScOFBJe6Wvqj8Fj6cwlIhPUMsY1K8RJeci771odK7qchO0TF4exbQ
QWAsykGdOeUInToFBONW+1paMg0hm/ILIMBZRUQfiM8+5tCZdcFZD+a2ANK4
0/CZzZK1vqUUrTNUIqSNOUI6PjyOIshqbLhAr94SN50DYa9yk+/q61EaSdam
G15tB5W0r8wzjW3yPbqWbnvMV1TpvEXbPQ6l+9oyu2yAMR7kI1YXb0yVQaFT
oCDdLT82sLCHov1xbG9or82bWT9YGg1X5kUO8Qe+fDctAiiodYUnZO9vl6MQ
Qq0p3iJFjvQvj6hEhF3rQsNvH1lcC/cbe1H/Djz7G58Nqvgy/6QOdVscEWCy
BeHBhvxox40Kikv4OOhSsXvIeVqHXy/GWXxc6RtaGnUq529hNygdVZmEtOK6
aS4sROtx/nX7Wf0k3ve2Mx6KC7vAIJ7A15MlVOKvRLhCo/5oywmZEZEbeLWa
7M3ABwPPmDCMUya4hn3hp4usav899g2cmIrSdlPPjH788JM0lqVCRBKQU5SQ
Kg5Ps2N8XAB9qwOL9I1QLLfFSRKX9bDkesHQN7uRUsmdEEwchgCv3wv0hvge
NgH8I4cACJ0r/MdvBsy5hq9mZnVB6rytn5G3XILa9KEBmHjsOsAkbpcO2V2B
ERD9VqzGn7B9Miw2UcCeOyl5XNBMrQUyE4IIm8pInYM9ww/AHkrBDUUd1U02
aEqwuGlnKPVYtJaoVegbEsp3BR2uNl3e9KxwRcM3lGZyBPXGLup4lu1ZFCWo
sRcgw5jS2QX4aOO+GtTqDv25A7q4rFFYYrO5qhS1rS9zYhZrqmThM6sH/mns
8Jj7v6iOifn/lK2pVWtqS45fL9xolSMqBIVslHOW+K0C/y2bFpyzbJxfHaZL
trJQmJnNzMcflRLdKooM1y8VuNA4/9JhYpL/idWMJXP2j4u2hBOdPy3HIN3x
H2cEaY+mESjpCNLtObUMLR2sFe+vW/DuJENWH+GssEyW1osWVpiLouaFL1Ei
R9Z+1lziDXGrrmGXr05dkIMvLX8kTfX/dfkNkAH2/adjilrihHUjH6+YGSui
2C1KEEqNSI4cxYT0zZHkFyGdwfzzTJy4ttH57kMwUyqYprxdp0eRIPQxnXnB
p/ePFGMP+qN3/VInAHRTDLlghFi8954UFkIKz2ZuHoPPyj409SS+XkGtpvRv
/EBf1E8vB9ApZUxjV08HQ5+o4h5uq76Bxeqe8cz9VJ9SWVF97qi5cQGPvuv1
9/KCvFE90ldrUrfRK2lnmNGDP6SFJS12xfS4p332ck52mjoxHTWDFuECc8nM
NfcwItwTzjIyPbETv7opHRWWQPyjUtJMzwvk9oAsGJWJOGH+aPXuLmsXBpNt
PCTd6hWIEBdTG70ErXDdFy+spIU0wcN6wXjctRu8FMp0WPR/C2czlkcOevAc
8el1ib1AC/sZXxpMEIx3OuaYL5MRv36WFauf41wl/a3BaYnnX0IX8UPDJTjL
dOqZN8DPv5e43UfCbVp3NZpwgk4LS4U+hZP/9hC61SgW5SGlFCWVDtkuI97L
ZMadj3QUCCG+f79RrpJj2Omhvt/X+zepBAuzmib7JSZK520qi3oI0tkNvQ8z
JPJQHc7s6uUN1MDSvr6yyTn+VIpgNHPXcyxDbl1mkcLFriavioewGWk4zrjf
+aelk6mfNDAos9gPRpPt21WoWJzFNhfDKAfFNozm0ig6IOORnxWKOp4DLOsB
hih9kTYCTk28RRb/QdP1j0CtneozDbAXrjGtpDjZLGqgTNXHmHyJUvnoT3AM
JzKKCvgh3VAFkg7/WWnX1HH9QFOSv8qCz+GtWHIKEtbt6nS/2CYQBpmaLF/s
SBHvq3Nx34wRxV5HnmpwQiOVXJiMBZfBpq5BS5GJBw7lnjr6kJPTmfPMw9Z+
oDiKjnb0Yj01BD8s4h6UiK0U7s0rk9uxXYYLpcnNfBT53KuR5fONQog4Jx0+
m1c9v+iLKMJXsOfF83yRh0dNWNeB1Nw6UVAXM6P+ZE6PzDFYGdfJTXtiK5Kx
fgoHX3dx34f+1TLbayNOIQjIvQSllArF65jYTyH4NJRNLaUsftmlSGRgrZ2s
9wMjyKnOitrWwXEI2LoH1wHWWlDZBCmSUfGoo2hJ/hfRIgXeJdU7gRSraElv
GSUGiBVmC1yHUeT97Y48PHSytmr7+XU1c8Fenf5ZMlHqmWgZnhErtX1lTto4
w1liseldOqgyXnMFp+7svTd6KcZBoBVgM6goUhVCxp8x9XDTtsv6auAAelmU
5P/tbvLDSz0/KSU1qIOkDGQs1DT7o9rdZbGio1wHGNGJo6ou894t0KxZ6Ou2
zJ2ILFklMvUwgTnEQ7knO5dK5nIVfZA9pWTIHPnqh6WvQcjwZn44bluqTeH8
v1AKREvNPo7bG62/6MKNncmTuDiKaNbDiRMby39G0eWwot9kZdFYrO8Gooj0
BsdOVLQOnhQ7u46HmmVPAAiAuGDHhnTfMMaSZ9aTQw4QSQq4PhKd+vYrmmDW
JZEwy6YABPnnHOKf+FmEjxR14AiJn67dAKJXSDVHuDQMSaI4hYq0+16ZJFTO
HUEM4xgEy5OkSjZisU7aTe+VoEjME8LPQvA26HJBxKtwywth44+akM7Z/LU0
zaeI3N+hM7k5IIiZ6jjAgMW2Vk0SwDKs3KdiT1h0KSMy6kufuHuWrMs7Oq4/
5EJ6LpMSJJ9vHWDVy5Q+NlEXzdMf/boBh71LHNbWlql8QFIyB1mQQIrjOIb6
aMnagZ9FqyzqdfZHHCdcq6rI2fVscsKn45eIjCkEUUHjsa3NgWGFyXG3R1LZ
OlimgXRCKGqZFWJGbzzqi/u9LvJvEKgKIt0NCSVDns2wMgCVpBohNBLO9qtJ
7TcKD65TzYBSCgRk2hv9MDxAuePjQbqWbxHM+PlAJ0n6e6UNNNW1fEpoVjU5
H43bHhVCUKzAeQrpWLPQBCLCFSHFhV05wkRGQZ1tBB1pdAE0KlYFMQoHu51W
NM4TEwRLWdn2iCGuOYmgFiwoOQuOZ+jL8Mqb2ri3JHkoVkTc+B2MMbGiQxk4
lI6hF00gnIZdU8NdT+xdYLEVxBsvTm+z51/Zdi0MhAEdZwKzkGhvwPkg7UvT
r0csczVMGkB+es/dxOMJtGU7NY2P9TU+KkyTb0vfb+0DBblaNDGOg+JLXuR4
Aeih2pTkpWVfSA5+uWBc3q5azm18H/hKNw4NRal/7toDmj1j9Ad0Se8VR8HK
1KL5Q2HpJY3aupd0zkCmY/SCjahKTyN6itgbLJZd4l5vKWiPEinCy0YiEn05
9THMEk7KtayKy5obyIa1nsKm2PBTq/0W5A0EI5kCqDl8ddOllvXK3nyMiQiu
iyFGh0+yyHyIir1w/drnniUsci52IOlZT+Bt45F5dn27+javqUMaSl9NFYcr
d/LJg204dIrXM5i2hSyx3tO7F5NcgUhQstDhrdHZ99GPGUdW1d8ABKHB+oIW
rJ13xGF/5J0qoMYZX77VNU9+GtdFPRjdUk7BIykFwWbCa5LmvC2TpuNE1jqN
RpB9bE9G4oVS4zhn9r+ID01hWxH8CO3gJ5OYrQnMdf3bXZiOXVfp72GJQzgK
gsNmtwEFGRPzBdd7yEZRC+0dllXpjYnNLpRx/3MyVmdk6k7U6qgiudRSpY70
gMfphsZ1n/6v4k4zzRNr5lHXHx0uawyeQYxjxW92uhBQxSGda9oLH68yyREm
m6Blixut7OPVomAKa3Y8FrafhD9poEbVb/4vZ6qPvGCBWA8eeyBOvzM2BPUl
tdA7XuCbiyKTifm8xYN+Ae1j+VTMzZnPpBIF0hxcgedM7opyMqYIN+WGgIWN
H16GhoqdHfi6dp+NKg4eAjqMfyYRmZotIb1DJNb85fuGSMiT7/fjLboA0CCy
OfDdJfsZFkhL44L6GMxxzBOq+RB8AYZB46Z1infMESW5Vv6eGLtWI4+k7BDw
LulTSLx1GOp9DTfOjj1wYZ5SmG4fS1Jvee6ZWb6uZfj2xNv+IvaRMwbpRCdP
Z47Fu8/mt2GpT/Ba/Oiw95uLJAXKzwXwtOw+l9HU/77gRdv2Cvj1xwN3cXDU
F10DDXqcYzl0DlpO9/qJb/Spf36K5jEXIW3dKRkwHa9CRXSc2SbByl9Kwxk9
zHotS2CBltfRBrXBTHgOyJcBfFaRxO4akeHyjtAQXs/6PKlxR+mDH1Q3xk4z
5AJ8kEuB8ySGBmM9CPk8ESdloOecZ3tFXwRbyKMUhJYo/mjBgzy4dd5hWCfv
3HvLsD2fHvhTyQ6cE/qW4isjM9+GEXpadteyeo1XPMnZuO6kD+OEnnA6czg5
9vGHAn+vOojoIbWbNqC/SknuhnxZZg7IYOOG5es0QzxXaRlIxUWycabvLTSF
d8VpXzWPdDgU6g84W33eZ1x/RoTWNKO7GGOd6dzGMYl94WbRCZhuOr1Uzvzc
P6q+z3RiznMrooRbZqLeNQU+3Q+QnRpDCOsY3Ev693dIOF7ENkow/Inu/JTi
uLM13A3fETbgzeov5/b1L39DEdO7sKGWkYrevf+diIneNGCktoSwC8ZT639p
0dgXoDtBtggaN2ZB8t1Zah5GgJLjqf4+b/4kcZiU0yQwdGHIE1Y8lvgbcS+e
towQSgJN8I+EnI+7Ug4qFk/XM8ahmMeDV/uhopLErOxVZMh0IFm1sCDGkycz
38vo5fmWEBZ7b0mXCxozco5DCRmJKIUXScswh4y+7a1mmZAxSHybGW2i24/h
xZ1QnPQ7bhfQeJdUJSAorcr4R08c/PMXC6XJcddmkX7b9msbKuhXKnCE1tnf
jWIpTp4Iv9i+AxRWVPyjdzDEEhi7xEStQJetHo2LTwvL98/to7VRxZq/tCLJ
0nHVdQCgFCRKsU3xA2Q9pq+iX7dmtcPyX7SD2JKOpziVtpAfcqKBGdhzdVhJ
Qjxtp3ZnqZdohmAdEdpmhmKnIf9rfCEW+m1Ra/Oxz3WYURz8G0sJFXENEbas
7v35UMKDbxuYTTq23Dzj+Xl0GRNhrP6Zb46pXNMzBec+0XBQYOnrSJXF47Z3
SLpJ4tWx5r62d5XHFQgbC0HtyBqNQrw97iKI0mhauYlGyBAQYRjCOmOuKUHQ
Jh5kPeElBRT2a3igonMRqheLEx7yiPDRRpEUKT3cWwe2eEJOnH6MXEcWktlA
zcOtKaZfRwXCds0AO50Y5CZKUW2XNoekCgQcche6zPhkU/fo24R5GClp1Pna
sd+NNtI8INPbwKifEjELi165K26s/xEVwEcso9jHwgMci1uH3lpKYCqtzwSw
wAcg+otmHyeBhwt3IA0WOtwTmEiP+zZSQq6J+PZhBF6r/c2P7Dwc1isz0X1f
iez0zX+GxczTpMPh+C/LMcmug6MOm0a/eJgNNop0CwpkgBOKytnjyL3bnnyj
9lvFf2dok0lrAhHI4tZrkwEWZC+w0wmvC8BU/Yb3RGHZOC9KiOiigEkP+ml1
CZs2c0O28e6vKbMA9Sg+R1DGSwsndTsjRxJPpjYQdscNG59USxCn2bFrUqDx
56D3BoXUiIQjfqOX6wXex0alvxxdWbrE+4HzagNAustPZYKMenpkZcFZ5rhU
+mrivcywopuExqRtbxMVgyb7tksq/0hzX9m9PZ5VF4PdTQFtQN0nqid0RFRQ
ZaBWKUNAkgzlHiB2vclfD5QFi8b4fN//kwukv8w7joTS8Z+UHPUMJed1QCVn
yATf3wID+rGGzgfzuVlVICQPRHC/+E6b6nGmnv8zKLx5N4RNSl7GsTADe5pr
bg98oWXZEjo1FDkPGHvlWMCDv7l7TsJPeuH8Rc9InUGBNwswRTFRhNY/QpGV
9DibFZ4IRZccA1y7HXXHHmX4PLu6k1mYVaN8LzWjlW8buJC1rBIcMhNLIPEc
XYeqaWwvrzjK+3Q4+YWwi/xLrWYD8ei8OlgNo+AaC4eNOrnBpHc830htRQVS
JYepTYfLsM0yjNPeVixxL68cyUf9fKt2cdiNGijux5VqEMIIGm3OP2GU2pe9
tLS/hAzjIUsYP/pXcYl2O07X98IMhXBodXLoiSooH0fDVXsuJ5ISqLGHc4B5
eeFmVSQ15FuoXhGlnsn3GiHz+UEXryFrDs/e9b6LaUiMb+JV9RJ2HfSuUzj7
hPvyTAoyuTTx7Q0HeDmJI9lBoh5bLx2zTIvxFmZsATRqBrGwDWuciNdr7QUv
9LBju+hkg45/rIMQgSvgoPNwPRv937UfWtmCrZsxgR4YiwKy9ct0hKH2UJXf
zuL25cIlnrmKxDc25Nq+vmXlf0PpmX/jLAVjcHDQhG7TT39KTBYqQyFAy+aX
mZR+BmO295L4jv4CYX5WPtHFWgKkxoHicK8GjsWEEaJsVDT9pZd5HlaDDtU8
kvi+ORjeQfMYkLuGcfkkqgIxOzC9a9rgblEGuNM2QKI8Z1OV72gvE4FCLQre
TXx/oYmfTSno7gJ8oaGrxzfdyhb30M7ew2tEOhRK76VUWWQBy2/2Ns1ZB8gC
6kdsFNS1QSx6EOM69h4X+4UuZa92Oce9v1FRkHUCHCx96/171XmNN0I8mePE
S6lWV9wjhJiIz2muceyI1D0bQ6fp4w0Ib+m7g9Sc5UemK6Uq257Dkah8HWdA
/kms1x/KyJuyG+DRyLAeOLVLlVKJnPieHKixcuXnV1UpJrSf/0uh2lOtvbn3
sfzCDnnMGYfIgasLlGrEALfqAsdkDiVuFWGy3kbl2T1JUl3zOW6sLBbDSaWy
iD+CFBeAuaucQ00Vu0KHnTJCmdn/W9G1AmkMrLLgQrxt7CmdUY+doPiQslQ5
HZKNp3cZ1yiifG+pAklc+RvBCsdENnxMdDs7ePEhaM8tqtwsCCWQjyVT/fd/
6EU7rUQmp9Ty1BYTCs59HF/8bpNA8zMvF/U2iN/uUyEpCTZ7kuhQsATgN7uo
Gn5opagTQPr0+nM471X5t6ckPI/QkPokArqwcvO0Sz7Hb3FV97NbJGdb/Kd1
tGbC1q7bt5hFDq9N99cvU8Z/P6xWoztc/hXtwawcTzFayAuHgGOtN6ugZmAA
U89ST6dDle55ENH6/d3aDbVVGdUhN8wYw1yhBL/0VjX6D1PF1sY9thZTr5uo
JkZ8HTqQdssIz8nXY+dsfjQwEvERN3yGMR1po3x0VBMBrYwUfby/x+HZF4Fg
W/6kNu2/ZL/f9d9TyDiB6r9JS9r5vgjUJbBIZIKGXrLhoN/O+LZ0+IlupKbw
gxXxbDtn2bLMe7Aitr89F+veCk5oNcYDJLx/6zEuIgBkGw5NVkdtvJ0TsTot
kYnigwYJ3ozfxpScTmZc2u6+qPy9Dm+pS46Lz3RdF61WAa070eUcXukQkvuf
oecrjCxA+H0Y9ytbJzQyXQUv29i/h5TTTmiZOMSpvQZn8kgQnoO+uZjmKD9b
REV7Zqw8ppfolz0bLXBJmwRZiBq7zOlCPRjXsQzBAyNhtrZ5/Av3fASPZR4C
ViDi9ugbyU2mBEDCQ2oUf41uuYPHxQ98+1kFcU2UJPGyv3HuCf6gj1xc+ca2
g9jAKzwyqLjA8U+0WzuyUa39BlwujqI7mDHJ5w7H67fegOd5cOmzfRNdocex
KltiXfvohhKbpmP4Ol+ePlqQNJMphIliwxv4d+rVO5RYxGYENJx6yV4sxOJr
+Zh87LtDkXMWbzYiXnyjBe2tJrZg/KEg6iZkvJT3YK4ooPZyHEjzqOW6fTIm
Km1OgwhA9D6cxafgGO0d5ArCWfg0otR8ckh8cG/FJrrVOgwBUpsfAa1SdEiW
AY23qTs27cK4qZhueHG3g0D64FB62y6YbEJk48i1Y2JEiz8qCOroQ0ySEZFv
HnHF+zB6Mjzk1i01hUtR2ahlD62JssrFUj6niifMTfEse4OAryTXLceaGgfJ
ZD8k0MHg8ZwFeF7Ru6KntzRibf9CnTA1fEjCSzgLUSHFWU9rCkORL8ha1hC2
TFbJF6zXmPRtQnj7CEQo3DAOyXzYH/mPMCdiy2OI3Q9g7AKQqXngXmtWGvb7
GaRrq41OMWptID8EvPiQkQBwFTZ4H/BDFCa1NRM4sLzGLsgoa2fRf2wctXtY
eop22QyGmgFOohWf+se302EXocz/wWva0qYB+eKbpdxekamoWxBvSv7KkVun
sh11QGHfUmu2dwjCznvsEOQQt/XccamieIK28XOjx4IvKIxgPJQdfnQ+wnmZ
D/LhI4TWyQzpmBCdjFN6wpBaQhZIAOrJzZyuGIcux1r4cukKk9Vt5WqD9vYm
JU+R2iA0hOnPg34+HCS4Wgm3O5MjLi+30GgdDHXaD5BTbUm9x5I+id8oSNGi
385iq8STAyCnQddj0MRKmSl7sm+NLtJ3F1uKIJUFOfJcMc8hb0VQfzslfdob
yHRsTGxkjdD7JdZ3jfHtLFlMC4sQWNUbops0j08MtXSLsAk4IICXKhD4Y+9B
RayPedbLbm5PwSk7bH6lRe1x7wNxmF+xQh1K9AitYLvTYjqIHxPY20UnTPym
44TKFdSt9uwWOjlpMvAjpdZipbDPCWrwJDQzgDAYx2WaZbG01Ltt9/kT2rlg
ZPRZr36+SOp914t2bzOKEDpDgedidGAW7nPZbJT3DlYKbi031gqBnpolNeSt
S+7GArciMpVSxJRDl0aVVe55beyZDvKtG1nj67+oyf9gbF3sUyk/r3Ttvj1k
CIFnBVCGJ0q/FRe9pKsC620OArMSeRqM3wRMDVpuSWtzVq6ZVEiP488w7tOD
ImW9/W0VYTRPyyEvzVw7KygDzESA5lFnrSGJbnWo8VLtrMfWWL7ker6DjEJD
AGW2/KB70EwJlUI1Q2thPl23sANwDd5t/Zr/C3sguW/kYw58xghNbG6wg4z4
VWlKaHDCCF4GIV85HV4ayqCcSu/UmgfnuiRcY2tpKKW/DOXVIMhjZ47elZ5f
Sc3citjm0nqoue3KnpX5hWTr4e3TezedQVlsxu94zQUzdh3G/OQ+4UNEescJ
yd+9xR475Qu+lKh8LiXxV0dajC7ZrZbTOLr+27TZx2Hz6ryDTW174OnQWl5P
GIm9mTFzPGNr5tUIPWfHZBG1zIDkB6T+IiT8OliYn2lg8795zKF97IrfYXI9
Bu3wyblQgMiR1OdHITi+u7gT7daCA1EHMUTzIP1uFtgVm5/lbZetFi6zN02/
V+ty2BM6ExyIYxbR1rFNCmmyQf+DC+azW1Xmc+PyVr/Z38OEsGAhcAS1QPcT
6RfWd6W0fmawiU7EdXoervEDXWCgeTYdfxHAQlW/a0kBqT7rQgWUwOg7Noc+
xHXKEM4oBBBP0JsYM1+ox3scd0vgcQcFO1cISqLahnpvLGFmcYIBPOfx/Bmw
RxYUOeVA3yBQeCIF8RhTagelciVrQZlzRz8zqj1lXEidP+6I5YUR8lUyJcjX
ZDUvqi7Hg2BgbSOmpkjFR6w/3BXgNe2AnNVVE6shF9gstYjEArjfz+aBJ4eY
iGxWNtVmEhLOzpYyD4nbGbRosCHVsHT1Ro+h9VtD0CbvU7S3lqkSV+CSQleI
7v9I2TRz3n9HVvF84mmC2Fv7uJ/Br8KKNp3lI3fEi8zg06pZLpkdNuiV325u
fpIurZ//a1KcRzl2uZ0/L/BNgPJHcDXKgZJ+BbRCP+FiBEOaIRVuwptaPQrp
7KqUK0vBHAsi9Mx1YimabTcigPF94sMOPEqoPutXKA+flqzWgayF6QhS7EsB
niP2E7KBPGWWyeDYaaJjjmQOqBRP+7MsvwLK0Rdhp4DZgIGuSxeSysq6OY67
XdAR8Vgq+lA5p+tgIZe1V3BV04ivO9ycHmBRcj46ThPtW4Ejuaziyf8q9zH4
nzDcTc4q6qMmfz37u6hQTlhgsoer5rbgKbpwQS2QjBfY54LuahBvVAXCucMs
uyYNCO2//Sn6FGlPrpVfWR4z/fFfEL1J//lQ9/KJLvV7CSWIP3BIPt9uqOVN
r0sZSwsyuqdrgKr84jY/LyxYtvCXW85IGNxfYiAyoprIXOUdDNqVTBZMKFTl
hEJ42fmSwK/gpw0vX7OMyAg+0JS94lI8kS5Sj6KRpwqcLxiwOTjpDOv5RUWW
GLSoHx90D/HhO+evPOIaOTEscx/AKBELj81x19XgBDEebDiehyCrBowi4qvB
h2MZQ4pldG18s7bFO2upbX+jBlQVall342GMdWQyZ6lDZRL3x/UIV0XjWqSq
h2NB1FlxYQP6ZS0ANP5KhIOwEkRQ7AJLTwDMZ7Ru+qVaVuPrqy3PceayBOsl
6b0ekfb/lsKJCyWsGpAGgLtxqM6vhgrSgXFCcrZMBR7PTqOrZqvB4ekCmNWH
zR+qIvYrMupO+rkWVC7U09Ek+Ho6hR7En1reXiwIN0wgx/NWKd1cFdMyXksI
RqLf/7dZkyAgKXPYupECKKS3t8ausY9mF301CqnmA5lf/5DoS2w8Iv4TQuSg
r6Z0RHQxbrSiAPs2MrpC1siQcjcrCuT6uGMmi6EHw/eZRFqVNel3osNWqe6Y
ODBWgqEi85QQm0vHoxlkiTRSqfiuvmS9+ym5U+Vm343QNmXh5lEew3S7vMJz
Y1BfUy1eXQBQGbNUAwjqgeo43y4wwXTZYi5/4QksoAZGYlh8AAVZl/BEFY8M
DhMr5odGep1BVDc7NAQVP85eehs2dZ1RtHSW9Fx5QD43vloDytgArLL3jMSh
pLJlRQsWKUV5dPvE6RO2+Qx8+7eahxigNO/Mxjpmeqh3GtmwJI54etehaqgf
BXP8J4sVkrFP9MO5NwgSo4n4CYWuTaYUpkZ/oMsVQUq0ljclJBaRgeCbV7jF
2xqH75XGnlLjRYlAZiVNLOztUPxiZGb+GF9noNEfqCk9oyZyaG3AdeuAtOVb
cQqbwIrZC5BRg/VSVxZEx1KN4myzW1dEdyUHBMLSDGyLhOTViDwpCs4sa4Po
4t2ofgOBZESj/tYlqaywPyoGIF/xKl3/VK/mErfn+faCR5u3xe5s3Gylw8Q3
St3Y5ADgjRMM3kHQLE8ii1uL0LfI2S+quPKEtNt3Wy1Ny/m6QK6iMkYxHKVr
dj7uLVst5MqwdBvCsBdM9xWMM1bTtAg2x88HuKMW2NYNXVt+0LPYxEZTWmsH
XIz0+iw6gGaqVMf0m5RIdPkQehz4oYeq4Gd8vzXWxEjQ5bpbD0VUrR84DpMO
D4jB0TykKy/CbzeTERft98r9RlZh7gSAl0f+qqVuA6b90eYII3smaUKBEk1H
MuowLDHxDKsp3TKTIJEwlQEUVq8ouk+BtpAyBy3pRFVM4nm8p2Bx/c5wQ+cA
tj9wMNHbBzcy3b4g2WZs/8K1N90SEIejdTTZWqKhnFVT8I3F/UOB4yp2RIhb
P7Cy0SgAQMwBR6NrHrc8s3pUAsznA8vrCPyGqcMBX0bArc/voD+s6maC8OYe
1qY5des0R6v12Er0mJr35Kbg/Cwokd5uATD2zsLkfe6sht+LKBehqnLj9sfp
QzDpPblhP6FssipZCACpjSZA9ZsSoh/YdagnbyyFik2oSxdHqy1cBSRHU8JX
H/+nOCsXXgD35hKA8Pl8pfAvBh5CUL1gUdretDUaJ3Cm08+55ubymP/TDhJV
HCOuSZpTyGU3PVbgHECx5pd6YJ4vglh3eZO6f0vWD2loLToBHLnaIep739de
JoNiYeBTv0+i3wWA/DnjmDwcTU5LcaNcsOWRkBDcv8DuPMESs9AR+kecpXz0
L6JSh3iImH6EXT5RQCjWeOtjc+AI/J9rNmW3zHT/5cOy7QjryiMP7LdQoBHh
XmSYbWlhOEnajrtWbJXcky5nQhp1WnJQNxyEYQ6X38CzuypZtLSxwrBQ89Jb
GcX4olvaVP+nYcETphTsOx5avwh6c5w4AT3MOVvi+k47EBNSg27Pqdm2erqt
NcYopyK+cRJDfzJZtVEBdn+qz59qAf7Tm6AtCb4UYgxNCRJzOGPQkARjeLCY
zSxV6wEjPRnJ7/jw9xbEHdSAw22h1V2+lc8lzoDmuF4eZJIbsRkjZd46hUY3
ZMX7rhGW8uOEZwauGRjwEE3gbF9fr048eNFIVbv6vusnVk81hCSv3vQ7Ladi
DNLSaaeAUJTie0wJR2SKuESEJxO2LO31G2UDh+tZ5EVTs9Y1JfpnIaFLAbJ6
KWLibuCUHztnSrCQxOH5zCHzNynYNyhI3wmwbRwzg4hDrZ00S6CvaVlCgeQx
MZtqwTZs80M3clY5A1MX28RTKdUTBUGVGFqEhPOAeqOhJ6xDZx0q48GY+Yb5
44sYEeLggbCpkqJ0tzlSZEN5JX8Kf60s+FsYEEMt/XdwB/fWzbac+OM+3Ir2
czZXm7FJaHKVo794kljW4KCmf6M7FdrtJ5nwBg1PE2fcnOfpAvU2tirgJWnL
prcre3bhNlfUj1JeWxXbSKRK8pU4zlf+aYkPcG2AIP3FrjnVTJGT1nHkbtN/
9R96nzWelPbVds7ugMp6WF4elcFXg5ABE1HFLH2hA6Y9XhKMxxv2Cmt9HdpC
mAPtuPLHiFhTCSFg9ZctwlCIM9T7FHqKCKSUQ4+kYPgDYj5iHhC/I/K+IkPh
RpNedH15ASM3iwp/jr+1iFDCrCI1ZChkffHkfbNpwpO4GfC6kUEdk6HyWQnD
p2M64QsyQUl+gVtktSbfhgrit6pl2tgJefFvW72XtXTcWNtwjAEHQSXth75/
YUjxlNUg0jEtPtzU6jQZd+RCEXVg9HdJSv3gmDhV9U4X4tXf3Jl5OXf4Q0Lr
bLc+EfkHZM/pc943LJyCtJ62UrEJ33dt8CG1DQ9gkpvac1OBczBe/uoua1Bv
0uSK1qtq+Ri7yvENPg57dQ5/pm/KtmRB1I4VAPwehORL+RDln+KTu0cr9Tu8
yVDB8nPEHT8s9Cif/S+1sshoB8D2ALP9XNyJmlBfic/wU7xQLtuZxLAs80hK
4RaEc19pgX9fsMTpOLg91Nv2HcA28gMMBblNt0LSwSETtqApqEooiyzk1k4O
OYfqdxaD2NQs3cJ2fk9pX8ETDf/PXa985dOGi+XqMgmnmrmsqWjLqxEl/cSS
UuF1XsILCAwWIkV0DINyT9qGoJLiDJEEEhfS8H0/WwjprDbfDJ7sGPDFSNIO
TR6lMziKNhhXhZPxnw3UYHcLSKaRQOOXmEyMRmQZK8grKrkta9e06tR6c4Z1
kcZ3gzYMSglNtKzYKOsdbdga7PKskzeqNBwP/G7iTXd18bYiYUbF2TlBq91f
/gNtNR8c6X3QdLgPZg93EdqY8TBVaqvb3TDcb+Sx//BALMsH5ZB+bkQB0jb9
4X95HqwkpK/SHDaAi4FzG0h9FAJJ2kAjxq//gbY1zUEsTGEu6iTCoWlFHjXg
OIyf7KgvC8YZoRJhlwOb0UQ/MzqyTKFHmc0OEk0UCdLbZazeOa7abp3i1mB7
SVmnq01VRESQvGXcf9FzWwoKzeJ69J+29SJ0KxGaspWtY0RxE7mjtTCvcwXm
TfBvfWEjzNA+MomaEcw7VMFP8y4DLmlR4xteirAlxHDzMBZq9sI9su+qLS5z
j4PYo/O+0A/h2mNtDAm/MWuFWMMcA+zI+WDTUAytON6uGUa+hmghZVXLOxpO
Bo6bRmciyE1EYei8H3E6tmyfpZtEmNHClm4MUz0EGstQ+O7kVqHiBUy2tzY6
rh4hwteq/8iRRN4QEdWjTFAbHUiRGhCWjAewnWnPm6AiMHjfjrninQzva/8V
zf1hF7BSJ52BCi6n7/FNmF62walKYsgXbRyV0sNOMrWQNC0+7FllqiRwnEw2
7nnEbixTKm1CPFAzFeAghZzxxtugBdj8eYQjDwMpkf4F4hJVJBOZRg8HKHjv
9/DNpdJGvvuvYDtqLscp9ZmcIHUSl2Noe/PZJ9+G9AMl+nmWERwFm0zEuIE5
aE0zS1wEiWkmTaqBYRPYDVVJ+EbK2z0U1XxhX9N5ttAFyUyl8sL3G0FGbxSp
Q4gJwJoruRfgz1q2HVi7o7rKZT+QFoh/4dwhiPwlBwXtqgJbcxrepETlA2Pg
1rToWfDyuH17EJsPuSP1qtudvxGvgwKxJnjOnj3dmKpV1wM9kn4PBlqLhI0x
lNDZbpVf2XZ8KPIUnQNPw5YH0+CxC+c5yskGOSS9JFlSOfj/Pmp8ChrKxUZn
SEPm0qnzkSGXlni1Ij4wIWK0NDHhhnhhMvyiuQS+2922EKaLrFSPV0OIY1ZS
1FdmO5WeIZX6TI2SqUKTn8w6Nzh09bjnSxqrHfSAZWWcfgacUeDs3+CSyGnk
h7pqO2uHoYY8bn8ZrD+WiFDkvy1HoUKS42w7M0m6Xj7UJPeqtjnFT2Vl2gAO
pSAlH5nIcqEse8M12q4alAeyWWzN9boGbSODLpFFgMVsZZdJpbhidi61owK/
5zsX4T6RigDv2nFugFxnzns1+y3cLuSUAH6JXGPR+f9XcJefJ6EzpE3yXzvq
8zrvnBRpzVEkmSZyTPlg7syenMXmMX77IuhmN4uTTNTUXv04RsxOIcD1v9JP
FuLchL9ag0RjNUE+pkJNEdL176yR5y1Qp+LKQsoVoCi0W037PP20FzAj9Vv8
EskL4VRt/sjcztR+kvF6iEGZX6/5JLjZUZyIr1FW5d86I4nLYTNI+RAABdwY
04v8fLKLyCCGGd4PQiL/bV3v85wqdDjYhBo0JEijBCupabAbDZDe9Xx2BgIh
VD1zKhom0qkNyEdlpvmULQEsdCoYqAH4j4Pms/i4PQNozMdzdZHcYKYtAZ0M
nsA1IqAtOk0OIwHOSfrkN4HnO6009TbJryxZt2xbwWAWHHJYOR3CwhdqAAIq
4aPufRvkxp7T+6KjU6F+nbd2g2St8GGweMJixw/vB4bKej/e6TEGhirTe+vs
ObM7kZYKNQswPipHbAlTifS0sDitukfhy8INxmnEEcxPspBMk7lgpz2LGcCP
9XXLZATtPJDAmbS71vnMGiF8kXWlp7zRb12S2Zam9V4+H92qsbzxHpDUhifv
cJvodqLFykupTKkTVHpb1yn8mM1pSSwLEzdRaSnq4EQP8NsMLhS5GTd+THCy
qDkckemQJAPgrSSviphNe9GazsAysR8oKMtxV0m0aEz0YYQbgeW5OBt+OJFD
nTxWyNKRntzSkWkeemeZuzISIlGAeGBwVitII3IqeLdjdpWfYCj+xb+hb7JC
TDw6x4LdHu3KkzaipNOVrggLWYpeo0PmqpC7yHtMamnq87Gx+fSXsXy23mAH
k1O8Go3jPD1OK+Mq9NNkeClfZoepxFblYCH3oKt+Qk4z39oRidY0Oss+3KXB
n4hocI//9L/gJ4wPy0Bcgtuq2ZfIQwhNuGkeFI8qIZGQKwstf9Kg7mJuxwy5
RpQTzj+v2CUs/hq/WJv862G7ttMxyWrig8Rwx3/kg/yuDUVGfRu52KH19cZJ
ZmPTY7D3uHetrI9c36w7W413TxG6ElzB7Pm4U8/NTTRZnsCMnzZZmkmWM+iJ
ImC0NMWSSNZObCYvV3UZ1QCwBD2/PkoubtmnSAFEL6FshE5hyHj88R6UVb5j
qPzrI9SiKUs69PFMHiXHdU61/RyKDDrU3UgH8XqnQDmCj7fuhx9vCxYEaNsd
xSiUHS59wPyTF+ptoXRpnJoN+fKZJ/y8Xg4Anf89BgcFbha4Gskc7c/Ww/BT
/GD1597V5dhCdx7mah8fMNZYysZ5mLTsdgvzQYuBOv13m7S63g9t070Npxho
SViqCkA9XJUE8NbReXrlyBEBqFSjfkKThjMQLNG7WDfdX7+SYBCa7rY4ynID
auFUMaOIWea3Gxn7687mt9Jf/vjpTvSqHAZ6cizMhyii8sFYYAy6gQFFCNF6
SeND+YGkW+5Z64GvAIaSwvJM1uYpFA2xZlt5Q08UG/yAbDWO2EZDVRmAzqUC
UpQaQR8cMC2BDk52zD9reVWpeBAzHSdI1x+9jHTZ4GdRtCyoAU/4ixGvTqEJ
yWsmf6xw3ji32ZjRjwGeWA5Z3qj3XtL3mVLdU/JTxmCd/I4+8cAhd/CPihTI
AtJnj8IBljihiBPlnpfkLtNbhDP8lGZk2cE8YA/rLdKTM3z4ETvyJVdx1fUy
pFTvxVZD2Vda8bQBx4CttBcG0LGQI4l7gKzhRq8Oh6bfrVnhFG9zbzl4PhN+
hYhXFH4SQimz4Y8go8K0cudVAPcTYkM3HpF0GbIAx5ubDrNvY6Tp9OOD5bF7
npdWAwRPTEDh9gpNrqhWUKDhYwiKLjhDZKhnK9B8dOOcoNEjV/cLx+7bKh2z
qoZtWbn7NBRUf5nrhB7/Sdbo41JmtvF/IllHvk9ZQlKa+iUhar2Omi5igB0g
HpP7rdpuT9QZ3Bho8M0gjb6jAM9q9ldkAF4kiaJfdmZhsZ5f7pNfC/fOMsxm
HhTtpBnPCFC3oFCq+p+fRBdwjKhgiUmWiXAMnJ6YT0jptLlAT8g8aY/4ZKAw
zkcwWkduECkdE4yPFjkrAn0/JTwX+WjBQVokVjnZh3Jhb/d2axC5gt01nbCf
4CTMdML6yEuz24mznyoWMuSDH1QNUdys7bwMdiexoRwEkmF7Qby2dubALI0t
gW74ifnGCbyWbZAQX2N7iQIAnxecDzuAfer2wFWhCMgHOeT37sR2ITHST35x
ah+GfmQNijyJurMI2t9LuZF4VTULuI3jcDe6uRjREWMUK4w66j4MirAvubu2
obZclRkDDE9lDUEKJ4Ym59Ph4YTwTDMMpGSxStiBWvqAljQV8SCSHlB3TeMU
LDIAplL7TM3jHhOkSYN6G54mMX0AEf+ND16s1r8uRScn9vfFgQtEDoM+ER//
1cljehdJZnPoQMYk7uHs/oMOBZ5Mv+x61y1fvajq0MRedHZ3ynW3q13UaaZh
C0gUSFP5yKiuRpJsPYsAv62oN47sL1lr3TBj9B5OlyXVCTN47C2c6cg34129
J7GPGg7Ya74ZtBQizF4dpl6OiKWWVFhGSUcD9ACWGIx1RMNDLj/kEBZBs085
3QFThsYh2u4DZhvBSRjQAxwSQ63CHrl8wksVL0ECnGGfJ17zOmJmxdbLrRLV
ts+DAzE7CcBzj/RniFy8Gr/cYK3jnQECWi+adWfjiUgbwKCZu5cXwdN696jw
fxgqNlrZLSWsPkOWfasICfZmnEzy1fGpvEjIvX8HV7laSI/cuR4k7uEe1Bcv
vZJmbRFdktyeLWBmbu6CBuwDxqqEAiDMM48iYWQTh+oXFYXASU1aq8LugIVO
2PY6rBw30CHkeDkGHR+cjoTaM8l+kAqeB+cMYMQbEKAVGN7+n1FSOLczzw5d
jdeaI3qYeDmQ7twgUeSJwZF42JQLC3N/JPHjnJIQeXu4COT723jQxnqC0U0H
1bozpXIfnSunEUlQRIEd+t9bIDX1QMD+6N7AND/Uu8B6n7oi7WQPCIcjCcRA
XCkDRrj68v/XeyjgBHsw7paLX1eqQSXQYlnXL7aCnZzeVwcZOzkxs7N6o9Go
02RgAPqw+UImcQx3cPIA5w4BsrB1E3V//mM+UorA5+2uP9KNq4cxvfHnB//8
sEq/9o+e7j2Mdyn65/QDbT9yIT+TotVwYLcGh2vaS98tSg/51JKVzLWzEDf+
CHc/OACBcjBVcPXggQSse5svlGNUUG5cP16MkqxdWi09ARwM2ClWgvhv62h9
jS5L6T4WSRJhmjSFbesvS07QG1qsZtmguNHBBSuUiZx+HXFP2jn6CfhqIy+t
6dSVJ7FFQ65VQv4ahc8488ShfuBU+I5ExE2YB+Riqm09L9eLSBXvBWhR8q3u
eZuVmC3zA3SN0/s88lKJAY78YNl0K5aN2IX3Hb55ySbx1BjmH3P9R3MYEp/6
X+PZv06g9p4eAh8a7gnRxWbCRrL4qPO6Y7fbzvzrx5b47MR2kgzk9HfZQprS
IfJ3dDuhbV1pigs5EyBPXjmysCZHd2sPXWYfzXacxLzwzwNebBEP6PS5qJco
EC8k/OKF/nVuCrQ95kKUEomqfPD/ZSGiDgkBXB01mlL6iSURKQQdML5t4Ymx
S2WUcrqtgPlmWphtFzM+5bfCTHrvoronvX7Wbblq1D6cxAA3cdF/TSMUzGz1
1TvcTJaLLYrLo53K/2zFZxcoZE7SCjTV27j7lxyVxVJ+366f2x7kWEwUt4YZ
YEM7acbZHRO054vpHR/R8i5MD3kq8MZEjlKMETcqnyRVR5GfyHYHnwZe/RmE
1hkUkzAbEd7zmPVXoSqR3LhZPrTzWRIc0Ri0bzJwsE0r5zZfD6kN7xK+GucY
y8+oZZ+wRyDtF3LliqdjzDmnKPxBYgldvd1PNOnxbGCTqPxdf9jHxI4neKSD
9JJSadryYYoC7GKbiIpMU84CnRHdJBQmadFhK04zFOHUDs4GvdGQddcnQ4VB
Ttx5fGCHku5px6F9VaQ2F/hL+ogGxbkP4JoOLeSIqQdn3u2FPlokQ5Dn/kgR
GwKM1nGzd8Syd1NBmwrGf46htXrabVUOm/hr0b2/9Tz2CT6ek5VJ1N22Tez8
r7Ck0CjYcCKpr9INxqKfblraZi1PYTeBc+aK9kCT/1fpyaGVOlgp2zVffVos
7VMModkBE5adfNVHi+JSn34v3x3/lzfQd5W182dA2wdeqPlkQncK7CzSJOpf
CSk9Sd64Tk8mifdZwXIbBWoErCyeX0xCoCXspx0ewNyuEB1uS1f7+oGyYTEn
4BcYRKa5A6BBxo0aAS8OdN6nb968NrxMx9u27ThPeGX757KBSaQoFVxNATB0
91N7wNClpuRP7v/IRtgp84F/bNWL17pjAiI1qyGf3bo4mPjogB16IORezcAW
TUId1eKPxipM1rDqPg3q8nILrKquTM3dbuRQTpUrx2GG6tcibBOB1aAk0RdZ
uBI0sy9hCVp/SSPT5TkEwbjbKNzbjj/IesUqGjPLQcZ8T79RinIV4gq/n6VB
k7MFs/0jixC1d6HwYMR9eWWQkmXXPJejqfJEEZ4t6ws+KNm9DbR6ocdFJozN
rQHpKVEHeUARa2KoMbXlOCPJe13G2Ylgq4ocardTcrFKZNFFurKAzitVj+Ct
wQLIgJR7mtrd/OW0p61fDn+n/4qCRmfNbjNaQMALreo4V38s2GKgcM/Irtg4
jtlqgGgGCli+QlgUhM7x3aTyJAOU6VAUgrDy9LeTYQBlsg0KozBOkf1ShWkG
rcWM8ZDIJaycTi26GIq3wvlBWUTXoNi4zLFwbqO1bApyWAnI51kAf6gilqQZ
VElEvjkFi/XBXU8FfmtfsqOLFTYiZcJqlog5b/7zuyxWYAyxYs1kRQXZk/hd
R6jwfJ/b1i7aD5cjmlkbpqZ4OsktpwdWs9MPyXNneZtnpyDL7nQrozykukp9
ATfXY4uamFIbBYo5Ni26vO2Lkl1uQ5aIX5HDRvysHRp/OiPuECqYB/RLvuBY
nJOGvOywQXH9BHgJBvnl4IIF5wgxKMbWNkx17IrbwcBraxsO+XSH9jkYiWkP
OCUGc4I0LyMVnow8EwtIGXksf4I02ZwQnUEqIj9OIojQV3vCEqPrhSSyDa0w
t+Jh3Y7pGsnxdEcTc46syvM6eUGkaBHQiRtOtwoGfBxHLWHFxxEaNsmDj6/7
sIvhUnP6c63k1tw49fpCTKgQ7WgopCm2R9LRtHx5tBvnCAaQctYT/Ogzltq5
xqCua204HRRz0e/l5dO6nfLGpQ5Ga5CouNeBojUXI/JAu6ngT9g2vRXMlkX9
8zvL31BggAqHLkBkuExKW0aZoMn3WT2J7iLuc3qSIq4sW8mSeRXXhf3pyZ41
xHpZAV8IJorIdiH1wG1rvZaX+zSCiJsKAaqT+nCe0f1hfgG5Q2rjSuIEqyEf
NlsiJkimgMQ1nyNMCbp84PDWUVyTyJEgPsqDm8mJVQmRTzExm0P0UbkOfhOE
ilBKxn9TRBJL3RBRAShXwd4dqTMiEEqB9L0/9O9Vtz/Hv1BxEJsKrev1UR2T
oqzoSzAV0NzjLmjInIE7r1MySTbyGGh26s/TlvbyQVaW1V3B5EDNkqXNo24i
6hbSMhWhFA8sLHJrMY50JVfdL/R6sWy8xHzaebufmva9bjqQbEIBJ94ZGWOH
rXkxhWsSk2izmyV4HLVDqm+h4EZaTpyQyEEdskr/wQaGwVPoR3QHCuOSGqVt
/Sd6e/Hfc/nnbJhH0/wU7B+vnVm5LqC3jSbxBzIpUziX+r97jNAClyoMAjw7
KV0uidAj1I6BBQXqI7dOqVSNh8wUbFMq75G8/zSi3Dnv2THn0jgLuuRPwvrJ
BDTmSrZxISf6qp2I8ySOEqh94Mw3EwkqW51pRAV2xmlRmmefsqzAuNSyPVwN
v2QP6BBwbkEalpaZrxXv3hdeuHp1RzR0iIDBY6GuA3MhZkpQh6r49Rw2xEav
kFDofU2v78/DpIzrpOZxJ6Nk5583fuq8OzhJVmOYFqpJ3B3IKL/qvRPO4zDQ
fLTdKl1OzI241xVJ53Gv7X0oXQjk8JqJH+5EEbE9+Ufsr/oLZgoffc1UsIs8
UOBFHdigLVHUtY2CiNQI3GdoqZ3R4Y1QTIYvEiHgXtrxPOTXgHNyKy9Jsw0c
4SlUdUfPgzZ7t3l35A/+IHxpfVXyTyWthe2B1s9JfhieLEZ28XVEHjcJ7QwG
Ccv+SZdXogwxY3Z0qZjFZSbbU/QNJ5OAItOkGVMRSOGKzdJZ5/xKNM6CpeC2
gg/KpYh8Vib9W4phHcBto+lcZXqKVabpzqux7qeHRqleK2bhDkCuibIC8ZiY
UoxG2uTmDgzvhT84RsYNVLO8jKe8bVFb3MwNp5cxTdNW9VQViUsqBzQzNKOr
ECRk0Xbr00Zt9hjHHU6qfmUBFPAu411iH5oeDYFjTOsg+GBULVFQ3CZgmEY8
fBroCgktnMfKcRHfGfzLp26OQNcTJGx+pZgK/kvczQCJnUhgA4mF5nGKh0To
OemwlCfF/46Hftjkc9WnHJhdBrO97vpBt8+seFnT24U+hQ/P3TQZfAzn1p/o
WArI32oxV8x5vzgW0PVnB6Sfy/xjTtOATkF6XjFJ1qeeaxnSQSWHkL32wvMl
+0ibQnZYyHUfXgnPQqqbrOSIMG/xvaD8f5JQ19JPm+QtC0/gt5krhYC4ndEY
Ry4eQoifP4ilgwym+1YKkR2mzIUpOEN3ZiuTcgc+EytpqMD9gd/hHstBr/9D
zdTTWocQcOFDKrlvxRWEMlAtidT9pF+PPPUg/QmB9GUayWJl9EQy+ZIE0vBM
TKUb/VBiIYDsFY6Wv5Thr4Uq/EahszOdfs2to06PgSc+bVd95/Psr9ZSicYK
GuZjc7iczmeoCD+QbXqU3KfWWeS6Z1ab88nm/94c4JAzlrIrsNvrC5EbV5qp
+vqav1bT4KQTz8ivcheYd7DYzG5AKQ7sqKe5jI6udGa+5Pv73fwbfiDDUS34
YDJ6SFy8qCqVOqvhx0OnC6kVUNyM6gS0y3w3K2/keYqIM/oFFucZxux4f/r5
clFBCJ4fk5BTMZWK3FGy20Fpt5R2LIXZBzO5Yn0JxSWqGVEvkiiLxYz3KuHK
xm8tTFt0+gTTw8FkUmDujKlKbGTvv4FUqX1/XFbSgRhYgGayXkkqDULQfmt7
bvGxD3c2DQ3h8sO76y50ChtAgNGgPBOGwKD/0W8G6dX1R/Hgl0hM8h2EU+Y4
EW0+Cc+vZ9ps3s4eWKQivIlsL6yscplvrTTQBu4L5fdTQCLfY+bydt3+BUY2
p5mxcYQGEKyCl7p0RfeOTlVnmxYlolls6TlY6PboNP3I1yjIo0Wu6pwomw+D
m9ICG5Pakyn2LjJzlpVD4hX36Q8svs1jFCGmWcI+NqP2TVjegf+0Oynk9aKA
IHxPgkB97Yh+G8eXGY5+m/PM1bHpuhZnvIff+Ojcjz+bCEwv+s9x5X1wKbo3
uibiae8N/dd2mda8cm59buKj3aOEcoCEGiIGhmxMyMkP6XDbmo0a56l2G3d6
2ltkIdWXWS+jwVoWvMUUz26OpTVPVTIcp7IRnRflUoSo+cPD1SyzDzwqeUDm
6tOCDL/CuBIfXDcOTwU2RWaJCfVt2hNae5U9DPPsOZFnKL5ft0ahHQ60f0z1
iYqiZ0LZ+FAOtDeVKbyLYxHnqsknm19fyBiip5sTCdIKLJZvy9I838Bb1nar
cTlCFAkHl8l8On0jq+CAdVOqjpI1j9HSTPNZ8kltEnQ6FdhpSrwcwEkq1eha
mAXAgVkDPMhj7tS70DYS9r2uBtVdvImT4EGm/WgsseOmpUc8F25e7TCKRn11
i9t2bFrm43RvOmoJvrWFErFcm9usruzFi2HCCAsyZwUoDXsM/LGR/GnKFGQz
mRnuvTwLUrNk5Jf7Ci0Pei1hboQxRp2a4nyZJjDwudmjQS4xqKqjegO3I7xk
or64QCT8a33gxFtKGaRhZc6mkr6b1KKoxgwBOkVvJa0UpQPa4VX0HA++5P0c
yz11IYyqV9XpXpvQ605k7p/CbEkYK+p01OTTklrGfuOn1fDKrbd4mJnW+jU7
IqoU1OwLG3nCWQh2RPE9+LUQnbw1+Q4FZreJVVM3YdgYL45I/4J1xWyHdKfV
IK+N1enjUsXMhWa+y1wcWcWnEVM6hsLbq2u/+rKkHZokvDyzDDoGSVuAW2W+
G48PFTiQuicIH56WXT5nnDfe9gMHLKFj/l1zkyQF+mUMXMRlUR6lL5t+zSxa
v2qTBexxASinKvGKIfA6nBfAF+JbLq8XFc+Ilh4W3noOnnArkAhNaK3Utb11
Yt2wsOvkcIYgbVy6LeFBiX/porNUcjDG5cB5Jp2+Hs7egqq+gbhZllqy0O1x
e0wVettXKAjajUGzqr+HwwiDXiLL/u6Uc1yIGF6C59TWmeaBRpegUj64qK44
7EHY+S51qOHrIWGh3HQEn93kE4vxH5MtazcN/raZrN0oD8qaAWtyi0vdfd+w
IrHrW7lL33Tykvh5BWyE40gM6k0pmGOLibqnrkjeJ86twVMjX8GFISdTw2IL
/BEwQZa4J1LNwQy7znHJK0XLoBz/doIVolUOlnC7fU01bXPPZuWlMmQDkHi0
wm4ZkPYL2+jpFisssx0E+l9aSh+Lu0pVZnVdHr5SIffSTtT8dFXn163SsAmR
JblHoSdZuL/M0sijvJQZChMmPKKPelIvVB+jG3SzOVcwuv0n+PGdANtMCUcG
CnGjj9r0uoMoWcZfzOUOr9TsEvgWr1IK2felVe3g91x6OON/Y4kbi2bq6tKh
QVJQoifO3o8t5pJf4qWoCkgGPfJjVdiT+xbeqVlcVGQizR8tjwSwoYIlYFAw
GEtgLCXXr2bD7di8S/LjJnRGc3qpjxxeDu79VTKDOCHpAikn3buUfI0Njrx3
nI+7hPCFWQiL7994xykjMPOtSZ3RmZ+xsb3KSEs29d6sMFUpZXhani6e0Knp
KkKjATX66PKd9vVqXyAvu3zARP+pGvIkxsy/v5K0HcmOx9WxFEhxzgVxa1HB
9P/pBEnkkrrbTvU2n2jKECP92h6yakR7uHzAoKOj+KnyHnQ1BLkRT2a1j6Qi
NWkgY2LzV9ljv6fTP2FJDkR0rwshev0crTWnoNWY0SC8uCp4NajoJyn5V1Yb
314KBkAB8gHBPZC73nQOMtADToxAslUl8I0a+S5zFK5OKZ6/FjjOMs79EID5
58N46GNglS/ahiiP85a0W5hUwKt4A5jM0FnWKk2g32DuCH3Pxkf/u38c/W3o
k2ibTkHWfaOAndaVdi4m8lZsveP7h+XnJe9kdBxOwY7c05/l3miL/eZ+FDXX
KibWsPdgikQpCZpgoNGvRds7PdyVQ/Up7JVzt6tvWuDJvASzqFHNqWPTiZD7
bdSrrD6+cYqePfNFaL2JWVoe+MjP8qnwK8XmnfG6NBOwh/BL93trsmT9l29u
oPzVzTOKQGOWN/cEy00UhdwxzxIC9fFZY8mb9eqxzpAoyMFxmv3J7GU9dcqG
QbtnX0gT7JYMS46LSM/kA5aeoKSPTIRZodkLl8elBJjmFkupimQemz5igb3g
4aedtuCsWxmLzvtkoZOOQApg/7AUA7E6kfVEQjwJA9DkyL82bEW/XboGoS4V
oGlWKW43yI7Urciy891qo+OYjlaL5UcJ5fqm1H2s/xZDQUR1GFhwD3btvndL
rjHG4ZlsjL3OVRbWtYmOOEfaFaNH3V7e3vtq1zzmzSP6R+SHhFxyW6WgYECp
9TOmznO3wKMs7BSg6xZRz78RaqjnKaTsMpPI1QcdzVfmU1VegfhGwcxyXc/a
U2T7rcHQ6ZmO/YbjvDt5gldMNEgT3OURmxOggsszgbfh2s5xNraNntFju+mD
N1SNCJi9mJxSIqseqrVRqvLKL6gdU1g9vqQzPP9benWymeOaT6G3Sd15gV4e
QfELeKoskQfTIUKY2UFmoCWf+7aCSu2BkSfHtuU0NYGdXIXPlEkFIKDqa9ri
VyndV32gdrDQ+IGMp4pgnXQkmIvmz+031PeXdFdHEC0bvrEcW/DbzpejBC6N
6rqa8Fn6ENbAoOoim4VXBFnbRqgkI7GLFNbFeW1AO9q8xRnmADceDMe8qLmI
v4h9NrW95jdknPlC8aFU2bb387F4UaZSLehnDzQUZh3zW89gYOn/VRIl0sFC
WmDEVbnuSewggxs51zicfSktqSOULq2FjfluZBFglCk83Bht5zE6NgoFFVsy
IgSZvuQktT8Qo44BWeIRhW1fd4tGq9CFVS1AdX2AthiwM2g7FfIdvuTvcKu0
MXCEmOc6aBS+Gg8bQ726lizosPTltC9sZGALYrvtRb6lUviLI1dww4vNtqva
ND0x86oV6KzNFaDDUpjo2ixyf3TYmZlRX30XSXSdB0Iu+nSiqJvdbZSG23IO
2ghaNj9lK4FffGkQa0U/BBmKjBVLfhud4JNz3pbDpIjMQOdQAj7AEAjiQWNu
zyb7GopxVpmHGNK1j/2PaTkyr2x22BZ05P3dB5FPAWaKvfYCocqfrUsHmmCC
IUgsvIS4LELqHJyohR0KVvIih5LsJ0hJZ+BrCaAk7P4RyZqFjurQjPQ0s1NV
BTA6Z8/4dCgr8vXwp/jHN6KsyT/n8kSlb1gBpiMku4V/VeyJ1nDnMxQu+E0g
xXt2aRkBnzz8MDK+V8SB8TB6O9croirBomiGY+aaJM2CUrO9QsrnwSJT9KW3
2VvhNJZDXZ9b+0aNke+wdwH0M8JpVm074SKPw5mjz/2yNNcTGcl+T2piknjW
TpTDCXkSAARBvsxsDClURjHrspM7LFXETIWHn3MVumLVUgaOsKorsagTB2q6
08nAtisz6GZB6xJg87VAAyWlQf/C3K53nhoXVdpCADlpO9Q6eqM4wG4MYyJP
TENrs8y4lqL4rXo5gwWraJB3/0QZaMuafQT/PvzOp7RIVWGjBLMMi/9aeR3x
LKUBzkJF0aDhy/TUvOx/zxBQaNgMzlOFke8bzLNkYahoARdJsvWu4PI8pg9h
y2QkSOFhrd+PW577zPtfv+4lQuKW/OzlCfvt3rGTVG2GSZejcrWuaCFYXXbo
VDaq2VRpJVeYuRimeQBLOxkbZY7Ymv+gjspeW8mtQGMA8mkohkCLldGBumSb
Rji2x9LObra9Fjp8JoBgIqJZ6bNfCqxpJ4aNRn4Z6iSGfSoHPJSmiCl7PzUr
ssL9FtQSfZggI18cvrKPHocixOVrjTY6ReFaxPRWzJcwd0TN7CpMuwGHEj3g
c7xMTNdd7BnUDAvlZkn5WHxnA5tgYVNTjyflAUX6YDZls2XtUy7lMACkJX6k
JevUKU5VX0QR3yrkBWNajtyA8i3qbl626Q4mJTczyCrlo01tWCxefwjJxMXo
NywE2K1zHm+J3izygwU7X+Lr5CGrLUch0oqRcbTS5JaGTkf3Gj9bjgOlZOvR
lLiCq5vQQsZHn1GKyKi4GxDRuCNJlhDKecxNzH5jBjsRgWNtycHP5n+W080R
IDp+QoVxc1aJHn9TEu4V6XSAfFgA0Ty6V9ovI2wYjUyYHXUanJgQTfifmVwn
4LdzvKzBy0lDJmVT1IBy5HGBeQsYPdXafJ3j03j2bp763fkhvc7g23eNzH2z
5Lmnxs6I7c6lYqXeLzUUn6NKcHBuyT46NgL/bhJk6j+j4eP7wJ4dRlLi8oVQ
eeBExZLnJOFhCnPQ+qmbVYCN7QoIAS3m1zFzdVbwpVaXbdNrt/JvOyre6lVC
/ShnJKog+FRuwPqmtOQH/Pbb9gKVunPfokZDwpU6RhuuEZwifNBgOMI7BJuL
hmtvSpaynbzTiXksxOTc+6WxIz7izFnpPnw/cXFMhkH00Y/ZDoJc9r7WNONo
8nVT9ed0tNKZ/fkSfxiuMg4tp6DnLRoyFI7nxIGUJWHDVA0BpZW/QzpVk/9B
lkmp32CaIY2ZkgH2IXqXN1R+JcatYQLUwBho0Zidop0ShRhRx1GGU2fNizdO
4x6AZptxuWU/FwjHUG25FeC8JwW/9zTuXKVejMuvvNZKRnJsRMubm8PYMTmh
RQaZ+xMuusjJYoMcUhJgAWPilN9PsLmUyQCFNvw+9yerX14p3Rpf5QmGIjUa
Pwn7QmH4wM9tF1khv69QEZ4N3QoFt+6Rp2FqynmHFvvHy7BXAjfDz8wJNBU0
w/h6uefMBskmRc+Su7apjpT8lo1RQhrDRlD5Y1xNTVKML3YKXTtBJ2azaHAW
JS+gTgeqz0RX5TtmND3qPYKypkp1eEK7FH1g1HJrA2iIjf69fuycdqjHwUfP
IDzgKM1n50K778mhUK77rKGKLH0zv9icG5Mfx4oZEO+T4/cfTNh6q/6ULYFf
YmpQzr+81ciOusqYIkizetfRe0QM6rJyN+WP5d8ZbLljC4/hwFf4fh5I49uQ
9dsDAvUGRlRUAp+hqcYc3s43e1CW8DP+D3TwEO1vNxcFdcR0mK+QSmawNN/3
RROXzdnG8QZgzXue67MAWS4RZDtI5f7FNziUaaYm7rQtbbG0FkXEMwzNKi2G
OPsi5P8qDH2x8NXIpMPms90wEqZKUv6ByAxKzLGou5uvXzqg5UIdgDrU2uwi
Iq/wEzBFjIl6mRxFOZ0xXCfeBAZWtPWNbjGaN7XYB14OSF76I2VhQWMzUuye
PO0zvR7QKeGFYqz0kiwIjJaytggcxFy1F4UjjE4/qA8rGKue10I8uD/x8KnV
uVSM8odhEgksa98de1UnZbrnvCl28k6Lf/0G5i1myhIYNAoaM9Kj0jHjyZb5
+M4lei27T6/FOW4lXGpKh+jjwd60/CE0XtGAqOmlc6nR5DtFSAYcNO/RG7hm
2rxGCmf8uvYmFP6n5BXjEaeNz12DtnX7TxXWIxUDwJvqWLZ0Jc/hwejLGUhP
eT+4mug5vA941GgG0X/fA1MDnyMGFyQuAhlx29zk+guIEAgKrISegjfsyhaK
JQc2aB/Q+iFN1mojpPigh8q9vn7hLKXnpbQXr9IkDuoR3x/EGJAxT1QhGP0f
a5FLoJUpkdwzxfGyHRWQsmdNgLHUf7ExJqfOLWe51tFl8p3DZDQxCvAamjmp
jatuYyDmZPUSGntPrSU0BHbiXOA8QcAIQYRaY36ZbwwBlHBGEVWOz+Z52BWo
OzHaqpkkqL5RFIDCBHPjPUwXqVWbSTl+e9oLqli4OOVbkYARfxUrTZpLPEbb
spriuLDXd/2CWtA9/nMYZrVsj0fMDwAlsui87WQk39LwRwc0homnR2uHUf0S
pEfr1QPa4eFOK3C2Jbk5hRjKvEGQjbh2KcK00w6Tre03w3XCNHqNmlLOWyyU
qEIyDO4WjU3/gfYW8z5xaOC6pJAn1fjBt680skws7cfZ3pcyG3B22Fw/Klk6
6kHFcDoNoIC6Z0DtKvdI5ZamVAFlTtprPpkG+nSyGBjqX53R8ZUHiDEgPxYo
Pz8c6fkVim0TzY2FH8zyWYObt91b+YdvKLVPmnimSBFk9kmyy9P0Tsz+2DFQ
V+A8iErga4oKQPVdNaZYistgEGwLxmYXwtnBQ+45Yr+mlVtXUMSuFsJNakjd
4pWmtMneyiGdTnx61PLWOvODIaC4olI4/dUvNGp/+PwvEqXr25UmmJ6cybMb
YkdQFhTg1RvQYKG5wbRm94aQH6jhSRICTE+cvJW0+XEcoWAFO8+E0JTEoxhI
eyu4OGNmD/43iEF64dxvnMIvfOOlMcwnGNJi67TGiUwVnZdsNINUhQbK9B6E
1CnJOBpSYayznVLPQWw3e5KiEuGvYRf6TPf2muNUZEIiJzwuYzt9NJB52Tv1
Ut4EWNrlCIoNONusSglETnW7zPteXW1kYwm4PCO/OwzzYjOFXiWsG8mU5tw6
+nl7dlq+2kCRj01n6r+c5fAwdAR5q3K34/rvQE+0sJk7sJPgkimi9EON9RFC
t38rDldbYehHXH03jaY0piMCqWvukX3ZZEf/JsxOuCSAlOY7sSdNB5zvGmKR
zuBY2VDwguLkHHviYWTy9HaeG+oKGMVdMjXYCybb9OkJvVB6LYTLUThqrjl5
Zv8pUJZLUC2G1cg/fAoDwdISJH2MwR35yR/mYdZdyQgFPxgweJngs/GlmlJV
qqf8WYYttogiieKF4AbO0i1G5byyLBqgC34sZLP1ZN5pHsFpfRKdHTNUZa5A
teSO67bTWYIzPlqvzkZd/oPn3eLAzNt0d3CFE74Syc7tyS9eGPYEAqU9lS62
9LQ5azA2ZSJqZ1OBgGUMmqwAxrAP+EDbg+ut0Vr3lvuIM+rqZPTIurZcz/Nt
qMDWLk5fFYXNa8p8R5UOfEKxjzPZz5076w/Bb0M0lV/30AEIlgpYHLR7nFBE
bT7t2ysX4oaur3AGZ0rSacgvLuTjJ55UGBbpuTVqY3evV6kiwUbOetFauFNw
KZ3dRWUM/I5Fh0j1OG4j09RAMtdUwBhpC8wmQXl5K1OPri2Jzq/kIN1U0H0m
jTQ45MDjhVIIVnQCJDLF9Hkz/TKx2XiDd21PugwH22b3OO6yBowJZutr8TsE
UUMuwiz/SK42n0KqO6fyI4A5mdlmXAysHy2Ux2X1LfJUT+nxHlYd/PskP+BR
d5nqdOfmBGy6scIXbkcH/QSKbIb4IKGFt8JpEaETj3D7X0Iq8QTux+UzU56N
1yVrgkribdDpF1f8MnvabvPeIZYURtbiXOG2pNdMc9jP1kpD82H2LQcHPSzo
dPaU3+AqItf9m6muY58Pfc/xoIRxqGFKt6bEngHLnP3fdHmJ/LlHWx52yplg
xfwz2lfoJ8sn0YMw1JDF89yFXSUy+asQLZqN7REG8gVCebXcckBHqR0oRzXw
2wL4YxyCdUtVNtp2hrOOddie22ubzuOQvwRNu/ckoOK67+0tg5Fi5o+qg6DM
Ufxncu/CMhwo31ze0AKeTmUwgMLiHZwjDV0ThIe4PaTdbSFBX3gT0RXxRkA1
0dJMECI7wbyUjWk7EgEyum+qZQjRZUSXadm9Og0EgfKcDmUszQ8C3qOkoB31
/QnaSEpNmMSkh4G4qE84QtKwYj2csUK/zRTcHSgDMEwKALX5c7TmInqMOxHF
N9WsD8SSFkddKtBthfaKNeDqOxcPCySbLijmLMbqCdkWsjihhZru1FljsCEu
hWZ+MW1NJ6/n+BfHrfoKPPjUC4BBl4sehl4B3cFJBjMuC0qvxXcPtkyxjSD0
wTt9abWYVuueVUlTc8a+Manj84XFX43/RA0l+kO/SUiapxIpMmQBMgf583Sg
jJKFmLLdA9rUt7i6ruCEeoXTR7hgmUCDPhvSz5ztOvgv74CAU+ThpxvIPTIE
c6kghcTqPOK7POAV9ZcpIksOwidSVGu97ILFMp4zncyGxQ4FHjxNDzGW6NyN
P0Wz13EB8YaQTG/n0dsrqQ6dC/Gk2/H95DoNeqv5CfK6Xe9Qftw6515nXpB/
oHXnu318ev0rPU52jX+s9PEcKNsw6MSRCOygEIhApoibq+E9RnxFkkMwIz4s
ZOCmB0IuPPIYwLWHUjwrvfSn+cykTKsNeKQtf0XNno8s1+ysbChgfk6nZGR5
IyhReeYs+HU8zUDkZfCGwd7xb/Er3GApkjuvfE+1BhyGIPKzabMZnNDjklgC
cfqC6liriv6Q7hX5Eu7iVcMCmNNebiv3JlnBTZ/LWbab12ASpOX66cDYD9QX
cB0aKAv9WNiH0gW9qPm6H1n13cmZeKcmUKP2dCikD/Up+n/6wcvdVhiFZM4L
VTiFuqyFSPGqqO/86BRCW3zSeKhss6BuQBx77Zd0ETj/06Un2YmScL84rG6g
I3d3iQvHYLmwHI+J4jzlnv39b5IhGnZ3B7U+dNirIkU9w6mj9EzsNCi4Tx2O
zzpqNJ1J0CYY4rAOxl/zAeROmzaNNpD9IKydATBrzvVhDwRHfhQ6yN1CuhZ2
NBMqXHKFMg36BzJZSVmSn/9GtO2BSrXQdX2Mqt+AfhtV5MuGo6G+SaDw9gE4
N6PK+y/cmwTU0zur6FMg6r0tA7nmNyjWsW2HdlHnVEJMbZL3Zy24AlKz7E+E
ttJrWPhZBcRgeuA7TbynG4wE9U8uXD6SeO7SV2HIazYU8PwaJdKo4l7SPUMw
vJcOBxTmi/wgM8SWoOSIZu6vYrqfOQ4X5jenQXt1kVBWlB0nyTc3AjvgJ1nz
hyaC/v2b73TG5MjXCzyHREz9dRwnUKqj0eNtgF8s/Qpkgz3n6Pvlk0+ybqyp
BjKuKdi3dyjWw1PhBdsI+9z253YS02AKuLFkR1T8miTK7p+FQATgHnQDpQZA
53BStwcJTKPOp0hqt/aoV/AK0gQ3uB7WXS/vYwzVJCHOMdtV60gxY9diMByf
Ag2sOT8Dn4ls9En8GdSCqbSnbwsmoZBalaa4dTYBcINTIdsVICwTICLelOkm
3fmrAGevyfjURmfIqby9Xo2lviI0WcFaNjbAWCq6iIIJENuz0aLkYwBlb7iW
weyb1fk2zdDqKvFF/a90yMUy05+jcB3OFC8R9SgF6gkakYzs8BZK4vq/CKWL
jWL4MydjgcFGgZk8vvV3qR5UzbKZV8D5NQTNt910OazwQFivPkFbENojR7IB
52kELMrjCeMnUdOEfdFVUxipuTxFH/U/Y86DwurmnPMhsKgJgl5PMsanyo25
/btvrcD8CTNIFlMK+J+HZnsUBk+1MGK4W4Njo+ysnah/0xF3BFa5nPLGh1W1
3tL9e/J8jdFruJ7XBv1NvFEJpMbUxaatHm9F21j6W+ynktiqMNQb4//mjap7
+s44ZoIRSRoY/KCkaeLqYw25HA64T8hagf3ejPxhRtKiz0XAgZoGMGl+LqxO
vJRPMVGJSEGPDll68hDitE5/t6jhsDhdU4l9c+F/TvOFq1XnsjSlTm02uszJ
3ofn7x4Zjde6mZiGPTxtJGeQKlZ+0Q4oUKH8KKqur+9V+1DhdogOM9+En5m7
4DN0uTB+Ebg1M8/xdnK/7NaAv+HmlFSeDrRiB06zgVVj7yCpkH+vYEyKnw+I
TtafqJReq4UzCAYJ1gdY4WW4ZmS9ERSj4aE7Q8n7Vme8oRIPV70uDm5n/jMR
7LFWxLsxBjshlAnIPR/NB7PKT00YbnaTZb9VJrKfQVRZiSnbBPuJeKxuE6Rh
ddnu40mVl5zrm1Ehfa+D0XFf1cY/Mk/nou2jgOfh1oz516hJ0Nt2c8F2O/dB
PGprQWyt+W1WMCJ8tNcNbEfEpoIa6VAubdSqdnH0/XUvbZ7wcMVUYd38ml2t
u1rEj7kfiEOtsLS9K1UgrBVRp6yuwPgV97b0dgkNkqRVciy5P01+/vRpSzgv
0Ya0rXtszoY0Cni/u6buEgChJm9vonzWdZkNJjYmPLMDlIR6N1YUHllFtFCN
imHSTkPPYiRCC/f6gTdhEIcLRW0mjgrdm/b1ckyBNwnQF1nWMMgbfHCdTOV7
M7jlSsTAE3TkBvGqtDkwA/fyuj0TdmP77zpdaOMX5FXaqVNG8Hw/vVtQE4cC
Hrx8GDuMW6FqsqWRYkJttkp4hbO5KYFW3zwmk08wj6GCKOGTwff8efpwGuIQ
OghNaVNOAruquO0n6AUZnqUVAIzMwPwNrh0auEJHb1+v8hTH96KVQt4TVJou
SDfv4fPl79cBU1YlHQ8d6UmJd7GzurTEYFHmcPh+hYYiARzMMQqfBpYnJEWi
D97oueNvLsnXsKau6MdCb8QoilLWkZ1EdjU3CwaAlnXVux7HUQtoyo+HUcgb
le66qRK1qUSFRfQUOW15mTkzCIJXz1YwVhVwnjEBVsjD0jyyr5Y0CEWfVuOv
97tw43jkcMrmbycvydvx9GSjmMdgl0EUrRry826GLG48XlzkbchjF7e40qTS
vhwaJenbvFHn3dPSQ1oKmn3k9GvTuzGwDYHabP0T6mWPWuuiFQFXu/mgWugv
uC5/YjCvtQR8vpbDLtTXXB9p5J6uI9t7jGfJIuLVkZBq1DXF5gkjV5UAIvnd
XknetFWpODR6Ms80DasmKfHOu4ksrrUekyksxacU6ZqYQy8Ph4V9XYYtuwLu
chHAa3XBvnXDe1tlNJ6ul99LtwV/sGYVqK8d1NMhj/W+nSvW7BvDRdM22Zti
/U57CnrSckSINVxGcDYnXlEGIMb6q8N3sWiPmNJZV1uWvfp1zy+8tbnbseBh
c0Le1Ot7aT9CEbCmwhIYPbXaimmj8oAyFlgq2a56iruqueJGLkGOigArPh6Y
utnwtSwhwXJ4bf4CPN86kp+Qtk4cXQn7CSJNZHI68VY+tw+LQmo4oCNJu8Sg
9JqvokgCAk7jebf0VEf60HZMj2aTbbPuIHjCFgGgTKVm7YhD6N+I5qSIRoMC
3+1GOIBUnzImWa5ktc32t02j+3mfKyfApQaNUuV8A6vpaxKULMP1bAdMLa0I
bjUCnGtTXiui6drndGr/pIl2TG9MfDv8d0fJAduspoMtbSzTRF4RD57p34OK
sOY0rwMazHq8amBKYtcG/y6QbEHflY9Cet/T9kdDWOSUovwC9uLTeWEJfHIj
rff+gR+pVd7aBX8bE+o2eWy2/n18Pg88yu0iNeI2DYEX9K9FJDvwF2yD6jkv
TQK9Wl7TcyEwNojDg7TeHjhBxE9rPlHkoJ0jp6Lr09y5SiBQv4vKRzQeXkMG
1eGGQlXTUhgGuX6um15SddmcaWFmE0BeL8iN0tehsurWfci1E6X3MuBx5Y+B
s4T7qJX/oBwbXWY8htuoMyPgbHRYEzv8W4hF0Ie+9sLqeTY7zGjldTJ0A5T0
Xw22jg76r4t1GOABRrqx9jCzVefIKbud07erVZS3Hdjm033xgmHqW/jptnVK
KsztuIxcwRTX3TAmfwd1TfTOoHKKU4m1Zrj8wMPNjKkDwyDXh0cCWVcKzOVs
LrpbUaMnrHO5ff8gzjIt6fv77rkbs9XV79khkqb5A1Zz+Mvh1bQvYR2fiscS
m3mVPS5Qn83oh4k72G6s/x7q4fG3UPbilZrdPQ/rfKoLJHKrgAGxkr3f9MmW
R9L4C3zS8vvdYXsDQlmnaUV060mry05t32abNkKub5PsgE8Xx9O36Mq0/viV
SebBxWXzQ8xW0jLFOleKy1g7bwVHC+NQw0mSSFe6B5h9TfcHXUGummpzdYeA
eqxtjVD7lPzjxJ3BkgDAGer09W5LOQ3332tAaK/TAmreSUNsLI9ZLwUwVReh
O7XQB3EzjopN09aCqLz0aYMXWVuBNTopJ9e4IuVv7wRLl3/GCNJhBJxSMgMy
EZrtJGSd6iRRZIrbpUqL/EK10zBs2OJtTWZZp2yfKa7LmfF8LH0+eQFe1Np1
kmHBtyZw7jRL+SySOugGfUzLp/vBOxsjEm4oPjcwPLZJ8nRp/bo3BOkttXjf
Y0BJiDUAPB7aKBmwlztxm0u+d+JB1NAXO9LX4rwdXfO+K+XQ54bNU17+WZZG
PYih3SHGGpxMEqYNvz+qayG8rdnUN+YvM8SaZuKuBigj/39WaIxFETQZhZGs
XI/ZDI6ujx3v3cOTh2pKt9/2cnZpFZkHoVQ1dh32jxvPdKkB+mFZBrpWZtC9
KFdGBjQ+TP9/criFYgLVsNkIiqCEcLi9SVFuxEK5pFqvnHv+LgW57IStit8G
riblkPlyd2w2dNUz5CQzdSLFVdLpZdjvDKwlUtj2oz28jTGPGcBLqSHvDVbs
7gEUuq0h2WOJeEbfLq7/4EO55TTx/QeK4t8CpAAeOvM2c3v3EVc1MSoVTTxz
2fd6LKDGKSptEbLIWbwCvDheCqI54T7zE83OEpv+rhqsv10fORbQ6wG7jV5R
qsSoIORV9NRqhJlyN3Fe/FJi6EtYXxUp+VrjxDzJWPzvkT4e9hSI5er007sh
OOXKfJArJg2glhY/xVX3Lgo6UEcgqW7BAgdIEGkf7ulIj7zt0H2BbQ0COmbp
1NpMuiL+roTjYua33VUa7+93fZ/TmxYq3m9OvJi3gMOyfwivocV4kBqNR7XI
eUIMQ4XMVBOfI+tEerAyYIEp9uKXr3J8xFB3jl+SagLRdi01xpI3F0boER1h
bZ7fZfEp0siVwmMG3iCE44uW3NATk/uJRzfAVlabavaI49L5vIrgh/IwEazl
J+Y2dNm/qgRINgJQph496VDgB+FYAVrYBGQ1NSVS9QwYSgh5NpWLKy9qFiPk
TIMnC5o1iKYa83+mfdBDvkOUqQan98XFJk5faoTMZCBCCwIR34P7Z42doAFX
KdbWTuIwUTbHzzAUUP3qW8QIdn+/nzmFLKmvKfrjCOPFef/8GW6ewr6W3zau
qo2OBkrl7MQzjdb0cLz0box+Bx/HwkR10zFTB5s+XGDtQuqljL4PVTlCfhOA
rNqJQIDtmwfb0dfSr+GvQ++BAI2LeFT1TXhe0FmyGUxnRuC9bZH0uICuuUYX
X4SxEkG21oQuFbb4uBaQHHkHsXkBLHh2q3DZ2oeK8earZYwZwhSGoiXUzqBR
2f45+bsXlEVHnrUVsTAdo0vCnQFOEdEK26nKF5Bn03FoaAsZ3L/wMV83n2Sb
VW+QUjxslGPf93wpP32EEmEi3o0OyIqugO91bxiKakyhgaRTP8aXlh9n7QeW
jazIhSQzRUfzpde7enE/V8NPo8ENFaIupK2E6RtJPlxM6wYTQWHAoHfSFbDe
Hpoxq7hDBcwkc+UQPfRpbVqseYAObpbHchBwEov/LsMjKUuTta1M2vJtk6cV
wakqd6yPqhdumo6KF/g8iFgADXfdL/K9YgAFYJFyuvsqDpnwZSYdZgmuHf7W
x/aV2ATYxOMGKj0LYYJhIuGViYwvsb4Tox2/wWTCkxPHHmiKHD6rSPYBzZ02
+0u97ljrsfFFX1KNWn3OcCcIB6tfX1JEmMIzcHtkfV9Pu1rcJ5vUEWjuZR9F
7Zr6+pwwTTlI/cDlA/1Bk5OhwSCrYPIKQMxy//Es/Gy6qbAXBfase5ZgMup0
AQGYIzQmCjMyxB8kGPV+AElIP+p35K6H7o5FfFbFzsEj8KE1KaKYj76/nMZq
jTH8Vytuq7PxQZoMZ9ehM5lmRcy4O1o54sCzrpp+N7AVZ0HmMpk6lDVvOrnQ
FGmlEv9R6QwxVabvycVqDC2McDFC+lsYFGmUtJyb1UWw2n4uX8mqVW9WNtqi
s95JogMhzcw5Bxmfv+uIHnHcbf3/NxSgwGJV5iws5Eve+j/6RnyGD+aqTNhG
RFwfS5Q1eJKLQy6aYc/hDX++ADWIbqnEPtmmoMIydx0NnvE1XSg5kdr2JqH7
LzXcHiv/W6CjVRbjamOXuuU5DiNdU/qliv0USpokL0JHVccQ4GX0f64AQy9J
NkYX5qZXpFFdYiDcZsYY9buYOMH3VrEBTcVfJuRLjdXEz2gqO+b37GkMaIYz
TTdMCdNkse3tT/s+lJAlp8FBU5Aqy7jfCZtalTfNwXTxQp0RSmPSvPHU7M6J
Rkt5wKrWat8pLz0qhrNra18jAWU+kLnX1nwLU7XnfIopyWr7VTlbCn7640WW
C1A409YHReF1Qcx/izA4tR2nHhkvQNFrdTybMHwXdSIIxskjOjLuGLRVWyKf
JmAuivlnLtCytqxB7ddwg/xupV8kAl9Z9wlfXsPFFmcwTgzSeyFhNZ7CB6mv
teWSMfBN7KMcWJHVsXkdstYXhR0jpmsDoE6TSElgRdrq/GPBXK0Uya1Zsevs
4Spe3V9XYFp2hp3B1NYoQDomeWZJIqXIk/1Tyd+XwB5CWJRE/xOykWXpMtYk
JV1q2h2Tkrbow7aMX0IrvEuLXwD7IOMC45C5cmKK+FpVs0j2gF6+E0d90DLv
NLyCAKPlBi/f7LzlONhdt3bqX9eiPOL7k8aIrfs8LWk3YU4paIeaSLxaoPsT
4Q3W1J+KExXhLzVIiM9HbaMrRDaiEdYRT8XcrfXcjkvafjoDhX0waAGq3vlm
PBNRIxus2Jy8iTO9egQ5RR8Zh5hZ1yEDP+83VUQPrt56e9vzB1qWfN34x0TQ
b4n/EXcyGZ5cD9i+CnseGlSOU/5TslCuzauEGjeiybkmoXcKDnlCmIONUQqi
j3rXv+O5O+SBTXVFzMesr0KFL6luaOmfdTYzZt2xixyVsrVCPnZvZsgR+HMH
rSPxmPKCCo28vk/gq6y3rhtEgDktnnnJo3gZyGP4ZzNImWLXZ/QTPnFZkanQ
7xctOUI+w00PWTJCvRRzlvDjv56Isnbm7I3jFHzuvo/ex2HRrVE6nG9m/aNO
Ikl8KYgdvyPMPVffD60WkZTSD8Vi1ywcHR1W6CF7nGzeGP3qCOO1hUx61dYw
J3EkUFDwkNdM3JPR9v+h5tefstp4BCSNmoGbxfQg0xC5yWWn2/A+XwUh/NH0
/wiRq2TZEc4Lb3fhAqxrlWmRdZiXaHOPl5vPZVm+6TclY6V3pGLIkitErF+L
q6ALL++1D5IaS8SwlF7GfKJrwD3bDcRgSlX2NYxIMg49MPvZ3O1W2SCt3FKB
3G4F+zcdSqao6j2lMH55+oVmOmCrBLChV8gKk1BBqAqefdPyJsD7yrtbjkft
N6g7AATe7UOLOdURwrZQvTBKDAU29fVc12b00Ua9R4HyYOFvYzuCMxZ/QEok
WB6i0yeXGG7fjHYLuuQ1mb3sTf9WKEKJ6BADiL05fLGEPP6+YeIN7WtkAnjM
M2QtPulbBtwnUjqUHNea7ODmTa/O/5cNIX7r75E5MW8TPn5v6GWHTFiPNs4M
Kxrtwm9doXzQCMRoxzpkqQSKKlgpVRqr2KRdo5a4dN1hoYnv/q1jqUhgGaet
C/Zbio7V4UbhiXFOmRlSxSC/BI4UfUYcHcrRLHVom0iUzs9VQL0dh4w8Hpdg
76Dk8s1c6OElmJj1jecXWyfvBW90aq11K/m9hbX7o8/bl987vDkk3RtheuF5
mdwWmOcOR+qUCOZTk+ukrP8TZY1FFPKYXuATseUtf6l6NiDfM0STFYlz8UHS
D/83dDRahoEw9qh34OWAxEY9xzZN0Kox5jVD2Mp0xySSv8C0MPQ/GEv8NDbe
vv/op4k1Syw+odkcLG3GUeuD19Nw0Zar3RQ6PlnUm01RgYdhd2cSm9wUWGHD
qsETv8C7kqL6yTcqmKjufDdMGhxSH3u+X2Lqtla5govCRV5Q+SY3O0yM3JsL
7BKIlz7zLkjKi9jopQ6VXjnelizqWdU3wV1BdlhDM4jc8rI/UzUalqGlYeVO
BHFsvpnR1CmWaBuBE67SnWLy79peN93W0GmxTNBC2BYe9JBXDotDaWZeKn1f
QKzKFjyBi7h4Zjw1ySwTZxc8Pb8/YuacqXpZLSYA//lcSURcEfUTKONcNZds
SJIdECZdB2o/vnVoYpJb+rsoo8LtiPMDaQZ/U00SsHJx4p9cDp8C3RFM8EPK
QQ+4l6t6uMlyr4JN8jdJWwTRjKp8xjpLpCGJw2jaXbUcXh9LfFSZaEzCfUT2
13Y0zEc1Fg+R/K2Ws+B90AYEq10aHjP7RirXWj+14bU1ivJ8FBpQ6g4fylFQ
Lp+ItoknViMoLUBEX88J2yFMx0RdnCC4LR25uz6aFV0IFAsy5+i0mbEpe1H2
FVYu4WpdTjPqmdAgXZPtl7yb4j38xCY5kWm6MocyN9Cua9hRrhpqVyMcJmGp
fFb1E91K5c43ZnpsyZUXpZbbmBGFVj2utJTIF1oORbTqvr+tsmFfzd2Tm72g
alhy+KddjeHAVMTMvNXnhXQR4xFpT4JYvGRUSN8eL7iq9THSjhSQQSUPry8V
2d7tN2dseEOV46gZn5PGGJ6Ge4i7zTN5GzlbcoM8AYOkTsJfMS8MdeDu/5HE
+1DfwS8Lz2AfmwPvqbwE6mYWfx7gpYMu6xvk0aYpbpowrsJ5NhQv23Lj9DZ4
NStYv3HL+ZnIW3Iforywx2cjORgQ9bij0rFXhqh8fZ5DE1afwgEaKh3H3EFx
lqq4WbnrKFMUzpr47jDPC6CxFixWxRLSlWsMYTU2dVOO1juK9ccZXxtul02o
IgoA6Wc1GFtk2vi1DRjB4YCHGSgvGTsyLEXWZO978xG06hXLtOeXBKZIlVqU
m66tKfKWkPJuRkMYDiCx3lePLvKnUCb5m0hM0ezNylV7dmuHIlEYiTuSzjFX
hyT9er/I1IaX4Jm4TLZ/hu61NxwlceSRu6rUqZ6UcBKwphrY3WSyhIGk9+xv
zA31p/jm+WwG3oljwp5gPo2th7yBqCf5bN9dTWX1jjkXv1yBLchgFlQSnMDd
wRK9flRcYEz9vddupx15Ryq2dn5WpcYJfrfte12s46yRLiEVD4tXar4ErzMa
F6I71vkP9Qvi5AWfEJbsfzFRlC2vpFkvU3ABBQzcuvwwPFjftmt5yAcUlxzN
wKH7AapbgFT3Q7yb4Fih4L0Vmg5UaHO/PKVkfgcAqBPN+m5JscgyaRpQTPvb
LdVDZp7OH0O4ig0nFFyBclhCKVJfCV/N8lMcEdHGrGIf1UZR/96RQ//S9zUZ
w1OYvjveoc5xqoIdJen9NDOwhog/FKjeU5mbWAfrOh124D7FTjH9f6T9at1E
8jGvyJhOW2RP5L4chIbEcYV9QcrZ/JtjxoQ64cCJDebrbvfDBIG9uabeiJs2
TqFONd+VyE3ZebvXyT1OdmbKkvde6X8H7F4TztNfLH26uyWjpoSo6FP2mWgZ
pcW1JUSxUq88iCNWFkxnoLBpC6PmhYHgpycivELac4O08Gu2RR7smXP/lcD6
fsf3Op7Iu9bDSac74KxtLDfmvd3A4R0/x9b2P+MTGmSJxDdOIFdyzpVpD2m+
/RQgyjmOwZEfV0F1gh2NiCer3LnbSGhcxwIWTDzoWqgG80yrWjooBP/o9WRy
t2c2iw8BwbN8Rsn2NE8DeDfr2tNWWr4En4oh5Prte65q56YBROAKniJwK1Ds
hyfaO+/cChjKEnu32572X94JEm5PAYOXaVfJlLC5cziqUkZp7sD7Nc7DQo+r
MUabVESKOfqdGUcNUq0TfKeH59NAaOqIpWkwVkqmcaYbmv/9bKIDmNN0bGdj
rj/GYZvzFloCjgYkW6xJ1yoxxUSyCLtFOWIqsnuAY3x61H8jKubbSoryxe4a
d5KC0M1EbU4PNPzHpKZL9vkloJb69iq6ribksPavXlDGrwveKbABt3z1fSmP
uRZMvJ+fagwz5cN7VX/2QPHjstnJevOhezZHoCx6dlYtJZrRSa4N3IGNzqLs
5vQ+AP2MMXIP6cTzV7GCwgQ7fn5cH196qGptQElI+WZguh4oK9de5Annt3Y1
Av0nME3tsOhubSKgbrQ1ODcAX61vyzkYl7MfTMLj3E50FbW6P7EY5QXIZSTW
C9yYefJm6xIl1J7lXWXXepw/oGPWf91Rh7JLhLqe8ZUMRMQHIEIC/6SWIaVy
6vBg3NoSxH65vtDaiQuRiEdfk3Qvfiu78npJSESXPub1kv5g0dftSQEm1A6e
W2+tl1qqZA5MetRyVtTfaCBY94JLHiurdlC/7qmgkP5gXt3/SXwOUxIbJuXY
A/IsUvx9IZs50Iem6SOUwJptSJ9+CzQUXQL1SoKjLuhrZq4qQeqszKIj2o59
2ZBlmosO7qB+GXF/rVLKlxDMknYFfOK39D3SUccAgwkL+zVy3/P4qyyJp4e2
T7uoZ7onzncp6ilkBFb+rmYmNMZtCwYhQiHUV6RtEueUdxc5AlLL7j2GQKwN
EAVBf9nZJxoDsVtwvgnIyp6q+AD0Gb5YfNtiZhbyuoqyFAYTMZJ2WebHN16N
ujJLQShYP6MiNu5lgxKwE7tjpwiTj/JBWwWC4C0QDRr1B/Xm3cCG/cec4PLF
6Se4ucwjScsK703vpNdlJJrjGI9m70u5M5uJeVvwEcRHwheeQ+eqGoMGjKr8
KDfV3B1P6bc6YxqVSOIeWk5PW/NEetc7SEae6e9ZtB+sHTsxdXkvfwd0tCYc
agFx4KLMyd0iaNmhiXyPT5gj1je/4FmO3yAu93HV+MeBW3DphRIr/j3O07Kq
5gN6etw/Umnh39r3Mcp5gNAXL95ADGEVyiGyJfKtVLNgx+0F7UAOjxtNVk2X
ENg/PK6/PL4YXjWJrsUAW0FtCbe/g6laWCp5rIWa7jBsMufQJE7rePLSV57f
r3c8b/DdbLTaB68Dj0JysEoNfppQMgS5KmnA3T1v+mSp7doxhoFUX10VmBQC
emWASP2jsKXlXUDuXpa1eduzX1jqjlsFPtBevMBJQL+2JLJE2zJsmEckEtnV
3rZdr3r3g1SIOlrZXr+ax+tvJCQ7nOQFJN+ptYtecFJaFoiqDqvD+o9b6jmj
h2i6sZRyRKI7JB30ePWElkMQoMsMKWqALQiTU+/F+wCFGOal698Bor63wyL9
goRgLxN0FbzejtDyqKfiY3WaeceRnDeJTBPyS/YGT1vVHU/+1bweVpKCat6B
X/vqviY7ZP8O/mxHhCSi0jjzBM12pz8zJtJbrKzQZs22w5ktta7X+reI+dtm
urauj38AFzFxy1gvoip8bHk24XkTYvndycfmMacj+aHqul8DvEIhHSLVkYzp
LfszdnUkYirYZSJLrHqLcIIPYWtQHc46m2IQa2aPvnM6zqEa+nH1oyi/Y8Dv
wRNaVv/XKqFNmc9PZjFNTMObagAHpj+dEvwiccCOndQs1beVgXDsImp1GP/C
zh1DaQ0kIN52ztPFOEbg2iW5spK1oCo/8kZx74IYelKldOcn2fZhuc2CStzd
UjnK6FlEaXcEdLrQe/7JfbUqEG2Klsd6uma8trCVbHOiyUR41e/G9sLSYrSO
2keI7rvOpcuap6t48KYivTnmMmcsDnH7HSIwYYZxEvec2Nj0+9VGXg4SbcEw
LjpAblasgdYfjF7xcrfjhK2AJqfdA6t0k4V8K3yZt4Mtd79W9QTu6zhvegwL
i7QusZnncZY6wYfaQRrfA3FDYfqND5tg/ZYlts5lFDTsAiad5TF02WNREQiS
aSi+dTDIDyR+yHm08brfzP3tTtBLWg+YSKpl2YCEWz1R8frcW3VLpN+2MkdW
IJZ2BQyOBhhiofgTuRrnnOFjRs+aRdsdDOykF0LiH3LUVVSLDcCCYORC3kZI
wvRurvbxwwsI8iG4N9HmgAR4ephtGgVjZnee7QVN9AI8JD/Qhbt3g//WlRIW
HhjQhsqWvSLeKZWwuKTEEu3VIJMOaHq5+egnM9cA0/wwhh2cVUlY6CUXgg6u
Igrj1J1dUK+UasmusDsoYxDvd5ugKtmwVtAbHvRaT//B9/lT23FqV4yPIRk7
N86OBNz2FK9fBWpimYE67sNSz+SIfN+bBUDsjO1O4oK3aDOewtkRPaQpi7X+
zOwMjqQ6rjVayx4SeqAn1KCo8pBV9pMSLgTBNxD36hz34zyik+3s2OlbkBmZ
IQv1LWL6SOKsfhxRLeCUe9w99MOoN22w810518wMrP39pD8GesZtOk8Ljgba
4BaWhoSc3ZflkHYGYoXQOOfIZh4Am+o9tuQ7WSvBPc27944pgoqBZ1F+GHjE
eGilaB5z70QLZFbp416RaO8XpSZxNwV+RVgIfuOpDOQ3nuLkUE1zwwFI5Rb1
F/b4BrCLqyvZSh+gQbyEiq2F7CUkA62oPNax4BlCuQVBVVob6lSYY5ejAj6c
sZkAgvE1+R5QH1DCvT9NCsQED/2n81Z8WnQBMCQvzPokrf1y+x1hLrFCokJu
Kuwqji1DzLct1bsBwvFrksHio507Mzy0Cqwi04L7k+sOytSQavZfaUnePMXF
XFDr/GtOv1pKigwfEYKL046qcJLCXzm/Qj8Dj0jGYvji4L38vABWnlIG/Qys
ORIUDj1VZKIUJbpNRE9f8j8Xh5Kpqq670Eg8o6bHC/5+aO1LszGXGGf/J+Go
TnJUbuchB7QQM25l60ilImlv5kL8Isg6sTQaB1gJ7pYygvBNfTOPuqp/RiVH
/fB0Ghw5rC85J31/U00kRms9Nq6ois5jW7JGG/H78nmgVBoUaIfTBzhgWwwp
WX1l0MS1w1i7UCy9hFovzbxjLvohBroy2980H9ufSANATC9FzUWmxVObJqu8
XwtT1N9AdOID3VV7xdDtRebbChPEbJ1drsUcR5V1hyIgrk88wAttdJ0gCkYj
3N+tymUrmoAzswe5MYoxxlDwHK5y+IKJz6B5Y0sQLpXOCT/UWfaEl01tqWZf
tuDy347O8FNP1NXEL7pERnYT2CY3GVTeMifcuIXz6cUMSefl42gQUkPlsrmH
QrolFotkzGDBzqEB0Cca8zlf/2KiARQcu/nQ1Ha+t71qJFi9llJGfke7gtNy
yKCClkwWsEcuM0a755EUe1r74v7Q3vlo7YOcOlyZqM6VuCN+LGbRhVIu49TA
KSFeUm8LN5c6OmvjKVuaRCk77LNNxtBjMQZqakV+jx/ZtPqseGRymrZbs9RK
WY3yYuwwjB90PK5Cm7ArBwonAFOHsg1ZtJWOK396d9uVcMcBoD/95anKD2Ew
+x+z7heLO0bIcBnLcypwxO9qXUUA2n3pvtyDwGspf5bsk2uVMo6O1FxFvjRw
d2fe09kdybZeqkJYfoktvdqjKD+Jt1PnI7/E6Tu7s4SdIamXYT1DF0RXxHEE
kUL2ObDcpNj8zBMn7+Dvz3WpmpwcTyjS3qg29DdgMjOLAD8smdCArfPigAB9
eKtsT//PZxg3QJAAVIO+0715rx7Wgqnlak6lDaBVipSAgQojq68wAd/JKOce
eqbc38fZgXUrfQbJCERqazYegx5P8pcEs0fBkkBU3vet2c32rngT33Ws5hUv
f7Tbc/fYXhpMyBjvO4u0abrNqFT8V0nMQE6no/XHz43obDfQdVykGAjlW7TV
Hnc80ybxMV4i0S57/xs9h6L9+3sxgaNEvYUFceQb2Oki1lhVlMzh//OOc1qV
wcL1l4Qfky6vWeo2xxQK8oUDQ7wkWB4h/IkIpIMSLGc0cDdUGlHoNXY8M0ph
5g2IUsXhH5PFiiJgolnrAqaOMh6kCHy3gOGwQ4hN8gFoK+TFP0aIV6L1uFTQ
N3Zk7Qw6QN/RSo5fEIV5MMZ0xq6DLeyaTdRcxf9WARCwAHmAfPzLc7CDrlUs
4nYL5TkbAN75S1EKeEDpbw8x1bTkhMD82qozs4M/Hykd5H0M4OAL5Vqo2lbX
YqBwpKe1Y8nraeyhWg1h4v44A5QrRHnYrYFb0L6SCbmWKxF9hpNHwRCPScHY
devhI+YX24tWj3nlch2h9aDzBD7OsuCZJixjlnjP93f4w7SlQmfdL4ie+KfA
gZ0TZSGKz5tyjoXEokzlPj8RmjbsiNCdEYimMDHE3JZChrmM2b/+U0LgTpr3
9DnWM7r7iC0OsTT1s05eVd78yUrHKbgXp2IwO/CuX5/dN8auVf09ZLzLKDyr
fgOlpbSsIicm7BjktiBcuyTbErPgr3onlbl2LKuRd7LrKtAuWzp5Sgm/tPBm
Bnpb1w3oCBmWH7s+SWN6VVOUOqN6jpYW4MZyfJL64jJdx49gSLyjTJxEqO2F
cYy0W+quSuOyaZFrxjZQrXTaIHfqcN744ZZ652MTw2S34VN7o2h9gVnh5bxU
0pYA4gnCAa76I0XnPObylxPqYxbX7P6yJu3lhvg+0wX0cJm0U7fd1rumBAAe
/bQov5zJVmwIFYphckIHBBLCgRdSrBfYLKyiNkBvIVzvX6Zo3FIvlkMWpP+M
q0ODap9sj73DCzO24ijqyGOPj5gCMpMPG9EDBihWsvCrlKKinOCM/mQjkL7+
lce+/Ae3H1hq6iCvfIHKjIrvo1Iy2Euru2d2+QgrE/+aeiQTRCa0wmsqfVMr
LNx3OvEvbH0eGH64tGTntY/cS9l2jhxC5IRLaDR4xxDAaovwTRiidfSS7m0O
zL9L1uqtSGZnUxoEmtZ2uT935EI47wLYPApdPGc7IwLJnmnXgo+27tb+UOiO
fAPOZ8O7YoT9f8+W86aPuD5JRrB/PcOb+6tV2EKm4eGgPrpZux9UFg/cxvXg
bv0Lp+AzQ6924w2xxwPzzQTrGRRBs3zHrfmM/I3NrHW8dq3n6N79wYwJfRcb
mDrx/OS9/V1obwtpI+gzk1J9eaTwEIKfAvA94DRsjgSZxLU2QYJb6zC9+uzK
rVx9Obe9GDhs59Vjq3/p2b2b92e34yo3QGg/KtQVUGzfdWzDaogs/P70wqqQ
PZjpPWmx/9QDgAJz0+QLOGbc76fEtc++9tYq9G9DSo67tyyizGZqbU5Nsx4o
GxJz9LVyBZd+IDnlk1uUB1QWA4K8v8P+0ztcz1yZ0PBENdkpAjAeCYyc0fQo
JljJjhph8bHOxANIBaxlzRi2wbPPZ8E2ueOs2LRAT2BrwmQxYr9vxouRtHaE
h+9Zu0Z85yS2R6Uk8ZUs/CNlUIuqSYJONql+ZpDmC9HChOXBZ7hlMZ99hHvE
SYDM9zpvCDKWaHFOhYJdlZLbcK3i6wX0yN5WRWjOKa9MUBp6op5v8tWeM7su
AuNkr2AfQpKmpnAFTYxC8LC3PzDx5U1KtJ5mOR1XN9sbyv9bNTRHCI7PkVLx
P5Tg4woTlxCYKCymfH0oQAFHWvmjEDZqTWJXP4npMHfC+k3EB3cdtmIfmhQX
D1LZe5jTGI5imMnGiDIQqBXR2VO0qGpVD9wi24mxFfpqE0Z1R4ZUGPZVfUlS
5cZmWouVPGiABe3mpjGn9iuqXCaSsFoR1jAUTA7B5IpJyT6VCWPByVXKIOJ8
1TRV0IYPiA7tcz1cZ3LucV8FJqAIU+cU0X70zjiQHiIFGlQKUF8geRLU3lh6
GLe+fS32Nd6WEjnzSEK2VhGC9QCAtun4lphzAfhG4HXCu1shdTccNBM/j+xp
GoRP2L6YJKaacIyKPEFKrveLzTUlaLuqGHrVKFHGI6YZQodpFJRxm9feIeL3
xth/MUYGRDvrAIiyROwyqi6+lEGCpkooY+mlUgkUh4mF/mW0jOcWlN007evj
CLX6QC6olxf7+3xXVZFJjHsFo8J5XU45nTkAP6Qoew4mkjV4yXzNfzhEP65R
xpRTg01lhdiTj+FVcgA6XTMAZnI7QUylYM5Rmidylg+LhwT2QH9i1vRyLSIh
Te41yeJSf8dDdkmtZkB27k7+m3zFlO3cbmm1yWFVwm0kKOGKB+yE0KME4qXA
AvbUAESeF2AEERgceHHR7UK0hOpb1dwbM8+CCVxKvZ+FoNb+i7nY6ETKy/P6
6ZySGMnn8KBhkTDoRN1fKSTpRZ5FH6Gy4ds13cuhiOKnFJyK7yngYlwOMaiR
xaWDA8mO3cvSreKDvSJ+PuKTQDLR78svxqaRCjIuQL2YZPWi2N96GaW9C53f
4uDySLSsX/12DGyXMwxVjULIgzW86tvPFBG3kW0yP2WmxnXVtje4OGugQjpU
Ey27eYdaRwNCtdVcjgt8OKsKb6F6q9qSR6856YQGemB4rZ+ZehU6+md3ksob
UsAnY1K5pB2GG9RvKgBSzrLHtecLEpwrMWu5ihB01DM2qL2AvE16APeT4KTR
DhjsGE57CNR253erHSf1c/YRLbqYm202Qe/kIEIFT/nqFMHaf9yJstWZAcqt
5dgbAPZH9bn6jK+TkbyjBP1dUbcgQtLzDmgkXPQn6wJ9TXHtXv5Yc677Mioy
t24NHXbxp0Kf5mb9ywPCNXz0Y3r9TGlukc2e7gWTzWID15rdEPOxdlgBg++N
jlvhs1eodePo2wSTQBCk1T7PsNuICuEpTucDAXwReQ8/FmO2N7Z8YIqC/F1f
PFQTsisxMz4kII1N7Es7PNs9FGZxlooSU0vbX/GW+mpvlWdYcyLg37df9jsx
VgVBGjBpGEl5jpnTQFzeFddU34KqImbp4NUoyH+nTIRs2QitkajWZXwBVGOk
YbDLQ8sEtWzOujq8p0ynGHVrPCCSvfyjumOwIimNC6XueWUSPYMTFcQU4vEN
m/IpbmfiswwNRWA+1/SZyLpodHt7Nn3bx01n0J0YsF3KDd/n/AJwXx2pa03E
z686b1W4nwrBRwaNxlbQ9FmOyh6qjgy6qNvvBq89ZreofNYr2neM8u9jtmlL
BaLb8QJMHgrqyIyFFqkA3tfGZ/2yFnRkLFhpXf1GwabxKMJSuq3yIDnGlKmI
f8poyemXs8cxGg9qgk5IRKwzhbjz7WhwWgUmRqFbF2ZW8jwOMp+dbySiPS+l
2uU3L/KSOSE1T+sOPhyoD4BMAndwUMm4np8SgNzXfPqK/2kahtM8Swbz48sP
ZIumxZla/MXya5iSbtiC784/betOF48q72DXCByAFRuPetKNiO4Ux3ZxkD3U
1x4eCNuqIVQXQRW06LhTSlu+HPc6ESZJElnVkZvkoh1c+UaSdD34fHMA5mIJ
OxD0grIGFh9SyyPF44PN82lN9959f2ydYAaSwd5QrJ2lmWURFRbvPBTWaqUB
qWvhxldfO70UAmGUScnRzBf4srLsiYFYs9RUPvNzxrhy0WVd+pJ2U6DZEFzk
ZVmzMpRYYSZUIjZviBVU+NvTmQlsnBaTr1+bpXVpoKUFFSRwIWGWFAwpkCjL
zCQcgKVp8UuPLN6ymR9nGeVk1OHI1jJZ3gs0PsKCubAain9m+nRfEWF3Pepi
jMA+Dd2hrBB0k90d6/vqm9hU4Yg3t1IBZG+y9kxA92aaOX+OItObVkVAOndz
ErLMTKshcHL/Bi19uiUALBkg/9QAeTkhPnXS4ksNyLqEOBOYqsruNaRKqcn8
U2P+GNafXCm3zsTeo2Az0NJe4/fVfS8ol+IzL2G7s8Qngrbt0p+fgarOVA7m
aDlnf3A/P2cdKHanC+U5mNnKeF/fa34leyZ5NQwAObpb59Xkf6HrPrsUwO2X
1Z36MMFwQc2UMDmA8UYA7JosN1PlpAn5FjVyCIl2byX90ZfSUivumI5spL4e
rghmv8KM4HNUwXSEijDnsvs25W2FZnTHfg1IxORpe+lM89MSgaubRWuty/x7
pee9v1Q9G9PPUzbYuj3IrKQ4gZEgA7WnIPDM3rXPUIuurqmdlbFw4To+LLph
n72pXhUSMmb/oiV3IUA37g8WOVVnpK6+IFBGj8gnPW1uLpKDWt+8jtT6LoMD
dgTpOxKDPCwWRvjmlWHAgnzBgSbchX1uwdNfxM7PA06zzvEemJzgtv+0SHlA
Ailz3uBNVSS5l7EXsuhthtjEcsfiRdo8ESSl0CCbZW20NXMg2bbJGg0/DQlX
9hjc0mNz1voa5RADY2uNHUxBYLCH7l5H04cejhTmdmc5PUWrWVBc/sakfELM
GXHT5lrO3gV8IIfMVfy57usm5gHyozyfWGgiIQh/nzC2m8aHruATroTkiB1q
Qt9m/RXhJ7wEvmQStTfWDuWDdssdqVyVXN3Z6qFei0GTOQWiKJy9uYPylknO
uW4IwoTSDMP25wB8zoFvskPJ9OM4grB5+9E7OKIFwsqmy2ZtnZudXvhbUOSN
4K1wX5R2R19TpRWmWqYptAJiG1vt96L6Rt6s9iRLl6J0+6qgt3Y0jXtcHa5l
XqGqFOdr+F+GxVwE9mn2pWrQgrLN97py6Y5hw7DqdSzQ0K+JcHZUVyHiUm4n
yb/wP21ItZZzFPzDj1csU+qF7PGNoQXcW7IcyDJiGX8XhVYCLjkUgn794FIW
QLYx3qify8bhl+Vei2VPNXcW4GjhrtK5w/p6xjJ3jjOWI4ZbP8z8er7hvrhE
NC2hoG5jfYEIms7EOWymxo4LIvK7dW+uh/PUzCojjAszmnO350R6rscuOgFE
RJVIiFZsbTYl61joRr9LTPjREPwe2e4ARjqisVwOhDN7Wnnsp6Gd2y470GIb
Lt2OhL0qYfVgaI3rN/LT67Ju/ZP0VGO4+cNk6QKw5STegQQ9gdMrsiAbu5J3
0Ei+elY8l0Oum9LgH2WTHmE0H6TkRlsipdZeh3XokngkKntYYzBN0jYtW78b
PScTKJ4bh4edSVtQ2PBpFn6oCB1bzRSSSv8exemdebP/1SCoGUMtIjS9BQC9
lKGLJ2XmfKdQmxitI3i2gBlq567dSBiqfB3Y8be/8PF7Fq+k/PM1CKm0Frdo
SFhYxaHzIMJcuVFiK1sgwkJdfOJxn9qvM6HB6bkl+iksLmYlfQ4hnj+3yAi/
v/8uoD8E35nkVwJTQr1PHq6LMq+SGyxB0Zh6ViDxRJzUQEzLq13kPOn91tGq
+DEWVZo4RPDOSHhyA0qrOABiu6h+T3vbbnuRt/RstVVzgevSz0LbEH1VNWlA
Zr61F6KgtOnYaImeCgrE6JImIuWck2fD4a0EtbI0BI2JwupcRo/sWZ1qTqMy
qQvEA8rZ+Db4/SFwn1RQM+VtbgC1KJwtyGaeMN8OINOb3j8NC+DzPG1exhSq
wWOOXb2W1WHU74niMn+GUor0AIPuT9+K7xD/D8bL7XmTGTKqomds0G+dokdS
F2gvK/TRaZR89nKXCeJzhdtXKz/t2YKpWVxul6PvGVrYta12folS5tPP5Cs2
07Dv4rrJSESWwjt4UqxMD+VufdmRG73RBMBPpz6qzMqOJiBFAOz/Sj/t0gDH
LHrQ+l5/wvKM40VDxHJwwrViktb22WQmeEnwnY9T1nF67PqC3Hpyyfe8PuLO
VlSrOECqhGrd+7OnC6vb9+7YKdU8n3U9QI/H1PKGDCopBsWDFYyzCgHE9WJv
kObJSnxKLi6Jj0h1tLJro+AlYHmZB6NctKxT3oDYbf7bJ1qP17Wn+nag2ytx
qoBkqLcj/6DJUz2fa2AZYgVHj7UVi56yIDc5P0vgnn1jW+0TqMvbdFWqt430
k6x4OuCmy6MlunwF2YjrB+BQkb67URBDPWfK6BB3CPysL0naK4FukZW54yBt
/CI2T+knpWAKMYe9/O+zZ+jGQ/uYgpj3XwcfqSS54UD+/AHkxip/Qq6m7a0x
jen8ibuJixf2O/8WjW2fgQyN1eEMsbMCxpvyJT2EOwXkPgYpEifS2w/fyudt
pbcUfnLOyekNtOtpgkXvuAwyIF7C+Wg5QC6pitSySXngDEwcBPBqCrpa67GZ
cyl4xSZZPNY0P/PS4ouPfMMSa/DOUo1ZEhGIOa5nf+HNJo4WWQvelbGHgmU4
W4SMZGbCJjxkcJ8BA16osTurd6wDdf3p2lgCbtgiAFqSacXSDT4mI6SyfuUd
881cei3jOrm/O/venzsKaqPHm8SpCR1etRYkp32bpcF3gti9UfKrQQbLihYm
gw3/jOs2IfXRzyGpztYHlv4J7PxxvNo8vNveHaR8eFBypjTZlsVEtAx/vUe1
EUjvTp0ySroPM+Mg4iXEUJ95awQTBcto/YSIKXfzYB1xGXfjOeUgzQKmineD
9KJGu9ee9GAVXj500ZZ3XEKwtkoRTv1xTrUHyhvx+e38i3B9aCyCzRnad6oQ
JocbSZC4KF+oJGcj5jx5JNtkiseTn+aEFLW5upRj7psqdh6VSdwGPsfesmCK
sOvVQGqy7FvT76ZINbVFI9vzwnU20NKDXqzNTMKtcZNQnXPiGepitA61AdHA
Yon/MgQnsPqlI8r8Uk87GE5ww2IoS14lLntG/lfy/x/jLGn283QbXu87aE9v
zq+aFvmA+u6HaMJ/Zu4xSn7IUEnOSuOnbktOGVN1WURRiq+iedQirdEmnz97
CaOl3jI/QTXGorF2AEkQq9pfaZI/YF7z88/hpgvXw7XFG0BdV3tuWgSffNH9
wf36WxLaWWtsCYLptXPpgekkQcocbYkCBH2IKhjU3HDeS5sBttusG8tfB0vq
UaxxSEDE3Wo4Vaq07TNkHg6GosnIaYhxDG8u7mlnW/DnnRUyQG7ULn500ZbE
JH2yXZU7G+GUpb4iV6nSWWgNVvLNkhZ7PewcJraydrEANcniiz5kbPXbfPE9
8lmQMca7OBb5l5+Zpi8TssUH1TAEKqFbRPvr9xXZU8mQ6iF08PiA8Avb9zLh
CEhy/fweWZfZEyTqEUc54cHc4OaM4WIKlB3Rv9MyZ48o6kmvz1aPrgl8DiJh
E0SB+yWb2HCEmd+8cwDFtfgIMR72BxuDVZd2jRTdw6lczpLM6xvGBc+FN4vm
Edgffo2aAiRQw8vILbT3GF0bb1tfH9doRO7URgE80qfmzlgCG1riaIj2sKmg
ZUyb4yoEVFRXyUPU3nGltEwuXVDsBBduqE/5oXKzjI3K9lEcbkHL0d1beKqF
r8er37XGmHDCYb01Xpp7y15BxP3FyBp18t6UZDr3nfj9oGL/str1e+IT52F2
HHzxlsni1c4J8G/n2Go8/Xz7X+QkNFn4z1tnXYLV0ef7wp8MadbAgaImtSX9
ew40dKERDb51mKi+ArUQTqHVI8pZp67fnXiSS1/i1MS9j5pIrEOecwykDv3O
qbwBRqB8SmGfs+wU01aJx/vibZuRwZVzRdU9vhodD2rVw5yRkStcvJZZPiP7
t96CZqsgtmHd6C2kPwiITphCoIz5tfmznPiYF8BIYR18oe4ppAopHDnElCHf
+gk3ibvbLLYa31OhNEu2DrP5UNFf8OpZrsKXAk5rRVdu4BWPxlp+F/kw6xRa
bW+nqKMyVGBbUxEMbJf4BTaBddOModAgx39hhk4F+Cvgn5X5+WPHkYAi+fCk
dH2q8zAYvDXOaIq/beEUsWwIcU6/yZmr+0mZ9IafsnwIzE/XTC3RqvS6fFcN
UeVnTh2jtkXM0ZN93rzAvTPXu4lPkXfGCiQIxlKNdOkZWHmiOBG/aKI6zdh5
0KhTLxBXClxgRuVpslLpT4WozfAJgrJEx+vcO4lK6QaBiiJz3n6eF1BOPbAn
VRqBg/vKFYk9NW77ecPg2DyL8ijM7GFfGynQEL3MwpOsOI0PloxfBaw94jI2
SkHuV7UhYA24hCr6i4WyqogSw19wnJ0GpX42ncNfUHxIQQrpOeSduO0xaVOI
onOzAFtV7mPC/TTX1nLsGFSZg/qkBV5/396NYoo7VmOWkdeZlaZJacbk7QzM
tZe2VNyORLaFwdNDcOD2fl5y1dwyiXsotCjP2mOlipVivccjVOX6/ykDS1g4
GH9EXVFusIW1tsM4zyrQgyUwd/QHZyIYnEIBjuVnSBF3ayUufO3o+29l3oqy
C3BcjqLvyzNawSPkhwbjT/e//p+jnpsPq9aOIb/R+dJQpH+qpMxtCFSR48FC
HWO8ngue7NeZNQwh14mwZIBIQw5VozdTRMIONYeqkS74ra9mhXG7HEksvpc9
DOOeOdhrT4xyiJqXJCzuwrObLc2vjgPb9Y+p6yqJrKSd/4IjtR1CaZIn/T4K
/ZVbJfv8kNrs0irb3pnWKdlITch0C3ZDWoxgjj2w6+IlJG2/8fm3fQYGkU+A
Ij8EXir9R8+d+xN9D0EhXVSxeJlNLSRGCjX155C1id9RvUbLt7xp0AdBSHMh
JvOvmD+PnpF/qIsat5oBM1VyWhA4dUlMX//pddq7aklIpCRMAT9aoE2pBR6d
poxhf3QwiUHv5Tdce0XoZeukexrZU5cHEv8BDHtTfLOQsCHZw5YrGquKPokp
BSmruilqVhctaS0UHj762kewRdUaWOQPNB+KkbqrDin89skEUkfkFoH6GJ+N
U4ISL//9HDKUtS1gN55fW8LcAwOxl5EuCcqT2nC5dEOrJNK1VI8Vj90/4eIF
EtP5PCJV7K+qZhX2sVqU5Bq5jPwRX1z68SAnlFbkWg6XVyqqUjlocgHNYhE2
f+nnEcGHZM8TSTnVTH+5dQMVWTQtBcm8wmuXtXfjybtgxLcldT0LG/IJs1+S
EJsyFqdCd8cbgEy8GITO22pXRtqECRN2WH7JnfRmDK8f7Oxqwvw3kC/Ne0p2
rCG5R3lXJ4B4TL+YsDmk6mQqHr6HZeW/fWHYsuJtatVyHnlcNlb85jgGTMIe
byThpxV6z2xTFWoXM+CHGJgeAKRqdvH6RhmGoLV0doxUtQh1vuHXMvzcDXjb
mg08dUq8TZzrwSO1w5nByKSaq6H+GW6HPT1PXH2D+eB40dlXG/yqyjpY/cgI
rbFRAq9m+mApfj+1paPgDQH0Vq+vYK+tE/g5COdgrgUwNsqoHo5nmMwa1G52
N2Bn9+p2VouviPpeZpgqeMl1RjVruxte9lXxo6oU1u3kpXRZkbScGerdyvaC
j3gICMawChj+RcZl4UR98JYO3yC22FeMAuXOBaOC3hFCh3D09W8aJbDTSdaO
qfJlqEC2VNB7qXXKefYW45dCz+Kxp+iaQkgO5LYRfDsMzdfN+0wo7eHl/ZkG
oeKQuYn/mvGskq3ceEXSzXwT/NHD/jv0GQ+LXis9r+sgtwoH6N7b79rFbaSX
JdNWebxfiSYF3oZhkupbNYWR5DnPlAlKJDN0HYZJyLWVBny6l8Avb6ubTDHZ
QpNc7SgEEaS0xK2tFdiTjvQpL7pQWiP4OQ5ttEVZOzO4Q5fpQjeqHtVGMo03
MAHjIyN9T949MczdJnx1rXr2PN9MbxS9d4oH7XclBfIKEN9lzCVB/jJ4pmSq
NmbU3pO1huVaDhbM89TPLPdSvhcz7iM4rOSJPoCAkPaheRqE7a7BKNWZ4Op6
1JBmL5/1WKed8R6oB8yGE7V7+rB3DskMUEgU68GYrebsM+OfWLKN8TD6/dwq
uW32g3hGjkVNP1jCVxhdmhJTV7q4HP06vzPl4sei8ehSJMK0FIfPPhyAciYs
uP6+h1wfx3RFx8zBfxjaix5Yv/vx6HtYwJeLlMu4YPtcYdcYwVL4g3lF+MLa
g0cUc/PzEm+32HlcA7I9NE1YZfQ6KFhasBMB8gNyMIUaDuPHOruct6reumur
35WIYQxwlJtb9SBQR/guJLlP6+3ZcSnQ5KvAb66Td+1U1fh1RFt264xnYe/b
eIEfJP43yALojbFaROVG/KSFkimmoOt/Xe6mbb/zOMHZFZjddp9N+2QESCaK
uukJwchrQ/Ms5d9gZ8vNDYAYFGTyJi0+02lrT+nFo7Ybycu473QhSm8c3HqO
rn/UeleWANrJ++RkltbMzlxooyhGWASHy2h6WoInLjypvcEP7CxNGHvlhH8Z
ypTGEf0V03aL0vymAQhr9ibpuPAwdpvK/+UnFinv1weerJlZ2bIfsKjHgKsi
BDdYJyqZzof5tqxMLl4hqIR3MGbILBlqYByNo9iDde0sGwwyYGXLaYr9IerN
BDUH2O3pWP3pB1wbvwAExEp3mCP2l/19sp34fQZJhCFSSnCAclb4Az7TuhDB
/AVcPRDaiFE8fH5DGUG8IRj2fofVYQHe5wXCZeqVHU8rii2ersUVjd4Mf2B9
ZIJ95ECciF17yScJVNC3Jn5SFCpiCXr9ZYY+UIFHEEah2goZlwlxo8uq1bpV
Nc9PM1kni6ftY0tlhusEQFRHC7rnp4R5HjBHzXq4XgGh/WzlqeUkbxKP+CDb
KvRyAhDqGHrxw1V+R4jzwOZXuIhxmjFg71NdBdYjPqqBb0ecisqapJ5AdUjT
5kAreCV7N4ANgXIiP+hAl0vrsHVZFq2DJUolunPOk0obgRmYRM3Wm7reO0Jj
w47BpIxkFjgt4KqLa9U2NppUK7aKKxC84Z+ZCdDejo9Yh7IdyS0d+1gbE1eW
Xryd/HZMcRF1OKlWltNvQvFgg4gCohLIunarroDcoCQucZMEBy9OMxjZ7QYt
0Bp6kJi2TYW+FzKUN7FG+Agb2KL6S5M6yYmmSpDYmf89LPGeHYR1DCb4TTzp
GHJX39v038efuJ9uyTfnET8g5daJV4thGkSj92yZXR7CwcOXRadJjlP7Znwl
Tq70RkwpuQJ/ZPh8N6TyswobQ1aX1XXJSf0J+a7BjaxIIzjXZjbL8WHWD94i
v4z+J+FUpFPLRk9vzt6DGQSLm1lGrAeJ4fYL/M+dJ6Rwbf5apHPRdTDUYf5n
RzCbxBzbRBmnKX55gvSw82t+bwcbBgztu2mHI8wfPp28NeUkX6D0/q4/ZEy+
V0ULuRUNqejxTnL2ClD7LAZoazvTCNiY29xcoUzBGss0Z/u0XRqftr1SY0Rm
Iy0hBClsFTzjLXCBfDMx5081pUqSulmj88ayVS9yB3/dDbAzMCLaFMM+Ef8m
XL4sZyWDLL+31MGDd8M0Kj7hmIGk6M9PRL84lP8UUA2jOrkQhXbEUkuOH5qL
C5i/frj/PT9tECtAED3LQexoaFkuofahQfxgoTepYQo3zMn4rPzlFE2TrFid
tLmhrOC9OPb7fbchWR8yqy+7FR/MxWnRzKZ9QYMmsLxZWClPqwTJ/mZYWaOB
ZacYlevKRwYOFQPzJg00vFCTILijNUeLyLGe6yqkBTKxLYgKvOjt42wPUVEK
JxZokVR7BW4fj0GoFlA7WtvcbG0+2jXNe8Ju/tmHrcRJZoCuvJ/y6A1cYGSG
gm2Fh+EHGiS2DpoLy1ubdumo4DBcehbVgneOriCVUc4+MwdXqZfg0C9MHBeD
QaiB99Rke+5dx7oSppChiSvmj/bZxgeF2Gs3uOR9PiJJRlTK6wm85WlOYMsi
mmxGfLNuATLwnDMCm1O11Td+wwZOX3Ub12Njaggw2xX5vbjfVOFGDZ3Cei57
QkqKUcABTSpRMSVuKie1O+rvfuo5T6WTXFOaOOIoXOb8fTcZ2KqMIk5F2Vp0
ONCRX7G1+mo+eJEOyUs0iwQQI5+fgmJQOIvV7uuXMA5nm6iyMNkuaNvfcsNn
AtLcSOrX+7U7sMuQk/E7f2MWG6J71sGTVEpatZlmL6fIscOZEl4dInYtMQgu
wY4bvVKbxQp064KYpgib/g47Ucqq3L+u+bYOolsm5X99+dPB9PukHrt7hhB2
3OXdSMvf2YSBBF4sl1cAMx4iparyiw8/1Ez4bEzmypwEvHd6/U2KFxVtsJio
AQ0UHqUAjv4dbc3ZtZ1yTHvwwDhi5Hc9pUR0KYFXx+G/tocDHeoQA2fxnz3F
X/hepCrkJt9e+FiptjTANEguxz604Qul/Kx1GODbtzK+xS8exUn9LPENfRlE
PUjYj1v8CQJJwAyFOiVkhaCEqgS9QNxBbHFeUqyyQwEqH/EGUfCC98cFXzIz
I+VWMChJuTWcoaf+0ReZp6arzX5kfJMFlZMohS+xCFBxSoOMudk2G/Gohmh4
oT/bUgibQVx1Jf/8r3NGy45CpIzPHYPNj0AdHRQvw1OkBPEg9mq3JfXe08Lf
B4nWbHCVk7bD0p37WmU3oJb5ubSNZkqAAy7g+41bNf+Yg7brrM1UH89VWL0y
xpsSgBek0cnvAPIkHXlcxEGLlALKtbf8fgmHGw/JDSDiYLxuhNxXVdg6JOFF
NJwvOzyNpugRneMBUG7cUYpst8Lxkgh8Vs1KuCDJ0lU+iqPpL+ZwXkSVbxnR
2B14ck26yMBIFKt3w0b/0qSaibRMzKfACRnenNjeDC7JNVd2JGGcfLcefTnQ
EjUCbSyCUE4CN0L1+BAzJ2v8hoWi+aK2vQhm13LC7esK/6hngumUAfIWcAox
679tMNqxby+hzzkf54Ct4T7kaFqipB8RKPUdQhl5oEot1Pr6E5FKVzK4htCh
nFdbXz6+ypsxWTeWCDeRAddLeFWEv4VrUrPANbk8JpbXzXVxP4M9XZtFn3Fm
NvgBTU7cYAlASubicJ030hq5Dx0BjCHrP21IsXYphzAyXUOcirsbcRrF++rT
aOyeJ7Emcq/fJRCjSYQu+i2JOCo+jLDSfN0ydQtY0Jm84AVlU+BAyX9OQ9E+
Sp+DoD/O6WqPR2oQkOU7osNLaXY6yPv3YpLkI0+VCSfoljpN+hLkq5GpE4Mw
JvG4+v1mtUuxlratBQr9bpX2lEkYZSZlu6yzY1nxIgkoTdzpJC5zslQA125M
roY4UTFMAuWMPiD+13FBdYc1tzpYTlLbltdXHIL6njNuWyStIsOFfpB2D0dN
BCPmfQBj6JV0/HD9ov9Q/IDJsuYIqOULTCclM0Pc1FzEBpiCFMbLZccLqKw/
dGnVgKCF1pZKMmYLPKLnVjNLZSWb9/Lcd2f0p2HBYApJzKgD/TeZaA8HrNxg
hHK5X7URvnPX2qHFwHA3+wE99OgTeLbStdW/pyJSyT1gZoar+SKQyLab+syi
88wcKXAeWLndcnaAOQsWEq/siwHiQ8Rx9Qb9quCSbo6dAHaidFpVE2OCm9nb
k97PsJsQi1rWSOXHrOifuxkE243ALitXA3z2tGMzUdAPQ7j3nCMxdfJtwnlc
k1S6DCM554eQhxeqP+Lw9Fbqe+17B/ymZp8mNanG5CzMsItsjji6Lwu2xQs1
GaBzD01xizTK3OJUPGr+fTQzk0kFCM0L3NkLzfnhA0KfhEYVxQqLlhKnOwMS
vpo9WJO6CzZtQJSq7vaEHeeZKW+GLFZM7CTyx2/YvGEULHfKWzrfEOA4T8UK
rD1nDXkfj+HqCVioLMB4JIulndtzj7kswP7xcdw8gWuvx8YHW1BjcU1i5db0
6JyfZ6yYgKuiKAtfsy1N3EVhshoiWDWbeJmrriRgNnznFM0DOWc1MPuXu+kC
stPFM85GYLENatvv/KYYnOx9MZH5Mz7Oi5liO+stK+e+TWoS4W39Hf1+jp6N
rNAyOZHfu3Nb6X1VqS2tOELdyPzvo/CxpsNwErmrMZV31KdwX+TBbfatWMlU
tJpO/OOLUQs+EmCatbJam4bgRym6keR1pfMyiODN5jQ3ATCyETXJdtI9kDuA
+2nwW/pP45yp7o6Nbc9BmPOcExsQKa1Xd/cf1WZYnO2pjPrTM3DPp41GS5XO
82mGRxKCaVjTValXboilL+k10j+dUlOqMrjaSlZ3cNFdQ6g/4RSvoNumtqad
900gxY+Onj8xLmcnqYobG7Kwlphz3yeZXFealmlL5zJLx2yTnWvl17rR+Ka/
c3OKKuw2QCVWdHmsjW7RcZbtEhLnK3TBMLW9RGjFYdV0RcwWtwmeutqc3l/I
AaYxP+wSDfkbpS5bkOSS3py4mR5Phc+Rn2ZuoShjy9SdNL087a93mY/amGjy
i18yj2LIlQvJWYbaf1oPpBuu3u2hS36YS0DYig7WjM1DM9HcYO75JOHgokEQ
Ktwbdl7a1lJAdka7t0F58NQrNlP+t8I+MyHUEdXj223N1+EJdTyfjTG/R71j
Q8rLK1O3GB0gG00z6LsyhPQUNrctma5qK4zetx0lERR4nP9MY3jeVrIlyskQ
rm8LKhIurdirqMyERxLXzwEXszXsM35jCrULUlV9L+IgupV5dxg7/42lMWns
ATrmfqAxTfi7pGwoniBo3VghrvG4ZzOfxl3fR6n+LrPbyzM21vifUJkAeneZ
fKtilqnAUSq6TTiGdJPNizgsWfBEU79V6u1H3plTJc9v3N9doFBYKJWI+v3m
7WNwAKW1JogtgXa5Icenlu5769N9W9d6Cnt0uJFYrSd7LnRcRHqurpGjIePJ
wP6cyiKvypxU/ij30X+IyrzBI3GJg/axB+ebezAvvIR1GBd+CP7/B6Ji6b3s
3dkYLP9IXnLcBSlloZeHHQwTLfzJ58uspC7m7tax+nJgGvgcMVpswEBwmoz2
BPPLUSLZxEXicZB+5Y33CPrRiaTwOwYBqv/KjbbrxoemxmeZr2xDgOUABIj3
hhhr0CX03tTVGkIiTfGmU/nOKzlOBCLUDT25j293kFnZC71Syvhw5/YzgXKE
L3leJxmm7ViQ4S4rM4LvZolmDNQsVQI5BbhqgYQ2lcgJ4MCucNNgfybEjbXg
RbbBUynjZ3IfQf8VzbUgEvyK6HNoizhguCRAt1zzbYt82l4eLwcFUmYqf/1/
xvJBafTbjLqWqG9iyze6oFyvhobWctBPifPmOTzOs+RKd3GVmxkSaDwfogl7
YlXd2XjU6jG8N9x4n7r4VUmJfAAlWzoVXq3YtB31i5lHeBWeaS/fACeLUQtZ
zhmEyYrLu6dSBXsRBOwcKpwSIl6KH3hAErVymdxEloOOWynz4VSlVapfj+yF
p3vTcidqph+u7WUcZu5c3AsWUUFRP7h2ATa7E/VvXTqcfNui+x73R/y0aPSj
Rtimo7wD024e70HoQGGiGt6DN8IIAdbiIEF1OcOEHieIQnGazAwkv0ORKMcz
m46vcCFAR+n8l74RutUGfo1YJ2Q6yoVzj0Sjhiv1vQ252+BB/ijm4whcfEGs
Iok9hTakecFFcmQIQqozyD6Bxh57E2nFTsyfQKEX9L9pU/J/IrYu+PSrVT0P
iLGtbZfLyUjUxtyM0r2eMrPfvWXS3YI+xVu3xFPsP4CwJQujZJbGPMWnVJ6n
ua2U8iidALarDp8AC3gM6IXzaa4A5wSNQRKDoBJCMSapkX/S534of580xP5y
plmpWVnQBwKTrEvAJ0o9lZlQQX+k3ckWHv3Y8kaFf3LCGQ8vGf7IhR9/H6XB
EpP4LynbbAtgHllnsfyPfMJTes2FErZPZ2+HYBBlGV1KL61vZ4SuFtErz0rc
j94kXqAQpMWud2TQ1YYnAd5F2H/00tqvOykIfy/k68waTlD2Cm5Q4utvIj3u
8UWQQrb8Sq94q68RCe+GBo1u1QAoC7hEf2/FGriaoTdnPyvF9Yyl0Vak8dES
/9LrOn6TI/9wSacsrkLNFFxLYkFiz+q8Bat+FAxx01TfMSYysK9uC3fQA8Jr
52HANnCqoYsN+OntvBPSYLUHmwNl5xjmDKVV6KrsDkm8XSr0co8LIudtRKWb
zf+5xaH8IGHE2Yq9r1pFHDO1SBT2qN9ITjSY8s9xJrAdCGqYxQfSUWq+Gr2X
aKKYGiciy9Ve7gJ4jP0qYf0BYLZefwE2rydxKJvRJkzWuyGasyqo/rA+vHYw
pAWVW0TKDzvYcZn0YFjrhot7Bnf+je3pwFh6TpUiKMqqDEB4hwOVlRvx3sOA
YF+4QsVb85UyVpKvFszKMYU2Y3VjEN+rSFBJT+a/5H+i5VDBnmFLG1yIRW4K
rffVo465jizPQA57vSsIhyiwLmTAF75x2naEwf3VocIwBa0kRnSdHeBAh+q+
ODzrj9fbt0PrV5qmE5Pae7xYLcHec9lF0tHHv/DeNNCsLHT/JQqBFZLQZKFc
YAZqBB+4dPuJPegnssznGS2tIoz2cV0zovsmowVIjZwJMzMNP564J1O4tf2X
MtTyCqHiUMP5F42XFUCbb21cnaMr84OCvcaNS6t1sbfdhjpdVYeF8ASkd8pd
UKevhlcOL45JKVPs3L/eYilRfgbVR/1zqCMpxoNuYECcnz7Fwl3nRzmAzdC7
nPpPfmDiw/4XrgOb57xGqNW1wD+ZbAsN4AmdLIErW0rmiNMk1moShsDuGdM5
9x411XPoyoyTUTn53x9/Lncnz7FrQWgjfM/lSbLvQZ4GF+reLuYsZCkkB6UE
6MyYo6Okh0QX9SWWbPd3ktfMfatOfhFATkPuMX+TiqqvgRVpL2824S6le+dz
qQxOD5tyOKzrSNyXGT0EKqgQ7h2oyYoTZUGOqbmEPdDRIrYC34Sg4mu30U4T
WgpeGc23xZV+JJ3SDkn/BBLgXjG4CMBIxa0k6I2JYtvOlepYaGn+CfJGX8rL
v84TTZCO9Owx+KRvp/AYxz7NHGWK7+Dz0DTUpqjCD2ZW8os+uQozzH1Mg6bs
NGTy3coLL6/2Aq4JDGxv9Fiw2nigBXgd3SggzDM53rmPnhdX/445zV8wwTeS
/HTiaD7TXQzuSt6ar7pAU7keKedV5Ftj+KqQ9yK8N+OPavD3lQvsu1v6us1J
ahhARjV9zI96av6UOwRsNh9w06RL3J1qCWsDvCGhmpePzlvE64k0nvMvHDZZ
lpg4N/2MdYJPBdS93Mn3PEtabX+yUjhCV3xMmzLxHt9FCz/6BCyZKWe+NlU1
fyBv81tHFWsZuv2IOEJz8ryGT0EKLykhXGk6xpTCGQ411k6YX6XApk7iodsd
NLQ9sqf8L8vw8qkp6RlazGe6WULX2zBFvN56ctZ4F1qoF4/JcHHkbDxdVHKG
8SXyeiCBc2JAWiUXk4W/HW+VenTqbRrXIv2wYKp+yQAbtwPMbNjs1gZp/TZG
suFbagYzoga/5IpA/rFUgYBrzSjHrYv8WTkvU+ilTqLkfoAEyLQSCphGzhUV
6iObJbnFHAuj6h1Hy75tIsV9f2WJx7TE1DFETpw+67yEH9QojnNc6FbB6foi
YbPJlIlnJ/wi1+lgr3B4n2ryX4wkhhobk1OjuROffxQGy2IhJpUQcCa2k8WK
oKN+OBhw7Lm6mCBGR9qOhA/LhTBxCWz8gQWg6Op1wXA+XQ2lV9LiGdNo1+CU
8gInP5/DJIpqXIq6ltjZexsAX+jaQ5hfokynSH+Tn5/3G/pBsVdbw6YEWg4u
0VjavDVtioMJQzG8D0Gn1n9xu27EEdy6aXQRLprfQpQBpNkBkNJbplOmc6Y+
sjSrrDhcwOFc2XAX4079GXqp4znUCqjd9q0kBhGHKNkhPF40qfRgeC3TZdy4
9S24jCAcnx/vi2/3qdYEMyUCS/vk4fh/MQHJmgg6yhGsdD5DE8rWNosabdML
WYpGNmXdfh8p3R+VN/iwvowDMk58+yM9Cf8+6CDEAMZF86BqpxSeImJ0IPfp
vo+c/plk1eKXIqO3SCmU3EekhUceXwD9cPxiGjRx/r0rdtoj83LNrfbx+mIk
/eomX/hqQk7mZTx7PdzNi3YNslJCIYJlemKKl0mCR3u+m0TsWbvYeVR9CTTc
BhGLgJannQW6qMwTPVysqVarexjN8arW5L5mvtqU2jwSt/FUncY1a4Evd+Yq
tcOVPOYKJEf9R2OEOulMjoDRVIgI1t7Z+xaYSvIWrng3miVML0eKIbyUCKIO
AInG1ZAhGY/sXD7fK4f03F1VRCX+sOdMcQv+DBrm/TZRBADByXTzIcD8cR9R
RuEEhZEKQXcXV7ny0wzdxROwK1s1oQ3seUjbUPF6CkIRnXIPvNnBjY7TsuCE
9ovxrp8jtzWQZqavV1iJkF41a/R9gWh0Ki5c0nYoGmPrU6wCC0mIBQqW7oYL
C4QwPHVxB5wc56+EFvR6Eszf2LCrLxC42Ymd6bNSyIN1n11YSj/1+gB1gidC
2+OfL2TXKBQOu7Wf/4B+h0MjGJyaycEk5DiVHjU4K8Kkm4NqiKH5rbJ8V7LZ
idjWVAy18IKEv+jBbFqiwFJmM2WjF04fijuQoeq4rS4tTR3Mc5ndA/793XkG
X9Tj0NJkHn9hSG81Z2Y5/7y1L6d8H0/TiLh2louISOh7IhHyHql6Mx/gtEoS
r9o4XkJJRKL4rCC57lxVFOGXIULT2xKcESkhDv5Q+n0ISNC15abM3IKMKFPU
7i89WeIlwLb0QDudpxjg/WolFtAxbAKiiVbAJkd4JVwxNS7WCkDXqrIW7kdX
MmgI94WbA/cVcfdjjyvg8+j97G8yKEKP4xqH4hZ+Tc/23uG3CyJ6QqhJX/Im
XHgr43XwCn1h/qEnQPbJtxbcBqIwlofZI3uSTWML4/zFoVSbkbh9MhTmmqtN
GLgyAuMkIS2tSJeXCTMSV4mnWwpxdu7e/CphOYdUtGzHjVTddrrkU6CVDl1s
bKhnZh7Rd26A3rQJ982haoNqY+jOqGUa0PIWK+0EKqNVzEbU/VPz6yO6LUsH
ZwmjK1rWfyaMSWGw0x9SmMj2llE2BGl86itBAtoGuNJQQwm70sRl0GLsD8DF
fQVF+HdwpjSEiGbfHqhwVQc1EkMrSu2S82cWC60KJatZUXvD1b2vrjWtpOcX
MZa5eTI0u9PJOiYFtN+CFKbsEjSIgkRPByIgndmdWs91+cHwsvF54w1KLNvT
xV5ia3i5tYMVsymIvXzO37A/ivt0lyba34BV1Di4+/J4WWA8Qo2AuKs5+fFn
YhP/7DLkf+/80hh3cJbO+KZQB4DpjzFPks1B//sOuLCbvP3cCAUb62uLJax4
CF3HQmv16qqYrBdKvIzInUVvnwmIE6R/41V7fJFgvZbJuEDQimoyGXuWpLVy
A5To19IiuvA/TsNPGRGqilFI1S44cDdUCeZoskUHMRpU2ZbuIVs2dUbDU1VY
hNGAxDN83wcL6PZcI7rpVEvBesBs+KUa5y6fHVvHgyP4Mie+ep0KRWCADN4O
h3aQa2kHt4Owbin4niuAiyhD2U5vu4Pye7lDwWj9BRr651Yj8wuyThCpa0pr
lVrF/zjHnfIrmru/2KI8Lk372tOywis+shtb9Pf0dKhVFmAA5Bczu0T9TitM
avs4bHwWkOMD9hQF2RpCXHU2qg1C8nBhqgGQTPLMOfYmkPHUtvBygOtnV2bV
KTrYgsGuNMPhToXXPKFQvcMq81cWOlxXUqFb8det2NYXwu9A/N961Z+ytxa1
s83uuioFGknVSqwb7+k5bWIUSdD7mqD/dCntDplPLvFVhAzGZn5aCqy0mEFX
8P3ZV3Z79XvI0mRroiRl9AcFv9VHs3zmIbHewkpVO30SS4QeM3Y1sGsND2IA
NLVKHoTvBrTq0kgpRH8Njf4Yo+qu2BaRP9eLSVz/0qhrVsV4+VWmuvaEb3Vr
RXhwyqvsxVpLI2JIrroNHrzBBV2AbbBWgFBPGBy3Ma8ROOQ+Pr3BA0jdGA3L
D8oIsbHzf+IszOOOiLp9C5Y0bnFX5iwYXkMd58DNIZ1gPVrnpd3ZH7Ofkz2u
h73Mh/8wG1zmPx3cIC4L9OXb2wZ3OKb+57N1MftrHJPCJ11+KlPwV/koyEba
Qx7t0X5LF0fxgyp35GDO7FKRMQqLfKNZvD4YgiRU83WezjWMwkt2FltAKaz6
fBhxMzxxbdO2Ro9hEh1BBYXR2VZI7WKmmm+gx7m5dFQNC4BswoTZruDh8K2d
rrxzzWHQoMFGcPAyby+37OUqqwp9B6SYYTZZCGCLfyy6FgjURR8jmton3uju
pU2i2/NYtGvfVJdYrCiItHJXjAM3oJhpCTxY7LhDQToll1dG8kBGyKZOCNMj
d2WdSGKONmij+W+PLzEMZMjCK9V/5+qkAIDC8rK6blRYmEUDT+/MI+sepNFA
b6rsDVm3xwt5xAI8MjowoSUlMca7pfpTeQP9XM3x5cVFJzzeojdlVXWRrs2H
AtjXinyboi5s4sPrOflg0MN4U4O//FGGfUJe1VyootAE1QST8YDk268BTlzX
+zVme1cgNdXUsT9xag3+LiMlhbZLuo2WhxFaDTv+c2w9Xz3yYDm3w9WpFEA8
uxYGfdWosWm5mWlJMvc5cc4ZGYq2Pob+q+N6x7ctQa0zlQe7CuDX0woDnVIl
ebpJKCavVZr1F8QaXSyH7w60/iNgjhB8iEX3QBIXTS7Wxo/oohXg7i7IK71V
U7xqPFWpJ5HplkM7actNfDo18AJMCdm/ViGnLWZfEolqCXuWyvC7L749oKPV
ff5ph3SQsFv75lR+1KPXAD6aQ5caiC04PVa2ZA77vf36eo+LS/hxfeRF4K4b
a+nD4VGX4EBk9uVY2Ehpw6suMeEx1G2q1NC5M3bLUscmQQBepVhh3LzHGbz0
T40hAC7OZMqgn5v6kUdvVOGIONwadhDyiYoNnAQMjZvwAysuxFakpuAcCHtK
bCfflWDQ9cYbNKtq0BMOTwx9PWn+u4DEhaC32UAMtFid3U72/iVGL88Q2pzB
l8f1oIAw54hAX1y08IKlT6EFD6kAt0ZQlC6tDzppb24gO34R0kWESiiOUhMG
uPF6EITfalrDEyTqUKW6x1V6gBtb/1l+5E+sxYHnhVLoYHnlXObNM/HmXAPJ
ql8wk9mVGnJx9dpVddPaz9TFVKTfrphXGHg0nf3y57F1ShQDAH9eUXVsti9/
wm00nmSiwtwIABErvDCNVvoxtCulrnj3ahcqcyzfcRYCXORHTov7VtEaLlw+
p3XD718+euGRBHNIkVXsRJOl/ULZddeAZpKEVYTLjc9p8X4vJh+r1LgLWFkZ
tVzK3RFEFEqxuCev2zVUwSNVQcduNgLR4J/aJzAqd5Er9CAw3tdfz+aNsb0+
n7o1v7YFGdMSf0kjyy8G03zYV0ESuHcmhLKrGaP7jsk2Bgr6Y5liFe99XW7r
KofWHMaBFUWTK11SUZXq047p9HEMC3FFeYhIfdfBlrITdarP6Fsan1IhWp1w
Ek4WmPgymTVYnBec/A+jYX9MdWFxXhMtgPJrfrZ6qUwyicADitf2GlxXXNPX
tg1BHwl+h+fJvtkFA5i4ea6qKGZ7pPI8vKRjumktbT64m0Ng6y/74ybTxHW7
K+cU2wnOfBigoAn4o9XEPnsOvcpQzL0q3nZPY0Zj77ogUHrFo9BFTXLroFl0
0nsfALHF/WPqos8jhkT+G83AYShQM2JJ+GLtqEKVmrGKEygOwz421TmSvKEz
ws7kn8I3vIxZZWi8wTb8ztGlGrESMmm9guZCEN9vISscri45VUTOnc9ilKsB
Fz5vi1t9i57takF3SYlSny6D+DypNsjNdxr300E7F1qVw15CEprvqLsAAPfv
920yjTGTfC/wFhSZbFosWwzKDirBftODVC1BHFZw2ztm9Uu5SMPoiwtgG2C1
6qD3q1zoZsMkAZqrHlFGzIWMDGPon8eIQm0Ab5i3gt20c4Hvcj0EdGvZJ6Tj
suWufLSYG5UwEl5wRb+6aQrIsBUF4DaSrvsYB4OFPkvJdjiyeOwsMm8LG/tL
nr8+FZp6fKC6b7aclFDMhAjQMWfksezNKR7kwAK1vNKDpFVOv2+qqGRkAFUh
EwyqYZEvgiW3a0W19VkGhQtJHUHYIwwE2/SsWCgWbr/hWS94lAijg67AHTu9
jKAwRqBjwqRDJbWnWWKDtavUAFbr2FCthTodqWw4raosXeJT4mH4FfUe0jz9
mSaCYbmZfRgCXfmKBTAj5LyWPACNVyqOLF+RmGO2W2UdYHUODgzVAxY6Ooxp
zcYg3JTfrrgiXQFiRQbM5u25jYY9AaQZn5TeaFt44WpiGpubU4FB76MVa1Hd
3XA3+cj54FfzBaIfL50xGq/nSFGcVq+mUXZUE9MxfdPS8Qzm0jgrP2lq/cov
JfGOzvGN088oDeRghgZeb7dRWNJeOmiarcUuxN3wpfHTOkXTbq7x78qEuiRi
MdDTr+7GwkL4DvBhWxj+qrBuTv+hBJmAdWUGNOkgMKDiNKHSPjcqEF9w3DGu
fz7ujR8F7xIShCg6+1wOFeNVKuJ/AMXl1BOL+qXMZhTnGiKzS6oePY9a37fl
g42Mdrf47yA2JrocqvoPq8XdYptVcejggC7EC51Vus9fQvB8C/YJlYXxAIfh
VhOPHEOAdAP3vb730E78IxJBURDNnJ+tqiD2kQhoSW40eQw06AhUMyyCrp+a
ZZY5zK2KQAE9zbomUqYjufmIXgu8irrYHNmOCWjQYH5wGrLV30iCpCgQf5PG
7Mgo/ghXxLx5c6ViAngYVgG5/54gaFgIYaWE4AUCja+gYx1qILYpIpl7umCm
aqBfUF7BvFRI2iqCtvFw0bcVM6ECSofpTnJl/hs/IvDGvReyFuJCbrTruBdl
xYT+0Ajj7bkizY1oyEwgVajFbHZLYOFRcgyfig6uyP5turJdakUN9I22suEy
E585jxMV4JnQb003nAzYF4IQKl3LsBJwXQgrmJ0ipkFFpKdIJ16ZC/aXhWHG
WNyGG6dStYB5g7cQlEhi6bz1XzXQyqisZHnfrPadnN4BgBWmgD0TRnPP0oDK
eGIrsgmQsYRNyOBDkagobos97SZYjdItMlhzrqfzznbc9Uw2k5v6Rlc7+8io
2tZ+T5YFOA/jt88bgYPjYH3LyJJpzriPvuMKpr1XdMLi3FuMMtC2nDQJdg3P
w0MdNaE0j3BbIjUSwSvk05vnTTNNgChda7P2RGNkjZb9YIBx6OPPbto7KdkL
2VYzk1wZEff4lkmDriC+jgOgEbeCilt/Au/J546DLbUH4oghl5balHKc+p+s
WhT8N6fsUBahXxzi4AWOOuFeTsKwZ7DruQ11vJeGbjt9635zecH2Flo+7Fdt
kTqJPOoWQncbqwagM9EEKSWwkc0zo6WqwbqU6k4AjbAkFZ3/NVz+w4zaRhiu
2OHwRpytOHeX0S75TSSOO1TJ/xrkgyyz5HCc0yEVz3WAW6Ou0DfzgkR8PIHA
cEc7ynbN/nPWm64H8q3WMNI9IbloBUVMtMulzETT9ppjk2OgjtUSzQiTVYhh
kZeRry4gDpDvYCGT61oWWhuuEM1iKeb+gS6iUOtwiiqlD+fcFsMMxn/jtOqA
9b1ZpXHISiey9piskrDtGWoNvdCcR/CFwRSLuMuTJYae1TkVy+P46EzfVWYA
ZP+56ojrllhyA1U/GkPCPtvaW6GkeuZPwJTVZ5OFAOeN6WIOWRYwnsPYhuGu
UwM6F4BELRvIToi9m4ynFBKjpC3rSW7xoJwdVb0TyF9UlUHp4/nadrZDjPS3
zT4MV6JjsNa/ekhgo4n/MZPUNbIUGmIdbKoCjw/i/+of6ap25HdEgQeqwu4w
b2cLQeeuow7fKxr1M+KKLUGKQka7M8+W8Td4rLJ2JDQ3UOvjMBvtvz18wAYQ
YGRUij2a2aNTro3o7inQhurb87DETavwz9PXMLOBz8aJkqNfY5sBs4wXe7/W
ZYuRfrRU6rK3j004PLXjNDJkc1LGS/A40Dhg7eaLE7NsPsCBqlT53ruFJXrQ
BURRt6R1x3MMFhzgZfIKhGA3ydJeGlvDPxo405+huWpNaaD6jW5Gr7lAWKBC
P1HKcp24diRoJ/0cbmNhd9diBqTRTkelDXapFBfwTGRYFcfNQpH/UTG+D2Gn
NIPBc8xxUw7mNBYhIt+7oEwIqGp1c7fzW+XPaKTF03JLzf9xg090jrD9jiPf
2iWAWWKfxFIBBkJBLNepct2EWb3sImA/Ia8olLEydSUgtXR9emdHrT/eIaL+
eH1oXvhhZQCHuYokL7k2SjRVW1Xcz+GhMeTOJ3Yh23r1p51iWG3+ZyY33ATB
OFguyo5AvSxU4lfstjnGTg3hq0wukC0hK+S+JWC80SWnj/vUIbr+w9sx38xJ
Ff5MLu5SMJKUG+6YEoMQxLsv8fvsliMG+disFqlCdhz1SNTp2FtDc/AFgsE7
rYc8+z26e1rqGZ4ZBSfqrsfcnYdrRutdukET7GDOplcPRrlr3hBtg/fBJ50g
8nVPEM7qODg3/aLbqyNDg21Ykk4hmlmbEp0SOv1uiuPdADxVS9i51aAdma9r
SaCB5qvM+I4+h3tGrqBAutgUygUMfTgY1Oi1Gx7sTvvvIUfkHmrZPDUPUUIl
4Uqpz1Rl1rQE47ymcespqxKrTsZmhHFmizxDAaMo3NcnJ7Bm5sEKcLAYnRGX
syGkgpqWwejuz73KnTU0M6baWKarcVC9PhOJeoTCR4KeGnW5Dnfzcu6n9wW1
+PmjaVCQi0qZG+k8AbygWGs34Vgb9X2EcqjYsUdGg4IqX2ZJp7RQcA19h15n
uZskeB0Kd6esNpFdl82evO591MJ6UkyYfBnVzD4PyJQMRNc5+xji6rHce+N9
Jqswt4MTDLO1uw/tMnsg5gmUMEdXe7AmVegcUS9SaEpxNi7Ci8cEOkedQKWz
ldjDSc68vRHKaSb+cLm4zabS1KlrLrZleF8OsqlKSIJ2Pru9auaYvfeTdwxC
wm0X0PPyTV56DYun60Owiqjn3uejonSj9YwXiM1yqmtQrgyT1p+6WCpM82AT
leopLHyQDujxbTPpuixWcH3AFaV2ZKw4FQgdanKKW5lIZNeaP6GHbHQ7zfcI
b3krQjgLfuLLwLivt/NrAKxtpVxRh6HbaY8v4D4Yj/nyoPovpa24/7W8vBvJ
HkGOsvn1VtwMPh2j7YrEsZfZp7Fb3Xhx3v07LCk60Q4SNLsk7Z4yeNGrR/p5
zguZdbdxMFzbXOw61/MINwwSyECV7/C70zwSEuENjVBV69kKHKVHN9LdLwBk
UOXNlF+xwgWRV6zJ0P8SduaQusYQFwjvDO9tb5/Zh7uZ8HaBbscHf2wY4P9C
ExB77Fnx2LDrCsZbOymBQOng+/D3w/wQXq4WLBuF6EmZ/I5NuvDVmOevbNrf
QDDdr+CDM8XJWgwQ0YJPcmWkRO34bVFDUDuucV+jxAHkVbmM5DSotu8J2cCg
+ERVv1HwQN6hbE0pN3ySCgy2HaLehPFnZ5vu8iM3sDc0d+GHHvnmEAqvwB2Y
HjenmJu5MtwAXjrFt8P48IdkDGA9RF/JbyDa8C3IIewo3gLIIP1f649zf6BX
RqVTIfkbET2S2GWtprz+wPTRFIV0YOG7W+FulVJWM4nnh2chxVxa5LikkSsu
ZioS71iAGmylh7pHJvoYAWjtrHcpY7OZuy8p8S1lMQ6fKHRCRtY6PDrP2HnI
7BYjYjBNgolUxii7DkIf2yYU3pKip4SGSWvqLC96B/1wSDObEKnVJE/pHspB
LyhN/Zm2HP0s0d/fTUZ7CiIQt2XJOCX3cuS1DdqxrV7IqhEJEHCMzRFkWReX
Klp0f10Im9QJsPyQxtk/kRR4wcGWNtWq4SVNwqSTyXsqPKmJwMUKQcOH/qCy
jMVq4i5TW/ifPvdkxFf1bbUgGq1SxkXZd34Q/3bXwBA5xSdmttvYFiIxPUvb
d4yNtv/NygUtht4tyhgxZNzeZaokKI+QHAdwJdixtzk1HNYYYKGR6cIU+E2E
glVe+Txk+2Zb7tQfeDiiK76vKMtopWIEO/o8LO8N9HCcNErys8KE/P38OZXi
0kYemZPX/0HQtvjS4gXx3ldk+Sga6wE2tXX32+bx7HVXD4M1UmpU8UTowzLo
MxgdSeKDU+IevADGm8eWhKQgneyC6HvwJqjvGSYZs1cB/WuRRalIX3h/2sJI
dmkA5nGtEmdJtIsgQxlV+tnxnyD0aupuQIA+eFQLDNsTPVNbHx1X1XRGuGQk
ZzgjiTOcRadLcUqCGXOHzdiKGaBFbZC8uiU7PVtDvE+30djEZ0F4sj8Y8/Ky
mqThHLofpMxiQ9nY//PDL0MSOcfPE/qwX9PKQ2Su415nZkXCUdZuYwl8Ib85
noBxwm7O4PD+encue+fToaIWeyo+rKU94bB/Blb4joOhtHsickcjI7CUYLJG
E4vF+FXh/ZdSHUd3FOtJZigpvh1q3T+l5XWCyclLrjKoPlcXC8TD0SNkKrkV
RMLRzQYhSwrcnHGNNus8+ChHr1n0j+CU8XOdTAff954EniuRl9DNvcxpKL/n
yzFBwplJKv9T3n2UV47wGYXvih15IwbNIfmcJkJtuSkLAwNiFIx21x8CDelg
/OIOP2UqSZ+rL7Wd6MVNo2SqJf5cCzcgZKJwXvsFxKdDxuSHllJ9hjCZFr1l
aoIdBuI6Io2s/PuH6H9K0DUGGX+z1YEYxVaoLSRzO0hK2Qnz3sg1vBATvpVs
vHS0B8JB1/zXXSZ8ET0efVBvOzPSs8RYWZYWKmA/Bj40QUobP52lhrQGfz9o
AD0AsYA+uLlXuWNc3iRhx76iMnRUa3hGlMnp1kVAWcf2Ez2wIxuBrAAL6+OQ
GKwP7hRJgLf26hptsG/CeNQg2nvWHjnczyVpz8MGEic1tFx1fliU+OBwl2WT
awQhkkMUuKEPIO7mBdwDFRkL5o6MEXX4JKLo+tK7s3SwnIBv+yodl0U+gl6d
+LwrofxcygBGQnINwbcOZY3j1v+2UsrIbSYuHNLe+zeC0XBcfceADQ1KGh7y
IG2hVRygl+yMSXzJrLQtKQzbqqUAIAfZ/h+JhNts9aAKDmXZ+5MZp8drkycW
rC8lnj94JaIxFMv6nrVh3fWzjArMtOVHXdh6TdkehvFIsLDFPAD17j4f+TO0
l1H9IQRjV+2EShdIxhdk80JxJEC7OW97l31NY1Dezt2lB2lYZ39ksSr1zAej
Z+B5uAhbHeOqMSTqG4WeLY8YbwrKSbV8HnsG7hreePSmFh0YjS1R/HGvlK8m
KrSoDbRQnlISRtERHJK14FbmMXxCf6xDSyeLnwxIq7fzuwCN2y4Of1NwLy75
IqntTIbBAjELQzbnTIV//Y8XmgItnF40zCi9VuBkrx7Z0HczO7j2WTPMGvVP
vMj53cc716XLnzxznidDmpUTKpnXUFiGEAXgdsMQ54YMymAwEnDkcER8UBH8
aLqaH6xa0rBTYgGyGrMQRx2OW5/gRY7H3fMiy5S6fIzAOBSkQeQReVvgRT93
JIDi4ZG1mIDGUUc7WjAWKrhV2pQgkwEbeBNSFjuokuVRn80FRco54HML1MIx
gf9UxmfExE2JJZBMBqyeuvWeGb4lQBFo32t17AYoreDwnM5mfBp95b3JRZ8l
jq4gUaH5fOOZjiB6fO9Ou0wyqCcesoNRvoA3oPwdNd0szB3mM6x2N3jdBtcu
SaPmJLWiqc25tsrCw+BtCt8XdVZvSfXqkB2P++yQVhXkzOW7Nntu2Md3tI4J
y+4SqgGkdIP+IVCHBoF51zt8sXEGC156bFTlZI+cowFAhkWe7Zu/wnA4O+0L
ELHfySHg5uw3QlDjQkaPfso2SewGiscVurouv3k7dqUgAx1ksxFvGRs30Zv1
NszuXrao8i1IMuna0M+/jESxnEaoUu3Mi/YnVKC8yV8jCOt3Kc9B6oiC3KVN
dk1ePESGBQArKrgfUuCzsamAhUTi6P6WY4ugt72MIvvl0TlmiPorj+Ym2qvQ
XUYadZqofZIYaMqN+gq6zTeC+HC+189I2UCv2qcmyV/jwxtAcAXypT4FPTbg
sM9CUGJ265jxXsqCRsRvuyifEsQBag+3f9OlKMfmqLdMtj0Hwt0Vf0z8+MXI
gKknfTKPJtqk592tQRRfwgkYJnVLT8rJ5MpMbUoe/SGOBc8rPmXnnQVIU2r2
ACxyatiT+yVCgDZ2ygkcGeIlKZV3zuIpX30Uk/5MYVgZY4jmTHgOH9Pv+j1m
2lCjnnRJlbyoXxLtK1VHffwxJWwLTvGJxByo1/aDqrggciT5+MpNAzbqUW0C
H1Ud2h/nNA3b2SbVxDNbkcUs8WaSrll/CxxqOMh+ddH6tw+vB8xs/Y8yk3lG
6kFlgzjUCk5TgTB7a3ISH+YoIlWVi9ilJMtZsQke4CjZjQZKm3E4iJHptdQC
c7lv6Mo3pY5Swro9wAY5EReWEoEPDferk4aM8YZkY9X7UGGriW62Xk4VDgwl
wFkZxSWFvEtfT7g1JW8FYaCekUeZPFsAEgVdRFLjYRG2Urx8NeC9wTusY7Z1
4X5bkSi4ol0nonwmMmqSXzG60qnGXE1Cx7gZyTq5LDrqORxuxRagpoz4CC0D
DnfTixpvMkQ/Pi7Pn/2w4eY1wWn09NOJGSWFJbDPa25CUWE/Ltv2kqne1jM5
N6z40N0sYh0lPAnJhDDi6Xymu9TSvhuNUGANcUhRVdvdwuBzy7qB6wDocWGb
xx2wvVu+sHOH/KMIkS1mcZ18J1kIU4WVzkz6Z0qY+D2T+r/9WXkm/iopbGnp
d+RYmiUg0nAmpgYhVaktiJdYHpueaVjqAtBtj5eVVtrKRVvhyZAZQvpTVBWd
AYG2CAly9QqQdju1H4aVCjkLGEmuR3aaW2/TYUbwye84KZwHX5yoVQhflVmW
CERLk1kiiB3K0JyGjLAzRX9I/0OpIu2CvhsZiKIB1wwU0K8sZJYU9Z3n/2h1
E6DGyNkvcliIJjpl06yfFq0LNj6m3NxinAnjkPDwVyghUyMxs87GZo7KqNxK
qquNvh5S2fgnYu+X2t3GfWLKgMI3Gy72aOc4AVM2wyC8NNU+OXXW6xtUBmhb
Eqvnax+vpT/SoEKRDJrpt7lqv9ExxnkpAG3jC9LXaSk3DQg/vjiRbJ4FcjMk
KTUH67/Y2pcbFcNeRJh4jtKoFfXbbmPT+rzcBXEerP3JaG5CJkmRBRfyXo5n
AvysHBA6sPSjKaJvHqeyDNqS8IrwtiayhswswvKps5rfcaFAp+6++n/K49mI
d5gWpaD43+Df9fauX7GWQST7JF0bBD+tG6YysADGxgmNJA/iyK0qPVxSiAcz
U3Q8unuK68GoH/TmOpeIzRLJKXHHm2kprO4VbuAGW/DA9n4eMFN+zPLj7oYd
o3aLnxGnv8I2kbzTlTivsoOonSKf0i6XFeJke1DYexmvfasYMHx4HHLkubeB
78UHodDVzTss2yEOH0cMCoI4D7WzgsuyPm9k8SIT/t4LqC/gV+w1UUoQPyE0
rcyXR3JccPDayNpFl//rsVmvWQHJalKQlNdgIa/LuNtxpAqhVmmZkE8bqvex
oBj2qTq8ftd0h4VH1z/yQGFbTzTiz/FWa46mRzXGJBW7XgKQlIwmXiqVY0Db
TdnEALgQ0ji8t5MoDovZtaDvsRwkP2Et3s5vhBP/1hHXEx21W/2r/z/do+0o
xtF54R6RxXct1e+oRiQJ+z+BMJAVwEeg+ulPuHMMvIH/AT+HVaZDq1zUztWg
rZ4YqcFOmocCt8yLtxvpRrIljssYjEFMHRgWYpeB56elQdjtrHYy1JNCzE4i
fTV+ZZQtgldMQLgquC6kAF/tzPcoX1ys63N+o9mq4R3B/0E3BlS2QSfkLbeT
M3+RukeSrfYA7rci1wum6aIrrodmyXgDF4pOvl9MfGfLkJAUhFxYhayLMKf1
mLG3iF+5l5mSR4Ka/bg/u9s2I2B07bXOcDNezwQKQiclH++yIWLL8fQOFPpx
jeBEn25P6xh18jYl0F0rGZDegBafnTZLIepc3+YPVsIYU6nR/4oEQ/RgGyO+
HH2O/WKdljZ74wY+9D3tFo80Enty4tjef9CMyv93YKFKEgguhktSO+69CHG3
5XP0w2zv5s+DFViE1Nr1C6Xbl/Qe8ZJMs1YvzT5dbaOF/i/snldgqnp5OlDu
9nfo7mSAEErzITtE8H9oTCgFR0w0R8leLFO6JXZj9MbR/1ULHEuPK31dlX61
5czoFx7ekbkE4j6sMt00Honjq9bS6jn2PMqsx9nEIILSPCg8wZYTvoqtJK3p
wx0ZHm4mkigRwNmnidpuDmD03WDuONI+31+lgyCUcL8fWPr4X66PuQRYtpkY
+ta8Niz+yBEm5pCgJE+K6DclNp6Y4954cEGxhanwD2XSeG54mX+QA2YzZ9G0
zSXiTVkE7iPT+2n2yLIgTsuStajg5aFbUrBtwoUCW+kIJsNS9mxLbncnoOf8
lGo+2TRvzC0++3dfSpwOdAxvFMZpI3YphsyjcMV6RTK/lwGTawuXumTM3jTZ
HzFKfLQCXle0/d8PRMPYEWNpR1a4HnWZLj5pdPaQTTDy5bRMlEW05KjKNvHj
50VwN98VkrQKs6GobPij0cdNa2hvMIgS/0RUPDmnHs9u0l1JEH8df9MwcapS
YhW3i9n95MliEJqLViYVlWBgUgjheE53gSDC5QGNPy0sGZsQFPFYrqPZVYiy
SfpxnJ3OHCNh0dJc/+6zu2iZLmihdJRr18e1DJ4dE3LoTSUUkBIF/Fje284z
XnS/hBD9WSQttGBnxM6kFEBU148SH0jjm36P5pESbdzoX90URtKfZ4UDgFuR
yjEH4cLiLDW3OWxQ2qAsN6CFNcIijRhufbrzCS904Xl1s7SGh1Nr3MN1WRiS
Qj5O9eRjf2oxWyW7nKH0ZBh3ObbbjrmIljGQrFzYdHOrnet4EMtzXeUhpEkJ
yk4QYXRqPN/J95iGQCffLb1PujyqD86M6ytq7+tb6mo7Mm+pRmr7Sak1Ljnm
CcVS+LYZHoNBgfbLmr6TsTqKKkTYeIW9H6VtEj5DXIVd7WaPFRcIgrb6VNEu
ICI3yKNKwRb5HZ9roWq4Fcmug0qbSWBITkC1g0DcuWs9V4YMG1o2jHk8HUWS
KixMakzcWY/DGjRX7tPZYdsGw4MgGdyXeXe14BxYmkxX0ANbyhtPfTVcBsQW
X1dNbKbGlVbHy8cnij8/jMHfTpfAUiZKXgrgLwfe2nNyqZDvLqbDWDPCZzPh
yl3ntk7O+Enj/apyxkcgsQDQkDYL5ePTwkgKyVWhyaxsj7WXPGq1+A9TZogY
XbWR5ZNHH6zeFIyH7jmCejf7L79I9OcKtinsD3RisqhUjyGvw5ORie+x/tLh
5CMcJsQrd+rTLANW+2wekOF0xHp4jeeBzHft8/W1hJjzg6fjXqnemOTBWK4V
HXv+slciqIM6eEUSvrhvI9enVOZQLJxAHuciLn/sbR6pYh/8rLi5YLym8JP6
sdu/W8RRomkZZSzJiZMp3rlKufoOULNgajLlx/rKxzArv0yIvQPFS0Or2iur
Jk53cmRswQvJmTWI/YjFQ9yYl+ArU8NiLFKuVh1vsldfH5ADYub4lqGvANNQ
1D0LDyk4NQgrtScelfilo/iccjRXBw0DHD9S6+1bk6aJbsdLo4TBDH/l6Vyh
fvviWflXFF9Xl4iOzTK2TfPM1D8K2u3FsKWQAMEXEaTSRm7hH8eLPpGpPX6D
dW3HKvNWR+jEDP0z/7rLFsMTw/r9Ev4iDd4DX1SpJx3oFNWRzIz9OumMGJ0Y
vs65kMlmNEBgurpclpR+RIKfZxaFTrnRViMi+juNxWgfeHq+Jzbx0TQbfZAZ
hEQt7unSwOaj+50eHnvS/VCI7TrKoA2wxvE8TTzUAYXvVFxzl31lKBAtvM+v
6YWzqbLLaz5WIDXFSKrFNDRZhfVXqE96qdZ1XxGliWC2k0t33YoSes4wUu93
0RtpsM+foY3r1Iwbk25MHQngNMkvTkWjRXToV2+Yqt+QrPmRYfO8ddL8f9S6
aBm9NbKnEtqxsHQci5cywR/4Pp4+8UHq6pBle6kENLZMKrTaWRaEROqrkPoP
+hlPXpmXgVS8bGIE75J08xTdOKTFS20fmWlIDtao7RQMlLQ+1APb+fdC0MnJ
PMzkPXkZ6tDOW/eeMTZu/O75hffrwQ/1SYFNeccfLQIENuQCMVtNXsUSJjwr
afHWkvWEzkUqSoNZ6mFXtVtWD4EQSAk5MTz9yHRLmtZCN/dpVw3oiLrrVBJS
bFySf/5YWJPQ9edE8iyCR7LG9F1Da8/Vmxbu6v+Y9jGqWCguCA2mLOsFjvBK
f3TYrPu1qaqQPVKpJc3JvE9VWDKbr3aZWevbCiLeIC5exKuhPbSC1hOMps9A
Qkjy+XxqaxsZJQxm/8WmAQ+mny1GpvxXDcOqz+lYHQIurxVCqc2VhXJXgPyd
j7F4s0yUE8vs8Zhho2zsNAG+6+DeAM7i9ODHP4xseBE7a4y/CfaY//jCmf6R
8pVar4XkCQrWPZ4SvDVmprZ8cyH62dEChLcVj+ltNNtqzUfVf01YsLEgCwKg
99Q1UpgK+0zjNIs0d1gdc/U0IDW4JG5Jlwn6YHqWhaeoMhDpcfyEgsUbu5Hn
qq+5iYCm1PJTi0iEWHP1kES0YkGiTFB5G6rMUdpUXZXDftECi3fXVTyD8as4
0Hg+C8GSVVuy+SFhTvQtFWDFT1kosFAuZiRYdVn9QncntF3Sdo5f7dXCKVN0
jNgOQtKxMtyLqEgMM3haVIOdpOtnEvSB88aVptQzZXnCwveE4BB1ZvVjjQGt
/Jv5UzoYlMD/JnMveas56NrCpmh+3VKAOyTl1KyLW8jqYjePsJUGTAymtj+y
YnSQ23vi01glQWuupUtt5kGQzCc+HOlz4uxrJtA3nNPnz/3MAx2bzHYwlFpJ
agm7ZT/TdsR0pehBV2wqrzCtbyNUNEmYww72cBXDgA6W/Au+pqiJ5BhBkHlS
AFu/N6blypg8ViO0P8q2wxzQY9uqcuVtHMJkmX6oCu4rSibo+wwjmrkZrStr
QzpxIhLzksZ03dB9yuRg3LCg7opH1HKFfUYf99Hzx75nsrzdcJMb3VvMzNjr
8P5UwOi6hMSjNDMs1Xt0Rc8yUztMnQoC+sDH1pWtk5zDz2aNRfK0e2N+XSKZ
vjLdVbT3oJcKONqTI/VAl6NtyDNeLDryyFNvsw29ngj58LCRl1CcJ8r5r0Fv
h6NdEoKDaubIdXd/XMP0l9MnNu9jb4oRKpQxSNdt/AS1E+XrQNu0N9rIxggq
ytLjTtGvbwoeancSPcrFpCj5F/OSKo08jxJDCmCvZfVyKZBnMpxVvwssIZ+e
FaVvVmGaI6F75B5YGG+ZjRUMItWu/9Xe4UEQFIs+wWQbxXdF4kIABQZR4AlI
EsQ6jDgvNLWQOGFYG8YOCD167peffnFHOtuMQY72rZfS8FcjY4q08NWhGzWc
+WcT6o2h0Iclq2YbTwSqPMF2ssLlcYerd8hRd4aU/TwIqmrccHVXS7epiSF7
EdHTj3bJOdoh1+JcDyCPfFuoQFWf9cT2dOesqR9+bPzrVV7HHg19Bsr+WLBx
6Ev4XYB3xvS6ywlNvhF0im4ErmPvHQE57CroJB8hwy/Oxn85O6X+S6Dji28e
KzoLZ8IPLjJB8SVFB69ORC7+gfuWRJmC+7lHE0fPe2bB8Mj1oXHYeR9f2+1T
CuubcwDT8Ki3VZujJAKLDKX7fZI5UGi8PJjPIDIdFjxgduxCb+H4CzXmzuk/
o8DG+6jQ/CFEvQIR2XXd551uxBqv/GBHCNUJ7+8XyPlqX7BuaojnOSHdLpcQ
7lb9WiS+IRpo1u3Xo4wy9hirpMrQSsYa0mbiCW5JiUdpygQ7EvJL2OlCYZoI
4NS5WiONd7PYYv0PgOlU9Pwcj8FpBEXaJqUpw6rzGE27uBZvZaiWkO7UAotD
W3hbtF0ERc5gBVeturaU7b2UJyPTUDjHRcNY01HryiCyY3xM62EN7Cok8wfU
cKsP7oxQnQw1a3q/+hFaUnpxZmcYZ+kOqbExDAHwtzwgfqqsrQ+5D9oQRhwH
vILsQDE2rNV9ZPMOGMIcD0Qu6MTdK1FpUThVfZD1sPwqSTQx0KgOWP6p9buT
QyU/43ZS9J9b1IpwptYFDQHJgly0jRcQsWddp3F+VGncoTSJfitt+5Uuajfa
kDRPHE0TcXER+JVrsYMNCkwFAZODymM62fpNLZIJxA0i58gzGukCKzwoNmfA
V0o9QLjowQHFaQnqK6PuvW2Ic1Jv6mwmlgjSiLiu/DnV1LGdwzN3dXqnS2Js
Z79A7/ZsKrmp8oU4mzPslJpUTdcUKISHTaP94QnFVWYrBcviy9tITQFEhiI8
Nvy6b7hfg6WKVhUTjN/WukRmROGFmzrPh5YDE9m8aPoRnAhoBgYpSEIADiNH
mCLnqdHUOpc8GdDUJRh3X/vLM3eNAvQgesXc8JF5FJEuUm9OSwkaCwIHe3v6
s/G0BH+rV22oTh57Rj9VQAYEsizdr5tX9Z4dNRXSn0oY7uBII8mMG7U+2CsA
f4z8iXHLrNjjK3kYGj4FHtJMUxHVq5oB64IfZuJ9do0e7/u2FL+3zF3LO1nT
v9EtuDW+V2opVEASX72g9Pv2e9BLo7jOO00n+5bqkkOQYrMqJHY6/HTVrQsW
7OLg5pRwlUhlyGoukTp61oPLSSCPqp54jVu6czbrRLIlGJm7A1E8WmS/4ilN
7jyqXiRNL+WZbagtSjNNT6sN/toJlcBEhe00SQ9Gfi2QlCZlxuixrMZg7blB
zFMZVqpZPRJtsq4OuRjN/IXQjxqM20yNH1qRuOPGnj3Vo8sar39qgWSKlBzk
Yzb4I3FuNkuuv5pknJgSGRxkLnYHh4iyC7Xt7BeeIZ2HH/zgTIZ2PxFmcVJr
qRbqRfqJLnW7OM898lAVuLvYe6ohZbvFBYvDTAYLwtCquDP89CBJ9DWo7QGL
b1a0Pz4JmYMoP92t11c7ojyzAWQPu5V3rPX6EJ8dRIe+0H2q6/A8OvkReAL1
5IRjeMOCkQUKhVZsfuH6dSZ/IhL5u1noKKyDTxWVnFiRh1CxDFhb/s8YivIz
xXy3hT6DzfqybR8MdoLDQ3jls18Kh3ajh5A/Q7PEla3FiR58IEt5XFSfFOvh
fHAycJ+vR4XcUYRo7AT+o8DFXKh8V6aMoYtWIUQeZnI5pPR0PH4ITXhBmRbZ
m5Zu2n9oAO89R9quWIl9yuNLNccodtyPfdm3nK4Sj2FGl8wZcbxxWkLvLtll
1EyGuBqeKfPFh7ejQo9KlMtTBqo7aqc6nDqx1Kk6OV4Kat3GgvvhqBxa10Aa
hKcoR157f7mxRsceJZjU4oAMxdvf5nFhoAVl1Hq3w6PUSHp1gfyVaLDzqJOV
+IcIaNEvuZQb9BAuqR8qCoesTZPlJg7TBroWG04ep/CcDO2bi6JMiBgfSWEP
VLO/ScqGYtLYxBwjSCIz/b/EWks3rjSbYjwDodJwKzx2zO+jUshuq5rVhy4M
ii8Q9f9KRgV3+JAv5tLrkPkUaRVA5uAqgf2nfbyl2OeaSFwl4d9DfQ8c7xAN
5l7vD7eqALKYcvgTnIDrzFnfHOkznT6J7IfRAgwHr/4WWcK35WfPK24FmDiO
0YyjUYNvqgoaDa+e+mpu8Ak4+bIUYGXkNs9lE2FWbuk/cBvvd5Wg/c78sCvS
bBGbLYkNkUzGSBhCvPa2Z9EDT9wZB9fEV0x0ZxA55C75aVQPzZ8BYYRoN3/8
iiielfZyLrE43ZFG0ZwCjqbPoDYGSv6Hy0VYkmx2Lu8+RpdW7xwguRCp2oEE
5hk04oKLpCmCd0zsWk/b6MJc+s2y6d68Jk/XVILvsNA4Gc8OFHYydQXUzFTl
idRVWZPrQ6PP/AZYtmYYXq5JEvBjMRbI+UY5XqrGplTMU9E+GqxtNFO8k1jv
Sn6Bds//zhe0m20ZjnIN3tWKBVdYIr52uB2hqANJ19mT5JmRehqqTWwl2NA3
7PqQBOTRXbyLkfo+/+W7pSIwdG3YpjFv89O5qVoFJciuRe7i+xpv8Y6c0z2z
zzQ7YQKryFyqCHjRSXHEqyzoDZG0/0OeueP3uiGf6qWwFDzRBeW/OMm8Jtc7
rp1qtanNJLrjGRwG+KULaB/KZKFpqs9huGm94Em1RrFlM+yeVJhm2euVEkhc
FmiP1oGi4YVfCkO7vBb19CaEZ6dXxYp310F892bBG9IgmXVnWSNDGEbsRPpj
cgejrEDVWoWYQOh6KN9D+IHereFI3LlSegRoDHQldVu8tdKAAoEOeEgHpMq8
1A8AVfF2we+JpI9X/DTB+pQ+wutU5OdLjQT9cJWwvfqcV+OqCln/Fr70w1gR
LM3qoaUL5FPMVvcwBiMF+VnYXHjDxEaFVTbQO3VHmi+o15pjIIM2ojsf6rD2
bYsAhwu82F8WQSh/YbDbhiiCppFjPDIeGhy36LIi5FJeuJgn7zUV+H+BC01b
U3jSYzZtT1kyXqnhEAhxy3FuSUWKjY656pVRkTl3vC7Oljgzcrpd5kWsbGWJ
khICYgDGHWqImuJkuSUvYj0yr7M6heVAAXb1x+aDoC1NEw5LJrefeuUKPsuT
b+2L4lpy+a0QXYlp6x3A6XVhKjXTZIGuxY39HvsCgfVpaG6B057sVuelfA4Z
3+r3qMeLq0HvoMuVe/e1h+0elXbigHu5pGU2dFtx8ZVeFlFvCR1D4/msDNmH
6CBu7yjLGUQ4+Wlz6X4MCPV7/tFCVfc6EnX1XE46MxzWJlvl18LYVQ4chLiQ
McTHLw0fKVvZp+YEyiXZ3rrEd+KgWD9n79LShJ+wCAYN1fTWtOZIxzbvTfLm
Il1OCZQMYdWBqVuw8lCp3qFty1rLUEjvod0AoOSm2IvYTleoSF7lU346MTMd
Us8OlP+V2tzIJxRfSd9cq45IzKQ1QdBmxrcukEXUzCeEL1rkhB/LAZa0d4Zt
51WTmUuweI/mdVRwvnfp7g8BF4f6ik5CynzqOmmG0i8pfa5U8qObKX5KoUqo
B67L+I+r6wB6FPe0/UJCRtkEeY+Xt+kg/zQpv0VXgDak33e0jAZKIc4tVARL
2rumpFBBccuUMjyxW9v4r4kdXpl2s7MU/FrfBuQ9lIJbSZy27H0a8AT1ZRal
YgR3CnbTHruxmfvBMLj71WYERNagh7VqBFdDkElGPT9gYue+f8UV59LaGsqa
1clWE2Ypb+il0Fhp5Nr1YxTVAL3KSh7+Vx38jGg0iyc92DaLY2qWk8XFpuqe
/rozHhlQt23Dd6EO9LKKy/8WQbk1FP8Q0ir9h4R7fSVhIsoAZ11iHH3KgnPK
dfrsdUV7NsLFa+ZPu5Y5TbrzkMn+FtsAGcuCRnp2ogxlNVJa5fSee3v5JEwA
O+JbYGsWRWLYqKGbOLzWHaOfZU0/TLz5W5tSmTA2oxr78K9Ka/X5A+QPSxk3
2PZrD2z7CNu70ZcKZ/mLV3led1dgLAzalar3OGvC7ups8aw0VldPvytsCMTZ
KbTMI867BVUvxFwAXfpno/IPeHIva48WxKw3fogrRy3uIx+sx8W1b3sjcd7T
5hTIZPDI2ACgqPzerCi+Wos8/BVG4jxz4GGIAy9zmMsaS2flQmyA0J/1HMau
8tffwemgG0qc2VxT6r84FduUzsny5a0s7k7ydG5s9HuHgoqVM06ppkiULYq2
2KjPRtGPT00Net9eIJxugc/mxP0q+gepQgzmTv3zuej1m7x9Hl6GkfI/71cA
dWIR+vT/w+a952RId1zmFZ2aptgPxkA13czh4eIG8x4Y3HpvfzcpbVMHdyoF
rGJuZmSAcKlOeogK09j7VX1leNh/6ItemVChBjRKergiRIiESQACAbAyoEUD
UfXuB9M4cio3d65W8euGcH6TDvLAv5UORFEFPMvECdhhFZlsXXHl8Ql9BNjP
7+g2K6UrU7Rc3sFrKOI6S4kTmMErM2eu4JkvQQz+TYCyugmaMfvUlKkK72jp
oorBP9azfVu/3vDYnbeGSMVA2XFMttKFo8NJExA178lUSnf/kiPt0dhHrwFG
O5voR0RWKfUtsUPmSLbptWnYSo53XtBg/n4kQqbG4F1MjyNIIiWbyIqTD8nG
BivViYSs2+tCSf//0LKfEJ3aQ3R1DQEr3ttsN1ULsF8c5DQdTobodwFEbTmI
gBI6spxymoEOaF6LLuLGtg7lnnVgqt//n6NNjeTe2VEYMrgnalPZXREatN/u
b+N4ERqC/56J6bgprNyZnep3guGDrtPC4dpz7ABgzcRIRD3BLg3jweCvsvzC
rzYZuZ00UBHQ8WJEH+W1vQ6wD5VVQ/vcrBGmbVGPar5IYiTIKDMHQ70yN/bp
e7/8IpcmDKNrtGVRRE8i+wOwnXH/8dLIuOmt51usGbqU6VNUwvqh6ntddMIX
v/25Xv+9wpD5XFLzFpcw5VRyXQj1b5uSqDJovaPoS+I2Mi0ysRQmlR5qiiE5
zik4b3cHz5Z1Y0NSLYaKLaxaxFdd81WJHe941cgyfYk7a8GPL3PxU7xoliz9
dr42qjpUojt/8IrOoRbl7mRa8eEQwm2N+vNomEycqRbfWYS6OOiGivmxHR8A
PcQeHyYPluvD1DMIta7RcFFEFe7tHtp3pqozIOn554df+KYLdRATGVxJ4QOS
Cbnd2EHuJLeKlkbog5U5clNLyJrfM9EQ4fSbhZPYZ9j6ZD3KLGTH0qe1pbMg
lVp1XhcrXsSUHNYFi7I1geUKTFpnq9WVHhiQEFAklbi91BUxhPy4VVwYagB6
n6bXBEdvJpWGWm/9pVLrrmI7IS2z1t/dTJ4AzHmjDux33suWeTev0RBIbtG6
3XWLKJdnkXtUcsBq7CvuNCATGTSQW/h6ZquvEQiFAbmxnTfzlzbo1Cwfm9si
7I/5yBQKbhfRHY4Mfjh5d/5+YxORJBIVB1cplqiigbEny1BzM4cq1CFtGgaY
YmKks9swFpB5OZlT5g974fNllrECYzlCtGSAWhEhym9gJrL0gXiLpU+ivv3B
ZtTWeZhCJkEcIyRNZ/gcVAJLV4MmZ1JjOPcUaAyAcUhIZN86C05hVNgyoqFF
P73iyYO5hoPETCVb9XK2pNmSidCnoAzkEdF2+osWWXfw34Rdw5IDiPyMpnQ3
c0fn2Fx53QEdwEJ/CgkeBV9qHmcBu0zZ6SZ9xniOge2yu4u3gb9ti7HsfQ+c
U+cbVwsP/JuaPZkLozaURBRYAhRNd6+QIHfJqhnTp9YVNS+ntG9hy+PAm9Mv
AIkPv9r8N5kyBeXrNEnqQi5oNUALPxxPJ9FETIppZjakbmoDLQVgjV+BTsHl
44p+NuXNuyAgnIZLQh9HHCo4jFYIVeqtMfXPI3ue9HayK1bFrURvihlj5nap
T8MXSt9U7gZwctoqDQwMuIhuosZGTiKQwZaWMA0v2blmW4UWiCwT8p12c2ww
5Oh9/LjdknoegSbXuCzpT2Gdl+vid5Zo06Fx1o7QRZcw15NPzw3lMqnn+OUa
1KL+BQqOdq24TNlBllZeL15AMnxPP3uGxDJYSMy7K2SW6XP0oB1ZktWLfBdd
/yDRd4xypQtANhMr8HY65J8GnuYdt7kJgRJHMfihZ74JS0fQ4GP7UZv4ARuN
eCWJ1QEb59l9kqUWSFBkvDifiU/4WSVhA6AI9DROkkL/EJI/yp7xsiJmXiqT
C99NZMujth+Q1n8yWHEGDeo2jYSq8qNASWEZ1CkBoqbh2/qX3GaGDVVMjsaN
Yayw+QyQzDCo0xodkHM+1+gHPMBilW3JCOGvtsRdNTLIv7i/L6JL3pXBxI3u
X57R21FHOhe+luqTvCwq7LNtguPvG9561dv562KVCRH8omYPOAStG8/tOMRs
pLvawpP8tZ6beulpmvTOsV6WG7aP8FGT6tXZn03G5D8z0g5HOPi6dSaYvr5F
MrDMpADd/AfgtdSy5pu1auEjWMUJehZGjnmFv3JUOWZB8ceD7VOiU/sn4P6Q
WwIuogAvD7uB7uOuBvnK98BzvNzx0b+pNqgY+GKE968+eITl1j09oH0yfGi2
atXTlsVMrW9wdgg5IVub8ko5u7008fCayOLhgZZDmRb6tBqAqVJcpCxgCZFr
Oo3jYW6vm1Clr3C5c5pT9EOoorR9Ln2dUVAxwCGDyDVclgp4HBnjIIwAsk2O
8zmutlJiq4b1KatYCYLMGiGFVd6lW5Q8lZe6wOQpqUVifehx5TcMIVViVnfZ
18N0bPMVXszJZNApRrxE6w1esFo7X4UEXAW3OUmk9xIFcRqPB9nj6k8ftuuM
nJrvb2YuLx709v0UX9+SRzA8hwmrfmionkbKfZRfs3rRxdp3xKZN6tLt075s
upasulg25xu2iK6u+qHF3fwMXP1hfrVhHWj/yrQusqF329bUmJO6Y1y+gnCA
4J6ST6B/uws85JGADPzf967W+X4+ZkIpHKhgOpw78wfFP9Lv8cjIgigxiBtD
LZoS7tmaJlLXyFuW9KJ3OAUNwGRtOyyaAxl5czOjY6Vaj/C9my4DotpxU9Q9
SGu1kGmWk/DLAf10YzTN4JuiOfFQ7JMKyUVFzVHLyrbt1wPHZXG+zEaO49Dv
qIM6TtCcyPS3AQBNSqo8+V35aA5j1HgAja6//4im768CxT8ymkatVIGhK5kA
tugiwSEssClukHLM4ZMY8O01yaAXdOCz4+wEHf9uqy2JlTrs/04s/U6OnIQC
kB/o8W0rnPJejSkKLqhR43DCAZVJFrYnpHify1e04+0txNKpSGagQcpMAYEI
+V5zeSRjrCSZHlSDPB+Al7yW5ovbM1yoaq1njS3lAEiA9qvr/jF9mMpMjItR
YVw7y1OGwQo+VVt525EF0RM7R1r2xQftQQcN6lAfp7ho92Gz67KClvC9iEbR
hepgidefsgtUs+MmK8NEiqw/GjBBisFYq/pxuh+6+AHq98gMxT97Zfef43oC
zEUpiKxTe8jNt7JeOcXtZ2v65peJqsJ4w/weT4+zlY0aFNqizaeZxLp2mx2x
HO66v0j9BecwnkeH90hGZJCWDd/SfKIihYpiYSwIZ704KZpdBFRJ7uXpox1m
gSMUk+PtCUE8aGW6JRopke6IIQp9w9BFveT05D57MXK9uH8xesSLYgAhVJ+R
Gdzaj+uLd+ucQaYhVtEMZQmSmPmAvez2ZwdQE4Pwp/Q+uHFQMkMJh81DEdto
1e+RcQcE57KiqbpN9Qizq+xgmgJ2nXLxWFfqitsx6VkI0rqLYyE6zq7CLoEW
4HMvfI/kfYSYniqWc9s74S4pAxlDoLQWgPGKtxvOqLW+5ovf9/xgTOvMcPtz
emXjyZWR3ZZXCkCogZ+BDVPfuuXAQexrFu/qekMvCIdWbzZkpljhZ3fyyBHq
01U2vxJ0p1YJVT9aHtCF08MyotUuKiUY43WAxFoKJECbdKfIBSSW4YZXgv/F
0ZFKErhCvpJYOqabI6UJAnir7Xl4FLmS560IUrxD5FXJA8bpiLkPYxhvfoa7
DvidFFYbV8AluRo9UuV4oPhWjP9W/QFpmyT+M5pb1DztprfE2z6P800apk3O
i3mtSoNUQZJ6WiHrB+r4rQnoSQdP2OrhYc+6u6xRxWATp7m1EgpsNPjb8/JG
MKRQkRsI0W4GszbKZsHX/3G0+9nN3Re4xZNrf3zdWWbi1T4H544L7udOxJzC
MCD53y9yhp0FXx+fFllRRaicIIx8ZVFVdIZa8ynhz15UlvB88xogC3bp/0ht
cpCyZ6QY+Z70sNZIXQpEnpkNqZ1xwyylWT1ckxbIRqSP2bSYMbzZxZSLkUBc
h/4/WwScgdXJZSJGXTj5mPKDY2Em05MXeUleiulzGeg0rRVx9VK5HC9v07p1
s8HO/robY9CbiS7he5k3mnWdgMqdZGRh/21Glm0+1urPBnjC1n6WXxXNuLxn
uWkzD47F7zGc6J+OxB0Q4LUNNNxUWojOtltptbafXDjtD6KTrdlKQ9s86Ut5
d+Cru+jFEkAh242uCCOR1j6YO+aWnR/hucSRhb5NzdTUoX5XO3XjOG0CuIoj
5YZkNP1DfFdNOaZBbgbyq6QBEd1LL+A8moc3sxlSyQ6nHEJNRnP/EiqWB2kR
d4bmVAjeF5V0ztfG5gqrDGtxi88rh5g1T7LnUC7SHOG2kYW9nqHZjfdacwVN
lQidnOTI+LC07tPh9/1qnwfnX3Z+gkVg9sCtrAqRI30DghAiz8nNcIMkJXNJ
PqnBYhodAZLpVMFWJOUdZfl4zvfy3+XXtDr2rqoWItmb1zRveXjHwOUzNtVt
5iU1c1+SIWSKoXtzxcwUaGQfYPN9VdW/kF22j+QGoM7IeP3HA+CyXm5IPzUF
iVhSgu0MCYPlEmWiA6Y3+lpZZmBgQhmm8P6nbkAtfbQ1WcUEQhEqVcVXo422
nT6EC7JIykFIFSJ2nnW49nqp0aVMa5JL/hhgnzWo/q+oqpxoVZ+mvhSO87kT
pH9/UTbRkL1msJuO7arUy3TcfMRPhCQKJkMG9FnKdUePf7bphkEGxFTIYml5
vTxeF8gYW7IFLyKBqQw7AXfxNHTI9QN30UV+VtPzIHpz8lS1a+DKP0voM+/4
Y6u6CQUVq8c7hzCJineCrQcX6WcctPpQLcNxcn1p1M37ULnyfQLco+SQEI+e
LkJpO1x7cVUIsRB1p9jo6sKfL77mdYHLmx1M4VxBCoR247k48/RYtZDztu6o
x/5ospckpdX3gtGtJSGpBlRdiV62IiXeXD7e/kC7NzUTi5coh4c4N2DS4XJz
Wg4+S+Elxhem8P/6N2WAWU+4cPeoSa5whdPaOQ3oW2sIAxBU/81bINeyILy7
BERVntDoKnD+AvUGNqNgn5Swkt4S+rZbQrKX/lGWRes0YfYOIP+GvQBd4u/F
BYOgVxYa1guTNdZxkn8kuu/Jl1ux418Ud5ovaFlDVMCg0ljdGP3jz4sowYJB
54l9zm+KqE6cjIulVAmLXiqY+aWo+svHP7SLXL0bcodxPSUaWoZzKHJ4qMNJ
YP/i2OtbjEiRw/3+bQ/eCx36wXkxEgyMgab2GqBOQhwk9E2j7sVO4FI2QAxq
VCAXhN6hi6CvoB4luDYpW7KE/Hw/e7EeWqwCgHOvQXzIQFr5SAbWER/94me8
zmJni2D0AyR+PtktlK88qWhjmUqiL/wzKtZFkDgdHSTn+ZzhUfv/siOICU8i
L0LIQuO0DaGJTRHDeqN97j6wqFD7CpR5Di/R+WlzvoGP8qtRSgekEyU31kYr
sntTmptGt9MTsBx4wDRcFGGZ8dd67SXirVRJGZEvzVSn04f0umOKGgh8Lwr/
PKgagFNq2sFrsXn9chp84LEXzCU09umdNVZFnlXOYt8kOkS3WcGdr6LWxo/k
BTuiX7PyaepSuXCcsylpO9j8m2zOX/+lXZtOM/SAlh4Qs+jtGYZlKlzIwqFQ
KPfiXTWRnwOqxSEG7vHNum05ZOOHm9n3UQ0HaHT4v1Tz3m98ZConEq7jUohS
zetYO1Ilh4JZW7MoX7oweAlvVhdMSyWJIBjtIjF2S8zx7McWISZNCRfQYXeY
bcTJ5qH21hdGd9/qQl1he3MKgt1x6z2oBJ4rg1EgGDaL44y4FC8CCFfwZhYy
sLXrl38SSccqxH7plS76F9WJLP/XKt803anASRpAAe0S2Yj0rtjNX62NUxxZ
HjE2tvZkGIxauVCEd8JlOLOS+eJbvnCztVcZM0b/5oEw9F6h/vY5VeGnikJ4
UTtLEeVQ5OX7Z2LqsH1rZfZAWgw8e0juHOV2/Zxcp5W4SYoXLsoi8g1zoqlM
9aS6dUrlxwR95N4Gv3Lql9DbwjaCgemSAz+XeGeGilC+Bp75JBwymqotbxVu
zdNFAiAFBMPd3C0VxQNxAj5WJM/avLZRUIHlxcMjw+O5UbyvbQTgbwYOQ/f5
nbQgorBN6bkJisCPJFTnHu1A/maPIDONAmQQD70kl/FFASEp3WBmvs7xjrBP
i2n0yw0ilzR1BOFP55DZUF0RNQ5whTjz2JDq7EnDj1x1KsauRro8PNW9jWr3
GGIt1VuXKPtbJn/0pojZlJxLOqqGIfm/ky+rQGX0+Bzf8QPucobBFD3aQfIf
mz9HmsR2abRcV7caz2mRf0AUDrQNeZ2ni37WVwTQYamL+Hf1e56BMNKXO/zt
kvVeMshNrNM9Cc+GjPfqvUGy7RmYZFEvYHpsmeNU+Tgj7juH855YkFTF1TKM
lIjhmAXHM7cYt2AajSWPkwGgSYbdldzJgntQoP9o3O0tsctktl3oPSLQFlO3
4vZEPLpYpoK6ZqCe7ljrYjEXgL9OkvXXXAgpZVNkEj+gA1ZOIBkyY8J4FwFx
pDEw2q/MtXFnkIsx/v8kQk2iWpqFd6JLzBDEbeSvTr+gJYys6l3Bs0a2T/sS
k9R+BNd8PZ38wNn/F9Pio3zv9J2ib5EXvaHGw66EtxHaKMdnwXwWB/3stW2+
cEMVct3DPlrZS/oYCyxtuVbnTD2DCv8PI4rlRjqhGUhR3pBAm4S6ousvXAV/
KQr/d2Jm6atu2Y1UVb1RW1H2Xctu8MhR1+1NTE4GRGOjzPSpeFds0j6zUvyz
tQfhf0rlRCw7RBqYjuuqbZ/8md+V0XAv6g5Sq1nNZV8qotCOGd+iSy4TOEck
bkbJPd1V0X7Hch+cjATX1bx5mRv8JBsMqG9BWd9s/RJqiw1yCLAEYSQSF6Cn
9DYeYFEe1tE4MJLE+3IG2egAd0AOt68JV/JG4zjP0m+6UNg7Gdz57KYkK57H
UxcDieVzflisgwVT1lbtWJ9673jEqVJ1/H4PdvlhzvU52lnggYl8y5Kqtht9
3v7RvL6VPAWR2gOldaIIhYCflWsFYfZUlaPyTdRisxk/4B4J0rr1wd3/DCvZ
gOepFupPAiz8QC8cME4igL9FK2PyXu6BTw0jE8Qy6lPa7yb7dyFrm8EcSbA5
69MYk6sjcS7oA1gwSfES1aShKqkIUxKj65vLlMWmy/OeMScXk58ZysIW+/HH
VdaUycNPYeicAgJ74tkA5+v+hmpSUqYIaiIcXxV2nDHDSH/DlAf+HOtZMkEU
poMyu52eeTjvoY9pRCO2HxqlE6JDBcuSa/H9pInw/HG1/AuvfN8M46QVnlRo
n10ubqYe7pG5b+MlQ/nQrpsHwEoIWD93WR0HiyA5pkhTh871i3RY9p8mOtq6
IoKW62w5oqVicaUN6wbE7SsQgChzD0iemAupnZMbs4P0uAx3tvr/BvZIdeoL
d1DA0/t2WWiNKK5rvJReGu9qEAFiENB1khfinVH4PUYTbNjOqF/6CRyAS2lB
lL6jhH498+MEXv+eBV+oFNivi5WI4jZBse57UmacInYkiYdleNXTTHckBSwD
BKfjLioZNMjzXNZXOCSO/cPEHyhJz8HtoREV3nFuj/lAbxouYiwRRFg2ZMBE
eG9fY7oDq1kOHffUK8GSl1bNRgJQxQkD4WZo63s9rwvn4lV4mSYtgEm6T6wV
37wTVmiVrIJ/sYCfhufHpqqesqkA6q1XFO4aE6IMNi6+x7Xz8vAr6/sOzFlK
G/BhP8ru5BnYwRuDt4snR++4467V3y2LgrKCs36WURlc6hJ5ndykCZpfQdA+
vR0JXY8QE0yFgYnGkaY6mziub63ZmnmOUHbBYN796bHKozLvylzj2ZRqIftl
J2lwr4ivNwSJmg5lVXFAX/DopimNn2emb4BfsWR9sKf590gFco5+sqJtXFRx
Q8Rwt/is1EDAmpwYbDWx7ueHGH+08PLva/H/EvXxTsVmK6ISaF3BMzR2EDdO
Un0Vg8tSXutabjiYGdYs+J4ePRx4L8MW9VbOmo7H9SGqDjwHB8uHmgMk1nxM
pDAU9ZUdJxDYQkh/2qTpAIzh1f2us4x4y+nMZxgLnOCa6tr7jQHbV4J3e2mn
N7cICa/SGFTTupxddqb95Dgc3XFx1FX6z0dFoWC+67bIm1Zs+VdSrsjhk71K
sN3NHQ4q26XMx7w9U2pZAFoRlZrghp3SSadhYtw7GcZtLHjTsDB495TnJDPC
VEj5pD/1Q29149P4lcrqJ+row9kwOMFpn2M2gz79efHObt1hxQRHSv0gW3Cp
9XQWe4UkWhjtdMAKCIAGIhOceDBJwIBcPFrnEI9eHSf08xfoNhAQ585XeWuT
1wtUMGNtl+stLPbANdaAeJVb5X+d4PMgaRR2JJYUwBI1fJgUvtpm9kVlXZwv
By0TtJs4LoyrtBMqgTDu7CM1uQaBb9CrlJh+f8Rm1Ek+j2Lz/XYpo9YdasYi
M2iCItUhs5tWiqpbRavdD5MT0nfL8RkJgbsXPiYKFOCND4qQhmt2verYRtq0
a/Sr70tJGWvA0ltTtFiCD02Jh5dvLc1GKuSXM45stR2hgACL9a+JRo/pttN1
WCrCxpTluwTpe+/7jXqCJ9jOgToflbOsmXRFupgWAZM/MlgTh3VtHKNQnRxq
RsXGEDA9zARansQsYzOaClpOfloyaLTqg/IcCpbj3iqSoz4bsewS9dz0YoYS
vxwh8ZGFTD7uBlaHSDoezFC9HaNiyHTrvu7HhUjWTAoXtJgOx7Ozc7/IbMfZ
RjJyKWaFoeSQSplu8jKOwOfmZGrVhBIJJZSSe9O+sBJrrvooAd9jpk2BnZj/
Zzs7ce1gqWO4d1LKwaqNNppLSXTmMGJmbbfVqBwGMLSomTIFLsxVOH6hWJ7y
2Ciopi5AyZOyvkWau7bCPCHZIdFZceQrSROk7dhA+rTZHrMjchaNXxB99Hf8
jIwrUSAm/9RV5JEfhIbHXv46+AVV3V6RJx3NEp/5oIkNsgZIqXfTmLYv/bb/
GW4WzQHkpclyKpHDbIEYPI/KSVqNZTCuMK03l1ylQAiEu99+8co4AUmypHiW
7Azer8vRoyyGJ7vQvTpazLV52ROvbEBS4Fqehk4XcMizgNGxLaPq0INd574E
jcHL9pJoj5ubY55hsSpS39VKj+nvOgSKgsKymIV8KaKB/ME9axnP/smlj+Fp
lp6wCOS222OSXiBZ9/Le8nKkUK83+SyFXWREMEIFS0JVK6qD4+DegbA4j6UJ
YpmlevYm/fYSwj4JpLGNkqt1eP6A2R2q/LC9B/D5MPPQf4J37OEz6FV5E3fu
ied+ZSB7emOWD0v8OKZQwpFtJCrPzGCTfxBZs3SWoU581eIaVUdBk98e3QSv
O2+HU/zHvcfN5Grlecieqey5iBms008eP5+oY7yJeMEgyTftLfDuvSnSa3Gx
lnvRWCyMbJW5e28RvP+Dm69c3pXiJm44lbsEUo56YB7tdTl0aFLFAqAx23BA
aqcyLacq6L6YNnufa/n4oQOVyyX6ZMMy4PHEU4CWIbOiMEdHnWoB86PLzoFi
ihIWPSKb4OktypS94THZY3ZjfUuKQ0Egj6XlFL2CqwgExuJf2V24ms4tRMvU
jebogN+O7I1ZPbPnfXT29uwEKQoK0CrvzDSli04e5l1LgYKD3pXAAH6LLa2n
UMzS8oubKhPTRouw5wOyQ5pMZwP/VsM2nWUQSeWUcoCvcWY8d9VEZV99flVO
17XQFAfzqwQpR7RXU3DWyXqVr1YM8my8vD6MQ0RqlSNu1RaI7jBFiiLfr5GY
XgjpzROGAzepBKIwWA2C5QrAfnDY3A34xzWYCFHkXzlpHDobtPxFVwMXFu73
KQCPj4O0XyoYJkIE1mEgnyd+eY3Xa4HlDAm37MXUCzercp9qfkytW2wSEDjv
BF0GCcMzjk6SqPHPjHqFqLFsczIIGvU5pkz/Tln2lpXh3wC0YyWVZ8i54gFK
gn5h6MFZNXB894Hk7TqOfN+6Lj5SwBzcEIUKiHP/mfKfdBd9Kvmbh3Kvj946
2JYum66OW+LgQzQtroVtbxk3igneBVE37vrccjY5gVsO6GOqVdN+xG8ZmY/p
ofxtlcafQAuf/RfU3CuHQrJ3u/aPiakQR9EBNZiDiGRHDBCVn4FHtQTX6e1R
JMpP5E7x/c7/YNoeBnWq1mkGB3fiZGr2P3N4iNg3S7KwjhO2cA3wYPI71yH1
WXO0PEpYKtyu8sMrT7TzuQnPaPABuPwlR1YYgf5M5Ts04rQn1dO9cndIt/6t
KLkpAt4TXkgXLfVtdzPb6LdwP6vDl+NsH2Wyuzimpd/QgCFbt1AnluVpWpE4
gsqkR/8U1eqOIDIF+o2CVQOilL2qPZPgkfbrZ/bbvVjf0Y2SEvYi+SdRPMXj
pcHDOK6zsqO7yIsGgVDeTH4mRiU6SrwJzrP1h+5bjL2D8y3NnliuiN9kG96e
kkkaaeb/JGdFS9yG7C97gUoH5Zg0BbiKxs1IUj+weoMD1kPn//pE4Pbe//Lq
oYqO1lDeGU1D4+Ls/09LlNLVVEorKeeNBNsRtNLgncR8xYKPZ2iNiNYclJdT
Gs1G07V/e673rAH1OBnhsQuF11PxtJccyKUNWc3/0CXiPva3tpbn0GesfNuv
NONLeWuX0mVZz1LvyNatSejDuGs7gFnd3CcyhiG4dqsaARnLrdOeugli3OSy
6yF4yvPGtj+Ke/uVBwWaC30etlSqRqCaBa1mk/uTOfLCVvGCLRLurd8p8KkX
7EbjtJigdPCEoufOAb3OE6a0dyRjNVX25yCU5yqWLTqaMhm+N1LdUhHxsmoA
ueVvK3s1rztJNUNUJVJl1CHuMdqYSmhHeCB+8WGiBpt2C2k7iLR9sQwjgQRu
MlebfPGdxE56AAhcFHi5xKrRyE41v4ZJYJQTOM4pKtIsHHThWzNK35E0+df5
4oA7buOlYB2KdACBWHielnsTDeoay+V6fdk9ZJjhEfWQy1yf50Wsp7F0j37Q
YtLexN9slnfgpWJElsjZfdEvt6ThCe4yt3necPlgtWUzDsvJMZrcapNcsHkU
TN6lgxrjZhNboWeuAsncMZu9wXbQtAC87CHBg9wrCcjlXQAL5hFp2PfBDCS4
Nm1KcCIWFlgFGDMAk1oiV0jbYlqw2qH/hGfNN4+GNSuv8pAw86zXCEGEjZpO
wkUXt/tw/a7aK+tEGXTS7fjT+99Ok0b674WXjpFr02d+pV2TNZHMTF1QUTC2
+7XX+XhY9GTx1tiEc1Hd1oUa6iQmMKfV3Fbfn98pW2Sp1vCQv8L2PtBpzK6T
1FCxBPF07uD+ta2vBYaTKz63CrjwV3Ju8TaCUyL5ViAmyJCTKp2gssk606OQ
6SVlV2SuzhHtWtJ/HFQM5wC9Ep8W+uICiSvy5+yXwytWKxGT4VCD/pqvupgA
Tlyab6w9hpxazLFS2QlUSKN4hchqoeroaCbuvZXbURXqO/ALYZU4Y2qJ3PST
AV74RxVfOIoGLiHewzdHfEzlBE2LV2jO2M+DZTlxI8MACAR6AJxsVykMTbqd
WL1eMJT2UI9OBnIsU1u5bt0Vc3jVqH9ZiNAhaamKG5ijgElqFPRvdF8qV3G7
pbdyMHRhE5p3/mP0KW1JV5OmekjKicKgHretROhpmsPDAwkyoXbmUKnWnpWp
z+S4XWodhfVRRGq9Ql4hYHgy9pZhItnZThOPIk9o0//gJbfRzQjEe6xK/lF2
UtdQ5PwYXlH+EKo5IjIA9drlJvIx70CWrh+xS6yjPznXoYAvRzoJLflz0zbx
uIh9tpxppv4Fj/RTVob7uISLQZZoED0NPE6SUgl68ClvmDt3aXttX7jLAuO3
o85cUNqKO8uB945SlbMkcVRjexF4X4QpJhWFBl4vCKXZdkvAw4unu1e7k5+k
MP2CX2cask1cIpVCSkpS7XzQZJzD1jlQ3fd9ZY2bUnnb9Sv3LUDzJw3RRh17
gY1Dr/wrNE9mKO0bLKGAuo1+5VX0bd5OqYctMkNBSzi6EqbH1EtfX144prKN
cd0YL3w69G96CDEeIMpfbZpikAWac2FOOYozGc6XQ/vOItKc0P5xCSvXD2GQ
O0nyVXdXbfKwkk+RLJi3w03x+eTMUPkfMzOFt56DbF60/sR0Dzr0IvZOFlEI
e5Rn+r72S1P0d/jb/yShwY2C2KUkN/Do8ryBeAmVvOwfRga6ZSa/OZt+uIRt
/zsDcAwjeOodvgSLIfDCLg9V75eOe+PfTWhZBpKMgu+BW4xSbnruk7VYd0N0
K/tJ3DstXlfL0hmaV6CVlvOcQM/at/Lb2OIdVFcNe/iTUw+KZ5v6r6hVs33y
YPHaawjwj6ntIkvqGrlCuPsdUZpuiDtWZkv9W6fjvSn+tA9ObGikIL2tqEJv
j+Rs0UDxDrAHQWReWZyKLCzKfoCsik5OCb5wPfBtKS0HH2sMcWnnBbabRraE
/oCLt5CkPr2vUvnb3eh6d5naMI1NvpXOOoPcm0SMPzajO6piWSAKMLafLx34
4FuWQ8pl1Ok0taA9lC++n9juQEZrNKhTNzCUsOGCGqHyRxh5SRW+zM2Op6Uh
0RQPuzRpF72Mbxdkhy3whY6rDbSOhcU5+/1mUFN4uZ99+8f6WDnG5sqhXzNm
k3TWDtxDfWEI3S4Hj0fXdAsReLmyVoejIQu/XtReyBZ5oSHjMAhbPzzpwUAm
LUZ+nSauh3VCwBoLipzcyBRz5Q8SBU9wz1/jj+VSJvobWVEY00swWEMOzhf6
DQXalbXy2caILbnw03ZMtLGfhA/tltH427CYf5T4EWxaQJ365VR6CIWkf3Ep
lKNuOp2/kbDKV+nYdAsu3dFmJyk8Yxi/Vsj5A0pQnJ2dgBdpkj9bmrOWNy5i
KAsLwyhmOQC+uKNIjTxWeXG4H/LSVd7+q+kQ7/FSU24bLawXTFeLGNPxvZgt
SLw3HnFwszDk+1zUOfYzC0VgBICNOckgMzBNnDt2oU/1H8sOtHxyM5oGw1D3
EGfrsnau1/bANxxxeJZ5Lo7tJLnlN94UeQmm3HHba8rSftlMxrZLSeo8ZznP
+1rhxjvxQ0X22vZVA4i8w58atw2pPofIyAh+QR1FDiU4Hki47s3eP2L93e3e
J1TS9wDdLg34aSsFcrVxzOxPVLmGhkGkH/mvV0Dc184KI7RRhvgN54marazU
NTyhH8dd2zlcwl9kcjN59i8XqX//xQrOtzIxMcLJP6xquGOmhLk+AS0eMcEJ
NZ8E2/ALNDk9DghQEoJALno/946sKPTmnt/T/cLKEQ0/TGesSwTA1tFI+5SE
Rli3QpRf5BWOpyz8ewCHSYPdd7oqwGlxSHKcR3Pg/S+Z5VoHDSWgfhyhD3SR
lFpXJKwqaTS7iYvE0ITlvdT6CQgeveBxZtbqfXTtuEbfeCCcNSM8FEeletDR
Z1NbD70pL89eXq99oqE8uQZHjXk3qojWSB+sGgdyCpSvgOHIs0xkeLSGZoVL
8Tn3eU8t4PeduVlOeuCXT9bZyx5LL/CLztKiMbkkB9AZd2+3GSgxzrDSzxpq
hzB1EAzr3YfnpSFRmyyOZfuPbe6n0pzO33TW0L0whAlDZMnjuLobbKkHoHLU
RqNZwtj5yo44apVHahrKgLObRIAUcXtIyNM1Jo9Pnide3PPfNxS2A+gATNNy
xRivE7Gf8gVCKpKVSpctcnXDSGNi7T4jaX3tkVPDZ2ip+GWed1/x448NMoUK
is3kNT40lXHcmavebNh7f3gTxru4Rev8MuCH7fbifv23WwiUdd1KKc+mib+F
PYQ16YQqwEWGRa9UZtcb5247vQBlCuyzSF8QAE5i6ecXRte0MZvhfz51o5SM
rKabW8V/8zqwEIvQfUzQfzSjax7oZZ/BiFE4/WSemfOLd33CQyLaMjoB2UCR
Rkz+5fuT+dw0ue09m4MoT4WgT+EhrLKquWN0cW4NfqqeHP8JmVTdpOlz9N5J
/GqZ51qEOH1nuLr7dN9BJWR9hX1xhoxvyryC0jTBFZQtxGaw3fBxqqVsvIU4
M0lbSU9GSBoyNlkf1bMaRBI9Y1+PU6OvAI0BJaumvkrP+I5mTDN6pUdRaOWe
BlPA5I/BbgK1t0Qfq07QZVMo/0HYDnWdP4URZBes8eH2huk4ZmdzHlnu9woC
+5u++6CMFHdIRTDSTQ8jGYyA/Iz4mFYdGTsPhm0IbZnX96cV72b3yFum2kXh
rSm292rZLh1pkOhmZYcjsnRGCLl2BL80AO58UtTjIM+bSMh4+ydefNSKyIfQ
Ja8hS3S584fttsdM6V4L3l50X2bZnyOzp+nBLcZCgAhDm63/OfQlB1W0RsIR
FTGYLQnDYKzj7u0rUS44JgcOU98afM9btdZ2OxLvycP5Ed1bgI3zOzQkn+FH
lBzSZgImwe4bSkpb+O67ysYtDYtSzGt9o2yLG9C3yrg9Nebg3DIFh5Qwsq1i
z+KmZq0xahENXfEQVZNdtl57IY0SEXmzojRDZ4/XOGuT2wANkxsfKdHxqWuB
nq2iYPbTmE3TO6CaYJz0LL2Pq9RqKusk+0vAu+3BMnEc+A/OP7lPyWGYYrQQ
euKLOVPgWDN/YKykQYd6EXT91YOGAfqqGUC+Mui4wPYPl0CpL9rHreWnAxMy
+2GkijU7P8w7Bq6peGBg9RwG2V0deh+n2RcZ9v3C/0KymwtpTgWuRbqQVtd6
20n3JtiMSXxH+B1Qt/1NXEW/bMYCugRxTirHQBOmVN/KuNpeIUkcx5AMotpA
QJ3S0ti73Ki96iWXrK72SToMO/pRD6Ez0V1dTq53uib+QnZ99o5JPLvB22O7
r/jb1euTz8X32RXvnxhUdLIQaynGrcTk8b5cgt9GdxYXR3iMW4o1WwUOXNte
wUeZIr9hGyhNV9OAjocSwVrhnVu02WQ174qg0vTGDGQZ8dgAn9pgUoBAsSKM
sh+cTAlRYwn5IB/4GCKyldZ8yMMSYWsbSVhy8lhWSZggfmCENY3T0A61vqQf
9SZLeaipk+4crV6di5YcvZD8LMqR8rjQAl+q8R/B+/iitATgmvlfZ75IHZg7
9cAmOXunPurq/9uOA4VfjzqoZenv43qimJEjwwgQ0upQNv1nJxKc57+AJEgQ
QJM2RRJRXmvEBw9dGLiU9NMKQyDGePKPnwoGIDg4yUZ6pHeT6vJqxDK5SZRC
xTPTO2qhus/raeoDeJ78wpto0WuCWcuhapn0yi4te8BSYdPjlk0U+/6APw3h
eOqA5SrxjMREAy1SCcoNu1Sflwmd5GzBEabK7DZ3cpwf8zp/rF8r+OVDR1dR
xIxKFdX9eGB/XlCzQKnyU66jXYv1kOqZ9F/5kZDlB+Y7j9WyBthxx4/taamP
s4sqRUj8M5OmcSeXE6BNAtxLyqscQPVsnGnpEGV3s8OSBSF7oz33EZLv7v/t
s0yvso6UoZM8txjoxLCGgjaQmT/PEyekM8f8chOGTuxDyagPv+zDq+9dZdJ8
mydmsVDOzxU5hLJn8qjp0D8syjsGTB4xYzQyBmsSLle7zpXyouoqic+XYXYY
DgCUry8ETrM79CUsVp/eYf2dk9nijfMGl+YOuXbMHERbcs8+hPnUQDuz3rl0
ljfFtpbDZCpHjPFYkMbAYBNKdH0R554r4u25oLUvcYB0pZTf7dW/25nqpysb
Gm0puBMxD2VA40JuRlTfb2LnCIgicdATh8Rbl7nTYKaGWtG3t6UXe4USr0bp
ZVKrIpq9Jq5J94CBAYDjLumKIslPv3LHJZOXlIXzquhUkp+7Fqu+l8CoKhG5
7UEp5Qy//POPD31KUL7jAVYzKic1Iy6PdB2wwlf5r9L0zlMUN5rtuOf2FOik
hroJfJVeMyq7t8f9Elj9mtsJR45zlWsojihGqUY+OFlnRWMiKlJbX8PZaMtZ
KbskL3+eCUxFYCiizj+G+b1JQXHX6uJR6jzXkv6qCdcy0u6xW6heypy/UzJF
VF0KRR/7uPB+1tyVfNHvGAUXkOc5cn6AMq1d6W4pcFcgHgR6kGc4xsDdCjJw
wVKAJJeUDHJwgaibjDRE+NU7uw+ydiIaQluK6iXKJRi6T48BlvUqP4Mjidmo
fXLPhiQlokQd39XOe+0HMn/x+xnazleLx7eI4QwCmJ12gpODQb0wfrZV/EtD
WIEXb7+Ui4m4BfbtHNwrdoYrQ3y0TvOVdiDqNLAXjshtaKLXkrwK0prg1sRW
SdrFzCwz82hpDxWuhBgrixvvY0k72jQQYdLC8gDTA11cj5Lb3cu4mD/3XQ9x
qKK8u/WTYZVoE2RHehsSjqDDRiiu7fVa28OJ3PX9Xyh4MyF9396GQoHjuCBH
gle57HcMKG28/x8aVLyy2r4UypJRP6Hw693bjNtDYoaGpZ/RLqQTLOxsKiby
RjJMy1Px/4zk0PE8NLO+Q0beQAlHdWwOCDPmHNWkxrg8wI5lEn0SMTofJxBw
KjlGwpjDz0wvGVdvbzkuOlzacM6ROnpKOy4IZsEKOGHUd8HJBIzdkvgJpkep
N12tKtX9quUZtWshKDBLGN/XdALddPkrhNLCtQaZI/6Kgs+CAOH67muWrRzD
DXTw6Dd4J2NtBR5PMQx4UAQtgWJw0OPUrAFOqIZWEpbVTQXK/qmLwsw0DZem
YPyvuPbj9Vp8DuXdygf1bHLiPx+zWaEvzAeisTgTrqmBVtVGYmxc8NhMHIb2
cBevcv3LTcBbA1GN4lP5jQAHYZ/qDGzSssdNH0QWCzxJfwOffv+CLCXZMMeF
KvY3f5iy6rHIawlMfO/zX3iUc4g4Bkc51SeGlii3+8mmNCmIm3KAOu23ihkL
p0BiCcqHk2hn5ys/eQt+mwgcsPGbfaq5KS6JbnX7+uuZ40MDNxNAOFmqBck4
1AZUOzJEn5nkPeufFv5ARJU+n7qfSOj8Chnl8UKb+DxH+vacW+XoVDhjb/uv
VaDKwasezmvx4ERRrohYnEG06lhSL2HNa890DXR2NkYr3xPgsBazQfi4+ZXE
ezAZfTkpYIuIyxg4iBtw8hzyMeGoWTZjs6ewMdmnOSdXlRpym4xA1Y1BWbPX
mxq6Qx3YU5+hLUYv/BzoT/g85w2sK7D6CHD3kqwjqprYPgZDAcD2y6PYYv3Y
a+5MtiG1z6khaJj+fCyph9i5EKQavcM0i6yhiPHRKHxDDdCrBltUp5IGi8Px
l1SO/mAJw/QG9SAIh15u6j0u12zCuYWI/E2CfenYSHfOGIOiefHE/F2rSZiE
FXTa2NfSoDckIPhBh9nobaeS7bw+N1u9Su+KB4untl4lhkQxjE6Yp4QWfH6g
mfQivf5fagFNnisp54rW538KlcXxL9waDSUy/rFW++Gsdug0xCf0Ab4w6qEc
c4N4ABCbEo3yYn99OD8EJsN2VjcKTB+COKDbqqzhMLoAelTOlVgM0RNR5WQv
2BhSgsqkFfWHd8VSH8G+3NiUK8C5Pqz4oCUWtydpfnUlLMLiusxaZVNVPBHR
Qx2u8EQiq1GnZcE7gudLYMNXmazGYqfJ9QSZg6C+rdx0Q+JQVsAAsGgpCJ+L
AeIqLIzrPC9kzy04sIa5Doj0RwD7XsWasLA8KlGDXoJUtERJEgZaNU1jhvWe
dT4FF0M3h4OdfLJMGf4wXvjVqLlYLYpNPazVGREbJ5EAnE6y762q45iaYgRK
Bg/hAmopR4Ju26SvRd+kmmzwnYzCBwfEGTQhNOdINse1OtW8us11ADEQQqQ+
eTRMsh27U6L0reUZWVJEDY+uCRL0qJ6MMDsuJDqXRWrrPDDqBI3QDqfRbenr
mHskHXHOQY4rXx5gKZUDuG5YQzeUcvBHpphXEoeQUqP2yEBpA09ytpb/SKEy
Q8h66Lf8PoSQqL+YiCSJJ1I9jxtLyl2hb3E90qeEcv0QkyZN4ztSbICVfc2Y
YfxSh3C1fDjN+H58Zs3dBWPXuSdlCD5uBTS8PHtQjTCHTvd+SbAB7LBgkq3O
Bu39jkMp+4SPNeiY6vyzFxnKJXc7s3GS3xeibRUIjYqWUBEjg3dON0XnTmCs
TOPyfXv2HJgLS3W3+K9aA045cqg4aSe/3NpNNktiALA5IwbtFD9609hXX96r
kvNcna7D9HHp0O/PP9O/0/CZbalSD2+zZg3Nvbm1yXuHuCMSrX84bkOXF6Q4
FA0Wpsqji5kYDCa4tavmxP5lB/yZdwStNkGvymZKWMTaxvx3kPiMZuZREkKj
TYbYGLtPf6API+696HCPSLn6OC1e78tFZZud4P4rFaoito0lsv76nZ5GOPS4
NOHqeikgIc4jAH9J5KUSfKUHr/G8hxVzjQjuedUj9SsW/fuiBZpWQI8dJnek
vj3QBDSydBIx1s+adGXc1pBzb0Yp3GSylogRYR08C0wytB8oci4hONxo4kdC
9ekLSbvQalOXg6G1PUSPHeslBWASiAtGaHGQScJ7GeGjrUAMLI9FnhE6OGLP
Al/DX/5G22Ghr9dxBL5Qf0fsjk1wH8x1kmt3nRbjOh62SiHfn++BuoTxw+6F
pfweXn81CKyWfXsQBF/OVnUNdH3uiVk8Y+fVuReeIEYU03cSv0Z2Upu1Rxdh
I01jXFRTUKWjsHZDWF2m6H4mk1nJC2agOXXcnkNu0cXy3DGo8YMt3BXfgumh
/N3rSw5bUB5bGFcm6a50Gg2klkKj7omQAuYIu7FjQ24gnCcbfaFaeWeeJwnC
FqG8oeQ54ApVNpe2cwT1DRV8MfAVjofpeaKu08NjR46WkDXYyGq0kpAGY37S
Q4qq/a6SRfWlm/DGVlyEMY1RSayTCD8EDfpdnem6m39u2tMlzrD/z1p1O5RT
kBVxuAfr5jNzIQqq5kSIuAzxQQfU46eHm6lHBjZ+RD5QdZDiTP+ibAdxmn/3
KgTAX0UIvrftIBKCLfMKhdCVTWMUIOSa/Dsd+Svov/mgYNOEWE2V8cIR8TkZ
zIeIo60aw9X1M3eD09hFGVS9BOpl58GTqQTiQWFXr32ZLff5K6WmUwoTq5JM
GstUYIWZqGXyhfyEpgshFa5dNmjDmTO0juEZJ1w0GEOlbf1E8dtGRvDo08Mk
jwY0SSl0zkqEpJruZWTflv3BE1yvDSAhJOmmOAHsPAKLY6y8fOmv0RYp680J
sJeRfDocPGm6Vm5tf1dDQr3kxtURH9PKF6y7IbYyVWFlu/MhnibWxyVS7ln6
B3Zymy1CjP4w2m3mE9zxfHpNJmrfPF21FF6M8molk63QTWsqo4RuH+ktpnHZ
7xJfW7BhfHHTTd1xchS+8/rPntXk6qRnDuNoxxKh0mM6rbxurhxIcK7MhAJa
BoChA1O+89Rr/7lrlfX2NuCfuv2vmuBQ5XYjJDvFvmrxTpMULKfgEyabWRhz
tFaB75/P4QdyXanyY0XUoloIbGzAt4T23xrSCCcKtkEqiwHe1Q6nxgKFD8FE
t4TnSx03JceWCfc1MwkvwB6xL2AXeNz+S01OCBE4/IqWMHPzjQLN8yBNYxyN
/WfVyPcZWkM34kZ6Xf2GpbBktjGvceyJlmHbIQGhxuNAnuiu2KCFjpePZwZT
/JZ0tflHhbqmMYo4eQqQ3seQ3LKKa4/uwYivJq5zzsxXj+fQvv67BEP0qpGR
flIDsQF8kwCpYFlHQX6I6v0eSQ7WDNlXvHtfyXjrNUP7U+L7Ak201vd/dqPy
QK3SpTHrCRl5PlYvV5oPHbQA14x9Aj6brsmx8ieYRm/yzm7q2evL/Haj+Mcr
GrjcVjpY1la5agqQ/D4U2K3B0SJabY0EEcYLbZxhp+CxV56P3YTMyCDVE4/0
Z6HErCWKRSsvuzr/U6EixiLoPmxnUta+/w4DiprPkIN6c0hZSA2ED0qBQ1/t
xE5w9GT1oqZvgJ3FCA26D/GvGJKLwvekWYvb+24GbXEecwa7vr7HNmUJn6/K
Jod+zRcAN74CCSN/hJDL2ew177fhr+ZjESxgwPaN7y4wEnFffW2CjIjQzy8F
toDtWv0OjHrC8gyzXGqGv9S43w6xFAUTHaVnarPW3K9KdA/a4BhZR9MBIMkr
xk0EGnZAIq+9vF19f8IvifYBGj3vNobwOyRHx5Z55N87aD3bFPGK+KNz/p5Z
NXa8LOSXFxU6s+Dy5e9PintOScC80NVRjOLq7OwDe59A3XRBPzSuJZdPmrrr
y2tmQfDa5c5GMU+apBhV15d8Rnlj25jR3+ehipoivM7g/MsDO0lisFDnmltA
oNuMtb7ZDFXVv6aWTIXC2+0pCtjly7f0KzV9ZtZQ0roPmb2PLMiahS0zSXba
CPqOHiUZi7uHy3GYxL80SiN7qd4TaEO52ZiX2Lu86NKvLXZWuC6NpzPK8mi2
mbTH2PDWxkDcB05EfU8TF+maoxlsdLJ1wc3l71mE5aFlk5JzI6ZSx0sk0qTx
Cu8e2oJZq2yMdf7OlOp7NH0ivh7ZWghRDwdaKZ0NOp8pVLA4HV2JP4LqrTvc
LDcnG1knHf+R8AKa2rU3CwCFoQ9pRCJlaD173d5vyFcP12Ic62mC+M1UM7vm
IehQjVXLOWcMDGXhHN7AXa3QK+SMGr+ulk1jRSpE2AQIVQsfNjvrN8eOURA6
nthd9L841B22PcMbM1MlNK7cwQtHLihqFq2zKQHFdx8EpPqfRhVxdlAf4cZi
5KrXoRZ7Z/EEDo9waeqhifdslSrdNGS4ZABtpwJUaYvPn11fzD/zkNmbkWf+
Uf4ZSyG8cnxJLmA4ekahBPeQ2q6P8pgGFUvakRtMBoPjy8sRg56RiQ8P+w0z
ZPk8i8GGx+fwsvwYCtNakNlemCSJiMZNcdCrUxliYmkFLVWiXkosb6DfRxGO
/zAx97h3tiY8EfFnqxa9zenZeBczYNeY+5DdhkIaE5dlhZizR4G4G4sb67oj
wpZ6PFRu+hovQu5/Dz+MU3aDUqxVrL2ca8rMU69eczrBRSvbQ98yQ9SNI7yu
6xkH3DyW1IIHNnffWMU/HrjhWpv6le+hhcrc9+RmyPxa935+mxh/XA4ebx7Y
24EAzwHTPRIpgZwpM3BRsHGAJQRcepUXe7qG/0h3qraGVJY8WJkG4fwSviWb
HZ7FPP9gsBKry4k8l6Iu0gUUigCpjvzR1cbT0ETqBxBjAnbUnqca194SoN7y
4fcRqKTVPvs3auMRe8GtgTXbz8aZg2VhMFClfHUbegPY3SjA4UWtRahxrRPb
Y+SluuriLJ3px7YM7/FGG/PAIN6oS71x+jcrLw75bo0fJ9E0Dyy82SR6nps+
2zzPxq2HFcgippzWwssGrBTDVTnpbMH4WGtE+C57n9a3WgKOj4cdE6PbgpR5
KneC77FITH4TSsiMwS6nUp2DmHVUWUyjoHIQxbNw7bTxZLhCppUCkl64E3MX
bnLHh3RV+vRkcTh0Bs803TNNMRI427RUhtbEUphKxycUXUuSCt5NeDQEPzI4
uU7BEa8PiMGitcdOKN2C00WLhJa8DGpvGsIPRGrS1DIkX8BHmz4+xMwui4/7
6ynqDMeOukszpNydnxqwAIq/wfQHuOKh1Ds9wixophNgnUACkdUylafphZ2/
TzDivtq5rl6UX4Kz2CWCf0oyQIDfHkLVAs2EXMvT5R4H7C9IUBjb4rH/U6ij
fpRclOJS7g0MdBXh48PgoYOWNAoo7stKqS2SO2jvbVvIOOlGrrx+d/ZAPH4H
VAbBpX5D4RJJ0BK2jc2M6CUVT+5NtX86WWnybaRp/p8gpFZhHzo3Yxokwa+E
zDa+TcaBzMJSha9nXY1VSfRAgWjvQNgR3b1UcDVLHYTc9zxOeqxKgVmPib/Y
TtRTKXHaL7jUz5AvH5zfUp8hxjWlIF2g2sv9mEnzJkCvzCAmeJWQabkWtsnK
Cskzh5sAzj8yPzyHH9vjIcG7fb9lyoLfKGLfxqhZvyCm5IlEJXCGU8aG6GCD
UgDwmHiVkhjuAihuwaC/SQp7wP5ygQuSE14Eg+/vHQWWYe1p9bgtXktj26Rv
of9wkk/N8aNGh5pbjWw0IfTRa3dRsyoXnmy1InPdIJguoyCc5lkrqTxje20d
ZM4TbZAzWKuGrq7B+Gz1n2MduFCWyLt8H4TZCDKGZezWYRpWPUX/0+eU5Py/
kpizFjca3zghyAnHbgq+2+5HwyP7r3utNU4/vVB+Vi0RaD55ct+2tS2HoArD
tsgDwCUFAKQ9n2AlpIwDNkowu1nafunNuPxH3I3llAmDh9fO3kvj2auBapFA
djJzPL85GMMhg+VllGGVQ3EwFYXAC2Jw6/u2UMXf/OBQSoIvxoUkqiYxyg8F
v6VAFZuyPdbQ2pFfVU6LaslNS1slVfxBy/x73KWxa0UwJKsu1lk/NLhGqJPu
1suMvE4Fwtu1HDtGPNcVgRxLu4joLa5jvXogSo7NryKtLmB6cqrig5cvqYMb
W3H1KMy5WmMzmRVDotUdjonQvaWv04vRIlblvN2hNfDZkFeG4NwqEPa7bTHW
2CZasj/lff8/qvkFyKkTbgpnYeuxTUpc/N0BNn0pnL+3DAemUJPZ0k/CoxQS
mVvywRF/CTguWkUTTtqt9dEvuzYofLoSZdKXaQKFxSbgQ6mE1hkaAcQII7Xc
dI7bVQ/LsVSg/hh9T0xvkezI+TEhoiA/scT8wvN73MZzquT3GfgBnnSpAnTU
XCrNHZz1/FQd5KABhV5kSutebjFS5OIYB7mwS8aHwb9286uL1eTvq0glcBH4
+mlH/M4+gn525oxiXiaO/QcMPDc+YyEyUrJFyFo2x4WDB3Os2p6Fwei1KAVQ
4k3NYNg00AN84udSX00c8SM7lW/UpUI+WHN0aPsckHAA7Zeuwvw7zj5a1WGR
FJWOF6v1CmgsYNqj1XkMWrnRCWwCZkyMMD0rjA8wv8slUu/aULw1YYNVPeNM
XNUyZKIXDtwDtHSHkoOFMmD/MKBC7H7PvACqney5c8HBCIvZh/fXPH9ekv5i
ETrJOK4z4W2pbUAVQYG2/4AgzI/tLRB9FBGlIAbh7rHHPfEWxcMMWKgxjNkf
cWPVMAt7dhzznozKdjvXhn52jZtUdlfQcWpCliV1dU9lM38362QCXJW/qG3C
3IVeYOvFN4G34d6XV18Qfl9+KjKxyHYyNxXZKibiJ8+S9Wpsnj4XdGyQvCKN
9UeF8KwA2lKrh5ldmHL9zhBYUAAPJmkiAipVOhQQbvVXrBIBnwlOjnMtI2ol
PX9CJRzGvODoDShfzms9AOqwz2gMuMebfSXjH+Sp5UuFVbP0UQBwgS5vFOrg
9haIUR0c3YBjDrDXXlSAWeYfmqRVpDOLhQsRli1HijHh+9L5/ZUyl6kllze2
xUYOZ891z0eRDIhHDI813bwWfRii7KdofubCSylkbaTTfAFvanSP9gsBuxxt
SeKFIHJAzyTOSTc3kWR3ifLLHUK8KtsXuStjSYwQfONiWqNxKX8Fttu1Oxtm
xRMs1cgbsLpzWdwWYh/H00mnqpwMz1DilHPzaCpNlULtt5neoCIGAzh09uAk
6r4Et73LfdvVs+e7pEhMVKhndv90eZdjsvPTWYDluFq+4mtcqPt11eXECbjO
56NzjJONFkg1IMFQgpB4ySCUVy/vgfepXplFQVTh6xPeXcWZCH6PQ19Zk+Qa
9Vj1Hc589KoyRz3S6qHfHtUDEiM6ubULD6GES9J1JNQLJqBLqhR5PieETyBe
NAOow6OsJ3pqE3JDDfzc/8d0p/7s76NTABEti/RUsH0EAEkpCDHULFcMtVeL
CcsijEFB0/+3qIBunnwWcSTqXQfzLSCAFN2DQx8L0TNzEiUwvV5GB83iNq1o
uMWkiXl9udTnd0IBPDYqLMOP/4QFHAuXNPStcFXEFFVQyUVy746aoEztW0zY
NM2ZWxWfkO9ZuzKHCFq00vMJEZ7Ad9aLZ2xpaRatwBkEUIjqN7v5MmpxVRa/
6NorVMMNMA4g0DAljFENbA48YVR3d31IVSvK2ROqMRMbxHNwuv6dbH1mczsP
denuCKFdj5K6I01APs7pT079b8/s0Tv74OrczmhQIHIiOd+L9/ECbde4qqCD
wny526hLL/aLYkNhFbEoYAf7Ffo/8ADRi/54QwdbQ01THI6qPFc2xKMnrtah
GnTaR97RFzhOWNxS/aFT14h3e+Z+wuQg7pRpRF4QtCznulWulUFf6NZWIBF6
xg/2ijfD7OxFEp8bvvLbZU00fbyM6Es+uxtCB0JklLqrnphSE9XwqYqAPAwC
3xYUsGWyS4iQf5/hsnIH2doj91CG5S7C74ptnr6hLE7MFkzmp4NUFa244fwv
l4kEpE857rOCeaYu89h3NFZnxd/5YgqnDB/cxa9yHkKEhBziVkodzApuSsGs
REPr2RgkfYUEEvQ1vrWfca9JFrJE/7IE54ELScSw8Jh0Y/Gfa74waJHW8lfJ
SeUC3aw45C6swEapToEDeDY/L6zvL5+Rl7QC2yhfNNkQYN37zJMyqLjNXDkw
8OQ8FRoos0QaeVgMoMFKz6roq/HOkvpnWv2Kx6xrXJEzafYwMGmrZGvxoIHa
UzXBKfpTzndSEr2KMC8VXdP7LWxihy6TozvUe9OOuEaUdHU3MesA2LGUt15i
qQSddITBfLxpKzpWMl33FVySnt2wncEaOaMGfpmmGuFG5+5rJ9QqB5/9/gph
pMlyw3VEiUOQAbELFNk7i2voNehdS6d9zblpN95wuSGPRz7SiXzzZfQYmAts
2KNBHWiDEt1KFtEjKb5VjzMzNCWuJyN2fSuFnXTzzRcfLWfPbZei5s+1dktq
3SZQJzTWtnFQdHuJkMgA6qaV/bqUyKXCB3wxCe9/scAd3EbzqzTZquY0bB9z
JxuW+SnNz/M8E/bc7hvJickW5Z/FmoOdwT6vRqJligajur+zLznY3tl4TQiU
Ck969KNSGdIm9sWebghftkBD+r5EB8/GYtCYgZulhaZJGTq+qf/hf9vqzcVH
8FdK1DwEYPs82ZhsforNBc+PuyYiY4ep9roCGcN1b/QVSVEF8iJbF4sAtZ45
WGQgoI5/NJX+/YEaz+wr2qm0w23oTEPz92QJJIKs/WFghxAgEjFNIoOe/T/5
dh4KPWeA6+jS9WD6br8FD+uHXa9XqlBJpLy2skdEVgg2o8ehinAJ1/bQpolQ
EO9sl3AedXdR8XYdH4kuKT0wR+TAl4561ixZkVUH7DOGyGTQOa3gOwoh5rOi
cELNbwo1BgGt9yscJh2iT4bTXgQYHgGHuf+4VfJkTo8QGU3W51tyZAsmnQWy
h0HMPTCdtETp748u8+36VCF0i+dAPxa+98FYIJqI0buwhYTUSbyWt6ffSoWx
m8B+v3CMA2yB8ZhWmomYlgPC7P8nDyoL2AdlgOVgEEz6MlzJDm1A7A+wiRQk
npC5OHVqwFrVBPg/XhbTOOKI2+LPr13tp8tSNbyNxpYO7B6QANJkefSVnGlr
+DE3tuhWChSMWYMma/l3eAcous1zC3cIgAJubdi8rJ8l04kyqzFYvu5gE1ka
vaWZiqJoa0Gh1mpbvkGAiBHWOB864Zaq5W/TgIfz8vXIVvptgbBMrGkD42D8
oQZGHUBzbN3bPt6YPjTx3xhHKIQmemibwN7CA6ZcdLmmqvMNbGzqQ/imlXRg
5hn+07it03H+idMeGjdmer3QTimiBjD1+oQovcVGGwDFLCNNlrTL3BG5IDac
/xsWB28fNelgFGtM+pgtqAC7oO2MW7hblXQWP2/kXL4Nn5YpMifhcQtyGNjE
fzvNDQuph1r1o+62Zer4zboq8MwhQYiax9fKmD3Yxh3m0z2eOCElWEUV8TdG
9GMsUuXZ1/ebnpwEUAiG3o3x7VUKZ4WC7ZHw4S4dqaEUi/9O9a36NUKRHVmr
CG6hHWi0dYAs7V3HnAOf9loyeqWr8/cLoiMpTCB4OeioyGsnsRYMfytJnttx
GnIUjI8rxioLRsCrfqN+mHHpz0ucgryp5yWzxVXTNV2ZokxqH+Umu4slH7jo
oIwawbPHF7ZVAqb5OO+tZ/UY8PaiMftO3lcxyqp4UVh94ED9O3eDix134PNe
ySiNTGOrlCkiCVD0taFpzvhgG2FAdlTFqAHS0Y/RYLFyQc1ZA4tyGSQeeagB
Kpjf3ca+7l8Nvi3sYCNWTUxT2lwFR04yBJPBGvPytSO+9+TzDM8fhVIjUw/X
LT6W1kkl/krHbNyP/hV4rrne40YCn1hyPKKZqJf8KRNq8KkB3OKIRPXOY4FB
TyklkKpfZXI0aQrP8swfNmGako1vFbDoFHN+6jTWkSk8f9p8ejlapcG0E8UH
aQWQCMbulxeL4o4f/xOwBZv/sc2VSTUhPtmgdJtRmTEBxnguMwqvzs33yths
5Tg66KWK45RNH191MtsejuykM6KyQ7Kk7I8LplLurYn5cRuo34rqovlYLbVF
U0APlO4pawmbG+EvzLR8QGq+gTb2ZpnALXuUv5wmiqB5zy7an8pi25rIk0BT
PPHcTMajrp6S6FbrKW0gzFXzvbEBS6c8lDRTum5AiZdy1kgHP1OVSic1/hIK
wCTDReGvR3lj9up4nhoNjWAI+XrZuQeHR2nlTT9ELowoxQFRBipMgzijv2wv
RZpAfMFLuV9AOtuWVSTocE3dVERJqsa6PBiDB8Fo37yRizwFSlfKf0OpbnDs
eNb1LynPg9SCrB8Txs13GhCWdmDSMrY3GnGyIb+xNsYMPbUAGzHOrm1U7PL4
cQk+lKpDOA6vXQc2EI2SMCVdl6qi0HB/Xv2CZcA5iD05u8PI5a9rgCy9imQS
dPkpPHrHLUObmSCf/UmATBsdG3vXQj7pYwLMy5M/srW9xIj4doVCgQb1c6vj
K3nHEc6xH+UtznVcSWHHpcMFAKBmZt/bMhfHusvB+cPJYe+AftvckJh8XFCm
1KrR8peGGxQCGvWblIPA1z2Jo1Uq7i5sCwoW6YtD/couirqtqNNoUyH3FJLw
iOYUQxby4UHTTfxwiwBhZv+Q+r34xZ0fLWCo2tTqZD6Mhl13hC13XcU9+AY8
OXWznjlQ1AochZ19EoKDzv+3CGCQGc/e+G5uxf75oGrMwb1kXu+eZ8lPeAcs
gN2zyg2mcu7zShlYz9lhG0qvvD/FXQF0nO/eHdkxnm5Hj9UdkPajh1G+cQZq
tofX0yk4tqEKAbNNh2x3MXOXt43Fqcjo8zbjCUJuukYyNElweIypphKFr6GH
pYUOkoN1t8dB2/WvyekdSyKIx1SZXubGtXK1G8/j9FjwYEOU6ReLTFAtq9IN
we/57dQ3ksuoqL/scAaABvrA/vtUH3s/ACcwIN5+TECPNAPwuYqWb5/Pia0q
S9PFVb93vP/IJs16A3Sy0B1GbUvL+OQUgGvxV44DcWubNPMlEkMdKgds2wI7
0daVCfKJsEbj1fQ5OVDIZKQA6r/PXO+ZdWNvBL68ZNkZGJgA/McPD7/GxGQz
cyJw+eeCsI8aFehJrmXRcIdt+lnpia26l2vPHOh8z5sP1O+bjc4xBsZLGNj+
kF0hbjDeengHgW07/Q+i02PoeJh40b/f9orYW8RFcTEJ0hvhcMM6SWTDNstt
A8t9nxaylQvuGRE6YpCvBbezWv9jLR+e8odTYSVld2MyabjgMirJ0+JfUV5v
V2UTE70Kojxu/tIS1MgbO49Flc6gL8QMAkHBS9GaVo5O7kUJg05/BiFgWTHV
rvdMpn99F8zSQUKiRroUPrUuVKVSse6HASlniZ8ufExubF4r9ObmW7J6vRKE
vHaPOXPYcuzP+N4RiZ2gCXHuaYYLovIxJJD07/c068+rHJqmfS0SvXtb+soN
gPOUDQMnRA+/kPXgNTw1Xf5YvkI03WjVIuV0g5cNhN6AQsEBebav2VuaL/+8
l9Ej8YND0wzMl02nTM1StXodpGx0KUMwcQEWGIuczVNMHlTz72UoyKGQN6tz
ASVAzXf0oiObzkD+CudQ4WjPUhq24+GJH/KwTg3CnXbkjN+Po1euhRCFQhDm
wezchfFQLgMUeju8jl+MGcfm9rrUFNZR5lX57RC7OgwDlmIFWt3GZpSj4vJO
NWHZI2ewopx+hSCkq8aB7ob7g9XX+92hEYSQ4VuGG97RoGKAkHkPIPYCRosc
O811P0IZLZTYleKR6kOJC/Y8NLVxpUQzAbiQr1v881WKsALktIEjYBL9n5LF
UplHGKP7p+LH0FeAhXhP7uUL4Ulh0AfV/yaxDvWGbhkR2jmmSDcNAcXU3coq
c4n3l3kCJjDVOn2VMOaIkZWQ9tiAvrdMSCTNl0nk1Ysl1/4e2fyb/PQrp2zn
pM3a96xYxgFZFeC4RtLV5aQbsuJoHSyQN421sDTjOwf+ecTu4tXJyTc+51ti
P+LfLW3PozXQwaPkBWFnaia8QpDDxEiPpFEZ8aQNWNl34Au8pYRh+ZHrdibG
wCuovDAakEFmZYqclBscn1iD/+DWXRqBfRQQ22wR3kNYfxX9p3k+4Gn3HI64
lq24WcInPy5521jaJO7za9bbKbjISZP2lC2RUgKRSR9Tz6dFcJJ8INI8MW+P
EBS/MyE2EpkRyE9L4W5x7Bo8yC6zB0PW8vsGDmbU5xKdUVO1XE0v7blTV40d
tcmQ1sqPPHdWBw72L/UkjQ2BDB96i9z9RhJPTjaV20PMX/NAbI/UJZAacb+Q
JWz3wS+cnI40vZuuwZ+qUAf0eHhqhZDPco7qZVQRJ2DpkzPfLNZXjqxVzim+
/thHF1q1d+xc/TbUgDGNODDgSv7abawY9E3m/F/NkiqocpTY+P/W8DafA5cs
qmF4SdK15yuJe0seZTYHWz63v5NuFPWfA6bZwHzW3XSbqQRRygK/Cygp4+YA
v+UH2qBUkzK85hGTnDCRBDWQkHZuYKIOVNlbi9CRYfWWRNSubYzRXwNcm//O
j9HUBeDoHjBiqyraUmpqWoMZHFzp01qq+EXPUkKLoDpz1x875h10Y9TCpHvy
xOpcnA0C6R5QwA604axn845ER+gCfXxYBSDuEP7gdnxEOMRt9hx9eXzOOcih
NzkKnjzVGs2jCl3694Ky8H+ifY0R6CVFR2yrgRibhRrUjeojng2hTJYrRlX2
9QiV1BRt2tjZPktFQrUNCCPqBnOSTjDobU52aexCE+wbpL4aby9xt4S/f6TQ
l5jMr1ga4QOvZ54dc2t27/I0tr0GFiJU/XHc/0Rv1yrPeDpsLY0o7JBhgAGT
ucszNPbYkAxAVzq6+v8KVJ2PB88bwzpBbKSvQpTYEWtH06dx8PzKRmx8Ad1b
WAK/ZJqDNvDbqi+igZ8Y/Jvas/S6rfhrfAXssr+qWKND+aRwraydClPKpFnv
/VwKicEyFqsREUXznrII1lDYOWLPyB+exfU27ARMVVeZEIHq0ToYkqUcqgii
aTuZlmKTl3lnocFKbNsXSgXy4i0AmqfNXiJc0eY2MceyMeyF41by7bgw28VX
Y+ceLnJS49J4vfAMh0mZDMj4cWW2Zx9i3fAIrtU11FQMB8RKJpWJsPDfyH3a
GbDnMtye+PwIe3/knT0Ab6eUsRtD2HfFiqO9MYf64KDEhKBMwlIIs0wmWsao
PIgVoMTIBztjxfpTq8aTT/YqSVLl0+wL3qVVyoJbkOD+QzSvdTT0KKcy5CxE
/abk0iQ1afKi8ZbfHfur+JxY+4F2N17svoDFr8ORc/KGf0Q0QcwhkuzAK05t
2lx3SNGmPCBVr+jZzfdwYbeF6FFZE7xEQHDn7d2k+a0CEp6NXG22UdSzxcnI
bhu10Ax027gVAOR4jYhS39M8Cs5zHDXzT0ooXY3OsGCyIms+s+QTQZHpHnTz
dBng5ld9mBgtCXyS0+WP70efhQEI592HpJv2ZXy5UVQqlemfHHi9gsezh7H5
NtUrZ+/VLwdZ89a83FqgtzGTI9L/sLBluYeYj7FpGwrJnJsENff24rUbtbJ0
FmJkjHsA1qo2vMc7fdzHLQ3FnillEddHN0REM+7VlsI3EQAHNQYL4woxR1j8
oKet18tpS854X0SLsd6FjPrmj76JnBzUNo6UKQq29Yzv2nFhFEDp1ii44m2c
BfkyK52QDyQurpxZ7jbsRoZ3lHJl0vPtEbsweFSf/s774HVZL9oS1faW+gjH
BuAfW1aYXHN3WpPCE2VuvnxyZOcWRZVUyHFA3C40L5fz/CnbGYQuYKG8k1HL
Y4ZwQL7nOhk4vIbyGxsL19CAMjRAlpbVLO2U677Rw9JkOEam61twlflacsf7
6YR0uOxkRQ3qVzNfz3e4QEnvNvSFg/h9WrKfnwUoVpsFUN4Rq/ZeZrb1y1ti
5+VFxY2AvIRpwX8HGYAB0yF27AS2LvO5E7n9BdppeKVYojLbQRoiPsbJ5uXO
uZ7nat3cp6bGeyQXy0X6fPkIFKd/po2wpTnWdVLfNRRJ1kfmHzWNhabTGuoo
FqdI9nqNZYVEalPpXzxCwKhEj1OYk9P7harWO+ltGBzJn2IBYl2sySE8G4AH
85qrYitGkkyoSMXvK+3JI1FFae3cTc2anoarxbKzuxxxxSu12HW3CkLe5YTd
hNw8mOlpmzOdYOpPuS6Z1cypEtyW4SGWeFFuo8pP+pEPuVZXoiOREI9L5K3N
INjSosdImPeGtZGfavG/wWzUT2zX30GnIoC9Lig2ABjaANnvJL1yB1CnaaFL
kxyxM89g/Lohz70HXIKX59x55QWEf4iBH7maJv4iPVAQSsakg5Ar79J5qqoT
DKoXNR2woywcqxMAFxuSCKsxHXXv2JCFtzKjFSkVsiYIeMhZudsxYEmkNheJ
usCCauNF4dRz88kU8TdRvxMafC0H6Cr3f4WZX+79OyExIZjE8oIE3o9uesBY
40ECP1AteSjEyl92/cFM8yudC6JDbm/+lkpIBTh+2e+4OIkmFtUZlvJ9V7p9
lEvJSEN7axxfwxXULHPsH2KetJbboCPLmaLr6xYXDBxcqX+PwFqk3zsamckX
Gn1GjtH1BdAKjMEzXj0u6FFyY24J+ekU4FaHC7xr6oFr0Qd0i4wfh+pszum0
ONMm8j6VsEFY/K+ZDbpmF7p371HPHSArkRvABSp1rNih1Le/IcY4dyVTs0cy
l65YZxw7WvDnNqRWFoIILYuL8hbVISwoOwX2+o/ICgNQx45sRXn9FQz59QfE
ZGX/lcGPXlhUJrMI6JE3oqO8Xpxqjd+sQOZC9+3jWqFnOEoaNr8vvOZ7GqzL
JHFb7DZenyRiu2gTzv0f/uCMiYg554jU4xnRLoTyMqEQODk7WQICWgiy0iL4
b1CweRspjHamr9VRVIFwE0R4fKu8TtDIrQV2eu1RbCLPGI+RseSs5TJ9JTw+
d2UMlAqy1F48xHum7FYLAueEDz6f8VFDVeAaD7MXY0HeGhxUh/Wnpf0plp5a
LSUHqldnZiPgVZK9Pb5/AFdaa2ErnbiODpJEzA40VJWMOe5fT/WQfl+fbaz3
ASHZ9J7WpkYRRDsh21AzfYwKvuXLBxtIEkqZ9aRhMoVz4vLpU18yFe6bKV++
vGNgfmXcHWIj86Qw9h6ItBiwd7ruySJ3uxm9IAzfGfyi2IR5jQN0xccrvtdE
ExpMEV3OzJghTr0OzBK7+WBShJogxzx8R96USYV1VNssCbIiM78jqjrh5xf2
qc/Y5t0Cyf1UR2Oc/+p4S6TTMnFj0oRfzpJuEq+OQHhZHYNkczkp8JnSzcyz
YdrkEPi+A4mbYlcCqhaL2k0jhefucTFiAnBsZPntF/tR2bToU3ZPKx8vEC5f
qYGdd1b/xIAsGdkW9/J7tiP4k/HPaunkvCLCPqYvUOd2o1QayyFgMrguOSY2
Fq3Y1lw5gPWdEvwXc7c3bti+cue7uM8aDjFpaSSW39VqvBNriwOkzUvHrTQp
kMpTLerMp3bVNTt1Qe4Rf6KOtXgLcMxS/81kC0AzPtxI/apxWwBGoOU/l+BE
CiieHlcOxtFggMBVSMP/yMlMdqJvvkpocPtSSXX84E50bs4s41f8BNHYkYkQ
fFGvXX3fXg1S1T2csAeKHOzCD9nY4sSn2ULlB+PEzs2LDm1SXrSX4e/lLJr4
VWksbvOfFcbwp+8p2ANPa+wPGA4170BcRASQgvBt1VQiQfodMUqEFJsHFR2L
Vau3nvxWAaXhhBl7/azwLVm4aqWrzRCYHRVHJPQN5EFywXJtV2vJsAiIyeFH
wRxJhi3k4Zy8cfd3ZzjJB9JcB3xzQy6VLWHbE24YI42nNp+U7By+78RzJxiS
DFA4/jtQfipsEG4s2cnMnqk/ilOO2IqAUo5iPsRO1AsHVwF9LuaWaE3BALrL
eV/rdqBZAF4I0h7Pbs84sR81nem50ipEdi9ZiR5eqe/koIWVFuZKvMdMQMp9
hjLL6BgKaTnd63Js6L5glA1ThJ3HjSEOPQKx9B3JnONB6ZJkGg+rqBZ7DyVt
3t/n7vuTpmP+MdLZHR/oUBOo3lZswJgHlnZjzWdyV5lyDy5hJGKbf8aECFAe
gAAHl3BMbbmhyMpsACIOxlqFHjT+sfVuxNPUIMkGOAXN3pKIJu1VFXcAkKEO
2BHOrDAaOxn0FS760kq7nQAW528lYK7lom4Zg/nWPeWdYjirAfu8SsLhtxH0
ePcLQ2x0QXlzVY8MFF/oi/AI65ug0D15qD4x5KvR2hQKIi04IX3eG4rl8zeN
6STIPTcQBJWv0T8vQ+fn6z7QmOOUUKs09823fWSaM3LYSy403aJ/TVK0uvTn
AFtki1MDrywUk9UV7kOf1XV5XTdEu/rNQsm7dMbV2zhvk9ILvW++xJXrlrtn
IVOlTXuFAJ2GgyxZgQkVCRM0kTvOkqILjh6dXygq+LUyHpAcppNa4HcXSkam
cCI6TSRDLDu/s9ezcp7mBzQ3p0X+q66G8/haluu5eISTo7eU0I3MnuNYc3JI
sjQ3OA5lhn+LwZg5tdPZzlwN3nwnQQWtu6O26EFS964fSlADfuRcdKvS899Z
UBWPWS+Ac7gvk5EEJ+sgyLc7kWteQ1Of6lhkZVv5pQ3S6TDTQPjeYNk/9IKT
S+wwhtZVTS/pQxgbxBRYBH+BbQjOyad0GnKp8TJu3CUsKFZG6TETDjDUwr8z
NFUmYA3U0fEC2Dbe8kpEZxvsq3wdRi0prEOY8jN39oac4gFo67V2LrQ4AgcB
bsL/P2ONawOL9em/bHXBn/POOhCZiCd8chJSQSi6lA12WaZ6oyRZ+4L/yU2N
xOpww2u0DuT/QSNBvgiOePA5qVC/2I6ss6cTIWVXa1GuHrNGVg7rDodnBVUj
Nn047ycyEjDAyqPJ+XiZKGgY1DwQZE7aKWmMcyv9nNvwXqPOaCD+eihVkFat
TK3MPdabqwnh/oxZ5fEVBAhNIzDdQouTa1EE7IU/3C3v/6YasPAArgNVAQzc
trstCPILPVhY91V6KJv0cjEY0ncZf6TqX+L9dI3nUrml5TLlsY9uiyhlz6FA
Xc/IX0/1x0tkdIwhVdSwUxQvnWPxSbHrfEHY8PmuMRGfXeeGhaIYbf8GlqD+
6d0XMM5+1Q4bFL1LweoA2vbPpLiZuCPFw/kgZaJ75Rz1YEFe7q4i98VFbYuR
RdYnsDwqhX9yi7ITkrmWtG1Rgw6JSr0GEk3d9H+RUpWTRzcFSxlPC1ASxq7G
FMULdB5J5IuBh/J6G3ov5/5ApHgwWowEtH71HCYeX2Vozn1I42nKp10s0I1I
FYNh1/U+HY35lcpWMX5DjLrnXkLON2GF3F1AXVHu1XdqwXv7LdEnAF3tPfRE
T2Oq1OstEQJ/ofDhz5KTVvsqEBd10Dit5mBIWEfqaNUv0uhmMtAwgbeyCvae
/JTSxNmW67QI1NHYyhcxgRv9n3WfgcX2cqJxiNsRsVNBIbB9FfJYD51JmlAp
kaEO+6n5wjrCVaZS4QrDpPs2PCwlO6wWpReDMxG7hRpKllSkAyPDFf3VDLjH
3TDATntDfr1Ro870GGc4QrZiV2E7Oa4LovQvOVPcLoiizOAXGUpgPq4ecdiP
pt9TpwMkEHf5zW+fdr7XA7sVTY19HSfm7WeG2GFbT3mbOGO6ECiJ8CUXNUZf
7RqAD2ng/56lCoMecaDKZ+8z3CIaBJOxBnmb03NeTWqG0w2mZjCavltsUYjZ
nON8GF0kMiJF6sEW7XNY06mlKNRLoOfXQhlUMhJ1BKoYfbW6yRwKQz9NEe9i
SKT62+/tGZMTTGOFECaRc0q4LZ4P+Sj50K/A59FKrznDyTDoKUeHpzwt3GTm
xjjEV9uExH5GY4LGi/wI+ZnRAOE28xQIfB6XfOQJoBuGU7m+iKSoFLeb+PPk
wKupu06nM/p7vSxjrGTo58Gd7Y+7F+WhPDsCXaGFpYwbEggcWuDnbJKD5S60
JMxkSMgSCi/BMUoiBe3Ui0utXrqQFkS9ZTdbUgyBncS6RrHh76hzfknQZ0pO
IrCMpibwQNIeTvPLesAhe+gHD6ODUlLuQSIxMfAtA9E4X+1PiFGfrzfkwPSj
AfMEZnOdGRIDEKd1oI0xtKP72TCAdWlt//sFl8a4pkfwCHjHoZR1339tXNWv
sKqlCIG99ffkxTj+2XYQP5ihqylHf3bxNhKK8pYI1odQDEd+YRE5Nx/Zdw+E
gpV/La4dqFEGQWq//sSJn4GfFcul7p2gV20IXM2H9mKe8MvSHwnDaWcKz1ou
clDISKMsuTIcmQ7ubkSunpFRCTCDrAGkbfq+IMrxgNJ9D5WtZOkpRqtD0gT8
FGn+Q0b8OG3xaECVL9cCKUcNoFmtWUmpYJ+s2hicfAIhjWOvegFA1EbG4tyt
WeZUiigKXNnMUGfNEVqnEAzlA2JLEzG0BrxVf00ukqrgJ7Fi51gJC6UMjG66
R9WYqudMjoKqK4eFY7PXUPEPfoun5H1yKrofrIuVT1dbqWvBBtQf67YeCjAu
1E2wchKCqHb+UgIbpyzzQ8ai4gSajDwIjXEmk3+JINnJbArn5onfr/ocAu2R
W822paYGNY3u2+1EEweadpNqi9UATsJNGE1LamAA/S3pYrCLkVWiYgN9ZVgl
SrMj6c7ztBCFB4kiYs4DMtdpZnaOALE+8/8YWwizm8bwUwNhDkmYCEmqeHEx
I/t+sHDPk/fx3RDBGS6y7gwAy8nDe8U7uSmbqk4DWB90M2wVwbiALiKtAMwo
o/S9cUrCGghhc6+ynydS0F0Shs0RjlwUaEktweDe95q9luA4M1FLeKioNCqA
bAS+RweJQapbRgNzv6L4TCct5YD+/+U9gCN8TfHhQVNmAhsapyvbDb3HG1Ft
TKwk9VFjsfdbHN2+wql3YVxxdzPTnv9TcdE6lRTI8Vsc/soN8JuZz6/rFEqx
x31Mz2QYj9Vn1GviaULz1P0gB9p3man/C+eXnPzEhNKMbWvP2uGal6QtodrG
dZ0JgDP3rv1akbLhaxwAVaIp58KXW1Hqm2chllbQGdLDqWROcLVTZYPQws00
NLuxpdOB0AzcUcs6AZvktsOMFSaFQV9WmrjYUYNbDWZR83NjZli4m7/rgEIU
9l9GoKD719+ZinFoqjl+4UTm22vm4Q5SY05uzZh4YAFhrph6H4JfFTuGJ0aR
cXIgNt41pqH6ExMaEDd1hXfHv0e2TRzqtOPPHLP0NSAprAtlMayh64FVTrTo
l9IYfViNmtA1P2ufG2UaIUs6uonBv41rhwGUcL2yhrm5p2SFs2QPIaKHcUS6
HentMXGVqNoz0F5xeMC1Cmy6EzU7OS8+Fw+uvlw/tcctvI8DEjwVrfPktCqI
LiLbstLaSz11UtXn3nhu17M3N20uNzhyEvzH/SIcZIDIYPoDFCGuZeC9HuR0
GusUQLGikq+4lAgtR5GBEKScRjipukGQA1hwQUJqJHO7POyVWasytVlbnrpf
3/FXWXRqmU9uV/gmvmyNRY9mAZrdgqSZUNCogqsS0gMvU6DyaLwhGI3WC+jT
W4wsl1pMb5EIHRz8CcJJW5sQjKhkM+4axNOWCcKtQRdevwLYtRc0G4VUz2aB
gL8SGgpZmpXANmXUTaMi9aePdRyc9hMoxjaSX9yFvZeW7DgnaEu8SlYlYjCX
ytDDtdyH4sMlhrRUUG71RTS8cmMaXHyxAMRCbbj1DkQllFdifTubuCzH8o0K
tTKX+ViYS09E0V9SwqW5I+rPwhV3lbuwpWHb2GTNbn7OIzV5G6+MUK58O4GE
kXY0syOq0MOEM58G7WrQdRLzKZs6O4jefHQFOhFz6VabBC2tdJV/cDoCAlvz
iSYYcLsNxAzWQvO11a35LeVnJjNB2L8/Erv3lqWEa2btwc5Z13h7BBo0KDkE
yDkqDaZRW1OAJ05JyeKTTYk8x9/5HpESJRusSZzCYO/0rdtaKyXm+ztqI421
l6aUvTzdz3liSIW+Goy7sVuCNFuV6yX2fwYvEyaRfO1vkAsyd/d2AwNW76zt
/OMluU/u3eg6G17DmGn319DhzRxuI/oWS/DApGFdO5pBoQvGLgZxhZ6MNg5m
nzBbomHd5fOHabbFrgGpK7Q2+eLtyn4nPGLG3ULsLJ+/mBES+jsQ3K/ZLlHz
0qDQTb6cyKz2iAGUe+gB0TTYbSls+90GzHQzVNVf4T0wTeF6W2KXFSJmuCRD
xkhvTQkH7lQPBHQrEcWliZIaIZ9gcwJoaugfu2SOZH1e+/T2wL6BOrdzgPzm
Msw/wPTxnzKfW/QVKGRZLbjrET7R7CjbvwVDMwW/603iO5Az6uqXtt3uBnKf
PwYsjVQb4ErjxHWlL28gml2HqCbnjLb3geBFh7n76bWKhgCFxrBFFzbSgufO
n2EPekYVKgKJ+Xb3JmmWEScwzPz9sldwYOXtkW2/lmfRk6rONitiNgii/U4T
Zp0QpS4gorJbU3X3BAbfxxbblF41vNEY03/xBILlUyfg+SFNT/E4c6oLxqw0
ek6edzmiyaaTkZr6tvD02xbVKWIm4TgzKUfnBdfva9EFS8DE5OQUwnAzULpG
PFBXhiUxBjW0pc+H/GdjOqLqcmtgO+OFVhrQI6tiW637yZUUdcASYz55PxcC
R/TBibEC8gjj0q1h5WD3CDTKPDB6zV2VwkGhWW+y0cRlfOAYhnmci6TsAehO
1uZ8vCi9gvCY3/+ioZ7FKuw9o81B1MeYhJXSPkdwsg4M1E2Jg9UUWdFe7Z4T
c7rK04PQczoqyYviavpHIMwPuliI5O9zmIflIMxGjPlv7hkUq7xi21UADrMw
+1Vfdn2xZHPEXT07OA50mzpNMzwJ3wQB+Wedu5fkdv9d6oTJbeR5yYqe5qve
lmrxcPd7xbdfVGdbWL6nGc+CJJC8xS43rED7khNC4+cwaJStDStnLvBOvmYd
xWP3l8okkKZI8CsO3CDJDc1V11xACKy5INURU2RwbgWn4tlYsG11rhC8Faha
PzeloItqDg1MWRBNvCMQOlTIKdrzUsHaU7O3yjeFpAnVMbDoH5rNSPkgxCGV
hhmBI7ec1knoFIt9FAsHKIgCrqFpArAwoqqtrGcdw7tDUt0MUCi73j0/eEqE
/J5ZcALfcbRUtqlGDpN2X8PiMeUfE9H3iHPujqtES6oNwu/xhWygDU3gnSB2
ReHrM4VBn430iYf3TPsX3ZvJrMnEHvw/LTuDsTXnc5tmwImEysUk83g1RrvI
4B4mEq1Q83acwBw71sj3fUYrA+txpai2T24JnBi1qTuhMm7x2huBqedZ/H1i
e6E+M+sZmV+M5hpPtAXZXYw+3rGC9FC+2GSIm+StQGk60/YGrCqcqlbJkIUq
3wuLaF93aYoZuQGW0kAtX/wBgRxsaTYAeGEdR06T9yc+jl6k94S8WSSN0SdJ
hYWBdTgXA3+HkhjZr1D5q4GOXS+SWF2UHZOeUQ7kG1RGNexpfVANRXYS7VPD
qBYOV4c9FsT5ycMjPS/1ukAEx9UkNoJ6Nm+NEpFlyz0StfbaAE2yIl5jMD0O
EEajB4X+WuNMVk4X6WMbggfQxXzKBYtpgTYfGsiHmiQ8oxkup8l2dyRVI9Hb
HBf6UbkL9y6sjb1q+TJ8ZX5uqP3mT6ZL5PF3nnLzgTBOWKasSWu33hoiBQ66
zp5t7IciXsY7lt+CR55GjX1gRZFBqxf4ed3vc3w9/Kg0ES0Q/nY8LLdF7fF3
XgGyofenLzQ7Vt5JFTUSTMzzkJlRKPp7WNw4XWwwzEp3I1b2aSQdoTdKP3FF
nPYWAEYQCdRwpfHS8gfInM8RuZWOzIize5o12kuK9t0Who+squcD3jm5QVde
7IPVt8sI5bD3LrQOb3CI6FPm1r+RvwLGuCRChmLvoZEpAAiwKQSbCZEqyesA
iWQb+uq9kYAg7CCveuk9L1WcBX8KRLubm+atREI2DkT3Xrh7zErhHqoBLwQb
91ZsiowYFIsrY/4PJEBlq1odWlEnWr4m1B+L/eUNDppMdwfskvVMOVew106a
etHl1IiAQkxqzXL93B5+O161n4eLTbMicOS9wMSScMdQxoctS81jjfiBk+47
kJpvkylFuPDlsNdcD/s5I/v4BFqKAWBa3i4s7F7pCXvtUj716bs1HmXZuXzL
g2HQPTFMdX3nIGmnnE+N0brTrvwXBnfLDoeP4REcV8V/cB/WbKeNoaHnm4QJ
iVVkS7WAzUDId7SMM8QeoA2PvqjjjPtU05YoX52yKF2aC1W3QIns4AGp8lgo
iE9OedfdRu6LDegX+rcJaT4SFTkwxXnpyiUexH8Lp5sGfcxEbZsYJEm79WdE
r+GAkA/8P4ay8fNMf+ohNrTY5okAexG1vh4d0tI+uCBi3OHoB4ssOBwAcDGu
hiDPD8wtN1JviAdHCnE/1EoTJiajYvKZEfcHYJsT8sUBDsTCOS8fkwWcNQwh
RdQeoHOmvvcOi0iE+FBnQwpgNXzDWbympG72St+sb+RWE/UnKIqaWEGUbjRY
DafSYLHWftKhCmd1hLN2jSG+nRkSqXkkmurfU+3L7b0OlQofHDOHh6Gmxuaa
12MZUpd3q2Gik2TBixxPdqcjcuKlqlh4OPHJPs90y60/52zMzKjeF3zPl/FY
D0LR6MNBjQVOp0RrURMjLaJUuuIyRjGer6UeyicxQzCH1qInhuIqU7Cgz9Hj
u0cP3MW6tnHVeSEQC//6/KLjssZl4PyGvdzRfHjc7xbG4wQEl1yicKR7P5dx
YJieWXPL93GmpOmx0qWHuQ27lHOwFf1ze1bWyLahmELyJEGbu6bgEE4+I2g9
MrIpfA8lH8BjbOAdI+NnLgGNlACx+iOTaOvetPJeDyobLH6WHoSBBycTziDG
T9Z8QaCDG7Qw0hGL9uH2o17r4FX3TECajBGs/SfVYlCwelZrxp8jVfMsbJwu
4JLSnz1YW0EZq2iW/KDZGBG4uglOEJ4zHS1xckU1iXC0sMq/LX+jIo1pumIo
HOY+Nopf0cA1lYKSkpTo3vm9ZxPEiryYXn6Txk+nOhY+3Y8M6ButmsVooQR6
10hCyW4sLjasfl7julmg3Xg80abmZvE76hfWSZDmbDvNY5mYoruzQnaDmyya
uF8UK1eYURKNx0ZIcKwzCnqLuV7kiPuZcwzXtv4Cj7dYFLzWA/eof0SZfry5
WYy6Fr8Gv/510+abGaVmuRbyxsAqf2rYT4BpmJJ3AGWeG16W6QvcfEWw3/3e
9iWHA6XVnj3y5bLs0CGf2TMXZ48X5MadYt1cctHVYKYibCMU7kM5K60qSixv
LIHAe/8vTxiBk0JZvL5PohF9Nk50OiABa1TqWQjQvuGBGzAvZyiHr/w9+/9S
anp3FOKYErOypUXnnEAc0ru6zFpJ/mn9a2brr1wX7XpLGBibBwj/30f+BuLz
ZFAykcBY7fCWCRlP0XcKp1vy44Y65Na7Z/ce13Rc3AXZFE4NcbBzbs5Ir7Q3
EyldtugSJJHcvviLe5CJBYT5OIFhHsnoflY2DW+/UpoVXwG7Vn9muRVia8RQ
TBtUY63q1LzK1JSPlL8KT/uzQ4Deq7Tq4CxbaktpyCcaKvV1tBdTN32BIsej
ZpaXnxAXlDciBHIyWsGqbGq5YaqfMeJWTi/5GguiUSKEml6DTCRPK7I/R/fd
nku3dmMx3eZIK5l6kEopxEYjxL8Dn/tBggqpgz1pZ02GjLTsx0DGA3QyRmnT
4Kmmzc6jFXIBA3oLndFF/nzbdX5fVm0hP386U/S2epPl280P/N5REuMOvdvj
FeXiiecAExmyLCo6R4kufNFEhGAiTMc5T4OkcjZA+XseQqGhcawnYE8D0/YJ
Z0uPo403sLcKzSLZxnERUfDlS6b3ECtnSOm2RMNRKFuDTwUY1vdqVr4r6Zwl
AKKQgzqiUMN8Yd9d7KUtn61pOAAYHICF1PyFMGjMRg0GkmqoAbS6BKfBR9o5
4W1iPOKi3QjeqJVuD5iyWSjUwNu+kOyZnFbxnNsFTk2sEQ7UyXK/4A0RpbO6
9vCs+0BGyaZZVVpVW/gKMn5nzVK8eX4GSjwSiqR6O5jQz6y5DB6QxbKJ9cVg
mXEZpNszpuG4qYJi/GCzFYnax2fMYLl+Fk9r8SStHgP3xEGKOBVRx7KU0u3N
J6Z3fMISEvUPM9UV5MgnGUSWhnZ/g+cVzGMn9rEabbE9B95dcDUx44BYjI7z
5dF86lxGiazSncZYNsVgOcY4KnHpC/kD5DxpR26GLzXDAM1+5mgrYpOwsNNc
j26OFef8EkoodhYOVbVrocYwFv43ho7LsV0tGt+28HWbxfkjp5cFngOrVWn0
C6Y3jhmsqwUr3kA+mQGqW3v0lwLJbQ4/v5ShNqDl2fJl0x0tNVbH76OfpEhf
nyapZ0HsyCGjWKN/hGOtS6LxR6XrE9IZzGHwa+LwvyPewN1cDf4gu/FO9QMH
f/9ZVJhFkAaGAqZzlQGC1wPap9/dNJB6jU56gY5/0Dq527qKs4J5oqXWHFOT
jzX4tpXgyyxpMIlLsliocRHzpc7LqIVojzvGnNR1cwhoBHTMX6E1mHis0iSq
KtevqrvQMoQFCLZMdeO4Se5nPeeR6rlFHVqmXdGPYMNpc51YKRPZtWN5fByV
JzRztrp0muIv4HpI/AiqlBGkEhnIP/gD+DFvCY3PlW2Tl7dscU4GhlJ7gX1d
OUClDdAgourGlEbkVjflfZ7jtDfII5Pz6zFUe/PG40ehvGMauCkwPET346kx
UT0R/cmHhk1AcnMVcnPXdbtKoLM+vGOhQRif++4gG571EOI3Hya0uTsDqKvG
BV3tYT/UBhnIlmHMczIlFRrgFChB7ldtfOzMgLsWaFSxds4JCuUEYZbXSCbT
BFSGhyRj1SegDoY2dFYvMJH4o6gXyVLZNLVWgAC49hkQOH3Ngye3fuxEqfqF
iUWDlEvGtZ+iFVI1A5z9SEVdK+/LA0bOxNHQO4Yvq4mV4uFM6zVYB2H6Bmbk
3hWXmtzqUtslpud6E5pE4VnAG0gz3Nl4jLBbywIuuxI6Z0HU9CxatzXvTotS
HvQ554C2Cc/MkcdX7lVr/3p6TftapDL0RGd/RIgO4/ng8hnsVhAFgKKDwUys
f8qvO6fE5hoUVppW4gNjpVIx5wqktYIavpR5vVJ1b5WT4uzOMVMJzbdMVM5T
03b4W6Wfw/WsbyUBDO5ZVMJAAB313AM9saEwrE4/3S9hREuuUYJCPvfFoxJG
z2Dr0y1azK6DQZWI0L8O9sfxiITLRGit2bZIJnef4V5Ol501xWYOtBDXjSUC
YM99tb+ydezpOgC2r4wrh8BXRG32+ROzp69M9Q439vhYoMQueMqXeCM6zi6z
PS4bkPfWdS5XYwkghj1h5jkxIQPjHuaUeXxwRb4xW0au4AP98uUeYq3Uf/Py
+eWB98QlT7khZXT2N8Lq9WyFQWcGioIyNO6GLth2bxR5M81pK629Bd9zDI5E
UsKXyAMvNygdpjJAfxaSNEdkc9ZpywSTs7Dw/ZiiBs8VWxglthjh2LJ/owWe
c38XRqa8Oq2sZB9cbidCrlN1C9VNF+3qa9x27mpnmL51uZsNwtLX7yaJTCCI
1HJsXLd16VcFl7cuF1Z9jLJaoY3bMZ4rOeqSNRJ9dtX1U0wxvw7BnrZCsGYn
Xrkr6VPM2HqoCM4raEQikwe76zBMRVBvrDwbT2AJEqyEYbH3aD3Kwpl6iUh5
xBQ3L4lgazvtvLfmEhI+CqnJilkYy8eqYlIQ9uHOD/Xz/AfAHo47Fih0iJ2v
jZrzkX7dNQUnfhahYi29ENrxCcVD04UA9ut3wxas5XXyXKULUZQlH6x9YRtT
eV5FSr57/vT5H87M+DD+amLnAp1firfy0WbhIh7dFHFzT4Ew1esgWaHptgoi
T7SiisYx4vpTJnVZhYmlOsAwmKUTblVkWXOWgSTnK9h9zeh4jYxVjK4r9q2c
U8emBTmzu/KoR0pbUnu2bTNheN+N2cRTSfNagaWYtYPR1sN0G2eHz2cHoC3n
WwHJyLjXLGMFuI5sHxW7UOy15cps9VTPJ6SQVJj+JEcAg+fkccwiLgXc4M5p
COYRBXSFt13mU/UMRXQu5XQrxV8D9g/HuTQ9ntIWbS551Hn9Uk7TG5aX1wcD
5YNOGtb3ot3bPe3fTBwcGgdQaBNiSxSDhY/Fc/cDJeyLanEcVbshhWqovTuM
7fLoAat+eZg/3jK1l8YbKQSZlkdPDSuvaIIwtmbEHA+PlVpzE83D5LuVAt2Z
8v4VLiONh6urcDTt/34x4FRIVeToE5gnpP4JdBi4qCYbORPybIZfK3n5LSPg
/k/NAXxy+hU152oM4LxyvGv6/O7WxQHQ7MgUiT3yVuAThHCLXGsb76cQ2uys
0M7B76r1bjNmzyiZs83U/A/a+iJ4wRdr0zAdcZhh5Sf0dKpAanSWcaUmO611
8xO63knyRPrYGwVAV1e+KWHJDqMsNDu87aTBmzUzrGSx/5NUzLnJKPWvNtfc
Yx0/MIrRyMLGwmIPqG0E67153391LD2/ZtCaLnPTvlG5xhrXAo4LE/tt34CY
Zxup4nHwFJSM4jo5Cpgif2MNtYmGeXMrIXF3hJtnIq83ilcsW6qYih411CtM
M4XRstFSvKVzXPbyIT4T7XybZRxreo3pPYFY0nww/clAlJLUQ5Dq8+RO+XVb
eVu+CkfqQhzkofhaECpSLOKg+QrkJfxnrKeOlFnnrU/xlsuRcXeTCYB0711n
dU6FtFWJsPh745a5LSSgWQvUOzzNrM225ANhU6EGIb8dZOwv6DHyuYFGlIf+
RWB6jK5k7ncu4jcqjWp9tbxLfDtlTE2Xj2Nw0HKhesHZDWA34NUe0aEIQTCg
6AT8zBsFQXlbz+LBUfbf430fXApsEpiaXXqPDJ53j0fQI+Obr0ZIELtdT87a
YPg5kEsg10icXJ/LmkiphTzcjYmzfP87QXT8LO93+ko21HzQ6WjJF6tUzhgQ
fNX4NnSPTPEDp6a+OdtGUpccE/bRgknViVc2QUmftcsXVwODRIZU5/qgfjcM
hf5ehzH3hfpNu7c4IjBDQTXYglqwTjRyVa2xD1OoJwajqs2+7H9ayW14jHRQ
hJ9jeLziOFW7cKvkw8Gi3ABDQGhCRuO3qFO//fi6JYboUE0bPvl/rkP0MRWx
ovi56JzKyCfxFRSDSEyJQujXqc0zGWggl2r1CfT4bQzf4qUOKmMd0R8MbQo/
6FGt2LGvzJ27oxaLOQ7lIFVyhIVAj4dYIN4nVy6lN+nPLkdakJu6GUtWh++4
sQUpYN11307JsMrgsiD4IEjJP7Mt37VyDIIHpvjSGdTZMe6DULcz4d0nU/o0
Q/ZOzWxB0oGL/JrDV2y6neF/ADp+hDJFIyoCdXxIS0GnXt+9cA/Tu1cmQcYM
2gvdOQ3mO1fOCX+b/nvcVBVsoO42VQZZfkMrMMa1l5jRoNDiqrUK1zz4eHC6
D7Rll+mbhQokVjeVcwUHiBiIx9XM7a6qSfGpFdAwV6JeESm2aKHP4NwAOaTx
073CZKHiJvz+d5FOL9ooisWSUxQBVn6Z5mEJnJxko8xpMTUp5ZDt95Ni7JFu
yQXs8cCxdbtjWtTHgoOWEsjXZhlp6wD/Mhce+xmT/EfogFA4GGzky4JR9aD7
34KT8mq5/4MHWYdn5C4wS9XQLbihcKXc/i8W3w0dNXJKMFSI+C/V65lE8bZH
u//WGMBX3iojgkjBsA8PfhYGvRPLC3cJVraqynUrD5SXMZx6EyJ9Z8Dp+2vX
IREBr4QndhzRSj284ILx2C33gNXbOQcZYuE9XwdNTRU1XRHWNOUiGSL970xB
dv4J9F9Uj14L2/yisBtuyS0ZKx8kU4PYciAoYUYCGo3if0NvLqqLTIAMNGvC
0Ay8rdODWnUMVk6YUXDuvqhg8edWb0yygGpFXSMJHn9sOL4IEQ4KvGg6HvV0
dR6T4dsKVAjBDxrhGJm8eqeZsDTninP2XHK2/ZnYlE20WRObP4nppLM7/gPr
eLR9t5g0ivC0Rq/LRyu212BSUq/GI4CycR14fH0QQJplN3gMRQ3g2BKGUUbX
9o+4fxbObE6hlzJVRBwF6m+HCFzUXXjQljoyHSCVc7TaCEgHB0AZXFv5/n4b
E0MHFjt3/Zj4jT2Jdvsnz413Kv/N/1MAaREU4hUaU815JEn2ABd4g18Z4ixV
MEtwBa2Nbch+hviziclIq8uM8Fcehy2SElcaWt7hGvxFuWfMjbBpGEd9Fj46
8qOLmjEC+JL3EUNN/MNaIe5nzjxFOKRCtrnYLxXXnDE83QM8Wu6yoJx2ZwDx
NTrbB/Qjl0Jv36pUMLsm6JhB2pPlt2e/lIaDcTlKw856L5OCQRA7js58zXy8
Ivf8XoTFg9x1i0M/DnfZVZk4TJuM+5EWaixW1WurQWrA9zg5xmFY28Tpxlk6
lZzr6mb/8bAMgtvXgim1Uu2oncLStdkPp5VZmAiquWD+PVYV8KtlxjGfxTMQ
P7txygbenatxi/YoaDTlHpL+VbEX1+QxOUjBKzY5VwY0Hu5x/g3ppaZqJzXs
PUP11A4PgY0n/dD2TW4UGSalmX19MfNTtNIcvpF3dv+0nVKP0QmY5bJ2z3tV
1Y8JT8DQ3JB+ZOK8mZ3JYuY2fvvTat04ihD2EUi6umy+DWYQ3I41eSSsAVxx
dkj3un66z4ZR2SWNovn815fMsd9DCEcrIknAyvZg1p5AQsw7bXmcNpTGHsqv
Qdr3Dc26MHP7uw21FDPjpMZEHsLTpSTiSc2kSMLq0Vta3nesQLR+5Vh+npXy
JMQudp9dMZmeSuphMAe4uPoXqF5sXHU8P4w86wiGBRUEBVA6f+C2B4AcxBwi
OI9Yled+nIol9ffymsIDiPxxlsamwPrzanWdN+ORPWzyIe/Zq0UVFtMhSpT2
pI+t3n9k4+AIEgthd6PXqlOV1kU6FYjOtsxNl8vn5vy4goxafIOqWUBZ1gMd
IF5y094/Xw6oCzMQV+Z6j46jcbjezlHPzk1zts9mbXfREsakHKSImeykZXba
Kk1Ppl99yZGCFdHBGYNJtkNFg8dqztX939hUfn/PTAjX+vsuKRu0NI4zXJ2w
IBCFDSVKh3ebE71VG/N7uzNwT9gUSELvh13tKYZSz8vWOMN6MEX5APO0+hT+
u9OIbae00FBZnmDpOXeUnVq19Ytfm5J7QuPyCTvie5lVHF64jNetFQw3FI/N
JN1wmyWxyGBoiw823USc1WrYEu3XPJtSAZccVEogHPMaiUF2jHN9OMp131Lu
XUHKMks+glhdbVSsaKl+mGjuMFmJq64QEDhzSbYNVbSssTNBJT37t1jgCjhp
YGKszWZWGjnPNZk6xtN+rOcMjXfu/i/dL28HIxtcycxX3T5eAxR+IRac5+NZ
dcKhNgzkYKSq9ceFMICnz2rsN52GntKvoUwh/ubTi1Hq3ycjD4GTw677Ml9R
16XgMJ6nnEIbnCfY+rPf78loHrZ4s+Pu5Y0MgICrWbbnodw6WQrwVcBGRUAs
eCtUDrQlgT9OPlYxykr0BKT7O8TERXia+ABb6syALpy5+9GT3J7m8ubO7BX/
AkxHDhCgvManLvJLifaaxNyyO30OVn4FxUSbr24zc67sBNU9NvgiP87DCm+L
5RR7Ggo4c5a5Ivqx2ALPh7MjAdv+r4udufNR60OvZRnUsgzQsJYyicDyS0nT
4YMhBI7DcAUtwqHNQECZrZEzyDDXqasc61uLagSoTLw2sRnlbKkI30z/AxdR
ZolPwdFdeCad8t0jwe97TZDTN7JTtBA1whXGummfhoK27i04syXsiG6nvrP1
gdWJo4F873p5PLG6Z1X8C4jXEMYMYSlovAXXdbQwJuZtONVx0VSlLrQ8Ld5x
sNR8+SQ8JgQxyck+WCt9LradWYZasVqxN7Ku4dN6+BucQGMZC4x6/H/ybZ2t
R7SJM2wkSfW9o37f5/CSvDMR8NaqehsFxsW+PpnwPY56kf+jA9Zpd3MwKq8F
wxu1JqeTzX1iDucntIZiWbz8hp9nqyIb5l1tWv9QvAto6L4ES1jDFVzJh+SC
rGkYmGa/iic2sTTHYWjg1bcQWtr2w5CnINa+BPhtIvWb+dfcRnKOT1croJxD
2do93MXjQgPe4aFJc8l50brx+HuMGwwRbyEGpMUfcCG9mUvS2mFX2DFXtRtX
C2gcW69EnrwvA67YBi3WiVInrrkTrB3d1+tNPnuthNxI30ozuqZktCrRDCGG
Nm17vV6OMRBG8JDbPWGLk0zI+FLj32WaZJKCeitTTkPqvfyGzf1u8ROK7m37
j3C//FR5gESskfnZAEg0+Rwr5389+EJ5Z7zaEU88tr3L4uDrU32ooRwNrS9Z
PgLnxM2KDUflB4msvPx+o5J8B6XVFQF6QHbC8M6A/S88+3mfMLzjOpKO5Mcn
foV8bbS0G+xpBPURCQF2JsDYwkYebssaMqwuX4FXjSbswl5/Y6KoHV7pXWeN
zhtRg2qWwbNR1+CLKBH7zQsq6pC2w/0Cnno05ZcJ0wpfAG2d5pQ+V08XeQ3m
fSw2f0P99Nlij4CDajaUqYf/9nPPAVWaJh/+hbDgD9YQ+RcCxwtVJ3DnYDjp
wXBOeCWcFL3/7Z3oc7oj+p9RC2dgOKB7gy9jz/ppKQmdB9NEdvBWHHBLamsh
vIFx0pKjHDbDgbwuih2OxbiD8/jBkKzuoawsgOlB2iNuucRzhGS6A2v24Dkg
WaLy66O+a6Uxg1KNimtz11yFRb7qgdJIcz2atzhzljWukhhb5a90W4VTUY0R
1EbhE+/boER0CN4H2c85Ssoto3N9sy2s3M+rD4bhoV6pXywPtlHtARNXJeT8
4O35sbQUd/OGLvMmJ4Aey2K5Zq5kdcjk1S55dhKLTMQZKl533+BbEp93WplM
kbv16gejKRaK/NJv237oVNorUa5NRdAcDR39QtzeruesA871CNfGSfjx5p8L
W8OexkkmCoyJPVneS1o6s/cKxWNObhlQvHpFwRWCGsm72ovQ2Oc/flcJvElw
stw4LTM85wtr+F1KxiY5rDDDR4+rD9TgU6VKYcAXcUKdxWXNzSSocj+DCN1x
+H+iFhINvPxZ/5y/59wtvUAFE7o2q+HBpipPFRZn72NxT05eGrJeCCjk6QrJ
LRbv5sQ0TRSmxKE9yYNEdiqZcTjK29RsJQX9oN5h62FY5DLz/2AOm8lWmIxR
iXXdBDxNXfGK6bYwaTFq7nHSxmOVP+IFQ8FV6nMN6MqSJGv/H6p61Z/7HVls
zRyxo/es0ir1qDeEOwZSMG58fbIZ48p9eWe2YEH0VdqqxwiPC4vXmSos6b57
CtCl6X1NVodUmIqAY6TPLKoAbnO2TVrV7VD6ZDSnHSmBQF4aQm+L9Eyw7dwF
AkoFOn2MaI+6AEuSeDdJfsEApNWvAfbIYWokHk6AxUs4WeJ8BT6J89pxXyuH
xSmwK9ux5nUrvIXuZtAGQ5QXbnd8DxdkuGkizTsTuC2Q3R8aLpEBT06un4Kl
l+TIbJWtOoyOqQF/Ht9FyjTSucRShwmvUSdRhpgb5vSXn8QjfRmnJcnwsNyB
xPkTVNP7xwdnLEkw/v56bPIHCk1LVhcS/hsrB6xqkgbhib5ftqQZRmyk/zTp
C+3q0xKehRyu4ehzMYV9Q1MXtPHp4WKDh8ulKDtuegxUUADkv+5eB/8sfPVW
lxVEDIssQ5U9poKyngxh+uBtCbIqTdZPKITXZu/cI+cuzIwtCw9FBiyzIP6q
0setakseqnPVhR8+Oa2OydGOITNW4/kYXtrRkasj+iO+mEbtK48mRbxr5vSb
Uqp6fRRHEXaqBTK6PINaX5wTJiIudZHsfQO8J2iD09CDkj8h4BqbFIlpW2cY
jiRvpB4xABCJ1cDl74SEGJXWP30hRB0q3W1vnUM4neOwS3MVq2YNEmFwA560
SzdY0IAGaBK5HTA12SQ1m4gSal/MRbHCIIvhf7TmCxrsl51tr1LJ+fxq2aUp
+vGVvpQMJPAVC7MnA8RDM/ZzZDTHwyXndAX92N+y/i22H1wWGDbrDuy5rOgL
LAjiF0EXFIZZVwEb+vRFD67FMZiBkxPfY7UEuFwMHjyEceEaUlG/zdbjyJbG
0otmYQC/VM6gSNkeJ8kZM5DqRBncOFsDKisvsepMPjGUdpyCXu0OWZVAd6dS
FjNHuALiqM51DI105991NhSuJZij5mdKIdvDUUT9fGkHk8sCgQmV/WGNwOsy
oa9acQiNB2VNwyZRzS6nlFcxaoQmK81BGOhVTAHN4Ov5eEKuPANuK4Zhywix
Ji4Gqlewwsaz9OmfbII04/BnQB4fXNix6gs2soynFqEMP0jnm1VsgCnrpaKZ
LAySsYkraRVN66AfZOC9yY3Uftr6ALfANFGTveVs/f8b6yKeNm3EwMp7CD/0
JOiF/4vbx3FuD3u8DDK1jzvPdzpk2D8EPVXZ/WCatRhvxi1/lUI6yRgJQzo4
23b/AyZYOf765eLIE7dtoAmj+g1tqLShfMNoJxReeJlRlxSR60kUO8ZyxO3Y
4GA7lAUQu1tFy2pQ1KUQsDdkp9/G2sJgcmGwBG/HU1mlWHSsvO8+vVDZix5b
4k6GW37Y/hQhEbOlIRTq7o2EsjwtplRES97xJjky8VRWgDKBLKQYqBx/EQAA
1Gh5JZ4I4Gqm5zZFhPVV8Zvq85NIS5XExZ2dLO0ewHWGO2p24vFoI/3FlAlR
DU+N3sC9hEa57rQ/beMv3FW2TqJ1C6/UM/c4vdYFDlCPH9ZSfuSwi7x7NJ3P
E7CxKvPIIstH8TB/316Jbp4ChzCt6Wvla0tRkv9tHZcyaHRf1X1+CH2hl0OX
DQ2Wuu722Qt5gpOJL2NYI7G1OaFvgLR1Dy831uCo8rzJbKdfXqTcWUgjV1gR
H45WoRkL/mlb+49N3Ej3PBiPjqDEE5wnWo8YAsrL0B4bRmCsdojg2xKsNv36
1wPj+JvxOIA6x0vfuQW9saFRWgeznA6mi6YXR0jxgvVehQ0GPWiVQotioq1B
EnuNxZkOC2E1vwAJSYm23WzW8E/iwDwR4VqNYhN05+yx8NMs3IoG21uRgd79
UEPXSabfbYXMh5ttyIQG2MnLsBrr2yyshO9yjoaYJhMw7AxEelMk0rl1bjNZ
bDjnYfLHke8fCPmcpApiESFIt225Kw4xiDn6WeKtalTBrsaq9v246Ps3zVss
Cc6Tvgy4S+BzKfXNLLCqy08OVpmn2eEvdjwwDlymvYyVDH976TDj3Rmu4wpJ
d0LzoNi05CtFnbtANZZwu+DfTvgm7vlYu6YimLkZ1ZcWhcRx6qRT34Pd3s5U
cNe2xKPo6i2W0/BkregSsfgL2dxdsN2dEhiRY5TTvqoO+nw7SCP2rhQcE5dH
wnR/T3g87QF27qeoS+icM4Ild8gR8HP8yLw+F/CinnsDJxdOYFFCEFLk7IVG
3sOa1/TQSpdwlZGkZRhGfNZdUO4LDkgBUlWmeZ3am9RCoofYx9d2fsMoWQse
sb1UHp1Ez8UGhkqRU3gEQRH710m7AUtZKj1nokJ9BUcuHS5f0usC+hVdJiqm
HU0EOCsr2TSZquJzw2IH6ra1HDRWSlfJom58nkfrrbqwRMNTz+4DxGzB089b
Qy2l5IO1oEEUpEK5FRDXWCbwJyI9gMvbwfTPMgiNm2GWkg8QtA+AOFZ6c4PF
yCW8VMBCOwvAS/4NxrHhygFxqPT0GUtjguoAgKsoanxCY5Ltqj1FP39SvFgq
tOcUUDUU8t2of2IAdV/K+znQ91vPJf6SCicwPjCc9vAySNa0k0AXNu3/HCRw
uMVf+pgTUx1Jtykkgx/LcBp6ssx1eEqsp7xaWuIPCSDoeNKT3FSUPi8faV2A
E1t8XHzRHYZwkxj7X3ahrMqrYEO3NjspkfD/6PPekXvGpu4LM5VD3NO5qgqd
Dezf6r4UtNszcK2Ffx7P+ubkQDyNbNheAoEzPHQ7DGrJIYdqBjwGTVVH6Bzp
C/2HtfeyvsPDkvNGKsxayZY4QteZcMSl/11f3CroRk2jjUGOOVLpbRKGctqf
gvmNguvFLERpO691JkTdbbvYrNZig9laFX3r9TZbzR6buJQYlXGrkN+EZcYr
XlytQsu5S3NmGucmTlyMB0PJYrLupuypbIC6O5lFHEz+1Iy/Tcb60J/ARteA
WssjpLOPFqXRzhcRGe4aJw/HLBs1Vu7/FbuHrqTdBHDeUquVPDTfRVvdm08n
UQLyqxPyMIq+O5eYYtC+Gr3angXQRbSWXmA2gzcxVl0XyqZwDya34+kg5fWw
+TdEH2LPInyrNEaKXrKB9bVdjNw8l7gED4d/Wc8f9he84F6nMSgY1jsCt34n
q4g36EtoAqhIASz+uN5DCs0Cp1igtLjDrrHTuExE3lkKwJlPRXrG14dXlADF
gy8Dfm0Na5z32dyErRNMm6++poHuZ6j4QhX5TOQFO6T/eYilUeM2eulTRw0n
QtxadwPqmyHQ+mtuww1q33gIWEKgOQ/AgOAzGvWo43TxbwWzrXXl9rz2kn04
hOf1efV8dGi199N0YHGyt0FdoTLo4cAmkOMsYgK9DAbhybK24SSPi7CF5ZqH
zuzt/ylcOA+q+4yGxgOacjhH2/JtuFpupeHv8LQruuifbJAjjwECOB/VRfIf
v0V1lRpb0nWH7YA2K9GF/aw4u8GQwqbnIlfa9bmJE0epNCJbMvmtjeVzMCHh
UcT/eNMC2NKhSEFIGtXAuPqZSjZ+5RZV0Jyj9mzKf/VW5ZhHUdtdNJJf1Tc1
x+xIWtqx9/lU4Wu9TxqD5bgHskXZxyNGKD6szqRmmcVGXKxKol9alAA1gpkK
URxnEK35cJ65nZfunMRlpId1HlY7iTamcY1lMahok4CYHwLIjGcEwOxkuulS
1gSyNgbU0NZs0LKKMFEFUJ0/oX+uTrm6PND1yF2MomKsfldA8dhWpAJlkDCZ
X04eYLtWQswHGdoTf2I7xe/4+48QTgFYwqjXOKeAhjZm3RHTGRe0NdgxwP6t
oMyYoXUBCF4+8b1IGNG8BY1p1kMJTcrvQxG9qZRoAp2AQOKvnPc3QUc15nqW
vKTRtbXQ6H5ITEnIx5/OZojmpFLCStEvdWxBCI5EEOCev1w68y9UW7TaLOmV
VLSigu0Jv10Sf7MvjtjxymRu1rdu46Nue/LTyN3ouRgjWbn011dVy/Hok/on
iFd/+w+0hbkHXhsHe8sJksr0V/E4bNpfpGezuKVT0f13Q6veCX9f953cHi47
uh1mUe1/15NJeJGz3WWHeu8de/y2wwCbjkZ2WPwABQ3Hqltldwrr4U0rh3S+
UJcPQxPGjTkEPXWwdNoaPwJNI0qgnOwP7h+8j/zdkR1GYS8w490LRTqp0A4f
5dY2MMJxne065uiaMHSF7fBnk11x7lDVhEID5e3JSneqWrCwdZtCLdh+vmw1
ebW6oGBgSjXd1hj0CQuNTsm4+tl0YdWByL0AxOLXJmaIf15biFYSHyW8qXQq
kIQjGetZHuVXvASqW+kYA5b32gr1zPSQZz782ov+FqXXY4W8xJ4U2ik7ueUZ
zj0FfCcj3rbrH/WIjwimm0LP9Wd48AKAdJeXbSbpGXIrsgBWFLGJ0Jy97nIk
HvKBV+Kj0kA3gpCJHLjCAE7ozMIhTqSEmK6KoSJx8101FFKADuuXr/gMR/73
7BLbqLGFGEhZrQxgGyNRy9Kav1583iqIVu/qDoHGS7Zj0uyFFdT+bcyu3ptl
shnHQdTuuTYNG8ekffs71e6TltufH+zxIqrIzZ77d4e29bABQZehIeFZ9b9n
7gYYOL9fi7BG1rQpLJIM2W+HbkfJq00qfiAHiNy2J28DtNM9X1i9KTi+ARsU
cES/5iwpsmsDEG/y9HEB0l4gVzE6cj3UlUfawpmiQCKUewDUKUDXWo6+i7cD
9IwXep1vW50ShrSO1DJXlVuiZfT9SF0OY4eLhM/o0EVQQ7YOGYtAp6VRcHOp
hA7A+Xlzc6/LTXNz7ql5Y7+7U1NMeozpLnzXpQeMIiuORJ8PK8DXvgwQnIOi
apYmyrXATrLh0CyZ7absMAIxLiwMvYFRDGOIAzK2V/n/4v72LY4xvvy5Khfl
VCjFjBhCtYMYYg8xxJd5QVGsNFpb4iHE27Wjd0PDLmWBBUukCx1IlMttubyT
+P8H7mkeuF4bC4slKtRxu60pZERV08GB+B0bhjUsSxJPxqX7W9f1rV3ejixN
az3ANr1h8eVPc6htaJW4tP4Tbc8eHb11atza+binrmWM5Kl5Y/weTL57nsCe
D2zlDGH8uhdTaR07T/ROzcrvjn7pACcF1OySObIAEhEWKQHgvU4rEvtzcpgZ
4S+ase9pAyb6zhZoXYqZd0H8HTwjl0/M4LGbuyP4UWDGxbSkpZd3hsdrehvQ
JKraTyB+TZBlTW2jffS8ia+g6dZ6RVbV2mfzuKa6MA6Iy2H3OvMjKxSFXrPJ
NF8LP2buMFIFM7lXo8+eu2kNT+f7MNIXsBlc77vGDZr3ROqU6JcTQvd5pTca
zIj8IdqyKxekIhqE5twndKZKmtC1MgW9V6s5yCfEAS/Anc6Cug+XBRWJHWgE
h0bNBtUENb8OCFRVtd+I6LSWGhoTYvpw3me0QQPbwgV6brpArUVjzxb/yXvn
8vUxV0dx2c+8YJx1VpztFIET1hwTAjgUh5WgwbPcdIowNaRxZoh1UxHXYIZ/
kjfq4duQblxMt9VF8A1/+XL25lFl9a63HxLxB/uS64QVqQsmYD7YaBzboMQx
NOi1B5EBasAvOhDG5945ruMJmd8mzDlmk0bwUu0MIaUEw4xX6VLzN3h7yJw8
vmbuJ9kWHKQPEEc/oTe2dBpNUWGas1wmGaoPC3405jl+K4RP27lYYFKjg0m2
cWgUFh/BWds7rgUNih+t7mfcVOKokadVnRUv5HyyAQBt2oO1h5ARTtS0sQmp
KFL0KuZ8rV0psjKKGdNIWSnJCIBrqZeqZJ01p0GQGgRtK52NpCA+mcdn/ZLa
RiMOZFSGi5bQ5K1mmC4bmG9g0uWnbhP30wx+cHBOnc6RI6R4wGSsUp8lyrF0
cBh7uHulvJL65mL5v35Ka6QNUqTwjrpuc0QPMZzzhwx6yQQSWkviZpQQL87a
INfdxQqUN2rapzYDaWe//9mZwBlnWsFLkRgz5GGtBmdopxDyKXhEDhRykgeq
fyMxVvzBehpiZ4udkbKB8pWV31rEZ0B8SdaG38tYlyIiXaWN6vhFBk5LTgEp
sG//3J+raYW+cA/L6MVLSQsuhY6VKhIzKDw6SfOaXv/vyIRMs6WN/yoOMr/F
AnHc8tkEcWX2kTwlfQkxb8tk1OPb6yOgtWrQjM1+gzC3OXOrWnPCfhTHL1QN
tCSvrRIqc8yZr1Wu4ersol/5FGayOQI/DHTNVRoeAiUE1DaWorbEkrnZbVju
qpwAtDRss092xbBhez5gQ1M4VW+4c8ktWHXjGf4hSF/7CxZLAM2mXWjEtZv6
4Z6PHJ+q5eWafFsDO6cToBhtidBHh46+bNfsOoYfgwjT3WWLxxVaW3epdt+i
9gyhgUjzGDsn2ZhBj6L34GmgOWmWdfdGOT6Q15N7fOHrX5VOlBJjF1oKskRa
FjupnFS/8BF8MsVX3PLUke27cZW1mbO5Aea1bbLaYVwB22jqC468jBS9njH6
cBwjOwY0OCcPrSdqbozO15l5auWmXR+1x45nucj23LpeOQ8PmSk+4v90N7v9
It8YgqoXYwZSYwt8HHxQyNQSG+CnMDd9cp3ZUKrTohCun9JF6Mg99+R1VnD+
twBqKrbTPspIIzVjgCGBZYOtyQrcseuhL2vvOEQ7qJo+52qXvrYJuwhpLMdo
/2Q6myFlzO7IjPq9QYsJuQFBuRSrYm9dZN5kdA8AlUePLOXZwNS6YTZcfp0W
5AuO84kQeGBOXxXE3R688O9dv4h+6fFmZP1bKmSJsE4lkHS+eWDmkCsG0nnA
Mv0uaRpjY44/Wk4HpfDnh8KBOkhEN1ZMwjdOnrRkvGVh60hGjYJ0Bj/jAKuD
lgKh/PqMjbVGPPzdB6cpxFiB15+zuRpd99VvRc7hwkO4PBER15BmiaDKcPWf
H0qu0tFMNQ+WsbEY71uq0nWUu5nT0x5p8mAcAm/FoblwOv0/ygWn/p2jnyBz
qN/8tvUuOpoBrdmBt25hc4at7BwQVWr5vYZff+XbSHig4mmLFqTUyPb20qmZ
pyLXwC8CshedY6+v5n5yzWedaRTghasyC58we4pRwE94aZ187eJ92Y865pyu
R4H6cyWVmKmKcxlV4OMxvpu3ZV9vo+5QCpt2cJY2eY8STQzbyGY4MBLtAQjm
dOeEaOLVAZDD2lYY+BT3HUx3sz9uIehtTIcn3ZePa9jQ/hNLgDxUrhewFb5c
f/pzYsbNthk3wSqZwhBf88KEfas3XMSeZ5epetx8DvHDnnEhdUQ1ulxNVZxv
cfMlgQaMLyURPJG3WtihrXQepVd4SoZY7WVdT7ICdjQdZHkja02JydXY5NFt
syHjp+0N7rSFuw8DE39NhsLb6XN8OmMCTLTO+3mbUUqfT4XsjkRv1/ggaZ0C
oAlOSFGqZAsVcbBEaTZ/AGoxP7nsXcesg7EJOB6TTt+WUPNlwuWKmftg6yVQ
R+B9kFA/FcgYehpjNdhya0T8C3Kwxip087TEqyncpWhz0HQPTEt21t10myRJ
C7Tv34YPPiGjyq2wDNRb41aFs82FPK7Sqic+n7vhR/XWvKXYxqChrAWxOO9D
ujVVb4NGfwFUlPvAz43CzYpcD9/QcUv21k+QpH/eqJ80NJY07dqxt8ggQKmw
pPe+LcTA/gE3H8xHa1BQz5DRXkm5lZd4JcN1xmzSW4vhsYdM4W1OJLgjCR5P
VKnC1PTwB69UsAVEEoIu/uZfp1FQWHRzpL1LNjo34CEYHuya/xyLb6cN9Dav
pPeQk94r7sdNWbL7T/EvwSzDgit8qmMxbPPXNPgVuvljZ4p+M0OlUb0JkSWj
IWMf3E6YWXSE4qT/7+tkPCJGkDevlOOqw3dXwJ8xLh6mAp5x7I1oMtxksxbh
JXij2wLfPnttI0e3IynBOGr6P11OUKBp8FqeTa8oJ0Tfw/jLHQwlaWjcngGn
GwoEhPTK/afdiYoWdqXaGmLkkpts3BFVN8bs+VdBZWzXFOP28zX8L5Qq6PzA
UF4Udemo3ZD8B368d/V7DBmU/dSjqYbGkaW+yAgaOY98oPN+IspR2At+++Bb
21hFO0Iuiv4L2uX3HQoSj7h3i49vBuyZE+qmLOuZfQ4gB3tqYXHH6dk8k0BQ
cnZ5+lDa4Wnz/sbCH/BbYJ0ONUDHjFeYaf69OtD/lnPEhUhNYoyeE0amJGvN
20ebD6xInm//E/oiWxrXHTfrErBCMwy1yrq2+sU9kkNjtk1IisKBLwnU5LMd
BFhXfn1TpinErStUPyding2f2XH11hCBewXFmrz5mUmYjYijT3ey5m3Qmbfu
axd3K84qBgPltUN8Q+2l1OzAYxUObfAHsSSetl+NgQSNjgzjGlIjy8cGqORJ
UcVcDcNEUGKJEMsIqxpIhJdfC5h03XJaSDOBN/lEm+xPVPbd4Bxrztn/JJlo
j7GyLhAFHtwm029FsaejWMvhwNT7EaH4jp3TkCWXra+0QU9KWEL07+iFrLHp
k4L1jG/F4HSzZ/ydln0qr0ESSkB65y8he6OXnEKT8ad/8WQTp3LZDPa1R/DM
v9xQ/ikVgzhXredT6+Iac+XfaU0/2LlCMDxLJqdwGrVI5L/4rKuG4v5d7YnY
4Et6+BuC9ms8QFpojP0aCq3BcGGNbg0NBJywmK/0go8S8fYZAA52yUUFVkFM
ch0wSXh+2v/P7/aBhastNi9NvqVfnroibkuJutMCghiTzo1yiBkpB/AgDs+u
Gu+2JCvVJzpGkDp6WUbHGIyQCFyh9L5M7JOnDm7tWo2eHts6ZTqeNW8iWwvf
T/MtmkfmG3xRPLfvCb3WyZtU+JaeybT8iBznSK+PlzFE0frMatHbBCFC42WQ
dF5Jmgan9nkrw5J6ZC/T3jXE2Ie4DGnLpomoaaphl92v7U/Be1+vJJS5l5GG
zq3DriWvEc6MpFqsMxfjDDqNaaN14F6eUx1Fgj0fCI2ZNXDEtgqe8RQ/b4t3
SNjZ9d2qRqkVtB6571KgVmlYOU+WAhY/acaMc0PzNwAK2O9zujx15WjvD5Em
aQV1Uk5a6qokMyL894to+xKDxwEoIjWoXy1sSBYrv8xklwmZlLktcphSu9gT
jYxxQL6J4OlAwJfcpQPPssLW3FJjAzVk1eL1i9FYptFhL/0H1hZknYhHwnhq
VSReKt73Dq+MB351pIaAqVGamF6jqGbYKhpyu5/ra474u1Ses7HKpvCoHCVv
yRz+WrQnVyeKoNjbLu/CCQPEV/cjCyaVKRWI6lgA9drdjtCYsTq7pqAc8sUG
LyzDFaVK9NkBpZvbrjhRXci06P2t7xlzf3zkMDJ4QLWPkJ5QsRmuyMib5849
hGUsOFQ3IPPhxHqy+jze3rJa+J0y2C9TNS2GkfRWILUsdgZjJT+GdC+yC0Wc
yYTi117WYlx1HqicUQK/VewoS0nDWgRrkuip9LqQwTIkjUasaGU3fbCz8IMZ
Kib0tmFUEtWGSxpYLrajyCURejIS++e4VWXFrpWfNUpzPVg3f6ZDDEGa1ueu
j06JQDg4gX9/iEtOLDxzOofkr/Q8EPJz1DwX5iUKh0v/0V04HI+TJ3DEixTa
eWiGLnm92wRB48DSfIwIUHh661ofswr3B4kH+AMk9LW9vm/56IZDa/lCawDJ
l4h6mpZjfXSngg/tAjcQbhGf5AdLMyALbczM8B5GspgIxbNLIrNLbrvEr1k5
4yneHMM5z9UbHDu7yS6pnINkOfJSGZrZm98Kb0U0MLDKTh6DSNHHvVrPrz+3
+dpjzE7mFdw84SyNoI/laIHEh9swxl/aB0CqauQB+zHpk51asxnaGSzTf6NY
I2R406L9AudFn3sCL2bLltG89Pb7Uxiz3trLqKoUGn07mg/gH8O3BjNVddHo
zIsivWAlRAJz2bcz8IqWOTbML+8/Z0E9YUCP4BHUSzCpmbMkniFdRUUlzba5
IiONdbR+0YgFkRaaJhF11yiQw4QxYTGIBZvgee94TZ1zXUobk3iXOJhi6Joy
U2HZHXAaopcrEBIbqmMmFOZEyRwIrMyTpRZqdroBeMwYJXI3/oeCfRgmXETm
LMyCT2HR+/UVTo7DzApkxJRGQzTlZrX1GLLDfVUMbyPmRb94qK5ZJPnaHKNh
JuvM4tYwz3Ll3pIzFmlc3qEZI50GuqdGWC8JrAjmeh8dzlSAsNuVvsv7EsCk
TXtOcZ1e6bX8xpatu6P83UMWDbJWaCvEzBKeakTz34GOx4jgIqADL3cgGRyB
nXZRPEebOldDXTdRGqaqe0NngnPo+DhIzCc35oIW9kbT/QpmYtzs3E3Ey31/
ZoORFff+S03kre22hbPhB6Svu3lF5BtOWuf1gQHnXPLGo29D85Te9jti7dcj
VnQMfpVHMxvHkwVB8X/ZnFMji5MXceQux/aQ2QW/3xZDPUT21/yieq7TbcEi
jwxFcNo2yYybLJ4vy2FpoaFZxXC+CZCxeY2Mop3lsNOkwsCkRZXmp4BhEUkb
G4FpyGKcYfBSbnG/bXQpaTJbLLQzrzuXAN1BK0cMMCMpZUYvclFEmgMp2ue3
uVEhSapozL3b1TG4hG00Vnt3znJBlnB3H5EgTdC/yCz8mVJwAu562r7Etfve
p00KGMziDA/V0hrbMpnO4V1k2Ecb/pn1djapPZF681bqs2LpCZrTsGH+ONBV
zeBAlV5GDliQyZROEruzGHfaHR2ahdk7xMDbob6Xug5AZMRGloerGY2boceU
qXJ0Y3xG60QsRKuHHGekM6AFMUNPxKsWRrrizbfhD2+EiF5Y28wpnOhHJ8/n
sju4yOkQl2lYPdarA+gh8Qddhn90XEExFYNUgf6wWxxY2cIOlTt00nzsqXv9
3v7+aoGXxjH46NUoIYA7k10sh9sSA7F6vm9XXw5GW/7WXqBBnDBT3C3L48kL
YvpwiPFlpTv0bZEseShdjkwaAKncu+JhikzVHF1bU3qrFstmjE/YeTOWsRwQ
z92SkKVfURAxQe9GVNNKixNZ4uFv5mNRROQrJT+mfX07hNGrTPvYmouf8vBe
81fqIQi6USpnlH3oT4hcj4lj2HfRABytXq/1B+FkSWfPVzI/x/lWCU41LoZy
FRwR8e1Vmz3sD+Z5xCRzZWI/WXG4Xmo5RV+AAicvLqmREcJAQLTqru83nvXb
QrKSycWscjLoquq+RF/IxX+eR1AFJlDbwhmBsBE8TwwHotkKGNDgEJn9w8QV
wO3GOJzLdJ6NepW/gwwsR6AsHsZ+T7Czw121fWdXwsckLluJo2F3u4vDC0Pl
vQdMoE5BXiqZdLvkSorJIgsRt2TER+1R2Vsij5t1FNMPTvpYOsx/aX97YvJz
xExSe+OxHuyk7RLDh6y9g55CGQ7e1A/pyS9l3e43tnmU0kOuHC+CLUSXgBdA
V7yLx0MHx7gIsWM0NCGl1Zyvnfjny2CeBL9RhOJpBrJ4nxhcAhriM6hr5yW6
kjIs40nzaANuhayoSKyIYWW8hU/Ed3KhFzzUVSVlE8X0Bzod6E/SAo/94hdr
/3vHBz/rQxKAhM08VpzC18lRBElsblEVyz7MCJlVdc3IYaxKtnv9PMI/L3hX
V2l/aRqUAP0JirphhWvq2+WZBHURfMAOMh5fOcMY0sv9J3rIiSQ0oFvb7P/g
caWm9qCVODiaMxw2JpANGGOJlgh8xGCgvMVqbbDUYaLJMqNRBG/nuUOeHcgS
7lEP59El48pcw7QMopaMve/xmRXEsitOacVmf/m4mJkmydMorwFaNUE1xFpt
MOCxZTt1ZE4zAkd12pcN6YviRhEnhuCqYLkcYLmek6ZChkak19sdPM1RQ74R
CmICtaY4OX2m1oKfAT0P5EXg8jHEKXWXLmdXTuYTSJT2HhERZqvN5gTxekUe
jkZ18wj+7A9yS/ICIluJwrRHHkKuxqnTb2WyjLzPL5Avm96kuNC8mh976yvC
QqmYr72ixen2X7606zhLNhhbYHKH0q2huMO8xPwrUZid3+bAXu6f6pn2NTGR
nmKLgPaxN9LqEm6wLf6jyRa7n/T8LNfXpg4nySsvz+tVSYZNzVYmxvcIYMum
oQzZJI14pOkSz9zaYpi/jE0bZ5fjmZLlimgoo32NY4gP0K61RoLapjkGWHiG
NjyDmNd1beoazsbsEtbNb73gNqNRH+IYqOqmqk2ys8GgmsF7uCib/PG+l9bh
H9Vz5B8DMA4CYZFIKaHQyqqWKRc0VT7bb8H9LCoGN0QIiA/zMLqDu+nspsgj
SfWqUnSiA/b8+EYXfsgVQsGW6Oa5R22xumoHDVh1rME8YiEkZT99D265Lc0q
TWC4dhCDG/aVtrqo7ON/rnZ34lhDpprGjsBV5qCnIpYzKhad7iZr+eFFXUAq
eCw1SWmXHAsbKUnkb93m6qRRQZY1bpy+KJKg5XTd1FpXsa2kYT5Xq+IAKFVL
VOCItsnc6PstyBhFACOIE6p8Hz+qE7+CoZMEXEVsyF/4gTUaBdV8FcApfHEw
+IXpZBwPp/oCapD+NU/y0tLj6O8We1aKUv8ACOsfBEpa8D29ErUsVHJjxOq3
+fXOHsYddpX+TVlgoI69oRsob4XXhFKYGisrl1z92nJiFIh0wCuM1CzJU9EF
8IVyEBmeeIB2FrU6PlL+MbuPLcNPCT7OWMrYpj0zwGf7tO4SeUZ4NbuCM3hW
V/kWNMk/BCWrR+oE+Ag//Fo/yHM8diu0zrTa1lXrWahP9V4iN6sv6NaxyzvM
4M68HC05EMmqXzv8xsiw7E9W1pPKGRfcAJMltQiDfgeD4irZRm4qd/E7bm75
xd0L0q185rutbagBSTPeeN4VJtbX4ENZqAbdgHI+ksuGxZUBQO2cRHI8uTjq
SFnV70mpR3DBQ5b/M0h1MR+9EObCCBnb4/1kgakodkwhVAQ9v6TNbtLvOiRj
J9bFvSCANx7Nslprvqxv43kiN8IfJzubyHL8D5wxLROD2zzjVNFA4l6K5W7G
/xWeer0vfBcaT1TyQEd0enO8lrPAuDVuRRqm1kTOB+Bja69Uta5BNXkfRpb1
C72eO+A7ZVIgfJ5vlNZuEUZbGWi85GyLVryQdiu2gheJ5CRRQOGT7vA+J6C7
AR8BEzjW9kv3FX8ndt0Pkq5ncGR8Qlgr//hlEEAppvXF0OtXzSPSB1qf2i1S
A1rlK7ewHlQmU6oAcNCaQ7g1JOVcg7oMQuZCuDKsTMvkgsI8sOev14bkyEG2
2skCM5y/Kj+77qyvtxu0t6f1ME8VoXa46LYLSDOi6wNWSnIF014+jszZYV/S
JHf1Uy19cn5xUFJ4YRus1JM/GPKpTKzex2/kmnKMQxgxUWy0jYDpMmPuqFEp
ueduhjjIX9yYMbZ2pTLU7aeNMUDqtFAL2P9vBcKRtvp2p+wLU8YVf2DVSZJY
RblV1AZihS1hcR3U3zFBRA4Rk8pgMMi9XaUEhgBqlWd2gXNIj8rr3swDKa1K
+0FfH5B2TVq8Pw8QDS3f0nETy3IUPVqI14ZoAIBUtlQKXB8v13U2PGsqdyd3
6rH3MUyz/RMfNg2ZfU6qb48z7fmosSG662vdGinx3gSaeDqkQKMycwC9ex/E
8CYR95OfbIdmHw6leYFLnYLB33VFfR1+V1GfjvGFNWMCE3nJbQ6qxF/HEMe1
yvoW69EeKzOWEpWJLtRqiOVFbbWJWaQpGUQE6eK8HTBRJPYbhpv0uuhDQVcY
tb+bvk+yZZp3gTB7Pt3LKQYYkHkMZXumOtmE2fbkn1a52Wxnb9DP8qt1zBd8
V7saXEcrueGtpj759rTI2qpNXOVy9SW7yad+NhNVUkdIVdNrc4ze7EsFD4FH
Tj5cqUVsG2dX63RipKddY+4yrh3k1krI12UyNOA310U2otFlkBm0eZvHs5Fl
B8qlxlD26KdDcVZ9t+vySG8tPusMKXTh1Ow7pPLpbSn/FhhObJ1Lh54t6dQi
YSdy2pP8PQHIoi2r3PoMrI6x5hQhka+IqmR36Z8UJ2lqNKVqzLdS0cyoaWS5
2xowzxDwpMrFNXPzLjJD3fpJAFJUv4l8sNIUERgyCU2yRmmNjEOrdrF6mkeE
MIhb4Q1FikrdEf2mqqKYeY3SiItjnT4tG4VRgstPDWqQNqe2+LuTcQeoTqTG
OmD8zY12QAddWfGppK0fZ1y35YhyC+N/NobyfsA2IeTA6p672CCBZWKYE66n
WjKxMogV6pEgGs54gh+xQtyLIVWNh5mEN2t7Kq4ePHhTEcSSeDI09yk0ACSz
eZfY3UNcUU9fZTdUVZMQ70tuBkOJa4GpmyhZ4B/dkNPQcOqsIFn3dnleVfX7
hEQqIuvaGJfzhm/8Jy7KogV8PQHBqeihBBkBsbjbzmJNorqPaT515CAOmY8J
2QunElpLGtBC5jPTHjGlVrxkO8qjuCPl2/5i1kie0w+BoWvUcgRUuHRUi+wu
vT5rLjH0osQNyqMZLiHexlro4qY7zLXcxs7mhOGLs8fSgLTb8ZK0rBN/+eVw
OpCx/Fel1RDFuhp/YFD1ncOIA1j4yENu5+CLkSxkWYWs/Rj7WkpVDlwSlimn
IeE5r614WEwfvGKLklhmLfvLcT89af4dHN6cD4CE/g9UCIh2AvmIF2AwbkpP
fI4To2bHiEV3cuO/V8Ts76/D/xt2yIQ55eaEFlUkUFuqpwb6HIxI9aYQ3fOZ
GTgUJ+X9AJyaBXvGj7ECIRS+bTvtpCyy9RYIJwuDk0dnkfCP2aIiXreuFJij
TKuOYBeSaUTI6slUAoG7RCPNwuywlK5Eh9e1mL9T0Of38BwuWgEzV60XY0a8
w80PuvkjsGGn+h6YIDq3Sb+qlQOvBuuCHaaaIxCeH8REVP3v5OI6z2KnvQUK
M8ZlwAf5+jH3SFtipBkFNe8JlJT0aBlBydKm4KW7iKy4EMeBapJH9jrlnOJw
JidweRhFrcoA6KJBj7h3wJlxTHT80QPhjMmwhxt1eANk/rpOLdfFRWfN1UtH
XyTGPW2fP6lZzc3B1FRSUMuuIzGKN67nKig3WiBYHILF5BA9eO2NTSYEKukI
RvSCc2+xWALuQQ952ifauBVeLDQlkYAUgivVqJsr7Agu1e3FuQ/MYBVD1tQY
feNiVUClDtb6Rs8JmULoU8wwA278/0TbZGqryHNT3qSLzBJmWjmF/bs4P4Nd
1Q4ND6pslt931D0VGnjg2SSIcWZ3YIAgNfMcbEQ5R+/qjj1ce7hjsaAL7APz
SIbRu2ad1PuSn0sHGXHHdOw3NeChcBEgHUZS14ApWbARfTtGIaiRh8Jlt47Q
tdRvjyswdFShIgkv3PkIaGJ2sn1TQF7eDn0/TkoGbN9M5XibZnghm4VAERaI
IIToSSfiby8Ojlmt/WkoywYA7xq8EMiDURdLvW5/t7eG76GsLOkg8LlgPATd
+5CDQ5jahd4Tj2T8Q1Q42YS+hXOel5oK5Ohj7YS7yFu0hixs9XlUo6huDDFo
WT+CpewJc1imPboLfnm5UzUNw98VlYVcftNe5j1DyGk+atE8osFZ4VpjgMaq
CffdaHuou4ZcVb64WdniaJr2fkr6wtoQEh2gzo8U9rEpAPYsGZSdp2TyP1tD
SF1U+5oEANSMDJZNdTAYsL2TC1gLktJOIw59Um831aglLWyK5pRqxGrkG7Qj
biem9eLfHeksHIT71wgJYGSciahpPy6qJf5ZKj+cOBw47PLef6LvQMd9jaf2
CCX0osZoqbV63WOWuw6gEpUZ7hfLfsW/XlW7PDeatJ+9Xs1pedfui3pDeBLD
XIJ5rtfFCZ6zKh03QMv0rjnXf1s4M/QdCywjwWXLqn3LMAlT3EnAZHLltdto
eFVzrNDPxaQyS5OgZICM9ze3Bz+l1nJgY31DsGoCDAxkTF9dtJdQdkvjzdpX
9T00DFaHrZUfvEYt7UjTy8uMcFmYLVJetVhJmyRBam1WVdvntIkV4lUjJzx1
tsBVlIOnSVl2MtYIPYHD80aXTVTghCjoTiH6BCh0+vkZt99BO2xdrRiq1TgK
aDG8CS1hwT/w+Yg+MemUa15Z3WRTb1Gb3hEtNaJmkbh92CQcEwFP11k5WTOG
E/IMNjVHbncaPUol6VDkyJG7nw2l5dqF8W+hy/i5nGQVuJ2RLJHJQtubAN1d
68xa6ryYqoIyV41E9qqW1VAE/NqMFbDfqRx3qW5qn1snRbK3WnyYasgUXUMq
c/yJJcKTHAagK1vXzHoTcIPas5Z6LWBlqW4Mc13ks04Doivlmon3NIKEgZL/
s13zlq/PbiuaEJ05rMKZ+4u0+StwOSQAtlLXScKWXp7O6PbuPg9/3/+GngQv
lUdXCiZX05ub6Ep2npDvYktZRs0zzRM0DFra9l2FCv+hC/1lA+sQixFHzJgF
fhST/1KO3DMVo7QcDKHfQoV9ysmrPOpYUU/L/GrJoe1QQNXsbFl2wdabw83/
A8wlEtTI1zq52V5BvTIIuV3ulbR2T+yMZboJly5X5LoB3G9C6Ja+oSxBY9Yx
EaHBsCw/zjRPOeKpLmUi1JK2XKckFE4yy8ry/Tyv+leJLr9PR3INDPt88//a
7D12w37JtolOda7blM9cNLjGq1TR/NRxFbJLepnomBh9ApJ98qT/Tz8Vq8Cg
v0ZveptamEnmamzTm/lZBXok90kt/L91IweUWViQ2c67DrWe9QYvqfoOhNK+
0lX6F4VVI9CHd8ceeETy1cu3P37edHIrmZO1Siytf80c9PbCBCur6aoYG7VU
j1RTu0prMaDrCHAepp89lxn1jRygrrC4yBmSNrCDgT1MB1OXaXaBSfaPSv8i
e7TgRX1v1g5LPMrGinSDTopsIQxD8SxRpP4kkGG4wH6uYoZg2xYmbz5VkE5x
Y5LAf59gc0+Em3hkI5SKeAr9NVGKmwPXRKFCs2Uy7NmwxRGKGid0fczS94HP
+5kSceQqNtZk1dff6WIee1uCloY8bpBtvHSocS9+MUYLCbFgXfrY84R9kXj5
wX46DA2EwtsOnpNiedBd1Dm50KWevEIM9Fp8UPlQ6f4+YXLKpwOqO9c9EOtA
KwQSDrNzSXvJ5Dg3mRonAXLTyzz7bhyFx+6/IEwxI1ezeY60Exl6FQKmAopn
bCmlIflFMeKjvZUk39ygv7HMOyr1PKr4FXf9ehZJun0aY19u5WokyJ/eXSMe
gyvieId3V7sx7pla6Fxys1iu2wlqq3vY0rtJq5ED4XOK7kxhMk0CsTnzx7to
0C61JI4dHtdUmxf8enh9nL9z8jPBxdkrMorq3L2gjftWEghCqDj6zmwpDlVK
Q1Wx/D4XH09eTC+g9A0XVnTJyIEsusW9lMs5wx2XTXjypSSRJYEDl7C9Ncgq
lTY5ky3gwle19OuQOqqeO9hh1GcFQf47RPsOCB3/g4/R3rtngWLkDaDnl3Sn
65vtKskxqYAtRZt1fwinmU7Lg5sbEQxqjibPoU/7rRBYx47fIngLv74g3kO2
xbv9H2wqsGZ8zZmEliuhoxNPxtaw8wUe9XIcEpRFJG5ENuBPlODI4Bkp7TCM
TGx6Gn4RJ6/Uvo3dh4jJMH9ubux5sITHzq9if0VWtlsYWf90UBj8Z4cdeZkc
TeR5bgLicc0/PgnSQBG/E2P99BpoQBqn59Xi+JjIbfYvdDkoB0DvsiG2di8q
kk1gM3ersLabS7xrqxstIEnBheYHo8HtJXS2rFamSUzzpoC1b8OaIQCqO58i
rGCAlcfsPxUlAN/OLykqq5Z7XA8rAx0IFtwPJgukP1+Xy9EZjCpdAzqMxfzS
3ofskYDmestBfjZkBrCdHAu/3+fmttA/jdweFOVrLKOonvSIfSySlSMJJDxQ
p1SueMC9bh0j21R3m2/EnM1RUP/G4vf8/VwRqPS45vt3kn1jmkHSFcLcJV1+
yaCS1F0nBtfmvtvnVCsAAOUtxSSQrqVmqJuGveSghvjO5pzzTGIo7zSkUvGc
NWI3tSum8RI9SiaQdO45v7hwunPnXUxdnTQSm5S5TTzVe6MxJjj84Mv1JgXb
7LxzmvKDYiZAk7SHj/ZNkpJFFI5sULOopAOtNX9vsYEQpb9G8azJVQzjW318
E2AtzTSgDxYluzCTPrkm3xlEINWLVIzHJluhOICokjwCt2ZuWQfUcHR2SKqk
b+UuUmthUJWXlZzUgTfZoWngjwsUQgLtOXL1BgI63IPFlmqpUGQgekXL4Ngi
Gxp6Pqex29qbVJf3NuL4VQXL5NqhO64o5cbny9MiUQPp88OxVjOAUmGEMkU9
aqq9w5OG4d/rczzQnAiVE9KOMXZ3Q0QtYDK/xPxQZoxJzthbrh1Ld6N11o9E
3mQ4OIPqoNMNUnuc7QXxo5V61mtWcmfUhDIdK3S/B263OUckzy/KmQIi5t3c
BSP7HbKvuLNXuPU3lpYFRD0UA45VZQK9ukPaLY+Zd5LvvR1jRveNUJ3KpuJW
TgZpKNHv8zT1zVZnA7IXH+GPM6RNDsU+2Zl16QAxzBcQPQqF1wSiQab/E3UE
s4uvNc/AAtxPnUOIaui8ITtvLSr6kmnVna6VGzosr/js0d+3EUma82wSi6/e
EAQ9R5TxTULH+mmjaoGjRZlQSJvst2d3GbokzYNossj4mZNpi2bmDrrlpIUC
VD60WjxEEqhaLImx3zyEy5SzP9VXuRPQDlRFSMzm4eUUNTb1psWGGeQgkuRJ
0eaGbvLPnQnbnA81jGp2LzitrOFcUwJcKb+XC3NUpYhP+hGwUGaY3JGKc5Az
dm81f2FThxK9s0MFNybSB+LUNWsnQT8XL2qHcpVLR8RQimEf1CcsSmbjtqdw
2wBPZqeXuN3IpUH85turizvwgOA5W43WtsJGqAkfoTJrG9dcTyKYhe8au8Sg
e5KX8G4FzUT0OhnUxzKRhYL8b9waMmrDacwNz0rqdYs8QLSdHaWTwsV5lH6t
RfAJEmQn7X9h/VE9eHgdHK0oRLSnJWkttU0rgXO0Ul3rHS5oFTa0nheYFZCL
odY/u9UWFx5gfwg0VsDIzAzSTqLWNGFU8ZjYX6CkxANwDXfawtLHxN03l6i1
bBH/S/4WlB2XiWex6YeKhuJv+S9V1NVaNbmwNkxtJ4QPF7pG33F3QA8cZBpB
O8aRbp2m/dZjJyHNAa72KZgSC5VZp1m06ErGruiiHfyDW8WV9NG+GfNi5QGz
iIa1pFnjNx3lrRwR2pwvacptHYFMVsQetciOJEYooiIse3sq3sV2upvNQIoq
IQI7RcJGO5KCrcaHgGARy3vOxpRW73dBh69Em9/uhZ2NRITfavsfVI3qG/mj
hzNxl/NQu0HmTb2WkptgVGRXVMu7Md94W/UBtKa3VDQUN16bLA/y7IFOVFxC
awzgadyH1XIquK+mMO0vFweycs1ytwUhgw6GBbMRATDZWPHSYUWOJEPvhKfK
GXOFtreXmTSJedmHX2e+xnA5HxzsLV1OvS7VRjdyfH8ulXd47cjXD8pXm3nS
wsncEtFoGiopmpYrteoPvahLfymyh/rHIIfRnQq9CZBOg/HSb3d6URd92yFp
dh52+R/0gPUS9jqycLOXDa00q/tsj7kDgpI3+mv0le8jzLCkRt9gJHLm7+03
78xLdibtuhR0M8hPkZVa2pKo2mzBpVdqh0+lPiBtUjA5Noh37AfxGM0Rrv30
nnztbaH7w0ubogEp7Um89/itpjGjyK11KXjSrKCN70YRg0UUFy8mansBtPfC
xg28AQIqaRFdg2NOcdfe4QUDHoJvp6SUSBn9ubDrpYQckfbBQtnQ5bQ28+DW
OK2qc5qoDQ7N7BTIrMJSPMN0Akc6IeT2vjjEXwhD+poxEN1AYXqTb3VdIkB3
xly6q9ClpYLSE92jFjTN/jobm9zyxSwoqD+ZgPDu3+ufjJQyQM/Q+zCIFcnO
JKAKsAN91vKCwGMO93o7LCdn8FuGms3jxzAg4aWMI7Vf/2jJEBm4xEM+2e8K
/c108TxMie6MjKNX+dL4V2x9Lsp+W/E3NtZwc2iVyyBJ5uZnB/+xTXePE3TB
QQnNJLn+u1HUdPt8wue4CMAI3/71bSX4ek1RzNAyZMHQ24VGhEbz3d9jRCRN
aSlTCLb0iXqwLWwWdM/shZmP/9cX0c4hK1GnUezY1Q1RkRYNfOLJufu8Keiw
/6aJKUbp1pBOEUbwbdSXr3y/6/GwOzIejHVUS+UD4eV/kVtL8nikQmUb2wQG
8+F4gUnXyO1jhhZwSyD19InJ5aShHWqxs49vfKDZvYl1iL2a8/4g+k13g6BG
7YIo0rJsllycVcb7IrH6pDxwHlfvgtfkEYu8hzP/usmgLCpW1f/NHO/rIg6R
g9msCuq67aTvGvvmnWbehXICk4b2vr1eCdtiBbjyiUFZnZG/RW3AMO58OoPb
FaNriDtNdFIBt7WBluf98phMziVJ4ArVqGO4mAucDBZ9Sp2zOKMTYjHZnTID
591AsTPuSseyNgOCKUuSxK3cuKm23qhf19XrnALZ41wjgHF5i1RFPPXJ7gi/
idQZVhp4j6j8bZsD5QZ5cmAHXHcun4SDT0SsrhrhEzqWOZi742vEzmpmljk8
3RwGLC5oNyoLHunaeaUFIgIni64I4fy62bO6cQgcV628CeYBsQ9t7GzhYaUG
bwO9ng6lZWSPCbzFLKayXhdWlAWCFRzlcnKmAUUcabvXIeR0WbYrT16565AK
uALt9cKgkfHzL+oV5Qqf+ROH115VfPV2rnmmvLAR89IIuPIHoSgpaFSgpQJb
VGQDGvjDgGgCEBUzBpLfLeRuJMHPeJod6cCOjL+vc5bhKCQHFZBOFV8XzL8y
0tvM0iMdSfsxMHuE6x9GkZBpI51BoqSUAuURFU0RP1kdmWGiOTh6q0OWl5J3
D7ieEJTrt4eOqY+4YtXMJA56pWPJTYCj0TJdrcqSrx+6exq/PhhL22ZB9eW/
hOyLHyefok4q9215mgZs/ggYJaVBxyIEUfqDOkmlN49J0wAZe4vi/kbDVBW5
gb+s64qFaOMNk/ZDl6TxbB9eYhI+vcHJtiAEm5gh2Fy1eDjhwebFB9rBeSVC
dmJmkSpMOjet1wZaUtsbuba+BA8k7wISvC2ZCnsKUXVPBHK5iE9JvL3vGTQp
rYmVEds3Ri7AagThLg+lLq4S3haL6gv5qDwVL3XQ0BNGAtpS5jbXp2ultB3T
c31qMKH5r2qFpTDIVejmjjoGD5G9ON8QYY06CjLj30x+PN092SVAyHn3Pe/X
TjGk4oop0RMi6JMLeNJOye/MKcgGD02VJ3+3GCOvM12HaGTIUUpbYzH0exu/
g9fBy9g4C+cgowKFAoMhVqJCa5meU24FviYUSuJmzAKaDR2TYHZ+/IWCR+mE
IK1MvOBvezQEQNyIDt+XLD7teCSOFgo1xw5W03Vri7bmght23wJOXQ8qwr3n
0jNxRzwPzLWjsWMs/YcbbmeOou8m+wMndS46w8cAZZgDbdXa3HYgdo5nFdIg
tx05mGXvB4Uh/uK2SX8pDWn1LwOUYzZo3afx9Op/09G1SoKMHvSZjZgAWcOB
oQI1a/FyLDqUTjBjilN+9qRpBHB2snCnu8dQ6MuaPowpwdeTjIj8vsgiTHuw
djj5fJhedt8y9QT1HoKbaTCk4OKD7zWkBmo8gERQ4bfWO2xC0iNhyA7ljhK3
2Bm6JfaFIyZ4LCPLqcdlJ1Q/Em858+sEjRulWjToIYphYaELsLPPpU9GjKcd
BSC1wGOHo1Rl9REMpOP2Dz0iT+4nRxMiN1ibb3O6EKHUVTHWzfNC6sdC+6PG
6z0uzoLxZw7iroAP8jrsngGcxPpFZVg3z9cwWI7HzHNNcXVXI7mG/GzAqFKj
ybfsfHqIeOnduj2oZoAzlhTPelvMs/VaN+/SOEdmHSTXarQxx3SmbBzJ/7ex
gUnBLLqoRlEZu9iu1Z3nLWE5UNYgjcI3D9QR3l1D1JqK4sHvS+DcYyTXlpHu
UHjbhXdW79DKLLAVMbAhaxo2OGTTg8QZgbFCAKq07hh7gkicjR7amZjpjVVl
TwI6fbUwG0yZFXw11CyWDMBxNhy/UE4XtGoeTLv0hKvpXs47I6Ps7s9LvKnk
g6QkLKsy9qKiJgFF+tAlQrfznEbkd7eR9mN+3Jo9A2GN/vkecB+i5+je/08y
wuCmKdBbGgj1VcNdiY8DetCmehK73UepEC0I9pkYZGofI1V0bO8ay0U+dvSb
8cHireP9jx8KU2mc00WZstlC0sKs1wVZZNGK4FIpbCiqRVF/zDTMCpFIVSVk
GwVSv2SW//9JXb9voOqItRKEqMNYILO7uoTgVWS+btaE3L4aS+4PAMYudzbQ
AEThQW9XwSVIeY1eM3TGpblVnD/rEI3FW2eLG1FpRn9TXH6XDRLHYNg/JBY+
UY7oChBB4RYxfiZvFOfAdEvM+T5uhFGaVmYnqnA9qKGjRoLn8Zy5QdBfDSl6
CpPY7mQll4yhheP4wTwY5S6SSZCoYlBVXUmXwRVHuBAON3fUIZ/Tx7aaOfcQ
YpM+5I5N5dUKBN61y9LklSijYrO6dkRhufsUNRB4Ju+aYhzW0Vw7b2blrG+O
jX68LZtF6nGg/LWJaT/4Ti38flVNfulmK1Xg+4rsjB2/sOfDJpkwrhy2/b09
yR0iy5Z1IDOitzfXMuoFVV9k2w5BjVS7EoEvlP4Fu3bZfCcgaFPWMREUxuNx
tbWFJW8rehrUy4SSfTIzF8ChQKhp/ySjmMcb7Nm3QvX9hGHVip/i12Y0S96s
AZyUeSqIY5FLcJUXWUKpcWTudhAevYk6IHSgQzyViabd0UI1rRBx3om0aBFe
sJ/DtNv6gCDrgTyrSNrLV77Yt1SrTPNy7lJpBlv29gQBBNDS/UOmvCpBo1BA
TS3mRvH5KUVsnOEGfJE5WRuvzxtYO6/3mLEKAFDZnEy8YfSR5Kxgk6Og865C
wUYWhw1JMFTuEUCUf6QMT4mbHwFU2oKxF9lndqkd8LRzwD05m4K5RTS+kNEv
iTexyoWkOT0mCNV8ZHQg5q54K2pyK7hBMHi5/05Y8hNM3v/KjHDbdoEOeAgr
awC7to1umJ2hiIM3oPBolxlYI6GAHeiSVisODU0J5WXqWkQN1uHqZGamQJXt
6hQpZBIT+YIFnqyifkF/g2qcem41odX7XzlZG3NyQgcjCm9HguoSTlqqumPS
hSqiE/Z/tBsY3GZW4qG++8ZEPiHwHFPA3zeeooSxSfB7JUFZK5Yke/fhR0tu
2YHb0bQSXtGcK6y7xzokm/USPAnlIQi4TH+sWaA+oJ9tKjGKusIWKOTWdLAC
SqIUZAsQGGSrFha5jOxZ3wHicZg7VR8XEX9/QmV1shx+ZoSVgjOqn6XD+PHa
/SxEbTE81o6wlgAgYNSRLJfBui10AOGtrB10+l991/s5N1aTcc+uDjZx6MGr
oxpxDqTpMPtsb/ifYaOgVmmuqQLsfqQh5TcrQlhE2E9SMdz4qr70FELyGtww
eCBzb2B9eqHsvGmoS0rbTQoNvw4H0pdTuI3ZaQdmIEoczGILWreif89OYUR5
s0ebvW0LlBtwxYCQsFwTfUz4Wg4bNVLW5clecyDbKfQasHddc8zj7MVj0her
t43sbV0p3cQ1C6H+qmltEUt8yh0HaLK+TsT0FIfCapxQGID0ykyJ1OxNlxrI
9/sh/uVIEMXd18HIhYloYQ8Abb4uSV+1+5149KWWmqa9SHkEZtKgNLltBRgu
kCcvZiR9roaxN37DGKZzzV+GWZvpMkXGz0lEf171tinNOkF1hmoE7n/nlkvS
yYAQL346LqacBQ2EDl+kW3sCeTCsEC8nWe4oFVIx4pRqF7O0L8bNx7nM34Hl
T59Pr3XLHnXZ+/BpMbSBTshpv+ywckX/je6eQFe0GOJcc71XlgKfS1tCP9c9
3PMvQWffQ5izGxKMdr3epSxUd37asgayYL/mButCk8dTNUIU7WG+IRKugIyj
ataYVFTUcwGIcEr0Y71COnIQkxVgt1ImkGGfizY5niQT4N9XTLsgglCpj3tY
Av0FhC0oqIZJ+vOtDmVNjadp20R2s4wvOGMt7LUEUj7pm/oxKMZSGVc2Ntoq
5fmbaWXQwRI4H+u+/n3+qmaSb2kWg5lAL6D9nQ4hSZJ0U+xKuvLTMLRn6VYP
3bE3ijI4fxvb1z9jra4yTgX563yKdDYyrtYO5X/LsBML9Rd6J2WhiblqWHs1
3OLTEzugcKSaBctagsS6Ra5+Sf5+t+oM0k2atUO+6CeKWTfD7QY2gL9XErFG
GGpJTCUprTTqzSlze7E/N6G6fn3aHYoPAyG83sHctQNJjB4lq4ml8gRh658o
DAGW/YYW4iqhMAA5h/7c/yVXRpja7RYI2W7+W5GCcgo52SxAIPQQZjfmdgCm
mU58iD+jM/oqdjcDxVzJg/akfzhZ1Wy868neWmLBZw9bigKnlr+JXgbKtubJ
eHogx2Jq1hh5i7PVbCvqWDUNUTbnpaO/BFhGSFYqJ8VPTIUy5mensCQaAVt/
ziyNyPvDxucB6nlZftHj3YU1YpdS34mVWB/kBR0Mw1TFreDz7ivhPLWnefS0
7fvRh92wDhDvPaaLvA5gce+KlGicu+ZjCSMtkfVkzeACWruIsLH9RG+OTZ/s
L62pWbnZBLvnbOSKYokiPdIwPU89DNrH4vW1vblvLrKCJjKRmAD1QlZCxfBg
SlU/q/fqvoujR0Mt/PYBhcdzwJryEm7EwsgKbX3JXYz9n09pq5ItwdK/QZr8
8HUmU+/5+VmFt12Kmcl5cl2dNqoPPJRKiNw9LWOvro/PJbCTkl4EVtpgBTDo
xEJ099EUCfxvHDJWmDSCDUX9t8gtK8ly4PhCxdRIUUXuS8rQ5+6yVKGDJqzJ
SdjnnJlYs7cApXJfQJxXgqnkdLxLMJIJoZHuvfqkDPRe/H5WXGanafQ+bJOE
t1/KUrbM94Sl8jiaCVYVkRfI957vmIGyZjMeYeGT4xpxxgsDFCBfX7shzKfV
iASikhui44f7rjjIsKqS+w/h/qr5IraHnXTFJ8KvSw0ifa5flTv+MLukRVzx
obnOTqjonlQNm8z+YU1+YciUHwrZ13qgHBytSo0SFaR00FXm9oQZ09dmi3Oz
PzqyPPkZCVrKzGSr0GYSlhp+Ye5jepTOkHg2nV57QC/fUpEaT5TSydT5GCVt
y/3Vx4cIKSYVTlcstNPg7rQDXpM3ojnjT5S0dOM0upqrI8MlMwV+4g65XSDZ
8F3FISHKk8RfJd016cVUd8HGdrYZ00VOGWpaW06k6LZE9Tj/ih6gaRc9j2mj
E1Z+gz9J6QLvvAts+avrCgwIjGSG8tfajTa5+4zikpY4iC3PrquOnlBdINey
VxktUqfkd9pTR48+GU2yK4GU+yF8Sv8z8d8x6ALZL8Lg7oRut1Tp91FUbMNM
WEmej9hzLPD6/v26mD3TvA2zvPWrDbygiZ23T+csf/miK5bHjXxyoYPJe0Hr
/hZAmJOjCVnwGdonapaP2Dqhr0xDAwIXAaavQuwak0gIp/dyPgaWPtcRFOiW
TBJ29Hhrb4GYVa88YKlMJH1chgBRiqpsYWQ5Bh8axPBvFoKf8a+W2IkOqWLs
pI0nACWEevEQXDU8Z41UzcnfktNB3p6/1XAtoL9hRwl7gObusmfu/vnZE243
WV7klv5x3QiGxSbCajtSvGJiUp+k2f3OHIUOSV6OtWDLjizLy1EcWAbD3Quw
XZOu28LC8ja7wwbkxqTGxMVu5MeA5iO6nNTvjFcrH1RlDWSJYcNTHnoXjY70
zkqgLIWiwsNanOKeSurKmlOpkL9FFppc/QkB+U9Ws7JFzt03JLmQax2yO7wU
Xo1V8D1tZKEPRJ8FEUbbsxkjMpby0Td+RzJGE/jqd0vDLSBx3m0eB33i3axp
R/QiOP/TzXT93oZ9QizGpR5Y1CLHtcZgq9UJeRX+4oWJWAtLaE4yxpOZQquR
FfpxFHOsRxxsaJ6v106gMn6AkGgkvQUeGUy4uPmljvy6f4RVX58EGbs67RI0
kguHdG38wGywzLjQJH6AuSI0kKnwNBbe4nMj+Duz7OCDKocmAX+xMe2Dq0I6
+HbAlzrKEObUecnY+4mI2Ih8VfA2v/vWU7ndSLIrsi7Mzkcamq2aQQJvKFA4
jPiaI49RkoOE2FavoMUOydZ+ZCwpBoM3ZVER66LcUiGqecvcel2lbYidbGw5
6znFSiLaaBLeZa1OJjgga6y6F7PXP3KZr+XQwqIph4uv/3x7GiKOtcPZk46a
3wRv/f3QfIUCllxb3bU47WD0mAVu3bBRj110HoaDWKHSyMO+RUpu/+r2BEep
rJDukWuUyz7XNl2Aj2GGxaB8Ubia1HnqN3eP0E/PMHC+fVG8LrYmWkZjaL8c
EkTpZpkce/ESFF3YuuljGfZ9TDx8auCNRAgG781U9beAGU4uo8w65bdc56Yy
/of/eFrAj47O4Llayng/PlnKAWVD0saZ58vUIXm62vNo64DxdaPxwyP0efCa
9dy/wILOeHmeLc7nOMJN4A4lw5lfg2o6tRwPMhqOi/TA9XvzJXZmnQv603GG
T9TKrXgKEcJZI1ms4uA4uN/ahftuxRf7cujn7AX0CT5SdUJhsBMJeaYbOAEE
ESPgi6qOoeH/K3wNDZ4Pq+xRZX/AJFqBsUQjPtU2YOIhjrVzSNQkR+7kCOlV
vFXy1LE4PEsl8/YjMlSz8QGk0IuKryr4N0gbHR/rzpxVJFnm1LiTH9jNf3lr
Ux5Y0T2zthY4U9BtaoTYK8Xp4F9KswA/8l+PI0TaiR5K9jkH/iZfxN6tCpBN
3vZ3EXa0RQEv912gGZjx6PyBauOs0FceDfchikvWvFYMd6Cm4GWtvXWeqaAA
yHNXlZ2EeLv3ZEqUY95dfRdySenmtrZ/9z2yJw2WfGkXiXfqT2VseLFaiHTD
nJmhA5FEjVqkuhtFbrqiZvlvp+QCtQQJmLG5tH53Cj/B11WvtIDKFe8rbEz1
EvwAVl/X2KxsKShHXQNou3HXf3NdW04hywRac6AfN/gEQjebB02z0NTjoL3K
iIA0wCCMEPxnMMWaiRmlD4A/2UB0K+su5to4OSF8wpmGxNbaZABpEMdPMLLF
/2Q6oUvCXD5VFvU9mASSKJdGI1eQgV0Ssd2GFbmK7AU1pLMGpcmllzdwNIt0
UeVh+0TfdgGTjco/3ZO/6bS/ySZU4Ro6BgEZY8Q4s83rEd1PbJeaWPmYgfF4
OdQJTZbkx6Ax12YcLZK8esMNVlt0xmWAhhDEDN5JYsMPK6b+lKhlyxAKvjbr
Q+4eMZGc2GhkYJlpEe6dq+ZPg6TIUZmmp37qmPr0N/pan8Mr7wk67CVXQDUk
Ikq3GL98P5f7t+PNKEE6ZrY+lNruExzagd0hwaZGb/lA+6WKRk3OWrehAEOx
JmLFU8MMnFp119E0IVm3QqnB7xCaFKVJifaO6tEmoHI5COAFEHws9o+JTCUG
A8WqasFiSbK40o3kIF7rJS36riSmYjGaQjw4xHib32hdh5sp4oyv7YcikBwR
tOiVyuthqgkNF3TuwRD4lxJ3bbIJ9K8NwsTRIuyOgr3oxtLme0/C4Tj/xwii
6hAVG71KESudsSU0690tJuP/CDPlYIujvAVMVzvIN3VHUhMjQKPECexqrpfJ
Srg5AkVnblF7qeAVsNjIzZ8Hfm0s6SI0n/6ZlQ+H//8b7BbpjL6a5iMvbdrm
dLfskEn7Nr4ni8StZrCWhtTkPeDDzFvkmB3Kd7krmdQXfKbWVWeaPmJcDymT
jpCq+V9n81tIwz/5VJeitbmtdAIKDK1b37XNfpsgHbNF3ve8KgDLxHwvsrjc
Xm1aO6znHRwmFzNxxBNR8XSdPzFsozZLnNqkKBmXwtQWTMShCkFo5oOJi4us
SHOhE7ghxwuz+2kjEprdfUu3zanaoZfxSdlNOBjQr5XMJwtIC2O3raWFmdgw
quVEoC0ZgN+Mcdp8Z4IiW2MHRdexrUXe9SAfbP5wUtg3H+V0zYceLHAs/QHj
GuyQZEs/D7RQFqfPH7cp7Qa4II6m2QHVo0HkU/DscqVeo//ZhkjuZXs8YJei
u8yLDKP1oeE+ydlxHqperlgCmHCG4HuJwkh7pgvXKc6gbg5rACmN9TRj822t
XJFkwwhJJsIc+dA7gEgnxHG/8eOFyh+hxaQXkT4GYJMUdpVyLfP3L+XvJobh
JpKu0hByuxRWKXmlBDVEGHBPwBOB7mFvw6C9JphS5cNQ5wfXDyjtFQiP2hmE
/QkXwl3hN3JSmC+EoFideIAtkXVdgAuy1PG60NcP+rBcZd4LozLlUSKZhBWd
pa48Z9JcspGSKTJwfmTu07DgweeAI9LSm1ObbSZNV3K70vg3C2lO86o11rwz
Vz8AwunZqrKFrildHL6BdEBBiT0TaEw50MeeiEbPRAWOwn9flxgC47du5lIR
qdjxyWcr49P1yARB4Bcw+gdYL8JUiqeb+PGTKAPxE45rP2/5kUD1qL5m3lio
OXLK6f7hx05GMIIJUQEnGXpfz8VbxOoo6VYl9r/HAdcuw2Yx57zqbUVwW6tf
V+nuUcFcVTLcODMmj4BCOqOhBEmOdLGnn+rYE5OIstavdUQQUY/Xh3RgrXE6
V7zaXvJH1TUUesid8qNtsWIR1sMdXgYzUQDO0AHXDleVy++98+W2mP/oW7sm
feTBkG+YndvP/F5Llwg71vYWLHELiOAQfAxOspLHg3Jes7H+fQMvJtLFsWsk
50/BRYu/5dwt554sx06/UCQTfzPMxAgIndqSdpcHqc/zPQwfumP2eTxDc3V1
sek2bEvF0cL3cGxy5KklyOi3UDp9UrD5d/aYd2fuay3Go/KHT86nKtjcxyEL
cV3Q3acX3RrSGQhfx1jJaAI9dhgaYhogQuG/oJLrV754Ay9JvoGXzeG22rmo
S5/BKyZjiUPrFaKWYuiy/Qebhl16gYB3H/WfZD36vR8gBwgpiTXw6XIPz0Hf
xyeRgWT4tdBzAICbFtCqUiHBIRB/TgIKxD9cvR8ZIabzPyz+uAOmgladeiX3
U41bWu9vnUMlKDmaiRWa5tHtHph7Dv4TvCEGUdCXj4JRgKpmubtsqOEdYew6
WSjNzluBEfxgE9jeLhr9/h1S/gryAJjsvSaarG/qiC+XW2uEwrxnRPSs9hak
WzqANqdF5GH6sPFFUkpQAffuLN7ugb4zjHtXr3fgNWpRwYwcyouRG5ZrecPK
1VqH5kcdzrNqNUGTkRJYKG6BBfGjIZxD4MgtOB7jVXorFMI2GwRmdSXLORXT
DlUSBN4zJOOGKY6CnscY1ZdA6k77G1KPUTFEwK5kRKHdJOX0Q/rp1dHk+4jR
UZdc67WS49jZ3awEAkyLH95GrzIMxNp2RaJr9972dHOMPgPFbKs7/ki++BGj
YUEXrFCW1c1zmi6TkVVLQtxT/W0mOULVCmd0ADgDSDZisv3t7eGMqPr1e7VF
uE4mY/iZpsrdg0jic5RWEXsHR/p2bUQkbqEdhP2+c64FBAhVdnVwZavM/DT2
4n7+pi6mdIdb938fhnWDk4tMl2dx0rZDqtVQJmg6QUlq3y2/zXT2/iaKrGUA
6uPGHy8FMOikfddQzhBx/FfjfuTUF88hYPsLeWIAjZyRvwIoDxk38LEniXwE
/cZQdlGlGEaDf7UO3tYoRTAGnH+nVXf3ieGgN4y2UpZ7QAAXaCyLcSIqMrti
IQi0VD55jNSx7ULFFH/RE4OKaNx/BrjIqArjgNzhnjZS+wY3vgG+29DmnFHI
6JolmxuHLrdaD2cg2FO6w/3OhpZ1Q0DLJdh31zZjV+UK7JYHP6ilXEfm6Au3
vnWvaQdDmNkEu8El8PgIxEevtmkQ97BVJ5IcQRHqqeSOISkiLvwQv0nTW4Es
NJFfFtexZGlPxxT6ofMcgka+rvhsS2F/vnLKY/UoSBUYnmlgTsZz+40Kt6DE
gVNwDzBqtMm3Br/zvbd0v//vnEXSnD+e4F4ZQ/L88p8LE3u9JNeXANpd9HeX
C9nAcY/imgB5AT8tSof6EoYJ1dDua9seznqPtykFyObEULyqz+PBxTW4L7RY
CruzS39xJaByXOOwKR+5lOhAzh75uvGnW67D75QKrS/31vvvfWINHFCWbHx0
ZQfsxvLYp+HMR5z/I22Qyfn5GAvVW8r6kAJBhc0s128zgUiomhCKSQNDX9AU
GiNybb2upwo6n04JlqB+P4rHXMX0giGe+q+fnMVk+m+MD1x6VMFZJoaasCVg
nWW9HbOnSvesOu35fFtSMx/vSyDR/YX84cL4dukPGAJMUb00boMDPFIZKyKi
f+nymAenLZUKuMO+wv2Plq+Z5cNNt5zkNh289oiJONPt8nSxe9Ou0FpEt1cy
hXM9rC9fWafrTDoRuZtS0/B1SfM/Tqn+eayqzOo4i3FsZNh+FO1vRx/amz9o
0eTGKy2nFtbWMiAkeKyXdUzIRFHUyxejEdm/+XbxHq8nkaqu+eQhOke1kzZ5
SDf4PtpvrxXJ8Jr5cysY2IdFbgK57sV8i+SgakQoJT8nNlqwAhD4VdyGk95M
zSzQIYz4h0bVxYUwCd1L3t5EeJc3ARBZnWCjwP99BMiXgJfNvgIftjoRd+C0
ER4OrIcy5NZJgDaU3ffbrXvg6GZRqFLe9DCJRQmqfDasFey/FpLxarxE5VQ4
kmS7OqKpOCkbJ3MPL9CyJYlVeM4i0a34QTx2Bfq1argtNOSFQQun7excLlwF
zhzu7tE4e1SP3osKI53aHD5e8oemSV61Jsp47en4iCyr1aUECg3q2TLtbRRs
ry2pKO1Q/X78K8FIAM4fY/TL88d8o8JjcEihiq3sSYM2XFnFoVAf41V2TFdg
R7Z79KgRDGQtKKMZqS/AeMoDApemejflncHqqghY6w4Vja53g1hVF2abjJ1S
sAe7k8O/evD1eM7vsaMz3tvWCNcbgd5TYfmPKie7L3w1vJ/uxOEaYrpU1Ipt
kXmMkBnDE1rty82FOIOBCL6HYxtX4a5dIAp9rDJVYSVSDl2jFYfQ/Yh0QjaP
lEtxfZgPkEpviAc//q6qPhFx6yASVh6174oLfZc0mC44IAYnTfsp6HlI1A7w
eFZQ1YXyEzsEiu4BN96NmHmTmwM+/HyRaFQZbamitwcRJ58YS0+vLs+RzvaV
u84yRQTeeL/inOFQNXDorUtuRSMs4k84UUTOBJwO1FJ+4gXi+IDuEHLI3dG9
RHMF0LUa3f/pPAOgeKVE/qVsaGkrC4icC7zRFUN5nHDy0Bn6UUmCNpcVn5Ol
45HA+XrIHn67aL3DiQGHbp8wCjAvxKQeq9PmPZy4WsJpynt/y+Tyw5Cy7RJM
N9BAI3PHf3JHBdkUtklhlu26PVPEkNyS0e+464fEQ/BGNu5mzQCOs0xmDu5z
XQI+HGU9CEWF9CfSxD4etwJf/UD0EB2plTXsHi+wuA+9DpOB9x8ZsmfZcWO0
HosAvA1FSDQYN+Jjt1eXu0lJkG+pgTNm5/XPvZz26VyONw9VhrfyyRUMnXqg
TXBYm29TF/3Tszm4HQBi4DSGToJTD4u2VLYx4ROK9Uf6bw0W7LCAjZda+Acs
4YELzKHFomQSMq2NdHDwRAGrZA2NzAnCyAkhwVcQYT5CpjqTB++aQktatlXr
h6339KrSmBAZEh+dXKWXslpICMDqa9JIjHO6RJpmuomYh/+l7N7tE2VJHytz
VzIef7hL2cIOrZVaQqmh79V5AMpi6POGU1NYriHGtE1JI1D+2isZj6dkMf0d
3uEAswLtUdiw0n6lPsF5JzZghrh7B/hUef1Pihkiw9EqE+n4ZF2vY5cmEpU9
Fafv2D2UNzBJ+uu/WX7fiZQ1qINn1iKw+42WpypxbHnIIct/o+OW/risff7G
zxhrKrjWmoUJui+hZlhvClfaLtSuals7dnD22COuMhr2q5AJ3YPgXIKnbeNf
OJK2xm7NXptE2RpCThl7WLhd9+u8tY5aHBa1YvV0NmiJhA+EoaqsLdmMbypy
1ikAYPM+pjV8cgvOPwFJl9mJWjsCc5UAJEM7b8rMIYvjuraoJOxkmgZwR4qX
V1v5jU+C+mEWjidt9pfupRMJlgAPhzpCGaZD6HSPyZhnFZl/8l4dusXW5UMY
+Jv9CQmDRYQEZQk4jT66mO2riEdizSEcmOaHMzlSUl6iN3erTN4JSU1j0g5p
LxBj9RkL2yXwbXwkzrE+c7FHK18YmM/XiorbAOLquwwxcaYUprYMW326FZTK
3GuC+ldvBcUCaza1fjxtoNgKwBl7ZmhSrmZFTpV88HYaMA4FVfhtMq5S7Nl+
NzT2PGCyKAmLG5rr544SPdtUZ8npmrlkKw94mz/VGadRNnARXCD2kslVXQUG
f2byfGbe/UeRdHr4L+gmOm6o+mPAcj7XDBtcABig4R9QBUOEDeoW1cJX4RfO
TqH37JifkRveu3FZL7hIM9cNPmIOjTFnOM0yVx11+DwRurweCq4UrVxo8nHK
yHFlIYuxWRNAFwMQx4h0feiIfQNaAv5mL8kagAzBRtLk3wFusnpJS6mv0z85
DmJS/uRUl0+IxRhWOYbQW8SirH37vwfg0XSgAxzx89pAdE7WlxVeU4R7Mr7M
BXEuIjGk4VgfvRcNigIgD3efs2GuOMfXwdX1Y6NnpN+jXrMAsS1sXwgiud1Q
NqIdN4JyxXX3cU1+TcMh6ZQi729pWaJDJjl67JBDbfm6dHHL93Q7OuwiSdru
lF9xXYGBULOMIHL4mRtLrehb19SnphjjhtjztjTWEdnNqXHDL5vaQo0GKSYc
QQFpQpFN9zt/LuEq3ec4fA3bmYbtib0/GlOh7KYPFHesUWoxr4H48mPxMnwg
9YdAtgUH4r64KW4yPal6HzdC59VEBgew6/OW4hExnVzW4oPXVNty+auNC5Ai
dckT6JCt+f7bYpNV2Oia2KQocX23osF0b2JI6Gn6bYbHoDC/HFehF4YlWBKL
+KkuCGJzhTGfuIZzvUNGdFY8V07tI0pxly1kjp/u4t7NRWbS1nTp5f3ow9ti
LNYvsKAPlycqmEVBLBwO83cUD6L3wWpHrwvSP4vbf5UzK370Jyd9zdry9d54
gCqj1wpxSlVX+m7qHCK2rHMoDOUlShDwqXBodFJTwkFhGwVh1UZoeCFXDnQQ
dNicP04PUVK4gr23QSt6z56hIfD8lnQEYaNTS/huqYbOhZAFYaWy2hUPWxoH
IIG3ZRpxkqlf+ipeBfpvJkVjDNvdL8KNwWzVz3MfdWHBvxounKC+sS8kyhB3
ubIBNruOTDPGZwa4zkF9z6ry+Msiv0WaTXV3cRNCwokNL882DwQoIg9LVNvW
dJNoLgd8cXfRKbAD2ANJAYpAEJvfJ4sePgf+QTnlPvULF3E9IWOaA0IOGliv
Nq2KKarMkE9obLXbWzgpzAsa7ac0o/0raj86Jum92aANMCxsLt87hryweFNb
IvHEn8vJnNpEcfH+xcCBkJ89+DYLh05c7ARd+FEdq6KSWpvAAQmKoSXiIeYX
4hafXpfuOosmOzP0HXEMUNGZe+MINmV9fdxl0Fe1dtks3GMaYu4QbSxme4Gt
OLGQ6xNvkkhIQwHVK33tWOi9wGumiHTpYtwBZusA1l7DHGGADWChe4gY09BK
09BopFJVaM9DzRxB2YtREXyBwtM4OHky0JTi0BvbqAu4LBGYae+rKOED+jy4
JPufk6xedamVunpFZASCD0FpiB5y6NBjoq9uuMSdYLlfx6T3oiQysfInuMsk
Raa0Ok/kwByZeriyTQcerbj5tPYY3p47E2sJ5GKsJMDfc8EY6Up8gAMUdh68
JilJSOzzCCTmk2/ZkuRHcgs4xH++HRxYSfAvKJNIRhT1NXkh9NY6oAiW5+DA
BCy95xjMqp8nxmzjw1Vltz9MwZYeoxEWQ2KCJ87/XBdHkcYCnzACyftxCJop
xwiQ07upYb8dBgtQDU9TnD7N0WsXanYkYghwbl/NjaWn4/oHlHatJrNkw/B8
UzSngg/WlvZ5ae1DIYyJ3P+rtKzR+qeJHdAr8YHtBeokE+wMi+qdKdAU4WSi
R8PAgJCFRc4A4eZXPaANNgXmVLNFTAeCjGeXSX8F1n+NQeFNencFFsQxIdZB
Kgg9ZzDtJlGTX+5JN5WNhkcSIY0LVxu5ETnQntpZ5uU4MmMrdwmkUyGtGjGT
67OZzsCH6mCQtoXiUb6XzNtn78CePQsUGi+Yl7AicGYymcg3tLCAoc0ePPJ4
dvtSw3Yrr6t4R6NfWAJR+9culKiSx2jHUH/Gu6Zm5t67MSMHURMkOEvhkdpB
gnJCFouRjzKek46GKf6lYeGxg08StB4XckzA1rF1Kt7P8ELHGSLLj4mvhyWG
Jz+Av2N0OXUDBL+oQi3LWvAd5Z+py+qDj/lOLhIXFZjaJin4wsoOIkB/9UNj
adrHjzCMdzJtrlFjVEbbOE444HSh/ya3TC8LgH/LXchi7m5Cz3avDM3AWTJq
VvvljUQN73xXHTTJcvZXCuHwhh+YglhOZtnMrlnkVRdMkkWaNE96TAymWVSa
2it2uVog0GLBIknPbILI5RkAYnBTSXgHR/i1n5LDV6HsEVeQXjAZv0CHnlgk
i5wnXPadooDmtbaAdI8xsGN9AqVg4v6sn2AXEcRjbtRNbqW220h+CmOJu91t
k/wjwFWH/ZJ5DeX3zlAR9Ai1v24/WvIc53w5icLT1fNyfikrlBQ2V5Cqj+T5
HQ6t2AfhHoLgTPw+2Gy/WB49I+72TySbZzCNCCQrttM6gFUbbEfq6QRz8VUo
i4tHb+IaLn6A1bScccpM7gdltN9aTbF7lsNl3tDNM61Row4dRGY9qr6VFYzK
tCDk0OJ+FUiM8IDzjIiGHo+2h95Zubyt/S7Or0BtvjDMKPF35Rluly8oRSo2
D5MXRTbHWusYi/XXcSsMPUGknj6URBFU9vYpBlF3jsNlNm86Z14jQTyv9bIs
kiqws/T0gJizChExC7UkZ78LdiPO1y0i1cAYlYtihR3Kv+gPAovAEixEgCPL
Z6EJa0iDa5MoeO46HIzy8rPfBntzTWyOe+Ti2hsHeNjtqadDS0yv3U6fZHnr
aonX7PCYsFcFBJznWULil0N2tqKW48TQM4f532IW25ZS3fAcZeP2WSH0rIey
tVhbeUx/zgwLlWD01R/UGjTCifhbfcfyiDvknAUDC9vRgkWHxOHb1qJCzhk7
q0rOTR9+u4SRNA0f/tPu0iThfjeoiqkn6D3bQFxVO3i8excUHzkjjB2l9A5i
hyyRHQMusrx08bM8gaiuDalTefHBEAZq7HK4yqq/FmbfJSoRqnQYXZRUIZ8n
z00DTRpJQMjgp4+0BTU9YvvJ+RHqO26CzCae9bd0il3jpqLB6A3cTDOdHs2G
ZuRGpgj3Ho3duUSi1mSWnoJNSbL6boC70CD9v0vnmL/feyht+U48jZr3u1wO
cJfTBM5eFxh3V2NqucdtqrZpafvT2HYwAFD/ynMJ8rYCGuoSQiZzj+NwNQCa
L7AiHYGCUf8uAfP+6GVy73RRcNki3ZyJi8/QqKxXhOO5nr3WMoMgfOs+e4nq
ZfHzQIq4e6U6avSupDAC3BvsYf3aUIQaBQzYiZObW6GiKFZB7N5bqyyd7jV1
mwGNeFx2oA6DzcFaIzVsf1EOrPpUXdXTtPL1hnxLwj2XEWDhW9QMNzF7w09m
O5Dfm/dEAbygyVzweEkMYh7M0g7XY0h1Tp2YoKEFVsrRisJmuj6hEw3tGnwp
Xaf3WP3Xk5U38vIuEu8MBtx3g5VwpwRh6Btk4cOCde8RrDWo1Ywo1JjeA19t
tvGwACfJx7ol+4uGwvlAiMZvbDW7skDvrLp8vqNw4AHZVc67eA2DSQ1TFmlK
rtv+0tyxqz/Wa372w3dg96ZlidnERLrSaTVEwBYAZINaRUmpoQ2pqmk96GNf
j6/zJIIsV31WgqLnjsSKGWU/UtAiDhKwPUWj43YclKnw3kj4/giWEDJnLH3j
3rVsUCkWLveqWeUTA8+wtJ2St30soDAu2ESTIUUzRvD+RHfbV/eM5MGu4eBL
nKJGlR6MWn5yll1SkhB5Vw6WRVuAh1OyekOEYT7rWpZ6s46hA+QKc4I8JJYO
7vUHiVPw0q8lAZhd17yPnLA3hU/xcRNlQ0C6vtdualV6uEH0vMjDbqbQ4ezG
z/4CWASpm1rJU3k8Xc4JP8xsRRO1p42gUe5o2gBibHYpekE1UvamKVhmjcDZ
Uuxg2/FJQGlH6sRkNY2MPhoFcXYalm7HBuAYNYjvz4FnHBU2kPsCNty8GVZO
hsDJAgEolJ2aSfpSxPsGFqgdZuuN5h5KCvaEwi+89G/qC99djSqM6/QY+UPL
+/BEAFX+quQ2xjAK0NXtcVWPicd9Gb5hPMwXS83pnqphSOdKQdF78qJtj++8
GJCXoSu8Q60iHsKdIKJHvCIAB7gkPFYSanYI7qcCuvByzJRFuMTk0xJ7pE6o
bd38trMqgCVIgV6CnHXbSSGIQfYO/9miBowwt3j9yijhBYuiJBkd1NR0tSy+
VKcHm7oXu1LRlasHUBgL0TXZQyKdgfEf2LPEB1O+YSvQIfHzvNfPGzoW4juw
+mB4tm23oiG6aySJIW2sg+KRlqa/q5OwIHFRzXRRLtKv2DiS5cHlMI/UFGIK
EJHSA51S5iSIQku5wI/+0nMgy6gy8/80rm/O39K/OMMQWvggVvRVPJJj7tOi
/VuEaFHdhDLtJK4XH6Sm3/M5OKAMlW3XHbvOxOdwmK9+sYnfMgaKEoI1owsq
P2p1/7WEjOWk9KXlf2XENhxWAM3C9JlcUGprmJrcJ0Dsaaa0UkPohV2HSYnP
9zTX4deENC3Ft3RZc8aT1a0PxIyqSQ4kdwccqIuJTwS76Wm9XfU7oNTAYKUB
MYJkHKlMA6Wi8d2Uk1myBJxAFqkYPcfRNKcrnb3pNIxcS0bBw//bMGT/NK5V
vb1E+Dvhyt9QJ0K5WzmAgx8B04cofdR6TwJkrL5tt5DgMrih5Vfiriof8PHk
HWHRnU3LoupDMu+ClH8hL+R1I4NEXVIGlN1wUlYkV0KcZ8PwCVsUdlt+gX6r
xAwj35HlKy6mKDEZA7p5ShpEQEORecJtWLpq5LoranX+1G5KebANzw4ksReU
Vag6uLL0mJLu+VsYLrA5Jo05RjzRwJF4Tbc/TTdftb7h4BjdzXTagnVjsVPT
+A4Uju7Da2+koC7CxA48TpD9RT7dfy4yzwAX8P1o5RBw4TVhylAPvrOPEVg9
fMFLDPVHVPWrAr7jBDugvNKlstOZsHfvjG7fQuvnA/MtpNJxpjhHm7ovDkCo
Vhn6nuY/QyshHlJ/rTDh02lIJ2HQzzijoLBf2Nxw0j2k5drSfHgxz1rn+IWH
PDFPkDKU1vfzOSLw+tH0eV/eb244QEc08QzpcZOdLwdBQHlb2WnVP6GczKlU
KMX58WnJW2W35yQ4bg9qI7Z4y6R57H9PZdm7My+kOYaFQ3+DUG1e5DFDvyLY
QrYIVXGGXV8uW2ugZOTafDT+Pj1iKrMADGPKHk0gBPJGLEDCi9GvrPbbpbFe
OKhB/vApaAyKeNa0/EPv9INUN8uprWtK3ZphMayiE0sJfWQ/bdwD3DPX/ZSs
4mpyIzEjeaOECeLqYr/LKpczvlwUkLeQhUoXuZWouRJQSXGhex5COe2c55G0
Zs4pj2r2semZaw8zsCCcGPgmrvcHfquSNEJAEvsAHX/4Eqkzr4bsQpb4YdAH
lo6p1t9kO5J1rKDQETFSF7KQZPNA0aY9W1I9CkGhcJDCgoX7uQtEAlUBfzxz
L3hKqMp3Px2za2U9cvKfOlXhC84lKnKHTabVcVIev8Yl0vMyb7F8xfEWNZKj
2REEuKxRuLhpQoSBg76sF+0GYaGeB0aHEJJpAz2QofeG/tmpRLak9cCw9j0E
abhoHq6n3di2sliHz385wSNy9NFiJ48xxaqbaK4h+5/k0aym1tcfjazWZ98z
SBiRWfG+p3bP1zXKjsqju4whFwtap6f+cJAT38n0E8pQB0/ICqqWkj8S0s5x
Sti19gO9kKQIbS/AX/eF6xehHxOpmUD0QtPwkD5YvIcnObVV8CCdDHqYuyYM
7Ghg1nM4+s2TeGlQcSwjyaJkBV+Gnmo0M6pW5aq+dtEnYTia3JzzvSOW74AC
vR2o0Hc/BqJzFo+QIaOC71dHqAuyLOKT98AKJFfDDh/VbO4BksbPosxJTclD
rkfCIM2o1DzrJqgOPo+nqkAIx+278ylWBvU6ZNyU4bBEi5nG2QW6xT8zB48v
BfTGdr2D7+DqVOi9Ci8BMXs4Y16pE0lnrPFfHY2roVDZP5Nyvo/1jjntQedh
NtvkaDGJy1+bEmpTwlR1BgmwPzMTW7eHkhe5Zxl5FCXje81fqkCFn/1HWCjr
u03p6RNh1yUF6nIjH/w/z/C2qp2iB1WPATVki5WSImR2xqxlbdwOMnw6TQFR
yuYiLI5uf8B5RnaO9wSxzjgzgDiGSM4hZVRfWmVfuD8qKPc0LvyJx+XJwvzI
bETDGsyVVJjUqso1+xwiLP4DPGR0UM1E2BEnlYK2HyzMagzpIPM8yb7Ph8MV
dCCouS9HQuKpf5EjjSHyD7sngtPiYNcME8BgNmjgcarqpsVGRASy4aImHUIw
GaczRSGCP5Vvsq05ZLAfR6x8Zu+QB57dFN0UIRSrHDyKCJjR5PY5Gd6djzon
+BLPYtRtA2I7N/EGEnmAMLwhilj1i0DVxfcrZ7Z1rPKOBZOD6kPA367qiW/z
S30KpInOttGJMhF+fjLQUggZ4tqRtlIsIzGBw0ecJtvwYmMxtwSaYQ/IOpSY
lP3XmpGiN6R3UhOjWZ6YntSw2hubNjS5ijvrzWgSSt5SK0iVLuS+/5c0iDCJ
Y7xK6/ISjyJKHEE833pFtEkhbK1npBGx0/yOrIgSz1TkUim4unpSO4jbIrop
ZzdcXx+bgr8r9ss/rG6Ro9tboLlzfkQ00DFGISurziNKj6EN+Pts3BNfuE9/
/NmPiPivA6ao8I3QGRX6BYk/g+wQ+4Z165WEFMXChFS5uIeiwDvutNdL0Qii
rJ8qurWFIdYGvIvWqRHcTsxilzelH3ZhMNjWWIMQDB4h/l3sNAAqFmBPShCV
6aglnTvCxGBxv3wJJeiD6tf5ktNUpJrW9DP10yt4wrZX5nc1ofYdA7k2+HQV
yaLflVPi1+vBlTFvmbge6DTqRC6zpumKnmnX6Zv7G5VUVyNhwH9399TjeUH5
2nnD/IARhY9n06bTliwtzADkaj1JmEP3bHd3p1BM/CIGi8xpsKMm35TwcWQE
/0nr8a6hDcH03CmhWpgIyvCl8WITumapEk5TrqZgRhB0qD3WO6Ptb586h83a
UAeaBPbqE+rNh7lQv53JXfVkj+DYES1cTrOJjg+Y2rVqiNB6BJLSRD3v2K8E
vcmAj/DhoC9/jUu2Q4FKW2Urrkp4J5YLzjQ7RNqkoQA4Wino4X8Yb4HYFrKO
kUNH+tC6SmQaXuQbtr/iKTJaGTfQUpSX+y33Yu7Fqf0nebbbvVeAU7IxEJFl
xcqF/svN5WZJg+uja3ThXaLUZbdBlMn3bWd/sL4J1kD64eMVaMhKQkLYbG1z
zdE194Lc0Y4DJOQOKYGVMeugu+JTM7ZGVl3cFrF1kALrax2+sJh4M9yHlhh6
uoUB1CnysFY4H/MD2QW0Lgomt3yV0F7rxFN75cYUpO5NARN0M5lQZJ7gy92v
SuF7UVvVgTIfvKPjLXoKaP31OmYsvcA/gsDV59pMVQnPoqzOjByOyYuatIDo
MthcngOOecYw8CFFn/kX+S6RtPYUiPunv3wljAN6JH/cxjIv6c+qI39BmqSF
49h2HzhHsVGarieal8a4hkNGezNpHxdUvF8PwSl+F/yYdy7xU/WDxpAWrkbs
a5+0Zj3Q1s8ij/OJgcRwSR+m0PkOOk+cGTpX3do9diRfFnCXZ+OCPLvo8CyK
g/LMfkQnnZl0cNMp53OmRVxnR3fcMmJGg4bKgG8YMtgaxy1gK5J5Y12fnNVR
eWXHQWJT4gXKBvwUyi8BDQ4Q6I1JeXaUEAUDDTrZYWz0No0gnegmDOv3fk34
I4Wmz5B86+OONpy9ENvHbw9MseR77ha3pjhGcuaXbu8frqUveMLsUTvyKUoE
y1Qy/qiShCF9jDB3hmD/U+pV9wvYluAOudG0ldNJ1SgtC3LYlDmMKhtHeVOz
P8lP1uvWN8CgA2/92s4scuXIOxL5roCFF1VTQHTNN2BK7BBnITOD24gVO+/k
l+JUGxd603SjTOk6QeXp8qmxAAO7SykJhoLvpOVdRd0LMwGOy/jYQmuNE/CE
i03wg8A4BwQSk3aW2YfOutRqh2STt/mMqvv42XVz4Xoh/X2PK+Z6LLDrIYlx
BkIYPNZAkZdw5LQhH61WFMeOzsIiYRLDtXggMcC3kXnBMTnwolufyaVKf0OQ
GeuZbrqn4LC4iw+BKBgVL/hSGLcVzAc+9T/cBaoFUKyOiTpe5KEdxsvrQUSm
YNgkN0B/4RtxxKDV5AkNw5wAxFG1HqruyT9sf9DrHMYAKUilpxjv5bgeSP7T
bzIbhis6AHfFW3UKVq/mlkE+qEwlG7IV7oO7VR7A84CgycjNW91uUq+5xXXJ
Nn6rdBYqMjxvryomUPkLT3u47GBheTARWKQVVJiFo6cyZqoGcmW2JOmqHItS
ABKQeWWyGGXOrAz2+pGVqmhlLTMwE7OQsFiov6CuGpHENvPTvghwSj8L8ojN
5KnXNaugFzye55QVnkvFBG8TUv/uST0GMu6CyX9TkSkdcIByLMhIk8+HoLJq
2f6JUqY1oxukOiuvAYFT+SYRD97g8ukriqacnvkcDtfFQWi4urT9NrNIJANJ
29y7JyZI7zqkPvY7XRglITha1NuvPzfE3r4ZoiWA2GmdvEIbmyJJc74d5cQW
fEtMrvc5VBkUZ+waR075bGdVyIzodDfTkeMJxmdOv63eVpz50NyCXBdct7QE
OvSUYCOJ5ZMATWnowZZduy1N5AMCk5ewIwPgT4Kg5FsaqYXtq43yI0GCIqk7
YOwTXkULTvlFrg4tGjyWMl3+ZUVj7l7x2kTzLFWupXspTSUPL4mMDXdamfGb
XMmxNZWTWiDyPpkU2Ajgyxktr0HMCiDIaPdgksb0CaNTb86zeD0V2pefqeoW
TROcB7PnyH/QiKCPmqcTVwolDXOLdLEOt8ufR2tlJ7KxVa8Yq/Kz9HRqBbwX
CQ1if7JbPOFZdwm98SqWgdRPGlfKFf77zFSMWEPRipGWO5lLpztj91jMDm49
Iw5Tf4P8JI0ZeeZlCLHuRFGuV8XQIumpNju0iZ/LsWR87mEtayoEjRO1q/DS
/byNHBv/Vuzt6MkgpqFWZp+hInpDyVvIATCT+8qNsW1fUQV7+2qTMU6Nyb/8
3uRiCFngAAqX/a2m68q1ij7HkA6e0Q0zklhR7C/QmFB2yu2QxjTvOjtncQI6
h1m+EQzmHOKpVLdid0OTekvWmPnQTaVPb4ramA3NonKkn5yE50qvsabqM4T7
azlQZqnmPfb2LfpgZlCIC0IybqFfm0y6K7dBNc11K9e9hXKceBk4qG3peBdT
phIOVRgWa0dUOORj0boWj2L3vOLEG5PKzw6KnVKssfUeE2qIVyqadQQ/Bj3i
QZqS42GlExx65d2hQm8asreSEFExfv13k0U5/xDBQgovaV5akfs2qkr9WeZx
Wab1H1X/tjoVUz3myZDjbQasgC+SiOCgyXezJa4FV5sMFZCmces0hpO7FIm3
MBNvJZUHGhIIiH6xMKHb+x2h+6g2t/a5I+C7RuCj5yM4X0gbqnd4uYN2k7pj
riLp077GXBFq58LseXVQzLWYMrUahljR9w5HDVC0FWUFZiHDIjc+UeTJurUC
E9xpzy1SWReFH4znK3eFSkLCgAS0vJVBKnSGIMDGiah0datBWLCO0I0Kb1tu
YTCtGbE7rGVBYcCCSU76+mR9opdfY8DnWmFOXmO02OLUARN0koyCgdeQ45PX
86ROqcnKV4WO5oejVZpXGZxAlZMbCk4iPToowbDeZV1i/5kKydwvY7zN+vId
ugzBSterybyuUEnLUlhQO4QYv9S/3gcUanqiwCDGd2uMJ7ubx7TuCBzNbm/u
O13M2ELxTLgBImehlpzuq3kAzm5B2uokLXthL6eVgGl2JP9TB2z5j/+CG8Cm
qMDXEiZwk2I7KuT0wJ2gYQyfZ2hYRSpSvIenlF5OS7X1QE4zThDDEMfnUZSD
cLNJZQ6sNSS9sP+1LRYS75ZL7ErAKYV/koj4pEvvl7/FBoDYWbE5T2UfsGCC
EUw5YwgH3nabTanW5qTfEcs+LXPkWvboK1qYX7bPKaM7FKc/vOn/Ta7wE1Me
x1rjSbSiWO2qSp7k8UKzgRDwuNLtv+WiTZl7yIhbtRwllW4583n2tayyRGXU
cH2v69DjiVy53gszUJ3rxUHXdmMfxNQUD3urEmtLqRJGY0GsiCPY9YyIzPl1
i1sa52/8vV1NS6RfFFpS2tYmGD1DEAdtxm6cvmkF/qtmG2BZdjzlyybXwcJe
ZVpN9e/Mpa5/g8zIBNJpHffELBlYnj34YnjnHEFUUuyLM8z/MjVt92TlS7Pf
qm+FbApqaYxRIm7kp4Muru7WZAfYmQ3ApT3/KK5dufsd60EHhDqhnwTXY8aR
6TeZ9rHPm9Dv0uyupIhDls7BjSmvMOX1nhk8QIBq8XsqP+Hayu993hdsdppT
SfO2nedyhVCA+4IgEQc5R71UuFet9LJPfmM/4hQbO1FlNqRpr3gdsEZExvkO
KPcb8RciM8ObpYRO6Rhgo8MFeWcdJXfndx/cSKv3bO+Pi3yk3WfZb1bfGsjy
LA3605BTkpo/RIChZP9wa3nKl1YXSCYF3CzVXQGFgN60OZR48gVAx8R0zgOI
aNZz+gLDbNwUTA0CfWX3/nemUV6LwFbK0JGbEgBB+wvAxADhxsGOG1qpkDHB
0q944NyHxHaSZc5xa4nC5H26cTqxL1egi/AdFlYHobLcpQrMzvDYEECxC0nJ
n96u+sbBu3tS6kOBcD+vI7/sYJhTLzbSFhJQKrWmIR9OgvQjUS4lgwRQ7K1x
+EfVbM8DeaX7rwAzgL01luakZ/wrCw+2KnIuUkj1/LukZAxpsBS7bi7FJkfb
DepzgFdSvN+ojm57E8JVnBscKaEebE2MN2yNhZJopfZ9PbuSrlGv15pRVTQG
X+WSNF0IHoMaEiVi74DVgv4YFAaSNVrbm0GzepU0ltabXHS980e0tm1ylm6j
S6hE0yq5wSK6t/rdM10a5us0muYcN2MpXDrcVqQpJR5cXhLCb6qnCitDr74K
odA/EV3NW3fLm9ulbprA6N0gLHsUnRW75iHZzb9OtIxDAk2/9ucDD+7BPp0W
OGP3vbDO27+8H4Bixq+ORotniPWYFju6TPBXy9DsWxCkf40+QasGtz8n58wS
jmOIe9MfI4h+G7yDloGfGuTwxYp52KDB8UxCie8IMK/xlg7PsMBX3FhOptGU
//pRaTQzpa0igKBnA1MAKkDwUfXoKuZOdU1Lcjbv1vZkosE7brqoAdsNZWpX
Wy+LXHiObbAoyH4qf2TkD6J0n9IrxCEYJIUXLhQt7WzcuB/Pf6MpvBL+BSY+
Q65Kg7fBvlCdn0jkQfRDOxkx8yE31JpHCJsKSrzkiJXb7sIeKh8kQal7DZOx
9Xa4haIbawhMU3tEUVPk7h0CUA+6BdSxmgiRxpEWv2GyFBcKp46VIVwIye8o
HI+WeaZZAZx126VzPkEWgJMaHO5bdDkI3uxccKzjHf3ozisp3hXiAbUpwrcC
GW9dalyX/O6QV0DF5u0M9F6NdTVKw8s5MOfo3o91lGCddFc2YKBPb8KM4hfQ
2CMiLcQ0ZQih4WHfceDZPzZP7IIpg/5DWMA3/EM874VEauaD4fufdTibtn7C
D9lP1/H85e3zX3O+75xGqPIeC4iGurpELdHsw2rjUm2jXAJKeuXJAE6U+k7b
Wu75/BULKSSlGYvmI1xpQyuT/ms0boJyLHNnLPQsnVIPujq6OcKepTcknu/r
4NmyWLNJTB0+KZu5rXjZsbyou73UFdVnpx+XoTbEMeCUfOtKk43+RH+Qj8c/
UxflFKq+wNJ1H2aFUf9S9NPtnQE67tPZwt9IeyOxrHcFZsKKeAeLWtoyrHln
Jox22w01w8tLy/4uLhCzqWaxG7NjTd38ZuP2NBr6loesZCaQpv9TEQg3lSf4
sTT5Og2M095n4n1kvDKGaRnO7dN/EjJ9R6DaWjnkxg0CJ0cKGypkHnJsMcUw
zQSTS6mQvp4t8CL+lAyKy910w4lD60BwPv8RU8mMfUq+3mF3iTKdKHwUXuHp
ZKmRBJzYq+JjudjWP09fLc+38r6zGmo1ebdX0Cz/ZvieamLstVQyzVNZ5ZA0
BUgo8zFAZz3qMF8Ex6aW0+hQaO6dBVSGz6x/dAuaEQ81VqXo6nSYs2m2pCW5
zlOd17VPsTAZWVJj7rxYbY8JreihyFhaoHGc2wTNlT1m54QCgcSnPdV0VYJ8
ctxuAt4mHxM/yrzBUkOrH+vgXQHWJlQqSMjU7tmdAedRMpRbAP7AoXzfbtOo
VLTYdby31m2GbtXMbqRhlU91C++6ORZsAdWUAVeYSdba2OKWGvcBuGGUoASM
O+w9NvK/oed0SryuCmMHkDj4K7Kc5D6gpM8SdVobno2gIUpGnKu9HNXUqoEY
7IgznQVSKzHO1Efp8bSWarB5o0n/Y7Hw5ZhddK52DHjB7K0N4aXp1PDcIPT3
LcLuAbw6zygrkbqxyZKnufJdSfsION7xjwsesaHO/nXJxNOOgpYuSLDdh9z+
7geEyo+EDU9isPdcwYwvZuY2lPNkkypeyZc/S7nzYS9VGdJPtlYWdZBf9Pff
1h+wSIM3SaGhcuYixm7pfM3iGx2jCBVxViwIsLwKXC58XqR4PXpRo44gobj8
5FiF6P9cxiyDbp/2T4mktMmX7DdAaqbzAzWOypQL6WhAA78D/pTQ/RWmaCxd
4r7d5fYF7nwdxcPYUeafgcLdTil3r1ay0I73H/qu+b+E9rQhNKFDz821dHpg
BRoWVldINbafM0esesvfeeSL63x7ZYfql9L7MItX2aH/om+0Wv264YvOf0Bf
hW10G9YAQ9uxnOdcucdzMvdTUUqo7AWSBuHDeJJn5XIuKGuM+b5ZTDIW7Jh1
9ln3e842ZCddx7/ne+0AYTuCTLiS54n7gyVGa8JtM0GTdtmvjWH2miHB+D1C
5/V/2Dfp4DyWc9tFx1rzzL9n0cgLZsBitubeXDb2/NS2RbnrwuphBl03RsTb
pQpeaUEIJW3vSNW1cll7LXhz7vGvHdHdp5K/ljTUqwxroHlyzC3nlTmQRNpb
thsXV37Ov8uP/AoVXlcvTSGMTPjuOm2isG5PMd7tqSOK9iRQz0HVrfUFstB+
IGmTu72HmBAcym3ntAm9167KAy8ElwoOXTUevZ6i7IbGr+iu3mUx6JNDzROC
16Z8jcFGcnZUCcgRfMlnZeEIQURuY6RR7Ugax6PvknDzF0RK+B7PuhzkoMbI
GQLb1pXE0rYUPp7C0igDeprh6dxl1fn9ZYt2Fp11Gif4GNd5Dz29B5xNq+7o
yHTrZMUpDxrxMJLGDVxpArn5pe6M+qIxxMpQ59f5ar2aVO3hdyiSwB6YEwSS
gn80lJHd6gcWQ/68PcYz+h6Uz64YOWO/+5ixfUkGnQTXTYvtUN+Q6CXrtmlJ
F+U6myRERY5pKCbtoAD0n2MCcyuXph8+RMrzXvvwBM/KdkRZbD45gMfN8Pv9
Gf9EmM8gGxyla5C0qJoHQQuzs+SOqdcekKASxMwFpor5oiE2hu+FtvAZi88b
yI9dDgtJnJtHUOschKGh1LL52tDQAw8N1oFxKgfY8pKNC6BJ2Z4hePme/qY2
MR0r80i7HOjwqfcKvwdV7b9jU8qZo97IfpVh+47PTmn3trqNch3Wweb7mUlc
pe4oHvlBwTvUMTH1VppXZP15CN/uYrJ+aSuwQ/9/m/xfbBahzlymLXeM2W6I
LQ3uTu+0rh8usn+9ljOQoJ1zbLaVHkVSDj70kB8uCgOT/XDuZycTcYqIlGZm
DkCbRCIJk/N5RnRXj2XKlVee/26czfxxrLzyQqTo+r4E3d5pErBCi84m8yPp
dxWGZfiK7MDTK1WTAZVLbjndFSynOYjVRJK7QORvbfVdnvG5yd0mSzVNZoGU
Lm3yqrOrJYi2FP4Tkkyc5dSoZM+eViDt8hBfV9uez53wDr+BIG11FS/hKTeT
w/UP5IjWJc9jm7ifFiy9n8upFjPBivDerRQDaCq4dG2MPiojLSZ/KGTGsYhL
spldmbRu9yaiygMfBDkULu7ULlfCx8L5+ueFAzuxYrFyZwB1paTrdDK31nRG
Emqp5Axn8KzaP7R6sKBoePaJewP3x0C9uGAZrqlbXxoxdmeEYCwXLlvJUd+c
NOSxd0gVrhkejt5s52JKdn0pSYGlzxlWihuMnpW2wRHqCwwQDV1144znFNVk
t3RUbg7d5icC9/8Mm78A9zwc/2hQgmKfv5u/hoGnx+8Pu/VstuXzEhXYEV1y
KTYrAmR981Y+uVxF5PnZJuIzatwInSu5ZuRkNCCgJeS15Eg+tNqlK2Vc+goP
KYlL7XipYZ0oiBR+CMbx4HPSef4i0qPyLYaDXY1voAHeR9pVnSy5qVfrJChm
OCPmas8gu13DAFQAJQQhVqHG8iWizaumqxCVoeH2ltFP3mn1hTG3g4/tgUfT
bADiv3y+dKF0bRbJYv6juvNTUVs4MidtJEcoeZubYXYIT2ReQU160l8QF9HD
oJSkehj7PpdKTPkZgv3T42J3Z23nVZO7uSJuhh7KvokcUPid+FdM9La6WBi5
mDqNELZxJsllZs8Pk8uPshX6176TAxYOG+FXFbuuHHdEBS5ce3bg5J8ccXeH
zmGlSdaFUkLxcL9msw/Y5iI5iiCBUMvdCv04Atim6iigZuXYIhtNBDnovUBL
i32VlCHpLDaV1SqCSXrkcEWJPgbrxZlb83KL3U3w1Ivlyh1O8caPIM0HFSMz
PmBRLrt7q610sTzduo/AoOYGBgDI020mcuCoW5cnuDceLoxTM28gX5N6yFKI
+ueqRtvadmmx6NNaW84mVFzjEFfEddOWFmfpYp0rx3mLHTZB907P7ohP8Fgm
vN3QBU+0it8gVGZ8THslQNq7VyJS3EU0J/kJVu011nV5m9PY/Oo0RFhK6PVl
v0kDRcGuPj5S2NgvnmjGD/ilLN8P4Rh5SrlVbg3/cdFlUw/glDqfdvO+3344
ZNoQD3S3M/vQFmae6Jxd7OyMsF6bdUiSynlMcZpKR77xwqtxvIulQwmc1GN5
Bq8xLac9neB8pYC/cx7uSHA0qt8gxy9AS3J3QI4jwUJBnrTD0Ous/woDidv1
IIGuYM4Q110Ws5XU9g02bL9H2eQ2LiOLq91b9ZOfqpNnxcznL5Sgxb7vbVAR
nIAqIcm0d+Ih+skkYCZ8cJtqUIZ1CxvRqLk7szn5WlxDclWxp0pGr5Pjid63
wI5x92WKDtx4l6yCUn5REeUCh8geYCDHWLWavbwezV4ZkBUIEOwPc+ZP2EQl
BxTFDUe8JhVDuUjU0SnFamu+/GyaN1yDM4ReuPugVhDxsjOZTVNWmpdmx/Ve
uLupo5Ew53/0L/PR0nm35rm4anHaOzIoyWj/OFkqJf0BIwkRkwxBoVtaZ5kv
8IhejeEXh+Yq8RunHryEzb+Hg8whOIInLJ97RL1C1lpjj6aX//9quzTDvWEC
yWBL31GqeTz6bPpKGaJODoqnuYp+GpMmfzdyLyA/H1x/gMyMzvhdzt6AEa6w
CKlXwdu8FsREtBbxy1Qg3OzqliU3QqTvk6DRL6EUHZeBNTrXTXD93iyv4OBN
Kfq7qFFV9lFLUz32s6wj2/1uB1GcpINVCNrR6nowLkl1XXHFGqlVzZ+0fRSP
9ICVh3LTrRBYJihfOIjftvB/DWqnrv47mYkXkx/xbz5fiJlsA/xGAFJJ+lG/
vuheKs3FkLnvKgIZgYaxn0/jxiqR+a5lTDTz9u9oF+iS5jYF5EaEastRGdkw
UzkZKQzicyDHKY/fKu62vL9U4lSnj/UR74Q9P7njn/A/qweqkXap1l2jzqzi
4IYx9/+UVpxM1H5USJ5IN3rMwT3GNutIwCVNZLfT638CyKcs4eISS/ehcO1L
04wjzqwlgXBJEtBJ0nMmFs7ySRh5gHvUrr9zzgWfW8ctViJNnA2jKW8bAxO9
nY2gcyP3/3kIvuKuMJqBufRgGT/E0tfR6vGNS7Vc9wGNqy+/xn3vZzu/mv6C
82AmzEESo2+XsUUVUxgAM2kOOAdb7GZEnANUWG4SVcp1bsEn233wIULNJoWN
l1+vVSyzp3O0e1GJHy9U9MifUBQajapWC4jAGLBU2kAPJUG2qZOzSBXTzcsL
KWP/lPob5X9YOK9wJbe0nPgQ/cSZsZiaOoZ+lhs4SDyuULT/49su7JnezklA
N/swRRYNK9weOMnqE2oEgQxIldXjulEtr/jSnYyGIgRlo61ockZQi4DiDKIF
KjEjRAU+1UZBgjk+VfSBoikf3jYNwuFVDNdcLWbsmjCamvPbGxcmNrXj6tr/
re6ILRpXlsQ4N7yV3o3tD7saja0rzfMBANYEqGOEvrOuH0vH3+YgHUxaOPC2
9uALbJp+CtXo/8G2FsHmx4OFuSWM/mR7jZmWpc2nmYQMe3jlViWi82Mdu859
RvaWocvvdbq+0QnsYL2ug7fvQi2QkX2kELBAcIfy3kxfySC64TZ32FZOOE5Q
gRojGFB1fMf60WwHMB8OmzAFOpKcTiTIyl/lMoFhd/8D0f0lj7UA+FhF2xED
3kkwLNiVNula/betpzzAP/lqfraC23h5eq0mt0aZF3jHfQIJTcd2bUejjk/j
UtVr2eL5RII6NuZbntSMNsw1aArqlV7VBAuZXige7HylTlaHD1lU39XkQ6lr
e8bQ8TtTuYXN3hghDDJ5Spi1CqAn/wHSptSlFwL0n6/La10EZukRB5FAEUOq
1LJ67mUVY5ieXDEDJhmBrK5Gn1/5uHipKipmrH1JtfoIpMoeXpxtwCkm3pik
LwelUh0jRnqMw3v7am5V2h42dIxq9US+xKOpJhLC4PQa1fMHyCXe/Abg/OHo
i6pCSxXurvkVZL4Twh9jy71QlHhrjkbi3RCAYREagc4B7PxmJ3VSyspb3i0k
yjy7YtBdQkrmfMbu5XOhUbEMtb88XAgwfq8NysVvdQysvDnnKSuxPMG1+/7w
aN7CCeqHFUKAuza3PXruXkP/OWZR0dUTw91X+T8x3UVf6w87i+l0+9tTJGTT
yzNHGbLQYYSMexitK7N89uajjrfuKbrRJlPXpnNCq0qPp9EP54z8Drx4/qVL
K7tE2izp+hpnjvphhAgsBhpw3KczaVEDn1TB463TCkT5QN41eTUpF8KacJ9U
g92qihcRK7X/xE4PF8UqWkHlDfRFucwqbyumF7pnWaFVY8IiuNOIdC44ecvr
3LWfHWKa+LzUERhXRrn5HYHqeQ2O8uz6F/fuiYhG56CGzW04ovG8SJzLYZtM
Qe/Z5B+A2EgSvd5XtNn2F9jQIhjSSvhzYkGBX4pUdK4DDKvzZSvjzmh+Jooz
sQtJEb/XBJCXVlW7Pn+qOpffmnwFxv8aBR8LGIEmbmjO98Xta1u/EEA3wxzm
97oRaSwYppQBIHtQbCIMQk8SVce8cDk7mtUyxCcV/s9Eaha9QgI6cD7Jawhw
Gy6bvl3yQmGTMZfWcBBNZmuvvJ6kZpUBgvIlrX64txlNKYdNXmKnPQM7FcX/
0YkEPDq/VWH8NiA5pp6MiLnk3d1P/iN3TAfHz6dH0g+5Mie12whmtRW00zc2
r4pTkpSaliUo3152cM+ipGLSoiQ58DpJXLxKEzBoaQwdorRs9nAHzkRiXdpM
kq5sXuaRWTVMwAETfNKQEl+VvrAZ3oUX9HPca6mzvOyTBdDmLAVocpntLEe4
N8Nvu02rJNMwj+gTfzQ3bqtpau0wokJ/Ie0/r1MkSDy7tz9SqJ7bxRG/+pEt
1VAxPFdagcXkqxPHmavujq+cMQq9d8y7+wuD1Vx7f8cEU7Ht246RE9hi2hrX
sZwfL9Ci6a4uivVjN+C3o37alJN+wTYxn41oPNw0Iswt5tSm6lmK+KKPuzwl
yNR5qQtS4wT6gcCOBJecn5xuXL3wH6TJBv249/XvV2c+NfMTgLCrhMOera6x
gCmcA1vf4OUpSQhgAsZrY6Ec2pqXuETYoKpyMOufAEQ+ByA15NSxzNBlVrAC
Na2gJFPWdOlifQWvwlHd5GeitqdSnvgDcsYE3MMNLDlfOywsyQm/ywZwN990
ghRcK8c+eLTgxpZOAVwO1wcRsJkuV0XxCrVe+aZn64PlC3almyACNLGTjruu
PkXKY8jbk2YlFGKd/NUAf0QaheV6AHNH69LOiZao2hIz/H+Y8AR+dTIps0OY
XqF5Z8GGIZ6CwFzpyeSS38FVPypM/atGJexbavqyGOnDBUg3xvLco9ujyqfX
txdKfpNDg7iSpJfjx2gPwWI+L4fNJLzbgj/GPlSlOG1S30HJ7WjRZC+iIMT5
l2FJg11iwkwAAi0+nuZPyIT83M+iIUpGhCDunz0TdC71txgqa53e9Ee5Z/6l
MMUFGPYajxV80Fg69ZnjPNRgyjh5kZJoE5LSAyEAvqsb69TsB/XyTjuODNOR
WKjsZuI2HoTBMOqTt5IwBeMa3y7aDrb3tj5mYcrJn603UcP2rnXCbbDI90Pr
HS9/T9EZLdOVYtWySH9rX+rm1Y//ZQG0huTvBQEPN3HYDs4VPC+2lp0LUkKh
oEpphi5sczEd5kyOJ88HtF/eQhNcPov6xNApVIhVBeTCnHsiR5OEKE26KEvG
qH6OSRR2kCUc4ahW2AO/l1BN4CVp+kdiuIxxbDvDFX2sUyDjCpdufTobEgnf
19kEUV3Effq89iKioEH4bPO03wz+R8ivfOC5DzKQDZtT5zv7UQDTrnoy0A99
GVKa7EUumrx45RQ3YAbrJPRwVFaQcNJBft4pVBuUaSrk7knY69FE3d6FCrIS
qRU0HZpqzJByXKhtLyHtF+jZPDFOuuQkO9RZBTck0H9hWcrLkexBjx6LHxG4
Qux1R+Tk2FeRn0+8ovDbYiWQjOzltwmaF3Kp138+hwZ9LT2NROo2kyzQQkTF
uO88ZTR0bSjuY3ccPMUv1sLNn7udhjc6DoCrwnwb1u/qgZbvdrj9rdgk+XMd
04HxMkedwz2z5xeylbAOsBorMzKaY1P0kY5VN1yhhoAIHNQOCEHDvu8vPBCw
fvoxiWuQq1hUG8SlVtrrSgDZIiglrz/2ztHP/EtUJ03RsGl9pQouZcsGUrXh
OVE5zYF0jne7l7U9GMowyEddJG/89txrgGt31NRTDeFOPQGXZ9alw4Xr3ey3
B9cE7IQPEa9cagBch5Ryl2TC9d8JsFh9cDPFXzpvyWgcAh4rkNqhL7C0FUsJ
rUVw6U7s45m3GrN6bt2/9BQKUjx5qjg9wVLQLPKh1uBPPs/8511UZKUsJMJM
DoBd6pVS3z7kEb/k1kDp955FUFR1uUkAJkVgWUOxpHpc2qyPEpzcGFC92Shd
+DAbfJLzofKV2kPhtd2hImU9m+5GbGSO0MNVhUzFu21xq/u5gnFWBR+k81Fe
nUQ+2CLBLZRqQCccQzIRENxma0Hjnabo/S/dBQnQoMzrwj97zMZ8mimd+PB2
3dMi2wWCyY7EKQSDB+J9rDTHgh7EhtFH2thhpLXVdgrXmU3HOgpnjnSjnRR0
UFZyQK/S3+jqWYHsGnYvb5TOqqABGx4M1IC2dgkxUSGNuWc5SDiEBvCZJJup
kz7EEyOnq+Y9OaHi5ND2rdIavu9JS7/WbFiYtNNoiKkHgP4iwcXc0zqyCaWg
XHGuZpHpHFl7K1DGj+aVkNhprVpgC4eyGGmfTzK2T6BpghbvowPcLzRiYTF2
OIsJqhaOW+RuwFuUnUO4oQs1mERgt2I0HFVqsKINrvSCYzXGsdydiCLzky7Z
oMg6YDOsgFuuN+OJlcNyCex24v//RXABfHxd1vO0a3S0ysWn8D74itFkEHYl
VJivCudnz0nYffvm2jgEcRpej8fBu+pqoVQf41K5NPiij2G/Z9ftMOqIV3Jc
Hw73ajxJUDyv0+HvlezLBvEs/0uGMR17q+gpOhh8Y6oKJM+9IB/x6oZaknTF
Fph8MzaJHsweLMtjXyHiFSRzE88HAbuv7KHo99pZnpapUy8YbFWsXPn7Y0wS
tdeimuPoNgc9lDRFFhEz9AlbZYtmFy6F/rNstBdwgBFH3xegc6xtPpb6zMFm
8yXyyDz2wtgGuuzkVPnpvdAxm8AH96Neu1+DfDG0h+jJOWts22rYCI3RFttg
1kRq0zNWrYwYipf/2x9Qe2YskaeRRuHUZqGfrYfTkIbB+nLJNxNcvg2Jof7H
C+FMC85lweIJg91NBwaAsxCZVB5Gmxm//ei9NC90jfVOmJV9ksGVdqeoDYRh
S23xbebcCrsym6eJaviUXLW+bem8pfXTaiWo89TnVNUELBttciIJ3YIK7hCd
h1j0PyOOWI6hi6c7j/DVNM+N4NjIp4+7Qz7x8QoSfT5uIyqoa1JVn0swogTj
x3aA7HiA3vMp4v7VcLZGO+n8IP9DCF0t3nUUHKAMQ05nGgdKSZwWtnIexO6o
RyTyVJcq2YsjlRJFnfCGc3kkJPFdtXSvAQKG+uUgHiQDBG0gspQrRVj6Cpvr
ZeWu63m0I8iQ1euMwC0FlqarzqlSlmb3WpJp34o45YUw2h8KsTUdLUtEHkdm
ZuTebvXY16TKXVKIaaJdpiw3EXY2KrudtprVp09zhukpoREJUwfuSWfKB2o0
bERgiLRn4r7QKBKeOX340mET54BwJTSv6xrroMCvjQ7zDkx3w3bER2SNjsuU
LMkKStBpT2qsZrGDnBETL7SGgMjXpBaRzijZouHhh3qEqq+HYM11PkICH4zD
5a3bQFtzCHJ/4S70IGcudTvoGQRRIFpalOteIMLA+ZFsKlOFEBjv9zCT5mcY
xoOB76m7Rln5MrTSyymdURsCUFZxRCuMh83LW7E0VOZNgNeaWOnXN0a9tLH/
F5ddXud1aOWA6nopntZFC2hMyc5rx2cp9F5jHSJx6VW4SsnTPgPQD1PcqU7z
rQSdUawxAcVL5yeB6YVW0VQe+UlpapQYZxbQkNSNYkkkR3lnbxXb7bmWSnf2
6blrkXgzfLuVa3fEQf/fAH8nRtM3Mm2mq0Y2j+B1zHygDK2IcMshz5FAdraF
TYs4XhAiWJAQRvXfe5JdTwMX1xzqS/5dKqWgMmQftnHzeIBC1OidY955713s
A4GAxSoXY76UMfQHayqifuZ3fZbp6dJ6XKFo6Ri6grF1A7z/r+KUzUVEO/ES
sEUrupWfYnFE/LLDC10OUG9SwkbdfM3jTNSbk4YbikEaIKYDkFcXBUq6MyCY
kaaUc0ztcBjYsKWZXP4y+yN9CFn9XsY3WItvqy+HULo/yuDOK+E6fi8N0KDf
6Y6M/9EMsIFIKXKxjVvLqW4VgixWgrlSLdEqf2+8bdumJ88MqLvjKFpC+g4x
nIYxP5iQo9qP9Cz+9PLws8b/tu7ZkIfFTMcHqv4MQWf09unIl58VSvxBx6Vg
YIM07ABL2glx8tMVcEQwJVO/pBtxjy7E7nDIjkrXwqXl0aSSo1L9zoA4L1mK
CRgntlPj6trQAAjMO4U4WpXz7jhv4iIdT8bh6C1hyBknoiQhQ4y2xdaoSbHk
yuF+lycJlj/yIkIkV9ZBn2nJYjwqdj3jWPx6IdHs2PB+qJzC4EFcprWaDJaV
oNhpCpS/APtafS1QpWLoNbH6MKGBdzG5MtHVYFBR3EDtwKBuUxvRECPmaFjK
rRy2pt9txsZK90bvOQGmeGnPUau1oMFd+yhKu0sRAwyOeUERO/TfmmwhDaCK
nXAeRlihRY1azDEqSgZMqhPZQr98wS7KWMkbc+H9I/FAnW0pf63PooFTBQv+
mPXyKYdlHKN0CueS7smxaAACG28lEa4HEOI5mYidN+nmab2OXgetmTpvU76q
8Pt4Wv6+WmiBjpwa5MaU65YAujnj3AH2VK+Nnhtc6fwQLa9JiojJiDz6RYUp
O8BQfOjeoEOrk/MEHbc1FkBjO74IbkLHPTzhD4tps6SEHn8cdVgZdr3FMy5V
oEYyRM4bx7r+nzia4kIQ2/1QCuuhyPWOEpbT4eCloAQwET08lhurC7vRKELB
BBajW5bAE69WiXrjsCCE9fSFL3dk+/RpjGr4yqgEjpvwgdeaQjZRQ0Z/7V9s
HOlIHuxZHHlD9aWkmddeta83Cb8MB8Zmv2CjX/vt7ZooV043G8peKGezMnq9
c0nox+KqBy5n6ucPUDHxptrU3oNzBw2szVzwIFsADluP6O1Oq261pnW5e9iU
LFZQSTe0boxf6golbnIv8Iy83cKXKJ9gSWEGKQKYBWFdux0GcWb6hTJAxkdO
EoJ8R2Y6DYs4qZywUmAZ2khvnoAv6kR5WGYDgQqg7NUP/wJest0smfROdbkF
lPooS0CBGGc9NVTHkbrp2gurfaig5mbteIg620m+bzUpT6uJn8VjdnuA5Jv6
C2qL7nnZOexC3hTzeui/rz1dZzk7D5omCXJA4ooMMr8HmFXQTpFyhydaTFwY
T533ksdzEpmZuSKZ/cDjCT/TeSPp9GCeTC+L9kfzX1jViDyqm02p5NZ/3+K3
6omMHJdf0e0oeo9SM8pvOwgwkAuavCC5wHY+RH08S29USzet9jURNNXnaReH
JKw4UWnXx/MrXpmF9oWGzXBCzbtHECy5MuOICMsaQRBh/6ZxgGK9sg6+rrI9
0zWMeVbnAZ6CNqpyYaPSy7hltxk/B5Y2Jy/NWu9PqTgnOULpe24HQeKgoTPw
f5/DjgTd1OmcWDp3A3bSIL316wBSZOHUc2rh8imDBYfraYd176ozDdiLG6+4
gzWxpGgP+mc0CYaKX7dbwY1B9p6Szh8YcCVSkgirpUALMHQt++X1ljRSSU0q
WD77ylrrRzYFWJU7PBEXxvWGST1CpQMMJOPWYnq++pgI9SIF5PROK+eQGWxF
ijXKvrTbbkajuCL7LgJ0ZYLcL0ghiiNs52OayepDEl/Dh9CMXpzWVGrpgXnV
Y8Rgn64miq/wFAzCJiT/UKv4r4ufxtBoNehkAKiShcYHyVeYjYMDF/AyqnIC
71bk8OdNsuzs0+k6Z/thxRkIY1ouJ3v05B9q8C/el1QpxjPG023G4R4qK6ep
hSM7wT3U7FCkA5wXjFQFJlhf/DuLMmikY6Lm7mAVSBggysIZTMxLMqcBaedT
BQsaLQ25XO2K9KhSJbAePe0u+F8OBzvg7MgOnIewlPylbZaodqT681g/g/u8
8aZMjZxoPUJ3LB16Iui6GWkKSagH7MI7fux+Qyhhih+uyQp/pcS+RvHwjVow
13DiqH/5/KeIP/SE3giROqKappx3lxd2gDWE8DaVP5mS0uwrsZixfMW09TYy
ic7P6YZ9rZrqBSjPEzDCB/tS9vOCLjUDCit74RrL0iCPl9o5DIBirzessKuo
Y+dZh6hkpkMewAMVfQzDi6zuREtgCz/TkGO7mDUfwlhi4bFAs4iUhTAmc2/J
MCZS2ly3fMNdaHtfE+cz05eqQP9zyGjyji3rYv5yaKuUj979Ey1M9DsjbDGI
A71N56wIf4pvHbABLVHjhEVHN3f626xkITy7u1fKu5a5KoIeyZfTwFJueVMQ
mchLR7T5ttva7sCjZZAsqOawHwCUbRsATgsRYbGEOaG3JZpItL6kIg3zDd4s
wbiaLAS/7pc5MxsC8aoPR3uv3rf5eBtZdQJPpTDit6ExVSUE1Ra7N6WW6mne
SAG7Cqiv5YRSWM+y2EFq6OH8oeALYa2czqTFOmyYcIdE0Bhl2AN2eZV6il/T
cd01o+PUXflgOKkxz0YWtZLpIfheMNe7yaG5gsDcjZkPskjQ593KywgCqgRb
OWwQlqu3uPLNy2nzx4nLnDe4p7oHf5aDlJ87Z0liy27b5mpSHcZhDYr4iq64
LEYC696cgllTzUqPf484XplHQh24mw2VYhFPMSRsCVgE/m/4vQ/zd69CgNFp
FID2ZdYWIqdxcp1c56agvx5jfRnPPNd+pJ+omDjQ9HYzCriDJM/qyO4JlDgs
Of5uYZqlX/92X2l1/Yw+jYqVuPnyQ4pBE3v+GEuEeSX78gYNPlcp6mATnuM5
YzLGYfL7Ftp84QIyLmREVMmdbO+Qr8zemh0JAaI9Y4fde4vop5K7lGTp+F6t
hiefaFP+QCMSerrNANkKxb5P29j0ktzToxFLmLLUKOdBDXi0yoISxtm3a/PB
Rjq8F2VmJ4S+r+Z7vsKzQBLjy7RBAZbW4h5OfAZCHWtkFA/gBMFrVJc7eVpn
MsDQis6jlh1jh7c+XD3HFGKtS8Gn6dgowUZNF9/Dt58yHPgsEMWKdaRiyxCa
l3ZaMMQYJIrm8qOX2wWDWeIyOxFRqpPdyBhKrA73Ff/L5S6h/aRzav0LUvSo
zqWR8Z0yJUKrXsfbXVF9WNL2WKS2qJgsLDrvq5w5/yTxQwfWAJ3vD8dkHuX2
2TrjWNUuL4k6ey+Gvm7jU67/OGUSXvF3nLCgUwdau2xNofH2NLIhwv0z+9UH
QAa0AG/IgBnrbdcXCCMCOSXOX21xqvwBA2+oVBRkPI7xRrf8dWgLlMR6EZn/
7VSuqP07E11y3JKWxm3Wai35vu2IEtoe+JZKQ2KUxJ6zHLWQkib9metuN1Xg
UAU8ljTnnhtAH1pgD6J1nArZFZvx+kNYWs5WEGOIa4MIeLjM7i+7/WGRHEPs
QoRZ4bLZXwgP9eGn6X8EPmEiNfaqCKRt0H9fXpOIJcfLek3k4Y5BNbaAqNjZ
BRvhChi86MZCAGbs/1DUGyY4C/TydI11lMac6NtNtwse4CIO165GFGKgNjCW
Ot75KBvA8U29Hcx8g5DMndNrjB+wfNTsupTlK2h2MQxCA1aHWqqN5wmm3qbv
gBgcDhiqDJhOzClS97LrgB3VlMQa2V2KiXkj44TkSXHmaKy6ap4KU3PEkY37
1bAud6zP701kaxqbfjYOjvz/Vc6VVHuHtWpCoHpl7sAMnVjQMl0IQxNuyYUQ
3bJu708iZ7ZfViaM8q8evAswD3DO24iI5B1O//lhEo7uXCNSZ6e+huXf2AQX
iaB++mijixJbR1e4kX1s4PqdeCHSk/xzTVm5mm104Vmb3GgdCUjcpNvv2m1x
o7RT0KXdyY+a9wwdKIX46fXerETyL5eqn2mr49jVe4jwnlulynQIpC+2DIw1
bGg77YqEwt44upwJylHH6c5bdJ9IJ6AcE+BbzWuQC3a/XqFQhhFGsAXpeBmO
VFka+hfd/s4OhMln8/ZRHIwjHeGYdQI8mXeipy8cPqF+mg4vXvIy+rR7dORD
ENTeUP9OhuKdhS9absHEeUUndszpl5YOneUiYLEp1clmOAIqrqeTwjVugffZ
yEPxyNHylM9KMyL2WLaRdmW3grGtzPMNdeEEaCvWjlWEPeA+OqvwNgXUUE6+
QX7FI0KIGSmdnRqhJv81kgjyYvih7M5+AyRSX8I8yHihvDvp4CRNWXuEF5mM
WuIQ8wUlHM7F5gS8KrD9XJkFP0wvZJholNzvkG1eH+m9JwYHP6o3z2g7DeHY
wJKdocXdQPyLj/2qis/vDC+6ygJqrvHdtttNqbXfz5pfx1Yg5gipNYo1Ss0Z
l0FhPLcIBZ+FJOGAi8tUJI7tu6KgXDVvBNjklRbWPZ2F2iuzlWhjSMlZLLfj
hGEoMDTVi4rDEutvot6OJH/9w9GyUY4NQ8QSypY0+F8dHIjDzFj1Y0th7kEm
+elUHTeJJd8XaoLeD/lH9VfB7t3Qe5nsKH0t1TAqViEkF+vU9+zPiuZg0a+d
9JE6UexF7qLcvQn1OF6LK3T7JaooPF5ombrYu2adu2UfsBwBTCoWoaOp925o
qtqUC6Lu/4ORvAiL7M6lwr8kkt60JhOHJOBu8umOHAINGrN5XlGSZvDrvk2k
SUAgdQ2ERK+XpO9n2t18AQt9sN8Oev1sOH0xoYppYRhBLXnC9kqZO2MjJbDc
7k/0MvJTwMnMoMJcmBHtjNVf+1YD6Sc0ZIi4l9dIrfT1W+Q3Z8reIgjyFpRF
NkoUqc29Ngis9DYwK0nQbIfpX+Ib4KEk7rOs5PWgoDFhzo6YU5byBvxQXd5+
SwAub4H/qt4iXrk33VJRZ2AsmemSyp63VEvSqpMlW3Emrh0zidBAWhdFN/Uf
HIprC8kUURDKKva4t0nlOLyjnaybT+Wk0k9zPO5MNgph3JL1ke05u168EHXH
8QD0zte9SGqsaZ6gmegE/4HM8f/jmpcndGMMltLW+wKZ6s0SuogKyeVL8aUo
XQ5pD2t5/lAFQPkNNSrXzGIhFNW3I2ssNlCHG+1oyksUgotOjSQfi13Z1E2+
NWnp/BKXxQ1Sv9O33KmQg4SLjDgQm1hYAhuVd8k7kbU491cJYbU+bvGSsmGM
zWBq355eGXlSlWADBSJG43KBJ82hkzqLlxiC9D1XrSLzbyP4Ib7babpaqXiT
UAAt+zMFk4zG92QTuCQDn9q2ObfUqBxcnjQkY0COhIjwpffOjhb4oHeEpYJH
H/A+OHjE8RAl5TAewIaBdH9J64e8zVIAxzPaiVQr6idg647Yst/JIGyvOUIa
2lvvmuBFsgFWqNn85g0YpzHhH6c6V1fIhyYp/gDaosYmw+/lApkb9y+udEU6
iTz5JFtko+hIZ3mjfQv0usW3wJ30uPvZI4WrgzKHxkp7LFsNScF+/icp6/Tz
S+++DG7v7IqG4jNs0cv2U9Gi05dgSY7Mswly/dzFaKU0mI9fAOJDCogjHhKw
PiFCpnymHensY/tM9KfX3s9yJoOK0gbMvE2bo6jfYCLyQ13ebee6008IGiQb
1XhzyaXOgaVqqrm9icMGWoppd5nJSD731DBWqvKL/8OKeom5Fm11ypGCagcN
lR/3Kppl4L34klKxQ2AgK41A7RCMzXBCrZVW7mFfnOp73tnK1Z/0/P1ESyyh
WfSEkZMeSTWVX+fC9ZgAnAZVRHF/tE8kNuDUapzVzVFg+Rf1x3ypJFQ7bqeP
BckZvTV6lPv3iAdr773rX0kJFCD9NbhDXd+YCm/t56tBcKpmn7ELgDMQidKF
ayCWUHIrgYT9f6FG00AYV+wR5FZ3YaMi8arT4PpBZnZE339UvPc1dHrCmWgS
7W74UvmGEl1jkhnMgr0ZBFNDccbpdt+xNq4n36Lz++cUOhLf7l2AA2x4Wjos
NJitxuBdLdQG6v5oF7H9qHJ7UNQzEg6zTWyLpn4jAqVEKSUD/0+09TTz1LNk
v3RwDRUGCPPVolqklfXfBCCRxi3w8wIv55cBDtaxsI2f07kScv7OkNFGSkz2
BdcLkjl3GGlEzoq+Pzk8Nz/UKKKa08B+EaL8/sLplcEYKUxeeyBK7PiwyDJE
5nuiFYm/yrx5u9//xv9N0KAmTpHI0r/x3MvHDvcgUktNlbABJDemtcMDpXBK
NmSlPwOY6WmaKgp+TeRi8uop1zNTeR/jf3zsvSAS9Fr+d03MOf6PrCvSMZxk
PFMJcJIjaAfkrS13rHf/ATdZsesVBLXAMpFobuP3rMZZSd3wQDnfx12/J4jB
TfVBP6k/PrmnrHeX+f0GOkGCSkv5qWjXPXbij/lQp9KECLGJh+5sufle51JJ
Gt6J3PSDsrGbU0r/8V5Dk/DNmnWAsO/Vc1rxfjRfShjOVudKVd1J2w+dXieV
7uKdihKk5hRajkGOG24hpxlcRo4Ttmk7Rhcn/1VKKWuznI2RLFDrDSHadkFL
wFUbF1rR8ELbsq5pMqnBg0+F5G6VqV7raHav2NzU/96aIFgbEa+LKWgv2p5c
6VJ0L5jVKXULkbcqr40t/jfAFmlxnOAdZFy2hXGg56I+b4OWf3Vx0t+zZUf8
gEu4dkEweAg4WKafQBFPiVZ32/4Rp80XwDhJjBoXHA6maVz/cO+DbCR+IkvN
jZFY+CMVjIJkB+qGH0abj7/P7TxEg11hMRhUq/SWCJNx/hEXBvRRsqsuV3ex
AEHetI9VJa5M8qZ7q7mgFnkvGSzh3bqjey1VPfiuLkKrz2+PAe70a3kETO29
uFUbaSrTFvidLR0xk5ySp82NzeHajJcBZGx6UdV9jeOisVKbhXHTwNo2IhRA
D2jPI79ahR8KGiF8ko99vILQpEsSEvT5MnZQ0+4dRAojotjgeUEkPRcpsCeF
l9DPWW9NtIvZ7MUIIVXL3++xLUpCXT7WIhIqwD/nPVNraQc5cgQ2ChfErNLA
gSsL5yYW4e3427A5HAe1M005xLrF++0VFCl/Kt05cA9LY/uySZP7SU0616wO
5UjFK+R/OIPtbIHpU7fLCuSEdWeqmPQDUh0sKAa8MJAlXiLYo4FY/olgiVha
9mUJNpmCfvOpiAOr/8PYb8ZMsodK9jmf/tl+1uvHx+GlSpPy3wicJSqv3Pmt
XlI1Upt4AcsWu48BoXCwAzQIIK3oqtX5n3o1R1bA6p6SyJ3ru8NIWxXmaxnF
igZxvvd7tEqDHeUoF+KS80SgyklT172voXvm+4x5lxHLq0B4/TJ02gmWbEVj
SmLbzgTiz0XgYtntIcg8l3yFxtgVD0JXJD0LqXD+GRLNGWbVkA5ciH0SdV53
sLdxAjHOr52yHI4l2zPWVJd0EEhokqjyW6wlIovFB5iTS176AEu7qaA68Gms
PdF3xXxgv5dwOpLt2IogfwAdBIgGIuO+gaQua5Qkdh5hpakps7dxUUDibny1
eCPqFIrbNOrvnCCn8MkmrDJB1V8Pg7OaxLS0EEyXhETeuFKoXDSdfATk6yYg
0mkJD2/Plx+Ld4yzSSzZ7TI/qUG18rzwob32zf1dmsFhrZryCrkMHktWSfRh
fdsG8DRZqAivfZ5bLRGXxiwCZjhJr8HLvBwSHNA/oc6iOF063cAEGFMx/2dq
AFIhkmR+MD5DeYd8182P9DOy/C9MKK8HnbHrEsHxM0wwPknFl1FwDIQsgb07
W+jDW1yWfFZ0YnzlKCqWnDtsJ/2o2GL9KbdZy35CJVSonxKTCVJdo7zkT2Qw
IypF9NTwF+eSoIhtcRJoMO0G5erV9kD3l73I9HUjDZ0H9nzpyF2/AWnssRKO
gWnwQ8gsIGsLALlTPnZ0bQIgBXhxMc1bjoyVvysx34EPYFwhcHFN2XhmXfaC
sDmuPGweVA5LDUIMs5Sj0zFle5L6D9vnfcFZiaIuz6mU4x3cew3XQagMAyaS
id7A6C6/FQkcs48/u8CQChYoQH637eoFqfP+0k71/vJ0zjYCnOv1VrjrY+Qq
kDR7wF4jm9BhFmOZoQBEImKhmEo97MdEyNqinizoONsd5eF+pxZIiJY2QJgn
Ez8IjuSavmwvbM/9ADEvNGTZLTiaYGOE+a03eppfgcFNXEKQe/+0ueVMc3fg
Br+xY3hTjcYVuE1HLd1P4WckE4YR9MkSExBQfhCtUCUZvSjBu+edWvbcn/Dm
jA34sPAc5ZL4fc8i7jZcdgkqi1vEEaO1YgcaP6n4A4rGVlfXKnXV2kIg47G6
kpy59GoTt7KRpawOIIimBi7ZsbSf1RIokuyFa7EgFVWX2DRzjQ8JboHwqkmZ
gpN2e+bEPR800L2WnPrktjd0Yzr7Ok+oYR21InoKdpk/oF2qTu5BEf3HyAoP
QCX4wFoSsSbhHDyh2rI2xftBwq4CSLcMkCq7oeg2kYg2gLYD3YZfl6qGvXTr
+PP14aCimcWs5Pv3W6OIrPgS/759JagR6FK7OqWXJmVtkMwbYcBFbWQtrNrK
Qs8A+DQMg60iyBptJLuXoA7DRLugDBzOgC3r8OH5K8oiBoNROpF8Hn4vmzk4
lf9t3KYvCQuWKz3HFJNzXrLQoZ2ZhPwr5J/e1uRT5fC7SkpLaS6gTLWF3D4s
cYPFdaW9Dpl369XVjxiHSHhSl4ZBsTjqo0ZtK0L6tif/YISk9DFm9nzJIZDb
RhUgd+wVU2WZe3poZMIs2n0kGmSMfETospE6G5xijt5cq8Yavks7UgFl34jt
rQzGZBm7MVXxUf/DmUnqbfExbHyGQIunLpPbkYAQZDdnXGUgawRUc7HohA1A
iKMArQhcbwNtmeXdJW132E+mSZ6n5CBzTFCSSaLZswhhzZ6hDEqQGUSvaTa9
DwybFHd3dANzmgu092z8byCPrV7ci1tjvMy1zwKfCfsWJFuiUo/Kq7y7veSd
Gd94FCnQTYVZlAEihnnlm6EG/AIivWo6weJYW9Ee+x4ixz+PMGgdopzXD3+2
Im7kwTB6H9Uw/M4y/t/X2ZZR8vgrQ/8kuGYnNxq1kg6ZbWwnwlyILdP1Fht6
Ud6tzHPNgWzbzMnZKO0eltTeXfNiTLavbtWHU5J+autAzasgJ8x8Eiig8Zl8
ftoWYB2HsYozStpF0E9meJXgcPK+enm+DPvQahHcLcErQb5k/MdwA7RTMPSP
rDSY9tDn0Q9Jxo1yjVXqsPrn8lIzjFGkZICRJSUTYh5G5DpBZFYLzIJhKLxh
TMsTwXYHIJkzMAlZ8XiejoTQx2cpFxM5ZlSdAs9ab91C+RARkpWfvZvGZyrW
Q8X/eaEaDDzeXMcXWQCqgXSvZXrZMVoz1YsTNV1eJlCGT2uMSSF4ozXEKJRD
pmYrF27s7iF3IF3/IlhxBMfccCh6txhOeXTJQwAq2jy1iAmA0emH9O7M5bZn
TxMhKeBlDlIO2Tf8phbf8i+JtiDdsgA+OYGclClQUV96Xn0E2/+kfyC7g6ZO
gSVfPVJ4kmqiAwhDQ5np0sPCYV8likd5WucHOXILP5Pz0VZkWYp045nTKnGx
j7ZoO5LbFuBD5zmmj3hGASfBRUBgDxzetSlEHycjn56oDFPmlMbvfb1Vn1Qz
LIilEZj8Rmr55BT5c+i8tRhbRjnnWaBggm5pfAtsdm0nN/9dnhiWhdMYZZw9
HSubhZ0ZoBD6QlYfs9tAkdZl13P4yumDAGKo86U4i5LlJ6ua1RpHTbjzEaAB
AYNtNZdDzrim1IsYYygZ5JcsWhCIoPoSQLcdxY7SAXilGAY61S6vgb8mmkGj
ck/XazVLVwGsT3KxatZ5YEs20gFr2DpWVnJVteeZEdWuXBKPrYAdFV8udlfK
82PJ24xNo34QY7uUl/SjHJJ8mRicVCanKcIMNee3qJ6Q+LTw0EeqHxZYJvzZ
sRWDplRDsvKhW4FZdetnWQrZS24r3KlRn+O/8qL9OIhIh33JM2/4bhgV2o7L
39gcsjh3f+wzK6CYVwqhZ/J0yChBQJepKSnG+wbSO7fWYN77bMu9onv6EEcX
BS/1uS/uVPwBeFSYUX7CnIG5bwmYfLC4l5K+VRZRJJdIxbJk2vNh7674VvP0
xlOrXOlLd8jPkynzKuqmuAXV1EW5e/9SIf4ke2/QvGiyo+Xet4BQnLkrGaXz
kasl4rWnftk1N+v550nYxKkVyidVcwtBNE261UasBAtaf6ygNGmOhVaHp5Uj
P7cL6B2+oV2VP2f4/Ejz1e3VaU3RWNsSB6QuL6W/r6/z/bVzTkcUUhaYSA9l
RBqll6onG+NLsIlbnPDqyqAQ/qSx7mlmIN6YVcS8mOLBlHG2W17nHdJ9mOf1
tSVMMtdVOgR3p5HGBme5ifC+ETHnrPWsLqqw3r+70lVteYXHtxts0a/TwZ1m
fLL40Ng3uAc6i9+Q2mI0HBdM8s4UgZXLmB3aY494qtOvCCSqeihP4xe7AwaR
RDFJBUwNN1mjQZMEX5ICjfrvIxyKeas3f3zhgxsNjulxHFQmB3H8s9/km12r
U+RekPAOGLmMmYRQfxI8pfiV9ss8+06FDs7yHtL7agF1QAGhYOd49cUeAMX9
L0ZXxRT7DylHaBhP/D5GZurnAXCTSijgkprxf66B9EM+amIFxd7kmwzYu/4W
zHY2u/8CWoQgmqHp2b9p3opJeEctMTL76sLAZ02gUCCftZ8AAqET/g7VLKSB
XhY4k4Ar7umdizmshb1lDeWE8337bw5NE0JBwp06Q2JtMBrn+N22iLd5K/n6
ifimWyNwyE8CnAdwYLPk3tr42/Q9yTqio8h2w+g9qgPK6ODTgTTN9PsDQmwG
Wi0qfn/0G08ULKekePnMc4cXLxj7xu+2ikVvK2K0KnaDSveGHhG5Nx53+g5E
c94Vk7tAaXv57SXVXAOQ3eFun88u4ERoFSVucke+q5KQJGlE+Oy+uzz24NES
v6XUM0LywuQ4ykdzP/DJm5p378z1vg0W6x0TN9JrZA/oKddGGfEaHbimJqgf
tRxJPy69DT4Q+McZQxFTpUXqiNfEYV4BKYd5ef4Bd05AkzSmzWoPQ/rK/vjh
+CNtdAMzp4vb0mkYALGJn7PZOEyxMpaaCCq5MNLlhmZSiot2DCVlNNL5pOdm
wovDvdQdxxon5e+OjW+VEb2zIrWjnCoUVe1/Qb3DkdA79SPQk4RC/kyyjN9Z
napfWFxuCmGRZA+KJX5qM56ovIeYgxSwOp1y7yD2Gx0e8CcDj1OcDP46ynrf
Im/ToskItfCdnUk0o0MJfztKWhDGcfWln0W6IOK8SVtv5BWshWzj/hD+gHFq
QQ+eVv4M39k1YUkjTLL3nKgqc4aH1SlVhA1ugyY8ECeejcKyIZlR/mvnaf0m
fRyilkiIHzfZtX8hLRh/1fjN177AGNACTZFfIZ7oryx20+zLGPZBWiC4x6FF
MDhwGJmibzL8JHQhCMa7v4rUjgZOUy2bUDU3+bbVHjy0UjlplmeQgV6cv5/Q
qUYl2ZnVMidBUqEjge3/N/HB0vFIUlvrWwI2TR0X+NLuoo2AWH29tHCZWa19
E5gLSVpZe78aoK6xKKqoTSHr6x0Gs4uMsPiHiPqgu/JWHEoun6uHeZ+pg1zm
IagVuT/zsQ+1KrU0lStTldSpZB7hSBjacb2CeaQEnzzxepCVm32VmvUTGUCA
qPmybMR42F34kLw6I3qUInYeEXSQ4UzVYhaqg9ciAq/l+ErbfyOhUvxSj8Ni
3KXcsjeH2P392M0itXOIJVXbM30Y1I7Gtgv2FqVYOGEjAAg0aeWQD53vtSRA
cT1LAyPVEy4q3D0SzylxlYQ3zRn2dBbTdV2DLD6DP7OcCyVzcPJvVT6FxjPr
w2KXxa/pTUyv79JzE8UfAAdp9l4NNkSl2VphEYcg3OzBET3uIouoixcuW+RT
vwUa2CTUlMXWwbB5ibWYcAXzZNiYZOPSk5MParh3MRzlmyoC3WCVIyi/OqEU
TbEpGTJea3HR7x/8uWOuHATeYRnmMpehtx2pNvB+gR+2f5MxOacWdoWOU7ax
YHglRLHt7CeCbKEGdfSy07tQpZWmdshwHcHArW+WrwcBaE3YD+p4by1LDajP
X+7mQ+aJ0ijFdfDnXA5fYWxaYeUCiuDtqjdGBwdsj7EvuARpg0K+dNgQtNgH
LOJI24nhq61Z2UHJugoII0bcHZEXZCvbzTWlwPo1PtVgz//QmjjK4EzuKgl3
0KZ7KW7wcLhgBkpUoyvPgG0aR6yqoJcE2VupbhPfX4Zil5RspxiFkI5KSqqm
NXB6bpwjatcka1WC1cMgmQuNRgvR7pbvlYzQVG33aL7Xm1f2EUHcy398sSBk
XNs/MA8dvcXR+8pumog0I1HoVLD+dY3xktyhr0UMXEOBaXEQtvFZ2O1aTAmB
KyEDSWE4xJxd2ZruLjWLWP6dkVHowwt9AXWkSRGFQ06cv+KDLF4e1WWQg6r7
Kgy3m7/Z5/dJAYzpgNAx2wkgBFwjdujUUN6t6ut9do5M+nQN1PBPsLYZ58XG
T3Y65KW56jqvhmgWPqzBzclsMfeNGtKFHQppm2iyRBy7wMWbvPwMsZRfVE8Y
uaOSpPtOLddQmonj6YLCLl/VAUy59Yo69RphOk0QNgmDJcMy1dk7O822ISL9
udSBu/504iyoOHANzPAkBE29ppKiGHTPvj2wPN7HSqkyCkMuOVIRNhJ7IV/I
3VfQQwC6ZdqbKmEGOXN+QbbG/oVEVEVApKadvUsg04Hkg+fMadi4WWtdymNt
cZsC44ngdXNMjHoyOpW/bT/nCagMhviThWEkB55XLGfoQQ1Cl74ZpPjbqRmr
F9BD79+74vy9wu6aBB4l+NjAxNtKYLVdH0CLQXIdF38oKBdQPK3s68G9ERqe
E46hquzfhUdJFA8ObxNcRLJcIw2qhnXoITkL3FtvenjbNVksT/ZEotYcFasF
BneZiW4Yw/2SigxoUbaeVrThHh6T9pPalQrdACH/+Kjejl+UNps2TYgHaJSL
aOGHCiLUKluMSYMjmMn1nCHForFD0ae25ULd6SSuZUjSvZDOiqVuD9g8dHiy
FHy8/5eUxcIfSP4Kd7tgtwGQd4URUCU4smH3mJxlTiudeU9Hyvwejjaiz8NC
mF7tOxTllO1TTOVaKIONyAw2pL/LRSF6quoIvAt6D9UVU5+sFySqP58kCT/5
GfW2xu0+qIvF1m4GDrlUp1sVrFU/tQBB3FeV/wvIe2DY4awL6rmrzZfCjLzh
K9d6NRELB/RDEBdwjv18Jkc4xfF/+B42Euhm1h8BoJYsliBZ6oR3tNhByA/L
VjClXJbGwUxaYddFTSZzNwkncCzxdIzeRuPUtiurC0LGkcbEmq30AbQj27BT
oZGBPRxtoddK87C0SQnbRzxtPK5vYKWOYI+1T2v/or6dpgOW0SibRwZZwrMw
Wqc738DFx2z5X8lCoj9PXOfVKrpmQzVOPjxPW8HoclBQYaUmQ1BCTWLay5bw
8/5kGRIYWedXP+NlNEe7Mu1WqAavQqThN9ikua/MflVJKXSyKitSNEQPTZAY
Wu3jMB8j3gpGYRdw7A5ZyzOIwhYXlHwfzzu+LWJozOWdA0hivtE5xE6Y8D6u
9i7GztNOgtEdXMhc+eDVvpX3dbu0jsigB7cmuagay1t1j3/wq9mDlFfcEDlG
dTiXl8VL0IPyDlWFckQHpWjTv+aOFOQmbcUnZZAVjX+tz7EkKu7rAGU9E/5W
5WsTvZfQ+FbxanXVIF/hT/1obocn0pfDnVcvqjh5nK1wLY9+Gi1hCBoHOHSx
eBiSrE7DsxilvV5EeKNh3hy7WSsBfq2/s+26+e4qVW9r7KJdFeUuBdEvmahZ
zdYVmDH2tkpbXhrA+GO8Ycnp7Iap5trz1AqxZdrBtkBpgvlzKQcT+9KQkhOw
Wl8Hz8YDL9vACdJoX1FC2FL0E8WFp+tCrHoQ2aAQ3u3vXLoa2J00CwTH4/gF
Q2WeDATuaHvXUAdl8p/jxPf0el9kCw5YrDG4sDcyu4KPpIG+P+V1ZZ1nmo7a
/1ES+8fRw0D+P5LERxJPKMzaVaIjYf6IEtgv/TTAziH5z80K/PXQC7gM0oGg
iHhSxuIxEma7Z2gbW5+zKhUW7z6sLWDSsjUy66be98C4FeOSHkfdB7moFmy8
yhj+MGfSYBZAuvdP83DpIyQuFwsNv63dTgTp+xODBg36y6u9YJanVi+K/GJf
gPYAWByyv4IdAjhLbVfmsktLdKChz6Hzvtdvqur9/UPgLhL73awwe0fowRaE
w4uOnVS3nkSnZhpSHMRG0mx1P042JESygoWRz+WD5wV+Plf/XFoOtw8Bgk2y
dNAqYQngzAAwTFr93JwWBRWePs8aWUxIa9P4wnSBoJHxqKSPKWy0vxYVsSq/
cQ6eWPf25Bfi+EaebbyZV/w9+qW/XSa3+q6lDzMOFIm5mprviLOy5hEWifcp
MYuOugDPOClZhe2hJOl+9nbtNNkrMBjhhD+QRgMAJC4+bjOeIxhrmpKt+IWD
I6kMsdRm35V5Brp6X6UcStwBx3IgAmvb89sZVcIJMaK0rhDh6iU6okuHmGWS
twgF6B1TCowllRWz0I7b2b2IvflgaajoXGkAPyczAJULFNMIoo4ybT+H3EKG
bMs2+NB/TGu4gE3F+GmOrexV90x6Ci/VTrvakkg99SkDhxbU5O45Tz5idvGZ
rOSw6Qv99JC3ytj07AfCSW6WLD00THM7FwJ2qhSmKSy45qFCmfsSs9u+xVG/
UF/TwIpjvTwUS2otnl5UilhG5sp1CDQdeqlTfC4p4jiKAr/NbkpsMAON3syO
Z2QMSDRPfifUIV4RuKqf2M/ZP03uFxAVF+nRwPuKaEJRxfGvllP07KyCdMlq
C6MXvX4lGDnjub/SoTY4b0keM4zgRJ3bcKc1QSLdSggVLubaVBXE85a9MIIp
V69LMNcWaNYSb2Kt7fdUDIVrG5MNhqbdPbgprOTDXklyNJg5kN+ngPqURUSi
ccmKwwS8hP1b1uihyZi8bSTkH5AmGzHn9ZqXOwGfg/ZaRE8poo/WIhWtYWQ8
z7RmheDSaixpkPqaj0EtkHz6uXKhdWoYNZqLpmyUBJjLfLLMNCNvJxz1j5P8
xmES7C+v/u7lkmIrnzNETOrMJ86b7bWZWxZWUKCMFzDNdbjIG6fsMTNRwzDE
xwbBPgf4pe2TuE0PU3FGfcmfcqehF3OmMavYmaEc+Ipb0wv0o8JmpHQ4FIhM
JJL0fPOUOt/MF8HNC46souLrxzAfxKCFkMXw5CviB6XmcI8p4GzQZuE74ujh
PKOTV09EdmJEuv7GV4THq8P8g7fmeDL3armWfMnf/1jj7juUjbEWzjnxHNdi
WEJn2BXj2MhM5VT2DXn9gmJ+QM2UQXVb3tZVWro8jpjU5UagVExJjQR54kUT
MeTRcbknl9eeySYdeRrJDR1aljmAyl1aw4c48o9qI0v2Ne9/ot2J5aQ9eUtR
o0yjNhwa3KVx91mH5y6TKigys4gKP4L6OZT6v0Gwc0KsSB/GN4BojUstEpsK
RKbgJKrylLHsZ/R13fEpTKvry9toUrfOVtsUCzbPb3U6pguSBEgmUOZFHQKo
TX69bsWReKtr9dMsak600lSI3yMYfA8tJvmCjYHFXMtx7EaBd59/vHpqjgua
+IiHE4ssqoMKXhiN3+T4PLMEY6A6g/50s6VF1SYZzl94MSBCyNiaZ8rlB03x
V0eTlbY4yuTBhhoAApCJxy3kVS9q4bC9uH+0jJP/YxnG7IMdV0zQz56DvclY
QfZ5EJP0b/fPsuKtGf4xO4qifbUkhpDGkJ1C1il2O/DnYwbu+K7T993FB7nl
HYT+gkfu/K0/BzuOpOJNzvbgyzLtrTWuXhntoGNrArNz8I/5Yrf24egYmKti
UWJRET6VFMk+hZ5jvPj1vNRwuYNUD+cWVW4d+G+vel+ZjUAFJbCCp8Tjt1aY
zjB34QpSKhUO1NTGeI2duTO0b8Iw3C/TvYOW+xHfl9H8+9Q0dppamBR+WuTf
S0vH5nxjPUInHSdZy7HI2PXqnPvv9QEQjTFB3b5ioqR4RMYVRDjWSggdXaS7
rmQMQ49ybY204h6pfcrll2R0US8mm9D/oQJgECa0G2ynHgx+whcpRm9YRiAz
eazHcLKtsdsbrh/2jUiEx1KtLzTaXHNxZ3GiEoDPfWkz3a38M4xaaUOBNY1T
GTck+pKvQ/UluQRHYOHlZTSaATfKkH9KFAOAed67VlIn3o41Wljd+m5kjBNn
2SWqMxVaAn25EUyG9VvQ8zz+Y45BkovuadasaPYjHjAiG+SG6cCwK08iGN41
gZ1QiDVscp0GtBxKoiAJ0fs2epI6ECxegsOQKheFFACbZ9DerTmsGJUwRfR+
R/TWP4BErXczSX8QwzN8EWd90ewrP4C+iBw1dOcAYPMHxdXGR0m6DIQsRnpX
ZT7jcb/qoL6NJ2jWalp0aBqSJdevy+rPXcvfsO1nbnx8i7VB2DFLK4/uxm7/
2mg8YrXSpKz54G23Kf0Sd9/QCQBmh2DvGhYIdRkTMZ2uoLvXAC4RceuNXK8S
VnFckKKYIPTK30y6sTkVIogDaWDTWlnqN2/yaY7gGRkKhoA5SQi4R5fgByNq
5+pFHvfj+/Us/nVQYZIWm6p7AKcb8NYiyUwrrr/GE2rWuYJi5gEZ79A0BmoH
d8RMaPvITgp+65mtXbp7eU0yRWczBt3g2mIKCeebsaW6LpI63wo2OMpA2TMR
mnr75HLrdHcb+tJ565RFBzqMmqyWoOnWMXdGcmJcaReo9dsZezpWcHSmaOD9
3A1jYCIby6nGyr+lVejPeRPLndp9MXBRmEWyQ36SHZ0C8YqrQXZbLgCfmh1I
GNX8mLQLnUwuwQRrLy4c9PkdgL+QXvnC/QRYHhnp9ubCRGZl+C+JkYdGSWDM
Kh1Necj1xqMTVYa/N/2HkjmNF3n4jYYlHlDwyR+tdQYr/Lt+cL9sPgqC4K1r
78lWcYl66tliccdg/AdsF5Jd6HZVIusSD2n6vnYUcBGk+Paumg/siRWMtR1+
qRHLAmea0RZR8kpU+zGy8YpiTbbB+j8wyV3ZXkadjwmJ4e5X1Ih3JVJcLXjX
M2R0pDFiBZOwxVu60FiLPVaSVcLu1lqrqopdOGmjfXX+LinRwHZ4EnpDMgQz
VA1EBM7VnbRBFnCc8AC7WV8Y/ZPgoPDqyZzBQ0YUoUSAcMQLsZOT08fiTqRK
e6eolKrqv5IJj7kZqxZQLm8/Jvn+GiffprLcs+9XOT2HVYMq0Wl7ks3KtMhu
9t+EedTqxglFXYxSS4pPQk/KomRhrHOqownutePrKqIgcOEaM94wMLOOGJyk
cbPdLPKucvIRae1ybqb6g0DiD4Q2xXHEzxORAjvNnjtyCI1W0ncOs8SQZTYl
9fP01zjm00kIYLJ+263WMHFrO16R6y5oynx7ZXmuTcNlUVsbDCQyxTjn1erj
pouQ3OC6DsUN023lWvU1X+4gu4f+VhYFcHDMj7p4zgwsP4Mcqbr68PlXEJrr
qFLB6cLu6MTLuSxMWD17SNKWNvFE+u7nOvnGfti7yYNeabDAYvVlO2DK/HgN
G3wpU1Kp3Fl61bYIeV4dxasV/Kcd0LJNjQGyZUKbMYKu58QiUrigQhN16rxd
BVcTxTlAvvNo+dZOwSId2PziHL8/R8nL0sVMw8fzegclczU48l0wIozSqHLi
fo7TS+zAMMnk50ucXWTQrIE/2c3oC8c3gs1Pmdas8op5XDFGlZMUjXEPjfY3
3TjcAftEoIVeGvtS1dNGVmNG8psiUHx2I43EdD9CtVUU4w8d4esT1gmgJ2mK
SfzViDbi7NQBCKpviXqA2vT5sriJBkmlhoyOH3ltA8duDItNANRGi6zlaMS/
TGVaZ+Ioi+C7dMfe5Y4uO9PLNwQY8EkGNEP9xqzO4ghON3HwL17nAwcGNRaA
8bwR9bBc3Aj0YEIGxbXUp+BkxTxGK5lEaGxqenYnaMq1dEQilt+Lk5rOlFgJ
1aEFJqDbpiyY+tr/XWKJrKpF3bheqemi0Xhv3hPdbF3W92lPk9bP0UUmgnGh
2/t2NzF+PMNtvW4rk6Myr4/Y7M7UysJx9J4uwjAeWPYPX2rnbZxlNEvMDjnd
agkFNI3gniNRv7TTNO1N6BmgFt7lOKoAWausJ0S4jCIGO0vGkw6GSHn2sRBi
gDE/O3xyWNBGypU6rpCWW/L7G8OD7XKuhxn96m7QjF4umdQtdHDHVayUpvrD
SbsG63+xM6pZ6FeS+VaxRYpxydHYBXa92gsQ7q7xjQruUqGKnF/aWF1PbLll
dzIQjLhWFAs2ARZbKUBcOcJtsyB6nFdMJePudtzBhzZLJ0Rfg3WGRlMjrfqj
Jw8YjeI/ELMw/MeN9/cR0WRrrG9r+HyWXcU9cxbctZnjbACUz4O0t608vAhK
k5cXJoZr3QRG1n9z0HaMOrfqhGA3Kxkj8x+UgRKMnFHyXxmm802xGlqgkOX6
YCFqdiGs2YBlGFNsIxWPZWdXTYONSzjvPa9wPMGmZHlLV5m/JmKJF1pKXEcu
FVCTAAHJKY8ocK5Fa0GGKEWDHy/j/W4gqCQGwCU+xWj7VpK2aCrt7uB2Hs73
KHLtHBuiOHa2pTVeWCVZ4yZ0F6VjW6rfKck4tvXB84w8HfZJBUVvl45nVgMu
8Du/CgI4FsmaneBGuZF1oeWQ5i755tk0SYWU5sMyMgEvzRxn5yTj2TBDDEs3
iuWAjcSeS22EvSVRJM7cfjR6tlTOVL7SBBWRBvmFprv796FJ+JVxrYWP0Je6
nzUXNFNgXCQ/iI7nAs0oxccBhS42B/Ujw2+wnMdfMDGM7kmH4qzA5JMenjwg
Gn7fSyODv4QekyWgGD/G/GKzkXH64VIh5VzTgbB1saNCvVPRbYlT/BIKXrfO
6cL6YXWA/BqKOgZevck54w7siTm2AYaQp9lQa0JbLLOEn63WuRH37bIkHVgi
lRgmtStw+BWKUFNfI26GpgylV69zgSTw9qATBr6QgJq7iVlqIar8vKOloQ9p
E7Umit1r0fGVIv6+7fIk2S3AnI4qGBnQgzzIHkTk1Qg49LtoqhTl+OdOFkdv
nb5L+xNUsdffTWh4u39QfmVGUVaPFS2EOgp0SB681DxcUAYUPy1CVh1luE9c
X7O9EOtECuYTjJ86VJy6Jw7hGbbEzbACSnYePIx4xxbpb52e00IGjJeLxVXp
MB55PnnzZjuWWhXxbJZ7M3UogY8fa+/vzRkwFW3n09aS7xKqj43GJTRy/iMr
EfA+cE6WWQLfeKTrTohkp/63JMazk71oP1MWCA0plAGW0SC57rrV1daAbNck
3IZEUTNKh/UCfkzDHWcbPjW7nPbeLyi9DYfnyJ7vvWroexAC7QZVtqcs3dYT
4YyP8JcRSTBD57/JPcnNV2+6yAkuS6pVLfHXa69T2MGOgugM2SgyKHsS1T0S
Ya03UhgxWw3nuColiZkU0fwBAPaPnbjkPEu8b9r9bWrxnxd7OWat1MSbCmlz
CDfL/sUIKwjjxKfGBJymf9DFaP1mbLADyJ0eWY30dkhYtu/Rz1WO7NTkmbSm
+i4nK3oMpWaxZV5tlMvPfVadex5fPwPb88/B7O/Yy3vZAufPKnVqhjSWzPfY
qY28gfJn5jvrqDnqwgMWZWHGJVW1tO3pUo4Meglflis9FLCZR5yewZij5e21
Og/kSn2YPNnC5GszHPtWdZF/fB1XIdRNlZElYGptJGq8+jA5ASTbekBkqKOE
CL2zWzGBoVCqY3mAJpYR0lbKTE20QxgCSHy2nqZV6f9+EG0oqorEWTQxAgFr
oyKX6kDFr9vMujfsztMLXS9VrVg/yFCO3tOuIEPgEe6MkYGe8FMRk1HOBCX0
sf2kPjKEYTdtrOHWYYB32WgySeJmp80zIniI5Waq2N6WyVeGzA9IPQ7/2ww+
rNzcezhp7fiEbEx1n7C+aNhgt5QP9xn3siOq7IYdYjeocbGHVF1HLf17N2P8
7ymMWPNbvh89z/rcSLKhEU43C8apmKy6ODXVuTmkmZegdRXDt2P+CUlIoEkM
gfJfrtCBGL2BO5LCOcs3Oz2Z+LmKLdVMxE2Y1r/SMWV7/eVtzNXVx4Pnrnlx
SOjyDY2FdgwINoZqSqECuXYJQQoOh2x0ohmW5FWmmAPLe8UbAwEzfTmAVK3Z
H1EVg18YArInCY1Vm2FgN0fkIIrjmdjIGiH0WaNbSgQJ2qAvzTYl/I6W9jPj
nDwQuK0KgrGxqfL4lverEfBwX/ZuC3t91XoiSkK+qtgRo/11lvbLhw4bVuGR
K1D+2bS/LgIT6XWDT7AJptN1Ik8EQbr1vAYCwu3oTMhc6vMJ2Jwh3zcm0PKC
v0ZJMVu3jbf6cc+SaETeVMoVpz7lnIro+bEPlLNcNHlT4GmqJy/aJYNdHI/Q
34Mi6Ve2RpaXlJwRftaNjTXKzXEQtaa7Ho5jh7zGOlG5K/BA6MvjVKrmX4uX
mEo81FrYRuyrKPfrbJbUhlV8Sxlo2IqTKy7nbDGpxblg3dE2LH/UUUlmznfN
wBBbey08v5sZlXIAzf/r5qs+Uuzfz0OEd6Jk3UBMHQXNS9v9jQLX1AQn2ykM
3NrUKBHBKqqrWa50zHEYZJCPlNUVbc/AAlYQG4r2ui5S9g6OerNPetctFysB
fh0hgcgJI+cGXFXbnYd9UGA80/5ZPLeumw64rbjNUH/0GXFsR53NwTVqHuev
Z1eLtKw3cGKJUjkW+K/lC7+h5yo0pORr/DqMEo1fXn057KkVj467RBRt/mRU
CMucePloKHIvxOamKpZDsDmKMUpQvBwwXrTU+0CMQM8FfIokuhT771gSepbC
1IPUgDBr8LiZRJ6CGFvLcjDAVrpz0QwTFp9BxJhT8YnzNqeqOpIhyfVBHtnG
kORob8+XT7UANL46050c8F5e2sCm1lYh3fqsoWd7Fc1zPJz4dlsZWS59zpTe
ilhgCaVzFIoLh+DOtORcJ8gzabWPMDhpNs0ZK/boTGlf+p3UFajwTg6aGlrV
DD88vhdq6Uc0hImJ5euxAj0twd/y6BPfLYG2n7VBJYNDDvTD3S+oy65CbKSy
CcWGZb5z48ewvM6zYglbAltPU8ed3coIrv4GCIwwfX+QY3B0S8B0okeMvEkX
Q+4QsXA3TOAtkx3tgzcAsa4RYdwfjgr18zLrcLZmlg/TGbmapu9KaOdHm5gw
qVefBgw1DBh4UrB4sq4m9oHIFn/RoOTk44F8sPMIotR+KNDJxOv8wYAhg7XI
8I3bTukoxoCGH9o7+IfUoe42D9wnv+pNix+pKs8coLv2DqW6RvgC7RQ2d/BM
Gh0sxe0hefzOBbCzuwcG4QO5brvhIvJuU7KO/1kn7kQ4Rb46/JregjnmbPZT
eY0sAuORuz5Sz/fpz0orFwKUH3EpFb3EKZ/o0fqDSJjUcSCUyLLsCCI3qz6J
jYih4W3BEzoIHWqzqmUh3hqwtmDV/ZuM1KtU+kaabWVAjS2ijxepRaa90UcD
w4KHEAax8t2F4Mu4S2SL8ieOgYX6G3VRMH5iz0j4Ci7q06l42dA/Zj7jGi5I
UsZVnbhZ4hLvMtFObFzfcYPLi6pWDSxKBSOKB/8wbJsV/ZZ85NQBOsNoGu7D
z8HTXbPe4n1bUfOTMjuR2hdOB9ma1E8ZfeONRrszSzeJxF3Bb6NQYPlXigkS
Tbq3dWUr2EnbP4cMgpUPJE4Hf86g1ir915k7Wdj7n2DyHR7hygMVH7sSajy5
Qg4MIf6i4ic14v1+nJg5tnnmS4uef2MipSr2vV4HcCiM5A2fjduDetoQtaEU
XgKQmkdel0oxpD5c0YdaWiG0/YlgMcz2ujeRrwvo9iQl3U9yl0KgxUC8fcWi
Cl8lCukSyWpbq+fuZ28J9D4cWakQlSbuqqTYSAwoisQS+w4Sp42oh47TbjKO
kBhhQWVNHpBacjD1qBFtfh6Lmfy0dAvP1zb/TEAH6TWjGD4hc4qKMyq7J1pY
ItC7+F6FM0fKrmV4e7ccCwetDdAxKJ8NKJJs+yse3uCOJ1fhd9xofIjVYC0i
MzkhBsY8fkWbn6WzzPbWQKiMe3lIId8jGyuOuGXoYz1Qsp2BslMlNYX+SFof
ofbmQ/Dq4KNYHNXLQcdTc4ZY871RYKi5TvyaQx4F8BLycH9qczFd7O/Wbi57
3njlsa9FKsGiKScmsrlyDytOOFRXhZ+ggYfiSDBc4FR3U0vvn+Y1u4W93BEm
OgWTofN5sfbtC2x/EaFsE1VTMOTZIjYczIkskbGj+QX+pttkQhKwbocWxjyr
/4LnhZyWSkza6QxDEZ1WuCMBCAh2sf9WGyKYbJURr38PsLmFOMBbvTSWzHS5
zzzbp5qLjaNDbHZe+B3xQGG24NsZcHc4YOXXg7kqgMcL97tPtNd1no9xa2gP
jAtbmFwOvDYVaifbcaz3MPSgCuVabykVWXrPfw38RRoCKeTrGAMuTh9ZPN7C
BF3lLh1M7GMb70aWkTAvbtr4kYyhARGzb5g3KZe/D8wPzflFFU57yEFv7A8w
5Dr8m2cEFOuKdgFebBeOzlDDONkUc/ja/NofyrQHhb0VpmzSCW0ced6DgDMO
Fmn9tt8ti6j2WvN/X5/yCi3ullC9/gQfzUn+pwqTcoekJURuAeXHzcuK9Eil
lqyHTFUVkcfWkZWrsV4TfEkC9RQq6OXHgOWvm61q7BYmvW7ABi6xYaAmsDcS
uvpY31+lvEVEEjnwwvWmTIyYUYo0ySD6ywrSEk98C6dzarrv1CcMKLvnZfY0
7BBiUE73TPr7qU3JcZKni8bD2SZ1JlyjPaI7VGKoHk7h9ZsrUwMFA6ZPtdn4
m8dCQM42IRwY1/0MkkbyM1rFH9nXCoAYZcApUwggCI3G3xbrXrfwiMBpgA3E
7OZHiEyQrqfoCDh/PQi+XCA92yPXerH8BRXuKQny37DxIq9zd7fg7HBBvrpz
cgtpHKTNNZJwkiIaSQy+UMjtBhYWBPYsa4zHDA1hRatm6gu8EIfWcOpYptrE
tDBhb9GYDFd02hpXMt1qJN/LZx2MeGzHPdNs2rczkJo7kxN2jR/qoBs5A3Ko
g3RgDmoGu+o1GnxfA/F3GhOpr1TPO4roNDQdjV6utuECuPWP/HOFyfGHtWgW
LOZ/4+KicSj6de6LIftYlR3TDiWVL3Au/TiYfsrTltPmWVI4hC26Z4+BcRQY
HamdisbgAPYBOseXnXu2InBC3qgvdhC+smDy7N0hW1CL0nnLexL+bfwDd8PI
mqDpCf9pGdMU7Aw5u5wgzGhzPnSgSFAo1wD1B5/4qQyKebNOvP0UhBDP1J5e
hwSgf8c0/zBmR7yuZQaG0lFiBOciTVXxL+E2ke69B1ZZCgQ1wwHctTeIkeo/
F4juzWcfKOedyvjJFTxQO70LhpWXzEWBznTv7hlD8UdRoEH54U0tZwTl4vCO
Q2YoVKY86YQlgbhpC03kylmI8z0KfxWtzbb38wt9MTNdzN70puiJiI0/E1DI
eoz7Nyhw2AMPxDEv2edpvAoOKTL+pnHS4xOe6Tn4OwfezfWbdk2rJ5UCfvlA
ona0CH2pAAqdgwykL0p4EHEOCqDfFas0ef3/GXkM8zcAXUtgzBhRocy1ggKZ
I2G3NtPbLbciB6+hnFz/QEFFltQ6mwkDzyIGa9aPrlW8a0azjDMVx3MUD0OZ
N7Q+oDq/pLUzbaDVVvZu0OrK2+WrvjjdgOvbf/B79Fsd+3ZLyEBqmEUOs4J7
Vuo8HqgURmxAWNcVE4oFa14EwdCt3MDQrdw7ee6/1A2f3N8FyQqNhB1DLHtb
pK1bYfn6nKyU6sltQWlf1VaIsSlrTp3ZAdbRTamGkpqgdNR3y4jYg7XKdNoj
vLYwbqJf7Tq8vi0ysWkW49tV4QmoED6ZiG+wpl6gARSJLSi2NVrM4LLAWIjI
uG7e02DOjvWDT0af8cPYRqoM6CoFTrD9CAV0jWf4DAr+AtobsXSHPThCmQtT
qDh8SSZhjlh6uxLOqmF4e5tT7yWsnVFwoxvgTBBGthDPBriknICqeFyiJUQB
0ohVWeqfYJWUfOhciWP5GPNuYX0E8Rg4j8TEplkKpj0YdT0LbR0TDIBTQCjO
dxgNZEH+DqWClYl3PIjb0TjBHKMo8C8Hadt2RoG42sqWyHWIW8Y4pxkMsxol
oY9BlRF2ndf+Cf2PnO8Qa6u2HLB4Z/fIqSjlQ+UaCZQb3mZsevKgurzxq2+K
/7ZW1Zs2W53e67n/yfVzfS7OiMOCdUwg5jHR33gRs/DthW4YuYXkRyrmEaMJ
TYTqvImCfEOXnyW6rYahefIAEZ9HML0S/0jE7WbdF8bQnJWPXQYgX0KqL9bo
whbjb2T1MyMfMEFkw/5upCvRulZVTIR1E/4BTTqTrsQiUtX+hujZldvD4Ctb
FH59NPSLVhKE3sVJ/P8LjnUxLUZKfsiYOAp6SW3cvCouGM+qEvE0YLyA83SA
ECd2wEXR5zD6WqEKTB9rIapaCrVoWXne0iVf+Qrpuc4IYr9CthoGvp0NgVlv
u26RG1vLbztkhOCS3MZBCVX5sJQyqLnadMKBgMBLYS7Eb5prgOJmc+eM0Y8v
XwC2eWYZilunZtxgllSNqJQ6qGY1MeGx+pLl16ti4t1JShq4HXDPQMZ89qFo
z02pEJUrx2hrH4j2QkyZPr55euihBh3u67vcQ34uXo3PWDqWyckI/fnzR8ZL
JHhnF1QyLRXbj1h4eX6wm+qnFakpOm6AMBiU4YcwiFeVjC62RaHC2UBuecyJ
nkBvdqaV3B2c8be1ZsIIt+rMYeiwwoKxUhiFwTfiUi42Km8fxfCvSwaHTIEG
9GfRSHHX8w/mD1Sbcl/k9UjOmjoIa/m78DbxLp3bo9lmXmDrrVDxIKRwzpOG
iqj5Igo+VV7NJETL9/mxDBIfA60qMrtNpUh7mahq05A4BHACImnCtXSCYY0G
zAfp2Hz7BXPE0rTr6LFqeUAr7qe2hVBXka3AIqS8TpUobzGGlkI6MSOvH0WD
uz0ITnvmRSdWFzVNXZ+8fmPROIdFxnzNMxTy9ZRq5WZpzHgoRTuQIsdzsnCL
1x4OU1yofT5PBgYTxeyPP1vnYPCZ2SOpJUb+KhQ6/xrX3n5/EIAL9Tu2LMaC
Yo4HTpu6+gY9tl+gnWAynNbyylOHa6hiqR/jp2YSZ5BehtYrpxLQmNn0pPzQ
ChavI9JdusmezJpYorfdEfLm89XSCpTge/GvCCUPVupYTE4u6J/axvd73L3K
PO0Z+xg0Y+tC8hpvNBkeysMWwaEgEgb5k02nYDEcTPOXuMDbNXOifRGODyBf
II65m5vIpeVv/ukmZIOOrWJ63o+/TKV7uGiNvZeFq+eLiJLXXBjoYbTcH0D4
A0I+6WEkQKRv55f+prAXv1AY6yQsEw3OaoqmRbla8HZJwFEb/kip5hE7ebxN
/nGkey26QJ4J0SNo/Ogi2gY+vkKiwLj9NSwxAjiRAjtBQWLOoV/FH05uEZg3
1Fw3oIof3/3lPqmyMxbeS5qrw23mrZL2cYRiGtpCBdSgmj6bWKIPGvAjBqAu
MBP131wYhRskvdiOIwG166OBoBWLZneIe5WDazio0CLOMZZEExEn3jYLBfBl
XUP/oRC4xaLQhPkB+puQxUBy5EPmXTRbtET5pvxX2OAjV2Gxe+owDOUbduIQ
wJUQfdawIj6RtU0o9RwLojxVOSSF3lcqbAp1e6GsgM9KlCugMeicYunrRTLF
J3grpV6VKW7ob87wvLNPWfoUYb/A/vfGm4GBAnNmEOWUDowK3d4LEN9ha4x4
ff7Mhm0UrGKNmI9VwFqWHZHR2GMWWEchwdcBGUjgs7uCDdSZuJfzKu9EPaeB
YptePhM69u7jRXYlKBbBBUJ6jY/M8DE1Y6IktI+2OaOwztuSu0AxUnYzmxYg
dUV1VbGh3rCGf2lz6qHiOw2vNLreZSidf/gQ90srkZtOAcqjKhB7yw/pNCdc
UZWxNTxwzmynS2YxKri6EXVYR6YqWOVRbMtoQ5F8Ii/uHcbS7oNz58+sI9A+
fAK1x7VfEvyYe30qGZlXQOW3ujBjHur7wO2TLYLthiPgpXmYind7AzYCMAFI
c+XHnBs7wDq1UW/7bPLNqigBQm64jhnZQHZtXSpeyLnVFNvEbgY1YYWDIqOX
+hLqoeQOTQvxM2mVBcEOulAZTsTNXhYA3f7pPlm+Pmw58M61vQemhO+kmQn1
aQsbXNgZIi2nSB9yHxSBGSS/Bynnnq7hPMs+b1ojTfBpOeXQjJ9ZHgikklDU
OqrALG7BRixtTOvO9jfjAYhesBJsl9ZhQe70WEebBX+iq79fxLkaYUj3PaWr
7rfAib7dCvKkuwC/hyu3bqjp0XoEJPxtoETvD2I/W7y+wEJvCY3NY6/xvaMZ
stUH2A6DgPJ4QriYbUJphnwT122JhD+TLdoydztha7NDNVpziWcXzXPcsQQS
M+WZ2IlTNtJafZ7xRGA8AJvEshtvjVGT5vXRCrwI8JBegRTjyk7rLhj3LTEF
fc+QbomkrnKbGjlCESgDc8hhZ2teDU+mOcXv3pMMUKF+25aLvT15Fe02E1TD
nDZJRRzf9B/vZqO/yVcY9U/2iyytsEspZ2SGztcYwN5/3zWdupAEbZ8evxNr
86flgpBnCZ1FeUCsf+CMunUcExQh36Bzo8+qR6HYjKrhD4A87skc5B5Hohkz
SNJX2/vyNYkBzNK02ilpMAZGIx/cLr3aUuADlEv1Wbpm0yKUnPSE9tKLU+Ty
snP+qRXgn6YjevJ3QzFU22biCWptK2mv6id++3du5X+NFyeW9Ze9OXDk5sfU
06yV3YzqsHXTFF9kMQzlHcvO2q8E6hEaEPp0FC9qknYSBwVvtCoz1BsU2DxC
d/FUte21swbY4vOIth6a+HL2Niz1N3smdVqCsod+WPGS6XLorpkLGioWSZpu
sansfJlgVyGtS80sW024gGIyYDAAnDsFXvVyeCX3gNGg15jH0D0IxEewn/n9
cVtC55Wt7yf1v6QVA3CF4bR/nCPz4X52sSrB0GMREFGm+HpAA0dZo7O2pACr
FvoEodTBhbGWpdIoAvLfx9jTGet9GR7bWl6dULatzOonxKR0xheqcXJBxJy1
+EGT+SzARJQZI5z6z9Mw9nDgsypH1Qek1GJ+Ix5k+3iURXf0Au+VI4S8tLlJ
CSIqtLFoxH42aqyO5H6pIqkifi30ebw9hCjyPwZmLqAv+ypEtsO0mTvXMDqD
18TLZu6IDkbTtkKgQlHWoG/L4Mqzy9wq7TkHjuaEFBgDwDdn/uFFNENZqh7v
4F2aciI/tiQnrZ6/t9ceaXu/i0F3QPFYLI5T+V9du6xh4URTDnk6HvxMvO/A
vUQPA0ElLE98Glveg+QSPcNkac/vRPwC6HS5uAKon8j7Dd6z3UXjwvaxJUuz
G/GvwGshHLR1E4veXEB0+PvDmJDDm6wpi2GkDPsPhplB7wYpcMJ+NvovuNb1
9FP758IlDhrLrhdCasv4Rm9ht4OERxIGzZk5HMhh58YfaTyE5gfEyPb2qYTa
SSBOE6eaDlcX8Efy/TESIBeEm9KyXsIz55QaF0lpp1lDwsAODJ5yGyYFMElw
MyX09d8OQqChWmMszXMsQIxJKkhPfvTnjIC/Kn4/YTp8apa5Ev6EygqInaI5
ecO5eJkRtNJTseX/DNCm9SugJkRsO6qNmQuZGDWveJDnpqhtNyG/xVwJE8NL
vKq6ETJDrDOPNLze2npl/sC1CBHuDwa4E8F1qI8mFtey/vtmWi8why3nwKUr
yWmTX+AhKARd6FQr2FMuqUjdgUwNzh1fXXxWWlOpnwqsviV2f6aGyMjI6q5U
4anj8qv4NoUWVkB6h5ken4nqvLt5knIzaIRXkgBCJmK8+K4+nTvzFbBOFjPf
8s4eTZwdBQJI/C9J6alo8wZr2aPJgrBjDC45FBnNtbhsGjfLQenATS0xnSDO
CzU4xgw0Y1kHk6LKxPmPGjWeNSWgToBTgwLXHEHhO5la1jT9sKH+gTrcEjxL
UI4OGivXsim+0AhkqnjDKqg9ThWjuTZkhtNvZI3sGlNEyxvLustCDJZcnvQH
0FPvcrm6IO4FT2pn3ZNXNmMxKNlq2YoEAh/KoU/kNEIPcd2b1JhNRLje+x/g
kZI47N9UNsZuqqdKK6XAO8+w7XTW37ar42v1HyJ50zL6OnOvF/vG/5gzuGAz
2f1pU8fxZsWJr0RuTiDfbtMGGHFBw/YiBKCpFXYdM/OdzPpjw62XboPUyyKt
PKfqlpqCH/5OhHNxfG2q/7FsWZd2bBtT5VS8/cB8wqzo4X7oqp3rw1Bl4zF2
94Znu/iMKShiBzm/Cw8qe7hpbFh4lDQY5nyOGXzahEJd44HeD0rQmYiZ1zmb
ratySwiKZsKELztyi5sfhyO88Z5YekMAxWhAuBknZ7smzsgnjts4zT4BCZF8
bzHgLV+333GE5aNY1J1ktnSmRNt4kRw19PbcBVQ0kYB7bggw8owflTcnNJPM
gpXfICMy/YoRRSaFgkL1xhkUKeMDVx0Vkt8zBUqYBqd2O9wrdB79BQBpOhL8
n0u6yCXb6tfUoqhPHmlJNk9Gt7wncXxiUh+OTvAAG8LPoPhmBUandmRkuvw/
BDP93qTb/Ez9351mYd0kVx89LhL1iIOVO6rEaNX5OAPgGHKXk9ON120Epl4S
ZdU37zNtEMEC1qJNLdmWRNZvHymW+iYG50LRG7gx+QUoPcBgduPG6u1vMI2B
w6s+Gz6XvUvoyE9U9OkwVeLR2G3mlzLOwAY4pecfv5ljFIELIyFkEtGO5Xmw
Kd/tal2dSbwUlr3ZpjfvLYH3J+Vq9//QmY0eoh601Pri4h0CnPhPN87CdPkt
HUUUtSJf+Ym78T9aW8A/yiZxiv9uE3/sX4hMRtsIuVN5sHmrf2EXQAYTvInv
Jz9jjL8b+/eGOFtYyvcZCm10Jz5jCkGsYlzeO9C9ii8jAy+PRZBcGAPGccXh
jQtgSF0GVt+ab2MfwDfh85HtVY3zYyFlz3hfNfLHLImRuZKxyLqjSAr3M396
bD3nAXcwadaXX4/sUnlyFD6CAJQMBQ0luVli5QZ1Mp4bZaoWt6/XZt72ZBZ9
DRmUDI5uOIRn9wSqB+BJgmkGgC58wh4c9zDAoraYRK1scYpOOB4ArzJ8XyVi
bUIQV2NlfjliU0dsx6DKFOhYxWAgvkji8+KCmKndbHkv3aaMLLAMMAA0fCGr
guJJJr8aivCchon4wkSYodp933sirbP3D7b8bEajargx2dExYifXXCCi8d0X
g57uaxWgwjTmMkNZee00nUFizXBHrbFyAcB3JbSji1jquysiXWHWXdUi72pA
ZTTNEJxKjeoZw3T6GmSmduTbuHP7PJZwR1GTl9x2TMmEQ2gb8LxzpNyONHOc
l1AIYO+RvHs4LERFLdKot1RZPsGb95T+iE3a8f9sBrM3ZL/nkKwWA1yGNaOM
Gg8An0AYMI0fBWUECs/2gOqBy6gV+KeKhCIDyBqVjh8RhSz5JjAcj1kSXkas
IQTBY2e5knATHCGK48qhjFvAolQvqeGFfBT9hkP+iqvkJvX9jO3LsdNWLoSu
hnX294AryJFN/8niJveaxbqRlYr4nT8nLpBcEYtDQVXL3rFziKh5cLB0/gp0
fvfiSj/3ItwBI4oWtJkekdD+FGGpY0ldh0IfeqAwb+tOQiu1pypvgzK3nSb7
rsVjlaNg8aOfiuXf3Djz3rXv4G2cRCEET4/V5n8QD3yuvgL3TnTbV6F9Tk6I
IP3Tub18oYJ4JvsY3UoIjiIWjhwoH+9qjHge8pSt81YU6KeHjsHDPi6vAR/y
ccTd59EIwfWR+veHlzsqLZvceA2dftl6vO4WDiQ7TiffcK1pMIX84IvEdmaQ
B43AuR6cDOtJcwWpgpTvuXHtsAxC8XZveYfLPtlNeXoFYALYzcMYxnT7pfTk
onyN1fgQFZ4bnDM4/kG1YyQD6s3B8Gg3DGcJ1if+a4ze+IUipf1exo6Coge7
k2fyB3peXAdRNwzipX9eR93zxRh0lxNnuaqqOtj88n7D/nNAUKBeSXGfYZKg
4kJOLOlqWCU8uOUGnx2qk3RVTom2l/rtENAc+Cxw1WZww1W8Ag2a+uj8IaAQ
wP40nMWhNu6BKSw7WfQp1rGRW4stsUKV8w5MNhWhiEq7LiUnJmabfREn1pm4
2J74HnDWlaCVohrMd2VG5nkzQI1NDITKGL3mD4imxRrY5yWohaCgLRGWvv43
RbcGEkKKLRUgd4GSrIhdtNOachsstvYmYU13s+0VPeQKs9Ttgi1N0MC2+Ex3
qnHO18sudg5dhVkvYTmqns7mt4piXhzKiFbXd7QfesM21Har8YLiCGqjdxPO
fpDaYygOFYLS6kt40QHGNaG+0ZMY+e+E9NA+60/vvl2g2NVw4hSOKTFATPyE
VMt5l5SOahc1xbiSrwkJTv0O121sttJdNekzjN9BxhxxKdNCv4dKT3rSeqgn
GxBM8eJaP/j6y9Iaflgzt/tzwdEzDExaXIM9TOE0UKMsUHB6CV0sTQGFvnVK
4hbQMFjXX4MFC2baO6C3kSdRpGjRc4/gq+nr/Db1xZKKYZlID6tX8yh0EG5G
3Rb7k9aClTXstwZKcBfuhFJXoI974CPO1wYspGZZexojKuV3A4F5uTSjq3lx
XK7yGCaIIKxTRWG1+BiF8HQRLf/A+mQ5+XAh/V8G3P1DaAnDynllvIoeathC
IwB+F2reG8mU2JwrIpMpTKR54UtgYwz8OSD5t4HdRlQE5osPGiBd3yrzcoBm
LFPGyZKw6Q+RvkFPvg7TgQf21yjt/HkBUUrB2ojvErB+lRRNPRRsYSpb+pD9
IoQzEqPuxG2I7gg4InZGpfktrpONNADe82P8Bip7G5N1+gpXEFs8Gb4b7ho0
qPXp4+zN2qzZZTVZLHaTqMyy4lUDYfU08+/f+c74FGsjpMaeP+Bpwm4nNs95
yEbqnFHjlcLrn5guumVQo54d8s1MRKNqWaNkS+K96bwlih0HAPgbA6TxznoX
1wfsG4oLhGLuuY0NeT8tEygKpAtLObhMw0si5DgX7z+EJDcFepGstd9fmcZB
BhyKKCb3BbjyFDEyr2dRFSC+WDJ0/YRT29Td3AKZgs8Q/kv9f5iJLJEjo+Qe
AFGMiP1AOKLjNiilvxzIbcicwcjzMi9BZ1Axcq6CPdKp6o2O4Wl15Ajexxmk
MWQmekpFuS/Mf64mEhxBLi0XDYIGCIISPsDlGrHZ7Qmp5jW32lr/oEXysgo8
SDPdesh7A2bNN7dxuTbXRIVSzgtZjAnCMsBmRbU8ixrpE/aIgO0puy+dXMXg
qlwskb0+KIThKeHX+lylHdugNquIOXX1YEwfiJarAgqkPGoeu8redwc72BoG
OEzfr1R+sbu4eoDA+8/CtDM5lAz2467XG0pQF8szXvvAVm+V+9AA1kj/KdjQ
9eQdGkQkIy8AKbmKa9llnSyRLkmcJx9onuqWary2NwJWvs5FvyRc2eSQ+Jb2
tge7AgczUYAHef6cCv6x/orlVSKAU2mTUagUgHc4w9+U52y2IUdJec3E+s/O
Zagnoy0NGdO/wdVENCEBF8Jc8uRPd9M68j8tHS4ULiDyEjV6ecssoOuqlLZx
PbvEbsWR1t7CUmVzJe9X+NlMM5GQunqe5cTCfvYAM+6MR/HsHsB2XJPQ9yMJ
ap3CfLpIS+0OKgZKXz1YN05x4yE3f/ltkE/ETJ1Y7XMDoWAP0Q/agO5d1haU
q/+2rKP4G4NaDM2TNR+6xzxL6Kq0cVfHHGf7kL/aB3ulOm9S3vE97078IN3H
Qt7uH8FxCdrEL7fcvFTXhkvd3yS0c4yqVN2BZG3yVlEw7yroU2+TFGO9+gNb
EM0za2cc8UugBExPCoFIahI3w++2LTNlt3jBLcRi9swlsgu31FFDZ9k1Rk5t
aG+M+DSYt8cmmo6i4wpEfSP2Ac0BhfFomJx4/F8UBzmVsk2xTeoAK1kW4tdE
2F0Mva8+OSGpmi3G9rQETPsWB0h+n4DThRjcxnClB+9RPewjJRl+cbsLChZq
OkUybvrPolwt1X5O0EL64AAcS5xgawHzIxOsPMGZn6cZnz92MZ8o9WSMVJec
YNkYFmM1hqw0aS3ulT6JllRBceO75WGKncfWNAFwZVXbsJjPLP+86p2L6Nce
VhujF/jWBcw5Rbtahx3hLFp1kKQ0Yhul9SBttbEWxMlpq0c0UzojrSvSW4OY
mUcu6MecrqW7BR5w+smuvL6YFcYGmR3aot0kod5RzixCQLXHjN2VmTTmYluL
H+fplwcs3UlZSCV3OdHT2t808tRYbkB+c6DPHpO0dLIaroJH6zzHxYUWwG0G
fACEhCDDLsbyFKoROMFoS809mQmvINmL3VuYFPtF3zm49vOBDHLhcmT1t5Af
84vco80hUWvxYI19A2IKmr2ik1tMEPPMUkORmnk5vh9qX/V9+onBUEBJBuyA
KfyutN5DF2mtn7VanIZ/azy99avTSOXEYr40O/0y7JqFlIVBjJum4w36Wccf
MiGIcoD++StIqMSTjmFehBwkCghaLKJZOwlLzQwxz1XLZx2WFcltogLFsBdn
n7Tiqe3eHi09IutbOJRh4DGXHfOSxW2iU4wsrzD5l2DOnv47o9U6MA48QrR6
H7V8rJR/2Dq5vhGix745yzXPaXIBE/QuB8hrOEczzoOgkCzQ46XzVWbBzms9
Nj2q2wkyYjawAoY4CxrmV6edqpgqNI5a5kigqZgRyRmYmqvv3jxRArDrWWKY
b6dcADZQ3w8YMp0SySj/bV94UNQ5PErGiUsYDFJIVq6TXU9gtWOkTjAaJ+Lu
bTE6CbGQ6UxSRbRSBnApxj1qI+/0fANzAmSshVAJwQljeWFuN4jOmPqHTLyd
B7FJrToaDmShWghRWyvDAHqpxuqvp0kTlkF6CtL05/mSxsUJdAq8ZRoVaE2M
R6yKmdSxpwWoE05ixgJ4Q/+Qu4hRsaOmsX5BaAKTOrfcYIpCxiOd/r6XP6Kk
oMkfKkU1e4mrvZU8RpGy0ZM5PhQ8gj5kNvtoFaVlDCWggcRwV5tQLT/klzN9
PffCKEVd2nxrQc6PDRjlWB0QaYml5y7ydojmSaOI1yjP7dr2ZwHuwjKdcFgE
Lear8wmTZRzHDqdq5HjQLCmn23nuZB4GfirdrrMchZCHsk1OKWvS/yNZ85dk
ejD1f0Amy2n/WKf8fOfeRDl8wmA/IH7Tvz6bSAgSYoVuxiOTzklk27kiSl1S
oeLvgFoRMzYeFWos+zbrtvEeA7bdFjXxwGxGJyIB59aPxBzYjfMFVlus1AE4
7nrlqW5dX4Q3e4dLlCAJZg/TEXfFuWH1k7rLDJ17OgfVz9rn3BWFFcjHLSXc
9yPfGc6cXVmnVKBTILC3VfAXWArvlDs+G4LidFUPC6Ef0ScgPg60jxNWsnSd
c62il2jbkh7CJpA7bON0S+ucnXxxuIselMD0G0xGasaRG7UYIjYbclYwbbsa
uYjSJsq9F6yphx9jVqZUxFSZOUHSng6Lc+mD8ZKvuhVZ3iAFSatuOt4s6hM1
nijpp6hJBBDZRlp6uFOW4IPRm0hndHlUTIPRz5EF+vTajiPOhgMp/cYA3yfn
fgr7GsOUv8uV7mZy/wVNDmC70rLvcbz3AqaBccis6nqcRxCQ76L2/J90qugh
niQF9N4yh2udkELrApKYiWx7K1Smu+FlgSGAzK6cGEu1hnhUqyxh/xnIuoJb
W5cpCIPga+wwC0ImeRypFr76Yma4nfXXVSYLjfRJ9+DC2Aduvlc+RoALAquk
GDsv3T11iuIHro5tGnvMEVpsvx6dNiFHuOtA9Q1PtWCOUUZWTRi/fmR6TMaM
yyP8z0XqK6i0vUtWAwGjFyMijrYYoRba8mCLoWryzlBEiQrMAIsY7OVE9l/z
kuSHPCwsqPlSkXg2ufg8xAXIJha/MngRkKkyT8qRRTrYuB8Ks/lOjt4fwuvr
+/sRZR/jBgyG6HNYv98/jHFeN6pmXLizl9kGqddMnipcaXYpvIPnT+byWuye
NGFPUAD4qR9471mvs/QgNnQIFwtP+j7G881GBPgCb2QqQntlF+r0eXT9FPpp
1tFGjwuqqWFqul97CPLOapLWSEEN/BBCZ9Qx3bKwwUXrZBYhIPVnFgWWRRoE
M91c/MhDUtA6x4H/HgM3tMXS2KHKuF54F9lEhX1XaRHvikkgXihwPzHc2MY1
cGyIkLvURKcHRKF3lmWgZLwb3bz4y61EiS0FmBBsMo1pBo4dHKF76M5or6rE
UbUws4WYZ+3KmtFjhoA2Xw/Scwnp3NSEc4s9bMLu/v/EaGxn/YraPioIl2dJ
DDWOiPuA1r2+gA82Q9wDs4F6NDlkuwainbBO9Jq7Hb+q9Duqjs6YUaWRMC3v
BTd1YEpvXI71GnMyXaWDTGVtFkTgvewSS4wc20hUg5Xprlr0Ns+7U+s5y2Ut
NDApA11J3tV/MqWolZkRQoWvTqau1/DHP9yHSUJbUPuOHgU3Xq0OOtN8VT08
NictraTkqcyCQfIB5CIWaZBjj3iNWNH1oaUtPDvqkQgrd91/5UGtHfhQNCJR
f2HAMfrDawWaaeyVqYY0zfwDtflnoN7bgtio6X5mKwpNMWtlLcih6ee3t8V/
Ji4LgdGciPVNupxEzpBKrceLAieAJMZLyV1bfvAVRlaofMXBHkb2GEmwBfug
JmO7wWWan3HuS2agk9i3VnMfzXEmx46iiZzcloNFYujvt4Sj29Poo4wpCiQy
daI4QIWZR7j5mpCmfkoVu3Ixp+Hbrrt56Xk+UJl/3vBh+ZGfUxPFCbxU37wW
Q3lvjuZfZ8fV/EuCmCoKWZlfk672E6A/zr/Ts8idEFeFa5j7DE2A36t02uF5
5G3FsXf5dLZS9rsMOW2Vzr8uDZDicDRWJo9+3CUG4cU6U1wiCbmcjw2fAIya
6WdG+/wC3nqic2snUsRBbd7kxUVc8BnsIIIF3P0ceCH5DodHhSf1KeZyZVmp
JKGjMydqssAGE4ZoM7uN5KdeaTIoHyJ4mFpJe0FRVdSINA8dMzsBSIxBHyhI
wmLOVTice7YzLnuktDCsVeE0GXK1Et0fq8Io2cMhRijpC6JcohN0tECmICuG
k4ttDeXe9C8xtIGT71JIGwjM/oAkru9eTl9G60ybW0I29CIvB2D1bzTkv5KO
9z0GE1af0g4zP/PT5j6XvASusXy91lFLF84WYzskth3Z60bXK0tyFcbv1n71
Ta0R1hEUdAJ1Sd4UTUydL/MeH37no9gp1pNhspvSWqUJHiZdiy0ECkqfLbrB
rHB69Wam49p+QI6FjcV3jFvjz2INUNuMUdsdeD7BE59R5lnJHWYptEaXIeQj
7V+EYnOf9Jb2Nl11nSRy72QVFDDQ6MEicIlZIb0DTnkWuLdYyAZIOFa+T+cj
83f53kE+4GXLepieyGFVrJ80+/1kJCUYS25T5/Pyo32M+Cfi5+jR62U9Zg1D
aYo7aJXECTD91xZ649PBZty/30njjueAo0coRS9oxsZLbUqU8GKBiHUdoskb
VVOMFX/WO/EsPmk5Ckx1GrzcH2L7DRuwoL1PUA03nvluU5kgS9ldqjSvce0A
hdKExu+zDQKDEVNQsdK75+O430Ck3TiHMmN7udUaDXe/d3i6a6AdB6ESb5iP
IISqSXwIPYKrApXkqAVF6IVuCOOlQuNDnXA8xZFKcrGDpJJSrIgvVxp8koOH
U5z4JuokgBNWfrtCKdjRDgItr5uhrWF5wMlagbS7Nce/tMD1OzWQqEacMEnF
zTDxvloMV00FWQLunDJJmXh9QBmT2J6plq2NKI11oT2T7BKqrB6XO5OiRg25
QzvqolygumNM363guC7ifXKDW150aF+gUkaIWpvnujW7KOro1BsPeD71L2o7
FoWvtsTtzupvLxYeInbGClZ8THof+E245eRlTch+lL4dfG7TT7FxU1K6fmvu
z+/yvz+/mZp1KamtTa+pSYLkHGE+I47uWEAsik3z4X5jrotmy95v31oxjKmj
/ExZ2cfhGVcvnGgK41OMlB7ZzL4NF40OTJmzp6XYGPpJZdTCCpJEGJcuOLpG
6uO8e1A2vdZ72W1kN6m+a4dQ81XVthpk5LL4J+3GuBFr7YqlxyPv8r8bywgx
zP2IcVFjVPJSTd7yu0wvD/fu1KVEwtgC0xeo9Zewpj8krge7QO1US7PbQIxh
GENza43yl+R1yhg+jiSMbfcvE62G0f1Zc7wr1X+oM5kKrnithXJx+EuPtEyP
y7GF3OSOi7lgBIT1wUpkvY/Aur+2tK4MbV3GOzTebcIdIctf42/L5J7fdb5I
q8sYJVY+J1TRxwhBMVPWNLkfwhi//PXedlK2B1lQOtE7tzCTTiljgGeJY6Wi
FsOc9vkKbbahDjSRtAxaDJKHugsd7a3+anjfAEMsyZO0oy1K54IMliWLijhn
X0Yin7fDMYCwzPWnVCBgaGKwZLEFb20SYY0AOdwMSgFFaUrv0PFAuC7b2wX5
8xoflGW4SBU32gdiYSl3zNoneqnJTtcBJz1Tfoq4DV4PNHwUgaN43NXrZyZ7
8bVxcAaadNbfhg6TzKptsyrwcd7RBLLS08knDibyd6DyX6OCuGex6ClNmBit
ukPGf1VieS+s+X+YbqTVW/tAPhDlvFBlTyrJYqU1olOrcfWe2jjjUhqIiBZK
jth4HPLYb/IE9qhImgsQo5x4cbJ33JnBZpsg38yJaQo1cFZSB5/1tMz/Qp24
QacjFSrTT3/FjAOY/Ree+ADNOjnc7qzf7fywgKPxxF2LKWXTaiv4+htygND4
62xhJBttf+GP23P9Elk5Oz0tAGB2TfrQj1QoHP40AtYNj3YL8514pRG2d6Qy
gsaNn1SzZODT4JjEDa/meFoTICk5nvZwudFS+v1rBG0BbuMyTEpSZ1I6rPN5
+6jBXO1Qt+mItmOPBZM2fPqDvq1Nxc0g1gBiO3xMFjMA6y8NUA5XvbEC+9tu
clFcowzB4RskQKA5/QXlHpOp8bUdqvZTECZuDmttvkwcBBoiBzBRnXZLvGv9
c5wKFKiQl3yUrNbIHPQQ6tm0Ow7lqa74qeC8SRb78KIHe7+TP+/8Ma7znPbZ
V3yyvvRh2QNWMHjpL43/EoCqI79nN4LBk7Gwxk4T3Mws+4L8XCoX9iiAJE7c
CdGTKIHwHMjKep0LOFyYvg2KnWnTVJ/pSy8EggccMB0RiS1fQikZkBt3mmKP
eiybE5mLp3ReqNNXb/Ibwmaq6lcsrNBEF8DllKsliFWhOA66QY4t0b48/27m
pAmB3CiqyJDUFmyvILL6ytiBwqSDDU0w2wCOZB3IEJuGksQ0ot9iIE+d2cWD
R7Nag37/SGgAqdf1vhcyTI9wwq/I1OHNI2niIutETuQaDatj1o+xy1iDlxVY
GlGXbaXSO8j4aVZLaRVBq9FVAi2Gtow29FHErZXpuzCOKAgd9/ETJpz2m4Ua
8YGEW0LIJYh7WcehDcZ71wgqDZrNy6Z3+hV0pHTfB+HYPlHOqEe7SBQ8rMTN
39WLOI7B6I4Li93hFpnYXrkYxTSo8PBRrv8AtXeRVcoHB03TFGdi/qxyHdsO
ZzJ0H609ieQwChoc0rqfpFGridIYZ15shgIYj6mIf12UWoW11xjw6ze2WegV
RXZ8R8/oVYg1Hyw8nkOaJcj3OBuhlCNc7vyXqGyd0CzspOypm/+fMCDBEljA
w7rwy07Iu5zMHdmkjQI7UDLxdd4ePr7m+4MY/9Tbl2waXYkUHVXXvwVJnHiR
Xvw3QtDNA/YUdGSnpPxmK1W3NDp3tHowJaTu5x6LEvtcNWeO75X99p02gd6M
WpJmMxF/973R3qPCNVlWrfF3FsRXtPL15DkO9cTvMibttXRBUTAkcL4AogDI
RKHcfLR33Nr1yRpAMqLIUaVVJG6ealz59fxBZ/65Ou+DW7MuAgLspVhiAa1B
MDbAlPrPsULux8+YyWq6nBHNbILej2Yg1JXSCbm3IebjwUWpTd6EPYEc8Rk1
BP8ARNg8/tF3FctHsEvJa3GWYSqtifJhx4WL0E7omCqAT7eOu5tQK+pbzivM
N538sn3dX+LXqpBV9yIMqkwEq1HRTQxznEr94QthNcQ56utai31+/Ssph9uI
MLD5p6W2puLQGUmDlyYlkoZGz6I6G6dGHmRoBH0wpHn0pe0fnvzyOGAjLHxn
zc+4hXIevWb8KVOZut9Ayls6JGgTdic9Pl/j9Z6/qhfiWwL4WHBwt4mRSrPE
0JKEYnEP5zTKPGqNQ6+OanR0ZdZ1Hzlx8IzQuhk2DeV2MiD5KOcEI+Bh3arn
15sq0dvM7jKOd5RQQM6YsbTFCVo6HisM6Pmfq+bCD3RvD1nhR9pp9Vp/Qt0G
IrWqVOknJ+A0IKDSFnZ1vbktvoBykIL+KQ3C5VIAB9RJDBLMXyfFdsxvMkT7
KYSef/NZYWcNE94Hwb6Vyp/Co9XdOmgw+Yu30d5VWOCDL0Ma+D7e+Tsi47BO
fki3NSfprwirw5A/0s8CZypDL5cQ3Lh4vM5fPi5vyBaYtD7cBbnullZ+iF6z
kx6T+tpi6fCRoTnB7T5UHSO0Y4BW+oE9h3nzUS8vOudlpPkIhAYycHIblQt7
C9rtziXb/LoeB2z6KuNEMZSPFUDj0WViFYXx8WZtHJUHXMd9uQp606kKSF4V
2FE/cOz/Txl1aqubG/Zsgzn6+uD2/dopXrCHVhaEx7JaxLbiPFh31V7s64O0
iWApWj7q0rySI91pxmPedhnmwEdLGgNkVfkgiZDOZZclObJnIpc4eoATg//4
6Wl8q03VRX25qeQsl9HCrShF7bImMen5Ptd0cO8kdWJXsLtZ/4Q/Ouu8ayxx
7KAsZHPV0xBOPFBhdJrTZVsPnMyn5JjDgcbYDMb9eAcqV2OXIPTKMPR/taXN
tmMCT3xwkUbU8pUoDWnkMoyvdGBAtWZJWG6r75EFNCUlzHJ/Eom33YoDhJRP
wyXjVms4e7yZt7x+8II4layWzi+pTMH878Naev5auniqQvWv8yxirikbMdf4
a+isEx41kVutzEo43y9o0yL+cs69YTVgtqz7cQwDC2xyzW1rl3HFUKbWOvhb
zemxyq4fPIBY7heQjWvvycSKeXarHD3oWel0qiQs5Iq0tf2mHq+lH+wvhp+6
siycf7nPtcUxe8iKbUYGwH7PVN0M8LFsDq/q5Hx0mLFM1qfsT/HP7WANjbY7
XxEF9TRNJieomYHPhYp5Mz8wDumK7/xjLLkRvifeADssWk/ua69PjMIzdg2b
S7PkdYQDI6urPdt6EgJGa0xqdQ7IWIFlDUCHyuFpaiW64OtDRF1TeLyxEUgG
pqRpRUw8jj/5Y05JG6SbTOaVtTJLxfFz9v4GY9tS3xSsJRjqJXGNkQ2fgdLU
34NcAFK9Xu1y5lViUx8wXO85FWWt3/1bhO3Vp87A+5t6gYo0Pu1GoTHRyUjq
HeKlDVfl+z+NyVDx36gbfO9ZGh6bdWprS2m6JCkpOU+T5ssF//JZOYOL+5L3
fieAUQpIfEtuSJMe4h0Jm3xZ2/Yxfl44NOJ0xSeDcbvaZlF9Z4O/Oj4FxNzm
ypQ4NL3iSuwlWhLODl4TuuzccjlEoquH63KWzeHLvSIKuC/PzNPPIaswO9bK
VG0tv4H64UWopU0TnUlaAYsQF2RMl5F9542DsG9RhZyaF7WNOEkg9cEHi12i
7P8TJTUmb84qAj7H6sVskQgz520Zn3ujNgpPMoYrG5GCPAUdhRmsfqNb/Wlf
fQJviQcC1TI+mm5tMTWawZyjVp9pVyZwGWAEXvtDLCblnOZzmODTZeIjufJJ
vHITifuWLrU482l+wbqlQtHx1u2t1pIAqAgmRByPpVoNsH5+bKgUxrkkTxDQ
7DQTrt9pKg5lIgmF+FZ3vwbaMqlYGGoyZN56nwrog8cmQXh8UqOHILosw8do
kgua/tZWb4lvv8ZLykmDjbtlT4CEoZMZvBgBo/JdImMiMUVGq6KWbwRvx89/
eB19kARjGhCLuTU5+arSHZQj9PNdkcYRn2Qx7nkOmWWR10SUh7iYaEhM/hn3
72ZgjcuhSw3olT0wj9jtc6bSkOUCQK4akTiY6hGoytfnDdHeJW5JWXMGs/HV
6qcpW9ObrhIHsfYH+S0KXTUlf1elrZn8Eh6qoO+0wuXEKbyLTeXBjuSUnhku
gUgzf6Bcov2oietd+xR01rXXbIk8ambTGxbmRQj6vg7hyuOPE+4QWZLvVqxr
bRPkRlDo3yR1cWSugefRJE4s5TeiUWB1GcUTRDw9zlBeKDaFVehz9N/sk3Bx
31quoda0gOkFTDGLzCNK8SLzhimwXpZYHyGji/B4zBFp8yGtYpohaK21ONUH
nXihHJT8dSlS0kuXjv6jyM9xIvPyVVitiANTb4C0wYlsDK00+kFrrfT6aogU
SJhhfuFpwBhYNTMr4oCp9mHyy6rc8riO9yvoR4diPJvD2dYLFZrn72I+Bfep
Dlb3zuNogVqscw9cgBAcY7tyz5hjdTMcOI7GxNdNDsk70P+0Bm3NSA+ZqN9j
5a6bnwqfakrgWux01wqQAixEg/l8PdGJvgtXc/3HvctvrRa25HIXQhoZSXpB
8reeN5V6nrUoEpODqdLzfjWTjCqXnri9nrZJoimDtZI/bkRAInpL4fo8yDJr
gxCLWkz6EaPxd0Ud6sWlqRiQUa2OdYgZM41k8jxuCsjY/aSshMTJ6ufRcw6C
LjgfKpdBrvgfvgxphc98B4ERX+JnKPtNMVDoM3WHdBfKUsK8cTX6nqhM/hc2
4fdWO6Z2clrLZVnYvDDjmjz2WOonlUUuc0Hea2UKFzB/oXGt/GRiVxiX5t1m
XJRpDuvj6iusM8luYQ+o3jBEwduTh26t/YSlLp79kelkAa9kxIbBVdioJC+U
EJ1/MwhhhhFXIsAcOqszFEF6B7gyWBkmmVUmtJE+Vp4oDHF8PEzlWdoZDcDM
Cy4UdF6/tKpA4BL67tKt+DQdhWEkNcrV1gb1ps2UJApPYmZKFfNUrssqkz5x
gsTUXItcYVi5RfanQkm+2i/LQXzaqZD+nFfD9GR4h4nSKqPX6s8OzMinlHpF
b3AWnXA4+yEsQ7Op8Ry6RERdIultNi396uq39Q37b6DQVhKFbP960nNbZuxx
kYqIpUdSn/0LAU0hGuy2OCCQ9PhjT8eTLn0uYXDuXsAyUZGb0RrCsJfpA3bd
tJPW6hWBV5azFXwxLPZH4xsRrT15QPT/9yy9jaxTwR/+HOdTDuYZ4NKe3vJU
6jThU9LYMgjbE3aI8BGhgx+Ac70dIwF7RFYfRKhiF4f2/0Sh66gzqb3CpSom
zez6J82nK/Eq3z2D4mjU6Bdm3OsziUe52drednwjvJFmOXhf91UjV2TbxObx
dg1uIZWzWp5ni/7EACWiCutcGnWpB4FSfo1rZLZGT1qz9f6h726fDiEJTGZ4
eozdf848wWK14SSjzCTf9aE0In5SmgoZtK+cvgpnD7i02LPjRBbOeXUi5Bkx
b5CsdhnEJ8fXoeAnBQ7jqo3+7+B6mDzvgefEFdn5mdyOslfgMFCVNLbsiJPN
eo1OnxhR9TqCGZZ3fPYRqrhcyWXGJJpQBBM+rWw2Pp3ZnVbF+90fUEl3q5q7
2/Rwg0rhkC3fseUmD3thAtWUb2Ejy6y/GlzbtpZqX0t0mzmzr6Si34h/Xmfk
qCAt2vN8nKni2AJLViyXuxAz9nJTdmZkpIdSBXU3YfQAnA2c9MXY6eEqF7iM
bnf5IExHRo0M+OngOGXmPWHIcY6P3clSZ3YtsDUbzDeURRStDDvggscjm0ND
7h68f3z17xxI7XDroJQWRGexrxMFEiyWqcx2uR5ut+hOEWDWjSaTDaWQDkpx
suwNu1M+DxUamm9nq9xlsywLmO8JtNtyjYZtu1jHdGJnRwXmRiTxcjv8Cbkd
qWC7eeVeGq+Ug7Vumn2gMd5EDsfP5g6BFOUXYboXd8p2zw9QRPH1O20RUGxX
1XCYAeVUmI09arYVt+NJtpT+AogV+oKn86mm38svkG4rsGVg3vz2rut11JTu
avSRJcw5fWf7GsshLBP7zUXr74hx0LjtYHGcdPMKFR25Rs9OP4LbzraSozEL
sotyJhWjDKoNwwqSNAxOwPd/Fvw4+dMu6t3Mo1S15PSEjrOtHDOYjl8GWM6H
5NQ9rBlKfuigl52jDd/2YUWA24vt1jiiUaQS1f3s5v/xT1QMkbSEIr7T9ZMi
6vRjV4O7WxtCh+wyhsakH4Eh1KwZk8EtyqN07GY17NUzZu14tRkPyAGSn+jS
4GsDnez9Zsu9dL807iTOXNBegmAulRnGEM8BJQmdggGRFd//7xCu/aP8FCy7
qJleKkkh70J/+BQNSSIDRBLm4ApFG9t1IbzRGVcB1G9RcmfCkW5yq9gNXvn9
fpDi76S6mS7f9YiAx9a2z9zUg++eCvppA0WWUVmz6ySfR8acTQCC9P591e8b
aI9Uy7efgNFX+IRDib5PmFY9KIIKaTqlNNEOeWSykdCfoNub6Sp/wGAkt1m/
/u8I/9M3a6/ARXr4W9RGdLUt1QV0QYx8vkNeVCjwirr2bWuBcJzKIiV+jql3
bcpODtU2T3QXtjj7BYY6nvlutWDdsW1zuFxDQ4WydPmkooxY3Oq7ivOLfANG
c1cOvew4ZsNELkqfv2OKtqG7inpLJw+R9Ew/A0l80JZGytS6bRvgOROXBsll
LRHP3F5DYX/v5xQ0c+Uqgfqekb4JvKM/HFz2ZwhHIK4/5eI19q4EGLemgq8q
Da9kzZR21Xb5uncgRLYHBB9Y2QJO8s/edRjGn3iiL5QHTsldt+c8rd/86MTE
GMCE4/hGiJbhyyptfsvAFXSI3sJQUYnWjsnWpRE/yKvzrUWqckDTu5nsHz0O
StNIa5mBwMTNRVMZrG5Brf2cmguUg+OVtQAQZX6fimhqRUkc7IBfqbsBDOue
CDfhviFbsk26SG/EkzBG/1cSEsZ2KqhSt669DxK2QwiLK7CNQEreRgMLg2mW
NXLBuPqpXIQ82GAy6B0xxaqKqEIniansPyOfrOu3WgT+G1N8BrWy8M1oJQOm
z/hJ4qhicnlJ1oPz8/Cy8LCo4Q2fuFRGrB5SRdzuX63qxDt+ZM/iXIUkTCdz
b5QPWDdnl72h46eYYjNqRzJ3UNkxsLHVF/awL327KpimgXT438G2B1sdXLLQ
hDY4asgRRF6OIZpQbhEPX/Re8XejL+j2bCEVkSiBMEDvb26nYA0PiGt4dBY1
JvWCWN3OaWmlgapEKOwQl2iMklvss1p3KfvDHKneo+ZUXRaImxl53RbcEY5l
FnfsPc7i68THUNIRuR+seBUI0G3G9gtjGAjyB6u6d2Gp7SCaOKtqWt4gc3Dx
9hlB1g862FbmIdlWM+wm7bRyCRXJYsoW1xYMkKBnKHuySEC/0zP4ZDnsrTXh
aCNtwDA4J5GGtvC/YZLjUXNb73z0pNuA7cmchvTcw1kE/zDKuhB/w2X18JhD
l2sGwc32zjv9xDzawoSIYgoOK0gHkKBhTHrdzfoE6CgkGjDElwEY3f29Xltr
SDizVOKU12uUpng304QqtbjGww+NwTAKmj+AQhGeSkQR/i0ScMsXEvoEG8bV
GgnjMbhaM5uUpV7sP62PkXf2PLDLBgvFZA0+0/bjxVq08bjkWspG6lYW+uWN
7WT8tM31Dls9GWkdZOchmgY0qpwEbwGWXn8n0TnTkaWqzbP97PZLI1mknNge
LfzoR2AJO1lHMyGAPLe433EIzon4zSGCA8bwxl5CImhV6QgadzsuD6ZkDvNj
x+QcJnk8sVNva9fuapKKOc6EnZODJiOLGkXZtXFkuZPrlPgbrKs3P6ZmLpGv
k6Ogp4cec+M0ZiPMeUrc8EyhhjfwrAbDYPq+oj5RJMQvbmZsUuHBw3yb7lMj
ilPee68owtrXOAXAA26gTrcOoXH2QQ3K0DQzElGSqr7s2TZPvznfbrXnnEVk
WKhEAgB3MEDf4rVYI6PM63yZNBTs/KQRO8Ewwwv3sTCOeZjpPHphZrTImNO5
ZzCOMQfvmHKltOHjl4WLfK3MIoSC5nWh/3nYDpqfWOzeo/dHXz9I5yXtdFgy
OOgSSEj7E/ufdtrAVfn9n1SYsJEEN5ybEsCeWWvnxUXYpQgEooln4vEHPT/B
E1veflvPvYo+9Z2Tj/TgbzEAHSh488Jaax4T/PT5y3x9UeAgj16HN6YrAjJI
KOluLEa/W/bPAn01VaKiXjminAtb4JVKXlyLWI11arrt+XvHwPEB9lAEnLu4
JEHC/Ht466BTd8zW5hulbQViC8B68PuQc/FaspSptLeMCedGipngjkj4jKq9
rOCgbttFhWOXPyROfhjW2hu3SiSny5Um6O25yCSAPSWqD1Qq9xCZMh0XUSO6
Fwb9DFGBrac4BWqGENUSRG5IV28UJfQJI5AtnmmH38e0OFGR+VPL/rKmpARN
M7BAMbyqrNkonaaowSeUw/uhJ9XPQgX50jnDx9v99vXGnaO8ozGPZrow6dzF
vdemsKZ27JXMK3Rk8rc8uIVCwRJOcAms3TZKmvzFI3yDf/g/qMjwtydkFW29
yvj0gFwbjwDAlkjDRK+y2t2nQq8a9lZE2fvaSdxRrnFeqUhqywAttHYsp016
1jtJ9GKhE0RNFL5+cWCE4opwSGF9B0tTMoO4YhKnJ9bn0I7iLOy9T4xQ2qTV
2f9n5mTwLiqDOaF2OUB0xCXjnZo+qe+R5LqleiBi8GFD8Luo82Ek0Rj1Fe/n
lzrRoc6zfhf4TocLoSWQSffZiIuRuf13jj+sHx0L3/ozHO2XIfedtT2sf9uj
PT07XV4TQO5DQsG8MjFXNI75ZUJkaxM6/d3cOapbAvdZ3vQVe+kj+VVX+hVO
sPDxIY3A58qeDUv73k5Ek5ANkLCLrSw/2GmAn2qNzvBp7eo6Y8ucl/07Sbri
xJjwR4MYYlEMv7OjdR++OvW9gNPe+aO5m7eSiTrKWomkHCFpprxMKqsKG0LI
u1Q+ScAv73f2XhzB32fh7gWRtR9fUS4uZHItQzJYsZ8NAH2FHL9bx49nXjNX
AE9gnVKc9OK9cKMdKiEldV7F84BXc+Iv6/J4EbEIgKQWCHxmCOAiKNdSvJXi
zZqXFKlczq8ewRopm/e/SKajHJfklcHVSlAMnVFVA8uYhjxgVohcrTbjJ7vU
vkFdLFnqil4L/VJM3jnJ6CtQEK1rzXTQFc+2lAf2gkSsF5W2nc2mACpIj1Rq
tXOqmOWpNDUbIuzdC8bLvzkEHS7RHzlgmZaXUJELyTm4cWg7tJkDWzQLogTo
xqMfFNZt0v0jjp15qI8VJEeVEPiHoYSTK/kHBfdDwFFidPJTrG5niqOXtwDZ
S09VV9GwLxlbIR8k9GYK25qr0qFE97uVIIKNkUhnR5zhHfqkZwQg7PqdmYDh
QwFX34m3LT5/Cf8JjUhGorIcE+do60K/1uj70YQNzAHMiQMYgzybGVxYYStt
F/qwzyS6Q+Ef/xWX2/ijietODsRdSIMabofKq1HpsxufyWdLc/59Z+d1brbd
eFXSSqEuJfN/TA+KMX0GyPlTzXI2Seo6VetuyNJ/YQSQu3mJtf2WwjG6a+nU
dJnQPP1A2P+kacnlLKcNaQjBjehXvI3BpKmp4z5dsxYZMFRmyNjbPDIaOYMM
cMN34muhCz1XHcG+wj7X2kUjd3LN5fM/S0MY7trf4ekkVo21q6p4mE2XpyDz
fCjffTarEp/sna0tEY3Irypdskq6Mvwcf1UfrrH7dfJHCgXMdhgXaFCF8qTm
sO61tu7U3WxJHhldW/RIICBdyLMzplzfAj5fC9wWO1Gv8eZTPmIU14KuEHei
bQD9J0UbUL6YE9Gm6GoeY4SHEI18uiu+m08+raBPYTHdI61pu2OqO2N/ZoBq
lbToKspLbgG9B6/MtWq8vqW76jebjQHOoFAUVt35tW23SFGFP5HNBjno/qze
4DWrPVHH/OVAFrcgYdgpTNLsNS/0O4lNwf/XPDcgvn1yaTycC4jbUAlZ93YG
Icho06LOzZ7vfCxC0tywZucKHx8KJA07EA7FXyvrUgbX/v3sJ9IoSWId6OQi
YLU+0hL12prMzRANXOP3LsJdXtYv7Q92gZWjw88A2EFgO9Tnhpi1nBoj0g0b
S1p8hG0Fa+oDGt0+POBkNAuN24Xnl36f0g1aVOCkLhOM9tOwKCWKpaKFqeuJ
nVQBHtdqY000tQInuRwOO/3Rhl+/9Ao5kFJ/W6DqupNN0ZKb/6LgWwdLwtXL
ZUHGWld1QBNCZGQMXBla0aoK5Nuu/9eJ/827BQHJsfwIXVCVL3TGFJxQqFkz
TfQGhrBfk9UmmfEzi8FGLQp1OkzhhjiWRIcic+htC9BziouCAXexLLF8uJGR
lRCZRHEWLPHz21IGN2v0pQ4smsXCGzg0eNZrt3qvXDuETgAKl8Bl0S6iiXHj
lVfIwKzQHSeJqnUpjuQjFxjUxbEMmYjGJ2clacDb6MB1hyjQXtpra2FH96+f
JsKUvzq4+Cg0Hjz0EiRuKryRPi3vwDYKn1B9H2HLgeqtvRkpjYqJwS5a1nBS
JiqR+xfI6Yayi+zmlPj9MSDKP7dQku6M3ObHGVH351exhFXn0WtmYsxh5kFU
OVkPOXqWSJ9tJEQqs+S4IU+25fUatVLiy86TRgiodxMQEMesHO8yj1k1GyUz
p0TB9/wVzhCRMRjjuhGHtWaNNwnhBHNwh4U6tuxjOhGDPSagMTD4jNosLgux
ZL4p2KYJh7CZUN/zOeG9n418bN/wRUHHZm9QFFNSWrY6+NkK/D/8K0MMmNoG
7yJDYdJSbdgRVXMfcutcYi43vSsTE0jDUDQjww41UELxWLBWe2zPxwRoYXsN
8P5s6CryJcybix5Kp8g4ByxbqGVoB+GsYaLv9lUolXyoaII/bZecXNKCADP9
zzBWKteg+NdK5JL6e2kudmfu24L5GLZ0DNMU/z01aC6YXfkmyEdqQ/G9MuRQ
SSf/Ch/8qxb3kIfFLYp0reNfTVsCVHk0RAckCll8QwEnSTwiQUvcg0D+PlYo
bQSqYK4sbAwTgsX91+wfvWiLVGCu6pg78GtABDcv9dL7OQCIC9ZyzE5udP1m
GbgWQz+lgP1JuHVbmnzy4DFjScd3ABWksIlyO6rBf/uAjgYmBfpxK0OCV40i
zbx+EkkfOucECUpW9I6McRA+Eg4aS5rIfXOVM9mFY8r9t55mGykemK8YZMqG
emRALxOB40eeGFou/C5XLa9a1nZrHaP9r2iZRpY28zbH6ksNBLTxTr6xH07X
aLSf2U3MRxEuOmkDgsa+e4fNDc+LTx93Qv8WuodoeF0mDMDSoswyxgvybFjU
zQsDquT/apjcunBL2uI3wTob/9OZykSjlcUTnmLGKzRL2t2TkTiqyxzKdlre
fCLjoLcMeokHbIR9oaXx7O0bCvzaXd/y1RwKcFi8ykuqxcJH//7flT9yJfOI
DK1ovaSKejmUZYqgRHwJ+nbCqzOCCaUEKvJ/zoCMeNPqZGCr2vwYKCFT83UV
33R8piE6SO70Hk0lMxm2ZfDJDPrnsrgX+sr3VsRwr+ig61TpyzbeK2WrYZOx
0ZgIozFcCpuDY4kw3+s15qySibSSc9lWCU3XxncFZR9vcgsVaT7iLmyvl/QH
zD9qQ+AVc42mALlUGD8GdxP9ATyyZzcN/zAMYf3ucZNNgF2WsHu4BleZFO2N
CQXJvfjQjF/Sda+DwwXlCdV3hFmrt8WG5vcYVYcUuNgbKclOKOElKame7KlO
491+CMvmUjz6kZABX08o/B0NVNMWwRGA8HKVzqn36g3yzAlf7wpI+QOozx1v
JSTnU7uRhc5bmu4O2/ezP11QWB7zlgiyKsNv9HcnPslZMPpWjKwftBXHjSSn
qN+alzE6Bre24TLuEoMRfB35GBaDNsUpttksMiwUMmgb93VDyXBWuD9ECzu3
iT2BwZPVnotXnNfhplkcvLdRLUJ5OR/syCkdusfPVP1J78XxLnynEYmo0G4C
NA5v7TT2+A2PhEOqYDgxPlv8yIORUAfP8hnQnyuxZPZnzCFGM6f+7NBPigAh
B65BfmF1inl5O4ugnGMznKRAm6xn2m5qCOjsagMyxvPk1ShKiIsK5Rqal2zC
4eN3GwQ377E2umygmqbhWJ3eSzRdp+brlXVDi/gMd1BJcaj94bH+erE8nlrE
oWdZBcXKzvhzu62L+JTg0YNTxpyRQeQDovEGqJi6jdsW9xYu/z54DQSJNMZg
sBnMGy83vNwX5hfa6/p5/A4P0TQicesLeaQ/CSBfT9pBJByGYk8WLGNlBDMh
e8//BrIc26luL5Yhw0bSMRQpY89p9VGQBQkp9Xu5bVhCh6gIp+sI1JNUM7SO
w0A9RX2ZTytBxyrsnlqN0csoQ8mLaOtyHL8TgJu6sP09WMJD9zuy4xDzIey2
xr/mAkhWnn8Hcz9c2JrE5YOq3WDN0XrjYo+IRNXp8lNStg7+8KCJF4aGqrl3
FxtNUflRYcJeRTa8w6S8q/zyJsuS4evwx20y6ZGwUHHKI8/5mxL0pTq5XAvz
t7KNaZ1oX1kT/GJqHlprDIyjNIRVIk0HZevfgsiQ3finF3YhYjF6rrUTRLZy
VGiSrmd2HYRz54DzbzbCPzLkUVBBr2/XRcA/hJ8yk/yBNc+pO7dAT5//V9ds
Uhk1TWfUFMiUVphZKNaSeOGev+XXMaF5IfaMIagx4QohseRBhCgop57RB295
zbsw3HEFE4yfna8wpAhEFzM6CmIUeQzQGI1I/ZPJzVU0QaeEVn6FPkVzrkgk
jf5wGogJ+wEp3jIu1f1r2G4Wv/8t1/DkruUTstkAd+uOcs1+qV99oaJVwq9y
LJt73VgDELe5cv8HgyLxkuiXmLxDW+I/6BFiMsZagQfo/QoGq09ff8N6W+RO
wJBbitVBBbgUXwS0Gb0QoT05eDRbw7DP+yCsoXoZe1Hs9GDyioNoPWra7Aak
sn+HI7UUC36LyHHZhB2ef5xghKZMPgiVc8hXa+2K3Oqc0dG5UlRKFJsZv2yK
zvrT5JR/e7csgl9w+kvNmjLoRm8pp0de0GHexAEAnwZd0Zc6oBfFY9xiUM5C
suPKn4WDNfrmjXW7bEpb2gS7fLrYFNwYH6xD1uCBMvFKHc6GZXXx99etd7BF
9af6OqpkqxmcoZIT+M8r9RwXMV5s58OmlBio+N1EV6YCkGtboGDPJJx7qSvx
qqVi3T0u+NWewovpL1bc4idkh+IrtxyyUGiltWlXzHUpFzPw/944hbSPnPq4
q9QjCCTGwOs1e8kqwMgcIC2D3Cte3ViBHpbnRwXFCVJsb8kdgwVmL1oTvqu0
6ZgTC5RjCOP+oqW4OD9QxzZB/rEJIp0yZolrJdgJtk8tt30OvR9Vh9ixORPN
Yk2rReW+FUuUe1wIdwsB4Rr06i16XXnHu7OuaxHYNgATw9BVkiCQXulNJ3z9
UubLe1CwW8bCtxcN+UlHHH+x1rpi6iaQfBCdmb9az97PZ8B0eHAbymG9lk1j
Sa/B5MJpc6xKCGT5DMDyAwFhzlIV9UdLffpVA/jruwM0cX8+Yyj4rTU7uzlg
edGSzfLgy9hPE+lpaF8IpJ9ef4Qab5y2XofXY7WFd4d+A+3YTHb3bsAWvVCZ
8FOZte2SvsHox36b2E4ewbX/hVm5C5vR2snauOn1R8CkCzmj6b0J2tv07PLq
1woxIjXFDn7yOFiC84a5auSkAHTbQv+KoMNVeI4sP5wvj1Pq3CTOu+ydjRkL
LN6l5ZJl8f4pq6/QDz4mZA9iB/7VJKNGsdLpACkdlT9p2vdyxFsuU1/l9In/
/yR42d1ziGSvdjNrxDD+Dzw7+avHd03PR2G0fbpE+N5aHMRmp2Os9hyO6YA7
XEHUzl2+guiX499h6uAGSTw/HYXl49jyrNJ+FgmXidTnP7adkQ/+UF19284b
mdLvi533EjlN7eOgSIonjwab3CTL0RBgIqX6dE++VMDgj66NZGsJoHa24jbA
1y1r4sND0J4ZUb58p/BjpOCjDq3tt3tho4qiyBiNvo0Q3nn5W0q9CQfFYzak
JyZEEz4FtWvp2+FpMH5K4RvGh27JYaRpcK7vOW3hImLHxoHgj45SGHhYJrGI
cLDdPeLcikMq3JO1v2UTDNIvIRIO6oqVRq/cU6qfJ08TFKXyrs/AB+Y7X80Y
OlCbdURwuu0u6QQmVGAckA2eo3YTT886CrTSgJy0FQHxkbj0kQnW5St1K8WB
eqE0/xzuyf/rijfrUfdaUf8Ti+I4919pL54R5+qRJswZwO5gF2FRtl8EukwL
P2rRJEItHYEyfeCTsjJtEG0c7bU16TWoYGST68C/nXpJzOgHqKnkMDEpijcA
L05u63hr0CO83jy7KQAKUz8GlSJjvSuNdsll3QUdCTOUgsEyxnIYd1Wph+NV
5r/1Hx2dEq8V69sQ66W+c7JAn9v8c+bmuiyBFs6xUCpnX7tOAkJxC8rSJkq8
8aH/y/fqQ9uewxriOBXWlgX1W7tBySC9D4T8sIUDHIv8sljTpk+u8u1+JQ8U
G2EM953GhQJnnKKT9xKBuzPIod4NGW4FJcDm5pcR8jtLDDozq6/sKPMgCjou
o7zZPjYGXhrhvZlZP+5yktiBVkXUqbAvnL4LPOMjnhkDdVDWStUDL5uwcqRT
823q6ndgtwEnc+xM+UVtG8J4h0l6fnCSRPffEXNBiByLXgRc2A6VFOHAHyUF
9XlD3qOr5jgrm/NfORmfdnQdy766u2oilQ82+1IpJFLEGKMNQecwWew86Ql9
v4M4ogftIQxxtsTKC4L6yN5LkE1vjFIDqE97p+8xJt2bHCWJadQWh1nweP4q
0kKMMi1bF29FrpKOs2F4TKp1Bt2tPcshrqqniH//Uh6JTunh/yGIe6yedWhj
6yG+cPhUbnoelEh9zMPw3ulbJkTaXrLYZaeHfEbaAxyQ5Ps4L5v5LzEwBeVX
8WXcQ93ZgNIxBK/jr7vx8sBB9iXYh5C2mesxRkAJ0WTfB9LOkbaA79xKtF2+
DH2jfZZ6DL3A6KPmkMU3MydrA3AP+FCPKUK3UOysGkdHn4qvgPF8pPID0pcM
z3C1HuN5yDFFOinkw6qY4v+c2jDDKttwRzCFC77gliEjL9qSCI+htSFCpKHW
2LKdY1vpphiuyuwGdZk0VfpU+V/mWybh2icU9PrqybvrDhrI71dl2pWL3DDd
VH2KagOQpQBSbkmQ6jfElk+Jxjhu4Fchs1lUqZzAsUxl2Bt4zLVF8hWK8Hba
kOTXbYxGpAlHhTZ+a63y8N0ENwJJX1Ql/830IoJMPQ8Eys1A2L14R+LlVr8k
8Os44/137mmt7ya+VZld8nx2kJTD3VvCGzfeY+o2ZAqln8HBKYVNZXPW8nv9
NeRyiumvh3WAS+vYUtFNvsh2/490lkzRH9Nipa0lO32FFXvbAQKJWEBFjL/I
aQhCOfr4sStauSscQI53/HEQBzn1VLv7M0++u4w/BxZ3+Ll+9y9bdp6x0Nhq
Hbs/IAbKFauN3e//L3GrpxoGAcl8W7GHOacCMSTkuuRrJH6GoT5UmYMSVZ63
K2VB3YIUFzWBTusOrhoxEIB7yj7NSp+5zghHY2XC/QV8QYzrKwerQ5gRz8iY
/aRioQp4lYOU7M3E/gNfjrkKNCVucim/v1wT38KFTtVz/ZZwnMUsjIrGjYG9
75rCdz7urvsPadnKoRjFgz6zW978gsMZos5tiKq4N6kXBLxH7yZgVk2+eRmz
fV5Tmlotf3fn1gXJR46A8rKJkHX1MyyQgt33Hk+w4Wqh6ap+j8+YoGuqg83g
he00sxIthrP4odmvVzUxOjOGT0DF1orkh5/a1BGxj2tGzenSktIYFLPsNs7Y
ZYR9eBojRGAr27q/rmYx8vQ7LCAo6VwUxVJXNi9mXMjIRwzIGWcN9rCiUg5n
7vOMkKo2rqNaaq+WvAEY/919L3qEw8Nu8p29DMUAV0ZmGh2Lvf3k3ve5yLb/
ZZKilBJojXPzBAqSmBWKaJnwxGwFJQefuuPAWftDqUcIzUjhNXBsWm0kpK1+
0pAwoyw3j7AIJ90al/U5AZxUXtDdKegOcKAi+gDKkChaKVkz+MirgTu2tkLq
VTwmqNxSGb3cGI2EKAU1d5WMDXLvbhIta8YpRJ18GVVJ3cIkk+Zh/X3HZFf0
nOJ/xCHuhHYQXeRz659cjAc5sEoELKAT62IJH4HqJFS2ZxZ4NDRv89jWFwRN
Egcozr7TGghAZcOZKT1V+L3T3yy9Qzvd1vprrHlmhSAtbiy2tK2hMQ5brfMe
4ft9cRNqLN44b5VIWBC8MNwYUcTZOgO5Qq9mVDebcLHBNJxiDOaTPFaA7xHr
+2VhRrnAwDscnH934Oew6LmyW/mC58cNpvylguCVVTXkGoxI3Tufvqt0ey8K
igZ792IjBiF0uIM5XBfntXVOeCEZuIKQwAYwBUpaKXOwc4xTAdWSD6SZh3gV
sYM6NTWYJYoPfLSEPDO3qLDGvrX1DGbvYcq6/2BKkG85AGTFX5m+9bXLYd5I
o02QWUQI4k972nBzBcvmabtivg1TgK3OhD+17+ljmXtnE1LaU+VYEmbO45vJ
k8z9+3gQKYHgPUvNslzWhpQ+945t2gfRZ7w3+TGguf5Upf8zhrjtGPn3grHK
fzGefB8RqXvG2siGrHTNOffL7Sn0OUc8tvMSNhAtpbCViB5W9UUSK3xib3AI
wbDJ+Yklg49bCMQMIBRCAppARJJ8qierDsoktEYZfF26EaeOTpRrzr3VJNBe
4kbaCCTQVArD3UDkNA+ImBnDLF1hZx4DAovh5Ode4VnzamS5TY32S7qishda
yyf9RElS95swaKYbmoeRoLeUHnu7SeucuYah4JdPF8egmjrFCuIo6JVw/PdT
0pEw0oXQYCypLX4NySkzrKmDXwZWWz8JVGFljpsJ9DYqR1tHVb+vSBZd+GEX
NSwwH++Ja0fMyszzLjJTl+6Jh9f6KzZJ1URhMHSm9FkVwcymC7OT5En39ZMn
/gjv61hMelDsZSGOITOBEYB302KJKNFsTYCdK5JNZMlV2vc0PHdI+FKNmFq2
507xxuRg7mhIOLksIUha3zNL/CJQ1UAygegkPjayhr133GsqGa8w7fplePL+
R68a7kwXD4MZj+vDg4SBk0dk2DGnVvkduOIIDTEDZOacRUyYD+10Ga1k/qR8
a+5KO4CUIPSav1KKoGvT/3hvll5mGtM0NqmO67dIOU9vjVdyXP012WEv1GY7
pmiZsmscMd0YrHlrMHDoZGCU00NPi0iPMStuoE7vBzxxGn4qon3b0VcyUYQ2
QcMErlLaosrUT9rCvi6b+WpyTz4mN/voEb9/bPDAyKPqwoLGc7oOvt3G/vkx
7lU/4ngs/duOvoRdgRdlbmYk4tcJrmdv3bW5bWGyCfJpELYuSZsQOnGo7GKZ
QRZ2r5ZiBf3NUpv45IpHkqmNMgSPO/EGDnFUvXFnbre/UjTb83OW6xhOMrLP
+1z3dllW/dYqQRCMS+UWVawGKLnsws/F1PDhh7gqhAJoqfvXCpit/WX15niF
KCLg7Sbnta0KMfkKZURfXmkM2ae2cak0ZrgUd6JmFxQpiE6PbtVi0XOJPeHP
BAH0RaOkMD4vnI4An4IT3Sh5ut/XJ24g8pux514yVibJKDmVLcZNtZLLEeGC
cw8+4flK1OKpBKbyFWZz1/4i1LwSntSYM15HVqVymhcORHIxWq3oNkn314QN
k4kxa8VAJjF/V0O89z+qfxfPs3OrU+YuRvE/94O1biTmVs/P0p0zrTyASY1j
8vE1+E9rtDWJerHGw7XhyC2uE0vaktkkZomX80TwZLCcBDQm6e2s5MGHN10z
vp8ZAbjVOag4WET3dpVYvhmg0Mrd2LT2/hJMJXVzJ86sphUE4JyhwFdXNW09
k4AxVRsQepkyUhlcsADzMyHIkH7LaBl0d9rcrrQffB9NzmJ08uUitXNrsdd0
D/sAwKd9IJuti2fOg2CT7277YNsMP7WHq9gBuJyvoO9RR6t9Vnd8CSWJOfly
k1N3w0vcUV0OZ7EoJ7pWI2pQwcHxFz2gc/k6IT1Pubw60bhkeWQF07TZlFyX
YJi+TywN2TM4Sxq+T3pZqotlW3efJ8A1CG2ipE7F7Bu1Ae5A4FSMYJqLgoC5
0/X5q9av8TC5FRGk11UI1VglNy6yLpWAP+PZAtIsG6hHcXMZ8+Iq6wIryuvI
6GemNZ/wfRL5AkfpARodoSgT4UhWWsz1TeZLxwTUSaEoE3bw4xGsGM2xv4+r
9e84wZm6EWoXtPdByjlpNVvwOwsUE2/WBDAlxrYqY/5ySGP6HvEVBLLWSfFS
ty1SojLgvxFG3c3saB0qc7thJju4vmLMbLu61HwslH8h2y9ctCrONReho/kj
BBP82f+kclJPJaUiCa8j3PVl9UaBi5R47eN4poZbg8vYTFRx9RtllosPUn8W
h71zoPvsktVoy3pmprd96U/gFRK76+aEXlUGRFyWqXmFPnQnOB7mm2KAPHaI
foohcjj1iacAnNGTwHilvDyz+7x5eaUlAjby+DS9uYyZTWot0Hj8cp57M/5r
Qwq7hr4b4HQDWMwdihEMtnROxxxTuHikYKbilmgijSDZeEvWWoTcsbgXnRcN
25rMbTgLVqhbuVecWbxfLfR4+dQq+EBoVoWG+A2SGh4cQCUO9pylJc5UtAPb
wV7rlRRJzMLL9B88Z149wi8ayMR4fn8Y4jqXRmk3TFoF5HxXkPoLcIueNRzm
PKDIZhjIMPa78Wf8LbEh3CqQEzchAJH+TqvdWXcZqTfiHUf9sH6YxHEutSRm
63FsLk/8aKhdgVGbzYVAZ0U0lfAZFm2crdKeYvvYhARtq+vH3oCj0UG13MYY
y7H23lqE2+v6vnkTJ17oFs6j3uazvSUyzev++0DiV+pExEFWUnRkFT/HeUyh
+I72gCGu8HzWXF8IqgR4OwUoFPU1WQRtDOcA4gsmKmvkW1yRQOj8S12KYR5H
AdWexM4tCYZV1T75m159Mof3VN5jeSAf3N0OXMWxD1BG9yUiJ5Ga+CRG9Xxl
ITL9Ma93SrEBrfu65rabri7mtpQkNBPuoLm7367AJgtl2LsMk7nvsAQU1D5K
gZMAkYdeW6jVJ2wHst4PGVsFVONu7sfU76oaovZDr0xMxIjB9vgA0cd9C7ij
V9ZTCe2b6bMHOCWC6LIcsDCzwkW9hUjLW/j//qiRVa0qYKeX9IOzbEdJvcD1
5n1EAYNS5hkqRN/0JK54cG0wP4FGCJsrK7I/gAOV+f4g1AGeNnzst36PjDCh
O5EcTcArV+/G36tUlkujnRzEqQILHenRP6x9sKoGaftrWpujm7uwV+Ji+eGq
hc/tZjPdGW9DWkMLhdqgWAKVx/6HyZX+pV5eh+n5I1eou17U1Dmu+rYLmvqn
2Xzyd3yPuKX1KhnaMw+pKOJIw7Ebt1kGXHZHZjrqGCyVJvxTBYc9nuxzbPjy
D7qR98BBo5cbRugzLccFKqzx6d1vIqfm3qtuwopxIuL+NV/SH+ko8UlfStvL
t8kdXuiYkPZZo5f4+BMu1JBgyoATDpICQR29H/KXuCiOm7nwcrylHYePvcLs
EGGgkau6YO5uSE6yKyS37qrnaQ3rf5vW058liTxCLbMX8RPDI4HKI903Op3F
mmBFUlQS7YXAVryYmCGYx3ulZfsynQoiOMXl/Z8XOGFhUKn5YXqqquPgIzCB
nrz/XzkDpivmTpEUKb4TGzC9WWdg8Lm9x3uH2lN3bxApqY14kOICMTxeulN2
CcjiMYLSNe5EwYrxaMEuSF4dtf3sb5eJto0jXk11L1edVXJhXATzk2emv8x5
gjem/gjBwMtn8FfWQU9tB/VtaegjB7jNF3I95YebDRRg9oM8hoWg6OZ9t7by
UzebHtEHyB2SRYwUTg4vI0NmDhOMCrnb2VdafH0zsZa7HxHqC3tWEmv8F88B
eLG/FQUdeTlEiYcxKgjipoH9iRGJdusC7tKzi+IBTZPBGDgwpgVOc8OYGfXG
lZnx9AKd83JNyLjgfVetuOBQSdeBHz/hmXFby4ad48V7DHm99i/uwsepxwpt
LpC8vwithU23MhITUrpNtKsk/bLuwHFYlO2BHhlr2dHUIFSREbsIM4NSfzYT
nwrkSd6wSYGcKM/pv+tXa3Aik3KD01tb4RR5mYr5xaHXEbRS0OQ/9cO8uCYy
j9pSLmv1hLb/WflLQafjIg4fWtMA/fDNaPdgifnxpvORcIShYHD13h96+ztF
hb45flkgPgSg15Xze0utUvDj5yyHplcu43jka5DL6qUqLWgZ2ZfcRiW3Y72D
T6riGq9kP20DxwzezpKWnCYNXFghTODEpxLvEk1WDaimv1BwfKh1KKzyJFnp
ZCjWQdzd/y4g2UtjML8RK6E5/4eKlUcBXaoJRr8ocMlICM1AKwzXFTae6Ix+
NIKYZzRx4zSBIcK/YtDsFMBwAXZUHQqDave92HpTtxqzjlnBA9ibIVRXRfQy
MS2FkRfYSNW7ZoOqoLvV2KXNYCkq7Gn2DdqQy0MHlCR74eBsXHIJVn4oqfC3
JoQzaWtJrU5mnXWMYGY0/az00hxo3RRvSjqwAhK8yf5bKaXZaMu0SzR6GcxI
Isi/XavWyjZjuJw/mypIgmSglrbWFq6duNzzsYcfHMlqN/hwdiSDAufdokr9
FcztAGP3xITmlpXW3mkW+9vksPgmuabRQbGN6CC8Io6BoSiBmS0Rn7lTTeYV
tTM6Bve3q19LOpGmkQsjmNKsMDuDO3lk3o1Hs9I02ZAh5v15hImEyvCpcR+g
HhaFprnYYqhawODebGQTlAIcPyED2YzEv38sThxptncjeOF2xZRDbFrkiaz+
putV3yjGESsBqO2VfOdUn2ZWGDAwtVAAb8GLapEckpArfA/9R/u1Nvf7vzzN
vYSNHuoSBWFIVb++pGzMXslDNBwY01/wYMzlhbWiHUAvVACGrV+Y0l6LyAyx
tg1uJVz5TZFNSMxj5bmqHYUvLfiuohII3oqy5lS/zR+/011WrrV/7yXeI6Mq
YAhiEo+q/oKM9+V1cd2CUtL2A2gx8CFiegeKapUBY4N2nuc1rYBDt8SAaGob
Q3NatzrXhcRr9L1O5CLZi7XAIZj5ZnJmRCwjp7eugZEe8UWvNmHra5dCm09h
0uOsw/BPqkyIG42fIMQJlcf/1sHdFvv6Ddj71UursdCo6YLpVvFmxP/kqDnn
f26cxzKPh0DksTBb3EnEMSnAruuPDf0v6rEg/IIADRjpMZ3HbjOKLKvfjpnW
5Xkn07SNcJi7sLe+2Pz7ri2gzhEl2+yOjnzOMPVhg5d4DceqOOYXwR+Fgt4a
8jc/KMtH1IzgbgUs8WDfHBM0eqdq8txqqVPRov2stgi0F7Jqof5za3+C1Pce
eBiF5n5H1qHGKehCsG1lRgaUtsosQF8p3nfwLEUwfGEFQIfRroDcI1LfUvhC
yry0fg5iCmUVfwUMYr3PHAQ7kMLc98D/JbLWFUgDkm1ih9x+LmWaN04DJXtS
bxeI/E0qrcGWCfjD4ZM3Rh5Mw+gITPNUIpl3bFU3wNd2Ht8wEaZA9puU51eI
HuzhrGss18bOJ63Utf9usBHdAS5kbnEO9NWILH/fHfqojpDbSo3vGNiaWA5M
7w+2zqDDzxiocgNIyB9VdLVLuiuy6zJ72mEQkZnJX+p0tYljmMNo6eynFjKD
PfXFcRUlscodAr+XOOVBZVzQyoar7kYiiNDTG5tymfO95In5z4S8V+TBlUfv
A2vQmzDRm4d1TQJjJ+t84QiPHDUedNwXAnmdFkiPE2gZCMwCQf8NGcW/OqCP
dSXWoKeYtGZKWfwtXBFljp5pm4apSnaHj6T5HQCJc7BgV2c3jkLNlR+w2TSS
30kjFfmClvVtWPZDTSQsA5IwkW38sFdgaW9Xs7yzQUnrYroJTcLtCE10b2Sr
mN1WPJJpOCftA0niMCc5ss+67h6BAqE3A0v2yeOJ0DCzQ2gYREB5gfTaR32P
y17ITMS1KRiMsK4Q52DEWR5sXBfhizWies+2gy0ebgNLbg7o4URXf7MLKBPJ
W/AfVkQkSJZLL+dBYA/tbQzOHEhdgODRE4JbVPNqkGVxAVJfYy3McJzcQcaT
Npl5X7Jb0VTfoWtCWp5IQMUz7HlSUZeLkZQUUyLrkCYdHTkHRPOhqp2kIehK
IGMYn5gweQwlOx40b85+oguCpxwBcc+KJCa7SXo5j9Imnl40U6iF1kceQq3E
ssd7uUgyMEFGlE6dyIlJn80rJSGNwb1uy/HIL99Fmq03qe6BwYPNClbHr93j
ti7yIf/MPA/HUXjyCZilQ7J9qO4k81yCklvSQAMyE/Zw0aJ1gmp9pq3HCxgv
XhIfapzNngefUxhrdV6Il5UgnkXCe6WMFOtLs0ESJ+4Bc5KQpUR+j5KES7jf
Hpu+/qLUwUMt9TeKl+fGG5KPWJiRB9XKjYKt7E90yNkEQ0hHKx0Lxlqe8k3J
CwhMqFZcKQzMPhkmvS6+hXDa+cW9Q0uk97eBjihAIg9TGvGqmCvLc5QdL+t/
T9JlUYBFrJpRx3NaC7zELR9S7PgO5ddEUNunobf5/aF1oxjUj4PptdpmQG6e
6ZyBN2ElBIuNSriiP4kEOz3k0bEQFMQxBocB9M0RPmGAM+hN+GfpEVX+lZJT
q+P5fvVNKO8gtq9/H+KQ7dQLdSsnkrHbClP2Hn2pZfdoVhEHlueMhyvyRneY
lLWEeDvMYx8MZPtqTDHGsl6+W8A3+uUWUi5slNAznehRiMO21+gpWDpVOW2T
1p/P81yfGeEArWO/hE7qmrunpK74c5/8agalw5WGvJzVVKK5qLvh1Hn9vHVJ
JJMFrb2qp87TCohNbuGUkW4yjkPjUjtyLhlvGhGaaPcp0Japd30bmvtEaXjN
6VgeLXKRYugJk3eMF60r8TE0OoiRTcLWo8bvsIOL+qdOGkoHOxP2aJXzKMWj
sgS6pgIPlWjQhM8vT3//H1stbzhTlLNLh8qATGfpTYteMje5uIRDf/Y6WxOB
581UiPHWbSOLJIxB5+/LfHo/IZei4Ne3zs2gLqcu7xJAfzcQduTsX3J1zC/g
gYOB0n1VLvWm4PNP4Afjgkka/CoD+FUMGNq1gXYn7EaA8JzkD9qQOuegtOj+
QdthvHYSgMBlE8zt8JT2x0cHyWmw5AK/HldRN8TOpcLheJzn5NAvwDo0+Wpu
34WWEx1UtNllKyM4x4Jb13uqR0Hij8hbRKiVhXxIkjUVN7P22xPgsZY4ap4L
fYM+YM4JoSieh2rP6C+V+cA/SNToPme3QYAZgGkewdCJStEMNe6v7cn9dsWQ
xx+MuQ6OpjTA+WKMGSkHPsc0nYYIHBMmRA9OBBxFGk7lCxPDyWsknu5kjQ8A
h9S1FC8JC6wy0skZqPOPQ6qCUop8RA4HyXthJKi8GgJyaIn+aOMYC0ykG53q
dkuohjCb3wVOl01UCieh8FDoLhq2z59bK6CkAFElCyeg5vEX3vMi3qoO03kW
4NFwOkXDGUJHXMidONKNCxRZO5l3ulP87LXaoPipPm5uYrpRfMsF21lsaU9g
Qx4urnmtdiNqrbi2uD/vqZ9OdvTrKkuaXPn7LFf02Bj9I8vQVv3YZVM8zbL9
RTFWWdq1sxRzBbasnzWgj5gsy6Svw/nlhXqlPG6HFQlZxAmXPmMbbjGFz/UB
CmRTnDWI/wAXWaRNcJNZkA8ZNSMxT2kVsnuwH6UwLn6ou8gwL1GvFlBdtwsE
4O/1ftwz5eT3LVlOPPdtijxId1O8S3BYfhqO8r7QsbG8TW5srVSbIScTIv6j
JZ22+u2ewfGlFjRbjczauY+dtcJRfUKmjkA1VRYTAD/7hAdQLikHn+HvKy9R
jRouUPlodacDptX0KNU+tTA4QQFSDIsqa5m4+geTXF/ZkdH5QVGT8qhhTNpn
Xrwvv0EmxI2r8aPuPNYkQZMnznUzxORCgbUKskApuyQ57D/wU95/4rVbVH90
10ChWEpe01Rth9ULPdD0FIIaDxDL71LwtmYUf02MOr2CfZAFcLMq3Ku6WAhQ
krtI0S/MltbaUq3UhbNfd66TvfCSlWI8BS6tSGlVqADKChTPaM7RkWYhZCq1
gttvtzAYZ0uLnanrT2mCXccleGJr6E+qrYLRXOGANWJ2q2d1xbEOGdqBD9mI
UJRNAS0ANzskKvoHohoEWxIUW6ewrr6UJUaT430sJq4zDh9IL4yu4McAT4e1
YvzE+GnNswMphiv9aG3SGlRhsHU/EiApAzjYJm8PN6hEDFT3ZYceFmUf6Xc7
ggAJEe2VP4XrdgUUByqi3pZhN+PkSJLmZxTGCrL8qfSBm2hqyAt+cXkg+BXU
8N8oAFkGOlmoSTEQlji5pw+8ZOZ+gWgnFrXv47ztOzO77ktJwZAW7TuyVNdk
3MMaWqANBl7c2Nn9JHq0td+FnVd2chSuxBj3ttp6Ijy1MfYe8w7y2IS02aTK
qi9LJKlrTpUB0Fp+zBMEWEtu0qRfzfJRVPWI6yIzxVGxK1xkDZsMyhOeo1T0
Cu2Ycx9vwsVRg+dvElgK3nNLg7TqxxFyTdqUcTAiwowClmPX0B2ZJ8BprG4p
cEj+DI/BWnvPwuZ8fAiRFtvSFqk0Y29ZsekgxR803S9WCZWORLS95AiMecoo
5S6kZp75Z4+c4PLxCf5VM9sKPYyu4qbfix0LhDgdvPH5scuHxq597eCzK6wN
xCBKR3RnTODKZEkiobom1YjDdDIL9DOrEiQvOlwo8doQkUEY9TMq+ErJ0mjW
Cood/Tg5gIY7iTA6TGP+Eyrw4AycY0GyN0aN3CNuihIE0iUp26u0GfKefd4J
negED2PLH/9XmIcoEiBj17ZWTOQgMOAD+5db/Xvyro9kQ9sC5UM/TbpT7QAU
97YNN0vV0mjq0OdFQvGzMRidFSjZn4l/5PFZa30tRb/zPDqPxy8CaD2uacoP
Uu9GBDRxBlbrT1Lam3CXNPj4t4Hw13kzL6/mER2foDHiBkfXWowuxswOaaN2
OJbsVQG2pHdNsz76E2rr2AKWR8UhxBLo1lB1k00Andj7Aqc/LUI8nSxD6Sm4
/wHn+Bf5txBHqHdntzoSETyXFiymbRnnD+3qk9XtUPCz+jwKsAvevejEa5Hn
9Ms/MTBbT6T9RWXvJhfc8xNENJIzixrqH+JOrahAnaCtqJJuE1qtUoFgjLme
YAYo/9x9PoUsEaVTwz+xdg822xX0sG7eyFwW5BO+JcWr4SIuQWa+8Ccz+ffQ
5HbzONmA/NEHJpSv/WurEpuMRG5mh3ZIxON2VrUQGcFzf8e3GMjBZs5TG/77
zcSeQ81cYLE+sUyLws6iHs3Jr4quhUV1fap/y8G19DppB5GuMaV1LAaZ7Irh
6A9d3SHs213IpUujbNeiSHLjOFmnypdgj6D6bmiVy5VyApe8kesMbLv7Tfof
QbAPo4VTNzrrlHVHbuAWbjvyoI0CnleWmGwxkD151IRgLIqIRElm9weRpFqR
am+/EpcsM1iT0nqE4DZgKc0xGvMg9W9tZ31LIi16K/sbUfx2lF1EmjYjir8n
1VO6No1B/si+XK6eFXgT4ZcDlsahHYkrFczGqaMwkWB6lX+YvnNrkKC8+3s6
sfKmL8y1x8Xo90VdLAMMpCorfRsNrSmWeh7L4nINpMIrkGmJAn2WmGQRX+dU
SykvtweX6bLnZn94ISm4o35KY5xGok3bITVGHqBPXfnmastEEedwmN9/5O+q
fjFueoPnb6WTPZ4TFEj8rOPEVSn+PMJSAcVKcLvkRnFRLYuoDqL3a551emf/
PmRdwZILwPr6SYErYvgZKcnEV7C4YsNeqai94D2U3Hnojw007bav0UGstoso
U2KNsMFDcL1UlmDAeblP/4Og+ggTK+7LfrY4/3dRoWnH2+wxcna6zS+09kh2
+AfhIe3I28hjq/duZj5jM1OGAEf+EqvYDoD0b6qfRxDs720zIZoPzs9qi+Wb
FLx2ghvhrpNNPzktCbwoZZ1sEXkmP3OQCLzaviA1PQVSCK6j837lLHSdTzk0
+pKhSfXpw5gK/CxhWsIr/bRLPJOB7VXg3UNtLzoRwfFeswR0OvvRiE0Zs8JS
U0uXgnLofaOJMvz6mb82ynb++NjfobX+ktyKhemFCaBSCsug8D1KKQOHqlQy
RECcofFNgl7ZMrEjNStM1q2xDzeD8VLLfqJ0v2bC9tWT0KwGmMAkMTpfb3BG
sHIvus8yOZCNmVZALQSFYUnugJFPz7FKePllFlRenN4hcKI1muthSKYPfZkH
Y3wGOpvsf6fUCOcNYhmn+/lqiGH+9PFRECvkoqNAjgzSUmdXPvpq3iY6LSlw
BfnoLzChw7y9od7FLAtkbEKA6YCx8tUW63Jj6P5NATokKrHULQ1+WgbDPGuw
JOjk1UDo43eRQoVnG3RX5mRfeCzxzhsTM5qSjyl1/+fCf8Sd0ELm0g4kKABw
c18Sy2IIAL4ACJZBsDnH1JqMnZPBCmYK8J7eqPKVbMu4NbNj1uFKWCSlgR1W
EarycoLOi3JgRWNoH2bdbo3/zGa+yB2RdvfMjVh6Pw121MykjW4jCt9fpcmS
4u5eq3MbPQqP7IuiZJWkYZnBxPpwdHMhzSolzaOVnLS2Npo/4njOkGFkVQKb
Qek07APMbGnr1BX+KNQ+T+OTR9iJDgC2RgEQAx2vv2nTgsR9Bznlm0303osl
NKBSwgmtfa0DmeYX0odooDvWRhSsb/ip/f64ln7RZsLs2aA7+R5jpiwK9cig
rh4311raE2PDtAU5fZd5utdQ1fP8brBBp3p40U+NslHX0s9XKqy8+1m93FnA
Ir7teRTW+z/bQcRuTKZr5vY+Z0bmuWVnaDls9QEv9p2s21s0NW7p/+QpC9Gq
f85nXN2RXr8/nhnJcVFWQk65NzaYWWulhD2TcWtr+nbn3s2rgLYWkKhCgbHt
mFyOf5fB853b34K68akolTVnjjG2fvlQbbe0GKWvGeUX+/kCA8ILxfojd549
jLRkx3K93ZoIOlAq2uYW/cmqOWMgeQ0XjcNrXl1gXpTVFbRMRHf1UzqgwrFn
LQmww8pbzVvpQy5LJwxyYFjQuC6pT71nieSZIfH8dHbq14KG0BFr3mXG+CwP
SDNdSSORSg4fIgt2cqNP171TjFHYiH1YzWE8uKeBkvMtIb4Rwwz7jNQmHpqg
YGTuf2MqHZZ2eS1amBcHBLM+jZVjNJsolTuuSH8/ajLNHAKu4GtObbgoOIUR
yqtLLjiaHQSMSgX3gzxOVeziR7LYP+VoUQo2JCFHkxMcs0jjzawEXttAv4VU
/3Hl9loJoZYPeYNH/H/VnFY6ee8BA0OP1OiYqCizeTaorj0hfPicXZ8vYs9f
X9Fh+lXBiMwz4UzkrrGoBtc3W2lDBaDUljk2pRfw0OnJIhBvLW0usCofTulD
kIau/KNxDwstuEgqnPkaxESEVV9N5EPhkdkXlqmI+r2cVrv4bUrsQHKkKfkl
ovZZIMwPp7l4ofqQjKoz+OYcoYuu1cSLKbKjmD3yN22VFtwMnXr6dngZZE4X
0JqcZPV5itiTwOUDXY9m0dHP2Wfu19zUWpr7+H6KE/sI2KkjYuiBhAULb5gw
fQ1FYLmaYva0kFMLNzwdOxYtjO8CqlBhNaqUtfmVwQaPqPZIHHGvp5LzYhA/
sk9BhkZv30t+ieb946nfTcGeStkcIeiOJ3XFbWBcwTKk4EZj6jI1k/sO8/JX
MEXqhX9cKFmKgE0wqU3uRz5cIOPxPURuznEMrhyq3YSnE8o2MwNotXrKnOlT
rVv7kji2TiVtEPkoP/6QC3Cdc3KhOFKhkd7Q/6urfXoNGSFB6mIDeAbRxDST
vFGsg14oGTbz5Txn3IC0DKTPHTo61rq0QEER0yfrEd2iLFV8OaRvKKv/drxB
jJsr2u+0OOf60q3XAfij9GTiyZdtLev31yyH0EK0amThgZn5FSO+x2X5chbb
JYLqoD8NEQW4iKOLiyGKJoZ+BV5wuZl033S+tESGKVx5mdQXr3y1tG0c87pw
JaPIOKPDI3HjGwU6wHrt14uWuf8KHGlFeQrE3lzeAFvoFc9BjCqvZ6fGH7b4
nE/S5AgJJtspueLnby59GvV6R1vwA0aCBRl5wD4lNXYLqICxQKg26Bc8I86A
umlbLPL2qnQA1rPnTCIEhVM4mCmYWCWk1dyWh2WQikQx1UFJ2W0imX+2lewT
gxjDR0VI9yw+JqhKDKCpgpFMLW8cU3sRVUb5jSRXzHZycH3rotgNUjILLLP6
6Xlrkg6cOmQFJbfLOjnH6/+7PUoX44TC9jr/de+e1WJNJpOt7rQ06MKDyJCO
p4mW+0f+7GpJLxSweTU8XGZ2+ofHoG+yqmTc4xYuCkBfk/ghSCDwN06SgMgs
gyjYpdtDPu95YoqBaHm1Ae9UN7oaQ9ZRmRELDLoZ4WyafELKbtjDsidR6ifV
3rog4VIwfRYZ830ANz27hWBZLlhNCdovK7fQqdpoPPvg83p60oM64bZjHDTU
jN5oTVhVznA7d5lMWDl1RL14tyh/I0hvAPNNOEcMAW8q5PIjZv0k38Z6dUcN
weL0nuER+rWAWoJoGYSMlzJkWdTr2KMhZzcB0ELLu1va+bzQUkVB4X5+GaSe
M0jjWhGsDSb7aUyk4lOak1TiscvoUrYKdx5i3IAdieP/UlHUlYNRN9vBf/d8
eR7hgSJx74el6wEg3hJT5n5nNh+Jir08KBssK8TSoZMdYCZqSCI0CnisNIfw
EnClEnEnj9f+XYL0sohq1HHp7GSW+75sfWsjYR2E8jIAINfvuVIVgNxdW7s8
6lixfN0S4E/JpKlEAuBaeM1B4NFwcVSQDYbqQNKkvq3542hKg/pHpIuLc63H
zRrwFpuuvLfBPbbC3tqyOg+inJomAEZVttOYhSngGd5CWXxPQgvx0h9h2Ko5
8qRKZDGqTqXNxEhGrK06qkVGd/Rw+p1flcqb/wgV/C+W86JUAwdShh/HLNR2
gV8tl31hoVUA/gaA515+ExLm5xNUV+on+Hnl6m8LqRyLau3/n6mLNNdMZPJU
O2kzMWRoFFAH1bSHHxXf8jchflmeLSjyT0yhFitZE1gQGiqFgWcPy+20MoZQ
W56Gw0zc67ql7zYAHvzhnsfwFhkUGp7D1sJUtm9Syriu1TNA7NoN3ZGDCSuc
lVTT82kAibXwK6tm4gn1xMLS3Jl86RhvWQI6P/zGVK4JE/k9pu87T1DDH1E+
8QHU9SKnVVXD8fQGb+ZsO4b5MG/PVNCIIgMJEyg8xHJFE2Hqw/dwt1ZSzhvu
pVcJZrzK5/BrEhcW6qXC+aWH8leModXRtKGazqaCbtDIs8SJE5NGEe+rsL0/
Hg107WFPwgLSM2oPgpLYlUX+ToNeJkvM0MMFeTj9jgkK8Ovp/OG5Qzf5jxEw
fxWDeedf8zaCZ/cuhh+gXSZqLmHwlBoSTSOKrMoDBhDOuzLn4m2Tg0IhHXka
Bo/bfuGqlW6ZurFuGehPeniztV2xyfnDuIEIR4AQ6B/hxkCB1Q7c2bbz8rzH
tErBAo/JjBauYPAXsYmkz6+FqTv0YWnBoFO4p3xDCMEPKLA+tSpraW1ZU6JE
jJ9qpJ+IqJduF3QCUjDWTt2UWAjehx18yz5rLxmDff/6xy5/XoX29mD3N3A6
/uR/0djYQqzNMd1Cd5RA9xUkuQAWqN1faYEkXLv3UBRkmQNodbaWMyAgJxRd
bSoNXSw0UUFoPMG/HvO3RQXOAkqneOzOPzIuArkQBJl9cmNUtvSKE9vS6F4C
T+IlLRL0ackJ248w78p5pALAm4MMLIt1I9hZOrmTMe8xE9mlA4sRT5I9EcAp
XEfy2RfdLQe1DtrGy69tPb04Qb5zXHp4vXjrjPv8CvOYC0CE/TiJ3P99u0f6
S5KJ1GOV5ghSXYNGkhsMRl5qDpNdIcLEjFiwVvXE/Bichi2tZvOU+7zzsWA0
yW3d/p00vZNBT32G39nfq1MtyA+TX3/WR0o+hWhP3tZuA/sxFBnbxHwE1gZr
p+zkH5dWtyU25CPlH45Px/c4ddMduVnO3PD6kvYJNs45Msu6RosMpoky7LDt
QjvkX5ucXHKiFbppHCeiVkHq7Bt2m5mQaZqaSzgvIJE6eLkaEcezeNXS6JhC
navYPusaRKqIKSWfCv4UgMGX8R2Bj+kygR2yr4c4vNd92vrVm42UFbkcEvuH
om31tVS+ktJ0UzU+ariibZiOoOxs5LvuLE4JQv1baWrllmWFxS+eqtK1vgU8
iGKyNmcIxme4YkVATl2OVTDTXVO5ptS37Jm6/77Og7Q7wm3pdlmpeUvqBcdk
rZWD1hyuFmOVCcLUq1f5rS6oN34RS4EDu1V8o1tZX90ixPZ2SpVzWTTMSQz6
lRNU/k8a5xi6YdxCiWWTziOlZUfD1MDtAUOVIKXmcKu6jnbp/TzQGy6M7oju
7oOwwTACnz4mFJ/obIS8ZcjD2xdq80WEosjLQd+aaDEa2bcxUp/ML4B/fKbX
YZQjYQ9suD4ByNk0BeYwWHcsAkMqUamtnopx+ySMJDrRlFCs0341FPysNAZR
PebJz0msahZQWH6WArUHLL/MjTmhpmY2CqLospmDkWT9j3XNH+xME7yRlJF2
figZsm5CnMCzW6nnGtwvugKoAPubsUq4BIjkKhr/tm5mIkgoUH6A8xjRA2Ci
uTc3w3xVxo8crHGRLzm1HV7mllnWzDPGpadkjID49nn1j7YzAsDgliw0Tc66
HYi30PPc0W+RS4Bsfmi0SpgXmStcNt2TFvkLAGDPLG79cjqgGX/nJ2lA/XIs
yc9n56qcNRN62nG4uCbi6f4POqwQQond3DXTK02VkPg1yDNpM2ODjlLf8Af+
tFHy5lUV3Fhprhkf5n5WRINYFmOa1epoCT4BSWEBUGLycsac0wAKSnMj/dvA
yqgNG0WMMQ+rXnna2Pj69++KiNKXkms3XG4MwUEjunjoh02p2pRLUM7BqN6F
yC57kOpkgfweQW3ZU12mbFHmvuoFJxwYeVMymwzVJdO7+UlKubrb3dxDQeYA
StZEMW3J+7lMaqau9DsxAzQDz2yWsVPntkGsBoYQEyE7OT/iWpZ2jCymY0g2
gYhvH3uGOrIaGCKQiKx9PQUpm27ERDSfYXioNQeeReV6ZtCgTN5ooxguezk7
R345H0jm6k7DlvtSYS4YPnBOjNyU4FoSV6zBfPLcq6Lxr9MIAzrC8O66EHR3
8Gco/vXLA5b5P7JunyGQpIOZPWsnb1PErWYjZ17QHFrWcGtwtBldCsG+z10Z
LYHLRhoMl/znQwiy9J1kKBjOORC5DqOfTG4lGy0GejUZWxbesmOTqYQYjyvH
hgSxvKijOmJ9NgNkrCarRxjcNXJs1hab0WxRUwsNWTdZoOJXTgZEJlQw3R1U
OhZkkJb8I0ajlAWWMTL4Msv7zwKXLAlewrGdYJYo1mh9RH6RJ/agagJf+os6
GK0k+FF3UhPZRHysSc3enSpq73gQBKEnaz6TOotgRVtP4wrLITh4D4IMRtZh
mRN59UljGcgxj10tPhrDsq9qiuX1coKaAiRakoNNBRGLAYCTIX5JaH28qZU2
NzTTgSHQts78jFZkW2Io6en4xYzrn/uICLlFSYYrYN6jW0vNTlpF71npqk1r
e0T180+UfJZ+9dcUnDnCQQawwN7SZqstx1W1ykhpjab84d+fPM7PWqoY9VWy
qfshMMc5ncu5/QYky8so6vxk8HAbXENO4EtEnV8wLx5RXYmzexzLZLJaMHt+
84Rp3nEWvPx9MQP2IfXb159ws3yYZu/m4MkFNG0owt6Klx6b86Hr/z5R2U58
2XpxatY4AGVpLzwQ53Xcb/D9zvf6PkIAk5pUMerD3BVMi18gb2Mt4nBV/jvA
tVbZ6zMOTxdbqD/fS5s+2aDAR6puIYauxqHAS7Ax2P1rxsCNmg1jCEUoO2F0
eWzma2M5SXIqkyvCPWuLeJrmWTaQzWynS0tQ19sHd58yMG7dIM9367e9jrHO
/70EL7W7T2MGnixR97P6HAZ0uHT4UfPi9w3q7Ph245598BwxUBwLicZ0Zc8b
lAPLnovYs/4gJgQHPLCULgI3HdSfAGeVOk+HXp90maewalmQ1KMGg4j0eb/I
yUexIp2kw6Jk+kBsbjmzvZqDnGNBEbuPjL3IaYQBDYrdrilUCp2FGxl1dkf3
Q1mH/Suf5KgySXa6mqfrLH3XukHOSaDb+pXafdO64CDhhon5YrQvb8B3wJvw
ljKovGtWAUZI7XNSvbShcStigdASztttgeQ+bkRKFmcW9FNye/TfW9PWqoi3
kSxTMSdts9m+7lSBhm6hDraIIjcPaYF7HPIgY55wo6Z1qYyNb5C3jnOHhbAC
KTcXNJeUXf8CYrdxcQWA7yjKY65wvYB8URj9wr8rMLNKXXsvgDwQ+QdDi30P
AATNVITS1jCUj6Ar09owd8vX9Qo2HmzRZUSndnW6+y2UL6JHXq6jSAveyB7J
F7wBvoPYw2KsjHb37UjQnaRzvuANYdAhJbjihW2qHmqI2lYmGaEWq4YTP+rz
zmCf6tYqVW/rT5tZXw0hOTpw7k7Q9sHDLMvct2qDs849FnBepuw8s8Z6mu1d
s/4R73eS71FYdtPhCJB2XIiScG7LjLoyPJALofkajh7eSpyBFWFHnntTe28s
7SVnQehyyNwiLCFhK2rCPBjJC+AJa5/tBY4jFVgxx5gQO4q+OARdaUop7nju
f08kURX90ESP+5JkdoVCVFJ3wy6K/d03Dk3plQgO0NMdYhE/bv/WexP/+iTA
B5CcElzmfe01FYc4zxttsCycoc6aRvXeyRnbsmLDSSJSR7DGGnReABhF2XmR
RkBWJkBJQQReLMBg1iRzqpOMm+wFqCyRkeSH40VE/DVHo2DByKUCAfQLN+T4
42pSaDHJC1RZBe/Z6xbrLTBk2wvgybhUktS1JZ3bDl4viXfMtUZKxks+aHEb
2/h4Y90mA1JyzCuhxSdofZGngP6UMW24w6Rx6HWJR+B0DkI59tHf1b+Nzja0
ImdQcwngc9LtjzLVYrP/4QXzyFXK/dJFNZ7jJeTWfvMEqpF4crdcRtG6TkLu
IjrBDJZ2Ivm66waGVysBz04rUR4rRwomAQDBV227Cp6BGLwL4PkdNAL6tDCo
BHTz9CzY5ZJUGyoz6JOyw1WQuSY8WLkY8rr8oMDTe4GrjIfFCp8t9fgz2wmQ
Yhx68GnNBPTXoCUo2AlnU2xAgRsp9JefIv1MBc/7M+4gj6vpcjhFSrx3LmMw
3txewdewkSFbqsp56qMrRyfTMMaOYitg48rPduIFqju1ZsgOpETYss0BkSIW
XZ2kz6/EM4vv7JLtOlU08DGQqccRG3dhw82yD1uyaezy8sBbfevrIIrUB1dm
Wo2yOE2OG7kxUPvJxQGvdwB2Z+ErdmKowyB3MOWR77QLfNelEXkfsKbe3+kn
tDqJekyZ6id46+YS9/LybkEOcFmUdNe3An8KHHTPbNfexAXM6pUR8WXp9ewx
i+Im0TbJaHgHXC9PKYyVFURVG2FuD/K6L0z/IyCVQk205oMpzi9gNjI8h49u
YJhsDWP6MbDFLOyB3kG6G0UQPgyuy6S7rEbA0VGdMGrmIZkZkjGLsRcYHBuW
iYlRZe8tQhawkfxRZUkI+gjWy6XhRvwNnK+mC+S8NS3y/LTVKtoEEJwD6/ID
+yh/Pknw9gPvIjXMKAVIqGBgvx2pijHSVCe1CpE6A6aE90UPvDP4GzqtvDyO
8oFubtHqtG28Gg66TYgVexTMfR8C4UI7eS65h8QvOg4RcaURzRc8pkQlxvMi
CY7yF0t6x7mrC6Pcey7nXeeC1G+GPidMpay58REaaR3ltHKme726+zyrLHvd
TkKAVhLcbQia7ucvZqoEAFewYceB50mnIruwq3mC5Km+uSjqZNtduNJ+O4EE
6soDRd/0UnJn74DQp3qStIkWSoKcILSzHLVDdWNt4ksmCnYtipuhyS3lNUuX
jEcWvCyIdJtgTqabpEEVIaYWcSJTwaFY2LB5M1868WrDug8K96XsHIl1f/Z9
hl9GU5thG4NH5zY6f7DKH6HcFhgPI5QwHesoqeUwo4yy7qONJdvyhIAX9PJj
fgz36AVxI+q57Ij1l2UxIvVp/6CtSw9Im9olXwcWfTtJxgxFWwtBkF+iI4cX
b0y5VybUU/auRjKN4Kp8hI458/UIYm9YhWEuKWeD8kZ1lP7/+6o9FabZmUfY
Bbt2OAcS8LoBP424fa2SMuWFscpTMkoxTWvNkjWWgRzPTNceDhn0DwTNuTah
8L5OljLj/nZDcUJrkHZVPfyzjXVsxf9+Uf6WieceycH+WdjKxwV4yU/JUr7G
3OMu8KZGSkXJwqcAOQjZxDTTfZvKb3ouxQGJ2NPJ0whn460ybYYKyXva/ES0
q4AO246JjrXw/DAc3vkCY/npaxBo3rVGeROzT78TGJIxegSOL0Si1g0bGmkK
Lae+IFFlMECsRgN9/cDlBZ16Yykk3LAq46hcuzUzw55FxQV772cVC05cezt0
kt/bB5z9UNkBerggNTzJIVM69m6tKSEl2k5VhyK5qA83z3NFCFni3ImaojbG
yeDoegmv75GthVQyrqaZaoF5d5lZRv/tun2PhNb256jXMf+pN3jtGu2D9ah8
f1X3pm17m2uTLJVncWNeZ+cWCYNoFanPvJj+/ymEcr79O55Ir/hu1O3f3qvq
+ma6Lhz/P/QbQy4Ztpsb5MJpI8zonI070PSfFvjdmGUMuJ8RBJ8RzirBf55y
0oHsKYZlDc1qpKli6tp70CwFo/Zfg3hfYTCXcJ9W6t1n+N0+MF65dEG9rRn9
5J4xm5kR7gDDG4zKsZj97ydgNcLcZwvJPEKcnny0KrVEXuP6sILlFe8E5Pt9
8ljpTTw6u96oqN7Zq0WYEIiLUxLqfJp9JJGSX6mWfsdVx1ItOZRnq1caKF+L
bvO9KXX1WH9r+JA/cZVdItVG5JMJuxlKShyKBR4wIsqNC8E2Du6HOE5H645k
UyPDaNDrdTDwIHeB+lQFMb4t/1mNgyltQKNWXsqH32wTPvRYgANcsuSMLEIx
Ro7cu98Fv3GLYLTvN+WWtvEirDIRxABNrhYqb9tagfUSZioFrNN/T03X5dd1
DCiI/Y+RTvvP9QtigAi4qVLAZhGZRut0GyEhv3SMTLmcJu92YfNYHCuCB858
G4NUx2dOnYjA67XxDGljZHoKmDQ/uhawv7Ad1VubHpxaM3suwx/50/jHBYJR
9dzHvZisuldg/jJZ0h+NzHn++WeFdrcETq5LmldUPtsF1DDNM/pzohx95kfv
HWU5s05BqDZwuaumDxDkxGyqBj4qPaII2pNINAShTT0/71izRwgfiQkyqtnC
Sh967jw8KGs2aYeDPP6q0xGd3+9yet8GSRjIABQS4Vhlk2R9C7QhHHfVO1TV
rBzRoEn/6FsUwIjNcJl0Mzebqx2Pl9XSNuj8jZEw6qLat3GK/QyNOur4cMhF
Y3RBF++a7KKypRwADY1N0GQ2nHrT2Huk6OvtXDUEDO8TBJMiM+Y899EI+QBu
ATKBey/8bt5zN4udNcQgvRarbS7jWaCyjggbeQkgbC3BsNnGyLZ+xu1HbTZv
8Gf73zE3Ki+BnHKSEZ0cUCEiOuu1fpPIevdmp9I4W+kDv9Z33VOA1Pm0qh+R
A5LxHV7mVu9tQk7VJyORqQqok74VybtHp2chaMPB17jyDdRQ0CqATgFrL1WU
mfkZQ0KoQ94g3iFceuQxK1xG4sKgFpDh1qdcsDIm+G7odTRJy3taDM6lMgn2
UNdkERjeU1tE1CBlQge0OVbOg7n3S8+bh87h144909I1dubiiXGTWZzbNMlD
rfnRXdKm7yORkV7+t1AeGQ5u/gsAcwQmmcdn8n+2lXOeAJRfkgrMnHdcuv4U
ldfWIzHSIkE5DeMq13PO0ZBbxITqHD3CjsyuK3Z4n9Kh6vvqUHsCMM/SZKk+
ALN40abj6qkwjcSfwm74bbHGKmxb8AH9FTWmKNfjU73U68Xtq1qpGTYNQCfI
+dSUuu5pRSRKEiQGc9GsG6qwd8MLyuyWnXGYGWrIatgH78iolZ0bGnp8kEpI
rJGszZreE6nkN9xFhClQIHrrEe/GD1Qwd+K/GFOlybIzYTQwrrvI7+akD4tD
Wxf5+l/16XLk58qs6uDM6692j6RYguE5r1Qb23seXtJgLlK+32ZIj3FzCpTO
7hStGysLLx64vnDxf43IW0bLax7Varg964vDqmeteUUq7hmBVxN+lwS/PKyl
e/0Ta1NbkJplfTEuoLTNZzxQma1k8+blsBbcTALOAGsNcWus14hTZVaOvlxp
TtdcWSNZC5nXUPDetXCQA/fkSdFSGc7WfYHCVaI97zett8UqPZjbFSS//RbB
ACnhSs7kDU5rpsYaMq+1tsNSRD+O9PGTuC/iYAOBfdM6mO8d8lf599W6zmi3
+mcbn5gXqgvvkS2j80gkVrTtDEj/6jrKefNYCOJeIcc0FRkefNJWLcVfbJfv
m/3ZLbkMBmpF4MxNIohgMelGrU8mRPquJTCCFeID8mFRIaph1gRXHoKeLlR7
FkIa3lI7gF+2o/BpRM9rBknsOm5QIPVEw2O2gqZwzErxgPdrKEwOTUXxnyAq
cpb75EDoYnoY6PHBKzNH4Y3KjyNmtMmuXKQwfuSYmrM7lkyOEBa1r1LWXUOD
oHWdN14kckciCfxiRkEhhaZOzn1RRB5QxM3mcebNo3iM/S+BQBaFtVEnYnUE
tbLusbJ3qCskUF18og8NpFla/e15dpa6gtLx/cnFPzOEMB/M1SZ+TkOVoue0
7ENsaO3/cLT/yzroX2g5PhMUP56G6UVy1s5N4TteCkyWvQ+gXvtOcih9Qr0r
EEAPNOAqWwZv0rG6aHoHb/cWAy4oaviKv4lkK45n8RfI2m6xwkbkwzahCymH
VKXcdQ5mfTT8VMcbyADq/6ZzGScKlOtLNvjdb73GF8V74c32Q7poU8Avwa9H
Q7qWsc9PHHVlDejcvuC+gaJN24ERU8JlFp3y97zH6pp+Ueg+ssMiQk701a6b
MgLMBEwJWyP09W2V4ir1f/+DF7GTsKvIthPYLDmXQ+utKzOc2CARqLXn9Ecj
ga56gG4/g5igUEIDZrm90z7mFZfy0OZPKyPr8PGTVyGR8zHFY/CXwGq9OGb9
icvVWwo6TYPfsgGHpQh919HynNtc1vXbs8s1HqVSJQAvqphLKzS0ZqZI5ing
p4JPNsI7K2tP2xrwI1LR7702zR447UoxlilQZSZTf2pzaE+9oOsdk0etM143
7M2Xleiam86qB26C6cDa9D56TO7dCd7Yf6izykEN+t9XHywrJH5IWrBnnw6H
HLbt1RhLG65n9cLT5Pw0Q0CaEFqEECACluLyG4bqQbHG9CPjSD45Kd5n23t7
aR67LfP2HpmSD/YBwozVl3+tvGeIPV76iTNxGpBdB0wohwhZCK1nmWqyoWOb
jTqnhehKzSLBM7XU4PGnc0RARAJw+zEMarLzYIVA3zC2w5TA8WGCGu1c2K2A
0WVxB6zlX3a4wuJPkmklPG8uCV7Z/HzNG6YB7zBBrirg3Jz0OELD6tHySbU7
gC2Er0dmEe58/Zm3iMqDHoMXM460w9iE7Di8GtnCQhCnuH1UxiYKZlMpSVUD
dm8cD7yCexrTsr7kKgS74qCT37tmk7hDfx62j7Kidb9QshVxoPCwYdeqKjPh
hD9ZqZLxw1d0pCNZaNSVprgCkJfQDC9Bm4m1tCrAPcMoo7Nr/KIp9RLCsXdw
NduM68H1KDIRs0MyutpWAhT4xNXhkXkuWfg8owgPBMKr7CVGqIjYzsUELdGp
TeFs70iFI+oB6Pt8DRGq4MzyhD2XbLMCK3wfDybGmHsv3JFykBc5+mbj1tj3
+wDehVfalYNsatphKv67gkv88HNFlO6PbRTd3wI9Ps85tFTTKluCq6ZoxdOw
xNzcjtYv6ob6+J8Rjtxb8G+d+LRrt2SUtyGhMlINg90l3qNAyx8/LEab5wmC
iTa6RmxcyNHPoSOpfevukDU1CZFHCCfQXSpQwK3IWWOikn6obswvemksIp3R
L80KyiC6rk85p2mtqpJ1A+jWgCD4EQb2rhiGF+OExrHT0ZoZFMpmmr4n+imQ
KJ5KcL/XQiEWG9AesSx4YfceU3/VlRsxptspfyj15e1oUduvACttjkfHTzdg
ViBh9jnSVPvka3HSIH5Vy2CxvikqEm+deRyt3K5e5ScszgTdNHRYhCg0v0aU
JvggnZol/cE15sQE3/rFPGg6ia40nzvp1wxQJXH4LoGRfSYxqD3J9dlghb7b
awfg4GrGlYtZ8O20WmN04u/9vcgRpVkDIc8FEZ79VybCPN2qaZDUXogGQpk/
xYZWKSyq+BSsWQq9MojzeurouHV3Xae0Fx3BlmramMB6WPeAkUo5cFjM4UcR
rzozDj/R9YYmuJlxAaTsI/AX0ztd+lWuat4ZUCK1ltAEZtXW3herhCqMNYq8
3pwkkOKjz/2NtGwDI01jb/JZuyVfejbBXwzIwKU1tVx0H8TiBLAAimzH/Yhc
A5osCjw5g6AY9cVCEp9MaAg5BrAj/UBK4SEEQX3vxfoNKntuDDFOiyAJCuHN
SzYEkOYsVID9lwNxIV6KraZjbvUOonSrF5Yp9kDLbwjD580DEuuoO4nn1lql
ZI8+5nFP+OqYwlbvYtnhCLMWsk14bmMPwu/wKy0+FaucXHRDd1SXhe1HgV1Q
VH0qQOpoGoCkc4/1SRTWLLUdWI0Y4tU4I/rS/Em7+TeHbHOR20fqHlo4rcA+
A4mP124X2qHKiROvuN+K1BhToqnD2A/ogvHnKvGu4PMwfl29YfGzLEvOpOmJ
HK1kOXtNmlV6tdaDwF1dI0dSNNq2+MZT1+doEOFYYQVYfR+BeY4X07SK8fMh
VJKjVQN2dmRyhFsFBEuY2JMGS9zKizueRZPtoXzNL1KbeZqIrpfcwMjkP96B
zeQ6LLAWGJ8bYx6wxiWyl5c0DkFi5rrpRxr6QKNi5nS02/LF98uj41xK5RZN
C8IcRVuUGccS6pF+Ok4+KsGtl7CRRKpH47fUQd4qbf8BhDxzS22kaga4a06p
c2alpvlgv3B5ji3QjQsVwIXk4CKjlK2fRPXJ+URxcNEfj7ohZWQl2/Y28j5R
NCdct7keyz/cUj4U06r2pMboKGhQjKvLy/i0HU8rZhO9d1dFuTW3EHMpgy71
pHb4XTkKfVbEq4YuwKUydUIqbfCVodon7XFe51iYFuSzkTSMG/AdDUblFlcP
VeNeFM3EO7KvI803teMYhtkwBuSOv9mJLtH7oFW6J1LYEnyJFqu67SSmcy23
ua5qlY1uFh+qNKoLm7RC3CZKcSw5JXwyn3fTIKCVFXJt4JCK9CNtlk6Py9vZ
I3byevcgDfB25lexDeB5mkh30OstaTbtrzlGbf9EEUw9IVIF0FbUJy8rwGmD
BAqWLQfnLgRaH2359DIQafvGBIjYyQVWCJ8wraarxK/MJBSTbt0ueif0XVyK
fNy385akQ1Mh1sEz0aWypItGXyeOXgXoKozdiU1EOFaDWcOMHJa2DNz8iGkg
YM0Z/99YhkzAij7lMxdmL2zTo5h5cuE+pgV3fIoweN+BPR4TkTVLmoZVPFHn
tkkaChhIsSzvq/xLw+If7p/P1iSaEm/Pjkve5VKuyHoiMwLwlc2yHy5QF2fH
ZmWoAHwckXDSnpjXzKn9Fk+dJfhXzZgjwYUvT6ZyV8RxWAaeOmA8RaVm/rMq
x8stqbLaJYR/b5i0aYISmXYuSIs2WYc/hVv/KRbxtMIzHfgRGGQ6l1IMLv+u
IZ5w14ixO7nBvWkSugoiLCXd99A4nYVpwYrfPzcCtkv4v5TCp2U3R5P7njkc
wUxLW+I2Ufq7ODNQ0VLXTikgt2us5GQuHiqbzckk1sBaouVvL1u1X8RnItxw
T2cZpTacZrOosTSpEGJ8TyBq14e1vxxa45SpdzOzS8mBD5MD1cFekMrrtp2p
A6QOt9+Cc3NhKFgeEzAVTDtIIIbb8J7We8l07vqb/RqCrZWMTQpHOjIvltwB
Kf7d1g5E+bVmgT5+IyyPe3aik5TmnNR8tWgckGWl8jJkTIj//Q3VVKjX1/Tl
+v8w/2I6BgPQ3k2PHmCSbHM7FGPQ8dqDHbizDZ9m7+xM+1plkkY1GqPXtkK5
CC4GUYxm86NFxvs1DgoxeIVrg8y4FJpj9VwSogRArzNacrJd30Yo9wGQsbZx
ByPEG/YKpeJrXKt1srCk2IG1w/7W8UHnqC9A1qfeuTa0R/WjvbPrnRZxmEWw
ysEh+SYkbih5fTJbTO3ySKoa1gyP0aKuuI7bFMv7qm6eN8vpx4I30uw7cYeu
NnmJvnAIG7fk0MNlB0n+/vHbrvIyR5K144rWcv2bmUk/XX56ITd5hAiwFOLd
GfKN31wRQsR2ycyzqVHFJFsoceCqP4cKmqTE45pc9DttPmvgQvopDQ5qDYTJ
l+qa1cKf+TeWoM3hHOUf6dZV5VkuWOSRYI57zft8OAvcSDE5TPuQJbrJ3Udt
hG3CR4VowY0XwF218LEz84EZS5g03RO6brr2hCpKr/XmGOHKlt2MbIHDkHtw
Yqz2T2dmyk5hgGP4NM6zETEqF3MJSXk3D/efNjPAWs7+cJCW9Kc7Y5jldWsf
OTLqzi6r9/nwj++2mTDazgHTDR104jg02+jSI+lvTRJcIbvhLGvG5onYmYwr
HNaVlYhDUJVBJ2EgEmXFelaOEvy3AIGeDJ+HSmBtf3ab6S4NeyJ+fKzJG9wa
LWMGta53ukS0gPlCctgSkanpW6dMTAoH3tPjLz/OYlG0T/fwLm33Z8GpMhMi
zhKEXiMT/wXQDEjqtIFMayKP2iTZSBrvUiJbMJMbAV73e2UV2kyYv2zp+vIQ
vX+BYormNOT1e6Llzn+yZos7Y/rEpk9du1Bx1fHKwAM7LkEXhVYVmWJaesmC
KV3EsUnmKBixv0TXRo3PTg+ioPG8gJSvlurMI616b7tLFKbBQ/xciuh/0SWa
JdpOFqclmpFvmGNEg4Wjw+o5MYL1sHjKz335QSvA7hf/qnZ+bFnci8T+bPIU
gy5qCy2NJTWQERj7KcV+a37vvGFL1o5tRFJTAlIMKXBNeP9Sc4gZ9RKoQ4p5
tYUAyrN1/0NHfEjf0Cz6nezplalSHr2XofZDG3e2V4ZaLzohe0G+RLKhUCGj
dqCPRCaqlqsR+/KMOHmk16rieNdarUoWJ97Hp4BM6OQ7g+CNCxgmrAGTNBTI
vyq/SHSMC4RAGcOnkN25pNxM7yCMgEE68fF/y6ow0qMRKHLJCuEjd8UhYWDv
PX0gCLvJDzHvn36Lt9jEu9ipJ4c/f80nJasjGTXoktsyqC8206Z4BJgFrg/2
CN1MQtsrlCGutQoE/Nl91PbdvhaphRyFkKnjp1s6wrpeUB8Z2Ay2afUJ0Ss3
7896nInXojE09t00MOboteJoqxFFECklyIP4NhKaGqUUXHet7uR9dfdaMX6i
cAiGgqsdK4qCsHxpYtzBTUe0Sft8FsT1UN1rhY6Wy+6Q1pxGmxM9Xa2SSs4l
avv6xP7oChOmzD6lk4zYA/SRPJb2treBnntykafk3mCNXAcDtYptN54PI9nQ
lEXgeVTupWEyf3yEtLqU1OxhBZsrNpXP6oUacPDi0OVf5lA7en7Xo2uzTi8U
eKdmU4ys4dBw/rA6L/ny1D8/Zv8oJwX4YZnMP26xHQTlO1QGs4FIymagL/1P
rrGA2DWJEm/Nto+ao4J3Mo0M6IDFxcTBOoXcumEnmXNIhEKHDXGKbw0JXrw9
JrMaL5z+6MEN+oVtfKKl1x4RntAlQbr+19MGWXbtSr4euKP0lRGG0fdifT57
pO5AHDuKijt/Xr1r0FyaWCfjBlo2EYvTwDM9dyiwFum8l6sRgED4p1WAoN3w
BHMJRggfxa+b0MOKWVLoOloyTjAyx6HovaZuxhqkBD0xzJuUhXrpcqb0xjkf
H6c+JSsSCGHlCBlVYAr7q+1FFLSfl/+HdpFtxYm/RZwdVxhO9C3HMFwJbKfr
WqfDhf/2/9GHszmSmHROkT/1pcw8ToyNje+2d5ffLhn3jmkha+18536fgChN
HtZze39OQnun0rLolvKQG0pQWbJU66AqrokMwjnmHqVENamus4DlVGX+4FTY
ZyieJQgOU/RMjk7+mLOYC12VzCPva2T5jqoexwe36i07JhELIVTYjhmDEVzV
Nv8SgThqJM9Qjxb0f13WFbAtk1cvkmT3vhWzdxXrTCLWjiPEuV4tRKdd8vh2
WaXueGAgdxIiQ39X8hXrUnlWNjOt5/MsVFn3bv7wNiPXDL1hpg4/SykPobOZ
VWuDNpv8Zn97XgNuaANV3eqHlCjjK2K49HE+HfN62tgYP1Qm+k8clUGJbQsa
XlEYP4LcjTc26I4No5B5c2eGWo7Jyv8txVE3Pm9CFmPegQP6c1blJ999wsAh
rDJ4Ow25akQLbVcRO/9ixe8N1qSbrtS5xC2cRQZhGlC9+Xl4SDaBR07ZHHVB
UWUZrKM4yCczFNXHPje1n/8WaNRa92vXvV4T8LvQBBxnZ55sGrIrWV5LtocK
hydlpa/YmDoRJ06cTR8eAsF7miNslkPBRs93i++oXCqnBlC4s7VamAAZUjdx
YXwIABvjUuNPVdK9H/2grlvofFiouOFltubp4C73SENHQkTqVsnWNeIYo6BD
pMNdP6LZkJyYDAadiTyt3kHv1fQIBjUfzcKwdoi2WVLrWBxHZDEt1yi3XJ9H
ZsalB8h84ciugG9osbStDV4cX+fIbmdNHcn/CwdqXFQTAAMrJ6391Z24iiqw
cizK8FF7ccca2nU34kwIuvjEwWIPWivfpdRmleycwcsWi87R89JKv/knrVO8
b0EfTegO427UrnCTmweA3Bu7maE2otP6UkUiT3F+lEuccRtStMslOxbByN/V
zgzwC/vrAUeS8xSfOc9VePvbUqzxWVURObpaYtG7Ffri8c6hMbRID+aTx3KL
IPfKzkdwzS27D7PYsT7Bb98XrdTmDebtIC3ce6bjqpv9mRRZD5qh2ObnMlJs
CjxELe35EOqXYZyjbccM6vbKTpv4gHa90fIUZULOwodP6k9roRpjpWCPojX+
UYRb2EFePshP1VOensA97R3FcSeHFGM6d97cLGrxzTsQyjfuIuTbldZiLCxP
55XuFeXR5Bg1h/CQkTrUf78mWqJ1OP/Mtd7Jg8pYF3KeFxE/0hGQ5tfT4a94
+rdBTHHDxLcQ64Vcal02KQTTrTwkWxXu6mZK/Nh5FJzSPa08Rk1hL5DXWXXp
nbMSDOaYqyyHwtg+fnuM7sVWxxANsJBm2jru+As8OMrAKibZzQzcPibNG+QN
/XGrdqhbI4ct881LmhT8epCXQhsWO+1NDK/7gg9L6pL906kcvVqk7+tk4LNh
k9JDykCdUFs/OSvpgotOwUSJiJ/FGoa0Zu5r5QtN00XBIHXyHHloGGXEtkTx
JxJvT6tzsoCdhnEH1RcxtM6TEjSDR2/Fo5Wfxdff1GulN400eg3J5po//ygZ
W7K8R8bc/gztaxTyFxlQj0dc4mtagWFrJLPfJLQbTxkTNjXlawSUU3dsLEXl
0X7j3wiMMEXv2rrTBjY4gtjrrozKOfGodR9f2Q0ebQuxxx27CnxS4Tc11TTm
8IUgnAdk2ZyZf3eqJ8DToOlOX8dt6hHdoApLyBcc+cCIwTv8V8p/Pg1ZjyZt
E0OMI7OERbZKrkLKxapcJNCEiVprtzplwzVHFiw6qEyFR8cUQvJeufY0YnaC
p/rq4RtSJVQP1eDBy7F8Iw1O4iJbrtzmRPa/sNLV2kV2LCVkfyNmVlwJWev5
ih+H1yFBv9HJ23FD+x5+AHCzDSrfkcQXq6u3uJ7s9cglGmAcUN9t6SiPm9dO
OFtS6Zuh82TiU1wPd4hnWqLK/1QrGFGY31BGRgTioW9EQbC/K25+k1ZubEbd
txouYAC9/xTP+aVv4vgtwAvzpVY1olLkzjOnC0r7ItmahkEcbawQWXAAsuGE
kd+J08t6oX2wSwvsw1T+bxt52HeSdSV9+n707T2PgXDITqYhuQ25jM6OGVlT
DukSDiEZHZe1Trs64khV1oDc1zx1PUjdqYYYXyGXna+asW8EwLYcIxVJecy9
RWNtNHG+5V5g0fnWt7toubVQEzbEBJiDcneEJIDxq+StJv7/UqFPRi4Flp22
GG7HyqF+zmsNtQaXGGO75KoJCK73F7UtgZvODU2IvMGvRUH9+aK5mh+s0Bit
RX4yp7+uPT5FgwfAM+L0VObVgObrp1uF5IV1yqHFG4EisDYJOUJWNF16nC3T
N+1sK6LnkiZnVhpSRjHRrnedxYJLZKVT37W7M2HRn26fNHV/plLgY5HSe7jg
kzn6Lmeq/RNOaykW5xtsmgQHHzRakGywT9IULlVe+U178bcgkuO6XMb7dUGb
uxZOJyzm/DG4+ZBF9/QYFROKrS+KIdvePbj9Q/ICwcjXA5z5mdfYcvcfaDpd
K5v9btvAhE0uQe0o+yMG3JQwCWUS0B4Px/HaDVu9WDUxOTbUJNTjZsiLOyV9
TiUrah3YRrzKDNYt1IkThvygKfjr955uLXI2SCW4RqNzP4Xv+1EyHWa2Gl72
McQhWdNh35C20KiM96gelQRFduKq0eZ30aPLZ3g7qPYhxZgyfU0iYMus1I2p
wFZwNEYWQimhE736j59EqC/kLxd+U6Jg4XqAgLjjsPMDm4N1AODQadkawBKB
j2ADn9tyAwf6c/Vn908HPRrwIq6J3CneMAbkS0gSNDNtH3zmOXbaluqf6sAh
EWIRvxvEK+rjsKKZjIL7jv7TiClvvTYf9QkeJRpFcl5u4AufOxutFx/BzFZm
YMKENmvMhFfNA9A1s8tFB8MtU5dHe00u1bhoyRMEs2rOeltSOvbXQNkvhbMj
g2lbvoG5fOTg4O+EYT3A+yet3uvv56Am5LqypoPKocLpu4chTRhx5Jc5cI4Q
ViHi6/ZCkdmuDyqikm6WO+6FQqIKpsfuc/GOFhgeCw5AJvGK5VG9MxUyAHeT
3o7aS3hRIjow0PQ4K2KZGYz0czy9kYl0uN3BwOZ52/sAT3jYt7qj6Z3+9/+P
lVoG52B8Cwq8TB5gvpLAkYPYjYGbybj8zHjKYxmgTRFEyGGPQBt4x8TJ2Bhy
VyzWMlEvXkJ1gUt7EmnQ1JNWGQEJ/PC7QgkVhJymX750PhpImq45936Q8x5Y
+EhD6qMSUrcH58sT8riLFRT35He87wPFnGfN1drHv3K2j01Xb0gEyRM2xGsh
oR9n8SeYhQ8MD5wWj89R8cbNcphJZoaME7gebJfyIUTo2dhzfVXPY3nQ5V+F
h52cLSglxb4oldXfQp37JnJ6OodfazXQrXkIg/AQUvNWvfrmx7flnQkPElf5
zbOGkYVUccHMKNZAu5/bBTxGMSqQdjxEYzW67PZQbrBpOHQU2t4vRYsB7kj0
qfQvZXYBpCMVXB1v0i3YFloa0paQJ8TgeXs/5kYHUHRzNcMjtx7fR4A+RYov
nyqqgW01kHEzlQQ6jnVYEJaj4YeXrIZvGK0rrDMIYLOM8m8Dt+l+RRMsU1bh
TENKVK/2CVCPAHTmm7D8cw1tfC/1l33RaUYZ47qZHA+Md8tJZILBCZWGzthz
SJ62iAX98AvnhEeyakX39ABySfCmi+g+vsFa6jbrvRligtVOPo8UgD6Gwz90
6CUvewTRHj7JBkr2JT8gxZZy1/jbjGI2Bcs1QH+1Mz64BSm5MlOoCkUq6jEd
ZIBnq09Kdhp/RTd6/g3+eFqkG854LMLUkVGvCmtR90UP+tud8l9BpDG2Qtl9
Jft+InZmEs9PMIGypPq58jxkmTNypCXFPVqxfwN21KgAkDGmcyFACk1qdCVr
hTaCAzBaQtd99iQEuPhBNd55iftiTV6wVuutE8UWc9EdFPdBX43ArIXL7TRd
16K7KVczcGgY1383Z4Z7oWitxN1U8944UANA+mNmxaG6RN854jSv8mo74qhj
V0Z2h23qoG/UNbAjwR0mlqBSAnhcNmQJ8mpfHYlfcCAT3ydhNdLYKh/qAe13
JYlGMBIkvK031cQLzYPkLY9RBfHEikQ2PqdJZKyRXWI/ZwEdyecNctUhhKBk
YBAwm55QIF+/18uhYTviRMzio4eFjB1HKysKDapFYManvXfTK0i5AGt1I7H+
eZQ/zZulbr76VzY+exeSuaYRNjCjmZ0PDVC9JCa71jalKYhr22UHmguDi5oc
QCNY2hnn7GKdRAqWVPGe7lHsp240jtBA2gSKE/AzX1/qPSjyoKDo1OwqC4zv
+xrDpGGxcrQrXXY5JolxjMZ+YrH5JQMzr8zqe3VWOWmpPgKk7/iY3AVN3Upm
o3ogqu+0V5iIpV32M1oYiiFkdldXvDJln5rUViPLq7Y0PA0T0DYewMRg/lP9
f9xmAsIFY+uBd/xPnM/AJAGVfp92dfgOWmwByJjvbKhQnzOd2Dmg6KILf8xY
VwM/XGi7pJMN7xao3qCklPLg8mTaXSIK8+vBuCrxFZDQajTwYDO2ADZdzBwN
eoI6rtLkCS+5BC5PFgt9iHX9FF/VCO2/1gXSJLobWceFk7kWVeFfzAKEtEAS
zlrsLk2SEGuqvQzpoQ7Bf7pa7EP/8XjV9BFuBVAoL5hCr5EJ/LOsnulDSz/W
i4iaIu0QSJKXMaW3ySTXpdu74A7rae0MV1dBlEDcJtOGMf780rSFK7/n+1i1
vZHn3YwrktE1jYCaVKoNzvzJJJUYZ8LiR5Pk2OBJCFbqc4A9Uw+gOr2HH3ZT
2ymlFh/bpLxo7xPpdRGIiSW2ok43RO/NG+re1wkVMax3yhgmDjZGQqMO21js
n77n8j8M8/fkiHCA9CcRpXnQXpnLTqmwCVmHm7pj9Tbple668S357HGV/Ijz
EO3hj6UoTZKEqZO6I44rz/82YRE4It41BvBUJfE/RCBcNJOLmQ6J3DVEExbo
+TI6rYL0rR4Dh3TsilVEcYFPgk5B/yswSCiMRs4b7vj6MRqsmvKveMx0ftBQ
6GiQCJRsvcACgLHsd6ZT4wrPglNxI3RETwIkW5YN7YkSNiQgVfhFmaq2Holn
9hKZBZEbCNnOv49Qj7DO9rosqVQpL0j1YqseM7U3N/4clz5taNZXO29oengj
tBVLoH4ZtOM/cMVj5wfxUqLhrVUbbEDUk3RiOUVKS4eP7k3x8mmf3nzOZI6a
tOSAZ1w+90wQzfW4YYXfl24/z/I2cJLQOScgLzMxmsxoeQUzwe3RMD1ca6IE
iiMOgPh/Uemv5lVxOwTaEw5H+8VqQnELEA/5S9p53L6HRS0PU33Lo+6/AJHp
WnPcGTONXCrFa2P7zFtwnvrmdaxkNzutHweuVnbOJuORKH/Umb2TvDEcg6m+
X6gUhZA+it2h5e8hsfDfHB/vBb4l45wLQe/Yyx2b7Wq4T0YmQ7foeJ2rPjWs
tSTteMmJuUfRGsCvUXTboAxHUtiH01szDqAplvXs7OaRdRbVOdHgO5ayyZ7Q
+j/aSWJsAfOAapcK1Exb62bsjwv2cBXOKZ6VDR5SWLMpe/q9aEkl/ifXVvWE
CdlRdFrSFY/n4st8sHX5mKyxFaJUN90rY0lP4pd61WPIEkM1C2iG29kj/iZz
7k6nB2ibGY0ozHmrzdWhK5MrpTpCfdvIulL5yhxton+zqlYqjofhkaf4vhNR
Pm1zMPHOVccngW8yYmnivo5gGiT/1znoGdA0mfo78o+OMzm8aQCsOoEVZKMk
0A4PlRqkRuzX5J5hgR41b7+d7+nX+1wgCVfAdHjqErThMEaRtgVXsSiyya/B
K+oC96BTcyB8Jd54PeHHTn/aHXHhP0IdDT4XNysLukA2wFL5HCrroSDKz/oU
E42a1rHjtMU+X8leHAFaYAgcK95xlS45YrMFI3AmMRLEJYCjGv48xOumm83S
1of0I/Z03ehVg/DOfGPNXdN3VwPxb8bwYF6zLrwqYnr8WJQ6eOSYj31OaypS
aiF+8/G6s/BTc0XabNTCXxWrRzI3dX24DkUZ1YHMp6eVIggbcWJxVMbJV4Vu
sQ0vzXkEeycadf8tbkWtJ6jo2zK9eJ/R3+1RAX1Hgn8h8nUv2CqsqxNe+C1N
vpok5a5pMEu/AbsBkBRkMR8FFgSOwnOOoTg47yjhdWN1FUT8ZDRhn5zRZUun
y9rCX/dlMF7TE/wh9Jhx080CwgPlcVVT3QeCSDefjpQW+/WEh0s7gKixmDeS
lS1mGGZhBZttVQ9kk1RwcViYxyZWEag6x5SrsZwbTnuNgYD6gC7R41uYKPgZ
BptC5hIsxMshcY7ae9QZKoNHb3KfCiaNf07xbmhmkjwnkBlZ8xQSMtzfya6L
qkiCZPR/yvO2L1rCfgd7nE9iuUOCFg0FtqoEv2M6yNOUm8ySjPUrMqa/uuW/
4pP8r8iLbE0NaUwJqlyXbroLgFa2kVawxp9pSvXPWHVlFzuXF7MmWo1hCdI7
HF31jFjyY9WYNe5/ANnbTfkvj2letqWMfBbztqhMCDELxxUdwSasfh7XQPSb
MvYP5SzjqOCY4g9nXgIIZrr+4SCLjs9dlsXEr7DpAj1OIwiB57SOB48XQv7E
RxT8Xbif7W+LqwvDXjFoyW+j/tI6QJVdRcKLXFqedMLry5kC4q2OJ6zAj0Hm
B4oohD+2qZjEG7g3v7ZE+inw0GsOsyfIknTEB6XryrldXyQlldX9yU+uZVtj
mz1jE3bxuHoVixcrChJjJo0thdmFbPtO5O42slvKrBI6d8+4Jh/Tl71Xoot6
Vgdm6t/jCpoLU0/mJF61V1CFrALurgLJa0MxibXY3ppx4iNw/+Oqb/0tqE6q
L87RAR6xHz7hgd5kReSJDye/RV5WIKxzcqSSbDYIUjii+rirLLYIBq++j+3J
lGXgTYtq1Ta46cY3FWJYWnXBbNEOV5amIOC/GjNLaHGPt+/kTmg8rxKQJOhx
obyICosl8eNyGRzeItOCQzAFG1wOyO/m/7ViQC1JlqgS03MzjM+L0/Cs+B+m
F0tly+viomEU/B/wNcb5xGjzG6oVS4IKuTeMOx5QwfgLsz3VRxOjb6nj+kNm
gkOY748a93p5rS/N/vDBveKyd1mEkp5gvELaWudqTyk+DP+ARmZI884NVeN7
Crkgo9UZs3ukGCqgj/wPQm1yrYbQJhCU0utU0QppAub8aN3cuVUwzRfmHVCN
7kjYAsGMlD3iNkpEBn2CHvHrBpoN4gS7VrN8Vu2dSeFIflmVJCBk2zFCMjno
G2myXL7tJQF4hO0/E045IoyUl8srk8qCSl7NU3wHYd0hb/1ZQbQWMKcFVBbz
zMbgq7qNBthkaGlhnJCi8dLodfX1//Ghf+eq54bf8C2nKtwuJXpkPBVMxCY2
tdGJgycQKVbhvQzlAjaLf13oJHvjkKS1XmHml9rtTC4J4Wr6QIYTzls0FCZ5
bbnE3Y2PRDcQMee6GEE7vBlQj2qYFyiHaLMNw806L+KHUPeTFaA2WbUGI47a
ZOn7vtbL36mEYHr1rUhBq/VhnQvNXWadtWkU03f08/XsuDhBtT58cNZJbE8s
cMdaGVas+2Vok85iPbArRa8NW98m1Y96Ea3x36/bZZJWUCKfv5BE/vx6gruD
4t6MIv8FDUDeQGbq1DVIzw593UpI6zxPLrxaHMDRupUyS5z6hBY4dobyoGQk
og7g6VdLgVGFF+HhOwLFtFYDI6oTetsBgXulEXonAhuAAx0mOAogxzcjgxj8
cQ0/ttT9F2IFbb8iQMLnrUFRD3RewQ6kMs1cXEz5jiAzHj4Kt8QiVNH3Tewt
EY09rKAmBs1J/YtYAoz3OdvMX8KyViPwkMnGy3MihtstzA1syzde8DoSEGbB
kt34n768evneApZhj0Lea0NGUM4uJq/YS/EUWN/Hj/B2BS0mdQYdiRFGmDhE
BTrQB30PwxxyYunYYKMv11XP2wWXD7fKd2uRO1tHZrvDZ7vwDH2BCRKsqDjo
QK2xy3mp3eHX01V1ZahOZC5MBulV5nbt8eLfK0wzvCkJLaEH7H3MHR6gQNhP
bmar45zNpCC2yF0T3tH4axIy/K+jJPGvY+OZNw7OZIN2hyIe95dYDQ876hSU
I2YvULZrfUdy5xPSexPF7IknJcPiZYm2Frd0BqqYD13xCCi/saNdrAJ3iADq
7KdbKteeKcEN6OlmdytPcGp/Iup315YqK2x5ETiwIMkS4+xbzJ1AsEZvc33d
LrIXBx4SObACftxi+V1HgTq2uMldiv0byFzGg7dEIddlxnTfzYS9AlBWO0mo
TcCnnpqDO0pKz/5QYU6bgkY9oa7tYIfDjlm3hos1P7fff/A5HsgWbY0GmY2v
6+ecM0egOIoxSQXj1vk9OJANhW1jiiQ10iUBZM617sr8z0ir3fx5ajB8tqYY
tCJ0w6tQejd1E6RWVEltWnz3HliacMlFkGysZNLg6S8D68Fq9jq1PRPT031w
WqhU86d9BXy48WvsAicySRcju8q3eT5ioKn2WkXfemjXCyjuXzCS4qBKcRw+
RWmXk0TGt9KKeZUgUw/cTDw8FeeoT8I76czHy5NopBFDxTkWFSUxbEUVkct2
hu3Qybk/ri9oh20UvhgswLhviWiyWcekB2Hgg5689PWrkvZjNlLzM7pnpy2p
v0/Jlwfv/kQPhmsat24tlJ0+SNLsbexmujDxQeyOsgt1GXNrvsqG1JSIQ+VK
zQsJFU23bP4OCLIiAETeS4S8Vjz/H0prTlTjFQSQgsgl3P8dHLXO/Tr7eiuZ
W33Z+8vqIex2sk+G0B48oje0l/DCFct5cQ2PBz9ADItRBXJqc4HdJSWEQF5A
cmywz4K1NbXu3WR2gkmBe+L6p4fEJON3jXZOppbL7QzG1CvIO3afZC7zB1AV
SKbInjmInbdEb1LthTlZssu9zbQ/Ycju+8M64SkbLVx5H9Asb/UI0fX59Nch
C8XEX4WljJ0hQ9DbVdr38Qc53uXI8Mwwqrm42Hih8geV1U618QIPce/iDWVP
09zbfuboZVmtzNkG9ed4Mzm0aYsA0jdbcJ7spjNW0ej3Fy+yCrb1ucb5Pzwf
NZqdElLqQ9VV7w7jGepXHbF06tH8LoT72vOjShd48l+p/VhDmFxBTUIFw6nD
r6JhJryRaIwuyDX089AAVZ74W7S2pnnCL7yFZgGBsgh96TSNjntuWE5nZ6oM
kqILb6S+02rDfbsiNyaqvJKivaW/4QiVxDQwOJ2o0JgB9BAEm2CpE5TgiJLC
f56ppazYkxwFN5FBmNMn3to7XoEhj9BMKS5gn5P1VAUPswme+QSI8gRfkbsG
lAN3EttT/efZxVZYLk8tPW0KQuUUEWQ+satOlx5/H6N23chVK0+BNDZLYErU
Ti2zUaWj9HxS5S+vjjjJil15WzHvzGJB/InGFAJs9/PQpBIEOJxKrd+lF+2s
HgswO7PIzo7t4fXCvWWdFFC8zMQR05HF+kdErM9sE7haDxqk92tmPZzmsh1/
NeuVm2mQvycctIHxgkvsWMGH4rdWR8vXjRVtuS1K9NHj3A+8g/wChGwoSGfU
exdaHp7FBGw1Fr9uer93/5+rMn/8S6hYSF9YigkpYvGS9zPHZXqIrSTwt+6o
KQJYO4xnnpte691rNp3B+ZCrG15zmtnhFSz24ZP/yeEPXGx23qgG9CiVc8dp
O3VYa1pYBoM3eKnvp5dy2esw8TuKVQkZnDphnEHf1mYm+2N/j7LQ9j6pVAqG
q6bYhwKRBqdKEK7wMbNuR0IxNJamWA5bManKgS8LcLBvA+L+GMju2/+Ia6sH
QXeV3XBKM7EwzXZlUxF9+Jevtkmh/8RUkvZBU/ffrmHMHGBRGf/n5W99o0z0
/mvLbJJZLTIYTR8HVReKel3Jv3HqFsNCv7/RR4DPNBIgO8CpdpfafoFurSOP
NclTthGHYWGomRMDClKNHW/VCBBign5Qz+C1CL1YKUVn44ohCyE1Kb6F06OF
h9cqTXqKQA+khJZBA4/UF1AEZyhxATOp9TPQwbjNZiV5OeAgQIMvRajr+7lt
qxEdPmFp6d5ut+rkMy8rWLcKHODgD5jRxTDDXocwEdgtC2z9Sr1STZSPgxdi
fgVBEZbP8s1wG6qt3q/OvLQm11oqXYCYduv3MY9XVYB7WUitO/uzgKg9KYtS
eJd3ely2RAwf7T2tpvu0waMK59MPJxShXSSaJoDuRKEnqT+x14yYL3F7ZpiJ
farP5qKRjK9iSJm+T4M0F/kXSdJgVVzAg7AWsTAWa816O0/VFnK5E8IfWVn5
ia4E6yZA36pkDNNPOPCEHBDrakH1ZBF1ZdfgRkeMNrLMDA9eExpq1cApTHDf
ARj0qO8dcC0iaiowxTdn08vJyopLiYwtwb8nxa1D6mgv/JeLMQzgVXb479Cj
zI6a9zEIRrXN+4puBNtWGmhEc+0JmtM6CteDUgasa7zir0VnNjJRykl/N48t
kQR4sX5dddyRR54p4HNnNQeFufkuu55CykjHwLjvpIpXpfmoo53VVI0FPnhl
rsjJJrClNWLzX9R2zMbUq6DT1u4vk2s79/LXBjdSBlyXRewVgABlmB/+K/XD
kqmRw1cqjqq2rczRZsSbvvVEIiu7VVt51qOvD2qd+3ABjeR8UEQQucPKeN9W
AB15X5y4jAwrjQ1wIspgRqHIZoEgqnBOBzsxpctNxFlLqLoAs69za1KYhDjv
q6Bqx5/MHnTBKntknwjU4PTBaWwU214rlxJ4SMpTLyCbAJfMJu6vkUD4zP12
d8ff/apeXpeXp07OUPOCCYm+YdjHHPfoYVYACg/ilt1Lq3CYjkMzHbluSBgZ
FlbCE5Ru9ACCAP0zHWtyFthD3jPPlrxc/k6thEQTOO4I5TUfcNp6teN1DKrZ
Dsv/U0PPuQSggaU5WErOSvRV2+au7DQW9GzoR6DZ5/KI141SAEuA8WcP8qu4
pd+ZQWuPdqyqav/aKes0+ybZE2sTdzfdD/8reC+Z80d9jPvhLQ5RCL4cJYoP
yn8Af/aOekXKzQEabVsBteLpHyWcazx9oH/LBKErPRVgFs7gXaIslaxMw9+s
NDFa/02jAj0SigV7frFas3lcJ0yeX4NMdgNVULCHlGrJvKda6nrkhAicOQXj
4iDajHafP+aGtOh5KJC3junxcDbbcnfnuJPF4KMZCwtnaulKrmMQ1bi4cXEk
XSST2nn92U5VFBqnuWIvtgkYD1iX2c5HgT1ljK6pb7i7/hshUfrpIMyEsKan
tv2mvG+28p6JnfAYAoQ/qtXgjmAHhFeY6X9+NgL2vM2oiU18njT7vP9vWOrh
uespVah935ZnjpgIqzsADPOQ9LaeGZmmxsiIFVkdCI8h8cCyyFs1tUe5TXna
g1+MzJT2VGKogzAsw975tnTk3cEuirwIc32wsLt5jtj+aRf8YosCOSlV0iJv
cW/tW9sbOOL+4F3AV1+aIC1tLtzT9YEk9sSFsDFPUw49FFno3iCD5NbPGKDY
p1/y7YXTqZ+zEUY5poIUa9AgWCJ6LI6FN8zbxFJ4XS8VQuC/V1dP1HBSXmTE
CfXZRe+qCfr+DCL4fq1+aVcB+KM6HIU96rCanOjxpyS9/qD4axZFbGRxy+Uy
iZ8PHaBGQA5XsDTmvjQja+CdzCPWIML6e+gICFmTIFmdvMAu+r/VywxZ+5hD
H7JPkANLK+9DBOvetpYNGwFSqSRU4B/7vzo/ulWgiwWInp8KkBKKOLZS2LLj
zwrUSoMQi/F9vWMgL7qhFUZC5OpSP0IrAXj0XOwiTqlJgQ56kZhWA/OmuaRU
GpRlPENIa1E9ljYbr16MvXT91AJ6Lb2qkNIMDGQo55iJtJn6A+yO7mrFXE+l
5QXLYxE7rhuz/vDXY39GBRamqpLXAlMZc2v3k+155Qj9YmhOaBp70TXmwT55
Xjq7uNXOEnR5HDCiSso1l8kFv34Z8OkOYMiDXoJuiApvUOizZDzhM72dn72O
inZnkAeCW6tKIs4poMWM3dLXDQ3oQDWUshSRltFpAFX7LP1IL6pBVVbM7qR+
nls/jRxiMabcG4nFjqlThW5OE2t0xnJKGzEcJcHuPBcnGDEvuryVt33+taBS
f43k0WQv+bPoA7NtoI5AVwC76Zg6cKAnSWo2kGOQQTiyBrpY5Ed9dCUTpwDS
NNXp88l/TTiBbOYbN3TFlN7Wehq7ka01N+lDenu9WtKBQbTgV6ClVCwnETof
QHM3LEnS/Bw9FqsohyFCHacfz9TUFeGtiqdz9c8uQ/LKGnjU2lKhBwj3h8ZG
MSJTrQmHprMMwG7kXjYiP4IPr6IOyPvPq/qi2Hq1rcBjRHRZYn4EIzHomDfO
+7c6MEyLyhRlPZ4pPXzVFTEBMjRDIKDbhKrFs2H1fAImhShtprRazoxgyObK
Pe41ShzPkE/BaYLLhFFtMNSOefr1tARE0XjJK3/xykvRBodtrx2DAo5c5Vip
7NOuw8aw0w1MsLS4A+/ASDa5gdaKWh+INDwXjJnZ6lDm9Vq31iulhfjHHzPX
0CjogUrw9M8o0MBzFiB2HdwMJAhxpJJj4onGrYgQPOsTl90zvtPatGaAY/tD
hOechhSaN43DEuf2s5d/HV0wnHUd18JNPaws7YpUViTna6WFOgUwokaMlhEI
HqYu4F5ROEh8xSikWeP7V9kQf9jZSZDP266i3xcsLW1ofXLgfey2MCEyXjVO
PtwExhqLlefsLiRvkwUUTFudxHrkZpJIM2EkaX5RvreEBget5TeMS1DMXLzv
zmbJGx7Jg2pXa771Z6gmFallXy+Aomuzeq7u0yJa83bBUFbTq4zqNO4xlOgg
Z0N62yING8oOI+KdqmNuaLdusCtconDbFIZQjBrCXVGzuOu6MaKOydg4EtLX
wNBzBSy5e4dHEqaY6tnG5FqQhRFKVClZTA2Gy7eWCYYIVyVJGG/by9th2/m8
7U2KlpsTIDPzsWVi48mCqsdZAmnFVxJx/X+zTcCLXYwnMlMBYlLtrd+bDp7V
TLclEbsJMndlTQLSox32pevzwmMLVw1wF058IWODE/We82CtU/MPLUaDiZcD
T0stolkzYB62TzgE9jxSl0JFQVamaR5BcAhFcrVR+ABhwmHGR1pIpc9zcslP
qvwI5rCdOnXLhTVFAsN+auEqEGaOrww3wvUT82zq3a5WpvSUMgWwEFioV642
6r1G1mhvc9KtWQcHxrTPeCEV0KQBlMaa4EeI++18vDrjbUTl3rEY87BTC4dd
0R91e0AvyGGunJ+73ZEk3FthcrWtqMdcdQ/89G/I722NtkBcTMiyHC6RCSOi
VuJ1f8VhYJKvlPEQRKKMeb6hC/YL6hwLuW004MPwnlO3ehRyaSLq6XsYcE5n
hc9b9ydujanzMzd2f2q61v5jeqPR4g1HIbVHeg7xkXJNK3LkE9z6AHopKgqh
CXF0Lr7vglYIaq5Z7zxexY1uoseg1DtzqmU7gKhJnq9DgT6Gm1uQXP50USMF
l3liRi+SzSHQaDryD4ceTNtjeig4LqSYFD8/LjWQXyoH0zzuNyEVyMuCRyXF
VHd5mlGFD3BK1czpnpR21MaTwNFDeZGU5upY/Nc3TwxVeHkRyaP9fKeV0N3c
qLMkjAlgXanO4BfqMAh4l1sdo7qIOQNimI5XwQSUoAYX1r84I7BqEJHYrNEy
mo/rhk1pP2ZCoeToHOpuJml1Us8j3NsLt8TZ36pNcL6eK9whXKW4a/492PLc
4Dahr+YZeBr7+o2YTDzH2+PBjPvwipZcqqR0Hz0m56KNa+nigDhD0nQYBXLr
gICpG/0BUomfPH+YokgNHLD5aZ5mww1oUubOc9/PUaTHgBqLLfST/CDxje4k
4mL20yREyODwa+GekDnyCgGiszAA0kZb6h/n6U5ElicPTIS5+VUN59vduZ4A
JlubVR/2pg1cCCoFZ94uCVejmEn162DhcJFgW5zf8dSgby4vtOvXa0TGodXH
Xcbo+rBJJgK021/t3EhAn1J712A1rwGzhwfK3RgZpPrmqfNJV6+aNXhiAgK/
gc8vnXxf2XT/V11JWmHBnL+GyuMCw/vLyn6HdhZta3ScTvHX+HdNittseDco
3dJhmlwYRJswa8CIZfnD/C25kWekZrQ3MfO2ftjZrzsqsk3zB/uQLJuMkWuf
5WWA76CMt1CL6k2aAQEngEfTx5nsmSZo78/rF20uds2AWBAL4tQc4MsosJGx
8YfEoKV+j1Kl2VRJFCceRoUfPkkjiQZNbPMwcQXcRzXTLscKZ3MR3pvoCOPx
6CweuvpEWSQ8lw822kaPYm2xKepnhQl5k8ivw4OU80dhV7GeuLgcKtJ13XrV
7Xu3eJhzqtv8r0JCZp1NI0NQIFfKe0lSLfKiOhBDQZFLNFkNTKuxnxQpzZu3
r0TT5YZr5UHoPl5FoWoC/B+nXZfD1IVxvrQQGYumeQmvJymxOQa46fgJ7U0H
SugzX8r2PwrgNAgh50JQmdrsDzCrD9iF9HFYOKloT8VKKE23u39eNYx31AFi
mKC3MaJpKNKHLLtkN3tLoQi2IbNEoyU0lL0D95aF1h+tTZztezJNItlBrXPT
Zm/6bjOmiwUtEy6MQQzjnOEDDiZQG7LIHFav1SH6v8C5ei44BozPSObBsy1k
WQ6nV55r2feTr3o/xU3Ppl3lBJbaaksvOUZjJ4zSDWud9YoQ4w9eSmtgqOgH
UPuTO/Y+0B1dokbTJirNm7bVbXx/VH1si7p6zkVbDw+H7IiqNaVWB68q6zIo
9BSEWUjCUpMhSzAykukJqvzm7cm7EGvLGxn30EnnKvIrivRH2kgF+FMFtxn/
0cCiha8dW8esI7VdE3hgT+2T8Y2A/x6RY2vRs8wDA6vugnydqkXFSlv0NqTN
FA/qdP7IlalZ9MTYAed+yKCntjFFKrUkO4nXNTGCQ2bPrMbNFxQQ507K3Flp
01LIDXlivJnF28Y2BhAwCLEx5luYHmErxUPXjeFF0mX3ycVvJkLUlr2JW6hJ
mSAGmu4FPbMez6jcWzikdfbNK8UBc6wvpdGa8MMOmlhZpk3VnkrmFhh3DULk
QbvBmSRwM1D3Lx8Qf5BTdNpGO8yrlSFqN82Xx4/EyMrOnwNzZl6SDSh3AFiJ
0Ll15FMoVsi9bjSB9TBGonfHRaRySoD/BLTQ7dC1trebn75ET15Vb+PM/H0q
Y+JCSxCHTOpFpgPBJNc/m6SjKF0sjeepyA38+gPlraCcI02e8t59UAZFbyxY
tC8pbuZi1H5FbWED/hOMThM3DF61MLSX7okA9TqqDeMlmN64SHBwsZ/47YBo
ZNgW8rrl17ofNiOJM2pBqxfJd/7pCdbo+i2OYqRdwJm3sLOHqebipPkiUgaV
kv7zQsnk+I3T2o8wfL5Jy2wicV3aonO1z+NnF0x4gNDljIlh6p4598cNPpiG
wNVknYeeE23QAt4QLU0TAoxqvglmOnfzwWQZishI4kxl3XtwO9b80avF/Mgi
RMTZ4riF7GwcOJok9LMAbfu682FHGtwOQlzta7Hr+GgnTDkwMOTNggfyA7zu
sPAP5g19qsaaxqmzJ7MUVuGgBbBmM5CJBmH7ewdnC4IASr5dl7tlqyoGDWgp
0Wd6xFke1TDUNY98Ft+iBcO7dsuTDVKWo5yIIo6fUSItJOR2As3cxZHAwMlS
gdZZqhHh2BMZ7M+QAMZZq/AKHlhPPPtxz6vXYaFZJCHBkm/WLMJqYc5QpvFq
WytHbpZdFfkjhHqaDy3lt5D2aZDIZKGBio/HrRpkvbP5d16WR5sqArpkKdPu
nKrfFCBq0dhV65W78gvYuOVlaBzC9qi9M709xk1Y5EMCLQBNAsZ35efdBdO9
Bdy6+BwD/FI1Iff3iZ+fixdyR4wRnQk+HB1+9HMIHuPSCkL6+r1hioWmqU7n
SXMKy6m969S616/Mvq/4el4N+wKKtInaBD/5eirOKg3OuiB3+OtAlqa9CUfq
pcePRHOWEiJh18sXPnrhBctMD6qqSZnL2GupNWFYYRgx3aFy0xJ7aq7MICy+
3holJWlnlIpPWuXOtNnnmZcLLvIloedZEgu3rcF8bc+aCarAOYBTIX4Je28f
MddP4jEbu8PCIwMF8XanbhgBAaEY3cpWnjOh4ZF6OllYKJGYcONDLJT2KyS2
gfIjWeXU4vZN1WHxVnjqUATnhfiAhZ4iYi/orGHVR7YMxdiuMgyFHRy1nHTq
eKrLV+ZpuzsbXpN4vlfQHZ6C5+qNvjKoKYPuFqc1WclAFYD90kV3mTRk347Y
ZLd4SpzCsBbh5gVCpPwUXHvT3F3jt+94iKMVwRDrhFzrPsBnSMn7t0PrrqJx
fToGCqCvcrl6rxxQfJNgSGk0ROseFk3IJhwTmTDPXMh/T+XVfeWOXz0noUr7
hHpXT542yMqxi1PQSxEyk9dK6oAtna7t/z7IPlmsGx1uUR8iR4LqiRvWUEWv
Lbev1uk2ZUI9mm8I9aizlhEBR2PY+jANY5ypRO/7v2Uup/gqBhEQfwavQRno
pi2kXL2yfM+JUEh3P2OIIWwX2hQHfEKBhfwplUxMhjLP1sgRae6lhYk9VBF4
EmnTihPddjWVqxDQhSlcufyvMpDGnAOUCx0ZGsDumPwWtHssScrlSpb1MAX5
Q2bWgJkIS6eOz9lEuEgQ5LUE0gXP5K5210Xn2lK4t5iHo4SUZ+IDOv1jvY08
bSj+UjXLauhS4/h9ikO0wKBrduPIursVNIfYcnOGJ4GENTrhc4zIsuun5MqM
qZyxRdi1peFAs5PdoEZiaiXeaDKrWLB7QWUO9bK25LKwuxip1oC3fXIGTD/9
Mslqc9nsr6mIx2gqaVdSZCpcBXtlalMv3/ytxRwcFpUPu/Fa9fS9p1DpHRuq
yF/wi1emMFOrPE0SnILfb1MHydJIcNgGOiqdUFjSeu2cimdMA0sM9LoNU2jI
p3DC51lwA0rW9DIc1WeqnJSFBF1H28zfFbPh6JSRdtY1EPIdARk0TzVVYeYl
qPdkTeFUlRR0dYAf620kP7HrrQ5+t7fZGjahOP2doQSscyNiKMYFjFwzQrlc
W+dcPjFvTZHxBTTQ6w/4p7njmv4NO6G6Rml5qsP/sKDI159XilqM2Rte2/S1
W//nLNOJRlT9RTo2mPIdXW6pxSFJBYy7NczXauAqC73MOfrtHdMXqwtuoPSn
SQpW6V8XhKC1wb4aBDK7C7U11VR0dwgie2hYHg3uStZwtCzNr4uX/cDUUyBe
q0EEcojYhlvfvTPUFu2LUNFeRmdt7tm13wK8G0/h2Y1Pv9PmFLw9BAH877cl
rMy0JedgYymSI1uK1diT6SNqtoTed/AxonkfNRdrB6oU7q3oTfVlX5adNntU
AoRF9u3XFicUPJh9YqCchbQKDJpXCOFT0v1TFa530OYvvLCn2mp3mByoo6FF
AIVMJ8DoTflFXeCK17sqN5d/tr6Dw6pajPhnVucxYsuQiE7mDi5TP50a9mPu
L7pqJBQVrmMzhbs0WxNrKQsluk5ONlQJamVjMT5J/Ek1ZCsSPg+999jEdpPJ
nzro3fEhrpvHw+H7cIiHWBPrtkI/2R1b0/LtaSU+l/szzL+IvqM+j8rXVHpG
Gxg72F8ZVEmKMzraioeT73pkG9Rr/Kb54CNT5pZPSRMP7/Mt634eNGWqosVB
YRdDky+omvA0v9Ew5pY+EPDH2iuQ7bQtC06qq96IPMJdP9yY+qwz73ZGmDq/
ZvaMZj4qiqPmh+BjXIMGnucXoOuZK6LrSrOqGyyU0k8AUhWkp0hY4R8/7pEM
eiR9O7vMsu6DmZ+Wx2Eh4lokU8hodo5ie57Xsy6Ubxkeylrm6FuHT0pb918g
62b6D7DuMqSfHgRVFgi3qCEt9kn3fW7A4NMui9TgjMaIehusB4t3O+5gnm51
V6HAscMEaYUPP26pr3wOxIQQvurUQ8CgTZF6MkheExCNLjPPQ9nmpbzJbYbZ
YrYyXSmTSKFhPygbReoF1/tdKLVo7aI8GDI+vx8IeDrx9S+QQe14SzFYT9UF
uhvX1Fv78HtxFTk8JpIjsQJ0jq54L1StQQSOR/IeYAZSCsNDy60OYo6xMPx+
jC6eEPgKPyDlU3+EW8v6YDCAzrEihaLA0YsiPjobJxAGlmda0Q3KbQ2nUde3
J147WzU3UbmSwRNnKPiwpfzv60jhC0E/cwr/nOtTZJfywAlTz4mlex1SPGGR
evuDRvT/tGXBrjy3xWgLiiSX4RqrC/Pg1nyJoDA58rIwW58ayj9ORlze96hk
/TB2WLUERm/oufhJuKB9hRTLgMq8+0NfeYf3320Wstgd7AKtjGMbOz1Mgkz6
UnVGZdc30ooFqx+xInV7q9gDbWHLXQbHr3lxKtPwG1FlZc6U/dNtzgdKsify
DbvS6ib/ZYgXl/QJI2pN/rOZTbAjs06GV3E9zlYwAY0ofCl9Nzub837FGOc/
KeN39/fxJzCaqYKH2YwqA9/V2ys1fGJz1pBgV17O4QNDnPnRpybZu/RcbUNW
N9s95eiCRwIiuDI3nWa6jUiTOIe2fiTLBzl9+DPKnhnc6nE34mDrXUEb2PEh
aLT5qm024VZeJp7WTyQ6S1nGJsrOYSiGe7obe6gbFcfEOArN4qoNmwZNRrtk
PQBmxxQ7dWmXtBhn5AfqWNp1FQlLHKH2A6maFK+5hKvnVDf1LsIDeetCVfXC
dqlI1Eg7TvuXTyTAqJbqDZcYNe9D4YPFViSqTJZPdhkiXLXfvhxcWtlA8b9Y
/0IhFuS+KSA3xQKrSngKD7V/6osL9e3Xzzl04Wsh9LThpbReYXUdHEhVlwlO
nracE/lKX9sevRK/j41mIh2m3RNEWpB47MguCpTcd2fiy2ERl0cAjYGrIzQQ
+qyQPd/WyHfnG+7wTfC3a8j2egposQga8FuHEKcw6vVsEHuJOV0WO6Oq5o1S
6plcGv8o3X0UdecfH1TTSlyMMFAvzBmA0SOhM69q9evAKopFkJrMfOyPFKpY
4RsItWz48buREdXewondhYJWVMA3QEf3CUkNCoGsnth3e7cb236DW+ZWd1lv
YRiwD4GDF7x+IhnN/3iwZkdQxNtSqUdQR0zFTulsQlVdDd7tCJ+lC67ZAwAQ
L2ZV2efRCVk+SNuiK52Jx/qfG/NEo4yt6DJwF+3M78XrhsZfc6dcqdgcAHoF
uqsLpOJ6SJRpVSHujNK5o/oHkdHG6uI4J57MlBG4Ymu2d6S14JrkGPAvk+2Z
hHWDYhDbczi7vkQuajjvIJB324G7pg7LQwuZB+rfaNUYm1nfUXwLfTZmBhDy
sYNuGnFt32zVd3y0+ewUQUIOWW9jV354zTSQ6LFUxEXAXvsZBN6G8gADgcOS
bRrtv0WrZokM1exA6AjGeN6F3Avb+vKIn3or14rW99mJRwAVTGr9R+uulc2L
YW0GX9iZvToBC5bIn8Hqk3ox5I4QHP/pqrV7BlTit8oKbBmQLdvqH5EkH95u
ePKobZU5KjUSKjkrRu4sFqdhBKMUiDpThEDQyU1MNYwhfKGCOHiGmA0UKvi9
9Bi9dt7HQstWH0BSgqwJUMot+FXXXe8c9PwEGsTq4BD9pQh2JBoSi4Chscyp
IAlZ+AvFErNBJQe0jBlAXpbJd+XuL/wUNxuhIu3KH3dMZ9yQYKoOF19jVGD1
XXkyW5kMQMM9qxSbjhvv4mZFDEZdvy/JENlzbgezEuEAnGJKRFxpFh3U8BeD
rQjp5wxyT9JiEpRiVo9OmuFmOHYNUOdE7PF/cEAFAawAs04qOJ268zf3p5TT
8MlGDplCsOUdfiBynbd4hqumF1RfEZC508gZpLgISapHe8sau6Nnu8YpH0Tp
k2KF67o+smoFb/8Rb2eQ1e1WS/B3vfLuOwhR7AjOIR/nJuh9M4/UzVUp7vP5
qiZQWHUJxcIMe0ng7MWrGhf+Xm1oV9gpAU/+VhvRN8Bw3IdmG4gCEAeTT8EK
r9T14+QGOBKYmuhGAuSq/NqeQUgkUxBO3ZDWvXh1RSDCUWEEJT6Y3lCJzxwy
vMntId0DmRAhGir6Ng8Zp8OTeL5pg2+hM69ZQn2uyzOJM3awAcUVw8xdHsBS
e/bPRepaadDXyfVq5h3jAOLg9vV10Y6FzFuBKduIQ6eo2mVhw3B0hD2VfYIP
R6cEz0i/4R9+gbylY4i3Up0BKMbPtzRY5QJqsIcTglUFuCtDuBJN68sFIa5R
s9Dpsx6tDy06SLnXQd5WE2lnRluw1x6xEHveSvUEJP8VdK0l7D/r4wBh0tuV
131UUOtQRhnfFs+0KgW73JxmfftBxp6e08dvrbp7v60KyQSk9Tz8yRyK0l9t
fYN9+pxIIufABdsV4HZ7LPDuUDLdVCZTv57Ja1yv8DKm0EIBB5nwrh1cz43+
Cz79RkY9SdiEgt4qpgH5OG+8PTl/6Smsoszry/XqwuhpiCfCEzSwyvgXLUCh
fMpB6U3Dc1ehoS6QRiDz2qY5Y6Af6KRvi7+2CRI9LYfDoTrrtAJzJ/y7/1sk
foW3DmCvqSH3sJWlpK7lTAsR7JWpB3XdAHRJ0xpg8L+ZwOqQN4Ye++bM0tu7
DPNJH1Id8glxZxgEoj/X3bIz/89TURaeqa6SKUyGure72GntFrhEiuuEWuXA
7TRRvVu6q9hJO2M2LDrsULGhpdfZtEcEz/FXe+UHRNrRT9jggoD1GDXzNPmb
ZYamD+PdWPgn2GxNZ8mUQdW27od0Ir+Vt9PX5klZfAhEbpSwMyTn6aGGmhSb
N/QiSiJLv5YtQ7gJ/KxnsNH5bZUBx72j1lbhYDnFcyPqNZ0MfM2I/qxmNZMo
jCQvt1rBwFuJWACccszTrGHRsbhjPYJWxSEkdZnie1n3IOi55qCoRTe6W6AX
wOy7v4AsN1uj9mBsnyoheDZOgABhX2ftiE1RU485Ft6qxp3mSQXD7vLZS9e+
lCKeL8/i1LVZ4YanotJ8L9RLfaz3LixxYoMdkIZaqbPNpZPukb08YXmbKzy1
gK9yWFa6ATLJcZSvA1m054Ddb0ygZWPivQM9uqalTuLhTfPuzSAyeGN3RbOe
XAEJjS1zPT3Q/O+ldBjkzqSCXzl9/5OyQ3iBN3L+oriT8pgdsb2WRodnRJn+
d2IZhqmsZmtalM0fqskGmDxg5akT3gXFzG6dI+8QWG8ZOthOPP8P8/kHsCdq
pQklTl5zL02dNArixh2EgZ/Kcxy5iEc5+m28x0A/1mWozq2NiR+QDVaxbE/2
tHVvGB4253pO0MS//uDy/bqjmgFEF0nD2nW780eNecpcCxbQFTbJA7aSgfqC
L7pi8HvmZDPbRjiO5wrLB4Ky9N3SVFMoZiU5UiQhoaX6RpOmu7frg+4HvhHa
/kGuRb86lDMhbMSdWE3j2unLvFROJU2DN5iTkvC9xvGjumle4aNeK1d7S0qk
xUVAoGdH88OdyoEVDJ09D4hQyfjzbuv/CMDFOflsJSh+2ZIw83SWAMAEkBhp
Qh4KS1djwhXqXOh50ZkIvLbwxBvdXxRacIXo1M49GeemkbBn2XVvMmEjzVnb
OAF8uKBRObaV3EYZvTZMaZuD7F1UI7mtyWqkqlbr++U18gZSFt9WsMisV9Vv
63N0sKVfksXXt03vYCSbUNS04Kp+8gc/nysYXqFl613DB4MdulEElO53vMXx
j385sinti3+4fivK0+e2BmhT9uyYe2DYQY96QyuGfUfMUoD8enjmUnfNA8YL
d+O3vAkRH4b4TC7ZuSNsirEZiuUSYlO2Q2vXm48YXcDjnEgeevdqEalIFcY2
aRVVkEoTyPxLIoOxMyQ1EnV7QUzb+bL9ZjJj3e1hSJ5oB3irZUbiZ1fSw2UZ
Gke2lMRpm/yFYCETBqkkcN9sTj0NJC5tNHCDA8asagMlfWfWoU4y6c80VQ+V
4/ilk2RTj7fcvsDokYmON5mEfbYNhsIueHzhiaLhXDVp/atQxUXnbTgVWaaY
bgLEvpwNk3BECotxkRKWP3KPQa5aiWtPqSd6T/vl0drLu+RdhgRlY+YgyLgn
cZ+UaJsMTZjWRGg55LulUKbL1c9yDdL8jzhz2V0Yb90ROzx4qiONoPEaP2AQ
U8pC9sYj3CaOUZCH0PjVme5pLR0/RUrOi2DZZNe81hbDo3b8aXiT3TGRxAzW
1ryKC6QRn0ZtIBWoyiL3hhj5iEFf0T5sGhcw9GJZGsl9JUqXf2MUugQsy6a5
IBWdmHDg7VEmoed/wCXz6GkgxWS6Ar4tLBXrWIJeGlH+nlAvtPhPLp1rJxqB
iZqCuAB75ImltI5kFM2PFuWPJsp0xwca+wbk0MNM4LvdMmLGgU9sydlsxZsk
5O2sQ+b/UU0bD2aRuVkwseZtHRo1R1DrXGefkDVBdml5NL/ffF/ub2qYg+ij
clLHsepT/Mk3qyLNj4QxbouBotOGDZYyQCX2nX+cevZcMO4OoFLvOVgrlF0j
NgtOWkY2vpNoGQniPd0S9TS5/sUUOdrCyiNRE0kIsPTpJwURVMHgUZwsFCVM
nJON3VDZtdwjg7kS9gvBtjHpFf5IADfzWE8gv6Y4VjdwbMJVvub3BzrQRL76
SaPJj4IzMlfECUStkevRaKmpGtQb+ivkeYc2Wh+/889zfymKmCpZaO3XOWve
WFn6eUvK5OBxtOXJ15lLarmc5rENmc38V91OBmgFRCIGsRnrih6nucU1qJa1
MacNTelw1AcDHvd900E23CWMXW48H0xfBheUwSwujThHlH1hT7IgWlivc603
Wxn6w9tVuw2jiUgNvQvsuB/ZT9Wb0rQ22QHWNXEW7Swu/v61omCl1p6EvA1Y
2Bsevgd7ipcST8NHtpTUB+xxyoMsp8s+3RwMKevc329ApqNsjKcYagUzSAo8
wt2+LrMi5M/wtoPbGqWXrXzwVeaHm+e1brCNKqPPmXTlOSByQYzZGDS+7htE
ArCI0IrbpWs3JaRrfwPKLF2avc2DvYVLE6vw/oimEvAkG3DHT94EMdphWESr
XHCT4cwShvhGSd6ryeRNIUEflNqKjtKGCPQI85rV/RjzXIHSUnziGllSNohO
vO+9HNm45yh290/GDoTF6V9nRGsPu5eGCjRWwgH0KJkpgHS1Kb8x/flQz7AE
Y+zqyt1lIpYQhqWVjW1L/dCqVSPJ+DFPkbx3H20Qcy5cFL8XucKKuHM629PJ
9JqigkaHziQBMo0oYq4IHTu+6qNOePyfhC/bnrz04hZLb1zg/EWV2676RdBc
y0Pu6nVUNYXsQRe94BviIypzx8qpTrMrhcpFpbmK2KAgx+xZrFG10p9JKBmA
0XFz/CqBtfTH8MNjPjXdsiwRXQ1bTvnFlTbEpJWhcd5zb9OH0AcH2pH8JU71
6No39mPrTv+oEEj/abp0O3iytlep9LOc0jRF5fpCoN9J/Sxs4Kd0KDfBD5PK
1jqkA3w1Z6bzpkkcgzXbiV5PRaGSTzrnjvrufJvr2NnhE6LKaXy8AdEGx+LX
k2M4PUfaFglvs6B3Bq6G5P7Z4XPk2K8m/QvrQhlsIfUD42UFAhSPnHOtrsAq
NbwYJ9CFvEHs4WeyrzZUmWVByyDV1Z49MD3qJQcpVbdwqJc+tiNpM5cGUZJp
fSDj2wOb6vdcoeLuRvi2cj8aEp7TbcwYMjNG5N/VNE0a8FDJl84XMWlRXUbX
dpgMY+xEr07IlOJGvzz0i5qkar18tT5AjMVmbjxrX5OtTxNCUkNNdP2yOipv
j/ONxtrWMqIoxLZxJTZiI5IsvtlA/xtdm8+3SBAhIlWmqnPm70dxUw4IHjCu
XeYhU9RPD1/jacXBCskLWQ0/CcEwAEAOPjdydjb7PDbMQQ7XDN0aMVZL0422
04/2HS4jpkEDHLKQAeyfZl9ocXW4TcE6rFSxslsINWxNUAq6lk9y5juFuwI5
8gyH/EnkY8TRZCGgP6564uMm2ca8WsYD0OWWQb3H15eRqoeRswBMrL8v6brO
D9V1H7HFMllU8Te+veN9IEr2RRnjYhqmnRXP3EH1eEfPlWOsa0VYAQGGBJ4J
iZazRyweYNO+QRjNGajHpaq5YX2+11qbc9x9LlAe9bq5pNhz9vWAkyC9v0NW
UIGeahbM9trVYkOnui5sor/v8Kb6t4uZ6k7cuX05lTLadgruUbdbXw7F+Cx7
20M3V7Dp7iE4lM04QLklKU+9sC4nqWzWXnsF60DW2Kig5zIsPn5mHdcgI/9I
zWp33ALttyFpU3zn7BKkjt+1J6brFdgoswU/kLk5XBWKy4vj8fKeaYdZBOJE
YLb6kMWTTGWolTmXrN/25/oDn+qZhuseEUBsmUuWVkFlQAgsGp3047IBuyg8
suYfMZuZlgwj2kRvwCrZuoNWDz7yiw7G/Y/ipoqXWIbZhihGQiZzfpXscZDA
B7AVGqOHDmQaPCOuD7jJi+7nuHXE7gGTCyaxeEA4G2QddWm8ZhlBJW4XpZYy
7/czuW5Ebbqt7bRVvyfnbtKUhXjJra8NRfkjqnrpyOTynkV5Yzu0bGYyEUI3
GPUH8jPn0MsJEcdla+ZRcUffppRSgTIAKWuqWjrvJrJSoi6iRNIjcf+iXTaZ
diXsjLkSw6GItpaIb9GpLNaexJn5RWkjAtHyZATpQyxrLgn8uhZxfZxjVxKC
1E6OwjDMlp9lnEB+5aRVgDyo9UecANSsvyQiSt6forh0ZpDMwiA2XIJigAyg
pg0CuCgeJGBmREOSSQQGSC6Yq5DNopUd7c85tYVRpwV6nBv6xEKQDTtBVzie
9fBPyusRAo4LMGCyJltEgq/Wz2na3M4DIv4iFBnNxr0dDSiupPoGOGtJDt7z
yn+gqxiS4/FNebaxjEV5kndr4zOk6Fi0i9g/JzjXdjQYiSVp3Vd/jcDOGWIi
epJSrLByFBQP1Gpsy8oN/TwaBVJY67LfEe5JkauZ5up4FgsCpqhy7hbKFKTv
4MCP0opk1AfQbHvMQZFMi5OY9gUomM7Zx+4T8SYU6RNCaPhiiT7v7xiEPnlj
1c4RMFEZtdKpMIVtzbRVkl8qdlWBx3hWd9WgFwa2DqC7d+MKDcIrmPFS2lqf
wftnl4N7s1cmdJB5LHsxSXFIGxo1pMEZq4PAxrm5GcHbg/YWSQW/6vkpYbDq
LZsji5bcf38dCgHgWcLp56WqMPnxA8uqeAMbpH3catoQTmyYETdYrHZAuQ/r
engwD6XFDttL++t1Qco4y0PIrOHBvesNGQ00LueeJLrERtt73sBYl4jnz2ZQ
GjfN+0L6lyiHayzlbF1d+khNhGeKzEfD4Z9CPcouk0+ITN1Xv5VeaEXdqNaR
NpLzgYRw0Wi5SmIRgOy6C4L/reDAvvNWGFh5XHN/+LNIjZb6gREQvKLOpTIL
CTJf0z1XdNXKu23Lx8ZcmaKjB5+JJIfNTTpgvBkx0XmY4YikwjoH2xhmNKSz
SkvUJIvD+RvnbpJ5kUZw4yNRMPQTajCTIusacyBDbJBOmUpufXkmi/ysivlG
tnHuLsK5mPDGX4cUuMv4gpo40eQgNdMaNRTT2CiJrgGate+FJIU/XrP+6FS9
pJ8FF8/YXbJ/VjCyfeO1ntucZziNanrKqyJ2ru/JpMSLvcMmbyBpQ1Q4gnds
6Q69AmTdTkbup/6v3i4rdjcDBpH11q+l7kJ74tANuMji525Noa60xqCnholN
hyz/Yd6U+QKclSdS8K6hQMRUZf1Avn3QZykIjv9+k6uQMx824h6H+DZ0f1Rz
utbOel0O1jEGkwMViNj5ZsWC/fa6b7Lwl5YaSalMYSAJUoT/cNi7s4Uiuf6P
U48xEMoOy4K+ONnEz9hOudIKbw1Fsn+i/TpIROxnfKnPDaKuE1Tp6kZuKsgU
NfKvBfpxoFA/1Q8e/tJY6b8Qy3ujYORtQCukpmShfZk8wlFgXEsUn3MRsPJc
a9wf/Wg0Me88XvY7A2K8pE0DbSY6M2D7wtaEjf7aoCeLAnlNu2UrUt+rMCVL
SfdC66AfIyMY9PxoD75n73CKEKmg5BT5g67MTKkvpu2/k2k4xci7wDeQUe3f
8yWqhlJP2V75Bk5Hop4gkyOl4aXLpZxfglz7p8DTCSDfoWNWu5jCz0TCsQWa
NGRVGipPu7zbm+siR8sfMgi2Pe4CDNgDyXBcZx7abh28CQt6EoKkGKDiPmdJ
BjmAQm59cQ2brHEAdJEo0d8dkdKHegIi+OZpRixtkNqC4TKBVIea0oI1m0jE
YIv3lwrGX1nkNn9ZcHyRXe7KSBRXtJLHcffzFQLMA5WVVYQYkho7tQea9F3M
+gR7Xt5N0stFDdVOi+7zbVV1bnbXl9b7uy3ZAtEJACXlLUbd8ZAcjJ1BLKra
pv2wJ5XEsHbpflBoVnlLp0mMSasEi6fVjzmyPfZKpqPj5aQl5c8MzsZiNq8T
4xmhMJAVUr70Fc7wx0H9w6VlALhZCE4YoRZJgBk5B4/eh/6wb/jgSSIwPsCu
1hfljnS0jKGygFbrvzKi5BVaxYbMeBiZWovLoi3fhbZW63X9JsLMsOVTuStB
0xHIVqmC6kFKD+dloflBW6/aiipCnhUrF2cVT45EtcSjCOm8ZaqvSX40xcXG
Z8wnJQ5bJ9YPKTA2ui5/8LjogF2784gNYe3GcQK9GAA2tYkvf1r/iSNbHt9T
ARTWNkkPcUmGj7ewoT/aLKc1E64nC3X6jcQS5N2SA4T6ltXyEz6+3lznDjUw
QYxmqUpRWyV/8M5+7Ady80X4ULCdg8iqDbT9bM7uaT7KpCjYDHkQBotAnquV
rdJPMWtSCUYVZ/EvemWbYOgzVakNzfIFhuTgd/4GvO9vYECiGxFI16CeOIBE
aQLmAKyBI3bYODXpqQFE7OH7O+qdDuwfuL4LIf2OKvtdkNvL9+9gyui6QAir
23m0LsPF5dBviFnyhjkyx2+BkVOPsy1MmbPpkBBxVPIBb3IrHEIyhlhIiZUX
NnJZ802yg6tiKeAj2n0VK7XK4cyzPggE43Byvsmi1c6HGM/4SY4JMhBnA0lb
wqy7ZLrfTDbD3zK7JA6+0qNFk8VS5qFk5ANxkAIKZHReb+CBWxH3OL27RhU5
+7u9BUw82vnL6qaIDpJOzf9WctXWe5VWggjRvgWYNN4LcdTgw7++Q3jKdYFS
Yw2vi7Oe6dWZ4ujxTERs6asJiPeGkbd6WoZcgH+tjNCtCqAYdNwOpO9ikhHA
v6g9Jtl40AnsRQTu92qNcsgn/zasBhejnbbrfbDB+xnvTk6h4NUcZl3ET7zm
itD8ktDOjnnSA3MA7X0kqkgkkMbHiWMoTlb9IDJbZa09eE6OIFGsta93Wbua
LoKL4RKGsOr9wIocqLPHfnBB9iQdmV04fsdROMP4Us3aXvFkJFL6hnX8fqtJ
rBFTaZ2V90iSQBd+CiJs/o7sdjww85aFwzp/c4Jvf8hWW/Y01URd460r0glG
AHStcomJpqWt+1UDdEHL4yGHfTZomTPreIJRlB7ZhUR4e5orUsSaSC9ZZCJ+
cSLkveZKAZKdLmofkRWfM6Kuhh5sKku/Ut/EnJsDAnyMy56uEAulyf41Kuco
ImNLZ/w6e1Y01heVAR2EUe2MK6A1DSBMvMMXImrrHrRPetykDgNaFi+8yAfS
1rorHQi8hiLDwUMsImtxZZ7k7bTV4bePP1lh3e3oIhUEp+yB6o0aFliSgEQS
r/qN0VIC8PcAMMl+zwPtgQ3zZBwTbEhybRbu2/tStEULi5tUu9TzUblJQZv4
1DqDP6efIKCR07TttWMfsVM1CZq13g/VGdKfTdbU7eBBpyDAQzGB63BiqhxR
42L8qSv8DXB1nwbqj9jCM56eXZpktXhR9BlxHbXMSolpJeS2kMGVQ6yrG2V6
9M5dFBcgibqOEMD6S0BmdIMESxvNbKqlf0kL9bXpX66yBZTPuOxGQbZc/igP
/A9YlgUrjsXWHbcrLDmX76MLebmqSJhzLYTuX3GJ0D7hOYHA/6a7Eqpv1X1l
w6XbIBlThqhRGEcdXy2NpuS/qf4ZozXmcO5ZRC16992E5FuOLo0dpOz1ODeQ
htFyv6nA7kgzPal3WLpp6KyNp7Ozx/dPRsvAp+AG1nBxnMbbF+wFESUANU8j
/3xzIndSehBDinsbml+oaddcfqrf2Xf2FpVVcqx9vOla1RTE9H0IAeAWD8kk
oUKJq5l9CCLiBI99Keugn6dVeCd/L0c0CKHfaA7AN43jBCd1QxkO2WDzgD7b
KUIaLGEgf3//VNnBSDc+ENVuUw4lyeFqfGew8HbzQOlANvZTJmrW7hE9siPc
4qsuJdu4Oq4XW7TjlDkGEfi0iYmt8JK5rT44lLVo9wAAzi5++czi3szseyP6
QEoc1NMXHbRBu737syQVc2w3MoPVb8Y2iVm5bBGUJQDShteRRlQwUEWPZ10h
ru+5AaBvHeILpqFlAlt9tWgICHPgZ/yRa9ydiYhH6TYvyYkgCCmax6+ivGz7
R9u7HMrGyED28ynTVR+9Z25seIF6yzKJsLivzyfQnVTbQJcB/GPYxB6FbBJw
lW3qMnudidU0BN5fxquC6/VJPgyMGrqEVqhGQDsm4sZSL+99mvVYy39LC/g2
r5BqJOT/0dloMbauQ2yenLRsappzD6F1vja/YaTxxo3C5+Go+DQPeUQTNuLO
Fs4G+XAkiTaDSMPAj+yOg84O3rzihUk6duOFVZhBV9Vpxl6LC6AXHTxXrtKG
cafAOGQ2UMuuOrZaHy0mjFg5Lhq51QnbogsJEUzw8GNc76XpuDvcsO/tK8fU
hJWUSrvfPjo0aBHxTs+CWf5V8oHBvMfhgqVvWSgOYrc1ePjCOuarnP/ZkpIL
Cj9Ez4uPDccUU9BbZMV0MHb6FtJdXwlgUvT5Qgx21uYyMGk/x8mM4ddVHidA
KyRSmNzmv0h5TMVaM8XJP603OisSQsMcZa+wPuMfPJHPtn8htaQgJoaGk3vv
pxCr1xM405OHclEjAY08oDpmoBKl0RUPG7KSGe+eGTf1305dFlGICyDEdNKM
VR9kYg6R3GasoLKDJgIS8Di/kXc+F9HaD8H1FsmHPrTM8ogI0t63cWd5XOmj
he9sBbe52Srq0icdA6PBJ9Rx9Ar3ZhxQ6ifhBrOx3FKOKNTyqLz4hUrmzRnM
/2rm7vjkeByw7YdPX01nw3MCN7mgTD2quJHCbeNztOJp6v/La7BVP2kkeIOh
06IdZzZocEwYw/AekCapX2gdHM8z0XR2h22aNtbnrGT6ewAx270GGUPmHbbv
X16DhUv6PFq//kvAZpYXz7l8s5yVYnhhYFYifUU90fceJMcWGqyOY1QecHev
QgOWdBN78z9A4VbKPpkUe1Fr8nWhItOiJ4m6Yyvd8eQclZBuFF8XIdV8FdK0
OcliC4uIulezjFy7JvI6jI1Fl681U73RDcRfMmGHLYNHh+dmVzQ6zUZVjUb9
StWnBgeFnEaIXQgitd6JAMXw/FJnrhq60S6gnTr6/2MKuPuzRNQ3I2S6na49
83uhdmfc3LsjWZ2HsLtEejJke878HNjPn4T1ZXn5UifWZFxIPr4MW5reLYt7
0hjrJOmI+lK9iuuRFTSXTeuSdxkTLjU0YDZwb1fMmFQMtL85YgqopX41+Oqv
8o93lSzOGhGo9nfbLCOhNmiT8ztbKffPu3v5/MU+E01L2LHyFVE4ZojQ+RBu
EO9AvWxjibVjbVfZE7cVP2m5Y4pT24j7czkMcMdxGRpFfIfndA8k5sJ3i/bN
2lAz9all5SYaO8A/yatkc3aHvUGquQ0JPZSDKucSW5yqoECS5Cn5DsSoRgCK
YtnqBDXgW8dLNLKwm9KBpCNsc7WrxUae5cKeE2RR3SbmyyVH5gLTna2hVqwF
H6xhE45NdQJiBJ/jY2bPOnjwX1yq4ecQR+jdhcMmEcCRCShaJiQsxQ1zjpyY
CFe3HVUNr5Qdcj2Q5BuTG1Uw8oxGnBS1iaDyxemIk6MuQ1se2pe3LCtXJOSV
AVJzhF3F5slSvJ/UrswYTwsBPGEwFPfgWWaPXtNZeJ6ged6J61fBjC1ypw/v
QgIfA4Lt6A7OuWo0X6ryBgiVd5/Pqe1xo1pFJqCJ7dCcmUS1TodYmruwC0RA
zeWtsmSv7oUf9k2IqP1Zlj8nZq5XcbQguO4b0iT7+4mqzEadagW5uftOcuU4
jMhCdFoPM4AHqLiDr86mRQH1aA+qLKvFC+KffO0ERs75GePu7gH0gbj8h+8w
C8kpqV/E5Xg38j1kVASVmNwTcq857vxFN+HUOj4TeV++GS3wmWR7aNsPyDy9
Uxn6LwiQ4yFVJzmN79dcX6eahwOAqLi8PoJe+oBy3XQBMV0pN/VuGV4/fECj
czvM0voJCRDTxPLw2PvfzXm2jcEXERCcbdDGnH28kvgPJyKHGfx3216uv2E9
7j4DceRxInFBPOcG8sizLVzWDRuvJfVq2hm/kPHQAsWXNfGWw4XCw+mDFzjU
ty/baqH48N6pynhnrGbTvG1smX5Xce/HdPFJjs8TpkhLZ3IkPG2ZoYfaE7ks
h0fmZ4/8Txm9WPNrmJe9JPgurG2nKfJREm9BykKxRADqaqHD49ZvC7qttRw8
botgpG3uqnKlW/5F0JQ26JFhKBUlnLDJsww6GbtVKfLNo/UThqYTLKG2bhIe
frTF6f6/KATC87zO8dLhXjxI4NYiPvvMYrMVCl/CyyKLbvfA/2tHY8tjigvv
beu5WxxjgpEMSFkKEbFYCo8CLqlnnBO9/Sfihhfx2wN3eDzbYMGvg6S2p9yr
A7uNzNmZ1Jer6NfuuFyEmsJs4DySNoxqQpOeqkazAHpuQ6nhsmZw2rl3/hYj
V4IWc8+QPnJCRj0jg6y+69uchSEV99/T661pCAwzuBkxWfY/BJ74PxzKp/QX
uIFaqc+cDOeVnDwjMitO2a6ENK1T/n08kqdFzKqMSQSNCVbhiQq+r4NUCK7R
BfhwSdgSwPuMcCd9h4AceGew6bRHNdW7g35y2ElhxJCLJaZpzUpWTMP3XFf4
YYHYeadszllr9EtqL2WZSTsoTJt66msdXehNcs2buYKZA0XlDszKTWhiDarO
6BQzIDmj1ME+1+MgZUG63UuDgdvGtM7ScgpfxfmpfDJBLyeaLTMQhXrg9Aq+
xATSrhL14PWyq0ngXfWyoL1yPNd3GrG7Hsm53BsB38UCCAEVflwBNf42YKwx
LnIXabTijtQpMKRXjRDq6Iyho0MOpJxSsyXo4Mry5dQFyuzkiTMkTH3VtgJ9
/AZtrs+mvTkpSSG7K8sfn394RSJSnrT4/tGRBqOFhY0Vg+Ffb61glXTAmMD2
nPoQDH+hRNUGiwtX+PwYnRtke6PRVeeeJvjTzQD/MHeW+AM/zQhtzXsrwYGv
THF8DTqsrGy5a8KVc7nOovpr+jgpDs8qaj/5zLindLwvXV/Uyk43SY1FCeZr
nQ0kG5DHJtlcihzsZRjNC+Xu3v4oucaOmQplUez12VOke8aoqlxN2R5zElSF
gATrJBLtSs0Hu/eRsvEnPeBxq2JhYuO8fd87HfNwHbG/K6UH5Ipdr+54kLWm
wCD64hVEANOC8xXoxbxiF7WfmI8cDk05n1N6UIaYW+pHUw4oenH3iJXWQzwl
z7W1SpsyvWU7o2+pFtdj8FCs6Cezde7+6hSaBsYbju0QR4Yimlo9ziP0IcgG
9S7vrKTQVLNFG1nEIemueGnmTxm9q0zr8WbhDKJQ0EH5ydrQnuBSERxE/f6o
qQPsxOYbHlQciikzEkbtMO4zPYdQz4oqQGZyl9CgtqT19AQaASjoPOOMs8Ow
bIl/HNeJmuKnzbgDkTLhrZBZMnFsPrJbMAqcFElzOVNQ2doKV6D4qX4vRlIY
WDwUf1K6w1o6loEM2pVTrFlD+x3uqJLzh3LR6eAlqRJSZkdKEOfD2IqgtNv2
7U9zXs3+zZEZX8F4EAHAlK57GWXCTX6H3bdhJnBTFtQwxfm+AHRtlidla87f
JK54Z460x4wPb7IAu2HJU4Pv30IK+q1TYRc98lM6XVrtDwO1b5H+cNUfwNah
Pmdkp9sAkkADn6Ds3T7eZ8ZRj6zWT6TEiGcw12tvH5HQYGLX0tdDjjBFNq+q
Kw72S9jCWcUH8yeShKvZ5pllc9dmgm2AewPPJ1YB3lon6e90rs+6pOHj85on
Mp4/nONsn9LiPL/gLgmJ91jm5eVd3Lt8c+FbuvcgUtbXgH5aqOI6sJvZmnWb
8Szzn5x0L7sO8komxuk8TZjUDJ/crRdqSpXLg0lpNrpuRw0NJ58uzYgka6r1
0wJNa9NhkYet+MueS0x5i1FmzP9+GRSi0XuDnK4KEUDxSYoEhWBV2TgnbuLJ
b2CGCkmk4172G6XNjgXHrp3T8HISOE/ytthg+fPoqaEU/n3XZmicSysUIKVL
03T8avjCL+iJNY7nCmUFKH5lmz0qPEd4FH6AUILv3/EoKJ0eVN6xnh7ENYrs
gAt2uDk9wN/HpPWUeW9e4fHYTWLY/vICKbpilBpI6ionaZbjWGFv4C32LqmK
PmYoijCbBIT7ImPeFM+SQrdlqIE5JKdIE4d4EFpd3lOMFFrbJOshS+IHe2l5
mj/rgYMdxr8G1nJXMnInhF8vYn4IJeFpGyyEExXsAQK1AymBEjZfGEzsyH7x
EnXJI4JANtJmWeLY292uI4nCpPHiCgRx6IzEIqYqpKUskmQYoQ9z/vQ4DzwC
HJKuA7At9y1NSGuiEkXfQkNQfmmkb6/Am1Dr/sz/ESVrBbDHx4pBdLobRb2U
ef9/IczPxow0LRfNUHdjpt77V7qVa7Z2ndJ+D5lTSuFwVlwzJgbh4wFJjWQx
yHeJ6ikgF7d3yjlRscfzd/KxwEMNP868JrF709VL+dSvOKhs5rBQ4lBZHUuk
zLikHc3T2+0+FqFzz3ERXwCfZT4Mx07FMA+4oJq01lMMWhRT6cgXQuGFjQg7
1R3QCbcSNFPyRDmHyhwcozYJgbNpl7v4B5oK88ugsHzzrjPHtioHX1tud8vK
8DCJBOoIeh5HJiQbUURVF6c6IDod6BwDJmZQ6XMpoXlmQA3xDFjxaJIs2hl6
Rer1xDy4X+CNpSJafc5DdGh6jvRJ8ROX7SSKU3h1e7QHKZ5nxyCtrKZMebXO
0sHGT78Y/8tKNilWtwPCjwK5qW9iLX7lLfCGsVE8nfJoNwME14Q4ympGc6Vt
qimBr9BiOL0PVtstE2YLOssHWEo5kd29c/7q3IVlJ0EBwWPaEce5h5HefFa4
Eu1FdrlF4gYtKy1xNoGtlLyHnarSyjkYWlzD3XOIAwswZtJ+E3CU6PsRU5VQ
s+aq6AwyhZ11jfOKghQZBdEtBTAAgmPaU0PFvIrRGwEne2r3/tpGSaaYv9Gb
KAhCSO/qQPC3hMvZZVZiGVcvLExG87lWiEWvWvNO/tCau6SdvGBPL1zUST+4
Ii3iTClj9E/KVv6Nbp8ki9qmErx3afb0/EmLfuU2pnOif1fYxpdf20wH2jxn
gnxmnx9cxxDnjWjruzMO7WMithQpAeG7SgxyFUgEPM1XtS+OaYH2VoarlzHP
wRH0tgA0c7LbVtOPKSwolADYtohbyIApOVv8JGGv4FViHXDiUup9gXyQs2zF
qgRhPgY6Mkvh5PyBKZjN6Veu8AAvM3l7BuUMKkP89cZKy1l1BANDzp5l0OKX
32c22H9/TUCHtmseMKPEIiZPITOivKFXxWMCh735rUbNKzyjhda4mZNA7uuZ
e4QDVBwWILRezehhZX1IMuFNODKd5TCzW9iTb9D3Fb5Bv18twTpI6aW8ahb1
0sfdaNGU/Bs+qtjosEV5MCo0OYPFBLGnopicF+uooIzTAxGn8yECNzauX0IM
STL8+HfIsn5mjCSfvGcvHjHgPA7q9KItv+dxD1v19EyXtD0LeyQopO3QfrKh
O3bBSmVi2Cf6kPh4gNHQAbGOvZBxafmOQwaRKuzjG2heBWFBO+Ee4Nfw/8Cy
KkClvUPqucGgAMZu65glIH5OFYORGzrXnkrW2ekM4F7hXWyabWav2hInxvMr
iwj42hddU4NhFE9lyYJaGh1Azc8urOT/jjZ45pGMaTGNfDHzjCq96+YsOl9y
3IWcwrtJetzJKJZWkVHhb1Xy25YKRCJACnz1J0ky3R5fTb0dJpbt6Kw/txEs
ke6XJVTavXqX+unLVRpNDuPHwjdrQkeym9WnT/WOGyiFEJceYQ+h8/snbQJE
QL21rF7VyIzb3oWp6tei09IetPRcYXruJ0su9+3APSnL0kzd4OMokz84/BkX
Q97xHSnejrE6VdL0QnF9d6OqYEjlpLOI2TZNRV1QQnjtBbZyVQTh2awCcJ1v
si76VoSWWmGfyX9TaDk39z5nD2nDIoLP6leAOkNiVpD+18/0lNWM/eyK125d
1KPwVzzsqQsZ7FNN7JHEvBn+SWPsY3ZVRPSi75eICh+NUKF/8GgUrQ1yznn6
dwq0uVGafLbI9mhsmWUb102rwyIxnqLAjgKLbTdEEG+YFKWgtztNvSMntBdY
eYkvQvEkDReMmIZWtD8S1Tn4xd11htwqW6T+zNJ2Et1xFQ+PVCef2auEEVXE
S9uzHKSqMqY4igwIOCgcxgTbetcKCqwCp2SDvHU6B7jkOKGEhhVIdP6DUyLz
NRV8YFo+a7w4EyB83Yx2Nq9BpsJBrUek4nHPUE9bHiyoowTpD0py0U83Qnt6
K6b0ntX8ekiiQVv+nycvp2M5P2zLyJaT5xcIiQNKiK4YxTLy9yHk/rYt//nv
ZOYxAzdJDQoJTIBVEdkpglmrehEIGJuI4FdllsgMCUMuaSKT95uqu0Xrqo/S
DcTKGFFjkUhEavksUEKzbNbnSJm25VagqEryginzW9odQ51avShhawDUzmrm
BYqXLAfmoJL2PV//V7Fe7S2Z7Y1TJQZiG5xLt0lFjNjnuj+ZyGL52ngRNbac
kQc6WFPe+uLOuhaWVQ7y1/gCsSyPTWvpcxfNWpOoB+uzWJM9ZOVavB7C8IaP
qYs9cqDS6jgvCUQQ48xtT6hkCwraGwdXN5s52d9My1I0HasEQfJZoRzd5MBA
EvxZVdAsCjPpmjR8Z+bnNzAjh0JXHUATeKIt1R0FVdsWKk4ywnarpkgzCLDS
ooNthxdAftDJP4tnR/oOwbKes7Fq+z4TDqU1iHN6/b73OQNYoy6tTcoV++UT
Cp4cHKXen7BdAYfnqTWwJ4HewjnnnIuiznn7uVJecEFmi8DBvtZ8SJJS+34t
IOkPzkoUOMROlIkMiRjew1zvVgs8eec9zF8EGPGnRZgHaUQbcu5T5WCsKweI
1eN0YaW0pHf77mB0cGSgAwXNn21nik8H6fH4aHHrmGoQWVRglylq5QQdN9Ut
ZCLTqZyu+h7slrGnhnJwjMT3OA+wgnw+Bgndj5aAPeYXIBPj8PSuwxLUETJV
aLy9ugp9MwNwLlesnK3DPmmwVJHTsGFXcPaYRRfKq4xJwNeNF0LTZXPeoGoo
ddpuYwB21hUIKVlzFwK1MoxSeG+n2KAo2XquDAQHwa70Y4pMS/GhlKoC/xkd
fjZuT6GGmTOaiMU/M8elGaR67b3UV2J/I+Ls5crotWPfF122AFhmqD9Nlvck
ztbrNtpOoNAFS32glhDrv66QpUu2Si8FxPAopJCspGzO0o8hKosTEuenpbP+
sJo8ddt4+xV3WiWQqUI3KugWlOp+is9z0pk0/44o/H3y0RJwD4rJ5DKsymu5
U8JNDya5gofymxj6csx7RAIN/2e8SpIYupKr03bRExrIjXQXiPDAndgBSIwy
CetUU5eAAkK6Kmf7cm4pBIauh1X9GybUIetQ9AlAaSDQ3fBjHiNHQYjUHY88
L4glSUvEYT3+5rmjBtVwBMY9FnWKhCwF3vmzm6N5o7YsEkYUK0s5Mxe/qaI9
bacFK+wLU2aF5Q9P5obgTrIU4lo65XI7YXJ+m2VvXNJT4ugQ5seveJW6x0Hc
VBzthkUMll/hlsrjx0rGYOpartLypg+FM9tp89gzfi8PyXG0ue9z6a+lMNQH
osCd96bfaG9LaUyINa3D/vQBWA7mBgZdFEY8Uy8D/jfZdXfrgyoqjZuFpeIK
kw71r/ubTl3GMrzAFHQkjdxageKsRhUO89RIqhhHpr23nW0LUZwZ7sSbyS3A
tJMaUuwUjHnfzDBirTbaQyqNP1f86zKzQIhZWdwr0/M5pVEbfbf4bqzAhVAZ
eqNxQG4H5BWvVy3K79eJGQcHzwfTfK0ipCzNdfLm7/VI6GFU6ydThGil7/xA
i1bTKekcShTmibt/k9bXqSiT8wg00RVsNzIry2ozmDk6Ye3AtVIib7ajwIO7
Sn8okQ8Omk2ZzgazDvBMS+do2s4Br/GAIqo3WfgYjZ6lkX0SRbIHkX9Kekuh
/IrWfLzHIw4QIVlXcR/2NeKtPtp4WHx4EDY2vqYg6qyvm18hvNWjsY5eMl4U
bE/o17oAe3u37UT8kGJe0I1lttUU6LZN4zAgdxeEUrSYj2KGUueCz2iXaKhM
h8oOplhJIBBhWgBL0vbLzpEfl/YAakb3NeXIn9rY989XSuG62KTdwCY+8+PS
4+ebWqSyCtuoyCgKfbNavNaJIwmUd30u/Gep024mGw+siEM+LdXsKP6prhh8
nfHGC2ZsuQS937k2MLRJwS2yeB1pbpqn9YDtp+EkRZYCTyoxgyS+G/QPrYul
zH3h+pOMAGW8d4QRXzCzLlPmS1hH0amFyTcxlF+VwTQBhlvsZF8zYXsOFCKm
ZkiJL03Efm5XdMvqLSi0jSiRoSaB0D/ShUidoBWdJH8+ac+ByveAsbjmoQiv
0i1D4s6vxvktKQhbQ9MCjMlPT5qvOvyGYXFalPJqzRzoVFLD3yeFdEQxqmp7
Ff6kAV1lVUf243cZPfA9iEf0WTZIYYD0OrJKUQLW4XQqC+0vMCrXoS8yupuF
Bwvl1bRRKASSUCA+l9s2homU2oCLAq6WNqdszqlMk4fQxUrHWHQsdgwuRwMv
Z3jf/CrEbXhDxV+PAn6BsIFKwiYZ7mnVaIdJFIczGGXrq6bHMfQ1G0cs3lgM
5Vkbqm44xk+Dmoylp0ms8ktdjv5D8IsPUorWf97vHNkZVRRGSy2qfkc06s+S
sj378//sFGUyccWmzc1erKBisC+CcDL58zbBz+4iXWQD3U+O0OKYtfUp63JF
HnNp7H6d7Cfg1L5KCUlh207SVGH3rHvL36pAMOrzp2UiGQg31M00X4TZ+C3S
JMI2JXbIaVWzk1WZ584opP0TsCrYpXwbX1yuHG/ekm3We6w7jVcXz+OlCOTY
mAtuSBYkvqz57DNCSVh1n5NxAT1tB+FqzVXfT9f/4kbg5xrSugLS7Hifyttp
85fBbICkqNE43OmHlhVsE6Mb7bQmOvBaup5TkuTtHvxBuA1lNETXDisRRPzu
abEvJao/fjFbSaTekSaykYsYeLRk7wKbqBl19zu6Ay4fPaLEPUOaAXUkCQjq
zcqH6grsIDKQGPawHFil23zasmcnkXHhu/LLthjF+VDcNO6/XvEmx1yXkiF5
a/7T1XmOKK6elySeiDIgPq6KEpSkaYV8xrbEkr6Pxa/wJN91/TaHy0l49SOF
tew3mshUW/dJMHa+IOqZhMjScMivGsM7jTXYgcks9XN6r4hpAAcZCtjreztg
NuJpaNr5sOiGsBuqAHE7zkBg8Cu1YDCc/vpcKE7cVfYXkn826KqelEknO7KS
Y46M1758og2s+6qzfoPMPYwaL9SqHQBzE3oF1YInJtEdkkPYIBrnvfss6il9
VkqBhPxjeRwVZnF9PE2A7fFSaCWOcQMZ+FPcOSg6ipI2+T60P5cCo3vFwlTm
H1X1Xf6lX9HwIWmuK+syFdqBeTIVhXnDL/Q3MV/yoXiWQj/pCqYJ0queXY/c
b9YcOcsR+bfRJBBHBWEU80X0DZP7kAEuUlQ+EsOAr8Vl9Wjf6XhnwTffArNz
TrJAEhwvRBr0qjURBV73Ve+ryu70dlNkXXQXf4UcjeZIF+CEVQFdlrNu8rt/
VQiPh5ivWr0ET7xS8eqsJTTPqG6MaKyH4cw9B/HX6tg70EOYD81b3Bkaa7yU
8OrlKssWxDdpYIzGGDkP+sOPCQyT+IH57oZwykAUh2ex6z/Mq0cYwV+6B44y
MmQFCQUPIQhorSFig78H7V+mv947dA4+H/6RfducAFbMACx3uUvjYhlsYbuO
4BNOxMq6WdBvkl4Kns8nJK+wYPNeF4MFGRdxDyA6/6+gg8ak2mNoF1faUCYX
mkztBlCOUc9qgrXV8WiT8au1pmwlqgu6Hy/AgE7cQ+8agA8xv3nIWU+Tkzai
D5LQUm1EShRc8c6W2fRhl1yXpE5tdG3nCkf2qJe91PCV8X7rGIRwoUt9YbIk
QIWaK+mcypxkPKCnheATxQKZPS21Cn2oVIssKNc2fLe7TNjtqWTgIQOwuOBM
7GmFQotVe+Q7IoJh+eBFhBKdTzuoiINrKMAvW0zu73UK2CZAeqSL6vY3i8A1
4fMOi6bsQn8xDHsH9HMz0ADeh7VA8KpBpnfa/It34jUT7Nrr6Q1W2aXD3NN3
ATMZfutxTnI2eP7qhGZTzvgi7WwZyh1t6cYLA5I05UfVBC/XtPglCJQkvWrn
vet3dg2jQHz4cUw0+Ek6fyLV4192FsfRVla4eJR81t5id3585h8WXUvvqpj+
55HGyoNmtF92ZEdDIu81GNmQfoWljVpCh+s6fHybgXE3lhgn90HRyLpF1xb/
LALXA4IdJnfS6Fj6CpAq9A45sYv4FJ/yggeDvYWZL4WQSm4AMdzszOTTvACS
a1wS/XOvQi2O6HZl/U8zaUSA6fLQgFfkHfvn7UScIQyx1F5ztM+KuA6tNwSO
bR7spFTOs5ICNMcxdT4ztfihdc1haore158U3N6ygBOymvHrslC5LPFCNowr
PNAPBo2ki1+t4oUc7RAUV4SUhscPPs05Hm9mct6bzbBdL4luKMjpqIx4bNIn
rVbhx6ZieDT1DO3ju+Hdlw4LYKYuU5zXMTTdOsdlv4LOoWK/mTjWIQ4IFTmp
67/ChQWYhe5mfz1DJg7fGyYU3SrelAi5xX658rLUzdXoxIKdyXnHwdRqmz1i
btOAFnzWjZFv0uFyYqjbb88GqWbJ4cx2ttN7urpzsk+RNAppmO+FvBgfTVEc
WBT8EzDFvk3sXU4+gmvGPrDBZBMlJkSocp1lAHEVnHR/EKv0B7/t3/IUFF9O
HBUjateCUj9KcA0qQ4s370eHZRFDWtAHe+fs4SDAUkiFDmQqgnjurmlk7cZ9
gKjdN6+v2eOxn2q/Eqk1RLzf2Fu1V5QasU9lkPjeUdpCQSeRIcpRWHv/UZk3
yvxDlMW/570Q8dyBaOY6mdCUrpJzSuBXWRl5JVYC/7WayT7vdbD9vsBkP8WY
jmYpEgdgScZV6Fmf2K5mBhrA2ApzqmEGXt9Xx7Dg6zxsTi28iFKDD/BVg6nt
d3Ddirp3YBPbK2WLC5VetmvoB8XNJkLmXgXNnKyxrJrkppherKAUqnF+CGBL
ZMPb98G2Aps+/w20m2StwFxlV6/ynoesmKAdvJUKqADqxf+4jbsK+lyBrEIx
FG5UdRMAGGi/hXrqSk1k7DJ0q+k+aTu6fTMrvZKfv1jReXpToMuJJNgLKWtq
zVliGS+KYRRnzY58Ra0R73flrAXS0F45BNW1UcAU4CIt+1txUa/uroVmnOfD
e4K/skrKyU7fe6xsX9vb6nb2oUVByFb3IMxB9IZaqyeh6HoYB0EcjXW9dvZX
WYAq5Us5A/giHn87wIRR47SU2kTDFSIksVV/Lr9sb32y08oX/vfLbZhFsPRy
Uxcuhu6oG88Oo8y2lPGgECbBshGwrYJEMvHqq/pIzDD7s29rT0+WLZBt6bUq
iBrYFS93B/IBlHdp8BKQ/c5O2ORMF5uLw4ap3SSvGx5589srKInwLHd8M7ed
IPnHXPYU7pgzFOM6OrsrBUQntx2U94KUwaoatCckuwSgnOz7JzgJI+64NFd7
tiG20Xm9jCaFedUWwgCExLjnp45+QGYIiF1PHi6nZSM5lTcUSlK7TOQAQxvF
q7Uyet32FP74y/JF2E20/al5HVH/eXXao9Y9zqolTlQrlDbulQKsLZdlYuP2
62rBIXOqNbtohefVNXrvGCNSb9UDklGb3u0C+8BWFdBfIrVdTmQiN6J3CiVx
Xkcib6bFM5ZkvBCv1nhhRPPfT9rRbimVP9PdXY/i+yr9KGQGsrgZm32GzWcm
sfiMp5gMOV4xKIeH7B8GmtWg+eXL784lDZ2DAhky/N79t/WTnhSKtqKFi1SP
c5xtVcbg7KoWSGKpOvWAvtzeqktYmmD+XpXfDX4PcX4lh+rjHUfB2cICAki6
4wEh3DKMT8rWR4UB7Mn0jICWwNk+UWJPOXgHUkRVtapQ5Gj/x3qnYK+euqJf
DyI4vRylIkaSFfK9FMFvzbAqTd3qT6apwkh9ASXKSjxEtKRW4phqcCTGXohU
y1BKRe5DVZKsdZ+bZKzk3ZmFxEJkv4Rx7KWbGbbMym70gO5E1Eu+QwdebeGM
bbVHUtJMbiLkXGTjKjbYCje9dFkkW7Rz1l2kOE1OrO2sbCiAQfMhXjWENKhI
V1x36yJOdTBQY8tSWzR5N9ErWgbjBMlP2Ix5Y5im9MZjC2dAuLrrUPU0C5i1
XHfozV8IIErEU2ut75dqWB1KaBArn1JmGRBPhS6khyjPwkjGlCODUQOlJkEf
y+mwkU05lsNxoTkqf1egq+qecyCUnRqMqA/gf8C0Vf5tA2HZbr35/vQwIq+P
WDnhVd3Lx5jDTNDWOjMRpSNkrsgb2K5lSetdHrLYk/046rZ3Y1khk5UGPDe2
KYcoCjfnZekp1PQjjI5JLinP7misSP/sQwMxx5iqdmsGvNtZLw7yIggeSmZB
aCWt2+MQU+lSf0eNEmbX49ewMvfdE7a374Zchf7EmUd25uBrwE3QNAGqIJO2
kQksjcrAaq/vWjwJKlJw3INfZEj1QtHpzY8RhS3b29lkyKTmQE8cEtU2hUx5
NpH6RC8SwN2auXqTtbaQx9e8YEFZoZ/cU3sIAjsMdyPX7sM1oIag6YgS6492
sMKFPzb3cNQBPudrrp7eODJqJr07eUiyLPUqJy5WPxBQjxNTW/NH6prfJUNJ
ZmpEQ0U+DW0h9ur9sYKJ96q7lpSm4SjcpEsE3HMXtEM8DfDguI/n2UgTiit7
Lc08oVI8a82Fxq0JaXG3G1zyARd7fvatuiGDGYgNg4axEVJA9E0vDqhFKR2Z
Yc5LJqq7KWAMMnJ4Dr9dIl/eIjHIaPpkKHkeRkCnjSbHPn+HxjvEY1lc9S9S
mAVPXbPLzXIAcjD8C7yumQoQS2KJ/oxBpdTSC8Jn0udJbN3RcWdxjvxCHuS9
AHOveBe2QUXxZfaCmxVlVOFuUEVL0rTCiIPWF0dUi7MoE1+pwCQ4jMtsm3Ih
N3lbt1ipznlc+C0qeo+IFGUwEcN2J/8clu2txy0pQZA37YvfhEJkpcxGQNFn
8Wx0gRiGnp5cVFD/g54MeY6njLawzpFcGjg8XU/bc54lcj6Gv0DGPM4mCQ3F
YRMEssnZ6zAeZwksUwe8CAwhapjHcF5IY90/1FA3ZyChughzjrdGL3sjeULz
dEZAHAjtaLNHh7EmXFrfVLHvxB1ffmriIrrvWqEsRqb7I9UcESe5nQP5eJ7B
NVtSIG6HvTm+3/9ZUlGAVslodVPL6Bnh6Sqr/M91kD76ovVQh5B5rD5J2jx0
UGlZAUK9Qx2yRwfGodCNu435Fa+8Ln7d8w5IvguJMNNFwyungI/WNAPfyWKN
asDRI+qnwgeJeVWU7B+LyO6MeKfE5HCbQExTT1cYx/8OM507R8W9nY/kZU86
473W9syiSHJSBscA3zikbPKz6JrqwmRFLoWypXSJlltZpqZ1ibsj7vWlYMff
9YuvLmBvpcBgnjoiECVY8M4CO9v03GY6z7JXUvl8KCHndDwOe8cfXV4Yh0Sm
moVvQQ9pSNs9OP7aF5i+9CX98ZX+yszTidSbZJJJooTM5O2QMVmOOJjKJ7bU
JR4gRG2vx6g1pEok3Dqhipz6TFiubd8D8gYaqkdfcIpeN53y6nmpl6cd634M
pLsPRJaxbIGkhIBybUHr5k7cfDzr2x+o0alz0VYosT4MWbNdus+CgRVRNy4x
yq743x9nvSX2dCjvVxmwgJBisZkPrjcGbYrNjGLhJ0Ktj1Q1Q9QgWwYxvg6c
1oOoZainLQbGtQks9+ZUoPOP0IVIVdSfwAOsyGvddIMygK6S3c8hjmeG0u35
I1asMPdvZrsA+GzOztgMYqj4YRhwAEgXSSbw4WXeOOXxcX0SiWggt+SDZ0gL
XJCVqmmx1y+Ahoa/3UUn4pDqaKPUDbZ1ViY8E5OynygS7c7+Iz2j+8BscZvu
dZg3O7P/rv3VGReOiUVM2dJU2eZ32vzIO4bUeE0P1jCmUPQ2z+Sf5wEoTRlq
I8RTfZQwtGuT28WPuJ8lNMBiC0RFQB4f2XLJ06BF6sVlm6mj1oeGZe357D2a
JghIEopZrptpahfK9ZZrq6d4xXpl6as0mHDm9azZZvQozYCRdR8xDgkHBwPe
yxbVBu4GUlp0IvhEoXcgfHTEu8T4iFXX4qUbW8kljapukXmrv/gs9m7LHer7
7LsqYmbmL1gkY4zelxydR4ETZ6z5bf7FHY1kRfuEPH7QAYbVJO/Tu+XAZIYB
jmYl5ZdEtknJidzlYDeGhM6jNqOX5AJWYdk2Jgd6xWB1JP86d8l40N8rqmoX
VPr3mve+4BdbTrh0Gmra0EBECxLgFP9X39+yYb5Jw4qX2r0T76Sxx4f7+s5A
YiSdj1hhtki817xyHqqkg5nq/+ubMTOmpDvrmndcPjJOcRjB1ZsEaZLc3ukr
fF13iYeCdbiuRlQhx5RmFAhISKL34a7DrYvMYyrORWd8nJlwMbvp46tiVUO+
VAwHhenUX6oEvHUAoiwJdn7HPD3KYrgIxGJmvesOlnjrD/KoWPzkQI/ob/b0
hUfWqwKBv6Urxwxs8shNjbMMP7n0vchijVhN8hb9LyOurfgjk8NyvbqOBpqQ
Ps8UneddVVYAi+71RLNZYgeC4BvE55KRPvSMt6cMMexm9xGqYLTtvjr7CVQY
5u6SCAZUc9W85Y2Geybnbe9j00lu+wp682Dfr3jU50apGyfL0tqrFw/3zBAU
qxJ/63IOSFIdDHBqxdtcyGQHGtVqWHZKTCNy9Lh18K6ySAYvzdNMQShtuQYC
WaXpgyuF4zr5VNgbk/YpxL2phzHaG7ssyrW0U4xul+1xUoSrEjxIdKk7MRmk
PSeV+7IFiIJUTl8awcS+7ob+KkvFC78t99O3DalCTrdteDe9KDTafnvD+6V7
AgOcFVi7f+2Fp0r/fyyQg3Ia8z/QKRceD+5Ag77Y8ZV+lxaJrzRcj5kb+Pdb
TaQ6zZ5pz5o8dniFK1X9PHv5CiEL1SqrPA1/7q2OmG4cM4Kd3vansaWve1Cj
VBzAackEwPUdvjCZbA6/SBrheCiVwsa1sJPbA7/AgxJ2/vjleT8GRu1BrZKI
NSfwlKgTx4XU16rO+pcaixD267RfT3N4YLnZIScZjxHy0EaFALPFOYTH/sIY
h3UZMK7AX5FWUpJfuPhUwbWQvR4wP4NZQdvV9HGABS5HR0lVOAlU2RX9MCpe
rg0KAJg7wok8lKsV4DcAE5i/FT/YCf66R1nmclNKc6URWWdQ+NYgmx+swvcb
xP0Dq7epR3m9gD6N6AyQUr78eh6oOuI0uuelx0LeViSBr8Ly6xy9VLDmsk5E
wuzN1/WsLxuvHTH+XwOlCxJ/0DHFhIBAb6KVtn1pkzkWxfnlm0k+hpUHN5+f
/tIAnib+Qnux+8tx7mmw5T5RGqATF4yFGNARQ0LDZ6rwOFBZInRkYWExTsSK
vtJyPz3yvEmTPoBP56uGnY0f/CpiKFxGMzg/Gl0A0G9ZSOrGPbkG5i7NCA3P
sy8a7yb8oeqORpG+8JCBpSTWysmaT16/bK5B4Tn1CDBBH2jPW1vJ0zzEHjus
135zbo2nQqdr9tOiJLewaMkKNhGgHC7RyssdtQw5A+upwOpzQNAKlkRlgpmm
/hJfqZO0AkV4guAZRd5tMo6GiktqbieNsYGaHJMJZ7lVcukKMuKb5tBPYK7Z
uaUoT+fOoEhOFxeunpOPCe7NTmpZ6F5VT3eUJRmgr9D9oqyxp6dbVo747xcn
kvcqf0uJo1B3c3WqFpnv3zXFKq/SlRmUzSGp27YG28CJ/n3/vWZapuoMsB/V
DBSTn69RGFYCW0X2igwPUOPHv8xRTe3eATmDJFTznSXixjIqCn2dg06nnLuI
xx2u2FgRv6WOzrKClvsTXOAZZOiRGkEMeLsYrr1ULEO7N8WBPogtpywv4r6O
fyXLjgn0lQ9SxACTsgQERJONeZUql/9Utz7y0bhhD1/OW6RebJh7Et3Nv1Pa
N8xtynAiHomeyEuY5C8lVj5JcOxflE0sPyYyG8yBc3HgryGXw9iFI0oPUKLG
5lx7QG19eU1msbHUY1M2f1TMMN1m79zBpvwJgnKybY0g4os8WLhEcctoTdVP
Gs22j0nFASFzpndzTdrZZyrCuJ/sT52hk0AZrzR4pgEyGbRUyOvHtMSh8mVQ
9fVvjaTL49kebi2t6mJut1FHspyvpTFCLatxnWl/tolPvrkT2FVSdqIcDpTe
8Q4vFG1d4Wxz2/gnVrGEBJRL4llkPGXJmvy+73g/xdDrgCkGDVJ4jkT8YHOe
3jiOjmoKx6S2rg+Upnf8EDTp2efPjL+zg49ccCEEt06XC6R/XWaZPcyNZMwM
10WLsLS7OnCBW5gM97yLj0Aee2WAnj7UhAwm+uwci+ny60dSqFvsXyVr8gvD
zlQa9LBz83Zu9an+MaIYpY3uM1vSRBwCvQ+ifsQozumXbNiMMVPoMhc3FXXU
fXJ5ayzV1SgCmWo0x8DjVuQKOPIPxJGY3r1TGowsKC2GzGCbFw42YErqgIlT
s7VCP9Zv9o4dTwymTCupxaqNNJb+29ip+Auw4arUk9c5Io8AtH0DcQ2lyIkM
vcRC5pVI6MLSiecLT2ixD2ebe3J/JJCj+6Zuu5bXFWovMU+QrXfW/yVUYysc
1x2XhiyZA3oEeEac65Wp1pLRNMbt3GgtCkQmiVGix+bGrzMGZXVFGA1s7ujy
OBlRnSQ636hSiAWFQJmri4MgaAm1IfmnsMiYE7/ymeS/LAPlYHTp4VJLaNnZ
iKUWB901HzDxnTY9+9m9hjc4abNuRWFWpmFipy6C8OWOIu+nDyHXqV/2upGa
HakMkowQJj2CG+KAjxDf3HJwNQvuYlvVYabWHcwd9YaXCBR5j7UMlxHXdQwl
QqMoy4DzwRiIeKiLq1zHuJ65xvbxiirHb3VkDg5FHvosAeX1BWbko3BL/dyL
nxEGqfWDn4sCWhjjKXz277w/iYAmFOk+XS+gr3Aiauw6mJpTOQtpYxRFFhqT
xuac+1xNoM4c294xT1bob87IVooy77ccqH01rlzRZH9rMlSpSVy9b9KXaGCO
5t7oRNBgaKC9hdOWdj+W+KbgKMGwEVhkpnlxNjafm7QWCt9nQqDKY/InD6xp
areexpNKKI8LNbjUtg73YhH0LzOuY13JfQdKbxKMBPvON1HX5S9gaLF3WPGj
+p08vcvGkWoLqhC/wVl/mEgd2b6vRvYi/KIkm4Mj+n60UsmWDMP1UyFJFsiP
8+TkV4iL/t7a71xf7dxJbUwP4ySTq9sH81fXNysfC5oq2WlRk/84NGihfFkb
aQBOSFjsgg3vOkgd2cW4Vf5HN7OmxmqsNdtkDIP5/c+TidzHkO7fID3ptgD2
WUWNF/9l3zmiik3KUxnWYt9b/1s4j3uZRgmEZvAZCgpnopO20dEBv8Q2DUHN
ofG6vBewxyVkmXdo5pAglorN80yHWakGTp9hp+BLbwcNNzG9MidL4jxtcSBv
8OpKHzgD2OdUfWOsyIExDWw8/QXvRRyyKBJSwCISS2T2ba4q9rKVz77qYFMS
fiUvY+pD/3hmcoZVGFMMvk09ZJ2YOVfB2cQPRxClnNxhLyaWUYgIjL2UdoKl
sqfc2qgUkuvKVL8C/4+vq3JDSjI/aUyi1S9Tlu+aHtADgDUN0QBCvVMY4lbC
h4tQ1VymbdVpXHLrsICe+2/vC5zGC4DbRtLNkrnqdqjYO1oGFaLb5rCqA43O
j/DD2zzi/tUZC2OumWRjmM22+E1aw9J6xpuYzIYkV+SBZZ6KwQoEP+PZDgrp
rYASdvXezVk7M3bQtVLd/5mZoJncID0AGrq1y08Pq/W1eH3zdH4yR0UTlKg7
D7yzTIH5/iRAWi1hNPGcA+CvKq99NT4NlqfcmjSjkOPtJvsCTNRvALklDp8d
+p4jpSC2rwBjp6e+zFyudoVTQHFHI56t+28vHhrJTuy30022ZMzGxSgmIbiC
zLYRqVSKsClyVTtEaKMIkiO8HaLGlnloN9IgH4bKlh74otGTY32Eu4e0mSwE
qL2bIo281/nEqek9LoB1gPJx8Ti450Dp4EQnqMoE/AAmfql0d35fN2yHOcXY
yD4dPQU7WU4scAR8cqvRB+dNUK+0jspaz+A4LqOFDhBainb8/ouaq8ToMaUR
hwSpn22qhiPUO1pOgXeVgeisqvlc6nPhXID6bweb+lRmWn4SNmZZYNtEsv9t
TuCrmmi6pKrjgm+auGEKMsLrUJ0c1oKnJmEXlYLQfb1pwLjWFN0J2f8oIFJD
T0N7R997P2dICIh/r0zHV5JZFroFiBdAFFdihPdK2ahyyWwUrSrolXyvG2RE
w6AF5g8Cjc8jr6OnAwIxy6g7Z+LOX3TdRAsDM8wgKJ1TD8xaD6dA020LcsDl
JkALxkUtwQTx63HzMJkeb6rkDZON41KDoKFP5qMit2LbBruWZ+buGc4z9m6M
/u+HiJua+V8Eyy0RaqA3wVJN9SNKg+2mdTOkPqoaY/fl6mW9SpD96O4vQZ/D
BNbm+m2I4WjWrE7J0+kLxuurJNlKbuNaS7j85DWeu68kAHgM58llxYvTGYmh
3/qdni62dCxUPyquSWRCXX4aHY32vpsrzBVmuzLF+JRe4E7Lr2Pq6pGluFfu
XFEoQB+GpUQYZfOG9AeH8z/f8kiBDzDIJjlyprEvIsNSjD3AG4U42Oqvp/0U
RNHlIvmskeQq6b/L/IkFro4ySrCrYwI8eP0VKZmlaLYDlP8l1Ur0jLVLWh5A
WpmQnIuPYjNn8NN+H5gqHloRvQIJjc16E6w8BUaGKDhw+lYQ8j2MVSKVOIrW
eHd5pcsfUmqynNEy+iKO2xwaO/9+1eOaoziwfy+8sYXOZ1BPznmTvARXGhPi
KMbzEGznIw6sgzuLC97uX0feZkxhmkC4yGaVI/zxlJHOyo75c0sMnyrae/0x
vLFc/uV07H0v4REOHhyFCyb+vhGNUQvKXr4SXr8idJNL4vBZhpiv6DnlJHNf
o69fEJURO6gY9mIehxNbtCncM5DrJligrTIgE78cdWqWtkSy59MCSkGa0qlf
zH/0V0G89bGFoxEn6I5Y0LnBRIfwSgpjtF56T/A9xhlMdk48E+8E9gJJUIDD
BPGpwGW0RFUdYo4u50ZO8clUqTtY2JQ8zC8flycigm1TNXhKybUZXEms2jAY
nPJdS6jRw99vINLgV/u1JdN0lunINHKmboNr9ctlbMucAAvqcF9M2dUBAF/S
sH823pUlsbbP62xtRG6Pa91JDBfNJ0FGoKUpa73hJcPXdBr15SdmHJcS8L6R
dUmljAwuySPSM2d0eoTdYgfzOZvQ1jONjebuEUDAwSEW64/7gi3ggFEjSEna
TClToopv4Oo7nbxiLv+BdnohkikrqIHN6uUzexe6m1bXtj6OL5mhlAJdDY01
wg6Ni47DeHIbwWB0zjIdB8gBcrbGKkpJNbSLmU8Sz3++rrMeuyYGPpfdI3Hy
92VkRqhtttpzzup3erAdq2L9ropA5dm46Yoq9vUe63j4K13WaOkOHGiAHMXp
9K/S6Tue5pe34J/f8R2WUM7mY90ePqBVFQlDaj4EZhtciy7PdsBcAdEYGak4
WrN+OxY5pvm6AbQjOaWhQR7WFuyjoiReLzkYjJqYgWqE5BFxxMpXaUnlZwxg
SnPP32bwYG5/b962TbFna31WHMj8yZip366NdpF7mL5J8jmIOfY5Z7ow5ZN4
X2uOMCyzaTsKfdVq0DC7g7wI0V8Aj0rXzwxXTOTOPSrgsY0761BJ4+jsz9OL
NM+gwS//h8/kNjal8ZeYG+l2Iy6frcq3Xtw8Y68YVKUNn6Ug6qWbMlRG/caA
1sLudkrsuijOl48LqZllEIqAC/zJCWopVwT+qQRPpgcfszetKg1HAa/zFR+6
RmmdfMtvZRQka+0oQCQivSro/GGqLvN+/gutJSGYteVIBv3f99CGLc9+u5U6
7QS+3rH1nIQKTpScf+Xk3nCvBkvNflDk1ouKQx/NWrpQm67VORCFbGGCrpc3
Tgfjk9pIX4HK1/j1G/JFiPZ3UOYFE/JEh8a5ykyYkFX8wzDOkl3bK3Gbyjmk
5oiB40POE01Rp0hCFROSlXIZHSELDxXA8z4qTP4VupFLJUI+W1CbO/OvmC+9
awNHema+0mXNtu6XZ7w+Z2RIXlSVCzHF/80qzIpQQvIgTBiLjaLhxivs/SsR
08HG/+C4Ovvsmaffk4AnFMw8DS17yfw8eTtnuexjSc4cZAq2GZZdVtTEHJ5b
YEf31KNQXS34OwTxaV+SoyHNlRnPVIAdscSDfyajVrs24ajO2CL1RYUrxG3R
PrbxOn4bufFxrvTrvEGEDRIJe0lrJl/49XG/Y6NVFxLuUa6nIcyCo+QoX3kj
e6LMEWfP2X0fEmcZf9kUr2SSiPkTRi0ADNYKsC+35wGri6zrVkFL/mkZj3B0
ieNDkm1e+mN6h82g1pU/OYnwWMDP1p7VZmRdoRetSgTKX+PD7ta2nnnFXyGC
MbtCR9PuccpfjEn+UWXyLXJWsAyQdlQXFMqzWJx6WGNtFSHpB5Ae90KS+lgi
ydFlJC/AYy4RXLtcNFoICXIJ/Cnb1rKlK/SOgaZEqzCoZPgwExSDoDSwm0iv
uhCTvpaEaslbZ9aYZs31cms2bAIY871CHKHD9ZZOecExFJUfPGvA3m9vmVW7
qlE2gvRXh6pG3dgCiGFl3dgdGyR5/wCCod9ZMdba0AmfRMuM1vVCXYqFS60/
onZ3l/lV4IZQcbYRkx9LRjCxc27uMGHdJTj7hBjENoLuK87glBNrZoA03kY9
w10cLRrc6k+mX5SB81qOr6mz19EBrjLfUTrYwATzxerLIOPQkS+7kGIYkJs1
Iz+K5r8jP0p9lfdbJRXtKUIBsyVs9iH6ekD+wgrzyeBdNlGrlG1E9mI3rUEm
nu+NhCLBC2qBDx3XSLTXZKE+yZkj8dUD0P3TSIjB1+2MPdGA9f7eK9K8K+4G
mae0GcSCVolEa1fWCdkFdGsyO1CT07sADKpaCmxjqv1x4hId8ipONXMIq+NS
gMY6UoYau/e4ZOGkgP4UkEDnvDZoGxW2yOxog3Tq1vLJ2C8H6gVJfkJ4lfDF
bgP/YHQ2pXMk7yB3v4ENqMT2tjixntgGupM2YXpitak+f/ZW6clE4HOdLD2t
cqMVqOObHmMaDAlQBNM5SWyUH4CLT0xfJVYfXmBZ6bRq+ebiBpA5LKDPTOji
wiZnaeNVlCEGqgS1UM4CBtYGbQ0G7kzIf5Tn2VsvdbxiBNPU1CiEvb8C4jjd
IHgnPhBjjhIUeXXqbgSe1Orfurcf5VjKg1kHlD7XJX5AUgDFzGukjor6M4E/
flsT7XcKckElAQPjlqHPzuz3JT887mP8K01+uNgP89NwovWa+tt5NmvOs2A+
tBEHBRPqVUDCF1ldUs7Yh0H6L1Zp2Ta38Mdm0rYxoPZzoO/rzlocKYqk+m4S
EjMHkowoglPNIrRQ8t0TGwlByk4Jy9NK9Mg/2J2xjUr2oVbM0/hyB4MAYPFk
rWx5Y5HOf7IdJ+SyitCQ/R7QPNqQ489Yqcm9+x/XkEhAqsnUYtLh58kumoMA
SXCn6fwu3SLwodliuI3V42oaPry9WY6kCittjmlH4wjrVzJacZy0XL3IXqw4
jy4du68H6QYzRTqpz0iwZCaPqTVJY1LeZWCzl7daw9o1a/mRMnP6+ab3b2mJ
mhDInUto1FCELsKuuvoptnUEcZc+VkHhLy0iakhrYsc9QRCmfVNpE6oBj1qH
j9H1QDJXff8H5Yd3btcZi/SgCPnxMu+PIammAUmv0uhm3QgPbv5Q+u+KRGrJ
7cxIlpCIIMhW0NG3cOTA5i0uMTO6aw4vzRpZN7tvA/7Wo28YV2ij2SyRx15/
AHo/L0kN8fcAExt56np7NEJSVNI3YvU8SqusFJw/WUUUf7Tnj7q6uHxJ0tTf
cOPQu9tc3KQmlaQRl7cHLnUmgpKWhvBgCS2Sn6nx/lGCW7VFip81Iacym54/
b9IZitEwCzP8kIiXyWpdN7cAoBdtygoX5laUfEm8xvwQyZtHs76Tpjb2qiQm
nIJvUxwnga53F8qf0frPgmWJR0qp8DVEI+5kHuxOunHHclB36Ev/fX+9o0bN
vZTaIvlDkVzqHZb+k5GniBo5opbTS2d8qel8PoHCs9DAA7PyVasnh6WvGvb8
gqAqDIo+JrhAE1sBWsnxcs8Ol8q0wKqHlTh1YI5OE+iFGFsll9hVlBfxYoEw
hqpKuPlyeyZkn0zxJolcdgPRE4i/DftPIRDrOZJcbCBxh9oyDi7LMVRCxg+F
IqIzmC4D3YGxqeuk1Ytb9By06TK3Du1JZOI1uYy8GChtQKb54rwyEINqXJYi
0X+gDpgTAy/10te+kVoada2yTVT+6GCFJSmMyF+UZmHutcLSFfqruYSjHh7A
gY/emUI9JXX/kHytQzrV5g/6+5jfFi/BDheVYu7BGfYsZHh4E1oP/hhOX6R2
LcmCqIjx7XNx4HvIZIoP5UPEdDoraLd8CJl1mVPHcYeDLQisFXG4XPgwXySX
g+48OxkNuOsjiLLrYJB2Sdb+ttQ7wgROOWWwbMqk1eRwoFizCAUQLDc2qrML
8EeFG13C/EQ5OQXh/1wVEhJT/xyHvjkbuclXV/n6bJ9pxKSL09I35BXtlop+
eHxB1Ufi/Yu11F/Df4ynSCmgb8Jr+2MFHuBSEDSR6+D8a8yuo/TKie0Z+DE6
E2mifQwc8S8mdwKarJgD6xwPkKCy2ZQeD3W5OUhMnNndaVwj6IT5OadoTHJn
z4aKHch8qy2b/y71j3iGxdVKL3XQoPSfS9VdswQOqWLOO3ig4jCr7N+SPO4k
YguFePf87x3FN/lFnva3pFZg7LpoupWmIjuBRie2LvJbqHkqz32svFin1zKf
mVq+yChk2VBCFUyb9TtUDJkeaPTTRVGsAEIALpQTh1qDd+hLp4DvGNID7UKq
CZMKKh0JUoahxQX89SNRpwDWbodi9fQLzpxT0k7FZ4/m1qKj/CdXEc17Hil3
cMmKciVqPhCbbyoQuFB3q3pKHZXmtjq+b2vHWUqAFYeOows3cXHbEcQ3B3Gj
cd+tbf9OmOdgb8u6rPIJDXP1sFwOvYSPkt9Ri0dm6APDbUibBjHwCNRy7dbw
xO6ixMw7Gjxac28Q5OzV2FGfe0CB2kaZfedC0MlgLy2nYNf6ZgPG1leU6oo2
kBbBxr5h39K77ol7S3JjucfqQYOJiOt9dK4h1PK/4cnBZ7+52MYjTpasLC5p
dq/zHBvyVDWqj//EWw4BS6eE1gZ5zrS2LLUIg8LQu+K3AmJCwxjz93A19l1D
DGZk10hSoeGPNXKrnoi3hHFjfjd/qJIS/kKXHpYQ2PRbIFmqRPhzC7E0h/1w
gv02PXoP3PJ4zfpDtWLHA1cmM4AZbCIufeDlRrmFVFPGWjq/Y/a/lnLK9e00
BA50YSjWvI5+6hbP2aulCBlvxbwRNHYYw45M38/CzGOarsMXIoRu7gk7lzvw
Yg32qCJLTQjpxYDA2vQjM1jbX9GD3/2oLEYgn6geU7eO0NGnqmbFh+csSe07
sSSMgcs5rWiRr417vAetxcUG7ApNAJ6JB+poPpIFrgHI4c8FOxFlX34PJwy1
s4X0hReSyb1Evo6AE4H+2FEeZHZRFbr/YfrSv8U4Wmf4XZg3PRZu7xSnU/Ix
ZTZQU/QK8vgK6Mur75P5TM26oYvNvjJMd+gu33T/bwlB3JG6tlJQcijDHIWr
LuDuqRUEZuhWrjX8pPKakah/nhz9vZwbp8VRHhF+/e2DmFDt+pvg080R8Xld
IqD5LD655vB/vNQ8rcOsjrt1J9qb9DheeLEASSX7bSmvPPESKBpjrF3umLgs
uTZ8b2x4u8I224xxBfrWDQXXOwCdspL11Nvh7KsxtnsajkTjixmogbmbB9MB
QL8k9lIIkaCKc52PdOEOx990NWSlT6Lo4eJA70dmtF5LRzMFFJdphVkw0Jtr
DKaTsjgMeytcnZ95LSdnDtIfInVuEiqmOuxCU3vKeaIMdNZ0VDBOhLvS79h5
qFtJlCnbybxWTJckV1ZF4jcs0vVelDc3g/qaDiqDdZv045kGfkJ1YaALdHU1
bLs6vqA7NWUR4uGbnhgH/9oyeGv6pZPC3/oQuBp1Us2LgdZzI68vNuGErpK2
1tdVdFoROeAR1VYMb3sBFtVYS3h0QnrEAV9AqOzr3oRaS5fbeXeX1SbkDn0N
zYT93+yuVdacatfCEsNeKuWYBzBxAQhDwDD/xV2UgMqzkw3wq+KBEvwQzLUb
/0wO1oZMBbgYubGMdndphVGG4PAFJn6A8fZ+ucDq3lqmvB4vbXX5gDpyQ+Tb
HNe0TRT7jELO/a7gm8dyaOfdXSz0sVBaaSlA1IhV+7AxyGHtw7wjPJI4zT8B
VJRvmtffc+/o+Fy1P7amUO/GWJUTpiBKCIQLinZ2PYTSdWEANDX9dwJnQmXk
paQ6u4h5Uh+WQgUSxJF1av1Z6J+baBOBATotg5Ne6RYwmhMKq+0nyJM272XR
WprU+2z/jsRNfGtzU/jui38qZb4jCyqavnb/PyqCRdIJecCHu+Fx77CrfZBM
H5DkFBbCsZrV4NcqA/AN6sPIVvM9rBJIvPzNftcrhzkWsQib46MZZ1Pe6lEw
iCEt9TGEVoliQHpM/c/QElYdJP+goWNShgDYfWRdw6CKBu/c60nxpU/+lKuM
dLjcPTgDqSCZ46iPpoeEvju3BLyf9XZ7vOCsxl3xsyeBS8xPV+5Jw9MldNz+
yi4fC0q8njKdTaDo4N+COw9iAoza2qz4LRm5RS1CuH5GB2gf27GiBI6vjZrY
u7lw0jiJu28q3f92aJ3fX+K9bws9FIVg+o7Ob2Jh+sRRvfwaeDa6jA68KQiK
LLsjLvANIN3VazfGZWeuyEEgn7x2CaWFJr2y7UEuMwZFFW/Wk4pC+Vqcvu7K
P/Ekq8wByw6NrHfEE5XjrZL4o6q4iUCEabkGSr5BoZoUko743qFI0tQLjL8b
SQTCQmcRGvJokVKDkBDeb4/rVt0TrbFoIQNe5LXDoLnLWdgobe+Z5URMVAaU
K5TwrRa7YPv8LBi2U4EITGEtD9kuzpbwAmtPp02Tv/A9W81GCkf4HTM3Hj1G
G1ItdmqHWRyckWcSOitS0Kau3UfEr3BtO1Ll35NV4oJDQeJH4cuK3glO5W2J
nZ/Diyrf6u7v8KS7A2NHbHQePQxzrTRLDKdUojvUp+XOsxBrNgVv7+KNkOew
Ipzurf13231t/sZfK/6rtdkeUZqHW9NpDQFWg4ECzYUUaXaSjW3Pxhy8MavA
9by/ZZw1ycwnXAh9QeYFuC8CBvsp6yn45HISQgXuzyhPU2mQHhTIHUS3r/C3
akpj24kqVpRnUb0FRv4aXNmnxoxXy+CIk0o/PK+vIdqMTOjEVgmYa470gksy
K1+kNCKpL5U/Ie6dtfk+czGDxBj3+rikG1UpEJNxj0YNa4mmx+L33KSdW50Y
GlXjiqB+2fRGnAipExX92EDELdcTVA64b3x2tFL9WzIjw5AMO2yK7ngxnOiH
bH7mTDIv2Ywe23xDPy2lFVXq/NdD15EnCdzrjCi3UstVLqe+n+sUeCEDbVbQ
bucf40RgYIqy6TJISmFtoNJSddkp0CjGI+S7/bk/Jjh5qtjqlj7qZKM3CvaA
dRDATH3yMC4sOH9Et6C1O8hihBVkAOkwpGS5BYsMSycFod10EEM1DNy/2ZSV
0PwaRJ3N//kkteg3GtjTRl092i8rlRQy0WFOuGO7lcmabtqZMxgNMzUL/EHt
K7kag5Mn4M/kVD011zGVMDoMpLfa9K9CSQy/BKExqTvH58E3tOIoxSqhPzet
Mlq7KPzGGaKaDUB1J93oan7aW/sSodVB6HaAu9T5gA1wNz9aZYtk4KgCp0No
LSsjnEJ+gztSlNEWOiMV0UUvy5Q/5GG24tEw+ZYKRe3vPpoCtNvHSpgwsS2s
7rrBif1E7ip0tzOxxiupPX1JuwTEbxUhE5HzQtElnzMCCwNb150pRmkaozqp
xb0wizRDjU++keiVJI9u2o5J0ti0KdTutItlq6nY9+1dzQ68tJNvk3ImxprG
BF4zYRAUF162p2Y2KTdTsx2V6bFlCZEvn6BjBxYtQBzSvk6nAJcMb7YVViKn
RXgqZcIlBGCsBtqNFDu7Y3Xeu5LowZfXDediLuS2RcigkYxj9g3Lk5RinXdi
FIE+V6Db6fwtoafre/kuyDl2BaWxJbQVQCiS0Kh742NG4o5oafHXP6h57F3U
vuA76+ALICHJ/k8guZbuB6CTNJz+9SzXKIAHtm7mZT1DhpxMUSHzUHaar5e+
4a+edZlPZ/RRR/XPIKjv8Enn78se+qe4mbMf9+/biIvlgwL5QlPd9UCPMF+I
MPOhk6/azpKuSiSJGorFCNLsPq9h+8C/RqwN1aMY23ZkN2Cf+jBtp2HhGiHE
snx+KRchXvlZgrlTeIT90Q4AxYB6gpPJME0GJ12BAR42NPqauIBBVKBFotUH
bw9YjBIp/Yq1A/DMcUcXExayM0BnXocz/jBCi9CrCfPALpfBgaLu4dE2kIjp
tcyQJ0BFemlBTIRS/QJdMZ1mSUfMnN6auVpreOjMKo6v6ihUrIRFi9wD0G5x
Ud7Tr/R8h1efvUSrunkgPCvTg96hw2O25wB8DqCBa7XbPZrssmFQxgToLx8C
VlalyyjJv04Ik2/svHrDq5dSYthQr4C7ICAIOvLeExWnzMn91y1kMgqhHOJp
aQwyut9fCdT2DkEJEsqsDxgjaeMS/UzhCi+whaS+ffdw80XNiFjjPnTYGjBt
Cv7G4VQu9I5hy47H9E/RDRk5XR8dLVbZU/LWdH1Q5873WwLxcK0wVmxwf1iZ
P99l5JVvUzpbAcicPN0F/uwZKln8uFtF+1Mf84vl306FRvmewaoXMsB5bY90
sED9CKI7UPFj1cmzIckcsTrNGx6yL472dctgcpE5oAkap/1CWNq9cOG3C246
+TiuxlvI/QB/E6iWe2dO/rxnqYv8jZGsI/OA9oz4NCvIG4VMOLJ22aTz6DjQ
N+iW0m5HLu+kpn3XXlRJFwrJ5r/u/Q3POfeKWV5D+MgkOGduTsiiP2hr0st7
iMcMNcB5msh9+Y1EBV4mHmcpIZsXarpMsAqZTq12lfK8p+Ppi84//KLGfJhr
9YA6anCmcA3iv1Il1wGx0QFE9CvSle+FaMUevhXnz85GZuJikmxQEslb7tfZ
gv5qVkSDgs/guGYD0IhVoYO0hArHAXXqFGm4zjYUhztCVPMv4cQi1e1e/bPC
apqYZkJsMVAOl+RWRtSEo2Mc4nSTaxoyBJIFRZH0WEc58ytcwC8OVrYR7PqS
K4TnirvhZOI0FVYeUmhUEDrybmb1CImm1YhtZulT+bd+QHY+WD5gvbtO2+V7
Z8MwTLVE/WEEsRtHVMx9sz+oFr8/6tVAE6LBLZEBHC55xutum5QbqH+bVNyf
hoRJgCiZM+Cdr91uiy2qWdOrf3lUCyLqphs7Y5ojTWCvmrCYF5YkXW2gaY2E
lt3I8M+KcQPJ1/0a8pjNzxfTf5lCODJrZv6/dMbK0v0gStjiJDhrUbSGRO6f
IekANUHnSi68OMmtg39EhAOo96jtNSW2SG7i7Py/pJIqQkKQJfMur1WbFxVj
e1lKX3WXRX6cftE7soQ/+depApnLioIHIdn4tCLsZe5hGDqyi0N1Fp3Cikxq
EkMhKbz82en/207ALuU9KPYPqEq1PxhoU/JKMvrsTOlX+gkeoD3A1X+h7PjR
3+T4jSCMroD3zlG9fdK6kHnGfTgRBlmT+WLwL/ZZy3PTAdFy7jshOxI5eurb
nTRB+PKB0RWPC3f1sv2QY4nHfNNB2G00fuGI3gGINCI5xJQCPWtkd0zqO43C
aQKWuBLDAVlZj27i3nUXfUq2RRsqxwrHybEEVmdu1eR6ZAkkzKlycIhPvdS6
n6LpLlxSQuLnJjQfsv/pj2kzPxJpYOnWb7qropSJCo6Gp6TAUdAnQebfpQ3O
zJ/7NXY3Qe6JVFlKM7rCf2QQ6gZbxIyVam/9YiQPPKxYbveF4bZa60Zhv8Is
f97qbILPPpdUf7HoSZbrzDrgxZtusyQYGutm23Vwi5iN/YXpPxQjM1l/wFQ8
iEYuNrB5y6QAxlHJlflDwCaQ7x+5iH64MZCohGRpHj6AqKq+iHKZ5nt4prKK
EAHDYPWypz7TpNXS3yvq3TGMca50660nRU1/ia5Uq8SfxIqV8xSD5C53rqJu
zH2LW4oHdegTr8yFfA1P8rkblg1/e5tD5eoQx80nOdVvhDeS7o6/55alST7y
Yr+BZJrX9b2Po2hJvNAuTB6cRexJHtAWqE3ik5c5VIJWVkxlI+RAvv8oDVAy
s7BNZscQdpaUqjctjNRUstR+L3QCM2vGw1BVJCEc7M6ruXUvB1gB04XfxvKH
lQcxUXyEX46sQ4EiEyh/FpgfjsMEiPNgIFWI6HJZxGPMsMQjcI6N0cIszpbS
8bUnP5osnE4+6nJD5FDhYuJLbguVMCFvphnfM6RE1jLvDwFCsf/0jDunnMtO
AoAWoTsFv7Wal93Nl+q5Fxxlue88A22eS9RKiM39u1iKTPz4s1iEuYIyfrUS
jqUA4/sF5XgJS/x8ZoETDLF0Yk4RS564TOU1vBYxEh7SohDL/84PdnH7TRzj
JEZUbfwlkUNXYjsv4XNW/Q9jfyjd5VFflzUvaT6bKKj4WOBoU/mng1FYIMJF
SkjfStv/Scn3NdKdTpMUEmTr7mxmey1k8WdmtTpmPMmZ13Z5jLNPn2OJOV9m
287eJhBp9AVpCBViD81YjpeL2ZMnp5pL0uYwPawcSo1vWVHvinYxMARs4l9G
gHiNzYAAa3uNheRem2m7EwaWB4kbCjEd5+w8bgU6NacRFbGoZSEccxWCqG8B
erVST6Twr8t94cz+qSL2XiKIna6Gz9rkPJ5DBtlx8FrWmmoNXgC8qm/1uAoN
NwDRckviN7b6/UqbSUbYXYIrr9DUGW7+garJGfWVQovq19G+UpQJGEx/kUjl
0UZ/B9CvLbzX02cUrHZwZG8ML4CSG85JfsAL4HBKb7Sp+USpoRV0+Iv0/Zwe
yXA5I56WlKWtEGvBt0pWNRxOISRh3NtaaclZzctYKOvJee2dlTseYfnHEdPB
SKSZbUUkftOmKLw8pwJGbT27yrVJN8cWDYbVamqC+EfXb33D2t+x7g7Osda0
XbfDybAv2cceUbLLRIzy0ZCg3Mj7hxq2UMTSV9cuGw6pe2y26xITFQKAkU7+
if6NMq9ENt3MEdch2cIkbWFYPgwtJgJskVn4NlQlHxaGGLQjpDIIdERi3SXS
0GXtk8InV52Ei8jEN8FaCn5wl5WFJy0+wT0pvf164b9Hm5uSvtxeq2fybl2y
89oLdChbtXH3wx4wWHTiL/GDDOSOp5kKCK0Hk4gIcK/EgY/XOXnKW+Qg1hR3
/qhxVCGGZwORlvqkgtLTKZxkp44sIvBQ3gLv1arinNGkEQA+edmJOgJu09lo
SqkTqVeIVJdtVaCC83V/FzQqCjKtllFdSdkbYXSrRi5t4ikp2CdbQeOx/Omb
qMd5F8ra/DEwC+nN0r9sMkqseR1tQbSlmg/Wnssxv7FDS4XjSMVv4PHDVivC
VmbzFi8mVmwNye0ihuP419C/3tyv1huI7SuXVam4svHkvqIt8ArGHaid1ixL
guW/1shksVy/M2OaF4CagohBrPxTIuNqWg2hUc5swdv24teQ0qdTq72vdGPN
j6xOFE/uIEIoT+miN4AmCWjc6RpstsqEsOvcgQpGXLJ2+rAwiZmWUba+nJAQ
As8KUIbu83rxKrqGvy1lSWm8vaCNcMJQL0JcWSBL0FKEQijDbbxctL4F7KKd
ygJbw8e/KJFEPzXR0HcTM0a1y/phgmxVqxAhY7sdWwrFngUvgARhGNnxh06m
sgRq5BSfV9iNjuwc5SKcGs459v7CrJEqwOSMd6Ma83sN4MP2FVNyl66VpTvi
jhlNCrPvi5IFTHEBiFcTLOyXqKpFrDXC6FyQQfuOzsR/2JeCEKTipmZgvpyF
jdOv4bkqcODJTm9Wk6cpv46p1chJgEOBcUoYrKPT+4ezKjjy+0mU+AtG4LFH
wsxdkuE7DqAKj1qsxhRKy7c28orzLEF/64SRj+U/Ab9QAiXsSljfN5h6CUph
DQhzw2zvbXfy5UDXIyidId6wTkTOWxU5vJacQLysQYZGgtr50qCDjsFS7wRA
+qwt9sFMETTZEeUoBsm9DukC+NGvi1tp3Ikn6xLf+n/fje48aJt15+D4iJtE
a8rpwrBQWtiQ8yxghN1ZElgXSj+8L795BMWr6lFkOHnk0BeIWaFs484iGpYR
criJL0/IOulnbNSn/Lrn/BqjImD83tYRiDiv8vmt3f6hntfkan90RoHu8KF+
u8o6TAUDjkqZwlFlSH80z7FhEDR7MR5a5tG7R/tIVE707jBaqYCVY2Nj+BIl
Gywb+eczio0QdIH4rsUt3s63G0IlyeqLPLCDBivGbrcuShLBYixXcZMaLaJs
oIIhmZK8qkCGD+WiEfGhb7tXGMHaL8R+GpKLE4kfBr7B3B96BfWQBnUBL4rM
cZPtxE9X9NmMRbubLdki4NJZhTf4W02+R1BLLBgCzfxHJ+JlJ4K0cNELbiGu
+1WO757u3B0yW7aGeyeTWG4M4m8tfkv85KD8HQQkDFEPzbz9nQFfbb/J2PS3
dH9l3Em3p5rH7W0piuV67tDoCu9vd9cs9/Nl2CZZtmMwP12qqYFkBesRzuwg
gyLB/ViiwTMt+NrKtLGyBPWX2LbGe30OW5kvoEDYafdtydrAIifuUTgoQX5d
MEBffXdawO+eeSDKTblqbB/08ZXmjChxB54Ov+TQ2qLzA/sGkBdcXA+Sre0K
Tj1P5qK84RGarggC6XGGqcAmBOm6U/NqQo0Cbl/4i2pPJS3/iRVJiQsJ4fK1
RqwYhhem0e84bYVY/jSFcHuc5sMkfKUbtcO/HOXxOUTQ13b9Bvj8y8KYNJSO
fTbao+UHBhwqvMNYsV//1yFDLF/SBwlIUGTsJfMut9G5gNM4FZq/2xtvzJmY
ML06x5lBi0fVXdVFx4fRc2ruizLulgrpqKs/DQBooUJyRJaJP5wrrzjzB2gs
nWCvSKhj3PkEfSZo9XIKP88WFrGU5zTQTB465T4VDuBixYHGTgeGNSeaxnhJ
Wd/ne13Kk9euG+c14wNASP9Liw+X28/v3P/Hmueq/WKJCPJ3Mi5hr9lH8hj/
NmgcT+ASXLwknmA3yby2XVKx6vRT2y4NTtEsYqR2oW4ydmeQ3UEWXrCSycK2
5d3bz3vaFXmWlJieCHg0wpP+zNaaUfp9VSTQ+D6LbDQISi4IIKbqRlQSGk/7
Kf7tYRWKU/TTS2nPvKLrWBMrdy+GcYhaKthjqeFxQFlPsAfShvju/fiDjDpB
o08b4wYLCq783SQzeOGW/r85+3PbRmonX4fyyNfv5tziEzmXdtS4noMyUJi0
Mfoi6fXkaqdRu4jG57BFEXaexjhqOW4YSI+GpNHUJjqW+iEen3PAnauLQhVE
KtdES7fQsUQPf0/NjZseG2A29MavoNZcWlkwfg30l0aClZjkggHR1zSqokk+
5nzCofrclnBN22pCaQjxBhnm+2ohTVXLrp+rRpUAkxqAu6c3wN92vLTa+Gn7
Z4thc0yJISKpbqnNTV3IL+vbgjPzMf5BHH7pVQ+x4CsQDX/HQSww7pgdZ/Gq
pxBhnC0osp1Q0wBFMvkfPVEIgKtXWzbaNgheGwXftbQIYF9GlwddtejC2PRu
8g3eusQeZtn6m6Z+EHHDPALFZHsH0JpvjU1JnlKy2+GT6yboh2EfxQjgc3rG
OvsfzjAnHvvPV0n0rQw/oYlIOo88xHZ8Awuk/Y3ytZgJDrq5RXPniL/3gvyz
vzugAOmm6bRcl0XNR9kkR5S+sqBdUwbqQDrzEZFV0QnilTdAdjnb4dqOL+Pb
yxE8Jb1ds5Ru5IG+v04KSblfcnTJjRe7Cr0t0rwk0k7SooZjH/e0ULpLMNoZ
lsgZ5GRAlBbhRhcvNLXQe+ZnObkfDEjn7ATNotck0QgpYl5MY+RqlNLgDLsj
lH5cVc8CyZUekHCZLdnhTJAvetDzrvvusseG/WuE5nu5X2r/AWMFb4uJOp4o
f/Ihn71Jh/IofO70zyIBw51VkO2Bo52lxXKHcywKm4PuyXCKqVLt+nqpUemq
ilWJ9u+tLKNY6isr4FNGi8rJ5W2RTNbTL2DWpexR7Mby/23gEJcWRQc6gqhD
0EhazvUUfteTwf3YERzzkT02nptfl8S8+TnjsardcMjACBcO6mIPeYdvFSBh
AGpNXwdAorWdG3a+McY8O467auoVmQxC/Sc5qSS1G8mn3i8uCh1GhFFc7DNO
Pxz5a9bJVym2wsp8QCDIvmjdwWX/MhiVx8WoumyTcwgywopMjbcFAm4Em092
TaEqnvGFeSpUiOu8FLK+4nkjpYKyjFWXpppUCNEnjZOpukmnQdj7FNi4a5sv
GfyDMucWAYWDBy6SrexpCXEyA2J9rt5Y96iFyG2xmiOrBPrA13BkU20i1A2u
J7ZeTRFxgLvx88OZfB2drpyITgDOtdpognXPxXSobhxI2iV3cWDVQmapplgH
B1Dod4XsYXlkMA9wnfN/P1lmiFaa5cmlD+Gfy5+ZcTtOwkeFalXvlnPhHVgy
y3lIR5NaR9XCTlZDHB14xPCW0t3pJ9kwihfPcoXUu9C5COFAPLefjn/Eoza3
hOcL71MoM5/5VXJDEMrwfrzH61D37IHCgTVO7JiWsTpHKkA4Ku3D4dMRUKsd
rbUamMJ7erp5821YBR4TFLXCCz+8uHNpRIsQg8dVha1sl4k2aeVUYtcuYjRe
ZAAbm8+FmMEg2tBVZh9gDjkUaxrjEbQ+zsoBYYEJgnt5yAneyL0itLroCKRX
RnfR/pqn2FF9iHjEuccIgtb9sS5gFTApLovsNOudIV23V1pPvEf8SdsCucPK
G6tw877xks/SM8F3pmP3NeH2qeK63LR0ikydwi+FEmV1WjvnwX7RqCyrMZhK
9UnJ/1zIBeBks0Km5b44ZOAOOI7uYOkFuIzTd1MxeeTPGt0vTQHUYjYq12uE
ggoC0HpDy3Bw6QjKN5s12NqiES8gTu6dCgfO/mbY1eSy9kTymqFGJnvNbsbZ
L7aWSpuoFnyKgsNht7hAVltzojHfcSQ4iv6E5LEfbbiH6GaA0Uh+oXfVFRSw
yIj4RgHqNLvGa3cEEPpx4TkWRtzWSY0ObAtnDiKtS/8HMqbRrFJqGKhBcuxR
AnFMj1bx0PVosXMgNJ8YptmbpmuxQUQ69Eiet85qQL5100bIDYiH9ToLwZ6K
O9cobmZqY69SvUQTKSkkVTKlIy6uH4894cz9AA5uPkJoLeqSTF+WpdrXCfwm
WGuQCcfKztYB844I0INHQ7/Ec+3nId2Z2tgALEiy6KvAb01Ui6NeIz6aSzZV
hkwMX1KpEHYfEt3Mzht284zc63pnDq+b09G1iR9t0E7jn1SyrxlhxU06vgSc
8NjJvEETMuixAWy2OS6OFnTGO+X3RH3wnPbk1umLEtpkN0noz18QEFq8OwDA
iv06PAzqi+TCH/RpBGKHrcOvhwl8d7UkW/1AtNyYiXdLwI74ety9HkuQRW+7
fhPRea5HaO3Hqoi9H3E/Lh0DjKCcJq/FUgkhmFnx57DKkoFwKafxZMGX558r
gt5nxaEzqnSvetffXj+Gq4oypxA+cldvAJULUNDuLrlHAhWYV19XA/h8LFu7
I1d6dN4DlgR3OeKtSqRt5qd6O3ldkyDqdTAz80Nvm9r2Ne5f/s30Y+nh7olS
qBlAx4roh3gPsmSF5jS+KgpK0o5apuwV7ol1bMJf5jtms/O4bw/VrxSQP2kv
S4a6mkDndpx3dPgJGh8VWYM6KpkEuC1gFDxEHfjlnB+zSWLshfodoYK0BXKU
OQjAYDeUnZ1U6iuUbYcTsRYOTzZN9z5SC2GTQYjQAodg6QAx0ZdHqwRp1gRI
wVR+qVUrSUoEYZ8ynqyOFY3V7r/fYuzjS4u0JhWluqwYR9RV9sRrhh71pM8c
ZnclVmYK/ZbZeNWLQXTZXnUTy8mE8P0WWd/tbi18xyymdHL2mkXHH/HXyi8v
xe9FxIF0R3spxphaTJm7QMRI/tF4kX0rS2QeRLkYC7ZZexq430MUfZKYInFc
MU2TuL7+zc15MclugmWmojkIgFN2MmGCY/QsVCobG8wdmgyHkGwcrkDy/bTc
0+mLSh1y/bFRSKoS0O3cQuBhKpXegu7O05he8nVe3NeoZ9sWATbbUzp5BAaT
IJYqpazbah1ZywnZa7XXPd/GolpAT81KZ6CIT85+4mksiZnCPLASidD2f00G
TVEoc5o+wX4s8X9p383B0FozBy81Fb5fnjK/caePUzdmnca+IRR0bAPknM1B
FIqWhrfBasRo/dbGsxsvue5e+UGu05HnBbUxV0riWMUb9fxn3Bhrt3TTv3FW
S8Qv86Mi+kMaEX+cP1nN9Pju2WKSk7nYkdqtV/SF+wxCn64k31JkxdMyZEox
BTcUHpwoii6sT0DYmumwUkGKHHJtipO39RB2xXy2lMldUcd2GBzIdfozW+qH
aJbepJYDrXOpuzSSMQtrB7tGjIdzIVQG8ZBVAUaK+apbB0jFRfyzVC0bZdL8
KH3gW1LolYMeZ2Q26rvUWtRKrvml2MmHm4ZwCEgM5BdCzUXLK1HQtKYpr9LP
b+7f5arY2//+4/ZbeVZyJ0rg5KeWWAwms8ruLtF9F0VhOhJLOGO7IXfpl4Q8
n7Pl7d+Ay5GJ+LGUDAzAoosab77El9J+3w2Z6fs3hyoI/gjf6kvo/TJ5Q57f
07VU+GGzVK/XFnBLPUNDHPdmGWFsHdAuj4NgYQ5K03WH33q/pwX9KLJ02ve3
Efg46Fn1cyzF865TaSKF4yzkLNw7UEO+d50l71YZYmmN5phaFSArMaJRCoLD
jepKbcJ3LPgszwSjbw0f1mtdIFLkGLdiTn2Espu1c2kLc1rHRh3O007H6HZt
cic5xzgjHLtriJmfNyn5AG7eBYhlVdfJAY+BU6C5nWshQMtL11Ltzy3HSFH7
Y9zylunIG8aeCyM9Ef0ttnDDe5uC7VwHLIZCqpPAvzovxaVqAtIQ4kcM3rsA
EthvMAn3b5MW+NVMMxK4N/9h57/gqXdhKTKQ5ii4BYiCOisN3Ue/ORUNrNoo
xSC5IBz0cr8sCSQzA9KNGd0LDrF72me1BCtlCV+a56kG3VWesl24AAMVN1NT
R2fiATbzmfT8E+c9tstvqFX7d0Rz7VSWMKpkhPv+VqDDqk79GrrDNsfBby1G
hU9ErvdFVagpqzCEb+RD+CdKsOL7/Yr6dGB7LF2Rokpo5hzvgOaRH20YXLwV
M0r1+qLtokd5LVyfhQCeHYSuydiLRbbx9pitwQU2Ifo6VA2qtJROPGY4WYXL
vHU/1SZtkgeCUTNI0b4Iv0eRcIoQrYIv9UIdX2VIb6eJL99lEDConbTXtVDF
auxawY4XkFzlkkP6hMPy8sphqYbpyABHXXy2Yk6XGIXPhGSRRrjGxMIjuZxz
l2LEuS7t3X52F995+GUAFId0zbY2SgWCC8PM0OJVQsuUO8TXuYP/bHmXwpe4
uxadOFcell3b6TDsAPVwrmSFDcXjRdPd8eHG3BaCTVIX/T9s0yw1bZy8OzOS
49f3TvFCXY8GKrlka2BfJGkGnNYYzrxFVZGYcC+nNwY8QOLBXgJfDoOeYYzc
Bd3N5bMR83yb3BucqX52Sf9p4mLhVUlFkMgYDzAdXKiKLJOBO0g5gKIweC5g
nl5V3BQ08A6r09gS81P4t5XpLkcpi3/rxVx1slcVTFtzOVXqbvL0TvdhZzem
MZEVXslM/Dpwu31zoweCO/N+JsOibKhI/BIxDDSXjMXAEDJ01auyivF4KHQU
BQL7usfEbmjj7o2IF1taB6XuK4ZuB9baaA37GhqGVJop4HhQMMWw4UCMVXql
C0Ulzwbi9IsBiH1e2SHvAe6oBhTC0bZLBuR+PrQJ3LNgLU8r+acQCgSRQ3Kq
LRp7Fg+UUNSXZHN9GDrhufOZIh9Wp/xeXrpc68TrvGN2zbYAa5oFHG7F9/Xf
tlacNN7pmx3XGfBXQZESTMROaA0ETEwqifwJVnr9XYB3LYQTKZtizX2k8ZHV
NUhxCbs1Vd1QEw6Rb6V7VywGVDj6+8dKeBImRQ+TvW21oXtn26oLiEt3vGYj
aRqJzHCZbNft3f/woPHJG+t9cWUtUOFNLpH5m6nl/4O+fRr4+locNIeXAujQ
yPH2IUHTqQJ2OudvizVmRZz4Al4StwzehgnrKc8yna74N/au8XLGXcR1J+15
BIJx8pE79pobUMqPTdABjthWBJWrgCzcSGNYeTLjxfdBXpHLuDBEbMc3CmTj
AkG1iqVFeEQZECrA4ADwgfA07aW5SaH8o1zZu74/p9Opi5Eva5TRtIr+117Q
3yTbuAKgyK0oodqsl/1aB2yzmdc1pHLU/7AmvDkpRi9l2L3d5cKR8thb9nPY
gXCNKrXzJYR9VMY9Vja7JgwMPfYZNi1xt8N1BdtPRsir6Z0ha7es2E0+/bdt
B5DDeADKFZxvZxE8cl90nazr9CwJIyPsuYZuavQTCM809OLN42kREWVJQyBb
ZKbbMjlhbfXRdRMnoyGTbXLOQpaK+0Q6F/5+PlD7dMTV3fEY/3xQK//LeGxy
65ok/plaXpUEaEWY/8lKfoRIuhFv9eMAycfO5v1IdR3jPWS/JJfAqI1vCR89
eKosem5bhKfQjIwIp8qbHU685H5wGXDGzniA7PYdynLo29S3EKaHCINJCfrO
KYTP3A5/2dVWk0hR68GNWJw+Ss1FJumQMQazRh0QrTgv9b4CP2cEjtUiKEs4
e6Ff8SDF5T1KNha+EmcRlFiIDsKLbzZtBvw6r3ukMAhBOgbPlEC0VwQ/8KUG
EeIznh67+U5XykILpCX112HYGT3u8NVS24pg7Ga1bHnqeWn7QixNoHNTc4ha
J78QlDAzWU4N9VvpeGHnP705+qsNFnnM60TjYbka8qAiZW/rC4jZFBb5xAhe
4VUfpvTP2bxhYgiQi5Qy2bRrBY4ZLcbF2cF3wwEJtwkAQTiQZf8miOY6OL9u
YTAAac7o63YXK2BnVNB5EN8qxZi5zv/fvgWwWV4giGf/90qUwlKHQnovpvn0
FCtyq6w+Yluj4gEMzJ4modO5iNP/XW6zYSxPpZ5TzADomykFzYbDk8DLisKZ
QxdhPQWWMVcg+8acdXtPa4DNPJZpF/nxlBTTe4CtPR9gutnVqwFShZIxifV3
fomxZFFef7WJr4/6V9T3m7o/39IpsyOT/MoxqUUbzz9d09TbRc7Bdhz9NqxB
BG0JPqOhvSzilE8Iqp2GCmzXJNPTy9ouvl+P8XHHSriUYIB6LhklyV0ja8cH
qPR5ibl/f3ttN+jjsNmxZ+cWAJ5DBovAoIRN96a84WG4Wmxi6iYNM5+U7r8p
IhNWNO1mVC6VCWM391fMDJzU7o23iXSsMh0MrpQI7MjGhRx84vXlCYu9s5Rp
KpFK+ZMASgYzwOpHtUKpexsaQrAoOuVcfqz7bTAi75B5niRK6cWvXtp4uR67
7j2Z6sGvAZMOTxwytSR019qXteu84VUn+C2XNOGqV8k9n7hkMCBC62PCczEL
I24SFu7v1akfkblxKLezCQ6JxhIrMgKWMTZyrV0hAZQlcTf4pTdQBkAk6o4N
7ldo3eS/ntBPYB4QMSAsWTF3LXQSGlJSgIc8ws3ADmLPG6yXHrTyk1UmB63u
R57N2HxLGcBBP9FgQxQ5o9HRwkWLg2R27b/3c5hag0r1+eD2O+tV4+3JwckT
v/Hom5C5gEz65r+rnuHJXQOZypov1byb2lYnvrHXQPTR7zvDVBh6pSh8jW8F
nG5cEnf3miyG42Ewbr58JuCKrfAFspT4JR/xtq9Nc4y+QKWqYpQOoenS+49l
EX82YuZMvUFYQd08pKOsKY/GjXhueSQklRdK2nB12QdFf3dYIRVmHWffmTu2
r9YXCHJwqrlW4LQ2oNHis3ZINiya+h5azGBnYSmgbcbk/LZK02L6X5jsYFhH
I08JYi78fUGGCV/mow+TFOR5s7lZeT6VwZ4t7tiOjjQCtHv9yHNCF4QzeURj
qqWGlsOhJDKkr/A/GqCftdK9JndeHL8SoX7MeI8A9lgAu32kdpGM5gnWNMBz
X/MmL8Xu+4Gobm3NZFgmeroAQsMM3KY6t4O+j6fGMOLg9xRCxFtqr4iHDoZO
2Ixz03I8hE0FWDTVPZMvO6zZbRuMWiwmFurZBLZZq3XEOblH6uEj80N3KLQJ
mwroBjhMgeiKPF3yowTsnXz7ccunibyTa/jfCwtAIASWmT9dWeriSdoMSaDH
ij9WEL6a23OjOG2nxPiKkKZU4e+TiNEyuS9OYeHLX+9Wmxg1Wk2BPMlJws6c
iKC0cK8c+ix0/la3iOwmWwtakmhc7fFspB9HieXob7kXy19kMYWDr5lS2TXX
XU4XhSQZm5okaFVayJ/gBIgRt1WfqxZAVusneL9PHrPlIFrfus7JDsVGHHmH
wBHwJat6tLAuLbkT4ZsosiuGIxWz4Z528RIun9xtCnZ4Q4DWQ20lJzvhxwhF
aoXc6tvxIf5+aoF+H7TYzTJSM/WiZJ0Eo8qtug+Rn/7FV1wD6/Q45i38zwAY
TKkvt0pSl9pg1+JlHwaLqj97Ain1ybnkRpbHO35uNQma+x/Jh1lLVXZ0PvRw
7cz8VAciR1kzuuBQxmz83vuC9VLSMC7Ha90hXekKOnUsGbqjemu89WQ1aXR/
O0yY9gaiszDm23scvP2CZSDl9O2ZtXoUbbY+CW+1NkXMQk4UmJCG0wKJ5sJU
O5TkMlIbiJIOBetbJICxaZkYD0a0Hd/UiWuPWGpjjUJmPB/mLAm2A5H9cHwA
XcelLv02LMogzeozFNwtPSZj1Rnus03iK86ss8vk7cVd04QGAq+PvpfxX/nO
+zuE1wvRdwME/br23dAh7m7Vu9dQO4f0WZPoFVT8yncozZFOx6CecElufrBe
JV/SrO7UKqr1nlSX2dcH7YZEIqXcw+eQMcutTx5uOura+e/r553+gM21CIO3
DFpX1pg/yOAkMuDFmv2eL5bpmFcapX0hFYxd9KAn+eE3T+8RKR9pdxjOlN9R
507eZcAY5ASOQ2X8gFT4HqApj98jGssue7p6ejlBY0IlQbRjBK5dkrMxoh1T
pWCEdL5fO2FMR9HduSvS56I1DVcg38S3wBRDW8xhD0hL6zCRINyGbkNL1ksj
OQ5hgNjSOtkoD00vBBaizkuV3c+c0WIrYf6YRL6XPd+8QOy6qPWpC+N4WL7j
EJmHmt9N2IYZPx9XB8INQDqYCccUg6S2ZJJb1fPtc0H04PwTPLSFbTWEDkLe
U6GW8NHeruJVP71KG7dg5Qd5y/bqx8WybHvY4Vh82CFcHNZDN9bMMaOVvYIU
dpPpztCkkWIYjfYiFOtf06WY+kLz5AOSdPJ6LvsotfFljwlAxRFoh6S4DyOs
zTn1gu9+Fo6KqMfBphl0JU6W/ZQita77YC/EKwjYN5Rx5eUgEfVlePk/Efl+
nJKV+YqTcZhckG5IzAZYItFmMYc+FXFBJwQqblp96nmwTHOhCcIPiUKnNzLy
5YIdPdjhAGq+VFmi1JCKwO5hHYhaB9zK01t4ugI+wHc4a1NE6vLYGrVqGKo5
S1fQgHi9IRsI4f2j4DIUmwrykOmnJBXlwRdDkzo7mgq6BlL9+gNrByGsqUqq
7zCgU6Vy2CWeTiQmzvpK/rBmqXmYWV2evDO+xCN764nnyhyNkyhD/N/QWPq/
IVufOsXoqdU9D6XkvfWfsjefkfmRPeYNvUjKdOOGCtNWcgnpOdoCuxMwLWxH
GMk464X9wOBSlj/xjcQ+NSpQ5e2hSyNhrRW/GSa75FS0a9+3+Qsate/9/QdA
TlHOP32tP48uhTewgyLn0D4llYxgLJLcYm67ZLZZCT85D0bpGqhiGgNRrO3M
FfSVmebwf0mP7NfG0jRaXz/W7oQuDAeRM+O5lc79PHQ7f/8aVHlRXZxebrus
lXXRs/9ebsoZsqwCHlYHQEtJVxojAx31rWHlIB+jGIFlZOBx+aL/AZWmuMvu
5W7Ar2jK8r2+fyiekD6wLCeGuL3e/mSn5xGB7ldq/EyHfSB/MKR0DvGg5lvK
xlRsSXLbT4CYUWWZApv4DQa+5xRWKt6lrImJBS//QeT5cNVP99Y+DYuSzvWB
Q4nXWoLfR2opT5W4C+7ofoWOIEkHJKBEAlOoho6DRO2WH7GarnN8YAhLka1H
8Sxj2H0CQAwoADbCvtNcl7Hc1peeL1f52LyzlROGmkSmWsydy+GFNKmedwfn
oh8jVd0HHAA0dQ78ek/L7CxdEVcrM8V88gggom4iA3CiXWl5fUZP/kHm1GMc
/oDxyg/fql4ECkvN7HKECARoqvOUcq1BZefaby8SZLQ7JuWm1oGvGAyFE4XI
X9QeTu9tfFfgH9cu2tOjL0OxPS++2VmMmcmit5ayRfXcNhP1uRM+ENnpRoVn
iBSMpDnUanPyNSU38UT4bC29IBAZr8zkSBJbFULhP70Xam+BjxabTgE+jJP7
WD73ECvvFzRTNHaE/ONHmkaX5vrM2Ic5LPnLYB7O9eiRrDYVKFTklPkY8vox
X0MbGkUhkhKuhL8K7oMATwvPGGgYCq9oS1CKsBMEswHFbU+sxUwQ3XVEmGFg
wGeMZhCy2kqHXuRn5ShR4BadmozKP/TsPFfl9Xtxxa5CQ6oakEXJAAcZ9ceh
C3QKIPA6FMMZ5zancXMh4OXPshdrQvtmk7Qm3Db/1Htj35FUR48hoMB2Cp3w
OBDh4O9RFqOMENTdpF23PjO23E9fMRlHtYa7rEMPc9TAW63rea+BhcPV8YZW
+F09N0ccRC0BvcRxmtcE1sjWBbwKCjSUgHAY/SVbsXGDrYY1E1mT1mYVBxJY
ChvXT6Rr6LMadonzKwd5gsiRNQDUQzM2wu9QC232j+uyh6/FPaySlkcr8088
gIvmjPx39ptyZqCt24ohuXKwtMxqDibvzbw40z03kq5KzFvK/gTk0U8D6yRi
4oquSA+EekrzlkEAo/zhRm5fhLZh0cGcKxctDx7AFNlrV1kr8FJcBYXoftTY
OjvH9AtFMZpmPeLAMIZ99qFaTAjFai+ofyA29MjRpyc8QIag1K+97yE3ziDU
LLQaaEHfk9hUifH2Y4o0BHqEjM/3OJvDtRhRUOO6+8SqD8/qxrx4flcDLzu1
kA2P4RHhWtKqgNKlydYf5p/Cppzc6T4qz2K1TvLVOIfXjv+wX9sgkaL35hmA
bijNujClpbr3zYuDel3a/3eRgm3A9tEYko7pZ9PaPMhXTy0zu+ylteW3zGsr
tpg/WriJDvS+WE7Vb+2h8PStN+nEwByZFwoqi/tIDCk8mOarGYQo1F7WYiKA
QgOEQ3uah6dmoiKVSvJgVPf4e+5YWybTRSHfwUzbcUiLobLzGZavlUNI55FT
tQiwzheQ8byVq/FDBqq7dRTP/yu+SF/Cm5qvbucpT1ft0bblYvk7fbYCrpET
1dT1fOcfWHAUi58cgSZsP7/A5JJm4aAT/bhJRNENwloaN9o24Ha5tOJN2pug
Y8yoyt0YBwspshAuF1NtmRXFQCF8gDHMOXVaEwzT5wVNbjTbU7Dp1Z4fWNKR
V9glEwlvtvJaPgOh875xe4swIsEJlzSNOsHKRTaXt1QxKTX63gjBzBItj04N
AiR5W0GaXlwjKlW1fzPQq2BnaCYtNf0dSjHdF+ipStEBDFuItVvqaJGSI/R1
1N3Y2A6c6Agc7HxGhxw9Z9VHUO/iRyO8igfFM3ijHMBvHttkR1UO5O9tou9x
ZqAVowcq8VRvx04Tj/Tefpb6edDs23xP1kaQLalnsmC161RsF+8vThfVtLdC
cXU4iZ7dfd7TNut4+xS6GwuTAFLwwXSnf9RZzZyCVJLC6uJ6WGSIU4QA2XjE
pZjKNGpr6EHGbIJK9lpVQcDmBjyVpvUXDrebzRw6aeMctaR179MKTpZRJpTw
JcL5Q0WbD5/BQNo4z/GafbazSCO7wnZHAU2J87ZcowhbGjIlXEeY6US3lrGT
G7MtmDEex62c256QPic8FKU0mcLCtbpOMIG1ies0LJYZ7oofCBmswfF6zFII
UFC5nVfZa6mj/e/NKuOeRrAhmTix0KMbYbXSLQNFgk8BsAN1fodzIuNGD1+N
atQjVh8HrMGvcEcsM840ps6I9Kmjtfd06T06RS4/afYRXTafQlruJfSXT4rq
vB/FZ+SGQZH3LjXELbJKIVhc3IJmn5Ja/1FGBMUw0mPRAVYqWJ9MiykAB1by
HziumXFW8P9/PGNGd2PHs9n86+qmNSm3vGJJGNLsUc1655lwT/LoRhADPCcL
+fZMm1A+6yS0M+qEjBkvLDsmZWXk4YK1MiVPvB5MKH9zqFiMGx7BROcpfEXu
lUsfdW93gcRTItkTYjFshJTDKONpOwZHFuLILtmePjdJDniBoq0Z9N3fTFaZ
QkujbYtfHM78N9CChki8ZnFLWZdl6eFe5d6ZUfPpdVYcg5LhjdbY+NhRiAJM
BnOeWDx+i2F+JYaajBSRxtJppOlhCBwCS4BLbOtTisjEU8ZV/he69P1x8q9Q
hwF/N2h1y4gWqiueYNkNDbSp4NwWC/ymuqkFOQ1yAmkX/fEYpaYZTWvV6EMW
A/nyw35aVAqDuK0t56VJWNLuq0f99eA3S706JjmfTC+/Q9EhTr+F8re/L4c5
wMTICcq1V+JkO2SDFCTSmy1HUZeGqXHchqLKejWnLxNWvvh+egwfrtC5R214
oj/UEghvauxwxmC4/1RuYovC+NZ39grWilJghYwbqxeJcvEuZflCVCmC04cU
IheH3TqCaoV/8rByWvKbZtOAZ1KMvdezFLeljkFBw6N8ZLI4dFxOE5R0FznC
1lNQ6PYL5wdek7vv18QaIs86wAxWADQBtgmJoAORqCc5wIT7phBDosFR7oix
tDdyqf1kbWtCdQfmqgSKsDHTgWv2y/hEMbOiAwMwNCopZzm6B6ja1lnncqDY
n0HtLP1TCfwAhuLLVS8c5EVsbkQYOPlsagjgFSLZeskKXRdxj1Uy9U2ZgS+j
V4yuMEZb92v5hZ1Lti2fPhmkAQHJz7Q0/I+7choWsAPy7wq8/jzSCH6qFB4V
83Cn0yexSbEGDBWc/jb1dZbMYi9dZMZdHTgok7uRfVD6czFBB1qsAwPoebax
p5Cu+OvlSF5Fy0v3XmItCICZHi2WLb/6qhob9yaPJOmhvnZGtNd6pQXwwWNV
vZIgjCHjMsuVwagCU5mfvj/9LFKROgusRe+NnkMQpF14F27U5d53NrcrY97S
h0pgCo8IcrIZ0tYoyEVUvWWoOeAcsTVuu3q6m9yaRtO9R+9qPtsPynv6V/IY
DxY3QBem7MBHGjQenH5le6W5FxMP15BefeseuzvENGdOn5S/OVD820pcgBlS
gZidbZ0QJDFFVp9vPpcYmfoksOp2FWbC1n9JKmg1zNxG/+yDx5XpwhCfMcFF
yUaroIER29BsnYMfTDxQx2NpgZ7J7NSOaUS04gw5AXjZX83ko7PjWbXDbu4s
bth4AxIIt/v7lEWxjTbCRxzAhGp8y/zCcl3q1hMuD2rbWKFOIw1Jh0XHbE8H
MCbko+V3c2hOrRqjIJQZ6Uf/QnGsqxsVk3yDeHitfxw++b5GEGVjdB8h7KPr
7hv77eAmF4raX8+e8N4y/VEPHKy3U0/+JS4gJg1WPbjTlpyprFZg8iOpvZgF
gSJKmvyFwSrwEn199O3KrHmz9IgmeA/LwEmvoniVYvTgGRtMTHsX96J5tgr2
boB+isfw5Xp9/EDqd4Va/HEc+bCigD5BklLJQRQjjV0R3Ai/dGPKrsFVRojY
kANduQHvfmu+7I/cneOS8oH4JibvCgnBDmd2rM7dy3cYZ5k6z/eoM+9vBEuB
tfYlp50fpjIfubKsB+ZI7+RjIj3P7xZbjyaF1JwWw71nl8VlVtWJPv8lPO+a
XgL1tMpYU55BLsD8AZR/2QvzkFmM26yj9VpgimrTeMf3Rhgy5nZg7DwAReqX
j2xkvpebt/Ey7cra5XSWwLw/4X5P/Rm4HUmVF6kwAtf/3r9ng4K+x+ZkIfAe
6zbrV81PwZYgyke4kff9zkdiw1Li5fYRpDYighsFri793vPpPZzzxoFIS2OB
ngzPkD5jU8MDnfbksqVESO3I+ohdnUIiAAlJB0dM1Z+mlDjw8+sTdEqL4nEW
R50ZY2VzWrKPyign5lke+3iC6QergQCwWUUSo6BG+BrgTrm1BtZHE5om7sVW
7fXnEYxZ0lx7FCF2GxdrQ9jnD5/KZqLODQ0U5fpgTDIQH7htX0xj5H65w4KI
Iniws43G2Ogb5PZfh9oUAjVkqA4xrWaw7YbFlyJmI8DMZguKW07Tp2PNeqoc
f+Syiut3GSH0/NEHNj7iiLWaUAWgd9b41apKljz8Ojki7oEPhYLcudDN5ib3
7BROu1WY38BZQth2pDKkMTu6oZtk1V4VrvRze+5KdMDwQKhcmKi4BH+KEwLr
zNIqGbK55WRDsVOzP1k1inYcbCFbvlWfpXmR9cqCJHTfb0cVLe9+qZ1j4ezc
p856zQBa64rHZ67ivc3bVhdRs00js/wbhY+8iuMUCSf8eA/UxfH+MQYWAX5i
P+xdpLSPYyEgZxf+fO7XDkAnWFApGOBVv//6KxiOK4Ru7HzaILzPNH63CJf5
90LGcoKgIG3nIl0kQjldYeCDAkXcoSe8CbTCb+BQ5N/TPx2PMwtvWEYxTMhN
ua1w34lSJnafryO+6jVqJ5ifU4zARDhVW9MjnCyJxBEqCRe04CC2wUWz21V6
/nukQOOW8r4PfRGdqxP1I1KT3W4oXkJg60XfM0Qc18IJxbOHbIuXOUenxxXN
/oKe23Yy9xbFzhzYAejqNBy/7MuNMfwGpWtJhWL7+QFQHSPdW1B593TL93kr
vHPNgC6HgPGQoXyenbj42vljkTFkFyBtb0Sc/cMraOpHwv4Sei8uruhEgM4X
PUQXnHsi926XvlbBgPGDq33pYD7tnHMXSCi//5JzqgLc0wD/1pIDk/JS0c9E
f46SSLM5D4RKFNPB0gYk7O62NoCopkXwfq8zuFrbg4vzrnpmvss5RmZu65P+
CMWv/f3+nRj73iQ+eza5/9W0mX0X2GCM5vd14hzZOVqlVYTNjWjiOm5GI4yB
Ro1utkidWhGCiVKn3GEV+6O5SRV7CRqxNCfcXb3brWy7zgAxWmp0Z9fPio7n
NXSUfGWiVHYHbDYrbjN9FQV1RLa86rbSio8Fyv0A2/CD6tmzJ+4AmmRpPv6Y
uTBBQHL+ng83ea+vUMtJwHrbA1eaJTGx0Bq31TH40xT9tJmE7DHlQqrsUmnE
1UQsjGC2Ac3CycSLfqlbGHG9BajZuYgBER7kGAkmLWG9gfWBs6Kg3sPHJU40
BY8YUho70XvtEZB0INE/g5cUBvSaUbTRbKA9CsM0E3ayinGo5kTSJhQ6utIb
cf4aG6R6hWTmXCzN7UOG8fzsxYAggHb7GS+NddrrXlP/Dr1B/hDH2dObMaMJ
0Ip4bowXC5SYfSh+sXz+XrkygnWyzURxvWM75DMJiGzbOU09WnbiLXrU76kj
9vflqjnCHTWJjAhgjMvvKKFPvZGWhuagD9vOFfIi9hOrePzMYTLOkvhedZ/W
B4gZWqUb1bTOkZTe7G2a0Z7E9gIpQDMg0W1zLAL49KDXAqFjEyX2JDe5ZYq4
DxYTP0Ic8YVem7bXZkwk8VKHDSM/NaT2vuJ9XdiR2CKuKBeTMudyEaIYsH1l
fLHNPbjhYm+zsKAGhcewhfzrSCnZIuPL+xGJ/+e98X22wnTI6lBdrsNnSje9
rmmD9D//JeyEfnCY8begTuO/KMUYtbYDUhwnVoSiN4V3QQRzUMiKgj2P2IVd
VwiPHJ7T2jVPB9B7/ndiEgQwfkC4Nc7JkzouBpyh1tv4sTxErkLd+CgLABZ0
Z97KkQuN3XR+YbQ9DlEaeVokt6mpp0AL5Gs23cQTLUlHjsYNEZToScvEWYaJ
EBTYMy/9qfE+/kMl7KObTx/oIyXJsKiaOMjGIK26VFqnqEAoVYP90sV3mpo2
CcybQne6LEpbS9QqEw7Y5dTfNmDIAApGEolr557bGXOW7ixdtOFWEO5RyVYj
4Qt5TZy2ZtyzUl+nh9h0T0kGbEcvsRUeSX6UwMq3HwkoqPwHlCVINyMEwUTB
UiaemqTZ/Mq038uaNgPt1FHpnBQJMfILVx6otQqG66OIn/zuu+bLjx1NmhTW
h7VaaE7qyh9SFj6qsv5vo4LVdEMGhtRth9AXQTroGw7xSW9EU2ivtsPRrl89
QS71VRWxjyE7D3K+FW7HD3tVJbijTJ/WJhF0LR2cxOEDe1K2wxwKP7Uo1BZa
Zr0Xti4LbEFl7JYeMBT+SDUMgNusjUfHku/v+BW++d/CY0bQ1DdktB/QTmZq
wAVJtLwrcd/KzykmsYCwIY2cH6DgHE593O3fdEjQOgHSutJnmCLRg18E6qjJ
p9vRtfuPAnE1TDuPmwNAYTUTZiqPegrFrNufUUVzNfWNCULhu8dl6p+sL/jH
2ufkCr71nDgcm2OHFmKv5VOpxmCuf5KC7Wrnpl4hwmdC5YA4Bn3DPw9HO2tx
HoSe+75HD5hm1c35A6NNPbuisv/R//bL4gxmz0x0795z9bbIYRr11dkwbsXx
ssQTVnJujNs3FupIQ44V4EQg2iehCOEw1LLZUpIY5s2NTx0MA28/RXroXXYX
4WQ3ji12+oq8Vkun79mKGNDCbYSY6ugiqsQ3bkHW/g85G3FqxIFLXBPALzfv
DZOdu8ccieewEWrHW7LzXHmFe1Vr3qcfIibVpgN3OncqMJF13Z4yjyclnH3M
NJBPSs5vOY4uoDnT3Qz50QHfqala1T3cZzj8umY5x2UE9cFHBQQGLpgKdL3Y
Dh5O3bkgYXC2LiNATV2TMvmo4dH3bkVmIqz4FHUJGb0bM8afSYnLq/gtpke6
2xSnoIDiAu4B8GAST3qTp57hzyZcnfaFmOTERsO7STLXRHnSoFEzyKAztsU2
33wglO54zL5/YPkIBjNPmLaT3+aZpT7krpWX0TQJ4IfYBAo1tajfv/VaZDWu
QKE8A6FfKXdx1+//MagKIxyLa5Oe+srD4IVIcY4lP2AVMkksY6sJjyF4R0wP
k0fhbF2kFx3sK+ocnRbRL5uxs3xKvWwZJjQi3xiD/71SkdeZJVt8ffZYi+o2
LgegvLxrgB4nruNsTiGwYfmI6XKCVQNiaXc3JWhUm9exPjEabFeuqVBrxALQ
+tLSpH3duse/WCq3QHNNkOyqeT498FA2TaIpAWInaQWcnvsDgEy5HqNfHvhf
0e2u3JN1wMYGIkht44rFZ+J8WtRVx08xodx0lw14KVFYg1C37DrHR63czzfe
e0plgtOdxwOEGFE3o+PY7RkAP5oDUFqtPZIotnBSBc1uU6cHt9WukflReShv
xCXlNMPQieEYZWCJbHvyhyyD+qVfPcnjb0WtLFxyA4tg1/INYE++JGlCzCDd
Or2PKGeUKdcMBqmMRTIuNFlQ7K1zo175MQz6XE0guBhqvG7AVEuMYfkHATgP
0y7F79NboM3x+nxF9hhsN0pJXieK/YkpCgnoXwsIxhACmIbKdfAYb/bQUVJF
SoL0ChOw3OldDH/TJX9IpVAhHhYqya3ydJTdNH9yAytmj1WOAsXlqt820kFK
W+UZcVNcBm4XSfOZabxoglYqoAplRPW7wxEK8BdVnfu81gXJTVUjA0y5L3xy
v86o0tVi+u7/B08vxWJpPlxvZCXMCbxxWofh5xV3lsPIG0bEkARk6IEQw67J
5yokQykvRwfvOK2sATQZQtBRu7JTP+2U/k03bd/vQ4Qf1E5P7NUpkvglU64f
14ckhzaN2Y5y4o0tTCxBzX9Z8UqgLM9j1us36wifxccANKpC9G3nOCj+v0fB
ur2DeJgkxrK98k0T2tEuXgDVCKQygb7qiEADSg8YSkLDotUUB1ONPJ5b/oa0
fw7gGfuiglczU8SrT8+k9mjbzvA7uMvpsATXyn5At/oV0m6u01yYog+sEy7t
JxlyNpiSzbz3Lp9wmK1os1UQI4EUK/fnC0xNlhEh6nU0TbQK91qAhEGoWUew
OHhB0QU7saCyWkELNhwyAVssooKokl2qPclvDA9zePEHmvIasj2Wso0Hgge0
mCECwdliO1N1aN7stBNSkj5YUmCOoRPxZpyyYb/P0i+ah6AeCUjHqAeTwTef
LjPhtgqj9UZIpjZf/P5PJn2DHsj8Pnz+Z6wGkXGVl04BvdpDJYOL8/FRgSEQ
peZH58W5HL1lIj5kX/VYZ8OHTjJ+/GHuHVnKZurIMwy1f9fYjPhmeB2hRAS0
Q7flviTxvGgCWgf+enIFoiwSQB3eCh3oNpb8R8q579sInZ+Q0d9yilTnZkLy
WaS1o4c5+0RMy2M4juDnkbKp/ZO+DrVkAqrYiQZrrZcjWC21kD4/WVN0dXCa
IYozOWEQPQ6+q8/2FBcIQ3jhAmEDSqdKt4iSzT59FTXFgLY9GzetjjgaPIgy
GkuMJAdeqwC1p6ZbnCDHxYXiY6ynKO+IDXeut1mmMn/iw+/nC4vNiIGBvJ8M
/jvPf6iTAGqQ14FQp/8nkE0SCWvzTfytEsjnle9YIaM2R79A4uirwQLf2hDC
x0iISzKcRrL3MGbycOvwYSWzwFCdxnzh3HK9hKn2E4+NbZCAVkeIM9Xr9jmw
DVS3hmFDzz03vW7vAangERONhKo0NQ3+StUDEs1/vfpw8utkIuhzfpPEwqOH
N7ZWGCRuVrs8Be1pBoAlkaOfLLItd4WI2nCR88C5Dyz9KjtXmkUxgSkbUDiK
7giSVYlkhDqcyqvq6FmhYXkDkVWE1tKcsUBnWZwDKQpQkaJ4CtQ4nxDLSMgy
4Iunq+7fJmXa5cuZRzPYCRIoF+ZDZT4qJ1QFk/5u0KM3AEUqwe18f12Ni4hj
oq4/QdRutTv6CHEUnAyl+hbKm10nIEGcC26awqaMgy1JoWcxmRdBXJVlMGiF
9r255CaXN5G0MOSApTetrQhPpzbIbpYrn5WqkQ/MqQLo9Ky8Mh3LlclGakaY
p2WNzoNNYdB0JD8ir6lnxcEbpTMPeOZWZ+cQkphxPA5hrkdZhjhAbI5xHBwH
g9wsYK71CzEVH6TRSMKD6njAn0y+dPdfBNNuY/ZWx/BIjQdms2JRcujXO1v7
CqJnqj4TYlsVwVqRpwkfKDownbr2py59d5c+nSsXx/xJpM3yKrPBUFMjjSpb
Z6YiJOlFQkrItjpChTU1veXV1MdH8mCYjWFiZ9vmn8YihsZDXVfS6GbLTqOi
qGxiJoyRAQdRYe9cVQA3LOZywT1wH4TOEBbWqHI6ksSmoz6b+JK5B4gioZQB
ydBkmKb6LiKuY8qaUkDZle+aisTGpXoN3qdf211Lr9KSFqDewR+ZFHW9xA1A
rjGDdEqgwWpyzCsMrQWe2XoyAp77XK4LVTwLoahjd0gIDFQ7o0ag8hWcxg7y
Da7pawD0QnH4FQkjd179oBCB6m30lpWtWWtTfBOA1dFYrD1OvY9bKzvHaKUB
kw/7hJ6j3A3kLmqgpXPCvaiIL4Z1XJOgNbZ4nM/BdRQZWaxS0OkMZAyvCTPC
85MAjDDJRC0+USK0+aCSL0khrZey+FHGqsrpb25lBSPbPYQjDNlonSS8JcNc
IS833HU4NXy0Uzbldv51r9CQz/O4cpZw75o7Ms/l5ey7rz3gCZwVxghRHEOs
6m8CoJpXPO0oii7lEOqCSzZ6kH2Wp43KAKSJnPW3K3smaeXGy2UIRkYyZfA/
02rbHZ4EJbSt6+fA3Son2D5q9/4o2i7XfdjgRhBByHevRAAAOmigkcg1FMvd
AY0PDdvb3uwahCezLXzYdoTjjqwJWjux+AkvIGJc5rQ68yayYQoPa3LibOEM
ZV4w2a19AtyMwR1EWPdUEAD1+v5ACQnybJF8gQ4VkFlGuV8JnvhLoCJTc699
zN8vkJrkQBFYOBIbghtbHw3nzZhHz1H5xOpb2fZUGEQvhve/6nHUnFompkyX
sht8Fs8GiAFdQf42tb7fg4+TTzI3NPWWOV4RGJ6QH/EEITD3YE3uaXuTdBJG
4xu2OuJw8C5l5rLPJgxgwyqAtenCjwpE+PvP1Mh7kbDTHjaoiGIvOY6COS61
6g/1eXExLIBP1WW1+UHk4R2c1euYJS+FumjxVMUl9oKLvjbSnQwaUf1jxQYB
zBG0FMLu26HJOukzxfgK2v2i7QIXR3FrSdOumdUFdKh32gMtJAgSamEewAn8
FfEpRpE3dzbMaoBbgKe8a7JGR0Aes+kNSZC3DBGIpjMQvhfGfHLxZ4Ag3r8b
JvS/7eFHrtSi+ujcx8TGC8h93BWEj5NKf28e6ujklaBk9t5K1NJCcuzKfsut
H552OaSakBE1t2rA8X1LLjsDOhOfpkjW/Iu+4LG7HeuOmZQKMhbmyIbhtuRY
tH7YoYqGclxA+FtEGTdVFhvMCrThsyVXfQj86WwxHv4gn6DIZeQ8O/zFCq5L
HSCDXpNwhmDCGMDQUNjVhgHtKfCoy8BsM9jXCSrvwzFe7QKosYO5T5s6LCfx
8tMbW80FJdK3lIWKAoE48XJCnnqQbmTv5AdpDaa5pw7qbKBvIU9Pxz9wH0UH
eYg630GEzS0RWfKcpG88I5YYJCpmbZXkxyeOyobB5VM/FnZV0+KOagzhGq4R
X45DRkrb8X8zm00kyQODzmdj/ZEy02mReSI50fmYOx7JkT7aE7tdVq/xqYLh
wney39Ye8JoQzbkHPaY4A4lHqPgqfKJJ8NRF30Rs8xXK9XGAV5nMc7djfehF
090U2hqtSaBz1iYuOUgLfobFDkQvTMpVaTCZCu0848qOUCQDgiAAKNpAFx1Y
x3NKOl36yc2F1q7PQVFVWN70Wv3bc2/lJ9ljrcCe+/PqYpYkpLo0p4CRjgN0
Jx3YORqAUQLgTP3VdpdYEuEc4eowFyodP3+KGduq5GpVNSyAWbm6U+yihTwq
D5/cjDgcXGwWoW1jU+7WW7Hcl9B2adn4nnJqbJYnKAcSFrOOVwqkETCcAy10
/1ikS/cyP9Ss5rmTOcivy6Q5rZhuSGPYjqIU1crsxIGJTgBEjFGlH4Rt4kAw
zALWRx+Ti5wFHax9S/u7Y/bXBFcxYJq3656lHbb31HEllAWk0sMYAA8uFH49
0Ov1qzan1BpMByMqkxBohLMMj+bETCgRGQ1Wry+fUt0MJtcAstbCLhaqWX6A
2awZG+MLj6XsVPKiXWWIaUvLeCIVX4kzE4cZmR/4X6dfTM00jqQKIIk2+ekz
NEj0AnnIRkGekl/idEPkIDpEyS6tu9ICotA65qwDreFx8DXC2qMZIZE1bvjB
fxPplq0bQ6t7wWS8KtXjtC4a7/Xng03iZH37fEJbIP0gVUdKwtMAlVscMg+Z
KWTuztTu9Uk3AloAouN53DTCv9tqV7qxCDo2phvPOk5SfI4zOISqR5AxE2FJ
6Q8gJN3Mmn0ltkrWV0YEJMfPdaBImmsbFdx2ElPxeV9vZrD2h1BbmXQ3MKUh
POtcmio/GIEft+hIGf8pUelQ7BmSIP5jX0t9ayfX29WM13hXcI0YIBs2LOC5
jNcLflM4Oc8yytNoo5jbMAxWdVN8LthtwMDBK9KzA3/1k2vOyf48q26u4PuC
vUy+PzHf0gEVnVYXeZ3gYW1Z3IRwTe9X6SQHSTySBCzc01VCLunyUQ/os7kH
9NjtfWd0LOFmGonYFOKqja1A0T0YttmXMYnr/mOFpggoqXOFXlb+TDEJbQoo
WnFYjlvq3NB9IhZOfk+WTeHHicAlLTZb6pxR8Icn3UdZljvKYPxtWhLMY9EL
KDR4mUPlQ70eUEQXejdlbUoL3ns9IfmZLFb691TFetg2bMkKTgyrWXdRoXOa
4J7x9es1xEYBBcKkM0o0NkgjPRalcgNjCL+FYemPLTN3pIcAJvuw73BI9pYd
53CaTYvI36gzyxWkp2Mk2XDNef7zEbSeBOkRsHpI7Ox1gBt5N+QHfh885pse
B0n4L5ex4Avk/ndoJt4QdnSEpWMjr8lqzTWQSvtp1IZYdaHyomlE8d8LFrLr
f1970bF342UdfHir9eHSp7o2x2sKQJ/tQBglXN7ouYAdHyZUxvmI9dvInuLx
dHZupNJmN6iGzlhdcpzH1x+jaXbUOSzGEAh+aogPFdw/hZmMaPEE3pFlZHdq
mGh5xFvwULIiltYht/k/Zs2vjimcEnhQ77DJyb5/wGuOEB5xfvhoZRXHYwW/
Sw8GSXfrfEzTBXcljQdronF2JfbpyOTDY8R0t9+62WKd+4893t6Nl5lCnV3c
zK7mciqVcozSGDpGb664fxZxgv3w8vIQQB/tFDDaTMLSspknjvojR9IsZzwP
zCFzaIRoxYsddZV1SiKuzIbePqqftvz7EIH7hnwUf2njX8UWIh9hdKkAcRKb
GQXrULHKKuC2w5l7TcY4iUhH6R2JMFEYRpnHhloUgZGUfByjxwOn8Ydg8FeV
/qqgcwkCXBabmXmPTZfIIIxedLfA2ZCRVntGzdWupQGuZAs6yQQhQqBtEl0v
wxFFMXcpKWqtKzAineW23iAdjc7toVCt6751M+FmAFUmhezG+Rczz0caUCBl
rHNd4/3FadxO0ykCeKj3tIjzYQYKh9q0cv1gbgr905Xq4e/24YOFKcfqM2R2
EG7pfDskmNNLiTrCs2P0CMGhfHis0Cv88UzUBif7OTW74YZchD5+wEP7yMU9
7cru/ZDvCUYlukEG1FPMmxNbYN5CCKUKPJco0OiApABRPB3MzsYx4pYpLd1/
hB8x3iTElkaHuj66HceXvsQPU1FU6X8llwvf8eret/q1dRmIVxe8P4qP432s
FCqVS3Hzd8nqI4L/UzX98pnnFJuW1EaGDg2uhcNCfaGl1T2OvOjVofoBClvh
lOpudq+/Fp6pwv42IvJ2EwS+OwgAVBdOt/lj32qsi3U3TGaUkN0LdOY7KSuN
16kI/S+jJyumuKOkHTZV9YCUE2A1AuKMP2AA+xp21j28fvUEgXjb0MJp/FD9
Q0g5Jg/JScebIFh6K7YCXDaEMSqMPyEBCVgVYK9W/TPQdsRGVYB3/u/HnFE+
y/dqkc+rWmQ5yBY3RmjtOF2muFhVxMmGcYm6OE5lToPJ8pGuW9XZXtNq3RXO
IG4ovMVT6I6RWZf/JAw4XBpp80f5vKGvzeSFpsfed/nDBeym8ghn2nVbHOCr
i8/ygATJpp6e9aiSpQt2ZmcuoBBOjY8+0+qZ2S6kJr5S9CFeur+AjJfvEEAq
YN2f8toawAeGy230iuXgGF0Fb7Bpi3w02pIuHrzeAkuWDdADcZ9pKhrNeCgo
lF1tqbCj3nUW/X6svtEIq0MLjpNKEYyvkyBdFvisU7P06PnVb5kJrnTbymT3
g6MbMGZpxz2+65GVn6dNzr4K9QOnZrgRAJcwG7z5C1258mgtmWnSoKaYS4pn
Vp3rBYrt5K4SS6CP3pgfZPUsy9nAb1NfQzbPd2ImUIu92QfTq5M7lia5ohTc
aSiikNVuPvsQ7UiveKJ81tplEmY4qtiFecbzwT0hkELedZfVtdRvGH39nYgf
/Q9A+uRL4z25BunJru+mfHHbTqTrf1qkaR8etkAYLitcmF4OUAXgDqb3SVB4
xiNchKuKW9LOVqlUg2HHnxalEfO96Kv0PYZORFaaEH1MX/NDYQH3lyUJQoQ2
189sIuRoPWR6hH0kBQEDM8knviybs9MzeZhZnUydkJPPegOp2UNRCJYm+Cko
h0aQV+KcU1Di0OEqYAJtN9EtWK4kq5VlR1D051bH7+8UwCMAixl93bAuFLOd
xaEXL3Xi/TsmqL90UlSxZwlF9P/AxUMx3Xyl4Lb+kdn/1SjkK6rK2NtFA7r2
U5PE7DYJ/k8hIGdmKsuEVMG55giK+IlDcfibyIxnKTi7CifPyzFE3JJfWFrU
CAmZqj7zDFMs8flj9TJVkV6Or6pHH//jdVAKOsm22M6U5PXubAnEISr/iXdJ
4Prr5MWBssBmrVQ3KArcUMTBtKGSXj4oUDj8lWWW2BvVbhHwtTeXeVB0cuwt
ZySv16F8pO0f9nWqUFykFrrrHM49jWGjyyDiZ8z2a/IuBkNdkhKQV0oL3GsJ
MF5g6ZqEYvCz5twhSt4jE9Kz8FOldUfvUTOBiTK0zM30A+q8iV3Exk6NTsfb
pX2aZfpCR5ujM1a4+3ldkBwBtdDFqZN7WlAX3uMYALk9tGwNq1YPcpevLo58
QZtzAneXsrr5sr9zzy/J1wFEx+98jrS0CSu41F2qSDKkIYSG9iEsigUODkPP
F3METTjPJPYTlw5R2I92T/aTljVf/iZqmP0jGAcWqVD6VEkkL9RKXY+h78sB
+Pi94SW9pV52wbci6VjiUoXFkkCIX7cmYmPlfNosi7kSGTskDz84jMEXqaAp
ArRz+J6bUBUSrZ4ZzOqiU8zLQYnSKz3W+dC59YTDSfU26B3KVIGSxcOh2vFg
KlwVUaxGsDBYW4x3/h4cCHGu6PcRziWhLkFh36bM6JM9xwC6STbR8d0eFn2X
q9caAbTPDtuo4kzUQC3rDKiz26BMciv+JzF6wjpLERVtDrAiAOa0yHixsrnW
6eTy+Z51UG7lOmXVb4C35vbcS0A0n04IdzK93NSLyuhvl0yM6xbmrXCF+Fdb
ZxVURwZLw9FMXo6xj232eB+lJi80ch0k6pOGNX3fSUvF2PSLdOqUVL7GuGjp
HIGz1iZObeL40fbLyCM6+aaeKN5BMaPKIUPt3aA+0McHNE+bzMVnPbZ2yzfp
D8lUwDP0u3uM4nSLyk7pfvQGFC1n73WwhPQSzSstOBEycvQlBTqMzBaIdMIc
2QRFKmkQC5UJcVjtKWv47DtU+oYT7eXlaQzt9ktjgdbQ0hwEjxJBlNH5Js2y
RBIPBFhG1yDXF7JsSnfacYhb5KOmoXhJ/GcI7PIGpBO2Xr76TSaEMBy/bAAU
eqUbnNSFLmExIqjCJh9BdlyrQ5Q7G9FoOsTVe/pGjypuYRpVt03fVOBsSvCI
3He36LoAwXBQ0zGH10pW/vGjkd+f05JwdgHxw88lb/GgkucnBazTUcmPDADP
GE5njKY1/d5jf0GPwPBpnGiQ/cKlKEnXkpUP7jRCIiGds7iqY7XYn8lYmySR
T3P62rSIt5pdRugigvyru80Z9M1GC1czZs7/OAuwHn0uuKtynPYRVwwY1Bv5
pGVKnl9064X1LMWL2YiNHDYlwggw6Nbj+Q/h2sCyWKNsjmIzfJq3YtvEK5Sr
1nnny51nlPa2H3jjgPh7+AAWNXxrWCgpETnTFnprM+G0zOWJnCgUnvDDsaUX
kwVaJ3iDnlTVe1Stq4nlEi8o0ffBPqxSPWu3TWw7vCbvnCnX5ZS8F7XvCMId
Ld3SHtct5x+ZRpqDMZ+PlDS7HsVM5HQ1qOoePGVPmLygfMZ86m0eG9sH1McQ
zuc27Wn8m5OiCsf11vc/HqdP9vI5IuKHSWtExZEyGX8PqHAslgwxyNI3wNBs
jQCk/4+o3FOUl82sjchY3k9Lt+SFdu9ODCKsHPjBiO+0UJG/8uZ8C9ogicwY
i2CpdXrXSksbKj+AoJrMnUBYXOcY4bTlrPZnqUp3wEvAUtMY7vY9z/winaNw
FMBHRIXrX6C/RNOt5M9ESMMTrW7hHJFgqbD2wuZ4VMzkDN2R9Ik4MJKPO+XN
j7QvL3XFupHKgEwYbGKSZahTiLxu9dfxsqV455EaqZluMGDt2WxqipvSZPgY
qTETirkfE/8ysX8OvRXoK4/YidyDh5Yas4wnJiFoZegKZ4iKA4KtsDH+nMmw
3xFE6AJH61cX9PueH+kDERJzLtj9wFPTlAffCZBWhiepYfd70qZX2lUaRyNP
VsCZABernccjXiH+Xt4P60iy6zm6FDpkuAJX0HahXbpHFpnuCY3NBiVUGhif
21eM4TGWLA8/9ztUGQUwlNFCQVxq76tE9hwK7W7QuHU9RGpJ9ziCGTOLBdB/
c6/a3qA32vDtWJuSsU7FHYTYaik9RCIqPLuoENZimanGpYNiJ61ilcbKaHR+
57lrsrCx47PYLiAUmyhjq74pj1lzKk504iyVMJIexm06EO4j/eW93nnUR8IX
eiOeS5urw0pXQVLM3MOxW8AXS38ywI7vdN+2sN6/28i+J4Fx5ItpCjJ+cRRV
JFmgVQ0+tXoDPvEByeoy/rTXu2Mo3CO+iM41ptNv1XxC0p7v17H4SFNsYAhN
nEQJF1JbkdTX1iBYWaCWSsF7PQZByqIaGNsV0w2JUHNnkFspuGFq7tUzUbNu
ssV9AZ5D9iGoIqQR5gXYbHDdvhtHrx9u3mqTbBl0600gQZ/8KSK+Hbjpk0/2
InyGSJeoXzydbL7qEwW8uuglVh5RbvPtEi+gXR+z6hxEmVktOuIZNLl5u/N7
7ef8coh0PoY2IkNTYTPVTe4pu6aJe45ueQtgwfAr5rY/XpmQ7shDU8ELyQNK
UQVGBOpj93tPMjpv3OnDrF2FqLQPfDlyjJfZg3Ymh5Z02PeMYsJFdjawm6be
T5zUohCxX9VRTQqtndpHPJ1Xb+c6EIN+HAb6aX1s+3j0ardQaMySFWiT8WX+
QLGLAtTgNXdk0+6XKQkxjF+74DeuGTYhReUz1LphviCNLGdjTPaqYp9N6Mre
3vpt8svvgeZdFVEfvVPiSQTaKfpZ2Qpv2J8cVMyEfr1b2hFx4F/pl86m0gf5
I9Qx1T0Yrb8DKqXifQpTV6lA+Jg7ZxmgeDvIc+X0JEp3LxCjbR8AyIH47goc
9D4IFdb2t+ZH8RsMDNlzGP1HwirrxP8iEDxmugGSBkheRkR6QPyGdypeHblW
fETBq4oVg830necRnrRV/5FJHO1EE/l3fGjXnX6YrtrFeS+VM9g9JAQet7Yg
fyP5La4guNGdz3g3zAKHxrxdfTQyEx3B0AVuiFvBS6bytfaNfpOqhp7S8arF
F7+qgAha39v4FqeBmVIKdai+hy2ZE0iPxYs1cpwbYEth37UKRT9xStEvM9xX
k9VFqX8VwOA+uG2beX9Rc2TlsBmJgY88y6Ps1pPDqzMjKhGcbXsizMsKTsQq
Bh01XHDjUGg91eaGtYzQdLX1MugoVObN0HL55wFisvx2B9GVSveUVjGZBp51
YXKZEIPcNh17IiBQ3bbVZaZ+WZTwDl913kDM7k649+3+ute3QkxP4ztFikpX
twKH/VyNvSyqJ6qZ+DqWI5AVH5x8cU1dDsq8NkufmShlpGhZxKyqJRpEjhxE
AMxAYAwDTOhjHuo7HPqSNfsDeM7G/KLcemqJ7ge23WPYeG3G0PQ4ncL41Qlz
LZRHziRK/+NUGUeNPkJUwVg8nYZ2yfb9xe/V+8mRyRsjvT+Dj3AudYyd7nA1
kVgkP9j+4yElz7oiWq5h2HQMTEhm5lRRCnselt9oFzD442rs6/6G1OXgfX1X
mgVpkMhXFgl0IAuFynR9SGEoNdbtnUEMVk1mnk+k0Mz4SaWs/17t2yIs5QFf
9TW/c5sMaG653dveZQULyT667dV5LN2yp/XrHk6KHL4sjWOKgwlowz8dowj5
zx5iRIcZxOa9ixW/XVDfIJVXD/I/7A1pxcEgk8zR3FgXmlinjYp6Ucr+NKTI
4X/78mYhtzk6bmMsVBsdkRTyseC//a6BrEN84zQJbDaGQ6xk4geIV3gNUFOW
msIJoqeE8pJqnBPtK1jYN/3XMcLgbs6kHC2+ZOkUlaZkFUF6iniCaDg6xxfr
rPCSN7dQLMhM8iWYC50hLx3kdBPQN94S5kNrazrUNBAzd1lz7oZSkuU70Pw7
GhVeF8oYCZKV1KP1sGL6Y/DmN5BjX5yPWou3bEZHNP6imnTx5XRoDwZiPN+U
PifcxYxmQJQ5ybwAlnIGtdiPhtHdLIzxnN5oyLeISLjX/fFzQbgFZsnos8Tg
hNMLvAomoooyL+xH2uk5sGCnx+8jwJr4/avJDRl40viXkuF3pE8uWrnDPFOu
Vp4Us3Qn0kXPEaIUK+MEqZbAXmPQVxuCNdfZT0xpuCq1DvOj9b3Jp9N5yFu7
byHiVlnNik8mFhRN12+U16//Weoi8CmTcQZh/E+dB0ldXVMRG6AgzYKKhW6T
3YNds4ans+NAnPuV68zMHa7TcyE2f53EyKiQa7X27HPbb5g8/XZK7QvKhYRo
KszJlTtcyTFJhZoigXv8OlyQP1QZb4+LoOYiOK0us0FVj/B0xuYzxyDO2azS
v7CI9ijI6pQWXRjcyK0ioX30e4UcA6gqSbZZ+l/YHpQNMHNycesvtdrj3aPV
2HqDv6IHaqIasIaU+B0FacQGSGBVSbbS4u0vubd3Q840c+rnwBGbqATWK9ms
gCNHi8MRF16A1eVHAahd0MO8kF7qZm5w7NgKRN/6WST6DILw7TVIPE0D+c2O
wiJw5f0uWN1BmQUoD9+V+cvYincPs1wBciZl3WbYsKmCG37Mgjx5US32SPS7
mRni8pYR4SiA98a87v4qTPW7efRLNv96P9bDWj09oC/J/xAiKQrpfrPLxn7y
+D0Ul07mlGzxz6SCMCw7hUHoEGjM+Zekvq8Kn1YBQCX1yI3Yhmj4dyPZaFr6
XkhY0gQGAfhhVY+SGhu6u6QyAmUO8Gvft5yJLTAIxu9BjDect6/0/GtKLBYw
GR+BIeT1o8fbaVbbnR84pbfN7MKShsc9BrcPeeqc0FNEBo3dD3Vrwnbx0hE+
z4R6vG+1D+rq4bKe/8RN9DHMzSG1fIxhvHxwLkPF5WUBNvghtkJ3747FZu0I
zVKowE8git0KcXfZc2HS6Z/9BDXMoYbc5KWtVItu2XoDiRvvzCCtNLyRZiJP
04HB5jivbpFYCCyUUtcuh71+oOfHZXhCs5R7BsYVBGfLGVJBnYz+JR4SSREq
1jKKiFWL32c3uyv5v4o/+eAG5vYHsDAWaKpAru5MvCy5XFSnJHrA+ZsvAhZi
IYMX6aDvgftaAjmddQ7gJoZGDWBH1cEKyWQKDpVmZvxVbYb6tZl18/2BBy13
55MWNcaWu133YlxnBq1lE8Jx7Czx/JXEE75+iIuk+KqdvEa3QKQUePKd59S/
ib6ghsbowqvzlc4Nsv4bUune00o4Y1pGMWfE/8AO0aITxXlO4xnZ7GS8RJVX
FG8RV0b4TAcXXK6I6eXcZyYkXX32MPJtvECE95Fdn27Tw6xSaGL0P0X7qT+n
9mBBAAABuQjSo/di4u0U0ihRfeV9/keqvYa1Hj8noC/vSV7stZ7tMwYkcq/y
BiMcwYa8nFLdhSEzjWYFMvm4vSbgi1ddDUxJl6VCjJnIQeVvLUTMFwR9OUcU
hfHABjdeR7qzAFCcA7hLJ0firC4OoxmLqNnJ96RnQJPUT41eXPGRLfEVpvpp
1Q2tjtAyBc7z9ia49xKNWS9Z9uwMxO+jGp04RFJLZGawEIuSqjN1oXWkK0Up
oO/+4kEE31MEpWRDbIKOr/Add9eHoYT2TIqCIIDzBlQEtpMmSynMYG5odFx8
EamAgUTNbhJyjCqir0C4W3YbznmlXe3iTAXf0WK6EnCXfKvh6YC3XEqb+3aD
939E2EZu5WU39x5nWORvEoV8e1WXavV81dPYu6cUdNbkFyGtEO8WvqaA3ZD3
cLvm5UvVMn3zvYtDGeZAKBByPghxC4cxc1EMOBRViPN9dTI/3Dtlvn4GR5VH
9mrJoCvdCJiQEosjMouwNPBMzkvYAIO8PiArns1x2/cR2xGqRwNzRgrrUY1V
CDcwP5v7Rkbc0kDCHQd665/gs4NBwu213prWS1C4IJ55znSuD6v39esI3xEs
w0+yGtOGqWQdAQ4rulWV8ATtz9NiNrbIQjMSC4sHCgEo5KGuu49YgaO1RIc2
/cnStlmidMUisa+AT/iNFUdPaQ8fd4auwJuuOCXAAy7NZ8y2jlAYsmxUn2+l
ZU2cSkR/LvzdyHQZn1RRxOo+ZbNz0ZYMOurX2jM1OT6G8AKNNCu2SvyirLF5
z24WRus+MRGy8HtberLhayHXaUFb29cp/6wyjZKXwlYVLKrLmuQG7QHP6Isu
jOEOGgSmwKJ4d0FLwp0rCLrC3/WG59kGAUnyD+KaP3/75TrKyOwWi9vstBIe
mgiAN4rJypxsT/YtKijoYCQCHbCamljfbzeQuVlMY1Tl0mkrbtJD3pCP9raM
fIka2E3t5USqscFDjcgDSou68I8VNHJ3gAPB+Z+lFKWMHvgsUxPRWeln4oFQ
pLzI4XhShBbDPSkVtxiP4Wgx3MPHco2AkE/NVJjtoKDhUkE38VxAfyyofItj
jCRdPH+3Ly3Lo+GORuseylzioMzl52rSPrFO/NYOwVnYZUnq0F6vAHmWXZrH
s8/ptpqhQFaB+HTzoCSCju+ygc6wh1NCtE1IKja6yWiugIMcg+pD1YgcA4Pa
9yHRQBAJPaV8dgxqRT8iTNBdMftFcGB3YujSPKN7ttaEsXtEZEo7Osus8DCp
xcexUE8xVAwth+3P7hVodMOflHKhpWMDA3C/t4rX+Cyo+gmhGXtfwx0vADmM
FUxvzMyIOZp5j5DphzmIgZJH5P+VZLDgvMnmQHDTWOOU6vwQi+n8DJagOR+s
iAMwICtvw6BOg5pEWerxZQR9Akdh3+Jb/Bj+8JvJ4Lboyrl0PjdWm3EWDoq+
5eyUYagmvI7vXOdjlHHk2qSNrCIjGSSPAPS/hoONzUOb0GSePpAwZxbhDmpB
ntHXpVLeBsuWKHzTMQdnG+Ks8wzJtmyYW/VMj0937itAbfPwK8CgOeW3Zw6S
z4+kj9RFF15Se4Cg7x5b5Hzljsn2DmALBEP8bwu+sJzlGMd96QsuWbq4FGrr
15Cr9sPi6rfCPr/8EPfjYN02kq+rsY9D9woGb8rEHnPCzFNHquWCnrvZRKch
jO7I+8PZnJ0mEcwxZXM9FUQMuncHs0553pawzw0MioBAKjREKTsiZ+yWi3bF
vrRMK1hX4aT3Z4Igdux0Vm1ZuqVxRKwiGqLvG0EqofRrXfp8seXx0mvgu43O
xZtBWPOlpMHbrDfZtz1GX7Mxuts92h8xe56nzEIQ+8ax7soV+NXkwntxT62o
/zpC/2shRHEep5o/1aybp7kVXanFFIkijpD4khJhMaJjpRkE5S/T84lDl8Fe
zwt4OE0Pk+Clph/APRm7rAKvAcdTv62zpOuehKO8U+bI6/eFWUXpMV5nmM07
iIEGEaxd99rrLjerNsH7e/DViykp88db/NjySMhz/uGwH19ewKWPu1IiKpvX
F6khSYHYVd5xzZqhKgAyE5bxdTtTjxHHifEWYav4k3sZNb22dvQEG8WZMvaP
ZgxOox92bvR/UB7yPVJHDzS/Xlvf4VKDRywcMgvng/Ge0oOf0fmShd7oJegw
HiDHoC6xif3N7LOIEjc05gskRttHriaS5Lo2nm+Wag26g5dmk1zJ4p1axOX9
8Sgkhb/2Tq8i7PnE1ix0x5KaT4T7OLzZTcB3dtcTmEwGYii9A56wLDvquuLD
TgLq9IhgPTIJG5fyaRKLcun+3daJOsWiL+np5ZerA//nyMgZCgVAe7hZvw/a
H9e8+LwxL9tzqzIs0FrSGw7whYbAT6h/79YrAZrUXiUC0lfQeJIl3BUjXCXx
/8eNqjGjOEzNd471PCd80EDemMU9hHjreemmovhY6ZfqYbSnQFO0EpW78zhg
18Sp2TY2qbxlJd/ezv1EZwrVBhPL5MhzVr2YtUko4IhoMl5cJlzjtSgQpJzB
Ta58GZKHnje1VKAIOpKrNOWtrWfUrKS/2IWT1HcHcyqXygope9JMql5qh6QP
qHWLFdUtb2G4IFFYoV+p/Nd68DOsrkTeeJ9O1cP/dk2cdXPRFrPrLIjEMQvB
x4aii4f5Cbs5td/kZqptbmFXWFRDnwaM4Chq8KSWokKOKxFhak19iTLpUweN
g4HtJDyA0orlyitAmc15u/mLBUhsQw/m1aqcZe3tdCK0ojeuqg0c0A67qj1p
8fEVtRtfa5CoIIHwvK9iCRm+gKefp4ErFB0zMrB+q8c+nJbudl/Uc3FljE5K
M0BGeN+xcBANPV06ztuRZUQUpLihMto87vXA4ITH0mz1Vst8lmkyI4+MileN
W+5H/AVQCjdVfQV/ldKbrF/uFkyznHCksFVTCs3ibgJhDMQ8k01nlzmNX+Xe
jCt6ZRJbPg6/4zbvFpiQ2jedLuD/yQYd4wMLoUjCGDMsQ8SmJdeIS3F6NanT
jAEGh3+4lLjBgafOYXy1v60/lXIWybp2DA6Z778JTFLt+MQQuIMMoAndLqHh
0lhSLbhR15J6KlDtpNiwbUdQZz9YrqUerdzq5J/J73xS0Ly6N0OtwRkS9Gil
lH/03qjiB/Rypkb7x6KA3LzWzjXKyuuZm3cdYqMJjdKPUSDCsXa01M4hfWNZ
WXQNP5RmOoz88fAQX0vWHKf2FRsH0Nd/9Ph2BMztHcDIkGoxVnNOmKRkqhuX
Mq5EUW9i24B9pji0ZqSdHb6KoV4MdLbCCifEUxfQZl7PZySlqN0TjTBR9SFB
06eN1Xi5KNO8o17ynYquSVvLwUiWnBcDaa6tXFZTkEMbrPu1DdtZiFb6CNJ4
ufJTcm2pFkxSXPjDmblgApnevUxOoIEK4VLlitL5KYe/VDWHYaMvCWmR8EkK
dC3ZrZcQSo1JuPj7goOrvrFLnv3hsn7sKH0TZ93NG0AHzjakGu0/s1Z0yrL5
QvuRNt/QrBPRJG1UMNZ9bbTida5Gl1+m115U2o27BCbHiVUESpvaiDlexehc
DM9zZKsyhxhk75dQS990Xavu++zIv/ppbV3r6mrljTugNpXBrrKUJcXVkzfK
Vu4nRP0aXZoEVb6S47GyTizjuE2LRf1hPwXbSO+uSWZv+ervovazrx4KNUPv
9ilnLiq2gvBHnYwZc+Hcy3zvmn9WJH/BJJfRzfT3pevOhcUpERWXnLmJKOv+
57a03DDyQRN80JdwE6Kv9Rtkhfs/5bhz/Pjruzq7GyMG3M2tiH+veOXLeA2C
Qz6TmXHW6tfiSHVBEXrj64JnI2ZZoZ+1yjL6KB/wMTP3twJRAWKc6wZ9ckco
UFTZAKvQFDI/l26ErWYuM5RM+HddlNLWAd5QpcmZE1QFnnwKCXb4uebqFYGQ
w0ouZVxSLuOIZ0Gu6ikqscO1uEKouaig/H2WbwhHYlSiZXR+To7rYxTWA9aX
VlO7ivNNfjF6gYBYexCp34bc4s67qh/WgcgUI4qr2n/lZNPWj6v1KWu7A6tf
HSk5S1QcQp5ToFSXRF+VeTV0lmdSp/SMPoAQTk+d2dA3ao8sVCPVssecKVnh
1Y88YMfuLk9lnrOaqKmtUXoqfXbF1PQAE8R1PI6z7K+SQBSut5R39u1b/obr
GNrSTio2/cENYmLYqv1eJU5DiPaiZsjJUi85K9tBvjXKJqi/5+eVI32iZ6An
Qfn1rYlLiR2933S0TSn63d/f3zL6+ANt6YU0IgZM1OxYAlwnbHhslE5iaTJC
1yvYz3ESzO2x6lf3Yb6en3uVISuQiUtMJ63iIXYV15qN9j7Q0coXEjoCeBKk
07pyA96b5LQ8CsyPo1wMOU1v7YoSHFbByyRFzsR/bXJ9fBgQwveFXnUthmaP
u0W7uTxG3u3ULNHjo/9KEcCX/wngKnQZMF8aM+9a2Ox9C+8kmGHL3m9UwmRZ
2Ukv+Kegk7F6kbe7T6BD3XdaYRQgAEMWrYJ5ab/AMQCPIKvI9NbeNgAmBHkG
ioPxhAZKY/vDWjRc20aq75xWaUZBQ9spw7IF9QPhU3O5GDcdSqGAoCJ/GNZI
UP7r0AoKjxv8q2bOehXXxey9Uwcap9aXu9HMXcoqkAW2N50Ihp9NK37CT4x5
02O/JxzUPfe1M8wZEjnntjnVidhA561NZ/WS0A5CmpYRlwS/FMHYJFnBP9/t
JBwhOixdbmeYfdrcRxENsMwBq3KVfOhscuDSDANuoLe4F9F+Q0SiN44Bzi3B
2j0p6bdm50Z4oKzA8kPh455gnHBBB7uY3lrtNUzl3bC9XG/AsMDG6t2V3d00
a8Tj6b/TEkSTOxNFNcN4X/YaEvhSHMe90mWheJOo3EGYAB/eaFfp2c0GATNY
MxI6vtrvNCSIxlw0DzygDz/1BlgzOigGkiS/EKLmBRrP5OpAw83Q5lqLDBer
3jxVdXaQ9Zpi0hCtvPkmjliry5FOvreBt/jaBqRXUF9GCWhjsj3EU5EG1NZg
9suCo/LnTc91rdnLB3ppdH0P12ORsiu32ERRQBvLiX1png0bSw9L0oMNvU12
0oMx5nIOkCzw/7uipXkSLbZzVpeb02ImxJrI+jF2ioNhxtBOM+ZVOvox3BEL
8KUf5hxaHRW8P5yxWVrIHd0xJDylc7xET3GjAnnP00POhGk+zenV1TMdqUeH
5URL8mbTctqE7TT6GKAM2lQzvkeK16AWOpXrIszTCYdpP7IgW7GuOEMTSJ5k
Ttj9PBL6+NgVbDHE8M4vTxcL6DZokP0QndTzaZ3X/Zb4dWAQ7VSesHSDVqcv
Je//hpKpLjROD3+W2qSJ16VwVZ6/y4/dZROa9ZJK2ZY2A/iLEHxuUdJH2wcQ
yEqZ7CMu6CHiKq8TnCkVAYnTo88/lzqGycKhf0rWI2Tt+6PU1f0S+LREIswa
94c7jeekDGzlfFdBYcyT4rHI2IqTor1essZ64IzyMLEriFfpLoeiFs+2dXmZ
+oD0EWtiUkUPmSdCNak2E4J5DnEoAna6gsULUlquYPfxsvS+DiByxt1j73Hg
51/+CFFf2M0juSkbXBzIZzlfcucMOIi6TyDGVpnvyp1VL8G2+EyyG9T5+kij
eBIiuHt8Gr5U6zumtMa2zzYIoCHTX2GgfjSxTU1cmiRVDhPAS/a4SXpS/WXx
ZaCGK/wy9UAAFY9J7ObfuzSH/ffRUV7UpivYOSyFWTzal8YkOh7w1YCcvZwQ
JBhxCPCIA6AnNtvSBug1XKRshGzWn1pCR3Q9xEYuW3On3fmxVYbiFr+T8vaA
mMaLKU4RULOFO1HVHj52vZaMrUXwJq2u527wYdhTpMgtSHC6MHA9fjAGioL8
jmfzMCWoyWIGMBI2lY+MsFxoaLoxliagjUb9tl1V4em5hvt6CrR7HzaO6lxt
X86r8oTRXizOlmljl63p5ihfC6pphbzozIsvPKcvZHogw3Oci/BNNWcO0JEP
zjUSjH2hfO2L84u1satY90iS/7JoQlkRUihyZWC9V/QmZtRMNEa5ygHJM2JZ
gSwbzhYg/kwTpkYtRhlBgyPZQ9YG6H1VhdabIJJKHMZkj/tJ95vBWidHr4Yu
4G0kXkHyb7oi+v5Va7ASAFIS8+LmBl0XhN7+zCMME5T1FMkfH2WJ5LKCOJc3
pfDvceV3ivk9d7blyfiNlaxRGotflQ0MXMO6aTkb5FYdHXelX2HKwOYEfpLL
qqpdx+ZU6WWeoyKp1VxwAFyQbnEf6qmLSo7GDfZtalOOiwOHSYgZJiSXCxBd
LBqJL7za6dHlgyUzoa59kZPGfQXt18vFkXndIq2vS4HSoIU3ItMLDikOGsey
C1Rd5Bq22IXsFRLhMbo+ZCk2nsJoSl2df8zcLHF34SPzMyCsVRupGMqCFnLQ
XwedlYMsRK9D+FeWMp23cwN9n2yXDxwQmnlrQCvLnFi1amRmmSD8XTJCrxaR
HrbSCuJBiUTvkqpC9d5wkx4vV9iAqlwv5AqK8xLTcWsK0o0xnFOXjY6OFaap
ny2KqpgdVoOI3ljMs0KAEWpA+jaCxrdTlz4eSFLE9HVzHX8AMFTjfQqmfSXu
8bSvNlZB+Vn8T4pEEmyuGhwubypuL0crxjLva2nUV8IkHtxj3ShqBRgnGeed
FbP5Hgr9z1m2x11GmomVTMll9eUQX5OvXgx6ra4f0ILq5gAKoeDfsvuX9XFL
rZ0YVdch8j+vlpN1zQCIPhKi8q9vEa0rduJYQnax6Q6YDFGbhNfRyyRhgrfZ
iLjDnCw0D88LAfS+IhbLANdBkUIjJICd2TQWn2rvPT3Y7pjweojx2OFFdhbL
rFs0sTAO5/wZImrDEOdxbrJS8e/eR5jrVwbXwL8Q8lx6236W8PaJBivXNb5g
SOTuzThJdDnyz9laXYxDBLOLSeyoVoEDhypDOb7N1LAl2jXTIvGZzCkV85ZM
96RwBT0NHNwACvDqVwJdM+Ahz3UJi4AyoPV4SzLtBK/qZmhmwObD0U8PpWAt
z8n+XOhswsqzjyZYkA+0utV1MIvUFMAQAtziFi/b1WUmRMares027597hU3Y
+VjfZFpZroz5Z9BuRfhqgQODKCOQaQ8yjReJkQVunGDJ2d+GEVOtmfBhEcMe
5wx4jVlySKcE+BhPfA5SkIJ4VZpvSVdd6feJvmJxMjDaaOfVIaHaiG0zf6Yn
NEq0BpXnvy6J/j0PL/BE96fvdL+fSl2gctvVXUrTq7gKYTp1k2kupK1fves6
qAUE3O0xDb7kUPoPLc/qS654i1ExpqwDALyEDJARaublCFvUJnbjjY7UzCYD
Fb6Lm8JkkJgO5XfdMU9c0NPH887/hCx+zhxhK0ofVcOyAi5ssalCII/UJxMR
s+17wRhGtaQTJXvI3Iu+iFZFlMJgEniLhKaIRpTQBsgtUCqbMWaHsFgHWdnj
OF6NJZOaxZryMHnLo2lXm8zdiLdj1ftLj7l9Z+wZWR97iHjbqbOygtHGD0tm
4sw0MqU9f9Frk9BLwn/kU9mpbq75O6My6KO6pdrcHT6yFlPrMv7Vtt2YhPo6
kuhCKPtlkWLL+Ccuf4oyFwTdORYKsGuDSMw624cx2Ln0wxDxXOzEZ/m9shvx
qgXXEBEyqVf1bKBaV/bO1p1OndUn0tqLHQ2UU0Bmt5PMyaMmY6Aus3rTzYS0
IzjsfPx0PqymIuQebHYd5pPGpArKG7XG2FglFGBsgJ+s/oQbIEy/w0nH3PCZ
JwekBrGwfp9QhX9kOkOWTLLAQs+7W56OtWi6QdHe/8Dx8V3dtaRqxHd7uWVm
eMxgNaT3vijPC/fZ/CnvE//pNC95RLBy7PMdVVQMnanLdeIhuX5sWVhIIB9L
OJOvRyV8EhZ2MvrZv5guOQzL+sj7YMPGJpO5lAo2frMjEXpNfhxcCSg/pBKN
cgbOBL5AA9Ust8z1ewaa5BahvQmluPaccWqFEP0r9Ygfb7qGgPsp7ynlk8mg
J6Hn1xHutD+wF3hONAZv2dkdQ738+vXQm7iNyHVhx8nvvVESbNk/K98tvezz
RNn9j7N8ggbqYEne6u/zNVq6tXFchoTQfnqvu+wLbBB/be69jDvEkwLD5x64
F8QtWDJXKTqipsof3JSe0MP+YkNw5fCRQnWgWjOBzGhYzMuhu8ebO5bj/uFo
uHD6uK/yzTanqVOqEMBs2AW0JBfld1PSkEAgG2SmJmnPmEEJFYMLiQ9WFQ/O
Q/2Qs9PAIOqvEdGJy8M1c1Zz8Tt4lcnTuJ4Km1eZvO1x80tQAHs36NkRaL2U
AFMvKPEvbI8uIEvmgXh4QFO8+xK69dhknA6mCzDYLTsKl5m/lbbYArSWQSMF
GZMd6BLvSotdb962lZLtERTGEHMCEZJnhFfg14X7bT3Vxc6BcAZ9BfWmY6NT
cNfUy4/QlHaX9B08o8B3fJhYox0aDs4hLQNhwu8dMyyAT8Tjn++O6YgM1W2E
rFswxBGmKZq7oXBVzlsvt6v4sLb9qbWTmvPN2bzL2AKGWo/B42jeOUN6H65B
PDWMKSUcIZsQrqdpG8dWl/+KUGGsrwHSrwhTwR9srfkCLaPOKb6RauI+lo/Q
ltzB6mQZash7FYfrXYYz5VQ101yhJTzlPgiOYlcjnJYdFrK64dRwO4HOWxrM
tTo3ZyBxZZR2K0y4wV4UElUR8k2NBh0FtbhO8IUeINC2VbwcTRdBocgpr3vO
SblfvKIyAJRWrFoca8hM1ed8IujlnAHkncNoZYod9Kuf+R5sWGtUnvOUK9X1
acufHAXNctaYZrIvs9aMNBmBJ3FPm8W0mvYj+lwiG7uI8QuiHyImrIoXOI1s
/b9Fuf6hlkHWhNPXSfCYv0O6ejauOe1L8Z5U40zo5tvksLcmYXguYZ0wE4YB
zm+mBbosHqHkXLAdmCOJA5QDctJHzATCZzwmrSCggvnoRmeDuob3w1zsZEuA
oHMeruPDxJ6J+drhnosAyaQebW9FoY4r9fS5fvDHL6stRdz9S9InwaUuDGbf
g4Q9gg5SYuKTfzivdhILuarnl0bYS5CO2VfJnMB4+SnkCm622+n4fK+7PURS
mdAwUclPnqa+DLT3g+2o2RBmVR95xScLXanx/39rjamlj1h8ex65NJXSnI3g
qkx1BJDHrbMuzwHZebAoZS/Rhq2UsL8rI3xK0HKuRX+KzFkt0zNlvHyfGMqH
qXpBWxhg8hK8pJlCMIMTOC+L5Miqaft3f+Tt7H5dKSGYi2n+GXAJ7MmZN78L
Z3deP6tbRmm28km+TgYBuYRznDgieKlYg0LojFoLrqAsNxvAQXHSYB+sV+sV
GeYRUSQHKjtIBX0spvXclp/F9AA1Nsm7gA4CgMoXF2L72TuIxmEaupzOwr3I
Rx1SjhmjlI4TcLjb7XWLh29Y2K2Oy7xDnmMuJEzBH+86sX6bych/PvSrSe1i
8R3uf4uMdELmAPqCh53t6qcYihJTQM400DLfCfhT0/bKuXhlRvKUMwzAOKvc
QVlkb8JjPSd0PSTDVeNCJecLKiXG0EYzclIkvO9J+5GYvDJUuSk18rvliVWS
EruYQjspIguZ4DMH6ZZbbEhmP2y4E/1WuxVwR6bQuDg8vzkG6xV6DWHbwcoE
XCBUChKYyXw4gqgI+u9eXahETZFbk9M2Y+7rYIwJCGkevZkL0GASFMlA+qq4
ecIwQNqh5y4fG9VRALyvbD1P+3Q2UOWwF8qpg+6xkHpNNgjO+t9GEy3QWfgx
KgBgbSlJ/WEqz9DRPuvq1gS7Wube3j0iBi2+E6FoFPItdwrUd11F7fgx8Reo
5oNG6jDO3ATbygRXmkr5pqVYdg44T+WJCTsc5vphKY9n9pFHikMNZG+t0brb
r+0Y+leFTwc90zQOaPvft58MnXvi2Q0CLSTlOwmD/DFzW0M2JqaXx6xUkWQe
HbpCH3uv7YlSOINfySFQC9pwV241G92tf8uGns/hjud7816TROizBYwLs44T
nEUg2NhQhDkN28JwuSYk1nLx/Z1lHSXFJix//w5opU0jf5nyn464FVeGQGlK
u9v5qF1AYurxbi0BhR9aNXkenSNNc3F1oQ7pUGBKDtuqZozLz2GQpNSkY//M
I1trWXDjzh9HZA3SFCbUGWU1tmkELwuwTMeboy/WMbKrvo4tRgdhGRWKlcPu
BYXI5hU31H/3Qwv1EWPZhCSqkI3z6uTEZdZzgAfrqdz5lOLvoBPNOSmi8QEw
5ZrRRfqz2G0X1Yi820+/TlAoEfmYSkywUd9izBt334CRd7qq6P4QGGWSIMkg
xcdgEp3Y222t8dYpTPgb0ij5Dndwf2PoQtb4esJmc02NcPwMhgdAD4ao4IsS
C/mxT84GZDhR9cVDM5yfb4UXf7XL5XaKwsPAa+5gqhMGjWr3euUMzSaWiNAr
zuTjKUlllZ9qz3NI5TE+2bSJB5Lq3/vU0RSrvqLk4tct0VRzQNCAa0tfEJmG
o9BHuc3w0/qcw2s7smD1tyTLrPlVv8OyRL3mkOmLll8SET87B70fFGn8/CuO
le9tEytaNashwMUg3BjH2CSPIKnXbOYr05Gc1VDp6/fpkiDNKB+GqazV9LJk
GoBISyO4j7KFwbYAumlbXs8GJXLjjR44Yq6BLrR+52aabyRQByRs8IvMj1WI
0Um6om1TSa7o61jybmbZeTMR36mi5cBAKylfQSM6TZEsGKkS+imtKxWoi6uj
kxV6ChpozqWvzJy5uVaxLPlNFI1dDfoGZC9jv2yTY6xailK1E8OLoLO5kJvg
KZZyrhVt3Z+zOlXATpAUILnlQbGCZPNtn/whMsdBnxpuRYRxRXmDAAPAXm8/
tc3lbTf9AIH22blBpBjKzTGTo7mtT2hJqKCar1zTFvTRBLTmhi+d0ng2pDYa
qp1JaTJFGyZD8lAcE/7G11L+c5xqJQSbDcdlaK3VpLWUZBhdLQBh2KApzcPn
VtxMmqprU3TVfk/SxHvjTWO4xQBeborkLH8dy4VreUKoJVhVkfEba1Vl2NY5
Dxb/b03mKbPr6lHkClMxabybhqgGP4dUniaMqjSfwtcEsMBISqD99L7xAbgl
DUjVEnmMEDsHYi6sbPU56/NDh8IFeZxPFgGhY/lilTjuBuetVM7pA6a6uv5k
f/VtWDBkNWqr5CZKEp0zjBSZ4Y8IJxiWN7jf0uH4OWT93RVgEMa0kUw6aTvN
fK+0Xa8tv0eDJWUZmTPK4yABkeHvGE/rMOI3OWJzolb9Lwlq6tcYPTikhAzE
lcXhY8mVFhk8SPsI4PBSy1j5Fs6eZxff7/eV5WHiBm6BEXbE++i+uiaks/X/
wEkYEcFxx65SktIwKir9blwMyBiu27rJXLfUT8K+oHL32pJsbgugJPB82pe/
CyEo7wCX1R1d1mclozWO4sC0YatNw2RGztnOFO9P3kLap8maiqbNO2Q5Wnr2
x31mXpeomxHmJ9HazJXHmJlTVj1E1zcc+7BWYz5C2PDypBL8Bqdvrke+Uie9
+HdYXdjo5CiA/PPREHd3JL5S75ui2l9MHB3ny4faLrL7UfXdVpKJJGyR/8O3
/vBmLfQgFIAPi7hhFNKI2VOcGFZJO1vB2UK04ikHJ4fBzlwTSPISd8zVTUUL
u3W4kaWTrZhPb0jxnAUvOj6N2xHf4NhF3h9mu3QrOH8Ww2QB6CUUk+AcxkXH
TqaWKNic57jeFHoRGLNLJ7nJ47wAQIhLb8V95XTvSJ3csG7HV9ecBRppsZPG
u51CxHInFGZ/pvLuGCzJiXxRM0G2kpbbRiG/2hKrrR3dAaNcqUbxvgxEhQg5
6WyW9kXJK69PO00TLVIPaXFRwYHV8erbI6GoOalMJcuPJNn4iMki7J2TsTXj
7zLGnFUMxl+KAh9PqvGOZ6lldSLQS2V+no7lhvWkn0G34c1SVgjndKVlzsHH
hoeC5ZKRR5fFBBo+U5Ih4jLx0F9mdTh35Sv4+L5g9rihK0QE4OtaHXy0ctYM
R/Zm+fn1g1aqzLwoGBOz0dvMxM4k7GD184T6TJju0y5TL1ui8+xK0EioInRJ
S8Y/Hf0iWvccds7JXm33V3/BHdItk1vqQjA3N5Ad6vlUkeHoqvJ9LSCn3RNn
X4JT6uZIn4j192QQfyXdZW8s32ZPTg9GQ9zB4hehA0hV85bVWevdK/5sF+LO
FfiYswfthyw3BDEz3LvInWRDWLvZZ5Flw8FoU/3gMJsf8LsetH1duwaLBtsW
oMu8pZan0txUH6Eqxuf2/Z5lbBXEH5KQxITZxZTljTvylPMONQxLuibikaWi
/YV7n8myz6wiv6uVIDcqcSh7A7BBX3Fwl4hDCmrLLgSP/mvJ4SviaXlRLJAu
YPHDJuQvK/5we0FdvPAVA/rK1K9FT2T50pd+FDyhdIQR3MUbF+MeAp6YBTy0
nEOJgZka1dBim6V6EhyDf959W2m707QltiIk1ZYKSBb7aX3cCim6rIOMGcnd
J0Cx9Dhz4MWwWBP4M5F9oHSrxZDwzuEgVGkZBnmbYpxIMWI/g+dIN5UA6nOk
AYciCpq4eKoArw8o9tPEMZnp9KZuXx2jJg3DeT7EKjeoXmzu6XIFtZRZsel6
G+7KQZNrwd8QzZjl3UV/WLzt2X0HTM1a7g3YtTyjZdnIaMPy0p7gyVbMxiPS
uTQCpuFnO8IkMfBVX3gpKWJNuWXSnkyK6/f5mBlH1mXnwe8MAA2grzyYej9E
cz6Gw54hEIJnO8X+1s7YSUdsAomlE6CehH+ZxKiCeHrqjIkPGKpYstMQUJvl
Ue4g/JpXiwntieYIKWpROkbtPwrd+UhAePOzpRPVhPo2Tkmpl1HF87xR0fGm
K+CUuue0Qm5wOAiUOwDAZFlUy0XyNaqoSRoIoHOpBmqm74rWb+4jknwv1CNA
/ASjedcoesaZu5OgFl0od792Wpr+7tdtLJvgQhC0PSIx77J7uMy3Q3Okdy13
bL8OrlN4Iv0hm6zNc5m+MJ9uo3QiD6KrIkn6wb8XWXoRwZgZvoYh7bkT+nz6
D1O4lRmeI6MbwCVedZT2LFejELtFtQ92qXoQshvFmNHeHOA1x1XFa4AdHN6U
EQaLsaKj7uOWRgHb5vhAlZ38fNQnlbRdh4AxoVJ9bYDGxcGB7Q9SwQqhsoJh
yHYBLG7Iar/N3xlaPjoQjxBTqtWob8Y0R/RI9zt5z4EA3XRFcHd9kLse2OB3
LHQChUJxw87iQqDKOeORFlhl9QTmAkiAA6JzheIykBy6UsGbE8UMr9pZUiaq
0xCnM96FUOR0BRfWFo6GD61NDXRLQSjT2S9NEySsfF7Y6nEWisU87WbKTX6b
1gLSpninVNY58Ai5hAUFv/isjgrRr4b2UBDpA9onNUz26KAL2vj4ArQXpNFA
gXVZfayVnqkf1U7ESx9r8cTd1Jw5lzOCNjr3GGdR56hcQLdZfRDFM+ihxa3u
0sVLEVSmnp7yS8TIseTmn9as37AOHYHVE32DYjNDkhhqhrV4+q6iFhb+VuIo
6UfNSpGvq6hIS0+1W7MKKK6deB9pzq1JuKe/4IkY+pyPHmRV9Y4bnSTkUY9k
pVDfYuYFcMZOBC+IpACJBZmEz4hxT8A1EgQVk+NcH5D/UUyI/K4H9lcifgk1
BuSKALln+xCJi42GqkX1/aoIJzxnf654fcB7MgA9YtyXA4BC3KOdCoKGzVkB
hxPTzfpxPqDm1T+pY+F1sR9+rXVwoUV0O3fpW1UcOQ4DckPyjInCCS3adasv
T/vTWT4fIAkf2pbj0Wu8a4iuvuQvFIgwvR/k6WuQPzoWM6fmActjforGfSTu
WGvkTOY3pWGi5AfUerULbJxmmsPeIqGbQS8270OvSZgk7LH7ER103ouq9j9L
Sijf/jaBCiZWlbYrIqJ/gzJ9tlhvLNnEw+bQPPhITOfDtY0HNdULbb02TGdw
TdpFvHuCWBiQY4X1YQm7VZWkMVJ9V0x3BZO1XI1KipipJQm1ygp3jnE3Ivsy
ZWykuG2f/WxxH122/UGNkeommXlSMERFuB1DQzvlVwHd5GBN7ArlXO0gl9PY
+1ugGvX1ubLP5pR1rd+JFIkATQxM3sxoAOcuJHSj0EpC0eDK78qtlhlUn6w3
A3krscZADwD86DEBhko4dNA19yoDp0sX3VqLEYc+/tKi1pZJrOKjWEGpx1PN
pi9UirV62bApyVnRaiiJ1a5SpaoIZh6OO3wQcRXJ4EdemSBtJr4j34vMyABr
aWcpEzOQuJZhyv7i0jKv0eSdqaBkczEaCYFuH5ltmhJW85zr6bRTU8hAM9Js
beAOJlmez/BLTOu8siWCunALBXGO2a7pRCTyGdbXVMMT7VX8m34Rg2jUsHTo
+TEe/VZaERBPh9zwhxLi+YzrAfM5veGd46DxQxp7B7aywevpyd1op1jAjPAd
r6eYfrQUCrXjVI986+a+WX+2vBoFgLzfdX4hT1b6uUTX0HGbsGnB/xiZvnVO
Ker/XQR3kJcywNy4UrMuOz0ohY5ytzlJVkUHNcFbpyOgmjzYJC3UoUlVJH6r
iPFmOmDiELUqH5JqTTi04+NQakVcg6AQBCXsgZP23e6gQlLXT2jwTRrpmQTv
QsnM7tioD/VqK2lvFvVBAHA2E6hstq0ZJEax/d8UAQOsDA96uV8/eNkVXvch
44AZV4fYDNdhgPajj6dqOR0EbQuozZEq0rARF8jlmQXgFQ2iUTUASJZZIluC
ZORZGHzBFFcrxYRAiaOs5DcNAlB9z+Tva0JtlsmRQDtlIR+sgAQNXUQ6vFPn
qg+jhILT/N6vWbCnfAFgS1xJQ7VdETwEdmYDNV/WKHUjrKLpCOjr4Fm2BxPo
kRxHgT9IwDuALQ7aVM91PWjT/Xz83NPeyxcVbD0UHS+rR0jyomsad0Lz762t
sLiMF+luLDLwQTVBf2zCG8d1ejQxHVYYmI+9glXmhTqkQ3or1X8B+kQ0wGdn
HQbD0ftZYjPY/JQCUT/22ZunCyHitKtp12R1WjKVW1sopI+yqYChtHbORb1b
OAnIaNxlVfZDJ1d422uUsjDyy2GlnP8HgHl2NLtY1SWUX94XaQnbiL7TYkW8
MQBg7X1L2HtW22WsrWKNeIPoylNYokaUr+Q086eYI9x/p6Le1p8vhswJT1I0
hwYpOKjt6D1NrZv158pNMZaikkrMY3FPQZK6WR3xzL9Z9NNy6RB4/BZgLLQ3
f0RTmCBpH1M0Kh+2MtzHyvi/TKOKONaaO80U7KKxB9URbNTvllReRdGVSaSd
3pCdvX2HeCrJYrOBt1N6m7xGZ7jFv0GPVDUy7aV56qMlgcZwokOSIvdVNmNO
2iRzYxJT30TIJmdv0bPtcwehwc/Ebm/75yNF1d1DzSepKgxC/u2iFWblix0Y
8WUnyyrpi64DYOhoG8zbvE6czn6PoDkokjFjzMW2TifJfGs47kkuzEkCJS9M
SR7CMrHfZQ9SXHnu436XxwfOQsrTfABGkWiwqmryaiSl5p/1Gi1jIysGIBjv
lp3rrJ7VP0781Q7NpPMR1iaqAvbStkVouoAOFNOlftibGwiiF5fN6TU+96h2
rB8Qv73sJUajk1GDE5kuw3az/ScNA2uDhRH/B4y18j0iGQFX6BoOEkjzE7PY
pmTmL/XLjN8vNdp+Z5AGmEJvvz+5tsKXvfnsba9IKzVKmNUHiIMaPRGPongh
XsKBhJx95rXFDWEC/jaXZPiHWcUnNGPcBoohvyK2VkBNRMoRmezf3vZNBUao
1DPwHgiNK9+FLQJsiIHLudXVu7Qg22Toi76yK82+DiKBvPfJ7/cbcg4s+9H1
/4+btdDBbWhPr/rjmDutQDjQhTWySI9jb/lz4K+D8+k9044kCYrLnL+RqMf8
Z73mzENbcB+sK11MWaPDiu91Q3WYK7CAC8Ood3KuPXReJ4pKC26RiuRwwZAE
tcl0AMnDoeGzYd1jqJ1/DRi7RR2fS/tci0LWHUMr9Jigc9xaeMNSd1hSefMZ
CeHlta+oUHp+R/5GVSuclVMX0cN5/gx2bfO+P0ZFuT30aPqW+WP8ZDnTuJMg
JveI/sA8bfHIN9Y4szlFL5JTnBwN2cBwnsl8CTlD1WESCWX036m7DtVTsBbS
bgAIE/tjoS089AapGKYQMRPhoBJxE0lxQW8hQ1Kj6J0jCjQDxGic/TOJP/mM
sy/jZcbtlvaL87DZmmH8Yliqnli8gceousAk5cLswFM+OktXE/Wc16v9Bz5B
MRYjaoo8K2a4vbZCkY6ovQb0jUsZeuQBRvxktwZkRrfQgtPHAMINxCEPlia9
BNViAFyvpqSEPnuB9/DnHijZACVK78hR2MKq3EPmngIDaetOc96A4J0jdac6
uguOkpklV+kkyEIw9zWe0fEY1CziV54PNESvLtdFpXCRYgDKqyrcsxAq/4jX
8Tmv7PdUmibIpO7bjl5hURTraGua2AwS3ZbIfw70Bo37cG+Xz3et97094ncy
W3+CED+o9wDAQwEX9Zwe8xMueTjP/fi3lhGN1/ttilFlYyKo7dipcRksQf49
cnFsLXLbV3d7W1nNuBO3S/D2QZQ4MfmgZkAB3BOsNYqdwREgu63pql0MQEIm
gihmlYedC+tSbCBEa/EOHvuyFtKKoQX/3u9ELtjEQtr/+NicA+8Wp04lD4td
H0ycDInX7hs4PCkJgzGLplX7CCF0vxXnvutzn5Xm2HE/rHaefhaqjK+gvp+8
xWJbkRxEpl9ZaleF1g5tMFhoAuzneQNAZYfvNITT2iH5HwLrnM3TY3KAv0MY
E+/qF630kHzVzkk75DlvsBYHfZ/rNK7jX3e7fsBL+dYv6ITHBLEVn6qZtv5Q
hAmcVTcav+8voLyEeG3z1r60tRK7uFtZnSjWjMi0Jre4xKPKNCZfzi5zNlVs
MIbQZlKzTlYayjdErmNmS8Wb5f+oXu4pRlv+f/NJSvmdAvD6ivzUC2bkAmK3
oGNGGXYcxxkw3OfmRdrZiPvyy2NHFgOvcyNDdJCmuzMnyUiUys3oARittV1v
amzqE2Wbqk6MTMNN38vcaxjJ6r+fT2V5tmI3GI6knNhueixrLFYPstY4LnhS
jYE1wldmNePFBkKig21tk89cfk7iChJp3k4Lm+QyO9guJK5pm7FOuGpf9SUU
yyxG8BVuFNevz7vIapBNQqiNaubXQZWPojh1V6Ao8QW0ZhO6wc+pw70Wdtps
cjBrs8sxKqC0D6tXMTgw7pvSZ6MUhhwk+0u+e6Y8SGa+TouecnZmVkJ2E3M4
itC/XaVKebO1oJRpfp5oagePQCka9QswD4vM+c2/bKrO1r2q2GehEFjcX4g1
dB3dxNDK0IAn2zFSZCmlrgg5p0n0DxO0FmI4lU3u+JBtUcOy7n2zbQXNzNBl
5Ke3btyYnXGtcCArXZpLzAFTkFbbzB4qMAuWjlyECteYWUG8KM+O+mM3t8X2
1VxoK7IR18jIcEY9iwtOELF26BjJoWezJzXpVaY9Ocls16fNol6pOfkVjD3f
sNOQ3p2lxcQ1fe2wauZD0iQGo4yUVlFuFnoxqP4Jt3fnPyO/h0uJ7IAAwONk
WmA+7VfENHbd09/EGhDjG6RQImnvleg0eSB+Y0DmhSG8AcMm7UXwfeiy/T5y
64Mi89oU86R+6M3IpgYTSc4q8WO8CD65qevy59Rc2wUc3M81qXXHGZAfZ5iX
zsi8JVoMXhv6+7s53RUQ1i076K8+a+IOBT3ONd9Ue3Wk1m8pQ6XHxN2UBHr1
HetS3t2RUi70iHLC6SYrJt0t50QajikTGiN+jd6pKOHMSzD4uRKidwz5oNNA
rSgr5JCq7he8fKGNiUtTaziMFFL93YUsGCkTeA/UVulQeuyabLLrVZDjWaBL
gGk/NDz0rvCfdoFT54Iz7idZt6l0+WiIYJMGkjpxCuLS3mrpdKZ24Ek85fvt
HkljMBtIL2ZKkfhxdeJMtRbkHWJi5lv9cR9VeSzy3Sv5igcwoDGnCwt8qw3y
CFvi9hRAEC9Xrbq2lf0vJ11M82QaNeWjaqdaolMmwnn6FyuRqMjMiT4x9hQe
gQyskQCs9OfLIatvMJuYohhRtAkZwVLsUm9VkSo04kOl4TzfzcZG3nIipx/t
BiJZ25QRaUynC3/wk2s5VHaPObUaOOMqxgHQS314x4fflt4vIwezgAuK1t77
o5HfhKqv/63UYIzVgULF7GdG+xFSlBc5iLGi3T9gzxeQ4pXRycYpdTSpDYkZ
V15QkPmTZCngrujYzQA+35w1+wmfxijcVUaNB2swaZsfnHECMiBnLkaohiQk
7WIKZ+wPtnDGbo0ZOtD5Ng9G+6O01ww9U67f4W6/J6s5Zu2Xwr0k9VWFfTZm
uGX4tOml6/vkxhhXNX5zpDly5Bv3bR/D2IBONs9BLloxvkSDpzv42URrbYHL
ZBRfUqes/p8CgK1BiZzGdZyMaedSES4cuWiWOiA6w2E4JIstKRnEhnt97DkY
HZOQfxsOAZd0PsZyjLv1LYegBcLF4uL9JKGC2zuRBr9A6i9setOboe9NKaAP
mLXSqNYwVwvQSjenpZK3uJaMsh9tmjKpx02KyLsF681+51YIA+8BCRrw71kn
CUunOpMavR2DVJse5iMzvSGkmQqv36SQQ/8OY/kwgLEye03Ca04cUiAFKlOX
kmZkULh6mFQqTRrvoFBy/Er8WtHaaRlk22x2f9wBiUT1fLqzbiOvQNiEQ2iB
ineMEUzmvegaUJglXJBPYLMSJ0ohyXd6yvFdU/Jbggsr8mexAo7ExRPQ5Np+
gJj1ABx1KWTsk+8sv1BE3vtV3ViAVg9nrea41Y4BnCRIgFW5h7Pp8+VIuvbH
hpQr1J5p1JcuUbrlEkdHw1h8QGOFGaVfc3Xp/2v66wSe70yClZ8GxX5iWd83
1xkoGNdCyRidkhQL+pgkNYBrmcBPcA/hpgjXFdaFIPiAV8gE8Npl8mQnzAaU
G2NaJehqp+yJb8cKphKoW8WbzVSIBP/E3CJCffqfVb2P9DyNUMjQsoGSdzm7
PRc8S0HYZopcLBA2JkQKGzi6ugOqsahNCZ/IinhjiPUnjrXRM3q58VSHJzZh
31ud5UyNfmeYP4GckWNar3fWRFtzzdXt5uLJjCevZH1i7xELClK2UCmEwHDN
2ujdqS1rVA1eE90HOc+0fQREEUXvfm618tFjuBL2pB++TS8XwEzrSiX+qlea
ulVsQhJ7rp0cYM0p49N2nClwx+E5xbsE2RsaIfBQDiID6SnbefMCsZoEsnjP
I+JUMW4rxXqKFU6+yCLBS0hzQs6gEVVykG/PO0K63FJ7+BKQKCasEiWUJEII
puTAMd2uSKa+1R4YY20cZahAulBr62O9VLK5xDxwY6r8wCrzJd5Isz1N/Ghv
ycqmW113d3BRW7fkjJSrg7/hqSUIexP/CHnmWaukTSjostAT6x1ajHbf23Ua
kUnI9YGcc4vz6fXvhdSd665GujFFA+y7/tIhBE2liQwbBN3n/UhxWmBUuh7m
vU9KTmNWYEeDeXeAVuUsO1JmBbOdhtS/by/zL/AFR0ir6gBKm6gQrGeOEPbC
2lo2uRIeyzcdFnGb0xhM2Z7LAzGagiIbjFq5tZvdRjwl5E63bruRRRTH9Z91
2D2JPji09mVi3hrItsPLLZdtsD/07vumur2ozc+MINEmGYr20UfTSaOOit5m
2B5bYRYDWfnjGFx6vVeDq7RWs7zzQEqOAeyLQdcwEzIdvTSl0/Fu22fsXhCZ
PPiFHs0+IFsnjqfMg8MDesfPKFXd86dSc/Xgp9noI/WezF7z34seMouWXmf6
HCJ63RZ24E4KCW9IqZhzmpKqCuaWPVdmENQWTcmK3NCxFE8FA8lMaHKcuhyh
vHdZbS5aaaJvkBPkSLn2ehmmeX24xEqpcIw7LcY0l7ydmeS5d/Vt6rI/NVpG
iMqA1LOj9xbro97/0WL5AETbXNWDDDK28n2wDejgDwXAWBgehBxRos/A/bj8
xt5GknUxpkUKdOM8hJlLTVXIq4HLLpcdIWT4m5Dxt9D84pyp9rohz8AzO3Kz
IjsHQDjT30PhvfH+cAibWnmdATVTcAvOmBFMZx70zkq/31UdpEVJOrEWcWum
UMQmTyqMP+DB9fljhuXBhmJW+xMc+xbqV5pEPfzgx/OeIdWtxhUcODsdQh03
NXhnIJJAymwK9lzYf7/xVaHDxP3QkgX0NcxeRF638JIXACQb2IOaf8wTomYl
joyaqLLFPaBfTSdGRGjmFnV7XwOIf8mlvHXQM4vTUxSP5muf9XNVwxC11bvL
RkcnZB3ISy9Y96r+6pzyqAWqQ0k2lEVUW268urgByNntXunExt/jUfJjCt7h
l6ct9cDf3ceezIBFY3gXD7TeV5Xh20Nfn7oR9TB6lwhuDmXlyCA6Q83vVOWu
10jULGJrkOXOuEXMAanYttpWO7QpZUigmqtgIVqfJEun9VMV4PLWFzWGrbv4
zeBVBz9j1d/GlqXebjmAbOOXOZxeI+8N98CNuG5h6pGaFvean1vl9z7wgltu
ZW/ZB1qODqpjuziR8frNd/vF90GMb3R8fWAx4ib6KK+7rxUEUfFebq4qFnnT
e9Tmrf6fO7bqS4OGXHFrSt09uVfzu8ckBc1Fk97PKQR+OtmZm8pBzb805dY3
f2Xn9wsgGsE+YuLl+90hzKhD4xgAojW1+KlsGEGQS2Upnb1q6HqO51HUaMjj
IXbcI01jGylPp4h0DKOaHRLvHe4E6JnDIoMz87zeblfvdQYw7P1d0ydayJIu
cbxm5xQWd4aHoqVezQaXuilzh6OQwjl9+FJwl8It0c0qSK6QKTGd9kc7gICt
iB1boRvxkRNKHeqGV7LY3Oi4sJ5GMVIa/t0AbPrgxci16YTmV8CTotE9bxyS
A+zPRvJ3WHn9t/PR6nHQntyYPMEq98cGf0pwttBrkZIjlGxf/EZ3NYEVZUUD
pSV1GFBzT3USA6J2gG2kY1T3N3rAYs2nQRHscWKH2GuAoNQ0/wGmzgNsqQUq
4wU404OeotjLcJDFr3OTi41JRbxs+yHZgfVl+6zd46xYlxNDpnoAX3/ua494
aFi1waoVJviH1c0BepPuS+6mzYx2WoggcPy0snFGBCLmCddnBxqo7sMpE4sf
G736Jpj7maFk2YqOhTMBdwBhQSRhDX3ZyYGjXjL/4J8iPe1ij2LortFv9CwO
/prJwujEnGoyLcv1UF1V9e5iFsqKmJjfiMBJTRuqEDFOdMbByc+to2ZYNE4T
GwjAup/hBsZyAGq+nWPRONSZ3pmvHkpQiFQZwSIZOOX0hr3bWGeLbBFKgMUB
4WVTRUuwO0CpNJ12D3yRKjMNeXpePhoHjuU++6Di+216XOT3X1u5+qkZdZT7
sb9tCPppmyrL6j8A+3evI/25qITVVgbZJjyuoz82dP5eY6PH+Yu5O3QPBA/2
0QO3LEOncRxbbsSRkGaXdPkAnyldYKaAprUNUmLM+nXe5sungudDSHMO553X
AGiRhok7RCjYtpO0XqDGXiVDcp04dnhN2ePsNH9g78yyCG+W7mZRdKl+BuXU
44dkK5hnguUv2//fgTV5GwyIttzZSziy/NbD3GvLORgDOy9eZ/CaKNKbFZPL
RJqKCEBG47QsI9hkj0kDkdDPoAwo1h/+5+98WhOf0OCH47XzPDUph/KxLo9r
V412FR3PSCZFVwNdUJcu7x+IBNfvitxWYLCCQ3fNYBBKrFAfOObQwQ0Ajcv/
tqKGKAY+C92hZJOVAA8Xfd6YnJF6r73Lq0Cs4bOSjwrJj1canP7lCnKg/vnf
8OA3dJuTehZU8SFqSV0UPRDFJzz/NZkLXjjEQwAalxcsI8NEEFs4/3qOF0pl
roKdOFD+X4wrXRoSlVn2domiwRTKA/UVGjh0LlcOaKdGW+sOX2z8O2S9hdxg
pF+3CBqjIJ5A3XppDKPdBcOs7BqmgGOtbfhjaZXYbUIhZ3Br5Y503QoGQZ01
oWpOaijwioHdy1xklvkYl4/gnocGr9jZY75s5mEAgS+8ufLiV7yFtgsFY1Nk
mGtEy0Bn4onf77RBsAiM31OVL9+4p6Gz+f1G7f159RKYZeGZum077HlhgtoK
zCd9y7ai1lbFBtRfU9hKFdQxirsHaPmpTMdHj1L8/nfqFdLZ/c5rW2yvbEOo
ASmWHIRNu00V8Qqbo8uQm8J9EYvhKZumLhJ0/Y4MFTyGu21HhxmUQZK/QoF1
ExyIDjQ1NWGucIHdn0Bes5lJUHPq23REaAj+SSbofgvNOaRAJp2XjbxPw+RS
GImchRhhqZLaLMnFzMWMRDA9D2iPySg32HpruXf0i5IFdIrHcab/n53x/vgo
xB996LjRMwCH5zO9I6KEeaWouH09Lu/14clVHlS+qaMKaw7GH9oQPjPfRtu3
K3Rfpn9S4szsjsgUN0jv6bxkuQrX9yGrCOywDf7Vk2heDhlvXvAkopVlq8X9
+8tL4KyqpCk6cRRz8BDpL00zRCFTk6miL4S+/JeO2HvITM7+p0yTwseA0e+8
v8FFP5gouKPCamVI2R57p6fSEt0hET3vlkJGRFAXw6ghFxltA6s6k4Y+fTT3
PfbHaTVRX4T6vTDHVhY4zReeFtow074VEGqcEOM6gZL32KSWiT6fW4/uWvN0
Pr68hqrrGYbYsjTXG8+MUUeU9DdSF7yUHxwTzhArs5aHGH7KHQ2JwGpglHhe
EGZqwU/C9xq50tvkFhLWu2oU5PKQw7RAAFJtIqTOLNdsuBBILSHM5cw4wLJC
tjVxfh3MYZW4nrj5CyYZySWJtjD+E+QXxN5QLVwOA5iNCoAqcG5KicqNwtG7
nttEDGdk9+L3m1CC3MmJtoThqO9b94K13EAEqeL4exXNmGVnl2hqUq25jUhc
b7FNIZyZlSYqDtCgfeYpRH+MHMQOfW5WB3BgbPWY5hXnJQf73OEA1pBg0bnK
Oii4ls6O9y2AI6MJRdM6H0OkkdtJB0Px8qUHzQdk0laPH/1zaltspkx5wY8q
5dRUNL+I3+fr/pK00tOPD0CgUV4NMP1YXIydCjIYSNvM0nWGKi0wjv4wXc/A
yW5yjbEYyno+LOTFim2R6djcdQ3+H9xaZA30rG6/KzabhHOabyKQYEGqkAFD
tQMOPNTCiDhLxmIyYH7X4GRzH/SfnyS2ncLjLkgDfDgMp2Qg4W3Eq2exArR2
tvXcbcn9EhiGwniuPjGmSQB6he7NBUxMmfdBPmUmGvp3RvZg3rFAhMtupzH7
CPOtE9IJrr6rOxX3sJQuwYFfDOSfouH7hGTvqupGMM72BI0g/6n2yZN2jtFb
/iWuHi9ZgZbAMfpxPwkRdG1McnomJX6bmn/EN5dgukMdfQ46qfV1EOhW/Hph
j3Fxsv0TV/RHxWXjXDQjze+NmQWkkES9tD4h1xZ9fyjxWxIUfALNSrW31Esu
3R9FBoZZ1mSQXGCB/NNAQjYKx11/MCjI4pKEOxRJOtFhEZW19s9YqaOTVcNV
NOG/CJPB8vAc96cCilc4XscUArJlvzKTIfEkvvyMBI7M/qMCb6ac97rkWg3p
na7+hzhLg1Bma2RNafwAkyKGH3MoZ4EXe8gi1t/se7Rc2BnvUIcjzTEGJ5VM
TEG3tthmxXQcWIJUEu/dwAcUa3i+NdDbCnLq65ygGZQSZj/yKVL4ysqTSI9s
fDwnC25ustJbmTjjfkQIGi/hf/vxyPGUkysje+kEaA27UIh5RBGf6exjMtSv
RcmNlJQm7/4MutdMJpPMssoHEWq7Zt9Ho+gIW6weha/6vrgpgyMG7UlK08XQ
H8mRscvI2A8L3feduS7rk+FrafOWuCbnd8U1l9ktGTvIi1Y45rAeSg4ahxQt
YYgkCAOqcWhyXChY2kz0eo339CyD4sFneOig9jKpJaHurd4zHlGKC9rc+3k1
FI1KGBNtm4mOfdGjf/KXk2M7GjgS/hJRyi+wAWJt8/P1YA/LMoTLiQrqIGq0
Ku2TCpbocFPvACKJdIXnIfXKuABE7P4mExM6294/tRd8c2KJ8UE0vcaw/p8n
l0+NqasYxURTh8834XLQRkbuHs1FQpJLArQWFtUmdpWvAWYSSHklmLCHfVnr
aN1Yso1bpQLGyFYrhH0BhAHZunWVswLdqGs+aj7uf3Ifl4ZfpX2Zc2muOMnF
710nqiTo6kFyL3F007pfPng5BxyTxpZnRuSvB6t5pqk8NJs4pjn2Equ82I+j
4L8L+PQ4G2Otja44L7pKcTUBYdWXAp5SAeU7yEmxGejNPKjHiwneMCSNuuy4
6XhyV7qgbB+8cMHjvR/0GF8x2g2FwM7F2ZreRoA4OQzGu3dUUKiCr5vsvXvy
m5YcgtTXEXC+kCVHEdq9UDmgbijjL+Gcvvum0weTLpzddmsMydmgcJQCvhaV
orkUQd3s1ne7eQZxhNRGjXtlWyPUrhrleWVM0q9veUB0Mt1LlD/zwwWSS5Kj
VUZxx6akr8Dj9rLq6WGecsVR5vLm+fWwiMHVZ/fg/wnOUa3L7khvAhllbW6+
gbF5HmwA7+AUB1aZIP54jToBtl98m7zAwDyX+T95mK2BdZalxmPK2c7haD+R
7VRBx90/AjPbg21miS5gaHWL16T0NYOQaYtQTGgLK/HT4YkEnBgWOdh19C+T
t2tJn3K4cUJdRjzbSXBM8ma30fgCZ3S/QQGZheLKzliCyGalok5xXy3YOUTA
pR336En2351LKrjK3E4u27KvWisv6A9QgTVz3CJ7zDtf+c8utTbJr1LOSGt3
kRmkg5R+6OUT6otBe88VdZm/efuyiz/DdMKF9Ucdtnx/4EGmRDBnSTSVwh+E
vUO7Hz2TcyZ7+VviyNoBxi0Yy/26mF5n/4VC9YzHWkAZNHV2rmKYwFzUXoUO
E0TVXZSGfRRkTxUukPOLwEcdb8LIUvEvnWY24S4Utq+FG6AQU2pem8sQRG2r
iZJvs2Jna6PvI63v1pQZb0KwGiloRK4x7FoZf/Plu/Ln+o7zWBalyqApv+Ak
RGqT6uHONUd6bRpctRPkFdgXYjlntyzjcVz7izh8N9tfjouj7xKa7R6mC6EY
ZVb4jSJzEtbpcZFufy0iPcvKWtEgL/zHDQclNc1wkfSl/RLHe1OPs5qw0jCJ
KLDf66/P0zuieGfnm8Dj/10Q039rOlqkGqw8DMfEjR6U6RWr1SfpgID7+/ZI
hCD8/Tv30SFIdG6PdRvVwhmrj8tVohpPKnLA0pXEwwvYlJGCarrHbCfZ9766
YPTs9REvbcKwjnUewlOAUwnoFF8d8RjnVjIydHaKiBzBsvuwsLUOEliLjOhT
gqD/rZI8RYdPm2Ecli8Cn6v1A2eGByI2Fnq0BkFfVF0Z31ufOQv5vzpJUD/F
bdqwMZelzQ5lpchi9aF9f/BjNa417SM35RLH8Uk92rp25tMNXkVebx0l8Ag+
lWNNCQ/T5RZVcjbXmbdy2NMPZipHoIKXXRZaNiq7KKUF5+cOt6k9uRHreVnF
kNEHcTOvfYl0U33K4Z4cOumwYtPPqsF0e5UsCGMWWrwo7T23qG5gF9YbbwmA
ua1weYDN/pnmTHZ9rIGv3eZftwfEJxsrIgeuSyqyUex1TYVua1K5rzOVlygJ
recunjk/koiXSdGUR2U58kGjww9xHmsJ/kw9n5FK0tl4+NGx8Fy65n6Zg9l8
RonMEBCKqPWHKvrgMaPjFhpWnoDre/Uo9nYMtQTfS8iTZM4pvDZIsnhCKgV0
oOv3Z4ZZQxtaGaaYYA8h7XQMcrxURSev/De/ldDp+BMhO3uQ/on4SjZoKVKY
A7+XB42LvANAKqSokU/lTBquDjTQeS1lm4C9paWyYiBwDrkac5EBmKjAqlKI
g0lwl3ua5SFKTkXT5Y3i+SfuEQ1LFEY1sqyoSCDytyjWZ9B1qNths9iloo4h
CPMhtlVkjGamXpzItp7xTK7S+oecEoWIMcmJVmzPQ03p0rALPuCn45Nqr45k
ffoGcqcC74g99eplvtymp4/XiYnN+NppWVqxSF4bx+J2sX9jpVUa5k/oZFvI
B3wi5WnLY9Lr67841dfwaJ6ZPDyYZpRsuW+rCWOBfyJNIF2A3AWDmYsHUW+L
EPp7F2I6spugfzmBXzTCMFDrknz5cgxyTYHU/qr8OK+CKaIZW7lPLGA56Giq
kpRmw3G6GdE4V49A927DtSC87HGe2HmiayJwPTAMA0YI5XTsGVaTwY3EvOLE
GjS/zwcitYqTy4jYg2yIUshlKwQsiZS1cl9yn1ktGP13sf2nFPUEymI/grNf
ZEYmP2yfI3eU/qeepK8F3K5IuEsG9YUFA6pjcX5FVNe5HFzwWQP0M2Cajc4G
SOfCjj7aJCOGu1pwZrjPbjPkRqPAGzWtGKhap2X56bNT57lHEAFGhH5BrXlE
1CZN9Z/xfHVUtOmSripT0bYbi4pUGvyi6xd24dSmca6YYximmOYfLaXTzyQ8
LgdR72d166t3omEv0kF5Dn9gtCoDH3tC1OqfMxbrBRzA2T7LqhFHF/klZWKm
vqaqbeM/F4qD4d8lXcK5DHs3Qb7f4/V/wY/0210/0mRphWLp9f6Je0mMJiXX
nSoOexqE5EV/3zPI6qbPmx/froYtHala21w935kvRp+O52zvXzNhyInTU3Z+
RI3OQqhtr0fhDLnYBOmn7dHCqt1r9XITmrdtepxazMrDtu7HQeAJF0Y/FjKb
M8ifBGlIFPdmUnc53DxsovGSf5hFqeMia73PvXXTU6Zi4Mts4ZEjzDSbd2Uw
Qeo/yhkrtV/gj92OT2X8GHNpiY43RsvT6wrfb9oC+WaxdesaKTXNb70axK1c
/BU51M4s8q08OeCKJ0TD1HjhIZgXUtOXWKee65W/MvBMhWE8c2rkQMaw+lR9
d/fEg9HRoWuPUe0rizRdLc/B1wvXb0m6Mjyrjh/vu22Y+9NNjeL+zSqNW4Cw
MCMUuZJ+ANGW+c5NY4/XRoWFKqN7ZXe0ernjWvaL7JrLmGwkOihbp/5WAb1f
OHzK2A4y68wf9dBTFBwP2vcdgcpN0FZxQrU1H61byC4cUM//3v9rvTlNAmfY
3aueDs74BxCuOHjjs4WnF0PDND2t58IfO2fXYK88jpXNPCde4jGgc6d8qhAV
uj4tRLxlW4sYV5GbYofArBnzUbYC3y8Ihth3aR5qyRyL/1g5Mk1AVyjX1/FI
tMnol6fEuOuTL34JRRQIsExmiCu4ZlqFbBzDMXbkXtR5V79yjpb57HMlB7FM
PBeHXYrXmXg+hyubnBKrQILXrahJxH7okTaIGrJqtDy/pCpXfSSc0BTFEJEN
AU5mY6ZA8uhc1s99MdveJyJvA6ZWhpMgb9Bd3GMA2cDHBT5HTkT7vnjFo+xz
5fkKJbnn7gPr6t7NBgCYiwpttsPad0rmD1D0AFf3b94Pr9lDB9g2RyW2c+qD
YjHQxsmQlfCBNyuH54CYOSI88DYYIBvZebe3huYAm2LOoewyHH9keoK++Bp2
7Jvkji5Lr5cOgYjS8gX3Tm41JA+OV3FjrbzR5rpI3ZNXRZCenNt/DOFHTNYF
jr4vJQAqLTJgFjAJ7YfUt2B4VLjv8/NrxCKACy4n7VRcU/POhpMDx6lNS+mg
OE8+OpiulayEFx1GVnFhWPr//Jqv+sTlehtNrzNMS5wZ8JVfU89FB0uoJlKt
MJn9v2pY/QLcIVTgkLJHAmopxLa9E0ZyFmv/adHo41sToKLPwKGrYWMVfYDI
okCCyaDUvoyXcr1lhGxKKooooK6fb2ryug6P9EOTnOgGFrtz1/yRyLqhGwGO
V5SJVMdhzQt5eucdIXviu0VsfWSPY7XPFXKJWG18EQu1Zok0t7JgC9800vDe
STPcWe+A7RzsvZw1Nadn53mxtOGrrl3GScBt7NwXol7NSWB944/rGp0sQ3IL
iXW5SL17RxoV4LHOJJPXRa+yDW8laeNAx0cJ1AXOzfUMlUlsGnelXJ5f3jmW
fFO6DbeTUGmaVv1i0zLx/Bdl0z4RdZv8yfUU6PF9PVzcK+zwOMSi0t/DWVet
hu6xgN8JICBvs9SwcshX1fN465iQKGxPnD0X/4ib9Jf8bgtGATUzUUdTu0ja
rSkHBgMbzDUzKkK/zeR1EDoFrUoe8tdTvPOZiqoY44G2HdSommtgMEHfkZ0u
GOyca/WL1wXv6z3XQ3GSLpZgZMnp4xL3AtLA54Tc8qNEsa/9ry1+BLzElceq
i13OJxM8TUAZqYlvWPpAnoubMA9Cmi24+nAYeCojueun/YtTOj93b4j3xQ17
hHdOe6GOrMykCBNhgVCCYQyOLnWwqknf32pSmbcdwIryXG9OFxl2Sk3cPwEL
ZfsE/5j6cI6Ype7CJ1iHcFSA83jqhe2Ylu3J5F0h5EYwHKx1GbQbSyIA9db4
0a2vQIDN2OuboTEgn9VxGDBY86cyY3G9sOY9RuYao+7MMIqxUrF5PMkhKN4M
BwGOdbH0DMRoustgEG9evD/o5uSuHF5Hnf0JD1/N487+9LC6O2FkXq81qgbW
YvoQyc3klTdwmbyFZtPvWCSRJU6Ghk+UQEQLPocpt3neP5K58uAHdIIMe+qZ
gRzJwtdRwqiptCdmiq24tzW3RhXXQEKaM+l7SLZ147cNc1r1ZcVMJ7xpaN7n
SPSt6VL0mT8MOjCDqFf08p8MkP7RaHl2VqGo1OvADHand0DBAsRA9VNJYEDX
aYyLwMJ6mKlwo/QeheU0aspG1JjFCq6OY7/Ot8ED2/KPfwY1oXtwSnpqaGu+
x1o3kNRa8EDvssEe78NEelcTMaVhq+3+bIsjOlVRH1Y5dYcF+Dgpj1ED9Z4k
58S5tp42c1v9QYE1AXKLu7SEGPMHU/WGWwaZrU6BSD355YBOnL6QUjjZ+MSl
+lVf4QFCGKNDJ9k0iWlYkE2Qk5C/UwaSdkScLlpfCjKjijC4PqsWHnUGn0LZ
EcSOt1lb7vN2yY8vFDw6kXq7dTXO1309ULVnLpfc3pWu/NkNVFtB2lVYn/ay
27lBh6h6qYQfbvcJ7tbMRSkS3PWq1mHt/0oL8r4EJcSU/f/d1kevMRhd7ZJK
lV5TocYEMqkKPL2AmzOUHp6Z7U8Eq5Ol9JyHo21H6Bx5JRoU0FY3blW/xDD7
z3xcbEoXtUjwuU7aa6IHneMPjq1bZlD9WB3Bj1NKnmRQYd2QzYh/3M1v8102
bni9uJFwbjcunztqxqdTGJifnYqGRu7Y8IsE9YaGYlhVOuiaRoUEUBmILIl4
KhFPEi+HOOovM4qMQqESS/GPbExM+vahjPjvNbv7dYDaHEjCpP1zNQIdJUpw
gN/JLBrVlaA7mmOOsEeQatfg5xPVdQLFYW4xtaBDF/02P0OzsVSI5PGXB6KG
uxgAluxaxYFn94O5WEv82UyaAE/01XtvUpCatfqwemwrx4Z/bNKKos38ssNF
J0cg3IfO3wR0PdY7F1m7pSpCcDgXpwUe0CMknKxr63RNY1agw4BKi5Mi8w3V
9xJ7R2pK+gKeIDw9OszheTR+X29irMA1fL0TFVfibN5enPeYzedSpK0dPz/i
+hKfpvJyVb++HOHKXmnO8z04tGw6BHnSvKafehqf0LhPBVfSBdrch1ItpXi/
/vLHXYYdRKk1/zTO4vTYq+nwVtHBuGDc25iIbzm0Rzvg4El5Py4/6qwSCFoM
GTuNWB+g2yY2djw3KqdMPyKICMX8z6dEJVp8FX48BLcNXd1ftvZUxVgzUyVT
dBRmajiGRH4QOheGPtaq0ONQqup8VaYyAKTiJ7hOCf3PykvmjCDmNqszDUhV
i3CXjeWy1FpTLMkWUZ7hBOlSJ1d47MiPDsn+vEUOTS7jGYmJ4N37VxWxmkpC
qjtSv3iUpM94ZfHK04RmBOgOP2pDD7bz/HxYuqNGbFTm5Dd8jUKwRT8yjrwF
egcuy8pLwVV6/9xaNgM9GMhcob7UztXpeh+HWVnt8W5v0qZL78BC0dL+d4vp
S6sCACzwVYevllKHIONRlOmJv4IzGM0UdOnq1SJKY5ExGLwrMIy7tCG5jPGa
kcn6Sl/TuFQJ7I02CqBTTGVTj+H+4FAqXAIy+BNVsOBbJfjtpt6zAAtAdtcU
CGxXRM+ViuAgfFGqoXyrQxIJm1+VqFI8vJIe2BVIh+uLXvZK1DrCEekDRF5h
q8+O2nFqGL6499uvlPlqdVsHUP5wfZ0uGpDekXjbo7J9fqeIFjMwtpDYRaAX
cYA5o2EeT30Um52nBfBSXmM4nxpefsKL+vscu7UvJMDmPaone+RXmvAafhak
oGPu7EPNLBrJWcT6cY9s8GRlMLfrJHGNUqVza7uKEYdHCNco4NVn5Fu5rEJS
lyzdvJx01XUod8c8+2zdAB4xC7ZbSnmU2RjEjMAovHkhAFobhXbMpiiUjyWA
up0achJgmJfvQvgolQvY4HoqiYtFKi72dCj2PACkdGx4UpgIIceZ/RPx8+zV
BIWhTvnnzJ3Ft5dmmY+PqugXnrCQ/TmbVPzSc79kaR+SIALmRia+Eddzsklv
ojqNoGiYtC02Gzf3HFNDmMRTSLemoYEXiG48jzynoeT7LxT2t9Nv49zVC0Nl
+u6loG/xpa7RdMCTLnoLhweimBP7pvAfcZvW1jAIcsfuclMga4dVIBCJcKHv
OCjEFKemEQTuoZJgBjtvw8Mmcwp4qe+Crre2LGgsmC2cAUeUPdtDvi8s0Mjh
S3JrFSPalBQJazzodUx07SIhoEGjHfMJAJdxrrWmjaurTR9oRVowhJVoV8Rp
CgZyoGbabtV6bH0ReWgkk1IUqcjs0BzmDFZKiLTIUtwYeGQXVMmIMBpgbLhG
01ExtVtYz2N6hCMw9dDb4BRIbVEOXKO+JZWXZaCP8XOR6VpPDSs9+bh58H9C
FTTDilSN0P0UD0Vpn/PemEz6ZXs=

`pragma protect end_protected
