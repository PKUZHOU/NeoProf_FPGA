// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Xy/jOIo0BI380NgI4nnIC2WJ9FFzmxK5HYNXjr3FyBdk1GDwAjgLjCKiv+Nq
/IYANfwafB137MlbMQAh8nUUzXmKIfz6VvZDdlDD8r/8v5GakS78xE00HGgS
EpPEGLyRdv3NmLNR+H3ylUmY6McGXIR7WGsbeXZbpoZDKwPY+NiKyyI/tBB7
rC1NnBtftEc7wOhgF+6xe6XB7xZgaM2/scFTZ4SMSk7/FYgLZSZaqeMhLgny
V1oXROJZNqCRBB3eGap3HJIB7Irj5ns36ph5cCDxfUceU7ZcVx+NVWQT6B/K
bXpqXNZN35gVBw54D1y/X3FwwRy4HOTbcxILbeXxxQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
GsmfqOqT937F7JCQVWKbmwDqo+T/m4gBg/b+LIdcEQjkbwvD0AYouH76XyR6
QBsNu3GRIt06hvaU9XitSZm9uOt7sELzNnFQTiYG4S+1IY1USoAdwaaWg5jM
RaKEULNPgejhUhsfKfE3ftSlDd66HcHLxkQMxUt3KM+uQQiSrNPwSUIuhfCf
75DaHyoBO6AAp2feCM7pLFpnNyb928cexnQrg8I55BmZ+Rqcl+nDM03Xv+gt
eacaoznpv5f8l1yPcBn56J/zzWIOC/6UwQdyggO0fCAHoW/Ud0mOuybDCHIM
RUK32mEuUI+wrcJrNhYbIlBDFrV0PN41538Nw8X1gQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
XepD/wtbIsW7TlMaWes06syEAvSUt+tMbJF9SlCt5DuAxMobCne4bU2TxkNx
A0YIJdAKPsPh3OjgXEJTLsu33GfmTAYbV/wd/vR4oc1Rvs9EggGRY99DZE0n
0URn37kyrNKtmGuoCKrCaJ1T0SvgNPoSCAgrXnT0rfrtezIdnIXRVz5VWobU
btlAZ4Kc/tlvLfdJA2/ryjgd8xAaoTINik2CPl/CQNerwpiBp363ApyP5j6u
iLwb+MeWptSyzc3x37mWgiEG4z5XCF3GQbvcolTgN9RbSsyPQad6c4qBTjxi
FOi5NSrYSVgGtwJEd1ecI7AWlQA/6WqBPTc0V5SZNQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
U9TIqYgR/XeIuuL4IkAdd8llH4Q2pFoZo45jraVCW3tNkDokGt2ub2wTUEJ5
qyaVlkTI4PBpfevAAY3uouaLGOqfDYwQJLd6AR5V/gTtQNHnrR6jXqOz6NWq
Ht8FwKok0oyOQyRbGSoaaR3vzjIIMAYkOHBJ+HXqvD5ygfbAMUk=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
BEuF10W1iFYA+ChvicAfniMl7B3zILPnab14i8YCo4fEqPZJSoe8suW0cboq
3H3nCaJvjRoP3roaXh53NWKxGOrWQqgtNsVvvOX/8nZvJgYAP0NqwyTuaavN
P2R0826/QR2ydMowjTi7wqlTw9il8wpf3wmj3jx+kQa49bMlOIAu4KUXz/6I
aBDKgy+zcTuUASCp2p71vPEEuQJNwVE+VkcGEsGz7s2NFC5ILoM86jkvYfZo
BurHIMnBg/xCMHDmKoYo30N1KLvar8s75OFpEC3zI8c5y8zqfOsOK+LId07I
FYZpb6xIsAs7cfEjpeRwSXcKsMEBDsbPHt065ZrBIUz6Mt1duJ6FkbSfyr5U
2O7jnZIIdMVHCPWazh/K39dcU7+Z3VnmuxVmiVBbG4Qeo0ubj+Z06Lq6y4g2
L8HxTzXaSJi3xACeED8rYyVYWHnaKunozx/ZPtquASEFPtDQEGfnNgGL8iid
Iy4KvpONbVxFqhoEf6vqRQ0OlKm1nb4M


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
MVJMjoAi+lPiTYOIoE8n8kM2Wj2ODk9lcPrjUD22n+zt4dQQP7cjjbu9I6CG
PywUBwsxGysvFQjCn5RTO4AKKk4jgMq4vdEuKOISI2XgKNwPucL2yS8BvBQH
u5g/skBrvkZJHjCT0ghLe9u8SX5IJFBtEh3LkawHgG3VTJ+RzVM=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
PCC6K3a2qmHqlZdiDzTPXkbpqJzcIXqyOfYEKtrDNhhbbf013GEG52IzOL1P
zBHdBHr7TlXVWfp8ADcsA6xj0Thj8opBtIYsZX4pw4IOpo55awHfAA0pKRWJ
+b3Tj3Flql6M4d7r8b1R+COR34xjSSjCHhfFOXc74ow7S5jWYKs=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 23504)
`pragma protect data_block
cI3Xn3RsjDA8QNBOmEc1T9pBK4KFWXjplS2G/XdBBzXsUBC3hr34sR9/j0+D
SD/Rp0zXoDgE+zsorylo7MWatxBqqVtREeHUXtELW1pOpdEmv+G9u5jSe9e9
dkF6HhwgLrV/Owqd6LzoWOWQJWM1LAdBvnyMjbsdR9z2UafN+F8cPH0TvfpS
WOaJsi2F37TDJiPLCnXmoXq/3wacyBN8hP3mRjJTs8InGz6J78ePYs7JOwq0
PgBvdmFsKDUzVH1U/3ERp27w+flBxnoIa8WqYy7V8jEaFFOF7N41KE9mOb3h
Tp6oNgmPqoWvqYhQez0lkG+Cd+KuRxKb8J11SXcAKoa2IFM+PzAQcM7Nn7Va
YfV6L3R5jNRs48/wC+TMQpKCHtY8AyDMTL39Y2pzLYTampUJqRl3vteo28Ca
GHi+MPTx1p9DUAs/HCI/9V1ahHTv+AJIRhOc0ASf2V6YI/RHz0RY6RCRBb1A
Rcsu2asntRcPupnwfFHMI4W4k8tiKPipghMQRUmib6XC64wpS5UdRmUpnxEW
P3XxVcJdLPNx3+mwDsrwXXXIn6hDF0yPYZoFZkraSc3WYDwYEe/Fwx44TdBx
EF7SYCn3zVn5QweTNHHa1pdam1S7YPrVLSb6SMiMWAGEGxssylvTdaJu8q8I
Bq7HX0B3KVFH2g2Cdzxx3ZYQ2fuPCpHDQSMn8ZwRUuYXZW5gULNT2eyM+YOS
pvm/LX+esp9Pgmgop5efeNDhjoeeUZi3WwfUqS6voZE9dHqKlW2hhwTvkBWi
HKFzgV1hu0+fF91MVaCN+atYC8n89pDLQfVYBvoVE9D5IR6M9MEBIKyWcnA6
Z03xN1NPuIx6DRJyFXAHLO0zbk020CTGpBLcbCE2rbWih92D7G5kWsBzMc5w
trsuGBnwsyt47l1msAJ62pDS6DIJifIQrSHS2VjsCKxVMDTOyYuVA8ZZVXZN
RvRiQfimwGSkWg4jCKm424xSmyX1ncgCpvWmof9lTLLu3qVB4wSDbRLYM4gy
KuldrSbReiz1h+RPAR0LcnPPYsoFdBDhp0U1mJSvONIqagJnCGb9C9KiXdYc
HUQMVJ7cW70NnLDruANxYVAL2CiK2ln5Zj6RZC6sc2bAzZGxc2zZNFV+zpEg
vdQB2jHdct7OBAQ9FaPp9GlVqf7Dbw2u+mZBF4a29L/vNVf8sMhXo5W/hdIk
hy3rmOpHN6SmftGRFxiD3uQc8CgJ+WBHMQiB7PeTGD5WP9AU0AeXsoi38l2k
CenX6e7SC/SJBLYVJd718Ny1O357NPhbh9yOItYgZLmIhkFmaM6mf3XqjtTr
3RKfteD2DZpLRuy0wNFO8n5BCs6+D8GYJfQLT6Hr+GxT4Zq2JfTAGN5z4F2j
mseIlOyqA3GSf/3Zcd2zaKJpMOxLa6+HVYPvONWu7dZgo+dZV/iGEx/GsPZU
gDjHioQFbuWvWmJcUXzfq03S62m8oQr0xltz3hAg/RXVhgK7jQZqH9gxvylt
tcJVdihNJo+dJSRP3FTK9wR8A97FLO/B8jmpEJI5fil4KlMrR1vE17Ha01le
YPjzmaeCqtDrl06v5p35MpT1uGULnidB3kTiTnJ4Wv+1nl7pRZzR9CkqfvPY
b/MvnCxfdaxgFy1clPJ0cHF8Z8TDnEodgq/0Xs/hVCQy35wKfh6P6fn/Bzyf
5N4ngwfFzzSf2bO0xQD8t9vLP/AS125ci5kuqPIeaeJBtw+cTji5Tk8//P5J
T/Hzbxua2kuGU96OtiNhTnVW8wIgQT8sYqIv7wXFQB2Ko6E1MNK96QzC80iK
g9jmcME9rN2gR0fxYbkykjCOuAOxWC1BuGfbjj5AS3+To2waDIw6BBAGQm/x
lLLXXTX+vZtniJ1qOf5NtZkpb+mvLtxWIkFnNGiethJ5+X2oTSNV51DySWOo
8av51287hmvesUDum5K+pLL/AwwrwXtLzjqwZ0F0Y7/svNix1+AstJcv9SPt
SDZ7UeWCvut1HrL0InD29CaGUJ9RHzQZgk9YLdyYdSME1RulgZ1PgryZNQi3
ftzYuCtn+9BSyKvI3f5iadQfXcrDsXCZL7vo+fixRCGmq2tQgA3EPCyVwN5T
OqcYdrOTzlgEWoyJ0e18PFKDuJYVceE3q2IQKuAv4/FSQvGeNPOq7oc6qJLg
vjU6IM+ozjf0VbB7w512xfOyLWNdMj2wVpf/HQtoOxLJlE5fjrRRZFwU6E96
aITDRDcIVia+Db9nzDPm4QWayi3a+JzDtmRFvt8oO9CbynJl8X5oRnFRjQ73
XsdS9Ebm6e9TCklwoODj8MI8cvgrP/7LEmlOm6rn/YosDzPNohtN0m29tjlP
FlDn8a7s6uynhLnnC77FAn9YbyhZrFcl2thQgkYTGyCzSBh8uFO6Mg0bYJoo
CwAo5LWcHLZJs59axxm6ARbgPFU8B0l/wQSDHPGmu8VBJrMRD/tv6PqMBrRd
JLnUnCGKSb8aprdYnEiko4P0yhgoc/Isg3QBr21BQrv7iQyVlqeFkAweS02F
TSG4+nfKpqQ3rhtFLgLNY0P3gqFVbBfKlHctJl7LS2SOyXxfjWefyF5dISDT
99Q0mMy2oAMmVCnyaF5j0LJyhZ3E2QmoXBWxCfS8odZGNdbfzxoI/QWf5iKQ
DXQgkPaJXcl22OD8DLFcxlFsTgNO2HoZt0963O8WuKDAAJ/4ZPtplb+wgx2Y
wRZlcIsLBpDza5tzNsOnjZ45iQ5wlZWbMmZbpAuzupcZ6qbnmQoXqUBCV0ah
NUb9BQlrQegbEPmy459lEJbHkmGElKGfmAhyIfLyFDsgBsD9Pb+33NFuYlk+
H5JpR1KB8iRsfZ93bAwE/ZborMylQLDlto/thrZDJ06HVIStOihDqHdcwBNy
LoJFtbuY1BxKVfUZpIY/G+M2e+sKXfw9G4mwKP8VDTLc3wLg8sJVdq7SmibV
yCbJZGfE58A7zs5MDPADR9NKrqxDeIXhPTpOPoCCNm0SdyDNwNSt4Ka6twXD
7+6pIkQUJrwjdUG0Yw6E+dYg0E0wCOWr7hCD/9UChtALuhW1pt2o0uR3+iM+
YB/3X/BwJk8hfrZo+9BZ9AqJJfC82Qn0lIc9WRQyFsaC6LdgGJrKONIlRk8I
xuGlylf1ipTe3yibnUu16AYDiXpLg4BJBErR9sdWCrR/MUe6/Q0AWyqnFJVc
ppvtHDPqPfjXEaNUSBSYDO3z6FWHEv282OjlOAbGXLvhrv6w809j+Rct6PsN
BZM12d+5gIwlpo9vepw4iURk6q3INHmPBLMNibgACC/7f4g0ddxug//fOjz2
w6xiP424Pwr2y2OkH4i+vW+OZfZl7XbeFJrxIhs3xb2AgfMXYKx4Wdbbm/Gh
84i/V9Ahff8zszVbJy76h1/yTl4/CrzBsBeZtKocx5pHmvPjLV7bDh9Q09nq
whkOaen+hE4zTn6B1zm8n4vLO0U+8ttGE3+vaRmszZQ/gIDfgJc0kGUfkygO
KUFDwT45AsuowMpYaRzAeUKaQYy9TNmJYWAo5vzpLn7ihwK5ErZHZg+1Myyv
y1xa+xjeRH1tlal+5C3uMwNpgCAdxZZXe9vKiOD0qiGLoc2nmZ+RdRrQ0Mqj
jbWdvHyyYtYkDKZ7waVTSlMbTXVEA51mA76sM2fW1tJIKjbnEAwPaZ6gND5I
kRtQ1FbN4/47Ajkj5Y0Ot5Fua1OOe+G4qcac9azOgGpZAo2wUXMxuUG5mbUO
iq0Im95vr6rcOn+i7ALRW8kbjSwm+u1mFKDeJuuCkB+0tOjjgAi9XeJcrM64
iRiNTm6m8RoF7nrBDOspua/mK3JL8ZQIaTIRdbrfIMog6+znOharGMAlzMDr
14jeG4xeD5a51wC57HV78Y3mdJ2mYEocPq0ekVHIi+lUinc7I6AgRAsb3g8T
ycwy4qlGizmWmhZhEVQPfzKsWrXU79sSeA6wH67rFLVSCpLqU1Le6DwxhgUg
SR4xJe0f3jfY5+2iduvbfB18sd355OZIM5FGozkHQPpzUFFC/hCRB7AHrVxZ
UQwJahiVEdpv4OsGdff/2fF2AqzPJV6bS2ZJB7qPXtNo9U5xFsSv5OfRqCfd
Mwgm860CsLsoJYAzP7Rxin6XfnNTxqePypi2Moik0H9oovkTsZwjnBYCOEkQ
ucde0HpLkIDvwCMRh+g0Ar6pcEe1bpdYwce9/oEGvYKPErlc2yNOIOOn+G+r
N3NcB7VmhG7iEa1M8RlTO0WR44p5qzKW5+kjCiZlt5ej97Lxo6bGT5iUaj0b
K5/lSJk/+5Edbw88foxogmtiiz0RqNRwEUGcey8+ovfr6x3KDmO2ko8/pbAr
cUTP+veTpHXCpD50SKxIMP5Kc3h/mizkn0VR2HuhaMUsM85SJi71UVe0wA27
5mayDl/odmTsF4Jqo1NmVsFsbeZiSViB+bleCS1CJ7QCjp0QOxt3liLyraPy
SkcmKEDvXoU9Ru4TJbAG8bcAmQXiA53NRaIaRjmTMpyNt9pZg4TZc1okKvyx
M1g//tYJhFM6a2g0WR+mCboczWmbRjB0uSo1i6FClwOvztbQyra0R1Rq2Emj
uHZ296T9ldi4jhTVzR5pV9zHb3BUgUxUL0jfro10RuXK9FCZdFoIEaF/bpmV
ddYJhhI/Qo8AgOkD4PeAXaIUn5IfrFZYItrjU2I1uKCOWBTVMURmm7dj+yTZ
7ff1SrSFtnapYcZVthqaVVslLpgdNSfLKPha44sYo0x1IgdrwJ+xVE5aEz9S
rRau7+qXLQFmNoudVx3ld9dSiQZjroDAiRubbPSo6faMx4t6ddiaw/R5t1In
mNj47n8QxFJuW6LzKZ+bou1Es5XbA2AwQIr2Oh6xp5vHMaxaRiYWJ7aKmbz0
JJ3q2LyqR4ciOSwvYcFunKKWj31T2fBJG4GxyzxqNbtB/poFsudpRxhyG0SJ
93xhx7k1ebyu7SsqIihyBAl9hhU/0hZkqpZivI7g1+vk8U8FY4FbF0qoClxs
t+7jQZ6Q/52++ablDXCmV2oAG1PqCwNSJjYLXKBjNWe2C6CFvkJy8c6+8vZM
8mOAj7nRpdtJy5O7WuBCfX0Mcwm6cFwn5oUsLRXm++l1C1tbzq9rxoC1Av7A
HFJgBqU0jkT+UAI5xr0JAndcuN2U0pHGrsqdxICpEh/EjpGMzpsP+uNJr3YE
H933iTFuGQBcy5n7twbhhFpt/bYxWTNpRT8rouxmjoqJslmZf2BKQoqpAYGL
DgiYA50M5rBRYhjXbc42J2tAYRhYWt0Q+7AVEN7E9spzvKI/W3mep3+t/zOC
lJsls+F8xDG7+hz0UGe1FcnBvXwA1t/HUT63y29elol6f90P+joPCkWcqNry
YK9nx1zLZwN3tF5oZIsRK05Eom6DbBT/BnFKr/BtV4XPTr0llu0OGA6AQYJh
9/EZhdLhnDLEFBS0OX3viZysmMtxZfi59AEETm7mt/JmoYX4SYytxNtdzyU8
M9bcToBqXadr4UTMtPOhNHTTdDWAc8YFlcTeTpcO8w1s7sejheyYVufoyvhz
FquBMp1MNsvENnxn4Nx7MB2ezRcFnD4d5ZVY+uRgaIIADuDF1xIHIJB1w4YM
uW6+12Obn+Zu7cUPaXicht2mhjFjqmdirox0vWbdky0H/rPKBTIacLqej1hH
NEAtgvAnSRMF7eop8sah1+I23lKvQYOjVGxmY/h7WnAdwx9bPhI8gmMqqTkP
tbnB1YpVdRRx486PAUZsqQwZsrVlu97CS4Hs0llj+oAha+HwfBwI+gN6wCd2
OQfW0yz2gqm0rBka17bil80FOom6L+EVrNNyBkstRe6kQVQwCTmBpR2SxSVf
sl2uA7OD3HNDEXFhkdrimNqyrCCoRzIjewsiH7Y4TOZ1xm0d7SfK7b8fqTKb
CitF6nDtmy2ZYHr4adf7/RqP6bjST338aEVix6omaFadNcxFh4GKQDKDI7BF
ouSC4elt4b8HT57JBTUjn0d9uXpxCz/mossK3GuFrBkGjDDA/0SdmNcDOPQ7
H4xaSeu7x2m9vrZZUIc6/GziPw+v+5oWc966podsqpoVrS+OgSDpVy1vrl30
LEM13wF0MUIGuUlMslC3j5osf1JqroAOAMOHVu07MzUduefW2rMRgBqIeO8X
yTLeCmm1LCYMd3Hg5Uz+XK7IAhoOE0e26dstrOVyurMLYzZB+yQd7OYlSOwA
MBXP3LGK+rm4nZegIAouPJg+YfPNvc1gyxZtSc6SecdkHKtudt3hRggNZ3QD
s0j2bfPjl10sTzO/P6ZUdBoDm/To3ItwuqUNwCaYTUxl1wKxqPBU0ASsvkRZ
xY48OJLk4EpjZL6sjpGYTIsNSW0A7lgS3EKokdStfFp7AoMqLdbVujlGU0KM
8BgVW5gx8P2qinGZXlmXhZ4RJuR+uslRBQl7wXmJPEm/A9HG7SNCBqU9oY/+
TQWlENveNNgzsyhqgniNi6AphyfUngGPwNyb36ad83qWUo0EfZ8Tv1aFTMZN
OcYGHkooPeIbtupfegbKS+sWzimtu77zj5qp1GVX3nCaVO5kn7IUdLPcyCzr
kFUE0Zhms7o0wQoZds7A1I++EK2ToovPTlm9c9yxRDUHKl1vo3oAuvZAiPVL
AuntnSZXoNibhuOzJobXSnQ4nmpNP16UK18plQX/Pi3gN70m0N+ljTuwp7FO
c1hynCFRYIPGYDBlTwkEj64b5hH+CBueutbAQ6mDs151BeCwP9pQahvtVjwu
SketBlAwFKjosfwnv3poygtUiOB4ZwtNKgViKVsMe8gRizpV2ep4W6ZAFIBV
XQ5S6gJpnd5hjgPCPIUMB6dcTCzFufIvffG1dFoix24i8qyruFvrMyxeVi6K
kOh6Uf2GGfceV3XafaOXcqyV8guy29Zz/5ZIZuPUNUeyNvgjbElXVuCkIWzU
DyYjz+86Jo48auvw5AHfEUYI/q9P4RntkQVR580rx5SPpI66a3+w8TGwHvNr
cVfFdunljz8PBqLTzGUwcihbC95/l1ALqjdBiQ2qVdQJiqS2dmT4bWAEt3Wc
FTyKfzPd35OKxZboWHyf5BkgVUWLFxX8esArMD3KX2QnXcIS4apInyyGNyOg
JqedCLW8hAitXAcg2hYVawI3lAfzTh2ODV8mHe2Z8fYBqbCIBhFuvYwGv4Io
8IDPvwfvTold5rpP8AYvgzuCOO/D2v+JlJ4u7lqAHr1la/PTFrCrqjHy3Y4B
kX7hIxNtcGS7xl4PcLVaTeL9Sr1t6KGipbTKcrdW0n9N7Gt4UKf707Ln/dIb
cxmRRCrF+OsgIpGwval3WRqaiLrqoTscdkml7tGx5GEBWhTifSacAvh4JPoI
HIYDCxnrUDOhhGH4GVJq4mPHSlJest+4jyZrFlL7VtqIpT+wQiAvz7tBaZPw
3BaQB1xB4xclU0/LaFdlBc32rYob3kFZSjlDJpkYq/E9z2V84BRxYQmBAN8J
ERFHLIZlDxBsZ2KVy/n95nejzYYl9yI7zQ78l9Dv0GHe1bnKrdBMCCg2c4LI
GrkhRADP9E7Vuxa/9Giwk+/d5m00VoE+mzRG1851aNe/8S8sDSA4iAOvZb3w
IwRvJqrpiIsocO2GlLKE4PjQ+nSSLhvdalwhDfOGKCiqxxXmJ1dtbBpmHnC6
mcEA2f1Y8MR5nciKv26VyVGkj6Kr7+DkpccAc2SKe7EqEGgRZItSea4TlSzm
XXmmIrSypMV4jWscXJ0g1ZqioNzTfdERYgWDodwXW9MrOh5pV2vPQ7enrQkE
0iv9xf7zesO2N9HXRimPY3XJpBsTMxoBMFMTEMkg2Nxhn7XOAsqs5rvmP/Pw
ms45bBWwifaKyrhH8pDOmiaKSI0Mz040WB0ulN7yS8k2N401wxpWq+MAWfo+
nbweHequZfUbSXuusPn5gHdIpYpDSjnMMrFBsrW71luIRCn2PfVWFIYDoEpO
8NU/uNCIEr0ASduMQrrBtPGm5kc7awq6h6QdJfcbbUCgTyIZ3TvnnYjYSQTJ
PBO+hk8kPujaKjZVhL6D93wn7E3MBPxbaQoVQq1Ggmtp9vYpp8TUq8fdLif4
ivlllIqoXQmitPvzq7b0p8vUcAnMc1oQ3Mu/8wlgoQWWK22Ib54SorbITTRS
3XcghQ3hNBFmG6OFE8RgznLVI4wTBjgqILO63/3AgEbLadR1Tz4I4UNn8L4M
nzfLTpl6RU6X2YKwWjlPuFtM3ehrKqY3pkbqbWKP9i0+uZnoT9gor4Ay31lI
34G8CcNzKBUyNA+OBBq7PMBweXZ1HyGyhHwO9qUykmmzwqg99u+nzpXXkNOc
+uioAVg072YpU27jw2kTDboVd10AQzVf/A7s91xgVpZN1c7rzgdKkfjiqZ0j
jxUiK97hczPFN/NzmCFylyQGy+5ELFUYHPk2AJT/4gX7x7Ip5KI5tanqk5Ko
9CSt67ilXm0KqPwBNPA0XaprR+cqCt2/ESUYjsGKXzDqyy+e3bkNb3/hTAgW
05tPDr9PTHZ0YDvcUY2xQtmJLZ/bhdH6RzGvfRQESzGk0ATybbDlCLOAdY85
jf4LlMKqAijG9W9rTSDnUU58gY1A0bWorN7OTJkp3zZoLG1aqn0hHV4mA4+B
G7nhE1AW8tE9w+sHKfvtQzf3QHa5WkG1453wAST/23VQHnqMP4zgcAyUezDz
FCETl+9TCkmIfcyaOAhsnDl2CAG30DOdG2g1pz2lZxA9i3ysreed3t6VwWiF
hZZVcqUkGS07UdN7nFw73oijYfBgpoLQQ6i+IsDzpDRVYHhbUL1VWIn7FsnB
xM6nBjPiRTUBrvshoGWXPnL1nS6wh28YFBsyI4Jf+bt38J2CHKyBi5llux3S
McJ1jSZY4ovl/OR5Gc6xX8lF6BAcNqt/OMSRiTI/0ULmUhiN5UENSV65pYo3
o6SzmlO1X4i1fe8d6+nNiZh8rrCnSJpvypz5+Dxquq/h2FgROA7aCjuB8xp3
3/xumqWOTOPUkO/lPeDaK61IoHcb/o7mTuVsA4CCIRzOV1ybTjB/LMCyo3lm
jV9Yr6splOhBoQEVNPI0KZbspQgAKIzSebMZXNXMqVYBZ5xvfMg+pwAq6Gk8
CXUqO+rcN5QabBTKjPqaxlfT/+k+SxkQRdIsB/hsIecMeuW5KYeIJqiynzZE
QbEvvT15jANg6E3c45nwXlvf5yFfPScY1Z9xO1ogQ22x91Og9lZ70VUoSzNP
USnZiyRhJyEIts9jiur/cE3ukFmjKGIfx3IFl5WXvWfnN/x0wXV26koH9WNr
svjSEwJOl3KapF3KFP8B4ZKmrjEbFHcFszJk+Qhwe0xP+cm24A3+Kd/dmCCS
ZCygNpVpmB0qCfKsNMhfWOFthdu7qwMqCOF5fw7lPqbVV4E9N7Yh2WRZ9aR/
o4+O0BsgJNqjFdCkiDq2nemSnYiwDfN3xdMOKUgJsj44cTbPOr/XDqM2ggeO
g0F1gaqTFcnmZBdfWNRRloHuX/7VBksNLmWwP5y0bFKpMoPFaaF+Wzyu8B9S
XOLbhmTDoy9o/+/tU5k7NVchP9+VreDK81aazuQVhDUNGJRw0WJ3y8+zzFIO
L22QFa4QGR15pZ/gLpfY9tmLdAQrSb9mIftO8gm+PTivI/Lzr2G+bQgNlGSe
LEKxrV17w9ADyNwk3xYHMdiA9Myzwh6QYGyxFIdfSmvvoz5CyDz/yG2EJn/k
6gyYwv8hArv2UfihhnGeAUJdufWqPPb6v9L2BR7Inq57TNw8RYsxB06LN75L
mbjFni7p6ug4JbYt+CgyiUyG0ZvcaJ6CY7HR/QSSGzFmyE9fssYKDFUeIlYq
POevQiBXywhw+qociWcDXsq0Qk5BudvgBwkRcghfXrDiQdVchgKfR6hZAIjC
kchdxmsyP4EJmmRomSywXEu44INoYhwqb+914EzZkWNHoFlVy6OXd9Ri0x8Y
5KX/BZI9wqWjiSky6/VI2cHgDKMCSjUINfsXGjicLW5r/7fJURyB0w2hDXCH
XQbi+BkH+F54JSF+beC+We1yEPAoEkas8R5odGAGCdlpwZ6wF3uA4zWRqQoV
lfzfJ1+8ARly7Y4yVY+Su0lkd+fPlNngWU7sNCivw2l+OA3+TSVXPQHPvuPR
YgqXb99TuZBronjwaEE1OgUmHz/l8VplKIW4wtnuuSe05bV9ZdMYKtHr35rN
GTqeCiHWNVZ2yHk+cvSf6ClslxZtwMq+4/ftCChTbYhq09PCzPPBjOqMwUc+
HgFWU+Ug4+RX35WLTNuz9lgeJZQ+qwVJZauEIkj6nAjang4AXztyCJ9HOqBR
ExNRs84wGHmz9435xA18HovK8Et7xnJnFGvsD8IFNEYrUEx2XVmltqxH9gje
bzdm8WDWkvxQmLot8tRJGwwl09JvKPLvJDW9t351bBNycm0Kj3zoamVb72zP
fYpPpROUuh39cYjxNBxo9XBseAVKhr9CusRWEVe7cp6fh626wZMD6i2dUCru
+wZy++SQvc9OyuZFew5nQLQJwRRRd07yuftv2RV6nqQzvSjbPIoTw2witNv7
EnPA5zo+vEIGA1cPSV46QEr002kVOm32PmP0XmaujZej9IygH2V1k9VRVYAv
ICcqLpl5N+YK+6D+B2f0w19HSJFY9lh0DoPkNIG5QoFdoVCnSTW6uN2vG+7M
GHdofhB+NWaMpyJ/Nv1PeGqpsHcZqdY8eBV0Ez4/h93leBl0mt70ZSBDnucy
sjd96YT6YqlsE6esyxZLnXY0cwIZf7HXB0qIrVVaLZppJX1+AiispNUY61Ha
Qjnx9KL8sFSeykGwfGW56nojrg+iKV/YopQZcdF53bbmclPUo/inLpPmdj4j
+aviVRWYYRBzJ1o3DAc9hMeMiz2qD23rkFXYLGagcZBLcogHPe3Ek/ZmFeZD
RmZtDi36vr0pJy09OfmsfFAcxm653MeC+Rxz6Tr2CK/57wQW0N48lYk7UeNc
fUtqEa5Z1OV/kHm+0Qb7VFr+BOqrs2O5DJodSl5yKMij+Zf41rgyWrfyUQBw
sIbvjoXnAvHvXskWCUItwMYdWfFTfzGVyQ5RidDdl+XVdTQLQnALUySjKfAg
yU2KrnOPn9TMcvioTuHyikDJrHb/QC+L3Ti8nYwDKaXTxJ5Ehc5erreDAwDj
68xcbztYtls+zHmeEPFcABpyyZ2Dh8sGEbw3/bQuQUjYAcdVv6gigSMeRU5Y
al5wwZ49an+rZXa2QKIzvEdDE94FyfZZRS3R0C5cT4gL/76SRslpN0ASURzL
a+zXuI49v1giw9/FpqxRqLvCF8u4zHIu27MvuKPtz+wDBNqpHAmyJIwyNl5I
j8rKCa5HuO/rZa+wKYPKHMo3pO1z1/ImqqqsS96OwfwWG5Lv3VTmam6P4jWk
HmuaW+Pj2nxImNOwxUJWoSns/Kh7A+LG/QeaOl6ZAGunpECCgf/OgxH68H5L
VBSglyezW4F+Y6bPdBt/YQ+bCdyIPHxqyD1qSpEDu+LjHHAdRLOO4hZsqquw
Mn4xjxUrA1EQ84jyjczzXDy7xYm9N1MYpplTn+Tbo0gEwgf+5Ya7JOqXTfb4
GHOAAvFEbQm59LEMDndR04tGZ46fuC8Z5g/OjqsqMLbt6X3tp8mrAWkfqg+Z
SPyzeWAqZqNPHs7a1o8PAwrz4rJ/pxIJcXgCiIraKBNmTXb3P+CdT+zz4L0I
8uUW5sT6X3b/8orKzbI7B+81iV0iN+NVM8eS4t7i+vBo/2gg8ml+Im6vXO8V
pYi/af84UdRBbyzyG/sdvcUOtXwMB2QvTg6hCgLq8t7QwslrZKciBpP6dTQq
wqu6WOscrxCZusf2v3NQPxzX0gFBB6apqTnpxmNQ5MG8BFCEmQP9Cto2CgAW
D0FME0YiQuwhRthEQska5yvH/6SKDNIpYehlhPfUMEf93i+e1+bGdp84ZDLz
ZvpTQc/Fs5UNo3Jra5FqLJ0GszM2rCkGSRWeZbvHGIvsII3zUnPBvlWYCBZT
PT0ASMsS4DPDmWOsvrxIynP76YuVXR01LXqWJ/lNPd+jcXJtc71Xxa5sqPYH
WDKLu2xvo2b1fyRYoT4WZ1HUk7iB+pWTTav8FDoYpWz6gmEUf/+1KihLoYfI
kjmoHL/9Bxz3udYgb/5evhQOz+F95iWKpNjC35QNdB2k/S0RlDvIHxcqeZnJ
jHiGhdztqipb5Q4/10tB+Ssj60g2ztTOn/ApSUyC49oupIx4BUkSXCWQ+RuQ
N1A1ghSDRm8eirX6toeNm6Av1xzZve8Ya2+8i9/MeN3+zLDP5XEUEtRBjGxp
SqE6yDjnMdIfsB6phhDatMk3DW5IAxGaAm2wuFpd8b4iz6+64FwSUpw4SGGP
jDVzfDqM37r+pVfdiRlbuGb99wdjC54V1QLP3Ozi3ZHBItb+Ym0WDPYKxcDR
CxmOOfus2SVmjzNr2h1LmiQSG2zxyE3LYrT+k7CC40zISpe9ZNuONNaViRho
UfvkY9hspSld1pbl6vL3etsAhUnNj0GmAfX6xshRbc8F6yirHiyZpWCWDlAW
wJaReFUGG/GetO2y7LxE9bfBUt47XwnfIGRCi2g3uGU3K7saTaI9jUFAA6OW
WuMoXC0zQF3ahm3Gh6jp5em640kLJA2M9u5Lw0JS1VhjYrmSdhxuC3/0SRoS
uEUWs9fuM7x+yYz53MhSpTRVi/flIEIW3N4CVvX2xbPm9f2LnKDlZfhxZsdw
OrVTR8sGoiHOZirIbdumxFvbkNk5pB/zHjnqRMRdDqY57fckVsglMjRxXyJw
0wYled7Q7y4YsM5C5m24jOSrqefUpsGJOJ9V9bNpThkraPggDWCm+1pmDLwY
byEG+Eh3d0A0szBqoNQshFa8Bjqt1oO2bomyxhpBNL0sOtrFB7joGMIaYOvx
FqMplcgJBAVoyrHO69Z0BORrTGCIw820owpVgVDjw+nPUeNnWZhqahul9pi3
AVCuwW4LoGQvmYEYiZedtn6HbcZcQuT/Csv35xYydFTpv2/mQHpasrDusTqc
v0aZJvT456IlF0cjy2x8lUNOhmakX/n3Cu+EYhlVhL3xQnc/bbk+cBOu77QC
vVMazV3MGjxyBoxw07Y4zTOrWM4Il6JqPAzayFcxiDuIn/yL6qLsKbJ+ZdEL
LwfA4tBngjF2KIVPyHzs+2fxkZZBsoXYTvRrDxTR//3/y7+M3JNyJgwaK5Rx
iN+JPOJ8kcmBE20+UnJ8+quGh+iHUhzeXlSAYUKxsmNqjgcMx7vjtcIIS71k
x92Oi2N7GCDn1WMQtQJalW87/qAbLAYIJ4TMfCArpPib8HZghT1RSCo9JQ35
e+fs30zWCUkXsNmuzDLKh7vqPBVvzWhxVAPizSsqxDXqLCKwbk5jMT4gUJH/
1SYDImosllW6pA69fmoDtsBgvLvTop7xU1bnjg8wOb3WZMhYKRilAh3h/UtF
YijDOBewOmeiFcM4N+cPWdj/TNxinaYMw6NsUV31M8WUTFfnZojKMgsPFCFh
Ddp3GdnJIJv/hkTVc9mWuUcvHhVYgM49+7sFlzR8tlIHOAd4XYCgp4QKKNlz
ZqgdnpZgHK27CFZYUaYg02dgGhnoZOd8tbVwoaQw1s1M5iysQTdY9OlXf4rF
7skfXCWh8Xte/xOMaEBEpJagxdrweDTnFX9fK3ek0Je9IxnX0or2Mh92w6jh
o+hw6z687pbBqmT823ezk7uDQnmAmEk82vjfWG+FObdbu6JObbSPggrnhEAu
Dyvm+FBdoPerOBojYz3nf21v4CNkMeTX8gIPoduEeVlxPza99f+WxBqSFkVl
4ZOlb6GYD0bKjhjClD0kTi4ZDL/wPSimqD9ubNuu/s/B17ViLPKFEsQG3V85
xaqSuPnSBWDiWIC3E772G5t+1+H84LBL89fZIlO434rv6R62Uf8/f2mpQOC6
Z5Xy8nSDhDuSxDRKcfamaIwAYuxY7M4IWleDloSifZb6JIIb+TXc7vGwHAb4
6Pa3ZJQ6HwoDL1KWr9JdmlucEnDbRii8er/4yw0cIkRt0d9hMP1kY+Xbmhn0
NIwyCzHw5k3Yjqn0BVmEW3wZAFgFCdptuFhWyWIaPwgu9z3F5tLI9yx6yX5J
h9iQt7xmBuoz2O+v7sTClSezHgWCTNzSGyDtfgA7njjxLbc8jckOe6hyyrIu
/a7LlHPlNfr9UrUK+Lv6mTRexeP66e9dc/fXjanz/JfX4KjHUs6YPLXfVO9J
/rInVAjGFDViqyki3j7NaAWmZZfcFLZa0TOvbSXOz9twXy4g+F96VOwVMIBi
yyINbOdTDo7M15fu5mSDx4kLbxGVKm0Io0/OfzVMUMoIHpAsLhKv+t6BEsBJ
sfsH2vzx+EnOwm/Kp8wpfZ8rnZy1xiCo85qM89D9Yji0baMPN2q7ZZymSxoc
Uyq+GvMLLf9O3jTLT2cGt9KBYSQ7PtudlbWi9Srn/irTndV3e2H+ewyBnA1t
jq3sAIOHkop2XPtNQbfODWgz4ciXfLj90Dq6z96yTQX69Sy5uefuFRRlGkzL
mZgENsxHmejcauKE7CR4T/RRIBXvvbRKb4RKcvCqn6Xq//NIDK2Z4A76r/N1
HzZgF4f214/hzri5thAOzXMpiNvIGNOssWjp/OzyySa6onsdNyCMfFSPgjhJ
xU604QPA4m8Cp3YD0ZHEJk2pe7I2arQU6NaqJNO3kATUo5m5AHHtZOErVxvq
L/6wTtMbo2TlmQCKVP+VoIfgzvEo66krIeZQkY+Xo5ucE3hMLt2lzf3Xe5w7
xzLmrftClMuocl1ngdLm3Jk57FmXhIwsvuyke+EEGH1qdJSoxzBnclGuzzWu
9p62j5gl19eItYg0esREh+d/t8nhD0yPxXC3yiVhTxMhD6AioXDSeIVK5Zik
WEjjoSAeXewZnTr0aaAw/9s8Cg6WGshwcs7kk4t1RRe4fzL+8xidyU/5fCDP
BQIs3+ReExWf6phdb7G5NX0k//5kAtjdTDroqMBURWrW4GjQWHRW8USAIkkh
82y/9CpxpvvpZgDFvMAdQcht+R9Mrk8Yv61JPsxMbzSlyXYAIYZqgUY2Jzru
0ioJcI/Qvs/JPLyYKTsgDt+03OPCKC5LTyTfBRjFzgpknc67SaNR7RXxdCnK
xNGtVK5R8aGXSC9lgKZloiweIzetcWPFgKiy9EoYZoDKWMCweB3O15rAMzuL
BSPGtTHv2x1cvp8hO5bF4P5ibfdReEVMZHJmpu7uoiQ7CtyBgFP7mNCXBNZU
8kkj8hMMsIG+SsTLlTwYeJ/rQaBbIVPhyHWmE7EpqpE96Cx+xCHsxunojJWB
GW80R2NW4a77NLlgcAY9dOSHgdQezF45sFLY4RkWt12z1r/428FwfwmwZn/a
jHtoqAawaCGOTc4d1TIOIT0CPkXFHP4XGXb4tPx2HBbD33Fg+PJYT3fVeKrz
1PdvblUFUJ1g/qhb7ceNTChq/jTDa2himR8wq4BBme+fGsEfQa8+4Cm4Ycoq
nN485ViO6pkjmfd2By3tVcejZF9Iu30ynPZ1XnYpHWBM+sR78sjOACqh92Gj
Mmlcbf/DaAPjB2kSwfmvzIq4c/uj9Pmo9ecpVhIZNu97pMjPrMv1e3MR0Ity
UZ5yUDotW+Zy9INL19lv36EyvsrI8cQJ50T8sS8yWs/yC4W9HpVPXFlt9PWN
1i6wfb6V1HjoWunUHHwgv0MZqVF2GgpEzYpWw+TJwszKrQ/iKbHctXPLZFMj
ge0RNQef6MUkvM+m7Jl/pvAcxoV3M+qwMP6kez/dhA5IatGkVRBUXPcIpzd1
sJC0R2HhJdjwvh7vEeeOqlsMLeXkjgPQefram8HcCoNOrex383nmwATvqNTw
sbwUxn56zgOSY9PyVx1jb/szmLJ/QQmNQA2M69A6m0ibIY2azCAc1mn24zlk
8zI+Ras6SIy2ocXaV6RB6nvddw+wcjvhJXMQhH5PfjudGn1uVVlDcZY0H851
Vy5D/HkIMgCKiRPQ4C4hSQtrsRwSoXLAofW5q0MuV4oKo69qYtGwtNwoBAxd
vmVRznmrlXYO3b2OPpXQva6Zba5RwHz9bhlEQeiCZNjmsr6BDrsFhLK87IUK
MUbamuI2IQt4+KgOygVle3H1VS5ud4LSnOnhkN9KgHnMAObuMSxSUiLApBkL
hxFd6WBxQ+ZlgicW6ZplGOH6MxYtYK62S+WIhMPjYXbNgvWMQfsxUhl9uLkL
zBUqsAZorjtLMcdYud+uLKLpmjCiXTr+gaJO9oL7vEApkfE0j/Rjhy29p+da
Vo6+YrU2zxMoZ9XqOf0qg/PO+6rTqaVY2iVrjgDx/A9Qn7EwxiI7W6A6087f
cxBzraO/g94v0TYrI/PfepU9hE8ntL9XnwDVjs6R0Dud0+O+XDVMbV2RJjXp
OIeQymF8ohibXkl4hLLWRF/9m0xwBtyUKBf89b7q+/zo4j+KSkauadb+VO54
S/ksbIljbCjyRj3ncr7B82vWJtGAutDM9VZjd+2kxabPeMr+QjyMKPGtHxHG
Ad2ZlBJhKmYKi4Qyh0UVIcLeanTL3PQ8OSGz9A595cUNtTKJV7ZHNV/QPNZ6
jFSb+Xrx0/IM+upC1YvVtBQ26Fp47z59YElBtphf9EP69A6xrMyaCYNr8lmQ
KCrHfaf3KD+KJlbx85svXmv60jEA8UwAoR4+5CdR5Yoi73yJQSjwqis+i90k
y4oJ+3kYmmoiytobo3+wnWvI1N1L6Rj2OT4Tvz2/DhJRG0n/dg7MN7Neq5pj
1mk1MScqFhNZl7S4CdM30/9+ep7Xed6WGCVHJUV8FyWcT4orkMkSKvnQWhWC
eDy1NIx/7DwShyWMjmMHnYFH+89NgR4Vh4PrG7tR25ixivAOMv5pZheslaJp
i8BTfkdMaknNXcH32Qem2zDH3APP1ah8xVdxa4hqqzq3fG0GUDecjRfGdj1p
Brre/A4aUAnaK6U0Q9pllxAhtVRV6uBxjpDpkj12RxAd+62YJWt15I2KDeqv
TBwcLCoWgC55+QCcKmaIWSCdfcOJhUpIrlidXpR5Sp6finogshZ9JUNS5wKo
4uncFchHlmmrJWX1qQDwV2Lz1M2MSwFvojC0QD5iRXFVGP6op9X0JviEw/IJ
QYnVA0Hz/upz57v/C0oUfJPkrAQPvU2UNTaseDKehbELLzTPTdwLGlTZNXQk
2FSzqF9c1pHNRaiuwM5EKgQ+3eb7cckAKgb6jYaXVu1feOTqjrG9B/tXoOEI
ltqMGWOHuN3nZk0P1hOFfFu1MXDg448AO7VEqk8Vl2Fw/QOw73oyqh35UXU4
C+Bjhttwb2CuYh/CCBsidkMkYxiOSCMP2C11cx/9+ftELrQrztdX/ajDKWCV
q94F6ABn1u7oU26HVE29miiPZfk50J/byiCsSbLQCoc6iN1S0ovlzbne1q3R
WIbRWz4T9fFkrcFnrWVbGAI4T1NBBhBS6FgwjuzU2eTtrIqNq2Z2gbibfocr
RD4pwfQW9LD+ruNK+gd5Mvj+GrogbDSHVJgYS56Q+Ra0AQs25fEESw1PUZae
uI5GF7aYZYCBk/Vxd7p1Z5lhGB5v4Si0lN4qEx5lp/mhsJtTkoiNNSSAZr6V
4n0OCMGxQic3ae7FxeCYViR1CzytU045qtpslNlLFDsKiMrOS5wnZINUkUVK
iIhQdIcp27bGOhBtNqrntH7g5DcOSnC9UO2BZ4JilCOv9Da0ZCTbTzn216S1
AedZPPOwD7etfF/VwqwJgyCHD8Rmom3Owxtv/+DuImY2+JPXNaZ7JRG8X/Gx
w2x7ed9w30+SB1qcgHS7UrUvtdxnWiPNJ5aDauxXZ7qMUKgmc5ATRYQa8usF
cM7pC+fDqLRp8IY6p7zsE32z1zLz292uXQbOcvhW0gNCsQaUwO/wmAICK+pb
RJSci/vzFPNY6qiMNwKs2t4of2AiWPB6f3pgogUN4u7OOKy2f5ujMV+8JACL
mCXdHGAWFV1sJl1nAEvapBZ21k1D1SQ22jVyQGve3lxskDRdIxphVNxHat/r
H1/LZjaBJxYgdbb0dHYL4k+affRbRUkLn0uqP7kyzRgOO91Cro37UeTPdo4w
7fM3bqKIREtbPfx/9qttf23R2ehs6toLIOE7cgQQ8OiaafuyHClrINyGb9Vc
2rkdfQASjmXw3Fsm5FK97nGcZ58CNmDJW5f0joxB69ia9xGpONqw+iwZvaFE
Qx/5jIwWy4zRK9C415Ff6xczkuU428G/7uvNGOK/sGlEn9jsfs1i95GE520z
jBRoEEEaUKXau8nu2KrdBwm2F0MXFtPmYVUANpW8N41j1eDBcmnYuSQfFE7S
jIFwrcNZb6kTHXlaPKbetv0MKLNVpguchRFcYyxC4l9aHDZZthueSYh54T07
mVxIrpkBOjc+MegFy0foPUtpX+8a/O/M71DTyjkKmrBx1a5KGaNz5U5aem0E
+0qBuJur7x7blZnDcD1jY4LuI/9vklNbCq64GfhnI7g64KhMwyI6vZBxmvdc
KYlYdlHCB53t4+Tpe3QQH+Jxn6EA3G+SALSdxfUWuZtSk1sbH3hIF338wAN+
YOHijGFnaD1CXFy3+XYWFFtieEqu8tqo75dd5D5M3kokML2tuBSp0cfoaE/P
k5svDslQKlXC9AzZ6d6WA1Bwt0hzY1zwyv4jNn/2dyKFwhLrb/mXQ6u2ly2q
8SlqdPHLC2EHSaEa5DxhzhPqaz5t7p62urODwYntB8ACjkv+nHi1NIk0cHO5
kcoP1Ch71ackyFAhRpMXU7K+yWpKGw7zhTsh7ROfCW91QGO6iR8o9IcvjFKM
wzbmxEMHlWzD27jq4lV9ia6c9wpliqsXe2qQpxIJuzgf6e/Q59pYUAT0Pr4i
4V6fHMuLn0kWBTrx4fICCdX0ITad5QM8kZAe0IZxcD9cdrOLTm6H2HJTrbk6
Wx62J1ss7toxO1ZGxe2kou6nH4GH7pk1dQ2CM/wMypbGlu2UrqfFCzgEd9Hz
QGZpMmwPBq+vZPJVj/JYdMBk4c+rKMnA5TB4bbprRrL3V1iVuVOvDOCRQ4xn
Y+6cnDPTxV5qv1BLt89w4MQ+w1yi049pgym84qjxtmEPZiJ1jBozn68j2Inm
MdrRapJta/jePfN+CD780ZzilIY01jvyL6nN+9b6KlLSQH2zF47Y2cSWjt58
uSIT1XcuGVvhqwOI94GM9VzfBaMS1jhn2KqLugW5CE7aHTEiUy6nGiAtzqMD
vExYkg2VK2c790H1kYsZg1iDVpfuLCNk6hrMOisXLvyuhrv2k44RyQocHp1C
ovAh8jqo5tQJil6TGdNuukpgAnFuCmJDQCZqmpouvjTermJ/d8M6PlovXjLI
UyxMdDboJqotIdmwGyD5mdFIoTrfJmyvWaLuGxHvphk0WSfc1bMrr+M3QPv4
/7T/tu01JdRCU/Qz/q+ZH0aMhbvxRlB8sftVAwgbzsUUUQE1R3Lcpw2wGkd/
JkPPnsTOYssv1whmniLzNdRVMd8cP8s8Cf9TRMLRVcDPLe1cFjN2Q3fw9umc
ljTvAJXz3m5S1XDoaOseKNDuTUxWGNZETgOyvjukoOoHofie/ytKJ4IgaIP9
ViQRdoDNgwP2dyhFil/8gSQBSiNk6Q8z+pT3hWIIdx8RQp4DGFeVKpGtwTjx
qfrcbYfd+X5lmB/aftHqXnWA/7s81OTIwXY/LPECUO562snWHR9ls7o6AU/4
FZcUnUDOu8ZqFx4fIQ3x2n62jhzar0TyElWYFzoPC/qm+w+fvkRtIUkOqbk4
o5hDiGGB38Y2m5i8O6o0Z8LHXu6XulOPV0f0Rrs3AmvHK4I3FUoKpf+l/Ty7
soE04pkBoMWtiS0BVuwEenzJnHQbDmt1e0+o+aQGmokvJSASW09Fm0oDDb9V
sjFrTZ8fOSNDvrgNQZzot/NJWwQYXQJaHfTqhQh0dPv/YDF3V29NRWtwkbIh
mwVlVdN+1UzjUn5xW/RuxF0XRxfYzy8jht6YOazRXML0kyYG9IxVp2MslvSY
O4ixLJ7S8CRwW9UP5f7jJvywplp3iZiJH5/+CvgBzgUjwbx2Yz7Jq7lNBuar
JZSsXX9eUSwh1s3fH6E2NrUxImx4oqHXxfewQuv+NvHnZrQYHCWPeKhrpl+4
Zei3kjAT4zffe5TDHwsrLPZjoQrm9F3L2fEhH50dfpa3VDYnvuKQsffl5gJ3
xjAXM+qwb+CqnByAoTBPs9AKD0jjhZlU1LWdRYn9Bce20fCkgf0FYKz4uo4w
5XEDvvSEhmMYoLLmLE7w5l21yYMLMXeXG6pKYWV5Sbtx6EyOTX2dmjFAe6Ye
Hth7B2Kr8YQ0mvpDKNpaW71pneLKd8GbozbsQal3wrLg43udi60/9nGVq79b
9EyWM9tR/ISfF4JgF2VWcV5JCYJb1tpQzmt7C30veitXrQUT5JoRlhLw0qp1
c0d2xRsF058jyEfBVZ1Vnq992a3m0IMvs2N7TpvSI30MN622QoUAQr1dwdxB
k2qvTwMBFfIJCPn6bA6/kcmF4AEn/T2S3G1aTzhenXnMdi2JI8xEHzBOOb7e
e2fAFR6hQdkz2RAngRu5kgbnBULPEe8B8IYrWAz4Br8bQY0fszDtmOYj1u2+
o4OjhcPerG5m5mhmu6IcIr+Watqz5+gDG2D7AmwlEIRzujy7iRo7cqa9aVhe
wDbE4HYpZhxsI6P6rBQJ43HqmIB79fnHw4Q5kke+0PMu26fuuCeyn3dc7pDO
x4y+65sYfG8z40zN4Xytk5ez+2KwVl35k95ziSBSkBhVa4zhLaTEr/7t3+JL
nPGrPgDOUm7aZZzRc8LCNqOcS/+vQS4uaArPjWhOBAa4w2BSbhrmpkAtnrYf
ORO/9j9H1l0+jfe6swDvO5JVOBRRHV1pI28tehPdE0OBPbRLC3MXVu4tYfk/
Z1OmNQ9v8w0G2kLol5rJkT77ia9WFSbPycEqHCF4cNWZAD9jbLfQKlbO0Hpr
VQMYm6Svg0NMlJtEiUwISkV71JOHspQIx4mT3aenb6LjsN6xbGfvsmfO7qov
w1AA2slyFbvQBJiIwA/oFZC3GQYm2ZQq7X1a34mNSL16IzI81f5Rvf2o2tOX
Nc6nzwiut66f6XS4skWaj/lVoldTTu5oHEaXM+Moo5pfhztrmiWg1KH6QbJQ
ZrugTbiZ7L0TXddukenVZDEe4V8taPqSrsflEIEDb7UHY+eME+pR0BBMvA+v
bTTQUJmDC0LJWX+07J0WQXZdeQzq8EOzmV2mU9O4gHPjKi9vifV/YkC+hm7v
2WiBRKm/JseL+ZxiqBMcjuGan6vRMfZmyHnR4F5bkqq/JcTFW+rbjS6nEGEn
Uyrjbt4TuI/zyf9MUWRfLNk/kiz+sgjxIyOm/MstUZKg4C59To92xeKVqHzG
T2EFEeDyplX9SZvEQTJcdtnuWQo4pnGuD2S7y0FNrlsH6hSxo+eT++XFKCZD
o1OgkqLyrs61T0ArV1P+jFxkZleIAl31bveAER8XUkiHFtszc/QIiVR6bfBz
O9L0kQNIe541MeQVLbp9oGzFKTVsStfvY9cFRkyu+eazkDImI3LZl6jnyj6y
Iq1cei/9ZG1d0eBPsxNeKahS9SbtbatXcX5cRiIDul3xMdnvugbbaYC2ZJXl
3lUauUaV8+6DDERzd/BT/wxFokBRD/PtpLaa8+rUjFEyYc1iddGQDtP36F1E
uDHIdJ5euf/nKyVI7PpYyjFV5aU2kcOJxaX0w4zXEVAtyh9lXpxD3l70zENR
yrAkYEbyvs8xHRzrlCw0ZDpTgu3GUZOg6PJwscxOADzuC5BS/+TLRTyCB+W7
uWSq3fnga1oSnT7L7pis09k8K1p/rc/IxdJ4HanYUb0VNvHi9SIZGDJtBHLP
cmBvOVVN+Pen4CyIgxWzW/epylLTj3+GTBddLlK8dHjIfeHuwdUwUYIR3Mg2
PqwZD3tYduvWDwsaSnj4Ky9bYuVARicnQb329RXBUkT6haJ9kzLnoHrNSHp9
91lR1PXiV2/1m0HLtj1gcEtVcL26mB8M6wULxHcA7nkkdbaTeSxZzGH+nS84
ftKxfEzMpFxFHM4DIttCfvEHZ/rmfdKKk7CyxYEKUppTUX1qEn3Oq7O7GajA
e3C7DdhhMN4OcMvIVNxJwoQpbxis/Mva4SvOhpo8QiYM66WG5C/bOc7p6uyI
GJAYxDmBD4eUiWuY9Chw3+ZjNHkkHqv1KWR3nXu2zEbZRgjtHnHfBZH57WGN
GoqAbCDahFKlZyX1rupXGSYLS5ynsyhyObKMrdtuSbo3yBi/HlZgN5jvJLDq
Z0bgGqr0oiHZsAbPH6l+HpFhzbAacrzy9SjBENB4aXdeIiledHURsGvsruLn
Y1zV1KcUHPzqq5SywxVbPUKpl08wynCxFHETfuxT8lKXE1qjLOYQQF8YCrhF
Rv/fL8NCZZaAeduh2vFJcbO622nhnJKX2APt2lGFpAmPsltd3paJTAs9jyyR
KBSjELEaBVzvQIwORg5yCW0kVQO/CSzCbw0eXtoMBejUSSRkK/YG2hcTn0z4
AcIsJQ0yxKUr1dlzZCZF/M0BsbmYLxyMYv2vfoXuGVXoo/hDjM62NIeMvMLc
IDPDWcKS3qnhhfU1IqRlLlEFhxnfoOPQBkdaKnBrxpz86E2k43u4KdqsF6MH
/Xf9Uc1ZL+LZAjLAgt3jDKC4Ph88Xxn5rKOMwZjZRxIL6NPPlf69lyxlIzRe
yfEtMwQP0IQdUERHuQhwWE4ipwPk9YdtqGKm293i8K2orLQml1L3RtTGVXoL
eCmZubTifMFLsXG9KhppPdruMB8Az4zdMSpjZdtFuo2PAIwqeNMSRAFQnNQ+
olisIUODQkZG+pKAKOLZO1GHCmv0d/rqOPXbJppPGqJtOO1b2AS7D9ZVrmoT
Q5vxQY9XPKxTWon02gQilOMPNRlqj/gd2KmCpzJqdh2Z6hzS2nFi6yAJgXcy
NbXVmlyk51cIvEWvVtTbd9iHCn/3enSdi27N63TNkKUFU0Dcwb/k8Eg+hO4a
QNzfyhtLXSAD9xCyji8fgnqUMuFj3xw+vCR0QCO5YXoDIbJFPEhD25lXgyhO
Q9e6QC5sUhp3pFB0YhSj7gVGRlw8dXQd4BIq3jPU/0DqebJCoySVwyqvm1az
EM2LDzaGz7VfqgaGdz5utZoLd9COu/Ul/UOyOF9MPsB4wgcjIplC2UtRvvM2
9wV1T9ZmzOKdBEje1E4cDWvkHdtbAWqiArQq/dlme1NY6n2DcBbTwDN1za8n
YFOmOSRtPU0K+WGcj9nCuV4QmOo/Wxo2vFFOD4bl9sTig8A1YLaPcjKDFoZn
Y6DXvS/PDwPT5GNIka/bGNsOvWsv6gysx3CkgZCrxFnzXHYH9MdCIBybmB0t
W9wSd7yqWFmTgDpaQg3MOyJ0Fd59YV8910yeLScID3NRqXXeJ7ELx3lHN0+J
uMXZPr9pBbp2Q9IRbK5QyATCjXTRL2OrGggVEukBTlJQeKrSvLuPlovJBrsy
l+yelq1X7YdZ6zsaAXUlcfZPHnx0oAS+aRpwJ8i+ORlkz7vJ2zvgIHzX1LU2
lEsNiPnfUSX/n7Oj/d7cW+R6OtxqbSa7PMRLCowrimwlMxDENyBgyyVUbRuq
+WsKteiFvg6/kVuK9YKQ9MTLo0e/x31Smidab190kHB7Fu9/o9YKFN0v5ita
i3fD8l8sQwaOA1ZkVViJmWwYx/kM+rPWHd10TeT70VTnhHSFChBmz/kbkAbN
YwLtuo+JHAk85BggOS2tNhKlhSYdXVoRXb8qRMrzRkPfWVSNlP/La8fsXPBW
32dPlXphy4JJg210ulHajYu6968y+nVaWepLIYg2UNTHt/wAp/Z67V6eG7/0
nAW5A1YFtTwtELbHkFjHaKLqErX0Eymmc1i1O2KDwqHQ2ygk4eW8qhhTnlb/
4cxeNODpALreX9XjnzM2wDUzyn8tqJ2i88vO5oDtFdGAv6WTbG+DfYN2M+5r
MolXAHD9LI2j1ZDvaDSOLQvzL0p1hxG/Mv/zQaPA2am27mYnik1hx47UGGuo
c0fjuXeUT3F5OjBosveA1X/LvOCr5pnzOBJ1wkWqsSo/4h/WurBrgXmbHuqO
q0pH2AL8D7wjbFpEQnhfX4EY1js6tqQm16PfzMXB8U/Nj3KuxPYnwcEUp31+
ZBIbxhF3zoFqwo2EUk9M3EVlNzsZqZjX0TgKM5tbjiqiOHyrbbF2elzFl/J/
QiZ6oNJ2Fc+leI9CPsnA+mwDY6LGW4VspdJbP2+Cu/T4X5uHFwOzbqUzxE4T
uTPw6lgJb0EVkBlAaejcmnuLfZxS9oCYiyof1Up1Fdt0tOEQrTh2yIS4S9BM
876t+myYqN/t8u5Gb1OaLPaxUd4j84MN/GGR0HvPW8u1HvtwIx/ei9Zl2nat
egNo4h3KLMd9AYlJ2othMu6fw7O+ygDbIsc0h9gwXsvKx4hl90OiBfD5w/5f
6p2Y+kuVFXGQAQlX0YJzXktYm7oeZ5lu+CD4HjCc5RDHxAeiFpFLl+mlFJTw
C8C8VOoRkMPqAkRUmiuAKitVerv57RSLhUnjGDOeshwTXZJIqBW+2XP8Zia4
zqsJNqttoO/m91yrgxGw4MVcarihUA47sLE3/lFcJBKkOQvdgpYA0P8jaYml
CIB0LXumVnKPBEyR6yH6h6R/Lcn8BlaZLRyaCS2INzgGMnHP1RgVKP+V4NDE
gfWlIfll3ABkiw9EuIko96muBIcTM/7X2rZ6YIrwpHtqDkudOPWAWHxxqcB5
1reldzf0i91+s28AR0afkskhggt9aFVkIcYMYRH+mtXG2qf4IpEJPyp9X4Qr
tD3ebqjfDLFKfBVgDB3CkvK6otAnQ+aY1KOintep5Vm+f9JbM2jRD58Ee/Uz
eOq1wdFcp7YeSRh8dpqNt83mvLYBTQwP8Fgd5wNupgwVOC903Ouk5r3sXaW1
CMeNBQNnmo31cnToYJyalMiYfaV+iGIYyIi9MbiGl9QglJciLg0QADarKq9I
uLDPjOUDC8WGDdq0n1/miFLTGDkJAUg/5Dx3TMPCqDb6R5RqPQAUH7Leztb5
vZh/aaCxhKLu8VYVXS20GyWZ7b0jnMolSsjbiysxgk/ERXeGDxNRtcSXmpSJ
p2rHrSCjdAwGWlGNrS9A4/rX0exOqfLYUL6LTjKRPrTkBFGHiWL56FpfdNia
Il9jP9gs4utFfNZgFCMGYGWs1pYJ73iKaBPzKbpPFZ/fCx6vIRpxwOim7+2D
QVCSeSgLQlkAm/cT8VwtBKcNTw4Yv7PG0TlUQZY+7FRV5ER3/KsDQLZ2nY/Y
+bsMRFTqnwILhRzkEeyPjLeKfOkj13pVCGlrFHexOtZe+w8nOdzxap1q8JFE
WoHLZo+OJWcJG+R9WCrYlM3LO51gfp+1VLGU2c/uvEFXYZrpgN4tANdvOjdd
eyje6E5FHDBKpj49FxNkPPzOQAAL52ufwAmkvSrRj9INVWdJ6TKR7Uu6gXoT
K8mY9XyPIdRlv2ORJ6Nm+0BtHYzbW1kMUPgtntu6Ze7lVMgLuBr6d7+HTatI
qJXXT+t8tqdDt16i5+jGA6h2ZkFIsBKBPyatcWJ9ci7AG/lyZSRfGExHgRgg
kStUboiTiA/OsIdx5/Jn46smrL0vGiyf07dRl5viUBcvi+hB71djUr4DWlP6
/mRMkh56dGGxb8mcdpV/oax0xq5Ee7LnBIGsgWCDuRUAcZx+TfC6y24Za/kU
75p3b3RfcBBLN1v0RT+XxXzcxjTMp6crr0oG7cZ6p4jvcfk8vdGBP4woQRkO
4TTGTOgvKRathDwMTrsQkc6+lg7lGvTwCbThgL1ST1GKpAYvXDs1umjE6MJf
nDo8TYcTSNaIgmno2iJvzds1uPI2DsYCvq8ijocOkSBT2WVHSosIVNZzVnb1
kOLnagrnXocnBbZl9eQIPs6e4yUe4BEi0jTiHU2kPq2PqK+To5Qc2TK9Pxu4
byQztYQoYwJYjH2JNj2KkmEm5rnmoy68iu4mV2VoKYIO76bancV9ekrMlaU9
ZDJzHp6WlMdW//UbSVvQN/1fKUCBo00jTiWCSJfK+R+Q22XbLSM0hwzL/3xL
RgLE7/9tk+VI3lLhYfBBnRId2tj5bTucKG9ym7Hh5+vLz0DWkpdx7bPx5ikQ
KHEobUquSSj3zJI/FeaGN5ckOadyn9DDMF2sKw3EBdRYtRNVZdnxKiEWdLIn
mDC6xdD9cyxxx1eS6wtCAWYzoFjOeHiBJc5K8sEZwnELRyA7BgBlx8WCTPqN
FeScn5zLrqnKIhQyWYT0eyNws5wHTbgRjh1ufuXSEjR6rnDXUHUGJYQRx0V1
K5p2bKuMCrcGfZIFtAOqJjWQatmFTr1uTyuDvMKgOzUpNamIZj0iVq+vc6i+
WMQmRjVBYEcakqRF2dJqqzhrM+HstDYiCsPC6eP9JsGYOLjexYQt8DpJcNgK
ff6DMs3e3Oq6qGoQIT9MeFKHZysNIr482SDzsPsjHYZcy/yp+XkoY7BEav8d
A1zSknsF3HJafRszWD5pU8SO43BlaCEOWBjRSxfEGA3Bk0ZApKAxIedYmcpQ
nS2g+T5e3Dep0r5CyX9admU/VUxlVZM/2xp/ZB2C4R4E1JA4IxnBtX/AHXOc
rV/ayUatSMNtLx+04Dj8yHHg6PDTn0Nf/LgI/IsjDcVf6KTqsGx8iS8YxHST
mqViMeGloGTTVMTp4LyRraY5eiNqX5H3vWuIduNyCEOCr8K1j1vagTWlLjT/
vnrx5PT6F+qMWOUQaKllAvm78MNXfgOKHzzuh19W3XNewGXBTjEfjRRoT8BR
glre4JUf5b7QBaIm2RNhjJQxNMUp6HjLQjv82cxrEupY8d2ZJU4dViXeCnvn
5zkX/wEX+9A+Vxz8uu7Xhx+Xo481+Y3fzjYIeu0F5xfaX7OnvFj65fLGnqmf
i1a7MagRrlAy8EwIdyFZw86Fggw/c64TRmaR9DARjApB4pWz5sEJmd1nDzGk
/zwfbZ+gZD45YK6M8YnEKg+gBg4TBmK3Mltt986MHcGRGAtsZDh2LoQyaSOM
lSNbLZeT611rEzlmjrvIoWFi0Li1uO2+y5dZg9NaSR6xUh2nLDmCgmKsVXPr
L1KGZvKfaUCiWHvZzhJM1/SH4IUHzacaeeJRgPz9wwNbs/JZK9m59NYXrjp9
938u8F7i0oF2NwXhTJdLhKVnmTtAhvRx+pz/kMGtEF6S35+/7LRkuT/Xnhh+
dfeOb3aV2pKsPEht6J//7Yxa7Yq31rbeJVY+qn/2Tw3GQHc92K/e2aRmm7ZJ
qulosvxw5AL+MDJnY7nc1uF1Og0vwDWP/LaZ0NzVEuF9QmOwQ3tUi+NoFHD/
jtoRCX3xPnEf6w/ulAtBZ7VgQY5P+J3Ymn5qZWpHcoJKxHgDjUUDrxgQ3wKs
RzkrL3Wj+P5Y3A7eDavORrWy7KCEzRrpaFteoa2PpIFlyRYTbd52lrmSlT7o
rsMUmDmKdLUKHRb/hrtC10WSlUZuSgXxS2F4uUliz3ZBe+0krvPhlLnl+559
/ihSZUdUz0ECN+9bMTlDLqFb1AkAwZEQ9RC44BM8bTLeLSAIPhWa5YN7UfvW
V4ZYf5UTQgEmyDV/apRtSTjQToLqzDXhxqEjtcS++x/igxEZpLprlp5IsWek
xAUH7XhlIX9thTxOpuMHz06GFqLqZpENAf2hmkkAWQUmr0Ofw5EmmQ5yolP/
5LfO/KN+gid4d0KU+xXzdI8bY9KKOR5QevUniXUhESTpTBhL2kw7MS8Qh9gE
F6sAucg0zKqTQPBrrT+XlUQC5mBZqODsPJuZuLgoavtWZOM/mlHhaXvY6F85
SX4voGqKlVq0yOdteufZVCCHc+O90Q3Moei0gX3qyLoIu9wAuSUUuzNtY9Jx
GHSfN5iXBGvdlr0gTYhtti/kRVEwtPgSprK6aYefbAZhmHpWYwUtlTnZnjfu
fj6zd3Ler5ewjx8IiPZzwfMu1HVIYvu5Vr/DZFUNA0QgduS3oumsKOFhVJLM
USixksFrZN9QxqKWxv64nb+hFe+OePh+dc+5lCxDRPXilBGC7Xw/OGycfx0+
kfnopIYIgaWrjbbVs3Ms+SimUeVv/bB+DYR+/YxYI6+PNtCha4jKAhEncY5E
DkDtos0/Ugi3YiQhl46CmVXZXu2yxI1p88KAwwxl/+nFZCZLYjRWdBePfCfS
RcBI/Lv42rQB5imtnIJrgTaJQRIoBeNsx3T7zOw29XRguvI2U52gLHEA77Dw
NilKJ2XmXwUKBxo05uVxWqTI9rYYu6wTCoyvK0Iet77f/Y0U9P8yL09/rWOm
Rl/kRu2/Kw5L/0f244/6qPzU0vWo0codjhaQsBz2B9rTgqSVQRiEt1H7ECzi
KLTs56xbAQrY26W3AhmmK/F6e6y3XZ+AFWNXaGTKDRSOWRPQjFU12EH2wAy7
4jD+dcRf59ArFY4IqWBoOsJ6Mjv4AQISZTynSm0Nw9iazf7zf6LtIcPDcSs0
RnD2fjOxnujHwrQcsl9cn1A93uwQsL6p8uPvqt/HN7997VozyIfluAxMKe4Q
SD7fyvZuIKgidA+RLzsA2eHFSiraFvQWytRrrhMKV7iXphhg/9PPj6ohR2pl
GE8+Sr+fKa3H1i5/9AwPzrXSQ1/slOtM/yKX99bqCVFDh2nmueQVKFw86/AT
R9kHljTnlmQCrhVxHX99ibCP/wDwwpjL43PKXkve8Nudkns02eXd3o325ihg
4apxKCf9FwrokqdP+wfjtzqVlo9Q71zDywSuPuRvaDAfXDgBR0GGJLXwP+3U
ApcGW+yIw1mNPYh/Uj43bchaNcv2GEaEHyY3H2QiQ3lmwQFILVtuquavZ9Wq
8AxkD5EoOD3ZR4+hfhjUDHDt0hpO4YpNxbPrtwY/2jK7BZ0eflfBezMwiE5x
rSLZ85r6Mc4YgAciBSTjJnkHyvHrCijPqlNSHanSe0IAggHOh1KjhomNwdHp
QZpGSjeye5NoVoZqBYX9BND/y0ErrayFjDNWvXvl+Ruu5gteAc9UHGpdfEdl
4hXkL4B6E0OicadqwfpRLek3+ly7gmwJkTkcZVQAT4mPZn10cXYTsepjAZx6
33IwdgCpFaWG2XtfEq/KLOHCpV+jtK5WY/zv3bzXvIeMAFI61zYupnYbizf9
at8FGV7vlnL2Xl9/Ko9METnrtUs2dqaJahNdMLDeRrTtGGAcg0+IuTfD6nmt
/8Bc6TR9dm/ccthw0S/6SQzClCT7mGVybqz35trOmdr/yKjXpK6n5F3EB6xB
WidGdQ67geSpbuUZW8D8K3OyTTeQrlo9lxgaY24tBJuLRkwB1g+7v37E3phO
L1VcrD/f8F/xEuWWR1xONxPSWUb7yFKsF60sI8RGQNEVtNNlPTGB2SrjtfqG
rsjdQG9koU84NpNd8zOQ27otpMJ0IGCsl/6gcV7CdaN8BVhqJJ2dqdOQo/Sf
rQBWPvcFwcAIwkHQrKLi8r4Gpwgz8iN0kb0G4pw2ODfNfsSOGusq0hU5C557
E6zdlCIXvfSWllXKQGiPRRlTgHMyAqmhdJuNq+Za3FLnu2miXGeT3cizqWEP
N92NTkV0OtTxgLwn72MDGENTaXQseFuiZuiZXF1eNAu+TcabBChv5qmOMZt5
buIQ5nvRdJsJimceeOGwN6M6XeKM4dZ2J/srTYyA8xO2Fq/wzUj4IzNDx0pY
OWsOQt8GsGZwJWLHtnpduTYZyXUtsLHFOGVwSfbLhj/YPTHrhrJScWiFXZfu
d0aHaPLLoG6tYqaki6Kfx6izv1utx7aEEB3rJlVCbgjMtr/qYCSC7SH6/3gA
66kqOaUxaK4y7SZ8IbQe9b5wrGXDlDnkBvOFHEZtV6pg0jhzvLGrEffRkGdN
ZCPg34EpZ3fIEGj8J+WcskKacq4Fgwx6X7nOWTDeA69ZSsfIVKM5uK/3cAgd
bTghiocglrcHa6gJDQDtTfkqkieU5TrzpqPZYDc5KN4X1PuneWO/R9JD7KQV
nWBPAJzTe/DpU48CQj4mJw6bTF+kvvP9MH+k7Jl9IvMd39K3UGeuR/TV/3SF
SFcj7NRp6L4vL55smfRJcEfRdT1bw1FA8A1QJ4a/LITvEOfhLHC8VTU6U1NL
U+WHJKec5a/zhm4dK+xREonDCzDbl0Ryu7q3VpuhPAnbu22ObBJjVenpW+eh
cmGbTDRCsqvUb3IIbo1Ww/0YWKsM+SpD8Q8ZkXPLhygez1oS+wVuAn2FkJvm
Es6ot8ZpxMjtYsazgy7derRnuerhBT58dG2OAYbO6BK6AvcwDicSQioiMAZu
OhCnnZ9w0C+69l6+7M9SStXBL4SHrywrgtNRt+AtxkHfEBCG9X7K4O4GT3ZH
1u+/daoYd/YmwBsPCXtzX8/EKnZ1LnYbKf8Z2whPGjl2Bq/cD37jYpqhxq4G
9ghhwu9ZN8TNd6fNioHdjr4GwWoO1yzzG/jNKSKjos2RxSpLFi/jK+rwt5JT
hnzaKX/TFgRyNnUuJUsxl/Q1MrrjcFtvaV3Y7cvHXwcvZqYuYKhx3sA/pz79
+ueqCeGLrMm3/IApQqfCQ/kDBVZvZtyPC1c+fPxTOXqXoLH9MY5Q4lsIerSw
bKBQQoNAANaNr9zcrCXrmTJpNdb7UlfjBB8s60xYJAenDAoVJM/OLQ151BK0
n8T/O4LSyeu/d5BCm7GlcOqvw+oDMBWZw8+DVtoM+YxrXmY0tBdD+izyHhRc
9dGuLzszmsEB23uOK/OddtWJlVSeh1u277VW/nOmTwpp+7lUWnCaermioUM7
YKYDIo5jn1QSkTs7eR/wqOWTo+RQ7wfTv1sO0BNSqS8QixW1uywCruZ0mltp
3IH5jsckpzAIPqXZyaN3e6nWRyxghvjuoX5CJQIEMpxiqsI33oqhb6GXRkC2
RgtktK+YTK86skxkXpfilyKre2Nbnoha90bwd+V58kYcLaN7Qz2vcy7eWjHL
E0pnWrr6/3GR/eDQBNXHnxcXUiMetfgO/yzdkleg5wncn42JPOTKfdl5nSjH
A7kUdtOUa0Z4ymW8PVH1/GeUdPNsS5ZJaEAywjpsbWmYsFiEgRQP+4mp0e0D
4ZS0ZckK8j77UknPv915YYIVvvhVlRRVsZag1GjE62KG++cnHIoWnsYhL5U9
hHXLdQk6ZctRqrQROoPGRN49nbP7cfU4sWIEzKkGsARi1Cweo0InKUA2Mrm8
kCylO0Jajfonh1Za7oUSJ0LpewVWvTgtoNOX7+U/CeaSqeAJ4n2Qp7iMDnHl
8e3GRoZhcPEosVN+dJtHMrAg0pNz6WWm96y6N6Cu6eA0NQMX4pBre/iaMAQA
nQo5jcggTIvUDS0se8hzV0QjJnO+iYXmLu48xQPlz1Wwu/5lpJSrsbK70/uJ
8DqeigXYiZ74LOWC+p820RfTgzV1S3hZwAVjnmwi/nuWE7MZzxDg9F2i3s/H
QiHNh0KDp3sIem+l3NM=

`pragma protect end_protected
