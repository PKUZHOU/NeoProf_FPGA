// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
tukOy0iwhRcvqGhI/PBhGxGPOCWq6tVsnVQtImdvXYFbds3NewdFjH0QOC5V
BPUbaMZKH54wpK7iej7JcaY4evT5nhZUTNUPsreBYhQR2vpUSQyheLXk2o9v
R0XXu3FxeCI+CTLikgQWHj5yp2vjsrYX8cv4A5xuRdeLpJbwsl4DMN46OIkH
5ljJce3TmOtYaWsx2dH1LHqt4Ag5QdBbCbVQ6JLEIc2PboRGKfDNgWrmDZAf
LBHf3y+tn5cr5bFQcOJnxoKFSJ0DOIE0Im3uJiTVXQXwVUv4V1bTzFbkoAE6
BSh7TAVTYHO/E9oFojOYJwJW9z2uf2NAAcpZrIC9kQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
L1LRwQibXD7w/AAGJeMqAVLTFaWi/Fa8QsF3X5F7TIfnAUQZrAgTvvpOD7zz
mZ7wP5qJu0/CN8r+JJsjgFN/03hAxBR7snN4RIajBVq0SFIIbvwWPZkSAFBo
xvMMa7rAAH8uHNW9PzzFMdw0BtCAtia2hFTtG/eleXuOs5QeRWbQUOzLXbVp
mp7ZTt8xupGU0ZFVg8/SxB4SK+xsZNq7Wx2p+ZXVwsShY6s88n83/Z0Cx23W
fBAfPfanBRkhIGk4riPYWDGwtuMpzljcNj/lkEtnYVDrF8MnqPXISg2g6FIL
Xqi7eruTsaQ/YQIiojODjANgjvxcaACrkXAdi3wzRA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
AV+Uy7m8imMAcD41AbaNxVAc5ZqqftlIihtEnea0Hg0GdIdTWwpysHGwPMTt
unI2gQDou5Eg6IA+N+YLGndKFZO/z6nW0GdQZ0KHcMfORUkCeql/QluCI5ew
10yAvHpblqfBEcRQTXaxLUuuGMbFF24imP/4dlyP/T6W86jXsKULl2Z1ryeM
z93spIr0na2l4AatNWFEBEkb6PLPL4/hIYfTWzut74eJ39zJknSdOMnOd51q
UbDTc59KVcs0+G/ErGZ+woC79bTYIC/S35BSRQLKV6ZR1B5mchzFWPqsXQ4N
WuV9fDHGqP6KCWmzTQwIvOIIbxZVMPwE+ZyV84AyDg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
cThc5OGaGDVHaDvFCCdvVMsRs9cBkEgUwIOT6ovawrl48YVGwf5yb0kos8Qc
1VKZnc75jsSsnJnM+/0/v5Oai7TgqTYZW9ZigIc4Ay9FjwAld+jOxd5r0soT
SawJtVcD50LX79oMLyhzRUZoUDlMmTlSKx5iFxnwuk5HuOnstJo=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
u5m9mwf7974QgG/iW2/z4hdG2t5HkdenVKgaDYCKBpIV2cSS/pw7IPT37zkn
pti5X5phMIXRuqftfzw+5qSuDfNQA2dol7s+76j0rLea1qZS71MmNILzV/SH
DhewL2cEDZ6UD6aSCyDcHyghKZnDtJxaXabtMg2kDIv3T3JXG2iXiq6ubM6v
VIerCoqlGq1nebO0rj0ORTUNQCu+WbYtIVjfRdrhDEMY8xOesVsqV7mpOYdb
zxE4PYMIAaUFDAQvGIzrF+emhw4tYQ3BCQR4l15f6mfpdE/iiI8Ab+uRS4WO
MCbCQZKnxecBb/5WyW0r4fbWCYZ9Ycptb4qy4p9k6QNnZUDqv707Iw+Vwi+B
aLcNX69VF+fVsKqFzy1rbqqu1yeEDgz25KFf/9OQ2OYDAmcmyxs5QQLtMMOx
eKpI/NFZlqbR5/x91G67ZVGJAQs4wJxI17WtKjM9la12zR3Ibt78aLBkcen7
EVDfKYEH3sQjZRGfiSWfMC5qMIUHtxIm


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
JZLmH883uwWRg1KNefJtp3T/iUBSjzc/5GkAMZauIDNvQbppQ6RByuD3nRLh
XwDMUdex2c6mn7f1pDGrB9bd7+2+Czg+3Yj95OQ6vnmH65NlrNXdD7VDY4ia
Z56kzfUO+0wksTrJ6v216XPjnLu/NNSY4YZnV6W5bgiUd/aGHgg=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
okGilfumKQ8vrJtWJ8RSVi1XwZ2+sZkQn2sp/2FUrdkbdg+1gxE2V44MyQPs
4D7Km2T3BE7o9M7Gh2CgrJzZi2R/WPcBx5hhCw6X2T2+ceyP8gccjhe344/Q
um5CiYxY41bYE5CbQny/V0RrQTfFantWH+4DYdXzWT+WpR797xY=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 12512)
`pragma protect data_block
i3I7pqskq1iY6QKVDVxEUgOnsPvAXDIDV6n38X1fuzSk1vLfWVat3V+QH8yV
dIOFS7T4+lpPU/Bzem0mIP/FNgWxL+85ktQw2L/J/17F0cUgJrPAoz32SI48
+Nda2hV4rVKQnF2jX72PFrXa2XGQ64EdkILxFaB/IbGq7NSKACpAR1OfY0+X
EC/KaQW5Heiw6u64HpTNJCYmT/189Cl+9r2FWmyJqMqvOMCrXyAZI9WyK6gd
K5r4CpkzHYENE6tOWrkKtdfPT9aqRTZdcRp3Bv6MvcNEgHfBglQl9GK1p2Dn
iQx6IjFZR2mPBEZecV5f2/3thr/dsB0w1ZaYnqfdbBpGKJczQdVsThdCSYyC
805Ry+3IaovpPi8p8PjD+XCivBv3D4Tq0828w5ec9+1SJvnRPn8ObIObIX4r
8D1h4iD2l7H/+hWT9P1LIkyZtqCbUapo4Ngc1HvwG8zAoSw+/jZZ0WLuOi6n
iLDs4LLSN2GZd34/VY7uZ9VRC3I8G1BmGUuRW9Re8RO5Hi0MdGxM6G+XXJTQ
6bFsN5Hs9rpuvamg4ESXRA5/0BCIm2GR1JWKrEfiF2C6Ay6Vr0vKO4z7171S
LpQUpePKKJLIJwemvEwfR7tb73fV/W7r0MXgXOyUfDxObxu99HqpToW5cC/p
fuuOZazFqxeKusSuIhx0ikFNekEDu1ZJUL5OKCshbDD018urIak79GNr3F2p
7H+Lwx5f+lkharxitlaiLfuiEw5VMCT9scLAOnl5uTxx80rbhwHwQTZ8Zpql
b92NxeGFBKkZwSjzEjAo46iILTJzO/Ktg+puJ8oSqNshqlrE7R2QpYBHxQ2k
5npn1MCvmr2nWJWyssuBw6ahVbdgMmG7UKD4zs1+4MJHgQ5B5UK/dQy9xHDM
PnURnajtqEOMf1cM4OsnwMfSgcZJNbEyQyec2iyiqZRb5pzc9o8oKe2qI6QM
6rGCDIeoGEF+qs8yjWZbK/Uc4ZGZ3kiDQz5/Mj/ZXdh5Zm6QsykoTqVtv/Dq
eFrwzKXQMqPJEu795YwvA+pJfHkiR3JGLTyv5tUp57t3q9Ugp223aRRaCB15
qhgFLYXDmOHTQO0HprTkcqxqjlFz0S82IuhMG2nY2sr7/GHH2MBqev+FwzXE
QSPbiG/dRT9VcZ9+SqESY0/zJmBMIRRq38NRLfoOWMNyzwBaS9rBWnPMIvJe
GVuTMwuW3EM1cOf5ZWzwdv6LaQySlQNx9kLyBoPuhj5O2jMayOq7COO0ySrM
RXztnCcWWknh4KoXPRlzwPvNnOgtgexGgImYrjfruh5Po+hASbALIlJ39id8
ylt+WBl1asLeQqvcOPKnE94moqKiQqZ8ZoyU5RCwuCjzGVZFm1oHoseF5uvy
ZeGm8o1HMzHzIauDicYUJyTmKy4lvYvFDU3ZiCCXdWh2soosYNNwwcVBTiav
e19DIGX/f+m303032gQY8a5e1DRTR/Lq10zE/BFJin/1cIHFEjx7pCIkVPrU
AIvF2/Tyhlw5kF0maV7pp2KWK+LFH2gCO3jk3E0hY0qF5uXjuiSGRsGNo0SP
qoR/VsCMe4NTgZNG3s+cXtLWDgDHUHszai2ZjXM4XON/1ENV96n4rrSJ+XmX
C+bA7RtNRum+Mv7lBrCZZZNtS9tm8iGD+9ars6sUFZkxq2QMriMCpoIpODYu
qA3ntDEkDzuUGqjJjuCPbqAaNoNUFlSn0xf6DXAhyvq9a7aAk/rO7VFIHjqC
6GTyz8aV9Rn8xhaNdJjuQPVIDhLGKDK47UPShStq4vewjpUj5v79VDoFqBs1
gLJAFKXqX+Sz7qDiezBgRJ43EDVkQ2+d/xX99v1iLlY2EezFm/hGvyf0bsFT
XhehJS+Vw/R5Jp6CoiOJDjwje+bHe58aY8qXE0Pu81KicuRAJb/CxKaiW19e
itbhEJIT3s/l6YIGlSTgH5npHDujgyMEvqbaC80XOMI6m22rRkdrt1A6dZ+N
5xWZMl5Gt3vXnPeANRGV1S99t6MKlTe0XlAMLYGUduDMCwJu0Dk62C5jgfFY
dkZVL/3DR98G6vb+rcTfAFqmYDauyOtxAnrGEtrrOIsrEKtY81zjgnigoJtL
p8rmTFi2KN9k0xdN5ZslBtjzLNCkw6kQ77T0s81esKCSqo4sSWYufobRNk9R
pmJtt5Olk7GVDeOEQ67qqhPJDWdXp9qZZL2jZGwU0L4vsLh4dCbECoJSOwMF
osH2KD3S+eMua1S8YIgPycBO5L4pd5W0uFD4AFERzhSp3tO6eKoPRZ6qrtop
QDOLa5y/T4yMRq61Dp/civ5AmTsTM5H23sVEyrou1eEo56o6V+VQGFpm/iLO
W3hfbL3swYBdKj2PXWso57gm3iYuT5OGFiCjHsdk4G90Jc0IYY+QftCvQdcA
Tx1dIWLOwGX/oixsWHLnaGwGCe2X9PPjo2yl5IW/hmZg7TqJeTg/tkMQshJe
c0X892TuWMk11p6GISzuDFORyN4YGOzp1c9fumj8agf7ybBVeul7iHC9bgHq
fq7rM290gku5LlvF7RkuPrBdVhcq1hxCTJrFTPeRDcIOiyFBpMLncDvvzK2l
FqkjaOHlCiZjzrEdilt6YFcKhUzL7odPFHNwBXuwMUE+E2SSwvzFTRkka/qq
uvLmQHuXsIBw/gnoxJ4V6896h25kLe2V7xxnMWg7nmZ0bYI05hisShJyBTlZ
nCyltkwzlbKc4k0vSe/8zDaug8/TDFGcgWVuE6KMAi4cM/qUAplLptvsRM1J
2nBh/pEpHdSfCikHVxqk8pMoPFEMrUfUTlKEw6E1Uos4krFA6wXTC7O383dx
dPagxmRZKZxPl3GVShhPdcW7uFfPbZIKejR35HhdbMPfv3GWJFC0rlwrZCAs
bhMVGX4p/cnXXQSl7yYsfODaton5JrC/uE52DYhF6gsU07R/+c5nRw+zkVCr
4cwQTu2NwRxvttygyrr34RviPvt73Rs9zmP3LVrfLHPUIf+2M27da0U4yg5A
sFpbsTy1lsk2+trUwEuHhYZSwz8wvalmt/NsR5InKzcAJilf5GCP+my986FX
ojnxl/qEWAnfoCYhVyromTeKzzgUvkvpn6/Ofl35ajUqK6dMFeYMWHwBrIoi
odA+jBrT2y59M4bb2jvMbq+bO6zCfxvM9qyXuHJvavlR+jDV/Pfj3x35NpqP
fCcaEkOfTdwY0B0+y7qZqaJY5sstCgZqQiuUAmHsx+8qvCRpnaAcz4bUrx4r
C2JgmP3gx7loK87kX1vMyOY6EOuMxKf8qv6YPjOF8eAHa5Wt7NL6U04a5AHY
NCAhuSIpwmWwrnREqNhoKR5HDwvbbRPLxHRw4S3paD+kKMrdDVON4B227PsZ
i+XuPolGY8XSk9p9fK9TIiHkYsQBINVRjzpEfV1gnD9LTJkuF5k0Hq6FT1SO
5+DC2bsHMJ4zLTu9diWb8AX0XYHB4WQZ7xqIZrrDt1/oQdupFYKlXptb/0pp
XYHNgMqemHa4c061WFa2EmasJxmi6GAp6+B+E0rgb+Vlc4Vq/6QRgzDOP1ud
unjO7unWdL4bBAnMKpJ9J4cwhIcj/gVRNCSjrjl22W1bow93z2KQIzV4wh3l
626+urUJe84JRoTADqOzhlwkwev+3Iq55Hf/J+Zsy6+VYqbhLHcTdffehK81
TBqH/PG9b8Aag8jf0u6bpoeJBpvK3zMtlgH+zYiEogtsB3Ofm2eEQYRgqlLS
zcoem7G0rGKiGXF1d5aCqjMqTj9YDBifTHR8Ln3A2GFJPrCL+ESGKejZnmtG
tRq8knYG+jcusO5j1e30+YHOsWAhX8AGRt45s/cspDbGqvhlOJXXnjv4m0BS
K72vzXOUvBVb/EQ8q9Yoy1oGqKjUDhVxN67yDeIASSuer251CtLrOXjlkbGv
oeS8ddDc+FUP7rdVD41tsDKoz/3y3PP6RrrvqgX81HYCpRUe7Tcl/K4kLagz
cy0E4jUWVZYlSop8SrmyP8/6ETcOLgoeX2uW+GydWsex3riwtIQrHuuBaKOA
HQIE2Unj+bOv1ZIuLTVAgx47NOwu8HIiLd6QUkTa3uPW6YC6XdX1s3ZZeIIt
P/6mD7qOkX5h3ECTakhz4iNZ9I1dZknRpA8n5EaLnlgE3xP8MgWtcHWbLdX/
l+wXqnz2+LtlmosvFmfpm4UPhg0/jJpuBTT2ONoJrizX9kt1uXH+8iwfkokF
6zBTEK50uKENLep6pmtbaMi5dCSnidQgwiJl3OQisrh191HWoAo9GEDPDWIb
wZ7ryBLYAvP1SU8sVe6BtNw7NDNbU5WtOVTSEPzWDgUKk0fNFPTSWNkm3IXZ
XK85Io6AJRA1ruphGwoHFl9J73PPOtH70qnEJUJg/v6SzhD7Ey8eLHZxCPFG
74K0n5wMXPQYCR+ThugA4qqMSRj2UHoyz0XL3cLNla9xz7OpICHj91ICBXPv
plkRRTc5RPTCZMlr3ZRlxas4a1W98XqB5Wb4b/LCqKCVry68PhfYqzEb6QSD
0ZbNf6kccbeEAzYTR2FcaDeawLnv8n5r10LG1LtjB9AAqoLsd775Z5bYsEi0
uXATSXVSTVpdIFcV/c9LcXUkFAWLobb1JSYeOpPIxWTFHOJ3PpG3wVoGPmOB
3knKr60amPQYHa2s1AJP9w3G9VXJlcqdaEap/ylSZP7+eUwO38BX0pbe4lDp
KryUKgeIa4zf3ZpNdQfL4D5jbThB1P3UsHMcE63gjHWbKDmPvIFZ9NbB5P47
DRQGxsfd2UcVgZiMRGUra2E91l+TTUnqm6VytKl+oc4Hl5HfAOeZjeLY1Gbh
QKY+DLHleLC9rKJZRH5vcM7/wzxdh0uPFjmfu3ecfXQ4PGWAyDbbtjCMkFFH
563VqPOLSqCAzAVDK5OrQVlLaPVODGAlZp3pmqpOSsTq9MpHrPlL1XCflm1n
CqWsFl2Hf6kmdAT9EiTAMDUt1ZFUj2qgHEYjQ/87umtB2OzRlbACvS+sEP7r
4uDMwuNhAMhkzhyuT8ysMkhWQ/jEml3z90ExEvKQBuLmlksfBoAXDliuXFt5
Wt4Q1+K42kj0qd0mlZQqRk+OYNOaN3gdGurxQROnOk4da0ai3dxwHkBS4/Vk
hM1oSRepHFFxaj2WuZzim322GxubuSOuzLn3jVxgqkULFwSv/jqTUmUv1bCX
D8b2bpAS2/flnLQrzCeFZp8IuvBTi9KVfpnsGWyidu5+yroSJ9igaqLe/ICC
qjuu6r+NjIlWCDaL0qQzvehhyolQJfG9Eb6WGaXZsXquQny+ojLeEyzyZwkZ
0nuCHb+5CgpKVbsbnQsPT0OoaDgt9L1e/uycnN6xnguZHV7IsqQ8A8O2n2rV
VQaScBghMNkDtCQ9KLgIqMi4oAsYDZ8oM/1KOctXEfHkDc+9We2mBXr/d6il
PO5EYYLWlB6ByG29Lvq8bOPL1j3KX9mhGo3OqL+LzgLU0CIRp5A0pZIJjVYZ
VZO5saOOYBc9jqiG6TlnICTmh2dAEHjwh/LSVxRN7EtWoCEeBkTaXL073jym
SUHuFrIdnF+lHpoP7dOdX+lilC/3XsVeNQQIFL4uxOYeUwyjNmWOhDK57tSj
6+yH4mg6lr+1/RfqZVqJrj8Lad3mFKRi+YnPPyee+IqyQokA/1dEEnaQ2Eeb
53cryiVlsqEQkGXdUhZHjupED8VZHhK0tfKUsRAt7Gp/GycgBhUvwp6wly43
uy3kI6fhYpwVMy74AxLn6gM+IqQ1sHPH1ZiBHwgkI12j3Er347ua7HATqwLP
CzpozRpt9dpa9PMZWkIwX73cuwf3YvJ0EMUVMdJthafgi3FBrFmF4PJlnx7+
BaV4EMoBTyIl3gaAOIuAf66imE2iShBH3Q2levIZE6vne5O5h7OiF+2E2GZK
3yEAIRWGFSZ0TFA/XYv4LrWRk7uepxuHcpzEuDftWPHq6uAplObgIEbXEYAw
xbPP1cwywGNx6F07a9p2PSRTCKcqW4xuBggBeivODuYhxCfMLgRf9REyl+FS
8q2fpRMj9mMkx9klaW2XJ6+X4wxu1oMAXq5AiT99U5tkHn5Jopz//B2cFAgj
QVCwmxiLN8ZfYhGRbSBr46l8TpzVybbIYuASC6JO0sLFl6zkzTlO79dyT/7W
vS1SN71O1ebaQVEsL8GLOxwo28Doj5nXGy1CTU2a2Lh4PKjCMKTahho6PE2Z
0gx006G47SBRcSUvfMqMwhofA4qbRqDwx+009zfqSQ+8fWNGXih3wTEF+Z4h
MW8rSI+5GG+qf9BeuAygkYPW++XcART3EAJPEBkBnFusMITFd+hWeK4sWQG/
IZSmg+hLSaUusHjKLTI/0XkTSQt92P9CPRbpJPcxFZlwnv7SMjmPYD2Dni/+
pCEEWFJ2eU0WoVpPKErXHnjiZrFZcBILg9oZbhCsMYK/LKLLkBJhEpPw/Z70
5C+5O3mlRpWQ6Id5yHNr9zyKTWW/mOLwQl7xQP4N85dUIt3OASybewv+5pEm
oBddWabqKXkJMzAEb0zXq9gs0Js0WPFrtlaf4x6sUDPNeIW9pYGHQ5n9RXou
xmbRmUa1ktbaZyzi6P7Yjg0x+CkMna4aCN6vIfqd1HlKiUwE5tKyM0+YfhkP
SHKikIhsWrRlE4/18FAgDTriquqJ6VMyRAbCaq0sUC5DaU3idGi4priXSSMB
XhNg6n72ZdPIy/B9iEJkXRn4iV91s+Zj5NqWDPqm4HXuWm3vYUEFLfmkYRVd
bRqZv9ecqAwRiRvXi4I3xBgF8JF/VpW+jV4izsm3bCZU4x+YAxdY9tQ/rPLm
tj1jOAnqg+QFW/H8CNHJHC10B3RLltw1Bxg/o8HvmZF/RRXa5YQrpqnie+zT
zLFHLKDzBYGuEgrKWSWiM05p5J3u0UGZF12nna8bNIb2ERhVGFfATE6oEAK8
VHwGF9JR9ZL06x0XMbPLYlaVQbd6AHy/Qkf8mgDOTOuzPm6BSHMyT4MV7TBT
8iCuyGS9uL8C+E/QEfG164uaGX0+Dfqsepj/wW9chulQuKTCONV+DPXP8hTT
ssQcYG3WJHaDKMtorajrmIEg70oawrA87ibb9Y7wLRVl6hXwtCnEmZgh5ZjL
x1vQunjmlr0r29YBJtDCWF9Jn0ZVXOVwI7LI1LECNyHiPBC7zixEP6svIJaq
6ogrzIbcLv1j5Gvr6W9kakP6iaCFObp2Uh6k8RDMJQR54Yf5/q+r3iOGpPuo
Cv1KK4RQdGzezfowrkKIz8G89S9vViNHr4oO8JusT7JjSdt9GGtT8RVLlqHs
j+eNmLWYHVMwFxyK05y0iErC03EvLMlN+012QPdJVkU9AD7gdj2pXGXL2s3k
2w98ilnmijpzAh8EiifzGL8ihNGYdz0cHTn1ZfCH4upfP0mn3yxOz9O2C4B9
j5BaQTet+iUm5h9/T4cisYZVZIODe48YuGWRGXt6jVolDzHr11/dI+BG73Mq
e7OtbCFybX6XTzSTK/qskakM24r4JIh5V6r/BlWnxMgpH4NyDdGbfDK1WuxZ
W9Yaneqitn6roVigU/YNAkDaJSwSovhIvfe6ZrNEoBdo9M4msk6H6d/Iyc8W
CqPqzml5Lp79vg0YkhtvOXcwvjFz7mngPMOUSJ1JT2aR2cjY5Pr4w+yITrbC
LqEVBGi2jyprcpoBHr5D5xMs/ZeJtD+pUACPzwbwQhPX1A3H2ZtzYcdNeSBo
IrbK8bOw6UV7az4zRPTkCr4oQqTAC8rXNc4THn/cqZJHnC9JkpOeSSjePpRy
p7ozGuhPNguBh/BvB7m6s0hX5DEe0A1GQQlcB5CJFMTthXwg3sEF/mzb5tzM
VWvs+0nkiw9EOWoCze2/le/SMCA4bwFfdKWemddd5EKJmxA2Hm0/melvt1WU
NsEs7vduv9nur5t1wiAu4azjdJdFhnKDhiJHpDFnHS715O2EdVh7xirrKp11
KS3RRdfVALsfkM3ku9xE2N8DYsbA5lBS7x8OHlXhy0nV8fpgvb/otnz1Wf5C
9tQVNseQkeiaqi9/WOuim6Cs9wtxPKTw6U2oxxonlg2IpauuYG4G1pqbgnQ8
D5CtM0Tg7R+kn29MHrNpGtoyAuUdZrMycP86nsb3qdOK9FiXYG1HfYe8GkDC
vV4RubshNsr+ZJdwnJsIHkP0f/MfbbyP1qHrI0DvZWviXFIH9ndoTDTjNGaK
sxk0o/kuxedNkK7mnTLLn/bt3IPwgG+wPBA8tKkg0Be3eVaJ86xau2ZyFGoy
suG1/Lz1x7mOr/5sMf60E4Ikvu4AtjOZHhDukJQvVvhvTPn0CCGbyVTSbdPd
B1W4yl6GbvHjCtylg3MA8RBaEX1msRjqumnBsxUv/DbJe++3bArFi9p1B7Sc
di9JKHIYuwkmEluiJ83XpzdzMmD2zasPdShR0+uuAVu59XXtsgWSENe9AmQL
XjJPWDqOkNiBuFUAlzSrXfto8T1J/4Hsp/udqNNsmaAPavdm00ONB3n2bQnx
3OOnbn7iu79AqRCJT/tuv3BCKuVDixBiOcZttONuwNWeO/dul/pw5MvEbR+U
/KF8Pjyc2CVVIb13aJt6MG3cley7RUkSjYWdjrjj7AEOijucN88mwd41J47D
l/MueoozLJsdww3jkdYVaekeRPPA0YA/2n3u9ErZ38gce9WkBuMgeEwobHPP
PkzAI+Ow1g27SMFKppPpXRoFb2jJnsVxuLsm5uUSaL+f8I0KdXnu6lNS/5ja
NoHOXWVatM+B8Q8yQzf1DKOkmvOVplEXI+fn3da1qjp13MxqNgmYAfOigCd4
83/TIJLWsiURuxRAn9Pz5LiOB3tsZ2VIlV22T4J/KPdyJoMMqOjpkBCtPWwM
jL4zRTS1RofcFrv+pJz6Gw2gWmKmVOsU79KruNxiBNIkaaxy/m712znKwt0N
6VjVQlekCbEK3wGIBZeVyNSmLfW1V3w+cSKY1XXFZTOOqzOEkOSXrxNB9iNn
7FJxOJ1RJ/lIV8SYK2Up3D8QBupQJ7SE6kH2cc/hSGJ7Ng5iT/89fFs21CPl
EgseZfqZkSLV4hOwV3ZNKJB1iZ+xP5z28xQPGwVlCiAjQ7Ug2wlN8Rgs7ayQ
ony19l9V7/Awr3Jn3hHnMdiGO5xhJxRJ9qyY0WX5jCn3wrTHlN/haRwE1iRZ
vkT4lGjXKQf+1EL4J1i0ywS3laHuDR6Hx0nULMB3qTG5WoIHzu9mhicjnhF7
07btIRzZav+k34bg0QOnFCoOAEXaMoVwdubOLmgEZWk3v+EJXT9luZGbeZse
NoPDSEodSewWgzSehagb5vL2m+NGFfdG12rPD0+Cy1nEFctDiOpnQDvhZ46X
FEeja3jiLUd6zXL/qRiuejoSKRgnxHLMfKUkW6rTKk+bYvEpQlHPqnzxpLgX
gXElwyjq4AFxYl/qpvdz2+Wtu1hxR2hILkwhQ47/z69mCbZnKE6Z/Ki7taLF
662dHLP5snjQFG7WB1lRlv4PGN6M87Yar8uv489S7U6Tql1fltD00Gpst/OP
K+rOlRWshYmtyEgyeK3gQnWWH0b4X8DrTHF65z+h2yESXl6lIMjl6FIhQk3M
0y6PncYsO8ZgE38qiISocyoGN5KUQneDI1TrtmNj/lhaaSZHcy60uCTdTQGs
FeJCAnDoO8TFJwqNKG4a3D6lV15cuTERM8sxT7nGHweSS53J12KVujmnYjSH
+F+HohAfH72t87IMSJHdDuwcF/JzNyD79kI0J8aoZw5nopqKrvKRTTww5TYN
4r9yUVJYOvygnKSRbaUwIkCXa2GMsWHgBrP6mZN2Bct7ZLJhMP8y/nc6G649
qdZTgqAnnvFHxa14XicPidVer4t7gcJ2pOGXg8FBbxuuFob7FZjSB/S2S0oQ
eibD0oKSZWB1Zw5prDQ2l+iEy9CH+0bC0X3ABJ8fi0I/1AODOYjdhcaSt2Ac
r0tAwaMrcKZUOuS1oaMLWf7eTdL47WZRLFQMwAXQMWBeAplNvDAkhjr5eZEY
xBA+cQlJWoD0zd8cqK6fite1zauDHKYrO4GqAkdY/J7l/i9ngC8F0hBDbXXv
xVqaHLtFmC1/pIdOsGqBVEv4eAZeHCyVqaWLNejEJkYfZ7YDjtFUv2gghG4t
DP24hQXSII7Z5l0/lF20PhsqoTsU1we4lL/FeRRM4gco3v7Wr4h3x70IFY/d
RsDvhBluoHprcrgnRxm+wzTthlUxFjMB6YzZTo58wZSP6aZkis5WmO2td7pr
+P0UAMKky4eX6XGYkVnG6JmZOnfBBoSlUGWcHAETIZAjEyQeiIIZg8jsD1KI
osarlOwnBiLiFpEuG7bNjE9PTy+Dgq7neJezX4sliiw1cmt+vbSEbjkAcx2j
5RSp163F/tiDp8zfqIUZG3s5tDRUQko+VGcgwU2TUloVWRuj6Z19WXLWvPm5
/5OpK42Pbce5wVrL2CFLb9ueW3IhSdmb7fJsL2AaItkUcoFqQVBlblF8xOC0
XboZdwN7XYOKIsqbbgjc0NAlDpx6bjLkXEW5Frf+sNRab7Sy9ikYsdJM1j7V
0QPkrTd4BJKIXPbMg9St+DgNAvKb5/HNniC71NQ/fySCWw3e+iO2sBhhtu13
40FtAK0L/+m+12qnS2/3uyPTzAVV+0qNjMTDexyhFGIFY5PdGxpjjnRBJdiY
2s2JQtZ0TI7/ZhX7MV7DDBngmULt+BIVWDX3Iuzpatip4QJalJ4kCAMGTyQ6
B3axdFSlWzaJkKJajwDj0WA3HIgb1+tX5gyr9qlmul6vXhidZaQA14Uv+RZc
agph20FyjpA2GYgA7GihKI5ZxdC+MMoRoDXKvPlKDdVDtC1Gm6LTCNTJmdUq
aSMKMkSym9Z0eZ4HPASwUizuvtnKqM4ZIqDEBnIURAoD/U8C7uG/4eTWmN64
M5HTyIM4Hvtwzm4+OKEOV8h9NW9D3hlxr3ywnccYgPLltflhxwE03ih+yGoQ
zWVsA4o2z0G+uZuU1vkrRLWEry85UJ2NSNI2wK9OJFP8UlTtpHFRfXsv1TVs
2qIeCbm0pz7jtf+iAtg4dnr9D93QYSqsgzeVxBdTxMsXWJU3T/XSAYeh1kY6
tc0Ry1AGnXJujxv4OsGQ/zHagl4WUqnHJXeePIQaZRvwB5ESdNsPgQ2gD4dM
sOA6qSnNOrLCLUxmInrELLCF+VUi3nli8g06/BrFjPl8NJpsD8DIPOp6yFCU
3dGSa+NFBOzafDobWzBu34GIvClzFBBC18Ey3QqonS9qUuC9d9V/XbIfA+te
lOnxNhcemsjgp8fWlBxdt+PhQlWxR8x9YRDWlQzrXEWJYvGFK6Vxd+U/YN6h
xcIfZG1fpkAK6l5s47JfuCmQPN2m8sL7712NJPK9qp6TH909a+1TqYb3nnB6
CeHaYLGtwfXeh9Kc7tiCF/PqyjiBqwbzy5hp5uz6ADyP8gA7NY/eGDoqur53
LVG/Hh4L3CoCNrwp/VQHnnHZ3KVvivJq5SuFcbHDRnqVENVHoagGaR6O2qYv
mXL6HXROT/FzgYnEwrC1SO1StsZc8uogcsjRa4TU7PCoKMM+F0F53Af4zgBT
5UfExR7Peh9rHRAYtqQtbzAV7PuhsBJEsD9TmyvfPPt6wCVchsmrgYvOg6ET
7aOLvKt2DkRLuB4VKiLD0Va+f3Y3frO03B4ozky9dinAyvYy3jVnQQbZspa9
6gug6joODuZCbINsAQeCDkT6btGPqRv5S+vZRkX9rlAjFrMuE3UyFgv8IFxt
iom/glxhtvvTFo4MfCLS03xemEks5KhTQQofgKLZTBlnZ+NrxMhBkKqIitnK
y8vlXUO/jH+2+z/Z+7TzxFLN2ElP5D0OwRO4WhfOm14quIHaXDSwnkVFZbyV
//WEwaJHyqLdAs5pQdS2eSvmlSXdePSP96ZmGncBPV85Ge08TJ2n8sn1l597
/bVhgiFLBoT8be1aWSdwlJJ/+Aqnt75uSdD+ysXiKVTpKoqe8SZDyFjkRxC1
7Mk5MLOdWQH+vzIC0gr01Z3jS+obl3BWuo40Q5suz24ltDty1p4ExnQ0+E/9
UP/H/AylT5kgIHeJ0LhfNwcy8eKbrb63WdEjw2gRIwqeYN/Sf4Ed1/R27Fbq
Z/xlQfS9SUm2lYshUkiVquHL+G1plSeelvjRYmf7Or2dLWmNxq6HIbuOHe6r
MaSOxm3SXL9isGF3hZBPBgYCBk1LlZYjAhUCUz1siJALrJTEqfPC2FR2aTRR
wK7guyDwWu7ivXb8/OWaeWAJE5IK6DCWZ0Z8Q2dlg5Ebx0GJPOhdGhKip/hi
Hr/cnTmirqpONsVUzxbL1YzmvbnjWF6cxylAtUDkzeSR/+3+VA1AE2WtS1eu
oUMNWaz37eKnqg+ZLTNLd88nLpvsZMAFoX79IvAjBkwtb48tKevmlqJGgPK0
OhrXMr8wxdBpZyckuKLtNvCPUM9AFmNWZnzQHujdO49oeHib9TnkBPQx6Ip0
5WYMGe91gfQVlayourtmDoBIYqEAttMaGUi+paEJJctex6Jhp5qi1lu8nA8G
5H66NH6ek33eMkLpZQJXmBFhl4SsNrzfPqEF5AXwc12YoYeEoigH/WFwjNUx
8wZcoQHa7NLoBAZWY/ler87QzaWEWNx0lU8uysNRBwIk1nBWgyLCXmtYU20E
rE+UpbzSt5e/I0gGXMk5aDDjWbwZg64Cq0tqqIlEBdXgjLC8vDJugppvxeLr
FoJvM9ktOII12pZj1WlPJ2Tlafk4V3bwcCd0OH6bdBu14GWZIcFW9scEvytr
abwnur/rqHtByRIJArbMdttnljIgcArf2QCxOT5RebgIH3/C60F95ieIpTW/
N0xobbFs/d/7cynFQkckWGRgjP+FWgSfjuvdIxw0+Ja5YDZFprwGUTQ9GLQM
NDgJUSMuGrrg8FKc+x7LJQF+NvLN4mL1681efaL2cXbhvn4MKDSEvX47mIJA
G/rtOiuvhCBmrillDoQS2m/dKhrOBwarhzwtR/KjwDKfzAaiGTg2fK32wouK
k7QY6DkeTTjyeFYqxEfBftjChoFz7bFydz+YrwWf6PKNFK50mgz56+oXbIsr
uRg4+MIYgJ61356IAPwGfT3M0Jc3dZtvTGlqUFJ3Cyq3ChxRFNOc9ujWSYfj
/3m7NohCa++N3qNb6bTP9XOnh9VOtc5oZbNF14FE9t1uJ1EQxClUse4js/vZ
jnENhbnKK0mcH/OIIel4I0FijW94+RxVJs9bl5KA7XFPtSP8E8PJUnTHbFg5
tPxoIhIz8bgdN6LzB1jWJmwqx/VvGcKJmzLWhDxalt4VAP3u/u0QDcbQYas6
Nrsa8QazmBjUM/NU9NWzWUVoHb05XdbGDPtOqsQ/PXn8L55R0YQsGMH93z8s
MCgHDaJeWy/kH/7Z/s+F6LfKH4Mc2p+BJkfAtXFruC487/WR0ooxi37nnjM3
rHzgANNuXDLCZbtznerT+QbZsoMX2CZEpDe8ZbPiDjAzwFnFC9U25rAHzid6
PPPI+Vnb8yTPKefkyDhAwqq/8e0fE79sznsk6TmK30PBS5Vnf0V+leQlXIFO
+EA1syueeE2hXjpGjMKRGgH/DgHhunztov5uC+7JkHASivHpeCyP2OzEi6Sz
iaG3RUw3AHj2I0jgKywW3B23f5cFz3QslsQm96bOZRV//Fkqpcgj2oDfTTGL
yr4s/2urxWV8suj+n4mzk6w1+r0J6LkLW+v2d4X5nIPmzLM2IG0weu0Lyam+
m0xCWA2eRkYobkvIjylVTeWSnlJLwM/RF4GUpNq53SdYxOsl8mHbRaaX+QcP
Cq0MCBOrYiqQ8Q42kRpDwD7zGV3Tgq96Ftpmj2e/5YNqd4HUsnV7JLpH+Z+x
rWRr8JbpWaGXm9Dp/2fN+8ybhjKqKnzRzUi69rWqn6sCQtrK4PNGS5P2eIS3
axstuimERVoPffxItMOa7gPCxITv9QW2VpvZpTA9pB40D9J2ngL1c13z+Jt5
N+SNVUsvxbl5r1N+zzPGk7oG0+GVg5xElsGFYvgWidd5Q3o5EgVtcpDiyjSH
H5Dp3gdGH92pbur9SzLAiRXGryjJHfAH5HAjBzmfGSEVo8m4TFD/F8Pv+nIk
Z7gIo9XYBlMRpvbOkJvVYS5JhkvM2Rn9YI6A4l0j8AccNncrfDx5W1mxBuO3
FmvjGtMrwwhGtZUygSAjLxy9itWiwdS+yQhFgwjfQ1BsBqhABL4EiXmd7dZA
4TC74BUf/PsO+ypQZJBH/qyA9vgbXKLUNqmYYFQYgR8QrtJIXcc3BY5hZmUK
L4Cwpv+LKqPrsiJ/MqOM/0yjUWAwNMVYlKB6kW5McQpq+FmCvm+c05mcPu0h
2zBF/ZXpvvqHgEC3dYXSGPoAczoktTgbNexInmYgb1DIGzuSQ7RpjIo9+6f/
bJXDJwo9gI8nPF0Ms3dhtjfbZmp5wl/rv6O71c+hQO1IB13dVekyaGgKTJOJ
3sexMivYB1bsIRPxOWlar+IZyru73ZgdMlVNzlWSWoHxJJv8l2QJFY0KeYjY
q0IDQXM61zF+BIvcPA01jhM0WAilS44lW/GKf+HGNgHoDgIGeZqUK/QMU3cH
/A7g7qgqPn9bhuC4aGIcvvwJ5TSKiESD7NuO9K5ZOsexaWxwWooTcI6eIJbC
HmDhoQ+S+3IxGrBECLz6OEqT3Z8oofBG53cZ3oZXJqj9Od5JWWfHGM6SadTU
aFTRX0XhSkbGPofIIhP3fyHfdbI0s/BFruXRfJmxC55direyLgSz3GkbCIGA
R8zgaBfhk6yYZG79DXhohv2nkZjY2twSLqhxnKrDVziGI78pfY9Q5Ad9TxF/
2j2N7ssLqhn0xYi/14TMe1/GXu0kvAXVYGexF7eG8ZImzINFVV6f+gsE6Wd0
C/w1+0CzQDQELBigaPtQlmzHjBZkBvMikI0njs15Mq91p+YYRxt9N9xARb9B
VOEjC4Twz/ov+dK5gvbQ/nbyfrR3HOEzckFpYnN753Nq4kT0dazdCJRqu6y/
ZR7ZgXHFaezPhCrOiIrmquIGgpe/dtojziUOg+jd6LFIKJVdwp/klqaJuxfS
49b/hXxIEdtIr4vxSkJpW6OI3qP6a+EGJTigZfKMg6SDHiTQmtQX1xOgYIlT
KIOggi8X/I9Blm70ZVTCl1wh4JpuckOSbWmrA0pDIcHyWlO36IniOoj9BwE4
ivEA67Lde23UnIt/w6gLoJ8X9TKry4aT83otJOu0e1qeW7W89/EwF3rO3ror
qMdrgr2WO2+U8aVm4jIDDaFnvxCCetTwVT0Tw8FSFS1y5h51TfD57aLolMtP
ysxcoWWTvJJ49ZPSVyp7Kp3OYkn11JvB+0HGcbRvrfn8Mg5sNwW0z+zrSQUH
KBDjF8e6JKMBjKGXWiTztNJK6myind6pnclYjKLgQ+eFlayKTi3mbEOn2g/8
KTQ/jMd2SbRUiTB9+YHAXADt9lICvkzFnlSPs7SlvYmlK016zvf4IaFY0OX9
Lzr7sD98FaqV0wyHpg8MOgiaG1tk6Bnrw/LaOl3h3B23MlCi3Ib1TQd10Ptv
FiGj0NKAE3Q1harQHh6i+RM+YMxOt0uRrVHMKbcojDosJhKR947/R9frmv+O
G9fofF/Lgso0VLsShj1n4YlmkVT1TmIaciQsbVE6xYH6O31BETVwq9LzBByR
PMioJnrDOqEjrIqwG+AcoJMMsaD7MaSN1+PHTRFl1sja+6CZxAbRrn1nKkMI
AqbCm6mCuKUrTGx+kjdVfK7WBkZf89/M+EL4VkisoD3om0lgXTx5pbKaN6T0
H8X4fkYIJvGidSVFhEiPiIZ821v+3k4Ak5koixLcPWV0HDKerri5UaJcBKEd
NxwVznBxZAYLEa8pp46Ph0VlfW0F0UQ48TBRpcwz/xRUXFsVfIudHtpiTGXw
hvXN7gXqL7LRCrhEH+MNFweCRb4usJnn7sccyrSgnWkDO6wZPRLcZpT7t2cL
qstPH+YIVRkPTIhGydNhtgx8E7p2gnIahEJXQUwjKlDi/thHT5qda3ClRovu
LOJ0fdlzLVIu3Wy+qRj8CSaYDqMVmS+vrxUkVExdIga6E+SAVNd98FBuZhdB
YwIS/R++PgL5dJbbUnWDx34KbyUO2uVYoNFolrYleH6p6CLcgI3u9IRakSKj
R47hrQEMT+gZsKz4PjRNuNDH3Jk0oHxglAiWlwNVTOZxSLdUbo2pXNX9mqM4
CYQcoRr2Ra0m4N+S8HXqpPiCtn5c25l+Z/+Ou/phFHrAdOhDiKZgDJJu3klI
/ZffeYBpeK7/TPITrmu1YHRPvNKBYNq71C5pAV/BZOjBUMe/rTG4OsIp7z9q
l1dD51Dzu4M8jBORx6WiUyvSCR+yL74BsFT50WUKARZ59shQ5ZOxUyEIxAUk
GHjyrKjBSSe1gaBwP9elTS7F0yOPUM4Wt2NMALmn0z8HDwAE2JICB7qoDKog
nUO+E76Xilc9CSyh3lDqPMeodMwHnGQ+trlqCO9ML0OzDuZRJb849ISTFvt+
IHeF8GfkzkBauuxRTLHS7YAaZbHWu047ze+eAQJECpxfycLyWYovJx5o0sHs
evJwmWQiAD1h441KDuaK0CYHP63NzF5UZHsVJG3YKPU9OTKpcMeVELbB9sR5
jkRvOye7MwM4CiSHKWo1rP+lPlftkb6jpM3Wncs7RoL7E1JeznL9rYsiGHjB
b0uEDEA/rog4FM7VFdL/b7rCeA5Xz9RQrkLN8pZAJ/03bHmvaAEd8bMcc3W/
5C4=

`pragma protect end_protected
