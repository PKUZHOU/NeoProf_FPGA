// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
QG1piTPrbobjvbMzILrUmHxHuVTIqYszdg0Iwcc78HdGdEk7/wGLCAYhr0HTxCyH
FV+LApX23w2l+y7XiFjqsFxKuC/jRWLq7mAGlpjhfKa5u4NaAocE2sV1AQ7rSUCY
HDBWL/piZgUW2xAJtNF91JZPdK1NI+cEc4qX+ivO+iE=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 9680 )
`pragma protect data_block
KONSWcFwb6Fy0HgQDilhgZuEv161YeE3kr1hrV3zJ/ZVYygwROcyMI7qDoSYnDgE
Uosc47IwdXrKYQWeiDNwFSCC6VOZJykst07IMeLmhuVlIviT13X3hiH1VxHzF0Hh
NAtuyjVCVw2vtA6PxogGzFdSw5dfqcBb6ZUoQ0bRiMa1ipcCK/nkAecBSKYYeqOe
cJPWk2LfRd26rJ0yt5TESyS+ZJEo3o5YEM4FJ5Oh/DhCj07VWEbP2n/HVyzwl42u
L4fLDoFwz9njuIlEA2DdNk01e3uM88pYbYhq1GEoAFlwSwTPBuRKEbYHhd7kTv66
gul6uGEOcjIMSqrIoj40DVTtpOYjVwWvobI2Gkf7msaL+ehBQFcgdrDmjQTyaQXj
ivLyhJNCXEZcP5QPgjHQT64ueTbOfz9EZiFejCeK9yoXFWYnWtzjKfX32ILILcKl
cpZ6ghxsmlXLv942BNNQCgP8J4Jj6oES6uS6onY344f99vKkq4A09KMLCMwiAgt2
UzrBu8sAj/dGrdN52wu6dPLacri32L3CNt2zSPafzSsU4NZkcKdIX3kInMpB0LS8
m4YzoXIKllVAzSWaF6fpDzBk1/VhPMGrVoPY6nZbePuf7e9WpYv4+BzTgrPrIZif
X9zvT8YyYsYoirP86cksoaepEOcO+B6aTjepli9y6UjGzX2suhIfMuAOfk+9STFu
gdXkxmu95gEjQMVvk44N6XxhjpHo2sMuIkAKjyr5/Tk4unKbrMtuJKbNM6/63ohX
wQszKO2UWdtOvSbHg0XWrAN1WvGLcA55PH3HJv4AkyDGUUWFh/VnNYiZjicXuwvD
72zzghQWhB/WqCaJU026MddRZ3fzotUhPFwB8wiK52t2/q6Md8Zt1rBYfT52ehDo
/3o4VM1MZ2ojX6zzhto3sz436JidPSwiCP8Pjk5amzFfIT16XIKa4o9QWUor28PK
xS6Ig+nXQyBmqRoQv3URjkWsPxYAg9VOf5UWiQfdqAUJ17yQuPEkrKihX9KjZCi9
o+zk2sBgq89SEGd+bChM6UyI+jN8BDtUPUHBuiGK0FFheAegCWiZyv4akKhK4jlc
KHgUiWo861qsooI3IzzHUbBPnNnofFHG0lNgElB+XbskWESWSNvuwdIKS1cxxDak
mLYpVFHs4bPCpeHSvvgw2n/VQIOx0rvVvYKPUsKxkaPmeWOgbeoYTiQGbsGWd6nY
WvxYCq8mcbFC9PujkaclPbouUNJVvwfdCaYCbq3BUksh3R4BcmTR7WHvA/D4Me5F
30j/6ySBNjWQiVJVsBJZrdr7Eil9B6h3ibKPgsP980veKCmfiYpzRGw07r9fT9J2
TmKNKyAaAxENbZ8rr57cEskZKa/+jI8n5U/BOjFdHndP9Eha6qx0SH1Mwq0DMbur
oFvFPZ/LFa8zhj7Y0kZHjIwhgcgVHmrjMhnFOOjIebnN+5Mkjuq9W/pVmGhO30Le
9IWD6XhZWA1/Q9D06qW11GGEt2orPvAPhCU+m4mvkjmbELHCrklJiG74MnKdk3Ab
AvdmDkkzmaH1/4pgQW4kLOa48xgNXSoVqLugrlXQ3PBeV8IlXZ2yvkafceMHP59x
HNMjpXgsZRShjvQ8OF10cg6ho4a3Qrx208ciWQojxKnNogC0ZBBzLAhghSm1snch
jZvgmCn/5L+BzrclqUaSGcM2S+U3Q48trXO7YJaWZr9hbtzXkXWbjUjTRYLwe2a2
c0CTbLMNoZlQZU2re4niDFERxtaiCZl99GSJPm8kUxcM71AMc6z6YCVsQAkwCrhT
afJxS/grSQnTJiNz4Ufkp90x09wWx7z7xziv9sNSgYZn5uQ3rlFPGuWyy7QyF3N3
deYM6pXEz24vzdAQ3HDLQdkLs1StBRQzHLHxa96Ud5dP0XdI0Wt95FvqEqfzqyEM
QhNCwMHjLkcF3sHHvaHdwAt/23AL+lYKWQ74Yd/ps0xEOA6vcWWpke3Kkg260gMr
0wQgoyIEuboZv/gXvDCscqGuZTJnEngEVyy1iky7k+nJJRr78+zopVJB+trC0NBI
DHtlleaUCGdYugg5qa5Ii1pxL8SKeL9d+zuVCqY5FjPgPjOz7sPoIrGi7B+rCvJ9
6S7jamapVMr7610welNiHvAnqqC5ApNw4jZoMws5/LUxqDf4mFuypwn8/qqz9JvZ
wV/dqkXOFtDdoLmXX7l2Bw1t+W4Uycd0XGqXfMqWcH5gM6ga2ng6xexsXqZF1ipq
fumFOybj7pXSPeF9vF9lpGIV2akOpNVu02H3YxkQEnL+N955i5dXxEDenFezySaT
4ggtSKPOuk1l8mz8Pds+w6gS3qP54Qmf9MA1KusVRhnb2BVcur03AulQWhnKDFVQ
319E3dcmvZ+Mp34KnOKSUqHXCCDbbTbG+3Olx7/r5+3t0xDr24osKtLUBZzn2aGh
41L7cahJI4WLvPSuwfIeSeIxvBaYC06ltQ2BVFYy8U9Nua1M/t6f1S0TyJFhGcF8
vU1MwIII5hYUb/4Spq+pRFHDpnCs1gwVJbYDwXKJQIUVIWC3Inr67Gk3UANQUBF0
JJX1N0Pn61DEOHseYroFaBeFYPr5eAyCBL2C2pqLLqOkHdrSqs2kap4RMJlroteI
GLWMGWSFpt1u6TD1ujWplwg3t/rW5K+xseGDVCdja3Pc3A6+OaKp5ba5NOg5QIot
eV4gpLoUUZ2RGGgDMLN/xm5NTUQz3JD9GnCMCKZ+J4p239V7rv+GolbYONr2eRjp
pd3Tzv34YAu2s5lcUNLdG9bTxme+RWvyzsGGakbFzKfk++LuE9ADsj4anoRge71W
tXAYkbwbzp17Tcm06lPcoKSA8KcV41KbabLple8jtQWe5IpfPus5ANnSQWA3JBOV
L0/f1Edq1b5yddbxSGFu8iYe0auI7WBc6UmON+Ogm06vHd9cjgAaeThAh8KcZR8t
XJhZ+9K1KHzN55iMsSWgNmGHDVhVYz0nubRplMeQ8H3qEtU1raBra5liLmLsnhuh
bEhbS904YBSP/Q6h+BM1czKcmXidFZyVhrtemK3q/mD9gB1F3zZJgKRAyXGbpfTa
OpycdlkKjF3PZFdOpXZrlopKUnFsh1IbbUMzJXJzeiJ0v0jhbOoFLOuN5HEU2Y2+
Ezhn0nnllPXfNB6vQPcq6Oqg4WODGDdIz3wLQIHnXc+xW9XZyYURGUoUZNcgeSxJ
aWzOlPTYQY0hqgzN2v7d3+LWhc+oSB/eTqg+GD41ZtGNkUT+j51n0/iqRcndwyOQ
0p0Y7XBqghOfXunR6rErXfxBQBzqyhjWnm3nSp3luaOzlcVjGZawKNfZtbNALBO1
WUGJZH4ow/0xIofIHh7hZng+D2PX6SXQTD/BssvAWE+A+zg9ja8gVVnVNTwSvwT2
yB6jkKMK07tV2wtubEfrytmK0WwLpOlLJ1DofLE5LCTV/7pWJto73kKlyhmdiJhM
mX/C67GTXWsAtqWS2YreWM/eG7LC4w2MpMHyCBadrzoPHIF5V4U+YHJGWK1JMh8w
AFwdkAd0Szlxw52OqVl0ZyTT3JK9GA6FCWzeTc59/Nfe2iAnNpdTdva/LKI7jhzC
3QYUzxJN9wMEG0Ot0hp2heqKbES/BnOzi+iuHmsyUTbQ4mQmdw9PI5gSbZX6AmNY
hCN3iXDCOwsz3NZII7xyXub6m1OJEzfgkckUlfwiLUX0S5sS1GBPajN7WsJ2HHIQ
Eb3ZomOC1Lmn+uXpusr/4ep+PL41OXKtVH/hy7AatvFtCRUrIGyvhgDox41lQ4HX
GdhFatjlnzJcst4oBo9lFqREUf7z+NLQfnPgoncD2NDjMjpOZ7d3gy4DJ6hplh/D
yVgruLcVEh1Ea9Xmwh/s28eR4ohk0qxJIYWtATB7EJfjGRKWPXYNH+rFUINGMIuS
U0ziYYpjcAIjFiXZx/2Dix12oPHK1SA8BynZ4TgQ14ka6tuM8/KV1ZT9azx/BYc1
SV/YSF3BHC0KgbxKwgKV0sGOp4gH08eySNPbEohoHSXR90C+UkRywc+UWxmSZz4l
vJ+P/aO7jZnKMsBnv5Lw02vsZQFy8JMs6Nk+40ifFGDAb4eO+PxMzEfCQd9McNUQ
1svvpLpsWN67tCe1sqgLx5mmIWiGCz85ClscA/86vgiB/XO2kQA1tTOu9KphJ3IE
69msbp8XkeoBX7RLVS+U3U5rW+B1Z3WkMrB3P/6Dd38HVVC6TwmOZcyIoewXw7MD
Fy/8sginEbNUK6E0z5MFKkV6F+kBktgunFOWHx8E9VAUB0JSsVFSf/oayzvcYg19
F7Eonlirat2gm7yVsf75nU+bkLf6+HIAz76JMUPpOQq0CMbAdija9d9LC0aOhK5e
KQHdo9tESYTi6lXJeYI2WCISQ8BRloLVuZTUh7cikX+uPE8kOGaWzrdFcS+u302o
hTUVyitKqLTUgvgq08lzaX++zYWa8RfQhsh7El8w/8VxS0bTyQM9rjznonuhRPa0
ykd2xLW6FtNFtGqfBFGDxmKiIRkB63nIhJASyLD9Xewd5TZPLv7COKraofssY8Tv
FKbvSLhypm1iXNHZaeWvFTl/on4w7C69xYblmhKz8mAwxdmuSt3cZtwmkIHW2iiR
mGmg8/0atxKiDiB3TfnDfXuzqeoT7zJNCAbSLZlAin+Xdc2tEgCC4v/CY7cP2iOX
zycMkuFreqOtKlYjZ+2vJStySwBclfMQ/sTARGcLh2ZZXd6jItJrmVjEsqvurOlP
M/WLED1txwt0NvMgEsPRjEslDRW4Ory6+Fzin7oLDj/fqFk5sjx2F3/Cqmbu4lvU
BxEC7aGH+u3VI0EEGPNAeJoO99LyPqvXV61U/BO8Aq3GqE7SxvykRpNmRwcyO+IB
0xa64Hl1DhDH4PFXMj4RF4Wl1YpiUJxOeYKvr0m9ZBvlbBtKhIYlNQx8hHBtlmtT
+xmtYTpvSvhZYmgqE3n4PhXMK1qnBWGDhH3gTmMo9p637KR0o3Be36OkI2FFj+fQ
I+Ta2fW9/yImdJH6n+HmhwRL8q/z05vGfUeUiscTQEejYygaovtbLtCjyyn+ppK7
Tu9ZeNioyXVhHc0SgXtuoU7+PO9B3SBE0xdBtmJhw/aFGrflwSJP02WlepEI2QYq
ZZcT4vSRZ1gn0v8qvYbZSVAc9EXHrLu0q0w8qsnJVTjWLJIUsTxDTYU1nnyBUeJP
AxBL2U+WfywM60Xiqd4fGwM5kLkvjEk9IEF7RLeh9pDu/6Zoj1wj5Cxl5nM5Gysd
EIwNJSf6rlCxB52ZQQ+PCbbwJB+lX/++fLwFhb6j+3mfzSP0biZM8s2qB6dSnZc2
9496BUGH++A+gwZDC91AJabRH/bEFvifUgy4XDZxKUcRYLu9WZ6qLiC5nAIdvtvM
vRr/RQ5bFs6J1eZfWu/7zVmAW9gVfGvodE45EE5035cvW81FuZaqMx1k/bVu2wta
4an1n+RT+ppIcrl+VeLoVRGly1hk9SVaAlE28a5w7yoEbeBsFEq9S3/+4orxRPMk
G6NxTo3CZWm7d9bOne6KTRQZuLkHehOeXGgrrOaLmSVFPz+kp8x8GnaJgjyKjJr9
kl3VPWqijzuCYvJqY38dHyD5qbhkkiuMKrY19huP43lmsVYSZFeOmONuyJ0JR7ft
VtnoydWolwNjPV/pF2gWoencJZSYZd1+3rR0o4Kb1WOsnBFW4h4aF+bbwNBQdvEb
aSz18uYcY8nVvT06L7n1atqbPOvNkd6mO6Lvucm4ERoU67m0BYM+T/5rS6R1ZAzD
za7U5XhThPW01d5K+5UHi+3wpKsMjPegp+HeG3FciZf40b5T1sMX89uDjATSnk0L
gMOTLwXNO0s0P7x6XSJzVp13pn/D0TCU/xaAuA3pqFjZejE8PalKx8F8IozgoV5h
Ba2kmLg3gJFmWb6+Jc5LFCO2ZGOxu502WtblBsi0S364JrdMG+exZ7FAJyAx+/3s
n/plsGrsenjX06bS8xDG1MyxKNtSkqeFq+JvoRUesuMjimq9LZRa4/wk2pgy4ocT
yHGKlpQ9386q3YsCHP9r96jIMQwpFIbQkZjwsEQrEq1cOP2Cd18W1hzSMFLJGLBg
kemQ6cxi+yhzPXZFO9R35PwKu9SaWAlb0GwDX5Q+3r+wlkyfBNi1f8zU/YyXuOQS
v/YLOsb2xzhmMG9I57b3Z/lao8WIocM/9OYfjEdIT95/CMksbzrrrzvZ1qD4PzSG
XJ0mnNudRhRKnGSbU3+mzHKD6YT4rrDUxxpbSJO0e/Lfco3Jsnkxzb0ZZpv0ODyk
mHm8kybERHL8Oi4a54vicreZf0+WyhgQl3JjElWX6PK4ls3XR0FrB6FtJhqoIBFe
KhL7MlVyBmDj0/L20TUfjytxTGmlxZsYbdpfyF5IERkeMFERPej2skIqcgXZ7VtC
tc2cx1AaOqrK4a3vEE5+5tm7DeUpFVAsl8MhsT8rmvZL+ELSOTAXpOxuHRjkNXdQ
hkEpL6PhwkHV7g6+kU9Sm7OqGeEPPiYYFd0cnxTMa+oAAOUbGXsC4v4IbltwcpFW
gPdHA2zGGKQt8FgumTfLOumizdwJnGhB2OQ3w0Voa9SvuzVRye/eLQc9k2ZhLg9s
eO//aEnCrYTkfYahVa7IXYtmGT8S5uV1fi/y/dn5tZ2udmvtIF52Bil+jybAESoT
MaYJ5Qj75MpS2lcE67FDmqtWjn97jGc3UaMKLjRU3H6F7ryCWkgg4yekBl6FACuX
br14kxLiUR7KImi+njU8+DizKmObTLFp+hBhntj5IziYv25ab5saqh2bAykvD8VT
ci3ZxW2RH9EbYpEuJZiojzqnJAGV3E8+bxsORKOXXSicYak1GHryYvceidQEV+MW
BW0uFuMEa3CsoL6Jg7shYWlLrqa1vBIl3LJ/jUfmovUdXSIorgxA/Abr9raVKsSM
qhD1nQtG9g6c7ZMOB9bGloQzjqp6uNtVUXFqmI7C3fwaS7Jojqt7bQFOaALpf72e
StFt+0U7CFYc6MIjS/8wlJ8waL5jNjRNVbzekMZ7wVK2+xulKCr7DwKDS24z0/Ei
hLD9WqflVbFyU1tGJOIG07d3IPmHq/cAXWswTbi1Si5A/xJJQ3kj2/t7al9T7Z8M
EiwTQqcfpnYsz94HzhU9urzcu44eU3fFSO01XajqXE8LB2YYVzZKMkJ19HpMZkXo
a+2106bPUXG3nK8JOVtLSrUQZn8Dg3CQ8NX5Aw7b/6OjYoDS7LbOq6AUpnBp4u2d
cgtiwVQNQcBxbQiP/4qoZi1F7iTc+Xkl50sNyVsiSZIjf2/2rnAQku7r6JkAqy1E
xW6CWYuw8PIWJGxIhXhNtk2dSe1kJ/1S7Y+bjdBG8b8FPN+5d/pbZb/zga7rtJo0
GA5NsjqSfhWN1CTLgPx57Gf58QujbzOV4qfmaNNMZVx3Ugx3yD1fI3EOyrnLXMN2
789VH/O2zHBKSEqirnZizroCrsx2BelwtyzCjIw0Ww3TpgiMvh1YOubhttK2TM4y
K0IneXtnxpDw4kzV1dSVqnaZSS/1YFHmq+8UfNWqd1U0066tAKbQ241Kb234safz
G2X257FW6C2MEQMKx+BFGjOaO0sGlol+mqD6X2Nf7OHgwSH56zBq45Y7/jn7LNjP
aLh4SugsySFrEp0KZ7P6KgeTrsClDbJ9mGmiLMpEqWRljxo0sxXEt9m2IhZQ/mux
M9MFqiQEUpl1brHAF63uTlE1cDzZJQkQLb2mAGMA7EEdwWABg/Q1FQTwVYHsNnq3
WsPSH0TgKaLqDdcZY5uqbF5ImXT4dY6Lv2jp+0jDcnwysQi15JZY5DfkkgkIPVtf
Kt3zRdgHoeklyXPETj88KA+gMpStujpSdyGrOPbIGIEfAwtiBtDqpuqcUOPkWBxO
s/n0+kQ51YefqSlC+7N4XIfwVR5V2mypRNrE4ohZ2s5r78cLyQVbJSvf6UL300Ha
Pz1nHjTLazlOe3eB6pIFHuwpkE+7GIJOmOknJiblSWcR2YxHhnkNMaR2xV/7eW5V
7f+9552AI+9PHsK73nzd2KkrtptQg1eAw5a3GYtWGVZcNhgo0LaysXvLMxfBCKWx
6qVDjkSwtUxS/1hB8Cc+X/EZKIl6mANV2Hmqc1ABtPyJhAcrWlskJsZY3Nb0EntB
xFKcDuokv9hOYbfln13ZagVMLQneu8NTWzPCq2gDqVwVyVVMQ8NPNnJAZOOZzvO7
cwBA06N1ynPLMmPr/gCmCnsO7K7Jej5c9G16mJNdt0LbcBc8Vbgm+3z9ZrO1vAHv
1VjAE2S7yNqGe9uKYIdV0nIt55wiUGmcCwkSta9eGZJ2+mEK4bQMi+Z8vs4rMu9+
+pePaAUrMRH4Q/WcOpXkvOWfb3rjARHrO67l/wwvBJ1Q5OevO6prBWLvjcQwO2XZ
/ZedBHO7j2W0g3yFfERu4TRbiVaR2ybtTc4OSIbgV5AH4cexfIXHWFsEGRzEB/X7
CU4sfikKMXFFWdulFSAMnmke5EhYnHYwYjZmXK2MP8U3VQx/BHw4IX1PE75mShdw
02QvcIuObHZFXQ5NcwDCFL7lcXzMtyEmT0Y2E5DIDfLB8SGYByGo3JQKNXuBIukT
khFJtr62veccUcPEsgX62WdCtWwNYt8pWOgxidIwv+42aIFc3/3cGrkbHbK5uHie
j4kove17JCGe5V2K01zXyzEuToMIk03AscDt4BPhsRE9zSjRy5f1TeqP5SFwkniB
fKFy6mvIiT/PnHDEtR2o77AaMTT+/dvMK7pget1rjTZGTnnjr60ShLRhjG0VE+3h
QuKCVC+rOOERlrAHPsPU7GJy5hx+zvEyIdYLkZnTJ4NMdW95t2V545sPhK4qF4tD
SisJrqHEkaA8KODEHfku9EDkYaflAImpfSBsT5/Fsji92YdgD8IuV10CbYjNvXAb
mRs6YUMRzU+OXtjRW19Hiw67/0mxgMU4L4klG5WFetJMYj5qtY20Bwa7hBp2/Jmv
ZXqBpMNtJ3tpLy9pjCff46DHdGXGppzqencAmOESFt17j5llZU6475RuBxuC3NSQ
rZnpe9c35EPerQJVHq2/NTGABlYhyQ3/JBzOhnfumenr/2HwQOMu25ZjK7D3iCiZ
AG17uSoCiQjy64N/vjgnZejKGKIJ2JxWPe9bFfogvS1bv4CGkxZBbxN70aDE741t
qJEVipNpCewrK8wgFt1Vjc2nLnz5l/BzKJ57+5Fx7YupITUHntnASHuJ8tr6ikxO
aTxY3mJMEbjM8z2ov9x/TiQGsFsDCoFHTE/myubC7FPs1wmgxI8inSiddiGx1Jjs
hhQi/UOdFPzpslEnwNCUcJeKdbxtk/LPJ6HbH3p8N+j+BI25xj0yStZ3p+dlBCYi
SXBdvIzBkKiD1L3L4wVVht5RMAuUj6UCK6nWkEgl0CFBD4HaTTorerTdgurHpjfG
LttpfaU4Gz0bTiNR4EOMisu9oYqxF6fQ1x703eh9SbpRtuuZrgA7UCAeP4auFV3I
NXZg7+BKPqEz+jdp9I3jOmWgrzfL1Iik4721TMj3KexENPSh6VeYZcns3ae9tAuH
78H523D2EN/KTK9F9HGidwfgrT8PTus1HmHMU80tBZkn3FxKS6XHuG/o8G3ow96p
eAPG0UKwxzX1s1xX1gd0vRELiAKu/zKYpEJ9p6RCaPl4477kwvgBkZyFCbXCShcB
yDZIxQugw4oRpeSCNoanMbDO5Bd6ozXoC0mqCUgh3aQLPB0V1ocYpdteS3kwrpAy
Noq4FgsWeXNlpER+q52eKpIe927JQOVZSmHydL5eU8zY4LN1u8LSdQoHDuzqQJAL
609qXRC+ABZ1MwSDj2j6N6WKvvjYLVifMLs389QTuiQ48ldcIL5TRuYAq2UiroVJ
gUZB16kBBJUUL223q39pDfmmRjULFUYhSBekVUsCAHTbLmkZj0DVj1bg9VUreAv2
UMxUEtNgPtQzluMC6D8OinjNz2BwzeBiDRsoFC22O49/MqfpNGQkZGxriyzagX+w
w66pxprHjPlgvOieUVR0qgtCIv4B1NlffmpYR8oje4+2ZXnSTO5YfSBWiDKOEo9g
oRsgesKxWfTBs2EDWamuOQiDlPXr1OI0QL0mUOwdNsz0+qX9ZtqLmPccdF58e0mS
pUV3hX7GnzdjzbryC1wfdH1uHPmwYyGlWH3WVMf5kSlA0XNSGqYl0ydTjKTW5tE3
6lwd0wUjVi3WI8YI4MP1nzaERdkcRzo9/8cfw0pjQo8USXSIPj1wA/CGG47DnXMx
Xvlyx0xOTFYVk5Tg3DBD1SHnqgI7f25WVvUUpMDrxfRS0+/qgZ5OaMHcy7wLzFjP
kysvgqRlqUJYTaEchp6vNkUmAU0zlqJanT9NncOVoKnXSzoibxSPMEgdvIavzY3d
Lk0wOE/F2Nv30WCao3BFKqnlg81PAJNMrBeB0oMox36f+MGm5ZxS1iPnTHdRqbj2
0HLpOuoEeAA66+/7kZiL1PPKIrNwRRFWP3oTKDazqUbQhDHSVe6y2PpmRE+CZCHR
/Koagj2+xar/sx5iP9FtKFzjXTjhRPxw9JIJLNHwh4Z9EjjQlodU9lqdtuafPWei
ZP8CwYf8ZnMrQulNms+lQcKX6z8JhGt6bXcS1igeMrlwC0UIdOLkiYoOcADdQ0ui
U3UOp7s3ubw4M2izIwCkks/Pm3tRh7su+rnB5FFZBUdoUjkWtqrolGAT5LL0QYcY
iXA4n0OwRPJQQkxgvgZll4wRvSMBA/x1KQ7JtyqAhKOiqoS9xqt0hZelGU8SYjgQ
/VzzSotQFVkbWdbDU6+ecobbhqfVIyIbyIzBrcA4VPjWbLj+8B1smZqCzhYnIUM4
T6X6KVJPnPAdvBGAAuIcybSN7nkxSbtAkhFIv6tIZ//Nl2oJuBdsK+ieoStuB9mo
Db7B8SV2uMe8y5WiMWf9m28E8aXY5K7KynrPgYGbO/6sgYZTB5jCca+CnP+j/PXw
qs6TYmGY5SZ9UJdyIkP4srzrVLRn0t/JigKPGYISPAJ7n1QIZ+WMPkxRDO11vwMa
+AKA6k0IQlgnGqo8G9wZl3Fvj43wwh9sJMTOIHx08xyBZ+dp34H868v1jrFcGhsw
Dl3CsB9tBWYp20VassJNCd7P1z9eEtfAxndxAm1gB/MaL+PKBoILjsnBz2lBD3ym
4pnqP7JIbakY4XAr78nBV41B2grxer3iuT6TECOfk2QXof0fjI6BwCc4hBF8Io4U
5MahQlh/eRdVplbtGa/JrwDhLCf9P91UeKPpSfSXLXSbZr68yfqLVokqC4htu9rS
bH3JFwCuZ2xP3GxvbLVE1YguvL7L7OiVfCbNvYHH3agEFWyOzgtfL7xAuCHnuoac
Zdv3YrMjxwjdukXQ194Eh69nxZS06VNvRWt9TgZAtVCWNt62AaaE+m4duWDz4ugy
o7VQovgA/rM1n/zf8Y8ibVraYaBqAwvyCUikiy/lyb9T5HuGol7hMyGbCOZ29o+o
NsQFR3+sMpKqCPxqC2F3wsfIov7ois1wpzryjeHiw1lyk8by/zCLMCe+GMy+obWF
1bU7j2s0Hp1LD/LpYsXxP5HrgD5YN3S6VbMYkef5DO739Ea5BE5gnl5oJEKJ5xJS
AOhqhuHWxn7TWtpitGLfVDODYyIHL5apsXddPOOmfa7htjdBEM9Bhvak+NdyH8Nr
vDPffdrvn35+u8Tav2lbOEAtfYFfLyOViN+7mzloJY+8+70yplhGqOPug2S+IxyH
eRw81+7u4E0aa5ycPcfxFMT+CzdXX3BsZNPxaV+JgJm0D2NJNWmfEVJZn/BBE3mf
bUbi9VNn8Z+0YsWws3RVVHBaw6Jcf+A2L0wXSLBRMeLTwJAFJdCwAiqRjXlQP8WO
LlxJ838SOdqcUY81x5f1ZWeygggcG3gIStp4QhegeVi751ayD00Ggr0fXpoc5++w
mJLaC2dIb0KDmbNtLMdYgb5eXmFjmjgaU3lEPUes2P3cW/1z95dp4HGnpBeCry6s
KQkVZXHH4rvfZlSSVgqWkih6XbfRBsX4V06t61Mhp0SAGX8Safn/CjEGfgti5xxc
+5115d4jcoQ720kCdjMRX/z7cFAdVaKmMnoy72YYTIsHaDavHkrggmgme2d/+MBO
viR5ESRue9+wp6XiEUaIZvpr1fItaRTJkNQ8f+76S8NH5Sq30660g9kP29gTiNw6
aq9usYiFI7m4OSaTaCoDYlLriyfxFjLWXHZ1nmG4KcQaAdBiumo3ehGLHcVlqxcA
2K3P+n0e+iU9Gs3a7tt/4r88wvVbuCPvthVK2s61RVp8q9hTLGDniZD3pHQR2nrY
f2lnbpVVj+ZOLOTu9P7zD402JZX4doL1zGca2jcy/dDubbjUcYDh94vyogpMcZA1
kNw9fQboQGm3qD/YCplKwItUpDTkYit3K0SwOPjMqiTJUsg6kb4d8kAsFp6V973g
OKSctEeN4Atl687RSTZwizvUlN51tc747Ugcm2dEhoFKtMkKJ0elLRgDlXqjKxKt
BqWky5/McLwnDmCno8OVTVMe/iMv58lvSD3dgysIeQrDIjLHGL/IBfkmBefHErtq
meOMjZzaNZiPQu0c9MbRW9JH44cefBxAsY9nM5wJLiwFS0VQOX1Plja9rvBCbk3n
1gkhMMs2uQ8K/Hi/T5qGTYGycY4QzAqDEA86nQ3wcjxFXFJTccTehuq2AGg72S/E
/qrQi2p5a39D4v0U/UvZLhQFK0+zYSW8IjELN0BK3JUIvy3HYBi4X8Qjf702GV/t
ZbUVRQeFE+ArZxn0niQ90FIP81Aptmxj0QO1LJ2/9nNMwmkns0QbtH+pdI5/8Xrw
EZTO5J8sWX3MDwEcTgfRuT6W7FY74Cvfmp65xiFflFAeBULCuvQdCo8TbmuVcoXy
qfsdebHAXcilVLdESwVwAUOdqlAZWS0d9LwVROFUqK4=

`pragma protect end_protected
