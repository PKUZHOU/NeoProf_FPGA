`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
CPHpAZMfYK65hfyoczzx2Z1EKYMmPgXPJJbTHzferx2SAB46jYw7ceYVlgUxLxRE
UdgV9xSs4O/xNnWf4HHNB7NT9uUmz3AGnKu4JyHp1T0h11ReRq4w661an3gx+XNu
AllwnjyxYDlT3Bdedb7lGO4EAS/3QjPpojGZI8vg2+w=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 4096), data_block
/UlKDOMGaG8GRPNPbBuQe+G06ftZze5GCGBPx+NsRdIT26QNFfaGTUwko4riW+Ik
A3HfcTZmBkL0xdqaXvmqUsO8Ym9E1CxdF/fOeqDaxA8Q04z445hktkZaUwzVsyqt
M+fUcX2cTN8iFxAbVk7fn55lIGha63wil8XREqAsOcDrSUhXcemv3sG2aU0j60cM
LxIFUZw/jPq/A17owvIQ/J8s87FfC15e21nF60rVHkZAmUQtB0SB8omkBb7HSBFg
F9j3RIRPriD48ro7Qp7X3YnnbZTJRYNTzrJcA4Sq3tK2Oatsh9LrLVeQVmnZHQ/p
aLRTJcaBbGfLz4jYkg3k/IJurS96/sm3/KOIfoP1oW4hidJfEPgnOkUdR5lkLe6f
AIPUEu5mmf7wWvqQZB3PN5esyZerU8dnv9Qdf2ioALTzWJA7UVvtr6qCTi9dhBzG
rGU/+ZiLMqEifx93LxUedNYLleE4qnfux/E8TLBGgrIPBstdny2aXcXzd0g/yF8C
LxTc7WNFAsv73jvA8urjA8plZKE18/RKt/OTKYmmyyRxg65PTtV7ihVpNDCmVPMx
B/KKi79pC+Ocjwlhsx70s1cRKQI5aciIANSueTtuqcF6EAFN9rY/wCrrYHzkF9vn
trgfQvlRSnpDvDECwtyoak732Qz4F2F+SvZ3TS6CxbqO94DAL3IWs8KUolGIYhZR
M9l1cFJzkEmsPB1uF8ddLNdG9wey+8BW3pwB98xU7Mdi/rK/qtevkQhWGr41Oj3K
qaHjgUNguZm3fdYCmR2wYLnBQzNllJoOsG+z4bb/5fZqlaf3v8hHXgudnDX1Eeg9
FVLaf/wIzsPo5q/rrkZ9HSudxNul7LIsHAjVw3kDPly3p/5kKSs0z34MdGG/cka+
I03iaN//tVWZGuxclmRljXyMeN0pUZcHrIK5Cs5TFmUx1RZtNJjPkxOUwmnUo5LL
cOz4KHKHLr5WrGyMQamcSVrj505U1FMRE0a14eMKEmoNgKYTIiFtttw0FWAxxPfT
EWIrCz5Jz1FSMRQrGbXcBppRcWSKHzWowEBirxBkmHCqVHIthF/o2s9rFrxLQyFX
8BMzSh+D4rLgjvbIS27v+UP1zJBW7+PoqYu9XkIMNJ/6Tl5ah16SqSEQxup4c7A4
u6zZ87j5I8NoaGHPwWbYQzwXBOkpF7Jzj12JoO5ACNYpfqu27Eg0p2GI4Z6vu7OR
L85J7iHsuO+zbwjTHHe8mOKdAq7HwxKvokDF+/Vd8NHyK98y8w2DFfz6489PCkZK
AnRwd3K5gfjyVO5+XXm5oU1VI6VdxeQXY0XgWsBXZ3OcYl8menh2/oZ96GGYJxH2
UzMevHcTNC/C1iVDWQ6jkHYkgT03M8QrdGXyOG9oaHQpRh0f79pkLaqkZpS4JjAY
972DWXg02K50JtoQBtII6+vjzq3obpI+n6/LBrQsZN0hTfHV0euliPCWVNzVy+ls
8csucoycGskUrETRJXnxsHGL1AIJnzMDMCq9MS/OjEVjyZoiel4vTms+aKi0TRg0
Hj9BTGc1oePH3NMraWo1m36ZmWgjF5uo2U4ANOgACeWT2bvlZ4bArjQCimy82qi9
FP0LWD/lb59MZ84RFPm56LIcGc8Vem/PDMXxzRcElNYb0PTk4JWlvFL/vC6e5NIX
K+UbqnEoapkz66nqsRC4SrTtB1+uztkF6NzJRp8cAoBdipCpgUf9FjpaFVVM9gHs
6qQmifb+HPZeHRoToLUxaaMp5c/qdtzmoRmk31C/JFvud7I35Oj0MD9fZB7S0cWl
LiYatud44dyADSC7318ORtrx4LpPwOCkNYNF3aJnxMvdzrCTPxp5j1RzXfsbxbdr
Kl0AOIT2sH0LYkVnFEJiUWtvRWsD+q82GZ9dK7xcN9KvrtpzHqekRYR+fRONAase
uvyFcyJRgaDhT59StVEzfKhen+asjUx/QT1V/DK76kxCI+kNqUCqQSdPm04F0pyu
JIRieUK46dNESqG/JrJGqsEq/TfJnY/JZ46JLnyqx3Lr7gQs7it5e0nNMYvt1Qkd
5tyq9GHW7lhCjkX6fIkcl8G4DMvkNLTnwvhPInftfbq/hgHHWvcDfR7dj4+69/Sm
hocEx+12Qc20HEt3B1Rj0DeTBYUydwJxiy44GF2xYfG8mq6qN7mJ80UxnbN1s8Rp
BYSVVujUY/2IyH3nhO03c4BwA//vtYQDDzlrZpiY/rd8fcZlLS5MXq8HQuDnbsq6
ysrUnk7sxjHTHUH3HcSeMb9oAiWvrOCcwAFDGFKzNl1W8lqm/4RtQI8oBPyIVD9U
aI2zQ3qFGxiC+NpWBHwiGsWh79NGB0sEa2AUO1ovD0MdyAbFWVvlwK5kvABKHzZE
MPdD7SuBYX7gkdBMcjC/Gm+Jmo5DKhhXpKjp7jb7t5y2Nwwm4sFEId8UvDrOKXSN
Q3gv6/ANHE/5HGBp8vvVGbzP+YRExaTEQzi4jCTvrCO+Iup0fm0AXM8woGqC2WD3
+VluRe8R4K8l30GmPHZlFLqfK6sqIRTnIe3iyaGxXFXa9oFCLrf9fDkwD8HX0WSa
BdQ5aTf0moXoC4vNoXnyv3QWp78MwNQyX68kQ+Vhlecud/MC0dVbwZzZsnQYBMpV
pFd2gHXrWQSMXuS15FWh4OKg4ZrY846262tgxoJREOEbbdfxqXeSP+Law7jTeNJS
t5P/hmQmWR6Rvtgh2qh8UvaAlKscu1SsfYZSL82xzySr0F8ZZR90wLLpd5b7K06M
rrxj+4BVxuDzYROD5IyABUxK/7gaIYkMP0TvKyqh4aj2Do43DRGaC8j5y8mnDz0r
1FB/7kYeFzHIafaz+6S10UaqIPSmirkBquvO6YuK+OYF6YK7hrjwjghVlMncNESY
ZOb8+gim/s6LRy30t4Fub55kU+5t4r8I4S/fYnMXvoycWQZEORkY7aV5tupN1mqz
Zz75YzFzddSvthE6Svw/Z07lPgi4GYwgHBrOdsBV1+HBVspNQUaeDRt1RgXpr4PT
+xeVGJaSXHgz++K5PChKlyqUiSV7tmiW2nF97VZQ9b3RFaY0hdvS86qA+Pb9sJGt
N1N9oG7oLrHL9DsJC6XW5VSdHXlVnzu4BtUPusfLNuxvng4NOWJ8V6UToKQlsnPE
LxPZOJHISdzrU4k/ksC9mh9AjoH8VFQlHk12uDhm+uc7AehAWZ/2xI6GoLkP7uhr
4XcypvPNfJCHLxwkehgI+pMOEXuGYRa40j3ehWuS4Vz4HnC9igepuayc4Q6KBn90
d2lYuC/ZJcVsu2O5tGeknYWBn+T9Oa5nglzNTTZgm12ogTpCN3NWLGaEq7bd51WU
XwC3qsc46QelB65wIA0+29NlLVagTpkGlduaZl/INChUElyP4Q5vCQpzY07ged/A
kKb0CNIfynTcLP0mEiElgK0zRZpSPBqzXXqPKE6FaoxF+EwD+M7fpiSOOG7EfoBy
zOS4KqmPJoMs6+gus3cELA0x2U8sSWtya3uZX+zXzKCvr7JNq+4nEydrwGWJgT/o
hobRGLOKTAa+O+Wc/gGW/Kpg/QxWtLijzd3RVIjLOESq7yrjhH+6jXYpCgskOF1M
F0wz79wsIkjbxc153VVg2740erGjKjLgduFZf8Ao4uvew35y4cFxS0skftk7ASOR
qP4HvhUU0+HgLYPaWBfmKSB0VGxF5lkMBqAWPSFuX+AZuFLiF0S8ttGJc4Jm1TH3
x0bifDdY1SZUHNJ5XzXrAzxHlCH8Vk4bnL5R5uRswsQ1Tb0n+YMgoli9TZGQaBIt
0i0zWMWLaAOJdX0WGI/zRlIk7j2OajdRKUwWD8/KsgfVPQHml4WfWw1SBKWgQx8S
qIe84ldGByUPzQwy8Q9RuiWK8nFmmGqirXDY0hv33vpf+neUpQrIeC6yhqltkYMQ
hbvmVkzOPSyzy48sq2HYu9rE9rwDngpPjWJfrv/Te6NIgs2gH6WvtTi0pNGDEL2T
0GK/DrC8BYh4mujL3xfY9qNz5nFSmTOsDc6vibhPAzA9AVzJ0pLvNB9hTRyWwK3a
9QtWIA1/VSP/ZWnFkPv68NxGLtO8jpEiDE4eanxzx5as2ad24BfTyZ++K0mrxR8w
wMJkPt4qCPXN2qUpN35R7yqu9/oRSnPZwrj6oF/7J0BLXPjF5qB3whoKFsnACY89
RJS1fNjGET9VkhMt+kgqEqrlTAKnk3S2MzX6EwlOPndE3WUBEczMZHT0yViWDHAu
eeNa62yS0ZYC2YQDV/R7km7xFQXRqZwYdoINS9sbnvsGRcK9wGlWXMmnNKvp0c3B
alRaVYbYMeUA31M8l2/XWAz91RlAZ/Dk7NbchJSE0dWosihLTNS5OEJFiVuDrOTF
qI5BBlA0KbPjI0rYF7MKB5po1ojR9Odxplrp7C8kzJj4nzqsLaxpVmmfGQH7NqRL
sWTrtlYZlmpNsWbAj4j/pB88yp8Cydlw45knP9INIZtQBR5DoVb12l4ZkHFvUYHQ
L1dSZqM0XhXATmTg5WPuI+sDiW4ignHrKmTD6wFv2PEUQ59P7mtahy9CEELXgpH5
EyXIKzvEPQLEt01mzuAk3IjHialbzPR7HxDMtDdmYZvyqJSxHhIieRaGNUCUlNf0
styy5OGC0/H7vzJZyLLlqWCscXxtBnKtPCJmh7R0dJH1lrqPCniVPnrynW3qZrft
EdiyMqOtJByV0eu9TBBOGe1f7pjALph9r8o0UaRwzGqWmZx6z+/nfTYw0NvoxGXU
SRFSRm5jy4cndYsTp9p5j7uJ2rR1HV8YZSaZAPwtV6cMAacZH1iMW5Juhi9LfX70
TuvznFsmP1sqNX2EAJOoWWSZ3pOJkwPC6Y/DMTfmJniCN6slH7bM6oDj8aDrVWap
o15Qoq0LbqpSU7iePWWb9idZE3g3aiUTxehts4PKYswt0cZVsxHnNb45TEO3pjwv
xgS1+R7upBbBpeNcfMKH/1d/HKzn2B9GdfhNLR+HAMjRaiXXgSpW0wbdvuX6nwpN
xZOn39e+ec6i6HazKpj/sfj0IZ0tXEYs9sw99hd7b3WqC6k4MHMgT4xyHHTnXo8z
WDIZI/AMBpxIvvADiPGBlB9rMHqyV7H4Y/lMHlTCK00Cpr3g9kCqIwlO+YpfKTTj
bBZj9UW387owuYVw615YRfxrFV3pqlBaSxD71tXl29To9Iy2sESuj+Xt+E1FGIXm
cT3XJ6SXvM/ai+R2Q64xEVERRcu/Gb475hVVP5u23g5pcnx3L9jIGBMUr4JSL4zf
CSgYanPhJ3+1Zy2+NyL6gJROGc24Vw2yX9GqnpFqp9mTxb08dAGLpbsiHl6QLbWq
PIIAc5ukSKKxrUoxnMJeW258y8R+IpLks3KT1mMh3/wrDcTGp3ouowmS13bhU6Ag
5QhWAO3rmTnW09nsvIHa6bJvrKDvWOB/rzWghWUor3aLwY0zp3euhYjfgByos1uQ
RV5UEr1cMMQMZRVc4XEF4w==
`pragma protect end_protected
