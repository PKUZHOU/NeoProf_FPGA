// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
S/UnQv4KP3X+87ZLTiEPD0B1QmnC5WQtIGcbS12H/uWvwcWEYJFPBomPFEQMrwSc6/9+qrxxki/z
EouDce/u1eGIs9lppKgmwSGvlZlYqYVznN0rn3n298blqxkhy7psRxJo/cVLTxpc0MF9RzHnKBHW
fTEaDdBf3eBXLB/OEfa3ZZZtqVW8qT0s4bWBg15FmIK1ba9J2s+ooS+52ZB3WGLLs4RJ8fOgwINH
TeLzgMhxt1bg7ugE1osG5pF5wkQ7nH4Y7x2RhTCnXE9vp9whbyUqRobHSM0pJTTzEV3x4klOWqJC
app6I7493qxIHkXTq/Io9bGt+Ru5PkgdQM1aeQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 5472)
xXEAf8iTIWqkQr1g4EREYJOkPmgIAVQDdqLef5CzMhO8e1faXlOVsJ47pDHo4Bm1Gwx+ShUfUd9m
SFh9cJSBenY9v8TlyiaRs2aq/qlAcH33qMWiV6Up9htDRtV/xI/uj6HrgxiQwvw+iVnV9a//EI/y
+A5KHUkery3wCCVLAprNiiJHzazTMtj6kd4u2jcFFk6VAIGEFc3jTB7Zic4Is4RqZN/Fym443FIe
YIHgieRuHJLxzlg8gbQTp0ir8QFjZEmL400EhjiWlOHJMgodIcbnInpowjiTj9HvAuvTWEZ0Krp9
BQMprVqEuiM+gRX1F1AE5rcF7azAmlura4L3TxHSGt9CSM2GljZhSxnXRwvVrR9b+SOTNSRY1SJ2
II4it8DKzMviYqOwrndgkkBrIBcaZU+iZL1k7Jw3aiO/irRyPDmnFNXAJsYtC15QWLSwE3FIwCSr
mVnP9atBU1yoOHy3NQVvPH3KJb030fbOyXuCLexNVEsH+kCsSz3uzsKWEgIOPJwdtt6V59U8E2OY
4wiXzQ3Qzdf4lUHFudVv96tGKdPI1XKMdbJNIQV7Dx68fq2mlzXiLpi35tA4xgSxVx2LZOAtVOX+
k3IVcAnyrL3JU8iEUEt7jw3V0WgNRyGCKJU/QPlnAkrd2qQgKrOW+EhCsgvc0ZtiwMRfGnIGBko/
+6568q9EyHAO/j1KuFghgv+TDGQ8gFezxffjyeoak9OE5Y1TWHjti1qPrG35t4sfCvPNysujjZeg
+QPbcrt2gGB7JuBhHg/zG2ak/W1W28WZ0ZiBYKmpO14nOh7e3P6iXGA4Z7vUnttVoUua9JOgkz2n
Leiq9JiCW/PUZu0apC2rRrxbKZLulPIK24JvSCkKlj1Lje8OYmGOOf9F9VL3P5CNIQtz7Vz4pNI6
uOCM0B/Q3Oe7yM6eB5mNKo0VDu696f/+wjitHTnJ8caBf47RABah0ShJEWFu544Re8b/lDcJBht5
KioGtEz62AStPIJIJwinsfS+Y04F/WmSn295UvEpjA/4qB0ZfDGaFuZCtWQAtzye12YDd5cQqsqp
StFRLRcWLeHZ3/7liAGVxmgrP7zojj5eYgol5LIe8yugHW3U2OFjHxl4tsZCvq+cRgxwfm+VklG6
nCFswng0P49qTXWYQZuUKqZnHeqsNMff3dekFbNKH5BqkAloBc983W18ygEFrHC/17yl8YABT/Bn
9IrUvteO7ruSkptIYCBpd7GfxvTsIDdWAm/3LSB8HWXHFFddWlpjV7utW56Kx5yF0EvVNsOOiu+e
9l28ChpsJCd9tkNHj3wD5RE4BkYT3/zO5WjKF/5kC1jL2z+OkHpxPdQNIluMH30tNT6G2ZhAMDBa
qEqQyEtN8pUXbVR9qMJFEY9L0q0xLx6RQgjxwRU1K/0fuyQ+QxQO8sAi8YPzXEWJ959YiWYx2oF0
765AtPHooRsf1dJgtCmG2RwGkYK5jWA80nBbIflxtOcDJOk1Xl2t5OToLdFw+UqAQyO1f3O+Tnyj
9dt5fdlipLug0Zl0Tj+1/embvIojHOqynW2ceHVVBEgKF4uOkSq2o9Zwj1pq56QF7OBO74ws0fe6
gHMOytkS6z4QDYZpxucVISU/Xd1K7Fosr3pbTaWDrN78Mo72ctRmMePLotDqpWHFr2s+0KL4FKqK
ACQNuSH7T2pbgN4KswmrcOA9WZJjGILEuEj+AIECR8u3LI6he9pCabop+eNBLX4AEyg8KPDfUYJL
S1ABe0VXgeGGXYLR6dUwudmzio3wK5EXQz/YJ8NPzlzT+vNwdh089FAFhYKTO/EKUGKEwl8ydXuK
glfbI+z2mX13RqxNy+M/evHPiH0bXjHolXTsdezMatgCu36jelx+aPL1bY/UJwaT1MfmW58LekdC
csZT9/ZAozE/tsM9zKyRzelSQZXITDDoBjmbErpyolvwhmXLJ+5ZadMJcovZ//Gqqlnbio+IYTsw
v2jDPGp8lOqubXbTS7l554xSkus+jVzSwJLs+GWN2Ls3ohwzgiCY7lQDoBfTp5WgXrzeq0ick8dL
Pbw7EfNZ5JkyZFbJkYnL9REoMQbaPkD2IJnNrkz9dIzJ2w0GTDcRmt9Ok/c9guw4VrcQYutxsb24
nAfThm5l/g4RjFzMQYmx78Bl4O3ZIjvmAPgQttrZCT48C5ZI3IMdZggrbcYiHul/QMD+j/GXaAdj
bAHfrWf8vFTbURXE2+OmHQpor/9rtfhGUXoUvW4av2GS2NbKfnAXVxUcOjMIbBcY/8GfZlJf6e0m
VvYRAZm0q2lKTTjGbEojn9Wigj/W/wE5nzNmi0NkVGty1VTL41ZuWV2Huthfad6TCURSY43RejS1
lyxSlMKM+q1T1b4iguPbLHwX6G9kbLVU9MmGhGTj+dOhnxaCBIxGmDkpTvaOD6CXOgoA9jfxJZD/
L2d2cgP45tPg5G9ZVsKkeEgSW/hLN8uX+PwqHg/KGnq5C2sgjAQ4IIO/jyBG7cEQCcWoanzNwwnt
UtBvWAriBtWF8F5Oebkas+5VI+bwVpuArzzZ1rPQnhioHf8qnRphxa/pEVs6hOtc8WmduZcR8RB5
m+kvm0Lt9R3QN2bEX1wIqIxxr0wBgW8iSYUdxzipbQglETMD7vye0WPqLGlkayNJLSBV2i3PD4TB
KBA0hWXr65nXhDRwi72s4m+4R0KU82Sdv6pO2irEpiThbaOpAW7NcyoePSeGjPQ19aLecQOD7LmD
7Xx8VnrAHZpF3go6YNujXPy6/xK+0lV3ezFlyuM2rTXPk1ycQ9tx0c4zqDuVoI8MXLsdO3+ZSDhi
J0hoXmMN33+WkkWDyGn6RaCcEQ6IylF7l2VUXRarbpXRYpWqxUhDF6l9MpXpLquBGPWNngiNGgua
yepiT8hohe8oPginnfE1u1rRGNuB6FcamL9gMt8ep4TsCQ/qW7hjAbDTeounkCe/Z8uowyrYln5l
oKzY+N8qjs3cRtRoBChhO1iLFZdra8o5D/MVgh01yd2JQ7fpwbosT+2DbG6jBPKdch71TcGOwfSK
RWSRpKSBtNYXkriCBROnyJ8nK1UApLmJ1dtthmZTJq3x5yrjbNQrATmFtOXJ62xorTlFEI29zKJ5
IwpL0KDhqF5X+hG9hoZdZrJSjVxNME8vZOJ/bwzxRPaWcmANWHM73YP82nzmR1T2OJQcMWZCSMSH
3Jnvy/fop4wZTBrUM8JVtw5/R19iMo5anGhRub9gEhn4QGA+cZ3Sawzg1B/uH9nqO2p9HZMmbK5f
2909QruDwDnUfSLGh0wfpsCjYd6QAUW9tPvSUf/VtLuk6zfh7nIOS+OIOCdN3dCHmv96vGJ5DBgU
tFPdATaa5YshkURdMUPcTguskYzTXGVwgEMAaUeD0BlyHEgZXXboTWeQs+JrqS2/V5jbUJ/os/TB
PcfgeXAt/kIXf1EMmOZ4uBJ5wq1pnzsz/yrzrt8BwSFhOQCZmrfV9ASmLd/Iryq1VRN3WBV58kn+
1JVAVUggT4Cd2r/PUpKpCf+0xDoO6URGKylNbUmiekrk4YpC2LQicspmNp/+5uB3VwwO+/pOW59M
FKnmfY8pVR3Ot3KixKNwd4ClqQQQ9D/tti0kEt7F9a7WNK6rPGGfwMAm25ISa40XR2msD4FxMApO
5XSyirCzOxoNoUIv7h87M6IvewkNjzQE0A4Lc7SiYq7MEzct8ZqN9/iAVp6A3m3kNHcKgftezI3N
Tl++ByoXQrPgrcqNQ1W4ZekFi67PugjN73Bw14qMha+8SGdPY2twHEd7xJx5UkPfloMXjCl2SBer
MMiSzLdF4IYGlG+WM6Ca7ztWuirZzlJfn8XvBNxbUPpnN23YDrsf6L7gMu21v/hmzskHWu2NSLQq
xWo5iP4eg2S1B6dzpQA19yw9+JSKAQHbBR08XM63maaGl5X65xgWpZRchWfyClWjmE7GWywvktSt
qdEUoXiQySnbGI71rAqQ57qmx6cwyeXEvnc4499R91IOxUZz9Mjs/9TJBCWiw4FRFFe7yDGWpj5u
UT84Jf5kgNkQZ5lXKiHfVp3f/H15fCuJlPPp1+BALZj0wEzxJ/ycpYTEYIXVWcblMTAR9v19qDdn
OyuzFfbcsQPvySZZjkUnDntsAY7S3cP2o+eblHy1WBQuOuVmw9IgwXzcDaE4+cFOk9Kw6fNYFy5s
hhHKaFi87WrVXSHqRA1G4jStwfRBjAJQKOPdRWTEhXoyhbeF2gGPRS4zQL8I+LUWKlc5bze4IbWe
oZmMeCc1dg9RSbbWc1B/mMokSpYk6XXMO2FsouTfm72iSpWwviLnf9A94FQPnTJZPJVZhlaPY77G
pMQR6oWfiud+TCZrol9jqajoGboZ2J8qppwb9mZdHOCr3kDBekq6ce9ljvqgLrdUQiBtH7p09upv
24joLf2LVgPVVMqSq1X0GnwPge00ycf8hI4kcnWoWNYVZig2f1RKh1KGY0Lv4xEcmW9AUaxQYanZ
FSAGA5LslWd+LyWuFSPZUZrSm4tuYOR/jbLOmWHQTTZZiBwftxF3nPHWeFlgu7OwvdBK1BijJyRh
FMz532++d3sGyIfSa5GxO+LwfrIlhD6novG0APN67PVAQIxtRl14mp26OLs1bunCeWTXU9wmxD2P
HFYpLjfHJvKnAiyQFlFHwO5tlSu/47wFAifQcooc/MgVdbaz4665vuh2+ME3JFwgv8lUTRsZAQqx
mKlNq0AS+W2b9yV8eKzBxLfkcDc61/68cu0g0ovb3VTgO7pUHD2V8lUfDRDiJCSmeYgkfiWXZrjH
UNZDqj3PtkkZ228IdyyYKNPrmdC5hbuQXk0/u5UiaEHL6vWsGrBojxdp+MZpOJRrGI571a3nBrqO
B/2sgHcgo4j3mUr1u0E0JkDHpnpOKUK04Xpuh5d4JLTNa4ky4mUWviBHelorYL5lMttR26KFyX5Z
HQHOVTFsfQCxL1mZW15ieZQsBoEnO6iZJEGRFpLXOQ+rNxMjOrzIAgy8Vmdh4GDN6JL5sbNfe5A4
ZdlmVQw7ENeD0PIcffAZv1kulVqELoDrdQa8CnOfIkpWRu9Xr1W5jAA5Uuh8jloCIQsPKOdfqN3F
qO3bkeTgnmVZrUPf/ChoOMirvuJ+JBvXzg8Ni6hvRFx0xDh2QGSR7ONwrAT6F7nkHDMymBbgpE7/
HUeitziPZuyowxY1MsXmbGzTbDPzVN1E179c31YE9dSZgMj/Fp8J7HxhffABaqLu9m5wz2otazRy
w4SG7N1NZKPpC/34M+SRf/bilhyDlQx4c9AF8FAIoKzAsheeXdN46ZS4+YlwxTwcHnJWQbL+I2ep
X2hHBuRz7lp6+YoJOymctplvPC+hI+LQ/lJ/J8kfVsZrj/4cJla+Q8qaLO96FPj86zgF74/TWeqC
sX3JrgeG7iPC66ew63CXZsjGGYMt3RyErcsfQfwlan9iHguAYF4aTrVKBeyhbtWAARgo6BJ6955J
rVfU67tLR6XBTwLte+dI4EXRJ9g/Wkl6EOLkB+WUgYEcykgzXqTLOLgkmIos51VfBwdnyiAeUTdj
TX8f7JIrEOCb3zEtuwWLqNB0GpD8BylTCfl13iDRxabTMAQ+cV/a6JoadcVNDrm/gP+zuLdtm341
+ePR9SgmfD1am/1M7Rx7tNdGOHxdurjabGS3grH4v6zUsIYUHtlqWOQ5zQ9Duk1gQ4rXw3MWRmNl
ukhldPMoeW26yu5hrttWpycaeSyupjxb78ld6Y2Jzy46l254NQaQHs/s2yJjh3US1pnK7A2Zfceq
/RPM4KXeG+sMOtKmZbWnE4Tc+/2z3rPq8wPatAQ9gpa1v8xlRIrHP8vIKY+cNleYS67CZxOp2TpH
CvAshPvyB/9+Yrq0YB5wwKuM1b5/TA5ED+O4bDLDnK3RaTt8dWTJbzVUIDLQn5mBGOf1gT2thlt0
DnyM/LG+lRSgqw9GNcYmT0NEFbAFCSlDwjyussRTo1Guj6E5o/DiBcCdzOJn04hkP0cozWxkMmHv
oGjhVqcUf0ZFBWAS+WKjQARiO/jLV/+3svDF88iaLoQIh1coUgqd+HZ/tvDS6lVsFxIU5KPa9g+Y
6uXPFcrstpKZHRRu+5HEMIXp+PgoadlPUqJeI9dFCtWptNBtoJTWmw93seNBEUiWSMfCqEG6lADn
zj94QS0h6MPIMQCI6c1djKJy7XNaxjyvvwptMxSZ6iC/VPrB+VGBZ1+WuP1AovzaXEdKJtRFB1XR
Ka2yoeQ9SU0Wr1CC4njc/zFBqnj0/ugUoAoDQgwVAmpzKhMLYNN6I8BxQx1Pl6CPLBrbylkLpb5t
s6pRYcqFH9XIf2PB8f7zSG2juleRLB3mN5TcHIVXm/eF77le4T+JV7zOOzXXn/B9zVtTS22WGDqc
v2ELh1Kffujg3Q6m4kBtbaLbwEgLLqxVrujlx09Kms1qLLmKMfFmBbJvRLmZ2ZgV1IGwEzxXHOu+
Z44aiAtyNAv21DrIOKzrjTLnYPqaVL7ynhckQ7qP2k4A2H8E01Yi9CHRxsqTB0Fl0q+iDkgYe1zG
uiVBPNj3TgExU7fkC3pA8x45rfe+G0UnrDfZ1w58up/MKi3sy1ZQGIPPRLgsYuaXjeCzk4REmvrG
Yla0hDAvQJHV+25DeOPd9cyQl+YBKjilHn5371R3WT8Tcr9gW0nYKsvVbhEq5ifnI5NRxnSqrmts
pWjet6Lr1BYaZMQwFonLGFXdovvrVDUFeuQkLQEoikEWcWQg1FbQ0yDlcKFWX1OMAkbCl0NqClL8
aKyEwel/bZ0cpch4tG9T1nzgPSAKdtJ4+ipHxtuBMd+09efObC+lfg+QKos9/UPYtIdR6+e6Pwkd
BPC+u3g/gIrepiXxstoaTxhQv1sAJiK6fiyGDMLfPym/ghefhTWHRXPBJwHRrGLNJR7C2zZML0Re
1oG1oETZT9IokiM6jWLO4tucA+8MshI7xq9rav0Ha/OzYmzdG71lvOk7kulP5ZTySA9wPrIzgERT
Uyf1dMXvID8Mcpyt9k9BAImC4T2iiEardiZGkyfsdw52ooqy09lqXSSwgsM5gJOxnIYRD1iQKCaF
1GdMCbh1o/ScmbVhZf0xmghx6mQvz6DvhdTKJsZx9K6rTdG5WPWTUALBh6xre+39FHWxdtat/VxV
UykwiLhuo8bW+8JMfM7WX0PWepfZby08Ald5rk9G4cBS91mOqmBNO73mwixj/6y/OVDogQsGBGqy
gAWPuix8z57ZR1k49ZQhPbaOiG6o2HOjLoaWpKIAtUnBjjO0tJAAJZTvKZrRvJ0l0YcsM2ntPSW8
`pragma protect end_protected
