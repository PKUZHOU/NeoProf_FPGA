// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
Nc6iB/vlMHId/l0ydKAhtXW04DY9MOIA+aGKNovF0WTu6UGSO61YdTtn3PpJUFUe
ELUWSLATmz0radpxgpH3l2YwM4+av9gJvTbYzvut9gL3I9wonhUBdKrdL0wNKgIp
SSCstU5/u7fJ8rF0HxP2nJwiDWvmiLH1S2FRUde8dN8SE+AToQ1O4A==
//pragma protect end_key_block
//pragma protect digest_block
lLN7vw/+Bv+eXklzCCpo9ZXSP/E=
//pragma protect end_digest_block
//pragma protect data_block
OtS00BNp34lsfhoauCcqrzK3eAr9XAIZFqsV1dcoEZqNi3nQJENb1oBblEhIGKMV
FiEZ36AOocIgP4NvjjK5jsNGS7w2GTY/8sY0gx0DjQFK9S8x9gQmKpMLMRQHmOxS
sqZkpN27Gm4HhavWgUf1CsDzJjFI02VicDnJ+UprJ6blrZ2mwDJ6PmOIYiM5/1cJ
WlefV1/G8o2Jei+VpaK2IoQJUMCsJWlEGlp6Kj7p62mDLbW8rdgWJzpVwKix0H+I
qiCsnGtSuJ71s0CCrJGh1vmqseYom3kyGJ4OaHvofXzGNOXWzfDSXXigDhUYn7hc
SniwDJ1hWgBWvBDXod39yq1EOXJkaGit7z2lZScv+2XgYusYIWkqp30IuJe8TavB
I4u/63fXEifra/uboIk9i6lExvFRMvf0ISFAcO8Tz7t+usoai7syGoWMpxb0SYuw
NmZ20GmN148F8DHbadBLNYOi1UYReuIDpjkgTeeougCC9qrfY8R3c+rwuManVgp7
OKbWNpxpXqSbTfjGfb1bzKDkuyEF8B7m0pLelrG4od21gGnQDpgvaNmVJDstCaXQ
KNitbl5doTsNTYmXhf9mkcVHbQF8MsWoCWpfDh84L0PEa69i3JfBJdhZg56qd7MC
ikc7U1WzLe8+mIaMHVjOht1JelvUCzoWMAIEwgWJFslVu31ux6LlCZsNT2xenp2o
cVfrxNKFcFitMawEyfmvifdLr3K1v+dEPpyDXzwNrxTLHSpr2ry2vkJtfS4rIJ/O
c7hd7sNYTt53QfsGjTCPYW3yBV1T+35E50YaXBwcXuX3psl5o/pHUof9EalbDGVg
vRU1zpL6e0gax2Zm57wyopfD5fe/6jSRLt3H1yoA3IqPJIu7YND+NO8o55rBJcKh
LfoJNSDzyiSyodjaLZzdiglzMNcXmPkP2ujspHhOheajs51BML7SScmEDSDSiwJV
WOoOpQ+iWaYkOufLrOMUiC2L85KnP5DjUH0zWWk9FJ6yM6uOYOy7U9qNJdmhNV+E
fntraAtLXnf5RFGc4t4EeQpugrGPbvJNl4V8eSauQ6+rLv8HK4C1ySuPLOsuVLF2
DGgHCRYQ5/0jt5eMLgCu70OOWzig6VoVqat/ytJz+PdQJlA9oaZ1QFZwXz5CJGR2
ygai8TbVEltU7+jvAnot+rSwUgxBkkiocPVv7UcwEjGtm8/6pdu1bNyMgVb9ls8s
AqI7q1jfdaDoFS9/5y7P8a2nNcudy1kd0RuVM+iToVDhWdiJNJZW21cuZRluMPQN
SdUk/0qr74E91AB6YqFKHKSDo7scu8SU6pxcRotLAChhsOoc30cTQbHtXAyqyhAB
wS2+4dDovpcsSyHRScqYH4lSNk7p9zyDZR3d39oFgGTXPADC/MIzU3ookebTlBaE
fNvUzeiwZ1nKoLSxkD3TYcd7e6UXlrV67B4cg8Nl7xJbshzlbfHTdve8sSEKrG9e
0o94cLt9+SDoo/qkj3Fopr5gyKH9JP5YjfCf3bacutRXIFVp/7hbXQokwH1NTgUs
y0ROebnGk9i+tnu7CRMQbWXg4TQe29vavpLgF7Ar9Kby/aO59JsROEY0OQZkHk+r
2JzB23AUi8fY0UxwWV58RdQGsBQ1BHlMLSbsvtAgfv/kJJEV1hluyuejCM8nhCPM
bhagH+iZOwIyeGPA7lPsoa+WgMc8PqOU95onzOmhbf5XVgQGp9pjwMlbRbufTnW+
vUJTYvVIUaKN1wT+/cISrsWj2qantZNfN0PZCbm/Kdvg61tK2UuApaegagKOw661
TdAuknwWCkrOXqIAo7ZjIuEOYXBRVeAOd2gCtKcCBjwAK/K2tmOiA9X92H7VqkQ2
+poyEbi48bLT9f0GaiG8jbcYJ0QnwDOqWS9S+0uTEDGFjYBCa4RfPma1LMt1askI
n+cILeTTnUzS+nnt7OyxwZ9ydABIZRlbY7Do6jaOvb1vnbYk34ldKNYShCmwMEcv
lmeo1rjbeckrnSxap0kDUaWl922vNwrQMIuhUig/TgahYkAzGNE4eL7Z2/W75i8g
pVa8lMeznfatybpxD+RiOPrDHMN50xwsMDV/2TtkGVTae4E/4QqJ+QdKTOZe4VqA
7GK4z47v7QUIh5l+DSAKJsu8p1CF71WOETqTzKUq99Yuv+5prUspc+0pKv1Eo1tT
hfXW5na7bzsNCGaElGa/AhjWSy5YrXoe0r8Ft6lQN2pjOD0KDwYHNgGJNGJ2Z1kx
8mbiP0mptL2Rz3Q3VlJlVFv2fmZdxxDdk30SN8Ls7JT5QO7Zn3uUGo+Y7tC39UBk
tA/iZQfG/hlE5/DuHFxlsz2cSKWkTdq9XzhWgVR+mnUH4zEV0KJIetqsGP7Iio2t
3AHjk0MWwuk9kqm5BAWUf2auiAHEjlnpivcbS9fs/AAVJ7M1MwKuc0pA/Dq0bMhG
D81/oZEL1zxWPNr6UCrTF4XdTUnNPcgKpqDW5xOGJf2fDfid6AkruaMRSWAh4sqx
htVjWclEIlmy75ttKAmrI2mCOWLCSgL5UNV+rP/o6OkIHLUKckMg4vFR9JDtBfET
CU8ugE8tPgsmoNK970M+todkFKeRUUGksRy+Q19z0vfLuVtw2WTVutOrpQBnGBVW
TBoeztg3YtpINOuvl9A+t0tHmgKhlbKcfXxkG8NAWjJiKcup0A172XMvUr1u060M
tPpwRv+AxGFsT46c+vzyIW82mQHxtg25P8eBfSloypui7fneG6YgJPAbcJEyZzt9
lb4Xyrg7hUOvt+qEMgs0F1uxsnTR5HGDGOEpdkEnqTg4dwu2MDuWx37U90VwwSVG
wWxV0d2bd0Hp3kHT8rDYZD/IEKY/Pq5tCeBtedd92O06/oGXlva3IBKSi9EBqB1d
6PKy8N7OVvD0mdgHIBBV1lzJznGlgrG82CueltQc/a2UA3X/73kHM23hDLUcEcwX
d+lCmi+Hnmnbz5ZeDBKn3j0pmPvXg3C2+5x4OfYXxTDGQnSXRx1PyyYF1jWhTLiy
C4rCsOneXMaoHXCiaKorvNrczkcAYoHm2PcNy3mFuLKrsrRfXUX7N6kiQE/MvVVL
5IHf2NgWfz6L8i7it77qu5lDQeAXKLpDa/fStUIW2YOL1s/C56cehNhq2ZlvZsnw
cKmiMNYwJT5EwFD0PT7/1xJzva7/7XdRpvcy2oWDQ7KVzQ7wNPcZN/mbrgiVcPm4
FjTXnwAvJFyLQbNACoai6VaQaHIPNsKatDCDRNaliELYXF/x7tlFnSSTveFWGhBq
ue7CpHAfYyJV083DlIzJGrQuyOggUWFfB0+jL1aKuZgLf1w0QTOvAzy9uCHfYDVF
A8IoGzTqYY/ff5L8cAO2uyPplTxESnQ5JGmkvv7Qz0FFHj9f1v+Vz+wb9DFFvPOs
n+HyIF4Gy7b4tXR3N/EqWZam0QG9v1LqaLu/GvJ7iCEh/61D5D9dZsrPtTtNJ42T
7ixAHDcfYp7eU5OQFrxjjw73o8IKNqKI4S8AWBKC1nQMJmTfVchwjW+ds4+yTyAv
QzU+cG+spZBPBBUM7CM3eSicY+5LubIVVKw3lJ0RXNMMyrjP6aNj8LpDxnO9Hulf
lxC6PKEO5z9d1IfZ3RcuuvdwU4X/wdB7QglMap6Y3HnuEuJJ5GbPJaNypU649cJw
Eo+WhoQUl4SGe+F/yq+H2HiDVZ5dGGwBN7Me31yGviqBT4Nj8fBjTePy9BtgPTti
h3cfhjnO20kvTjiwjY0/iRlg6Xp+ZvsGvH8DqPhnHqjM0VHiBiZMPFFjtt6z8or0
4rMtbpUzMEEyMq2esBLdPVaxm9kwkYgHFDVYe5sHKNl8aiIvEXS/tIr6Q8UbnJMX
FEQVfuWAOeESx1xLlAisoEMAMTQBYp5tV9NgJarp05CN/FwkG73RSIqbB6sEfIgl
yHJ9DVn/ggpaE7Ekmpp7nmoiZuSWU5t/uH9T7glwO7dq6GK2WWZKvHpQtmOP5bgj
NX1DKInrOeGE7/USfOflSBmDBsgD+CUUTbLq71B3kEkd5Chs8Ea3hKbaoLaY+Ci4
nB4NcNoEuoei8x9WmnOAoNXgWrwO8Cx+3yJu/3YCyhLh3LNCWwV+OKMZgK8Ab0s6
k+HeGpPmQy6EAxz5otUXX9KVKRWXGSO90+WIZl+VliGhAJdkoqT4FaVh35DMoqzh
vJCqukDw8XNcoRDRFATovJIGG0GrePRaLrbJ3tvnrT30qb0gVvZk0ziMvqMeOtBj
/YjaboEshhQ+oYPFZMp1igFiupuqEi9e2NYjguzrr8M/5FnTt53NI/QV6yp7wGR2
2lROl9AqW0azKdUMEqWZZzDMz1ol9Rb2zERNKKxec7yCdWKUshjmD6JC+uHWGzbc
Bj0o1jKmCNI1jKQDc76R56V3Db2WCBc4oXD4yR0huvKNXh/iuwRUApw2FBhjRb6T
s2Fa3T05q+s8xnfdgVKQYS146w16UKC11qu/xd1c6h7RT25q72YkrFHZYtfdtTyZ
9LeTxDbNMz9ASqQnoC5bnS7UAtPRrrE0LPAH7UcHvNvaLBvJ22UtiMpNrCCSmOsh
S1BWyR/XJRK7byVXYy9izaxgBxED1WRLLfsQoiE8lE0QbmFM9OCGG0ObpjOMY360
RjtY5LvX1FmPsOOLn08F3tSgNG7wXuxRG1AZ/hWrlh7qdZRPMWQ7aSU38i6HRHrx
e3Zg2GKRewEVhUJN35D8SkTK/aLskFlMp3eOO0jyUhQsIWCDBSA1HbWz/nDpaaRe
ZCjkgCm6D/9Qrws/fbWsPv6FdV7mvtUA/P4YUq1M4NP++7SsbmHdqrR4nx1o3sXa
sGy2rOhSpWsSJfUMIg/btPOv2c4aiqvF9lo/YPu/0MNyXMS7pUNPbdd++EfcJuJk
g4Wz4ZhjQTZpqAGen/8BukDTSM4/FPH7VbsviK9dgwiM5pm5CrnqKhnR5JlYZuyA
hN5UuLRGAGdqzqOy9d0RpqtWGQiVq2hUCiifiGj5UAOYXGvPta8V2uPsUPAM+2QH
Pp0nxtmhB6CWk9ZMTFkIBojtZYLOpaKrEnTBuikm+/F2Ny6vb2H5e7d25HSlZmRO
Y2F36krG+Zd46cuV8DaJgtA9eCHwl2Jghgv3AztDp2Q6FScHBNJ3I6F+P3wBRIus
szrfdrJGZjNfQKkWi+CpWdzQdeZ20ZcdyLe089qx8AabtideZEuLjly/I71eGkBD
v1IETnEpUpJfVhom/y/OItx3omZvFF6n0MUJ2ORw4bLtmqq1KPcghlgWUO9Zjh1b
0JjsxXUF50Uo8ODRgNLSmzzqRJrJ1wtHibbbmKzqrv9YE8LBQrkb0qvl16oLlkfF
1854vu7V25UaxGsROsvVd294OWfMilTEarMtXMxPFjWonVX17jhrxjjorNuwQ/XN
1gbxlYoJCphte1gaNiInl4ByYYRjJCF8opTBza/JDdPRCb9tGs1ucR2N30qfMeKo
6YCo+/QT8h/C6p7qB4qdrRzVV5USVAR7ctp8z+W4ukJ+D7gThkEc6mCALAgYM4m1
DMQCppDFkfelALUN1yQKn0BY6gldne5x3190EZ0Z4P1FK4cWJ1ydWdMx7WNbJuDz
Hd+IkQpANCxjuFDCVgWwIA0nx5XlSPi5yLL/K3IrNE1cPRp7JkKBrdCh6gZr1BW4
hFPwsUAjUWJD1kJKmHggSVYvC41J0hzenq9NwLeh7f/F6USSF6eZm9ciiyC8k9yF
859bQGTHDQRslsaZyuoaZdKlnRkvEa83j0L7Z3oa+0D8oEsxCQ3Xlr6KAaOGPLtG
D2d93BLwEs30gmQWn4Dn6+P+WXe6Ck2lH04vMjfSbOSv1VDA7BQ2HSydNho7o1y5
j90JCAEp0CrmKkmTQLNNbq1Rtz2zmrPf7uSnBfGHQAq2Rvhrq7pc2kppY5m5aTxe
Erb1zcky6HA5YcBcDU1K0MpAmA2Y4MPyn+NVHzIBQvqevQUisFpJSoKhNHKvPUSo
O+zxu0jR80tLuAyICeul+63NsE0dJwkZYLE83JrHWjzNYDzxBOMkkWAdZcxVuqBR
w/5Mnxyb/ZpcgkZO6PqaOLvvNq9LER1YmcbCXAgtsF2Nxf4PjYGik0OKU01uZksM
6f3jGUQ1N4zQfjiOfIDRBCU9weL6vGs2aI2RQugnuTPoysEbVRpgCsN6NM8juNkn
c51MgbqDQ1OmtmWxOkZaee7cbd3t6+EsJw9ezrtEYVH8/Fd9UIfuqe3EZbkWkwpq
XO+zHOGpwxRoaurbYlNA4rsJExdc2eCPu7mnaazr4P5EO6RSPLGZgL6ZIVYvudIz
7TTnWdZEZ1sw7GN36RKAHqg6+43ubAq9mSm+yMitgNiireWTlNbkhjU9EiwlrHcy
iIqaDg36MradFxpvak/y70G2hc0U9t8JFql2L9nQPcFx8XZsUXr6ZpA9WB3A0VbI
DGsJVm8bkCbKP36X82h+VbBydtXo+rathyxEmZ+bIx7CI4+pW6Oba1SvAeGsYdRs
dRJSN8bGtYsrrr8wpHfG11b8MejlWjbqJ/1v/NINaYSSLTN+6iJy/TpcFOhZUwiY
Rk1dspQ4Km40LuemFaz078jEZLv6Jg4s8LnSo1cCeXMsIzJJIpLqm/pxzsNyCYb4
P4ghcR9PafXF1ppw5g/EgB+hLdKHjdM7nIwvfzrAtLCbXHFHMBloxKZ+amHbhZ2C
ufno3oaMOCXFJxRfV7oD6aviQRMSpksX068zYey+jqpwd6PJE72FhMAsFgZbu2Fa
IsZ3XTZExpMt3liJtDuWsWusA6F0UP2UOUPJpPsRJYBDyb1EkhFr5hFCS+dPyiPx
nArsBS6DrQ5mvvUHDckfmeJ7b89I63scuhYSB0nMxNPBQTf+GqHDLkHoSR9TV/2g
8SIWux/nPFJe6910B/043B0eVilqwLARXDiDNkKcjivbCjwykICfkYErwknq/uhj
elOnoSMdlHbGGCKSmh8rPobSmQJFpcT+r1tjHmK162AfjwDM4Tz/MlzA9pil57Uf
r0zdWtTRC91tVYblNcyegOSER755G6I/quGZI48Q9NSNSikSrEUnv2ACODODLl9z
GSPE0iRlb2uF9kUkz2B6p25g0DWAM89Ia4Xjx1M7YAUrrlTClRZMILt/jtk0smdV
IMmYjSILpbB2ejtitGjmBsVjrPLKzLCeAHj8hwpqsiqBWiDWYNBYnSqchMRqUksG
ihxZ4xfdXBGrZgJQ47hIMwCH18wr9kZiw0eoegVxT/W1zevFGM96OfQbpBLqZoE+
Pc/1yRu28NcRiuYQr2cSPzdacuo0ygUaYjthX5bQIOEQCKsQbakjiDSSnI6alTpi
JtXqwAP8+IXc+ndEamjKfMLLTMPcdemq7wlddgUKdPI9pDV3LSyDQI8OVRl5DchJ
Evj6aJMk1mMB0kw1jfky6vRuPbM/e0m6nc08TbLZjTihZeZRQvX+PuJtA8cQj8Nw
27CC5vtzBrKsprQ5d4/lI/lzxc4wWRBnLzywtffNYJXwj2odmrhGU/20N/4hHkRB
Rdjwq3qzhwIo68/OyG5ltkX4K2j28kw7lQJoO2Rrdc6djwG5q+aEX3ddxNXkX7oj
sDRQxyNI7eUsyXXxI7YeEVY28AXeE378Z0heFTGjK4/tHcoHxVkAS833V4DtlWDG
ApCZejl5D1C4UrdpfXt1i7HBXxnwuZ37ZSgHSM1G5oHF1f0Zx42S2M2bkTquXhOh
Bzu7T2OIwhg6p0gAikw+fiDCRyDlVoMeencqMmFVb9NXWC4QmpYS6Qr7hs4JwBbZ
FrJgAj4MBph6kQNgrRYtBhhuXRP00Fm8O9u06fR95FfM3Pia2GZJMQqocuK4AZrA
04XqOuChpR3Yt2gOsxq82vlIa8wpYRZ5VNYmQ3tvFe1vgl4WJ1RHKdbrsSvFLre4
xn+jysDnxHywk7FaG/b7lRI8HlBWObom1zHLwfTBIKK2QmQgasvdqAzZNj8mTRd3
NnSCWgK+1rQB7yroghztUkxEwRDo1Vhm6OGX1uFTN9/So3tv9jeOIMpWo4iKgnCI
DExuzqy6RP3GfTdxFygf7T/WGj4C4+9cArNWgCZrDfiEZ829xRM30lNZYJmPt1qv
4hIZG3ziK9ZR2Xa529BJT+4kXy5meAzgfukbxsMzfa4Hn0hu+O6LS4FzmomAkhhZ
7PTLeKiRoBGPYmyXJob7zqb5aEDpTzSYnaDAx6yGtuPcD0V7pwYrZfVUFeKRphC4
XuI6Xzu1Q6nRb4KmyvU8sxTbSSL52LHynztEtrhYMBE+D19uOpxsSiz8MjHjMfBC
8cl3812chs/9YiOhSBbFPNr95Cyg5Eof0vReYoCxTHrdFsSIRRmlds6K1y5TE3Yf
CTnau9imdbmDAtBckUunCfcTtM8s6rfHSSY52lnW23oLe7r6lmats5khKFuWdJFF
KqkB0LmiyRp3MmCUqEtikJtv5jaHIQbwVtLcgYn/ybMmJFXO/j6akeUMCu5lj76K
Aj7T6+52+kszqBWpxTfEp58FbHll5uSLcon05K61sFKxuWOEGCnTlt1QcLISMo13
8P1pvoNvx5H4EHiXA4CqvsYRMFlf3Tt7EU+QJZizhhajJmWA5t7whmVhHM0yA/T+
Q+E1ll7mIXjT2TfK1crMqcIv7W6XJxwKgyFzmMDxZ+OnyVWBLQl6w7vy0eYpflNY
uP5sRB6ATcElW6wxKgPSYMRfeycdHuk9CtpJM1bsnW/TjFaK+S1eiVLsP+SfDRqx
BVoeJdagq0HE0VYxr8eMVnbsMrA+fMFQvNRe0dSlIUdM5a6xXQ09JguacDJZwXMW
7VZ6NwETXLSLq/T0TIZl2A0/44Zvtke/+/KHG7ReaCLQsefIjlTNJY8dGqUYTsmi
n31A002F+FY7YbUU4K0tClOLjbgy5jS+ydEurRHuEvNvzuJRn+I5lPLGlTi9TiCh
Igxli7Qn3gvj00K2HRcnRP6ZMtWIsHFkcW/JDH5GGlrBKeKKAUGjhHqckKPCtyAd
hCFr7w+RdEjC5p9tcrBcGkyLYYzPoNakPSocy6uCtWK5Xk3uY3wQXh89hBvtGG5Z
Rvq5wcbLc/ymA87hNZ22mcIpDTfWPcW5ACuOpQZFRTfWpFiFwjUSTrts0BypLV+U
oPGvV91tnFc21Q/x3O/fGtzdCVyxTQZkO0jRSnODWYetfBmm0GrQwCl9x96gvFL/
aGYxO6KCrDoAG6zlzjvZ8xdqCd4FZtkPK46b/85kpuXDxh9tvGvMMmQPGJ8+cx9O
BBAdENQJqq5tX/pY856ETCti5ssIKa77pqMe8d9viVcakeek8AUfFVQiunVN7FZO
4Uzasb+UBFSiaPN7+Su3Fcqw2kKpDTDXy2nNGTL8Cc8Hu1JLU8YxLtYd6HfIu0YK
4IVngDkE13RZnHH6ac29139it56+C8Lb+CVUXL/ziLJvOUzUWpfMtSgM1wbw9LFD
/RSBicj+eaGtc83ZYLPSrFVd0bIZIVMFwx8wnKfOM2UC0WoRXxSXISzVGFXVFD9/
TkB4EymrWuavS4D02fpfT79E72vSJ8ez2xqtePjZPVZtU5hA/aYWM+sZOWc6Qm6n
Fx4/WtICfAfw5e+5NB82PFTPO/P1L4bvAPv7jhoRc69Nw1sB2JRimet37BhhqCZ5
9URnV4ofOizuk5X5X2xURoJCsJE8uP9sWXvCluNfVh6MgIVK8ule+kvw/xgtYToY
2qXMT9k9Rbfs7TvF9zSAlqs+UOVK/FH9vd7lxST6835a7sWAeSwvdY16iw15t/H/
LcY56sQvzJKbUIaV50SA9ab3TJUHT7LLln9Q6NmKaHIopZyr18kUYYaRX7nBqyV9
voK6SHEmTpsf4iAZuBzBk2TjTkYxXjPnGcgfEVVgZRJESeDn1nQKo4+b/MdVjhPI
5fghAM6mfERDhNMIBmUInDTq6hdTHNY3PfjyWSglhPkx7rvmCPLcN2VoucLZiZPS
71nv30htdrKmE419ntnKGLGwlyiv9tgC4LiDQDLe0eyLXjVEP4JujcxVALFvRds+
WMO9OP7TK6a/SUa8hxtZ0rejD/SY1UdkFjum4xMCguAJb3C+C7zZhn7WEsk03Fb0
/hGOLxvHVYh9BkaIcLvQijrELif8rUQA2UIo5ars+SPX/VuZd+S9eDXMuuzqwkIh
4/XWWxul2O4pxJxqB1hi4xBUpXS5F5OIeD4i+kh4dMARwxV1L+71EQaIO5wlp2AZ
ishhpWIH0RFOzn68GizWKZHdSc9mFu1jPCRZJanJ0h/jUjzvYYSrcOPeRLG44+LF
2CpovBu0BCxL1gH3AEULD7Z7NSKgk9aHOiW4hj+qfhDOnKi1V/NbGuOS3N3wIbc3
tNWrooNHytLgRGS7bOby8MMBO8PDeN3Hd6hyE0l2ukI6wgUoeDWVzZNsi55Pvx0H
1nEdQ+BKmIdFkKIKOE3+sMccSRpKmObVRy2WOaS6WxgNrmTmmFCTsfv55zkXQi13
W0jl/mRr11jzuyfFAbxN5qdE/8+UeBEk1CpJbAbi0PX4I8QcZvxZ9V9KEdUSfD30
xLje9aW7FqzUoXsJwiV+EVXwspRIiTc6xJbyfHrG4amnR03P5s6QWbiaEznvcpHm
t6Tf17k92wCxvmgD1+bp6vMijPSZ3xdQ1gTDinRjC9ayOC77nMz1ypammw9VYhzz
qrONfAMYluMMiM4hqhvhb5e+hRUw32Z/KMQ285fKLf1fbJABn6KPVN1c6s34QWiK
swV1FrVgG73fp/D4nB8BLHZvL5MtI9MkHuLe3yk8mInpj3nr2WO7TdbcLzu1RlBL
+aDeXU9sZ1V6m339NYttnroG6Bjh6MgWz6Gr5Upu9ZxRP6xd1dmJncNkOhZsC+s4
TQezpFI9YeN4QqapS/JpZJQDA7i5k44k7zmjy6HllQdqYPKTiUL0Ibc//TgxMvae
UEVrhIgXeKOvEZ/G5wHQEzyDP62k7vMp310aDY4XJtUNDSJIXw7fhRHBiCQTCqRj
8CYUOfruWgodsJOCWAMafQgbSSvjdhQekGRegi4QfnnN0CzW3XD5c7sRJqU6LqDS
/NyTTByVM5e0rWBxV7Pwo3GnwI4ZnBrNl92CgpW21xd0ZCgMCCvb8HGnQvYzZoA1
KX/xrYqkfH46ZWxQxLCVT/u7a+8uHX0AfT8SzytazfIBynzS8UkSiMj+TxtAbEc6
5M4CftUgXIVW+RfT2R4a2Q9BCV9O65S1t8PxcQuZ+bU04jBVaImtl5vydFmpswGW
NWvjPwdi3Dw7F8fjAdsWNFxrZwmzNF0APYS6Gn1fQ1I3NJlhWMgresnntMD/3ae6
GoOPa/y7lA1zQIAlqALFcHAFBZgkE1BSWrC9gNP/Pyo1FKSPBhH+BdVd79lWAEjz
HUBHKj5H2B2OmFTtoiktqb/JcM1/DPJxiEDIVBevSc4vz3bU9k16YMVdzyPq3Lvs
IzQSDWe7phsZY8O6eNJTJal0s6IdgFNTcadG1DAFQspe6+HhEAuN/VEFg0uw8SmL
ZhLV45Tq39+f3U6RG7u7CFdbtlbPShmiCNrqdLa+L/U4O+756JpT2nf7/k04FhD+
JO8ap2nTnSwkfIzWsJrgiDMvXlHdrjSg4b/tVruQtZLJwtu3I18zvf0SrAlWjjuU
umgPjGkEGVK1gJ2gGuiVlOAvw+i5y9p21/mgQCr9HHy6ypd+ffxP5Jn/U8ygrgwm
3m/6m8RzjCY95TUNzxTPc45hcEt2NpQh0jsy626UJzNbQXB90fKfjMnpSsJiyXeL
7o6fHhR7v2TSvcCysbSgTXs0yttVeOMG4rtWEaprRBUPOO4GftVIhJVnmciM5DnZ
hP9ZqqzHcZWzdGaFgtIium5BlMqnoono3rWyfocNcdDyGACeNeA86c6dUUyqAC3y
/yQfdXGiEMd/uEqwEw1IjDAjVe1dGRisimN8cNa5HAsSGSINoeooel3x/y9J5vH1
rO2OpQHC3L6B6VCG9fr2Iog+nqWAPWXgsU86N2rS12D6ksxkv0C9CajRl/Pg75ih
hIoDt+5JBv59Je6T6dozPT2k8C8lIDZiVfbxVoj78T413zo9y95LUn1IlAleU5FG
YrXgbcy4ZrDOTykisVZBM7fWh4urXTGlhR+3OpwEXzJOJarvSlFE/QrLZ2iFoUkW
5zpvtDGP09hLCK/lHI0anzsZrqvnn1T14DomAv70G+L2Q6H3jSQGm4ibvnPH4GaC
yB9r5nW8BxUk9Aipiw9zq3ncYLlvZxqISaT3V152NtgogwwfUaYS6imc/3d6Gu0z
zkC/wm4V2lEXyai3Vpmf51r/RYz3XYG8i3EUsUFFk0oHymCd46/G0FB40YxZb8Sy
RN8WGNsC8Ov73gHhox3YETN8EnTzEgo8+/Owg40Ab1J/4t/zZuK49KtFp5vJ5Zrz
pK0AgDuIxZWLqSB3BURx9Be7+Weuj+aOKO+VRtVQa+pZa7nUzaFp3roHGSCPFETj
Mn11TVDF7z6KqngAufI2hubgoh/csQMtHFaPH6ffH2j4O2yroNYX0P4L+L43m1OU
igjaplqtc9gjtcaXHJMS1PwPi0d8PBMLXJPtkTA2AASuWet2ukvAvjHOW1825H1D
n6bxAgbMhD1E17jyJhUyf++Iudw+qDv+VrXQjY5kiBCDv90cjtp75a7i8W6ANxbM
Q2PVYQ8SbOwm6giBKhEPiHZdSw/FUjuzn5tyWu6VYqAX1hYgME5j7qcSg3PoUJAF
8MAIK2vFEcHoNK2ow+MddfDs9AAhtpWukOyQUANy+XXK/v4aSEfYk2a9Nr/m3kOl
VQkgaYfhxTqgmn51iJnZ3fSJZNmO8+OppUSMncIDJtuUVvnZf6y2ajSjxkeDlvef
JhO8j24gepyaEImM6ITubi6/CYodvOZJ0M+t9iGAOtDxdovAQEzz2kBwDD2/RF+S
wJO/NbXkKTC7tmmPEXzX3BUbV6f79MwkMRDJk/xpJyTYzlU0EDYD5BmuQjanvkiz
0wMomcGum1Ot50gJ7uyoZnzDWKsEyRvSORxZVcU+vYMQs8dcdmsAzoC5z0eHI3hR
orNm2gLCHKuufbXqMcWYDdTAhS4COgDaQBU0pf1gDVh3yiOzjx4cZnYARepz2Fxt
i5ZNfthrfNQBTmOYS2dFLRx37SGuIux4liQ5i1oZJnzds+GG/8nU4lJ6R3viLXJT
UVuX/P8GYo+ZrpTrLg7EUKuHlANdjUhndd9/dpQgiFLwDj7noxt8KT/66zFl0Vd+
zdgRRReK7QyqrcfIQPqzD17qt+Zbbret417Gr4eIW+XCbkYT9iQYofPLChWAoVKe
alq3Yv7KBjeOsSVi6SytLiDLq2enb0fuf9+jepMaHFoeybcTeHkxmEGzIOGC2YT2
vlO+WmTYO4T3cL6PRDZn5Z4NitdnzfxO71gd4eBmBMTyz2ZYNVkIYfAIhIFH4sDK
fGwDK9lNJvoDjSdcrBo9TJzat5UJb3BMeuun7nBtfgDljOz+rVpAZ//o1wOSxbkY
XtZDyyFtz6x48sU6oJZhizzg/QmfgHIb3tt15iTa2Vj4hiVStM+A14urYRZF/NjH
izxGZDBreDEvwZSPIgv2yBLqNGKvtLz7jbmxpPMg3LtywSiNGv+o3UWtViD+zEsn
BGSXwmbxK93McCZ4+BvJKBy3R+TzX2joJeCKFZqY85IcqGS2XtJAU0+u55qNMMXc
V9v8CgQRYhoaSCKZXd6H9+mN0eFY0a7xGDOkitc1Qab+u3iPqr4K9wnIqzXAAfQo
t82BoGmTkt/5mLY0mTGvT4Y5d78dg9TN7td0uEQMOlu0TUQ+RfuJOBV2dxlspahf
FaMZK+6tdMVZZNCN3XOhnA74A+0ZeMOFFh0zw0/cHgOeOrViConiZH8AUyOMHn4Q
APVg9NnIXvwFKOZlRbsBbQYLWF/t2o19Upva9cnJ5/ghucOTH9Kl8RDG86yeM9Gs
tA25w9HyUkmdCMzgg2FuaBL4yC82CvH/3N+pb3aAAEFBX1rQTvRRHbEvfqyQxwr0
plFvVNrh83JvznHx0PzvrjQbSH+f0Xevnw/1b41H0Vcwnbf8vXjKcLE/JMN19H22
rOXEg9OOfo82/K/gfPUoHySnevzBecmvOfvzoGbulKsePPJ9YzMQ2GV0+tc3h3Oi
CSj/9GjQEMXrF1qAzDuS8Jh+zZGGaRdiRY9L5uZwbB1ZdNJWlBWHxl4ZoLXhAqFC
SXMSEmXBpezzEKrMDYGVlm63GlxWarTZY+pVrXrZQ0JcXjHfDYrCSRsV+AGAN3HS
3djx0ejPkzH+dKqGbsPPBQr1T4XDCEOMepcq6q1nM+9f2SYRq5vNlbQZMg4KSFV/
xlkxCA/AsMOEEImuthKvsqqB8CNrLzdSHo3ediAoc0wJ9R0MwyfWjzG90cuHqFMX
K5DutI336vu5kqSCFcJh3paAQqqGsK89u6tkcYawnCakYrVQA4aobLXx6rEbzuKE
8RFu/G0SMFFQ+YWAF7Fmin1I8vc73u1hS4l6dPdxl8k/GIMGHZjiV+LGJL/D4gYB
3ekkgX0B84bqTX1RQul3r9+oAx8M0W9S8E+07UhbJOwyhp1l6U91TPHzSeYNHmQy
KtFSjwMMOO0SGoBhnIhufN04RxohZLhrmk3uEak1Ygm1ckH7Cn7S19yUuuzIc70h
Rq4aksiPeXZTq9YsZ6a+Dag8mGRe5N4w3qZhvfM+5LjKJlbJwe4hvOK7KpQqK1Uz
gS8WXTSwRh8n9P6PXCx5D/846CVsgvz3m1Jms/UakcF8AZhlESiy8E+uJ6uS/oOq
0V8v6F68nTLGYpudLrDRNtznSG8J5ru3yHXiZye66/ivkhaDL1kiAjfrk9vd12WZ
8hcU8y94i241UpeDwboe8IyKDnq20o2ijgA8btGMDLP75He79mk3MXvXNhFTzYZr
BnNo3JUz19CNsZqoRCfTPCVmzPy2rTlG+G5w2vTnfOl1yxWO6/WST0XjuU3VkvJW
scC4hexIbZN3JXggLsjI5mo/hJVWjtI4yvJW13TtZGBOeAUZzs+pmFiD0hnJXlsK
53nFxZvSijWvb0TOR9TTjitygbh/cwT4Ws5QRAnV3QUlbbYvMGw5v6iblCIvFie1
DgRT/xYKs2WOHHe9JgHdxH6Id+Iv3gKRPF/+TCLSYmV1GN70iINf9szCsaGBgeO5
F60kq7f5kITqgvr86R423jauiL+KtqyZXM+gFNo3SpBbuKeUvlnOJbbtshpbaPNB
NwIcslRtJuz5AAUNsS8Pm9YuvTIG990ff6vhdJzpuI1qLuCiIEuxXW8VsmC2qKcL
kAIJJ6IrXbHrzXX6QiQow7sOEsRz9s1bhR6PYRe7hplo8vGlGL1Ml4JhZRwgYzsD
amxmTu1kn5DPhhFY+MWXs4EK3c76rAjaAG3hZRWR2OliWPU6UtZ3hOgieT/0/AGx
6W993I/UrQzVZ3HObktKfg9A0o7m48/kKr0bkvx7DZ+hZ7PLszO1VuPp/zUebVnR
e7OcOuaGfbZxnNrx2xpe7RcelZp2dR1uWUcFzbh36UHAEskeoq9Xf128ibWR5xVN
FjsOl5QAAbw2E7mbyAqmyjXwZB8RfXrc+BZUHrp+on/BoAmnSDlEE3iPN3j2lA8A
IMe9jFNMsh37p9Rj+Atm3Cu1dZBG4/Or017rO+5KoTzhEFOEm8qinov2gUsQoTN1
9Fnv2JerSWs6dpf17qtAB/+UpZFPB2QUqJTQeElXwU56p6Kn+lkzd+4cHBQ7H3gb
U4uoaMZDAYpHv/AYK8izqVIH/O0GO0wUX7cH/iS0aSMl2QhyYJl8luAxzHhLhaJC
hTnzPDrkMiDD82c8pmqhsGbuXDcI92whfYstXa/qolUSzPxMtYFY0I1ufjOshlmY
0TqdMTCS1Ve63QuTLnL4N1prIIncVwJvsmbMj+bx6HWgyq5OdrM81lJbbPk6e6Fu
LP8mV5Dmxq6V6hs4DpOCPCSyJSQcXnyKveJJpdSSTcK7rSpz7P5TiR0PcUasRVil
lyc86n2obzYcORXExYlR4lvk51bqTanax0H865oGAcMuQ9ZJJ5FS+0b8STgHA3ac
21lD67pAscWlgksBsu1gM0fKUzYtaR7QHDRCD1JuGf1LiDg687SDxkbXhqPvaJ7v
0e7CPMZ7jttb54Cpowz5s/YNPHpO99Jl7fv+tMDsbZ0sErIOyB3KS421vlUmy/AE
L5tyEl1zL/vt6z9pwUhoZFL5Xj/Gi7K8rtr/CaVFtToc5wKAJCjsesR7SH3biLZa
7FrNHvv/mrnn+dNWddSt4gt7wlKgkFEzwheTSqUWlWhIadrVbeVtxbGIAg4DyVz0
n4g9bIpxOx/fdMgOGY+xMVIbXHm0xxv3B/BZBp6g7OjXRKCvRpZJwj4rKvMCIDUb
15PGYL+ToZFojQhz1Cx4UAIVUwEFN8efJ6CTGvu0kNc/WU9ZM58v8rtD5cSwyf1J
TXegrPHz6Y1MzAXpaleGgBuz9qpHrwkG39Rrwu5T3VTdvdCEqgwZzy5xdtw4oZa5
Zzkop4hGiZqceMJhybtmvmeCXHOuSbAyV8vxA/qexeoLZNCVOGP4P5BhnO6O7m8h
E2ErY61DjPB+aoVz6FvvX4lsoAcYl/Z70mUDTrHVn5zLjZpL25CT5xGZq+58FEh1
v9wWCjcAOUXSzO+9wLw0WvhCignSjjN0cd91spJOVspXSPT/HRQkY0JmB6W+zMxS
fq8ajXEyfkCFnl97fjp2tgZ/8dBBiFxFjpcZiXEZDsbEwiNaxKOg1upkMVJBNylI
RPhzmsaQwBnve+6NX3aAFLgW2afzkVpWZe0crhE4oNUgwcoBGDpFHj2apGsxBX4I
MHPJuwYijQlW8TcdRQjgr4RY3TjhgCsD3UaAX2fJ+ZNOOP58f8fipNGZgZ3pheKd
BWIoRc3Y7kC61thEuwyz9D+drVcl6xrUgquQZ5FT7Dvq7vRImfE/Tj77Ei0KuMqV
VGsVB3sqGeMcgKodyu2bnRl0jqkJKJsaRpT5316kUx0bOvBTEWg7PKZ4l0l6rwrT
og6xQLofWBcFsNYV4gFes7nj1VgWcZbZzEXIv7KSIfXOJctsrOhgFwm8ltdrTKIU
lnm4p5UrvpZ1LlEbYOLnVvJi8RT/rfrkYqc7KbKKTL02xag0uVIz6Qke4hQRkNyr
kylYwRcfXvHzpG0byalsbbRW0YOM6NIQMUXTGwUPLTyU1txLNxo7HEIJHf67cVtB
9r4zWWZoucHPnmj+csmLY+kywuAIGkBZ/cEAY7/9NzlWRy7IhfjeAWEJ/rvqiLm8
WYepsLAH9YTaHnuRrVNEQOJBYWK+Fy1stfVGZVDMPV4cYGXkExVO3f2YapNly+r4
1jjQQdKmKo64yfAGp8ybwhP+Dth3aE1bhmTf0IpG4WByoKd8mH2fxCvNaIPNDkw5
lcMlqFEtLJhf4CwJHrxiRomTjuHOPDoHaIzbc84jJHdxXdUxoW6K2F5rej9xWwRE
s74DlgdeuTgRSiXOpPNCHxAVQT/T6mY3AUj4J7c8No4WjZ9JmRubEkOEIvUfHTxp
UI1EgCeOyOLEeTAMMOYqifS6L6ekWtasTXpDh4aQM7ie1sRGvutWKLgn1FSZWiSl
jiga2dfRYFKpIftsvoS+qx349B1HPxRULyUYvapQ9yN+ZXL7tXxMpc7KA+0CgMgj
Bj5/pch1Ifsk+95G7U6YchnVSOBqN+7Iv0wNoxNztww8QorigmAF8zqi21LJa5DL
xDbQlHNLshb6bfPfc2iEFSFd9gAlznR+OqO8L+dnthtKb9agUWe00nsa/EF7/gmp
ILVGR0E3g3/HaGzGa8z1x7CLx80BcIM5+zcspYRTjo9r4oTbzO+o20MaPDlmr4rK
pl1Y9ie31RtqW5CqHrWkzjepsFg/aETFitvLjKaI31EpXfKZ2CdACMsWvYctYGic
8cepwObk72X9eLU042y9lg5BUvFgF9BHS9syxHXZwUZkpgEhVJM5nT9rVsa//5zO
tDpJED0QYyOAsruMXdPS/G8vqDTf7qO0kSyIT1ACduld9sgOvoh2Z0knht162I7/
Cu8jK+c5Dajzujy7j+XqDJcyIcykzOr/E5r+3K7SOuSUbHUe2Ezc7yJtp/Kp/KpM
da8doD/aFirIkc5o3JVs/FsAK+487K0xzjMEi/y0J518n+5zqmv3vHuFevupNSFs
bBG4CmzO767iBOHmBejxVsg1PF0K7921eruLfxvI2myeTKEig9QUzphfOvt8uz9V
P5o6XiXRux9S9A4NCEoHPlJoeMAikKGQL1wupKOT40TyWRCtPK1JHK2Lt+5kUqwp
xAv7X+z88xNJ6iTN9LrJE011A+lnKj2+oI27VUAty4oG6BEuT4U6e7pESlIgCDDM
EB/zxDFAtnT5QTs/XVIIzACl8BWO/cgN2Zu+A0DBC9N2s8iomh5GUQU8EaLj0QlF
+qFT7KAvluTgK1pL/EjfXqz8oUW4kE2Ta71c2WsZniXs27wI1rvRgrYJgEb78Y80
gMCh3GdbkNobxOP+3vGRNfF3ojPuauXBTjQbAIvEwwZzbZPfnQpo0aJE77feDyNT
gIF1onqnKNnp+4Zu0W9YUI0/VKbWu3XAj68yq9e4RptrpwcMW1xPlMWYHMHBejI6
zYgg+vVMLbwhi4aJ9fNKd7qntLTPKpqA1SuPR7fYKt6Ma+LPBLC7DiMRJiND0IXZ
btDfnHXSlOfDr/kayiIyFlhX/QNtF+V1128/49ivB5/SkeweUmmfuz9zUr/TtYQy
VOOKaiwloguRcPIiTipc3jws0u7WOuCL4v0qCFoHtwpthBEkBZer5gPgkflNL578
tXi4Eu55HXpvHJeuFwdQVVAQTIr3vBrWqa2li5fNvntC0Fhk8pZ2lBHXKEkD+lAS
LaebbUhP0ocToV6VJjAq6TO3z5ombV0R9+HqxbcpYbh6h1OlRFTTuwL17OJQE0gJ
gpnt3a6LyKLT0zVaecuSoRtcm9neaz2fhKpMPeAg5u6czBjHsp2QBi5x9Y/0P7FS
d2N64XIn9JmcfjmM+Hz8jd+aW5DC5iGVDQOj6wEdK89ViFqbX2R3rFmjI4MmQQdj
nn9fq9+ZRuWkhw5lhm5kBwrVh50gN2t1X1lV8gByQIstl+gAeh9zcKSw8OthI99t
VS7T2BxfcCGN4WK1apF1Nb0XeX0RQ6b6EdNjDvIJ7v2uK9teCvwvFDHaxlyvaXug
cXYQ+42xnnXOvPVrdLPzZQ5Dp0h4r5QR/J46pt4WeuScCnJJ0h1i3JJaUDWVIYgW
sPqBRyJ8XLUP72jVMzJOVmF50ZQa01B+BftzmLCAEY+HRzyCKrit42PWAFP7V7TJ
UmdJTKpvgwSwr+DJlbDleeqx9wUctJad5ub4FKdDQyNk5Rn8M0aLiTYombVAG+0l
GgcH5g4A252Rlza37qW7GJKTG2t0/0p/t+AkE5OSrptcuMzKAFDYaUuW11kVr+kq
e4nHri3RN+VRCTMJhZzd+D2Bl4x2qNKduRcPMWDrYOOpfjl8nvauM77DkTUJHf5k
HSTisBr3isoVEFI0OCNzYMRvGLXno/mx+6Ueq7te75zWvLglM61n+Nk30+qKBmVs
qdSJ2eGdjvW9Bmeb1q5wE+hk6S+failDPgdhKOiEePqFHSFXb6XmQoSHZihJ4ulL
Pfk9YiilM8WHZZ7P6wNexZ7jSCauaQmpyIgItc09JNBO8VcjV+3wNidKCEheyIuQ
c77pKdTtTfpSQVeWdwh2Ta2Ou6k0Rj66k1NNQWZTE759Kc8rgBUyPpc7NtsxQdwa
bapROx9TtAVCjeURnBS1NjK9OXakydoHxQni8BeeKtqsIPFzwO9zbV32iLWvBBDD
26gk1NO15LwxImE6bg76/SotVzpZlEeS7CsjCZaLe67E6uRM7xkf2spoeGdClJhE
tcn/VUtL0wvtDRJlpugYZndJ7+rqxGPW2bQ69Qcyu6gRYr/ewaDbDEhIerLyJdzG
+XVMbQGR2aF35hQTGYdAwQFXf86Eu0F/2hjamf7Nfx9TVxcm3BkOcKBpdhkVha6S
QiPFCZqGkZOAMcW6MiKxR+wUgfXq8ji2eEEZOmB1A9pTPmOgbWgYh03lWyYtKyTP
Ssq280dpElTmemCDxZRxDNfnLVD+phNWKFsSaabmhIiAga79l3x2HmHSQpCjNl5e
C8LHErnrCDyQeXXmxpqnA1mnnIgpmRegYBAexmHzQxzTHe0Epf64sJLLbYQriYXX
xtkHzAARULF0UEPWVoGuQA+++OhgNvtERA1Jcde9MTaWjo83ZE23HrCcbKSO2fTN
P3qbnqIPj774UvEuEDtJIOZdiniXvXXGFS74sxIcVL+QnQev169dSShroP1xKRET
dBKY8Ij3fMzLymdSc3JM5tx0kRkNuOzYzFHBsFr8VW3qbSw4oRNZ/djvnADDKmtN
NiPc3zCnZy8fMV7Iyu3I7J7hAbWBlGj2yGkxGrfMOTnOBodMktApVi77sMWUiATJ
wbFzQrMDoAxaUo1TozK7fINhNzloZtHcV2sTSGC9TaK4eqeSvtW0bKzdaloNeM4D
edg8GOjP9WikU9bQ4jBZMnu2UYQrQ+JB+ehwWIdUGow4o9Jm6aQaz6f13LntPosF
QhYR/R06pfLQY8vE4Eh/QASc8Qn+WXga8LnJaS2sb5luy9BIzATpA17HX7LoMC/s
yEZNFmOz0nvjRyWZesM5oIwyw5Fpa/CN5S07etEAlvTKOM+CwZs/NcbNYcMcuG5Z
HjzVLSCy/pG7cG/I101tZzAAv8+PqpMjurOkxFVz9s9j+3KgPwrUBAshH+siOtI8
YU+ha0CJyoL8vHf++/1R0OWyYLNngXbG1d0Vumxa/RkiPbBZPCpRH5xIT3cjtqUj
SYqPAnYnKcQG4izrxs7jLOAxIUUUNZqm0ZkS4RywlXp1YmkqOMoBnIyQxNSc3I0v
fms9Mg8jFn5h6BA5PmktEE3cACKePCaf//LMa5SRnjNqKK0AR/im/Oi9EGlap5bX
zzbb/niSwa0SPm3F5cvPb0Zz6tWsv2pdFsDV9iUnFQ0TKoohueMjzzPUUaIXMTsF
Is+rW+FGV8PJtAn+j9rxAOKvjQI/6BbWhCw3Bbqxws2Cx6rsKkh7d0oUW1YZ9WEv
awOmtRnGniFacQgMwIkEQnxKu0tu57+sUBtEuNsArcwosnEujpdXJR6CHPL5VJbM
Qp9cJog1s9W4ivY+6Rw05CgSNC71+ihJrayot/pj03uJZvrx00uDfjGfwAgJDoJu
FUXGeSsGns77XLD3MD4lv3mkkQ+Ne0uHSxl1HWDwv38rBGS2hJOvaaNDwUEdhEMf
CxhmW9Ebd0ycGWnRnlI70koD8n+yHEurk7myS3xMhkV2apGWXZqZIJcpqI2z1iDY
K0TaYA6bv6i4LsVeHnqVAIK56GuZqoq5HKwSGgDQRD5xZwGq1Sabob0omvDwTacU
4rSpELRUWNKlMthJFvni3K9445/q/sn4/mDFuBzdWG+ByjodGjGb2VDFwYwbCqVQ
5uMYatcQ0B5usuMCerEiwLHFU4IAYzgXZukBBoJmuq6LgX9cW8lwA3VdxJFZ93V/
VqwkRkY0Kt6EoCPP4LPmiiSHn1xTN5kVfjnM1ZTcAhhOWlcuGJ4qI/oMG9jJNIUX
uol9iGabw1vMhMGEyKvet8rzQ8kk5ZpdKA+HxGd56aIx+pi8gkvGAhR3cDL2+IKe
E766xBlqvu+VCinwXr1mAN6MQu2zbp2XusRVUeIx1GYWXJJUWZCKBsgCrbyPPLwJ
xw/RHyAnfUU17vCj3XAyOQNCiYeglHORVlZVifcFdGOdMBwU8TieYMRKrlWi9mEY
ng3n7oYjrpbc/YDXxtiP6uL9n6s1Ynj7AyabWtiKAn+LZOsOU6mDlhSAipd0pyIC
cXLK/rCGsVTd/wW+AzGfPxKbFNchjBlpC5TSiq0QfXlLE10uh981OSJtJXiHQbFZ
PTEUUy/UktwNQ7eJu41PwvIT/NjxwejFOXrLmmc95EGr/o00tzPowCwxMCD8hs1U
xg7wrdRR8l9BorsZ+mee+G4XnqLwJzb8q7/UD0OLfEMKyTO7dZoWCcUEK1lDv87K
hkIEhUoHP0aReKyh4LJmtAdv0dZvi7AYlEfjBSYnt3CF+lUJVw86/zMYr8an9B44
FVKt6Yd+7kA7imgmG9dvNzzD/okuy+KHIvx3spHS4SdaHhtcliOVThuWWTQD8dYw
WciXjkV13ubFKvQDOL6tWltOXX9HZtbRNDWLhR3FKcCIt38ElwGVhi7xI3sHj0oU
bs4wW8ZX4fSsRikeFNET8Tu+hd3fnQsZ9BRZvBRgujZNocx76rZHH0STGUV7IDQw
uwK2gEfBth2f0vy7DGZCL8vzGE/e3G7RWHZaEo58y85+2hE04R0o9nAi9+GgHb9Y
7xocE48PHwfbAG/Tdyd3/FE8RhwYGo08+VQx0V0sO4knqvDpi2WUA1WY5lKT8Je4
7XTywK8kc/VPVaeklExb2+53r5vep68tbvaDTqyA4Ox4k3CxvOWMiqBSacpTuD+5
jyZyQzVn8ZPzk+NLehNUoSZU/B7H6cmGR8pI8SdIX61tlu7pRP8JCyitgMmPYh/B
oje8QgXd7n2Qc+YtIvnqZvucplEI0gEPIAvRDSOMlx4qRAJpWqHBetgTI2iGjoSL
ysgM/MMDNtFCSZiorPb5Pw2ukCCy+A/BUlratpgzVxU4SUEvqTkCXIfihq7OSQGh
1X6N9W9laZkwJ8OopOh+ahH0uDWITFPqxu5X/O2IaoTu8iTSIMdq15CWWgaA2yS8
FIa/226LSu4t2Cm7hnxT8va4zkRsufsXGruUzpiAzab9lxlFtZmrKt3mFHjrnsLo
4CpVUsiMCzcbklXQyK+yZqM7NNj5Z8mlod8nNIkxUplnPqpzocrjpO3EkivimuhD
7IZUNRXsSr28Zt+MjX057DfixwAht3jK/tYjakZB/1RAYujRc7WDinqBfiNw4ROw
WDcC7THFcKile/XIkqHP6amiV5rAGO2eQbBDxvHSxZVlHB7p66m7P+ZJ6FBXBXTJ
4UDZ/Mt0Cj/lKbO22HJznprIX+fqEWwZAC7HsTCsP/aTqm2yuoBYUZyTGStTZqMU
qITsOWgYatPVRs6aTCkDEEs28hFzt2Ak6b7EfVlq0o12t1ACLP0T4C1nfcDmC6mP
9X8z2/Lmpp+yhnhkpgMTRsQqRzxHIFazbgD64G2czKcMFVyxtHpPGgZULPyKEq/c
mqqhKOEKc2GujEGOBaiv0ON1q8m2aGXBDzkb0zoCj9jJa8s11BKT/u3e5ESGnEm0
tzxoYFmK7rtsrOvy5j3lwBmP/GorLZTXj2J2id3At2T9Jc5blDZiiqhCtcnscPcC
iA3Iv+KEHe7PH1bXYPYgSQ1q5j5/Ar0ZqKAJ7exR6Lbp731aveLFlfo9RglzF988
trK3ZCV6bmXlK3aZfa2IZTj17qi7Gmw2dHLjbPYgPXW0BmlikhUBPPM8dLApE5VR
Bwe3MSrpZ3ppYUb/J9Z80Lg9UDDG8KAC8BcFyIBs1DKU3cUrNpehR5qMLZRgTZ+6
z5IVnxnaPwfdL5lwKEEdrXd4YocmjHyP/NmtQuTO1Et26QIvu5w9dqiOSmCN7802
KeOOtbd8cs94TpQh6zfBfLvKfMSx4Ro/htCbDaL4wq/DMtEUql3ScISJaM1vk5vC
e3a+lomL3pnPTRXq0ZAhQCvoFXZggKFbQYLCt3armGRPKe6PWkI49in7koWDk4wx
cQosSqTdvdmYJfnogSYMtLsgfHjaZeK2mvC7+B19O1bnlSdtRnymhkseow/0OBjx
iqWMljlQ2OqMv5To0Cugg8wLbhfMDKFSQqtb15AfZf+hNU2e6hDGvg42K8mCQXOM
M3U1UX6TUxu9RYP1SPOPDn8SgWMPSkOzX2DFdchSTneAwRaSkbVsvL1F516LlUAU
wT87l7h+e5yeD/N13SVFUMz4yC31FS6iS6ejXQFql1fuDWlG4GWsMJ/cv9Y6jZwn
uOSFRyfcmhQlzNKIl1xe/bg3VQhalOJXSTyxvpQOulbiOyZEJU7OJmdvh0EeYq+Y
QekvqgQwue/ibz601XM4URxBJHSKqtXbw0SNSvnlK3UAL2/RdMHlx7BYCnRYi1Kt
tFzzalkpGugyY6KT9cksyzOzIpHTubKb66k6SK8UrIQBdlqrxQ82A1USC47JQ9CS
+93y0NgJpoRkka62vmFYS14vWF/vhxnyuzwhzJDuSPkMyTMUUYXYGox/PnRFPoCn
bYWOjZ+D4RqT6opighZRa6KRFRpQbg8WIMr0twxxzxPWZvplSE8KJFMQsKxwc03u
uEsu0Hwtj/QePbddwEPQoI2Kl3P+nhtDmEA3MgD55KPWjaOZvMm73AlE7zzIV6oI
HnfX3RHNP/Bc2/ANG0ciVsj8x4lIu91mKwBcozvw62O2NOAhfkJa5sF30roc8l2Y
McUMy+/DzNcU+CbegAMPBNa8K/b4++w+PqXSf6FH/0S34ZSVaULCRP/eKz8H4xBj
4L6qNGtse1TN5pwFAj9OIG0Grl9iz1tBwZhmizo7QYcbw3VgYFNJWhyTUH5U3j8f
edGqKa2cvUGbjIL8ZIu9df8eIUzh3gYdPbxtUbXvsNhjd3oC17RuyuGI3+odL4Ix
Ih7Z2ToTVo1bL7icRl1t/THHNzDUWg7EjAyAtmdrjVvcyo5U3eWns3pkmXR7qsOz
h4CRSxAEvv/zWuwDKcZFcX3JBFzDidJuU3NLF8/hsoBPpqsnG8cBzP0W8lRBOVHX
mrMRVcii/ljA0kQIjDxhZvAmZ2zjWm7TYe63ns1rvo51NhHXuYZU/KSmRT44a0zh
C5Azrgza/Dg6T2ORnwUNPvhnh2JTVHiJ5EGOiI1u5EnBiSiw8Be3g4BtfjXFfk3B
77Nttp2W3ZY38iLub3WQszfKcc0I7WGZr2QostplwXngK99Q/M8hGxvx4p02ahct
Xiz6vb3vNmMWYr55MmdrovaR6LaqsEQpCPIqmXMJz6UwUCEBrdNeSPD9zERoQVuA
w0GZtYJQJOzOcrpP/F9nKKeBdAPbWFgMlruDe15cgb2PZxJ/osZwrx/rr5lEUPzl
J5FSj9Uj7rEp7sWeAbW52qAvt53vNaWew1J3C94PkBv2zn+7LOA1w6mWR8kto5tP
zhH1jgAvbvXmjie3V1d91VsD8zy6wvZOvH983QQA2jyUYegP3dCACfIsM03dv0fW
q8+UaG4r9stDGKGJZCMioTDjSA0Pwm7CR/pcYPNoyLsdBIgJRVAPDfQlcfVWtyuO
NBWm0sFRBl8pIEITJjG76CGatPYhX3docynZTyc97UOza10PQssIYjeKfNUnbNSK
6GVUNdgRj8KL9W5j/SrKbI+pzY3ma86HzPPEKPgJmrfwoC8MjEn1gly+yiZs/Ppi
fzCb3f2nAaZWsdzV2lEEkR1d7XkmAWQDsuRFyLZwRPFGjCmBT5/LLky1SkHlv3D2
RD9zt5Vl9Ihc/IovbG+CFfqe+OT3cgpxK0K6lzZGOGHEEwNTHb/J1IPItfgyG5U1
Mwok2JCm6z7wOTmBgu2CKoTC7ZlCkjjkREj9IZa8TNHJjQGFJpcNGXfKuS7zJd30
eLpskL5QdOyL0tO7UNmhG1RI2W7UaS3X2l7zrF865UCLtoM9NlJw48iXZOCbPYdt
PIfToZ8TDjabgA4xPXOd6YUD757XYhGKayRM7N9H6/GaEMg5XU4CrW4Ho0c8r7lf
FulKRJffRXOxRnEdukl2OFfEShsDsHAjnSCyz87se0cS7Q0JfiGqWDngXKS5ZiDk
kDSLZ21KTFiIFrM2egp+Xdrkt+qu+1exooZAV53oHSp1NPaimpQFP4BaJfv1CBY2
jDCpUoA59ZbctMWs2SwDnCmZe+98yc/LTWJGWAiDmfzbJP1T/+/k3jsjRUSJampx
G7C9dTG0+h7pVIVFy/t18HTqzv3znEoeSbhlOjRlX/srsfsDRAUinyX+AL98QwD6
j6QlEIYTk6Zph1IkLmR80qi77MV2+7TVHJVvfg/Zzo1vA65mqKfEqQwefkMFf+0Z
MzP1b/PG09gPfW4LbMKu5dYxykPOTaUP9Q/xMYOPhH3YLg7LHnlq8gKzM6pKNRm1
aiUDgkR98GMeFblQ9ysKb+ZMkralP94xPEw4x867hf+7fFaAiBEhg6nUv5XWlJYP
ppvbSEZOoEdWuXsfOFNfFxAoU27J0Vo1cYZOWh8tRRydYpvZHB/t/YTkY4+bJEjn
SJZukK+qOC7ffkiahQB7UFeva0UUTUA+2xZqJmH5tkmykGWHA/TBVGD9vM9VEL7W
LbeaNLu/7axxeC7EsyJFEnGM6UCLnt4jGlz8HIeqFTzvKe92JfmRuZnCL+sJrMva
SjYcj7NrrVANYSMJdoIGlS9si/p+bDaWkL+jwL3qGlYvENYwVigbh1ujnWi/kfXU
XyHeT4QS301prj7MhNuJzPt/yEME81B/eOFXGq8ZOZEUIpg3ohEEfpP5YoL3pma/
Lbz9jrv31PCaIx0mT5egIGeQXkLFIw+VomWSmVbf1g2jfmjNsULbZDfqM7Ktev3G
R0L+DM8WyMJXs5SVYJ2QNbhU7d8fLnz8i1y89ZeFgNI8vWZYwjco2Hm92I1HPYjF
bci/TvCd09hdBdKJCX3UoANL6FKrcyhNfT1BWx+Eo61TKi2ltqeANBhZQIo9dB/Q
ZumRbF8CdS3KpuyMOR7LcSJWOJcw574VG76855ahfE98aaPMXoAZcgbvuRzwfxuR
XoYImuMBJHdLx76B3QEdQDhQz+4m+3foS6WeNyiJXhjO7Ru8U7kfhCSt0WGfpjjR
KDbXVHYteaXPijsF5YvCWQ7QFrbaJL0N9nfdpX4T03djvCf23BzCJUYetCLBVBE/
C9uiShm0mOdyuj8qSa8qZdCp3l4jn4xy2MDgjItV/momh5VVcwxZIR1Vfj032GyE
+oObVA0+bC62s+5mdCyLrs64S/AFhZP7yOff51+y8t255E527WJFQFR94hXNkBug
8ghmmhewnWaHBtonNsRaJbVPIHIVNQ/j2gYnkKLg45U6erXs44xsqCQKuYtJuxfy
4r7u13X2H8MDpgXycsGjsibiVFkc2fOEkKIAADNTluzsOi85m3iwq4oGl2GDSm+r
dkxdap+cJbkGNsPUL0r07B4/LTVZu+YK8Pz10JiNeFEhjcIegw2q2mhbsdF4Fry0
KPsy1B9adap0tsb17lzCjHHQgQciy+Yr1sRPu/DmjZ/1Vea+QEyCChS9/LOeUoR8
Lya9tzz4EGbD+C/jmABNKzYwT8fyuTAMTN5k3d2032D1ZmRD3XdRJ2O4s4Z2KjyE
ZcByGfHrHyHEz8gB1KQkcbvrk2/n8Pdacq0Nz/rObRPzhJeyJYwuj61+Gj/1v/IT
W1E6sP+LCy2Q/xO8NcwiCDez35r6lfUwq+xWkeYgNP7f66zd4Xk45qGInZk/4Muh
TXFSb9CoKR9RWnUd+TUjt0i263VH7b8cy+5FuRmvISP3MOOLT+OVRSth4D5et7Dx
OD/SewE4vTa0lNApToQ16BKVWyvbIMGv79YraYfC6feq7S+OnZVJOcSrJhnYT061
2MSduqlLg0QlQuXVVfZ6HI01hd39G4G6wF7Uz9ZZ1OPly0dQvRAH7J3SQg8YQCNT
aupoSW5/eXkG4C5Pz8L1tyn5RQxdivrMjKHD5TrK1ztopg3wbHtDOkwoT99Jk8mX
aTDGLEBhSXotdzySPiBkShNX1rBGnB8o3rVNBP0jqbzgzn4Bxt7XdgslFJ7tIHa8
YDlfZk+VGfuJ9Ahpt//QBnMbVz8bzk4ctc0N9k20SSmBeQoRF2rnOFzt/GzaidPz
+Zk0YIZdPOdrArb083+YB5581rnw8uoSaoYEjr8WCVHSDBXGXSooQV/ytR4Q9YA+
n4h+40uuwSwxSIMgmDzDltp+Z/SKvHaNMmfLtWZIVw/c94yUXyjJuZi6QCU33iOm
1ZAqGOr1Y5ayMQarvbjkeYiU1FgqJ3SN9vmW0k7jO4fp/H9s04wyQ5E2ZOAssoc9
4y9/CNyeqH78Z4B10QQiS0gf23XOpKWbI4nQ68+UfcWAWMe3MWLysVelkyMO7Au2
8lYykjrXqzTT940lREwXjzVkGQGtqMoVhyH20f69BSkLS9x406WqsI8PhKh0bCpQ
gvE2fNnwKsljYBU+2ugUm1ePZAW5IdPIf7hbEDfzRwT9mxnqlQo9T4ZJx3EMEnzk
q3dETmi+8/JVBzYNqSuU6u8KNZcttPod5KQDIFVEQrCOx8g4+FKKLQTXSIVKGtFk
diJfOVifBWemujrN8Vgzkkp1t19QxRpXLOoQ9VaL3uSRAABDaPMxkNHjZG5D5mk8
4JdRJBAEmCHiwFUxOIc3XUOia1KqSyfa5xFUNv8PITKgpOWDlN/N+UzJVHXTPZwH
GYcFiAeksP8iDozW7M3KUIsmS1cV6f/N68+jGZKiXNNSQOFhCMbxQyfy7c2AEiMG
gpQoRamnJrFUgy3J9CJaCkTE9rDVYVO0w5lo+EENIRqlSMYwCzAVnuZX6sNiz1DO
aCRX+jAH6UjtbTPE8Q2ittKZHjPa4/iyY8G6CNs3lJMAWYgWxGS8cDR5+EuPIwQb
V1sRAtOn9g4E5hKrPEziikfARtQ4u3hUOTvZ2nY3rU8PwS1SBny2x1cYsFnvfmId
paYdj0fPoPoPSEYBOUk/C2W+QMEKAL92QFrcLoQTcCtjR2Z1au02hL7PCHrtqOoD
tXftVSwqQSh9H60jOlKYzsq0qlWJNm5DvPQgRagMnMAlWNKWcv5oSQQrLOVazAaH
zD/iHbrMaXJCVLnfPYBis4Qg4reEh2jHpIHha09+RinkdFjAkpLZuWCVbFZ6wa7D
NIhzXEsTOa7hj0IKagMclQsKFHSZWAUvTorg4qgvWeDiUkXc9j28N8f9T2yg3i2y
d/06zZNQ1ovhBW2/HF/Lm93GWFdbgbJPPniBIsYLqLZMs2CN1d6SJsrdRdGyABi7
gpzNqYAM8+wj+Jzb4apCdAWxLpi982UJfn9e/2zRtOr4MF6BKfI+yLjuDb9wx6Oq
vBWbubWt78GlX7sAb9gXy3OGXCIyyw8QylQVpUc6uSxBlCaSo/rAw4xMuSU0yRLM
/vqYGwav0hvYxc9NwFLG8bpQG/lo1r7WNLFtiFrYMkTQ8izb4unHgUhwrkid6KKk
sobiNtqYjGFtCJ2FkjzaN7zgibnEMwW7FYZBrz8kbDoxFlTihtSPMG6n5jxo4sv0
hVjMnTnS7SWsrti73RJ5z/tNUOnz3OH71t1pwjcLmu8ysmIuOAzsQOC6RQm63Rqj
EeqK0r+ydW5aoiW7e+R5R8dD4CJWP9vqRNnbOKIf4zhehmXUiQFzK1i/vYt0y65g
hZjIHHDh+qSdPPsIg2j3QOUjAVaRcaTLf4HQilEQe9qpiZW7UxS25RkX0gQ6i1bX
9xDdqxUWuSgoUtldG0dm8564ERrAppHGtXTxXTzacj47cNGDtkYVQHBq5+skrryX
MMaV1ysWGcLcLYAZmqLKSQVByoGk6xcsjCu0ovp1nZRPqq9Fs0GoP36wl+IagCkt
5pi4e5TERcg1P7fZuTdySRqoj0tsfRiQo/3fJMUa4yz3vLEno9TcA+ONGkDlrfFS
w18vaNzec9MqNTlf57DhmlbiwWjGPNR+oE/kgZNj98kBlJiugM2UiMLApfOK7P8X
dbDfP3rRDfLDZZhwAEFZjIhw88xiyysNzkGfB0Z0ts1TqWS94eTaABrmgiVmfvRJ
u7OCjGKMi844aY3WHTzeYW8B0XOpPj2R+OfZJfAZeFfEGYvid6fuNL/tRWSiYZiZ
gxr0f3GsVlx57CK7XCefvoWg2jaxSqXK1WhTGcsrrCSNoRULj6LlCqjhqVDLRKzq
Rfy/ZxdolEHkdOE8VK/qfGut3xKIeV4//48ni1wvIahNXIHGE3LEDZrwcuQUQRMS
qNqgZTA2W0gWOigCifdvOSMeBaI3MbHAt8r/nYhhDv+9QYTWkfHUuPcY8+UkGC8j
Bgs9yEkJZTBbG7kfQFaTTAKoya1qr38MV7uaMy0HRfmmtPOk7qaJBNmRuiuJe+Ul
YX2FK4BJJVfHFtL54k5RR04HJVmDHy3DXaNQbe/P09GmHf24MMnvNCx2k+WxoKvI
yn8qXkvKE2x71NerAQtgO5w6JBLRyq/ZnaYhfZ6kM0yoeuFSdhZfEw0fV/AtALOi
npvkFAxPEv/5Lr7cBZwHTIvcoU7I82d0vcJIpSV0YedzV58/GT7c+HWUVeZZYyII
TSmak7IMhbrdPlCcODAFCRHYrp3fIzdgURB2b3QOQvM+F038zj4NBPxYifezQB37
1+D1mXQ9OjCmPCsO3/JedlY7eq+B3hTwd8Tud5dpEAq7SGz/oRQu/xHZi5nGPxmf
7gBFa4wn00dkAMUlOo92IERn16FvJNEyagPnn+yAb7UsP84fkOF5i3wrp6NUlD+L
wFstLL8VSTSvt5W8x6+KV2SGoJG+VcGgVLZsgEVOXChP1cXZ6m52TwykDe7fv/uG
V5EQFtO4M4HdvlXTLWQZDKeJ1U44WdXwLyqhHogddSaS2yQNd7qce5uqyoqHBhj/
/zQLT9Th9r3jPLAb9teXpbwxob/6UNnbdNVD5UFPN1pCUyI8WQxb1b6m3zC2xRN6
O0BAVieQxvwotaAK0ogaxNDXi4D+I22UYR36+aI1RlXASL37iHwOO6D6J1hVQ4pQ
u3Cx0Af+vS/3od6Vj/Sf9caV1kckOU2KnIhefkGlzEh0HSjDCfG2dnTD+efxDLhb
C038pHZH+mwPb+q6jOl+6biSZxdGzn2rFLg0z5h55Z2db/p6AC6y4SSWw7ksaO6b
z572/TXXrDAQzZtMrxeKw3wq4VbdMd2SaNrqsYCGKnYuQ7t05Na135mw/tcLO9Ym
wQrdnxBRGP+AgzDNif7Rsl4bPgmVpJUYCGnA/85XsGYuhzfUUcsJCCvhr9Hkpo7/
GxTYsEBbkwguihAORi8PUzADGEk6rCZLrebuy+Gur/wFJpZkvkyNSVLCySTDMyMW
6phJQ2B28n2JK1800nnhrbY6MjX4/GOwuho3XjPgcOMLTnh2nxtWDhm//kwDJjfB
wbXQT55PZdB2k6q6OuhTRyPHId4vhwfUwrP/NBa0jZn2plXdpdHJ0V8AYN8264tV
0O6rSFfMOhjBG5zlRs/6HuWWip0FGW6ccniW8c7R270Cz9PM2vNRYI9LMxsFhvEu
pbPi8Ips2yf7ZlO7kutxLiGyboj61ZJMInQxejtBpBmAHiuk+IZOAP4EsZkIQO+E
85ewGX/m0NdcYwC2yw0zahslJFfshGZcvDxr1PYvgpN9EK+RTEmxomwZXIb98f2a
hCeNjqcPhcQMFSEHICu8kyJSjj2jDxPpav3oi4l7ouVbMfNo1ModKf53EAt9A9XM
W0kjeZdaWVSvA2jnS7HV2Gs5rFjXA/jN5jjcPHUBw0qfMNmygRWcuL8WEXRDqOKD
lmqlLcgE7yUvJgawkXgBh4eBN0Yw6FsBiN80C+TQ8kl/LwLoBCMci6TMl2uOv6rL
4LeXqR0akBKer9Y75HFQuzBmmfcCjjYbsRyIcVIcX42axxBXWfwckg3IzfcFL9vZ
bOzDFWjJZFqMS+/j/DuNfnowcoXfKbXRyDIn6skVmWc7/l9oYATMRYSrw/yHi62/
5aW9Pb7VS8BPOCuXY0GsVsFpOlPXP1/syWT6/vLivOp2fqvWHd8dDyz/G4n1WzVW
aZpJdFpiMMRaHtgF8iHoH01FhEcipnnGNEV+t0/B4lIE5c735TLzqoF5nHyPIwZS
2TX7yMqKAOkZ3QT7xG9knp2hLOXlRSU5csGAdx4UDaENuU6hQpsFZZ5/Y1M2yuOs
uomPjKnYCbFbeAdJ6F6LAGYDc7v6GNX+Z2tooQ/I02IBZpazAN7rISfkxXgp7cge
cVdxgrPVzzCr3Yx64g6qKnk32cYzhjywTNAYwYwHAjC+zB5bgYB0gNDAppodFWUw
vh/63bOAbdndSD+p8sx4oxBV86sMil2egcykYyHa84A3mRoI4TPSPkIyMTAqqi7K
AUf5r4Eh5cT1jPxVdVoOPRBQS9BE2wTMK4D+O3yVFG6pJRH157obJRvm6hMwYFto
9FhMGFPKfLOtAR/RbCeKazJOrfwtt521E9GZBPFAQh4Zw0+XbubdtU7PcjC6lRVZ
fZyNkFTArWAk5SlfXs3nZzoyAhMBFNZYhmLa7PS2ul9nWGwea9trtCeAfmjh9Vn9
gDnwdjAZMzkiX38SHHCNtwazcY9FsAYIHd1zxhW7ea/hmYrab2uWM9g+Db97tXqe
vxLoKYjXo+HOTpTh+XWXxCs7xvA+WDBQXBsKlngoJqoSyhW6021ZunnielFk3MEl
AT3m4PgwrgJzciwvvGuYacDn7C3Fp0Gx3RYE6eAjoYwVtK+rrzyhOo7L6E1YMIFK
vNqZP+aKsIyw3l/tVMGRg69KHTQ468bISUWo7WyIJeawCju+E96T5ov0MPz/mL2X
Q/FkSMDoeLJRjvixERfaV1xg31MJWh3EDMc8Em0Wk85llqK2xpZ+WTDLArjmLmBn
GHmeH+HOMNCLwzxMlz6gKRz7pgYiuOCm/kNO3s7pf/uvKI8goZpZ85lN2qa74GU6
EUdHnZPceoJ0boa5u5Ex1249jzy/EqsTn8wB2EJTZmgauJgtWRGVR07qSjIfegVh
Ee3HnfhYTBAkUPualBNcY4LkCWCDOv+aRmeBramow4XnbGzupCpT0RHM54+l18Yw
7+wp/GiPP7fKhlGwdFlkL0+Khz+TTlL4kzRKVaF9g4GPOO5NWwX7fjxEvDSRaUPo
9DkO0JKLi7xmV1Q9tDWigkJmoMmZX70bNMj58UYzxQ9DwylWMywbPqCgWqPp17l8
XlTqvWekPHHRxuT9+NVMQR5cCMMwWXT5NDbE5f7SnZGXUQP/tF2XlRdtICs9AQ9P
iOn1m6V6Ht9BzpYLH1zZ49twINxsCByRFozkr6TzgNXbSz+fpY4pNVmJJ6pnE1Eq
eWz8rN+5ur8I9Qir3CrIVzR9/5uSWsPL2OUrG1aod9ARjTIdMMqfZhyGg6IT0UvK
WZX5BMQoDZV98XqvdwT3fJ2fs3rsX9VtPnZm0m3RuWjJRge7oYbwrwUQCZxII4yI
8Hqkd5uZlJ3y2cVIMTDYqCQhohhllCeYMhLFOZmXB4f7jWI9rObaftN/hRC3gciX
gfbsnv+VsikrOgmCiNeKbh5/FmIH5Qg5sQCEYu6m1apC0EVCKvdnQ687CLq+lRIw
QEIG41bKtkyUq3faDCk7og4dWELWD5877I6cs8/0JshIebbhak6xPu9x/QorKLPL
DVnLmOAi7rBSSC7a4jX6kWRliGSIslC9pz5TtSsKXZhznLcx42daNiWqvm72btdz
PgjHyY3IhXgLlo2ROZi29Uh3vYMelEuY2TiPs+GOg9NDb1Q+niuOigG2ceky7Xmh
NF3GKsZiYsl2KaTsBOd07y+J4F7pnEhQylsCtU6EV0akK4unGb3tdKtfSe945K5R
tt6ya+21Yxvqgcl0njrG48LKZ+3SBmdTkk+1bRwQIGUcqecI13R1GP2ISxm0UWr1
liSfI/f1lw5uzBDpEAGg4EW7lSb3V0fKAANXETW5lOQcqP+RZ51/nzf0lEn/XWXu
oE8l+yCsevE8dd22tpKWtdSais0H9dnrcnC2z7Uyex2s9s3SI5+wmIIiK03kCqr0
j80r4DVZas3d8StWGgALRBIDedxiN22owuoWiVsaKzXLxdrWedo0Q8xek6zZo0rB
eGMvhvuXWv9YiHpenDFyjsf5LTqbaZF7HilKElq3T0UpXc+FeC74qtfBZ4s2Dywa
JYejIpCh3EMWzPVrcPrZnMlx30g0bYsJxRI6NzMdqh7GW1g3qjGh+MfHZ+Bnfuad
5aCwotmQPoUUvYnGVY507V6mLfbmhxw0TrLPHJSN/Vdlu2tE/BjQuagGafIdatIq
+zsinAosTe1C3vPQ/jQi3IgJ4IpPsMj9PfPXDp0rcpZJl+0y+LK6vDud3Y9p5Wki
/evtsneVAT+QRb7OslZyesZdhmub8qeTOtLtYJK+XnW/i0GyU+UB8/2yntoEzG6Z
3KQwDnyGPO3lAeVoBKbXPOxflQWa3GfY7TNeVzO3U4gDGlwYEwVr4J42ubiPdPm7
7JYJYt0L6VyJGN9o5PmgjdnYn8WqtlHxbix6atkG/Us204x7BW+lelputaT1w4Wp
h0K4wgyg/bn9Phonox+PtjCDi+tkGmhMXW45dOnubhzDH1F+bSj84yScFCgztOrL
VRaX8qHfnPRXkEJDSLS42j9EoKGqlv6U61oHZMb3JbjWrXdaWxwgFqbWHv7PnFUB
vOlFlq0L+78T4bb93BgooCGa/f3Yvyi9X4U8tGoeNxgo+I2Jqr0KDuijvuTo6HZj
hPm3vAilMKHu9bE0Bpv+iu7SRp36+5PqTD4aSpjrJagVJF/I+qPlZ+UdelXLgYlL
ZJv0DjItn/uJqqhKiiyo5x5z5uWLYgRi/L/e0S2s20pPmhkT5BFeUX48hh0cCqBo
7L/jEAOr+JrvZTEruccIriTVW4WfhBfuFWVPohyhiIhM7bc0ZhuWJHf+R3TIeGdM
tEWqYKPq8DGUeeG4KQw818d/F/ROzyD2cT8Yl9/ko8LpZu3M0OIM+CCW8syubksp
xFEZeTOE1vOQdJxrMPd+aKYCq7I1cUHc94AeJDP5kGrzkWVZFqWAycgy8siZgA0+
vdBmqPsicxqVQ2hh18BGAV98aptcKQuYhI07J8QjYtJl9go/pf4qK91Xyrl+VH50
xgDiepI5ELJH94zqkfPVMrAi5EGWzZWrxoQRxFyFuino6MM0HHEXCOR1qHoMWd3u
v8Fve1xFLXMNd9aVpSjYo4zCmVxJSilo1HSpPlcCV7D39Vevw6+6rX897RVLjMGa
//248LThgWwbql34oIuqQAVl8K5IImWE/JBTB1tYmRIc/PFe7fgXCakqTO1KM93n
hfIBCxJ6mUJ7WTqD+ag25EL0K6rjcmxVNzUQI9TXsd0pDTgVUDJAvjVdBiitRQHe
0nZ/dDtnIGK81Mj3bVozLy3kCvylHPl9rWVh3NxgsMlUNYDP6pvo397Ta2IThCqI
8M9foNIzvHb94eTj2iAF39kfZRrXBPcBMRGo5jfXA0+kx0bDhrCzKYBuLgb8JtZC
tSiQ/r/AkH1q1Yfr+k57fR5hWXgJZlCzglF1poMtq18ffQDfF9wz+rb6Vqp/B2w0
pRfyWJYS0tqv1/HDZnus/+s9Y8jAWrCkjGOPYWJMJw/KyjAAyCZ4PKGnF3uhHDnK
5/Y7AAt7koCIDLSiBTF1AVpmYMOHttShOldzXzG2u4CGMiKgv7hzESWjUwhi9qxA
Nd/RrsoL0Zw/DbgbrWz8zSSGqCX3jnACkLD6Vfa+8M+oEnmoHGZsBRiH0IDuTL41
ryvS1gBGmsPUL8R4p12QXFKSp8h6g67XyYSPSnpn0ge3+89y3d0BPShNjTXXfg9G
drKPYpFcDSp8Xdn7Mcv23EN++Ghf+CZJJSF7IjfW6Iml5qZEvD5vdyvDDhS9gkQs
bTNZ2w0oCNZ1ICec7QCMRvvrnZvOQniknPWygpCBlVsBuDKXPnszykf3PgevAZWF
9jy8ByANb45BaOT+I+K8Ga8DdegH9mGqQikr4pu47oiRaFfTmtjLIak102UoWMeS
0YKrnZ0t1jfXIr5LJgvycXuJeadXJERkjKDAwKMW9mnNf2Iv5CH50iBQ9iJvxhT+
7BvoF13faMe+Ok91BLx8cDyE5w7RAlIP6CfiI0kfXpOyrwQkoUmARHofIS9epIAH
poFy1pSY9dHQfrC80mywz1n5UM77DgeGH6bt+XHCq7Yfqia9uEwZ2bqejwc90D4P
opMYW4xyMV0/t83ScOBGNIiho/2hh1K6sOCXh8EBmsSlNpD6wIl0N6g2K93iuXYD
+cxYK3pCPEHDNT/OzsEgzJ4dMQ4jsnDLQl9fAsfVt9UZWrQ1AEbUxV/H0u2I9G/a
eCXjUD7En38kVmDHVRjwZ/z9Nv9mcYytLjKzy7kkHiQnbcn18cdesP8xQM4UAvJf
4C7iEz/c8nOIzUNwYR1Ap6kAH74GtJY+3YDZb4vzKkVPnB6iEo/Yuad/sXUiBdcq
CD3rgvHowLKRNpXubIqydav3bIRaZODILML0kuIoscUxHFQxelQfyKg/l3ciRIhQ
jVRBIVxJ6/Dt5GGxOwuIslvmUqBJY7VwLmatkUuJvbgWcRRu6Kq9RLREc74CNu1R
7QrUeTThSUhR0XSIpvWiY9/lF4d0P34zkVj5nPYk9OrqsAvlYlzYOXUH3xMgy2e2
5YydKAw0rvQbofq+VlOGm/XVS2VBlbmoJjgs35utA+n6o/CXAFj6qUQLs2dR4uoR
T3Dp5gjB1XWpGwQNDU0W1wRppL9tTHkPMCU1NzF/AFaCJa0y1gjV2W8tFlFoAagp
lm1eEvESTou/fimy1R0KNtpUEqlOKX+cjAhPAz8KC44ee8ygN9uMSTmST5iabBUY
4ODJ6MuIl+zh/0mHZplWPquQ3TQwKDGN6pKz8RGU0ClYNSbTUIXo5r0Y7iiOfenm
6Nz+O52q9UgQJLVpoqkTU1d9ZZMZPqNu4ee2uY5AU+z1rKYfGCrYEEkHsALm/OV3
TQz7LvQObSzbNFsN7LqXKrhitTBhRtpnpHeTtnKfSr5LRWJMBvrIjMK3VL5ungzu
3PcyBVYVfKTZ56exwsVhyzGyY/QSCpL09I8rk2CuP5x/nu96oRQ7EXDY4o81Y/3z
wM6BTzKgY0zZKYgNC7w57h8ecOvkjLiuqwTlUBrXHbb2+v7Fn9Fc28E712HqZOxS
4YxFr7/DGU8rX32erSYEMjMdLfNoSpAjqBEA7DpvOISfEQA4vKbay8xKNQwKqYgD
oxMUvtrixxlMh7LPkXFcNvmPWW8Zt1lzXGBr38octszgRFBqf2fzdwhppuCGC3PS
OPsysqpjdTsTcx8KLNYLhpRNTsR0fq5g+EJwnOWwmwKpTAmMj/AsJ8T4THoaklw6
QVUfO+liAikr/y+dpH02Ch0T+0bRNpNvLRu5UzmpeI4vgEXuSufksaAzgnqu7Pmk
Riyuwq9l0VkzHajxIWLvFFTghEtsGkn1+71xv6dWoVvzie4dgF7UGMYqddeSX1Ej
udLfOFvYHm3x7wFUk+q0xWcBfsfao0M9OtIm6B8V4oN3edRcVuNGfYt5GvRJljsf
jloTz6LxvhSpktPPX3XcxVkWN/xOWd3WgawKrZnpVvbXIRbxUKbHeZWDJ74RUXcK
M9j+/A5E5tEu3hm3lt3ouUQksTSLIdC47xwFGvKhFKMHWlQJCaGVBYS+DV+FVmvq
u5OhGV9Zbr3RQTumTh9U9gYL3Zs0AWjEmSneEcEfq8oCIMpA2lmpJePZe7rx6K6A
fAtEftZx+Pv3gXtJdXb9nM3+iW2QuyrYRDW+1ljmUp+UyAaDVSwl8UZX62LgcTzl
h0BS9om8ZNDojFEjIO7CFZSjFMp/ArPN4nAQjJLBQdTD46YMD7V7na4zFKoMjiC2
DiAl18NsWLlNkd0B4iKHRLcX/GzlXPpHy+Py212YvZ0IRjCX9U9tQZrkreWCTbTm
58hIu5/D2dJGra5YINII+OuDect+yIRYsTI0VQoVVJqahE37lPnicaKWywKvK2Ss
pj2178Lzz3NBy7WVaLfl2QCeQRHjKW3lCzAfnhjZAkU2hxKwc3Mw3bqmUn/ZAZvU
nCkvDByOBPfIrCqmUzEcSHZ8I7xvOQW4zmeRrJknTAXILpRSA/UHlhuNqLxJdwNN
9gK0WpO+pM4ILGG2TG5j92a2qHYYfFf0TQEuuatgCOCq0Wxhv6MzJkOlaTS2iwIZ
Cg6jlDWzQunnU7WtMs9z0XnjHeGH83eJtbAjMZyCmJTFnk0dWSEOesimFfW5PxFE
4VvD3raINQ5a/ppW1z8TMesRMuBp8onfJBqyivYmJaVyBgt7CA5mf2p+xObsNHT3
QDrsKyR3KUou1VQFS8tMxWtxTQHMs0pWPQAG97TZeY0miWHeiRyGvb1MpIKKP4ON
4HnmWez1asd/XBEA5tUb0qy3fz0JsHV8W/kAczT4DMWtMlDrAwBdxyTrbelQHFl0
hAcK3Hcvc1E46BVYXzHauCVHO6I2Gfu0IDwV/TT+5qjWChVkaLeTKuKs/Dio/uhg
GqfVuVOg1qr/lmKalgZ9JncbCfxY+XEjJRm5oGRO88lztqm6bbIR0alFIM/AXpZj
Nr4GOfz/cePu3GEsebMePKhVER8g43QtOmnVFFa088XRhXMM3DzVW4f3xpPHeIDs
AVjh+9HX9WUD2XHMop8cg5GdQZHxnWQ2OIRGbqm9y74HzHUuRAYgj4FVpqUBfQfs
eeEG4unci3TQ1vQ6wBSHNd27wR67XVJypXyypcpFkozJbaIznljEEQi3RH03JTFB
bUhfeE/c1QEdGDf7/b2K4xtUfQm2MaF/QilgyHyBbmQDcsYC+MmUTv3dty5AahpZ
2DruXpvQgmTding1BYd4va7JMHC/6xNC4c7368VMI6k5Q+n4oi0BS1DDJKg5Tadz
CVPKRCVG17SI0QPH429P9EQgreoZElMhmw7KuiaPvblWF2KNVuYmcljUslI9kKYr
iUPEQ9ceZVYFo8WbjLDjajVYSFKrmF5PnnMR6vx/xIhBNhkrg5ly1QXd4/i9dUvF
wlOFCj3+PlfxCGK75pV1bAx1k89S4lQbavdkVIUmM5ryyOM63nH/FK6sqwJU14rK
08N5KDUlOHH4R3Js3+79L8AeincBs0E2bmNXZV0NbK6zb0IF5twDuns/zOSvtthB
E2KNPCCmRofJuis01/wwqoKdkYeFJ+qJvFAsBUxjvjISnjKMzcwSfLQAblYxDMtR
xQ8z+2lWp/zvian1rUtIyxHyzB3gyhBPtigL//lN68flfnzLIv5TEF5L+MZYU+VB
zb86eKmDMvMEvNG1FBo5cX9nfR5pboNONZ9tRiE/sJ0VMC/V8RboUjoQykzEHD/T
W6JkW6d7u6FGzwU/gx5t2XuxC1egs2gkJXEES8Scj6QtXv6uIMMrgoMMO7oobw4L
1qb05G+bclco1U13E5LdLUl2ND0b3ZcHDFAdwBJIcSRJYNy/IUJjYFX+MVgL6eNt
REZCbMaWpoC8Ad20XYcfcYBd8O0M9dHrpPLld+pTOqjtvdz8fS45+eYrexeCAd5r
xMRV8ueIwt6dM8L0/dRr9AVbBzSkGkcuQwaiHAidtgQ03Wb+9iHULE5tfyIORzDl
ZX+7zeB5v3btEpcPi0ojQhfPt3LRGmJM5FaRSVK4ppDnMAfKPCMnwroV6A1Mt1zk
QOppnvfLlf7biwRVkJ+HhfIh6CQ1XTUTh7pdgeGFPwjamIzQtFdFETAIEModHMmi
KCY/Ysfw9ZzQIX0ufu9lk+2isxDWScBVnzkRey/7G1ej0DuHTX8tK3AbdXnp1IyK
6Tl9j824u6AUFZnR2u4ZXbXS2Ufa/aHaUaLFJDOQk+i/eAwzqPzdjEY8f5x88FNs
Ex9xQGXgTrt8daM+UTVfsl6N0ecJV2GlHzagXm7taD1KNqOZtT7dv/+qIhlHUpoH
FDqf+0Tiw1XzWPxt5jhSVLXUijeCiO3kv23USMNytoAgiMVJ2LXFTLd9skufPEZN
f34nNgLhpi1xwjZmvsW1o9CNss8my+bs84o3GUKOTHs96+GkVMgCoyXesBVl+nC9
Enw6pBQfGAbgi6umWhep2QsweLNhkLxcndB6y3PW43dh7paItmTsXvkGvE4Xtd/w
Two28bpdEzafdadGlaDvJhLFSZ31AU2CdfL9iNMKjpt3T+5NUHW5VTwgNkGtgumi
yCBKm13Z4cnjQGJIO1N3nIiiwajLoXU1cK+SDIG/lZsKpBBwSu87z+1L5qA5SMIq
XpeVHD8Pl3Ttulqep/Bp4rJO+bEQIvmxIHmBy+GGKxdRXox15m3VIsXN3UPYmYHQ
ZQZNCf3Wjgs0llh0t/+seSU6zCuu9fXLP3TxfHppfJy7hUtzv4ij5QMR3moHxukH
4n0R5l2s4o464OVPlrwawDTRRQFnpKxZkmIMuAiC9SXYsszRz5oWFR6ICVOcpHR/
uYWWBFTvg+feAHb0asbTXpUyxncHEy74mnn1FO9UZFQEW+e4mt6OHvVami4uw6Ec
ZZtBf5hAv0vX1gZj1gAtbgduWyZkuC3b8ryVXOP7mwMQ8A+RVDch7UI0RYwuBFH+
YnGV0xb72NaFwAYq7TghnOiHRzmL23ANUi9TYpmetSNZR9ZMSRAh0IwJDoXnqMYJ
hv9OjfE9JuZVgNz0XMtmZrcxJ8KL7PAnF6NMEOwwgkPpEl5VzywfMOmPQ2Ok6+9U
3NlrdSY2Jqn3ebE2ilqd09igeG2m0KY0EbeXvnIPDZgfMcvQgJr4C1gBns1032dP
UFGiYiYvrqNct+DQ4Apg1xufKVVmc6Cdb9FOD6yD77AVKMxuiCecsrYvZsbS5oTd
7exoodqt+V+rRq8dEEmZ3HBGjS9z5UxUt4ZVAnQ0qhmflmyGFFabjUv1gufMHGyV
//GjlWI1FCjqvHgdx0k5DYhWVuzXjdDTpxUnVTYRtSWHMOS5RfjNjivKFn6cxW5O
mANUmkTO0ao3nN4wUUBE8oRlqn5KhtWNGgBpMuvvgaZTku50y7zJtjVZxqWWDEWs
nKRUptaE34bqXcLkWICnJtslfXPHuyQMWc8PGrBMwuYPQM3SFM9m04yzjrAB8xaI
IqMStREMo+rqk/1MNqQ5CVZNlhRYGxKREA7zD0exKGhYaWQyDb9tj8TOF8uhQ6CN
URJ4al/DpBgZCEi1+MA4/et+ClPw8iWgz4WLklXqoizFk7/JJRRfD2+MY6+O7JWW
I/7rv82MvdmSDlClkE+buNEvY2xGUhe4G9375UPljZ032RMnx5oTvOrvuTP54D+5
xy3HXW88aUNk2ARegx2uHYIqmgCNoTInWojh1w05e2tOxY1kFrbPDF7eaWZw+oUj
fQkFqC5FLsA6xoE41wP11d9Pl34nAWkcNAvrflzQHT09T555KVaLKj02+KvsrfOr
VItgmv3rN7+kPfvIATyO9kPSyR5fmVvKMLPuJvOlfknTeJsSjmoGH2AR3tYwRjLE
MKPrYvWtxlTxQxWNPrl2xwVWNJ+PiZ6lI4snHUvyBaGsHbQCY0xxVfe01C+SO4Qp
Mc0Ky9c1cajShQI6CFT9u3Q648vWJ0XGjEE9bq8KsgjpmvxIgPmJyuiWOj3iV6XH
tSNnvRLyb8w0sU63Kq0mQlAnn7AQwm843iqkhMGTDcKi+6pA3vYuQ0YXTai5rlbU
BRBatw/3L/nrI3T5FYJ/6J3Dst8DcXo9ClA+UK+Fxd806aXUbW23rimSrPGYwc1E
WOVSWVGyCYpg2IRqLmuEUD4I/JMu7dzrRffvKfn7COldjIwrj2lldEBJxT+naUXl
aie/Ipb6KQQGoU4k5TGHl2zUBNK6zwCCvBFm4tJZ3IRDWqXqomzXAsrDgWk5mIqv
SLKCyEQ9KuGTtBjHxGooeDqe/KGjlx2szG82J9RCwT75DItvhE4j6PZ/G2uewav2
pI/ckrZSpt1maXrRcLygmjP10Rs8Ib+yyDbAXzmyQBin3kP+NEyfV6RHcj2fBy2u
zWzbhV8Lvp/fd5yCUEBjlZ36J1u3bUw7+Nmu+Pk2KVAPQvxLqkxHepRX/U0X8V2A
2olMWLBauHQxPWrwcUMZQzaKj0YKBPto3P5SZHehIvomk8ZWvhVmkFnNYIepTpEh
qpisrpx8FBskwhI0yyzQerskAfz3dWZ2s/JSabLQ1fjakD0t9sqHuIT4oOgLJexV
85ubVRxrwFJV43mJuAyizaCOmU7svQMUQ/39egJZAHpwYTaMWjQAPJMKrTOLOAkU
VUt8p+ua2mU3fcmncR1Voeg0Ew9ZC7SUYvW9AuKG8ENAEWvqFZWMEhFH+x7L6wlq
VSJ9q4n1czbRwJSe+AWDlqHI5eN1wyslQ0LLZZpmA4Wlb3Tcaol1A5rlva6gloWK
ReTQUHowktjOyI6pj3I8DdjBkyt1c3OOW/OBNQ86W0WSlKpyWSZs94YIxySb8HxB
vg9xtqPW2z+aeyyFx0YpDQPI8Atdo+eVlt1YvkK2rSGXUwLv5FXuhv9utMawdItB
bItnyE4rWbFy/BcI4qz0BB/2u+To5fb250nVg2/Y1Oe+ys4v4nyLPyvK8liXBwyR
nqYAv3wu3lySO3Z1AasaDL8PoHvial+35DNe4r4ZnqY6PK1lIID9W5MOOLoNF7cx
8rWd24WjQ4V2fBwQklobpkMthioMgJYstfoyzQKDlnlscqzTVEq59krNW05WV8fW
cm1HzWXiY6zNadyn2GfDVQl3DA21wFrkJZwJOlFKNU4kE4z0hjCYQcdJkWm3fo/I
Nc1MFs++fCnMoXRbRfxAnGcwdFoZrleKEIYqs5tDNZGkprxK/b9FnQUEeGW0xKF2
Hv2/8+EV7A6wZ5ybft8pnHON9TvfKpDdiaMPQ+5Cbx7dWY3w0DAy/MsiSsFvOs+D
cu3D7v//9q5gJqaqpIOBTBkbKVanPe9qcyKE6HWCWy1PGFMBZ7KJcqVDjuxbt6jS
sPbm7BZZfGAiESyXtjtBbwMhI23ESKScnsRqbo/vnJ6iNVc+3JMiZBRs+P4vRAYl
uocMpiIsbnb3eO/+HVRE2hg7A2SLbCUpTnDK3pw2ehT0xghfQ+uVGlZFrYxlctUH
ppkQc6NsNVqkwNm7ZvVEcGphLxMvBcPWb+aV9Gsu1SLP7BryETLO7NU0o7vRPhx1
5VfMuFhy5mQdnxCDATGeEQj8Sdbfk7KoNNwz4h4moPUqnvHEoXOH3Z3HRyCiHYxE
W6vhsMO8Qh0CD5rvIjaEunXEYzwNeAlku+hlTGBEiCInemIzfXor1RVH/RttsmEV
JZhr56TXJyeVC1q5b4ToEgUmx3rH6cgu79UiSJJnBD24LaFyAhHNPIsXtUI/Aj59
szYnImihA7swhaTCzrL8NIpcKuyuYO/6Kkm/57ZeFrdTm7PwJY3KPzwB6o4pNxi1
kgFRvFAF2kHgjBeHd7cSL3btXJYJfPv+4uD9urx/3dgB9S9TJBgwIOy8DjlU0bV0
5coBqieWu6EebKl91hTaI3e7jf0KSt52zhzKCN6g6i2ikYzZW6a/c1Pdnr4h3WZb
Wt/cuu+dfm2kHyEP+DlDv/2/BK+TJikV9SU25GolIR1k5c2oGgI+NAwjQybnRx64
OZz4yGC+tShOuMH4rJxdYlvk/sFjDJomEe3gL46Sa2PenQR82FhJoWBsRXxlhgvz
IO/iGQJ9q4oiXFkAK0/CjtmQj5iHlYuzojXNVg3uRFS9PfmJY3+9y7uNVPvkcSfy
ZSM9vEHk3PQs4w0RqMVLYhdTQ0zqhAOltXQ1cKIj8IJtUkCkHIiMm5DH5VRLQoF/
xsngVQqavWAkY+6Ea4vEtm2DYpMt0S9+Gk949B7m5cf2kOn0v7nEs8/2TQhzaEnk
VotgdF6bweyQx6mzWgXDiJWWAnOrV0hr8YythToeWe4jShuAAkC96+8tLbNPact6
HFhonnFzTUC1QTYmlRKaoBMsEXQ+5EyZZZtCUvNey9PoIpk1qYwfAf9i9dQ15tjO
AbM4kp8fd5b1Oe5MKIWzJmHVTuYCAaXF+ZabqLRQ4NyEjflU6i5ctQGyr4L6wPio
zh4zIYrPO/mhBwGsCEnJIY43o9cI8yv/IbItuR7RCKcTJUqjNaz5Mb/ZBVr4iBu/
tLO/Zo6c/U+ajucxbiTQoDDaSO7c5+K1qbAki0LSPovAEYp15Y6DxhrqyXSCS62n
2bONI50Te2QSwnn23XuXNrRDhxtnp1MKD5/H3IiRGzCNfzke9iNTlg+0+GBKuqsM
0LLGJ2EEzxs0KYe5GywU4921fBe5ftFbTJLDt+7mQTCrWmZdmoFDu3zCgqURYv4v
pE1N/vV+Bcte2GRKUOJRYUw2pqvOaD84qbiPQgppZkxWkd1bJRALs1AOLLIvgRf9
XHqzJcTKL31hZyFBhHKzyPfVpiwVIuQqXYD4adol0QJ53JZs19mL9LXlxg7NlOH8
pV7x8nIC6SqwlbWCKSNt+6HIDNt2i6zqQabqn5Qk6IfRAcrmJnBQGSXdF5bIuBWh
4yIvX5Q9VuvtQg9GvtSLO3/WqaxeB9+txtxI6hB4+uy0g3m8klQlALaleaGTYOb5
psqXSmvvC4eyM82GdIasPj3XTDbAPzjIpvTAftWA8pKPbijNVZehC9hBcvIggoAe
y92MIjo+6ktyJZBWHzHJKbhdQSY4JD6aLaPPKp0jZvDueI38jM068084+5SxkZJo
PWsgE5XnI3rSW9trOvLMTdcpNrUOO9Kup2fIURgPQNLUuelfFu6fft51atgphWps
TMmR8X4LtAgYixcwAiKYdtVFkJSMBDqVMeS3oiuXGLlpX8UEaMd9rhnopJkBruhB
GMfG53KyvyJv5z8V5Kc2Y4zv436fHFCCntxk7M93rKPOE4xvqJddl0ogKhboYtd2
NQZpg7g1G/iDqswDqNO+oLn9BR/yokpqAY2u3MP+2ZgYlmK8i6v9bKfAKGvzF2+/
/kPEU8FanlvjoJTxazLiSwq7Di1lbJa5Daonp3dcyEgfVkT4nDqqYYQVENDQ0mje
Cb2M0hycVGd4ckrFgaZb98A/TMwlb8KtTVTMeVgtgFAHiHCXj94kqzn4Envw6vMh
3qiDi51Xjaqfh0DmO/FWL8OE+eOpBSqxeoubn+WeR1j3uC3CZ7R6izqsJ1Rk4DrY
LHCKgu++MaKjrsneDR5WJ73CNBOKbrRUpe3YFhyuvXdqWqYdYPDVEPmtyavraRrb
aigdBHp15BZWC7BKfDoTDdmLwotBZKSUHlQ2nBOpXAygSqAzdDffh54WYv4rnRwz
p2Xz2yeZBwsSoWUCHT7c/XiMazBdSkfx0xTstJTkx/8XwLGStAAJaD4CyxZReoMI
1Y5LPvz20L77YLKYY/vZT8NoDNppyEBOzL+6280G2ciPuTJTbuUiIAZXZBL6F0jv
IOQ/Q0pKrgPnVkSEezwHkIcSNZiqBACWBzhF6n/cIucBBUDVq0BbhQscFphqCCbs
KIYALatWkX9O8ioMwzlIxMadfVejITngdL9kJX6xBBHrUrabtgkpfa0Hw3lWIL7C
s+z6CFyXdPB7lrn6m5j1ARlRJ2A2d9emmZJ4Y4mdflBCHdL6/KHOY9xKiwOe/PMl
DBr+UmJ9/ZyQIGZXSsfAC/SCNaNoGaYQGT6tKKfoE9FGB9SufQl0gfYj8DZDmwdA
L/xeB3wQguzurjlNtq3Nx6Qrai9pZLwBg/XttsZuhNWahhikM2oQABA8WrDe0iic
PmckzeRlomRyOWv7o5AJulxyoYbyTCHBhgQgAGvCKuwWU9jJg0or55SKn8PWUX5v
d6G3plIQt+KnOcVOjMSo9LI4oqZTtk0jYYD/6IXohBgDpUYiWJmvPXcuUsF8dqpe
QaVNwrinMxUOuawwzkT/TUlCBIDIZY1yQ/YPpFxAtgJDlo4FAtivH64BQ3ym/yBd
u9uq7uRu239Kq9GJTtTD2+3ND4T59RTdRpYlkXV7ohfh6BAy3DfZIuL5msZ8J2qd
KEPjtdxIsOrH1Wc03mCCYyt1Qqya0kd+PJ6g+Bga5WNTdCxJnCoM7F9S9IpoCar6
+ccWXEZ/cF3XazglURlH7zuMMgaBMSx0H8eiRfJG6wYU/BDNaDWZCzQYMy45k+Vd
U1NS9GReJRUhtem28etEhICHebVn5kymcC/CGNu7ednMGah9BVoB3FuR9pHKbjiQ
CVsBfxQC3ARz25M3u5xgvO7YDMr+6iSHWhIIU8glUsj48FVqNyRZwtUS6H1epTOl
Ej6rR0CzpYmYIyyi0jaGQiFyOIUsOhTMV4EEt37dcffpzzN5wv6WX0lkIgjhHnrQ
eLdwX6POYfXm9sNLJezLAHhiynngHPO2CZ3ysC/QJ1hQuBjCt71hA7KEi7ht10p/
KoViOIZ53txx2q0pcUlly6d99VT7P/4oulHgL8rKwKVN2FL3scmyy1O6llT6g0PE
Re02Zym6DYrV/LTyZxaHB+3xfWvu7J+qcDnGSBCYQnSCAX10vJWIuSHqaDf8eyN4
gPOw+A6BRxd0I595+xVzxv620W/WDBy24M7gb8r9vS9mBYCtk0ZJV5+pBZT9Piba
+WLc0/omVAXHbgFvTeiCqZxiOBv9uqJ+2SyB54gwlbM85FCTy8CogQeCNLT/s4Nz
uWiMdK35NjL2qw7pCjUhMwj0Z3Y32UGYZpODAADhO4GLOXTfqCIhZ6Hz4O4gbCFo
WzO8blsgCesezjB4CpIB2iTojfTEPKgVYidbn4rdRX6eHKNWUnz/alIir2KzzFJd
7pfB13HIfqzekiLNbnCTBWC+ifq6CNumsYQ94lTTTwHSrmFp0RploNFHB7Upj1oL
NJOT4retWiIZEAfNdN0+8bX2hmUN0Avz/z2X1BKmTFZOi63o6uzbD77oDnbOtjsd
BUzzQCEWvndxR5VeXzGxsZbloA0Z5OpG62kSu1TVtNdZaYKBsmRnsTgGKWDf2rvl
C4VRJm3/aXXUTnZObz37ukVfhXixQWlUk6jgLY8G8nHZrd1BMCl30hoIbMZttDJk
E26XaUM8BPoVtndl63Wm27IgTVnWllfGh98i6N5gQDKOarAnqfMJdSRw7VfFh1TP
MMyaFjJm1jJItxEb8AN5fFelMa2MGSYb4MfIml4o7BDYyqeaw2BEFMKFIwNovho1
T9bTXcg7z3mYJokBnFtOK3umjIQbZADTiK8T/axe1oLzAZZpWVSAkrHDryzWyJCs
Vp2dxTme54etbwYHbFfW0Dq1IBYtTgA2YEPj3zte3GoVXJ7SneZdMGWj0H6qU1Nl
5JMCQ9Eaf1BRly63pOckLlkAr7orubGx6n1feFg1+xcCjmyUxmJbP+x9aN08hWVA
/+8bzcFs/ELiFQULD1A/RlS8iMxLc3mvkKQeaMApSB5HmD02iPkIl+JDTHDxR/OC
6g8BBBQQD7763DUSSCIXgIz32YY/gTrcKgmyBzLQIYyyCJnMXypuODCAtfUZnoDk
So3e4R2toO9pI7GYIhEgrf5eH1uvmRc879HF98id8XwmOeFKv479b44RZNviGxOx
t9QsVa0KSF4B/ZzjFStDbf4ZoN1pn8KWj+bQ9qLC2IbAVrSC8oXnmC27nm1usyed
HLrtK2qUApcwfeTz/B6J4u0PO9Q2m1h72DliiQK9L5e+c5KiJPdZdj32kXXJSUp+
21JMRG30kVYMHVNsUc72hSzWUwM9vuIEMnF/vV2c9uSLtHZH/amGxVr1xhk+4dcX
HXjQRITO2u3iO7BW2csdkjEJ0MR8W/5D1tIpaZHatxxCcu0YOrawfwQGbdlz9MeY
TlVeXyX8OLZrnn+JvIIpRqXBTe79a0OCv3r/X84Qj1GMrngNyYWZGk+w/OuYy08T
QiMQpB9KDCwjUQNNUGepK5zDJ4qqYm5EgtV9VVDhQTPRMOwOuOR1KFtA9G5pfyRi
jUXCYzF+DtONImw+v0QRNGwOeK2U+kO1Tp21cWREWyNGyIZhdO7w+oIbK2pzShIV
ufMlFzBX1n7MyvL0VIwvr/piG9CPgzZpJbLg8qAe8M17lSYklRprvhWOn1dAIOlf
lt1xale0zYAsVjUcuihT1urHkkCnS/Zr8AoS115eoG23Pn5oxjMCE9fxfeHzyrS0
p2nVdZJE6TAh8g24zJurWDS+EtpeapCe360lRnDia2JTEFywIQQAL3hRmaIWr/Yw
vnFBEjdbc/BocCXlzQJi3F4HSHJse/QRcX9IW6pthJ+/006i/oF+WEVMqB8szebE
ZdakLL2sTfNneJUMc9wDd8vXwzEkYt9crCONYS0Lov67Ag0/WPNksD9qRo+R89hF
EexSRf61ANm/72lJEYL+MBOXOicRkHC/+CltZr665TF8HUdwTOeTI2CgzT1lCckz
kDk67arvO41mkso/YLks9/Rp4YU+Hk/K1ybpTM5ej94PIbHg5AfbwIu7NCVg7YRd
nQu/YFHZpsYP9bj6Ed2vtI8OXeWVbO8G7BRH0m9AGJ+N21Kpu5Mu86uCKZ7Ga6Y6
CMez3DqPZd51QkCsy6Wd+Mtz3LT86KAXSjHTST/DzGCsfjZq7PYwixOW9WKCPEaC
HVMhrcgAKuZo9QspPighrqQc7SCtIpe/ExbOtR2+QjOLDMV9td0fbRoK3tbTNoMO
dkNrA5NhD59DfLDC5+HAsCgBuFgrWWKQiDg0wRzB9d0ZqiZVtlOuinz0OAKObbXK
KEvp0AzLrpy5yPrNcowX0rHo6hJuHQgOt9FuSVKtuwz++X3QfJsCUlBYVVXfe8tr
3i5YVAFXHjbidjaydU+IlGz4n7xOs8P+H9HtZqhyac/a4j5MCd3BZLHSTbKb/Iz0
O/jE54rLv/J/VRsesi5soPlMchCuGOF102QYwvec5TvH+T0OcKocK2RLxAboaxB/
Ly9uoC91wSQc+ni6Nst+vY4hWdptZtWO1+v40RC9TxfFvv3Ojz1qBlRSawuFwv+U
AIoKFcbvYo+/sNd1OdzaU0Dv0lYTjMaDco7nz0TJBCU9oxAFQQeJb/vJIz9qiVTR
bLdv3SA1eY5gcgD4l+SHEVPpoaxE8JDYdLbHfUAZBrOMS6MzcJhEvAdH3/I1dxS5
a1u9PO4cBIXu665qJ7ImT/9r+DDHP3FG6+lEtdaH+5Mjx3tHJ/i9npKI85bE5f3u
C4jMdwFRnjsWeAPS4920SB/+VT3LIgCatKRcZ7u6L+BzrRYFMskA/98F8PazEryq
u2d+DUqbNcPl+XeMv7dcE3FQ04fnwC9IcEU/Xu57KS3ofelWVLNfXuLby6YIDUOB
laIZ5VgkJ62YH+xaShNRi3VDgiXC/TwY3qZFYpO/Te4DoMxbhB0HNzsVLyOvp/mC
RjYEwQqSdfDVtghiRwLMuH1KLiSUA0XJ0odQlhmMYsH2aZDZKpraDSabDGgxDGp0
NL4yGk0d9hpDFXVVax/c2Q0QjU/YydzIkCLwud/LBVpiwNTLnF0RoRX/fCyJDp2a
vGQrb0sNJpsFKVyupbsZzsm8jjixUQR4RNyXCGcitZTqPB33AuR5ahBbKP8fmt1/
K7fvf3kzxxWHpk/gH8AUSFcGZ0AvJXvy8pn9+3z7aJve2TOE33zPPk7S22ZRFM7n
OxOtGQE06FQMlNbPjtw7UvJGmD/JqmEDPC/jHNs3SP9/ZIOtt71V9gMNCuywE4Mw
vHHce/dNCbttKxfUdT56albNvobyxZKVL8qfTUHHDIEc+ZN0ob38/4J/Cuhdjbs8
y2Fur320jUflzVtHGp/qSwnlw4CWqULWMvkJVkYPAG2C0h++i+pn+0ro3VA2EuS2
ExinSsY3Nq3b2p8zs9dshIZ/tWnPNsRS9ozcUj8+o40upukK2jn2LYbbLVNjF7XS
s9S2XdpH8mY2MIuQjkgzrQhroSCbYh00jdhS3k3nQ544v9k0/XcMWfToqhXMoY2G
oOkgJuvW1bcW9j4M4StLqbRBCbBsx2xr9pixha6Ir4AHDBMwpFlHOK64gi73bkhS
7IGHxf2TQkF4AUUS3vmHvS3sGKZ0g12Wa7jQofQp9qKexuQO1H3/svbkvwctwy4B
gXKhUIp6wibEl4/cddPE+pAUaFw3YqxPGqY9Tnl7duKfx3N/V4yLfbHsij5+qCd8
tkM7jhFyThXRnaEdrtiRIv+NHTGkc9NOpr/EyR0dcR3LSpHGanPLzj0ztP9i5lyY
4zHEuf5pOuUbQGC8NaYpU+ghHyQZ/aWo3K4xwqvFNbYb5HWfyymMAkiYw+RfSnKM
IQY+1InciQMhYE1AL31gKTplwhx1JFRoF4dvJl41efIht2WVBELrFUCsF0HPpkIx
Bs9TiwwQbtX6IU59ePVjdkGMJTiHMH3XVyqrVz9uYXhrJc5FJ5PnREjEqMq2tDfp
36C+fW7ncby5oKxlQd5HprnC3nU036XN1M66GyQBf1C6i4Y7sslzroDhhQWioPX8
oklfwqrQyAz71l3eMo/3RGGw7hM3NI29YzKaY9QB7XC9Gacxge/Eg0m+rC6pEsJm
+D0K8Rz3ys0pyepCsO5/naEhsdOCTFYMWaqZNIggdMLw9XMKDIl0KyI10woaV9js
t8KBWbGM42K5jXFs1v+hSpRgeVaBYXcmtNLCW/sWnan/0E6AqnylRmfWlUS2Or3L
1Q9wfR3ZWregzY2mzhuv6Y/Yi6fl4wXb2zKl9ENAcuBev8hAzzhKT4qKpp2Bp7Dn
GVFXtfDutEhbJbkrNUD3vit383xvjFHxV9xBCJlvl6ZbkEAq6IQgluvAISEaNiX0
apHLKXKp0aiwWrk2jGYS3CK/utFR1+RH2Cb9pZqaI4d/vFiNYVzwMNePsFKPIc+N
ID6yOvnEGVQlmHz/0uwe18BB5dmIBFK/h+nW85RR0vZ6iWMmp8gkKpkwrFWTVn2E
ykW4EYZQEo2Nn7H2wcQkuvfGr4876uvDLJ6Bdu/0sseTNkZ0IinwF7fyjdmZPwWH
sgld24d1VcXvTiqBf4mGhD/SxH1CzW/IIDtoLQq9mhQ824+RnjP/Q+6SMEdOBHm5
v3Zzq/28bI648HQUFC6HtYLvuPbt4xBXcIRXRq3ZUi1wpyqFtAMZe3fIJGiIsWLv
elm7FGxIvdLPHX4vdHM3d96SgE+Tf/ezgr8w6dJb8aJg19oPHAepFWTOTKQuBDBB
6zc6eu+qC3qXCqU8T0lc4ypIrKrL5O4Csu0uH4dNlzOWPfZVOKo8GC0uaJaieGpO
b3nDHc6YSHnBcJ489Q+D+E4rNygkRYSqWxsAMJ2/zpTEq/JxVwTL4XLKY6Bj+c9F
yr+KFW6HCTHj2DM47WmTG+yDXOf4w8mIkQxySFwTaKTOTQGdUjP25Pwq/CxhVFA4
NyevgdfdKt3wnV1oFEkgkSHAIan/KFxCX08Hqz1BSsMl39vQPM+SNi7XztJAwZsC
s0AeprZScQfMBaLB1GR1XZO+/5ouq3GgejqhMb2b/KhJqiDnGbGks4xJGb5PDltj
O8nohm5fIWzUoFXuFAHfQ4cCcB7C/2z1zlo3wsH32AXxrdWtFuth8EmAh2HAi6cW
R9PbBwtLVmUqpygpB5w/aPUxLc/eGFRV5jLOuy0fiZlXy/8ogaRDMMbx6o+rYzaj
FoiZ8cpAjB8Fmrcpblry+z+1V5SBJDqrhpjPUIfmVfcR9aYG9v7297KJR/M1egDz
oeKsJW38IWXcwiaJUMy/ejum5oGDg+dCpOXEL12CnbHulwFYsInTlV4zCCj25AHc
phUdH1d04mBI2GwEAwpg8Dm1NmRupEV1kA76l11gM3YBNRBec1wO+2gLLCZKXtfe
yefSklzv5zlLWQNQag4G40ICJAiWJcmYumOZFM7u+oYKKzwfvdFUg/YQB3iTsXZd
AKMi/cLdpHUuKslw5gBXKQMp/ayGWWUBsalRPP1bPcsemMo8Oq4O6m0YF4CPvHHG
VDW9TBNfwfAqhwmZF44C947rtkb4A2inqfMGA/2+gWhwdJ5hv5XJwl7UYhL1Y8RB
Zwz26Sxp0SUuhOejWtLC2u5kldXNssesiBG5493xvXfD91PUp8HhQu4cCpYtzkln
xX0E5oWcOaf0gIvB5nconJPYVdaHwdxdxbT3uan43NLhAmC8oGF98vHhjz61u4gQ
5pkOgfneKx32VXrHrun7nSMwg1UB1E99dvNn89rsFYYcp1IjAY5dz52lvOluTTzJ
XNAubHzyAbpmLhUxC2JztAZzZ18pwrnLLn+q17ccCc0WCWJdK2I7Y/mS1vzE8Lac
qSIxVRi3OmN5CPmwdQich0CozXaLfbOlJfO+/guignzW4yqt5KynawqkLUpSr2c6
oyjUcAljZtKHM0PogZazjYc9QFUJjU7maca0HCkiTsU3u4Js8Gdu9+/GOsJibZRf
vFG1flSb48/ABFQtb/+LLUOesn2yvsUMY4VT5u99YMSJFuf10rYS42ySwuhjpFtR
bSsV8p/BMQRvrUB13016tYItfXqLpm5q4KWod7QvOEGyNEGtWMziHs5jPzZDP7xv
fqiEfxOPxxZZXSNnCvW9FG9jm675DeG84aTttdQC6hceArZf+ORDW71c7VUaGmAO
MzBerBcIhaH6uFfR7OBd2mXeAVh747SOWP4UuuTbK9wV0jznLaapcdZJIZqzpyVn
mhLMPUMc+xEOLGmxqG1A5+B2iRCsD+FH/5uXDVNm49d56H23q48rS820vXuphAwF
rIjC+qJeM8LIe95460P2HNRODP/aSsR+wrPGkvPUrY65rwVf8/01XZtJjXRhNw+o
NAbS+PBpuj24J5LUP6LqzrIO+v+AwtedXVhT4EnSTPdqxf+9/aoSWlXRzC9dWLHk
pdMxKUK8rK1JI90pk9aEpLgZN5el2yuZV+JYBDd+DrhYdgNnZQ2UjPlpnSMXc+Nv
enuvTdmT9egDm8AqoVD1GvzEyczIhLNwpfqAX0RKzACSw2lt7pcGEGKs5IO+oBG5
P6K5lpp15MiaKJieBjHeaC1v3eOCS6aYqj3crG+DeoF29bdP4vJ21bcBnIaoaz2l
+IMz4Jlf3ph30X23kC6s/QBgqnsS1z9Lg9izYDbk+hwczVWHWIK5y4v5ZpVZpnfh
VThngyoLwgibOqrx3yEF5Giy4YuY98AGZrvWb6awxOZyc0NNDPZl7bJ16sMeLeQl
lm+J5JZR7mY84FhwAf/G8oFyTxVfVLIzChgH169fOwyLRSOS4d9eXeypcrdBQji5
VtJ95El9ayIUUe6HmBaRR8i/TOclfRt5KnOWOcI0AqVYvIkfbvaucgfU9dzUIgkk
dPLWaIJGBt7chv4pCi2DYg2/Xmj1KjbIfA4vyrT9qVqXQA5GHz3CdqkkQjcxDtwG
uSBVCHyu/oxMO8J0zN6m4HvYU2UKuXS/UIzr48TzVF9SgGztyHaGL42DR16RDVkt
Gk9lEeIW/VZD8oLkzhGqm8BUncvKzPhVTaQft3j317Sp12OfVt1K56pkWG1Vqu1b
lzfXy/KzHuY0gPGzOh6sumw/XzZ3SekDhPLx1efn8DnxyKbP0EyQCXVyOzQ2rsHS
EielJ19vR1VEfWtxdbiD6HezL4a+jWoWZT2IPtp7eZDUi/AaXg8Q+TfFE4oAdVO6
VxkigyMLNVqjDNCcfjWi964qA16I4UzBr2bblFVlvAaWXv7hDwb0tWe7R/380He5
puPJ6hsc2UptR8itDq5Mq3ocrrXKgk5Kn/I7QRjioPsB+D1eV8dELJhChHWk3lN9
0z2vITbCS3J/U9Z7vlNwUWkLdYVa8CmefKbvHM4AESU1ggEWFyG7il3PZkio5RCQ
LQ8r5sHr3PzfSq0kSUmsAh/2G0px84dPdz9k8DSKU58k/ALMCb/pFJWh472CXJyO
7JmGDvZggmEB4TjWeqi70GpUrFCCuhGElsxsGb/SuHJzAAA8zCYwOp/oqXABrmdv
HPo4C1KTrxrE5QR3HJvCpKmBSd2FgRJBW3U11/dwExADuQztrwlsr5MB3OefpqpX
dLY1lD7MVoPQY0HnLVx4NuuCrMpQf8BXBgoXMeZjkppvhlIRMWrwhJDv6r5oFqEZ
3V/m5SjkzL0EE9Brvu6jWTxrLcwcOLOwAgjsCIF/mwTmWNRTMWImmOSnaQn3uk/e
xX01Q1s3mUq55DJ5tvbrW4frIY4cd9nstZwJFpPd8Tk7CF/goIVSGUAVLYQok2aj
64dGhnEFS+l2lyFVLDNQtcqKUwsyAAPQNF4/W2EGTDglcAqNr3xuUI1W0MP/guxR
3T+8xWbAmkTN5N/2zEKQ5Sik8Zt1usTDxV5lyYjB0d0SceW8Hsp3a4txav2w+r82
Kfbx+6T0VM4khTEtxd5p+02ETjTAWO611JB5C2zZDyS30upNYp1SbzlDRPn4Atcs
Q8umiv0ofk1KLoh0rgOKex9wSHfUC2Apfdts6GPit6AYoB1aHtN4SOV0mRJdXMjU
xeHxHNc/D8YXVuG/nl8jBMDAJ2Pdbz5gLbZbfojXsDwSjVbu1mLkORL+2lsCgD/q
6FeMj4drtEasNSx0JJD/wyBzfcKSpPNQDfWhYNEQrh2ZZSXEYrJS4b/2M1A6FTFP
aAIWwIqxvG8sC4j61IoP1ZeYMA4uzW7lAHPzbwaBqfUtnnKSkz8YXrEivCovRWRV
pSBe3189nMkHrWRHHQDuO6olIpUIT/G+QL3WbN7PqR7yRbp7upqmIYA3rBwafzAP
mRG1ssCVBNwQFPKIX2uh4W9NP1xLSZ+x5WVSZJMYpLG2pPtbvNACDLN1jY+VNkzp
PamkAD71xfxu0zOf1BJcRpiVo+QnM0qttt76bqzQ2ELoTjBKlOUfHa84Yqyw5QzC
l0AAjn1tbdUbqfWnJkhu+Kj8Km1Xz4Knxl8Btm30PXsPsk6F/pDFuTKU2VrzhQYX
jsJARZO9amt0klMeVB6N+LEe0Da/LqsjO1qqPFiCXz2P5+2sItqPX5r+l6rjq49a
p8Nc4sXsDebPrRizsWvgfecWwHDQgRjzxL9YN5oRjYbPU2lS7z+d89o3HvZvqF6g
lexMIsn7mw9ISdZzKhLAOa8XZFTw3/qpGHOn+FZ+nMtCBZG/6eUzl4vJhhWw4Csc
7epf4UD/bfEoltl8lBobbEYl1YfwCzM3cR34/38sAxcrAtYrz3V+5OYV+vVeBKNr
fTyEuDSV6Kbti5boy7KigERJFxVFhOYQJmCk2IPfacNlcV+rbeo+CMTA98kU/hd5
osd9goMnyVNc/jcevSxwZR+ZA+zgSpkLPvjx4/Q11jDtzaQNbLYzVwRRBij8SESQ
YhlqHJUrp2eg+SoJKUJbVQervadf+5MYhzWvUvsOb6l39muZsTvWHfyZWIjMJvF5
DDTo4v+dj1GOGoquxMRCN0C/j6L3QLtCNleaICfpAKRYAKjwH6m4CCKDA3UXyro9
a3qsd1lQ2omaoedL5zEjesJeTGJesSdJWjWlvQuCykUPr6WmHGTAHNxTILJ9cSp9
1iTuQDEk+Cbc2WAkS7DlpQ5+ZwOWZP1ulkZffcRDov9bsTvjt3SdJECt8cYb5jh4
MWOZcFcdMtKe9niwgqjBSE5IT91J32DGbDf1veZCZD2fWZjyjU4BYWN9unPL7jUF
6h86GILwpAbt9EGcMZfR8833UzC6UWhvD28oS3ao8K35Fjz3YiL8tNQiROIl2yHm
uELfnjPHKgXfDmqIyqpIIPq/U5zC5lgtTv/ccSPi2H/whs0MmCRTeSjvU5EdT+1+
vfF0C9B/7SjVTUBh5YtMSscF6dXGKhpeMWCQYH3S7kh51Xbm4W53w0dNyZnjvtrW
loiqZoGjQUD5AVtK1sl7Qf1qfdeGTWP8VkNTfxnnrP9YzWIVxVTBTTq0VMi/k+zY
cm86if0F4wdbNgoKFP+woX1884xdUBkkdbqFjJfzM8fEoVkSZwXtj2Km1+A94J1e
rdqho4fc269Vtxmt1smL/5Ys/Mp/gKx8z2cPFCwtRoXF8rYNUmsMySPGSIcpZFj1
0DWNvvx7ZQvOUrN0vC92hhZrszOdxibPil2MFDTnXDCvH3Df5aVk/3x94FhJbcZh
wEo1SNn5UnrRlXKS9bc5LrQwEMEXe+0HSSFWIR+T4/9yc+XRUciPMQgJ4sbQTOjA
muWGPprb2idR20e06MFz56YpQbQMF4/d2K6rCw9Bl40nuzY/d7dEvEo/HgWBNF0e
8YNeAHtohskk2YHVY3Iy3hqQiD3/jNEhwOzSASwSwXLy5Xhx1fmewq75POu6T3l0
/wRgKZoMraFTZVl73bd92h4uucqcFzQwsoP1DxQqbWTJfLXU8ipdWMhf2Onn424x
N20Mm0EMIVAXUeWCi79oR80NAS+jyXpUE8vF9tH8QlAkUvitt7xhwK4xzys2FHsS
E5/lWPhwEXDjqwJH3oJp9iPdKrqx234ojb2AdnmLg6hXtIMqY0QOhQ3OW2a0xcWz
0xgwUF7aRJQE6pqdQQfNj5O7YJY2Vem5exjSSM8uk7eivuLewL+nIG5ZSMu1t7gs
ZsCrYi6JZZdqGNLud7otxiPXoPu5GY9hhbEihrM0eGo4ZMq63CRqFrzDjlW239SZ
UEJgws+XYeWJ4wS2rL2mD0g+jBbmL2Udf6rxDqhUiB29A1dKgRT0gNrw4iWitZk0
TTyoK0kQ2jnQcW2KwWkHKWcUY1Oz8iCDQRHkNej1PMFtYI814yipaoR7WNiDkVym
OVo4BQxgunwzG14ZQZrHai18W7muGO0+Z5KzIA9lzYWP94KHc3SRtjGlHt23Tz9Y
wBPoJWfpSf8QWtBZKT537MgL+QNfZRocamdChZiQqbe4BJqmAhXPtFiG6bThJNyd
h1HklrxzonTRJWBSVGEEO8sQKHJxP5FEju4XjuXf4p2Da1i3dfEja+PaC0ArSJMU
NFp7PUSJ9VCCsm1iJmbChHm1vh2vRmdQxkROxdzKpLfnXmsmG5/2hzgR7GhBH/2w
tFqAx8jp3EHVggAj4+PM4fO5UOntybAwcDwtLa6cTuZcC39irsF6dfRfh+LHkRoy
yQdrC+f46wo47wVO6mGKcpqv9efXLTtgLdJO+NYqvhZdLiA7hFnsMozZgV7+FPxa
3NpaBSbVlWJWjCOjIeOnT6aoJkb62fxweBdmhNhazD5R8QecCE988qDWNiWkEuDS
EIW7yJ171CrcodBOxyhgkbdlSXYL04v+MEV8NtUQW//Hsnqs1DexqoxttRxYGCYV
tp9YPwJ4/kGXraRMxV9YftrEGbGCyMwuR2jymy4qYUgLwjfdeN6t5lQWvFRUudsl
MS/mUN8fq+ItlfPDwHEoC75GhK/LZtNex8I9gechsiSsLceqpdB0bXoLrls7KfAz
DElp24TfYGWjELpFBe9bZOtXf0IBWtreUJ6y0Rk5/7nfiabYGMdPArz+fXCAOEmG
5tVdKGWdOOLRTpM4hFHtMu/Pkq2tNXPhhe/4PrLMpMp3n+sODuCaRM6dR+p8S3LG
r4Q8vdfk0D01njMQqzn+9XP4Dg5clZuttAjDTjja5aKA2+nhURpfz/HcAzBZYKLi
Oh3+YBxf5VATc6xo56Cz6ghc/E5tkN/nAdTUKfPbbk+2FCEzf1VS9b9vTNgg5agZ
jLORxb0I2AoV0DzufupsVK0FLignEtwj2TnqSxz8lren3hjUSQj0qF5v8xX8CDyD
uCCqgqiUjNkwsHDJ/GhX+1lKXhl7t5rIDvz91cT3crXVXiOPNvEqXmVoU4NsvDq7
oVQ7sO392sVvhqAKyb2sEO+Sv/mxr3OZU7+UJgQnP28evvIzPouHx0aRVDOaOZho
sAMx/2fW1j5bZJ1lF5h7AkKrPXYhOhZWr6FFTknw7uQrQGZbeAECJzyBR4MTOKXO
JPEYRVG9turAAm12D19emoNYZC2I1bP36B/BSP5wab7RbEmdJgCvaUkOSYMBoHY8
ikoKcDEyGpY/Huqv0NYQX9Zhv1nH512bcRZPJ4AHalWKCkr88M3xpMz6dvlDZ4Oq
bxTs2Ox7nJjYx4PMZFeCBWh9JJJTHSpN3VpQZIoBdw9giKc4RmM3XeWyh5k1pngE
jdqsavICxOPDsVmlrhRqnG0qXvi2ehhbRM1ZvjXrabPeNLBJ2DuREBmXq9gbt8XY
EB6f09aPShTaJKFFr6DFU+sAw+RuSvMVCY9GZuN3pUNxZ0+kF1M2+saEun3TYFSO
Q4DQfvwalRhwP4T0tGFTVyBc2KatyeosfKO+QLnom4E2rAnPJLxk9l9JvTRc1HWY
kqtuKW9uI0t+dw9/akaaGkYKpgYUYjXnP3iB+vjRIMjxjW5sxWL92C+FNWsQWP8l
mvDj1iR0gNL5G2GnmvildrUTILHZ2xFZ2fkxjYjSMpXWP0o543nDr5H+ur/HmLc1
QVc+WLbsbHls43NKiPhpIJZfdJO8g5Wo7o91wDw/3zPeugnENDKLPCvkhOXvc7/K
0BBRS+vcqg1Ab/kkz9NWPusRhuHrRPogS2LbJ/s8XgyqIukGlNbquHuh8t8OXZI6
IJ+aiSd+EBDVoFZjt9hcranFcChtF8P+ZuaDpatIuY8TsJWVWwrZFf0WVecwrewt
58VsmR8PBilY5pPZEKea52COSUGB2wablzcXgIWz1pV6LFXTscyqNIdSw6uh52KR
3uWUn83EobqPWtZmqLnBlN5wghnqVsp/xgKNNvvCvs5Bc1drK6wzrUI4ka+/RtaW
6trz8jHtLyk3lXgzqP8H0JooNQBPmJv0qhu/icGWu/wG1QVpEt5S/HT9jPK2yheK
+Cwli03mLQ6VLoW9+gkio5r7rRUOKxa9j9BF+m5wVZwNySI0hyJvyFdgiX1zeCjC
FoHpeBpT5W/WBpS/vOx6/HhafZ2CkPzTbQnilU1t7LVS4kI5JwkCUO+K53wwW1Jg
LT4f76l5fT/yRtd5m/WlxlkGnp/x4fy26vr98CRCCOjBnraaTi/mpOgi+2oCbNfy
aZ0Al1knS9qQMNVIq3RVr/2iFI8PO91YObR0GGd6d6DiwuWWL/DHMAAe9LS4zyDT
leW5OaqFSrZ5hUHyKB7cMIKlY3u8TgTMuj9+iMxOlXmtJP0Q5FOJYhF9ay4cFEhv
17MmW5VUSxe5dahChGtnZRGY76Pg23J3nT7RZW8XfhoVw23WESSR95e7RzYUkYN7
kPz6C6+S/aVkrwY4X9ZFlcBDajLmNzyr8GRO08+TMMSkNwNgP+1g6aXNADq7vY7N
03IEfNYYrSAW1B1ZbVRhfwKluG8UHdmnogKBw0XP1F5z2NuMQ0kyYrFoqJBYApBC
WJyjg2BXS8hSAf0LBauEm2yHFOn0kvYLGpFItBGOXVu5WB3kGj9qSra+/NGYwdTH
wGZrmf4c6R5OjwE/4lWtIwEeqgP/4FhzOOhvcjsLxSFbpCrnL9WAut+BXabKdhW1
1SwJzOUZ16rCyhFdhM3rii2QXtJFCTkA257UgT4tSbHwnquXKAyBEUOXa+OW70jz
xJi/1c3NYHO/l7XEi/8GlubUMjh46v8b69EqzZzqRuqbvSuVm4vEn9dHOXxysHEp
yp2IWlc+DJIdGnDLLHxhytnznMOW4YG83wAntBBGcYfIBg36+EtrfDrWrcPDaCxW
GMIn6oMNvJKh22+LkcrwmiW4335CKWaXnwuENFVArRe2dYSwtnwRO2CU/h/ykasz
+8N4uHzaBmpgfeTTIgYkgz0KPsPXyG/JBfyqn+RjMVGgysafVCpV0kj+tyIkuq/0
c/7XmT1+JhySQribR0+ge8BqdCKsQxPHFie8OE70NUAAh3kgqtiEaZOebg6THmi5
LXMYuL78DO1xDd/3e/M3ZIWTZhD9WOF8VG2D6I2ljcdXxnuHQtB6N3eIBJHOfXkW
ayZ/3GzvWXHm28MFumJnmf/8SzpLXLzaVDXPb4CK9iLNFNPKRgAdcr6MJh65lqAi
XmzPOMnovfYJzxzj0lhUYWn/WiI9EelDDnFbD7TqFL/f3OdkZyTx7g5QlbiTXsn1
SWnK7O7xZ1BoTNhe7xwUMOGFseipIZLuc1mhgqisCo+tfDVvDLuXCyeiJbpDN/oN
dgezTIYc36NojYRJ+RQyVOyRzaOOZJnmTA5Y3c44gk4KDNuzaDFmLAFsguUCCtqB
qKZOb3SD3yRsOdcqRuaiCam+3Eh0ItxZuQQdN/BpSNwFhyh27bEdXhiwgMuNVSCp
9GVmzBrxCLqt4R1AzJe6bWFz22IZU1iBUWBDp++oRxBn+YZ5tz72MBwsb2dsXfbW
2rJ9AMq6IYLnF6ioA61mV5AFPvVnohvokwZ3THpoP4DY/kdRaYyPppjlgcuwFZi8
RIVxUMjHR9H9n85s7t+ULWfU7LMugafoG88zG4W21LgfRPLnrkPjpFOljfMw4PGg
gE2loutyfqDT7M8GNgTeXsYxHFHIbDC4V+vhZYbvfFZQRUSiISiQ4/lZDRJHU+tw
jkM4Oa2ry+luBAvW5hMwn3d8jkdRSpHuTpozL4Vpe+S1sYSnp1O82kPm7SYJ3FkK
rw1Fg8mrxaTCYOWLH9JsAzRd2r7lCJA4KvCwMqYUhFQLvAmEwah+9IYHSuL7KwYs
gEyPx9WtR7OF5u8e3fePsD3LnmVGhqwyCpBxO3+Topgg9denlDYO9TzxuI4eRkYB
Y78fw3SSeqb6gFYaGCt/4GTmlBT4r34SQr9zsNOEEhc6OSvoV/rQhDWEzixeZLJo
RmFWkpDFGe5PUeOfTS35/Cyunv2AaAM1HPjDeKoVj68PJJAFYMSWoQAEsogwI7ZE
DPhLPkCoe70k0oBP5shR62WcHXnaqIzfjXyTNjQsFRscoZVG0jrVl4sH7AiHfoqY
kb4SJJdiPljIr13iLleedOyjkDLrgYgMtd+RcYT49cOkSzcsA+YWVWQWaHgpPat0
KmGWaGG9UiM6yqkp6jNL6CDO8DQ56qGMBrIhJlmbS2BD4E9PMDM2IVvoWP5RvfsP
LFSNGNya0sYwXJNGtqndQJtQbXFjMVcNp3E/IX0yAPZINIJYATRuGNm7af1n1iay
AgVWRkvF6BV2J6Sa7ZlYX3/zmVyOewb2GiOi8XyoVMnuuGZbaYXpmgOqoulEpMYv
1t2NbMDvodh9H2/AouOeTu0m1Yi03Nkf9Sn/E11Cw/Ih0yeNWXphuQy/NZM32Yip
cJnuwoUFEYA1oAW0v/UYbd1zl3x2MRAViEsn6TS1aErwC4GA9ydMigtClY2E9mbc
faW1ajdJcZdkiY451Aq+j1n/6ti9YNNd8wMMBLKTSnGguWlT8KRi6nLzeb1pStKi
bacTekZk0lKkZZ0jcNr0k7WRc/NyE/6nVCPzgs/FLf7EQ/UBq5rTeas08D+nGZ4w
dfw/ckofzoHc3t4IBsZYqtQ+e8a1IRDRaHWowqHZflFmGwcPvu1VKgrQWxHC08/m
SSiSaxDkIX+XrRzDHFr2QYk8lVKf1W6kwADY4p8Y1YTZ3vcU8nUvqKXwqCgsFORP
HxG+mvkWkKOW9GTZXNBmg7vrfDwylwpPHwWG3gkFRjQMDV69RUqMj29WQ3RFStf2
3LUfbUVX9AO0pBxWZPdMnrfDx79MdASbcqb/rO+GXDE8FtREqIcMbbgu4TLU04KF
15zFsTNB1NSoaKi/RqK4px+mQdjZ6CxS0vG5BkrL6DvJvl4GTGbGZQzHNGEE6QQ9
DsIF5DH7SFDuwhru5GX556Brin99hR5Ayb8IAmLb6cmqfB1GzbSEKw/M5mo1/lnU
zHx/mxotHwyrkf88Z8oo6dC2vTkUWUVPKDJpkKMYlHdJAKCtpmTdhm92y4fFAJml
FhpMjqlhPnULGW64fUEdzht8CyJW96QJLtR5g+ErtGjHFshOqD7NDyuXlLwAe/mI
S0SnfNI5btLFKGfEqE9Pan0uVc80uLFhG3aGe6OGvnrx31ZSK1Et84YFzPz3R/C+
Xbc6WnLV1r1RhY/NwZbklHfYowvmLlPvYkrRoi/AaDK344X8Bmk7iGLNBk/ywf6l
WbqZ6MfDXOs0T+uZvrkz1abQvcYoz0Y9eLmMVN4Y+oU4ZTd443GPNpilFfppgqJ+
9ep5LAY/0x2G2LK+6o/kxRBZxvf6iHxp2P97oUHG+JAHm72UOIJpaGFRAmk+QRh5
WSytnPt+nSA08XQmowCnTaaaZ+KdPGiMIbJs2CX5pOrTHBrUXs2I5l5WSIlviSL1
ZoDX8dMfp+t8LmJi+OVbR37IU9wDUBVgv+NRIwP19/SQFAzYM2omtp1yYVZ5SeGN
mr/+M4i2lVus6blOkrbNkKO/1Gtmo25cOBKABN+MWQbeUJ1fHa9YfmVL3I2gxHsk
o9D+W8pDn2q+DmYZ1NndhCJgQQ0pLgm+YbTIOpITcws+GTsxEgVxNjkmjlcHwOeA
kGGVwB1yuXFzVwON7CsFjUw2q9eP/gcqLFY3KOog/Fvc0AqxczWYSO9mFdWkXUqW
MrqVg6/QZ5yq+1UEnbrDrieGhmqtNQlWa1TLkxptVYQJs4QKeZlSKMIRW1bvKxTx
o0DebAsbYI0CZSthIl6nR5EMrnJTUaBqk/wMi1TfegJUiYWAjAYljDuGxbRtnCqv
kcaO6Tdk5bZmmOiABupA19fPP0N8x2k95hnX9xujPMGNBQwmxc827/UBMK9+M7HZ
e9PZBe6gwAkccQ3Om2wZhK0OfdgrAz6Jzx43tp+ao7JfDPQsYf5S3a2kLzF+O1cz
+qM4b+7LjMq1bjLq01ccGtFxt6d7Z+Z0WW//vnRL+s1bFbjD97c5ks3yOg2AKGBn
xkpXcNx9M9/lZWOozMlg2xp+Frff6wI89XWCEQ3AtQP5493SPirLEbKyz6EmU26N
WYu2bFtVkYMzusHMC6YbEMeSpAQfmhtfBiykQXc4rRRcKdvex6hQb59CHQgvOpLs
Uy4v+QARZl+GQvmcOu+ud0iDkbt9m0/I85IpzFIOlKMRI1P9qkyWeC2/Ee2ToaWl
ti8qAb25Ssv0i9e9PEb87Cg88d32bxbbY7w7DA2UtnUwU46d0XLHwQc965VD6ZTP
oD62VBx3W/Q24xt1vb5SdxlElERsjW09J6YaAMNQMufMpbgXoRudPImxabTjl9Mk
rmHHgstX3sujFY47i+vw72XUi51yRlUcXkrPkF0jvSESj/JU/pU7A9dgC5xOvpYE
MeAvxJMAhpqwpGT9pq9YYhdxXoFr7nAGbJ3YBCDy2JI24/L6SNYHgppKMFYoAYXz
QVZllG4+tNRJPyIbpM3FQU6eqBBAn/5y1H6KdERfPGDuZC8tP01L7A0c7oqPOBXp
7cP2lJKOvmm1cPduhjm+W7WoQqtKy4M/PeSQaAfa5EErZ3uQ8jhxeazEtoouA2GW
p84w4zu/DumQbE26q0yKzn1do3jIimkO/bFXpzZd+i9GfZHllLW0j2k/93uUZpfI
UPekao9BdudhVXKshRecrSNmtbWJvD1t/yvpJRyNlBqhhG9SLJNAdXZkYGE+q0HN
CtBpteIs6I4e21/VE8nTLpoigdgLYGJMH50hIUvZuHNatLkGQC2IPyX0kw84LDlB
hrdYBH/UPq9/wCEG9RtqRnVq0Qh6pAuqClVbFmpT7CqVgVwyzmLNrlavozBKiJPc
Rm8deK6p5vxrFwo5EYiy58Cvr9ha6H4pHYTzOxx8hSgzSClFf7wVQRtrqQhd4fdv
6GYgG2QIQVqIoesWytKxI44kLdE36NsL5jsTO/rnshPYvL32p2ayZjWgWhB/uE1H
xHA6Xvug9eym92G7RV9VGhXaVpPvD/4SP7k4nLNJmUxl1/jaqjrPPbr0qmFQSqCZ
B1khnDlEWEUfdgP/D4DvgyUe0BYyceMLCBb5Tv5pfzGY62rO1fZk1bzIfWV3Fly5
Sg4kgLmG4eZigHQrn/LZWdaXo1wbXiIbepysLYOzI4yv/oTXk8qTmgDP3OGzokF6
SX8GcoRCY6iwjHgzyDJAAZHrmj+aYxbRl6Fzyx60ypZ/nK2+2Ry1HC9CouPbINU7
+S/WTSzlLWF8oe5Y/lJyOuVkclXRyLVN0r1PWxa/wMPcNV535fC/rM2s7BrD1xuW
L4GXnaefzAPBt0QLWApvPjFjbUYrLJrNuWShM1HIQxwJ5cfzwnrBKN2yNJkItVqx
RMlAZ2MX13/zIjxl7bHyuQIrwf4tBLmYsjpIKzu1uG0YrHTSObr5Su7CivOuhySn
CE3zoUVCtQHU5ko6yiT0OFR2y4rz2UEbYSAURfx3fTh0YgLiUq/cJv2Ku3f1njf2
m8GKrDWz7rfW0tBNrLpbeBfdCOIMOmSgw+FdmOQqtcrszw5tjQYO/49faeuckYiL
GwnDptQF347XO3aNuCzW2pTmMDrMMdm2AFtsCE7N4h9TW5SOjzfl3o9H4QmYDtCp
+xJNG6+GoSSz7cdLmqviQCmnqT2rAy0InpluD0i+mVMqnWH5NdhCQ7AeZKmqDjgn
v5OeOEjUHY8bzjdbDbgopbMqHfPM3zz3PGLyDRXG6YwTgfjjp1zCNXykXSaEEjQD
H9IbFDmphj4dtNu7CtnG7mVlEvJSMXLaqdoR3IQ6f5p4NXFyNCOAOgAPeZq27i8n
up5retqe10W1VC5jlVvCrKi/XIZwl+kAiMw6mYreGDGJngdM5l6pfezoI1uB2Uo/
P53mwy42+J6oeZhAIULKHCWbFJ2Wc/pZvF8mkIQLWTCLjA+8nAnBxWg+bDCaXwMM
hpltQkd07PUfvpLN3Emw7NDo3ITGmGkPjjz6wylruEPVbqSSfyDUnJWAQUsyG6Lo
SdVcmWyA1KJZCvp7cIfD4p6UGRROJjPMRoNf8ATGz5mFoQJVVqyLhGesJP6Z6SQm
HyeL0Go4BkbBQz9dkUvOTGHfhy+CblwZNfBJH2Z0OSaL40/MfKqmwsmwqjiCCS9N
U/8XF6p8CaEwC9vkrgHjMfYDYSWyadVGuwsZqTyeEsxGkLMFpWI3n8gxOdX0VpF+
TeXGjl3SblFNcqW++XmUO4zDUTqfK12nFzBXUyTqsUMlfeHa9K59s/G+MHJJTo9M
zJAKZJYMhx1zOhQazk0K9Eaw5uauGIqHM0a2nWr9iGQvtMEOUyCBgves02Dfuf3q
gR6xkP49OGRd1vNC5WqdcNoUwEzCnlrvYA1hvezSe2QvUY3o7pvAbIDdRlM2x5dE
QEDuMLlFTUgv0zJS3/KYvsCyESJlIbREMlfj/HOc0Kc+p+S9dIWw+zoxLA5prsF2
PiWuLRf+oc39g4PAJvpVJwoyzuTDpKQ48r+hJdljLPYUe556Mo3DfSf9JCblNwZ0
4PwotByOATg3cgus7Tb++ckSXajm1hSJW7EVoEyAk76oGP+AyUnRrwvkPIOW9h7y
yrh4y2MAFRhMgXW0I1VB1caXhxeJ1YFM+q/5szvFwNAk9HANE6vNRt2U/3XKbqVZ
9/HHwnzsohhAxDuWbowbwnbyxLR4MCtsMgKQwb3rGxjRNbhoP5uHv+jHlkoORd/j
S/XXTVgw0CyaNITdim8W9cvfQMjRizfjRV/MekBeh491aEaMhCWqDmbQ6GGorllp
gFXDNDhqNwopeQgFXdwqyAosTXrNpHMJUjLZGTyfcUz4oyecPd66WPuFOBFStA6e
Bb8A71kHmFUlreMrC+9yhRb5Akk9ZyjlSyMgTnLEIFeQm7agOFD1Z2m5ytthkCsK
tTVvvA4vkKuzdad7ldnGyfpqP+70COOmFKk6amGVD5v2WfwOeLK/LeavK8t3HE5Q
M0P73wRdmc/sCjJYIQBzWTrRwXV3DzC2u/VpdzYZQq+bUXTuALDFLd0bNvYShiAR
V6P0uJomLnRFBBdGWFBy9AJZj5wctWOKeE5nipDcCJOvibkVW5kUhZH7VA60Qy2f
SlC0ZihuiQQzmUi5VocDKCHW9vgVoPJvCiB9BCLaL1ntXxBS1+LklPCa3kncnftm
cE5cjbttYQDRH1q3THaebgQliooAXHv8hijlucVaU5DtS82V5O8CopZyQA5itcai
3tIgjsE0fzUGpLjGDOAD8yewf1+upnpmlu27lmb4wOe6vgONZrnzj3UqHWgfm8wK
PXnIJn43hXIKg7sH93hFSPmHXwcFf/V73biV5YZ0j2K0OZwvDBI2WUrpxlE5XuLD
SDw8IyzSbDz9mczxr6cQAnIGyJSp4sDNspU07nwx68H8tiCgr8r8YelK6g6TBy28
axOcg+kzQ9K+h4r4g11Oxe2bgBOCuPojaBEZBX2QCowGr7m2JRmu0SOolPWQJOQS
n9aTGuglcaP/KlnjsZLgrGKJ/dcpXKb7elixKoF+whZR5WNu3kL6QrkFuwod659n
lR29nXXmoVtpzMfv5m2avtOgrF1SJHEdL4spxz1bjEYo/bhnbh2m2AXFv2W/QAJB
KyOuECFTYPi5X6GJFSxPgnZEUiT34slvqXCCk+DQTzWJ8d+mJurSGSwZK2WTU3r9
0FbEYRPhdQYQLDVkms2ychvvvVTZQqDXZs4r426T/9NUZ0GpoDgKWWTl5BtLIQQu
21pnHoBqqXdyYrHOPFXt1UCq5rjLJliOeJLXMc9uCEUcOFNInVKmGZf+XeqCvHTB
jWxVvuP0QvQUmCxZZh0D0dHdkpb4/FglbmTZ+7syTY2Y9YV2IgWcQgcVeNMp+Lod
NhGP+LPa/qc7HkIo4/b/WEm6eYZGi7dbva837+hzwcCuW6LpkjwZv4c9i6rzHsq8
AYa+0g8H/l0ZfLolllY2nbbYEpsdyRkS4Akd/EXdgA0mB13vf+cJ7CgynxgmCPs7
5SMlYG+lr3ng8Eu10yYCk9yXGB02xWgAhEdZwACv/eKfwmsRNWvXcgH/vUHFJvHU
RkRIr6+10Pg/KOw+PyN2QeFEhioGhLByOLbBKcOjXBO4xBthYZvbz+0byeJxln5y
52+znX21/yIMNm9rq0Q2TjzVkuJrvYM/CETyvTDukM4FEOpsEXfBbAi7+5P0RzyQ
FcvVvA9ymmH/pC7yQy1dyvLOLJE1lukYZSEXvVIjmSM0Gcj0gd5+hSjo8jG8Fdt7
56XU+//ThE9aKqFxrPOrbf1NPCKqevvd9CjMFq1fKf+YebpcQrKb1OJlIYktTZQX
o60RyIo9Xn5Hp5c/4nnn4gG759aS6nDyw7wovVOU2o5qaR//lJzUL7DemoslPOyJ
5zP8aijDNELilTdX5jF1Mflw+AvnmRWzmfs5RpDQJ1gC1WLXihrAYGjDVRuCx3ME
Ei1Uo4Y+KTfkpJq8+j6BvXlxMrnbv3Evdtbj9b5Gio/C+Z18gKFxUNixhJKfp8pO
kz7lcV820FPfnLS/ZUG4a4AYgQCXc1BL1TQveVYwbIv7uJNYUHTug3fJIq5QzjYY
9FTjO437OnrmOHXHrsQZdAJIe9KVATImGMQsLQWu4dBIjKSYbnAT338QyMwhhPN4
rSjSlOpqaWIymENBWCsrrs03wrgU6zvjDU8BxUEw3koQvNvpj2SdFKNYB9jKLE6R
k0B28UcR2bA2ygSDM0EYBCntyt6TQpQ1QtB+gpv2ctuqnr1azi60/ZrpvDm4crj0
65JKsA3HPaTjLcVqUCWc0txoLM76H50ohUQJMHtDXuH7rfjZVH/kdLk3oqkUKH++
Enz5qknuF+HOLpa1dT2dtPXhKxMkzutVog/dXaLuC3ZObFN7bK11XvhCpdSTFjku
P6sswgmTsKlwlsVSDMD2aiB/n1oKXyCz4lHbt6rWnup4EMIa/MycfPXMU86KQi7u
kZ4/TLMNXqDOrrc1ghD8If+/OIs/uhyl4AJBuh3ujss79aPK6pYviqmWKte7tPPR
2iGPQG2lkvGdI5ITLmpZJxzcjOyI7ONYchingiSJhwu7xYixR5nfhrGYCczB8f60
v0FptF2lc0IC+wtPL8ff25QBnl+ow1+BFk4aJbq0hIUEAcymXBXn97nKBvJWUvp4
fdEXKal730lF0IN71Uz+f1D8xI9xIFP4kES+veyb0RZ0uTObHlXshe6o6qf1bElk
6EFZ5UEsDbJim61MxeZ/2P/5G253zWJzcoum9ITzdF/mXFTvx1QbOzJRfmRsSSQ2
SAUYYNqFnisF4T+uULPLpQKycWIKmJfsvIwSVMUKexRS70UiOoWGiXrtBBcIFkww
KhXuGvt5HYvLIjZbRT2XSF/h6TltjAg2qLfxbKbXrUp3oLsc+uJB8hbW6kwI7o0P
VvUs6Ko/8Sz0PigHdxHpb6IV31LVM9pFKRpCQTV+h+dD1Z9TCFPPaXYb2i5ldDMf
nZxVQ472vGBktgN5uwFU/o6fvu36t0VrHStOuIULwbiE0a8Rkfx1R9ycyyED4wNg
tpK9yqXFI/YLFpGh006UdPTG1MwvWeGZFiKrroxOftsR6T7KbS+hnBcMrDkADEhe
+x2MDWqCrNZ3Xp/jJOphHjat5en8eGqDYqbyl/IIaC2QypxbuSpm5OangCGTDMMz
kU6cF7XRjXPTPk8jZ97RHww3snvAfGYniN39quoGHoH1IZnICWoMb2+Z3exng0gb
Q3cEaV8HUwQNDiu1jDq91B2PjLobGxzkczDTchOmTX4zvRIAGcxXu4jcNtxUyaAi
Jv//l6eFu0JvGNj/lpENjj/nKQ4C3VJV4ePmeGhnbqozT2Kw7Qi8FanbxGfulim3
nRTGBF4gDT6uayXjSGrZDCcQzYANuGZNvrENun1oJLICLts5F2V3buxp7OgZmfZQ
pucQzunGLgNQyfyxF8TYEr81tk7ficVnmBa2Swdg5aPGLSgoHdamJPMAxMnhxeag
/FPrbs+HUI76z+Lnenysvu46Jai6k302a/auPBGvI+EXfEvQ8lnmq9fgcVgL3jM2
X7okH17B1x6vS8h4UQbNLAlI4guxKlveK5Gk4qgQjyBRQHH/S1Dc96cfiEcokiFM
gBSDlNKE5fphGHvIjnrSUz8x/xvi0gPj5u14S0/RKmAFnftvkeG/As4DkcgQsn6c
7FBIoWXS6Kq76jBamOfhZh2QTlWKT8Dk+ItUgmNuaOZJS8y/Rm+k5ZYBDyDZV7G/
NUL8gKyJrvDBThnwfeQUP5pfjzf3hgnDGxdvjw1k6uS+itK6vQVfI6hvsGAJSMua
mfHE+E3tKlpDVhxUGfuZ9o3kKyrArsV+WGIZPNoLfcwve/96XNZHcEwIJKioxpXw
azrOuCz5r9r18XA4paC2jHLs5nvZk1EDto2ornsROTVCwlWx5z/VUwzj/8N5K6O0
+lnnn3HPI9+5sYXlnYYdbRQKqx/Hhc9DKE4/Tk3ojvjjNnlLqvthJ8G1adPY9/fI
7hBnmikg7IfM/6Adft1FTu6zMFkFAovdc2Doq7Upr5k/B3noO+I1sNuEo9vriu+c
H4m+ozZrm+r82zCF75ijLdLDGOVlj+xdFLhxenVfMMg03icss/O+WPNw7rJ3gUNa
fviHltFIaWdqXKYegoqaUWbfPZF77lOmzXGNguRHFIeNusbMgL/pdwZtiZTE54bI
HItVasSAWmvyLXyqBBBk/hjvyzPoXo1aQpK26YNldNIlLtMHx05FsqjGfyzV3ekG
LTio/An88ej7p1XURA8pWDjaMdjHu2SWK/CtPR2AvBHK8QIQEReYEkba+aRFr1cK
yXN2qQJyIhF/QcLFRO9N2O71Bk99MDusBWHQpEYF1LsPMI7/eRkB5JJtNosBQAVX
ZK4cUpGegs/f/6tuyWM2JPy1KGGiv5/3qEpfgg3iYTWjwb0X34EvMpAdx8sgmU94
DQsbJrkLZh0d0nOhcm4pP2hHobQoHjNb0yhPZXlSBS5+GKXdUuEI7NpJo8G9G7Cm
Y0WCnsKKtLvj+O6aO6vFQmYlef7BkjXobNBr4WWihkRqXC0xuR8PHFUmDz7o2a7S
IvZ+pW8ixPbxv3r/JmgKnGFL2tEW+jxAjkt6ap0fA4iwM3nYRq/+Scq35fb9yp1S
pZ3xADGZC4R4goam47+1dpA2A84oozKSqtXqhVMO3ka9UPqxVdZITaiOATfFSrRC
GFc0yCB0nKFk7xfm/D97DGAr0sETxaqICMujDgMtygyEzgqKu/xHdLr+naPD89/M
kzDhIoxv8FA6mS+XUUGJSiUY34u3rN6ZFrs2L7NhXv8p58/DqxbGf/HUFyozlJGJ
wakUiwoYls8sbb1gXWlf/DydXZoNwi/HdBCgiraa1MHLAwGYB0AGu9VF8vUmxNy7
k3CPXcIH/QFxkqt2EFKT8Pe7cvDcodm9StNbcjr44Mj/yvOAv1UkBeMfsheSSuvA
B0KGmvFTjd88Mf/Zhea3E+CJaExwOR183bSqykAqomipzOPgpo0Ab8ecOrykuuIp
qg+tokbByDIu4ValBmvpj9ojrtl2zCc2lQQprC9L6PBda5v4ufgbLCuUXELiN0i6
hvr10Bd283cLVwN3Qr5NfOoS+HSmNXyU1UZ8xMh+Stu4j1bt8jr6aLuJ7wSVvAVV
GmMw+gXWnMUMS6xpGE3CKJFz081ZCgDtamTGG/dsGsAhmhgKmpVlPo+uCT3BO3UD
8h6PZDevhL5rgReYu/RHApJtsGrBva/f7hP9uX8f3+MoUS81mcKT0QfA7yiS3cQv
c2nL4nMRMaQ3oaDaPUYMkBImVCFNKiCF0Omd+RcNTKmiqlO+Cb5w579Dxd7eKlVp
iTtw99JBGiMQh+dDAhiSKsnj9zboa+YGdcGDgyn+20VDmdQTyXNgLojFNo2i3/cK
9C8XaBeKvlR1z6lTO9eq7/QsK5wQvNmk0/aMxV1GpvaCCjk/eMucrCX0r1uh+ZGY
mm5/fkMz/5nsz10ecrfblUbPwew6Yt/Fv0z3/EbEt70xfOsHrrZyIYDVNl0pf0wb
56+J/smfXGcIkDkp69owCFRoPYLSoLPbGkp98yXDCC7j/sREEwLGGp4xeHfxy9IU
7AOmAthFaeim+1LRwHRErKzZjkVs3/W27oivkUfj/8oys8qqbNxbw23R0bGOV8EZ
dj7dO0DEeU6dMMDG0QoVMgl2E6SIC+xywkUexYKLBLgh6BnX3oqAb3vl7dv/ENwE
NPUZ6wbpjooLowMGXhXhbFMIyELC2+3IttFqrxTxDnepWq3ZlFCS/hftQhhH0zJy
dhvh224dHl3kYRkZMX2bIbLSeIAmnVZH5kGks37OLD3RAZij+DdAVtrmFtOygZwt
FChzxv8UZ2lLrdVmD2AEZpFk+JIwiHZt91SwHvECeN8zdWwVUJzPpHrOd/ItI0fz
Bl57j4y/xj+2L8OxqnhK13n3aQI/24Sg0fgpn34Ez1joGA6BkKHbv8Lf6oDYB+Sk
xxf6Z+7lTgReEgf277ThsDSqn+aNRIs7hBe5SjFNwRzggODrgNz29FabqfGrOpZW
m+zjiVaSU8USCarF8BL3GBsw9j+2erXFUA7ZhrER59W0Z0GbCdIvRSfntDmoM4LF
h0903eE48JZSjwFAfj2CfPNmEKnmW4fYcy4xotjra4ZmmgrVveDMWYQdKQmwDJgp
WUmNcTTfbQCrdArnvg6a6ewsdjzNQjr6rTDl3zx6QBWZ6hn2n+scPy5Gz8C1ahAK
bUsz9vMlmi7eJsGpQzHUgufNWcGZT4zv/mVDJqv4BgAXeuwgZYKb6dxTt3c+LSXb
O58PGRWhC0i3FDxVlso5v/zBFB34HNeKP81Cmtda59KYWrd5OyzjBwPLby4YQUxk
uZ+6ZSmeYRNX0Dnanem8bvrV1Qq+TucWqMqy1v3+u5Mc67pSLQpSsizXWUqRFi01
YBiUnr9PTvRE+4kEcZ0mgkJLBeDkf0yMpzYkecRfsoyVKIeRhQ8zwMCe8cjJAkQ5
Z0yT8xQovD3CPBKU/LCN4ZmXwkSM0oGUkOxxmfahVFXPMU1nC2+RUYBHAdxlCNjf
fOCuKrd0Z+B9Bg46ZxlynIhaGUAe/KRxjilwGSFwllw9+GkLUBUAo0INV6aPw96L
KMOYLI4e9+yqzckjdjnULfun5j1UmFW+hFbVHAeMSLflEBDUd07rB0fB4+hx1/C6
7CYkk7dLPhymgdKgQOztwBoVQVoy5L04LF7ISwnu3M66qjlJf8a8Zr5f7wFKDE9Y
xXtJE+t9h/mdSWRrPdGA5EpJByUh36GVRvFF7K9QO7yocUdtydRR+1Qy2+GXe0fq
H3Vm5bqi7XaAaXy1fNGOruXldO1pCj7HDUStE8y4/cHABIpNm+HWnOAn+/i51s+W
795keZ1bi/M80AY62mJ0IhEse+xpfDpdlzW+jClSY5ZWiJaotrjuPa3ERSdCSRRK
bU92gWJR+tdRRv1uqiG3HEkwuCd956Zfge6zY79ZazzTrhPJYDlr9nSzYRS9FTId
8PUgmCuUkZD99oLvZ5r84DZYbA6/dS/FOOrfqncWXrF6Plj3F9pRIPpsbojQjWoF
k/ZNaMR/BLO5nEqkiwTf05xdfz9XK68KqGHOMA7Kwq4+Rn/VzkxRyzW0qP4A5rEH
n5MtxXjoM6p2A5+7g4fLgAwj0QpSVsO+nli9jp9PiKs8XnmqaDIn8UWEcINXhbS+
/6pGiDZYYsQDtlSP6HQVeTkQETycFxtnndAX4XW9ikIe24MSCZAb+vXAf7eE3gpn
bCXHLYjU9HkR4hhG2op8HeDh6G5C575b8EdiDRI8dvnEANCUzjwHmCsf8yQyHcTq
gV59t3OEnBFCZVtJfflm8+Mi1PusmUEiK+qFDASJQvGT5FqO17v3W5fyGDW4D4Kd
9iaRD4RHLM26drRmIq/6ex/qAAGo2s3ykt6fTwE/QAqLqC8AEuPDYydCAV/XJJgD
SMy+MzxXhGtQdV75iRfHrzlfNtxYX5A39dF8KNoePREbNrcNJKBq9KU7oqVd4SvT
w1pJzHRHGLIRH2wZIJhwJWMmRp6MLHf18Qk5NTHdfps5diHQ9Db5xJsRcaUZYL6B
wwEonXbpZmN7vwOo82qTaxIGIQPxnIUJceRWqIn2P1c4lTGxk/x2m/71qxfdFRRW
J0LsxeaxX24et2HPZDZaszRWUAGy9qdbtuRuPiogstnnY4OOysKiJECN2bAN19ma
uteyGUnGdcnIqaqWbHi+1u7k7LA7fk/ejR+NSKOQSFnqAWNfSpNRr5ockc2q5Enu
dRxpmPOj9mtLYo4Hlw+V5tNJ3pxYa/6asQ7EoqiLpyJrDEOKPEkR5wH9dtwmW3NK
If5j263Wm6ojTjXV0QdDx/N1tcgP6b9m333YzJ3EwQuZ3lpLOBQV214AV4j6OFF+
W7HORe3o69TqlkQ0Vk3Go39MnNCfgt5ZVMhZxhuzkS75/hdszecGNcDRCaF7+XIm
42gn7X7zENEq/tM2UEioh3FN91enjKF41vqRagwxIx0epgmhfxdu+xMgSRSu4D2h
qnY+PecQh6kNz+anfk1sNn7R7oVFSC4m0gZh3OvJ9nJyYXp2h8cUsbqBf5RuLkGq
voFxTq7TnVezJIeKDFvn+B5WV4lnzCLkVKaTQyCln4MkRe3Isc73Eytg6NMPgRhC
LzPx1jtvxeudArUrYCfRqdv0c17ktJI6UwkOhIy9vtY+ELn0AI+hBzbe48uG8NaP
ZvsQlCOGHQmj4u6KfffwB/Z7FiurspFCL4fCsCyIi99mGFtr0jWVi6P2ytbKVc51
N2Um3NphzsA8nJs7IliIftLDCG5kvRut5h+UyvUeYIdVr7wmqNSxJ/XrKCrGSgds
/wjS0UvFnvLwyNcuo9inWKuXU8XJPnIkB31jwOz8LvvXrk7JPGgVs/vZi/VlZ7pI
st3/fswPP5KF48IA6TgK/5mqD1GdnR7jvX34eIaS5J796CcKJ/otzXfWqhTOB/lp
dL/bXZsBP5cVgQzjH3t39YhdTqYGvLu5Q81h05/+TY/Du42S9+vOQmYfVzHTJSvT
y7QCZ9VHXWGJRTZEiiV+QjVavC2P9MUjGBeUo0ysAMm0e6Y0ATwuZqDh9imTOiT8
Py05GDAE55x2GcBbD+lbzCOnBJoJd1mHp9bqqYC6kcYl19qxIyN+XnfMhfaen+sr
ra7laN1O894jCq2WxKt4Zz8lHFoQYQqWk6dJtEfmbKeGQndBPQFBjiraKqf8Udf8
67NALBBf9ARVKl0fro2lZ8ui0MazVOUmulrFEmMAfqRSe2wJP8yEEVBjl/7D4lGC
W/AO5fZTW80COIKSC/dr4IOZt6/elBUBcGtEN8vCCbqRQDYVDRmrXVXKaUsbBJO1
ujp8jKUQfwjw2kFN7Mg4y7oLwCIIaEx4I2eI2sFRBub0uLa9FmrAzLiONJHYu4Wl
HkFJDD8tI6uHQ9aB+24Vm86oygVyJrm4hPruit4MsKNfGabZ8fgArAOLZkl6y5OE
SRdgpgdq04CUBBcsr5W63hZDOvaATr9MW9uP4B/64dsvNNkdvk/uSFeJcUNxwgA/
IisqdmIK6IzNmyQl9FrAzM8UmxIbzyUHNV9RJLb+DRO4UKZiXRDnLlpVdR3edcWS
sa5y6Y6a9J1zBLqZfW6nEC0xZw4fOwsQpyrj48WnZE6nJPVqbfjkojnFuFQ2lH+v
55oZ0X363gUlTViB1tZoTrWRlj7Q6LHt5iS83PXIaGictuo1de3gqt7Ll+I1PP/3
cefeTXWDre0tt0PaYAHabz03RP7hyjOH7IO1VYeJOqVuM/Rr1A43BLUB/Xf/euVu
ktKBO4NJv8w1c7I8JQwgNQ8RYrTK3Tf5yIyUhepYa5i07rRV//FB81F3+suLjCaP
+6RCn/38hS49JE2oI8/rak+nrjmKgeN5eeVBFgJ2SjjfjLxuwdu+LvqG5u4Y9Dcz
S9zh+MCmQ8l3gTbcCOXTMe3+zQLU8uLLe8AKUzi7uicrw6Iiu0QzxQ8XumTm5Ydk
FbmuTfCdx8hkcERkDeecd5eAuj+9MEnxvCqbmEwan++aYueiMC+v8ndq/j6LE1kO
5ilHavyOEFY/2uqVFYji+syJn/+6pJGcC2ZUVPk1BzZgrwBYelhVPYFBhucDpiPz
ClkOqQKFypArV/RuM6ELTDUfE1pKL9WYS3JD2IE8YQFtWPuJ5MLpcfWZjwJ5KZFx
XeaKS/MaPhLqN/eDnIUG2UuMoZoRZBFkHuaMLSLtu6+fE13ZalMj41qN04h2nbxp
HF+hvu/SKP9SDuJ94XNvRtbeDEzGI5JG97yumgR2p3pOt1PTMDGkDLY4Ux14UcQ0
FiyGq7Cz4WN1LCDtfyraJR55Ct240J8tvVXjuiRO9PEMuHRRrhzCVgBLaaNBZ5yN
SzqyVIWy1VMLmG14WM5VZBy4L9zD7z0g6lulZitgimFHJSk5wxSG7HI1m2k0fMe6
nZVGzXIbveYGBBsPg8SGF7KU+i/hYIwQNFCylYGvg1GSkpdLN6u0aGWcbUmRvlCn
6gtFTJnsk6R2b94K/uVsZVYQkHkFGhGYtTP5m0ZSiKsoURnJLBEbG9ue/UftzbLf
3hNDadSO93JJvvkybVBePqFBu15NToTyl4HeecDeS6LSwfszn17mWOYlxe5xs9XJ
H23B0Ialwu4Z+dNpct27YnvqNaFYEVWtGWJ06f/kd1j8lzTjpvrXqkzOO6/IAxot
StzPW6rNvXBwgLSrefDeZR2ulnQhY2Pp+kSPciAVXgSd8kM+Sql9P7YLH5yLvCWa
0EiLTyXUIzkCAzf1X+KZbLrS1Z6ALH230Q+Q7Q/O7OgXxoMRCrYwQ5p2mVnoMMlw
kpLBXT++RYKNilN6pH/TwhzydaGqGPYOv85vTddYfgqo6jW5+2CpUSQl2xDk8/9v
qey6jYzN9DsSDsq9H85UamqtSTMzZVssXGZ83uT0ynOfqgxpPWZb/vBbTkH5Jhb1
CtLp9RPzsYZqzzGphFNS0A3aNFlNdatxPd0/M8+NybTcwEhtQS0/3SgaQLkV+XJ9
xEGjJkOBuImP8qCqXL5g1QPuGJEmlleKK758kC5cWc/Lb0kbWqpCmHoes2N8/tsx
cCSgeNpQo6HiS/p2WpBQCcFq0gqbk1LvTNfIoHkhQbRZq5/EUTV/vOApz3kxn3H2
2rBwOAZL44laPomKH6o5r3mFPiRjNND67M6DJm9Lax6XQSnajnpzGcWimj5XKS/k
54QtP+4eLqKxrr8NaaxLpTYuunfhUcIbIVljHTqtzBP2ls/gsuShhYbhFGCdl29J
xIfXlz/eQSjUhA976GrdSzBfxMaUMGTiW2rOy6tktp2wmVHkoPsKNLwm+sUDy01C
vHrXufMt54RogZq8W6xhD6COXUdMYcLVvPPRBMqCy8YFNzzRYXnbD74sAYPR4za6
tn/0Tm9hmoVTpPG+Qd95fJRdcyl1IBxxrXoA4OnAQDs3KGl0YOESrBZKCcNGmZGG
6IIzyAF9tqH/bfLLADCDMnKbJCTDuVOrqJzKvXGGjV2jqOHSfvlnQJQWMffiQqvC
G46TpqO6i0stAZcFlfHIS/X6x78YdFUgWtbVsdf7qPxGrhOvaxoBoqq4MLLfAfuR
EqHLWQp/NKLgJSC9XsBXZhUZmti3hZBuU8qCzgaAhZRzWlt6HUZzq50EmOAs1dxn
jqQbOCGA85flK1lInAyKrRKEMDIwoeDHJJYdfUOYeia2w1A3LvTdrkOwEuPYuSHx
n3Q4v8J1n5nUmJ/NZsXBdloGX4b+TBKnbVCPMTU0PCsJstihSRqlpSiq2Xsn1+/f
/7vsfF5EoLFMoo2Osb1FZ2ZosPKf9BNljjHhpmoEnJ8ZSdKbL1JGDMUfkR/PoJRw
z1AAfHldtVw1KA1+jnI9OGGLSRqXiUi5FVzHQW2fyvS1ehNUrgDdy3AXyosAAUmF
T3w3WwhWOnKhEvGcy+koXgv2wk7nupWgZ2AvuV9de74Rf1uuHmwrNImqxxzJZpDl
EoPJqWTk5TD4XFH9wGMAXeppPVckVdm1KSvtQwOOLkHd6O+LsD/dCWeOr26VyiMb
Z2ymC+xxSeF1fdI5TdBZ99GvgAf6123M+lb3GT9NR7btjOYSnieVMissLbyrRVlr
8G/JlFNBvH6w56rOJ9ycecEsXAappgCilB+Ql0Oj3tzuG/PuXtLUewQMe+7ujA+q
AWhrm/hlBSU2bQJW3nBXtrKp7d9hc58sT6KF86zZbGYhD4w287Qq7je68yoecW+2
ku0YZyiVpsKvoyrxq0k52y/ojL39iwsKK+IbN4wa3Q0fkM7McrImgYsdwsvARkME
dKRAFjW49+t6RFdR8yBVKrFHDqBCoYpFO7t55kAUY3M6nPRnm0meNUuA0wdeXXvs
knAPSH6Qh1XOcY6bzx4xTE2j+fmxzei8AB7XouDw+fF0toHEoVs5IxhNNa6ndauR
8ymCTjoAL5RtViBjT2hdVTfdHWe2LTpfb1DiC0fAl2BXy59grX0+xbHzpRCda2eE
zeKo4d0+RuGCxD9cLncfuwk2bxAQPOLZpULIuZDhcLFvbxuW//ZjGl7cLzQJJ9HQ
PDlMCNNFJEFurGf+cpHaERTK8rxw/ERvVX0s4Hvn+y7cSoIaAl6C2XkFyAS7OfLF
tjxRSNsrAVQTfDIINilDhG0wMGFJMD2bfl8lw6wmT95902TZZ99K/1SDwD8dsH9t
5H1R+gnU6Qd/ik/P0DhhRrjF9LrKE7o98F3VbfrP6KGGFh0kHKSjxR1WPNZhvi81
uJvL2idf6hD4JjcSeArvGvgp4GYUXECQKfaL5gci6ZTdWnPQfY4AFspfs9QBOr7m
STBfPWpBT2MwUg7pQp4l4fBKLm+SQgdQQm3ZhDLdnG6W2Lyws63+pAm7rcYK5Qf+
10Mw6kgKRmHoN5020N44AdKZcicsJXti/auNipUwx2REQ6Wu0SV1JdJXRQmw/1QU
bTdIwEUzcUYUyQHopAhLhjQvxx8QxP3ewb2so0SrPKlruPmXwkUcLh2g4y7uqQNm
RtrVlcfF9C9Wt8a0qFkNZxvhPR66Y1LtuGkBVG5TQ+Zuffe/zMJDCYgzCSVN79Qk
zE6Va1W9I4Px1HTVPpIau/CPu0rJAbt29kmoq1HCBRfnI/ZgV0wESCSqMaq5lhMj
f1uK5OSKU8b68hl2edw5SgbndCbNb1dn0/zsALTZUsIzJt9PyCpBUGjh4mYhXXGH
zwwvnbs8qZWdDhy7O0pueeR1e6HUhT8ybGwtm8Wl8ycvsGathPl5xTC6ZM2rIdeC
8HWYE+/o//J2P1oiNki0rmLWzlGmL1XiWB6qhfNeonbrC1+/X6+eaouMoxPsDguz
h9Gt6DC04SLwccgq7Q+XiHaByF89IO/pZDozMc77adR4ASRsRYvx4HcagfiE/bTO
hVaULLuWHwkbqPgj0gObO0/Upb0EEO2V/wkMhyv5jasO9qPsZ9S6c2e0ytDV0ofq
b/Zh1dG82Kv2D/aKhUrQlr8YFswy+LbQ39ak2FEEmtESqwaOLKiszk0fH/1EZ7T5
8yqlEMY1URde/GIneCGsemwUPlQWSnjqj/Z43zeUGdnNT/0Mb40je0E12w8CQs3O
LCMXG+QlThF2ZkB//2u4pTuCMtIp+TakQIc8JvDldLBckOM3xM3Z5WvRraVQK8mM
3LdSeSukGTpp5NynkDwuufZT3gj7J67kdLM0g86+sSj2/yvqGX8E3MFDUsXgGcEq
+h3qoF9zt4mSYU5P2dCpbvCuX/syL2J5xrCUMVB1OvWneVvOU8l+DzETuBV5PMWs
Aelcz//Zhp4cUrTIGDuRjMRAc/c/Jge6otPLuk4EwwqUyh+3bpAtYo0Pe/wJPZqL
eJh+MBNQPhuXU6bjjl7X0SGUJ2nHSvvekmt6scJ5x9r27nCj5LMPdG9TdM3ASo6A
E3RAjW77Vu1KJN1gX3Lw19vu/r4nsTN13KJ4nEuZbIFFRqwi8jEKYFp1ineEzt4p
/SQRfGUSyYQNO8u3va7BWrbGuYOnVfSLZaH0w+Y3tUPwnUGByNxVIYupJ9hhk/UV
22WRyi67cNb4kSLCiU9EyHJc9ntML4Ef20o8IdNXjzo7Cpa8MblQNgnzjCzM1mq6
tIVHijsca1Jj7ZdKEtLbUoRZmbQKcGPFI1oCYX2tundDmhTd3SKK/dMKGuEXgzxM
Hv3y/wmErKDAuhn861olVFTBDuBfBIoT33d4kGXHkT8+9AyDnWqtHXlSTi8YC/RW
DkNabfGsCtbKHsMRyfnd4FcVKQ57ewZ8gUFe1mj+RFEb9SGRudRHY0ZjLTllfhUE
IPXLS3B0AhAYOf4TJIgaUTidDYAxmnOg+LafHR3xid++7D4YljxYeYbkgyADlNNw
di8lGE7Ycdt3b5Dd5pMqOlVS8rHu/Jt2qOcaRv7nX0myJzry+JsDXopcjnAPbFJG
Gi8ma+uiFan0es9oK9FYVksF521AwRewmlVqVjx5z8OkwtW3TdnMCl9zxFrQgajQ
oadv4UhIL/bBDBPO6NpkvWvAvK1QDc0YnCuXoDIZAIA3DHU9xtmCqg64kUYCTjHx
fBOTv3Ef0Tw817raF775sXj2VUqusx/YrOEfPyDQ+uF17KOpQP3hFGLams3rGmBd
ZbFgxzjzbu1IzTTPvmdppIAT7FD+IWVsD5Qa/MaR2fgMNWCpYifuMe9VmjwDrYOM
O4KUDSP0Ii1koPzj+/fDJFiYzVJZvaBPGibDiikphGgfbsIhhkC17fRno7wJY0O7
hYdeLo/VZGzNjyH6DBTzbk7HIRIP6Dlu6qzU9mltkhwXfF6Thh4l+gByIF7wIYRb
hruUXItgwaqghGuBEqKpkPaPo3uAVVZpMe0ISWSzA9ZTMCAxmqQqWrDXjlRbvV0T
vVuJf/Ow8ZuaKzXBjNHhfuWwjfxI3FMLXS25PwWEKfoZonTmhBmRc0cwpjoDRKo+
2OzbAp+bS1F4HT7nU5xAL6GFbJqxUlGtUSsD7arf06SSORIxGNV6gV5OJW2Trcml
BS6irUhSgccRLgy8vxZu7w0TWMqsAMo+BBvP4J38Jq41tLA4NndcoRptlMghNugE
iezb8SzRByVRSzFmAZl32+APRpwO26rwRIqKmF1bsw4bxxTt0RVmy0AbpkicmZTH
gJORVQpfpKoas2RaHEUGCaOKFimUPLil45o+SPyLqF9PidfoWU+ouaOUNFk2W3R4
18cdFyssFjJrrn+/FO/Un1T4riXAoRCuq50z4Cpm8KzbjLL2Qybqkuc2UvFojaqT
h8P4S4MIUq5laNMJEaEnKvWt6GrbGDlcMTtwiGChQM449X0MnB3R4RtWBd6XlhEo
fvt6xpXO98JrX7Hnc2oQVkjSZNOe/6Ba9Fijbx6MnKbYclH8DHh8nWBphn2uXPSd
8qJmGNlemkYe4QniPKo/nXNeP1Jb7PgodN7utnjmp/IAMVGtWV7Ku7P5he82ZCNT
2bFlfT4KPUTuF1Gc3cDgurpit1A7BEUdrzPXW7xVqhv0Zz3WuOxS3eN1LfnrUINQ
ALRMd83coIL1lJY+Im05uJu+TgG2+GreZ9CZFQ0Y+ZBHkq/6H1OF+HxTwStOq0Ea
BvN/dB/Sg9UZC07NJsqpbeRrYAkgotvyh5T50QNzwdTm8jZw4Ic2k9Ql/7tLAnAJ
hXDG7WDUhPLREl3Y/IMdkF5qnPQDMtKLXCQdczKq/8MvyLMZZILS/apXWlU1XBRV
gs+rtysXO+blAUnLnke5DwdK8JwuVmgUNvvlGwTbTrDP4EyxVOmikpme8nwuzlzT
LWnW2EMS4RWwslFQOlBQhcb46HHCR1wG57w5Asa9YfiQqyO3aQlFq13nZwublpoE
XlFcRGEMef7zHVbMiUU8MsOPsXT1h242Fj04IQZ4iPbi1vBWZOl/vLtzJJi3HK2L
JRu1zB6aL+9KKorKwfccuTZAXkDrzRgxMBvfJ0DaktRnz0mmNHeYc2SrHLPw6UsA
B4P+N02TyYmPWHJB4wbcqaB94ww/bt4HLrrH33hAVZD/3GZFj1xfxA21oA1RZO32
VxcdbI+5EIdYtLly0mxFeJ1BswZu9xrLUsTlO7aSNj4OyLy3wIEgk3lgIVyTtUvy
SciRg2S6fzlXJKQ+aduYwjVTj81V/2AEMI5kK1+dd43wEI9hkMK+oyezWvvZsSsK
p3e7gstUMpkChHJb0FiDn0ARXiczi8qlXWQZZcsMRUA7QH2+vHkM4/b8WGQTir9B
DgjqYFCq5gGpPOJpgK8/lKCy+JK2pi+4uEOjZ7PMxel6mrVTehMB3Yg3DcUHZcM/
W0XUZ0JvQDTHu2NjX1N2VfclOkGM5nw+JxYLs3vO2MQh5SLzqMZ8uTQz6QSZFWl2
my8VP3MrhsFUSXU2xnx07mAB/Nnf1WUqx2eHsJLh3OhvLA3zBzal/mJTa7b+1q+k
fZ8ZDTJLL1ZFy1UdkDHDvaokLflKVSkx/YueOFtwBgDrhUj+40ASkInWdGKSam8E
YBnO7whvMj5jSoybGKn31jC7YBj5S8Wo/1iOWrtD+ZqrWTsMpqhwNkg229B92lDO
rnyckKfaBTWvodPSqMEreMjABRj3Sinm5CoV8lgWxlelWzbPn8ETy14lK6bx0tOH
QSeZAb/kNTEZviuh3UxEX/M8Ex3GG7RT2SN//CmWr+rl6w5BQ3nN+e4l+VqLg2Pw
nknp8KapaSl39i62b36w0K6+u34QbEtgr4MFfJ2VM8MAzmcE2nqYG4d9DM8YajO6
cV1We0/UJu2MqHmYHZlxGgBDS7Vxs/oA+wvgrTCa2qQzauzD5yoVLSy4/X5cnTTJ
bJUXRssm1nHubBH9WrgKtrzPNEqdS85Y1BTuJib2wthM59huKshJxlyeeqxeMjZg
khkaekhZqrY6BwUzxEymJKN8aVctLK0W4W/8fXeJ8fcgDuYI8Ue11r3pZlFDfBON
wbRHngv8cAONBsZH9Fk+vgSbZ1WTg89OIZkPNKDQhpc5vA2fTFcL5OvTWeLSJ64L
FI+7sHY2U/svEwYHPmTcTmgkiAZa8Kok4ZuFgSgWPhKoBmqXTwulG5BreYtEyWpW
yjWTsMA1g8P+kaCK/Gsc8vvEZoLYmRQPxl+hAHlNb1XlMevALt1ZI5sS4XxpyhHc
ccJjI8FS4UXKBvB4mIRRgCR31KZhGsHdUn2L6m5CR247w4ScqkuuWaJP6TR+y59T
lrLzZZnNGM8oeKCiBaDSNDZOQ7Ze4PwD6l0GfLQMSArZKqwa4vRTt9ZIJ6beT9nc
99uM7iUnn0ZlSHGMa7HTKF+mKJkG7HsfWKupMbyxB/ucTpNIREoAA3a6x31hkipV
vOODzLfXKvSutG3ie4kFzTtTlojgZa3XHnlvQaqF8Jh7bXX9H3RcH+SgKoI48Pli
jdI7nk1ELb26/Pg+CK6K8kxO9RyRijUetKbHavyNu6xc3mnEiTcVfUU5rHK86hV5
hxosL/SvPtQFD8JgypbCrZxgnsw1vGuP/G/bohbj22DSPn2v/OSDV44h/rX05BPX
jc0Yn0fjVhHgbNzObWlUA76jwr3clvRWlIjy2Oq+Olkp8vVxwhv02TBdy2go0+Z3
m/0MNubyVBeuaX+qQzVdN4wCMwSCAIZeoaxiglLh087IHg/5dCXQLGhU9WlfKSoM
9aBWTsPTLKJfYmmsynT1haUS/WxJDvKYhNHmf2h+o3zVwS6BKEH76e/RzvkcEkSh
dUzTWWYdBYPxQyNs+6sSR5XyALf3n7VBdRzjlyBs1DSMZ1KDhmaKu/Nco81VC2zQ
N0nEsuBm5sTDjMWWagj8gWtDHeqz/86BqaJ7+zFDNlf67/O/G8JdzewHYoppqSj7
6JCPEjafyEkD6QGJYJPrLmICFAmg6NyZ2gFjHFCQxUXGBnsjCu3Ocur2kgoZRFAk
WH+6SaeHFrAzPtgVGZpw5f9871Jj8zx0+946VufcEQ2bpXpY7/qSy7D43Ay+/IJZ
PZ05TXnWc0k/sSh3F+2qXnRwwCJBeOE6ANocVtkqKccFVjQ9PgkB6k29ggKDgIRN
lWTpktOpGk0hoaEzwkOvKyIzrcv5nH61vAL0L73PdnjyP1JI+nJzv4fKAaXQVvyy
iVnBemoinfMK21UMwVvfHaeIxs5Nub/Q47eBwl3OToXCyJTIM17sxrdlCbNoUYo+
MyVh2xqZhVg4n1AY58LhmyLCV9Sqrip8/SVzMpZHrfjhaRLXPO9XmVxZhQEdY0PW
u3ghXKV6g/Daeg6t77Lk9bB285EjL7IENY6vVeaS6otGqVXDVXWb5m2zaDYovhMk
9Z1GFfGu3qo1G98rpmW3Uxn4ePd6IdWg4wejFAjl9T815n7EFt1z/6duzVdXxZVH
zm8KaErX9g3uJtdGuR1GuHVkNS0ixujlkUcD1p5TqNmFe/wZIE5+SEFMNNBDSGET
y4zd+PhU6FILMJCORYcOFb7EN9rIvHWCfr4Nv42ju0bC8mA6V9C/iZf28r99pBCN
/aHCj0FkCCMSsCKQpUntj9H85PO9WyIwICuRzNHBuL3JtvwdU07SXEfR/GrZqSZt
I/1fel6YqE59sI1KJIjWItV4vBNMvNKfY44vqyiDeNQqcYhiMnPfF058nrD12mdA
1wiYvWnMPl3hHT45OsUmDI8e2a8/h0kVJTHaazswDw8n45oGvwNziEobJNqTlPQZ
89amO4jn7XroevJmgOZXHwPW4RWt74CpYRpXAJcAWNIZJmjlYD8GEyDiTn18xIHF
352svaXn8+vAQutiBalMCvQjcjguLsNBq3mHog4B5AD9g46YF1P8TDanlLw3HqnJ
l9rgVFJBoC8sE34F2RS4pXdcKsl53bdp2QvJ97rYrdKyTCGFKn4XSDe9b1kIrKlg
svh6uMBheWb6fege6qpLeGLWUqxcq0o8UAklsKmAgivI4lOQN26oamBQdPkeY62E
4kfwXPjz41ENrWVlaxFl/Ne9FhzrcGeyodsNrYGE2f05R4TmBTCFBV816QEbpj6p
nIOYtAv92mHNE/5cqpQ75HE2JYrzvy3Loep45d01KVs0YytOoGeZ1G+xbemfKjXw
AoATByZ96GJFTwibL/gGE4mmLv44VtimofAcuBoc4KYGXKTayIMqQFihjjmpDxAC
A8qFWt8wRR0XPuAZFrjzRYhA9vn56GHViUjpWsuWkEDSrN4nXh8YMEM6E8SrvJpO
67ftg0O3VwzzE2hQ2wE8xNmp99FMQmodki1k+C1IQ1lnELv7NFhtNIeZO1cg4JbL
giWSh8o7gO/UxGjNagoMJxP6UrrWy3gTWRovPvNwF+nMZmkvajTeUAuiQ3l9ke8C
KzgBzJp8kBdhZRkhzlcX1CufdJq+0aBdD+KfS5LxOO/nR1RJ8Q3L5oZiYrQwu0uf
rXc77fvNz45sJct/vuXhEKjMYmYXBJ23aTawUTz/eqvNZglwHVJb4huWFORsRLaw
LRRTr4pc/5IHucRAktU5IIlB3gRN9HqE1KPJYTQ1ucdgrmvf4AJ612tUbMK3EbaL
5tdzX1q/swxOvRFPGa9Qg08M1Va7wg3ZRhVpQKJeQnrybYpIXKSnEzyPoDw9NmI8
LjiKMv09cIdrz0S4zzTR5gr7+x++qFQUaJiovhAqkeGaZQORwCZCi2PT+xBDjW+E
SY065gj9+Z4spx98kNCFaDjmYVLOR3lfLO2AJGPPCheQTpjdmgcJI8BzImI29BkH
ckXFpQK7ddsfgNNeInBG+liZH6sIdgVHj265G1GKU4gZTSMQHcpqrv9nafriUmzz
sb6K99NB7goCQk8JO5fwCewkXUobTk82b8k5O2LoLiAd7xPMLqGGOZF4WzRmgxCG
w/OsgRFPVhIqovf5W0kXdDuAVNCyoUAcMhC2SyCtlRhNivReu4rR1MHKs12GWwKZ
JARiIFPHVO+WJpqABQS5C3wAuOUIgQnODHkovJJffsdeBLhDEv1T0iXEK8UxYFSN
+ufWaDHSQAxIJMrB1jpN4rnRkL9ocpzaYcCIBftKL2A93V4FfluUAyC+CMV/b8jU
f7Deb77e5lUyBDO0tXaFHCfz7wFm+C4v4OcywSjV5/odpjcJaT7KPL9zXxRZHMXy
L75KrMWeU1OYmgySMRzr3BHTYxjj15syjMtomTKXtxx/Pmgsk/aKYbPTvZUZMxgQ
GNyfZVFjFrXSFz4urV/jIqu0bECyn9LvidtiyyO18lUxNXcgEeb8Mp5JyQw4lNVQ
ssJLo5nO1q7WSn8QQ7WlPECdPplQlpHnb6TWUnsBUqyKIMsBTsVaO13aTbg/ea2N
rCfYUClg2JN8HtudE5/GzBVJ4t0t2JUtjW1WS0klloyyWt4fyIcx3w5o2MFnASlc
UhnLA0Aa5RVHuJHslwFp9uZzMX3WBTpZSgnnxvRlo+jUGTIqqeGPVa+GSEq4/2Lc
+bYi+qtPOZUEDpS+PViHXCABeZdZcErydnlzCuUlKJRd57ufWnTZMWugalc5Rzxc
hFEBV1st/4FkvxjJFBx/p1CJVi8BJDiaZhdYROmhh4NaKkjJV7PVMFTtgFcyRCOJ
FOfXhI1uyS6eiUQLlptFL3tzDi8y6e/4iQspzr5dyXWXhYdtZLmGGCE/kj3WePAt
go+taS8jNpv24lGaon9J8KYhOFPgLzGMJw5SHME9cwrATQGRDe45JT8eZlhOrU5s
wNUbt4dvLUpe6n9ZZva4mQGDqUI90pUslvbTykoX8R4+Ug1K2yZ3EPdRBMlX3FJF
wjBcT/APHpQWqstsLvLktSIdctqkV5lqi4ebSmUodLRwKAVBIIm9xSK1qO+ocXQr
7n46jx9QoGsotnSbgPa+uEiTJRL73oi9k9NJ2QkeQcExFgXOqPNWRTxEXgQCjz08
jCze9tFmOnAXP0SrZER7b//BQIZ1s4sg2uFwqhQiTS1aE4RV9eGSMmVZflLFOjim
KpITvAhec/nY43N/zSHv24vJtIp6efV7jB21gHYw7ATFoGiqt0J3k3NRcMHkGiN9
pOtUdv+hWyg/8ijHTMCG3/zx8pab9LRung97Jf1GDqzAqeasAsDaN0/mvEPQ0igB
MCuMrUM/xXyks5K5UPnmhQ6kgHld4FV0Q8TV7sE6NSn/F1st0gSQZA2CCBZsJQMM
5+mZo+ZHt28Z8ec1s5HC2jo+ln5nzcfC4j8eES0i+C44EhgJTI01qp62E+mDaOGa
mbdR61pWVKOi6zRWs/Zfemt077ZoguR7lQxTwHvqo1/4r2A3V6122MKnM0NIqquj
uyKP8vz6l7c1sJbf+DwzN5TnL/v5rzb85C1+H96EzkfXCuqDiq3U5oHpF60vYATZ
fCVKZyN13tlmGrdbHZ7jfqkL2dJjrsOlyCXI2rLghxaSdPaUK/lNDsKURixNYObS
MNzHRXo2lQSJcYLVWin6cPiQo2mr0lw8K/sNqcLEy93yeJs4yARzCeFVri5NCdJj
gVQ9H1HzC+J07zRv9zcHSihllEhxCJKrCTqi3RY+9UOFMzL+iYV00iieBHL/GZUh
pkc+N1m/ncz8h+iom7Qrb0MLCl+UuVLFcv8COld0afkV4QuXNrWcpLv8t2iYjqTk
ddUSrt9XEP8VsiDeXUI9naEaoWOpvJdaIbB3OoB/5Dw6hpHHTj6B44/Ad8I3dAex
nLuxcpRvLmdlpTCu6Ezbdnq5nZ9nBsGw4sepg/fvM3OM6YsG8+LBwOaamqsOnE8W
wWZKW1Q37ruHW+eoTuyrRQ7mdnqcPJBeplOWV6sMTtEvX7wbjyLwsXskdwYdqSBL
5G++MrRvwbVrCOawJt1+HP7P0edr9k97LraxlH71H0tdvccWFxFo4ous6OygzM+M
utYQKPJc/al1JKURqEo65Bpn7r8a744G9M4WIgIWzFLZSu/CLgUUlWtHuxXSeMKB
Rfc/bpf2kscG5zXe8X77MKKS0WTSnkgXxg3Xr+p5d0DeVn7jaH1MtHLCyDsU27zg
PZKna1iJbBgzMyST9mJM5JMZt70NPDvTqai3WySO1EIWujfvrAT4vvSg0ruzzZtT
pyVOIJ1OepyTYfx7ti9LJG0qqDICmA/KmcurkIdF1sgDTnO0eMH7LYYJdmZXks77
KWCB5Zg72KZ0af3PH8pfVBtywgKylU+1ozmU820fBOXJpbsFbnpwsi1qBpHQe/9e
PF2HxNC8F1UuuN8+TQ3ORihmG673LlrsfpO/4dIFnYmkyicr1V30JgPsYe4u2tt+
MIIm95m1tVn0TcqQTRqPxNfGwJvTBZ6iyttJBoGD7EWOQYrrBXwcCvJqAimSsgoI
Ii9RArJgdRbqIihQUDWhbxflPuIZBCoSyYXhtZ4SjbkcFxe6Wv5AOILvCqxD1AdU
7UCg3e6HAk/xuv4Qsw3ivKjo0ooa2jhgcqC5fnX0ZBPg7nB0KluBuhuS+MTq4fb7
KkyguzsfePbzdBQgpSnYhJa3QPJDvLxR71OgNXv6YkXfgdvb3AjRfODdmnOH8Tji
ACaPe8c+sz9cOPmy3uNf7MuTJhP1yfDfaVKXYbHj0VhG0LHR8j4MsIZl6I+HFpel
pZn7hgqEhvzM/W/IN50/QxMt8WcsNmjWfO/JVJZE7fdQ7AZrOAzuwlpO0ZXLzqBP
Q53GG8MJ6RzpC3kgcKYYxaKSjzRaSEfFsCpfnDGHqaRJOQZCsQiEdC1oBGvK4k2O
o3ZpD/2wKxIUrwvgPVh2P9JE9QKJAXxxhBu0DBDyYUVzSORHE9Sr0kfAxfMi756M
kd4+ZTi6lEU405e08kteHfAuJMvTuOy3UwbX5u9DyiQVrYyWsY646Hm8bEeVkLW1
Dl/SUQLBQk18s1GqwtndtitwKRsOuuYT5rqyO9AjJhrO0lqu5NPDB9fAsQC0YDwY
4yWuA12dGvL4KWF30KwM8UG4nJtKJpOAeXjfD5Ec37nH5rDRIsI+7QIYJPRdj8Yw
XvN48LibzsoV/casEHoRwi4+QzD6Y/QoRBJP9tz0lout5LNwYzDghxQ+3KeLkyzi
GFQM4gnTglg5PljkDP6vrsEmQu4+tIp2RoPavjIkwGSoCmTICsKdZhafB88WuDkl
wqw2uC6gY9m0Ug5ZWUGZU2YbmH5Ki7kbN8WxPUCJSaa6mkVscVmfHQ9I1/tFLace
QtFjWeaIpH8InHMoj7eIEnCSpXMiGAcheaxMzLxFvtgj3JKOKitn/cc9m1YXazn1
cUEIrfvTDfeiBGtdF4vRu8j1vfiixL2t/rNEBDTNYnpCUr8DoAeOYBqdlAs5ctCL
ZZ3lJ0K40oLaK6xaX+HJobj5dcosN0V6Qgpt6x6n/iK3yF2FoX8vSyTWmK8uWzq8
WQrkbvGILHojLxzrfH6du6f/NUmX/Bcp+aaPFHydHQAcgUjNBVg6YzE5ygBHpL6x
mCfRvm1ADI7npgicEkixEuV2Oj5U5ku03QHcmPjvt0kdirfb3PXcA/MIi/obHUlm
3xNks3B1lSikmcp82mDmsssHbS7VZpTU2Tde7vNBNpPnKc4NjWVCA76R/JC8KAt0
OZ3Ty21iGHEKD163CwVenSXnVLZrcUdtFg8zuKWCobIMo7as5+kzO7TFTOq9OUHA
Qjx7PGmPdlL5p4uy2rhpH04k/NYpH1RLRVG6xPPZBTdK84Ga6wipmN+qp3/qGRZ6
91CUv8Ijf1GEpYbKaPT5J9HA5xRMDdj4X9b/QEUd1n89WfAk4hrvu2JgyBinGzAy
gX0YFTdmF+KpnzA53gtPSy4H8nEO9bgRi33m9kbfzD2rhj1FHijzgUAYtuqa/ODP
Lc/JgBJkLDHn4pAJwul4A/FmskDcRBYhvp71lD8x1lSh60vJ+YvQ7rWmAobpTSoa
5hYCdj4/fPshieDG76shuE/sbRqNI8BzQ1UPCScXhq8N5W1B/zcc/dIQPyuJPbpi
+L8GGTwqDtYlNY/1xqTL/MUQj7n/M3aXS/n2efjaxp9lk5q/cMRSnAOpBlo5kdsf
vai4ZTBs5Q9yu4KRNu5dWgjMY/ex2oPVHDnx94N5EWjYipl2H4bi7cHbJ7agoNn0
ss/PUeuwEOcXuTIomGUmWObTbSWAgg4l6GB8LJoL9QEkqijcAowELX+VTm8QshTZ
dVK9H8eJ6wUxmfhm7JrhnoP4By/eRBt+9rkGkp/iTshiDlZB/o8xi/SbuEZcIWpu
JqmyqSGl6bgYSKdyzDcJV5XDxHwBSCPBxQ1SnJm4oN+OGu3Jcp6sdMpURldX8Iwy
cA0kwFcVvyplQyKgXWTC48Ka3DiGbT5TxUf91D6GOE7etRyyQtHNAMPW2V9KeRxM
C6LsozNgGtb62WaZF0zbWv02NpxNv3otG9hz78F7aoQZ9dFrMh3T7yvwSwGQgVlx
r3XrXJySeYh2MyJv3lm1nzYrU6aEPQ0l+aPZMsQ94K9tFb3/vo40srFfQXW6zdiv
x8KSRvh9H0qipqvt/SBvdf1Mkncc0gj9qr7L6H3N5DzzCulH2RbD0hqsRcfwBY1b
qnO3dau76NBMqI8Qukp+7CO2QvjOLgEs3qDj6WGlyaC6bRzJc0m1hC4s3evVE3or
pmko9BPvAabZbiidXLRoR3qIJbpu5kAtPWRjbxCvefQNmx2OkcsGQg0a9kwOouAn
RGK5+51rxYQ/sv83cNWXxWGpptIuZTjY7CBVpRLJ1jhzJEATym7gChqY7SM0f91w
QFGDY3TFeYCzDlCx/0BXp6IcFXGVBHD6oS5L6YwHPeZJxcGttkmNImtBb/aTyvyp
9nkU+HgedpAQKucQIVGLuaiPYP0OBS5lUHnk2RdWCVC98wgPkqtC4ObhYT5nbBgh
Ue9AW+PN9myWekUg0tn+LVtLRX2Ee9NrPrdOULBYs8cNezpncP7v931SV6AD3rEL
wi+dcNM+uo3nq92AtD7wu89sJsHp05OCZDJ2cfOoPojt2XWuKpDSWlrwR4PT6kF/
dXncRVPLNWfA/hKEDzE23Te11p/cf2o+IwKc4wroMOBNV0G3jtYffXIuVHLCxOa4
9Mk/RJHJROuEP1/oUzhWOHiz77BOkJONJxjxxl3kj6g2L6rSPEcnlhDvV3voeJTq
GTC6ZsRtrXpTJydQDjBE2ukxjdQDDu0pPZ9Hd9za6nM09g1T+ZGd6DrNXvXaQDw5
fcPnE/xYklHAdsB4H4zzifEsterkM0uthASnL7spo/T7WYh+b+up4dqO2YIx7ga2
dc7JWCrx+gb3h760nFHw1lwg3+sLEMj+tjaALHMMDn3SLPLTQw7W4MYp9ZpBeJtf
wWKO/BKflnFZ+/Mgrnde74oJAVrzzYCGB5n6nil0fZiSA9AcKWEspPEM9NcDTT2I
Er4AdH73dvdpP15jdc1O9AJv8sBA7Sk0EaQ8rCTKic9P9YGbBpxEbr2eKnq6NeBx
BGXagGR/x8vDTTefS4hswIVYNAuuJuH9+VSGEh3EhIXAH7+QOz3jZ2uYGPR0ofSc
8CbxUWL3HeyeVyNMphRo/EtLVXeOtvVt3493ml8QIRALzeSYobSEwDkrjJ6kQrwS
HGCJNqvT+sM0AVfZAk5RPnQbdNOUcSK4QFG+EwFmIB4GMx5ekyRpMOPSvp0JI+mp
gRYFHv48m89jvLF92oSJOZyybuOmle0KZo7mPJe9tVMu7iZtt0LONOuTCoGpA99m
FBszXZZL2M7SiT/WkROqYOJIJQmHrbsKf4ZtgNGP+FN05yS2Qg5e0MZVM7XBxBbW
KymQZRFtbRLhqFTK8nfjMdAJYxt0odZ4MX5eNYkrm742PJsCxnP+1UDIICYPXtf6
iElQN9h0Fi++ZvNjKZ5iRunHSSdz2YN6LJJqgGFu6Ai03yH2XhQ4rv44aGHr4LWd
7QzNHZfmvLstNSqEss3qkKhFSjMpmpZvGBTJPaXIuU4l4juAZzxsM/ZY+gHE4Deh
F6lPQ3vJv+TfDw4tp/A4h7JQMqmR6xKOxnl0h1UVH+XGftAkoRFhFfwrj0WTGiPz
hEHDrKG4ECsr5dyy5DWtKvP5+egDcn7zhxRv1E+UWTs7eaFP0zs0rqLfCskrfuCK
pet7kCdgp5rF0lN9H4nPRtAAdoJ6oBDR5OqXt+rSLDuiJ9J6Xsa1zabaxMGSzTIW
6QVJb9+ee+eaUPs6S8HZcgDggY0yLrylU0sEQc6H8NGnoAYccE1SZs1fxr+iO2Qj
CuPFm1QQ72aRmi0gJl6HkANNFhtxy0Rn0O57to80JN5C+sVW36MOPoya0luvpkml
W1ugIisHmtD8TCC7W8xMEgYg1mlJln5vGfR+jT4gra74/Wpmqbg4H+QCA5unfqMP
Bum3+wNh+MuxB6sUtCjTECH+McZKCwvMSMJJfomJqa6OiJHwYmXnKbGquiqxTxmA
IZFACQHiC+XgfepDU6HIeyTTqP+cUAYAS7Ot8yZ8ROcLN8zKB7jDToUGAwU58aMV
b+d09yGsZwPdeaOxJrHVkdwAE0T3mPhL07qYknGstgnoINh4dtG/gSP+YnMfKe//
PzJAwJv9CBSukQsIpiTFGyLYjC9ogBZTLOoyzPmpkShmS9b0tLgzbWnyRWiV8Z4x
xgGFwatoa5UTxcwUdh9Ozb6bICHYRNS67wTND7w+ZHdCF2hC08T0aT9YaE2ZHhM+
S+8EAm80Zr+Vx6yUrdUWDqJsm7pE+JUDZnbunmzkLZR55zz0x381Cr1x1SoH8FLm
eUPQXFgUAMsZ5Dkr98nTaOiKdD67+dmYuGWF7TCxPQFV7C+KwkNKJn6CCVCCKSPe
5iDlKQ7LT/RLqz5luvk/hRTY4mfRbL095KTsk9bx9WRScnCZabJHcYQTGf37HdFC
jL5ktKl8W9nvGAacBKuMu7+9Lq+JsS5X/wZZnRueX4DcPdxgTak24MYC7MRBy7Zn
CQpFtEa3VIyw6EOAr1U3JpAGikF3PTe6ZEyixOlZXoiMdSZIFvH+qU9tFeYLupBU
jacd45Lsjx5LYMaXyoN+miSZd7tLIs5STWt4l8d+CPIE4Iru1M0TULDmKfTKTCQO
e1Lrt/c94XOMlDFRkJ4MEr3JGR5scFWmvduwh5A6K/HWP1S4LjQeBl3iZn9cv0sb
NmpRLG9P/1W5QrEPO52j+0rZKpaSlE+rDqdGOVqteOnU5wPzq2e44VCBf/tgKGoG
p7Zb+prRESya7355Fb3B5b+deGql2dPQJBwbLEK2Gq5z6x6TUX+ZCq0WQqlNDkwV
J1eE9rz7bZz8wMmz+lz2aevF5dUopUK8/ayi7eGbD+dN+KjJlB0WIHlfC4PsJZw3
6totQgO91qARMmFImi7eYeNmuTAV7hqCfrg0v+KeY/EJXXnMimAVpEc6hxtogiL6
90Y05l25Qn5RrjUm2tM+GfXhEh5Q2U/lfMh/9KEn1hPLzt1aIoo4ACkvWyBXp35x
0SYWHGF+OPjIVhUbdqcR1hUQ18mRipW59YY0zgLmvlr0mEWqW+bFrXZz/oJs58pu
+RKlXYBU6Scs3Jt2LrNx/RMKbhm8oz9OUhxC0Z8cAgGMBYF8uxK9FiDoPmB6GhvC
3TNMIFFWmr5/IzE4L5ENqBa16tTUJu/1H5aOl5bBQeYmhb440jdtEDqD6NEG1mRL
GzPCHKNBuSWGvhZ2GyWWeYczMSCtbfmBWwHJt1petn4dL88Hiwubs2UdJpEgC3GA
Yagc5pISpFibsFZ5kv8Mnx7Bed/wmCzT5pA8j5fB3Zyd4o6M9hLkKZ5NY+mP888L
4wjxky+FjghWLpRU2jakNIzZvxdGPVyXG5D9I4iN3TcGk2vUMdJ7j7R6Ah9IenzH
uXi3ulqux/iyJxpIHvEjV+Jm0QoGls2/3uaEQO0J27Qa3i327VENY4DM+GXU2332
ALDGSUaAgE7/wpUL5aH5ESm1OxfqE8cfsM2v534MchCwdXRiLpGAVNH4YFNtJzvA
zDv0DAKoWGrI2kQRHqy+gXvdRtrPeWQ55ZSebxDB30kea4LZ2wqNptWzVsfQPZEK
8zbPzb9cdQBgEafSgJyreVlUBJCdae4mVE+lxWaoU8/0LhT5bAdtiCCqCHm0PldV
rcG8JThLAY9uUFphyA3N71qPad8fPmVz0uAkfOrnf5ANOK4+TWLsNIQWgXE3Qh8C
t057+nS7TeLO4nKloNjPbCgrlpCCB+UH/WOnb4QJrRmBfohe/7bUHqJPj8YUKSfp
zR+fcVJkfp4n5KHDJLqIjS1fsOPwu5nZ+TfbuvL4JAHSTUGZooA9Xx/3BKzq/vi/
On26+UAjxGyYaYSdEyZhoQh+8rwQCEIINXUWuG0Wj7V5OFtpZTixeaaPzcRLnt5M
zCvzZj2cKKbQV95tfQ9/+jWAOcyJ1/iQtad4YN8Yg3a33/Ioo2gjJnfpUdoF3LbJ
vJFVA8I0RIpiB6V1/40nOayYKbbVUX8c0NmYCJVq3Q0G0FGkNRfV0h53c1OoaQmy
9Xez87pzYsMdVpjsKXRjFG7Yapdv4Ogt+IaArPoWumomxBn4UrsHFrHIM8UPdWPM
peO9uKHGssvCa/Im1OhyiAi9j2lcSt98UBSh6AwH7IknpXY+kKvQcde2VmIlPNeZ
YAowwhrsxezsBJyW3oMTndKKvb6SsSW8hPxZrx+6RfFAUcL/s7tFrNZL9tQgtx09
GGURKlhcJ/32GkB5JIcD1LOwu2NjTfee1Ve8qBNsYzv3BvdP1+Q8/jmgxkwIj583
OYf27zJOG/+eillHksHpx3/i/9LAmo1waA5R3uh735W3FMuqhyns4Yhjf0CrD4IF
K1lQP3TZi43+T23xOgqjqEvt30yLW8ZWDZIrmcCz83J4gA+BFxvuIBxw8c5mPxRq
b3nwqbRs0z6fsqP9PbqExyfvXV5NC5X/sxqP6/9dYCR4dNApfeMI/LYi5rwK3IzH
SzU2wVGHKvgv8CnaOY3as9r8CObbA3rLGNC8IzRqKJpUNWOGhNbMJYmaTDsniaU9
Q5RHa0Y79QdkbXVvdeay7BoF2uOkV1lqb7JGzZn/YLiOtfH6Foqxr0zOCiXV5ENr
QffFrEXa3aGWehoGY3aO/GDshuXA5ie7KUmX9Oj1SHZ188O74YU/DY9Drj15Cj5q
BiLEh3ch9EOHjqTGYqs+dPOxd/YiVRjOZ/7vTiHavjUG6dn/SAXgoxCJC/oP+STv
kij7yELelHGV5tjAv9tyrl4qLQ4uKeOjxmXuWBQ+mEa0Sl0HKdph/q4K7ZNkbxV+
6Dmj/pKdrz4y/DMbDfSjk6nrXB3HH8FgwR0BYVB9vyi283R02SpX+PupvhwyjuJB
HdS+e2VE7vAcujpd+pZ6dchRw9wvbx4+L+pYGYeY0jPkLh+qXBY8SyJKEgMBm0eF
qO+i7Hv4bYXjamRHukzKH/v126rg/MGUa2lWyJW8UxG9Les0mJ3UQBI6udGbgG89
ZXCtC8+dtmcyG6KNTQNsnaY3SUom0yvPcMmygRjbijnXvE8wXLJgwvpc64WY/lzh
AmpBzB60B4q18r4/FdBuaxatjRRyaeNLoXzITgbYwrifEI5o4EMTSfNi2fM1rxrc
W85GQ34tLUOM4Ishzs9hFuN6b5sqXHrwBk32p1k/QNAUYZkylyaN/hkJ+wrhZPVi
en4DwwN4PBj10U0JPXPVEFpcHc3Kyx7/8AWf+DGdJOg9dKbVOjfVXeHM5B0jZMc6
yFQyAX2SHl5KWXoidYgiMqypy77+JF0+z4qbPTUuhU0t9aQpqJtlTtyZ3WcODGjM
Xncfsl8nAg1qnjjnb4g9u7R39ANs8VeOT6TKG2soE36OVTACAZgTiNiiQVsOvwER
LKKeshhyH7j/eesNke/b7j+Y7BWjZ27yZLkpMlGep+uJnOsyYuLyF+SmzRI9PTUp
mmiV/zQc9VOoYzyzBWA+2m26oOGmdXxYxBvPiiXvZxduFeNhbQ9POK6ppnifr753
j/SldOcFFOwiKCijNmC1PEd7QPq5lu2K2kC2NUv7F5rGPmIApJUP36k9WGen1fEp
a0xKoerr1UK/T3LyEIi+9XNrT9YCNsrNrCi8OPZUmHZmIfyrOT8INSZSJMV5Ybrb
97iyhLXQDabFcYGu0uYlhj7VzB6QWz14XdjIq2OX4Sp/FCSZYbzS9fAR2lYnW+0t
d3ok7u2ihMbtJmN2T60wrAkIJtoo70kGOzI7sRM/HadsqmURkIlAMrjgmzlVB/9U
mi3r/PvNJfqZlZKNGqYOUMuBVKqb6xRrSg9MCkJ/2dnYP8WkH8YgkmMjs/TfG1ac
E4rQt3NLt+ZuJ0mXUt3fD6f9UJS1gpqc0/9Re1LqsZzmkA3/kEATbWOVl+9U+2nC
s6V7Inn7v0AXq2ewN41Sl6xN/n+Abg3NCgECvPMHmmYGsOMwrEgUaaQCnIhhzQ+q
SAyJNq/LkAQsR6m2lqRPV0Bucea3qEslu58Hcaquf6wCN4DEhn+Z2ADCzHYmd2Ry
JOt17j8DuV0IWzIMMA3Br32JY6WgApe1D0FecdTop5Wo3FWromoVdknqpXlHkLMB
N7CNLMIFGK/D9/6sbTPWWvAZTH18HDDz5yiyKbRA35J+E4SGpj+8skJp4DYcsdZL
TmvlK2iI1tkPN1xyJJpyTu4FhEX8igPy9SJKqGWQWQwrKBD8dbVV6b8Ib8X2s+D9
F5Lds8Ct/o3c4gOTWnIOu5a1QMPOTojfaJjHapsYSSTEfGAHlBG2c/XVuJc1QCkG
zoZ99alPEZJDZzrO2yS9V05AtzAuqGUCUpGcM0rcXG225y7HM/LA8vcD8+6a+dCi
TEAMOiTOcZ9VJuwku8upyDJSiOwQAbpnV7gF9KuzsE+b3C0utINKk2R04h2AohOH
74eluYtwvaLSdC9oj90KrKBOWUEl56ACEUkvda+at/AQzHJBKfWRT14zr08W39X8
d4yf3QNi1MBgzJahxDMX0N8VI1sx/2ZccUM7LGMFPndOHHc3XQBkHNxRpmreFCqf
hKXTUtGH4laOptEexXHm9KPyLZtkwgwtTW24wYINS2iUxIijVBhgXE0ivrQMP2fj
3pTwq0s4Nc4wuEH98d8C80PwVcMQg1K/AvBlcEKDGf7/QScRdGa13UcOkqqDG9n8
bI+347QdwjydHfapy1ESYbWgpv9FbxTU6vg/Ep6STCyNqTkjUepkILx0HfwhKyd+
X6oei47KEeolSq/O+fm+DLXe362y9XDDgTnQoTOryDnShZZDmnSnjX57AyGJGM9b
xfXd3rDtSU+I1rxki901o5ZKDijkEGz9uxoNrLyq04kLcB1eIQr5e1PTAZsDotQu
8BSTdFHLmWjQ2/avG97zpMnNbiTB5WL/0hnZXBkiCEbmjjx7l17aE1aKgeug+Bz/
3uQgYy7dCseBRtyPSINqAzP904dSz+Uv7c1KXW0oobZsg9zHtDNW8xGLlVJE/sYT
Yl8v6WtGNO27S5JWhUGUtv/UbjjcUwCd8MxVDGmIH9Z1dcKEo7BKcjuVAsLFqr29
wjPNXzgB/0pI9Kq4jWqcS7vwDCf9OnurnAhl0EYHV89SI6YEpiJHu1Gc0p3yUjXZ
YYg4R40LqhkDN7shkkiSYdy6Ug8hJ5A0bPoRHY+orlvYCXodmuVmHklau+cD3ufV
AAGdsOTW73+WUiWDuK2LWfStRkNaSCxddFVDVeRsWOKW4LcDtnTTBItn1u/Ojq7e
F/tW7DyrSVtNDACHJuqNwBiucX6BZPm33n/cn6S4cIYcs3gUA1rZRLCvv+pVKOZ3
yEjCG+6FCexze3yyW1NYZ+FIn0+OdkdaEC6J/A6q+b7Ulde1nCYMZMTbpamv2593
BBiYOqEXCYMQAWhXkc5c54kzCJP5IrQbRtFfAo/1oFqU7qtLRnHztZXpNPf7gygt
9j+Ar6UaVb6B4rmpzRUmXz9x8eWTJ3FJpqSva2cMskXXMpv4Q8PV+sUinP2tpjSO
5YBHK9DkUH2TPpUSVagfzXqspj1UEWEafhlhZo39sKZLVTFJLkPxfIp0YRZV5mIL
qMyCnbaAYblb6FfO8fXkPAulilWJS8L9TmtYHW9RjhzrGKLy5sFE3X9ttGKozVid
e68wLPozWpD007ZGdBU3w5olZXritTPo4cOrS/98a2sx9NJCJw4mNAC9Pv8BEIcT
u5OeH30xzsGEGWHKXMnpLsKUDTNffC5EeG39BEv5+HDOXuIoKhjYXdXMgp4dMrSe
77BujHYKk+1o1i1sOQsOAXMj/hlPUJUC63vtENWUScdpPWlkUS+YvhByu6xIK5yf
W2LnmvNs62/n7jakJ7+QOPi+45fuzgPgZxt22z5GZq+foQ0/PZQJkcmpuYMtuHPR
5fbhL5sC9fX6RRFCh/QAyp8IQS6Ub7jlZS2evk9QPZidNPJtJKrNSTadHGE5/iAJ
YOImmopMOxeWhfWabb/P1s6UNM17GtVdIBEMJEZjHKCrpVdgcA/1jRzQI7lKdJD0
FXF0Ak/I1H/etl5GYl26z69OrGYNKh74LNgB5qZXOuCT8e6vF+RVG8T/64Bh1OaN
SKVoFNnzUZLycl5BFDzzKCpqgHps5F5ga8rOLIGFJ6djKf68hp2HTY6yqEF3nYDH
JXbzRIoGT2MbMctLj4eD83vqteY5xkTnNaQrpytgv5kGrUvSEiUsDr6ze0N6wkNU
rumpz7+MjLMhKuyT8PPWubzlos5eh3aXOPyuNOYLvnMCrHzoBUf3GEM2kPbo5LQ9
nxw1NlXOCRTPJw6MaKQ93j82daK4sxQ2qwTsrUSbEWRr52j6PBuJGLiX5R3w9M3R
eJAZu4LVlPlYVSKM+M16Yk32VTy5fUrrC0od0FWaXHehOosEE7uEk4qR47t9f27y
F1OfcQjUnMo+2z1FNBkrWq8goWDbQrGb3os2LFhXPp1JdKr6sNtwK1E1sT+e7IDd
24d9+VHj0bQjRwS1SrhB8kUwdbDahoUxohZyszCYvRn5CfKL/+0FSSodl5eKQOmC
iLUpEL+sMt3u6b9AydPpsZb66BRp8fiK+3S+4i2g+8RgtHFBuk1Ai64g5a7oAy/c
HHzAhRk6Hm/XQMKChuVuj8D5G2eWBKynLtx2/WjmRYlWj8qznaUIAIqPSDJLs06Y
QWTQBYh9mC7WVObEwL7USq1+hWOxf0RyBh4QTlj+J2Ed99gaV92mrj69f+Z3iHmb
H05oJDBPz28iNUCY8Rf+VXOxUemt66tATsypcrq8RT/dUO5Xr1mTqXid+2+PnBMf
7aOX4nReR99QnVQKnEWHtE/1NA6Fp4MIOAZBrVnKM/o9FC0bGmS97qrCR/1riXbE
eXh/qncQTLyHnN7kWymtmvkSMAW94xOmswoZNKQdeYOPQcW7o26EiIrMGtSIkcd3
7KsM3j6Gy6nadikEGqDsw6K2G6piid4eUtecptWHrYkKbEK2rQY0U2NarUHTy3Fg
iiEN5EimNSqbFOaZRMy5aIxZjuPu7/c3qbNc+C18UVLXdW/hCKRmDaAbGcIJ0lIc
ePhQYpOM7We0MuS346Dem7/M4ax7Hh1boTnKeHtedSPRAt5ggX4dUJIFx4rRieBr
wkRodISuQVIYijVOzb2qrpV8YtfOKfQBJpJ5tzjljeqf54QgqgJ5k0cnPXRktWqF
I6aH95SsgMrHU1gCoFyz6eMiKzvjD+638DWO0ATDQJ+Q6QmGkTpQ4aitaazohHYF
a4pfOjB3rvVkHoQ/xVMU0XImmYyAGQZbtK0fxOeq6hWa1VR0jr9FeTrZofIoQOxm
5fmwy5fohb4VJHQ+XmF/smpP9UthrKaZurgBGGSctNvaBgvgigVEO3Wv3dka4EC4
5+flY1sUFk5uok2Ul61vcudsxlDklEZhgoV6FFhFZSdEOHP6jV6VKzE+KDYzPcc+
/05fjxfQKQnij18mUm4c3iRgweTvaOv86cNM7v/Uw01bEj8Bbd4O1kg9n5X/LkDG
AVA4FWwnT0L5fUceudyYMQwbrhRy6HsUB2B/DsRQOVQlKKTuP5/baBMeRPEfkiQg
899eRP/s9siMjs5m/LqLAgK0Z7SukGCAyXTFDpAuuckZKrxQF4i+GPsOQhmyOHk6
AeTCQutLJOSCd5vZJj4MBlnwuEr/PFx6lV9Ep5N6vslCwTxrBXmjslv5H9hy5Ze0
QlM9hbe8ZMFWxFAo6fKcIOhlOm9ZlMl3+WbYDxTLQVY2aIH0lohKncq5ioZYksr7
m8DD4qFywMWxeb3EUwKGIiv67hsRcmhO9ds0w5po6UbJJ/Y+XUcz8aFYgp0yrPV5
YLfHGSmBRw+I2stbbokOyOW7VBjU7G2Ku2aiNToqcPQxNEBzLp2VssjJAcrdwtFE
b9LJfHkTnd3OaigW3QRwCVR3NwWhGWvGdovNuCazcswAiUBvqx4vXTl3bzJLPQwk
RmuUvFtQaIAYBGRPUmIwY7X3rMXXLVXxSgu3pfLxUnz+zr7mZANvY9ZP47FslAc2
r6UccHobvXjFiyti6pHK4c2B9J0rGpQFjBeGavU3frs/RJeI09Ck5P3wyzMtZPuM
bhlgA6iSQp450DpjJtG7kIC8qJNCa6m50V3t+rrOQL3aOb1jVfvxzzeBj7Q47d6Q
jxeEAFJ+B7ue6ra6Gk9tytaJJ+tPgJCb5SxxCvJsp8Yhq2Df1xb2/q/n4wIH8wG2
CR2PNGqX0xb5umWK9jZnxaWjky8p9XVIeU5Sj6C1/5o6Yp8oyGwl7md/7sfuCpe4
1h9q1Rf2OB5bopPLw3/pAu3J877aqdotFsGhSmfYdCjyTR+HWdCMkIVRJU32N1GF
w8H+0mRBHfq6VUAFFuiLpuX0/H0a6r+JdBsSdS5fVZaCyAQIYJKN17MtUiMejYAj
UWinjNmc3WeCvnfk1CSmUyNn8OByjnAMQ82I8OD/gwTw+mOSpj9yFdRJEETvuqJQ
5gUHsEPBJc1My/J/QPJeL4pDFCwB6crIpTTZNznCY+m6/LBcZWdlmiwzNo9OBpII
yQpN00hyC+Pl/dTc2tjietVXpES22gw8gl2tgiIpZPCnbjKyembirtIwMqSO3veh
Q1sFSEvw5+C6n7kjMMNa4hDXY7/5jLeY5IaT6uXbdEGz0YsXzwvbeqo3SoTmFl3h
Q9DRqyj7/y3DM8ZGHVFvupsGWi8WiFbzbn4vicg+xmhkBL3ueqNdVak9Y+oYMOel
JsciuDIALjqvmsNkWOr+L4yzVi3ZDsyyErY6+JgeYGoQQHXKvbdMbyt209SD8CNP
XkgVzJ76NTSkRBB0vIks9WSpf+5z3x8312u0TLLI88fMg9hhIWVw9dFhYcgcVS79
vQtOrmgnm3PhdqcoY0jMmJhqovB+cj/Ty9HDhGXn83+Wqd2i01oxRMQWiIqcWwtq
oCwK23QabHcNs4rwt3Okn4fp2OgF4VXVfbyCzZH3xpcpgG1T6IWRAWsg87KJbY6C
ybL4u7qDoAyebgxI5O7uyOzyMwTBc4VHUTPCnyuxMG0DkafixOKK5ZTP29xqnrHJ
b6N+kU9pnGR9lDzyrQFNDGi01dqoPKzsQqqlkKfHi6Z6sXjEEmFN0E+y9x/kOrAt
2jnAIV2T09mXZ7GbB1/Qov8U05+SCanaK+mg/V6FnyPvI7fNnR1D1pEVsMVdq1v5
LdYWnWTS4rZRbiIQi/2OsaLFuAy2vmeUNk2DaRMfkY8N0Z74XgHx4JTvFKIVbtJj
HsKFLyijy86fo8IQn0iBeDL8zjKPrWm/stEjRuWK1ovJx4IW4Ln3PrO1Jy5ISuHJ
QY0rfmvBM4Txeh2a49zZRTOkFTJ9Ek0FbT/n65omQMAMmqv2ZHl8G4Qlv9QPxy2x
0LlZWln7LFxyoHTIHn0xh13pn56mlXoES3NEsAIsTm3I2n3hRTIM8PSFDW39F3vV
fhfXhC/XbVVXJPEliOOIyu3E96gaugguN2kMHk7rUs33/LnLbYGq4mWPwGoNX065
f/wzJKH39DDwKVkLyXRh6tkATqJFrfy8QL6Yo/MgIoOsWkDX1RZg4AxpuEdJ0Y9D
ytRhREhzxqFt2fk6nTjhUcbjQsYUti6hPsSWCVrMGDMTY02to6yT8KWjKbXI2V5w
4r3FfsmUgkjL+NqZm1Nwv6jZGti/2iuhUAdXUfE+cBB6Nm9mZqouTbKZ/L8iJz5h
8OApT40mcar0PtF680tSb4S4YUHwg0TjyNgsDJZfIVkhZ/tqd/3eWRvULFj1LQ6+
W/dYwltgDjg6jP/f06EUKRllgJTb/KVkBdgz8Shs1qSDeyaY0oeP7/t53T5opd6z
kecR6OuT9eyOwJVJk7rnrpDdIQnHMgs8YMI3NAdWZir8NsitvY+Y191mLs6NYZaq
gtUadOC4VeHDGkQtemGc4I0MqgY5X+6/+Ts/Apwm42jZAgiC96hDWMdWQrLYEuw/
+o0w6G9Zkwob/Ubf26dZerZoNKpZgwkMGoobFwzE637Ysx7fJ0EFy5IaOHMIFiUt
0dPiR2PXiuzeQFbnnRYtaOmFvo2iY6dlqFd3z3p0N2sQf1K5Gwu3xP0e1inlKKzT
wTh763bt2ZrsKRj1ErxdH6OqGinqvgIxFxZnK8a6uahhd6SY0EUJphFXUpVqLL6a
GxwU1yW5rjjNPmE3oCUzMKO2x406B7UzoSWHO0QlKosiIlG51P26nJt5CJmmW1qT
UsPXmiotrnSd6T54r4I0S8rbWUypyzEeYJ+uHmoWV+PzjUfxFgodt3asvsPtKAz/
bFO5h42keRQAjBsJ2LstlesaUogF/I3/kAXAyLWxAl/AwTO1P3hgFumrfeB1uofs
w94SkIfOwjBBFQnO8X94FG6eKgjjj+ghBOJy0XRb1PGmjx8PksjEkuWziXNgpa14
Y9eo54QrYmgrzXEvoB+aftZ+3ezSCVDcjraAmn7PHxN66wtjAfgKJ3Q/a67iAs07
15N7P4dz7NJGof465mmBnSyCbI/HtlB7k6u5TK0H03SzZ8PoZRicAyUymfk7+HNR
0XDUk9KTywXsqUbiHc48o/C5Up2fCk55PnkhZl8i7wKo3OmdtJqfXPJTF72c3pHf
gy7O2G9y+7IOQsUxDFFTc7Jlcb2Q1R29zhIxGDXqXQp0N54ceyCcKYtduf5HwVir
V0LyCTMjE9Hp1As2XUnyxnBVWMlRuIdrauhTD/i0pgaZbeLLuBMSP/xyu6Iiu79U
YYEO3cyrKTI8UE82+K//7ph3fvcGTf7J5h3k81WjSERBr0s3isER/cW+TD+IwzUo
UpgV87C4KDXZbw1/OMmdAoJk+1LTTvxSDYHs43Ka/KzkG997J0AtTO2Qk5T14mbw
U39HYclHK+YS053anBp0QIUpsiWiF3UbVTA4idemwYjJtBkLwfnPI80rZPDJChNQ
0qnLvgYm686loPNTDUE8J6xExhWLAA/vyvHHtGbnjP223zN78/g63v4mvLeURQTn
GdqsPG9dunAjo1F0y2e4vkgMSspEX1miBDYPl06EmlWOQ9bdCjOOv4+IN2h8Ru75
fxum8ez1eR9e/qc0u7gW6ipKywc5BhCDHBbCg3NFJd9AOwPLMTbVanOWkuKOaMam
JXpWKryW1mwDLwruARPs6SoipZgABnm7nWvlEg3FuoYFXhDHITwJXbBhHFfq+N2v
aPOqT7iDXlTPzCtgSNzvEW4LtT8ozNFlyCq1Xs8MhbjHSt9qVr2z9pk5WI87Hj6p
S3Cn+Jg0Q40ohfwR05ZEhgHY6NvWb1PKY0C51kWGG7rQ8k+AxCLeK2tV14baZrB9
uB8ykEoMILZJXBeBNzFoIxcxAfuDCQhup3NczyYONnKEs4OFH4rTlkQlhSUrYAm2
qxLZRd+D+R31VCdBdeycP+ITqf8XoZlHZMZpPuEuVW1BPtcXf+1xQAC0eJhK7ELk
mUnnkJcsYlCyblDl1+NgqQqXoEiR4VO/C95z+o9ZKacQNvrVvOsXx5/wYqBwdyif
Mf2uqrwiA8AcsDV8bhllYLlep0cO6HklAXix/sKjReMF1KIMLqO9KxN9ULAeyGrw
/gSdN/sabvZe/ALz7THnQr6+8R+PcqZeZqhTx0Q+yHwPhw83ERecrYP1YfwEEiss
xDJtgW9HCuy0C0ixNe9yAZCYt1o3oCluPPP4lsgM+fdEeyox22Omgrcew9XFj5Hp
ywbUykq0lto+wQiEycu4jplie7HZQmjHwglCkFWA0rzTh8UJF4GZVFE7UWpuuc0K
iIpC3yuMvahaUCg4vztZ6Xt1aAWUKbJOjze7i/uQBvTIT/Y3CRHxuwOI2PzO1EHY
sw+5IUVh8kflaPOngeAwKhxrGv+hHwkML+SY1jwWO4tWbo3SZsiHMI6gvfQ8sDrS
M/PtqillBnHzruv+De5hMOKv67CFYaXmmfh37zGoGW06yzkyyYmpJKLU8iv6/mIV
UbMYYSUOmy8F1VGsSy3+n0wneSeU/Ynp85QNVZpbvA5ncLj4WC4sZR+qE0KJxUvA
zCfebqCOsuCHe3S7Arkwpzy8m61DvLhFGHfP5zSFlFeFqEwVQ0zeNJkmSf2zcvr2
SYTKhCvIySOrl8C/rRttrpHvBArNZ8gDiair8pTRkjL8rSYhXXFiMwh1l+HHnONg
p4yxvjcxo9bijm95lpy3ovRdfIIt++Lp8E0Fvxo2ELCbzhPTwjhLm41aDzkhS2R/
3lTjzt/YbkKvGj4vMRJA/mWxp95KwOCBZU32/XEQsH5gnX+BIw3HlWSqRAyZpLyD
HHe9g19FZrfCaz5MvQ/0hUZBxEEjjqbVDeR0Y9xghJ7QbRlx0tyeLk3B2ikoXAES
dEnUGzroNg4LhIlptY2+fpcgRySMA274sjRPS6eNC7555GS98IEkQ3jGb9IfwEWB
7E/AXVYDDykW742zJvZu+A2kngT8HX9u1AdQCMavixnf7Je6fh1N2Mf2ahCbKTZ5
S10yaWLN5ZuKyFPMbTUA4avjHVXlTfToUZaa98o+ZeKq0lS35oQckYF9ZFFcwFZs
F/s8W8uvlYrbaAYZ/tawq6r16WVOXxBLfg3xCOZK+kulnBXrfZvIkdwwp6jC4MXb
pBK+nt01fbvUnUv33AELqloxSG+ibBcPjOk/9oYpDQJqvreaz0lRC4qKz1Z+wC7/
BqqlghQ2W7gCny1iR+KqinDZG01ZacxAGnPgo4tdMPCSUjWWWUFAKPXNHCKsOp/u
iSiOY736tXJ4IIJzykTQczJk4jlop+gXTXcLZI06Ls0R4QI2AxXhIamT5JUVDVBo
isb8wiikyhJwHqI1SC67iQzqli5RW/1LPVdCyVITwOLLjGylggOJiDsxiRbmi/mh
D/+DuUD/fByi+ZUeIRfhr9AJe49Xl8tRU56ubHw5fenjMMWDuPZ9yvJZGLZyxdK/
+09feGIUj3k6jfaLp/ohseiuLMtcy+KWkCoCoTv2Vja5rl8KnGIlyOqriQnMdLjc
Jkdxrf1f8cWfmCWpZw7QfDrYMFPKonjp6tsAb2sfkKb3BYg6uAd60hJu7WiOvhNJ
Vdgp5l6aVXlRaKDv4zbA6baeb2uNFlHIjUppGGqPHmp/QRC4PBVIT5e30/wT4Szk
pT5FzJ3XzCVZyzF2pmBS3ojCs9s7hnBV9csPGiB+Ek4a68+GFCtQ35Qo2boQuqd0
iK8K522zdQxXbl8LouUzM//Dj4FCVczy59wOB6eQsUTwcvWrP8T8M3S9uptL68sC
MqMwq1sYV0S/NUvP4qoEhtbvDFkiIMi3POlNJ4Mxj0T1CycNlY4pDG/yweVva1zv
+8KvEJe77n+Gz5LuEqH4YKLqYppqDiOE4WXB15DEU4gMynraZNLnADTD4ITtRTpo
hwxeMLQ7/T5T5OD01hXXdOK1PcV9VAwZJyyOEl0nU+Cx82MOM6SinzyqbRcUrbTl
YWXTSCKNw2bWwAZEUZHx0pkIcZ1BBRGLTpqJq+imlIxDeRLbhX+nqUpvNJgxGOoU
S/9ISEfVJL2hkRgFngmc46lxyBzpQzo3Co8pmVTCN3XfpsVWXAerisMdPFZp9Jg1
wxb+mHND5aBNmTVLAn2byD0yWE8Gv8agJMhP+4H1Ai9gM7TspFSFxo1fZsnkEyKa
mN2uhGLz8A9PbBhaxWvYUqkhrhEkwWeT9dL8wenR8L5FoIdJCGxNv2OTYlNlJqng
uSqf0r6ouQjeTOBeHk8Om5UbgjuikVMO8KHj+vUvS+/LwQJkg6HMQh7xX0FXgoLD
mUsVwbJrRoT0pW79nJzdkgQPgx/ctfbsV6tSar5RigbNq/d9nGDN8V4oEzAfetEh
9Bns/VBrnLYABoHjLHqeY4f9c8oBznpWAdir6CnCZK3UrMOsHS5IpApHhZ7VaMq5
KQw+blBIZPV+cTpp+Aj36gOMnKTYuQ9V6x4DeghN6Nioc4JWssjt32WQc5DDwtV6
ygIJzkgMZNYkemtEV4NkXmQ/WvXRNwTYxRx05GhH9be8V2MHBd2gMzizFMgAAfsY
cc6eBoWlL6zlO2YfRbaSwqfpVArArvPGFUqVyJCWSxtPQm7lpsG6R14OOZghfTUH
aqO4j3Xiu3zl3OG+Hr1BYdZsCpa8CanwTtJXXATeI8AGFT9Ka3dY4zNlv7iWnfUD
TKqWBaR87//FyXB6oNJ02Jalpe7QXjQryheTFFwUgd21gL2BBmmJf5AW0BgP/xT5
XeEVmoK3G6WpVYbj7yHwas2V8oPdO0/N82H5VkS51Lc1dtcHbvcOlfvJ3z+5ibwv
/qEd5pkpCLyKh1o7kE7bpj0JVDKgygDlveZpsg5VYmY/YC7DUssGWEOGleatpi+A
0/yRtD09gHXWFrnMSc77FwSk8Q4KdeDXMjqfgU+3l0GJxLW9jMcVH1Ky97vckMCR
mm10iVnVpHieILXQwuQJr57Hh8ch3FZ7Yj48a1jhrszxigDbH2fvOTGbnuc8R2/y
Ud7blhhEZGpQcsRHNMYhO5c5RcOv1+X06zlmwYuX1Ru0nOCCttZVbC3TkWeEuxrT
seElODg2gyiCbFWQWNptyVFnCyUDjUalKdTm3A5va7wJMTYS5+bfAHCu48uG+cxi
XPExtyZmzBkJYfjq36aZ1M8BPgfaXJ/4ZH6MaX7h7SJZpDQdf8lWorHL8AniiEh0
jBqOVcH/XjNIIREQrfOAnVzWMZVCHVAKJQ15JNgxmVfPhEg8s1zubKg1kVv4gQke
rqQYhuCcjHQZNoIHyYFHQI2R/g0mPjvYTR9aQMgii2WE1Mq/GkJXK8DFgtjExEMX
3D7J9dn1aXHw/7rMrXxjT5A87Tc1H8414uRvJ6y6TPcfC3P43jvVIzUzRe4Y1XlB
OWkk9TT8HFiAlRHozyULnIx8r7TkPqpUXlQuvuZlP+R/h5RDeT4tCCgrI9PEj4bf
Qao+tjn40DLxzVTKEOV5VlGNEpQMBO0Gv4g6FijItUYtPKbkyMdGec8JXmeEzuV9
qtqekuWZcSF/eBZFq813sEuKgZRDcOYyU3j7yuPeyGTlYMYY6cflMbopsfdwRLnr
xmYXE7qUtl23SQzjYMhupL72MpmhLwfwZhhHuOfgpppTRX8rrZChvzP1wjMPkYzD
A0BSQc/E7My6fHC2vrvE+AT1zRtQX1u3yzx8KErr/abW3GJDeUDQNNLA12sUKWIn
JLIUcFNdeKoC6iQm+ym7tDhjnUOMZg0jWRcxhoUzqK83xYnNoM9vJNxxp2o+iIeU
4T79IGstGd0UX2dOC2BAM8b+/dbYhv/XQB3VgXWRinWJypgFqOazoTiReJC1e5K4
Fw33aUU6aP/NUZB1Oh0eTAZ+utvgV1wQ2LLq+QytzVwJFf+TFmWIzBQxt0wLzRTL
Tld3E08ZzfurM0Dl1KsVzHrFYOI4mBf530BcOEbJvtHWhztBFnJ5Si7AzWzKSxal
DXEAQTRpLkURCr3X/NAqSONdOghMdP9SMSVt2Xm8mfpH1pyzi3JznnD1Ba66UiRb
Jaio7xKAooSIzzpfQKHAVMEGGYRKOM6r5tTSlrnXqeYPAxw0qo9VdUh2Ek9XywOb
b+3EwAS+2PofhEO3jhLr58XgBwvYY3G/eVGGWUvZW65hMVo1o6tiACyh5L4+nSre
dLe31vrcD3rkIkaSGr+9aTUxiDF+ZpBJJ1mPU2iH7g3khljfz4GEG7uLsrHn1AJD
PLbVl7Xy4SHUwrF8T0IRNB4BOYcb8TkhKJP32i73RDReKbQFScklv3FWgDMwmisI
hqZM+GlLPGlTRSSCBkOMTPUE8msHK7+8RRTFscCx6vYvVOLdxzFM4Cg3Z1XMkmri
SikJ9JxqfzA0ofbysEdKBnxq5KSG2kdKq1bHxbsBjtKV+xdLTEfKhQEwPrglbwZl
0RTsntEVKGmSVzwcyWvTX0CdAlo7y/3+seqfAYPdG2t08F1TjnslPXMYkubxq9YJ
dezlufoDb6LWDaaJ9Ey8rp/BvGcLordSO7u5ZTutvzbf3/yAwPn0iSYPq+SxGEai
quD39t3vUsGTLTaAHuh/5EGnuEBDGYjear0ShGKX+5JIBLPuL7+2dHjv0N/5G3mj
tW7my1LwBeaO7EocfVXh0TbTe4IWcEMmELYo5ospt3fjy06mQnFNTnOHPJqiUEUw
WYUdbolkoO99+XA5ov9ubWkb0+70cKTT72i/iso1dJ1KBczpviEy5ZGPcBteuI0y
JjEsKIDeVlpyDhV+qEhokbGqoMxEsETZRGElAR9bn2jGq+oB7Jy0iAEwXTMUYLby
L7+U/0gWDRes2VdUNUB16j8z6IBcQVfdOGOgq8I7/+tEDwT5SKwyIWpFiiMMcvmq
303vWb5UjqeQypq8EH0o9uhEpBpv/F5HdvGBF0Jrvd/JgYtzKnvHWWeqdqxUoj8X
nUvGrk1PfIz5m4tGDjNn2nl7cupWxnVDV8RJFNNA0tT2kCMMu3GTwQyDfNNPpQjO
iwwIkU8bJ51FSXwdYfjMvnteT6IZyb/BMvsm5cpngz+iDihtX4rWX4QfmSQA/vuo
rBSvZb4lVaqGtjlBzkMkhf2ZME1DPDXJVtfrMCviLkZf10sEHCZf6FgLnxnU4pC/
0qqqkcJlDDHKCW8iJKVuqr2/ivRPP5MeVgnUcBEuSwj/bllQbBg3YvJnLc+fNypv
NSUtppZWXmbiKyUqGjMoWa5mCWQWQ2+3ylODyf+YpFYmmuDtGBr4J+n+AcYMUNUZ
+kZQaqUsZuUbu6gUAXOEGgRh53qOgGgAaUmo7jlv2eOKWfu77url+x/1u4Dh2XEe
9RhSFPkFeNaRhzqZTz2frvhAaaAi0b347onBo5T02nfwEDa3SQkwbU6xxlf2+2Vr
dRpOQpgDQpYdp8lMRlw8B2wkJmUj1LRRnHzSUZrHGYyA0aVFeDsEb9IfIh73zaT4
UpfDPOjPXKfMOa/Fc34RYTgZSIwRw7QVtmBPThs2uAauJBEt2jqhE5gMDZV8SbkK
Apb+rXgS83dBLJ9jQRrCAm5SstwhmSwqezgwwuhcaVgHgFfstqlQLw2PFFAtgRDO
TwlEFl6xGdlQgkfz7uyYRAu/yPiRwpIQz6v9FyMXVGZIhua2nqZpiWtkoc4q8MPT
pmv8mQWlEFEofQXD2TnrvAqDqad9mVOvum+1g750mKCK/yWphv9Hg0YqVB9FsnUk
dGWDIxALns9jVY+VX6ZSEwfbm4cHvdxwzZowA4iCj2FhfYuZjjFHlgEQ5hVpsvwS
zJvrs7qCLl/sP66OxEigeyKZLETCRfTna47sU97Ne+TwTIN6tA8no4YR+djyyQmo
hVwjN/2yP3yl8WsRdzFj1GyyD4jFTg1n4Ngs0UOOjTe97ccKml0DpwIVwpY/tmci
0jRi3Sd73nOJxZVJnTDm3pqEEpP/b2mtlUvDjDwjH77oho5WpFwiGNteTlAY/mlI
HUZtkj8JiDVbszQP1Slbl8jwJQ2Yc7u//enh+YhaUgjijjoYfkA6XUOMQ0uCeP9u
jCGP4+eOqJIphm6RGXCU0SfouPMj7qqWWfubkEpsysJUEi9QcJlwPu6r4cca3W+B
xYGHmM/RF4wZgrXHyfkCqR9GtCqve5aomwKu+1ofb1JxZi0xKeCYpO47bioDbkvd
kjDo/dcPRgeDGS1/zPuCbwznKon+aYBpEUeWuSJaGMfD4U4gffJqe86JwskQd/zz
F4MrjmiLHEKtmEWZuSk0jlT0j51Xh1RXeHS3GQg55swrVBilKj+lhIFeNWd5wTOK
4uOtmn96k+zMOk0+i6qAMv0FwsXJrvaIcmiQ796r49gH1FRZnJJM+T4Ff7fnLs3s
NdL15h4/lFMdwx/h/W2IA4OEeGpKR8yNvo9RT3E9DpE3emyHcjFSg1wDIG1gzi1/
jAk95awsCNqN/E+4FjPOi3eD3Cp17VkNWUAjoBXrFhpOjoR9vunPR1kF2jgT10Ph
BxoPc7T3V2j6KdZ+01DI1rBEU0RN/KqklhaC9+laqWhU1kUsCT/5VeIK0FPxOOmo
VFsICXTGmkCc1MTEdvibtIQJHEprn+1xruHn51HIM+r2oxtqfkg3LA2huTIDAdey
TiBbFyEH3CKoEs/RTATO93qBv8wIR5/VKyTXb0ivAaXoKytM1WU3CQu+1hPfT7S8
thx9rBxgvxmFZwRLgPnwGVEA6ijZIBpvePsys6yzeacDg4IpO1RKULgagfJyOcbv
teu7S8JGxV1fuWIlWfDvCmyaqq8jG2IlWqOEb/UcrhqQte0K5WsI1NEbCV5PlFtC
74ZajZq36cY5ntzC4bW3zO9N4gpPa7sSXh38p/a4uHaWf+mILGZNPg0foee/T+89
SSkfy6qE9NEo1bztdcSLCEnFjmloaLMGUQNw1sDX0dctxoY9h+jaPEeXL27HL4TX
iKulJRRfPskT3A8h4EUtcqlqv17maOVOMIak9nrqG3mytQDHEp/z5mj7R0TbV43x
F1qusuI54svbkIKACwM/SBNcbiFzUo/zM2fkDE7tANCuJI+XbLt0ST8ji0S4XcyT
z+/3/GOpp5ZPZgMk0CFtb7m2pyVTfYV9MeDJ+2pCpY8XT/9qdraH2WqZl4c7yD5w
MVkZ3Uidp9KwbXeQzhxMiM/HVLFwPBL6pCQdzn4xRvMSAxZBfRuiToQla78Nwkd+
iY2NMoAV90mb98l+eNzAkAHcK1abBUPMdk8oprMCyzVFeBun+BBT0HNeNGTcvjbd
M249xuZvlg7d0LAbnMZ20fpEwZTRLCaqMU/YnT3214e90eSzWa/rmzAZS61vpZmI
ZuoUixb9mGm7jGgbTbuz+W62CaBuYfgdBaVuPGxIeHNYKX2d5j63Dh4W98Xsir07
HWmBNPAHm8juhmATzimrtICaWxyvBAH1kF5RWaR6TbLPFMxtKtsVfStKkQaJ6b8K
JDspcxUkXaHdriCdtVHbJtH5yYg+ikqixeuvyEwH/2ninJl15INjqZklrXPocitZ
EE3npBlLvnnG3WBN/KJmrCvlfwpVFYDo/X/6Ikdj0qDW4dR1kDeKXSyPg3239No7
d4r44T1YnK6wTULxBFKIERizOLrowM67BzpNP1hNCPsCNCUK3TmkHc9EdFTqy8oy
gcEfMseJ9h26jkmsb4hS4WRAbmvG1WcZLssa//ODjssoHiaKSn+wd3CUylN8EiDH
vnMwquWtlHSQWZmOXDC+A4qux+j4+P6ZK1bgoAFH3QgpQ6lAsDctwxTXQX5rWoaS
NUamTLjZvgvADg4ZQJ5G9oyWWjAsLqB5DQsJBh4BJg2jnW/sWp9T/0S8LkKEvrYp
dgZ44FBbber9P0pgBSPP84YIlSE/4fYQsmZdPnVG5RwPsxdza1Bgzzhjj+NoX3q5
69oWf8khXO38+IXeRxkLLuFzuz8/uwLfDbvYdQUhPY+Iy078FRDfQSbK3LAk2i44
TBeWN20AR2evAk7jXJt4+jPoInmNztQNLnRSLn1x48gbg0jRdMgbyuhqBJTMtjoX
mQZOHn1O56op9Kk7+9R3xElka844je88L8TzRM6vRsJPSnFlE2hBtlDH5d4Q0Frj
48HJVRRuMU/dT+baZVFL8p9rq6vmiJLlmGVxVDj1wHjknihkNXXxzhqcm6RiuRbp
6YpCuLdtGkvtBMAtzFbpT0Dz0XdObRwhaSI/fU9KpuyM0mROcIRPNySFToz8ewHz
WKy2R+BaQhyYqfSfXg15vC6R/LnzGf9T6LV/aZC0Z9z9aFo02qhw5gNeLZJDyeKu
xSP2re/KENQE2uW9ErV1BR+3UZ3ZrEFBf0lgaTGJMhkRjQCOSqOCMBZognQZLdze
cwXyeEb8+bNg9N136Q22BXVlQ+Ype/Mae3VM2X1MiQRiJBp7rf86pbOyvG95loTk
BZTsfGjbgU6SWyT9GdgpAYj7kTNoW8zw5oj/s2pHjgju1dEBoY5VebCpf+XOUamc
Ld0K4NxRiRlLn5hNw9GSqDHlTQllBvwbTRoFMk4Xgoz55ZYfV3cy9FKAb4QYa8Oa
DjGH7jPnbILBu4WYb/USSkznZB2Oe8xNFebXMGSwgw6cG5HsTqNY8Yrdz+G7Oxhs
XPlJebfQPZWXFgnI+vtTMwxVpWhwXT9erGtBQNE/PwoAMFxn9pT2onF2+qTXDb6G
Vj6iIxZm8k9LwHN3NgKvwHXHcJVNrd8HMfPl/+P7vYrI/V4R7i5I1hc92i/71qpf
QdTfkIXs9t9904pFeaevHrZIEMP5qBVXHLfmz/KEOLps3nVZ0PwYCsn9yJd17PU3
lmZi+P20e5BmI2c9QQ0vw97wHv+cJKn5ChC8DznNqruLDXfz6heuI+rxe33y/hnE
LLm3BroYtNDKKyiK/hLmGvOTWFlptbaIQcAHxv6cT+4gLsY038qbkVG/+cCfIucE
hVDASJKv29Gf4aEBA8BltCf51vOzL+yB0dWQ3sqMb07bdtw6d/SIA3IXL1zrkXXE
ohQ7COIsx7JZF6ZZUPqufImmnG/cVsHx5fHcuoUZq6Rns0qRgr7w86I86R8HbxZH
+aEMeiRzUYe7QoyBSPFA3TEDRnK/oFkSIm41vpOmEetO0PUniewQ9TWHprWCuqxJ
bzdrMcfBGI1kdvbgyTgdNplPcLZvnsaciVZ3fknWDIAnH7UGQW/tcWIWqpzC5hT9
9mDVN8+bsHpNqqCL1cx8FPbWtXPsZpc6e7Z8p7U9OAzeKnCn+fbwmWdZrNisyQRS
sUv4Bp5Zcsr4lJ1vF/K3+l76y9Vlnem232RCddb9YX69bj0ALSBGEin3sLnb4IoD
7Kq1YxLKii4cQMqSI5HlF6QvwpmiXm9hoJ7oK2KVFvPlNMKZIbZ5XI4VViinCili
lDJdSlG29ZLgTve3zIe0+nLcmmX7yxJTm3ErF6ES4jSDiq8WZMoD6jDaRqzzg0wo
z5INOzeXyvCbBAQWTlxq1haTsQMSz+xoj4DJhu5YkdnTB64pznC60sSFTzDnTKzv
Jf+82tj9rajZAS1OVeNsm9uQwiQGyvHaIzPtzTRdY5h2pCzxEzmCAJ64mDoCOxaG
ILJdW/PzaiIRvb6S8iAXPUDlpcdmTnzhYJgNTBfQxA1MHTluD+8nrNNruhsHwter
Dip9CVKucML1Q37qUIErgzPLblOxElZZNoz0s+nnbIouXrOAFV5rZA1mr5igjFmT
ZF/A6rSi+AvcmNDJ3mpF3Hu+RkbQrQBk7JXAEYdu1U4kh+KFYwulX5SW1PJbhtmt
Y5UP2W6z5QXu3mXhT1arrKMuDtlKT5V2Rh0DaFjU+9LzpF3BM5YjuonYTD7VSEfT
yNu0tOLo/DnofHPbiQcIF40fc9R7yW/Xtk+NsOLrh4yJNsxwvyg1MaRglInM+qrC
X8HxcDBXYYaOwbLIZpMN5Smvm8bnw4QMI8N1kpCzCtT7b90Ia+E5B7GnVd5xansE
T1hd1PWcH1MC38glDibHF89nv5HTERw9ND0fO2STD6ZJvzFcR4leICDfZRdJr+QO
2iwZDqC9Vk/2c+Tbk4RLustCVAPG5+C/NiKc8RJvQsrpShWimwv41ETREcZ3Ikg0
I/kExBSdWIrGfnkkZMR+vEcUoXwqEBIeSALhO7QWKaGXOw57BO1Rsqeq/qXhiCsX
/stzGdfzMJfe0mUZblXPJNIt6phS1Obz+N0XGwwbA0++yAQZc8fHW5eADbpgK/dW
joKpw25j26tkYclGEz4Rm2DXHtRLaXqh2j86mr8Vk98NSWSbaOQwesvdQYDv7SWM
DPwmsX1MVgkljtlpSiWYCooLWX3TcZHldHBcT3WVueSb+qka1gJtO4coExz94SDu
m78WTy3twapctXY3+e9p2HwTXuJC6r9X4oz7uSR63mqZQ738l73wT75NbZqKSrxe
Rv0I0jonDBFEyhnOoJ/JztnnvBtn6+MXuUGpDneRGnQXI6/oKNspUCbmgklsX50L
w6d4zxPygP9ov0uAvFccx3Pl/o3LU5Or+lRuICBgcqpFhU2k85sA2IMzfwgOU7zt
l1vRpXXZry0zy1fIlpPz+RHDoWx3gJ5kuvuklJezX/qnSBFjZpU4aMI7fKpUgUTM
oykk1NKjqlOfBbHRZvoVEzEYJqbPeme4s6XZl4p/7XCxY4wBbG5FdYPaBpBT/qV7
YUbR2mM4OUdvg8MJ/M2x6Kcq4kqIZGKghduJ5iVYbdnSokAUuDOUZI8HOgiokXCS
qZJ8YkG3IW1wspog/vAMz8pNltJxbAojplQcwlsjzp1mdeqwcEgtzHrteM21751O
ZLea3yqyV9IsBBMMpvbfWkwjY0Xvz7f0ib4o2ot12xQ4JQ7jZ+gflAjE6a7rK2XA
bSukUBFacGYMcCjjgf4zlq6mU0t+Fpybu3IRl/uD/GqttKt4MBUYh6pPJmfmSrkY
I4DLqVGiF7bCqeD2/3OxHQfuZ/Q7LkT9atyVyHrG7iJk5KXAvhEjDeRMDRTjh6U5
TIc8w6bVc4nU7UzbYsHH9rTKdGeG7Uf+26ETz+OSQqwE2GC3qU1yLcj8ev9/6J9+
Z8Vz14a+yYrNG8JBny82npALh/rqdGnjKmJpswdxDD/Xq9th4sbtBhRBaJIZnAxe
Jab8t4t3L1IyyyyZ1Cu+q62FuLNuOsyBhvo4z5pUuAmrYthe4yLm4hZXMo6nJAj3
IgvqpyuwwpgrW6JCvfC3Wr/gvp+G+HjcRlCHrdug9gNUgMz+XMSKI4o1ZB2mHkK1
EK/PnjYbMHnAjmvwJoiOrikXVJfgeUPNPUSoDO4Q95bLfxQWjzPq8rePp32w7uf7
0kPofuKA0pfFk4x4rIhCPnXQOXUe7TxfUfQIpcJLJNF3QhRP/LybTtQ7S+/T4lA5
4OWbaYw5MsSPXKq0+U30+uigTVT3LjcxEjgrMLz7RFzbsvzZ1AMTjohrCHu30aBj
pMlB5K+I7RlZVsU8BGqntnXLRmgljl91uk26xRC/tvs3pSyZAagtzA3r+FYK6oIa
skEqkKDlZUcDobsU8dWlM/jr8UyVxHt3AVQR4RfdQKMfX4ifcFkp71DNQewb4zzz
pI+RUkHjnNubspVvQ1jtFmBAa6teoy8LRZ9nXtnf9EIzsBdODQJuEtH7qkIJzcpY
x5lkTJ834RDlnXIZopZSGeS7ytdl2F0VTVKmkBPAKF4jNE0/fEXDyj2DQ0wG9w+z
9pl8qQT33klHyrONUew+J0zlEuexQWEK+CZnRtya9+idPAzkfSm3w1YFWkpUuTDp
RlKeEez5T1ccr1rKGrvLGwsa7bFmMq4xZ5ujKRTqYfqeM1uaqC4gMNfhKZyXiVxR
7ss36QHWl/TleJ8CD8g5iaYo/beT56mik7gcIGkSPW0rc2GFBK8LVwCDGOhG832T
72bjoFmIib0PjCqaehSVhsaCRjMy4HiVSgc+Vop3wNho4rLSyx/LW2yz1dwLdkow
tCuLhS2mQnT4NjImJYZruvAwH/A2EkrPR2gRAQ2chs1L+HL/ER2z4wOJOopPiznH
Wwrehc3tATFX+DU6XnmxEE7DfYRK1P2ysSFv8gfgtk2UIjkItCD7/6t5lB+SkipX
xbMuw6ht2rGK2bM66xHy8tnQphotm0FMx1IBSIrND4Dykbm8YsoVJbDFUZ+PDxOk
Jw1n/ME02lci1htbiDVZOKx+nUT4Cp+LROdto+E5IXf2yPwEsJpBbymSLM2+KDwD
y1IiloqVXNetd9BpAKt/bCEeYdSMvnLYn6nw+odYvlWc05h7QG77MLDs1H+LJaCy
KNiUrnPisR9Q3z5TbCn1kC80c6udIOx52b9D5c6ff/2FC5MS5fmcM8jZ7re1NV+k
X+e2PMcM6jT7/w9jHQxehZRJhsPCZRxj08F1sCSTECJ6dLirC4CSwGN2Ty5bepyw
oJlwQSjqcoKpBZz0CmWmmqAv64TitDl0pZ3JvbV1djp0dYMW0DkxioLjDO17Bjfz
kuOpC8WS4Sa3I92X47BLhwQL8NsbTc1E73V6diPSqxikcmYBEs//fq2SbkEwvNJI
l42fiSxr7qBGLqYoB+qYHbq4wjeisYZr8YfGN51teoYeImxHn7fxddrNkdhpxOyg
5xE4nlgtqgGOvxMGN/NcEZ3bwPHKSkWRkeTCPJt/jtwHD/TXwTYurXn1QdUYdOPc
Ym5rOZRXz/9LK8wz35R6OpP2u4y04/tNFUUb/RxStlQxwgkYgs3990c/xmwHZJY0
IDz8cUjC2+Jqj13IMR0rESH8bc3egqFaPZyXl+34c0OYk/wvPAuoXLlJ8CyU2BXP
DSVDYOeEUZ+fS+4HwE5OMnbwiehTkZtUFh9GHM5Cl8YLB4L1GLdJNn7bNKbIwahE
luuSw9MGMpw0QZBltqvprlqtCxGrHYOPKy8gjIvMK3xxgMFUXJziSM/6vHHUcTN7
LOn92xLCaN10+LGNi0qO4K2q5aPAxFqFsv5/i6MN0tikAx5aaP86SjMKhsgk37MJ
Txyz6hE7FHes69/abfgQyUkijY4pg7KfXxjYq78n5VTaOI8OZjdsV1I+VT4iCiWm
HtMYS6MiHFb9wr80AZqDDDIRL9IjRcD+uQTtLLNYfLQlhuKsi26iVMjiFMsa2vdJ
5ugyDeC4ffpcWGejBUH0WuMQQ4D5lOlZdempJyjiSvw+ANAj847VGmGHK9rHChbJ
HbANNlJQTgbGN4NujoWfHGRT04oHtIm2ogCYssZ997fCqsLqT2sk7bvl9y8Es1Ld
A04VtfB6wnNb5YsOu54pMF/zKXIkWT4N0DGW0Yx6Ge/VPX3Dz5H2UbuN6I0viafD
MzPgzGAL/+4MQe8cVQIHaAxiAi/CUZu7Etj//M1C3pXZbg4QHpdBTq7iUPIME2/n
zPbyUApQKyuuzLcCcAtj8497uJXfvcTJLw7iJgRxtZWagXFs685Ou+isdewViCkv
3hlqqF85S4bBgRWaGBpwtIJv447QDkr88z6DgGSjXeA+9+zUdh3tuq0r4GVsRZNl
WIKaUbByIzvdAegyfFYFpxFHRAmTWshe5BfNh4Sg9OnoJrin8wAauS2fqa9qUda8
Ez5lO5jf5eqeccD+Darzg3WD6vG0brfEK3QnFcJ5YqJmNYh9ef5mTZyyL4NIZWeV
4qilo2Qp8LO16zAIozxsmxw1ec9wdt0dFc21lblCRV29ZxN631l1KXljLpUJ7c4d
nYiVAVOo8qezQhz4c48cWcEvf2trs7Et845e50KF1sC2XXYUObNRhLDqiYo876Fw
dKPmtpo1OriicpI9mzhpeOUPe9UctzpXitF/+0PtFuVYFiJR1Y6MDd4Hui0dGcN/
5yWBucrfI+BQ/MPtA7IQOIapHEy5JqGiT8y6YBIJVBI6bOcoaqLOJxKeI1TqjOHC
0KnUwXDF8gYT6bpn6y1lAaf/qjySo0fwn1h6VjvbL1DWlwbY7TfqbrC8GVziJgsU
UzwO6wrG8ZbJQQFhaLEk2VQZpUAWeNOmPcEHCKal8CV6wyOB3/7Lm0fW9/i/BHGV
uL2isOd+QqfCQBPTzOdZimw41RQYgT1ApApsJjT2jSsUrbcWY0WwCa4r53aBOvE0
TzmCq8/Fa2GLiU2UPGDJluaAVgoF4mTvNFA50k8g4tfUZ+QnP7jaXp8jpw1mUvNd
xg4VdsxFHNyUyTqKDfosJbNlOtBPkjvLozg/vFdAh6If3S0AbCMhLMk1uMT2Aj/T
86FryRYnTDSpwj+PlpObaU0gFYG3NAfj6Cjg97S7Ig5KI/3PUWPjJXb2JvKtuE5S
eFb5bj+P4OchfdozJWsYajhl0vT1kE9IQAMIcwSkiTJifOWumFzA3BvAcDzZ0AJE
XYj2bj2677E0bjkt1TL+n0OqAaPPil6DIISxg4UCBIgFHVil1HVYxagIYBxV9sXb
cY4gXE/TZRNEjNlkifJLXcoH/XYzXL+VMaYBecvTgeAc7Uv3tdTb8onFwVnHBC72
AltFpHAtskWNc1kaAezXgrhpjlHDfTgMAPRcHhi1I3S8EH+OnV2Z4ScCTZWcasRf
+KpmWjkNMEme4ixSSBgu+I16jd4q3OYTKHExUI1QwdL8wnFxr2wXR2UGM50lQHwU
Ma8UE2gLbTRH8GjIU7Co8vj6URpXJOjW1KJ2jLBS7iSrXZqXIx5Ncps6NMaDboKC
PptddStf/7NOltX1BtTCtM603jKkFkgHBMn0nY3++26yTlnZ9LXnTJtwohjDR07n
KgaDyzpchilCJ94LsH+BVeVw2lugUrvqRWaCNZR0fK6KB5U50TEL+Kwfrjk/HZc/
eFk2aFIgHl6PSh1PhO19QfxYqC/Y7OthCFAcb22my/W8jsRtvmSiiCKV/pHzCQ28
dZAzMm0qC08ykjQBoOWLybT7asEjzP9/f7al0NRQq/EkXrblinyhy9/F7G0JtSso
yqHLKeuYxoofWRVq773S3+5OcNOXdMnHJvPvPSMcWY8q8tXrb2gtBp9QTQVvR47p
s9cu30pZLyUOR6tLQCWfD5ptynuiL/gLQdLC7hFvpwY82ceyYWzq+TUUwdHgrsCb
LqK3ZI4fnwCK8KiewiF6z0Kg/7tPon7F7OkzekjxBdIRq1NyK1lSP9lVU+P/fJfH
lSKsISencHZ1hetc7SIszMcofSbZu8o5OOHaEGZ0W9blOVap/VPqNpuv/y9I18Ea
hNsAPkmw7yo4CbEWPID+cWU93VMYRa/pgt8oiWEGJaGzLKPrLYkzeb76KIzcdi4y
ZyI0GvuTi3SQ3HHkxz3NzyisHKqPK3nUEfVZIHjRaYFyaQe5TR/d5a/k8dj12fhK
O2axcvk4nEc3KPYB7s39MbKOwQ5loJQEcKeHPYxuvJXvrXhVCQ1cO9j7hq+TC5UE
CeR5XKbEEVETZGBAhCytnf8oGwTmSYoCYborDsUCgUvGsgkj3hRPnDapusFQP1t3
Z1CqS9R7SL8zBC5fg1BRq+lMkZ5ntACoBw610vsAhQsCztG5bJ9FUIIupHmMEfYT
3Ex+TGVZBGg1nLhAykx5zfxnSQ7U+ziF5LjTg8B8neSWVBDeqdl2aNVSwmK//Xh0
ckxcBPtmuAbyCnPRnA5G93ZWQANdUQMXHXEmlLDpGMpbC6t9ex0IizQLVZyyIz46
IdwuzlmTycVlTR5NrmFeedw84/1jQ2TLz/qUpKwgNliSx8DJ6l1xJVJhgA5ZjcMs
YR/Z7ejjFWT4jlvzr11NUoGeUefJSJi313K2mFnoGoq6Ck5oV7RAvDpTlZPHkuML
Aa6zzR9Y9l5aORDt8oHU5BTf4QO0yf5Ol4NHPHuN07G9ZdHU5QqqiyMgLaC6RY/c
nRy7orHWEvJwfmwHrn7pFK91szPY2WBQt0OVSR1oQdwj+pWhvJk7j675Bf/x805h
GA3KcIEb3cMcEfVSKMAn7SV9w5Tb3CH/gfkhqYD34PE6X/kXhnOtAN4FA+KDArdw
JeYb2aOLpm+rT3WeloCTc7Uxj6QuQP6nDbl01h0tLCVgriw03oVsrWh7wOBZJbwY
qaSb9J9t7R0rTrDubUqkjwju9Dr5SEcov2oZ1TJLdGbwl10T5TqpC/9tk71KDnqs
I33LRTFLSRC319fZ1js7l2tSekvmCvAsL+ldAOiOp1PB+s7NyFy53gfJgZKo3Tjg
U2c7cgFIbojn4v7Oa8exHQ9dYDjeOAlYzHnXwtw3SRIscd17oXayPh9qwS/wk7lS
feRa+ZBRyhYMMJ1uFkz3Iwi3Q7XTwtG75RzRvZCY+n4JXK2WWvszh+jJpwpki5Zu
ZNkainmYLOyZhGTtKApOBlA8s9XtAjAnmAevwHGD+B+1rNFMNBEQpEOVdW1WvXGr
Z+K1NI4nMbCSP5CIr3TJf3jtDfhqAWppNNp/SEqTDaRxZLvwC+D1zs4XCGWRfc5n
fAN6kCPvYwiE/93i/Dcu9zNNpU2yo7ZSUDPxpCZ2QRh065fr8hoLBgHiEABeRp/n
TT8VSiUItP+srHR6Z0DAnwxh5RxYGWTRpcHkH80ofctf7GsFN/DS66vm1m/6nQaZ
fLaLDg3ArFIH+sJaEu+rcznjaeXzW6m6HghlcoG/F9zcBlF+9fXmc265sCziyy+z
oOXgr8rm2fImbG+T4XkfZfj1lj6Lvqi5BgiRVemkoXTqlvRdS50ohkr0jj5kmHEv
HPEuPuC5jIE2ZiQD3waNTFYY5MQQ0R3bX7pWCKYnJrw/FCQ5hhJvX36J5vD00xPf
a8pU8RVFysyDELYUTs/I9ArF4vPPOz9sZYKNRKscDsN+D2aXaFbrysem1WMm++C+
ZsXK9dzbtwjagIHG1VDvtSFxwEHw+KRmENFLFza0WDSaOK9UVtpepvk4+bJsYLgN
XKt97u6WU1lCLgNDemol/KS+1pWdL6tEQD1FR+k75OtUk43MZ8quNTWQxbJh8NfY
3Y9geUjU9oIxPg8/3T4uFlEjVI28S5eYq8H8yio3sAAoNO1CKz39wU3yHjRw/OU3
0c2PR9vuk3uBxbuQoNwBE1fV8on7CDlQETmwNY9o2suqnb0X7KMXGzFdrbuH07vS
XtMdaCb4tNW+IDVzMz2U5t7gtUFRCO7GZ5cg4a88h/lU6AkVmbvh3mTjlbpypNM4
sTx8XrFJG87wECU23JKYTPvcfclBcqvgo2TTW8U+IR0Uq3yQm+fpJCBvI4xkXeVV
cRH6n8BarFwetdSXqUcEQVFGGW+72iUXv+u/EpcXULqdkjQqgw4gIawghiclq5Y4
AOpPfPZN0DNuLN/GIXgauHUxL9D20NVTuC8n9He9rJj0pPVTwLPbOxTuIKBpYjf+
ntCVvVIP+lr0gmXpV/n9TMu2He/xbLajj4AU5FWZ3u/3yMDf+RRu1PxfidAkNwzK
pWCGaNHUEBVo745Vi4LiFtZpK+DMVOUP0EFmW0ly5zK2BTCNJEmOMxNDfBGxWss1
fQwOtldWj/nPsC1AlREL5um/GM2TGRSBYfPnA9ym7nzhZTduGS8lHFRRzYh36mTG
4M2GH1VM5kKeMsJTGuEbQjJ/tYpcARymzZKcFBxdxQ4oz8enN+Wa47O3ZRqfoFF/
5WctQp+ud79fBxe9NVityjuLArEp/g72WtAJXubLDSKgu91Umr6OqrtZanT/as1O
6ym4NOxnfZZom23BJs/L3vCheVmskJgwtw+KHXOd+3RkXijxHqvLBGi7hESExbR4
qCtkx6NRigIxs9C4s7pIeBPeRQT8TpiL16iFMcgdoBd8D0SLF71rma6syEFaWs36
iHP8zS/iwjRNIm+kqNCJf4c7it2TvSapwKydYIV7p3jLTp7hza3IGk4Ke6k2Go7j
Bsgts7wGXKELl3T6D3v05Pg5CW4ZBxuVKA/GhXUuQCacIYbNZ05SWieISWwRcYn/
wlar9J1qiMq3kMOwABVvwV6lvHqpP3G0Bwbt7FoqAXSf4KB5Exvpj9YPdaQj9GoA
gGaEpFSLZclnHMgP8aPHUE1AimaPaiSFJZaHSHb334sTtdsuJVZTX/kZckYolj3w
lhk9E6hyCq8vZ9re2ZGlAxrce4VfntrL5k825h+F2s7IvnLoOs6DnxgmaZmyp6O3
wQuaEONkRfcLwAXacUI0o5SQDaNfJyKLJUmKdRpegm511PFCfDNwDTO5hnFEfO5K
rNSFcAmK/1YNCBPqlTT0xsfPhQncls5Ii1uLRt+c5OYVQMqrXzgk4EUJO487Yfzz
1Y1McZeyDLcLMHQ3YwX5dWepMXqvCc1M0L9zTKYNsK5RLiwwiVsVSxuFLrqBMDrR
KXE4qogSNwtnAolMJm3Dm51TznNRJka8WmIFmfvwNFne+L1d3QlD9DfrzS4ZAUWL
qW5rkajBkrwbn+UGLgz4ucnPO6BcxckZ/uW4/pcZpKvup7mqz5Q1iWdLCPCEul3L
dgTEuXsM7YQuGEoEk+BTXand+Dj6Kq0WtZm8zhIOOxdxcFkGiTfa2pSoCuq1fXAM
VaxF9776HU7hLI41tYKChKk1W5KN3FQefVoMVh5ylQ5ZEai4NR47I/2XlMeH29sn
/Fy/udvqk2Rx82D6tG/JEF9Zquy8oSk5avPaUGqboYHtrwOQ2Dv7YYMY7yAT+EsE
gQozvFj6f6p0iafWTuUOOyJhACMKrI2/n8jBtIOveeCBTBEhFLQtpxsHTqKwAnvL
QOJYC0F8NDiVRk4gIA1Q4OOIKfbSaLa0pUrIqN4RI+iHQXO6acF5W395Htfr0Chb
fdNdrpO1h7Sy/QrTNHl5BEMNMhbxVnQO0+2Ym74FmIG4WlEH5gVXnqJeisuZY80Y
07Dz/mgdk/ajBCeBYUh7HV1/RgnB4s2g9on8JOFOyDx/3sh+eRxFhoHqP9IH6QAv
ViIA96TtTDE4CsB0T8JASmJluE3JyPchoNLXEQS/wjE17PA07fDHG/dGLeSGn/dI
q4axDz5D+mwCpBTClJNJ383W2D98d9NMD+HyC83CGuPKOjgefxTc5NWrCljm+XIf
pSxTczWQvDQlWPSIVL1EIZahgNQiYKixPtIhUs0r9AZWG/Uq4p75RQZHxLc0hPhQ
W9Lsi0FLGte9cRFLNI1hEvZPbgy7noS4ifMQ4dMtf/M4dorwpwKIvumvxFvS+0Tj
RlEERZnyv0gEeTz3YkwiwJJcfZG6H0o7caT5nfFuTw3L1rIUMLLtTcZM6sai8EOr
Oqx4smqbA655iFD54LRddS1P0oQA1YGUUcA6w4tvFO0QgLjp46S5zn0mRAeHSnEm
Ft9PjCkFYp6nORuK2paLaxEQdJ5jvxLtm/kivUu2Tcr/43Yzx7gGlsDHSRS23Mvl
j5UydX4oioIxOE4B8qq3+tJ1+NYZUFYPXHhQx8rXm4EOAT/wWSc62ZGdUzXqsRdu
tmrAU1PGks+ZZ3SSgqdX3NXzyALpmHflaefzvcmOHVomT5h/caZB6MwrMod5i5iY
vbAndIXUsCYQ8dHSnZZBPDrv9+Q2BLMBufAr29KRGUbxU8euB8ntasm3jVsCJTuH
Nru+swLRaY8vDQJR3qallmEVw17+/BuaRca7GXn8ZORsoHnlDMTBvpvr0U9OpWyG
3xCmdzV9GDLjNHZOkktp/sE/e/PMFc0zGzaaeIHLqQt232QEn0YPeasm4+l38cL/
Z/efrmlWrkVPHO/Lco5w4V5iOPwln4y/zi028STKq1f6EynvRFA8k/tRTmr4RGtb
yZKx8HJXV4YqRLc0BVQNK5P5LPPYVMJx2P4VVXyzUJdvKkDm/BUKWbv/dnoO0Omc
ySzhwCq1V0TX5ARqvylSmGIFyAl06MxWj3y+xjONmOjwkWI0aOhTBtthGdAFAy8H
8pFPxecHKQSjvk5ZLpReduQeONPKSf+mn9T4ydg2U7CQ8jUN1wTJdmydEzAqJtIw
YonCyvpJk9pGGsJ5Ynln5jv4VbOhbkTM7alwMJmbsQUuXau2UWIzx+Glb69k1QLX
kWyILwYqLbuPbKK8vBGr5J+2RzksJlAtrLExUyPHi/dXqwsBuWF2gWUk7amuwNVW
EPAa2Zlqvvntm7VoJMuAPP6nOG2HVmVatbZbO6pSGsmwNSa478dWJ4LOMlYrJcu9
Iy3NFFtOYjhjM5aybXceluJnybF8+MAsFzxaheUmehWFSGQxXMYCUUqH4HZL+kWv
0qwdoW2acijPz14uZbzittmGR1s/H6U6Ci51IgaOuUhEf72onPuoTmraENOmQ5zE
KbdYQZoCm2wpvkgYL7RrAS/VWg2De7B+ntj+/h+1bNaLbzpmgCyVsmD3ltF/3Y9G
JR6LePnof0OIGNPmVqH4r5xul0dC4aB7p4rGCFUi+PpuEX1AHw0/XQrlq6UEHHAG
KNXCaPc33veAXFHLBgBp6Ld0LSDmTK8uBCVnt+2reVooNF83lnKt7CNPpq/zOEkV
MI6ciBzo5s5CGzvw2O10dyNIqfDUZPRahmB3pJn2Xp/vGHlzzdxWaB/DtYBOR+S4
t7ReFD+x4Hrrq6t1ipxk5JdXfaMrLJjFLO5lww1VSiy9zOc5ic0VLcP9Yh+PTgwx
EaVjRneDn9pgFkyKHMsgui/KPJ3Kex8Enu0dCiEOtMoEwrWhamwdpM+U+jwcZ8Yf
AtRE7/fPv3m3qveWRX4yrZolhQmz1EW5kktNm9ulivzjvYXb4MVd0jehrHa4/TPS
LI/vFowczDUD0fLPuqkac6MfyRfKnsCJ2FWn+dQp/aL0HF8wVDIUgifX85hO06bI
wB0Jb/30uocCgxDaEuLJAAfloM3d89FGh59TMGOreqKYVZmBT5LbSAAvbOzhffm4
OPcN0R0Xbaq/2Jmv1H0i1O0bjEMUtb4k8QPPjxK62+35Ew6Ev9wiaOBo5/Sbhi3J
s09wNQ6QSE9JrIjrw/j92JkrJyoBRQsFpJsknfofHFeUOX/8LOlwRJusQz1Z9vaU
VbbpYlTRhI9Nbf0mKDEhim8G2TrpLKiJa499e8lIHtGQHEyFwX+ukbXKNe97vxNJ
m3w91FQ6Rbt+I4M+gzcb8LmZabTi7sJqxKgcmKffiY2CKj5frt88HDTYEfOO9UYl
+V2/0dCIbTlY+b25akzPu3h/smjo5PGsicTd/CPp/G1PNy2FYs5B0348t0OPtxsy
ZP4tV1N2Z0oVLbs/TTUlLmltJzMUfb/z7BmAofDWDPrMFbe5dcH2ESnBGhdv3KhW
ERuXzE+0SXkT8TMYwKlPXGHvduYn5VZjR5lFKPFs90FYRXxJB0vsYLw1brCzr+fT
Scua+8/5JTv/7hztS0OxPQIPkCRInMqNmRkORb9T3/cO1Z3exOUQ81tX7HMrgHC/
4y9eI2A3ciXbUnuV8FepLeiCb7zKgtXU8K67dgLV+1Sln5jV7G6MHaKO4lw0Iawm
wcdk+OfGq6ofYXndy45YyBucRnqpMQ3x1jkvrQ7Onp5Hg7SEh3YGFoMcCOYcmGAq
tuwbheADoEIf0tsaQs5UTivNeAP8Xk5NtEyVXU9lXKIbXPXN6myyLBvjHgDf8JpA
DuqYQ2NTFqIl7arQdeQFBjmTH7bSI4mx1KNW1E1D7+j+QXO0kTw8csX+rxBFts/p
GGEhH3pHW5QQZJv48ULxkGrJ2c7q6m1K6jqsatfI+w9hJVXu8zaaQK7KK9/AM64M
PnLR2YCqmFr0qeAxMXGNN9jiYY+Q/BlzVpn/Iw/MIffVAA+w79wxAClghzxFJZhe
m99fXP0oYWMoBP84s8WiyaXLCJDR71GVa66TcEpZynNfgFJTRWnOAY7wrhx0xNXo
A8d/AqEExwOo6G7ZI9Ra4vffeuObCiLfErqO4HGr3pxHNOkF2oP4MWYa84fWov0v
Xi2NRAGv4Fp2kUkQdR5OkNnJ+64vsdOp0HwVy79arJqTlGt2ncNX00LIYmNsesis
wJIRc+QzF1JhXvn/KE91LGqfv+CW7l98icdQeqmnZqsPReqs/WZSVRyQvueN0zVO
nfm7IoUdUN66BMcF5e76ptbJEyWR1/dv5qUUGwTjjrFZxFANaa9DUkeSPO4nRMfW
fT5m2hWuMpxx/wEYDftzJYc+BtdkSRZNLXNSgHh8pWjzCjp2l59kYdnaXL9lBpNd
SRpAPWxGIsfTZj3iOVsKp6rLWgP4AQjNCmPxpNsQ8S2Ba97hlt/opGFEHUS4/Xnf
FSoNGjacJxOxDHrLahGObx5Ww1J1ayD0uFN5lQy6aCvBvZOH0fOhY84rdF8KKcvE
z3NEGQaRQZn+bJX4c+gpsrU1IPCT58FpnScIfSp77liBCwFBdXJgiGwcPwCdSGbQ
7LVp4Z+ta7MOPcuHISfWET4U6f29ppBXvXfJgnzhaQl68dPV5p1RSkM7cuQpXekN
L6SeEIWrSMHZXRT790qvLJ1X8hkRXatnE8o6f7MV59V8OfAGFkyknVFlTMcVFat3
xgLH6YduHE1rMk7nIcmbbk8m65Vn6HHPfuqglpau+NUYkMsSgfGJDw21AEXrUn98
yDCFJ3HSZkb1k3X/pZKpIGBXuJt60L4P3zqOD/XoJKVrWo6JqljmMdCfpI9uEo/1
pS3KQ3N5ZyfRkHgGdYA7K7mDEtHepyDqt7qGHQ7bCa8qbikCoiL+3vJzHG3Jpc+X
NxVsc5Y8R9CQzpKqyTH3bsY0RhzJDADqC+PzRaun6Zq2T9Q1kpjNRT2RQF//5Smy
kE07Dm39Eo14rSIawzvDyvmVcCsP+ModVhsbp9z0Tba8zj7Gt5Sv2UU8uJ91fhji
SklQQV/jEQEKoorxmgPwsfiI5QEq+2bOvUYL9dQPPvqstaxaZls0BGkP4lSx3QJQ
9FoeiwJCeTX8jkL57p17Igqoy2TJsKv8gfCufPhd5R+1Bmj14GnAwbaKNRd4l5dy
hqWiKKAfmosnDkumDyJDi6RN6FLS4fHYbLL6VtSv7fyYepEmr1rl0kdBFbN3C9HH
EggsHGLPzis5E0TTyeQ4wJh9Hb1lqwB3MsTnVxNDu5EBqTSRhxfjyD+KTwoNJyQt
S6Y6DvG3gl7BN6zKg8wegnIder0mwtM1gyO2vN46zh8HT+uYs6w2weXYbGMVu44K
IUHOZZqgtMwHGjhMAE2JLfb/VdiFYYD4Bz+pVIjBSljM56RYwPEAj+Bv/eqJTmxg
TkTh4YLfXTOXhwucXnnFiNlxNWr2G428WQE9NJKp54UBcT45lA6v56YQjdqXzBEf
zrg55zlY6L0pbeC7EqviMeqzW5PI7tgtnSP26ekTK1alD4PlOOKSE5it5YjrCTPL
WzMLcmcRI9HtCazGLktYLM+d6NepiPkSC+D8RO6DjH2gEOKswajKgMyNdJkN0OT/
3I37eKfO5xZhMIsgZLmF0owylJNDHiXnZ4l/7k5abXE5vxgwdU3K0C+34ad2X0i6
WrrXbPxSqVl3WexVdvKfTho3oVJ2OzuLPQmsUMUr32oPvDtgbUVhd8tj4UuMA/IV
RQM6aLmsiEhXXsZsxov2EwnsswIKcZgdyLnPtKt2tqOdt+sRwiaLgvMLxBddCDJK
j0a9MuTzTZB0tM8pgrFzBrlh2bgrKUS4cnOV05kOuUss0TJ8MVWyxS+KYK4crjWZ
fdfktc82XSMEF1+0xgRp5mL1WRaRD/7Cw/oetN3OsYCktoM4ostQ3370fjx3OJKe
1bVp9HpQhzZBPH/ak3u46dIXwwExbmEqR7rcJsafV92qZYSS9U/TnmBOQCekVMFp
DdAEjUbYMmhCHInUXy98ktTLiXODjznz5XZARxYJL4MJo9Ly8IXwajA/Aqf50QvQ
XaZYvjTao3stdMzTniP3CTo3tG0/ktEUtaM2NyCNF+OHhFEOR5v7iOrPmhkjmnYz
hntlDTN5EUD83BHJYxCCXCRJuqLotaJb+GesCe3KwcLye0Uf1+ztU/XvDlcrI3Y6
Eo0lMHwF3YHLW2cGC36z2YaapglfO9HYuYspQTUAl3Zq5Hy0nmtUrYpYHaMZaodc
jZfG/nVZFbeRoj6I7RUN8sHsSZt6+ci2vdnlMIc45kQbzuFPKrNwMzNig5MjLtqH
NdZYIlvgG34i/nzzcwVM/2NudqsfjoDBMFRczVvmSSmYBMWUGzi3SpKE3cH4hoCd
Ep4ZlU2rD1U9McGLxJphcPM+BU/EO/Z2WaYopsZg9R1kDTGgoPaILk+J6EqnHJdG
jqKXmFKUU8qCXfbia6W2ZAlrXzfyfaPPiwr/Oi184KnBdfJ4Bd4gteB9UGfuoY2h
1lIkDsVuP3KzGR6jzQxUX95xJ8nhSx2UyCkPtCjQQNVMfFt/4OqSCbsSKLKbbuRF
m7r/vcTWz0GJJJP2PiXrpZ1tLe0W5vXTKsvsxjq5SiG7JonFd3K+Dfe19MbPKdBT
YnBJkYIKc1h1hMdoMr7B9OrPso/e1CLyPn+rtng+ixAbbQ4n9vEQISoakEg97k+p
rTbMNi8lQcowbcJOSug/Ku2rVTltDvyVFdsuJQg0oDeIa/yXGLvxMOxd9NjJEBGV
Jk8mkFykTywfdkj446/bFL0fLUf4vAJq2bXLEOIr9Y/9e0ww+MKQkF3XWDLeNtZk
JBd7B7PPnrJ4KfvG4o5Ji6A/QL5AvFl0/Tp12kXLC38ei3uTctnkJ4VJiDw2eNof
DvUeRQoxsrJwAffDk15w0OmdiQKzWi6ubRHB277tDLKu7eHM186jbEXAz5+hjmvr
kYSHC1pbtOm0EOZWYyi2PSVEx6Q2QXdyU1mUlL45BtKliE8eEjO+zgyY10gtJAxL
/VY8SRl2dLtxjYk/cqKbtY+piBnkI1xefFXQ4gCPkOkkKK4g3FRg18H2xqBOJ3Xg
EaHTriTy9d1FvaC0AZ2JWtSD1pobLWL6qzieVgv8X/lfSQEjrBzgznbKVudt/VQZ
nkBkOat+38zEvitNiMWxtAXN9+i1lNW6q6mk24oUVLqnFsmQi/yJudlBZVuDSQMB
JRw5UzsHFfqz2kqxUZbr4OWsCN7e7oqWtXtF0iKdzl+Wgj+bQvBI/3bYdXyPZ652
xEjctRo3scm9W4BArj59Ho8srE2jDOsG3F7tAvjuLwV825SMICGdTlS5VG1ffaXA
ke+6cR6sP6ilMG7NNYuMBVmG71pUFtVsdekqO/3hWE3Tb8Yk/kTejmhUIEvNbf5r
06FzcE5m1p7qrfqtjSIJTmbJi88CcwELK+Z8zIdGkXeiovdRm69O1+q3McqpnRp5
epH6WQnA6VpMLuG0dhoN9+YXXeP/I9WYYzCbC1zrCSqV12RLCb9DaY88vBl2mcTS
mPkIT/s8MMzhoD2sgAURcwHd1rJMYL+ytoBGXcgOBnhT43M8XZEiGxvJJO5WslFJ
GAozgi8Y7IiXdJMqBMn75TMgFSYxYCbLRaRKTROoSeWbVL8bl6Es+Dt8nH34m8Y2
kYqnASjLk5gFOHRwwe1pbw90jNkMocSNZBZgb2H8v+6cCxjIY98WLftHGeHh6Tki
3B8Jur7vqiVvu/ZHsW621YuSuV8d6Jf2u2hvpUciecXDJAE9Rh2ITGOFqZEb05yy
GD35HXMD3gM/BUECHnuq7X2xuEdE8TK+Dy16HtwxanBHreshH+Uo7+eJFsqtKrBn
rqWhr1fz6IgKt/7GhpJ/nRiRhrjTceqgrEIABbUns0weGr/Tx0hFnOf6tNo6CaaK
Z11HswN86358atAAA9gytsH+2eql5PwCTIRoM8IEpzHYVAHH23rYfbh4pyRnKKfm
eThB7FwU7GMRJq0OOf3VtVWheMtIOugdUXzqy5rgLdXS3tQ7bkXfeOwFJzTZ3As2
3NtpFldW3dOlsf0V1HuWb8VNg0HgZeZ1+3J3oHdOrcQk2KTwTf0AK5A8SL0uqg/5
ofy30R9cE0GN5DnSvFNsfa42FBG4qLf8E7u/nYrehYhi5aJtkl8bpolNh/wMNeJ/
HE2Dd1zC9yiwKqlrDHtd4k3tDy0ZWqHFA1P/NXqLboo90YZD5Z1imHNUtIh5WB+f
7tn1iglVw1Sd+1m7BsM1//HeK38/cCtwrLpWLuQyaNh12jl3jEYzAYblET0R7Rbh
vcsUWwuSNX5WgHW9FJvIUI2AfF+NzXrLwrQy9drl7uahMeFYpnnthqjYb1pJp/z1
cXxkr9HFzG63NwVVzM+x6KXyKcBz3VZt2O8Yc1XndYmNi7OOENmd5Zg7nchkbryE
ew6a7IuoveEZUqYMPiF6ypDVswPEtkwspg8kSJWa0tVMc5vHM306zHjE5Fv4lduK
bez89jk+5SzySqNrKuyTOypIMaCqZojnxbMi4FeQ90LPDzihktU/4Ov0fKXPaSkE
MBbzK7JWjHzaaU+V6zQHA4sfup0CPIWYwUgLZImbZCGLMgwonh5xKAKveTKI1Lr/
Du88/4YkF3GK2Uo1R/ZLCsjB3SuWrwEx4fcXuNsf0+Zjim3ZilByPSIBDWOHcAFQ
gneg0HeldlpYgdNdlTtwlZTMhDEyuHEQUnGBaY2wnZMN7utvQw4EvMRT6ABBFeDX
e3dWMGorsh8P7dcjPz0zhSLQhlX0cgyBVyKaTeJwYNPHMz2ZWsbGopqffPs1h3Hn
VrQuHOwyRPYsQ77fhR9LM1roK5Y1KKOo7w0/iraFrFDTErC8KQZSLaqELfsmXcRE
IvSwR/ZPDQiqyJobShERlaAnOe+jeWUxiGYcZFWubcZHUGkmX72GC7JFUh4rBT4O
EjR/Dm1mJUQwW8z8DtFv7t3ESKzpRWylmHojVYgPiibpJvENsJx83Nj85K8tU8gj
M4DIVqDB+KD1MAg4pjbDPfxmf+JL5BvNxiyzIGfknzj1ImnJJjqv4R3trM5wFtg3
ndgI7LOoUDQ7pNQMYM7ezyHqimSeUXUrlf9LlyBXP41d/MgCBGq6Ge1724IHPnwk
PrEaeGm6qIUx79SHte2WAvpLWqyn+HoKmvoFCO1kwFNa+210i6wqJBgtGVC8eqU7
lR/Xu0gyr8Rzz4L7wCRf29X0LqRgBh8z8UyuYXurPFZ3ZEInJVu5XCmPQ9QQiTEE
EGR8i9qjXACjP3m/q1kxjIaCGh0ryWoGY/D4UGsjBS6Krai22HRlEszKAi5bMMcZ
XOGGhIfGFhSSviRWGgdZrMoz+FisDp2k4Fx7l3k5Ircn+jq5E8ZeqbEbrQBIpnXx
OjuY/MyFsEPvrnNqcFvLbzB1xcNyT9au1pirKR0VYIvhjeoCti8eCgBBdCrH14t7
0QkVkMnAyLgWnVdf35KhaLPIZ9+5MrBYWnO+5sjTkxOsOElzACCZRBDV9KOtd2fa
CRJOWTcy+eH/lX8wpyi2g58yO0zvUyPFXGgmZHP8XTUxsjuCpeQJL9wWxoQ482s7
2IzFh+3yN6u0IYHciq9azjUSkxHg26rqHPTvxIP2OjkmZuXL5yqhiBhX5DULPQG9
0brjwO4QqE4h+C7BWTce5uTU8/2FfBkghrsST2wzDh/rh8xnKYunLxGSjRFTjRQJ
Gc6FiM9WrGCKoJaveXqRDBLcQQ/ikYIQ0u86ZTVkmRkWkR4L4iXaZ15Sxlp9C/w+
HWj4+kgZ8ZDwgdGFmnM3YHPmAPBbN+gNSXVXt087pFL7n6lhINJwALBrzvfbFWV6
VHIrXmPkBr7oMCz/2w5/MsJT0Hj9hK1xXHyWODYEbkLElYTRU8x7psc3Q2cG/mMw
cIgez+D418TcbZRTI0XgfAOiSC5Sjw9UwjDSDesHGZntj/jhEchsrxZvh1fgxS2e
6t8MkOUFfuZp+0atRUEQMgNbI1gZh0hQ1HyiAFMC9T5yNIcQ0202YRYSafumZ4zk
X4KDSiZIHF9Hq+jM39WZEO7tTMsTu5+KYTJ4SF87jl2S9SMvYpsTRi+ZR9UqMtKQ
XZPpYRL2nbJxBo+mU7yOWOrkeTIEzz1XlZw3C2P9llAvsCa7CeB1yQAeZKK8/vLS
T+jmWCVbzYiCOtQwMpsLZIBL1qinH1VEZjQyRg2q3xTO+LH4INR+5KIqPPQPgE0e
IzfCte7SuBIgJbXXruaW3jzLRK+C/Dn92H2+AJK3Ri///6tTiNwPK9mHdn68xTC1
PoQ9LPjpUbdnLghXCMhHYOs2cMYAVMMVeTQfxNcYHypfPeW3Q+f2E0rNMbn6AH9U
X2vxTeUE0ADAq3WQqMRv6bir3WznEO/JM/uf1rRct4cT7GZlYOWAK0o/ipMWti46
QClO4Tozu1ngh+1xfTZXgwzv45CyUDcniq4g4tkvM8eD520mBGIDtT+Dlz+o7JNP
xBkhe9dIamoC1DRR05EFhxMNYwS3eAMWRypI4ZzoGg5wwCiyNSV7QWAE3W2WHhHA
+A3sGprLX5y+FZ7D56c8TV0pGuGgfsxh8dF4fdYx615ecGi9EhM2bKKX/Gy+EOuk
5TF1luBgErPasH3ECjJ+qIIVVoLneKILvUmX7B1DseqQVqmvNvvXxoJmsgGxVzNP
6okrtu6t2c/jaakgeEQ2sptLgFV9nAiez8a4VKIhWQ8XVval+zcsqAg/8M9qm9no
rDBjkF6//+B91oPxOGv7DcWN/UquUxjzcnEN+e2msFQpO7IaHDOGiiwuF694qH9A
PmW/6YJhTdloQkHeynZKzN+ytz3o3I7M3tV2b7BZv4X28ra0oUeaHC8RlYyxtNrh
NyaNA8A4AWQvbJF5ThBCcCtmjIySUw1P11MoNLMNBb9w87Kt/3dxZDB8ODy5W42c
VmUQ8CK09lBV3xjmKm4SXLgppDiubAg04owkyti38Z+2htRHTd3dOfU9bOCXvaWF
t20gOckFvI4mAz6pnl7TPKRlfQIz0NZDic7MesxHmSwjesswii6dIsjSyEClVX3T
T9f8BRiF3Tt0YFpU2lEjijZZcCLYqQzn78xvZ+zzaBV/38122G1Oe1tQh8KX7yyD
83kVyUF0lztL5rDyFDqPMMC1hp8xu0cLdUNEbhjd6D5MqDcb5y2wC6YdMXeMckm4
uCBewc4y6jaAM1YsZVEQRBxu5P5M/0MFRD2u4zovZoO0lrvi82kA1SFabNjYxQ8y
s8LAqlmau2csFqZjf4qGo8XPYdvQ0Xp/PmzxdtleWTn7BB51gCuRJJfQ5DK+0ecL
UD/lOqhsWofDGxUTxvdOI2RC60IXhsc/lSc2QrrxKMmUw3PMosf3Dbdt2d+h/IcC
OZFGMVlq3zJnjEgFbUdjvdSZ6tcHOWUh2Pv43W/zoFFKKkZqDXkovN+JOZDM+IDg
4RsU0ZTvRnY4JLGBRd4LOadVN7il6a1m52wd1GEbnYeQEYGWTBoOgpUVbskJokpo
9g2ljCitXz0AHgZ50I1KoMd9MV83prLG7/zY2BA4ly6hsW0InkQdOpfuJJ0rPox3
NmZPTtEwnrO/bzBfNcnhYKpTXK+F23URz1JiAkkeJ+Lutca+lnaXVm84nnx6InAs
zK4yTxiEg4q3+ZdLI4fns7MFrEpqJKBypY/rISowMIZXDFZ0CyM7tIHZ05NSKTlW
xRrhXrPosnVw7EoxDM4vi2eJ1eJUpDXkiwnv7sXBPHhyCkpaQgC/WDsP8Tw4Pet2
u8arqjNyNH0UAKfMnKqCYokqkyv/9xb8lz01Atc7lFYI71NcLf7aslcPnU2dayTj
26htJ8vMrZO8UnDEJxTkf93drPotiovePyWcVsZbqpuAfoB5Nc1dawagymO3FIJn
fnyHGK3WeKxK0Z+wY63mcvPk0kKtpxOxkHziPao3XNOO2lTNl7If/CooVW9zkjXv
8byllsPNJnCVXZXLOWjR4I8WcOqCecuxfCWSFQPkOlZuh6FoK84DLs5DbVFHN2i0
FwJj1+k6/qSCZPpjGQ+WictnPAYNxKQP4bMv0Fk/N3t8dIEbxIijhYuRsKNrA2cG
8W6IY7sQgEVveG2bqUyIcRdU1dRVRi/P6nqVIHoK0BBw1NQ26ZV+mCYjMM9fVK+4
fwxnaaLroSnQBxsQdtcrZr7k7Swzh5tm3xxdALRAHKMv+rq7DUq2YRwAR+2mI+QV
QyplNPEq1/ufcKKMyfSwJWcAUcPxtN5ytk7+IXk1KNAKw1cr6bzZKFSmPfOpzf8q
XwM9jj4hhv4j37r7Cl63zSNAliDaecJUWK9PEl4nfyE5kWqaAuwNTSftSYWPETJo
YHMQ+YVtn2Nx3ccwiUENV773gYmr921b1lnRn8kiojINvIB++ZwKdARts+jggWog
LSytz1AMqIuEW44QsWOXbN349wmq7KwTOnykUw+CrPo2BEu2hELTL2zo5iXXr8p1
WHAzmvOnGiBj9FiPgLwlEdFKI68QPDxoSqUdlR8SQ9qUHoZnE5NpHvj8HDNahve+
r7aXONfQL3sY6fqTSGuX/5sTcLVRRY9oN4NwQPhU79mF1aYCAsD4hkQAzIqHxlGu
Lo1z8ji0W3QjNb8EGMQam2eX/PXzWpInIrYnIMk26FTrtY6VnFpBITeQWJ4PTYN4
7WxJx0FUlQc8wpufGlK6mIa5xbAKhYyI8rLJWVHzWbQQXF79HZTvZc7ewdTjZtvE
1x9LDfohMlB9gkNTnnRnl4WuIvnqKXklSyt9oXb1CuC6HcujbYhdK+KuJPT0YLVV
RsbA0Xhe6TDr/FW2bDGQqlQSbNC9qjtDXjqhc8fcK7FiCnqvzKnFRuaazhato5qD
ewgnxO6mj6hWU3H+istIaNKdYCg9CHR7QQGUgCCj3hlV6JaQzgko/c7sFohKT8VR
n4yUurzakOrQBLezXdYMprfy99kBMtwYnU58w53DzvPlYTcP8wAMPGtfYAWMhkKk
ZDMy68sqYDqIv24K5z/GAzDYPmSBfkiyrg7eyqCfb9fMGKmQxD6ds60UggkTXl1E
i2m2hNXVVax3b6wNqQ/HG17opaZS2eSngVO0ebEAhFhUWB027cLoEyHijPOHfRIi
QwIJ9JF7rCfQviHpVmAi6JH0QFT/u26tiELKwS5/XsOvciRMHwsRRe4FtFCepg1L
a/gqLpxyNTsFp/BKM5RRyrVFwaf8a95BA9UAu+/qgKVvHaHNBSz5dBSu8nwS1o4z
Pyyje82jCKbJFZzqE9JOjTDdP++YHpOww2Am/UzMNvzdiFRvE0mdehTYelGc0ZkF
mS90Y7ierEZB52y+KM68OhHXF2kikOv5w/rL10i3HMrk544xdG5+7Iq9hps+ZgB9
sGGl/RJ2e11x5D8297ZNqWGpY2TByShcRK6Xwik7aVi2wVnBFYBzjz1gpqxcgHkS
WOsy3rmxA2z8Ym8LQgw2criIyccSKl7Bjzi2VrTSIHtYDOg1LSsA2xb8XjH5aYtx
oy5kUkgDDxu1xj0C6ZsKLw3JVTwMf31YlspPGi34wH4eVkgImh1BkCgDF8ybbYzC
zXSvhKY+5lTcFrs/hGPA1GSFH4WRAk/gIMwBBjZXY6yeyq6Gtn8xhPCPzfxGU1sf
nLkeUWDgk78IhRUPGmyr4TL+h9ITFKkDLbvxTXHA45irKQlY4VsN6mYttqhUvqR1
MGKqy3Jmfm+w8Dk8XCuRmXbgdrgI1CoCu/9rSRL29gNIysNri5aR6Jxm2ZquwDV0
NEfmzTi/pv2vaGx2T6rsMr4xtwx1uU2pl6eCekId9X1bcfiJMy8k++uCYT+EPKZV
a71O/t1/PqpgBNiZFQgxF+8n3w81/GCpk2paNgoTEOg19bPIimQM98V8rpW2/CBe
pVGgwOjnnlANa65jVD1CMp01UqJ/HZ5M09SeO4ue3SL1t2PDYkNbr3Q04VbAYbpv
FlyaDRn7ofVQKtqi8j17TLWBg3iKm3+H2XroUC0jJlcEILID7W7mYpYth5Fa3nua
P9fOJokwDNcqom20CHMEow==
//pragma protect end_data_block
//pragma protect digest_block
SgsR5OIbNklWW3ocpj8dCj51Kic=
//pragma protect end_digest_block
//pragma protect end_protected
