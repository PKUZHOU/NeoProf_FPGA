// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
JyB2GWTxZJTj7AwrePdd729m3fly49ywNM1eXgqQr8kpKCWT/0QbwdsOgQ39
yFOOxyTtS+MQiA3mhrTYtf5enG3xwMuoLt8vCFR/H5BRcvEl9gANOE84lP5W
1ov0Wg4bBMFeiupqDuGH1YFNxdVsiHI9bpbroJXdxDmR8widKjZCe48gQl8n
5PMEboU6FVnZr9HW/6jQZKidhtm4Srv5BWAl96FG0zxqUEKybEZvPqGfzlh5
SHeJb5bfEVIDAajj76Iz98pbmC+ZR/Zy7Oi0f6cqv86Zm82qg/kORe13PPpD
KPT17OxE6bql2lWZLF1aCsve20wRzAx5U8uMJ18Osg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
M4kkFzecs7CQimv2JIAagJJTapR7koVrXvqZ9C+rEIXmEIwWSRkH+B6JWs3K
3CgcM4W7jWUHwyLpfyo3XxzatQpCEvguKcquVo/fYdA6dJgdKYL5aEWnhOIF
ssB3f7ARGdD9mFKbWBaqTDb2qTG0u11Q8D9mvuoMyKKcMCKNBPBDrHkZMVq8
wlU2noLUPBnr1mMA0t0eTKxC6ar/TtorhuRoriL1zFXeeIJjloNEbeyjYPms
wgKr2kcfJGCuPEZ8H1iG06GO95jRNxXzATNNIJX1vwNM/9+AUYGqc/GFqbAW
EO5v/g2cr+BzNdEkqC+MPuYjTxFDUpmNQXehE8nnAA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
VNIGFUUi5LJxa/2FJ3RBjiWOpMd3hotLqB1tKM1BJc8dsEE+w8ACPfw9DgIl
5ItEZW4laDlS9+gM6Q9KH6uUxoCVbePWgGRcXuh7dTcBFEoxOywWQCRqNn6G
4yyoQV/xn+IArw9LkdQG+O/k2Ufs68khmmcs4elH5YA+h8paHLHt042iJYue
MMq30cbBKmFYrBYmMP/RI6FuVlsqZBPVQV4raM4M6IUO8Yo0DEa7JmYKDQJ5
Rp6Im+fZ9+cDnN76Kiaahkkntjn1KBi5uQnMWcS/yfCdV4Y9BUGjkxiWl9qb
OctI1+F/nBIi843dB2wgnyjx3eHX7GCaRkJpLwXiLw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
QvSvJYZwrkRghZ58U8DQoC1zhHVK2bsNPAVTViP1b9Uy6QWnUgD8PbU29In9
f2ZkJOBsgPtzPdpgaxXIM9UySA4lOqU+yoqSMXRDsm0WNGJGKRnEhCF0i1UK
eSDBlu44UKlgO7aRwRWnsPcoLp9cJKuIfnIux4l6My8xGQ/33hM=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
mqwvmp/1B3jCYiG29YaG/mMUwtNObilVHy6ZDouiHLRX43xaNSTCf/h72BDl
Fqk9qfRPy9JFt+wj+ud+SL1fYzKH2JdV/IOZ/sQEoFx2QlQLlXR1KE2Gm4wv
KCzRcrUEM+Fc7NUiQ/WuucLLZ4UX4CS4rLx0mwytccsNh7XceFw3LAyGZep7
CccxBduS6Z4cVMSIFZuh0MdCKFra34paVjW4MHO6Dfplc3yFg1tIbAVLOMpv
NUn2vWa6yMjR8s5RDiucWx52OCMfRgTacIj/v28wqbN8k+UFNqRWme0w5qbH
DP6WXdU+LwVN+UMJhofE6RZDHFOqud3LAzw/hlZI5YVcjmqWlwS/RcwQySP2
8MWjaYKKFROdkxSAETCjYghj1cu48yyS94mZyGUK0l85/wm/IIyRyz0D5hIN
3Q3YN8iAdtzzy4Dnip2vnELSKlnDonMO0EChJtygkq2S3MTMBGtRiH0ltr+M
MK6rYn0In0bsZ7wvKlptUVbNuKjLEfgC


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
m7mtLAlSsH0U2kLMaNTF39inue3DsR+BqSXoFlR8Av7fSJ+cTeEyGCHNU/M1
nTfcElNpcdFtTYzPLYNL7FDvbjiVEN50TYJOn5wADC+kAdNdLS5iUGbaaykv
irUpqq4glVuAK+Uwtvy8x5v0IXdlFB4xNvAi+bbqKxKPLS4/hQk=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
p3u2G94HvJ2Z40RFZI7U/olECrYJrc180veb4nKxWTTNBvjNlhdz1hDKLRYI
Gyg3ATYv6iroxe7bN8/ox39IDjRtOjWe+BLMDbibT3K5yOQOUOwsRZ3dRGGT
jT07Hs2rOKNSKLci6O2oUXIWCmzQgXZUDwT6+RH+eSjg3/QNORQ=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 6608)
`pragma protect data_block
lvrRzjWqSoxSznTJje9DRu5oxOHzSubcf7mCnJDz889bo0FZya4HNg9DO954
1yYPB17RhNcPF9rbRoiXbtN2vEapRzCZPKXw19FKPVo3jcJOjiarVc/utjbZ
De7o1jsVR35nPv55jqXUgP8Dy+HwN4bj/tLYlrtwokiXp/DQp4XS26GS4W3y
rB73BDUxUzcplC2Spo1wR50l7tb7n16MNsfuAHu1EYu59Rqe8ArpBqP9o8U4
TOdY0JoU5aL30TK7Qbf8s0wQYyAbhN3YnABHRQ70Y4LxGcAZGxmTL+yBHTlC
lmb4B9xEkBLkt0sznraZtoHtk6T+vNm9gLeoQLF31CieV8gkFUtN2HZxiDd1
OXbYKij3+xB/LEZZYcF/TKCIjQ+vTlDIsFNayVVkwFpmVkk5Fa/V1vaoWFOk
OHoWyWbMAj9w7AKGk0EgzM+b81isuPSxF/9gn0KVxUxxMkZZEJg+A52U05lc
Tnp25cUVuCXQVBLSK4i6QGaGbzMoozlHg0e6aRuVL1nm7tgF3b7dviwEQkQj
Wc0cks4PS9Ess9Rtzrt5XpVQsKhk7b7tV1kP8AQhIFRA/x7yxwXn0lDfV+vJ
JNk671JbiDPtWKGEXLp+gCkIGdjxUAcBJbTdxyYdJH0zX6Liyxid6gasMj+z
6IGPsN8luf+lBabgyGOPR2N+83RiC2+jfr4hANuGeh3dw+HKjCF3CJ61Kr6g
yZxDcb4dGl2QjgYpHYPr2T+se8rVVUrNPB+gjEdJge2oWb49btpT4uasamRt
mHQX8wEfXbj6/A0eIkqG2hYENm1GK4hiqwhD8AVc2wqJEakHoAyE24ncgeLB
VIm7Ou9sqQNidMcyboddZlhfFlX0KGuwzo+oSMbfw9W+GibCgw3ZWJHynTDe
+dict3HBkh0dvd0pDgnRSjN6YO1cHc9S7Ke38YMtcj78hW/h/hlE3S/+p9Yg
Nc7na6esQSMHgfzC1nliCvw770sHtHzsStcXD9SOsgV9TGJJIXq+hP8NycNy
vsMvlxgVWQlSWmlUTrr9G0n1sGNxGElQALNgWzkG4QZpUK758pwMvkOCrgmJ
46GXhN7RaFbwEOrLfRsHE0Y5FfnL42xC8B4eXTr1QOa/xjPBVeP5B8KOoD2N
qqwB07IKwevC+TqlZ0zuz/IiwUeU/Qemn8J+YMjilQTM1t1Eb/z+F0cAzRvc
Eff0A+pY5GEo7cdjFke3IXreD2O/jm1AeLYFC07wYHhsgxnCsM4Hip3pypAI
vVFgFkQ4lFokZ+qkI/6v197EULC8HMX2wtiKKSygdF+LYHAPEvX1oQUfJeic
pdaENXnDpgmtZdWOByZ+py89P2f5tZMR0QXe/GXQahW44H+BOymDJ5pciV3F
jO4JF7MX39yk7QAB+2Fk9krfkUM9560RHvHso90Xesh0jSnObBWEZSmT0O3Y
W5VBEQfIOUXXCyymRYfI8AWCl45Glz/rW4xGf+PcHHR9u0+7K1Ff+wMzE9Hg
2qY3VYpDs9z4gB21eqynmStDzR4mPHc7OAc1lE8YnJqCUtxO/TECSEhEOGBQ
byaLSQWzKmygOpS6swscnGrsKH0cKmZbSw8clVDMtX8kTLXz/UXqbcvgt5J/
YlTmtXtqRpxU6qLd3/n+aGx33PRhAPEnDXVFmJyC3n/AxU1NZ6kzGCVJGWoH
3G/RtdSo5+UIMKsmIlMjG5SyGBn+kGvC1VSeeUrOC9cJ93ROxWCN9yjV+Kfj
o5pgaIeM/YuVgRNdZkEVLL+6grw1LQI0ULW8VyrsR7ZlQq3godzn8mezau/l
VhQyM8c2zJsUBh3KMcRhRD1+s64CmXK5Uue3dFFuy3qLs5IQmgKcqSj5GhWz
e5isggPk1CdN+TvJxovxOM1Y4SDb4yYWu6z/DfIdcSpPmQSrKwyLUrOPStw2
wzRkCFg34q2it+x57XKcJ+Y1FelNC0o1N4dxzqteVDJLSR1CeTRWa6YSXRRS
7d457CXHHPkEdMxyqEXLbebhrTAcU1P+CdOjPxBj7PGC6lx7I0PJnQ83NQtC
CGv0L5ykCGcbIz1Ti0SIps0ppkrPgLAi8ZSLLzHC9BalOGZtIYdMc52224wd
1GU14QnOBW9kQpSmWmzwx/PWS67YhOEkAD2g8dUxVdPjvlg92EAAgbLWu0VL
jqIF7Rt6es6DLDHA7RAC4JFpe0ga5VhTwRGnhXsMCpz/6uw0CplSwOXqAY50
Ofq+9EaVcdPpYJ33i/Pbl8xePyfFqeNy1AsvKC/Nz8bK4Y2IXzulpBr52KCB
RhjBnCOrbhGnFnB8x9pzuYhY0r1ZGozsBHkQeGXY7zYgvrAv9Rmhc82zYDaZ
Gn+oB2/ZlHiMLlulLqV9GYK2k4Wmz2hOydvpEt1cGo5CHfTQXAmjZ6b4V73T
zfmDuwl4gPNfrUz5JcpwNYo6XwQGQi76o7x9p4jINIkTorAPhY6ZdOiDmH5Q
aRdt9E3IRNJJSHI+2X1VtVNhPKxnlQ8abkGy70vdheCqq0OhFGuo+p4UtAb9
2Y9sm/klqAQ/Fk45lIRP6hVbcMZRVEPnfqdT52VAM6SwgLFLFEFcVrlTwxkO
7EDOfgsauJkIC4e2vlz8D7hcEDKCHYAUSFZHOrtNaxVp/fhQyBnkvl0uMveA
Ah+w68u3bxbaCVRhYGTfRvbxgDbhEC1PjaRQuPuJAhDnGFeRPwpo27TJ2ABm
1K4wr565KWyULlnT1gQA1CS/fVB6DmLNS/EPaWGVX27lUwuw2kuZF7JK/iMq
R/8ZLuAQrJ5iONNxY9Rqk5bFrcWzx8T3Ti/V1vkNK60EPfdcsupa4r7kxlmI
MeUIWeY25j7KoKgRlALZO+ACwhaklGnyVUwZBIQsbc18F1F6MgSYhZHRdZg6
32qnAKEmNSgWYafqOSC+kbxR2+wdVyRrgbZKRK8khep+i3nLhHyuColoqBap
lovyA8v6ilNHc6ZPKc2MpPlDWo1yPdX9icH+Ga/vaus/W4AypmcVZMimXGDV
qg3Yx6N4E43lBOejdHe3+sJ6GRzXBTfn6tgoZAVbaW/KzJs5VrFMV7/0e7Ui
wm4tfCt6qpieWIMc/bAz0SvzKgHXRkNxWjOYeIE+Kd17cH/dz6fMItltPhmR
xk71ai27o/utyD5foh+1vWol/DyxOf03ql7idaKKC4nn8AKbmrKFclvEEFef
C4LkMQ0A0MlrurP6K8XbbepZGZi0bsZOrHgg9olCVl4pbckFIQkjaMd1uxM5
LB28CLIcBOrPPU441Y2jvP8IarYMO5pl8pNLqyXDqqBiBjPUBXDK1EG2Ivzn
XJGHEYeQs0B4H9pafWfagI5tgU+YdRYT75C6zkPgMdDqKq+dmZeGusg/LTOH
XNzm+gKtLxLUhGvcEUjNWaGIMu5fg2eKWk7hOtvwJNoA+QI8b70LxV0/XVoI
wPwadeU8dNcE4jQi7SBDNeavuwdyQ3qNBnma8Bj775TiKKwgSQgGFUjSuMf2
9WAly5c8GR2UEgOi6fluDmZcxSTAg4C4RaEIBGij+8iCfkt0Ffq6IIBrwvC8
IcjT/VtCyd36cB3iFupKwmW7H5/QNlmzpBUtFB+TAQE/YtYPO6BZp8LYk1je
It+HwevXKIZYBQNrXK0YUJqWHt3crnVmdcZ0jO3ePEyG7Ofw9hvDf5P3UWFy
nKQmgDiYPntwIyJnrQLUtMY8WCPsQkzNOK8o5uhq6ErrYu96K8bfephxHz4I
uTXibcl/Fs9GrclKlnPaWR5GMBBAU53m2J7GWLsNxBXqFj7Er5M85MqA9H7z
mbJnoI6uK+OSvMW/UwE0eTENRJWQw8FyGFsEvkYc0GF+Jlr+e7zmHq6Ew6jB
rFnr8dpKI04/fMiCQuZPcRn/lnJLqxrXPmEKh5s8b5Npb5lTWbd0A3YQ+aGy
meeBGbrW3ayyR9xc5zLPoaFQa3KE5pvPgjoOo6MFnl7mEd9tdqv2g3Kror/6
S/GxGWPpQEG14PFFUSaZ1T+Gy4C5F7BzQh+JAfVa3HHpHXUK5EfKj2c2QT7g
syGbiUBLNIAOORl/2g9fVsshiKbvXSHgF/LGWAeVo6ykp5URwqhBLo5sYl/7
uD03bdQ+dMi0jNwxbrvHUZVhJ8crwZMBsuccRO57J2A5QIiz/1mdLUiuHccy
gkcTnAagCXC4Pomq1+O2CnBjolXcJavUMSXeZuELw0YlC13CslTerJnT5D4W
bRLrymEDJDGiJpWucmKnYi69aXsjpMcc9Q4fJ+0mZYPjXglbZel8pc5+Xgi5
qySw/FGYgRZaox1ZvHJ1y9hhFyeH03UgrIE2UJJqc67IR15gtZvM6uAav4y8
efPZCM//z+oMX/IPwOKXdJQ2jl7Ncie70sSMp/UWh9HU9dRo+UpSvCstapSr
K9DEkE32UGzYPsNr2lW+hvDUSqvJX8G7lsWAr9K/Ps1dYUKqqfdEYKMiXYPj
EhoyPxvVc6MpfS83EpBW7r+6UPm3VKeSZ0lrBZnTBnrw4X1V6++6XFo20VOs
2Ac5+QcMUsEgrjlvyDaenS6GhBscCJfMGUDEW08+Jw5cXirZ4cRWRw7SAuce
pW8TTcpvCWDla7UOb/getS2ky8QDfKXu+Pu2Vw8gk7E/I5UlvzLWt5lvp2Ej
dZ33lfZXSV+VQnks0bafyv/DnAyCVvbNNPj4w4PnysE1F/U7i1xAcKCQgkVF
pWemWbRN3/a2nYgBg7Nxlfxukznp5rNCFQRvOIedkKPbJLwopb4b5p9zn6Yx
SLsIRfXfMO2cSBfHgKGboJgR/Z94tGb6fDRPj1JLf5vAQgSEvEmpiXGFw+t3
ABUGO7no8xrHKva6MNFIVgTF6KiFNwCjGb7tcCzunXBvdmhH/5jYaXDfJ9qj
rC0rJ9cNWNihOrALRzmho9vuokLJeVHlCplyH/UwM1lLzFtrZogkgNZGszNe
t/Q+OXwiwTbEvXTjzXjKt5gD93sXdTfeoNy4Fv0pUMa9W2NKVJUx8Pb2apcN
76q5HfGR/IbuwStu0wSrDI3QnUK2ibiwPRuW89WVSN0IleodNgo2dO0G3NF3
95yWfdNLjKUoU+qWfc/F6kNO0+GyW5PqNMo52koHm/mVPKq9EMiMuiMAE/DR
ADD/QyKTmJZEOCRaIBiiMN3qj4Q7XiOrodlcpINZmgpAr0/gW4b387wypwpr
G0Rs45jxWvHsSwjynfWmtjEj2YDHm5XuX4K3WY7iYvf9PfjsW68ylof7TU90
/DlBfc9pEeMFCSay86HatEJ4XKcY/nszzcLKr3PhcwogIC+6G+GScbf9FWrL
tcC6yXMTS9GkYScRKQoyLQGESi0xkNbaoJVD/ppU+whv6yPFqp6GKHD+yZrq
V5vXEnKt8pq7oTEG0GZo8LxPLSZRFXojjIi0ZAi+hkxYRCavI6iiwRBuIgRT
qEBuRZ9zu5Fki3ZBmTFAjfJbUQ8RoIETT/iujrMWSYIX49SDZah2zPvJHa0N
jZXW58+elSqW29CxP8zXj+uZjuS2+mVbG/haiziSCA/7uj19utmQnHKfXtas
sMljXE/JzSu8H8Y/zTkjBrFSJhNlQpfOU1uQ4St4ppcSeb5bU8CNe9k7kted
Xf4i+as+zMTwnQXexFTYR8ESuR4DuFVoB3FTNx+moYhBkUI+tYq4vmtW0vtg
vUIyq9HroMxDXZig/2YMsxr0BzZ3fZEkVM4OB93Yi7qak0UD8h4JcM9u2tBx
nbp7V2msK7/0T5Ssb3fLiMjgE6uqm4Dbu90kE8vwQmbeVctzXKVLj6knbHyD
PB0BGJCeSIjjubgLDduDu/RGjpxeW/pJOGLyTVZWtnoaNep7kf4HbZ7Nelzf
GDCI7pFKYg9C3+0v2zduc5CcUxLOt+4CFElsllCmQoMXlo3z5ykcMO0u8O1r
KAY+J2g5Q7nEM7YeenY5PDDgA/gCIFSCwL2MfOQEpvBE9cuOTCU3iVagdhqQ
WoTrIa1CBFNT8n0SXGtCkC6E4mtd2LMjxzQzP7F8vn1rdgd/58SrNKbkd/9J
qwsyi0QXXignR8Dnnpz6IGH4CRkmzI7ob56FscRLtNEATTY//m3DwEb79MYg
lk56r9JvAMh7kT7uecNkLNtHeYSFemFzspwSC3MPf+1xPlvQFEuesaos5LTm
NIeLcltXIP3O8KLNMa++RK1H383W5NuOmNcp3qfgMInVuZhZCyviPHP96E2R
QjOrGuyhqtlX4AX4DZ2Qr4cp+4DKez5o5AHgcom8HSzMpoLV1dxmf0/9Ro55
XrBGBI2peTdUokmPFSKvoyErA3fZ28VejUpAfx+e8zQjeDyED9cuHgpvwNEr
ewj1ZfGDvi8lncnuSLEnAhd0pndfSM1Lhlv11zr7ABRH/QejNXhm2OCrTDC3
cLC+Vh4Cl/TBdiq9w8FhkJS89l0BOo7oyVaMmFHfeMc/k31zR7p4HnY1+qN4
GyEpP4kEiE+7mXDPRBPZ+dlb5QN0HlbCFM089i4c6bxoQhxK/Jzsfx+CIWWg
rp8u29i4daPUGNSm5wX4DDxADTTXVEOOkop2AGA6DyMAaM69s54+RFCSMYJs
vllRGFgN7iPx3dE0wD8LMXrLGcMiZeP5kbIB4Fs54V9w+tYpDnmhrZg/f+FA
eV7Hg56w/dMPR1i7jekc4U1sRuZu1TnzpmFLZee0OzkwclkIBwIWBrhwLCP8
Tee137J3PGSndpFoe4eZW6oAygD5kIOMk417ZSPC1VPKbklAg+l2e+ZKUQPP
XeuGkIp0pSPhT6zCrqWqG0PRIfyW/+IwXO4ph9dZWIjc6hNH+JXhkFwcoV5k
OMvwynwyWdpXJv4TUtJiyPunRP5SmlT3ikmzGtcoyy6iYIkL8qYuvsK6eFIj
xfeNhEbZJ51YbsOyNLswMUQK1HbPnCFinbuju4Q8iifo+XasK+YsuQ1KoDY+
WDShk1ovZNiAjyaH/071uKWRww4oQdJcfVEz32JY2jmnzEitEOF1Fhw3Kuvv
lbsPVv1L1Ad8Sv1HiO0q0s4PiBrOlr8wG9KOlThUPsGEHRs1UP+MV9A6vPyN
87HQH0EDKO3MT1DCssH6MRwmMYBvVTt+iJh4x31nKVu+tr+d3m5jsRqIioSa
5B+xzohUe2PLjIlNtMZqZt4AC3/ellQlTnctiFzY5JQb7oZG7TjuC3TRfOCZ
p0EU0SVlG9F6TKFV9H/IoQvYcIti4/GMiUy7eVUl1OiNqbLzAm8Jhaq7QNCL
sgWx9ygtoQRRz4ZJFO7EgYfWtvynhJJF2uzJKRaeCAGlhdd8vBsgENWwM8Xf
iQG7wMJH7QB1tgW2seYtMZNBn7Qdjj4jr+wWTfWUZpDNzNg4LCXa/pOqF5fm
IrcQZxZa+VUrrLewD3npmmElOQJ2fMwBKI7i0kTm8XEDdU+nZ9tWecwUcU1h
/YAuENzHXzjSM7tcf99/TzEackAYYkjmSgNwtEVnBV6qpsJuTiXSlUP6vHpD
3yUUv6jnk153dNcuXmtvJTYapz/tItdrn0CSKyhmbaptY13hbzZrVrrivI/O
RhxgdgprpAMtRRrvTtvpCSpOnxoCQQ7xUdXDU8Otvu96HunQxZ6NpcQ23dWm
WOq+scvkB/qZT4N+7x6H5ia9lTO9J3nWZLG247aBwkSSO1GFabFfZ210HPAl
WE3ULTSCZbnm0iZMDJ4VuCaq1nyoZKmxQRoTeIAjnVRxpk1lEQ/y+AOAhYm6
29USFQxEm9EtHYSDsCbL0LW3q+stUfx3uHK8A0RV2/a5bLa4hOYPwTwgUHvk
Msox7yep9qxfl+IZEJI+930bh7+B12UFRhdUuDCpkNiDDlQgDA7X8HT+9otF
d03GP5eJRf8sNxzdfXFyBWeBoIVCZcnQn5jRUrjVIfYEvc7xsuyfkWXyeQ68
2tb6eTA21k0gdgo75h5ZIe8UODbJjLU3c3CM+Lryg87MRa3uW4Yb9gWYN2+T
jo6ZT0ecGCSUBpiQ6J7M7zmf+CCM/6UKmx7Wawf1Z1I3ATPLEN8Pc8LGm9LT
Nr1pZkgmZnlDEGQ4r/h6ijAeTpzMfPwaSx5etcTbA0qvtISHVDuD7H3wU4h0
+S0vFQIGwY36pTZinpWdzhVvTwqgAl2wsBAek0B6HaeOitEENycyVeIOFNj4
/M/FW69EsOaZ+Amb4++7AmnqhVNCDrhv6xkLISCkZtXAo1R/7bozLukohGaU
dAmRU5mkbjbztPnX+Atw7phew0CJyoPDm+rmy5nJcD4rrhoes/yyHPSGF5qH
OZYGa1Oq6YeJmuNjdWBKbeQtHybhRqDkN5AmKVACamqAykwhNx2cLbqskzqZ
NuOzL5aiNF0aBTR0MLB15o4E3aDhNr1SdXeWt5XJ62AMLr1vwVvbF0TrO5SW
x5h+vaZkxO9hAAbJBMd9mj/u7PfwBqSkEKeYonWgg2w6RKy5yWRPkiByTHVx
qtyWSVwrRaNthf/8+W1qKLTQG++sKfGQNAoOuB2/JNNnDZUnNro2OhhgS07D
maCR1Y0BPQo9kBBlY814uFRKQ7AUu966C7ucLCCsZQcH82ZoalEDQosSRrkl
lTddDBACMLWX4suYwM67G+84PNwKC3bTkFD6lBAmKWRsaapUJknzTuEqH5jP
ZSHJWvTyK25GpFNrDFasY5lqd4pARAN7xvO11DhLaMgH0Dk41+xSlx5lfWC0
PFjeaTvxdi+lIWOKDkXRlAEP+FedrfhuxJ4X6zvVma2EA5CkqbsFS13N1jGu
NInA5qp8IHfSIomum7QPmENkop/Jtd3aWP16C24vLWda2EwRnfYJ5kIv7Jnh
G4sA4P0DCdCP7YGfG7YCjp0rz5x+t1NxbYOnysm0TeePN5WnwWk=

`pragma protect end_protected
