// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
JDTz/t7OmjblhiWw3KYLjar05fPR9sIu2tk51lPycry8i46cP5JK1mJYYUsb
rNw7Y2Ksd2AC+tcuSu7CP4TOg/1GEYUkPRVn2iTa37a19ybRb2S7MbPJXB77
J1+bQF+xP7FYzD6UNah2Hjwk3NywCXkUmOPHkSNRWFoRa6LZ3YrtClQgmIIf
W5uP9PtSbmf1dauSMZpah7RSXc2Z7riD6E/G/6TZRNz0tzrV43uMwbuV9XWU
bCMxmSnUZPW2esWEZV+9R2NduPE39DHCw+JW+VF2ZLSxAPiTe+AYT0BTHYdd
YbZoYTgrbzsMFKGpKFJCOnnn1pkOZMpr1rkqRdu0ow==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
WyWL2jSUANwtbm6z6s/rvcUi6mbTWxK96OSzIslJ84h3gCY/pVwgsb4ir790
WclXKYYaR8RcAlDqp2ik5FKSskDmh6AgsTpenaV3jGdb40WZb6uzuBIyg3MX
/EdnmVrc5qHS/JhbXxp647yxY2KfsPtFNspyUp0kSEn1Ivxp4Bkv4V7sDZ49
7SQwv7L1dzZWyFCZgL0xq+ploMk47n9fFfw0u4S2wwSjlbG7V/dQe6pd4m4w
tLoHbtiQ0K57xdlrECqghjeUFNhUUNg63Mq+aUT/+Gaxxj5w9LOkVD6UIaNJ
tfiYuj5pFY2qjhtq3wCMrRz+i9lOGt6JpE18sswLew==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
StOr0g17wTQSxThVwy+tmUIYJZ20LrgIAyBFVmmFgBktJXs3FthCBGY3twgX
t9Vhyr2cPHtGCbIdlO7KIfzk8ksIyK4Sb/5rqPdE3zNY/W7DGxojsFshLl3m
ITVKeo6aakGul5npkICdHtvm1UyqnCgZ9X4f7L5bYAudjBNdv++knhODBrmb
KKiqQ2jcwwZH+N4t0AUvHFoSVMRh8W+4TULPQ1H2i3Q/abMmxovHUraPKAns
d5+0im45Z5agP18fw5QotF65zPGPw6pcvmxR8/cqiMSrnE1vQvs/keo69rsP
NTdue88nlDoIE46hmTdY7upQLqnhXa18U4AEbpvDEQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
NfwahQ/ebFA+wKMnGlKdyH9sQBwi/HfBdiR640RdtULLLxYGIQzFLg5JAKEN
ewqcG57AeoCBLmw9IWWjevBYfI4yDXR4s/Y5XwsXaM0w8glTaSh9w9rj5YQF
aYDQ8LgsyGAYUPkGqNKfWcSxCE+dkas/ZdMMDcZgKkU7BqfeEWs=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
nXOYbAWgJOifrjUEJXaxiAn1hGdvLxtQXkUy/oTKYBNxLQIF6/mXQAlnFhg9
+oPFmF9PthhntsJYXZnhDdTRsUVCwQjZaiJO7HkaQqGGpK7S5W1bgT5S/JB/
8ekqYtYdhjWMlHnmQVHAOySOUh/FP8ZU5PTUU7MvimCrzWGJ25u8bFWSl5K6
156fui+NfG81sht43n2CcB9/dM4ukv3Ex7Zh8RtFuwzj+4oGrZJsOPx6tBUV
QXtT86ToULskgC7oOqiXLK1PTEOuO8CKL2QO/HD8SzEmBsyYz/w07A+GtELD
Tb2OI1OTYPfqBJ3owwjmFDVni94Owa9+AMA5hHRHobz8uMd02KUe4g5m8W0j
/uOyU7fLG8In5vhsW0UF8zF7VLOfsSeGnN7CQFCJGQcMNWIg+nLmHOJtI8tc
7gbZC7EhBH4l5ElkHrhQB5weSfUUFMHH86vZ78XR4Nnc9zPwXlYwKC8kePXs
z3nNdINMEQ/z9g6nFTTQFohq6wgzsUYi


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
So0vCrzN5DF9micFx/bdB7/u0Y1Pd3jaad6oJO+qUDRbAA/qPl4bWKB0YEp8
pTreM7r/lQCucMeeWZ6vDPTSgTDHGBcg9QL6AngTYYqWMk7gy23yLOt0MBdb
Es1mRvd8KH+AowjSKW7SG7VgNYa3DyF+AsScoFbYzotQ/db5NG4=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
XeNrOKY3G5gfSWTCTfbPglRIKvT12mU9dPQofKEpibLFoiP4byo1THFuDpO7
02iMwZmq/o4/7dZr2+0IdiQUkYuqmhTlHkTNBP9XEpaTs6Nv6+vRJ32UlUvw
KaJEVnvE9aU8Hxt4yR8U7q3cvr2TBkWvtBILp1w1QEsZUzpCszk=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 8000)
`pragma protect data_block
8QrPhE7wY++rRYj9slm5NXpyXMae1MAr6dAnQljKIxKsUOD0HmFg2FgKg0+H
8k5qpC2zV+TnDrd+qDumMYB/o8yjBaed/r5viIaCJmun9RuKSUekpFUZxzVI
JIt4SNtlZwg8JhAsbNxLWERgWErpkq+ayeQOfLLrIwSuMDLgmWZI95iJ1PbZ
tKqnbM++CIJvZFUeoXYFwgMB0M8Gb5ZvluWobd9TsH4d7FctTcUa+7MKUoHh
MpHoUqUmKcNZke7zV2Ftp4nRqqHR/zPvAAy2NOvcUMpPX/kJbnCsSj+iHhtd
vwlwpRif9C/UkDwPuN/K7xFDDxBALt7mhJN3Id8WLwzvfKYF3eqeL+/Kx2xN
H/qi7iqeLoAL6zUkkkvU2OfRyNpSECNu2M8vhIH6q8mLXpZu9kdWb7zBBLqf
MdiD6bsYEb+0uj6E2QWuJIfxfM6GA0S98yQ4BpNwRrqdiRqyAoZEiEiOLTVY
Ao5W4YC2Smj0bnWExt1A/1lIuGTjH2TLYyp2Yq3b6jTDI4Vgjr2q+2Y/coxz
gZaYU/R2r3A34NcRqU0ei7MpB6pIg8vbdIcHX/4p1i+W4JtdRJ7j5O0/sK8S
4HTqfXALfnpSICVdVzp1JIcfANZU8tD62NQp4e92KbsBwc5vTEeRmKRqLKaZ
YuuarUxm1BuzDti3EiI3qwPfCb1ewaGr0XALxW7Q19Tav05F0IWSbH0u0C9d
klkqUV3EfdFuGYvHZJs0zKCxxVFxUCYDAFeedsqOECNleKNEU7Ut19jzkDd2
sH9XlyruYFpPwPZHSp3i1V8JuEgjHZI/43iirXe2sPtWouu56QHEfEoBwxsQ
yXzxmSWuyV0mUGT5oCKBI5Is4dxawgH2dMXnpTqxGmxUkKjABj/Kjkg2PhQd
SjY8qcKo+hT658ODCM/YOSqTRxTwPlgC9SRTsIrk3jX1I73dZu5BSjgDhKs3
LIFBhR3bAHF42a9ziea2qMwr34lZTjsQCbpSu6hdXZd9aF/G/nwCCxCxZMIH
RhXRupOVrecqlS5zYG1uj4HjJ/LSeTz5sCNXKgafTRlg6rlv0Bbkn6dUt2Pm
U0gb2S/AhqAB6itd3Xn26vWHTRfeGFJEDnC5g8a2RgN2BQTCMtRLmjqRf5su
dTsyEpaWy9eg0ybykgYQOW2SM1xNkqOKdDFWAKrJNn8sWAg49H20lpMUj9pv
euatUVeBo5KeOiJQ3JbXLeoLbqrLZdYpHbityl4g/90IDt5ReRkMExb0pkB8
peCW5a5CdBNT1T0WsbnClyJy2jqAkDFXRBeuWWpg49IbtQGGot78/TnxoZ0v
gzMVIe77yr/qNWKsv0pbhaTiADLfyTK7JR+ORtHh5LzNmokOWtuBZzdjU4kD
bm0o8UShvVB/gr+i1g+Z5cgfvm6DD2dF9gyszLIdjfT6iB86Dz/5RO2x11i/
XcqZsGWmyu2HmpLtU/4ZPD6g8SsPyWG7RxWkMsIaPIsh8M/190Ul/SssI9tB
WvLH5HuYJA/6dsXdU+fbYXwRl6fSTWRjqPnKAhI//SPNfH362qmnDLQczKGh
gOSaCp65yH6e1flZrVwrZLcic84ZSVI7g0+fo7l4qKTB8HCY07CVydgXicFD
rC0aArr4jnSTzfLZZULRQL+u3g+mZEYgaZ+9BsO6Ai2a6fhahhrpqjYY2hAI
E1juzLlZx8EwJMd66eEB1UKMyusOGg4M18QtbkjLqk1MYiDwAFYz2xG/pLBa
l0HivTmeD9AsWZ9M452LZgxTkbxyk+XlfCt93otC+j1a9PzgF8g2kYfyDV7d
yN4S9oLrvmph1K63+fniRpoNVbEfN+LiDjk9k2Oxz5C1j+rXIV+8vQThmWeh
CtdN/+ikje4t5vq01TAelObsQsIkkxq2YqDZVrA8DiUMIjLQfl7e0hjZZEHf
A1OxRz34acCk6kn8BPqu2k3mMl5rivD5xEONyhnrxv2Q8SAbCvI8/T9+Wu8U
U/pgLLCKfyuWRZZ380nPG5LjhLV8cNeFDzhaa5NnlgmyixVOuYTnWIx+gfK5
AhOD4iCfsplkqzEBC25FnLNNnadBqlMb3SWZHGFgrX7DTKMMFQ/GeD3UE2Vs
FCN+LU0al506dAb1dEl8uIqtUxEQ8XaPEfh9XreIrfwqroEf8FHH0yBDslku
Mt8HmckFaxhbXD1WbExgRXIWh1CIjxm/kymzMFLYtoZl9oFMbpGzEERlgjWF
xcXVbGdJdIquC7uAIdElrjOJ1wnRdmU2SSW+ZO2FxihwaJGQQgDLn5zF5pzt
D8ELOYvMHtwvrEU9vg0gbdpRSM4jYknzsRJ/JD22OQItVyoCrx7iATcalPPX
bXqzWLwm7HGgIs0xxGQ77OAAYscGZ2ZZh1aekenG61SN3WgWHYI+0Zs/qBLX
2LmD9u88ZmTFIWAhTAY9zIoV0ehsnsAlArhEF365ziAVclnPQ01eBeg4H84B
on2ZkcxD+/K0XLrj7D/L69HCBabyoVKRMfhh1Qe5HDvImqdhwBFclL7mXwZn
AnfhGm6YjQ9q8W3NF6y28ZaEtD/Y6HYfFuMBVjChDNgZYDaubilBvovu8AIy
ohLeg7zwn5MImTqGTyKmMBpOrxONVkbG2yRGZBAAWuNpi5IxZjkceTwX5BaM
WK+xDeWBd34rEppgEM8YmoZVBq+9Z6w3QM555TGvzLxOyiVDXWTYnh9sEDP9
Pxp1dbRynb7M3xantwC4s225OSGsGHBwloBY1vDwnWrt1aq3Uykt0JVWSn9T
d45LzvC2P7Mt1xVvZGDMypanvx0fgA3WJBMgWfaTQ4+LBeSqkPzI4qlccLuR
xWwusc7fydXULvwEbxohknYfTho3YMe3lfAuPqxfijnvKK1826SfCafZohmd
F5v1558coA2RlGhB5xBYiK4OWGx4TgpbmmuZ7+3C8UFo4upL3ODPpkTQM7aF
nl8pahQn/V8G5KcLpxcjElOiH4cdq2FC62il78dRXVG/pqSu+QxFVjVI5vQ6
BBknnE9cAb5RzgYv3Adirxf/9umATC7OJTpqJIlWv+Og7Ro/eIcAZ0OwzJbi
jFhe93ZF6klAzXMg2a0rSPe0glVghoBjjFRSnMSA0PenHKWTN1k2gmNLJ3CZ
z5oydDefjtmuA65XpcCJcHc61IP4+O625fWHy8erGG95ztMij5dmbLuehUi0
ezk8UWxItaYaYf32/v9c+hixTFf1HuQ3qIOlCoZko9FG+jhh2nqtD/oQbO4q
uewemV2bk36bmwXSbn96KZNv3U+EB4MSzwyeewjWRXQACFfCN3TP6xQ98LP+
WN5/5hehh53OLxyoSQmDP6x05qZIk+jkH2Qlqh1KZAR2F2D02OrwqQFcipcy
sYAqttFMsY8eS8r56fDbw+hZ5OAaT/iB05BzS8QJliawWly5i2zCFysGFEiV
EGBeV66zKqnwo9RqVfpmu30vVoysybK7XubPLIQLSsg2ayAkE1EKcHoLf1nd
pikLdw/obhzHuoFnVUufjrUrAKqIE4QOO+eHN8fjPZUB8GZlXD+klEMfL8qW
+1dowMqrgf7UDFuEkTAwWHdEaZl3apXFujvX3FxWGkpmoSHjIwkcs3AVJoLF
Ao0+AyOp40DfPukbMcKNJ60fsspz4nAgRfZvvplGJ+/NqFstdzw9JmbqmZHQ
8VeglR9sGfi2QGZr7XPqESHn1FzvNX/K5GJEvBg/klriPnioUk5frb8fnRQ2
bMuKFEWcFGWtHfy8DYmem7jKEz6uZiuqh5da5CaqGnBFdKlKCKWPGYpHDD5n
hinap1OcY2RHc/gDQS8K0BZuNxk8F8QeyJ+qsbUA1z2HrNQ58e2a85STuVCf
CEWUoFIQc5S1So1AOkOkojj0I8JnQ37Vp8aYvpBm2Iei723qNNDPqHKp6+Ly
ys/Ib5XeTnCs6L3ywYW2qjb1fC8kCrnAfyhPQQqUHTMPQntZxh4qi6XG4Jk7
1TlGW0JHVRGQ4Qb44Yq7DiuK5kUo5gjBTyyy28XucjxlFdfMQSP3+sPiUvXt
jYCPpopkjN4UgiohTvsCC1/fjozgja+MIr1I4cTH9kqppLqJygbhPGMtpwRf
ulr+mWl2MUJi+O4+qIkDa2icmvqtiRff9klkgZSSYyVf567d30wq5cXTbe5I
NxdNoJuHivtJRKyNxfHwc98uvvXvDrTSdd9ySkXVE+7XORHncZNf7V8SitNy
pklN/tE1V70aoSkZQtdf6xVelc5NBXPGLZ7O7af6wEUPvq6TwssP6s6DIjqc
eaeVCTQb6S4ItVnpsJGojqCz62SzbviNB4yZF8wIjdOh7jmOl4GRFma1Eatp
2dicnSaBg5dIrCHUUpBqkKTXhYTuS2hnIPBLhjZIPWqzq/xy8pde36JuQhMF
pjcOHqXldS5LARb64hnhQtU+Rbg2YcmIWb7fobu/6anGRenAck16UNGH/USJ
AQ9jjbOqc8zwjCyK5N2HhrMq2vJe4WFoEotrM8nhE3Z7unGESK/6W4BspavA
msBA9HuAW5oi6wYRQJWB7dNBDn1ROERku04wjqYWhRLHiQQz5SKcvSgmkxRo
rWTLQTIUS3HsaJjyIrXO5P+W2OvRuC8V1jY8rRBF6VrYqB4GUnyW0TNVj0MT
Kt0reVC34fGyXqj1McZ5Rt1pov7zKBWvgPMijMly1HxVG8QsNyXv8xbrbS5C
PsJzfH1pWxpDgmOBDatJxTVuh37O95UbBDIhfWsztYhdElgLh+ZzyT5fevzd
z1bhqfWPOl9sRD/KOcZW4ExF34xZoVJS7d8+L24DoRKl4+6DeSsZBJZIeTLJ
4WzQog/V2eDFx73FVEIZrkqCRAYAHrVQqzRqdyFS4tlEzXu8GhiWz467Q3lL
WvepWfwpWfXM6Bcp3AZPWWt4q4H8VVIxF8UKFtu3yUgknCsnyjB4EZIu3Mb0
tGLV5S1691R523sASwVogsCIPmiLRLdJmDffPCsDObo9o2GHpUvMCLacfp6M
pob2FzyuNsytkSM9nv941dNR7xWsgoofMZCCO3O4UAqR3QeqjmMShc8RmV37
9IHWFJoJoawggrNLXZOygDPAESobyqr3F8oj1KBWpH6PrHZfL7tG5P67Pv5h
Ln/znUkHSIWSlgVQDvEbfARjzxs2sEe/Tg8I3O9tgJfeu5wRDjX43LvQYxb1
YnVa68INfg3SP1LyQRSb25evqftdjCUEEQu6Uybq9ggpsw+B4KvgA4iZSigV
nylkc115t0wmJjG4Cb7KDEDCa3ksLgmnf6jGPq06UQhaG9aKDASHldk8FFmW
wh1ZagsBBuCftyNkyUcGbf6HIBTQRGq+SzW1cttEZLhXeUeRyn+gAzjdM3dR
bmDyZLcjys45a1BLJo5umCQVyGRgIRqzK0WO7NGwJEr8ayazVCYRrxCyAVTF
uRKGNFiHwYH/4Iwag18fZn/7PizeVl2/WwypPNtMF4FsfcLHw0FK9NAnah+s
3KbhsMiU7c7ZXW9H7hL/Od8FzX9yF1PiUoUCvD/doQHHomU1W5DfCWCznZK3
1FDZsaxCZk9lvjnsOCx31vGxfQikLJLmECIUDIc6afkQMbA0s/KIkf4FPAZ3
eY70Z4d9n3Jb97mVQyar023lJ6FKkmZTYi7v7X+84T/Xj0QCy1TPvZMSMpNk
37B0N573KTi8nt3LK+38cf9qPGrk1QYcZgKFpCUErQ8qXGevCVPmgWdLVidm
n3wP2lFohF7OsKgwQdDC8aL/7l5qiTHPtIXM3T2hmhsVqEXqGOCfk38f3H6z
YdK7dwh7qVjaTItlkVy9bPi7XkAqk5e87M48iZ2SbwAiXgqZRN1TfZV3Hrf1
F5cRXD7usL1Zq6/0zNGmc4VXw+BN+VhT29S5h4LkFgZQe4sEzaj9zBaas3cB
J7hOlRyYZBI70UmyYEZZlYlOblKFNbCQBillLytKx2RQHMAqHIYfIkCIPLyy
veH0Xd4rUWnQSCA/IvKoq4+dDWGzpXTtNnmEd94A/ARXnVR3geNdyEHiq6DR
jaRIX9tOvD/jvqfVWOOSScVFZhv5YHcivAXzQ9YLV7aYxoXlfeX8n/FaJmR2
C2/Y3SMq8wUgJcpfxd/bOeYzV/GNhcpmE1zJkcoQBseP+rrTzWYv0KoicjZZ
jzttxLWk5Y6PXFs5iOqWeLJHBHkQpo3CYUwB5TYLe0J+8e5VWc5KmNtUUqnq
gzAUf4s+l19V6XjSX0Mo78G6oQw688u0y4L5tJyWvUWSDQrZD4OLA8MZpdtz
NP1lhVU+Sj+vjcrAeAYSKzwUl3/SVkPXD0IXp2XqZIR0DQGK7dEyPbhk9kNq
lUQrcOX+U7t4UoqsAW5u0hVf0Ro4DXf2S1zXfOZ4DmcHjICcVbR3M2o3pB6U
sj2CFwDHKIgtGLuwv+SneGQF5FOwwlZIyKFzooIDY++VYPH4UrJ0tMJ+8uIp
BZsU+VFTFB3FApOUpN1cZ6y66OUkkZ/AqeaO8QPTIV4GpvIWwLIyik387MZk
jpLscS2gaG09ZzSfV/m2OyLd0r4ZzpGaVcMCz1C1NUTZ0CEJEKj2oQmtL/ep
HJLBu3zfOKTPLFX3EDS5Wb89isnqo6QBNrEe1GqmzXAd46yN5OAt26arlRVe
DkklZnkNXN0Dtw4l/wpMfv0usv6X4xBwti79JAjB3tWeUgo2VH4m4fT/5CwF
tHpKx71NMXrX/b7sgEdJlQIOf/4zy2OO/m6aTyGONK42qTjycpqV0Q35gn2F
Otz9KAEXvkZI+rbKC9EsFXeTJJKmHTjQA2DAicAgAoCkcKF/yga14NRYa/zU
djSSG56gtlw6kBPp6Y12IT43/aCMbITjCmbVG+HDbncoaFTU/a05+yl+QYEp
+FFkRFa6sx4VrGyI5UuPOlKr772CrVGZPZkQUOpg64+3DG1//XltmamKlTep
BorsutHQhVN0f2L6XioZvX+Gxv4ryvC6SAmNAUdazVSgOAomifSPGtI/NVNE
rdlYUoVDZJNc3Q01c7rIVvKD347/PWSgCgGsoB26w2XT3IU7MTH+6HZCsrQn
+zXZB45hlVrpp4Qa4dpFmu8KoB2pvX7z58cBufiYWOkxJ7Go6436ulhfqec/
/UK1qAs7Gu5d4dg8JQEcfcs/eAmOkUzscc292Q++B2lVXiGGz2ayxFQvTyQx
zH1bbvNQGnSF1RA8yHeuUSGD0sUKSfXT4zr+/opqrP/IZ28Y/GysQgXnaGrv
4OY43RZbXkrNaTxHPaI1U60E4VOp4Sh4q0CFnpwUdwjSVvuGW7n6ZdyV3WAY
V3sHWC7z/wl1BFt8mcDIMx6dJzEZ3eHCF+LTuA+A+X+w4VgNCirEpLf9RVyI
MosagBqs4JaYVkN3RIT/q+EQ3Q384at90++HQV0bveD95EGgG7SndFkntUKY
0NzeYMPYNxCQt1kBwl1tcwRiKd5r7ZN7zPHzJSWkvoKR0dKsLrl13yhvI+j3
D8ky3W12ILpqWt+1JrbSKj3Z58MhZe/68YWGWXrfieH4DoPrJhwW5ZubZAAY
+gTeWWCiE6KGfBAdzT36HP/QpKPff5emc31lk6nZxhHJnmGA15IErCoquTfk
fkc8Z46zHlq5VFtpL1PCH/Xc5BNc21U3F8zSi6XoLu4XOpr/QQyBMm2y87oC
XkAzQe3HOmruY0B+bfcvW1jBKlPriVIQG5M7WcWArSgnLHlVEvUUZoAnQXDD
C/Skd5+Xe9WMIgeruJZJRnQEZUgZajIGZLNjkbS3Y7j6YVGbNjkVSoWHYgff
QtorhzM/B+t83YYCYsb2vrsX19Fvt1LEbmVBcrPTc1rSozi71BDEZcsgRO6g
yPXgrBT3b6G3jZ9kT70yHdywIX0G7hUy2NkGoUTzObK4vHt3o3Lae7ecDapq
dLHAZpPUm9eaFERrQZIvVqsVdxzctTGuY/kRf3H/DCYZxjh4sG9mMKpjpMMC
xnyPfG9b6vzg6OFI5kowanYOcSrHNiCTD2dNZcZ+9yo6GwNNw1OzbmbTxj9e
meeth/oD6HGg0d1LEk5uTvKa8RziIvyu1w7888PJPAdzY7x/EE1sFNBeRDoq
HXwEzeFkl11cedHRxpnTMBr9sykCj20ua0+tbdyQdT9rQ1b6BxyomJzau84w
DsvZ4DKSRalB3L66nwuSMl1H4VYpvUXfGqvlyBdyfHZs2lrmEy/A8xrAR3eT
77YYE8j7SXtK8slcP3bgOlkm4vFcgsfuko2kaik2ZqCOiqufaQOyJt7lu159
73XCJrc5FMgb9pqMOWc4fHP6kIOSdgff//fU6Oeuraof/6I423BptiCLUIuk
dWpZvE7pqPOQyWjgbXaHyxKVxPwuNpWYLcbq5BsmbWz7eRQ3WRhao+o/y9h5
r8TAFCtk9iFZwxl2PsvuAtoiXPgpT5HnU2qLZZ6Vj9l7VhucVHPlec+jZjnp
fQRMERHg0CzCaDdQVnq9Wby21Pg3Ags6gR3gvhrlXf1BX2cR/yCuQ1C8Lc7A
BgiHz2g8QXtorwPIUk/ZPb/Apvd6ri+uNXiaqGuB0h+WkKneL2q7zN0DqfCQ
EkHMyBZcvfW6MMyZ2AcMqHycUFBP6hUaQqA5tOrYRiFOVKIXFoYx817o9Wyx
ZV9bdzb3zjbEfH08AvPIV5IYcv09h8PUS7JH7QVuspYkk7C6CTjJiINzGW72
L+crv1lWz8nc0dHdhgaR//qLuqFDMn5KEKnrscUTdxbPL/nHqBgPbuYMhPs4
Gr0H6NujLS0+6LAGSi+T2p7kqXZvLmRoEiad7bFJa/QohAGB93SoXpy6aH4A
2ZBntkQ9jZMDsUQCc5csCduwGm+tSY5QQ9UMJSQtkkpLOHLKIYoiC/0qb/Ck
/zNIqmLCYFhEl63bxUoXU98RcLS9mEbeLHfdOn79I4IOnFGQjozjDhfEx8A7
TkaKNWGk4zXOgEWGobcVvJPLZ27mXPCuCTx+Iv77hLgFiGoPT9XG10tcaDGF
NaL/THn4ErTlXMx2+6xR9rGf3lp8USBCIhF3YFmAVnTViYE5e672qmOCxX8N
DWZwK1e7uVYvGqeLcawSPgZdwEOCKus3bF1e+z5/KgyZbdKZfZ4VWLHyuiiW
offFBHu8H2CXKTTr0CU/XGpOjGn0h1gklZJ3cE+33b2paComGhvaDU5uRjpR
Gnc1gHlk2PvEpzVqsMntv7upD/RYcaMpmlHP/4ObcbY1lnjXQ3TvbuDZZhCK
TtWBEZSWioo3cttZdCUYjX413NnF4IFmsUwtllUjAmTrzbOVG8WF2UqET0g+
K/2UV31xMct3ehbhi9kJTxXy/yzDCMaznwfDiI5ziaZro7RU/C5rav08n9bo
Zy7tYsWFguWrrrWBY1p8XlYz3tvqCUcy6AOA2LTOmXHaDTYuJ+HBKHNrE1yZ
TyR4Y8/S9ozl/ztcgWZkDmpxv2GY+6aRTxlKV8ewPUu+3mHDXWwU+J34RrlA
eHG1pA69sCLU0+fAT3b4xa0xRHT5gJ5hO3lnqbMx4E8jOMAUZa4Rk9Psq8lJ
k/mEnFKxb70povnjSbotNhdbJGkUjmr90MQErs4O00/i/72YjogO1y+cjcoY
DPabGu7amIPsRNWnmZYhXRwm+Pzroz0A6DN2vcvLunyv4zgRp40RfVpkJ4CQ
+mUJZIH7GMCi36Kl7P6XRj/AQhPc94b26Y2MtqStgMfTrhdR2iVt6yIU21JV
ZyNhB/QqlaP9krIRM0Fva3cmUuxac3m76C+jFZ0dd0prxiISiKSm3VHXFjzr
f1iwOFB5UgsmiLjWt+PEjJPHXBaIURNQx4Kx/zNeW3VDLWzUdV1TRz6AOonY
yqYNKs+qNCqTb0sQmfsHUQSe/gvQJ5RU4+S1UhoMMN8+eoK7JubMgmF5+ohe
z651/FIV2vQ81rwdy7ORzGkw1ODkblWqw+MKZMLDNeV087LE1LMSZwpSoF4w
VCqnHoLV1keqjSo7IdBP71I2FKZLjlSkQgbxGeXa3YJ1uga2F42Gpipd4ogf
cwQsdhSUn1ER43Zq4A5oeb1EjlAmQv1gsSCkVW8eAcQ+AK5w/2VED4QRigv5
ef9MBKkDXMKmIPJyX3bTZX7dYShsivgtiXJRl6e1YmiBsXLshQOaWs+s4ThP
KKZXv8eALgAVX8MBEZHu2uGdkSRnkRAR442YNRjD1s5yauJjXNzZ+sf0Z07d
fMTI9Obb149wGyOQOY1aImQ3LzcUCoQvLceq5QlOTvtdQnwcjs0qC+ukw0Gb
BvaTllK8Wv1XqSK/OGlem64R7npP9OUbbSXVC4bZrvVG+q6Vtz/tlrUSaxa/
cESqqjVmRMl3nxku7FztwmDenHHZDptDHtcqFCr5dIXBi2b+5VloH7APARwW
3L00xdIDh5FV2AshJe38it9Zl0zQzp/4MhlSUsG6UQ088xIxEOTuObX5auPa
k+OrHn5DW3ujrMAs7x9CkdNl6Wa9JlloS2eKJhgt86MDwIdB8nlQn0UExUp8
DJuPO9yHUfpiAS3CfJXPlNPkDkB11BV8fFECHSHEcsruoVwQM+EMBWOjetAV
ee1tBGkVMUVl/TXbKpV+ec7cBFZNAKoOMzRWtj7QprUOSXDjREEna8U99cNL
xbKGdvXJcV0veQw77kztgCdrQlaLQtQXaFTcoMpjuhZ3m+suI+KL1gR6NFxv
XHDxhawpaa9lawG9HQn6Cx76x559HLq3vgoECYbi4DxjRHg=

`pragma protect end_protected
