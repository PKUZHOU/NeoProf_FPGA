// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
PUOWOzyfpnyhNndF4+C/4t/8YEjMXjCrrPOSajEkDUikkad6G/HhECS2Bw7iy0JS
ofySaqc/Lf7zK8hjYQBvH1+GpNCfy6EDoY3cvIF9fMv2SyzsO9WrnSSTrV0HTuLp
IBfYzmLEuTFMX5YKp8BUg3ZS4WxGhXUM5Drh2ab8O/HQ5+4F1UwCWQ==
//pragma protect end_key_block
//pragma protect digest_block
EvR8l+q4z6nF/QphowWjyL6HOkM=
//pragma protect end_digest_block
//pragma protect data_block
x0OvNMSc1LekYMcWfFg8AA5lxH6D8qwt79wlb1yNMeJppL6xIp2xoaJEzbxN0sP+
0u+KsihhWqJpb5WQrGg+ACY57lgIQx5WYLOz7sbEiKQhsD0esJzGIA16ufgmJNUT
Br5dHTqwD9rMZ67scoC/sCn5nZ/rQ9835j7Q0XROxtxmGzGdy6FORDTCnq9+hqQE
PjRaWEef8aYisQ+gUXfAnFWzZsqpvoov0gO8ZBsfXMTl57LvvEAJh8MBXicYuvZv
Bg+1yzgobXiDOt4g0/25GnHf914Fv8zVXvYF+ozzXY8BzluXtQeKtRSf9cfSww8Q
ULU6O9IoNBx51dCPxWbERVHxzugGr/zDmmO7HL88Gkle8ZTO9MY5V9g3K5bG6w7H
Fl3h5ooDdr0Bsc2BLkRDX2P6aCrKOy1YY7LPD4DIiF21Ug/nZHr55VLE6lAEZUOt
a8RTLcLN0nCJgVF6b4YnQDnknlj78eL7S2aVEdO5fai4wAF8Q9Jgn3JlbRoIkXpv
6vZ1drv1sN8eOt/VAVPL4BYRDWiGlhc4q2wLxRAYtGmecR2/2KgFeXE5vwtKMrxE
/YY+L5OzLX2oinOgGWR/cX37h4TcNphXwQvSNilSsuedIrkeDgzhYQesYQtT5OeS
Q47WFq4IuQKNjtzIF1TUzTAZ5UsPPxr3RkixZlSuTXzmuxWn/Nsf2xNfX7sYr21Q
NFsPscjjtzuGGYMZGrtmktwCfaKdKM9Hnco6sQcc3dMrxJmj9ZTjmdoGU4iaLzdi
hG709SIoPWQ846WphwufKAd/qMJglzEpPtq/kEMZwaTEmZh0YxIHE2b0iHVcwr/Y
8uN6OxrM0RqIMrnLvTnrWuP5lc93R5evbu/ssjj2KIxJFxFsyvzVbDPJyWmTGqpn
YbyFWDknFzMJr+2FvvfNtyRUgnzpH7ibdTaFhRfEGa7KwPNM8gMZejHon3q+qgMQ
dQCRf9QotYtPXP15vF1k8y+/JeN3PMZRlg3Way/TZCVZWZ0cUP2oEmeezS9t4LJq
aeubLFtYaldz6Ftsy/M7zEjPq9rhTVrDrGHeF1ivnOeJB1j9kH//zmMqw4wV+QRO
+q7khbWWAXypoJNGdycqfAJv+zeZCD4AsczvnxaZe0ajglvKzMrhodWY/FgiuQXX
54fqXAxis0ZKGEZwGDtXGa5aABoLq9h4o0C2/a0ERfGds2IIJioFbEVYWmKBEYyT
sfU9nmLkIe5JcAs22Q+YgexrwlgFAMIsx1xPKWK2ZklWMvoLmxFcxh3QYUcTabnq
fw9btkpXs1cAW8+YdztX07MfJKw651745t14C55lyXp/a2RXueaMxF2iQH1Vvq8C
aJHuTDpOGOw+4WLCbtEM9VTd5qRNT/LPCdjB5+SPz85gxBnVybeXCkChJ8eOD7t9
apoJPxlq0PgQx/jWJlMtT5CCnjjyxxRRwmH/dreSj190Tog8b5gqYTluJkLIpFbW
Qbg3xoO6JqwftLa5rAngLfDiHGoT19CJf+ZyZaqzU05IIBhmFwhgYOf5oDCYBdfU
TG/7eqcTSKROJOt2J8dhxs5EIsHpc8LMMs4oVSuuk1/MjCwUGe1ZGY3Zx5g1Ziw5
d0livveo3s5pAJUQiYcDYgb0JV12L3DF5SUxmZ9i3OeXi4gr9f8KjpL0yC/Orqbw
PC3mkE4Jxu1qVvwHM8hikDKByCtU01BYeZM8gBXrPyFwE159RrUd67/wurCYp+mi
5GLglLnRBVmZxCw/j1cJaxPeu3kMmz91Gj4OmiZBbiaBvbl0r6Q9RisDCGHIaTmt
5+5TD1de4WkErmMzKwSPJBdqiP8nYKb4CZghWPDgNpaJRgTp2XWgWcwMbX9JBwBW
lw+/YTIL1RWMtnhpPr6rZRWbAJCuNMp41nvKlrKRpSzi2XNwulppgTXZ6vg38x7J
XQ3EFWWodMmO8AWAWsZSQq5FOaubFvJZwGJgouTK+gGc0Cry5hvz9OK26s6imTUP
mL+55/KAe39z43BApatZlPUUNSL8JtxO2Y/X8D3qw4OBSLfAMMwhSswf2+dcD/pK
DiPJAMHTb9l8ccpyKq3B4eBTTw7zy3S8SOPZH0uzas7PDuVo7d1WCa6qW8J4MnFT
2tUXqrWV0G4iFLFBKHolol5CkDUJrvWh2PVIjBANZzwKDlQ/UzTria0KaWdtLhYU
J4jf6FIOGNSbCCPaAHHYCLzueh2fRajO2ABaktfL22PT6bn/ZjVOkr2X+AyWJ2cR
6O1hHqa64690TELwpJ6VLgwMt64dw8vvBL4SmyGOuJsQCfym2xy8lKuL5e0pWEyd
+NCmyRa3AEJjcsKlcyO2M/PShq/m6aDp/4ccnmhoQnNALVuIRLyDs2aaL82+0vGc
vOYgWhiDEKR72zcUMT6Cshv6x5Gue8ggUzY2W9IWECcuY0VaQLuDf74025F+lnRp
R3hsPp1hLwRWRrHpq7PtcJH6SGxiZvHnMNYN/ISYCQ7pkBZwPZEVDpyX/JG88ViK
IbsFHI37ubS3did8XCWGaQLi7GsKbhDiw/w7aeZqaKIWwiuKhSpCI9eD3Wd7XieJ
B1Hmf2jfP/fesQV+ySzkzQgwi0LVGqR+rxioG1Dldv3LOay/s1XfD7iEyrixL5Ev
kSr+KJFV4xKu+rUxJAsnzhMeX+piVRi+oo1VCMcbtfcvQ0AFmQnod1ywDA0Lms9R
osPExZ+J1/0LjuiGlWMEtLh13tFTYTUIob6rYaZxKLnLqQSxcfy6J8zcfkvszfKu
xan3e768yoK9a4kdEQ15gvMBYj4PXrZsOkaahLu/sRBUSLRIS5vev1oXyi78IFRb
6KTGn2R+wJqlaXenDsY4aP+Mv3oQHZWGMIlVUYD31GaB2MP8B0x801NL8Dkdq90Q
nFhu8m5avQ5eJwnEaxhcG/KZfzvCBfwxQxExhsNAczw0MDSMW5aF3fPFdGH6KCz4
kVBQMaz+GCfdvQo5Rh8M4YWuV9TptqxlGur3BIDj1HJyXZZKf9FkWVy1SsKoHSNl
FlZ2vnKwv7XE9WFPq4ZU4iTphYx2giQ09zAa7hFtlpLqIGksTLdxl0/mPo7LLzZX
G3wp8/0fU0BtfGQrSpA8FpQKryCtwDbMIHtp/Kh1UrZEmOxH4+Q+bZGa3W3yx1q4
UfiIWFMoKd/jsUn3aShdh6AveRKFWQV/PYfGtA4+6v3+pCmabPNV3v/d9LJKc1IP
//TO3pvSpbhbMVjjQewqYcLj5nvKgSVxj5BIwCmTeXqUtgPU0cbvDTDwXNKvaO6N
NK9UOgjtEaRQUbOWwkFjEVvWcguvBf3VgeRs8v3zSKYkoDuleQ0qW/zUHMT7ADBM
3q/Gkbhv9u3Y1GJSJ9gUQwviZrDbQY1rrSPxxGvPuMh8Zjm1oLuG7DDrWAD7+JrH
UZ47McxwaCtVnUXqQoSHr2n0YNlieCAJO8QJuuknBwAtDa0OGmrB3PltlFxGGVWZ
4NzLNpsDfBB8Xyk4W0GAMbpOhEC7Ggr3KH0zKDrPDlRVoYRRqJW1kxKx7s/Hjf/7
O5AWKlbDOBVv9BXkyEgqHPDuhSWTNujr6BAo8Bxt+8TM0bcLadmLwuy8BUVUyjS1
hGJPh8hWJBYnCS+iBV0kBpGH/ubwgeQiFrAV0tAu91BHPFeWJBzoQf/MKN0UuWDF
c5NBVLw8QLUBQa3b4ieSdWd+r+Su5k+RVYOxhL5gCGybcej4OWstn1gPqiZKfYB2
KeaZhCr25mFO+U9kkvU44k2EPR4vQ2zqkAp72OVsgSE0VgcHozmU6WfjAbSDIEFG
8bd2PtlY06rMydb+Y19DWL/Gv1wx7ijxz9SQwD5i1j6F4GVBaC8oiFsibc9RDAdg
vqH0Yn3b07Sm8N2/UV8aSfnrUZzUZ6gzcsSGPTYfNKiTTyFV/p57WiIgTR3pSc/f
QZsiPu+GAMwEe3FEVQ/tIxNpP4TcTFQ+OO2EdGWdaX/AuO1EfYUVg1IOWQjv/l+D
buuiPZ2rhoqcxvU7lXcZdJGt/YFrW/wfE8KXpnqm1eg5N3JbaA9ZDDAFF4CSR5dC
eNtLZBEqH9YdcoQgXZlKErvBk+3Ou9z+VFhQW+p7JAf8kdgi/NZry7I2JC0uF7xc
YH21T3LsbXygcGoqPH1ILrKfs8IVVqIWMUjeXjjhbLh6RSzISwA4koDSYFOzD+4F
jWoU1foZZn54ra6FQnI3ntps6w20CCu+KGX2icBcfWIMBwqQPS2bx8Tazg4WOUAA
BZBFYV8weClm19FpmZVcZEx/ytQWcd1Mf3AirKA4Zn77MEbRXHJOdgsNkDBexO4s
Mj1ZKSZXSZCVvLX11hR2bVauN59zcCXQe8gHpTKagHOjLJSTxuyOZdPjaK62718p
DnEPE+fRE2cf5tFAr0V3SLwUG0Omr9IhTZRH0UzYBMoNicFaAXNhqXc8UkQd7qlk
Ja25ayOL1byyxZITcnDIinFKs5dsVLWFZgAcVkGyMykE6+tCzkwOJ62aK1JbI7fa
FfACcFpNHF5PkF45s+s4wJLPVxS1eb8ONKAh19lgUiGaglVBq7X7N62KJ2q+3She
Q/Ij2x26ECb2a2Q76QrnIKSrbk6N3m2N2M9HcJSJkXea/r5mN6gXNbuCodhOAj46
zJ3mIJTyWd9fJXjYuYOLdPCel9E0N0jS0WVPxu0LMS3hRZppoGduiUW4TyjSPtxR
lfU0KDanQTbh0sIvyheei0RTPlTY9rNnt7UhCkwrO4jA+Od/lX9w13oHYc5mmclq
+1qFJ4WyKJi+UiVZxtKBMroAiNZ5YQzxSggWNnOXvK/edn5/zkOW9CchsDeb+gmr
7qk9uqPsZ+8bu2k9OT43ZjYhjw7yz9K2l6dMe8VfgeFB5YPgbS+h9LxJYO7l5djM
dbmjWLvN/5hegjY/gYFhHQqRyzhZKmNEE9Cv3e4LnyFaDIAQoyx28jiiA+zpWJkc
4ib5Bt22doVmBPMP8JBDYLXMEKUoXwNzLfK83U67loD380EbCuxzA2FBJkL2CiTS
fZGOK9Zij4iQomJc+CFJuYbdq719g2UXVDF50BNIWbDBSELl28kbl92BEaNH7F3h
TWsLpVITo4Zbs1uk9708mo0gXwZ3X+odXnxiwyoLDIfF9VqT4vKQkbALfko1CNnI
V3T+4YF+JPB1a003PDaWDkyf5RXUOPW277uWDXx+YvBZLTC3fZ5FKoPtPK85mm4N
lOt2vwvl4VaEi4IHur2uZir7jCnhEx35ctEiMZiyy9yIHaYx0476yAcEf2jNgzKv
SZngh9P8nUPf0MEKuSYAGby7Wm4KPjSE0IMQafqKFc0x9mIzJtdaYyHWIKnIVQO1
Ky6kKfI//qoCGmD5xJ/9gcUc+kPacUxFSUgBIYjtyC1fA+vpVfVV4IuU5oFYXcQK
RmjaV/XJbxVvlBgwvdOtJD47KDd7/OsXoiaZZCieABbraWpv94nzhyN4vXc9oLz1
kKTC8Cz8J6k8lYhWTetE8DV5VEJRHLiyTgj7s0yI5ryJ7KarWQzM6AiWHKx3Ypot
+SUezXdKgBfJ1NhlAhj/zPb0PTWIYIEniq3WELb2OVxm4s/zMpxTFm88lF6Vk1DS
SnVxm6YBPiw873dvtah4dRGr1EFP83ZLFQm8vyTEGMZYATkR7SBTP3Qjim5L+l0r
5d2lpskQ7vxl/XS1Lq6h3uhr/LrLxnwGzStp4cPZhE7xoEs/++KgwKOErzPSNpVR
+KGdgb09UH0sPKOnHWCwJ8o2nLzg7gpf0iKVhf5S/R3QqgkP3jTAt1XLvvY18ANz
+4LqB2vCD3xQlM2MkMg7vpK3aPx2FiHimTLJZYD+1ur+pSp1Nh9DDDnGRrdGPleI
XoYZPa/9hPsl9/BEUlm0iTMUNyuC3rZiaVsc9X/kiHpa5E5hc9l1oWdeTe6WW/43
Uqs6fxtgFHOFr1+3cUm2+5Urhq01KPRFyG6HgDyNtoi0Dx7THbPXnlhMo36z+qg6
oIMi8iDBjA1IgJNwXfwWpKLc8hJnvKyjPHBBOhh5rMfuE+6K9DEnFVTEf0OE4JcD
2qwd3s1o5BW6mnlfc8KHe4MpE0Bw3oopeBIhEY+2VtMKu3n50v9FsL3zgPpVtsix
fCrU820aQcIP2Vu+AVtt1KY6yY0SkqGMyhzLkAPofh5gDSSl15PzEoUpJ/olNfDO
yMUd6nVsXxglrb5qZi2H2f7SupmvgHvonjsCvNxHeF+ts6EhglmELXSUTVCY+H0q
ncI2jypaj9o4Is+b7XYEsBgn89yRZXyweLboHyMO/dRHv9JGCZiab+/Qpnpt4qPJ
WYOHI2+lPrnhUQp8vxH6DJZ3X0HvHJ/Plfy3SqGmArLyuGg5450YFDde//ExNLYl
GAIQ+0i290fSzJPAsVdmnmenXTCzmKOJilC8HZz7j8m4byeBXkhLAE0GlJVSJ6QX
7bXsX6bjhWtoSxtlO6cVNtVmYPTuvVb2o/UsZ3JYYR/gx6uWEXwRqLY0F4tSyFSg
LuT/pet9UDv9cQGMj9KV5W8irou3d7wQV7xllJV2BxnAgRhSYhUudBHumPnxYEyO
kE3f53DPuSf4D2ic5XJh9KQPy8k9NN96J4GG7NWrd5JMl/1VAbclF+vlCq+d7HjQ
cxVCIu1XMK01/HEwn1UQbf59SAujQcLW4gvDtCeJLuIkyvx/ZO88ymsiFgPvvUr9
kRAhASvBDkfRN7s3toGrGwaoK6IeZQYio0swJ2s0J7yFktjm2adoLT/V6EX0H1+4
0zlAom1bMKXHCMYfIxskh7JQbHKpzjT0RzUD2NtmQxmJPbQDy4hzCU12WnfnrY5K
+9nA7tzL+9kE4WfhHC0uu342SwyL+DF/e0EF2JCqYT0oF7zgUA5TA+2/8IjyUVXq
45gfMAmeq3rpWtFs8xHj00Kq6VLpsr1sn8BMFkGdsr2xcOwm0Znt5L6VfnbvbX6O
1m0fpKWwA2hKTxzekvPSw93fyWDH+qw6oYDVXX2zaNn0LMRxYSQF6Mw04BkkVWbb
iwFkIdYtF33MuZvwaJKfUqNp/Py92mk62L7/id9py8JrAkso58BG5m2NBKfLNGbm
D4X+dTT6/gaq3Xo3a+P24CoeaS72leOEEm/6p7fHZiTui+ivXRAMfJY9PrPLwhup
Mo1anaim38AOc+djptFsK65IMkxesOmp1G82M/h1jQueGRiGSJUSW9H6zeXmwmRC
DCbdTU0V8LsqjVh4IG8bXx9bBHzqFkuNz4+o00vCPJl46pRRllV2S/PMhnRyl/2K
Kgb9Pom49AGSHChhOOMoX3T1Zct5y2AXzDxlj4i8Agi6Hl8unep+nUp8nITKg3qs
zWG7TA7IJlUImmIi23/7521XyiKLtDhXXguP5PVkFyqi2nNJ2A8iA5AGo3PeKqT4
mBVvPSJMvShJOG+25kbCucGlS7LZQTo8hLSkqXRXnrtSJpqB14iHJ3pake2Qb5eZ
oRbxn18e0WWxae1F9BeK6cg8iC7jwY0Z2349V1dfX7Oifzqyku1Db088+jOqFHsB
O8pRZDEHRPCjVlKz+4+nHuKo9kLhDBhLg2rXboBeyx7PJBc2o/cim2MzPRg19vTo
AiU7DBQFWjXrAF5DD2/F3mpXdPaZYBUFYPRAvS4ILgiB2P5HEu83wmXJ39H07XrP
IMIoJ94xeSBR/JSMNv+2UMmLdYbPDI/0gkJQa6To+lZ18ukcSXk70dIZC+qIQC3j
HnRDBzEPwBumn8yxJbvVnIMfq+EjAzQf8lhJ+uUACSA2UUC28se9tbutj8uQkJcq
SPydaJGZiX+0mjxOddE62rrx8OlAAsIwzUIURBoLiReb/2tGeugmYC/Pxza8BVeX
r75JpJH4iD41eLQt2zT/bUa1D4m6CmZBGQO4bwEaAoJyNGxCkBPX3rE5t/oLUwli
3vkFoYpzNDI4oiyR9zfoJlyqIQO/vUKmKJYx49aZcXkKQ3q4APv1hYX7XhVw8hWo
483TQ7J9qdc+t1J1iHVZr6krPz94XNrGqvS7O6H5qES9x3LL6wARxSJjmR+3ducF
I9gra8mHu5IE6eFhRcpdm2pVadGWOsuCgJ/M6a6Z/T5Xc7KhrzZwbTOe63rSdbBL
QzVyvrfLLuAwuuQGwitBz/cvAkhyrI9HsjAzQgTsrgQYpt9hU5lmjNOHxSjPkHkY
Db4G3M2ahADcJ4te5NChOURbM331BRNmBPDKU+oqycEKJZLk9rdMWn5aiOrz9ZWe
CSVLm+t/6xmJ+jdLzIeGTsYoGz3eK9WEGcLA2/xRFJ0Bu3TEk0TI5d2YQ4MSaiCe
tV8FCRgqMGEbRH/FwWwvH5XwxWCNdHxE/1CQW9+WnjfdF0GsTgWnaoKj8Hxuf+KQ
a6l/e8Rip5obQiNbMqkQGXdPsZCLljVIqVamH5L+Vl3rhL98/+x5ROZDPXsUmpEK
ehA6cKX+sbLwIZPqYVuoWOyCdUgo2L3dl8kyA7GvHktCGSk81PBwY3g3DETndyF0
aEQ6rrU0Y+UAyxGq4qM3uqPGP8b2UqlzEkeO7SOzxxFZ5Em2yn04u7rnJVBJ/9cl
vmVRvby5vf4Mq8KFPw5aTDzNLcP8iFCo1FgsC94R4BODTf0UAgpvPXVIkMb5Rm2D
xpWtaYH4kFdqn8QV+dMF3ENBfUStBVfKmMB78H1/QDIz5E8EZn9UavTcDBCBlz6O
hsLMq8bVzAJZsBiwxHSMGVEoiorKzsxO11IcwssH8yFNe1CqKGPYQe2GcL4pRxIe
zAw8fTaAVakjFT+8BENn9q4/w9c+wPAhoaww+2YCrq/A7plzDvBfm75+RTR/Ft/s
lFga2bu/oIISepWSyU5hh/6htvkyZVEURgSHFcBweqe7COySOP2luvCP/FrYOGUX
8wjYQks0gzkcAHCUAUynWY2tAWeXKYDfb6gHyqXu5yN32dEDqhzNJ07ckBb7judI
dkgOAqRVVklvo/dgxZEXCCxNaIct9GNd6Eh2PCsos+MA5FP+ao2Bm/854yFdhL4S
Ryi5zox0NH/U7ct+rxKt3dCqNYUGiwSEf0St/LxRcqSzE8CRauFmQ1i+aMtaGaUT
q6zFZHveRlnK46dCi7DrXNG1BYDEdc5fY/yUHlVP/66JBhBOdu/aKmCIZuYYY5wn
Up8VhgJVCplyXsKTvwshVrhEXZTjQAz7MukHx9ITynGQaO0ZvdDiZsYt+FfXiVcL
EiaKoTC9/WM6mzK1bEOXa5XBZqPo3d90h0oDn0klHOrBiXPHz8Tj597KzG19PlRF
RRB0Hv2tBUfdnYZqQ3nuMnLIMYhZlh3xwYaY88RqnvITmYVdKb4DGZEsBh7CdVcr
OdEnKH33GKvnLG78oBJOUmvZOv9jllXynAoykwiZrh+VHNXoVep+eXdLhoIVYhoi
bEfB1kg3ZEHz6lIbtkxFAgt+8H52rb4VmIz1iaNTR/HjZ3Abb5pQC4REDxg2h57z
duVobmxWYNVUsEf8ZO7tZyjYCZtsk3GvC++qx5ZFUuOA14gRDXfjJARATG5bbAKV
nwzPshr2iaIQTrOC2CRz5Pl8ObSOdZO/JsIAJARTfAioQ010a6TLXtkq4QKO9FgB
yCCjcnOV34yeXEaEUje9EC7OwZ0rqCOdjvZC1KRkDUqqp97hPUeYtFx4Qc2gZaJg
fWKHcIubt+KZOXBB57HTNF08Oxm15T6CTytFDkhgD/EDhBL7G82OnFNzg/X9YTTQ
2kSOeep9pcqb2oQ6YUSaglGUThRbZ+qSYc+Wtoi/utTVo0yyF1tKWMbVhywHRlb0
fFDbV7y2vmN0qx8BBynnuDNW2SCHDw4LZFmqcphcFqFvwSiToY0oNEufvXF2LEmV
LKx/1/o1GpPKrrHUvXYWNEDGFQ27DUydNgoQ2GSZFG1k6//rs1UPabt23P6yVW7y
CHLdzJBWWIkBbBgstuEV8YZ+2b4c8qK54D5M6LCqhnOnEGYVc9LJcw+TezAGCPja
kYGtlSGKuUD2fa6YXJkd0Hnrl3H+eU8k9g6I903f8t/ruuNv9ItDXCBs8Mao6n3/
QKD5sBo7Uz2ZPaWah1Npu2YQq4axiSTZVEMTrvKhpe6C4iyYZJsWR0NckzTfnB0r
5KEW4RoT41Elj4ARh0kmbdGP5bXtk602sLY+EZvXCJ5sWy9BuGJ5vtBqIww32pAt
aNtmx9p/82bu2lWMKvwX06TwjBhBcTHAJsRonE/G7Aj0/acduytKMHqiYu9j6ryq
NS0nzTS43Ym/rJhBiWvaXCcgfj0V6NqjYPgjR1vLhLo4iQHcZSdwlzsGuQZ+f05c
hKu4CoDfRU7r/cL87Sxl+makOu/9H0swiz/Flv6oShOch722jAHYKaLWcrDxh1KL
yKWpQwcDzI8dU9Tb89de1kwQD7CiNpVHBVPAzxFJzbSwpGgv8WokhaQCRYAGKcTd
gz7oEayCWQxhy+C4eWun0bBf9qpL73a+caZkg1EdFtsAEezfX2hDQUj2wxMHTwrd
8JUzWYkias6Zn5iUEoVJSfJOmU2DYrqpOzSBQm4A1qRcX8UprLMaEqKRuc5VWtFf
soScsEJskQz70INCWO9e8CSX7Jln8crfYRTQF2nRXMJizCOtBL4uhgxsi902ox6I
ETV1eItvZMmby+zT971C2DsfZq/NhAjUpKEVQB9HTjliAEneo8iEkfiarKyWyVi/
ucvlSqirOOz4eQvs9025lZufWtM9YiOUfT5lS3fjSU3Z3m+QOnac1M+GuEN5wQCK
4qRx/3oPeEbL98LNJe7NMcJQqTOMZzDPUq12XE4/Lz8+0ibhTNjN+72zJ5AAmpar
ZyXwjdn/ZHHnRELQ0bSDCQiSx/dMwXBBqMVJ6QDglOD2LR3C1j8pq9SXfSA+fjA8
dWLROSp/9VFxuv4vU3WccA5aElDaAG9PdPb6L4G9CPAsYkkEgKV2cvpBVWzFkNpw
abPig609re3BgXLgydXHAdP9fOIns8tMzGUtpfFgp5D+ZAnaZU9GESNa5mBZfVuQ
xqySXRMFtx8QqShDyOfNIrNgI/1MPRGHmOJ9EtrzrdVIBgLUMo3S/elaKj7nQteI
bNJphNpDUPlIypZ+58OUBncv9AjkqA56Db2VFJMPA0ee/wxxlMC+OSIEZMbyaYLO
gzoBKZd3KPpuWjQ1FsUafvnNS2WA4TeeJagv1jIsurkUIrzgJyPfqTc0zC9oZsFl
+ABfH9/8Qn+KgJwLfHMGFJaq5RAh7JRl2xrtTAfV7KDUp5iCnijZkHcK1tPJ+A5s
GuyZenzc5uwWqjvAUl8dX7MSziIlr0W1O7o8pH/RBJMZajp5uoXDXcyKxqO5D2Bd
NWH1pvYrxgZssAaEkdzi+9ikXqrGn6a+7436kRp3447Eb/p/jt5QHf9wlAjHCQUT
pOWqkfr1X+8jnXsBiQ1tC4AYnOMb+V4VaRcchy7P6ds1qiQC+jCjN7YCJwHWbMUm
YD3gsC7QE0nAqE8f29Z2IV1tWd497bT654fbY5hvmABB+cciSw5Oq30CCbGiazEm
7kTfezP9a1sqkiwUGTn8XOxSX+Hxts405ic9PlqkH8FN5MTOW3Goe6fgOQKZrRMN
UVMuAEUskfLBKRKco3OAHU9780jQlGAVt4UX5tAssvnuoT37my64GZ+YAIt4TNJy
BwV4awFxsWE0gyJ1yZLblBUvp6WpfBCZkzV7MmNJ8sJw9kt7vbMjSGr42sdACWbv
M6yA/2cwvHqeeCVMLLAjD7AqAEdpdriwnoT4BuCaIO2eY8KzwHArTNVPDF0xy2gU
qWOhtOtNJCnF+u6uFwftF+yJAKS+o3cT5b9gTLTN3VjBLaiuqyiIj+deGCDJh4bB
IzcFRlkWeN5Oac9JfwzoQ2TkxYnER2o7hDN06fULRcZm5lLvDVbTOJ2wgeh6thPE
M+y+1hdvIITJ3A/T+4Pz+vUTh272vrm5U4zsVlilUcyqSUVhmHPVc8eQdm8LfE1N
Ravn+IFf3R+WFa99O1vfXcmvSonGp6XUcXfS1yQb09U3p8G2wjgdIgE8E/mZGzJ0
lrCLHi6suZm2vR+88embAaTF9VsjtivpfzIGzHr9p0ZU7O2Y3aiEme49ackrpk4s
NaLYygq/pxsMqKC6hl3LU1XPllj5vDLwQxKktn1m+WXOhxz2KrNpvhBe00H2wo/K
PYEr/kS594fghe4aFxh9XCMsXBEGD614b6razH7hdlow0H28wtPZQisMoOrjsoSb
yjx54q/CaVwyIogI+/3qwZkItcI8e9l2DasKmVBCjce/eO0n5N6LxEEVdzOi7qN7
dehLKBp6VvW0DYW4p5mV1Pb3jAQ1uAt5k4+wrN2/vfzcLgXwigTHhQOjX4uS15m0
Uco7QyzHYyMvgTP2GCbutaVklkKr7Wv/Jzq121GEx41UnbIgJINUUG8nyJWo8k2L
9IRPCSYPqckl4oVs7Cb9+EzZ4qg7aJGLFRsKO8S3j19JUXdygIJdPTx5Nw8+tUqS
M3Xo4gH9ua/0mH6tMc7CxTcU6IGWhzf3UM+7qx7/S/i4vERTBzw5EMcHBiyssftw
s4mrcyAeYrB+CqcOuw6H+mfLxqwN8c125wov1/83fSOiDqG7upMZSlwSWAOy6gDK
e025VwZwooo32h1D84sgKxQn3aaizcCdMASg2Ek7SXH1TmXrh9g8hXw4S8ebUd2q
ZoU4SVj+DaGz3Q7c/Ht0oMqSVNaBFiXY7//dAX43QC8wvNhOMmSDpZILcSY7jrT/
vnIyT4081Z8jIoLjQZbvTLFt7gMF+yxANROBI+BfUS1jDP8SyLmo05+FVPW4YJ9J
tE1pH8TLCOWWVJW317lD4ERnfnr91Xyn0nWzP98ve+vQjmvZFo/YQLcpy2cF5hoc
qgsIlYh75Rd8y7Q/q48IggeS17jYOFVAwgH16VzSNMSF/HmrBk5OsredDKhJDcgh
NhXkLXfdzchO/xJ2iUjzBJZog1dXYm2DBNGsSapAc/Cju1sIHfimlK/anlUBb0Xj
604RpkCs5Ii26d/I6BWMcmziZH1uy/egDdE3fcwuddH4xfMbK872KtYug4cOSV9Q
9Dk8cA2AaL75664jCuVAkcToB7lmK1uv9x4jBPS41gMe4MyUmyWtHBJwpnYKrli7
w/XWWfx4uWeD5AK4X//0nFIhy6xR4Ceutx+CpzFGQHFaUY1//AZgx4wEHfjb5Dxa
DWTb5T8my/pR+Wc+Sm8yKgx+xdHI4JZVgye2MYY1+Z/b668y1BC4DTi989ovahHB
+ADZg8N4K6SrOPGp0BviES08RfahHbsJWQsEgTTvNEHE8cAfMgDHU4A0DtqncVbT
x34QAP3Hf1nkHKgEbm5skQYmzjGcxoG8/ylyva3YkGUSjcS9CQ8umtq2gG32V0Mc
axqoZ9aDvmwG9InpDwDUhq77eE/axdMDNNcT8qZFSGQrMEy8SfMsGiPXWG7HPbyn
oVHtAvT3v5wYFk4ThCAgIhn3Wu26eNlCLnDHrYSOnDrc9qMwEm9QMhjOAh/he3N4
8FT6xJkUJhv0autbCBbCcjYErTn8Z/v31/ZJytbru4zZr7Lzw2+B0TnKwn80JdgP
KlFtCAkIr46mHosbMIVhq5AfTAK/VBP/f0uIjnprKmjn/OJe7JpdG4bRogjr9Jq8
qgKbNLJ2F+ILPkcYhtsRIZfUixyuC2rL9dTRymDlyv8vMSlJrzRTKCjstxU52nYr
mIrepkiDkwm0FLyaIGTLiL20exX5nCvJPB7wxoIBjSWyt5BIH05Lidp/zBsfdpO8
6ms0lfi5jUZ1A2xvT2vieEUCdi/k2NcgP+jUk0XQJmymKPpoT6H2KCGDbcl9cDya
+hNMSNNcApUNbo1iRcQS0CAM41B6q7RakjksANOaf2+Am6qA505oCgD3l0bwwKA8
gQ7/I0LG5zkAFqMjn7pEWMATXEx78Z3iXFY7DnWRHuR42WWB1nTuVTPcX+Y478Ne
X+cAJlv7pYWSj8nmmN7Ptipzxz971T7G2kSXQJj/phxFZTsPYHLo+woBnRk99tWW
+RP2XIwK5Vfr2aRTvDAgirVMKix3dVSyVu31PjwGkvlMhV9yz/oHdXWSXZ7Cp2Zk
qiYhoflOHAAmkbFSxr9I/g7stNhSquVeGxATkLcf9YdFskSRE0Vo2VzWWR7pdIX+
GidkZo5W7huzTkLBLSdqkdgk+A1rmCiCGRKWyeikz0EdT6yxPfGF0SzWdfFguVPi
aX4DmjyhYWP5oB25eY6VIUx3ffatZ6Ju4QjLf7apFKmlOiqfKGmM7m/Z4CgIHbww
SMIONSfXV5DqUVXO7iPr3cJqlg8r40Wx12lBch0tr04QTyF6qQXpxy1HUuLF5z8s
xF+g/qkOFKnRghzO5XeG8QLwv6jwRWtPjq4LmZIQjRsVV4LoeH/gRankdu0v+715
NMKJn+dBrXwQEveV6YqpaLTB9ldeim2DX8VBCiWEF/CeLy59yA5Zk0rpr+JCQGio
/5BOFhPOS+PKvcEsVkL5Qzr2txsSKQR6N43WJZZi8aBmzaEoYgaSLc6BDTLAxx3g
tSy53hRbL0niuVAFnZGiVVLMJvH7LWRPkUHsgWJ4pyR6lBJCNOANhce4DYyK9Rnj
8XXUqWfuBEE7bjw3UtAAEDGLoQMWROjvfp90S3J8FyDUu6B9veHJ8cpQSDF2EVZX
cgMlmfBZgvLIb4QwgKlVdLu7v/U6z+SoO3LIaraM3d1bCo7bybpHNMkIeNzTTvuI
jlvKQTcVDhYG1Sa7kw6EBxAbGqmqAayGc7mvNBK3imaOoVe0kgzK51r7x9tOJPLD
ZsMXBm5cqIlHvUJz7pJ+0N0QuZSoAGdTZAkAs5EutmjgRESKeQgzmOTLscZVPikg
R5cxNlWfzmw6L/Pg8MxRS95YwtLyMSXeRaVjeUbWdQhd1c0vSFW5Yc92HH81YTQZ
fuKCxesT/2tWl6I85mJ7iyVNseYxPlWju41Mu04NGLZvT4RQX275YGIE7nfsyc8g
Z1gOvg4W2Z1NUIV2gYOCMb/vs4Ej9Q555Y62i5SiSCZ12VLNP+u+fVz6sQHaq68V
nIvnzBCTYIWRer4zLQ6+taPobotKlSy1RW5ywUD30iF90BXNRSBY/CLqJs1KZ9Ch
D/9NzNMXfNqnvQ5g9pMtGAX7nnhsH8kZYnILkjiHuoSoFv84ZfzA8c9gM3PjgXTF
ewFLTbH6SRBD+TLO1JGp0Q1XK/S6V0NwV+nK9nirRdPotkjdvkGw7Bg/3XTo0nsf
lcE4av2M162mt/DwPG+tN7jRtqif85sZO5njWuqbK5Q7wZv3hCFfAGJ28uxCm6p/
Uc3yRsWUT1FSwpDiHXgWs0CzaYH0BhpVtg3VO1TvF6OcxIm1GJrsEzRJKQyG29Qq
1mD0UsXQDXmNjzOVP84lyJukkAj6ZSih+o85YnFwme3MhuD1Wt7tPrZijS2yElaj
HiahOQtCSeCM8O/C6e60hoF+FNYBBo2lCDNXTTzIoSQNHq1665zjtcZwC3pnAja7
YUBnXcExSlyrQSZKtZuS8wIWC+UCbEMFrufG1TjfdnSuRWjq+XgcY1b7HFn7k/DC
o+jKqua1vWsyt7bQ52JwvTEq69NwR7PMQjNRMjgRwQzp2da16NIq6z2Bq/ZYj2Gd
HpoOaUYK0/SmzpLKlyRlqCT+naWhBCBOIwXAEya/TnABtd8isMxDiF9jAE23nvOc
+m/h5EWgw+TCYKlJRpq2spJvcfjbkcN/t3m3uSdSHQfGMfrsG5Juj2NeLn7wOZxd
FQRKM+Se1vrwkLxdzrOhc2us0iFeRxZz3C7cfJttSw6JMCUqXsInjEir+bZgYor6
jeK7I7YMY7yNgP62/vIiKH47kWaXpEw8Wd3dxtzc/c1DocYjTwpZhTiZMPxBxtM4
lbbx5wFXPFQ0nRfMH4X2WelINjyz+pbLEeJDe/oJcc74MvVdpif3sMCU//sYYcYE
2ZVfUo5Uwwf68GqKFaNJpHsVA2Qx+IgyyIc93c6IPie2PkNGbzWlDQg4IyUIGY40
r2vjr4iUNdnt9Trpk4j1GLHEQAh+J+oJSve2remjln5K4sV3Oc3Iknzwbl4AGomS
Snr1Y/F5ugX8GttgB78IqhuLrkxKVaddNSjhww4C3LX1ar157XwO4iZxvsf24Xae
JLLC5v9Y+/hb933e9+r4cwha+h/zZ178e6Djza4kc1oYeC/4WBuIBAS0qBWOqC7p
8AN4MAkNkaNvZOqCA3IdsULPSme/3Z1aCAxY6HWnfS4ZAwQXwdnU46GsWOCO1rvQ
BlBlBM8EGZn04SgJ2LHIBFUO6a6A3HYlQUKmViCItg2qPEd/7UwgYyEPxAts36MZ
a5lDyp70erjf6G7SxHIhAQbWzdAVWkpz87f44n6gPIk+XupP/PGnsx4N+2zwXz2s
BvRa6OPPQqViSwdtbBxr5Zet7hMNQFvRDhHRVYCfKkiPQshL6SDcbkA/uc9iwPOj
AwMMBHbDPAp7qvm7Ollx69x7c3iYw9AoF0veLWcxk6HiBBIJxMRkRqPRjkVHM0s4
tKTIJDS76fWvz1EL3p6/2ks2MbNZeoDJF8Ul5e1iqvnJPdu00TmqT0ol9G/SmS7g
mnZoYywXrqgcv1PvwKhHxJ4P+zznGmdotvvMYX56Dd0qbNevBabCA9WZoOXqVZgV
oEt1JryZCfbad3ApEFq3xt8LWfmMPbSS+YepUZwaGDxFVWWi3BT6kQ9cWlwSXG3x
WZuH9580DKMete3x9sYp86r9KAAb8jz7aCWBRymn1cJ+Gza57b1LAP8NmfiwtUpG
hF9hk0TmH14OZ3Wtr/A2G+O5lZzxx+45RvgZV0rrVzO3q/CZL2NhgsrfOFohfBHk
M41jOMUg7Ln4Lz5HYYQUPdOBZpZ7y/iAowFATxy3joPStauEdig5hCechgpT5a7+
reOa0vrXtm60Ywew1hVMNeMu5DhaEb0Zo2tyio4eFzDtHVU964O5Mlvggk4xvHQY
x4wZ1um52Yo2NDw5NKeGgFQHIqroqlRiSyw/eVvspJaxDh+t1xVW8SXQ7FyO2xk7
bkoFI4MW6F8LAf2Pfogs/me8Bam27bclyFvQqN4qDfw+MLL2omG+zFOqVeCWi2Mv
y1nbz0kKYPiJSayRjLv86vaDdlwV5YU8//3gMoUXtiVBcC7zEG3/P1DwmE9bLLyU
AXedp7yZKcjBk5cm3DLTFcGsi3MlhmBWE7mvNz8sko4VCCmmrOR7th5PRCiwwQil
fYJ4BOZClI7Wi8Kyuw58MXQMjJ3In05MCJqvFzIT1uZZae6mdAxsRps381CU3In0
jCz4TUu44O16mTGJAdv/QxUf6feyF8xNN/jeEdvgj4i/ApmHMADXSUGwBuryFhLn
cNMgysQBHGkvDiVgUKT2elyuRZCDRngLnxRz4snn75UlWeRe6TCBOMwappYzR1Ow
IhPyykh9cssG+xNB/Qews1DlxOWstmaDJG99eB4gTLCx7x0KVXUbAH5omxWiZKnY
hqtApwLCq3klOT2ThJTqhObPysDExOxycCk+lZjVBpj7HCayU21bzFutA9Y0FWcR
sq+uzHOIi6yJeK4peSoCccLCFKMz2vP6nFm0Mksxc/eIoqFZjRaeTnPnpfP+6tUA
+R4aAlnOmoWSfX3rAVJ3GBIPgvY4RKmOl+LZXKJJnsSbHl3h9Y3Y+0rARIGFL3Dy
fUKXOfTInc9sDm/ODhGDhPBFVKXP1Hm5G/2Xy0ut53PUiL6D2CUCdw+V4ehrp4rX
B7LvVw4Pyx4KZ0UqLUVwBM47mTdn6HiT3NIec6HkY1pwOKxatk/OJZLlyrkkHJ33
rzd5l05AP8J/Tc2pgmeEk/VZsq614j+wn2RXgJ6iRSncwCOl95kocoQNRgOGJAjU
KiOVIO8Mw4jwl5dnuMXDpGjBRLao1WU8P9qJFxycLhD5baH8o/1KdYrrBfkv7Cw2
8gzcoTAey5rQ05p4HoEcXR68tD2OEvFbodtWOKiZuBkWzCmB2KnroRuhXif1hFqq
ue5E4GoiYOlXaNIPZGGUMWWp8PPGewEPa91hEZmUv6hyzscHyCvZ2Lsh8MRu1rHY
3Jpc+N/h4g5ycpPp92O12NoFB8c/goaArjbLpOsXG46nDJO6GrXwe4vHR8Ltiocw
26tHa1vxjlwpE9Lg5Ki2pTSQSf7YvrZh/WdCn4ZdtngPEQHKe90jiQ7W7HDKCDPs
Nic11CX4SjFcfTNQL3oD55h0A8eEXQ7BWQCaMlfA7P3+0+UITu2lk776VWVHl10A
O6PZGgn3yALiG4EeVpI00a43JYp1ZvptuzDkWsjY4sVbPjEQmNf6/zKcJtR/+yrk
KUnny2+OU7SL4gIPJucVnw3jWSloBvTQrdRSv1aTCwFUD7b1iyIeboF6ha78f6MC
0yAmSxQoHDFySWRxotpxEzbeFN766OqwdvgUVnj9NLQsaCID/janHIj+YZeDjbid
PnTmiIXogYxoEJdaRXSu8j9572oKPe3Rlfkz91B4dg6QXWF5h/B+jwY3tB51Wx6L
tfiFKZe6+JY4EugnPBMdmx5dyzn8sua9oAnQgDAEvyMj8uRBmlYvRr/SXvj636aB
rRweMh+4rAFAFB58amb3Qp2XncKWGNw1ewGPPsjiDnQHL5sw7BK64nRp2zbOr8LS
nqgT2+BzfLScjktixSPHwnH8EzXU4oN/FbneGCOeMqcuRNHaNxO0BnRuqUPnMqDP
MUQZSVKVPJ3smGQvBsCK1YRkreF8zTpRautWsqoBggAnWpAjz+NbPe15b1QEfgLr
470PTfwSA6uEbzTyPE8VdJXvrMkpt8s3nFhiubkzShEdSxbLffQ+eljeH6dVhNy4
ahD8+So3xJmzBbbUHLvcdxvQb1VkhTr/qqA2djpuidz8YiRQw2bV2ovhNMPiKKE/
F74Lxt/eUHyTTJ7ML96Vio7QCeplu8uUl0X3KW8KV7RGv1xvdBWNxIfha8VgmKHt
8WObB7iuxO4OuHBsY6azPhJkXXfYqGCqdaKtUX09FUW6Q54JH/z9kPtfN7eMMquQ
Y3FYFrnbBl5m9sou4TEVCSCM8qlfskqvDmQDoxSxJyKDSX6T5WpRaJR63TBGHfC7
O626wtuUnGji4MMic/27fZWlhHe6atDu3cxdnWELS8i3WlyVe52TpiyU8c2GeFOg
/EVSiw1IZDAZI9yCyxU+eMhzjAYK1loDDQ8B34qwppTdP5mqvoc6G5N7DRAaVvtP
kXWGtRihBS8dK4XHUZ7fgsiIOmb6A045YV0bd+cZijG6E9FO9H4E3ZlmCbUQ5nK/
mtS4Ly35IUz1jZnkvt7AAcNLUwMzQ4eaGZ8kJyIm6gkOjyx6IPJ2Y251zMLbZUKi
Y1OPRFE/O4qutgzV6rf0PjEYk8begFrBsmYwj9HHpb5Ti6Fi8xBo7qwbyrE434Mg
onZsXrptAQsyqOth+uV5nfG6g2XX6+5ADPlm5WCQdTucpFqdkwzxi/HhMs0/4VwW
uwyQFKLCLk8qvGmIucp843l5PrLNgRXvMf2I7hdfKWKo85hh91orcon5Y8OQAwI/
ljGobYadM+wZfIllL/GiAQS4ceag5Dk9RoI04mQLh2gdu2Po8xRmGkYBPmLkdU/2
vNVstsG5ObHKXWiYPH9CKAfxC1MWDiQxSW/dxoPuKPhUgty684LiqOfKQtW8980B
rFkF59VeuSnZVOxitFqbxY1s5UBp3s1Bm2/utECk1qbO1WhE5mUFHnYNMxTqSYxP
MlqjBbO4o3M8EgN+PkGjRO9z6Wu9hU5ftS33NMgHBaui9i2ZO5cDGw0H1aSLyffL
eENuILyyDVyTyz1CrO+3qh5E7CyRtb0fWAKqmMvRcB5vYAE1MrB1uCg/lLLNeEYz
R27v0+SEyu9GhtEpE4AJPPO8JoZ40A0NdxOZ5Y3/H/tgea+0R49Ux4w+XZptqN4Y
hTnH7jPB7XiNBBaLIWI+41/UCynyd4LilXwazlT9FdIaYUPMTqo0fS8b3Tdsaelh
LNCXdwgWn5BBYpttL7x7DAOiYT8RR6FL9gHWZbIx0VaYDIEEyGoLLszWfc3vbNKQ
JVT9qRGne4r5CZN45If78rquxN0B8akpDGQxob49+y2bpJnXg6qAb8RlK4NNr5nZ
0vF5GKK0Br6IIBwJEm2Bcvy5MAZ0Ogscz80ZgRbUI6ctqD6OXCkmxRQkrMLlLxHK
VotVZ47uKPm6V2PL+H/pWuOQ9kmkAd7Xo1IfcPUKDVvqYA7DhzJ70UIFbm72QN+s
7a8ZPvoDiA8bHT3U4tHuUwlRMZWaQd6zJJmK7SYEPYvdxrFNTYe2jSxFmwR8loXc
jxHQvN2EWqgpDeEu7e5RVnwyzik3mBYK+z6To6QF+Ru1ZIiN2a1dEg88IOBXNEJT
e46/kEAXrn3eBnvy7zo6sD9fvpkF6ANWW4p1W4jotBDTlhuOy+Vo6xa/IO6fVWpB
vwxissoDnT4kmBqOyhhvtcDVpENCjBnlXEJaSXQuR4cMYEWsrsIhOpTuvvmeX+jT
QNDHRtt46a9+SXtNaRPSgcgCn21bnJxaEroggYYW0Hl55jOCQB4G+lepAnz7XwVG
oNDV/SC8vvnHcr17FCaIV/FO1spMWYofl96UxkbItsQhIuVRWx3exgFY9npqmNvL
bVW0pCFT+IpKnKexQ7/B/3XRNMGTcy6ndrO3SINByWGEn40Db3mEJH9F+mXEK5GW
3T7Ex/g1v63ANBacryow38xTj1JPDhNaT40w2mU0xW/Xy0H1gdO3/tXgZ6XOIAZi
zNr4ulG32hOzHjN9xoOwSeiPp5p6zD3GEIsaKC8MMnnWGIhDbMviWaWgYFI/JC4E
ZKoeCKxQPbW7bwwYrnURICSmqdgbzIZG2+MfQSvqxUAkou9CxjmdIetDC9PYaOft
gLB7pm2pBPbMM1ULEFJ8ecb4NHvACLxqe4dh4cVEhnpkYq5AQO1xDxDgc8kjFSyb
mVEIQeZDkuupryRKCzrig6nTqb32NG8wszqSiSFapZsUaoIQqOLZThM0X3rNEbfl
TOzPMIG18++T059TzM7WcgWuXW4NnRzEQh42jgLEFim8p8PVTQVWqANkGo54f+QM
rrsA/ExcwBwNqHph/a2DlHRq2UzjYueE2NIwxU5F54fewaNLaElDqe6P292LsKKl
Ea/ctWKnZn9vm6NLGxaL0WZhVBnarRMXb3ZejWnkOUHkwyjl8u6Ds4hWO5X3VSqr
aeYbGOuA1zXruxLbiFoqNbutmpRtzBmgNvLYRiojqQjdjy7cnZ7JwH6H6nlFknMq
q4NyOcAjCTbuKfoRGeIrsXequ4iOyVKAbJIOX/urIrmVN9H5jHLEDavXWeQoIZjc
pOUfRjeIGnA8XxpQ7hn77IlDunuCjK1wnKJDwKQ6PQmdz6pNDqz1kjtu/UXAdNyh
dXn8B5dUSYrX4z6fhbQga+I3XsJqMXNdhBTdyCqDGIEpXRTQ88zHD71zNp7NgAsb
v4I9gykN5M1lKHDlZO94L0D2TMqnonqlKNX0PwUaBRruKFVgzjHO7f1V/d8BA+Q+
pFjHNXL/0FKs+DJyt7wP+k73DJsRYzjlYoVu35xDl3HuOjZZiElb8xjbu2Vok2hC
6mBLDafi17YnDYZVPrOhi7pJXR7R+U5nizKDfKgaKgCWvh4HOvxYq4eEqlslfIXy
61+KxMrw7llTD3ij+wtGlbq4pRUE/SFeeQiJxMVkecj8JzF25q+1LHn/gPOfCFfI
6TsB6GUJE0YUvAmARJwNxYyjAXUekVl5rPlgG1/Hp4SqPP898iTLJZYPBN680WEY
mNGM7lNLF8XWcfz97qPmg2Q8mCybDRnvGUAQrBsELhdSVjYUrdXsH0NMjVIvn1Aa
T/fskeqcvh2r+36PCh898AZiBDM6A9udjyIWSnDUEjI1SXTdLGxM4WU/JdTjUiT0
4o0LvyO4kuRoGwqC8y/UMNYUIJOpGp1ve8qfHzD4wN98nOCUl4Wkpil7VAZv0YWZ
dTIUX/1b/bCfkfOw+Ur/aHPsi1oRvcK+Kqv9sXm+yboQr3AsJrenvPqP8I7RKL/f
HuGixEatteSdRLkCAW7ZZWAhV/4XktY8PecfdyDJmwe9HddtFX1w97HqQYkE0uK6
oCjzAjudt6jy9ENPD20Rj51Gr1TLXjqXFErwrmXWHm58L4kt0b86HnxoGMHc8RP7
Ft1TF/NRyN+oysiJrF/kgruTU8EfO4/2/BGazf8nSIDcLFhsJF+ZP8ej0QJiI3jk
8mUxF6Qa32+JunvGQyE6QwHfY4OSLrZpkDOWYkcvA9LgoaXt6SRUlUtNZOu9okMS
JheT2cMmSmfvxDdaFXvQgSuCZ4vdlaFPnf7WSjtbPgxWa/WwYWoMrkhIUeHORyU7
nY0q+t3/8UWTfs01optsQZifWzwrzZgtiAhnMdH4ZhfxrG0Utc1/jbErzHA2VZhM
JScX/vuz2Cqxn2tZMG/hXRM4tAEXnO+NECzWn0ZF77H6ZxzC6v13THcjqDGfRHta
UW2JyHlyofRViB71SgITXdOiL6qhnmiXIp9JlJBSRrr0foCmNSJEbX6oY2GjgDL+
0amLTJAcdrvc3MSBTLnT/AJkNMgN8Lylr2Z6iCN18jH9kVcXPleyE8ue6D+Zrmjw
VxlIYG472kYJSCtYq3LWSdg37hxQpkr17xNL/F/qgJLfS4/YyPuWq3imk28NXuEE
jDkXJSBMc1Zvd5ksE5dyZm/GSozyaurI/uFM5j9raMlEd7KbkvGWexPJlpcfX2b5
rgrret0sfOFfkQFrrzD0HjFhwxTYLVzvM8ccMQicgdoXSnP9SymQMBDH1zvorZ7K
LshL0jwrCfxA+G/ivtdHYWQjgBSLjk6fenkTz+BkXe90tLtfkju3wzlG2vcwTJwN
YVi9SRAPbaupubLVg1hFau0hFs2TOCfbu9RV87XzDz8uorRxG2waD8piFGk53tIU
5F7LKaxsjHTD8F6vbyag3reyCflShuvZoJnVr1+zw7jcwk2z8cf/iD1+dpQM3mBF
PE90qXnLD8D3AaYsruVheVcF7AAWF5grkI9Gl8CRH/u1xagJB9hpqlkEno+/UieE
lU+w7sf8z7oYUaQpb0ictmEEnMC0nFCgoU7C6UEOYN0hYrosMErr10f4lFjGZ2N4
6xy0oTikkQkKwctRdGRzjFIeCm31sVYvftqpxipwnZwIA1yyHYxOZnGz155IiMTq
rhScH0HJI5ZAhju03VMABXnMEmhhCnlwvgPjKCSbVLix2gm8gIiBX9qBhOrS6oVO
H0Mu8QgaVzFeediW7aRQBx6n61N/5c1tbY0Ta70UZFBy4NP7XrqgiFJqLEPlHF0N
7uRu7/U1zm6c/jDgwOwiNwSON6g3JYwPZNI6UTiwylLzkQpVwoRuImwc7vC4O6wC
S4SJfGKAm2z/YUa/aR/7HZjczHREkqQlcyq4vD65/ut+sEhXphfIpqIDUkVExe9t
9VRVpv4cz3puKNJAGiBqm4ijS5CLJ/IL4R8YFpXTS0y7eUVDegRLn3B3EBr4J0ih
DNvCdCOIKgqWs3RQgnTAxxAQ5904CxtaN3ZPWuwUITAFIOJH4cE6lckVDyh8OuzB
O9fpRQv3+Z+DCW5bhucBt5Z0MnFvjIwz++07Cv3jMExcDAsZFjk7ZJAy/bYz1SUl
D7NoR+riBYNDiDnwqyUnZOa8nITklik8ME5uuLtSBJ+iu5p5Pa2F8fCexIB9CEHl
TtshOhLTDHNG0T85I+gBn2s7+F+YKyOpCSOT6S6zmTj7psFfBhpCe1Y27/zBPNjb
sgDMdf5+46ROY9YVa8ZsDi/Er6NK5MaIYY8x516xlfj4b8rNtr0U5VG/enk475y4
FC/vp7Qdc4+i1gv6Tu03W2K6qZvIGZfztXuSOQcEWqya2I7TcxFGqC6E/NvmJnpz
7aUqUoXbrzq02+AskOPPPFtl/SlzrF3Sv0fOA/4ZtwwiQ+sl8vBiXP2CXx+tzoR1
pUabbHAMVOemzoOJ+wQYto1zY3QKKel2k2LWPNERzBLsOxTOj51dKwhu/d3a9Rmx
8kyxaD+XEzPA5pSCeEVKbq6a73o1nJA+T0s/a0qjqNcP/Wh1QTSd+AUBU/TXZLO7
aap/XS739wM+MTr5bMlO9wfSidG6WGXhnHXuzx9M803V3BitXXKzN+49jilOKO83
Qp6tyrM0tOON4dQONeyxE64/xgMkH5WeiIw4j2P2YE846GGTlobYuhbUTj6ZG6Ru
NjBtc2cZjlMVY8c/ES+MxRjK9IiYQo0ppz4KUxwmDjZ4etryCatFBN+N39TBthZt
wjTsOiN7X84xz5Dp5B8kA8PkFBBBvgiAYJnJWQ6yyTPbiFgyuYiYE9GdVuXpg6u0
nnyqX1yACSTHTQ5BYgyBeErs0FnzqOyiHeaEkLwSBrsT80kJ9O+FDUCOaL248N9C
iLz6cUgmqxcLwY+j4pDIMDBkd9SVqS2ZrwloBYUxJWq5/K/eeHJgfK1wmPwR9LcD
xn3p778AZ1vzqIkgtkid5+i+0hf0xt2lyVIXzXbYcmkm2oOHar1/TbK4BEgWb8U8
v7+MZK59T9geUeFUArhvtco1kn9rKcp2UHOV9tqCW20NT5AXRkr/pT+kzUPJlB1a
MCewwVYUBhEewrZLS98+h53iYHEmTTz8rA9/bxhIV5HU4gl3LJvbmUN/MhggTdLF
O4+qn3AkhyCRojW4gNzJqLt50+BoOUKcGXfkdk9DOaYgZfMZ78k4JVVg4fCXrvhM
IY1ObCqxgQL7tTawSz5xIs9BA3J/aeTtFPa77k7mYVFECNA6qJAwAnjm/laZ5kBv
2hUZw/bkjE9Q575tBS51PW1uIyCa5/+j7Nf2CHJu3d1wlp6G6XpxpTQ6cbI6E+ob
iRhNqykI+hq+yKcnXxQBdhbyXMl9PNEeox6cOLAi1oG/gXZYzk1aHYXxgxjWundo
KxWGiZ13Oq8nRh/hOTFBkASOgmNk3hPeeEretgd0Cc/Pc1vJ7wmiEtlLN/Tmn9LS
wURns25iF/M+rJzK2mEUK1a4sN3XeHjYjcvJjtC4jAzcE0+ZqOqnDmZablm5Alk+
hfggyoGCkIiQAaiGvPakmUf9jn75EghHkelcnWwQGPTFu5Cxug5wfUXqKrjjuMz4
dmQ7I7gJt0RVSoUElcFDo/P1cDr5pSyiHvPmxrLniXYtmM6Aqpw77h8oC3QvlpvB
RCblsWhydk5v47UWyL3z9jnLrwFsZw4CnwxeC0l9cCXyigdkRH5d6yYEK8WGVxeG
8u8nVKbP5vSn5EEU6E4llU1vY52WHN2Ag0vo22xAqRUEsxNY5VI3ucOChwu2KhrM
LtZBpQUakJQEQvkWuCKq6TCPF1+UAcSBgF1Fs6uXauUhqQFL6mWQ6x5Exg/sxXmO
ANgMMVBaxOrIG0F2lF/CrX4aSLj9wYkzyIIjORuDi6yqbaTAO/gud79OF3T0y0Ln
0o5TGUKiZYJGL0H87Z2pZHXhAYTZqW2p9KFgV8IemdZTbqBeyJZ7RYcDIlAqk/Yj
3VjuacM7DCy3m6LP77lvp+mvDlY+CVKHDxIHsn3Q2IueWH8KiJCDkYkRxhR3+S9e
VthdPV6x6AgGnfv0pewskJaBpzqMVZ5xxp3T0UGmlnlTW2BPKtwPDBVClXKoS5Jn
daBH9v0lfYc4M0fQ69m5CeW9f6LZcqFf8EJjkhGADLxaOjic/Qlw5ncNFVBHu9AZ
MsdM9prap9wPVt2Ix4/4E7Yt1ao+QC5xk4C72Mg/zFENCbMd45Nx+a8w+3REokpb
KIy+CDm45r8p7CrHq6J5zgPbglv1tQFTNYMJqbB9dFB3FY0HLmUUSMbFkTUuYxZ4
EuArvWV7t5TcVraxVgP1XAE67oXYQ9lQSgnT6I+NQ40unEC/x/2F3U5CudUvE5ZC
UrpDUfLBMgUWNXBK3IeTieyhqki8fArHcAG2sMyKw55Wn3pDD+nT2MH0j0Cn2lI7
lSZtDQlnEz7Oi22dnYmfU67IzIPTnDYNaQAHK0Ejg08gviidy7Xs+KWUN20QVVKT
Wj/CEJijNvi/eFSBrhvCzW9ODud3cTQtf2rEEYRw45ddw6rHsKiRy2sU7WFNi25f
mVaL7IEI9+835c3w6pcjoAlNaAHyVFT+XW6yAvzXwFdBc2dj/qtARSZh03qwtdv4
cymprwnS8Mmn99cyhJhNVdClt7E3QCGGoZIUPlxveFnMqVVLgtajAeTCg8sSzAXe
YDel7MkM7TDFOswYQa+iO2rhx1XsYf/sluBw7ERNmcHpBsMOxknkosWp7qR/8P6K
DXB9hmhxjyIt2m1uvf/Fgci3u+cblWad0Wfg9YJJ30ODog8Cx/ZJ/c3q4Lpzy+tM
vOBV9XC9EUoXXmCwULImkS8jIJrdOVQUFEQHMY6zkuUouCF/7mYTTz2qeNbaxJsN
4+mLFNFfLKW7I462J9saHKUR9T4NxWpVdd7s9OUZgAcOHvdfLeXr/aI1E6tckvK3
FQSELvy2Ymc6al5nh+9LqBr7onFjIt/4k4tMn/GDqUWotS5bq86e2QXzVVtDURiG
cwl3/IhpfiulYmyD3qigUECGBHxc2TpucaV/yq0/Nq0Ol+tYuRFtBvJ0/mNLW82l
fWwEcuXR7zT6ghOq1DMUtq2DcGsunub/+iQKOs0gtZGy/wcLrwxNrPk1Lr5pZDuk
0ocjWhFPF7Vp33wAbyJHnukCCDRsKjf46M/15nfIjsZ5SlwngwtVXS7ej4qgtIJG
EvFBC9W/GgL9Ub8zbW836OqZHECaQhADZvfAJf18AgLnIhKhdrNxSByqLFM579kS
VC04EaP6KF7ljGHPs1ukujr+boYbXDweiLk4IEleov04z/QkH+3B6QZT7xfExrF4
lrI6d4eyy8EYRUryNZktD6m+aVKE3TXivJUIdHq2fJG1qEqyWFGjkZEMBPxvlJTl
/n7wBipZyDHNGNiaM0wob3hCgi6nIQlRt8leMtD8JKLqm3wnd29luS5TGPBeJcBu
rJZXnejHm+PRuJ1csJzCyoGWO6OjEfnmvO0oKBqV872sSdNIZnFH5frAYmTVsYP6
xA7UrvUHbF+8rD+idQi8FjaYuiWNZaOK2uTm9NH7y19D0Bp1vKv9fejS4X8XiRIu
jbIsK6IiVxCmGXBXL5GUOGwe81kVexHX+mHLOT5WPjG6u/PxXomsx+HneuQbiYyx
gJlGrVnq3iRisFjmBjhHFv0KG3KAVPgFTZ08erNrsGT0xpERDF5DFotXRK08mDSx
bu3m8kuGsUEd/GPZgc1y4LO7MN+bn9VvJckStCPvZ2Bc8Cj9BJffBH9LNY+BH6iQ
uxKhZg/xrC88Kt9qKDIanF3jmRa6eC8CwWz+0nmPTW7MLOjUVghdTpMw4vvD+iCj
H8Z3qy3Pr/nWeji2CxMULUP0uPeJV6eoa5lQnZqEGsFBEDt3M/n5gfxHYyShXCyF
cjvtvAuIbQ9QS/9AlcW7icJc+czfVc8e/3eU1qlOpiFhLSOGJl2SOyc9ll41kMI5
Jo414T9PQ0jpIEk2prv4uXa7zJ9tEXC1RptfJ5xwXzsCmCzCubPHrIzBrRGW3l5y
NlrGuBT/P513G7xsXyoqCYAtiTL2zvfMr2Wi0zVCE6NkIDbXl6laSnP87DNZDS5/
FJg3xr/3YJq+bF0WhMaq/7aZ0imGFmZ9vlIhkS5I4xe7wAoeYkp7FMsWy9A9q7Pk
fviu1PNFqU7GDau8rz4IvVDAjbCZjCM5n+2ly/ghw8uimEntvnjN3slKrK5rvh6b
KGJ9P08MxXhHEh4DRgeqbbV8Iq0j+AZWyWckrKzSPCpWYJUThwvQMFN/44nwcBct
wpKLLminZWHaVTVV/iiDt8W6nrIBkbTi9g6n2K72ps90Wo3XYcM6mlzJnYs9MhHd
p14zzl+k/NFCzYNz2BLR4BMltBVbq/21a8kxoV7F3NmCxrAF5tHweYXGIXUSKN0o
vfVcy+xJTNos86sILmE7EIJVyUOM3KNT4HO9NILdPVBGPN+OZd/GM2wahU5lpgpU
p0QVc3jMJpS47spjt+QivUuBzeN9UwbIDnJliJsoXvakRaw2PvQ90o0tww3cDQUk
yvgym1mYSHbkUp2CXTvMHLkPyYBfPvKQ3EGwOK2XNYm5WC3T1MSu7bTqF592+D15
NwS3TzYve37IehO0gyF4AotVHMaL5AyvZJl3V9RX6cQCLJ+W8d/Ahsgc+IykAic0
MZDfb48zdHv9UTjlhu3VEyYk/CDqLvB87Z6pipO0WZ7pYmvsfuhfPGza7o2g2AX8
suiAKW0Tzb73/YYFzV6CQC+D1lq6nUEO7f6+XuvGi7wDrp4n/aka9r7A8Q8zhKu1
djc8mt69FfiWEuRpKRokINxfli29OL6Sx1KmscCHbF9cXEGAtCaS5OqHAGeXliOt
sAUK2aZQUFCK2gs9mjKcQN4SI5tZPyCCnkbOrdhzE6q0kK0BDdy9Uiad31birRqd
en9AR13d/kOCBXkopzd7lZubIs19Qxw7J/szimAgwYIF2gPT6U14aSZd7Rzv/qSu
c4LstjevUvZBvrV0C3+SBI4d+XXu+aXydP9MUfSOj4qldITD+lXnDbJOwCg5Dacl
AUtOQwd+0nttazpk9afQUzlhKxI6DekC/1O0l+tu0WufM7txJYR9Gxszz/XH94I9
zmjkD9jwupr6rzxfyJ88gFfFVdX//rkSZ6c1AWbdLk8TXvFSuhYVPiwSQMX3KZsH
SpTQX2Cr1N9YZjd+AQTkOJMOQOAenE5Ym8Jspa+EMs4zDMnT6SX9GPTpIYjIUyyp
VJW4XjR/vKOGbNxKlhHCXSODhCredMLiFaNWzxrZCSRHCwWsth03zH69Ztfkq44R
pOnShAu8tfO3lgf6I42kwIcMY8vqxFmcHNWtY60jP78mxJEteLVuwVeP5S/+82Im
8FpSp+GMChAbbH0GffZobV4t+D/doTSys1ViMttKxMcIW78H+wE9Ad7D8zfO8pVe
/sSDIUrr/yf6CEtCPBTaWnzOSiDe8aXUoddVr29ZIs3ZgKqpn4jhnqCS9RzfRDNb
ucVkufAoI+NsBeH2jpmcM/lPs8t1GzYpSEpQg87TJodkqE0ZKH3GTMsF+woGdL9K
O0kRyZ4G49xOamIdxZlTjdsOcScNpQl41WCI7PwlOEzHsq4IcxMDYcEIHmNTvxw0
qgSw0TXb/zGZeyD6y4sabwWbayiZkJclBHAG6/PWoxGhB/kzXlReIUtzrWBJLnBr
Vzc6GUrxwcbrxqz/TbL2UISjC6rOdgKhN8QDvLl1i0r2Xp+LtDdaSOfAzMrf0v1g
X1nTPQ9tiIMwIshZez6fAenw/Oh3kUCLuvpcPP35ACxa5anllk/ZFbuKXC3emm34
DknBvH2bAoXKgTxNcVu/EcUSuHH7IBkXh/Su7hLKCMZHpjuLEtxCrpvuP8QItMyA
XqmZofOzH0HHa+2F98BvcMSPhpSG74AhcxHlrkKC61E37sEZU0m+rnoj5qFGEXzN
WhOte3IjWaQFLdQIuhN6eYz0nvEEsLQt7wQD9un10QxN+hgOJVRKYPq9j2qY1roI
3dj2WcV4NVfw8O0DHc5EHEge6tWCefHOpOl5E62kD4aZIyRwgH8X8n2QXHC77wJS
2hWk4lwWXpw44KXz07cl3OQ7ia3oyt+NWSEFTZnrWhpeCciKpbhdH9x1pW5OaWcD
QeMS/JX8qSC4f3OSAgQEChHGQN3uRNv64kZcFtG025UWhyM3vUPOCjZ3scL4CuA/
E7nz70JDlEXjoWwkOi8i/copZZenL09o4z9GFLXi9UmoIdwvVOAqnTgdMZO0FyYr
HAiFrJSHm1JCb83GHMmvTPa4IvvuAFgZ8hstzbjoKGpNjtS9z2wL6Q9aHfXIcx8x
M6WvxN1VAgs6U4pn/c7XQV3fO+z53Mh0hgclfPTKNS99o8YUzX+8BXq+j8surQB1
Z00kcD9p1N4RPXPQ+35lh9UUulvAfqQqjmlUlYV3ojVO967h3E1SfUwg34Natk/I
b86rYFmgiSMqPyWvUgtypJ3bB90rO3vUtKViHHeVTmeswpN1wZjiefWJnQ4tf3E5
c4kVP1TamluFaDzltJ79gRn9U+h6y7MF/+zQh7tuIXBgrEAT2Lh3e8nIPq9SGQKS
/NE5Fc4gsrWxhkMDlTOwVWAcudvcjvJAdkZht4WM1yq8zpBn/uzTiH0uohP7Ouv2
6OVzha80xbunVfPo5UbIas3ziyFv1O+QY2mmxN2re0G/PXunxBLBqPsqZxv5y0av
ITAe0a3O13w11QuYGUGTNsiGQXghWslfcIUWp0QRGCl3IPIgIhwrJGhkLvq6tX5U
xz3+ym4qDEqFoQbwDeYPwN6ZNRPWYewofTVVswP5FVG85JLGGamohZFpLi7/i1vy
khsuwnuFlJTOJwsTRgDjEgCVLNbjLCMFA3AfcoWZ4f3B+rCJbcQkCqF8nDFShho0
e0ZmifzbXJtiq7ThpmmEph2kphWSW9QSdfqECnrEWPNydh10kIqbTdvZ2/2ubIPP
eroPdRShG+jqsibz8l/ICpIhaenIdQbOKjCDSqaT2JT5ElECx6Pb7GmSZPQPr98R
3H9x7aRTV01oNNmFE8D2AoccjE4azaUcgf+8nXR8meYSJ4+rj2Am1ejCwQcJfas/
JVt7tscXJ5lCXM++azohWwAMcW+LsjJmV3aaqCaCqkyqcnN9wqm0Uq8gGyAYyg3U
G/g7/9yR6+U04i0Za3caEjKcNmsFOEvWkaUV2KhUoqWGBoyvspJoTTOW+4ED+VQd
g9QBx9DMPz+HrsTW9q+XvSzYgKc+LbozWn6BWkO2fEWiTWPoTSbHujv9NLd0BnwM
/5BMvsalu09dS+Qni2qeaXaN+m/Yf/Pn4PJp9uvfp27mFbDb3gI8trYqej8ORiYV
OKiQsp85EPUE4Z3hGCB/1R/1LUu7JxNQKG8Oj+RZqibTRWPQuyZqDFfclIfF5eXB
Bkrtx2YPfPbortr7xFMrzC+8/omikjSdyy7UMC6+ZJIolG1Hrht15wxwoxbTok0Q
P30pJrk6S5OuiR7h92bdu4Cjan4ycCeRBXNtmCar7iukPwtlEv5xm9+uCKdKstbx
lFXFrwL7OJeQM2xBfn3Wo7ofw+Cf39Wj0ClbjgODkURppJUtr9Vnvod0Od8ru2U1
NiF9wDf2g1PMyMYzyPQDpQ4UAkDtc3GKt/yMYzV38NdesUKrHUksZxqlKW2DPvSH
hKFcDRMhf6kXxE/bWwLLkDSF/Y372NGM8WxrP8c0S2nI/KKadCTPpnM2bUOHwFEZ
6mlt4c35aQLynOlgkJcLALBJxnGrCYiU8UaaK7QyYi7RPb8vwodlkMkzmDw2XTmD
EwDiIIAzSSU2UQL0JOaBTZVY0usJwhy4ln3AQgUEKtFgYGlkBk1UukrUm58MO0kO
yiN8LW306s4ZnJ5mNwCu3VJs29Ql7nNpp+EUNVTZ/fXOiDj9tpokMHDkVaxf47Rt
aLKUg006T58L06Yrrzq53SLKDuFok/AnP4VXi28Z1VsiudqeqCksoyBnq3lU6M2Z
wLkcFlX/M4LJgO7b62jS6yzUJg506bJGM9muWSwWH2gwKrSjytnW9AewZ7od27t4
bfA6LiUK/SAC89DLB4uincJ9LjXFjYfUn7d7F07zSBmgq1ntFpBMkwTQzp8lha8D
xSmesxqMn7H140crt2yLGAfPPNonpDlWhjYz3gV9sxh+6xNbNGVb0HmYXas5Glla
KV39AeZ1S+P9DHr0bUOR/HBTVW8UkuY+LaINTnTA0M9CkY/F9VqTA8zGuLOa48g7
VUDhQetcpYrbzYW1rH9LTGqbH7g/2/tmkHZ41pljrD84SzzYvE3G0ypkG8buEhNw
qzaVMRnVhHx9n+/c7kTdgfANiqFhpD1aO+YlWFXnmL8XW+zkxB+to44TBKM4f6+X
NWR7vD5fYmmwLoPQ2xAnMd31YzgZLdwRDFqZndgBU/m4Pr+qbBkFZULHzIbSusU5
V6g0/LCT3/rbLtMVBoAaNkCyCypqdh2RTy/4iyFg1mO/cg2fr8pHu7L1Mc4WRXBL
wg8WJfzbjQwLpoTmXZuMz9sDisQQnFlRPhr3IVwFt5N2UoXuUtIDRxWlhcEVSD7O
8OUCWQI8VpXWTuv9niQsYRqk7Ifj0X2zd96J0BkqrWvv3kACJJmmeS+yGm5gnmdJ
FQ+ZoTw9EYNHyogo8HZ/WantKaXPfsmeUkWSSD25+ZkSDpipfNLf3/ZNHgarKRzj
y2vhkCpfShBlDR5Payo2PN2fdJnAyTjXsrCSOOF5EDEa++UiqA1Ngn3qm1uCYOA6
kQOK2Cb76Os7OnAqSKwIZgBU9ymfupZAsanxZ+TOy8t5KS1XV6ggrf1p9+dhvRwf
oAr174NIFfLQZqDLIn3uFl5yBm1MzxfmLXIlXuCSPo7n1XedQN0omzPsaqJv+XIw
9TuQAWh46LCJVbzntcZnUShVFeRvOVhOpcBgWTLkqtx4w8xCqvoUk22wIolP4cv7
EZgHMVB0JP4Mv4zEdlTc0Q2Bv1jfcbZGB/+QtQ8SuN87yPYsz5CqRSfQwL0jRMu/
dGVGpQQLPQ73u0eWPY5DYzm2v/yB353YaQXsu7VO0i03H3w1DumAxxugEIs5f/t6
HpdJKwfEhHTXijetEt23bVsLo2U6t/tr/dBEINc7e8Yty3Cl5hevcvCY84WyOKhX
c9yRrlZMITbPrkwBgliRbl4sq+Y3QDXTOpIL6VASLof8pe94JcfepwDMNLV6XptS
+5BmdiVLrV8a+dv8n5dQ9ldYfGNpwQmglbzNNu1NNCgJcBNrfEAN7X+WQUC3OrSw
uqH+tFHZcA0GYmShFTu/cXPfeqjPrCK4OdaGekrqFe5nN/okrf7Coe7HkQZeVgSS
rWm21Fy55CN7+/XI5l/xKMp5yh7wotkfKamP3TpjozuTb5LmFBCjBsFA0TRSACl6
KG3cjSPsds1yqNBuIQOdL4n8Auz3xjhXpwhxxTik84M2KlmSHuQ5PUjBE0HIcRI5
la425OHVVfXcrhBY3tMIWFj/QT4vsckc4xYXwJr4ptr3frP8w7qVsfc36sNF3Myn
fOWF4tWASV9PiRBVE8wNQTF8j+maaVGdGnEmowzKmEWOwCLaB0wED11x0aTibYJU
lwGa8IeiuMF2b4BSWQy6wYw//nAO10uCirNAN4Oav/m/oN11LwzSR/pN0SbBpQmk
/7oYG0E/BIffZ9AlkU5y47iQVE8U9eJyRI1auwFS0/ZbSrPa1k7XET87d/gkqfss
MlLCx16FlTmaW3E4SwiDG9RP77WFneBmPrgmSrPT++yLiRLw+FmMms1NszU0acq7
86QF8cEGnHtweZKR+AkuVUTVh6fV5Np6QYg//691WIu7+Zkwb7yxBos4wAyktWl6
8DjLSRlGR1VavOQwEZpjVFdBWGAz2YHM0zLZFlYkm5nYfwjHtKxs684EVaNB1deg
SbLqlNbxmiDhG2rQWHLSWzbvZUC5shwY9+QhNbalayVp/krlKPrRzL8V9tT4mOMx
H63y+buRzqsM9Gfx7T82jqG3GxRsuwA4VpPjTNligAMGw+rGbMNUL3nApfzSXbg5
RTaVSt/O0OJufe5yiU0ZGIub/L2aoJPAmFdoBMB1jaMRPD+CBWiSfBoCwy0yQKdq
faZjLVhfQcVheDqS6ppV59k3XEmbX4Ug+J2J08Nf1/I8GsWEW52tvuRz4K/LxdAo
GKRLmiwQdXI27h8CcUVWZuZXnubZFiJoGWXbwvd5LHRIDPPSpBpP/Vy+0cSnRxpy
HNi+2boTIDb2S2m1+PmvxCdmrbOP+weM+GxZ9JJVC/AtRAxUNZ1oi6GbUM5S1ii9
xqeiyvsYAHcnzgjv3XObyBZyws6R8nO8NJiPwI2ZYkEKfhMXR4yrwvpOLaA7jQxR
VpXWRavGhSCQvfs3AEJ0flyISVu8VDRCTcYig8b76J57T4GnIR3lUP31a9XroNBC
DD9qHhIzJgDU1DNEnIoUXuzSV3jeO7G2pFuLEy1YKBgeBjTuRdmaWHqgQoijRED8
Yd05TwLoT3xiSDTsW7pUjqCNhmBQm3vlGAwuLVt9V1U5vs1YnxTgTKsWThXVlIwC
QUO/R+PgDtdrTp4s01rg6XA1n/MH2Y9Nk0u4N/J8sujsV3x0cGxIFOxNaBSxy2A/
REYV/A9HHRKXXRgccBsPFQbN0/QjLmkCWzMOhkIHE2uVbi4BrcQw+HyA3ZCZcNCX
lCmnwEqJ4HZkq1jJlhe/nR80O+FQfyo3d4nB8uCHCGl/hqObyS4sUdbmpn4LZnR6
zczyEq4QWp7tQBXPz+K5wUCcwVGRhaQ1TxL3I9QL0M+AUSCsFS+NUxLKRXwyYTsq
iRFaYotjTEDK1OPHVLHIF1evEhdEgNbaj4Kt1hMLGJsUN5Bzy/w6ivKvriV3yUzk
HsSEXmy0Gga6YgGt3lhAK3pTbio/FPa1P6bbsQQ4H1QyfjcCBLAm9IkgHI4ZAV9c
7AIVFxZ2wzmVfZmlE0nL1k3Gvhw+6GRc9i+5+RLMNWJHdZao6z7f64kFQLwx32au
nQPDRnnTIItF1wDhyrgwjNzzvju2XFYw4j+0oHFzru7W/fKaWYN5ZQadxbjvnFTm
eMq/ER0oesOlqsF8bW5kteJxJ1n4kZBNZns+9bzDzeeFh+bYr6T+jwH/S2bGZYo2
DNa3pJkQ+0xvXS1BoEnsVrn3gIPMH2P+SdmHhg2hctO2Rd5bjF1oxYORwTwxjx4s
5Gmon2l1Qwla1qF5GPLRYPrJ4K70VVwNEJC7OSrdzRuAgJqTu8/oNfVhYHBWsw8U
y73Do+V1eRkbsP6i8WHzPptnSUXePWu8RzCexMoYSQ4/OtOuYmjp3heLzgud+Rg5
Kbk+plVZw0jb3INN/yRSxMaob+xEIIwp10434owpJUfccbXKtSCwSiXkgEgsjFGl
KMuyJCx8qYvB4+dc4IuwMYysgxtLv7Ww+BKaC8Rn3srX8OBT+oI8R7dwP1NjcQ6n
jrE7X1OSeO0x2BnbZlQ1M909FktcdRhcsvvSJ95KOpqrpTa8r1rorkVLANRPMa7D
0w2dnTGeCWdf4hXkiMQqabssfKOQ9wAwnOK69dOUNbHIAlehQSj2plwBv1qf5GRE
V43wqSVdTSh+s1g2smRV9BXAeuJ5xkiI/ko5DjB/5T/4e3CPMxcESedNOUwQVoxH
WBngO/TGP0jsri5MVVvrc6ogmm4xFxPilVZ+rOe493ciqOG/W4+svxBaflnwzQrv
nmNZ9YMSlKMBrV6CeUNnohPyEew497klrNc3Srxy40MW81Px71ven+9deIf1Zr4f
qcjRHycS2xqn4UVFZ1I5JFcbWQ4s8tXNJ+V9f03vbUyYPwTonUAkTTfMXV5Ja1nM
ne3J1RTBPbhwwESx5xDcgnSXF3n5mUUVRIY+2ITJopVhm2LsrvSwpdgj+zEgG3SY
/w6CbpFa+mWV4RrM0e0d4dmZznKcBrj27ZRQEaUCQiZen0Qazwp6oZ2LrYbpsVjH
UQrIxyNyzMrhmFx66cl7KLfX29hGyTNv7tbwEbb/j4k3wdoAAmqTyD42F4ibeWgr
i2nJxcA6hkB/pODzp9Zn4cQLFuEmllx6oS0S3tFJXyC38NYIeC2odhIqc0rchgnQ
DQfGHEUFpoOuMnboUIcdqB6PAXF3ffnrM7Mw2COiMOYLR4OxZzXn/QpBkfVxqyMU
gcFTXG2OL8PSC0W4D3+/17p6JuInLb4Ds+HSG/5WHnSdgUmLKqcTQtOSR6xHVILw
SLd93+i3YqH1RAY7C5cMbSKMrbYCisl4tR/q5zfFjElmaY8rIAWhyWoGwH2FivMx
w7uq7Z0a48NNiiLLNzjZXO9cufvNQZ8ZlPwXOuTcCWlA1cnYE4qDJs8iI5l/3maH
/4SAA0sFEococraXxT4lI6hr6c3O7BS+ZnEb8SPGmotD1nEsbq2HsdUCDbzktBP8
kGwYaqUoWGio4f21RhMpyobjepkGVYmvM1GxiC8AIkUE0YxaNaeBL/4f6gx4MJ4N
xoYRtj/yuZCbcKJxD8DHat0bDDEM7C5bB85StWY0dxiP1HeMS6sXPGzFpavbO1Wh
AVKcGX6m6kPg18zJQ8wEYjgtxfH72dS2wzF48dT1bNwYcMTGttkTxR58wE7xMLfc
w632/aUVXr0k1ofvrW6i0PRDnrEcXsvlZcpUUjtNPaTkJgOxI3v4evP96Zj4Ie5H
9GbVkJK4ubzYAn1XabjxFO7VNtI8k41c32ZCOO+RNRozuFDp0wcee89wmZikcSGr
DJ+m2C0jd2UGGt6xoLv9ecIS1TYXYu7QyntTHaeMdO7yMZp0mDNz8cpc6CUoAMaS
ft6tDc8griL8wFSf3lWv+WfHww9OlxXw9revFyA1srKXNRDvo+j5l1dKKQhut4eA
g+l+ZoKA00DTYKKwU3AvcmuP8sE6oYW0ZJ0SmGR4oLiAoygq+qBMPKLXREoti3TC
UFx39StUEjjgxuNhmLSfpJAgIHAQubyecgjkgaY2qhse87RMIU4ahhXKBWP8RmLg
pLY5O7hCNOVyVO7vg+SJhA14kwgnHVzF9YHp7+Lao4nG8rKBrFV37ZrHkVt7XRbg
cpEiBzgDNkD4gJMbKlfuL+13N/HX6gPvYfebromNYj1KnhnTFWW0kqJMy6/LI+cp
u8TeJUt+LGcNjWVCGHD/Y/9wwsGGcnK/o8wLtyFjFZHc5jA1tFQrGx4CNYvL7c9Y
RiAsffeIAbPqzZyVcMoMDR8bpJDdHnvSzIX/0ctHviz887PMk77VgGGOgWHcs8Ff
2iA1Gtpe3u1o0gHhKl+rdhoyo3ZPSi6iaUmtV2Lo+YTTG83q8wku/O0klmblz88B
FP/xNYNbnfSmSEtUIFcK9SYKqjEkdduDUgy2TO2m9xbWx9xEcb12zmstCyVWP4Gl
Jw6yOR3bambOxsTeRiZ2cMIGbJ9iKKtHA3WvOnxBOuFKnkjq7Ftvh0eegzj83dO7
nxG+e7hCkR22BocRy4wtgSdoU8NDAg1tKZvMOdNvTU+W/EcikaSH0jBfqGaXjIAe
oEuWQx2eTtQSGTz1U1640XJTxOotukIEewAF1VnzGnlphIdm1CbnFpzCPp38sgk8
KT0wInNTXNWtvDihrzoxCn4NfOm0uPDFGuUeZBLoOpNmlAxGIPvM1cc6wN0i0i4Y
SuJEDmLDE/tpBFm52aRPqXENyfdpvwpDt27KuJ51hNjvSDLUXV/4laPqzfPQPTpF
l91apU0hBvX6EehaPiBCJnfawD8X8fXU7eytVEe9mo/WjfBye+aTc//WzFRp0ZGs
mb9BwhVa9skidSuN3kTg5Kv/YEswJiuRYNTsWVyixo2T0MH7PfHnNomXfVZqNTvA
xpDwtYbQ61g5Vbc6U2BGVWcCetLGvfDVLm7Q9dusO0ya/QbfYmQQm3kHy1mnVeWo
Wk0QEnw6rVXlkkfIy96yy2i9n7wiFo8CFG1y4nbVUwQfxQXOhWNvWn1DxVnx4Wog
hy6GaGGDstMsG+nmJcf5amTr0yi9MZWa+aveuz+o3/tJCqTLm04Ko1kQufLCGyNa
GUtTZkBTzFcQldGqLwKN2GjKg4RC38buLdTVJ1dvqmRAOjL3/bZZUjPjiAHHJ9fH
p0nIolPEos6xNQEJtwdtmRt4TY9Bqkjk3DWJVNech+U8Xqg99BgW/SbNkBjqM/4V
ZRRvIurn9GawH4w/bDATWboWa04jhifg+7/4i3a+Ep+omzt1QExVBQY+qvQjRWrG
7a4UZC2wOASiydoUZvqwGWVzeZwO/9kom9WHwe51OSAOHAcntKZ4iKHWVJTsbKp+
s9WWDH+JDpSoQq1B0yBY2/DmWc1YwLokagWHI/w0tv5k4QnjhYEm4biAxLw8lEz0
8Bo6+SImqm+DaKyNKOF18oHuwLDWLm3tgWj/grhP3l+vunTEV9MAka9m+/IV+v8g
UOLocd08CuCLnmcaYgQD63US8SVucwqwHJhxAkxK1kKl9TmAI1JbaNUeLFHIHGDR
/aBsRcno4KGaFInjfKwbYRm0ctO9JkswnogTHCqPi6CPOcakAtJjXB+BUmDECtBL
+kWd8/VBpSL99Ujiq/S8sWC6X+yPvkLIW0BVb0ONd9K2fRFGUXK9+hrXVaTgcn/V
2x4MFlrH0/rC6aDcowAxAx1Or/XcEYlxFK7X7JSrcnGlSyrx+Yza7APaLxyWuLKg
xgLJXcwnHlS/zgHjPbjL0CX91Ch9TNeM/qlz/QgfCMvZ7Nf7KDuRUDAauuHywT2/
lgnyHiK9tFWblAfIlsmp4B1fpeOF6LlodYTBQecBgwXhd5/lSvBqJSSK+sPwDjOb
nww/mDGUklUoSH+HDdsiSmeMHzPQ7iF6UyYOQyvO1hqRrJlUaQ7L3Y/i7YQhXM28
GXHo45Y5IUxIBWtoPvm9COD0Tj1lht0LhX7GS1It9zjdgdPwe5pWfIrjVLx9XtTM
6mm1XrvshdJ8Uz37i0ktR3uCDuRphDoY9iRf7UY5Ky2xLDW9zCkDn18wEUw4Vwqy
9bx7J+gXDw0a+8YJ6FOSz0pr5fdU8BBrm2obG7osZpaVa7NAZE9VkMA7wU3xwuuR
vxa17TiOrv74oeWCTl1LYf2P1ek9O3ix3KLSg49g7t4j9RQoEECobrUcOPAWxlKl
bhueGmp8zATIY4BmjDguYnv4S/NCoSi1qbQbw2RDwpguo0PIKA1OF2eVbjx1PHJX
i7c1tRF6dbidv8ZYMZ8xr0kit4BPkkWgW2vZyTi5yLvWZzD7zK5j5qHRrSgrzRnY
KMmNt6LeXWAgYrhqJgd5i+XZ4NWgcaeNf9HVoFOB5qcZloMDowyaU1bnh5Rgp9yE
wCM3qweOcklTr5cfu/xtEjycBY/DsyL6y0Pn0DU/Vd+yq5ojiQfQds3O3CL32oNf
KNywEXe77spuP39FVagPc0JZ6rUY5w7xqisOh0U6ami/QmjU5OUHzzGqFB0MUR3t
3E9SN8E4SfhBiwiEpyF8vokrjV7n6P+6m9/zVh9ajb3hy2EgnfgN5spjxswrIxTD
i48KaShyDRa479+jv/KdVXr64V2hZh1A2r0JUlkk9zDWPVasqpPqi6PPDrRSOiNX
H4KTMjf396ZrysS6QMFKtNNNeHWMVQNAzq+jqs1BOjVgtpIecSfWctF5GEX9u+EM
3RbjpKYOMaMwfylj5nK+cAPROf9xk9OYt0XtNYjclYA/JpliWSFHKkVcB3XD890m
GIwyuwz9xBW/Z/oI4neFQ1hC8E6ImEK9HQPHfgLn2ssI4b88WHrseDbqVq/zKr7l
C/4mwzcFd2IPIcYg/en72ZKyojAvkxtEph61mmOPNbWApxQzmokKb2srxy3ClgIl
Bo/c3hbpso+8kspiHSNkpjUtuTZmUF+yqeBKMLKePRPvN8Q3GzS2PWAs7UyFAxoU
fXClSEB3b/nlHbZAdKB2FX06/r8lPNqMNMHZiykUeCuxNJOfC1JVLR91gjoR8+er
M6/acWMwiLmJ8J7G48KfOIfvnN9tArFmc8s8rxY1WG55f2o4KZVdvsN/jer6By1J
amwaJe0dAAknvebZQD2ITSVONjEZ4XRemPiv5B8SRt7tOPGBotkxuaf5o/yeWkJE
4wCkq9Hj3xDtmZOfydSIc3dbJxQ69sPeXtOA5YsnSW8O1xJe37pLQTCOhK/V7msI
ZjZHzA+/q2vR6/ajpNUqEuO5ob9Rpyd0odaf2eddzqM147SttuK+M8Njv1LIY8X7
augdEiIYEFYDF49qOpQmqLkQB+TlGH7rXQTiMWBgkOfzrZWzEsBjy8IXpN/qrtzp
2xaMROBB/J2y6ikBU/siBGIRVEL2pIA9T5YAo7x/QTETYDtxZ+oB4YTs29ssG05e
zTQZzVA4+hgUxsMcl91j5xeEmSRySMY0lcDbLRsUmEYeX3ZLKhssg1Py38spedDp
HKccgCS+ZuizuzVfNrgSSfFIDrcF1g0eKqCtbWTLB1qUgFo1OAYqbPs7dU55zyif
7ABc8XATs4rsOHYi41RPTSHsR6vK2Eez3AU43acfMUkH0/+HiGiPNOdWWK3CEeQR
bRVLuHNrYO4PvDB4cI7Ux4qhN0VDapJ6EGlhRpSa6CI9AcEJVoq3LiVp+Qx3+3A6
X8/JIdrvpmHBuJTrVCB43Ew4vEWPg61bqHl8xz3xoSVHXElrU3Zc2zLFFN0Ay48q
HnH6SwNLBNMZMvT+5KD7a+wR+wh8Vzwj9W4/mmgvo03lM1+Bd/FUD0VOHsz3jQFa
i1CbP7AufEIvx56ReUgS1xTsy1Gfn4bPaIHZSvjqGCrCp8ieWLMPNFXJTLelW9Qw
kUWzT8VsX5x1A0/OeqiSxl162t61Rl33bkHvWim/aONELGtcV9+6Y+gE3AjxU7AN
JZXXAn4NzbA1pcu8ZchQMSbG6v4756EOe4eTB/qeApw4+8YtWSN4Z3liM/B3+v5E
kyoQp8hEbIGRNYS6Plrw/tktc9y3u0ihoxk1Gmjh5J+hq3Mcr96rBgyZyRpVhI1S
8+Xx4hoGVVy3VHX+qgGdZtWMEHRcGG06pNpZp9gu2adnsW/an+CpYT0hFL2G6VUn
Z8wflVY+gXv/KkPR5tvQe6iJ4dY/l6O5pHKJwnj9pRYZldE9e4JYRyGFcduOxm4o
jXZ9QsIGh7LwFf1Pk4UyviC9yv39yrmCN/uqCvIPi0A3m0OOV9BRI9w0OPIv/2Vy
N2tW4AKg+5pzMIjc2ipuDMcyFDhx7BRJXgpIcO+cWRJzBSrqxjXLm+PeyX8vCNDq
77icev4dztYF9a9IBioH1Ziu95OxyEgvX5i853E3z1lU7AAuRJOG5qNIA6eFtsbL
PkxULcW/+WdH4imflRAlkLRt9xO/xkAOdZz1TEhNoqorR5Db0GzH9opGaYiZV58r
RCdvcWXnCd9d5D4z3feQ7+rXPwnuU20KcAvEOZoKPrBQkOh8NU1x4tr54jwcfZ1s
9wEUGjGHRBU/eNXEWTYHHlyUX1QFRxn3D+9OdNf+IHX9/vvcsW0h4hyL1FVjUQHL
Ixhg5HO5QwuccRKM2xWnU+p4YtMbqDy6NblQUUFObAA/jes5ZBpigPM9uTRVFeww
cM71wbrCBBJvMiQzbupQuxtTWLBO5YwDhBJmlqBZ/wTqgDlyjEkTB83o/yb/5QJL
IvYbd/eqPSDphfPLUM/6XLjtQiZd/05aa7DfWd5dsErcYp1KnW3UwNycbWf7KwbP
S/s1oTxMpAKPiPrqoYLJS5wrlhQQpeIgDglZ5NAeoRiiJsXTu2C+f1gRk39ZqzYh
sq6bP8XaXptBPBV7KPHwFzWsfMknhnY9fn9+NMnlESjvWlUO5Qcl6LJmZ68nte+k
qkss96qUH24et/UqpYmjpL/SCwRyfrm/imxqqpd88D/7sK0uroffhjTSiu4N8qKK
De0qnhe8vWyAIi2Z2x39hAo4eYRG5h4C2yi3DeVoJ4F6aoavyZS2bXc3d8hNSNDa
MPip7pq0zLzv+XJ8fZfa52D15P8Weyr4Y+9hKSTPm2m/BX2RBVGf+nYD30OsiTSi
e+4bAN+xzzUs4d9Uv+HzJF1kagdG2viWspa5yT+OKn+giCy9mayzMjbiMmcD94zV
i78MZG5QHLTcDWKVREwxdE12bsAbHu13hdsAFfczOKiNRXHPUJpyeUUc85tZA3+R
EufICFrxuNxFBZdErbDliumN60270VUFAeSmjT89W0/26BxwGGKBz9D4W3iw2T47
DMZsxVa3B76n4Z65o2ZWVQEIY37PL4vPHWI3Dx8EaaScdw57LmMcj/91H6QTJ326
R4HqQr0vrmhQrQVowJpQKzhnlYeLy1SXL7nWKmynayItme+lwneGFdDaqAV83Qfo
EVgLl1aT/VGQ2yqFEhXOrKfAMuuDy+Fy9OQgHRjrGasDjViRMOrxqLH3WmooAF4d
faPp1k56jEA8Dun6jq5uQvuS4+DTVSyyeTUlSG5rPaSJn9ubBIq4BTPdBSiPF9GU
A01e8xLqyeLIbABgE+OdvIYuhaBa+x04pFzhbioHQbp2UKENj89laHOFwkZUVdBJ
p6v+ykeP8lVFZ3S8y1NwoM1ADuo+KkyAcjEQgE2ORrlavkMBTeXwmT/0Lok4cpNy
ehaY9n2jd995VQvXgo6+ea5rA8Kz6V8/iewpjMo2uklHYk+e71Ubj454W2yxJpbO
ffkXqulgvqqp2HrodZbEHx45u2jeH3XbmGLlvmSNrjfTNAbeWLl1qGT8uvrx7etD
2lxv1DO/uPwaBcZrRSmYN7XrEyGbIK1pViXk0lasRmM0vZfd41iQwVtrF4hE+Pod
dqzoRWUsDFALNSwshRA9fdMo8mYiIvRcXhbtDGagKv5yDoZL1KQ6hQpiZkB8Ue+d
pb30KEWPai5+lRUrj2l79MOhE5Wh+rnG3vT6ysbaeRmmcdGtCTQhUyG9wIaVzBkO
sMvRHDQinZm1dFaiZ5BY1lyFgvQZr/Bke+MJQCW/Z9LDVJKRgm3zGWfHuwfMzWg+
yvlQGENL7s83JdRwBaQyUDiBLMEdVbcJXk39BiB80WrtBW2OvnX/eTNSXVNbqjOz
A+4B3riRZefz+RV2A7pa4ahnw2HsR+Vmnd8Hwnncn+fvQvhaPRU881oAWN4pgT6c
zcm9OJFO7upqWYEa6f8of0kuRzDfjqYy92HklWc3FJyLsyFHTm1MBBozBLhTMud9
goYc8/eSR+EgX1E4zWvdjFuFxi9me04lCoAAqv2ZRDAVUepjByKk34Z+M10QR1IK
rBedqZO3hMh0YajSyU9dCDsKp2+2GWpJi1ijLxvnuugSwh7HyS883kOQjE1n5vXw
2SFKXjnhdPkdKj2J98s7GJSiXQAlSxWCM1Is3DMD6QfKc3Tt9idcQnqO5lq9YBwn
3fMrGesjSuh0rbXpwimf+73GW++3H4VCoJE2kf/x3/EqbZnOQIN+eTtkVGyoHsPt
Xbwc9iS8qQhq92HM9/QAplyC3u0Rc9AC1Oi01rrzju21GamEsF6/4TepTNclqgrm
zp6zhMFRf9mKM4+jYvDTpYipmHv7qVKPC0YM7NIQZT0IRhqHSQY66pfj5pd+nRcR
SrllKybYkNqV/wIK6G4fEDdlzs/Ta/aixh4s81vG9ut8Fwa/tvGeruPBox/rK+kz
bxfeJToN62r2Ye3Tm+9BC2cOP/L2/IqaeoTDv6DKwuG6cj0odWJNX8/35oHuAyvZ
HFjtJ3vgiLGQw+O5qsE8+ViSpFjQyadZB2XDlKHBFLtvD8tQkEFGFGDSFmZfv96n
K8h+SPuU6pWNCBak5AxjJfSGrZYMYbE+unKIKL8YXFhbBCZuMMnipPPfWpMSQIOK
ap/lntC02kwYTchZaRkfGgboomcWa/LFnefz8vG11cKoAIBoATSX+GDRbAviIA1p
HuNsnAAdJpTI87go91g/LmYmgLlV0uQir9z+Z1PsdJWHBDb3aNhxTnog5KCZqrsa
v+aJ906p702oT3FHvHDzuqzTAv/oKl30xVwRNCVI9Em0bGAa8PB1KxzdlpUfRAFT
2iIXKy00F3eGnw24x2No+ulMKeeR5XuqTUZEOMGtA1JGL1zOZhNCOY/qp9qEUsaC
E/SuwyVX5hZxHYeyJiWdHjmW8X9FjABmwdJWaqJVP3rkyyY0He7YXlUmbfogLfP/
P7c5KCzzttLZvITXMZigNhyAcpVErpVCQtdN7F1IjVVWEz25jB/lC068PMqlJY/9
EQxJvnjDfnb3rxOUm2kHLnKC6wfmJ8VnHaInKX4ZtMkYCm4vz0zAzmYXA+hCBUWM
XpdKN+F91+O/xrce5uLxLtPW61s20PhSh7IVXzWnCHgJnbnHt/WKiwt2yYikU8mT
OwXl3hxUnGw45hMvFg35r2cKYQSA6Vwr0WQ8KhEVuoCwfG1JGPCq6K6EgxvSbhQ2
NYDPRna2coxmZBR/kDaqyQ/XXKc2XzIn3e5m+oxSQ8QqVmW4luoYsFmAd3zsYKcT
csA6ipkpMsPT5u4PUeh3v3ybetUZNVoX6Vp/3FJSWCF8AZWR4nukqJ9dNt0qlN1P
DKxRPNVfpJiiBznwwJ3bbJw0pGyHQHrRGixOPHFcm7bjlkg5Zs+pQesUYzXcdw/f
reGbqBJx78rDcUsAY/tAYWzqMrMVCJ1CIGEGTPrDJWzNI2gmoe6a4Hn9I0WBM9g4
qDqErHcuy/gi8nuJ1f3igT7Z10QgwuHGDLG3dIsQhtVrx/h2CzKn/M2vtGTAxPll
umDdLykbhlonC9qcS5r96AFR6wbBfyXHUeDGQ9PrIldCI0ugYUeL8kdyF4mR+ZhR
i6WVaFdh+/N0KIPtuDxzTTPnnL0OYYNpRjuX4VHpORQdOU0bo9KUG7d66DA/ApVj
UKMw0ljvOigXusFlJ/eL5m5XOVLtscEL8ZmVi623+qNzxW+cIwFy4FhlGrQJGzCP
0G4rOOwEuXXwuIKNDfh58TAI7e2mrpmiY0KwwxsB/k3KjVdkzutv6JcmPZciYX4w
cMN+LWvaPKO+eG/xoB9aOgDm21j7ZogIcMhpf0RjUJ78VLu2Cj/AQti/mBYCKodO
NGkozl/uIEz/hOSuDxEwMHwXA5rytGwF+HOt3iLJtOmBWH4SIe4PlwYxm1S1Ib2S
3yE93OfNzknZLc6AJKxh6N3xAZiyGatSBqWZJZXsJ26BrviemHygaBiK++kF0ODx
cmmPCVleYmG5vSGQrrYiX3Aq5g+tOADZerE9ZFGVglloSf9/wEuvtOo6adL2yVlG
Ns8advVHs/yNZQ19ZW4DZE6kMGpZVL7LDaXR/Tz1yuDu0dXZSPa23Y6+LeyZYRcB
p8DPw4c4yEYkE3UvARKMOw6n2zHkmCZFUCpehriW1E/IFh8JO/oOw3XPAvAXkHNn
J77/Hu4p0catqWq5G6F2gKe/BaEmUpyl7OmGGO8QGcFV0MC9rMGIycOOf8ET2ZaZ
TYunFP8xxK9/c980DFRO2g/5VQaJLc4U/KJK1aU+Bq1gYPHtAivJUe2504vipm2U
jMKUvl9C+eldnFw6fSUP6HfEhFZzeT+OdgAbA5nztj4OHZjEQ5uDFQ1dCURBO3fq
WbhOSWycVL5UxGSdTwqK40ykBGZhZSi2dWz5ExKj/B44ivEv+4XHtokw6PuiPJS/
6DqkP7zPOhJIRll2WFXOC1YKc0/dn4mJlcyCuZlZfGksEY8dh8MD8641V5/iLQEb
zxBnfky6XJxIjhqz0eWs6U0ZO74/Jag4s+f2+tbgC94acf1SUUFObS+j5inHfqD2
6vFlMyaxGI3FKKT0QNboT2D0oHDVywNh4pE6kcFak2YcdIRJvWwyywIQPIS/FE6O
r3CgGT1m9UFb01BWMM1QY4f6Dq+bzP8vLlFlnjs2TVfW2i1yjiqHpKsxuYmC1iPT
lct/UNzNdvkZSePJ4AfyOl++d/b5E/9X2JqYR83dVaH4LUGukBsPjo/rFs2l8euK
Y0wZWx+/mVl82/pAOtwElfO3c096sl//pge+VHbeod8hICBrDBHC2QuLimCV6VHN
wOHswZvLt211C4Jfks+5oa+HbEOTzmhKwViStTOU6gHJFmtK6V1TXps6UCNtfzan
nc6cfooMrjTPye/Ewf5wExq3JbXtsJftBCVCA1Zk8GaXqJ3YuBGxnHZJ8fIJwHXV
e0FcuD1u3O/2I8aqirPCYQUUM60g9ggVC5ykegqu3PBKTNqR/P56ZGloJMf9rWRz
X3HdREuzy0bXLdzcWaX/Te/og9lZq/yCwfkIL2EwfOJCX0Fu4F72tQNx6F8OEhA4
8HCSUfAZSTTakhcBnCAiP5k9aTTVWT03r8qTI2/3LyMxfBZtwV09on4o26ZY4VTr
cpmU+TLY7L0pMU7MU7W1epovj/cGsDfqPtMVdecusmX6pMiefdtUVRKc5un4ERQo
qyLVUnjIJYcRG+U8G0CQLQMA3kJ8LwSIVqB25g1NwIFoxSqzjwFsAmyIylPUYTQf
bBuGBNfbvmnTIVfrVWh/BTrP2lsB0T4YMBHJYNTbj+RPMF0ekYCFYguffgCDtUrS
1r4hde1O2pC8xSo3YeQQAZhThph5gIFQVpwflpci/spz0et0HrhH0rMBfT5vH87u
7HIgLDGFwIMasZUxXLUq15ILnot2HmBZo6dbp6puNG/D8/gRxHkOtcHpR5yEsi4a
8hvIhNHZGVClTA9uf93egldu+ZdqisnYflHOFl4woK2ySfx1odb5zwomHjHuwwhU
Zj08DXu9gLDdczoq8RuA5fzLDvTjSf0QyTlQw7Kxi7+aF8OK0OuN26DAGUtskZ/8
oJkDhQGzGtXsRzJbBGKf1SRYItB1ULMnEe6rxSICIoX5jymwH1Hg0uVeNWTr3RRI
14RKf2DZhteqBJmlg3/hL8M8kL77wBYOYLXL3Bdmlo8POKo+KPA/PiKzz88k5F3y
nv62us79MTW3DDHDNkrhlJJT1dfDELFqw4TbOw1FMjIebCxqksSM8nhfgDjahwar
at5xE9jWfia1kyBpDz8YahuF8f8diX7qZjwN3nlxFnWSfrIG0fkVru03kc4MIjLs
djU8CXsjM041kt5qUdAbyMcTrx5CPkQDhVdvRNPx2e7yEbL9E5zfglyK4sKLkAM0
8Bb2tn15cTJTgrRqe29Cr7jx2AzYXBiZ8GqPdXXefGUukYuIlyiQbVYUd5+vSKq1
iwbWIFHkLVnHGn2JQa36gm+KrlTL1f214gxGqzBjAd7M+KOMyDLVqA51qmRGF1T6
unlWFMOsrOSstc7aAesYL3Xt2Ed/qJQ0IjWJZ2bVvvQyySSeKs7MBUTvZ3RSnMmS
CIjCkb5fyft03KAudWM5tH20cDmONFZdx8bEiLMDR834tPhi445IZ0TICCQc+LiR
uGQHABOCFq0EUBshsFtjyurqp6ohkcb2e999XuZi6B1OeSUEN5msHXdHdEu5CDMz
ykxKCY4EmbLoVdbdj2h4kaCixGyI5wJEUwFFugxE7ENePWa5Rc8cR5SLEADp8Tlq
1Ge6J0RQ9WSG7bMU0vWJ4GXN9xeMrGzJ4UWo9iZZ5DtUe4CXm4NVsmnA6vfnzcSx
ZfDKuvq/ds2LjMtXNSovhWj1CVGW8j5Wx68CCk+B/l6pG5LdKCdWjD1VkVcaVdbT
sXEQT/JM3q6Y/Leg76R+QU8BUsjUjdyP+/7x9JOuwMRFyQs3EEO9m0uAVTovICxU
LKUvz0weUQNacXQQubv9lW9L/2uMogsXveB5vU3ge6bzEasjGweBgS1ht8P/Hvyh
gD+4Mayz6d0l0HjXnfk8le6JDocuk9g3uco+CeZVjmiMTCNuqj5PPJG33Zd+i7gc
XeEpLmULWdyN5fk/Po5GZIiCX2hQUJvDpVE6mGnGtiUoL8PsE7TSQRJ08sxUUIE0
W2npOVIahiJUpP8BpQ33BswwdpoMQnv2/OZbLkZW4dcPuHa9H9ahlfXkL3+/zEYU
nI80dBlKTNvOrgebXRw3IZhdJMWKdu8ulEeUNPg5Ad/u7X5YuV/74i0hGRcEek0O
QOIvWS+mkQihv9hAm9aiT8SvgFIkC5gkonB/EdHXn4M2kG9Ewpv9j6o8q7srCB7t
+n7VOLG4GvnMXfzKoJy4rmsUzVQt7pIFDHj+joF/rJPUuodEaq1zQRd75/PVgsmD
iXk6li8+KAio9mgbDDq/owLl7xALaCz3kiia3DucN/uGq7cB71KZ6c7Gdd/ahA8h
jG5VkR8u2fYaV6gek9h8hcGhTUwbWrpLzwADOD04YvNLtwV2StB7nYrTsqIdj4lr
BHHZo3oEgfJLTLod6D/BkwR6qn5zVGHhkdorNLDqiZNaIm8Ea6OFH18Syr2525yw
4jDC7hb9+zvC7m7p04+7NRrDowOxwBPGEJCfAuUejAqAaZOnLPvVVQXzJilKy8tf
shmNVH7moEV4X5+VRfXGvEPmc7/AzkwIZC6wOwAlA8OlmSMEL6HUP1BwZk1nTUje
8qeKgMYSoSBalEP5xREBw+pc0OMYcKC8EeC1fMwlO4ZahD8/GlyTbD+gPoS2xXNT
R5azrGeRcT27hdkvVykL23RBjtOo8VJJgBBNfVX700ySRCVvH5R/5unY+peUCA6J
xmozTexWuN8gQIzkcn6WrwiRG2znTGt4F+l01gastC6NRCU9f2gXn1GaqDDZLaZ/
JDGPZBw79upnZuHJBosSrNHuDEQtoOCKH4aPujraINFeWzx1l4BBkrhcCJiETymM
S4IwxShMaGW+206OEPiivNWkmWT9rwd6cqMZMScojpHxuRijYHx575Z4cMlx3jkk
QQ9eHb+Y3NQHMjzDM29QYuyP8x8v1B86D7yiB0Z52y4d5TMmMSNJlvgN5qZ+IK1E
FLcmZZkhWQZlJY4iJCVJx+whG1hQLNPnS3WzN7NvRMgfyJlspIpcN/vphl2eDDSC
iy+dz5ftNqv6MD3UggVMfSlhCYTmjHnORNNxg1V+EdCJfbxYmFJC92R1CcmL7hU9
1iaXF5V2TJxRrjWoytKQf9sSx2QhbdW4+um4yvLhT28qLLyYJykl5Am7yA1OPdV3
hjjwLRr8xtm8NekH2Qbmk1hAjWtKKe0Da6hKkmzzC/HW0hnExucq8fSgejLgVV35
wuiDjqwd/x9B1XdlsDeNhEV5XZw2/WSOkzOTKhNVIDQ+ehcL3akU36SgyZSfOOKv
J4BbGnjspFbyUnpeV25mrrzsnLwdO8JYazd6VTfK/DZ8cEMGXUAK2jlZidHJvfDJ
2JEjN8dI8GqPCMs2jcLRRYibFxt0tWlWQvrSDPLboiCqEnMFm+7C/7SeQoUkZvzj
DJJLec0grU73pNDco07Q21KV5s0bRzwLcoGLLw4pYkZ5quzXmjzVbPL+crEyZSSv
/saT+hR01CtFSacArV6Bp3GV14jhdnTQ/Srm5R4uVJRG629n7KGrMwkNMBQ9pdRE
a+uk6MnMoouHrEfJS9iJ0tvg/D4DktSQHSZ+7p88UNioQLT1YvUynsBY1henk2wR
morfA0vy85rBJFjsqGLVPCD/QQWjteh4uA9B1YRKRTOc3XbR/49w3bgrbww2xvHs
S7XtkT0yhlN/mas+75W/zd7XdqA/UfynrAsefYfKevpyuqw3+ri3NAc82vOk8umF
RHuGcdLEsLCGTJBxbYnH520vOZGmLehM0PPkTmZq0xVJLZE38+UabHMRNXq9J/1I
3+FQn4iZJOZHCyCJPCtZkdNtYkzVCx8QOZaT7xpnizjjq9/McPWwjBzhup21boLY
ALjJskaSEemqyjB3BFku43XDveDRhkyEPjtPKOvWI1fnUyGWmDtsZ2rL3QzP/Rq8
+waUeNdDXz1ylfHEuADbKnhlMNO+KWwP3Sya+qVsjnyuNQiUOP7/pnK8uvS9kS+K
A4kxhpxxjPdoOWo/1Xo8Zc9+fNxFSPGL03NRgu2/0Mrw3+n2zSlY3dCWlnLVmhE1
fndy4bJGn9ayojUik5runLQq3rpNFO645MNKn1ShaKOTazns7wsStG240+j8TC4j
mtUUsfdLHurskXQojozZ+WyDASHEeP1mt1a440+pVfXWxS2EjF7+H6gGUfOHusyM
2yrWkZ7FCHF6h5+CkPgHzgpajY+0/Zy5ehe7GX6XdjLU3AefvXsmpjJM1nH+kIqG
I9h1xjP9u1ByFlVLpQLiXaYbd+zBcqBCuP5HZhD2fDxaKDv5ukPPfYgipXLYMvwO
xJKtmUsNw7bhhOV2tVfMNb9ET0Y1HqA8oe4bRHD3ckqyonzy52QuAuVWVHBoZ6Xl
DS1nDRrVKJVd0PAInJksl8YB5B/kDSXFjhacKzWQUQavw3fOxEL9JBqJLj0BnZUt
dyX0XECU/cXIzZSgSarKWgkzlJ68tBe0HtdpcYqQRGu/KOmorpo0niqzbZDV2qFA
JamnSvtvW/r6ULStzNDfolbc1oJY53AXGZIk7G28yHc=
//pragma protect end_data_block
//pragma protect digest_block
A5WK+GVZ70t4YszdLtLRSXhUjYU=
//pragma protect end_digest_block
//pragma protect end_protected
