// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
iQfegRC4+9ACI8/9B+UEpbEoFus0ns1YF0Na/p2jsa4c/xhL6evsaPNQZbZ/WmqLESYYbXsCNyxz
0JK0GuUcB+9WlO6rX5nPQ13dJni8wv1djbqp9cafEgO0jzuEjEN4gDLJ1PC2V8Y9tpAX6QhfBlsC
vyU4kMzQWxC3fORvFIaLQ9Uf/hJVg9ZlK5aIznlz+u99Gve+nykb0e/lufpK1ImvTWi6BVChYyc1
hBkDML2UMhW08eDdY4OlgCnc+P228wrDy8ptcD6xT/8UBgo8SndmRJwFY9zrrbcH8QR4IDJz7GDT
9yez/fDN+BydNZSeAPhryJRYLmih6wHHVoaZJA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 1152)
Yzy8cAxBu71FWua6NLE9V6BdShz12/dulEsrYflY3AJQAUKXKsEW1btMLY3opwMe6P/w9f2x4Loi
XCb6IYhKfbjfGIRY0DJcPs8OmN6ujhg0irUy/zLo5BRzw4YW1SNeDVwSjSbZtS+3MAdA8pfu+34O
+1pX3hroq6DTdTAD/3CpYmmTVDBpS/D7NccdcFd+fL2pSf/K6IDRAhB82jXiL1DcczdcCSU4yFcE
rqcvLjiUx3nLdbAxygyhiG4m4EJ5fQSar+24kbKD4KmjRrUjaRuFiXB71/3zglNN8hJr2SyBfQut
Xf4PAxCaL30GsCmBB+phCYzI431Kvht1dh/ODq+XwDagU9F5VEjhs5dcwsgSESEoIz2lhL0A0weQ
yIWZQkg3VZ6TM/TTG8cB7pyLzI7FPhupjVOCSoV+pS6iqmPiq6P2QLu5WoVKQ2vyZY86d3b3wzA5
7Y9OdtRf6+5G7cBWKOPprWiW+MLn9E6CF56f6HcVF15TI88HUv4/ukMucpIhvQ5JpkPqTTDbvjjj
x535ubj2b1p377XIDUMCDMQfu/MGLHWq+2YhLo6BAwP3bEzGQekdDeny68K3C+JgVA3WdGO10hOW
FJUOX2p3H6BcL3NJdm4wdnl7YqdjF6g7poHnuojAQPWQI1KW1/YAEiL0mNo6JQvDt7PsrfKAiEUh
CWbRfCsTmg/WGyR5vWzVOUA34iiiMwPfFP22sM9tHUGL8Xy0sQ2UQxop9tqEfAYHk6zaN/FOdRDC
a3aXtUpM601Z4y//xvkhSxltGuPM4WBISa/60hRDaQ8mGBO+lnMrMTyUEBX3pyVMRBcsikMawT48
f1eCxPaz4SpmMXIgCV3FAnAtJkARByTugyPbAteHWzGcbzeXm78fxzrF2Mbwe70Xntb1hIr7KxEK
O3Xo6RQRtSmNYL/ZXPCjtH4wJG8DFiqezrA1ZFygq8R9I0soJmJmPW6XPGKcC6BmcWisd/eBDsh8
9QaNcdHwhxJZtwGhilrGDzTC27rnekVYM8MMMHB/DKUib2xrmqHzqrIXvDUUM53I2UajAwxaU4Cz
zCw+s+2UzkMIpV92KVUXEe415GCM78k6suuP/jgIkKUQdUY1Qjk4TWx8SmDGG2AB0lznie+C2zbQ
XCV1Y0MV8GTD2WeIbzY4EhK3wzstTFBiW3atYH1NWz09MmDGrfwgZjWAqVz7HPjTrFyLDQSRvyM7
UEYTnbgiZmsiKkVryKw+MsBFgsf3hhSAZ1i7hdj85qcWoZVTLBZe7sJJVLudaNET8x1i47EqcbAW
u6njgKixnhDx0Rz7Eyso/5lCLreIix/Ocve1ztaWGzIxgEHGcWw2P2WXmaJT0EaArSnwrxePIZ+g
ELN4XCeHbanVofQeC5oSHHshcdHmCx7Jg54Y0gmVudZy632oigtqOOho8qopX+3Xd0aq8P6nFXuD
LoL1fbpQ9rdNTph+5unL+Y+NAhlLO2Sq0psFoM8WWdYGbeAC/yVJSlPFKIMe/XFEJyvRRunyfpIz
rg4Nrau421dGiDkj
`pragma protect end_protected
