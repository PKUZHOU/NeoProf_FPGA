// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
sC+AgPXUv5lRCSohYlvFM3nzy11GAErcororOYprga3elnuIvVw4cJ4MqxiKJuYX
Qh8NHKIpl8YVn06mu5ytwiwobFzp5EvUHDKqOc0C6VRymH0ujEFhyKrweSAnkxGE
EyFOR18jaODiD/q0bArKQPXWv4oW3w0EtdYt1Ck1xMc=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 8416 )
`pragma protect data_block
jJMd8eb6/pcxDqST3j1EcMV8RORxGOldnVVHWctCX2970EF7Hha4SK+ewklcRYoi
faKOHiFGCcxDrAqMB18d9oax15jTpTlHQHu/V2k3+9+sBkn6dFLhxloOEb60Wcar
dmW/56AISDP2ykZEyihXz8aDvrnvjiWn9/qO3WahWYj5IDIR1lOAsi3XYTxWvLgc
ZohSHnFK3L4zdx/E7S2btBVShEXMfZXK1N5RTm19NvrXilVaeYoj75zxNyw8cp8Q
6cDCRr37rx9W/d5OgTXpPs8xOPNKiissn5D6dIcT9fEmh8CWSZWlF7QjdTVx7gD0
Aucs53BZMH4gTSXq5BYKj/NtAwm6JuHeX8zNNzBnUHi0D3j1jIwGT1QawyBZ6tNj
PnE4I+HWj/pKygG5kshdTCQc5KQxbYIiTQoLUnnjDRgm880deuSYOlsbC4eD15x1
LYJQlc2wUpUL6g4x525Z4+AW9vvOxycy1Wy0u/WKnoun0wY0cGEFrluXJEeyJJD7
h3JJ8JVfS9KOJFzXqhxEX2EUPCdf4p8H9UwtF5g2QxJjgMR0gY9EgGgDu7/CY53e
C+7Uk8DBUbH+mkp7GQ4Hmuxt5G9eg3BMb02c7Rb0UMUXJ3mnOfYBo8QgOP/+wjxr
YeeVYbReyZwMzwwOPTRwPbHOdrY1eRqOHyImemk2LmqpFFqE31gMRXBk/9RK2/2T
+S8fpPyqQphPgHkJ7PB6yOfsCu4l0TmdFKGOJZ+Z6W0zpIQMq+YpJs4IsZa4aDHN
ux+CiSI/bnj0WdjwQt7Hc6MmH8F1G+Lw3LzB2Qf01cG8V7tiKUlT32lmM5Ux/yjH
atn5fL2xS+2qF63U9rQ0AjpKNfPsbM1dz+MbYdWmj6b0g1sm8j7FLDV9zvLIyNfs
RY59XDfnN2hjTsRY4lbHajY3/8AOuHXnXzPLAo7Dq0J77TwQyNkxr3cVeMVIZSDI
aPvrYuXnXLK5JIaMZtd+RlDTH1Edw3BkcmElTi4tXoRB7p0fPcy5IxCVDmp9uRE0
JgeLb3J4xwQFGi/dkg71ksd3TIBDzClE0mXQdTDhWPKE+FxVo5ekubVR68U+MXJl
kGIEinLvdOxDZIo24rGQUjqcqelk1Ig2Uhe8HevjbH3KrGpLtZDp/BxznlFZ3lTt
Aixv2Dq9XFrRC+q4kl7U1Nuj54BMziVeFpp75o2/PafxKyCycgORYCxNx636CeO0
qptGc2sbCVGPNXlUM0l7ttKwoxfv5C/ZpGIrhhP1AvZrpINHMrwRYB/YpD8SXt7D
pbLFhOfbMhYpcvd9X7maBZTeYMllpkCxoj8Yl0ZN7SxwVhMB0uFnjheHEfqPRrzv
VT+YaZd29tf2JMPusZBcPGYgZQ7ZJwA+cJTgYMBQPGv1e4VzQVMo0a9jVyby7NS+
feRU9yHR8uUoG6+GqQ/1sFqgagSSoqMWBo6phzp1g0TxpK/mGr6UMBO2IiRuVW/F
3/GzzCpDWydPqlPf6pjPFMRPwPX9LPMeoHer68qlkYvZJ8ZO0IjCNhIYAur5FZsY
Tg0w7fq4ZChb2f2iimiBS3cP6y05H7fFMhuoKmOVJNx3O0B0mYBAygj0bKOinO7b
G6EOddiQyVRfrvhKwuA2UBpYf6KRoWhccZQSotzAB85MTlDZarrgG0wRndSdR2by
tLu8fDMOQQtCN8MgtMT0eHbhp0KS2BQZQmCnzA7ZGx4S7zrbc68fbHJ10ZBRzL7N
fxmUWXlD9CjBZKctl6ewWL4y/1gKpilv2FLwrPeI63HN+gIBzmcD6P7iDUkCGTwh
m3iP31mhadz9gWFv59t8rmF/X+aWcgwNiXPJpTsqAEOLcdk2djMgSh+N3ZRQtuzX
vTTyzRZZCcZCaMCUv4IVdWWF+w/rf7GQmb4rYDh0mcGCv5DEbfCCIv7ooq/mw2jy
LbMm/euVTzTGZMOB4gRi99ZOV4qEmlNrlbNd2N+fxht3eUBlBL5UQnw3XZa9+Wz0
5cWREA/Q1laIUFW2CTa5WCLXrWj2hn7Hnx4RUOAzcfXcdFZrLxQf6cZShYnwk7oY
ULdQzydSBQELjYBFRGtFdjcDhr9W+J8IQ3PxKU/obArxPRR1cAfW0qth7KbmE+jg
LXLUrRxI9CqYdOE0GJSz5T47YkoHYPz13vP1LH8bFSSMRbFlH9owdtagqweipZKT
sBeV5cB8J8vQ5q9DvusVMj9fb1VCL89n03GAdQTJSHmygSLy+QAtWYC1TNfwEmDR
CY6Clqav89c8ktAZ6dT08EtUMxBz+5GAvig0Y5gxyxfJvviNB2ZDHRpoQfTPyO1I
dG2V8L1/XnzPpBaDb+f/lp4gC7UeWW7Atx6ptaqmN+8Ye8CxnwqPrGrxrsytoufJ
aLdnOVu6VX4bCJ0pVUMDz1hQPxJJXhllKQb7lP7Wq2AhFVaM06XHO0d9nuaGocOw
1+Cj/C8BLUX5A4ym92JvAg1rWC/r/zNmffti+2zYrj5La+9cT0LyctCKgQwk2BeF
gAL+erBY3m2l02Y90sZH1hkTGfEI94gqBxRwLb5F8hPuTZh5EkqhmZFail00t1FD
AHZz2EXxzPj/uM3v2vwuJ6E4hAyZV7V9gVa+nAIyPvqI33/qcwXWg7vlJXLCwjFK
XNtpy20yEA4R2RxKCMBgil4yfpVGh+kEenuTpz5ePj4D2uvdbe9jNtwcYNySWl86
I/Ubn6LkmNGNqnp2SW61q4FT38QNAx7zxQcVr+YNoVXPy+LSYg1Dpm84tI9WWqA3
VerPlKF+wFC6tqLDfEJ5XP27v1iyyujLEbiWxmkcDUCAtxEEdUIpI52H0RsSkGdn
xGfKFIOlyBoZDWAuKKyh5LXSreXkMUlaV8Agge5NGpdLaLhfP2c1+UpUp5spQobY
Ev3T2ZoOgCoMqdvRjyVU+7/q5eiQo8lIcH6J6UeTnmswmVsdBHqB/coPv9SY5KYb
cAKiK9D4JySCqn++7JC2OV/k19yPX+lKp2ATRAJwpY/zYCGkGG3bD6EcGLNPasyK
S7R+fgBQBFiNY5qT/5frckyQJWQkPtU1I21XIMR/wYmM/5Zj9vBrGeCZl3i6rN9g
2jwRZseN6WBwkQZWAz5SngxK/E8+d8kZBLyrAXH12uotfH2wsG9xMy+s5U+etnOn
wBHqNh6pq9Is2qKLmuMBouYhem6KMCma0lLnaLqhr67JRtrfg9JVq/mSmbKXEc8K
EZhLkE2NykAnwO8K21IgeEjwhEZ5lBJIhxRwslHCjM6QcLDywVqmerYFJS3Km3cf
qez1czim7VlPmJiqieSNdKO5PqAjWgJrkKrkPkYd8ALtc6QcnIOyaR3pNVZc94ZQ
KLjoYOuvAaimTuQ1ZzaCZUugX87P87SrH9uQPk5oGlnquIlEHhSIGqPvxA1WQscU
imU/ybYCJ+Kt2kPQ/FD5QjtXBGKaPD298mU7WDdPTCwhizClzWjdRA1FMGRREaiG
yDYeAwzy8w0RmMViBbhvKG8NRziTXrd9AEGuZbIjffFQnRsFRUfRP6QN5cs+/WaU
tzuH4YuFWU059MfD12bne6BH4bNworGZ8900UrVhiRiBkIp+Ci0L06az78S6QqRA
ecsoGG+DzI8C/4+h1raSqN95n1xvkmmh8CxGbWrX7mg56wtbZqeqdTPX7/XarEDN
wrbCsGwF9pFA9QzKnrKqi84t0HDC4yAzBr3irKt8WjpOfVC7zjDRMsacrSaL++X0
tOJVpBqUOibV9RDzohuMM2F6Xjo/sLvC0FanRUJHNGXaK9pTuxcMiByIfW3A6aCN
zBSOQXAArHwie30gwLcp0WR4ayIqBYS+0ZTvv/5bTdZuYT2Wd7Mq6Wo0rhdo31/X
9mpeX0N3YVOnNmAn6HpZKOUpys16vJ1NExTbigcC5xOsK30eZuaNbiGt409yh89M
ZK+TpwsmQHtzlum3Z4kPlnoK0Ak/7zsmhfg1CUieVFDBnWkI9hCECzPanRwBQF6m
N9EFEOpFodyy5WtfvaKEkVWds63Yr2LSif3Mjmf5SwedurlmxmtgvsjhnXgrXs/1
mKOyvtmcfeD+vU2GQhlBuuJJ/EqNINMuKc+yHz/oct0lpr77DiyR3cJteDDMofSF
euiMVAlPOrjoEmFqFMCYBA5QcVrtXrSG3AWlnJFXHCI21beffnUp794qQGXaq6qp
g6FmipPPnp/IBBZADTfF/oD5pjmB9hSmhb3djzf7KBZfeD3B4nZ8wxjCbjahgX5j
O7RGLshohW52knCkhycyfvGFTb/YqtYyif18fQlVQ8WxikiiUQGgVzwt6nKEW40+
2XmihiNaOhQLOq2xfk1MgqHr5aqhHqjl8iYjq7sSNN2pTssd/4e4RWrhJ0qPsROK
AMwtRuIbuptgdWHuT2gwA6eqnpUnev5MaLLJfNTOoMgDeruhkh/2jAFZpyLDVHEs
C0bP+cffFOF3Z6tJq1zrQe4VoEBA8mJiQqvGNYna7MTUjx/pE1BdwZBtENie1jTq
u1PkLaIGEaIUMfwl1BYslUHyZjcJhaNeA9aYltiyEwygTCSVzn1T7HDjIZh0yByt
Aahn9Qc0RrWPJsal6IPtI6+B7rE61kHo6Jn98f7wGF3X8RUFJSyjX3WrcJ1rYSSF
vfUTpQc7zxsAb7Xp7yUZ/kT0RI4R4pUiHI4aTtaleeo2oFqgEwCizLEW7recmNCE
Cr6CfJVNp9b1SgP9BJQ523gxFzAJJcGkilTnczVJkStapSbV7biE19XeiSTUbYwS
h3g99DqmImD5WQGnguQeE7aGFv7wU+dnGgX3y0taTZ//9uNW8aRB1polpH2k1R9S
cuLkjIeMF+wRz2nLXy4ZkAVXBWfCAUQDT9oDTSfUF6Y0VKPDUio6Ga7Lsn9PPLkN
rlHySnYMzGjnqIj6auh7G/Oxhed3gJGicYnc9mrrVDrFFFNIk1RQ4sMiAZDln+LO
OLTSzRGfuu7WZIxebPDDgFO3Jx5YX1QxJRJnhaN6ptLj6nnmCsP2+gqJw5xSUNug
TvqJozKYaRO/cN9EGRRzcpIcCT2y2nwGww+7cbFfI362IDj8oRJO7WM4rMGVtMoG
gioQlMJdmOyJ9UYuHSHJpackFY4Qf4nxWeFgtcjK0zdGwDtIR6oqibqfxjWjflcp
AOy+O77l3qS9NXZALgofiTPLXoebfz9rPTLvUHOgnf2YH0fBN3nGDBIA2WApKNms
eQMEjVGcdq8uMeB2abU8bOtTyq91MY8AJT1wqiffHOtnaJfzZceswV6jmfJzEvI+
yQE2H2ZsHlMb3ObKDsSBV/DtLD8y820SNwA2ZFkN9vQ2/oUMyfEY1Q3zzBU2uQPt
bZjCsL/SCBE6ETVVnSMjGK7Nt/qGSv3QmtOhj7CXn4l2DpDQYdtw++RKAeEu8wqV
1uxrPkDUH4+C8SIo9OlmA3rUsMIeMKmF/uHYIFgCMZJWJcilZdmnyF01Sh+IShj0
Najd4eOA3cV22OY6MbpHoBF/fZ0VHy1f7Cj5xkWoH+BVwbI9gu1eZUk0To4SEyrY
akLoFftuUoRUwDRzkR+Breup8Q00kzO8BB5trhchLLZC127Kz1lSrujYkmEdQXx4
v+wa17wdFnEcyLU4euMA/z/VRxv/Z4hpKTsZxEjRNQ9PNpMtnUxEtu4Hsq9/lmb/
6PlH+ROBWkp/Row3HjiRhxCIZkFPXaoSzLXJHnJmgmoZnT+lgLO2KPaPogh3Zqtz
o72MyEUPNBM2Qlz2ChGzDND4M+7xTebOhcfbtdKoQRpwoCdfgo+Eqc1qYGPXxNfQ
sTTHVYEDDwf+HXShIhcunAcOHfoU8bvSlOK9VszKJo/2nR6d+udn2ul7C6fC3ujY
f8cxs9Dxgud6eiQw72fQq3ok5l5PoQ/hBBxWUvYZBwyClB5ZthVTcqBGMDUelA6m
OoxlauL1IOHNGxqTlPN3zKzUahFdni+WRw1ECDS+YbJE599S9Vck3E3ZaHHFLVIP
aNzxS4JYTcoxXHvkip++TdCWcGtzQ9L8478Ixr1ZSpaRJSMuaKyXCLM3Pd8PcQJL
J9U5w/O1+EA50EduE44qJNlAgCqyH8qSOKtgo0lnCsz7vESzalKxb5MwnegO1ezi
Q2/0tj2gPiiRg5xv3HHAUt4gnmaRdHF3cR845WPHK8SYwK5EKAgOL3FT6kD6o6M7
lDO7hEmX753WR6iaWG0akwZMHTuq76GlSTWDLN7mdrBH7e4IRRwnFlEsq7lmMVhb
wqtGTk3EGwnuyJPRDkjl+xX6dXiNgvjzFb9fGEkGyXeIMc3hiYVjTOi2sPqKnn+a
oslt0RUHdkP+IwRk9C6Lt0X1CZR7rPnUie9CqAHivolaUXD0n9/zZGEeriI9xHr4
/NivHAectC987VoT6fRbcDZjRFZ/EPiADnwuLjeR1vAd3B6G595bcUhKvdCFlLVt
cfQzxyz28hsgO8DD0vHEm2Pb+/I1binEiXAm31eiwJ34hG92Xa1wWrb9+xeLp97i
PcoeRZ6X9Bo4zfDTsB0+pzUUUWwloXJfoFDOK1fftYKyhvDGdoiyoeo+lhoZT9Xt
0tfDuE0IGRNMFCdyyPkqOQLzHcceJZu6Z7xYs1tWUeNd/kPsZ/0sHFslmzM6JBC6
ESHKAHUoWBImpsvj3dnv6mw1FajziQHT01qnVaCrAPWmQBnCc13jnGALAY2J5ze8
El7QvcCyeNGli7Mg1uiJWhP0oUMEW+kKCoaUmS5qS9WUWi/9gGOaRbEpnAm4Arin
NSZOUhTb+JjzBMH/kzKyqGdLxgeG9F2PefPQHA+ql+YzbcQj3IrSMC8pmMtXwk2t
5NSoff4/jfzUUCa/11qKRHtat8/uMTLJwxE6O0b8ye7vhg5SYjv2NMnsec4Y4C0Z
jqdndVMMj/lV6JRHgibijsqlvo/TQsdn3Ghc23TDuM+NrMxOeI/RMdkfZ4vY52I6
jzCQtfYK+DIzSOWEw7uD/7CNQZ0zg38L084VqAbGUv3ujdOF+ie2feDEJMzWNC4X
U9bwaIQJDqLY4wQ11oHc8CW0mGbSS/6ZJnDFdSlQGKadngyUIz422dSbPWtm9wcR
4mdUYm0LoKkPPaExG4ZzqDRO5PtcKDG0E0m10S35vTDF8zCfkMd07p279s5+2WJT
H/OF0BSHGZZucb3VGYcldHbq2TedKSx39AWomM2FPlnL8ZcKQv3Ozc1yrCBMdwx/
UG6qP5XHqUZZ7bBzMCcfgZUI1KOuvi/htorZsWAYGfvk+MQgJLPcIao4JWMxFNlt
du6dQegebEWpdXu7PQEKGi7ekvSWpHDL/7ztEUHCVQe3ei3qtGdBtky/YZDf5IEv
t7kf3Xo9BnNFPK+bLYzqvBxPX5I+uAjMYR1SqfKV91H5Y5PLqbV4pjx7W2vTR+Vd
XnMp3Wp1MaPm70FCYcdD/78CRvJMyJ7tvwkyVbVR4fp6jHfwFSdBLiDSjzb8N6yx
w1lqd8WgIEor03gvz36tQt3dTsrfqV2Vsv+V2sgYzsHk67EkR2hjwB2AMGf7PsTa
wca55ZX0lhyeOkn1N/p8yAhsXTsEnFLstdLFOitpKg6HSZNsoks7xSn3eetlML1K
vefGgbkD758cOisVqIN8hOKg90BlqxdvsnhhzzY1PxZTRocwd/Heo8UgmkebwzWz
N2ocn2WH4kxAn7hqHPL65rbwQ/ky6MIj+ugLOy0SZv9s1Th6TiG5/s9eSWLYt6Qo
UffFmuYks/5KXeKKjvZOB6h2gqoVpMjfj97ZTc6CtI2DmvKB4ldzhZqa7UgTMt6Q
yE9AouF/A9E/8VZiEWTOOX8qTf9qLVQ/tODHIhqoEtsY2lbMsLoprWw4Tp7qKhyV
r0A4WLkBQMHSBPJ9K2ObaWyNxRS/8CDJeDBpN5iSpp4WAm7KMWS9lr1+cVymnaaF
MSKA2xlxkdz72hvo0s+h6zH+/JbkuIvCLsRjm4F6x/r8X5DCAt3GecHoFrtJJUhG
RM7/invD58x4uwAxPH5IwA3/54J6rUMHYE/f/Wfqcd++66ASbCJwG8xvcFTTqWER
a68BsTOBC24WSexw3ru7iLay0wtSxbxrM849cP3lwKZAa+T9H5a/F7nv9cBiOrmC
iykoUiUXjO7CtFzbXqv9AIXSmnolSFziWqFH1i4Qf7bSiNEHNvdQ9pw9lG4Pn8ej
mAKRkgqn7OLq+zWZOpRLOezVCW07gfwwARHe7uXIMVTNhe4SVr7b6KobmBAdEz0s
/6nwCItgeD77Vlenm7NnXPNhjOtOQvo1UA8ry7EzlTcMgve4KTK3K1ofgMG1Qc3K
gvPHl2xEJxC+ydui2SFC/xrl35uAHzNe2mKLOmOUTJmKgs8YENSeBUKuj3zDrCf7
+8q0/0PUWrvXjxWwsPxJD4J0bmBUwFsHYj1IWyZRQCQKpuDqyLY1LzChNOzieEw1
dKzrfsSc5ehuL+5BoE14TG6Zh6qjA9Ysl2+4Nuxfi1jK0KaMiqvMMoXfm/gJmcQf
09S4bALLiKGeyX1GtI4qcVQlgDddUjdIi1r+dzYsr77c4GDiGfFvgpvmdduPmer4
c6xgnIHMfrT0L57J6E84H7Kd3yS8CWAuqjpIGTC6ntXgvYb88D4mFvUMp3jAUkXm
Yugug3ppTrgoCPSo4XJGVInstd7GyCXqmzewuDYcxZDHx8ii8HtLQ+0A1V9W4PRW
Q6mPY9/kvGeafLoQqt4E5sH5BY4N5IJG5BL4kDPZSwfrsT7sjZXkTIiM9xv8/hE1
5uKEGQcpqX3tpBQjddGX7jGr5yr5ME4rBLoEbYe461bjJko11J2jLXvxpXZB+usv
4pnSC3VH6OdUZTO1nq4BNlTSxn84odJm+AqbwAsvhCaVl2noK5ZPLKw11Li5T4b0
ovz1iKnBuZrjStMMGTz30Z4LWReYXO5RBOt3VXDMRtkd6UvnAEzg5DyfZZqtKy4O
o4bb+fLf62TtByeRBsTAjdZZYD0vpSTFv/UXg40njTfrb0t6jw5gc9RScLj1S3Cv
vlfx4l+zQ5x0AM8k4wCLgHlkSr3YbJ3uGKB2y1XD+40IpSsEGEqu7GW1uKUFzR8A
DcbEde6+RhgOkv7Ya14jntCE1qCcn8T+ZfpjkJfs5LWduNgvLddRkDP9MqUu7Ztq
xpxOKcUzsx3vlMrg+sD6cnoVAJbQgv5/qTUAX674nbtgPaf4qf/vi0w0qPwiAkRB
Snem98MiZA57oMJ+aXkSbzriLUQWAI8hav0SpQKRGJ1nYUZ2s8qedHIV3EinacPP
giHpTAHSp5Mb6aoGKJFnfcR9HwZvDJTq1gasechcrZrm9HIaqkVWSrruvNhtMQlZ
/IeVYa6/KLEQGsXN9SD2mImSKxih92PT2Gps+LdNtIWQrf8qwwuZ/JszG48WJi1+
rCiKLp2qVW9/fUB3e3RMZArRoCkGRKktdKlXNMvIlfepByiZF5JC0F6UPLSy+Eak
+9xIgKT9HUsvBJ8flX0dAuNyMIN5DVLoX+GGuy/Q28oxJ6sZzazXg4bTNnkMp+iY
1rIESaNE3Cp69dTxaab28raqFyYtbkVO5NTQxMamOLTcuYOM+vgz32DYhgYNCR1s
zdwvWw0+t7Hw2SNNmfItUf8MeJA8FxQDdsqDlSuPTx/innrm4PR1h8Q06Bn+yVsk
JVzii+1etdA8gmZouauw0daucKn4YP9j0evKzUyEfqV4Gmkg6DfYap9JPsRCPE/O
nJy/8LT1XVwu5e10vHFWB/EtP7PHYo75CzJBdfJn+9/lQWwtSboxYR59tB/+NvpK
ydaI5jTLJZrCnCPolS3xzR3WP3OibZ1x5dcpYGeZUod4LxmJVouic81E9Z+Szw9G
BK45OGOPuXGoUKK+KbINFOvKEK1jTdatFueSu3z3hclzsu/BIsdZqUo+LyAIpidF
qIUvuL6UcS4M/A8RkQptHYW+N+u/Hrb15mSj8Eu7uc17G8Q/I80zNonaRv9RSV6P
F+VNm/he9Om5LCLwKwNEnoXCpMCfT2BVhnMK3+0MLskFsI0TY5rNx/qPQ/VBrmug
V2Lt76tWQhgXn9bz82GfYujai2luwwylSBex4Chc5EMxbEammbU2+qKA5fGQsVRp
X7AUnvrYeOW7fbsqR52ytklROOZ7ESkq4GhF4lBUBus4pem/A3jigfmk+zX/3WRs
SGUvDWIzXfQNq2H9Tmo96hE6C88EW54MJuuLwzYQfXloRhHRHMnqQ7MZoIs8esiA
6CEUwgsNeBnin9RSPYsy70LZ9riE09F5kY7QV0DLyH17LoD44UuKmnGSn7VI5+KW
De1WWr+dFLXW9Bhe2dnNjgX6Lz8vw5eEKKslgxzGil3WQrYewnlbeQ3cdM/5Z2h4
kvCSYSwfL4LYJPfeQfJKHJPXxE9boJUgQx9pzUgbLfETq9opQ9JwBMIu911CvuQu
jXDulXT2NyT53SOs267U6tUXPWKoxihfexRpTH8anxvmS+FaWgYd6kVQlW/FQrDG
8y02I1eu7FqdAjITdWAGEPbaeWSCks1shX2uboTBHPq50P0DQ2OhZexoUhghDzHk
9ZMq8vzPvbZdbwD4z+JG/aPOWq/+DagwMUgeItlWsB9h9Mm/2sZrIFYzLnQumjFP
no16V8Wd+cbrnI5/F0ZCZS75cyllfRKYY/H6m4+nW1zkwx0XH9ydDh+XlQKB+8Iu
YrXmvZVjqfk9xqQCkpisiY9Rxzj1WemkDwMZK2HEt3G36u5yhPGuBUdura4AzgEm
OoMbC1cQN7tvcDuogYh5idkdIE7Dv5cYyfHOD92qNJbKyKAsyIPnaXuGO5rTVQFp
fTqf7e3zEPYxxb+m84JkxQIGn0fyPJWYsezFfwVr/Rzppx8Jf1m8fF/38mFPqj5T
1uJS0a5DyYlN3pwafK+3lR91tBq3I4rNak4EUy7h92YzAFpZnQTocawQEZAfwsBr
Vlfgh/GPZIa+R3GBa5qg2fT+M4WS16GO137pw2F+HulKsEvn74b14AHuPlSfVBlN
8nmajWVlkuk132c4pgNSt+UHslhUYiPC6CVXeFg29oG+lduYzcyKUpfSKEQCyiwO
psBN1OqAdAm410LRA2tvVIH+OMtiSAkKcnawWXsFy2KCSGlharXip9yuEnSKONH4
pj5ARly1vf4QfX+sJ29F+oem740KdJFGfNQduvq7oc98yYPR6Tm04/gT2N9oo9+I
YwAMQrcylN85AQLBhyC6mMNoXffnrrHyUGDv6h1qDz9jm6E1zJJKlika9+k86xIr
MpSWzQ1QmHBKO/n1veHkuQ==

`pragma protect end_protected
