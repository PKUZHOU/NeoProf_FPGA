// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
sXK7x9SkqIcobUdwDy5MfkcQBHTvKpo0vgFfSb9fzRsDEi851sX1YcZG0xMGJfPI
6PECJHPaqk+AXcPun4izFTkTnggT7AhnK2k+k/FAw3vudqZu/WDiq/pr+ymRSw4e
JvHthVrJB++Eppx7R4soGzLi33dubBE7nadamRdrCzo=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 27536 )
`pragma protect data_block
tvNAgenaY81PS4sPjeXpK6iipIvzhlYwrK3OFbr+7eDyLF0r9OJdhkZrUSlPnSAM
xtFIITbLPvssCG392zr7kf0XI6x4yuQNC5DT5nZL+Ux0aOMN422uUUnBkxk2Jxtk
1Q94VORu+5cFFEO6H7+Q4Q4THJ2frisQE+igaVyDzlKroFKqZKPsSYVKGZ11/5rF
DavMfA3VSt1Ko9Jf+ceJjiyWk8JICeRQrWhGL5mNbz0Q/pCxdWOCE41EugWh+W/e
N3xsSPjy84PzFqsDQl1aBOmoq5WSe5vUcv6txinDb7FX9VLE7DNr22nWHmRwHoVv
/nt+4FkEOrIWATyKoxmHsr+dusDgvK27GnS4/7z6YpCk2zgEiekLrz0YHJAv8Dlb
YWrIui3ENr8Rg4Qht4BHAFXKLtl/QnMyFk64iRxzR7ADCP+YRr9XedEiZMAme+Uy
9xH1FJ46toyQELd+GxNIEf5wtp4Gn+2YfzJskNQVLxLjspoT8341cS0cyTsJinGI
3qQUGHIk0Tn31QsGmAu0CX8P0uU02krP7WJ72TaVa4r7pzxrMxRRq1tZTvv9sPL9
ZsMcyQ9iLggBSrJQdnrsYJKZH/pLRy+sfrEmhcAPcJvY9W+6gw5vKyiE/ER4hqur
pnxSJUMSvPpXaV5T76RXsbjPHiaC6v2iBTTF8bvbmt1CFiyPgFzHCU9FqLzBWcQ6
L9QXaRNKx7x0h4luvMJQR1Qsqo/mBWAHi93e1/+ecOqCnucCJwFaCBNU0oTMLUqB
VVrNlpplGuFHoj8RYOX8rI6oQhawLVF06FHw3A+YyQKcEuR+Cd7aHts64btX6x4x
5X6pkPm+CDoLv2Y36G7DPBBjsXznaq2Jaqf4dMgvqhtRgsonVwCePBu0lk4WqQOt
DKKnXHbSIgrtOesg/VllHhYk+kL0Fh3TOS94FAGE8NMei67Fq/Tlmhi3gvkKdWO/
5GxdtongVuJE62mcvnA8Qng2ri9qZFmj8qp6vKA5H9YVTCWYaCyiFIc5rbxjZ/kD
EFmUcCh/07Oqcy3Aho4nh3LBwfwy10XO1QYeYwMLdWDwVVNpJCb1pMshtRWfmpcu
Nf/2vsJBvQvcfMXllRutpxEnSkJEi7sUi79/i92ScSTm6YGUqwo8+PKDhHFYMlMJ
UgGqbEsug7bOqmjBLihoggWd6K5X4yjHuyOwsJ7rPv//iJaxAfanzo8Sshgs2+63
iIMbbtPDBB91nlVKYDBoslih6j8nV//cp1FOVNcYroTjn1bzg/wexfuyX2V/W7SY
3CboGy7aXefqXFMU5wxTNOb6QAdpvQFTDfPkdtvfug7JrvIWPZEQ9jxztawHmDZw
kxx03EPBNOKb/v1WTlLIr6YcM6iwEogD5liteutGHWuE4WCQQZE/UG8tTIBlQQ4d
QtxvaUt1+8P0gDuEJzmFBWHZ30He1tTUpdwEAevK3PaBxSCI38lz/Bji+NSrbsmG
cixxZRiMuaMD0cJjfqWSppciH2HWNpLPW/nvH5CKIUpbE9UelG5FrR1GKMIISK8c
gr3FoZRKFxmP9Tt2t0/CCxPSceQVJk9uUA/C1lF6YcEWXecErbydmJjJElNrSOTm
by+PcNF5MhA5QleRsmu8bHNLkD1Y3cCYfTVOgbS6v4V05dnQO0rWa3qbWHmNyi0z
evVEB6gWqlQXRjUeBFSQLR3nrk/LkKfqKRR7kjMpm9cTHAyH3cnduCLmN0CDAgGl
Q1lThgUTCV55aAh87vlZIkT1nSfz+lhsiiWtc1ThZP/Cp7ZE3+f7l20kizH4wiZf
7j8kuz7nTRAhc1jKLDjfeL8skCeviUg/hjUWFVR4e9ZixfA06HBImgskxokI6CRI
LEmWQ8Vfc3Yrwyod1TvTdvq3HcCHOve6i3+Tizh8t2HEeNtAXA+Ewp5PJRiGMwyI
BHeyzvDFvx2X1WolEp5efYAWgmbwSfFKmR/KR8ubeAg4lM1mJRz90VB0G6E3qb32
dtLgg5f1spex4lvmlb71E4jDmSmZMQ0RR52InGHmxPowVKKSL9NgzaOzTQVupeFe
vgqhbNRd1C3jGaXTAZ4v1aEZUpuhrwbYRW5MDLC3JdH0e3LDznjbO2Sh9l0SJB8Y
N0kNdObjVT1CVnteSCPHdPH4a3sPVCVTGcKP1ZM1uXbRmKZDwCoTo9+oSGYrlIMP
+rCmTMwbLtR5RixmZhfIiwJUbNRKcYkdGVTDSHJwa3HXDLUX2KKreZO1mkDJlr+q
XdwgI4IrOi+YevQI13T8LOOmR0Ag39T5So9a0KV8beIq5Fr+74moIh+Iszq3aJEx
UZmpLZQMpH5flLQNkD3si+sT7DnfEQU98lIaxjT6gfUfK/nunydbhUNqoFkOMoTo
SMDfSvae1vpFmnGHuPCFS9iYup3p5Yqs2Dzv7m/lUvVY4kf+5YP7uSr0RsaKb6BN
7c+CryA1ybod0s2a0RLaFATQ1JhQa/CSVCGAH6bWWqY7SA+xf5f8itBGGo1dOHfx
dHuFy6hnuAxGT6PjHAL4F1EEYh04sjhHe0FYRuxtIzvJtkn+MP9/uyvDHBE85AF9
X6VcjOha4FDU+pT8+o2Wsx1kCOMfnxmBeycLeJQlLFd7Ps/N+IO3dzZgRNHQcMB4
IcfshRFP/lKO1WS5DH55QmBQWRG51WM2Eo70e35CzxgGfuTBEPr5FVXkQbGMKySO
WDeciH2eEGrnVvNnlnP+u0//N5Rs5urR4YY30Zf2lkO2MwTgDSQpakRyyc55WOto
4ghWbpx6SBGEeyVCJbsuECKkfcv51VFIzB2LtWsDBesMDa6mFZz7QiTbDgL8BF3X
u7mmC7pRAbEdTaQ2pGxrAJTsWHWvV4Fqap1YyCO/hUo3zH6in8Fa5HHIEtzFn49V
Z8Ra6IY+Dk50s2epJ7+gsDc7nZz6zZynRfL4p1oAWgFYVLt3JNEsoKKbDNGa8PFD
ja8zY6mTJWKGdzx+R5DLJX08lvwSBX/jUiY5iAa94ZpfuGcf+N1HIHn/2CE8O8ul
5bkUU5PMfcD/2PYyAoeLozdE416d/AHQeFoDdZlezhh8eXbKnfpxjzRYpVVoT4mS
cF5FpPL6XDOFBwZJKOzbMiq3JNAS/Ji0VDsM3mjqBilmfH7SsI1rAFq0YmCmwQFY
PS0VGVc8925RuFehyANOvV/GP5/Jm5AyBSBIdd78DCJzhM32CyyxxfWaFa4huhSt
K0xnsp++DWm1pB6WJuV0uNcfkxO7PfgPBcIH3JGYhwhX4vQ5FzhkCKL6KYLN8dLr
HgnhgbRA26tlpcS7yTJLg2cNoRtaZH8z3puDEC7GaeEvLTFFGdf/dLA8V8NyR7LP
wBYlMRPLKZHg4ragwARO+6qCRx1YqXWdcQ+xr0pXbYz+AKGWJCkYZtnogkpbkL2q
zqdNViHjw1s+AZvXV6bXeshu3ei7AJ7AEoZNZJx1JExrnW29XChoS+HFaWpiJq2e
9df2IKYCNZF//77/MlVlq4IcEAxNvP9XxBa4k7euay6bnC9fuml+M6NWwNdmpDJ7
+4a60KS0Lki04D76Bp3rteyDfTV6Nmzu8Qvs9r9vkBAhUXVtG9qqu5VeF9zRgwRl
TWNvYi9M9jjkP21ujWJJ/Ga77c7Nu7C1q56ftC3/UCKvz7rTuEG8OhI3WGIpl8Yz
FK61XAIsRytl8LlfPUSfqy2/5GXizGvSBJwvXFeed6PVmbQHfxguYqCZ0sQHyvV1
HbA4aqLdWjIRImIrY1d5rhaZztplfBRDvVvQnrAIl7S2lw/W52wUv1jUyixEUZ0H
Ik7O/Winmv7U0vOoJqGYZZznPxPTitU7okNSCrKbgv6ALG+ZU5LJdpmT/bNOInEV
pO3q6XV2W0TCUcvsuZ1undh1YYAL1K6WAE4EZuxHkHdM8z3fYbStFRNEuRApA8qV
92hqxmOActriTujeJK4AHROL85ReYScbog5PjmEg2UP/mRxYuBKo58JlUdC0q/rz
SE5tnFhIVJZr9XqvSdngYQ8L4RW7pg5VcOQhmIJSuwPJDnhCGzIFA6qpjXxPsSc2
UpIhkCOF/0KeCnNWQEznqQt1LQrU/JmrUj/1Y4Zd7gLo2+Rrp1k/UHAcIUUwKmBt
5xifs2dxkWOvHa4EzTU7FXRj+SqzSR2v/Coqy5RBe4MYZb9YH87/wlDDyzI+TETh
y4jqo+WRdQ7F45lGZNTTTzTxQ72KZeUOPotPFx3H4rrh1h9hEMrj2+a+gKvbnfC2
GP5p+8z86Lgh4Dn34de5OQDT9ZCUA+z1U3ow4Cg1DpeioVF/Sog1wodlRsdhFFVe
1rKPOdNC9V/vNzv4d7WvKnCPrQeJxx4fogo8kUIAZhO/dy90zdNqAdoiqreBzrUt
Syp7kMAW6NqNK5+OSiSJwghfPCRJISnVUVfAJe9W1gRwr7+bOSS4RGXOt0pAS/B+
aTT1anhrGtSvYXaDUbwn2oymhkDMwlEg6/MIgN+96/4Rw8qV6KLHapN8/1iR91mX
4Ikuax5ujjELSE5+Ux9jZ4iMpPfvgZuX9+wbry6lE5L+/ZuFLLUlj7WBmLrMvVA+
qq8AAxjNUN5uxjIPNMfBr2pVcwwQBkIQ1nyK+mHG//p9vvxkSaK/bqRHbtwE1vzw
bzfbUylMYNUCu16si5jXdh1im7EGiguo8F1OBn8f/EV4+Ui5LP6BzjlN93P0vd4J
8k/DTI4o4CPr4bp+fmWwqP80MTCigry4b6GBkLfNbEku5ulREROigngxtMPRWnN8
vCTF/ioB2jLL23yNgW2N/aJMCgUKxVTztBt8O599IPyejGXeNT0T0tqi1q4cWEUR
Yy/MN+83kU/Pv8qi7okmyqBw3jSDEZ93ocYh4q8gA/xPs+mpcT2A1rtvyAgxrepj
HJYYD4n8XMlggvYNtT3ESuc1EUqTzWapdWOprNyJozFNiBsekI/rjE8Oe595gtHq
fPLjz10+/vlE98UwT0C/PUFbhMG400SQmm9Eoa60YIZFEcUDk/ovOucSnObDS0u7
U2Mszi1g+pwP2HJPGofm1FCYcEKlvxgC8kLHi/Gs6oVetJmfZsW76zQzxphnyOK1
bAVR69tf9jftJ0hFb2PfjoQPFieS1A3beLXgq0sz26TBRSjCMuev1GTNkXLj+gj0
+iL1XLB2U1HSL7qk0niHfqccjro7hrAHiP2DPL+zQBiVi02kRvEUQft+ly//sin8
12vIEQ/JFf5IgiAD2KNWGw1dEvjeSwcPGcvmA5sB5e1MIsEUgRGoQO0M9YQx1STk
gsUUhFWC59cK9YumvdJ6O0tP4WUh7JOzXNd8RJNkHXRI0dvgtuY7QO+8RhyI6gLe
GpeFmldnJG4DEsPx0sqg9fpnIW5skR73mA0C7dR6ScAqksq5xya2gPNV3NZUy6JS
AGOUb0RBzqJJS2FnhI1v4eMuSBA4HB6Hh0tBZv4aviQDPahLl03pG/kIRLSjdCtk
6ZBr+zI35IW2Ph7VUjrfZnnksHlZDaSKUfoPqLvW5ltgr3XKxZwTCN+iff1GcPMy
AEdcA1SB2MksN7qzpc3qPZdn3yEuDrut+i5jQUvqf/GhQAWosBr1orNWAqQWEVCS
+N81ZkhhithOZkzo6gsBJvLK+Cpp5dnfQbSzd8tByiQQpD8ipv6255ra06/uq7GY
avBOv/KYbDx+ZvzngtfVMOFAK2LhlaNLqG7nzuK8B6MVN4/CsHsUCHNNbKW58QQB
LMC98TVggDeL/Fgh5Yd5IqhL+NJni+VdJo6wvk+E++RybDbEM244qtwJIbs74gVE
PrPBgFjhyV0b8qwVHMxdU/zaSwgb8sxoRJHMcyPAck8RZUZrKe1EAbHBXmCg/eRq
APCfdL4GaNH2RlR9wWMGeuWUViio2eMuAmhc9AjoXM33mtSpaA1j7X4w8hKjvO/7
ztVbbqxSv1J7uz7wXms+MirG+el6BqqxVJ8Jdfd+vue4aGPLW52OzjCnzT2tn/bY
2PwB1KJgQx49cBximtFpoov/tHFWqu5cUDC2nPDRq6PeWb5+Qbeokzbea2OLdnC5
8dki1tSJVLS1VknaIOwuSmLqb96dKPCFqJ9xfa+zDfRR+XhZEcjcX09nJ2YMCUKc
5UsDdy0fck82R+ag2zKWd5n3pFYGHRzOdjlmhfL9Jc94UPJDSTWOUOwxUkH6xjqS
QnRK9kshGRmsDvEIwN3C8G8qRrMKbbHzPYEkgWbCfcQK9M2zICcPIeqqbf6mMO0q
pmNlhRhwxAUL6lqqXToxsqvoqCI6S7jzPjt5w3v2xi/KUfnVdTmtbBmmL73rUT+3
akefIHJKI5b+JZt/b6hwpejah+TnjK7uwAHDnzz1o8b72PF3wvpNtCCA2WbCv4X9
gb281hCwFyzvCti9xCY8z4g7XBmJnxYgnm6Na0r1yXzHLdmocs3EmH2Vqvs/W8gl
5R00GP1PXZMvZI6qGA2G/5d8U70g0OtflX86YaiQNnTuZF8PCr0rEBTrW5r3DgMP
RDPl3xKzDT4zuhJXRzw56+w4PpCVMfhH/uwnnwFCZ0DbKcqCcPPEAIrMMQsy1hh4
DHNK1d4juI4VI8wSeP+aUfMILqLKsqIxJoE5bOyDJlv123r+26Oe5JNPpaWLLZ6F
m5mvmVlkWy9vvBWbDV72ckK7tgt6XlDel7SH9Vvgs00hnp+tuTDIS+Cr2cSeuDHX
brNWpKxO/tadjoIgKXWJWnkGJ6r+JZdklTKEAmmWiR65klFbBruEEFOEapekky8F
5ZAMpFomkF1QqW8v0/NMjcQKlp6d80JJMq1zvDxk1CuybCIbePZQwhFlrITAo1fB
z678KCQb9OFIH98N2dBMR2IsKkZuHdmuELW7B4UW4GD7QCD74siXx3leCiA5o2kW
JWwtA/8W0FYCZwwHvYwFyypXlOR3H8XVPlHA/PZdfFcG5rxujAkieyWzA7X1irzF
zU1Ry3+s3E/R6fstRKw7qBooBpjLCMIY657jPEOJaGarV8PR1JgCCtTckJWfnPRs
1hJbrFB0M0Pg5uSipL02OjOaF3j41y8T2IKiQXeu865c10SO66SRo8yRR1e2ccWe
rtW2N26tSSeBkwMQ+9eGWWXlSp9Aa//UC2QAal3XHq6pTDMiOaT+sqsYrFIHX7s9
bKt+Ca7bpKnj3sg5Rs4vnriQXDHH0E2B6GrnbpM5hiqCkH6jZQLpFJcd9gb9BN9Z
W9iwhGihAh404xQVUXnGPAfokDF8vjtOQQJMY4TyW0EcJzZUhGjvVzR7f8+q72Fj
HADrrE+0zBFCO644w5md7Jlz+BZDfX6wyAsNtLF72nGlmpmnL+ayxVCFHcUDs10f
Mp5VN639WU7zS4PzKTGPNM11engred9WQohXQ+zeEPTjDP5xEssleo/exRcLgcHS
8LIJ0WVCGXCXPvXeFRJBqCt/DGE6ehoFzdQoGpEezw6WQfeWetW8lgG3nhPrajLi
yVwm3jOUgrqDrA3uvi9rIxDz38xvaN9CcFpVxluygsxmC/GXKe/kj1nseAQZwX9W
LZmv0xcdo6CiuW9q15qrTFnkzwS+5D1XI9pJchK3+EeiBexnHK9hph03dOuwUMu6
0IEKVQ1weE9NlOY7ydvatPYFihWM9x1GvjL7ot2svYTMnrFpc1xTPEcChkK5EcjV
gBROd8pPXQa+LQnwm8O4QH8UN7bG3+hRldi1CtMSkAJQ5Fncb+rD2XPBP2F8Y3jh
tLpWGXzbtxWIVjgsNSLyCSGYJHsIsTbU0DHAO0DRf5Lw/bK1gKoIsZBf74LR1Wyd
GZ+6BQraVwVnvzOK+bm5wqmY5y8ELv4cw/SYfiSGQdk9v1l6yZbR73FN1tgrzB0X
gRn8JMfCVP17B516jhERgizNW/4o2fBMPzKV5cmiu7hAn7kSrVYsEJmWGAn1X5nw
Tru+WHhBULzxPaKqspzmO8Gc+xTPfp7C+5CTlixpkEiJA5d9KmKcqQxjv4vCDlOc
G+aBClCRctN32dR9YupRc9s5hpi6kLaelATgOp8g3Vg0ojE3gC6ZEyQnRXOgZ1Z4
QH9OYKv10u2TTK/ZYSrhQ9ARcrpfw4KyPsZe63vxaiizbpWqc31jf1OwwElVuBcJ
hjUe9KjNgzkFo3sxAL9SeQMXMdto9v6lvNUMZnRKciiaYLuu+PhCBZzSesXJNNiS
NaHyiuyHwVhF0HN4A00qhzwcpLUlh8uK4ehb5PXfIBO+vyp1WUT87sSQAycBXyOL
CeaL4V+jRiBhhGPXOIyBA0+ziGBgktZlaP+Rj5kTGgoaQRbvymfeudfgIYW82/eG
2yc6BomAAmtF610j1sSaoHENg0naYD3a9a2laa+C8HJTERgdwfwpFz4GZxMO4KEX
ZmumG/ud1p9Mi2rUTYtdRG4juzcLaDFi5tfrYEK6twwf43o2tofcz31KArz9MeNE
eSEM4o7+24qQ30I7xLTXl5G/IUmYyt+w657HPvjmoeybl/VQ0TTTVkLPZqxoEP8m
U8OGcHwSi9O6B3fQ+97D1yb/LViD3oj9WDSHTHruFnTFUX0QW4y2gbMRRJZKmMXR
NIIkDDXl/WYcRgRbh1C7L2Hlh6Pn4B8L/BKzYbrD9WeOwyZ76eaWA72MVTVXMMcH
d4sOoZedZsn376hAkoTGJjkMHCoCG5T+1KUjahIF9XQ1tvbiA4hnf9fv8HdEHpNj
Py1zcBF+eb/fp2gkjbsgMxzp4RJWcNYilSUV/PL1InKd/aDXTNmxK1amczDSdB3V
d4ozJt2RdOgY8sNi4mCpQDYxrLBOWmvv9RbtZZi29egFwn3shvhw2jSQ4dCReAiA
nbz0evN77aE6vfu9OVBr5LrfmKDBJMFnJcd45hxrRVMA2bNxaPKkxLbLk9Kg4bKq
fKH+iNXVVPNYa65ud3zV1drwpeTpgAUvs2sML87taRZk0bL187jgjyK87Ti6Ufl9
NzFgt8Q1VFehLqTeeR/CIrgWA7RXL+ecoFdcyDuO8BawhQ3VGwyVQTvqQpI/Fp1a
63O04cGP+JY2YzwJPVnt+sCvwupnpxJ9UAkd/7uS8+pspkJ37pZFe0zL9hDCKP5R
mcWVTu5qnxn444VfA3RsGjwlyzVvehBzXe+fMnRuHw5zErv6OltZXQyqbKUicMqY
28UgeNNWhAsdwzT6ro41dM3MsBAwsajUEa2nakaGDEfiPfqO4cu2LPHeBSrj9SUP
ywhsF2T6FXTL040xcOscaqWN0aeLBFVW4Y6cgXQUQF5Kd37Cl+/DVmwgGRY2nWfI
02syAi0X6UWNzCr2AP0+qvY6b7km2Mx/kMHIrDAMTobT8Rm6ZAU/uirLFIWwMgT/
dedjO3S++vKFLaLGYlqa0YESRCwgE4LRwdMZEh7+tLU8FRFWm1Krp/+ok8aDn5FA
/+Dk3b+zialcGIYv7j9vsnwAcZA/O6v0icdOIbwg3oqBun7ym6NlG4RvzLryXV7l
RwHPCkMfnUywGZ2GTWn2YBsuOKMcVVtKkCUmH19y/zAFdXwV51LB2MAsCsXEannv
CgUY0Rzhmo43bEzMtR08uHkKGKPWuSaHor21t/DZLjfp0BKDviiEJ/pHMwTI6o11
V/6EQFwiTAyPt4Tox5srZ7X9LpWY2/4CbWi7CgRgcM5xe15tzd/0vg7YBL90S8kt
teag091aR8mrGHmIyokyAhNIuttd6m4oBQM9jRcvtJCCx0m+q+gndN4l2Xd9cp0/
tvdPExISTZ9dKOAy7/mBLs85qlgvc6V6Y35WQgsNXnAhZlqLQ2ZC/rTdTzv3d9ZD
x3kb11MuvdpTfhQWaBRqrBJ4JzYlckHkMsa0JxLx7CLpWWfzzXFp8wIYuvoPVcEk
2cll8j3QUEsSrXxWlf+jXj6iLbF3GZ2nnNeKOt0ybB5VZuY8ZTd7rpVe4ud4WKIA
5sOu/uATx7z/joboia34czc4kLbwfNvLidNb/07r4A6i45KOKOQK2tqOvWDnC/B7
n0i1L56pswVJjY0ZP2XSC5hpWjdCVQUNlIsNtJCviRWlg/YwMEx9Tt4ojd0e+QwF
Fr0kpPEjraBCNTkPMCZuYEqRataHLIWzJnnMIVXJJYd6S767g8BSOrKJL+TKutZ1
/Sped2Ov8xokLU6rlElpbX+9KNHha6V2IW8o6qIqYL6qiDjbqRyAahn44Os4xs8o
guwFKdHvJZiRtMbzdjw5JB+VdbrGa4p6p6Iu4d0YJnS1R6vbPMyrYeV8tNSYu04k
iKEL+LqyntrxbSi89k7iO/i5oLt4n+IIIJ8+UyTK1Nr3eb2nvvGxbAHJ2t0Cv4wN
PzNF52shjWg0zayuMojzSszRqO36XGLfN+YibJ+zTKJdyR3LM6hDktgkgbjC1IUR
SXmDAtmWMGbLWKBZtz+idXf7G0DsUxFU5ssoCNn+/HfBsIIK71Sd7fZ3N6TXwXct
R4hYT1VP1uWrcZYcF3g1J0+wf6p7zf/p5v7xP24eo4YpziguDzPNRvaDKsy++KzN
iLFqvjIfrtCpegEBtQ01H78+zWGoVFU+gngFUN1pPKr7yVBVgCG4DdE6VKbSeLLv
44T1+ajjfVlJ9LqkBauyWGxjYTapMVHg3BMK197yVpfDigf0qlJfFsQX7cpeapkR
Jt0BfAPa4rxXh/KveEhZvxbVombBkhoFdEJl0/7w0MrY+jch84WBG9yOMYMFsoXZ
U0Lt2EnF1Y8/u8TkiKRPwGYNJGRAWtctKcxlOiaJRy92WMNc028fNmxnuoKRZfOO
qYeopmVJt36plWvPHR6IkCqvOus161HgouVEWtC8ECiThzsskYLAjBzVAhcRF5VJ
cAVdlLXSrXCih8lstPbcjKuhzOk3BaYrGQdOUZV/KoYVLzaUXcYRUAFhsLjOgtT4
jAF9kP3FxsvrGhxMJBC9cCIGO6fcmM3PWw2CRv+PB4wbUkZK4B8SN9+UTYZdr2/O
5sJ0wNmSRSbb1nZT47QS2HFo8GqhqMmbSILA8dyiBw6xR50nMTGxiLiDvpUWYmtk
LL3j5yzPtBaDeLoj/uis0Q90fCT79VtEMZVEuemmEdb+lIDnrKuTikOjbnXYE+73
P7FRpuqooQbq6J9tS34Dm1SE9MRsveQZD66DWNwGupIzb7AWZ2hUiTfRdnRuwQdM
qagdKFLcIpWBlmHmYnQyE29AGSf4Rc5HWGyBa9XB/NiuLPFY5H+nKlmAMJkbLWul
QzU81c/Rf9GevhJPApghV1utIvlGjFc6w/g9XRkNV88XnnxTC/xCkPlzCD8CzrD/
WBaNPNt0mPofLPZmZLtKRXixXJDeD6QR1lpgsnla6dgnsCv/jTa0wv0uhQLL5Z0b
niXywYuqPoYPlObgDvhYPoMb9/EbPvWWfU/0WbSut3Q+t7ePWFCiQ9rJ4Px7ToDc
Wa9otlXednA7BVtjuLN9dcsDcGFo8FcJMsj06YLnW9vOiu74r62dFhM6JyyojmyR
/dMJlZhbKJgFtT2/H15cHd/vjA7ZtP+XLLdMwxO83sl/qaOSLZjznUJ+DV3/De1C
MIbLPqX7FzoyUnWbWqWRXmK9GCRrpDHD2dfep+3Y0FGqmrMW1WvMB60NX8vxOZkw
WNMWKmXIlLv4WSTFE3a12U8qbgEyZ9gXZ00zyRamRAEQBkjCaQytu7Bt8Bm6tizS
tKc/JNa+aNB9wy7+Yue2Z/CHhUB8djkSOrRcTVvW6zz/N9wqGjQcZBL7m0go0iKj
wNLIdUEwHrrkbZxgTepCtzzu697QO+U83r5GYbZMTz+8KQgFCE9nx+WChMP7Xldg
RQuJPBjI6zubYBRIWTDlA5EbFik6QTxBOy2mC0y6C9Bv6VzS359ea7Uwlz0E/dJL
4XGNGQdqaELINfr2o3gC0JWq4lI80cMuzQJrnyZzQYZ03A9+cFWRNofXhcvCO6TN
OYJYJ9a0RRUtAttYDLwVALlAo1+TlUlGh4rD2OYMvjnCovNu3nFmODDi9OVw5uS1
RkjDxp7mY/arDvAmdW0QnZ9qBrUJSgXv6oOs0Hhm8XEIX9V27fiKEaMZpfjPTrun
syLaqTwhmZ1JGFMmGo7AVwZEbZxaUi2iSVJhb9uuEaJq2GiJtVe5hLtnYvf34n4U
AV02CEjeNe8xv+IwVEvc0DccgLbM+qM2Xa+qatthzKnNRPxICn3A/mUXTaBdtAwk
waxekVmM7PdzETlv1LXTE2xYcwftN/4hwa/gj7ivvEKYMz7v6BLlfgFKlo/4I/Sw
FvXKpU6t4XUo+MWJOFCdygjYLXBeF933j5v8ysZPnnz9O4hN2+dtr14TLGUqz9kd
xsoAHQ4s5Fci71r+r/oMJ9JlApnBAKq5fWVQg5HeD8PIq7k0v3pSS573IjMi56v4
I37y1Fl7GLVQppWL9O3oGSDQPbH3YvxPvFess33WkmlClzUfYd5anQziDFQlB7/1
WQ2fTTKrMYFcuzK2ZSQPeoZzd1A4qjE6/F40ew/98nUVVIiPQI/9iiIwZRAWVkj3
nT2xE/R0jXoJgHehtiWZ4vdZsUGfY2C8vX0IWF02fbXXEORoyyaZr5yhqYzMEYXn
wUQTSqBFHbBPv+lvdPtmePtjbscBjeZEtbi2m7h6d0Wsawtivq9PrjVanLTYQDGB
C4Q3jf1HJ65Ep9+ED6fhPk5yHZIxcWEcsdcZxDRutswSfeS06tAkh+tKlXQ4qFyW
EeDFXLZB48PAUHmyUwmisTF3HzHQeANw81aaSYZEPmXHwdPFtYszscFBYWJnsH8l
AJQc36mfioucUfKHts2BR/IN15N0RvZ/WpzUHqd0vdoo9WVO04wka+TV/CFFZVyf
9kXSHhocNc0bNyJxC2gfgEjAxYHD2lMOTNlyqeOwnT1piibxRG5BEJYy0hXa5TVL
OZTwxR0IhFyjcQwSAyzk3h6jfah6Drw7JHIalwHPx7osNlJ1U/4UVUy0kKo/a+S2
0x7ppuWDxp7rQIsXyERzoViH/JTKiXdJVGwKAx8ZtpB/KsFj6hyrb2RAUYTxPV/B
up42hXacEhRNjV4LG2beT/pYjRmNAwz6xL31pbpfNv9+151oSXCGI6JW+cKCmIiM
Hr2wKsh3Qw6ZWLC07J+3jS+xJCx3C80o1lpySa92D1LD4+HftDAKkR+WbjnGb1+f
v6xnJZlVmVw0X7LVFG+eqdyZG4GcyUq2e4bmNFCl1dxSH2Xe149O1W/hF4NMq4Mp
ZtnffJlrbfitkpVKSOqqs8fIcKpB8DuJEm9G2s36MkLrUg/6P/DG/fZaPrC1pstM
vE2mqvkXXUYJq4NGyP3L/DIwFY+Z/McQYY1Lm+q9iwT46C/0ga/ixcCHsQLx7FZ4
3dG5bnIhGOVcqvVdQtvJIWCP2ljOsl5tSshgMGRqMcCH9vG5yWTRy5vHX5NQV5Vj
MoHm9xzi24aq/LykEIDvPtS4k3Q69CFJk6vX2XxmkVY9WcdGppP1k881k8sWbhdQ
XQDtrZ/uLf3GlNCW2D6VLRrQljXEngsqNFv9JNdYl3Xn1I5q/qUvZh3JgzDGgYaq
1/kzv7naG75ZP33yt8m2gIw0n4iyyV/TKOUxCc9v/zw/WAgCbhEoF886NFKnPv03
WK7w0pSOnQGR/dSNL0NzCTFq6Z5A1pC7Ltww4uWaF8g7nokO559ol7vhMytLv53I
krXvdxHtTxZcAadN2tpGONosRHFOjQUWPpESBiPP9dH2+J1evgHDPGA2tBHQWH+Z
5uH6FIGJyOm8qhKBMPWbhDIshDYiPfcgzg+b/ctcyfp6iOaw+9rJoeNOJ92fOKyD
df9mc8NACzgNEQkMENy0JEeOdX3/+/k+nv4v/2BNLh81f2f1l1FcSbeu5Jzaw0bj
2vz8BvnH79wIzxcOIdmVmzJmbhfWlUTGOXds+uT+7/O0Na3d9t4+V4qQdPs+DaJ3
r7Hk23EknRvQo4vhc0sZOYVn1oF1htvT9LTEqOSqK9HCeMp1OjqhQhgBvghn1oBz
w8+1eP2T9HrGCW8bzLFUKSkCL0QTz5oydJemrs0DBYlZFyTAH3sVVyyvXNPlUhk2
6nqJPliovFa4trFMDD3bypDQDzrAwfGChPCTf4chTXJJ0x8ZYW5a3wQecydBh7Vz
Mjl4+wICoaFo4yXNSVWOj03qD9xztpz3ShpezP6rUIaMk2rAezIEW+YOGPZGCJud
b69c1kuopENT/8u6aSjV9gZ7gHqKXFDyvqfWSfyi1Od+Z2i8jAi5E6XVXKpmAPXE
7r9S/+VkNAfsY+JtO6FrkAYpdxdmCdlHFPv6244SMuwzsnwEIcdrDlsOApWYzxJ9
qM8EIpS7U+g0dKjVJ/71z2tV/FOSThluqQMl2DuwJ+TQqzNf8DrJdQztZSZWZ0UO
gnhTTOWW8SW7RtGa4KdAxz4OuIMc2i6eVPRD+pA5Gimam2rOiJ5fJCC+gpoXOm9/
oc1QQxSke8qO6HG36p2sBxb2WfvKkguBLIcLNxa5nniJSNCUjW51Sz/90TiAADi4
S8Wu8lmwWzuqqpcCVJ4d8qb40M6VsZjMvcH1ETaoPAeH1WNXWkHVaalcmq9uXc/I
nhy3zbyr7+E+3f8yk5mym9naB1pPEn/UWlJLqQABt4y6VbB2bxCggibnjH/RwivE
hpoA+sE8xavczl+BojerLGklj+eIxq6AtEo+jq8QBGH545P6YhYQsnO+SWsFAW0J
+17P9MAVPvhQf0xbsKmtyw2gImvipnA8IDhgmJvrMtjtyhi2gOkqvD0ehEmjYoB5
gJdnJjIMIfT7jCIzLD8HlQCFA9pzFGYrpFlbBsjrHvt6+/hwvYxNchtv4Hespdf2
g4CsSpe6hG99mb3yAyDxVCYAir8PXq7rAWBeIHCeu1KcGbUn6kQrpZIbfybVeZkC
mJYK3RXbRDcgeK3QJIXa64839B0U0QQaxRkyKfdhnhBxwI62upVntJ4g3ITXXHmG
zd33r+F4RvHslGRpzeuSPFBMp/vZc33mt1OQOkBqRpWob+j71nmL2MUW45M5QnUY
pu8eF9/PuZU2QrtQpB03mpNlO7Ke6RrQRW/tWRWUNUA28w37yLkVspcX4uqFUVuv
QC+w2/WmVkaQcTKSK7PyKvjsAQObCjacnBLbpTd2/8vrDqqF3Qh2erBu9tUoSvgV
Pb348MO1mMrtDXTdoikTnu7z8kmGra3psnnIRFbPt1i4Q/w/OAgXfirFaDHBkLkf
zwrYv861TTqQRbMA+7HWc/npoP5m37yR6SlS8TH0h7oLy05zy/P9WnSDfrEj8/nt
CJpScVRbRg2YUaUlO/6eGbnRd8HHvgEDf+pFN4uiZBRLeaqeMncMTEB0TfE13zEB
dOvD7BKnmlNm/Erz5kVwx8V1KG132rWovINE6WfbJPpw2vHizPgQN0uXFGKHltTq
QJY3bc0yFTd9CfZFC5gTV7FyWD1oNivHeFT1SWSElme/7DCChQn3/9kozUSpQZ/Q
oxcjSNi2HBrC4FcIzuCb5oYgDC+I6hGZHW3NdDFXAIzj7bibrH2/Dqy6iDrozWyi
LThfWAE1AxOGxTOOkkjJU+QSjy9owifffPGmkaqBlResWgNSGfZ/15DVJpGpsk4L
SmI34TDgcnu0D5wrB46kYawKfIYYqN/PAA3isjP8n02fiWKxRRoCc0lGpAfcXZUo
IPwNaqw7uPbM4cFWSu3V3goWAR4EZUeOPhe0V7p15Mi63s7URKUbc5nLyYNuE8L6
qwLWhp+Q5dIzLjN5dCeS6BF8oTIqVsdrYZfVTEw6OGALrxgOpXemtvPSmahlyzmd
opL4LeSaUh6WowtOyW2X/K5Bx9N9eqSb0iUqT1KSyTHDxG2ESK7xo/ix4jR17r9G
wbLmU9WEjs/Ksg04QtvquATR+w/5GcdjAedNdmf66CBmwcQddqa4DlyWzd3m8o9/
JwO4fnElom+A4TnIoAsnHMdBohiXdeqCP+gmsYDKa9yNsO+RCBarzvvhpHKygC1R
U+rGiXNui7W/TaV/01WO2uliZlWPcbMpLfavnYFFfzIT0U2rp/evlPqoJcMqkRGz
Pp9Uc1Vq5Om3a8ZwPljYTOAvgWtaB5e2CAlTgm7EbbFvFfRfUzPzAoYVtgHlSEYA
PrK/vdU/ypzDx/pS7YMYPQN9lwe6LKzOdk4hVH3z+GHjk1ToMIaYndFAVzsjN24h
61oUQHgo9HE/ZUME7nNlwjjbIAt2cCqN89ijE2+lk9WXewZhrVPwywrbyLrHNLG8
QEkoFZtgODMGMZ+gV6fZ9tLu4ieoXInmwBkFrowLvu0BjMueGbUumtiw04r/nVbr
4DFQd7O0kB5YlYNTi0/nR4fUKe6DkuQr7+xTs6P94Rls8lHFpQKhXIlCwRUrr3AV
lhJ5JgfX6EmwdPfYz9zcMxeA2Ix6BwCwWOwzcgsHz/lmhJsrAfjwWrLEtgsR9Ln0
GCqMucSKpwlAjoDVY1vaVbdB83EoQbmQrPT66YBQTUc9u3UXtO/5xSy5P/+LJwHl
KE8vbJZyRSAFSUakQ/r4uSWQUTd5h6d+32XUVCT2AZvidF/m8Km/L0P8Dz0UKJl7
wL6s4FHCLOQva0vu+VOPNOjc6SVaQNXOdrOQ2KlZIlaU2TS2SUP93IEMK41z2ItF
jW4ON3or2HU1+fN4wbEo4/38iBuUCjKvmr6OI6i4UQnPDSz/2UcVxNPgbaoH2GVL
D/gG1wpCrcavNK1s9rgMoQ2Y1GsYB4GQO+131aPz1l9MYl6JL4yy2L+T2PjOY3se
hM4H7L/e7i1ugPJZnD14Ze0k7KpCiUpv7P3oinn/hyvWVqpFYqM84agG0RJRdNS2
4pSQe1CYPKxFdUUTfVl3YvLiDJLPczxIgYJrVqEVRBNmxINP9tratw2GWBpcD/dC
bt1i3V15kBjbkFqJtHwNq2B7TK27ZH/dBt/wXW5t/bSlnmDdorc4AU9RRfsqYckG
GQFXXtMA0XTGwY4qVHMBkIVTTgjhWmTuMYB7U2RKapR9JrUNBgWY4doEXEznelwb
arw8/j/ZPz6iFjc7iCU0/k+sZbMF3+0rzz0/vjM9Ygzh00b/uqyiVbOES7B2mLvW
R/sgkK5B8z+hLCSMGVccXQU9i+cBCcanPKSeSDC3YuhIcjcSXU2S0DPvUVQxu/R1
8ZKCRa8TqP6UNnfhY3q55w42m1c4XrDPmEA84UCoHNzBKKJXUlEoiy41od1rEwjn
33cNA2NzjmsZCmXdWHrTPj5XHZPD3vMamtXAyMxaq+spzoJhz9ni0rnz9o5VgkBr
3N7jnyM1wIc0Tre1o/X87X7hbWa9w49LRQHS02lAhfclev9C1F24Q28ux4MDu1Jy
Fu87fsKYy0Hp0m1/jhgcPlw/Zmtumtea9tby3lVprt2elZ/u0Eh9P97VznmSBkxg
KyQY30Db9CvsFhm/9xK2yKvMPZOk3zNPa+zmQA9DFK8ZIpmPMcrTXkDmi6i1QHgi
jZ9ra/A9CIdJ9bpcW9yJIV6ixbjrUdXmgjSVEaT6SGjHWicLbtkLO2tCUB3Vi90C
c9vfFyomI3g+jK0lfb/b3+QlfVbzK6t55tRoPIGfKAFfVR+mhGrtn0117a0yYM0V
5+kdUUj570XQmCHdBClmdB9VtndNvN7YGuREHpK3htDh1cTCw1+j6exNSQ+HI5yG
Asw+CdU9rAgF+iV80Fp3A3MXGcS0ThM5LvvEWro+FrtvCt8d9FOgyFqKAh/G6tNz
lxq16UL/Oar7dQTfsV4B3AZJNpszuk05szNnKysUZYSWZ8vWCU3s8F4S3zJTZt+t
z62d8Gn9KYPNnoQPsZZV7Ep1PkPAshrbjCFmc7ue898Xepf8ePqMriV1fm8KDYAt
j0eDPYb6sa95GBv8caqz6Jqq5n8Itd169X0LOkmUr27fP6IcHGRGjmbtj05vuR0I
Ayto0jxUovH1ejOWfWIIHHRQiJi6zC06HYuQkUSGCmO2x74kY3Hs6JMkSq/+g0cA
DOzbx2pyV5Ks1rL8kfCPvDM3xFPW18CLmgTrQwswcQVImc7cnxsIZQMgdAideWAZ
ktkaT+7VKFHxRMTiSc910xyOge16Yti4jM8nnAW7GEQ2sUthy87dV95AAXyP24LF
TtJLXG8IpdBG7sRCN1ljrljljf3Jo4uWBxxU2NRHn07gETN96TCrgWPN61akBdbN
xi1ecTaGsYJMVg5cPh9NljVJge+977R5/J/3PCOyX/HxA855DdYrcT+4QbvZtzBr
4rDoExMo3t7BDJJkJ2xNXuIl1lvVkAvNhwjaTNhuCdjoqRiNfAQ/ewvS9fXbGQKo
OKQnMg1LKQxOXDkZTcAV+Na4SyqVU1C9xg93qThlwpNN4m02jpRXb3NFPOJOOXYk
HekRixoXkcP2IsbH2NBG9veWwhAMBIdhButtKgg6BI/LBkXH0FigzuuBvPbEf7ch
QJa0lPDBS3y7XudZteyKrdm2TE+b3H25fnpClj+XeH2nnkIN8ZSBmbCfVnpWWtM6
0wqQd4UJWpTKSUVbmSeGf1OjFUGZgCRxwQwzDCJFxs8mgnwxmv/G/awwBGt55c8n
QVpITA9QJCOWZ/aeiEcxwxQBpby3yH8KL0w3H9WeVAKk8+M++O67ZYyA+uhii1ds
3dQ3P/v1MZSwoIYCBc3pr38bqCUyR2R6Y8ht26W0VqG6eKp1fRS2sJkP5bZPZc2v
UwAhzPKGi3o5Lzc1hQl6kNFamYFzpDmFY89F8PAQqF2MZqBLAh0nruAYTkt0PDoQ
hYHINmO/GZZRk4WsNNaSE2HDRB74uhAd54DCTu046VqQ7od7yMOtFYaEdlHThGGn
jkYLN9DQiQ1LlVpVzeFk0zF50KEYFiFA3ROta+JTaRpXR38kz4ewaF2Vx6Ao8ZpO
FrLGPEpNMaE+Z0BkEiN2GkkW7GCh4R8b8lWiGG9YCEvlaPhvF4942T9136+w4U4H
uRulFmdYPdi6FuXjDQ53RoMEG/L5k8ZZiw8RZmIkVhklawBe5+ODyvs+sGAtzMlM
bADYuRQcn2MsBeT9RwEIxTX6m/AbNm8+aLmqu9ensZD9dk03tTyiTsqc16Ctog2U
mlyD5ZT1qrTaH6LEsdzHIU5hEBZF1Wp9GGmWyiifpyyKitEfNe3DBi2NdU/5O1Ah
VdHdB1u+fNXuSuzVGBBXluNpbfuQYfmNlk2DnCqzN7D6pUQHqVJhF8OkQ2hyU/LG
5mdspX3a9SyILi0E3sEgnp6pB0QZIYcHK2Mbacd7qexDl8DgNM/pUtfet/65BYmZ
7zZQNSjmDS6LMb//6EutmECpUYOgqbm9Gn5fsx7MKHAOyhhSPVjudYG8r0jQg5jT
E3aOSDoGILamkGfoUmrXz68WUXWJ707+7ZTa/A4e0hMGQb9rOsIZ4jvlrWzgzok/
CXeUsKQINZuRNYtsGXxLG+59nmJlAP8LebfnbO+UStSwK6/+nob/+at7BDJ7VVIS
D7+3Hjln+Ivx4YouETwjmFjl/oDHTqq5+hvCgn+mE/Aq5i80T85nyyHPOFHZZhTy
7imFzKbRIYBrDKLWgZGzsrfChqTCSgb8M9QL2mW3+6h7jDqQyxxuhC/+f0Qe/jaI
GTFEGSjzVxcALnc/yFFitwtFGS+nL2AELuSWGm2VtacqvDkfG86rxYfsn5OyC695
PXgJaEHo9k645XVaKBf1XLHErthXGK3nR+xQBibc5u01MteKUCMoIEsouargG9GS
zNt5DDfbiiS8X6gIICtjAT4RUyhwOow36Y6h4FtdPQclqVJISl6Z3aSk6SZqMpEM
qrk9ze/vMZ/t7zX4eVSZ3+jf5SnJhzPm4SOy5yfad6HBi3lEl/DE29YDX4gEZnrX
8wle53msquf47iPWjcZhm57KsAHVUCMyr6l4wEXJQKDoTRDJmPxO+OeMZ9Bm1PMI
iOZs+sXWRlz1D4Xi6EeoOUEGJbxDqYk2F4uAlRAflUUu1/LfyaFTeF2Px1Le0ex3
1UWM/Pl7D0eH79YgB5j6sP9UolhQwsBQltyjHajCjcs1QLG7AS+zx0s8SkWXEDc8
dOaSHURX1eploZ1bZp7qBYsBudow8v5mezUqh7Y62Mw2OJXdrr8mLnMZqHNY6dfy
AcPu5YH3w0ZKaNFh++LudyOrOkpruWSiN7d9gVk3oVexER8wKJfHlvW43fB4qNPF
Gd4UIWtracjzT/fsBCsFW1C2cZT/Lie5SHjcTc1uq1COeY7wWgqwxWp1ZiRlxMCn
DaFuxk2ZIeYcnEPocehYCagW39YqJSw7Qr/B2Sl8lrazCC0AAq105hTJtut3Mpum
bdq2bSSKjwFza0sk6g4BHC06QCwy9v+CCCwtCdQZdltpfq/WwjvI0x5hulA7pBvV
PAJfGDE9eof3lUaww3k+8HtjCCrJJoa60X7S1Wx1h3TKD5KhJrMTpxAOR9n6vMMh
lQG9fUdWEstL3JAaZEns1j3MdeetzN9OcFkFdyKiK8+O365/xgv5HXlG6DHXGiDk
f7bNtzanK/t8YevUICxjxslcsjgDPmjsWkgejBTlkMt3velGWYgK0Vp2z7iHx/qx
BQg32iDAmqSs8v/8v4RrFUPheWKc4z1fwa/WJpfP35J+WOKqvxUp0MBPuz+qb9io
TFGHLlc297YusKjPAvtb0N88Z2Rd0R0NxWiQTjlzDth8CiRzJT42nl9hRCI9LHHL
KhQsLKy3NFI3uC01OWqs9zFDSd8cEp0NLLiGqVqheGIm7oce8p//CUDSdBa7Uxuw
F8x9glkZBDHv8ul2wC9ShimaMjYqp2tc42tw35bfxcIV0/1LozOilvQ89i0kUkNV
lMlUTJCTSssqbgOtY2zqUUHQO7I3knauINUcWjz199xxgnd3oBQHt+D4EaaQC/L+
8WIwVHPM3PH7OpiQCUGinLUygoDgZwweqoqTAgTe5yUC21U9/6Yx7JmUR7mToKiX
Wt05Wo/3te3tnV/qzD/WOlA0otkcAQNSXay5nX/ni2kOyp0zl59w0YmdhDMZeCj4
TyAU96VJ/UrE+DzSgsdaPaLcy1OopqPs9Jc0QxFjyx41FcnzXDoW76i3WMcBsmk1
WusKe7mv1nqTWqkaCjUbOT6ysPVzyKalSinUWvMYW/9sx0Qkz3UW/DoWboEV+OVI
/BJokFcPHWBcoXkukIy4whqto2h5Zhfjf61aG5EwbVy4Vkw4zlj2mXN9OcBpINmi
bByxkTr5sRuqItyqeCeb9HF7bngq9lBXohhzKJzj5IPDGull2qb6T4vdpvCEuNIv
YiZM9abupZJu1qPshaLSAd5u6d18S2XhXGQfU322R9i1/f5i2UtG+Kdj6+uANy5B
7Setn4EtyJ5vhoeH+va/8VsgPFIYLsLN7U6o0qEF/RTyVq1EbMvWpWa7hq9nhWXR
H+n17W3xPtlUCeyBpWt0Ek4wJ5DwVtkmXzBzK/NAC4C/NgmF5u7Qslb1+lobqgWO
qYygjBqyU5NIom0Z1lPJcBT1/5vgUdDkl7n+Rm7hz/c1TlRi4xM1WyV42UM6LYqZ
YTvXXrH3in+qAo6nL8+520SaGATejqw1EarFKBuAd0GW3aUWEswfB7NwruDPP5Zc
3p8nE292JZ/lGMo4BTh1j6mBfsgibXgher88LlpfzIcL/WSfGth+BBA8YCoMlc9v
6f2cdYmPqqZ/R7w0ioECup0mcQgR/SWyI/8hoDghlCryPwf6+QpZpVox4Y4ezg51
pN+WqgPQPIekt6495E9mQz5aTgUOyVJ7FaYhxOmW7E0unDzN7eebQiq0OJRLK89H
w8bGmVs9dDJ8EsXNlikcxfhGQJMUbrQbnpIJaduee2EPnGoEPq/0xCeBDNgmtY2I
HJEL0zbXDOsLnCE3dkZnZwVdggGmaD4fTeGEAJsY3Db9qHfRnDqvpFFn4R+sG3h7
/toOwRIV3vRfyA72cBxShlHpg9L1nVJBHBwa4ZN1UgVyrXdMisosnIHbHTXUeKq5
g2AIVwTnWwrvwhzOrYr5jCMMT6YEBzjNrQktWUl08kgDYatz3DuP6eet/uHbEz37
LAeYojq5JOHfXJLMd3FhukOUjxxgsrHaz+0IWbXkgcSnBlmYY2B1boLYk70RF7+f
BnSu9lyYnfyswkaczpsEgtzLGhvlMHiBdPI1jtqum8wEafOIT4wrh0Qt1kBaCrKf
EhLAmoXqe0rs5raPe8aQ2tG65ekecipoEHjfDhrpKEnGMmdEdHfogbJCFqsyRSmS
BF4NhIA/vb2iY8QVBM31RUWoG4FkIBF2fnbYoMBbQ/BYOv/lajSE9ot7jEn2sA+Z
YL2hL0teE6zxJU+lRQ65mwpTpNGNhbGaUSrT7sdf8TSPS3ob+rdmkWOQ/oh9sp4P
jDzZOWKXtb/ExfDAIGNtZevW3WPBRmanFxXWRD76qFpFqwo+XejQjB6zJjNmqH53
8hD+4/e0o6LlR5oMjdKRDqFFfBOoWrTALkBaK9Vw/lcenHlw/bqI+90/OPf4ouWz
/NDOimMMIpE9FfpWET7gey51lePmW/ywLdvVS0ixtSp9op978oYQO9ETLJbuA3/l
HoMiB6NnqAlA5QUjuvuQbcN5BV8iquePRzp3Vn/chguDPhF7sdQ2psRl3/i9hhEB
/aamOVigxZYJWycBS+Np9KbnfIMdtJyKNQhVk2J5sdL88GNxgqqe1h6so9HOy6x7
+UFBQpN2rxhEY4nntnKTp9QxBLqnSj1chjow/GwMCeyadr+naTuxeUtGMg0F0ri9
agAhEpSBM8ZC2cY1SrjRpHivPHsOxDYvG/XvFc/H4BRdMHrw/CXBPVXGeewk08oV
QeocqDRCJyUS0kMuaiMbwH/7NraKJYXPMBpi+P6HeyW57H4EIft3rIFcFK7aapKW
wPZHDZToXRcThZrJdYTSZvQ/+mGvy+DTJ3O9nvgmLLmfP2Eq8V+RZ5vLTCIXKybP
3/ZKkeDD0ByI5U7aKfSOwn8JCc8p3Tp3vA7Vy/7EoS1aCzYNG9T8auRfuzn48u6O
KeoL/0XJ9z+H9yyH/HC25aFteVdzilDzpTsiAYf354uHaqLzAtwch6xW0Z60FgN1
+jJ/9QKjpN7mGfvqDQ5SJsDpGBdKiQnEpyJcEMf7QvmWkXftMo8zIKuB6PShaUNN
HNOV6na6qjMpaJnd/dYoljF5bbAQQwPiPZs7KcAunMw+KoTxcqXE8Q082nM814ha
ApoXyKDUYMLDvtryVwfjwndap3edifHor5J5bAxCbuNha47p/l6tAzIZX7B/Aotv
jNauPoZCsq7Wf3w1RPfao5vWB9sekWV9P9CxPGwYRejthL3pWkXcGQ67k0Zl2VMY
axnI0J5V0RfSPuwGClon4lXb+wNjD+T/XmEWHUqLCh0d8wXE8pbOXWmNTXULEg51
Kxn8/OmS82dAaKcN0fKy82BY68iUaM48zRyKuU7/e59+JL5DUdsSkjnibyhkaoiI
Q/Dj0r6VoWUF5Ff9Ih2R0p9Oh+8vmX/Bk1yXu4RcUqExXEyYp0iAr0TzL6ghmO8d
O3Py3mDE5aBMj+92k6UafA8eaFeYRftJ+SiUYay3/y3gMB8CeieI+DdWqm5XPm/R
TAVPSgw7Xqa8Wkvyyz0PIj/xp3PDvKUEdI2UjcT/nLotMzT4N7eeOp+IpQiugJuw
aITmCH8kaZBfqTyKqFEnftnrn22uhHZtQxSJgL9dcZg1SJnSoE8+IcVIOStUoqXI
Lc7DLGigjppckcfDb3HGBQa13R3yI6u9++GMVnBZQrJ7eq5PnluzAdngCtoGsXdx
/IqhiSSRSwxa/aKWF/bYRg8BXnH8Tj5ZSCWTqzUBxZSWt2EZZ1xOTcfV2oa+Kxbc
bo5w/KbSOTYX7NKNxt03EbkKfgdTkK6SMbv6idjvSWapWLhWvea1wcscR6dLILO7
M+yNSm+YYZOmVp5otkEvmEUvQJ8YY+QSxPCL5PZT5yvh5ZPasMcC0gQMG2ISIe+F
q0FQucQQP0euSyc54GpgqUoFtLSqDZxxXatEIw2m+D6ZTXJyJlRy78TxlkHhnHX9
fj8ErrLXq28kRFJ6YTQTPCZjjIt//mICIzpiC8gXEGe4mk9ri98LeSN8ou63LLv2
i5L5b6gaLz/KAenX0lPzetdkAXAjkYx+iGZFEU/M0EnOiF7irezUd/Y2dqfgvoB2
Fyl+Tun5/EdEAz7g4HNOv2FxtrLoIjX8QKHADAIPzhIxh8cpgPWpi61Y8g8933gt
e5yV6FZHNTTg3rI0rcw7WPdGUWp8VUeRpYCzjcCCcy30RoHX0Vb7M3FsJUkBtW6q
uCorxxwJ7KqjuTjqjrMuDW70Gw13GrFGSs6RzW57hbiLEI1dd90DqREROorkdqQ9
7ShT4EB+22XYajcIbxSQq2aZl/JNteJNpZaG1SPQi2mfvCQLwvD0mUjBi3B4RRn6
JQr/ARTqLL+jxmQQ+8mdJvkCcyl1mnAUCikOJ5PkF+ZrU85ox7yUuWZnedXVyAi1
lHs9/3t8N8KmWTzdYA+CY94fc6HHjdKPgC2Im9wZg1WPVQ5ukP18FjitO5KfV6q4
2r3x1xpmBCz50pvXdYG0Esut1K1t42SJV6skn8pkDVp2JrfxwjxvdD7H5S9FctGo
tPdl1oEEa9NoXgfii17z1nXB/x3PaqpQGcDE0fL3sOOKJCc8aWDgRbZvPGAPqRea
5TXhu985QFilqSQ6TUtMsYwu/chC8rvRqpWc1cBkOs7eGrhFtv6yiUSfz5DSulPB
EUmupU6SBbEMjAqMo8NdpfwKfS1WhpPsKCOSANuX1tCsHUywN0Pl5dNVHsSScLCh
r2ec6llt2Fg0ZPmJfScm7ezFvWpSwOEnpbwn+GwwxnohM/CHQceLVJjiMFTy5aw/
nUh0hWhmWhIf98dLsh4ohpS8d40jKWaJc7xuin6NT4x0XbNNle5kSoa6vIOWwJuq
IEKNGnH+V4YlXA3OfIuMVZCzD6WMkaQ6cNaPoVYtumRQNcqsmIFaYcaQc/3K2wE5
myUPVIg3cmRM60dh3sAx6taxKNgn/3D03Up3DyWfkwXaqDG4JnI7FKr+RyoJkn2b
GYZZWLiNhelBj5MO9ure0s/X/b98or0fHPNNxSXFEz2O1TUfhJ7lB71WDn9OMELa
G+8AnBmg2U1HKDfSmrh2+d3kWRCYHVkxL3SrHseVsfmEqmBrXw2jjjZug/RmTYQQ
9xPmw0US8Iei9UoR/eRwoKJpwW/SR99GS9Z/4JcEy4fmjfmWw1EuPipcgXV3yJJh
MVg39kZWWlbni9NoBlXotUBsfrnHkeOmAo6VrMIUxWVkb34p2ims3G3At+a02qUY
6uSU8wybBIHCZao+6TpWAZbHYf/nwzQfEtaiEidQXJmhiS8G+ZCUOLwWgsCTW6BM
PBbBPZik2/22TyVFIFn3YLEqvvo7HqG0R45H5maapvivqxR6IZmQeCyiVpg94w3+
rH/fSc/WXz+AF+Grh0ZPtr66okgYSVXluocHjh2gwwOuAhHMDABatdTUn7d002B8
jjYkhyN2hFlCwlO4j/sRTWUXB3LU2rryKV0LiJ1y4nUqWGIERpl65+MmQoxJ+Hfj
5MJJGhrjMfKOZ8qrQnpZWxK/QnvJWm8KM/gv2qxNuL3uB8M9T7nP9ePJD5q7XsC8
e8Jznvpjr4xi5fj27oAN2UR7gB5rU+RORABtwI5LAcHL7qXK48574/3THYwIrtcK
xRZPdKsLawm1YGKIlW2mTW2PrvyJ4KK6XU4tIxKH4sV78DjnAhzh3C+G3MiT8dnG
R1Isw9Svu38PKdZNhC/89M4cbtKzCGNVyN0gHbcrj/mOXUucSnpciQz9mgwv5Zrn
4ss6auDKv74fqS+d2k+sXQ7pe6TpmXjjodrKlKGLF0c3vavgX0Yi7v8vPoYA6t4C
sEon/HUqsLLF1J6jgntO0UkOvaB715c01JlO3CVh2AVAv3LqO7RCYSN5GeAVxxvE
PRTElw7Wr7TU0f0QSQMtGXKFGmwj74X1CW4Un3YwM03RBfXr6kJj1AsP2WSwnoG6
spka75NlbzRltANo8K19YCtyZdCogvL1mPUy25rFC5x9GLj8N9DZHYkLUXEWEjgE
ek5EQzrETy0sgwsgvo57cDF/WG+YxOR1SAklPHbEOclMDpUuPOr5u/YtoCIsoJJB
8/fD/r44ynZooKyUyJlV/mKmFu+yUIG1xZU5+L8EMrx5cJBospTyr16RoirbWlJB
J+bNzLewi27CYQVBTAStbUjzq53uBZPIvQOF5x1MRf85+y0vG2YNrQ9eHrJQ47Ah
Wtkmt1XNmj4BfSjNPIDvjUr5lQMZKz5ONWVY3Wfvk9IV8kCl+MmqRz2gJvMGVFlC
3T5D9GnSJqJ+QGbLhbVRogkT07lYEyZTjvXPb95zyoQ1bd/Oowf7gzJkezEdvS3P
vSrqlNyDEdETF2arW4bcpfmRlhaI1WWiRPStHDQgDCVu8yNUYaJW9eTf6kiTCnsu
3ixUqS/GVf9X8yYIehL7KYktrLYq411r/K02eREZ9hLSShg5FLvULCMZWWydXEzA
bW1llcF2IciAaEN8L7dxGb9hG5TTQE6UW1RhKChV8yltd6gqOcn7ddVqgwaZkYUV
bneEZEcw3s+c2N5INMzFIuEixAxMl8VOL35PnIosJE2xfA24iDcebB6FvfXtz0Nf
uKqIUPV15gplCBYITJIGP292YTHrs+pp9fW8//75E/LEex2V0tlqSFQuQ9kHJR04
oZShbjZfPFr5LvPcUQXeSUtpe+Q6nLiz0Pk7wcPL+O3gt+nzCY4Q4fSMHK+kM/CZ
F/0D0jtbgyVGx8NY6Gg7UJ1zvtAToH5SvtkHtZxr+pj4pwbAyeS5bRL0PF6KO9rw
KYfAHRyAfegtCuOXSxPvjnO3u3x/ZZCgRa4ZgU5wzCXZ2iSCMzDd5woIldCCKpoc
7pUrr5l3NxT7BEcfWNtWNuBNn02TC6ONZ/dCm5UbmTREvyy3dDClknt91nxgzyvJ
M6lNW1C/5lcc0UbDZMdC4Lk/shXUsjRyVpiXqCzkknuKqFAM+7Y9HrvwVu35oxJM
ugk4N0B3tqyRPsrgbyJ/XZlsHvqI3Wqlg0pzfhb8K9+6W1hce3zrzMNauu23/Elh
8uaEIqYkFGmS24Yn/CN45B3a4y8ZwKgemDqUxFoPvL7DyRT3ucfws2xE8XnSd4uf
n1vZddr1/iWMccX5keFcekondy4CzR79obvmzyq4Nrn7TVmbS/0aiyk9MMkaTp76
fNSFlFU5AeHU0IgRd0mzv0wBr9FPTvZvir7LXinJXaJYmY14m6/o7XUSWchPx5Ym
Pt4rykTslLJG4/H8itI7LAvBCnoqNkhU+aFx5xu9aaPmnBPdIa0ERrQw/hD6Pu17
1gN7V1DYWdAoNZE0TEHuJaski+gcAixlytF1YwLxzjP6V0u4kI+qMGJ+ck9Y5CIl
gRP6eDzwboDci2JMZG2yu7m+ueiKYoKMm6VY0L3pFvYHe9HB4IlCgeMZ92C/e9L6
G/7JNN/vtblbSCPx+8bmre+cW0t8apKuBUAc14cokieUGDLUw1bEjqno9Jh9xVuv
7MydmIlJoMbf9y7lwXxFS9WL49jF8U5TahfKNJIulrOcPyXKX2f8kFBYWOfxX4gF
/JI7Zn4bn37MoiZjjMuVWNt6ZD9ZN8re3rOGQLOWFHsB2mHoPY+UPR/fDPCDepld
CUuDkRfYSrk+cxQNYcYFq6E4rZWOU/ID3zy2zma77jeeA8dGMsTy4KRmThRsIzcO
mof/vXVl2Gf1M8hZHTfD2TRbo2J94aqs5/CFNdsxMLathevJ4xaZA3znrv4GSmf/
9eRKLqr6bxEOtXJh7B554x3Xvmeb7WnKgmVruhRMF+80V4stxpebTKdJDx7zGXBo
a8/8TrVpY/Y7bqt8/e1QNUE9kEnigR5KUMFPUYuxtgPpx9Wiy/CsfUv7VVgTN3b6
/eOASlKHtTdBVXylouBPd1BM6QUJ+No+Yyf0snTKJRhnDLfhyifCAcdZVmeiijy8
QOIUFeoZZ9gIwTfCrQO3t+Z/JwK3AC+nfdON4veduirw9Fz9iqT5/IHQQnLyVfEe
RsQnzwLjf8uh5lD1bBfFOx/uET4c1JAsJYh7kb0DiRLmJh8XrZfYMCiEwLvv5RGN
cHi8o2tE3IR7Pnh1hdxfTpjdE+MxgP54Ppz0s/VhLB17xyRbxAt1kxqVXHCvX3D5
epSJb2wEP1L6YL9dVWgIg3fDthoayDMnmN1EF4lJ/iisTbJRbEosRtXdTJEpx7AG
tB50tKC/vyWrv8vV6IfP4S8c6vuWvgr3/2sjRnP/bA+B1fTYECBLRkDe/ngrch72
alV0QNF3ytZnDszVeOJqAnldF1BNiRhaSMVhDwxuTlIoeS9RyoSp+Rh5Wi3XvSa4
nn0Z4nWoiZpbMidHJ9nSrD8SBHpnx3q+BYLrBfDgd1ytYrInWP8PNCfd82/8x62N
8HyCPljFMRQ00PdE3pn5wD0UaLu2olNWUS6DmHCliHNzRFkPeBgNg4DLbydpRNQU
NbbFhQ3PCPSFxeEYLZCyAClw8pb3hCzP6mHcdcnofRqRjdNaj7NNGUWcS2CFVa+/
CPWzrXaeRhPjAeZkZREWmUx+WUuv9hd3qvhgjlIcaAmTaDWSpdhECajWluGCVwtK
9sTRqaYDOF3WAd/KuJPKH4iG1JITVPy9tt24hOpXzSX61+fRwF29PJzv7lCMNhjZ
IXAazeQguE4viUS02fL5+7r9FODi4WZggj6nkE3K+2TcGwttnjQaxhti1YDohHkO
k6+fXGxsohZ6NAyglNqIYH61G2dJ9P1lhPkmnxgEKBOfSm0BkmM+Dgjl2xWMtuhT
BEXd2EAlDmPxtXZOGg7DQU6cXQ5T1C5kdr4zk4usb8X16YOTTHtv9Q3OEvXwijWt
ACL5UbuKV3cjEPbfHKy0hsdVb6Bryg2HdzdiIxZtJfGyaZ5VhWcFlYlD0pwSTfzu
C+JQQWkoRirZI1g8sN1lUSbPrtm69CdP1MT0DUdR8+2Mp2//ew2BWpuCfXXyr8rK
dsIdQ9lOvn4At+NQLYCJJaBCCgJu5dOwR4keDbII8TuB9lQNGChbjbim3yi5ATbG
38NmVmVJFYnEydcEYQgEFCBVKKtbSbcq3EBvfSlFM+I9mAbiPuKLYJx5NFvE72vN
l+R7+WqKPHoBjUUlWOJWuaRyIDtBU4TokaiWzkSyumxmEZlknDbHENW1tPcOWJXD
fNbHrnogUqw9BxyF2rgo9YA1lzSjU1EdBkGT0zoXpt5GYf5rhwtP6IvMnDN0u60Z
mSriSTyNalRMP94/r0hzmMxVbbmLv3X/vgubpKXTdV3JzPp3E2mTFOfaAPU1ukF8
IHB/rGbClT0t5nNRdnZh7+SbuHiY2ULEur/2R0HWhKJuCTzR7RooQei9CgNpM+xq
Lz6llSsa4+OEuwYWF80VBV1Lnosgw516o2z1zb2o0rgTSvf/uWzj60C2Hc+IKQfk
2KQeDDOrHtf8PzIOALcXNT9uy/aB9T7geBJQxwyxrgN8VNn6LOJd6fHcVXP+NYHb
gStwTF3a8IjkzDcSevFRkanW84bj46uZvflQL9npcBjI+EfnxJSXQ4aJUGt2cEPk
0wmHNa+F/BfCdJOeP5AXHcYnE80sCOG6vRDi3e1eM2RyG+fbsVcabIpmHj1kgVpu
AizAVwHea3viLKKnQQEoEmZKvjPofaiCBxA7NqLUjY7BgePf9qgCMqDGNXkzEUzy
kMEf3OgloEnjzez2jTRHagAgwnhtcJtxCEtcrOD37QAvToshtOAzH6FuMySgEl1m
5hysHYi6od1HY8rjHxpo6DV+97qTodC4IYKf+Jsh2mW2m3okWa9Hn3/XoX/UnSiV
S+75NGF5D6l19WdmZzzL5dpWlaQWy3qRDqKYNkoKzPJP8E04kp9vkXeqwvCQnC07
AkLApQD+zDed1mLISNwN5Bpy6qtoY+mHcmHGT22FcMHSiYlYlAbh4/2KDyga00Nc
pIE66SxnuvVj/oRU6oWB5+zQG5W2YG6QdgYtyyySGPBw6lF9urJnRBc2mQTzbMAO
vNBP9FH1S0r40fv6y1rx4bYOp3Sf6L8cjk72Nvb3GGKH2SOcIIbhszBKid8iXBYV
euekcQZeOeCsRp4HWLur9g2R1yZvAe++sRa0bYgmMKa4xVJbYu32w3roP8Xp+5oA
y6RP4H8ifuJAJVXiEI5idEZXBJz1P8PvBxjvIA6Osl0X/IC10S+MCL3WXaQjm4Wg
4kBA2cf6qZKyqN4lZui/6Id6x6Mm3C0QIIWI/y+NSxmshjc85h+LkeV3uyKzJfI/
ZJws7Ux46c1u2P8hg79TN8i6W8tx30nC5nXnMB4rpfPHSYZ6Mh95YOLYvrAziCwP
Qws6bMl6L4oAuCMy76xnJ6jATDTOlpL+HOgw91FXkRUlk6cOnNRy10xCSnxgg9Zq
ZkNt2edWV1AJzu5fFRmIwm+aPE673QSRsateh6dtZRcSv91BiiBE3T6pVBz5X6bT
EU/XOSx03t95m4njYsDlqcOwXWnk8jTus5dsFiMYfTOXNM8D7PvrwfaqLG957Apw
5uID/hPYPR/8kFnYAoxLz4cjgMsDB5LBDeqvcZ+jT+Dvbfv5Pc6B84N2V/sSQkLv
plvK/ssmZ9ZxPhqtTiuJJxYhH6UL1kagtmC4wWe99AEiSoNf1oj6NNfVBdqtP4eV
zuaQ6l7ye2sYPz+UOAgPxzuMY7h1TwGWPQmNG9kHX+uWhtsWeeweFEEFQIrzCQTs
QR/Na/8CtX2Gq3qRQDdHL0H5Xrqkp2Uq2GUwRkD4E8juB/wqzFEH4BgEx2o2r+pa
h7fBDJWUzywRidrjIN+lrOwVpg4FXkR75JQHaVSXkXqtCO43wFGaVmb4DJp++gMZ
UsyhxV7VHgNmGD+ov+welLY7Cdy7I0jz2rwdvzK7Hs3Eg1lPMF62Hkri47xj3KOU
n1RPf1CRle36nflVYvfCPGhdVlTupTbi2lUyAjUh1twdVfWUofcUE3cY2MvQxt1Z
FHQzmUUIb476RFLVMn40WI6tqIJ1cHlbgFmkSP+YzeFibEWFz0R9yGlIt5BE9Ex8
IYq+Oxiu8XeAtHw5w0JxGPufPa0NlcWpOzj/f3cPJMZERxP9oqwAQAWOCzYxr4b1
7OChqB0PifwyJdCmrNTN7BzJ/GiXCrtEOt4seRCIRSt2Fzog+F1LFyuizIdTAMc/
Z+zUW/hHiPRrxhVppv7GmybBFp6EwbIRVA4dwAmVBHgD9Ut8FvdyHEuVskAXT+cY
ijKBlevfJR5SlZWg8BhRyhBvOzmbyrWKl9cCqpKrXJM0p8D/ADI2XMmKcI667gCI
bvG+3Y25PUtV5Jjrm0WvgHWFmsJ5/udZgcjoZXm/SKlMjj3AUXgAerafY5ouFblD
iZiQPGnyEoeFEt2+BqBnPGWD9TT1gNPb3yU5K57dIkO8KhJzJnyehu4VtcDc6GzC
ozTMITKST7wMeslqmLewcAxbOXRza6D3hhV1g/FBCglg5VJF9G9zxfZUtqPc54fa
7+3aNOnxTDZvi2X+PWc9l6Xgz0v8Tofk1RHROmcZn4c+ZinKJr+qCo89hEftsSLr
NIOKJEcBeeU2zwELZd5u2Lqjy5kClUPAZljSR0sd2pcQQ7939wWDUsBs3YfWxeE/
yqk2xW5gcd68Y7xQ6RIfYl+iCv/JWbYWLTXww02htZYR4VHv4Hgc/3HxgBfhXgA8
jTqJjSP/jcX6oGUh4F0g1eU5yMx+CiCHB/ClT35Ism55uHDPFbJiyu44jxoQw8pl
72Tcm6pOwyxytBpo01+FiyMgJqKfciUYNKMNqDvZuQitNYmdATCDmY4COzXgM95V
saVzx9Kd/NreP9lOsNp47br9vuU5OicmYccKkcWhYTOGWcsuWEFZ2g3giPyITyao
ctqRMk9DsZUz+Y8Kl4IU8WUufFJi5XRpEjRKsFosZgS1ZFR9f3SXwomTen1S/26f
daVSjsbHaVZZuWpV62XqQDuw//oDG5E4spCSMLAgydXVtE/COddO/YwVkBHObTsH
2fwqq0P8GJ/tEV61MlgmGIL2tqhdmG/mkjNtcQg7jWR8vdMjN4w21cw4wj+z7Qp1
M1pX9n0xON3hsDo9AW4leneQN2+GhsIPnTfWAKW8puwmMfI49dKRZd+hffFFAG28
1p7pOvLvqB3earKg0GoQq1PVqKxvOBN3HTBALvmo5YvPFWKi0H5cIxh0+omv4j5B
Lm4CV4qpRo38R4xmZbCXDrqFkhzG6aY3B/tSByJ1MEKP90iHfSwlmA7QPWoG8eBd
MRnHCW5MewJOUyifCEpedyXUDHDKlEYE++ATBDWjpmITJg+8yFXdMBksC4jCjI7P
xYLDp0dAqKSnoHWXbDN2rmKtyBdl8InAFABgMoa7tXzdeA1Bg0H7jgZIM02gRD8L
IalNg1pVl5oes2gVQOJTfsuOvbip4gErsqYdsAWp43mMv0QBZ2VgWRAamehJOBz9
Ibg24gsz8ayMSx3PugvicHz/nwntuEhe9bNqzClQB2jiLvw64iGPfp3Bw4YuvG7+
2vKvK5paatcfozodso3B8HjSWCdYOYpUAsGyZY9N7O6GcrsjrX3EogA/zzAIh90J
FoNu3PLlMAvvvCbtkgw3FUO9omEtnMy10lzQ8SNJdhnrIYsRjUZAdz83AHuf/zWP
EMy7rnLoGAwsicwR8l8sXNVrZcoJVM7KnE5DrzorbyOuRlSkAlA2+h+QbFzX6gGm
hg5NvgSxkzIRW3SnLbAmQ6zpPT2+zEuhFLHraox1YmYd+dCFJCliLZ2B2RILEZfx
TZzZyoyVAsvLKNDLWlVI0ql4qm31KedmvkslzlD180trYy3gVIt69nC6Ceg5Iwfp
RGT63bwBpIWMj1xpygW4zYVlABM01cTMDOHW9jvheJ8MRp3Sv2oZ9EJv0M/BNGhY
/ZSE+kErLZ5eZZH60i+nc5Dxf9MX3hHFTK6br4+wTKtJPOquXW24VlKcrGJ3FnRP
KSwNQQ9jPqkHjlXgVVffjQOTs9B9NVHr6Wuh7MrQsYt6dL3477E6eWFhd/qqpBIf
1Nhmrcq9LIHWC2DjAfRVbXSP37slLhKdTvH72odW21ALEN/n1SM3OaCo5aSMpbe8
86fywD9e84aWWPFTRpStID7baqs350KrC78Mn2zGMdrQQJLB9SMn72lXfXYqNHd3
NijDhDG3bjJOw4jg7edKO2mJOhext6s8RXGrVm72vnQOASfPDGrZD3MMRGIzKVnn
ydLNmK62IIqmhlTVzp/7JGx4mB74X2kqYwVXPZ3Mm187CmJehcCGfMahFveFV0dq
CJzw08LiMPZyUmU2TvGm/XvZ4Ip/hSa36QQJe0SG3x1RpeuSWefovBjCOZdu/MW+
nGmSIMaRDt1a4FnveBYAHaY6kYxoygfxVmzEI+Pids5gpCKef2PNKo2sFtwHXa7Q
qYiP8GB/CL39FliGDE9wq9D8HtR11L944rWginydsOfY6yzcXf3HjlTI+xAJKHK3
wFQMhougU2i96dhvaBTtTbU+yPqeG0vfnPgxssLwWcM0p12i5kwt3Ra5dEmMDzTH
uuY38IpVKSQLSVlkVjRTIbqg3BVXO1zOU1WDNYOxbLaycaWuOPG+SwliYCrbmlA+
RW1un7hPBx3osQCPY0JXyqh1n2OhtX3GOeAEDdgqGJVhIxhYlJQYme9q6DYSiPuy
5ZZAroraiBalGubLFa4GlJK9xv12pxVaDkeqn1cGQe0GmsIFaJERezXCSX7fbS7K
8JIPyW+wD9K7yjLUvEzp4bemDkGIxs3Kt1dRdCPzmbcsxDAHZraJh3DkWDvO+i12
nSHrjKrxh9LxV3WhkGSY0Efz72lIg814moVjvJlephnepVZfPJDPKHjSNvwFbb2v
uOFz5rYsHjkJK1xPkJmytKN1feAk2RB17WLnLBh5pGyGR08dSiN5TZgsKa8wKZg4
Hle2E02x5fdj/fk6YNLSvviO45UvRx3t30PuOLqzdktEw41htGnR+am1P5QiPVbj
U2HKt/XiKH30U0qhRxwhszn1m4bstEGmHMkUAa9az8ybIKMy/jlwVfFbevYMhSGi
MPEQ31/TVB8yqkBjbVi0FJ4KfccdSNyvI3h4xf/GREVixpCeU3loakIdqrLKWTf5
3iDPniwJ6PF0Dz6kgmBvHH718Kxm71VVil2Ar0t65UuLk3LYFpmmy+trXikGcdiU
2+Fb9VU7zT8Hekc2VmqB2DQeW0LYKa1ior/4EHF/uufKwF0IckPK7eZpE6LYC62V
o49fJvXw4u5hSaLnsLMsy5dAniYnuzR9LKLumm/raKDXR5L9JCxoWS+fIB9uX9bf
5sSG4hpjmJPYGixzKABaRKbSZKiv6xt8fqXjtWZ2snVMLG3ieO4RkpoTbKnRrYbs
yDMOSOrq+XDwr7/miR7BU+0V/zda3m5eLkLhISotlxApFNM2HgR/y3LWj+izAX21
bUzLHBmkpydx/51ky9EAY5zvhsGyCkt96yfC1NX54xq0AZkngD2qJ8X8u4IyfbKS
d+25zW39/MF9+FTEdhkEUhDltU+4/tU+FfYaVlIbAyY66y+i1PzJ2wr3VtupwzGS
/xqOOcEZN8REw2erUcGXrSGhXfH3gjs9Jwf7Zft/TXBctLMDxjxWSzGURQlyD+Wv
oxVKzcm9uljs/eGudExCa3ktypELpIK8pwef9Er8NlTVFYdgy+Hukrqi3HtgPq/3
XGKveaunFauFd+tVA2wWgDGZKuacECd78Urcoehbke55GlOyLgM6qXBTsF0xoW8T
GU3Edyoz9bboQ49qLAscQ+yL+ccYYl41etDQupQ3D9ZkLyFoRwzjz9+OKyBGEoV4
tnETTduEESG6g9qMAfil74eEP0+Uk+MDxZPWbMkupDYUGD3DbkSwtatwbHi2iZlD
IGSa3GgfOeajeQLml9hc4t/ONruvBKApoZvSNmoT8NUdTyaGTDJZCYYGX+qE4KhC
ZcdmplINmXep3mmPPqkOsa/4lCjRqbcM0cp/OujcOjUu9ZHBmUPEWm/+TX1xbkNn
NQVBpR7qOPnZQWDtfacpbTgRY5yxK/IsfwNtV+tooMU7ehhHD3XivE0okSvUyYT7
hZKSHRrtWqScCrMO97riP3PaIa8hM7Rs4JdIjA5/ZCJ/A5B7IJVRppc43B4UCWAg
6MIQWwMpQJ2WqLjsDHX3vqOBq7RWmdMzAmwHphRjzdRpcTGtWsWL6yvDn9iuo9fy
et0fZG06cK9DK3PVkskZc1tK/X3oNWKXPbYrdxB+pYm2HKRykrVGzFQhbmfUPpFm
MzWLG/pJTaETYVjC1oEl+cCakEOfk3ipO9/x0VWp/TFe0JlEvk4bccaGTROVzPa6
BXkEe7XaqQtmxgxje287I3P9bg8EjDCc87+eiLVsRkm6oJLUayl/kOiaSFGLhghM
mmALzjr2dtPoUUQKtq69QB644G7kDwSj9tet8XJp1MVk5d12b2kOzC+b93km/+08
754ikrs5XdcuoWOv/J3gNwm9fPkUP0uvlBIiT1x/8hV2swvwC+xu9L/5qy5lsCn1
MzmZ5+H+Sh/2NByylXfRjLuQ4Q2ALml2C2y53lkt0eyXtgFdi1BdA9mZUTO24F49
SXXBAUtlhoY+nfclJaeAzRxVRQVDvBxaZt40u2MfYAfgWqf+xb/45QMcu+VyERDn
NI359AE3wQmYJKMf9y9qDeOmewZrLQBjJU/KBq6x1HaMayvb/WXjKx7DeA4RBGm1
l/RMZ6ODBd0mTFFPNf344iDUmPYqU0JWMee40H2KK/wFyvcCEjZwsRSiajuYZrgp
YLeOO6xuKf0YqZ5nq7HKn9+W3u2Ucb+ZjfuA0pTCB6NTiwKuMSau9exwYUSC2YPu
jJ7LhVVqMMXVcr1TlJc2i8ccVGoccRkqUAbid+vA00TqkoT5mcS5SD8rajeTq+Ot
KlVDA5d6b+KMW7aymRhgvITaVpaAO5OeCAV7Q001X11klvlci5a46LIbsxEtIxzD
5T3DxPWpTVbXfthNY2g6NTg0ZZO7KG8j75VJKUMSnf64XzmrbJdPiqgmZqSdYrdC
nl0yxxH4qHRm9Yj2JlLq1TdBvlKGSJjzEGUcdtKRks/pBX/djNXYP55s9eTEnUm0
kUzs85ai1/hv8Zotlg8FmgLhZjHkDlLbdGvy2aTBmEkL4FvO1U1ykZ+jRFFLPt8x
s+PC88xs9ZVCN4cklSZlAcS8oA+4RXzN0Js8rPIpcNFWgmB0S2AqV63EwmFJn+Ma
xyKAkT5FO10GVuNxOvU2gmNjNYE+SSukvXsiDTlgj45SjtGMC02of/0mLEBqhglh
4dBaXGtmTnS8ouDs0/JPSRA+Z4NHTNY9pJQvTfVR+YbUyb7DrzPBW/DUscHj6oe0
4sotOTA1v1B6cJmi25o6jg2W2MZz/INfsEzOvRXiRBayk3XxzmWjWT3KlH9yfqEf
Xbci/JpTrY1+Z0PVqticpc3O887fthiM1rMs2oUTHj6wHiBsYOrngo8iroaUz/yo
XJKbP46YEnIrY0vrfoTocYuSaS3NI1xvUustPYZZhoJ8oDI7Qy/KoUMfYC6vFhR2
pHfgv73CGzTDzGg8a5g6KhwTwau+kWhZpNyDy/VTfRYaWYWndbFToNOyxH/pO8l5
t3BHFyYnc7pijF6x0G20H4jzP0bjm+n62Fv7aD7LXIy7bAoiG+dN3WFrs7V4wkUn
FjAmw1/0Io2Td0RIyM7j5Hgd6HBFqh2D900rqaGre8fqHOuyeK+aVyccLdxwcksE
zHJY5dIWm37TPdpu8PhpCMgrzVav1cx1bwmEsOeZM2D74llGmQazhxVFaXNhyO04
gz5U2V69EG7AA3Os0YDqaaySU8ZeJfShYVMTGxGCCRw=

`pragma protect end_protected
