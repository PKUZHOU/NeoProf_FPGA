// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
uk7aAiPMuyDG9LCBla8P+ykIQX7RSu2isYUY5U/a3futN/TrbfwntimOEjr1EyVPt6QY8moSvRtO
103vGgBWl0cCL9PTgN0X1Vf6YI3tWdHNNTVkyKsZGCxl287Q/Aataisx+01YOvBPYaZRy4vHejpy
ct+RR8Ly1QtSfbRxd9DZ+QmVcoq+N/3DwGix18LyYhXpBl0zMEiKatT2CQPAa8KQOCW2p3ApdiQ1
M6+/AmpJAv/E32vYoZdCpNoYKoEcSIG1ia/jQp2vHQnrTc24bQtcDg0D1fXq8bCEzAICxTEnOYS8
XPqu+SADm00pT05/xIPP/FxVLgzX7a6TrWRIuQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 8496)
lHYfVh2KQ9A+CfekPY+zx3pU6XxlpLK+8b+uJiAqwo6tHviYVAWrqxoho29TnugT/9VfFj5U60rA
50nKvx/zzWKTIL/wpalOkaleWFS8tt6RALH9RonUncyaO/4nZDAjMmSUkJO/Rcx225bXm2Am56o3
LdEeXvY0IarwIPVlsmrVb+Lz2UcaFxb/y1rgcJ4MmKtQRk35XpOQHHfzerTuKrAXPYzZlcLM4eL/
vCPtULCmxoBV7Puc/uHPeHTGKF29iAlI/0n/DNz+1cOkAKqe+EZ43QDTUEwOhqTn9PY7MlJqdc5Z
vbaBGjFuP+Mcra3cmW2BZQUQVJSrRL2LLrM4o4FpGeheuZd4bNYRKSrs7Ulph5l36kIefkRiTMyQ
oYgp1qOykqbDN2YJZ2ryNu8g5rfi5Z9sfmHQUVwc3YaHDSdf7cDL+SGFtrKOER3obIcCW2eacXni
Nc+YemcD6cikDkiQHeeo9XFNJjDS4g7cgPQF/uhKuwXtqRMn7WkJpMfMxtk6yhnAfdaj/GbdSVKg
uuw5udAho9PBTwMAZMoLKHUzd8+EGKr8rcHGMULYk9yVZCM8bHRmcsHqgAsOIm8jqdPcp+m5dPTL
mTP84L6KzXSjbDCvanaA25INGbDjVsCvy8k4aQU/g+F+ekjbPOA226FOvlliaP07HNPjva77Up47
HKHMacxZwKdqVRzndN3ZtM732Xu8Sl8aCALhN88b3SR/272sQBp86Ij2dSca0ewvUa+dFZdFc8O9
qKmYRDwtgqaEE+0nxdFwvvK0Ujj4lR9We4LYMlf25ZSAVa0tsnCqopqanjeE36QyvwyO+1Yz5shh
b/z/MzThPfd2iQ3D3L2DBaWK8+/+IUmN9wP8FUJ5gqxjoUamoiCUS+ko6KOjImXo0hs5JZ2CB8Gq
KHgfRWhC7T98jQYTcLxFhQY2Y2MDwrmRqdWAHXYk+qXzVM3TX/+hELt8LN6Lv31CBHXZCPBECl0T
3f1DtC4PdSEajFMh4d31JKJ4j06FklWdAk2gyQ8hr3yJnV2l5emkCN8haMFSmj9n0SXh6ip+D84p
m0VTXumuHRhWdzuTEPAdnCdYKf32w3wiQz7SxwOa3sCFgZnfxIWUVga0xrT8PMniFhNrEP3iEYtl
UHUwvpFuPe9IfOxJcd+Qrbc5xTvLxFPyboxkkXfUWfm7CKrtOzw+jvIfVHSnyvg5qkzhCcZJMMGP
aKTuhj3bU4kWj5OG0Ez31CGt3TwFus1BZ2iFIFo9hwiR6thPfguSSM83K9q2Cv+cV1kbfPH72K7Q
AxUQfagLpUi8r5Sz7NZbmoF9LIObUvBW5/mrBJZ22+ara1u2fMjuNh8+Tm5luUqOnYG6MFBpB6S3
za11ZhWgI5ERFXA621JsNBhKJ6uZCF7/H7bBJbTTj/65GZZwM8aTkmOs3CvIMytBP2o9MrUHV2Pi
LmpcU6xhGhuclQc8KHTOXpxh2Kc3t8zJ7zCmk1RaUmQ6sdkroQh4riLj4lFOhpu781KqDtienek5
UFlzgidk491duf0dcwFsACE9dtedbsM6nTQ37aBDI0/21+LXFNxGiENyzIEVIrN2x8cVj+VUXY5b
lkc1OD4Lh5gDNq1aTIFNsLUlSNmRVlVccfkyp94yj3nzvwP5cI6uUzMsiOM6nsw6H2YIgTt9/HmY
wRMk1ZptRm342+o6uyiGSqDjTYgJ5kSVir/JnlWSZZKcU7MTpvr0twqfNVRvnnSpIxBt6EWfRs8N
rIPVdsbK9TUHnqNNC/ZLlvhlhQoGruxVnivkkqHjNIBdYQYWsoRWRNkIg/bD0g2SbTjl/kfI2sec
px/vnLc9TFS8+tT1Z3D0n56IcQEclmGmJWMZG62Z8Dz7OupLstdqEkhFSSKhctENGtwDWrHUg8Ds
178y6fBE3vPJDUrE4jNoGx2JmaC2z04SahQ0DpsE1JHP1kGS0VciXFFDBuEEcm2ilrIdXGP7yAd7
n1Nw0jEHKcRk2NPngCDe56UcphnoYe2lC6Ky5yRz8sTv+CXZPJh+zk8MqlrrzfASxFSDenzZgmi7
2LJA/tEAP7eoBNk+Q8gN5MR/DRWLtTkv1hfdGlHmYEPG+F7aWf0bO/M3Ovz9AiaaCBYMlt/soIPw
VcQuE7xX+7lhbxwQsYc7+UKCMjRL7nvAfu5a44O//zBNgO0tOTpMCkqPJLsQSZue7XEtUqkJTpfx
xtoLeLElPmHyxz7vMrjEMJyOECMIw+YvR8MVPV+E6CFWBWxNrb6fDl6nRcEHdNTffzYosudoOhOP
GhpYG7Y2F4PZpW921EeuciPcml7rKCzTEDyGjs2DxRzLwMNh97D2SjzSBfNGfiIK64DyyY78fjPY
f/cZ44zydCs+5dPNII2ZnAAEOyVEPAyGx37i5+Lr7BIbo/YyxaTXjUvEuJNQFFjliNcFeBakN3rK
/tPXPvJQRGuDf9D72NF+vyxqVEbh43Dpr2CK5/Uj5zBgrRrg7CNJw0G6UWWAir0IQ2aAJaxM55Ca
5qxcEk5n9olELGHo711KKeEDwDiMVc6EmqpqrhyAHgfgTcaedQ0QpPwgNCTI+kuV9TFG48MY+W5A
Iukg+VOB+6r19p7+0u45J5O/0awilQ3se0dVaUW+98y5zuL2/ySdXTogLP6hb341GYXJI2UU5Nq+
zb+QiZ2oWvaW0nM7SEk4rz5uSTxt/PKY8E17YBZq/62Gm7NCpPnN72NIrpEyCzcjwplFZ+ngJijl
GdUEdTdehz2M+Qq6J0z40tU0jhmq+jG/ZsbcBTCJtCk4+TFPA4RAXl6xmg1knsJmh+O7anwz0FpB
x863OuvMaQnIsfltehjo2yEyNdjI5pmkT6z19MBSsQ9XLalLyI4KZ3gqdJdg11Ics0ADa08TgJtJ
6qdxAaHbyRKFjvKPTatsS+8L7Nnoukr48gPspeUh8suwrz826tMVBx1DUSmhOgklmgjUumx9QOcU
u/P0l3XJ9oQyiUfDiWVvvYgm+svHpB9WeKvTvQp5NrqY2JAnPvZLNW5YTW5GBgagLGGmw++nLh46
AXIFeUKjVkGYhpeOkFAx4/ooaAok5ixZTBn1nfNkVkrT90rSDGsCnTJExMEPy8fk0/nuLTzvLOXX
TdJvYtqfKCcDzIdEKllAxKLhyZK5Xw0qGZFD4yJYa6JKgKpcFlPcKDTYJnyCU1d2yFnjyS5bIeW4
XOEIJkagNqE8LTzwuBEOHmqEiE95wwvs4I0V3W7GMwklh1DWjeS6hkahrlKGZJzz/dWgdLoa12lt
foY0Bvydl8zmu9IUMyQFvrifM4e4C5TopyxE2jrYh0TCOxnhTdSQ+rx7AA68dEsgqH0TbU/0s4Gc
gUTDXlRYiXDq8qacpiM/8iCCHL43g6DdGw4nTrJ52GWz0JEotk9JZTXT1YowrN/dDlxOtoRpV0xB
xnnYX03AOZqF51Qh3FWT80b2tjq31yT2wetsQk6iuriibGG/iHsqdvUL6ukMHaeaCMFtDghaO8sC
fHgrKuya1YpDK/pF8s/aenlczfKa14MG5fOenI4sgbc11yOV8aCtleuUMHL3gydydRKkz8vqxMVY
ZrB9YmlA5VXnRR0GwTI+XXGrGd8K03oGKi6UQoK0EWb/veuV2ELOFKfY7P2WLLfckzF8qYAmorhG
v0+ag9pITgJBxtJRiOLOa34PR9PlzdYtYxoAxWMf30Mh/0BVgsPGxc7w5xLahmZspYw8AaEvN8Ea
VWrfsdXRyqm1GtxkoeObotTxoyZLwP3Ukcw2zwOqTxULp2MsEe+j4TxjHGIq3DgrunybVx7zFflm
cNRxLWtyNkMqru9bPPFLdw9M/6V/wJLubUI0aWQ3YKzHpQXqkdHIpuXfzrFY9f4XRHQc/OPH8pNu
tz4GPy/f+4oShFSMnBuEbt3srTCvlSUvUVDOji4Rh46Wz8oh2iIEJx48StjICLqdmIXHcNE5FD40
nbydJcPzwwnLXkCq54CkYrj2m6cJehM9GVW6JLAxFlmpWfX1P+VXwedopcNk0pOnRzRCJp8dzOOi
vOUwTshgvIBJ2z9wS663WThlOmbnljgrHb8ZHqXgru0OXkTsoHhVqiiVZRtQQ4xGm4IsrWQg9ssV
fFN6ybbH+nnj9bQ+hWmZmk6iO/q2gyiKtcklxV2y/fWQX7bqf2pdhd0zh5IcCsPk9YEGE8J36bvm
JGkR1NUC0uomjoIeFmcHWI21u914nJw4gW3CGbEZhsUsiixGuvsaucux/1paDkYDs/8L0fSyrG2X
nG8kQXRumo3fzm5q6N2tDKCJGP4T4tJuFvvlo+a5pxP+GcIR9XuDbAt5ufYpPot34Q2832MGkDX8
KGw1dY/FMdU24YCywprgYxF/0Uz7fGeqe1XHh6wHGKnKJRNxr2v+N8WQg6/i6dBrt/GQ3krBPKkA
SIbI7vq7HkZ2G031bT1tt/9lFymbUsi7VD1uyLOmrM7PniPPPPVmPkkZWCDTF6sKTY0Pvdg1xWLn
2/lUW8wbxDUTevFAzHX7Q/+IMEQaPV2M7En0WhBNK5IoI82/9oJIp6/z2AwtH/QcVaJp7+QtR/g5
7JGiVe5bKuq4ba8qBZnTQLNeZXusAePgk67PARPlXF0dtL9R3kIkpBWYOnnbAA+S8o3Uckvy4mBV
odCmh/3ER60tEX43/sVZ6BJyxBg5IKoLOMN/NxaSE/binZnnI/kNEC8lgyEL/7U1DlODRqoih+Qh
b9H4YlZn3D+8hV/7z9mqJvlVY1cbYg8W0q66oz5gKWGUVGaWtIk+u/Wc/DBbvqbWn11wCphHQTCz
xjpTYQIpbOoMhgDNj2ekQu3T3GO6TJpfbeJH/AnOVGxNEzF9/m/SzJP/2JN3zOzDpQ/LaahFXT8+
EExcv2FOc64VOltMcNOQ98F+K8y+ZRCeMNEYt1hDWUhoXTk6lIA6oOEDj2CfAMozkUoS/JAHZcvM
ZKa84g4n5F6qicA0jOjQpOCWvhszEGNuo6KrasMghax7ZhEisAwkW8y+wsZg8pj9mDPOTn5v26fj
haAbFh6sMMAVakr9aNb7+QehqNSLD9d/pBD5xLjv/SyE1rXFE30bp3oIt0Pq8PHF7A9RKff+7G+A
hJ3Po8bAXxGS4hk+I2qGXopBE82LgN+3nhG0Fu9PVuFfr0sQ9qLOwD8SZ5y3AK7pr1cc0cFfyEF/
g2XD8eSMPJBUZVRpdX1Ixd1ASebeTGVpVN/VRtINIB/cmVCVtIftelo9p9FsCghuTMubjXaY58Mp
luVqvWw0g2xIu3cGiuSS/V2wDDx0X4iwRz4hGcNOi5GpbVeIRsdYqrTk17lYGASboQtMvI0L/IPQ
rbGhV8gKIH/bTqhRhfxs9JCQV/6yOMma1Woh7Dpm4eeEKPflcgpBLR3e87pVZHlOgx6+76o8sHtB
In3y33C8fmtHj2I/RKZWRgKueqte3tr/VDMF+PsaBuTscdFTz11mTOAYNgVkAh22Nfcht86P/zKF
PT50MuzXhRqawrDgvHx9Bzk1k9bysfEG43F/I6SNBd+J/2QyBSFbKxgRXECf9zzxI4Zw/Kf+VTX0
i7wk0Ws/E2KQJo/9oxdF1uZe5T11FOqoX4ttuI4Zyq4mtEngda/oUfdU1YcxEi4Fr6Lm4uy7Snkq
YwvdgYB5b7UlhhbVsACMXUIOJZZ0ldlkMES0ApN/JQcew1SClvxquRIrqAqEG9Egux7athk4nCeI
/w8r4SwMzIkV+PyD/C0QL/drwIza8tgTv8jCUadSII6SOOeYuEfjfkwCLROa2aShb6T5xLqQY1jV
9tFhuUdP6S1NKjFrkNVvcez72bKBp3a0XTb9WOg+32bUznYb1xtIk9apRJYDCJj1EGakK2Bqv/8e
fp0o5zoFlFQKi27cJk/cNPSi02Mg6daYMBgd5cwwgNAqifQuPJeLX0bp6pCbBPLJRJOkMvMC3IFf
aWCSqMjj9NV5I3gJ7c+NDcwvdawwDTTRnMWv28YXUJs92yLAABKZKNZtI8kGKU6rh9tXv/BIv2zL
dtiwYZDOv+/WaUftyo1sJz0E690XuewRZbG+eh1PpuDOUuZ5V7tcjbYbSd1ZSxk1DFYTsNVdCwQQ
oHHMQA4MpXIRtzlmfujjW9gg6Tymwt4vUbAKNQyE1ILXFFkRFhlH7TgceWV5GYL+ZWOQuqPyBwQj
7FyOa2nS+RURMwvVBJtTFpt2AZdO2CrTN7czGZ4c2cHx3rGdQDDrRCJ6i7dOx8gtNWl624rwWUxy
ZLyxV4QfswnTloqVdsfUOBBbbOQq1/vqQm6Kju2R87fhYsbam8NXkvxNsj42zbtvnAfGFEWzyRQ4
BSqXIjAaZFL3i+CuWueC/QXtoairdhBRMV8cYirBd/2TZvzoXrvCo9TnReBQ/84D4fmcHy6EUHQU
D24G4121evQ/RU9iw46eFUUbQ2aqAMcrguBOoNBu5HUQrbF3uDk/Whq5BsnVEVtliDQz6CZVdy5o
qtbreFw9/H0OhHcBXTu5b0mxVPP0LH4GnbpYeZ8SCZ+c3gISPw4oa8seaIp78nLWil5y1QVReMg+
Z8bmHZUDcGFisTi+fS/XZDQI9uWhfbtCwvsaRfRbpSjcBdhZ2b88EVl4spKZcH4uFqWmQc15VFB9
ZuCNovvBJDF3CrjDNiU4K38BBO8Nku9lG+xo1PTn8vUm1L/pihHLwk1+SiwE41rIK0xE93viDso1
edUD/HeZLG+ln5aPtjpdR63cWsK16ZkKM3aWo0k1awwqyBI2Wddt7twQegCd/SzaDGG6giMKAEbf
Qedcdxnd69nsFNIb7CKKr83+3OryKasWFfQULxmOTpAnS4HxN1JqxGEf1orDQ2kChutObWsqNzM1
QmLVKzm5jv+LmxjCZlV8w2LRFINVNiTe+lf6xhv0eeuCRd4EqozfTHWnU++Ha2AKcRWM5hRxHFWa
/Jtb4dqSYNYu+UY+szkCa9UcvRqjvievAQ9UW3AtUi7JMRYnNx5QT+9atdinxk+ZlukVImwuGsYw
dQplaFpRll4037V5VlWhqIspac9Po0ffQxs6OhZpcKs2phLpCySPaqLl0u5Gw24yt/kGfG6+UYQJ
Pgj4pU50vKJTrasto0Od+mewx2/TRlJe2BvKdbhE3en1IpyT0HmsMTPrdL3vm5qq0BbPTBk/ohOd
UJy13iFV/EXe2dAHctMyJGVvsqu92BUWIzJenfFS39yz7is8M8dOuYqDvt4XXs4FXnib3HRfmv5S
eVSXx8rgatvG/rOSPZNj3Wp9EoAW/W8ki3SQ16w5mAzVGFaICeJO9tsYc4PQhpvSoa3K5zEGNkRl
2rbyd1fnImYKoDy6DhOqSQuVH2lQIg1jWD8ap2FSDXyF2vdZBPCZPck1pi8CI+Rdk6FIoZDd91hT
hNQdWMoOqQ+6+st3XW6SbBN9V02dWoQWZReMMv1WEZJ1Fn71kiHM8H5PjwExYSNXNGqvvSTnVcxi
Mujqmh+3Pz8SUmtpxY7BjL65cO4gCzpqo4x1XUE+SveUP9yi8fa9xJq1Pwj0sjuK0GNXpCdDlGUW
1IeDkmexYB/Ewla/mlvPLnGNvFrtT+EAD/POlb184pwmgwCggMX3feCAphjv71WFa9OllqcD6krX
YO4W0YGerev86ITBhUcikgIlTnvJM3DBLJB2QQl+mm1LTuyNzv82OsG11Bmi8uRrBWlkJv79YxEz
mpswH4edbQ3vmn+J3iCIeYDpxN/SUZHtFwKcOm9TWqt27SfVr5ZktbzuY1v3XZ056yLizAGJnc1K
YjPfKaQIjuoBhAqn4Jz+FGRVQPoPn5WlRDhBIIhWdUUmqo+n/gUkxdGghVc9pDwnXiQYq1GuBqRC
kFFTap1Jb/y9BTohrjLHCVcHnHNAtcotBAQb7IM3Ib8ip7axy8Zk9DBDJpJ6BEdFUlAt817pM3fn
mQ8f7sgKIt1afbbqh/WmOA/AntKPbo0EkLy6XpDcWfgPFahcqK6iuKuTqNxSiAhLm6r3Hi1GJtKt
nDk4ALR4d+6VQPlFCaGUaxs6AYPVn9gZNUJr/D4uSl4fk8PVAzlao3FTayqv6k4IuqosUU1ZPBFf
Qsm9+9H6BU38CN3mdM9coQTa8WPgyMcskN3Im8gqQO/j5wUhwMe4O56o3eMXW6g3HBD1ejTw0U3/
9PiygxM1vXmnEOjAQMI5nuIEkIE17ttxXJkMBba/BB0rVF7hn/0gOAApU/fOnIBZPWMaTJ/YvIl4
MFuIIn73FBV/lH512cQMKISTmhAoPt2KP6rq1kj7S0hg8qqEzbUSCpFN78Wj0lHqwrzgY+IKVexT
dcvYE9SMj5SZO75wY3ZZciF+w9K0yaU/0GPjqblRrNtgOwMxb6qm573QPc+F6jHioSDuAh/qZ1Zi
CFnOIXDUtBSLMyqsR6atZwyv+qD0zDMfZcA8f3HgLNXTNvm0wf933WQsj8oA+U0kBcSqk10mt2z3
nNcyKIoPklo2iXdtxti+DiYtpJ0K0bknntrsqNSnvP763dBu3dsYpaMdWJynP3i9PPC2ZEi1pwDj
P9uRF5qjHY+o7Eh1REayBO1WU/fV9ZSAtPmpB6S+DkVqi7RQeHorX3oPfDIyYfSgUivMPGZh14bl
3WqbTRnDnnJ7aKgW1JB86elskwiq2i8i1vp3+JWO2vrST2iOVE4MvyEWx0DadszZ5LIDvwqSTXdY
fOFKVnM1r/RJXB39wcAA37SCW2A3454NuYJpVdZBGJ89TUiyQ7KsSYjhSRJjt0ggKQ6RyOeq2stS
SbqgRfeEkgX6ABDLE/aVb8DzK9o6Le0OTiSSnQfhJ8Ys6hmZWlprK+n5F7FhyLfM/0qXubjk84GF
VD8Vb7cPlnv8VKyuS7qnDhOFFGF+NqUtiH6u35+xN7qmGCQOLJd3a0KpMf6G9s1l+7+Z02Se/ePY
A3BuGeLjKa5HeaBWrYEkBTj/MTs899ngy/9VXC2068TQRbVIvyKjlrSSmfE5FAwsj9CGBG1lTZdO
tFRSygr72CH1iGDMzcez0KElXVvuydES8MfpByy3VTBuXwBNKIRz2NeFJ73Qoy565rY7FlfZ0/7r
5ku0InHFfjs7vgTNJPUWOV6hmMOhSBkFIoTG4/RPwxEHEfPDof4VG8STknBPQkzOK6rRF+hUb36H
d7cVzOjWS09t8taPbCF5wwlvX2Wp+Z0vMnIf1pbY7C/ZuVFGx8h7RfCiOV/ysoiCzVvCys3eUtUz
tvSq3fYJ8jQGI1h5U4Xzsv5L7hszxM8QZ0AIZe7c/NPoXcHV0OjZLMXuaqiYPyNNaQfYYxCyVPUr
XZSX55U4c7Pko5m2eQuhgUeS98BHouRz150sRLjUQ4L6PzIXtYVCSSQ9l/L47/+SR3DNcFdwyDxa
/+RRDrd+LkzxizDu2wZsQwdaUT/OnnkQ5ig3iqCc6+NDX0//5Rwrl36DQRzNeGEQeBmmCOa6UNTX
XInWRjuVgijjneHMnnnJuZroylSA4sMjPTYzMonQXbdmYFfuLO26r9SM8e1AkejFSh8T67NzJgYm
hAcnokeWShEismbGtPBtTibZW8l+tH2o8QNvV2sTJvtkMuRXz2AZWq/iaARJmTqcVC6zZmF63Aru
hzcNGham1/g8uFAZNY+2uSWoGbGo31ZocsgAnFAcR1ervm5rfdPx5xDHf4BBFtQrwEs0M4NeyTTx
HJZ4xgMCn0i/xvNGoQc6JGq4o/KzuAxXvTE7rXdFLEkVwB7aMbTV/cK/vpwwvj8jxyc9YleKG2h4
j8qSKCoprv6BR8cRx0g/FRhMVs6prtEasJKj8WVmhhC19PZXXVaidBjtLK4YuxqG9cwHHm5cVOwD
Bt0VfnFVMZ/pOELf+nm6Ws5aHx1rRV8rJDjcZIh3HCcBYUTGv7Rsd9cNzyPgMRKcMMBr0/QmXeWa
sFRMv1tAA65MElziRobmujs65cjL41rw7DNeAz1Qt7Liqj8oCyqVKa0iuZm0d9wqgzy4P1pwI7JZ
OH1Xldtj9RV3I7d9lg3+gRO0l64l74gjdZ/BTIL2WSz7ndMbtZuBIucKBm++PRaq8nGSMiYOdvOv
VNa7EGlV8KQv/D1+/Z66hH86EXD/3maJyp6dtutVNoOYHQn+859C1svtxy7fl7kWiZ5G+Zx4igL3
kopYQYycZrS7AlSrjWaHl6STj0LrJ/RkwZpAT2SmGXmCoKlNWYdjcjf0MpavRG0dR5o4P6TTSpsq
XWfQ18lbwEBXHG9K+EwmX3+egwGgbQvQJytefVlMo3QzdPe65epyc/1AEhzmxg95M9nhMVigyjl4
0Hnm+s9vTeEhtorkJ0i27QPfOVQCMc92DwsM7kON/WX36GdYz9S1gG+kBWdySIZsS6og8d4CM09P
ZeqEuEgy1+VujnGvm/h+gwI8I3sWZ9IFM9COlXKlndfuXJ0F0EisZXCHO6oN31OH1ZsvmhQ0s/F8
umyQWa7Y7ocAZF0x8kBhrYPYM+YcdEUTxY/YVDkvkQ/WWpsugbhSagZN3KVrtWW78pkd9LWs8BcT
TP74SVdgaNv/caIRfQ8YlLh6J5+YvgUQOaOPOsmyM2qQD8EOAsSd+XO0f//T3ZAlh/dlu6/gAc6C
YxtsWdrMSs0UdrMgUJewEqQJs9vwPNvT9q0sU8tpEO8gqGr6F+dLd8c9hstznGXGKxbF2nFShNZb
bDaH0UcOHV+A5IvJeikx2/vNzIuTImLecTcOQqkYlcYvNDF+7CoiWx6ucGNaNACBhKLlVoXwHRKL
PzWXJ8yxKkoF1WNkRsl+JLtg7ljB/cxuEvr28PjLBju/2KOiav8WpAQr5wwaPbaMStLVy1canle2
bxLffgaSxcWUPnUXq7Ny7/CviNEJ3RT33dg+8ux59AZrDyiy+OMbunk4ME1y1R11d3LCT0Rkozqa
HSGVKG1IymkbG6Y4bbCB3yRT1pO5qkU1vcpyiP0cJcZjlGjvQIaTiP5I/+e94tOrk8bfy9JDqFF4
sU/H6a6LeG/VRbel2QKZXOVfH52kmoEep8lSNPuAnBcK+zD1MwGklRLUILIYsl5oTapJpYu1CM2w
2wWQmVa6/qsvtrCluoYDwiads5TOjgb8eamu7tFGIT8Vb2no+tQpr4hWogUnJo+lye6LqFCYVi/J
H6aMSeMfzAHThY7M5M8bl74BtDpUEPWEs8pKV3leCDJWTagNN/yPm5gSLZrN/AryozmKaxXEM9zO
yyBJQrRQgvfXlLtaGSM146RKr6M28EB2805OgzHeXAM6PrvJ+OV/ihfmh6uTZ4g75bpSKetMINZJ
uUYbQ+e0jOjlEtIDzZCjWgM0bUkyrN6dOCyWtiAjq0cn2Y8na0APEyp3NSqpQgXDydAm2xsZvVjf
qFAQ
`pragma protect end_protected
