// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
nnQws3BvAxSh4Gd8xSleEPMAkigBX5R0V1b/YBJzK6J+BWats+ZBQLy/fovXdCQ4
iIBV3/6yezCTFcw0hfD3jLJfyZw2O+5RoPhvicYE7RSUH2M2+dWWUVG4ZTc9PtUr
/EIT+PSb1TQxqqpnGgKfYF/ye1UGZtj5DM6O/AoJbiCZJGhW1DTPJw==
//pragma protect end_key_block
//pragma protect digest_block
ZK8QFseebXnfRpKdQNYotpcZsto=
//pragma protect end_digest_block
//pragma protect data_block
dEYwDn3r+qOQZRWRro4UKaZ+0zVw5DQ1eygX9U/AE4y47NjX4MOHE4H/VOHe54JG
F7WGaKKYWzUhbsKMJxH6P6iVvA/aUSiTY5MZ7Ee4t2r6PIfytlL0VFpJMtUjhbAT
08ahnBhHOCh2wsZ2zdEB3mZkPCo77vutCdl7pIeheVXXHKAmFSkTRDRAAbqNMNTj
rKz+uqgwAS5PqXmnm3PmgmgQlzMU3NZTnKpouUFRoKyD2fytMUBbu7VInp/C2mii
H/ZbN73jj14uslKEG+NbW/IKO81lU7bJ68IilQ4ub0/c1ASHgG23ot+Ebc+nvKyC
1k6B2uqYLPWoq5F/J3TOEwJ5aiq0p5KNZlQ2E7zOVkrMMXx9sCqtJSDJrIxQ7jK0
7aqRb9jKfFXgaxhieksaWbcZ7UaJ1cwEqVKtob6OFGAASQKajZOxmE+S8McKLWkk
DZ5e1aeXI4Di0A0R4XGsQKItCu9YSEP+R+VpqkKeUHPorP/SYgBAblB3bOuyVeP8
i8/VPOeZhBy4VUER6rNtkiY14kqfk40wMznF/EfmZ+YsgoaR4bvKPi7VyRsvEqo/
raXHxxH2hVbtieFLH+uKjWKmh1W5XSSXkSca3P0qSO09XYXiYQjW9NJY3k77+5iL
Nid52aiv7unKJV8aO9u6Ukz8tvIlmBHlH86y9NHJNfvxvQzjbvGXNYBIXlTdlkJd
xJzx2h8gDOl7mrkDoSgR9SBMAsrWd5uJ3kYJvRjX0qOoFy7nD9JYM3Cre3PUD4wH
WoF2zcBCeFahb2/9cSAJLmrJOqu3X1J366bcFkupqxXEArVx0otSHqx7PMPYeSrO
U08hkjJgaIVMULTOJT1tRfzspzHazwYFMpwbjhdmcQgd5hqvusz+AExh5/Fzs+IK
TnRz96yqRlQclcTSwie54imYuP9ossZhxn6SHwVzH0gycsU07U9wrRnBbdGCfXKt
BE1/l2YZNbDGj1YPLKrBRfL43BkCniLLNU8fHyvSF+6MYO6HeB9FQzkvYcaMQ5N4
bvdYPDuu00V/RSmA+DeLFHFd8gnP8Q0KoCtZ3hq6kPQXXnIFx3I58aDPhYr/uqQj
Ni6ux41ZHfkSswgC/j55/6UQ7PFUXK11q/WYCnrQfZ8jCucrTQkIu5bUNj1Sr2j7
ot75ubtL78zgHqCZDvQkQKrYsZTFa9hfi4celqa1dOloVqAQGtmHlYC86qyhnEJH
6ZEFnpmyMGPYk9cHS5+ddmSwYFn7zy3qfftMdpp3C/Jbau+9noi+Wj/5hWwr2xNE
JrEjX7OQM8Sbnzx0BwupLZlhSpizold4BOhm6glaATltabc1HuNq+l0P3h5woEuu
PwGG0foifJf56UFIwOri/oHh7qNx4FlUlANsPKLUoaZRmfyZGrUcpJKkNGDgKh+C
QBHczg8nhQJALVZxZQl23BUnt9jtWJACs7HT7N5lFQTp2BiQ1D7CSBqrYAFA2omI
S7q9oHomGIBzbiuO5GupzGiqR8n22+eq52iZh4Wo5jEwxYab3fo0SZeAUzGXtb3T
Rkp5PA44JXeBoSPxGqd6m8M3Z7kyb0viwXj8z/pR7IVhKHLRvDCtJfVXkaH1G0+w
z2gDujHJljjpp0pRsbFvdTbm6xPxrvZNr3uto90ta7fjsWXT1STbvjheOLD+s+yl
y9uJJKD5jNFuQ028nwpXNfiDSNslJUp4nQnZm0d92N3gU8sQ00fdk1ZX+QaqPzbd
MGeXv+BLJzcoXgX9hcPX6zmHLk7qis4BpqdZph/SHdtVku4edNpJMONH4VQHR2aF
oF2IcwRMNgtTsClWyxMKskVBHcfScf5OSKD0CgZ/9I2EWnRY9FMoubGtszohQYzH
xgrDBzSZO1LlGaZdquh92ZO04JQ5RInyL8c3N/kh7wmmGfX1PeLGHnxvwU1P61pJ
5d/QFgrtUiFzkRagqMeFV6p8vzg3tOlaKvejLuUYxXLsaRCNN0cRr4vexvUTxhXT
VQmBnbuRSEri8SG6zPJOX0gonVJ8fS806GrKdXMKeurB28v90nTG/4O3x+mubTE0
VG6qgsKSQaR/7mYGmFmBxkaRlfNg53ydF9+116JEfnieJC+5+lpHE78pZ1+Cigdn
kC5RDWCY1p/nwz4TtLeM97+SmDE4NuPMXgJOGN0jVz2V5z1kwnhlj2yGPlZoWS0k
RQVWeIOni3uaX47QvDEcls97JJ51fj4c0TJeZxLrE/Py9xRIFSwBMVeCvZpEqeiV
pDaqHGk5KEDVTYNgq1HBulClCUyCQ9/zaaYIBSrlUftxE705ouPLE6XDTTrS8pF2
Eu/90EYxcjMOOyj4EY1VEU7nqZnJ6/+zOCGNjms5RxvJIWKRVtfYQhI7RIZxrjFW
5zyS7C++tZ7NYJp0r4I3RVvuvPWjztFl5+ziZeoHRKY8xot6R9c/YabI9iYbBwnx
L9VGMepFa3pzoQ03YFNSNMQdxxz7YVMMVj4Qjh9G/Z5eabJr8G+Y11ikrWlq4uY3
sTASt3roSO8vfZwY9oA/WPGD+T8/2XHK5F/sSeYEhTUAIXrUZxayaX49/fCPD7mT
FoNwiK2AezY9NHU1pSP9ry17oNVb3NuHvGeff5mfGUBIE2oka9ojqZrFqsK+id/l
csaUMz7Pt9RjQYtT8l0Mzc5dhdrdFC6+K4DwBQZP7RL9/vL4p+QJrPPnst0uho/v
zCDt0KKouDlg4GkMkoutgjeejqyJ/6CqMcu49js9o7f0HlsmmTKB+p3hf7K0doNW
CPlGbBlyzMoazGOyyo/0gchf2WHXWMaSRAvtMImcxxF8kh+BDXTdN+Q7WiwUqmcn
OupMxn2SpUkJQrjKRmrCH14SE0+2aIA+Fh1txURdo+mnKf+NJTJ2GrHVlJJcH9OV
m9I6XLoVdHpUTeBCA449PKh+buTpWDambQMfe35iVGlyh8ChzAFwWLnopE/rBYaF
zb6B/pJdWggVdcvVb2ljor4IR5mUwOmv2agFm+Q8XTK4VbNqEMmd2zWHjAvXa+cl
iO5SwDQkR0Sd7GV8KUfMfc5BX9AAjhVvlUPlQ0hWXMBlh0j+zH57NsHbfrRhNohe
U/7Nt3gsEb0OOyMAMb/U1KCN0+VjOYBlyPRp06NGAdTu2JXkW/YvCk94zy8ExgbD
W/IS3h+bR1NF0ZIr4pZZt/PI9M2p6uoUYs3cI1Cwj4wiAY/LMpdO77SqEXeLxarm
SEzMpZlefFXtbkB3GiH2Fw0nOtNv6bZS2WbX+zqNRRs+HB3Mrjz6KgG2f6bTXfax
5DbSlmD9UkQBeqCbwSEm8e/wfp8GJk9NGllr+TDje1w/93gdhpfHD5AYIiC0zqOP
PiOuvgwhvhKgFS0B34S9N1/pajKI4mP80inGYQi2EYBYpw/UzTMWMElvqRopDsn1
iHb0U5RTV4PE4mGNS2WwW304NA3ivGAuMrzp6KIEknokDgWeVp8XSxDLeOZq1mwt
mfisQb61cTT51GMBjO9snWto/WTOK/fKti5eaJbexd3Cr1G2ORBNSO+cfkH6D5j/
M0KhLO1VujNmTqXMdDg81yiDE56kX2X65idFAoUnQ/Bcu8y7ctYBROWC44hx6ubz
EJWaveBkbuH4640M38x8Ls4pV85tCAFM3mw6EioyFsLAgmkKdPq3qVPlynOvL0Au
Mrh77VGnzvy7qheG6QDU17ZX79SmmdksDid2AfSltsLLq4qjtMHyqkZBop3ezJ/Q
U0P7pwfmX2bcV+qXYlJAvirxOv+Fy3niRqXBT1bIVb/Sdaw11Gr1M7detWC3BIer
n1ZrGu81AZR6bw4IAqvT53yu3kb6t1GvUMD/nOaZJv+oERes2NqKqBNdrMw5dihA
M7FVuk+Wj0CIBibNzZ6uq7xI4EzduHkvywQ69uKE9cR7m+qlNNIlmn8TkLR8Jioe
7v0gQOyolWWOXtE69qPQE42dHonmlC0fX0wTgy1Lrub4bmZDbFhpF4DJ72l6buUh
DVdliKiPUk8g3mTGxW/Radq9RhldbzKjvWb2FfsB22fwSw71RpP+08mZOfJGVtFA
OkwdRwxAX/s5DGZWVjFe2Fag8huvIGhHzXapOuq/waIgOuySAYvu8aMYcpXCGLHh
QAlLvu84CRvpT5yDVv6PYRS8X7inFGo+8JO4fL3sUdp2NkhFu4P8SivcUIdeDd2O
sMyyhmjdtGEoPWmRm+4fKT27ljDnTFc0B5mB6klUU+99iKqwAPZJe2HmBHwKsq+5
kic06da/D28vFXuIHfI1OY0PDloMKgAEnlIAvA3fhu02rj43oWJoZ4bVwMJtt1W8
W8A8vUmlH0NYMmhto4osvLalDkbMAaaUtR2IW5cgCu/uKAEohIyDCkVZ9qXGjAi/
DQnv/IYL1WNqGupNn8JXeXIumAuzK+0sjQfcfe7YggIYfILLhpENa1RJVQNVRplF
Nn0DilLIGGsglBycGJ3fTWyoqL2aGrAYIZrLpQue5n474bN5hsj+Mn69FIOZPLHv
TJytViL+Sh/z55BBXU4ohpasLlSYd3DOISQ/5ATFWZE+CvlCvcUKo5EAojXVDD3f
c74oueIgBrQk97IagAgcD1keG3lyohpySaUh9TOogPmxUWh2A85IZwCZLOwDHH27
kddtbHZJNH9M0MZQowXjy3QdA1+WMWY76+HaUzSad9/1+jYCjKCnMPh0BM70X7F6
dgWqH/5BdfNFtXigAvmA4Pbf23jiJMdfH6TAfqYv0//zGRtxLyVRf5BPx1ys8pog
x5Ghg+wAsCaHL1qTqse0waW8cb2jjhO1yUZtv5P4eUPhMhg5lJ00o/yr/NAOZ0x5
eR6rMyyO5wgBs55QmVwbDjQ5YKxX4xpi0nmqTytnRVIOKYWI5cIn2RRwKKNpMe89
E3E08XyXAM5RtMzsq2Za6rIDzAwn7eGHuI1xRDLsCYB4p58W7+3jf/DesUZZhZ6b
h9hbCu2kMcyuroejvob4wte924wFxenE8rUPHCagTkIViVAN10j2bbOL0eL64YgW
oJLWzXflSv7YikPMD1KIkheixo06X95c9gqQEzVmiLDIxfy/v80VhV5vZ6GLviUe
xh/ckD1Rz+V2uMPNgwrNa2oFDoAm6sskCics37ZR481LCAORywF6nR2jyj0rTv7m
ihG3txqjPQvxgZMjWvYzxQTloLaquWiP1KWha9a4EewbFiFP7klJhYiDkijZwZlW
rLXgo+KE/Mrp7JhnMIK9ndudmrreLTY4sS0Nq9WEy70wqGoY9L06l9U9XCZASWNe
wmjkwKMZ/GaxL8per8w8Hx81UKZRMGRXJ9MX0xet4/astoqcW/sB+3tVsAFK2nJy
6y/uqRYPY+ar6H4xhfnedGnzIrmwW4iD2vBliy7Ms2sBRi9N9eXEqUf8F74ZmQpQ
AOkekrXnjrTOQ3vDUrsKesDxEeFJ7UzdbMrDNfIY769atb5nVRRBEyScSPowwg2u
V0EsJhGZ8gPf8MpOBuPmtxmWAuFhuCHB5jGdAn4OkrIlVkqtYmDzy5pf/KxClNgB
4tCnIW+nvEGN6NUITPYgNjP1k6SGRJ+lhEAOqkDPWMdaAsxS7QozirPN2yW1mKy4
lsTKDUJB1pHwSrlFfTj2Qq/6cLrfjXgBupQYlOq+aDyK/RK46zQSKdVRZF8H+Wur
22E2GStD2Ufx0aYV2iYjoP8RDwv7YndWr6HJRE7aZhU6Xv1yelnGhNs5j99/Fj9a
qZlreSmV11nVw6MfiknG378hBhmLjUDAh0AM1KMU6M6cHZzj8pLjyxZ+SQcqkSZB
LZb3BPjARPWCrQyzzP6OJoipfRsLkeYlvtva/cfgOme10Hd8NSKWb94PvalxrBLL
foUFKmUfRYW5hansqflckAT1qCaUmYeo+Q7sb/FO3d30oJx8TBdKG8NhifkhYiDe
OK1VlVqVxMPu6eslNHPb8QgAnJ9wPdUNbzsjzx+xKAQrNeoydhQfhHgaz+Tznuvu
FTp2HoLfsqwJ1z/JxKgiSGNEu6JGEcx04sc4DXRPOs5DiWbd57umHCGojEKQl96V
gUF+ILQ0pJW81qUv6IckI7U0MLCHIRO0qYFUfC1BoePLeivG2hxf15rk89/hOCOg
/Sr1av+j7DgvzlnR6rOg7c21hc8oy38OV+MGJcnerEr/tVz0msTNnX88ZT6g/dah
4rLZnu6mokI2luGeoJsGyyKw8O4JpHTCs5+DCYrSm3cqD7gjHpJNjNun71l1sKqH
lnzgOuukjE9I4/4QjJS7VcTlMQNfxg+80GJ9rwDZtIHLQfEplp3n6MhxcrvSxDPj
QIJKvUyKCcFM6Oot6dss0NWWmjS2Jk6v1xB81ii13pgxtQoEhTyY/clpr3QSJPVG
0l6qIvP1DHpVRu+OqgYmmSzqxpMWR8YljGgYX+UNKyV2wqe+/5LCK18Smx625n3Y
gqcpHzgovseCgVgOuCojriNhSRdBVhY92xVE4SYPBqwhrTPG1wbVNbfU4utY7xwX
bWHBt6r2J6fSj++bXr2Li8WuZ+sk/qY2QH1Do6XLdZXCHuYZQYKXF35+JmoVZOk+
QDnRc+PSpYVMcvRKkZtfaEX2kUvjhIIv8m/RqiYJElBsSBs8ltyCtcO8qLaQm06/
UMPGVlBEa7QUYxcIh6OrDWKyYkCcgFtbNBr5VBGrWgSBDkiADZ9ndf5OqXr06wkt
DoXeSzacoL4bta3YVXLLLcdSVUVqml/lAEq4Gzcsi4EjNTlu0SclnFpbdaGBnpoy
AHiel4GnjgKo1FkKAx1l9jkyEGfaIaXxC8CCv38OEHNJkQC2yTnNvtCa12uJzolH
jRSBPLX7CJnmH2MykbLDlM79wCabifxo2izHzxcGFyIUOmUynPJHizmveVt2UEZg
8ccGHIViTYcPfR+qSW7LJaBRrZoCKmXtZ9/eI13oqZSW9nNM3O79OWjW2XV5a9Vi
UKlikKC9ZmaOkYk0oxcNGk4W+/cKGpI54FaVvsUQJ42QcB0F5o/LtKu3NHKawFJc
jRRa/RpJA0iB0y3UayCe1/1hlAwZwG1hKWMKbFoM8rfXPwXl0IbKeNFl3bKyhVBZ
nckKgoZ0XOW/dCblITqzLOBv/5m6kkblqSqjPW+YLTMWIoQPIB3KIM/aOateIo2U
9xwKXVPlis1yhIEQOrSt1YTLxYmUU04aysK2CKDO6Gl4z4h+3FXi4N7prnhnHKrm
xm81DSLxRS+hKE8PEaUUpNRPqBTAdLyGJRNCuy5OihOKWi7Cq88QMx94vwT8ofpX
KDn0aqhpjL0lXVX3Ad6Syq5LoEPzLahHFxjOUdMeWLk/ixPq33KrVWMcl6FIU5iL
ovWLjRvLpBHEBPO1X/cpxRkXqp4rwQ1SQGJ2JdO8DIy1nV2M+mya9M9FvIWiLVoY
J3rVWNq4TeNN+wqsK7rBl0G/YQjNMpZNl2t8FfxjdMTT5sp6F2f879JWina6wKbs
bLvhaWq8lRLr4JLVn017ubFSsUb4+XVxJujvgOUy68e6N8cVaH/5Q5HWjR8vEzr3
IYA/6+9M5kI0Bdjt+VjJPHF7QeKN5kxWJCp6g3Q/Mzh9GXuipzGetxTNpNU8gLF8
+Twfk/P5uBN7kcyv32vJkd4eO1Z6GchYdCZq8Ros/bofQsULIGJ5fTceQfSm3aVx
NEd8ogmWafwjGSIreTXB1s4ktFF2amDqjE0Bc8Vb7FESJBntKOWm84As70xMgnkW
QxBvAI03fpZfgHYGZovWLSQLEOjM5BH+eSx/hRBzCg1/2/RxOR5XqzNrtQJviKWb
ohtGOVoMEcF4GQ7Y2+BFOZfn52CAQ6E/5DDxRdCAbGXoxRiJLmK3ueMlf1Xoe2A7
1h4/8GTtgNbpiIFhUJWG7TvcwxQg5t+XnFWXDLuTvuH2bg1yA7t7pGzxMIKI3RTV
tXMidsoW7f1mTfehCuyfHm5y1ajT9ewUz7eqvcc7SYa1XF9GoJgrPNJv/7s5MklN
XqPh4XJpcg56QfDVaNBxcq48hdeaTJ3GSUV1YlSyvIPrczqlYyzGevWDfB3cDcva
tDky+gl3qvRGwmzBvI3Y2SFeGkOLiltPDfvNPvo0S1e/FlIhXmqZlDjVqTEPcbHP
NtZ440rm2ns0hAaz9IEZ4c7IOf5XFL0YSUfsocsMpvDXIFNwntOQT2vKX3JG/t75
Doj1AmhvL1ESEX5D9aoSC8CXcV+M0l9GA5AhVcKN2hpu5qNKFBjtSguC1Nw3/JOe
ntiAyEVrO8bQ7Bhz8v6m4RYZ/re6Lv3AmvhhHveQ6LuBZkW1JYrguFthIRhGbNOA
/pDpBhDenECnPKI3iAyfntt/R3UO2+jkgaP7g6OYuTZ+H5xfr5JlrNBADh1teGSu
s7BvgehCX7dyHkOegdLJjeultJKd2NMI4IJbt51Z5YY+4YgPYe9rMudzosPPKht4
OGwF2/F2JMu2XMXvkXxKlWEULEFFsDNqoNPaXQBR6hn1A6GI4+QxZLG1HO8SYQUu
2Hko9l251FAlWkMrUVdizbE349e/3ciLCQfcMgrCXbRxz6MY7K2T7f12v6Z1wqrW
+oUtxXHGhq2Q+FGQGNKsWxw1iRVnYZM7yQ3OA73W2xVvHIqfKH/7TDRONmVceAoS
mdR0+i3S54F29j/wSDbvNKW53OZwuee7ed8q/UqgDegdPdrGWrmiS8JwFkQNCMMr
BN+g42cMMdSiEx63Dc7xB6l0/zrAJWM96qnmljflOFnSjdSnPaZKT/0zhHGCysPM
SeNLv5PEdPAxciZhgtS+KaseVhIa3ZIhKDFqGkobtuz6AIfYpQSTJiPjYxLzBwfL
kBVpa+e3Z3EYMVso1YcyuYnR7X1GFeyRV/lD60bJMwSYcD9xa/WwYFkFoJ8ifiuj
Fy3Eq6XDrlbDuPW97AzqQmyawVkmEb0xbQta7ffv/sJLwLGbrbnklWu964TrF4k9
Kvx505sIp3JmF34UX+JGCQSPjP4unPblWdYsqio09QNa3yniIBv9a//NK7gQFZk/
F0k21mm+f3tY5te9YG8k6c9P8VVODdn1gUksIqQqUAfHLhxHcrimTzyfgbtg0g+N
rflZqgDFXNyIGwBn2HMvmvEU0XQkdslCPilvu1Y+MiKoWABKER9H7koCxZD8N4d5
5Pvqgdkc6Rjx0f94SCsB/ulE7Z/MF3oBhIELMBeHlzUI8GY6kLpZmtCRLzaEnI86
1U8Lu0TowbhRly6jRnUMrUAaWk2zt+FsaWuaWTXySITLaXTbOSuapQFy6KjCuPP4
oeHU+Yuo3cKR7Sw3+Udu2jtjjNFijhLnh0uFdtBG8IijLXKaMqpPupWMEgkTyO17
kAQV+n0nXzdOL8PEKzZ8da5jhvJN/VycLblW9DNBNmWGk0rOiXTOLHcaBwoAwI2w
jb8UGx1pjQniePE5w8gMOxyAEKmtScNl3YLpgoHdo12LBhr9FLnZb7vdbzE6xaiP
3pOPksfHRtqg2XRxOJby2gbzDLZoWL2bw8Jd+iSZWzxkgfLWgsNFAIXPii91MxD4
Cy9Va5nsa4uK6Z5j0mFjwgjIDomRdkIY2BvBCWT6bgD7BEVEUti1piV1v/ojNwJy
CqViuuqAibKuJGYGw8nHPZInKhLqgR9Y1At8J6XseOwmDFyDDw57JjhukPMbW479
nVWpskfGE4H62RQmHp1vqdT58pF5XcTxPFWUIC/mIQtXw/1iBT/oIkTGnEB9mYTC
4hvjSroEnCl7bj3Cqh+yWwzZvYJtRsY48TBX0vQmPQ+zWwwUNHa8QIHxrkIAw4AZ
qdzn++7l9rMegjOhHzF3jTt+qVaso9LPCM3Db+6+md50IajG3jJ6Dxv1t1fRHenT
R7VFcZXHhx87ZFnfN6aX71j4hNRdvLw58XlgOnAkFltW7rsXVMRsgtWihMuGztHQ
eXNHLthq5bO9VddO0/hYyrDsBycdKBzNoE/vK3aH3Me+ocUlHAUDUws724N2XpiQ
t8kfuD6ZmCnnOkTLmDm7QXnXRcfJdZnFUi94k761Ce+8Dsg97sqEhGme5u2YjSM9
TtyAJpmUXAm4glG+3DcEuZYaj4+Mn6YjOewzHHrnG4s6BcoXMwNcv66uv2HlmFK3
31HciQhJXlCH3Hlp39IEChL+wGo5CrYeO5DNoa+3QXRha8M1frHgTqcnLHrsXi7t
t14BrbU26pGwmgRwk3Chgo1xH0cdOc3P1Jy/3xaY9HKB2q08rCKOQhfCe+yhXLHk
Qq0q6WGQFXaXrOpUDezf/QaA2n6cnyu52aKSThLbeNhEsmSn2kbVmE2qw/fwilwP
dqdSjeoVIxTTPh4vTl2MQikQbLD7nfwtvO2yL4ObCxJaTzxgafLOzGajDG40UOpN
/TJ/Z4UbYnp6W6V1x7g5rMVGpOppBX5snDVizf3N39fkR07jUY6yOYdNN2emt6JO
uteqE8HGTvuDaF7Sc1++3Zc74myjpfyo7mDjQR2MrLeqYQo/ijr8Ajjcz7Q77kCh
LIkAwHivhlOPjrh/6L/2E63PMVBidyN086XigT2JerMWU7e6+K5QIX+0TUSFr2EN
hLXehVgk7IsfxrihOjVSTI0gnzA15Jzk4DI3IdPZpR3vC+qPK62wftCRLYQN9fqw
8SgYHrVvvY5/W4Fq2rKyVjjBcnhNtHppqWloAeJteGIQtMXq5V6526ZDxPgp6jL6
sypMuBA3Q1chuCGzca3h5MBQNnrbNAlB2hbCtSN1YFlLj7xXveF8ELANTKLKjzoO
Sd4pAjTP7eYZ6oMUpoYV/Da+8MlpSrKG/ZCTHzbMqcvS3Qbl7vUrsTGWnSZ98yIz
jrRCAZKl4NbA9eUUkGzKd58Ercq9iwZ/lXi3aAxcyBTMhhIhzisBz2JAVpmaBI9k
JIKknHdsmg6fD8PTdEANprI+15Cw7TPzKR9Ct3Emyw0WpVvH5j54a6OraA6DDBFx
1fqN72obT8p4Sc//0/IiGxS/Sv8hJxUqCkU4V1YRoyjZYxKFNacVY43bUVp1eme1
Jj+Yvy6XFpHlu+0+haybAkLBGtD+SlKQ5O68UmOqdeS3Sp5rPOgsdV7iFeks30dt
aSKS6LQyYFmbDgUfvVQ8RaJzIdk92IdgPR83PE6TOqlr0YnDMC34ubEGVrf5l1D+
+8p2phKPjjPzjikW20BcrVZZSGOhsfiByhBbXNN8R8CnnwQlovlbNLBC0ygGJ1v/
FXYkHznyJrbnYV0p5eZNJIZ+47DeRUkCj85RQJOUvJurRrtshvtpch3DkCjZ11c7
+UYTkOKu2Wv6vyPNx4Xvos1CL/FrqFc3xCEzM0+rhfLvLknHafcaYI+PQo361uOX
LDVEKLjg6TmxKqbLDFFvI7UqPy3M7m3imGJ+4ioC3mgthNxHkgpG99ea4/THRPnd
+CVOEjYt5VPrczWEavNHHgoW9BnvRi+xE4hSWHM67WgZEAI6SrH3ohkQYLN4oegi
MmlEf4tTuIez42LEXwHf47xDvN43Rl8LJ2PTuYlF+Vw84uMfVn7vCIgYK/gJXzOn
s12Loej+/TYlBzlKG30FiJPNtVWfez1hv//kdcaq1eE3xxStVeG3D+VtHIFAUaxc
XRefaOaiixEtcqdDR+E56T0oHKqOTNyu71fFb4ObtYY0NzgShjVWYDfxnCOtkZ23
RVqXmIgQDrXfNz7PqsJ64sKR0Zyp2reD8kQhO+x/2cpPwv/Vbp4aOJXBYoUAtMM9

//pragma protect end_data_block
//pragma protect digest_block
8TNXq9hlFO+x+dlyvcUYE4smV4U=
//pragma protect end_digest_block
//pragma protect end_protected
