`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
SXcrpxeLG8i3Yz8F6C1LGM4On396PJeCdC3xe30DkeSFMkvHQ/9Wd1asTL2uWQQa
eCBJKmkryShuVqfU6O+WvhJcsgNTeY9ph2MahQ1S5kXpUmHLtYK4CfKs/wvij+mn
wqRWFu6MtMHschzS96JchhhahydUoVXAcgGNAveneK0=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 8576), data_block
vc3dPIh35sQ9xgI8Y6515XpMWFD6IsWkiPf3olNx/Y6l66nV6n8iJQg03LzIky6A
rLF3JhVVSnjknp9hJTpDjOOTUrrgcXSHlV9U7zijsYh7THGZH9IDDGMY3xXpe7ZZ
W7L/6xrjuSxWB6K0+t5sC8V4V0NyYD8JoWaGOg4A4WGdh+fsq/29OBvO4Il6fFLz
K0KiggdXwBOcaCeRaj9caSTbRC9GzXPm4HOc8jhExT5SsNWHwMTN9tlG7uflwZGq
5FXPRA358Fty+NaxyTqwTeUeyt+aSa54xp4yP4XDgvbvJa6DuQle59HaA1ryGIuj
cVLAnAlcbBUC0c+Ez57mrQ8VccbnGl3U5FA8oHDs0a+LZo9f/fXPmrSEFfQAJZ6q
HzY+QHuXfucbQgqDIvHW6r3LQPE+xYYYCfxMDa9UKtMhzRtPQyb9wIJUMIyTDLY+
3KqSZsAqLmE7WE33uAW8gD3dnOxEARVhqqYyo2eHLnnr3K96R7UokcSv9RK3MGad
YRxtWkfJdng9oEX2kdFb9Z9g9SXdKT/1tK0to8YV4U/qmuL8FyijlF2JyNi8LkYg
wtbMHoOp54pHRTRMWBrfxkozBjBN0V8JWuFWRsQwFEnJjrlCUo8NvNMpoSjZW8GX
lzkF+7u/WTMhMqeGRR6i5p3lDo+QM5D0sPMhFzXNZkNSXk6yHxSf3XGr4fN34lR6
dBzuYO3w9NMaebwJY8LmvGO+1SaKLXhebFSFMdvg5TuaJG47THVXly8eshltngrN
hkaAjFrL42bmGbIeAxazkW6/iaBX3PxThYhOySvL1IIxYyF45OW7B3K+BE1TdzOQ
Rfxk2kWWfuDXQZjnTKOOfRWSAPWkXYSV5CwDNqmxCZAMB7dMeULxXQR64urwv6g/
Nu6ORWsUZQtKqYhMemZUGwtueJRyNjLnigLc50Nf1XGJKxvtKC/FWZDRWakxs7MG
n3/5X6CUy2O/+VS5GMa5O6iZhceXCQOkgOJHeIUE9noih+kBmauT8H46QJoLe+FN
vja/wHCYgT4SgdLjB/YyfPHkfjYK3/80Hjzzz4dPemvI8sgcImUOn9+kqXKoXsht
SQU3NWBKhhuUqolxUlQmkS8DPxomG41CkhigAHegzXmFjVoCBCccb95UaLd2SEeV
6OGhDtOqjQa8AOETlNPwMu0e9zR92ZX51M5agTPHBI/7O6vvH53P9HS717SCAlWX
4dzqVvrseqtli5kF/ZYBfGTf2EBt8eCdriwcDmDiLNOV0aYgzklrUyFBqE7zkeNL
rb8fw/DV3T88yWuGGAWKXbcFpurjtx6Jb+o6DkHcvjxX322A5/qhHRg26IUd0bT5
TjSlcgkawB6p4ulXSL/uTigcwZ1vBXRa6muXHHvF50YyLO8qbRMtSonYkp0EE75k
0bjwOdVISpsQ/CrA2a82UH2NnZcBrPevVDQb/oqzJDhPiZstbODwJ+qH2hVfKVEI
9kpD6tyjiWu1bi61IE38fK34lG5Tl+ANm39ezY9Hzzw14n3YYjYWeY1kJZzS9xoW
ZuyLGDfYK0+h642xPkZsDg1fyy4WK1pYgU47V6I38TggCleIwme/9DORYVKUxJOb
kEsTSqpNnv867+EO+C51i/6YJQ9vqrCMlEMow061i1Qdyy7U5wGU4tMRCN6E1n/j
Bx1ol+kPFuCoCgPv7NdlXwSWZ5pLTWnwKyF/EVTw9wg9q1BHp5IMoLCOnqqXV3J1
vJ9Hl1d0WFQOwL6a4+PTkfCg8lQV9wEjOQR6aAEnuOb9+SZJJNzgNFUfNsU6KSQm
UDGQJbWfXfIVY83XwsBzu0HtnwDZaDtD+qHKe4/NxinscuPUuVQ7bgeJM2xYdavv
CPTG16CXV74jRYo+6YSdAe5xh/wCKHyp7bJeOWUBVULCjaK7TGA3BWRugMftDYWP
WQlboksFsS16Wfkp2mgImZfFxpXdeW10AgCXAPtzeHwu8Z2CpfoRJgowu6UvIguq
/nTKqvCcGAo4J+/r8mWUKKPOamDLIW3PIBzt1sw70ytWKWSmipEiG9vhfX4cViXl
+4eN0LZkjCeIWHd9TdlzUTTFbOrTF0Bl1/qMDqqtYbBnr/GjLPuxAz91owfiR1Lk
tcEWKv7OdKEOBXOa9NxAxNQgTVTbbitcC0HrbK0ZQyfM1eOCYe4phsXGtU5BbJrJ
3+oY1+vIaUWwT5W0TWJHiaYh0KIuGXMN7g+KYRz8qna0voMLhNTwDmuDP6XWQARy
yTsI5MxxPG4FLU2LK6eUuGlBojXkPny7g0dtouxyw0DoMdxUSo3emaOzfdzloac6
nqf/msDJy/g9vVBPiobGU/9LRbnCeCLnSymCbsMb21d8vsDgEJ5nD4PgmjHdB3+5
Is+z2gIdC5Dxba8KgARRBDTQvFPRVkFzwdWAVHbC9UGU/kS2uHGHW+VEmQC0SvA9
y9lF3Nsx04lH7AU1XheUqDhjBwCqd4ttNjUWft7Q9yE8ebVOSm6wuebvgN3SHrNn
Z9mGg2NX1E3jgQuVCBkHTd6pTbBwSbMsjDEmq7ey0IG2K0IVIiP0CNWEVePqi/UN
tHPMXxbwv1iFT54nIjKty6GzhGy8NMBGDzjSul9q5xcL1rnLR/AhtLKOvrovz43p
mqLaI3nt9XhzaoCYxUwJveCI36ezgNiLztmFfW9bF4/88z3QWwKYsDda8Ag1kg/X
c4DSm8RVk0fYEOXxt8BqtpyrKQOkiHoby7JdvYB9XHD8n6MMcpRxJiSd+vebngO2
Vj6g89008N1wL8VrO2EboRT+AB1k1pmsbMNoJkw0eXQWEULrXeJn/tketQgMV3j2
q08iOVNZvASAqjj/GN0qApSrqPV2QkqMKhxZpj3jgqOz7BXLGga6nkZn8HRUXRmZ
oxcGiP2QRnjW9fKMtjG4VwBtJW9cMuDIB/PWTwZG9gY8aqr65y4DxGFdtPquZtB8
H5yJMUXDWCG3z3CYdKg+p3WFjT51cwrD+pvJDqq2mx+W7/VOP964dfVXC7Kz+SrZ
Tbmqx1gb+2AOis6wChH5WLK6sK5QpIfR8g7X19cls7TDs7bBxlNpjcKOqC6fzOYW
xphCifPsMphy7DVe3qzXLwJHcRmR70BXB3DV5iSKv89aVNJfnYFxtJ77bIhcsvBl
uSx069MzzWFuYPX8N5n4Tt4ZiJg5Bp9Rl7Ova+y60dxgZtCyEh5bA2D7Rzaam+y4
PBNedwAMqbXD6ZuYg10QFmRom7YI8CRCj3CocDPM7JNyzrLWwS/+ouXmGrzwKh33
hId0qbdqqYJhHDbQzmvzKnQhK1gEuN3u4vC7ijs0DZWMJNACH/G/hL1viE3rfcxQ
o95GkjMNkJ/xiLliWtAsOX/12t3u8DJkuRgttybRSbFy5gHRmxbkUXg9IBc/hBoj
81Gvkkw8nLH5ZWq1rTXVam/CkPwXjW6YeqSXwdA6NKpRw8am1brRIzvd5XXMMggP
7/mFU5kmDhlnyysFBzJ/8s2VM49AHLdDWz6XPiS2QLInh66Y32OHdqLqRhPHwuMe
X/x3jkzslzIn6O1hf8CMD4Ljba/RM3j4h6v0szlP2ApfeiqlmpjGhsX8AFEMT6RJ
kMJLE74ri4DWznUFZdwETeSfdo1L2WRj6YEQ59IXvmNAfxOlt2Bqfpkb3o7QDYtU
Kfzn9BBFF6xtF650r0UPthAxB8mZoNMAal2+oBxci1xCYysNOD3NkFNHV+9+d3lD
Hqm8Lw5XKuT/ORr5jNVOYPgfRd6zwaFh81Y1wSDtQDF9BK+f49rZyRdWSxAbe+ro
FDUTO7Ki7obk+0/rW8zvCpqTMu/Wlq54IbA6C0zucHzLxNfGL1f68dFl21fg6PH9
c5t/oHSOrWqwSv6vq+uHTuscQ5EafGc/kCbXwjJAiozrpBkXE58V1Ptg6FfWJLNb
3lmr8iodXY+eMASSYECuumYQ4nyM9k56ilIYGtvTdlEGCOymslfge5wxtJkNamnq
GvRvu0cchVXS00VYIJqQpmfWAIie0oJ1rHgR5LWyaYZrAouo20HRHBCr85HpIQXX
dzApTgHNy+xZdRI38DUhw6qw6OAj496ds6Mzk46FymlvdfLapP04ha2Rtdi+AuQj
+HHMe6s9wCan/qL1bbldvwIpzBLYdzBa3cHoZsYYKpwGj6Djy6+lH+GTSGJYvRwy
yqEHHZkXwOCgN0rfawERAUPKjEXckO4cuwjg9mPbDx8X9RRF3s+Xu05E2tAut84a
J2eTpaRa6AA/H2NLwpFLZVvMgXir5/jnllVe7nMj9H8DsVH3mXrcl2uUbnP75X8C
QE0pHZX29AfidhPl5EromuewKvpwnBeR5728/YEfhaXsECk0xP+W53FmbHAUW/P6
0+HX5/5U3Xu7tCWR3pv3wYKyCrzZVQjOClXmKYuMgw+CfNEfxGGm78b9eMAvTVai
Fy1YBd5U8uXhmF5r0xA0E5cGyhNmFQsk+CF/Dh5BmCfJXitrfn9nCbAWdGqD/QQQ
RV4qdpOgr/q0aTn3mCrQNlHckSTSUzAtIZj26FzMOfnYrcBiiUEucHKoLnrGU0sk
6a8YE0E+RQClFLEL17NjDC4jiHx70aF2KpUsvsXgcnKLsGdTHVF9TUfIjEl3mGds
Ah5BoFw5Y6TS2YCCJ1hDoswKabW/WRdOp3rgg+Ws8TfOi+tc8h3DoK/frPa8viXe
uiCGQfHHpeB5Kek/V9ne6t1VW7IZoW/U9J6D70shvlDY+OpF/vZc1Dy81iKrZXTv
BNTFoswogAkshQvofcj9G7oXfUScen+LbtL/u8Z/9VgYvKVimR+3vY3wLg+adOFi
UsO1NykXQFqqqRdS+/CFTY2WsVPjV+HnKMxq5xVXnbxBe2B3eDae1GUIkHCEK71m
+ZRBjQdikkMTBEKrw3g6hsjp/vPJLl5UtbSfDlfL+91eO6DrLiT4pLjl+nm+N2yM
m+Zskzt9n9TWVOBIiZJHa3GMmFvbSSIzAzggQWJk/tfdu9uvvBPE5wFlelpBoWFj
72nFUUDzwTpchdSOM+4JZXLZggj8qUwWFiaW63Bn9x8sbG5muu+w968RaGtXynv1
AklXYJOAWgN8y7Au79hCybU9hE0BNqR+t7HRtEXfnf7MfN/976Le9pw2FbWuXsuW
XpivUjD+8+sqK2C1v5dxSzGQaUsnpcYvNwDnAJ6niI5eqPk7fFbY4XCqrTKOOph7
8iM/LYBKFSxdBahAJGeYHv4TEhR/uyWWMoxRUlhk5mjgebuYg8wyG2bRpcIZheUL
VMpYTkrQKp2Bg9r9rv5WDwliSuHDroBNB0IB6A+G/LIEXpzvvGqArHkloGCudG8b
Hh3qzXmINo1+jaLwD1JDdMih8tqS83UKmEUvRbSg/x9T051PC9X+STpQkfHKJ+C1
ZQU14vtzzWwm8QPOv8dokHJEjvd83/3aIUYMWb6no2Fyom1LYDF3AFbZqF6KNRs5
hPLEtHwLGIkCpvtwHhG+JPGKm9hZEBB9UBqZnXYVIiajkvaLQuE+e8YcaBXyrzYk
lKO33lQbXCSmAUajJZcfXbtSdq0Ztti74rZp3qoHYyDYB+XSjAOTUtbKd2xCFe5L
T3jlnNP4x+e8tYYx8uNNXDsHLOGVOGcuRA8mjXE/xVH2itdzvNy/YTbUqM2nwK/y
FGAZNVQo34XoTIO01p4ZDTWU139AGVvpwFRp8qQiCz1bqNtjfSklBhet6LVZJmrz
+7vGva7SoTS6gShTVKu/M9tzDKpiJf0QpUaM/uJGqmEopJO0uwR/0EyJj00dVu6k
cBh8GIj8KTvZ/Mp2s8JpyzvN/gdljkdLcxC5+PiP1jydVlNYOmrONvFv7VRqYtV1
JKGUkVVKjEWrhLtpThkX00XyGjhXBHeppUrOeyQcRR6wds83NlJQVPdm/az0mhp5
fQwFh9APp22R8dLY3d7H3HjyVEWbC5sJ06QTkE88uYrpLlyfeizDvuZbxX44+Hfx
ojMmlFdsHvOX9FHGPmcpixsw9ZTwld2Qi/aogCOuZvAwKnSzjeRdFGz+YF34k8k2
3gITe3xH1Qp6PTlqrmNBbNe0iKvQR9yqNKgQh5kbG6oiF6lYjCVp/hY3sAwc56kO
OMuJBv/yUnHFjcYmTCVtW6UP8ZaQgVt1F5Ra3Cpai9hpGMlRVFBGgP5XTo7n/6/R
yjaoeJtzJ7q+BSBBdftrGJKRhtUnp+B+vHr7a6ncKFPl730LjZEsSfhbeDiVeX8w
WNh1qqSoDYOJ9cj/0V2A5ujE4m5CUWLMU60na+4fU/AAilHfCq+yAX1ZmUhvCOMU
vdQjLg5wd3wXRJjufltfzwB6qKWqTugE0zsukW78WXqwOXs9dIoHWMmIWl3le2FG
9hh5j+AFUXcDO6whlN6ObNooXNDk4bWX9UAXFgNFl60wh/HSCjk9USy4NBAb9hMj
wPso5u8uy/9jYEbW2jtzmm92yv7LF99WtJJuv9zID2lp8tJq3HcYncKZEfO8z1vy
jt5Qj2Qhv/M93wYMQ+bKrVVYvY6ChCVvDrLa8O2y5ZUTq5TmcdIoZo5UGo46V7ZY
M3AenID9ue8iAQGNsKcOrPAL8Nbi++FtjvFGB7Hpo3xi1zwyspWlspuJ3o54utHC
x1lPDhnyszHvA5YUHPQKsjwH/Wvuvi+lZO0DgBTaznH2tsF7U0WlbsbVlfhMTS+x
4LYIM3FWgmLrRlloOl7KLs74xnEuX1FdwCzGl+F46SXXQgKff0N2ja0XOWByVcCP
dJ8tfM2upLdtze66C7i/A+t0bFqYZqPN8axmZQvMgK/IsL7KA5lRoDuYg4yFIolj
XzC0KLy2ZoICU2EIUeyg+eFjOfo75rjXqxXiXlNjpMtLTRw0ME+FBAo48uh7p/Hw
V0zKH43msAm0ncam/IhpBRqeBCewXcnSyiyGDtWWUO5b4WUP6LkXOBHpwnJOY41c
L1DpJ5LuVtH+x5eHPAl+a3VvmnSeDAqm5dlksqBrKzS3t7Zu4Us27zgCO6+eBCtV
f0KrfgioPrzWKg9ePN5PbEiStzobLmYd0aNgNj0vP/K+5F1olHNN8//jdD8BE7Qd
BiW7+3mEFYp/0Hdc+gaW7nunhz1sStFiLapdWp3kQ0OUTVVEIvmGTxk6h696Nu8o
Dzh3B0HMcZXbuJyrM+x+UNAfaLoNG7nSeycZsH8u+QCbRu88KtPRA3CUCZC5Un5Z
UzHO+GzUKnUT7Wuup2i7N6zM2WucprLVs/207w4iOuTbZQ7Rn/ZEraMVcrVyd0UT
UwguKCmN9TncouWozM2eJ2la3kuTyV1+ceCNAb+lCOVJXXaJwb+cJcRA4w95Qbq4
trR2e6y/2/RMgmO6WrYOHfck3YibOQmMXwIgevz9mOyS/YPVoHQOgxbF5gs0SK6U
bLzJGaZezMYsD4eKjxXPsBXJ7U6Gf4gdCOqsOs88xa3RMY2BKHH0TYuObP0JFtam
3Ii/ii7ZAMfWtXJoeGIS0HgzOBtG8FX4FJyQbf1ovlDOWqYKcyiK9ZdDBhhlXxln
6j9+6rYUzGmlxD/MnlPSoCT2iHNe1picuc0yhAfwKEgga8O3TKrLaOD/2dW8C6IZ
ehWUhOpwSvDY4buIv4IioAWNAXhpea/4W3g9xM5c79CvXpAsp085HKC0JCvORdyM
Yp4KlTsThwiw0nXbwnGf/Ao5OorzbDsdvYCpGIAD8IxQPvq9yRzBhBGDhpcA0bZ0
G6Fbiw0nDM9VLnYQ+MKT9feL0okI3FvS238WzGMm0MCzynW2gU4Bum20mslxKybu
LUnlz4brZfz9BPd6sxuhhY8vaMDL9+pthxTyW+KRsbqGHSVu9zgtZhOpAXkiuzEt
9V9ekRoM5v9EbzhgvXc04rUX71T+jkUwHiZC/LPb4d6Z7Lk0nPB5FskwiFm8oj08
ZUvB29+EBEd3X1iMSvC6nLtdNI2ujhgC8pOJ/cM9V/96oOFfQ78CpqWt0IULFlr0
OHZIjc7ODajUWuZGe9823X7JyoJAmWs5PD3x/RT6Y00TG8T2Jj854JpT3Ko5z7n5
4BVgn/7oaf67XJQNBBfdvaMpSCln9v3dbujrhAcCijk9a8LGc9/OJmrQYvg4AbUE
Zrd5wgsWkNw9g/W+DqbZMY9fBwpdjq28edrHAuYCQ8U33CG/A1npAedS2X5rMpXq
2pLF1lCDPIsv7X2nRAn73j78YO0EPRdt1Da2YBhS36n6Bt7tquWtjcDFwNwA+4rc
1qPm7HWQ4EeL5+ZW7tTBoNxZxGjSFwUlZDjMkbIUfp23J6Q3qfO/ricYUZ2EVMH3
OZVaNFeqbI56IJUfGIUCltXk6UnNL5w9umDe1sHyEJCH3fORjWwm8T9BzzV6q0zt
tpX9Pntpn4XmU8h80MrD7R5YIvCL1e3fM9gqHhq368NOSZHRJ9KJA9figpUatDbN
wY6aXSrBviO4w7uhqeaz8TjbzwpK2JMzE4MT9hTaXoz03dd2AKDPk9BCojqrZU7P
iGvZox10OvqqIzoMMOCnGcyngX5qQhBBo4yLwZiGKtqg03HYDZVPEdMEZKod3ZkQ
4pPPYN6DpeNYyOy4rv7Q5VmZQjPeqps7aHvwJwXOH+79yg6jCaLyeF1SvDO5CX70
9teGfJUn4J6vxgvbhI/xtNWa88AcCAQEORox+YBcxAxy7A1y9KAu22i/PcsWmB5d
EB0ENz0LHtYksXjbDBLUYcVkAl32rw9YFTywkoww/Y9dzcsNPB0Kpjg2U/jpfUT+
Cz4dGcYJUWVzILfIKZm3KEjeD718KxPgzvIl+STWJMEiwixiJ3uqdTLzDPEpq94n
MRwLEWru5D58cDfW5+0aJFcqcb2C9KzZizv3UAnfU4Tyq/xkUlfcoC5IkfQqu0l/
HY0tH+PD+3oP/lwlTSMGn7AkmSxy09wKgS3q3dzan3a4PK56HeHb9Nxa2iaytlLl
AGjvm/7QYMGNtX2Ty+4Rh48gVNodEPM52SBwUUzUV+NZJ3Ppwap8vQ0R/EySSmlW
7PqAeo13jqVUet7BdNYp3iJQmZteLHRaPzwtvyNtgxf/qBEjvk/BPa+yDuo473wH
2J4w0IkXsZ0uDU1EG1KgguA749T3ACQsSy+pJiTpUySrV5K4FdidnvwXH3tOJrh0
5BPpGBE/hW3mlmEFznspkMwprvGRnXqksVnGeKZo9PY+cQ+PK6+/mdNb6zrkGWKO
7HJdKF69PmL5PlQOx0peiX8VIDCivlUB7+84ZdMcNq3BxWWr9XojmWdFEaYGBFYl
m/NXaQUJ/koTo7wWqa6wCnqBWHmFJOlbEFdz19QDBZMwMB82VZdGi1EtX+THNhy/
DZzF5Ciivg0n63ibMrayqFVrShz59nEVMGcLbDW71BunCsDXNVY/5rIMcFITtVO7
tHHRFdbG6OZFVd4Fs0+cnGO14WJY+jdhp2fhR7BV/heYESoQA6yjgJ3VKuIrbbKs
ZvnMci0LMxeZL12OGIYNfukaaFT5r9v/p6k0IdSn2ibtzfNq0vVo0HlyIeGe6L7h
PIr0c8Nk107EsGLrc3adOM/fjb09zuRJrbG37wVRt0Dzz/1gCyjYY7refbsHuvyU
eVCKSDSRm7oYOLGdCQ9DEeh/c8AYdvmBiAyaeLLx8ZJr9wj9PbPtTjVSRvgGvcmo
7e3ZCPXg9CPndapkTbK1g3MMEYX8Mf8b5s1Mzz97Yiwm/sQWHs2BdDSbe9qMKX+y
5z8NF3YN2VvQ3FP3AuiAh7euU+VFoZVLvgtPpNZLo6/cyJkcbtvzjaR3c/5scytR
pBFSS+mKnzMVmaT7EDg4ZBj39Jy7T6KEeT2XySBghC+ZvW5qmFsrBJQEsNpwwwir
7edvms3SMMbwPK5ScAzpucdqNaVw1G9Od6rB3IFhWBOQVS+RqIwxjASvmKqXcxaz
ISFBq/pPnAGFjvJQvPUz+Z7Mj0Q7dkMI1gttfdd0OZBZsnRkhCYXCZzH0T0DMqt2
hfbuGe5JqxN2LzC9ZUlyM9q7OVMK0SbI+2r8MYErphbyalqfjK8Uk/Ie0lD+1HfE
trI0j65dypXSn3DwcMEAmtlhjrvBWSazp2Iixg7Rva7PGehEIBN9bc8mn6WN2/r6
V41iw7VPPpYqZ9yU3IMeQ2MpJ2pCe6BGA5QCxSGeXJiPEAfUjDSKrOqxUMjwLUkH
RBBmjH27MPL7bzEnUFa9+J7UH1dVgWenQxUbMCKsE57EcXcohUDBOAJi9t4OoL39
ThIYNxjWoMDEE+ZYSbZfTOJkpQOcwqqKbKTUIS0eDwNguKS4qHH12nXpcn541IU4
gZgwUFnACdrH5snOKReVfIe7bMHz8xpr2DZPG1kgRQA2bC/JgoGDy85k5iWZpf1E
YsApHr+gA2dkCaPHnZWkWCbpDGsZASc+NdfCfkKtx06MNuAm4T8hzFllOmFMSmfb
eiePA4pgGYBG9adIrtjTfN3RnCue0CKu+g4VcnlfdQ74WGBoJOO72wBznXFDJsOu
jzxbbHtfpEl2IyhZQDVWsjOpNo7mbyHCWDm8Q0JTgsHQ9mNAbOSoNHCpLfL2gjkg
FEnUBdPxdWEXoA78za90AQOQZc+It0xpZ6lR/ayHpsxvx0OH3J3xjlO6OwjBx8mM
GRimW/QCo5Be9+0StbCC2pZKxCpUCykxB14DXTsabzTrL+AAAtFUOVpD/0L+L1lN
JcgGOU52dmJblrlcaxGFo0C2rHOUvMh59EOF1WKU/uEq3RjLD/3Wf1lVIOu54G8K
bCgmynbTxUBgUhD7JIkqM40C95eYOS80vLkDVEVc7z8pJkB94/6fx32y/DlEyOKp
IwZ+yQfoij/KgDSFgafA1h7AI8Y75px4LMTpLKhML8LAav91G/WRNtc74glCt8+L
qZzb9rosJUZloq1xtpqcGKi3x4DQ/sJ9NrqD4dBtXqUYZS0Mhc9gma4tstpyZPPh
WE/o4TlQBuXKGqOw2pFrRKCwRK2a53f0YD5tnP+fIHF2EdQ+tcpITDWMHNeiBgv2
L3t9l7xLMR4Ife79ELpRllURV0i2dyQ8yJ09OD3ERhNcwAwvALmGYotFrIPsAxPm
qnJDxyP4k1qD+LAWTiNl6qISa65WhiwWMjsxNnLxryEYvQ2CHhe47JcLiNJ8vLpD
XuRK+8ZFrmPpUt2fUPzzcGn2n0cZBUvoK0sPNgjiIUl8c9eVN60izsSZPIN3g8i1
4v2XGJNB9aEpeziBC/JHSHRPrBB5/NvbZVrJpEUZ3oCXPvYQRZaaVFQAXkHl8NrL
uXNf47fQgrTP29npu3wUFDOm1FhDI+pDb0PdNmJoi71MeYPXiM1w3tyjuXzOwTnO
K9YLvYQX01gTE5BN1+IThse0N0XR4JxdwvZ/ir1+SP6WD5SO4D3URUVay1IXjPIl
Z/JEl/vrA31Tjar7loX6QlKJiWu6nsFpNmF7HOmCbt+SjNkMC5owuslqAJtoHT2M
xIE6m9GRKo93SLnrYaGnzOMEVgScPaQoTY+F1EdWumU=
`pragma protect end_protected
