`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
M8zUiH10lM/GdqZXj3FRLcfxROc1lMe8p216V/lBPjqg/agCHU9fMUcI/uteogXA
iEKf+WCZuSebDL0Z0whYEOWsGjFdfDn2GUP8gTOMNiL8zku+qUm0VRxFZF8JLjCK
EmH4UaIT6tzclqmpuXdy5KTpaRPpZ4M6UCOWoKzBSug=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 8576), data_block
edgv8LRropfQpPxvsEipQqq/LMAPrpyNOUklIf77BK39MPJUVKnHIoyScQdUaLSX
c+H15a3yISE5fleTCZUCnEGfGOe3IelsXI6pbxYsrS2gsgMmqCqT39yoj+Y6E5oa
vF5+eqZNqqzRnblFc1yLZ/n2Rkqk6K9CzGkCVVjVckd3XdCek0VgDbstu0k6wZ4x
XkbQRPZ3pnUgtdCHzAgT4HUeA6RRJvGBZ0rzC6ZOK95lmcOqytyo2klD3P+VPSlp
c2PWb09sUjm6eCMquJHSbTu+TbUlSNT4wacrQbbCld4IqsgW/A125srBcJPUiELz
SDv3wlg6w7ESLIUIlZGyrnBjuAZQxV3s2oQb/L1ZbIIbJrJua3pwD44/sj3PPPea
QM7xgMyQUwywnJhLPvofxIp4FAnKwNx4S7EZzXpPWXIvLAIsIM28trmnPw3d+FdF
+PQtr53DrCGhfenemHKGeu5s0SOYvIo56OoRbPft3synxKyBYydR89HqddILCu2A
ltgNV3liwvmsirEY+lfp45yHEbvrajqOHh5cEPaLFNCg9Iyvzt9mrv0BQaea6aCU
Rt53dGGZrXxvGmlUA377wLidOmJeM0HiRNbnyyczqmJLwHecg4EYYTFRHqgcxecB
xAgkAtncsF9sF4ZpgNcoweGpwxqJ7fIjfbbuoIrq1qi7yuHLXQ2tN2AmKabFkSd2
wWcPCIkvkbymsnLWim93SJt/f8J3ISHYJNHUY9N8mlM55IOBDFFB+tfpkrBo4mt4
kTYzuWdEvYIbz8Jy8RP7wYMX6t4eHRjmKbH7MUMWQop2XafFiLMqU3OgXAmUHNdN
PY2lwk+nekgYfvwtXjlhBrCkGjl4jQBAhy1VDw7CGMK58nEvBSKxbP1jNUcPoryq
BWQeON1ibL+A9fDpTbj8NZUI3smFF6qWzG9k7/8w69Us7HLKdo9N6saqziqiLZS5
PJilzQNfZc+ip9V0rWIfzRuzits3ipgBqq+21diswwd6dE/75g8WCwxjqMMaz6GX
IbaKGGg/gCEdLM84MZ4J24OkD9bVhXpFWE8x8CwhbMN9mLfbgJGIpEIb+CxUbbwA
nepJE11BXbyjqmPO5bqbLalDz9T0yofY7Z0A/ACYsfXbRGGGrfKuIsmZ+gUfEP4B
W0ncquHxw+54xi8LVTcak9WX3rxDWW+yDufUP8YqZZMjsoYpOJBvNdqEicsMS75Q
n0rlRbk0U+rn6F5vHqMWxGfRJ99fYEkiG9wdJy4tUQ8yIWBS+CJzTyc8bOObFux5
YauFh+9A3dwaunr2fwoThLWjIPRy++frFf5k859S5tScCHYwLaNhW422VVyEyNux
PG2UA9wJGsGXSuYwcM04QLSSi9I1nKeQ3euZfk2V/kGnw48yBKIQppkfxwmThg4g
zj0TIqzj7qWCnHYilz/+ohm/aC19zgANNq1nhxIIhDYS685s/oNaMiI87QuMz6DY
RnhLHsjrAWFinotzdJoGiuZbJGqroAMpmQN0bNe+l3ElXXn8YhGgdnXaxW1oDtsW
lAMmy9H7XGC98dzdJCnlRUfcjii3/2Tv0ZxbhkZg1BPV3HMSsek/Se+zlP/9VSJY
76jezofDinMT5TgJ65qityLmCBzDofTTskhd6Mq46o750kbmNrEKxsOJgWoYS6En
oADKOP1VFayOfeG0qE9g+yUJaedNUoTRsQR97Sqy9tSBwGnP0R0k2WBjHPgC0agp
pSJABIPWOEdj/KMLLPjZdcbaryJvAgfGk+fIg4M8yCmyTNOIfCZcoit7wtMywQz6
A4Ykl263VqjPCc4NSwtgEydqazHM25rQoyHDaKtF8AmiSTxxxosJdnFtP2o/8KRA
w4WgieKK+qUFtfJ8PqDukHYDeDHDxnXp3MG+czlHzxEI4s1+VUwld2V1AvJui1gQ
sJcDMd6CeLyBCWMTVlx+B7jqolpTyPAuxJGN5KrMPMHs5qtSFlCDt7Mzt7WDUZm2
TK35RTLoJFLZ772YMKUnntTPsgSQA9qD2pHbx4N9/vi1cDBkNsdpSMmT3NJm10pZ
DdukOD5YCOCqPFdQ1XVouKEDLCsOIW9SBMEhKExgnyDUInkOaybFjzzLsmXfrEuK
U/p903zAMK+2qMMNH9SzZxMuXCX6i9A5eZxMAxmJLtmz+b3ZzZ17oN8IPH5YcoFn
UyebFLVZgjXCIiWeAgOaMlyoZ6mocfUJil+gw1u9/cQgZf30K+wqFuiyo1esujUz
T437aLgjnhWcE3vsYhq29qHqPM2Kp7uv+m1F7eOiaCNAMSU1HOu80+40NrPax79j
AyD7Bi2HNmBLrXsWTy13aWRDYFjFgQqXFYV8kjJjUlz4f+JYp+8J2A0ulZzemNuH
T3ALwe3WMpfRxBBRXfjhoTEx2ECP5jG/w5zyhlCplwbIKZDxiIUZveKAjnVXrQTt
5kr520ck6AjoqOvAxQu0+pJTqRM+dyou0XRfcFZ9JwtIExoUPUcAlHy8GqZl9ot+
dQVYleLx8otDzG5Tyo2S+WQrNptbhvfd2jhw45A+5Rr3V7eLwF2n5D7ja0uRKgmA
xsXWmKtwqpfjyPStVscddWllHohJxaqKo05YPNQxhWG7vWjMTWQ9YGFl04JST8UN
CPuWH+Uh7J1IQgiy/ZrMBpmls6ZwmARamvx04mbn0K+OmxQcicpzEWydEzJDcau6
1FEYj7gvqATK1csjQFmM0VgVPd5hqtvQNAmLzr52YNTy6a3h1mryqIT0id6PpWqn
/dWXxZ3Cp7UfWMdc6xOrBo7SVMSdDWcX3OdazrHpKJ4lcdC3NmttTi5SZiqgSvM0
EdrS06k6/tEKvLg0hdSuZ2rhHKo4zv5FnEsnSkO0iXR9mxEFLTUce5VDbjpUVkNm
hiBWWc7VPWdsB+jnx0hQ4F6lrrTTI+5GO/4TzEz1wsoCFYtEVAW7dseq0/j6dShH
PMkJUgZJxlwnhsdvdg5d9ZJcXXNSI7liJVCe+iP2W8cFmvIG1esYb/l5QxOtahKY
ccxo/yDjxyWa7doteqqywEJhp3CRRYhDviAut3CKsdMIe1XPglHKMKRGDMb9G1ZA
oZWFyQSw78FtTf7g+jFcfb80MwTTr4kWVjxmje8Ssiq4W+tE4qZMD0+kcET+FMBx
t9wD11IUiylrodRm7GLSJCLK337kAoEPcb/8p5QQBrQCxeoXIDTnXmPrSKLMOwLN
t/rVPNW0X6DPcjIcT/n9Vrk5pM9FNvFsBvFjCN7O/Fz02Y8jv/Xjq1SAsGm4RdG7
AnrGp3sm67yx0NKc1bwvbtb8qCUuK57lgdG2AYcQVmZpdgEOJaqfVGZxrmKRNUvB
rnrdrOvZN544MuQR9ccNiWcIetGx0Kp73hDuCml7wfID+LgJsjRY5uANQ4a43k0F
nB6ZfPgne2ddLhtm/SLpiQj922WfoSOJ0VJw5EYK574IUo9vOB58ZSaG29s8JB/G
eK708s5czNY3iwMo0rMk3XPNvDzw/eTHPiM4kkHnCibzevTBBNPUQYsh2JZZ8ayB
t69HxhsX0ke2F4+w35BAVZbsV1rBxS15e2KvtjLLDMbZK0sXxKzjAXskoREcXIgp
hcAl1uMIhs7+mfcdzjekrtcyIn+B9EOAFDt/TQpoea/2WA0JLiuh7J638dNzgTqV
pHRV6maF5aDyDqAqnr62ZAJ7ujg2AdcrxBgszKXi/OtgXwpNOPmLPyjkRZtpQKlH
vQXLyuhDdyiaAXbt/0c2ogNSFn5NX45JO4rlfmZ2EB4eXipVm/SIGgVgprrIzyMs
v19l90hE9bxr7EjQCmcKyQe+p6vHfu7BUYVsfvAyusbQCRm//ZZE6NrORAtYqLNt
AuH4xttEqssmqIUvqbSyA9QLjHFGXY/LW+iBu99+LLqZHREnhA8stECnBr5tpVQk
uFOF1vpIgfnzRiR1EL7CvHyA5SVzkFqyAaWeb/LH5lVtAegb6I4lv9WO+h6pBUUB
Dj/CTBzK1Ygc9DKEfRQLhfPGQ2cGN+eObDIbxSMTdbkiOu6alS1mhRYCcOOU5IYL
WigX3NHH/2Lcgipf59PiLcuuHX6lAE7yapn2DCCnpiiZP122mh6V6f2IMq9ZEAol
ZbNvnnCc4XlcBr/srMrvdcgCfKPqDFbSQfvN0qysHG5mM3hl5nCPymzZA9gzgmBp
2mB0XVeq5E63RxDA70x5V+A4b2sqGNCxBsy7l53uJZsAUK+e7aO7epBvCyTS+m4h
JiKatLUQr7a+Xi8KA7RACIOGN6BoLNQoX/jtNl4q0A8ftkQdzsmP5jESumIgvGpt
DxsXjl8AuLzRzhXiGRJ0F9mL4JvKvAogTMTBms4TIinEcQER0bsohUMRoDLFka3D
dbYW1YqbF4rDGsOKa6yEeKWVn0I0p98Qy9jg/0mhRbfIoI4WjgR9dFsXJpKIA/hB
pkpCbPEx2HKEW2YvxK88KpoLzPWP7hhjZgpvZjHXydcnUu2Ai+u05gcuAC88QW0z
xglCNyJt5cCGmpCAKD22ihBHgEZ4r4xLDgW4NeKGHQ2rpsmjROE2N1QSBEEbO4fL
LqZzaqV9ih0puJDz6UIZbDxlmViTofVzYnGp833ThrvYAUfBJFmD3Wco7wdcfuDs
sFP8N0kc0i3z1mG+WSbNErMJ1PcLhPG0gO72DQlaFkSOYP73fVJPRDnaDSRa9M5I
udNxW9DNLv/QsKXKeDnOezfgGL/KFcFV2tpHkiheI1m2OKl8zr8QttzK8OUBFlZw
Yji3cDV+zUTvDlI51r9xQPky+8rBG53jwhdLpqaUJipLpwT6jAgkgSajo70ny4Os
IlGqILNYuv9OCk/72HxWWDykcYW0zbfEeT7RiUQRz1BGL5/KfaPTqWwXTGCtTDIn
I4ru8oO+9flfZ0EO5EwKxKev53OLsziU6QaLTscwO8AFy5pJMnBwS9oRz6JXl962
Iy23kCsVNNbiIAL1PCLruTXQie3wR88ecVdQY2pFlq4yyaEylX9mbOBb6t0BE41y
gZHIPgtcgp56M3G8riRe5Yu/15RWUATEIEzPi9vLPCMLrNjzFqt1W5YuYVLH6bbl
Qoljclny2z2cnQt1qFifT7XO1csg7sNJtly0aKE+XEA+wkkVnrK4nMq3InPnejj1
KvXVY0rXMbidbAzchvisRIjyYfXYpq8O3OBEgIrf4CCW6KshthhFy8SWgRx1HoDp
TfXXjV759WMDjoonBqBXR+SWUEQ45Om/lmmd0TipVZWMt+kS5x2WTCIPexKXIIJV
YE0K6F7gwST0+NVE2XScz93PeKub8fXHLIWQo76F8EHwJ6aqEyKQLHyhPYHuKXpY
84+twuVSDdfisTmZeir7h6umBuJCx83uYa52Cu+MmppHHGsrox1BcWZgf5i91q8S
Q1em/vQH1x03kCzhvaNiFZLRyYFN9Px2OKua0JWiBq2wJO8q8AiUnapXvtZVWG1K
p9Co4JhMo9QMuf7AxYXUQRfPBj6vEriJpD6wOLwCQUvPTztqOxEZ0BSGWDtnvGI9
CbQiJxJAxZ2T3lq95DlUEUVw72zIOe3C6ufGcajLl0teOW1tOt40ytG1gB2may6W
VWNbmjhOfefDInF7iXMWVJyv8G6Aoq65gx1maCnMNTehS6dv4nPkURtwhQ6d6IBZ
cxsLy1g36yZ4DPwmw7swbS3mcCEYN1hBRSPR7nITUBhe2+6N6p9xYGHyEtyqT81v
i/9w20iibiLRkBjJpoHVuu1FxGQdfWwvL9IykVaKuc+xgbp81NotvaR3obkJCkEl
hE53vg8LPiacPWpXWHMm50yA0abKiC2P1kmzYpPVfm1WTRYfgi7TkFlAVDF85do1
GyMSNHk2CH8royD1bCofhC4l+RuwGDo2E/nRn8hiSIAD7htlM0BB9v9ALSjuKmdL
1rMPx2EvVHVVrtRCJ3W10k7TmJAsnOkJI0gQzFs8yeGC87Mewao6nLqeDNzS8g6W
RmlxsTB0GrANh9/suL18IxVaEDmywE7+/8gD6W5/xvaND7tL5iA7KTBCIRR53mup
38/7IlU/3Weup6iiDf0HPjsOSpyuda4JPQvgHus/NhfJ0EzZ4j8kO0EtiZFtnUHG
HpwHnu8ZF7zoOdFow+EsNhO5Uc95uoPesRp9bTZSwTf4/nyreISsEE2dhs3qSl1k
X0ZszIjpy3FMGO2nSg1qju58BjaCjTk/3wEwYGIiJ3J+3owQ+E7HChHE1LdytfaR
xzABkcOluGjtru/t0waVqPVsTnRhHzZJQN/xF6jBrbTNLfDJ9SZTgM+qODUdAUAn
z4mUogn6QBGFH+zM/Rd1xE12HHMzOSfaDJLOwJaVDzLrGxI2CPQDMabEIWBd9KUy
mi8/CLEMMJNFHG6Icpao8MI7jexqhAcWIHyISHbf8BhBPpfiAK4CiDkRHglkmxlo
jX3kOIdvZzfT/tr/cqeJP6uwiIRVGwfXNvuLh0bZWn3W6eczXcHsycy4eC4/hJxX
mFODiv6XyxOiHTtAJNZcZRkxP2KQTd0qjRtv1fi8MMutLkcPk6FvjCIqgEltVI1K
NPj6al9zJhaGu7jZkhoObwMFy+yjFeSNHIvblN185Kejy8lIcMx6v40kB7Vg6/a/
9zn7fbpPJHERhzpB8u2By4F7A8qRgbtT2bnWjjJumaaT1hQrufR+AhSUAR69lIcd
fYCJSem8kSGD85DczCj0dnA4WJWRj43MIE77v1zgRYYd1PjTTVqD6wuDQxLqZabc
xfWolaNefssYLdWf5Ps6ZAO0jP2cZc8O7GVVt0/zhPSV3Zr/TMoRtat4EgYMSFZy
bmuCmqPVJ89n88GOMr9wj08kNaAiqbOLxS6jyez3a5QYwU/hMtDWQnbtbYCq17zP
otRdm9XMnnRlap+znFFW6PsD/4L4+Jb6jASdZrxmyi7cvujqIyoMSeVEKRWYoDvQ
R1OcvvhpKOrBad/EBl+mWoltiAEdpqUoehCf1vlaulY7vAUbTkCCVsbG9MiZeJKo
hKEuSnXorqO9W8YMJEj7tBpEEbga0zqX9Xio12km+Qo5Bo6Dli7kd6/M1k9n3xyT
kyxy9A2UMgIxN7IFY1C5fsj8rLO6d0jQDS6yHJeB7INjgqUyfoiq7dqrtehfB+7J
gYAqo7ID/5zuD0iQq4RVxTKhsAQ+nZbbcRhERpzECWQXCwEfw2fmdQ4jlLoJoQVc
txrCVNDhsMAYtc0xctdhMQXlz9W2oYqPVRZvi7HLZB8wfQYx9QvhI/X3FLJzowNF
3K1N8jqcLSCyk1zfWJT11a2Al9IgvpmFuOyY4tk1HKaAR9lYeWRsU/qL367ecrRZ
/rj8CCwIAUG2qEgmgSYpASGCM5iiPp9/1t7fESnh9dZ0RoAzi0zjyU5mdjYl9M4V
68DBIIvLGjkpZin7+CGUjR2EnXALc9FMop5EAU9S24ClTKB7ghUdAOIMCGvoAwSb
+KpjBY0RdS0IZW8bdd0wgjyR6LrNnQBf6m+tyiU9tehx1PjTgPFbCktYCkQ+Xo1r
e8JcHJXtXNkKL0tCfUFwSiXUTcNYT137uzHUZAfYY8Ma+EDExlIyQVOaZ90Hdvm2
lTCReeBP3jX59C/Cie6AEpbnPXlrlgp+sfAhwEbKkJA7ZKQmi8yAgB/3CePxzGsI
mx1b2yEzTJeiDqDZpsuSHG80j/CqABnSJ8vy8+r0NITyXn6QDyy5coIBZOWUhXxz
Wt9e+GhrBfDhCL1zrd4bXhGT4V7NHGK9gJBIG0l6mtvV+U83+vRdR1zsPIn4ftTl
fviCL2KMXqd/0Cal+D2orn78IfE2ZnCCRyiTZ/VHffDQExWUlQgCHWf/B8nV0tC1
OilXolRXZQulTM/l0ESF0/EmcsXIgEBIItBwAUTjYJf8WEl23MD+JHYphqm2K4es
s4m4loHwMuPYne9j+g2rRRC82lIMOpeOBA5H4WGV0iT4eSqxsJklBSMBtzk3DEt5
uJhvOpaHAo6nDmnhKJrcGJ2CbcUlqoYuZskztdEmWN7NyCdbb4lBDqy5z4X0YUsG
qSywyr79A56YyllOgMcf2uCyyBYGQgkiHz7Uz+OJrOoZeeLF9tE9sJUc5x6X/9oE
5PLyxeWiPhNokHDbkn7nHdmbKd5MitJWWF5gjmWZ8QWpqc5bdPT6nSCjmtGAiil6
hsb37RzleOKXM01B+G8TFKwh3yr90BnHd8GCrf29Dqcbh3ICxqSymdpgFeV2ctCg
TnCeNBRhOFHz9tRuPUMzI14fLoOtOcvkmAaddXPypfPNMmjv/8R514eN8xtf2cuh
TdIbXfLiyxEbQ4Hf7rvPulfuZHkJke1yF99NFj1tl6/G3tiIRV7lb969ajAEJUTG
zd2bARHwO/UhuXmhKdkG8Ss5PEI7fWLYlUQ/R9moNip3Pe2hAv6BJ8xO4K3f8sKG
wYxE3e5gaW6iDbuBpWjx3wfv4+EB0dbMRVxCSN7595lw5M4NbPN+qqiuCNZzlp1D
AWrzYjfSZY6BwfD0S7dHyg8NCYVMxlESO1PtyxxGOORdBnVTQGSj5PNEkHFcp2CY
yaK8oaHKxqOnM5g2hFCr3X4d5YebTx/cvF8ZH/B5/B+KsTGaxjFD/imzAr5dKIRv
8qu971II2dZbq7ZmHgLZoZOS9baoMjGUZJeVI3THUlNTmZd0RzfcDhoyl6Arcca+
PbZ8dvAkA3/L9XbSmx9ULPTr0+TV1G9gXs/pbXaKF1v0jZzJ9P5YsOWXb/2CtK1l
ClkYI81YTYCPSkyGcxygFqa0//nWPd6yScNH0wMw39KyMsAT5YI8cRr3Mp2pi5Dy
3+eK/EFkifxAzqHXnZSTjZLJQ2spJR4/vBLWGcvmjpHVBVezyl/rAu9X8sS7M9Ah
zp2qAwBeRRjdKcM4uwVx/uJMXQ1mnEBDoRtWJf1gkFiI5gj8xLs0Ph5R4FbjkQJZ
KhJ6GGZ8HwZ8//hnK5jzgg83UpQwpLklweuE5p8PH+UmObhhj+/N+VU0eAUgB9NY
tM94GEKqB6qJC1tUq0fDCnAaixyvl3KLEDjBV5KSAedLgkzGCbxAozGUWWEnwpYw
g7q12t9vfs8VtXxfPVpVH4GjplIxJFvQmU14iNhhr6Oo3yV80vi8KlSX2c07d5Ht
cPRwFP0ncXeuu13dZWzLmjD4TBsP1NSGs7A5gd8QrHwgMuJZaTCT7ieiY2TUzI9R
9/wYAO+E/bFsqEpIPXq/efT5rCa5rpu1jN191PkSzwMEx8ugVYnnI3H88q7dmmSs
9sVQH71v0RQ3t643w94AN8OFGVtbysxgAQikU639bDTbjMALWIwt35UjFqip4vo5
UqOPdd+AHQQheLtKklX6/D0D7J/kN3NEsSqvfUbn+TtW1LRK10UNmsJZr0meq+4C
mW6BAYKjU65BI7oo1OrkjMmKZGRJIz+CQhP1oBHojpkvALPFRRcT1liS8ncjRXe9
MpWpWodLxjOf+PDEY64qFEEZLmGYjAtLoXbxFu2F9n0EZok6CiN8vosjuP7pjDiV
GV30pAJ1F2NjfE0DT2kKVEsQIu97mL7MQpBmNL4jVpUOW5eVFDrj2ycQX2sSRBR6
mjCUkKo07Yer7n5Ys0rDHtlAHOX7xspRk4FHt3u0fway6f9VjxLN8LNKHCGDmOV+
BT+ZutkgsUZDIXT7yWGL59ZiHPLKaQlps5454P4GBuWPRLVRLtPiGIbvIYK7JBAz
OEjrAyj66z5bDg+BG0xZlMob6tXV43UgqEt/PW8T+yISkErBaGa1kjzmwvx2Frbb
YV3I+7uQC8ailc2ubKC7xDIlkjzbEgYkJqSra+6iHRIuij91d9NQeR2FNqWNzf6A
tIOCmM/nQzNAtOzYaBsIQqbaebmg7pUxjOVl+vymFiYupYMDstfUGykpIbfGdHzq
EkGhEyHNqhbYg+nG+G0++wvDYaiywAGfTSnSZCyd3AZY6538lHoV2zsQnzOdYWTF
OtMjfqBnhx07YHQE13HOES7pGK53Nx5mz6iljsQbfDpx2eXBwsRXKw3vRV7xyFny
M7yA6hTxNohFSQUy44C+kzDf1oND8idjrJGtxa9hjePSGBP9YTspiPb9R148T52S
3wMC8A/AXpunzvnYs2X7NEoOAXrDXeQT4iQRTZ7f4z8DixjAXBaUlZzezh5O8rVU
+EwUKedlVCHwZNLQIvQVcItbJAE3AH9Nv90O/JvrwrXThGcNqMtAzNlRN5fCYFT5
ze2xLkP0jwsSQntumVY6/kMZLfgg5RHmFNmewEqbR2licy6DkJh+hwz/efbypLcU
5k2KJ/TFqujeQIH7p8WrQ813TiQApPVOv4ADzp4TZB+U5282TUsDl0CkA5O+GJTG
SF2LYE/vlstLYBOxi88JYCfwgGzgCwBYcdxsH2T4DDHmP3nVeTL8xZphWDLFnYsj
lTwr3fiTWDzaRbCN+b5hmfY2yr2V4aq+PBjRveo4wIH/jzvJ5g1/GgJktvUEfpOX
9SGeD14gJrkPzGP8IUTVcoF6RIQ/kLaYJHdIlHyhqxBmMSemKy8thSlmP9fzCNO7
uPStSZMqLl63lk3zyvwi6fYlLDwNJU3mHo5rzle7+5UP+A9sH2enjxIwXlRyz/vS
AVRL5Z1XFwalPC+TWkXCLx6YbU/pYK84Y5rLg3hDmoxUa6p+sYrycCYfV60Q6VY9
/pmZ3cEOQAjb9B5hR+KyAordl4k9c6p4C4rqwPYFNo8k1AdaxWlVHN87XIFdjJT8
sBV4XWv59gc8qTynbVLeFbifVSpurpU/gK/8FrD4KUyKnXI2araA58UsoZBRJLBF
DjyVbR6GFrVGxPtMHjj3tHN1mw4eXhPA2HKn5LF9F1yfhxEuhuTw+yneRQbotHZt
opT9T+ErEkBwCv00lc534NMImHW/1cqCOthpo6YvIiMbn0apsdPpdKwztJ55eaPY
PaKkAA9hrjQTm1HpouAaj547IJq66YcKDwENGnLpyuJoJ+Epf/Dnd4kyZgLB5t4G
DT3RAk2Vok3UtgVIHKbEr12EYK6rhhiGZPwDbVXHoISWFUeCuLLa0lhQpz8C6nTk
UN6yrsRDRqDVe/kwgo+vW9kMIPORyVjHMNBN6qRgAQ5BXsCC8BgzSho214a1I0oz
zgvc5/U4ZCjzVpjwDJWnr3JN+eA6f0TrxdCN4qQom9bKMc6RM5Twx2LMHvekVW7O
mFERnsP/wvl0CrIj6mSSWfmbX/LYJ6PwprhiphxeCIn09R/y61flei1Xh1QrBaD9
js6oTyNhKJgqIl09jLJvpkNFGxAz0zjafm/QUHFcTpMYOixmNLz9IENXqebN5DAn
XaLyjHKfbf4ffI5+/mKd6XwIjgHFamqdfGg8c/Dagdt4WI6meI4AK+C7aM5S67ty
vW0WRgTTTzESzL0NwvMBg4NGYCtiLgfkriHOGUtg/V2la0fuvj16g7/MqcKfV8Kw
yu5DKz43I/t1MX1ixVtgko3mLM/dJFta0o9uBSyeP9E=
`pragma protect end_protected
