// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
Tp7jCNAgSOZrsTYBRRNgAKHVcPY+M8ZrdXIkI9fR7iwReHFzfLHDek6MR9keTddy
lSngoGsG3Siv+dL5NMI9I4mSrc8vfMnkFxCLPLuXPKVs5k2aLxsRBq0fJCjz9nLJ
Ij5bR7r2Rh8U52kZVPANBVlF1QUgaNNtIpaY59UjoGg=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 99808 )
`pragma protect data_block
9k9SPtqLYhg8PELaOMz1Y4Zh25HTeSt7MEGQ2q7yVzVMvsy9peoBe8D8cV0ixK8I
rI+goVJ9r3Ja0f6NgKmib2bcrzuNOwYlni1ovQYuUGlFDnAjba9VSas8IT8HPdKY
uIJ915BQTNU0KkKVbrWP8e3+aADbVLkdj4wxtCQWyM2slBxfpFBJmeGlCoiJ+n0X
k1+8jQrnLKU+8hKnonXekJM/myfMVDAUR2UMyZiVIHS6jPRb42h4TjAvTA7EuJiE
RJJZVGLzQ0TgGKr69/bgGJTfKaVhzATOQ1Ee3uK8KVKMyJd/tk5RKWKqpTLccjXa
YK409AMon4y4a3OD+wsmOen5hJ2By3X3l1nLdENMvJVrPmVhUaRLskog7yzqJ890
8VBWLyNFDBQVTuaqQbEDnXDBqb1WiIL573jPek9klLs3JDfQwW8vccT9/rZYpK2a
q4EgOnf8CdigxRoDTwoFAuaqjQ9X5T7UFqQHo4uJvSzCP0sL2jIJzee8OQVz1RKc
uVCxJ0xl4jxEXVE3z+hCm/4+zEYFUK2HHtAZNY5CMduLBb390Bt52xih8VY381Ds
GMsgV3xMwxf/ELckiOkGFKeDV+bGaeaLvxy4irK6vlQghNdlnoFg4EQdgo+VaBCp
NXEdW4FlhhaQXs1QUNeuB8DoCHppvOlJMy3npwCif9WbChiGRkajCEBvSu3PdD+7
KUdCx0SQCqn+ytxIfDPD9Bizvx4Pbq5lnK/dMie86PE0vempd9zEj6WKT75YyciR
AFrJHjL+bTH00389a1ZBfXONLU9c1V/98ZDVImMJAyR6ADYeN48BV73Ec0jrdPCU
5i4Ltwovs41F+npAiPqwM3T26xUHSPGM/a8tiP0mmS42i4Csian6sGNrpvZtauLf
OtzvrlnG7XFErw0bESUFsArjV43i9tXyx+/+TbQStaiDWeolY8nAJN4RShnodyvJ
hvHMXg4pu43yMeB+RCh7/yZ0nGd/fOYpptTaY2KFEAZkBdD7/9BdwO0PdMWFm+rP
+/yKzeqLaIzmqja3xBF3ZMRTAIftMXfSGRXOCPssHafk2FgpvMfoaWK3CL49HWpC
14jciqr379zkKiStP6xJRNQ6NVok17EPKNZoR6v/1ElVYsWqcqQ2ZX15Ym46uk+M
LY0hCgqL4cQ1Zo5AOwOVvpIrVJlPNd/C2ykLWum9sKc31yBl3k3PqluBFH4de+5z
WVOshNys2kLvFWAsApJWUEq7l3zVirNMarahv3ORiupkMgaOIFIaQRsDxHGpu1gA
xVqq1GxHsvcVSFPuc9aTx23u8HwBxuW6bGEQ6BjAam26J6W94MoGxN58rzNr/qJc
gzY+rKHA7eAFmECIFeo1f0EDAGpaRz3wdRPw8ri+k+GcZGuDZu3Uk2jWErtySWGU
aWpLx6ykwyBDjaZisFylOOClKa5JZHlxOeqZHnp8dvl57cZwiNOS8Ri1xrazrIpy
qo+WH7S/L9fyd3TyCySRh4HzdzDsiCXs/Z6JVMQ5jiA5Slyavf3QrE4hAnqDbhE8
Dd4SqKANgWb4S00PjSiKJJZhSTMPND3jQ+BPDHVHuNRmv9AeFFnxrEtiPJtDiLuc
2iEUUP8kCVRP48LJ4irKbhzOnPsqcgaQvcWmRliImZ5Q5Xv4AYN7rlWwBL2r55KG
rdZDoXFCwyaQMIpY/+9QSvZUrrT2yuLjgwGMtcop+PgvdvDXvzT/TH+l/hoeqget
oDuk6af1MxB+Vsf9/z4AvpzSsPf9gSmwuPoZdplTq8dXAwU4MUiSIvBrXtXC+EjZ
tbJLX671Jqfiq7NOO20kCjzQNIV/+WyM+oUZfbVrM0UoC72ID69KMeYNI0ovj0DM
LClxAs1pljaTlcvwCtmx1TBFR1M3/pXm8H8PtapxqXCGAI641By94IAQ2W94p9sa
Y6nrO1/C2QZItBEftamQiCWeIPwwPrRQCIGh8rKQzJ/v8ajBp/PFBTfoNsykNKZm
15gk2XacbBCE/Da+fweSz39Xpba9z00i9c7lrU1floMAQ6V6fu1f3uLPpumoD41S
JhEoX7S4+ycawjFPHhPodwSsTcqtBRZrf88QZT6K3L9AqdvBSqBrSH7rFEOVEG3r
0RW1Ju3K53aoz+I2QY3moSexJIxBKe3iLSMPAHS3ySzl9LBuouAuqAU6k46kXjjp
4dsTTua4aSmKDnALM76PqA7RUX9j6aVDGikn4vQh9byVlBAUaZpcbw25HcF+pPlh
uQUDxl3QfyM1qPUQArkZJvy3X3N463Q+p1J3UOXP2EMHfZFqAbVUhWV0FPRySvlu
vGLYa7l79zHke5eTP+3PftCJorS9o1UGKcspY7CXi97B5rWvtzdzCkslxA+7+/lJ
RkGwt5cj2BPrgYlA3zP7+lF2UUyPTObW09tYhYFy4Mq5P+vkIcjv/W0eCRjDYbmz
E8E3pZJ1Vzm5OPKPuRch/b9xH5IIdaF+Rum6pvi9nzFy8JvkIo7zdRC2OSvZScMk
ZCfFhb/lnhPMF+Bn3REXEGe9B7vL2fLA8Q0/NVLwA6dQtmi3KygME3Fn3F5qg9x8
qBw/mh3MGtT7CXVwVk9VHlW3G4pmaTUm5F/lZD+VXEjeymlAiYYRAbvZj4ZTl4gQ
ihfAeaUfhipGgxrhwDUgDvYPyrBeyGJmwPzRlRwCFzehHdHISChqTaWoAzBCkFNp
RypcGlZnrPfVZtk9E4Sf1MKsaHg1dqC6gkcgkTLV6XIK5A1kpYkgXLev8RiAjR1C
aDDCYs9tj4ZyXgMnavmltwERdKPfBpcWWzzltLIwUX2vQJu6gkh+zFsYrr1iqUQ1
erDzPoF2EAbQZ2TCuvCsloLpL566Byxl5i0G7/M0uz6dPcwNesfBucZ0ropv+sY0
Ok7rmyDNRJqBCQDwZRDAt72v4BVlEfOdhmtjmnit1Nk4ZXPkdf+YdOXnKbI1r8xu
QdrduSxTWX5gxmH3+I7xQFYEWKsUvCPxghVn3dT3oQbVwQ3VXJeBmQQPeg/LP2xx
cnorgUfmNBto7Ut4SVcNbwWE8UxogUaPCkzxczHXNihRIfHverz/DSSTJWADdaYc
oBvMWaiRhkeRuS3qMK84iBtj31GOIsugFUPkLw4KfLnGfHgWk+TwJeRwWS8pUBZG
y2lQxACk7Ty5r3smm7S8huF+Cy+ChtfBh2eslNvT4L7kVkXSgtVu/3kNC0JfRv3F
y8MUS0N/B9hN8e40iwkPzbFa8eZeNKlokJiOTNmBySj3kqDj7Mp+/PVlBv9BzymA
0USNA+yWj2N6TI2c6ae+q9yIf4DAduI/XET9oxNOIqv8UBLijsbf1+R70jLPbc9Z
9YiPRP7A6+hQaAH44dqPIYL6YSUVuKKwckAn67vtvBPaNao4AJQWZ9X97QWzSnPl
3FkhSZU7pfHDbYpawxPDRYWJyFZhFJPh2m02a5IJLN2mIKqtg0DOAt8KeMZvce7V
/5ioqzw2VLEk90Rh7pu1waIP84W6xANNSYMt5xyfbFQh8p+ShYeewFvnTUMXmgjC
gjbK5SVFD93y2s4NhidyIzowColLpGyw84Pnzj1JIHxpNlh+VqFTr/kkUK8vrC5n
eLc0MLy1lJQM5m8zBWytXq+RQtsJS3cMQVxuUN7qC0T+nB6rOYD3Dz1yyC3ur/ao
Y1hz7b/KfC25BOog0peBXoe8iPrH6jhOgMHb6B1M+S2WFmPVb/pN8BiUZrnOjK7d
F1BLQkwa5oN4BDxw58lDBAQsRPtFUUWZHDt/9q2OPOkez55SCaMzFd6wzTmQzK77
t7w5I2XN+c0vyDFH7ZppBMD5zZycdbfRyTW3oio/tVSwbdbdjO3m4iTTTwLObLFj
poZfdEug20N+RZFpjgyrRsQ3CZw8/vEShOt2F5Dp0KADVb9Fs4f6eNWChJ56ZPgq
ww92BmXJkPVwym3t3aQkLB7/00ezDYQLqC6FObef7nYWCHw/vq8zk+BE2occ0xgY
xQm1fRXIh5TlD6UQTxuO3ps9V+548j970x8n1qg1WmAx5Te2yBvj46I4o295VNgi
1eFqzsQbFDz/QSAwn3fjGprH+2X/fZpS2FFKEutV5p6qc/gKII6MNit3ExU218Mv
oFprBXDt53HDOkKVIYLE6GUK56HRckg5rZdJ+9iAas7+9SBMGLDkQP23+oPqh2x4
xdKo6J1znT+rzm35rF6Xo6Cck8JZXq5vAAx3g1Z2ASNt74JymIkvum9xJBeZpG57
ZtIROf9ec5tsV1RqFt1ZEswEm1r6nLqV83ecYfj0EqOXQZmGD5TadbicoedPiKCo
b8z/YsHvemE/eQ44PnZK7eJFd0bAJyOw3xgFYbCsUB7kKxvzvcypcXBDQpehlsgq
OmRKl40P4yt9aOnJWW/L/LgUKudcXNgcNv1hsqDwpPFUiwXbhSWQHtwrqTlRldR+
upRVTGhb/Y9XjQSPRYdM3WLLkZbIBAinRMI/15wBLy+nawqPmnGpP8LH11w/j88i
z4goVAexF6NCw82F7bdXFXuwAgjzcxCOF915Em5ZvOzfYEQd1IiJo0XGMtp/c2Hy
1b91TQYBNIrhYoppYLCJqD1SBVZDAccXcBM+LrAH+PjxgFVlIeVqh2eiqjBU13ZE
YAqRqZOC5FSD4L9eIof6Lisxek1RHsT7FK3GO1rIbFrMv631ByrmmiXo4K+mEDD1
sGFSTlrxzrOX3YGaywuFh3vVmWGO03u2EZhs1pKHND6wxjdRXJq46VKbaKZ1jamV
Sbzt+oI5VkQ/PJt404L6KVjF1PGw0dj6ureFea09qSRdtHC0JG3BkOOPyrq4DgkV
udUsmen6Y898S9RzVsRp+ucCwOk+SdQn1eeMK+3mWQCDu6lPMtRJWNUSR1vIlemW
vhP2N8PyCeTygXSFFx+wP9dgT2rb4TKq8f4Lt2sw3fRhJWFsBXEhQJoprQnUrqR/
8Uj5R7u8dAU5VYcNrQF4dBcX0cAPOyUImSCoL1PQ7gah7745RkvnIrptUWmnzSiC
TaR1srbRFg+tnxvblTCuO2jiEmYthdbbeQh38Xzg+tpwwT9rwDwAabnCActZbC3G
Ig0rRUTXxg+hqoJGSyHYYMm0YhGUdBP1oBibkoH9hyenbTXwH3TH0/Nx/21ytb1S
W/HlDcjxIbN/Qa99qzSPkX7QuHt5GwMImq5m/qr6XVRefZhFvOIOyjmGSeV3wlzf
bPa0VPVxbwbfBoPVyttpC2GLNOeZr2x3as9VYdqkcbNPRfZSi2V3RepvGG11qTG8
2/RDMkVtuIcdVvK/qHQbNZoTe9f9KiLFndwXcbtO54o1IYibo4CWBmg/K+yYL2oe
iCdFoAz/9ogjKuGMiJQ7jMu5VaziLsiIm1XPsYukPGsZc+avfOl8v2pXFDOWmvs3
nN6wlRxv+RxlmQRWzXADBydBCkDUPUi5xScmcSN/0PU5wiVfPIr4QR+1U9wPVmv5
LFCqYShSMVeMiM25/+fi2NvN3tnHkKKktqioqqGlNFS+zLJXnePfFnaJ7ZuYsnfs
9WpIi4Bqnwqx70TZt2YDEcebEEngz34upZA76d6zTQtFwDR/BobQfauyS/u3uetB
u7+dOgn4K4aLSU9U7NEoI9/04TYKksaZ56AJM3TqqUiN1GrQxDa1GEjnDf78QC5V
vVZiMF4bezaIeqFEhOAjXf825Qz6iKEo1E8sTa4MYFxlCzp6eYRyqf2pTfGzqfrN
4oUXv3BxvsGqV+f7xJdo90wMjPuvAXuPvg1tA6yEbSIc3ip3QMsZXjdPuoqxzEjp
EhZM+QQf6TyA6bMmvAxSWw+UanJPMXxrl/PywCwbpS5PTkXb3ULpmgSPDmvT1Vc5
uN9PZSTaKwODPWmEB5jYGJ7CszRjZxBNCrd9H1vF2G4g4b8IpEVQwJZ78v0l8Ilo
LAeOMUP18cEH8NjmAyjpe2iC+oxHum+YnuPXab5os8K0rJ3tl3yn1gkKVzx4Cqxb
O0QStQrAHco+XT4m8xTZvp7tpPCkV7cycdopBvAbbXaoUbLyJ/y41V+C5aeZqKZc
Hql6/xcQTJaRzoK7iih4Pz1F0LIAHcl/FRSJ6KlsNy1ezyUXr6vfI/xN1ZI6z3gq
2Xf4MmGvzDI7/BjpHzMIbWCR92Q9SFozS+2PszUPt4OtEfvUiV6ANNk8yidOIwQ/
9EHyoeHoQCeLaXSRu6oB7DdXxIAd2g6UsRnG5v4o1i6orfK21o65kzTlz5XtZASE
AiK/wYHVVH0TWq1M80LrodPwKetMLfhi9OFUSxNmO0AA4u0GoNVFI2qJK1X2G3uu
AeIp31Wi6LeUyCPiDk0kYi557wz+Yrofii8cwsgNEDFB4QxeOYUB5lGXYEW5gVLV
P1CORv5BzWSIgQsZNcq/pHJ9JF5CkRl1qR4CWBKKCROgz96e0RoCtoXHVFxYbva5
M4R8DI4wrnZ619woYvWA/flLSwTOEvtwwhzk1Bzq+HHiiiSCIqcGNGeFp6qmWxTI
xSAzYrK4ll64UUnKg2FTMqtHzBKbn860XEvcZ9+25GXENOPOFaRRtX+5RgYb8v7F
6hDhvuVkUVG/jVPnR588+BMgQZEZF7ssw1vN/dNq2YGDyRZXD6Q/ftrEDR4W0mdF
WcsPmzPTj56lNqEtBhRpJdOjtN2ozrm9Es+7C+Q0kn0PTI4Py/cMTGioIabaBjCN
U7BMQFATkWt9k7nmgLMac8WU1Wf7z/mOFS0J3lzD2R10U+Q/eag//uIrC+2lvhih
x+dAr5R7gW0ZdXJ/ZDLa8IL2meXnAImvJKWRw0Xt6j++Wej4jVogLYBXKMvSPQNG
34mU65OSDDEC9RUMT7i4VgeNDRE41QRY+7f2/2tb7RGsShZIULslxqd0pqyefd7J
GtijxFmgq0NS64iDgLFRsKq/cpHK/JrpAMPOoexabFtpc7nF514MIBDMQqP/gSj+
E1A+2zb0P+H0rP3liHBJAZ8BLIYMEdDJETnlI6y4WhQhdJbp3yDpc3tNRS+SAyUB
0qw3L6NLLfVUCD94+1MOrcR6Qh7SKqTFU/IFOG8P3kU9uR8FdCHBbr0nfqJMVaLQ
kxhYFi6YQ3rCsG1pGfYIpmKASwcP5Rzev058deRNn5WHaABCxVfitF1zXAhESXPM
ergWJNybIfv7k83aoRTj61/QTuOys+/wVe6zF7Qq5ggu2jyEzvloghKardNxpBIv
MEVQ2lzCYoqDflVbr0yl5Ulh3S6QJjuD5ov5EyvVivy4gOL3emxael0ziBOqHASr
vbOsWp+qlwa8ViaTe8pPhLb/dSXnubOmkMmiCqfPGDlIg0QpgPzlTMGqXnAq3hRt
tNuikMWeU1fjvyukwktpYSzu2FHi+/ofxl8/dR7bbuKOiYLLJUnQFCNOzad57yU3
2SvvpE/bXu4gg9LPudzDYbRwsd3H4BmLftvDGWVCh3g5SnmKVmTxErPtJO8urZd5
p2I93gx+zxVZbSZB8YMxwjkbazGC/gGDDH1FwEHHwRxM54xFTkJkx6KP25te2s21
JduWH1+4keIW+PSKdFpWBqgjidstjyzPe01tOYmPp0pKMz9zbPlbCL337Xd6+5xf
VV4OvOw7swlhOEmk9Cy2eKLjMJGqOOXGmxG4kx3ndcrJRcXcRXo/8gz1KyBCNroU
OXNT+DO6yRrtOXdfa0ABGJta0GSPH8tK5nGG61WWQxuV+hIh15dbpEBjecnAYMXE
auyAYSfezCjBTLKt4aXKNM3hcqBeyFZiCT6a5gSrxd9pynTtRqVFqHKCgKV5mstw
J72Pk3KfQz2cssYqJsHCun+CTFrgwB8WFNDD33T2Rp6pe4T/6PyJcKjaI22rF8Q0
VNNVgNAOzV33X+bJexQWMawTwR+l3YtD4JAw/vntNnVmIOqoQo4uXSUL+RhvWv0r
rI2qpTGS8AN2SMY1cP+PWKemMEZolpqkt5sghNxYOdbQ8R47MNii8VPx2b6J6i/s
vePW5XG7d7AeMZZl55v9XZpzucjc90pO6wGlAFNgB800bWu63R8Wm6NdD5ynkYfK
14ES7h0dOQBPYh2LatYVyVwmRI7mDe3QkTtxrXu78RBmpEUm4sWw6uOQJrbR4Dat
n3fv+204e90is0MdHADNDz1NYRkFlGwHhfiCO0H75IieHuGNLmeerrJxoPSIw5AV
6N2H95kP9PAMVDbrx5ZUKLBMDW5x0WYWKx4Cdnz3SbmvfAa3pao+YNHjXO5bFVvR
Exama7KusA1CuYb747hj53AEJC/alIHbDOexnIkQ7MWgVdLxz3BEkbBDqmN2DQWa
9q62g2rNlMdGBGrG1zU9U8R+stWYIyaD3QwdBod46OS0RO1fopGx/kqaVAaw/+jb
8QW74Yh1zH/LKu277NwFLdKOak9LnUWjcSqEq5Ibb83kgZ4g3fBIwxzhwtd8o3B7
LpBRkcczolVAlU/mwYeMhp+A1Gluva/YF6IpjZ2zpZdnnJaldlMdcxaEVQQO/mUc
F+zFDuT6Y4W6fTrKHCJ6msYLNsT4AADc1jwjTlnrnFvi//YAhh7nnhB4S+XJYUtn
0Z4zpI+Io7Lj2FhjnQYDr+yICuZonie+0iBSScuHuZkmX72WNRLKzsSRoSnH0iaj
D87kq3yM9ITnqZ6MkSBRGb8ne/lo/YUNSQZI57J1CvXhr/0HL+P+7lQtqnTt/7/z
vCx5ftg0L1qxww5r+nV2jnV9coc0ZVJk8weCLPTyZ5tzgXFn2whdpyqr0WMJFo60
tROsxMs4hEpjTXH++EVzFwQqhzOiPG/oir6ew/ktPMO8wib9k3cMqiUJ9XocXkqY
LdJI//umc3+TsnGhMBg9b6cLIXazplw26RjTe2/VJibscMkI8LcR80UChNP1obu7
eXCU1vu/izmnZ2CgcUA/vl8iPIRt2m5sDjZ9OuwFnw2wIOmkLW+MVMGPvWRKz3mI
RuhBzzGzRDg6oKNCKJHI3Zux1DRySKh+0cV716jWB5E0sBqh3xwMHubQUd0R0m9H
58m1T7asCUyC6YTbage0+wVRhOAN+P6GhDAXbeGUBPFfpZ0uT5pUgdbvqmbUrr6O
19aWv+FsT6kR9JwuKzFXDTOZE3BEcVYtQ/5eiwgyOrcIUrH7VI61lHD34MDmGrBZ
WbNQN0aIo1KdYJFdpZtxtbGZN4RCWYqj3nTiGTdHGNhV/bh5qOf6+3fzhUpLQdAu
TXj4NVU7W4azBZmwv+4obc7LdM7fpZjQnLMmU90Nii4cSyRQNFGpOBo8Nejdidm7
elkoBax744lQq43XmHPVJYi7IyOyaQzkg8EqvqqTr2I/j2MyfSjNhdsgWK/qui/C
fl1TsCfflJ8kaXvpgd/qGXQwlnmMrSeMa+DpEDazmkndSmW/uE73ibxGmetXFW3E
MENHeSaGgsnD8f5ofEK2h8GP4VkW1eSYJzw9ybTw5Ek3miNXwwcEJSjlGvokYdgs
QoPRohI2VqE5C4LZsYqyXYuH6LYFFXPJFRHEcrXl8uxs/5jjfQkib+DuLg0Mwys5
oSekZvQ1UJBATiB/7XkXmjmFMNOd0lU67vWSeZ3SdogQJR6XMhK2vzFWXbEyUEpE
CyDXsR1Br5jLKvYq4wBgiIW3B3N8sE3RDssZTDGfgpUh/NHcBfNxrUB9TdSBehE3
J5AHUECYn5e8phwDHgFTq6ydeh0a8l685tct4c00fHKCG2BYbRk6aVtOItQOigUg
h286QQikGpDKW6t8jyDbpl24Nva5r0mkoF+zBmjvFZhrBBzYrjQuRYrW2tFw7PCe
AVhwqNbXo4YEc7LtBiRaMzVf64746B4b0vN2vxQMMk1frL+eWJxgdde9rL6y2L0O
T9oNvw2dZWjLlY4YJtzr25adRqhc/fniQgcdC8ybKkzChu2khV5uniUzAOkTc0j3
Y6gvSiA4EUHavQFU9d3D0UYxEOEjd/NsZhHA3g3pvQidoyM400WZuhrxxZlTlYqM
5Hbg6b4QBm38E9nsp0gsOfWRuWRJUXu/Kw9KSK6n4vZU0YgV9gMNdUH5Pm4VjjKh
eC9i2Gf12FNGvLd5O6eHD/Z9wrEKNQ7NpupF9fw+baBDKFRCek+m7Ct+xDRgHtQj
Q1Ex04QLtrv3ymvPYjqvd1RASWWobtjzudPx9LxqVWhFL0dmrC7DjK8XJdoq8liw
XhWlMbsCOlvxVpR2pc80a2gooCkxylyXNZYU5bFYH4bQBsIkYi7vZqW426ki36Fz
i5u+wvY5OmjxxqiLjg1EEeMLHZgQg4lOqGkLIpzQsxDTqUdE8sAZK1hqYzUW2zxU
+mepQ3QET/u/Wm4SSU2Hg9SwFZwm2MqnneubrgJxPz/tcdG8hkO9aoJdifBxGMZP
LYKLTGy4kIlm9SQOwBuhjPUZiqru1XeNDdhJMfPMV10h4MjNg6Pjd2W9/9QJpXvH
6/7axtGr1VFR68SY+i1ywD2NdJfjBD0O2ZfMckdXA53HQbHJ9pqLEHxWCodq/TGa
BRqOb2CwiB2fvF0wM3IypvTsltIAgPAP9v75ZExRd4uTG0hYWyGhwMV8XjmLYCyA
P18DAil21Cxx5tP89t32uByggou384sQCr5rTy1/VGrEbgkc3QJT2JDm6Camo/bG
NxZ1bEQN38P6IH6I8fQf9Ub6FNQjYoIgX2S8t+wwuXj1uWbmSy0p7fyzuaEFbY7U
LQ8IpweYnK3JmybFv/QNMfSsPfL5LYPEesHgV7XbmEjSGtXyTIykTTBWO98BAqv/
Jvi6DZC07EqbxVOY4XK1qI8QTFBMHlMaMPkgunhu+mcaiD57TfYZfKG2zHL9nJnP
PN/UTtsQckm4mw4NPwdgajTnLd+YQTmAx1c3UJyPk6UpJ/A3uA4XGwUkjgqdMhdR
D7pylvZ0RNCCIpc6r1xppCTt7kIiU/jtLGOWr4/2mlQ2ry+YXC3xC+MYkeNh5Ngw
Q4Jt9tSav98U5VFcMfgtsBaWT8yuDBJ6xQYC6kZaLOISXR2UvNMX+GePlM1GH8kn
lZBGEffwN743FAUkpP/vxM3shsGglEESUCns5wMfmHb3N2Z/QQriveyOskioevY0
3Xh/7Gg/GS5m+Z6oPgbd9hAiner3Ki8G3nm1QFp9/F+hyPMd0RkFicKA21we9HCE
aoN8dMB8qWt4ABXRc9/FTfwz56INmK3wK4o2U+L+/RZ3+GZRrKyIr6kXOujF6KMq
REXUaiNPNiu+y/9wdpnYRsXPiQSxMDo0cTkI4udgDENgbBaIw9Ee5Vmbx2JAa+3U
d34AGPuQ+4/3oz6dXjUn1KOKKL8FyK/zU9wg/K1tQ68YH1U5Le5dUObc6Bb9lYwU
W+VOkcPTp/dqUWxcDj5TiRpJk3ZPAG/e3ZkHKIezk5yXGBMc8U8kzBmifsfNkILR
p9A4xBvaLZo8eTmE7TmW0qnoOerCJQGO7VOIQTzG+n/eu+g0oi/rSZefYjhWPWlL
LHMOS203j+aXYtzHOkXgc54FSbzKl7RIznZe/rWia62S9tcHbWFYDRZCylz1QRvx
76m9tGLv5nyJGAnQlY1m/DOfwwED9WH9e3VP4z/LFmKatzTAC0Fwjm1FlaQPclj6
4+rYhiKGdn7RMRPGpcSk2Jnf1tM0aYks5MYKIf/NGOrLWuSft/1hsgCvPDGa36Ci
ZbkUBkwiDFIngjfl/WZhz03lKZf1PoFwH5eESeLhODJOhUDvj0/Hy1SFlmj9xnyS
f3CsnqEPsAxT4cQkEdTAw+TYkT2nFEUv2Dx4YRkJ6QxximzAOApKOv4s0FS/GQg2
9i8gyHnR6SvmYFuOMtisiiWVofrKWn70KtJ9LRu42yvU0fT94bhJQgECN1rAws4t
3swDGTti50Rb3AqsJTwp13shWiOxTmx2i3Bh6kC4O10jScEqZIUIwOdMo7yk57bQ
ZoOTIDnjmH0PomzL+V24j0ViS+M2Kykqgj9czvPJO3MHmyI/6K1IqiTipyhEuIro
sofIyRfOk8F7nEHugstqXEAsvZ252IH/ygsOYTBAqDtF8Q3HwrJy5qMSlytLFn4M
GdmEkXjCHN2vcbuCoDOfZQlTl25kpI9uTKJNiJVYSUkFQkWcwLhcPqwHlg1iKSU6
OneK7mIPLYmcWVvzDutONMcW2ShYkWJn9Ti0JMTtUMGIJ5puymn90BblkNpveZ9Q
mSgH3L7ymqIRBp9nBXGVaNT4weShADMISmHJLnAqNfzR/AqBU6yUO2m9di5E+T7h
Qd83yZlWckKZHJCMe16jYn1wDbWS13Dm/1kNwGnPsy++hbeUQDH4Sh1SaPP7MSaW
vIdH9zFpXOMBrlPTiOK/a+RR5mBME2TnEIvOGzkv5ksmJdPUyAHnP3RwZ80dyjIz
5zBOeU859b3ttUxlK6gtiWVhXLnDcBiXlkYs9N0anWwD7VA80m7p7OjJorMCL+W0
IIgwTRnxfnoCW7EeinQx3WNCsjEiPK88eNTrjzOf2dkC85p16NT6X8Ifq7n8D8jI
ODouqvTr2fnOFp4m6g88GiLZON6b+dtH599vkErE5QDbzhq9JQgHnPemx8L6Dwgu
pHptzxSsFGul7hC8uosggm3dYLd8d6QdQs4BwgSYV0UyZXKS7cF4OVp1E49Kn8cV
ufq94WXCOc6hvI1pf4vRb/ks+G7eWPNkBHuGjX+774K/+So/i3LBx43p4Sa0b0yL
f/UvpbX+U9syZNKSCvPQR1kFFvtjC8KsWr8qxGXwJE557mlBdm8E6/EieB8xq32U
KdP552e5TJMr12E54/r3NbctT4+oqXd+Tz/zJLIusqpEr/aJS/Eqq+ncN+in3Qwd
yYjZCEpGnBqNAAsDyFTrD18L1PF25bKclMHeyBZAwNFJoJo+MHO6dV//Jqe80FEE
kdnHgQjQ7d6AIogaox5pBwO0XvIg2/Bjrp8XD/9nhBjhe3yDttxeZLJisB4SK4d7
JIY/kzU5cWuSs0CyhUQ3NusEN7B5Pe4WFyR7kuYQ0tu3foHOqze/ssFFFde9AgLy
NqBJuysI7aDuGnldMQk73+HzIIzIze0z5SSaZ2W0kS4s9g9FU5ul7s0AUeJhuQIV
A3h3Wfpy994PYOPbtBQkBSsvZGDanyMnne0p9xltTlPG+yOCt3XnJDFnjUpTcmYy
OKxKl0GtfRFb1OX5Jwj+SQkJ4w9VSZpueRnBxEbpQc+MzkpC9z/Yrwex/mcUY2Z9
aJ/1i0RQtJNJBoNUoRUT+/7/0vJve4TGEKOBYU4QCDpsHh7uUtjk8B4ST020BVyD
UFjOiAEWZ5ENvPKjk7f19zAXkbFHF5KJZrWc9LYUksP9Q0+aL8HrkDQ+2BtoHIbg
uERiGCjb1kk1Zg13r8o+5VIZRH/H+4Kttoa0EKr6YKoo2wC9SRQKSf4oLdKpPegh
AkyQcJJ49fgVdpNSHyCSKtfNXxCvd91ATxgv7D/jiH/pPlUvo9XM/ftSBB/u0y8L
t3mIEISk2dDwUZKgoUMeOnFCwkFakkJqjrazfbCJ/geH+DoAQHHFdm9+q5nX2eOa
8f3V6hzdlqLxenUNb4DQgQdoNtAN7swD2DZ8kP21/HLpf0usTq320CWbZKGdQA8R
ZqDnYo1Z1pkuU/dL8Kpc1jkXbjeNuDMjpmz5xujXj8Squpxp1kbPsJkCDGC5jCJF
QuagY3Q00sc9lHtXYwK4DWnRjZ4CnL0W9Nwgs+xXmBgFO57m4Ks6kgFZJKzVwBwa
jOseAYRNzRiuL1n6+63rnlZwGwITPJ3Ys/ZSuSx8UsCLRYGFF+ghHG/515Sr1WHH
99SkMYQDZ/QNTL4DcNqN2lhETmuI0fCmAMVYdVWIpfk6UCxj3R0L/OkjlTrfDUlJ
koTr+XJ8l474IqXC/3JfTy743BR94+zXActj2zxR+owZp8PQ9+Vq4LTmK8s/9Qhf
S8jpKkT1M+/ClfrxMxQzgYUgnvlsalIENRekN8WeiN0ZnJihzCZ88tTSxmWsJLNY
6FD7Zw/d8D/R2pP5jzpsRXWyPDdfg6QJR3Rmd61CmYUgr2ElpHelG9IMvOrWJJtt
xPAH2i0vtcRfpDUGpRmzf+1eDvpTmW7KAEz+3GvGeMlPvRZ1jfgD57EeiL94HuF0
UY9Lu710yyETw3dcQDGKBr00C3HGvwy3xuT/MdDBm9MHLjBgf0Xt46zKzVEdqxIL
/7z7pZLkGX6lWEvtZCw72Jn/2iz6DWfoPCLhMmSJYJeFD9BpwW46WNP1ZVTuQGia
eWY2efYT83DVh14lqA8rf6738tWzN7xShnHIMJAjpvThFv+PDRLnswbv4xyF12oW
RrFFEtarr6gZgwUw6jxGX86wbeg1n2Y1c2JazEjMFoEdRJytNvjmoLSdL3R2FE29
YS8DxDcOYMyWTDGZL0WfjeUbMNCTH/8lBWaIhojA4gjwJSBDuFXuCnXNUwZUvc7D
LQAvWZkxpvvIzuHus2jbF7hwlAkmKS45+nqANgx0NY+gWpukI1clZ/L06M/lIsWG
yGmJHYfVAvvsq5byb+xUxgRt/Q8yNsa5PNPugBe6Q4acJYHJY11VLWlhQFxEI+le
YJOBM2nO616gNLPND0n9bRgeJccTe+skiMeNiUlPkib50fqEU9VhZAh61/7it/wY
KledBrBJcbl34EST6Nk/vcMr9yMff/ja0QJD8yIrSaBKhU01i1m8tOQEa1NE1JGB
hr11DicGB75ROVCZ18QOccgFD2sniQVUyUopLyFhu3uXlCulMifgEeACuSGJxq/9
cTxoaDNVYBlhIMDN+M0p6EVAdN5VsavhAeURsFjS8KE1OOpIEEDU9EhyIUSh2lxt
XwUpwNlgsJoFXTPimOxZpwFIf9mogKe1I2OEYg8mHl1RTnPu3PFAEf7DOrdU0GLS
NEIBu5AcZsbAjqBsgdkaW86cxJGyO+kqu2uJ6NkolS08bQ6GfaLPPvfjsAPAo2o5
4VfMcK3lCyJWkcUOQd9yQ7vXgtbq8jtaGZb4GjvXHXOZdWqy6XJmd/gEsNhG7yjD
Lyl+YAw6BF/MqEgzpVmMZJk3QWVsz4w8MANq9JUhEzm4zhbxLJ5z7HrGmtwYimAH
gHAt++uokR4Qa9yuxIKt4P+0gJMPjIqdrBuZh6fXz3S/1hTLUZPdl65dG77m5gjD
PeYvEzUiMGhPkMSmjprMP3pO16S8GWH2nPiX8v+FMPyL1zIOYTqfFT9quwOzAJVH
iEmn/sKv7oBEcKBfjYx9Bz3entbmv8lTqkGvIF7DBdHIwN1vKX3vFA42O3shgqAg
6yeXCfuHjW/OULsor78yajMf7Vy/PV2YQ7FkQHtlqTLcmlGU3Xn0EGzBouVsY2zS
pnEzSFHb9F90cZFZJzE2ObazLlNGCGnBnSvIi6SLWdT+NUbOMrza5OkSKp51qsbS
hITMwgMnfPCs3d0Xdxfp7jAmDd5qTum4xRcHFuBDH6j1Twquxo7VghFH12kNUPRV
zxAKxVPNV0Sb3ND33W7sSlXAqNAUzAhRGCE3QpHZO4CZ/WnG6c9H26XqwqSA9hlN
Q1taPnLD48aXp5zjHkiZRswrtVdQtwCtuJraQ2Ik9iP0bKYDrxTz+ltFPFAVto0e
AfuI6yK1bFkug+6V23iFmRbWh/vMxxPkr63B/bDYfsbzbML87+vi7j7K/vYjrSkb
H3Vj4KllaeeXamUsxeM2FmUw9Q8lNI7eQyNp3x+3KWpAy+wnO+2icw6UBTVBQz/G
NZD6fzmZRpLf+4hrenjB7CuHBmSu4RxjW03dcMBXpNVKWtHhlw5TjQTdzl+SzYZV
02dbEgN5/dpZ8gKwIGQC8RRsP5rwabIEYgSuL99yLcUhlDsLKqxgFduLHoCsfHqd
j/MEUrJYBH4ZdKTuS1E6ideCIWfysQKcT5//h0xWK7gKXWnVkS8+SAZipoMHc9P0
MPm09O3kv03GPBDy638BxovxPr12GsaFr/ZwJCsnkcMwOBwtcFt24SfFiirkde7N
aAOko6qDgLbaY8rw01e1wGLVe0SYT7f9Wgn0ss0RAlRuXeD4SkFgryut6R1bFMQp
+zkXKnBoncTEs3GZ6jRUOqGy9aOTGq44tIEzUI6hq5yvoi93v7sWb48coM3Y+iFC
T6VGezdZcp6XlPTrhg01K6JWj/ZEcxOrlguMYe5qrXKMMmd6TkmPxgPCA7z8cxqy
Q0jPXCdhPPbgjGcy3J/lqcl1LkPIAA1QgoJ5pAGGRSPhkgv2r8r8qZGfaWtl3Woh
5uT7zoXybpC7MVd9d6+XNmMACiDVmQmKc0aylX6q1UmOkOQgUWo8PAXJDhJjT7RP
fhJPBOUhSwtRmrIQHcLtAx+VlWo6tPionLz6dMwGF2aFOvDMusn4Vh2XkTh63TPf
vNFCynePKKS9YIWkBuHxc05Z9QUzTGsJy92izJWL2EjO79O5ys8fLo8dtj5a/Rdm
u1RY0D1cnbT34MHq8SS3COGwsQc4oqPvTJ37/oTxsRU5aFwMFaJTtWmXS6ZsGMzY
jjl7PShuyhfLZM4T0AhqVDBeUw6IaGYhNGXOxcpYSxfTZ5IunEN/2rtAOFVJdZty
pd7Bpe4VzW36RofNsX0ijMYFBB+nGBaXnyfq26AFxZR6ghJHUjj3jegpsTVBt4rf
aI8sC8h5cwuUZD5ODVneDiI5ESG9M9ExlbUWJUHG1IZOxTAFZHHTKStP41IQySmc
enVoxHBNQPfYJ/DTff7VZvIrTThv+wu1vlxjnfjh4ehJUaW5EJdP1oECQG7nfqcz
h6fVzWVaroW+NerIzBSXfhYQCmyTXPgJH+bPquQXgdTqs5SOQtQKIwyg9SK906mL
XAEr2l2+rTajZylJjiMesJ89w+TIB6ePQBmMyN+6mdVhy1Wo+sq65zzozSRhVW+G
1otLxawQHOGr3JU9Sy5I+KYg6EiFW76hAd4b0iSIszvvzrvLFHL3UZGwNDrzjfI1
xZR8FBqJb2i8rweXzGX0BSfld8p1pcMh/+OKuKAhFPEh4SBGInJST88TA4DrxjGt
msmHGFE5qjEbcG1AwdxY8+4138ldsukwNPpXbTwVhF29o1BAG2oZJgD6XUt6k2Qv
MCugFPyb4R12sVceWKT1EbYmFkzXM+EVHxactHTJ258brdK825r38I3Co6tvkgQw
WSErUeavoAL3cIyU3ulD/8sxeR0yRBVFmQ/TAIxPrnakK6uGEBNKCXQpYcDGwsHx
gBpFbb+hxalwWhpNLGvmP1YYUAEqutWnfU7BdNYRtlBwTg3+xzMRNXb/mfvKvS1y
MiAKrlcBznCAyBLF4+ZZ7xVj+7NLue3OtN34/YTjQaLyQ3rR7ORZt3QjhiBXR8/t
Auq+kKzxXk9QIMLkWtv8hrSJNwe5gktdLguMzdVFqKk+r0YfpRWEIOKyaz6jROq9
xi2ROLnOsTXH5bfwt7IDcqg7ExVYqASgvcgR0vFmoi8/kEniSRvEm13+85W2HJQo
rPC5d1gVNXXK+KPbj+CHGnYl3Qa1uxhT5hsS6DYGr/6prcr2A7iaaEwyTboxM2/g
6v4oF7xP7qWCeCBV73vgzh4gK0PqQmWpHLXTGS690MDM5v6NkS1es/qAE1xIMNdF
69R1ZXbuhmoGfiq+55rxU3otZ7a2RvHH6bvwCKx6PVuyYUdtGlejzFyRbgvtfTkO
XjE7qMqY8GtWUU5ENCmsjFG6T3QHilpSxXR4ts6yasBDUzCkS7HslqEbHPygQTCd
NjFioj+3YU4N7lE3wWm6UgnDp0TLT4PBgsA4Km+/ns0ExlE6XQWfpiCS8zJPB7tW
2yhtTST+TRk07L50xtKd6E3CxLdCSWocseqP9E8XYTzB0Ed45Ei0q9ViHrZikQHI
rUNm4BrTLFN2rpw6WuQBspBSnvhaEiEyHN5uescVXIl075zjpqlJJp1gYdeFL4Lr
pyFGlLcZFEbCCVqzx86azxHQdQHBQ9AjVbCOKbyw4lELTNSNRga8/gRf5GQmpFoj
rzQMHdVKLnQ1hUMMeOLyb0UzDlwE2TG+6iPtPjRtTXTNbvOm+Q8HS4BIdO7DH3Bf
u9nCZYXs4K7Qb6BCirq2IMG7YverjAT3yAdusce0Y/vEq7MOKGegMCgs7O5dLqbF
RHAa1k+jtf0vZUoydl8y4ncqOUjltES9hsYj3bq/8ZgHaRFogyjh+j3UTs1cCatt
GWry5kafnWO9Saw+VOgomU750G3NdlptmIoxAPPk8B9uombsXz4IojFC0/TJ2dPI
4oMGl+K53XsScoNm2++pN/vFTZ938EF35pHx87X0k0lLxhDzF1d37MxfHUVoTguQ
GHmau+CI0Ys7ucwbOehvKZcaVykj79q29HcGax58yUVyY4W9aPNHwti7oY2SrYK9
1LkXXUi7cCaYqc8v2ZftDvq5rK38qOsBPhV1sIBS0lMyTm/mB1fDOA9ykOE8S0d+
z6jjAKFTbf0Lb67mkY4FZrMlAqx4ZtlAfv/8tGetXhRKDYj5QxRihTsjKPDhZdbw
9zrE1cf8UC/MeplchjDjs2vAjzHcFBMOzpUA4Ix3GKKP4870komf7JaiAolIFk6z
0UCqrKmvXGmCjnT3yAnYcKvfwxaQhlh7X4aF4699nukj7Ao8ilnOYD2ZDV46KeTu
y7iFjzC15dkR58wdRhTKsG+h4ZttwMchJRB5/yA4P1cXb9i3UY38mD4uEqiKsA3A
ZiB/jgL4Gkx+A4nhE8PtN2XVVhH6F0y0fb1uKfVSY4IICN6BIo11vKwdT7Jw5FFf
RDdO8L2scaKEi1k/iIrE8V7UfQPw29V+GBIGtphqKWVFO7fvtsIF1vGy7sH9H2vo
jRUFs10PRxKDMtLWs2/kQObplS6g7Gl4tYiXeycxDZcmTwkvwRksBCqDKncl5Z3c
/fhwKyWjGOgWrY3jq6v/0/J8Gr1GdhtL5fkyiyXQuJSZVJOx/UGAvEvb7OTueyyD
/7fswfvka1UjcpJSYOSwy+8hvctWqI9NGL4sv+rWoo1e+07TIS2whHIJMtozFR0B
f+I8BaKzLwohgUFknSfI+EfewxwRHZ5LKL+w+yp/KbLDulgpckYT21un9BXTIk3i
qj06nzOWZw0tqSPXh/hoyTuC/GCYDy4rvAaAVflj8fvM1sJ1+DMWTUqpcTBbFA+4
4flBWrRybATHHdgfJ1lahkHvnChNnP9DcznoukDQDge8+kj6NyyarVTx7hm+9u9e
J2+D5/OQyYuUnt644LdPfmyt68Eao4K2DvaJExDmroUr7/K4ftCpteDPhAf8NIjZ
zFp5c54/t1w4Q4MaBDeJhEcsnY1GZ1vOMoEs0kx6B27x8GQLBJp6CK3NNC2Cl2Tb
cAthqXIiYnDQtrc5pjIkpK7KSmoLFNePBrZYghU0sQw0BZAj/+JT/1daIJ+32qUg
Uw97EH9BckYfuXeJVkyz7TDkm8l3NlCYUiMhvJjPdls6CMkp8veAJQcCM+WYC6nK
IBEBe2nfCHUSeulP1zAJ+p8f8jQhnufGywQ9w/fjYrR3aWwWYAypNg7wuLf+96ZC
ZDGaO0EWw/KUV0/oi75rGEeQ3gQWin7BijFzp9kAslnzSCnAhZuh5KOUJ+/J+UgW
N1kKVxK0lrZV67UV8eJ+4XDM+QQJomd+sEmxEZKbF+Cs5oNTrDpDecWulLup5Q7c
txKw9T2KtnPsIxCNzp7VCg44vRKozUISu94D25PXyndgpCTQgBKdyNILrcFzRk+U
1GyCjZav86rcqXhd6/O7jNCIbF5j3lxeHd6pYrcPM12AQkKIC4sZqpu3e+6gP0Ii
fhXqYvmYQx82hUBULRbjTcmIgTkBBW6Gh8mflRJhd+SGzVDKSJ8mTOxXzVxp7nBP
swD2QdIhuA5xX6CmqWY8g3s8k9oU/unQQWldt65N3160UxAwTNJIU+NORoWfg4wG
1m/obO8w1xrV5in7aCxTF0YZdMBb6DQw3yoPD1Sh41La2ybJ4/LRjZqDPWNlTL5p
P8TGBA7CDjUp/IpEwZ03Tca423BLc98/2IRoQXUT6OjMFdulmRT4B7ge8p8d1nqs
bN/0DGANQN5WCaR9cHRPwFwC8NlnQAxl2/lSr8gSDdrAaDqNc4iK6+G6OUVymn+G
d9FnLhETRFXE4EoEPHlTTVQLLNUtorUgxfHyO+wN29kHT6dFpZbXdXZ37L0B0/Al
lxcqu0gj7aOby5uq6vLzQ0lZfT1mm0y1+RWHVmbG3uRmtmD3R+RywiXQTalSSlpy
S8EJwHDiS0rbBekzXyMHwUUA+emNhYYySpSsFgHlvD0eHMp9TT3o7OQrmforDi9U
QYWp6BFYbtbDZKkxFotE3oE7w84gzQagTmCjG4uYxexB3Tr401A+oxCkPJWCJoqa
7jpx9Lb3VFL9EoBEYXnbyxwwyiQQiSbifV1LURnc2C55jhVqHMspcjPGeFI6Z91f
tUQG7Ck+bdQqy227037r6pTLSqWen8LLr+xBtW/wd5q+XJYf+wgW71O70JrzSgO0
y3s8DWWdRmcWYkSthdz9fWciVTxdC/zNS0yv1+B8wC+81mKb4k54LStx8IzYUWdc
QBu/QNNam3+q0ASHrdE78oNwFUtljpQCDGG1Aq8bb3zBc4Heaty1v8c6LjJmURaR
vwZMOJnareJOkWZgT3TIeCqGJzHSk9kAS5O06QqVpyMa0qp4KP31isGdZgrv1ixh
X5pXiVJZ3i1TEFM3J8975W1icQT75wNB2D+vas/HEg0Q/vRmNwrSDi9KZsfLE4fX
vty79l9wq7V9SxM5BLWnVD3ocLrQyqeGd+ick7jYCeoX0nw402g46CnsEqXtKwQo
nV07HztsjKF/to8iZvmEQuzvjsV1LmySY2hLd0CFPDogRZ5MVJIaMKk11faplm77
632HwhnsXZCb55k7dn39akq/TlNB+dL1dOAVRivXHD3yTFaW2Fy8jbSlvEKIEKti
rC8e2DtPEBkBn+Ef5IFjNTXSErQ0GVjTRU26Q5XtytWPVB1atNYbkzGUxsDJa5+e
gyU77UrxRvmEXDQUirSHDbo2tGG+fXt6FDslTU2FAjqPzsLm7fjo5rwY8oFSK7k0
8PDjeH96f3IdXEtCwIflUKYEOOwNtRd0u00LMLe6GwjiYWsDRZ45UBzxj4EDvHlP
05W4qa41r+etTHh0nLnI5v5plfvEsOQXLm20hPr4HhMRtPi14rY7zB/l9CFfkzGH
m454EkD/jld6TyNMI5OnyYafts/fahv6dDt4bJkn5jqIvIG2yav/opk+gi6BAlE4
SBgkg4HEec0zHNQAQpqRdsFWWtx2e1LnmmwAoRLZUUIoVw6UdrMsruH/+avAgyzo
yY5OMefpJG3SRhroAJIhIFLfRShX+WMhnnogoYE2A2/2q55krmOuyUVOpX526zxt
abdb1kD9/HVY0Bvh/J0TTonSsleWLN4qk4zhE5+8n3lNMuruBNSet1zMoNxjC7yY
RkNi+ywcAhSKiMmHi7BiQazwTvQCK7dvtu0juRxzZfvQDTwYHFZPYZ7ahfA88TW3
aXadyncfii3fx7o9lJ45unacoZGHKI3pASsd7jTRgqL0q6AX8Wweym2gsxXrI4/a
k2T3VJcxeZPVAbu87wJXRsHyb+QHGhUM2fR2ZAdRnHSr++4jXTZqa+8Mnt+fBbHk
+ZoLEzuJb9hOgpEIzADQ7iVE94Z89/ngsB06QjzrnVOFpdeVrH1U/i8rwc9GBx5F
vfFUrIdbtKEO99Exmo7s2qYnyNiJLyVj3A+mm/4qG+zu58ec1FY8rm4xqIbN7iLg
PWtV/iEdiDD9L2aB0V1unbg+0VMn0Zs+rnieji/3VcCYOS0UjP3q+/Edg6xwMdLU
/cnagz1UMRcurMn4hJgR9isCMDp88IK9lMlVbqw6dJWbBZZoFAkCVq/olbEHVYME
CmSexf3m0FoADjwQYFXzWMBM1JXx0bjkiGwcAtP0CYOmmp8e9KpBlHBs4zUOcfjt
W3Uj2syVydOKAbgoFkcmfd/6XV0R9s/dh9trXmtHo4viLqvAnhbHjPU5O1KUoQfa
EoKCw0HgWrOfy9r/HrEMxDO5qWxIHdoTfdHvIj07BVoKBl/IL4jteBo4jf+HKi7A
pJhlgyHt+g77roQi5GSFPYoMeVWAESysA0rs+iOu54BL5lUdSi0msk1wS4YLBJoM
vuUMH+ZskRu98zdbk1zdchqCpubyBq9LGnNNPJ4tWGpDpHZ9W2HAR5jI7lYntrPa
RTDTP/G24sG4siP+GI0mq5P799FQ4VZ5457KZF6fkV8YFa9zpb4eEcBZkUPhARhH
SNyV+jW2hIX7o2PAwJ5t5oZjj1CnMSw6P601S6/5kHM6t9D43+SGS0uGEeB+C1pW
uIEXCgTHhBpAP/kGiT6a+1f0hs090G7+2S+1SDwbwPB92wl+3jN9vNf5f08Q718C
8O/XGNitv3MrqAjH+GuqVmvDvfLvEqFVMymLl+p92sxAanK674CzTl+zqPXjUudA
qT721c8cVUwBFuev2HJCyvsmPcCz9vOKCX9ieoEg0/HJzCe22/eA4ZUwt5UIGgXj
7RRLsBY1ueQp2aAavpbI4KZplZskxrHb4X/vBJhEHawfddt9zDJN4DcgRNkee86x
3Gcyz+txrjgPAIeAygzdmuAYDVvguJ+/JoomcqXp+HHpEzHtb/vKH1IqNg36Qgi/
/S1JMpNl0RYO2XS7DV47yT+du7rXzMxUyUY5x9/SZGA2CO5c50FLbpwivMwdyh27
Y2Pkvyk4uUA+O8BMW+1nrHkYftjU89x7rYFFNO558KvBk9TeCzs+h4nnFUBaq509
hAwPwaBc3o1YGWbG+O7eorxgkEKbholI6dWfdDv7pmKH3LdUBLsmCEk0mHqnNjL5
yHlqpShVzu/rsCpNt/JWj8u5Rv2tvFIzDINAyIZcE8Ko2j4wqXXdpQqGGsRGi7tL
p0ZAcFJuBREXMcf4Kv1CpzOmD9Z/GQeby0vI0XPiHIzYkamf1UVpEktguqYVH+xK
HDm3+8HjBq8FuNf7i+UJg/kHWj37gibtBQP5fLrglnf9VQkXRvrEBoDtkkBv4mje
/ueo2qgb+YyRCPeqbYUSV4Bz9Xyf5vCmm8taMFSoZGjkm/Q5lodjkvER17ODB87u
JisyLLg/iE9mIpMLqy85LqRZnqLJIQi25b1LqzUAZ0LKRLELOR2OlousGZRKkDtL
i3STaOq/xgKX2ADGRRd7e4FvjCQK+Olo3qdK2zUew5srCoBwVMf4a1JdMOtDYAkm
5sm0bbfp+huB4G21X56F+IyuTfNfHD969vdaP9efCKtDxBzdRt0I/xz/Os4bUrzi
BltESpaL0pOu2T1q75eCtI9Z0mBJ3Y2JoQPT5p64Ge/yIJvp6X0xds3UXUx0z5mT
oJfflwcZRXFvht34y/dvyvO4OqHHHwdx9rctP7VU/vx7tMnBCKt4UnIbrIohZFt0
iGHxzYc4VZH+7IJwcMDuCLr7PpJ9oN/K+4C1g2avXAb8ySixupR6nCCz1SGgEEmu
iXxAxyKZd3GDCNdqyEZMDnraHOQn4tZxnf52ykIrlt4jELHoB6ek0oT+jXoB5Y5G
v5ZtHqjpcjeOQfA1iDUqgGl372AOUuL09q2CO0Wc8HmTY04pMKyg0hTPsRPZ5yZ6
2175JLGrDQMyBQuh7Ktu5sRwGn3JKtWKcmj+6TclBLSptcnk8abbzPrnGk+2Zwpa
KO1phEkRkntw3IJw3m18RWJvKe/8pS9eBRzzXAOfYOrtIBv9/jP+9aocP4Y+4OTz
V1692JzB+6CIz6QWGHWff1LN/6dvUyWAq2ZtL5oiKkCtminm+cVKOrPRPJ8C/hm9
p7W3TDK7Ya7UaYRxSDFnGIRurz7K16njaXfwcBD4pB2QWW8DsjrI9ZQekqWclnXl
vN6LY/G/tLnSQPY6eAlxPLRhM9HNG9H8SqAM6Lr6cevrqHA86wSPzOd4L9izMMd0
EZOZIncLYBu2Y45fL7Z8ijTMhZWtk7CbRSiVj3hcTvw8bcP8aARgZtvzrygWqpln
MMBPpCfPo0aZ1pwk174BloXGVJTJrBLGJvmsrF8womuuX87dr0cSfPUEFVHs7TJA
668Cz+/LoejvxjeA7gFoTFjfVVZJBglkrbzzQf6SVw1aNgDFVydUQ2p+RgXVW5LC
jNG3AkEpSz9w6F4U8tyhBM1zTlTNg2qZkh0ObI9/kge06Iq5nO9y9l43ko8Xronn
wmE/ViDVKOcGcRFTJUP8e8B5fwu0HGUBHBH5O4NPlHmQ6wTfrY5kn2ctQq3DDPl6
KPHj8EsmqwB94pCwW1Y7aWyIPGY70utrtVDypDXvJ8H/wqKQxBBwKsKxD3G7kSiM
IclB1Da+1ZM1r99pLT9m3v+DDPHDRwMrLK7jWp4ElENSE+nNDxsPHbO4MYq3E9Oq
EAypRFy/pWVwtCF6Kwc/uXP+1a8EqAq45jyzKWEhKj3Q+IdKXJk0ub66NSLesJGt
SF5t1LeT5vuvZsoAzBlUYn0JmuFkuRN/o2b6u9f694lRz/8s/hxdsQruiHtqx1QL
EDJ8uXYHFy7+I3iUqnE7DZrmJA9BjzkoiCqAUAd5uFTE6aRXfDxLkHP+bE3WD5i2
5lmJPYrMrVMyadJzBVv6zqIULJ5jWVSL6EUhDOlEnx5K671XkQt+vHkXWVfMqFvy
VKTYtEePa7XO107anofaNWnBz2hNaO9DyfttAjaGNit7uci2AIFI2wJEMSUx4Ufd
UkfhbwSjORhsOkEh1GWgvbNmwtG14dA3pyEiw3EsRAlgoRcp/1zAF/Q9etRn3M0p
/GPvgyNunrufSoaEcw2m2uxxPvqmm8vOeGLUzRHymSxq+Iw5i5vAyZ/fZ0uFNWth
M75Hh3UzygxVXKhFxnqt5Ty8ZKgMyrj2bY5SRvtRxzahFejE8ugJNyRrf/mMVnOG
WoKmJT2rZmp5RFr4Z2RYGgubnYJa+UvmIZW2CZUnoniilpJIJobcXOFy/2sfFEys
GYjaHh3OTTJZjRpsqWKc5ujrECHm3HUsLnAurXLhK4pqjA3uqiyf1TJRO/8M6p05
pCCQOD7PXx+hNyX3Xo5JD/kE/BOe6qRMagOStwt3bRvaYVSY0HVuYYDuSIyEpZpw
ituAPvAHnesI/B3H5lkihRztT5kSQIxuny1mSHQsBvbQztAGIIsflNNqPyDcv/1e
M40BhyqWGAFgTu6xIyk/3BzyKW4UJhbeq8G7RzM2EvBT+Vo2EhMBf9q+KrMHacuB
XnFti8L+wTRCGl0xmmQc15CXNjH3yV22ij4Vg+04jbEkfE/y19XHruAsnmn/dsAv
vR4tqmNUN7x5o0TsfsAaZ2tA2/ulfDUoY3Ats2QR2r/ASLXcSCIiCi6cd2nHLMs7
39+CAABrq90o6YiyF/aQT4Vmwiv0tBN9yTYGjd542WxaVdzIHh65MSmjv+tBEQyC
2Zg64CKkQVqijbL68fD1dbnlE9PUDV2ZZ+FpQYLOw2GNdy7NGPwRq7qPmBTomzi4
pauZmdEiu2pNMZJx1vWQBC0wKiPfU6MKRUk1Y3jvpmyEZagRMexQz2anEYoJG13Y
vh2OQI3OnbzxYmMXfFDvlwhVyoxWEZJpl8sbZUFWxKSSiIEpiDYtYjldKIma5C0C
xDR7SG36Anjs3b5BKoX8DlYHx8sO351YDTddCxJ0LbuPY2E7u6WQA+MIRH4pJBGz
1uoKpjTZ/GT79tTypt2Rh/oR5DDmR+sJbai5PwCyEM5lOr1oQ61R8m8xBnOYch5G
9KUnc1PSfmD5XLCaVYvcSw1nvX68a4fyymWgphk3WBZdPrCwQVAla55NYeifJTec
Lwx51xYSkKu8gujf2slRK7zciH0TGMV1PM/5N4/AjGVFqwTCzM7SczbUohVW57Xh
ragAv1c1BCXRQxsnJtrlWUBkwzhAz8di47TQOcUf+nU0PVU/9eO+ZiuxzI0zsTzK
EQpuv73ItF1/Qc9FzGqUMntiOu2ZGwwBPcLghs086+qIgg7WDsoP/hq7N0dbnz+t
scKt4PPtKKZ2YdqnymRzmD5L1xMQFoiNFFbajKHqINesbnvm3OCR3XnTjAsQDm0x
qubpxlsKtJt5o0iexZ7aRR5AqZQbEnMjREA/xO6rZVEcAWvYIJim9fSbupjD7xwm
UeLMNd8YsuL9v36359rTavCl82tfcWP66OguvXGpCr+oXztBSeR+U/2QxPSDJB0s
gfRJbA+MfqNA2aitvE0ejSnikvOiEWu8XgkUTDO4RaDFzX1uSLXgx3Brdu8izHfO
VlONar+SvgxVF4jr5gPcHJMFcR+2q6L4Lx2+YTCC+EnTFSn0S3ZUz+fdr0Z3KI/2
d4qSsVL2MbC4wG0LnMTxoBoP+rOmEPv/5SoPXb8iHaTGOKtfKYOPiJWie8l7rdWt
IFjBeSVEFeLENwgBf6UYN4GP8COT1vMKyi6otIBQto/tUm8U5F2x5woQjCeC6+j7
5S1eJPT/JfvLHkx1y55kDSlKBKUWekqBKbFq+zTc+R/l5WOmapl5lfHV/jRmsUvA
3PpawhZYvHqTXXsRlyrtC7jvEgvvRItAYcIL7EhFB6BVbXDrADpBlFV11IJIYRhH
TQL5VqnDgfFVsV4/4fjVbCn6kBplIXMi2x8A22/6LGqpqIMJottEauK3fHmoPSkP
Xff3mfOfVxUtYmFV29VWN8WPFM9wEIH3qTjgWXBDEo+KRKLi30QKd9KAR25Bg2eh
Tr4YneiDmPjoWdk+E5qnxBY1HKJUd+xOzH5BoLwqxqccUxb5MjoXUB+xTMglxbjv
nqAmvtf6F7ZjjFqQSPV6O9ExrtsBEy/EO//gRHHYhfqmbp0Uc+lUVVMj/BQ+ORVf
E0cOKJUIGa2Lt3cvHbTxxWlfFP0iatSkjmYokmA6Pb6xsosumbFuju11E+sCnbNB
8qutp9xu+UxBIatmTBF3E/G9C4B+/GFtb21G9OKrhtkoBRg8DwYg3KLsrjp67rPm
q9bgXnPTMIfMDyMvizi2eBl81GY18XEJd+c6iOU3dLIJDBFXJegjAJsY+bevniFq
F6HwUbr+vvHM1cNUrQg1wCiG87cxWr4UwonClkt87cvikuLQA0KeqeOvivJsB5z2
Km0nju8DnlL1hbrYFalfDjqVtZc4OHarWOEwr+MJzMe2+nXlNLdTLrfRyplngXAd
+T0cj3/Lfmdq5ua71xZetvDOagoIpm5oK8rFPC/E12phN/LV+FIJM127MnGFr7d5
PhJDAig8jI45gFNwpZ3pHYHuxkoMMTvf4RgkI2oJJMSHFGpe81XZvPpBl8sHU7hR
z/WG3Tl42WSzbFLR+QL26nym2eiBfxQbuj2kNGHiJxqixcRF3QX1Lb5XVi/ALwvp
B/Ba30wjMH9B7E7zhuyARkaLRoyd9zpo3mfBdj9AfEOfyk0ksDGpwdDcPBV3JgXy
mCkpO0NdtlbtwMo9MvcnFnLcVbHu4JHQOJ+FR/t6WvX5R1oPREFkMuG3NAycCBCK
eERPmyxVCcYm4rQ3XWtwcW0LdGTGwpjB/UFNABijmMH+w5fe5lau9a7r9zgl+60r
HcQpunT+jJt9Y+J41OEFN3y4x5nR7FGD67D6za7Xc7W3/5tXJ1HaZn3uNOqel6X2
zAPMyHu7JRrGdk7AbrE5n7kqYBd0bKGGFJ4UjZ8+gN62zWXK+L7o2GPyijtgUl3l
lHbA7lm7zIgfFUNhE/hMyU0/olbcD0HrnBuT/DyB1AdRf4Og/9elDFrCVYH+RtN0
QqDJSmDjzcvPsUqGECKZl59hqIkrk5ZvyqMXKmyYdhpcZEdBEL6gtheoHxjgHskM
ldOJphvSWaSOreMwRzeZyI435GQ604tv7oeO6gplACYdZCU3+k3K8Ron6IQL1OeP
2BELTvXXSv9cgeE859MgkYXBFqgz9/4M+tHd517YbM+yjedAZvFGSvE2x0Kb5HIj
emX1Qjrp4xjVx7g8hERuZ40+JERwUzq/0ThqtXEWJgoJT9CV4Ryx4SsfN+UtJ5w9
0QbeNUg1XdUMocR81WzexeQD59erybO5rAgmG0/AyrRqg6ObgeT5kWaPSuZ9d5Dq
YpnhQYC4B7QNZ+dFJ9VU2oCbhrHbEvNrFDaB4g+6CABRz2aOGGr5Wa3yM/faf8Wf
QDxdWM6EyespEK/Cnby3YFPux78aJtssINt1SSQzKp4WdyQuuHSTjcB+v2pGyN92
S1njx+Zs+7ImJ8nEigJNnX6eefwQB4Uk+XEiUdD8FKU/v9uIaAe5dbs4LtA0S8Vf
uTNV0wLdWeEeZbxjJS5UzajdAn6hePJIGhuY41fVi2IoC2/F5R8t8y+miqNpUo7K
nR0u70hLjfRjSeYHGtdwlmVO+MgOElf7GnouMlBQF2xX/uwz4R4gLK/nMlebTBDa
xcd5XlrGmDGfAeQEDTHCDlhAQSYgKpB3P1+Lo6ZDhy5jfIyphYJ56jKZ4kMHEE0e
szkhrX29+V2AroNCxjvUHuoLO7img4zdOqK5PBqGzkOupnX5SNdOOCc01uHT8aYH
m40132pWUZ/7lFE5hkR+7sZFj06Bysc7ehFAozJeIUAS+TyOG8vAAYTiqtMEHMBC
KlKSVz96k5KBtGQusNvzOe8zygA55x8sNqolLnDPzy2ZSw/Osq/58APF86D/ozYl
is8U4vaOcmjNH7Yy3bWL2CG79XZwkOs2qIA4WUJ6s+oob0pvAJQEYzTNRVjZklTm
V+TAgQao+YxBhHzURMaXdK/zgBl6CMKJVAcp1DYNT9aGCbUOFDj3v6dpSzmDYJxi
4OVB4yUFsf1XewypMA6HjbJndL0FIt71Yruj0d1rz5QPf421vZEVyOBRfMIdctj/
HPWWvHJoixhu1IxAzJqSPitKGkgHr1JJY7FHFhLsMMLFcPQQPBrwYrqGaLXOtbrT
WckXhLmC5CLcJAyJgdK0EEPKoz2XrPo2SZGlpH/gXGVRSUdufg72tyuVlQeQ5ZcK
XwKDuVg97y3yDQzWYv4EbXQ0q0kMah9oov9ROkwXV6AZJJmvrHQXi3vq4q6H8kwz
PHhGFWY3PvbPNwD6iHybqAmUVl3UfT+n7nMyPPuPD1+yvKwceQEX4AB0/Pdp/QsV
VA8CNb+4p3DwzMOEOjDveCCr/1T4CIVde5ivjJWqHSnN8DhB8o9TyFTtl1nbyGlk
u31DUDLy1yNzobQToNnrOk90bdMUYluww3r6JYqSEQYjqjzpzg/UEtEMqG16SasV
VZC/CSAmJmeUZhyFD/jD6cW+zzT/jVZVtgakjFqghjEDoW9Ot0Z8PI+tRoehwMBX
lYdf/BI9AbixXk8FDy5+10zxiRQvtT08vowCj1XfAU5RBlYLqLZ0rMbaaciOYFB6
lL9d/WGGvv05KozkK3Z2soxtBEvGNE/cbcgoq6ARRJguO8b6fEoA3BeO4xtiWc0F
Yxn7HGwRv///+1vAJqr5u4+Bwy7usiBisnzKaZXTxhWvWZj3SSeOWX7ToedYQxOF
aNyYaopjoH01kA/55LMMOi9x6X9EsHb3SgCnEHK2IYnKE5gZiSOByMILFe434Hmp
DAIdOVz0vAt6aVKsjloVX9hmADII/P5aI4rnydidFNhn2AiqwSENxaSbkL8WXR0k
Y1/aBYhq5rzxjCwIy48UD6urISfdtTRbQIqquBLq2crhsSLnCq0oAJCvrPnPWrzP
zKfh7ZJGDxQgFGQnWTTZy4ZrN+z6dsGzqyvE1AYgGcfSi1V+VmmKxqpPgnH/sbnT
j1WoFR1uo9ljTv3k87GrjQiom6f8bboWQS6zsXKSXsh2t/cq0MbhpY0VRCcKPl47
LDoEaTw2xE+kM3dxWawKanMD7DwDtDzWATIHEXj/n+jfkje0YFonb41tuuDowzO+
M5PJ9VNK/2qcaEqknrXpqW1B1kegv4zsSr7Z4bl5dp/TVMi3RfXgydCJXWZlKtu8
w58BOgQA8myutDJGlNH/aKe4Q0ceXX1pNTCoJsBlCi+LAzuY+m5OHwSD2IF0D5L3
JAD70zptpq5rJ9fbfkfIuJsIJUkbJXsY/ERU+/kb4FLnCCawrJDzipsPOqJtlDy7
jm3yRF4RJWdZv+JWQ9N+MXcR94IfTRSh47mPGUXae8p5i7ptCok/N5MtIR/nk8w+
oBbLezmtMk3vAXIAf2uEkME/Tzlb+gtZZuYa3SRoaPpG1+rT4zDFYekExCJNhc7l
47cqEjcgJMyE9f35Dg2pt3awMJ9f8pl9Pp5J3jS4N7A9KMqBiTr2g5Kq/rXabB2d
AGMocmpqBFF9o/J8y0iLFgpQrlfrxkbL5LwRS8lgivvuPDUhjQX9St49BRM3FL9r
DXodgXe4yKbLX579f8fkJ43vPIj7sjYFMCWXVSBNXoO1NvRglCWyW3eJurrEj3Vs
CX9DcDtFylZwoRHoaE1GtjUbY9EO9HL/VsYTSzcputnsdFcduJ9WtEK7g9byHHmr
8FQYwTMxfeRLnUsxmF3DxBGo4cLppwsqL+SpBF3VoQiNNE68zDPVHFduIw7iaSoY
t4SCA+/Mj54Q/6zoz2CbScKkbNyjQDbIaNgjhUnRwmSGnXloqW/4qQWGUsYJ0CIy
M75GDrR8BNbEeMiWj2v7JrIw1X5fHucgdvARRwFrGoNj7SX1fkTvD+qNU22x6VCF
QmcCDeFwV6rWQcggnpjMs/16PIg3SvBOzUZPBASrOwcWt0MXlTmR+hScWEJeGrsL
6RndnPgzBhnUdsM8cajL/VTwmfEJ0npH3vUiXS7OMeJmFD5WRR1oNygMXjAdVUf8
PYxguxAhykPWooFZolWe3Uc4pa0YCrJiRZQy0LoLesZsWY716QoXfsWUqXdijTMK
PifiA0TJfoNea27iq/bcH/ScZbvG0UKu1WhCwUVPCLnjzINyOWtYFaN6XMmRa6o3
VuyBILvRULu/tjER0oM+6fVLWgLej/yx4deNes2HfeBjM2Q1HPadUlLf6MVUmhhm
rgSiNsKwxMD37tLoAqMiqHUIgN4Vc7rDTifKKS+9A6jpfxDyFLWRAXNw/d1O58kF
x5eKMezMK+xoZ/Ydi/lejCESoB9Ib1URGOMBvp4w/o3X3kqMFAHfGZjMbfRRPPO5
+I5UKRJjVRqysnqLQiagUopjznfwLDIBGKuqzDsIvLK9RNfOojPQc9oCpVahkQOf
UH+zmf5zhSjPHNGFv7dJG5pwZSiZ30zETWIumFT+X0Iwgmq+/QcyuGgwQF4XXM8d
eaTUmN3gNjocr2hwdwENn4Vjor6ENxk92CpYfxO70OkNqc110swoUWhYA2/uikz4
2zsDIwIjdr7YZbRWcBuM9k1WfxZwl6kWt4l4X+CRMccxOXiwXkvDtw/PmjaX+BQX
/D3QHXuV2iYi/WcVJPTifl7Iua0bO6vZ6LC4kOe9yH4p1w+chS5Aspf9l+to7bba
hTkzDkUDbiRNipXl+PwszmdF3kf8svZV1IvUMfxN/sc5mCVd2segkTZgHhQPRm3e
Ni5dBvK+H6mITu7nzM4+tKnc6rvV6PTXOyXrX4FLnsgDlIqWB13vJ1v8XVKQeKXY
UVL4BXteyZWBd8tHk8+00RNpPdbOYdRsik/A0rS1XC9GKGmkA/WXwkkAhbDvkz3E
wZcAfXeZVol9HdtFsDhgf9pW7l2iRFVPqJTwGtRQjmWrHGl0/kzQAx7ibZXkWbcO
sTb3wFYR+HjIQ80J912MIWwcu6JcPuLQTtiyd5EKFBL/DDxZBD71MYtDme2H+Ywo
Uv7txFyRAB8DcKQl5bxqzLogUnk1lwtpRrSBtkHtloG5lR3oSXAm0iX25gNGXadh
p0uNKO6btvGEikyp5Aeyav6NAHrfalBhmsSSdh01hWEVCi3myoT1gvXEigixt1I9
0lQMNoPTqBcbiDiQek5IoZpjmgxqheeIViiF8iiFbeljGT+WH2wAl6Gp0sAT56jI
A/i17w0xU34m7vZJS4FwRz31CdJkMSwdxqyrb20vdvZLU+NUjY0/VwObtCH8wOqd
9kaNShZn+o5Ea5oCnx9SOXcpOXPdoHZhUJv7uqZgjmWBReThhcRISBvJb78/YIzT
X1JVgKV6A51dgaucaXegiAsHOgGbgZDLr8J9/pzXPNMW3k5SmKxC2r17ZDLsMH+x
tHUbXJHOUjaMITasLetVLOoZXVwYYm8ArJlO1vgYlE8Ewo15sEVY086hjOZTb0/W
zUDG/hcdkQ3CFK9Fhh8juCgD6MvfiVw6nXik0vfvdyegKPmEZx1ho60ul2lkDm6r
RoUhufTxsLqp2swoBKKpO/qeWUTjLXpRwS2+DQbxa0zCfRe7XLi1xhB27Fx49HT6
7Bm4i2kfOSeeFLYtgnKtGlrNQ4QLEgk1j08OobmjFkOD1lw58/FCkDWSmKePbVks
/DrlfPszvWWsX8bo5WeyrQxGYrkEW2Khz6LETAuFcwNhW4VQie2FCTt+K7Veh7Uy
rquO6JmQKqoEkHlFI2zZ/h452hh5JqGGQv7aIDDkWwY4873OLmqLFfpUnBOIu+O1
7Mv0UN6CU8pOGSzX8Y85txW/kR8xoZsa+0rvEih6g763v1skSxfkCyTtE0c1U0Mj
DztC9+Jwa1O84ij8aYnGZ0A1zCo9yrye5rY6vmzTsVycJPPFKVxHu0Wxwn65po/R
vl8Ujt0CYqOK4YZ4IvxAWzo6Guso0Pisp4zELjivI6Wk5fXGO35Rf3qT4otdhgOq
FZxDYGX6G425u7jbfvaOwzsh/RhecMHFuOr027rvStOM/S4SGwz8Y14+AV3INEMh
FpasRJT/WYT24Gqa4b1FVcnIxmpqL7AeowPaF6OC1FMz2DHzxhICVvDYs5KwNQ2p
bM69M7U/3M24elCoT3N8G1AH5WeBP3IX8oKo//W08eQSkDOeR9Ok+jpZPn9KXAKL
E3OwNJ0+9TpAVz69p24ar+n70YDMuGcxf3CdlqjlHvt/n0lajDZbKjcuEh30EBrP
jsC9ycIHetpCtcryh+57CHF7OXcnjQeRkyXvgDPi8bqftLYTftGeYP8Jrapq6wGB
URMQnCygFLjfu/yX1jzRMnS2UklqA/7DymlXEJqIe2FEj5L1HEVPhPVj8PU21BIw
BN68VkfI8+vhxPPrAIZXHMsQAeKkWO0PLu1TUQLrBWR0d/TigKXD4IS8vySDCpGf
2qoRrFDeTmtVF38bhTixde327JbgCe8LXkc/7hRL/9j2xbuXRZCFHtmoohCIpDjL
IuKn3ZFwNQj3wEOdmNSZJct6FCyxSaMt0y4GSBLholvXg8dSqBCRbyul7h1bBgDp
GlGLuFaqSDYaTwXjfqpqC9PGmwE8gA6J8/KwNcvEx3Y5jCv4k9VKkakeUrH20cBn
U38NO7My1MXoIt4JuJOnAiSDZ0jAaEwXdUspU7wtfu3kkvTNz/t+I9vp0mfZPGFO
Vwjva74hpe+JTtR7zFUh5ustH8bdTOFndjAnZ3fvF5Cztw3Pj+y/sdTieGQ5uF6+
lSTjmDCPV3zBeF/h1hO1PWT3rTl/L5CBEzRD3pZ1FeajwVchyvKDyp2in8YkI0W2
OZq0GjCbcyty+wzqFLFDrGjPZN3H9Xx+iWRcCV5pbDlUw6dJ+ZaTDrI0Iuc1pS4v
6LeKiqBGIOuSRobNVRM+oM+ZiX4PTUw8zY0TxwGT+baoShdCdu+/aS3x90FFuJ1/
TwgsRgx6K24I5/TqdV9Bocvo1FARoiJI34VPELMdz/sAi/BmObzmuqVZMibK/V7c
qWK50ZWZKnVRaEH+/QJ0o72rJkfAKVDO5fnxW2j1nI+7yyP4LTeQlqim73FmGllN
iPv0Tx4wJkVvQ2Q9W0OTXdYC68ZtPIjT2mAYNcKRGvEMcK+T9q//tryKJQ8yFonp
5tlaHbJL+eTsNwAZnhhW3aGHhE0aeugwr3eihR+8jtXTT+B/LKJc668nqJtJEzqj
UxGMEPaRT2evNKgW1brcI1d1tkbwrqsFt1g+e9Zz9HNMPSEXJV3FmGDy0/8cKWVM
NqSS9Oy8ebdxNWW26GQZ4RK5NGStIMmfkDzobXtEI9TId8kWtLvgLPVWj2gSIeak
aeECrri52TpccIr9D13egVipoIUAZ9fkCXOyP6oqN+kOadbSASWRvpGc88wslaXi
kN9tylcV52pK6RRfLbnt0QpkCIeFD6QVeCjZUXykdirYgK7VLR70T0HIi0X1XJ2p
6L4q50JtQFjNNc0LB97u/jctSjQ3G3NUb5xXS67NIMjKcdYpPLl3L5srNKIZPfZi
Fk5SUM7QkyakbiZD0dCAqDIloifcdpBDYGubPNT/I0m+QTz6wrPDGyj/hPhaVlAx
v6sb7ZECBmdNdaNyX53aTn2x1HDWNBQS6MyJUT5dlFCLixi22nmji0rLKM2gQ5G+
dF7pXArGVl+G6laU4Z+1cvzuHxBDYVkC1FF3tfhpjXhcHZrhbxFULt9SRQ0VculK
xcUUceJnXuYFsZ36+2piBEfp8+2u9dCAb+nCdoOtyaULL30qNGzwGzYX63SwJbuv
pyRSDtHv2OLAVMDccF+t0yO+utBw+zk7onO5lJfiLmrVQun/EQA+2KCrIbuKRf45
Haiz1Ccu1Kb7ZerNYXBDnyAEOAxPzFNu2+CUj93I9sVwZNUX8C7wscgk78ayuU7J
O6U6xgfkl7HwC4r/LMBBJm7gzcEWBU4yPaKvfw3nvJykmPBf8EN3dILhGW86ZWyO
OHfCttdR/nbfMAsp1711Csj845LMeIK+IBx3rgTMwuVlkJdOu7Wl2GfNhmGp+XwT
AnZcbhODL6mU7QklJmPzie4BJDiANLN0tAxFMAsv09eD9+TA4+CKp4PbABPyQwXL
9nFIIGC7w4FqVFhJLDir/f3qXi1VcqMshKIvtwpB1ngzilIElf9ZR8qXfOLaioDp
aVgH4wMld3lXG1OAWzgBtZTkw4iYQCD/UnXdyPCU0QyvtutFkxmyoU+N1vENgEFi
v17VGErgLG9K8IiTPhCzYCsC2dkUBzDoO0uBwjd/Yf0LG6W+pkvC3w5mOJg1SpT9
GNyxErmwF/9H4r3usL8yXiGUcrcjpRIUP2MfAZLSE7LGeTjeJH6nkXGqX7zKJUAv
ctaMqQaIuuUExVR+C5CLt1TTvQ//nH34zUbrj/kjpHaaCs8tve7RHuIoUU2EaAlj
VFMJhu82CgNJE8SLGbfKQ1qEsJsTCCOJcw0UAKV5bsw8WQiyQNbSWCldhVI5DNVl
ZBlkfb7ppu5mmVIgM1hPZaK4kQAivHFsyOtHz5a/lH0VKZGfVZU4M40FwCdlYVDn
gLwuXMeMz4k38tok9cdMb2z4JxKkkAWB7Mo3wdzyNBRTeN1vV6ldyRtS53ADAnsl
zcA3IeB2KDtyIoYP8JJLqAR3YDtdcngeKuLbaMhspDjBS6HbjAmgl0ogO6BelTLJ
zetbFn1U+CeR2igYRKgBf2/90WtsccVVDggMDRSyK1u0DuiOz9uTzInNXpkvz8us
nMnK8O2yYeawvNPGvvEUzHOG5jkBuI8+dfdGi+T5Bi6sPDHuw29zTzmZOlMgGHOY
Rzx5GXJpn8KK3l7MVgn8wLfu2DphTbPHsLbupM0v0x3tjE5saMcEYX9DJycdagYU
prjbABU48/iK/G9cjh7BvD9W50/p8K/TnA+1T0oClsxTP9hUXIv0L3hqv/nVuEC2
KEmZXJ1fYUjyVP8/VB03Z94Qkir+lsRwD5b541sEjiKGYoBJdeFgBHbt6bCZ6vZk
clYkQlL4E+pFh4D6FTuqMrwn+RWljzbXNSaXPYX6NqKMNpDV+/nZR+4/rSGBfwxR
JAtzfL0SJAb+UvMt0terWtXxVCp0Cgep7n3d3g/0H+koLcHxVgfbFzZL5YmcGvbv
N3kbJ4FRHXMbF44MbEaeQ9ofHv9w5kAmDyN4sKpIMqJAI3nB0o9E3R019pBSOsSM
lrVbQFQHcdK5nvanv2og6QSheegSUvCwsZLOswr5vFmCvCpvGQ3VcTACXmama8LV
MT9XyqGtHm/wltdozrmJ2z7m9dV+wAV7IVZCB5bwPAoHMGZVdoZcsRbQm8YAvWxv
eL0rP8pFGVRYEoEL+IQ9eHVtXn5oFAxeaoMLtSGyyDODq4ZZEDPSVHFEOG0ism/D
2KyegUQ15ZXzbFLYWVvRmGrMLutkwmTKPHykryorIGNS+xG/L0SkUUoKZNe7EVUb
NpbtObBCVxJ5/djbOAmgIX0Dh+TpBnAt1bgRzox/R12n/KRyzfNSLMeHWdQoVv+0
hNXbCB6Mz0DdyfNVEAWNbISoTJG0xInQSauZesPhHjQn6K2RFiGXelBPQfcrDhAM
JKdl+UKNg0X1kudRJLvgdXYXyx9jBoqXyyV1ujwbfDsp+wxpPB9o5hlcO97wkDhp
HtxSR9ua1HYs3gDIOzUfy1NFlbrPE2O2PhOvt+O4oO8Tc3af3KwWmolg+eRwo9/F
WjktfO/kCURMujGbRAAxkJtm8yd/sIMqUDDnrvYhh+Z4L1He6jIY1gG1AM38GRyJ
NHJUzljBRLiannFJ80/ETAn8UJhainVArJejU6VEzSBW5UfyslVobzX+tZXz/MJg
RWBWy5YC7I0L1mVIuLj5Np3OVAjLoo6Fric76upiZ+sWx/sq/lrRhcaPBGobqR/w
gtykVGIs5bmK/ripQv0pTSs8xw8zh0PRKn7dAqgAvTeKz5Suqf4L3oSQtlbBvPUc
PGvE8mqY7mzsyIKMkf7Al4sUoM8A4kk7pOWn6Yoq1zD7lnTN41lPkNKhOcrY6kWE
g7Tt2P/PXaO6ZVSJCitKOS6W/EwpItIQSo/FCTMMlvLY6/8swr+rT3kdE2lst5Cm
faWhDGzuLKy5x9aF8c7wWI+PAmC64er8wVANNlAgO/UtSe+1EryNf9AO7cLglI3X
f3UiZIJ6goOU30AVCqx9E3rBrrZSJBcIa5nP9LQ62EtOv8ckehEIBC7rMXLzn5ie
BEFZRji4uDo7qvmwCHroe7MtQZidLnRJBg0V7XV196hoIADzraJD0dJUAelx1u/9
vi8wLMmrDttWXwmAJfWWbGuuxEw+wAGaIw/JBZiH7/zQ67tQOA3YKPYwIYyUnWfV
XIXEUM5aKkb/Q+0eJNDzkxGLH7grJDZFYuzKP8GXMHYiuhO21bQQCFXNvbKC4Jjj
g4vdpp69Kl9pzuwYgkF4UtQFqIgOgGrYcbnASJGc4BNwQYSOqX0+R4zjsUImLjTZ
rvZTx6cTZbLpiQeDCnlf1uijpHa6HVphIPyHQXaC1iPWnFYqT3RAm63kFRlj2lcb
eRjJduOnQvBw0h3b8hE2B7Ef5YFDIxzS5BTdcrjnXcN1Rc+v0ESiQF/sVbKTY0En
+NZt1ll3Lcv3U0MddslVslIXqwiy6vaYu1rw4rL4PI1SzFIk6iH5cQe+RFsv0pzd
Qth41hSufumKdQyG94vumPd2QVo3SE9DNEiwBuIlTFymMThBsku9Z2++M7Ip6lk2
bMadJatS6vJqmNOvunW4mfp4KkNoJiHXBFlGDXGsV8EuzddAeN/L70badI6eYbH7
jsvGK/YSLegK5y7YJjN9x8c/0LsgSy41vu4NnO7aYKO7OpztXaYg20VDfqhZ4QwH
hYaNLc8wRbQn6rFXCGJ9SCAAJtcxBAN9oSeuyiwD6/PYJCf18wASe+IZlGOQmkoP
fbr9v6Zzz0meaFGoHgOr6Fh6JCnOzfLIlTgC9uxyeWiZcoBN6qqazj4Eg4WsOAnk
/XR0zJWiWaWf82kLntuLP9KxpIS+Wj6thehCesqVgHSMkRkzxSxDbEtAy0w2DPG4
WsO4QfjOLS11DlDGC+Ys6wB9O3MVQpJvotitmmc0//sZPnLSA2fKwyZDKGPczm5T
Rvi9tfAnvA1Tf0GZfkwm0yWRo2sjlN9dMJ226FG6+pYkOWmgAAdsSW06j/knCSKA
FMowssxkdThCa9w44fvLGds+cAJkS7TKWuMAQMIT45Fv2UtNLjQoOq9EIOQjvzc7
Lif49K9VKcirW12yvMQ7AaZ5TWr1X+zxm7gHvIXptB9wxer5yGsI/qcFwjDCI6Ww
kbZTbHcDozu9+qjcRQ1yf8za7an19M8JWwav+5h6g195F1bRI/hUUntZFRZ5ZTqN
C6ZOdPguJgrjkHLeSIVPa9UG3zZlOEPYLP4VR3pB97yleiEFp0dGWNzbJvhQKwW0
P2n/2c7/SmVl09eSbPJVt4PMuFq6o3zfTiEhic08p5cPp8FSSsZYhPZFUgAVi89t
Ltb2iWoYkoz4mTzsvzp69/f8szvFMjzkrnUWWR3Oc5l0aHQkxJS4utM0nHtr5mW6
d4mbU7Ph4SWRqJ7QWWrVA5Sl952xuHvUoE25QNDXp9flhLTzYiZAHm2hEMhwm1Yb
oQeIjvlALdpAndDsqExD+RAe2OSNGo9KBw7kt8KpKhfD3hwsH3Dn+/4/0rulCa4J
0A/crh/+QSYHrv1P28n8//K2+eDNnYdSe4rPsWeVBKztqUXecmiJY7kLoPCJMg/B
bwDKZSuEzPmTlMwSMTm5KphE9d1TzYJLp3PvsH59yu3jF+B0ZbEOaWf4O++Fz+5S
75vaGizTm3DHHmkc3RmuPqev99VfD7mqqaM0Lr+LnAjzlye74hUuzoWTRT6ewR5t
/aJA6fOK4VkfNZS3hrq+JibXqHlBs7BW6hc9otRBoGPxmgo1tJUKpHhIqyXDhzJ0
Fkpp3f4b/LZRJPb6xrcvKZ6LO2XfFurJ9Qh1aMX2+lG+9RahUQkhnt+piQl+Y89s
x9yXVY4NAMheY9CF8QfPSYy1cnYI8oPs/QO3tGD/zkBJMi3l1iOZTqQnxZQyg3VZ
kxL+Hg7dJicVPswU0lRoTyYDNnlf9VDOyp0BFGB6B+Bg9I8RljEaThw+wpeZ0x4d
YgSXpFQEw5+esD/fC8Pc7r7xY/+No9LYJLjbErla2g8aObdlpNNYwT883JP1Vr9X
bMSkd80DhI9JOD2Q9LmKyRZaG9iOeAXqSw8t6svVLje/a7Wi/UgqE38e/9rcK/F1
Tt0FyUnglRE/sojx5CztNxmfNpq9aL/umTXsZ0nihQbm/hkNwyTfHxNOB4q7MGzS
+zgzCWZRbuDHHWo/vYRYTXsySUlJ4S29Ry01vDzE2GUum4mhxnob5I9n02fIpPO5
9r5c+GytL1HVrUNfRTTXsQv/89hVzuOR98pdM3Y28haWrrBWMfDtkBZGClJ8+ECh
pSBv8HRPdIeG5JCUe5RUR6MhAAnVH73qkDLHpkNxU7NFe8yxJjQyNkW+ytmu58oe
xfeJYZeICjgjFuL/EG892BIfRbDUDxXTyjVShUFj5EwiAhtvNMvIvzVR5estDcj/
412dveUku9ynZls4h9BB3+ceOKvEzrWDeiTd7ao+p5Xb+eMzOyBDsqKoCuvWJ+/b
WVcacE/MYcTPM6QLxL6Rulfc9wAgn13d218wqlIBBmMfCRzwS1vRWvNTfEjtmI2v
+yetG4aAn9SuDFMizm/2VbXFKpuK/dsUGh4SdJZ7TyXQXvK+6PHbHQX/AGYk9yWk
RYtUc2Bi9LaIEyla2PS0baOoqeFjsfn/e1wfSa4ycLTW+jjE0ZvlHdMTa3phQyVZ
amSPTy2NTq/pVEPjYU5L6hSUjoGy/5Odt8npwVbwWBpgBKekaigp7rz3leYQjxr2
yn46nEKXRLzQXqO1+Y6gRsPw+I5QcR9J0GHGuBWIxxAbc27O6Q1GemqYlsBQjHja
hs1rVg9YGKdlgROUvxqBWBD42lHw84OrDSjE09zMsPZAZxGgAjeIo9exn0aiDPLb
Kv09tya9RSCKy+0Z4bBHSuwVhfcB3auxG4DDnQzBeolyaRgEbKETg/KfWA+5boy9
oTJjpEMk5R4uITmYCrK8OaPy4NmbvYXQ/TlAD36jLiRRo31U+z40+idJo6hvp25g
Opl5bBs8H7yHXpsC6qbhOkR4/1yAh67FiOuO1L61F/j5E6l/xbZARsF2yI5krtoM
IbLqCaKVu2B4b75WgOC91nqGibRzDjWOd4LCWFar+CrGyK8oYV260ABAzweMFMa/
DKtW0Eb/vI1dQAUEuc+rFVET106qVplNggmmN4UIZsBwiIw69IGxQqYI/BrOe5ID
3jWVwlE6fjFsNj8ZFt9ugVB1qKvzqg9hiwhymau/19duBKE3/HNNOlYk32IAP/JS
6+BmsRX2TftCeR8hdA8f12xRHoZqgpMQdoRI1uvCWxa1wlI7CKOcz8CsibqUNwyD
Ug5KnQlpV98uyJ/wzsJU3U541SSzuthfLOpaOdCAaoNsM8O/4lZazkI3UVYXKVNk
+oYOx1ryQmcMdbZnphTt/xZZ/XppkSu8i3il9xQd79waZxCUrMIZV0TyLhdAxjyO
r1vRBGsg4aFS7KWHrWuSGpQu2SrMaWWON03Z8uvw2licIseJUTYx0pNCR0xf4NTV
JgJMXLpE02cYyx5ai1atGHqdpKCCHwFeqLRkjQmq0gxdIoPdZ+hWSk6TjiW7Ycpk
7RYeeYwqDxXJLMigvSvQPUrv6YzXh2iCk0QqlU4tHJDx9oCXdTiM9B2cnQTqauIb
OhFU1JxSMjXKOxecthJIzEz2anWS10HtPUeZrHhSlfQcR82wPo+C++8MetZWhBhi
H8Lsir+WBIJlBBdX85SOxOH33f1Gdi+fNAVZaoa67pQ9hyf9j0/Gh5gHxQUhw9RZ
+H+FM+GQLqsGzXc5mZYeQSr9uAbFRxmX5U36H3qVL6Mm9YxPT0Fcs/1KyGs3/uWl
xid2usedR8nSiu6r+mbSg/QaLGx0Q7i5ewVdWPfj7zd3ID61KW1cI6UtIGAewcuo
R+E+C24RzA1uxHYRrkhNjQLBGOR0jvCNqgC9/7T81a7a1SO2g9B6s257EjHSxJFT
HIS2SGN176jXnY6jB5rcyLe+A0OPHVwrPCUyM7vFjpSiUD8Q3j2C7/5dsYkk7Zae
+kMKDUfcPmdKxMWkFTn81TWbxpLVdmQGo5myNfqJtVJMLhwpUS0Lj+E+JNOut1oz
v6B+zhe7WgBTk1oXp5BxYzIb/FLrbu5QZbj/qAQ9KbD152DwOZhA9zQI9A+xTqHS
kUEK3DkM9VDNr7PE4Iwmdixd3lZEbqpx6zzD5elkb/IxADs3/yP1hCjw8gB0SwQm
nuNxAcPWO3pIvOod6uSqdm7ckkrFewPdsHRIEI0CFhqxiYxbCEimieKGZucCKBrW
L/P1iE7RY276ruF1+Vs/0b+KzW03BtftLhyDn9/2cMvzxv2oEK0putP1eHctORxe
bsBIFUecme0XCDkDqX/MvzGBLoHhw9M+OVI1PffZPYkID9kLbquJyouP81fK2GNe
Iwpbp8N22ucQ6C/tRBKyGGlZyjcZxX0r+tewrODYawou9c0rsWrvRn7cB9N8w0pT
48PN9O5BUAgbwu5HD3p8Sac7IxwxnO5qB5U9zDiwT4Lpn+Hw+uO1CMKSCIh/jPnP
5AIH49uY9ZSzLQASfQAU7S4t6sIIgv/bkEYgCtExVGnx17LDbd43ClnTldqVCfly
yfoTestLOLAUwXaFFrFz/5fMThPAeodBAq/2LuzQYfFQvgTTH3B6hWrsQnlcYJxb
YwenCJ0qgwBDYP0gbp4B8sRmgRT8ZLMiqPJ8/8UFZAnhAOyLnq8D6D1G1t6nAGdI
whJwYm7t3mnLPUf2Qqsse+ibGvLYhlixS5VBCyIOVKfHDLNEgdYZM760GTbJecNS
h2L1ANqzVhVrT7/M4HxLuX7ZIZmTDx7Lrb9NfxzTizRywk5Qg6N6zGM/IbJIGXUd
jU6KxtG8+kdgvJdhISugop6ngDbbt/DvT9dmN1sD/AvSPNo9cVJ5C4uT/b2ZcTJ4
tcqHZ6T4J6VSkuS0qDZsz16iBszsOpLCoVSuRiaK7lI/U0RPt8pl0OELtGKFUOrS
FhLDswoHB5GlS3XyPVIRVpm+WFaeu5+bxgT/PRk8PGn5VSKGBog3yT2s6cRM1u5o
TAvBUo7PeEjam7+dRMlD8A3JF5sVuGt7Elqcqxn7DRQepXYUOiPbOXCq8HpN4jms
j6cGpY04MJtFbHEzQffNqilFcVA+F8Faum3YthlHryy/rMo3o9MYzG8QnlphKN+u
5Ez+na3URhUlHoT+w+FZTAQkQWylIccpHIadv61BCg7FOI0bax31fd25aieiruYl
P1JTQe/IcRBguOe7/pD46r0FtsGt8wKUHXNcKC9JHzg1iuhv26APYN8x+ksCq9Tl
0d6U4z78NFGH8aoPsCg5FE3QUT5Uj+qs1Rc88ldKfpB8GRtgMs4Hq/jmYaeV4GQu
Zx76KeDOfTpOdvk0KhCkdVpbh0Ba8eHfXuDapHchUqELivNTnfWar/68W+EfIXJR
JjyRcr4Ya2Ir2OaDQslD0njvPB00geltTZZoiqufGZqydUgcNbSd+MCI/oQuQYGe
fxaG94d2fXLi4pzFpA3rzsxfewmdIkqGY7scLEyvKwJy7hho3QyG1djlrWjONDCl
xESY/Ru4jw8KxmtsOseANrd/XnrxPLt+3rTYJKJ9ITbgV2XzCnndZ3a82FD5eq1F
2Twkdgl7OF2+OO14DJ3EVopk85vIV7qk9tWhGjvIWK2EjGqYIzMY7QRS7flFLVOf
ilw63PaxQ3v7IywNt3IGIS71GbzQeXDdeP4xFjytAX1OkUtgLFgznqgjwfzLXcBa
ZJPALMh9ungjwY94LeH7sHdnO+o6zKh4qDRzeX1RDIXTyhSnF2uN6aVrlHKKO9yB
XbU+i9qukh3gTLNoN9+P2y0MLUZWFuKi+8+A67mctHQoX6sCVlI4dN3Q0ODOEhwX
DTzgZvyzgd+4fdDxhuVkdL0p3Z/mmZ0jv8tOo6SQeUt8ST75b0Xl3E4xZ+9DwUZA
d9IWMZITtQGOiT10NCZ4j/mgVoWOeFRcW4GIl1NfZOuQKSnBCmJ9SpsUuWTcG1nw
ZZoUQR9nOrBWEEwHpavRJFoUlK+NAKo/FWqs8nBZARb1gqH4qHukPfzwzWna+a+c
MJUen85s5qhtnA801raDVcK6QXaqeNN9872QIhqh63Xs4Dg+c0PuXNtsOTS7wDbT
/cb9VHNrgpRdR8mrbQw4SB4DBOPCa6G/b0vPsf0+zFxK7TZ6NVFHEmsa7Rs8ymOU
KgP0EfgvUaXfULhparKXwi+oPN761SIPKp9d2L26emEXk0aTFwVO4vpAFVAoONXL
+rCU9EeErVk01SI8He071cM9F/EI5eN3IcujeNdmmiv1I8J7yUvmzcqsrlkeS786
bwHql1nu27AEEML4D0mT7JE258dzcUrXn1XsKDjqHHcgy5unX9BtBEKZuJzVK7/E
G9Z+KwmOunU+W8oXZajf2hKTM+V5mXtWb4rjjXLA6rWNukYUrfvZZU+fhyvD6GTi
JCcgE8TNriovNnfMKKuW+NQtlGO0fbxGVDUqnKUdGpTJZYQioIXSygIr7vScjvIO
3zBI3l4M4vIDMcjyHiEBZYjC3AvGQVAqa3UbjLfnKenrzeU7gsQu3th1OFPgy0rj
Plf2fZfnaKzU9FQXezWLtWEKGviFLcp0ugx0Zu/s93lFlrasrRWcdpqVNZ5t67Sq
H/UVcpq4HWSychxZaqb7VfvP0V4HCzNAy3HInCV+KW57H2tgf4tEPFbtYyn1dfNY
9Z29nuckLtRtus3yPRL/QlzvZcWBGE2Id0m6SR7ccpZMOOKKBKMSEUjTxXqor4jS
DgS+LnJk12s91/NCwvRfjR1sACafuk0hlaBsx9OEH6GXXdJW8SkPRT3WGHAMQX57
FrMUxYaCepUMqxXkMdiaxNVZJAKFi5/mrSPp+040N4N3STunMgRWzW0//rHxRDEK
65pE26fgSKmw5jvtf2Mip8fi/2BI3JVnK5XxkDr29VoxPqxLnvt+THwc9PaFSKMS
i04g5hsgXW5BBsTfoo7Sxtmwpcm7WaJtOBvrA64BM9b/PnnT/Qi4YS3wpXtHKZ9E
QfBP4mnxxj4/7X0djg3m2JUOzzcqElsObqeuhWZyMkrYVNmUrqYq7NgrEHevQMtp
XP+5KYkpJD6/EqbuiF5Is8JchjTXm/NlHPuSuRCrCwADt3iboQNuKLomUPTU5dMd
kWhxPqacw8Ru42O8D4nXcNPVMvYYSompOlX8sZ6eXXmd1FOIsYV7SvwES66imzjG
7KtMmP0lnZxGAx3Tvr4r+FQd8M66yKU/zHwy2KfpfS2uXGsAR0i/w8W49eg15yWI
R1sbxa7Vx9LTU+XmM5Vkf4Byv8p64H0GybWTDKi0p4N4FPihXhxyhEj1uHpEhGcu
pnW6PDuIDIsvKWECas61rycGxUX03YPTOWdtO/vwzMDmvENvNusH7/7+HNRp/qw9
FJghGPkYCYUL+KH5TOHXWUB136WqRf4Abvqdl8vMrhigy5va/6dRUESYGftlchwx
3teav3gQModlVCarWDLi+n4Hf7TX7aNVDkd0p8hPhPkK8GJIelMqLA8IDJTYpqTq
kfAQ7XQ098cU5MXseIAqprpXrTm5S9Wo+eyXdthfngyV4BpOdk+N/jHTUAQst8Av
stGpIWFAICEQMXPE+WV9frpIfi2rwgZ02XHnzpyCutScOU4gg+p+cZ8qrX7UC+so
1Zaca6vY4mSCScqLZj3y6fIdDa8gvIfoaHFxtGCg8y7D6+uAL9TJplvNeTtawNCQ
OD0T37vYgUKUgqI4CWp5LzFU4kd5aMWJsRY+gq5tJ18YsF/ZJpD3hrrZhK88L3l1
GnRat7LnBAiuPA7/vVPvZHKNyx0McxPK76wEfveb0ho9spxBZ/CuCITaPizyuG4H
q9vsQhe0w317z8GFDkEXUOWriiz50E+A3/pXQSsFHfNtQXdKRumiyGXfovEWYtLB
3YadIVFMqUr12s14v3QYnLSCcWhHI/AXMVJ6iz4fo6B7VgXHFeXU0uE7rR6UUNxH
p+Rag/N3t4m7ZDip3bpvmgnW9PayzcY2WsPZk44PU6uX/Qlymv5nrYBEcFLdq9Dc
0WZfnmWiJhwXQbRPKtsyylC7hc5p4UM57aBeA4wmQ0BbvWXEHJYAchowj8EH4AOq
o0BXTO8beekwvhaMaQfIux15yc4ohzdJHZr4Nx2MUKHv2L0PEvWuuH0qsF2Xg6u5
Z9xH3yvxAn8kgOau9HMUckX4TYli3C4iTML8VXl+eBASd8qQpdO0LVyOsHAugKb3
38U85RI2YImj33JKLpnZLy0JnNKueG5XZwpyecF2B7++slfe1cV0bo4yDOa7RR5k
XTAq65DIQo61/FB01XF36srQvZf2C/KeZ3TB6stCIgjgSZrmnvnYBbCYT5o2VLzB
XWlg+eerXHe7prgihSQamVjt08psVUXo5XrOh0R9wYqiePTHR9ayH3Dk7spwuNH+
aCPHuYF+RsuXwmcRlJUWXAqK2fwzk4luVsa3e3K5S4UB/hX27CWjQ0EdVL1iKPLB
tDA6NHLyHj18T0h1Icp7YNLknbwsk3XRXI62M6PCz1XXrUdsBOaxxMJac0/he4lQ
kKsXUhnDyo1fNdDXhZTBdShp8916QXBjCjlA7ui9T8ktwpiHpx/OYhxWERor4LEP
cwmT38R3uiYuTXTXaHE2+4ovSXSmBxjDaf4TztXiLjhTbZDa+jv0j5UsTYN71ZKZ
MUINYNEvsPYD+dJHoYKY0vTKaS1cnrEk3juC4OhKssWbEzNyth2vdavNUtvRXCgl
q9u8uoKxQeL3wQ3PEiiOdfgQ4wuPDAynKWm0hqt7Jb4++dXGvEamVv8LKhRwsByJ
aBOQYm8Aiq4l3Kk6yx/ShCsIl+krf1owdsMG1tiNdRkXc78QtwAFvx0rj/d8CMyV
n+co5WqQW/t3eb9ZwZ95FLCCoItRdLRj9UDm8MBQhKV4kwxjUFfZ8wmpPEAE19EB
8aK9b6gvAUvBQxxWv7PPCQYukPhXvG575wOfPy2Ssixo+c5e9wVGoEO4CexlobWu
KowRLTghNzgH93V3hM49TvvjGHgMg+usG69xZvIOPFBVHnSv12EBXIaGSOVOR4Js
fCEuDsVwRFzFi51uv6f78bTXxi1axjqsAQnkcLpGEAEslgFuPYCSwq6e+MaI9Si9
ZPDljEX4uHThdv4W36aCS3750BQktKpFR9cbP8ul5oZ0tX81GDL2cJ1q7k3k/mJW
atBWDsMxWedX5Ft0GDKhU/B4HguhqrZSGXcJxD3RnY3FSyhvjC/4AlOn9nLsQbb4
JvK65gjcoMsRqOcAcNCxmx7xDgLMraYbFgbXIsbHDjfLXhHM77wsalLDKfa93iY7
EtQCDAxYiLN/oL94bYqZj36/mpdDG7uiQwpeBGGb84tNf7Q26LYpn//efMPMXfzl
NnhbE+M/OJbmDKi77HbbOnNOwahAqs9mIn4SPk+IMiMk8WlWUIm7PXaWbO8aNbVn
vAZ7RmCLIy5yRLy/+IozNxHtCNXRKv6pqWM2t2ULnc8zY9VAMETvfRA287F6aERc
Tvq/1PnIZZ2iKfnXZKxnXm52KP1xQHmqk8VJJ7oV1UBeTECXlVjUIk3yG1QIuFYH
hf5ySyGVdTd8AUnAkaaItxoO7W/KuBSrtOlkcZ0XhDpi1m4i2OAhU4prtJZyCzQ7
n71pGF6Q5Oh4y+4KiWEt7ucRKl8mwXIUdi8m/MOJss2Sv95+cTOeBtgj9/kHwwba
N73TG95UGhLi8hSUv50mm9/8+1SGeGJW1HjXdSw20ajuaA4k0w6F8IwLxRnn/rzo
309T4SdkmDufb1CihwCYlZXuly/CqclarSWrILqZbyd5D/z6gPfOvdnZI1AxJ+bN
vaLANlFszU6NxyW6M172bqcj3jlHltzD0qEPNEcE28F1LsiJXDJ1+P0hgU2MgD4l
4TYaUKKEDGTVmPM1MgXEHwVkwT6RJfR00WRL+YmNgoVU/73/iTG5sQs57gKJzoco
czp6bXp1gnUAOTC2ljWkt6BQHBFS3aekobIdS1wSVwNOvMki57PxXSDFVRIUexlZ
TWVIYL5cXhzrxZsJrcoBilnwCO9r/tln3SK7+UCyvRY+yvOczugs0f4EIQMtt7ZN
ZXzx9BQaPnY1Lov35G5IhKncolGEiOMDIkAVlrSF/uA4NnOoyasyTjq3pW/J5Ph8
8Rqk88p0u3PahwJg48dQzPU9zPwtF/rjG2HfFfbKxH8hiYu3RS8P4M0stfZKNLzU
fkGqpc0/7YTzmq5r9QjFRWlXboI5NS8eF59Qq6y5vPLOgSsLc5eXhsAw2ZVfa+8n
C1g8S2DmdRg6lxdhr4IMiZMnICRYrxIlor8nl1YvsvXnVpBgxpdAyD0200oBhufG
5X/qL+5XRSDuXOcQzMKTTjw3bQDWHDyo9AaRermhyPaB8DAprx7nYm49H4gIos0P
zDt28H8TbtHUBGKvNbiTb2KS0ckPe961Ltv83dig/J5yhSt0VVqqsD/dqCBC/uYo
DdAO9MUrH3OD/ozgxKx3YmXabHjnineQbjeDT8KSHQ2o0qU2GEs+KubTgp1hRE3U
hPjki5f2B2ACT/h/1wG3iw8mKxrN0/9rW4jNXlGzBaDv+zopY5wdzw40dccNREcV
VTVKWpnHhdBwcoxlBHZuJPUx2riAl+gnKu3Er7f0Gr5jt1G1FUe1HGe3R8ROr8SB
rYbsC0xMrdP/6euVutQ/iTiOEo7xMtTX6mG2BSGtpUXajzqEel5qIg9oqbAxaR5y
7zQGA9uuTSjpfjFFQOZKWzx9jNozhelrUw9qyPXMnWmYzcCfot59KqA6b0dzvUx+
ZoOM4OrHEEfjuSFMbIVFriMjQqmdtIWgJuYSvn3z+eg5LIZ7e4V4+jmuCek4lmGI
5nPTBENswU5zkdSwzoFh+KPTjrX4H5VEgBJ/1RECNHU/INdTKVQs53b4yzzB77RN
t2sDTcoZ4+iPGYAEO5FndJZMzMwKZLk6rbhQSLL4rHaFKwfKLkN2I4MJN69/wTxm
pmCSyeTmXn+G1rr9kD1Ht1iKC/maQgoa4n9hwhyL/tZV17aU/svYlyzyqxMc4RHP
mqEm77xR99aPiH2bf95iTPFSDOpirrQbKk71rJC05xzbvgjHVo2EE1LlFdembwcO
XBF3PMF2xY3JZiQaA3unYgAPgazw8rBTF/uLgF3CCNwsJpvCHqEhLqCxD3zoZo6n
Xxrt978NFayUrIKcdRWCzBOW59HZdqNl9+zlM9jV5Ql4CshKG9irwM0YxPyD4Y69
7JVMD1ZTzj8MiQ20XUyNzBWws+C+hIjLG53PVRyp3m5vwazGa8rMJoO//tJSRISp
90Gj9nwG/qUzJwPxRgLKjEQ5uVj/pKzTkGfp9ZoI7bMkr37KPGl35Yug5D6qgOnh
sUwnvoosPoXPuVb8hmoSX5W8h1qdrxAqujgDo1RSwwyiWHDTHUn1WcLpH/23Ku5R
lJ5vJ5+tSE0tVZXAXzgLFw+tF71zoMFYhG8broyUIFJWaEelG1019bL180Dwv93Y
y7J30TVDNWX4lhoWWywwhwC4dYs0qwcBbvJVBofK6d3iZTMd2W9LUShrFIxcKBuc
Xlc1P/sMfIpZt4A/yebs5SEPd0RCBoAKVY1mzjiYvZZThYzDS6S4Mfk9lZUaFuAN
Zka/tVqqPFOCLnn8lSmMiLRnuzloPH+VHgrRo2vzC9OPY2oOuJ0uHRkrclJ4sSCi
161LZD9b14hIHiWyfD9mfySmUJGEqztQY+l+Z3u25HkLv75o001GMhz00GC431IJ
p8ZrhD9xkh+W8ELtJzJTGlUQ7RVK1UNY6t9Pdop0gw1M5DjhvB7FU+DQpeCAxFW+
egO02DYv4qUZNC41heWndLFuC+SPW5x2DAo5ous8kfpZdxiQYjYTCbTW4cYB3ag3
N4IcRQKlO77W5Fen8Jk/IX7LN6e9pUsj3jxXgqdyFMcXoQwAseaET5mWuuPiZaBs
Ki0An1JvDECfEaqOT/NNb0UYL8NibhHqhe7p4QyQlxxNZHgdI6FZN9/j8cGF7QTK
+xB6M3V1h7aAOUZFnMH/9UTGPDk89w6oiQfzx5CihwLDSY2qQ9J2jiM/bDlj/n0U
fnYobNi4JTSV8/SsDLbgXhhYOkmaR03ZQVgLfXFzREnFKYvD9lKV3nADhFdEDrnb
2wqpg8oqGePT2N2ih0P86dgu6MexC3oWFcB7PdmLgm3GPknVxx6WR6IZpBLzHl9+
hdqgG/UfJ0oqMoPm9/kW6NvcNoiITlPGkPVvomY35Phf0mcnuMf+pjTWfZBH/MZ2
mvynJrjE3u0WLMw9Wfv8fVtTZ1824CnuQUw/RSyDFguAjum5CWSA6TX28GrnQ1Ll
iz7wPahrmvyk7iM668VYsve/AxwCyMBSeuM9r0pbmqOEkZJ2vXy9tSNSajdA0Gpn
0Xx/streioETXPZaxFurlmZkaMu8OuYq2cDL6X7PLeuSxuZQq3B6HUT6k1D84kYV
M7Uf1CX4pt4hKGAcMyDKzsMRVc7tw9YCQtYQ3cx8p1GTB8sirpLbeS3PgeT1LsP6
hEAzH2ZndI6LgYMq7SxgQjkVKsSAoU/IHL9MmbWOJrUOonNq3tfNqu/aUiKmFTSS
x7qanqjR5kjbdZPxdXTHuZ+EKhYaFe4q/eBfyIBRWsZ/diXeSFOpCAXuVX8kCq6e
X3c45GIuEjf8TTdoL0ISHjBImFD6qHn/bi0vfBkwbXdnUpnKQgm9JORbCdlOWrw0
+AA14kUAqFEb8bcARDwEk7f/M8SSZd7DYZ8X7NB8D0CDE7/ltzbnhBnWrorXe9SF
S9Va9QbJXNmxBNCALF7asqAt27+Mt2njYUekrdt3a8py1XAwpvaVz6gy6GKrTTTu
YgFOeXE/pK8EspSUvI95cB0n/bnDGJFSHW8DZKMdWFDn+zc+IcFa2cGV3a7SdDTk
W45inV4UsiCWf+63stLlCdVvsKv+AiO907+ovXrLNdVGfgqcTKLNsvPQ7cW+DVFC
8Fb407NyPpjZfdJTH1kAQROum/eDfxCNa6Mk31MrW7DTOPA0hAYoO5iutmA2OtB5
d5T97BXvsFt46Bzev/onDcbTHSpvg/zNGcq76Us8F2MEHoZTU3QdKOVdDwNl+j8c
++CCzTP4a/MBBgyr4vZlkMEQDrUKS4KqVyYlG1kBdILzFK25MkNAnMGGHM57UZUU
9OW+OzdtYtGjnvaV9vLIQMF7yVPXmThVnUvdx0jWW0AE8zEgHJ/XJOll61Q4ZLZs
o5Suf0XiUbr4BSSQDmh3oNboapf4/hFMPXGSuCe5UTyTC1rSYlIhqKjXFDUhsuqL
m0+1fXgEzBiWVO1cwF/XzcCEAFLQExf1rizCRy/JpGR5qVzMpSlvtxTY8KVKP8qy
+NaWP6UW9sBs3GLS5FxMe5ZPacLIDJVb2iJ00n2mX0wRj0icDyGZk3s4E99irCXc
KUBYqzE3VlQWSvcSePzdfmVGLjG2KS1T5lLAiojeWYvWQODdTY5i9oDMKe9CMOdt
70qIL28wnN/xok+XPbMvoU+OjGRD6LTigzD7NYuDBdwOhtW2vkMRrktBPeOsv218
G0AUgmZVdUqgBExUynLgfKSYfaljBCFGeTY8rFAj8U7+RKY95UQBjpjn88VAaXD3
2wu+Rr7FtJaqL21YBqZSUrm5EhuFBEYnPLU7mTuF/OFkNUlnnNb+GR58h5sak0p+
HR73sbESIHq2UI8UhCtAh3aSqPrO6amrM7mrHAErIp4DMEz3RFR0bLNdc7zBvBTc
iAXaWjISjhIzL+n2vYdvGd4yy1JeIkbGfm7Izqu9/gvclzr9zg27BDL2XLWYIplt
+UQcizAje8Fv0xwUsx4XQ8YmhqQdc7fCTbbY1XF63MPiBvFlPA6lotB4jDcVGFiU
JdEm7rEmPIWT7ygtvSz1p1o+70j2eFNN+9vq2NWx7Cxw+cs/hqUPdNK8vBnFBb1v
iAUGzghdOGMVFDbTCpNGHg+q18u80sxDUSJGoTAtW5i1W64UGCJ6Qhov2jDn5k1x
k6aLcGfXYG2/AdQRRj/NX3uc221hR5gtvmEy5OKiZMRC8aYz8ebodUDKyTMrArAI
enG5/xeiHW3x650u0SHo0wIgX34C8IiJPRNEfEVoFxKH/M9LAUmUGPAkjipVf8Rm
rv9U58Lz8b0Q7Yaw8m9ay/oRpz9iGL9tXp4G6/9CpBR01alkuxTwqWzparKxMJcp
pLlM5Al+i8MY6sUnMqXPhqIMouF9Lug++IseM+KPMgG8lVXCe+TeyXULcnMT2GqJ
S9C94LgP1Bof+keuXVATl6Oyg2yH+fqmUXYDbmPlVAfMixyvXOXrmvwZ/xzVJB3F
jMe5IUNyCuXiVqgB3mimblpNpytJ5wuPrpBPTxiqagk4mDFPI8o2HbRogXQ+/yQE
lUg+n7ll8YQWPScPePgwo0j3L1bmQiIKKm4JZwUgecX0HJXHCd2e1o3LemwBMvpj
nG5pt9U5VC2swtXiH+RUTQp6BCRDSUOdtfKR8KOUDhhbiEAY2PZUsZp8tfhp7zmP
a9t+iY5bUXCkIOBliQ+dBFPrr9K9mjdxCWpuecaElL0qdRHBbb8dliK3lYZtV8Ng
xs2YPxjM2ah2QJ1T0mM+5Noe3SYnbX/MTa90rdp78lV+pXAQ+vWAmRcQcDTzWXk5
2RoddwQJEq1o4ladm37uYT0Sz+lspNLhweOlnkqUbYX4YwcrC37bBdexJazKIk9c
QjzP3Sb+obo9pNGh4wR73RhIFjViwLjAuyJ96sf9rYUEJx1FryDaXsxtR7ju3afJ
CDo99BOuKc707Uz9wNoKSZa5oleW8qZoJFzEVQtYrqLHvx4aYqJcpzEjgcASfC26
UQzy8kwpyUUfaWV1V/Wz3cdhmGKmqn5lSFpv9UIVRgqK2Pl2GOhNaZtLkTI+UwNT
yZFDws8PQe6Pu0Mm0NmbbQ1noQqgf01Y8GxISndul681o2tUeEcUQwMl5+5k0QLD
szyGmSX1x77IGyXhuE7xnFgrW3Aw31KwckIgRssUhdBVrWrOf04fCDU2znHdhZe8
GkXHLDSHWTcLZxUE7DZg66C0Cbz5AYWQ6D5r2g7tQM0tt1DaaFcy5aPYNRzcWz+u
+2My6XCKw6ZcjxnzevqhjsfJvAN3pM0xBREhUnh/GXQ5hV9TQaceQK6ZiOVarayz
MOnK+ebidcoxzDm9aaftdfuA+8DIPV4++kk7VKy5eE+T7GxxCiPGP23o6K5R4V8C
IcLW9m/yVoynyQ9UM7EcSZikBq7117j8bwmvSueItRvfwPqFj6tSvB+9oAsunW97
j/clsypMe9OD3pX5e4BDj25iV1vIjX8l+bI/zneHcPb6XY4oe9bSEIK82dFZgPTZ
PaOqNi+z/25kH54bAIKZeBYICpG49ZJEzpVzThKNykV9t3LBK7k/3cfVTzQnZ0qb
9vp6msGP8xm0tocm2mBm2r3wtvXLNO44S+V2R6yfkK9+dRf0nmx/kQ4z4p+vGUox
330tGNCmzBbiQfQxVhk8krPyyj0z+ziffGcwMB9MArPcUX3A4iIcS4iqaPhtK68Y
WE3Hm9puTy3q/uvCYoxfmUbFu/5m1AkoVooWYRNsLNDn2e8q4PeMBRGo/WQk6dRB
IfQ1TVZdCRbgSrIZ2m/9eyoBLqr2Yt2cKHFYI3wkO5dtPgt4W/7x3LXQTCU2n3x7
EP4fxi6dMyiHALRic1JQcZAidjJWfgIG2+RDCK8MEoT/yC5baIIPwmdsoOTC49fo
qtgt3K9PQ8xuNzm60cVV3JbcyUQ6tg+Hr+Ww0u+P3l36Cih0/lZZWuBDpbNrqWve
S0PDTrZoNAXM+pkm9UE4AYXyr2BvSTCshSxR05Ncx0t1o+8F409yKC218d1+FaYz
F/swCLfvTsfxXS5V17ZV/wTSsWPPCHcGKgwazuN4nWJdu6uVcEjqgyVyUmUFGbMt
86/zjCteNpkhd5k+OJr+ryUG4FvWjXwrrNZflJPJZd+rHXTgzNprf32teX2vuOSZ
EsUSFpp4jHIjZ4NS1FPNWVDeqFYU+JVtYpCud9wT2xvxxmaoqI5xG3F4QY45JsqU
69LGDYGIDRGrLXUZedoVQ8n/S81AXC2gPQoRvQY+dfRhhgetU1lk34HcrJTur5ED
7fWEKyss16VifJMA4e6EmvdlkfjuawEvECJkgIB/Xfg6Jg8407bMpyjos7e5puUE
qZXEq9mPLHfxkQfE3dc2afTUlvDKZuvvaBgGVJvDS+/I3S6CuCXK9UVaFu8Dv1Hg
M3t5gmXy8Z6UnkU8oRk9ElUOq/k4NcA25ccDtpgFn6xxViqDbJdQxNs3+qd8J5FS
gk0+dKljCvoabKmPyUO+eJqpTW3tlSWDs8EKqZ5FkP+2spqv0Ftoj8QqzVtse20p
esdmarL5yXvqAA4TTlyL7n09RYQdHRaM23/zIfIGo4S5c0Qaj/yMu4w2jMb+cZxw
bORPp4xGYJ0hyPBZEzoSgImt69YYvlPlMfEnVfRJhSnxZNFbqbnuKS9Ns/jkrnmU
yjF5rp9+IZxFWz9/mT9MwgqxfDbQK9eZ8PARHRbBmQLwwL5ICRDI25mutc8NMCT3
GCeFDa7LVtjn5tkxO4AqWeDr5sFKP1Mvr2tccL4byHpsSCI3EKqXSgJwVoK+IeMk
5gu5YcoFzN9TLHfa6eXpsAmO46bldRr0ELIxirnCyaI0M3sMH3EPp0LJOdXX4UAy
JlRqzQ9/mnH3ft3PikCIvr+1FyM+0bYumn/XmduSzJ9i4FmAqo9mrFGiYVe/XEy3
K1JQFBO7WEU71RqdA1E8GXDoyeSmIlw67sG+DZ2Bb0gKTMD+mb+LpML9lfKAPoBW
7Sx+ow7+oDHEUDn+mWAedufxAC5vw2HfU9d/BmJ0u5HiAV47RzkUqUYm5SZRhSHU
WTgbXWGdVu/IZMMCU5JYKcC3naTotZ5NLA+/BOHaBoN9gaIq3RuYFMyFay+WZ6gZ
JubOz7TkcdkhtVJMWR2bXbaIdwxxCaRveqF168HY1+rxN9lrsAeLAKVt2I0r5Dzb
kB5cx/USMkVINV0i9OE8zguANacK7zGXzx8bRs4IBAGfBd2uJiY+Mv7FbswDcdXR
TNnG/gcU7pSGI52IATBz3okiSJ235zRgclm6q4HaGOMgt9OoYVcCIuNNBYJFyxKQ
Qc/xxrrkwIuRaq/1VVnqT2uVvHeu4ap6WqN+xbxb1hjUbGugGrhyeBQLqCI6d45M
+raoTaX2jwcVAFEQaxrAlYAiE4u7T8WmkH4YF/m6KvZ/5jMuoU138WERdFm7jspx
RtKY2jZCZKSv2p/vL0JVLLjHaYorVXnrEpjgSIC+UV5+ZFBb++v1NJiL4SokYnRX
mLuwqhxTH1r+kzX/nOi3ee2E9p9NKQkJSae5MLo5hjmDiW8zayuEllYdOQsfrTib
vcs1t1Oe9fA5i2ZdeQn7u02kLB6+ZxkD1YM/u8eFR16u7Fy4W7zUgupHvREN4KIp
sVnHKCLuJWT+fcJcXD10bqWVLgwFIb4nfadHFdtf63U/Zrhenjw6S9C165IbmcOb
0snvEAViTm8pUYbQFYFU4L+qtr/S/H0A8/ZZS+9MFaV3qALbhm20KpOODUcrHUuQ
CcA5mUdqJex/p/rSycBxNF73Ji1ldNHN8Ct40LgWIEMA8ejqFk9fFpUvxPnogDO8
30NcWr1u68QSXwt2Vng7MlAhV/WvsqjnCeBI4hDhE5eR/TJ7nRbwxym28Pg7Xe+7
jFyRA1pHRZBO8ORJr5FQk6kRcD+nUEl+KV3so8v9X1JUK+hqzIQei7w1p0dkOJLW
3xrNwQwN5R3Saa+DSKB3f8dv0d+N62+f5juW8q/yVgpBPj8f3fbyoC/kMTfHlWf+
clLUgNHlHqd2k4yQvHeYYmM+FyQu/2zBDYww6mOlim4XFyWaOmDwIInpr3fy0MIp
7dCGDz9vlHHGNpxtpAd/zMQ8xV34cCVCZCk1gimbqJb7C8lq7jetUfCgSJcVwnUs
yq0OHF7B4xoeGpNzzEH6ARUJy4Y+P5FvA3jpdgqzCw6JtnXNvw2KFzyZjcb80PMs
haCmEdKoSzVmAuvbDu6puzFGJr7llmtPIEmrTddSmkN7tjwzaLDNDWrxEAvfmwsW
TrVlhZ/JNo82SNGg/pNY/GUVMhkCaHqE805YM5blHTU+8ImBSeJ6WFG7EAPq17j3
EqrAMVT6Q6QpkgZWLLrwWuIVoTpNYQEGtSGETwpxG/X74dfRZuSSRfkelTFmumAp
DkdF5COSJM1u1lF46e7Ih1vpv8nhApQtdrmmdCBCY03IDCwD9h/lkUAZAU+Je8FT
M9qdA6SDY74a3llHzd5+M8P+Lx/33QMf5E5QhrkuzQTyggxiujvmz0gmALIIgcfX
L94WFzD9UwTbu2NKBjPjAa4eL2aD3QRwmyqIk5VDRaGxnlSvc1XymEoD9ZBR1lrx
ChqfG04OZCLF5WcIsK3Vb60vEKPCkjrkOyYvNqfUFF28AOoYcAGZwp0xd7WrGE4J
I4NS3te99o68lMiI4itW62Tkt0Y9sIKuniTMAaKQWoYJgDI5ogRtL2p4vbndHH8U
jEQ/SiwVI0WSsFgzEZQZJnkuBTFQHZK5Mg4IrnBbgZi/egQWHWXjcWqxFGB95Ru1
yrY+hLr5xB6LRUZDY6kVjbKlvZlVMsq9VXuN0HVzK9WUKZhleYPPm+N1gkvDbsJ1
5Jlhw5Va6bEBpOMV9+47QFmjyYjo3SHGozyVShZxvyt2l2/6YnfwS0hoKYWkz6r8
cYjBawcj0ng0xK/xYl6llUznBF1ExE2MWHDHT4qaxMFIWRa6V1KQiYJ5ofWLF1FD
SoBwxSIWPNSihhx4QcNahe3Zgho7sg6PGZyywU6EeEx5toh7mJSDMphbbPQsw78N
W10boN6+bYZP8fOl4e3Y2h+4vyiXn1L+nZ1LgLYgqStsvR6mORiH76NDw0IS3KaR
bhJkVEplKI3GVfa1Fw5BPgK/AhHreavxr8Ma6tsGmsjJtsUy7L1mpWRvqFHhRM8I
MGmhC9fmcGvBhcDAPp3VbQJQGJPy0uvd7JjdK3Mxwgbec7qHJuufouHfIv3cSa9W
Z/SgY6uWUI4phik4Kw6CPgzNeYqKDJ43RX2Dn9mukhZVKmuuKVVHgrchd7csinl2
IYU27hBKnr81GoCNiJsl8uVDLZMEyfFSAmwU/TX/IluaJWzIjYt7KzUJsxNfbUv1
lU3OmDIOjlydPu2lbdJS/iS0zP3LC1J4fq+3P7MZfjOpqDN4y5VMy3tm9OuzrEL8
B9auGLuakUWznTsqYGJFH0BT/zRof+bZp95cbFPUddduXy9pyspPy+yT9rasrnQh
TvEHCUvAYHmsw+lq3AuQKO32ng/5X3ux6h8K2pSY8SO6QUPe5sUCzwUBpukDYQn7
P15U5jwvx3f7FnMhfztSvXLhUmFc9PIaWo7I+9Jhx1bvsTmX6lwYd36/5LtgoJvt
12OOSt2gnKzw1mZiSQ60APFGDuIm5y0k+zGrBWLzZTWabn8U1/I/+8Q89mhgnDEt
1AIzaGPG9YY7y/ooREKg5eRwePA9hXe2+fXp5OY18A0EBVDElbCI/aLRZlfcT6iL
mN0Nmh+apenMabfTilbUkH6DRd6kO7JtaD+AXtadv8jEp4Z3mdGWqpWnoHDrDIo9
3HjZsREGc8VNNzgftrlOUkkBU12GJt58ze6zxFAAJQWUepE8sFo8c3Iur54eYELu
gD+9CUyVo6ByY8q6ZmgfR8H/TfXaRmmGiQTC6su0nvKhmnvfois9FDVkc0RE24t3
tTuO/au1RRSSRjLyy5c7THF9LqVysgxexMJOoONf63XOTIXQaJqzGifkh5zFcMWu
ywsui5pdE+tpFQtyORLPTtFkH6tU6SUXvrDxun2YPomo9qHWF1cpddOSC/QtddHx
mBxkzN4z9PviEgFCTmWcOvAcxlVYAZIAhLRu19wmad+jyBcfJLQL3l75+cKqfhl7
Fzfv+c8cY1EtiSGxmNctvwlsImf+GS9jK1v/tPXkvDrOymUtFzsU9CUspHd0D5IY
xAXO907VX0mVo8h9TFMnb9yxuy3+Aa+kjwjro0FtiSh5fNzvoHJMdlXsr5eonetN
wemJmg1qORdUXE/cMtScyd2P7mwBoIEr6lHfq5M7TazEwxQYrTmwEncHQqgbmjF4
VbwWhCHJghmKT4BpbMF+GIdVCd4LapGU1o7eWp6C4rQRmVXaDq20DIGXPpVj447l
v0j8XMLUO64uLrLJf409RM6blEQ6MxhQ77H7lJo9sUsNagd1XqZaeUiJrsE4psly
1/eeHMczvMb9s5ChEK1RJpiI7TAjFU6C3Poi2GWCSAcbDV3oQCw1x8W8M9fUPiqm
0XiROTc/0qgvZdBVJFtY4XBydmvMo/Nf/r2KRq1cTVylpYehPLa551B+tnLEN62s
+50HztBkdP4fPzrGA0gd/YRp5enkhTOi8EZlAzRVPORMg6hPb+paWMyLiN4rR8En
jtfDuFEM9h19JiqPaYth/1LmgovYG/mltQHV07ltIEPlXjhthUrcVMsTeXYNyCrM
3NzpaHWMOPPIgmMq0orRiC9OLYFkjasln7FBcbKPqxSVOWFixUs79a+7cHewM/g3
xpdGLx5xT5O0nbIIEmVGS6aUVDneS+NX88yCeKh5Gs/IRlgLfSNojigNoXRqL/cg
iRrLGxBWvK9KIc9SzdzWKtkucVdZNSZkXM4xeax0BAB6qNEus7xEXKzXzZxyh0yD
HDPhxiLg0Yvpxr9YHFpjOUQOU4yVO2ktu0Ewk+qyMadtMgOc6d3pbeVVXTzk2Ftc
R4yGf9jkseChs3E5i3GeTA+/hLfgJSnV0nNBFAbNpfm7n4IPnS9oY42UBvLJ+zTh
eCXW6acywVrhICLBrXDfRUE84ZNLIf8Y+Qbq97SSAEPDgF9aAICH+L3umIvv2BT6
hNB14fvn+zOMorIkU41pGYmXbUc5tiN+AAvW8sR3UMsBVWfCAP+LmdEL2Xn0brwY
Nchun4UBNgqpb1X6KhRC+00XmDXvaNkgwOZ53dk2eiDIkuJj2RFenAx4ebSJ9T7u
Stty4yd0RK7XMKTs/hbF+CB0it94btTxj99z3LvO8DJ5E+rZzOInlexncYgWztc2
MKQ692fOK0nKoc/g1AR1DiixavzcwxDOZ45NlKEFomnfi3sFbYSD98HQKt/GGUzt
m6xH+kd/0LDrwzTZaUWXj2RY0pcnG6Ef2L5b5rgCWNgrTmeIfjIDNnFhJ2ihlyvU
1xXVpLIJHZ4x4sKJpguN/WglQQfsLbKhRIIz00F0/rJAA3rk6X4wSch3GwkWhIaO
/gBuevntG7VCu1abHuUftsr8x8iQGd8PfB6wthQ1uNvOBbcBqpS2X6KpYbeiO18v
Wol+/4giKKQ2SQP8gT1U+Z4XjnmO0Jxs+AqoOB8J8Valw2soNR+hWiJuBAf8x7GM
ZMfkfZvWFlGdAXKg3Uf/HUVqvdoDKOJlVdDkPmP1tutNSjjjXjMGeZ4ZopvFgJO6
1pF6YZaWcliQ5ao3TRF06NpoIxk8TUYcVVUGPMpimaKvKUNFAT+KqXvH9AX+Iyds
f2q3FugIuAPlqJ1I73m7Hzg9hHitxAQcSellujEPxFqB72fyGzY8OBSGMoPPCkB6
f6LvZZdqoEC/6CcdZ0aY9YjFBxur5hFGICUseUgMGsgc6Kujz4X2ujKiFw5hpbkq
V8WSkmsMm5VitDbOLT0vb4Sa1UUksf+vlLhlfQ5Uw80IzpBzr7T9HuYAefgTyYPS
BAPKVq/6gPo8I3H1b54GBxOosaqsTSVCUySDzzeeGJFhiwq4nFV0S2GhoRnnI6Qx
TB6PLTT7TxVU88aotYcTn4qnDktZBhIdhKbO45N+hIMzUXyUqgORr87V76dblZob
dcn0K93cR/rdibG7lahNHfFWNVVuVRIjEZ1/7lB36eLcJdt/Xduhk6KZSQmsl5XD
tYSem8mXqlH9rMJVycz4TQtsW0O/k2DgpvhlhE1938C6ZMFZQbetEdiTVitiO7S6
+T3RX1QYVoePrsbgVeNwPA0kSE88BoX6D0CWXmHC8MYrYLVARmo2+kq4W6bsbEdX
jIIzH14uiPeWR1rNteLj0/Y1mTzPTG89Tb2jqYYsWx/5G4BQXHUbyYZP890yICyC
O9IJF+PkQc7H4BImh7RbkkEAgw/7eEPf5sM+yCf1HHrBi72/m+k2mOa5uI72n4vD
X6R5L8ZV0WO0PjduUZsNi1lR8ydNtQnlVaUmebdilUAw7VZwHn1Cfx+PxZ4bExMY
X5UxqMzZqzch3A0xRNj94uafgW4DMgbrjgBA/eKiZsZO4H/gD90cF2MIFUZs00w8
fZRiIt+rNdASvOgjBECvA0nRGq8/kX/xtuDMWoOnwIT6ZydLEGHYm/5bf/RtWLM1
cFWNJPG4MybtVWwOhxE5GtBVgd3xUJBHU+mnPUorai+eau2JTHQKnGpoAa0DV9tY
h/39L3agAaygJuxYEzzsg1oKcvoc5LMkWaEYJqcWFHoUnS3WE5tU7HhwcovpvaL2
FXYB/IPaPCthjttCPg7ekQVPsbIDrw89Oe/QTW7iBfB6Be9ThrlA3RxjFBreTLcU
TpzrDXtvBXaGc3pGZY1ocVgFwg/r2FAXedwOVKBjFbR7qYsRnP692/Vqc+YPlaNx
URMi1RDzH+VCKQGSowxY4GB3MF52dHeNrra5F/h2CxN0HsTXkAHjRQ5dsGi+5nbk
ecWbB3roXCSDJqaECR+BilRn5UD362HEDQtm+E/iAz21zSRFDyt+W2BuHPf31Ez3
6Ln9PpveRFJZBSnEn0ykWhrghczFGBAsSQ2hk6N3w5ISHQG6DNF0nb5s6N84nv1D
Eu9IQIqkxacgmcoFw7M2lq/eUFuzyRTjrmlii+sGBT6OTa8faz6mPRjCR+WgbNby
440PaUKUhjSbM/J8ooQJEEd2nBlAZHG8H6P1J74h36YacbAS4FFmUD+jkOXArOf+
wzCjnx9bC6Eh6T8bklkceF5RI0Fh8oBAj5YChyNSiFEb2sLK205wIInHIxDNmP9D
dJHkHTZ3jQYoU4svlpvlmcFh46cPkhlT6enOBCR+jxzmGTGX/1vck0zwIf0fmMM7
/KWfknBANlGNVuAJwpT1W0MpA65sAQau73QLib+en5zQwH1ksyU6S/ta1K/zN4vf
DEBcmUNzlRZ8jDpcmkKiIAU6YcEaA9Z6UsjaGEgy4rKSvadrV/0dZpLG8snXhGVz
K6sAqgg8rvPYNRTJy3Q8h84jSVTZA8y/A9AIIPQyL8M0rpbnHvE7EMavY7tGgtra
5Msi8jgD6YGJ30EPWLQvK9dgImdlD66u2rET1jMtqK7FXl2c/0W5rM1imvAu6Yu1
C32Dcqc8pDHZePXJ4dD/Jq5kqRazOL1GMpW/FKsHR8GO9wEzqnX95kAPss5nDxyE
SfXL5a2n80N8r6D4gp2xrSKLlR2r7tzECCCUg6RsDPp2Wlt5F67cdLbvpTyAq6P2
KLF4JR5EYgmEbsXLMITYP+afIfE3xifZRUqU4A8ZyqSPeRVOQ4KBwD8bXr3cubf1
XEPZV6PCnAYkgOvrKWKeGqcy9IrVo346DSqS63fXidk8imLimF6/UngZuYU6E1YJ
4Q1nJJyjw/ZpKsmkMpAMOTG7iJQmczDNonlx6ykUZF4ozi9MlPl7BNbBySKuxRcy
guH53St3P9wC4si0swjlldA/mOU1rmk8tQgrtCpqKVoxU/bYNSFwSgkA4shd6DQx
G9fK4tOwoUwX+y0pqSxVnv25xU7Ihx+BUVradLsV7YYpUyz/AIxiiw5TKbiOrhGL
c5rL5osQsPZvswTlRUwuW7o7+uGfYpdOnqnGAThieUOziQRwzN7HyBeqPi8Qkyzk
zEGQi3zEy34V4Jp8DPhD0OUVBBCgeAytJWQo2fF6/U5Wr4MfIwlwHjnuu2Qn95Ii
MHp01z9o6KVLXi/VxxNvRQ7IRuUOjhnMh3MbvEzcVKZAIReZqLPSFD9MdadTozNV
HaZcK9u7S5xTF346ACmPS9FUGW4G+OMM/BeB/duhUfmBsVe7ORWSbMqNRxWpqPQo
MLVKKZm37bspJ7rSc6BZSQO2SsGJl7CoSD1BKke5erWu00XpF+yUJf6am7v5Px6F
T5lz/Ciskjo665fjjBPk8vfBj74+RK2ukP0tyum6XjfGHREl6gfl2JeXe0Gk3RLA
fjpGlUzE12vcBphuUxGrCW7AOY5/ZI6kDYZh/2q1S3BWmbc5VVoob2gA2vwPTpwc
feYChPZg6Hvhg5wSVWAnUm14Ra7UgcmaJ7pFEz20cXKsOJ9ThNY+s/GqSpYkrEaz
9C3lRYIDENoeIAsJbEr4p1/+/LQfLzhtUf0nbmLdh9/VhRWbdP6S2synOKr7gb6Q
qulQm37RiWRVgrh8fSEJLtc96uU891JvCgGn6O/q8dYD62yup0xbwMgDi4sMDF7H
6AYoe13ccBOUQme8H1OgYhu73gk79zsVHiNr2XqVvR52R0+fG6Km1sE9aeeR/umv
JWwivQvqM3KMzHPpOfYLIoxnSNcxV/gq6UnbxP/hylNIBd48+96/gZ4LUE+6s/iE
Zkm2elCnKTJj9YAlbeMGkPQBeyKp84hUQCl8eVjIf8LAPwQl0LpTyEepDZI+S5ex
tABQVtghMYua9zXv/Ddmc3BgFaXBeBTP5AP6mw12wXzbX5leBgmCsNlUvo45o1T9
9xXE6HuYXjLoUdOPPMWqzB/zVZHBw+Dyr2bYUB9+HNn9Zrhnf+oMlmDdnnXXgSuE
yXNchUqWOPTCdE065rNBYP7ruXCAUjCTnPPtHrF/fqB31G4LDU9AFcxd6Hz7x5ak
kRfM5p5w47jHjYsBWYD47cyO9LRMLvAF89cdladD0m5Ou/LsHquSgdQX8Ynge8fU
x8nfbQh+NYfC+l8vqFPMsNZZOerb3w0DDES80c8TdufEA+OXY6WvOJqWg62zNbfQ
SP2R6UO2Rmlp71V6AKEsAgo/jkQva5N2w0W9XfxlZAkUD0/cBp4/CCARdjMwFuzB
SMBgH9Iy6I+7RJApUTwbY5hmE3uVUCl+8yxB08oDFla3ZLPeMLjGHtvrFYIIk7o5
NC085PoyIU8MX9gYgwEdtIIkV01aSvyrJtsdtb7EELq9UBxOnw6qCeig6MaBXdIA
AI3G9uLW+5BPHRz+Gyropid62vONKdSEZrBziwpoOh5j1KkSbuSGOyhX+3roq/+x
zoHm4ejWIgUiIQDpRg8NPCQ5eurd2uHIhveCznFR1BHAtYHv3jof0G1MA7zmF5AV
Zk8JcoCAGEKfhO5EDcBCYG6jXrHEC8ZKpfgEJ//DaYXa2r63RGF5Hxcp0o8JJBS2
BKdJERPWYegpiBwlkUu8iB+DVqTYQs1GAeyyE1RStzr7e8lmQy2JlRVsixYixAHQ
dFm2VQGL58J+dow9cIo6g5PCrT3z1gfz6+kKCPeQnytcTzt9RTTkNydBQg/q13r8
2nwvGB1ex7iR78bxjoeftFXIqF32KTKZR65mBB+WKklQrYSfh97ghyinBCZuFkpB
fdkxvIWBbT7S+Kj9WK5+chjPsvJ2CHs4VV0Mdwq80hxTVA/UHz/ERBgmUK5aUo41
jA9IFmBPwx7/Ct5JSPYM8uBlEeSDM80b+XvLeyaQJrqUopv6H2wKpmapxnSSwZTf
/tAYHDIZUgKHgfLk1OPYszTY4rH5qVzz2geN+1RZKEc7hYSBJZbJa6QSxV/Z+OKP
tjIMu65sSHB0El9N9vUw5W68SXPf/TC2KpFrNj/lGKyymIpBKHL0c56fmxgnz2AS
laOKT0UaN+V1kfV+yCCpRYZP5zMS/Yez1rFH2XysVIE2eDbK/SUZwVB29+IbJqvC
BS8vgZnAbAk8nXQWi6hncCUGMCvnJ0OJLFpoCx9+Gd1ztpyqEvWJ0RibJ9a1EHhQ
71IhEjr5oVEHUG+D2pVAkV3h+0G7QB9ip4zIwoBqZ65mM4ue64965Cr/g1eE/yqy
hlhZQNYBMrd9VNKG4nsug3fMpekozF/PgpVw2Y06L5FAL9D/uR6T6M+QHqTpSGsM
gjHwF51Vribu+8Crzef5rMZoBaILNLzbDP2PfjfdqhZdbLkXyW+i1VdQGU1/mrex
Gx1HtcwwBcL9lQOWa1VXFJqPxSFIlo9Zgc9SzfvK7eaEIMPxYiK1cz9CPUQ3mkzX
PsKPAfLi76sQ5Za2aLtEhI5/jQ0T77YGqt7/YrYNpORfKlhEhDd7fkD4JZBU/xUP
BS5KTqEaiNb6gJZuliwa2LR2Pah2IYomQs5/zPu9ozEMVKux8R3Z9CJjgRwfDBgl
jvbdqJsm60Sn4S/mNg5hS6Z+THCGxyyVA3igXJjsMCrTrwlkBo/VJJnz1+ZRl0VH
lDUK8nutTDsUu6Uq4KVYOqQbZJuBP4ACQ4XRtT32SOSdRiDLfuHP8cgm4NcHnu35
SuNiZLGEUalhcJoxq80rps83NAf4M+WL+c8L/sVw10yk4gO1FIdlV/V+HZDTqZuh
YYp6pGgzEi0fgp5SyAEsk71HzALfk4zcgYctdcR/s2UXOD0tdDX87qnPLtQO6Tx3
L+PlfYYLp5xjIGsmiyVjAL/O9eBQfidKjklaQ+XjOvwcP9NvK9x537hIDIGd4KlU
pzG7qfLFp9tFZTPdSHR1iMglhRk/48Aq4xylkf068f1xlDqFmW3Y/PwvnDXFLR8l
bfRxzAb4JlD0FpPO5orsb+fLh4XW0zBS439VbSv1qXZ2rHA6olT73qxI0MjfifOr
ebqjyANh++DAfkPkm6CJJvomUbWiY8wSArrpgA/f8aaAR3ll9xuAlF0nHHm77iau
9qZESHlUh3zhNh/qMl4m202aYrthjowhhDzb8ht8m9DpP0bp5DZ95+LpuWL1oWdj
iovYNxUtNhTRKIA7xcClYy/lK6TlRaRlvcuMRx1BPn4dy+Tf+uAItJ8fNQBrqus3
s3J8LwKt1mxjQ4aaN+589CMB6NHZyU/YVHonGrhwaqgtO1qtlYSUHqrTx+wcYx0M
5OFLP72D7S9Dve+aHg+aGELtUuiriY06fD6iS04wMc54DXY+ReHIFWEvDvJ+DdA/
7EJ0RCOkeZfRC6WMgJou12eaUKG1duKQVGnBQosYb3ANJjrt9SI0s5WICO4QSHx6
a0jBVCKWgWL0U6dvntSohPTctW0niwMEFdqw+fgmUUxH8VlG2PHvG8hoRhnpfRoK
QBlRnml0tMG4+rGreE9awOCQ1kzmQdnX+ZQ7Y1o1CmXlLvxmiW4ELTYV6aZxW/US
GVCWw1Gbvp29hPOiVk7HD2RLI1WzKHeQfcH/hULWvKRl42fHit0r/BqtcShxdt2m
YAqRmVFoEvRa6vq//7+rvNSRTbAuEchqFog/VNMI5BGCnlAzr+LYlnSB0zTI/L2b
r2nsbQHMjSenqPxeO4dH6efjwUwWsNQWFGDAS3R9UK/Oo3Vvc0v7L3kf5JebysZb
ttyt08n1pIm+eMh0mgxHX03YkyzBTe0IowQrzuQn/Z33NfgY9nI91orYYXtgzPT4
rnq6fDXx4OqMiQErW2Mg8fJzwgLEm7L0gG38xtQrSYYVjFkzxWV9/sT0CkwnDntN
Srjaa9xgLxNSOr3AKwra0k3tISPIkISsi/VgK9CqlqrV4iR585YasyYzBMmAyTHq
pUeYw8M5TnnIjfhCWG/l12jDRslSjUsjFNXI89L82SoOA3ulbyJAJRSkA8ccPSls
i+64/VgVWkCCUJgJOAWSIpW+7yp86qkW5O8tW0MYIHRDv7AYJ5tnUE6MDNROAD/S
Eqmxh6ssDxmRFB86/oig3/c+P7bTiw6h9a8mUuUpCBgbql3etx0IYZTbKEsSINe6
SBeNL0cHCMTmO9Za/xFfciFEntqBDom3xsclOcm3OLV4grvQ5MoUpzMOi2i24PWY
30B49nQHiASut8Z8U/XEUfel82LSEyxUN3CW9Y6lWl19/lRWKGnhBsC/bdUWIWEB
YVg8/3COKf981th2nGYroZSpMYiWV8YmHr8AliH3JpqkhiRHeFy81auntRkB6ina
sDgE6q2pnMyYBjKx+rgHUb0Hc/yJxHdL85aZj5NJ3flu7/hA+NvrvhYtKOP553St
n7Ff10rITBpZGrsSWgVU4FQhxuq2yaZIkKTtMJE/oi14PE3fOWTEzXyVnkGv6xkG
hqSaA8eTlwnIhm83ZHCqh3WpG0sT3R8bq4XMxwG7jZF+kP3CZob/ApIQZQYx3EBe
Ozkb+GvBa7fv8eyvzxbVfqpzU+F54rS9Qamo+w7JRjz45TRENzZGspRnNCRqD4Oi
5lCh1QkqStXBhmwIA7NWpavn/pbv2leHb9gWDK35crPkdL/tSCYybs478nKAjz49
XdWnzWVDP4KkAytVXi7xbx42P4SDZLDq9Up1Ru64znmVIKLAb5RFmux7rPRSgKP7
HVUmBeCX5reIiGnjHrul2C1Bsz70Vz2u/qCvdKbMDhiGfdqeI3rh5aBPL4uJMtyE
Ex8mfHPNhzTP872QgOCcxwY7gatcndURSw6B+D1zWpMvMpLmFRI5f7W62tHygAn5
etfstt6UkZP41JOF4qVEraJJzpzvZdbmP0cM5X5gPTTF3dG9860xKI4mLNtijJx9
jQIoXtwL6AwaaPOWYCgAiBAUP9m77AxjyVO2Jkl47qulc67HVEvJCvtv9zSHFn98
dtk34e4XwMba9yA+GvekwuG5GKJmNx+iuOZCj+M7O85iH7Yirspo7G9JpTaSZfNz
7QcdBfOHNzmDsgB/aufumCwnd7lIPydJSgnJKsmXOemXQ29JgKb+8cUL6Eik+WbY
l31LHQx5Bej4hHQB7jx7DRbrGQds1hrJWsKMCt2qjJtnW9dCZsbWnd0l6C8R8A/A
hXGnctt9JJ7vt/TSFSOjxSdVwxvtswZCZEuepfDSX79XA9nGaBSs7LB+gIhvqbK4
tBQvqWFzRgm5jzXRix9185/Ujcu4aCAIfAm0Z04VmO7SfGaCstTfCiw4WrEPhEXS
BATEOyFw5cnSDHV9gp5MWBF8aw5JwyDZsmpj9n8jstWigC5v7nBjQdpx4TTWL4fP
xDovi8G9crPnQbRJuRqDRTh+e6Iy45oqMXdl2PqyN0ycXCGGLrFONxGlBX9f3+i0
A3EL5vnMEGv+0NnwwM/5bVgypfcvwjwLtWD4wAhtA7PKG2Glva/GoGWJPkS7d/r5
Ph8tmRGPfB3aG97CpG9EIe5vuviAJBaKP7ilIq2nlxQEAsjQ+h3CgFwYehXXy3yW
a1cznPMscmwikZBXQNeTEihWTk2Gd5n1a+XJZjsgHf2VT75pyCCTVkMXoDQ81qOJ
aNhm5oERbP63/3TfIREN9Nc113OGF/83XM4PDor6MNT4R2pEePaNV/z5F1GhXNo/
MFW1SmcdwG+ugkhAkQpKnOLarJCla48Wp5j6m7FdCqJ0iXpLHjqut+0c2prsvNCw
U6WEyOFB0niCNqWCxUIK9q/qnPvVy+Q1vtCOyzhFeh7XgaXAFAZ+ARargqYKgVQ1
kr/SqO6Vazytj4NOCcgWyTwuvx+Fxa+0/VKFdi8XDdozaoH5lZskhBMHXCYTTMA/
tPZco8jzLUe2DvY83y8F3i9wwFIJE8ycuNS49nRWVPUABuyqVCnoTaEGgXUDzagm
PZrpjq7qPXNHSa5VByKEezB8MmnMQ4hN4WsgCBOetFvraA4MFd+5pdeqBHM8OPVf
sluORZmlF1X9zzLqXASGZgoHjS2wpE4DrwjDZ3GvctuOVykQDVMrFsF/JSWY0ods
2YAN0B3X4KX+jO2ZuSo1rxtqMsZxpgpWwjFAZp3kcqdpniwBE6dNpyitjP9lsJHg
30fYnm6IR5ATu+AmA/18OOTlwBNXTT6GJPpYc7CwJxhOpAhVjE+4j9ZhLifvXKyk
9vB9/KwCzFoalZpVVwmG4JlbkQk7S+2bMBkM/Vt3DZwl5Iv6XFX2FFspfhCrbS4A
Js2axNQM1iZBBNgze+VS7q15RX5ATdLWqJfrXyXMQSSqcgZEMnPGjYq3im3HWCim
ya763bdkZQHjUOdpN3duH8q4U/lua39CG/8WJlx8izD7DOtuTybaU9G9VckBFqks
t23RO1mg57slL3sr7uKe1PvAjxaj83t9ZVvLq7rBCHs3cjFGheFPR5vGN2EMO6ut
C69BYadePBz6LaJgdM0Y7zqN/EEBLvQEwQ2Q+WTD7hZaxij4JmN1NiTKj0vjcTKt
YaakBWpSw58FFA6guR3UOboJVhjO2feXo2wDHzIz9sEneSyVoLNzCRfKCGSpmu4V
t2G4TkayhaCGRdbuQWRmO4TVlpoCtO4LjPS6ipobxFzwEl51lVlARfnkn8CX3grh
lGKn+aytkg+F57YeP9BqTw93Ia5yBQ/6yf45jdE7Tqntpiwai93BLqRwIeAq4dmC
z4X/PAJ65DN/dPF1XPoMZbnuCi7Xt8DDsSZVhZXwSoEvVJaHn5WHoZVVLMRM4njD
Dor7MXqgGK9Qag+R5XRdua25oRyxctyFD671eFKkOrBGMPjaHaNsLBlF942E7tnm
VbI/idD4MVZ/ZjYUo+kOluMEjhMPm76OHh8Gmxbp+qZtvEPtAH0A9Xwm2KzUEekS
0sP7r5+f9aDumERKraLYGJbxrwYEU/kiI3orNws/RGHBKAPibtrWlbYV5Cq4rkiI
1C4faUE40uSc34MvOodFYpvqXcCevbSuheYIZ4EwG3mYRWu/OC0Qcwux8aBdkRxO
qb0IBzjM+ZrMuksFIBSRfHoT03H9/OSgH9akoZ3qt7+fIBPgKQQjTHVFb/+5KwYp
utUA8U/S6DOwA9TQR7ZPeTIya41wZs8SIAVElkVKAGvL4BthzXyzcXtBZrbHYb7N
WHVXE7Fen81S26yTcemedX1i5SA7PVIyGYEa2UGHqdrGMBSYt4Iw1okqCVN2OfMa
4PzpG7w8OejTvTXAysB09JAfU1wPztckCtAWzmbt24p88ELtaRKg2fDlnY1sIMRN
u8IGVIznx0t7PBMzetYNvxzxilxUHHTqBPebY0yiNVUVpgGuvmbR4z5mUNRqw/5y
Mw8eOcc0a09N/qthEHkWVWKxm8LuVbBtgC7KVkvZbKxq8z7pEjyo2iYu4ImZkkNZ
DJjuLO0Dv6q3o0boh368JokZsm/w9Kk3gxmfe/6s/500nOY9fVBD6ftlCII6VWTp
SHQRQdfga7S2LgI4F9qq61gbaH99uIJuFFI7DICbXRqJuGCIf+r7Gy+ZTnpugoXO
Mm5x6fk4jNAQVcPQL4J/5g4GAx9PH/YV/cQr6rFUcayPyssgrqbNExaye78RJDgT
54B1pv0Jk49pvrv2JdLh4Rb2lpIX1WJ+CwQ7TFQszPBt6MwDfhjNnfTevLehA/7G
2Z73AJ62QDvNnf8sesxqYG8gbxYCT2Wp/97cFghGrP6+e5jAyGenDfCCJDQYngQ4
4SJyC+QLd4S4VdpO44/rz9R6GitssRgRDKneuCIrkhnIWjl25qwGdiNbcZP4iMYO
HY6b3GtI1hBmClWIwf1rC4I0unMtucKC/uKYxFke9Y4C9mTNT9RE52f6f6z7jmdZ
i5zoski6m6SvS0nbG/5WGGHdXWuJY5uzKZFO3rw0Bl+1RrTDqJsFfvPlG74EycH/
uS3u+ftnkDgRzMPv/N/Q3NHq+WdrmnZoUWktToENx3Kqv6L7k/idEHTCmQavl5nn
iEdbAQJ3DRZiUMiNJhdUYRCkcxYhwnKrfZe2F7uZfF1+61HDZIsymxmu2ZkhR+LX
BOuin1G5xjbn0JlcZyGNSVFLLe94JkBqApHQ1bcCQfGfjS1DC0YHf2murpGAYNG/
6YOWXOvE1hWcillXz0CT6Si0btQGFPweWi3o2yP5VKCF7lcRqV3nt5nI2Q/lV9D4
4/XfZ2PEVoJ4L3N0WZWceWYbZBQQ672JxyTsg/4McTyUNEt7LKdUySZhyC98FH3J
0g1+sHkU6mFFkQE+qRkRh4UHMbwFewhMK+ljZBavTjlaW+ea3eFzAvOWG8Uop5k7
fAf+8v3VcJ2XNKxb7BqgSx/2kXUeNMdl2pblm+phdAv2NTy0gisvzMlvXc5jr/Lx
fDW/PguI5//aYpE3ZvkffeSVvI6Y/9uElIIPblA9dNXDH9nACroEpGXgQYc+2o0S
PafJmJBD1EK0GMbUasUSdzm4FuMXtj5HyGzEoe3dbB8bPv+PpmU8GRUhtQx5yz03
WFNOYD4DRF+vGrdz5gWwxLfR5zpwyFcRVOh3flk6weKDV50ENUEDngx2XUA7Djf1
aViHU/mffkZBYkOoIMuVUBlrCGidsWWGIvrapvwRnLPZvW52SQAu9I5jxaf+kkTr
ZFmo8qmSxZ8+RK4iBnRUbcibOuTVuVp8omTp9p9ZdL3+SqXXNG4BUk5f2tT4iATj
Fo41A0/ZDar0yZnHv+VwFio7GA8iLt8xYZCw5qKmaNibU5+2Zz5C0duXww5bdC18
/TkQFieAutx/PMLvL+HbOg50CvTETeWl3QqG3Ab/C3TCDEaVXHHV7aYNskbNlujE
7JUQtfFPWwUfNhG14iisIbRQx5aQlqVrN2qIU4yZCQ/jDPStlqJhfNJKbGloDJY+
qTksHl/gCJ8BbApfHv5QgPjE+V8fI2UTWp8sFwhZfQt8icRvfWYYhObNF+z3YUf6
jdz8Gk61JY8JxzKMYE7UtZGGzdKd+mPz3El3uQGEMS9F8MrWEY5BRfb8kiL/SAzC
KAhP1N+3RM8c6a0OPe+yCYJMOB8nL639INFGUO/Ma3bMI02kxpT2gCS68UgzlMqs
ElbZ+R/OgCaf1+ZwuB1sdwRpVFgXPs/bPrAFKtMNh6wB12YJYS0JKPEpkHFt2xVZ
G8a23eGGJNkqzofmhyIhstfMa6IYod7a1g/xc+mzfpg17SGjNM+uH03D7xV61UAZ
E7qk3Nkex4egS5pks2KiS5EZxxjw8yAPR7R64C1lr0QrgaAevV4dIhnnIxyO6eT1
LuxQkKkQj3UGRyXGm3SPXSRZxVvOVq8n8wW6zJluZTn4IplAM+9bDFCwZaQSxbjD
bCaeuvp6Gg+0ihDhFIGelUuIi1UFxULZZ+CYYDQZX00tvlaJVBPR1XvcrIP8bR0s
lsAmG9UeYNSfMOkar13PNucxiNXzwBzksKJSbwR4eBBs92OxY1r+1Kr23IX85SOS
rcveQAiqaVfaoNxjq56LBrL3vIBBvgvqT0+FUv2i2pp6RAc9XfMR9zjB4bypwa7R
zdETYPdheetI/pnbNKDmxLGqSttzQL6+xrFWGRFVRQZGnuGR9saWTvnuM72CaY7R
4WExCbRisnQnSALdc74tlHRSTpLUPHBXtP1Stq1KWa23UL6e8bYxSpHp1iEkHslC
yhB9mS/ESq5Hw5QxXU5cM9oySqIxahIsIpO53zRVZesyz62CcGjpeNvIs8wgUvZL
0cvUdGRbGYCrZt22uYLYvzJmH7W7jl+CgbYguXMw5mFXogzUq6EP5KgjgAtN4lAZ
KfMZncG9psbWVXj775L+sq31Slfh3LTFBc+44QN5R5M+Yfk+NpIWRi+6xgjBScaJ
PWUXNNp3Y+iSIZikLp+gVVStly5ocJXEwP786BZ09WjL1lA+zhx+EvB7Zr0q5UTt
biXvLwPQdelc83UL7jQprII3+jDTAL1w2KUvKK3HXtLZYpm/ONZgZUzGqkyFGSsJ
5zPx+OHno0IQzCRlx6MCHyCvrJb1dL159QblMs3cwooZIYCqIFXH5YnrA/UR7EN7
fPlG0oCUr6nd0zM4jgnTgYKf8AGD2AqO0lfBwWSlrSy7+z8kcl3h48bJzoNKXm7c
7zMSCcwr6mgmagdE+ejHK+KQEH9L8MG32RH2JfNxxm1+ridM3E5iyhjalD+jJ158
DtnN/bPhedBGXJO+3UV0JvQgxZ+4nBVVD0RinOhBKRK3Xl4WLKTATVMz5Yvo5StJ
XlZ6YUhdexKHcOSGV97wp6awATAZbVfXc+qyRSBadM+ScaQqw5+qlDntSoo3SM6V
FqSapAgvNPi7FsAZhZHDrn8Pa8J+K9W6yZ+ea6+RxJ9bzVJUGh/xTBtR/4PLSsTd
64pJX/1vGdW2qwDz7CMlGCCcrrU7zJdbNdjmVZ4jAKy4zJYoJzf76cw+tTVF2y18
ReZGlz1V44j8aN24MTxPpSR0UU0AAoL2QCOI/9MfnYrFEjUPH9te1MLoPkQtPtm5
IdBiUxK4an2kk296BdMSWtU8tWuUYok8+3Oarq3O3OqXYK4/RHKnx1KfydpLMfnu
2fh/Zlyu94GLjZNH6ToiQ9XR8qdZnhB2HiFYEkLXhdcu4gdfupKcx9RB0RqO8ONC
KsN4lr3o6A7ph3fbl/O8oW87Ymq8oA2LHvASZiLWxcX/NHMrE8Wh2eUcf50bR+Ft
fHnx54KSCBCk8H9rZDph76qkGxWr9fumuhXgMNTs2Y/wK7M2Fz8aoxKmMDFvWcuR
LYGdnNkTLNRDR/p27Cw1IZMUGazDeiP00DX15v6a8DfuD1eofNBzwUFXY51nNDZw
BxQ4pm2Tm9WfDLWqr4JNngSq2Sb1/7QOPyihKiCSHCc9K2iesHwxdUdR9mk549C7
i5lsEIX55zY3bUDsLF7RnJF3QaRRtc6OG0EwXwi9eA84Kk2Ifn/e+cTT0YuDt5Po
SouMaERC4zpA+/plu1+PFSfKaJhRYKVLtHe5t+f9XPepJ1Zr7CuEZ96nW/1Goy4C
BM5ZDecCN/QlXTujqU887S/5LC7XARLEQqKOboSfzePjWT50FgoIj/+QuPbLxcD8
2EAI97S8ezq1+27Dq4Twtg6NiVp0dCv3agq2j0lTdtxj4rr8bUgkHQcFU/w7oZrO
nIhpPs7a+gQTqwgK+43mypRI/0ZMEJBT270WisQyYqIGD8TGLhiZoh1TqtlvYkuT
emvHUMitBmT6oFbX00Gho7k4UpuLqnNKK7gx7GO8rknDmJ3gWInwAupWAbxBAJmK
SNiTjqiCkTPvtkRemdRLDm/0CkL6DRgSBZ+bdT7Bxn695W9cJDZQolAORAfLKGYR
t8fj6tb6v+8GXZyR0Q9siQB2NeHfoLZrjvsvv3RF2j5kSehbzw9gTepdgomeNiRJ
C5DwxfgVMv46Q4FFHR5KWw7c2ph1JWyyGSrDMV9JQlvD8+14mRNHUHmqtpHhMdZq
z6h+zjtKUUFXFhzSW+mgz3FbpD4scQPEHFwGSNOH+JY7hDkaFoT8YopM3CAIE1wC
xbkSv+tcy9UVGBqAguQDP0xiyGDuVFtoGHbcDu/4VrvaXgyaozTRJta6JK8P/Xnf
FlPBIKYGTQkRDUhJYBaLy4qpbidxE1Wz5MQ6fP3n1YMBf8bVstPq7/gwd4kyzfSK
1JlKyC9FnAf7Dk31x6424rZdunjAKQPiDyz48oO0evMTUW2ra4jIYnzY1yIi2tV1
U0XO99vBiNVH8DA1FuEiLPlmy1ItTVSavkqx1JJr4aZ86TJsPj6SX4lUNRYZnu5/
WU4B83aJsjR30M5xMJP4EJallsGxZ4U+mIHdtzm1tssYGtG0H9kQdTP3F4wGxk6E
pK5XUtZ+DJoqI2UyZ17/baly3OkGyEo5klGQJHLC9ifBUsMLmbyodD95wwb+bTb0
I5ishFGb2XVsQlrYJX5KB0VlAAJZF93I+j/oc4QsiSuHQ49aBrYivfjgiu2wkH6c
rAILFFfV36f9bkl1MkEyyMgWFWIlOj+A3HA2Yf4aGdyI2YYRisFoLiSCsBNzVzY3
zS8ltdfkIVfcwS3zjs7dweON5kJ17Kxm72C/PYQAmD6kfNiXOl9LbYxAmRm0moKp
9H3VnTyGmOnfy9MAnK8XMiI3H+HmWWqmKgdmAhZZttXJm/m60B+4joE0r2tzGj/k
Cl9hJcavBoDAuA2YM96nWuZo2Pqe9DQVjxJabIGuqg1D+dwCcPPBkCszCNLO5FpW
fMoBBbktDZlZHKP/13gw6xeODpTkigRJ/VsffPWAOmr8tdYbm2FUgVzCUvN6q93c
j/kK5AODJVxR8Nbkp0ZhbLjbsr/c9vj75HVyzMX51WbevGAK7mR1u93DcrtS94Br
9CVtKWP5KNyXpY9WZnNF6XZbdLGueUxsFkRZ2tw9HxOnY5gdXZVje9kXnCxjuX1B
I1FSioShmPF99PslyCXlgAwcw/H9QhvJ+bkcXp6RrRGFL+kXFeJ35FNSlKx6eztV
bH/jP8OhtvrRopyPfRF+AoebFnS0V5lZa9wrzrg86SH7l8zcTc7oIPcua4h/KKta
OZrXPG9y1WP5yyxYRDB6jAuAi99wyowdPs/3Avng0qqWV0bQAP+zEW9COU5YzWSt
PLUI8bdUh+B5PbreOdh75rn8wM8eq1us9YuqgZR9csK3R/IV5BBVok0A554OAS7D
fur5TXPlel+04DCTV5RpoOuymqM6+v1qAOs25Xy1Yb6btQAieRMIijBCXy8ubd3a
ElF4bzbRM9MrIb8zB7P8c1IkxW7DEHmcJKE7Zstiu66ll3zm66cP0wc1bxxEE3qZ
EsgMTO0TzsfifU9AIKZjiXaX0xnx8g7F/4C3aQzHckgTpUTRMK5FzQRd3IcJ+RZi
B9I0hjNVlfQZ59eVUitU0xfn92KMf78taBJLIVD2H3z4Nfs3AW354WriBkJtrE+F
Ke4MZIiE/o971atQyzpamrmUOR2ggMlBaE4m0z+7ZqbbsO1sjPH8UTKFPpDALm0e
vnE5lmJZsreIo+9nB2kxHSbJumeCUeuOOMK6W7Aza8CwOx1eZaWv0kMPoC9gJMo/
ojMqWkzSJTIxQ/XMilKlDXLXBGIqytwZ7ZFKSjwn2TXO7zc6ZRFFlRkfuAEvhPsE
iyLWOSqHDsPD63gbk0CmCiWHWb5OSoYhPMRGK8HZgZMpc+8dC+CsXX1wKen4YYBE
9YUgMsPBvaAreILadLtWeC0w1dv48kK8Q1MzxAykE5R5lF1APe67PSv2mPIh3Jph
KZqOqdmS/jACij61SKXAeHiG/Gb2y1INKIOi7WGfB+RdsiZmjOQrW1Sk7vfGOCbM
qdSbtAXi/AlwhG4NYB+mvzQXUXk3Gk3S3+wJw8eni2nmW7l3AvrW4q0MSWshdn1Z
NZmYseJn2LN0uy/AA7DQaanY9gIKwOsNFPUPZEXSntznedps+L0QKMV2ct9rtjp0
7hM5TPeGb9j37sIm41oj75U+qHdZm1O2FRB/5FInCvdKm5YrjCQQYcGCyejQR//P
OJRFKznrYgkZHV3GuxQOxlqlP0f5Xb8kcY3+CKFACQRIZXsAhM0XVDW7GDMg47Cq
fG2ms2eLEX43NeRfL6pBAtkw36XZnSQtPKmwwmvlKfPaCXugwpzSyEwNJCOpW0zb
kq4HXmc1MHkkO19dJJ9ZaDBGVA0PhUKaLz9ls9FySJjrnj6Rg4EzDrQHHdV4nu4A
6DcGAez1uTxe7jgmcZA+ftBc6vXU3zrpVcaxRrE5SDQs1kspbzK7fT/d2tJ3HEWv
sEfc6vlEC95kNe9LbVPV6iJAV2Yhw7rjs0+Q3MYosTX8pq1x6PduClEoQpnUk4hb
XaGdXI6aEq3M7UPjMKVQKf2strBrWcyFZ/y9eRlFXTGlWbphv5PDj32bU4AbFRkS
SwbMH9tnWNju56Rq7EuqlgkmRyfCU4oDAsT0WMLwzKJz7a4pIvwGj2KM1BMpQUjf
Ts4OUxLsBzS4jIbXIIWgvl4ZlTcnGC1GRUI0VIPsPKGIHp36+GhOLxlLnJvLhAND
19lvhXTVsdfMSQZFBmzQ93+NZNe9sNFTebNi+kYYIyL08T9ZPXo4k4uHVWgSgoyo
tsbz9B37i9ctzcLMW5y2i7s2mpfsYkoPCgaqrluDDg16kB63VHC4gkny6EqJ22DU
+G84KQzd3jSVQQ4ETEEO4rUjcbTSsOWZ/g0Dd5lkCaDKGZfqqK5/gS/LPS9YxfHL
WyojtKFiOJboacLSg838HylaNt5j1/VAUtXIPVNz2pcS1fMaYxd9TwhGDAGvhLbd
g+2Nzg/hig+AI8BHUhTo/7JJbWCtFGRiTYxfbAip73T2TpM8SDS6KwpfOz1eY5GK
e0VHb7VfZhhgdOXPgFunWs6BaaHnz+GHU0XLKW2CnfQFScx+1iecrm+g0frCo/7B
NPeyXBS5i0o6VJnrkIp0xn6CylTXDvM6g0zHkSNgv8VBo6oXlDy3Rvc7nYZIt9Ns
UdgIAR+ZcLaceHY9p2W5/GmJ8sskU3JAF0Qv6jvgTsdU8xkEGdtSadmxS/sPjWmS
PYhHNqEtU2GNwVUBKe2P6x23gCewI0aQqf0qTMRBedvm1d9xYa/YeFBkpDqi6nHx
Hg634ZhieX5B/VnBG3V+PWEVQ/8VtaSTvL/7IXBiBlyWHARs/EtS6Gejo90vTzHK
Rm6/ysBIGVn7suAKWdDYJb2ARjJKH5mMJ+rIPwEjb6oYEithe//HKyKiPxn6ldaq
k7QvetyWFo8Z+sQWxXCI+Ylq8Msr5HDbVOHOQUwK7o5ELVYxwbCMvVuooVsDDMC3
E+IlslzOdposXNlKX1SLLAt5sMq9bL4cCgLqxyNu2YHYtDVcvC95hNE0jABAH+rs
6v+7CIDGvw2TTse1mClD+un0j01RU9RX2menswcL2n7v6gAQjnEtlhU+5mfivM+f
Vi7m2OcDCnAgqunPVYauCRtr6btsBGAs7xOad/84X4ELdL4tbFGjSPMorwMbjpie
dGuMqgR5KK8E+CG6d4gYDetiin+xFOjLklM65jRxw2MxoWfL1LHXVJQJCmO1pRcK
NFEXCqFOPGnI+hCjbA9IZy7wa4MTY6ulAy4kpBInd9JvANcbyTjhaxZcCYzMqV6O
2PZueSw8eAOjuKDa+CdIvbPvs5TgaTT/NrQ+Ivu1u5YpQHFvL5kD+PGqmvpGCnux
3/0ai9X8ahPBaHs3aNU0liuS4NVUnzEyiYiccRV8D4B8Q6pZ/D1OYncmwPvmoJ5o
0s8TFJe26DTk7tBV6D4HatIKDR7x64rVPomtsw/9EKv6BtMFkLGQur7EeGuweazZ
pk6VzffCFHXXQv9jlp2yBfkmdi0oHK1ZjR8I4ZkVcddas9du6fTMY1XSYUjn0yCJ
R+GwaL39vvat4Z/AeSBFyUDRoNEP0KRvUJ5QiK78CuqiWZOAcWDYcEvU2sPMX3by
mrGmEyVRV8T85qRF5yN1ehJA4RC/oHkUVCXDFQey9iIDIb8fuyQlNmdsAwVpcKWn
hRsJr/7/ZXvhTk1nz0oubkpd09L39wJhXqBDnsC2ydZ6TvAKjxrye55ZolAGJqZZ
3+WUBQMzOJuIcKXlLb3TwE237poT6F76s5tn3W8EtnWJec9kXlUJCxrlvVJnJUq9
JGov1DMsQPodPIWoGPuLEc31GGRWhqBTqFYuuRnP/lawQfWxGT4u/muGSN33m9MK
hMuhYDb8aftETJx4IgXXQlBdHtqaYuWblM3NhexLVg+ZzSugUZRiwG+nRsk+fFMQ
3MYAwq4lLhZdLCTp6Du1Y7F6R0zO6J2vjxMJKZQAvKI6UhpVNY26bFntlVahTGT/
npX8rcd79/OB9lxXUxZQviOJP8mo+VmL3/sJGhWRs6w/+ZQ/gpKGPOYIlLVgi9kI
1z8jxsNfPSeDlweGKALsf/x8oUgrskT/39b70913R4DxmKGxtwgIJg675PVb2lE5
Y+LY5pc+KB+BSJmSxWNtwA3FeW4x/eCPW9cFEDbXgkWYw/3iIJ2YhPu/s3JSAdaY
cGvOyBhasRiqEcs2MAtA5OaWCd8pckuvnRAOPvqmycf4LO0d+29WXeSZ/Sd8PXsD
hj9gDeb9O1u6Kp3H1mJ4+TOon49CLHPY5VQ1W5HCv9zckPUadZSWb4ZNAPYKD5lD
+ws7SHxvoEC7UBQKSTcMSmxf8LebbItlSFFtGjJNnvETo25YmgYz7bihnvkTMWYc
YXugp1yfVRkz6pUTeg0wUgwtyV5CDhRPGlH9TzgFbBCYmUlygDtablvpT/jCyHbr
wmyv8Y5UZERyOpGE/L1OlyLIIyOXWBqdMRNHUX7REnT3mg2J0GpAYWTVJ7wRMdTt
V2u1dSTBmsJc1PjzDFjiQ4S2d/42LbcvWGdatR+Ax+CxH2Ey8C3JAfb+68Yn4rmm
NXvm2b+O4GXgimDAY/SFQFTi7rYK9IV+gziYdIbQF4z9yD8zXXorZcYGhYtzkTQ9
QlkRuEQg1lbL4ggMTRFsAgXLplqfGpEuHKIv7Z2vE1LDl/+WDO+uLYejvx8wuqTK
D0V/nLUPqlVftM/mJMAcVMihgrT97aMBh6x0NUHhIk9U4LVUQ40e81o0DFkTnej9
qM+u2EfqCSlAkLtTMiGpaVioIzXUUffcWBBZ3tu5oFBLYd6eiNP9/4QB+mMGuKfQ
fmpY3mrlNQXEx2T9kaXLEo1KF7/wzQB5EfZEGhN7zm6gYsf7Is/wPcJW0H5cd+/y
LK8MpnlVHz71GZwJaVbpomO13DDdMrxglkmU6OPsqC0/RE/5dziMYdZ5cdxUIVT8
lLE+Tj4WP0WPSLn1wBGXUSjhdvSLU8qybC7Em/QgogU3wghZ/ADtKk1riAAF517R
Xuu6vGXkMqoo1BV05dH0ezqFiYM1731m1v1Qaf2Kvs4VEncF+PBIvw6ee1g2cXPW
OGXJVLjdU4YRV73D/pjWpkugf9jsFuPHW8iAtzJkVwo7zKheXE+e5ZEO+tbQLXpJ
A2mdbiC1/opJiAtqj8JKLZhKNg5U9lNDOuZoMJd9E2CEjPKbz8Nt0nwHucPna/SJ
sQbgP4wZfSqXJ+c7bUusFnDcILsag0tOtgMzjkBocxmOoVQ+Z5nsyMtR9nePEjtu
Yvjldlt4J05277oinPfTxh6kyqjXDBqjQSdOBI6MAKOLi7kd5wZ2eBhszeCNOrsK
5yP3vQzp91rpH37SYhGTh4eg9syJ90KlRbq1yQa0XfGaGK1JDTUkKOoU8TdGHAS5
cKxeZKtOLawQvHOeCP9pWHdohUqaWzxuvWFlbgpSZrNwNQl5/Orhk0fi/ja2hqY2
nNnleshX6uPdLPMIqS/AupZ71oKicy9BQwjUtqHCE51RCDRYdeh5Ja5kllEkju4b
os22q8Njt4ucFPHzcTWabp6IjBvje9Tv7r8Ukwbusi8XeSbAS5VeDUFX0MtPYobK
gL4ciKuLNczcJ4Xmyb+68xxg4j80Er2vMIKYg2rrzzVT+UEAYx4fpHPXGphFGDjl
7G1+PsayxrosHR0FkZFA9BGwlghD/GLiVxv5Ix98WMPHsHcODgMbdHen8LkTvIjM
Xugnth2lxJr8IzdgJHxQCneYsuivpLcmbWV6UQRk9/aB/T6kmLH5VrsLL0ydx/Vs
C82RMCsm6EvjIfvlSxERlrrBH0ZzrUYo7nj7OCVXGO/aVrDoUekmR36iesEvRJRF
98TT+PCUrCEexAg0lm2eJTSUlIkwjyV7aPM4avP2XqwEIc8rhFSCPz/0CZQN8xYk
6rmEysHq7qaR+ZVVS2It3tB/ZzaLiv6Nv07xZomUhcg8VtTHzideSEg8q3y9mUZr
0eunAHJGkc2mYkvaEGU07X0Gm4a4zuJs96nS8OfqV9pqlxbT91cwh14JG0LB9UPQ
Auek1oH84k70OtfvwlDtaTTjuZk/KDzHwnYQaWEx0HexdMw7eINCovgoC3eqMSrx
cfFpjdxcSVq8xBowzQ3VNXGa0WZVlGlvlFo9hjdfdZCw1v4718+0LJg0kEus8TdD
U8K6+xeuAmzqI+1v+rhCwgKIlfSa+lh4oibZOs/TaL17sklvAnnoVH/LjabEX+yp
eJtNlxfzkDhsiIyB7odzC/HYPKnudL6maUViiJtv0u6vNGvyJSq1gaGUb52d2A4n
NtWn219xyNd4RlY83urSjzj2AO6pcLZYCYmIboM/FbFWQMhXbQUVI8TiWe0a6UzM
4tP/lnJYP20gI6en+HtU1a8WTB4CzXlyk8RJQb4imIpeBJPoLyA4qwtGxc0pqPKq
Am1F3siZIG9K/1XysmMpldpjfqaXa0OgN6nIP5BUXiHim8BD2/iVj7upDw8xFWiy
UZkbLWQGTPSuyQxTfyp4GNsUJTr2wdk9Uc2s1Shzg3eoCoxo06HxZU/oTHvPVPdq
Cly5v9VJE5qWt00qNiHnu5YmVinGHb9z25Z+AzqOwlUd7It7+VM3BTv3eUYqjshq
gflW/AmXGVtbTWOicSrSe7kV8WWOOA+sRMCaUHpwnJL2euB2UvU5FZ09YOOCdXXi
BUskkC2OUOTh6WbSMc+mYCsbrmV27Ke1xQE5t5ONAscenIhHRZhvXF1VyAOHlRds
+fioDxw0k22IKXGacNC5llLTX2LrFZXU93fpIE2pSH6NRFJAcZKRBzpoBgwCjNtm
eP06KAHqlguBNaCfNhXEI3Oy4QzxR+btb9bK0vMNp8sjW9XneLO2UYIjBbJfY3cl
0Fuc+x9YDtmZi37pNEBUUV0BGxMl2NZCytziXPf+hmhM+xJ0Yoxj/I3JfBMlPyX7
yEGJsR6qaCdtr3zg36hiH8HKZ8ilfb38WFKMeyS81ErxOQGqxQixLf+9uuVlV3iH
0l8YRrNMrIW+095CsJCp5ZeOunZqFp4HzwBQ79xq6+giScLa/VEiuLNcCgyNkX14
mdhKg6TnXkq6sxLRvN2jgsXeAVmsJVV5HHMYZuaQfxJ9u8S0+Po9m5/oQaV7upxW
Nv3qWRXW/XSSxaKxLTZub6IH9jel9+ykzwGUh+tQS566Mltw7vY0kQPXnF/WmrwD
lrNmJeLWz+gup5IDyCUEwuE+OD9U6lFWLiI07GeSknLAXZFXAGp4FLIOSRXTxW4r
8GaOVA4XXOC6j+PFlhUoYBEUDGcb4mHMAP9pEiwRHJhXWlDSAHGhLUyi/cVKSIKM
QuAFLI7m72CifKRR1RHGTTQHHLSZGAogYl5mMumGqAixG8h7kgtGlmaCtA+9sj/o
seP73SJut/atPSHG3HKsY7/c+VRTZzTjnuq3UfOqq0OacOB4lqpFGK6R+LiXgyUq
k1jk5UWaIYWc5kYS6eUHHiYVRRB2HuqJp9Tcu3LZIpQ6IRmp0SnVH0A70fRFnc8S
nx4IbrRLF2rrK92bDizJdUuosta9rZBuMJPKTIArA1IOB3akTZurRVTInUxiofpI
GIbygRbsgq2Dyg7wK30y1IST2nTEBlXXzDHaWpRj31zvNaigLxcIbCukqQUGkIXD
2VzO0L6XzvTBytMNxOhOjmMx1pbZJKhZsJUQKP8drCA8yS4icWzCk8kwujBlPZSQ
uavReJqY/pqmJNiZRUQzfA6tDdJz7cgVCUmjkjSx7XDUt27rwakGG44gYNHIqH8B
fQlXHmSt4A14o8jNZzeCbCM8dj0xY5etzGpqU6TiwUZNZOeAb4XijKxBQs6Yb/p2
P2SKYYLsuAv9MQ4KYFsmE770HhVzta2dVDXU8oF0IIJy1UPq8EBUU8rShhmMrr93
Nmg0iBnqB3YuV5RpYKJETYkIo1JRJiBKdyFnqpwaLgfGYM3X4hS7wDECf/FFoZKZ
++3chw2MxwnuVCX2YMySR1Q1Sarsl6G9PZogSSgUF4+AeOTq9pFARmtoo6OPeH4X
6ZXp8NaBQMDFWl1y3VstA7OoHIQNlva3b3GGEHZNkFgH3GIgbpqqEebIjrCKY13j
c0bcR1MiEAO/J0dP5WGJ8iyw7mYex4H1G5HUu52mmAH+3EIb0t13pmxB4TXTUdjY
Fj6nrbiUae0ickhNMSQ4R0DPVwz05vVCn2ZlF04wtTzXyIDqY9hFtZrI58krv1Bl
+UvsRPovg5vmtQQdZGCAYL5RQYzODeOyANHqwBsNbimWJH/4LFsSnzPDNpV1P2JI
cg8lPqGPK8zB141riy8/eUfZizKdy2BQ6YXV9zY1VE/K/e8w5Kczjy70m2C6pcbe
L4v5QryIehkfo1YPyC10FkGUCasakpDpdcPr+EKt+a1RbBgfmPzVQSHoOw2rYDlB
q0VtmOxHyp+QaI3ky2IKbrx/59cWOhX2t7P4PoRCQ/29kpn0hkxqchlrHK3jYb8b
cupWw1mK2eT0C0Ywl2hTJhy11+zzkaWWq3GfMVOgW5zPKpkWFk+aIttw0Dt/3Jj1
jeQjzA3d3x2vUgDR85mVApvA/G0FRFc5G9+aSq7CHWuXClH2OdsCwZ6+aW11G55n
jqkwOHPafu+J21d5mjpfVEyWmlXkzCHqw5IZBBlBpgADDwibKU8TF80c0CS1rn9b
6ZBhW+gspUp4xoynhj5N5UJmk/AnEhfb1kOfHwrxFiI6azhlgxsN8nUlz3e9htAu
nU9s5sBB/bke0bgs1I6bMnOU+qhE2nFw881ZgKV2VHLryZakXbFkCuYHlEzVhwxX
ODpt5KxrW19qC19z6TD7HcKnhRJIKmNslvAvfURlXEFRJFPl/+E/fMZvI2eurnY6
rkMZpidbIOQNlpdyh4HUoNOk35YHPkoZzkifr++bDl/LpwJG+RUQc8seqtBCuz0D
XRBNZAFUB3ZKmN7Cd13mHQMtZMq0aUN+iht9Ctnu2A01FgBS/NTHbSja0dRvkw2/
tE+OlSGfp5Nz7RC5dYwlBEyaLr5Snjzdp9OEdDa2ZdEoNZnVI/dxEItVlE1Y4+l5
fWhbO3Ccu9I9Q8jGgvSGVGV0zWgxr0xtBL7Y6VA624+57HSOeDwUWe4uqBk6vxYY
KncYIgtqSqOt6C+IvQco6eyKVzCQ5f3Er6A2uyQMsMjkU0vMpPgZ37+a4lWSzK9V
lYB99o2Y1vzj8rU3FOuQayfGUxzri21jpfHlFtfN8XhbXTlFXb0kirE1dfVluJpI
In19yJxbbZt+ZbXXs17yIF9Ok6PkE3iYLxEoDFNfgRV2JUSxl73GX6cz8ipIYWX/
nW4tlVsgc7RnrK6glsgLsMvSRJCfSGwimp1dPYLdxKoCgeiipZ8LWhHDk0BRYySK
MNtVgvmN6at/LB08vKCis8EeQEFeI8iO5EjSIf+wR0Kj/0DpsVAN5O6GCI5ZMhpz
LD8uBwBI05M9koAf0mleho9C34YrLl3zPJShmZpKMErMhzEMjxXphgQh87FHEWlF
NIs22hp6yh+Gp2zaspat50HRehwj8IeMgqCOY4yyZsaQyMJqgcRcQxxUye2/M1Ko
YUmVS2sqdOM9M0jUppI4Dp4Mx3oLebKRkPbQhlyeJSnieZQFQYrA7O9c1i0Rrxvv
l3wRsBSgWcYEBZR3RGQevV8V9SG36Dl0rjesi4ztplIiLewfQA5A3Pb0aEmLsXEx
KdfuWi0xzYejNwjQ09BI+16raxLx+gT3vzYzNAta9bV0mYkfLYXQXTpDP/xQP2yc
ku8uuXQd8FYs4EfgJVUQNLBXfusPQ8gjggwlYkkSgDa3mLQRl4hc4O+oBQwPg3Af
K1J6CSllbCPjkUUEFw+FUfYc/Rm8+VH+V4a+I91OOshBtFrk49Q9QqEU481+Of3S
JOabUKflMa7BvDccOnqTPRNZTgQyBTiObP/qKqRhGZ7jhMxFfRxlkwhy5Rz8G0Nq
JFWe/yh2fBdjmY/LbFHgXo53XbOVPpPN/ds8oROfy6YC/xt9A/9IDHyN/S2RU80N
LkekNahJ27BF2b1BmxOVrQ+O1LBTx5bUjGXPtTXfLO7ARMuuJ6yIc+MUNZHMntcl
0Crsv5Nb4dYOkosXN7n9+3upOGskXa4GPRhw3IYFUClhsIQriyv6+VMRdTdYR1gI
pNp7O4oQ7egKRC3CNELwIWA0i15RPCBV8kT+q+lgLI5kXNPWxWTGXI/7iLthq2Ci
L+cQnuxmAaLpZ8DvWhnAjc4w7lNTkFVOAeIRM31NpHWDhfj4AtIOhnyKirwlOWyf
shnzBIGS4gZsW3OJl09Rnf+en2zANpW0qE1IWRZ2iusTKpO4WNBFWe1acGxGfrol
3Tqy1wch/UnFBeBdzqSJWM6z97zidkrqJ7/fzSJW/gyiln8FW6yyXeIhZTzMKQml
aqmZlZ2/c/UJmhetaKEFw5GX0c5XUBA/co7V17RFEocFtSTyLOuFo2Y8y2DGxCsY
7AqWAnN4tWTmFyai7PfQapzKDvizaxmGQPUuv2A8QLIYKgwbjUkYfqPAJwZv6uUs
/zoBH22aK8ksZ4xkNQjT/7/G9dbt0KKdWgL8qlJ3RXAbijk7RAXM7BjzC2gZOgii
ymTxkgNZMppkHWylppB4vcaFRvtX1EfCSLzckqezr9eJEF1Bq/s2+g5xCAqgNK/U
BB9dBeCv7efSM06/69i/xyTvUpd0H6p+5eeaoKWS0SwR2CYxxY6ycq4DQpvqSpeR
AMkau4b26NAQCFqDQhgHI4m/2vzB79cetQjz9jvu3SA06cr9F2+O5V2OiSa5k95L
D7/McUB1NAoA3Jc/AsKv/YcA1hteXZEynPPCwJzZ6QoxXyb9FU568399MVS2qhzt
9jPZyKwu+uhUwi2mHBUIXXIT3/15XuTmNBYfh0mo6DqFi2kbGadniWLbT3F0dmRt
JJcF6EErWLWoXKCC+6W9Uu46+MiqF758VuNQlCvRJrnQKzI4ETCtnqflcP8LUP4o
KPKntmIxmD+jmrVpaS2Az4XrdJxcY8xMXGxmKOIbrmDk/JJhiUsBkcXYHOiEkfoR
9mn0jZMqjN4WykQRp4lElVfevY3lfwLz5twhoRIRDXYkn85eL2IV7Jv+ko4mkyP9
TDJKw6Hmiku/6qvYs7Ih5kULj/y2jvClpJZfS/WSJiUlKeoylYCtxabOHlZLU9eZ
b6Edutpqtif/n0TDAS6F0Q/VZ/0nQ4zQJYGHouVOKdByJ3lKAPRWXtLkJ9EPfjDD
WA0bxiGlALOdugK9RowkZYeTVJdkHyCtWdtCPHEg8rS8EDeU6kbN9av3OBtbYS0K
MJTUYY4Qx+a/vZ5a0fImOES6Bnw1ldDqMzh4OUaBwQIxvRKQ9n3pC6XtCzb27oTz
clJeXaXjOCAduYR3178STyppKNG7xBMtC7S2sqDPUVZyidzD7LRDeHS5+LrY/pq2
I/461Gh4olKGckBbDb6FOLUbZcHnV72MUmFe8neqEQ6U4HWkCk41mHqHsKyTyt4I
OZGIqOnsZlnWANQb029+5jCQdY27DdReAjNGHTgGdUK3zkq1ql30oaaPh8NcJWVZ
GH7kMrluEdmDlEP28V1zGrHZ/zmmRQOU6kIzN8UHYo1JfqR0d+b+0rRjaPOTOHjg
aBVC6kRrft2V+5vwY/6RWO4NYU5jw1SHYoxgpghROX0aK1sSIsL7K+C9IxkvFexQ
B6qLqNGSBEgHeRiwOWV8ZQQ20AKQZyDBUNUl6l8AmM4fju+iEr0146vMAq2HUCHu
hQ6/Opj4mWQGVUR8C2iR8sVO9yLwnadODb7sDYaFbxYV6Y3mjH4EFP8t3WnOuBqV
Dhvy/+5VpePLncNP+jMyTlHdUIQEsq8qmKu3yI19lQ/N/ju7H0WwgqfJ9vuMHJsr
qw+kOGb1AuWIJKJnfc36Zkpvswwv3Qwk/6xgRp0kyf7ycY4MLvf8ohvEOSUBPJFc
fu7+q30oeg5mtuGZ6TLEjiQBDahi3QKLPXbcc7uYKJyo/zyQieF9JvHKNcDOPPxM
4woMZhIG7jwGi9p+uLgS52Qry/vGMmzzay9KM4MR0JQLx/8RfxQXgdHJKe2SjmjI
Z6J+RzszqaIDdpnOve6tpf1dbZBqPscX/42wXmh9JvN5EXPRse77Zu/psL7BjAZS
dooZZcORHOfBvnH54/Yuw/FGDPfiIN+PZ3x5VS2TjvJPLsASb3jqn1dQjRj4oIwt
IJrDcen2F9cMVi4CBJSjwTgWuk8hFKIPI+8xQYK0nUEZ2wn+yYcIwTCHUiwqJpOT
fvFL3N2e4FMdn4oPWqqPI+9HfI0zLiD1YReDajMYmGZtb9pgRhyZhQGk8hJjXr8M
25wp+k8I4G+V0NtNro7mU+fGzu1aCRP6yytOXe6UxEdiNulJ7FmM4oItFNWqVRzK
itsacqjyBDuwJakLTe5YQA9jz1GJFdUiJjHnCuh3G4/Z1m6cyN/ln32psc+bAoOm
/ayjrj+6pYSE42WMyW8algqFlCrQGB51mVqi+1Xv2DDYAeFY52HvnfzMkHQab+/s
F7QCCU7iAePSeoBxBIlgdmmhsaykUmDTV37az20tcstWxAm1a0guCcITwQKtEeot
rqlvBwQMf782s+96j/zpG6zg+WQ/k9OzNrMx2ThV+DaVwHTWpV2xN6B2p0QDr+Zm
jygIIutn3JTYCoM5UqRvQFsO1wUYNQ2CLiuUssyjsZT6JqYkFjWlJENzIXcYNDGl
XF4l+TYAhOYPsUSUALWLDNT8P7IwzF2XNlnCckgthUVoTt79i7Qv4rQE3DHvVcK2
9gP7QQrHuekcA+f3s2BUTHjFZ+0zsAg/OpP6StTtP8L448r9EBGrJNmYkjl+JTHI
AUVR+V4AXwB2nhJ63lLphgWPlpFyeLIth0mahsP49s7oN8pVv7wBhlrhFi40osU7
obNGKillFqiXYENAtLFH/+30aJM+/X1GNwHPTDclRG1+9FO8fucB9y5Vqo26Day/
TU9gug9D/jYmFXdaKwbK6uT8x3QZZyifAmwx2uwctsCGDmOHyYxCMGlhjMSrOzBy
9Gb4zsieDnpCBJjvh3DllFKnmSmw0JGu0mWldhK6fx6zrz6G4M7lRJPo5USlXCND
1IM6I95Wc7JUEb0uDfUPCTRKbiZDUY+bCLjxHzrJQPJSFTbyKOC4gfRKG6ML3YXc
8gaNcBeT2HGdQci2L4FjPqnCFSfRbkDDZtD8X/ZUH/kwU6yLpSsfzAMcTxt0HprP
HJXdfLxTq+x5C5HVcJ8k7vblKK8sVs42e7wK29n7BhNu7vdTQij1akAXEt48PftT
dPVj1GSBSCpErcxtNtj9ZqvpMpbJQ55Fhe4IQ+6zPLtHYcEyQnhmNAys4wcu+rEd
sQUgZa1+FnfiTizw7DGxpdM2EbW/20yjugp3sjBc33XBBs5LM+fZ0JApf6fwbShJ
JNMe35Moz5qylmy3i9cxRDX7TiQzaGpcz1PkLMZsnLvC1iXo+pNq0zDxTdWFjB7U
UE42j/w6HMitxiJA2HoFRyZbXQqysHOQuqF11E8VXa8js0S2vWxSKicDwtO7WPn4
rlMMiVLqr2V3GStJxQQKw3rYTJXJeZ/+03YK18Iqs9s8VSdeG+7iOjnBYXr/Fs6c
t/Xlty2DhHyi1uvw6pZw5cclQXa0UXN+Q09Ce05FJTT7XxlAHAAw2X//Dg/t8SvM
BMVf4uWkD61Q17C7lzV5X3cpwKaieE4S8YkA6s9RD1fZAkljvJrYu/hbuanvWF21
wlSGYjhJhVClJTEE6B5xmmMmFMPgAhCsKK6VYc1GDYzo2dAHDf2KQdA+7Q7yb0vx
PAXw/y6UzmBdOCdnv0r1fOhmZYqIUY/MbBBXWu7xM6D0sS2pTN5d0ARjzEq1LMkI
vPQu8KMtKyqa5AC7hg77bTIhzgD/zYMeTTjJ36rs8NO7o4V2mLXckt+5GuS86Bpj
4P7ulsO5pGb9IcUkG471helQWTHZsmlK5otQFs5iDdmo5M44OdRWFEayi4u0/cff
Y4vQSWLMdCweNrXFLLsE+ET/KLQ93af+emN7ov1qLkwosomDZOjK9MbRk/+aLE76
DJpym2vSk7FMPAAzgqxKErJpmbzZD1JFwiJsZJM/1KGa2rYmd0XusQMabiI6ZH9y
gbOCshwkv4o0Z64bLBIm+eurdFtgxxN5pPUVdGH/J8zPUGx4XJxAsTV6ef0VAtqw
u81p6GIeLStZh5SJzQ1nKcQHmGh+36znm3aYfYGR5nDteGClxLricLn42Bvs+mnq
mQhsmvTqzyrKnttLPYC0d9mbvNuZl9MdOYYR1/rteA8mrGyhJ0osPCK8wNygqdCz
vaIKI3+/vrcCjOOF9UE7K3960eK3Cib+lskk545XpbPf4x+3wHUKry/MABZuceu2
UjtzcgC9fXaDEQqDUzg/fbOfcqV4l4gZNrXtrpujAE6goeo5aajB8XIUNqWenJge
/on4sJjtUyUM2cSrJqZd99Rz30MxhcWbf9rrOTzB2SE16YlMTur9DGcOZ+0rYirW
kvdxVJSrWukOqvPwNGAv5hXOi7SWpi0ykh7FLnNbDvob/IvU3gTEZ8JNYZ9xcW2H
+KFU7et5Ps3pykAGVBVT+csNzrwKfXWMMUqNqqFZfxWevKqyJoALBO2PaK8Zz+u7
ISWf/w830Ex+BE3RouVpXVxfIrjx8mG9nSv4zKBaD/AjUYlMb9ZJ8Mc2pqh6Biut
8+UHRQKFJDdyeJOz9D+gJ97KXb+5IIGuNKpIPqvlQbzDIrrW2eH7Q//CX4YCa1Xx
BiXxkt9QryFz33cwh8j9GxXjM1kPNgyEM0RN1tJxBQXB3pt84JyamUkD0M1ZCFvi
Q+YxIsTKC3345T6I0nAf6SXwCrP3TR3dHA9hr7tuaoRoqksJZY7T198XYc6KAvwQ
+hME4IWojuSrBSGORkTbtq00D0/rann24z4gu0DJFxRSxwRnwgvPoo/oz7oGKbvY
Qe5GJYHyaqPcKmNpyFSPMKWfrSl3pZ+XsyvluLDlBPauR0NngwrmQ2kamMBG9raa
xswN8v9mM6sJF6LsftUGVX7ajdVL81nljoGN019OW/1iASZbIiSZeUDA3rvIEM1l
p+TE7MX9popVD2oH8Pnsqe7oJ/3VH9GJ+7zmm5Fz894CCpUAx4LjdXBf01/Ju34g
vr0VjfvhekVxAbA0evEknye3EVw5EiyetfwBslcCQnPO8sjmskD5g4GQkHbq3Tg1
Lc23JGaqh5YKTsV7qEjBOhrO2JY/gAQVxsef+h9xvFx3gSHD/vLUGGaD+tlZ0UH7
a5V2YhfvLI8nACfDFTf5+W78GE8vjlXNmydzYvN+Ac8QvdNAUE5F5qfn9BTVbQVX
PMOKKJQMVY/xaU2j8X3Us3FbGulyb0n0yUP78NF+HobCy9v8XnkcqjhxlTlgptrj
h6dI6ySct7fDTZm5va2d4t9KaySbInxCKRAckS5yyiLrUc1JSMlbo8sCRx7Z58kY
wMuLB7J63W9G4YzdvZ0hOx8TfqpCmrPZQrmCJ/Q7kWZ4Ttf13ErtzdufPxZG4Ygt
XBcfEtXaKNohn0bHb+ODCkj2z/GrCmFFitQ6FWqIOzmvK8QWRpZjsXj/TDfUpci3
bU4Bb7eE1bn2+A4dtdegfiEyv29Vu5ty5RUf6eLLPC6SVpENvLZ+/BUtE//AdmMZ
Yi67tTBgtf/uQ6Te2lXnZ+k/VXXfoQlsVJYN0mfO97KGE7TULwFQZDpp9j8wkien
S7kJeKeXPS3cjoL5Qnv6jqxCA33W9oM/v/01J/VKN97GufJXZwwtygeLbz+gaGmT
J6TlvR2zqWGidApgPIlw9EX9mGsYDnDoRsD9I+5p8szJ0uIo+Nl0NPJnzzHs2kTv
A5bZiDm/fDUzVOgWnF6Z3OxJ/04ns1MFbV79h1y/vK1jX1eV4LxHiQ92NqF95tqg
xKpdmaDMUlYmjU35cL2MQ9/fPahEMCAeqevpSnt0DkY8QLCkhaldUuAe23REktMw
Njej+GCnuo1p+UFVuGQLgtkpqLIJQVL8UFjm44b027uEI5N8Hu5H7GIDS4TsmCb9
gnhES+iFiAg48dwu2+8TDf1bXWUE9I46J4JAa/kZbhz2Z5RJFjap7PwUhwdUBOEB
XRWlMqNJueO3lZoWrV98W6e2WlmnPXmg1m9exzGPm9uoEr+5CxPLFDlEDmOKESOq
OTPpCkted6Tp/o5pDmoR+0d/mIPZIFbwh7S6U6ffp1VUFShqOIgKlXPc6cvS3ijs
Oo9ziBX0Gmp7oZy86nHpUUrFbcFUE5GCwZwQc+uiImesKTAfFRy6c2bIrCrwpSnU
CvtTYpVAl/rzvWVgsv2JVsYFlsmhAj96+jr4c5ZQ9r0oTlKwF/Zz3JEDyQvHYMgk
ic5hkTmxKgNpqDG4WbVCdBE+OG06dA0qT+jorIaGGYLz0cEijXPQ1D8gklBlId6u
T9wGD+YP44m87XA5QZMFsqKc4+gKHrvQyoZCsX/aEeSmlb50Fp6ialfP4hrBJ9Jk
fiWlE1gXdFuobBTbkzQ3ZzDz/LEKUKCkqSidtTp7+MwM3G4whN9Wm/uzoQgo6mCw
7C5NkD/wHJBmMCUufy5BjTfaH/M1qvBa5o158/B0Z8f2NB1/0cse3TySuxV18z5w
YgSFvPlmEj1RgnsOfeJtR/4bbLfPsr4k/nFdcMvscmzEUl+KT3ve61Rmn5zD3iiE
TjmIgFn7v1pVF+Aapl50xZ8gIopMXhwVBM0wE2E3MPMw/tfEQgJ0b/4dEgL1BtaO
cKkAubuQv5YLCL/9Ke25VTNnFGA6C7J0mEzaeLbn/24Pve6bwtAvNSjZOCLWTzlP
Y4WxemLWF6c9YkCcQm+gd0R4vI9PvXXENG9TjaRzd7F1q8LnqxGB72+aJd1ScdkH
VrM5hNIvMH/0WSZCmspoh3+/BntvAHnGgCOUebpfPp8bfOctNgcYsFs1XZXwTo+/
jFh60h7/b/cZQylPZGb3OprVbb4fvNzwK1i6IzJk8FuQvLGAoYbJxuQC63uoe+h0
tSWA6ds7GkAo5wYuC9dbUNvLgJJE/JzZtZlq13lMVgCSkY+q3uvFNrgs6sR20UXg
Yiq86tQmh6lybByrkV/Ecy4b7icrxOatmKucUood4UuwwdxHfgeUk8Pd1K85TW37
PZgxZWlhTsEGWvJO2giYlmAAmnwvUgo6Ppech/9c7rUYwbLIJOyP5j5W7u1qeDra
XgLW5oC7FSlWJS3KTvkhE28iUYm+WDmRsRVsDldbZgcBQUjuURV5epN8LiYVlhDA
wja6yl4MBH52NBWdERNg6d80z6pCzREy1NVxK7Na9918rW0/5xkSUeeHYBBg31n5
lwtWljW36PQUCUYxftciYcLdhjHKGJLUNbI5unS65+g3hh/gTHX7NENaUhgxxYQh
07i8McUW9H8DRh/4Fd1WyHlzW+G3x39/18yW962ABfR51mkZNeyGxy/ay4/C6Bx/
CO5uswrmT4DuQEApBaIsLsUJ5gRHoGHfMPCu2UoLrunyXq3omfy3mLHnzkPs0Diq
YSaHHFW8tCEKkKr6mqkg3lMAircQcSfrV/spKf9RDSTvQkdz/unErEoiIDrtaL2d
8Kcp+8xiXU37+y8lTSbqSRcCCh7YbgPvfswfsbeeyxQZPpfxs3tPXrp2oiQZMeqj
lbS3jIUUuEzQQskRaiowiQ4C30lC6obpZzYqp6QZZa9qYqezVNQ8F3Ep3rtSAyeE
HCPy4oKAhCZb895eyn+YdlYh7L8gqnwWXB3vyZ384DxM3wYonGQqzxWuLnQ6YIjx
ydW8OYNHVc/dwZbbqE+hFqR6JrSBBC5bXAoerbKta4pctQz4k4hdCC/1KG4vf6Ny
pakolwgngACg3CrQgnt3qfqmmSPHb6oXfrhXRL8nAragFHYoUW/J2nLMxrs7UouO
b3aVPu4Wn/9RS4Ca+SO2ZLkSYIMVr2uzZWC56GH2OwheDgWEdAUpCGTlRUAIDlCG
Z2GpQwutSGl0tyEBe9wqnghFI2RibU1I2JO45coxWxblqMQhMg0B3QKBVRUO6wAM
4vjImGqCHzXi6rfJQuKvpcH8xNwIjje7xELtZTC3lcdSollxohHWFjq7lWXpVERX
zu76eil0Sg/TZy5P/vmdZmvo+RXfR5BSq7MY2YGmLT7WFZgeioGPiSI10O9/Z7GX
XJhxlXg0Hsd3uBk4jtFR2R4kx+JzLVJrHsW5+btGfdftIFzmk9/txiE/V8N23TM5
/uV5YsSRKtCPHHd26shTaQvEH88B4ZHG86bYFXJwg0cNps+3otjnzrGS01+SYUkC
Bd9/imDdgjj8W9FM7hMLNwaCZ/GXbdQUCiMpEw6SejsrzlUrqpKUYAP+IoFyQLO5
BRUBtK94NVitQzuqsZwLubCYk/PnIVPkJ1S92IBi5jkEXSoxz9f2aJJNnet8e7ot
K+4WnCLTGAp07czczURtb09vHrFUIqDpAqnTpc2dO4b05D+sJ0PMwMPjFhcdkWcI
Zy4OqOG8QPxu1Gyy85py4fcsZ3rUkNql3ePukU4T6XRctUS9/3cxdembSE6N++E5
IZBnVIgAomXMQJF5q67k5TtkDBfzYh1WrKk8dmXq4rtHmrtAObnChbLLv8RzHbp/
ngsnI7n8kfedhQmu7jtxvaM1MI89y2ZQfAhZDjGcgHpIjkPMK+E9V7dLrQnuFnZv
oDf8ppZtmDZpwv5ldrh5NywlPczMevxoJs4bdQXW3n09xfZUX1aQa4SiximXaWI8
fAn3mF7N4nZz5yOv67jx0YedJ7eJm1/cC6viyH12DqCwHALm7fd718QYNfvCiJZD
GmFYGj4p+GvAL6KfTvPhyQX/lkBddXTa35/gG7Ync93R2lfs104RdZKoF9bHwxn6
C5dxyvSROWkybVjgfvJyGDD8ZoLdtWoIJbOr054YM4Y7Avc1hFe25mIUcAripX+c
YEyaLS2nhZ1fMgiBUCa0D9JkZEG9V1CEnx/MwAHpchpyWAfCrDIx0bvZG8P0mhnD
yIoNx5NVXD0tDs0O1MtGVxzZc/TkBAY9g+lK5GkT2hBT2YO3emZBOmUSCDI83r6L
yZo2KAt2HWA/flhqvf5rYRjTuQyzU/QYVVgeWnvmmOt0BG/1meMT5PQAfyO1yEkM
b3ZbP26XAICFuowhU6XV3iU1mgdjyOchRXmNjsoATFIOPRN9mkQvG5lS7Cb20CHY
vtSJ3xWkRCYsRtzoRy7yWrdVHPdrDHAExK25rJsVF2f0MXnnpGs04SDmU7J9mbLt
tRvlffLEA/6+fQXh81keZHjHDHJEFmTJrm8QgzoFolWxPSTMeJS/Xqa5QdecI7VZ
xJaHoY9mwSnkE8I5q0V35zaAuxq9lm51/r4EBRNLiKiX3G5N0E1Zi5oH89UMkMEm
ToscxnAjM/XOuqNi4NP9gfGrVufnVFYuapCRlOUxWbaZaPZijoQ/gzW0AdFHJRS4
9Ea8l/MoBbDS1cEjvafPBdf3R4PCkEHkXNqCUypRsts0s3NC2Cm/UGGM4psTXx26
7kAxmZjenTR79SjJ8cnQHBgDzLc/vXRj/iio6u6e5L1gDIY23LuvTcmbjpVZBM6q
+cC7W7BSU+gumMS7gaj6hifV6B4aUNdTwDvO0P3CgkcrGXe3UjoymCb/Wdw8qoD6
ilLo4atpcO/sEMfCKkGswhLjHWzLYzOBhlb+/So+qbueRHSnVUYnO9feqULp2UdE
RY73pPTtmc4Yyn0Ry7lWOJT5aCYDPtHTNQmpopMuyWmavfbfuERPIEp8NHhaF1II
oIS0JUOyDUktBF6LHOtAWlZG/ZD1IURksXpEyb2LUXG7pSEr3KfOVOXbtiLd6A+t
oXeWECukTy4rNYVyQeaMv9UQNkLwPN7jSEXfFAw+YBZn24NDGWwKicbK+t4SFupp
EeQXyNOeueEL13M2PG/PQErqY/vkND6zd9ohSvlIUc7j5kac5jStqx4jAfgyuTUU
3eWnHwJRsMfwrAy9J2wL6P0bf68u54P+NYiE+IA2HYW6YTqtY9n9cmV3AQYUkNtC
pQv+De2F3P4f9uJaPj0h39E02zNSxjftCafQEwR18cx7/CQlpJpE4kSKbAb78mfU
lqqpPgB9AmyE6YVl1MZXMzK2cpXrHehH9pehyVHCrZpFTrjZGEQgf0RSzZr9FWeO
K/jC+TaBSDB90LkmUVwvDWCMO7TqWUDNRbyEdp0KQ92mhByD+tAvBs97pOpAVci8
DJ/h0AdlpQfEsQTVAOob3UlTKrNH7CxwG/WsiyvRQQ9ONk3NULddiS3p60crIEeE
wckUeU9KgCZeRKVPXEy0iMBO/370RWDDMwcxKBYwqZUWpWE9vWcfr33HMMpZOF61
G1qRjqitwurswt6NS2hcJYGqJI8V6X4lrhuwZYkdUy+rV57RXzaFeuM6naLlfwaX
uqJhDGEfGGh4NRBuNIYs0GQwgWHWIl/jZEqmWLzU0hQ0jW5E+H9ntov+QC8f886G
1FM9k6AnpvzH+bfgfXO+Ee9+udezHI1h6XpAKTOfkRQFuaz/+PjuFJwm0iwKFZYp
1q/YnsTmWwIOFgphrTnNG/JLgsVnQDBcLqDQW6bLWM6ufiD5IhVjh/SP+Z9WxcGa
MxzAmGr9PnLFLfwtBB93zo++xqsXyhySApnmD1bVahKsSG3FTbX7R5cfMJ7Gxujf
r2YlbMgfr32EfyiT3Put6wvz/o8dVXNVxxDcqT6CzLVCYmP+SDAp25kwMkegMTLO
jTSyAWbEWqlpf1tWnw3I8xSPJJ2/URMFAtJdNSTMDgwBb9TVYrCUKx0WcMVD8D2k
QQl+SL5NLKv7EfUD+3j/X0amctR3oFGfoGBq65NwaKjMLJzIlRHXzaeyXz86d/+6
KE/qiwAPX03/zwIv3YDQnz7PAYnTFjwwxxJa2lOl2mFjGRXEd7VHkT+YL2BXbN35
H9rvQO08W2nRyW69qt+HFB4RFA0H89CNUQeovwPEfutZMPmYmu0eTLV2eiLtn9UT
zlnTmUoEX937nYSiFqAmBjlJCb90a5J4sLkJe880DdHlkczBZZMqWZQZmvuwsgXK
6R5DkaCsVaWYursaFsFHe5TqnAiGFxEsqFp6X5gWgYmGsBaVPGb71rGq+wVwyswn
ucsBuMy7TKPhPEG01hTVF4RF0TZGMm03g7er1Ew9n5ohfeET2cizlbve/VkBWbO8
yRgfLpzg+UvEE9kEIfHXw+7gLzJX1JgXbpNrDVp65qrbMfB1WZiHyw5tKZy4ynUt
ybltdZNKbbzaCwHgI7IIZ9+U38UUaCDaVEQnqPmgCAN714Qn+XuNQEZllzzUYg/f
zITgV9iZB/K65HH/7+tAeZly3KDJz2AIhZlVUhv89SRAp9ZcT3fznE3L1o3KCMoQ
PFyDxaCP57ePoh8apq//TRrOlxPX/B/JcDCfyVE4MrDsbqjEWlARSgAW90wahE42
8ZbYgLE5+MJi40S0UtwBW1Ra4QNn5WTyhMkmULaL3ouPqvHZxBWM6cimRED9DfVi
uDUe4btIbMqcwj0VnazA3TJYsgENNYKv/zclvtHjfTq2o3VOeJ5E5e2vVj5crS27
9QoGNKhvDHXVInyz+4zcUW+iezAEJV0CRV7IJElHnuCNDFzTx4LtB6D29xV1mou1
0QnSw1tw6Q+zcbjH9Sr16IO1lcEiYw5mJseoZ1irvYN0lj+mqGQ3TNZluml9hxjw
cX8NJK7J4ESDmLaDqO4M/j131DnaxH1pFdnvi8AJicSxBTAXKhU+8ZqgFXwUb+m0
2dUHI0FtZ23mTvYb3vQzbgubhLTkMy6zlW3EadqgdCtc1rWMGNqMwz2U9JaOo3cS
yf0tsqw+1e53XR12M/gnI5CvWuHYxhIPaWsn+tZBPhZSxThbHu2LtiP8svdDmCi9
XvQZtO/odllUabC67jJpsV3aeRKrM6WLkDTZG9jKofDw0ggNPWPynBADWK39lEcx
COOUfujwslYIf8HJpSmkvwmECvjTY9/mfAyoVZPhv9zir4kOKThBH852ODhdBWeR
8lbI8v6Cqcl32+Iw/37sfNnVpzKwmYLJQ8abXg2PPcKhtf7ZU2JrJemPKxRZptCX
1mSGGEmp3apx/su+h0v/BZS2eRb24cH5NzD7Q4fVCVIWsaORmyjPbDhwyVGG16Na
jUZPCa2FWYKS5PO9NeWTL6qHz62gOXjLLog57VhpgSz9jlfMMC8MsbSKPvLlJBa6
IEy8RUcLsi3fl5WUalu4yLp/NQipTgIpNp7+oFU2W7jOf8hYE2I3sJhlgJW60Hta
ypDnfIpFzOBSZYpFs4EMlOpX/lZEq2pRtLNG75rMI/iswI/y5NsFlS1f45AtnqjC
ekKTIUUNU3nG+4O/tYXDT9y9KtpfR+eWbzxmNmpZHr+Id/cOtXVEhee4vo2tyR9N
vXpnnqVf1+uLrjQ1OANqLh6PNTnd4ur71zipnGWPTD5Q9yPm3YN4YJz3e6OUp9qM
EPNllqr5oaBHAttL8v6QIETetVstYTq+dUH2Eb0oubv2LmIiXuc6piB2uwfOxEKH
AG5+VpgzUndamCGsUjyHIak+Opc1xfvhDDTaVgTo1A1BTM1sB1FcgxkOOrVPsQgx
XTB5AiK0FyTruAFQNgmRJI+QYjqeqT6YebMKrrDekbty0HMRWOWD2ys3vQ9EKnVo
9rYD9qyWf9bwSQf/jCBYRi1kr2XxL85s8s1kS84xTIwRFlNoT2U+wX0qum/ww770
ev3CRWd3a1S0ivNgNIrIXVdYolZP9SqCMjoo7nVufr/iPFDGBum+fURW7CkpE/3r
RBdKLbyzCQoPX3Ac4neZFwROc8ZM0t/e+lisxcV5bg8Y0PtU0AI76AN8nr1bIxyz
mvzT3bq5OzuISVDugDPjURsi7xFTVcLNMYJVmfeUvC6EO5f5B73ws44uG3ml1JXL
skj3V/o/IM1PGLYOw7Aet8BYQMPhdhhMZfMqXBw6ePK25+4pMkrGe4RHLtc9AOhC
VjEynPsie77lBwB4DxbSEk8E0kjn4yeM1+PCzhtBRwDmxmsTYARqjTy0pGX8ZvpM
QHvRu0IqbTcGrBZB8WTw+mujz2TPRtY2lVOoUgMmht6WkuwjKmFzHPjvTWZ8kMhj
yiVE4EqWL1oFSJ4kALW83686aeUcgRR5gS+ZLT6rw//YaqAWcEnrzoL9NZUnJm0p
+CY4L0T21ywxPKL6GvrpLM/B8yM9nWPfxigGguFxSUc/BQpFmHpLxFMRzv7jFbCp
w91mbqmCL6cFXnC+iewH2tmW7WCiCFJG2oHMInG5vOGS9Nj9Xy+2oS+pSn3wfBu3
STTtZQKWDPxRPSaIAtcxgf7Vp7ivAZxdifbZB2pZus2dq/70seAhdj9JuKM7u2gO
ReRSxlN0r+H+kg/rd47+X3Hv2f3wYO7bjMVt8Z5zwdWwCh3L8Aap9TB0eVX7oABy
9DzEaqIm9G2SaK/PBj5cl/qumoySpZ2WDqmxL7JBPiF0B1MdBW2KuCHkiA9wKxda
mx5ODtbujx0KtxhZeJaUWfvh9YYzx+II4ZccECQHuGFhgKBGdy+jqZWzYe20x8pi
1wC0k6fe+ZfCUuBPbsP2EuTwcD94DRtKOSXbjcu9ysOxVEoqbX64uC+BWD+oIhH7
ZzQ4guWE92BhKCGWbEpwg0+8bQ0Gc3obFQFMdsl0xfkTiYkfDZpxBS5Fw9H/JKSJ
RdO0nZtgCEE0Ue1VTXZ7RdRuYqExhVAvyvTHZhUhkdE0H45sAUqwkUIg7tWrdvRY
DZoq//ioqnnKLmCeK8tqMfQwXGgIBPVJCB/SAFMFRPZ287cAZ5N3MQI9u8jVNrKB
6wVR6yZp/bZ0ir/H5W9Y0XP1FEbbBR+wVCW9ybd92hARTl1D0en9UkywZha+iLU0
JhXK/tlgbXwT/dGVeo5EfyT4Btw5IKQ9lT2w3XYD7UVp2YQN25MZd3aMgJGNzi8b
2ov1JzjUruJ5QQSqo5HUjJZWC+uTdvl+lWwwwVAbom/Av2Fm6hMCRV+n426KWuLq
kryliOnmLGLcf/Fdv6iQB54rdSxeS3KeNCnsh0l/iHV74VZcZDYYrP6pGt6sE0WW
7ObhVuiMX/t12dbiSSVn9ratJnCGzOpE7UOuTdyBNT7ytigUIvLSrx0oXyIfvaEH
ai32frtXX/yoRRftL0qHLJYVJwV097U16ljNtCvULX8+jh/4mT3YOXJZO0MO+Woi
Gl0BfTB0Z5lMuBh4Cx+SxWkCLKmEB1gKIvCL+5USKSOzJL9sBusjSky36BZhA6NV
+uCCWqYOrCrnTWaAb0l75GjisXl6SwQEmKATcRTNZ28N6sHkyz/uAnccXEW2sLTn
5sTv46B5h0IlepxxP/W+/pkgQmPj90FUA4sstsSdOHVf08j7wPHSdutZh0MkhtnB
j/3mKAcuPXDiykgBGCVjqk7HAGAMSw651sY91WNLJs/YeWLpIfdHMZabpAgzW4TW
BTWAAzieQvsn/2tG0z823STV4MNK0wPsS2O1tduNRnFEucVqdO8QKcrz8hycmMyr
ISOmPdrhnryOcvaCERratFBxTxuEfKCd8O+jgBRH58xCYr4HRZ/GrDxoBAtJ4X1m
F/X6y4slmtazJsjGdlY0N9KPGQQaH+Jngk0XTQuN6BPfCHEfExgxhllblPTiLnVu
c2xT2xzcVWt0VKnsIVuOOOy2j1YqwP1Qdpy/83VPxfS/uThnuzfHw+EpTsZ2uZ2l
ws6XwLiURt6RRq/FVYl8RpJhf3tLbvnHVr0pfmQuD5KwIAnrsa3ZqazZlbqeYzB3
DTrKV1gYeFZiZn0SXorRy6a5omrn5LcWVzY0dcZoNe4qJI4JLAx0Kx+g4Qo+I95N
ugu7IVcdJ4mZOZ5QBsaXLipPExlzLthebrNXcrIxLBlJ7wFQfrIdNxGYpxVv2acE
ea53FFxLHPgHo/A61UT3REfFvx4AAKnt7MlcEUgNzbM63DvfnciaRedE3s+dmJ5l
Ecqr9RXSwnvlYJOxhBu+QgOubYw72kQTTiaTvBn04Ohaouzi63MYynlBnQTtfC0d
H7rwS+EN9lY5rqst8y787zGa5MC92sAao/pB10dBcTzQNaMDN49UYmjFNPotXlhv
l990Tu/eF+7c0wNJqjCjsW3hmtE4pO4BZLH1Yb+IK8d3Ns6t3GlBly64Ynavvlt3
Y0IXqMSKXpE2Q8XyRuXKgtu04eE/ogKKIs2xyNcF3CCVsPzaZjPR4vqBDBvunpBS
ecoxHapuZYj4WEktwA7FNfbwplw8qtz+YIysjpZ4Q1yanOzlEyqBPxq7MXkUQZYP
5ydFzQVJZ9jED1hKKh8OF7Mk0zkjC7KagiYn3+jcLkHkgE2E5HkJH2xHCZ00W4hb
jB7uiZmZ6D6a6stqzg4+Av/mH3hg9bexeH01vbA+e1LCYK2VqxVu7eWyI+wHANn7
FXg1H1nCstWXg63v5BujBk7UGizhk1ErKwoyfUS+T/SyTDA343ddnBWwsyyPti/D
JsoFyLTh8L8zkNThlfRRx/VhrFAzqFF2eZl0AbIMhIedMSaeH70vCQt6W2iCrc+C
rOVXtrgsM93OdC2PVC6P3voKPSMq8aSx0lliM1GDptiuMB2p/b8PKe53OhpDB/oO
rkgPypuPyP+qyh+FE2PgP6PXj9OFc5EhVZxXPdLAcaBP6cKcRHbT9KKUl8TiiUFe
EuzQrYs8bkGhm+qtsp9K7yZDs7HDSK+0KR4IGtSvc3rWqLvQ9SiPn+f38Sv5silB
SWvLjTLwcIw6VeSXcfweJpTgUr3bKbCmFwaC+rgkUiwtsZUhuy6EsiOl0QqUTIwj
vlkEmAECVRYfbXD0+LYEz79rgaFLZz/CHOETQsCd75gIeKR/86VsVB2WptlavdXn
qCSwsPP65NEqJDg3UCJzpaeR8sct3tBtjhyj1m3fxAI7CoJ0wy6wggdP1PR/xgkY
OWmfK+CY+PjpICiqqkugBUC8MWPCGFrzVzmTiPO0y/+oWXvyG1dU9HHz91dI2yIW
8SGJAXy2x5j5CBxJroqwCmu9qvM6XENG7eoxnvVQ5N1mF1M1gx6orCtjk/YG6733
Fy+qt3T0CiN3D1rnFetonGsjlRLT8LpGO6ef2XRi1yS6f1YFbxtbo4y/4vuOidtH
0TwVnlNhY/nlzdagTVbUPruII45d15KjNC3VGC3yAwxABjrqF2vci/BH8/TNPA43
LNzzm5p01g0aXAujAz12PEcJ7cawHyoiJN2tpXvnhWCJ0cFGpaBhX5SaxkDboYKK
bFhx7K/7HQbY0j9qkJ/y4dHSsMKlizQhhnce77J5LD0tfwSJRt/wXj68OFP5pbX3
2z5sX5kLeLad+/VILZ4SnNsHO8Peg7HXUDEaDdH5tNV3Sd71oI24ij43TjdXpZv+
GgdWP1p56DAMINmHACuDnf2IMvFaFxPsp8ndtRLC2EO1hE/DioUMgc9eyKGaTkIu
OgjI39GHIQtMpAmgKqOMxpPoNTcIMxpg+8HhdWYGfGb+Hid83fwOYl0Tf2NbvmBF
v7qm+62NoOM5KRNO8N4rQNTzfUH4LrsdK/Ijnc/mKzKzuT+5XfgTla9iNAvsVopR
A9qtpng8gPBKKjFCKV67lpIOtURcRADyXpd02FwKemJdyRK4XZoo6GSVcbpDrWFx
z15xWQ4Ao1isctdkClTAyy56F7NqGqQ3+HIrF9JW7GgKrYr6jDZqx5MPo25t+NsW
gxqPBMAiSkPfHhV4iBcDRaVjnMU1NDSS1pJ+UlrY7ZElOaC9DuqT7Br3ZsKRCBPa
YpfCvk3C71yQIYYHbuD+bkuK6Tqt1g9+kKxLFnRqxVQnjI6Xrt8th81irs/wBYfN
u1PqfJngFjtKZRXEdYIVNLWmV+8oPoOya2v4ayuWuKSxfCrywLoocbrZ9+MYOtdy
T9y4x6PiTmbAA8YTBEDTlfJCPfc/r5Ge56fIM608+jCY4uO67+YgOEhdkO9bVvHH
ygqDSP2xXkozRKShWLx4fMho/kKPfRWGmVRuejoyqz1sDHjvuvBYpQwOdWiYNVNT
F/cDJ73BiHWtYzsYFRsu8+9zKcq8/p5n+kouoFmzzs5lf0+QlLgSTl8RJ4tfHU4R
Lg6P8hMBKTvNVaSxkA9egIhDAdaMbElVY8rt6j6+VkZSobpYM+1NXPTu34awCCUw
DZRSwesipkkpGTfUW9c0YrfVh+7KGz2v7RnDT2iLTHRLmEABJWON3Sz7aPPZvF6r
bXcYFe6LtpzTlwqy0UqLlkBLUBWL6rs7/P1IN0OBZLq/1x30OvwhAn7mS/r0qFNT
V70E7fdJvRdxxhK2PYQDb7459ldPGa5I8d8eqWsC7UfRr62aC14veGpu2LDpRnEw
EfeX9ck5XZOKcfA9p+EjN2t/qc19Tz7+gYZ1uI56aZH0gneQUpNEXnfKZ8Xp8sFE
HcF/SS0dI0930FbQVj5doRfIUmr18qD0emVi+E4pnSpUDmNSJ9eT7mmYD1aB508+
ggosUqIqMWlRYeGhcMKrBpLwNv+2SG5DivZ3D1cZ2lK6BQihi6WhMfMbRQGzOGNL
krORf2v7MkcCvkhpmuk1k1qPKX3BvqwGDu07e+O8IasYpVp+Oh/1R+1p6asXjMPu
1cJACMJyPxYjKMMGHzWSS5dg8LRGIrtMcQUguIA9BoOzk3z3sfudgtbNFplRdxCz
vKf5CZ+ir9NGTzhPJ04tIQ0ev1I9dQEEULf1EIu3g1VzpnHhLG2BkOaaZlhe6128
BtX6C33HcV4BBbcCAlwfcPUTiL/RFxKio+Xz53/rRt+55FfuI/qkyM2ZXfp38QMb
Ku1Qyk9Q8pAzayCWNLONJWyK+rp6bf7Q7t7L0rdoRGHLx5nGQRwsnPnKWEvXTDAa
OGum8jiJeS1SxN9go007ob2zCjl8vY146+9+SAQd9DexQSml20b6bj3D3hY8qSrg
rkE5013w7NwY4OBQAWLYi+vKy4I0IeeuL8o2rV+jdiIOYGHFCIld1vsezW44jYwb
p/MDaM5KG+vM9vaI28JYdhVFL+rfJoSyyystiQAFik1bi8+MYIX1BRz25TzQBv2/
MDjotLhLRfPg4dYqDVHUVGtjq8w6Imgi1+ZHTKV1Dg0KfCOkc7kiJSymlrD4ZcWf
V1Lf4AzVfn1NJa5hOujQ0p2OiyJNB4dnO1WXUnnTC6ItWS6Oh58JOtHlR+nRmDpx
b92zC3axSNyuQ1v7kfgOHrhHFBXARKPy4bk+VDTnawm0zSzoJp12uhkOVyIRPiWb
kH+uPvH4XnkPNnc6CeY+q2fB7/TutfjqAHDSf9pCdjEXpDutHdn74r6gFKJAPmcN
PaGrxk0PsMGz8ociySULkMvm+jlZH8IhPiks5+hKihQ9H5na9ETOkDZKi/0JTMxX
m5EUTl0LYBhZRGpKe4kPONoSlwuLt0ZIi2E8KcRK4oj6S4oIiYW4AQ2hmcwmhpAW
lHhQuBqHg6VNDRPYq5wXOYazdP7Jh+8QuS1Cxnj6e+ttANGKVSimEZFDKDuna6pG
b6Pw+L6VkT4myaRjzWOoktuJAqWKg4OJ921QyP56fB+GMC71SHBo0iLpyBWvrgcR
RbSZB8SEiAKrwQuDAJHq6zBC5KhgYbx/XnntDTjAVROheI08rIkfuoy0LYJ97U8W
P7C+3zIgXz/ltFWQdqFY5Ca0Y3sWZecY2GMuz/O77WPZ1Ggmi88HJUXu0nEVPKWV
YpX8IGkL2ZBZS4yoEQHfBnJQ8KIPbpPTuhYrWX15ts7GxaQMqp48Xibesto+X9ZP
QMUF+dBUtfuMl1mTQe34G6KaO5cxPg/4IM55HZd4g1Ivd1UurlKXGhiHd0C/S++P
JGNXVE1BajFKCAgIXKHNWziLTOVtjK7MiP1lO+YcAPIGuwiPzPDWcUcoA0kQc5ri
qqkj6rnbdMnIu4Y5juBFuX73by0RxI23fvlwsc1ll6nuaNnlWHKNk8OTXrRPUFLY
q5DKbQQCHfy6Dwy8rCAeU8pvkrxsXKpGIMoZtxw+D7fr2SK0g1Yh3edHaFoPkyiA
jLayHSkWL52peloW7PcQstiPzaFKu7ZQiIGibgTArYZo/4SBcRm3sYwz2V3InGKy
VFm4YPbNc9w9fgGv+EHbmUByCUcIDuI5+b+arbF6c0mxG7yra6bUKJHQB1hibXp5
qtk0g2ldj68PwhFY3EoLiKwb65DdIXYMt6oCa4JzcprHyIsmv0p7j2jjdp2uVC1D
89HhuC1QZolv+ce2vkocfFRtvIYSZpFzdFpugR0QU5HAfl/uSO4kcP5Ty/J9PY6W
EU1Z+QkJcXtHkvRuKj/7OWsJlHkAtg3skFeMjHwgv9Qwfuu3CtSZR8DEMBsCXreO
0EfYBGCUPeHh384IBr0gVL3X3Yyd7N4IoYELkCr/NAqJ2mUQSxSudllBlpfn5ugE
XVucHwfskL0dgOBvtHDOvOdVfq+WDOTDlX4tIEtdJJFxdqOI/E6i3G0TSbWTpNmy
jVzt0c9T0XxiVpxdIXYMPLjBr5zdlFd6VLNJfR7pu8Ymh2zbfwEJZQYWJjU3vmSm
Gt85IRqtPoEo9M8x41QsJKrhb/CoOCbvx1AAcW/MG+qSvri43fgjTCMZkBCrcrIV
D2/Ff83l7c8owUvj8X49+mo5npre0vkjKWcWfD3Gf6FEpQwE2nJPOCh/keGYwIVF
tW6oKAEW51Qvp+rbTfco4dVgVoKv7teQ4JPVe6YLmpKNVvdcQcD5DdMRihfGEUL3
F59/oZS+XO+2yOOr591FLTrXPOQ7XrRjCiCDowuS+Z45eXJOe2rffFXbf83jg4cy
3dvST9K7brGVemMZxvReI53XfA+xcs2iqJtwMJM09z+lIH698PqKqYW2rHdrdFxV
iu/RKjlhcSrAO0sI7+d67ZZUCar1gA7RqOCgO48JCDjH69Dk/2PVIbuDNm8LpUWD
26uN/qwdQ8H+5QJbNhOclSO5OwvL8NL5aINeNC/QVhqEECXa/yYTNoRN0nkEFavZ
pcYnambBmREwYvPpDc36pS8DFF5WYgX3cNbYg1QsihqyGCFA3m7XalHmc65Me7Dn
x4FuTEjMzd+MjPF8vPOV2rTkGBK282uNIBxMcrpObFlJuqmaGcDvBp20OyeZxMJj
96fljcTDqMV/fV9Q50PZAjDVZpjt16tv99gu3RNlj/ghrlW9Ie53kM/ikHkUATX2
qdfPx4GYok1dF/89IEpzKfoZtLbXmG4coX7lfJqTw7ZVor2j04rm54oaWB5lSFQR
UW0JwlwtdFwMqgVI+ZkhGfz7JW66DHHQgagzXS+0bfNzSo0yNTxBqgbeSMvteAYs
gfYUXd/BR7yEY5D/lBbGtB+lnub4gyOIU+CiTNZwap217s9tX1OFS+tCcwiH5Agk
Pdkmbpn25MXJy9kqbtTYau1FPmcRfVXAV19PE3qJPFpJ0SqKqKRRznkG/OfHh0v0
1k/rbFEzqcdkZBSqe2OEeo0G34SMAcYsu314GFMLGYa09SxvzFriCAURy8AhVBmh
9vlbH3SbTQnrU9Bz5VFMWhZhsmGOcX1BNQcP5mICWwg7Ef/8G3egx+UJgUrAKamR
jHhN5v7iz6NWQp/akDFRzN2oGVKjbSEb4+vagXQyWH+Cpadsu0CfByIpf5l59Q8d
6yNUR+re+p9cqNgXQKCh5z73X8LCnx6Nnol5SjCHN7sYsWgwNrs1mr9uZmyvebtH
vz4SfaA4qLEHMpwwAJCdElNnAQQ5C7lx8z4Uv08qq6EqPG1rUY2LRV0WPeiFumZF
5GyPh12xVSc8EVm7Z2LERkcHLpjvw2Xl3lSpdKVl2gZdPzpQOr4DdKWbHjXVVidE
JYkNdtQWj/7xwqpDvXgHpcXojtUl01jvZFIFnTwoj0DsL6G0XGEpmQvhBTv3sYh/
nGLjNfsT4d07s3VnWzBmFrE8TFRWY0oDtysJOO9gljxlRQjjDhFVrzNiUJYHiYuB
A0AIBAsUkW3uuSq7vrx2A04pSya9i8pZ+2rcz08kFWhf4lID3TgIcBY3XoAPaHMe
vXGv27ikdqhQzNphtJkjXESdSiqeMpwEmBcsdzUy7SwedQTZu8vvxvTlPCgNfUyl
fL9zftxAWKCoaZF+B3W6KwCD+TxLgemW2uslQ6EZ6seUT3dTfi6R3pY0uLX8blp+
XonpthhjQ6twmoI0X9qUdv+QUKUVFQmmfxHohXWu0WY8+39VWSDL/91yy0CmJEs1
0KHVZEITj+WlAlXCSbdDpJZSD+0s4zS468rtJ0Zz0zn+w9NeJR0rochJ/aXPQGmW
D+y9pCZWZGrvHKLm6ZF97/Mgqvw3gg+SpLbMSbd5Hxny2pP/vAm540E12BLLTKWW
Qc4XeU81W1Uc3MuSWQm1C6M7iIwITuOUZk8BVwpb9149ASvxY8r1Ecb2nDdeumxH
f4q99ccEHLszMSgGKg2pMnsMseVGD1MfP3DXKZ7Nc4jMcZseRt+2monVFfUig4iW
HphrfSIaid89PPJH8sfUFA8YqaxCB8l2asdffjePni7MlM++L3Mf8rEmW3Q7+Tv1
g6MDGVurEpZor8vujcpJZbJyFEgspKhOkUA0Z3EXPrRfUMbPvnqtJQLLwCKBH+U/
kjxDj1Kwfcv7Zzx2rkY1a47zk7/l3eiWFXpU/mtLtSjRDm7J0RKwjA1zfuVKa/ZY
WSAfUqfdU0qSEhhf8RAgCZc8X/3HyU4DB3IIVHDNUnHDhjztrqimQELnUEiJW2S8
6vZJqnuluipSMIUpcGSN+RqoHmHdGleqBUllBid7KViDHCpJ7QuINbPb37q0LYjY
QTFxmUvz9bL/9LUwiAdRxCHmA6wjHo8QnF+py9IfXanBGteZbyb9XsviudRU9/Af
tjCuZfkfrbDPFqvvmWASpM78FOI5dF0Ilodbph22qNe5z9qHl5tFwlXKz2h3pThR
bUT+bDirYL/HDf1GxcnF8a763PcJwfLGKQG8tEUyXsMsbfqI4sYd6rHrp2qYtXuk
azkcNXUYxXEoBHY+lHyY+wtypepoD1oFYKgp7OYLnd7noqao2m4q8wj06KI3cVPH
f1kOZu6yGDKiWJ4/H6I098kGMA9bSyV5o/CdaoOGI8i95GvD1HFhPPo+6tSIDOZK
O4UmnF/Sncwo8j9oQIHlBPdgB4vuM87gK9Hj/KM7D6MS/6fO4xVdkk9dwqoW4+Zd
Ige9ibFPEauupZOOx7Fsq5ACsIe2WewcgbXmwLONbonHJmQKBiQFyNFm20H73s2k
oGplWV64ngn4nG1wbZ7anT5A2gYUsaX4HteJ2uXnjjXiQbSPK0k7iyvf1CQmXuui
BDNakOfxz0k+eVRF2dY4iUD76JRIHeCID0SDXDP7y9qQ1LGZ4NVnFhaYuPoBdUM3
5NO0Jit2fOlIlxRiDQd3nhwiNJavaWK0hGPfpLITnQQDYJRD8/gRtcPjuk49rfnL
8mUNG3nN90LkkGpJ8HvSmuD2iDk8sQgrYH7z5BGGwDQA/xsHtBkpqci6IVl/fZaG
gG0VcscFeTciogGCgWM4T9gAP5ZHZkXsoyU7glO1p5exX32SptdZNGYT3zNvC4ky
9h6zlLAniqg0+5lDUpHXixF28G7GaSmVuCwF26aL4sU2HQBnAfWeLNdJrR+XOeL4
A8piVV8K1RfW8WOAIncyBVRr6lvA+Oy2aio+c5t3SeeRix1GFilv2OAkYGLqogUP
lmr1Syy2bn8zdXabncfRHbjehdSqdKV6kyJz9CqpZ+Q2f9ORTcx2RXjnQxa3Zd0m
jXUHI6IFs+aaGX4+xQ4rwBdkQNgV/+jMKvtMsWPCfF8iiAPiJpMaM5b1F9uHP9QK
DXA0pB5XOaY+J6bT6xwhdluIAHAg17SpsGVI2X/wLlUaVVKQdCBelZUVaNur7YSB
a2AS0nXHw7pCrzMqjso/+6ZpV+TjfUngz+t1wm06vtAIQXfZNVUQb4c2eDrfy8m1
orZ2wnnitvEYXl6Ai2MsfZgkxB130p2pZg2Ux1HGPGL+lLnYzD/BMknaZyUs3tv2
ElJrdHEsU3k12Wv1DWK8nMgWuHBEZvXGbtejC69+DpmIWudgTXZSxnrEqEfXnhu3
RLfCow7uO60d8AjJKhlJb7JTikue3zwMSyvbn47faTd9ybY5Xtv+NPAWTtyBVYuj
e3yS8Xphlsnc8Os6KU3X/TcOgiG8uXbrER/oQhqylR1yG3sOD53mJHY3hGSwvIOf
CXQgqOqyrsIkHBXbnUseJTsCou1IVSxxqDbMH5RoG2v7H4Hw/u8k1VOCgp0gcvsz
atrjWK/7v1T0JvFgtidLRKxWH26OuOnqiUaXh5mOzXqE9YwH9hKrtRKEC3Eus+EJ
j7M21zKPgA7U2chxVPkKTfGrG+Ahm5aN2+1kogTAzmE3aZ5oukxgy+bFDsEKJ8N1
7TW9LqrSDIm8KENtkCNNPQJe4dB+lAsjPM5pgkYBFPgmbBIomln9lu+W5mwk9Mhd
HlaAN3w9yZFpFEDLpnXe6sJVsWuZ+IYFb8AfK0+QmbJgxZAwN1qyAVwcwW0MuqZz
pxOGEc+Chm/7TStzvrs7pEyXYWlUN7b5au+GXGzBWtRVblcYpZGzCoxcYGhqoMqr
X3SRHF0gggrk3LXFKNqyGyQOVUdNRCqeHZqhbl/vC+RLCpiXeiDgjQeciMasoMd0
xhxsTGK5NE7nQjsbNvncI40DuApRE5T7JWubqzFtW3bhfcuXyCNcEJFO99z6h59y
WsOkLYx8Cs6zpUA5lWcq+4AhGZ7WnyqacLQZ6sg8h6K+ydhN4pnXM52LrAzMCQWe
gHsNOpFka8R8/pWuDUzx6vdtOZd9cGmn/m4eqzg6ElUvNbVkm/ODfGd4y/288Gwr
mGsq/VZItbDTHwdWINPnoLnQ8KEAFnLvoAd+qRr0B7aBSWyAjBNSqYEepLczd6R0
+9yq83QgIADa5U277gJRz4harjFU5EVZTZ8hgSCe0oJIl4h/rq7QDGyyyc3QH4+l
hAtrIu/PIEyJMdKrUbNcd0Bjf7SY3oKoogdfyNw+wCmqSaynexyUVvFQQ3I4Tgn0
F0gJlLqndr6RoFyKTKRsP/u/2Drf+vCYlmUBOTTMAnNGUfpfhc4rU4TMDHZux9lz
8f74uczETyh7L7Xb6dv1t+MfAp83+WzEzVNjZhfEIdjhK8gxADpufR96EcqtBKhR
XhbJsienjfj7GcrMERZvE1nJG0mf5sYhm7wxxIt8oqwjGwt21EpsqcJnbmClnsmc
wtPARp7rELW+cYqZiSs8bmmcet+DE1bCChbOBwilOVAc37tvF2uuLBlbglek7Wt6
BqrIrX7pVQMIdvjmDQiWHVE01CUgaa+FIhQ1nUn7aif+IrSP8dNEAN0gQNkbLhC6
DnGyW1jZZV1Et3Z8pO/0olv4XPa/b/jYhjS8sUchrkVjQ0AWdSeP5j8KVf9p3CQ2
Z3NGwQKlE0s0IV/79Gn/8UwdM5iqcpKaZZZt+5cryKwzRXD/wKHwYZhCA33gDvCL
aDrBb8a6OmycDBjLIjmA4zGRP5glH363Nxk2cpVmj9iqvQNFXap53+D/+jxy440f
kzsGsyfZfoagj6gbbVPevnrcmYzmBav7rwauULW8g+rCMpABhlJ+tfbJV22sIreR
ylsgKH04LDUM8Jk6+9scTkQX3Dw3F8eM5T8FEBcQxJPIgcyq9bPTmRxyxmXV9hOM
zPU8xFZFNgZ5c5uGi5xJtta517iLTmoiJ3sKfVexnZoQtOTwKDb7RSHYys02eSIS
MSv2aMtuG+cZYV1Q6AxLgbjicC95odNgC4aTFK4RhWoV5mN5JZaXwK5P0SsOrvUC
7agDXMusqhdsq2ONcBTwRrAuxAQXHZVh4SGTFs8VPADIyMpAH6swJZ211eurA4/s
8ZZtFeU7jNKOfUs03YpsJgmeYmGqwftcbABnfpULbbmOEbF8aJfyf20dAU4HG3ns
UpAF9sr0Vz21EhF4Dj9oijaRt6IMgLdyPaPB5jczPyG1uwr+llDiW3zKZv10MKmP
96Ffk7mYA2mkmrhQFIzubp4g8TDZlBEG9/NveRqpmd+tuHcfrBXkcWrDYM6IZoE+
m7GZ372cqhXlZVguZ5HhsUIWodyGlaCjyXp1wUBY11r2X0Em+2JlW5GZzGQqlmUs
fl6TUxZ2Gnt8uIkixH3qbBO0kSeHA+NsQ25w7/jCy3cGwmRMLKB4ivrSjTXSrh1R
4OxkEB0aNAuXee/AYtEkAVAMO4yvipEkKyfCtvoNjPAm9qMoBOjc9io9yYLkH8ss
YWjRvtTja/04LoBnw785nBTwQk6biBXPOScHz/KGvPGgyj4E4bwzSpY607WEJ/fU
1eN0TpY7kw+xUX8MFBLsNpOLnd4lxy51uD6OE6j4DD+7h0HDXe92tFXrA+3ZAimZ
LR+Wy2jRa6WVYCEgcxHMjNTTGYnBAQ60rg6ksLzSHYpJe3IPCvaKqdb52OLdWEz5
r9R2IJUnQYxG8honsl6JkfF9cFjXhlxrguLXuQjbPHuWnnGa/B8wFnoUVs2HWlf3
hOI0F+pfI3VTqWJKVIgIzp3/7NiqOpdwH0T0qi8O++F8u93ag58I3be/udwajG1J
LQJUZ/fcwjELID+kACuus90+hJEgCdAXau5cHel7SUclWX44FJeDSqnwq+gQ9SBs
FfVDjgtVbGvFRHxN7jdcnaaQX5ziAQ7+M2/KLs3/0njDrhJ8kUIzqyw48+sRPC7G
h4WHhF2MLVIXb5iIfmJWay1APlNBgO/wsIpskDPxDAtdiDDGGSFTSorbAYDvGFRq
6S/ZCLX0KTUr1EKQbgZJdaooR9Feup7UMfMJg4fSQzE76Dw5GxDVjCSGnPH4Wbs8
u7I0Pa1qWVkHfjMaeNBRfRWwAJSpm/zNXONSON50a+gc+oJ3rhsAdzTD+K/bP5oH
kgbXXFz6bkdwvN6ZDaPCk+pis2NFpLNABvdNzg1MP7pOM1a8QaCypErxMXiPA4+P
bg0VYB4KrXDUb7Au5ugKKQzpnxSJHSM77FU4jpDbpV9vuuY8rGHF6BTrE125ei1I
mqxC0B+GyHtoN/LEg5E/uNTMbrj4ZrTlu30yrm1tixpNHRU4JPr8fp3qVTSffow7
8YoMDSvqGORpDcsTrv4ymtdRqkOuzevZ+JlzNuQFBEaRrzpTiNKO8GpMCDDEQ62U
YtPslgS/cAybUkFUnodN2tCj3p5agFplNDNfn3Tf++ZIZf51IE8R+gNwrj85nEgJ
5lDJWM7waie86urjmSk6xrOFWnX4CI0OC+6iVQjY+mcFSXGP77sUwQDHya0NGZLO
mOX9s9E4VIl1HjZF+X6Vrv9AKJX5ZIE9En4p3a7njuhwY0pfroThbClxXqlMhAXl
cSTm31iPCD+C9HxwLQXEkOzwNv8tiuXrQIRo3fs0+RC234H8PnVvzpHafwQ1yZEL
zPUlqF4+u+08p/8wW1h7wE5DujpzMfPajtEXgn2IhNbtvAyHjSXOz/geXZ6ChKuU
1orTudU3ieCjZ0V1GNeeDqm0aY3dxzYEXMA0TJ/F06F8SNNzjoRrRGHCnbjMD8BY
PVJZkSrK/pkOlNzDJWjJchQKHmoX8K+q+QDhtw4lXm1iqShEjz6vmKPwJR//BhQh
82UxiSs/SjUB4JSzhtsuVLnTWOqrBN/zagykkabTHDHBgUTzUF5psDPUkV38NeD3
Aeukddufoz4Fa5Eu1TBIos2NZShAfcjvUW7ExfhdkzttLuifKlDeebkDO3iMs4lf
hyBTK8Ke8/pb31746S3zVnmFDrXJBdXDMJTrtLkJ9O4Yv2NaoOwwW9yQi2XoADR+
wEo1FkQLAMtN9KY0VMTiTeC7Kc1/yxapH94Qoecmol8LVwvAeig9a/h0ALAeYU33
0kEPUDyAI2T63zUo7UlDxa1dZ1Sn9evX15mBQAbcRVDQsapAGd0ndCw0KarLOMml
AdjFoPQrt+YHmpsnpIGxAu/NdDmqm5rrMFLHdc+WCPDzVfcTJ9cb6Oel2YxOQlam
CW5ra9ds+VU5MXpng9lr/xKCKlPiGMLKJE2wfaKr2IQDO3+f/bhAWTRFgXRkQPYR
YTpDaM72I57rNJ8xaj1xLc2o/B7arnR9gn1glUKOmhPCYN0cdXVZvWd08hKVFSx+
w1zRm3iigtai8Z6PQHE+1WyPTV2ULmQ6Bac1nD1FZOeak11enO/CcAIAQjO9jLo9
omHR26QI85l343536xGh6/feR/Ts6udiCz3FSgPfVZ9ZNNhhWhkNj79e8kSsU0sL
eG/OxITEAnrMUfs8YGH5UoE+6jYDmfd9I889cmzsOeptpRxdZVdc2aORVMnsDWIe
cxuhx1mnaY7ox4cgErchuL5xt7+EJqWk/AdS74lW1u9gm2KkMNZWPwOHVXQJXhAs
G2Zk8YCtsz2FQ8EJ+KgtlcPIUq7IhTEsienBQWXKcvc6aOK+CKGhGsL/Ae2tK87h
ha+6NuqxjUxMJyxIbGy+fIFUHtdfx9qDv0ybLjwTiJKpSkn9WnmnvHCZT08rWaJ6
zjPgAEElbImLHYWT25YoMdx70xwS9chV65xYBNLpHCZiTrNHq4gEGeGsfNzVWkOs
kaPUvw930wztzmyaQJ3O9JD1EA561QGexwIMyJx85NJhNvlyAruNTJ+L9cXENuid
Eh/4blttveQVpFCBKy4uRsPhVBepTLNGF4rZ9MzVJGr0b6DQ8b84IBdH1h5UWPki
UoGwKggPvoZjLDEzhz637wTOzl26HaF8K9Odpwbp3pC5mMf5+YHM42MJD0wpN06U
QHRxzEOCyHXm2oUIaFmm2MZ6oyhJTU7DePzOvSEbP1yL6Yv3NQQpDNaJoLoOUNvR
bRCo9/q/hK89MogYij+jrHgCfk419uSntR/vh1YebAFxiJdVU7nrmfKMefXrX6nf
YitqfDiksJOAq18hOzInDFIMpjOfAtAHBtXlStT61Mjzl7k/mTbMRyOmv4dIF5x5
DEFisHMbdFHTi0XQ0fEOVWTdGLmHZy0azHs0CW8OnLE0DvB9tf3xNhhMVLdpWGg6
DZahDgVmy3RXwzwZtXrkh1MU4nTqm5Xvzqj70Itun9Pz3dcIG6otml/WME99/XBW
gWudFRQkUre6D3HyBmWHXJeNGPBWPZVW4fENRgrMp+4jS4RnLSoDPngsHs+IOwFh
FpXMfpSvuMQfjDyhHqfs4aF5ZoVBADnxg3JQhTqSF+LMmQuAGKcHmlQR46Xv+59x
9VKel3vUiLbYZs9YJqbEi7Dv5QoFDOZ8IuoLb+L23d/DyMN9l3n1J8iPvsir6wn2
SZ3Z2vnC/eQP3CHJUucFOAFhtd+HSkwvsMPTuMM6VDNgkND/etvDdyM05NKsNZr+
Fy4e+CA8aNj2rFTpkC7gcSANLpYgA05/tDK0iMxtZPo/fhiFejdNpuyHZo6s0Kh6
fYdXhxPIwBE08X9UZf2LdLTJhPt8rCHRD68ukIhCpBVy38P3O9l9Ae/hmU26fE8B
E5hIRaWjEsQBk3RI2r0G3ZLq9uSZ3cr94ocdEBzStL9lge7Y5fRrWXPDwaQO0AF1
XPe/1xSpuY6266JM/0ZrqG2DiDdSkXlOMNzSUKfypsHgQHxitSuL+kOlrp4gvu+H
2MkoX2zW+KKAMeB1GvhMFldTaIgX6e3ga9HiMXborZzpz0pdDYFZUX1SZ4nIkKJn
Kph+y+9Qig+cPuygQyE1NzyEXPk2i6pLP/xemln4TkW8IP++LTi9skZQd9Fl9ICK
uw9kcbjBxjLEdEYkPIYZEyGWYnvZC9VWPGf0da3z/xVumVRZUepClpsVUfCZNerK
R49z7yY+xOlMqetaTfW1yo4ePX5u8ziryMOosfJ/WS35If6JQjIhHpe8BuXUhLNS
BqFbOh8yE+hjUJoowmiIg3apJLpkXjZ0VbqaXINLDX+FCW52rUxmydp5JWQmXE80
lY6vq6FYsGtKlOdmhyf6fdfb00M+nxT7AkzhE36iXkbMsVCahxTZ/uIiUlxU53te
dQmO9IVoJjp4yEo9/y7/iwDx+b5hJq6rXJRpvemIUDx0hjwPN3+6PRr2ihkhvjW9
gx8nHs0L/9OIBiiwMPYBUeORQFsSlEQmGQrvfXcR0bLBNH48tfzeICSrI2E/77x+
aJHGLBnKtHApIuODZczWI+IWeeTk7s0c6Hgsp4jEWo+Bg461bQHdCA8bzN2xqwLX
pn7Tm01rrEqGmHxcWbtF4UJxeSU0euIjsj4qvruW3m4sE+If5H5E//E8BU6gMJ6N
YUKKbHM1Rx8HM4gEZ8waW0I9x/xJaNsnCSa+pHnxSLoOhP5VguxwV70BAm2aCYdF
zevuYKU7OukgBkWkXGidqINNlu586yyYNx/bcoAxoKJHIJCVDVZkH26f+xGzZUrs
x3VBgOx1ukaYJurap+ckzBaRdnZBJBeyNQ/wCmZ32t/vOU0ExYjATgDvJLaO9l3u
c0WEYU1HWp7dKSuWwN0tsAMtcOfCvT7kducpFIn2MbIG7RR+JHRqZNSEXBZt8VpQ
v+sxl6WcRJgmAefSuhzer6Y9Fm+AvGF8c9lvU4xwtVx/Kt76g4hVJ2lzp0aeS8+q
MZlN71Y5Qv8ld7U3dxa1onWZ6NtqdoaIAq2KECp3IhsJ8ijlDYbKnzoy3is7iWPe
CnBxx3UA/29uaK8icYla73wL83EQE17SZKldcekWR/wzlDWjMeEA7e2qFj/1ciwZ
C+eOH+Zd5evEwgNZoPszkqFXzezWz4wDRX5gyHcj+mGbYRYn0i8ed8AwcAQIopKe
Ky7x35mLrhdkb2yN+cjqxbcR6cXdNTpO3iUCy5A1wObnD2zilt7oejjZkrWT1WQZ
MG3vFrt8hZfMBKYlhiZqiOlwPJK7jmWBdsZBtFfD5Fhkk73xp4KrbhV9kEpfkQIN
C0r24lN9jef2oh2zm2+sfNoPFD/Q+cXSMct/5U4DkUxSS7ZcNczuvD14ua7b8zVd
Jm0X6FWr2d0032Mrr56hBh/gKQ3j+XabNcKI56+kJNmED23lTyDXxdjBqG5Jo2dd
JQp2x0OXBUQZtcfrZ7APUqIngjRxlTk42pEvfJ26YUl2/W3GaQeHmTPNLhL3TMr8
bxVGFOY7BqMbyRWfkYRzkxDI9xoTiuoIWxTEo28PIEMJX7Q27fH7ft4dzTZ7ucjh
UEnA6MSp9bf+zTW+JtFbEvrFskLaQ684dqNJ8ezKQljeaILudUw744Ig3EP6gvuD
IsTXpaPbMqtsQwZV5M+Ah7EduClNr2U0N95gnGDLoQlCpc8zDSgveOKpBGUq94At
tAYHaamUS6Tgo9e2G3h2c8CpR2jfsh7bwRzDhMHCmEZe4xq3vjE7DeSxiZD5SRkj
+8fqCMbMlPVgRqUrbpdume0z2VAV8CY/DqOfK6ECL78Wn81wJjCQazFwNJGb64dG
zpNbKkbB16PYW2xMUPrJ+oLegpPQmNF7u4wjJg4MjB/BgXX2sHG6hHNG74ufdQQK
pvACMHnTpF+5kocan2H8rhidtvsojmpQz4f1eyWjFWoLlxSJCYgiDWPlVlPSq773
ZuWc7q8ZbPhJ4Kuz9hbsncVPF+AeDif5PzjpJExyzalagRaPrLi7utdEA3hOY6yn
I3IfToEEcvkAsC1vdXt6VII/rIeg+8uyIY2uhoPp1ACmvSNbulvW3S7/bLxihJpE
v8wrc6tgOizLRxmhrgG6vEtWWxG4xkEVxRJgac0PoSBUzBAYFlcnAaT6ya0WeqzX
bjvniOAYSh2zF6K0s4jOp8ZSaOjAvSdvMzJh/VI09zggj/nHKtvEDi8zpN+N4exC
ZnlWcxZ3Z/scYCGRF807rBF3iaumOD0RmmwtsSCfstPCzKhlwnMsUs8xB1LU/PiZ
PN3n8hf9tBL517T8uECNIRIG8zRc/46XdUROFBAr1mji99i4BOUzfwSDRVkIEAKW
GC3lcL8Ssqf90qCdk8aGRnE3dZapAWnDUFLsEpQC+3CtoAcxiE5f52mg4d/UAM49
vmpXPpvjjn7POXWQjPN/ACvCX9j7BKHrmJhYsxLf2FFUgRg1QzhNQSbC/G9V1lty
95LnfpFLmQqTuDCReCRHCWUT8SB+bIFOzOO9PuJJm2ULQRb6Y2FTSmYUQaoilAaZ
CJGdxFegCYta1dLjvv6O4APUj6StE2n7WpYrynEV1/iZLiR4czMVHLmY6p35/ymk
IRcexIIA8/0X/uxQSDS6U2n2dfbTnJoy5U7JV/IHc7ReLoNnn/YRMjlTr++kCrr7
+resrBJYHlADITBHfRYl69dys1TxyCOAEXySrNFgr2BzlXk7lZKnV/JHIMVxRpN/
+xkROAedxv/SQdlMxxZLVPHN9FRiZDMlzxY4qqrBeEkjUQ4yRAJoXiLR3xUWIv71
UpqQctGg1nHmDscW+qhnFmHgqqt+qj25GAWTe8RG2k9ZhMYso9WXB9lMZXmDBVaU
KODdB6qCXE6PZy0NmXx//s2prGcUaLnK2Xo4bC6ulyEKxdFPrlX2UPutjl3OijKQ
qlmBQiJASB29yaiJ2JyzZV8MunREKsAguoKchZQU5xNIjkzzyWi4PGgn4gzD/iY6
5VZpS9XG5ii27XqLgeR0JwpuCCDaqlu2G+gfGwf0T3qw0nP6BZ1vfmN1i4z6mCMM
1ZyX+xuvnu6CXC4IAe3zjEEeaD4QiuqiBZDhYSoXETBq0PK9Wvi6CyWTSG6KQMgK
ndJL41jnVr6UMiR4T/+GlwxfuuxyBK/es7LyPK/UZiMmGaRnSpEwzhfkNVS71suh
5vXMLiwvxkcj/cMbddAhC59yOUQxNQyLhd0d0nMdaO+5fn3ukVd7ZiPrUeRICdxC
6qG6VrJ8KF5w5VLlaapLmmSXx3AX2VVWXkrfMWxIX4J4fYjOodJuhoi/3TNIWRvi
3SAfUHGa298YqfRU/m7VgGhv6X8ItMpTpRscWW6mh8OTrHUW9C671XDMzfzkgwgQ
69KpQw50aXK4xCWOdtM6wEpTIrGciJtyvWafbEbrEg/l/zN5yIqK2McitQx2DJ0j
plX5dxgeY8ubGlIjQtjRghWI9td8ofrK0FZGz4ur4B/8OQ9/KRYE7CrqfTStSdS2
h/kgsxfPLbWVI/959HclVNYywS2MbdVOVCrtUnw4pgxjDtOeqOQWtJNy6Z4/rVmo
eSnjBBOvYJTt8XDHd+cFM/036r7ZhFfv9OG3FTERteeHKqGIlJO9AJQCqAMpY5kn
y3iWVyMyHwQRJvpX3lPboXJy9OeN8axqqEUUbzA5B1ZFPkky3Z3wXLtOkjOteKpV
dM5V7psHnco+P533iC/qBwxht7G/Zq28tZufVlNzChFLAFsGVYS53CJ2+H8X4/eA
6mn1259Ma1aRfB4JHB+D1eHMW7Z7Pq2SXCL0AkiE3YdX77OybALjim5pSmkTfNOo
wGKEozsUDvf0MVs97am9G4kldP4t9vcsJCUKvwm0D1i6qcSDP7DU5n0AMxo2vzIK
YCvhW3ObXeGjEkhRN1Q1mrgYoN/p7fr0UnF74L8drBixLftuqKKEJARO/CuGe6u/
+I0a4Ed1KCNiv55AXfDUbCEVqJEzn5+vsgGgFKVLue+oBbd42yHIUO/u0e3KalCn
1uKVlJJ+LhAxcqRps2wj/pP2IvWY0ZdNQ3wySA8FivE18Q3+eJ9MIW0TuIf3jX98
4v3ubq06mj6p6PhkJu2z/sFI9Tze2+ZBcdKdS3Fo0o2fPHZYb0sTyzAE5X1c26XZ
6RxR8quGYigh9cveul2/94dj4kZKdZ17Vvh/8V0dCRGZ9i7Fh1cMu0disJTrv2/D
cQS2C5ckqtJAlq+ycIbjq+SzX2xSwp9Q4xtBWFQJJUwpsemQVJJxABDSPXX4d9LV
Kbp/Lnys3Z+XF0zpk2h0n4Wr2nyJf1Q9og8e3GnEl6bwGnm1XStCd6JvcJgzp3yQ
ohhY4D9BUcW6qNxkJzwk8At7nul/nJQkwB0igxrNotFL+tG0etfyuQAReAO+61Ic
aW4Hn++jhMscgm4xYgslo9wd9lclTUInSLZDie2hfayQKsLs19YPsCRmoffNUkQ+
vB8+rBRDnRW8evMybzIeMJZkUVFBrtgkjhLvjtzWb/XDV5H8UGIhYDLMkm5yA0P9
FZ9kk3t54yySqQVeOstThbgUeKNzVNBPrvbMOa70mZV3vlCPhRjV+vRm25T2qm3f
et0xomHAjyfsejsD50uN00chVrw5HRgyx2/nFTqJV3abkV2xiEhDdgQULDOTJYpz
vLVQ8m68PABD4zbUPaYU2SlD+SgnnLc6Dn3ID+8R8GngHOowJ/TysbB5eMXcygoq
ZNnxdgQE13ZEb9pHLS7DWjxU4TChX+AciUimRaq+3YvOSh1ozf7Y/Rdd1JsJsTPr
Bec5eRJD7tDZDCV/lYfhDHNyPaBa4Y1zzjK8bIX6+zFQaJPte3kk7aPAHNoKlfV6
xQgNHSwj4RAE+RgaUIJqk8ANHBusj86zVjpD6CerjZiEEaOKkaCFKVN1RkIoOB8j
Qcljet1pEAuP/SISwrPCq5gcMonil/ImCl9plVMb4ZI5fwaOMKIL9ysEkvodFE1i
EgFJiv0nXdQ3Mk5mT3uOc7ziATaCk1JhCyuYg4j14G0pNL8qlM9gaoJKDn7kZZUy
1ckk1AhMwYBfSXM5v4PXaE2GOF0xnkPbsq9oTD5kij8vx0oVVDrtvxpSuQ5XBvvQ
yRm7I3EQiFUxn8S19w8EIH3ocduANze6RV8Z583hGCzpZbjWOD9FNHoyEpRwuYwy
BLDMSdz27rbMvsIB7rmvCzAWATcEc++5Dn6xc7eI9ch2W1lmPHqwMw+C0UG+truu
OfH7yzabswJs2UKh9lqwU4BIuRDzDwzRAmWuACcMfW8yYZMayxmxBNcyqw+saqrp
mnC2cKOaZFIRIjRVsj4Ilv75xuTZY0/nptoy8G8NQJ4rJxudJjmrwNOkbHO5Du86
tS/XVkySV4Gs7n6D4lyjhmPGIxHJ2aF7GaIDJjHtNpmvaPsbpZRUWbSIEZXpeZNy
0uCX3tVZJtH2NK/N72x2BUl/iHq/GN+Ma8CI7FOuBOIh4z+577s8+mvCD8xESqff
+XW2mPvkIXHQhLAPnSi9InfecWezDrxq53Vi0gpvs0WHfqK8/ISZbe1YRtv7zirK
y1jBIu71/K8pZyOTNy2eK0/HKt6NrnDNCpVFzyji9aDD2TM9Z1LG7syE0qjVuodS
xeDC8oMrP78krP6G6y+puOmAuipiiG1lKLDJKLT2gTD8qd4cgGkcEB3fzVutRPp+
SBHqGzV5ey94vJXbF04+5u68Xc4tHZ0pEh/sgOKgBiPi+wcXkkKX35uOllohIbPm
hkGLAKDoUlDLBbAHpw5f28NymSkK73+NAzZtR884Tm50+NLNQZsxt2bria7aQb8i
wAiE9YqTdOdqw6fdMIEbfUpkavPdYVDA1bGq7MKC9YLk7ByxQst4hBY1cREGz8Xz
P+6pHtGjY7A0P4YrQg29uMINYy4zIEF4oW0D6jZrhpKBOu48/CDHrVvsXM4gmc4P
8wBpAiaKMVUUuFqi2MeNLTBw/uAFnXJug+38nhRzsg8HQLs0mkChUTfgfaHN7SCs
LJBd3AMGJMgRrT/38pwBYC4U+dg6b/I0kVLEoGwmRhR5/PvJCQd9qCubRJFxOtG8
z7OSdCLPaKEDOuK4tpXOQLg2p0YcCZwdutAWIBh8lhb5SrWU2l1oPsgETz+YIngP
L+9u4Wf+ZHgpasNEJtcjd3UVZFLgP+lPgQCS9DacDIEFX/DP7XFj6PtTMdWFNonM
92FvMK+Jfy1zL08Tncae6NflZ+gX+8s0pQRBM0fsPI8osPX2nHY/GqwK1L+vEBuv
Zl37n9KFmDc3w8ZnOO72ZXNuaHRVFVa8Y5jl5I7HRHKOaDWTS0ljaC8CGWnnrLGS
XeTDZmRHqTZY+huMMsKsOKonzR1TgAEtfDQXFrFq86q1aNDU6rqR32paqr0Q41lp
X6bpz0ksQUE1IMne5tTGAhCSMDH+LtAv1A4I8tSct+an5//q/9e5fHQrX2OnYINj
OsofmFaL0amsAzugz04nzAtKi+JTVFUv02fF4TyPXpef/dqS0GkqtGGi5dJh/Zeh
9E9VHGtagr2sm9oukpLw1dkZu0eRP3oVnUOcqfBeLZnIijwoyOFaN6X3D4Xt0KDa
uKVEg1B/EyX6H7Jt4S9a+uWFMAwQ5ikVS4b82PJWRCGCUvS8vx4g+e4gY6eG8fX0
dOTJ4XR4npU8xGg2UHbHHraIN0tLLX23dFbRg7oZ+xuGxoZUBKq4Yjhh01qLpSzh
aMqe9vCWhOHz9+S9ZszNGVsFhuDA+Vx1g1RJyp4jG6cceybjW2E1n6ZC61bZKZV9
hweFCgg1jExJS1GCmqq9486YvZ4yo+DlfvjxFKUVwNT9M3DZkHr7tTc58omVgkiA
9vSymSy0lblUPDsf835qSGrqgTsZraZEt7HTAaDNSOmZ8TpT/xrwrvd67hSotMjN
RUrkZG06dpF3aqW3KgrVru33nOoSFsOGoCaz2XW7WDCYwkA9MS5eARtEu5jd5DfR
CBh0afubwcdiNCxZbSuoVjh4ofRzVEnaIYQ2RdSLcIhJXUpNIx0yJDzZIEJr9wBQ
T/F97CbwlHds/q0YmrTtgyelvlmW2ZrUoYFcPMkqqQFLR9YXhiUo3JmTbG4pmQh2
2pstTrDYhGdy9UGJyDS2FmfsQZCP4xiARRCQU3a+T+KRoSqLTqnVXtb+6rFDWRBr
UvLpSRngruGzyHWOhS2Y1d3lYqoWCC8ZNQ0ne5k0fam699qrlzM/9viPu6p0UlVK
KvnJk0mBQcs6lRu92rrFf7ee4c1A6m1kht8c3U2lMJPQZL/XdCuU7hCNH3qfb3Rh
JiMjyAVwSlZ4BZRm5EUC5HJYrKJVbmbxGYTOzjDkUg7sIXT5N/je3BHvIoyEJ7sj
SISeQ6sYLras4nlJtk+8zKBKUt8q3ZDn2E8E3oSeCV9GNkyAvWJ5MkVUdBDkGC3E
htxaNbAEqregoy6b/qsGaFF8UVrXQBoIsUHW8RNUYleYuOxvY1jhCqe6F5Zaxh/u
ql8sYFYZqWbqwUPmSvEobJwipAvgg/WEnwLgxjeKR1i3dvHVU8Q0A/u9DGDwXfe4
vkNywcbHOF9AXOXauNPiTdjdih+K06nnm/LCQN6uL5z6+AKIrYGdWA0jL18ib3bC
vrlQSBb5WOCLLk1HgfRvxraEFJH6pOcj7cbNcTd6VGf91cisi4cJ34+VLBOtJ5rw
vw8xDDqG5sCAcH8b8VogWtsTHgOx787Mof7Q2/3aV6Ooxrlnh+hvibKaFKGJspi6
ucV9+ZMz2sIf+urXKZmxtTF22VxEo0tJC4qwxxGu2mF8l6WMdp6rTB4mbXHUsxaQ
LabSw7B29rdbqQFY6vnjE/ZeErUHOyRBmv88JW6dxxWGLtJV1va8cUYz1geQ1jMB
lxQ9eG1jHmyYWfx+64QZmx10zjPfH4CLxkO+lbxCKExoNUSoD8X35gw4xxE3Vh6Q
i/cFtAUIN48HZ5V3rKlbYIj0jG7+XqGyanqNkPnkhKpA/mQgzCSQ6gbathg/SvK4
m/NtNG2LdHUN+jlbOGed8vQaNAJB1VdyOSFAsS1Dz+DcR31rvFsa7GyNwUAXnbml
YCFXGIu7fj5lPLe43EEsja7enmcoFRk+v2oAQyWkBR4gqqZT+KVLC7fp7FLCsgiG
T7GUTdM2dOQQPYLk/XXvY91RZRD+0YZOZK2vhZYfKN3Z8ce7PReLGJPIgs7ng1bb
aWfxzXLUvmgVdVX1hettGgRWgM9/m0K3VnCHOtrL2FBCVfkT84hTLMGiPqvFIyAf
MyHN5ZYPi/qKrchi35kZx1A0DjK/a34GXFfzXXtRYIYNcfMlO/NbzOjcYmwAdpJb
3CUB9ESOi3sqhq4Xy0gHawEr2bKclgTwnY5/dHZ++pHoey0N6Dj4A8GZeFccXyj9
4snrkr0w/nhCgVLovWwGGL+PuIP0DcvhOSMSrOzn0xAr0MhkF7WBuIz/XU3qmOHJ
38E/Vk36MWj3nUoUv3AvGVQeG3XqaX5acjC1W5mdnNzjG665SeEIRcIT5W3gwym/
16ILIyqxZBp3Do72w9FsNlOSjdrDKuR/b8q2WKuPKxggv/yS4X6CeoVC3L8jmDoe
wu67EG8GhgsjkuWPUaUvxfCPw2GbafFOxkHNJIM5JTczMoZ3JbBxaueeU9lkwEn7
WbEyUaaNf7uGsLKbiphFKuZVy5doWb3tWqdyZqxn1hwNOzJ7H+ufIgWs4B4rmKo9
znbBUyKedrQ4hAWRz5psCR/53PEyskmeZsQBMa0uUu5BP9TheNM4pRgT5D8Zq4SM
jEuZk2r/KTQ9/cydZFvKFeZXobiy3fzhHmQgCCKFQGNhYyNpmxJcW/PQB3MqziKC
iLqEtPgq3enlYbh0bMdk7vIe/euOlD0aMb/YYvwZ4aA4WE+fC51uq5CifoqE/4G/
Ik1+F2aH7r7ax6t87wBxJtfVyax1dZUYNnSicR8WEVuGLTGTuiChkqcZ8DGqLvqE
aGIrE8GkOSLCJi55J2tHQBN6q8t6vaQmcqcjZYIHjUH9HM0XGE5vivCIFK/yO1CE
RwE6A9MYkN09YPadFCD4XXLVeOgdlkddssiz2S2gIWRWuPDzxQDWeGR6YlrU07Yq
zNkhGBcAns2Gfsp7NA8A8XEIYePX19ICTnggm306vWsGMrNGjQzggeQGzemvHeLH
7g4wqe9mpFAJms9BGOYXy38Mq2iYQMX726PEyORefK3/tdFjUbWyYZ1Ejbef0QCv
5/8WzpO3LxWyX0O6neYVkb8uarOCmq+IsLiLzj9UNCuAr35l/Q+oNvnS0ajHv3YB
gxKh5rJpD6Pvn3dF+cLd83wpJSarHzbjhwHtGa3XoOtb6ZIW7UvoEpYKX4fjxKiA
+m/sZ3p0PvaGzyPhBhS169+QY4HhzOkhaGJXwdAykirG70BGFQms1M1Y+uqqAhPX
pA7gq/82e46jA3tnQ6GkkcQCnk4YVslUp3rgL8zvGnoMhvxdEbNvT8SWF0n77Vr3
fQGGKylgFxxMOXr+CEvvjFaURFm5W7QVA8wrzazxn9Q0BnQTvkDTYhgS+oiJcyxF
lYReIwpc3zKOGKWRa36dslLAOn2GiJTQ4nV5iUoYGf13ENmrlTPn/i0hIMGV80hW
la44jy7JPnWxoc/ErAmHmXZev4TQwyHbw+XCqkO7S5zHhmg9q5VZww4MOuUHQ849
66Qq/Xv6Sxm4ebigvPzlc3wT6o9AcpdWaBT2y0ymS4Dv6ZT1vkX11qs5INh5lqWX
QkBYK8r9ZtcaFkiDdLJaaID4gr8BzA1OfXMsnM74uJZhDO5MaPa7n7P7zDxWowu8
dAt1+y5f2ihoCObh7ziaqkplwcJMagjYWuF4S6gsQVVOljOcDVGoOxz1YVIFwbrX
pE9FrNymP7vAD01wrytWcEMyDVPBMUAfuhVjCv6cRQdTR+IPKo/nxyzD3ObacDd3
h+Q4tpjOycYm4vXg5XnrkX/sy0JguTMYOiDImRL2JhIfMvBXDKJAcI7JIHs34Z0R
AI6PhGTx8Zh/QBsqjY3HUu1Luqg+6f6ZPFufxbTHXmALOLAFrimSvCSMbHS/Jde4
3k2QxxuA+RW8W+nTVUGQVw2XdWq0U9szk40e09sPr6/c8inuxuCChk4rpcNUxiAQ
bAEc2Ik4etUtJVhaWsGuD2LcytbhYBtlskFj5/NCVbn0qy/SYfy7RZ0yS3B47cD5
tdnrPT3RTize6xRKuyjLtO0hHbJh00XtBarDgXAjz3k76Dr+RojifgFxArMveI6/
GZSNjS4YP4ectj8jcHurx62bhnrmg6gD9kCX66+r82W5WSBDjWGs4hWWi/f2r1Rg
htaPF4aqmA/fbbN8G7cqpA3POogvjqXNqqIW8yx05x3kcprzpcSaBnAVOhfUGM42
/0afNh7pPMI2+eFIlTmuKh0s9oWSJHpmR4TebYCRhbRTBrMELzJONdB/V/25czLY
/tHFp4Xw0fWTD8f87eOp6Dd8EXchHLC1V7gHQ6exHsM5mlsJ134fn1gyGD3q7og2
Kpw0aJZZrBkY1V0zivG8j1efXriv21H7ckOh/fUvJxzQ+T6qC3cHt/ZWvg1FZ/Ci
R4M8zjbQCqCd0iOUFAMrzXS/HYkXfgz2nc/+u1Ni/OZM5YuLaaeH4fvpd2JiDn7t
fvM3BCnPOUeNCnDTPwB/zL7irmktiv/2Ttz8IKNaO12hwkpVoJg5ygA6ojSCcYBy
jynhaoabZjQFlNlf+EDmMX/zMh/2k0loC+9Ju4x+2eF8mAifzViZFYNDA4++cwX4
YI8BZKR+0m6EzRBrRd/W8w+PqlOgjxCOONRAbAzHYMZKmd9si7bX1HDiM1EHNvT1
hUIkeVr+TJzobnZLZKZxgQWgwu1Af0MOoSgoSWTXZsXhDK1Pe5OaSRTNUWjo8YjK
qKJiRQVFaLDWezSIf3Lziwdhu99mrgoG5Udqxcq4GzhUYuZAZK08fgYrlU0dgoo/
VuK+Di11E8sy/4sY7ivUeX0udwtDiMVUpzWeYGpTNzv4jJBALor6pZDJg4rrSTFz
q80DwO+3yHzXRAhv/47qr6dkFWzEaeQZwWGQGmrqYNvMgnR0AyI2B5rBNwBKE4a7
XAHUPNoLgqj2aA/md6D3xjLzFGSQBjXrG2YJDTxqggg0bn9Av582YBwpldpdjd0o
49Tzvoo+L2thSgYiAflbYmxruI2ecIunclsyVSIJy5apUy9PjlfBt2FiMyZsvADh
QXGHVKwNgXvwxUVQnjc3S1aoxjwt/5hfc7pqDuaR6s6i+jaM5OHxmBoLb52aqRme
tqQn/eeTRyclqlBxOBEcyM86nH9NvZWPJB5s/VURI78/sEP5jez6JIL0/PX/q2jA
0nY/VZjI9ZQtXw93mpYEsZIQdsgjhjkHb/s+7kOAKhrqmJ8Y/Z1dW/gE76Q8U3K1
y7MKcSg0WCHFL7QXiwuVmK09/SpdPxaUZ70mWph5fBqJ6NAYfcyN/dBzDe6yzC1Y
XXv5Bf9D0gVts+PNNQqy6uDmaLRMVvWwN2lNUsXg7+okyt4WHcPT8SCnA8lUFAmN
0b2GUL1t5MaUa8xLI8FX/l+jIcqkngNaOBufrrEdBYOJp6l0Yeupg735plPGJL4O
4dTSVlVaZ1gbhMEZqKf/gIbplqEIdI/GD/jIFStBNKVLbtiomL2PVtS4wZMKk0aT
5rFsYV+WX1BGQptKDLggzNsKYyWJlAm5xZ+SMxipX8uhJUXw3l+xVZfyaCaAXaa+
cUmiBwcDAI2ookMCZ/CSi79x+4E4nqzg+f/L2XGaHg1TBO6VYp6QAOMuP6Qm9Zvu
HPz4RoNRdEAu+pGB1yNPkYBqH/C1yPZT0ZPCzDty4Lb+QOuwaquYtrNvzmDqStQl
cIZxl6iMi09H6WZAnvLrkwaWCx+YJCPlmLiLKgBQqfDUsOlmEzX8dKtY9tVA4YSJ
ZhLJLSz12jdYwT3DrzCZhE3OEJyRuwkeYsRcbSbQv54jCs/tGUWyzGJNHnx/D+TZ
hcogzn3/HCHtzI57oE4VOvtnGNokXZmb6AsWqd2XonNA1xCVB1nea8PxuCJuYGv9
0wlvx3WWV44hSyRrhDhigAt3MhMBKo1O1rI/pXsMxTBes5aVMqkom/pMeKZjKqZM
Q781VC9v6LygAtS0GivQpXVcwA4HPUsm+HhIB9WF1qeeD1jfaaYW1WvVUnz40IUF
fXRtxkA6Tm8MMJCFbaEOPZ+GQ3UqKRchJ9669RXMalYiqIqYae8Ckc/tfHhfW8Yl
UAnTIfOf9/ziSpc9yGjvY6mPOqfxNIA+uFEUThFGF5K470EeOcfOUBlGm0LR3e7H
g3q95RFFO4xauA4PQGsEE8+TDrI4VqWzRHT257w4Ni0Yf3489EwZ+FClzAJtpRTQ
vS4ke+GLOR7Oj48DYsDS4sx593KyT8xK0u/gB26MzU1D2IczMUOyyp9wFu8wufnf
YcLY397TvDMjaRI3EzljLGwfWxY7hlw+v3lIUq9T5L+8uQuzFMt12tfROG73h5Qh
EP6xTovgtKMjlL7GnC7gMXhrTgKvxuhnWHpL9b4sJpOA2hLB5wSBFmLyH7TKDpSP
CA3YVD76Y9rCXZW7aubLNs/cncXzNrJ1e3LjoK5wqX7CLD4ZzvUEG23v/0VD6GW9
4nJ9S7SNVSP44UXMpQ4wWMQEucrpJKn+AYeH+8pVTGpk5ePqWyk9bMOdK7JvCvVm
AE9gJfTsu/tWBJ15+rm68gMGTvSumUn2v3/Xi++CiVvkY/6JqXYMnAC3xXKmG3ig
L7JBi4Ej0XXmstN1nFyI7Ds0K5wkQvLw8biNYOvKTrXTCO1wsl+is1+bYQ/5nTXM
0UDSnRsCiTdONmgxFFRlhSuWHz/OVbhcvmV4W7l7F4ZBiiFZLK5Xcv6b0Y/y874m
8/g8lIAkDedNj3OKp7JU8xWeRDBsI9tLQkeSKfTzO3CkauzMfXfN4aAHI8lrxms4
hjTdF56muxQrlkHBNi0U1ngaDEbWqGXoRfN1d6mkd6xQyIghHMqmu2S8D8iSAJCn
aB47SV3uajNPGeWaxsnc0hodVfOTMSexHl3gz53NxXPaJieUiLEOyJ8WXaR9wCqx
VZl3256v9iDyDu4XeiHU44PNcCrjlnt+ldmpk3dLWHTHRfjhGTZK6IutYksa44En
+sfp1V1JlYZXDYeeunS9RPjoOWZ8DnaGVX76KBJN3Xn721LWQv/VxPho2/Q9VKdy
Ii/iggB2wL4jUQj16FgDW/ojrLkwIvdLICsEkUTriA/83jKQNBs9zDz1USiEX+2/
iFkA3t1tL+UcRXzEmggI53U/kE1hI17wnYUj55G+8Nia5Ro3yE2TiMrlJ47uouc+
kmy23uCBtufipbDce08UJcVhhLGNxiGz7iVO3uT7Lk8hXBC0ltfVSwonpVImbejw
c9AG4csRYV3xiu0VrJrIYMoj6THWEhBmL107TG3DFvnmQfoeKjophz5PELULDwZl
yLnRQLtDYtz0XztCgYqcLqOmdYU6atgr92SaGc6OLXL3Mc2KOdewQlN9kWjAp7fv
vf3JmD+uNYs4Y8LvIvCPVAqYJ6SQ3vOHN+UL99UyHABOJ3VOg8V59JNIATyi4LhC
hOf5c8yKZClumHC4GpRYVEgaRb2j7yvYK+iqn04mexp/wcX/D1O66OC3iV77lEyx
GalLeC3Xf86oFwTX5k7vf18m3r9FtPpt68vDIoCOZy1mSi4fpXUyrYmPpmlXH/CZ
d8ESmQnntY82bEBSSTfW7JhklYH/3pc/doxA01CqBC2VVJHC8cTXNFSK9Lf9mN0E
LTFFRK4TL79p69K7oFYebgkvEfzOLx6iQsug7ii353p45Pwj9wsRCFizYZ24Oe28
lY9y+qVlAnV1Ew/Dy2HW00ufqmsktoSL5BLFrQzsyoZplJcN9fwhtV5u9zCcAfqv
jCW4Xw4OTNFzz/AspdcoU5cYKh6qOYniCfqjKBVPUiQeJOgqdtBY3UBTqgiSC6i9
csiydXIjusohwz5yvZTTwvuo0qZOvgG6pLYkhBKVKfj6yPXiT/MjPLAV3ZoVH/Kg
+89B5mrnqoJzd5RoCiyzDV3uA69BrPg6ppFSDftN8+iiL7DjMywEzlN6qxrTlky5
ihcDWh3OiPmefHNnVrEFyKFN3kEn8LjMIP3Y4tMc0l03VVkNtRfRnYY8UJmHik+b
ZIXl+bFHLjbqyk6CydHjr0xDKFbHO2vzQpEtRy2d77jTzAW9OveH0tyqP9SBRgOp
4lW1vdRlYy3P9+84l9DdTGuU+XGIaXF+Z6re/UwkhDFesSxS9JtcRvlbRaSz2nxL
9PplDagY/VEqHxkFIn7KsQgXcqDRo5/8HylQwFYZkkLVYN7dfMNUdUfSt6MMCaA8
8LW1Ba2mmceCiWP5Sh+TNGVQPd90xcEM4ZP+w0MnNv+BWQtEi7Tak4CYmmiH9EnH
G9ab7sC1fBqgzvDrPmh0S3/wU9P2fwwmtAMXxzMkaPRtjIEfVKtWZQC+DC4TUx43
spMOvLdtd1Lxr/8SFLtwTtSsK2zZOXORN9u6uq+/TpKBn9llWXgGLsd/8dlkN1mH
ZoFnXbKXa0tlbfpHSpCvTlNUhq3RzXceiBINTYL3CkZjLfEZi7R3MzQ8kSATVekJ
0oXvdUMJXfCvSoZ9r5jZhxjkII8Iin6/7mZI9CytWHA+8MWYLqT2J/PooUzWqZsk
oqQkjt07LROl0RWhncW915zGm84GOykx1UVLrjhE1Xbv2wma7PPjW7iAvZOww+A9
Am7E03kUksxs7fRpKbnL+phciKZyxURXU302qZKwG4V9rGVtOdlrM+hOCvW/8ItT
BgFC2qxA8vYOgAIp6IkHyl+E2kU8USPH3lZQXdqbA0hMCTgibHKv4CngfAJtOagN
6LnCWYVu7lTFHHxxAq1/X11FBo2jn/dvjVN52OXZHLairl9m9NFPqybS0+erHTHE
FH6cVyX1+ca8ABpLnR2IR6P0ea1PU4I91W649FYd60c3U0VPAwCZ9irvQ5vLFq3a
3T3SnE0Gw4wQre2W83kFXKrYLTDtRYJdMpf0gAQQzr1xlZjPHy/fPe8QbhLgrim4
9xbj//G3Fw8v4917JxFUbExllskFJ+z20kgj/kEQbZ37AWmqVQs7TMYyv6E9Ezx5
tMkclMcihrukggwRSZjhhrcGIukTInwHEThoNE2r4Rk8e2gKVQN3xXFr27tvMoTW
eHYY9I46rCfRbXrvdfoa1WceDCGmvMNErcyhYewk7qDAb1lLzaqCglUMLYEyMg67
8HfAKg+EdIcxsIHF5B3KV9GeyXwepL/OS3zzFn6wmkU15QFLzXJeCgJtkfrzMo63
+9yv7q3QQAOR0DaQJ+sx9DlRjRDF+FXe+tQIPz9mtDR5leTM41GNnKNiM6ItFexx
qOjmZo1Ok41trhVHZNRPLjVvAQyFS9WeyZa2L21mqFZF7wKZl0HmI+FRmPsQr5dV
sx5n53Xly921r/rs+6bx3LiBuyyswGGReVw1dFxrWFOzunXcmLsrCkZzvKamvgvi
x2/vnBgbdvlo0KhnmLsuFo/b47atNewx9A2G3tXM7VB/tG4HQyD+fSbbTyXJR+xm
GSJ1jPlpQLYCtdSCNTVl5TOMkyR9DBcO5IflBh7htWfib5yxKZy64x/6DTQx8fdB
IvMYZKwlF5r8ev/k2FnLWUShYk0lBgx2admdEyetK2JGmv6INX8C4jzjEJ6iGAns
mE5yBFQu3qKzKyIMyROq/6kf4yqAaG+uRzl/n7uWyTeri0ov6ZTHm3mH1s2yQpc6
EbDZKznFyh+89zimJOWsEG10hsoKzQd1V60C24/Llu4xSxZlqjoUlKqlmvmVg5uY
QWaiENB2LRMxDiTrIjG++mx3FrYoxvQV1wzyNUb+nRwhsu6ZAtcbgWBVVsvTvQ4I
j+SpqlDgmQWOOBv7vW4wS5akafpe4pgXPqflXvgbtuC7p1my/D3c/uBWb+VZf0Aq
5523Jo9Q0K8Bm9ih4ketSylgyoIWFWXNodLz9akeVw+2/01cVlgc9Iu7ioQv+fEE
bIYHxyDJ+sKjYyiq2sPV110RmC/nMmmNdslTPwvZ31T7/GRLH6i3ZQCGhr/+lD8B
xNhRfFYuXjWvKzty4obfUeTY0IiScoendxWmXnnLdoe7v4m/6iy4K/eIihdDdapO
mNyIof8wT0D7SK3bUlVexOq2klJfaq2qdPo9B1iUpzhcqVI1Xake6n6rcGkOmgCT
Edqtc6UurXgtRA4mOh7/nTwaFM6+A2gZ57D9wyuCPSJh8HL0yOsPHeqR4xpoQ/VN
ShhXx73JSryImgnPel+1UQUXPq0xtJ2BMhuLrbKxhERHBXiI/Rjz0XwEM5Yu9Gbc
y9vQ3YI/uSg/1CsP5WkgWuYVpX1IJzPsJRxztMs593Lj0riYMByo+KK7Zdt3vJD4
NWmSRvEY94PnPSOQbTWHcRyimxWtKJyhorvvyULBbutgayyKJrKyQzNZp6Nv/K4h
9nnSKhcjLC8jcCqrgc5iWamUrLyoeiFi3awxg06rqG+B2YRSLYVjnbD+Yf4kjz0D
8uLlxBwnft8kQML50yIJwrk3d2vB6VKCerHj3P+aWbf9iYiEArNuCNJWoBeyKvFo
+u/MaCvLRqMdmuGtJkHoDLBHwzUJC5Wv2xNObM7klYbugpVEs2sQRFpGts9PqBSn
h1w2LdveasBGYMSLOeYH0a4neVpF8xTrGCVQzKYqq/tJyVxq6w+37OxxUr+UULTX
DIay18CVII94hoQamO/P6VyoLGCNBnjGzrJKiX0oC30/46IcuW9SpGVksezOVNpC
VPptpw3PcMQQRVm3eV3j+qTCy9myLBy6puE6T4K5w5fXn6UKBgYGAK+qyM3qri8s
UFXcw1V7l3PqC3fxEmNaaFXV7jGKt4VkJR+tBNTRsprrZh3fJyEQNJ/RBu7NE4dH
PIDr1/8H7PWc31Gm4/TFWpFJFQ5UqXCm5+pHXPud10fisSKTfNHV7eVtSgYL7+WI
1TeJG5wXudSc2cHtc2pP0SmtD9v0y3b9lYMzcyuoXTfycsXYZDG3nFpcHs49lxj3
bAiVNkXoqqi8cJbXZN9x1SaaJbQ5RgxepcSfiG7JC9PIsERVbOLLhGVmhO3iRcXh
Y66vX6SWIC1g/R9Lazmk+3CWeaG7vnGr5jeGdGr7aACvi8t+AjA3R51L22j6uyiz
tpFsCi6E2hteEQmZZ02p47iP/v7dopQQI5iOYnFYALiV0SPnFE/HZXgJnrBueCUu
RfpG9x2FW5NGbpkUwLeIXzgiRODSW7FKAgulqOYIkZdmKrOk5luqreZwXyGd1hf7
NJ4Uv+yvpyP7h+qW3q37gOVU2Vy6KWoBEICOZQD8CVlLB1HQXVAQpzd2HtPNts1Z
QiHHwjjcdlhXMpGu41e2APY8Jmw6XKMEbQ4xV661tssPGqWoNeYxm1oIZ8qmQWdN
Qt6jJz/xWhaRjV8DGCCfQefjkaxfAISM8BzzlywyrEN9xrNIdA7hOgjfWH6LRiW4
9IXjxSjUjCtQsq/eePlkT7/nEQl8xWD79NGva9lUJ5I+9GElGCB0gL50t3yXlkPY
VXbjdg7IisMDfnB7IzcD8c+nU90YHlvLkMQHD40WvLFImnUnGSb9fpVPCVUsadN0
9FKtZDEswUGgjzmPuuspaKRkWmOpVCCh+/1g9vdWW0TNQH49Ix0zK8XEoTPh5hN3
xyXMiaDoz3C/Bf5jJbV7wK/+M4vfglXr6VunSkYJFmLKhdJ47em+6kUr5Mp9ONMP
MkckOmkL2OVWDq6NJn5D9+oOyEN79FaL/3+ZreIkxBtN06VESIZa+pvlseIi+lSx
iKeQm1XzhUiBBz8QXTj5Q89ldB5AO8lpqGuLe4VDSwhFDdZhccNQvICOv3deDW+X
OpB2N66vv6o4doZYu7MX8lLD6EiMhNEP9F0sNdkfJrvATi+6BMPot3cPM36VxNz+
EMcA0o2vYRwNBjL8hhBNbVaiZ5TtOGFQkV3pTKtA4WEO6EKbGia+sB6TLjAkE4Tj
y35rM68cWbG1kqtJUCsxTPzBINb6L66dHTRmi6nE6PdX2JHmm1Day/hEekH9dGVU
F1KFmiHvf5GY6s7Uso1V/v6ZqMxsMEGTPKpTQNq9c3/7QzGKe/eRro7hZAos4lW+
w6yjAyud7qYyNe06TwAs92DvigVlQNXN0ouaZi0zUBTWbgWa2AsIxZPIVZq6wh8x
BS4As2pQI10zAbKaoioOtlkRqAkoXefOrxZQgwDq3TkuBsdIT/1XWGGaTnbgpZr2
gjlg537u0TB9ZygzM8cIAEY6pxxVfuv2AyuoPnzswt6tenC5LTLU7oQCG9Ev43eN
eNgjc7tTzb4/+PiWcGc2JDB39iCEx3qtvRT+xBe2bKygfyUgUl7mCwEa8LkzBC8P
ZD4n7JaMEmr0ZKP8xDZQBf/I+k8m0BxM0vL1xFVRMvx4aiwXWElhBm5IBmlv+lZ+
ip6lIVgNLBd+cIb2dE1C8M9C07OzeDm0r0/l0IwtB8HPqREh+z2FkxV137L15ns9
K3kPYHTt4s+QT/z5i8jfET9XpPult64Jx4VRLzybeqG4vHobR/9Nxh0iPkmOyMrZ
hdkyD2X27MtwEDdaK7Kx6gF8AHYkd+t/ff6qyVdsj5ruT5qd5IovWzjEI33Cd6qW
WD4LYtiRwQslbX8GP8NYJhuOZPiPljAn8MRoR+WJqrPNELAee42Mx1KGl1Suqdxn
8xPvX6KByVB3dbeg+yMlKYrlmzb82r1Zz1tjfRyigAFvCO8y9xcXl3LEJ7A54O3w
qG2zFmaCeG6OWzD8ADKIUBvd34G7Lr5nVkq4o2LLzxhHh69rWZlu8sLgEbUrRJBs
Z4PrTZ9FJY/BOtcKaGPCmmqflb/W5SrWgLqDnnW3WQRm/tMJ+iDuWWUs2bp2tuH9
GmM1sT4JKS2dazr2Gjm8pUJkFuF8Nifqb3IGWeBf/A6Cfen2zQuLq+/m+jHIRV0x
I65jkvkqQjbFn99iNCPDhL35uX7yNomWp9rvQ95qpEjtW3MdpTqepuxRGiWMW0gE
fKG5Kp3iIX9JMteQ8QbZ+2pVwLcqYomvwg/41fJ0yv0R74St//sHRL8YsCV+ilbX
ejAMVx/VyZ73LNgaq8RdgRwWM1oAzKGn7n7bzIrIZyJaVMesJyiWGcGz+sRFMRzY
m0T29Z2fvDuDhuRDJZ867Od4OPy9Z/0Owf2m9Fg2e+dRWEjhzQWMdmTk1WGYs1Wj
oqr7JD24FxKT6PyYJp0LbEs1iqoi31TDgZsZLdcIneneu7pOtrhByiR7fLku+PMZ
tfKJ1nEijj4wnv1Bs1jbed8wVt263An8qfry+J4tzFG1ItVoJ35BWUqFkfbmRCS9
vszVuHRm/rsbnKeLORSC5rw8zzrO4cnARjpU0FHvDFmmu/bOGlZDnJLVUMjxRwHC
iHP6HmHPdG6zSYERhf9X/UZ+/pg1x13ikLFPQxlM6J2+YhrV9J9JlyUOYqIeXVvm
oXVKFqGnwpeHK4aE7t1lQnQuA5AszYbeIVoUMtUou6UuaSsjjB4Rx/i2AplBssNx
8NPRT7fu795PtiZhSjgXOyBSUynfd/X8C5wI2Ymaz2jA1w6ZK4HNZWOLlqWDU0Ud
x5TYuMeaj5xzMgiMkKj3ovWShVXV127k7c/xUYKJJh9iaYcQIHTdY8hitgNGfxz/
4Gtfgf56ji/nVWZf0mcT3383BGr5d1NBKPWrW3jiwcfntHlSFswvLRLbbSTmn4VB
bskkYKaFy6fczcLkxX17Lbiy+JXrlBzJC8j2nvzD+fySWK7Gin9EoERTZeJWGgWM
fCR4UQmrYnKFDjxQsDpi+yHEJoE6BmIu5srAypxR8kGusgIDFRHGxasNSZgpZHKG
fM1rKcWDfezfXY/VOMkuyjlJ2wyvo5gahbMj5Z/oZ7kto1uLLRuozhAGee19q4Er
HYU1Rz4YSkuZyLU4+rpHSLoMj7yi51Gvb/IOusLJtpK3Mzs3KWsMXt5adlmF46Kw
cJbEqqX0q4347vrkhqAnwYLV89p9fHIbpvoFtTFuDRjiOWBP13Dc4lXTb3ri4Sjv
aCNYCJG20afrYWAf9RLRWq1dSZ8Pg8GFM1XrYE1HgP8mKGoLUkFjSOhfLKZORpCv
J8WhP0Kx/YBO8OCe/keI2mMEW7b3oaP+sW+NyuFnCkzwWgnZQu3nDDpfp598GdIP
dna/Z9FkEVYXGlObumJP5DHTA8zoUY4FUfHIuMBmbjkCkOxHOj7pKmlYRzOfghz8
cJ8lr/D1iwQhdZ041ZQQi2veZsUxE3XH1T+vjaXV8p1dFUL4UOLbu4WaRXr4UIF3
IAMc/z8iaOjWMka9cPl6RDkj0ZzkGg7dwpPMZ0v0ob09DpzrFqWCIdqLlnLSm1Qf
1vhbOFGySIHLoIDsbHiMZOetgY5eIb9WSggAVqzdCPvdFkJHhj0a9Mxku/hpbe/i
Q+16R1ONICeE/IddFCkBDVmmzkpuHZKN++umSWt0wzVd8nUq2XE/E9vx+JS9OROr
PzfYR5NrqevMJw/RkvJCBmyI4qWUvmLdj+yoRoveN9STrVFkNMJj6EtcRrsAZfbg
5lnhC50FAGKN5v1gQKkHCBIdwie/ogyBfTT2QR4Sp/B07UzUA2BJMgh/GK/hO3RC
ts5xsSXfSpDu9kMD5qEF+CTqKI3HjfKfo692rVRX2wX4BZW0B50ne9u4wb/ySlj/
uTbe7JBDYRqFBSHncGsuoW5iu8nHKq0c0kN3Fut8nP2MqLAKHLd36o25Q0VGcYl6
AjwFGEAC3BYvfFpkrilMu4t4ITJxwMkT7L3flaFd3YyB8+C+PZDzm5BkhsjT3REY
IwRU2Kf4DZWuf8ApUfc12udlKCcMSJJCWcRiXknnQHOiWW7LWTshobCifdU5YENA
xO7HfmWfZjIuVI7CvjQhHL2Ssv/bRP1QUMH8xN1bWNnHXalrZuSJLDpb8El137sL
WZkBEhYn8okFUSLA890vl+F8m+hLXxinnMqcfJSHKX1TGzQnR/+DQsLtwIiQ9tYv
tZhgTUXRoIUQJzRKTrzrmQEBknLjW2pwQRxlqfp6e5arIP+/fC1xOTOFghy7CUcT
cwrQltZQIa8qcng/bSS3J6UlemhDyWoVvsyKxZTcK4MWcSCD1dtfivua4pDgMGh8
wpid2yyrXgtP20+GM2GdE2XQQq/ysDIP/CcSDCuqJxw8TnymiA+sr/ktB5Byx4yf
1p9CHbzd0SV98fPU0jWAfUA4d9yfrhpfuBF+Gn9SYtz8hIhv0s7skFEQ3GXrC2RM
1yu4S5hLM1VWjIQbS75X9zk+whpyIN6pCgRZl3YCWCgX2DC7dpqBwNTblrNscE2j
s+XFYXUfMrWC9SanVRoTR1G+mK5WLzz/gImLcNLM6QrrlsZk0cDV3briRfZcw76o
zTmmWaIlSG7XXY/cxUJdVRef4OFLJOq6Yh10moYCVx3gEtTK9m0H2EfTs1Cizi6C
FhunhWOKQe2fR5ZENONVTe/pkYHXnXJMZYCn0aSfgWBg3gzULS8U/fzar1z0dP0u
8tVYeVAaWaD+2EDsXUisxNg5yIlAEP/72Eu21dWdtQFgWn4F7RhwA1kdCYpSjGD4
Q7vCS3WW6uUikZCT/QXXzoC4j2bza9E8s2XSJiclWjt41RT+IuweJ/R60sd0o6C2
+kiLlSBIlKYNSRHzh7qvadS4otSFiTJkYXU8G2133FvX9GHxw6b+2LJWHx0QipQj
JBWV8mJyMu8LSMZuRP0ZrjE+PLBsY8EFWeh6kQpuAgxowZ5RWGpHCaJ035QpJLRA
bUW1Kjjpcxx0fPyklj3EA1Ni4Qr65Kw2xzxioggIk1oHkiYOFLuhzQFr4xlkk/23
0/L1cicNMrr2d2l8gXC/XNV1MhgV3T08g7p/wFR9e7Lmd/ABC9FKTCctWc+oCcc0
8M1FmeMvFlX8oOwnXjly4h/hiP40ylrBN5CVBFPYth34h2rll24HRobZ3f9p7hO/
QB937yj0aon5NCMdfoLrbJ7+8fYXHTLKTehOUyXPg2z0619MzVjswhx8OjzH6M+4
ovxUMcDBSKCgHvG0Tvn1x6Zb7aD6c0xeFiWxe7JvWlbvhRdC+rsdIAUwHPUUsjkY
ZpkCWPqftpN6aQFdQbgPwRVGyEnaGtAQatJtsPy9Jgdbg8YGDbwoESsnVcpUEbyj
FxbxTbZbdwJIW/THMpKHEsF/ixV4ECpnq4sj8x0KN/CQD8TysJg6xckoVxrDB5bi
6tAYMKDq93fxezaK5aMIRBgnVvnfDt7IDUBB/2egd9GMAHh1cB+gPe+YBedX0rAg
Hd4WPeaL9/Peycqi7/LVU9fn+Z4MoaAm+SB+I3LRTB0/fIRvDs4/4lWNEnjR992w
xUukuzDWdbgw66RBzsXPAO3/kDgNLMjyi2lW+9EZpTpvASLmRQsB3dauE52G58GB
Dq5aSxcLkULQW/SjHRIiBE4QsXRY6hGX7vWqJ3RAx/HvHyi9C+u2a42VKJwx7gz7
VtrySPd5Li75YchrfaAdZg==

`pragma protect end_protected
