// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
ImHZesJNMA5IsAhGCkVt/9/BlPTKuxlqwRUX/4V8Cgem7aCOkWy+moWz22WEnXwy
H+WXog62LSazkn5tLMOFNk4tEBliqFTPsEosLXczCJCbxsTV0O679iLCtaZGudB2
nuHOa+wQrQCE7B+5zb/orf+aRAtFg6jWFHcV1+xTAqs=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 1344 )
`pragma protect data_block
cm+1++bT0PMn3fy7+bUuDeJuzAHhN8N7BCZWQJuPVvlSgu/QqMhOiQDT3TMmWadm
ib9jkbKV5c/gxkWvxI+vJq/2idOEEFebTqdDG/PAE129ah6cRQgae199HTujTRQ7
TTOrFbxIUB0EFL52OqNIZGEuWwzK5Aju2euML4D7VKCcPDnotfe5F+rU0WBGZzyH
vM1anUJ4lt0GwVopH2V3ojhC40Tz37RV5rKaW8jjFluz3ZeOVfXhzTEhYWnPc0qB
Nek4rU2xR3/pFrpMMCPQYOd1oxinCqtvMoXqADJRjYN0YTf1sB7qRVkVwQaswj55
8tbe3WiYvnpY98pf6JRG3UGPMH4kW9PNpudOVusAyXZmon1h12+YzM5kDHPe2cd0
4CBZO3dGwO8rVkT5B6UC7ePuAhZzIgYZHDcc/aqUpW/Yr2Oj8kOljGKelqGSj2Jz
18GkEdf0XfZm0AAdUSaXuitMYylIzWw9YMKoeeeNLLq/TiQgkD7yY72nRkhp+FJl
Ch/sQt7LM3OXFlMOLBm/aQw5RKceY+hUikk2hkPOYleLGviFZ5EpDvxS0BLPg5rd
f1jjMJES7mB4ocCmP6geGiqB6ID7KqKTE1lMK7M+6JuXHQrXQE4DzQ7We8wDlUvr
Xj0pbM5MtVjLXVHSkw9IbVASwU14mOb5F0gupP70ACy9o4W3RzRaXhIwSVYyQU7J
SZn6Duo9bdTlxo262k8JwduTrCRnueMlSP1zdE2ghwpJ9mgGPWklihf/jOJSGfb/
b47Dnd4wVKqdj9mTwqw1Amd5epPv1rXfx1f4O81+vN9zyIZOdS2LpfcMmmoUJPat
/UCFuOC3f1bSBFKdwQqgcyvdkznjGpd0Qeo51C+HF8ULAm/yADb9ENmrOy3ZbDPu
RKdhHtwd1IWwliqB5WE1Ar77b+M1QTjYh2D7VMys5HE1XzPWZHbodXuCcn4x5kf3
xn26mOZcrRTIRcWVdzyp5vj0dNORSXCShY799GTrDbUco+KBhSn0owKjJUNjccVQ
rkXCJbFOyaHaxqj1274pYvz961NYHfxOkdcahwokMuenB9ojM4sRwsDChJq9H8n2
HB123UugcjGLRjmr01RFsZSfALsJCtnBty0lQNnmGmKjKK9BmkVKo/82TyFm+XlX
L5m0vHhQ8wZPfZaCFCUsROJTYyeMV4MusDYiLIXctqW1lj34JcCMITIfVpZvR2uj
SkMlYMJxowpspE08pkYu2oYvpYAIxvIBP2228XMIOFh6mei/kJyhtln7wnUwa7Sc
ok4kQV/P4oW97fkY6AJ8gSec6Q38Fb/ysx7GUse7+VNGj2Lb09A9BpaQoz3b/uQR
U+CZr0wF2OH+zMkir8MbKYHCeSfneoCBaQbNahF9akt6sOKRsc9nJuk6vD+uOKu2
hfSKt8XLCJrptIMCXYrJP4ZKR2VFZu5F8Ryp4mEa/klZ9BGxw+FzRcWK9z4vU9+Y
u5f9miUXWhTAYkxcgfp1w6cQYb473KcLX+HYtwPZAvJa2nWy4p+0qxG3fqrw3oLb
UH6OJ0qJO5yDpNSpRQ36e3qrtUEZTtt83zp2Y6TVd2nhaTWKuwqpuj7wlKeiIoiw
7I/cE8EC9R07Rskf9F/htMC0EMbtin2TaWL3QBDON5YndKe+n14fQA2ExngS2D6R
zI0ZT0jDgyGPBJdX5e3Wnk8AVJIjCCbH/eHFPpiVBPRtghcXENdX3O+SVbV5raek
IRICc2i0XOtxyP94aSjWbCICEZzfXHEhr6J634E09w1tJZJVoNa9eSDfwil5c8EV

`pragma protect end_protected
