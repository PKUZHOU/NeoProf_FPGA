// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
kEJmw5e5P+xl+kUWk1Chgb/TWxfNrkshxCLZ4DCy/ZY+ir2XhfRG1xex4kSCWL1pEUFCuTUIoRIc
U+TcyVaiL0Q9QO17GIkCmaZ4wytHyamv3mK2CwUqHZEW/gmY9t2SLXoYSb5yunU201LxF8sgEqiZ
hlg26CTOG4h234smartzkfQtjCPnCpTQi4ShqG8esKWc7C1Ay6lib/QmFvW58js4/Md926wue/Dq
QQwocxYkO5T3eK3y4mcToTgslrAw9YOAEQ7aAqyUD+E3EdZIeexri2lJyssJWbwl/lV2+t/Lh8m3
cMUAKXxNe2QcM0KpFr6xn79S+HGfh1GYN05csg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 8496)
/dIXQ5cKi11G0VA1LMxZXWC9YIHUL81CPViGjEthowEOZ2UVc/PduWXi/Rq6ccdPUTUi2KFCOB+m
9sRA/1sBwqjSU+kE/Tyua1uKEq+rZUCTOvrvGwx+V0NGu6HsrO0EuS94EC0e72h/vvf9evfhiRh5
j+uFVv9HLdP9TvZXjoOSPDHhwqKRK+jDPYcIGgNEm8flOoCbBIqI3OzVSqgwVgPCXzhmj5W/20wG
o6D2WnYXwhYoy6GSs4FoGxzxDYhl9aPU7FBckoMJ8cA5AEwPBYbH2dlnfrPhRiZJai4rL7OPTHgM
ZvlhnU0k9KJpBxjughLjeusCXkuT8eIo8F9qYxEvii3LXwgbKIfGc9ewEZUYxqf+wc55plqUL1u8
fUjqOL0LZEpRF9l0fNbL4pdU1l3WAOpUgqBIkT1vzB9DM3mvzV4D7Grv1tjHixk6qMmlFcGMVNk7
efo3TchYFnM3z8UIce8uEkokC6AWN6u2OD0Xstyphw0t3E+gfVHBd0VIwlqHkw+GxQGRBuUV/bVd
YUrZ2EAgLRPKYCE+oUFr2aId3csXPBZNaBdvJAeXtLheONCiUI2sG1VckTXr3N7DkhBc7uZ/+/Jm
iuz5d3XFg820zq5rSYeeSBP3+nOvTjaFCNc5E1ZlkvfkCbw/fQA32/K+4hdI9dxUoA7tK08YgQGj
cfDNUxuXEVngxy7ZCg7pt97PMYuVgOFEitwgwEpt878gj58sga3ov5JLnbym4nVVeibA+94JlVQP
7G2MS6IxOEvkAQlEAud2/NRPNdZ+FIMEoSy44yJ58jhf2Bc1oaQh/7ZyLAaug8OQqXN3RVcaMqVG
CqdpEh3DY08SAzZFjpsc0+PWFxbglYVygXCSgun7E4jIUbPuWW/yJCtNIntqmlnvquieELimOUkv
TmjFLaYoCRDwNkNRJT/jRKtN1HMFBw6afrlcTcoXQIKBpANPsmsLjHb3pH5gOMDHWB4ebNMF6WB1
k2XZ4bDTUYNxE1XzYJ/2LJ/j4c34O+0ecH5cI2L+bZKkYJDJb/bWrkNa1bGxLl5jl7yM65NrmQI+
XCpMYeza635W3Q+KKQH00P25I3r0gqg3iDESmiXhdzfNjDm+jsdDfViMPH1aXtHWpVfSFIdCDW68
vSpYYvh3iVSfpPsOcuoz/7O0ufM4pixWZzmR4tU/IWdWHvg2LTnkI6YJSbOjiHjc0E2DZeEsZx/1
JjPY6CqsLCBfIxRTxnrI82QUkYDJtOKumbMxnoHAr8RldduaqWo+yTl2s2+tRwZz176BySVqngfE
zGxhAK4IkyIyN8tC1B5inTu/GoKgpwJ5o3zhjU3orq0Ds8HLTR7pqavGBeMCgfaM1a07hHZQdpDt
qXxT0COOBj1viQBBNyVOstpN+J1UY9W//qV3jc5KFVS5qm5wSu7eCS5/ZMCMpJRZBchL9FEszja8
jD/NF71rLuRzr5iENmzSE8omKTmotBx0uDDONVQecdOPUU4aKSxvr53an+pOCtEjEL7mgRhv4Bh8
R0gb0Hsy3OYVqPLCkKI2oo4zl/BQEauq+05k8YoVGrPilJNP5myyVtST+hPU3laFt8/QIk2RVfmW
Nf9/3f8Ak2IIYV8USIY3A4H9Xl+4RUQ6Sm1oWPzMiOrF6r/GmxbB54f6SyV4vNF1uauxhdu8kWsS
aSfE/1OJwrMkwr77wLNtnzJm204FnBqDOzJg/Nn2tlIawSA7uLxO1rutYaUSLVGgPB5YPwHKpnH4
z6nInIxJx3Kg+vz+uTY6DUQuZAVOIV+7vNQtFhuVgqjKmlb2npBUDJpJxUwPYoAWvXN36H9CxzOs
niMXMOinis1d6pLvEfZmFugTbXaae2TZSZw2qFJUXQ4qPxOsAB7L0KCphGkjXE9gdyTER6mwzFYF
b147DGw9YSyYkhOsB1wsC1bm5sWTBLxcOUqR0fQ6BrNe5Ur6inUlBltREm7x3zJWxJm/7c8iW9nM
QKbqzviqA0fDP+Vl0q9n/24P9fhDp4W3waYrcVL3nXjRN6gA7G54Dr4t2ygn7wZzHbEyIE1CmfjU
nSB83MmN3NG5E1/HK3biC5LqBttRU/zp6KBe9ZxoxNqtzL6AEWbmHsr38386hnPQggEdSFpMXsEs
Jxa1MMSjThcJPEl3Hxx8aie78NOKCSdz6WgxliEU1srfCw+BwsQoNTFj6tfe52/0J8phkpI5Ze9t
9q6SyFkukmebRj1VkcyeFIegmP3YkWNLpie8mx5mxBDeGIpRKSm7/cMzPZ8BBRJv5Je0E3esDLRf
BfY28EF16tsn3E5XhOlPl690xpiu+FrRO0Arl/Ja1MPIwWK2p7COn5W89QFk+5njSET9y/4kRr/W
VxirS7v/NwUoUHcneZoB5bpaye0SNmDeWP+A2P1Cl5Yihx4sUCJAGYPrWxFkGvUZaQeSpBq+dtAY
MXrT/oPouLUQ8+pi0eyYDeOXxoihHnJjiD9UQZQY8G6o/9H4HIxvV4ezsJFB3CoI+nm2KcT6G2qQ
dQxnM3a+eNKepWqJ9+3z6VmD2EEtL3VLI8yubOkrRsmRaID7+q3WZtlbWdxnAdkL4M1sRTnJjH6d
xqhdy8vN8Mk7eIuCoNEFMpDCkSFaCcXP19qKYE0WxFxYq42OokC88ojgVEQWoqlUsZWy20E/+4Ka
hID5CS8wUbQvIEoVAt1xVH8w04Rnrirqg7/dOeEpuHYM7vr+ZuOvrUh0ikvngaKATLwpTlrriE/z
vs+jpVMQptjDs2qV75S/F4156PzhzqpRyWFwQ1f4s3YNiJJTJ13pSuhreV8pxiIRyS9QuVCo2Cl0
j9OlajeTkLJDz3qKzcAdI3Un7jTTa4Z+UmzJnSG8JSIJRxAMCPZH090s1JRPNe/9ML9nNQPChy/0
rITZkDs+s6+1taZ6ryTqZtATxYGzuq/197WwKOVnm6LXvY+sUkVJnDoHoSkiFLmXO3EtI916LjkL
/RGLnVg6rRIi6CCHuCevPdGUsCQYBHQNGy1iqyeJt/Flp7pIaVRUHqd5PWyux4g8n308W9PuVH4k
9iwtw0c6LTRjZOfUcWRSIX4HLPa1TuWLD/VHttms2SY0jdAOixIK2S94bm8Ow9Jw9An5HiEeEQhX
zTRJWqk6FQh4riUqUtCW0jCz29otMZhAQYnMPSVAeclhxsDg4fHXa+82sCKIkBqexhpPKlKaw2I1
ua/kr/6TTY/VHKbB3iJ8Gw5gO9GmMZiNSa0nBJG7rGZKDdMSyM99MvEkOv2zvClE92KsymFO8MGj
0cisU7D8ISFl9v8wH+lbaB20npGFysZ60P7lGhjMbxxyjfVY7E1NyUSbFrB5ywo9tndEwvwxqiJE
Xo7Rw2OmfS0jfdR6oug0uxqNH1PBRs0rD/bMgkNOD80NkjnR+Q+2DaGaoPk1zo2N/8E6RPykmH4o
RNK+IMH1lmCMxmWf4VcNyqpR1lgk7giHcP4CuurR1V8jjSutGm4P0hygfvjJVcjQmR4Pq9obU0hd
2ozpX8AvudlviD+YIa6dQ6GlKBM4lQjmoOUF20bBK6otIUlchODvOKxsFGh7QCSZoGdTiQC5MRM1
jg4SPj5gbh5nsrkxmMAURmqDo794brosMFsLPn4D30ak/Ohhw9eZrzOJDRYODnSJbTOPAmrxIIyD
vongTJWcKPMhOiMEpb0EfQTY0yVAW2NB2AY3bqwEkQkBD97nEwW3ZLgr+cb1IU9eIX7eT3u8kiQw
4IVd7/m95T6n68SemNDvQ5FW4M/k8/R2Bjah6CAPCluEw8VafbK9F2b9HQx4XhDPyFbm0n5dfU3L
+ANqqDLTDDPDLnmhO86CSYs4BJcfKA6o8aDmRAmYxGwKQatUBvNy49GQMyAnVIbRfQwjJ/VzDXwk
4k46m1xlZd4El4Uelj68HFCnVb2vq9ykxNSoFllN2Mc9w8uO7jqrE5/2rr4Y4wOxrbN/u3zdDvw8
oHvZa5edzKeeMG8/GcX/SGi3x+XVZAAQXosv0lP9KucbAp8hnDRZBTo0op2o3r155sb9P7/eyyD/
ZrWCv3PTFbdFuZ4fLKjQRnlN8LHmVzTbPbU0AwpVe+oI0U24uKVObTMbKxaEL6ti9k8MkRtnQmVN
UENRBBzt/G+DPZ1NanRlMHbyOpLXAN17XJv00MblZd/2W6pohgH3IEHS3xmi8PzakPRfocqtOX8t
TtZgqeeTvyinGz6QLLiV13uG3mBgiU6LKLlCFs8bnjpYQ+2V5tRVxcIv/owHPR3Zj5syNhPasy/y
gXGS/wedzvdgW0MW97RMd+FhLnCib/0FDP6kxBamoTWqfYg95IMj48Fw5jF3ZgSsapHlvfZjxp8D
W/xqC2bdDU5/KjBia+o9rQosGhwjFi4ROMsUQNfSUCkrRjrwPmHvg/gZiu43+8Ps8ZEhKOGuDXt+
G6PeE4TCUKEVoyYSp4ROeoweAPWz0OB41prp06/hKU2okU8MiViEeXUjQIa7TsqSaw5h8vPYJnmX
VAqzGMiifvapDJH2N0406r/Tt5VDezE9Kn4SoDzbzcGPoKtTBN4AlrU4Ys1Hce7f8ew49hcPw4IH
t2gWjSqKcubD1vMNCgYr4LlXP+Bu1Q66IQfNxk6pEUc9KbLRcp/NkjWSczHaXdY49KwbJK3R+kcQ
FP3mu8h5d6WFGVf5e/2tZKDddGzoEshxrjwubnbUtgUEAbVqW2dvX9ZqAifVuhKxXAMNW8dTOoCR
U4UVWiHZQoN7anyaiPx6TYBdyKG23TQTPBWKqW9ZKW7uD3MV3ZgmboK4QWSaUmUe+/JILGsR2GiH
dVzJdI1l3AtN48hQ0+XD/MY9QGOa7403tCCgZgTqkDkTz+rjMaARHvXUCejUjM/QRMBn4e32wWcf
XlcMRO002kzrDDg4rj5gHsQVAn6GEQNbbIIJNGZHsE3NHptigSmsP8fWIJHoS7N/vnUGrDZ3Mz9X
mWTvcHuLxs60PoIf6Wi5A78ini4qBQ/OgunNLi4pSnBVxws31HWQWrS1M22uNvSih1L60pQDxkta
Y/iGgF/fNhakWAfwpIoYYDzVYrv4IoAL50R+Z4a19bWhWfMrPvReUvxI6vNBkGsad8C2eXLzbKar
hynZC+BJ9zQU1+j0auzx9Ilaw4P+cPztfVT8IX/nb2pShktr6zn54bFWHHulCugX1N61v+m7w59d
hNZ6SHCkkUgMhmk5/JvBTU0RKEoAAOeezxgGUP4AvcsDoG503EnmM8oR21Ymlgj8W1DzD0wvIqZw
8yBbo92Y9XvJfGhiCCOqUQFHEdZEDnmagRvSeYY3KFla2bTcGmYwYRq/5/evS5kgRPYBcCAZhWS3
B0dCgd0VsxJT2Hc0CdX4LZf2uU7gUm0imxcbJHe0RYfvU3XOqayxGU92I0ZbEtLKaYaBxmNkMGvT
22RJYsdZUiuGyKZxxJR1dEX8ZK2+HoN2WkGDrQ2vAndRU/jjE2T1ei/5x83icowzEaJY5NnfT7KP
V8oKR+f5eXTRhz1un/wIA/W/xakljYNEqP2/o6d03wdR0C2F253UqFyWSRWc6OUzPKqKuOf1zzWj
SLoHTQjt70tcGnqL6IT1b2PKQQdsYZAWmYs3q7vV5gx2tFEAKGCdxdZNVzSERnZhO92IB2+YD3ya
6UHhZQBCjxJEc2lDnCIQxN72aKVPH57ZQYH7XN3WX1x3dnvjJlH0/bSyOjNkYvXE62sD5vYc8uQI
QBprqkLMnnxdjxf14o2mKK8GMsXrQOcmsgVfsDose1teRC7RbjcYtoGPnYIL+Dob7xcmR8WBpuma
Z0GzeQ44WiqZW7t+24/Rmz+tXBret4nkU5gwTq0EZ49wC6LJSM7XJE560TbJn9blH4wEBCDHj/KM
/jAl7gj8R+rcRxzygjnqIeDiSkXFrEEOAbvGpQ3K6ip7QFT5yBt+fMOqHJhrY4eWVKZPNb7aAt1V
CmKOtQkfh//fIis1vKDG5FmKQPkd7drhPfSqBtcYrC2nvBNoDs7vDBfo/adJ5GbZfDq2ww9NpUsX
nSY3uTQpUfip0fXGbJo9HUeEsqpcniaGVisdiwok4jZFeMi53XVQYEwLxitVGq8AyfQuQIZX1vMy
34Uw31ODqfMnNjNhywasjnNmRs/czZSV5IffTaazwBYjXnSlL6TGTJNjj0lj/8Id996UvAlpnRL0
yxSGup90edaWfpDsFareWs7iSAlmJjkF4zsD4GBNg7c9H3BbY1pxOEZsMeGgT7VT79Zr1vo4s4u/
iEEDcNqlQ9E0Hhk+K9nrWmsXm+e2SlcJyjygNohFtLpNjdh2152dhm36saWF5mxSxNoMhBCmdL5C
7prbzFObetfZbmtAj8cphw7MvzdPrNm6/YIRx5squ2MdcgGA1xkQaY6ohT3FUHce2hQbWKnDWxrd
n4zNoAFTSxWtBHXpJUpYSfSoKGc/p9FvaQaMaEHTO7s1iqWyIgb0SA6YEF0waBsbP3e+lRg1OIis
BDmy1f6IXpYhghgfvLcEc38JT5AjY1ljaX1+vssA+Xr+pGW16NNeA2fzPDSIxW5GLwjyIZ2D855x
uqVV4oWqWtWPYLfiCuizrfhp6Y3g3SiTp5MNnCppp2tP7v28JkPFbAt2gkdQUrF0q69L6tsmCeVs
U99gsMM9qGQfmKIEycjB68bdvB4bowGw4AaqDzqxpdPZWh1/5tmUqIX1qBN6YqrQruEQ/RUsaC2A
1DQNFJpBpkShbwnDdZfUePWde3OcXdk25//8P7MnqojQNEVDXyk6Gfg987CxWBK/nJT3b559mKO9
iFkotvTCTmznHp70nRaCH5qxc8Xxqdlv8acu+xG6p9Y0vNoMuMc+OvX4OcVldIH6esOyJFjv0ehF
+cYihIOEe6Mjd9Y5D3xjNpqTdu9KmiKsZRcl9Q+4zD7PqYW3pDYvGbmkZdidtGFyQxLqftJcRpdq
5Q3RcX+vxlM5+09zpfbWE+At//dvVB56+PXJRGWD8S30WQ3UNkP6nJoRXtuRFEH5Cb1yqXexx+zK
m0ljRPrv7Dv3qTxZ7zAgAh2mGtyv/wbq7rG5LxVBSwZPd+8ZNi6KRcMmZp+/wIKYcg+CHWZ3Jmgz
EjiU1eCHIZn66mmUZuCo8Fh9TjdeS8sKfEZtjp25pvs3DqpxNbEtcmjjO+QM011Aixv9ZIeL8iio
BiS0PB/+qNrp7RdPh0ILP8uYKaXtrzG4vm2y/ogcvfjXaqYErB536F0kz71Zhu+XAH3YU6uJVtLD
OiVnShfuDE5JWwe9jG+iW6wnUIx/Y/IQS2Ozhez0wn+9fPa+4iOWXfydYCYoFWHAFvB1h8WVpmdg
OT7w+78pNgoLC8oSCKjD/WxiUy0/5UQ571TgORDeW9Bx3RzzRfZGP9EmcxbuLRncGnWJohIJUOje
B83Q+AV6He8Dwukgfuqai4WgQZJher454UWUVXD6fu6NsAKkPFdz0JNMBGojOzrAUuesfyYTHSln
puNsyRjrHEjyz0iqaEZd0iGWDhkNnmjP+qKLw+I8DBj8+qTeBQ0Ds1Mh0MFCRiN6i1IThq26ErCz
3C3GZ5WlWmyMb1Q0LNW77e48Hwl9usLII/SaZvzlHXmZ43iz+tmxCPvjItF/1wRA3cdRKL+HvFZ4
6an9S/9NIp3KrZyN8lokvEv55We0wuw7FY9nAUtYHWLioDdMc+5HP5Z6LfVRjTSaJLln3wfqR+J8
7yb3YzzzFFYaEy/L7ecVa3w19MghTIwFHW5FQAnUqSBEmj4HJnGQwerdmDe57RoMhFrNxZ0hVbjQ
cinsEVsK4+DnP00ikoNjq6QJ9EcEAWTSWsvgfugW2aG01j2xnOMaKDxr8Mk49yBVr5fhJL1U65Gi
LTkh3vRfCs1LCNdthCiSnhSm8q/jzbyi1X4tA8fF/OcrpAvd2WBBKRS6ylBLjthLrQhY6m/zAUkK
XqOkOPP4xE9Sdhzv4k4qqzEZK/qhpvJwrwl7VtugY+QSdXncVj21SC/ZPgWj5SvHSJDrIJn1gp3x
gAHS7ladzJJcA4BfOjyE80NtcPDsQtbTYDYyOAfis7kwYyMl/X+3/GTg55hcnJ3EliCo0qtzSO18
2KdjCndqNSNc0yzA6PS5gQcXSXovOBPYFFk2EZDoI3Sn0ofNR/qujcsugHSELWkloJkQv/l8Hj0h
aKOA+9cbE5seCn5Y6r/mSsBamhj7CsnfDM5/abh+KJN2lXrr+3iJZty2ADjqCcjlKRazchY7StBk
ixIXf52qwSTUQisN1gff7N+9xmW2w2Upk8r5CGvdhcTdewDBkmSo+/0y+5nuoZ1/8ra3ZuFlVToJ
1zqjRN9EaGIrnipTQfHqFoQy/UOekkKPUe0WkN/fMxEx1oEeVrwyn0jjMDHAMJbTQ9iScEvPETXc
ZOK9A+JavK17U3LeSvhtg3Dln7yPbaOUzIaQs8x2Y3Tr1pQookupmVAnEpYhnrnx+7ecOqNr2Vf3
8sLUu3iSMCaqqNxa7DhGNYNCfrbL34MVx5iGrccpV3znj4LDvYA96LpfAAurzx0BhcqXJxsWoHJ5
SXoJi20PI0NsLw+DCsqSSSvfJ+uhERKp9weoimHtJxe2fo7ekoKUPOhLW8sUX0k6Pq68KgXGVx3l
fCE7zjjywfMOTVC1hT4sTzEp5qfaFNzM9sZO9uM0u+hM8ywer3rMbJIZWGtjh0mkoPGICuVrhAW7
8L/a4vOMOVpX5oUBT5DZeQMvEPg3ibjpQrVO1ApyajGHTkw8LocMg91A0rhT4W5WodVcwxbDzlvs
clAzazmImTcDOjbL4/rB1bW5NzmNncE7bKHrsvxgUXudNkkTyhGKcUngJUwnU9eF+SrA4mfk4Snb
KZE0htkg2rlbwIta8NEGUgaIxuma/FP2DGOfgL8bncTKixp6yfdGLiIppDqsD4rXQqoZF/iMOa9A
KpJGePVRSJlfpkb4puiygvMNiF3X9F6rRqp8LD+bw+PdDFO2g5p4/dspkz/iEfaH73hLwr7NemnL
ciSctlZ50cz6pLeaHXP6Z8HAeTGe0qE2hiF8liGZEAvySLfpGsYNxl55i/bJ2W1oyCWJtZZmK4Oi
x9SqRpu3TGwKthvtgKVY4or0QRjla2CF9XDhZLn5WU/vubNs5lrcR5MYYsQue+tmXEVdUdf17a5T
KF5ars0tRZ3qe6hJhX7K+il1OZ5LfXyYYtHEy0ua0GdSPo0qbCn7OcSpBsGoPZ/j/aNTa1BmrN/z
mR1opKueJKN9StBNLyjDx0II6/tp+bUCNpcsJ0oAz1JW0QymB+bWLvhwRn1OvBZS0amyjqC9EPuO
tuLhflGXWYv0Xz82/EXNk0i9u1rWVbX0uy/vpH7wxZRC11oOIPA0dDVe69cnn7pQovncaT5UMBZz
9rY2LbCVLERdaDCEiZ0Kj86rcXtWwF7/ch0dsQeAEJR1TB39CjF4oOzKHE4x3dvQez2+xPGcGwpb
Ta7eJp07E7UgqI/wnciAdXAFHFIRMXQz61e8SOdfiRZo7qo+GVqfFQy4/HODavlTaFgdZ0Gvvjuj
V4ulc2XL1yp72LRoDwyoMIejeXiRHNdKBBJfWlcSMt+KlRPeLgaSjVp3ijQL33F6Kg/LhcxwunBs
RTExmJ+jRgiyCXg91MtslsvghVy0GK6JJ0SajnuqS30yq3qhiflqVgp8vElyhkL8hO4VTZFSXlUc
2hbMpwBOwzLoLxzXlhq2EVNlHJXOp3W+m9QB0eJ1smIyP3q8E36/9mWT8rb/SvyW6KNkuXEX9X4z
zPtHg7M4maZaJOZIZ+HkDj4VwQRssQg3SERg2CtQYkqIwNE2Rgdi282HWhgdpHZqie4jZ9qBqFV4
7X/i5vvRyN3hIduRuZOOu9LM0WrExfiEIMyURAq5DaU97YErFkN/R8AsYHzbRmAC86QbcKYcQMGp
Bc578dip/CgMqKraqyaD61jrOrgBwrCZNJ3TLbxHyf8Trl35MIMTxC8hTic4ejyXvRRM5yttSaVL
6aC9n3npvjUhNj5gD47RGAjRP/sYNidhDxTqxstJP5vEJnLp3z06jKCKPEwtWALZ/3JR7vo/D9LI
0y23leGCpHUCx2CAbeN2p9mrUB+5gG03Fzw4bULTxffHeGbPg9eAO8s/eNwmzargE0sQcw9AirAB
ZrGBsH1/AgxWP4g3r412aYL7f8SsRocvWjabpGGrNdU4lK7aFRc4xxDo5UyhmpPFi8ugOYYIUWXg
haSWYNXRwiBPQOMM1SxGroI41XORrv93za05uGUHYM8bwuVzCMNC1mH8YT2b9PKid0kfMSGGbWcr
pkuphthlTaEp5zrMIEKv3AQB83GxRJHASBQvQtitBrkEU1BBTmZgdRI3ovaBbRwVgXf+uEBnTx6n
hytK0As72ltELHA4QbvMBnOV9QrY2aWkOUL0tuI628p1/tcp+JLI7V8JrV6D4Es7sA4loZM4/uuP
Wb6JzloJHxLFkA2fKHC9CUZdvbvKGM+V+vSzRTrH98XsyfSHKdirS9/j6IXSoHi6w4WwI3h/qyCJ
Ma+2awPM/0XSp8WnPmI0DujBWVrUE9JoN1Xr33qLfzWh6Z3Ke6yX9py21Bc+9NGERrPCQ412EGLW
aiLIaIeeqejVEQIEH2hG6MsRIA189KDLjsf7OrQf+GRl+d0JN84/ScT0Ma86GD/he3cR9ikPbwMI
+xpj2BaCNglelEsDD8USgEyf9cAQFyLi7w7kpvVchdcKWGoD1OPOtmIYptRF3jN2HFtE529RHEWX
87MXCvC1pAzxamygU9j1QIMK0XLgt300c7/Kb15DH+iDtO+40aP7zpmNDV8S9ExcKVxEnWvtl0gD
AYtAxg+zNupGjInuKBcMNbHOHdK4D+/vsvve4tcpe//pRwbzYZvry48KuvGjM3r4uySG0dakStby
uJdsSyGysE02NapxSoYmv/kPlnFRbDNNeY48T6a15+6nhLm7+uFRNtdlK8ghgCReD8CiDQr5L2B8
P22Q34r0UPv4NRmW63hRX+MvomruLEChhEhXIXE8xV9Zx3XaQdLkWGIgMvGrEVrshtv0hJ3SnJhN
SqQF35YzrFMLCtTHVtqz1iOYjAJwO0dtUGbaY5E2Szt9TTRPkRchui3jZuWwf9mIB7bdhE/c7Ji8
X3X5xtNfWJXBJGlTFp5NfDm9wUUpqzY8KNNDo2IIl9hBzRZzyZlSuggsP5DP5WUU7nPh0FgqyFmY
nW9kDeMIPNz+1u5FXa48v8TTh4Xoqn5b56qXO5tNHcwP28oMOA0IAeab6kMfeOIw3uFcy6dd0Llw
Lv4i7nC285OW1YPquM2qe4HcqkKzyvcK8+1wd3HIWaIJhmofcg4yqWX73NruWQHwEAcVg5Sw9mP2
IIEM
`pragma protect end_protected
