// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
dX9VFluWZ+Q55lIaDcLZ7RZGYBRnLY89V+ABzy3xs35pLMIF4lYo3nF+M1vFvE7U
hIDqi7xec/aqHjHWZrVcTtLobPtk0QqGgyTsI1iJfOaHtz0Yf+SlNTDne6TZjAiv
6hOiBn+plb9bGbuYFi9LOxV7ph5kbHHFNxsOUzN2gAQ=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 95872 )
`pragma protect data_block
6X2snaA+mjnoIsj9SOuB3rL+0o4ax+vQI7FJM+2tBvR4jReMkXqHzUQcKE0bJC3k
D6ffzhMVkHKQIZHvyD/1OLeO4wkG5P4ZKBtwiy0dQP27TfBvbuYKEs7n73qQtrH+
dJByCBCEz8E/2nQpKXCBinaOZGHWxT96rCn3AotyleUidrrQjAtoChHzvCJqJT9X
lqzHxgMWwC9KGlI4bSmReXBZhqjr1MpgdG1WcECTc9WH7DVIy5JkZux5C7N7bJta
6N1gFYYOEFUyIs2WTh1vDj9ugwW1vD6Qj3wZ8QceDzIS7Uvm5gtjaNTrtntxp1OT
PX3GckHqWVKojvYPCKD5lqMsvdpqAZfmtSc+CPJ+98cwm6oI2SvMOuBe1CW+6GRG
URWR22zBKzueYS1VomZal9TBOrH7PAH3qbrwzZq9TQldJQXZJM/4CYGxa59/boJK
3g22PRlvkHP33/DFdOJzvM1Cf+x9U4FOgdAPMdMSsxC1s1M0ZBsNMCcjFe+q8kN/
zED0IvNp0wYRpK5okL/mBn2+dZMDeHUakHwPWQaGyJ8LFjccxzMsSTz2hUCIMFTP
bfUyTTvrNjVD0vKLwKK26EFckM0DBSrTMQwteuZtDOkrGKanlkQmo3rIoMsWTxv7
8lpTAN+zHp5LF2mSehMHlE6Hb34tfcyABzwGa+oIgVxwVRCcnccZnKSSRyFy5hEx
hL360c6Glqo2m225WNN3h7zdHWuiDXQNgMUM/HgeDoNa74sRTYDV4q+5rtBLauu4
am7q1e/4WGJ7L4OG4pCCGarmqUEhY59keS1jQGiwyZRkXEDNWRA9vc5JVyQ8X0w2
ahwDlIoKJ1uEOZ4xbvN45zSav1OQAdMsX3cHBFIllcKm/8YFuub7m3Z6ySN1Fdly
KBwPy/j9F/IdvST/PZTIQPo59Ip9HZdLYkTod7jD00Vl3TgKjpasEBkwLYSr8Jmc
oRpHBVDOjy4lP4Cuxh3LqfQX/faTFFerTRFdsEjPEtCDevKT3RuC+aPjPzJwTtsI
DMFKPvCpCcMNlo74Oj3hyO9eCN2afrk4UbAbSlC4h3A/TUEBqk+FK47T7Jwa835r
XTBVUeMndv77TBK92n1WEOC2Sqe/fyGdqp+1UxXpRnOzQ4gAdmcr+dry17zzRWpi
QyiXlqwA4T7Mxc/+tpu/pXROAZs/5XhikPcUQHDu/G5OM0rcpnwdKc6G+zdvgEVE
GLCo0yQMvYg8pbX30DBXqXkatD76/foKtEw06h++3rCiPYKnKDM6zLluqqzWhlGb
tfS5VO+69TNfyHbRUjKJEAOiRKupwsMjK0OFa1gDZQhk9I1qyO9TMuXjJtMvMTV9
s9yhYpNRHZRLuLrqb+kcDb89i4+1Q0UdhjTYA+0n1IWxiTQbRM6OUJP9ez8xihlc
pS9Ky7DrljhEx8LOCPV2mh6+ogBGY8JRGCRgMnFto8IXVG+GH/llAwCRAyUB7kb1
gBEajlRx5jWVg5Ryhu5Hs8/ApVPetmVptu888JUWUJAxz3Q2BC9sJwSGW4ABxMM6
UjznQKAfs4K7cGMvbP4o7MPBRbZsFfUYXEEvz2b8BGMPLuOTwlUjhpTaPqukUW7J
ByZoY4CMFnyE2ANE1W+4NP5WtR7bEHOXrbz3hoqZrm4E6LE4AXfE6F6rIZqzzJjN
EVh0J2dR+++MvCG8vh3WfV1/Wq1Znr5Ome+1Og3ZwrXGfdi+uEOr9H4b9KmRKwRb
C7ZWVkOXe19/xYQkkJXdnPXBcRuBJR4WYTLiUIsCvDiotx4DCjwwMhydbHeLc+i4
ipuTbuLxyE/ALIvNCZRSYCKcAaBEqGmLB12RlZO+/X1zPDemnOGALIdccDnm2glx
eDHS3eYkuwlQpUUKMR7yeeouN3iIFWd07gRFu8PYlyU2eZ7SQMWIgx5ABpsjRBuT
ZeZXcjbwvg748ZikyQHsB8fK/GY1L3z5sWO8VfNKksNLUcUK7NfvEZscIYi2q1Xe
Jgebvu9PdIktpo1g4P3am4NGpWj4TpNQA/k7pjPL22WJP6a8/mYGiopyWT9ZcAy2
1fKSGr3MjqGD3XUYlnHlNHqNseoN4F9grgMWNHg+YvyPozBmzMwtQQngbHi/bjdm
VHAbbcXHhZUhCODgVb3mjvibbHHINU6FCkMKM67CPVUMyf55zy3bdMXvg5BwqzDb
Ne8h1dTApKO+wYZzINcUlYlRQwJnvmQH+VSv8z+BdKB11cU0SMFunzx1omtWUvxP
ntQXNWimyIuQwE0EPB7nbhvb+//thVZTZmrIN5JA2olUjt0h/qBvhFOc43rxKLJd
8MN/6fVkYzP8uGSCwi0qI6QvjYaQZwtwRi8QxssZt/8wuluwG8I4rrcvgos68xDv
jQAJo4sCvfl8qT7mVlIoXUzGGifjIgByrrxwN1cfzCsLD9hKMki39KhoPxuiG+KF
qD3/8FD6rMs5u+EP6M5ewAZKBO4pYhu4nRPMPFG9Gv/Qaq4TfoVgScmvFzJetG0b
7J4fgQ2AbvxKiMIE8q41rRXyxC7gRBVX9W41eq2zSAnwSPxjgfW4BJounxpkZ9kT
sJRBKDESx8Gdw522uRHQ1aczMW4Vt5Ebgg+M37Uwctg86EBgG5df0Ez6HfHrhuEj
xCzfdvRgQrmPD1l7rxCmNFsvbHQippR5ZkEc3XvucR+mtfAlYnqyjQszkc2d5Nm5
ks7dkT+9D1T8djEnYyv/vKCauo1ch5nhd4ANxvAdYet8DYhvlzOUHHMaDbfLUYF8
aqK2oOduPYk4ds/gVQUIncajw6XvRJFn3RqR46l3FXCBqV+RvoDL9xUEJDQOTSb4
9EHQeZF9iUy1D1n8lrubzpmW55STIyLt0epi6n+aKrxtZKeZ1UItPA0vhu47Soxg
xZ8eIPZE7ThqaLz0An3gV1kM7fJ0lGDiJcwOzsm2pljzUJ0inqn4dH33vxqB/GqM
Zpa1UvC46gtuWs3RIXpYc6dhSg1vR+Kzak+tsyCrAuQnycgHbPsMYUtqa/Oq0/xt
hnpqVTfpysG9eXcfdEtTlJdLdPx94eBm7CI0pN4DAHpKE11geOD9aldvq0fTpsjD
ElFUL+5E2oZ75gV17+dZoiYoOvUaffF8iN7eLtWBv6bSmar+Lk3BoH0fb0LTFMb3
rCU72Jwl7NUthrs83lAC2fFN16vw1qpSkSP/fAUp+1Dh7IhtfEAPkuH+6RJPW5yH
1DvM+XMwOLHoHaovh5tshOEhXOfkWqlbU74aSs50PubZBkSpdQgJljVBWa6vISBr
NcUhZpWryg/WirL/VrO8o6JrtOBav15x+iZIUx3eREZQs/EqJYl4PeZFG4XWJR7U
jtgaWXIfDddFACO24VKUfKtVH7vWZ5RseFsbO+Rfbcwuyjh881NBfsK+ObYK8UAX
rx8iAXZik6HHeuq2534Wp7OxVrlQM3wOO5iTpHGtk1wg7cBRNwGLOKLasMgnq4il
iP5ePjK2GsMcW5h6JKKGl6b85bd9+c00lMAVB4BLjOhR92S5IF6fkd+alqqKMwO9
Puvr/Sw8RNqJ+37NqcgpJH2p79RYBfF5K3iN0pn4Ah2OSuy38fmKU79voMcgvFke
BZ0+2fmHaUFswmi7ob0QfoSP/dUYJwVCL0h3MDGkMnCe9a09Tsem1HpAEP3RbnST
5G3sVAq1ODde+azTTW/q6GCnb510E1kEcMF5tpXdJVUnY3kWDVJmqjCV/i2NY0l8
MA68Iytkqxu4m2q+YmPzAMOIY9NE4/JRUDIYEVCgpe8uFk79Y9S2bWYgfCf8Toxl
qBBviSQn6SrjJlzWn5s1423dw2KoX1ifp8ABgP0hOWzO8RHbQIBHlRD7/b6Rnzhr
DVLYfhhxRlkvl8RBgIVe1ySo/f7mI1OBAXf3BsOcWZtHFDmsaq6btYMMrykhCsRn
8HwhYgWcOYYIOvu6hjoUIxO+AHG5Pt06Zird01PWyY6shim5rjzyfTwAs7DVm7yF
SVjPhPomRwu+rDtp76IhxDS+ir0bENj1nf4KReX4lAD3uy1yBVHR/oOvwP1gPFtR
DX5+KQgAYffBM5btGLFSV+118+m/GLom9kfCKBGm1XyVMvzxdiyAkjtXhypGSf8R
qMIMt8Obqp/GtMbOl6mkmybddA9rKoPKYGjKWSeBJoh99ChlC+yPCnBgbu2VGX1p
USNwY5bWMYnzSQe8Hcbq7HNX0OWpxeCHWcYuTZHA2IsfOH6Af9G6xcUAGZGrqaea
qZBdAa2H3sJed/b0/VH3QwPgaBgkW0CTvG+HBPenzirRDqosqTSaM/U6tRIJKwfp
cMA8ePlt5CfaZj42bKGDkQDcyO8sDTu6VFRsS5I+Duik9aJUqqa5JwppM/y8S5qm
67fvicBAHMgAF2/6r61286U6nmk2HKHhDp9V2mPkDCAOdpJtE9Pg0orx9+yZ4LeU
yEfJzaVYulqCl9DU5jVSPfuBcKu8Fu0CJ7ZQeaI1KgJBAfXxBkVcRFvDTem2pOz4
EQR+PQX29J67qB5tnExLzYDHcQmoXqyaU156XQm3377Rps/F8ybFRCJ2X+Mj7Io/
5QLjXMMO1TZV+KPGaJG+cXHWVwhqHIG7LL6MF5FQ1p/NSBDW5Ek6pnlIo1eyCD8F
VZ4Lm/Aw+tdPzOjNNyplKaw3CrQzYiZXRHM5/u54BnQSCpr1cBVX76WmZqk5wXB2
SXmRzDyJgk/35lO9T4wl/TcJLf4Hd5OlLbSbVbjtzYHOOJvH7Rqs9NEkIRsGIW5W
paEEH1GhbiKTRW/vY5E76VKBpFnt1ew93448sLYLBO3qMZIm94jwDAefzEIsNxzb
gKv9Ua6g4YppEi+gNO2vHg+WH2upF9zns27ISKMo7dvBxEcSr4qKEDwvOgm2ivjV
lYodZAod0p7bcCHxfKncxAmKn6yILQaDdLP/iVaVS8iz8M9nQXPcFkg74yXbx2Mr
Dvqc4Z8l5TCbFnnBrKcV+4PKNClVWfMorhf8eqzE1AuIqZZMxaq/t/Gc2BQiHkXf
82N1Xvqh2ewSQXwhZsk3Q22Vd37UCAiWaBME0vSd8h0LZCBkWODp0addmssBRzGK
A/9YMdBOsx3EXSiuybJG7n3/FL60GaaOJNCxDPKiI/tA6E24Tm2o4ZfHnuKLmS/+
XMKvTEsxasxu9ddsKJi6lcm5N3a2oENFqlLq1JI0BJSpLSIrZ78SQNc4f5Z4h5oS
QNU9ihCVAxcc6IVGqtDYo9stdDGFyc8DVpaL6/z4UaeeTtlJi7I6nJZcSzBVYPbf
+tjhwzPc2SUlphY+YdNgrhQPdy3Ngwj5NZA/rgFNGNweZBoUmfa2rMlsTBZs39Y6
c781GSXtugfU4M8RADtw7M4UVFkMKJgQR9EZjsQeyOdb2D+hMqCNCwwoxaTRSrO3
jRF3OhwY9HfCUslA2KAt1o2tXGQlGQYaTx0LK34JxF6VUj+y0LN+VJy5baT8U1Sh
GsmslPRe7l4Ah0pDMLORF7LQgtTYhefz/ddpZbQiXLNpXUCeP9iqGtkD2LbD5xgo
8uK/Xa4VyVK/MWRkgDhK0pQtFwLTs40uPBNOE6okGQXeZ4BJ2pSrrDxI0kz1VocX
iSd8t8KwBjzrK3DdnoVMx9eA45+lI/p3ZCL7aAQ2OtU4ishZNuVM5v2Zrw7TFiF0
BqlL2LO9/erfb8qYePAvmR55KORVpEAXk5IHgrAr/r3rdpsgMz7BOJ00rTIymure
0vD5IjMQwjiVOFBscUSCLRzr/PV0mPMzxFKE9wHqqBORMGPDRES+EHya6027JkFm
mzo4K+6XU+OBAikrL6l8Gjm0boJ0EV4C00ZbKrvs2vW8bNZjevmWLo6bwcVQf6bx
wrz+0FIWYRUZZX0gU2gpEoSMnT5GjlOeGOdOyyS4MM5D4HwqXhtJYI8G1M3I8VeI
ADPCcfkyv8DnQs+tQ94vzfwzwVcJ9pOLEVKjZRjiaxqXrw9G1ptXVagNZx1pTRbS
2URiSAh8h1BrfYBnrNMh5r9Km/D+QyEMF2yev7YyJcQmQT6gr/kMNCRXen3BdBwO
+67rWD5zQQyKRzMEkN6RTgpnSK/JvDUIjRdMo4d97KHjC+d6iWDwBDa0nQK6c4bs
deGFV8kcGm6dri4Lwo7Q0WDNy96ndr5ZXkUJ2Dr86lFa8kBPfE3F0mWcia6IcI5E
o9aADHWL9ysYh+YdTQ2C8gE6kH8ZWzVhJkDW/9+pBO9dL4TyEJSNOmkV2KSeY+jO
caLjNv1NXMFZW4fFENtWbqnTPFxTO9u+zeElNX46YxW+3sbj7Fsp8sKUxv+7ggsq
6pqOGFTfAzlMyuu+P5zxm7VSeYIDpzMP4SdDhnk3mj0K+WVwzfkun5jvNXoL/tk4
CRRFIYTHcflWMzV25IPuR4MKL3f9TEE8/625zHGvh4rxbg3uUiwUimAmxXYkE+s5
ZesfUr4mGeMRnipj3ajCJlQqpdNuynox9rLn+KVetgpqKQEwoRWuXbshmFtuqENH
6MXRWKmYPpv2xaPaxw/tPs6KZRnWtjXxtUZ2L4K84cVIM9dG4DHavV8wa2dgZfRl
1Fu2eXaa48AcshH93tAqIb+tS8MMIkEW8OfweZy/0XvbtQj/VthznnFweK3N1wOn
fSqdRyyOaphGr7/QKyA2MTzzC41C+oUAqRAtcvcTMINhRFYccy+OlGD4yl3E8EJU
OiHX1QqwON06esh8pyI9PNDdna4XOxNMRxIzO+ZBPUv18t9EKYULs5255y0PTziM
/VKDeYSvrtxjku8zoOFsyZkiqgW8hEdc7WXzMIQnIwCbse/hT8ixnbooIhyB1lnx
q7UgrY/z7VIUnox9NeS1SHhBXSCd9q5eFsioZJQqGWd9pMhcEszD6de5yHdNZ5z/
ZRm1F6lhkzqTbz4O/UJNN17OslYwqV6c1Nw7pgW9V1fCUWG4wrK793ACeP5rM1LP
N6Rr27Xf6orQsqtU9KCsRb/PFd+gzfHyBkQt9b/A4XTVHgnkzuTBhgeIauWG+5Iy
a7tUNa3wfxExZ9jWa832wWlf6Dq2jjlphNUepoZSRjAJYSYZ3u7vxyDnmoxGXCYg
2CyFWOlQxV8rL1rhd5Iw+Eu3Wiquk7V8PvKF4lRAMS7sZBfNylWH1bIzZX2LLj+y
PbtaTx13M7uHVFN2IyTPUT57gQ4s0ZaA+efuihfTawvPncVQlphTUdrowFw88kMZ
u+Ivh9usNPdxxGvP4Ao52Eka4Q8CysG8jO9RVoXu6LynXXRrt5f4DmcOm/RIhzYu
zNgemhvmPzDiP/lb4+leV0FzAH5+4vCOnZpuUGOA0Qvs6Ec9kAWYFEn7vHVD0WJH
+vpa+rz96edBSFQzyFB4LZsOyk5gw8na5kdsLBGn5uQxiN/4cmOHQy262yvYqOvi
5MFrti3CwavacTjzMNZO8hQlDmqdUiqo3e7nszHXOYK8AaWa91weUqt32wDkqsGX
J8J+bh1YCrhPmpTsdPRUkhFoJk6m1gjFpuWYVWKiTD5bcwZ3fOyGckbHPZX29G8W
5Lb/2EFKIB3IxCE4U8EySngc16JMLQF8dVW/ycbcZTdy7doU+pZRhoeyCX0nohL4
doYkX0DlUo8m3zahWjN6mSAUFmKeQPeZ5/+GIgJaspE/K5XMOAUfs3MZjCJGRitx
iJCZ5B+RAtatvZ5ghlwqpki39gDcGjstk7nxB1hg01NpJkZTXD5kf4SBIxvUVxtl
nInwXuRs8fuzDzigM+3OZSmPAiCurJwUaZ/NBWzavsSK1G4njh6BcGj/ZoP3H8LI
eOS9HVYH9SJxsk/WUnv3HFfhX5ntIFxixiPbJzIvNvw3WPuzRzI3aKLj4vUUS3BW
0rI8agffusmWv9cMrTDg9Jm+bNV4UI7AUu5oBlsR81J1pg4LOYxuhyvRPmoxSca8
6BB60T6ypRBdpjq3Xg03pPkmba5UNdihqjqmdUJ6CEzVHWSMCo/QS1On+1oiAFZm
Bn7desZYDzIoLsF48fBhbAThZXf/dHijcNp9brld1Qwb0KQF7llOokuqFOTe61HB
t9cSVMT6bhTgnx4FPbX/LpfbYWb+TiGmSLzC2adTSQu8QKLH0rfFckcX5T32JVp4
/EEtYvKXCE6B1OhfiESMZoB/fKxFikaiRorH4WCWjWv2l/XGcaMqVotS/tlcOLuL
yF7y3B9fe3oZTWnul+shgMpzVHyy+IwMzvwijsroTGKgb3CwYcDRzw2/VG9e3mJq
8nwHvL3vimT3BRhNdRs+HCE1uCXXtQL4yIdHVJ8WKB0iGJf/QqIuiG5ymEwUFe1n
/hT7r86JNFnP0UDkpLfT3OqVO528OKRTv+A5jbO0Ctkt7Ju9Rybk5v78/s++24xf
j8SAcAmp6kJyGbCsuXIDeoa5Ww1N99zLK4Y6A16yWO6mmQ0YmdGnB8IEEdfYbmlk
DMET+RztomGelPmCuIQkf2dFW0mSQD7kmR3cj/lt5TDCh69OawAj0xecv72/35jh
VjD+EAoUYRXvZyaz31rmOqDwrdaq9bgfqUI9cCuRp8D2LzEsAc3wigM/pHWI3jh9
xk9y5Aql+cz1doBeNUo1GPoKp3dnRQ/vMZgCa/jObhuA6MQz7nua1gU5xZaIQPS4
uUA5F0fMVCF3dZKGf6yew23wueA3XKj3eMSciRK5vHV6cBgQH1HbmBQc6zP1uPK/
6cPV7/sErZdbvMFuXQLbXBfnFbt9WiIc34rNiICkGHcBb4fk0Tq7k1MBdmCZU/VU
NYXofeVsFpPZ4rleudGGxm6WiJzuGmzJSxVhfBX4L7jClL01zTogA7hTCnYgg7Oz
mcYeJMJRppSWA5Sd1sgg5bEXHxc9MokJParpKxsF9sgbj7HOELdgrPikf/NBNGIY
9q9Hsb12tmqo0ECM61/RBfwNTk0QXckv/H/s02pLZ1NsM7h4BDDfivbP9LOSaMpS
REAmzgTpDsS7nNCSDmy0DSmn9S5IDgOGjEWwRM96RkfaHtaOE1OqHX5618eAqMlH
1kRhw1QdsHZp9HcavR9RKl1HEx76HRfBezfRPZ2NkOEdTbQ7vK5XiX/EFjPrGIZS
1phpdZ31cvnvB6omI1g0zCuveneAjy7+lJAwYzsyAmpTd8pEOxEwBjgqkMre/zTx
FuRl913xXWk33/tjeQgGmJeCs0h+EW63GGSlZ+OBULCvbiM7ukkkmNg0aOIn7sQM
i5pX7z4yA8AvsyT/dd3oBrEfSAgPH405ru58WRzhv6QYX+eqbNa8NrrRJaWfJbq0
jhFoaRgG/doWbXmtyMIlCGx6kKZAuHKqKlfp2UWgrE7t5m5blMD8B+r6fMKnrot7
UR8hxDm/DUHkxVi5L82mBtyNG7xALJXLdQ7ryfkfRsdepQrvLga+gFokGTgoXsXH
xlXzYxh1hRlDyp8Vrf3WS4zDMnAJL4luiYVvHhVc0B4uNV+9x//EoWUmQpWZz86i
SllaQkl0D6fUeJcFr9RnAirvUGKEscY4Kpk/izdADrAkAtd/ZZ77trFTWonRxHFr
+hMJ5x1Zr0lBFiZSIaGNiEWxYFD4zTW15CFxbOJ1wn7EiS3wRw46lINiUBuIGGtl
ulxD+Yr/ygmd57Rq2/uvIv6uuB94NqI3HAKkwA8DKmuF9WNBW1V8Opl19wc7Z4dG
u6wMSFnSI3WnibJuzokxqFb5LPn3qb3Y4V40k+ICFg+IugEzV3szjQTEBeK+qqcc
qdWSKsTbx7IXojMEF5Meu8mGmKSyWGi7j5MXGnttDX0SwhSiIAwMWu8eWqJoI89h
iwBCqfyWIiR//pCm+T+pLYOBRY24UtIN843tJ3udAIyUNgM2kFqOoYZI74Z+QC2y
Kc3kQlwhvVxTvB51u2Q2MuubhfXL8dpeBJxYQwM8fYkgU0ABGvDGMUC9oiwOIVvz
/oHt7nzg6sRnGSc+l3gT6lVnehB/SHlwHXBtHPjSMnNzlg8z5J58P8WS1PTB/12I
xejrm1r4zhdGDH9yNGn6SLjivm2QhBXVu9TRKeYn2FIfzl6+vCH+m+16pMn4GBOA
Zdg9TcdHNX6k3lysU+wR5qBkastarDrTGGWB76K1a5ENPYeiPZyWCkuM4gE/gCgA
2DhtLwP1IK9JCTXFEUl5vmUb5IYlyogonhV/BufhUMgAFt7kOwFee3ocf4bjqrKW
9LR9ZbI5r0IXryLT2B3sTJHdOSl2vYW2uGyX1bHY/gOHMt+D2eumcxqsrphJiMXZ
rUMossy78hSPS0ObZ34lUi/0FEqo2aINr+nEx3J5LNx4VlxaQzmB3aWht/2vyVMQ
ob6AQxEdS1oMP0TdDrVXSmExlq0M1cozBIIWKpTt3+eXErveXIaBS+n/SwBa/osf
6SvdhhdHkDasevuJWWwN4NPagKUcqpVID544iuloeEbUin/daPUb/GNgGGIj1JO7
m/0yAaCjIdCD7ZzX31gqD4VeExbFVRnp8F2609YWHqpGZpHVBcZCiPL0jVHgbyVf
3PrjMKrxklCPyGaihYWU+zQ3bE5DuaGSOBzJU5yy1PeHDq11XKiS+rJttuw+0E6u
RDsNucFh1Z4Bb6Creu2OFK4lnGQNCKEMyEriRVADXGcnF11Jo1azeQhMB4Uy5PI+
atHJsHyYSz1WN85knVx+hhf8ulTSmDsI7LP9giq0Zcw8cRB4gq4Tc1NQsB7GFfL2
/ZvCdPsjbrhiJXxKICJ6fmcsYv688v2tV/LI/bMjUcQ1+ZnFEwWRTGNUYjCu7ZVf
iGlcThNZW6LDEWEYHE4M1YVNfCGe3/0iy+5cVSBjgNdbYVcsv/OyL2Ybwctc8mXM
aznAN7JfwYNvim0qvOXXHe/JoT7fXQP85hkWpdkz771L9UgA+oAve/NOBslb1NJN
7ghy/N7Sad7CIkgu9UicbMnGNmcIgDM5gSP1+n2o4uEMEes4qSSLs0TvBUQUGFLm
BMNtSvpMWsfmJ+4GUvKfKf/jQGvfEPZjN92GfTnLErew1sD9W64YD2HUtlSjdbcR
lH42ktgt1Q8xjWqXc2d/mG3aFXJUa8VzySp2mL2lo8SNxlyPpuEmbK3BV7rH0ePa
Z7CpzHSwESHnuMXiuLpaq7bzQRNSO2xnF66uc7zhvTz4NQ6DdXOsVqmwvLXkayWp
anXWH+KndOlyF6Pu+6jvO+xK7PQpmMNcuSULFrt+arVZ7NL8eD4xinNs1YBZNmYL
+YDWUxG426EtkXbrGWThqqf9uQ+VBpwj90cNVDcKTpwsJeZjYNFKNlfFTspjLvR5
8IJnidZHVEysfDh/7yARISEJwaIwiwOFYvxpGqGFhfdVyuIbItxFkbfn3MrBjAj6
8XxvdvapsQTyJNgAvX+SFRr/yGIWE3N9Tyc67+VJO7GsKivVzzCY6I7PkQCtJWjq
XKOZkdTL+YL6R0kGGEYtRba/1rjxNhDVvlK/bfhFFGeid5MhVOlep+kktRDc4sTJ
kbw5CSPdF7Eiar7XaJvHOvmc03BH/ALUn3ZpluxlZahxVL4bCeN7YAN+IzbefqDF
diBlYHpIKI/BPqk9SdujJh/SDUVOzUbWosrOygRDzaUuleH0IXJ+cR0ri2L8sAPT
sYN49nePZElWSmkWfdBC1sEi6PIqcvliFckUOvnyLKe8bC+ZrMKoezetePi1cbMZ
QZq7Dm4UxyHz059WwUhniYnUq5Fb86Byw3ujKSMq/kVJX/lM6yA23+2879YVijHD
OdyP4ZfWQaBwvdMI8+w0yZGaJmW6I/eltXn22hP4kOdkLyrZwAB42F3Aktlhmq6p
03Q3ZsfHTptxKfWrPJ4G9uj9w8na/wvL4XPsBDjaBYQozY5cmoSvh3WpY+O0h2na
h442S1VaJQ3EfwEY6eCwfP0ICyplsAG5jCtF85gTUjuF+Ns+9FCZ0YvKqc0yIucM
a4YlcV4X0waCk8XQQ8uKmwhZe1Z2bGJJatfJCH96RAAEEbs35fy4JaCQlwd/IG3Z
4KZ1SiJMJDM30vvVosn58zV/QXqL4RrFIiTluK77mMrzdKKjAOV4caQ9XAAeZLR2
U9Ki+3R9I2Kmau6TNgin74SfcvxmbmB4Hq1+Ye9XdI44FUQcLQ/bZfofI2Dh1/RN
pYWmqzM462M5UOC+CznrR/Py7H1mC/Zf/YFP9Jo0SUDi5iv5eiTdW6ry4lMM7vfa
PqXJcjehLn6SF2QpSqanFIBdJfdJJ6NeDh/8nVrRGwWIJg4EBGPlCrJvADMFggJG
SPM5hLv0weI9bXXT3YozxpRdhy7QHasyIC4/PZrOoUB+ZZK+awVCj5WHdyhXjPoH
0M3KpPGuQqbwoRIEqfvzdtvAipx8eaDID2DaeEyzxk7v3pMbVUAmSFW0rKU+8xbq
wuJdi2DTalLFw3gSv1WPiTmeCm0ZPYS+GlMKgCGFSP/wOhQHiD+9jBn+PHzSHlsy
lLt7DIo3PR8YSsNiGxbtyy3p+rL9uTHkey7mzCZ818KlYaNFLxrqEsloYMc9vY34
YOKYqjKZ8OZSKNkdviyAYHi2PNkt3JzO1kY4m6WN+cq3L4kDCd9uqFPnMC7mCYs9
COicnVDsfEzKFeaCnmMGC8oG6cx5hiBOJT6482cxCJol6zQDxVD2xbiVspKsql7W
dvfWrH6phtbpYWO7n6SYiqr/Um66+FzO7ORFv4jOUS0J2wgYL9BWOROjynLuaq+I
GSA96atZdkiprVu7Lal9sgwDJYYL0TlARwxpGgjbyy2tnYMbNeGZXL0L3IhuBcYa
s7lgPUQPesEuQ89smHznl6Q8cRJDJZ3ImfrvPwFEVshBB34JZt5qfxL4edILz95z
H3QxeWVxVloLLDYGmyqn1Dkeblbx3LzJ8iVt4mGh7AkVkgk4G2pEEqrnWWDMf9WY
vM/5UWOEY/cgmGkYMEs2pC4flAWMg3jnKnSg42TWdUcyXH5aLu/8uH82ltI55Z5u
tCoCZkTkn2xmqoDQaoT/EnBOMxUqjJ3koT+UCBO4A6LP7/RyD8nhZ8v+LUgTmDzi
M8/fPBqCP9Qpb+WiTfqauW5einOhpsvb41c6mM4djsjpwaaXas7G+nKTLkc9N4ko
y0xFrtwAbcrJ79kvn4SZWokI9Z+DrRzoy7zhw2MvphKAelu9pt9bJ+nczWhWDt+i
l5ErR4Mv4FtEeLDKm5rxj79zFmISXORzv1Z0GM8r5nW1Q/vKqO2jwgdbogJYqs0l
mn1sIvkep34DfeDULWfm2BmCsc1tEd4cb/cu3EUBDOj6W5gluIa5+20o0PEem6Cd
lg9w6X3qVqOKckjjpsloFZECX0J/+w4tmeJS5TXYj6dwbkUqdyedQIgh+vgmQWNO
6mIUn2iK4kkr2kFW0OBHV1qIp7Twj7BhDIAA6kmkoxGazF372ADAoscXNMIz5aYV
vdm25HkHGWMjrqdvvz4ZS0Wlh678IHal4zYd1yBfVpGlI0/lRfcrYijBlaKA60vS
TjVzD44UA23ug4BxNPBQznBktihkOFSaf7rTH7BjN+9NuDx4aS/I+tww0G5WCjHV
j3jrzbkDlLp7LBlruo/hqaVEi5yNTSKMU9sVmvbAamgfrGTZDyWV/0pjszT0zHGl
Hdw9CxUTE8ZNl/AbYM1T8z01AmXUvuceOhkTzCDiosBgQybHjZMhHx5pYtqNKrPR
4gQSemIPB3J+8vqkdDUZ+hXfD+apO1s781JwYu1xZEUkCW7irvLrVEJ0S55W5YaY
5N+FTqc4xIio9wFzbaSA9SnuElq2LuyUskaJkn5a0LHCzw18lrSPV0sXcejXrR8H
EFaqZcoJptQEgQViAmTlIyK3ch/ooJ3OizYOFbteB8plooOqiLYfhaM6XLFwKynf
AsIhvhhw3q59bdYPFetM1oAPfh0nL5da516bbCQc2eStcOJ2E2fPG7N3ZS0SYbsy
i1T4k6asIK3oxRIE1fjCtwvLFDSWMr7cxrcU/dvbCcFvRsb81VV2BIt9/1JZvkpE
Uox1hUz1zilfjY768m4+8PwtoC+y221rcdAm0ErWL+EYpKgTBg8UsxRXsQ2Vy4CV
pFLRNLwtVhJlM2l4tzUpi5pFl/7QlUtHExZCouN3hoR07eNl2gzY7GqzUEQ1oQI2
EnmJ96v1cpOflvp53QDyDSbMez61q8ZMwVxHrmxfR4GcLi4XBph2SYuUApigjtB9
FOL1QZfBhN4OCreD0ua0jP/8uYRb+L7XL8PMBJoVDC2GsanjGw0N2vZuywHHZr0Z
jQvIbjYkqy4Fifkca1Qa7/plsqIbzeaDulXd3sLmw4CvymreHkf2YbKV1Dr7LxEi
D9vfSM5CEgMGCP98SkUf/c5LolmFJlU/Ioy5Lq5B1WKvZFf4l0LEChgRTcpU1WDH
omxdkZ7TP+EfbZLmlo7Hlh4QJ314u0gr0EJO70qwuc5UvhMk3uuBCP43/gZUhfk3
Wu6xICi45KFIh60+K6CwR1TsWQaNJfEQlDWA2bARZCIBX3RGrOSSYAcyE8jDf4VX
FznlsHi6eIwrRL6/IbcE0FPq0D71adu4pjc4V1ZsORZ83o/Go/csIwyuaFhlGYSS
vFageb4TEAmlO9Vvxfvgfg2u0/b80JXY0sMpjWwkWD4uuWdUz5kHfssn7nul8o1G
MPYRatfFMNGIDEI7Bu0GiI745EC0dV5MoMeQdljfpGwARMvDxpwDuMY/2q5H6Dc/
fuWLvblZRZGDcCoaxnnHFDSEX/Ge2N1p69UvJZ3TuCxvKBeufjEEnYKQDSK84OFS
ZhOSKV6kkGszJlT50Sp/0aWrahzL7WBAy8ujKLWLqz5D882gIeu3w1l0TV2PvxU6
8Mx1Fx7AkMxsJtapm+EswNmv6J1+RU7/Yp8n5AyU5RYA0l/wFKZAJWPDXqfRSOdV
/nZSsuIdyxRGObcoRfRGHADt7sbZtX8a23NCXL15mgEyTU2xZQlSYyVYyrYOU+yk
4TcRd7lx30wSkJADQHjnQsW/G4bjCk8DV+PBtuZvODA0soGif3o+uZjGdMxx/09p
tfctmBx8PvbRICsa11ZUKjnKWDHw+U9FSF8qLWlIDF+zepM/cJUdwvmtGxN1aeDT
Jlb41h0CdBNMUKeZJVGsXbdIBnYWMzwHkIN0sP8nu19JU2MxhH0LmMGESTn9wS+S
eH01UsrlofXjP3Chnc1fUJc/Z21CnEiUk63d60aCvQqaZ3znvxSaJegi+eL41Xk2
lzGFm7XdSWy78FTAM+Ztv2i+HnxhwkZmnsYvdj9kVyD3bxcK9afSr1kxNBFYPO+1
ExNYj6ftCfSnCNsqmbXgLZFsoHVHg9ok3RynKuG7rZxc4n3WUYaE1AIPX9yX8HPg
GkPviNCgPl9omLIJ+wA8uN3229e1RSWgRj2Z9ldH2H6scQAgEjsloYR2iuziDP2K
oqm7ZoWkK/924xIN3EFeEqiHfacrZb5lJAauqKOC3v3BCZJ7d0+6ImKc7M7IPAD2
KIiusqLbQAlNQYW4W41wafylV9OSFg/j1+ubrw1Kq16pBuBiyb2D++hP5dTBqOmY
osqvW1UDDQCuhomxdIvY4Bco6T1ZeK2AvUyhnjY6O/9G30e4zLqHBWfU9u/l9JuR
IUO3wpiRYaLRivdDQnNmLZ90FxH/QRRNlrb4PUm8S+lHo5GaySsUlP+RJk+ibNOO
WqaAn0sjg3ugFJ8YmKw76qzg3UrRI/PGEohT4H4t2Rx6Dv+1BvfNfVAqbsqRq5MD
6jYDDkjtREc/ZvMauPxgs3IzTdqd9hv/FCwyDlJBKJUhTLNae0nW3M2mjp8LByc4
ymiD/FWCUFCzKN2cAwfUimnEw909lc7FX5LCs0WK4E2K9adSTfthivlSiFGRS0S2
Mj5w4GzzvclNl/7/yNXPCsMUnsg8SCeX+sCSsT7x+psPlD0x1xPLoKw+LOU1X7Fl
2vXrgHdb3FOmR9YnY7m0MuVtGc4S9S/OpiWqflklCZSAwq5auYszpyU1BIhXMw7I
QSocwFgDLCW592uI3uhyiixG5nmcBIzIB1MZSnTRYly1OsgXJE0qIdKVHcDTmhsk
4UsITPqWQJKczccNOvUkBHgM1Sh69gKwBERkx9ckmX7jEXdOw0VD7wQMvzo5vv0J
IqzyDAilOWuKwXBuSoCbWLGkUIwFh70bPeRWOmfOq+uTOYyemYwQmH3A9WXWbOKa
LmnPqgDedmtcFXj8B2nmD+GJlf79ipPIdGNQ+9OZmCuySRhGQsjbnFXnfDjWgL0R
1PWopMMXNUXDAdm7hKe7OTba9qYVaLWRclR+TzOYkyoGqQkK7tzeTM/HfvQhkJKQ
nmHdWQdBl/3H1lNBvoXz53VfK+1ra7f6Y/FqsD7S2NobJTZbbjRMlcwkzdOswZz3
Lyas04kmxLx1KZVopBwDGDqqzhkEX+YREDdUYfFoVr18z/AjsBQLWg35GTuVZzGt
NMmt5OClrQWrn9WT+tY23+b2DhQKzUP/goxaeJ0TfIq0s1369Hg9rsrwpSi4T4yY
xQTrLQK8+q/Unzxop7vxD+LSfpBy8Fy3uGsLKG1ItLkqhT4LQ99IGzS93xVKfoQ7
F9lUCTkbXXUt0S7aZ4RrdGoUn5jZ2qFJOiQxemkNdC5GU0Uxn5zNbUCZ3dgcVcrA
cQpYm14vrH9Nbz8l0DmC3x+GO6jS8ypcIsatWFCBU0yS/og2zO+YBvZ+kM1UI+Uz
v9P37cocIjWsZsVwXqwgPpALOj+D1bZvc2fXmVkTg66khEitwmIG+hJ0jCswc9na
50R5rsF1nbDadAXgRGHl8X4ML5G0F3Ev+HcZ3D+r5HItj8vG3Fh2vfJ6dn7tJXAJ
TSnrsgzG+G882mwuiyFu96Xa4KsF0WQ/1PEjNgWP7wapyZgrpd1ty0Q6Uxq3tUy7
CHQRaFRbhXYOJGx6nT0gfdYu0pdCKYLpfwnpSZfh1o6NkATeIH90oHqdvDBT/3/X
2atmGX9FcGT5IZHjjcQhxBTTEzz/00Cxs18RDI7iIWeUhKqa0+S1xvH+LwOnHAqd
vYErDIlrSc7BxJGYurGA5iGXvBHgCPZLM0+QVRWrVzRGk4vrndnOy7EO+bBAwI32
IlwZAPMWBSSj7jbgbeJxo+NgBfz7ToHJB3sSKRqq03RVTh5Cy1/se3UcPs2tgWgp
xAm713lSfHk+HLetWXe8+1tpI1w0xuV96juFol6LfwFEa9mKEepCzIc8gvWUDK02
YT9mg5VkftJF+nZEhEZGr996bmykGMLwkinpQeFWLYA10r+nwfziuwax7a4rZF/t
5oi7ebiuhYKQChby/SH9WbwN5I/wKQIO7mCMMWrbw2zKDqwkyMGoUWGPSWEp+gVy
H4TZqtXNCJ+6D/83WbxsUia3oRxveEaaIxLA8ILUiKV6vFqFKOazTIJnJ6UmNS9G
S5Sn9nwAQ09zenH7w6MPJuFCAV2Mp9bTDtio85tgGTOcldPoFap4TGPwla0hgpjJ
0Btv5pclCoirVvU1i+Q01ZPZn7Nm6PfYi6sne3uSplSby6w48SbsbQSpQQ5Zgf8G
8BhWcK6IUzQfc9FpjUMftwblASB4VUaGMPyZHh8ZVLfOvw3Y5DsU954x+KBHtGpq
dNghyAtokXoLHsTsEz9sHTh8QGhGm45CNq3HZTW6MYF+U4a1+WlHxQV7801vSfSZ
9x14Fd4Sr/1hiG3qtlvn3VES2NsTPBjJLQ54c0XMMrWA3nsYSpuN748s8s5f1HO8
GB6dOoyfwLIhxivuinarBesELJCwh/mYTz6V+PY37fS/Rq0s1AkW78i8mPKj/igc
RbXOkOj1cUUKSQXKKvCGae+qw3n0IPzKbKzTSN6IFi/sSgEDyPj5vkDVzZJa9A43
Oyl0OtjNG58EO0aJJLZJ3JjllqPmcwHd3mBxUc/OxPHSZ1urbxAGLs/gl1ksY/+C
Qzv8lgk1f66g3iQV3SzZqtoGENqAa+Bin5MowM8/M5vX1zILE7CSN9Bm1ugdSJJz
6SviDIMPt48t/Frwvxm1Ckzp0RaboeW0lNQjVOQ5E1wO6CmMY5xYfBUoaWQ6HgGe
87w7qZD7GW86xjKQzfMsbV84Zm02gEZzdOjn//CYNwPblsPf5YF8hIg6qV59KuXR
lnXKtNFitO+BBNktlX0eH11uTObOThx0NtAwt2Xoh1Zrqq7BCoUZmDeGEEhDz4bl
qO39upFPdf+f8TyfH2ufg7RKHe3fSX+m0HD47Dl5eB72r6nvuq5FdkHwPuWusNJN
ILOPNSbO2aS0Tf0tQNHLtSfD70mwnTQ2drNh01j2fcvrX/1dqxdFlglALmQkpTaf
fHZoaFL/pkbqPGFnok0soNU5Lj4qre0fuzGuHBSIT9ckgqvBOoLAuQ52Sr5wa6H9
rz7fDXdPQO9B8UepOo24t3HvZXGl2E6uM8PBmxkvhW3DudEE6oDem/7dMvPZMA5z
YwWFjHciEZ2avwm922Kd6fMhKqITWNho2mmbx5avqxb+sqrDu9jr0YFzubUkSxtw
ZyRHJyKLweLTGWUqzqZ7fJfIGYi4TDyMN1I2kvjbqRKmw1nVha1IzEzPkX+lN9dQ
clfbR89zN1QyRtAhojHjzTQbKJgkCrdVDGZZN3bffM0YOjkJptPDoutG2rAXm2/v
TEm0E5e1J260APjgM/FB9OLZ2iqWFO7J+DIa6sdOh8O0vQfsMKO9xq4ohUVYAc5R
2uOmbb3+H9qRN+jbDCbvhHj/eA1neM/kszi+QmUUB3de49UjrBAsDFMC910gjb2x
JipyTByhKmEgI4MOwIZfCOXA1sIdnIX5lWvV5gbF4KGPMnOsd1TRtcqs+cfCHcQs
M0/SLp+z3qyfcrmfhw4hKP5YZAHCZmByuNfo4HFHUZBxO7B5Cc64c03NGAAfzWXs
HVdFAit+sMmTIM+UhSsFraV1Huf9epiUGKYMvvBKWsgOEoehLyaWRQQvoblQye4O
aHh8nyxmQa+vD9NbfyHQHP4EhZVLpcGk9vnpkw2lScLBO2qOisd3FCVICbqZ69Gw
NOx0jvGL9jFZR6n2F3KnJ9lwQ35c2vAdtYhU7aF95aal/sW2DvmVDQQ0vB24in1T
P1Bwrtf9Cs7IpBWWwqwLyzoAVpOVqZDU7LyDUDhLJOBCLiUJM60KB069dNr2i/Ka
KFkGX9cXUDrD8Y4jeg27mzcvDNdkYJz6nhbTI3Qc3A5NuGFR0UIBlBSI4KP+ITfi
MxR0L0rcIAP1hLe2kJFnvacK1RaJuzyz5kdl/YQmm7ZBH3C0H9iLtDaK1PdsXmvZ
5ze/8pKKS5B2wkee679w+j7Wq1X2EoLKKbJXiubJjhC0EfImBOR4Q7UWzPawOW28
9P7E/T6U/s7w5HrFgloL5rX7Qk2ARvo7/ww7QE7Sy4oj2n/MS9/gXQ9OFy/ckZLb
RJVgp4CsHDemUC7gn9lkBB3qLRVKB8JByFcE/kBsdjTHPhB+4N7T6kEM77FKEBwf
EBI4Ue2sVfB8mfYLOsjE5vjaj3Lms80JsSOOBub65a2xJEcZyqBeAVYOuxHWOJs1
pPXUzvKHzFRuoLOCZqRxxbX0VvyiqAmXMxKBlSrOoTg8WBgOwveYLH1ZGG/oMv7/
uoBQCnNde2szQmSQtbYmYCrZEzo2U3asJtCQ+1duORdVRJBq7yM39Z7rLhQpAqcO
7yppN+4Z+M9ntkE661bNIlf9/4guaXtx9mREk3Ch+RvyCGXp4fM4c+ESURmNYZlp
qJKT9onfayOe9jY8GfW0gkathZ1Qf7ykKna7zjnFtZiMaMGmG61o+IDRsIpsJxFF
31JlDWcyQ90/v2KPJ+M49TDImJYCVZ4OQySYilj7C+gi5fXzshTUmiubnG/TeZJr
KwQjHfeOn4gPnNnKYiHHZGqmzZ6M6wcY9zj8U96qRbEMwc/Ne130iQRYKAgi46zo
daCNFq+eRR1HTnxtrrDJHGqQ6oqrax7SeqtoNpWzPsK3dCcylEWLMga52qU0xVv1
bLxJMgNsTkCIjbiFT56Kp4KuyCbckDrNq60wtH5RU7IofPWOvZugxDCO3oW/I6P0
H2GIaYrI743nmgXC6VwrpTIduIaGreF61dYfAVTmgH/BOmttXfboEAwXbFyciasF
rnhTx8SNqmF6xI+SqMOoPM9ekeKnQ1ZuKCghLlL9weY7/Pp0kdEqOLMg9I7jJGJk
bi6rT/j0lu2mZdjYvnEdcJJHwCSoS+mFGHwStgP5epfpv7AXVncfYwmkneBZDDV4
X+oBhorHCRPGbf6Ea88/HznQVCFQE+PhaSCuG4l1ouykQb8VF26Vn/5KKWGxlxuX
ro4oEkvfeXoY2mbWzWIYhttUdLRzz8JdDdpKhBa2rnsStgL0UV4Fo54unjsfjIaX
MlLnV4J8E71DTevilBjBcSbDaDvLl4F7MmLie7ovRvpeecjAeehG1O3+05cgrp/Z
GonybCUduxxDmXKha2Sopf7yQZCxfGCwKis8N8LKhKd8JHzutz5jHFgFHpMEsYQP
mQkesnfq7RsDM7gI9FSnDDlzTptItJViptt7zPx8HFnFx7ltsD32sJC8rhKMx7TY
hTBtePoNu8qdrTq+6KHIq+wlLY0Hxvuc5fqZ7rA/k6FQx5+n+JkgLKqofrBZ24pF
Z1qaR/Q7DqTplD79AqwFZ0+OMo+Zb3diZXGdRtem/Uz05J+RHMm3NpSRYfJyoTbP
pKYNmzgFs7OzMXFwsd9dQWughREoPj9xOUhKGOKDjKkUDO1/M4/PY9bxyJA0TSyQ
TkhogoXMdWwQ1EGiEzXao/yc1COYC0tAlAsAsfnrwsDrSbJTZbcVyun8z2EavolL
4RbVTPflOi83C+X861Q4HIEjfQlyVG0bJ1QhEdgTuhhKF0mon2UqHB1M4SmdUaZU
5E+HJmzyXZlNePQJwbvM+QLcdLPA9NDl9IHmriZtkOU2fZegJb+s7FNzWhlN50FE
V61t7DOt2mU2RF4F1IGrhI/d1ClM/jwXOhynLlBFLbv0jUdK9nesjFXofwOyR6MD
yeL9LGX2pe0Qu06iwXsejkwbf6fb/F7UAfjCDlS1Hw/OXTfhALY4bV37u+2L+/Or
uyGUfj83EtfAqSQx1LWu7qty5n7zDpf6+v9GvEjWzn+2CmzyP69Yu+5PP4mTBPbE
E2uh9Rm5ATW3W+0uVfNZXjmzmbB1QrR11JcFHvqHNa6vvKWWMT7S89FeDIA6jJJu
XhGOI0IthkMjom2iYWC+zDUejU+vveI2/77UCYip0YOCTXx51HK7tumyvwZ/ApuY
UOiOpMwmaK4SX2JIJGEPFMUeUjHxPvRtn3bM16Cdqx2RJa1smxBkU/IUpmmex5U5
Ys85fkGOVzsxcJU0py+al1fNGvbwkGZKHrmJHd9UvIV1UuMShlo6XwoT4SydIkcl
CwbgrB7t23GzX3cU5HVNJ7NF4RHpMJHY7HUfndvHK67mUW2HzcgEZUhSNR6nIgUi
r3JWEYMzEDb5cEs2oRQwa2gIt+A/EIVTF5zWJSnLt93+mxkbtIP2QoqGS9Kggb94
6XrIuS4rYP62O7u7YIFCs6xq5MtdegzzTtiPEOv5sjCaZZeiayXOR40GKu6mNcW3
Smc594eN5VewRfcdAXDgbGd9loOf/4UhQuaGyym9nGEFDOE7nBTs97WxXkc/FTg9
P8T1UiR1TH4C5R4eFvUZ2wJbMcLs6BiePMfoc8/+9Yb4+ExFrphMxGjPC6hkWF9E
utDH5t5/VET2lfau7e1+lfCOknEt96JhQdxmgCFl0xnonDqScByk8OXWqnnZj3wh
7I/2E/Z7yA911aOM0kxTZULqdkcmdTVcS5ZDwhoja+CZTU6xJwdwde1WOhivfW2Q
BUoBe5+2M+9UnJ4oiPp2ebrIFf1bJ//KBs19d92n8yVdoaiL4oKOzwzMeTvLalln
0jAHKK8ExwfdPUSUfoVHvSY31kU4F5vUHFapoc2OZGBid7R/1FPeXHE61oTKSsaD
YPMcxJvgWK5vR8kAHMNvuQOAON2Dt4wTYg8dwtfzzA8ORurtupDhYF+7g6Oz6lXl
j5i7zQwT188iXE6+6YU5KtAQOxQqnY+SlAfSFj+uPQzShz6y1wKrlqObX7AzCLZV
VWoJXguUlZxPkAmAGoyTBVAcdztkpr7uGs8J8t8x1ul3WsLPjjeYKCAwQZPIFQ1i
TufISe9wFDP76TVhv0OUGj+ZANDkjq2weOaC6RafHR2zVfAkSMq3csLFmk7f4wof
y/EhYAXFtXyUcltekoIlxLuWYPkDa0rLBaDJn0OR56NsvVt5ZWFjQH99gseVjvJ9
/lgn8A8MWlTCu/+LpkKKXLaFfMGe07jXwFW5vr2axvJ4ZU11gTOY55wLuZ8duoN5
f+tCl7EFatNB2rmRYPqXqZtLattOOOfuYfA6SS24MSVqKQAJMQ14RA5C1eQbkpYn
9yB0X48RKgcZyY/0T8pPp5+XOX1PUdqkJ1dYi6Lcn76rHCAZuYRLBXMg0Mw/nbyD
IEUKk+o3eltl95NGPcLpJVJjDM9WzufEchkPzq/ObFUYHMb/+k+RmritHFkL5Kp4
6E3l+vc7DvwP3oLa9rNvC9ZJdG1B1BpAO5LVOz/nWEztskcVZ+d0Gxr0CJ+AHxp6
DOQyQcwQaDPUofhx7b43RTCxZAq3P5FORdKJiVZMItmOlRQcx0c0KSc9SI1C+wAg
Ei5ad5eS6orFSNNIyCYPd44VBu+/aSRzKOc2m+UytBqeb+YFCTdbObjmiwCPxnMs
47ULkSqmQYPc9UigaJ9W/rbSpxJSrDgyWe3YwqVX+ZUYeKOGJIqX1Px2yt9FgvAc
eZzbN5vJelI4qV4pw11TfnvIvGQLKA4Br48ULU3/C/hbXVmsh8a0KqCsHxB//EKF
Pfx9x2hENIhekdFcd9i/Rx7OehWdqzVSay1eRvViRa36nklVhRx8gaL1TiqarlHL
fxscrNUee69K2lrrJiW0HD0zthMNfTLpalKcxjClLJtQKKqHYm1MNiG9JIsoTP/d
FG/SxARHMU2998p0pjplUHECyDFfddIpCeTywMPMVJymKHVWsQHZgLubk2wHuB4l
1c4SxPTjNvwxXDihj0dKVqD2Mc0opEYuzshtmyoUbkT4jMZjYl63ggGn95t+/CxV
YZacHAwb0OepDQQJgjWsBp7qY849IfwM5CMey66BMi1gEpnGx+BgTc88vD68FRyP
3lberiUmkp+13AEVEz9YuacKobkBbOmjIwEi0829NJZo9K7Q/9Ln2fOeCrwI9gZp
GbuI05L2r/pcMqF7qV6wMo+J6YMYgAO7QFg1O4626iCmrD8NyKUvqWd0nMrW6XUO
gkmI8xALE2Tc6GKRzn3dee7fo8lLXjgVC3XHX3a0akd3NIoUQw1273RaO8IXb8Am
h4vxRyNdjItAoe9QmB+Pxgis+9ifmWNDHLcW7mFmJjkOHDOoCVzK9xAXKlc0OeVi
I0w69k1SntDydUuzK5bPpoU/gRCYzcX86gNyjFF1HhZYQyqvYqbRbwpVyGYadF31
l9QwhcEnIJ/6NUey1gLcFfPiPhoPKlhXe2KZumBH/fEt49Sv0IQ9xY2Kc9+cfjwe
n14h5QgHGjIjOpF3qD7mz56Sf0GNWU03IbH83zvHxihGzutOIxV+G8n6v1l3VbW+
W3LYp+Xii3FoGU7Tu0WQ+mImDPU+dFOALw02hYnEt5sq5dj2DpOfHcG6GxnaOgAt
Wu0V58sdZFDXiQNin2eUfniZbhuPDeUg1ogL8oB2Sq3KQoVNpTXDbsUrKdBeK66L
98MFwJKRNZYJOdVYCLJ0EnbXfspd4z2r7GAsqN2BYdCZvQoyroEieNQJwzi43Ani
epV4DsoyNxgcxCFoh+FXP2b616cgZHrAf4155uW5NCg1TeBdY9Y9Rm0UribvnQpB
knSoM2V/zn/M3ecc4KdcGQP9NfHcV2BaPO/NAUxxojhmOlKZOiA9DzATDVVzdmt4
YwL6y19Mp/4p4m/osV0/hExxyQjVKhQFmIhZIfZFmUCACS9dqn23c/um9G+3jH4C
XqUDasRwU33+cvDEUcnOZxzHVdD/BGzEtHFcelt9Pza64l+R1mcOgnNkzwwfuFO1
7HlVjUzzyzJoWdoqwqt3FW+5ruoO5PiQJBHLP7yvLFxUO+JlJy2x6AWDW/C9GGY/
ri5sgbsanTJ30gLiBGh0nTn3Im8ilfTw1hGe7QYh1Ajn2x4yygzu2G1nANA4N5bo
xsWbo4S21WpQw8CG1RkJgCD0E040WVlcUzCsA8qnan4nxUD9AyC0cCLc36vnk31f
RlIZjw0FImo5VqXH6QmRfL0sQpeyR6hz8JopW3sv1rWCSAxzusrk55c0egLcrb8r
jf+0tmHnxvfP3nl8Sb6qszDBKjoZqdV7LiVk/CenUjtmhHp8b4Wslbo5CPxwA+w8
JWNqWNEl9t64MWKiRKJoGV3SV/jsXJKcmp1vQvcxRm5UVVTRaZovYtfbog2XZoPb
Rho1Cpb+zA/ayoHytTr6jaTHkNPllFZhb4aw4ZsuJzzFsiyM6sNlKu7/8X9/29EN
8Ze3Ovpvmk3E5N1fLiawhr3oNwcFb66EAMKAdVq+MrQM9OUh7nfry+Bhiyx/gaWS
cTlJ2Lo/6jGOMpiHrQeNk0iURAmwxdrre6PvPAEBsFxj6Ac29ohLr0N3UXrST1Px
sCBqcniupwZsXplsjr0VSwWSizhXiEQaPuIz/oEwN+Oxar/xNsW4LhrBJz0R1/Tu
BryqBJCVzdHuVsKkpXL+BpjtnUSRgdo+LtXnOMzKIJalU1gcjIA0re0vy7kmLwa5
Drt0YF7vYP6jAOKmesVKmOLhpRNBWBYHTPL8dm5yKgUm1N1KbXvLZJhtHtv1oiDN
iXdlvvkfAl4mCF9nE9J0isVYXE7Qw0jwRObg26KwiVlWsak2qwxIsYyM5BUFkEfq
Yic3LWkpXzfZXKGrGqadMD0zIYqU6hlsWerqW2JMwdHQL22j5xMhiLUD0KZqaX2c
9z4bGu3DK6NjUPN6M08jnfepnNC6dt8fOMDpPcJr1QXGqzSvUwMfer/VK92LLok8
9TXnXogPx0wPCPzSgHyqF8FTWhCoFu2Kpahh37gpq415qKii/q7g3Ts7avdtZx8o
kZ5ORozAyKK/30kMXkPOzt49cZ+qDneQJxLQO77ttlFJ7cJeDrtnTFoWtZRekkit
2SG3PvOlepfHj8HbHjp40BREnwar+lLRbkGPcsrDTL0SmXThSmehQ/scNkiNdTMo
rjfhwDG9eptWuaymxTUiC1hYU023CTQr+ahARC+WB4cUc+d66Hnh1fSn95VVoTZD
PnV488s2XE70b2Ay3yrcW7ATOKr0oCA2CX9Bs9ervyy7MJi0F0FyZaUx9Z8XIFrT
L1UPZh0eDzXE6UQ5VJsXBhdJCmkCMcmPwh3N5NgrC+UVx3i6/bs7U3BOAtGtdvpi
PM5hTpYUj1K9OpTjDpjxHtJdxMmduIB2Wcf6xC896JRLkjfkNwTjLIz74HuxW9iN
+wkXW+skR6MLEo6qqX/2I884VosQo1Diuj/cmqHKZsPGj8fyW5E0WYfTWNJUoUNV
mugIWf1FG5cYkXWzNUv/S47WQAXPbLRWwdE0p48oox07t2PtA3XII4pJnueaV85L
2PdgHh5it/pwNqBXyDgQ0W0IkOqzB6EZwhoJHgr7PpIqsxAHOwhHryvU60NT/iYt
dd4c8ESYw6HoEoLX4iSnXuY9diOUZ4fCzyS7iC5jc6fa/zqmZMxAIaAcDRdQvcj6
pQBD5FQf5KN+9aiUUlwHJNyKIJhVpV9A9G5OB6AZWjShgPVw452XZEpvDavtXQDC
YWHTP3Xc6QItimEPrhg7ra2DvmRka9otARk1go4RffmalbKXDWS86zSjFxvqqOih
KjjELnH8tc+Q6ELk6T/SUfqIyNc3t5OqoSD8Id0mYEGx3dHTIm2qI/Fi3mJUxVnj
7XKRVzW+2c0Ny1OUPRQx14M3BnMXwBQAUkRe0e6EkR1DVXqtURf7OuRF4xcLdaWM
MtMHXUwHH9ryRiKCOKcshYtxEWPG9siEYMtJHOiThmdwwXLi83XgNs4GD0h6K7gJ
KyufprBImeVtdIEYX7n526di5O18lwhbBk/Kkp6FCkHXOu+6djnvmO7YUJQInXE3
/uUvUEI5hBKZ2P1SAvXvkPHrdh3KMSejHaFDD2fkmSidZg/BXohB3fio3EFZXfd0
fU1DX3TfzRhumJkk5XH+qL9P6VUG2mrirwcIo7QE+lwxiyKcXP3ZWOjYE2/AqLWs
ffwA7GK51W7em6f15BvfDpKfrQX78NF+ijKnJyQIgmdcClctPUgvexAl9OGiZFT7
M714R6aVmQLZZOIkshtHr1ZcFQAUZTw91jTnJdkc8bpIhQm+tZNaqx15W6QYmM5i
eycvREFEfzsRrCjWlEF8BsUFn2GLbgD6pwGlhp6mwPhs9Tm5dYCaRj99q43TR/UV
J/xmbcASabB7SvOGX7XmbLMByEKQisibtRlUOrh1G8AmoMHyKLmOOLTlOHN3YbLs
ql6oxrcEiksOiKzijeQCsZ3vIFV46KvJGyvpQsRIQ8M9u+64ZWWV5LQ9ItjpR4/d
WmB0TumixbYAySffT7w9PP7BpSZVqZPSKsE/QeYyIWm53hkZPioPEJjHhPvi4BuU
BrZJHnf9Ssm5Wg1bg9qIHa589M5Ddi89pjrrj70ejZW9kqZyIN3+cuB0ePmt5Yrq
aDFvNveqgeqizG7xeECZ6vKEHSULL/YmukZzMTirwDVoqGfLkhBeA+jQjIV7Tb46
q50Pze24XB2VpQbwmZs3HQlt1ix9rN+cKmnZWwrfebA0se6BpGrDo+JvvPK6EduO
dnC+ihr++PaUWzkn8iwSQAVdXkBYJqrdqIe5EXpJu6jp8aEB/DsS+0o29GijYqUs
57CCl/ZVgW7zoSBqro5wILHNEJ8CJgWACTDIrLEJzCTwWSg4QjzG2JWuh4LHfQv4
pmEAa7YKhisfAPMbX/M5c6bUNAjXxVltt0Jwylvxd02JNCcR8EC2ndUVg1hD88La
dSClat7ukIz5PVzDn/y06UYMXaOfEDjpG+HPtLZEh86NcCgg9ScXqFCZHhe/bNUU
zMhSo3mrA8opb4+uMSlPO7WLhDTPYcg/pndpHsVx4M4KlnhOYWBQStSPYmu5IQUf
cYMr93mEejB0y8FvkHJFnyW12ZUk4pvwxwnbgeiUdw8WIiW1xy+0wn+ZtzADK8/+
5ih9KxztO0z5ErTQrH+RmfY8i59DUnrYnNtrsLHCdL2IaWvdiOVh5s8jl7K4P84L
N4G8m2NAmUnCjUcenAPbI2wqOZSnM8dzqyqy/Q9/yJ6SeGLUZGpbku/bWih9JSDD
X4QhBkZhB17EHmgweXIsETJMyNDEZrMamt1R/DqlYonpI6AxusZkrA/IepQexQso
UlMhb8UlQMfXBef72ieuBlsF+lbvJkuA/6Uy8X+E0B95mXczbUFZgvn+cKFr5O9Z
tt9Z8Es04jsRhg4ZnNUndkAPK0QcVlITrmJbBWBITtqnjKuvHNQu7Bd4bMAzVKGd
Dd/FKSoCK7uFVNiAX+Y+/4N032NFOt3+tMq9VSIut4ADjaZSfG8CKE3Gmd0LYK3N
4ASQ3o+XbBcjKzgzu8EbAMMsvSVHRaQquPhzj9bymh0CKqzxeakAkF4146SyuZpV
IxZ+reiD9LhtfGUoYGrNKktLjFK+oNKSzFOahmOxlg8OJYyAl0nAMccokwy1G65E
21PTMIC3bOrg02gFrdbbaDwyGbpKkwxsCKcb3u07wJa0DrpyvsiBsLzzptAWzQEn
NbHhZzyyBEfks51VHxsFhGVUvn6HbLh4yw00wZM/dC5YcIKd2BiHsUyOIv6xEzP2
sYGajsANgkuAOPQum8b/kSOkZnOES/8aC1V/sjB6v8b57bnmhVIDjl9fcQ3+IY2q
6FKNvbfJqQRH8tnOxXUsxzkX5ewZTPwdWGxxI57XUdOYSuFjhbcUkTs29Z7pkk5w
AN59PiWi+wok75t8I0qruT5qzCAgaasAr9IS/qXUNcECHFPiZhJfBHcObnkUAiB4
7TiczOjBz0lTkeqlPmb8OAjcLQztuurdN50xOoqzQ5UQ/Sp9JbEDfOm3y2wgY1yG
ytBN3Pbo2D5DpkCgAmp97ASLzQKC4jnttw5xZhigpniUUcNuf24RIHVScdpRxPgV
mMUI2AeMD60WY2jIhvrihMLMSYRn5bSV1/3BrsN/epKrpGlc+QQNkmLeAVcKXSox
BVFtpn4uq9lHNH/YJtYXoKg9Uk83KkdKRLEjEIJ5iFCaj3+RK1jL8i4N2DGF751q
BlmaPL2ai7dZ6mnBzbZbG5SvwGZdcHlDTHAypP0lG7vF1Z/sZay7Q7r+7r6G6BPW
A1WLnNxpIqzen1Dieg6vPflsCzJbuB+UlXaY/BqVEyEHiI4JESPtBaX+zdDQqwyW
rxFZ9LNg5V71wnp7M1ltM9NrgXBHdNtQa3DTAatBMt+w3ZSoIkn+zs18IuYpY9SY
pKF/YViq7sV540/FuWS4zejcq3gh+t7DISbvVk++MpFAOTiQ2zHiKTJMOxpR4lBv
qVV2AgCpxDDFThRAa1icEKTV+2OicKjcQie5p7eWRbbGOwEDADYCVCe66BkM8aG6
DgPJ8a4SMGHbTJBLmUApWD3Ml7uede7dHlL5bHDRn9ealU6fO2nxHPxaBnTEvBLS
cMUzf+SPjjm8zkwebJvfQ8WPXNyxySGcfB5Xwper2UfiWW3BkQkHRHEn9WiJvFhW
qXiXeebc90G6d77uAF4FesI3VpY04ZRzDV53umNMSC4526yRHMk8G0eh+RZR5gGp
vNdc7afut21q7aHEbwkyaa4nSwd31wFmGFPbUqBB1sUJkcBAOBGnmzBX1lEO3HfL
w8V6w2anS79JaRs1JSToAHaTOSlEGG2QyoGJcPA2cpm23x9CYAKU6DVyPSZPCH2e
rPCecQV5gOcDCjWqTx19CNyTERz3hT7XAiMFqtzg05h2PlBWqn9z0bzjD2NcSBbr
0tjH8yxy33Ri+WH9f018w5x9B7X+27Y/bk/9GzNxA5Za5zN79tQZf6wtwFC8oq6p
4RtcvAffzxFEU5NZICV5GNKlY4oHyD79v/yiAL7Jg/RP35XKN8wzHJZKscZoGvJk
11qNIvTSCOrt4kwhdD08WgrNoC41parRslbEB2NIRrNql7GpuCNGYxjZBmBXaDPF
DgOWDftzIWYTPEPu5JrvocA7la5xQdzfD9RmhrKK65ODAzO+j8ebOOAY2GQjpSQY
nXFX9ZUszABVwKirODdbolq7qz/NNMaI+vtFqMCU9OYM8llzf3zSDnk+eFaaSHST
dKGIORNnMm2D1HoH8qDSs+qJvu71ZBDvj7sgIpbQvRrVha1kUPhDMHxtThejxLTf
WlCKaip1D5XszZa0+/iuh34s+EHQRVl7KsIbF9vkFeqH4/ac0m5DiwkhJ4rkuKYY
kB3KU9vPqF/jvnbFrkLw1F7umiRD5JbsLHoxG4QgNEVvImRhTFACELkf0ItRh6Fl
JAgGotKqvgshB11PmOSc8poTjp5wHc8pm235t5UqWsnk7Kf9sfoYRpO24gWJxUEZ
Md495EPyDuFMYYSIdHLkLeu3ROD28nZQyk99tbRm7+IT03amGYnQTMTw62tkOD0O
4qFjHXKvWjvC/tZFEg08wBgV171kw1RWh/03ucaEJXiPUIQLGdTUwV1FUO7Mv32H
EjCW18lqrpiohSnMFMTGH4nmSpRvC8D9UZifsgoQ8pS2tCxVA7wziEzxoZbIKCLa
gp06PktjQOpibO5K34RllTSGcKtFyZHKW4Vizg1iN7Zkpj+5Z4Y3gBwZ8tzS5taz
hDeEg+xDPmjjgSoRTSdUJBU4bZTenrTWYkKDG09tTzIrKW9dWyIJ0vaZVhhWrrM9
sN50qk5hH8zI/gPDUfIBGwdPMvhCCW/hZ0w82HN8n/JPj/es243mGIxWu9o10i2y
UvebYJpByiMfh094NSt8vf41mIQfZ2SHFJBXcYeT3QkNTZBbApYzXaUmmIRHNyhT
Wnx8tZxIKQ3rWkVMaXqhck0EZNdMx0cooGaL7QMCMQ6XRrL6YDp63yVetnz0d101
9fuTHVTpcFu4l5utYE5/gdLo9Cx+MMBistZCstU2mLN6xNnzbIE+drja8JKYUR8H
OJ2Jvfd27JtVYglMSXlXtG+UrgX/UO9+1fpNr4LgTCwwOLC0pQuCCRGgInAmM4Zk
H0FWwvyRgCDtNyFu7HwjP8eRTforQPBAvRIVRfit7oDbj25EABgDH/1Hd1AEpeOd
brtCo0d+JgprXg0y/UYdhxQIElsaR+vmsOEMV0B+NtEzJNs84mXKtpW8ff1VfusL
n8kvpjpM8dNIOuUtTnTRnP52+nnQwILCHUAtaBp/+9rbORlHBjFjo+cfeAmKsn5m
0zaXYtXSeV0UCaVc0FdgQ/4NuX9n00rrkKjg3kNVlEQxtNiwDtpwG1+g6Y0Oe826
lT3Uhx2bkb9aPMXCxnJlboqTNmGN2UjQd3mRF1AQdyy7b2IcARVKiFQKdo2kKTSz
dznY4w2RREsTUwD7fJy0iBC9a/DKwowunCWghyAa/879m56myV9lnBbTn0CpfuEP
A+5yrJW5+zDIdZA7acgWkwCwOeLV6lokbfrPcIljBLSmXAo7NFO8cWF/TKQEm1jd
aLDraiWl8Th+n2YcIIXkskvs1qDuqYTKVffL4GgmBzdPAOZft6e5SzNUS9XvjLAp
wmp/kQW2eN/eWu4x522CEX4wb+SKx8rUd4p3YvbyLpFeau4qFmsKSrRr8hheAPrR
yxJxpUdeD8PSd9xo/waEVb5auo8+esrnXlfGYiAUHoPqVcjpWOK6TqF+Rq11zrki
MnHSJVe5YMtQT7tzF+TrphHH3xvrMEovTad2iNzn5ME5TfJzdluVqFJoWTqABlvb
MfyIYkk97+B7BxdvjKWwD2RoCgIUFl/B37XqcrRfKVUntLWkiHwFW7bk7uBKnHpy
A0Jn9jDAB6PXazszKKPm65tLggPSRISMqhqOeNUqgRCc+Ly0ZD6PtX253A9w39Aa
uiX6RqUNcu9PS994hZZ1hDYl+0WTacGQIwfBCO/vLTz7TIruMJ+FS8eiizQO6mzN
NlRmGFZ7A7fpsXKgK4xgiyhczQjPNiP+2HgtkHN4NRjKXSj2OZyY57x0x2iVgvU2
GNIzL6ml4jbdPrbLcczJHJ3XcDfs4DoKm/9O/5U8ZV519MNb6zDiaHx/t+EuA0h2
IMVbso5oYr6mnK0WuPW2sp430VaklpDIqhbcvt96GLnNIrG5+Plcj4aB09LEtU7B
r5chHqI+YJN0o+GhGgYcGUYE6jSlNNWPfjFgAF++6A4dOCDNKT/UmGLEBKLeE9uY
z9dG5g4RHdhJ1kXf23Ev20uypz7b7nbeMhskvsdtR1fKkN5Gp9lCwsN9tpjO1he8
8A3b6xu+5TwzlzKcw2JmqUDzlTT9bJm23KGjoxdBa4x8znNRUSZ5HGVNtDx9WPCQ
3DxLxydVachjkcJmswzIDxGUAmxun5q8P5LLr1hS3KNzHypIC/vk/lJiPkWFRMPO
ABE2OxfmZ9uMGvO3XnF/xDlmwra7/09b0r/vkYzYIbZpPXf1Veny/hiW5NASBwoq
EB4ud0sOovB8P+bWd4O7TaRjFlnUzOxv1Y4DPgnU0ClgpOWpp9BRFIst1g/ZKW/1
z1oSagIUuom/MBCS98odrXwbujlPcqtyh0HWLbyn/aIuXBAiWiUD7ZgvnbX3jVBS
+vG3i1Dk6hyMakoIP1fye2IrYQOBIGgsFgpcifr1jazUjOqniy1pCIuFlHUy1qhM
ALAjZoRyqJZTX4ZZE5ov2g++V9d4mtCRtpqT9JO1mvTmt3EcKfJSyecA6SrZCEVO
ywq0XWEwXyIrK1IJk+Y0iUlw9/FnC9ZtdK/gHdgr8tBdBHnyc6YOdM4cWUhqwpNJ
WhbQ4FvR9uZ7mAUgtGoYJtxR03V+VRwm3KUbDCqIHZs1xwRlok2kLA33Z7f3PG4k
CeHWbcmq4nJC83jGg1Rd2PPRx7JkAD8UuYZdXzhw9taOialybPGXynF7dZyqpXug
XO6Ju9VZ86eGB2hpLiRLL/lsOmEStenG7xrpAA3JHDKE/jQR3aFoSS2Ogub8FZF9
FgZWtXeN4T8OKCvIU6UxBcFF5oxfGjbfv2HzDttjTilByyO+sMXX1UBt5sdKSWJB
DuJMzTEAPI/Lv+O2pVr5/J2suadWbMYdCe09QjyrEgh4C7S6sPobyNW9tduBHnUx
4SNAeGW3BPPKphvd+9+5gFsIdHLLCMI0uBOO0tqCXwhp+58xx/rvf5/O2U3xSOFp
PNSrQ29oWQM///Nf/DKzELlxyXnJ/BZoJ1rEfyZ2FB0QVKdndk7/tcd/1eR4lfap
y9DyVirl1WQpqwb0CgP7FYQjA+8F7sMpzbWHk9jYgpgsgYIj3LQEHv6YsVyiQkKE
th2J/qDQAy7dXxzkH9NqWpsO8q2YXqrSB7rCjBpeyLe+13LVvIrax+kYNaVkey8X
oSB141f5QO+fAuHWuPqCEwxQL2d4l/0Ko0oVszyb1UAMJES/H8ulGMkK4M9JfJMk
xoTvfQ49RWHwyLQoXhHzfMFynv5xYA47OYpDZM96V6XWsv6i4RFfBQX8BLCvBp4n
6zPUK8L7A/hzcb5KwQzHzfV9pHJjkRtXlpukIWdEjRaN8ZEdQnDx9hyvIinphFWm
megbtRrwPAbVniXn1+PqTCwJcOxHlcRz5mEObIz0IEfJXQrYS9ZBrkspII/IVmNM
ksRFr4EWWf7pTMo0YGWHQ+w6JK84FzT2b2m+PuQpU+XYZBfJ1sJbUqHmdqmrLkD9
rDTE0mQl33iPBN4uq/cC4fKYR8cF8HmHDN3LMA9/i7CUHoWyB76O9sBWiRClbIc1
8xpqM4l7/AIFv4JQpfTOplMqRWTG3/FwO02IhpsRQWmKrSd5NstWqQftRdV2kBLi
MiaIAVh2dw6NjQZnndoLCb7oooygGe/5oJ09PrEPQxiG6JjmCXWYbOjHAIY6QZnI
PuD1MUYDRNJRpwk8jrYLkygGUtyELuMr9sh3OFPdxiX3KQ5FfFZ6LWRR1RCxhleZ
SEYyAllA4XXJOVS813JrLVkavlZ2hkongEerXt/F1ixFcXc3a3VzRs0PpgSyswGi
02yI0bV5gZuE9W6bmsyiAaZ/5O1qH2UVcZa02xAiZdb80T7fl4MDB14zjtOLf3U+
JFxEjVEtMascP+qDPlMWOAGxKHVaESej10TXPPO00RaSZfdVTLo5h/Zc9U8sXWmI
WKmY+R4k5ujfocMh35BB01C4TesEMEKv224/j6JFDiBuSb25+j9MxDDIUbYJCrbB
E3JvIU/XW2oYXcgZmVze5jLq6da4b5wFr1sNSTCb8Z4yt8uUp1WW2O/UwUAZU38a
zwSdrP7tPe5qM8RBZMe4ctQkPNq2FrKuS2XPp5INrWcFQazmrAviLYgpIk6i+nQW
jqkHkRuPLHJbGVhGo77c5H9qPNrNeZAlSf3w6G9cOyTUPp12UK4ZpXWBus3KLGWZ
DsNtm3kV3i4AX+4ffwGh+PCPBw+ws1vUz0mpsvntv3pO/P8QC8KpbXV4PG0G2h5y
lYJbACUUc5InW/FwNGxCyf+XrCeZ7F9HWZaOuw2ADvvEj0aJgM4eT/kIfkie5HP1
yHBV2q4NJehGMrD8GftAr5VShuyCvhqEAwESTK0OxRNnuy0p76PupFShbgmxoMHi
NX6KchYAkncKghdYa6oBmTT9HyHtB0tyKlMBCPE3kHdxkWQI4dr1wT6RO+r/ttf3
rGc0dIqcXTQNtK1igSu9sSpnWDLncI00CBm/HAAuKeraC9ZYy6gjFAIfWp/Ix+u2
jBXrKMoUaYsPElZIa2Zux5RP+2DX/kmrhoSl+vjJun5Je+sxQGIKQuJDnc3L+71w
pPmbfnFSuoRA55fhTjP4PlHraetQV+7Rgb6fTnlv1j+WWgEFX4RKvJpiDzIczEHe
eQkjX5slhbEeHEC65YFF9ZD95cjqT+pyqhMqDH2Nz8fwewZhL5v1ze9lMK92xz6f
us1qVkeuqYU8iegBNhwvZvPFRrhNx7CgXBP1JAyRCaPQn+4DRrFJ5V7OLnIuri9+
+bZ/G6H19IjmFTnCYBaFhAdUPSVtmhkCzT2WYizrPbhU37hgacYDPUD2ROagFjtu
cEea6gXxFS+7bENk5+kU9m9+CvcTpInSApKoGsTN/o6/nstSDuhGzYRhZMYzRDKR
Zmwj8sB2U0dGgWcKW63O/q4EGMV4UojK4zZkk6WueQOFebU/82VzSHouQ+AejHlr
2SESrCUI1cNcIh+EczPRHOypV+pBgtv3X5G9WaOmu6lB5+0BTY6S+YxSoNQiZQ2f
DCwHjHDygx5Dj5JNr9ywGJogYAhLD9hxO+Z2VpLjNMrqEDgU9IGOv1IXjkrIVlhu
CUEDgimbcHF6+NjLB1t7izTTRqfieaJ4hv9OTfBhQUe+81VjWSBimmrURoE3wr1b
x2VCVTsVuvUOTdcyC5VLpW5F9wjjbCMFw0dq4MEzWEkYiUF4WFUyfdBi9C7p0wc+
wCNjE6yY4D+dFkU/rbgbIpQkdtJktoPmQoGMVWFTOLTsapQgYARGDbABdYxXpACB
DnZsHEerJHdcvXixB3JYpUHLwvxDaaqUGH6enwRcDfQR6FjX1J/NBeTfLnMJqzGt
KBzEKOi+fFo8FJCjPoUB9G0cyW6Uupn5kaDHdVV6ygtDcZQUxW2eZpfDEWp3eZw5
xpmnVt7Pi2oBO/lkPgI6LmoeLJeKpMuJegchzBDWadWQH3mgMCcpk/TvnYmAuhCB
AvhubV1hl82r89EIZAyoeYI+28xghvZTtrYjAZVRS/oMGbxpVQEysgmY8mtm/Pek
0XPaiXCtDI8KzNAz71y6dPAaITG9sQWCsIwLDSiC/YLm0XGK0ks6avlkZp8QLpnU
TCtOXw+wxLl46fNQuCbVsEwHw29ubMLGePzC2wB59mnv+HTyj5Nn2vSNH2Kv1rdE
u3oM42MRWo4EFV3iJWzpDrMzFIzlUKDXyhZu5mzXj2kU0d9exwsmcwK5C9TvFiIV
xx2ElYVjhf8IjzNI5z6I9znxXXza4RYjvaWFCTiyzR7omL8Wvnx/BAMuDG1WbAc8
sA2FLQyQsngsVwtbZ7sZEnasWEIfP+rbqZ8eHWOU5iYkZ8ED1iauHHzPQXyubWq7
1EjTBasgyUMabakp6FRI3zF6pphWxLmiy6FYvb3qeqeYYZ/uiSeVlqx0p1xELA2F
BFxa7jPiFzKKFWB6tp63k4LKOHSO7bRoP6jXWj4w1r3N2de60TIRmySd5NV/4BEt
kbv8+yOreihMtmVFUeJS5qKyj+qXqSyUSY9WRQ9Ah5XSJw97igkV/NOXez3Ey1Ug
D0oNZR2o595VELzTGNbxI7gAq/dB767zes3XnMbLbhTGLpHC+08F+sF569AzRWtO
Sua2jpQ8HemQdlOHw9yyQp9gLhZA2fAhj57OvJi5Cpyifd+hmi73/qD7rnnq289h
8wr1k4A+IW0717uGt9vFoW/NcJRUUdhQXMpBaLLoPtTtiB+Gn0s2MgIEkywiefBz
UQp24gII4pt8xU8tnkt0Cdja22fNwxTggAqb7nFgCZCRX2qyTDwk70K+d5r7gpCh
54oocjDBEBBRPU1/KDLhLbf3TIgBmIKodWxRcgm399+9gTY3S4j1GtxGAWUae58T
qcb/XYnRFNrpu8qDLYBeESdwINYJUOWK3Tq9IVPjnu22w62n13n2o1+9moUceAgF
KLmA0S2iTj4bUw2GEZHApfY1z8zJd9jV5paOAKZGUjfSx1PxMT8785I4KAXw3uVB
Q/FA+lIBpDfyIqic66BuiP1y4a/0UqpYuhMsxW9O/yiuUAlb7uZ2FeXpkpkwRUt2
9ed3G+r1ETzwH2VxXiHsdNZ5d2eyPDKJLK8HZ+qvwrCI5BWSVRRWKHDqI+EPkRYJ
ntx/UaoEFlres6LzsdPKPliXS7VSmKaKNkXYaEG9JnTZ6hQzTWwICVGMwp59A5yF
KZLfg2vWGZvl94XNL7mYgmltUC2ef4YBrQxD8jmP0kPJYIvHm7rMVZtKgPxIGwYu
qIdtbYDpfbitb9lJpquV6pu93ZhRfkecA1ifyAK6bOdXjwMCBv8ZilkQ2nZhw2OF
SZcV5c7L1zR+YvT8NzlFuOyiuXzL5ITGAylEypx8EYrt2jxMWmRiq6r7PZkHPlp6
mQY2e9A3/qxdn/EveMqu7tqSScgysP5c7MN/FbmHDAlxRTjTNQT7LbftM7W25srZ
uRJ+TB9wqjuNb1e9LT+wU/wsFA4zeYh3SRvNmrInuMHS/TZu1JldUMzEtm05BgcK
Np24ZplWjj8r4X4/U+gVhQ2zmZPxTTbU8aKe+VL0CY4tl1kLnofXz7+jO7tvD/dH
TAKMRXienFjLR7FG3wSEyG0lEB26dL2JBQ3vPwTMw2JIPOTTV/GLgYczQN8Y9bpV
lGEcYfEWkraTM6BsMyyFIfQTpvevsNmKy3cG0DFikflYhvDnbnUrhCfWOT2O5TDo
zXwQ8PeKK3jTT/MrsLnWE0n+7YYgcVsEXO4TEWcsBPPge8Id+epwMMS4mIGV70+7
gx6ysDcO4h7DFZOKSU4MUH5XS4SApcmSZFgormobKxqA0viV9Wp7o3Hm0706JeYQ
lInrWQS4BNf8TKHgQUzKlMj/gLc/ZWqD1jdxfdlByKJ/SqFnetTeu0JM1dKGT402
0cBigNUaxEGnIny3yqw+9WkmPC+BRrvp8u+I8aI/SoJnHZBSzFyG1k8YRri3zFB7
w/+dI67bW4rDzZAQLc9DKjmti2z/bXr1hh6PhcdyKljfCwtOnVpDsbJrYhGyTlDI
DzGdWml1PtuvOOvWIA/TyWCVRTWJx8RxfEnZH8iCit5MyUWHSQUIcMgIJwdYjYWq
iYLhlHJt4155EJh4SjkLUWPyfTuAX7SGyCf1Nf06G3fpZs0AwEhi7I3j1tvTmtLd
dlhHWjakK7pA0s7bS7O+UrpN/LbNbMFqTkUCxxzBslXE5eI8gJLyXYJ8MKckXktB
/HCcEyx14tA7/lYKHRsw82NW3455th4Xh9a9X1BIp/ps4IpwuTU/pThXAZepSOtY
8x+0kLvIJFONshD/930T7MBaHyFhwIMEjZV3oVrMQFbjEbcR+EDq58vv2t49851k
U9ugTkbdBaP1PVt1K9gcHbpncyGwzuLpdpn+2/wME/dFSbmV7EFID5EoMTnmnb5m
pk5zft0NMIp7exMbzdpZZBe0XT7YBojbTVginw/OKCM/GZHiSQW8mylBxr3GxKeG
qZKQeE8PhdKrwW5C9wkR4LGZthCHYITBDtrHA2SqQuVu3OUxeGyBBrh99gr14sP8
7J4PFJ7xsQ25zYKpqxeUmtggdlwdUpueZ7AEe+XejiCorS8YcWwoAeavq/mZG0yW
1KGusrY+/CS2IaJA63arheQg64akGP50oMUc6vJOS/B1DZHy0bk/74Lwg8i+kFHX
E5PIPr2sbTp4yGeUnK7fyjzgK3CMoMJlqrJpPzC8HXZ1Lcn+QYWLm6ZU0OTSqIbr
1ewAT7+iFK4Mx6QsV7LC5446lZp2cOvFYP9gGAF6R5hXjHuOuzNVc25s+ELxDLF+
82BeYGCT/NQ55MSUCsd5J46QW+/UiVq12Ta9nN6xsntrWsYBeJuxDqzKG4EHE8KC
/bHvFs/qX+vJav2D6Htdo77M0iqPK9tJ2DLDBg1ahSOMz4SqleCSxhPNRcL5PTXN
g9mFgH9/Fkt4xgrZietKso3R5aFRcr7ihdpJEoVTY8KOK1vppPFyl6BhOyTQqPSw
tT1JfyZOYXlPMIvYTG4Z3z60+QjNhMD2Vn6eZq55sWA/Q4gc09AsW8vIwOBO5kRx
Nmi1gw/koJDKglAbpc/UClsGPexVxRnzuFukov24PiKqwp1S5zx5ZQG1hAHoroa4
RflWxjKkgGI1PzLyyU0vTNcOwfbqAs76Wyfzlq23i4ANybClVnz2muB4zN60rX+7
+l0ZPoHPIcHIolfzofiHptpPjkPFtG6p2YNy3Hkb+t73Blp3b9MKL/HwC5n8QKF7
GMUcgzKRhxXuDQX3gqwU+L+uQ/whoPgasWxEox2baxInBWFpQfdtL25JbuIWcK/n
8IhMMJkmmsR9prWDbMtAe08qRJPZYG/eocb5D4mgXSMIMJ2+MmuO8Ffzqe6l0JsI
XPzns7YbSUr03QoY0vEzswoHrDi1K4+o4wGgL2JzWXMCov9IkGImJq3qNaqwhfnM
Mcj70yy+bWXnLRr3lugZuwBtfNrUtGAo1eo5mX7fxrQ/hrYPoY0Z2JTIT1M6ldAz
6LCN1TjLnhwOSExzscfKtOQunXwbByrAgwKPMDgizfOGWNGNHFiYLxCJJmIx5anj
lcdXzner7+eZyjzy7A3eRTU4fddx4H2NnpXHNe+sfDodf/AvSg3SFWcP/zYmI/q2
KrdY3qLFnu46C1GwpKIQdSEefzv5d7BbdeT1Q9R9oSYqDPRo97G9umFP2Y03t4tD
0kTLl0eRKm1GxAd3M5kdd/69GHYVjAaY4dPnIL7vPjRgjCMtXFMvOGhRXPAnjROg
GTQGdx9FQT2JJdIqWr2hZnMy9+oozwWHrAIA1zNpUXBZRUafjhUSDoncz6g29q61
OW2hxquEXr5LBd+pJO3IK01Ev5WiEd0Qn+WpbZSHOsyAPPOXY/NoTCUs9DpAhkoI
9kSrU2D0VNdeivOzxIEuM6uSoD1kZKnCsb0ijgQ02z+ZmdFrhoFe25oxuaV0YExg
X9lHbsEI5yX2Wduj4u3s2Mn+ivMOAiJ/utZLL7db4wfqWaLR9qq92Be45XqPMbxq
4J0C6Cad7mwOXVHLICA6k1TTDARloZuLBLDJVBqTylCb23WMiFgkqesghyH4u5cZ
pfQPZWRpt+WWQijtEnqzttOgduMtUP+0RhHzpRh7xI5BSEm1uiihOIrvHMFaM3bA
W0R2rroVavrMX0R8dayKw9Fvpco+UIMj1p0A0tSoWPXP1wGHLA3lTN3d8SqjJQSw
8XYC1LvyQ0crLayl5sk+7mzoPZ+II2c12bRCjwgCAcMbtSxsefkm/0tAXZW5ryTI
3zDdAGtimJCsO+NphaIJ9vuODsK1oRFyzc44pqI1KKtoJKmPtEI2yr1W+XRydL2q
T+3D1DN38saTZCrwaALvauKtXV1I/M+KS94wQCM+Lpqw8AkAVutY5MyYr129TZzM
cPJ6NqJqGo8WXpsSyryI4f36S397J3wbh9U8a5GslgNEQAOK3yoIraM8xnGLhg1f
5gHfXEL0T3dHlEZbpn65mtjI6RO6K3PyjN7ROb5VjDUqdbqInxFhXkiSmjmbL8nb
A093ssUojM/P1rffTtWODAlcWF9p5tm2yIQ370IVUGKF+g5Se1lgnLSlYTc/Xbrl
IDgBjcFdxo625guKzocRRnSNEb5vgGlfBZ4M5HTobpP7q9hNn3mSiRBNY/gLyz2G
3hSKkfNdwmkkHUlArwBuSMxrhYLUGbjGpyrEPwRQh4OH/AJQb5TT0r464q4L5JfP
HifJ30uHQb54qFtXfCBP3LfxEeCdhw2dAFnYKirWi4kCsweLVqLLJVKZya1mgcZD
VAQN0NhNYi8H49BQhzxtSMCfwbzxgAU1xJgYTm61aw6sesn8jyvbzKp9IWRYANqi
FJ651lpM/PRHCfZlG1GDsYbJ/Aa8QALjQ6hJ6HFX6MrKoeFmZlyMA3pNmuXX9bMH
zQmr0VCMSOKPmQk7yaC2UcQYRwvroFVb3WuGVXKZaxoli5lnAIcEGrwVd+O6gI+a
IzF/BBjDq/pnmPv4G4lCjVUX/fUCtqpn7iZ0LKMXlJvt34V5RpoYPoJ2S2iztkao
MYU0EKYDnlMMhje+xvssQRXsOOih1fE2Y3kqJyMWezE6IZUJ390e37VQvRnx6l1T
1U6ouNvLofROhjIiWeYza2UUROr7egpvmBCFpfQ8wNGFPyoG3dW9UQp7qnjRYGNj
eN22PrmsxhoF0Tp5RPkZOkEYZelaQlVNpi3Cw2+1HKtKXFij85VqCbL/LegvJCUS
k0NGERYo70iU/71dJPYrUx7JFHRRnTfb+8qTreZGXYMhTd6HjxQmSGWR6UInIKtt
erqBvZHqmYvc8HS4orS4ApSOuOJYG50H75Y0MpQZXEb079IxgzS9BIQVHtawb4dB
/rVfCZR9MHLv1rhQZV6rgbe4r7LbpM+A0RYmlhQxyHjk4du4GMfvIvu4SqtNWSjK
P38EFPgpKWeyCWTneTWN6VXcrQ1yOu7jb2Ls+JwEmDNlirublKygogq8kyBAy442
DAKkgNhSAozGpFzvtunN4V1BcwwHA1tL9wTGWvgwlyDVMe3CqUPm7Ux8X4mdMqKK
+g6RrPrQ21fa+M/EIrxLffXyOYMeg9OIXPCYIODeIF7vLtgcQjDAQxD+c7Dq0UPJ
Ltwj6WajpVJJMK4O2oAuAJwB9QyohuoJxr1pQGWmGcuEX1DklVPzbqGgoXOYG7qX
/+92LVVr1k1Eso0pEtFqbe09WCemqAatwL+h3WGGGFFk1/2L5H7O36J6nmTbTgIr
ImwYHtWe4ZUTV21kEB8ANoVE/MngLHzoBVRFHmhC8n4th2yub5Ed/kupOauh85zG
/3p+LolJAh+wjLU96AtOKncEMlwp0qqS5G4GizB2GxUkfJrX/k36hEIwFDcBhINB
2xf5Xjvsb1I2s57b1fyqn7AM83E3j6o8qX/3luKWPpAvKOWxvUjhHjeTdnLjTlyA
4gVr5y056xFB7byhmETAXrdnK5ZApK2y4pL14IHlgNT+HvB5E7G2puXhk6WuyJl3
2hE1OuHrSscNTzvg72A7ky5NFUwyPqxINpovssvfaq3O0RTDHZwfGRJv/cjfC7sH
Ia1MHT/mBh8w0tzpV89G1jgCR8oPjk8u56bpyXme+blpsfpg0hoRjwbXceyGKhbb
Fu7ZOWZtHt/ZEcRf1ytE7qhPXwtGU+8z0ih457sEvQc5OSkAFyvNedHu/ArBzUcX
eQEozJX++YsB639OLCFa/wzV1Qpia+i9K1yHxqc8oAewK/RQ/adUXw5At6J0sjbO
GMi4brsaQbnqDEQPrDtTWLR6hPSlDTseBjAmghzmdkMEYn5QXh/aNCqNHFV3Hm4e
adJEnp3IIYRYXR7M3jM0/FnfJOEYQpoT5/X2dWe07OdxEMzRBmxJRKao35gTUdeX
QF+zZHK9VwX0fe4W6dUbFFcOSL12OVBGqQkgswrlxIO56uGGFhJWRgmH+dF7MWNN
rypHorvPMsShJ58uVg8uaxHc8M3qxBX9HLjoRlr1u2/oKEDcLdaEIZSSRw6KaNYU
kg/aAZDly/xJ8Eb1VXnCaBhirDLELpAbrTbYM0QOLCz5NMOmlNNiIXqidPEODisK
nnkwG8AlELg9A4JHYqs7CYdWQtd6sucLIeC2gv5iT56YTbVdL2snZNh+rLgGzWWI
L6DczY2WLkFOdssy14Jct5ApXNLH4kkhkhn2cYRRbI1fRLep4z49kC5WufTDnUi+
O7cWcJ0iF8rmqDG/KTC6XYh9+WHEeVsFlcyD6QzbX/KZ+778JaVt1TKGcKUpfC2H
+HU8B21qgroNxZReaJFHf5AY/Ne0k0+6qke3H0Bpatgmlu0lb3PrtyZvCCa7OWWg
rDxK1jW+dj358zUXkWt8nrTWAIVCod/M5GsTFWcHJViYZDxDVkRjqt71CPUBRbFn
/Kf08c2uh21HF6f91AYlpGARAAVJdkkOnYAoFXzz3Sd1nMpV3T7IEzQtxeSAccYx
hzX0nPnAQMFBQrecdcpi6wRjdv3L8Zq4Jj/2V5rxmhoaTXISAmUFcZYz1yfuV1bA
pFcY3JQ1SF0ndgv/yqi/qHVjDun3xxq53FhueH2RRn+N4D7DDV0Dfz9jG3Yx4WNO
FclW0PVY+Wxt5XLCnPHSwqTp28p6XfjC1f+Iw4fc/IlsmFzpgNm1xeWyiV2lXngS
8U6G2WGxA7xh3d7JNFKnrfPfZfxLQ8PXvwbVA9cSc95/wjcC2l6l5U38HVeN4pFh
E78lHWG8r/WbkgAHCyqA9HhZyfm4KZznKldslQ/QDs0U+i+iCOqg197hh+P6w/b6
nlt1lcCUDHLWTpQOSQ2xdMc+zzmnuORcbyFqw8LP7IohPssy55l9jNM/2F8bNk3G
4B4AYnaz7CU4BdmMCPog37ssr5upkXiC4px4xBfq33OhoIcCupqCk2FRS44RRM5Y
uGr6L6yD4hoQEtOTctphZkMxBR1orHmv70JDvEH3UeK/v6lBiwvbdPRtGXlAjVRo
xBVwcn2GZF2izsG8z9Yk8mayYGpUvjkHa75IzkKkX6ICWmgwmLvv42jB9D4WJbU1
5VegIYhhItuVqFGGWSwN+41n8kokfqbHWLX7HRqc1NA3qz3q2xxA810aMBoFp8eg
4EtjbzW9amCpb785aTuOTlimOrstg9BVd2ZfKncv331Kqw2JNIpcJqgUeT9GNC3s
cA637sypcY7+ecy4lNj6fV/BuxYcuunFyyzSdnXLtAmvSQFPFyMmDgJY8bdsTwep
63TvhbKhxARuog8XkXjmBip4oTVSK/TRKosINvZ65C0UxCdTcPUDO/Frr0jHUnxS
zWWsEjLvk8ICtb08aibDS3GfBRsiKClQfAhDN+UVxzbKGsNs3va0905J2QXCUPe0
JEbHRQNXFz/Fxm56vT2DiAL1is2z0C8UrC0xRax1Bv/rV0OwlHrnfwxOruCIoth5
8qGJllDBOpSlRrPPocA8Xxk5dJD9ClpagFr1Mx/Jh7x0QGEPeAfCFREcxcEhT7KX
I9Hyzeus10AjPc3vQZu0t1eaj5ua0g4IQajSTiNOfUhGDbi2fnOYblZMizxcU8zF
4qkQTnJGggxC6rIqRmw2f09if4+IGKUsQnUoS2jgoUmz6zPiRj2IItgJFZye/Lgx
Tu1awuCUjSXEnlmiPSp4QJuoXNFq1MbSkHh6RGwKEw5d++mbuiqAr1OHZViMnWRC
dvy5McRt4JNNbe3ZjrMzht98JxT4gfNxEcMzafA5fCxpyCsddzwTfzpqMn3Ysifo
LAMzrW3t5Wydjc4aGDuJQKaIUvykTDAME7wlJz5hPGMXsq33OqVOE8PULUTv2t6K
tV0o3wkWKay6JYsBEKtytghZpYDW6IpKD9zTgB1jXTYT3SiIExHyHusPVSXDjRnL
YlsMsDKbCkYnlTgyr8MIEdFudmfQQWIXJqFYmKncojdgXtii4j+mYdZ7s/V8CsR8
vew1c3T5kjPh6vcDu/hEyRSaJ83CRdNet21RTmxQHo2ktijR9QwrzzUvHIB1TZhS
hQ8c3DEIOD/UjTKHCG6YhFaYWEgDEhvRSm3gac+GTaj2+BkpRI66voeWaG9gnbNy
Y55W90n15Qk5jpUzX31xETHpBv8XFk3zT8SdLCMzgaCqxDlNIJghegC3iBUlUtsy
Y5d7G0JKXwsAM2ic8u0quzZioD4jrf9ZVdNmpeygymG4yuuCYBfy/Go/J6O0GaMF
1iNdox57vKeCSlsEUlEUF4S39RE2Kn8XqFlix1SkFU+kSCunpmu9safy7ecB3KY/
+LmcRzWS/u5XA5k1+eX24Y63dkO6IgpItKhD1vRh3yP7l2ugPZBlrnh5J6JjqftF
BKan9U4rPKT7FC/0Pr8qKEvjcnSNy1PFu4XpK42VbyhQ515W5DIXl59r2RraWhNR
9qN8ZKhDiT/Mt7Zj3yG7YM8IhdGHGYZbpb9b98Yaj1OiEV4wosHQFAvEglcAsJXi
3kzZd8NbIllNkJnnMxVF9Urz0rmOJk/q+WpuQ9Eqv2vdNZdcTjfHL4bQEEhbmmRY
Y3ubBbTEpyk1VWSg3V/vSBzfMsruVTOJYUxPV6vIpgk/Ji8Y1Mc9zR1gPN9ttJ6Q
ymTziVqa1wpUj1b6pU5QerjQ72CBAbeDvsNnNZvoQmAKWhSrs3DHGMOnpao6G/6x
K96n3V8uPBpgsr6dT4wWziaAaFaku+OYHtmARhZ1YsTi5jYAs8Vgdr5jYF+EZzem
IX2fucUltJ8Ry6OwhblJptIBFByosZ8whiD0K1lPo6j2yNF5rj9YtZNNsGzpt9kQ
kIzLmxJIw7wEruPhioRL2Sm8XSUCFlSmIP4HxQ1oHhkQQbJaX1JlYQIepMmrbsqa
Tama8WLRtCo1JF2rX5zE6KCLKF8j3LSD2x0qL0fuN5Ov3Ts+T/6s0KMxpxMVgok+
OkLv5+WR5n7I7lhZBEay0D+FHM2fBcQSSWvUCTwTQak2FG/AlBM34zbtEvWEhG46
ypvnAY2rbUdS9dnJ1LYXcvfxmHwL+t4/ur56ACm8xzPw/J9D5xeJfUIsfDYjXY/d
pX6FvOnO/3jegjwOfR+1Oz5e9OfJZFqe1VZVGpgmjWhPKi5vXkACXC1LmtqS4uid
ubozlZRQJ4YGVb69eI1ZaXNU43oDI0VsiWBL9J0F6xZv0Fo0uotzaeulMrIHa1nj
HL+AV5ntVx9Al6Hx5JiwdAjigOlYyKm5Iqtjj3SUkAiVS32RF7ygIHXRyqYqmasx
8KpJT4QWjbUEee8v7lIcKckeIMy7vo1RMA3rCrSQqqc2KJvrgVMMwf83wgmKnD0c
ckWD63IoDmaagw3zvWwU5M7GbDMbrJ33Tm1D/eMfCjOzi2t2SF2F5nanISG1jEOy
9rETTMhkRgexxBkqXXUDWXgntI+pbJAUPXP/JLmD3eE5KCQLOha40/LY+EV+bU4D
N+kbq0+TcvKco7+jGcdyQ/P0fDzRCbIgZE9X4AcAyve2/dvzE79Pen7FsFp9XQ7H
mA2ZoTCQ7WFv+8lghGVmzsgjGYU38F6R69Jm3Aj6O0FFFFlhAd+4fok1qDwg7bjG
YzZvqJ4rovKxY2kWHhnUmq9wiJ2XPRVL9wAV7LtU9KWW+qp3O+0vkZjdsLrfMBSK
giwJX2ro7uM26Dl8J67Bwu6KVujag7zdYapBVrsNodosnXIlmIj125dww853JHaW
mHoQu8hjBw4qE8tM9ZNvH8PfBUbQ8trWjJVusreehk95+At20MSZxJVqsKFmNFB5
zoNdpw03xG9oO8eJNKBTl6ookG1tAQZBGtJZXdvbpkVafOQSI59njLbqLH6H7VwV
BRMkYLLCkFutdTVWSavJ1Vn7tN7nTDdy4pfeohIhMHZttalBGg4RGR86/ZZfubVk
uuiqcJE2Dk/meqieJUd+WAlcWwiHA/izFMpUKPaN7fSay2oLc0M5E7ORWZQJE415
E5fIJQmoGKE1cpPfL3YQAqVj/pkutx5EkFqgtVKxi1Bw7r3eew/EeG0Q/7o/ii8w
CGrlGaYpe6Qb41SmMzaNg4HpPcIXI4qpEU/2MdO1TNILxDLlHGZw/95nvnIEQBR5
w0xXbnRqXLxAU2D9hyjneqfjTSxrL5y3cyoJYG88OM8h1uNlLMNF4N2YJhmEXqiy
bbaLGdPNH3IpvAZ8AOlygYiOsZpqkBRzY+Sxxzvq1O/laqRB6IRr5vATy6sYfex3
bWmQYQVer2ltsXEcq+rCCu+ubWrUOjNcNplg3cIIswhkay3BRFCJFp1fEpgWoZqO
wLDV+SbnWaY1hIGY2+f/DtylT/GWqFZmIInoOrGwwxor8hWD6wSvkbVlg26rktGt
U2sLxX1vdecBHJX05oCBXS0ijBimxWNnN85rmqeP+lYSTuZQFf1O/MFEQigjEn7z
tUgh+dz9HxY9yqjEr6116jBm64gjXaq0dASvVYIiSocefB8/G5f+/IAKihFfutRY
6Lraws40PKGgg3mjSGuJ3nLp+6nxyxMyg/j/UXlwYq2zG9+holLSJxyJmQ+oV88h
YYnFcaY8toj/7SQ54yg9WTzyF4MX/5fSC9wQn6HbBT3T8ec0fm5fiBI1Sbkf/qtk
Ro2wZjRlFkpibuT118t7AuTo3HH7audjMdd6JFOyC6bLBvjk77TSKQhssZSZRnBR
R8KbD+pw8B0plGNbLuUr+0KLZffpVpbH0kyVTb/71ciLuDmuAgw8Rf3E+oyY1oNd
Mk2ot6Z/tC00amW240JPzvqf58M4h0u/sNklSsQ0ynrPWm878Kwa3uv9BNEdTAGm
10232VxjLT//zmxzmkorv6G7sBhvLFLuCqDvqCeOTwIUxLgp3ymrlXivhsarec4Z
SAuPClah0W0t+MYrxeHV7I+AirtOzwQJF/uMIn+bESQjc41sIi34Q55Udgb4lwru
ovo7BXdKeSnoNGHTL2aa/8n6sgzsO7maqDBIAiIGLuKfMBjAGNMRs2S7az7YLSZi
A3e4zBEu4lo3NlevsP1LEHEuSiwhkMTvDrzbKCaMMjOXZwE8YSWZj2gK6U+eIwlE
A4mr61fhMoEw+niX82GZTtoNYYcO1hhmmwYEGm8vVEPNKrA5ldapnutDiD3S3e8G
APo1ehCUdpNV89dbuDFtYtPYbki9Cdw/xBDoBLYvBIJPwvmMKex9bf5nz654wx0m
WrPMSMtd8B7ebVGtytzVfyWQ/R+jg9K/GlowStNw7CLFMjMIwzMTvpHOlTRUPLSz
IM67hQvWXdqRjbsmUQUkPa66osOCFoYmSOPDb07PlP7IqmWZgcik+Ql5WCl9++V9
74kxT3MZcr+TWx9l2VBSqqFFa3/vE1yQsEd8d4JMdLgqVmc/APlISzkBqzvBtyPQ
iIkkYyzdn6df/ut5P4laIestZSk8EeVrqEhpOAQ0ZgYLPhQ5M3IiiGrNLJtL+Wwh
aESgWjckrXlHXLmRbsk0Pvgo3owViE1+gwOQZLwP01zZHLuyoPdfkoNULW2sRnGN
ekTHUZ2+T4WG4jqYQLq5+eBhPlFAwmE5545TkTeXyjws68mo+YKNUm4xXwS9JgC4
DOC2h9QlnS1WqMSOifRm2I2mj5JH7jomPD1PDdPDtdL5ipKtndD++6zmYTPMsLbs
CIaISXlU8Pb33vjUyQnBoCnfr08E693di8NnBZIMZ43SuDc0AmcJGByznB6n348r
aHMlQuRwJPjeU3EWjfhMzu3/Q6rRUf5OBMTobYk+f/MhGMIGPbuX9/Cu/AYnaoFC
vT3zqwasryJ4oUMQYsOYb8lMKniVaGUI4pNm0/bHRah2P9QZFZaJ4BHLRdfxp+Ry
1/qmz0QkEkCvcZYWIq4nY0Buy5juM7y9LQUtwHDrsM0iWiiuWo784qgeRatixXsP
fRrOp6BW2IETVcf2OdBNw5dmv6lSZbzhhye+c0gRn51+6u/BBWf5GznQY89YR1OL
vKeYAQx+XBWFkONKQqpFfNqk31vRcEEMcBHbZVSe+EHBDRMnQQEFP38zK1+9fTTN
DQwh/f6kTbmQrBeaUv2IL3Vp4DGDS/rVTBso/2wNrpyFJYuUPZgAYuKTlIoYY7ec
kDvAB0awXORNu7TzAm6iBR99K8cAWFQ3Y2gaYgBaZdj4+lMO0zjBK/BpwLbZPlzG
arzgqK92XA3NrFwqdwwbA7NblB8avrL16OMMv2UGIhbS5t+xGhX15IsOKCHtVscJ
2jgKTm45nT1/88k8V9jMNvrMxjpvMmqtQHEeKMqvX5SYPyhXjHXgT5HausBqEyov
Q2c7f5muwOGjv3qC52LkFzCInaW/UdobNq8sx8gBjmvcC9zT0ui63rpZNALnxQYW
2y9ogwoiMwdQq12gCFs/fpUlWdwMWEG4gIO/m7cDSqrFZePcN1F5TIbgXEH3xZw9
MRgoy4ttgWMMLOmPI6FH9J60is5jqrIgGrFh2pr6LXhaGBewCZKSkZywsCA6moN8
92oX9YcqbVE7gLzba9kr7SKyxcbgqM7nj88NQofH0WbklgbgjlUrJ6NWeGEN/yzV
HOyNMyPdSwwyG1+K0TPo4pQXp1YQXwnu5h1zjQ6tXEJcZbi7uCgEXLj2R1FZsPU6
dtmXx/uxsLN4hMGQXh3mrEMMFQx7CEgL2VYIY847GqVyIDHvwTyXcR3EepDoKWMY
BNMK3FwZqBLKBpmONMWgqXbHAETAqdkPSQ1YHGmuMuiOvOSCu59PSG3eCAek1Hvy
T62nyI2EKCs5PM0ywiZO0MFyRpUh6zaXGZNB23n9pTUs7LTAFj2TE1wP7Tj5xiEg
NpKpess7z6Bd227TZrI6Rc1IQdA8dUkUj3jYYWQPqfxgVWojGs7XFKMwTYRPE8M+
7/18DN3T7hSFPv3kxWUVxnoOHSNWYpGmi5w4DldGMkN6SoTIILFj+ZS0c6uBf8hG
BysXkiTfOkWkAzZJQngL5IL7K/u9HBTjUvZihJnYBHgfx/skEPEYXR1Aoo7wRTjW
1hZ+CwCFV+E0UCV6Cv6ereToGKEM5nuBIu4rLvop/3IOn1rE0ZdTEoPvKBhmkVfi
d39al16lqCXyS8M4hKjbOOWZEMjN7GuEW+xudjvDpA91qhzkDIKYbdGR4K+ZGf59
t055uY1hU4FtKYlCsqNWG/YCMpV1uma4x18qJ4t1i8cwsw2VAe4WjwryCbL639gm
3GptupwsOU776XZpGIlC+jAy09zdZFx35k6gupK8onC6EsbJPFIoracJPF6w8D5K
XkNiIraj1affdu4yZpVw8IBH9wLw/fwfsei0BN6IC+MB6SanwCQ7q1NuyYJ0oZ5T
u1QZZYpy9Se5hmgOKvlYB2vU/pNuK03koZkzjmqkT6x69V0nYgSKqHYUBjl6a1DS
yBWJ2Ki+3DwWWGtdJSooYl4eTceYpEi+OTlNV4oX6J030OCOws3I0MWSujhI3+r8
bLP3DXmYEMXfl8K9PpjEzlQn+g8m7A4zXKiBsDOPPEsu3LhgIvc4XlX4+UC/pIvb
PXHtOLMuwngerW9Ct85tTdQzbsf0j08wKcqS9xBHlnyoUA/Imrf246wFZrEOqM9J
Ox2iAYdiSplDYHu9LZ1juHcAKHi/kIUP7M5kInRF8GwzLBdfHUbdueWk8SXblDwS
wYMSYpYGEi/b7inoZ0W7FkPNlFePyui16bUkz1Azk+bYjvzi5WDLzA6JpB1pvtBN
2663nRdrZKwv8Cy9N6CUscAl99iWsO7wIoD7IyxnZ5xE07lAmvKzXFyNCO9aZamS
r5tq1O4liW2xGFkfp5/ZGVoKNuOdUIbvaoKJFTLq8P6no+z6bqjP/Y1Qq/FZH3+T
RXn3By54LjTYZzLIgrpszYU+k7ZfhNFPlt11HgB68oALX8mI28+3OnKYl5x+1+Ie
CUWYrfuRT9TwHQehfv5rXN4nzjB/42UcMfasGGa/zU6gh6j6XX2cRASdrIi1WjWl
DhPvrqgltwlxEuKecVhF9hg9Hy5t/ZMEqT93Ce+SaoerCs2fP9RE8C8V4fky3az2
t2njyMUDsexbNvhuyswthHEVHBTdqPLhHHa2eriXRMr4WVu44ZWLOJu61l6mV1Gu
jxzlWYFN49ZTEBiWrmoTp5uhXbpK3yVIFoQl4wUqMCzlzWjnHVSzaFbZ45ba8v2A
COe0AnssJQZEKH6ovTTbfC3pQL/SNJCaPVXtNdsx/ltCLYNO3trkUi1NMpsGesfG
KgT5ZFl+bnv8XhR+igSxGf+a0mK6egJllh8cRrurUWTBTS78P0COoWDEq6vtuXXA
U1lixYuLmwDMu7H5U3eI3EUzwjoFqjvwZt3m8yH500KlyZfEiZJ7wW1opCuWawZK
cbGbN78tw/5oviKrAu2aGnFC/eT5dA57V6OTa2PLVhBe2IsV3DhpdjQvswbtXFR2
BywR2Q0l6d6vHMBlqITHlx4y0www8nFLBBoay0ZlH8iy044aTnTBFgreLy8mIIkF
AtCj7XDnyxGXAbna9/iXsUR1Ckb4kav29EeJ++UF5EGDMhAayR25fFKauihzzYMa
jr9PpzManInnHTdKVgrAb9WWl8c2We1WAEWaKNK6Imx6nsdIA5rQu6KSeD8lGB1Z
gTYG8zN7FkDxvmAGDnXxfXIxddixQB3TQjgXBbGWxleEKZQCdh8Yq8F/AbVBEKdg
/7cW3ubSRTrcbYoTZ1mdSlLKtWgytjxWKQcGD89lDcp/kwd5hCJXwg9afK0Kfa2I
NpdMNwgOz4nGV/0KwL7z7tDMD0fUivjqBls2IasR/9eVezbJ209weACPCSxn0s5n
IcVaZNaMF0f5nKsc24OZNv3TWS8qJHOg1lwNmZ0jL0WPAiSmF7igtVF7X2Mjy+5+
WzWH3IHF2cGBz8oOnRXovcX0Jwd7eNnBbbrShA8xVhsr+sd0RxemhGiBQnfaEY5g
FxPSpbdQNHf05RijfY5mttyjuaHYM2P/pL7dDA+btq67MTWQK/Vz6lnndLRFMWLZ
9o6DGOxu032ZQrgN5YIA07UO/c5akNQRqCpEm/qxnHaP/WfjOCaPuIIocS5o/JhM
UJmj9yGasVJiYv7DZSI4iA5nKoCEFB+X9uDKMcb09vwrMeF/T7NaXf2hiY6qHPUe
6lJqLVjmjBS4QWV/u1DHiSZ1s2O1OJUONAPTKOUwhjMx/AcwxAO13LRpSxv3EpTE
dhc8kuvY1rTUdbo6J37N2eNVSIRUZEEHHKMh1M5KoWlD4unCjCVAcoeVAENyIJFf
Ewct/8RyrxEj29DLCaJPCNoEfOez54QZ/82b97u0F2YMmrafT+s1F4WDY4tjxX9h
stB7PJKxExiXjCDGMhGTtnGmOCPcrr5+gJ94PllQoVOMwh27lshQy/LiDBX9pVnN
2E8vohAMBIhwvycxjjb2L8ejGKrPMuSchnBmjDCEexhnHlskEZMF7wwTse2CszYn
IVkxsAAbHSVZZ0fVbuBzlsJEtVmJSc4xqq4hz8tsMbSePCHhQHSu68ojQsDqtkju
tPkjv4tuLs1SD5mx40VC2lWAAi8gKuL538sA/WvTh3rG8wm4brSg7pfQCLP0rbfe
nQzxXCqQrYq15pcIJFSefe7T/hemzmLhcu1IKrPSpJ3wJ0CmJ8o2/wPcF8BGmPyg
bKZU/6IITHwpjOdz9PKkIyTVyqwWKd3iX9ndYXtaUe8Jb0dZIAb0BDfXAfylRoDT
idcmLz08iM3tdflbZEgCN0t/cskQLzRdO4QpZBePZn7U07c4hsLksYCzBUTDqjY/
qjYvOWnSgQpBTZEki9amVKRJVyGEdChClSuhuG+w/hOwOz/ewSTKqGDoTbVBOAYo
Zt/zp0ZXb4rHP5xBB5rhNl2ZJ8ROLlDn/X+/MoL0DyBUIar3R0lX9cbnyZb0MWtF
YYwtMVciuXVxV9fRf0LVeCRnL+3CIfGL89in7Gv4U5zFIeFLeV0KUCCgLoFHokfw
x8imdFG+XMQ/R4TRJkZqWLFxN8wvCDhlKLs+C8JzI2pEZ+zTbnXdabvZ1i1VdYM1
Cpk9CmoDBRdjR5ATTvMw7pIRaJyutUK3as9CIC6kePnBTHAEyyoUJnJY/k0BSRKU
iGsz+WqcrTTJlKmMZlWrj4/nSAk+C7CtsS46+VFFjlncK7qdC3Sd85/2PPx/BMns
xw6TZ1n3jtq9SV4IICixk/v66t+APyB/dzv8mJv/cWP/vHjmC19nZ9etNMxKRcVX
LDtxpy9vfUmvGCtYjPldcSPQgfQgISYQwjWGIV6xdMItYlqtrFnEOpKrb/Ly4YdA
QLcWc+HJR1jKCV/n76R18XM3ouN0N7Ge/ySX0tE71VXj2wpb4cr+LkuXnGDQmvzH
7D9fbk9vr33nwcVMiFgCdV9yRGbivGlJ3syAw1d21lNUxRGf0v1GqDynrs47ZQdi
2erxIrNG9VYlFFa//LmOwt4qkVHopG0ZM46mTdnTrvNHzzsksNuy4Uqay6QhQosX
oXajXm38pgD+qd8bwvHH+LtZwFbeAsMjXIvX4NqLjh7NXJkYt1rgklGBgoAfhcZc
yfYZcv4UJsgFS9Hja3Nas74HuJrfGbQQCYO0jVs7kPpKinljKfd2BYWirvt61nLy
HyDXvEBs0FjLWmD2arsk+JdaWtkS34hGBXazxICPxs1hkwLkhVJOeNMdm9x6ZGOw
BpPjB2SvYSZ0vVYBkz9h77yT17rRs/OarYlgG67zs1d1sRfzKXvQUGkz6nGI9h+n
vvvAkbw6/TSlz8csu8qqJZ9L2w9gXu090X9LvIDi8hqC81dEJIBnRhjnud4L8Mvy
ZWFUjAYwWPuuxSJOp3Z17+KNSGxtGGuwjLN3tuMUhwje9yzlj7RsBkOZdOM21s0W
0HsrRIEawrpQSRxRIXEOD+Ce2BHD7OI6X1dYlmNfK/hBauyykL0EP0wqpa09ck15
cVb5lJny1PmSylThB4BpKiH+Kp8A0HmRUNyFgCI9yb6OSYzB8KzojFNE68dC9T4N
Xm54IKHrOLJjBqioCUv5KWN/U0YH3F4yxnVtYJvzc6ZlVP1fre9vw0gMrgXPDoM3
iYs9ieLcCoqAqqrjQ1Ipt8i5l51fRCbwnGK9DOWJJJX2nWcdHGQp1gqCLD+clF4I
B+dosu2ZUYezXnjzmlX81TRJiFrw0xvamxIjcD3TzAABFEYySgZr7e92lHV4OsJ/
Z6g2rBeMoQ2cJoNlX4T4NPPgTuuB7R14AieQiIerDsM5lA2wpTp+MNrLetXU0WKH
nGVPeWJiIUJ8W6R9hBDWE9DS/DF9NYJUHnKkN/OTJ+bSqUhRW7EkGvmSQUnCo8Hb
i1UVVsDZozd5Tv7WuawPhkJyxdjEsEkpHZE5A8ZdZ+3ybKhM3Uw6tKRYjuL8nbmM
VUrQqLgy+08/cTpDdOq9nu3zuwj7/H0pzqu4Sj8mJJKl55fpUS8x0jN6o0eT8ohJ
a+1xwSvdnsT/4I1FY4dhEoj9TIJKV74i7sV9hRydTSDq6rpgkyJ72XIHpkkiXLRm
j61we5WWsDSL9Bxd+2hA6wGQ3KDUIbUZFbRDQjxlJ0o4Wm+mT5oEj5jJzA2OWyv7
AyoTFetH6VgQ1ZPEHBT37xUUt5JuToM/PJORLEhfFgnYfHqXiavWbTL63GW7TEt+
dutMJG4QRFLTQ/P+hvRHxRk1Fwl+zlETVOWfQ6CY8xwgP+m4VlHDLO9oTGBha/pK
qBHHaRdb5QnovkqTB4gZzMC/JoQOLngZOppD1El3CONYwu0hgnOTOp7OtJuS/TKa
aNQnNEJITp0Uic6E3XFQ9ly369J+c6ES7+yyAHvGx+G82nzPhOlpgzY58PsA3+fR
NHMaYR5e6q6RJR0bCUPl0Me992NAq+mWXB/zPPTYEUCqPtRz/WVmUNztfnqpTb9q
KlC0PP25GpNGbO82uhgc6eZvhPZ+ikch0333GqV2t0BTmM39xg8MyEmBOW2U72f0
S4wpHZNuTBkSIFheFF5c3PiESg0vtpZdY6EK2jIO7kScZz6VeUwpUyqQRqJ0/Lwt
GRHNR6cicKo621if8eNyrZ00+oYVOwRXlwowmkUU8ZDnZa3iyYudo2VCrNXTYahU
eyQNOnejV/llbvL9uJjceiNPslX756wTTSoqWPYiqHUZpZTBnBH4/agW/nkcUx0d
7sh4isg1YCIzZ1F29etOVhKuQ6XUasTZ0JFlgUbARNdMcB4B3/qjeo094dLdJesp
QxCEL07E4t5xC8444jYTQ3y2z13c2paYH4wfIpkYgimt3RdfyFTJABJfkbFWbsMZ
L738PLEGxlKOCb8h2CIfMHHN5LHeibY4zF7G9B817TRcOPEbiAip+G/z927hn8VN
TJyCJFkjkvta7fSYlWhfpAIPZixzLktlMR7lP1D4EzwWt90Hz/N6XnqxbhD8VF9K
KA1TFYNSmCrMJN+kyDR6c7yqZIdeRngglqbQquinawQgeEftEjCJSwQ6N77Mhnxa
eQbPQFcLHWh9ZebWSIfjc6eSQLSi/+l1/lsRECsHJqxx0lV5YB51k3NlZPILJh2H
rMAlpbBiB1Py47rki77aSL6Ddt6FDoIeBiEAj0yggthMcejjwEVT++DnqUMQkB+k
9lF9K0ahvnhoJQwRkvIegDfJifqXLxCa83ov4eOF6ExReMQkJv9EcEg6Ba4YSEYd
HM+qcGT9TjaIz7e0MDmw+v1dw9ek4mT9njhtlQthF0LDT0zqEdU4+OnT/Z59zCOc
+alXICHaM6A1WlksE5HJvTYP52aoWZZZ7RkIDiiiS8VE3Qrb+zGfM1xzEy2TVxkp
7099JfpB2sd9/j/vM2S7le7BTGyOa6wT++KQWxKjE1ktT+Ts8986Es3SSsALL7fJ
XnxEEn6VISm2Pt6ieG7jlignoEhvo+MmJOAzrqxrNuvhbBkqiBChZm6zpxqZ5dmf
us2dRDv/KCWLYjEkJl60VZMOlmgMfgGBae9Dl0qR50uQ42ScGP1fUp2gyVGVGCKQ
PufB3gVXFjl2Guf/Xq9L9HL1ZcElco71CbS6y7+1LWaom0B136M550W2NXITmxvo
w1PUPkYPt8HxI573FjlgHklaDwAz+0TR3PdBJes90bD4mLv2qHHmziSkcmLMIhDu
CAMT2kyvZgpkdfQFl4K3vyDesmhPvYbzpGpCy3+p93pqi3urzLzylLq/J5KxTcWl
zLn7uQRMV0p57uuJkJdE7tR2Jkyvn3N/m9VYMpmP1hMrax9Fbu7TR9xOMAn+wcM0
dSUHhFEeFig/ql5VlBc5E3J/wxMQyCw/5Arw+ce2V1Txli/j6NMcxNREQUaH+QWa
C+fkbo/e/IDcas4sI2O8SOqiENv5zEuQ4JVfDEDsaexcrPqYMvaw0gFepHnIlsjn
xsW95EFrAkjEi5zlMJTcnk9P21V72WO2/ev8Xn8SURq8hTYNxcNvpXsupZEo2iNo
4Gmdb83wlsSOOSdC+hGIXoQfR3ZvLBt791xtK32J2XJuTzufzEgr1vxE+W/lOSBX
nxpKI2PAxtNyX5kDAUqkolmrit9i7bWIm87SHs3ikyNyGYiCzMWnGjRqPPMymFvU
XwIMPLSf8E5bjyhpLEhQhizP914NLnm4iQdzV6M8++6Rh0eBBoK7HorJFBnilRr9
J+Or2CyFDmEAUG0BlaBQOAvJ7/YJgvOchc41CP8oQHnFnCYlAneO2jGNSFCQlYwp
OyHqIKu//776W/Fa+o2GgMENWSFZriEwrH9sN62m4oCkCI5c3drSSiye+FQjGdOX
03H2lF5KOvIunWtQBK9ynxkTMcivO6dTuX5LsWd3gV5HByJbIRqHw+aZbwQ1EPiI
BhAYYaI3jZq4I8sXtcDpeO5v3f46m9kDPqVh2ZgsPFvXdVUIKB7eXYjEL+rDZGPh
xZSJJv/kOa3dwh9bXXJ6V7bJqwXizjF3sk2vVa6DofzIwYCuOOxOjRU/gcoko3bn
FKF3CFyrAAatKEu+4HctVQ62Y3Kv2JnrnTq55KuQmCze4f+L5tBg/fIdNzPfP97g
I9pSw18kVHwYitsLTHPIifOOSJvFZ+d2L4pmoD1deR7PqQubE1uK44NDD1WiDbGh
m/P48MtBevM3h250xPCeS/vY6GggZdr6ysOSo2c66Fnm9HYsdlOqKFw3/9606Lw/
AYv7Qjgf5MevDS7JHjywGjfAOUEkPsgERmOZ6MikXhI7FizAiEj/YU5W/2B+cOKI
47N6cbXXdbMLMadlSiEFx9shJBEhosyCg+1PNBjieGG9ivwF+ZVzPrNtg9HiPj7X
Td2DeaStVomSktAPB2F7PL72pESpienrP04gfUiuc1pAWzceft3FVOw7YFN6BLH9
ewlQnF+XyQFFv9TS/6CT5aqlhEx9KkAImikkkJdVBLzhc0cYjDH53a1UjjnIZYmN
dS/VY/RQfn0bc5fw4VGjSoMgjmfhUQ5BW2/mAgeO0wq2PcA8NKNAaMueIdmywiLx
10HWw0hhek97udh0GPrYCm0n3ZwTHYGlycYQkoWzgYK7BVYOedNgb90i/Lo6kzJQ
s/kSy5wlNZxx6E5h28YKJsq8wrexBETK8/viaMIGhhKSWqbmvdg6BDvP1bEYe4HI
TXK7X30nsM6s80dp3jm0j2d1/z1CX5pQrHG5OI5li1biFNXeuqARqwAj1ggJw4lm
gYHNArCSex+lr0favZZMRn+dt/9kVmJH0LkGowxUJQKdehRmwNLM5V07HtOdvAc4
K1pxZL1uHSI2oOE5oUNu6vRWfa9Ll7crqXwPfiHrCwzU5YIcOAk4QfaOyWYskp7U
OzFqVvoVI8KDjWRYI8uUA6alSMD9uKz1tV1VdhJMdwM7Y403M9E9gwiJr/MyhKJJ
08OD+/9t5K5Q5kQrRxkEGtqjgdLO6UnFceO9nLV/xQei4/C6bzwRgRN02TJ8W+hP
PAj9ukB7NZhEB5Vi3Oi6AiT6B4VmBr8YrsTs+4QV4jpD1CvCvikL2CYfixo6J1R2
N9AJVi/u6ojljO6LWJtoOxbnfLcLsJhKW8LXenh2FtyqmRrC/Xkz88KpKZuBVTSt
bB6HMqCVsAQWcsLX1R3+WXvWi9y5ngB2F9Na4RszPz4kFGtu+XsfjGWhGN/VVI6r
+mVxoBj5sKIQAQkyUlKV7C13OCFGs6dSjjt+r/HlCqJIJFbboXb/GA5iU0R88EPj
WMpoI6L9w+uhnlnGx8/7Fk/oEgTIA/Z2S3t2akNw0QGXJXpkoIaYQgEM16J5BFwB
+5v3D7ZFarjcPZLwikLgWXpEsWuox1kiSMxeOOiSyO86DYitRvVoE/145MEFL+qG
R1vzNjUYKHDhFrHv0lN7TrQk4QAgi2z+M6wkiv4T1LUTn3+ab/KhA7WAOL61fU53
Sd82N8KV0BL0hbbXNbF82IpE2uLSC46OAenAJI5vdGaM8cMnXcm916gR+tY48heN
6EzTDx6PyPYk8qydt9m7v4KwzHr3SwYq+E1i7H6erCYH7U9OJVJ/z+JijapOyeP2
z4hCERf84SUaZHiQA2d0EJ079dMrz/wiVgZsV4gpBMP4mSavUfExxMPDkviyGXGP
tQrL+AZWM8gCANfMLOD/6Or3xCUqM2f5iVT6CAxrcaRNvYRHiOgT7ZGAwg/10kxZ
E3Zmvwv8XL7e1/9UshSJI125lpZ8ZMgxLWh7dOPM4Lry79hTPv9vHt8ygRIDVN1T
QMJ8siU03aqrMHxu+Mvded7Hv81gOxNuwXS/b2DoL4eko9D2U7gKjEdnp6B3xUyS
e8ZWenqZjzxPFdgEsT5LZqE9YXdghNwgbAaAlD3APBYKqTR6K7FK2fjcAK0FbeTu
Ggy+xfTbdZwbFjnd417IJjgdqQlxvKw3B6V78D1eqZgHsqYtLNZLS2jhmWiFA4C7
nTzkF2VELHj9mD3bZsUzzCY0NpU9zAfNjN66fk27Ro1Kau+H9QuvtGg1wxuNYnVa
tV18BUBt9K/XHrKcDS7Ls97nJUGOvTFQSvPuTqo2yQP1f6H3MHlbaMBbzTfGj/uP
mOr0vWdYQEGqXBfENaB31JCfyb/v7SAt3HFphNeiJDlyefKqGi88rDYSlvgAg6bo
OutdBh0RpbmsO9yh93FKVlvju6PdwQCnSBNvy2NEUEcIesPutPvekAIewWNr2YrL
GF0AQYBaClVJmYrdY2lPzR+/mA6565tz8003GSSb+CpWtrNwMK10xea3eafHVmGJ
wkRy1UELTrW0EMaYs41lPeaBHGF8gqOGN40MOdXS2T7V2VJuVZQiPYMdxK792y2U
U9me48hKmvFTHX+YUCKoQPQmNGJJm4NB4A+tf4fAjpEcPFLBAqA168WPGwdbLCm3
5HToV7vJu4W7rhBs/EB8hRcVAVv1430VuQcZuYcJPO5Ebi8r7wuZj6MVrOPl0MQG
POnbISHikeOsvhmxD2XTXwxhgTv85q5elHFrwZNM8BzEABKiZTnt61EF/hzAvKcy
aM2fu46wkXjwAuCgQYjVzM/oFO9t4aLMoqR9FFvPcZsLLqv+w6BZIc1wq6v+4GO9
TdSBbC/h7/NwDadFGYf3Ftc0ki1qL37DG/hfn2Yz/vnt8eppEk6ndcjcp0YT28Vk
LgDaqm5k0zJ9eyxGUFtvzYjE+YFSssp0tZZLNUNOp5AOh6vNvZdcXthQxFziKrw5
mozGtoOskznE+KbD2k+eNuZh6Ojpshk9awl8VV5lhhGkxwMUObOvvhpR79KjVEnw
/jxa8PufzgFzRy91mTkpr0gkeHEiNfYATetfa1qc12WDMLEcWrDCJCDMW8raEjpg
gbzWapQBvI9t/7we+auLwdwJY2ogv5i+Hk3qZNxcA71gmTCnT07lDNLW9KBTfE6j
LWBCPm3LN/9HwVCuNVpTH/cUDdMHfnPrTVGmN5LTmtKIZH6USWZeXzqBs/2rtVMB
RgSN0n1wrXy/iKPjIIL4p3e1SbPHhG7sDYfIl9mWP46dfwyYjdFval02kOjiUaWh
RXLJD3HaxhCF04mr9qxRYQ2bb5Gg/yvvdNqiZAP/cZYkbpBo8kISrYKFdv19twDy
A+w85+YNIYJoMtuJVoA9BCjP4eHG70tnPSQxpHIFpOARMWJsFluP+xcqqDNcFQ7q
SMXbmpJfAaWbhG2ra63eC/af+cBjDRTumkfLHM+oTkNnzSnZriyLpnH/92S9ROO0
/HgXfh5WwJetheXJ2kuofHhqra2FHePEjsjNVYUhZ6yrrE4IdVqs39M31Ne4krx3
g0MbDiXSRQC17rLpwD9OMHuL3dCXEKQrqdSQ+u+1qJRjAv89tl6YPb6JI4Unzv2p
hAh2Cs5OH5k/5LTEO2RoIPeysyyuuX9/Tgi/gc/f6eSrXiXpNEWfvBPeg+rQmgmE
NzrDCNhR6XUw6AZMiW+t1BYAFQqnYZIZbDfr9pXE59BtFY1mpftUHlGKPs+7ecRr
a8ha3NsyIecOhEYQbHNNRZPFPumgS/rkuYLOvSU1AFzjxyoEGEwZ+Y5bwZ9G4EAy
NfGM7GdEMuH4y6fYMoaTipDk9oPWEEbmlLhguFMMq2yoLhACdwmt4L93pDnr7I8Q
llF9dMMeR+7r6ATfi/hTQc21nkKxpEAbNflm8+srFqNpD967chmPc9hMK/g+rS63
fkZVUB74SfNxTztPP7BI2yPHuhA93y3QbAEQsKo/L6xVCg44tVogWJeKllNZ0zpM
ex89lruiPaheMRV1g4EVYGgYqKsXgs39xOx1rUTTYzQNAAJc0szeFgGJs44+XgQF
5RKXriwnDzW5UrkqdihHJzU7hZWwINP90yQYror9kFA+ach1958xR61j5DIt5HXH
NU/LszbN7mMWmx8fEUrFsMvuxOVG7Be3Lv6Zth1fF3ds8cYpGP7Hq9pwJ+EUni5M
teLP94aA8rkRVoHx2uEMyT6GBa0Xl8rF5I99ohjoL1y+eI488L999SfiQkjds7/A
NCgcsROX6TFFXzRwowW9+2w9sQF0gICVkuT5XFq1JtrQDSEKZ/eWCIZI0PHZEVBt
WwXjy5XNOOBtSVCZVRfjoeLpNsW2LcbLYdV3JNHGNrExb0CE7L++MO5V9ZSizhYI
Ncb38MbSnjCJLqLPjbJOheS14Ng9H7kQHHjCnBJ+nKC8AXTbjdQw+kU94fNtuBzi
sGY30/NHdSlkf6CulmYa3/hP2zg5g6PqODMPI8DYaiQJLyn2x8pmOpAqOwfXWhWT
sPHv6kwZSOqXRIg0ZvOTEd5x6GhYrw48N2sn/hilJMLEvZmU423QfIEM7DPf/rVF
nm6q6r05h2tbW3c4UcjssyyhSvKW2RLoyiQORk4TUv7rFqbH4rqUZXn26z3bMKeO
mLPimVVf7KSltLkhAMtfbmKmyEfuD3+EUo/G/s45yW90gWQOApZm4nJWyDaF98F5
lGf7PdNwRpBW4MKTg7Xp11ZjeOw42mxnBtEguvU/5YqqSwzS24fWEkGwVANAkudK
PsQJ0Mnfy7dTiW0AkPBfWbZEgpPJslm/j3x1Te8zX3i8DJYh8T4Er3Sp6XGwCptp
DYfDWtJVinFI5CeeyZHl8T6IAHCWUCVZ1R0jdh25ZrYLjqrYsOFTmsUxA3MgXEG8
CHVgXRgvuunbmQU351NiK1+V9yG6pqo+9DcxnwY0ogVvEVhVofewrjIWPqjdqVRC
+97BgX7sDn2FAvyLItNtDqmoluD9hkRHb9SOPbpFXifNCmQ/HeLneHDXIy971o8O
X7jsgUuCoLOwXVqFUZ/693Mq26YFOEpo+vS5W52WYQOlg3YyYmkm3iXvT0LhnKAY
L3zAnXBr4mRN2lXK7VhMvIedYH0QV3EiT6ooMsDYcyHjUj0kV6e6MB+9p78ax1dD
QURsuquwt+mnrDAcnjKdFoI54IUXQa3g+f2iPpuXXtPNqBY7tZMaK2yuPJ7b2Gb3
onsS9v+k8R/XNITlZWrkzc12BQBuf0GTG3CpTBKfLdXmXMmX5+wV6oO8MzepkpKA
fScTy3cmD38vA2iWOmmScuJ1Oixme0Gg61+ttEahXjlg+rx/ZijuJUXOkCkefNBM
hrIEmYiaf/OgnFNLTqokWxJp6rGg9Wu0X1lmoCk1zsIyIvhLlGRrDVkgVGfDtvNK
DAIQaIviAAokdTguGFKkqe7Zm/YExluU3WDmPlKnl5LWsoef786y9ARf9851fbWU
tfC3oAwGFvBrZbKez7SXS03n3frv60/TnES+zTTx3DDBqLrgCsZTXTUH8slULdB7
xWVjQ9m8xncD6mO4WlMd5ic/35z37h/lcH9uzkO7PNit/32yGqQL3qgVOIOoOgcK
CS2aFqjlF2vx31oE25KLapmzdeMxWjDpoypUS5wHgVB+6tZYKG6V3EDN6nTQgFow
DBJrZ+WG9/dvp2uWYJUfbXVpyl3/uuOvG/aLLQiT02UsOjEI+fsb5lCJaUpF79+1
jr213mG4miECwinrCCxKz1pbssy3FvVeY6MjAzB9XtKwm90ppg8c2j25IKddg+As
7eS+n0Zx25bepN/cUXR0TvKOsfJZ/Tb+DWw5Yn58flX6DycOG8CP6ai80nBO2mQD
fHiiEJy8zvK1oP1Eku1HarxR9Q4hKYkViwf9aUYrU9pXDYHzA/QcEpMNnf1EDvyU
Ybft0Ka8qsNroV7DlhlYI8Ag0YCw3rGM2YcqRD2nTteaouZqpJGuGc84DA+gyeQc
LpjGnyke9dVLpcFaNyiPT8VspSs+bj6CWcWPzFWCAeliUzPIRU1bXH55CuSAoUKZ
C7P2a/o5Pqj0Q2PJGjJcwuifPDdCTvjPRy7Bu4qZFJsAQ7UAW1suAiq99oZSLkTU
5gTgTnH8THV2GvIlu7fn/hVQinNU2eG6+Ft5TKUXj1cJv+Ml/Ah2RV8A8CSBBOMa
n+wOIdjmlyEOMLixMacI5ugvaO0vFWlATQsX3znSsbAKXfo5CnoDhCYHT56pYeXP
Xxq6I+sjIjhvog9Z1kkpdV533DSLOEVlhZFFec3Ttd0K0BGfh7w484hJ2HG8y4fe
G5Pcd6tkTsqymTkZXyr9J0Oojd90jMNx0v2ofvUU7OiEARMxMYaqkGEKBooTF8pZ
/eT4hNFidpfdlGZhM8dUKL1guEGTVCgoAbQU+fKZzkV5OjU85XBZ2NpW+tWALxbV
lVoaD1X09bUdV8aHqv06pTSgeMpbG2yYlpezd8D+BIuJ+7hPb+wvPVHeK5DdEDqs
j4P18fnjEHvFTjM/htr6isCJdbkWnwzaUlvP9qB2SDWiw5cZctakGAr/2Pn7xl1U
hB0PFH0Qx2/ouS2xA1WWuKdB2RRLMTVQwSIB9cGOygZo6+yIbhctFXVan6CDZDDR
UV5ud14KXyG9SDvpPAllHOUnHMHGBYOOf1p6ujyL2QnSXD8e9UinY9FUSEilQ9/6
pZsKDG4t3ivjSvllayrv/CWlKBOqyoGRlVT95V1nacrfw5tUfKeZO2M1ZVskH16N
zR1KSK87nQ9COU82ZyptNilJDR6BI2bKLV6GaLGFAj3Sa9S03xFZYriz+YR/AoVm
rcqkqb2Dsp/XriyGV2hgeowpJZ8wS185RWz5zfwb4kbulK9bJKXeX41vRrXecXcH
nkJfYb2wLIbJT+71jDAWKgXAMUvBhzHEXnU/ruFJ8BjTmfw2Rt7ryaNmco+iQXS1
MNw7UZXudh2VX5eteMf1jPp6OJkTDpAKZq5zVgeYYyXEAk5m5UdP5OMiXdgl32e3
rTFhdlxN1avyMB37R7KeTnnHc5jRWHyZtDFKEQKUcSf5GreAIMM8KcZo642KgwvR
Naw/9VeU3Myu/fPMFePI7kln/Y7QhApfq5idoDpCCNVyO2dmeg4939drkfilw5F4
AiLM3rJtJDQQvKCw8/XICJzttggDydQGK1i6TYUnh40VxOZEuxxCaXkMvH9MrhSY
SuB+ry48bAy+IFS3edp3PR7Z6mWxy+LUwgsYhTyaWyUg112e3VvXioHV68y4WIIz
ZklBMYZ7uPOR2AKC8A027VpJunOG9DCc5Vw8Uj7qCPnMj+/qGPho6Gevz3SqIR8k
7DFuxRrch4un0FcZ8ZxK5pROkyTkbBXmbC35PpSE8kD39ROkFlVXuNTrbbILGq1r
UofETkI6t3RPQ4RbaQ8zItliGY/JsqhMqCJ8KlH/+c13EbnCfDhD7sKZ54Nua7bC
G78s5HAkXdJHToWW/LbNzRbXrtkd9DjJ3RI90hA0dEJdsLt4Dm8a+LIPNeHB60h/
4/d5hIDw7YM3QAC5nAebbdFF6knw7ywR8YoBDZlTfgR0g0e56M6iWlzOgZ16Dp1A
Be8o6+qyMp9+U1FlskInX4LRgg/mQAlVvn0bqGbgCj4yp+0byQGpoH7NjBTRoQHW
Z9Z2vEGWXZXaiRHIX11izbpgE3jzHgm2/uj9/6KYSgnnJXwHHKKkXMlRU643RBt9
EdA1O3XEdHCOOkQQF1AXgNlFygVedM1pIS1MXlc9r7hqm3fHxXONIn3rYXzBxO3U
viOtNEJG7KshbCbvuRVh2Fw5uzww+KOxXw+nuA3rIO/pIxLXqKHNNUsvt1D8nEMD
llRV4088KRj78Qm0LPS9dl60zV4VDFdIgKFnRr7WK3g265qKoUxvFRyNgoJzvSDR
rRo8dh3hd199mLhTc03bAFKiMjyC71wU2bzNGvZfy6EuIpT/0v5+l6O9gpxZod84
lvBkSWvJWDSkwbEyZN4/olJCZuNCOEBL6VaERdmBQirtwbm7HHHDbfXGdPFeAezm
gYy+8ymAV3CnwU6OGT6bS76yqYI0tCdE9xTX6GMlb4DXHpJuY/+DXKs5yKy2TIRZ
19t6d2SFVavym1XKQCJX9bD2aafRH2zJtb1h0TDLHiUTKA/BcEzrQZEqTvlHZ0uh
x5IdZXfrSFs9Jars1d3xrQfSUxij3DD+sGWJdWvqs0Yt1z9ISkMhy+LCQjGM2Ao8
Xcz65I+MPne/tjLPgDsH5AUcW1gG+yk+Bgi5+GT+i16cUuBE5GeNzfUribvrT6RU
tlblATuaxIobvhyprXFhqDZl8mi4o1lim1ixKAagZkcDcb3GNAgkIPN/SWgBjuXS
DJ4EpcoTZ727T84+2tO1uVCVPRswoyOyAWNNCiZ9Y9QzjEDu2r9unyvO9P95b7y9
Ml6h7amlOEQ5/UOT+XP/iFx+RDpVhRonMfne//qYRxJLbGAcDJrb1SwKwZRuK9SZ
bEPOXWCTYKRqGFgQKE1XS+Tzs15IOJ1QNkjeG9ofvuXgk1OjFyDAGAx2K+e0ugIe
sjFdYItWpq8x2CTdcQTckKh+fwW7GEE4f7QLezFkJy+EfUglfPLLyNOSTOIsls48
icmHpXwxQMkE4TPqPFCrIp9P/Ll0blaN4tPfs0RTQao7Ye3m8MtIQ5Cn3RfIM1Jc
1Vbaq5vO6NkjnLQ83inx++7Oiu3HJYV/1EkvlUWch2rE8pHOzI//t5NYoACWQXNI
RcaBJkoH7F4b2JQT7aHjRiDD/uGcRTLyXcRIb9QtBybeoOhg9BcVSGwpCvqWW53v
In9S9zhF+ek4O5xVN+h/ahOvohjeuBmyco3Rq7y74vniwo8ZBLANKrrCfAKVN6H3
RtH85IRBU6sR3KbIKTXm6chCP8TaLq71EGONIvYvwlnlzbeL6+jDbPPtOzihBxK5
yXpi8YKyNsV1YDvPzxWC9s67LXLD3GocsIzLZhkroZXkWgPPPmTJWHoW6MuEmYDl
tEZ5YKueWtizPYY9EP3n5BFPaggmdT3tSVgSnPK8kiG8huutH1ynv2eIw9n5zKmB
7CMT4UTg3CPSsh5/4nqeJo4NLWgXaNyCZAozBmD4LG5zYRWeIbfJYCW2McWlE9RP
KfEMsvFyKyxTzNvCODYSIDSRbh4W5cmhbqnDaQzDmpryVe6+d3uki5Mu5lr8lhqs
V6EHZCthRgunjAMLz3rmwcrGOfmwtB32IWX1ovss+56cSvwqhnKrXyBxnUFxCCOF
WEmq0dv5wkIaTdm3yx3VotgQrghpF2gRoJjPp5UKv4nxU6YHYJIVwsgM35aVb2CX
eHuvma6on4C35mkWRO/NtQgCwEAWAL1FsDfux0AzNL2s6nhO/qFSD1GNHTJHe9lg
ID2iqL1e51ibiEwA9HeS8qlYtxBRes3C2BvJXIpoyMQdmmvq1oelsv1gBKIYtZLO
vGGhRvZFmnxEkZ67f3z2L34XtgUxYsC5OCS+YMZBB92SPXZQcXNG/jXupgy7aAtC
BygkNBQzPAV9b7KYaO9k9+OJcxS+kHrCaQ2gMmBPWhjCP5hPz7FYrwF1zx9h/xJL
xnbLgBlKFYkJmWYeFX60v0m8ttbbwnKPQHOgAhMrKSXDShx8Z641XG+zTvWBYlch
f3bvyON6dLeaTBf2mIgDK44f9zOxSUdNQ7IsjN2SuY8p36jIqMQ5J2QIgPoai/rX
BsRj8PVZgbiwbdpy1nBV9rQic92jzU3/FMmJ7x6PDP4jubJavcC8HBUtrgTNa05y
DFyEcS8xaFr7nZ23MXIvBBznHULzLfOh9adg0TDyLrQ7wvaHOz4v3OFigwrpa5Rv
OcX3WhqC5/R2YJrjDmFveJaawbADtUh744yPaTck3Q8pic66tYxO9jKN/xEaFnQP
w+Ud5P/+AM4zBKXROwfJl/xyBtntTqsMn/vBEw3a9RzhSirHWbShMjZQ09U4ezFr
GuaL3QSYr/d+IMQIcvXsK6dgPH7tzXiTfs0RPy3TuDl3rZOHISA+PtXwDlZNRAec
IFkZqDt/QdUT2pC4I8eH0pHgS417ptEApfalq66l9QzJluV2lmhKIgIBwXN538le
EIGH3k4mV/9YHairOeP99aVyIiJF/CXHAGMvGRqaXjUYyPxuWcnpKiNijhy2D8ZD
jAJlJaoOqgY8XLnEnpXznUL6z7I7RM2fWiydI8WJeUdmNB5d46bsTaKIPePJ5dci
J41nCs5upY+gOYR18Q6sm6wFYrZlpezf9lEF79A7vguZVkcUvYTIHb3qFL3d2/nH
FOkGVKwuuY/Ain41KXwcXiv5kgrztRuJqnmWBOSIWOcHThYWk3krkGUsIyv/ZdOu
WkvsOp+7vVMHhehEjBv0mROBW4E+KTZW/7fafJtrouf+Cn0b7sqgNdpos+tplCHS
L0+/7J+bYu8qwfVApkuUtakcQ9BqklqRhx/PphUzHSGlTtq94Mi8XxHzs7Ws9vLB
eC642inpWrSiBTBuaYNczmOC3OntkNRSoZy3Nn3twvjMGr3a7+YxnrZHRJUs5jmo
oN+66ktLHQciKdKr8PKPkOgRd3hIoWj6wZy24NGdOpXPd44n1L69DWtRlLlvekLU
9YtxrR+1yP8OydQnAG7DsFYcOtpLZBfS3hL5SEC+625dWrROrHp1XO52wgXK7Nas
KTycBQdkRyU1d+5bx+PIPjQFAZjaUM6iRJkNHgDBAnyc/NiLgA2emBfFRLlysdFu
74brdtM2hhmVLcjYY/Y7ngp5KUWixvMBQdNyslEAndPlRV+Wc0uaKdv2h5RSCNFN
FCwRAb9fJ2Pn9vTzcB6Qd1kWzmXgtTW5CCT9p1tVUBKupt8+2UhxhAtxuRUhEvY8
N+Ks+2SIPK9lWR0kh8ceHzNTh+TnhihXiZ2Keo4j8VnTMdHAgPfd/p7M8a/Rpfww
4WcGn7YZQ20od1Ck+D9AKbWa24quZlx/AxrQkGuK85cyaPGxuike9pcqLPZzU+8U
KTCOxfC6gPcIJN8dDyDiuZHN875gKWR3qp1RESOiLwd7ZKw1uLS5KwxBEGB2qVtd
jZIoYcfTnTLVP5HHbf0GCu2cwVjTp7nJYBhTioPmiQs2aQbpzkgIv2Ir46YaPZZ2
nhWuILMt8y06J/dkaQ2kcGMKeOxZF+GC5Ft4bTM1GVqrsGDd6/Jd7WSfZTpA/5uq
RPVYOVqf2Gb4czk5C23dJqqvnlBDrODXInNzIxPLZcq4HhsDHrN3et3ti7NfWCaQ
iXyZaHo1NV9Zq4vfMl6ujs7d53quuYUNXyr+xWKoj9yRs6n+QqW/UQy8ZmgDmPsH
iKwao09RSUAH/6SRsNHba5i8mU4R/P8Mo7VO4Jc0uxBYSp6AMFnwQ+27sYCUjZ9Z
3FI9PgjYzwnhRovAzeG/T0zaM9hwh5Litmn15/kyl9mh6x+7JOgc7OVNsHgGb+GU
Mn8MgafaBrnQ7lG0dBppeK7D+6D4f9tTLNvpWeTRT5eBYKCsPXEZ3Jp3Xpb2G8/4
0KlzXKZgSNoScYJm/+1KfaFwShUmB+fOH7BEgzXAFQ+419WQRNByXCRBr05qZydn
SLDNZ8jqyR0qbDZsgKW4Uwh3FK84VKNjbvaczxqp8EMV9giRClZs8ViZxRYTOksH
TBPYqXk5g1qbl/+VkgMilnvoh7CCx11bXn+Fad8VgNv7QE3930MtaW+ACDrXqllf
Y+oXsaCvJdlip6iQL6glALg/anATZuFsfrhkziTq4t7ydjdlHduKGT62QOjXkvZL
a0IjavsVBv43m3iEhGb0CObgRVEDKwLLiHXQv/ndtcxdaqSbjRqXRtNlP67XG0O8
ZnVa2L+mjSJqzqVNoGZ/yyO1/1cXznV1nTrv98IDUHRilbVNlK8GbsWo50UNs8T4
PlW4fIcb4W5NPEWrt79A6uchVAJ40bpinlTWeVZMl0UZXFvPZkd+xmKYuCAM0uKI
WFRsH2NI4Cig12wbWPAL1fWO+jzp+DN5LMjGl3O5GN06AmY3oKLPzDcJ4SDhE8LF
wyb9zHrYN6OvDZ8ItDc0tOvzj7CU9NRbrhBF3UU2TXFfO2vJxPTABkLJMzl+Vybp
odVtEv2TKBxIi/mvpdrv48RcSHe5u/JPy8JrLgxOOEMPaDJt8wVmZOEqAuLzehzr
Rt6W0miduWhFDOaoWpDH8tt/P5FWa7oGqO6U35fNXy5V3YI8ktGRMf2rVWJzFuWY
Q+tEWM7bjzFGdQQ/ZEftEH42MSSPGSJJ2zKiZiIde4VZfjxo1PpsSvvmPfD9tAcf
XV4YDOIh7Rm48cE3knt+ckVAwKtHwWGtMslqP84NVlMwxkJMnp2IZjS1Rq+soBsq
G/nLt5H9BtrtNYZN9oETP3J7WUNK1YrEqYhxDW5jFU3s49KilpLRp5TK0uXLXoFt
C5GnwTcNf8xhwCSbxU04G4PGQeA+9DnCfHHEimxfaRda/gVvIl6qq6EPp3kdKcju
vDse/NPQEei2s8dtyGDQE6hsU5rqsAjrN5XyZ+J7CYcH8kWT/jwMWKJZVUL4ec5X
AvJOrpwnEfnXfUIxGOkg/7MqnoH7Tz4hGxIZip0q5YpwcLoqgs1JXeWQ6DN+bcVJ
EAGIAUs2fJt6xPRN+WPCu+m1jaWVlO0v0/jBrmMalPBkER6P9ve4prKb7P7OZ6tV
2s0wZc3IYVpgNvZolMXCePwKO31ctnqTQVNbeSpcnFWZxcHEEw67RWN1AeSvm0VV
jtMdLB9ymd6j+me3oWdnqbvjPPArMJGJDMvZ0um+i/V7/VZCXjz0vgNqQ/5hmvnY
0+fGboSMU3FV4wAjxDTr0BQF+z9t3z4bR0PAvCjbI51dc+bmDQl/ekX3eFzuNr+T
7Xo0UhTdprMJNDbUjB8dm8rG/avYorkDCFIwlosnKRXnBTh4HJ8frdhrXXpkcDDD
Az0p4qxJL1/0JW4+uYYYoZ06H9BGatzjsfTepz6m7v9u2cdZ1XkI1dWW/Av+L6Z1
Of3oIm2NoxM41xhnRU47e3b1bOwzu/A37VmM5XYtX2CGeWddnvQABpfNh5hEloUI
/PPaLEm0cTsAWg0AfFbruu8TRqg5pXhszNnYcSk/Nz+fwYvG5ix2ESKoL91IfkD9
DPg4kNIHn+fvGnzhv2qTjQoy3jRFuPU+MTfgY/IJY3J2j83bDE6o0eNMzPwW/NKn
QsxyJE6N/cx2Uv0EgiKSsTbfRR1FP0S705DxTLmWeEDLmZc9bZTa39UEXP/IYf0q
eNdMDxd51W0e+OwdoNzLopIcybhNGb3SKrKy1Vj/fbY17J11ioHiZC3HzXPt5TmG
TAOqvjiMi37N/b1B54kwL6uAzvK9jKHbgt3imVojivFUR2DLyDTmGKu5Dug7Q+ds
Sa9CRz/rY037OE9fSq7Z3i3rX/Y5wAhH84gwpqY2eVYJqDP0+K+7blt4z04IiC0Q
8tjDmW2zNaJW/ghb2kpoGb/37JMP4Ttp3NelZZDwtpvJvigdx726mCzpy3ar5qJq
s6IZScsk0K6h3OVQkixlXbGGi9bdt+8j7bF4HQiDsfVEMyACfJjmjdUKxVDSy528
0zpmfyG+TSmvncYCw846yyHd3agWeSOTos4ciJT2+fb3a176dMSv80k/TNw5OuUV
nDz9uj4C6s9YAYIeW7RqBySPzAbGSRU0MbClWJUuNvNpahsrQdorQ73Bh1DiHi/C
bzH4McLfHRbs+WdItkfhEMkEfnYxvz1doI7sVdnH/q0+SqSHx/8EG3lcLGINafLw
cFyGvHzyiwAMGITJE1O1u91QDZ1q+JJm5sKYkl6joqUmmiZ04lhJ4CJLsGlWc2RI
huiVL0E3U6YZ+dPiyfDzVp58QN0Vdv4mlXTNWpTOIqP4dj6Srz2BiqK0rXt1zvN0
UpXhsm7O6T+0xiiduc9bIFVvagjey5x+GpEaK23fRv4gh0HSf+d+ftcsY8wwVlLt
u54gBOMOsTyr43VI9r5bcP9hxButgJoDrrBnzPk3VH+M9CRRzzDhdNDTNpDTDMFU
u634iwnyik5X3NHQi5xsFkv3sOdxfucy0/OlIotCNPA52gMQ5svLp7UoolLS0Ifd
zK2wYemr7EzFSKBQgPENoADmqm9ldkYSmQH+38J2UgY7sr7Yli38l9OPxu5Wr6KY
uyGOQw/5yUjInYYt/+mE+xrjvr65tbJn42EG8TOZaz2oIJCoGtBU82pqktap02WG
CYImRATDqIgjcgAu03PS2/BN9ZUJFVrXQKJRQReDzVtyMKUL82rtQ3dLPcGHLMmr
p40xJm18nrNj+9wxqkHYfSzwGWP9ZUEF/UTgP1BCAzdWfFBusrjofyYIeAcMDGUp
/3kgwwIEXGVsDtM2I5BZkHwf3HlABnHcVFddleYiD6ZYBzZRmONQCnV2/cfkrj/s
COMdlXd7ulo7DOJyhQKtwo9fVPvfd91MO+xJjP/i19Xx1VWWKcQ5bfFjqVEo4lvI
zwXa1Vpz2PkNI/4499hv/I4RhkqXPDfWll+DtNvp8jjswWsF03Vaqno6fIfHx9Ty
aYqAWVzeXlFJcq5C9GBke8QzvTehiv2Khf4d5zVZvMNaPhw7mCsgYa7Lxqsa7Z7o
h6TwEYS7bvHoSaHxMz+3jnDbAaXsldCqtAsEbbtJkg77W8sJnHnV5eGpJoJyA0+n
3ASKsXvNqEWeYZ8ZEwiD2aNbbFctgPTTJZnizibJtNqE/h8qXKI16yP42dB9DSpM
i1Z4erJ4+6OX9KjR2XD9mXxHPoykajcFo+sK29Yho471Cgl4EayqROBHr+M9w3pe
s2cEq9QoX8ku3oNR7sBNFbum5+fQkOnHLCySGp7LQDqdOsAqJ8v4EsA/A8RhweKf
kecM76MGHodTjQtEtUNOrOnQVKQuqQANq/V33/PUDpYwIk5o+Je/lSc1Ix9w71Lz
3BGczBkFgEjIceZ64bEtCCfx4wW6WnN3KOn3pQOZM+WLHXbS9ixA6e/OCWbRpkVx
fMUEE6y6SukAUr1ljg8CjxjCWL8V6f/l7J80OibaOlyG9q0uzyJFywIpVpXG0LiD
zsWM+tYdv+6lOeNC5IuCWO/NQuf4ke+lhjsFY4TeM/U4+zWn70ztBZgxpGebVH/k
F/5HC/wapF1kjpVoYro6I4xlP+zfwx5tpCWLPs4SJLLW1yg+sJ7CGTlTU2QalAQm
zhd5ixUnW6vptO5S8LBChwdMcQSMFjsuqWycNE537x7mFgcUGUKnZn8AAzpLoNrN
wDLMocSwZrLoFTQHACHJFtRRv5fBOCNLoR3eFLo6K3F8P3ajr5WsB1uc/sHdfPjB
02sDhtuhAcpvFS5dKNm2+9ltJJAi5McIkxZhqAnR/Ve5AhbZ7aiEow50U+viG0J9
JUnuE4W50bDztCPIFUWoshccxaRxE/0Ja9MvDNMGnGo0J9kuJJBoW0M0vIBCYST9
xFzVRhRlVpuaYk+X3gM/h3MxjtOVd/30OiYoWHFzbjue+IxkY3bK5/3qnVsZgnyC
u9rVHBRTXAnpS1ptS4YtjTI42v8AuOUdfw2vsaPPqprf4sR1724mLhfLgXsQFSVV
sTs1qCBSo1uDEAuHupgKR/U28SLRaOcQB1VezWruc4xbIQ7oY6s8LDWswffQFNgx
FLOOJlEu9WoCaYJ/omlvvTtGBfhFUdEVHBfVALqbQCPru46xLK3zubKGrnhCX11d
qtyQ9YFLLuUvBssLZQirAk7GF8u9ZDDZ9Oo0o7vDZEKFt/ki1kh0gWPeCU/szwnj
R0Lb3nsAXCMGT72ND56K8Qo2W6VlM5Hji0d4fbOF/98u1RcZKINLUmUm44aCi1rO
9KWtJdAfgqSzw1jDe4TWDoX2z+v4S7CJ880+/AHDUS72JCQ/+HdcMM007OBtkYPY
hA0vTcvwfuVfMlBXC4qD5ZYbRULHuwCRdOHZoKx1nzNV+lcgkH5nC4Vkew+5vU94
Wk+qXVuUnd30Llvd7PAByGTJID+8BRf+nRNWp/lP5CvofwyMkdHsyIzZBsyH9309
AaPJyxuU2KfwTLocMLSrHWKJsFOjMwg5AAeaerzY5llJO0kNbmUzQwBc34pUzvst
5Xi6eENOsP3RiJNX9MUFMp/3gyAulgx2buY3fyvaA5YPEnfp6+5RmAqY1V05xs+v
+vP2ySo2JeSphghYHne9LVDnV07im6EEDK/kDTjPaQNodT4VNXfUeIt8Xg6M1yYg
QgMenDnY4PPJvh6MBN0APbkIc5MuQqzcnD8sWkNN+M3gt30MPxcrWOS47n/xyUQg
mCBDanXGgLboyWiV/2uYjynSSuqfciCMyrful+dF/0la6lfTRrxNMtY20Xom9JU/
XtAV5mNYDBiyyvDlkTCYBzRlYx9lIij/TX5DzXbR4l/TwaV35cx3asVMSgNbYQ9z
1CVYuEnNYaWihnIYw7fmxOe9ymA7rInvZ3agHI+40d6NqM3IJ/BF2Af+v2GS7U04
eNvkTymX7rVwIwedRrGwE9HyrJSVqcBZcYud04vsebjb9j1q6tpHPS5miscn+Avg
ibPY46jqAtccin5Jx9Xpwgl8Mdpnqe9Kblv2cGVf15S378FhJ7JtB9CevgHfgCCa
oJgUFq2sej2+L8+aPunoKxrWnClnE6ivTVv+1vTnFVOI5epa8RLwoxIREIQGQCpz
a7GcYNtggaM6EelZqiQlSRWILj/ppkTm0kbX5Q+apxzydjZzO5m64C5e6C0L+BVp
1/XMwL5IZ94x//3ecQA7mNKjGGviHBf0+QN4Q8xIKtw4NW6qacVtKaF4yFV6XmQ7
lQnLAs2m+T5uGhIidvGO/Yy6EKxEeA5DGRwCM4+8KfdUL5e8aqzSOivyCG6AvcNL
LfA5wg8Auncx2i/zo4S0QIUNxUUKVIpOEwM5eWGqPqi5ecvbytlCZCf2Iivn1I+5
NeLIPfOl/Vxa8/IQDAwimrB9VITn7DcNfn4j3SCGKAT5JWXwA6RaJXrk5Nd13O0f
/N+P7q9cHPgBq2LIDbGLKihTFkts66V3J0YFRoHbp8tlpVcK+SkdbGD8p3nTW8zU
zKoDzxLRlQhtSeNefrT1gW4g7/guFITwOAS86hSpvvU49TcBZCOI5k38ZRUVhfaK
2cEzVc6gUsOgIwNUoSi4D1B+e67eWo6qPqDqYPsKGbct5Ug14tzWj3nnf/ZKf0+0
s8jPrIoypJATR7wxXNQ7WokWoLKc6gxC3fiG2eyF+nMb7o00t+1FufOJSyzO4HoE
rAWBWow7xPc9c/Z7rySw1D08J4X1L8XQZUvIxxhGhlrlvU5EQ37C8VKJBOrMQuA+
8We9mCLIo7A1B3IAgo0l78pX2QRhPGxZbnocwxqPLUT2fztrbqNMLjXvdROvlhvc
VL5GGP6moXna4WJDdXbEb4I6pE2pS+vl8YfUq65r8VtrnjNQOSq4Fzriv2gjjqXJ
l2bbXHOzygqMjDee/vfmxNF3wxEZ9k2RiMNOFzU5Pc+lHp+GF2AdS+ylRUfq2ory
0+NIVpDpDPKuZphfAtDsFwZjMGbw88wl5IfX6DHtL4MZFbr2GpqHVgD/EvIc+ir2
FSSF4GnTzTbLCTWqrnAcV5N7bmyoQ7LZU5atknv5NWFNSi8OMBO8yss4fEUIPAhp
iAh0usBOrT+J4GHGkDYkBaySP1KO3kThLW+nv6oO9zu2Q3stY1/oaSPob17WStHI
x7TNrsbS7H2VGfPIr4+SNQKsWb7Lr4LCNtFO16/Sx/5udTa3RcW0sbFw7oXjsjYh
iQ9pL7m3ppadGKVMtF87/TeYQS/QyEB3VLsdAt9RUDKOfoMSJuMBcTrUmmootmaD
8QOEzeL9J6rKs1J2OtLy2Q1aCqxX5L2ucpFafhxaWwzGVCT6PLyzyOhj6cCG9cDs
Iek14kDqyorqXKHiigBIV4r+93wnp8orAHw2CnL1vu7HZOVPG+Aha6LLVBriaNGU
jiWUcu27puew4EfEDIgI7paPEEX67I1VRberIt4E6NXF5oIqCo7LiFYwfQxWdBfY
VD+61o1zCjYe4KUuoEVPA3t2g7PIAc3p80vd5ofTsZoErDaO78UnkfiRvITHD2YO
GVqN/iYSMVkKVQmOl6I1Z6KSxdK67FXiTWa7gEQtmGHKpuaqn9LVAsqFjjWg04ka
9G2Jm/o6AkcLxnMCZvvCVuLcqsvNCJCNblKKv5CKdBMRNGoM6ydsYed8uCTwKud7
p1poPju+cvvyJfDgUWshKF5KrqRFVC/Gv3IDobz0tEWkHlZzTm4JRQU2E4n1TSdz
+yEDOtSzr37I1udlPrTsZYfsIWSg3L1Nn0Y/zEBO41Ul6C5z2VithRYiNPclFt3A
Kdjoy5+uzesp/v5OnTUMdayyvWYu/03Cg7VzrMW1a7ChlY5S5JOw1NJNnRrKs3ge
ywYaj1kHU8h74GcN8ixeg2mXxDab+lG0+R3dquBnPEn+mm5LRjOq+SX/u6tBbSUy
sCeQ4hIl9nqqq6Jn/cEzdwueUrgL6pgWvL8di9aR3IuS7g/WG+HDzZw4jBS70BJD
2Xxs62tAsqE5/wc0KT/t0IAJhAJOPTytL2q5PGuv9ht2GNx3+zQZtKh20dI3euk7
TqHPCCNVjeTSac1hDNhiQamMUVCaKXZIfcbe9+AgokqLkN1CbpWJheunkwMPwV/r
N2J6bsurkwx4wm8p0SoKShGirscEdu35CMO2NgndlyE31nFU6w3uXrBWsYIluuzJ
8MFqZObZ1uJ7EfFW479sViN4XV9ix8Up9Y1QWz46iavWg6NnHD0bI42sVDw3PIoJ
k0tUFwzekW4AqmFyb/gaDEpE0VgbmMiUPVCdMePmXZvnvkQItxtzj3Mjn0Kt4Bgk
nyKPQGCyJ3foa5k8DbsjSwgCyxVI82oEcf2MxgJP4zp4mlQPwWAz0odWVgjZqRUV
xLL0uXYCigJabJkip/o2cBwOzWHI89Ys9MV6/Uoj/6c6/dZKrOiyeJlyOz4lkMzt
zeOXwxpPweXPMl6S6PvdfypWmph0iQdRn94zk2h4+GwGs2/WpdMiTsonV3PejvQ6
PblJG6b0kEbcRoJ5lDRLQ1crdsj5twJhK9voCQFgMInImTWGPqnMmqUE696VRwFZ
azFN9iQW83iiZ56tDS3huURyuR6u6KH9YP82OGkKSLMz/jB5LpGpNF9kayLXNswa
Gjttn6tUcINjqOHRIy9GdT0fycBpSjEkf9kxL+fCUfMRqSteWHCoXY0t7fSMgiFj
eDS+FfB16t5pxcS4ySbfFvXziv+bUxhm0n6qmYd8PeIrFi6Ig2yTPr5ASpGpVKT9
ZD5jVP430wakRIF4Yxk7837b15zXdsBXPXGI0ErFyPkADFOKDzTIX+ykLO1418bO
/s/vJZUCVUn7O5UIM6ACV0HGlmw8OoVjQ/NhaX3wfPnfThs0ZL2ilWjkfhrvAG9/
GX8JtJcVts90ag8VmkUOkpzbqKmBax5eAV99E9zbnmgYuVJ0mdfaVZAc38KDBY5U
YZB2vNJzJ+errr6bQlGPoBLj+rOKE0iTuDCMgvHiDvhjPj8J7kL5DNpJwrjO+DqM
hSBVDS4kFfjoVRriuT/x6Rm0xX144A1cVvElVZXrGxS/tRge3+fijPki3BsUm9Rp
JDdMTKNQ1PWjmijVzmbbIDzfoKv0Irdbeidzs7HKoJ8I2Eixzq9ddywQaJjW8hhf
tI7E/68zPrNxUdJcgnZSGo2JN0LI749LuuIM6vUZKHkFKCW3Sn4wFc//4SIkTmFF
t2r2CJk8noyM0q/RBzIhzPWaGrLs3YzBq4Kbyj2rl+OtJLBnj7zK5r5OltQr1q5M
FC1Z+GcTseVT79ALhOnqGnig44OrsPIsUjZcj87dkb0OK13kPn/PnMhETsaKDupR
WnTFvrmadATu5FNCdWTK3Nsy4tflGCbp7Chw0havMM9tP6ydZidc0vZ/BPWylaRI
e0PiufZP9+WR4b5RsKyRkKxP3Z3y23krtGlOeNgB3u4DMBDHyPrzY3DI5/tEWJL9
cGrWHzTT1J/ef9jv3k3BWG1KWOTlDtw+UvJsPN6w645rw3NXcl873we+LrzO28He
eWwJf801xahlOjGtZxjDkm3TcLdCEAMWlNuPAxqY2x/zAdQzQ3x0u898VAWt1rx8
2bZmLs7c4SXJVkNsDwWlnFTWICIhP9TsrKGmG0LHA6+A8MQw3aOze0e1WavCIUPF
z1K/Vt+lVV2vGFDdjgUt6hEr7nyadj5QLlrzAQ2+NC+Mz6tJy/hvfxOBrKtKVQhc
X2XmqKyNBvYktRFyPRCLXrrrpNsNDWq46FILVI9HBq32HCpUFmNL8xl0Ck38d6sH
WvIUaRCkeJutaO7nuozHWdUvoT/IwZ1jVqCIbifmgKgTpM5TbEMOzwKGZHck90OM
R2kPvmjFVXIYYwP5QWHBVZOhFxy3/lxhgiwXDCgeQjzf4mrg042wmeW0DoZChdYl
nT/fv6QSpPqEd4lmuhleduksvNUmm5NQS9j5w5T9kj+E+ZAkjLbWfn2Js6QzMwfR
dSf42r28z+CCE6sRUeNaqcd0j854zgU55fIzD6ZVr434a2OUVDoGEZSP3znX4oZS
ipRIdy4f+ZOnON+ZIcxxAeOCNpBVXbdIAuYkNRn9rngRuiqOyNkzVGPhYRUbeQYm
n/X+X2RsPyqP/tbIE0t2Ho6KxJjbNkxFDnlyUIt5vj42nOvvF/1k5w2yC6zp8zwA
DS/92jIHWnGQOFjDe1Lv4TmTa+VrFZT2yicB2U76X/93YHca4kGJdZ/sDNCtfjED
AQjDfQaBwmUc6R8k98frJ8xONQKoTJvUS2W1H7vvjBmPkDArkXJpYst8WwTL9+ZU
gOy8wTuoBkP1+PDqtKTRQJnkgMyN3B30mIkhH4uKVkzdJ9BTl3QcM/riJlZfEWTt
ynHQBACEs0BC9juBjW8PMqPNjNoscGx2WxJPQgt1m+ohvWJuXTwyEZlVt+YwN70x
oAydfGc0d5ihgK/CdWcvnHm7uewaAihocvRFDLPikRPmvIGLW7Xk4hTqvNTnFz/B
WrIu6b5S7sy+tlHr9c8OOOVA/GmvQwSSHrNEF5bcJxw6duOfRKdMVwzRl2EnZ14R
BY2bPHmRQt6dYOtmZiODX1NinKypz4DomLwDYwEOMbfBMkNEjfq7+GKoLbPYDhKw
4uUNKGGkVzx+oUG/xpNDigxkjgLZF2brzk8cZEv7dzJ8zwsKbsOsRQ72vL1I72f4
qLZSt1JqwI7LvNnQhtvUEbAkB6cp3FYq3PIST6Du+bD8H/SpQJJp2fAs991QqVJd
t3sWEVobylJEBUaldhW/hhU6Xn0ryRWvjjAk8xYh7iLwZ1tPl0jj4uxdeaDKgi76
bFz0S7/32vj6oNW7RuOIbS9MLRql+kEBc40tiRLrJvMFNrDxLKOBtv2iosFxB6Ir
Z0wKk0/TgaIfs03/0s4bwqhnfk+RqEqAiGOacjRSGSb6nxTTKMt7AMxRWfhSyxs4
LAjl0v8p7l/2M4KNQxoJcMQ3ZCktWG/PR3IrPpLS6GX5rUtxyAzKu/5AM0JcURV3
dJhA9dOdkGtLNGMQFRZdRztbrA/tuqbS4191yj8icSfpAkUv5GRAllS0BVnaqRBM
AGg9fde+6IgAeBe4aKbYWM1M4lefVjH8CgBOXqo9KG6Ovk/7EzDI9cQTrBZBsnd8
4tO8F0JRnNHKU4al5jqC9UV4tLYNyn3j36lIL7lIFz5UT2kygKLpkwPn4g5gWkAO
aRl0jrRF/xgTsaWmbIGBIPz+o+ldzuSS3aZcH2pZjBmC6WLQ7b8Gvcx+aSnh8jrw
5Q06n4uRGnyCm219HqVeh4QbOObYu+fOJjuGDbtuZ5Ax3EwWJmsP7ORZIpwtZ/bK
cermcsDIsyRmHvKFkMIH6WlxUdUpYvQrN/nj1UWhBtmqOK9Ya70QcCopThcFgZuy
G3aIBcfvGjb0MU+snwPG5XZZlno0AKmdAhg+Vaq8m2ZUProupgP35I0LUP3mQTs3
dNS6Fx2PvVtCqyfCg+WsE/9gWy0Q939TUmXK9oTIOUcugQoqXfRNxGOYzb2Bs25x
hQF9tIGom1zkeHsEefQLuAYr1cNji+6f2ukiMCd4+Xn9UVQQFCanytdwgcG5kWE+
xq5hr3omhxUlfZxL2yXtGJnAvE7zKr5xRzBlTatNaVIWAX22piHW2+fh5twfEnah
WuHYx+b05p7baea+dqaSLl+vCCLJRPuUitJ5qDeXQahjbfR98b1+PHVL92xXKfW2
Aa8kDc/y283BR4SOz7C+3ld+QOoTfyzoHbcyYshvtaGP/gAG5PNeXOazwNsuIqoj
sREylZJXRtQ8lAQB3N1O9Pa4JuJxUui3yzmGFUiQi1rY4azXm3ONry1L2ACy8SY8
H7zfRx2HLUhSuKYn9JbvARVO4JY3LpecxppFFeF+D9ZvKvTrTe43iQVLqJkdIDrY
laAHI+GdHt4l3O/Z/fiAiERToTSzdUWpyIxwwdTqaW3pM8Wj2bURwfWNIBXgVgsF
B6jpeT37857ZIm5gMqvKhLlSSp4xd8zH0ECoGfDL7uEmVnCLCiNzNi1OWK/1wEMQ
Bp34tzKi7fZTd6j+34YHiEKk//C3HDTSvOn0DunX8MxVv1WG7yVm0KCXQZrpKh49
eawvin03DMkNrQjNbEVYRumbg0i3mKzAbIBKyWblws0cfc/E5Hr5hPSn2sqB3kb4
Z890Tm0Fxhil1O0NXttcUF+6qHUInDVFSomEkj1eyrP/8ZPK7cuPGk8VJvt0mMm3
hifvqoztvwypZueh0/JAiV/vsf7+9s+FlZlEEi6YSENm08il7LmvXpklV+DIdfWx
oxVZlF+ycsCGeIvph72/5mSm9Alhu2SvYgCLvEX+aB5xo+l/rULOavIIxqWQdOZ+
i0EOMEBsDSpEDed5SvetpEBdBEwFSl7KzyhSxEl2K/sX1Da+toztTpwOHq4jvltI
k2F3qzK7vdIszPzd5CNNFWd7rwi0BEbZSqonUic2fpDGWFj4GlsHEq+7nXJl7a4Z
x2vTcbPLoAr2h19iGytwMEGrP8J9nx1LChAk1CT9fbCx2VXK/yLhblm79qOJg+6V
QQxoDP7LufnWFRc0O+/tMnpEu1Pi7uSzPHg3ln/vuj+jbCuQaPN+HcruLldsR6Wa
f5iJwaQxZZeBTx7R899tOYnJfzrTXuA/6WYOAeiSsdkPuWVkaHCEPJb/15WjR0GR
Ckbmo+RiABlONhP8jrNhsuaVV2Hgkmsq3f2hwdPIbaNJHVseWl4KZdkfy+Uf29l1
UzbCFENLtMAfet6jwJV6JNuyuy9YxztjFQHuh8H84/0/3n9IQjyZNuwt3fYQOG7K
2x7hU4ri9GiNzcf64rhgN+UqRc90skBfDBy9rvTeMIR+TiKJQN1v9HIbRyEEtE3k
w/C/V3uhN0ijbRSvxQkaezD3r6q4mPIzBzlOrEpL+bKoHGbtqN0UxvhrUTcEa6IB
qP66xfsGb4v1MVCmkurwwjTxPPBb2l9pK2+uLGkRrgcAuIiSqJ2YxD/NZj0qo1Gq
jm7qEBhaIJhwiDKhuoBtmsq2vjU0ntA+siLPR0mJ513+QwAH96Cj8jy4TKiP9KBX
C+2P60D+/RkmgE2nx9wpvpj453QljxlURViEFC9sN16uXjxilJqAc1peHxiECkQT
+5WO60DVBUvZZLdiHKFkdqpBCWrPBZiolUHufycB86wkqj5fPgCDGbhccD6pJU6+
QVpuMf6eul3eX2XXM/+aolMRMvs+r7Rit41GciNWGTG1cx/YL7bom0/Vf1Vu/sl0
W2K5snRXdJ5x5WvRc7Y24sGfenKOT5xMeqYUnmp8dP4QaTTg3fUPLoVCrftax6ZD
NMpy8HINYdAQplvn5acSMtqdi3VpLTEl76yYnNSH8+Gyjjm0FOcTOjj+smOJ6nNg
ny0PY9sVYXrTN7WQ8WIT5dCtoSjX7NWTgR2m4LAW2wAW5WiHV3HGq2s332skL1wB
02dXVttpHpZVgXdgyOBAdncmg6LsJZkOK6qh8QzNvC6Jw/1aIM+Ps9YJ68k8o4Na
SOZCmvCKd/FLLZXonkAz++qlBJc1Aa1jahV5PRiv2+IZXei3upJvI20MScbgrvng
H9jtZbgqhkDei6TFhS5xTJFrUH7RqJnO/ZtIc+X/LMZdMCXMxa+bZIPtAPraw83N
9zFGMGNIHOUszfae/V6PO1CneYsArDTSD5EqdzdldJLjnU4M7mAo/QPqMo/NRMxP
Wf0WakNtlH+U1cnRURznxUfnOCCPoNy1gcy1Q8gZokrGAC+wSdVQAqB12T74NDH3
hOjUa1PTm83xRYqR1FSyKmutspSRJYqvzMitf3CYkXzWT1nrhfSryJCD4XziOjcb
6irc4uzkOMcD0PXROJH2T33CR8uvU0jFWpqvphQJ92s6wJ4qw/oEnndhPvEVULc6
fdXMRPobETB+5L8ibp7Zhzgz4MAAqdEpyBR6nI/vjC4vdFDF85Jnc/iYwLgip6JS
HNr+HNHjpHdVO2pV2HoUqUN+taWHmq43uqP8rwLkIlGsA3UvziWTt9JBez5SEZ7M
/8EYY7hi9EZCqCQ6GhUDls9e2X/0TaGnfl3fm0HKdzERJf3vjl9xVSh1kU5k9dCs
JnS8IIk+hfWQBMDKSCs8TLAUKCde4E5KhFrc5eoFXvj/FC2qFVLdfvVB1U2x4g3F
N1/r0yNcH5ZWF+qGlv+E+Q7FxSH6GABwezovj/zRGSWs8UCIlHlButhyrfDs2bJb
lvZEHmO0OFOBKNFRgxgN6CtISs0WwwMkI2ukTwH9AFie80kR6J4pE4gtW4dZelBh
JehBObyRwrJ6m2z/Nfqx3wtPCV2kluAtjtMT9IV5OQYsRhZvZ8oDJHBoJf99fGrA
4FPh7C4eq7aDkjz62Vy6AxS8OB8kaCp96goDIsY2Z+Bwfs8ZXz9KSfaXDcvk+yaE
4n9wQGIjnjnZeFzBBKPsBGzxWIiIrmM0C+R5jqD01LM1VOwCM1NrDX9BFFm2IIt6
yxHdFyIV0/35R4Ko6zmY9vFBT8aq+pSxSXmqj/X1hlM2i/B3qZK7lrEiIL1xtP1I
DVLx8wiGMEvtfSY3TP5VR/j1Q0Y+8VwmA8jOSPDnKrlDFIOnufEfBH9cYyorJIs4
rHr7v+NguxI7dWcPzZTaJOxMGBgNZgC3YV4xMYVEWhj5jgqXUasn1Y+d5Ez04iT3
Bwtsg3U45WwTFabwQBy/tFbst/qTfD1szF6GXrVSuCuDmcYE4O9PY5ufZ8c5UkpG
v1jm2iaQrIn540dVoIc4sSCWn6CvRUpvaBo7TNW5lp/HRfUjm+5ofZrRb0AUhCCG
SGz4VvzzAO76QjaTTgqLTQVbT+Kh8aGNi6OzOob2tVPi9ESz1CzIO6/vdiwkEE4R
/QR/g7fw6PEZVstXTY9eOMy8a+boFnDIuk+Mf0ie+VWlZwbBqq+A7uaYkK1NMsTg
SECBE59GSZbYiVMjPU8WfWTok65KXyB+mRaZnq2zBaMav8GbcR/MBbyQ5lTOnkMc
diplD2zWww35yaOFaMBh9QqQmPouE0cMPj9ak0iDuYiroUZIihiv6ME/1LURaAWN
PZS/OSHAtJrKOHn5seo4qovSQL+uiFCLZyFYundoiJxfEnZqvlJmZzSjxEx17+o9
AB6SQXPCZHm303AJpOpMYSbop7g6j+36gVq+qXYeEBeSTFaxsiUnVbpL58fGg6Iu
SZ525osavWp7Go3Ut5+lPY9l+hMsLOXX7sE1devJZ3e40DjoFefZewRT5lRFinPe
Kjwwlzk78L3ITxrRwQjwEUUN7EbyWb/H2Rfe1+9QZMIcU8fPbIJI/CIChXFARuV6
3mLfi0U8xTjrvcHozIai1C0Zyy/bHSqg/45SCBxRWZDqqZgFskCUThsjscQClQat
sCS7he/EW6vaGMLHM0kbdlQVl5O3N8M60jdn+md5sDybGuiRmRVJHWcZ58RZ8wWA
3c+o5RzHH2Lu8ZTXhENR1b4Vgf1IzSygq5ZsdjncLcvDFbomAPNs6nhBMaB7VZEk
pTSCB+ouAZ+8HfaDTjd0mulU0kozFixeJdiNMzjxtvcP9wMoMoRvLblCRjFfv7jP
MS4b2tzrE6summtvKGXcJc1++uePWQkDEBl8wi4fhYMePsQBlegd4qm6lKdBhQxB
4B4g+HNfkqfwlgTUok45gGUqfJ97qI0FJ6S4HvgAuugkTgxWa//RO45iwAi5ePcG
sxgQPdEegrSpv4cGTPhFaMnf96NQ+fXBzvtcATe8k5+6GXpU3XExqEa0YCiNBR6I
e28GNI+HIRbehMA1kIZQlC4lmqYapiKqjyj87b9+M02RnvDHT0NJPfsBOKVhkVSp
WbqpuHnkx360LqyKJsNA4B6bpN89eyORslhukQmKNrBLSyPxQJfzoWrxXu8yOUnJ
JFuttI0Gk+3G5RfSuVF9ykxIsjWXYfaxMeD9lt3pGOKLmT6Dli4K5uvjsifr8zOS
iOuC+D5cJe5CJ+4oSxNUlpGi8b0U2XP4ZHbZwSVfAbTww/jCLy0htbVAl5s+xMh4
rXnBkLRSuhvDUSbQS7KzmOMPyQ6/fw1NrHVSsjMWjQJT+ojVnlhHHXYLnzFM38jJ
01XN4rtuEM1DM3Ktbcq47wtQaBfQZ7nI8Z8KVy90tnbvZ7PXu9KEmn4ey0wfSGKS
SAL2CApP2AYiEyQolRilwvEQtNYBXhEZqFW+nTUSVQHilcp0WlxljXwpwNJg2tLI
XN1VjwhdKjw6yYMQoCHLccq4POFM7MB5ufPhGmvt5YV9UTWHIoDg1LUIhmTL1bjx
Bb1oejPu6tBif1sHiFAJw7oUn+crdcIQuqKyKSVygUh+W3IGScQr/wTxPum4Jiil
T/YUYKmiZZMKoYkTRai8btDhWfBqa5W+4cIEvkyXmUDxeuVRTpI/IQ9FZBWuou/m
pFoAvLCv56TG2XHx22mTfOD/FgrJvqDIUYvssabxoCUwg5uyERGPFdLHim7Az40O
yYiDXD4OO5YLc5pjgrVWcl3/QVqTviQwTKer8dqCoHAvIe4KW4atkVvGs2HisttH
/4vBhAOR8fylWCXQ+WRyF/QnHvBHuRecHxU64qA2Nm5U3CHOBs3F2xmNAHWAKStf
b4lFtydIgHsZxCkzh0uw8az0vskwcesAwq50OmzT/PFAMTOomzYF9J0WT3H79Cpv
16Tfn9PGc5Y1AJPCJ/a05RPXlb5IsFANtQgtABRPUMGQtfVrAttLQCTiVHc+w3HY
Vy/MgWNIDwwlbMPmHIiPqjEr7Uaapz2TGbP4CBGceKR3LJ2NwtxOCkvJu+buO7ES
R6+1YrVDvEUUAiwVlJZCqsejWMZHdzO2Tkjl8T550XPqTGPJtwDBynF4cBfWK232
7jhjxjLgADm7q5G3x5GThw+YF442+B5kZkbvEdavIPn9yvjomhARPJAtPHD2DamW
o3eLs03Bc8qBMqVmkjH1eNEEkMfdPBfMdw/pnvQgwSK5eTTeuba9qEsW6KU7VsY1
1Tg0+WiC083hwGDQnGo1FbRUrR/GuZ/q0/iFZ9HzSbUwPMqskyeC7ajmTa8Be8Q+
shr5CmMbYHAWVYNzEnN0/leErib1mN0vJZn/YMpEN+9iB8b5hYrHXlVQi8IDHaY9
+LdJ4xTyHndI5YAfa+b9pqsAWm6qmML31J1jpo0tLpkOUVol9aLYsBd47VrOnSMq
efS/MLQYORgeOIny2dbN6k/e//FknzLBHNJufkc85TQwoyRDBLRM+1fLnu+S+rfI
73Vq2+4XPjkQbsXbxn4ZghAPEdro1CbSj6ECLTEo25SUs2wl4vqFYev1/szA7emE
2S9gnNnhXIlopraFVLqOETxKlFG1hreX2DEntF5+PP65a8rRh2873TWBSWeCHAgF
qzd7fCAdxTPMrSYxPkzVYy9Aps3eqKV0x/39tS096XnZ3gmgDTzkLMRVObZVVoE5
Yg/CgOXOKFpb11s/FYwkVLNlk7mo7KjNqBeSdYLDlc6FFbS2idIREdE0ezfK5WXW
sjbiy7Tb0CGdqjy6dzxHA1HCYLBRa4ywLnYyixTUq7PBRifuy79W5xTb4z7KW3Go
GR/rPLg3BMpOCcD6tR1Kxg9seKzi3xeqwRxX8ejFdvPZfWMECCUNG5byiQXS8v2V
gMZwRqVfmJl8OQMKUwBHPeH1dxJ4swI/D+hj4Mr+kSO2gjeXEC2NBuU3BgtUPzSS
kMuLJ9A2EwsdHHWleDBIysNfx0r0po6hIl71nN2gIQEeOYQTPU+4ER+CGPLh/nEL
TS4o5Z64ih47NY9hh7EYjaGAxJ79/Nj+YGJ8plCFGYgU/8xdOajRuv0ss4GqvOGm
1R7fedWzzhV17KPxmpgtndaFuEOAyIdmkAxkW+f5dw2Ts9o2dZsmyt3Wb6O5FaPv
6oGE0G7SyZ1VLsNp24n24EhYxPPQ8kl3TWuWpvORmcl945x8WiOQ0Irp/ufc8FQC
KdEVOecH5IQrHV44wG6+9VT1+ilsaKLTQkUNbdnYYSliD1MnOPDWkn04pSM0Bbxb
0V+QAcHZ6cSQZnuNuqWC/dn+i0v8sdv5vbSSyqTdiHKiCsapTehXlWw9JurrB3OR
d70XHB3yd8l6Vswu7oA7JEy/tX55+02QgsC5df9+x2ETOuf6pQQ9MzY02cXelmwq
G51iTPVgL6j+xYl8xW6GGI54PMPO/LJoqY8h0pU78PSDoOhfIV7E516hiX/ImLNj
MRwv6PPIN9NiPPiEXh6mWusVdIFMnWBKV2hKUwyd56l15WryktqnQ6ilP7aG0TnQ
X+ACvEbB4xvU3EanASUWy7SBIoYEmDSH1eXvsp6y9x1p1tHPuQS9eIyLGwZ78QVF
I+qzRY30/jKSiCmaLIdoO2L2ZTwYl/ix5v7E4M16fHRTDTy2uyvJCT9TF+b7v6D+
lRDJ6HLy0ao02/+IBMMdGFDO+UI3aDVpRKx7ppdb6tJjfZu4+Nsx6OsDinPB18PK
65SGMe6V+BZsohHtt1ZK/b2AfnQGMmqdvgkyUJaRvsBgmBNXrwg7NzyJkYI51Ul6
f2n2qV4ub/ojbYtP5CMDVEP4QFkYhXTMNLC2YSiloWdgu1JOHDEys8sMfUjCBSxZ
+wqrbm72NnZTznS+Tp/SVvJu/ZZycSYGuGnYLe9crJkpagguQRaokx3z9RR3tRys
WHdo6LDCdYv60LCcIhPQ1awuatJoF06KzbWJgzw2yuo2T2ogX3RUemfA2hjkKY0P
y9Sx2BtR8tMQxPqdLT7TTZXEWjRxQ6cJpvNzXhbttWT8mAw7Y+JhOasxfWlINYHL
Av6Y76xRCiv6N8JWeEf1Q9Fr+0udZIR6tX8g/T8VKy2Nc1fBfKpwNOGIMxW3wWlx
w4Tam7BaXbdtrgS5oAJBq25udExW3UaOT2QNEK+0eaQ3rmUp5OsbZrNIAn1LJ0o6
Wqzsd+H2K4lJoNTazyxoqw5oTcNHWqyhooAFisM5PXCsAQtLh3o62g7TD6+4rVaB
CGSNPLSMLyWXPnk2Aj+R1B1kTWnSloi1tb/jA0SjLo2Ezn0t6RydH7UNgVjrt1Yf
AGmPex8uqeQLockMKQEPBiiczWFVIZ3FTpc02eVeDNEezKiLcotF5fwOyXbWeGqf
u3OhUaPcb7PrSSLuXQ/X2GEoc1sW8MxJ/s5zoRh8cZWVmO05SBDqBxwrm9+59IBk
RJRpojH/tnCl5rPDz44Bzf2T7bZcKF/n5VEdJakGyGpImLQYkpaZaPTmTreK0AjD
Z2WD4nfVVvQAyGZLOMShlVMK6hWjU9GSdyhXgHudUd35Hu3a6tp3WBfseBZ6DFfr
djvCeM+0tYeKoV6+lwQTQZ3Ndz6tzGFb54z46OLHR7KqQdEafDkNiljuIR4oJSHZ
8Rj7TL/gk7IG2/suFxSf78sgrjp4RI/sxnka1rxtveRwadS2K2WoxuFvStmhhxkz
eIPHx/bXgC52IrQb9MB8m/lmUyRqsv86PDhkUM5WIuH9ca8P0aC76seVlTyznpqJ
UMKD2FmOrygB7S5ObaYCOaNd2CXfx/tsjfyI05pClami3eY8CSZo0Ph2lJpaNr8w
iluIqzcK4siwVyKD5bhp7Ywlsi/xXiiJfmW0/RNSAldaLnEL8dqmc1TmJuV1Tnyl
GiAZBtXIcbxMSlNKImPPuX97mXVldaO1ECl8/+bFpGGvDp0fOjy3u+1AjAjZWYWs
e/uRKpRSbOYGe2NKT4Ip+jlvoTOwp7gw04ZrlGgfXPU4FHZHZDuBAUTsPlVmcm4f
zCZc0X1dkwRmeCNoHL0XVSlAtRjn0jLDlSQl5I0DAFOg3DZjNRnsaw7p1yDHARrh
xGkqepY0ekbUNR67rCZKTWLTg+BKc7mM49JaNI8kw5mfU8scc7JaYLUvItiMAKqp
MMwUEMfXI0i4U0DMBPlxF5cr2sDRNRMEUNiZzzP6JhqXfxHY/Xrd/C3i0XiOXDHX
h/XClVaZwIhVIlzXQRRk76pJyz7C4ubAepsIFtGxNgdjNKqFQLoYszWzCcXJQaJP
3kcg8hsAhG+76WJGTSLdAq99yo+XawBGPJq/oE47AubLg2w330OPhRBE3sEUfThD
kp2d2yFn2xn0NFWm+/eJvS2A5IzXigyqwPM5pEnRR6hI1kCfqv8QiW5clVMtXRRg
ERa4Up5Pt0J3hi4RBQJ0OcDtxNhDmEcwZW0nfAimneanf1Qzen4YMKHKO/dyTzc8
nEr0MSSxtFioi98DzwD6MmMArK26Gv6cyl+IXcA6+7zwPz2R99I6YJ23d4b9UxKg
y0c+aKnRLCsPu8j0nUAEZ3q8plzFJ1TzhlYcqhxK1OiDcgVhezxXsMGhQaXxvPJc
hU0A6iFpZVvO3XGar2YZObTYQF1wqJ7WmhZhmnxAiAizhOOQ+OmI1dWq8nkAJbuh
nVNX7Tr1zReDyFNNdY80vjsQbNSeTvGmSBZiiO6xETNqjLhA9Qf0hRBrVjSQPoJV
jRxL28qV3nB/qU93fiZMmaazRXf6oEfuLFs42jTthUzmGIRYRQ0ZysNUIAFr3c3P
qiB4+UEo0SOzIl6egkYFnmhA6sqrctdyvIcAWIhN04uF40N3gZdivkB9/4IlkQiK
8tVSXZ6K/vfV0toHzOoJpdoQAJwwJAccN/DkPLcWxSadIl6C1TyY8kIWSqH3J7a8
FEaXTn3MsCUeu2GGsXkJWJq8S0TZp6UZl8h8jeC0QBYaVKl6Y9wVdTVSYXQGrYH9
k2SXGeGvdLzeq6PD5NISCgMC8GL3pm90JSDHXrDqKZoP2JBs+sEOyzrmquGe84b7
cCs8K4RrTbaT3/JWhqrbTUpqFByLcNjXWYvVgMbPTIaBUTy7xfHWJlCYzhy/JVhD
accU9cDu2Tp1OSnjC7OxOPZ8fMtZA5lkcZrRHe15fAAxuVIx0ThyXz1Ahx5ZRifY
suN1sTgKFsk18TVNo87ee0SdSn0n3bt7gbgRirzv2PpA4AZcVQ6Dc+g0k3/4AUDJ
qHlk6aAkVsfCxG+xjXwr6dtm4sdGCmA2kqzprLS7GAfxqnOTuLaDnDsxczSE605R
1izg/yia3t0qEGcyQW8TIV6AmaLxBngfu8c5PX1F0k3EIRR1IRWU89UQrnk38HEE
t4Z6pf0gl9JebRgrApZ6u6P8hFblYlQWNyAGLUipw8FityYLXjq6wKsPPVvluSJI
p4VnNPas+Q0RnzSiDAkGqYCwAnrnTkdeS93Oq6c5oyBUskP3wKUawDjS45+dT8nF
9KPMdVgnqMAkuNdFee7mLcP4FM3ZwZmuQz498eVnJL64ZQLN4gyVwSX/v8qMKRfH
De+oqrsSQYwTg9NJbSfmEKlV6uA3k52KwxBjwrOI4N5oupTFP1Rhfo3KdYxsdlhp
y5vSSKDSepdAPGUVjsdbtU97bjQdYPlVeMCsdbiYZ0s7MfAAsnZqMf3fthdxFRef
mZE5RRFSm83rbplvZxZcnEmjsCPSzgMinAxlcGU918ZGRJKwWlGjocP3P3wNjCaO
5qzSTHujVUw1ymejPijMOeNnqu+KmvAWlMnvzGhC3Le72ngTCoV2EuqaJJ/jtS2J
BIP4YhKNqIATCYy2wm1DUy3Z/FtoCwOpbBm/dAfIqvO1jCi17LBkmUvQWvzHWN6V
fY7VPr0FXWar4a8GvgPjfebh8ABfriApkZMkrZjtOw7iVNB6FzLb21TNzNFLReir
juTx/8NwG/UvVPNSEf5vbDv0q206XdilRRRfo8ZjdOkAjTUo4fyRwm8at2s88+FD
Rm9STRDrfDKGmCAX1cRk8YpwXRqhJ3clz/g1UsvluEDQfJExr9sZWyQau50PVeK9
EqGAFwMLbew0MjOHdYc9Fr1YKrVPEo80zRu8xVv15kqBItNrmnKbhYMW4ej/Tqeb
6wI1I9NIoV6MVq1Vs08eilEhsrIGtQox0+OwGbxcTiLYzqCdqzJq6xALeaJVH/JE
SOIXbvrTDEfWgsjHXDBDq5cxhE96DuEDidzHdrlDjhpqDyohCzpsl1YPO2wgLFlI
SWxUe5ttgKBRY8T6TWIrUukvoYQLUNKEVPL5Cxu+rxanrUkv7lEyx7TLUO2WNeFY
E8vC0WU5vHWIvpy8tzoLmmJb6/iQuku2lHgqiPrH2x02TVo/Jb9w+sH2abU6qD2B
qmyctiOTZJ3LiqN2Di4D5EVvHfnDOJgyvPAoV4/Sls3bLGx9XSCy1TyZmVwJeaD/
+QrZcZDWJTqciwUaZbXXk50WVe3rGUmREd8apvTUHvZ641pLvu2ixIL/2LmeObXf
xxMDfTB9kwe4f50CXTc6G99TIQLaCTjp2ce9kCdI9xLK7GHwp5TcnPCC/D6QveeA
Hsv3RONF6/xD1ehhnnf5xpD/OqrZpSPwJFlo4oTEQ7bH1sxKppjCB24YvP6fR6Hh
vLoFVjcy8aOlQjZK0vSJ8nfKtsE0Xr8IFwBTJsCuikwXSnC2kGQS3THgnR/SowCm
mpQfbNaI/Z2YKQlDQ/cpuNp5mgRBHrK63hW9ww00/L+rP3lsh2O4erXE81sESF3m
S8aEE8atk7uGbsZBQFARzWtyO3Vs66ToyE5cXUVASZUKdKyJ6B24ai4+TE7ZtXqE
cwPlFsbRS4gR9PB7YiYRvf0bvYo8GX6I5bLy+ijaOFtXx9/cJa6agK8jEy0biLdI
jcTVL3GZICJb2Zo+DGW7ju2ZYFRLsd+mT4IzeeqdbHA45530gq9FsgI7nkt4Hmfz
62ur+pAIJqlgbX3OXzdMer+Wm1Nxw6qgHOSgotFZxR7TvtulNwCehbHQgKIFXZ1F
7/CI3TZg3rwxCmtRPc9nyQXKZUoNV1G/PHGo7dwB3E9jPFtNOS1EErAsI4XH28ts
PrFiC1oWWKddPWO1erq0AkFhkdZq6JH33NdHjSCbjwZPC1DDtYMqrEmTcUqLySJc
HTjECz4UaX09TnU1gt2ozni6oXZ5NDoKgxfmfiy0WF3dxVqeixX3baQhSV0rbxT4
TaQEstCa91RxQ91C4s53MQ4JwwQTgNIN4VZZpN24yazg+eXRgzIPb2VaOdXZa3Yh
l4w+eCR2qmcGncksJCR3AqV26FM4qoWKHiP7AtvdZyMZ7YFeGVK4PY4MEkgRYgnw
buu+f3HkLBusAGIFankSUO/exPaCow4Xokpup020qPpTLtHx2l/aYskYuiMTDIHx
LD9KWnDQssNlQ+qqdquwU5v5PDdM4MOjFj5VR02zIP3xRs1Ols5LLPLGm53uyvQl
yT3yJhb2k/CnknRwFUlwY5uzAexWPCBajcNtqZ3FyS+Yt00Yzb3ZZtVgLwhKUIUn
AuslWSps3wjB7WaK1o9+Jua5XhlfG2RmHWKywakCguo5UMBs8FpnlXrxPQhNtkP2
jGOv4SvUwXQ0GktxpyKQtcw8ss5cCHAxRsTCG/I3ZfTpS7mFe1VSPAc2WWsVHw8t
ARWWrLohH6E1lmkgLQvTIQ9Hr6cOyv1aUU3K/Okb+CXE6Fah9xUoG3tym0Vrpa0J
M65VqRJM73JA4GZtP7Qe8RQS9ZVseeTIm1jmnhmoAn3+HuMP4ZHPnmRU4an4g44K
D2/rA+2REBCnjz4L80wFTF+4dnhEbE9xwyLQxqDpESYVjMZC4Nw0RpwPseSDwQ7Q
w/ny7WbrtY/IJYrxhLtGTM4h/CS94OE7f3xqpJuvl/9JgBMFnleOB5SdiecVhCUP
Q7MJN+EtBJ0m1gKaev09tPqDFPAknXt/k7WGWn/kvJrZFqDiePUGIlwEdpwiuUYb
3OGkyRdZDAiEmEkr+foTmxauHHONu5RkrM0MerD0+gW+V0UXgaI8NZXlOi1Mg6Vg
JL0MTTvwJyg3ZfEkqwrzgSY3pwFboze5gigRjuckAWD+tVmpGRGjzEfiROQVKvYW
v2hthglS72yCvo/ZrNmWjxZ82ZcavrFP8zbME1PrpN4e6CSUdHVWDBgbcb3MnCO+
5ZOyEHnQWeS7vGMqJRpwqzOccbK3XhYKL7WFisrH+Gswh9T2gOR5EEgQAMuy3p5M
4yIQpoDK7+/Gp03uMB7vwLZGL3557hyWV6ClpbtnRXqUW0fQKowkIOeImT5jSiTA
UndEexmERUjua1T440/TiWs+PEJw/TsfyWQP5oV4mb5YtoChei/zlkYzqEAlv/ds
LaPFCHEnxtCmzDe+d1JDiRZYW7QN+kMN9mDNOj+ylYzjf2pgYZanrfvo+ewBETgB
mydoFKIwixzF3zqcKk7r9BXQsg1vHemAVaNwagoaIAyozGMVOOweBMzP/jDWvOOt
J2/TUXQNODR2tO9KX2NSM8uWge5l68ns4kHg3IH/00LwclWzelZucIQgt2SCkKzl
cPflLT1qS+WlMXqxZvJuvNjvD79x6HkpIdzgyk+AbNEm/S6k2335bMK1pZ8KUdun
GIyN4SQ7sy8LohLIuo4KyFNe7G/ICdEDsLqATGHLRuTC1GblYMIFE+aiCF43YDe1
YFjrvp+D94ioyBItd63INnKHipFK5LHySOWH5z/ZvyJo7ByAq8T6O8NeKbyLAhrD
tRlcSlssRM8/utT99BCt+2SRbWrjf/1eCqwxylJczkZKykHe+VyDjbhl5nb0+yMh
J7h8es5tK9VPvZrtCjERCBt5W233k9PwopiSISlKjnRBw1OEK9uAQyqmB/0ZsNia
pcHPe8j/N+h2y0o6ePcvdrsdQCTLh2eZJRAmkNrA63TeNcTH8jVNB/DoIn8N+ckU
9rko2oPpS3M84CR+Ew+BanA885dR2RO0gwjRZwA5A0kDzS5k9rpfaK2vOqgOrt8/
czcOua/Ti6W0RncV/lbI+CBCdy5tmHoLnVXQQjMXhtpU9Sd5u3fLJD42cirzcCdh
GthVyA1JJFGmWj2rsaJkydN/djRu1UlCMcAgJEoMTsfxUxsfVQxMKxDdGJkaEUaT
d2Z3c5xTK/lRqf3khp1w/MpaMGVrvt2vDHe+pimDPem6tzPqGaL8lWD5ZJdiwumy
b7I2FqhHSg356QCyzKT6o95qtCi4Nd86Cj9SGLD4iUf264xk0T+F4pNB7Wwbk53a
Col7j8Zn4uPxK3XB41e1XO7yOMXE/Wfm/JrC78DRXnTXqtO6o/ffbwzu1F5ylnw9
6+U1wPCihcDz0Bn/ysJvmF3rDTi8RM+Y0njERqiN92tbgtod4PJ6DSdmKxGDWuxo
pLdU/TMcTlJBRiBq0vW1KC8JUaXziRCSeKn8D0xATjj8/n/0Z2LHKLHYrEQJTTFb
Ytp9CTmX1pL1xTnbxRWp/GKoS4/pLvfnVjngX+c52GYhkoSh/PV03/zrVdhc1T5g
XGNBKNFmGix+Yh7Qr0TJsEpEUj1dbC44lfoXFhQwgQCQistBqAz7M5tRrYubmsi3
YihntLWAgVC+l5NNsupShFwNrg2S3UbeROb2RFJzcHDjyGTaIalZVDz3an/FE9/W
U8LrYQSrKysust2LvLL1yIAYyBm30GGFst4Jq5WYPPqLv4O3z09uQHzrbd4Qgrwv
oA6yN0uUf4l/I4m4hV5iWWWg1WM/WC58hCzlwz0yAh+YRJZ1QSW2dvqDGJcfSpXL
AIKThFkPTJzOTuunOuYUW5LvSv4Ztb5JCB0bMQW3Rj2zmbk/NrewZXkXBxaGrxRr
RMz0b3Mqhz+R1nFWHrmD39E3yU2W0Kt+rD4smAOshUK53ZudxJz64SFndahwImws
muCfTwYN1iORJBm2W8HcPcgqBscXVVPrGlQv31vDId30jUGBI+esra8fzjDR574l
17NLzWSnqEO8iNwaBddFvL51YDJ/gq+PnHKe9iwxqFX1fewRy6OgENLmWQU7t4ji
7d4HUQJWvBRH5WGOH2qOj3vBZiQBwk8knAsSwirrsSne9KDNlc0Wr3Brsp0u2DqO
zzcKmou6P9MhZRs5LkqBzqPvlGYhi0PJW1UKrKYYfRtV1UEzO9E+tIe5F8ZDd/wN
vHLdP72G6sjDV4/hIjmT8wrgYJX3K5jrJoBaVEV5h4aQmOL8fo1a0Txfz8MeMSKu
6uxQh/VRUPf/Qvy4ONqY3xnii/D9ssR4s9qKkwws3xBCwQEXYbVFPz3OU8WRnWUd
sElQsUbFIrM8SbG3fW9PdO72Dm7zeFYwMCbF4KdF7WdOp6KfWpo/PkPfhPG7/Ggp
wpSI98DP+MSfUbqXJPmE+mlVPdX3z+huiOG068OiS6GTybpR+UDtd/ilrsUYvcGy
rPOwCZ+id7k9sH05yiVFQpuE8GYIxLh3DLxG8B/PbNpDhDZ00/gOb5td/06G9Ds2
eZ2pLxKVvcz3n1KtZLlbOryeFOlECabHx14G19Z0NNESYveU8uV/0wQRsrAUvLeI
gZkbcOKKtwkNPZDpJuZY3iDrrlke5r2Eyrjugxw/mS4TYuXK/SlYGzG7EPcGAqPk
k53GmT4xpu5Qr/WeWel8IeoYCTto3irPppRN/YHZDXsdEyMYH3mxcP+Z1NmfRfPc
KERBgqxuh1NWZnln7D3It8Au4aHMKaKqox5G3QzuHWeOyEyL6um9dNUpllfe0m1S
BFMGrmfDKsJmKwXcS2m8vLOHH/238t5qTCVuDaw0OYK77eHtPJCOYgbocMz9E5Uj
Wgdk5FXPMQvhjgEX6gnbXyFlf7yd/8Owu6KzJJjhk4eJSeCM8aH+PJkRu2zw6fEV
FlslWyXpfznDs79KVXYVPR8pMZSXOihsW/bPCWpkQKda5H5zzKEFdkPggVAk/gM8
lHkBTz3SfVuKgpI/EJIR5wCSGH3vZl+XLTS52K99nRSzFQMWsIH+3ahvEKaWSVAH
gy1mEh5MpWPztLt0X1y18UKRMBCxlWMgRN2mj1i4glTdrP86YRpXGgirc7n2MtDe
Phu7HKdXrqt0mHEKjLbEHgOnU6VOA+HJmG1/Xm1B5LVQiLAZA6fyXB+dzzGHZuyO
3RdA/80dzfBEj0VOWQ328FUBJINWvpX28Dnt0N/NH84K08BGtxWkk0cyZGwHIfMq
eIO0icbJVWKPZvAqUdTvCv5eB8y/YIOcNP/WYKqi1HKF4ONxkIraEHhMLPl7q94S
+7mnXjmkiYiT5BrBWnL4fSKz18x7eQYpqwzZ7ut03hw3ZAQ2MXhTMyoLiwvCrSlD
yDN48NCpZJf43HCV0yza8W5Qga6zB/OYGerXdX0E5f2Fz2veVyFR0cJFznKQ2/Tf
HQfGqL6zQsPyBCMcWjFIQh7qaZa4FRA65qnmLSGJ8g4jnga+A2kpFTEb4/hJkTEu
JkNxyMmFbfBA8TAC9XXGl/lflWrql2ubpT1zrJKj7Gy1G7iMu1Em47VAz1Q5S0N3
4iHsH9XLClIF9HymHg8vtIkGPYc/vXRY5dP0UMKya+oSBVhjCn7ue9XwuoOoGRRW
RLFotynMUaeHTnilkgIpz6QYSEINGbZYy1SBTMGHQa75vAL2/ntPUzwk7UxXQxrB
g7wi12umUSynRh1wA7nMRmhpQjwqWnV2Fv6u3qumab2V+8ABMLbMewJiYmonJdo5
0n35zq5Z2AL7zJPZyvkn/Bez5ds5HATbazuhT0VD0Z8GCe/cNYt3OeJH8KIlswEY
pX+kQDfa7aB4Qk0iy4emTeMRSJzgcoU8sQRfg80eP1D7uZ8i+cqxMkvUkCNZfon6
wAulYN1nyG3+XCA4wB1e0YPL2PblsRxdLOPxtyBTdZjcX1rP3Ticfdb8huNfPqCe
Q82clo6sH9BpbP2z1L9BQR7cUa8D4OU9OmNNvs/WS3kL0otrwn0EiTPjv5hclg/9
O7kCZWu83RGwrw+4Rzl28dQYGml2HuKtzqmkVRI6eRb8m6dQHWWj4s3CmvdIicHJ
mF9PT2L3vuBbBjdeei86U07uZ69v0ziwbyS/GXknrCWvJlJZWr6h/mHtS9zj3j2x
tSMtODDVMTnmQeNCBi5g38wAdfl7JlYtCPzczUaMzRqYeJ4E/X8pjk+cXX1qUKCe
mMP/zl9rmgDFj6ILHbq6KKArSuo8MSxh/0EECPZRNIup+d48FIoe197WehmUobHW
+IKIKtFboQXmtxAOgjufxxPf87NZyQ91LL+07q3a8zX33PDn3G+UvLOqzEeVgKYM
kqGyqfcTl6ht8myKB+n3cdwAXoKSZV+OOgpJd99cB6kxKFxkS5CVZdg4kdnVChbR
VtgtrayJyO0I81KL91rRUVS9d8Y7oypqi3Mxf8TSOd90asQJvXvKpmAAnK+SzLkh
PjLHPUfqONBZ0PpJhOfI90JdfAAlMwIuPqbaLaxhroz+EjmYN2tvGXafD8fIHTZC
yVjSZ2zUTLMyIQCJ+vZdXM/pesvbB/mAgWnrpAtugASx/5qOyYsCi8GPa+r9STYY
y+g7SBCw6DiNh0LtNHIJ7k+M7oMc8M7fv+agjLh2gOjD1G2y6A/IQHyzHYZJK3qJ
fNitYBO97BPfe9licNnBgjPKDLK9ngapt2zuQHBUtbdvOibEMsuGCr9YPh9e6Zdi
4QFd5xw3aeFy5Ja+61h91ktndnM8RidXEro7FuULTzTVc9zm6DX6tacjhV1PYjbg
PN//g2MStqbLmmTjshmO03lliORyHPO6ntBiLAXkkYWCGYBTEhn7QmnDFegi2o5g
IJMHWJhqsTV8HycJAyGZhdEI/68EBXV5WdirQ53l7u5jHSpx926BLjFMxD8JH+sB
D20G1DYKwkeRO/3j+uqLUSGAgkd0FGVFAFFmdjpe9/jceXZEIz/ticKwAyPqn6ET
J18tHEZGiU3fEWLvyi1WO7NgD4o5QHTJw/4k+9ao5Bu3A8VMI6wXp/RyAgLu0PX2
mws77zFeSakyQoc/g5cahPqa2z6/A30sVPFc2vvR++fVbq8VbhDxkItq5DaTEmuf
xpkM4mraJxxSC7qvH4hk4iQb1bkhsQV28+gGbVPNv26ahcPCXb4PnXVQzLrQJvDl
v3B0mY7An7Idcc7cpPGCphSFE2F3C0Q5UXv2t0mdg2YBERV0Dh+ks3jcRsmSGMij
VPmDQL6/QxY71p+6rOPAizXj8hWtRxNzApxrcKrOmc9tyzWycl1b1w/udNV2ie88
HLhwHGw+ASiyhykbtWrRxgQJZuc2PgYVaHZehwupKCso8stxZ+QVvqR09xmhGpGj
IYfhyWicqJjwjgm8404MEjjGQ9xLBHR0Pf4VQRsCtUoUIWvIc+xGvX1HlaMW0Xgn
0LwGi17LiVB//LU/qWiLhHc/N2V48DiQLnl5vRii5ooTkbHk58BvCFjStbKkiRVz
10FUcDnhkxV95l0a0BRVDJzrRAf49MWh6mq6qp+k5t/FrmXKce+ykkSiKwKj6vrw
iwaRhqGD3oV9zqjWELMCKQ6uASdGolb47RxdYqGX59ztTI/v8VaZBYgzKn3YnPkx
OQNmK/JaMrYUexf0Iay1ERKCtCgunt222d837UD+oILeYlcyqZ62cd1tYrt3qAEC
wxi15Wl3RaU89H0i/azVEX2iRqi6EIIPYAD5gMU7OimmNstC198vi43eDZJyIBlq
Q/R+DMIJLFWi7C44ZQ/4wczBKm+2+oHbcWAk/YMyp0U4qWXzA9ltEhQoOa1dONA6
Nchw22KOJYqE9/SxGIBLc9Q+nleB33xZjGPgVxc6G5Z3X7sI/vdN8DNbhUjX62bb
wytEzlDUeaZK3dKhg5QnfkW46pDMKPsSR4Yr+tl6YwPZ9FQnShV6DwFhX0DHmxWm
Esu3RBSIibRo7JJpIQsQXlZclDsFzysPKORDrvbEu+No2dZXG67lutY8n1Qv/2GE
aVtz8CqHZvWLBQMlubhdgxDgBR0wtamqVxbh/OFTTKz2sU8/fL0T/DgyZ9npZGFl
OLqdeJxNhbzex69+v1SDH8avL+ChEQ+Y+cRaf26Od2OqvHBm+IetyWeKq9rDOM1r
TOIihPPQxBfxqLSST7jlo4DMmonIcdWaTg8ZblcESm1hyYQ+n+BrwHXQkQVrfniI
vNz/Hcy8QOzBbnAhlUNavKuhYqZwky3PAziwfJMVlApNzmAeov4tjxswMubwt4WI
FZ7pJSQagEJ3Or22UbhruO8fEtb9eeSwNEfFCzjpl93hb2WkKcZgCqJXVDXiPqBK
LUgozEVf+Iswt+vKXIkUhdGY1lgg3pW1E6p48B4JRGnm7qInBCsCXwwbKe0otyXK
c8HCgof0gKna6Z01Xphvxb4iOnfeHA+GyEd6yWXdTiL434BegcmR4acaJMGYxh6x
AYBDwoilt31d61OIJqBHF8GkEEaUIfxtseXD054s1+dq5WxivT+ctJHkjjf3E6+D
qU1+y3X6Q3uknh7JIFfXd2sQGL4SAPturWbhNw+vZp2ZV13ISOJ7PYeCppnWPTzv
mOECRSv+ypB0B8xisH84voEbvshKyGhNvaNVfoq3HlvgtE754KMo9JDy8m/HJOwX
Yptz4twm1jPNtPMKtPbWoD20TK69mn7VnVXbcttSA8UHPec7I4V/us7sWeSi5pEl
kDQsMF8DYOW4mvrvKUDyX5DOk+0cLa6ahsT97jTgpZvBRf1Fc3I1TfhaFagxFEtR
VIs0FHU8+Bc93+F7dtHBnd+G4myYylM9BpkVQJdP+BQoGWBHdVS75PoK8PytOlJ3
JmuZQK0FIlXf/ybDVljVixSlJkaABieXhMsd0maX+HZKxNOEczX58RzOd91TpZn/
U6X770OcIKHbviVwXaOi5xkPgOZ2JY7w8gmgYvlOxmJhUWXtG/T9or0ItAOK8Xiz
lwzt2ZzXP/7OfC8IlaLDdboHq/DHZSuhYbVvh7Ezz1jP90rp2U3OkorcCHZ5a0Bo
oS13hHtLN6px/XU6ilP34Sq19jWcvTQRL2O3T7uUaO516hnhMgyDrTKFGRf70KoG
eutWeh1LWxVvYfBqzyxIff7AvfjzwzTPLt/ZoLFHWrwU4TLL92qsjo1E3wxqonGN
ziCdzKwy+7DsD0u+rRdup5wlOhsvX3CSD+gaZ3WudqwnkqdXARWK/rAHI+gOVn0a
14VW9qlFufbvQoA2mmC+ukQPcCIEGROyPbz5kgG50tDcHDbuJ99CJibK6z4dgSWS
TKYLeWIfqAix5F88qtTJagLHw8AC9OOntnXiRC1lptS2oobYF+ojwK7VnBn2VQMH
UVKBPq6EBT+dUNgv8VScwCEjAjczCNuW9RgaolB6J+XARLsbdK9q0Ult8oTM7KCZ
MqmVz5LMwH1sZsSS5eHBm/4wRF5SN7cgLnYeQP/k+tC7RoKsupdPfxubWLY9AbvI
q65bd05XN9hFRcVQiuHPJSygrbZp4R3Ize/Aq40fvYOzSkkCQIg+lu+XPEsva/Cr
rGGiWZ57D5DqHBD931Q/6fHmLAQ06o2XF0IParlTkM7bu8MJNl3nvhEaC5SiNv7L
tVxBt3MVmgBFq/T5xikOadWGxlhZdLNR/uUUvCwanby78yU1lZQR4+KGPTRJsHw0
UEu7h3SQ9m6kCPrKYMsRpd0l19iKZM4cS2I/X2U2tHwhRk5U4f9XxMpSv/9KeNv3
hqoEApve+3agR6U1AFki9YwFBM5bvClvV577xHHxY9YivchQxUqgiRSGY8U5bICb
HJRZhEQb8EvkG1CqjE5FU66balajXfDvxcMviaPSBMpxeUExn3GhU6dXjrRAF0KZ
YViZGzCtqrrQ6wS4ZZazCriGo6BBEzRFl13fKTLxZYApwTzI/8SfBKsjIBwW74ac
Kuu58o1m2rkrmH5GuTai8IADgIrMGMXFvoiN9fucD/dzQCAU7fyb+C6P8hOvOriA
j7WCqEL4c2CE2ZeWU0r2qtXjA4sNWnBe1yq0viQ4j1RULmf9CAPpm/12mH7HxYD2
fJcWh/X0mQt4/5/ip1C6BRxiSCd+qI5GsD5x3aG9RZcK03BMhdn9FmLEhlkIfnpP
lH8gLRyUNo47SFPSEcBU16U89mJpjja67nu4op5LRxVoKtOyKuxLQE8tQp+Lq8/q
GFaP9lrz7Ys9+Qk0YDDBGFr37T2RDVE+r3Wvpm7vefPqAwF1i4oiJfvxYU+7bN4U
8hKd/RfXW0VlfvSclkH13af2l3GkQaQnZI2q7DA6kylnvqa1mI/T3ZiD4USRDe7Z
FmAYBlpIK6k/svVEJXRu66SnqMqxO6qPkrsuWlHxRkzTnibM3R9E0yG59izaorO1
reQa9ZB53IoEeDLYB+cj/fqSuIJGbneIITlzBtg6SUXa/NtVub0Q4TmPREDk2Dpn
UEai8HR9lkoyk4NR/PlxPtVj5JNr/RDOJtROHojt2ZfZWfqSNkp1nS9pUmnKrgeR
wgYuO4ItDYLAxlkC1sH1EBp7G2R0zHPyqYA4aKtmlk44tne03cTk148shjaTLqCe
msAGc4alTD3Qij3TwxLvcBpJgNiyjnuL/h0T6JcPnXjYFRdZK41GBymwYSwGkQF9
jKEqmgHpcRlKQj7TRoyyuMcwjO5vUYwqD8IH12ogQ+Q+LhKkdWSBG4dkq+RnuGi+
5ywlqbAOTQUqLQnXQYop35W+sUEtiQymPEYyfzus7C292hIUqPSBzgNKwap2L++s
gHp9RNBnWCUK7BxLhT7cou1YtWjt/JQ1fa2BTX7peUkwV5UEP86XQxGu9y1255y0
Psct20pgbGA+BumQzEPCPVt3Z3dxfzwwpWNXEldkl9UjdXZlHzBgAcucsN5+PGv8
JxINSU3xOCiz5nL42BoJ90eipwAWK343kza09RPHFxf3pm8CFEsuzT+vsAhlk+Mo
h9gWbC0nPZXr9LDpenz2bPbIS9mu4k/aoVDiN82komi1JGkjkVaAM61/KA3Or8/R
HuS8unPGbI/6TrneiWbX41pA5jbBdUaTAcWv57mQGccSWryPdmZCSdxDK1i90W9M
wYLX0tRWOQgVfmSSDydlC19a1qC9x335mbcPbMRKL6ycrkWg6XBGc0cuSxTEjswh
MqQAb1YFVxkzIh1mD55sfqXZt9RNIkkSce8fOk3C046sRDtT2XVmV3Pxu6ISARwO
tbydNfJoRtut3Hs0MlgQPlr0lwspB9R5FKkMBltljVyZLkQeuoH1TfgP6dQTisjt
CtfRATuRcFvnrvEQ5io/T7bTyS12wx05sCsfptYJmyQH1yg+D6s6ZjGJH7sMCQfU
/f5r+lol6BUjLHeq2GeOyEXPZsg34YfHqtUSG5L4RliV3itye0I6vq1WW4ZjEJ2U
zVeKqqwPq61VbFb3J5pnzpOWSM1nX5tWi8NSH7r+jnaHW42IORw8odg+21J9/+Sx
4wS/cYgpE+HNBHm5uaF76s5JGgQh6cciSAQrhw/A/PNaO4QOH7e19Bbd6UpRPNjH
vhYGif0bHoGCD2pdh22HaT9UKvpwollNHXMeh7C2HBKs0B2jyeu7oRVKQ0UQZ8Yy
bUODpscSRMIMyjii9xEyi0i9bj+X1K8o7u8/ILa2XmUXfyLOfMvd8ZUk2r/4jLDX
dyu+GVXf5ti5NMDkK+mHH4hy5gUzM1US5aPHT0ekHwnq1hlq+kNRZy08eV7GmqiA
keOJX5NYrREjL2fiPsV5Wj1x/f05nNveZ/di/K1i0svLSQG3RPvPgiRc4YqenvNU
JvxnsrvYPf5pp34anDzMZs6wPw5FsRLL4szBSVC5uO6nAJwpgaLQPW3OwFTbVTEt
aFbJRvpfuqkB7yuu7Il5CPpSc63XC6hVP8RqVwIfs4IvLyYjXrb0KSr6SKHAkfX/
kKtY2/em86LVU24xVUhbmJUmmsrCdENtoMLXWIi7r/Wu/RdOnQ+KsvwT94I0s5Nv
oCnkdcSiqiZXLwoi9y6Rb/YdhyHh1TUvPSz6GiAbGi9xLYYIxwL3Hf8Jgy3GsMEY
VOQu/232vSKXepqm8gES8MkKJL3N9K02GzoY+vHb9fMS/hUYl6r21ERJ+bz8jlip
hddN0+EuTKSiKHZnwMV9cAKe4u8NFTRalUCTMsOrV6kPT99qM0UFcmeAF1qLvFoo
HhgmiDZDTTomXSI4Lq7ASliboT1JduXNahQXXisdEaXuVKEnM/fGSPuG02MIW5uA
TivJpjH8Ax/QJnmTI+OwCDb++WLrEH4mU8S/Ydhf8yD/7qPjB6oxFbYOzZ22sFlC
632QX86tVLu3cu2me6Z4S9KNGLr6Mkes+mATMxQM8PiaF7pCXohl21xmK4JwUy2M
BfQSNMQ+6Fn8OtP9iHK5DsfCuhxCCi1kjUMSl9fM/wunYn3VqoOuMFiCI2ZuOYnl
V+AiVgjarU9aJnH/K2b2KiPDDMvpmIciC9E+1zxhVdjw2MArkRs7krbVeADwJaCd
GNiV7Hh6VqR1KXAQsndlM9OMFMQByRvd3xTi+micmoGwevdoqU4bVMv8PesQUyPV
Tp2UzM4oP0fa7atzBn2wwJShQfyqL9HYru+wE1hGXRlHyvEZ3F4lfju+WEsRcOv0
VYt0HibisYN/Pyvu9NH8BuEH1HZFWFWUzf9IXLcC3lV/X2kjjtYguv5LXPOU5eeU
1hYBPmg2M5EofHPBb7S1q3XYUzQbbKNCLMcdYkn9EDhCVYLRmjMN0R6ZSgHA6Mlt
CdEA0PV5xm1sOi5U8wKuKqY8ev6jQVMf2CWpkptMjGti/Pcbvw0LjBFCL5jspmEf
ErUyvaFINTnKD3WwEPZByaj0pw30eFXltBQ+zu5TSafzLW48uDo5WMTiVvjh/Zzn
1EyADky5scmm6WX8VbyHnMN+stECHwwgrtDR1KWN6Iwv3/DGyJzzYSvMJMu3YC9/
18ZkW5nhsbCNhs1nhITJEq+CwVm6O2Vu5N9WxOR4QOBl1tqTDo29ZcWmNxJwORwo
vZd6Md5/mx35eL7hdrD8F4WX3QIYGEFHW1wNGDUBXvsYmukj2GOQAneRNrqq3W/7
NEgQAWPGU80xrB1J5gh5yi9vsyekOCnRNGx12MY0bTpmu0QO2UvVpH03t6PUZJrd
XVoZ50qdodycxWNXeO3D4FG4Kfo/pG1sUPHwti7Og8Ffdg8NfARS8M85c/uJtGYi
NM0c36FP6sUSIQa0/P2Dipk57fGGJjGcPxXvqM8kFbGWT04wi+GglUULPVd1tPAw
Q8h2bmFS3osQPPK2VnYp9UP8TreniDAq9pb3WAuLrfi0mO8hUQKeLGpk6gO6va1F
jrcveB3xguU+WZimhyJL6+lr1aE6MMEQa4brPDaHqwvh4b0hb3IjI94YCrf+FTdN
suAwxttAyemuFQW9TegxPNhBNQalOIOFfxNE9YYAuQrm10ms26UpCkV5lY40R/+T
m2UhyjLZcvyjJg90jZ7lU4IaMdpeMXf1iMUQtP0xH02jFriCOayJbBcPLnfDYesD
cS+ALXFb0n/4HbiRPuHVccMkL+RL7LkvcOW4aqc0JTqz5bCkWrYPzCZaglkc5dhg
vSEtAp/kclwJnsBOxd1TJ7fEcx9KLGlxFo9CSrxl3WX3hOu6J1PMS+hZ5Gu7IEuD
InBlQdjTHZN2MXxWNjQa4QKueIxVznUt6ehj6fHbnk3yu/t0Uq5YJkc8PdtTEGaZ
yT53NR5GG/Zs1XFm+iDu+zbKmgaL1hT88fhcVcgSFv7Ssli4QHt4nLRT4Fh+dzOd
XnYy2ocpL3fvn+9bxTjsoslbiP8RU9perk1VOn5EH/cTkhnLPmNVnutp0VHF/iPD
6ulW5wTj7x5lIgu5TbHok/Ftucx48j/QAXacIwdsF6AxOQSPiAyZpUmP62V17zqQ
dtla+sCBEzoYDTMupNAro7LHC1EOAZIL9V4FnkIZRg+adrg5bun/TRgd8qt1M2Fr
ollCUJLu8bJWDfNrY6k2KcA/iZHq0GxQQjPGi6wVQ1/aBVhkgSIPFV9Ynfj1O9hD
ETrwIC9PApOcVu82CZugYkHw+fIlD/dCbblZsXoeOlSR9Ee069IFU1o5oR0MP9u/
agTaoMp0ZEoWl2+x2CiH/A0A1CxCJzv5THFP3NucPWhUhIAHHfB3wmxuwnMPexBE
w22T4CPDeVoe5wag62fM54FtvehTxMzr9t/61bYEqf9s1BDFl3A5Yekn2MpFwfjy
G0XIr9D02y1fbsSWXBesxQTHlInPdvSOXcGHjNpY0jGISGOf3SV8w0wUDdTdH0qv
Pxn8wbtYXR1GWPEOb/tOrS661AvNyCiI9Vh1H5SX2mVCkUq1L87Of/b2J5Bf9oa/
X99IJrbBeKIbiSRWMFeqC+zIX0tbywf/+NNG5xhw/eprdJao2yxbGUPF200j0rNc
zqDbGz/kSrxpRwF0qUk564uVnVDSKNOKMq1x7he79i0l+tiDzVsVrSkO0VFwD+o8
z3kKShtBzQLD5avbA02crO688kGWEHPPBqPxVeJEvTR+pSm2zDXGS/Q2LEOrsnSY
FkjVEi9oMyFiyGAg/qiEc1Ew8CK9QzYkKe6lcZkItQvAPwSNPj1ci92CVBzmUm2f
5BPXGiQgOGOnUbGwNfU3DhOQTGPvUSKDQY9HslgJOoHYlDQRVc9Yihn8gWhgOUIQ
vVbeOsUmveEbJ+d9rKyteL+NtKAuwkX/4SQIr1ib/S552HBhctGTQ3pc3j922Aya
xcWAdzNMUE1Alxl7fNB3YO5FO/LDo8TZ3/yDCcfKCx8oyaOD26pKWZ6ZjCfMf4NH
FA6PiRkiM6ft3UnWqzHsTz4K+I4Tyd7W7ti4CKuR35q6/yFy8R5UfoLbtTaete8h
9GLgSMjI/cCZIOUFCBtcDjOZl1G220zxREuGrsA9Hfe6D+VZhxrCinEMZpxUwZRY
ILg8Dkq3GjrgMmc5+bWEU67UO31M/31iMOiuTF41KjH7GOrthf0Y5yXnxQYfk+L/
9yiC5j9YmrYLighL6mjPQDKOKC/lccPXA5yKDPv0UbdjVGWjAoqCSjT7i8s3RytU
byZJgv8LuxDUYcv7dOv9PZ+51yB6Fnt6/fioNXSgJ3KfD1T/ibqe1i42Ho25x28Q
UN6tGT8IyZ+Q4DlDg1kRPH+AI0M1KDpZoVrX33f2ReKfsOWsJA+UBGpojYB45wsF
Wi+J1BuqJkI5JMOt2le0d2EapwrGUfeVW5AZQfnUKfWLNLkYckwWWb5VSrbkQnwk
26zUgPsJ5WJg1wP5Iy5/KGe0Or4H6eM7XidzibjgHGAOrAbX4va6V7O1eYWIw7dL
Jyp/MBorI13+2zNudk4s1Kpppz+nxDOVzdLtwMlOguV/CDLq8V1rS7N8qM8pt09F
Rq8WB4pt7W/Sz7VfjQy7n6XKhWmbYwrkcIz3MnmLvbFOxW6yRz2hlEr2kd47WSkj
KEM+BCojVMBqorCHD/swlTEemMT+6fedMqMy9Ar9znCyWLCYVPCGftLrZ9zKP1f/
CnaWhq6LS/AAudh2c1G7vb93uItxAHB51IEjSS0r6rbZOjugfh3cTBpBm1DpbubH
orhniORTdJUwcKWDS4gPkWGalPPZjwv4E8wRokvIHt/957mQUshS9lFzIN0j++Lu
SwsjbPkbCrKNe/6ZPv6Nw7IP7ieCjP+DbKdd3eoYDVC7FFwjHf3XPuWXqIpYn58L
D65l1bARPWTXloArtlU0x1d5rW79O5rOPEzMSkAZ2EKi9ksuXVIX97ykBDgXw4+D
v8pMEUQI4tmYr579KIFCBXtrDF2q7Ajf2uXz1Md5SVBrxed5H/aaqWweoJk8Ones
/9QrmMH64rh5kphwFJvZEjlV1mECvxeLo2Grhvw+mrqtKDK9JGJpFBowHPRtPwl7
VGbASDKdkdVLgf3YNmE0wFI2Ipga0PPKtwpyGyk36fZAxRKCac+JmsGSqcQ+Hxz1
SCqcXaDfxMV1pa9/aZI+8jbNXJ2CWaaeKySO7n7+7LVc+rP0UbwvL9I62WwF0SBX
2YcEurevV44j7KHDtgQYdBMt+k67TsNKQBwGzDGsPRUB8esooXSqYhX4Ez4R4vAY
1bFTPkuvnOMk/CqJoNtwtUN8arV1ts8GeMSSFtpPSpDvCx+p0CpPKe2dYEU6ynLz
1hljdsQ62SUeTgumJ2rFYkhkkoUxikSSEwVYcZsdaHnHJrdVtsArBk0NiJizKz3a
r+0zTw9M+SDuDqHBv3CtGj8QQqJ17dC1AZTTL0fbd/K2dSJVd3yY8YnhS03DWwpn
rOc2T5qdcTjXhVSl6BCUUe+9a0u19sxkQva/t9GeS+5owzL8fT9b2mRE/T+hMsiG
ZBZ/cO2a41OyXnApu0kO4EElp4g98Mi7P7ZbPUZM9ezlIpw6xfR00SYCYntxlcGS
WICSbOdmzoTvnCiWigyJXcMW6Wasvkm1t8OgkZyqHsJJqh57hMvPZobvrDIFwvWr
gTxeWqxAHyR/GjzyRtUlEj13WVAjvH1lwNdt3KnX3170/VFMYkysu+JALdR6s6ef
JCvel15eT3IeG3iAMni5YWceu/bSLZyvadzq3CKr28+XVsd3nzifWy6rwVqTk2+h
q0hgRfc+3ZF/pm46qRazsjK+bcQ44l7IWDl7fSb7Yqre7gKrI4n3h+UpTXBv0hpE
qBbgyOtKscdDeKxpJE0CuEp0/bRW6THJ5AdrPIZlqVWSbrHwB9+8QV40bcb7nkVA
jsn9GXaElJIJV0RV2AlM435YF1tGY1y4nE1zQ4E6fpRJ1BqN4lTGaGiwEIx0aqvx
vnFxvNw8sxYp6dF/+KkIoCc83z5Q1T2Z1wWyLUPF2RAsgOa+/pLcJLojd1I6nq4C
qNGGrApILwAKMOulw1RZOD2vbxyc/GqaRoV+YEB+Dy8jml37VvH/iPgGorogFSzD
tbDc93WCWdtl7X5PAthnGjBYJuSOmbKRhj4gXfeTvJJxEkX36lHdhsCzDUhigkqd
RcWai8DYyADlM57PdBlApWMfL1dzJfuOpT4wUBhKXf8fZ+tKZMtoJ1TrZmclwR9e
8EEWdYCRMJ9RRT/J7GYD2XkHxLiNILli8KLZzSPrjNuygJgZsrqu98lkGxznC6gT
3f+XY8gxioQecicj2pAJE6a/VU7uxrh+adAGmdkEyJtSlZ989IbyJ7Fy33AzzhMB
krBJGTcAdO8TgGuA0kbEcV2/tLuHc7lZ78GXpOeTVSRcZb81JpVLd3SUxXsts2ds
B/KnZd8q3SqWSrGEqICEq1/YTRJqN3vA6kZwBnfOJnXC/A4J30JqU44AYQoiGf19
WVD1Dcfo1Bf1pk+pRavDYKnkOj1cdDGEmIT09a9EM41KwsvbtYCDuxOOdgYlpUhs
G7/9JSgy9KKQvEpOWLJGoeF5rgmcsTvPDbS8HPcg/jbyMM36hGvmkO/APxvlIf5l
AWCnujA+3Wr7h08oUKsd8ELMzOuabxZCzlmWF5afLc0h/7TtTXtdWprHa2LJMYc0
rpSIyfgl6f+9TTQsLgLRbB5DYWBkPeCRRMlQNKhtNyv9LhwHX/L47DWBQ2x2Sjrn
jQN6hmkSVzGqCazNC9GDkA6fPr2GcIuzyHODrpOsHs2GepZRS685pOVpYI+k5GVx
+z6FIvl/Q0MOnFBbyNiKhzpN2BYPRFHYPorjcfVkH4TKXHZLhE3KaOzqgqVCPoZf
hiALCW3OLA2ZSbWLbDMia6lG+TjloQ6q7EWDfPDpcwTvgWPOD5j2I1A2EegpMQCy
PeF5w4l9n5l1kXMMgEqPZ736dlexka5kpM0NXA+kIkp0Df/8mSNnX8ea+e1eo72L
4jg9OnEtJYjaNdkV3MO5g1Kcwvsdm+V5ebu8+T/mdJTkGW4Ojsyplqs8BSDWPKdN
JvD2BxB1SweQUgek6Ht7FQH06atJrV40KcCF15jT9BSQLCBldDV25TO3/CojekF7
GVWmIx6zGLBzaxkcbz5GIG3KP3s9LV0IO1FB8qnH6nSWnEFygbVSGr3PyfIXbWDo
Q/p5/eRpCid2ZiVMXe3q2VlLG4sRMnvgKzL+W8NzMwukl6v5XrrkDpJiHvtDLy8z
FKaogL1mo83V73pey8+6pkp+KbX6xbMXHaY7bMkZ4BRPQWAyly59K3qs68txnpnU
S7HMw4vD879Ypjc9dXrg+JajChbsPDkhkvfv7G5SjGN7GzXGXnMwsrz7b4Nrqdei
nYw6SR9DlClhND2wfo6hp2L2fMJSQLAMcwHTDZN/W0S/yI3q063BXpr9yR6OpM/T
9rT55GwEWMFdx+fixGxcrHwExDWiiMcdPnCOCPxTOpkHJXNdF983W7VAwAG9fbVj
3FZdzNmJZQpdnUpsZdJGOjopTclFcNegIKdONJeL/jSZxwr5YuIRULDSlEsUcBQA
YgRG4EU3MuX6AK2b5rvmbg5F1aA2yVqv1xorOROwPaHqMZKPAbbYzMu0ItQI8kAI
1bXU4MiZ2XSJYTxk0PGPyjFucrpzrfXgPUpMclfMJ+rDJz3/7BatuhuTiszleWBK
Rp16DZpK31skyo67O+tFlmiOA8rPJoHX8xjHZF7bifkuCPwmhxctlEf8A97p6zCu
T3Qe0SsK3i33lLYOe2OUArfjSyGy44rxvWS/vRW/KHNQOvpfWgwSc8/SH7h4ilXM
52ok2ek+S8wXtcLDQAlmVhIFR7VUaNKTqlOYcPDGp6N0cIXXvQoQa4P66JE5Gyga
+fpyyjMx2GwTVOE2D094R/o56rewnGaUalf5FP9yoJsQdxoiceG+ddC6kicHzm8R
V9QaD5pI6KRtlsO0xprxTu9Yx3XOJabI7Z8Bqx/sQHTHhceiOJC3LU/Wszzx+RkD
/BPEkRaRPKTvKKIgmOOuOBVKTgJQsv4+p7qvlzfPejeAc9ix+ObTrpG4SlbBcx0Y
V4XROGiVMBKbPZN7+/gRsASchYs9Zm9KMNlmUyGg8ZXA1x7KJzmucwrnlUIsYxv2
/Wogvgy5klReBNRhsGdOZiNxXipQ/SUUnuMPn8z2Pys+1FSYBQDtrRXZchB8MzG1
l8Pdy6mn8wd7eZJwfsUuOJ3tJq8D/DylM0lUuYwp0hhumsmHTh4/X4YwC0xYdOZY
Y93EEiaGBMLGgfvrFalYcW/5hVpS1h1bGOeKRQxmPKm3pwpb+4ZgZcvo4B1pEQBR
KYmSXH8Lrc1NdGXw0t2pVxFlY7MweC0g5hSSGfsAP7cqshST4GQ8mV0FC/l+aDkK
JsJsCc8cbCYFmtB/XW2/1xIQJ+CkuWs1V+mB65eF9koXDfjJh3dC77TaPijwV0aR
4w4XVsprL2fD4Atz5NUHjHBw3rTwbqzujLRXtm69f948KSo10dIO+3LTXK5JCO0l
DKe71vpCIq2FJejegiaVdowe6kI+G1SA+6NwAvz9BAtpcqIqfG1w7zssvL+QsPWx
a34asIiLT+eeIctG0rSM0a6UamvvjlIyXOL2DuWGyL9r0XqlY18M9J/54GcZZUGi
ks6YCwiA9OdhSkimB2t724XGVaS3bSWUzSMKy95McF4xYWKZHJmEt6Xcfljwcrrp
OERDvh1/X2xLYUME8/EwzThLeSe9JMhcEDHTZU6VjJyeTQycNZggr8QgmaxU2ylO
OXOJWwSKMfg14GtB3+Z7o6RbB5kgdNvp6FCfYu1SR++blzvBb3uznZ3/7jX8Djct
PbtIqWFhlFQUb5Y6YRT7QS6D47XiZm2aY2QkT1Obvub7x/etUKzjRZo2dHy12Gnn
VYgDVFwX/kBNjKgawa6E7Pxx+lprWqKY8v2eWSD0zYlCCMPDNOfjhmNep8KCxZ4U
5ZfV4sFh+h3CjMgcV/gi3CGD5zK6ww+5laJx3wzsoYSN6rN+DHuw3UUrAYG2VHKd
Xwi5DYS9Pw7jvt7sZ/mYhri6E+E1VCF2k0cyuTbzZ0sooFrmJvNcfulP3eWIjWw7
NbuhY8f3zWY/c3IbRbs6UhYlQ/XL5L5h3FhocaScz+3ApGRMusupPp707ThnVDGo
Bm6IsE6LKnCZUisdAHwg/emHq0O94C+s2Z0sdrmXd6Ts9VK6o6KM6Alffke8JFeS
yS1pUP1KXaQc8YzdLhIpGcA+WSGWHXsYnUI8sEYXqNmsXBcMsbf/cfXX+9BAERBp
ugyDJQ4DwvWSqBJyo6a54QlSqKuVs1tyv1hfmT28YETIlx6S/FY+9d/4bD37r/kZ
PtHwaox2yXvEiCPy7G5BOmvUmpw3Teki0QJk1ewutr/ULFt6UfXxwvpP4cTNblGd
xaUFj7m36yaPbq3pQHUYu66Nxm7RT972OOOf0cSDFmAhVTqiTE/HY1tu2cgcM26f
4OQBleGMnldir/rBvLBEdD4ETNQfixzIpssdhQ9wAvijgnnvaOkQpXTWMFMg1zRm
/i0sKJ4V5iKZrJme6ZeqZ3EGiyLRf1+S79flWRA7zfsYiDL+GUCyOhaBysv8e8k1
svzx+W5tDZ8vYhjXa5GSP7IIyM8uLgBwbKKJ28fE1d8GD+mjzAKpAN7r1jscvAMa
CIDhfcaszh1obM9yeSqF3TIRF9my0dlmtrvIrb06N5k/Z/y+Kf3ccnqWi4Lrq1GG
hbmYP2zY6W9Hss+Uce+Tn6/4+KeOi6gjV+xLd5yqfXXFAECj4rgLVoCNY/KrR3ej
d4GvGK3UqOdLhkq/jHoE2aCYM70K0VUy1P1e+skneHY+O7zpRmK0/OVX9XmHiZXh
fgxnSiksyKEE7EpZIVzv1MJRsw/bv2sQH2Cwv4awV/PiuKXfaTdBvyBfkeUPADsw
asutUtXTuDGIPCW7++hhTpHtSvHDJp5QixohdljZh+jDNVknUF4VwYQZMfQTj8TF
D3R5/3HZeliG+90cGe+KvlW4L9zOsziZtX4tY2Cwz8k/J9h4Qo8EKyRh/4fyll5p
cEH8LpimtmlR4lejpcQuQZnRh8gRIt27cCn6HVkjy7PZDFI3PTkDMhdQnjOg8ZTi
Z0ohx4bgqYV9P7+4ATvWNqDsmR5ym82ntt9XGhrcyKXI9QaBPEHAR0W6z4fzISxZ
t0d9lxE3e9ZzRqbFi06H9O3nEFNGmhUCMJf5CdKtBjFQQDp4yWpNEEBL0yk52ShU
3v6KlHaHbRg6JoxCwhSdPXWYOJ4ZaogV2dGcx0JFFUcsmljBbmN62R/+BzLjlcDj
7/cG6kjCcXqpd65tY6sSAhlVNzDuzv4efgbIONtl56v3V/ZJgrIV9AoIG2AvqLxx
4IluKGSGiOXs4JT7ScYMMmYHWuZPbp9JH9WzkoSqA47zgxjJYrn80oN6yRMmJc00
YiaEXGAKIs9cyFQjaVEPWMo868SoYr1jjgZRWQt8QuGmntJfXB6oZ2jD9SszXwO3
1/xXNzafhwUKdIweRnXmEaDdXhvTVFoSwxKHYrDQvIeXGK3NYclLD1H9xq3Nfyx9
lOaPbLDP3q0aOUrtvVJXYnK9NZRf6rCG7VGLdU6ZeabKTEnw2tDr8O8uxU2YohNQ
48AgZWRE3p3B5dac3apfz/lHMPf3H4Klh402SOddnxj6HF9LntBldDvUYoO0gkCq
4v1Gg2YFs929JB9U7coV6viMWpm5bPvhcIkN3mQvmLDuvq8vgcPmDwWmubVb7FGs
iP5zNWA+lOd5RXD7+LTZ2SPwdq/uAfa3o7DdFTFW8HGL/NBQTWpXqTFnrYc7pWDf
srx9zRSCrcpOxDscTsUxmDtQtog6WSIvles+ndLPLias2JIQ+3p95zVyzi1WLf+2
wG78RxAZFgr/0FOsIaR5i0SlXzkg1armRuYHOhOXiKHk2bilCyhPkAztYNdrWBhJ
bzz82WmMptQG0Tzqh1ZoxHYuth3Y4qnOETM2B1yCQ38+ornN3kRP7DShwstNfFaM
FvhrxJJ1kq/E0tBtjvwBLRAYFV800qEUY0w1RPLNqBE9jiIjYVc6YijrqRI/hEg5
mPYme0MMr1mtM+9/qoxsoe8dWwiPrDarHzgxdBKOi2c6AR9zV2vjPtt4gxjHeUh1
SNyD5ihpnXqpTJxYRQat/alKalDfd03j5B4E4Tmzvxy2d5AAiACMYWbA1gG6QHkE
p4V4DFUhF10+gypYu7ShTMA4q+RGbMAAcrCBwqpnLfeejBQ/11yi471vV6wo5szw
gH7UGDa4B3Ve4xCq7/1t3M1X5Qfgmat56CqnuNGSsu+lAj7mANQv/1O0/7d6A2Dx
k816lsucCz+qw/Y4m6LHZDgya5WvGPSpa+JCBf38fq+T6HBgPvwEcisSesOPhH3p
pi/BGZ2IGSTxJQtjeu7NmH/tksHal6w6DJNy21sc1N947g/wl7zLTu0akNxw54H/
x7qWw7KM5ypkQ5cEinArlFRlZpAWF/xm4D30385Zm2uFfabwwqG+xV1uqqDTjByf
rXfFdNX/oFzYXlzr+bjcBxx99ELULNjGN2XCalDfIDth6EigFaJFjgLPR2o004h4
rs/9AuX7mrpraDq8IIqC0QM1cFlYv/QDyYRwPOj+TrGOD7bNY08ReUx/bgp99ZzB
tcZhkmYqKfpmtkYOvD3Zpa07IIoGcr+S5Sk2MuyxDM/L9Ui+016SE6Yc2LiUfWAN
Df67pbuEoYkSTLia1IGm3Od21MezvasPmTncPPPwUFjinjBozjl+8HfTcaKrfle/
SiBnePSEwvXMTVf8wKbDnF8Hx+lE+GW3qeit7XCY2klJxdWIroGeA8e9UxUIN68v
DgQIxpb09BKTW7vk9k6kUkH0ARfmHKTw4bkqkHYBmvbwjtNK4V7zhSyDxEJgdg/V
wnidS0L/yNC9yMqU0VCWjQ8dxqT5SbSb27z6ymx1txz/TcFJe6p3kWUmIf/Az8J4
EocDK+mpAjgEn5l3otLK2+SpE5k4L56qmtgSC9j/09SMMGRcoAwJC+NVEqvKxDl+
Lm/D/xUZKNplhy1gLyUzWt9uafv9Hj7G4ozEYwJ0V19Dx8qo8fYYyf5Ns4nB2wn1
0nJm3HIqwNK4Mjvfpu4XqWEYOFB4nswo9sThNmdMEXWelwNm/4nJpqpzIsVTe0sT
54sqxkHc0s8SXXAqYzjtQNv4h0DpTmo35883SAmNspqNUKFMlHSUUQJdwKZuwJjJ
HvzFoTHbBWDqmilR795kSiMYvT2uo+shTtMcHjWFltYCmS5FetAx0iDhZxZjngix
091xes4j2tG6sI3HWg6kDA9fBxuAyhuMPSdAFj6+kfBMZ/gvDwDbVH5HQna4FRZm
uTZMqTnT1cT/mkhiV3egjaXhLKn5ag9H+GggsOTy5Yo76IZZQvXUyQkSnBzQZK0R
CSs7t0fmrmAycgCwQVK0YQfXa2h/Q8+PjrbNSRRM7zksh8HMHSV7sgD4FfFTaM2q
26ASOhLfc+t9Q5zzyjJiDL9B6aSCJd0/lNVhO7YbHmfP8l1tlvF3bNyVD2uActxY
aWwxI03dT0LbC1+QA+tjzQBRKVevwXHefLaDrMtf4Lyh4zvVRKLq4Rklfjw5vjz2
jrHbT/3PeqpG/vgMBjYvWFu7v2gY7cBCvZkDq49/zTphFp7Mig8cSRgGFdZLCcqv
FGH3m9BsRHkaW9BFSe+QYc7Fu74us8sC/IKcOBwwzQCBN+ygzrYezG/vSLIHmHb1
nFuzDLAVEGasUQqXo035CUfJTwE0lVb5muuAMsufVbxL2oCVl65qJ1waSvVtUky9
/+dP+XydebCPqFAIZ2Edr2KOkrItaNwybkAkvRzx+WKxUe7pKUZs7BL9U/W3z+aX
HWNqRJ6C/1MJGOezSoCo9lStwuZCpSEyDeWEjEwiJoESNuuhfMeilPe6yJEXn1Dp
xyGxvl7528w0qTcIj0lroGst9FRbXPKv2KzJ+qK6kF5CqzlaNJxC14BdpZpLYOpM
p36GYFybxLRfxUVlZDq9ak5nCKpOv/QLI5HRB82Z6/BcqhrG5KitsNZwRunJ1Isq
+IB1xquxCcQ9TEHKYvwbUzmsoFEXN3nD2jUc5Wd9HPDq9RRMi7VcU3iVcJB+s6zr
AVX8qN1VwowUWFI+GnVuOb7IIjpAt6lBqsGPvggIN/M2JLTBh86DYnqMg0WX1pFO
aYgr2rx08gSnbbasTOV5cyaJ6kZakuGss5kE91Cb8N4JoSWXOtt9EEOEHF20i9qs
TrGJem2Uk4CidLQGslYVL2twWwAvUk+sJE/BaoB9+eBulY7FFUJIAipsh6w7UlaN
m62CxIf9qgFy+5qQvhPiL1fYnsviCJS3105pi0qJuWUwNPq9fjiAbqdk3l/KiLYN
r4bItJQWTXZ8zKr0GWIZjrc+odSstTPzcxTMOTAfCXUypbnoMZ2hjaPOcD4PKwA2
4Gic28TwtP8r1HHZTzDkxOjg/4X6hjjy6FLle8Y0GX+TI8K/aaIMU3tqFsiw++UY
Q8ukpSSSUQlVMqH1/c7Xb8Uk73OCLGvI+yR3IGYxRHlwVX0r8dylqkOxrwmOp6Cl
xZNeB3B70RLilVbZ1kkEWDWAsz+OZlHFG8r2VIhjkMnJHW+mThI/baS8fHoBgIU3
YlbZhd/Spll/7py3p+JsMxgo5f2qCmfR7xSHv5vXGhoyPeEUDsXiyd4D8hypfbo0
lUzlNv5cpmr5ZoytAiVgU7cl7L93jlff8Sw+pFGnGOvRZ+TUyG1QU2Ow0Y86J++y
d1jyTyN7GvJg3/0K8mrIErv/vTEGIvMQTyk+j6y9ezpumxMC29pv6BV4t9HJxhWc
KKrgNhfc7YdJSbAbJumzQEUxOzpwBEFy0lzb4RsT2tPFevSk6bJv34wxDeVISZ8+
6Zdi2jUKxkmL0jRR/RjmEl20PsF7E5RLOWburVI8vHuO5Kh3Dj0AwT1RLzxFy+y7
7A4nVgfCbs2mz9/MbzJK8B1wEDX9sNcj9zCIJ7A/d4KySMqiyDfoIrPjXOBLiuwb
DSfFTaV0GIZPmph7Hm4sHH4CvArVksqVXIy65sJtLE2JIsBaKcKAUlq4q/A277rB
kTwc5UfwuyKaVYp0uKKYLZLZUoKxleNXWoZS4DTpkhzI9YkHa4TEgtCoaSsUP5zV
8x4hVjuJVsWV/2H9Dy7YKCH0NFqylugo0Z3QXkzzEFPDyRyFFcvydIHLC35Hnv/g
bXPeLYE1T5V7yy3Pr6vqBXISD5pk/+Pja7+xw44IJTNXibfmxo5XINhVcJRgkfn1
UOm4BZYPwd3OGVYSK2VsXXdZ3CfPWLTre3EWCwk8eeZ18/Lhn8o3NG5DEfOPad8+
yKzu4DraLmA7YV3Ev/8NPv3vitzAaMEB6JUSbD/1W0DBv7c4aNI5esBj0fQkVn4B
6KjrdfHJXTziUZ0/agloeMONoNoV9tm8HVF8UivlQxkeZ6bxOqvaL8QH+BhEakqD
TVFpa1RWBn2xn674ekat11w1uTm8jxJMl4aD0xJVH2cZIQCYY6QzsACgtM3LDvc4
PzjtyZinmZkNPddSM7G6vMyw8h8UY/HCaCNqSYRPhV8UzFBp/7d5GKVWKWL8Oobq
32BIgdYa49E+EQKOlLCF2BKQH7lB6OzQjcHU8j9jrlaROCYdlbd/tm/9i4InMggi
XyFxGOs1m7IhOH6ygdkZCqIPcoG2MRA3BqCHOE3vb70U8LJxDbvtYS6rxhibibGu
5Vy4UadCa5Au/oipHf6z0dWHMVeBLyiz2FKQC8j3QmQEVK7gR2U28Ez1z2cz+i27
GJclTD4U7OxBnSrXvHIOn3bEnXMoX4onmB53UkMQ1ymeEbZOjlXTt5ovYiyh2G7r
vd/xmPX3bY9XS6Qsvp8jiMqaE4KuwxK4lLDOzw+IakU/aBtIrg8HTuWZ8BePZJmu
jJekKiTgQlbme2F0EonCSrRwEXNRtJ+kyA9S0rH/zZrj+WhZplcHI1BKb2NBhUuW
eppjzMaEwsIj921O//c3Y878rrxGIytodbJyKZyqktNP+9z2zqRXK9kASg5G6dbd
OxL014Q8ajKoW0z0jHtUU/Q6oFiUpEmgw3IAQB7OclVx7uAgRni8A3cNETM5PEk4
DKHbsvKb4bU1O3W0zkYTKmv9o8vYBEONeJMDo4rX3SidVDPOZqbHum6wuuruvMGR
MDPncCUMxO3bY7CVQRpLTYq0z43SZnJQ38v4PE0ZzhyId3yl7NAE1NC9qJqEqCrL
zPfNFrizJb8CUIhzHyPpi4viEdRWAZPFH9pV6nrjjVOzMZXvBF8KLCGXysgHS0/u
diK+E00NnEsmS/4JqVC7JyAoSM4rOT95/Y/xvCo4rgpoF1WyPUBMAY1iSqgkeWka
WB1j1+TJpEIMVMnEX3eqyleZnhtKcu88aEqnEvRbkTDA7WWZakyqG8d/x/InZ7nY
dBxYSRDHCl5D4rlMmVhyA1PvNkaB+6x6iz+gFLI3M3u8xASrIfrnV1smHT3gL9F9
ZYQMS1x/mBd5uqM21fQu2t5+xNOK/kLrXnBnwRBksqBVqEgeMMrYwhQkoLtEJ6X4
UGE7N1v0yZ5fjpRnM+qYcIwHAtDZrxMKDZ3VP4mLg4LtULVdWaQF3eCxF8ATejup
1tTGBXgaHXC0JgyMV7VvjCP2tHJTULsEPuswQiylMI9tEzSalH5tey0oevIRUe5k
apBOZqqJklkDkWNHxfQFkD0S490O8OPE1DmR1VZ/yH+l5lKzfcCiWZ1q7UPw/E9t
UVvAstJBmx9IlENHR7SCYxeFjYDZX/PgyyXEm6megnghHdsuakHNrAv+ZOiw3Q9K
Fq1Ir7hRZaEYtopGga7cqUie45u7ytfeDdv/C4jVfddjNSCUz4Q05ING6VoaJ0Mw
UiUtGYI6AGmAn3ELAzWvo3jMUvJkq445ODb0HCKLOGJRPDn8sM17ChVy6nOF2M14
QpgP1JHdvVQs43f6C4DfJWBMMzcfCbfdC0J29Peead6+hPVgtGl97brrXmPc1n06
3MzTbF+aJ1yTFlCwSKSj6m2LilVlK2UGFNT+jdILGm0ICjmxYodJhSVLpeT1icJ0
5gI0iYUBO6cIT4O0j3PDASwlTIFkB7bO2MS4nt7hq42AG2XgP05lOGlxrXYbYQXd
rg8VQHH3DiHTrcsmeVD11pXls5MzzvrfNylhQaV0AyQ2QXaByqw81xe32+OCF+nd
VAfSU9TBm7xGD7NVolXOmklEZi4Gkweg/AGs6F5fLFEoRm6eNCvppnPJ9Sd8/tFX
iLpwlZOkx01kBGfs606lGoTMki49LB6SBH4IOQV/JgGd+vTcBUTA6QulQfefyfP/
eqHFSsocp/namxptFJIqx6Aj6KuUmo0VUQHt74WtM7Ca8rL7BjhHZWZNH21q8dRe
E6+7dOqtb5KchpUw/sJQEcz31aG08Rh/ukNQ77XY0eud1gfrLrenvjM09V2reP53
C0j2WEHLXseaE6CojlJrYAtIYNJzZdoaeY4Bw83hAw48fhdD4oxJtge8U3OnsY5d
ELUnZjolxPAikCNZpKWMQ5HcTJ7O5ZLjm2KbH03IeSZ5VYdhNiDuyT9i4WlwQZck
0Z5yc3q7XvWFVZebSHfXLrGd4NERdaaQrNOn1fWRhw2vlND37tms3SR9F49+2c48
7v8o1uRzytHn98hjNcavGiPQdETT4nadiLXeBla3BrxcdagdxtL9Ldm6K4U0ut7J
ESFHYzpIvVKVPZ/EtNxolPS2XD/pwg1H4jCCtDy5kIc8jMwDza9o/NnkJ7xa8kKa
ALfpEdqreJdVSEK7ctrNZui3xVZGeH70+cBZ2oRlWVAN3yRyJIlIvyEq4fLb4cH4
0t5bqTxkvEaVu0VQttP/UBMxh3/umExUslcogoJsF1RBrhN8Y+nQHBgonyr4V0gN
nCWAqgimwZt8Zebi8iO6DkQv/AmSAaYm5rEFWbmRvIDNPgTSa0c45nVsX6BJZ/US
Il1W+LjVqwxamiRcXz8/JaQ/wQMjaDLXcXKryKvvfNhRmQwIPWfXsbLF6gcH8yGW
GpJC6ApAngckDjMppU0feoQPHyv5/9MDnj1Ia9mkjIEMkfmfqsNdBA75oHb9cmDi
Yo8QYVJONkfRFzSkpEvX4rdpqGy9cobkKhqInFX02BqfeLJ+i0GkIM538hAxSn3A
s44zsm3nB4JmXstF3G3ARiN1Y067JnRyQ+dGvGGJSd8avfgY3c6s94nwU96Zhy8T
fW4AHsledxhpgwVM0rLZuo8rUrUU0cppVeuR27ktem1ryNEA3+RILRYeCOzX6g8i
jH1YlDy1Ok/afdZULpOskLbJH3HBuAJZ8FM7J8CZYuYF2rBHymSjMRr7AgRL425i
NGuSAegLk5SeIui8IFvXhEt0BLs6H/oNoH9w5duGSze6Y3PpHDm6OT6HpLZeOQup
/HFMOHeuTjuKKeK7U0VcP6q358RVvSk2xhew9+X463BlO3grycZbaIJwTpbOZb6P
xRbtp6TgmGwyzqxky1tw3j1gdlqV/FGqNokaMjtTIKc2T6wOd4SSy24GQv2AtwNw
SSR46rTw88j7/K6vbMbhhm2Ok53VLSsKB2qUToMOQpKqnSZpqDWZxeZpojoqURzr
hhmj6oSNy28jBj54JxnzYgtadVVgXd0T9zrb8t1hm6kJRodJQB6+E8pBH3JCEllk
+dX1aQmAD3h+FWHEK+ne9F0B3PVQdWmHFP0P2QLCW8n2FusUYungYCoZMRtqYZwB
bmyEepwUTIE905H5QSvqWQ8NPeNvNFnUE7d5jPDeUksGZ+xWdylFbnu0JlNG3cQD
qZPRXWLiOevMrAZs/Q8vZcKeykHZKXpFFMhghdIh5z0XZVq71Ov/vMaj2O7Rm1nJ
dLKIkqPNhK6mZjZK66ZrZMzLbQxljMRA5fsL8cJz4ssyLGrzRMwr36/7IZQ0iSef
+G4r16gQmpQ6OPBKOLm6/dZWQodp6gxnqDQRatxTrxPjoE4MzWxXgCMFbA2hQQRW
yQJ6MPgtxhcXV02Wn3yeXZAMkC2kk4ReloiQ2yn/z9il6W5c6aZ2WmMnJtuYJ+lE
B4ns2Zl1U/Ktv4LLdAmcBddAapHAI/QjOwHJRbE794XtgKY22mkXLwPx/dU+5Ikb
Nr+Gi/nRTYwjt6UBvJdhPAmNthvZcRwsdad3SRYSJAQn38r/nnfSJEZstpZdxq3B
72UKRVYYPZga1AZIaNeKOc01fHPweMeI85TUJODoPvDiPLzSnReINNnZE3sG8q1S
1Bblgw1DoRDCb9N38V95na1TmH38RknVpXTKU9hDpK/V0TXQwgr0/tliw8AsJIgu
UygAstO/HqSNgj2D6kWB/qoGHnYbHBf657Rs8MHf/b33I/giwHqknvTtBM7gfotl
36o8CsCUvwcggBnClITfjfJ/c3VH07m5fMw7mu5wTXW4Br+CH4Q+B5yWmL1GC5He
btbilNuyfJaDS6EeKoCDBxYCbVn0z9QIEUDKflXYJyDCqGmbwCAh3y3fbI/Egm+3
0/a8+sGxezUFiSBzVffD27PrQM91dPFw8yUQFscVSTBS9EoJlT6XQelXu88kbJ8h
m9aQVEN1Pp5ukS8I5brIlizxzsHUe5x7uGc74U2qeg6lEwmynB3C4UE9FNAFFXmi
qf+zmI1R6cvQb/baDTekkaBYH7QYZKqgH/KtrHHWyGcPwmsKd3M42/l1gU4RWTPw
QrE5Pohq+TtoG1r3djh0lhQLAYLYrh+LW+PC11J6zogW6swoHxr7IEEYb4wG1im0
uRY1lug00wzW0/oEhf7BPW5B/x1GcePNT0ODVFGUmb9NwqDzNUA+OOT43bAtcwo2
Z54Nei3IVNbztr8NBLr7483YpxduvCQ0orfTJYbkGCRxaMRDTszFlY91tg3OeMjf
anp1uh8kIMOb6ib16YC0RSZzKKhEll4YjHjLoe4NxhBxAKbAJlGJjaHsLTvcMYuq
Eeau76+oS7IapnWbeTu9VY1ztx2tXKKW8FuuSzaNKNcQUr0KQjYOhLEs6Ppxub5c
6W5ceLj2CN5kRQNPzJlZvKCEe8Rbnz3rJIzKs5Z67Rxu71Y4yojLUZl6yVG7ES1/
SckFdS2haaLRqb9Dt0QyWJuoUqvGq/XdcvvheCnI9e8BzzTCKgkzxMBEcNHpFzuD
HQNf6Uqv897qSSC+sKHEGj7yLVOfg2u3rRWE/RxihbM56j20igqDBmK0iZMWiWfi
NjH+9jBQTWkCgEynB1WARrwcG6SMqqoOHY/d4xG1vZ5dkSPzctpJdb6kyHFqd5Y2
4s2aUBnTewavwt7aSftXQecpeF80j2Q2KcZPLPVlU6k97Y1+F4HvNlINuTthubcL
iBrIi/JCnThpXMUasV6kBZK0KNtWAIC5jznVCodMJ4byPy9JEG6X0vcCgbPxxB1a
RwD9PTU44t3QnmOBFKOEESYqyNvxfN3AwrGfpQPy1eLNTONuuDj/mHHnzKpC8lcN
58MZAeVMsjvyhEyCawann1NM7T2yqd/xn5HWaniv3AaWvtB9QuwFJ/VnfJMc7N/y
oI5tE/2Gzi8igDyoOt5gAK1FfiYKwZEt9YEGp0cv+4k8PMscc7sKIwfszCScBwJ8
FVfM5MJB4po9MMjT8+/WM2c7BoiobvM99O4DOrkh73ypuWtLWeCV+1KhDfYxr3aW
eSAPC6em5qypez7XgfxaTCYb1/2ZcZTYGfqZvmYGqwAM7KiYhKnVQl43/VzixQ7f
EgQD5WdRzwv7pbwHs8ztWPefJybaTUnhqwD/HwEiR4sGwdi/ZxK+dCxGhRLVeOYa
Hr8oBt5+i7rTA+Ee+KzKPaB7be0QY/0V95C6+rv61ve1M7elnxIU5/RxKBykhiu6
mbI5bKosR5wsn+FwS9C3Se4en+dIO0gFgZfiV0LKJs2/5nHpdeEtFev8nrdUeVoK
BUDAp0WyH0u+914BBPCrAAXlfEi9Mdf8FfBIX5JSlurS770oq7Svo3QhImAQ0B6Z
cdYyaCgxPzb8bpXjtdjHiQqkfyJKHJpik6f9Di0zWFN/ZmwEHD2oejQwu14fSFJH
5aqnFPDyyFjw9LAEKyZw8JRIFvOdcQUuRRZMfVI1j2EXQn24QuZtlzEO1VBTmr1S
KPbppz0OqnOUznTsOUH5nldDEqUoQpWLbcS2aMG9q/lmEMnSW9hpI+yqpf0sUItX
ul4UxS6T45rVGJXf8TCC/WzuiN1C14uSzxcoWVbxsyBTv75CaQwB4TO2GP8tU2Ga
CO1NFxbJzmN47oSG+pazM3yex3gOPr93PrKzXBsb7pbhFy8pnOA0PLaDnzREe30+
DciHcO9MOOV+BCPZjjhQR/zVRkDWR29Km22dsJ84l82nXxrKHqja6947xG+9A08R
faDBaYtcHHeWluGUbHhmWTGAMGk43uM60KSCuZ7o2CfzvLdvWgWJSzTaUORxhy11
9xIQtM4mLtfmWmpCylmv2ufMjrvHjR+ivK5I9+ypmnCWoiwahNmYsPhDqX0ZjisR
hD2McaRbkdaTc486iHEcEVyEf++gWT5PacaibOZheLc7gS/bTDWLYzyK1OzvyFD/
eWQYtULhDOoKcXd5eW2zmUZ2JTsUwVWbqq8WkMORBeAhtbCLij45GGGiGRzabcqA
eXUIUoop7HIDDasVSA4lF3xc1MstoC7k36wv76HE0Rfi5R6Al2nsSyBLqA9chCgS
RGxhq1MQKWjyKmYsYRwcoXhlh7w4GmSZH7H7cGVDBgyzzMIBkLXdYX1lXXhNqFWl
wjNbwSzw6JRvW8JZSZf0IIVqbLACIVlNnNPdbfwMXadKL81Gbgy+lQBE+05hv9Nj
R4yFhe0nM7wSAvPCCrJkk3RFMdjXYDtptKZNczSZy/LTVUQSf7OLOpVcsIZ3bfPv
ePo9oGZ3VSaR9dFspOwGmm0jFkzFOMCSgDU5JKboGRU+XPIIEceOombnICwtEk0l
22wz12g9vGGRtznNSky16hMWmU3+RUA/k8rTuRYHQYrRIQx0REWW6k0DbzisBOZ8
EjsP0RqgPfIxEOwsd63mC9Wi8YePBVK2DBZPHQS9wzZ2+KBW5qqLov0aJXGW0y0t
uf4YnNukg2Dy/jGgXfPW5Vcdypk4E/9v4NgzxBhibiZ44XP37FmHdUwN7wMhB9HI
CMNP9XaMXtBM7utNOt1/hoHtb6+VccJT+dmw2tnG00bjTgJTtBUMnTOB+50/snrB
N0SOey4tKIld6bdHCoesU3KfWWOW262/4Aqnwo67dDAL1/czsaVOvs5WfTih00e6
vxKBDE/jyJnc7k0GDcrJTiMdnjzPKzLz0uEusIgUkjrbywqqoV8kRun8oMcmg/tA
Do6zH3GqQv6TxWWhwY9LsyDkdGGvNKaiKS5AvzTFDwbcJf4b/D4jV2aW1cMEPWBo
F4h7/ontZ8ZUEkTjBOoQYw8ksRBwHVQLlAKxTFgo6s9vxpG/ZzR8MZLwdmCnyZ1U
/4CqxM/Go34nnhu4UXpV7nKgvsTY3mT66Tv2hlF+dz9tvpR9dUD3Lb7P+nTQ2dpX
xHSkXaisDo+BPHkM2aB8nY1FVG2RD3/yK8EfN5ovBeY/5zIvJnND/MJy0msLGNr1
7zKYNsZn4slexDx7d+LOIwDzBPiDreI1pYfi85C2CPl+MeHp/stpoDHWrGO3s0Kz
G98rUlxNDM7ht/xNtcpILg5BpmgtxSjdGuticNaNlX306BUvgSORJvnGoqYQA4P1
AVTz5B+P0/iGu03NyshAyjuPUzQF3K2Rtuwy4001sscbeOXpKL6FKMdHc09J+8Vu
h28nXiqHNNaqAoAWimADK81m+Q8DX6GoqKjkM8heOKxv8JakzqVys1cQfd7saNmb
xKk3H+HLvCv0qiafgZtpIfzbNiyQHAnJnGNBg7xtxmtH3/N1h+SxEgp/bGCUveVV
kk/SK5bv+aMvIuZR9vd0LaOrjfymPbIUJzek41Mtc1NYQNB6scAcQi4gQI9MZjDF
Euhj3newrtvuX/weBl9/5//WzWfjmmIdUt45HLBcyKQYFpf4PZt1a7QQ0S66ukZJ
WeCLc7XLgPqLWJ68UuUAZHykB1GgCglEsUG5rVORUwITxaxRpXHS72kx/I6eDzWV
8z3o4v91PANtTPlysCNmZojfCFqtyJf9Tha3K+CuqHpL2E59pnFOYVV3UQ7/ZGOM
K3gWdXH+kq1vAcWsuJ7xVOc/HIPz1lH9KGyV3cvdYZGntiY60OlWlQ1mxJuLBxFF
P9mQLfEjRNopuTEKI8gVtXW6dEgdWn/4QX6deOlbykhabN43HVb9HzpcpBY/1WGJ
qC32qfYamkURH089LraC+5t4UqwzrHgcnLmJ13h47NGloESBZqNKIC6DdzUVdt/e
xjmZZHjCRuxLXdjB1TLFHt/EXq1v11n0JFC/Pnhnwkz3qksHaCvSmPOKfd9za6xz
ygG9kxGKLyakLimkC+VjvAUVjRpJexTgvRvSwrcEb4renL83Uk1B/pMTtFMdq94x
CF7Qo+6xi8mF152WPEh3j+TAzbHVAsh9x2l16Ij1xjuPivyC+BW7PwySxs+nhkJj
t7a+q/LED7h/yh0WYQMJxvsYKtyjhTQlXpkKeF79cy32csTcs6Ldw3S6xf5QmTeW
V34Jj0xliE6oLhcw3VaqPCx3M0yJKbeL95AQT/MNUOOls6ASI8Td6h/RcbZyMY4Q
qwvn2UloA+SJXJuoJWm0wEES+3SLtlffXMkRxCcUAkvLP1Lq1p+NGHXGZTTtCSkY
k3Hj0UeD+66DLHSHRKQ337gcmrKRx2EWztrBDtSheEKTsZZcI/uJLJ+yyZGUzC6y
IqDbgYIUS2lY4TgLm1pFpBq1akBm+NGXmSsEnYJhsaLew3tkLBzn9N6URdYjYp6G
U6lq382pXqzI6ryqrRYXDNv5vJ1UISR1wLDGanb7fqid7HdKOYslmlB2/kUOl3Vm
fCNpwzjduvs53sobi7AAPUX0httE7AycEGG5bxGqL00BILS3xrK/QgdE3KGOgoo0
qop8jg9LedtPvrIjcYuJbEsuzmMDi3k1bhtrP+qtPWzSKexvN5zpmfHuH/xDB2gR
vjunykSZPraHDiXrDNXDUGpdZqELOcifWqrq/lQz3kAJR+YsKLAa0h+mzYk/Zudw
QGIbNwplwo8HJFMTenYX9DjQBt8Cz+F2XQf1gwtFyMhs+I4qxXPp1h6LH12hFwDw
CReyk39A6wvWzfl7ksKDGs9v3QBlg/52gGGl+HJMKeRGlRrTw0L8isx5Uo4BUUX+
4d9MAGWIRl6lLJCGHRtZZbizWeCwkORsPAdypRAPWPOHVP/poQ4HGtJ6t5xeV2RX
7JIU/XZTj0s/1TBJu3Iy5u+3pNwyx0fd1vpNH+jk56bh/CxyHAlDaMsOiZ+UXFBS
k1JWHcmloFGV2j7+eCjXbHnodqOg94P8CbW0TxWkIjImdn52c0EINNf+7kWZF/mV
2d8lCYl7Hli6Ilp2iatfar7QzwJ5rfUuJIiGxlZLBDXPvGugQ+VZvF0UKKQAahTf
EXShCVRGlsTICen1DxG0ZxbBDTc71/rgEA+xFP5cUDlXrUdFryK1KMC31PNP0EvZ
cjdx+uZzHx4skmejpoYqofi7d0UKSzMP/1yExHQfITd32HNa21apBhE5vNcgu3Kz
SymGqXiwAkibhWe4KyidNCla8sZh7ohfasQ27RtolKYc/MHQ+sbL4CuwZHJclFaN
uqLDGcqhCRJNMiI/BeY9A9BjGNlajLDW21xc8TX6jB85rB98zz3jwdxBeAp3ZX/e
N7Gw/ex4JRDev3foKvd7UMgMwC854QgfEautdw9ynysebM6uoqCpp1Htvu7IyLxR
fpuE97YiW43yWF5nHMh19AjyHdQvbW8nkoRws1Irq7XhrTi3ZrnY2UtL78+h2bCi
+VM8sK3MtoBeUN3usNPoyWROE38ooQur4X6OXR9zgCminv955mt/mE6NwcOCAL0B
pUafDxSVddJzvXuxkmEzwYVius9fFTFfjAWtwHXbvvveNyA/fasQ2VInnqXemzeQ
IuEu2t4doguKjkHCu2MO+n8omAzAfq92KHVoTZk+G9zyNoqp07Qq4osnaZz8/aIe
E6pF28j1UEqeQrJyN6YgkYTb8i+FMAIa+dpdvf7ewHfRC1xLQqVh+cYYHO2Fk0j7
XloN3Dr1NwFtu+OfuubUU7ugG6al0kcUnZga4uhHcNoB+emlqBmEM9HMJ4XbwfgY
aRXGdHhCRqeJzZW40xFYfZHt1DR3YChcSKVsdgvHgC37ErtlOKwIJVZs3lwfVWiW
TZjHTs84l3tHs0q7EzOxpXJmSif8TBoDhk5GLv5hNri5nNAFe3NcT5o2YLhRFiy7
UHO3uoCDGu9UmMbpe7IgiY7w0bsVo+lRlmbLSKZrtvsIb1k4ZyfoYIrA5M2n4kUk
rZ4W5jPxw9E3tpfu+AKqT6oZsZyy2/at2jcdv8UA9XZWB3nP5GyQphIpD6FV85/i
CYowmgNP6XLOsLB6VwUQ6HUYyNwe0mcWj4bhjNneyFr+obEi5b/OtvYnaxK8wZls
ZA1ksjKb5QiOIFYo2fe5Wmc7sWgC0FFkN+J6JPOVaLaFM7QAR0PvDqk/n3d7zLn0
WpR/zGdCue3p9wQRyOQk2n4Y6Tc+dX+WbpPKPBI19D4N+f27fKf/5bgIbcF7YChQ
pySA7YkpGVtPVHiap1K/Rr58Z1vjZdSRjauWa7GlLDGC+dPIoRjXU+8Pu0lP3JQR
KaTF57ndU1QgH6WXHCPf1xZePb2ePJRFc7wu+vlPwj4bLMBvD8f2XulkaNWbBjRT
lRGZ6lkem5IT0UtccvsbR1iFpQ212JWquzutLwfd2r/BnAudJ8JWE2TOEiBL3d5d
+d0cntr2FuYWP8fhUFpnVEo7BP0+clUw92As8AWvOwtf1q1Rn3W3G7I89cqT03Jt
mWu/9HGUZE2OsGcpOzja6ssiYUy8LsPxNxs0XOZKrXOhx42/DlIXGdZ6bnDhsWt0
jJs0aZfIWF3icSUnUTZTznTzMHuqy28Uw25aSBDaUaSxlRYQytmQp8ZFCYL06wFL
qDpHyVv8g56NSxMZyh1h6eL2IoGFqxW0fAwxjxQd3v+ZXodesmwegFjynPF70d4t
sIKaQSkOkg+Z3VCdBQMjrDmeFTAI0YnGkWUz8lPTuWuyVN+zIm7b1lscBO96TMSo
YRtLprD/wHI7CFUbP+QtFG4Vj4iSL8AUb5J7krWefPojaIAJIyRavzf8rWYZLmSw
pXYN/m1IesyY00vf/x01NkahYoOBXT80bczGO0L5i6Tjh6Qt3sPVCMTj0DDo2Jjh
wfxTi6zmeqc6LseYfSdCFXDP8px/dV+KA8CD6HOExJg/vOIJEyYF2HI/GVAoipir
nUwtG8Gh36Sp0zlv1sGgFLF7sPcFtytmgKXbd8wKDkpVJnxXGfF34+7L+jnCxVQy
9wUL/ZFMsRCdrfohqoOlefTx7GMC36IMpUJVLJYs4g0SCIIVKTfUm5XGaVGMqxsD
uBh5bDdNuFabS4zA96sRdUtTh+qNyHsuae2I6FiNX340L9s6QAsmcP8GBGePDrq9
lnG7yNkHBbWnHdfH35KLglBW+JUqdDo+0L/AVz4HLs5vlnUEXTqZhZNpROI5KskK
A8aBVav3aUG9+COM+JnYZEwsXC/0bZng4D+cgt4VtqQqnpjEJb2Dilu1Vcvjdr7A
ZDb5n58mFWHWtdKPLN6WbTq2MLwF6P24Wtb1Zk/MkAEsK9jufkDSIzGXBfLXPfkZ
TIxez5qDk9+SgE1VRYVgW774pc4aG5BK2QlHioX+i21rBvFP+iVZhXz+vA0l7aup
9X/XN6l0dRrm4ER6D+9Sa3pMrQIAR2ylr8vFy7r+wxo/mv6pFbG7ys6UP06X2Zuf
ape0TNZI6lvk6HvXWQg2mLnmekPyzmOKVWttlvllZyQZnYE6i9XLeAmPhhXQFzba
jgajiU+Wy+U17k1a3/BANBvgVfTLhDzvbFyGbM5q4lfo90SuVobSA7g6Xdhxmc5N
07I5X2te5xuNZcC2PX/isfINS0A6KOkxBlIJdVtZTF26SOI3F5sXDCVR19TF3oWR
xwH1rAy44Df270fEOiIGQ1v9EfdGhIuo5rj2wwQWyMOmvFnhDxfeE7hdSfkXYm+t
KBA3XjFrhOXZiRW1GhaQQ2u4hLfDRNeNgFsTn0wU9PM/6Qr1N4Iim9K+K6S7bRSf
J436E6qDRgwzxAPUKniwp+Ew9ObzddBRacmRFfJr/Xq8ugGN9211ysRTVh83SxJC
9jqEdKf2HUCh0QzhxHFAhnwPmNzG7V/JqJGcxMkwiepcbycG/mUDK9pVpFuCNYUa
jvDCOtRxBTdfUwu7h1zwIS8pw4Eje4mZsizOKyegYpgVD8/lv68JkGXO6N9tSzpk
gjpoyxxBIehgu6AsLtmBUVR81+HOJlfj2qkxZ4piboBvmh1kaFSmN7wkoIvMLrMB
QGplNHbqYdPCE6FHlIyj7xXZnQEqcttNlcFTU+hPivUGjeXNExLl4+AHAXOARmYC
z4A0boeMiVU6mHQ38G8JyCf9A7fdflwjZjne8FEzy/Tw2oQuuFrCn5kdXJ8cp2rF
2GZ9SuKwYaLkw1HUakBPWnYRAv8T08jTAd1OQkB3UctULC7BEWwUapSBwHlynA/6
l4u84P32T9Xkr2A9JU9DXxMiSH2sW7FBOdNRzg2p9/iPLCiOCIAj/KnBKhthxtMj
VAnjlfhjyt4OA7C9YreaWRlWF7msmqFupxNwNeEgU8GhCDq+A82NB954F3PVc6GV
vpKMg6qh6YwzMOPPRrOJhQ6+SAfLf8xSkXBSxcMholPtjocFe2FbukVSYI/i62Qn
XBmtfKThhQoSzwmw9pfFyCMvsBfPcrUUlywCKA7uNAQv/JorxHgeeYsPY4LtTs2R
WnJ8JhNdJU8Ae5Io4P2O4yb/7IMd2AonA/HOIH5J5Fx6BDA2DaiH4dLIKA2uapu5
gqZPALuMSs29ARVj6BZKumpJuSOj9DSWpMQA9nL41aE5Ev0TeEEApw0yTLTQ+RRO
sIirX1XOQm6BaQcaVMzclvAsiYkGogLX5cM10jqmYhJ3PgJsNd3/u0RvAUSvk6KY
5Ek5drofrbYJlR+BRFcKqIq91DqvxbmTO3vBT0vmw0F5H4K8epg/qJUVep5QwdJd
kcrGMrlh8FtiJJdgKYQ0orf+rGqeSlq5oQV2nzmAeWH+jVmyvzJIpRo2c8Pbbdl0
8jRS4aX8dEYZdAs3LZQLjf4FXhAzdDp7mE4Wg1UyLOY2MbpfdZs/lmTCJFU8QOzX
m+loc9Pf4vu51UPilPhH2mNrWDsWxpv5qvo4/tovE10UULGgdiPjUZUTkM/YFZkM
1vixJL0BgjhAn46ujYlhdQePuQjn98WSJnMy1nJXqI8TieAFH77SFkoM7eFCp5+u
shtVWGIaZnZ4flmO5jn2HzvYI+G5WJE7ASWgtNfguZGshxsRzMJAqUnKcjhRtTxW
JPK9mbKUPKETrjIkrv8bf16sgYI/WdgW8QdxUQlYsfC3xdBwa62j299Fpb98q4C7
fMHjK95wX0rs4MLOdkyRm36gvKuvsWo/mpOPqifwhKz2MlzLGVaiLVc/Gb5XEU8X
V1Rg8SctykAQNaD9UWOR/PpMHn+GHXczQLIDtDKRLLHGNqAR5MTQegrbpjONd1KI
2iqgBtamL84gK2aeVQ/x+yD++PLAHfbpc2OB8BeODWW12XRM3N3CN0pLvdVPl19X
c4ju8xDHCNpfxiXCgl1ZEQncPAyHtwnCHxD/uYtJLZdOV7P890JaN+giYNB84vl9
c5w0TrrM7DH5XE/ZZE/LpKvUGwnzwjWXgowy06yhwQVOXrYfwurl+m+tB5Tb/KU8
pviRDbFIK5C9TCVUMxybwSOPclO2kX++Cw05QtxLx6yBmQCO252p24a+7j9dVWRB
Wh2O+NSP2Q4GC9/qDNIIiL8XMykx6X7Of/rrDml2H65FAoXIPlm5c+hkMBnBZxqB
dzeY1q0gY+D3oYJPuI/Kd4byuOnuc++tcEe6P+iFPb+FKOOMviexLSZLXU+AV+gr
QBdegET1D1OxvX5QlsNJBDff782zf2TD+XIL0DLP7BGYyGE/KVYvPLtD/lvt7u4/
I3zupwkukHdSdVTO+ow+bJYqAjP+S71wrPBlnMrLUrMexMS64iiPdPajeUU6KzKR
UC9hlX1/QiSkBp/cBoqjmX4Pv79/Gz81rNT3YFFnmvchoSaNILkQsX45/T3Gwn+v
itCs+DLYRaCe2w1ByFvMY90rTU+T0qGXSzDUHtR2Ru9B+xOOxIog4+NvQNEwtPyi
1CEs8oV/tLqNkCW3CHf4G34Uw4cvoe/TpBfXtIhpp/lcqKZ0FaBhc6EAKFSvtMdL
j9yvpdokKHjJlPlAW6Rlfd0i9bU78X8WCzVs4aCAmd+iRPTe+n0Q/BTXD843GdxG
mDlxcrTo4BnTMvHK4eLIDPutykOv98pWNI+66Fmt63sHqI1mbvJOurCxtLUCzqSo
7m2TCUpsqeM2Lsc20VBwCOEEhDTmKNL9HR0wCTUBToRe/D2RifYDZNczNcFwtbHT
OERCcjKFWbA1jTszQZ8UL4XYvSZOJ7RjZGon/hncM5TGien/SGkeIh3V+6zpOQeY
i5YeiMyW/2bojaf9oeKMFs2sG5fTvSepSF+TwvkBhSMKj+askcAMhG48Xm83migp
o2qVxYVm8i5zaV1HSOyedM5Zxt/NZG0UvY+Kyl+E/liX2b/kapmtT1P6O5cZXxlc
FQcK7fOq6vQYR0IX0XnnFKHPJtKZyVFPpaeAyD3fZt4ZxfzLKk+XMvt4JfaovhG+
2SpLzO9rOB1CyktJNKdS6rCYHbQakwlzKCgWBi/XMBbqQ6ScK4KGBIyKJFcagCZJ
2SwTid0qBBNXxyfsMZaUVAxsvBp6fmz5LEqzlTPsNYV4vjRBmPKC4f1IcpO53dHM
morxRP5mHqp/82JeLB9OGPSRedSwMdOXCNR1fNGLrTDYvsU397aCjR9R9PxjD4w3
uOo/SbnB3gRl8p+zY27EpvB7GaeDYCfEtLCzESFX6pCH/ZVcw7fUt+yA3q6QD52X
TwM8NlRjufbms74+L1ZxAgS3KoVQk4vVHTSAfeVZnjgnKNszXIjR9xmAAZk7DMO1
xcllcwFucjPvda/10WDCVtkH2ltwsOnGh74x7hUYvizMVvVlzwLUxZkOUxDSGKeJ
XQf5UbE/rh+h7vSnV7byaK0CIJoplHD8hZ8AF0iYqArWJ2aL1AWgFrpTBtScWkIp
avp4Lisd4xS21Uitvl4y94s2KX9tuLbuDRYJg3f51MgORWn/o5ryR949B4fm+98s
v2UwZK20hcYQXAH5l5OAYD9Mv64xgrheKG7Etyu5BIJvVwz2JTZR8cSdrpsOXSjS
m/pkDfdFBzZUGIIvmDjmizB3rERRPFRQNNPsHSG7J8RzSy6JON8aG4fF42/rUlTA
ER7Z5nQOe28x3FHpjof8FutjU3sjFSewdx5IwGp7JJpAvDd3DRo4SDixPCEN5Dvg
lb+x2SNQTkBOqI/9T72GdUjfg3s7oU7ZJeq8jpyGqQvsLtGnstGSUuW7RuELnNVZ
eMMn1fDO9eLV8daIo5cGWKeD4nlblCBxBJ+srQPMCMLL5g39ONRrNoYULYyJBLdD
IrKhkAdVfXRbdkS0GMxu5Bjp/2eGmBP8j0XNZ9TBsLZ2VjDeOFlgTNwRUsyAbjUK
ilSNapH8dG6Z6GIKerTam56jQGOJGKa1RKotM4ETuaPf0gDCivQ/YZ81uwujBZJb
tBrVJtbbjyLjq3QIN99GX+Ty7sX0ugzJtcaE925aXV1O0I3gZU6/vXH6drTedgkh
HtxtrUVWeL9ydBRJBfiat5niPN35KkuV6Qt0TpYylWu0yEss75TpIi2nMVebO5/S
RrJkMgWxrVW79KmN2kQRFuNCVUwNlRkW+UKM3fwY+qW10ta4QWTerv43cgAfp4wx
XSvJM0us3MJJY8deNJch/IycVYPwD2FcqDWmZLLtgNi71TjJeaesT4X4D526nDLU
5OdJxcFsqGOircf3Fc0BybB1+JfaLRkm+4qF3ktOoYncKTuxzY3lQzvHbktQODv3
KFtxYRdH6e6pOgXbaGT8OmNbDcp7BUmFdrqjFZk61zM1GPaEqAkReJlbPrCFk+Om
upv/M+KNd3NN97G+mFY4lA==

`pragma protect end_protected
