// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
a2PLNTsQyS4PoQATxyUTsYByQYSQlP+zIaTiVi3wnKPrceWoZhMQYddqdWiw593P
ZV6bKp1mK86EKO/dnsBLFaJieZeZuBWSjf2sFys+uNAskh3OmZomWKhWVVkYcwzX
qGDkA5A4Wg/CYLDQQKcADDipXOSm2s0X6gsA+j/d1YecmNE3qDl+/g==
//pragma protect end_key_block
//pragma protect digest_block
Gc5O6n3OuSprRXtOapG+TMsPhks=
//pragma protect end_digest_block
//pragma protect data_block
wudUwTd/SJX67Tpax+B5eSFFsvbItB89QKHuNtuYFs1eTu07UJRyKqvPa5nh150G
Xz+CkjsH7W+3ko2LLoa66qyTe55C+JV3H7TQjildrvan+uYf9fUQu9UR8/DG2pJK
Q0A0BKOzFweRmct71Q3QbIjIzkcKm97ANAK8Vmmtiwqhwq3Kn4kXnt71MNNLWS4Y
5lqxfSjwu3vQEY5bldKQPuebh4POPEhhazgnirax4qZ/y1UWE8UWgu8kYPWNurfY
g7I4Pt9N+rKdT3rJpN7Zje7rt/nnTkLbijF83Pyn7GAb9lns34rLXh/57qs7xIV4
an8P1OMiGVS1EbVwZvmkHO3IOOcSFjepxfHz4+OVphMF/GDF+WpmKtJVtxIQrYKZ
FAPa1w0kVe06XNwHQSbRmvKH8AV/AFXok9cWXcnCW4BwZKio9QbuHcy2c65xF7v3
g4cMGHg9UfeaN1lZViDLlDXNqJ+0oJV94ub4QZ2qV/YZgP5KnsKw6MZFHpGMGPt/
anIx8DRpyCJuNpob6zq6FFVnH3LZ2+yDcyKe5KWTiB7S3M9eQq1lMkzchvFGzBPQ
z9zFTD06iJexY5umPCdddvviWx5z4QUjq5Zq168YF4CcgfEdhMffMuZ8d6Z718Wp
ZOZX4zrnVwKEggSt9QFyVBbyYnrnST8tmpwYmI94/hQYfMgXQTZzS0EdK5e1DsEh
meNdWKVrLbaHTH+/AL785as2F2hurgJw2sZkexJGqxNFWoPwT3wphtMolMg80eU7
ugVzTVFyFAB4W8/yoLx66l6U82wclS0d2GJOi2qVKcu5SlH2dC9mAaN0g7kCBh71
w1VjTCO+uRisCplssmlBYeDcBEqdnMrSxzZLP/8tinf7V5OIFl8cHXViEVEkqg2A
uQdbvO/+n196WksWBD5iLzd10HZL/fLun0OtTg23hIFwkf8SadrBnBryHRpVlQWW
v6vSTqwjz/XaOqYhOITFLHVRwYsHs4ghDkPUE8f1eSqTiHAn4pB/eYL85cD/hlhW
30YO4mezVywx+T5LT1UncMSGT+/PQjYtRqALcDySNg8tzVCG29f0HbhBuQUmR9qx
JDWqQWZhOumf3f020KFerKUCAbapw5gBKmh/DK1yGpXC9BoArbtH5ho4pJaFSVok
AKs6oVnogGGzhZ/EbBs1Ju3K+bT3co8l3EdtduIzyxN9jjI+Lwbxs8MEoLFBPF8z
9ctWPIwtobrLRaUwX1bMfgPVoaw7vEkvry97sQNOvj0CC9d47HiKLl7FUM3wWniB
PBEvykVsa+MgJJj0wRNCxtH6TSsgRm+YvCmFhZ/+ioxVVlPvFia6eYmMxwC5fFw2
Ua5XzYPBt/FfLoxiyKJWk/7CoYTsVy6hHhy7fl6uaY2DDkirLNIEAFF4XU8xzDqW
az5di/QFVCRmUrphBxqZjPRav7uGLZjubcYgZDopDJnbS8DMSZhLJY/XNqVvvRYv
lYuc5/SrFZp7B8CnI8ctJ7bT6u1gDXZXXqBjrQMujH+qn7QLU4opbPQTMZUxbIWG
8j/+F9BsOcsDNtLpqFdQWurT6ZVR/Mrn+YtaCFICLf7sr++bL6I1QrRxu5iw4JsJ
ERGkH3nT3rJ8b5Jj8J/++0C8wfC1FZ9Ec+vYPAMtJcVcOYntW99rhy+rfXA1IfEV
jPF7qmIDJEDa1pauzGppLzEs9Aga97LiLkDsA5XHW9DSs7V4YzTHbuMbvJVecyex
zcsjT/urNTYarYP5+M64fTAEVBjBOnKp6i9YAIDP0fgZcGYMed6rKmW02ETAgpxe
kAckSD+8bHXIN4HzbbZpTS661/Ynqyue0/b43f4H2r8rsqJ6o7fZwnKCY35yCBAE
CEBtxz4g9WOD02OpIvHAVivIZSgv042Y35NP8mKSgUeKT0ADcyo6Ns3K/1YUm7np
GQ23ZHkthKRU+832nm5M2BAUvs2KsU7OuIpLPvYXS2abpznhNuPK4oyOjn9n44oZ
AVj0++XVQIfR1epWLwrd/WICOt3Me+8juLKNSe0sG62Kn7mgR1gNCaBWRfSGF0XM
FFwm+FmV4ZxXlHGK+7qAs/l+/uy+Yb5hdS4WSDeOWpZBOs/BzGcLF9R2+gE+qLBu
Pw07tdW88r2enBzQ0JnlXmCt1RMoxlNrjx1S/1aiQEkUQZFDwEywyzHzWOq9BU3P
goROcMW6CTVaiTzVBY6svVTng+Varz4ttn28q7XfL9XS+ZpK+Gl3OSzi9xDeqWAa
6BcQYdWg9EtDxEEamqw4O6vryJ6jL+DW6Q7ivZeQqbPh8fceYcAisM7tUzJOwjrh
cOBI253WKRqP4YWKOWt+eUTkZCCLhp+7bcOiPahobdJge6Y0yBZE+lah2ejnoW2v
j0ZrOifv2IN0XBVjMnZXeXJYJKDIRNRrTHNwi4bkVpE8tG1utP+rvDfUqIG4iBKF
OxzWmFRxSSiw5E0BdO0CJCchbflsdTqz56mPoZEiQPdH7YCRPnw+FaT19efwzre6
ZtkwY+Oft0PawOipztsmoJoa39t1xpCiBM1iy9fyQBYAWk01YE5qWMTZq4WQlEiR
0r34PCPLvH7djLQ6FMKP9laC+O8HUyA69ysPoWWYr4+uDcie2a33+E0/Ugcv32Zh
MbxrDwI+jT0g3p1u+Op5QYKjyn4Oo9G5uoPBjfzOetD/hSBUBRpJ9DB35UVjI3hb
k4DMXjuPq3DA1IZrEHf6HIjYq6SdChYZzGtDoDlCfLi5V0T/8WWkR8ccFz/hxLR7
MfCldxKM6x7m/OrbuXUeJr0KZ14RCNMk3LzoX0UHj870DKs/BtS70quk9pGSBuXt
tnUaF48OQZu76YSexOLAZSSwVEymVcdsXC86C4LT1GEcwZUsCAK8xxnM0XtjAnv7
x1FZZeAxdRUbFeE/9vXKU3zuK2aDIGfYnkr3i9Bu2DdCYFWyHklR/RwHTzIznoLb
DqX+pxFwhXAs37unZ3+37rBVeuHZx40SbX0Jj8ujU00rYzCdvrw0lmXiRMlf2M2d
xQjiBuEXZ9p6cvrwhpwSykJf6O9DGVmVmKTT0143wiEaAM80i3xOdYBCsTjh9nV4
6JEiPAJtQ6XaFWM3DYK+wdM9laYL/kG6APXEEMy9dEoQGdZMKoI5lgGysw3K0aPR
Fb/3N2312XfUOz1MiyzUbmc01Tc2IqNeVenBve+oAEwAazG5LJK04MAZXb/rg6FP
xSk8wYV4CA62u9oWR+cBlnv0C23tbPdr3Wdh+aqX7k+D5Gxx6/dfclma0j2WSW9J
+zrZbFSOXmzAok7cPfWD+aQ8KLqoOSV25Oe7wJ8NxL6ruLjxxR49dzqfOCuVZaJu
QmZYy2HYyjSf02s5nvPwxHcRYVRgcgGMxChkzFRinBaEAPPZZ9cDRhpQExcZbwbk
w9D74fgYukJMdhA5h13mDcgtTnIQuKcvymVgqKoCf/I8nh9XOAHL41npNqwop761
y/A8pN7KduJPaJrZnJXo2uYG/iz5MGJ1HPeX7HJZwVw57dau9CLlVB9dWYnXKCdo
mZVgXX3f+pLF3EHZTQOT7isXYwhr3BBw+ryXc4UsjGKEXGeJMdotw8yi7wb3UZWX
gkJFjfyCVvLgLwSCmAHn8GHUg0sZY3iyZTc/gD/j22QWL2yMG4ttcnT+0h6Lh6tn
XsTqKa8ELxwIVHCCkwiuNrE+WV4KvDeORaf4fbv61x5k/vLT6ohB8w5DbfR+1NX4
UAK/39P9gf5BoWXjb/h3hwR8h5ugquunOhFiwufzXNi1UDBM8t5vg0iUfGmF3QzG
fVqSyAEIyjDBN2XXXBl6vdopmUUyXEd7CP3uu7kq9BRgk3FZ5Q24HvP0SUte66dt
9qmSA7ARzf7cvXTXNtfYuJ5sypAc5S2U7hsNbOfGnMRKiJtleqNzXcX9wHO2Xcj6
oCtAcggkR0UqRkpg82wRwLxh0K6dX+AC6tbrtynr+dkwo0BpsoUI/RTe4RT810SQ
tEQwYp9fCyo2sM0q77wwpaZjjhSBxtRVwUj3WJrpUBRTk8VH100/0Gnu1OYgcKqQ
JLnljjFvHoikbxG3FDsQob1ZEnFZiCx88NR8jMRK2KuLdZTOc66VbHoy9YHxYsZ6
NEiiSaUMignQIKBU/ynIPOboqubfN1r88o1jqo/Yj4Jlvf1erU0CStTgqEWNNVKv
F4K9uiEdgPdTKbEFq1nJgdt6XNueWvJN4/9R8178Kmzk28e0DUq3/tN/wyvCO1t3
W7HiDbLVHBQrB/7DtdLQ4+oqPvWHcb8QtMsxK+d/TEFqG1oCUOFt0b8scPoUfdYT
7UmJd74JQigXiAF3zl3ZkHlhtke07Qb69+HVsi4UM9nl2qFXJYZs/m7ymdhlhm8b
27TH4Ork6+Efb8vq46i3fSmX1Mxta9vlViQ/MALKBkkRyqHb0slZRacZFGXFaucC
HnpgbRdp5pAwqw/oQRISQCthYfdTImtTjU++mU3z5I6lWGFDK/t0nm4gBqvGcQyo
7tSNe+lYumqQ5tIlX0H6Q512LTrHNoAe6nUk0GUdQN4sAq3MnpXktusirVQkoMTc
bqsyd3hkFjRHG4b/zGIDussir4YnQLymgCco8G+A20xjIM56ZEky5iFHxTaV7HOF
//1FEamDEbjUAmuuSJW7pDiIwWOnJxMzvgS0LCSHsiZtX2icjMSrPs2nIKvaNZr6
Ke5Z/jWFcNCNt9euAnHo9FNCb/e1d/JHyvB9n+4eD1Xur2AzCeo/3xEtXUeAlDcm
hIdrYsYnxA9jYD6go/DSOq8VRkI0Y4u4e4gsKWSeqS9RA9xJBBOm3fHD1/jN4bt0
K6sG1PkEoGWP+QIfHrAxfvR+go0xGMScvypyAx7xY4vo1rLgs6IHnMd4PIjX1Gi/
4HOot6zIxgC68gHcory0fRg4L3uiURuKcp/hYRpGl7VIsBQcPbyxonmlam0N1HqG
PvK+227/+FPG8I08G18TEnLzmZ39h2s/rCHhBOP8PTU39/URPz2B63fIx8ifEk8f
JPU6GiNjcxTAmg10qiTHUTuDo4E37kIp7tj2biA7XBfVFweVMGy0PMWvePsl1Yp4
Eva7qVvfFuY65SDIaLQBOeKq6nwfYwq4UXsfhGcogKGggt/38slTMbcieLnSiaS5
vGc3alOoPSoIlRiwm5pGkGooaWx0i6G+du+m9SFLRV5UlVpMLzoUZoUYOFoGSX9M
/S4104BwIx+IDk2lv6FIBOhe87DmCH5l17uaMkBnXxYnER5/9mWVBwe6ESwq3Ydl
bxokTL0/gfTB2CJGlYmVYPzFWmEQeSd3gIADpw0uQxWJX+dmHzQpYCpYevWqvBN6
xEbOPa+4K5H4rJ4MNzo9AuwV5mWCpEAQqL8axAf/le4MhHAixKnmhkv+p5WCvNeN
VF0LW+FSTm8EA5naeb8rNq5Loi4WT9uyMx8isvd44uiGLlLnfZ22XV+F8ZFyjf3Y
udYCXZkMpQTjpu473KquPXM2J2CLvqf4s5J4QiSnyRTDNVP1bECsdgLYg4KUZbYv
NJieHdlM6KBAg1yM3EMjNeBQ8UtVFVdO+8Ed2Qw0eA7FWNRNXaj+8BG5iWEDMKP8
jh5ng+RYSPI+BWUYqj2EHWNno+2niJbPBRQjtfKvjxWp8k2WPPi91uHnJNfNtfdT
WUDrqLkcTaYPu9/ltTMhdAeweW0Rla2FN6mJaGZ2EIFNpMvC4xSUsTb8k6vFG3QO
DQHqNGCycefshcG7rpS9PiT9LKYmoP0yiD0FDyWUcm4xTCa+ZvYp/oopEoS0k9k0
14XOfGCKJmLeSBpBzgX8d3CHMnx0R6HpUtOUoOsV/g9SCbv7OwHH9Gky0pNHVown
NmSBMyE84Z0XvA9icApjsA506Q+zAdoesKlLuRAr+G7dynb3b0EN7u2JXX/OiPWs
3XNPmGy6kAgYqeRcnCImoF3XHC9a/yLE+MHBOwisOIXIVDfc6hVOXZ2DYO47lhBz
gc56AFyuZk4Zt4EOiiyC1FeMDqi3jZ4WjITf7grlnRv8afRdtkgUuqfj18up1dKa
iojE42G96pHnEbfIkpRZaQd12Z/yagUftioPWWC4qWBwXlsFKJKiz0o0uIPHOf9o
7H3vFB8TI9s+mCCUnQ7LudtWM7vhhIQD3nHvrz20XgjYJ2Maj9nxyHfVkz1dBu6R
ZY+OTumpJCGStT0c4anR+AwJ0yUB5mcYBgX29PQB6zu4R/ZFIlOdyTOPF2V0AEoX
AgZ5W381GeQIuscKeoOhYVEMAU5sgLLY0cKVfSFM8WpSvgxvYlmf3oNEZp+6LRhL
e+UoNawhJBuV3xaZaxKFaZ+6z55EyNtSos3U7ocT18ovQMwJQuGL8mDh3TWb3VjT
9LWXLILGS4FbteV9xz3mc3PcYvXnCh73Ey7hx57WCALCH84omRjVf3Kvh71p5RMn
0GenpJgKB62rEdXk24+U9vvdm5RPnqQ6+Cwi5gHQ8zxr+lkmAG4UG32eu7JCK1v+
i0pi1q9d5ZXJR5Z2fyjxDcfXkj/8fx9qXDCgZ/SFyiC+7AcqVVrpULnKHlWudPTW
lle5+TH1ZCWnpGSGb+AyP41kB0dPIxazktKjpibjd+QXu5KyZpgNLgxyOfMWFol0
6jJQqxfpPwCP9T4D9SaT3fma/K7G8qu2uFuQpqovX9Z44AChJgACAIvKz7Oa8Sej
XtfMZ8bqEHuTk0WLd2a4kIK+8qPDk00ciDvIrTsbrtUyyPWxYbFeqHJ7rRU0ivpD
Jt6g1JifLhdn/XAonBP6uT+aR0sY03jlWjFC1l4GHtlp5RuEMwImnrVorZKby7Nz
txc7Y7LnT2Bf/Qt9kaTGX9Tj2lHfPiq0NS/AZK6/HK+AS7HE1llt9bvTEI6FlJKT
NYsP+SxEXWKGSgudP+My1cNoI2bQjWri9wfv3mXAtwoBmjOCqBjHU62+EAuJGK8T
TcOnDNEz6v628Bp5Mzwl/hJ9fh+JhpK0T+/MpDRW/nJPnWp0YM6gVq8qfIrOq3bW
4qGfB90IUhwwy2U6tg43DWWl84nzoBycqEn4jj3SPSBvjAekOXbkeT6k0RzzydSM
N1IyfTYJnH4fEuah5QGm5OV4hdpPcXurBI4UfR3GiYnUDSA/pJ2V1L3LyjjtPyF9
+iYVfZEhA6EM+QZ5onrdSg1NzIdCChgE4jAIkS8fNtc9hnNmkxcOhqe9WqFhvKZS
V/2KNd3Ao2sGasWKQpCb/9LzBJfG9gTwXVKo0jRc7FYBeGJ8G5ils+4dIhj2qjr2
ST+RmoK1IvYQtWMLncguaHYgsG+i/4IVK3kQ6WDYpOH9eYbtlgq1eeiXGqAxDF/A
SYGxz+gefnX4BHnDS6o4r/NXo5fE8SCadA1sw0fngmv4f44pXJA2TPPS/nj1Mqi/
Xiuh8VQ2TZ0cTH0xPe3PdU4Am5PsO9LiM7YHZXlZtmiyoXCVoRnK4a1YdFfSjAA6
dazHK2pYRBa6zjxHYQJJOXNL4MQ3/w1aGhxHx9QtyYmt1ck/AeMLi1Ux2l0DWXOT
ZTVkIbVcyXPyFHQrOtfJpT2Vkps9lqM0/zqmR+dlYIRevF3LJksNhVyTPmGTMVnb
ru4Nc5HFXCKClpjhks/TFzVtcF9KD1CmqvkXHjVuJh5G5X1q4XNK3TxVGuhZZsNd
gpS98ddVejZRmTMV4DJAEU0b6uMzAwznbLccat7dQCmAuxMLWnVPBhHi2Ng7vKvS
HIoNTvRL3s65yVIEc2woCzKNor8nb6Zo1qr0dDHv6rJAPsPeOSY0vIY6cvo5rLIH
SLjq406zUk1P8TLyAto3GPaHS9wLZkPoiRFiwPM7OK6hzAGut6WRJuhDi6aC078A
ulpkQjJKkb2hIwLZ2G7bSRwR6j9Gw8nJLxhkiaKSzDPZ99QFEzdbBVN1eEdQvorh
Jv2+ciOMi3kGDNeNUigWyfsVO6GtEk4MOC9JeHnSZJMQOfyVjLT/JWolnOWSoZMn
Db6QJHOVMarerq20UAjGdA0yxnFhZ9c90figWCZGsz4OLBwDWIcIqYnCGtMHHz44
6aVex1nj+npAms8L9o7x2ZshE6SmwBIB3jjWbhRS++F4Vh9izc1mcMGUGnJrKYts
8EKOj3T1K4KAcA1hgTadeemJQFbbfL2Msi+xwqP2ASGSY+kwaeHmBxG80eeiukwi
iRwZsN0C5pEa2bb1SCLXrsPU+A6wFcWBwRn05kNDZJ4z7m2Kdghfx7IyzhwxfRyj
P2lRGXH13Gcnuh+U3rzo4lK/uFlTXjZrJyOg2CdtX+MAS1EjK0ZwgmJirVRwwcX3
akfKBZCtR3Uv6O/FwVlbDNRr6vSacDNZWu/eCXvU2S4+ZAJS3zvMXQEsz1g7e66t
R1pupLSLbmxYahvUxoY8fOIvqUboEgrU/lvvEJNYwzRBqp9NVqEtzh4qgFSPysck
LoWhoGttMRrrzQc/xzMqXPFwhhys6xdNOZITKT4k0k3aOQo2BA9wrPxjN7KcM4j2
AFfQYAn5CX9P08tBwnDQnP3BSrlz0sycRR0HoNTUD/vcwKxd14Ly1IeL/+RS52Yw
W6j2fYUT1P3VqjOXZJaGC5/Htgm27asQEa66tXD8ODlfV7E2h8968oh23CJ4F10m
lW8ANj+QjaV03M48hkvOodSvQJTtujT/J1rCSaWGBtRPfAWzZcQlOHnaLUCknq5S
vJ9zdw9mSnR1hIajrYOHfk6NStxOkjHKT4KmHFqZu6jpHH2KStomklAniCreC4JD
pNttHq3nIqf5cZhXmEnvtqiSq3+wGp0SHNB/Qph5XU+tqNW3UhqYDuUI6kp/K/5m
GJ/Vc/yHUCVP8N3QkfpontFdeVx6wqN/3FEAX38GZaUeVHcVkwTjgkwEExky/SbB
M/VPN7weS/M9d2at0mXFqGx3UA+w+9voA5Ar5KUebDREglJzdO8IJ0VbUqCDeu6a
CBQ/7B6SyoE9FfYga8KOpG0fC9A0RIpNSXIl5g7UTtIjjXC5wf9aOeyeuPfhbnVV
mxcpYi4vI2Btg179ULz8L2s1zDnpjWhhplikgZu+9Iyehpk7abUMd7HrJ2DLLZG5
+MfjwThodHlE0GbfywimnSjRkNjF54iIMLMxVk6349nohvlHauemNl/U4wxM50oR
MpzyX63uz4mNSse/T7xJN6r1SQ0QUG6kO9/U6E9yNZf8E6k1Y42w0A50nFFf5rBr
bDYOw6HRycH94gGZPWkBt2/khNyfAdm7NfRSmdIsW6PGmhlb60MIJvTU4Uf8S2I2
5bCPuxtuxKDbB6TfV8x3xSJNZUsmiIqnaS/jxOvq0kUn4rf+HmPi9vwjAIk1DNfU
/3wWCmbnCfGk0tNViMtB76Qsi3KZ4ilRYg73VGPgA200DQ3qjXd8ptGFoel0RWUf
rdAQhVerrZP2+U7RGjYBQQc787Gvfj8Oceui9Crx0fcZAap/1Crau0BQ5L2hxiWy
OzgXN+L/vSmzKBFCdroEAXRUGtK9RxbnP42ohq/aqMYueDVDwnLuc+w//KAFrOd7
ypS7lFUJ/9NSAtt6prv/UPLipnU1K8GqZfhA7YzzeKf1RqfD/7foQowSEVdFy5A8
N/C63JacU5FkjHkZP98ZX1eP6cWfYq3F7G5J0P+A6lC7gwUNz45rXLfnTQYBaUDV
/axXQOUwxJ0XicXFCEL7IzOucrsK7PyPWzmzpYpaaWT3Yg14MMPoUbPUARkDiahZ
qbO2aLeMFiuSBYJemIUcbB6uiH2zlOcEUgtZuRFR4kiIpugqsB7RnFCIbF2r3Vba
5QyGayzh7N10SJ+jXYz6lvw/n7nL2/aigDqoSVC+EFk45wU7O2XXOeQCWwMZ0CbD
8527KBOPWGdXKvu+7cdtbQhgTdvfw/8lWTo0svBEv8C0tCKNFkIaY+K4T0dj6xyb
hirJVArOFW8wUFY+FVChpcHds79ZT3dDb9i3/p0SPzAImLxB83G8zWw7JgDCSJCi
PtSOTCunjNuj+g7IyVru8hy+HfZK9sKpePaKAM38DIdMiGE8koPkyCDZxk2lvGjR
Lpd6ZtALlVrHJ4mwz9fGONMNqhtmxm4DFx7eU5x+2eUAcpaudxPcFQyW8zjLqioM
v8DEupRo3DDZTWzOFMRmFrtFJ/5UU13jt3WotuzpbmKpEhPf3t70ScdyIhjkVYyM
xoH2ee/6/bqaeZO6E3F7dbKFUthfD7c7K4DfYY3+rvMe7I664h6lMfj3KFDKaXoE
BFH0O4jASNSCBQRLbygSt92OWEFXGlawfxt9sOKM75eYVDuUbm8CY9PHyPB2x5yV
P6EyRYY0UoNTRTaemUaPjEnp4rsPowgGOH4mY4+HkUPoKtuTo7t9GPkjzKGSEDvf
u20RzWU/sAIj1vWI+0PMJbbKDrHOMm9038Xl0nXte8qOroNWe7TU11KiASLfKXd7
sjfxEAzs486ZjGRYE5FBEdIZq++Zu4B5+TgZMxyFGpxkiwb8HueXCVllMkfk29k/
pbo07NqP2SBc9gz2k3IZLrxWR//H2Inmp/daTwfaHXY0XrODRKwh7VsPS1DVGwDS
v4iqiCAtDPptAoJbPJWVr5qbsr10QBPbANup0Btrn9oUF/W8CA6jbLhZhTgS/14U
BMT6t8iQ0xUyTuRVj7086iFNwb3o9w+hayfT2797q2pJWLau+TRxDLdZkS14lYCL
bHafyzksF7pfMPpPwEb0oXp+7E1u9k87ZPK9Aed8gXG6poyeam7A/ia0p2MmN/Id
7YQ2OzwQ+f1LLGOQUcmM9YvZqDg3aElbp7xIk2spSxkvFe7XhEs43msVGxIZDywV
EcRloWZNicx6+MUWjkx1NxCbiLfI25nr46S+x1C082UJf/j114zX8MeFOHI+Tm3e
+/NZf4ICHFRF9Oe7JvYlVbkqX2fxdmFmyfNQ0ev2iQGg7ihhbR015AVwsnXBMHLZ
WZgnx7a8Ti/FGebDWmdKnt9JJqmx5KQwRooFsjNdSe0pBQNy+xqEGQcCd2TMiFBe
EA7ClPLI+P4oAVR3CUPyWfiAGICbHvggk5dv3jj5zL0Gt53Bh98RdfRN5n1ZkW8I
IrIYqsTfkcqsfjL8Rq7h1fv0/ESpM7pfbiHwRGk1YaHlN5vraUSCt8U7jT3seN+l
R7PWy181nW9W+99Zm2/tF0z1j18bRftaqiSCK7B8J1naF/jXfh+O1lALSWYnelbk
hRxwFU4gdRQBWSAAKk+3+ZVbV8Z4qrqxiaLyOLsHE9W2NKZd6kzpypTmFMg3u7hK
H9seFkr8Ui2zMNDDhPKHV7+XNnOis/E6/caZvN0ZQjmkDERjFFdUDVcSZqiefqSl
wu8NLNHH2ga+BA9oaJwmTDKDLaW4o9V5c77qwRhxi3CR2oFDuyvZc8nmT34bbw4j
Z3SZCk1MziVFDiVQ3Rnc7W0lmAYBgDfQJ2OIstax3mvMMxB3QBod0tNcUZLBxydd
mlRN3F16oOVSPY1lovHPEA+WbqUSmcs1Yu/tfAJnDCiZquo1vL7pv50+SmCLZ0Ue
6M8qjnrpMpYTbxXB/6EFWx7k/5KrZ1gUSePkA+wV3aV3SCMXF3ejp81VFYNTlMSX
SDAHvvwIhy5mycMRFCveK0WuVrZFV8SBDDyumsov+POoIyAFcqQSb3Yu4Qc+lYS+
OxuCIOcjSBhawn3oW+2B/MHUayggWmSLHjva+CYGzBi0Fhow+F/dDwFUYBwqbn4r
x79uQ59ewW5K5sMeoj9Plv8oq4PIPhc3Kt35AAW70rIKKmWJlC1sjQCPAR2wEImI
cjb4ctGz1VWkFU4hbxaDSO6aUzA0yzcRhcq9TCrbEMnX7r/Ifkik4f1JwmTAAycq
UzOuf0i6vIUErP3U+/j0dDxBPYYpoTbKzxFZoKhO5EQdTSyaQTe5ueG08u7WjLqv
vbkxFCfqmUWax+siwngF/8TRmldRqzPY7hfMc8kVCP1mUgNJ3gIoT6InKeLySSWH
KREn6UNcKFR4XstJlEUmdghqJAbj4UT99uxa354t/w9d9f5PlexmGQVuBbp+uFi/
UpT0+OjalUrkfmpjMyW4C7c4Jl2zdE8iaddVIs72ivgM66FherEayOdabnuWHMfI
M//jfN4NyTb+gf/0XHlqOsWX77uHBr2TJ+r/qT0vlWjrLwuyYGiock5HxyELwXW7
7nqekyhVCvkUUZM2Ub3nWDoVeo5ZZR86Sqqv3HU51zR5df7C3Z6qf9/Gq4vECNWa
dceGuey8PgfALeFsE7StnLJqqGFzGD80/8P8G7u7ocWDcRmC9dOCTXjDYqIH4uE+
+uIUGAzWMM0GdxMn0cIIsuy+r2DaeZ7UgZ1QHr+oe7GzmUKz4lT+0/9LTpjNXGrX
Mx2jY7ZsAkoNMhKNq6JqoLaU6tSXN8BMm5mGvYcVmza70BrJkCQffNTAxdFe/05v
YuUjMgrVrtVweBIb4apGjsTCu0fRP/ACR1MZNYNhnklNBsEhkpF12UxUikzTo0Wz
AgbznePUBViRvhropN+MD6U0t7Yc/el012rD3MPVFynLDt2WxPbz4W2PVaoTnnKD
q+XAFBQh2ns/movg1vvyFK2x/jjNBtcKZZIERkvE/8ohaIXiG/OE64MXKMDPEkLa
CU6bPeZq45ux86mZulFH9yNOxXVMmDNZ8jW0q330O0bpNPeMgbFLocmUWyLQSgtT
ES0WaZ3UahtZkKkZbrhB4yurdXOiCW4nmmUFtHi7j4Qz0bvoDrfuTAeSpMpI1e9i
DXMkGfPNdFfSeMLHEavcbxNoCzalzGaT6tMvD1yX7c3e7bh1P6qhRkL9+TwXCEcJ
ewdjRCSXrwv/PPmNY65wmCDyDLeAVdOgLtdircEqFj86boIIfi9ZoC9q7uVGq8LU
HTRdPumaM311fn38Xk2AWQUEzWaA/eP4v4vENUNqHwyUnKFQXLCjNc5Y3pr7agM+
/edee6HdV3AEI74+IEeMyLvm6+bDhQ7FrSHEE4YtrQVqB6OdKNn1n4peGu1ljdoH
VZ0Um/fS6SXHrGhIsvuwk24Y6mMeQXX/v0EvuPSVdnE4CpDCUxpMiAfI8XgvG0pu
Ts4uQOc0dQBUaIxiBaRCPBqHG5KuhcGHZPdy7o3Ztiea3CR/MLRkPz/3EVwAzic7
jU/cBX5XlLqNVI+rAI8eUugLqNLwxa/ayAL3fuZbQWThm0+oj5m91cmdG5+6CWAI
z6oU5w9T6oCBCBFIsKhjex8GHx8psXWbOKCCzsh0nU5L8YcXaoKgqyqR7VNSmRC7
zhwESsupGr0aTUgtMdO2lg6Ckm2RpSY8srN4yItin+jqW110cq/kqwzy2yRU+Kpw
Jl0ls8ZgSqlVOn4aG5qO4DC//JKwPNibDyjD4qcwWAump8csdtHC3zd/IgZ51Xas
sadrPz/uBJJggSxMlrZoB3gTD93RQv2WvT9/3TScjiG20kP6T1JJm/Jp5TdPCj9C
ZJMlvom4A+RbHZseKUvnvoAurdwLUtuUCOW/QuxKv9mswd8zYLw3adHZmyENv3S9
mq6S6hVrjmaB8huK4BrBKhyvNl9UkWBXTBUPjScxc+dYyZUTkgPKNMXL3k64VMlw
+Vbjoanonhlsivk5Ck6bsHDCrFlABRM2M//QGPSmEHqxVyOnHiKo5pwnufcTWkX1
h2LLWnjOe1dlY+VnFfkbk+Jn/HjAZSELPOgcgM8SnxQFVduIBfPh60vJWRk9N9Uu
ePaUEjMokEeuZy08os5uWOGhjpCeTwvNa/59wGuhSlNwZAB9E0y68dd9JtPwGzhq
Dl9sqqz1BJL0OJaUMs05/pX4gRyQ5H2XnNUWDHYG8bH/Yp9ckkDCDD/u01zVeeUN
H3PEwceKoWha1d8a9Dr6u3Y8/B0EdSjoRClNturDjYoJ0RGUJarbMVIlL7TyCEZf
ZTCIOW0Kg85ksLIKvtm1nVBovEKgOoafBn7mmR1zSdXW+ioBeuC2tvbC8wXwfyLR
DCHWZhrHIClEPBVue2J7ODEz/O8MJ4XH0I8hmdlg6qTB51QsTtx6AZaaq7M1bIUa
8BrWipk2C7KpdtY12TZNfv65yZk7WmkOQLDcja8NBGZjbTBklDz79hjIQJKn3rpD
K2rAh8KNi0seroD3GqJHoL/3VBqPhW5yx6Fg6R03w2vhDlbb+b+Eklw/WV860QHd
YS1d1B2yZJdQzpS5n/scsRph6CzZ9n7xFpHMoT7CCszr2iRZNEl++lNqdSHJg0tq
heLwTIlf2Axpx1dPC5zUz+9aiYB7m8GwsbGGDDJJ5aSA9MdPlH7AWlvvDxi0Y82e
xWVOudQncyOHerHbsAwgag87Y0Vn0ZSfvXSEjJQFv+IALR2TsY0j6E5VI3+YDuMH
qRWat4sXGEM8qNRs2bBzD5y5+9UJdYcnvuPFB8cGG1iPD/gqp5DRS7Qg3Ducc/I1
oy08gLwGSgxXBGwG+xOooVfsYam/keGdx41bTIew7jTqH+V8gpUALJnLJgBqx6bo
kcVXix+4BLl7URo2vrbJqO+ZEMZEk3mYrSfKOFfeCi5sAjSwazhdVC68WwzylRNX
hLUzlCg7nQoy/4Mpl4IgwKrw0I4vRWEMe5350pK1EzJdrU9SG0TLriv3cqXGkKN7
3oPMFHLtW6/ZHGbm07SPeGCE2b3Pw5wMTrDMGka+5GFfsyzHCTn+YtKaFbX2PwCp
ISjsb0/3RVBrSliR2GP7GP/1Ri6VkcsbfbH8VSWpIHBgo+CVS2td1qXCe653Y5Xp
GgGKMNNc34bPlTfYZ8tX1rqnP5R/GxV0FUZOSK4x2P/daKBSaP7W8RMZRCy/855O
9PabtyS765rkrwkvoAqY5u4FmhJ8X7wJbPHcXXK9+d4=
//pragma protect end_data_block
//pragma protect digest_block
NVGYfxHR3INuZ4JL69BkvuoRt8w=
//pragma protect end_digest_block
//pragma protect end_protected
