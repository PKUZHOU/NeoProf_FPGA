// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
32Rg/VxcbOE6dg8QLPWOqnVj5972K6nEB1A+g6UmOzYNxJzW8SO1xD7PxAYOSbuk
avXg8rXxF6NsQQwKAyNv4vqTVOnW/vRjUsRaGUY2o5CXlMGXA+vA/cYtETXimI1R
0pq3dbc37XG02Y/uexmkmZQoqAcct2CJfyhZPhiuY+k=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 1584 )
`pragma protect data_block
CvBSdVZekbIJgVTvflVhdGPOyD3oAr6JiZQ++5MdMXs8ovsP4chYzVMQJ9S+6y2Z
I6JqVTdRWwSr/Y5yjLxT8oEqzCZqR0bosAU2cfQPvnUbwqbsBNbebFiuRdBjljPb
b4e2lp4TkJMmmeM70oUv4OkufUVeHxvxY/O6ZP59GYTDlpbnRffvKeBN7fFnRjnL
6LZrrebnLBEWHSUGrfc65Sn96wdDd9Sfa4/47CZ/qux94JFAmbn0Xqu7dJjS3Drv
Xshu58qPo+mCcF2NBe1OhszagRD5mN9mCrtsQL88lJ4HPI+ymXB0am6aUfZ5tsSk
0VRSeGgBsFF/jsi27+tU0a1vUu5BVvCVs7BAEEd+wET8vHs3GZ2kNKVV7K5SzOFP
QAHcvPNIn5ZW25y5Mj6jtpjRXcArJcXpe85XLTeAyb8bT2rDx8FyK0qD3aJvb5S9
oZ707btjcNNI0o3o/yv3Jy3dQhSgzaYJqEhktIqgm559xpAejBsMIM5jxEdUqbnz
7BjA9FqAuqvrQddeGHBAsqho5bMgI/J0s5DP6OWhCeWhECDkSOpoM4UpqewlOKEp
1hpJ6f5hv71pfoG2jasChI3udHM+PZZj4nQPCE1H0Evl3QxsNTBrszqChgHRfRpy
9Zs+cNR7WCaERoP8So8yd7vKLzKEY92qr6HbqiXVtYKUfvNlRnZMJ1sLAcUvdhGB
/pkBdQNKgyIh7oX5CmMgPVIWQptB0cTFUlKB8ciiFUmz7/1bFOhWdhdf1nRd1Qd2
f/A00IawURuX+mypMy8IWbESnAADaTsEo4YTjKklZLj5+em/RmirfeA5T+fhWLhC
qx9XvQBc1RdL4SBUY84szTLX9L8qBQXqz6v2nNEetc9Ou6rcUiJ4pGX/6JDRXq++
46KJRKKzXjsB9zSJT3hneUtAEDGBJOjuieNG/qIGi/ecAR6DuI8iQ19HZsgDK8Hw
vYUb29Fjze9NwnIOUUICEIraTHHmcTQNFEl63DIz4u/vKaTOaVOhZmxUGFv3Liz5
mSFfMD3faOQ3LdrGe+e878NkEOZKUCVlb0gdkDJKgKU6muK0dWHqOo8uQjBP4D45
6OwrcFhZ1UZuhz8WoM3u+/mWKzJ/11XXjgvgKKx7U16ysMBAJZWrnPjVZzC/VTV2
Q61Pz0Eq2uQHBGoVwL0rF/8EVS7hlkECh5HHCm6lh3OBP0uHcxyRUMaCRtJwWzYE
nvnsdT5jryLAXQyAUmrlAA03Bc310uU9e9CUDLAEf3PqLNu79FwUU8Zs6zKOXu3w
vQpTdePGxx0tXyykN5Mc+V5eh43sBkr5iZfdaUur1NUs5hoPC4CluWRtVYvm4Kpa
VCOexxfGNc4PrfYjjrCUfr3ESgqErQ9BYw2KzFbFoGu9eX3cEq6mW6NevmsDgPx+
Lefbt8L37+SI4PHFNOL7ZJOMZrHmLQ8fmy/ab4sPMXzcjO/BUJLI16zebq4Agyer
2O1eUFbYnsfInM9WE11cZ1YqhS9PA77QoQ7o2SZMyrRbp3y+Jrjucg8IvNd6UrJ2
qnufv5U/NFhFKzvfcO36kXvHsrlVAi+rpDUkVPoeOsuu2Ic7h/qoSaMWNV3ESJQu
78fX9HBtw0iSbeDduEXazdV0EWucFPca2x/eXueok7pfQHRVwhNkPbtHQjRHk88z
uVmrCcNKlPixeSRYhTSGej9sI0/Frxf9/yLNTeORQXiYDaAoWGdhKa/kpmGI1fKL
qnEk/xvFclFPZO9Q+R7sxqgANtOPILloA3whlUr0nJ8tGkm18j1LlwVMYnyGtg4y
CpHl2OFsj2X6VlWNuIyvVy44QMIM3LUIWvNWCL+F/Usj0D3iVtVFItQEenHMjORd
mV0wLBJlRRv2DRWhgWXMz1OKX0NKrQL+wYnkuLxV8SnCSy2iUDYOgPbbPXeF30Cx
hPGbwxzd5rmCU68fcdm7QsrLdWmomLKCZvhlo3fv8pk1zpcqdD7NFrTqb1jw9Alo
T6VY6bdncLsGegnVi0nA2lB+Bb0r4lumVzTSUeYOshRCL9nckdMXlHGS+pxeORHm
zKG8DEaOSZzFj4uEsmU8FvYiIyybfgJ4URIew8yOCLCtZ5YT0he2LjTBvb/jX9Wr

`pragma protect end_protected
