// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
EMDCYq+LPio19Tby2/huMna0Qc4oIfj9S3sHDnC3nAoEO/RJ12OTATxRnLqp
4cj3/tcamp1vCVrblQdfyHxIraKQUc/dLXKegH5i5hNNNTonyu51ku7PfUtE
U4bETAy1/mt6WC5/lRYvIWbs5tDboYHspLLe42MkVfj5dliGbZsYtlFaB65R
Es2+VR6a/or2WCfYva/oxztGpOfBifU9rJGxzLSnoTNfXeN+I1zfJ7cyHQvo
jP2AxBIzwLQKDwK2EDoDFfM96HXp5tHOIe/sfZGPqc1vl7E+rNYSjSzkYCjR
JIqWKzVmi4Q2gR2EwGhxZLaM9wi2Qoq3zYGK6KeF4w==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
fK+zrQfzZmjNj/gf5+xchiPmWjyN3+4G7bI86O+MWCCOVF/qZ/SnYh1hWvie
Fk9tcAHfCYyRlfyb/QVHuO5y6Aj9rYjtLZd61t1fM8RiT70J4OpA3+eT+cLC
U8axaAoBoCuOFD8qnD1aQQ0PFEniBDouyByHwxbvwg75szQ/c1tAx7am1IEm
8WFcNoMlEycioC4ZK0loIVq3TbpdlD2Kvwi9fYW4plx/TaPWxNU6Fd53UoNh
56lVZBUYYukoSVcJvvsHIsj/NeOHNxva2v2u+ahOOGFgiKroQH1WueELFCLP
28nylNoxf+Ckz8b8HhMP8AI2fsZAcnd6U3BYk/ldPg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ApKz88NT57pcDl/IYem3bLZKPQxiGCT00aMTXbI9R2eU6pu1vOskuV5VtrMT
yGeRBbrKvEhVJkm13IesMvLlYNo6z4aoatARoi4jQBxCffUSGGioPdhRe0oc
y+E44Cv3qojOeA2P5iyQXyZP3l/BF8tXGt/Su7saNUJqaGWgVCz8Xu8IIAKw
JfDKG4i9gGt2RsfFw92d8tyUjJjIKMwFjjAsCubJF4QuhdcDgnzMEy1rPD4R
m0pc/WYmYKuJsMMfWrMuKErG1brQO/o1sGcRf/y8vgMyljkv+pgWXgKVKoz1
OHehx8dZmON8pTJuLKyMglwMWUpCqxtCWiD49FXTow==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ZHTUUhOYPOyX4onSFddPW1nk2ZvoUhLo89fW6WTXiXFf6m8+BlT9fpcVAxcz
erjD0FKd7I72D3jR4FZMpY28YyenxoiY+DkKqRyEA8nr74tBlyepzUtE0cxA
pIeNB/qUt0T5FOclPwhaUR63Zt65jy0hmPRa5FMVuRB3uSXwojk=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
uiuAQAoCTpvHWNZf9q07zlTJXilyIB0/UeY8mOr1X2Si2Mp5H4ePmtBiFsz4
RpXrUr9JN+9m9HjaDppKmJvFzxZrBubsZDeYq7ZJmTTs6SGl4vK896SK0szc
aNBdSW+z//h85oqwSNuDNzzKYLdfYXo66H6lvCI6r0lqzenTH1TpuztJArPN
IXDQS0O7B4OgyJOnPfAFhQaIUnZVxvR1Rn7TcGZWydxO0eqp7KwTQfInodio
WrCQdJU8SneYNSxwQJ/0Rn6cLc8B7NKzMR95Tut2/XeVJ22qu8NQgsJ4vB6J
8B+NA2ty2GkuhF886N+C/yTN0tpyk+4+1y/AOe4TFwh8mXLQMXIU3yT46HWa
ezWkzo27we6DcYgUb7y9JdAJEXoGPUF1MxWgKMcMOxZrP32Vulbvdxb0g9sP
1Z3SBTVjvdrbGetsQ0Ul5g0pwKWQfNbBcLpNUR7XFUWbdSJNjj5e1SLptO1f
KWVKCZbz8g8t+yd63foS+utg85DW6dTn


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ukL43FSTFlcFB6xGBI7jwW9r/fPpDOUwshwBNBwzdysd/xnAqL2Qbxedj06e
EfVNjoElZ7vMy4+UwAm4qZmYc0uo9tkVS6ZzcZUOfHPYORZxF7dJ/qF8k+Pm
/7VKyrW73We50ZSIZQCb0DBRSFxrqy78uLtYciQYqd7R07l5hR0=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
a3rKwNGgw/5To0rH/ZurVuw6UNt/hmKFUSZ43y5SlAGC2J8JX0Xx2OO5CKpI
HtvZiW2U6NlbXJVLtgqDapn/qYG1JG+B63Z13xO1oh+XQYiWsH3EWuv6lLZp
KFRWreaqJSMtVJ6Tf92h3gICKr8OHS43ramq3idmklwzPlfsxSg=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 21072)
`pragma protect data_block
iSWlhNIgm225Q7j7yfKfx9XhQZCfK8jSljf5pIGLUV0w707/vavTqOErEKC9
BWWNpj2TKUuy4L2Xvpg32yNfEdtMFimLj41FAoItaZi14QIToTeV6UzYgU3O
zsDnnoLd1TtllCLxt3mbsX9roTb3ThYjzD2MetwyxbZWDdxlGIClF33tjNcj
iBV2mQH5mxXKaZDU38yDt8KmDd/1Xt+wWzBmSaNvJlNIFSU/OZ9tX4AUozqX
8xVW0w9jfVNlUvYbmEL9LBFdY0ynd2ZbvGh65nEMhG7M3twcVrqbzVTLIsw6
DxwWZ6A8H/z7zdh4tTX0wR8np+zqeiOvcadKvBqCXb1xexGVRMnHfHxxhce7
GOzqAorsZvttdh6z7E66SMk5PA1D3t0F+PpbfYC0Xna7NHxcGumqYuiJSccJ
PBQhlLiSJkE1bmANGzjjvwmeMZoxMQ+271r7e2SndlP8xQ6H6PsWvbfLWMVk
khVwB0DEWOo8fb9hgVmmRXBQI19nnWa7LhSeH9XAExbkM8mwIoOgHSr2aHDe
hk8R70JEzLeVtWLtqyQHC4uwORecwlb/UQylcb372hVgKlWX8xBHA7y2YCtZ
uPwkxGS6UoqT79FbtZdW41p5j5c2QPRz9mUY8DpDU8AnJAXkj2sG+LTXh1N+
cehMwu80BQJFlUjfq7S4EalIJCKPIrz7G268bceqs4dGKntK4igtWlwko+OC
us8XATLTPZ63Ps4cgNyoCib3yKgKSvKcQgMRq9HH1nHWX3ZtNN3iOlAJzXC3
yDhRXi8wWEOyYCMMVwlUKGtRG5yHvDKmXpJlzja3ofbG6gq4MwmTS+vNEdIz
D12x9m4OH0X0vFkyQ50g9JlTIlCOkz1LA9fj2V5lpy9eNMYnqOScM2UzLllN
PuRD41ZKpimHozwmFIU5EUpL89yCkT9l6QgZXlpir6Wm5SdsPynu1lGOdgN2
NKiCao7YT3usizvemHcfEm9FuGRIAxxz5QoXWjAkqs4JB033wS8rxat8phmB
ghszITm6nN8T+7SdAL3LH+LMpxh8DTBGANMB67aQOdQZtPDlujRjfMGdKt9t
H9zO/eaq8VCVSODyaQQ9DPuUXkgDUvGfyccgZUBtsaSWxX8MWsdinIbI0CHE
2JBL4/OC0mFhVUOFEfbJIANc9A9/Cn0ZNCKj89hEeTiIcMlYdyvFRk0tGrDJ
2C5bQw4s6+Yg3TKQd8L8uYb0InrY6+kotP6tvfoJYejhzSvNXjP+eVpjKa25
3Ue0mchKPHh3S/6iLx8zpF3QQUBH1RJCQ4oeAP3QqL71Cl14cLHYWE8NUZsd
uAQfJ59JLhDdCYb0GgrhFRxEfULu5gcC3y3CdExJ6UpQH357qezbDon8MH/Y
VmBlGgkaYnUjsPORFCJTNF5/E/rZXFgs3Pd9CxgxBJxzwLU9HOBnNet2UD54
uG/02fUOWfNopdZDxh2MCk2aTr5YCaGC/THxvFho74UMK8aaCORNQucTvrkb
xwmhnq6ibI9GNGKfJnb+DqHVc9Jk5Hb9kS4u/TAQtIwJuhfQlKW8X02ZFEct
Rt2qzydmh2wleUIu8HvjBBSlXvA3kmDIx1VCQBGkJZvCD9QlBq5K+671Nt9K
tWvIAN8F/V4TBlOIe/R7jw9aQWJuDCxFH29JebOCxRREjMOzmlGmwOgQw9PP
vXwQUUY5SiMWayVYGwn+F6/AE0jGsSDCWogZZGUv4MfjhcxhnXkYa/LR07V/
+2JKSGuZUDxFn5MYJb3RrPwuCVMkVCKogK0Wbu0KGB3K3jdCx3hWV8RBPFP7
aSF62D5zWF8RHrPhsJ7YnfzA03tTP+sPv6MlUZa6ucgQH9TLO3MAxGw/axKt
wOwTK9fAczzkvH5rVYOsDqXPRi6oYAKfUMaZ8iWSIowDrP7xKKjq0/DhkH8g
ouv03GKXw9vcPcRLb2btmbxrpuREsepnu9AbBKiA48Hbes6fcM/HXpx+FHoQ
/oCiTu4XOPnZuxi6Uifh+lGIId6KLlefUxd7ISln3IZcmBC2EdiSdNsDN6vZ
GJxMdP5bUgoutRW8M792sCNI7zF8j/4Bp4oExO14ok/yvRrL3JC4HsnmWT98
3obnjJdvIIF8UJ0tNb7j0l7WnLPipGSlh5V0XiQnWoQ9S/b35xgIhNuunu+f
LAX73jeknnRgnWRL4Q6xqERIJ0b5Vc7A+Fe/vLI70wnaBzWzQwFRBwi18Zrw
8RX0vdUi+MH/lsGvIBk03TWXtq3f+evGll7gxhYnCzc8vNdEGPbO2gUJWrhg
Clf80qT1alI8WvPYajE4bECDzdxwIO9U5uWSWkFgz8xujGqGKO4Y5yjG6oei
hCJQ3Tcoz31KH+nIOrEj7Q/U4NqQaVuRWsWJ/oCVRNcbmyyuAQchKrgRGU65
uwb0v1xEfPeGN4p8HyJEyYy/MxIvtWPdsWn0uvmZ2GQGloR8X3tJva+mGGZ+
xfcZtlORtteM/P4CEF9K6d8yenuYgUtFaLN9dFP2d9aoO4P5bEmdHPJ73hya
8OCvYqmLvtdcmeM89ul1zUGIqALCF/axD5jbq1tNaaRX9MTl3fiZTrErw32n
Qf18OEehXCtfCxkfFzusTxeqSu7LblVT1UMAA/uaqrEbnIGPcntrls2lT62M
ArMPQmVVRu2EOAvGN7viw4+6SKNFKaeJyPw66XZUDZJ254HoxoXjvAfOQybs
2ibCuV26bVCVpMxIu65dcvBHhWYQzr8aANLhti8ttsPDtkwUe0c84d4Uj3OR
P46KGkWjIEYhMD+LVxOYz8FhEc+V3bINj2SRjSwZi9aTp/BPE9CiurxmhAVb
pWjrZW7I3IzPKa0CUkRM6lt4rqU/tHd8ja/Lpy9fae0+rEU8u/yKf66WDzKu
d35xmcykOhC8UkNciiN0vSAf+T8TluIUdayb5BhBtLoQi1g+28vWNLO3EyCC
GYOKrjFb8FMk7/U4IDCk9E8OGG3QuZmseW4zx+O9w7gW9NAWNYRdpz1RiNGS
vIlVhq734f60wrXJdO4HvjhkR+ZUomLLFHLW/Rg7Jk1x/r5t8hs940XB7ouj
FFD/MeFzFjVJ1mbmorn++lDicCKSTePSNYTzZVhpZOI1xZSXlwf8WHwhcbEJ
Rl//iwNz6ce9uTdTIou+U4COqtZsESIfxruQpzdRTC839zv5bXF/AmVSGnLf
9X48az1LVtEYXp8iSw5FybFATOlQ2CD7ahbCBewWmjTVhM/I9isUwYIlhOgU
iLx0Ub/lywzKuJEow2X8g4X9kpWMyPBWzapWKRvXzG7S9xESmMalDOpgWxuW
BadzYBLmGLG4Mjub3TOmecEcWL1eY08/1P8PZPPf5dgvxMxlWNtKSXek4mc5
GuyT9CFayt9cVQx802XR3qNwz9pAszyhyObI0ezzr+A3rgYr8yAtA3pw82hU
995nrWq9xL/EqIysGM9DRyFsZRIXTG+rESkFM7jJhbRhUOQXk0KpQ882ghCy
pRueAKOUeGceBJJATQHVn0AWBL1Cu5vtPHqvzU+2bzyu2Yl9n+wcrurNmcqc
rZJwQlZRY8/jzMw0JZPPixmenrivW4xi9VP9Poa9mNNOijUDaHdb+wllmSBU
hgHMsqHgj1WiaezKkKa5bkv2pNfcGuty0zfwiGt+NfX1hFsf+yY/86U1HMPJ
08LuALWgIoLrzoNPg4GkWbAojX7/SYWUJjzkwO9FWqqitHvRBeCdYcYT+Hjv
FWflLZv0fx2fiEDIaACIPedWQPD4cNXknpD9nVPb8huF0lHWgZwEedJ2D1WN
P0kI/d4eH41oWGciMtucZUKrEygV4L/+autqtosgITlaq/z2xbMoByuFBD94
aGV4soP3GDeeqVnkv5uwJTer/r9pUgwxQnjhkPTtomJVLAepds5Ylr/6d2Ni
CHPe8af4mOIZz5zJm653GmZ/tidRn0uzX680XDXfN7cVc0N7XLefIM3lIYVZ
GNEXQYqlFw7rx+XlcmBOnP3aoNpUVp3Rl/+LqKLwU5cFj5jAetNRjFqGn5gj
BkHPX5c7oWwq+KPAp2dx51DsePit8RSMw4DH0wfFg0Cy1X/tcDFMlPz9r4Cv
oR0q8rrEffoUef3kP3+1zRdnvWWrpo4Sp0Zv/ofcQvRKRHomSoY1ImIZ2z3d
zFOlwfuQ16lk8ZkbIcLkO9L9jRYqm9I174AvijVQAjo9c2BJMQXzx4+/ihX2
GnH/t5AgsmfrEffqD+717uDPye01WTtS+2ue2F4crBYq+Iy2b3BIEncjoCQR
VXTJs2YcIyYTsgO3hNwftL1Kc3jtaJR72/1dRpj9PIqL2FJG/h8qzXrfeiDa
fvESDupsIMZO/IwTpvnSr1lq573g6RyNxauH9jByRJjCD0iV+8wtD92XkXZt
VTcSDCLGpcLiEw6McfBlst864NXZklAyduSkaCPTH/Bdw7GCeLmXjh7jSSKJ
lQfoQUZcot3qQDgwUvL+SNdvVIYzxua6wEHAqZNULQ733iwzmLGinrMyqwHl
U3fV37JYB/PoH6K6bfK4Luj0IR1Cm3zsF8JV088esBxCrduj69JLWna9o62X
kIQ0tcUU7C+3J13gFbhiP79GNMxQPXR0i7+nRPpU+77tx66d2CQwfW6NGim/
2OAKSp89ecjOOhr2FHJq5APCfBs7MTRI6O2T2Ix/Gn+0C5SifdUMHfYSEMPj
StD0jznxO0mNwFGRNESfbiUa07+ZNYzqk7TbFwMV5A7546gC8WhGbZOJZeSv
l3m8mG40DAjGF3GzlwalA1P2lDxtsEryRkTlfNKnZdofOgYHuj1iyMs8Hnao
xYMhHZnXcbVL9Y6MLZlXEtjh8ydmbLmmmAdBCIcwayV9gDJlKsaT7dX8jEXz
chJ0StRKJdwXK2ehib0WFH2XPuBL5W4NpzLXLtXWlsdNWV8g113LILxRF7bB
TCchVY2eJW6EEMaRz/v20l3BVm90u61TDyWaXOAX8GppR/cT7axeIOig1aLF
U/NVPg9I1R4qdPaPZLPCys+EYmH4aFsp4x1wfQY4Whir4B1Y1edzWvqn0or1
8BjZMGZUDDOCz6p8rd3ZVhtCZ0dU6lRQmvZK/EanffhdIzoYjDZA20HyTa3D
ZDoi7GmG5KUTbbbNoL3ekzemv0a/SIFXUfOxBbTyU6xYd9iKr3thkg8A+ItB
dMrLjlBisjp+6NMycmN0mTe9mV5NrZwLmhhzlUQy23ZnjCAUmhceQSbm1Jt+
ykTcJRVRJKHRbf/tfDdx8RCufxj1RQVQbzPtQSE51ykyQ0heZJERO8sE6GHn
ZCAls8SH7RJ7NibXextHXQ4mOGozAojz/1IyYcEgmDM1uK13sYGTzyzMktyU
Y/selZNBrc2lNylSndRSZPNDIrbVBMZYnfgkYaHpZGjpBS95t7N7yFAAsIBO
V4CSR277CKJ+zpdM0XP/gkEzw2dJBsbLyp90QnQKgGGWl6nlG8zj96q5SiG4
6kWSmB8LOLDNtOYB+1FVPUJ4tIizrHTwi7yTY6jbE/GaBJ0tq9Ff+nkpApM8
QNDlTyTCIxGgRznAfwdQavUJ3FyGJiDnyd8CHBuSvfl6/nvG8zf4J5IAjdbA
fLum43aNFx2EVAJkoZo9MZud8zLCnJODXDzfqwf8Mp8l1uCFvBHC+rxKFanp
s3VIr3a4o+dfRsG457s8nt9UFL/andCUgwVHylhLliMj/c+7KiKpccslQ+29
gQv7NSQFn1uqjcCfbDvXZKNGg9Sse5Qlxx2KqXoYDUXGR4/7jLMB6XZPPPkz
4bKytRfyragWkhmCikOPe+M7edOo3nJXWT459sEY9N6H00U0GitwMzWlyoRK
Uc/+xCmlMCu5l5vyDRDi1NznNqzibZfHvPMY1xeiz5rMRgRbvEmzq7IG6ss6
0PJM/qo0NT0WjdtdivDfuGgxUeoS8tRctFCy1gelTifwc+cS22S1hCBhZItA
QTJ5JVIK66r6K1kKZXBRwbyroIQ+eta92mmUTK97Rv2E1d7JQ/O1pJ/Mc0P2
hbjjdSXn6iGRBSfdGTbbgfS9Efu/qu/K24d5wDW80V/4wdjdz1jwlclkHHxh
pU2vjXKb4oLhkEo4weHm3OXSV6mHl2VUVUlmYRHh+qnxxXjC0KhXYQ4EpHBd
EJO9n6SYMmis1u/30PsAlQKnPx6SfhYz2lW9v5SNYIcqadTkgb6BWtBi2NuR
uHZYZKKfvyU5OsYTZk4dDDFM3vKecIV8/VX/cANtBqpcBgFsGeT4fUUqndlZ
SlUQRHuDhxMP2s9ka0H8nUQbiLafonm4VYWpvlE0PNWv7T0hC4Ay4aiBkvn0
mSP7bvtenhwWQ6bJSTHUkE3tk3N6enLkugDTPvDkTYATMwpuEsI8Z15sx1AA
PJaRGYggSkYai4zjIOWvvjhcZPInn9aP0R0IYngL6y/MBtEZq/wAWvdRV2OX
iEyK4DzLfqYWFbQUNvA42pcLpuT7kjw14OfYw8Qdm+zSW6H14G+CMBIazGEU
nAMAnkWLEsh/WMrDEx47UaxzhqA7R9EfZTi496Kx6+X3GvR8T3UE6gnFOIcb
o8vvfrx2dFDSuMgBzKgezHKYyNJXQKcUcIyQ0pLBMjOANCklB+dJ5yjBinJz
NeSLgCI6zcsWrg32/RnU7May4/GJEadTzrLtWK1e1ROb878EYn3tQTr/q9at
v1TSMOksSjUV5OCwDlcMTr4UHLNSFE7EMGn0X8kBfOj6RFcrZKphQYGLsNfn
ridLvSArs+YdJtVDy4qJ3ITPqniS1zURnZHX/K3Q4SICpwQICcVaE56qI413
PeFSGy6wdOieICqfwubLvOD2Qlj9Hkrl/Cr7vfzTZkoCZOln9IET33Y/X1Nj
+279xVxoAwIevKLrpphnHVmyJWSPFaG5s8OWcNtuEpyg2YmR54CNCTIC0FjI
4GksYJ2xQ9Cn0qkgZk4iBqKsdvolb7inUB1QutqQcXOQDyTsietVhnsxwItd
ICgWzwyexyQOmNWmJb3UzsfRy50k7UXlXIoolROWbjh/CyacFSPt7iiR9yDE
QMIEv2FXzufPxYP6alqutRDUuQtEtVSFa8g1i8ICd7PgNUBxj4tP+dxJ5FXq
7hOLjOXdP5tavuIqGw857JbFywKIXMLW0TwngO5L7pEKfw9ZQmBKA0cvN1+V
ZAClJ/7zE7N6FacSw+VRvkwBox3V83XcY2JfHX0NR0HbmyGA7UMMjNVD3gAj
VEZ47VVizzIx/eVz8sphPHFliExF0zvnadhXQbXxWbMMhsCWX6SvBxrBEY7V
4HiSMc927nut+r33ttvP/wC2vVQxa6rORJAOu4M0ttbdXF1KiZQFdNAxdAgN
CZhWphuiXlFCdIJbwIy6jTVRVPH9ExHK9Oh6RBESsLOqo7N7WxKEVZWtQv1c
g8awtWY7GtnMe1+BDRm+VoW9PQe2BRjuPqOBZTGzeBKhVUBRa8DHJO95VXZR
bZ3Z5jVrvgV7pLlXLWvRycB+Z+rxuiJ2uzOw3oEV6KSwzaHSCMuVnQMPtUy4
Rpt5OzxEaHrkbi3F2N+jmKeyYmxL9rt7UV2il28ju6SuQttKc1NgDs6iewRs
xaa3aUdpd6prTw1ewPZ59em+ENdyz2jFkf+2ll0TcSWpDD2miRMTFRdaDzr8
3BmLryGVgZCfkTHhz65Nxw9lzalnrK2Y/UNivgXDub1fZ6gpmhdHyuM+kA4l
N1I9LXt0bcak5i8o5yBi3O610JC9HmX4YXgy8RxBohMkSIweOlk8MUCm/ymq
qpDWHUAQEXGhL69aKrgteeH668mO4Zyy84URDHEBxFsaBRiLocghD7RGvJo7
TvUeoId+3qCv81QuIPyVIXB0VF0yfopnYOwvglR8QKscza79lik/fQbKDGZ6
x0dwj1OhQXv0o9YKa22LXUcqGc/Cruysi0gzs5UL1ejAqH8uUmqgKWTcEglK
7XMPzRVohF/Haf/jBCtvLO/txPdCLtu8GquBpKrr+9/6sJ1sqICYMvgBT8us
F9igA4UWQ0kMwJcxuXBPdYmiOsGjqf997YIaVGTZQX24hsS/6JthbmGEoEAG
zzO9xF07cjqA4KV30r1KT+eBydfZH5mo87Hanr383xI9tCbUHUT5yCpe16QU
0wfYL20R3JDGG68rt2KPw8gm0OssYkBQe7RPsxD1agEf1Dico5eBpPi0CITQ
yb7/KgkgJRkurfLCUNW/a8w9w5R4x+o3FELQYXdhe4fqbWf8oyyjGs5NEVnq
wkFLWJjFMzndasQjw4cSnjcM3WnJIo9qjtEgrZBtQQjc/xrNbE2oY+e9KxBk
g9pWhDyFC2BikX2Ga+T5CK54PIMrgS+4TX3shjvmYg4f05VAVPLEuVxLxBe3
RvLEJW0xbltHbuHc3C5Cuo44iRoKgntD2eKzJ7xXtQkhI1MlbPJ+Li8HOOfd
OUAH+mJvLjjE7Lwk/izAaUGt+wjJ6BMMihOiZdBU3njJS2GHTTEVsrEMC3wg
Br5e1fLzJvhJvc/Yu0FY4SEBbGjUUUMRHXnX/zQSpSrT00p0nnQVt4fSDni6
1z+52sj7FnLBPj66z/3ZnyX9cQRn8jRCJSYz7sKLefkGGleQ8s4AoAqM+r5B
dLTKSyqAsfykDBTuHVkXtdJI8Gisca/+j4mWScDQ5Gtz7PEBCzYOvATdV1/E
3b4QoM6QD+vfqLJYG11TGtRxsyeB+xKZ2XQ1fV/4TJkWujy9mneAFvx7/Si/
bTxVZ+WHYX+n5stMYYaNtmOqbsVv53YHkoeqjMBTlfngosmttQyO7Y1qy9Xh
ZjI6FYYdYKALZuEz7zgsdWijRVVvNTgi3Im+6sOMWcqi83NKbiLu7xF0at3O
1QaN5V1EU4ijy8zbe2Xm6axSzHar4i/YOiZde2k4C4a0SZ8H1gNF3bc/qGKT
FgS2BpUtnlQ0HfJiuEIQPZeh0SvJreiu/WRNrHPMq6MoKXKEee8dt35VmGgj
FF7xANJa4tPMABgF23srLNstMVIqd0PBcP6OZxABzHcwKfdimsNrdmdcBYsG
QasFUc4wgqkYOjbAa9FN8BvgCwipQJDe8orAY9GxypByWsVkba4aSR4qwrmJ
e8sNEgbs33VK7HVeYehxWjyv8+ezpKyVZuPqhA8lgtPworWri3anzvceBvFo
/qDZhLGQiYYo8KK851DLvBrg3or3TJMcDHaIZbf5vsLMnH1YaJJ50Iufksiw
fO5LJL87l9S2M19aLveoiGv3zd3BEJs39IlXMIF8pXT+LOSLF2c9xrTduzOr
RAskqyHReI1zELijZ/N0LaDu5ZgS/pBY6Y7Jx5X7K7bmyxJ4iOOz/2yRXjKU
PZLiWrMY03pbCXvgOBS54jw5pPOFuG2+x+lKAZ4XgJjJaTYz43wZDQ3uZcqQ
dWd06DnZ39I65qRhhlnR1/MB+4+9z4QwR5HpmKZqXBydfxmHbOcd7rkj/Tmu
Qq5IQhHPrvGDYPvl9huDQEvnw80fI9quBZgyeLRtbqkEaYe/DXPzpHE6yTFP
OwnqI+qg6ZPxIBbIbLyilgckgXoUS4d32mYKMCegsh/CQWbyOelksPiSO/W9
xyAxBWYXGcHh7yii46G4q+1dQ5wZ3OkPBq0ma4ro2nPnvYmghrErK+sCK1aA
4EZq7LTibVgIDqcumuvjJzbHG8B5kezmA7dzUESkgma1YCc8wEdvqZIiFF2d
p7w0KrR1gjlsjlF5ikCyp/lPxk8Phxlzhkq2Nx/gpia3ucpxLK0e1jv/iNuH
B9bIH5KxWzSmvqAGVexuRfImkJMQDwhwBd46EoLz2/4uVnUMRNsekYQozj0C
GLnAKhKCEozLu7CffATPfIFQHjyDLUirCF9foc0a5fIv+Vpqfax0mo+kBQ5f
sED9zHUQdeDYvMUJwLP0XDw7V9TAMeX1dtB3ETSlC17+Xjvq364ycbykl0Wt
TJan+MSzUMMBloyCkuaYS2eLOd/qsI1J8iJBS4qNgktyGD/gG/blrvRMjJep
eviZ7VlWQLia6O7IBb52w2HJhrZ3MG5un/SCjWpMz66VjklZTlwYDOfBzdCd
qtu3nvzFsa4JoEerDk3XRCD7W1fFftUENqkxamZKzHycP0hJ2tqz/eD3DwIm
BFoWt0zaZgWU5XTUnaIUMGLEzfjfwLjGoOMxBw6SBfZke35Mou1fCeOHbALr
OBCSapJ5bjhjdzHke265KeG/TghKYyOL8mFLCGzClkSfZA+WO6Dz4mzGcQYV
v/tfj/a1p934a94f295ARecNEqeJMBSlu1qy2OB6V4UXUUiftJLRXwtgl139
SRYfH39H027A1rk4Mimgt1JGxmzs5ChB54irQpcq8qbeiLAg/TERCEBT+kGA
GtDsBm7sjz/RRM3N0u9ixWGVy9+H9T9wLR30xsEtNLpYSnb8arPdB4UUoZVA
9sJpkfTT63mI81HosdeUolGXg1rZktKdRzlFq2W0SRB19RxEIjBYs6C/MqAe
Cr9w0jm1ykmvkhy4cIFFdeHu19m1+cbWifCDbBd3m7h8JXeuAxiogIf/vI7w
NFZawBwRDCeT7oNwMIqUV16C3AwsyeK+vnMaOJo83zWMjyLDChh0gNKA+2Hy
aWhLTLsTQNbCsiTNht4I0VcrBtwhG1pqB10R8i+bjcQ5u2/vNO/yWHb8sBEw
xl8TEnEeQkqOJ0PwX8svDu+f2b2Ty/hYI0BGKnJOJmMSexd2L+lVDVUsbnjY
I5Nk0rBjgRsEFnWdjyAW4iSezLU+wqYidT9K88ETMSRsPvOT3H/nDUz+ESz/
7bMSwJ/Cok0vAJloTuj2ljTvha7bX1kEiaat/DEbt9qWe8NIBB69M6m3qfnK
SFdHTPtXTlPw5TC8BO8o6DKtOsRW3e4NHZICg/srHYCsB8WRS1G8ULyMs/10
ad+qk84gZaxcHephDKMHn0GJIiZPj3EZLCy1QWyx7ZAGrE4KbXAHHoNE6hoT
qttn1PT+Q2iV3Qo7O/8q1Gt7kzo7vikoM9PmJ05wH1cx1e1YY2yIlxPjv1ek
W0KB5XdzwA4s60Hr+L+k5RnPl2Xsdw7UNW613tSW3zKnxuiqLXDZmD81wL1z
VzehVWXFbmmvI8rAaTkUzIsQycPhpzQj9Aj7Z0TzlUVin2nBrPwSl7sPXNo0
qd0+z6Yei4z6j7Y6mbXkUpLqDmlwwnpUl0wiDQTasHhzP1J+o6CDFei7HdFp
aDRq+T8srDPFu63sYeP1R6aq+V2q5N7BN2NBej42tlAS6bAll5YSUyWLDrAm
wtxNmcQHhP52VWHLhLyMl/x4X9U6OoXw0e+aGxegk/Ro71+I//FKEx4jMq/1
Z7WAbwAHKXJu3osLrTgyjF2wnoBZmiHweSOM9XgCvfQg8z8M9PrUE7y3UaVZ
lSbTwDjktiGC2VuIiQfu9fzuTZTn9T35Jq/uC7tUtRP1+DLV0VQMgISMdYgx
tiP5UeOBucT48dQGejC8EpkZYj6mW8HYLINJYBn/ED5BVnRU4qc7OayDEM3e
P8kgagt8brzSXJQaP9QXmgFfa0+HUk5ktOEIOl8ipvFcVHsGADuRcD7NR8fB
NhlSY+XaueQRMDWda3dIEH7iOUDGfnCNBijaoPbS+I++Vw9gufH+2YuiIlC5
43edY2dRU4M/neQ/AsEXDlUynUDM/kT9YqMKJ+1Cgt39EbPUU3XWWihCDemD
RmhhtFtrK8q64HMX8ujXGFGzUMHzg6e3LozxBacxVva4mRJPg4EDf3DqkbRH
lkRyDZ4LjqA/RkByLvAG5xoESsgFjDqdP9/NxCHdX49cLV3b9UZzvtyTDhHc
hSsqv4JIcHSZImpt1/CN1gR4jpG2iwbUHd69xE1/ulYDpDGWi54Ql8WLPlUr
m6ctTbBktwsbT4vRRJsyeopMJUkFH4DBEzzwY6J9LXYwjIgq8wVK9ILQW2ho
tzG25IPQIpxRHzodfJXbSFNQHr50O6r85kMmRLCL2KI49ptP0z2XW1MxxDRd
1DB9pbAwqP1MPZKBH55s6s6xXOMHuaOb44ZSy/+Ypu09NwLvJmbKB4tDqhVW
FD2xJ59KrHd8mAK8ljrvxCRHE3PJYs2L8GVkLdWy9cfZUS7USu0j2sXpZ5v0
0RS/gPz2Ae6bZzoAolWGqnb2aZ9biiPEYVBrqc6mVQJy5dsV0bXI0oUUA77x
NJ17ghm0snzHtYeJB5FUiXqk9DTiCKn8iNv4ZG9BXtSkdQPAHyUDmREvfOKM
y1HH2YosVkrNBhhMjN/6DuKeybUjMvIdRh6WyvKmTciEQJAChorVnYjjSF1O
E4JKunFV4W6Da9R/ysjaGNeIwnD4KqL6An3PKeO+LsuAeSowyIwvpC7hu8YX
LdKB+YGxHV47pno5bp+kmBBuU5sQ6olsnAmAWM5Fr2TVIzO1LyLMhoFIO51V
Dup1aX/AZGwRBIID2CQsh6TgHwWnoW4cY5fcwJ0Ip+NoWE+cPAVJbb6p4L63
yM2cPOtARH1V0T13silr7wVxoeVI2lyXAtS7LkJaV7R32KKSltZUCkgFUQfg
yBvKDy36CEDD2rDV0WGuJnBQ3J5tVOTqyXbIiaRFkaiScfooEMzcl8020IiA
TRXOqxvxLMFnGRC34NA6PXrDd1CwcfLOEx6VHXBMsu1rtvmlE4oteukENj1B
jbERCelDRRMYZk2eYAPaNtHQMUdDEg0ZSL9TnXquCuEINLsmV7aPxxRg5CLz
NqbZh9J23OZOJPi1tPjwxqdMFofQfOeOitsmWYx0D5tGn5BcTdCyPbeyuEkT
qt4+jEammRVmafIDSjSJmwJ4M38J/52n9iRuT4sbBRlnQFjsR3zJTb5guUbB
4nXN9ckCS5f2dj9J3nKEIwhaaiAYScVVBOeb1LxPpDAyj1D+9wzhGB2yikkR
OYgdLZRZsjgyFC+Qc2Z4jBzPaE2CMruFOJIFcAcQ9ingVuakZnn/EveddBAE
4m9s+Vx/E+fs6yi7Vfm0PZ5K7cOqx4SbVxngxsc9BMgPRNeV/ztYh0Sk/uom
blyAhJI9FlYr+BJ2AAowyIY23Fw/XNJWw2mI17IW2AhXyg5AvlBh7kGs5FJv
DGCU/RnUxBWRthhTLceVQMojbyrdQSvuOKFILVshighT4eBj8NhYURpyl16n
NyChKaDN8r5lmfnCrl/syr4vNE9zBe9X25hYMxpqDq5v9C27blgb2NIZqNrn
IbiSd2Cd86eR/WwN1nbUxKW4aZnJGDm16me9EeJWi5PNkimN2UzME33i+ccb
30YBapAnapNDKxeTpWb0bs9BbQljI6w0VqU0PDEE+2Q2LzZ4XKlMhU2LKJpL
A0sCCohzJ5C+dQDUMBS3wDzw69VDr/aDJOX+g2IUAEaYNB2eHFYHUazxdwsJ
ke+Ksol4BkeKtJGr0lVz2AXFiqMnW+RheCWClHsP8gdkWKKfgYgCV4cisbOo
St91dEoEEhFHqIInGcuxtC7MOJwAqoJpstRisehyURJYiLiiPBvMfvLS6G4P
BeYUcvF5l8jRIzN82r4PgY7IwoH6XY7lUbxtABPkj1wh6w3BiOqUN+y/K7P0
AsgSwX9Pe4RzkQKtmtkMA3qWSaAiEeLRA4NGtZJ/CdaHpaHrl+KdwkuEdyLB
HNrEqSjgkGvcB6dcbFlmAWSkeoLZjb6+DXw70NkZ17WjopKCtb0ioYGpxYmg
c8Rtq6kSMyw+O+LMfBem3pqQgwmyrgHUUZImLBPpkHHINno3V9FL3Za4z4ES
8BbbWoMfXT1I07B1zRHnaQszVlVw3P1riPOJ9Ks5T0Zd0QWMWbx/kpuctDix
/DH5eL1pU8948m5+xw65GMsqRqnB4VU6UfWxY35JgQvgf56ghksA/ICwv34T
mDg483oi+d5r4MHLeNPIQUl+mD8rsKn/UQTpt0Rnj1S03aUA3k9JwNDELUA1
2g7DF9b2U9jylEV7Zf6L7sSRhFI7g/RpTYjqejimq/MkVPEj4ftB3vfFIOh8
khX6KsD3s0WsoP0iGUEFUciV8S0MZp2Vo67+AxSA50AbUIRZrhqGy+nJDuPY
/FvrLKeu7ZmMaHSFUv3msy71Bf35uf7oDsa2X26vmGjVDuPL2xFy+LGn+SQ6
epT4NfiACskM9L7WJcT5LPjd2jj4rddNr/42G4nmR3e4u5lewhs8xblAJOHx
B1FJqOecfJT+0YT1V05PtfPd87nE5NFUDQvi6WaADSfQDcofqhj9PlgNhSOf
UbZHfQ4vD/uaAiK+ibUEN52qlaMsVAcROHNQcxTlvXLNej26VvJvWOc5e/Ar
i+DjRjpybMEApDcORE49U4NRbaeRYYSHD0M1LhBMnaTLbBKFdLnZPrcVey8H
8Myea4gxtSfHD2n6AKVgZzvFUR/DBui7f0ytXdFvUVb3w3oDfEGP40qmk0dz
Hw15NXCNkTD4h47zySBqaYPFz+YnKgvxWY4HJy9pNwkYm6y4D1m5DsucXCoD
QWwDBHQ4jcx26ushYl8X0qPfIF+fIOXGC3yVMXWFWQ89k88FraMmPrlo683W
J1BcYQW6N6JSeKhRDxz1H1T9AWnbjEIKbrHz1l8AiA56RyqnfYFL1qEJnCsk
juoamekOWynItdnl2S6VR4ezzVG+Gx+2qw98YFdtulXGfu0EJfwQNt53sI6h
2jIj8ugdK/XYbCncfLsTPAT1y78XJ558Tdbuh3MNyAaM0cW5WdDfO8ZpqoQa
RcDLrnkMfe8HDYwGHLkeidw+bGduaB2Hl982KOAmsXUJ0IMbCKVYPys4N2PB
ZmsmbNibtpvI9EUBldUyriB5Yc6ZVSNV7jIxxnBLrf/B9zsHtZyN0inpbYHF
I90e84Cf5GGfgNXE7GFh7lb6GX9p0fQJjL1QF3C7piHJO/5k5XzsEYRoQxEG
vV0LjklCgdavL5NhKwvxjte99ISueehh388KS6MIvxJCHKKNSi5dT0FnG6qt
WU37ZOGb4+/bLRfWgMiOm9soWSyinbaVA71ghsqSbgW3Rj6P4IeiFp346iOm
7crehgyO1ji/vaR1Tsel199VeiQ1d9cOFzruPXeumn07khC8PauNKr5x2RSo
sIyqqUB0I7EkONxBna5BydInEThPT6IB7oJTco1trga/xH8SVzGpoG6BCoTe
8aiDzHXMfxf71XnX/Um6bThaQNJU0xX0gtGvKGAqiDrcyDUpXP0RO4awS33r
yyJD8nVjHxzMyZVJZG0jfA+SCtCBLKk2dX9U1MYCervWO1bo+Efp5GJx1tz8
IN4/XNQHwdt1a/y+DbYvMDtB+WK3BPQX1UiO6FnBY9yh3vqZqtNpC2sLak7L
STooIIwKhMyoF64SuVtmkKQtc0K+Wg1RIhCfl2r8d8d18cpJFtLD7T3mGdQp
uMEWrZoW9l1OzA9tQfRa6rk8oX9jOup0dhcLZYWsVkm1onUXgtU/19COY3SJ
GteZVE34z9Ctgcl8Uk5uYOZFDC69OHTugR3daRl7YQQzq8Xp3XM9DFjAmGLT
PM9m4DbyB7JhYPpmohjR/DBTMBx0PFcR/f8sFC0bIyDMeTVSTcJcrbroTKCZ
utagMTfDvopDm5XA7/A+lLEWAvgp2uRO7jW0NQV56pKdBbg0grAtJvPsFoD7
rcEinu0QfAj2mKAeRhlEZdUUqd0GD+BsBLifvvImA+6uGTDVkZwiDbbiltZG
mRaQw0DRWTPtnwG8wMdpOq4xq7QfDr+itDzlEVTOS5pjN/bDaFbLtfzxYsf5
xg+SZ/HF6+gsyyjSwIBHO/1hAMkdxoHsz3GOetfiK9OQYPwMXqP5VeJNORLE
1g+7bf8wKmZgWR90AVaDaRu1u0ZLrxo+JLO9gktQrdJr2c925KCsQpw1MW5V
OqtPBqCAK+Q52OjM2Zs8ZQXK15LZ9++7KmmW4jGdtPPt2dqOiVqBpA9aFq4X
+hPJSYipOl3jq5NIgT9yYxQAIFZ1ayxHwfNESDrzK1AJbFygH2ZM1ucDHE8B
h/a7MlP6uz4n1lqrQeVSmvQ3TWK6YOiI4wG95/qB1xAMdBZ5hT4UHkx3HxSz
znLb2cw8IDa5JF8Obd54YwEYWcKeY+laMTIo1UrCwdc96KCjtDUz2w0+uQBl
mI0THZF41vBMVHdFT1hXb7rNv5JoYJbrH8Epmdozn0/inHesUlzJz846M+1q
BhCuMPuHb+bthCWiieZc4G/0Ui8zvSTN3eX7JpGK++IQywRTq//L7DUu1Ruj
np62u08EjkXywLhSK/hHNst/LkvZd42wxALRzcA5Esu9rtGbRx/R0Q0CQLQ8
73V4ZJhBEndbb28dG3E9l1Mq+whpaEMCJOJlJm8zwLwbdiDl4c1JQhcu4nKP
d8TAvNSKa3qi9Vwo4aWu5Hcf/ISulUi2YwYpMIAvTR7HDiMMNqBnVjLHJxDl
vFG9Kt0AXxDqF3Gi+1SgUuhZMZlgFu0dEVcbubMFwS0sm8yP4c05RJwO42tK
TUhPV/YlHAVfc80hQgDWlAkLT2nfiu5mLlZho4fOa1vo5J/8rmfigwxH0dEN
ayDRL1U22uUOS4NqJxXWSeNrzxssvGW5vdsKTWZZAcSFpRyx8wDgQTdD9Xob
Yjy2yKB17LOO1Z/jOXMkVY3cTLouKF1CQGOlYF73H411zkV1pyUpLTniGahA
kAeJwmDNzTx12ux2wtOo0dipcPnu4GVBromFa57J2GiF35I2cIr1y+x1lWtf
aY49OxYxf+V5F7anwXAyqg3HfGvOo6QW+SiG09/yALQsmxyfjnkvxaiF6koh
LHlz2zjNEIVIaNPakU/9Otx8SCjIdnW/O5NEs3jUq+WTfMn5OlFbqqRrPyh7
GkPGNAPKQM/RLM2rDRETWSTxHpORKpqMBHU/khqwmrDz0XuQusj/pWIANsmD
rfjPTUVMcbbkQlh6cqx7SzL2oDfk4Y5WGpnYORJFbrSRsJPDblt/siKrUsvJ
Dl+rPtjG5UfVn4ruN9EoXdF1h6o0l3jL+7dR1UxYqOf0J+LWi6ai0IBzOB0p
uflkIZj/OnzHe2XHnRwsWpyKpMs6eHEk2xWSBoxXKHCosYdlIg53h5I4NXld
QJV1cbu5jvanblzYYjA1PKNIukwByRicDFBluwhylhhCfwIV1rU0m+GQPkh0
Rhz/TPTTzWxWmfEfNonkvWtdepfIF5s/5gkmAVWQAykVplSh7e/b1gREkRPr
7FBMERrizz2bpYMxDAJJZVdkEDwisRxEgSW+iYoqQ1TY9Mx7C8efe/1kZ0Tw
p7PadJv5T8Ka3t+jbxLQ3qwtLNsRE+w9b6U6AMI90IUurTOpwBCnlekGUgEl
qzOPAPociu+mWVwmds2sQkChxaUpelojLOA2o5G7go82pplkIp8T1XM6RbLU
kEYBk07DfWFjBJ+7wTCchTPASENYqkznLHe9KgGfOERRGnj4NtAKAZB9beF5
JoBJTX3P0DsTQik/Kb08K2dTbEvPpww2E0XXTmhuU16AUIpKkZZueHamM8xD
wMas9GtIbonXydjbBvKUZsLXG3gUfX0NXUEmrU6VDj5i6sVMzXc1AnG+y9HB
g44kD6N81CoipzJYcTqVEhfuRlDR0jdhunDVJBGtQ0a7YF9drF8b7C7XvkVe
ZaYIsFOnLkBC8hxMLnPq/5Rm+48mRimbH+Lydn/NVL6YqdCcq+yNu/0wsbIr
3bbrCowyzgbrf6ldjtY8avii1+pZDS79eQsF8n12RRSWUO00FGrtRcvck9ge
2iECk5C9Gl0COci5Ctpu3Lq3TQPE+5oy02Geuc3hNuUSRSPgdQbX22yLDfiC
J8nEavcVq35PZ59KjJHsbAPyu1Db6rmaNPsEKb7rop151MXKrUzZq8Xmjsn/
YCjXgeCWip4s0gxAtbPwRCxrIzv/ZW+rfNLCnOe1T89xXSEmiybkgAK8av69
K5MQgvFqYdgYeI3yAmCyUFSJ2XKEEttuEufUIFmqF8MmjY995Iz3/5GKKEoC
mZy9YzyMc8U60wKaQWXDY07a3oW2eUXuceX897IqrrkvfAbNUsJooDwnQkDp
i9twYBz8HrVcO2r6sNG3kF/dJn+7YraOeJO9XTOAb0viJ7JXRgCoy1lrgrwn
TUNsr12FwhduJHrMQ5IKP0SwqkhV6mHascyhJKYoL9TogfudZqKg8A21X35e
3NZQFJauWg2stU38M1Zt8Bj0MkPDKYyYBbGboeyfXB7y2xBpSs5HEFma95NB
glkL1JJfLeUUY8PRPG27EShMkLFa7LyuqJj8cH22JJB49AWuTnBv8SyJpHsp
1NjN/BREDS0XoY6225F8tzeMxipbedL8eOt/6+0pH9lJ7+PuCDTIfqkJY8nH
P3/7FgEuGXnll5U+lpG+nLOg+wJ/hMO5YfaniD9EWjBSuaQ4XOjthnX87+On
1CALquZ3hUYJjQWuNZICd14RT+uzK10Va5XbMorQWznh9y3JrWCbqb2NVpF+
6UXb4deYkSuYrNoFdRAxof/5iCk1ju1EtuNGnM8yiL7je+Ask0+0j0SZX4w5
6ie9+5IgupkYFJqNXZyo1kizLDDHbTz2O5hKeoIUA5OfdJ6dWM8+d8bk9cuw
PMkeftMH1wu7xjItxakLBhOKKxhMPOXKk3pxeJcv9AAo63lUKx1fK/+hwJGI
zliFY5asW5pM1/7KCRWICXmCOnZQ4Er1XyMeXGptyAsf+nzRIHvTkSb2pHrj
K85xJ5NAMVuSn/XCdhAXVSclugVlHvE/Ms0AFdXmyHPeExDn0BFtt2GLdAQW
Rhk4KWn2ehQrncWcEsywn3X5oRD1jq5jGlDZ51n/7/mU9ssHjjiotbA+aZ3a
u7L5Me/Hk2fUa9d8hKmzbcRBcaIvDJgEvDJhwNwJAQwt/+u75SpNipBAJzuI
77+S1NxKDrCxp5a/avoXPzg5hSjOrzejiGvSky2DrCHgsCR506UOAqtNSpWg
UWZOYTyUDVPqA8OY3lWk5QaN9H0ilcVgJn2edboadL0vWXKW6O5HcEmDt7a7
BTErrcikYr73Qs2pDn/vfj+cUQZpdLlyKxQvaRhOuvoBBpdWd0AuyoFxh0ft
XYGi3pgQcFPgXpmMRkrAQ3Ox8kBeo2fqL6+dHAoW6gDt9MyKY4P/+CWyX+6f
Phphv8vw0Jb+3mCcKzMblNMQ2fo6gfoMx9QsKy8xLNJCTP6k8JJnQSthGmzF
IDMOKj6/2EMzPjziQBi/270Wsuqo13S8G2I1wtCzxuAo5DTj9CIuXOg5pJ61
088jE0XsBV6Bp9fAL65O2DMrWc4/+ww7slTs236kNuw/Gzlw4mB0gehS7R57
6t0InX/FBnKd1nly7Ehkyk0wzkDTPR7U+/P1lIdm77njtpw6frPMbTNjMoNv
0fdrHcgGunzip8+yFjMAgGWYR9i1SqZFL2m1VTL22iNQjQt5ez/17TEwZEUW
HZPpXLwk6zz06EY69OyRqhK22LvnMUdeJfeB6JYQTOQd92nplFW8X6c1Tq9b
K9ZYaqnuSnom0TFoDUU2SAlRlk468rzdgun1Ff+bqBIKln4SIzrTDah/wvUq
B94Y6w9tJPdXhKyap/1T9FjhBmQH7F7WAAaGDZFC9U/1CO81MmWr3/fX0o9g
nxTfchvc7yw7Kn0sd4oBHYpFlWxqsfGX7B0TuM03tsKwcPJ4G9tbm3lV4MsL
vNHMWUDmdD1GfNqIMhZgiY+9t1Bc10jQkkD207RSMaw4W8c0HFN94mJSgIcC
t+m7gjQj0BHMVU5nZVGvqhbr4esJ8M2vCoPuAxTmh1FIpaVZhP0gH0/PR5hG
4KT4wXhZxhaU1mWaLASovS9BGrIAZy0e5Zago1r0W3LwijAIC0btmEtOazP4
5nyx/3eHoYn9mjjNg+im9tp6LT7i7Zl7iFSfYbAW2MI2JzBpTxzoHixoLeab
qctWnGP7cnQ+bLbjXv4POe4ji7YZ5ZeEIqVZ8hCn8dNODImunaC6/lvcgYMZ
ts/Di8xvPQ3MH/YwSLIPHraMqwPxHnu5WJGsDxnKxVrvuHF79L7m+AZJjq3Y
2p+AMHt0Rq5lTKinDSBIMb3xVdKRxfMsdOg9QwvtL//VpyUmRqDEQDLHaQy4
D8S4HGZmEH1XpQGBOSA0LH7nzh3aM+kz2YL15rTCp+cCXNoN6YfNKXmVdlXz
z0Nm0DrRpGvGY1yj60BxCS9ywQtbXsgM1XukqhtcSm9KBSAE4mnG709M4Sc3
jYi7XGpOtK9SU25Ttt3ZYtzk1LaQPv27OOFDHWfP+hZtFpeUs4yeywT6By9S
RbY8KVelpR0kq9M7f72aj8j9GRbCDUiberkfROWOBb+5rfmPGi+TvPGcpkV1
Du6AuW6WPPixN5Xxdqolh3LdTqi30LMb6IAia+pqieBwcteuBuw4h0kFxQ7a
mO1QJeq5I6MheHSuKP8DCgmckN522vnYdOZhy1vVW2L/1p4YK3DH4JjjuMvz
OFd+0pwFpraaPhJZumOFXc9hyYlgAxT0nOspvYiDsmfxIwMcjhkwx0LozNl8
1Smuakzyo5p/zZfGk8wREnShtEjTvYhD4wfDUztyHhPHWEGZ6mMlXRwhldgs
E2mL4LQRL0TIjHNTHC8ycn2irPuMXneAAXhgg9SspU3mPXKAPaviJzbUHHug
lqZv27ehlI5h1xl5+bOBYZiKrN7NbyJlKF5cVLSv/5TH+rVO+BghkGsZB6Qo
hzygu/lN4Q6TX9f25Mvr53LYg4b3Fyz622JKZVKYW5mq0PDUOprsFXK+9S6U
Wninr8c+zvd9Ok9i8KeqZlNKQyPX0IjHuoDCWTKr/H5gghxBiRz8lRsEFVpU
K4jyBAeRqe+ufRr/PIT/FUbZ6y0MjGkbiB+NgmofuyR2ujOjxFPbptcMymj3
zFvE9EszS4JuWgcnyKyAwpxelJgkgi5+ps3ONtG9LvL/F3R5F4ETX5E3iVcY
4XVyU1Q/c3znkaABNuX3LAyI6cB68khFW+ESRI6TRDe6Hx1lb52NLntN7313
udw3HUg6ujcgBr/cWQ1WVThk5iXTv21AkIdHrfe7l/mWXJIkVqx3FAH9jM0A
aNdtHNK4VCXpwtBaXXy5XWO7L7B8yyC5PIHNJbVJ4Lx0pbmKIh2Yt5MiaN3m
HbuEjyyzYwdTPTzsebUYS48Cf6pFp+AOUNZCu0DHaOiy3M1U/OJxvxq5eECB
X1ts3JUctmy/O1YShTBDZLMgoRkPYKz87N+NGN2mVpI0lvlT2/Nb97GeuW9c
A+FtEDhyq8fWoU3qFmsAzHjGRkpPmf7VCsXVLxgSL1+5SrTOLnP2/vbmtfzO
iZxBnywq85NayEUDQAYXsIlFeatOePpZ/qB5g79C3jcwYTkzEy8duTG9E/Pf
eSn1R4VVb+YXWxuvfjkWHVJcIfvv2ONpTwH9lgpthBSRvDEMa8g5I5Qu2XuQ
/GHLn2QcuKXvScT6QpKiuZ96VS1eiXBzVP7dAwpfvboYMhl6u3Y3BHuIXN4d
9nuMQ9SDvDUtI4tCDqYevYByv/NcdN2Nuhced5YPRit5sZ1aWapc2HGTocV9
oUgWQR+U1OAImkLu0D6aX1B/W+C95L2gULPB8juRxjZ/Szfl1VxF/IkZlF2C
ckHd2wYN35lDg+bdq7eX/zH9cB+GabpgdiBSgPZBdjXIAlL7URGkO6TD78bp
MtnlUA/8Pc1lvJypllSJ6WgXgg9Q0fBySawGEDkjUPml5jr0j7rHZMu0caqx
6n457pM9RWYVAE4Iu2YPLBchWgw9y6IlFzmJvu7WMQUrrzKa1WAifoEF6Pra
ntRfZgVveVmrpOePlYa4xMoNFlnt8W64WjkCTkHGPFrJlV3RE465x99J/3Hh
id56SjPYEkbKjRlnj+PvtW8zUUmSAJ4/LZRBm1ZJCRGRfG5yj9dNwpjyECvc
7jXilXxEvXDShy5exJB6WW+5EfdLzRSBDpQcOdc4R20PBoRLBMxsRtJPxpJN
dZt8XlZNsaFcpFV/LP55HGF0f8bOG5ibSynyGy8qXWTZqqwCc18YHqDn/Nok
jCqI1nhBayUs1txVD2ajQNbXa1ONmO516FsuIZ2HQF6/kmoxT8MwoZ031Ezy
RtZljeV6z5r6JV6O9VFSrWmtT5Qt4r+u5nqUFL9pdGy2Etii4T5czOHcE6CF
RkYGEMhkFjEyCOVadhnKcbN62Frt/++dppO5ycUm7fHChVPE/i86my0bn7d3
rVyUTq8U4Tgx9nyDvQUfuU9Ixe2+siilgu49BL/UwjbhmPie0vfygO7r02KS
l5p0uO9DIHaJWBLtIQkaqyKmZm1XpqnCnwL6kZuULbYecHvnlx1kv45h06MH
dr1BJy6m2ug58BW0LXwchvTNzi+Sbw6a2c+JuCycrA8Aj583bDnN1L00SWt+
SMWeBt0RFAG9TEj5XjXl39B2g4sEzrkfdI2jqCwpz9OxkM8S79Gr9fYIo2eY
Op4Mos0p7kASWh3Zfk1L9gIESLegwuchL1U6/M7k1l1I+r8C5PjkFK/i5RYw
5WlCUZYiLswi9OcY/GeVy+XfY7Memu49naC6RmTj5ink/kg7rdbyaISylwHr
FBPqBoKTCpflXJ3XAIjxmjYEwPTDPf4DqV/3+1ScFWiIs9Ns/L4UZ+r058X2
7knTphDSTngaph/aLwjS25A+2uMD+xA54H0wW+CjcTLaAC6ABG9NxI8cTnjE
7lwcNUCk1uqyKQaJH5HG4RQSYiJ/wAmXvUSmJ7fRPlU42WrmdndGtXl0Ka8g
EZ8V3xd/mP4W3j2lt91zzLdIBSS0hLQSNhHWiM122XqSORu/6WR6zhnrKfuT
vMGCDPYUxOxH+Lu83I0tLkyFT44au11jgW6pnfa0Vi4UCHHOYHq2K661yL0m
Rq3yIv7db8PrjeuuVfqX6F67y0gZPeI4gsrQueKrwToXa9NPs9F5IlZraqBf
rFoIxDFOTxtttq3bloDbAZHKl55BPvfX86Grr4YWvD8xPcz61X4uc2ytv5mc
ZQaaBosGywJSKW0CJ5HYGqOcx8KF28Cf9mA0irO4Xv400k51C1SOQIoaObCZ
OvcmPjkMWd9DIciap1mfMcOSdkt1qhteNApjvjkE/LcSwtJc63xPC3h3zl6M
lAhLDyIviDWW4nJT2Ro/n/cYduOJM1RUGYdnCopiGamo6ENOHYTWxEbaf0Ag
qoBAtkDvz5Z3O2+Iad04+VUc799qSB8X4EDYBlP6zJC1nxdDfUMjcska9Eu8
K4DmJoUQH5gakvb4vzDbdPzJk51KsjgP69UCTxGl6tqJtZHDMWMF7Zie3r+C
oEv4BxgIVofWjoOKdUC/3u8xFspfi1zbtBtClqJ+14b4nDRTI0ELzaGVVY9G
YKUh0vDnSky0CF8/lXUTHoCVV7X3wc9MA53HTt51CmnoHHcGsV75EveELuuv
rkkL0LAJ5572IAwaRR23++vdpMmIVFbRoMdB9Y4UBjcANDJyRJ4RHkVPpQ2G
X0UthiLKHE53iheT8jDO/AodKv3oy02AeOrLHynkaPAEN1PLODXyjqDcOCf9
yvIreePNKbHduU251PBQJN1xBD2gpVBoc6YT4p/M38ex7jktMza44y1apDmU
CjxWA33FJJgIEUSHwMK6kb8TOwx7rCZkT5oFbuJOhiOLCpsHeDMCtWvQZlZu
HNwatiagDskgFA3MijyVkw+l1YxK4DFHU1rX7ttQa7dF+L1bcrvr+NzaAk7I
kYXAsRWMq51xnbyRxxpDTEpCmUfHm/cInZdeKocgi2jcBdNRfIA4FMGsjjCI
e8KV0qTRWwvurCsbDclCvk7o88ABNAG6CMa/E5rHlvYtXZ2Ko6Ql9tOuuf8J
Ax+Q84j2Yxbc3K0ao1igJFmXA9XhSGhxeP8bY2JQDg1G0Zhi0je3ZUz6MXrZ
GSv+119expnRsZYaTPfj2EGJO8VYncCjfTYHHVCJO0AlFdusW3pMAZPTQ0Hg
ZdP3dEJqpaGf55aQsAHxt1qd+/ZXd7MqtuB53+1bDoFvK62awo9H13oXiqqF
Qe0RLKFpp8jMSG2rXLkStpH/PVCfMH9QrlMj0qnL4aVGJysi7a6mo4bRKPz9
6NMMscMIwqf2wucX3F52KsQVmeTDEFlzFXuE8hD3PX7SbyFAH7f6DLFJI2Z+
2nQMm0TT0MlzvgIxm12P91REWH+7Iz1pPL5V0V8qNK4uNU08UmigaE5B7hko
05trfOJL015RldtAkVqgcxJ7p2oFiol6CI9zyjvEm6XggvpWqWs/hwrv9xds
X2tt3/k69sicfehnIGfhEaJhcO74dwfbsHaaWjl7FGynanZ0VckzeNcL/4Vt
oD9pGGQXOYTXn0I/zJOhENXpTeu4WEne6eWwjj+hSgFOPBywcfNSuVpSfs9B
XE9rIw96OVVXDwTDwWl2y9Bkh7jSwAIYcSX70H0NArwsCVzwKu4tpWc0ql4N
45PHEHytmU/EN0Oa+heyF7zb2T3hy0yExisyqqNfVnRb6eGtc6bITvmHHeWO
V40UHfy5g+cqcZGvuxqQE5POELS4mVUqwo6xAX85U1P3NgOVqL5Bf/n2sxE6
xt8wOFfc2YvjgJnH3aB13ZL144h55vx7l/yHh3XqR7Hnuv1yKqh/4/yNcWWL
A/QnfMbop7K3IgV8EhKq2LzlwjUOlv785Svvc3tJoYLPJLQo+oB1jmRqDu3b
FNjEdSf2rTg2ju6Dw9JfnCSsePfir5gmLzkWPUMhpTC80lE8InzLhg38PxQa
x7ZRUphpT0kL8AK5/1hNSBC/uU6WAqBHygR9Yy3fvVM1HpY7iWfpHCbkZb6c
yhn4d1s2qZfawwZINk6lAPqnjxlJD2ot5vqUxGYX6q9I3Kj5yH+eG90W8UFn
H4V5m5TGIpyTCXGuXJeHA8zhNX1VAXYs5LnJ/x4h4U+d72YBhOFIe38kpIrj
VPsj9DjnZQp1vCswBLayN/DPCAmmoH5lvFEpVzxOA0zWjpx0i1Fv0LvZa2n/
z0Ne3cr7k1Q3bvTLRoJQTU8Ye2TTbqqAvAdxZfAgfS+uXyppPa3fFqKJ0+xD
qSf6m326G4n7KFKLUND9aHfeuyBzA+kv1o4s3/kS9HP2DPiP+3LPLWYNHCE2
2KCjtNEU1FoIyj+xhfMArWdGZB16kpVizgaLJ5KZvELWigt3Ru6w2vLAtsNZ
Y7nZBgzXHgvVQVEo8o0VfQeYZTRYahfddbUnYSKKKZ1GMVZI6pywKFd/PqzZ
myiWVH+/D/BhyvYl5dBuQ7TX3hYCA+Q1fTNL4BnAMbjucJkJryphp3McHD8m
kYwEEhIiuf/5nUb7bA9eWfQCjGUAVK2a3gugiEd9EPW36eqEyn4i/NgjiuIy
wPtPJ/CN10fntTRMOBWwAUzrI5eQZlr4p+pj2Brt2P8YHi2wNyIiQsrCrrEU
V2pGWjNNwk3QHq4M4TaIJnBwTij0IoJ+Ml6ke1e2OceVWl1ry0INN6GtZiIH
UBly6rn0Hlt00uHEPlggA26xdzDNTtnOh+26qOClnAKH4rnlJLKA2uM4eM3H
8VnCZ63zK7bQbCJD6cGc8+Sn6Y6Q3SBvps014luM6GBEMdAVkeTmTBEVFvD5
Fr3oDpeEaLczImLo6VA060NVRRErK6gUS+if5wL4QbKbMa2bdYQBDx2XfSNC
THX5zpKPxEpkgCo7cGwuji6tBSsC+1W6mGlDu64Jx71EXyybyAJcR8D6+sja
NHYCkA27Gb+RizkpEYUEVgwHI/rh/QFDWNoN2k8h5qucglo8Fck3CyTgLQ27
eynSpvE84wn9FyHpmeAqWBAgymdbDC2WGiaGrotlljUR/fb8tF3KCMeXQrmz
vsiaQPjMMXKtQ42SAHsT0H001ptbqWPOaWULr5Ag6oELxqjDW7ssOMjxCxjK
f9QC8RFzXJmkmngxL3Ze5/5LLiJIpBVNPxlgS+4N1jVdUYVFhjpeR7y/hLoZ
fcmz+K9ply1Vr2jl3hb1A1gAKANW18as4bkN5OiR2Np5L3pwPKn4gA8AXRpN
eP/8Qhxn1vCnTNapGVkq2bNMJcXfmFA+9Dhn24OaZho1picfyxThFfUtQbsD
3BwzfUBfgjbLSiSRPr+tmXiM5tLTTV4EDJNfLeyyQdGVyi8cPrMPYDVmARjU
f3ONcF+NYuApvJWBYrUbz7d6ZqfVUI8oTlC+wpPlD79j9nffbyATngV1af4h
1far+12rKLQ0VOGIylKMaGfk4oZUS3v7BuHn63ofW8YQWkbdT9sP/kBJNTPo
3ovYvDwqxFg/D7RPxK0qlHlSBZZBlxlILMfDvE1m5c8ANjVJMGxzJX3TZtJK
l6Fvr/yt2RRn0do6iaGToW7BWk+39MPCFG3eINys39jcCw7yQuF4irBeMAba
pmfmhbpxtof9UMTGE0KXPQJ7eoFRfv4B9AO8ck/exm+n4mkCBgG9qlFLb0/4
Qmh2KwTw1x/u7Kj5zHOYtExMj9FRxie3i4IJCjKmI6xVAACHYT7GI+R0tEdc
G8QN8bEXA1lIsXftYo/6l/80sjKIgc7fM4OypD4dmyCYQhU4llXsl2IrpvWs
1Ccvv8AexpTOakrtI4TYqcZOrW171VMwNpM0fFIrYhfSiAIBHYQCayTgDmiF
TOHLlm7iF5Q7kpiz9paAbH4LWH6/ORwPGxq1pyVNFZ9iQh0g8/7ZcXIywwpA
yw1/5LY09ELU3OiUvO992+073cBwvFZQ/PIV9+H5JNj0hVMhjp/9utTvcVAY
gL4VgNp0GTMQS/Q5qjy79ktcELdeZkyeGxePD2XGWft7MyZttuGjUw8wXkgS
S9IoJpU/f71fEcFVyKyJ4rJ95p/Fqvzy2VDfiimO0o/8Zpaapan0AfVTWGqQ
aHWLB73eLNbjvFq2hYz99a2V0nb1slokenBKXc1QQ10Pt5G7TpHoIz5jLpsI
VyFYf6VkVkGT99wbqWNMxgGwrytXRZYGC6gDbCIme+2V5dQYz63/dDBIMhCi
+cZxLw7zj/YO1DXrp2rYrCc5CfAQJeSgILhA8Tk+9F+VItA2z3Q2SznDq6On
8ZkgSo+lfXTkcLQB+QFx7jY3OBxa2u0I57wx5nItjAE9N+6NxATUMjGbVSHp
2tfZiVt0MPnXuNv8gbT3LtS59glGJuq4tvJWVIEXDh2Cw7K2ycQ3gup1Otew
cuhQIHy0pWmQjrhaA3RNyCv++nYJ1VAyNb+ypD47XqzZGa+gqUz9uwZlVlrC
Oc+GpNQ2UgqurNLEY/oSx1W1JZNqu5FXeCQgNzl9hs7IsYSiUW/GUTVzqIko
4tW5dQeF9zEz6m+WnNV3mNBwaAq7kkxVoUztvYyjrWYaxYkJ9kAd3voR1Cuo
LagnBeMfCFR7QZE7ogUoCuDQH8nv/r2KJ3zuCU2daDOveCJ6lbRUGVSx4vm0
uZteKKTy5XdzohBOyYUSacSB3GQay2QR9mJvH/I2x30lfWX7Bj0C6YZPOUOl
IP6J/bcpqCObl5HzYnrDMjkCX1A3qKcqWnlP6ddM+qSnieqk19NKZRh9k9eB
dKIX0RdaupmIahBvH1QrZ2WE3No1iyIoVqxPTdPvsxMvXieRSQPV17YWbgU+
IMZahS+ub5JS8TYRbhS27bJ/J85I/HL88pXXZx4LNkAlMqTbbe7WjfwHOfP1
pUl/sFBn8eIcscJqOlM4bwPAv89ZWvp2I/gVsJy8x3LpFo67ZGVMcZljrCQE
abXI7XRR/zDTOGavupqtnKYAL6QJp09dzuuoRhiYx65V8waXQOr/SqH8KYPh
j6BqxThVQS/9ZAa6lWBdRQmTVKs1lyuLlxT5ZFMSYQJZNPI9n4BvTL++Vv0k
Ai4hI3XtkBp+vv5unmMZH6eXk4I97t7bK4xHJznZXr6JKzejvPEcRsQAoIQx
jdwzM42uhMZ6USVxLPryZtb31EqwvhSJy/Q0v/fuXxY2NUgfoothCoYIsthf
yT5eZ1pWjJUn1ub6wfdNWzF4aBOfzuA5mayY2qQEgOru0kgIgsDp/b/5aOwH
2AM5XFRVljQ3zbp0xqBUBSVvqTUs9/bfIWR9thCNB8yh1bZG2AFunhd6nvTu
0w9bpdGOmw8VBaG407sMZJbcGrMWWfOZ0c9DQoFAglXEeM+xPtfO0pihuZfd
Yx+tX40aq16EJ9tcA0mA5r2xJOG3umALZziEInGn2uvZNu+sKqJkz/Jaxm1r
g9aBYNYBVV3IsMSjStko8WzRhuETIsjii/YYP2dAUqMEx1iFJbMgRAMDSSfO
ryPSu3WBqMReLg4R

`pragma protect end_protected
