// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
hFzZVNRjBw/zcvIkYia64a1mRzBACqz9I6r+M1T/pzphhGw2T/doKcPicIAmzaiJ
c/de2QjadiD8JuePImOiI9ncTp6tRgNXKA8v9YHCdfPE4gh1Gg8SOP+aINRvdTKy
UajhKLOiaJBxCQQSQIGGSFIuDt2OrLh2Wka6Kx8VSLSqkSVuZoFSUQ==
//pragma protect end_key_block
//pragma protect digest_block
swb6XR5W3ExMEkjJdI1E/82YEYQ=
//pragma protect end_digest_block
//pragma protect data_block
rJi9F5AiXG5Mvi4TZULlvmgmFQp7DQmslPQeW9Wb4EtqITwSMNVdnnJb6dPgumbM
SqXilu48ThGjABWk/GDxYghxdPkCqBbP8cxiEdcntASl3LDo2QiKoAlVkIwBLGMz
oXMi576cppqLXy6ih5+895FFwsF7G8+aCJW5Jx8gPmwVvX8c5ZrzaO1RwgEKbMSD
HZo9aN97ByNroxI35eFuRlYFc0RYRVgzfueW+wln39oEdmw/uRV6Bf1/J+1jXnF+
XGoyp0wMx0TV+xNjZr1ZwKD12bBRtM/Pa7GvEBI3UDQGAuB7KzP67hZ77NaGZgrd
UY/owS887+cA54gjGPjHyl59g7nalUNLAYF9oeWdeb/j9JmLXPHQGkocJOrVp+p3
uP2jdYTonOa8koKZ5K5/ZCXgdIFtWVi2KreekqANqqhbLU9Iuwea9zCveZe1+MCC
lSEKegYNSkN/Ws79xtUyZxQBOpSIL2o7yxuTWXMNdtBGEkOJCVCOZRTmsFo+xgoA
WDp9ZLpR+llq9KM5wqWG0QtVkpD8O95rv8zcgnRNXC/BeOnNrjewTbb94m6HQTCr
BTT6Cl1R9pEsKhG/Stq6q6s8/vd+Rz7hjHyQMI9Ols1cTu21Y7M7m5t9rZefdX1c
/qqTZcxIMAdM7lnnzS9Wr5w9ZxAAGB9+jVg63F4fs025G5Lc/uALiElQWLtaERwr
JNkr/412WRV2aoSf6jxjgqp29Z4KPFhPRTsxg6rW7VazMIS+95J2EcyG9cyu+YsM
mU8sNnVZJ6cCSnq80aKiLc5krmjUSWWnzhRRhQ/swC+SgXmEthca63alOHg8Yd0P
9AyxYvYY1qsgr3BDAvpqykS6/og0iaNfghnBEFSHrbhfxea3NZsVQjLvdBkpfiGm
MXNxQHt4FUzRSYBbSJ4sFOQPYMYsYWRGFafx0DIMCZu7w7zsrlCasSc9hdFJC4pO
bDDBsZoBZIBxn0cueLuyz5T2cihkcY0ifyNYWbC8PzZc2pkl8Dt/0mPOMJ2moljq
laDTT4XYDph1Vrl+AArcX+OugSTBU2KdoXklTdun6hPF+cGEnZNv9jA76pJnOv3R
n462zlXhBV6s9J2F9c5N3VeCnv93Z1N0LwtgALWNWSBQ1fFemA8lk/0yxdzM57rO
euYQ76KivFD9gKO8UFpDS1oq2SbXo9mRjagGtA6YGXehQ66VambXewGj51MTftHa
BV9WuWowzd8wNrt14fGd+I7Xe0rBo2m3wXRokHzgGBABjQJ9bY79ogmUbDvb+/vR
TzCxbrzmdm/Sfl+CQ2pyd4n+mR9Rk7IMhuvwLYzBWyIMVeERgq9ReWOITjOS5q6l
6M8wfxlOnX4W86wDj75TJ5zXbrztXJa+vaaOc3HaqDreD7zVvBDnjHnAPtQ9R3Zg
1pb+JOMSYmL84k7Ge67FcdWyk/ht8dX7zdcJtSgUiaqToyN0RyCNSsv5/0/vteoQ
OePudAbJRg0nC1El86DNbZb9a/5TLLkVrrFX27j+F4yDkNZIiHJ8tq6J8XaFN6fi
dsxMeRJ5tByzQJ9GZiM7i0p0z7OBFgqKaWMYqnun1+Upj7bnij64ivRBQiEzD+HF
+9XIx+QMSZcfl+OLHZehXB3DjWTby7mK52Wy7VxpScEiv7qjThvjKfhw7eiMiaYy
uHLmSR2dctd/NL4xlGbEOUYTqaT8R/fYZphJK+dOaQoR9MguC/b9zev1JyguigAv
ZHc6e8hezbZIdmnDRterLlS+Medb3w5Bg1Tpcu+u92D46y8Nk32rURPZ7idxDIU3
HANyYOun39qaF8aElsJQsHOPZ19J/NuabMz1+IcGmvijnZzpFdTqXbERZth4qnLh
vjCZD7jQzr3CHSCmrj4Cqt+QAcSIK2pqE1ZpgFXFT3BApQxkO/r3WopSi6nQDYI6
NNMZx3YfomTpZcyhei/bKyAQlyiT678pJt/88YXcrize45HTjIUeeelPWxiaS8Zt
G5lShzIEh8RbmnzlN2bVvGxUxaKNCFCtnVn0etd+W97Z+lqb4tGB54OSxntL+ybI
RZarW5OK0KioIqGfAQXywz6coUEP1wZbouWqjg3Opp1uikNJn7b+4C8oxujhevuc
yXVhdnSnaXn4623c5iZLh9QCOliHMLspl3YqvtuZhtAE3IqUDQrZruYkbRzSBwpi
f+fWTYWS7wj/LLpcF6JIH8rbOOTpk69Xq/XnfnZEq4eyBGnupN+0lgavhuJ3rvDm
nGq40OzbRy+2KbSopPHVlqGxVXa6oK5xcBKP+6C5BtutDtRHp2UKy1sckRkxtkx/
jxvvxLY8Bzodi3OySnFvgimlVm2PAFQwF1rYLKs+rv/CsysfbIydpkWtmnop9QRj
m0E8Nqzmz52DvZNOS6pimkBxirOUrBNsVb+AoJ60ONYUWWeBcrluhxmxebPPwHBl
ZJfp/bFJssRkJx1DFgF6vh3/5AMRrRM5ODAaukB3onQ8707P+xDRW++69iy8uV2+
YnHM3MSjlafNI52xTWO1YJWY0Kp8r6LHEPMhRlnL70i6qQMG8gdc8F5H0bP1zD+m
WndK4euWPe2Fb+ETAfWAh7x4/IhByZBO8InAW+X11nU9YIkRw6UQ0Dr9KWykm0wx
Pov/eGPZ4E8iM386YWoXFcRLQoRJj2qdMSDsnYz3Xa5Nu4b/n8c1xoYG6WSNfQyo
JiZ0IPvXzSgTxl0M9V/8bPisaC8LClCAUyNoqr3F8ONKZoVwZE8Pe8rUg+58S6Sj
truRKtNr3XJcHzIRh9CEMA5NA7om8hQsfcVXO6gfxlgLOF5B1TDZkamQcERlmIxo
/GMhVETgV5gEvVZN5RWcOfObsr2StFp6g8wMq3w+NLtT986OcGrdrh7L0iGvLWEv
ANRrngJQD4yMgU31zk2yZ/1byBB77BVt9MW0WwFAAlO2N5pY9P3aO7NBOqpb2g+5
lOfzU2d94f6U4ggGNqOdi2iBny20HpvDJT0cmjmM0JHW5vRb/CnogfcGLPq/Ocr4
MpXfri+/mBstglnWzCkkdc3iJ0I3Xk+aA3eQ8LzFBy9W4tvfvGJrPr95meRoi1Tg
hsJar1Xi4VnCPDHmkD92f6XF2eOKpxMkaCSrM38RuHrdWwua4ukK60xG5eLhKWkW
Gk576Vn/r60tPPbGP5ayuAmUz2nKB/F1kwieAwdTjcpaqoEeHBEmCtqxNzf6NUqD
pMvqs43IgDpFO8Ie8U1orEfcMOgyPjSzSmj94bh5EFvH0ZJ028fyQf056/2JyWVG
vKllxp6rW9rAQMzZa+4xxUtQaOGzIl4lbRH/n2QMUQ4Qq+WW6/Rs5WyL/7ZzA4YB
9NJxzhZAFzwPuwdtWMSOBY/k1VGgVq+vai0mtS8KuybAhab4+JwI66yZtPKHL45S
yelfV4BY64cHt78LSLHDJHB51xAmYDm5drXDHBgFgabms7hrWlG4bE5PWBx9p36M
qs/MT+z592f0UTL99DhjALRlEXRZdCmLDyN2UYiOSwEOUSwi42yPHPRfgtJVpmI4
B+xtOdIpypJ6bOodnBJ0WeR3mTZCX5hNRLNjcTyFWTTkqSjM4EupqK2hMII4UTy4
qxGK5cWi/p3Yt3JvdcX1cfL9Vq6i9Foc2Lf7jqhMOPGc0t0jCcjefXqJuZWSZGjy
l10HfA+Pif/aZUax6A5aK/7zjMF5MuzuW9AAB8xXrRxNmCB307hfdr5S+tA4j0cH
5asUPkSAOeCvj4V0ZgjVGVv+EJoY0gM9HLzT1mNqB2Zs4BUdzVdp2a2zUZ6qYitq
vHoJloj3hnfAwlPtbderGQVhd8mucQzhsXs6xFd7GY8NwI1Qeqhm7SvhVY7DRxsm
S0jn/5KTFR1PUDVuTkc08k8TEnDPRjUfg584I1QofPWFxjapFH8ubQVBTLHWSX2S
j+sWmxcpzchdg/3d2Rn0vzDo0iP4v/iDQjnSBEb4MfmvfLInniGoCG7LgssOe7MX
gF42skPYlcPUE8136sckJWb0Lbl59+2aOQQ8WpLr+znOjsrmg3wvOeI/B9ifNmML
bqz+hyJwpOCalDk42ezpLE1OA2OYyqkR5y/Lqd6eeSvijp0yyC+Lv7VHUObUt2l3
79fnI0DgDc1lCdtXDIOJ3k0iGxby5AypOQbJXRMcLiZ+H6Y+mIohJJeokrTD0t8P
6maZVQnrZQX+WcOUurbTFIZDRNyBz4KUM42vUt/m1Jlfs4tyctkwXPmMBIa7lbiC
7n1mHEVKlgsHkYwe9mKOX81qgQdh2jty7A0JM7D8kCdck+GkE0LSPDWVdQCheyCg
8SEtsitAmKiPvWQrTASZu5c1YiBYY9lh2vNErkV5dmzguIuvYvmp0KfVa5gBigW3
pKHiGpyr4u0QiTJBoXAbl3y7BQRstIg2AKBkolocPzwEiRpHBrkVT8C1O/BMKApf
e9DAEd2gHdIX9HYbw1TynmKWtwv9jStbpeuAW+nIjSpPZop/Ujm4Q1VzTVsBTGJS
G6+wErbPv0iOA9AZTS1PhJLU9n9UrOdLI8XCC/UflknRkXi7owDrqbN94ngog5pl
Dc6Cf6Bl/VFEdDUn95MD7NTYwA+c6n7Z2xjDgjD75xG4HtjPK8GmPYhjdF/cP1Ua
zEqPLYcBzKj6oS38X0b28zA0nL6SDNPsa7jgMgk1zr9q18AjE6xRcnmciHKZux1l
qhLzUo0hShwhwaeHd6UJG6vjUy5IGGiKWVYc3ng+nJ5HASR5UMwCVoCmuezECcty
JTkqebr6Du5T83JMV1u4bDl3z8M6Mj6kl+I8HsZikdU61UirA0bvxqz2EbZ3cUMm
EG2v+EfRs0vDidkwvPCZ1ap9O3Ztmwcn2tNBG7rEBqhQu+u7mAiS19KPtGnXeFNR
9R7uYqPvKTU6XSQH9Q4yKgft8hiv0GSg4qoecmd6kFUUnVC/G0pnFvIEPjwej7C4
dxIxIdXISmc00XCQKh69Gz395GxsDckMIPmNUmwe6ZUKYGqsCvn1c3TKILR6oI76
U9VxNNUS/QXFgCAu9G2AYzzRVeuSfMoqJ2iqQNCCaJHUKMRdHEr5/wRbJPV5ljZD
jB4U45n8SphDOpwLUw9T0DVGlElSc12S7ykbCxEhxfBIf/j/DaGCbVyFZ1WzILyn
SElGnxcvfPDTF5hziCxvSUpN1ne0EjXw2UyvmkksuZar33XaYrR9hS4dpZQ2J84B
B3+3cdjiW8eRCjePavST22/iuY7HDTM5XWcFBQs3QGVb3qPtcsRb9MTdnT772U9t
GOnniTRy51HgIgsIAx36jRNwlHSpGzCpGNq9M5CzpCR7Fs1VFVrfmtjoKEO2iKMi
gAiL4SVOkV6oETO8aeSXfI/ZCIkL3e53JtdhOWwGz9RkbtUdUx8hkCq439coyxqy
tSfdiOYIH9fLUZBf684PBtx93vSWBZclZApbr6oCpyQ1aOSjzUjFpHTiQ5eAr7Us
b5TTIXfHRMDli5fjcscHkQN4ZwMeeYeuEXxXWQOrL8cjz0hc2I7n707P0QnqAFCY
R4VJ5OlLhfhHZ081iBrtEl0beQseGhUgzTdXo02mhU733Lpnz5tWMpQqOWzR1sft
4/rktR8ZmlzrqWBK9xzBlYDmHt0ogzYXXnCVmNakw/BK2n9ARcY8ziIzntv28+HZ
t1YtGm6DkoBTdPgiZfsL3UG8mn9j+lkjmp+O0W3Z3zOYRFV4wFn594DK1r2fSA2j
cBZ6e7wzm+zGtreAqgDZ2xLSsbur66LVd9LMw4La6J2ZXG2UbZfy/Sh9IYI+vjhN
plOE80yI/oZ+V+QL7mwVxZFfMnPBtFNXwTxI+0LCe/kg7KA0iq80occqztvGGM5E
KzrhnDx6geb7Ib+g/FmOwolebMfvmkLlAF106PvfCehNsSR/6Z7Og1FUiXgCLcq/
1BxjU859fRTnnzOwPCGIWsitntrPcV2+X0cXEJZFGGmfV68yRTt2WW4NM8usktCd
O4e3bXDoWVA6Kw4oLWHYBcr8LFp8X3hSXhliOZsXs3eWDLWsWpmae3nbgqX5Nw7x
YYtcmY14L9ljwTPcWmvkoNOded6cJkbtbw+Y5eeMWpSD6WnO5Ym8nWpnCjaAxXtQ
qdjWR83Of3YcbZ0vgEJm6fbnrlePaqp4rcQjzJxRAU8USbdEk4az0rcIX48JerTA
sMypWU60Hc8RmhlH4NeA5OaN0sDikRDIhrw/B3Ci9HeYNq551oFrOGfNwXRekWIn
zGNwcw4pQ49g7aSQkcfuzJqq6jl9h+kO66blLAiiWFQKovmyxXmyr4HSVw72gUJX
o9kkQkjBcEEzFuW1sHadXqBMMSYxMwDeZBFvnsAkgYhwEjIIyiIaSjwYsN9fDUax
sm0d/yWYlDrEtnBsZi2T27T8U2nHxlGdYbNZFciLNmVSjDsP9IBCyEPNNdjq1zpc
TBz0c4ORt7elZxhpQXlGSBhpWZ0+cF/Z3Czi5Bup2TLIELyzy3o1h+11PYWx/Rbv
lFS1NZKRLJzD4bRi8RNYBr/rwZYnD17diojMxSWsmlMBu9lsyriBVmMCfYUKsvTt
rkKv5UFWfA+h1SOKl14z4yOs/bMUqrC5IEbfL7IAJFtH9Am/WxgyPKxbBlaMvsyt
X2Aw4Kk8zuFcpCI3oK/8jo5FhLMXHXK+BckVi5mkAwv/eViQyAhe89MCRHMgZFbZ
Vl8FbQk3ejG+GJt/t9yc5UZSQPljdZhvshfVcUhZS3UhIsx/whe7JPCL+rk95e65
Vrz7PlgTR8NEAVTNWh8shA3E3p3XLKnJ5oXGMUvlgXBBFbQpXma9HNOHwXWkXNXX
3E35LQ9Wi026PaKGiSvX6IvGQZG+77k2GiLJWGau5W82CbjTzyqn3Ers5YjYBKEt
a8Zwy6S4SJl29lVb9E2WTdvYmcmPD8PyU7JSPnKEBSXGc/PJU7EuXxryS9t2Dd0P
/GNifTxFgyI4ZF0bCGK8Tfh50o8t5eOx2x1yB7YIVvaLplfb1efAmlWHts1abx5j
gf34fcDx7emJ22CwzmbF3Dd54ljamGNTODdV7Tss064bROrzZLusHwvorT7oSKa8
3/zRHcPzrHBjjWZCWppoduNzbOJqVNYYXOzNYWlBXqbr2m/82Q4nD4F1SxPWKbJ7
DkSnVcxXil2H1l8uC+VhLHOBC8Sl6EjZxKkt+4tGavtMuyWlbzusY5T5t/MgwXCh
4P1GvU/2W1tLGOsKMjjpLEOl0+7zugtj2NwLofsdHUC8k3Dsec9UKVa9ZdjJHdT8
gFdD/OCftCLuih6cL9ODI0pJcNleZyWNQRWr90EPoOtu4bOgjxZnE4oEVzQDDrDD
2dAnwROuVXPYQpjyi58xOqryTcjz8WrFxET4kzs3xfqF7nFN05bfuwk/uB83XUwJ
OEtYiEORLJ/+ob738jirP4gVWc4bHaZqQ3mfxxVlhAqVEK/MQyIsp3DAye/vQOXe
EPV8zfy6B+DtnCK0ErRqxjhDYS/Un+DGUbLNWDY5VxdurZiPw2uMzjnsHOv1tMyq
6s9O8hMwFoj3BigNWOiADupNz08PAxTnbLBbOrcTIMAvG4Arv6ltHOvZVrHdvRbx
5L0Jb1JGrQzyOtDqKUq9O+NSizwasKbqYT/dVBTYYObj7p+u89N+qu2nbDcaWMNm
zcnfZVIw1pjijZ/JzlcFnGy1Eg59Wl2AeKRwBDHXrU807PDQHt9qGETovbmxcw/0
X09IgQVu0ICC+BT3Ukb1jASPBOf8yRfVvgLUWe013YhWwVQp4gnkJebulWJzixj0
MeKZNv/y6lY6ekCydvKLAaJWkiWZ+is/bevgaW9O//gpvYX+8CQmh/mTS/ZA026q
C6MIPTG6JAfsdEx7OIvwhQMQDlwJ0MiHlXH/+sFnjv/MqsiXc8GPtes8/dL+Gh15
ZFc4VHhyTcsvEKFDASIw1ITGlBKkIcpYh94+eERgEi9sixtq77PCCycX03rhCItv
rkdsIFLhd5lba18GFOF5NOWoQqlDHiMojo0bEmTm5HN7vQfKfTD+7NOVwCrcRKye
q+ncIB5m8NOIzBea5Ph+iOuL4JkCvKsWdgAEKPjoSBLkLrgIeDn9Bx4Kol1SL67B
LoNx1rYKfWteVw1GiRuFZzfrZjHIgGYMa26esm1c8bNfQ2o+Ld+bQgdSSNJ2N2Ks
FujlL4P7puX8RnTQWA2r+ShG+vasSaxGzR/J2AgY13b2cQ4iLVT9pPhMCwltbU/s
K9hAmzJcGm1XUOkvJSizLBbSHLKUdSYpdRHZ1VhAfNHD9iIqPELDmb4gDLCWYXbY
thkrfUtyQuJSqFU5F4n1ZOCxtw6Ho5qjmkAL55/RaURbbNUI4lzLBED0hikkJCyH
3wIsD04uBVkdFsG/37vnUYOZq20w/yOdTgxNodB6sa0tUQ830XTzVhBJ7WB8xSLs
Xi5x/zYWeY7TlD1gVJAod0VP+8+av6rAT8TxkJDPcY88iE/Zgs9nyKTucSrTCqfb
sGT2El0ji54z9Y1t8KRbQqkHwFHvho+wY+PEP8gVdFzevZus/l4paz9f1QbAOQZ3
Z9ksWTnttuX1IOvPT66UXIDqxsQy916BkrkV2ETwDoiDI1EOD5n8mAIMfHUFih7s
5w2R3aDSd4wHzAJqwa9QL970l7FpegDLYaW5iTwxVbGkBRnZZh/GxEKz87sI0O8R
A4ohKge0SkezVxxHXp9yihuHDm7GCLs/CLdPTt78vxjSiQJXB/lrOCu6d4dAu+vp
6WC4xUOjkHOKPhBQG5OZq+I8X6CxTFcVPxheaYM3aPU/6oabGdDIf/Prl6pO1DaB
hnMYwyc5UzGz/7b3Y1cL7rih2sgkcIAQpdln1+eX+lUO7bW8pbIfaublKtnEtELs
qlRywkWH952j6tsdjQBieENKvNThP1gVbE1bJem4Gf0r4CLrD/KgsBX0+lALoKwM
6I5f90ZKLXND6RnDFwIKy9bVpebYbuM/GQPz/m9swWn/pJsXd4gtd+diIh4GDbzW
Z9SsPbGYRjEBN9xqATKfMoYmg0YTRS4aAwOareYOpYjHxhUPtL4ePYvd+f35KVbo
HF53KLRrDmpLt+EoCT4I1X+7IWOCsNTeP+Gzo/aSfzQJMTrZmGHuY3LZMOPS6oGa
2llgyBXJSp1swfyOoOW7xRzw+e/xVC6nJNeCbJ2Nb0VVoA3DDT4syFyHus9IYQDb
+68SSwiabLZnlvcqcQLx+YKmXJk4O5NNETjN6Rb5JMFT0NEiwVcx5ouszx8tVLjv
6ESXWhouq5ZDQIs5P6PIYCK/CkwQEF9+rVdUQo8Dpmpfq8ciR2WY/3k4ifem2WOJ
iWa6bhEy5yuiiDSGqwfJVw7bgrGvfnHf/OVjibsr7d4/uJCYGN2s9xEuGgwp0EEA
UD4Krn9FCSI3WqUro2YhjLY4VHQTv6YItS3x9BwFjqpKsQG9HRJMCtJSCaR82YZR
LOhmAlW/xF6NEWdFu44lo2sdn7vXmlBBC7PFmvA2GKxo6w5UVP4YzNIFrqhcgxhy
lurZM8ixK883gMyVcQiX7pNLcy5p2fg4+3NSJGtrz/mnM++Ue5MSEnOK8GtOi+VR
pP8yWxw4IW9EMHMJGeIifuFvE60FgC6RBEnbamskafKgTCM8fkSXYfQVA9auFCcE
942fdoVE1TR2zcM9PeqV9DZQcOcvsDgBKFzVAiBdSKHe4TLr2vSXUK1MsRYjXUvL
3KZVFErndqJSC292Itk8R0VbeYnOTEGIx50dvTsS/Fg=
//pragma protect end_data_block
//pragma protect digest_block
DGTLcMLvsMoBtyynuOTxXzkGxNo=
//pragma protect end_digest_block
//pragma protect end_protected
