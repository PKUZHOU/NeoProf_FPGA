`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
Ky0NUvmclq1uEwLAYsO82ST+ZkhNiC/bu/OpnAPlbb/qphq5hQzvlebD2VnWPgFD
gYp9ogSg+r26EntDAuDlHtZeT+MIysP3DU/upp1TF+TqMpcHjA+hXdH21Dzl1tmT
3XPBVGY0tI42hQGOQhDFECm/mlFqV9M9kfIog/uqLUI=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 7120), data_block
KyuvsLF95eBs+uyt3JMNuP9OLTkYpXo4ZF/uUlPxN0AXYlTjhI82eeySgr1bfWWA
WO/5EPOdZqrb5qOb2X88PrVeizMrK4l2LEYrCQVcppVeSLMShA3rkg1np+jSGxuo
FwSt9Jx/Ik6v2APb/Eu5fWN8K1Z57yiP6leGcVKdhp3hrL8K5scbDEXhY4wUNrW0
5Qo2mCneO2SJfBrqOU94rpIJ/bbPrpZCo+wuzipQRTNlSsXeg7r8DSlqntkVDBVW
+6DWbDDWLf7C8ghiyTRpiNtpJqBOrlx9AhGwcOJu88O6hQqIhm3OZpYi/tA5d8yI
+nJVn/f3hZ7xIjv4qP54vwPL4oSz5h6w1ZspeL4XAIatR2CDThqdOFwVrTrCVV1l
TXIGjJTln4u6V0jAymViiy/0NDD7YVbUpkzKgyqz7aki9C4TwO14vN7fvP6L2Lsw
azMB2znT/EDTt9Zn0kdGZLKu6Vr4+PlKugSXTjdOy/WUH1KldxdZCzfGVJOEFq59
STfuabVbkLsg+trB31IU20Qi+EXwY2yCpJ9iGkGyI2RXyiw3iIBYhHcid0sGHH1l
wwBU/typkEkcosxnQMXEChtOubly+3bWiGHFuwlFoZl7brYjUJG3PviA7UgoIrTI
/tDvE78457T/iZVKMWeFaShUaNadx2EsqfxxV7tW7884UJpPkziPJXbBuxZGitDQ
esvQchUlE+7sdJnnpTagTJlAQDvfNjvEhbtfqr7Iv1WCqzTImm21zQPfOzuEZznN
Fvx0dmXtlHoHIs1TXVZuK3FWKHC8sUBJZFVFrdHO3mS7QmfViLr4BCSHEZvIR45r
++DRjhYOaONTUZJSj2bFwDOUdybT//Bzk0b5IX5JHSBRJbeTFM5ad1utVCRpiiBw
KyH26TSUT+psHTz6D854vrQYx7Oo72Q66QYZpME0uK7WzpAdpS4cRatiR2j7LPf3
ZWc08qjZrFcRrWmGVQmwbZKWdljfl8eW8gSv4+kck2aZceUaU/j/pctqxaSeYqpR
Ox3A61a9mUuKO7knNK1J1XrhQxeGv8lC9kVeX3k8OzrbgehTis2tax3fyf85wRNo
rKqUZs3M0Pp/3J2IC7/m4exmXrZtcgOM3mYpASTIR26q9XUbh5GYJK4HEr3XTv6M
CCvl3T//pOoeS1kzCqFfTBxWZXMYiDRcf3WfWa1GvaZRwA8Uw04Gv2UTQABYeAYp
s6BS6TRn55Kkw26lMEwktdpw98WXI2Eg7RMXTU74OhurfH6PAxgH/HD9AZjjw5nE
MI+vgo4ReDPCWK/Ip+NNpoO9qSYqOzltCuHU43VLrZ5kitYsvjVO9HPpt9+gEdzc
boRccDQG9pHWh3evLM0L2w2lG3AWVauJ7OTAWssdVyH4kjPVO9yw+vc41mZ+5Ewk
+ughFDaFaFX3Fzd/xDU4imqclPImTfYJdK6EliyxE8d2bx9rqwVtLyAQEwm9Hmuz
85ODmcxHosHT3wzQheuGMX95xuZSoPZ6jYOMMIA/e97h43qDodVarpv5AmpHbNWn
oy3V2bx1DlWHiL1+y0hMEb6U4/u+bhMOILyeMmXIdAHLjPi4GdI+MULwFL+8WAvq
IhF8jItJhEJ+TL0HbgU8QVMcDqVY2n2Gch/Z5tVdMGHmEDxh1M/Tpx2Q9LBf8ppi
MbYnp6SasGwsiMtAZguVJDkQUvQSnVtVEJwgm1wu7yr7/1f9kikUUKMX29KrjalO
Y0HbQVbjcl6NJ4Kq2lM17j/gNAOgnkPsB+5efglSl/rX03f9arhC2VbHXM1MfjeZ
N+O8tTnom3mZYTtdCwQXIf33yBg7PgEyzytlZIoVgVazmsZZHOXYb8dsjaoS2kp6
ch7Xchum0xRKNk/1Y8QhWL1MviosT4pxUGBhykuhaibPgHSnoynUw5LgHpdE9hYj
aRyABKEY3JR+mkq9GfdjJFsqB6/rw6fifhvxVJndKxuPY2nyku6ZgmeD0jDqGoTY
I3zrpB+T9+Rb3ABZf+/2dn8G8iQNS0yxFYiBNRVljnFOIimZ5CDNSsoOlmf0X33b
iKcDeShd6wldISAX8XGBogt0X70HSqNWdWCXeOFdc5iF2ervF82fT5mINsG0Tccr
2DqnL9ABd0p7frM8hCDoIdj3fW2URFdPyUNeT62iGjawlRuLHP+aKwpkRPh4I1Bh
AJsNNC1X9/jYV9NpfeIuCT4/y42n+qcYnBEMhssTZIJVmudkC1ZmP6GKgRbojspw
8UPTSBc6hvZ673vFWO/OLBIOtLdpsSddAwa6fF3ckSve5ItlsvEJJ90MyFpSMKxP
0yVRHqYAIpxmazbYqz/EAdEGnQpVZBEM7L6fJvIpriGQb6/taOz8BHti0qR1Cxeg
OsD3ejXFTrGRxqhJnRIP4DmPcy0Eg8sQ9wcP82WkMb4ZgyGOU6tIld3o9nFswTLT
J1TCa78OGMM1AfXoB0Bx1N2uK5DDRSi7UjElhye5zx1a+SV4YB7uyeE8Txteq9pR
jQqJ0r3dI/BvnuxS14Yc5Mb208oP242tFX+aHVOUYJWefLsYFApRTD2hg0RDxvga
Ckizq11FPEPmt9l1NzU0QIDII0YOLHhYPqC8GwCxzmjUfHWwT2NEEOUD5Mnwrbyg
nu6KUFoPaGLDfeRbRfHeRP6hBsOEMvoZqLfFkEF5+hbVSpOJM4P6TRLRVf530Q9a
Hs5xES/KlBgzdG5T1RE+Kl/PH1ptCBF350wYQHOo7cmWqzAHQWEtZ4haQxEOvkBb
b8vokx+JfTfGGuElmQCJR4MXx4lgQyc4jJ25LCeclruaDZqPcS1XJTfo7U09+Meh
t+mifCL8KG1U/pVktxOXdgvRuU36xat5Kmr+HUpXkV+ZPHVqQR5R/pVD8koW8Dw0
kPGo6UT3Doa8FBcf99ivN++M6Zp1bmq4m0UbXWGCYE7u39aIWuavMyo11GAQskwr
sMiGlBcO/V2MuMf4X2LT8hZEfDOfsgf0YxhfBkzuFN924bjYzo2Vb8i+wyjyVlm6
UETrVdXe4l7Svm+yzu9YsufhFBOSJQG6mpA7dO006oru36Kj5vy0s8Kg4OZslCha
gOZECQEwK24i8iyJ6RofJR6M4M66wJs4KVh9hphSZedXo9NNVlpWgSmSVltPkViU
vJPLiK1uNhGowgUhG6oCMSk//gVYNSUK8hNNjPApQ8ux/6D4/WwVYdcKMG+szTRq
fcvLTJoEs66jmcU3JcFRaa9w9xEqZhtnhQg6Vswlk0ImYk3DvlftwH+vCtrqAXRB
iANUfsdCKYzri9ZlICO39eW6v/smk6yxOuD4O+b1m7b7RUbxjhUjpMqB+3v6RN4y
Ik+717TG67wqP9x2q2DhA2xge56tTtupFj9NJzn0ZbkAOfiE5Jw7fSavkpP5nMe7
96EUg9eTh0YPYyfXS29V8Z7oZjqEmdpqRfA76F+pbywuuMMS3Ksis3+p+kUqgglG
k0Ju4GV9nUf/X2X2YE7FgsozBj/JMN76bdhMmmPSpzouxGvQycHvTw3k7dGJ78cD
7a3ZSKk/obRCgl2NXbImDIBLH1hFULT5XboE6CnAC7oQ4biq0UySQaJBZVifjE+e
DKPLllHKuWd5El8otM/VcUZUh8s/zTgpAthq7riwIIdDBj6yrxpSm+rdVwBD84Cc
2kIKMU2wAzAJkHH3s427Zv71Q0ggWxojz2/9WPIIoNNNdONfgFOE70Rwz0oLOl1s
HhIyhT2gNyzKXKGVWyMBVc8SFZO6sH6jSBl9vEGWv6Sahz01mQsKx7jr+V3SEese
QMj6T1PSPxkc2kxCyU+RoWIHOQQNpuuqP8ombpbRKiMaO/eJrg7ojH/zD1zAQpty
HXdQ7whQqcjuRG3Zc3p6zEM184pP9JKvQruv+9YvNKYx9kzeKxBp1cneRr/6hq/B
EJWRYfxrhPZG+PmMA3AyeMHLcqA9fNGeZD7T4tNJ2MqChQxcXXjvMGwkPl9X4QK7
/kI2y7a5fiqleY9tE1apA1HDXaZ0kPdT5kVbXor/sB7y8urfQhok7nbYqGh920L5
DzmI05dACEjVjbYHYmeYkJgcyMIanqzuc8L9/2Lnm/SLdCOrUFv3lOqaljd8LMoH
/oBMv3sXuA89fpJZ7WlRCoi1rhrOBtzOi3+eJmt2Y8fHRvXx6Gft3Gsu/cwUpBT3
rX4jzz+spymNAiSHr4udu9l/cH6LDF1YLNxsu8IOqBHve2HwooJlyWuXFDSFNyEV
DYngYB8+P9D3RGZRChbmfXOqyxAsHZdZcQkUzvI9kbvRwksxcpYO3mCE/6KYs+YK
26mIAnhiBLmI/FiDuTBhFQ5dArZZeJ0em+DCpdGKryiVjeHGohANQ9CksjeSdXZF
9DVlMAG0U9rnrH10CiOVvxJ1XrPSLMpzT0QndLAjn28aDfCRkcWSil04wrkvy4tb
km7DcqXPcHxiU2sc4O1a1nkq2D/28KFDywQitIFHw9IlIxKtIOYcIzLc7VXBZjCw
uugF4VzRvuy2uzGtzzYcoM56q2+ooKXMsV8+f+0cqj4eCHTetK0UkCTryDaZqrjk
Qltxh3SNfJgwcXOMQFL+fp7GeYEy7csilpFw2AhV0FZCPqbTO8OhzUTpZTs1rgeI
t5y8EWnnYrWEc3h2bVcuVW95108SxYYkkeG9WoEJROi+1vir7H/lP3nTtP1KDC0J
jQxQXulh+seVrgvsC564E/wfz80io8WoBr2LXfq32SPGjI9GK12vglKArRHsLH8T
a/K0mz/eqdAeJD+0TEIDibB7VEYGngoyVzoKUzifTQkeTPk8wdAlb/3G8usWEzJw
GkiCvUbvuKBM6sJW8hPpLh38fUP/t9obvxPSsQoW4LmpxWAPfQ7AqxJpudW7aYgT
e+GXeCCrSUMXcKaBTAZhIzpUgeMO19PNngv3nhKMwVQS0M5XDdO24vpRsjkpE3Sh
doUJ5i6AxIXVWC8Q67cZNeQIEPDy6t1m+H6MLS9IMHJDO9WZrKzq0oZlBG4l4nyT
NNY9bedkBGiEycc3zIr5qe0ctToQ5K68UbWmBD2xFWVDIZsNmVQ6QRU2Y2uoBGcM
PVHsaVHlvNA9rFHu2PMHDaX4aiNVMWx0y05sElK166ayerXAbg96Nas+8ygSVCjz
1MgJBvgNukMiUAUqBBaXpxMns8OUjieC0QdETwwF6eJA8fwJhw50Z6NQZc8YoFFB
Hhe78FzUs+UD9u/jaWISTRgS2gE13uRJTFvQZr7CPturQqX0IZK43B+praIumK3l
YSxsZps+FAmnTzOkKZ4N5nlDGvhBaOzKU7BJ8LmkFb6GG7KdOYN1m4ejU95E40Gb
+d9YGO4MgBsyMxXhUQUby1IGokumigVZJINegSy4YHoLFvVyqkVmgNRk3bSmZKQ9
Z8e7vqNSp1n+7SuulroEPGNx3vLxwVvOEit2I6sOgOLYQ8VO11eGbVsFbJqeCrIa
ox5Fw47Umuc3KSGfaYoDW2ZAju3P7Rd6PDC5kcd107M7olN80ZWrAJIL8NXE8JiL
PrGUvUKyCu6yLiD/B6Fkvf82vo+97cE4Dv7RCbSDgnn+JFBjE5KzJIzx23YckJDp
yu66LgM53J+0eYQWApTBJMKO7BVQ8/VzyuXaspYBLInRnZK5uZGJtjW9RrXA1c/S
3bcANFYTcIYs2nkr6la2ETcsUtJhXVxBkr/zzoTUIqGYEueTYS8nHTRzgtZnUZH9
eTh24x70kJlcAtsskGQE5Pe/filsub70WwGKf67J7anS/m2B55Kyb/DXMSMei7wO
ItecwBjvxmHsqbnYukiH6JR5YrPskP0lLF+3QNFvf9sFxjJfvI7Q3eBkXjz1ZBtl
pZkDgQwvd4SS09s1wFIB8g97tuDAp0/IDgHqnf2lGayTFhGoH2BOjV1ZE9JIfnlS
pIjptpNMchGjkFHkd9s0NwmnewVEUS1CE5pmH27OKmh/3eozPlLPoKTyFdb2ybbj
QksiYyCmezUtYicbsXepq6/vcqKP5HY+C6bmsmIrB2HmGWqHNdqIveS03UV0Pq+m
BgBspJjNgOlQRRXQ10q8jnyUiYnUEYIu0ufeo5c7iahM8E3PMx4LkoyneaVtqkq0
feksV8fC1XPAAp+EGNkbuaoabMUZTsH0hWgvvctG4tktwkwOugak75eBlnOm+Cpk
lIl1hZY4XV/PO4QkaaIZDFKUTgynVVBq+zyONyA/85JAWib9NSx43gOwYvKxaXEa
ot7DyKZOSPsOpdx6UE3IQszGLs8Yuw46LwLOQZEhtf4YW7knIeCf4MM2HEiXL3Q5
/1sdD154EwxIdPj61w0scOmqKY/ZhLf9dYb24SFld2Sg3Qq3nvCLaZgKVi+/89JO
CCnCZMFqFTTWnWWJaG1fgecOvIJmZlG+rYfpDE7LJ/W91p+j5RWuVNFh3rRTKAnR
cwT41CdpZlroO5NF5sXkeBsrmVVyhqegaVNWnHyAuUv4CmW2zfG5GSCaG9FudA96
QyIyXK5SmOGSmRNKnCefzNPsd+2BzPA+QRLMPrC5fyNVzmxDtFYxe+xc4PFOmJam
7jpq/sbm4aeXtXGJ7A745JxQI6SiWhHq2FRottfxE5QkUkCXIuwodXRGFDz+4wtj
WXQhEPrkBmNMjfHuhixsqUsEiPzYRQvB2NTsDef8PjUm8Nnt4kGSniiwQz2ThgvH
Ib59sm1Bfoe14dcIT26sS5VXeuJoo8F2FN+43OcJLGf7MhN0znnjrk8ldCLy63JP
xqBnNtYfGl6oK4wS471lIwBKYPuSu3RUfAMS2eYkCaIGp5LcJdh3yBcqGE2le6zk
phz0UHzmymWv5ETtDw2Cj9rkzGBvcUxZCfvUU4KBvbhJMXOCYYwhup5u1R38R7S1
7H26LpeEYIZ0vK88rUbx0uZ+mQ0XTjaLrnTWn0HaCIVM1xTtZ8Q6dsII2hhtPLGf
2RH+9ZBSoL+nq3R1+JcdOaxmDIVBBv4Q+q5+6ziDbRmKL5+kHlS0gf6rJP5UKQNt
jKrU+CRqep3p1Hj/SjSOzfWNs2jRA4HPXriBoBIDILQPh2QP9EGz4UQCrTX5GlQm
U8xx5Erlp5dnNVtsCnFtWGQOQBxf1Tg3KdA880Ox5L4KwvwVEXDlkZ92Lvd9Osop
+6qh2LS8dHwH4XgXd2sJ/jWFVArH/XeLr2sf7S1yHQC8VRBHR+usDSi1sbBXgKQy
trTb2Co56mcHxc5fCHm1t3awfzjR+m8NHsX1ouGtucpW1oDTi3Sr6BfKawDPq5yL
1dpiyNzMJVTID1svo2+YriUvU9RRcSl+Q5WKIXccvQLpoDpF9PCr1ZfhRL/Vr/sI
N4+/L/+hl2syP6YSRfD/bQt6BXjoZKEu49E/pZMwBU1wSFoWJzjdPGdRwIFApvcF
MRmetuNqVKm1lHxg76ayH+OhWTfHYjBjcvC/qxNrvGDMuz8BdJj2OFVdGpaszYns
/2FQghWe9b20J4bMGRXlRn/FyQHaQ0/DZuqbJfCHCMarFgwqe+ykABl4w3xm3up1
JWTDk4tB71FOysGchvSvpjenhJsqYsBAtJMlNc9IAtbGqGXHZzlfvUWwhoS2+wja
I12pB70f/ZqSfKtBdgjfBzJFcNdYOOq/vjgcly249lprvuf1S3yGGF0jrDIJJf0X
5sjvGb0Dxn4jUZ/ZQfxUO9IZJUWsZP6Cc3lwX3/uwnZVtGly3wsX20Buxx5nujTf
VvnPWeedcalL9LuoB/JqBetk4u/zDtHjxrkPclMTUK47CIvXX5QAoFZr39aDR95a
3w7//yIek/QNCPSL5NQFbmJ0imsj8Q054TasKTSqMXcu1oiPe10QlOj+mm4BiGOz
7axQeK53EDpwr8XcakWDSDPtBMtDZCGdQIdAkCKcCa3X7WQp+FAShKb+ci48684h
2OLrYfve7kz/KRJ+jadpfN24qePDgLuXkn3mCP6kZoPHY29YXE+NkFEzBLoyegge
YHzbNV0OUC3XEXR5fZfWOqWsZGzZwjMaZ8U4HR1g4UzxeZxtgxgtxDeuwjR1QHCS
P3p1WiQUHmJoOp5YLnhvH/2qW5Xhw8MgD2hMtXSQKAs24y4oEro3XTVyii3seDHs
DHezFtxqIAwTUgra3W3zOmDDWHt4hwMHOIvAmx1VCC+hPIEQSlXrBJZ7p0CzC/8i
1JmSaNrBoTNHMlc7EJNELOIW4njl346Pk4NmCQnbgYm1JhR7jvs2eGiNmSwzvR3v
RrM+/fw1KryBrusrXY4982DHrKm6Lgs8QKN6+D1rv9mtIcOsPf5EPM5TQZ/oIqf0
cnH/uPU3eChObKaUhP//LrTnA8equ2bfybUYoqibGWQL2fObjlCw8MzTIhmFZ7W5
ltpm8irLnv8tXCA6eui2oqtFCXW5IWMyDuN0DpW8XnYb80gwK5/3dVY6e9Vweuvc
OHTcwLnUJDYAbAxjz3F13VDMhpHxtFLPzLBx7vZw1ffrR3AC0DGedO1/xUCogveQ
6jTIto92vNbI9jj9+7x3ecEb6QH6fFroWcr4YHx4xiZZOagPbfR76v4JwdzdYT48
6unY+3urJpPj6CepnznaNQ6IzSFj/PJIZGaUqM2r8/5xQjJPyX4uRC4YkI58WX/k
m2NsZ0pqaLRs8VIpH3WRm2QZqylwb2G37ughOD22jIdBhH6dUpY0+eC1BvFTImMJ
VD5TssNgKbuPySSDOOQGBdYdeRB+q9uJvF5ZboCKxGcsIBie7hJZZ1ulMWGGfCtL
PfJDRaL4R+w42zhquWSGMTJPyJ2sLIvHyj6LBJuJoV9bO375VyZiYIni+P8Svo/F
k3y/EEJyUBBgx6Ub19dAeaL8qctNi3IrTd3JgWiEkspTl7Z21D4Im4lzAX4g1BSs
FmikhjuVhH7zA0w4XIm1uLrynikGZkBiFKI8FzbkZAQI35iZckWhgGqeojxA5GN8
l5/FyQf3Owx+NqCAVmOjjU+J3uJx7ImLddk5mezmqIGk0e2Qx1WZUgbBdJ6TqA46
ZDxaMepi8HlijYKOrORtgmm0ELbwJTsolla5XF2HmVib3J8wO/t3klrnagEgyRNW
JjWMBOfWeT2p6LG8pMa36uQn6Bg20o8W+vUK9X1uwcRH0meaqJfLfgqj7a2+YAjT
4L11O4ZFnYG1JKYdOeRQ+jLri18bgWyXqvmvFbXNRvF+au4ohpyS/4jmW13LfUh/
eNtJtci4maDVu/QZpTOabBl34pCQZpyj7Tq10g0KL5iITqE6x5qLL3YBkqZMZ2JN
fC32NbzolN3RK/it1qTMeTk+f13iL1VK5XYCPLU5ymkdWepCtWERCEkS9VqdKxQD
FKjYcrFRBlqMrmnJPSoQWDSaUJPkJNvqv8GYq41JFcsK9kvjcFLPTufi1AzSjJGl
y8ZaPsDojpiXUmsX3jF86OsBNLfLyR2VOK/FNsHEG+LgNskR55EMjx1RwmN+kNPI
4QGj6Nl7EpXqcN3l7anKRfo4848xdYsNUtTYn+gHj37Zis7ZsTZO5jBciCsuovtF
ZgUdQpl2Ubz3W6gJgM6mCA==
`pragma protect end_protected
