// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
GmMUq+9Cu4opEaiTvTFQdu0Td+8H848tenhH832TrRO2tfswRgjFCjBT+QAkzSPVnIVv5k7bd6UW
/qId8Xnz0LyHbzh3PulLT1gQ5v0CAM0BYAc/x95om8CBuej4gufjMT1LZ9RzTuYiSvKPDhQU9Xq7
ltBhyKdwvGn5saaT+nVO5OREwb1Bvv68id0tpV+8LtO7VUSYFkFBu+ehSgrlMEpFZtAKLXSMiDLj
R7wce1Up2UQDMZ1BTfrhdnZGkcmR5ge32IWdNCfP+Jc9mI/XLqLr3T7t8lJzQ4b9XhKlFlh0KTAq
eGQdvY0jy/W4PRkeXduzzgf5Sj1DPQ9ug0EsIg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 11280)
kQu8kvehzt5RZxbK24UrpZ0dXK43neMPYsQs1cfGmcmSuxbaxqCAhtpLt09i8VJHD2u7Q1sF1Zia
7Atcd+T/TJsMtX7GQsahNZCBGWhhzcGGxqZYQqcgIay29NSVXlrRBSJawelWHnFtavOoX6xbANNF
MfkhXOc0FrWUgjsxw/nZ0lkjS0IgAGWexzdS7LFL4g/XT6AZXx/lOKuyyTQ9srpAchh8c7t00K08
4JbwKmmxRxhmQ4TLWXsZ5acL5MHv96FiFa/DalXpiVHWaLCf0pXK9WgHTcG3Oxtz6Ymo6R6CnZX3
0tpLeXeAb0owpDgUauszf/O8eHdMTMpzVTIKfP85GOT+t/Xm/FNyioilDtsZLkgIiQ5tiLOQbNeF
8xpFBXTewB20dahb/8GtDJtENVQjN2D+n0ycQlqyXZH330H+jMrY1lRjVNRHSM/WGKQPz47zDnH9
ImEAorunlDKDY/xsucTPd9+ZOepK3i4rmAsQ3gghoFTtVamlaZO65OGe2/8tiQCsGHQxXMqnNrjd
VvHbkpn1ZAQST1zxdx3NZWWnC/46dgYeENAbNm4C28M4JEhrQySEgihz7+LV5w+yIeK41wL4ifjz
NJ0IWrVKPWcz8CD0GZVlZjtGXQ0hdNiQo+LkWW+3vqxQZoWKejpHQIE6nIc+ltehe1s00nkmYec2
L+54vqhx1rvB7y2lW9UlBByxePs8m7Uqr70TNyLLTjY4oXHygflqGcKDpfW1RXygg8cVDU6Sjgy/
9+MukOI51Sug0UMbmHgb+ydBvbtuE4gPgzylCCv7EMhoqDflvoGXf9ycFyrMMG1Z451aoHxEtLOL
zHMpB7vbTe1xCOkIJz9R+bK1bqNd+NtP8ubgAubup0E7GgoR9rY7/02nFWO4zCq3A6Vxaff8/Da9
FfarfGNo7wqvztONYQ2waI+b4Sfrm3YJbmgoCzceLapLCqYTSDkeKGe0KF+nZG+bH9UV+YJbxYXw
5JcCFPaMzZscAyB9sYWOwPWSOM+plQuW9tUoNXF0OC1/RFuZK9GoJhOVOwCdv9/7DN2XcY5EXnYD
SCj/C2icELLhwgDMT0/kUkGZL/yiH5KrntRqvCvckfAS0oUbYpCH/l9gVhJcq815uoB+QgTnunW4
cEZKcXsWacbUI5ZCt4bubb15CuwUje/8XgH424nIdBmMeRkxjn+uywYITFpJMCZ+8hr03QGJryw4
W6nYKcM9HnDVISJsDXk9NTdrQrEFYlyDHYmvZ4h3im++tor/oaCal2TXK8BiwZb7ITzWYAtvqKXH
2kqgPMIoPRzM00vUlYbgM4hyyDlG7WPhWHGEuIzMxRrD7/HaNRUp2QGLQAZ3LlW3vi0VBg8QRTAO
HDjvXWXh0MfcLOY96SSEG4jQ78HV+4CB4s+Ysf2Yqkxz35bOpE6TSyC1nZIuvFVP/sP3FhQqyg5W
eScZEISR2XTZbbF3vss9ulCkBXE4HfoYEmDpb4+zW6U2lu/3FEBW1J2YRLrRgqsaU+i2eCRUmUVV
X0AcIZLL4WbIGAWW9pQ7tAHFd+0kxnU0HiKPNrIXnKoAIVFlXO+ozMILbAv12Owx5kEKb06jljtY
46IW9Btb/wk+7AMkYNuc0gyjPNwSHIAU6iKh0UaovMw4bf49kcicykGPy3lf1p4qxhscCn9cUpAi
eNpz2bwyqjz5/sWXXqcXs2JZMBATW8idkj52hFOx0EpHH9uFLAVN+OSu2PPRo7/fJpIOktanDzOc
2rTpR7TUuLXlO8rFho0NlrSHRxvksY7dalIw/KdgRAD/n2u03dURkWUBHvEwAFVRNRKKrx25vGzb
L7uz5JS0kku5nTHmQfh4dRrMQu0hy7nos3Lwl1ZaVc8WepbwSZNLGCLjzHAD/kEKP8LsHANJF4xc
O0JCrGoEKA5g7u4t2SedeFN+B6U6/CH4kbOEAxXQw0zIM7eIiH8k5NURNYk1uxoNzjL/TBNFulrT
Gb0pC9qu4tFcz+hqmDx/hyMmOLn0Ro0HF9uO7Y1EOeOcH20ze8HKQeeA1wpI8EsrOrwxYh6zbMx0
9Kc/NeR4Ohd3tSEH+R3BEYQiwMMOKkMYuJzXUdcH8SUzr4S4V2a8tXYGDhwz5+D7zDfrxCdwL0g9
yIMJhQgA7Y/FLr7ekqz4bxc2se5SgYY1eaMalivhs9z8Hn/xp9KDNXZv5l0lpwC3WjcJ0lRYhSQO
HVqI1nmsJxIuvUaDmyt8GeF7b8kvJjUZ6Yp7tBdS2CL5HNwQMbUOec0360GTkrzzKG+VAQIGqX8I
NkKv5aDYprOj9AaECug3G7nqWRVGmH4p9HF8+B/FZ7bF39aAMRuqZ/9+e95bRdFVPGjYe7nCSh6E
GIWEB+uWWBqkVFG24FdAJXRIWUeRUCKvCqeqlPYLdPkJuB+/zvlbdwpfN/ZaQy35GJid3FyDRdXa
ZcL5t8rtRCPAYz7HTdTBW4+9uWLwo6yK9Z7TKox65MTQUI3LZIoTlyikzQcejVljScni2WZlnxE2
5wFZ7pRY7ONTCAJTL+OdWixUZBRV1J9weRgDQJpdWwiG3Lw+6DZwjz2NLdf8F08OoJbeK56iYL2L
3S8fDslO3YNgbsM33GZxlZOpPUw/Gl9QZgOzkq/SgCNkhkOLE43e+zqULJRgTJn1JAyNtC/R3IzE
+3rlWTQccGB9NP+Oz93BiH9bEzWmURPoz2xXSn+g8z3if4ZwqDlgugAN56P1bDdZRRfu1UTPQhG4
1VMUNio7boC7t4kjLl1Wb2k/hAy9BBDHWu0ABgcZLLdf+z6ee1c1uy/9YVCSc1ep5GUccgBCoQ1j
f8M9pj+cL2+LEV8fx4VmfVY0GJsJlUt+SYLvyyTAhMD+/2ws5lpXtRtTqkUY7eeC3BFK2Xconxrm
6wtla4qYWWr450AUcwIFLvopiBOr7sbcfbpr3/ENxUMhvxXbMoYbFhWN9PtKkqddBROLl2jVRa3J
/PxieDOmcS8iP+DwRLr4PWDaei+AIQpgog3y0gYMA9w6tcEESVk3TZUHYjoHZO2gL5/Ruh8Gf5il
EHZAc0Be4VUYEZRcor5jc00M5Qc+5/Gn79tSxYmIOdPJcIfPtUVVSkstIMKHe+MuErL0mOd7qBp/
jumG9lUbYn9X0XLzHT8mmrBHOLOoHXxuNOk17c4kashu7atKXH2z9hRS2usd0d6b2B5en+v0pzVE
LU5eG7y9TR7Wq2eNkQvY3ary2oDKer08XACb5TpM/jrUp22XuxSlmDJtGIUE14CqfcqFUg/4L/qH
jfEBAUDhc5Tam9lg8Z2onMMYG6Cvrdge5NtGh2KaMUMWqA5x1H1ouOf2GGjGt6Ap8nXyXHxz5v9T
fNb/Rf+NnxKywkLRcCq2j7p9HFQRh5Ang9ffJdTR4tazYUkmmXvZwFjwrl/+tPrc+0sf4gBkkEtD
Z093e3I3yKmWRGV8H+/Ve3PHLCeQ+RNePXJxZ6ETZREIFOGE//90THDtitC/mRAG8lDg0YvSfZWa
Rv1nO49hr4un7ybh6Ok5PPtX7MbOmTgosvdl9NWXiY/vXAgUoUNuDESYVkRbUvOMtDxYOQsprFeq
r7vYHQSGzkjRMfhIJPQkSFhPHRRPz8tGtNVKVL/vpWmZl12s359WV/fwzHztSmX6hSEpEgIoaiuw
6JupAf2ZHf5UJ+eusPLKWVJQfhzS4u9uxyNzIItx6VhGgXe0P7KtDDd8dfge3FR99CcznIA5xSRf
v1OJST29wz3fgnMCAz8XJIMwMk6X1vK8/8BquryLzxcJSJjW6S0AaL/hpizyjPkAUe1MwYMkykxU
2WOSSi23p33Du667xUcEXJtNCeBsx8J0yyU5GqOojiL/qzYaDlX7wLXWiUoIREbGzN5xGVujEqKw
i6xHDl3vRg2W1Z/AhNpSI97PsdNMe6+7p+aiHKh0G/X/F32NM74QYbscAypdHyvfvbo7/Y0FPRir
ViBqElt0VR7mirsYATDYpAWrUfiX0fDBkdp4LjUmOsP140qQ9DvXlQxgj5EvMwEMfFNZF4q6nKXw
nrsrU3Ianmoxqhg5fX8PF0CRK1t+VX6N9S3kuHnZGAWtMQBux2AZsLNIIqIrvbPLx+k/EdkkG6zI
lknKIFEqzShg3FMDEJPaGAaNLECZmhDTZlTSDXaz1Xn7ubtgN5IexiXqmsc4SB8Cg6z1fyC/p3js
27DklPCeVdsul1s7A69AYjtazIyQAW9Cg3gvzdiC7mTVDFBpVjZ9DxGTf8GDK/XeWikWyxD3XfD/
cU0ySkGWlKgeIo8WTRpUgGJtwk+lmrRrW0QzVf/PAegE0OP7GoFIljCjrYspvclqiP4hohgS8N13
ZNL7BeoxW2Gx7qbt+yqEnFKB+W2fkqvehUkNhbNF1Z4Hl6jDTc+BMNNr7523nuP7bdkQ/Xd2fqwT
gdek42wJbJqSd21yyiqE+d2qy0Rxd78Jij8JqE6N2WtJDfuRIO8EtVMIjBu7p3WcprpA8hpSHtRQ
5kHgP/y3+GsXUCTl+KDhVIZtrL3Un/egbhb3qVperiazwNWJ1VeST0p2V9pGBdFY3SXqwagBISzz
P574TJsD4rR90fI27jReKfsGNNaqz/NBj9tG/kmhmD1G2KJ02aiud+IyDt4VE8vJ/rrcnSEi728W
i+Oew4V8wxQHdKlU6CvQZYvVLMsEKdpMtXDWeh6ikBjvNNjQZiVdY4PaSycvFfTGKyconTS8/5kL
GRpU4Tzf3OUKjZn1pNt51lhL2Z3We2/JbYspHR0c3BvZcNA26dpDZXUrSaAa+VvLCM/BPu+C2SAQ
rmIvDt1cMh90H36gN2uU1uoubg8mT8Fv9C8FsgxfQeZ5czWrqcm5rxPbgD8E+EZrvFlJaFsLsuYc
jcCXtt8YVEN51BzKI2i6EmNSbktf5VMJhodQhOB75CCyKxmWJFtrl+Tl6KXheAEjcbBl5WcV5/YR
PNx1E0kRwlLMn7foJt2b79++472FmOYwvs9wNpl++5aPwO5rvXda5HxY4OdFZkMB3uf3h575msTI
fbMH7ro6Vn5hpJGTms1kJ6ES/SjLmYtYatYEt8DeahyyByUNT+gLXlqDXuoC1XAnsqGIZISXC0C5
pEzSGWESPoAglwMHKyxrK0hmDYFis4GSJal/xamdWHY2gsx1wfhhpqpRcDZVOZdB77kaQs837Hsk
PU8VYVbiSPJUpx3mgxTNC1TXxlovdKgcAj6LfWyGJHa1OTpxbeCMEfPyFxyIJ6SYCEBG0aqLqN81
6+6ejHPFD+lUsW4be1lEleWozqpWtOP/54b5dcsGF51Wp9HHF2gWt2wXKO4EcOdOByQ4AQ34bjT+
6aP8xdEMuDIbrZIS8nN2fiW+B0MPjAaBy8kehZ9Di7wqAmfMmCwMS/u8PTOP4ilYZu7yxdLstLC4
+zNgEcmMgg+Zt5B0gNUYcWSp7Nt7fAWd8jIzKSqE5L74Jd7J5ozy6rV+FP8xNnKtgps+PCFJQ+xK
c0F7oR3tzMLxjeO0SEOJvJujdjauc3tLTi775hHfC020tk9qis79KpUZ7/1EcX2lQVcR4i1jwXNq
bZH+lSmsoat9gQPcEpG/axGYxU3tPv/+ZRSetTe9mld677SmcWJUkfT+mmi0hI0XUxGv8PWCrU74
9hjInG0QDU9laSDk43lgdtPnHBp0Sh1lW93eD61siP6OI23yXDIVNFXLwNZABivnqr5Fnoij3Y6B
vbRUYVgskJbBnqdHub2leK0UYynFROYV5fhJalhudlUftu8IntNGwUnt1KAMHRp3lEhsg5FJnvUu
BEOwQ2mTY5hKcRz6l/cbMvxQ32vt0Jwv+0YNx2ss9a0JcJfDOdBzf1kgcElie7kHQ6xTrtZ6DMhi
IR2QSVwEisQpHFPyieIikCEupuuo+4wAIpUADg0ZkGrjmCbpj2ArzTY6UoDRmaUb4t9rSBoFytpT
jEmo1hA0QgnYWMMVTY9PnsGnwfk41gvYoR1A5er2osHGhTNK8oPRyDL0eIIxc/ivc4BXTphT+/ED
pf9hzXYblobZgOQEPGH5chz1d8HDLd7yAO/lW8vJxw7iwLzeCTf1WfaicJUK+C3ipHgT7K6nwmWR
33OdE3gkr9p9jf4JlsEtbHS1nTJpkfyJPvovlW/CXi3sS2AEvFXLMfTkDlaGoPHQNrXGRvj+4NUk
2tNh4+yNsg/2HplBG/Xq5wUddzfA6MP98kUkxaGRaHVWyjJ8dUzDXZBqE249N/sQGnhZoz/yhOlx
FGh3m+0HfheWOJlkvG4ZzI98l0dmQSU6Xp0W2fbr8fSK7ItFYctKUWODjoaz91IFoYu+XpXGaPX3
qBMorbI3x0nyjWISal3cab/n+HtLUbl4dDARobJfKodSacB762d8TCYmokap8jm4+pB0kfUV6nYE
9EEdZOqx+owq51CuoZ6FxGI6qmJdQCAFxk5k7R61w9lild4VcoLCQ6cNg8w3PjLGEJEYXdVHCS//
2pa3u9gd/SdcFMdPt6/EL2e410EzYhZ3povFvwba8tan+DdzmdvTWSL2G0UlGHcbvzS6mmiN9JqT
XaOYqd2CWonrJzLYbExIc0TjmSwI07nkcDur1NYZ68ImXWt54+uQx3SAYu2K5mC/xcwR/Sal8iSY
zYq6lMlJ4wISnx8WZvSkNxkxQ51izslQLCPTD9pux9JOEBYEqBeXg+qL3pLqGZATnewKy888+klO
NQI+juxLpedN8iDQVHpBh/UyGGGE2yuyxzD59rDVs95HjtD54+UbMzzRBxdUt6MwkSRcJxyz2Osq
fxM6XfPRTZ9MnZqVrlW8IBL3CkPa6Jrw2h4HQQcZZRSfa7/lE2NIcqiJrbFs8b5Db2KxTmdEFApR
+IhdedxJ3wsRfdjGlatrBCnltt/weszFD/B6IeplyurJPPzqOldD5mFyFc1Ra3gqEvVTm1CPlMTx
1+QT9DDfRYyms4pHnplO+UBXMdcBM48UB1A/kcmj36zHeELL8Zz50XivQY49w25ZGDDTKf2GIdGS
16tFEqQmQa9oWH9MB/3cj0J3CACnVfmS+ftd1lOuYkOTlAyBYyXhP5C6wzaqTmuPKErr7u5Jo3dI
2NX01hhX+EWF/fWY23XYEvXi+LDV9LxxDOLGrVIAy6f0Q7VIMRDZy2TJxOJYx0SlC73OKxRkku9K
xbPFSSVSWebODan2bpqkTFDlmGsL6aNM9H5CuAC3i71HdGf/2GVqgex2aYsA/HS7s6MyAmv84jeK
NdWJjD/ecewwt6ehOvF4MaI3Yrhuy4S89Jn3KCOVjyvp2le36NoQUWlNr1Ylv4qHn9dwLRWOs0el
OE7W7GhSA84DG+jA1gWuJXJCT+h+o17Ii38K1Rmv7C3jTJIY/IdQr28fugVWIy/+JkV5LZYHZzWh
B/zx/H7+1TaGNKGysMFG8wvPEIYdLffT82BHOBBDZneuq7EURlEpupwCNomkAs2O9YIqEccxq9g0
upism2SiUXQV7luy+T7a5qS49uBq8NMEKsEPAEurThrnYgQag11UVm78si14oTspBGJzqV2zrCQo
BMgBGEMaN35DU9JKNeZ6IqOPCATGzJWzlVtggNhfatsWSUI7BOY+FhXRUc4H/SwTQg+UxZbhd5yL
hRXAA0HMjr4YJzA+ndh/uQOjyMKiri1ZbuhJ8P8EMJO5JdkdqDxt7Fnsgdt//+rQEQVaMY6zcNlE
BWLIMhIgPYP6nVNqpQNNX0j9geEDYBThE1/cbtHipog0ral2st+wm2UPCvHWgsYWtvTAkGieNByI
x4IKvCj6KtkwRIkB56PsHYYX7NZX2hUWwAEFTES8AbUmt6K+k9Q/rXE1mLD7yBLPH8u/Kol1yA0m
K/fcKyiRaGUt6gIzsJm7PSAPcT09LTL2vk1+TnVAFbeNMWXymo8cK5ef4wlu45vBzZjdw5lCV5Id
8JHJFppYjASobKK7xRg3om1juLJtelX6wFf6O9YWGNQ/6/3574D46RMc1ntiMNkguDcmsok1m0KJ
FJW5lew5Lle1hisJIZzRzMf/R3ys9vlBMPQT+i7kJgF2v1EtuMzq22/QXgiSkcJIM4HxFUX2Cu7p
ZIzgK0TAEaTFQOmLZSGXBaj/tnw3Zj8PlnmLJkvG2qpxuC8n6X2EDhb9LUkFg6toQZvIdriXsrgK
N8+BFVumJgDIzvwptQKOJAOqV+Dw9L1F9J03ptuutjE1UaJN8SLP9psaUBgI9D7LKxPGSNhS/z/l
FdDncIBDew0Xpcy5MMmNMgWXTZXzxh7uEpusPMSH4l4IeVvEgzSYOShkNN0TIJrKSXh39NMxwBwt
cu4XzoHugZRHl0tO5FRe+FDVCUQ8i3E3kTPUa9hxn9WcdvSfQWlJRqLtda50w2ZAxmgKRr8imLlT
iDsP0xy54pPl2uLYou5XaWeVUrlF+kncvHFHmhlv5xDO0WGJUFGx0qCO4hy7dRDuVmgWznozW+c1
l/UOHKjhDvyWjyv1NxwwopxqUELwft6U2kOvItxBoRC5mbyPJrYJPveCOdaG858s8WJucfTfmr+H
XsAhl5FGkawFlheqkDrt3OkTZEFnsi3aLv1K1pWygqT81F/fF8rBu364AKUy5av8U4xLuPVjOn39
6DwnFZOhrBcQwWA6uDAOMzxub4bxof6P0viRl1HpdeDgVofCKNtVv+k4OWT+0wLUhWr/m7mFu4It
XECykCDk7A1lQI71gMMroLlIND74EowCWw89YG+ooNGOQ3JHpjmkaS1+CA/t3nmPMRAqA5N2AZA3
rkzrTViFMiL7wz69iL+bk/OqFt49y6z7a+oMqo8H2F5loEodzYJGzymG6NigSVFxwxh3i3b1qT1L
eKKuZBiq+OF8g6JHw9GDjJnwEdV10FlEj1bxHZ4jWZecEp77UoW1IgobzAiyWLaOhvfyWlD2lV71
m9DwAOaevtHfhEkAlhkuthu9WkTx7jFyyzrK6z7vrAfAk+x4I0xEuYHpluZdU9UVYsei27mV5JXs
njXL7WkPhEo57an/U7oTJyf5bdLJZfWAPyhnY2U910QuzyOLTa4qoAUSv6VMjHNe6nUVl0p7vech
GVvp9PMN14UbDiewIm3ShGdHd6HNcwcCMwACudZ6nAUbjKoTjqlWAqDJMoR7bxSLYN88b/ckIaMH
awCtqSJzEV0XK3E3E/4JgmTd0n3ApXyYY/m1PU7oKVW/8HnFnmnX7dWEgsgZMl9Oueh5TxE5upOZ
ZCkqLb+zDWuh3+8GhoysOdAcXw7aWzttaCJZU2MS24LW0hKPw4pCEFBuvZ24k5vwuIHTVqBGRlaj
XwW+cLjAER/NFJfowAyV9UGshR5tjsG+UC+9QuHhefDZwgNBkwfqoPZ5G1Nv2S0IhzLGF+A1gr6q
InUJ+uU/wsbjl71bvpDtbnZRtKqzG46xi3AqegO/FKQ1OR0z5ra434zfVjF8do2U3y6240Ps6fRh
9NvHb5FMJHUvIcEb1XCU9t2ES+68c3L36T95nJfYbPZlUcVtgCHPJVY1wtIPltptxiO07Dyp7bWG
HxdkeeI72PXuGE5NrA+LwamNFFT4xLp+gDIm23N+n5SnJbrcVjFp8YyriwhDZHzxTBjuLdxDgzZb
dWrpwwhZFJM5BKaLmzrDU13w0UKRFTr1wrbyPpIvrxylrfwyJ+YMwbh4Elj1Ygho9RXqdnlFAmaL
nOrcktke/p1lDkVcLIFqD/D+nOQEXvh68CSLgdQ8ORo3dCb9PW9C+OMlp6eBeH7Xw5tAHnxb4Co8
fl8Q3px+nlY8M8wRJoEDJG6SiUiqVVxj2c8iQUpIKeua8rA/l+XZ0wJnaMUXLj24GfP+9V2ypPgX
lWd9x3q6ZKo9h4DF5iAJ/NpjD0cpgn6YYx4osjcogL1e39UXwdBQATGUOw2Wnw9F7PMKcvbHgnRN
fegCeEjcaHb5+WqPUkDQLGmsUkui1+2OgznUVh1ihUV4qsgwmY5dS02UviALglIpBlvCcTiyI3e8
m7LfGjk9n889lMc3hF+K+Whh5TcstXXe+jgXK17NitKuHxt3WOeB1uS5katpTcdMpakR8qXU+p7V
WusmXvMojDWGO+qo8tzZukxehXOKHLnAlkkG3bHd4SpbwhVwTSnEDM5g9tlwaAaN1JUCqZOSWUSS
vXYJ0jnlM39xT55k+YDO0BgQwKVDDkJtHQvDf6ueWU3IMwauaGINE8YU7KCML3KIVVWsiZeeSxyv
4nxZfU3GtX+Ag3XZeHbKg2iE1/BY7aZjTW7JfzJYkhAtjSXGNYKKUXOKQjE9BOBOWe/g2LcYuIza
PIqE/MeMDtv3HrsLn3odqrA7QWmYWZ73dfMtJHPwWS4Z3XyMPTGWY2jlQTLgTJQ/9dig2GIaJuQp
yqaEX3WaYHKFVhudyUOU1UT5J9s170g7PNa5EInolvo+Jji3PWHzNrA/Ux9xqfPQV9oxhRVFE7Dh
rGcuNeIYzCt1+a/NIMk0Syg3KPvKWa74dRvmuJOylSJ1PY8Lnem3nbsmNEgFou9eGQP1KuTclLT6
oRXWl6GyplUS58CHupcHzKUQCkwu92ORscy3tUBdQ8qlttWULL8BEXsfdDpbbfuSmPMNi6x9x5tn
I8q1x466txOtkXlGvJdE9YuTdT2LAKxg9ioPFdcf/Z76Tzc4czTzqa9ViMGYH4whDStfgASoBdEl
4E5t6NdzSEUMbF0Vcmu0Xs9N6lskZkN/54J+2h6znE28vFyVhe/oSOAv0NIjnJXYRbRQx9S08Kh6
CKQ8cfzhfwXX/l33ReHSHcjV8sM4rQWZwrqBfAoBEqcZZJzFh4Sl/RpJPA23kl/KmsQh6V/Hclrs
Wg8j92Bu58xhXRlKoDETzYQwYrbQyn6W9mDAHOSSUI9aoqwiUDRIBiWbHgqXlARkTO4nh8XF2wDj
8/0fgD2kKkG2YCTwna25pnUkbWysz0sbzm54RUxt5Xi6X893SfFKlCHA7t6SGb0BZIh8p7gfLH2n
rhjNlYrk2ckA2ga9JKNMlAQpCcqFO/ZXZEuCyJNiKkf2PdfPojGIlDQIgY9JrTeg1v7CersT/6Lo
zQUxcWEQq3fj3DSmUhKlwMedjuLRv2Jx+KMmnOlzyN9YQeFzL9MpaxjU7SY6LSlfqMpvsWvBGo7N
C3vU+ed3mGRpLeZiTR129Si94QbjIF5DaZO8yozRnFtv6l8z1YTyDT8aVBL9D2PIlrfuGaI6wvay
0jXTscP20WWHbCKzdceznxQHfICnt5mGcP9XVq9sLwDFWLtyaV4cNOIL1ScJlI+wfU5XO8Fyy47T
H3ZXS9UZsPRBVcyo3vGxv/YNhnFItpCohXzfJaZE7x3gJYAPVkMZl74wD+c27cjcgn++QaCgC7ek
dOORvLUIX+yMVJkOtjv5BjDkFCphShxmnDsq+SoKaRZzcHgkQTVE0tH7kBtJ4eKL64/I7PrzLGEu
0bhv9V8jV/sjBD/MRg4c5+KGxZKFtOQ59VKQzwqiLanwWzaCO5Y28p9xKVbrf1m+ThG6Ac50nq/z
GgZAX11QkdKRSY4ipwz25JL3abcSekWLwtWY1BxbdhuYuuom4LprCt83RRup4hoxdoFY3MHOWEcB
7lXpSuR5fOcwA8Z3yUVb75jVh9hQv0YfBZsv5MoK0KrpjuJMLQG4X6y5im9vYmJ8zy0O+XHPQ5VX
7V73bdSyrdfDivxLEVdjWb9DaqHD2FvOrt6X9lzAlk8bpMNR9Hjx/ug91QsYdxjQKuLwStgYC3vL
sPbejdk/E0F1XXwj6qZTVezYCqpQH9o/YhgtM1MGakXMILqzOrDMIUiLOYhbQhX0f7yb9He2U9FS
FHpf9MI7wj7ZSAXoPDnMoUIf3jIGatt79N/Wj3nuLp7h/4uFRjwiLl3pIIZkc9FHwG49DDCLb8bu
nUXlvVNMaWrE855e6bhKGODQMVNItWinqrVIj4Rihk2L3Wuu7FH/e6d4lOc4st4rrmjGTTUNQ4xi
GOOpw8i6coYPJrPYCq2NL/sH0IeY3lDSRvyDrlTFgTrgcbAWscm1OBAXMgHixYWDjnDvChwflEYB
XYaAW1kUdSaopbD8uMz469HRONDr3VRCvywzck+pNYFCMMdKdeVFogxbJ5THLKAQ9d19YEsAqUma
2+JL3tXYw7U+hZXv42l63osIf0dgEnaWHsUqn5yHXMljO9KfTOljFuvWnZx60ZsLNnXlSt3KF4fA
PyKgLRqEcmrfyZ46qsQ3/6IGcGoMh+2O9QDc9RphDS1627CLpCLUkWW+ehNije2ePRJ/xEeE1FKh
+N/TmOtKkO6wETcsF7ag8Iy8hNIKDczMjy5ZPfqQVEp7RqbOsJHbREmE/0R/6UQ909qrj2bT4UZ7
mFCmjupk2Ur/doeL94bJY3rHDaG6kOsxnIFehPLbJP24vXKtLNY4fuxMkR4CJlRqt/m18faSZ8Ej
g6Wo/ydkJRo4L3cZgF6YXOw4zIJaElZrBKkqurF4HXwkvrjf4gsKgcInPRiSDMcYoVytjXsQllaz
3LlLHqaKML0zMXpB0qmE780dgmWj77hZjmN6U9CoZxVPCFXtLU7zK9pG2A/Ojoo+k63vvxoIpF+o
ERze08llG7ljSWt9/TuHev53STN52M9vIZaemCJnjg0UdLbyT06iaF6I4yqix6b8e+joHxC90sfq
iAmeHyZi6jsllPZIEgMjjl2MTyxeIVqgNN6YFRIsdhJGQR3OCQSL+CfZFUOCEzfSTKce/dVF0Ih5
5nSrtkywTXrdHDARIJpG3wcxVPCSfZjVMpDPpYBrWUc3V16or6/XYC+zIJt3LFjUVMOJIlsq4jX8
rI+NrdAeFgnQTbGkFla16WXQWQtd62LEEKLMUmsLoNQvrMUA4+MlpavHjbea2mXLcC39xpyI3+Gp
IkSu7C0yfcG3fKjQDoNPks7JW8usXtfwTRhhqHcSNxxh1AAfky9yW0h3YTYeWkGPkg2Zppuydu4s
VMmvjcSH+IGVZyPCE9dTDoLKuhSEaUVWBwTRtJJnZzAjGwbJ+GBSnTjE5gBdPAk0owaHkEkQlyPD
fNIW5dLRMdMV2TpSry0H2kRJqcMQ+OiOuWjLH3YHWnUInXKkKGnD30k/Gycjk2Yaovo9aYEXvoP7
TrntTO6LES4DSIwZfGniiJOKTd5FBrhPqi6Z234zZu0zTkLsSIYkXFkz2WftxJDmZayLYEdtqTU5
eLolDBiuRMmh1Nbo+hxGu98DJnrYdK0FRmhJd1ar8txZEb2vN1wdfU9zwAJh1LHzaESBZid8iu8/
bh7q823W9HOG79ulLtTiGmyBLTdhOOfCLlgmV4veOeE8arNVQ2IYSxalLg1UC377MLrV3Jxtpt0E
PEKLd4pkkazNZL34frJQDiW1Tj9QHN8BgJNw55VcS6Toi8GKPdZsbnVphfUreqRYZVjlinvcuGWZ
Go4xOY224xvbjzqCHRLlw4mFO0m6hSlZcq7OIqgiziGnnFGNasKUYydfGPAPQ9q2I0W/bdAyP7dc
KP3sM90TALnsq6/D6VV5AQYCcvn3nrxdFyoeATD3qcan+P2kW9P23y/f7xkWyRLL+u4Vdia5n0l/
Zy1SsfiIGX4KHDODm8eeo9wD3734uD58uo44rR2AOAdlpFFkuB/z6kE8VWV9pu7xhRIGajPDIr/i
4WUB7iiHXhDxCsmfzW0zMjGgp5wAED4ZyveJxKHqHPQKv/DlQrp68PumguS2RXzdIzzrXUJPlu/E
tedwOmFu5fMDYtxbUSMr58zaEv5qrS8iWe9roI8vkZrR4Sg7hTiupkKbJVjFIY2AVvCRkHLY9Z4m
KEeevfZ7SU2pp10RjSa5F3UyzhHC+VjORDeLBQiffdU0R8d80R7AhgrqEhpR5xpBFr5ESCXxWyrP
LeDuDcUtehzeJA3LbVYPbHvE7YiZXtdxQUADxuM9ixO5tfGIavAw78Ap+MWpL1hiAW7hRdzoq7Gq
KB9u/bdcpmaZGQvhasAUEz1CwZ191HuLWuYQEWbxKx+NHHqrMo3cL31/E31RR5NBC5WR7Q20ky1W
Nxv9apHdsKG0TjKnCIZAHhHSmUaInCyopaKRpGS1eizg5sW+ac9z7YCTXh6KJRw/gagDpQ6eQNeo
/Fw91DZ4VNDlmcy7R2JCcs/Y4kI8Dr8bR+ClZJ5KxoHjEu81qyau9mWPotM/PzwOGA5G6bEpmlu5
0z0E7PQozXs9elMwBPvSctWnctAOfvQO8/BKO/S+MHxoF7q2G5Rk+ioDloJ4LslR8WBHh27XlItQ
Js9x29+QK1lFMyLzKmMMbf/Jvi7bbPNF0o1Tq+VI6MLUn3NPCzIJ/sg9OcO0eaa0gr5+exueJGM2
LaKL8ebGYDP+qHNhNJGmIRuTqLwiwxheXT4OQA7ul67/4ypq42Ll7MUgl1kJc328R7+3QUlJEJ6L
ODtn+vby3KCFZVhtDHaWecNf4lq5Lf285FH6CAsTRIVhhy9Q5+iltys8EaC7Qph1TXfU6c3SxQ2K
ji4a2wkWOADXqu6R5l+K8ObouMqKlspMs9VYv+ulheXQAag1E5eqSzUPMpg+afbV9PlSIG+tUpkt
ATZttHXbpwr0oyLwsD4jT4lLDcWDLbSoLcndX+FBR5yewzGexBUfwy58HqLwLsSA74Gijo9ptYws
P7Ju2smsU7YCCI1U2peTntBHyXnnIGjOifa6w+aWGdJ61FPWxdBuVcBDcU2C5lGU9Y+tGcfo/uLv
v7mZr1m94dv8bTbi/OEvzPbA+KhCizaqTwD3AV3sd/E3cjFWpTqRS9BoUT6vd13CNDs8e6M4N1nl
UGTfm6RrYJeJ9LozZ7NV3e6r8Vow4w8NYg6WBGHaeck1ETKyJg/y0EAX6gsIcIluVGUOG6htSDee
nbPJgtg4/UQ6nP1bxMolW7adA/VRDONeCt6fs6AzcFRbFX5Bej94i9FuxOw8FENmPoERNCpQho4H
xZ2s5G5DC3ZG5SGvDp8NY+f+W1JAhmO5Lr6mGOmaUP+KBjSiyW4anRgmYpMOjz4DEilGzPZqdNGT
Da+0m5Bd8c6CDQG4S47DXZ49ORQF64i/v20KIsM4wbun1/NslAZ3XNz/F7rXEJMkUsgX
`pragma protect end_protected
