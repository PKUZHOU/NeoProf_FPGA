// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
qSLJ8YtJvqFIYTKEFM2tydy7wca5K2wmUlQMIEW30+4o4/Ci/cjQmMgv0yCQG/1L
I34Avhi5refKhsJ+iokXewRALljULVyrmu5cllimlyIkbEGl5A/aimCOh8Qce+yt
WX0dVDxi7tnPwxnox18Ih7oLakXxriewx4P5naUXPJM=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 8496 )
`pragma protect data_block
xZu+nuzmYdr2MHi8Qe6cQe6Du+VZFA6ErBNl23JfdK3usZ7nlaDm9JwruJY/QOb1
AxyKkRYnClAEeOKfUyCm4750wXCmDJcBjyNo4Fp74tQWtQDCiOfLdhWlg5cVsTrs
g4XkxYED6SMeebaPdOrriseawDjACqkbuLIzGpGxyPjn+KV/W7RzEW5FgdYsSrw7
I1IgBPggquF7r5dGlhoJuBxPNc02UioakWWbvqKUkYKHDYDVChzG5XPD7ka9jd/y
MwXon8jtLn8QzzbcL85y3ED2C+FgQFHZr8lAOn6ItpM3VOpxfuBOepOl7NzuiW/y
ko5fg6/eA6zh/rxnPr0tqw7Hh9Yx69+axwV4kxaXuE/fcyBCzkYyMTAGhDgitvcB
vdk+pMqKHJfbCidBDf3OGFw8D7GLA7+bhca4qfHj1PaxWUAWaCDJr4wtn4Dg5tT3
De2zR/F8EinkwD2dTS/klRhpaIHRy1MGieTV/64eMCZUHqLsy+z6J9/MjhpWBBXm
mqk67dmbgJT1It9OWALrE7vhXII8Uy+ZrjmMqBUJwIdici0VIMGmClAV5zvwErx/
IFYD9QWQScoUHHlqYRUg/bqH9Tl0gDQXaU1kchdSBqjJOmuG08HxMrCrBAMs0Z71
V26Rn6O1bynaLGXRt1D5aLYrV5QI9+iKWeypjl7YOneR0i7+g38UaN+V4q5+Ac0G
DHAN2Bb1Xz6lbOK5HUZniK98kk6XFpBivoOPnxeiyu6OrKnlZFWJJvd5ITDFU23V
SiSOomXM0Q9FJV1AYCcjklwX0Na2OQdnsNCvJ53QaJf4tqU/ZXeg08pdWZWetAQP
CVku0axqft3/jb2sCDwsm3NWTLdJKOD+kVTJjQ0aVMGz18bhO9LoOzRe/HE898R6
tcN/nyFqZsrpXBxKHC0B2hqPxNOy53TvhKI7bmYmiz08b2mu7H+E0WhOFxNPdGHj
AlHZhfh0oXkD/l9ZdOM49KzpDK01CixbPqZC4y11bVgmV88R++6Y88tNJiawRKpU
eun60MNvyRnISpo8dd/yl6kAHvHPZyxukzzmm1PYF1bXXPZ+8CRwubeBOVwY1n0s
wC6yUav9X1BUDaPivqmVNm6krhX+R2cf+fqt4yY7JGDg3351YrteZoEQzAJqaVSn
gsLkHsgyzKzkotOUtLPeHGqgPiglGk5bg4NF6MA1Vy5ghuHJ+bmScXSrK8zUW4bP
yK37+jiBcXVnJsbPMEDc5hFV8DEzCOh73aKmNe//WnK/X2XVLh34dxC9PoTG3yRr
Xd+8UhKB7aFZyH8YTy1vDOwTiryHdtLfKkvfRbc2Hh7Zr+5hLykP7mhD2eS6nTnk
ttp77Zx/8sC+WubiZVyHtvh5gojhtlhtodcRQwfFhtlEOfd3k6nPgHGJcVgklmvA
rDNmtuelCd1h94bjlKCR634pZ0U2KYAgCcPAWvKCK2VWbS29UopPaWvOjXjub7vo
s+xuHp0dq2Gr4L3OUC15ahpVexlICMCjLBvybKFvwpJgEl+VB+19cjw6rERx7cKC
4FDgY0D00R7wEIFOLUmT/1BCaQ99Jun7urImI9IcOJp5dKzhiKCXQtBbhfvsVQ3K
f7v2TTh5HKf4R86gv2GoAN3759VWvkG3FUfSmWx0DDUxABvb2TDIHJaMFnpppCLU
dxFT73T5M6VOUcd5xnQ4g6mqcRbB3ocUBOjm7lffYWxUQ/k8TgpkX3GRvu6acVk6
EAj5PILmtZVb5bEesD0BQfMN24GneqNz9lZiE2tMHIgfNBr57LxUeJNsdWrwIQGw
zcyHGmbqN8CPgFe/m6n89DD0jHvmlY13Q9VT7HCDs0CWgxr/yDQaiWYFaBd3qJh0
6rA2WuE4vRCbLa+nvYwYDumcyHXmoTDDyAUAsjnKDlCTUlAMmynqRSHzc18VdBxK
NJ5SAKKTZU9A2dYwhvJ/mn//IPuDLwDMQecRIjn3kjxQG2OeE+jG/p073+8okbLi
gpzoOe+8Ka95Hb4xCZ02Y2BLTBwHZpRqzIuR+SJiNssmp6XlQLgea7fviJiDV+NX
rWR3kjCVJIYytxdLQJw51gHGqz38dP+RQjh9K9k5SCPJOvwqdfaIeswwFZqljY7m
wyF9vp41bkMnfWIVAvzYmd93aey0SCiOFD1laIPWyarm8A9JyaKCAQ9hJiuDH0qs
hA4jRzu02TUgdLNznG8upesV9srYZJy4XD5v2Hf+pDRC6kidVEGZwCokVTaoGwTI
WCkhL8X4sgbA7BY/t2RsPewouqdgCgyU2iPJnECZaeZ+6jBYCPcomkDYlNK7fcQj
0ckPgZRoyQ3H8ghpc3CH5m09Ry0MHW7VWUA7akuj4jU2p11s+npguVnf774JTxN0
k6HNl+N2hyXy5Up3MwdPRlDWeif3DuapPhh1sjC4NoAA0b//quQUlZUOOLfR2/Up
P92AJSifyQbWDSptyFvaDRf6r/EClY5Xdxb+3Ib3Pb3g71ivTdbDj8zu+MknMSw7
roGr4etvPVF4IE6aBbbkNcH4Ahy3xxpn8y5NWZPe2vams4sg0pjxue0FTWvqDC/J
Qcaz5czb/ha55DXCucAUpxTPPxs4J5/yxKYNXTFr9ds4K3lzQfH1LWxAHKJED+CH
YvbyoNa1+ETOk1i8TVYYP1UAw54AgIR7NwHdpIlLIOYsUhGcaQ1utvOpZ2zIkq8g
SsjVSbYeA9iP6fEmzldDIImab6d0sXjgo41s0LDtKgP4aSNPgACoIJmxeM4ldkPU
S076dO9R/Y8J320LSjYtSuzgOc6qQXzMpdYlAbuPUspNpNFd8prsSmJSBICqLKep
QposIRWv/vZ06bEcJ51bjlLKkiexASwqWmLKLm+jdJ1sWDA5IMvNi2mC8YpE/ZvO
3k9CaK3TnZEnXhH1Yq4zNTVlbe4YtCFWbFv55lz10BO3g4mkJx0bH0TI8KWWm47q
QzX+o9WWnamPY64CE2ix7ox0wT3tYk8D+LLuURvWotGBJvpfnUGWmK/U13hgxyVs
2+oeFh5sX+ProGouObl7LC1XjbyiOpOGkQhndx7pVzu+ysV/5X2eiQ+qRkaulNAP
FkA5Hi6hhERem7R0VZTipKiofb/C81EVAuihEgVu8zNyqyaXt2yzC6ywRqSNulJG
mdaoGSeUvddKzMFbKDSsNehJC1ULMwcV9DYgI1E+4+SI+EQrj8onlmX3KleJhTBR
fb0fcwOp+2Jg6OL7sLPhfWJhLEI3w93QVhK1ODcfA4TDUrTJ6u3gYcld2aAPlHfc
8dUCdBzoSja9ShrJAl/v/VQQ8obaaxLrXIHYAVBcKUtIaAp0xLzgSJmr5GwAmxt9
sLl8qmoOWbotj/ff6lN5Cnl6tcNWo+Vx8NObVgv09KjbCDe2gINIADy9jhaS2vQg
oIqjBWTOpQjA+sH33IXWYfX+2gw3ZPAVYFVzab1eIiO0wiAYzpxRbEKhGBcENVXM
MdUsBKyN4We+L+bNdGCMGW6RQGC5UhL0MNGCIo+8Eb0NUXEuXiUZCsC4xI3XQIqd
9tR7ALnyFl+dCcJ8tean1G3HcETcrmzB6AXNWhVKgxmG9YJUKd3yWk48Pkj85sBv
N2hUpldOWdXpbYQbsYGjulvCF2IZvfjaohLV0RX7bmXDKwgf9UNMu2SuQhVg3/Ln
mPNzq9UqP3uKIWuOCYAfA2GBGGVbQn75oepJB2jMGVkSLmfX9ZaQZL77ncc8vXMB
2GqvG1wgQijF3pZHagSwhihpMemB3b/kWVnCLdnd+B4RIBoUiqiXuC+mpnXmd614
XJkc92FX/TQOpPb++Qv5ks0BUllpXuHcxUkoaXz/eedkCMX96ge5YNGFSzzseo2G
Ga0Kp08kK9NzRRH09HTsqjqP21hQ4SjOAy+lUlYv9Qn/tEQgFvIaYT0fsh7DqCvH
2fSNco0WOSQKfrBoJ8WffJv6T23Y1dCWvHcJ7XzV/L3r4MhT8smXX6DnNcK82+Af
Q9+/NgCdm+EndJNnc1xLCILspH90Uth8CClz01aeNGIbitTpL4t3to7Hjl8cFNQI
PFiWMDPNYjxgWwmU4mgtlpok3k1MB7zZLaNQB1EGvtvmKgrdI5RZG6GFQmNT9AQX
zdZM46svSWs51+DK5/x34V08z3jdNM2Ane38BQSghyHhPx1v0+AHR4kt/oGeo+98
zKeZvdCCZIH/dvD082Ey7dRKjQ/xuS8Dpp22p3y8H0i9IKBsm9VE882Zs3UhT1fb
MxLQ+oINU5UHSYop9o3QUupLPyiO/z7ph1RNAGRp8tK4V1EqxmMxJXcSvJeO8wr4
2Podcj/TI3Zw6hkt+yNJxorQByeStZzX/zjbE99Uc3icNYQk/HyOQvsirsIzEhii
sPBMXZWzsMOpX8OKNDeQ0L0+cbFnjsReQGBL1hi2ETxFO2MUh28tHTBgdD3Crp8z
LKbt1FGxVi2mflIDrEdLUbt76ZzPjOUVMjPXdq27rBuyk51vsCb4Oml2WpBMEl91
xR8Olqhs1maGlD6BMiqu8Ii7+TmqADjmOGaWPXIYNYv9UYw/ntKh9Lyjwdx6gcrI
Hyd4W/yUFEBBZK2V4s63w64NII8KniZSxNYIVViu7TwNgMIvECOj+tkrIWjsv8wk
uSNUe5LVEmtPBLZke+V5rZJdH4O7AuXfdGQL9JgxSQ0nI+E2+YIJP6iW062TlstL
Z2yX9Y7FYHkWwWNjn8n38m+QmOUttPmUs+yVV2sXHGroJiQSypzYvEY3LaElstoZ
iZGCCNnaUExcqFpdhNybOXYYB/BT9xj4KRXD37zq5YAZ4tyz5Rd9Povgasx2fOGl
0pZ5iNq7YbIFKD24za6zkfwacjlF7jouk585odVYdlNf/nWjrReJHFj0WHLkKz2A
Hc7Gt9Dr0WUmykmT1lDrkDT2Mgfy8XYBH2MbEEczYywGhpwfeYPEbBhVu4IhdFUc
3RZFOd7bSfv2M8Xd8ZdWTE5Eg2DOSvn0QC0ZW25TxsrzZ8F71urvZksqDdIUI1N+
f6hmpVxkJ4X8hIF9Ki3Adqj+xKSCpN81eyjIyFh51X8eouW76VnNS6guXxGlvC6j
OZTU057n8gHOvYUp8xHrtXibidc9dPLC/ZKt5rXujBWPhl1p4gBcioKcjadS9QYs
ysegtskN8LwDzWuZ3R/JBZRK29g/aSSdOEgv+ni04wajVK3MRvRzy+qIy53FiHYK
Grubsz7/CN2js+FcFC/UWZ6eT03y03sq6lS0mvvslqsjMiCXHS6qoKcU4zYaBdvn
NLbQXRlr/SfYZAKTY6yZ2MvySxfGKD9vNU3T4kLanIvlnnMbRT9mVvsfLb0KEvj/
0zQmPBhXCWOZ5vOfbgZonoyKG/TM5s7+nYikTfENxqgybl/1ajJWEBFHoYDFrDRs
Cfc1ok3eU2T3X9GEVOv1VDreahDcjJbM6T6LwEIa++jzfY5M/NCGdSSOc49a0lQx
Kt4LHVNwmglEDAGJ3Ic3vVRK87NdueaEowf1c5isYZHxPEwGXKcyHiuu72+qF8ho
Rm9MM/hg5MqcxGoCsdLRTUvX7ojy6WKh7FTxRkO11dDCZsDAEG3Il1fptrnfBsko
1KRwDMUlqq5mxZl1hh1s+LH8vfN9CFg8Qode+MNAhzRy90LC9HWU6r4SWm1jIETW
UNzhOwnI6px/o184/Qg1Dg+cnbQX16QOGjEQTCyrwt/ubHSUwCYHsxVPcAa/O3ED
w22d8XDNMDfY/77/qkzhBqrzHr9r9W/pZST2UTmVSG18BzBP4LBTiW0rVry7V+aa
w2GFHx1NY3fbUKgswgzhc2Usu5HBiETiXI5GGlVAx0Gh+6DlKUa5WW5dqVGjOciP
uHwSvsvGsYbPbrVUd4VaEppuoo7WJ2SZuagxxHsfbXbPZca+5HT1CHfhdUav0JDM
vWM6wQVGhDT+k+klCTng52gLr1neOXkRx3aV3fDBH+s7w62Wiw3HXzgABOQFE1gE
AqiAUJqSIDO+9wf52wCEOVnGWQytnquYSithItXxn6KkEewgtMXkYu+hK6RmXrEw
u8/dyH4AZjS9NLtct0WpQXkre1/xIlk0gkdY17saqhyRE4cjOn3xCtQALORdFfJg
oU5Qn1v8Qr7jfQpvPQ6tEqgiKLe7TYPpBO3eMWRTIcFUiEwVDm8DhRSeIvEV7ZhS
tGHKAJgl6VmT3nDIWk9q+CP+lSoC/m06LbRwnUgQW8FttbAAJPck8BHyAjkGmwSq
hkf1XKY+rODmLMGuiD0ZQKBCdVyNWOSp2xFABXkl+7rMfqydCmodDMJelFgrtcyr
lgH0jPK3tCMI7kXlOGWht1mNqS4mlh0iTx4c3S1eXAd3uj9IDeR1+0Fc2svOFhqQ
pb9xTurJTH7JHcQY6nvwOkLzh7uWRuzT2aiah8BAni69qAbLtsz3LBrsBPtLMADS
DbQfjMmuuWhHpy+/mJR1PJiClu4dxPFw0erD26FZQUdtUEjRqmcRqyk9HQfop1+T
bRmxvxvd3TmLHWR/tSMKCx/kZmXiy9QLinmH+sgSc92hjMlOXCjBn/zvCfWTLjUg
4TxYBwpc9etqFFVUY38XjRVi7o4H3UGyNrVTj5vRkPE8NDnAlLmHmMJ5VezRMNbk
R9vdir3ddZG6Dir5K2FrOUvgM35UgFE/yVhBPJlEA5fr2xwdV2oP+oNJcv5EtIII
HsmOhyZZDDQX4q1iStxTEPZd4Ivs48DYn9BzzSFddr6Plb6V012l86t6X8fzdqI4
OUK+psY/sSUUVzOWY72OrQDGjhs7va4gXAm/10x6eOSM7HmKGsMyvwyjPOjK2ShU
/78yvAJ0F6JVA8KE8n789hwG5g72/6/BBLzrb9BknsyeiYaWqhzYp5qTCAig0CWv
ShWhcvq8zhyoKvjY3hmwRGzS92MxqhdafUTfxmf8+gIVQI0HQ+hpD6U25Xik3iQB
xdIx0qrKjdkNOM8T9ENZIWYixmvlNOXKbD8Zdlsu3vkCA2Fp6uYvGR64ksb5tL0Z
hJphwJ7PlDHR+XwB6HwHcjHwgd7HOXX+JBX9QFrEj8kR6b08VK6FDaP7ABFkKK4D
wrAKMPj3M/nIIlOxAcn8ZojHseIceZsof+H6AOFuT82JAcTl+JV/uBtsf7O69XYX
VI5k29AehCM7DqM7CT/3uoHRWSCZ+jzbJIpc8hZv0zYT8T4M+pNy7uQYMqWaKg9J
C+q5wZ1AW5DKfJmDH/5bxXlrVL/xsl3DqOXYr9Ag/Jpm85iNmQAR2lwN/9HMuqYr
yv04v+hJIFhWF5tdrzdPlT2HZuX1CdSvrMcOkjY5Byb27H0tmZ9z2+AiYqKwqdPY
jkkZ5hc/ba94bfTTyy4NcrRdqFaqgaHLOQ6kAGQj3l/Q4/GM/WJxjQIcn1TJ9xpp
WqXM8lc+zVeTiCidQCLpNy78oh9uE7J1Po1IxqCfRNitOtoU1Xy1Zjrzeab5t2gi
nfeTHEot0uPSK4gk6CDEMs6vZJXQHO4qTH0QSjrl9vF4exNWVAPC0u0zqfJxZRtc
SEbVrUkjjr3iTcodpVaj3xyDrFA+LdAM3sxdk9ATCFt2ZQHyKhYdqO6oUiMIeh8H
IegIVm+yEDZypDxHuXAiKTizirOg3A41/1y1Gw35jFNeclrRZ7PBu7d+7a2sebmK
EXvn5qK83G/gFDRzs9rRoO9iRoE8QpdBw7FcH1UwlVeg7MygaEBHMjN4prRveXCb
UZy5uuIHr/HrdqTCxoiC/UHkNmvM5TPFQQNWXwR8WK9mCWX1QJObo1KbsLMnx6SH
N8bq+1JxyVdFRaZtsTUq/OPTwxAXY5kSakJd2RLTyHHaPrc1YR9/toI2Cptkvv5v
UeO6f0J1TT0ZZ6lOiCLDKkAtiIaUZhV3Ol+TnRbbcQSYBp4u4Xds3qfVIjECEdCz
4HUv9gCS86QfpXKFi1ytrYAcwJkBJ+kfrdl4uEbpb5I1tzItfMZbRIZosnMBmkNG
dBZN9L3b6Fgo5jXNm6qWFLVgCcT3a5yRKhxBTxrlr6RMO08WELLujWc7AxknFhKb
w6gl4Wcrr5dm4ypXKZ2lzfj8nVJ5OD6js82e6vUKo57nwQx6xvLog2K2OBnMrZPW
0EIt+AVVye1e1aSp/en6C87aWVbiEHDnhbVkn2z66kO/fgrQY8Puj+d9LOlZLrfe
FcB9setgG1NM+5qVeXqgxN5mChQ4xDznGFplHHSpSq8tFFhLJehbX8sjQK6jWOWm
MVkmg2PnAPYM+GJ5FLNkgzZmsx4sUU5SbqfvbDVbSFdWqM9zT5Q0ZSo625jkgXjL
6r18ULYQPFOYJ4/NMw7yogUzzQp2Pz39MkA8LuYarjf59paYr6ngrnBMoXfp/9Id
EOqi0t0YO77ryBDLMkthjRY05kVYM+38nEBZWIo3stXYsivGKQ0H4Pmk5+Y1Q/P0
SWnRgeiKUwPGcnQMmMkomevj0CYj53/MbZUQ+my3mmr/KE9jmf+uTqg2zPzlAo49
wakWK55DNSni3kFlt+TYXBeyMz/9vf4YgfUGKDKVsOKEBDobEMuZtds3KE4QDNk7
q9XyLW3mywhNhIPqrnhuWVKD/rk1dwkwpktfOSUN+846CWFLDn0J49DBDlv8p1M8
tAva+x98S569zTy7wF6aF+GDGy2glZvf0HdS0idx9JQ4IM7vb+x3QIFK81RhZY3G
6d0xlR2E8MjLPyj5a8kGGzPOjOVYAViYc/niyO87Btwjc/LQeUYywY+FWKNf86PF
D9IqQKKst9/lJqE9Wyo/SdCwElxJFnnebWzFol7sezQt9yHpdqtlUbA7RYw6XigM
I6l8A/ikc3MeB8WvwzpY6DslPJRL2LrDicRGyZaJRUVxHWUzL4z4YydxEAiJFCLk
SgbY9d8XWOoFojTfP92vKq0VFfK7AfdxRe1NCaz5N2TdlLd+o1eJEFQ8CQPgRVYS
bXkTvbDjt3J1YYhzW7mjrKr2wHTwjlxt3D0NHIvLaN03RNH0R92PMbSi8g9LnFI6
mQdr4/gEAy+29HJoR++ob5aQyQK/B1kALs/7YNEP4vMnoVxgCYOu+lmYNcCbiZzl
+Xymfwd3KTX0ZFjXt0p1QVIaeKdNGww8tJYOwECllljuwFdp9ozVZAoyhPsFqVQT
XJmsn77pbLiKsMbRwdg6q1Myranjm10gw45tj7cjgyIXzTH3UUsaNGkGy5x1S0bF
1y0vIX/gPJNrRYwx4TQMF+RpEm+ZAp7j5dq2BaE6jVam7Zyo9A7irM6MFc1PW5ZT
zMTK7m3zeqnrLr4mNopyal7Dyx3Aw8avC9tJKPe12xqZBjOQfu8yMsnWh//xZ1MH
M1Mf84q+OFy9YHvhQ1qZjLb7bLTbGNA4L5b+RD5lrvxiYcWNqcXlhs4ZEnEuP+Xc
ZfbzrYtjG1Dws5jXLotJZW/+zgMo/8zK36Lu0hV/5D+fxekIWQfwK2xPjjffzsfn
r5FHg5AUFl5ENZ4nlolFxralvxevWMKwPWBxp9fPvrDAoN4lLFGxhxsUGpOh94mV
JysvGYnGZoxGYE6QUW1NdLSTFV4Jm5jDHjwjt66vnTg45frdpnmtyMO6mA6+YoBj
X6ojzYJGIrBx3cCvSIakjwG6CxJ9UvmYYSIN9AnhwGqWegBY48xtaBvAbVJnpKKu
ush0/JFSz6JZbP8pdrdgeu8cTkXnlp1CB3GNFoJMQNRttKq1PaQCymBmZCgJko4v
re76amQPq03lpJZCPerOT6eTzgz9KRF42lzzTkXxaJMXdzhKd5fY5RK3t/zQxmaD
3un5qC+eJ+F4ODvckP+z6aK3hr7azxMnOmaVVfVDE+ZchxNWiYHBE7cirAcw2q9c
HzKytnU4URHmUrlts4E5wXUB+qcvlWn7DkQyx7r6JfLGY+5AGGqJCCs4Med/vY2N
oUSQSLSjlTbGRO0YQcaCZnsTpkUXADwOPxX1+O9VcPVs1gcuQzZSBhz/mJRxtx7b
TGqCmpl412uP0gPbbLfRHIM9+J5A+as/GoX2bIr98aeQP9QfpMwr5vu2AJSRGVZm
QtntgCw6OGx7GLXJgMI7/U+uH8PmmaAepLXRb/EsNAvQiN/e5qrPzH9X5dbAJVnM
CQ7r46OzL1oxaEcIJ0Kdt9PVOBWgYRzTqc79dqCh/e6LcNaRDkB7TtCIOuNJ2WMC
AWF+dAGJYDved3XD6p3HAq9rmPK9W6n5bpQvFRGrIja2cXOUmn/ZF8uNDxcPKwT9
RiNi/LopweT6KRLxPoF6HOuHP6b3JlS1QlrXITFJV1vHolSX8lHlbr1v/CEusNPP
wQg8DtZy1LI0eqDpchynxQQmtl9UUPYFIC8E/2Drj+szOyrqnQrwDjbqlmzyGYvl
/W3lCVI7LgwiUn8JoJolymuRbfqv4P81G09ocnJ/H1+pUEHL/g7rMOjGbfIN894D
aBJERcNB93KPNH/mfjty02v5UbpesJtbGPz1qdI0ge9YmtIR1+aF1Fi+QNmPKMrJ
xIx2l6BsS6hxZ/WVd2YBY8g47YvZU+yM4tKblPx/rDWvWcnZHGZt5oCqvtFjWWbs
zOgp367zw8u2/4hNfdTpAe767nJhuCy3NTMESYgo2vwrgZv4i4CBw3tqsHYXzkq2
l5bDzP3CvV4mAS5kG9k5lYrqYylkCOLen43FT3ELgFy227OLdoMQS1ar+JA2GHEn
lHkV0591o/ufRp3PnghMLW3x/+lZscxncNAu02/lsksFW/p0DUsG5rVjHyHMMmla
U5QVLG1unDN6WCVAGPQZavFEEB+FtToe5Qxkm+kwU3RX6cXxxJNTg66kWCLk9VK+
n82Sw1u6kFOnHCg/h281QYNRyM5jqtSlhC/g9zg8CUSaZm+HC8RuB7Iq4SEAvxnw
chpivkGkTSkiUANMrprq8fHdaokd7tBkDm4biVHP8mC76QE5IjNssJK3KKsj3TDl
5kna4q4xn9aDmI3/waX5xyC6DA8zg/icvKdkTMrG4Axio8MEEH3DI5ScPeW0puEx
YdCgnZZzsfzVEZeCuVsQCpCJyoBVcp7PO5iDskhiQNfJBQA2wsx9xWKBVTkJabZV
cb5RA835SHOlya99RCvp4/hk/EFJ203gl26tX8/w5HOrOqcB28evE9czZWJBSttp
IGNjHqARGDo+3Wv46dxQCxAHe+MlH9qCUj/tH2T+McuWU2O1i9vSaSuXWrDyj2Mi
xxo8djVGD2wGeej21yh9hPGGnIEHBFJoIrAdrCSkZCinNR9Gn2Ovlxg/Le1I8Wv6
kJghQY3/Wqb1WmflAgz8I7khEZt348QUYMuBQOY2HnbU5OsohTZZvU01cAxKhvjv
xvLPtiTc6E+5bBEHRhheOU1TFrj/WdJLcCu/mN3tUQVkuxNm+SgeP5Oy+fqtMZ7p

`pragma protect end_protected
