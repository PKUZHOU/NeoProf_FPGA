// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
VYeIhKxyH/mbNr3RP6+BKdpNMh3ZgkY5vPbMC8DvwKH9xLiiFeG3GaeDPUQ4
A8r/jqkV5A3usZ/lIlXzlxfTITYIVv19bg6kMBsN0T4jP15O0FENBYvZMJXt
W7OlaI5H6xdxaYWD4WD8WJKMj6kha4XKezXYRvo1CNdcDBcSGE85OF4k43d6
bAeYZ6nXl+7ZYh/NU8rIpk10QLH+wmHnKPZm9WxX4oLeGZe3VQ0uOkfLmPU2
MAJP2IPbRr5nEYw3SGxTNe/ZODGt3BvHpTXHE/OmSjrdZ41wHCG7zF1Yt6Jz
ZJrDE3OV3qrBHJnS4RsRz3kM4aqT0a7yWZ8ezrmANw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
SsXJSDLnYl1ysJVHWB+BTFYYYGCHBPGDxfrut3oIIJKFzKeuPyPdF4wnPgHT
2CCyYDrY9yPmPAbT5U9+JNfd3Domwd8OZwJPNRH1q1A/ClbXWgIWlKUO5DtC
N8Y5Jn0YM2zP63HgyJ/dIAcww7FuTtjWp6neiJLVriBg8htwmNFkJd88LK0v
KOINylu01IqagkgyM6hAXZKokB0DrBvaimsnpRXLPdUdTR/ov1EaJnK1A1i8
yQSCL7gAfb2ny0BKGz8CkSl0Z4hzYHhKEBUnMglc0npPE1C+sidFco90Aomz
pEYAnvFQyueDk3YNnOcce4HHllnLPNgkbSiA693kjA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
os6W552sUmJ5hoxrR5pHCSPVl5nfUxRmQVlag2rTtyANXzA8HA+uLqBw0IbU
cypmPm0KKCu+au4zl97usLTAQhX+VYLDgf3ddKVFwIIf7qkCZMXQKMPePKQG
1CKjopsHU43GrWRnNdT7okZRTirWrBad13SJACDKJieQX2nsYgVVOMG/I/gc
2pRXOShmZAUFE42mqhWl3dr6vk1cq31M9Rjt4chS83lskzM+USe4U2CmBRmP
ktWyPUCdx+3eYm1uI4ip5HuUr8wUgIOwA0hcb6Fn1E/oEM61axwPPEvlwTBp
IZ+pJBSMLbMTo4RSz/A6uPd1JYHmRtzKfuMszK4kTw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
fOyRo1A1C8wzdvSh/5XjOK8xVB6CZ/Q6/J2f8blh4bi0DISi7JF2j/l1RrGB
2j/BT+udy0AkCIAArwxF+DAWsIIbt3/SFy5FgZFY90Gb2FN/XG0dw+R8ZyB3
m7pL94uNtqVf5nb9DUqDdMYfsM9Cr6AWKHgczzKl1RK+ZtOV2B4=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
w2x9ijF8XqoSpNJodUXYFXAHijifHFPNV3E28IyDRzn5maSwdvlWkFisHeLC
XoKd/jNr31g6H798YDN6RIIkyXSzwEtlMzNIbvS2ssFhiykjKJtm5wRzhrZl
lq4Bfr4mN5C5ronGovwx7yUwFmhXpicn3pgGSFK8lVo022pGPWGUGhpNF5Bs
aPxmLLf7lvsislVut26lofAREFj54qWkRtR4z/pbTmRXlGWOJy5hGSbYhnPs
Ed5e0yR18uUuDJVr+39a4gwm3wis5mgpTa+gfEjUJ0ca4F2f37zLMuQOGvxn
ht4RN132pDdr4M0G1C0/EA2s5FJLNEQVn9jgIH4yB2VMOAz8/k8wLEsogPGV
nm8tOrvuynrweIe5JQMGQRkxzVbuObe3DmnpUt+9BYp8ymNUXVloRhf+PmMu
/gOhmEr29GsQK63xI6tsqKJ2ah9O0wzIYlXphF4T6xowr3YY0MxhgdlboFva
hWhOlJPTS4jzEmK0ldVCZnPIbykWmDNI


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ONLx9euUMjOrtx1d130637JN/eQ/zMxCv3H6bMKLzDCIpZtZkZt5B+qJViyP
Y58JkzlNdF9+Dbkmw7nMMvgFnAeN50EDjVYx88d3sIEa0C2UMXUyW+o2F3Hh
bFG7uWdiBGW1vqnJVFwuQxW4KaJ7nSNIgxo7cFhL9czxlWQmeIY=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
uskNllI210IpsazjUIkOipVQrMpGcrjkzsvwmqBUtH/Z59IpjDytTPfN7hMI
SHHU1eNMqiSK2HSiqbCnxMUCzacu0JEGLoWpirJCKW1Vgf6DCVici0YQID73
PNR3OBif6QwLnd04X5q7f3tQCij6IpGdiOqbAGaG40SHYIckHSM=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 144800)
`pragma protect data_block
fS5JbMbtDMItGoAxBpoUcpI+PFxNalhqbjMofwifuzKJfm9WdotL4k/OFd6W
7erlwgbeft9kvo5c1dUNprW/axNs2XpEJZ5N3wgPCQbWqW+CIWe5h5rs+qX6
vls3lL20WyVcQTvzY0GcflI9AcO2DCONMoVDnPn/ZYQNLWbQdfFgK1XRAn2p
JJW2Jwv0eIInEWkjp7kNd9HXcaHJrnaRm9RkbnxgxJnRFUJ1VyaTM9x8zZ3C
TjM+hnn1xWkFbSRoMx4ax2zmRgmaXfk5GwNuNpAe2jIAtOqQMpM8s2+slAWB
kYv1SAOyB3WIyJR1m+kdMiSlr+FDdK/zoML68M5Nmf6K16kHy7e72R+LrtV5
XlM1CPB7N2Oza12uW1uM0v7OG/fdiiRrJiYCH8RsX386RZUVD9kgmTMoaatI
a94BZZDe2gcYhJmGgBdGOExAOfyHfvHlL+4ZJzlLkZrGNz71wQLJdvAv2OE8
h4GaT/j3vCSOv4FOQHkY3DoK0ezd7itfWmEG9eUQzT/+3o8a60yEQ7MeeLGO
d+Fo/XLP26dfLoMSAetnODRVr7Jv2goijoIRgr5BkQQfYxP9IQP1Bc9ePgvv
qdZ7zVAO/xOBO8bcbbAXW7UX7uklF/2nDRZPhVFslZgPak73yK5vwa8xIr2H
V03/LMYQe5VqWIGd/LlD6u4jqK93oWKWK1xTiXRFSTmootaY1SjXZwX8wcbA
Qhuzva8FzmwBRNIrh2cqbYrUMprq84qzatlAgDK931QhJb33JrWvkKsqSLkV
oGmWsiFfobVzji6sc7yN3p5smkxFfa5txj89Zztjlb9Fo9sn5I8bekiPAXGb
+U8KALXzWMNnHsKCrkJGF9oQspyTfW6mkKx/9kPywrPxXGKBtY1CNzUJEiRd
rlYOK7HHyVbAIxdDh1++d0pNIy5yY68sGj67P7B3DScE7G4adMSwjWbg8Mr0
OFU/o7T1mfOVSoJLSPK93H/sQsnAoQVle0l2++K4R4bi2/3t1jCIqrhO1irb
6yNsRkQTnVesyq7QUHRYvrjKCsfHC3Qx5CIsIPwBt0WJ+W5+hhq+MzUF1jYq
zVwh4aMm3cbrQsy1ouW55yVQkXczHIagGRIZ6kkeu1/jCp4YxcRec1S0GxeV
bG8dM4Y8z+6BIgbfv/7BXYHThMh9aeFdgDjhHrkmJ9pqOR9wxU+AA/W7oWvg
dLNdD2z05fuZHQGiRrZ5sWh7uEpR8l+PObe1JttAa/BVFnRl2rLiZV+lTEgc
vXBQUzMQBd5fRxC0RGxiapT5RG1lgvVFOY9fK9isVkrJVCwO8Ow2l4ICeAyc
SyZn8/aRmW3RPXrsLrPa5XFN0YBkS6yx2AwMLIIb37601sgqZVjK2cUToVIZ
Nmcz17KF36K8gWezvRGqpgQPpWpNVxW7zLJO2BWRRyGkTOIWqVk9Bs64vEEo
jiyvCWS5tnpnFHzHDBYcZDcg1L5aOJVHRatLXAcU2XrXpAOkgyBz90x8s9/p
YAfMw4xY8ZAtEEzZioxgz52RdARYc32RVem0Ujit9nW8nKw7zi9MdwuwFKf2
KKdM0IP4sn0HonEfqSNpQ9U2XOivxdUK5HWZfuOk0W8FiWhgSBRiXXnL+657
u7RbdKGZjSL7QrMmhpM0KYnMZfja8+pMUfeL25+lxu7Fil+AzektnMPXe/Vv
ul7sYNNOy9pNW5w2Lcg7Su07GBk4q/gINV1+8jt9Y3WpzELuYbrQLbvu05mX
DUUtLuTDkREiLKv6J+meMCq82KAsSdkTEmTAgz6CAQab6YnTUYxNKrgw41GI
U2ogR3fO50G82tAhKm0zSnz9/GLGO+5yJeryzNNMA2htyi+Dc0lwPGXrTAN2
lVww/BblgJdsqVjef5D1b8/mf8EloptwPvtMUBoaUlIFANsccKn83CcGEsYy
6uBMV6feq3fgGJ0tq0deMK6LFDMaxkq5k5H/o8Io5wDZO4iptYJremr5YKkj
CnDccUyn2m6EfUKPZIusQJBYVKpzdhe3RY8c6f1R4/0kIOrEOPYxfcZJxFqr
ovOd71ZI3DunwygAaQzJP80MQozq0E/mahrzOFPiOV4aWtuPMnsuyGQU+0qo
LGeAdygiwfONZ73Kb0qlSCfKSKNH+/MwEbUZHyznbDuBvh9tcBiM+Wefq6bo
H0zVGDsu/WMceIQK1qudQS4UdQeJxdMNtqgrVeCeeY66Gmy9jlWr7b6SiC6m
HIVTeQVlk7SW/untM7vPCA0VrLl12KZ4OfE5UX23W/8yQxZcTi4Ks/UNLVSn
Ibd34iK8rZ0GhbX4LZcs5/fEMOGMBWxCP9HyP+MBKshaECe+gXxYfyr522TU
9ldF3SOKN7mwsMeZrSR2QhJOwYE05WSn4iMsvDe8xTRPt7o3O6EBtkknjKOj
qmwqz3ZOtaSBF6p7Y/nryQSn7MoUMEEmWjFrE55QmYHzexFBD71cTjhTAiZb
yBk0wlNEKRqaGLr2/mRRvG9pHFFEaREJJJKZWJ8H9Nx+4cpFZDfDTV0hmHDE
AqRPpTjEhDxZBhRkVc6lOhr4f4F/fw+jF14kS6/3rqar987Sxe7xnJKy3f9C
OI6bk6xOaY88yluYbMUkAFq7hUiNbtE1aOqFsXIwEvvYSkjeh0npeZEpQFo/
HwKvYfQOfPL5iV/q5h51X0KAISJm6LTq6PesXTQkE4Ryxjia9ay3WD0gKdSt
+N3a4opAJTggzDVqOxBIBZRSlHTM0Oqdz91SDYQz7hSFUsEAaYowLlWRBl5C
0bYE/5J4DGaF1sazROK86OFdlGqvWtZkFj/sfXdu8u9RPasjpm6LqTqZ4Qvk
Yat8qEVPyBTTUXQ0X3guFw8nFgMobOJYFMDYO6erBLMruNy3eaO9Dt2UXcs7
Iuvr/s6YxSi6yMajW4IB/mCH4GOkBI8A3xScrAS9rEQ0JBon8Y/Wcp4gwnqP
0PSaZPxfxd1DWUdlfHO3bZnxUbAsnE/T3AQMuHO+lqnS3rFcgObbYuMZ+ldr
uGTH78O8MZpaNFKB8ycWOezppf0ZdCFKRhrgOi5PkAVEpiHWRsFnDMO2FEco
8h1BYxfp94syxCcRnoPcKVWazwozs6cHQOySrrKUoQ4ZtUC54KJYXvykNovS
NPZ0H6fwh0Eu9/QYNKQTD0JAKwGZev3JdoiI+KJ02ipgIuD1AR2whITQK09q
m0WUrBrvP8RYJHe4c+xQMdYGWSmJxEN1dRAofi2wLJt3NkVB4VkRm1rkWYpv
4GAuwmHiz0HGNMQOWY71CoT119fRKIccD3OIJI4RGdaqQYdoK5Am1RHeOYrM
CY7yJI9Upg3rcOEPitgABjegeixOMBjL43nfM8ghWHwe8LzczKWuXtIcRRMc
7u/T/KuVF5MHSRpTgLPSqRt7KKmjQ3ioKuOnXw+dn2SJD5oQUskWxyD+UYeP
ZYBv5fHwjHbn6LEC5pAyHxxXVGfhbvc2dAdXYd1ZZEsMiAtZfvzc3WvFWUOL
pplF9RZM2360W0y+uHOjJf1xjOzfZA6RzB7cmw2+JjGdHRSzixcD5pKxC21J
aH7E0Q38DSv0dzMcZe3fB4ZSii6e0LGtaHi4ZdAklfpIoNm0WZKa0/VF5GlK
832+DeNolTpvc06fOxzAMkkd30yzOATmfb5cb83nCr42QKlG6mSw3nbO2muk
+Qn1v0QZnFy+fS4SnYViei7PRV5FcvhvQrefzOGKAuTS+4kW0c1hqO5Lo7dD
IeeqmxQlpBiPrvmih4BgXqqxmDOKC9S4srdYfZdckVqpdXJpA+ClU25yL8+M
5jVhd3oGFhIhomXHX13Mk/wy+EgGLYBUILSoPWHuGpy1/SfRAOeGjI6Xy5Qu
7FOqbyqx8HVmCwIQXTGEr2HIbCvmeo8szua//T0s1MM0SC2ZszvxufRzqw82
ss/ZsjXeNzHkIDQGPNb4nq0E4Ko88Ialk1YDTjaw1U23pJUUP/kco1qfPj3+
wqDfLaRS0KJN+wC+XAG1GhUtVqTPCuThglCvl78IW5cY1xvZLfPcoNnY+lnt
5gUhipxP1Z1Xd19QUKDR5XH7CkQmLe6MzWHS5QQRiJm05hPqUXj83fItmsG4
bUNmODkH3sC5ERcavBO0q69ErVsNlIx2yZi3n4/10sjh38bxWP3dC6nRDMzz
RAmTIk2O6jnNIwzgwxf4viQ42nxtPsXeP7OGDMfwrjK9vuFaqPjDRfGcDU8u
RmsG3cR3CRSOKEbqsk/JylzfPn3bGL/cjAgDgPneTY+lsrSq9ejmr7MvPWq4
cJUvZtKWJDzCOMifZ1+uoUNTjqGqN2EjI6oaQVRfJ1Fkub6fBJMYfGhYHzQo
5Lc9VtLaepNRdkDCkyMz68bTBJ0T01bhlqST/GwB6CnNLFzjVd+PLrm86gJf
SPFiPXdONhwuQEwbbP7Ik0n/Den0jT2jZWXB5tZ9NntA2oNo15KUCPu1XWu1
E+dhJIQLlw5fdJ1dIdACrftwnXRSw8K/G3+iH5v9VRqhCp7MOEdZslVtdfHu
ssq75z/3rgCGgGHUnd+07POlLW4pqx9VtPvJJuECIY5uD4lgzA8aBKzOFNeF
lMJ9SPjTRQJR8Hgwpdel/0Vj4APBKfLL7qccMqqA/O7CFHfF46gGQNuFsGGC
WT/7nTHf2NNn4IGzjVg0rupxgyh5g0ublnX3L37N/SjVGeLMUUdrlIQ/tcwr
Umv9NkB8r2YOKJlEregEvBMFaOLzh4qbCEIe7kwjBkZIFcmoB+JqsBOT/3a1
cnPp6a3YeJaO/5Cap8zabmwU9RWTFWamdf7n7P4kWq7WUinze10g9Vwxx1Q8
sef+4flKfmLefCbepOn23FdgXWcQCqiJgDIQOiT2idnkFVY7+N586FQcBOKo
dtMjK949G9JgEFTacxqj9XRxMcg2j2ob9F48a9gJDoU8WRwP9xMevBq/PXwR
kp67HV4ElkGPEm9dnb98oQXszvFklHIIhrm2XP8aAoXTTht+eydeTyFW3yni
pCz/IWvRE/ChYMAjsKvyOQs9T9FUFv4qsOJzIBO4tiqNg/q/EUxZQjlNQSFY
32ngvomgcB9pwNpiO/5gcDy16M1URt8H/EzqZG2mr7ZKxQGd9gIQBRybSoM6
dft7pqqzSXsvV96Vo0t0UIBqEfj6wJ5gJHArvgmVUgGtagvIhj4xBb+4sw7b
j3IXbRbkdJM7jP9b12dk3CO5ArKFB4WHskpwnkWjOf3HdZHhyhHUlKm2MuD+
1eG2zHInWUtUZoRpUy3wx4zi9/4fXB0k16rxULZg5/3X/4EbvQ6We8oe8ri/
8jJH0pJeMvTb3mnzzC4BXbBurMBzRsbz/3uNPcgJsuqYi5dLG8HI74vOL1El
Hdlv7w2BO2Agdfe2Hxdxxi8ovg2rKa4A8p3S7bpRvgRlkZklX5TqR0E/mIrw
vRXLFul2nhQbe6yvjtTWyNTlRZ+mZc65tecAShprlAKsMhead5zZr480fzn5
Jbqe8StuPR/M5Kn/ec9Csz3/ZZ2E2vbwxX0gZ6nv+CGB1TCC+abI810TucAn
moBDWKLziLBU1aQGLAnRBgkC3LoTlYGQSNLmkM2zrW+ORlDr5lond1fw5AVJ
jmr2v0X90NEaz2HqKwnUwFnfhBT7HI4lSPPDVX07UQy0DV692w22HvtyV7Bq
Bh8xBNBuqvnWZcA9kjG2UbVsIIvkmxaN0KnYz8S3BRuEghTxwYj4MbJdkJaH
Ll/sXccTW7k6bccE7qaEooHhcob43AVAOdHboIfxx7Im1WWJC2VrGB3xD/Dl
IEEpg5QF1WEcwgIxmmkBlbnGZ9kZNxauu3cqKQ6ccJpZj9zRRhGAjSsB14b4
gGzICBZzoZeC/jwRAh7mPCwJMEDQFme4z1G0fDxJlnxARGbJkQKzKmxZhZMC
YK/p0L28YFAhLiJT3fxxv/jXlEKA/OlYe3ui7E0Xz9rmSGh3scz+Xl9i078/
ZQgP7Baw9yxKq+3Z1Yle/X6O68+OFxXO+kHFSzPbdg4Bv52TreG9TYyB2SgK
rtxiiIFOLba6xZErdwBCAdgpwgQtZnaTIG7i+VRefi5GrfxTTwTkEZ5Vddg3
G5ZJSmptrS5sR3fSeqDczNg6ExMahSc0CInA4eHECiGThUSINK602A43MDiV
A/BV/A1cUyj3I1FkCM8etKr4x17zbwQ/BUpm5CLWF7/3YxKdTbbcf41MPyVG
dJrvWpPAtdGTfUbCxs7DKNNZ3v2uDRprkcDSgxc1+p6B6m9lEM75Te05Sft2
wVskHg5kc/NyyF/F+8dbJ/9tleKYrF0SuWIluzmwFY7wNQ49G52vu0vVXn+a
gFvvfvVCF+zKUxH9qn4u9j9vA6FUc+lCyIcNkSwdlsNBANGHr6A9OHkeXHsA
jhE3vxf+oTSOX/+28bqEU8Wvj6QC70JETupI0StQO6BeDN7PTCUILEe2bHkz
9bECGViasxFwYuPL22sr/lQtyEjyE81/AnIQphuisAcxI9d5PB0wYR5lZV23
CfBsFEim40w6sFBJI+S2cazAqb7fFSXzVPDMthq3K7ZvNVjeIEuwKk4CPMcg
SNt2Y0Yuzlz6xlPwQXE5iTbXG2yW4iBGABDXfH2sfkE5pxBfYuXOsNzXkVJJ
d5hvJiiAOIiigg3A2Enc7vRYl9hDzla4bkJyykozKSE5YCd3A6H+Ap0rIQZR
uXAF4xz1MW5CpKdbCO4IWFaBllS3ISpBv7MbVn45xGQzdqPCal48CprAApTa
f5rpYvGpQ0C6keynFl8kJXhRwkctQcpPa7nfSjXO6oRWp7BdklF/l+eVH2Z4
WZRxjyHrYBkaCSIVe4/JRwPZncIbdXtQJyzxVsVSozF2Itp4PaHEJ3U9mLkq
Bcrlb5XnA0h+4SxztoYC7uU0rBs/BU762bU0/m+cePJPkJRZ+BoGrd2xvnhE
4hJ9N7mDOKvOY/7OcfCmjAafJC77bIPqgam0hHBeqJTyHq4+h45el++G4vW3
RfENg7Se0vHO3pSI5vf6Quke0EeiKWUE/LPq8fAjsDRnSQHNcFpAwYop5M8y
5hZFGIhTYWMVeqehdkqx07vLD0hvm/+ewan3eHC4mBSNRoDAt91OVAKPtn0M
PcmMSqMfPn9sy17coWhZxUMvPrRq0rqRaz+lR2EHXPFWs+AX1LluG5ucv41C
96BgqsRp/vx3ONLe9FNyzzkS66dWI7Prs/qzX1Jp5q2cp4/zV/bNFffA3F5m
2IHJq9eTPCboh4oJSSbEN4880pQiZQ7jL4Wd2giKH7rzes7AhX/snBodBVd6
qhdZFy4y0iqaJDH77TrwVZjyICizsoZU6r8lkkVNrZr6lgM2Np0iiv5+VYDE
6y4U/tUk23NJDUwr4io3tBNNWgdx+nD4kS+HgEP4d4zLcRcL298XlNv/XEbF
AmTASAAXKovWO2nFSjWEJKeRtw8MEzjIDWpeMEKYqSkuo9w+S+nkjWUaNrXh
dtRUUVr/BaA9dFhQBVDFuecIKKSUkJKItH+XOg9z18PH4Q5daIvItfED2wiI
zu8vVUqd4udIMj69ezXak8EJNSi8pb6gyOR9u/G2QhQxiVrxhfEBzQD4za8Z
7OQgl3FE9ViLEjH8LgnMrqlpXp15nsQJBedh+KfbUwUkcCxJva4OTAFhwTo9
08SppFyyePLyqhARWacIsnyVEzWFN99geFjGeepLy2+ESMLHf4BMdW2yzh1i
8TZW/aSGmj5KTz9YQLa6aCZLLhl5DbBHol2J97fc2Emm05xcLvorc4DHamuc
nvrT2olnyoP54ZGSw2FjBDDEcgQSOc13bvIzcU7Z/2JlJVdqecd1ykPZiBws
+O7WzkzUbcNkyvzKk2ZZRJXjbGXZzWCKrX3GzU5XuUnTZAmo9nNWitEggXil
8U5TDZZW4Ga4/BFm4Eqxv0QoPkSL/sbCgLWN+UYt5WQoPMtBAPLRDVdnMnyw
WT/rr5M6XL5khTYAi6YQ7B5p0d9Iv6ADQYl5q0VoUl42XAwbF8pMl5NRLETe
cENMJbtp/hxTjTyw8jVcHE+spjXcXrDhNPvfFOT6x3rMI8HFtemn5SiiB2pt
Qs9aTGz9+02Op7Uu5MjYsVEczVHkKgOAY9GacYb0nS7Km4PNapyUOkMUzlmf
gvwHTfnVVuWXxqdbqru0IsxUNXMjKIU0PfMqXP2ChR0Y1VggoQjqXUuG/q/b
IOvTGnxSf3p/7dJ6nP2+BxZcdPbW8g9CRi8mwrqqI8DNJO3ANWtS1i/EnhKl
W5Orby2NG3VffvvYz2SA4NgyY4d/dAmYVbZTEMuU6p8/rkixew3R5uQLjWlt
dZbl3nVPjX7fPF/goFzpDGubOKYqz8VwTa28zK2KE0HW4hlX07lTffltVtvY
tA9p+YCRJrHHokgcYvifXMGPPkKjnfb4rII1DvZxbxg/QrtUiyyWKa6eaUNL
tmrlY2jd4MRh6Y03Y+81RvjWvGXiIOpBp8epGpOruEytRLF8ZspynSCPKP/5
qUUBf/BlCRkxrFeFTsi/odb9kbOnLCS+qWFTI8Uv63UV0bXp7+VSxBkk0uS0
Ocb5jMEZw4r8sIotFMUICAHbl2eNhKIXCs36i6at1ng3OM2vC+MDnDkC95y9
C0aVUW16HbLImytFY+sYBl3ukkV1HUFQq0c6uB61SHIAGwXVoRGM6IWObheZ
B6jzwqvZ/DPrGR+YFh6oLphDPhsk8vZcXqY0oT44mQxhNrDv5gQ8H7+I+XJW
4JP8gOxt4/YTy0NRhTUcYlxpBVreiB5jdKYbSfoU8M8KLE4SM8vMSqYT01Fu
yjBwDAlAVcCHVjVg7jbwzVhIN49nBhdhRJwgm4B8sni88bbBFQrcosoaFTWe
ZLfa8ZJcw2a+2Sc6EuSRGCMwv7X08KVkVPC76JgjkPY8Y8Qd4VgnxosC7N6N
scbynxKc6ka4VeMxEDR/6vnN1oZsMCbQq0fsl33QkWghKyaFarFtJG+bPf4w
N0tlvnqqHk+WTXoW9vI0i5aW9T3nQL4gu9bVotHP0NPrWjrZpOa+KTIRt7xw
WQjOrW8GChoUD9SfzzIAifdR7j0iTGGHRzIfKw+Ed3ruPWib2kRTjyWwA+WV
3fvma9xnS7HhBS+BLejQWenyhMxy0PN0Stv8DRFBCwSg+K5E5nVdjrPXTMIg
rti5GxAYkfx+ufbEbyG2SVam8RC2ZEJRQUgIPO8UqeJmXdkBR7FFI1SS4ahn
w3QvWJaKm7+FtTx/ou4mHprzEA3MebrxUgysx+suf0ikQ7VKQ9UCMxeLJJez
POulpU547/v04YmX4pcqSo71QplxIlq9Xan94c0r8RixjLGT5/KgZR43q68P
KIAwfHsmAAeBZ6h8EQDfBze7b42hqgOv3fpwdPI/hyez3Qx0D5l9UVg6C+MS
pAOkbO9ssIibP3+W6R/lr1phUAK0rgRFsnAfypCNDJQCacV31Z0sq5W+J/3J
AK04lP25IOhYgPecyuTB06b+zA99gFbXhp1wBhrueIRneVFuVRi7/ua+G+bL
P0tKmpR7/8VQbt2MvltS/NA0oj/Q0xZ2nV+3xJOwVtWdTqHscaDHjcnCmMwQ
5gf5AHigy/lLz3rDGLLdNE3yX+jhhV68Qyq3xJiVttN9podqZLP90zVuDYWB
MDJj3Yk0wWVeKMe4d8p2hloHvcw9Xo18RVwg8gIGpAcGIgN+nkzjIVML+rin
vFMTxxDO7JPJHoqjk4bV7KOr+nI3yqXxrUCZ7ntpKjM4+N+nSyWxbvfBtx4K
uhRQIaGR58DPvL9Z7AadWORi+/e8JjF8BZ4VyYMUCzskPXZnsu4bmO1Np77p
X13UfV5Px6ECvG17X9Xqvc64mlNhAu3weRTcTUJHUJsL+VvwMK+NGD8z63KB
lm4zVkjw0lOCIdk34iM9Grqne7bqOWybmSQkK4LKMciiswZXY7S1ZWuUylNX
xAHj/9NaxtcEj8j7JxdmdXM387v8PQvvIgeGhemdLfArH2YnFOInjKymyaSk
ZQc1nKRMfAoq850xtoyUCVh9XrWUAfMX/q3SVTlUFGOGl28DbIOB+R0E5OjK
50inPYK0wzgbA49OgsJiDTU4F/16kqlKWRRqPi/6/6qkN2lZb6bjrMnO5iJX
RgxFj3ev40H17xWPBH+ZcTh6Nm+9snsxQAYl+xnLr0unVZkt0FeNLlyzrudE
5JhSNkMin5vwCZkNgikROa812ILlERxmOBIYKXvS6U2YNguguH3YdENTIt6p
mKdXPcT1jdSvEkf+A17Y2VEkGqN7gHng5UPmVpLx2jzolsf7grd3LCGxK9uP
ppHv9dJaeAtn5JpTwPENC/2aJIek+JK+wdfSoXvm4ND2kQbXFRznP8cagGQ+
QkvzswEf+BdUxI1yZUAqgjjV0otakKYwUITPeEEellFrD9pyj5nF+4gPi86Z
zHz5F8cSZ1L24rd0z18tB6kUGVZuE90uAL5mHoXwaQACNpmrrWSgSCOy3vpf
MKB3Td8ScJZO8VFGG5toORhob4TmAZntLPqCXkywUhU98wZu1o5IhtbB7ilg
4QqGZJvr+mejBgIUEVyvV7gp9BVXlQAVoy0rAZHOtsri69wt/WZCtd+VsrmR
aJYDADaajcXwAFameyPob61ri8BHFn3mJPRneRBdQEhUsBqL4foSQM/kjRsG
pOuuKPV3ogZtGacaIEO5+oNXK8esw8zwRMtzc9aXWx4+mXHJYNPGTPjXEeA1
I7i90PURvljrJ1OqByepU7hbngSejomf0PkevOd31AqT1qSzgrkJfiuaS2hi
m/LpoOCxsCPdD8mQugHLCJ7swM7Fc46h3zdYqkZmTt9HqnSlE+g6K3IJTliO
uupS1Q86RcQNANxctmSXJqurX4bu3yArYKpfkJAOwDdTbBmKrKnsP/BGSz6J
+qojKwRxmLprcsUP1mYmAGqi2Hu7nncBSaVT+AO8C6T3erwm+50nlZ2xk1eg
waN7il9qgS/3tdKhnb1/cQGO0lrqAhk4B9IbAP9x4HKgkoQVGJOoH2et6I0j
V+Hke0O8Ma11+tua8SXfajsArvHgnpjfN1/7HstfY8Ua9lHiA6SmjZ+EQKZk
AmkYXCcAcdzbBYWRCrbH/rxnkT+CyLQdqxZ3y7EmDAVbGmHE3Ojrwy9+V0bm
Nkohp+PO4sEj8i4pDwHN6j3W0sm4BQFj2BhSHDlKBdflgReLDyZt/Cju6Ta7
jLpMNyVfQQXeikwV0GJhcj3AcAm8K+rB6eyCBMcn72R1rmCu+0GpUrT4kX0R
vdMQksYNEp17ZPnSlb45rofgl9y8Zsu5zlD8fN4qlLfuliTBaeDyAYRrGrg7
jL/v36RdSesX9JHM2GK+kmpmRq6QZW93q0ALihDbDRKl6o7BCnnnJ6RC8q4w
3PgkYHgFV8f6pq/h+/OmzuMtp1wl4f3SzK5guN+mRR5dGJLPTJJlj+pDQzTz
/MQ1OJpo5FSZ2PRKIV2X9UHjA/1DnJSBNMIoZooW4VfjXh/TZINkKzxXoYyw
ckc/FIQ4Gln95s8SSLHwnHxIwo5ITeS42N5rFmKUb+98dXA3WLbRxPrZQ+Vi
7fT0aSjw8xgghftHHbiZps65mEEN4oeeN0vxevq7mlR6JJSKdz39FkUNnCjE
8nKIziAAJcimtIUyf0+HhEdO7jAAs3LOZTSMARlaF2GAKi6I+xKHjQ/7qEem
RpTiXLeNwVKANwI6G13ozWr8Zsx2YZKmU0Ld/FbFggY9V8T451w7HMAuGmwr
cbkbwwOaZdCIY4aEP+0vOddT3z55IFIyOE9l/ysnvuUqXsiWti5/xL37yedr
ZGb3WHhrlMPjBU94hR7bz5s/YgxsqXW/1Li8hj+QtNTWvSn6hMrDwAIcKT+O
IlfwRmF1btiDKKYSkoJj1SEmmBEl5WE9mXrZj9Cz1icrm7bGnENa6BQXJcj7
B58dlgSKtl2bfjcq1Tm1CARbiEr+RfKmUsB+1VX98yvbZBgiWbG+qhSGOY6e
zhbxX32Bx6u9UcKr7nZ84jIYdpNMauU7NL/UJqHXKKxc6/x1sMqqv7UI/SDr
wBNtaeDbZqPVsU/xcN4VgUhFu535ts1rCgMSEEchnvSStZ5Xw5CYx7+yR4a0
QnKSt/NPLUgqfvkBhj5S+/4c50ww3Zre1BTJIqM0NlCHb/F+pC34bHYlRYJN
NOFErWMOeC+JhciCgph1ELzVIuTDrZ6Q16GCR6vwB3sJ7BVxlxO0FI+KQinM
zaQa6wTZUy9Gk64QejB3jySfBGcUd4X69dCWOKnj4eVvSYxXDIyUC4DXh03n
3eJg2JgLL1kxRKCyEHNWu1OqjGUhEfBDW1PEo5PX3/Z4GAgrLsrnoCurV5JR
5tJNL7AWGrtD/Xb65Ng5fiejC9xOFl3WI0pnV0NCZz2JbEy/7w+bCz6n7Q+W
Uk3rEz3UWtWxTJN2YdTUegDlOCK2Iz5IXGBi6jTt5yoRUB3qUfjNYgtuunxy
7L+8wGS20TnJn5q3FvBHX4bPCvj/S1S/htBU+GvbgqE+G4GZd4/eXBN+kp/E
dA/bCoEppAug2LXBRNEN04b5KeXSsEl3u/zE8BxC+hqFJJBK3Mwaw55etC/x
6oAnIfX6/9Iys/KPcd715xT/nVmZeVlETAnkpTBOaFDANc/qHv5n/u6ohtvl
/piql/GE2ElxrrmQO4ZjnZnUhTAzOc5fYZ3yP1TXFEABoZIBrAylj4dlyg2b
GlYCdbfUc+eL16wk8FkXMlFtvRxEOsgbpzebBLUuqPTY22A63fsZZuGy0r9c
0ZFoSFBXJ+9wGmS7Vy+aGb4OgcNJQP4b3lOUyorV5w9sQByOgKiTCSkG75FA
pn2pQ2oXzEAfPjQSPUZe1NxDd3LwLFfy67ejU1gdhEqDlV74yAJ0HHoDj6ZI
4795PawvNz7g+KWE0Pl5qcfhEbAPdpRlPB9D0vfC4VbYWOngQVafKggqlFYN
UgVoMJQnwtaGJCEhKRlBOGEuKEoCojwcbCcdG4NxiXOs/oSyavWa/6v9p6zS
NmVhg69zzb+Ha5jGa1+GFTcI6gYzGQPBUgD1EGE4l3evHSIoa1oKO/iulYMT
hyUXD/kv9TeODP5GNcJiCRkqYTND2yw+iIEgGVuK70MEMuwFYMbXwWyu7bkx
RXiZIbwVknAZPKKEPV/gHl+2NiyEfDasrubDL4A6uMnCYj1KyHVLU7ZdZFz2
8OPGJXFYhFJ6KiJNVNpq9UZA65GxqbjORL6Gj7tYLJwYEXwKft/71tgIljdC
Lk937Y7BvPrPv1hx7A9pdLYYWqk/5kkRJeESg4F3HfGBfpmp+dfluduH+XOi
MSc3shawQ1+sio64Sho4m29FDm2+bipEEvkH0VuSu+kelPI1bcxAio1hekoS
7MhzQdo1fYb4ALgkvnDrrZcjjGG12rPIwW8sPTaRvmwHc8RP6aswcqeR3xmS
4J9FnRP5uIY4Sw83W4dBoWatvbWhKWnXFrTh2rMIwqHUS8s4hBpFgw0O1bHe
02cjgYktMdEB9WnSwrFNTf2RY6+933NItDY4yzFMkJKjv82Arllpil1XeIzZ
G9j0l5iwrLB+diaMqyPoK66IJjXsoV5IPUK8gca1oL7XXXUQL+AgSMnq/AjH
JKvN1JXA8QFWF60JrBHxrflnrYMBXIo19mx3Yelb8SJV3l3BtOMnoZccD7Dm
Urp9E4vvf5uSBugf7Wtoq0awTB8MjUST3PU72hkA8aTR61YbuQG+x4qxH0Tr
k9uVLk3MSx2ykyx4ntwvSg/iIIOakNEOzsLH0obLiAMZtVKKWCdJ0g4CgePa
zGZoW2TfngS3ttYLOuDkf1XLySO8Y1spyAHCOSnuUpoLlKfEKFTEmk3CmN8e
5oWXsLOItrdzXRx5dHBPdtB8qCJdOHCVXH3jm2+j6F+6vABiTMsGS+rk0pBs
BVyTqoNPmwFIKm2KuCT1XF4FClKtSuFA/VH74U9ANe6n9XbxJSIBUnNIKlGA
2abIhcW8XA6Ve5zfdvjO+WlldKuoazFLiwC+U4d8rVkVFDEP7qjAMgZ0P+ls
4yPPnhVkOHotogEo4+lIu7Hth4EMGTWgvpEdqy+31EfSnoD1sUBOtH5st1VV
5R8A/Tq9jhWUO3x2Rbl2AIlXgbSaqJ3j2ubXWtzGYwa16dK3IBIVD3Ws596c
plHJrlqtd2T/Kir1BEhF6eRL7UvWb8GeJ9BkHrlZ0PQsqcx5ThtlbSSRP6xp
CHDqogcHjv9rTihpehDjJ8px0DomwAyDn3VKBXfpLKatUlVad0n1ieb0ArVe
JjKCZbjyxdm8bCKfqSS48H+/rPD0NytHNUjh+yQGkkTTT+RmPvSe7liwODSV
IGNcVnMSrO5e78aDwK58wDIexPqtgbShHy/U+f0sokBArizy1n9AbrPC3iE1
NQ2vDWQwvCj2Byg8abo5fEXshuBIC8Tfp2oTt0O23DA9Ysb9X6DE3BjULBxp
ki8bFyuwe4HiX0FaF9J1IiPcyUAW2BfPk32Hmaa/IJGYsCOvlYUAPkRmtu0F
LJZoJuYfK5IeHPJBWGwSQDv0jPKqFiaPZuICRs8rxfrCZHR0B+TQ1/on71nW
dQhdlDgKGuiyM9OhKDB4ENxIyELwB0DDCNEyKHahM5OMxbcUvRP0bXD6sbQG
j01og3IkJG4RE5gJ/ZqGHaoXjn+aC4Oziu/Mb6IumSMPrHkbaJmJWhz+KGmG
gcVHcn7qgw+JHUhlvCW0wiorcqXLevZ+biveswgXsNocbKtmd7qV+yYEOlRF
3GS2l9UUKlXIrrAQYbxZL3+7QKpWw9xAnIyJz2oQRE+/JTgtv0ItRJvKDeI3
BHBr9ecprO4Gih3XGgH959UpDBZgNmpScXWExEXWEcCQ9g3dWK5ylIIIk4Ud
rW7tBSTNV3ZNU6UQj99X/vFPTAiuwVo2kHe1FajFkU2P05q9PHm8qN9Xokx8
+2shxhffMx8So1Md5oVSOEWoCwrRrJerE2DJH6/3Ytq1vinPEhwGg0FkDiZh
2v0u2kavU8Zvf8ARezum4/bU5Lck2hPfEm7wloSd9u1XoG5ltVt2T+K87BzL
o2XKqHki09BFy4r5iCRpxrrG7JEcGLENbjdwIWUxkTmdum9QQEwl5hfx4q4y
zhZvWauNVPqKM28y2nmCtF6XH+mzdyC9sFdpgJXeC0Dt0hvGf2rfwJ4MUfUM
62SJ+kcd/n2NPfdZZz6MqI1G54nRrYbJxcWAv0a0Myw4D1LYzbQLpFyNWIOR
z95p5Szw04KyLXRFg721LawUGjxn3L6Q1Lngb4QzzImyfwjHU1zwsN6qJPu5
WPN9+Lm4HfhLZeUQ98mYe1xQ+bK4nSaUYPod0WGFeQZ7c1gQ0aXaUYvLP62L
Wqc5fcwFwrhgOzsngmTJFMTPsBEVIG1oR/Sh3VFbc7uybQzIRQMB4eT1Iid8
RX29/MAOi7RMloecu78ymja5IdhBwKGuJxkH2A/+deQqtI5G4xnlRIf+GsZg
yAMpvMkxbL4HrtFDwO65x9+spDpMqbbJj6xHswksdmnE/gsvbNrjlPLuCNHD
e+C4OxcwBDdv1GzdA0haiC9MvlqEQ0E6el8i2vEkkrljxDiQ7LCfZtRetkMU
m4rkKZj3zA1Odjtun8Oeem94ka/6+jvQAonOI1APiVxmV4+po5L2vWjOdEUK
yGfgqK0RyHlzNkkDy68yRRNL1vwRBbYkkVCgUp97gogRib0vee0A4MSZPII3
JvnvB5Kso6Vz4/szNNMvnYEN1D+vszMWJRgNL9gJUjDHZaQGjsonpZD8pIYw
BA9hIpgBbBnzmzH0KZOYDO8UAWuWs1Y5f1w7higCWhY7V4ptivSy3vgu1rZa
2UTxZMRf+bBobNXSzehhJTXE6nw40i5fxuWCpqItc/THsVnKGeR22/6J8168
Zx8ApVprlY/pd/excKmOLCSWMDGHUS9JVv8cSnog88EiI/UKmS5qgltVuEuK
5OWEvt0179h2XtmqGly0cTCfquOW8W8bVJe7E04R+cQHaXsH0FWaKuy3UJPc
znvRGKGJ/zgYY6hdYhTH4fsXCqgNj2/BvVZZmh2esiarBCcDxn9JNU/UI+f2
5z7cakjMGx3FxrAWJ0IGVIkTJMzPa/0yNvpg7QAU4R3X7xA5TV53jdBzFcSM
40v0tX6wInh9XzgpzO/d98UKLNLOeR7rjOP3KszInYEUNY3y4k0vvmki1bwE
TvvJOuhkFNR3n82BbX0qA3bLMXy2syui1kfkiEF7gqDGfW6OI7Xdf4VlOEXJ
unyHvFIVy5tpZoH2K2O2/mJiu8m/j54MI7Y2aOYys/NL0RinKASGhMmE966B
wOI4x9UOZv6qOWXySTEOgV9qlqjozPRrSrueMvGMamnf0fm34RGP3YJt3bjr
PCkxNOPzL78pcEbpet2NR7xqyIoRvc56ioif/9WTv7Lnt0Sbpyav123ngfgk
6kVcGs4D1KTUW0ltN4LMQn24y/h5K1HQXu04GJJegN9TcrQZH217ElXAcW0c
g4B9VG+i49O0lw1NTN9lYYkAiKsvFTMXzq8WAtfwh2wHi83C1FVGT/jARgFx
xd8nr6wj69+lwQKo0oQBTptsRlx1wH54LFgXXJx9sMk8JnvkyTuqUwfg917V
tWeDefWDRcAhGM3OTJfjV4OmJiwq3epKSrFTMT2EAUisFZ6A37Fj02SX+bSb
6SmBZNdx/U9skJzKUZuePT6azJGh3KG6nWKBsci5vXVAOb9m/nMWIWMy1V9O
qxhtpvjHmT1ofipFEqAfgE7WapiVXtrZdABvuDqqKGSscYn3W8qBxWSLGJDz
xcPKMns3xiADFGFJfcuQBYhY0DH5w+eEGc/h2SnsinSfWMcjZOKsTVL1FW2m
z2SvUnQbFL4pKiLjaaEp08SP5CmkwrJ0wwcooj3vIGqSKTZvHxS8uQsICRwJ
wXxKMp65Ka3rf0LJtuJGnKHWRXBK2L0yHqmQAhZYeZtOo8WodVpWKjyeFzxE
xh7zwFnvKsApf+SELH9zcauXij5kq55cPJa41uc4UVg8s1vD8tcM6z8SRWz2
dL9QTCfEdi1M3VqKZF5eMMPDqkuznmnzpWqyKPCHQxTV47jaQYrAYKMpIln5
Oc3dk6igF5vt4uuqR+A0KMrBUDutDEdJ2BQ5vvG9rIAGMYormeXjvpz6cSfG
syW+OsjePZ1c5zvXW7y0JK1eSHgDg/EGuEkaMTl4iGnaHIXG75P2S6iSORuG
7iGDxYr+RSIGe5+l+HzmmnTLOR6hZqRXlKh2RAo3M1LXqvkqNagrMzvEG04M
E2Mdmtkulwv6T5wWRsiOVePGE0ZyyNqY+o8Ru/DovtA+ON1I6OwZMQABNTHx
T/zCbfBSKAgCbIttd8mRxKad8xPEECN1ZQDMqGTzteBOA4R5lxC3Lb7AwOg3
8PfmwbiKpB23Gmd4yUEcnDp6JlGs31Wg1zhVihp+4v9ETqBd9YUSoeHbH3cY
cFizhXUZSP2l7XfHj9Ycw3UbojqSZa0RkpH5224E1oGpCYbKq+VootZRfzFw
U4pYGBqXWYXc/khrL3ODjXploaxFMbRHWk/8EP3ctdmZnt0oQVlHFI/RyI3K
Vgj82byi0u8PDu5Erw7Df30LcwSs1hrAHJTxc7ydAi1aA2Iq3O01wz3ul+TN
jWuVYYEeyH6z/ruFjT4c5qrqFXQZPMj8lFU5/Dz3p7qE/Ut/vfA4Y3rjKPsE
G0lW8BBtraiWst8S+BNh6Nx9lE7bYRmVg3Y8bBPNANL2YR/y0BIWTjMGgnky
SVknWiNeRe1AfIUUaqGt+1U/qEtpMjtbAetOAnrQxs08xr80KPDTYycdzCXy
9IIfmD5tWPLGryaQCkR4VBsiVWxeE3gC0x95/YC08dhjNRTw7jHAhJYE/Vsv
9ddjEnZkeCAF0AMFQMWu0GfIpkW24/E7qmxWeqto3BcDehl2QprkAsMYsIe/
pvXI0GvV+CKZytBO+mQzPDD9Zo3dcFchOljef532zn1S5+VWgU9nduCSADDT
CUZkfI1BSBwlZS6e1mPCMMXR47gHXDQQTHbhHlvME9C0lgyqVq4Rf3qle0pb
p2u+qY+zPoGnfnZ5ysX181r3ZPW1KezT8o/qL6NCeoGFmo/oEgg8AR3+ff/k
k/SL7cJ2CZEuyEatRDNQyqRf9V8ySHOle7LzO6rhcPjL8QeL/bRXnbRV5W33
FBRKeYrzSg8Xr6tG+H1wLtPUI8agviTZSaAwk3mxajbazhxIoWt2Q0LcvJgW
E+Hv8eb7B3cdT6gR06vzzOwtwC8kUQa1TPBeYpK7iRU5nSXACC+O22HfhI7b
JRD6QhjX34YA66amdD79+Vi+gLWHUehpRA7rS6T45fdz0nEFswbciB4t9I4V
uWohek5e0pnfVep8BWxUb6/CAc9miEnwk0AL8sitqd5f2MDKT9Yfp/BL/tAa
c3/lEXyX9NUtspxAoW/Vl0MkJy6xw1xVx83+bfFeuNQjqwEQ2SAn8JJ9I+Ns
wsovv8aY6ZZFGn0LAgjDOi4oUCQw8cOCmEKYd2kmJiM7ntWTdwZA+7+jJzgR
vxPu2nxdf5vO6HShfHP3EWMV85s4EfdANuhofcisTSY5g4SEGiZvSfjLETkC
+bxdYTRqBVEebgxnBROwyrjDFRn4yGt2tUDkhXBuAO6IyhlNZfDyNyWGGOem
h0pzT9AuyvKsXPtUSkgM9SrogNc+cANevjMOHvzWjX5tu8M20YEvibEeRlsa
skOgtCXfAIs1o1yY5NxwR7PrZW0x9vkVn2y6/89n0gL3Oh8jNWfE/+K7iWC9
y8KXBM4sOVR3JHo+7MmTOLAYjlzdilwHko5baBwWzXC24o2w0z1pPpyiTD+7
3LPuhcip5d0bD9SHltKGY6GLEG/L0e4/rWLZLJCMwtcyEpp5YUcrwRs7fCzT
jQXoQdz8CDCu7sGmxFaBcnJ6xmz4Nq2pUYbNv15gLM8xD5aQnhdRFAqRfY6D
x4umSCmBhzj4G7Uo6dy4paZvhmdTa0BxpjteVX3IntiqHspsaomP3FAupS8s
3NzxLkKmlSJ/8bUnTUQ0iDOseFXuBxbHD68RpzsOFB7dDm0tI6aGFnk0Si0n
+3RHxodKjtk/xH+WZtIInhsmrXaddjSVYMY4X6T1FIyIIVUMXucTMO5JTCwl
CL6aBPPUwxrLrSnYP4F3PbjHXGQ41EVIxTi5uZRRv2F1IcudCnUrDjFXEu92
QEBlPoohFaGvWddwl6cZbPeEY4QkKOehuC3aZfX1zDYlgrQhaXYkWmHn4axp
+9GxQQcD1LwFYgZGgu4Dzw8esDOzu1noOgb2/+qWpdwZpwJPDA9FPKFI8THd
UQh5EuG2jQuDEpjPhYIgCw4MYXecypNXdFfVw9+Ielz0lL9Hx2p106C04BZk
POiXQ7nQ10wUlUL1MF9Gh1DyEdUALGPX47bEY/EYFurW4kNWshPCsd5jihzS
EwsM+/haCaLg10F7yr3+vdC/iElp+yQvIPWhIQzzWpBWfpCcZtVU1cbVR1+s
3rLn/JY5fJHHrL6A+fKSWuXyv0PwZVtvIg+owkGVdkdFihzXI+8OhlcXHJVY
P3X3AOH6XFxBPF8e/Tm06rwXlhwGD+3RG46WpVGdOoBe0PqzK0QrE0mjSDGQ
MTbVWEq08kpwqy2/Xn4Azjn1wpvx9xaFU26CZ6D7HoVi0orOsuzgtWlvPcXn
FSO25IMS7bnD1aWSDcI5Z5055o5sIpWcUjDfbcFALLLvVNJmsl0bprZyDRFc
tQy6ZQWutvIeLhDPP1BCdYwj64E7whJRtVePa+okRyO+32gXZN2J8eGu4kz4
MxeucbdHKz2kK3vIa+4d4brGfKlLVaRMbLNAzblTFFCkhElXcY9pd2qEIWwW
+25agMjIT/BFE2ip66THLxtm1SZYBVzYBK9NhxLF6csUM2RWVutdCyvk8Oqs
WP5UaZ6LSPL1K/VcUlyI7CC638oNMs4N1ljyBVa4qloH0LgPOC0OMsDZk73v
srm6WO79Do06sonWIgwPffY9KeAnRfb3pozuCPmPYqGXEyQSleGZFRflz5Tm
hSc6/Gn5dZmQw0/I4cQovkbcrb8olYrZtwWobEP8xNahVWuhwJT1GwHDk8sP
wXq6xs3oXaQaCvPRRStdnLxqhgLt/8K8A8fXzJdD55TG6BIlMd8Yz21ZGhMb
pJe+vg9CZU2fX48rOGO6bwup/UcezKPjUiO3rbqDUIVRQ1hK5ebH6oPKVOwj
kwAZnmMSXS0Zt6DBBgycB8dsNn+73gz6h8mh5ROzw3rBrihBrecvXJw5sl5S
6MMz3rHJrRUPmPOCFl2v1suJuDkKYvQeiSdrxkLrBYt4bH28g9R8McJ9AOYB
D1Q7eLA/OxCi099sWC0Mck6713qxKGdxQthASzVzJ59sI7jawdCGvnVQDoH6
xvbAYsVCedxVBxQsa9Da+RZHVihijGlDJE1VR/FWmgwfoAjck/ZAw3vnqrHC
cJ8CXWJdXyFVlVJNLOf6/9BtJESJV6LItyTaNgTMcIajryRQEhs1met6t7mQ
LjBHSl1vjcffioaLxEg+YIL2SFOLqlVXz3HMKK64skdBpYa+QiyzlbIH6Dr+
f8FgbFl/GyogtMQ28c+r8Gybx4X5n38Hlm9T2F0q6HYTFANkL7VJrEv+8sHK
aoPNtaY0b289vvKPqz+s4sxkAfy0+6gwmEY5+/f4/7IbEkiCb9UDxwbshYZP
wy96xC9mnII1UJTm0rIuM6o9hzWqIabKPI753ld+0bQzcEX7cpO2Oj6JlFUA
rLgaF1snZLPwahVcQumeByYfg9J+FqHKngG0NfiYPF5sgWiPWGqv2CXntBJS
FMlncTHoBIl2Ckoj0ZI4laa4uVERjkSgk3fYQgtxaJF3TzjHuqI0V8LIMRWL
dVTbh02J59a1QZbaOrWW31yoMu3j4HIF1qktSxCA/q51SBLiZEtO8sHwh7/F
qE2f+TrQJcM+b5f00M9n3kwB+tu2EPJTQOkVRDxctYcHgPnFV0uETy6a9OmQ
5z7dd2VG2s7tdSIBmlWgTIZgbfhBzoZNKEjtik618c9qnwLdXUvWwOGoZ1ss
1yptujirUQGnleedD2IwvDxTGZW6YxAFTyVuAABQXWyF45QHjKxhM3faUzCI
OiBAULVaA8rcScfrNnQ1r6UM9fdxHijl/aCKxNI/J3EdTMNCF2oQx43QRvr4
24UonGo6H80DFYaEGxEd3HE8zr+7185ytk155IAtLiS/9JSbwzRvC/JOPawH
rlJF8mMl77mGddShsP0m+bC/lIFdOC48zlPgWdJIntA8lpLhHuXjGHStia4N
XuHpRIkAQkHWV7/iCnr7xm9HnCNYLdC07kr6mIZzEFbf60+sswdYdkTGXERD
RpBt+uzeUhgyKGPYw1MX+ktR+MmmKiiX3W4VyhGzqSvtRDSsMlUfwSEVvC6b
PPDu9t4q2/+86P2Nz38eLucBmV3o7yj6Cg5BFbmUjcbNujz7A4SLsXNAMTfJ
8qqkBtnYkHMOcbiLC+5apxYyGNSV/XUDk2fJo5gsLXWNezKXJxAw7Bsz05s/
0o8Dadon0CM1OyVZz94ReJRwSrKZlLYV+8LTZUqYWHgvu0fEb3SIC1R7mmmv
2pC1Obcd3IZxSYwayOtCyUzXgDYxXvPYo196fnBataoY5ymYv2k0qKrsd1R3
pnXFBIvuTehDDYCVRl9ySmjHEwULrazNd6sFtLplsCT0uY28w6YNAb1FUxxv
P/phk6qJNiStg8rFJuimkOCjN9xovoKENdDINadu1I0vZRE9besFDFaMEBZA
MG9JF+pj6cxmmGjx+UWLqetbJdfB65EzuWJ0/PnPd8V08q8YftFduQ9Nyo6w
CdzH3DVUi670wMX6ENmf90p8den95utHquDMV3h2xkD7sWqM+sAeXfa4/BM7
fh7xY0nRfi0wN/g8aJMbzQVje4QLHDwRjSAF81b3N6O278QdWWrGMJkakJRA
baydtRTxn5crasoecVpmElKxvDDw5NnawJ9YAMxxtswQV/AQJaSSZSPHMf/e
oGQyn/JZxY+x5YAu/vFP/qUmNFcfZtkyyV+/e4paTC1fmfIfNXV8Z8o840xa
0mH/j+276IjMSo7L1L9xib2CHWLRTPO3+ymdyqpaAlRsksuI9AjFhlt7eyYK
2+M5aJFKirrL9h/bsyxXl9ZIkKEEFdDCYP0avbfkdcnf6TZl2wYB11r6a7zH
aEx+MM06Sjv6zGahlmn/8pIjem7XPW8QkCLdCcNQj8nixT/a2BYkwliWOAQ1
IuR9kntlj4sSEwJdhXcObZ9JS5j6idSwBCdoIMhgSJFifS2lxtNtQIf0ogg4
R4sMMr1looLIl3FUG0JT5XS+l2yCPOLHBJOv/6h2Szwj1IW3S47rYteLkPQr
n6Va2MHkTodVBbosA5RwQ+5WOZqD3Hn53o5swAlChG7P+mbL87Ow9js2qWfO
NHDA7wTWCpmwoa3PR42MeN/3If8QfqALRPb6yT7kOk8IsFkebyaBDIJlqDim
yR0RiBj79NwKtV2Gd0LYKGfLAZ8Ax41zVN7YY9YusvUTelCIqkrc40mX0kpN
otUYeQEOBQAALl3Os4Rqy3zmLAf1wuVZE2rH/YDRtdmEpjDwaogfDZAV7PWo
UZAkdjPFvuIPgfTS4uJcFD5c0XVranZFqZcEM+y0HzhOurrvyu1USyDiHiCZ
R4hW7eYzFUQQSnFb6NvHlhNo1JBOVQiXWSQ9A4GQNomRQyIs8WevFDjMRyl8
rP3db35LP/KKWFQfFxjfzaBOcidhGRu2k2KEdXtGb+WU3yEjreZLe4j21SfR
mU6rx5zgRX33skUkZGLogpB2VRLl8KEodfU7GOQp4TsSV5oAvo+LRhto1BVQ
ygXKdOPCzZ136rlPyQ6YPmXCEaytmR2OlGtvv4svEAGDU467pn2VhBYbHbOu
E76GaeMCnoxtXPRxpsoAIRxCkWerddeBMnClg2a87OI9GtgEmPWGGXbj2eSy
J/yK/nGI/Ps0THvpA7rJGyrLBirEQlaKYsG1dACHsFqfI4ja5MNbuZcP03+1
xAL1GrKBsx8meHa1OJUV1WNeqlQpEOsdRNX6yE1phUkUZnqXKtYcVBhgMLhM
wdtIOuVMKgOV5ZNwiYJcx2EWC3nvkLtI+Bn1tbnXqGr6pDwD2JabtfmpUr+C
fFthdBWTdr3YKT5IfnIQDF6hu5DB/GdDozO47SyKDZ2+PrjP+dwMxMhQpfuV
SDrcLHF6E53YGM0VxVy8bfd3D1oJBJm4SWnUYYoc1uy1OGH9SFOQZ6qzpvby
yOeF2AsqFeU1g0oy906Q4DuEfgGSovu0a37HKBlMLX+LKcjHgjHVlHCX72wQ
WU8VwJznT8iDmMitx5PVbr30KkKUdyTHTsinK223AnXq78ge5fjeCm1vMVVW
5C6JQ/YnYH2TlpJYiTgptVeyfo7XrEbeiLk1KsL+hZwNNs0CBmvT8qYJaPDF
GxUAgTKqRiSzjjZSUKNJrCRcAp+BeWepFM+qawfMts+0zRIJVR0gOrnd3PuS
McGUteCCE4gVZ3QxE9u14DCv0CbENbmF2EOunEWnehlfi5oOwphSONwHi3I8
mFjOFmvqOgUrBu1LdjKTmxZctk0LGC0UVYwDH3f/SH+b9MwnAS3txMbs9lyk
8xi7JjdqswoOukPqkeAHcatNOQqI1DOq2bNlgV06VULJ5qLFzjPCZ8HtjcZB
BizlYAJeSe6TZ/7rmnnJxKEbPg7y/FOuarKr7Ul+QqDWvxkXTpc2aywrXHpW
LjpTc7l36b5m099zuorRQlYaeil6ypr0YnnOSNp2HUJGeGUcoebneawMCcrv
W0qIph/qE0Ppma509nbW/mmjlzoLxw5VOU2PehilRk0AJJTLoPj/o98Fq5Ar
Lt2OYpcz9Jg1jRQwsTSGpYGMwLWVqqryCw1XX/XSOQweOlTvxQc6232DLtwu
TT4kIuht8ZwCtjyacOQyNGaMc0fu+G//du6CsueYW6/cQv+elluTL4vNxwVz
IdbRYoRuW9a5wLq3BRHaD+UoAIm99/m49MXwpH1EbnyI3DX0LoBjNiUONR/c
r41qZbQnxKV0fidvM9GlDSj5kUIGeQ8XU7bXGAsP9DdGTfNO09k78OQMcLDy
dLSKHqvDp90FD7u5IjkPYmsLjd62hYSk0Ulvt8wda+/r/D/WrZ1TEYtITYgz
3gwjLCVVezTUnp9JE7Rmte2QGI+oz7KxfHOAX8H+CuaF5PbHthFZgx2piGiH
CHIwH3RROKq9qya7UzLOGnz7yxjqjJ4+kpjWROLObZycXJsjRXOzPlpN3jjl
Iz77/pTxKSawt/1hNcQCOvj/SDZQCfz5tJKNwm1wHWnQyae0kqZwO5Y2Ngl7
3vm0l2uJ8jz07sdsBkzdbWw3T7aLKd0aY6jA6rlDtrit6INu+MeKU+IiXy+Q
YWH8wVQendgHVlQIGAoUnF7aHdc4PiGDUusd5WZsva8ppf+T3PrL0lk5LhyW
6m9lCUTMV95DZtFavFdHACXTIo5Rxim2CBtqhzjCgK6WgbhiHYT+les0/0CX
2kDIlC5gx5DIwCAovz9TQx3u5IfH+22bJKHXC9C93UrKslJzNUlZq1ySe1zm
hiHSECJ/psO52yjafb8YWWjFvZzjGYTPgZ+pu6FcexImYtFKbMo5+/KA4SII
d54pgltIDjz+D3rQY92NIZhbe37wwIs8zPZpbhCT9vrWVdgLHYy7fuCP0eCf
OamZntnjm6NoE+gS0RLrv/+JpzHftjg4iU8OmRcsa9j7n5Z8hJvjXFHxrizx
zOgMk2n0k/bZGU9SS9cpo5+K4Fy3CXT7TrLnOwvmcPF8bl1MkMwViAYGYcU2
k2lAPEqGrLbQe4oYy2w0SdCqz9P4yM/e/YbBNVPbl+slZObTr8xwH8CnEXiU
sq/UdoE08bCZHo8kcM8KmQF+tbYSnzFESgRI5CUyDfW7kUNXSKI5O6xYyYlz
kHVkp0cfyUAArBLM6DTqeg5KXTnm4yj5AZmDWCvyaCJVVAFfwA9VVRhkjuHC
xtLHbzLr0viBAlOFxdzhapovoC83fmc8OVnfSHvODF7k9YYUkq0wuCijl77f
yKUzmiLguX/tCfw+55m8avm42neqbOdMAJrVZy6LYstFS8vYmqwAyVIl78Il
PyfhN9Qw6VcocrKpTCcG1FjhDxSMeiuFhIRGW//A0LQpxD2XonnPedZVRTMj
+kCVyWKk80MJY5DKxAMlX0h0IY6t3HFypYa1CJpk7PFjSQ+bnhfs3GIIjEO2
fyn2RLVoHEd5BwxTV1luQydC1gF+Byy9W5ZANp5b+jpI6wJNWsA3ll2l92WX
xxjjjkENF+ZuUyfDIbMt7Y5rltjVVZpZf+2Ba8xn/baksyynNGYFb5ENrcta
a6C0mEE/GOdQiZ/4nRXTihXi+j8fb7pxEtCKORQ/0WedtXBnljYcDNotGyCu
tAKC5RiKu3HAfmU3RB1IccdXmutoG8P6XogJ/OOXHGSuRhjW4s3ONtLS/+Lu
nkb4JGvo0WQSctug3y8JB4/Hmxs2mVHePXShnxblv4LWYonEzZzbj32ORfCu
VAigNw5k9o7VZyTyODPqLP0zSGSMxFnqGRCEz2+i9vliKsP16OSTRwnCWW0h
rNzH1GFO4zBF7o5kEql3V5VUzLMmZgujhFc8Mcwjjn0pRPy8Yq67HwPVc9+G
G6Iz29A9bJl2J50Mx00hBZtfz7umm1kjqsXol7ZMhqbSYrWSccCGP3zhu1u/
J8roOd6H/rfPCo65i28yysjS0ltJE84/tzKymFKw9aw7Xw9+ekws+LWDOWLu
+DfOaJCQTM3b/R2LF0ZXoGya3BgXSfIckENtW9k4+crLvaSU7OitUPySJsQa
l0ERMcTJ6xyKxMIMItzQGYeqDmW/v1CZ6qyJgY911X4XM96cP0iNycvwtHQR
+RUgUquDvYcMAI+bOyUoOPq1StEq+gB7cZYDVR4cfUpta/JQaWAoAFql8bvL
1PS0bdZ/Jlrr4aISWwfwfr9cJRlL6EABVFSNQjsuP7ylU1xaoaJf/FHWXo0V
zpDXOUlF8tu7Hzzu/J5A3uWWCijVSYgpshgzjQ/q8r68iduU3Q/LWiTSCmV1
ho+nmxId/cnmVPOm36G1+pTGi3q44eFHfxhvbKwUXAt7uRP7SenFR9+kpiC1
245I3g9mKbPLBWzZ2pQ8PaYVbeYTs3W1ZxDwJHBhhzwJk0WYx8Tsw/Z94xSK
hpj2RfVQ+jh8g7doJdxECzM6NUptDPv1mSExHsV37gBsYe1M+5Zcqr0bIvbN
ctVZUdhhDUWofCgEeC2iOGfbkOOsQutottac2nc235ERSkycB4THnlRklmYq
Rr5Xiy6vgemN38IAi3aV5QjulDQ6j20Fe01/fnTIuy50PPyUIl1oz31pI3ZY
dbp5NNRTbRc+iSpopzecr27bxVFahLnk4UQj2/MOqMeIRnbzVKzoV6Art4Pf
mXobctU88ywcLTN2ym34uoO4TIemNGHkN8Gw4r4mslNbzJG6rElpV+TzNbch
V2EWrGxRALA3Cz+wrfgxtRnXxfkDUGDjSNc4GPkL+VKfL3jtFTbWHEkQ2pxV
xw+5nfUmpizoKESEkju0NsZs7y09MFFr2XQHkADed8FfnZURlclieE7bZq7G
AZaLMKB6LeZSFgjEDZQrjTRV9Keg+4PTsPhDdakWg3c7c8Xifh/iMT7Byqra
539tnIXI7aAilqJNE7eei0LayFP9CKTWYhidBiTgm26/YdSZBlWOHvq8MLgo
fZ8m+1y3+j0tn6hI+hlfLmSXws9jhQo6D6yMexK9vz6gEtywXdUwxtaSIM4z
7BSje4UyAkN/kktYC6xPmOI7N9NiicFiK9skFmDRtMQ9tz2EukteIiYEIZK8
jteWi/tvjtY8bJSBfsagHd6LQQDhCW3cyXbBTPpMqGyOS+aGZBmezIbagKrB
HDsRXYcIh0uc7/Lsm1ZNRphC9FeRPjT3m50JmCJUDom7ZwHJNkmRto+sA921
VjqakzSOi/gxik4Gjjj24Zg5oYjqwqZ4TXOwF2MJObki2j1DSQldw73mwcQY
CzZnh4olhU5ja6Qt6D7cx33ltbsvLY8YHeaFWerK69dtSSCMvqEoNopndYiv
QjJY45up8xokmhKr4fOIJu8g6SAqRkBUQ8S9au+WXgwFfBopjuZFNgdXGPNt
GEtnMvyF7sKU+X/6p9xoTgZ5v8DJdB6EKkXBZkzVYeFOdqcpfNdrSaFaqccK
mqTw3jwF4ltMokamZ5lq2ihuZ1Z+GRTEDvtGZgUERnwVZWCklRMkhm8Lk36e
2lIVOGs9Qk7aen1Q4j/Ezp8NRxEZLlAQ/0dRy37JC8qBit1AhIERmj8/UL/Z
BVmVpmBFEehhM8W1lCBQkW9Y7Z5DsIbCzF7Qt9nXkQ3sMd6IxQcvZR9n4MYz
Siw3B+GqsO2LzT6GTKXvba8Go4wLVfpd3ezuK2MjLVpbssc7FhOd8bBuub2v
z5Epp2aa+MaxhKoxETF5pXygANqlfuH/xWXgLekDyJSq0ps+LFI+bxu4KY5Q
D9yXRikMFJGdzHes3w+/WrYB5ZaIg4cH0JRrTxa4en5Q9BAZyLCb278R6sSQ
bKTytEE8MET/o1UgloGj6x+IxzsSEDJBveO7zvU194BbYCK/AvC1IqKqwpj3
5VdsSvewWQiaBugYS0T4m6u68FUmbZEvnxu0SJgi5dh7MANyJkri7i9psaZR
rYrIaVTdpl9O8vD0hJLiHeQ3rLAst2aC07DIcskMmDNKnTcg/jnhamCsVDlP
/qnWKHqw5eB62G7QmmIcPSZMgwx17Z/NizauL88Brzlgf2twLxJHCqzntK4M
5FOkazBthRz0sxJhfRG4EEweKxiqnkf323M+NCKHOI/7EXQzC2KUS/EiIWm2
P4Xxn4IjKLE9zoBQGKD1znsWSRBhRQbI0qMxxF5G3LzBF+XUsKdWMUU5/Sd8
qJ7/uOOUEuJRbSMsJnNW/02EgxfOS8HrsCIQzutI+WHdCl+0T4t9aTPf+fS8
XdvvmCRrwO4sPOXPUkTI9OV0Eop4AMxJisXIehnodmBoz2KHo5n3D0lHQwxK
pZpK5bCW/A0be5RV3Cof89Esnp8rE+7UceXt8yJuekSFj89SCUdhYBc98Npl
8dEncPD8fNHfbcyJFV5S+G6B+m+GZazamWiMC5HvKv8A7IVeRQZuip28B81g
PXTdebUBPkx2hbNefqYAJztF07xhHAu4aILdn5e6EXv7T4nxVR9C9RFbtdI2
C1ptgfekp2UhXvgQ878Ril37a0/yU6ADptZMOrj/T6d6cj9aZMSQUqNbUn85
RmmU/3oMKdhozyMFw7sq3y05Kx4Em0MN8rdWNpW5YLDIgtkJEVRV3lhuduXS
2oIKd14czCLdj1s8id7vkHeYjDgLrB+IyWH1PKeVvee4Zy70kHYrlU70LU03
3pa+ON5a+5H2NkgiK6ecmjyTOIs3UJXrs/vVoNiiBEp1iFaX7A9QklMKW+6r
3iY0hR88/Cl+D0JTsO2wXO01PYRbgoNysq/RUNEiarfBrlkEu1F/Sz6F+8gq
OZBFd2cClDGRViF/7Nw7SI97kPsMFDxKY6GwoJq28E2mI7cflOAtAgozIw7T
Hmbou+bV6v3+rK+zSbPDtnfRjKIAVSeod3hzoWs8jImirFVexDUhlJ+Jh01w
S5xBn4HZNnmHHfsKm0+BmG5tRx6OQk/OFKshG41Vp6Vy4U2PTmuRvFuqz2Pq
6GO7yvPEkK33G5XDfKRPDXHJnq7BNQIAn/PzRWRau85IgdvxdiErBhT/Zu2I
5wBiov9owaBsKnYdbcYJ8AHxFbJU/Q2OJeQwi16LXfghUY91jGawwpx13Yty
0qqwKIv1dp2U4gEphis/8LXtNbRa7j5tXAc+B01F0IdafVxRmabB7kb9e9sW
krgBABHGbnrH3D2FB42m3f6mgOuFVsJYvz7cdZcIsl8/PWD37fW9o7v1kcG5
/brQjnHTvt+IdFcOKKRVp7HZmxJbDuPCuECaZ3/GaF7uVZhiO40LrpHY/nM0
q/t8tu48qXhpSqLrhlf6MfuDcAEIt5AXzJ3iLCkP0Ey2lPz6D/tDiZ/0n8yB
8CGtaEYsMSFPCcjnqCtokzDbQD1CqmqKxL9N/YmIEhm2pwz0XtkLF4EBrdrL
B1jye9mAQQzTmR3Cg2ryyLBJlpCCpjn06gZHyLo7dRv5IrB/QyMSXhCGQY83
6UFjffxFnU5RBLR54+/OUrB7CdIl9uHL1Vx+75p0HjXvsIowl6EklEZCGrY3
290r6T1LNF95IammpyWkZ/qBeG9cizPROpG5oukESBUTIbQYPDIAXbNeKvUJ
kDfI1Dfb4f43hBDUwPJXP2+NChagolOzdJnYJvRxga8uqEm9/44Mhd7u/tZi
ATqcPzzkT6Qv72xRrlFQuuix+J8nkfuB/6BSHI4SzH9MAkuHowGZLLLW1pKk
JqDF61BGyzYMax+KCvY2AN4hnPRrVcwgVebZn0Aq2158vMrqlHE1NlGl8iEQ
GSsAkmPEH/MyytrT97Okx56Su1gl2ZO99ndaYYVedyzuTQh/dmjRlgimv+/9
wsJYFW9OL6j9hcOCiexgYDbH5Zm1JjhZbePWPxc4kXBuVxKMo7ou7rz8uc0C
t4gLu1LxZdXrGU28g5TjO2De3sCKjCjoGtsSGoRrEL4NXzTd67/JKkjEs4Wp
R7AA2Q0KnLDaaOHz0uBa79ydonQkFYSxapBhFvqsS0e8H6z9g7/SWB0Oc8WM
oquoA2puF0Ut0EfAoN1eCZEqY1AtoqBinSxZu8WdZWgHlY9rwL5CmeYOhzM8
/c0wFM/tr5hpdk8eMs53H3ymHSGverBoyNfchptDFND9yjWKlrOF7KBRbO2f
H/ftvrwFceYVavGaEdoKSLwTnHk8dXu8uHxe1NZJt0JaUqnAPHFkbus8exxI
UdypEWgD/tftz+7vHELYr8YiIEVexQTeo0GqC0r/re7YoGmimU8NFEqESUMm
vQby0nkc+hPlMEneP+dOI7u/5IfwE4ihvobYLaDdPZcrpK5F/SPgXX9JxF1d
/pQiY/RUm/5Jh6nld3Se3AqKmrNHCNrsktibT4LA1/prKGEUZf9YQqTs4j/V
LTbGjfDO0OxPBzOusoY/azWHUB/E/Dg4CsVKqZBm1/PrF7PWi1WqzMV4olhM
cCH/m8ItfgZE/dCN/U7bJTr16iVi1aT5GDrHo66uj/WAl8NUf2EHAEkFIixf
skbtDd1JNtXlLFNquuFzEYc35eAg+sVQRe3NVJLUqD2goxX5HpBABMLNu3vv
JgX3vZ8EGI1qoSG1HHnZR2GHr5075/n+rL2eHLJYoS3XFoRP5+/+5c+xi2kY
PBWOlXnr7riSGEmpdQkc5urpN98XXVsTTfAziShdyiIEDB+7Ap+DoDZLRDyI
rSyC0wiY9L3mrOMQcm4is1KSHPpGiFVMahqtOfK2g4S3LktLQc8Nvw9VdkJL
Lg0WCXZ5hJbzCJWfMlhLlKquiNSgpXzfaimN2i31AwqVYqyyDEBgzZGte8Ty
fLKtliKbRcf4hyneTBV8IFSaqzEbPvw2VFDNChnHZuDf40TXoFXXYsILPXH8
53tMV0Dx8vR64ZbatG206EWpVkk3wDOwcQiVorI1w2ZYo00X/s9eA9uTAWNK
SfXydcNP8OZ6/4NhiEpC3j84CImQt1tIdo3cMtKCt9PYlTOkdLEG82C2hCGF
IOeZlBlBmWAX0A2FpGSQD+ryddy8rkJPUIe1Y8JEEjca8RuQTaLA6LenXooz
X+aPr6RwbcV/2inL+7d26TcZDQc7RlMWP3dqr7K+XL6hVOfruibXcCg6sAsY
POofxu+r5QIG1cl3FwEWZ6HYEuHxjYas0EzCEmMR2MtPUeHcq1NfjT6SOT7a
dgxtujGxjrQeyR3FSs8qXZEgaWSUMZqq7Qwsev+YHeKYMHmzExWNbrDNoy+C
Kr5WpxQY6fryXD9qf/V0koEQoO9wQSY+zVYmXF7yc/6lAKzfhAPoq06I/A1K
7FN/Br7T4ijn0bHEWTzT0L57pYyCBfUvJ+OwEi3BTZCubrGKfrxVfPV5c8Vv
ZpLSfYTeN/u9GxaWwv+tCvaw++oSV5SpMCfr0QyxelWfEBtdNrmlU+Y8v3+G
z/bCMtPyMAKCpJIhy/WFgjHMTfUw3M1/MSHsXHAXASp6ODsx/T4HBSq57Q8k
IV9/YQeds424x/ONq3pJ0ofmtx80Giak5DobWORY9Z3r3TAG07UkT91UiYvU
E47Q9yYLaV1SO5Qg+oKoVsEVnfoMCe9fFnttQCTCV6WNMnYitAGYvRJ/yAih
g1MulgKWoobr8C5FOIuyqKfhJPx6L3V0xg2DBUg7/N8Z/inOvKUoN/LC3KMm
GjgkZ72giOyHnxnMyGvV+MyCrdaKr1YUAIPNPqT2rNq51Y6+NQ3THGC5czbE
3Ij9qdRPUylpo96+7ky12z8kchVvey0f25Kb+iGvOnVe9F347ftRlqziAFkm
NA0coS8DxoJNvVVb0Rt07jUkIvC6eLjE65vVS/ZKhzIZMrbbttmc/PCeurfx
XL/0fsuDnqaRx4FQdqcOq3+NgRCAGeoFS/Gf+n2f49ZrPFW/TVjAjzl+BO0x
zsDpwlwUi1ThZf/0WCFkztv6/0CFbcE+ndrP4BxUyBfoKNWQ6K8/i+fUbWNV
4F6YUKc6BqZEIeajTjM16KXPDXBPXNtKy88CEA/cPFH25nhUMGxkvB1ni9Me
d6mSd02qj0cXnGE6Ok66cNOmVW2pYvs6nHbp2gIhGzeZ76TjRiMc0C3bBhg4
EXRcrV8SvrmU/lL21mOENQdwiMZVuVHCSe2o67GhVqcw4qUjsmzIDsTRRA/C
mn8RzU+zYYQwPhe+ULNerAQwpvpkHZVD0Uyd0s3cNjEMSRvkHJwuKLwXhWHq
gFDhFWfLfP/5ILN3InHUgzrtLHVTFclvzK8Mf4Vi9c/OhCwkBSpTap6MaPKc
2yWNDQ7o5RnfU1++m/RjfmiWJtG/LzLlb7NbGy8b1/GEeci6ZJiBZgc1Lu5H
YO6SibtGEd5tPyNeFaOYxQDQa6wJ1D0gWHNHoH3pHi001yvvZAZjtG54cDPy
/gnXzGPcJOTZHbZQXW5yaENU/5414cvpYiZaZ5wFFOOFssQxZat6nIatanxx
NUwcn85wWPzuyqwTrp0P+U78Yeq5B7PNDtViNbVmqGXATz9ovNORBrN3suQG
//DliU72PMBM9xZtK04bj9lfwQYb63PBgjUhoYDa1fc7cZrJIRdw+af+tPvK
s3mPSmC+55hDedkh0//0vFNnO3kjhH4bkJGanQAsSD6lorjReBJ00V1YauxQ
WxZriewaIxQZ+LsWck+pabBKFJwMKwwdE8t4HqtLdILPAosf2FQZsm/6w24N
s9uoQLM8oplqzaAaDilW+d6QANdoOAsP8VK3iU9qELcmr+TnHbLW1iLu1Hst
0aEdPDFGk7J3xZXhapP4cJmvv6awYHeskHytlhLwBM3C0HHPhUoGHrqIWDlw
krTICQ6D/mOB/Iw9Go9YAG1xZ9hWw1xHTDT2n2VzT/LkIEEuwNNaARxYnnhE
VmceJH5jMoP7Cr8NUU8RlQk66p3ekN9zS+0Z18vBNdXsReD1UObdLlGcHepz
le1Ighe9in/wKuhth9tuwIPwfsNdZsJspGZEED/PQbnw4f8iEA+KP3J12LO+
X4f36GRn6JpgsVv0NpgOe2LbVZBrDxdHnPQ4a5vIWwPdDv8stfpDQLK2HuWG
L6QgA4mjlAHOaRI7P00uTHK1UpbUpSpGm0yPmPaiZ8v1ORNQdBBFqDKeP0hA
ZqKSe8obIIypEQ6o8vsYFrI5d53WyEZAfrEA7u2BFyr/pRcbZvT0eja0SsGg
YUKtH8CM2zFYtDwm2IzrI/BeCZ7D5p/EpP0DQgfm4kMFguD58DZuw0xR8ALn
CmaGK+a18bnvoaRKrh9Nl0g46DcskI3jy/BDp0Po5Xq6X9H9KSIXgKChOh4q
i8X0KUg6XMSICrRAqaZQjI13PAFkh3RFdDuvFljb8pXaSbtS0U0A0r3fDQG6
ZrHhTlJkOjXamjdg0hwn/iT+y4b+S/wkdUbokZN2mz2iKjlOfRngQbkupriG
Oo5ovAYbEJaT5dYP9MKM1a3T9ZSOnNkQeUr4uiqDhif/GRCLgQJWMNQedAzT
XrVWs26Uu6G7l6JOFFpRt7qJ0gl7Sag45sdC5MtyRnMcfRdwLCcXf4K9OM9o
/XTC5fLGSbWyv+jIDexYvqmc5QxzyJzwuNOniKw4rcNrilFT1huO2j0tWIHX
apU+yv4h6Pp4H5zEvUCBwAhl9NkuwOAgSjDHdyg3mkOXiuNI/FAdLb1fFBbU
1yM1IH3sCi8OlYkgaujbZimJ6sdxQOYcAuPfC++v6DmNgkFnsowc4LTbxPhb
nfREznVOPba/gZWSkVuHZaKyaYLfkWFjZsjZxJJJCeBX3lICUyMPWOdr3Qnk
4r4goLANsKk7nMRum3lSrrcNj3UW710RSnydJBoOeA2l8T4I4XZiUyENePV8
6bEBDwPRcEXM11TjdLWK9e8AbZ7X5IranTlKKTqAnaK1yuXhLTVUzH3NLI2V
nef7ij3J5i6sqJ9D6pbYMbuWBPofGaunmPQJuvLsct72OP/YZTeXQvkq6gPP
wKxmo8nLCxLdTJB4XWkQLkW9j4XMJ8px7eGKPlZrIZI9IYy59fbz0m2XS4aR
UxYSp+CkHEPocDmdMqHB/Qe4Gom1cHBAudN9nKiDzvpcwFcLsVr+OhQSIGMc
QFvPhWEuV+NaoQMqrkykJP590ahEKejvAb4yY6I7Vf9V92h1D0i/kw0s7LaC
uMFRfOnHkPyMtVYGfobFZ8ciBZAKeiaU5KKEjle7JGdj0Fz6PJFk7AMw/Ubj
3+C4QIZVRBQAK9dshVwRaKJgpUuyLBKE5MfqjjttCC5pmu5JPDvVJZpuDy86
T94BMbO3mpLDg6EGIWI3vBkXg8vgBi1k2CBSXnRPVPuD9iT+n3P1tkeDhpNC
yPIuTUNHxrUSOjO0j8U+zfxg6b3WcbCwbBJcPNY8+GaiSbmYbDSQr1oZZLF1
M9YLNTP46lqlNB/BPy/3ESLBsTE89r86grqeUJSg+MNaUop8h1R8E3RyH/TM
o7XLFXJDNTx9qOlcc/rVlMR7q/3AjN76CvUEJPdwTs5BcumPpifJXtVJv7Gd
OwpQvVJT6hcDrOmlEkarnT/8LjkoBVQfgpUh6KYZkWXtUU2Gmdn/725KQv36
Zgcsb+1+3d77Rgcuf8RtcbwFYFFP8k5poka/GwLoyCDIUDhywi/8uhcD0wSv
qogFNwlV4n9L5rZlsKkBzteEb9UpQpf4nO54spO3hxzUiHZWgbdb4j7DPCI8
VIkBJsGzt6M01J4jXZUwXxWGjPZhZ7p32s5maytRU9wjIeVxa5egiPR7XpZR
l3Hd1w6n61gRCN9Kvu0S6qJOs3g7qNC4L5zQKtEYC+lpmROIld0m2wFpCcey
6iMkCbHWd25CnZvhEAq5enKCRcy+bGsesj90jSdEbR8ywYRhS7EHwlQwHzVN
3v7F+mslVCYasMKQS9iRoarVh+LQgnXVsZwf61pnMNlfKwTBsZkb86oO2icb
xaOGMEOxy5vVKJi92Sj3F5kG7ULTPe/Skfkvl26lxU8fsM3bSwX3qhPV52Xz
Y3gq0DI5yqs626G2Mdk3MnRYd1x7r4Cx6YA0Hzabx/IhwmA+2etz7mOOJ+ad
fgccpBOgA43oXTbSuLx0szZ7hcQlybgS8OPAFqqqFBxALSGGoTG98hKAK2zD
kKbilnUaaQiCUT2LfvKzpN49MMYHLfopcUICqkqPxc+rru/U1yPrhx5w63GA
+R1MnZFa9JgYkF5ia0WrXdKwBL673WSH/ehCbrcsaG1Em6BEsjj2uwr7qn44
M1a+uFAma1IdWXnxmPnpgRgoDV+Gm0IIxxrcAVHDL7LBJHRV/zWQWrQ0aG1G
qQ82IySWb2Ax+GS+/Nx+urQWcdY42j/8vZFvZEm/wBZYgt6quwOL3cia8xVw
WywyH9qyPYWZpMQ28WVVqy5H6xgBG3VrzFBEvVnfZjELt7l4XzWF3S1n6Iir
G1fZy1c4tLKbNEjvfQ6js8ZQgJkYNR/62MzrqtzGoNLlHW0A1x+ndKGHB/Ao
cKMScpZ30ASVqIY0QkYvWBrrLWWGCu4oCoM6wnQ3U5G1zWzdWi5E17QtRO9B
g0/tS9t+XvMp/Nk5ML4uwxSzrFGcRErHnmHXyBL7r1jgT0pRvAGFxHdAzry8
zJK9qsPIoHPFrmM/qeoH7144CpUl/aCBpuyZenBUSfD325j/clsmiy4FEvhJ
Klp8j//TaQd4YTtUM82246DrsGvjEaOtTTuc/15MB+pvZwkv0U2IRMRxSUTF
0dYW/15ST4akKljEtPfYcQa86Zjk2dpiS5qxGEo7xtvT4AZ+PgDZhp2I+bfr
a0cI31RhyfnuO+vAdIPkhd0CizCQmOj7nJLBDuCABH8KyqKbVI6YAj3WayiI
lsbYsDOZmiEqduSK3x3KkudlvNDxXofULNECloEzb1GBviWe8J6CCQtJnQ7V
UzJekGD7Xa1rLZ9DcNvnvRpm4X6UmTGTKdboKvKv+/PUu1f/ZLLZ3xrbZUkB
eltIkF3Zuu94EjvWTVP0f8y/J3V4ucOGuyY3YvePCL0Xx62eCBpBzXFNtxZi
H1KdVPuswA+Ziz9QTdVpK2imngZiF6a7Xg5sALooKHZ3/CqAWL4r2W0DHyK0
lTugp1Ye+q0oCcl/HL8Lwmqaks2qcC+saIw9BRNleh4ggcFyI72wSRrCPXAD
V1h5Q3DtsY5Ez6Eps9tamV5iIDgdAS73wr8iJC2zX8tfSoClZaWUPNfZ1zep
TxfmejaBdJzkefSpbfkUcLiInG40jBZxuyas637qUqpU79g9Wyzfm83eM0jZ
OcpRlNKAFuQOTe5t2vyd5Nsr9M2bWZCD3vVnGyit2DrdydrP57Y8MSOVP4uB
VWG0Lfoh+PubAOF+uqlpJ9t5Hnfdm4g5yZVIALVXf+v2Asazz9+7Xu/Hypfz
BDuxv9112hnmUqsEymK+5z6Bzc5ztlm+RHCF5jqLqUKxno/alraEM6xFKbD5
qVqzcVa+ANCqKv8qwlc8UHo5kwl/Xo48/gXClRPpXONl3xDc6Ee2KWtBB3M+
bU3LAB+0vbBeGnXFAt6EhHsyv/+W2/cfCPnH3qgU0yYWkRRABpLrtuIZ+4x7
bheE7Vv9rNMjrj/3Zg6E3yeb3UfHmOnDcN4TGD6O1mh8LzP7eB9mgcXzDbAk
PEVz9H+WXXrl1Bq2Zl6gkT9tg8jJ7OANugDQ7x3FCmGBgca3KJNQbsDDfWxN
b9DON41WqmSGkFm8mUlJftvcMASvO7udKNM8AYBOARqE7+eSTmO2CO7tMoUN
ifhV1TBAOLJBjlR2/xMCzokLWC0NoZTppUldyOJa3o/EhoOUeU9NckWRiwDT
Br+pgmyIPz4LJ2TTrBHT/7BAXzy7zCHnITLlw7O+5X9KOxU3NU7wg1rUbCmV
9SWiXKcNpAcy8fIThkb4YT+5jrMIVj/pFWQKIVbEZSlkgK3JN7bEeOSospbc
0NsydYyAf4SVK/TfSaOukAGF+OOHpGCO0Bf7r0GDE5nvODX9QaZKxi6IoYly
qqFLQdwoFt93n4z65ebvKZpbbeMb/npC9FisVWx2IhQgVmXOPxe/LtWa/Cx2
EzRrCXYeWO3+TQugyXlFaKr4/CGqviISIwd4zxNc8imlT8XB6SPpMYWKUPAj
Az/8+fkB5aEv4ejb40/L1kwK9egOIzExr5pncsZkIVt+Fqi4VumzubwKEJse
PtbGhi7xADPtjCUbb8tz/zkk6pA4xtE8uKxb7L3WAdj+T2I9s+vzd3nJYd3S
+H3N4CUoSOKnNBVHPmsIaStVAZO0kg3qBPupzP7PpPriCIfd9zx4SBoFenE0
QKAzuRopPvwzxsl6HoOzkmdQPWqhmSrSmlaukLk6n3TyM9vAvecJXiE9xEPL
8fLc43iigBbaa25bgFMorpW3K53tPXP86S5VyONAqnQgcnzz9F2v856D8JzN
0ZcbeW6g/WAH/ah6peD5TLsysN/ecENHns/VbnPddzKCzWQjCiU+YZELZfvZ
50loD1WZORrgrN8V3w5dQwn7yNAujdVk0wmf88XFjg9k4uoiyc7DD9uhQ+5A
O2F2O9sZlr5XQ9K8MjRhoNQea9w9ZxboDC7a4foXc1SQNdEH1IgaQi4EXBq0
Y52ImDwg903KttD4KSCSPEgVIGAU7CMtCSC3VBJb/VG0WQ7Ezh6ZYcHRj+qu
+VrbXqtp5dDqYbqUKK0Z2EGhI0Oevf8U/K4ek86bxPGZUF6YW6qH50RjuJ9c
/RIZydjXZfEZ9XZshfMKTE2jglZLnXgklOiBBzThkoTaXCwzthahviilQleC
xzVMLfQWxgg+pPcZ77PEAQAiwFaj/klaOmctIAt80PaZJ3swCHpqiS+zQmQd
kJgCmWlkpQSe4XtPeVCIXbFL4ZsS1tGpMymM1WNJkGJJM6Bn9HvKgr4Grfcm
hvOmGomPM+VAcaKXcOPbkyh5T7tPNlaVvsIQ1KRmYH4ByOOmxYbkoImDFbzz
ubWQ1njLWsVMluNKQmtH52kV981aojCtvkuJa8+EKAE+0TcJzXStv9YndReX
Fqm9Syg+n3ygK4/cl0EbjQxCXcVUtd1ub/QXMwTWROjqoBMSt78/zMAksoft
a0Fv6hv16mp3NDJF1lyLMlKcXdbpfBWDOFFLH5dcb1HLjLCGW4ehtVHlpE5w
VmqFiJDEVona20fvR89FdTIiWIYnhjmCnLPiLjAfbWdNdygpdohuQwrxSc9H
VFxsUCKx412M3XpHYVLcsiDGmREC8h16KIl1nxyJiuxszS7J+SRBub93j4Lk
wUkbuPxXZvpbZgpGd28s7X3MM1L7Wr7hkGhsimWZO6ws47iWGYFSCcu+3cV4
tMJ0NkuOvP4m0BeYVuw4N2/bueRpBjgG1YPmlPI9EJNyMNPgXQyoSoydu3mE
RmCin3JRs1KPpT02X62qWjZk+E0qRg3w+2ACpkKXMrhtBpIl7/iugWVMA19E
UyjKMKACbkrqOiDcMnFmq6XSykwh5FsQwTgmOLqc9IHCWNttc5GIPFc2AXP6
sQsbiuTCsVbiIkiV3rczOPoBI03C6Ahz3UAzkOSwSuQL36YCwwVCHiS2ah7E
hbJg9Tsrk3mn2xJHXNgUoIAOr2qvMXykF9luViZ8/XvcmcesthIqq/mSwgsV
2lYqQAin9JhIpTYx0TjslyP4qhuuTbaRjWW+ZHjLmwWAmJiSzfZ6HvPT8NPR
PwkR8bpGy9UkOO81d+ChLTXji77aXdFRcit9Hksi7D1QDvM3MXrF2zlpIWIk
61/Zyeeif5MBpEwivvdjXM289wjd2LyvmuyoZodE69gaALWLFKeJC1zTI9vk
yP1QxQsOHmUhUWbgPE9FsZGLgCCcaJw4r2zxsJ1qWO5LTxshw0SeUvbGxYda
mz1CHi6WwSya/fg5O8pE6ZFOj1y1uhYQxcE2m/JGwbNonEmU/TG9nlzTpEW0
sf1qwUnQzLGP79d0IRu1uxA1vx8B0RLsqSQQ3eN/Mp2IDZLz2+ZMA7IkbeY5
mE6WP7QKeXEPJ19e9p0cfwKHWc2iIAxkvVnJQ99p/OvXcvrcrucqIpwxI9uD
FFStQR67mf/EhNdkLUIxEyUzMSH2DLilNz0ZeIsvNCJASWzNqAQOsS7MhQgr
lPMIaMQG7x+5zlCbHqolbypa4KYpU1xXiYmnVswJDg8zC3ifTXrPzZJm6aOT
LMbMJIyZenlYjKyVM4Dx/SJc9roqBxvrlx1MPup9AGWOVbmZLvjpBhabDZuD
ZP5Wlc7DbTSgd2mEW5SepkgsU7Syxvu3Qdc7Np+jZc5HStVBqpI3vKM22PdQ
5+oQ4qNkvvhHzSvcCJgLPe9ufXJt63IoK7hthkkAU/4kWsUHB5C7LILpBN5z
f6YKNNNF6MNN4COkBa0mMcNY3X96ugPOhkDWAaaPb6M2mtHICx+0HwiMPU+p
Za/JGIZt1mPU3UVhqmUSHkHdQFwfV5gN4yuGRB/mXYNQ/3MYXWVKfQf526qJ
zRm5tpzjh4kQPCrEkDsbyEN02kOVlpwzzgUW10PuCwZDEK+55ftsiKajyvqq
qCOprPCO5CEOxrDYmMN7PecGfcCYwQnPXdsTNg5okNvfYJHrP2cnLDtSXP2F
5sZHoGs/UlSyjMMsYkoSZd83cSXEYc+AmAAKERh2QccBn7kU+4eJtnH/sVX/
kvJSYJukJJGOG7RgvYiG2GQbgEv+oLHv68qhZUPVNCQ8stTvRwfS2dn7c4ef
r94nkM/k7gK7S6/1TG4JRvETMAzhLjZpW9m4IYljlroho8Z7XKLwQ7OXcjWi
A+a6v9GOTpBIZumgKdMWSYXLyAYUY6D4vWzYsY38IDJ948127SPXy0ATTDdw
ef8MISWUBtEUkDzYrOsUH9TzQIQlD6JA9fYPWX6/TDy9tRxjz383Spst+MsW
KyYHY3yu7lWhdeBVQgD4invD8VM1uAWI7EQPGb/Xb8honBR5Iys0YzJeXyQL
ox0qPyGVlOhCwOlfgSOr/PFXyp+93Pt8Hdi/T1F9nlkBZ+m+6pGK3Bp3892O
mvY9wsEo/phmbcXRYHS59t/VI1zUFnjLNMYrlgHRaf/+pWCiIobDycrh7XLu
TUQJ+1CShoyydoWQZm52H8pxXpmrZ8CYfuY1WNxvlgOhSbMWnPGDaidFQw6R
koBIgW79abMHb2YYjmLXp4B2GFgQPtJZr1Gfj1Rx94ncoZsOHbijvshQWMgc
U8ZMGp7K4mQyZEiqy4alqDNIsW3zv90Y8eKDb9TKAnTzmAHPIWvijd177H8y
SsxSMIMLbVkmTMwUp5NO4TyiBp0jmv91/lwOirDUGIbz9+16KMb30PSoExc6
SI9ktFRo2oF78n2P+l/gIR8DC+pev3zt3GuyBJ9qvp0q9bSLPK2L1aocOqGg
vgDmD0/JJ04DtPJQjfZl4dZKIFzHFMo75TALpodE/DojD1NHK15v9N+Ywbsq
Cr/H3izCq4TCvERuFsJigT3g8YZVd/v/EOtjv7fQfvi1szDJyIDRBdoajrwL
aFmabtXdrjrnp67icqNs6mmFtmBYRyU2fyJlMNIskgyY5qaByiljyJs0C7yS
RRfuitLR8djIWj147ut0GsXxYBRj4KbyoAt1g3lUEhBZoBr4PuNHfj2X3Vn2
xDLfe8HsWovFhiHgkhtEvTEwDGacdkPEnFB/FUDZwClMHSto+tL96u0U85MR
Stt6pjRAUS87GjbZx0Wxgxbw0yiiDuHAY6FX06CE9MjYuuEoyN480tVFAL7Y
En4YACMY5cBnO1E1qjhwtxQnv1RMTPC1DV8gUonNJJVnhFKG32WzeIbGvZDP
ye+BOEUKarT+Oxb/3Ks7ZXi9KZ7qhJdU/SJxwhLhNiLa6AQqEdPTUGvIuemX
a946yRGOy8FFSwzebJMVxOpYgQc8GcTziW55CUxnYgLrQ7gYKatAXpXyOXRO
nfLk9dMjsl+r9NR643dKIhsk4l8IUM9YDjA5TrU1cfwAZe+EncFsWghOYPd8
hBvnsUPoiVJIkFbnqTKiOaHgJBN3j5RI30BUDqdwmcw9EXidibYFbYgGyMPN
ZB290ldqsqLR8j/KIR0GPTurcUsLwepbwvZPPZgzudxR0sJmF/RMRHODO97y
XryhJuJLJJ5b85Gbc4bTGrRq5vLO9TnA8qqahgrZmFrwYLL/iGDbCLi1pRFT
WhVcOY3u9wYkF2vpm/bGU9RoArvkL2d8uyE5btjN/Iz2ArND3xH6IIjikAAs
BjBkE+M9CuWKSjt/E3iMWUFEW9rRYZkgALdmmeaG1kou6DAmVQ2JOI3pDejM
TbgTHKlq7GpggyWrV/M7yy76fTbB+BfBzcXDaLnHf/ybmhA7SDtNuzC0n9fK
CfK1OfGOeLMij/+hbRKXfaZKTcqjpkWjXBaAPEM5OU3X40/o9fforFT6MahG
R6Kt2IfXFEtvSHiuWrYp0kic21n4p03vt9YcS0t8G9MPVKKAJZgEcFWjskJr
5gFKtundhT5TQWjqERExf5JNbZePp23LMAKky7snlQMTAiRNmNe2uzRvNZXt
UrGznS61wh3KxFBT1/sGwtObArQBEF7rfm+ty5XViFLQXlvPMd9DFydoq7/R
J78FRudIWVG9oxrlpZl4tbmBGE1vKQss+vLQwMH8rpHxkiIOo338dKvPkVEe
5ibA0jtFSRPScnGrW+UQL91Hv86B8gzVG9Sy9YENoYVK4dgvx5c4OeYMUW5c
3mYK8rs+rt3q1UWS9l4UM7YEj60cMy+WteWH8izq/+QAW8FPOO/bw4SoBZMN
SODtc/CO3+PLSgTHvqTSoafWriznRdSmiBl6gEUHOkodkeCvP3QNPNthYLZN
Gq/1bgTvh+5qZOePKth1WGkO6rZqXZP9H/HDITVe1UwmPGbq/31thDWjOpx2
XD6FMUlU9R8onejyCdj86DwP9YfkORA7JhzTsq15CnffcgN3Rl7ksCd058N2
IFyFFmEfSTmVfqvRUfWdjDWc+aeKrhS6UO8XaRFep4LZ/P8YFEa/ijt4sYZ+
uuHQYYxp4Kq/zHoOptRqgttFh1QObCjSJDgoZQMBA7ZsK4F6r/HocFEX77By
wROUIFkliSH7/Cglivyebw5f3q3rvdESGj9spDONhdgoN5G/bNskElTYLsid
LyUa/X+/u3vCA+CNplSkQcjg2868DRY8utTpbH28BPRkWFKfvtxEeH4HA/57
gTMvWONNEJdiHHys6KwHfrcmBv/7bGNgiSTDZ+6P59EGcb7vUB740dxzDGtw
ASHXxFTTJexZLUVeGhkY49qW5FBSpven44z6yh47pkNiOZDDesDBiP+Rgkk7
JbwWVKnXSstzZfFnQGuVYh9Ia31yq+C0eGa+a2OHdXUu7D8BvMKtKO5EbdZ4
icPAP7ylgEFjB4oyR4He+M9yWRmxbe9QUdMeOf+I6Yf4pBdNod0SIedstndM
e/uvS0UZso0SMj/Wt8aOIlyuJKY7IvYzjZ8j8l9eVY3lM2uiwsLmI61g9kQN
d+OyF0xcHY/N1/tbXZ99ZDFef6XYEfCD2JeUb4J12DyDCIkahkgnrEsORZSs
jmqUI5zqN7lpnka9oDDO+aNoIMOK9qLCy78oEobAR3YOD+jpAlgyH3QWq/6a
i/C8xFrO+Qwe8DKwN9MposLRIKKcb6LpNaBjIAMKRTMvBG88tIu52aOznyqr
pLQcXlbiZYul3ZoRz/e8I6WEKDPJ0mCnBTEJO2THVPRXp+YhlErzk9ACUg+F
nLlBDo4beC8aVJl9HTk+cR7QawH7KUdI7Ag7lnEqTmYeSTQUonZwrzIZtQYE
pwi/s/xlLE6FQ/u9SI/SkImWToS1BbaK+6mN4Uc+SzEzk/WBlAzsK4CQMDf1
0yUU1qcA3zQdmdbZR+d0u0SBdhJkgKqpBSwge/k+4txFUSGVFPc6JptF7alu
q+WcXWi/rsch1UY38h0IJHSNa9TAotCVIjAc70mRkkrJjhPB8eA2dQoD6f78
YHjmwGzy3ei1gkMVltuO5PQdeaE4//WX5pFteaS/Lpa42u6PvquP6PbV7OeH
a3SWs9DuzA7GDWULKu/z3aO8Ai6AUuVRpuZ9iXnmBOO28qWkwJzGXBjCUMbE
2KKPhlxsZSwM3mwGfVHFtZm+tJ5Za6woM02bjq/GdhoTzw2DVpNoUvtqlBS2
GQua7CoiOtBxCtDEgnBsyA3p8k/pNeXjPi6wtmjsA8h9SSVEGyv77hnPqAjR
UU/KIADCfpTTpNFm9LmeJEaTyNmMl1B3fU3jqBgKjsQ8RLm/Kvy0iaIR55a6
8nXq30bgpZkyzy/QiBO8Ksp1AAr/wFlcynKiF0p5jjtTrp8XPfGPkF38ppbX
VnnxHhFsoUTzOITSEn5WUcwB36LKFn0F0AyBHw/GBAYiGBYtMZHbhjsDN1rk
YQ2Ipyxb+Ug8dUDqlCvlXjV3NBOYWylWUHnaoBtuvP82/JHGMhvEuYgJ663W
lE4YNOEMfxpeKOTAERh/EwYy2/EGDsg8RcarWZdVPodNxF/illh1Td0iBmMy
mM5KG7QKHDpU4haBbGl6B3aBaPeschBHbmqXsEOeB5x6DlSlyf+nxEhbQBCr
Bq8XDVK1m7RnJQ9eYDzuTMwf9mglKMyrqh/TSICyVnytdpvieGH39OAyXi41
jfmZbH60OFivZ59y4achj9J/ZyLVbZa4UZFkmNKG2o+uO8wEkav1FofGGNQQ
F0FU0ziymM6oi1YOZxMpcy3ip11KSzOGA18nBQqlKlWvTN7S+njuA51jM5rf
qnk1FiU4xZekWbTtq8rA8R+RPUocPCMsf6Uf8/xAcYHjfYfSjqN79cqKbSQV
E8bpakICdDKbU1lPnFlyaELnP+VZWm/DdB69YkvyeEZIHR8EyarA8frtzM5A
KW+1fVY4onoNTvBmXyInYxjqazfysDSe2xL6srIsOzAAWEhAPvyxIVShFvko
CBJ8m9bsjBmfv5IbWhriI6Q2lyoon0B6IY1KdXdrb8T4PfWuz4rmEP4tDRQg
7Lwys7qre7RY+z2EE3uA9MUk5jeCPiXgFJsmhX3U7vF3vLcSCvE2IyHtaNK+
OUUXasTOPHv37Eeb+P62+xV40ifN3/HvmfJHwlbUyPPIg92elTXYdtDzWCuT
5UNnngzxcBY35re9QgKKrk0GNB8MOgl+/Am5dBZnNRJzQsaODus5PcW0fvaD
fVY/Iv84D+FAWa2ALgTv8NVhi/Jr5EvqrewpFJwtZzGm2CEEdEfoKAyS/wbB
NtuMtaOtMUOC5Bfm6L+uhqV8HDYxKSWBHkBZ2IgO22o+DAWJMdk9WSwZXXmD
SXfVcGlq4Blz4AQVrn/eGX5xhqeBfdXRwtzc5jSpdh2PcgKu9hQQ1zir21Ca
IUcp/iRf6yQ6vaHiCOMhCkiEqc7Or0xlQFp6I6bBlumGM+Q7MkDf9mlHg0JI
LN4W2Oobcj//GCjDBYhrBZ+9zdG39AEmWdi7xUIHRwiIaoAXKD0yPYey3kHZ
uf7JitIoSFkO9AR4+VU97cUpPP+VvC5s46zRYCN5S09WVM89akUBrnre8Ei9
Bsx2MngjIRj56mvT3mJfs+FRb+MjvtLI4H4W6Cgrprovua9PLfiSizKtl6sb
GjzWr12IUPRr69NTpxPgv+Z5KVOUurMegKXlsQPWRAXhXKWHYxjIkoaryApi
yuYwcL1hkWhVb1b3YBHfhtlUHmKWdYA8nztaZs5fjvuB3Qxgvg0h1KaVjn5/
xFTFrfHLG/7EAczuQZa3Tv4+HgqVhIm5DgkJu5jgKeF9ympeaiWZSeEc/4nM
VbIMRzyxpvKPd/0573/KZWCHlsH89mBWHjkITnzq2hyZp1pTPw4TdsX9uCRT
o7APuw5QqFuglEvdl75Kt7/iMviBOexqf11PJTwdeLjXl9CLI1K0sfApGPe4
V9pfQyVF2kobidGESAdfRLLORqNQ16WNYGWFkS7MNZCtA0vA0SVxv+Ua9rtq
ooNJC7FzujU0jDRJ3/cADrZU4/ySRPvtiMkJQk5qZphdRyCr08NmzkaGJeJm
+cV5v2gxAybxnUpr1GoJ3842JCkTikwUuZaknkngfSu+2pDhWsLtKs39j3O7
fh0NpXbxj5T8be7DwlnN0dabJy2YFE1SLrEIb8imT5Ete2LXzr/p1Ks5PaTt
YKIsLeKCxkXwmVDC/MOGh90gQzwQbWAjH4wtd54r3lrHAkc+973KUQaN3GmU
Z7y6iv/GT8mxMNHWqHUy4FwPHQRsUmf9aTAP8jD6upvsqLquQGDk0wC0v88M
Y5FAJ+mRMcuTeM6eOXmzQjBYnEWN49+nazuz6TUBc5TNHrQTT5ZZ0lPoXS4Z
7nc1eKe8eHR9O6hKD5C3mB434axE1+9YOfqRtuYtnI199dzEeF8vSolqdfbd
4rV7vnHLyZZGMTakNtoh5g6HNPCmVSPjkacZACpyCtDMl4xyhGMmDWg+pz8Q
f2SrWusjbv5mGKs8ZECIsVvJUK9KZ7gqsEbsrhfII1DS87P5/heVFJKwfKGp
Z9Xg5gVKZFoLzaf7y1xHrB4vX2M2im3lXaKtYeZFtaHbHy04JxYFdwBFD2hi
Ij+PLhlwBmFoZAdFwJ/3NfXDl64q9LCsdBYKn4jQcvXhK1BfnQE8k3JVSPzq
9F6k6LSQ/Z/w8V5QDEEWGtWTpVKmwCjvPdS+4lc/CwKdJSCYtBiTwo3rtkeN
b/iXLouhxI6s6g5hB/xBlLL2RfcHiPu9v0wZLjP+aL3eNN2N/LaRxirstdpv
PCCHMTex1pKGqwNBhMM97ROXRbQj38O3h4MmD/ggG0ClPN+BwkVbmvsXBUfN
TB/Y4CMWa2nbrkHgQkiYGlkWZpnPiXO+WzzKFoey1mjVKjOqKcBvfdBoIJ7f
g/NhlZxmuzJe1m2bWr7YklBDbHCyFHWNMV4DoOt8nIwW4+kIqwYQRIBWcR4v
AQMG6JuTNWi8zQjuqTagRsxXZfouYQ2MuvJzaYAeYodeu8gh79Fg7clJPfQy
aIcNu/ncCBh0aJBWvjU0YC9HAWefRDWlXtHNh9JitLYtVJiK1+sviZVgiL5D
jbiKcL0MfuKSJcMDJUgH8JBRRy5mYMGySrrzmFpZCqBb+yzzzcBC/XuvrSO6
LoJ1JEK8xOHVorUBG8HsJhLbBRsW1+ek1cRSeNE5UzChxPs+q2FuKk7SHhz2
PSFJHxLQP/vs6RHKSKzL31AUNNH8LYCnab5+R0+8e6ZbWknaCq7lU5WSVviV
j90JfOPOT94okn5oYjabWbbf4a+tQllttXxaEWq7YZaBqhb9VOV1rcLMfHZC
9wWM8vNafju8mEzbm1EqK0SGtQd/pMflispUub3jSiMStPK/c+7L2xqQTDw7
f/7Le7L39k6i9aaod01FLN3Dx0uDa7LvOCearWh0e9or/s0cqY5PsHA5cZlV
uiSCo1TyNX+PNGEFaitTTmWBJh3eAN5pkYgUst/hxXUCftP1Jpqh6js1HUsd
GRpOBVVzldiZXr3WUwTAxhYVnxqenOBi1RWFP52rKtbYAT3amx3XEd3kMf6l
JvTlxPNzd9juXHst3MLVTby/FHlK6RfGEx+Gb75SC6KZK7CYJ8jR1XV2XnX+
2VPbXIwn+CesDUZqC3L1oedHnUmP8B48KHkiayUr2jZnulBAGLz2L7dwQhxg
Wpbs5WUFy34EmQ4tvsZbPmUwvjGV0mYMSvhqUtko6+qFCGvifcXbFBl4If4h
q3IBdaTRdy1HduUn3tNJ9HtUA8OeOj+E0Odt16LxZkPC0W0XG5Yc7yzBmT9P
8KR3Yr3plzqofgrZpz86ulRDvE/YEjYDEp+KeRnJ6OrcBY34Je0YndtcE/sM
SrNplPsZd0qmfy8oKmGWVZ6vuOcCAdov8jTEX7NHHOj1WLK/5cluQF4RImqq
nS+sDhPoJtXSEmcR63i/TDuQGlgm2kof73JSQRdZfio2aB39UnoOWL5D1d6+
9gjyyVH9VnCTCkH8BnfDsrC7SUEFulnuql7zSAMARM+t3A5DeMqi+BrR/cTQ
CamrlHQeBunFgk/vAjf40AjFnOL4Q//VRUmiTu8ZUcN7vfxahzKNIK6B+XGY
8WAynKgmu2nobVmtHn6fe83w5dNKYj3Xv7z1JpZyOaRj67vrbb8+oxEE99/l
qpJqYm6r38SjS/nkjcUlqNCq01m2VoX+0SRnGPNireTCWxiZmHeQ/CkRpCNU
juXCkY3lR4JSsabTFwZwvyNWwhZn6/FHdmdc4YfE8cT+IWbFJdrr3LhsO9OI
OsmXV/xy33XQbLr7p3BRooQ1+RCpXHY4B4nBtxdgp1Q7dwPOaJrvfjAnz6la
li5PR7W3NcwVC+iLpdKkjpu/66gezIA4niNHs1UL6Ii0b7NmENVz4sDytjwI
N3tW4tDkYdK9eZ5OF4eZbM/WD4QjPUkguSGcu5UN88zcrb9cuJfy34WI7xko
Nv8FTUYYrijtXTIGOeEIhswjx28qTQ5Ef4gqRpQqHIStVB35NRlBCxzZTgPM
5Dy6v7ihYVMwHLq1DaiB4/ICNPJhFAVtrqF2/4ksLqOXXJbjJdOGda3DOcwM
K5e1sEjQWAJzBI5lImvopEzCOWEWsYO5n5FPs2iSbIJ2TZ28teSf37HO1RiR
FMYR2zSP8U4aLPSTZqb0Fd+/Oo7O6DTNccH1iiHGSg3qgloqrbT1BntCFuQY
XPHMxauKPNtoTvHBnsfWFZgkS1GxhmZ/O9b+IF0BBENfut6E6NdDL2W9pS/L
KC94z2Wf7ARMs/b//jCTmWHy1gf48nL+JgdP8jCPcDl/nz64bs7n5uzNGMdp
OuexWDaL2JOPbiLQxrxkzgYMTglw1SEkl0HEPSzTLeDle8j1JE4cPM+ZBTo2
g/kl+NgQURmSmf2xb+xdT4J89peZogPANoJ9iyfrXmWG5Qhhx/OeQhGBBPH5
Vmj0icsLoBhJNeIU+J5ty7Ugb1PBwpKOdsSV01FnyPi0mM4o+PLhb55li17X
Vt2FYWZEj1ghbaAEhNltpeFwP85BngS4I12qqhrIUhCQNxb6W5CgjXeHKlNj
uayX/HyrvOzvCGPH4A3G8anvJdPf+XHF9scr8kULXC8+dW2JXIlYNGXg3rKj
4jTtZE0GVA4b6ul52JYWwkZ9MSvvDmlk+/niLON30/MMILyq0WajZy2DaR4i
t/BXsbjjtfoQxdLo71AqonSIrnP+wvRvQAJdLn/ByCYl6pqPISQQcWgfbxfQ
psrJZRIDfHKN62jXeK+yQ+S8Edyzz8MR2nrIhKqoxbYGMo1/x4DL/O7HOh+t
aN3qqOIO8Gr/CLVFDbZQKx2W50h38AEB4mWgtKKQGkjGX+vtIbKLqP80vsOj
6x1U46PvaDauKzEW54KcoDoDcraFEjnXZjMNj/TUqsXRLVyJk/rFBgEk4+EP
/QjprLrmHxF2UupYQcPeTpNed9AVDVpOaI6KFOyGKScIwC4PmwnCw3wNGNJS
/sGLCsuSuqDrXFeqQkbVg27GgngZO5X/5h99OcJidbXNDXyhL6K2bZQR3D2Y
BmD9uolKZNmZLC3auiLKRC/tWZdhQN1wMMOctdcuxoVITxeNFeq9s7EpD9RD
16rroWJctDhWEaE8sVEtMB39/3/hYqXL2WD3gGeixyia77q1v6ffL9lsBa8k
qT/1R0aNTl4AVR3ReU9JO2QovgeRwB5CLW3mxyFrNaNFUmyNq94+97IP+ZSo
KjmAD1pfX2zV2QPHp7aTcWrwBQD6CTrtJGeDXzYrV4j8HUy0tM2zycU5UnXg
uJ1hX6Kd9SPhSNbgIJ4pmOpiR5ZeoCypslZ5nS8q/138QL68j3LVC5MthDfe
QihpqYd46EU9NNlaOi9Zl5GdRhPGnEvXSL7TVvhaGTi98bS8ZUzmCBW72Wv2
C4q8sckvRHpJMzHTqqbXfwADLkbN6imHV7qDDsargv5IED//m/82vMP4PL5X
CYGTkx9eN+3sjyD5ASUkcO5iM4svYwa5YkZAkdIAAjlon5vOJAF2cGP058fg
sWN9c9QhR6XVxzK/e7MGRvNxPYoXtQtvicaMrWtB1/01C1kCo5UOE7q/0YLv
ufitv5FgzMw+xJ/xnt/JrE0HoVYtL49uiP+toQrBHfb16KRlu974EuKmET7o
BaBqcnoEr6Bf6FGvWNcLhaQ/kpK9omgIh98nM53FZvxqiIEzvdQx7P6hbmU9
sQEzYju9CuRfkyMREvRhhTyMcyDdJPxhbEemxzli8jH9dstBg95QuHsGQ2c5
x7JxXreAGkFEzFvJGn9zzvFqiePXNAo19g3qxnbH1QuSphA0YXa02jyXpMbQ
h34R5OISX8q9LNFrb+M1rgFHMjp6ThtnfyrVwGLz4G2b/Yxh7p76Wj+AR1hm
r8bMAvQ0B6L3MBW/VA1ibGyDKOriYAVk/sNCYStI1opBv7I2LSQ/mSbbQ9A1
uAA556dMOBWJPKRuRhu3bsAHWm0hWiNbTISTElVZsgQhzOfQCDPMnTum38WS
KakYuPnMfik877mPNnAHY8kqGKYUByIOLSOqbI5KzznK8aDEZzuqf5c5YQ/L
ZbnyBDZtXT4juNTL8P6zXw3vravrDc4zTeHlQKIuq6eTX92e7lNyrUSnfDq0
ReD4dYwYZ4w6yu5xQpvLisxGjWJ6bftW102Q5uacGrwnE8RMATved36Rv0aH
le31IQyiv7B0Lf9RnmAmW+adhs6aRh9LOcJroxdtsUCpVhvZhjBisDPVmzhv
2Rpky2w82tEzC7+wsdRViTK1Dgv4VgrXM8OVd+S5phdPQeHuyoIOql0A62cr
Gy9wr20vW7jhDDi43dx6vcXXj3uiGWQLT95ozg9K5XrMXTXbusR++K3qJguL
Q6lQChHK79fwLpenHufuS035/O5ORHHkMClsCIF88MqaZsbcl3jC12D2XsWg
UQswg7apyWwUcnHSa/2BWH7OkxpdgTaV1BsxPUtu7Z9OB387J75h5dlFijpt
fB6q6pON22GpPaaWtfuoGdc/+TOQ+kuZH7yyoIbKqLRKqgx4iqQqqpCQiSk/
fkfzbup8IAQ6EWkOwm5lvcrzdLU0kmnOAH1pGBVc7W0hvciUhy8Flq21VB+q
1WNwUBpQYnfA7eozK35bwkzSyom/1E3zrnGHqhXNhlilVhQn20YniRlLweiL
4l3BooxBQq7zlsg1P0Lo15WtbQ+UCawbq4kP/vz83hhV6zFziaxYIGFb+RFZ
fzjFQE1mM5gWh1x50JmNqGns2F2bpBl8m0/GvQu0d0E8Cb5f65H7c9WwJGUD
I8oOP8nAS1IkoXIM3ZlYJX0MFGag57SqaWf6bjGO+LDsLXRn9Ek4mE0yHpom
RrDgFCrkMGLqVUwtoYvgtYXTlC4TkkiawKO5Okm/Mz2V+dw9psM7si3VeCcX
lA6xxq4xhDCRXDJa32Jrkx+UXoadTsZKGiw6b8Ud6HdH0WhYMpnV5q2Hgbrw
8iUR0egXz+6AOk5KlkaXfYWH4XOmg+kx88JpB4P0g0RLH7Lw1D+2uHYM9UEB
b7dDyRbEkVQA/kI35eXr7HcSdz9ISM98U521csMHAb8cxtDxzRrf2np/uVme
pkGT+9jJLTMP8i6odwRs7VxRw96xlQepz6JzQ0rZNOfrRyjOFG4UENbCNcHP
mfE3kru/RlhvRaeSqUKr2ds+zDlaXicWb3/mTVl9AALRjsPLUtZi/7pF6ZGt
hdwHqEdpPUM2QrmhXE16Xuaqwk6ec7GD+KnjY9edEEYxfX1sViRCiLkJBNM2
O8G/oGtindQmUVtYAgR0njJ/I1ZiobqVE7+8S1Ycg+o7KGQR2HUh6rg3BOD7
tWwd5eW0zDJXtLEUVw8iDPeCOflQTNQcnCQo3ejcIf8RLJfqgTZPnlpOReku
MI/fS0Dhvid730QPmhVL2iEUy6oFiPIXx+clhv2riteSt+a1Kj1rTiREdoAe
phuyymkor4c5OyDY76dGqVlKtE/onugwQRD7q+qxL6Rmlnq7PWTg0gaucz/T
6rnogu97kF7t2lnosoMWqgvKs1kVThTC+42i7n2fVj5bgitP1wU72XK3i3Zr
/Oq55UjJf4SGPCymUS+lWxCtlgvB0tYA7zfRqXCr/JXdYYLz3OScu+Fh0lgh
BlY35sifrxpsjNoI4wMK3Rp4IXsL8Gzi5mQftZGLFdBdVcVdJ/WdryeDSq7h
0pdx9ors/+v7TO0Ql6EV1SDoaN4FE/3lIOXURSfduGqus/Hb7rRStWQYusdH
zNpIQEqD1RuZlkIWH5IoyqGvwL77FMN4gMHpDqX8NhJfrlsHAzCNV/2Ib2Fp
LxVU+DPIUdex3aRLaf5e8smjvrTvzDPChsfjEgwlS5tOKn3UNHzaZFJ2lB8e
xZwOMzsYNjqlWcpV4DM01AuCiUq/LB5xkvMTNWqFrcWe2/mRI71ynZkzNABW
HAGTwlEZjWXrcgKDe6VODZB4zXMFDWRatMRthuVnKYCFDG29xRLLFOOZ1I+a
LjHS9oNGpbTtMDv7XPa85ZqZJp6YrR7eWvIv1RhZUYVpl4WXJ6Sd6g9NiiHS
M1kEbg9jVD4py+LZ2fD1bJEfCE7xXJ6ifEr5ibJCDWiOLrX3ActU/AhA5tVx
Q+/1RiRkE3eJk37e+owGt+BFV5SO+gqQ6qKcIBSOAOJZPa0PwgKVfVfHthdz
eGnBnFlSBPHOGlO46sWEzeqMJAjEbK34FTn3SfMTdE38w7NNwCFjeR3VyNZM
oLvYY7AL9esyWC7xQivu9+o+NemxvYguwnWUS1020k63581hN5sJbXQ89F6H
jOz3g8EgFOcikNqRnfow43Y55p3cRnmb1i8QGzwgUaEyjVsbZL3qXEDMkI5p
9yoos0mUNQvk4qO1akkjA+XlJpdTuRxC9BvqmDtO1GlgjzgiQXrBPOtH6gWO
WbG6vb5Kv5MaJThKEB0OYLHIKjfPHX/K6Ti7+0gbUfBJpVcZI/7emclkPFmv
TJKZ7eRIfljnbGBLx4OeTxKtaz8lPbSOJxtXgix9WWAbUkCyuKxLSyFmDRbX
NCym5/+2vNVdPqKyGitqEyXZUPhhNlJP8fvecrnKZ15XoB3IFjO7vcwIBdAx
8COpFQi+Ng1sX3CaiKcFep0qWxiMCzzl7zpeNtt1Yv5SDOs1Sx7sccv6IKqA
rzNPnLmoI9qZgywWXShWfN126dHMGuzg0sX9xlp1F4tn5gsPGTanBr6pqD3f
jLvrhgnoRcbL0qgZtqjJO/IdN7lMSOH9YET7HVUptVBq93RHDl9RGSu01az5
6c4/bbOcSvm3PowQqpxQ6blgsFMgV+HUcDohvt7kwNJpk1zIxmj9YSoQV44S
gigBZ5/25rCilsFvOG6q6HODNfSEVrbxuxvVuAahkEtNgiQNWIbUmn4P5uPq
3GGZLlOM5UiN62scliinlmn1vx4qd837FOf8dpF2ONc7HXV/URJ7Uk7QIsTk
MgBkL0Pal6w8pZUs+rovIIGgfgPPpYmJ8XndAqCvG5AsymKellYhafsNIsnK
w7oEGl1d2iltP6qfUzbJA3ifZrY0LqnvVV+51kJIorcoSmRG7S68polkOjap
z8Rhf2CGjR9Up0L3lMCMpxWzWhwnWIUGx54hfW17uzRvCA4d4yytrp0gKMdA
XIV8FLc1QX4bRGEuyYYDXJQCf3UzHjzZtPk77jYs2lmfY2F9komDwCCGPWfQ
IvD5VjP4XBFaC25lm9E+/5Ff3qT415de3rfvBCeJ9f16IN/khyDeHd7h4wpD
RvIrKJKsEhDCue6JbWtULyW5+4lIAd5TFexfUmIm0KZ9TikAvt/k5NRq0nj0
2S8ZZZZSgXrJy9UFTtNteu8dTR4zD83BTlg/hjKbLwM938u0PKlQqv2v+FZI
nxXKQvTwep4G2hlBPCmJuYEmF5u6cyLsoJlUoWNVTN0BjpaM+lS/F4NjQk4r
5473DgoMAUyYlBze5u8WrABRH1K3g5/Ca6Fd+3SGsIqShj9GHrHWN2LBESEl
mnrSs5SfkhqYB9pBfpRu7AaWCH3pVW7TiSjTClt1V1ie3qxQWwFBOPhWtsVa
+6AtLjMEHOByAiDwpuAw0DIIc4DGXsENzF7K+OdgI6I26l3g+VkEZng3SzwD
IU4mQEZII8PAUGAHZH7WbtmUxhFR+glwypCcqcMp/+7+PBl0es+Tz9Mi76lY
UKIJfHRliF4H5yPalrqX9MnofKyoD9rMeC4NjUQKAYN31AOmyO+cVIr0Wt9+
inJXqJjYNOn1JkpsPiYdvEbXOxxepoJ8wxyrw246YLIVGWi1MiP6L+P0VBdF
kcHPl/6PYQ/B3zV179/bhGPExsMz4VuJz4O8gKyce3iXgbPNAY7VaDn4yks3
eAnj5gKh70RWP+nGzvSNiynObZvlXYqe6stVVNX0NV33OcubXvq1tcoPQiTG
zwAIQklI+zCgXRHsaiOYCV2bEp1KiHlOFxxIqPLrdjlCYGzuVcytkX/vCBQw
9WS3HeOZiAvC0o4+tePEOnrq2vIGqNqv3oiCnK5FZ64bZbWVQsFBOjc+YNEF
yIhXiJnd5F4ZqmZyDa7WU86P47thThN6leQW/Ubl/ZQBoDt6q5Ch6aQKMg9z
EAqxEfeUlYadtI3ftoJ2rdNozyZSAOleoP965FcCVbuzZkg3d3yyNFP+Y1fz
rw2382M37lsOe7I0daQTv0f+9sTDu0I6mzYDF/ta5iVKiwJAObqfAJuyp/1w
wU+d9IPFCGO+RpSoA5MaU174Py/mgoOnVa2sbXUAhKcGfmwG8/5AA9pfMaNY
sFzR52zTJ1Y3QRdR8mLP2P2/QTdQAln1j5yJEy8/qmKUQWiwcFARayCfEw1C
QfrIEsKfVb+Ny7+XHBOGN6i9bnM2SpbXbBCMi5Hw051Qaqg7AyzZXOuGvZde
bqZ54aRo9y6NxDNalBEYFZAZ4y/zz4K6CqYrg58G3jjzemsFkt/dIeVcVcfN
aHU1/HPG7Uu5QUiY+FMoibns5EOt69XL8E4NFWb8DO57WZfnVlM7nkd6i5jd
OQ3bkLlGLT6iY5Nsoufr0j+Uh81QP6t1g3Da+XTYFFwxqA4SwCSwZMkbAUnD
sRrEDNJ/LrRH7hMCq2/vQMZBLY37IFKLBDpend/hdLacrY/jhlnkVshKYmJS
G5H5N72xYd7awybnz3sMZzpUzcMqe0p5+3ErCB9Sv2LS55BzgHMab9Lv65U/
1q3Aifevezx22PUn/HlM6Tt5DJN9b2SPhGkmfG0j2HuT/eg7vxRC77+JBRB4
FDGf1LbpSqrnYuvvSQDGEHpH9r6KJK5rN7Z4iFt/ThFNtIfklwEO1ddyg4TF
zy5oWWnfOp3NnYGQ43zMQrJ1cPnnec4bWm6boj/7TcjoLwbvOrtf2mwoOFsx
YqvDMIKnmS1XalkV0fi0cQwsvkBf1RkxEY/DcNOP4Mwtq1xlOelnFsPiyS7j
znmn4BnyhEJ1zFP+eJWBSXwibEi0hG2IpPZ18bnT/Wgiuc1CH5IWekqO5jAc
VJPlMzN7Taqih5lNLmUhNVSeXS7HajzF8E81UG/ggMzfkVKFlFKgkLniTual
S4OygVAnG+Kd57osO+O9jCj4KewPVu506uQ0WbzTUwLr6+cmJZ7wetsNP8GL
gMvJ0m6twUp88E5R9Djmj2UPSLvxXYYhOT9VKi+H6L4+mFtIpGXVMtMgvJNX
Z3F/CHJIHgnaANtEzQorh5UHiiYzEiF6BCEo4D+b9HPOHtRPQRMTkvsKaCNA
wuLnB2ft/yKeRAo4AXNGQIe9mMZJL/z3hvQnbTNcW6MMiVbIJide3gGnU28n
h7fjX51l8G0JgfDaWtUfJpZzyri7hgjZj3437Cbg53kbHWbS02Isarf7blqt
FAKPXVqB9xfapudYgZ6yVmQccwyoQc38BQcZFMJUBunAoy9ifU5c/TMslrBW
xDleh+vwXuIwYnVzdKnP00KBdmp8rcXPSzBPz9dhr1EvbkzcHWrJnSkXKa3S
KT7WmmB629f5Lp5wZaqDA+MN/UARAatZspCbAK3hyWiLACse2K4M5B+p//bi
dORhUZ2/CpsleeJLOj0xp203jQsEz4mGkFPJjY/aTkff+LXWB8wrDhS46HN5
y/Ejb6ZpEwTZTBirnxflEnpV0+sBkhlNEVX9zqLzbHjD/u2BwX+qrhRp6E2F
QitdbEU8dXigHbfeMKxoA914qcdsaYVmnEL4P+SWuWLodpWWx+m5cTWklLH9
D3+zprV3T+/Awh+OtEjlL0Ork7FTkQ2W6e4eIseQXf1OXeGPziY53XXCIcnn
UuguCBZmx07R2Oji1uR3EZ7gHCzg1nCPX3GetmMZbmVwslcD86m3SJB5mjUp
0MSgz0l+58v7PB63pwby/Lw0UJVeTeY+jUSNlUT7YCxt5V5gzGttfX8Gw77g
2zQwPNWlIvmvtjYxgGQF65j/DeHmZKtOjSRlD6EFH91oUr/IvJw5ifQBVsX7
/9NOFhFiIEq834E1NbvOB+yXPMoa33XvZ2oo1Inun5ghTeE0y78zj6qtxX2X
qYjt6t28dN+NVsESgTAIFm6lw3lu+H/SfoFTsSDVfu3/fpZzNlqOt2HsQHbN
Iqiarmj4DkDWnSjtZcEY8EqXPQTTS5Qj0G7eXiitx7K9H9rLVyhFgCv9l7NQ
qm4ZJl+tgMkJTSKx+Y705qTCsNGYo8pEOUQU4XKB9o1pxt7V1Qqq8/8973ps
EoG+m/m6ziJyuhqBr+01qQhi99Jq9ae/TRWeahCAvDbdllsGUMFmuECtQ0JB
2V7W+9lANyRd++jxzLf60BUxdI5CwzmCxV3RLS2ADKsPiNN7waSlzYVQhtyN
0ir4IZkRu2rFsXndoaBSpBAok6RIYsGmUeyuFHWA6VlkZ43S/5Vy/ldW7BHt
hfjRYPqNr2WfRNDkAR3NSE27qgT49oCPFl78SlGFcjAf8cX2kG+S2v+meAqx
q47zCWy+fejIfMxHKKYl+b7cIVPrLigoWVcjTC9fBbGW5+DTHw661jLUKyQY
+ljjltvAhG+OzuYHrvYv9Mm5TCQHTjEx9cG7+pevnnfSINzR7wO8TsLyAIoF
zsrzM5GnB8Pz7dBrgkckabpoPIdvApXDUs9shHYkqohvO2b6t+lqtE61T2p5
OU/dqD4jGvjnD0n16vEBoOROsY1ZccyfYuYnWNW1SP1dOYI7cshQh31FzWi6
HfnzZhvSfBOpGy7DXJudzqJfq+3UjiHE//Bd7gypKVonHfBTvC6TXCTuwNh+
ILxCMwMPvpqQHaCEnD15Tg7iDH+eiZtN0+keBHYLrsEhgeC03rQvH9Lqh8an
gJiWweEzxHdlFZdBYuHTxZxyBlQyq+lnqnsdCcjSL+gfGfWmkfaMJjYmGx0o
uBWkYscP1LY3Rh5tFAs36wPhzc3AYtTHPjCaSAzQyHqhVp94hEi9YFCmFhFP
81EPlyAdBalFU/k4vTiutfU7MMiLh2BGlAiAf7mXrFFb5cebfhLqT2SsQYna
shNKvLh+bc1Z1PBP8ZNy/0fkb6H2uquwXy4Wwxzo0ULY2Z+b1XLlFfdA6Lim
4edHjieUwxQkS/hYDmO/Sj+oOs2ZKYy7YPbcJ2/PKg1NWU+P8ucXX3DBKCW5
ONkVoA5aMidzMy/JRWNqnOSEjn0D16d+I6EygdpLhWPQhm3In6xoZ5sm6qNK
aIklXU743WO+cuauEav6aoPj5PlgSxRRMFhR8pNNyG7hkDFGrtauoAYxOBm+
38yEnAFSvgXftU86QvDaFaZZlOZtL2tjt7lFxg2UcI7YTq5xPDKijzbfPPvZ
BQEFujWTnhdOv99y9JnEHxbcWxkYZAZ6kwQfDPcdto5D0EhsCIPZdzOYdiZM
/6EdMk6rd19G2fZmcb6MeJGaraqDUk3Tc+KA4hTfmBbDA8H865P6cGAo4K77
PvfTM6USXW70WdUt+wrt8VfmYjo2f3Ja/D1n8rvSZ9KTUac/TpPOeLgUcDE/
OIHngzbpPqwey32dTl7XNwBxWIogZ8Q9wRb8fYkkZDBMTJsdPUoN+AV2JeaE
MS2wkoAVkQ5ePM/BgBgKluRf4+QleK48dampA7xe46KhtZW92LKUWpBgjyvk
yaLcR5O5ESJoOr50WFXTqNnfWOPUIGZMQrmq6MHxV+oP6VjDym4XA+2cH71k
D3ilI7+5Gh1einCWFIw6GIzu1Z0kFJwsSNddDrynp3YoYmnPNbZIsKIi5lVa
QD4nGoErFqACgk/vEQLDJZtBLj8vxqb/9657AaXHwsdbjVGxhaaM4w70jinV
7jCoskSa9OYLzjyr58fosR6m43YWpsbDMUiE5yXQ73F8DjXk0e/Li3iYoAXI
kagiE1GRBHoTe31hgTqrybs7DhSF4rszFkmSSRWoX8t3yG1oeXQnM2Bv1Hdo
UcFjoDR9cCwSDVi4uImuIDzOLhGp8apOKD0wSGSbFpWvkwFKjUCJMz0KRsnm
n14tR8GZLRDrxyi9hnS7tDxu5TBGiAV5aUuWXGki+C4Yj94sh/MAHKBdNRGl
sDSBGShccOuYk7/BvlwDp+1MzVKAX0MKhXVv2/tVZFt96Mn7SAvu/J+ztlsl
PWnlTVKp0ZAHEbBX6Cwfp3xaOXUnEoUqabMTnToobFOZ1c0NmokCJ5vaFrnR
+86kDQkH1VO4PB/L/5f9CQR7M9252ZKmGW6XFfwyhCJHsk+n39TUSTa2tcJr
kkrOXc3qm+6lme1yQGhoLOYuzAsgQIxUvLou69pocrMjh5uYqkvTXW1Ikttv
0Py0rusP0u6G3oA5/fqEEXW/TtgJx0PCD1zQpiMchiR1EQ1qoMYczVDov7Xq
dUgfetwepvMaq9707k/CKXxkbBJ6MjYPuorgigfxbo/f9WwW/ne8/U9CCfZs
bpgD2pp6OoiINToht3/tDVeHz3mMu5MFWkuG532WDUSTWG8c3ZMJersR8ewR
ebBZwuJlD4jL0NMV7Rze6mMg721q7linRQXd6t1uf+YxkRX8bSuz7b4N/2aC
vYgLOom5WRJDs4efVZ194j2f0LnrXiKxF+G0wL82zYOahd2h9HYOB7Hz13xR
zxr2uMfgWvMhS0tyK3I+FIIMlxJ5o5tBlQD0Q8TRYTr4R/6FOOeViJDQDKBX
BRT5pIIIWHb6O8rXAM1OeiIrhpxygWa+bd2fLB1+22JrevnjHPwExfh7ZL8p
0MVEkj0UZuwTZ1nUoz7P8vW2Jou850hq4+mWkKpPUkRvqcrjdMAv0pel9J/B
uVtUhN6Ymqtmr1yXJlhrgVt1iHfYsO4+qa27HGKhnjLe31MUxaCkDIFxrVWu
6ia+7yJuZFm/EQQfukWTMrlDUc0jd8WrJZjCbrd9Vkpibe47vTHaSuwhRB6O
yPBhqGpQfmxgd265Z0Qk/dRBbEtYXQTjwbff/Mmi0eqZXFcgZE+/TCDb/jx2
RtSIgGZH0GahM0LEEfIyA5gJn01HR8LkeuCFQzxpfYyiRIakib6ldwV2WirC
XxD6cs6BLmWMx/MMkPB0XPNoUKwEy2B/54zoVHr9eE6TMS4EFRv/+GyJMrri
1ttgRXCwf9eWUQwC8rgcotW+ZNDigcchszJh4nBuYotAUFWJT5rhHwmzJHNb
TyPiUIPPevPEgVxLJxm/NnhQQOKNxJ+SdjhM2u5ZWsHhNEd1nzjfU2mYo+5M
KcTeL1xK7jzGodcM4HvIWi5mjRnrqXgi9A2bT1cAqVx8ApwTrIY4qIy7MALh
3+wcFYc8XeFWhKnS+jhStYkX4S2+F0PqGBPz+5/qidPtveI6JHXi/9LRCbut
iOyHuydHGql2r4GKjcctdCFqdfK/Pw+WKbgmqVCxLq8TO5nlti53QHYBQLcC
Ty9ADneN7I+CxXGg1HnzfAuIarGYYU+0w26Akc+iOaPTgPdlWhGFQpKXB4fG
sFz/ejt1VptG3HkiBr9sp9YPqgXBo+YkrcZXIoiiuc9cfjZZqm9ui6i593rJ
t7GsPld5TAsrtQ7C8Akajg1sPm5kHTUoLODF0XoB/p7Luhplnh+B5T75PuJ1
lCGBvsRP5Qm3tSNma+bfcRaPQ2X9rkC2xHs2gAVOSCtKrtexIwTBEgdoZuvs
md1RBzc9sVQbqWxov0yNPW2noaOj+IFUF4swaiabVNlsiS7J6Tk/hfFIX3gE
1bYRRTLAZWaEJ2oPenBI9kYkbn+gdnXq+og2EdZP6OuX95QX/eRhogK5ttQG
L9lU07jBkkqhlS5T0DdCuE/34sidIVVHE7lDoIIC07/sOoMDEN12CuONgu1U
+R4pjk6sld61UB+Pm3Ez+OzI/6hoDCEpdOrPglGipfecOiHqyOLjqWTED9Xs
QkdZYy4Oglfa1kwqVhKV/jJPrqSN6eqaSmgWlgqXucvIAOy5wdpRxOEluxFU
4gzU1lh0evy5pJNAsziM8mykxoHWEpPGClFhZl0XWLb//fQa2ohYrnvzhEpo
o2havXcojCEqCtWO3lRnpQoVUHX9A23yXqnZyTPZw0oZsdxbSNjJfxTW/wRL
3PKrtJ73xASXZfFNTe6DLlDogCVKNzNkXAaubUry0EMTJzYeFh+hruAbPaGA
AkdcfHMYbzC0iFBv6ILN0fn9SRUDyuKB84YxvHoY/KKnufR/YVhRct5aanz6
Lqi35eANSmQipOdjeB7ocaiEXYwbh7OZQk/3nzm+AuzYnWKmpAmS0ydfiNU6
3jZWAvL4uydhUS7xXTWLsPObeugRNuCws7OkqZGoR51PNVylSiLzJfryBScF
EyV5/Z1+9scs3XCNHEYEf+cEcaLRBryOzWRpYL0yLqAPtMusWVXB0DnhDsa+
jq7+Q+RLcfkKoBQrbiosPMe8GzmGq/DOY+sluAPiXi5wTHzdPYIAJWW2Tjsx
Qe69ebob2Eq9Iuaw+CWY6tqtCKrMvUlS3713/2zdom1+sEv4Rr/1KiA49RPq
eu5zQjKZNHH5A9vHikQt5YlFUa/KElvL4KwisUaZbvl2x4YR7NQGIT/GVRt1
cwfLcaD+LnkKVQ/NTsoj38m560PltS8OrtsX46Z4TwP4Gpv/UhDiw3RnoQ5U
0/2cGX3TdwWmiwPL3wDXjuVtG2/L+dMhQGynsXz4q/w31Il2hg08STMfLt47
ontngkBNBIYJJStczX5sYP8WtAcU0g2Mi4Yca4qkuQmAmy/RxntuIvobf20k
6/wc4zHxLx6727ngRbsScSBpwbN5ZKqJhEGa3U4zjfj5W5E3uy/dhiPIBEDn
LuRwNadviPkv5eMKSQrmA7vnWVn1hEW2FlL+gntXn1YPkDlefTqn0v1veIJy
UrN1oheHQhfyRjSp41HdqpLpC0LTNkaKFHBiK4cuxB44kgkiAvUX0F5yzOm9
h6YK6YwiasyFN6a5GDmWNbj2u1XB1+3lSA41sBTWgQKXU92wB9DNiKQqkoyk
TWbmJrIQ69qV6lMxm5ROcVV1McBSHDOfcjAum1RsYOlrcMnHGLrQoHiXCuBi
6eIj6X4VlzKJWkBk1cAffBEvE7wzyTXjb0FtvBA2O4iEteBRMcLnWjgpcKv8
GJwW7miZjJPFOHNu6TVSHLvVnkH+Tgx9YQa1lRqBXW+cERnd3b80Q+UxbB6r
zEnahOgnwieLT5Ntvb9t2UkLp7I5J2VSmIpwJ2hn576hUsiV4Wj1Ez77tO0V
lO6asUZBCUBOT3USNsFjZ6/E/IWeelhx/bxzZ9L0sJ6W6PhK4zyuPv32isiu
YpWRp2bU2HAwK/Y7BbdyFfxNWM641QoCSxteij3lSsuy/H/04lIgaj/koqz0
P3Giq7n7qhGV0bFPiuH9gtYczSUjuwZ1y4HUQtUFw/76cAw9QkR8bOGh2lJR
aYeHpPnasNw2Q67LopazlKzpn+bfNdbb6Zgi2T+dKOvsgvOKvaaZUE3D7fw4
Vlryx1Te+PNkD+7hABD/Q8QxNb3AmJl3jqg37byHJhb6velKecCJRMR0FdKd
d4Ihq9MemyNYCje1yK+TZE9v9d1g5l65GGR32TIfGj31czUmEiJFpGBMVAcn
Vpbqg/NykiADdW2VxLrwURtAZY9qchMIi3D408nuShxE4rZwjh+HkDuoYFGI
/XcovJPb84n50xxAEo1/bfzqmPcx4yJdUfEHHut377YGMqWj/0KSK2sBsIwv
bYfUbHP8oQ6/1Pq9VMNfRuHmgoF5FtYvMZkBeABKQnnpNCQTCXLxOZ24waav
dRTNMDblQobxnn+EDuSYPW+8VsQeZEyotoVUn1w+lQ/ANivZic7PYMnRVOMy
rGfY0LSYIk9ybj2fbub2b35QPScYdKUcnh4vmhmiw7d+l1oAXFVwOzrTZvua
CkGZvt/dZ+Xjr3wZz2JjSDXfs0A0Xq6oCObkwrhdY5bVY3h0ZML2Hf0rq1PC
852UJBYAS6DUEc6S6eMW9XN3OSliN0friBUgD5QGF2PJoIOACpG4RqX1ZzvN
+u1JOb+G5gPC6rJxO9cNUHJrREHA2tLE+EQem5xibjijX/Ks7oMwCEHeaJOL
Kjs1RfF33jL0jh8oAtUnirN8HEmt0N8k/9sl551eoZLZFF8C4eIRqmybIiMx
NkvjqYJzi5c0QTzRnE3y9FtJxZJI8VZ8sy34ECX2l6ETZYr3W3odRdoEKKph
A+Mwp+Thwde2D9VlkLlrnG3EuUvTLxTV/7uT7J1TMj8GOorabF7snqd72IO8
zVWuL4IQgzoRoBs0CcK/+koee0RQ33+P78pxGUwwBoPaiijpds8v04dbHxQJ
gy98Ih1SfvAHNoxqhNI6JpNSzqXsLrVnu83B8wxa11Hbg/QrhiKf/5Pk71En
EJWWefURzkIXBK8H+lO0LHud1mMqMA237R1585OpgcYpRWcwjTgF2UxP9w9s
Rw0aVdUNtoZFfWIHxfzT3k+lJGg2Tue0xB+/7b5DrHWhyGYz16Ju5VWHgZp7
pQKQSpBWosiN6CiFHGyDDSTuIMjFgfL+zNtbWUFozTRPUunamYsbznSl2xnm
BI0erSgUdGpP7gpisy7hZYOKQj+1sNKn2liDn+Vi6kQAM6jt2FMajuQFhu7R
oGULWMx/AawOTKP5U7kyHYWRgiYQbMYvwM6DxgrgdlfJV67buUefac/CWWg5
YcwL3gTekYRFy8pcECkKCu5a+xt9bOWVgEoX2V6Ce2jsrDzgMeESCKHyGpAr
wYWZo6sdJgGVcjKW2WO6zs5/kxUEym2p30PuS7C3oEGEGc3h2qpQnvICqdbz
SQSy7WYMbpo4keVuAExa4lz+BrHWilKd6OaqSzpfLLX8e40yKA924dqXCDtV
97aKFZoSaIDrbRiwBfOTI6mw0O8sAlVmCgSMYbEbZZyNXvZcBd2IegkA33VA
0Im933J5/FrIZh3vew3UyH+BTBWjAAjBSCsLXUwrWEA5SXiWU7hTYTumyHDC
G172P/nfwXYuMYcO+WWHD/OtYA65vwhMRrTtvGUpntGV0UMz9AwX79RiuE1c
c8YVKLe7qDYkbahjKm1iI/Oen8/1gAyBHecTE9HTMvu9M7Y+/6bODYR4aKHw
R5WLl50aRmdH49AfjRqrzAh0XKwFpBhyRTR+8FTAlLHpw/Jfp60ZFVgmgz57
EvwhveEQFMcyb279Xk3ANCzT5WYF0xTPFT6cfpORTPbQf4FGwQSpFNCTqJrO
vUEFbDC7/9CIpVY+HpdGiCU6vyprdWbxOfqK2aNvrM6ACUi15mW6wGvh7CrR
b2ilDzoRA2T7WHJaMZya0UnGIRAhQEDYV7wypAOiCAfyirLepD4o92nTsVRA
leTftjvmp2WBB73i00WTJmI8TZ6dCbZQSq0oZ0HUgNfvcyJqu1dp/2Mrr00M
vtrGy3inKQWB2JQLJQbL6FAWtO9lDnjfdNXQHlxFy0ZzTZRuGfprjGNXIyaV
3LOCTw/SgLiz2SdMmsov2IDJMBnM+PJjA0KX5NaOVQ2eIl+dhRVsXaziE4y+
j2dPHJ0/rhiodAK3Md7D/ChvuSAjpCMhpmwh+ylAOoIGtP8F2XryGZBFfqxD
RbjXdul6gLt0GUDOZfIgfBvZVnpZyf6U5VZFH2hEYAx+yLgSxC8AGUCkDmiq
qvTNCu1FFUOy1Y2JLZmVfhyWPSb0hyyGXt+uvgrvRyVP1b5iEWON5IjLU+3h
mLacnhgOrA4Z3AHj2pB5VIfehHiQirWOLrrYoIO6om2ZmOk/h5YfESeC8tDQ
h0nqDvc7NUq178B2zTxtrPWDsme+MCqEc+4Kyd0F+fLYpU+3dmvNXNYqGPsi
IjT5fmS55MwKYPU+XKpWszz0kKlnVFowQ6ExjdbYAKjam2OJxkt03YU/tarS
Ed6qfOZGwtqLhGZziaIqWq+EJSZ3wt5LnUloAiZrU/WRuOiS0DND4e08SQpk
/EZ5TymAHWAMqb4gaC31hoQieG77mdhO1ZkiJ5+WMoPvEeoS30Dv0NB3sD72
zoxVS7439U2BOB+rMxHWGXuXLv4PWVtdPbAucGAnZAvS4fOZeJ/4eiFlhVeL
USJn21xoU/TGPD3PLdk34YwNFH/p0ryXidEIkiaB9S2INbeLYfA22ZL+pQ+n
95+/XL9cSr4v3WjNq9Jp3glBx4eaJNNIH/J7FJYmd3fV5csuY4NQOUFD/+bE
T5tbRgZalT4Q2reyK3F9EXipywNeCTDOyfI5YOgt6FGI5eNlC8QTIHu+8Z65
AesWwbQCWUxI3BICNRCW75WOnMFwwD0TX04ukPTyTwCnPDiAqBtSowiU7n18
JChzcjaqNJZOeVScRX/wIXz3hop0KAc4VNhvQcIxv0H7P1ZbQmMY+nS4lezE
CxqFSG42Xm3fMEK0JQqjsL8yeO+AjYeEJG0O9GIFn5oCFdWz5rciEcaR8FoQ
viHLcJYIovhSa0s8aNczuIedOJLy5uRedXqlI+Z38mOk0g43ds3b8XCSxOZZ
tO9hOesiSX0mWkCSzHW0EnbPtpYHeZhL9HHXSnzhMIi4wtJi+/twK19x/U9q
3bArykwJFT6GCJJT8TiA8UEhQh0yG1vPZ6utEBm6hXyEwr1nYF8yhNY49BGv
FhInIfP9cTHh1QwMsBW23E58lyHShAp26XJH0ei4fqn/XF/lgzMNczK3RQx3
kmIgWrqMGg3KMT+e7OqrTvJaEGS5tmYH/EJoEqhhokWDNVwGM9bIVtsbhqko
dXKzUX0OcVBhk5j1rvfvvwNEomYvkrN8HEi5HzT4UfIXvVlc6Mz8PIgVLpmY
TNQzsUSSVNXa86a3nXTdT2agmotwvgvhSil7W32S8OkbTzGXV68593zGdfxJ
+NxiiREXI/5kDgkRCSQP/236c57k4Q6g3FMHvHfqCpLQoaks6UNu/2psEz9I
FhHWLps7hXrYGo8ua9ZjbjCBOXPLOYjqg/pl7zfdee6DSg+yMnqW/OKOJkad
Sz5i6oT/j2ixO1jEkEVMZbKufmvFYhjAbQ8VSgt0MVd//JhiX/qGUFI7igA+
BpQzEFPG597YmgqtQfi0mvVmbUqtwsbcxmOmIW/pNPuziQnssXZcB+pMzP4y
MsPEqpFi/BdWxsD+ks6rCbkyWxxer0bmdgCC9mYlRBukRtPRqprRtVT1+GMA
clqXJrRmw/Ldo5a+Hhzszjp7KQtU9u075DWjzHGK/qO08RCAZ0W+DnjpECTZ
ul6+VQCdv/FRxiJfAJflmNdNZkd0UFPAHIzl4YTVhUFvF18aVz//xOKYq4H7
Ww5tJmyR3gBC7GMDsI7Np9gcR2MPLZpBhYFLiXQWjneExf5eDRVuUdAjnwL6
TSiqqHPAHf6lSQoGxgUyV5dHiXh7mQT+3wHKomqLcrJx8li6G2+90ozOyNkK
LhpWR/fpE7uGmUjLqCW1lot1Y2TDABDw9T1NIg9dVDiFPca7+WlvPhnhXei9
YTpXSCWYsfP/gTp2kAyk5wpFYMyRcclbW7L914Z8HyAGuTAlRFVhpeW/CBOK
z6KyRHxmk9mUOBmvkMnY6VLgSjiojpPtuvdskJmEp6gOeS7foXcnkwsutMyn
wvlSQ3l/Vaqi+lWSWJ/7Kh0xRsDT7a2+4SCVUFrG09EsieK5pwKBxUq+rv7j
bpzEGg2MGUmtGwD+VtKSlZ9iEjWbngiHid6P/YP8HpG5NQFk1EnY1/qktqCw
UacJ2N7/hOsp9MasF1AHQQQ1DWKAOnfS5lAI9dglhycixh6KdICDI1wVoudj
swp7020DmtS0MJp9wXCBfvM0ycrdYHeo1JyJoIN0WQIYI8nG0cJ4T9A2OY6t
D/hdzISP+qa7D/wQ6/LJV0pXdiL7l+0fthC0WEcuClzX/E9pqEjoX+4Vs+Q+
fxhrLShJTQ6BjvI5MeLIgXBRhSsXtg0VlRb/KkaG9koQyw1oiqYnytQo7O6c
m4KyDayc63Zz0BlW73+wikOV9fbbJ47nZENHYGsNuPh6cylaeK8vodDBVaTS
cSe+h4WNZU7XEq1Ur/1YoAZcMLefsWweyNOMsdVe1fh98qW1wQ89D3N/YICS
F9UA+bEZCBK0A1BX4vVTES9xWMvqAKY3nbFg+R9isWQkrSOuKl+iYXc2iTl6
pw6x8VzZwdcqLUt1CpvL2461cxiGiWbcYv1Jo+JIaQYGorFLvTGsR4Ol4eKK
BJDDCC6fTSGe90JJMkSF7qPnK3VpYg0ZqLu6RLeuPI2PO6b0SpiNWsiBzTRs
7uMvUB0Z39xxgV+/1Af0RNrf6gYCAdlx79NydZGYayh1R/y/KM5RgZnw70Zs
jBxpGAl3u0Fn11kn4H/s4apOSiKyRstcXHnZ/zXYC3mRVXvXR+vwEisslIGC
swRZD9uBjoTbGmGzvNkgF6ii9B3p6WH9p5iPpOJ92aGNJfhfxS03uNulewf2
pxeOqI2Ko1Ae+dRYEEoMmzsCIcLcIuxZ8jG5KDV6Pxf9bcgclHVq9D+qk6jx
7ufSjMP5fCe8RrO68gwM10zkDBLs51/UlFQ+3dqUn20Q4A32VC65kooT7bHE
Eb/MD8xAuq9JCisoJTtXcoIlSIsdukiN0TUf+t3e2gdOqgIgqmeOg37NmjaO
gU7vIRZ37ZSbzL8mnYy3yES89e91rRBjQfPLu4GeN6J+We5RPaPazMnFZ6tZ
KJW6Ai5zd07upD1gt0S5jMhkFtEw3PsHMttAb7oU/UCHjQFrXXv1pFVnQ5ZW
dYFFvRIaK5/UXZRtBj5hxA1MmvTahPQyV8ALKEpYbPWeHkdabuY4E/p/tmFC
nCleXv2kHVNo4kEg6UuC1ALFP4WhRqbjqlVRbIryLK+Ck73ashsGLFRiUOBd
Y4vyz9MgfSaTsmSECYUVPUfbaHrS8yq9AsnJxXEvxBxOCB3EH93GWJqJ0uC+
uZviI6wSvzbDfdebCfCKG0Beb/2q5GPI/5RuC2SpCZ8mgjY9Zf5yTBM79zi6
q/1o4vMLloB9jy8DFbxFVvcBr9yvE0vIyfmIo+2KiZq77iE0HlCUupTPa+rx
KBvFWxuBIYAPSKv8P38UZyKCUserfVjFhg0c3o/wZws6UNgqHfTcE8eGRqlB
ta0N6MhA1rzuAum4Q1Ib7tdbsmfUFClBhiDHdGIXsQjd8Pl5woIGwv45w7vY
RI+7tJb4crXSPiDs+cKNpBhZy3So1ynlwMsHDIkNr+hrHlF+BQbRIwQ5eB0A
IeYkPuU6PL/cNLnvnq9TAUNWEPjNoXhQ+wQYl408pcdhbTcz66XCIqp8Se/O
6kP+pBrC4H8uqMiroeJYJ/73S5fTw9SOMat/uKg9R7Lkvh25ynslwe/sbaZ2
nBGmRfQusfKmEf/B0y5W38DJ055JQL/tPEWvQsRfMSGSsU6ruaVyBQqn0Sji
MEF9UW5rEmNoc0zU9EJl5vEHLgBo+RceDLaQ0ilvx6F7SlvT1DJvvI9PJCpf
uuIO5P1a+TMjsDu3/gCPLlwGURQbBX+6cVZZ/dzCDxbWbRB1V1jqWuSFQgV/
uYPAaFY5U9+5dMjF3emK20yEioGEp56Dn8ZYc8vmd0A9j9BuAPTCk2LvHfsF
7Fqwgn41/T7trNLr86BNqM297e7Ur7J3+aISzr3+Hv1FVVD801NnwCDWx5uU
2t4Jac1ISxjai2w6LoukAheCL6DKbx/I2tiPXKxL9CHyXsDiuwTRk587mFsC
UoA7IDU0ZNnccf3l1jRhQVEahYlEiRVdpb6QIpD5eIaXARaesz1m/6cWHbvc
pdsZWUUaRFJoDyHNL81Iyfx15k2j1lbajthmx+T/mzSu1TYYHCcr9z8izFDb
WKk4XYh1EcKEKdu0tQZ9YXbCaWNnDEg88CXsnv3Lh8OmTqavGuwReSXk38CV
pfIJY1MpoKsPLhi1qWikFoGtyaUbqXLHyzElEj/6IoWnShjE4ht1WmN6abPs
Q6woIdKLs8W6oCF+i2lDDGZKn4+p5KYr1GeBfMfZVJh5iczseMV6MTwB081n
x3FVjj+HjeITkGUauHWj5aaANJ49zDoaz4ipsYeOKVrBf4kCD2HgMz3+f4F5
RNr9sQfyiCbrlVKsYXkfYLrIDsmhSJ/DgL989uS/RUydOVrlFxiQg+lKrYZM
25xcSH0+UsbQWmC1CMRH/7IKg0vRx1EClf9FdJ8rDvmmV5LorNfXR8GT8G40
/QTlpvcsTRl5ICSwsTkKrQWmIszcKoW5zscj6/R/4qg88n0BdOW7RMBykwho
5QPe1+rS/6q/fWZHG/zl5oqRwxqn7iZn5Qub4frX6csy9tBtgDbYZOYRQK+y
b1jZXav3uciQoetYPI0Chwvj8tRnMyzmyjFG7sRZFKbBNc0xgr2qcI/w5qBA
NYrUSV6fxMb12KBWbT1dg9I/sscifK3Z74E70irTkvyXyRwZT560b2DVBxb8
K3t0HX+0fIdIRFq2z7ttSXr7+mPa/trf9q6H5WaULTS/fBtz12VhWxpVO+IT
wLQalMUarDDvJpUE24G87k6qSR1ZN/oiZnmZOlBiFpf/P/hXjmSlsEwWDCcz
aNseiOIq4uyLBdIIKeL+1fMUIwJFkmbwkwyTBFSd/xuOnKxFPBeD58ZgKlIj
5BPNa/kBhqPHucSt258dghsKVtExmNqEGT5J2+q/fuJfD5WTVeGcqgy79IZW
yKRNwA35q3C4d32J8vvDfrj1ENmspEp82bjtoaEYq+YKlW3IysEuR1XDqrxA
wM1CyGwwEXvfsgSo41ieEEbFihWZf9oyt2pUwPAYzMx/WJfJHEs+C5ZV0uRg
0hEiuJk/7w5pP0A0os0WmdolquTiaOw3NUFtm3nCjNqvTSXRL/g13EVUC5qE
jelOXeI33PA04QL196BNV1BSvjaCx6VFVihd4pMWohiEIDF4424NTGDbxn6B
cB4HSibk9ViMy7eG6VvTXQFqCNgaTVvGjD3SmSDg1EFYnBcGaN6vivDUrL0V
kJ6lvk8WXLbVqsobDozq5Lz/V/CsWdw8d+TmWl0KQyAk3Bu0SADkW+UpZVa4
FMwnj76WWozhin7cgY4lrMwTgX+WXbfzd4X40Lto7OLkVuHdwMZCTl8EE89U
MQek46kkdAWt7Mp0FWgrvKsx+FkFnmSECCvBfs33G93o/Gs/HagrNnoKtJxv
ZhEnw/2BlHIaXR/i3UgL7f7+m5a4kzhYcSl69PZsN8eRrypDCwn4xlVbgRxh
6qQJj9zICwYaGswcyQ3eMA6IaYzzvAYWkm7keMutEfWqUystEkUq+aDShKPy
S6Y09e4jmRwP1oaPoymZe3AhyFuec1pdIWZijuRd91zHieRy5zq5HIrxVB68
m/HuyiXJBWJAnYBJnDgbe+uGFDmNb+aix69dq+Ma9IwCoy0t2nu7yADxMqtJ
SiNM1ToC5/+kNo79aDf1R6uTTz2f9xXkOe29dYQWVQieONyHkZOW421grMN4
TFfaE1N7YZEX1Jcd3s6IY6Mcd7cuyAdTGoZ2zPwyT8IU0jTt3XKyzadoNO4K
RU90GgO8OPPynzh7za56z1e41YE+IE3iVSVtHdB4q3FeLdzNaWjJ8pVA4sEr
jf6nePxFJxMMBj2HecmQh5mJdO6tWFPdw4z/tHY/GydAJJCLWdpLYrTqsFln
xraRawYtR1Jh5J6btNth/E2hTksnJqXPxgGi37nZC9Key0VT38lguIvY9JKM
Z4axy78sYO61NTcGa72LqEDFSAUPEBzdXB5lJoE1LDcc/0i8HUui4wnx/q34
vDj707C0gV+R2XzciC35piQz4Y8oyawCGP4DlYEg0/yL2DyO1ZuT2TMMd1ry
2M/wndcuIdSBt00RroovydNwUKL9dzMd5zKjDGcrtlSVHYKTSn7AeZiUDhMc
buMbCHB7Lc/ES+0sJUfL7WGICr8XXpiHf3q4NK9OiMFW126AJCiU/XZDQ7ya
AtXEEj51cYAwqcTCLD3RvMdaO4AxPbBazc3A+26bLUPfaqFs9IpmmfRQNFfy
bYRAXt1ZtpRlhF9fJkRQcmNJX4VprM+HgBEboaO1zA6BnO9QEnfIgPbAerq5
GmvETnTo5co7QBSnH322qAhuLjsDmtEfl56e0AXZDjFnDOeCIulBqD9PJieC
QcaMWom3licOYhATka5k4M7vMxjhCvQGsuulBX8unDHc3If797FDUU0ik2tG
aDaICe0uOMsf+QLTdtiddbn048PF2JatjhZ3YzBv8oY0BN37araksuvaoqau
Qa3kTNn4C5Bfc8hwfB6drFoAHFM2wdi+TffdkVCk2EDvri8KzGFuYIz//3Qx
yNWJgAgTedZ8n/pV+jfpejk38EtMgkvNCgfUjuR8Yuk0dqDvF5OG38Zb1NEn
6JlZpFfmwrWUNaxz0x6hRNdFvlbGWG6kkPWl14gZs5Fa5mi+J5MUHsEO5wx+
O/7pB3WXkmJC8j34crQ8GNPOFO7pBIAKbguCrS6h1/ViMcpeqnOY1eUXNebp
IXzKDglL5boTwK5KfxaXec6+dBiLrMghSlAYCjmOGA0gHJi5FwsI0yRm+Rjp
jEz/7vjLn1le+mKIMGde0KgMejBcvO5bX7pk7RmGme7bYwexBAzJyahZ4SR2
GAMzJKafA7zH/exDwEV6nA/merlMNwzmfEm/toonh/gHaE0iLJZ/+XnzXYOB
8vIV3DE1vX65UsTbSVhJb76atWSeAtV3wPzaPrQBLYw66p9JGuimvpsRdUMC
HKqO20EeJaE2Z3uBTrbhTV+gC83fRRrWj/PqCs37NKuV9uU4u/hSKlnzBiMs
34QaIzsUt4mevhIdSXTB9CE3QJLB8mnP5llZWBeqCmbRQpPQRCsAgIqqSQ8T
G6tudEabgWaBuO4ZEoKY5gpL+Ve12Z6sV25ZVk0fUZlgJQ5oHryvRq2NuCZl
5grszMPkMf/9Ruk2okX6qxiS2Dpj5Yy16+pLv4jAmcN+tu6M+2zwftoniGee
8XpYyOjDWeN7uoC9h3rgevQfzWPtiKt4eIfUkgoWZ1YpzytTx7UJgJHs5QOZ
+zrt6IUX1snu6ltnigftCwOKFm1N+Bx9094huE5vnnK4SM2joLDrp5uiyU4w
n7pR/AgrLfO4xNcwwgdNtC62E8TXpkS6FRpGhMPb9mJdaxPH/tno8NHzT+qp
BiTw7B472hTAMjUpYIMEBAGTEpm2AuvvyV5W49JE/qZNtMqxt7bItDEi8Uf+
6VrwbTq3A6dF45zm90IGfoeGIjZQQeZMjhNdwTc2mRMz81nnRdGvix95Op5r
ZzNwL9m2AxjUUM09h45uSeUBiwI68RoY0lLSuXXI8tsvCtrdHDg9a6FR4QHc
asHmH0Yky2xqDenEe/yUmN47RL2pxcec6rTXDPNjzdgnf8luwwHNUpG4Hjzm
aCBhD5OwKlGUonOoNez0i3GuCf9D2TGv9al+i2BH4ngKfOSr9uSYPxStwU8r
dYicYPwta49PADdXwGYucZxRbloAqjO//HjBzonKtvOrkjQa/B12RndHhoqD
uekrUvyJ2t2o6gmBCH2A0SUcFz//EhNoTv20fCst6YZ9vkmzHnQD+LL7f/KB
lTT/QII0jsnHwGtXsWWGwiw2xrSJU+Vn0aL9746Fj6U97ydWtGLaAOjmHQxq
qcuONl6WFQBHGpyLrljbb+g4o3Ul72RX7dgVrqWC7jnc22fj05rBSZkVBgLv
CqQPHfwPuudQzZ2JequTij7V07I2a2LG5gYP386AoM0YJtd/KXKII6R7xoKv
gu0cu7Kn3knpj8RP8kMneQjlrVPjQAywptjm8PcHR03mRXsF9MJbbEaUTIWQ
3JVq97b3i84lV2k7+O6XmX/pX0mat3XYCoBIK/tw8AmhprTfjfYLRO1L50RJ
MIfxHrrIwBSAv7dK/r3N+u7ja7yFs+CTJ4uQxVpdOCNI8QW2Mepy31tFGxC1
pBTQZcNRD5ExnObrqSBL45Ui0ht2TfzvvB+Lzz5QceYR8KY07tL744lyBe5J
w6bYzFb/uNa9+eF+8me7dn216Fr8VQCtmJPhKX2EQ66ZGCZ/wC8z5NKaaego
rpkNspbHY8qmwmtHt3ILsD35eyDBVzybx6A0qLTss8K3dRuhB9x4MNDGxpcG
g/1SKOVIic7RTZ4GhMEPfF9JFvbmm8yvFLrwBvdm6ThkVxWHGmuX5jZYpZ3/
tBLujiTw4xJxtEvPXQl601mNLbOeoDQr6kmy8efa0eUq6INyJO5LIQb57Ff3
2XrQ76hTsPoBbYJUqKQaluq21w2lcsgeZDaAEkcnmjYX5Don4NFSHzDYAVWd
IyL/0dUl+2WEuzSIwtrPS4FBiKBr8EgE1UiInSNIou0unHrlxFFGH1FT4ZYM
Zsrr2tQMdjqoYhTp3n15NQk+c1w6TPfFUa5j1f5OBpxuEnmvBeEXM2A9+K29
LRWLXmjFOXFBYdiVcDemh9uKIISjNitzgJ1CFOKKTPBySrLwAnJl8fgMPnJp
aUoK9oQMH49Zs1iekdZ5Bf4yjWeLEWfYcEh4Tos6gNv6PI/Y1Jsc1d2OQsS2
5/e8fnfgjvpqsmYDUl21gc5HuCOYhqYLuU+4+Wl3fWxslxUzgY68W0GeEXd8
UmgRBlC6H6ov61I0qBImMzHQrZOXtKK8ZbViruhYyKzTvOFyJOdHdJz0DOWH
YAWIdCh9FDq8Cz1favfne9yRTahhlwoSgbZ3GvLJjclhWMG9Oa0VNbs9QS7t
pplXYMHaFRht+5WEIdEGXwy5TOl+USZqRazTZSRXjjgcNyRCgW8gQjJYkRHx
txxeRFWpW52xeH8rwRQJczXmU2eyBcJ7HfWYOIHroXol8FnuDb4b57gIO7CY
E6lKeIOIAW6VASRLylzWcMMxUVI/xEj4PDlWDDOLBYwzO/tIU+91I+Ivr1NW
rk25MourenHBSUa+qbssAl41H9xYgp9g/XlLXVqMBkfO+jF+rSeaz3IcH+xT
QK0bOKnvlIHPhDOukEzXjpONDH1ue/Z+iVvPDFsl00qPuisdVLrsoizdOj00
kWe4LYtyqS21ijwvDUN3ybNoRs4HzG2n9EggqF2BT7kuYaRgPzzoFsNk2DQy
miqcruSIQwL5ic4xHjjpzHzffTMVMoejwlYR4MaGYpedF19iK4kQ2lXOL3yJ
Z9LZIkvpE71CQR0rgu14Ykx41kLp5+Eu1OO6oMIb0z0D6G9pn89/exB+VmRC
po1sUMnRzawGcbfufvyUBWUu3ZFVejcSBIm/xzbZHlK2AvIoQqnOw4FqTzn/
smACUue/QivwRTfJevqNU6yipjGDMwQtiorCjjd82M2OTkXbZd1crnJAEzUx
vb3LO6zayL7pomHY43eC4pxdR5CWfsaGBhIrKTErRCTAUKQHGMVs6JxoHJ6X
zNLQtWNwuE+UojOEGkgFJjpWBRfnocOcdqy1+IiJWcDyp54oiwQJstvMIxQv
+BahlxERaEeG0S/wjaYZZ2jjMtrOqhhUpOL77Plwk4HoJB9eYHbwpnYggpk+
wMI3OkaFeU5rjKEeftM91/G+faLZwCHwv3y6yBZE0RnPly+tyjKlWRwzbh0U
9IAnrpsGv4erl1f3+K/RWuE4tuJlZk9cym7pf4wW/GKoqqcW24ahuUVBppUp
njIVypB0VRZMrN08vKTIo90+fWKCCPOlXzPRVY558wQs5fObEuba8kbm9LBv
wKuDRwkfpwhaafwQKlzHAFQ+pCplFqnT+KdDOEk6daN1xDHEK2pAj7xjXFsu
2sEZ4UXULzLipZe4iIfwmFhnEphy7jeQYnnOjqJpSMuCXJ9IHy7eF3pGCutp
6RQJwr5GAzQ3ILTFY3czVQrXHHBd718Mx3j0cvsMoKr/fTIYJRDmS+TMyL2/
CElh/tPIFxCynhlAtQaxXofhx/NQxuolasd7lsHRpsafhlCd3pSK8G+cPhFX
r3+opCIZiZ+uYCNwDqo1D+os6Y2K1/K6McfScSKNRD7ZzgxDEiWKcD3SbszB
B25poO5Ll10/bPJfE9sL1rYRwVD6boIY/Kop32LSC6zS8RRRQAbPZUZwQhsR
38OBYJH7OiZgYI53KmhUwANb7N9amfK4d3de0GuyEh3F1jq2dgpLAxM0WP0g
XytedK0COUICyVqmm/fk3Zn/IKbBRHrjeX3XVltZq4wEFth3CsRma4yoW67Z
PDW4xkvaJuQC8sRRBKnhKDLva6Sk7m7I6uKHKlTDtxRhFbp+FMsyrNP24mKX
psFMctKWjiN7qcnjf/vzncAkiRV9V759ARG5WKwhkTR+2PKVXxc5iwxdBJTw
u8m50Dz8SmTvLmC7VcYkeKbZtmCu838fAoPuxEa4/8aJaN7M6kmtmfpePVbP
EdypQz8+bV1HSR37jiBDvjbklXGVE4EpcK6L8yALQHxiA2NhdBzn8R0INYg3
Srba2vB7JxVXIlo9j4Aju8tpET9dPncQDecY5XolMUSpL9ZjeQ7X6FRZTtSB
rHeHoZ8p6GJFhKkLpqsUOKqmZcRxBdOx/EQEh4lLGBXn6brQIxxzsOII8js9
3Ea+IOxcYd61Zn60hdN/YkJBOJ1uVzD+dEg88YCkHySMRnQbM/sXhyjtFCWE
oN6G+DDOCn8NB85gomaDFDsVzhZbLNKOwnbjj9DlIjEeUuFM/K5BeFKCIeUh
kcVgM/kT1+XPhvjuWIxx1ff4OzePWL9TAtOVd4QRvcqt1xHeXJhh6vdLkvBD
93Q7+9IVF+nG/t7lUq5XpWs85dJUZmTbmLwFcB479diz2GvwdNIW2tAzwtFJ
UZBMEkjVqTL9eL9Gn2SZXe/zfftpeAyLqaoSTRnEi9/1BFa+3Cc0cQjsetdU
MFJQuW653eA0u5RkAKgzhbyQ9tBbQ5G25x6GF28RBJaKXt8rDdTqMvwCcicX
6wWsdebm/jN5T8J+YDDTdKjBlS9f1ly7jUZVu/2i0Gi1BLDdeMImO3ZzPVKg
qTNDCC56anXnXE0/ji5cmq1wqymhOM8/U7AAP+sH0f8iVcYF7tLz6ZN6ky/K
AanzWKL4ldYf15auYpo1YGj5NnTMmRW6KhDurwcyyd3bpWFX9XPumVmKj/Zn
DBYOP9aF8wPqypAv4VXlT17F2X2evVJD1rlb5AwKgYtRgt7sD3w521vqxGXF
mHGZCJ4TwDNV2T2raqdNP74gen3QktyvAjZopKtMwOFzN3B2SyBalgyRLLEI
ULodci41NsH3XGRRsq23qGClYtyLfmKiHFkjm7+4Vd3iLzSqlS+SIo1sM/lN
6to4PalSPwtSVXLSZlhHzGPJx8DWjPJMvN8H6EWL45gv3tL3WBHZBz6T4wZM
P5SmpU4eVjGaO7RbDRaP8TGHK/uiyQMT46HAbs2EzT9Uz87M8bieTiG6+NUA
Qk31IW65qfTMzpMzgWus8aYDN6ivCvKnPUW4NXZsb0w3jataMMXGna7lTGgK
fB3/xlk1Tja06XBKVZkLtbmW0fcR3WH109RlwF9qM1JTXhzmJknQr0+6ivl8
EakuotO2zrIHuDx1N81rSDHiStQO6Tdxs2x7HgUvXx+BeUrjzz/SzCvJG9gN
cGiPwx5uCokaI/XwWN2+ZvlPkcXRHUVkEhoPEWPz9LZPCI81JYp9aNzDxjKd
FrBluRGkTuMQevX03occqYdy7jL7xWZUM5aWmUDOJwVs33GMsRWhua6XLRom
tL5CWO5zspbv87rE1jr0TfqHDCIbWs0LdVA29xTXZWV2sQOjbb2zzzeJwRUt
8/i6muo0ApcUxtJqY4NahCp7dp0YzFPOjZ+SE9aTWi/8Xu5uBhleeSOYTv29
nyfntWupvgaZEr/w/QKEQywXtfRjFyNFSvlbx9b3MOaTknUljvmn53FaMnCm
0l5L1uiJOjlyYYD46Vd7/xOhXYnWkyCzUsdc5YlSk6TPRKcZuCxVK70tjWY9
J6lO/fDKhfC9v9hnNF58b0uLdy4WHPW5V2dlyPjNYpnWOUsQjO904DsuyPaE
NY6Si2M5ocEo9d0nKTEXqm5+4bQQ2UyZM7otrOF3ew0WjOCoeyKAQ9mZFSUL
2avtBp2+qEFe9zRjypkIfd8lNXIEppZWg5h2kKtg3NkX0JrCzl19LXY/HNYq
NYxR6b8drrupckYy8K2weyk4BLIMQLu0yo0tmu6HvRhPrldWs8GdOAJvvNIz
MSfhpvrlo13bOOL6rjtCkb9ebHsP0jkoFkOrlAwNSzMlWwoeyWzxunjISNop
hu1GEtT4uCa2R3yR7VD7hXT7mTqBKlADnUb15897dRdkInWZyuwk7bITucKX
+kG6ap5NxrJhftVT9M28cHLGxq7VGO+MBslom9wJQEhjjgRuk00N4J4aaTKk
1DyXJXZAjq++WtJpWD9MV8jliZqCd89T5bPLrlxKnTqx0btMWSb43m7UnDt9
ysHLcF29lAmVQ8m/hQ9VrMhOjJ6fTWHYcIi388lL/FCMg/GmqYVG0xJhDRXW
5bG3enIFoocbVIBzLnr7ORipNglzUGBcdg++cl/eH9dRvSE/R+k/FOcG2i6M
UaEOORKaq2QeA8TGh061yPspf716mZFwFDlycCjMU/4I5iqyuQ1avQ1n0NfY
7iDSx+54mMXrBWeHnuAhQZVlP5DXRxW6f5Xf3uGiZvfEDPeP7j2O9BmZ+e8P
ws1Zd1uvS0iGrdiJ0gsS2lDMTJBzl7N6VcfgDW8jl07YhysJhlPAtm8WAlfo
O13EPgbjhb7WM/17nHw+BNlRR7fG9N6SZurfaO+jrOKhVFyKLsE5Zp/Qxaok
XpLfe3cTEBPc2Us8syWxYIc0GhwsrE0/d9KRcU27FYA92kGe2cuTfP8acCd0
gaPHshmjDqh+VszHtUhBjHYW5fbbvP/EbBlfMQjfTOHLVASywOXTVrISPYVH
hMD+yAnNXJGlL3jeyFRbS1tY8mOh+cjv3pkMP4GOeA99K0hMQ9KOPB10lM2M
J+OdUF9PoxzGv487yUaq0tUUgDQC5KzVHVjQqwgJbkC+1z/l3P6IKCv44UYe
/U79T1nAJ3QL/m6MsMtJSoMkiH8BzGZfP0sSrzCdkTV+802BoL90hX2aXRpP
Wa6VHKO9UB2+SDTLGwEMm2VqstI/pmqVohRSkphC5iOaocon2h1s9rLnekaj
0m+drgj0gmhqrbYCP5uDDuHxapyzJSb5h/FkkmV6LKc3IyjwDl6KrrrWC0K7
YpVWdgoUVTe5gACKEbag3vkg4RiHEUGVIXjBKlKWdzbiXClDd6HoORy+yhBI
bxrv6EzL9dLGZ0liT+cEkQNoWSonNYvKTyIvGBggDvMHH9VV4XYfJAxurUOz
gxpx/1gtisc/niTRhfI1VH20NO+vGaeGRDMeDNLYopm4QbfXaecutce4+WNg
Ad6hMnGq5nNEPIu+Ldo+x09PVP/jZlnQFRFWRD+xa14BkwNh0xGC38Ba7pzP
7UDP/2KiUSyHYguwPZ6B83kuTjb6IAS4rqJdxLPclNUAMpL6dnTexP5G3uyZ
mRRBlQmrqBxyCO7bAxFr+KSaOl0L/YKFRE8IAeWzQXBMdIsS07xxavsPl8Er
VBxiYO6BKSamD/iaWnAjHQOIbEJKsnDu4qeF/wiOiYZvWtfnYEFea6UGqQ4q
v3/9QRWGU7vNLJ/t4dysOEOKOYhr9I+7ylsGlnVD0in90LIqVxSDEWhlKUQe
8qt3ASUUHrO6EDzhfjQlGPsItVfYuIHHzSfE3rz1wGsKVY6hcFZ5bNR3DL9W
reuxdJ03SAhp+FZoZ/VtU35hHi4xkB9zLBglg+zeiJyuM9z3FbuNB5ZhRwOX
TeKTZ9C2oERdRozc4i+9qX8hDW4IT+nC6zK0Q+bcXv6BusCgilX2W7kY4kpn
lam5pFjp/7Tqhbj8U7oDEBpeG1NWJqJB7xcdskmkbVL9PmW1WD+Z13Io3DRg
mG/uarBVL8n2Xxb+k73/Oi/i/DpSzf8tnOFZj5sZMB3MDFoOnSg0AHRdA3tq
aZwa08y6FrKyuzFs6yM11aASrm+dTj4wdK0CHzZvCMwknSMOzHKMjGDilxFR
bpMCFC4vtvhG/GPppyUMygacw6vYaQ0JuDQCdLHO1JWLesaDx6V4VM3qiWyv
A4r8s70CU3GsrAyxA+Dklsf2F+lqOLnT20p7gTLCapcuH7uTnX1cR10K+jXz
Txf5uaYafrYC9MkkiDkC5iPYCYVuN/rn6cGWTu5Kb786UsIJvvgXzKJ7vMPw
VLbGSo6RJWyJwO/ckXT2wJZhWOwbZoce24AB9A7EZby92zsuitl//gBTB0rS
y5jKMU22TYnX3Sjr7kly2YU9qMn4uDK5+y2pyFnuGRCDwquxLjAKfToWowU6
cFAHCJz4s2wYsYxNEoo/tp0REa9BKcdnpO1gA+VQRgar+VHx/MZpK4sPSv62
WJIEDCsRZkC6fkZVM/oeGv2k5ImR1QEJ3MplKZ1lil+YRdxMnp8TUqcihkak
Dud8I7KFaTgPIlQBVLD5IeK+mZXIDWrIXHFtIX8gEdUi4/x8RXnmB5qcggSq
kvc1iywtBPrqZx9TE3Xp8zu5tzXC4hktVWO5xAourey6xrE9v4m16ltkvRFB
7HNJyFVZxoqExzIKrC5HCBat4zF7cmxgxEy/LPdF6gWrs70cnIap3tx6triz
bR1kETyesaA996ITiCSg2GFX0IyWV0n6A7OsEnqieZSehbhqKvS4xwrhDpNG
ntthqBKL9XjviQGo8BpC+lf7sScZBujiPRs7DGwoA6GgBpbY2ZpL34yrjBJN
I/gxpbg5wAHxLG8CFB0oIa5lQ23DhyUzh7zhEGuJd3PAVZLqw6lG5OPXT3gO
YpMhAnTdTP1H7TFQWbNv+kUhq18n76l4thN/vKZGDZKzZkOnlj/ED2pznZ9K
VbDMgZ1oU+QNdzGPwwgpebYJyrtOpeELc5mBXefOLDXSE+qsmganBIxQmcNR
del8p+gcaP879M/tEyKP5Jk3wyKPkuk7sYgJxU5EKmjGdW34hMh9H6e7mWNO
UYg/F4ZHhbeJDDbuIdbsmGsZzptS4mnVH1s4a8cbckb6GOezMf7V69CrPSG+
R+TvTB9PGBSXloLeQutUB77V6MZf7ugOR6dTD16inTCIBK6CO12bKgelkGtJ
sMzmsl+Uew2kx8Da2hk+monCU9uRsPPci7YfZkxg53H5QSbFQ9tVi3Lp0fLV
UzTNZeqbO82Sc74Gdl4Lk+D6i9cfhRlQ7Cx2X41keX7CTIuTlac/2nACAAph
0JL148X7wlT4FdsU8mKzjnlfO+n3YiTRcZzTu6cnKlJ81NDuGf8jCC+8Cq6e
LzafLUN1vmqeaxsp3XONvb+qAclyfgk+j54UQmMGV5ByHVJDVygsgnxG0nFT
CPdoyc4VCb73Mj0m6JYAQqT6ugvS2EFIczpHjPu3HR9tVIyfknGTbWl3YRjN
+1NT3hFd7DRAJHvQxI5EhE1OrzhqEVnGcG7ywnZyTb77R9m2MhX7e/lENqB5
33KqVRNjhHC6R49wShL2bO4D5DCVeTBJJWycEB6bb3HWQCJtU85HL1Zpp0Cq
eQcqzXIwKpKUcopSfi43k/csOk6FnhAENxjaZh5tPvSKW0MQ+thTkm5y/HPk
fGameUrg41+Hf7yIv2wpcBoEdC8AW9ztglG2qQd8Hrmm/HYyhDtvcQDAkRvV
sRO9leSjjNeowOAVi28ypgb9gdzz/ELfd7Rx+LRmIJrBqAzl9S3FllGOeXyD
mNLyIvFEyLfdUQxGM5ClFttBeFM/o3bnARLi0E5mby20+Xz4cP93NMxTrw4s
KaHshcHkM64zKDV6Nc+HIqQGzq/w1u8kNIPLbDHrH3Ltz/yk0D+wMP2tb51M
c6md3FrfYt+dlJJ3TEsh9HGU88SYXFYBIps0S5YAdlIz2LfdtFEW4Dxt2gHP
LMGepJ5mF6qo9hj2Df5DWmy+TrVYYJqQ3cuzR5odQ7BLVxTjF96+WIBJ53gf
FbyechhdFATOpNisXNIRFXa9e0FoiZ0uhVhBQ3K6lk/zXn1mJpGTUFx1DRt3
Yo4WJRWO1+0lstkcAteDPhTXWxNK9xPFxrkrNiVN9OupMXmecS5Z8OgsWrHJ
4XZbf9eVh07h7zZU7c85cj0fT43mbmOeFI5cg4a/A3C91zPT4W4I0QORdz5/
srT7j9LoAp6jFcbgc8/e7SXKFjfBJlFVqunQcaKPa3FTAlRL18A+kybhdE2w
2KGinmBjy9NbA11BxlyS2K8ucb/zn5fdTy8soyXz6IbBVP1Q6bTe9w/Emh3O
TsADd3NjWyk7rx8F3UlThJlpheVNCFP8idNkpOektWwxyVpIg4xYk54C85N/
Ug4dUo3QzKRVR+d0oUfwKWgGsUp2uUa+mxvc4kVgbf2ec37kUT1nQRyqCOkJ
TUuE7J6gIleFodPQFzVcSaEp6JvRR6LYaE7uGoXMNOX6He2KzTpfjLFZMqL2
v5r7MsIBzLfV6gxLTZBy+ic7gU5cqPFbJowAPx0i7xP/YkCUpKlzwqhkD37p
BiNd0YafjT/4S8xpD5oRWJ5H/+QvysdPw21w8AkF8Bf24/AUJiXZ6EGkUAKa
SF5aLlLdEAEIIVoViC3087ZwaQYhl5sLi0ML6DiqIoqavKgNKy5KGegSZcL2
lo17WVmHSpumLPID+pXU4L/AcxNnsDC/Mpqw4MQjM6J5SSsib7puU3kYdWUT
QoUqQlnZgRHa2hG8rPZu1cYPmo3QmYVL4VlDXODY14OBDPBNOPHu4fnASTGD
BnOS91efMYLPvVohJdNTq8ZLbMwRNAyAsq1SCTJGm63Z6Sz5GvTP62jsPF0Z
1m017KcsXuSnmAOVXACkLHt4jfi97rrctKBzrqR8/xDli55/M7AEUQDKcsO4
ZVDb96tA+JydXpj2kUL2kgsSCAhqW06VODvZ4qbfEq20A6YRkkrw9AHQBqAG
D1dIyGdCJpi5b10rUJKB1Ly0Tc9B4a2Nbljm7s/OQpqNwZLXbvEGKZwhAZAk
y+Ry3jEpGbjUBmeA5hHieTXRbK/+9l5NMXY/eXhtd9u8r/kdBOb9wMijqsPP
vRSwDtK1gJIxfJ+qV4LkPnFX35e2nrbYq6/5lDLFdyXOQHqG/wgU8ej6I4ys
MW/GYuftC6MXgioMvlfG6ZFYEks2wlja/ZaMPYI8/Pef5uWkms/Vu10y3lzI
z/j0yvHMiDeu0nX5NyPRJlN1vMLme/+p0YvtwKUilt8UQeZSwHd1Di9mLSqj
MLYbev2awkVxOTsvulfQmVM7PfKRAsbh28nQehT/WUMuMwnOkw4C78qrvW2c
OwwhsEivyYN5Qz9ZAZQdyH2alLjz+Kia9vKnqp2ZK8dyZSEUNcPNtQ38lzwg
msnLVKdfEgbTRzI3C5Fr10huX8DNh1Xo70ZvN4WzJKRIGXm/KkmBKCJHCtKW
TpbXejwU0n27zroRcxP507XSJpZlDYvnW3fDrkF1108Czu/Jffm5c9hwvSe5
Ofe4800g4cxctrllp8/4kGYb2QiMWGk2z6qhIs/w2Ko2cMq6vBH/OccSyWNQ
RdGRbGCU7reTN6hRBd6NESMZn9GWSwg7ibl7MBv96H/r2yBLSUogqepJwhG0
czScWqSqBvgL5L5mg70B44ZKq86zOk9XXldd2qphoazDeqsHmih39mPAc+NT
Cp5wWxWn3/SEUxsUhdscQzkBj4P9dUu7KnYwscCe8hs3iZ8fmQa6w85Wihg9
oTuFH4FxoGY6trUKIGS2T6bGLrGhNlcejfhRIJgKbjki+xlrQhwYqdHBymo2
ol/p/cPZElJQkgFf0dW8TuJ7oK7y8xVXqNowFC/w6RVBPiWeT9GfWQ/PqfVN
aepEaZfBJx8AcqCUUHRhHGJ13fTbsNkovB/Ydq0t9BVuZ+2UsVP+FvZUUHc6
ktCH60J+t1ThK03KpyAF3aQjbkM+HLQKkXBCPsDL4AEkq2O1jIELVt8sHDFJ
q/YcCehVRJnsyVnjMQ6zrRjMBKWXmglNm3mL90DTGZM0z16Eb2grE6oI3pFA
5ZNtDhm6ypilIlSEfhBVSsSGvTEiLaVnfd6fbCPm7YNKYJ/z39SsG7+3oPMH
sU41Nh6B4fDKz8O9e0G5mv9l5a2jaA3GTuN1fa+CYPAf8FkgYoivcc93Jvmw
Qp2UFhMTFLF5TaBpAhGSFTTBIIP+cZL/fDi8gExJ8icbKN2QaX6mQSOfccNZ
zmDs7EZNsgvqEwImdi2csOz85AwXXN4AXiuPE2Qlxm6kRx1dudmFFlnYYpux
sj0eRHiVZBpALCQBqPg+5bhwQ45na9thJuqkSFCPyVCQSp4s7YWdes01mxkz
h8rjyYa8BNTvm2kvo2R1utmwr/8rxT9bmk4l7hQGKM/xl5HtC+yfD0nUJkWc
6TfwojM2sC4nuKleHhuemW9oXoFp2wsddmnapQ5ES0bp//wxw7hjVJMiWb01
+ovu5lnqYUUxSWaioWC2rF7ZkWGZYRhbOyCfLbRiEc/KkrLWAicQGepw2Bqo
nGmdGyHBUF6Xrd0lfrPfMKD6goLMyRN+jNlZeRkKHi5xvnQrgIqOiDzMP5eB
QtW9/jNsyfXEflJFgWkHralLKGpSUOJ7hhyt/S69V55nulxS+9fhWsUz4Fo8
cIoF9wy0OJZpJnXkQnhO4cOEymWhZV2mT+lpAIRGuiTAYGKcdTfET24TW9hh
YSUbzStIITMFkupdN2ruihGThLll/NwgiwbiWZjz3MbNuJCfZs5bbVHAFhcv
LsIw6zhU1bXklB0VzcQhqE7mKsborZTnJFTIWjOkH9kvTjBdnchmwwcNJ3YJ
4LfeqYnTJCPoIW+mULUVgja3TAC4zodG3bTy0NPwlllPNlKrqs7jvFrY9c0Y
IRNIrFxMIhkz3ZFIijQdx9QqG7AfLJUHBCoVardGVI/T9kcQ2qe5Ow75HXaA
vbfkh90NL+rZNjLqxEhyDSkc9iMR9L8Ck+BPdUHICRA9FNIXUAApET88Ook+
ks7ZsJ1zwaWCO0neaAsMm8VizDB8Bggb7bqLWcS6RmS/NMfoUpdYGMudQDiN
CMV9J3P8e+oaAddoTiR+FWNlxtVjDu746W8je3RbD3XmflUL8gssQAxRrlBO
ontR5VnsPp+rvHNRjTnPb2+4BGYDwQH0KUl4MxOTAT6VlZ9D4S1e83jJNt8F
OhoqVy+Wkq3blWyGGunh+HT5byGqunfy7o/4TRjN9js86eF/+0qnwfiHWIir
HRoZXtYCf9J4fZny5dnw8CVWeFB8O5n7JfTPzC4F6RWFVCToNkKtyvnZKPyF
yV2KVIdCosSA2iEHad6fpy2NSFByZ+/yhWDIPjHVNfQGUGkHgdl+Rv7gKqEa
JjKE4IeRniyuxHUoJ4zXJszR83VoSWq8zNjcCHrssQzOrmpm6/VK4U7Z0z/z
P6tr0oSHH0CDsBgGjrw1K2L5dJqDPbJFJsr11QvLBQvUd1J8I3Xc/HFp1kU9
vobp28I9aDFA9CT0gbDQ/KgzWKjFyeAKv5aT0eu4/3xkbQ+CyvGXiAXHK1eX
WLANr4VDVaqvV/r3SgBvcFjADRDaFzqwkzRVd4+9475iWz9QQyANT4Ogab2k
CPqbwEn7s5fhcQjF6NLo9VLoih1hBtOSSKw0uxQJGp2i/L5vuePEgSPq4ziH
ZkwYCMMVYi/wuPCtVrFeHxiAVeXhCvd8i+R/hmCCJe7f4CEZuOIN12gdgqh8
xNwvQ6F3CYjzVj1e9Tg1Xu9qUsexQ8MRlzPhgzf+SLckStpyCpOMtJA9mbM/
59v8pzrYHxuEIyPgat6GDIlzX9mq57jNT1t3sVJjAClESJul5Th/YJOgPTC5
ZISEbVHduOY+AwRmllnznfnk0zkq9EG7m8zS0MiKpjlbvucKQHzK7V84CnPT
sWbyw/Vky/wJLtlr9zSGNzGaVU1+XK0l03F/PKjzH+bfXtJLPgwxfvtgwnSG
Yz2RIFOf5CajQ6zs0/hwnf0USYMlKkp8+TC+F+IsH0EFs1RgdxogVip9pJgW
bEOas/phmL8CoR8vBYXZWBVMrp36PreRmL8Fc0i8MgYp7s8LXEFZct8Vu2uN
Wp1oAIL6xr0HHWMCkrac0Q43Zo96I24extAe0h4pBYr/FSqfEPwMwBuN0+s2
MNl160OcuKAksTxSIeZ0oW0Lf+xu6uTCGb1UnRxvzMwgVHGtpIRDp97RIWmP
4RlZ13KgEPaCiJ9dhsE/D+hvdzsh+64iQw9hMb5k8f5eeANotNDBxwTa72QG
v2uKnlbgLut5zk7zrleG2Czleh2ArnYLIAwz+Uw2QH1YXiGx6ph/pG30CDCH
hG6hkRlFBgmutHaNc642jQqy43eBPMMs357bBLHn8/xMFI8B5sPe5vsACe7c
QfACuF6X8TfpTqP48KfJAIdLY1uG69TiCL79GOz5E/xH2q7lBjNrrtDEsSqU
FFITFOsL8GOZ8vgwcvlTF8mJSz2fmSXtxUKfd5zS8q9aQeeWECrNp3VJ5jqw
bsJ/zXJ+JZo6lhOzzeTrgpLd4MTkdiK+QsZAZMlgpy9AMdQobAwE4MW1MLUE
MoWJBYqo1v6QjOzXxmbPVdhTXlWF+H787nG3lED5Bis1jJsK8+xkwa+5BuqK
+1hwrk1bUhjPQjaS10zsNnfovHAXgZuMlEdI6sBP34nUFBSE7ZmPjNiLk41L
PInOw8qTdS9pnJ3/0RL22+ldyapQE/v5QIr0Y4xqMJTWoS75xuVlvbAAyesi
LvK/8OnNWCCgiQPN1ZW8hY0kPTDaL/8BUH2uEUrvyFkDP6VF6dpQVRg3oOL/
9JZp8eyOXtlqta0rghltuRvwC+cfcl9Nr9kyZDiORm/gB1VdzlBEKgEeKVLR
BzUrElO23FnQxAm2wjBlnTUMz4V6Wq0+bEw0LckrIWFV7rRszIxlpejAp6wU
IQzAm5oghSHKTmzBAZudnVoGjQquXTloV8+gyRDAB6uTEdVpiBNzowB2c6jR
XpzQNRPJ430j5vMcv8Gh61qjh9AJnvdaa0E0Ob8jmEenD1UjWhOw6zT0mAcp
snvyFI85/AlJU3cXH0AQi89VptU1Igj+HWZo2yWEyFgm3r/Id7XCFljY9Ir1
GpOd8VRwFoYj7RmXIVxQW8szOQ2cUfv3LeQu5+f9s2fDSVx4za6q2y0PGM5y
+mxH80/Rfp7MHeF88VTI8xBvjHGV5SETXqyNiTih4leIiw/shJlvnEtYzmx2
XIgkE0lnmPhmalIcMNBtRH9ugqDTsmcpYdZnlw4KdKzuWYRPcLeG1XfxqwVK
G18g+hPitt98x1GVQ+WaLMNEBQHueFnFKNbJcQfyC8FOvNcL0r0DjL0muncA
FkolANbcpng7v/xX59ZCzpv+NKaMIp55b+bCkXG2sDApt/gimnrOmW8a8yp5
VlWeTeoSqLx8zTHe6O651yDiCVkOfO4myN8L00RyA9o56rr2MYBxaDb7QFzQ
fRzZKwF+BYCg4mX6ehgEgSYJ8Jdba/w74FOq6GHdilvyye5yHLMe+bTXtKse
TjV5cM/URS+HkdmHewzg2m6VYRtKuhHApEQUGZEWpQJE8HIEbcH8ejroPyn6
8b2nGmiwONMzXEUN0XEmhn9E3sYL6yDojF75KFi96PahDvAJjqqILAPDY3fQ
g3L1oRq31hlGDDO4VW4b/+3oJh7eu0YSudbp+Ovqe4rRbnpUvjrt/H7ElpAP
Pqi2qIcGov3Kt5scUzY8HwvhUsEvOWhm/UtYnwpZtTedabYxfxq9QG/8q8fn
BM7wvQ7RHCPRL7CJxWiIHuVta5aM32HEhsf8kh0JY4tY78F1xb+A3RaoOa83
jjd9Rl7qPgdNAzfxXk5XDqaBYBOLQMRwJCVSkUOpwfA/q70ZyiIzWVaoqVxq
7rP3P/81v1a6GTZy0YCOvzID6wIcNwpFs7kxQ1ShCCTfSYcsboHnHR5LTn2S
zhTMO+7WLl5xbWAbpj1Hk3l4Fcy3OqI+btgBglcsGa9s+O2uQv76Q2ZITEgh
YDAJtlw7IIIfE5Bdfvroo4AkcvUYdUfKKLEnsO81zV4J4b9TEgYckLyzgzIz
dVPXMAS6BSdoVN/OxumIwUZNYSuV6LwZiMyJJli038BE+aU7LjHCbUl++QTO
XcsXfbGD6TbP9N9rrs1SGmTCIli6Sq6SpOEeDNe6OFAgBAKP5d3tBwpnk6Pt
zhKgLHgF15sMl3OTPPGjqbbg5D87M+pkpztSNY30GJ0TTqaAMDxYV02a4H2x
bvH3sCGlhC10mp4ko1T24zPJG2/RYv3uAVhOl7oRFl5Trw8LTe9ge+lJW8Y7
mtmH7J2iWThIq7DicDwKzre+iI0ufuvgdJYFtSydAV8/QiGrhFJwUeymJq/R
E3rUpOylvO+DpM6yKpBu9oSPS7/fLtGxczm4dRXCJDLvLxo9CLx5ZzIUlafl
VnxpegOVVUNjyb6V/95EiLlbh9Lc8Ci2mP6yG++LHL64OFCxa0/dno0ThdMi
oEyNIx70kz8AZfYi+BFDPe5YkqkK0ciIfIP13P32qQ0eHvqEsMjH1AaN0E+L
u7ACkQfH6CFDoYNkeuHsw00tuU/VlWaJjSA/S1KmzXOjFldUxgmQDnSCtJTY
YHxP51oE+xVhvf7MMuOx8yUGgfF30NNw6ElLI7wdzXi442k6bW4KcxnJAYHD
dCJFcIz81vm8FFMdIhpRDiMdQY7BUD359I4RUlUUnE8Cjgb+hqHwYNIo/xwJ
/hHX5e9tfybcgdM+PAzSZvPbvfCJCXrPtb3hwOeCiYjnbQxR0EJN8ipjAlkh
3KshP3fvlPV7jfIYbR8QR/P6xgWQTClQVJnKkKntK36ZGC7VgC4J2V1COFuc
X+7Lyaobx8F3oHecDn/9sPShYY/9EqUeztGy5KAbsXo6ZkixZrigYVRQP+9i
Y78pcgaPbOEpAP61ppii7uWw+k9DFlaVVLVD0r9J31QNlI4I2JJUJvKqEdZI
8OwbCR5qSu62wcJwb74MdW/5DHGktP+dHR8M5gf0RlQYU5EyZRCOURJQ62jN
k+VTHvxj7jeh1TpC95gxWTwEcpU90iaAfKfrA86Gru6Fu0xLRF29Cf7E6Dnq
t/s3Ei1tEVhV8lHpsBp6V1D3C3qZkKqlDwk0HsCgm2jxNyiW7YP1u3NtYJt+
R371mbtdDQaHR4FjpqBOxNkgSRi5yNsG7n1qOv8r10RZW6oZ5qko/na7EMLr
NsQbukzZjKfEuzUjg6LyrL7BQXHqmHnpf9lux0d+6fsEIHqCSpRqIksw+Zyk
Rw7zW3XZ/Ig3/UFFmWY9hFQbiTPs7yIXY2HNXY2Sv35ZdBnbJS11rbnOv6zt
HuiiXvnumpFcTSIxq8o2JNquODZhYLWdIx0xKFE8REMkwvDwTKZ4ch+Dav91
eiVFq+6OgeXRJftPRdJbYY0+7mZgpf8EKcfjZxdhjDn9753j3VNH9NnXX0tp
t8yofUkFQgA6n4IzwV8bgMC4KlM3a+HCMtVCXgHSd2xeuLrzyu3eUHklo7YF
N+7e4swaWMaRQJDx4DrLf7D7GnDe+lSZGEfMmeaYkpvKHJHUUIRkqwx0axy8
Cb8jXzWYx9wL/pqyQWkSagVmsny7RPuYFkrR2JKCaPfc5/YgaIzKydMQPetj
hMqemp5ZtM5ZiXlBCiHgHx71JnbWURlS/vN+eBEvYaKBCzB+cZoyHQAGrO9K
vzie1gppZBL/4X1uZg0Gd4cQrmsZyksi1kNY0T9roqQJErI6u7q7oHMe1dpd
c7gModOU0+PoK+GacGaFUvbq9o4sfUQdBmJ+aclIdRJje7lO6YCielGZI0aL
VmSErL0chcxsLi7B3CsFzGTIuW9pkYmQsMn4Hvcv2MeXHP6KeqAJpuS0wts+
rgZ7W25ysTr5PEytMKNH4Tmjz2beIHoE3OX8lRFon4hXe2tYT4vFQaHvYR4G
aGURg6m1UjKkwSH1b42IeiFql7OT8O5vIbxR63KZBeiMfUoYk+mesel7ghjJ
AHd1FL/eQ9dux0CPCGroT6cPHkOAh0owsNesgwJrafp25D6u/uEfDIRqxSTo
dFMy1DmtST603vPdjxeBNyv8Oc1zD26cbKcMZEE67c7C5UkZtpES9KPwLrBM
Qi4MG+sW6seRgywgPLq9tAWfZ23yhfSk5xWTSsMkZyNmyNzl4LTOkkjfER5J
x5WOVqxB23jXjgErLHAlS7t23uwr8RF7Lm6lErFJGoUww/A10kkXsrncq2C9
Fg0DIhnbuSx+fB3Mlyx3ZB7MujnIW4MXekFc4BlX28D9kSXW3IapEmtnFi9z
f21XvMY79Kih/Tcq53IuAgH3yRO6xbEh61a1k4b0O5Szx6ukUA47gndgc72K
Mz9hjK5HO0ReJcDInMJ/kPM4Tw3yuLnn8IsG8RjezobVFP/1Zc9xxC9DNwwG
u5tjZGKb07CjlxkFIJcIcKNGYpXClZrGQLMgx8NZRy10F9HlRchLBkwekVS4
CYdBrFSKY8ZdmTsh3qe7GcH15EFqCD2Tn5xoxBNdStHJ3lO+AvbS2lm0xhK/
/rkxhQlCUC2oCdUO6ZvUR88knJl7JeqZ8n708XjdT224Sv05qEowZS7ryKgz
sOICBWTZDCotozC0UtAkweWrMysb3x0OPn7mnKqFD6yaVc9SrnPLn6Ppo+wb
a9LIFVqgiQTwtAHCTbiQCvmZS1flehI60966EGvHelJG9F+vOwVAhmBsGo+y
n5bBiHJTF2mPG15avMUsKOghqcJnz2PxBD3FsiDBkZeYvXyxulLv/L+9wJl0
AbaroFayxGguUq6+rQG9cMlil8YTo4zffLt8WsBoFfiXYxauEBc+01GhbI0W
fwwL/WE0VZN882h0pA/YXZ8XDkPdz3CuaB7oJizoFfG07iZwIbedLRHWvQ6t
9wdgYyBDS6F1CEQPJTmPBJ9OxFZlHuvh1HX+ltvd7upCt3TMgeht5pxZvMYD
DlEUi3AOzIbwYX7PLpJwAbGqsMWM6RctiQ1tenco7g/J2YUkpVX/i0JDa9sL
9dHtKBJGhDr7QC0Dn6zMDX5eI2CNDnK/LFtmq3pS/V30itJA1iIHLVbXPsBr
cEoOXduzT7WIFdHy6NYmBjGrCFVlyDpROBxAKW73KvY1B5VgBEeibuXd7Iom
hUkTuV+ZL7feX3uF0xjTjp//mSkC1LnEsP61BGqBZHVBU/EPBRWQV6q6Cc6j
Hq+oF9NoY+3bnguRqsJky7MvdoHo+SI6s2Ay9D23NjUmZL+dAKqzM+C7/WEQ
ptsK6JreeH9E+gPGAgvAx9Wnp+D8Hsoo2azbrFSbt7jQ5iCAMDeyjua2reDn
FREEBw3zxatkZSXNyHmwmSHsq6NvpwH+qV0XzGRc+fIGBJOvhyuN9AigPhfp
6zdcvKRF7o8CVu6I6SzY9T3T8HpD9iJDtg4gYRkwhvAqBXpLPkiN6xLrez8n
ez0x7EpQ3uUEX7ioFEYzt0O5v6uJi8GMWIfjYny5gnd0LpMRckbWdaQVb6L/
h3KJDBMID4m2owhzB+u2TVkR5EiQRm7QAo787loVWEqU3d8x/EJNr7ExMbia
f3PGjmjREvMGNSohtFY8gHH2skWBYv1JSjdslBFGkxsCQ6Q/OYkXEF8O7uBo
Vyo5RTffdyhZarX1zIRI4jJMlGp7uSD3CAA1pJsoT7gyEg4S7Q66TW2Tfseu
crxFn5WJCPvtfLSzAMFIVu4N3Zb6IJ6I6INQ3R0yg1EXHY/HqzjFIi54SQZN
aYWbTiOm+4Jn/aN2P3jvK018LpYFLYAyE1MQC3gpWcg/PrSF8KHjgwgBrl6E
+VWwmr5LliforETZ/mcX0Yu6BPmx84/E7iT3+S6jaDFFKNJ5FrzHyaVoiQyn
abnDWysuGIDOfYLKnEMM/PU7wmfveFYQ44D3zWGFxakVdzQ+IA5YAMtg0FnD
N3n0rAOdAi8Zt9iclYLy/y/9qUZdKUTsxnHKa+4UOeffvgS/JHnUCLbGZZfD
Q6LBsIsTeBCBRCQwVf//VV4t+KL0Nb81f36J4URTKpdjOTVb3viAOqmNnl/m
RZ/5WETzOT3V00frIlZjXigLV6z3uAtGPH/adpHP4Ulq9/I0reLe/TG/um5L
6rKJYje/QxiT/rrjSx5G92a2+sNcukJoTwn5w++t64I/NuvFeMr2jR1AaskI
N7rSlBX1Qr0Rl9cpvqZPeRt/GuCsN3QJKkiHFt/+Zr/1uQZ+vWwUS8BF/TZn
hIYFof9miVjcTFf1ZMttHoxrVMqdqhwRB+YqJsjceNaCMlxxEGfT6RBL62je
aB/c5yDIIa9bQCdKD6+zzSD+MiTtzxCCTMY0Vj6flYhzJZz2KodmfQTk6op9
yblg5ZHXOAen2/YN3hj2bV9uATdngLvk8V294tZYeSnge3ZFwg2Fx6KjVDgH
HKKmSPHjHOI9luQBRLnsOqVKca+kd1TJjW0NrD23HHjhtWbOrsc5RqqIpNuf
d5IGQSiyXxffuPDpjq8l8CHpkoZaypGAITFtCRx+ADrSxdPXr+NcnyZnLdxB
oL7GPhcn/nWdhcFLGBruqUWwm7rs2a03t6HxB1nuo5Qh/5mZbcIrtrcBnq5O
uGsfK1sHMLMVgPv9Du+JlvJnmBgDGhnp7G9lLHF+ovsjWe9nJxj9aPXWALro
YEMARW+iw0An3u3/mecR13CstZQYfmcwk1zWJ9UcDbu4mrWQaalHWdyCiCHl
IR4QvtMi1YYuvJYE50lZRd6eLXNlXwqaJSToTPzHJnsNF2abUFp2kw6RoiwB
HPxuJjEsZh8N8jvJsF/L3WKb994ROeLqSrw+kLw2ZYFiSwNtluhPaXg7gLVZ
6mWq1nqt97nu98qkyz6EJuSBRdO0jveha0tbyAh8ovQBef6QrBENheb33NK5
MaoJQGExASZH/b1o4+FHqWCdVnKT5k87KOEKG6k2PqnhFHH1ueyD8TMratRh
5QAO1QwUGs9M7cJZrhj00+Ihhad+wwNf3E97x4tcas4PRr6J5QxdHRnHVFjw
Y6J1WF+Drbk8lqasOibNesiBV9jcOuhsjL6S00RP+MSYcPExZV14iUBG0Tqd
+0Ns7e63uz9V7rG/cT2bmr4d7rzAFABZK8NGqk5imSGcXeHvSYMQS9QfbRgO
q824QIGvlHy/+ipkxHtcBDg+ZDnhCRoCARMpaxX7zpwl73v5p5FbG61+HmI1
PRfWdnp4KOBr/yxFpjGGsU5Yr6337TKiPr2/RRbSMVmGgElYqmJ/FIfVStJd
vn+0NkbYUYiUYkd7lgwoCDIDI7u0P48Q/pK8kWeoiZ/e2ypenpGcKn0zmJOG
i7fYrRnEyP96MChmiuoZF6sYW8T5+FU6isVjzYB8cd4nHOZCkV5rhSGtg7fE
ChznHxkIYWmScoCPOS5riAasDpB42OZYq9qrLCx2VF0U3PIS8YzSZG4qQmxX
L9zN0wXUPN1IFTo5yNfNTmbFFWYOdQpkhFcifC4CWMlWaRFoSnJV0pJLREZc
c7ULtShz5TPrksj4Qx4YQQMCGdzvG9oYd10OckKsh/KB1pS70EALcaImb0Gm
NsspycCNrsFwtud4XcvwozmtpJLnvb0JtfpJ2pMaMt+5MTuIvcA7ZnpzNLXp
natbvV+llcfMXPeoWXgdIYWtq3WsHgFiFpbY+yEMUBpnpuRBYwW+ojgWlP9p
6LylRShBIrBPMBMHWQY66NNt+ZQdwJbi1KE/PHjf8OnZsVoDJbwxYBDUF1rZ
usk4R13RQYjfpd1qWpWrTRjCs/MQMRsSwSF6YUVgUaE9l7KG/cZK3YcQfFSu
VPjDu+ThD1RyaGyr3KXsX+4B2nkzbEGelIzVH8YTcU8ISEp2a9pJkasD4uoP
Xt5Z0XO7cW0hWFUR57dRg00e9lzzEUK929Zdu0fPNji01mUFSlLhFaEWh9Wa
33aIDZ8fPz/UX+2Yg9ZgaZr9jFDFyQuqlNIXfGieAHZYekTVtWzo5kpp6xqa
hDleyVsnTvn9CttmFw+PrwyFB/SKaFUkK1yVA8FS1ikwQwPISYEjeC4idA7h
qYD3g6vmlapCUmm/xPd2ddFlXlcQocBdz4NFs2aYkVTNAZNgmvtBAAnkclMs
f0eCXiIO3QYC1ZK1FrVuvwY2VpOqIl6iRt/aac4YMfmqCh3DktS5y3e1Vnh6
jfI7vISfx1lZARX+Zz1+gpXtgclhan6wS+FE+0RdmJ7bf8ENeCYdYltVBjDf
PArlxyfEVBTTgW1GhlN0H8bcMK7P7RyCHum+K1zVcxwPB0GXjv8xe9veXDHU
dR698j83SZU/1XgskzbTGkv3JykLAEyZA6+1ILDC26SAkru+0r5ml97NEuca
od7vWGtmEcELqTg1zsE3uK/wSzkgO1yc3UMi7F/XmL/Tr3o2UmAyyCvC3mz5
Tv7Hqc1zAOVyCiWLGM/rVJ7dORLbBk5+6WA7fUyHvhHnlzCBwBgMtIoomgtf
DW9AR55w8kYvzbp8kGJlTU2Jil40Cqf0A/ySMJzYhORdJLzUFERUG9SQ1Mn5
LxMXh5ohvhEj7KXLMJEZEtfO9WYCgMTQ1xb4j820NLfqIvF6fllK56t7lipy
ZkDLdTU6a57jlXF+/PgvuypZvrYw3xJ2z/OSK9825wKCl2qKFyocJNchA0Ju
Y5l1t+6ThPQCKiVoJPCVrgkovs8GFdFczrCo7tRpXtCEpxm8GmIMEkiM+VvE
vJyocSvpk1m8ovxX1wpiWhE2feHyCOUQTydhVdZCDTIvVjfVgIHfy4FvoTTT
z2eU1faWDGyOlLp87Czn6JQOZHE2q5YqGByB1lu8XVFZddw/GNNXq2kaBDpd
LeKGpZn0BpNroFhUG9Yreq2z+qrpqt3XImXPoagwPeGaLkKSwsg7HQpBBB1m
kVL2W7noLBczDVvYvYWpF1GlYRnK9wePbkMXRtH+TXViJaMFF1nBBSCLO+sK
nGyVR6LN3D1MJe2uimzQUAQfGbhsOdpVmEyVfcF4A/7I7/MWbiyktPQWQrE4
FYWuRF0cUZX6ZqryvhqOmQO5hOsBQLAPjucV43qhoKbyH40awo2Kzt+r78vr
GuybRkfCiQURHXq4vjHZdms4VCCP6uVS4T/8V5Egkg3j06e2c0h3136DHEyp
XOq5ZJtEdpZdqvZWk+Joi98gsrVrdrmVe4zeDWptp7y1+eQSqM4wGdLCe5NO
FK33e/9GGMAcXmOsYwXsKJ8UIox2rotvqzMMRAIGkdC+fX62l5SqGEsIyaaC
PowrTmY8qRCfwzY0jdqzQdl3GomoktFmAwkz3DHuIPfWr2NbQp+AuVtRLHQK
8+uxRfymXTiJqOS0I7SuN9jbneXiOxiA+bovWesDyOLqCKfw2mH8SxTGgfEl
p1JeHhR8qRMIf0XlUAWfWcyKxt520/9O8ZuVY5b4KsiBsUp6pAO7/BCPb7j8
3Hebe96PV4h86uVnGoSbc8JafxR+I084fPMVg0WFTiJ+U+q9kt4GGvmJ3I9e
F3xfaVzlCUbSz4Hs7qlVNNplKscfJx+ADKuJ6CeYtHAe5faaBqn7WkuIi+hu
v61754k5D4hJH0TZCBfAEPUj1On9gGuiKAFZhDKhx7EWPQ1KYwj4E7iklsB3
ZcFDx1xD1cWBirKYBgMN2k+y/EJ0oERoY+yTIvp7mMsbQ1KOofMlZr8hMEv4
rklzAPqKFoMzRYN8fP3JMmkxxxjPsSjA5DJPXJ2ODVs1ThxFRjLsoYlV+pFe
HGJKEngCVqIlC4CctHmpCuoRT4Ikk5IJCTzFwOaJ93nfXUXLZ4AVAYtLKMyX
inlcD6P4cx99uUv43zlcPU0XMBEILv/SLLjp2uBLl/mEN8cTEi56BlanKmMz
9QS6jeJopmMYqxQ33IgkX4Un9eDIfyE0Yg5278t7ypOwA2A1+gS7HkJGNdw+
nuROo/WdmxgI1dy4TaMtCLxIWixxCvRZFMBZskWBPBlwW1ySEd+cYEjwF5jV
kWWbW/Z91SnA0o43kk5q4a1LO23QIsZGvhAtPPqIimQ4F1GXItCMr6dmKJoq
1qpHAj24sN1Fp3g8x5bO57U6iW0HsaZLC3NIsp5CwDYdR4XwcEivRLcz6a/E
Fe5WCiVjST+QOdo3EJ0h6gO9caTStFpCvtSVIEj827RYV63KrQdUDoJW64aK
d31I6dXIndCPWdG4+gk9Sub0yWaVngQCcg6cicdPEzgIOQQuO9yrz5K52hUE
M0XNzSHJA4C1NjD1M3i8p7OboLTC+fyK/EYo+SuI9MEilJnoO88E9JluFFPl
m8sfWhIWV9rFvNc25E0Sx91aAH5brtms1gepMAn1XGLLAP/3Yd2EYOv879mh
Fb7UwWgflqPiKeJ5BjAhw4RjFC0qLBPs2RBCEEv5B3Ow5v4Y5z1kCY8u1cI7
n3B0iJQHELGZLRyIALqzteyZErxHeilV8kQMixymyQym+zMT557u9GR35zcD
D8O+4g5yAQuK2tW8AQ2g1devVEFWYG3htmpz+7JQM/mn7RqIl6mh+sQNuX2b
eH5NkngTI0yT3B3PnfmTBWRd7x4yRmBWvG/b6fLzS0AjL7c/x8emr2YE78w+
TPF1VuqsOMN/BN4IsIBA17tmXIN4ofeNrIhFr/wtb+p1jWbtmhQ/fRObWDZt
gsec5laz4XBm/8I37cyL/lTmBGkBJuXxh3gMKyD1Ag7dWzT64iG3Wj7rLanO
I44cEkRsr1HCRcPcVCAk5kchZv/VNPP0JX3IXtQPezmlwm+4KaKA95WsS9yD
W3H8rmZuvjfF/GgdxpZKS39mVV0YmtlgwBN62sOdl5iNQcPj+2+fSsVcJBOs
zPD1RfJnG8X+N2yEJgo+NBch/Db07x6qyx2NbKSQDXHmHa+uwCHDsESQYqHX
sJHAg6Nh3i9r4abVzH03G+hEv5LDbFuNzG5mK68j1+wWOrhV8TaJoYXMmSgw
nSZaRpGgN2tJKP5oFnCCCOP3xhz//mFl8s7FQw9SJ0/Iy9zyABzYBiVXX1Qp
XRUdNcBvgnSgmo5ESkIpQUOscz55+t5gcX2rmWVATelXSIHWZTUV8OVIOURk
rlHcqIiMDI6tBQy1LnaZlsTlmhs3NbZsCPydwhM9EaUbojoJQ+Hksiv8WLTJ
6nI6fQNwnASQi5jpM1TQSBxBy3iCM4yN00r2CGDgpRzTjAA5jZ2t62RyT944
cR8HUrMLweVIF47+Q1Bs1Umz5mqumH/OXJk23qbRqDfkJKHVLjNuJ3IQYtTd
yNF7CBxCOqgYEMAe5g0ASeAYn7qG9FmhnR+GbunPopAa7Xa2RSJF2RXFyRun
X7Vv7J2LK7e4kb9g/7pt6y7D9eAqo0jLpY0ZoKBzb20MkpM1DaGVY2lHJ17e
3jtIYFpvInEGjdantzX1etveydu2Hy6rcjrLDNyftt0h1jrKuxvoZ20s95++
KQFa2cUYwxS+Zst7slJlmlFg8nnkhyRS0eXyhxnIcmUm4gdrsju8HQcfvvxT
OOgvcCGzBTOqHgKC5MlAg2cJOSGOw1/ubROmlv1oELor06yuUNewuo7IdExd
HKIWZjnsBct+mbg4Nz6yu+3K8wds6aFs5HX1tWeqLDpd9XyjbeOfJhscJYXk
AyJRIlPvQWFPSRriRcRdyPUUEGaEupYlUaUMgpc7vAJPNXtWdTahqH341Rpe
BtZfogdfndiPiGEvuy0e9lE8gSyD3CE/7BJ44T1q4vxvCgD6z4ITbCV1V2Db
9iAAtS9fQQxs55JNq34gcFXRG6eg7mqE/Vpa5ZrXj5MterWPqj+nIz4uO5Z0
vy89tec4JsjIWPXD/kgLPufmOyudIowSrGCbhVWC+gdFCiWZOsli+C7zgyRO
RmWau1jIyqgrWCUFQOhhDG3aMRUkK5Mn7HEsSKM0sFGxcwzHT4WraxfhwO1Q
sdwgyXMBP3mF8LEZIlZXJuliTCT/wavcSm3kE0NVtZ5uVIv6tXdUgNyF8nV0
4Z/0Xw/AFB1VV1J0ddipD6pQ3v/4dLto10SR6eU0o1XkG3E0Ngm81z4wX/N9
AruEV8g/c4Za4IUgS28QK+6aeXnlAQbfDw2XB3juYtILuH0FTBhV6IjAsJw6
jbsWqK72l2cTXIyB/YDTP9PorHmXSpK4Q/CNeVGoexSlIdM+q99bwdxq1P/c
/YNfpXB4QzM21CKYkEZCyl+F03FSc3vny1ISTfxxRj12hyNwKUrRpH4LFv8k
jzklZZF30XhHgRePgl/qp6aEUidfkoVCP/awSA8XCyiItyYWBkP3W/Byzulj
jrrmRzBHZDBHE3Fm/RvBMUPQewx+Igldh5Xcoj/WZPIjfItKt2QEEi/Bkp3Z
IRuj+lfSYC0zzFvVZKEKACi/zeLJ0JKsyihhgmrf5fQVdC2kk0ZzwuCABz8S
eHxUexNbyR19RHJw57FrumQMmNrbH2HYz2BAS4D9ozjh7XaPQfMQ8sGTrynE
pndRk1/Kgj70t4BRk5p9u/NKFgxacsBa5GEMBUII5UIGwxbfw3rhYapcvgn5
h6EKes5UO+ezJHpWu0TNbsn+N3cJQZy4pZ7UefjeKbFN+wHGiwcWQjkgq+qw
tEN1nO/46U6NbSf8WqJ7Yy3Buk+6Qw5eS0rlG0wi0jGyy6ZyS4H5YatWA5CM
bOjeuvUcxAUBWMqtqC0vLdoWbFOwZmFnXLm6jWV+LoD36csN5/WuC3aGXDtz
1awkOUJRKkyzupjw1+xWVffgxbSzL0ugvtxqz3uGh0GfPRwK150ZvwE6kQ84
0ivzczVZ9hczCbR6SnSO2fs4O1bjBrV/dVYzrI3J2x0KOIzJBKNEozrpXupE
BNFwhwfq/CwCeGOBsGoTlzxy3poI+S2CwQubEa8n4dV2ZAUwv45gv7CzbzJC
mDhBbOs/bNk0tAfIVfXH1S+wM8nvKSgr5gDLRKNeLxdVvXwUOsVRkXZ4TyR2
EDM3V7Jd+jG3q5+XrPzdVpZzP7AzOpbCnxVXzk2H5U1W8+cUOqjBJEcqHKUJ
osS1LjxKDENy+7EYuMYBLgbQLDbLtvXw0oRc5U4kc1oIDHVmsLV+VjbomEMC
tvZj3FWzBtyFo/i0B3+E/oGUYNF8OZYWV1f4L2gIfPCNThjmj0iBtunmSYvb
zkGjlawkRmS40rqkgHH79uJ6cfLbe8lMVjxCK0C960acFsLbooKaB07E2RBl
YX3tGka/TOwQoeor3toVBDap3PGhVv9tAHto02JWe7Z7ua4iW8S+4BoA1A56
+Ades1kn3irAUXzQ6H2pemGPEur6O8ONI+Vq5LXHlVIWEpsOW3ERKCS6nC7u
zbatr1lh0gi78vuZYF/AqZnFUbyNsYF9m4bi93ZWGpovequTk9dvYzdNx57P
1kDk1WlaMeFoPhShlvY0DqcyVCAZ6hygN9znMLP+pxJbzH2LPllBcmjL+kTi
bIuvHv8+FLeeUFOy0IqjfUUaCAddco/EcepTY0F0Fd98t2CkLe6oDEIbzUFi
tDycyj1oe5JiaYkz60wsRfYp1JIHeYacTy/j5qYQkzi9PFA1b2SK9EinVefj
hiyGqUyT2fZmN6BoGBTBt8GnVeb7X8ZL8hyCBkP7RN99NwTkEplUAwpQHSMR
1s6DNoq8EPR43Z472wZx0qYaHl7kDg6IZ/FLoQddaVyEm/oNWoKGvAx3NnVI
t3N6Tm7vZ5gqY0N+BBThAAntQKaPxb77taXV8eLIcIRUxFs2DCt9UydwcCRO
mZKe3N1LchSdYYsDRMG9iOQMz7bNgVTYup3mzMN/nyIO8rJaX8ByzXlLkbtD
+++2aryT1uPb+wPxV9vaSxAFAPAy/HzFOy+gyjOBTZmrvtTEF74yHynD0zpd
CEtLBEdrr6iNqF9DF9917X2KOgSG1phfWQgEysQbJsWNbZ6AqhJ5XW1E1mj+
hR76my4lzt6z0jfNpwzHwD+xjQOQfeFMpDvtDfP+3WJxgzPl3jZ1r5rfML4e
BdVkzwvBjQiL82Sbq42nkfx2aouJMR10A7dUqE5+KdFsOINRknSXfeai2K7v
SK4qQ3dIa9lYrz6sECcHH3HbTYABHL3TBugQB3C9iJfn4nMTNrEQjoObgVFt
TYZk8m2QRmj/9whKKPkbPZHMEDH10dif97neU884EWCgJgnGqS8xFpmr4+2a
oLahbUQOlKS7MRdBS58lDqiL9R0EQgQOIWJtA0lhaQaAbF6UEvv8dybcKXGm
ZiZQPh0d+K/42XkSxCXFQVvxB9FPvBLG7qa8Up6xuB4caHxU9KBskmcUpYrp
J+rECRrw2JcaTr80fiymEpaaaluTbiQdZCvUC0hf1kBycgqvaCdOOiEbCwXb
b1iociQwNyTnWvLNtsuNOPFPYwJQy+N3cGHR/ucltXzojrfp46K7yyAAo+Ek
8Baz/pHeYHOPYS9drt2+zRzjI1w3rC2mbEOLYiaP1QuM9uJlUG+EAoisQ1Ht
vlRjlqyYKHscDqAHjxrF6jlNtESGijBijRH0UTfdNk+cxTpeBbEE+bbnX7QP
ZF0D1zkY3vRlzbCbSTG6t+wkGDI0q0ZQ4CCqwtfMubmT7MGdiD7uKVwNInZ3
fwwSaipPS25CevWU7koYkNTUJG+S/MVPhIBXaIH8Wvcc7keA8OddpKEkifzg
yYkcXoRvTVWNHvsZGq0zWRt57FQ7stLMnKyOwFAhr2jXEKwol5FO3VpDMuHZ
gJgd0TbF0iVHBNcwkKMzm/fhIpVB1edalkOt2ZhVIKMvsTeD86hOL72Aq5ZJ
N0cCfQB3LWBM31gsV6rd19qLU4P1VCxCBa7torXSux7HgevYnDVVVjGtzTuJ
k+D2ZqUan50ez/ZWszhgRX5B3GDQnJIBbJYVrFeVH1mAB6iSctv3hb84vtSp
wpI+MXGAO3VnlqWoLQPg1Bv4tAzLFuti5FTfuH73+oNhNagMcijpfeJ6KnRn
ZHPhHxlJNFPY2HuVPdVkdJBpO0dfcnJ0ch4eBIx/u5l6nDdHuSzDspa0sUVT
2uAyEgp7LwDN4Z+a0W5N4cLuwNRdjc39wmUgvoT6opjyDOjyXYR/xSl3gx4L
xAb3YFHApWFgoleBp492RDOnlqBZzsLhY6sgjKoaf6TnVmH15druwspdesNV
qbhCygpBMqtLvlD8waax8L1wByPSdmgL0pKp9iTkZjDoZWGtN9o/MX+yoKSE
K+dN4IYVbxV06ZI/RqU9Bqm+OGqMyT5A4uVNeCAiOmbWimVQ4vxjDcwWOGxW
YgZPbiZWl8QCX4H3+4qosE2V0LrX9YN9xgWfYn7v7sz78kNiXsr9f7gjg54q
nPqRwwEtK7eznPrB7if4qVHwlY8qPnUkv+okg7F9x0mrTb95LmEb2jSIfSX6
+E4hD8WBNQmaMSiEb/pu2t8EQ0Zcsm5w3gj+imrePSR36EVYWpbsmyS0Dk0B
TLUKPlo1JQnaKtllVsBqyKHxlU4j3EC8D2R7MxBTXuoLMa+PVpT1g+niVDRX
lmlQZh8jjZoWqTkzodwKX91F/Qd60rjiCjIauWxuja50Y1jsvUhRE2hzWF7M
kqfsgcfDEjOXi7tO2BMDUNe4k1EhgKIszALzMNqE+5dNOAn/vndd/e3X1tWk
04rXN9PtcQ4geH6aZbhfB5a52yGcDORVS7Wv4Inf5Yd8jEDu9L+LtW0N7iAg
BZ/3FYxpnYBCM6sHUhvhY39m5CmscP5XQjuF1Iux0CdsBhD6nGJ+gxTDco+a
1rR9w54AWuHwebSXruVBOQfKCJ+fJtrOZS08pfz/JMoFl875Pw7X51CI5HCP
Ekkqsd+YXn0qyCF4bOdo8yTF4ykpB1QK8JCOhXfUJqJVmNLERHYmWoUtu8K1
VFMR6zu/WV8IN4A3VL/7DYj4zshAcHdyWIXi048A+BsiVIjlDZaH4tM0DlIN
qY0AsaIKTv+BY2G5hI+Xj5a9//XdBmUxdYsZLy0YQLz8wVZCvr4BFN2673Q8
fyMKvyqVD5rpv4Cassjs5BfhoHyv90ex3XUNkorcV3Qu2p1HhGCRbfU6DP4+
cVQKwAr4RPz6LAW2WFC6KEKEcpuf9HcX3oDh1Ie69C/XUjSWoDAIFWEFFztr
zGtTCUjlMhep9RUg/GkbjEuYG2ZALNQU+fYh7qE2FUYeJFOZDNsli499pJM+
w5Eouwf/3EyPtc2vAHj9tzkxv46jh6AKPkoS9Q+3mNEfBsn8bRDuuBFV6dcG
wSyzt5q1TfGU/aBlrW1l00eQUKsfaKd9XBFI7HOiEpK+nqZiVE8v1uxkIrD5
Ufju5YAGNw+d4mdEN88LTe/2IDNBEIPeZYmKfZYkkyb4LreAJY4IeYo1vuQr
LKNV8LLhFV39lapuk16FRD6HCJXSX2CmzOaAyQEDAwrD52/dNVYXnM+JDfk5
Vw2Jia0rZATZb3jXiCbwu+yTeAeK09oWUQOkhcSFi7I2WDT6mGv9S1serpET
NeEBKGV6l9EnTIxrYfQeYq0HImicMtqExk5a0GSXzgIkJf2zdry1X/r2PCZx
yQGc8TC9eEojFGYH4d/MmOVMlLkkP2I/b/wLHs4bZq/x17HQuzLcykXwueYz
lfFN5loYTaonMkQZcLrbQVimz2QIndMNgcgV26uUJNFE27xGtl2yVHTPIdQ9
SyU47t4901Hc7RHIl0W1BJgwRXWSrL5W3GT3maKhdgR/7gSVFGgXyRGMmI69
vExTkXy5QClS+6m7HgyFhCWdYggi/QZmT4uTyyM0h5J7yYv5NQHet72J/tep
FBkYL5lvT38x0HIqFyegL0V1wIb0aahHD/n61AOp/Msn7BfK+LSGZyI0pnto
LaVgjnRHaxwsIMURMHdCwXwfWhRkvAu6j/kj2dRON4E3+dso4g7g+IIqdzLN
W0sNX5UdQv5CUc/iV/VcVEKaOT+/SDa4ztel0UCHnTmM9T1YGyzmMD5NPC8S
p08YVzQNpAiYujOUj7a5eifGikTgpXxo4V7KSlouk96c5vbQR9xmjLQnl75x
69tjordXoV+pQ1MN5fW0zl0HDByoMb7wB/hJ5SybCRJJOm/i87C3HdYtJStq
51uDoaqN+4DTNaz5jKUumTP46v28mM75ThIhLujuYF5ia6kUFcdnS3MZUNXu
gtc0Ll8YVBarDqVvsXEvKwMdjUw1yLUHVy+3nnt96zngYOeQUUTl2Bf/4Eqz
UMb0VDpLhm9oc//v0/9O9qEjdFw5F6F9B+HFEpweiyAas4QkR0NvFV/VOPgD
7J6qm/j7+oqEwRNk33sJHsICqvXH4tPrQKR6IeHHl+P9WULqp2qgZLGzfW7d
vyt/ieYQvky4V7Us7eFrW/+oKkPqBlNRO4+Mlzey+ihwCA8qBKngO+RFcJzZ
MeEFxO6opLG2vat6+HF7Hgi4ekBN76LPbrJRbeaT7dA7r7ZPpCQO3JudX1+k
+yMEJr53AxA8y9VeKuJSLQNuy0J4/AePm8QRWqZTUcsoD+GT0VqWRUYFMHrg
FghBFpt2aqL4hMQGuPRBuQrufHEja9Mh21NL53YZYdrcH4KPjy80qwI95EjX
GUj3Ufa55Ecu/JYwsgTZQ7JPq83v1URnk4R2ChK7IkHRSCk6XSbIfe0n2qed
u2ZUpO0VFGiY9ROR2xhZzUHFL4IAsuGCyU9H5BmfWXDrHm4GaVVJQ5XjJbfP
TpNLFKqhsBc8+Wq08kOPyfezuuzJlw9H8e0JPM1M8AbWVhoA3/1OKdpJNRBH
eXI7+FgN/LFm1mUjtINUeB9i8aVRcDmRAL2JByRxNLm7LCGMuPDiqi09XZMF
InmyZP/PP6D9SwX+GOiIb3ZmvRM5WYgD9tzNcmXFKJwOuRCCHiO2UHFqa5RA
Ts8a9ZdT8zS+Nm34hGNJRCWntNJbQAaMF9dGAXFEZYsAK5r1TB3YGkzz/69Q
VGUwu+/6sg1Lz/jNqlUkfLPbxaxXXWF2tILtp5VPZeqz7K9Ri6jIN8b2FYdK
3kTbSOeV3b0AFtMmhXvOe+SVbX8y65SPZp/arwtcj8REEyrL1xQIFccXDkT2
4H1flY2xbwUTBfSANIo8NBq+2DmRac3oMXlcbxS4UI0a6ZAFgOfd8BYwj/9z
iJ6zsbbY3Ha9G8hCA7aYMlrBvf7nSasYrK5uRDoZ/Xag9a5UFdx2OQVapk0N
NXGUgQZc25ouTZ3XUAxCyUPbUTgzy5s0Mdp6V4LVjJYYV4pi7r1vVHST49eG
JaY6iS1AQyulqGBuHri48WNcP7GQ2/eT4+x3XG9YuLZXhMGuqKvIFvV6KofX
oHchAGkncJlKkLoKE7uOAtjjWmvMT8L039wGd6Ks/2GyCeJYy76X9m/SeKH9
7JelX4zyLBNC8nytdO1DuLEpj4RwK5/aykij5doAbEiPg60zXf0RwlfUSKyO
fxLfBlolm4Ipi2dY+Zg//T9Bu9Lo9NntYH9FGGOXNhTOHBuxalQ+ItDTbxgP
UocYD1gz14yLQ+Bn17R0vMwFVClrenamCqGn2gTPGLAF7b4VA/lz2s4Ln67m
YwlbP9I56+55TJEZKC4v1GXSixUnAyP3JcMkGxt1vf13WlkmC2UasGugayG7
dVCynFEhFsMdSbxeGq9/EfZi9DGkmE+l3Z2IW39G01F48qFZNBKid/EqLGhV
063TARuT/6w6deeDn0KwwFdBgQDb8sqkfwJgCEqzYkQUz856RccW+uBBzXWG
bzBkwYSsd6908ckNm/CUtjHxN2Ps2XtG+wOwsDzKxVwGEvlHS+fOwfL6zffc
XGKqVUAOst4k71BV86MYuIMH2YDGbrUG4Yje9f5TfJTQY8mSzd4gdIks52B3
tc5DJEK5ujvpM5B4y/y+YpVT3s5LA3K4xkbE10SWZf5Vp3AMIcv6hESw6T+h
BGYlRHEMIjvl4ow8Kl9g/sdAiiHib535Mj7i6nzEcmFjhADfWys+Sx3A3N4W
UM1/XK4ke/tel+ARe6JYSc+DUbpi6mH+pEMJMKiWdPXIq4Ib5HG/a1+1HGSM
Xk7uIe9oFU5SkR5LZVDfUWsDDX5sX2xtzsSKas3okEXy9ybWnE5Al4Ru7tYR
MLtncmnfCjyecJwZDXqNrPC24xfOvl483/A5YpqoDlMyD/tKX43Ayb+6gnnW
Bsa03x40tXYGRNWbuEq97yazwZRLFYTRoquDqtgo1OuudDCq1+ucL0b31Z0d
EB9zlZNOUlJme3kk1OWztIPuQv5MHVf5DGveNKGyQpmGpCP7jnTcBCAm/7Il
9Geri26bWe5W8kG0UfzFfm6AR08pZXywNJC2c5bOsr2xhbhYJj3LEXvkiJp1
vkdeIpifecHK+GsRcdHl4R1KzJrXfZF9ORmPETq4Eo4KT0j2vu6yYgP8fbmo
NAT4DR6+AnA6wsotnesYhP1/NNnkCSx2SEVQUvgvSQOkMGXIEzfjtg2Fb6Tb
igaWtFc/Std4n9cRFJI1KpvP6m8Q1L3zurkyIl13JiUWcWNETvicTusiY3xl
SJQAdyz88PTz2UxtvZ3q9BFXkOed3/rL6wgMu+qrxruKkk5STKO74cllALmT
Ed+C9d8QWx/ogKOg0RV8i5WS2MUUIkd8aDh5ddBach4u0dMnxWG/3J98+jSR
bkiLXUxGSMCnKO+iiV8Rg5BKh46F502vMwpR1mkX9SKMQ6Tt/6E8wCe0fOpm
Eu48psFA6NsRDw9VcxtUXal7FTEwmVBSvGdZBp1R4jGYEeDEZIyIZrEyjREl
8DFhtRq8gqxzsD029i1sRUVea8hbseLai3ZsUXEacxStD9gMuck/k7v6jmG5
S3cqdhLUXWo3lAFmEvTqCzVSVf1sMDytuCaLfdlzkxYPvgWAdpjrKsTgiytB
Nf4Z3093HvWzNmtTqbWuIZ5uMoE92ZtaOjcMHpWyRdqlUyfPfMS6VbCZeCYK
K7SZYrn/Y0t4ameVA2xjJ3Q9AnXe3jb/ptcdoT7DEFFfok30V9B3HhpLY917
4RtAeZ7gyFBfoZzJwiBsjHaHULK0JaSADgXEyxkjC5+2sni80ZC98JWEQQEb
wKbPtP32kZGL0AJ++DJ3s+Iwq682VVnV1VzdbuRpPZ0VELMAQ/W/ByhQ4jhS
8ZqBtLCw0hPAiVHgzCG5xwhZ7baEIbkJgyAsGfuySHTmRVlNpxEsvgu0sVv+
rMxkFcPPmj5ts9apFBbFvyR168TNA1ejfrz9n6vZrbGSLngyvfvk0yx7ZqxV
5ehjDgRAt1gYIKHseoAl65BLqGAGoQX++p7PvNfQpA5OFYvJ4AM7izplcpO5
h2CH7kK6mueJHQ98PX318MBwZEyW3qw33QhuuOjbLKkk7FI0TtdSF2FubJ1e
YcHyxMF/rq3Y7z3SVO6yf3G3VwYKUXV9Y46qGkfZ3SkSDwYPXF/ooWMNSjNX
9Gj06xgGWeyNt2syz8HpM5YqROLHoc7Y52TmsZLerEQOlFFsTeYou2S3vvGI
qO7gYa5Lzy3FBA90nKJ4k8S7yIvPBqUo5jfY1wMNsy9L3xImU7RHTblWPwTH
dWWxrqlyEHPre3DEeOQQIaNc6T5uk6KxSUCvVrPuxfAlNecdCygS5VpruWOL
vBsRndFzJV6MoJjpHtwnxzX7FYizccnPFt58Gnb53bQ4dvIVlD2xAGr7A18N
RTwZVyj5Od+R+QVoD5seCSUcMGqU4ade6NQazrjHw3MKhSLQDIuvcyZPoWdA
lbvELQQuaT20TtHNtsGEf1H7DXQyXXqRtfla/CTeK18a1uvJioRZ2sQeV1HW
67zCYgFDT8l5CLvDAr2QwxKgUzTXSyGd3KMSH1KlNOUhYiu5OyZH9xXpn8qk
Jo3OkoJltJmwZVwVnnVQs93Is5q4/BkDosbmXZOz6C4wXcrHI84ZddeY2hyb
KDW60amNIEtstq2A7FFmlKcpIKMvXoRnR9tBLB0CLYwwXT0dSVc9LPVhd8zd
mZmLUoiT0Blbd+iRCH+xSCq8mPs2HFog8XHVqGVZGUPUBtnk3/AJP07XHc14
+gdDw5zpA6ea1rQDbbqUpTJG/K6ks+xxMytFOl67YLlk37V8Bk/+qrF6CXKn
Brue3mYlT5eKCYWKPqoHf7Z74ixXOTXPXxg3zRWQvY94X5m4uSwnhyPryvvc
XkL4Q29lBjYo1G4rECK2hFPb0v2xqa4XoJ2aq9etvG9osjIaRKOPgK3yoTjy
XTpzJdcBdJ18toLk+SLRjouSQ7Ak/pFzt0fjpiubGKG9fdkdwPflCuB0jtDV
3WADf1bh5AMHaki+ed0hLw8rhXRsocfu52k1ULRjt2DzdgIADcF8uYLVzJeN
M7TLEupPbqW2OWn1VsmedxPhWXuhSwyQahm80Pu2XTaPEFAJ80euVbI2/51N
CbDB3UQzbdwd4CgfbgqwjD2BkPomcuFEiNP1pg5NVTJGv7SPGA5ALe7GKzF2
Mu+WyBrqt1vkqpe+q8+Q4daDnIYUlwnhuNmQT+tgpAHBzJPl2Tgr1dEv6nlI
cRqf+jRPEC9LUQppT/X7EYpAsgDogrnOGOiqbi5m/OaobeQp1PSlMmmVnuyN
LxyMB2GzvcvqmEe+K7AA5ppbYi5N/15mTKbPZUexfql7vOSuzBvuAre6QzAd
ajas4o3+fB00FnOLZJQHgmpy+5eQ5ROSWBS6b8Gjkdj2Xjyuztc+mjs+g0aB
WphHYKyh4qwOmgAj46EonkMli2W0QdfedNTcMyaxyxVTo7B61xBGh/xEj8PI
Ko9airhqOrnRMmCaFb4j3ua6rZRAgXXb5ybs9bf7wOvsCc2z9fUoTkdsbjK4
qjJkpgYKsScmkP7s7KW/t79n2tFVh/aHeF6EZCbzJnNHv21WNqkHPsE4hcOc
p5Hp9unUPn4QFp2ijEQCxPRBIcIVdOUp9ObMXSE1GrgoqRio0CAIQtHfwfgL
z99WIuJR/qtwGXJ2uM0ABBBrSY5xZ86HLWIj29zMxrA+sXhya5qt0FFFQiu6
A5bhBV5ZO6F1CV2HtVhttGRIvQ4iyNtsjM2jlS6SP6eyEQHNe0h/JB8E01Qe
MpOQXt19uzTxXYwoCD2/1Fhxa/RiuH066Jcj6LJbU6BulOzDvk+0p2N1t6z9
mKtravdjcCDwd1f0A8WILskggGKT9HxCSxk6+MZbqiYv0r/e0wUauq2IShGp
ziRN2uG5IUiNsNRJiD0Qy1mOcdlSfLNDe/a7XGV+tdBVsG3CONlhqqoqlC14
eVuDe8sS4DKdBCLxDJ7xm4q6/RjhIcoYJenaJVmeT+Yfeau/kOhK0OBBvpGZ
RGbVYxsyzEDdEPvpkra5FtBh/KchHDUxza/VqxSMY15Fq3gnZaZDejYpIOJ2
q3w8GC6117XLL8B1oaW/zpfI3mNyNy3MKTSqzxGNY9LCJ+HbuCjuIQcal6aQ
ItG7Wng9DfGiv22gAeS/e3m81Qv80WsNmRfbktJ/OXMGj0KCZUaFxsAtHrzv
tYg22/6EpDcuuKoJdmqFnUU9f5WNeaAB+gBSzKd7NyAh0qfiOz6IE+vXSv3D
Y75+i+Bcx2+0KDfTZm+zWNZvJzYYfjQnxKp4nsyhb9bZyjq1FuWc4ECnE4qz
vi+2EESiXhCBis5V9dLXH9YeqqUPWhXyzoTmJAMbouq74KwFKCB47kqm5BE+
Bnx2klSWbm2MbBd6eDesPfzLc0VwOlPTYbKVvQ6cbsCLFtSTvk4lZ2llYRnk
XoLzdU/XGWHHqOTBeg5/tc3U86/sWSvMvFOwX/PCKh/rgUmUm31+Y2jfRpIq
+Sj4Zsx3G+v1fCbVYSP/sqOBehG5BDhZW7lTS9E9j9VHH3Umv/Lnpxts62Nx
MAQaufbU1wNOwsbIp7fvXtCr1tgcVrCgKriJKeGY5LNnIT0ncLGtZR5SWi2g
Y4czlU8tUtjWA8Xs0lzKI64s2sWoidk+aEzckThU8DhKTEk7XohrtO7aBoSc
bKzhJ0d9nzP7XT+NL7xLt73f+/Vcl6jCBXDL3BLKDMlFQ48S9PzgdECVCJe4
dLZu0eb+W7/1Tio3EkYZjBQRcURbK3JnE0mcw5O6rhdzhc/zCy1Jn/CYu15L
03TphN8psQf/JdRMiijvspa/rTRQPc7yw9E/2wDCMcnm3bU21eHLmPYzcTuU
8YDsuqdEW4TJZRtssts8Jwdii8jP1jIKqaIuEzZItkhBUf4wys29YZCcHaq1
+7yAxzfX2Y4r/HRkA81rKtJmPQuMbbfTTaIFn/8X8GO/2C/Z09b/Rwg7VCeB
ekqC05rcMCeT/SQpS7n9AWS/qq0r8GLkvHu1NimsT0Ms4fRYnR76g4A65mnz
QfAjanK6p1Lxha9nZJACKIvrDNNTfj3fy+hGKdBJczBHM0mPgNB2wmA957W5
CgLoLDkYei2w3imD94MEXKQ13Bk3L8tVebtFKSECqCIuoGabCKg50PFnyjb+
zEsYrVbK7MrS6kVyJphWxRIUMKFTh/3CFGUvDRnsBA2EYhisb1zCSIckT255
uTI3g1ML9G0gREG3hZASVCTgVXXUyMHno4LQHeJ5LhedN4ctHagjsS/hpdjK
+K67FKCOTUeeR9gRz280hNG+hdOIUWFAsRZ8o892nkiFqu9gLw7duTcS6zw1
0zdSeAcvfauGpO2hQ87IXuscuALIttPYcQepkpNCTOaWeybZBtg7CrZ1yi2K
52ux6xDNwChx03WH8lb2ZA6bdDQvOjJHExM8tAN8DkodP2f7cMUQsYQPfbbc
P/2HhbYEROC+pTSLTAWoHanHR0D8RszxS4ut/m0uzX3rWM5KFE4SdsT+fYbT
6zjHUbt2YDWvGFscKwyjqeKEYnZDFEDzrMS8qTaU6AtB3cARFPwDRQPKEoZG
TyGzN8tZk4JhioWziBHO/gFKNb/+meG6+ASMk2gwPTLpShI0bNz++HpcIeLj
u7oYzGZTt04CWUd6MPkZV2RjeIligxt7COKIu9qlisBdiGXesNgp0/BPRZxu
9knKzcksM34E5e8yKdBJQVLNR1SuWRGnhGpKRsiLa5URFABbe4M73EC6KIOG
dR6yqQG7HTKGfWQFMFKUnXBkA+NcLv0wrlAMeQOyZJ23UaqvbzRcraIFa9Ko
bypCjMbzc8u/9QC74Ox+cZrQv8AVH3nDB9Akffh3b4oFwLdp02AGGQdKxLtQ
YaBI90wkXyqrM+0KN6sU/J1B6THo1NtdQ85huirbDUifMzF3IE8jL1cHHN3W
/PBRPNmSoIHaInQjwTdK7dUdUgy4ZdCpzuhCBxRPkUG7By8aAwOL4hSVHO4I
tQyXdiBliFdGrKlDO45k95fvdK+5ZhP07FMDVgCdddKIYc/UhcY0nz9JWUBj
J+rfDV1DNAOcoI8A/ZTS8thupMrv4XlqkD9Gui9wYicZFq5Nu5dRAmq0MATT
4jVUMy7RtnrXm4SVYL5WDWSol/oQMRUuSRdB3Bol+6f+FsGRLsLxHdTE5BFX
etGFe2dkk7VEkojI1rlvJOFD2B/ImctOvrGNH9KGU8ahLA+PCS76StN5rM2I
LVq8PAHLF+QARXnoki9OmufvNIMPQh5pqZrJ1CwGgtBtG4uxwsO7//UGAYVw
XVFM2chhPpNCTC4jPdpgNWcADg2hCShzDjHqCOAjNGDlw0o7T7tFYjpiCYfQ
A5RpQYs6Q5ufpLlDyRF0wH5jseEZjb5/18WJoFyaQoJrlBtI5qiq+E/Qe2in
X0B6UMGrmZEZtZC2EHq42C+AWe3JhBFIZFa5prGJVFa184A8Wuy+OwWDuhMu
zfRqhJ08IvZ8O0QLvtoE1P3OR9cBGT6QBj8uCqwTY3BDdFL/JlX8oCoJOwTP
dSyLN+sAryJqXVMz5tm0SZVUs6I1wvSxCk1Y6i+hT1M2KDMTfC6cYBVc+0oD
60QGQlCWRNAX4Hyjm2TXRIC37dDNKDlbn33a9Cxu7cmSopB5IfoO7jfy1hrt
hHmOm4PaYWgVB/LXkD/ruca7fOr53n9O+8YFCoPGoa14HHWh4l55eQEjed48
Hk6E9VtYLzbh+XRIK2LTDmovnspfs/sRodYJsI6pv858cryQX7VDfa75oQPi
vkbq8DKn2wWrombe7NuAvqnPB1fJ6DT1155ZcOfZKCOcd4Pu1hBJD1in4Bnb
F4WP9Yh8pGLEuu01RqBnPjMLaSZtMJn3NBchqa1InGH6xs4CJFAJc9EvKt21
nXRsY5LhVPbD5ppguLaQFb+z2bssa8YYT8rUG3r/XwgiYDw4Q75iUSRrj15Z
9ahzo78xHvvT66FPjvPU5zJD9K2yRzfzgk/WL/sYTkaOuvYYUjGNIacjK+Ov
ajPjL32idUSKGMI4dTUvTFRVE3C35SBxXxU47mAmIdyU0OVG65PySw05mnVq
VPI/DoSOb/4F6kiZ0c/MBcZRW2UvL2a4GirNvAXdk92SwNkC9vwaCu8O6wUR
h4yKRAe7OENWbEqHyw08jPiDUv+3feh2Wo6brxNiuF/DRlOm5lqUMQ7zXC7I
SMybDtf2D5aah0dzGDBPN3gFDAKMLTmwyFvjdgANl3n90ox7lainMPN3zAf9
hgKnyTH4kzgrrDG0YejGC+jw1rom43XhDvnsGNea5euQHMsg9MU3I6wxYeos
bFBb6NF9MCusff+yJG6lHlV5nKZ0zU+UgjF/l5DPVlP0oNWK0aJc19IqK5C6
SPiV4Z2iCJGnjwzQr61lGtS3SP2XbJ0LjMRxq9fZEz4THeD9xI0q4umz2Jue
uert3TtMDRHHbBsn3JbmaauWDGLvkUrJf6+x3Gf3aN62J8mvCCEog3mlTNpp
KJ/lDXmHKdd8cfpA2/vwHkXTldmV6Fb10pA9z9T17DumQLDz8bAI44DrR7ps
4loPhfmUravCo4OrGNGwoF0ynJe+EQVCR710rp1Co+yYwdaifNXgCaCSnh2X
PYSf/IqxFkWCMCpVvz2uIvJrUaYNZHpQCA1mSBE2yyh2oKk01mIVsXOxCovO
+hfq9r+818n96xKyFhPWyszhmMxSxev/MOX3iliN0J/UGw9GL7tSKL7zSGYv
LBMR4PcbsfHbwkHmDMfDbkGa0Al8vJJxLqhWxUPSjAs+LWqlCERd33eM4gb7
7xA4wZJXt3nAt2i/R2+M3j2fLqY62sBIy8bhZuz4rWOG402CvpHXohdj6Ata
L3kvYORNt9Y8D5k4v6LaGCJIzV6UFAvEOQ4Ee9+UpfXQfdvvHzjjsAP9rE5g
4M6r5cTqwZIqy5PInd7ZklxY0c0KIspsM1n//HnFEFUbeVhHv+kxkyTwu5jF
TX/AqRoEt5lTM4aJEHWK1llLS3WaKBU78yT8KDrHz1pmMhTvwWqqGXgxWP9F
fHOYnITc1HPQr9NGAQtyeXFjaYjoaevTNeG84/LnkoMSNr21LyTmpcuSwAIS
kkzjF2SobYqLev05sCPr830Xl7oJb4UMW02twt8n4fOLEiOHUplm8/UC5uVr
v4qEOPcd05vgGO6KEgnz21YLAcZ32nWBqwIKmJMyP0rDDxb3Al+YD/RF0GdF
GUieLvKKtp6hD5vj0DG00ku1rUJukFVchO5TMtBIsuuPoJSJsWoxfmzqV3ZV
YcQ2KtfHo7VY7kabhEKYOko6JMwn34hnDAaGsIOll7xT/IirPklJqkV2OfZP
1gM4eIEHW3rZrdeys7bQ/UuUW/ZyeDcXLmZypY28QKTGGP1D6rHaoIS5wzQG
O40URuhPZG+c18Ys2jE23ukIZaW9eCVObHVuHMKPksaCHW9bjJNYC+41afm4
ShJ2LEdkXJOu/FQIkTWCKt0UJyQgOKvKief8b02ia0P/omv2SjdRe5rjSLxs
F/fZT2BiBvxXKIviiY7B5dmRZpBW+zssAbAMmeXwJmvoHMnWHpxJ2XvFrv2N
/+C2fRpiq2INkoU4v4C+mHBptnx9RPDUMBX9e4vjB3PLfoCmVdHcThsYluPs
GzrjOkuwiCrf1ZT9Dr7QDCWyZaXGmM94tAINE+IJg2ors2JkGLaGy4CPV2C+
HFunLy31D2YZL3kgHEdk+T9J8m1w4kWLOVsUWIFBWcLnluZaDWmdUDWG2XDu
tziQF42NYp8pesA+N5IR3CqtV4L9HXyEefn+2hqJuv7iNjjGRTuVBus6nf+c
nJFr1p+pzVYRpn2+w5NJR2XmHfjkGSb+BBVBKp7IuW897BbmMW/feddFjMLQ
IBiWJdcT/zutkE44mPFgLml1cOTXfyqE9Vsjb7IHY3Zx7Ky5aGKbjg+g4w6m
Up1SKEGn0lDu1Bdtv9uQVEMgm/nn9/eSj+grDFAlV0fhTJWDKuOFhs7t1fBJ
YwBURgU0Dj4e6cQFGx1oXcXjHwGD3f1/BP1aABwLCvvuNrR34Ny2JH+eW5ni
1IA12OO6tZGAuvgUugdhHYnU/oiDPggBDV0nykvjthVw26qTrmjeS1m0NhdP
R4f2T+Q14FZGJHeokTdIEQl6OceVPweljgRZKvtobCdQkI21OWS1sK9hEEg+
QuM+dyN0AtVxnLCFkrp7nNhQ0TmwHACTxahcVtSizg59HuKMWormq12Gm3Z7
9EO/hvE3p1orAeY9UZQ34e4D9xANFV72ZYXoKGjWmQp1hG/lrz9Qi2cpkMvN
cGXnRxXLV3dCPFXDPjwwCp+q1CZgsPJ1lCVOR97dzL8+FDwzkkJDd/wbIPIr
CHEy1xQkMjeoY03CxF2UykT1loFXgXTPMfyTIVArMZRdPj9NmDuU81+Ws5bx
l2ATMqO37xdkp6e/lsytjCktvbJgIeqclcnEVQLeOBh3XCmErDSNY4QVC2pE
tGjE3mIGoCquZjsPPu2zuQDo9InOu4n/4T+2fuUGLOk7m7ruunIzKPN2Hdbq
we9YEE2PPblazAi0yu6HfK+YkRMHKuD8F6r9kDkq+2OXU1TubZqwIemZMXzN
tgvzIt1L2NUW8MNAZR1ge/ubf0VaqnnsjmFDUjfKU/1s5Bq4AGCjTn0ubLK/
5pX4i1J3ySibrjdE51CJ4yT0RWEcfpS1XNW/MFW+GdT13SjcNcgD5Y88kl3D
Xkhhhfv3wV4QqMYUi4IPUY1B4+hEneXJqp4Ffr6nkoEi4eiR/uwbPUglbueu
Nl02DWxZuV03SLu63MuQqyIudlCHqZWvgymOtEhDIKHmjHcZimcFYI0qbq1s
ka1ozPT7v5H+9OqZIsnXZ2Tih4aGOnRsPbFj0ba1F8swYjU1efbKOnB+wpF7
vKHPQnuJpXdObfdcqk6F05lORfDVZIyPIUMYMGL6IvIqlzGWH0KcJgqTigdl
i6UKYfFH+r2g+1xDnfmxPXeM9NAQp/qNLCVtgvhRvOEYfe45APvuK8qofKMc
VxqrvlAuWHhO8VHYM0UHAU/qDNwTnwB/rzmNP1fyydhOEa5GQeQOuantvOZo
/nx9BLdDM8HwWk7J2t79XvG7mrIuGmUnfRp0byOMXgbb083P1dxYYSgwrF+F
P/R4xgok5WpfcLJ/gVD++7c/nNwNCfXhP9r0KooqdH3x2+VCIP8YKehp/WmY
LLbDPvg0pfwtows4qbDJ37TZlIVhcnmwYRF8jbeP1zMuT+XWQx3ys69EQcep
tTTKDDBAlqTdkUZtz8fBFhPllWXnvwGALOXD8s+j/cQwqa8NqyxrK30MMQZr
oSgcHcAEgRJCbtsAWwejHhQgCUhSa94JwJuYXMaFkz+wVzsgltdyK4I36QYK
MhnKgjoXP/rYjMqr1tzMwrNhL1sp7zb2V5kwCuRw9YDu32fzO4qgEhJjzSgr
C3ZJXR7R7K7QQaYIPqMYPpCGAIL1Vs/yfBaQZF3H3FBf0tCgfue7h/TteOpL
cfUvJpxvEVpt9vWbvjc/5hxs8qd6WM1aeRU0LCAc0WzA6YvlxqVfNzdEWRto
CuAn4IlpYxl72QGUplwOAymwvvqAFqbQY9s8A0vY8Axyi6WvLWZewPYQ0UL8
PZeUc2c0iqrcJkEsrGLAsgamOkoyRvD9LELJfCNsDCcwPe+IAiEagkawKfP8
6Tfbm1dbknqEIZ+iDintZ0Zi+T/+Qyj0opCQxUYFPYAtLvvsDL/z9NTJsmll
YjFaSDUE4yiOVCaILX3CD+ld2ap5chXXEd7cagO+YIyDGz05H07ST5tAxJCq
KTfNyDYVBqle5oIBp12/4Fh7CHXK0aARHwKZ7GmpOMEagrsLGI57/LOp18rT
QaMkz+u0QVVshbC01Rc3u3eEyloRV9bAw5qBJvEDqtC2kli49r+u+or8lE4e
bUzb3ZUX+5cqNpwjyo4rg8KGZrV+CkJLMfsnIRKom2NfZfYxH4/WyeZEcZzN
vBSQO4fCyq5Y+HX4im/N+Ft7CVkkr2YjplBMztddQWrofQYBdCUWrrWMAaJN
q4CWVOV9k3UZTXaX3AjnVgHhgykXfTW3JkhvrOMX+ADUCHg9olqtpwll1dU2
OCpMCVM6HYs+3gGQaX/u7WbH7woljf12+DvunFDBP7bUb2TUIUeOMAVr+ruw
9BzQKwSaKY9LX5fhIQtcQqd6r35f5o6KQpKybgBiXflJae1i1kNY2i5NatnC
q9FTEm2K+PK0M+H8pLVWxkUGNlZ18rRcUDfHGfUIXYoVm8mB9BMR7lhiwLUq
pCLfWF7y4D4nnaBhoM0Dcp684vEIQyZTsuRiW3KFT7BwC0Zx63Vc5unzf25S
NvdKUKSnfqfNoW0iOVC6M+3XyNfA7n5Et1BQdtgXv6X0nB+dM9GuvtF42IZR
ESicTVCGElGg9ojsG7DqopUFfBB6QTSMg3VPwDz636tktszo7Pl3ob1nq2Eo
6QJeFIsd5EhiD1pgnfpLV8nicZVHQ/W4r36wHDDAfBbDnJIC/qgl+IWWYx6i
n+cR+/SPDikZFrzkHi6OgR/SXeFaUvcLLKNIiXfw97j7zrlQ8SJJM0zTD+ey
X5121ps+Jop9m8PCL04PD1QSaESoprNNw2L+V54ipHRzSSpnZyCXZB9QKQ0w
Wf+XzKCHc3MdQZoIMQ0IBeMA0RAipNTTO7TWo67soNX2HMQcKkBHky4F1JXm
3zQge88IajiJr/W+qtrkKlfCX154F8XfJgmgcSlC+Oe7Uz7eQoa5edVplmgF
5gDR33HwBPRlZp+YyANDnFCN3nGf4Fjpvs17haTVlru01PeWuQHOUqs60BEo
mA91NKazFFBJzf6ggtU1SjTqoN+vIEfN4V6OpdhzU5L7oBcArgU+YFQqKdFO
MNCpkd9cnlmn7VC7Fsrzfm+/eNIQwvK47s/E0Wa5xX7YqP17898HkyHru+D/
/CnQ7iMpu2fUQgD7uDX3GFZU4HL7AjZtHSE4jZk08rnxFHWv2u5maiZ+BW3z
CYmK15uOxJ6qN2cMadG9DDUvfbx7bJO0K03DeRwOEkXy+7+ua/2Q9oNucVbs
3Nz0W1d1oqFBIT3FQmyQyxP9er8Q+t68ox3QgKWWWQa9cpSOKQtU194Xgld/
gT2YDiPCd26WpXbnZEZnxOewGBcBZi6JhpUKHB0ZeWVSN7GOAmIw7bPFYZqU
GdoA97dx8z/exOChaSc6dAlurRBl9pI2ZZn5iNwxqHcMkbBBPPRDOoBJp41B
AT4T0/KkRrYO/2a2lQv6zbHsGGlwgVsfWwiuEqK0kJULs6YH0eqaX85IKzMl
1kkqTFds5uosi1IZYxz7jN2RmbnEbEf1ff0vU+SjZjZAlPIPQbRrYwfaX0Qx
jDmZRNpn6vHAKxmBjSdzzHsNc/lVHjH4CbG5v8GKhVygKdTAP0HdbSjFm3+t
8Y3CNDy0z+gLB1Hx+fThX51AlCy30ZQn/lxjD6cqEkYHDszaAx4w28CUGszu
Hz879nRJUadcoBR29fEFbvL8mLOtZf986iWnsXyCcOsKddWJ1vVCczBgt8XM
rGsDv4Jq5ILAtH2f6HUGdSC8iheTJtew322GJIV7/pBPgUMyWtsQwjL4y1yB
/u1od16NRqCeca0WmQ1mnLy+xfMB2hVzZ8PgKzTKjLpEiNvkJDJ2IelOONPw
nG1uZSmta2ak32Ry4kpSTlCpX2c2MsGC6EE4TX+bdDxx+EY6GxCHDg5A/G0q
hXmfdEoVZtj03FtWPTnf/GyY0+H/liCmPtnNdRRW5AqIPcs3kYArokPpVwFy
cognJ5NEcv5TirzZhF1YrQn/ZloK8GLBjiO/0ULfCa/ee6mQudsWBOfhbxtP
l9Vb82tZSAE+yoBOZs5gkVCtulIRGGP8xwtdoPg8lm8umbjlRjklfo/xdz0c
Uyu1lUXZueoa0q29GZhVcaNKoCm/+2+068HF7PZZBz1UoB4su3WrQo5O1qjF
HC1b7nUN+npwoO6CribX+SFZrIua8vS667anRqdkckf66Tv7ymdfqGKBOCPl
6heFtgO2/HsZrUEIwJy2cxXeui1G/gQo0mMuHJF9eaoACwEgENnhMIOHby2x
oIJ+x0fP2K82wzQc+Hw6wWg82R4Y9QFGPdQU3TAPXP4Qw22m/TtM/sGnxW3Q
Seg7FqKXzhGNXfXbYreubBRnNwbn42Zpw4fH3itYuJ47uTPgTTARJdVGeN59
aWKPI8rFeyVOaiybafkk40BN4ieXGOl6xU4NSlADTBgPRXLUPSCKis8Jvg1z
3Ia2eLleFCHBFFM2UvTvHqdurlwpxAPhElndHwP2ZhKRC7FcitcQMTbulvIy
2FA5GC35Vomcxb/aWgn0QM4QBMO9VO6JGUb0U4oi2AhGxLrJchnG0zmxo1Jd
uMUfLnANL729kHIDTQ3hsXFzSl5q7YjY7B3WBl9p/XxE0vnjxr+KI3khR1VW
AkcgqdsTP7nhLDLrX6W2xxdDxN0pACFoCNGMciH8t60LZINCi7MmzTvHeD4x
wfj49mZZBeTBvzI8Ty/EcCjNxoeLT9tt/PC/uyzyjzWq/GEEvXN26cj17ntU
45nArd1mwYW8B7ugevAUNjSfrvveqQY9GZZzYLVmLMFlYcb8qzwbfooQsoOV
33+hXlNu+/pYzQVVNdrcMXav4z8ZF/gBRdsePlgTClFQoXEJ8vxaIW7iAKdT
DMlFt1yAjSh5AgoYFT3OCOaP/qntC3pD8jex0ai/SUrxHR4BPRmAU3NROtg2
iuQT/A5hzjXKgCsH4liEjZQH3FmsG0WkKOu8N2qk37BVXHRyIjsaAOisLXr3
Pg7nnMIrRdFzFNQY9+Vc61VqFbu0VwCwX+PASJFtK3pjmJE4hIPWYme/TKPL
1OvmfSa0SY4ikLv1WABeh8cap2xkCWLHfImk22CVI+6PtHuWB8wMNM6C6JGB
zpBtBAVRw4JIzOvlNGjCSHtV2rifl0VBHL+imaxM9HOkhcQZdoxsAhwbd2sy
fo7KhFqjd82KvCajekaFYS1eyw4U0XR+hniHZDmftIndMvSd6S1Om5u/iixt
lSF4vWwOqXDWETeq2/1ZNhoK2MBNQdNP7GAlojBnck3Bh6XYOV/fC+BjO1uB
ce2Rww7Gvxl7immR+fTTGW7wFKvv48RsIYbSYJy72xltctchKIAz66jQQLLQ
BKvUbT8oHbbUbQj1prdtEaE//L++IaixnGk1pDyElV3LfsKPSy55QW3pobJw
z9Bd8OYviqE0TdtI/+fu6BPhc/4X4tXSCOtyuQu1Ho8i5XV4r6UEZIfJr9VY
ZgHxCgt8uLBvqKs4VPtPJ1R1BKNxjNjoOelQ8H2RuvqY7HJeB+NtXjURs46j
aH6HMNw8oZ4zvPOoj0eqJ98Rp4tJTYb4QIk1uPGIS/EJBJmw7IjNfmBZoJWP
cvoBwB5Ky11B82SFWr+365CNOgutyp00EOTKKM/DOgy+ryhw/5N+ehW6tO94
loJPY8E/WPb9BYmiAe2xcrmVw2HP9mSGSEJUsR0uvBFUjNOD54KL494Lnin/
Ax3odwV/ixU5801QAH1XhA2aQKxIwHAf66Wj/GGideE4e4Gf0bGYNa2zaJkh
jBLkE5L34YLXYdjqqVKjZu9lEwgCTaI/8KW/rN8yC8yCPyQT33AnaT7i3qkc
GyRqsypZ6gG4kkYF8va1iPOrncYiYmPPhn5G1aYDvP4CC7yxJOz9kimcZvTB
JuQFBUSKu0rM+7a4+JMhFIoq1JPMbYody9gJznP7XKkPfgHC7dINTqO4Tng8
uOxO//pM8N1JYMEHs3UspG933tRMhs7GoFtFU2cAjPGH67FLw88Rsh+N6u0y
deXsjBGw7kaZC7HtzTSv3ud+Z8svw8m0kGBn8mXVha66OY5wqfMbHXiPManD
X5Po3YEj0JydPnscQPqFO3tAQREg8Q/a2/LuTgxaOyryKVrRC4Ghz+jQbG4H
xn+8ZFvN1NSmy66iyXHKqUYQqvJAHxvqO5SFDm0GJMjT2hBiDuGTrQSHFDbN
gS06SxbRdHXQpezbBT4ynq8QHyklRWuaxV5wddTmRd27QRaoqyEXft413Xac
PX7ZIoEckpdCuKIvEdf1klZSLG9M9+TGis7nPrMcj/cGGYrKu0zbvFz4bIYv
JHZUHus/or0dCaUCXAvlLgXslM9kduQq6kqYimGDFSRYA/9NZdI2FPa06/DT
fMI6bkySZvLqYyUsclulPCGk6DvxIXCmgwNZp26sldEXtq9s9VSnp5tDtl37
J3/k1tlf7jtQ469ekLFqxy7qlXO2HUHVlb7I5/3D/SkHLeWJ0poZ7f6F0ap1
zwjL2GX8FK2adWANdidptpXh6Ru6RHFSfSUIv0e3UOd8qhkvRdO4GqbeEf2T
FgHOfPU4b6ruw5fktgDwL87tRLZBRMuZpsdLE5ooJJPjd23iRSFqhmTWFEk7
H5pk51KD9PcMYzhJpHLam/t2nu4hnaLDJS1Juu9pPpk9So03DjAiiSN8hMPl
Uwp1eN2UUziQOsTRM/jSjdGnamrgodmPZ63gLA3He6UESVqd+Ca3BvCFPc+w
jzQgnwO/uHxpS52CMg8zUMFmh2QDjYfEcy+hBG7vbxximSm5mQ8eVpnvbplg
HpBbBtzT+fsQAYikZmOflFMbR5as0DD1B7AgUjc85AzhcKhyZgREsEZWxRQH
XqvmICHXLTtYaCTyXlgl3u2gVeQ1Gaa1mFIOWavzMltJ06cREwXHDqgISJSD
XXUyY7FVjLDwLOyCjDrvQzVncpPVubVtzYKWD/rDIVCHgTxWJkSPbvueX1Lz
/pcrlXb8YEvkt8hVGtFK05/O4c1OkuvDigqoSUyWcb47pKW1jT3+1+xebUMI
yJifxl6X/0vmgFr6XPSffOqfyP46gQOibAK7Z3VBsJUs4tjYXwDglps0iUUV
h5i85U8y9N3Zrf3lmv3bVYHZBqaor6mkotKyFBtr8bPUvWGzyMqRUvvFA4JD
vdm/7/OQdLBEpd6RE3xkFe+UnRQrsMQsUQWnQ8ty/I8algdyhQZd76RCD/FJ
Ig+J0SOHDWuZya7uRBRHiYWmf2k+4K7bo57kQd3wJKi53T3UYZLicPLWGvIS
H2c3sayNGTgQK+GXkh6IelGIGlD6eIeyyDoRXVxpz6kIYEN0pHQXVRBoJpUH
g0VjckVB+4lGmw+63Ym/tXIhfJT5Dif6bKpJbmteZu0HzNZBMNli6iUc7b3s
6dxbgAl/CBdphog+5sJnH3efiWk7wh/tBJivTazfO6mVnz7lNmw7+Sx8Oz4k
skiGR/+EeuTPfwMqJt23EsOlvJAlOtXEvlSQG3fnX4ibA24bbHiKQ7zg94I5
i4LtfZAaseqP1Jv1xVGsyh1Vv7o0WR/Rni7VcuogPSYZmLW7qnsQhbTHKzK6
l4csVzQuUlmFjFPVgC7t2Ev0yHMvd/QVUPw3xP/InNFHG55RUkhSgY+goawn
Ki89obYA35v1f/VzMngUdIdsLFjbhvWzhBBX6GUUjRw9F1ftWSVGwGDQXQMs
NVaIkOc+YEBo+CKD7GdcLXi1REmEWLy/OQAhS6zeKIUR6agmlLkDf1TEDiMa
xRhtdt5INRFOLYSpmRCh3au4oMky/gJ09LFe8criEftT9hJTrxLxjBcda8hW
lxxq0Sok+1IwtOwRMws/VJYaNKDXJTRtTBepiXVaNjdic1BGvWdd7E/g6521
QeZngqS2f6unWL+i82x2cVZ0K1A7VbkFM/4kdGBYgthbBu2ydD8tcvf66qQs
Ki3aVQdmFo+/CQY23CIACP4lgHVoYcBm97o+m6fnFXjNlcVsF5VLvauV7dkK
aO5ODbRHF9ZmNxP+7+VesZRqqqV58kktzNol43Qc/U0tk0eEFwla+Kb6Z1BA
4dJvK2s2fDLXLTmdRckvIK2uE1EZzS3ezQqLDkkkCiy0iO6RIjFr1eW0gbjL
M1cghVmUmgXmkc4KHWt7stY0Kbz3yNqzwBwk11lfBJ758CQp4fghn5QYlNIi
dgVKwXjjZ846ujRFHot8H5O/uu768wdgmxfKz3TpxAvqTzKzs4E9WND4xthR
MNbuKmlidHJ4oQ+0O2if7zpBFD1goz+dO+9Bs6Mid97rLkbh9yJ3zJ8YtyMt
lKDYSMY5mJlsW67u9XnTCqs/JreRSylJoYY5LIrhSq1uNDcA64mOTNNaTEvD
BURtgl8ubw6+tkALkca9Nt4bdRuR+H+1PhQ6uQN1HeccS2WJTXjWAIT5yxwo
cSiZAJPx5bZgKzpyWJPkB1mIVwuCe+jp8cTZWFfjHQMvWfTu2NSF64e3vwj+
uiQ44/SE8Ta2NG2OTvd2hruK5et44YSzODOv9CIimdtsNRCGcjDOuz8zZ0Do
DDpB5yduZNmoSv7L3XmMlXRVLnhcZ2tFumkElGnZHrQCCARSBMRjAt21KpCV
IzChbPxLqEz6nMMIj2AZqdkrF95W3i0UmSBSsUPbFDqEcqlLJIPNyYkNhllV
/UmO4mwUzGeSOrQ9rkAtanoNJtg54tsYis0DXR/c3ccHEreoGpoYgvxLvA1d
QKmA1KOM03ltVBIHRI7DwNQ8yungNvlrfyKmUuMSmiSmBiF1gCEIMfLJItwC
GLv9M7Lso/b2dU+Qffnwm+Kffnvq3bXojD4g4icJj94ZHD8CExbADrGS5Kca
+njWB0sw52R3LR4bVBe2a5ieS2YaRIR++il0xKYLOOJJ/T76UH3z5aNyAwiR
64Yx2dsQejqWU8BXVitw7Orw373AAYOcCpnwYcCvKodutUTRvNielkGfs1Ni
8ZKQ91uwH12uPJfFmP/uwUqspqhpzef64mjnJ5LB8HNyojhwig8vQbpZ6SNU
jTz7gX/PGFHDOGt30yDP/cNWl0NR6I8tM4a5h0lkuNx5hXTp8PvuJt/hn+2h
ARL6caFHfyb7qoBpYi2jWA7RaR+dCBH3g0WXzwGPVjK6es1JoiG1O+Rr7pyG
zf4x4h04KxOlgxK+f3wH9U5HnMWni2Aa0TZoqU1L02MYO9QlMAocAKokADNN
QbKPELLogRw8W9QQ16wyaT/kFsrOjWDh8/RqQLRawNBByXCpR7VSPlFEGK7I
oq6Ys7pA0TmxJR0PTaEOuOiQFIlMX+aNuk37ctNkjrwBLaxYjVvmYDEiLoqm
DuYAQMnBIkpZ2Y7yOxYkQSo5LZ6fw4s5HbW6z8/y9O5w2xJxgLO5XN42PMiU
G/hk2d2YD2ziQDWV4IpzdE6n/Ou7rQCXsmYNet0g2O8Quq3YU2s/xhOzQ5/+
5UCFLro+mn6yfxG10ipGivwYCj4a1gcDZwA+VkWTU/Ks54jA0POnBAi97wmY
q99yX8qNoacPMbVI1+ZJiQVbh4W2ljrzwV5dCb46BZsl7gLeqZck/pXVKzVM
txSOm9xBrmYuiIcWqCrd3DKWeEnX2gtCB0nFC0HIOs0IjnQuADNP9ctyJDGy
zuM73FAioQU80Ao9Q3KLqtYFKvvSwq8oK/ySbBSHBx4omJpBnKUgvCovIS6R
xWutu1hfQCDMKDQ4aa2DQIfoQvNlyVJMLsiWakFpLY6VR4LEgKaEiEoYLRPc
XsM8I3w5nK74RudiXtvXb2v7l4YtMsM1Pe4g8Aw8f70AzQFwv6lEwJ9RXABp
BATBfSFTkoctfpr0/XiPqnxpoR88xTjvZblREzTrlk/5p7RGtHLA0XQrCjNN
K1zAefWL7C1kGGiBwCf97nsQabhsUnp1WjdJmXqKl/Ogd13NmIoaqIylf3aw
UHDVXNEA15xpJ2s/B4ZC7n8eAwZCcA0jEDoqhj4jVWqErPpDndgcgK5igUd3
lCueaNgMaZ+uHJAA+w+AXZemaaFCZ2LnS+WT0IGi38xIIjNFT1f/T4NE2bq/
NKHhwyq9s7qrkx0GvvXmvLIkbeVDBB1PlH/V0TSVLZgfY3hPCDC1y2ltaxZV
PA5TOPFVEmuxgohKnNNN6CBjHXxb8w+VXW8+9nT473xvMkz3iHLvQq59M1Sv
VQBZQxHMIgasMvY+fk5R302N2dcVuw7zfs2XZYpz7eaxYfLjHHi3aTeBXFhF
0y32gqTO5kpuUhpddQH1FW9dqTQ1KPgbEPFYxNeDoTOxoT0AHSt+4sVgIjAn
IvQXlUSaEg7FiaUUK5eMxcnYVuzYYnlLXIjSO+Ysv0162cen8qSUxucMe7hr
Vi9CgbkebO4fxOrT6Fr+xl5six4kCLjicekgEfbpUwcDf952awuQagXH1cdV
JgENc7pwpDxdEUG976AWdpoDii5ndw63YRIxSVBdhso19a7KRsBiCRUyfA7t
g2giga190B4M0nkNSFdIwaz/IG5ATM/F8uIUhisKlZQWNfz/EGnLRYb5m//L
sKu1Zea4z01lbMZgpMwZqj1l2HJMHH7WpFwy35RM5RDogOjud+ePeH7j15ER
tw5TNFnNSroVCQVVEL0nMF/wFuklwqaK9bjLb/H4o9RtAxHqWjjRU1b3y8us
Amj6rfZm9FND43tQSRGF/OfBX9lExfm38qDBvdZuZjHaXYCzpu/qf2JNm19u
9yjlBX/DQVv/fJKeTZNkZq9jl0jJhaYXpxoATnFsWl3/xKyAYNwUEOFKAS23
OtbFxBLDhOIc94ZZoOwDyuvkr2p6WwvkKiuHQbHFSp/cxrOVlGyaRn7Xf8FH
wCPEU3b9lkoP/9zo1o3XqVNjEkE5d87rnYsKvnZeZPzqPbbFyHfxkO12pp8E
PU0B4b1t039tsbgLiAhfCloQPuzKSFzCkSdCH97AEBZ3qUws9EU/gk15COrE
dBabCUXUQYDYT4K97/rSfsp2eJADCypJpZhZwEo44uwQ2+uYfjPvz38Fxy+U
X13CyJ9pdDxdQlw1pgyZHkXu/12zFFFzIxDMYhHxVUDwoYxaBPd1HyCBU4OV
bY4m0fDf75QmSzlQn4yVR0XMHTY+B2RcGwfXhXVKdvFWTWh/p1eYlqU4zd7P
vMDor2NKn+UNRC1tnyQPb2b1ao+VFidFBB+w4tpnL/VjqSMN5w7vmr+BerTS
Okni1gDWO0IvCXmrlwLo6isQXj46gOgjN3m2T8VhI/JiTnQ6Ycl1jWJvseyO
hlKrR5NJOCWInHXCUCTshP5URuufEjIAKvRp1+vgYxknlQcquBMjJN7CRviJ
6lFHCqy7ygWsXvxYlwA8FUjy3lCYFQXjhQbf5z7CQKJeqBxBvkOB3NClnJP9
sIp1aQAP2a7Z5cbU38CAPbMOMuF3f9sr5+H1zIe9tAMRCmm+BdT68ISntZzD
lbn+X/dw0SSXTf9yChcKz+5K13NuvrQiVZ6IyCmgamAFH0MyCN52VQlEmHcM
Db+FgR09l7r50rbFDydftqK3D/Npceg65BDJNLSUrO11I23xjoOLmP7bhAIp
zGol0YZTlSBAAdbh4dljk+qY0R/K7fu3Yrmy+jd/qrmkuWAGukG0O0AJdRxj
AyTqZP9YC4Ixy0eZy0tTkiPO6C58G+BijecYLo/L0V7cdrMUYC6P+aNpl9z0
6A5aiawYof5+hORqds6K44taa27O7fAsxbxzLW2dG1feNpz+BHr0D3r6rus5
V/uJDKEE7A2mIiGo/b3DnTBfuYWkc7mf446f4T7uqLH6/n84yQk/q2E6+kVJ
pGpfVWEr66OM0Vm+cd6SXOlBooDi6CjppYzJzMS0Nl/kFKDbbjlSvSWom4Ib
fUQhBpGyA31l6CzFmPe++SfuGFInZ0it60ngMWa/nu3ZtzJ9xKStHq08z/lf
S+IF1JHdGuexLbJKQ7KDKptvn02IkHWdIo06beoDL7Q8LxFy0ChdHnNyrMcW
tLSfGkHGUYECDOW+ILbNYY/1ICzMchY94/zekmUFrJFiNj5wehaW1Uqst9Ys
iG1AXx5jLj/3Cs9x7EDOBNz9igQN1WGdRBsX55iNcCjPHjeKOxMqCICf0r4m
95HZvKm6ZClMMTEQ4nJOvoQKB67Y5bSEfCC9kPZo10sESKRzfPw39HmM9HCn
KagZoIe52XknMCuWWzGjt6QIXx1LCJ15H8km08kIcNZserVJtIswPt6EgWa+
YC+fbG3q1WziKTDb7eq1q7+07CWwi1jM8CoytefpBBzbNlR/+A+RwizQ/nXN
QgVC3Ab78unG08ClUANN0eIKbd3ZB332GbKg4m6Isp/IuFGTqWH5suExevVy
IoYAcy3Go1SKYv1vwkN+9tcvKu796PKp7BPzyuj6TcMINXpvr/epymrGW+jj
RraFkTs1qoTtO79eOwLhUevrJ8/TIQc+HrWi9XqfZzi6E6WK8sfp/dv5pr07
x4xVn2b8kIDzowAFSltznsPm8vV29W9kofeIsjnhayOW+sbnk7Q0ubmsa0J1
/e3oW6/gxynHKJJ+OgiPIXfY9TgLc4xMyEy8qM3PT4ySuoVkaDtviN1fm8hd
tenh5cephGqSnM2nMmAJBVV/eZaStgHnc3ZUHRwBmM5umklLV6hKvrAQ1fRE
R9QYlaCusPAm0s/HSC6UkGZ1PcJjYaS6kYpMb/yRCMXsKFoIATkKDXw8cuwu
d6/ohBvWqRJan3beLh892nkzxu8k8dPY5qZWrP2W6KtitLcijQtJZQvG6p12
FWNZYA6h8dPFNX+TZsMj3M+EK5UxZCnHkkl+Bws/eMcpsxdPcSkL+QLeCbdT
YJJU8qZJ493++y7PlkFgECHffM8mpztZmDfe2sdUQC25HL2X3BKpoqrJknBj
zggGO7JJ/gGIlYMUgECp23j2L+59FxWtNwgP6yqJCWvJrZEa1LiTmhqw1siU
Lti6IcJSwFGFYWxY8AAza00kvCXdQg4+aND64keTeMOKONH+9Bg/ezLvsfrd
jPaHNPW7nqnENBUyNpFLX6LI1cyUX4jIBcxOytULKU//W1hq/Nfj3lJ014y5
S57kYlaIRGUtrHd0Fo72TXos/UqjlQUaSi/5q4/4sNa1GcFWB2wwLTr3I3kn
hp4CyGrJwXA8hnOW6qQFYpyClMOSCEu05f2BaCJGQLR0x1IOFWOvzoqTPpGz
ahNROSLTckpOZcbn1KFQ09MmWxNyUuTexA1nq9Wf5MyTHSrHC4/7DvRbUFx7
hmaz+Ksy3DlcKbyRoMBsJ+sMOIMIIxdxOttyVVBSleMQOjahGeAGMTe9OLcS
7hrRgUOI3rmNR1UEKc74wCdEEFc7mCySL2GdTXorW3bEHxHe0S7z96mUlJOY
XkzkX8AimVGMTaeQ/SFb7sVxGKkJZN8kDP4hLHniwR/kaLqaF6CAvm9SJ2Z9
BfrClYgBGI4Qzl8rHIr4VzELD49GYpw3/PWQ/DpQuC68A4VxBYaemV/cgLFa
Ag3ImR5inuzzKksBxpcGd78aij3VGQWsgKWdOs6imgHUn/08gitVe+aVN6OO
teGvEOqCDNF46m5w6NnqvSPq65wZHKjD3/K1htfWubWKyc1QtqqIDhDq9/C8
LIE4e4VGE2M6CZtHflaXcaC4JecqUJ3fX7z6rDvDIk6+Vf+XZRCUrrlAEk3u
UADQkIa3PYhZsRwIefLNJO11FCDw5MOMDfWUV2qkcMofjyhVo+f7Ll+GxcSQ
ddryn5Mmmyk80BjIvOMa0OeLmMoxacTehA2xhZRhbZLpY85z5u8A2whmw7ZK
fkJCMgNqg4WALNXq1p0iJbKHNsvGpE4JAhU6wNjbh2kkht7HgaMb1BdRdcOp
oeMBEbDbCrD1/Aj/icEnV4VHB+cA1sOECzy3uYu5QlSZfjnkM+V1PONH+Hv1
huGz5dy/dMkWkUGKYMLYM9/MLyZistTw6PcVE1MCzRhBKeep5mOaclk6OFRm
TzOEb3xiacJr60WI3tNH480/ffSinWOJixPBbXFLq4QFWDB6uDmr/WyrtsVu
oTb4PqZeGyothJSS58QpN9qZMPQV3NczN0VBmeP4UPmcBRDS+LMCRBtwt0kM
PF/e1U1HMD32FSJ/ZWmjHI3g6FEM/RUEU0XkNTktgKABbJwg2Jy2utDC2+iQ
t7TD33DODrrdyl7OyFqMej6KViHpOva1hmQ6+sp95bVigTNTJwzoFADmNVIS
BIk/pvpNlxQy0eTdre/yt2cWq4+9IV+zHMFJpJdahTmlgoONGfRC/wjtHHrr
l5bSFzyFAxhB4QYjKnZWLhdfW5OVpYtfWM1I++vSOnYhkNtSALuKwywo4bYU
wJ1/veQvyTJauBWH1ZpJef3S8aTeq87b3baWvsy9UREAWx3+otD5JaNgvc/S
5HjtET0CmZimn0gBXVHky74eEyOwQ6b9vBJ9+wFYYwhgFv+paB18O08BEcC6
+rGxBXaJev1ZySHpEwplnb/8+5+2JDEPyiIvGWyco7LvsL7Hl0b8CR+pSdUk
cbY9Xrp3biVf2Wr4wbm1uW6vH7WLN7rNr0G4TJigbQv6LK2zbPGZ7T/6aSce
mAvPCoJXRC0iPagD9uHjr0iMisZXQiwt/0s7B/V50ahcWvRL7NMNrzZrX/6F
f9UxwoCyqnjDlCicRZCN6vVgO4Shmd70nhbh1lVZ9mmYPLCQ4HifdmtulJdb
leOiIv3AoeahaTbx5253+r1FxOrpjaDFldJTEsCTKY7XwEZL9KnkOISQZmGJ
ozMyLt3vSz/wmanv1GhCeVWV9qQqsog85Q0h/DFY5kiKSICRHKh0bqSL+7tU
NcqPEyd4/6LC9dqJWF/5zwRMZFMOuCginZo1z0HT4vrPc/LlWseXocOLYGzB
OGyrmC2p36BHtTmEV2qvqWOGEskjmz7vRVDhUSVihu68RwedAHEb10681fOF
se/wK2JBExPHaU4LVhfW26NSyUYwyUABJFpDvWUaOFmRSuuWfGgiK5oFASE+
nHURTeByIQXa6BYFH5zT/TGEi0/wBEKwheDzZU7W8l+vLd7ZvmRHtZCUcJG4
b6yxvV6U5tZh84TiWDhGwinzGkGdyMm1Pc+Lf4Jq0lh0r4rpyddwGK/mWYVd
8twdolQ4gta+Akyc31U0n8ADsbhVR1ihA/ehHBJ5dnwZWCqAZbK2FC9umakh
jCGzz/FjUObXOF5BhUb6zgUUjami/1K5bDbmKkp5lv5WNpl6txECt17lVIlj
0syql3pWR9btTGqvWjhTBIUeURBMSzV20EpSvr7SezGtIeJiGQffU1YQK1nh
Wxb00BOxKLh8YjK4vXzQsr+P+3tlZPacXR0vVu+c7AXG+ghYPMGPhkmt0n8q
HfkyW5TscNoX5AhDaSJ6sHQvNWTKzxiI9NG0E0ms7yGx+oXnFdpGbsA8lStd
HP1lzhijCyuJvdTI3/xZswAXYKN66RlMzIA0HaclkxfKmcftNAo9iacbXUkV
P8SnaaHywU93yRNwb4C+utBgCvEAXuWqM6vmknxGe570LAKph5l7C2C6++kC
tp4IC01JjcGNWqJfBe+CvVWLC5f6ZpWnVckcCB6aib1NAqUzECCUsnaHRCkw
MPa+s31Gy0n1pXJNaVRdJ9rQ785pnFBlnILzektxypk/Y+AY3Zi2e6kUOsp7
Whyrmq/uBISGKViZNrKtp6AkHKa2vWJspN99QGAXu+DLryxsDKLjv3iHRobl
X8bo2tihTJpJ6LOf/dpSLVKT52aoFok1hENY2kejYAMoky7njrMRp5xf8Sl0
VPl+luG/ni+fB+wOykSyKWDbcnqIchxvMkFwGbRusegr1UFeVonz3Say+/XD
uOi+YN9ZL7S5pA/ODSI8ht9I8mrhl98LnXS7/Q2kdMthyndxOd0kMPNKadLu
nJMh73u9r8A0JUEaRA/NLmGZuHn/wo+STEWvxOV4EtmI21LnAficdn2ZTXff
zu8R0aHF1RlCcjbY4nANofBw1jhdCauPcvSoLATiJbKXepAyqBZGkTbz4yme
5ic4jijWUFomC1WPMaV17qgAuBTcXbw9FSCmmQ/MjIYys2sE8K1dbNRR+EwJ
V2gtY7SyR2eN7qf1doCnhg1czi1CYjhb9myVSbVvTlHsIqd44KeihCIbpPuJ
OONwKwM6nC/bDjM7FRqdOVtPLeunl34roZPnz9ejPEL8Wjb2qgk4Pl/FMrlj
YiBTsg1tRJX1pNZm9Yh261pfxY4H7EZJXG95YXX/JK0o+rMjMkb3V7v91gXY
Po6AcY1+QpalbaWt2QFFCRSnhkVwH/vlipE/dIFFlcTKbWJhQVRo5X2WnHq1
TA2j1HwT4AcWzwMs2cmDDdnjfEwdFRjxJxsiCQqo+qMWRWUsnTmU3a/7G3Vd
R6gawjW8gatfPoB2X9CiGr84aG5MV7OgTdKN6f0kyXfPQ/Rbdp0Cjhqhb35k
NVdzBP0y+LnsES1X3g2pkfOIUQrRxsTnn9O4YRotznq/APZ8FBrkAotLaj4Y
I8HdcBIlGwPH5ZFA5ATEMoSlIeM6pePzsMV/yJjTm9jX32LaC3a34N2s2k50
4cIitldnUVKY+DPhfaaGQdAc1meoZ3Ln42LwwGfNnV1Gv9v8JWy+a02QEaZO
YMRQ7UeDRuRkfxQRMJbUH72+uCRJdsONxw5w08Xhp8wh20FWu95PbQVhHd40
k0nG0ToT3Jah2xVAZgkW+N4rfVRDWzo8umC4RX8jJlUSkmL+CrKsSRXSIheA
GvasxSMy/6E6vnw7wmwg15Ako5V900HUAiqa/W5lmNqqXzzq0Ge+JH4m+FvK
kIH0zZD875l2MiW5aGRdds96sFE3p7eVsRuZLaVlkFf7VewfeQ5y0EIWIyBn
cMU/nQqnrutJBP3kxbGQswxRjljr75vpPo5VyXtOBwTaUAVgGds625RjLygA
9MWK5T3OL6EoZy/1pk84yUgMC+S+wTw9BT/g45hxOvq7cD0e0XRFhOwIu4wd
ihp3BkMQwF0xKq1Uv82RHwaGQQE/UwbrwLD+WNIxZlMwRJc2WQ2kBg8/8DMP
dzf5GfSXhCi9mgdYwWTBMnJAdEOXFxa8pkBL1wUvuN5vI6LYHS4D7ub+JtMT
+fJbUi7S3zZIRhv6f3sfHD1HweCzdKq4FKAbbUHZtpSpQnty9araLs8gA75o
QwUYT8bCXjEUgBPC2SBkewrclJR6vb/4MAsghkXcihBesuz1hTOUizbPwhol
4qDXjFPYzKBrtbdGGoQwYrAZHB/pCGX8Qifl/usLchQoxGaddvgBHQvaZDGA
QJNmItP7avvlu5MsulbEB3JcjYCbUTS3DNzI8wtyjs1dDHgOyCtmI4cEOXat
0sMnl9YspOmtDeJL89YGGOk+czKwVinDvhW8jQp/2WJQ7SJnyVcmSF9ivXrn
0z/5ovtqzdJSoFBtEBeXJ9kOb4y/NudYHW+DMlA+WXWOwAKGeJ7ckSj8KlsA
agpu6xX2/uDnMmTzyZR7YQcC6oAvSW4dKEUDpe0W4LzT1PW46v7gExQ1J8bz
SbYClQZ6+aYWDVWt5Es82WakpwkqPZ5hsEuvuv1dOYPsn+AOUDBXZxgmOZx8
ufWKmYnyR+UennAeSBMsGUNtJ17iGw2ULtkT1JP6V7rtJKIbvcOuTSVEZ1mE
2UgxoQRhGIPABIJay61pOB/wdOkwnsJkaeKsn2AIrtZeiIRbZIc+SX8ac5Bz
nJNE4OI5/clSbZ6dUNeeJBm/7or9Z87mdmsp1XjCQuHWltrX/+RHsPgaw5d0
qYgNaXR20NrkCm+VrgFhS9jpRfQFT0t6RVfGbeYHllBqXIP0FZDMkhV7qu6e
ws2FOj7t5YsoPVbKVbuJAjcqGa11qQ5ZF0BdKQqQgPkrAEkJDfDhIVE7GzcW
TjLs8E406IuLZJ3Hk/G9Ad+3hA3XADpENro86t9g+ocEUrY3bhHsYDccmrzQ
CjLbmCWG7obnadPZIaNp+X/m08d1PbStuN/ESpqJM46VI87d2aZ/3TwixgZz
c/g00d/MMtwNYSa88IQpeWTHZutGD7WZNF0fCNlqjbm+ANXgZkhB+/BKGEqE
gqr+i3/RbguXSzO9t3HNM7LWflmCZIfh0QVdY/jZgLsPlWCl6/rZ5ynj25r8
uj+nDbvVtCIUlToQD1Y0UTP4hGh2gDBdJxyK5PoO+xLXvMVTUJcczthF4M+E
Fg/8lhcpKvzBw9joaTT21IYIotgOxBIhe+VI5ujPbg/fGKyf1JtUoa8gpkBX
7TQVgmAKqT8svMigH+wUHm0dRxnplS6Y7NG0YFXl+55Zj+hPJIT514GMW8xI
Rhr8fIq/Y2gjpiWYECmlgd/3WGIK92Zevip5M4mPdzaHwUyE+OfgMXyxY32L
neESmOPi+RlPLsThu0CEJROC5994MDobz0Zr7yodH1chwHmXtJVe/HbEzukA
48lZeLKzlwL7IihQnUrbuHJwTXWnLa45qkIGqqwdWsixE252v2pw1m3mG4fY
mS5HTFPbUagwOi+CQzY/YRk510OXGIYcfsNvpZP1MaqZQKizl6r0I20LqgwM
X+agbsdxfE1XW/nYoHFX0AbazE2MFjaV3HvY7xUrVb3G2qsDM35bchv75SMf
qFRLMZ+WmlM4OZcE9CIGm0MeuUdV891yyUTHr/uRq62DUmJ+A40mBMIPgHPl
+ymg8EJkkP8f4F+owRcRewzbbYs332hT2B0xJlw0cOnOcWCyaj4eF51VJ9hF
W95ldwTlCCOlBmdI7IRR51YJDbJI8IPUjFdUsrDylUlhz/hG6c31t7qdGuV8
8AU4G9UNbMq8G0/tKrBfBVnRLFeswyBNqfEBy9T1oGhLYYY9WmFVmsqPrQse
KlWnagzM3c/JQirWLq8qI2JLwqVdV8XmfAiwf06YZV6MiMls+PWYky+E9BXR
uJnNA3jYGKgqyQOXrhfsGuf4XtO0Fgzg1/OSSBMya2/IMiWKzzzfZPxDuiUo
N3BmXqvCMsynLseBtofhdFOAmT72P/63OILTFFmTs3bDhy/cNZfI4i8EPU/S
M6UOYqGa1vvpM29rOpaNzITY745ZOP1B08MNqDCSs4Sx/FO9vTBgTu478Mc1
OAxAjTXrqEjS54ydfJsIe8FXvv+jGpBbEZGCo7J70WzwcHIbk2Gx3OCcfn1O
wZSu1W4+zAVVlDYICIw8EIfPiNtDMeAsStweVavz6jiQRJH8hnIPUhLMFc69
R1qIRiYm+QaT+n2Ys+ddSJYQP6V5tsN2MIEwerbDUDWFsc8XxIKHWs2GBUSB
6RFdQqwB0lAo2qUYsHm/jWZ3mN6nhYrW81RrqUlmUNVcRxgdqWyZUd/xXKAG
x5r4YIrwLrn7Heao1I/FsEPz9dbwh+oHHLfOVNGD0Sx93E7oUWKG8gOye6Kq
J19SzGfTzFmXnTDV/3fTF4OjmsWO+xLbS/Sgk5q8HEiJ/3UNF9HjINCxrCjS
SdEF3zOmqLmlASvvU7Y3eYhf53WccKTuPzU1Qu+sRqIcU9vldaUciGTUAzpG
1zPq30ynPNALfG+LEK/SK4pbfPqOw4D6pIfsyCMKZkiaHiu7o/0Xi4e7ySCv
Pz5tE6br3NTVmGqTSC+Qcqv8SrrdxBFokkhZH8tTKdr813a/o9oQucirh0NH
cw4agEkmYWV3s+CUuPpFR65OPAIDLiTKnMOjWx7am3P1CwJveffAsKhjMpUC
kDW+zlEM/7SwIlZ8nb0pgvnIlHf70SJ4D/OxfcEHApWKP6qrfj5Bp7pEdzMB
c2r7REQ6cTe+v+wRz72N+T1ykPIM33nR+taIvYMyOZ604UuHrjMLdoSgHry2
+OYjwapPCvOQ29Z56F20UFL+A4/pt+s0a38PIUA36mzYQtE3f+Qp3zcqH7UL
1qsmmD4CYAH8ENaQD0C1KLokVerp/vDMyDoNlpqa771RWzuQwcimXctnPBPd
yFAiHMiKm9hVh4zftnakJO1FE1rkO3HeKN/EnRHUzQ79lxORYmDMQvwy7gsS
fDLkoyFSapgzzCACBFweVaPwluJK4d+4d2OkYbhcpQaJE3I3VBL8NFxM2GFr
/QrLGOhct9h7YV94Jniqzq5XvSE35Ag0owl5jdIHJ6E29COsNGoYgXWG+lo1
Ams969gJyr1o5AfzaVOC6BOG0YO/A7hJJcLQWOlgmhIPbUegcNzOvLP5NPsX
yWZe81qlw74Kg1/VjBTs36liTtlep7yENi5jl85A680y4Gf3ZZJpOK+61oPZ
UeR1co43b7TnoksFJt/pkuaDhvH0iihxtQ7UlS5N134WeqsihHum1O+gjTvl
aUKMYN8e9JvfD9aXO1Ho1pAamF+ufFiQvMJ1u6NGRsEWFs/FyRga5MeNNm1q
4hBM5dFukxyJLY0VWbYsjujaDpwur9l2RmWsVK1YDsmnf2P6eaw6bVgk7bNt
lN/In/SPyUb4IToEaaJCHzCEM+2D2ZqSlG+Km7uyot15nVamGh3xzhdXdETO
wSyBlJea2MatSzlQzom9DZlz/DAhHUX6XuUy+TEFKK0XVAWsjJbBCQmJ0aOl
QxeFotHdGV7JjU6mCqGwPwkWrFiC+VkT4zqkVgXK/wjhqyYJS+oo/gKtiEX6
PK4bLR6uVwxn/HhnM5NItD+wFKWYtEbhEoqrrCt/UawPxOsg/0B9J+fFUbIm
celdLpUqBVcFDEUAU8hyNmVHVDeCoiJsJ3/migoZxLs9HSR+twlsOg+GVbd4
5zwB0q5H+dxw1u7Z4wCkr9rt7hbzj3f5QdyltP+Yx0noDiXqNQ2bnDSn6xk6
BS9RnHAPX9HbcWUwLyn9cLRmjAj+hPIt+wMxLDgS0hFi7HIxyYh2Hch5SmEI
0M1DtUU/ic1sMmuf53Mrp0UO2p4MfOLZTeLBkC66ncsawpBqXLuWEvCS4ZJS
++n8S6l/RZVmu+JSKUi6d2oRINHai7E4KgW79AhUHeD769LU3DQU3KU7xDyI
scvu0C3tdhLv91J3sT6tYNQI2bvC0ar/Bbr7W9eiwLCaLbLT6mbnAM2jqkMX
xj5L6C38tQwrxKBUEVrsVJYdCQGgcYIL4+Lzjs1FSU9SQikhZ70hgpmTaUSk
+xWzPdmeAqYG3//Iro1R6i/myTJzFeAqhSUuyaRh6TdI274BCQyP+DP/PIrY
uM70EB8dgCUqy80nt1d15SCYy4Tqe1XUE7jr6bnf9Mwr9RbP8W6iv2sYeT5T
D/hVPEHgG7bj2gHszRgxsjsnNmtvit+1ehiQ4pzQbhkfP2DqH/QdmRppyG0+
6rUR2OTWqsxUZYSIdszDFHYH+TYV1ASxVgfdUtzqj9lAoYRA4aoJ/gP0s/8K
IebmR2Nb7pXyFUYEgExkE3tYMGRe8jNmaxHe1dnOx3eAijMgEHJr4dYWWOjE
6vUwnTSdaXNUItG88p9kfNdocQkk56GGUXihbo4asN79aJG4JXFKToYDj76A
YiyBuBteYRpiFW85UVab643KOZ284T7wfXbSGopynIhrxXny/BCirH5vmItC
6QDewgMggDwxGgPAvbrVOZp+rGYsb3US1QrZeojWauAiZRbQe4591zK6t5m5
TPqT4TLj2jCyV93cAUnzZ7fYreYxefdTD9YGekx81vP6BVR+ACZcQWrVBBUx
knlKRU5EKhcDbToVgMyuvXM45JexjOFiq8yKGPuedwvqnZhwhKX0j2AigmnD
KKyf0BoDhgnpYNIzpyHlMcVljZbSK8KoYzUb5k5lRLP5cIVqlHQJBmIcIGMK
sOBeEEqy4Hhre4i1LuhVlH/2P7ZHAAnWwGfY30e6pfZzWn6P/P7YqZrUK9+s
+vmVvCZBsl8a5CUHYUrOTqqQrtDRwAcA5Wk+1Ux2IoFaYv/efY5UjOqIMj4N
fKYPHT/8/qpE+d2zTNHOUqlT0UmPrnpcD1VAY0d6d9SzywXDxGszrvDUWLFh
V4AlWIFPkNzi9y4xBD+zmGyge7pL5w8dC0vy7uHOaXg4ByZW/2qZApGLwuAR
PjECYQvK4ZKdFdMI8Gtvno38DCEnvjk1NS0VLfrLpAWObmmhbzPBkLxhzc3y
pIgJwzN0UafgwBbgi9J1Cwt2vbFJtRGwjlLQOK41pz2a/PDtUNvLmWli05kL
6zmjAabTYI2P8qN6sd3t0Vp5zUKVBGdmDAykbBaxrCXHrBcZwBmzGuY/D3nG
aDEIWt0W+ts+PqgSDtObqb4TqjreDcFZ9KhkJ4WEgt63/Umfg2WGaYoQwhOG
BWs+sAEQRSYLUk4g4LT1qUIc7MPETe2Tpmczu3EwH6mbM6hnp78MZkafg7Fs
lDvHFTYO+aUztvYnB2zCPKqraI3/6ruFAcXNJ2VTeNgkCoAhtQOZJ/bnD7qT
eWigZyKeaOO5m4WDFNAi0dtdVnemAzDj7rgfWjVTRa1LcMKwYTrVknG+3w8m
TRk7jLLxERUSuGJWV4Ho25XRj1BQgoSOCC+uo+TNhKPmlu+QpBNAopzgSP4c
BMsHVxjimmkDtrV1S63+UuHTfZPz0YyREQRm09NEZ7ohhW76/BYA2VLFJdXp
6b0kOxCWv41VAkULosV//RnChf03cYyC8vAhi5nvc0pcYTaU/MUX63tvd2sZ
IznVRiWGpAQHgC9RvsdtkSG2omQBxl6FuaOaH/wZYSs9NCM+JtLSv0puf1VB
YPAK95gVgW9362PwRkEkUu3RYOJ7BsWb+QB2+gpb51VkR27bbOJw9Op+V+UM
oefu9/t+HmlR9MfmiN3dC0Jhi9HBMQkk32FDP3/yQUS7O4NwjTkgZMtnqSZi
/KV5ZSPjbhpcs/rFnAw2U9Q7e2csSZB32HfvJD/0Ti/Skdz1AdsmX0rPkXwK
2cqXIN/1GRWUm7Cub84IlNHYKJvBCm/iArfOZoGqyQrN2vFnw3IxP/QRaMmA
4o0OdVEFOQ4ZLfu7X71GaxXzgSR/MVPBeMXLhZHo4kWvqGnWiwbdp2N8XkB3
LslfCAUltId95BgtIdpwLx6F3BefJspaE09m7OJWrCnu/y2EGJHfj/1SrjLm
qWF9O37BOc6A1eEdQvQvgm0+MR4PNW+96+hVvzt7JA19fr/9zvDdUvad3i5P
H8P9u3N3htAxLRB/uYzBjy4ugGCo+DBnSjhjM8dLwNC8MZ/OdgF6A+hBkokH
tdBunS9fA5Ye5nJ+Il/x7eVjvYBt+G34RVoaI/GrRtEki1BsxZmDcQjxWNZt
78zYOre5+o35AY9GCMblehHolK3ZqVbHaIMe9HUBm7ulBJwvvu8aNAgtvLBk
T6vEuDZJlWxvJJtdf9qTFS2zn8cb9VSzDHISBfgnVA6gxCpbd/73cyTFtYCA
Cf1TyAS9u8CQXM2gITRT3NT3FCLYoDPIpcfu0UMjA6KzE3JAt1n8HVFjoVzv
EM0ikXEXl+l5PTlG8EpA9Qp1xuDZrEXAw6vzhBzy1HbsCyNHxP7f47Cgk0AM
K3DOvuRMJSdSi/IrQ+QcK1QDR6nZXE61x/LXuqtlzYjuHxd1oYArCvlQWYwe
YVlQ6raDznTCEoY4KD2mjtHlLlzbQ9GF+G1f7nVUDF0fXGxAWA+JgQf8mi2Y
9tjldw/BJrJJ/fpKtxVU9EjREkZT4rBXyIkxI8qGQf0Ts8RyckerK3wpPxw8
hFLaIZircZ7O0G252MsG4rRqoh7SMIa8NFoAcQjiuF9jdfNZefnrVMRgPq/h
crYh96xow0+jXFHtC1bj5Z9HK2Ai/6b78U9CU2L8JNIPQB3f+FPqYNyEjddt
z7FyfeIsaXfOFSjLlKfXFi/BezcUS247NbQQ1+8NVsBMhb2KNzsNpxKzkrwy
ybhWGbiMu+t3niQHdlqtdu09gcNUSenmO0SNzjTdWmkxN98haVR/fEdfuPtk
gCFgX26B2InEbpmMXW3xKPr0bFiuPHC4O9G+Eu8j/EUzNXoGpvesfJ1Ozo+X
jdBYgHy2l/LwtQ5faBLGYQ7lE10k2dCGYiNdk6y7Hu0l2/XUiNpkWuY/vNhM
hSyycHa/wQOL1Gw4hek51IEKiFTz+uvUNr/EkDUt8nb8AAkrSxNXh1tEAiac
9Nw9FuSyYL9VoGXfY397DssjrcUODKEqxccfFoYFXjvi06nnNT2ePWQYHuxc
vg66w8QuuciBvn6jUK1GbGWwu0GNahqVXJZtmVRlwqDL2gP8ICNdoUHbaMCC
4CtGRn3XG1lmQT10rvQurgoSNlrI3g8vMEMZj7LYAcyVlHmY0Khoo8aJYY/D
RPLy2yhI6ydbpNKH1n0xO8q1Tl1gAxD5CpPqtf0rw3r0ou4mgvFFIXdrnviS
7kFgWvSdkOuYfPYuQCBsVfJM1QT6n4HsVaUuX3Z7KjZ21iAahgFXHI4aDKwh
AaG2/54DGFhgJfydkP9wa2gylkbIatGuNi5E1xLlcOBx2c82V+6lJtVxjAYP
rm0bAbqHYrTy7anj8EUn2eLTHmllFKfhI0WCa1zBuQ0edIRogoClTXDSfvH7
aBMw9s5q9gjcCwicO8SfguT6swLzWMyRVmt+WEb32HXU/CRB5+tdi3fzYpaY
bFxkjZto/joOgHo4g8oQUbpYq0ho3rfuPVMwYAyAULnzKFeqRoIQaLtVJCYV
d1SPLCXkb6ouOk2/jkGlQ+lNYqivMsDZjwwwyk+edGfvMr64wFXNlOw51iTw
/nEDNd9bWfsWzmVXqxrob79qRge7UBFRF4gTv8cd6nFz6pdn213SlGKrHTlU
MLhVaEYOGJ515LV7AqyRJm7P1FerFgfwFI/fYQU1OnhHWhTUDFG3BBenmDfk
9dcOkC+5tnrYnpLqJBRj59EXt+8aXtYyD9ZcZ8HuNAJlBmFy+OiFN4C2fCJy
WsCCOHsQ95baZn1t3VqTSwHh00y4yDsBE1NdCPS7KfdNv+CFwQFA//kieyik
zwPQya3v9OKm7CcKfCMsqky7kfycprJZPkbjPIxnO2cmG4qCzu9ZhSD39NQr
lMEEabCR23Kyi6sycI22DIITN2qC4fz182dxgBrfdegNcCJkwrDI7o6MSlts
2WELLjABOAwT/zgY8eZRl9dFBZv26OfnVNWVUnc3IYIY6cBnMveR1qDp7TRE
8a/t9QWefobXGxuTrYLWVgO85XDONmpzqEnA+Ar7urYJSLiiL/+h2lptTq11
7VJottVzDl60pXShjP6S5nPIwioDFIsC0pOFT9e5YXHgnPaFhEHlMMAHZpNd
Wk7voTUp5jcVdPqURinDFKV2CcC7QoUJgkPgw6VQ5A5O4aD6yE7PcNB0v0YV
5uqYYOAKkU0nuwiLeeCk4ZbYEJtAf9zOPHW3qU6N3w0NBiAtdmiCAvlNSo6A
7oiW1+4WzACTim+nnMsWGBbF2WlR0p4r6crjkx1oUMJGy5qD7vEBWKuv9Ihl
w8mEZSkEBqvfTv4LLhVlME8vjOttqAeZc4aPb4rNbAoFU+qgsc+N0J1DAPw9
WLJ49x2G8tunP5jBkkzVSjh9LbhT7/VSchRq1osRUyqY1+UZjGC/UI7MMbvr
dFIYHOt+zRfEkCUYs/J8cZhOInTwEQxneFo/qHtQ1exsGL1tiOouqGWKEunk
CCPQ+2gjGoUKM7FmWAeykw05FQumdLdLtNTB1qxLHL3gdiD4S2DqpkY5m+aA
H3vf3UQNYqVxWP4g9VGntVqNIRUOqZIng325KUxnqPKAmYeYDbbvvH3djS2Q
6S804NAmzdDhdxIXpPGbqKNxUlPDCNwFol0ZiA9XpyVWdN28IVBIt3MgGUdy
R34fRvczV6wYR5vAAIS44g+9ImtAfV7tGwwFt7Vhiqydu2Wmsl5X13n6/n8K
JtgLPsDvx0aR1CaxAZV4PBNgWNO9MoUpKzgAphOJ1N1ow7RHe54yGi7xMY+2
5VqJc0/6kJwoHaHWmrorVLfwbc1VW3joBPCXqxHsPjKTWq+aCAqVNHQqBPBP
U1T1Bd3OiQCsrhE2gtAPwDqzj1ICo8RW5FD8C65pZIeoH8BachRI/VnS8bxf
doF2YbzgTNJh3Uu5CKc16ppt/5yNLVLgmAiaYrEQzaC12vT7MYmIDQf5qiLZ
YXY6S1qgFReWXaRa/1KyR/Nx4iuVMEiEQ34g5ZD/RictbJAfe49LOm2GdYjc
1OepwmmtG25e49kFGtunifKYC+bJWIt3b1iHEYqyYVBIkWr/JC8BqTuniG72
IoiVzz0maQzx8q3DbH4FDFU6ZoOq0XhuzCEBKPkw1yIvA6bc0QFxCyicpG5F
m5LmoaAfVaETO4LGugS87Hd5tcMFhBj/DsuZIqGyh5FWz1TizALVAn4awAnS
lSVgVqW7ZHVCn5eqEtrnaDYsmYiqSVCmVrh7JzbK9AaffY8oNXqq4LmUkO1f
2WKiWuot1XIh9O+FGC2c2GxUIuSo41+b/xQzwncitYrTFlahxSHFn/vdVqC1
kAw96bAejKeL0Q6zOsgL31i10WA0iaNFtoLILLulsrmhOOLIZLJUCduhPgAF
5VeLvDA+xZZmHvwGwOy2tralD6fMuT0hPwtEoS45hMrNaouu8xOBYnpaAPtp
o/ZEV3QK9sdAvJZMFFrye23zW0e6sUym9P93m/OalFsdubBReMBxS6K35ME3
ND3u1XmyKVlW+m/Pvrbg/QUMBUFEPFHtDL6ihbz6+9TBOjzV7Ys8YdXIgoE4
PdhY0WWK1ufCL/R1VxB43m5qaPPvJjredbZgmM/OgX9pUJmSIBuu7mtUeoL3
ZWQHsZJNgcyHyY0wS03zhksHI1Y1zFPslc8Tn/apxw0b3xWm5889ihTRvgZb
WZA09uGFtWp1k1LHhW6OAIoF3/M8hnEzPYr3+VcJL/2y9MUPXxpFC07cEWR2
6SShtfqXVQ7BlPr8fsHRdBlowpKQdlr1YYkdvWElfXmEnErp8b+xoXQSYzO8
i9sA1RUfzS0YLGJBMJWh76ywvW/6Jtt5hclgKg465GqRA6I72a4Kk1lV58MV
PTtKSDXJroOv97PdkhWu5KPlMephQEsf3OEJ3X+8bgibE+63Hppit+WFDob8
U8ViOiHb+Fxh0O3Va5U74q6MtzT42m6j2wRR/Tev+hqu4erjBnjBPOzL4UPF
FlVfEuL7oE2Pmn8Tw/1oz3uM+dcklmI/kJGxFh6yaiNTpJ56hSXsPxH94jjk
zWkh/tHE0sn0BWDAqZ2UaDmaUesxO7zql5uXJ3psP5z4koMp3K6FP2xJTWaN
V9vcVAoVaas++jDvgLnkKRgE5/tC0jKxYtgVxq7yJiZNDcIqR2oQFxwp1PQY
sVV/HTR3A0j0nMe7tBJMJBGeqCyOnqhz41MkWDxwhQS5Hlwn9hLf7/8k5LkX
VUYwt5rHPgivruvPBhFe1PZ4Idqij8VU10tSH9HJ24wFqKosbMidQmJr0y4b
KPzvweYys9pUVvQg1KyHTo287MEP9k7Oz/4VLnovfgfsWnu/PkxNGJncSoEZ
l1CHrkb4+PPjmE76G/LCKOYdpTRnX5OwWodvWi6IEV/WJaS3KsNcpbmPYPBN
M845EpkRAyGDRXj20+ZLs3XxsZM4W8ZXLUwwX/sa1kR2FSrQPSUmh8Q4r+xW
0FqaMLEV+PZPovWoeuYDbRhJzyvGYN/AoCd9KDlX5SKa3E8VV+ljNZUDxIBp
UJgCTjGxQyzcTHzox7MgudPMpixPnY231qGRBGiY9qsrBjQiTOaAo5JgjJ2Q
FoLyCuwEq3zDV30S2bhi/IMT1KVj6DeOpjn3FO8b+aTFeqpftVRjFhqMUhjo
EElnt518cT8jhweakLbMH4eVu4uNVejEoCdsqT19oK/rssYDJinAlpboqAXO
BWu8EsK5QsD0Bjfy8WP+htp1COMWrq3xaPEIL91BpMP0P0vbz8UUDtk8/FKU
zP7st3gzIBG7mQVeMsir28/cC8ruLCvC0KgIcGxOUiJPfwC8aXQqs9GjLXOF
TRDnxBVGzG+KWSVRCWxd7pJjCRhDBsmMHZ/hS58i0axzJcd9t7GbMv+mNGod
F79qkqencxciQCu/YGMN9+DSeZD77J6Rhr9EWVR+xU9+P0sYjqdsmiVobvsh
jLqzc0zwkkFHSM3qjfcMS82pGpI+16Kx4IJdwzNciDuIBKGyGx8fCErkYWeC
jMycbOIi8e8znOb/EczGzqdZlK1o3VKGq0P+45bVeYYBvJ9EuTRoDCYv80eT
PhT11SBfGPL/gOiQrgdfMd8vb9Cc7KV1PJbgG7GxDgVXl/FlW+sbZPtRRRL9
d80mWjL3OKBOORL87QfkBFCbFNTw2cib7m5eTbWDjXID6v6tXGgtl6BIgKka
zRdAYhFhKiC6xyHUD1djWjs4m4srJh+yjKeneXlp+hnUI6xXQ/eLdffH6tQf
y9Ndnzk9hqfEuMRXn6e7umx/Ap4CelI1zV9EDZBsEayyP2buO2nX3QCoLUtF
esvTrSp8kG4gPekNvELYn7lxQIE8zd20MagAbRlZ1cjGAbZ6dtwpmYMPy6sf
9/DL/MxrBmefAxXRovEjMBKmQyEsAB5OA6Ak1HlThD6f6T16497EVIMYsLtN
G92+XiLluuIP0l5LE07k/7uXCAhNiutQn/708FmJx2juMtvzLDX5zmBwD9VN
Nz8OBhXvgWJyjkPdZVb3pawmiXJT+EuhLlm7N8hPCFNcN3pRl1Eya0m9+N5G
EHfi26hpLDZqA5FWKed/A0IO2No30m0fNMg8OJqeJhAzGkdVEze/bSx+YeI+
hZsLq1sn8wwh5TM7c4vYyYAkCpn4HTyT3+QmzVrhHiCu7YR34ekxsf9Vv31l
/AWGneDZprSDYvcnfmbMHZVTxOCTwfQ3HkSy4kidaVNY0ann/OrcBjK1JKxK
Ly89uM6wrccAff5qXDMbVHsXxcGze9jQmNlcnrYTikArDlSnsnpIu/girYBT
5/+9q7tYE7d0m0Jw29732VYHo2qUYb4VD5/eHpe/cYL72yU658U7xps+AzqY
JvHjGwZ7sjBzNOQEDCldcLXTqrQfhgWGm9xQBQ0kaHMOIwH9UHX4f1n5VNAM
FcBRT/oo/N6NEUGmyeXRQpAf/xQSqdWxi/kxZwS1BdVyEvrOd/emKXzwdPaX
lqpc2O0kj1I0qjbbkMpp03e07f4sqOlibKRcL2Z2Wp+xeZm7ACq5JHqWUDRT
KajcXURtd84u2dERRD2N9R90TcEnRp9Fv6Hj0G68XOdI3dtSu0ajedVy7Lv3
YL16E7BRSPLS/IDzoMeYPcuI0VlJpxTRnJioLTnIDc14aaWROj4ejYYRsnMy
WA2wslJGD3dkOK4kXUAc/yowk8BA05gu5gUGplqvXWdDQ/Tj35L5lnlY6N6c
YLey7WBGjLaZjOIcHjH7mYJIsQ35X8PAbJTBODRwKsZ0sENaYMH1is3EufUV
4hMDR7c90RQ4dy1Rg6wUEkRrdawqcEYLTs4Fp+qcO7w4KnNLyjOkA/KF7cg1
aVHyJB7A+6+Tj3bg57ukx7fFf8JcYrbb/B+Dq+ARcOTIUh6hFRU0NklvgodO
Is7WkKZISMmKxm5GwArDgayGqobP00AnVcRpIq26JnordbwXYNqnxy4plVZw
9pMHAkblB1AKLA3SSbSLvFJQ0VulSW8kSxCLJmhvZPcbeqckQnxpeMHvToKm
1rLbP9z6qLp5gS1d68Yo//wmSsqcSZZa7EmyMT30ChHBnqP8nWetPXCCecWf
nvmQzERSNA0PLUHKqGwMrR81l3gEQN7oFez2UhMYphIC3g51qBRBt66wcgjD
yUMJ96E+i0svr1unYTX53sd0WJFne5V7KusNXlq6fAhzJbwOBBXpcV26Jy+J
wyxqWDLaMrdunM9ttX9rahOmytQMKdGrSN0q7guSrGPLtQ/IHo/jB99JZmWM
RQrtE9Ep6kyCiDsCdSWzBSer5NT+3F6/WNboIuXWtrcrHLG7zn5BvPaU7fsL
xNlbnnUSRAUqvpmES6yArss2vIWBLH5l9Gbn7ItQpc4A88xx2K28a3lV4+cO
WFQVKe4ssashIjbYDoBQA07H6XfAmcaAoQH7CLnrm9WtGxD5l85B/F1SJkxD
nMKaw/31wEIfFJdBMMcOgkG2ShAU2v0oae44OA2pXEB/hfAJ9cSQoIINl4Vi
leIBxZ7bCA+4sLe2jkz9BMxWXMWguu/UXNcSLv5n89ZwpxhRRGrySP7Fti8c
w/efb5Ao4jXFPWr7IMOGlShMiPGRVnjM0gUgLxkW5+p3zH7Vudi6ArdVtkqc
ngX2eXmV6ltJS0VRBO5CU0tLotcILjgAknYsBc0IqLsTyd06zDQVu1n9Phf+
E6vFZ2qsOc56nv0/+RN8C+QMS4eXkWLuln6/UVg/MIwE+iQrFtgN1h2WX5lI
HbBa7W0l6tdVpNunUfHLNdNqjr99/REb5R/U/ZJMFhFllwPn3yit9P8eD0DW
IiyNkLXbyYdGlgWQPYjfMRE1LuwBZnq2iXLDtruPotxTe/keiqm0Wm1+pitK
ShF65K9FpQLnQ3OBNsLbVZkUX80J89Z9sFbO/08/79RDtz0+ne4lZJKZCC51
GLJJxdaomzNIqbVqXIWjRkozvnYy2UQTXefAwD7fy7xgevtVBTtPSFysOmmN
EmVANpKDZ8GQoi1e5Y3GE02HSMAceiiyjgZo5nkiABzxipUIY8O3Sw0AeCLn
+fMIrUueEDEMrSdvJ56+DFE694VK5JktmldrVflnLd9sf0swJjUBzC3F2n6p
lw1SnOGoYfqSr53V6lh1qiYX5TvoZSu26piXQ+fKZuWru6hTWxCV/E2tndi3
M+ygXA3qxLNG9w+WnoZp9s/3rt7GkjY7bIjfCXjZ+lOA4qnQFcwHYajEpdiy
TPZBcjhTSwBmr5p4NgEUuSPKKXTQ3iy8heg68DCKK1ixaGRoNdiPrH1oRYBy
de44KVCiIyg0VwFYI5ys4RM2Nf9dlRcSW+6z5m1LCJUcOqcanrLxk4Tuxkb6
2B79cHjg/PXTPMCSBSnhgitcoDZ95y4Z0oomNZT8+7TKj0M0D8QmJDluT2R/
9A9DONQkwMyUKMWmIxuyucezYQ+CQYeQbsBqFWrZmKkrYD4NSM4YZ1NSsy0L
Izl6+MI/gttTYkYIn6UjoKY15IXnWcdsIjT58xvAloAiSCjpunJd38gvGvRa
mm3VvB+AO5m2INcZdvD+nGxIy8OPDjR9l6cmPdaduLHWgvdDIxtRNDgDDe8C
zQQ03TBkS+9CJj5NM5tS9mmqUXLoENCe9UPQ5Zda7w4zACCRDApg+QQ3eGfz
bRa2JXw7g4+GGLzFC5Ghcsd99xkk2sHNrGtDRIfQEHGdnV+N4qb3X38P04yM
jvrhHBM64liNGc33U3ZxNmfVcB9bMxhPu9QE0wGKwI07LWFYoiJWXD7dMRRw
hoY31ddFygQaw70jN/ya8EdjJ9Ny8xbcRLY9GgcrTAIn5FABm2gUA6SyAcuc
kMCxSHwQYz/6Adq/RuCylp4kpOvJ5wEZaA8hZ5x9n5Q3zvyWeQ+BDpaWALTR
Vp7QZ+G8rs4zVit8vGu0FeqspmM5Vh2cCdnjlPqJQAmH6js9od2c4sNjglWA
/S5dhcN+DPDJOi6jfa3H4dwJXBQyM15M2AaXuJJTHVpNuInEhprJuAKyfypM
8Nb+sMhIr64BIkD+J7dJWmndBUkMRV/IOHa018r7jOA2OWw4xGqg986OTxrQ
KqvLdsFgsKTZ8rrUDEbszAZAoNT+1f8aOWhsYbihYS+K3cpLA/M426v4h5JV
Oj0IUuT7uA6fnJdxLtEgQ8bDqW8/H16rCdX5BDXp0BXTIuOw14ayk7qyb3cX
spXyM33QRKTat2AYFh1k2zFeGzzKqWVryEYqU6Gaz2MTm4GKoBjw6mfanxXt
Be5L2tUc3O6/m8zTfV3eyvQ1wptgr/2hePFxNHoLHdzprZKZjEzYmGalsNpb
M4hpDFkHd4HaT+N4URWPpb09zLOe/XcE19qUTylWa+hHj/6AID9+6WNvPgJs
f+TW04tq+v2KoalDP6t1q0AgCUcXNciXzrxCK8jFwoTQv9AoAiX8XBTpgzYN
fhKB/R+AJ5CTdzjy9FXJLhjHHbVtCJFwotLkTFK8U0Fco8PLzkQu6oTW09lT
RBTUETsP5AFKOfMmA1LlKHkMaEDXwxlYqnh8PCr0+33g/IaBtcy1vmom/bSf
7/1WIoM4UAGEXIn4bNgrnvvjdBClvQkpzDHM2TaQe2tC9jynd0NfQZtbl9XY
hIkBfgSIm1yem2xgy4ck5QA7Gp/DGCHjE78gjqSgZHR2U9PAyDuskQstjRFF
QlRM/oFHwDSmohT+ErV7fGFlKTkMl3W5o3gzKM7GgapaON40RDE4HwW8hNfL
WbX7x9/a6NYyrot6NLWXWyTNiuHbjMsQEv6oS2Ml8gMWHLwhezOIh8FTrrax
iNdZROpuAervzzKFkgZ1bmaSANdL3xdlyfL6LBFzYWuMUPCeUVjjeyGWleg4
eDNaEAvajXQRqMiXP2bBGo4XNBy61AqJcPIsEd9HsV0Z+WFScv9TS8cftteC
dE27Zr5mVKV9+R+kdLA1JnJa2OIQwF0bv24Qho7VYPJp12xT6alPELZ/jHcf
g8AYDROPy3qBQqOKq9IONH1ZKhqL3tZjnLcHES5CCwdkO/BDijxVKaJ421C8
o8xXfPJBWCERBJFzh7R4WkIvxw/EJ2nJETuVMxxZA5R4hM6T9ar0PoPvGmy5
0h2+Nz1Kgt8BtvsP3rnfqgGo15MSK6uHQ5kRFcIENPA/YJDOS1vk2XVXVJn/
NTRMeqfPooUT0FmjW+/xpJbJIZ8l9wMn/rFCcQKaIo2ojqtRwJbBVVdS9H2l
d73WiuvClvR4FY6g3RvvibJiMTYrkkcTO5kQW6nI+Cy7rHGoVD6homSaj+jx
T2nPGCSaXuf+fmvgsA2epsV/yDKRqGjJlOZXxO5d8jM8Mn7BaQGICSBACn6q
x32xy7xP1vbkj27UMkQZVqTU+Volb8Tjl6Td/5P4fmWn1VaDguNWxu7mtjmP
dl/dXt3JFLUJohFeON0gLeF5/49rPM28CXPwj/eybIzncwUwoVwLs4ppK5Pm
QkbTkOy+ulm6sZwOTVwjKvHyX78kw26HqIg/mxHCQj/7ifEa6z48XHeL9nsT
nqMkS2BwLhcQ6I5ZZ2cIlslBXqSaVPWSFR8VyFgDwYHR1RfmJ07idE8oq+/3
bsTVfi/fkqjhmiDYYEsY9tg5wE5CncmI8Ra3Zj1L4MxW4T4+/Px7Na1GFtom
06r7z8PMUPnh43D8YFjetKbx98TFTk+1+a+tCeP0obekkvyGK7EAhwF8ao6h
JsCoeNyn28J2JcpOSHgCrbGXDRr2B2G1ltpyL5MZaqG3PZDFmid2pwiul9jq
qTDSkwUDPttX5t3gqqT8LGh+fy55APH0zLfNvGMSjlc1MZHFvaDPmAbxYc/k
Vs2UlZShxvqJ5Qc9dmiGAu2dc3++XjZJb4bTnG2tpSlw0I4d0+VZfd7Qe+nn
G7NN16UjIkEt0Nx9XuTD3SES1ju7geQbQCWUqAui/16KlO22gIg+YKVNWjPT
hYrZJd7ftrPii50PLaJhz+RESmHC5troFHdlHfg1loyepMVqU0uE7xCsvfsl
AW6CEFlbszXtL+kQoYTM7tDbPDUBVeuDF7mHVtEX+34UqOafpJE/qODnesvR
qxUPsSDqGeQ4VFnztRw1hhQ0d74kpPWBcO+lfBTvqQCF4cWZWW02IH+VVkBQ
KBBs/8ECZPVtnYVQ1tZsByP6QDn0oZKdEJNqTTPdmXNtT9oWjgMRPCdSXn3y
BS3+2iOFSHQsTzC2a9BrggxC5X773TvSLrKzcyvguZNnm1l9rNprxbWAaAOC
nNqyQteRPoGnq2Q9QrCyh/X2tR+hgfs6DNOQ1YX7JsPuTAHF/TrQtG4ghkCE
zPaYx9VhociHV0GJHUTk+80J1xHVqP/AZ3QnKQsrmVXCo+NE5e8Xx5zm3aSG
WQX7Uc1hGXJ2NmiZQ+XXBtkyDu1ExkdPbh+yypLAXUPIbYq1/4YPe9e3FgcX
RcgXi6BcTRwCJTRnsG2rCUclBw8L81WhzNryo1YlZ9qyFyKZb7Uy2N6+QNOq
9zdRNw/h7oYZGCLKVG9GcvR0mb7iqM+WQ1Sc8LKxHltwMIfs1uQkMl74rVAX
te2aDJL5I1QeNBCHfTHSvUIMdM/HoLTDvlWMGpS51mPVXKLOraT1J0Mm1Rxq
3fMgQfR6ac1JQPKuGSLRZgwUVnMrrP/DWXls68YqlaP2mhHaqKLKF0IEu362
tj/IlZpEik6iluOv/633yFrThlR3v8yYVWckLTFkMW1sfiEdKqu2M7zKXx9T
MeNfAy13qbliVKwHMHWYIl6umyhaSkVDXHLznOOgEXbdk10rKTv2jSP8i9j6
DF1tacbH9nB9OiGnlH5ZnzTdz6g7zg1+e6DiZ+QyMdkFVqq+qvL5w6Lv0Vef
QW9G0C9neGxtmGNVhdGXWXm0lohNb8TQFC2rHZJnOArgDgLEjPZLmFbp+Tm4
wPaAfUTQyGY4f795lMi7VGDrmriV8yDzLSXrwBUw8jvk3hzh+aMr2hPQ1r/Z
+PDWwNafQTxNYAxtakhJmq8Dix7yP0xVVMg6gnYCitTwYNKEnWFfvTXSW/AL
uj5ZbJV/+HkjdAqxrN0Iewp1+zilriGrDjnaPmZNvIFrSCuozcLQlt7CEFqr
LrkR6tBCXTzFgtp4s21+XTgoe7h9nUfRGaCtJMTPqkrxsSTNFr7n5JtcOSyy
lj8IAsJ9ergM2phNMRkZUJUBHrDHljwo5OfV3OdzX0Gj0AHkRBATgBjBGgrG
fAua15BsMyYA+oQevKkSz97Enzer6C0AqbVCKH5sdglBjA0/iDmTmWMtfnK3
eHc5BMVYxPRr25LegZKOnZF/+7M/n0fmZ0NafW+1lcIaH3+lTdw+qe5bhR/g
/vUNnhlp2LeHLt1ta0G1QFbKOteH82s6nOu9Bw9DOKAqtAT40whoYq7YnJd/
9XjiJY9uoH4GffUdQDRkEZecHx045UEq5vRjRqwSKcysfOFYEwMXR1gwpDFL
SCXZWKfEkFvrtCpZ0/XQWU+v1Z/AB3+kUW0bXlcOoF/P2ckL2/PhxL7OgmEh
MWxm/mSFeU06iIA1qvkRDdRcSOXUafEltrbUKMN9qrGKW1gkTl6zSisRkeeC
sI3PnMyrYmUd0Xd8P28NBItmDrWnYd69RkIDmZM/i73xRiQXXpNFXWClfw5d
0gxbfwaivOXcKpot/eJbjErIQ0HYWyS+Qoor0tlVpbQA6ComCmcsSVhHTb9P
nr15tv64cgpVLIksZbl8jkB6j+k+4VTKhCkYgRywHqka/8Aj5MDlJecBu2zK
XIa98IEwJc3b8diha4+RuhgxAQrboP3qp4eQ+MJkJOEnHs+8XmNQK41EiLWz
DozoJTjyzyCSqMG3koS0wbD7MtLXu0OopDxDKYtw7Ki7Hexhq6UpHqm30Tm3
ETCYpHcegiFx+A3gc9XKNzO9x/CSRSTtl/DfUboAAvkqWZ1fVeOLQ4SKhMMz
YEas0CeHOJlfI0SLdlJCln9kdz66uNsCI/kU995fa4oqy4bvmiqb8m2GGZ92
oPpE3XWc1oNGDPxPfZb7jwH7n7VNiDYUNJ6uNU61tBOBwU9wvF1SjNhOIwU0
RS0DKRR1Av3vpDXfaEHPIf/l+nRcdrbehuXBSN/x6/nTysxrPF4JaiDfonPC
yIG712qBp0u6QuhlbUcuYGO1w2N/MtW7qKdzK68npYNpzXzif6DcWKux5VR4
CIP2+DhtyJLmJmvql/ujzQW3FudduCcb64J8U1LNwIlPOGOhtx7QwSWfVl3T
cQk2yDDlPo9PAbEQ2rQ6KNL+W4wIsiRXBsbOMfZubgoN/vrBqDvpAIh0fyz2
2oXuSHJ8U2iLoJ+ey887AtYGC7ym8dktgemzrxCVLfmwoN1W8aNNoZ5dU7tO
xPh2d7PHS+fq/MnPYyRDjgUhtNS7p0DSlT9tAb6+EqHLwwPM46jXKeYasqpI
gDhyKp8msC6zs9kGFMSEYdGccf0yzADsMiTOlKwRvw/9nc+W3bljv1TfC51z
y5F5oQ11cXr65GUyPksAxAu/1SrhVC44CUs3FNNFHsnv7mdlnncBKG7HJmJB
53mDEnxXlgxgVW+XywdbeD6Om8FWPE2SbDXulg0xP53tBWaWWmyw9F3Ce/vV
eaPn7cYf9YBaz4cXjDTHuU7NZTfN5KB4susXuiw+CgikKKvG2sgyQwuiTlUr
f5Y7FVkJwfn5cV3hHO+tqA3j1IIwQrIraI+8CdFdc39dN8BcRTTUa3Pyxb2C
e5BDnAuHblSXzyXtAkYLgoehIZIPny0zmBMHw3r1lu0V81xBzuXrIObvS4/L
Lg6ECpAZ1AG8DiGOXMKRZKBbnj2ZmkdYMGbVGjmaBGGvw+S/yGhdRYaurFAE
qfvMzrDhpYyo2IQyWLObgqqkgcoY07P6EeG6Zerh12Gn9td+a6LY5ErZvUXq
Yf5DvuGiVXyqIXsiy5OkZAtr0RQz3mvH77OzF2Q22bHX3ECjqQm8bWvhAMfy
tKqoHNMCY4DxSswJRppSVwT8kd+7IJtKh+PGhdnfMoeOxhPXwD6PaDQGfEa3
8Ya8hh09d/WIhD3TMi7os+ip8yVg0sMcJtNY/pruJTUPnHJUqXIToXWOtW8Z
R1elO4gXUs4gDSWWt4tBpRmHW25xUjP4J1efOpG/LwKrHQRnG3TEPuOZatXf
6wuWX1xwD6VLfuJqPmL52Vpid1qBtWe/kHhFRrLCoXgxokFwvCjNYl6TttCQ
3m1pbamipdyYSx9LaTsx5NFYvYCoqqhNUAzW5fswYO3kXkv866N5736lIKg3
KvODmT9veL+ImplWas2Y43tK5PCnPSwHwDBV9qSxChrf8J+mppWZ/Bq/Bd4e
pUMNLQb5nD/cpylNW2cGgAVBa4iK3KuU+jP2KmJes1BmxiYrmVqNMKj8jsQM
rFczY4g8BJukSfd1tyjAT7JK8Pe04AzrCfGDSjjN/d7gSgstAAW+JcatWbQM
lJz6ckdw9jPsZsQgqUrxSZbCH7rQ9FtYDFDHBrblIp7jokgn/Oiz/d9k2DiZ
DxI6G1QVTt4BlS+eYq2UaKJ9CuB76+tWzimcXG9G1C5ru/08nTMHk2462S0R
QrwuO9ocJJHoYD8IWvMyO4jbxVcEP9sTpEKtA+LWTYuBGujhgem7r9i6n0J6
csQI60QkfBl/8D2Q4A99MRH4Uxgih9RZPjRy15/W71xTChjTJx++kP0wZ9os
P7At2XQliUU+mOQm5yF5TDbOf2q6GqQBc411qBFd2O+4FRPA5ZPiRc4JC+n7
5qVmI0tndRYA416QPTaoJ72P+KRP8GPJfQJqIMniPW/Z6S5GpqpfKRui90Vd
5oT/Z5WkcuB833ufJ+33+ZBfnn/xFXPxdopSKcdpyUmEYgDmFPwCkEPz8V5E
C4+0ZBiuwy7/wa+ePDUYQZXIutqK02u8hWq1BEk+bTbOxmSWEEpw5KuYgsoN
qTRLVvh4g55frzAM7GW5V+2jhgh87Yft+96U2Ped3XSQnXk34SchG/BJLJKV
hWsfak4Snggyu6WQZZGB7B/X/85/jMkMn+iJ6TsTmfUtmFd8rKLtGKqL2Bgv
Nm91MT9JDhHoThdHw/AHKwO9uPDuTUOaflSmpY38p+gyVpDSR+JNotYrBJrx
sNpmirG2qmoYLa7tLGbCt2p+EkV/IxW+S9IT9rDSHIVIDJBV6g1ZBOj+wJwd
Q0d5ai4NJ+dw9lT64CQTF5pBlZ9oDxXs3z1NMPZ2VcO8svSy7ob2QvwrGu3g
JUT9dCGGzbH9kjAUX/g+w37kDrct6AmFwGYCWOnpXtm2myZ701l5OnVWLVhJ
NJpHOXxncxTw3t4UTbYDMJ8dAqSE0h6VCh400Ddb3QWjsVCLaiN47M77oUes
jCdwCPT1Y8VceGtLziAFFLTcLgkN4g0bh06wHk3o7Wpqb1lim2VzHJN6T5Oy
V6j1YOfVK2LSCxja3BkXrPVY6x2u5esGE3m2kJLV3MPNPLcNqWPr7KiXs/pM
RmP0DS2/RUTr7uCxrUHjIlwVu3V+bxwvxWdGRZtr8fYCR/yDU2hQ42YFgXnm
n4vMrLHpH4wbPlUQC32jOkpxhv6Q4H/7pZWAYqAkvQrP36fngxtLQjpufNcd
aJq94k4ocaWD1Gyx3P5tOFZ841wdi2kgMQFgQoCgpEIuhkdKOSrDsCOGrOJg
Q/05Mnl9jOS6arN9j38P1lHQ+KlYGDfb/cVPAlVknDAvsIafulDySkSXgd1G
DgwE1FbqtO7OAs2yGhl+0/SsNRzWVUqQKy134FAmrqgWFz+zHSV9qITSVtT4
T1Fen8T5ctoNkNosxkw681bEQMG/VozD1/bamKqtH8O5H738v8/mAISJx0jf
BOihpmsdbw85Ys+yl44jd2htETRxQRjqmPX3fw0Cb2A5Uw8s3FT3+vblo2kj
qheXz/C/rsSQ9ntUTmGNubv8n0rD+LcPZ0ChEviaMYueBL/YPFMCkGYHjDhM
gEp1s1LjgdwqWMJXRMlp7iB+HPdbfrQdsJlpYY4n8D+l6Z/PrXEZtcrh8QlZ
/JXOR7ADEJHta0UWYJ3zyV914uEdSNPji+IGniF1KtbEjxs70Flb8w+s/v0l
U1UZhvzQNahu3ykKr0lQwZTaE/ovjsv81vVInM2pSgkOXuTPd9yLmOyYH52m
LESV/aIpQSVtZPbB4iWGD2ut3Hzkd5BDHoqFK5g3LF65FLy0EXrSMw0J9Bqt
3jPs7PkfGbQgw2zmaEcIOzsS0ZsjlSOjK3e1pRvSQsnNP0VA3QWMlZ63IET4
SP0MfauuBI7IjGJWM7DYsFBhONkHMB/3NRTYHIWz22oRGtDUuXqXzp/1QwPD
6C03p+BobXsVVSP5cFpRV14haBTkkuyiyI1+rPFWakH17XeZY/56Q8BJgkOD
l9wakiKNEMIIn59haPxHtEzEJC37Fvz2ZrZHBBSG4nNKi6aUrYH2kayxtx8W
wsezJ7EhQiqL5ZkShDZIZeM+2amVlZUfIyvoOnsWZqVJ+Jo6fBNOyV172vl2
JhXHPdItSmOXwH0X9HlOyEbAitgDPb+YcAFC3bnF2wZup+EN8FeUAp+36gDZ
heb4Hknj+APQlNtePm8d4Rf0A/UnKlKOJUjJ6tUOUFjQ5H4ejLiScxLwHDuV
oUIKARaEoW9fdmFHVxNIOYPfo3XE55g2Fups//6bCI8mgu5zjABNssZBx69N
DvsGPI7CrJWjFlSYkLQcGFFJBuSTZZd8NtToKw9U6Pl9bmDltoIUU4x663Xw
Gm86knePtu6xQ5GvD9AujBkIlTdym5c7q0QUHJrR9NRZeP/a6WX4MAwCtmNH
4NJn9IR6KBVp4JS+LJmW01ysRN9u5KYhpSN23Ks/15ywKJGTZerazJFL+LVA
RMJY7ooF/rMdY1ZwQyuq3BNDE3FtmBJWi5r1+3b8pVn00jmNRQg83xbo47Cu
1CSWb0GmXS2ayXmTdmJWQ9Qun5GhArizqz6xdTPTuSe8iF6OKuoEiL/dDfkv
5hjrhXASFbnNeWsrrRXQ+qyZsp2+nsa8rTgGWgDNlyeNeyL26ivA9bYI8ioB
viF1Bm5/TZ6igHRhheReo4AJruPyGcHIIDPQOsM3GKkxjYeNgG55uvLwyABA
8kGM7LhkNioXEG37v1h/zjbypE3qYCGjSKirxDQZlnGxJx6KugCzCYMU3mWv
CSrUm396J67HNXRM/9NS4l700BJGvGVNyx+R4cbNnp/ssM08G4tflPCjUtcU
k9c5ds7vl23Q3SmwauK+c2jJrSAG/z302gAuR7aSuSIgnIBgPpALf6bfmdJP
fm4gpbbrgUYWpNbsIw5AMI0+N1VW9LQqKnKTauNsM51SL8WoYvn53J7Rhd5Y
RKwi+IMG+BJoNZdiNx01f2zzXGKp/SV2XzjitxWVVp0VR6tOWsS2o9N0iT8w
GElUKqjL/5VzcJPnZzxh7KDPOvkdN2I5HDqvY+P+BvRUGypUv6SUH5xm32t0
iJTJ1nN7fCFkDxQ4XUVY+dYHDjAovKUGHDtJsVyZYmy6cv3kwx1fA5wXd8NB
2dXRzB93LeuA40YFVtC29YwrgWyY4NV6+GoCuZ5svsC6IddcqYFQCKvqlDWN
Bk7skbTHbfmQ5KuxOOQdVl7Ha8x+Pcizvr0UydEB+GFW3rT11/sCTLpyvvXw
N0ccd66eCtUQfeaBqixsxcXLszO/ScfS1ySKjcVRd1a2YTTA2UH8Dq5sS9Zd
T0sqiQ1E+I0eQFLymqT1t1gKFnaQ5s4fxqVsSoO6gjFUsHaorqVfVMpm54JA
4w+tb2TbcYx0tmxFLLuk65pOQE2Le9ryg66nOtnppoWjHAmOsz4PXTHJ/kb8
y7t96Ln7SD/hOKcWglGtNQb0TR43KpqGyKTIIrV2jWAWD+znWVovn6+2HBKN
QDwWHgeIqboFTNHkwwHzrIH4KIiX66jOJUUZ4j/vxokwhpZhdk4z2NYzpvp8
1i0+VY33wp415+9cA917EkNnvFCL7iXrI3dm6TEU3h8Fgc14SVRmRax5yZuf
4fiOoXJxXaMoTCrXagPxI4jAVWkdzYmYameXeTXAjhCnqp0/41Y7e7nC3Sfr
8NajTuxHEl0Fsvm/0u5e/F4dPHa9ybp8Dl3ZuVKEGjC94VsBV/wpDO7P8/5z
65dv1gzaZdPqxaQUScyxv4oop7wCe/rSjcEFRWz87RDw5t1t1WRwQB2hpbt5
SF76iOTjkm18TS66p1rACmklRoVszgJgO0jeCYJAVtGjp/jIjxRonlzmwccR
J8Ajwos9ByaxrhFfUzESVZnUYz3ht93zCF8C2aEQwHqK1ZJgmmkvarXihXki
7AxisabTTbQOECnccw8OZ1bFoxkLE1WpR/DpaRJ7ImYYEN5oUCg//uq1mHS3
jz6rxD/aQdPl47WcXnPvX4XhR7bAiNj5oQ6MI2fkAiY2HwHKB2IayrWjh7So
itCJcIg5mvvfYcSudreadeQ7MGJhwxLHKqTlu2r1nTO+nnGq+hHKEAlG9bAw
ZNptTGS15ALStmfsQimBAvwmhabJVVoicPoPzOZQ6puObYf5wa2Rrh1WM3Oq
GKY03d0qHjCVBldrM1Yq2T96Im6BfufMkEiIZvBMxbq8RL/ze5z9zM4j5Enk
IOQAmavfK90RLy/vRAxqS1r/SDMGw0QvhIYJzD/NxFFrXxfPEkOHAMp9tZ8w
loIH7aHzuxrYuBR8uuCv6fPm1jEtOHvsUbz6mxKxF4Oylnk0sp2jVP7Bgge5
93tsiPtcaQy0ezcEkbTY457FEd5yPLnCSJEPqHkv0q2Aa4pN6bYSl0eCf6P/
iuaa9wvu9KDHJl8GjUPEDjisnJz+gOlWC1U/wfWtlSutK1IX/11zrvP6PJXS
zLONeaD3qx7KYDyC4vIoAZIuz6woE9ywd4rrh6QVkEQY3uVO/742epGrNSaA
9be8sIyQ7ObP+wzZDq9T4neDRSsD+rJ8PpF6MAn/FeBonaXL3lpB/U4dN4Zw
I+fqusqR0IeEds6fPLuPMqOz5jHA7/ABVXFgzkhkQPee//gY7R+e4yAAJB2u
ZqvCdFvMDYoJEcPxS6P4oHJcxdRd4SZd4DR7YR1UqIPtJbkyfEj1/awC4yZG
DFb1X/x901xIXJsrDJenoFBUWO38wOdohdgEO98I+b0/gY5BHPaK4Z2WXUyW
E738untq8cvKVtiJwBx6UJESPZvpkzzXWip3TCgOdQEdXhzgkEDRek3D8lJU
oBh0hFGhk/3t/MHOknDtluLKn20g80+jrR8Ph+ji0qsdDrF3Uoc/ZnjBu4Lu
zwmukHq9k2AaWX7GPBxJBjSKCkrrA9/SMC55ssqDmnDcDJgmkjJjqzI6oO8F
2j18Bgwj8ziL3s37QP0gKUKKZe2ciEFZobaySiWK6jO/9cJ43hJKzexpPtPF
75Oa/cwVIPdYdbtLT3F1MQfoaRf6sNv/Zye2x+foXcemH2k9etFVx+yhDtas
pd/gnchbixzEvsGMCDUj1o4EsXhQ7+FY8kthFGJkdk8G4qF6na0v+3lHYbZ1
JcgnLvnv5x+RfSLU5e58jw0EOfZ7eIojUmd6KyanvD9DyeYUNlCM9FWYzDpv
8qzxD63RuY7LJOSafFYnPmjGPk2UsWj9Q/0ajDpt42p/2+lBGVpxTFYi4kD8
oh6hbepTJRoKKsxe4m1RYmasw831fzG30s76+Ea6GT3CFFjn+Dc/Ngwq0GKI
UCI/e2lfeHDetWBmiiC+7+Ijt/uz5GonYfQds3B13aEC1k7WqwoOGK7MGpCo
+UYLSd7JiHDtFnMxzJXes+IOf0RBkqjVOpMXzkY+TxcIXRU45LremUaf9orn
ZmqMrGpYvGkqI5vlvgOhamZAB9xnJpHVOHtjNP/S4CeG8djYuFnhrKzWVa2G
qukGqZWmmMGDUUEa8ChLTlpKK0StSLlt9oeOitIaFOMbTR5xfJlMRyTM4dU+
r59Bw62M89URnvV7Xy3A7JAuvS/IC/+rCbO76N6c2seapI33xVzw5raz5xa4
deO65dI+FXsiaVtmkgvkaWolaxugzEJL1Qo3k3tXN8z5gT0ll+XVUM4hdmRs
P+JzxB6XUzrebCVvKosX6yUE7GsGAmBg/2z3IFnojgnl2eIIkk+gcELIeE5T
uBpO7SttaagsPwo3ehpBUPfauHkzh6qJrmQxhhgGXzr/cC7fbOAFtCzlx2ft
lfFvFYq3uldz7BBu5O1pXEUsLGgtsL1+3Yi8mK/5LxcEIk2zjMaXJGe+RLsA
sYfPnNmHlgdL9GanCimziOYzUfGBBwpU7uc+p85SyRIIj8TGW3yv5u9Snocj
tBeg1MClNDI3ijg50c316ft/1caBM4YZWwD6kRTOk/NHaHntzrc9IlL4EIwa
Tdkay9dyp5/JImNYmvJFqYr3mT9KyZUu9GyZzf/sOhKhjMXllFmcbOoXLD31
bpQij6pxKZbL3he6L1DcH7RmJo9dqDpX63BVOeHXPx12uJuTkqdALGfhCT0b
ze11habbskZ0Ds6URDndV7zKakZKltgLTQaCkAaPwwxHFi4qYwVuSSmteA4s
7dHBsqASfB24yEwriRzawtfFvpeQKMLJlqQDgArQg8yzvKxNRWgsE3D5069l
qR6VHL3aYJBlN7I3H9EPTLDBxhdnZxpEnJ4kxQvOfkEW1/1MUkkkHCqIZ/to
7k4ewfe/4JMdOZCXBOYCqEgN2DyaVYeXGjWaEloB4YSUS3GYgwxkCkLjf1Bx
hP2+z7Zg/9orvsTBemGzdK3mAaD9KV1Mg2ONVXi6NK6uRBLPTTdt2WMgebaL
rvWgnY8s/2ZHAMyrw/tvHC18YKQ8CtHUQ9a9vczdHHp4qp/kmZJ80ErksqtI
oqY3GUdF3j59Ji1QS+D6ulO74grrpN4q558D9AJMOL1AZtBdFXo3xHktvVnJ
Y7Ie+B8SwurweleMlC8AZKeDdhH6MhPPo7XD8GxSSuHC2d745Y5qeQPVBCfV
JvlGAdgT8E018Htk2gn9Sga+RrOem6PMXOmk/B5+c28opx7y8Su3zM/GOwtq
yr5B89v4DQK8U9uUXYdXRsSAiVqbNpspPSwxLuci+G3ynMJ1LkfqtHXr88i6
SlP1BZyiTo1y8r2P4Ldl6SsJJf7Zc23y9FsqL+IXoEYcl9VPam+Gmewn81sh
SvtSxMhHlu+uGxR5D4g0aEbdvILXhZ9Esb7dyiVnW/H1IXat4ZDOt5nLlvLS
PmrY60LUHE3BiVdBneBdA8VXlnQytxwoqb8OUaxO9uXY5bVN8JfmKxBxdOi9
EwaLGXIHMIiOqizm+0cqRIDZRe09gARIP3cIF7NLyeOap18ThRDjbsjkdqW+
AKi4BLDg3YCgP78J8CZLQYjrnzjRxs4I9OQqCNDMKdeNNzJQa26p37heQ+V/
2HMWB0ppLG7Q6M4t3Z4RsDq8H6wGz5NfyDQq7xj5dw0lcmhIKGlbofkmtoOJ
K0wHrGNbqV5d80ipP6Y8BY/Je3cCSAC74D9t2I+swVdnoMHGr/93qHihdTj7
TdtvNqoJqPRmTRY+uyPapjdxm8dScohdewHyg9lYEYv3YMuCEyzh+LWbnQS+
PAQv7q7Qiqp+3L8/APOHSQhaZTODyRXUZ2sHj6XGXRxysSdnRHtyasPJFXIj
LLRBQk51gzBmbn3QmuBwtixI58U5pi7kOPANmF4bBob/IUF9NdtAEnMC1aYW
KKH+KlmZBJ232eZ0UgjPUOD4iac74AXK9S86mu1nIyQYbL/ZIIZ3YMTCwwUW
8RqQ1hS1cCL1qRPydMkjmHHWPfM3Qc2T7K0YL2e9f8Gcx5TAwR/K9R+EZa+s
6NRmrJkAS2xbIeFMYPzdaVX5OamgqSGQNLiCYIwAad+1ggT2EeZrWzfvPkQu
5VRNCw5WKkeLpf6IGy+Jbg5lrhd9Iq04v8nfkTzHPyzdIOfzGQ22xaIle31F
SP+fZTHXfmlUDN2s3CmaPLbSHRPRLsnKJxEgJlDOuhsJe1R15So5txtltoMg
x0SBDFj3BUR/4BIWRXmqbbFR0MnHnDYtkBY8oshUpiMXtS21J441812C0+xw
iEGEN+mZ3XGlbtES/wUjffxmqjUHTdYUzCXUuBd0K7LibfDd6uKDFTw+q4ER
UAljeyfGYLnXBRxW4HS9gDT9Kes9eINReSxORbsUDBVFlH4zXhwazfZSRTNF
GSalEKfSNstbH0HwezG0FA3KRHmBjEsO9rBcBxysX0gUz/MrjR6NUVHerP8n
AOkqe3Q/7awCq3svktaqc4gNvLZ/zVBLmaP5zx2sRnK22FJE/hcH8bO1ye8I
4Ib7IUtYzdJAHDN85aNz3BgSTXiqWsbYkhxd1KKNo2+6839EiMfeRt4wObwH
tXV5oF1VbhP1jXREXyj0/RqVQ1GIRW6RpcLEeTAceEw5Fhr55L6ldvomvL8p
Gd+HP3nDATCkh83D+QPgavw+wJ3Ro6vv56Re0x4EyroBxxvz1Z8feDTLL8ys
Rmlkd/M42WRpkwc1l+lBRMaFzEdfmPMUeyWuO7/V43Sbi6aMfVmUrG02P/oo
K+37lzUKekD2wjVTqzfjF1B94Gs4Jlh2vbxOE3bb6Kz7Z+Q/F8WeyQ3u2TPc
rexHXC6+hdO3xqiYrmJZkPpLKj4EBYw068MnBRZ48c0uXFcYc/zm1uXT1BJM
iDfpuNMapJZWCSbMjDufybM/NHvwptDL9PlV2bkS7tLBGyXTZIsm49S29DMN
jcM1/GrRwstUpVGC/ml9yRHxmOD2w8Yr75JA1cpqfZBZRqJytluKeKLPrLWV
5gXpJpnr0Z0D9z5i0hBYW49xkGYkxyFQKjBl0p9tZNLdSQQBr1Q772EWznXB
1u9pyBGlOft2hT9Uujr1tzokRTn/DeM75EZ7TqtRdve6gxUBxjUJYKsagRoz
rUTtM/n1ygM+BlqB6UaUgIDF6aSMC7CxszWAMMSsCRKuEqEwu/C5c46ni5wk
fftktDlyKO3Md7Qk5rv4OGK0N4UH8phiELsQRzX3UUxQmFdGox+TKR6o1k5V
sLdLvJPfE11kD4HCqigd8iWfoQv+mQU8OHZ2Up1R5ULgSB+j24PNMccQ2qlJ
eTqcwuX7zLEz2DI2M106Gi9vx5IcbRAedTehJ7+xuP6ctV9gaWXENU4csL/t
BHzef65YVapYgSEzfyb4EM4u/zApmWtx9NrQlgpFseo0ohlEYd+FsLczSFAx
jpzR5yhHn8YufHZRXVkoYl/dIjb2PzRRPePUgI+Rldc/zYyOEEY6CA7TUQfG
XXiOTR+zL++aG5vFUsZ0ldmYs9PysM3NFL9y1fFYyuxgFMbH2bElFL9RHYtN
2DMsQ7+6L/siZSnYMo3RA7wZx2MgIKMwUfgSmwsnz89tuoOFud0Yi03Jx5cE
0pfkxYrCAh2zU8yp8YqUBPQ5JHZGYTNyLXX2tFxVmJVqcOIsS+tYV9GxVvHq
pLz2KQSfDsu90f7+eYg7pE33XaKyk4gktUH49/cWqBYi/2qYmt4hXgFAtNgb
CVTA0oLDuKwnE4RUtTSsgDDCz38I0oD3n1WhDr1fqvPBfUrErIVl1zdMfhtQ
F9LgDDyiKh9PLFacRSFqlEXAY8+QC0NCjHHSIr8sLbFq5Kn/OYLt7HwaEjju
gAjrQ7YNBvFbF3rutbwviWDRvfjvNvmu70WsR4Ok1HbS9QbCBbQMus05pqGX
XwjcVnATqA5cGX1Fk7axhluiZVukB0MsIS4P3kbQoYRBLEpLb/1FpdOxRutJ
fI/Ey0VPGBI9AmNqLn/uFWXeS/lXFbrHucFur3FZS/vqADNgmwl1FZkWEfQ1
KeweySVuRzQ+o6uBBZqm6T4ERZEuqAR0r0g09WQQ4XfBfS/m3YVT908o72bD
qz237ibbCUOFZVMG5qDWZNnwPTFzjM4ukHSrFaf36zAvsLIZOPocj/FJKJa5
2tNjqCet2sRtbl5AoRYnamy+Z0jDpCtstyOk2NlWsDa7wHahVLBPKgcT2h53
XpRphIqTy6o3fRM4zJVyv7/YyZBpj+9Hk3G/PlpR8m5lGt0kvXglISMX09HH
2s7Aax7wT3sbxUfgBuXBmMLQpV/tUAQL2KeAuGIEfZiCIUEu3LQNDhQGQuUi
x87snpByhK/WRVrpJjZtRTwURhuWL4ruGaQfzOTMvtVcwu1372bL/QZ2UkKJ
RKrbZAaftBx63V6ZdqPnmwoj18satjn8ysyUGTgwgzupw0Npk6bFsIO/cwrR
N7jmY5/ATTcvmR48aTXxArduTqvSO8vXB7yxah8pVuCrpj5iC3K6FD+Qdt9J
YGm9E9LGTy9K2SoEYw/01LlZItula1oGy/W+yp/z+FBygVcHFyj2+eKjRAhv
KYHEwbKAQiGoqAn4SMhem3TRagnurL7Y4VIKFsQPom/CWjSNMMPLpZ87jHDh
Bpr98vh0piCPNxm1poWpDFvztK1mLMQIQJDsDcuhzgjacn95bh9SDThv4X3Y
l8WEELDHdlEw0xrv5DFiutT1u+jfztFJ3PO2edSXOBcRQTCpnvBaLI6T8J0A
tkNEmfnL1oIcf9N8b5SlCt08yR3gUCnb/otzEyoTcP6uaPLeVbFE6Y1wt2SQ
R3+D9196tdOL9cQWEUkyeo9fqV7B9oFg8kq2So8NTJQyeK+NUXjc3O/SvSEX
R4j+F3gMy/vRNtUTVQrGaQQOIqLws5PYs66TSWU+bcYk0Je2E/7jd9s4dk9M
v4Hmf9Pdnm+VUn+jYems4g7iAlellkDgUE7WMIzwfUBQhjx186Q4FNKhZHVE
aSdykpKFo8u0uGsjzktksSLvKNFq2uwLqCbbtxGij6nLwk04+qaFnp0OPSRq
FVwu3bbbaOehIYCjbv3egF8RU9Do7NtM72RqlyuAYmw5cmeU4lKBl7RjxP1s
/P7P6N+FjoBhGd7A/w8Bu/7EQFbWPvTcYW5eofOG+R6uFvBL/oqEAzG4kgTR
8EYGnZ1XeNf38Pidrf3fMHECU3meYjyKL2/wkY0i1HrTGcXrdB7acAXadwnd
Sp1WyLkeXQW+Jf6+3Sa81DmYj6JPoV0Q6LORb1rcwucqWTX2fcD4kBJoVLlP
udwyxvYT8+BP8lK5U005J5OTcaa7X4vcUMJJCiJ0e9OkOhU8h8qxWmQVdgaT
7Pg7kmdpxyPUEgIG/ydwDEAmY0fW1RMWMLul8ADUn7n7AAR0EOI9RH2K1nsw
FCgq8p4BTSJvO7JRtgEci0Qs0NlWyuzfamIIMqQhhdpkfhKMD/mgriKbL5wy
d5i2pANEdrP7tlhFblfrc+G7koSVcfl6+gDRh5vPZQKG8wKk8lBTtvPUDgJC
yk1UBBei6A46sf+xPuwxhjcQ1B9qUyQpACaNw581wLbHUi92shvpbNX39/+k
6dzgopVt+ggRBhTojwLaVTzL/YbqXsltL9crPY847bZl5x1PBKHAQ0gbYqyw
b1IZ5KxetQzDkuHaTCmQaeyq2yTFWOtAkKT4m9mSjoLRnbw1YXb1UQmeVDs+
U0zDzwCFhYVIX2Jr1JLDubkwejSJgnpxrgzupK1VeXI2wS0eFR5EDZ1s3UAt
CK3g1ocgyg1f7aN9ttniVJGeDYeP+FKmWdR7yWpQm5JlFtrsaXi+nrIM3c3G
OHbABSTcF0dXCFKAKlaBXglA8R4RY0JZHeTnOJ8x+nUcgam15BcGCAH3aFjt
Xaw58vbap68qg8RXz2CNne49A43NxM+c5k/hayYq5pVaQ3dEzcDjjRjUbe7Z
1clfmv9nA4yV4/AsSelDzS4gUEGlDdIysD9FbeuJb3Zq+2Ra+64V/YGXFl+x
wmp0WVZa4bf19qPAlQZyTlkvWqg2MKUSqxwIA7cSKa88zU6RFpFFTNxkSHAW
v5qsyVW+p5c+W9OeR+L4Or2rGSW9O4TTNsxB2myH5DDnDV8nKHPXO/jtzIeJ
SoW68mQBBAdt3s6NkpgA0+cd4x6OV0jJJrkKJ08b/slF+xzeoMNMBUrFEU5S
kftdD7bl4hJ8X/WQ8dGwLJtfQNtFyJzX4OimnDe8Aei8dvQCtIzaLncXlFsO
R8gtpP/Jvq+HrN7cVHnMiM2cVZ3wYgpMkLIjsu/lVkLhuxaE1A1odbDcfww1
jYIDfKSzLLMBn0dfCGWFSs+xmetu3oKsLxFg5HKxQQzNW8C0cCnYoJobAPgK
PPNWNfKNOQJuj0UiaEyCgLUnLf3prYCQ3xCyjMLDg54lugHVttvBMB/tCg0G
EtMwVW+Yb+dZ8dZPezCdVrhOPqOV8TArNEfB70rQJPg+sTfllXPqMoBxnkn2
2PmC8gnD2BUaqKGay31x8ElLGNJ5QBFUxThiicdJ7uaWPBJ7ZC+v31VzkLvT
9qmx6X4rG2He0n+aEQyPP1c8ejalnIPgHPYLWZvvXzwwld3spbFNHzGY7Gz2
SkHfaJP5+ZmVqMUGr9qkfeFEC2fCNdViSTo7z5XwxtogjHRbtRe86wVO1gQd
kyChSp1hlUatbo8+X9GPVX2HdN6NcfyPtlfqIq1Jfg9IqGjf8iTASw8VsJdx
jwexu7sTqzszvL6yn9iYNBkIrCrlYNHuiypI6/74t3cEFfTivOoEoMI3J0+j
VfwK64HWSgWoQbd3SLKqHOfwA0djrxZHZDQPWK3BN7r4p8g2/1xa+bxEdrhr
Jdas6vFMpW6o4I/xsKgXTb9XH83ihmtHEOGIbdeHq1zWdK4RvuNrJarBihmi
R3vPuQIoLBoFNgP3k6pKXPm7r7VNV+oAwmy4DfHwr0gP6YGN+yKrBfptsXzV
+/QFrluw2JHCxK6n2Y+H2fiJiRQPNszBQPaQLZaJ2PTr7+jxEqUBa2iAjvZQ
xjq+8mF0R4XPgqb0t2YYXdCG9iVOjndTBEgVlUtY4rwXLs4ikQMPY6fMrhYL
lSM2nrDikq4mrWwJcDSbqVspnTJU4htkZBSXDhUDVZjyYSOO47LJJyZF6szh
dvQSg14VEBuAjULGoQP7Pl7Dxnih5vrnxLYNmbo8GN/1C9hRHwlV2Zcy6szL
1LgSBa/FDyscou+L2BE/noMwKacWZaX+4mg4TxQerG0QHGU7IaJKOSJshzBe
+3KrSfebi8Vr2oK5hIOhKBK2iXVZePAk8kj7uEHbOrWRNfclpXkLrmXs0mSd
gLA0slXzogTQ9zfUF6PdVOzQsiR92PS6Ui36rmBpzTaWMkSli+qTT8ji+IkK
u4LcOlYp6wXt5ZyUBKHxJ1xviz2IfSHQHKbwB8fm1VxKzxJg8jW8o0v/7nvk
Wfu6d6KtmRyGngCV5mxveKeukPv0aiZgAa/VC+CvJsdfueWkFfdAnZ+sf6W9
YzoqGLPU5hrEbvIC8E9hvtLF7hL93bogTREy2eAzV8cje84Ow1yf40nNenQR
XROxQoKPYnR25rzhJXTTcISGswStUNPFPGQds0ArnlnV4eKGaxyDsDrh2EY+
OyFTzqBmIbnNJBBMZQMqDii0LnQl9+W4FfcWgExsHgwI2Ee/DZhf9MCnzd0p
2xgY+USiXBfQAikXswVmyM5+DZcy0RlvDhPHxtwj2QxVNJXDAZySi9ENOWd/
b7a6cbmNl8+Mb7negzEMnaUF4y8y2ZnW3DnYhQcCmON7XvAHeecoXA4fHytn
NdTcECnnUCTqLcmHGeJ3XkuY/wGQFsOj3coAU56Um/YHw6Eei7FOXUiBv9Lt
Z47cyC3PqcO931HlA5f5n/aUW6wqfnqAQ1thcYWLJL7qC1GXZ3yaXUS4DVIm
AZx/Rr3qOyJQdiA0pHMxMKTCQ6ePG9/qmccNNz6J/j+NdEMKJ2ruFZ1/Ktom
dCrX8c640DIclUzHfpf8ooYZbXY9UxvxoTiZCoepj3rmHs0S/hd1SZJtfelg
GEGeVu4nP5/6lglfvMIPJpmvcE6j75JJqGV6Pm+2NWa8ZeOjuekcx/JIkXFQ
cPwastS4pPFgU7JFwL5T5B85+2lMbJL616bcIc0YSScyzLEiFUTyj2JmIEjE
leZ7NOWS4QqGvO4XPxxKU+UuJoeg3WHo3D4FxXuKAk37pdWzQccJh0AwoM8k
07JM0ZpcbAAqnsZ+/e9zpMdsTj2TyBdoqnsUhXC4CBP0YBI8yJETD7t485P4
hJH6c78JqyzULaLO28syd8bFWTPB1BrMLepDRv6GdeUF9RmRq8rjsVkFLmwE
Zqea2yZIqWB5S2m6D8p6nn2oKIKmPoCfRTWkAkNCQTosC6xvd37vcpQ02yZ+
KVQiI4ZdF/9iJWNyU+8XmPZA43FZ16rnoXsxS8fy3//CEXMeiXraTB1KEcto
Yjbzsk+eZHIhvNmaPz9VwfUBE4gr2E0/c5J8SedvaZn/L0+7t3hV5SxOKmig
5cu6E/P9+kRN0CRYQA3Rllz4dJd5g17OVF+tI+tgWpr7wPgXLwzx2t8fmwIu
HPwgNeMbYXLSxyYa9R2eoLNuL+lwg+XjYgeEZ4DhfvGQLOvYV1g7efPkcbO2
+PoHDCeeavELRPaj2OLJ1SmcTCEVVCQz/Fh77dap6Q8FChYtfSEnuK2L6yzD
mJcPAYvJ/iUu9cozo2KjNXQsqUUqzW9wZCNDpkW1x5j2LXEO18bbQizslElD
JJvQLza3PHOz3nY9bkiq7izDYO6tcQ/O75Y2M8edkUPtPJDYDauCcBnmbwe9
l2/wK1vi0RqzJXhQrqFuXlQh/3oSfIgBPopPtwIcnmKwT1PBN7iYqOapBF9g
GmRnJRoWjpwf9CBZR/DjbuHyzLAJ++Zcr+gL9CX4gWdlpsve71niWO7XQWsm
tC1yNJzLa3Ui6Dx6Odkk1ST01FdJg3mYwF7ajeD3TTVyr+8JH1vbFnp1gx53
thLwEqgAUtm3gEgPWfgOYM1v8kYOSm+taw/16xg2kx3ZXQrcqFw2xUHfYT76
SR/gHNGp1KYP9JPPFYD1otPguyThWuAyZ+AulMeLoyKFKOJEMjZU7U3R3Mwm
uI8YQ3CjSrI0I/+dlMWjbw9/Pz244+fACa8DBGFeFFh/G3C/rldWN+BvZ/1v
O1aT3TshAudzn0eYLx23nnF85Ul7gCKuLsGLvaSzQWI+v+Elq+8UCeewafsO
dJ7f2lGRAcXGrc1M3jYjcsFZqOmiIZliY98QuGwtoIoeCgyg464S5r6/4c8O
dEAQW8qyVuoTrLLm5pO0dBc17fLhSl1x9OfJmpPYkQLgfj2pnZ+/M7KlSse+
ll8Ll3HO4yzwPwT63dWGvjdlKrmVqpSAsEWZ6svaY10evfeheW2Rmv5gxHej
DJ2X5Xi5ZUS57JIw/pbBnsbIdrhkaMNHVqiiPpl1mIYBKfOBjbMtzAIyNCJC
Z2mPwRHJ3aJEmN+ICvh1BKj9QXGWNlEfxQxD3DR4zaCg6R8+ZW5bZto1bif9
47mZfAoqJUYzjXbeb9mkwZMKTlBUta3pOKs75pN64Vs1fLihPTQ+8eU+tH2K
a0o7UYfygJPVBDfrCDZ8MxzSWmnegWDqvFT04v+dKga4I0RqNhe6ohhdLzDa
hXuUBYJC2AviwOnkbOHuiVOceQUENy/lFCKTFO3Zq755cL5cwLzrUQnNdfNb
UqCfOBka4rRWSpwX5yBiRyaVIziDSFpb0guP/LBBR72yw3yCwVvpfIH3C55N
wBgbOBDhurHBx7DPgDhbgZRCPQeZqvKN5hKUOt6U57mxoYl89clyOeKiYwhd
0rQtndKrtRnu1qZhmkdMepnOp6V9FnrgnOsboQKTpxethjKlLnHjjmPxQRk5
Q+1n/AKecdiItDt9y9rQCl2fu0rp2yRLYVNTDDW48PrfGiHXux65jlGpfblR
Ti2bHQzn61ghTOhOyZPM/f8xQkKnVBQh9lxjSSsfT1MNXSLkCAN90ITRl9LF
o9qmz2BPk0WoM5qjizqDLy3RcrmVtKnG2mdS2phtePQiosPphmQ1mgvSnBkD
BnGTi0CndF/5kl5Y2R0J6DnXcBNLmr2lN2UfCbdZZt7L3+XrXWGcm5rlZAlo
F06HlihRpO+mZXB4Bvb2u+wjbnT2KWDo8IxvD3bjW5QWBvVw7qgJ82wVAY2F
bfsT+dFOb08UnbaTxI4hZQF1hIYVqXdE1KKCVcXa1VAk59ROns8VjxV22l5M
Bnf6VFUqtfHERGTioIEJP9inJ7XhP43z4EpMweEDy0R+amgNdgxK2j/+6pMT
sJw9ze/6Cqjwwn4vcou6qHDb3yq8kWUsjuM3jnGP367IokLbUQpkU7DGJThq
INjd+bpByHaYML1x5gkkgTtO9VKuPZ7mLEK9lmwQZ7purYqDmsElUuXvu0Jo
1fJNA1KY1QCaT/1eK2TWJiLIUMxBscg4f8JGJWNiMCWdoyCwNhZifzpbpZ+d
qBXg/0wxJQnaSytlIUKXrEgbQ4UQQUqGk8MvNXDVvcoDarIddUuyBvvbQaCF
z+rGyj3XYyujnNDDqoW1rjD1iWTus7Q1Q/1YZKPKy0u+uLI+q8ncsWrxZ1Cg
IAGmKlv16grkajiOWrU9E7BAEx46P+FjlxTk0TYp/tHCu6RDNI/uM5bdvdaF
MFWyWNXgv1853mSAvIfTBAt+p7rVhi1WfWVo2nYCxMDVINQn2SC9aQll4keG
O9VR7s/LXYXuMoqzilPBld4BWvHoAR6uRfMurcJKXuDCAIcvfE7jI8WEUxmo
H2W5C2rjjwRnFeSbArPawgp0ixwxz8i5lEfugQhmBhj4RKNEVhmIQpZcKYEt
YM5mM5h8i0K19xQMyY8B4q6HiT18+K9p3WQLzQdV98ZRB6UhX6x5nBpDe18e
9jNPAjxcUtV0Oo4GsG3NW4ijxPm3rgZ4ILWxzUe/n3PSnNyTYaN9Le5HS/SY
KnhYVMUpuF9W3IFVQd8HsY1L11QDPK799da+f85Wc1eg5iiPJVOZbhYcRKMs
6ET0Lrqo/Jkh+YnHIKoj0bOE5vU8GwgpNNiKumXA18cmoWzzbGLSurHSs7jb
CEHVAYFH7CnOqCD6Vaxh/joFGxvage4PtNmcRgBvWbMA12IpX+5B+/kVOUzY
5fjE2U1wLGc2EXLpAhpL9RCSAOmKW37eIng10okJlU6NOuN3yB/Vsz6o+UUz
1uPnAXon082/5dNPHuzq4zoEwdyJmYiJMVt8Q+/3G4TtjUP8ocoKrHZQ1KTe
dDYUJB12mVN5JY9rrPl70Rx0l6Ik4zBIMIPvZqcpIkwG5g+aB9E0NuePc8Wh
kYpC08jb4n/NDMTJ9kNwIiCWMln56KWCxqdszuaR3OS33Bw8fk0PBqhU9VcU
0/aR3edRcBqrnJFOF8U+7Au9GJzil4Op+zR38RPEGTEMGrcQvQWzRRGfy76g
kvp6Nk6MaxcLHp42TGyR/p6ALUNdWDJyFEqgvf6zuX7bZ6l0VWA8p0A2Wo99
jEtkMSj2C6qJhHikj6nbBNTco9OXLy/DizJjVAp66SFJc24ivRQ8VjMVfNVZ
F5VZY329tli8u6aDYQB97/C0Hq3RfpzqTPlwUdlwDXZxLLFr5bSxamtvu+mk
H2f34f89bmUyxNuHj45J19Q2HOJMr727IP6XrrmVsE3mamicWLVeTtKaLJBW
yQlXON/V3uJtqaVFxOUru+kuSy4JdiyMQzLdLrW3Zhjz2swV7MiVqLSELHH0
vVjj/B2KrkpfIKOHmhFEVR8Ik6xLA4gBrIu7z8TecfISODowlEZB2XBnYkG+
mdjNexdoW+GADGK2LhmR3RAwNa3UnCZ5WgOw52aC9W+G999neqpGrsiuWLWW
DtOknuiiU2TDRt4m+rnxABL96eU6AFeCQB07heJSC6fXNXIMFVgPYQ4Bco7U
a/0cmCVaSwEQn8xsxKt4zuIf1LnE8NtJnlq63LMAWA09OKcs1z4cpe3obmhc
c9ASelyERivZ8nbIR5Yej/9jIUUqv4y0rJVTRBdVh7ZwF1TqZWzC4K+sr0x5
u653zvTm7j0V5wo3IFYl5iV9s+dhOHgZhobEedhG9g3wPKeyHOQ9yFEKezG4
3FyiHv7cJlWDgtjfwH4o+DsIskIf44AhcZXmMnG74OESA0Hu+qcWdzdH+BX4
tZM59W5Tb+9HhLEMWmdraWd6dQOAeA8IP8pQy9QRGLnA/40D/ohk1g3ED+P3
6w6Qa5AGg1SLPIy8jNZNEYdakS7lzfD4TXC1YLWetn7+T+9FpxoL/F8U+nJl
NphlfrO9l5yvfrW025D4cM7/7DJYGWQyv1C9Nl10YeVy5epCof2I07vBaEHz
R4tXoqJrD9soWEO8E4Cqi0va0mjogZ1/GUWoDcHS9KAxxebu24XUmW+yyKWF
nP8GIrXhw3MDAknMXHESeQ+ylXS2+RFtsh0S1waZZHJSYPraJEJsU9WBipdq
0biBq4f+M/DgLGn+ySC9jQeROkbtBLRkwPRwGLg4/9m5XPsq8jI9uC3osa3q
Q2ypozZWwad9SfX6xRJMETz0vcE/5sKDrz5J5SRWU3QjayDnEw1bt0fUhlWI
ROU6cSg1E6pz4DG5FwplHUi3bCyJ52vzJ/OlGskgIucHYKjsuJIV7BTCHLuO
UZve/YiQsK20keXT/WFbyC0GdjA95hS3kT5wKum9AsgLRiyvmFCL2feyZ/uC
KKv9cN6DdHUhDOQJpZQAb3bC5Re2g980Ed547/E8u5+Y032zG3LOG64E86PC
LvWQSM+zLymlFwM3kpKItg+d98nVnY9D9fVmllIe39YUWtp5BkB2Wi9NfK3n
l62M6p/TUH2g/CcrMFaXmFFkgXDOoW6DVaZzG0Krj1DfKVNpm7bLHbT/Mo11
+XUc9krEQLIQcXLIrUxrHEtCUSDrtg9oNNTz1VIfvpB1jIsUbmdLkwfark3E
0mDcipqjQK5HDVCcjWKBhQVS7L2k136ZDghwp+sVHKCtVrx1RVtKN0jJ7eRj
aVAe7bmWHcb+JgT3D36qUce27v9GzYa5cYm+W1UvbwSFIrv03ByX6IfrqG43
ZOtWXnFz3usKVPau/H7MhHEJTyglPlpPoebeczS/C1xsT17IgyaocCEfrmsW
jOgx+Ildh59X3ymG9OCNyFx3vQpOMRGIgAq3aLg2xVCzbPCKxDweVl65FmVn
e+ePsW1umLnhRWcQFKwH5wdrfsLDipNttBv7noMIrRbROYiuKRwEoCt8MbX4
zsTP/luXAtzBy9hLmnWFx3VuZxLFv8Ro+SPgXMdIMkqrP86jaLhN9yQdJj7x
Q150c9CMkD4NCTrYaMQG1Z1TESq1WfKLRN1YRo5LD5LEWN/aa6Xyj8YnPdcj
RzNJeamIbjSTzcVx72/q3Mb2AgZavMo6tnI1CEAlNPg0UEm2P6tof4GYgZIR
AhPHgCRaH2XF5IPGeJ5czFAjb96FGUrz8Pl1k05SxHcBcn4CTJ7yMtvl0Abh
qczi45PYS6XGaNBJEf+COgZWi8Od1WzJz0Tka5gEOUfsVJtHDrg6zwuusVZw
+BysEGHcECt7oCZakQZgVPyGSSBEXv26LZaStRB6ef8O7EQFHtscGDHRPQ3B
noEpYDalvosE0lmRrOnmzJ+uVQvUO4DN2REJAsAhk71UD0yZuam/foxFWIof
XwYEEgAzbG6ksoZW1ioSE//tCvhxMOQzGbQpb272ESvOnsRjF69w6gn+4yu3
0J1wxz/e2S85g8tgqqWRpqchrhp+WRfvTVh+di9IkE2lXuUHhwSuX9LWHEF+
xPu7oe6pV2QfkRIA0UhvGdD+YlzzHLl+md9A4yXOUQjmpS1jJlfXJUn5s2ch
tmWp/Ux5O+OETrRrxfY3wLnHVZN5Qbtzt4TjypOWJBjTPkd71PbURJM9G8pq
pAdUjhs6M7qIbPGn9MCUshE2Pkn3aVVyAB94hXox6jvJujeFINZtks84Yiug
ynZIs/1yf+DmLorZs798vIG0XNeytawmQ43Ht+iqetnGFETC9+fzLDvsL2mS
YVpNrMnOY6XAB6aZbQY22XWJVEYMtkClSVsOpitiWojjNTC8vANm6F+7Smkb
YoE7DAgKIUCUN+DB6Bp7tMGulAH0QzVsvVPOZgst9xgOLjw0VXXz4jcQ9D/W
z7QB51uuFBW3T6zNwQXH9nb0rusP+hYitSwtHT1OZZZn35uxST08nvLk+9cu
D7Ay/INPOe4Ng3AM1b1SyAOGeZZ+KiqjDGxcWLCcNGoZFyrmjRI4/RiTtfYz
8zkKqfwGV4pHQ8lyf8IaBCgZOG5vbX3QYWXQSPOzCS4KKZXymJN5xAgr8HAh
hOad9BPD/FmhntDdE2WYL4aXFQlthWZ4dLIrNzaXGHbeKgCyeqzBheFppU1l
ZKWburRnCDi3CgPbtHwhCUJTHLZcLPXnLmgEXRhamm01VBK9ZDgzv9Fxe11Y
K9xraFfziebDGfm7/IfJ4MmDKLNcHfwFOxZFzRbFgPglNkwICDjG9DEhrOEm
8ix3nJXg5e7b235ZuR8UBDhXsRyL95KWP+2GA0Auph/hYXfyRVyUF0PimuHz
NGjY+y3YCRoA1AGq7qqr1BKE6z/H6iZo0Wd9Ic9+wM8c6BxMFUmv3gVel4Eu
3G8tkK4D5FQRhE7Y5fH/aX/f9W/2f5ROmD6lA2Hqm/8u3VfRZUMpznNJPEEp
N9PfwKwXI5fVqrVblAj6Qq8GQNYDT7TecaK7ybuA3f8PVxgkRKhak2qIlfrE
7Sl2qDUjcURhwQe2YWHAykNDp2a1DQwKGQbRsq/9h8Dzbp8RqSwJR3ohtthk
cTG0NfkfWjiB4CHl/u11V/dR1LsYScUZIMWMf6oONKPRc/wGaNqI94g0eGMV
RMPe/8SMF88F5vlBgMwXl2eNVkmnpMoCGgtumA8D45GhaxHkXdgtaTwXdD/6
GiVbqfGwp9Yz/hL1G3ocNvke/yo4P5INQObpvWyC843HTcDT64Gb+odKp6js
KUASOo8BPlSfnhRK9Pos4WRpf08c20vPyKCwXC+uqe5qgXpWLNG5m6cFI4uH
CwFXoLFVPrYxWPNoGOlBq9DEOjcPrRFEyoNcJeE0VGZ+YFb/Fc22j4lJlqRJ
BhH3bQ61KEPjmb9eDtIep4tWIT84u+2PJSkbtK2T7q8gYZYLTHzwSQwkRG92
nAbqxXIZKVxBhfTs+Gph0en6CKhG3ykswDTTaIWTDjTxKqFwNXfBAgD3yPm4
fzOVjQ6QdgcLF9++aZce6ClaOm/AMXv0WcSXj8e8+rmLfFiz0wPyFlMVB+nw
QCwRyYt+LtKhuXRiGe2ZexHlOEcl00kwNiDfl7M9QNvMftK6+R/pW7dDzi6+
k++lKJ2xNwzRtKk72C0PutLjFxtWYLrtuUf18kvLB4XP1dm9GU0OftBaxkPb
rm+I9DBB4lQ59iNEz0+lzKfxpwXfG3dOFlywCGYqYG8XhgvC03FmKdL+F9sz
exXfSXgnFHLhjWOR11p/jbwDs/LJAlRu9y6w0PWCQqsFaCO37YFbKRir1hEW
hlwm5EnXhmAlFmYCe7gLsbSA9oTBPAEmZ2Uxa7g/pwFTaheogGNg8f+RARct
sotXQc8w1o2mzolJP+8g/tDv9yEruPdj58V1N9tS1IuYxEd9XSAosIPrfHwT
ZQ5QyXhYhtcxRET0HuzKkuO/GLbSYzQfOb5CVoLZO5COZQr8GqNnkApb26VE
B+R/JR6Cd35LbZOIcUPUDFdIZU9FEkaky/RQOn3paHNKNKxjg+kGh43ojFI2
OMevIuUcNvfn3xO34XjW4oOrxKvA4/bPZmRWDqOZVsDrLw6CP9VhJNCfilTr
mhPbCwxttHzqEM9aCPzAlIsTP+o1s/lUVIG9gQzpwHsO5FLycsPRPDTptcuv
An2JNDHtfEJSgHDV2qjbuuLZlQOd29UBthK7CJ4mCCbMlrapFWDQhbkpf2OF
a4jv+UPQv4o23tZ2ANGVELzF11K/AuxVGtIbyljOu2lezdi6sGYN6ejsK7OF
QbYKomFDinhglwsHU75pRl4MplP5bGkOArS7SMZ7og8B555xvFElFTix1/Ji
Nd43n3a3Z0Ss5UGnsFCmCjBxfpA6z8WLiLRh//vr6/r7vd4Ct+kfyUBvvpQs
1kn0o1wVQZsUxnSprMxWxINY3fcinLT3r1WJrgSe+EgKGqhVpUuy3ythG8k+
NqRrfMzYn5dKt3hncPQKLt6lNlavVT9WkE73fyo0aKbiKKO9boNrdboA4LGL
u7TWZ2GuyACyCq/x/D2jkweqOoyPjqJUDH/SZijtdbnsDzu1lDwianIulHcm
Iqfa2v0kxXLmb7oiuJvSkfhwRAYwU/LffkuyCsw6Nr3wz5VI+ChWd/TJxqaB
e8p++xGi5YQWK2Lt+MPw9snbvETgn6akucLofN6QrkFZk9tq5v4qkeGH7nqh
k9BaOS0fJvqZkmB3EI7nFGp/hxYQqsXhjCX/tbcv4wgQS8+u6adr7wXzxFVU
zqq7hIdgDqPJ6JgpjvuX+aPg6Kvk18oqkSs2agda74NxDXf+9uI+iou/WS3k
5xN1TP555GkMB2EEXWAqbyL2c6jBu4rqHX8Z27dXZdrhwr5qyZwzqJfq5I5M
E1bEjt7TxiT3Zp1kHySDDH7FvLncnEw+5GKITk95ylQAWRc/R+9j5yZ4nO6o
A/4oN+2+31xmhRQILh9zQPtM25L8LwouNu+lIWyLdXok/L1liVOJ+XZKflm3
3ZOD9vXcPmS1KJUhGw50K95/12zI8voNSwMc9Vt4RiNcOyiWQHV+5rJfh6V/
g0BxEa3fXAM46QXyVLXYW/8FeRdt9ZzVW5wBewOEtNqTISW3aYzlqVxkHsy5
+E6QRweNwavzvnmLvy6L56/CmLtHTXsAbQkQLv3TipQSMmppUN7vx7QmlodP
oi41lX92N0N6HV7Hd0GY1FOM8S8tpCvO1+h5cLzvfY/wbvsC6Eh9S3F/s1xj
g4bXqKSsC4aOfcJJ1UsMFBWxfCSbe2BwfkssSGJl+0zwvAQiBV7uOFlxmDh9
gfHA2wJcv/p9aRDZPXVrhzhzcQ2iVTDfaGK1WdxxG8yRJQZelMe575hty8bA
eqzOcVvUUVE1rskvfT4iPfzMMmp81OH8gGw8TZyHERJtxOyLuCCWMH/CPvqW
hPPLXUThhrlZg3IImpEVNivOIChh6IYXZmTD0Gjlqm1jMwOJJR1iqPrs9xID
SyKEOyvNjnDEUSjYpIY3JOwS8m0efMlu71z+VNoYlrPdjdlFsjJObbWMverI
IZGEAg/onDAX4zR2Cjxwn/CqeaVpjz43I8CWvcvAeJ7yj1gGvvF9QI8rv6wM
GP74R5Ouel9T3JTfGWbXYcZTePCKNM4J5HuxT+bXSSCPoW6qdt0MOAYhKZF4
ZSj20nwygDiyt6loPaI/rIBXACXc27SzFDAiNaoN/vmZkn9d6FVmtWNJaF1f
8M6qTWfimtIaaCzadrOBLJC8OTQ0q8V1HXVBF3Qihk6liHhi8FL+zcH+ZMZj
DiTYxwv2KUVwgYXO85ep6QKPrviFt5eXOKGtOuwxo1CIz3kYS3ceRWRpaCk4
tCh728jGtpV+8GYtLgYYuG51OX2S/w4kCm0pFCIDY+HVJUnJsJMBpqQ0ch3/
z7gyvs5hw7IGw81GCgjbWZyOlb66s3CTEPSm2nof7UAMGiPl90jGartCL7r1
VhCONQeRNvz8OT8fUjoRELYvoMI8rTXXqCqHp1xf4QuoCjfk1LF7y4osokHj
FnohrJWc8np8JIwUOCngFzuMKmZUuCRceMWtTl5Ui/gwoBzOONJq5iQYkb68
+daUnvaLW5UPfKZAPQiIHDupgkuh71cvG8Bgx+gJmF5PViprID3od3ozKBZP
28qmkEQJBtjjenuGXAE5hVRi676HcruxEsCSTclpH9dqdZMdU/wbtv0URTE3
INNT5P2/KuL5KclJ6kQdq5ESx/d35iZ2JAig4BZDNTVo2d+0daZyrOkjM+26
43CBF0tQf8mv4EbW8zeShUSxJHVRhiOIfozxYx6wyGZ/kSaoplL7mzOg24uP
QtxwmLtBQC3+OxmeQXYdlsRW/RqFQLhsY1Ltc8flp2brGaNAO7pqPb2tTjrj
uJKTKJ78JsbHt6u10Px0oYHzh9+1h9eJhUcS4HahWFlJIzy0KlD3E+E11ZK+
STAu8ADyvuZWeov5DjXtIJF+oD9TmzsLbXumnYCzZL/8ERGVL9LX7SGYZmC2
4vysIsvo4PN2HETLNylGAPDliQKMNB4wnwiX59wC+NgiPcxILur2Vm+Ir0Ea
iIxDAkK3GFozzuCWiN3NUKDaA6FKDIrhT/9JP4FQQxUkqwCx2mK6NvR2H36y
od1rwTBNsFXs6NE5j5pqNqU1lP3jRvptwL3KjdgcjX0wjEXktlwGv+5h/RMn
IikX/zcAIuvntYg4HyK+BPb2OVK9q0YeSzDU2BX+nmBR186N0gyqfptuTZH9
mDeqXRKK0ZSt+r3Lwow8TDR0opI9xBD+Elh74gWGZOFldRmqPf60XpRcnqLS
an9Jx+oOxQqwEnJZ7fnMJhZhefYncImPMhcsGDx0GNvH0JetsS7S+3yRh4sz
JAL8nEAHwn8QPIrsa5gcDnd5zAMFD9NPfy0TZntjk2j9SN53Y+e2uq88aT45
l4VvDtuunq5LY0RKOmsuaq3ttDtvuX4xBywZqMh3enS7wVi58yOoPLmdwxqw
YYv5NsB9ftQ6XIm/pzTvyl6enIH+44xKvMOCj5ivqM2BI+UHDPwHDUmq/6b2
WxZ+A0+mXQ7Wec4MoX2/co85X7fp5bTiuFUXUxEtQL9x/O/2uswZPsQPzo8c
VcTcY7zXZE0BqRdBlIGvD0G6AyGGs1RWWJUQqVrUxk/0JnxmQ5dMbyT/y4Dh
7TAo13N0/TqZgwda5O/ARITSfSdrCFivc5mLw6jhcLX/LLfIyNxOTv2rV1YN
Bo2md5WHuJo/EtJJC1knegVYcFEkUfd/TPQIkuiCyl8ih2fRnWhL3TezR42a
v66NNXLvBI0Zyb3+X+r+34aMEQEs+q+mjLh9fDqTc5JRnVgtm5DfUhM0ElX7
eSWUsIcI/qDsE2B8opR1kive94RHlLHGczPefgIWlR/vJ+uLtdiC60g0x519
DA/0bA04F4cDUrDxyXS24zBaAJVntQb74LyyAj0a5fbdj4fZs1miqy6Sg574
byNRVihXG0ne7TISTvNWllh6vojyCEkct+xLoYs+2r8GAn2+WQVr6qDIwhbr
iHz/+PAD7JbSmpfj5ZOimibz0N/QLzkRHgkzYpr0Z7V9wCQH6k+o5TU/AAIn
KeM/S5uf0gsikV5u76FU9KDUSYCjp6xfqKLL2pLfr4tDCRBCk8w/Rv9U5Iuz
rAui1yG808xCXbQtujTkPxw4TIDlvPc/jFDLGElHOLKBu+EBS8TLKUAAzWqx
tUNjfswZsX74Fq9+85Jg1ZTG8WynYVuzn/C1oTjYfbAECKKnG7jhLONmUfn9
sSRsNANbYIKQkuL7WhJUfLp+P0tlwFlQ0MskWkR7xb7naQnQn/0s+4NBzQbI
O/efdtWMkrkqy5ZJV/vmlxl/6btqHnVU6jc+9Of/jmAICke8gszQDJ6iPvKn
VHVoDdksBunc6QoqqZjIvQxMm1xkVBM82I/LvBZnCASitEdUhTt5c0UBn5Ic
Nwiwk5ngauhkcT+vYV8/JmExxlTLTCFTiFUFeNJVlNVegxh7+etYiPrO7jur
uHp00ZGK9EAHL5UAfz0Rv1f4Lwh168bz/l8JzBi8A+RC5l8VW9PyoITfuK2B
AtkgvDYX0OAj9lIbACOpZcnJlH2T2H2fJFASzL931qaBTCJ9TCYJR2Xcspzf
q62dUfNmcYmtDohdYZIc5sLhwnH9VOBYU66Hii4DqD2oPTehHQ1w44Gn25/X
ci8t3DTg3ju68jd8swZ4w8SzE5gyzowC3SvTzbcxZ2xhaYIMsG6SdcqcOt1p
DxJEovrw/cpMpFaRHDBHdG0mZ5YjJBC+5yBs3kAcRIno3IJjYMxx/ZN0C0PU
+gkhiZDsktlzm2DtdYv+fD0UzXPF36xXx79gCIW4BkkBN0wFSEl9dC6m4D72
kSmEGivofW4uOY1ap41dOUxKlsshjJMcQp5ODyhokVXNq5LAvn22RvRl5SMd
eYO88ferN4a/m6QFCU69l+JwCnWmMQBJsYOXg2U1Ckop86caygDjnTrHawe9
+9yT+m5mDir5nWRzbOqUXcqlmR7oyCYgOy7VALSlbzZC7Iw8BFdZstd0ui05
7VyMpkALBIU4NB/3f1T1qdtxuBEIN5h+RkXLMgKssYDuJzDOH57/FYyq0O5j
XEbBCw3xohfCPI+fv8UeZ1+UkkD1FXsiFEkQGSt/Wk040nwV83NWFs9B8lr7
/sVFqPB8kxjVQq2mr+eQnTSGjROPQ62dy1Sy4qoBu+XTaQZ0sAsaFAukVpiq
UOZHYYlB7VyyyNqozSPNcahFvRAr5FJOee/taYj2s6DVLuZY8xXRPLLZ2rZn
iEPmLnPjGe7heluNHM9qhjBmDAuviW4vxucp2FgZSCZ4/CBepW9AMKp1OKa+
kiMxQ5Y6pyj40PyARnT1R7MdclcqIpKZSXhMy+PaFDLaJiPzZUFsKZKv6nBo
J85b35POB8bteiTh/adFmu/MpvUYcrKUEAo+ce4GjemvRMIiE7Y3SPtfee2v
SvLD1TAdyZgCyLkZo+wKVE15DA3C/gvphBwCIx0h2c04+QCqGgdsd2mmr7bI
sN1O7VVdAhAr3MoJv/WdCJxHkX3pEzsZHWhNxKTJmZeqMUhz1vG/ep3nzQAT
LR8Mm1qnzZLgHtX5Gpu9ivuTZ0iJDiWKLp3QbHW9Vf1mIqOWoF7olSSPbECo
jWnP1IAfa6K+2PspkMj29A+VDmPG6ZwRUiUw5AaQJWnGFU+c0AK8RSAUjDYT
4Xk7Pr2GC7KO+GDX9V41iSbMBMv2Xxa0+NexLDHbEFL3BfDMMZan5mbj8Xur
GnXJA9gN1JCJE3YgjOgPBqEtqY7qv3c4n45qebESfzZEWmnE8fHnxyDh3RFY
hXbxLk602OSSWP7jATvtLg37vM4m8+BOKKY29A/g7Z0TvavvdzShwBQE6Tsv
iF/g42USZ0Zoqq9FhlNIbNHSSec0Lj4Q16nyAV6d4fmsq9cnt2w1wKVKDV1H
wgAfMdtURp+jeMYKZY3KZ0VLQ7/BNCjSXAIyBrhxUbP8KfNjgbXm/Fdubfek
zAttZ3Jpeo8OOB0sgDvy81avwvsenI/LMlrkIo469C7E74Y/2+QX5vIrR67s
l6o4a7LsEcmDtWVHUkV8OLb12zi3042kpO9MO+NcoiUgruIfM/QLgz9C/Dxk
Sa3K5pUpGCEoVM2NwKwUfWD7CduXcT0fJvpwqDs/2gLDFIbUQUo66XF6wZtl
OMCWMvh96Sggv0ox3Ew3JXv6AgYJi0S3n16iSVup6V6/Wk3FLyCZjQKvumI9
XSOYwdUeBUCJaQOJJ6dI0wuZsXc6TrNUwMzRhP2h7JsJEV9OZBBDllrGODk7
CzgG0TU/4j2CDxdFuR4pnac9evATWPftwycr8e/X/nAZaix4mtaG6q+TZnSf
AnPfACXcpJR/AejCe0U/vCUYmfQUz7qlRTKXbSHRASxEwkpeBSr+baROQPGF
vp/nmPI7zQvPNGUEyDEF3yOTy3XKpKqTyu+M+DgnTMsMg72ijVigpEJQwSh7
wWQvX709DjCbDcRrH6ypWduP8M0QdylvQlzQ+htF2lRT6WcC+OEZXiPSUL+u
OG8t5cGtv1d3o0ScmwkXgkhDIaJKQn+O81FSYBxLFGe+istXDYB3OwFb2IBH
SW4qFkjzbC5zh+tBqy5sVSPwTqDYmrjsaSaIlm4YCmbB3NnJ+T0Y/SfN2s6B
6+MkOAO+6xylbnFoprNpnokjBgoohbMzNFU0mNosqc+BsiHn6xcEELJBF97H
S/Tc2yTA8sUTO484XJly99pFIyAgLZpCJoo3xoUcKDTsCdwmZBuhxyrWfmVg
NmxpDb7CKtyZv+neOyPuHIwHR+9DKoMvOiaQSHatJsGByuFSKrHNSK5q1hVn
DuHBWgufWgqJWtAkbeJZFTG4PLxt74hTxZNgsq1tDIKe+3VidjvQiDuvcE76
eaJlgFMhp8x+1IQ9WNrjbzPgVdRF0IhhoSw/bCNr+gLNyEtIrVR+e5RY8bq2
59D43dCBlPjaZbrV71kZL2by4d5itvt099GAsJHiWHkLQGc52bpOlKEDSVES
HDnzgIEKc9HmTDYBwtOwmiPZm+CQ24VEciE21pJvnm+jyJRiGWIoMTSKztAP
CHSvJNi1dYEH7Sqvg3N1SU1v24ZJsqdiUqvki0aDJgrLUxkOFP4j9ks8QDgl
imddO7pBKvPJ1f3A9PoVlxfkK6E7UYbhyQAGFE5WVCQqbFsz3WM63usV7dwx
zlWs5D5cYBeFI2GT+q29wqn4WQiqwT+jccwUZSmOjhM8yAS/BOH+dwCLPrHv
pkBlnvBPoC7q+GTaGhAVhsqXPra3x3hG9WWM83JkAUnSXwaRlCp2SHEgF7Zn
QX7cPdTEFuTQBuDuzhoZEf+Vql/9VkJGbjnbrLO40q5sgpA6akoCqOtlOksJ
whct3+D441kMs0wxQJsNNwPNgSBSC9Xh/udIqgXmKAnpnELe1DAWRjip/4Nf
rmfH5Dvfl85MlYzJlIagb2UZyaA5iuHNAllk9jmKRrr/PSTmxgKJWrgYbcGi
Bh5bi5rzK+rq4k49pVKPXAJhJldGaMFLu4sp4KNPefxqV9jL1wUX8T1OutYF
/Dakm5pz6hghdwS9EU+6kNi0IfPw1fveDH7zWTc000HfbGpGkLkNkLZlsDV9
ZOUTWFvQVVSuo9w4T3HRWHipLDL7H5zWf/oa921xXTWQFOnoEY7sFexA2kQP
ACtaw7V1HBM569Q3w5SKLLGEgNoKrUUuu9t8JvZRTAGnzhgN75WVGPw5bDgC
trjc+tWQmsFmlno1wIbarenZm5OZMe1NAdw/jMvyDZG0a55h4oujK1gtuvef
v168DgWWSb84SlG8IMWEb1TW6Zk3h+tQBV77FDpH30Kkby7EnGC+tBSXq9lG
ckjz1q1oDwF1x1GU/QWgnjDFzQ7SnwX0FpCXh8qeZ80CzknAVJLBL/O5+45Z
1DPKzaenzpsPhwTDzYGpETSQ3vWNFuPdFx/EijXtZMRHhKvO5vIRJ2DXZB7v
xa2/yAusG2/GCvYfzGWMAF1n4EFcVSjf5A2nLNFJAxz4KNgmxExT/iUDi5hO
QS2Uz4QJtIWwPlrZz4l2tNzEl3QFJrCcR4uUe9IH0IxSpSkL884tuTcQfJv6
55zEwAJPPBsYhuDpTnFgg6IH0MLLjvGZcqVlGZn10t+hPcMCt1XOrwiPiMGH
0e870G6fubIsDx9wLAXHo7jrXXnhNOqbOO1WnjMEVYXfCdv6P5ySlfw0nq/F
dokkWcB07DhXPv0q7QZbLg2GAvHoLBZdYnwrWoQSMS13jwZVB26akkaOaQgP
J4INRfYsJIVtkHi4TuBc0gLb09y4hb2hP4c2HdlLlxyK3brvuhwEHCuwO60p
0hQ3IU/aGFVbREZhjoIBQf+5eE8D1EBrWiAwWwa/bynQ9GnDN39xiXNBo7pW
oZ+hW12EgpkoVpa4U19pdvAfekCjpwC4aKYXyAehtJFUKTuavSMHAYRHR+FT
3MHutQ5BFim9qZLYAASO9oUn0z2RZuM0Fehm1rsV7msQ57d64pt84K9j8iT5
xau7HIdSlREj2lJdF+2+QiLQTr+7iE8zr43AiKS2Sk4MHNj564qCy7H+/Ia/
hlysBm/YdcBgypruteycrUkOzMLYsS9b75tWMkgLwMHvAhXKZzA+4OIoumaH
4bIbQ2lvjAaJMiSXY9e3pDjwXWCEB/nZx/Ws+qhct4lWwa6dgGNdXCwwySHo
xu3XfkJaed7+up0ouaadUUOio8mgONwpp7qncLwz7T70xSnr+hSyuvUJPy7E
NaRDTj/hJsS4gzsDrhhcq57lNEVRqNT6m/NC2bSAh79TxfU0G9ZYr6vJH+ee
/TIGf4zFJQnnEi3L55114IeMIdwsvhBTdFgzwHMY2QU3gc7Pnbd17Rmt3emG
GU8sV+LkIAtxyz5TChg0OBIhuQnajYPmss+HB4cUVPEX0o8UUSGGo2kQGAIN
XPPjn7iiJtp8NLukflf7HN0j2tGo7gUgfVMcxvB+T53rCA9WJsq7WhJQ4Lv1
HqxVKlE3n/ipzFATPNVGqi/3NVEhYsqj4MSmgkFLGpHoKta86rN51BbOT3U2
BrNMu5Vp26drOuEjuPoaN1bnRS/1FDBLjMeplC330m04d3ROupLIsz0EzMwh
a8R6JWiDBTedr+Wm4weMOYKBNhEAq/tRB4nJB8eHoAFlU+jTzTnTh9hSzX1m
VrbSJ7iWZBH0vc8g7KdSDsEzxS0X/fKTbYNBepcwiGo9IpTBsTJ0UmX/I5R3
QsoTPBGXnt/vwfVxg7lInkNPVVgmnP57hXE5Gegx98GwwAOONWvaBhiEfjcX
IR/gn23oF9O54ofsGPt/MQ5h6me51/K83WGxN5MOsNiuLQcbYT7M9CP9D5f3
XHUrxCG9FKr6b5EPKKO3AlzYIGNkZOu+IGB1dSIrvOB2Wf1GIJgC7DHfzCzC
2VEVcM+rtSRweqGPJz2e+GSk5SOPPjXzgUIkZtb+UP5rKXtErXj1JJhrnpUz
y5CgJzzOHuRI9zKoyPnHQD3xJcPh8+ZWMEKLaxZhKLbDtVwKzKgqhE1pRT/z
whS6jp/tovOMJtNyxYseWrjLvv8IfhQqF2Pz3L1hl59xLIRq5cg3ilXItUZQ
Gl53J6dJzwkTI9n1tKROhulyOw0Fov8oGcPgkGN/dj0l0USuVRg90W6Yg10+
L5zh9dtjovAUI8uopgLX+rLF9hU5mUtWCc8FhmW88fICshb8dGqGbNBRHfCo
hUOAjN7cPfRDDmAo1FysKa4y61fZb7JhXJPYKPOlq2ozt0o0L0e0EXFhxgY/
Fb9t6dam3hzhGjvPpYsW6YOL7CgEwV4YyUE5gQ+/IHGQWagyE2TG8aG7Fltx
KM+3F7E92DbJNENBo9AC0GYt61bvSvfoC4IsAJR5l49gNCjInjLVpSV0Ulqx
zwB6vPzx9SXC8SRkxleYRAoS0LdPXJ3M58wkvre/vvADEwFS3Cr9M4U+TUCC
h6H8p9PnqxaKUs9PmuHWQGfdL0QYTpEcrem0kGYwnSAGPRFPM8xUNFv0YVvJ
5f/hB53OqFWuzw7deR0mcIZxxLktB0FNeObRWv/8WlACGANgu+C4awQ6L9Pa
fLhb/Mmb33JUYRyTOHDX9qrLd20eUbxs2MCuBX6T1AbiX4PgusALKEwe2jSi
Q8Zh/+YmtZdA5xvOnPZh2Wou7Wt8nUJDpyxdnp7a6zcDGdiYi2EzuubjP83H
4dgJbeDPm8g/YtaPvIhtMG4m46TNi9yRX452W2zERJPY67DG6gYkcQJGGWKw
VPqWs6vElo2kEwMInum8/NaPJsvFEuGGTMhBCjxbrMDQQukZn+TfqguUz1kE
7Qe6FCoQ5tVm2W8LqDqHiWGfM71zjuDBgZ0KpOz7ziRGln3Ti8tuy75z1RHe
1vON3yLyqoBST0paKjm2g7FPmNo5PxeaySShSTOFqPQhGnNDW18u9Vj+EnYd
4ozW/M5DYe6AeftZZwt+Ev5mTZxo2Hy7+osp56Xd2Jc2QOjV4MBF08dMjoTP
i2IdGX1HBT3ljdfs2zAH2XM5mgtnkOTLJTXTJ+W58xO5z1X+yT9GNZ/Lyp95
n8aX+TQP4Fow8t9759WCFyaFJXHBGFC5Bcvpz5VuLM7IysmmZtj24ypCmXMG
iApYSDf2ETVElvyWc9audLTWhA+uTqpXmjyq5aI+oh7Jx0P8Vy5hajS/Nw8e
eBSCufgRQPGQ5/hM4XZcqi4vShtXFbT3AfhJeKfE7DZVHE7jlBL7O9eigvVH
JWUMoLPnMfy/FL422895WTd5XqCgeCFs3s/QETg7IClxR8dwm3E92NyavT8c
nT40VvJYopxPPXHFGg87n5ZerfcryZ/fbnpz9Ynk5YXPCCOaBuaTso1oVbLc
17mjqOEz10z5gs9rJmj7GXG/pT4Bic4Yo2eilSFd9YdGhDKAPxZa6PJGkJ+I
2XtvVF0ZcRi6rha/1TU3ZJegC7/WApPWDmrFld6XID2Mkh9sp/v+Z7bzfu0u
syRBFBV2KnLSGPeNCQKc1kNhhvyKbvzKWR/zzHgQqNMHaP31OnoZKC1UGl9f
aalaSiUi0Yz1whpdEq5Ae0FL9bGDiFV/xtwwhPCe8PYcJlXEvf6bIGNPLWg6
vsea9ursBch6NXI6yK9hjFsj8kuITpOuqYuUkIAoQSKso0wyDRutMJlkNR5M
vhtO5Jf/SSbwU2NpdCtn11p8jia5JypW1bVz0uwKlf9WqxwF2BNwZP9xe9FS
HVU3sqDujJOdh4vYchcQ8Ba7SCVkQ7xbf7gt19xTNp33CH+6KUtdNBS89Uot
XXjyi+ia4UPbiWHYhUeMzH8Mawo8kbseJ7irnrR0cuwF3QvV8H2vJaAAM5DS
X5dkgTDKNuOZlFQWMpQ1pr0fyOd84GlUUfDkTKlIkWDZMLkVnBAeWeNVXGa2
43gwx0hqnqe90d2IhuRhtfkpJml3ixfkHxnbIsOtK7Xj26ptHdL6VdAgBDSd
4/loeCwlyG0JLDn3qJA+coj1HwRrlgtjQFNa+mHYVZx2v/eSZXvJd9T0Xj4M
OIk+KO8ViH1QDlbCVjPI5Nb7UaWk+h9WNYGODoZzuocn22h69n6nZQtQuLOy
Ye5if5On8FkawEADDM7YhFCB+ot66n53/Uy/Ei7KvyWgkiPULx0nVXCT0Ee/
yjurO3dU4osxnJ2haaMLVGYH2lpYtATo1k8Nf5/e6KsynFgpOYlpL7wDoMMh
9WvD076HC5AojhaY86veVCbmDkDBsWJE3es//NRW8/Krjz82F9QGo5v83HIt
rqxGSrkFfxMJ9qpTdPaQIGknJxXKPwpu+B7G5eGTr7agakumYNfMEiyaSGw6
eazw0P/QuI0QuEQucBaKL96ep4jZV/SGAzTqXckOjCMNLMCrb3kDfLrJNvhB
WQKhWaD00X7Ql19C4W6U3q5rZe3zWxRUIzISaJIlkSXO1E42Cb+EzPJYd9IP
FTf7exs3yF9fwZDhmwEYMaeDMt1VpQHfVxP6rAcvXMmGyNDkHxS4TtGnQIdY
+HBqdA/5zZkl2w+oLrCaKLvv1Y4I7EJTSRzrkl0cedgsmh9CTwgEb1b8nf6y
yqmzgXsqW84MITEnWIb7y1TmOwJ1+xmskUkiP3wXm6ExH+E0lbpnG06B30Lv
Iw9B7rNa1E3dkIrVrSf3hFag46yNJJ6JVNmsrMv50/6SH1Hyfa/vuO/4IX2z
6XxUrzXxajWpXNSs+8ghfTmVB61IITGgWIiQtp6kTZIxmnMuAFD5GYvjQvhO
Kvevg4lVu/wZ5x3ZV/xkTPTcKaSjuyKPfEs8z+8X9B/NlXqbF5Tf6otuX0cl
XbWiGje9Jf6KUlEwhjmHiIH2pnNja34eqbSWQmL0kJWw2xPYGRCmaNbX6zyp
oV8H6TaxRMpycIF6lIj3oQyHZKwhLiyA4AN4lVO9p+aY2tRe6atbHTtEFpT7
IRUCMxO/uKiCIUkFYLdxkf22d1XWH48Ib/LWSiYTSBVjR65fLozbqF1BbOnt
+9iikU1F2orlSGZDa46ePqweh7FwibercQYVwTQ/9xAi6yTNn9kuwRZotXfV
BeYp71f6zYJeD1nMnccePP7oRCLcjp7X5F9sE2mx45WS2EwxdMOoLSSk1Kva
v6d/+CED2HM/wzaKJcjfxezzKdxkDLdUpl30mcAmZ6g7DWohyxY0kv7KKlWK
CXU/p18DQwt3V8VFfWYwuKk+PdpeKZBqCyYpWTATnAG5+x4h+1KIPVLE3HB8
/3fO9f5EVYpLuW9zqGmOSMgCKyiNbNYga9U0Ogbq8zYPhTMcaZxnob8sE0pF
gX4/aKApjGJVIlqer67DuHZ1/hbyOaNPufLOESaBxZMTKbyPK7T8X+tzAWPs
jDdx35yUvGAEBqNEqAo8djj4CZSl4aI6ivMqvTaEbK3qj7eyrjK7mRY5B8mJ
IyVc9K0A6oc2Ewu7+KnSlCwIE2vX9uAXVk2e5oIHLNFu9/qlNBP1nInX1Ii5
PTmZ8rjR95NVaugteleUAL/bjAmQruMEUEfqBVGb3bpN/kGxRo4+84GExi5Y
YPB0XQ9Hrm4I/vDEiPAYzpO8OlW65Szi21a7bThRH/Ge43+EyOfTTYBKjFtC
eQjwj+DgHCfr0btbrulKfqcVP28qH2y3pFlCA1OdlldZZHuRw+EIvPUmTERp
FXBljiW5P3tct9coYvt2+gKfTfL8OZt4aTwoPJ1rMgV2OKMwC2L0nA2eFGJP
SYhMv1lLu8oHeDhS4tyY8GpIQSjV1MXHAd3qx1+/id+C+S/7Y30vcXqcuDxm
6Uca2w8CuL6Qa7cU5HAEbYpbH1bO3VzqYWWxfJ03Cr0kEXMMukd7iC+T/CRI
WRyJL3VQCDSJbhIdiq0QQjiS44oXrqaV6+hqlasDyCrXnzMAurqcuc0wxjgZ
xviFYGghcKt94VBYP80SPmR/pGkp9Mc8t582Plo0GLDIeiXHh9GxH85NZk8v
OyzrLC1OnpiNk2sCD6Bjt/Q/icmYqZhI+r9K7Jngd+02zXVs8XP5+16JNudF
M6UfWJc/j6itEsNJ8ZbVRmAtVB14Wis9hpkSF+94Xxx4kni6L2pQ2S/0pgL4
ox58imhhhoF4C2RSWTsI1ZFROBSGtsGaubUwR0Y2teyKCCrRS9vRrfBXAfIR
M6JEUmEQCjrp32h/WclAm9o1j0NKi1rs/GH23sDoQ7CkPU2far3F4Sh5L/iI
0VxX7Wojmd0trDkPa7kn4u6eTkdVca3FvGtjYR47efevtfUQEFedtfsnVEmF
3bhLVvl4m+kTDAtqddCrNPqeMUjuRsWooKwQMbtPAgLHGchbiWUo0CPqv5Go
VuuqdF37Fzwuu4EzniVkS5D84ZJ/JTXy8NVyY5eZQCG2ylffcWNI29cU4KY2
5nLuIbx0SudEDCfSHiSuifhuPX9lnxV+bWBjtHRVMfGNf35NajnlrepmALWQ
Ng4CciG8JoXXF0GYTRfoyImYzJo9EB2GLYeOSr8+7UL4HPP0H8eP5UpEQJag
2LQCIomoRm7TrIm3060d8nbhKLbcb3aSwHysXFHtDUcPL0bsw/t68PQbBcH3
D7+7jJSvdZYLJNC9SdsOahj4s1BfsOz94hqeLiBCTveU4QnFh4WiKvBHoi9N
fp6nK31dinYRhY7+cU564i9HCQCBxmrcoXLoBX7d8zhW+acEY0GCLW0UxLIm
UdgfgJMHuWgSd9kY2BoIwvQxpdOxfNLnefGbGXz35pTRgjdybYmKLFTkV6TW
D/Vr+YvMXB9bryLOBjiwUe15J2g3V2GvUeom3OxsWXq5FXXdkj1AzceSAUk7
V0eFHo54pIxjxd2x/cxPznObTizUZzDQy59AsAwdJG1juWh/LT13Fkni6azH
/8IJsfP2e6PxWchR9ltfMDfe8YAgXIkwLoLb8NyUc/bxCv0l1ajYdL2P6xwv
GrIcUkzLRLHCFO3iBVqWUVFwe7uCQK10h52AHAPpUx7EOrHtJeBquHTnlo7p
YtSverC7ZnEDJsKFmDp0T0KRnUuBPIAKoLYp87MXkyARRVA4FjMYHVcFdrqw
iZ59s7tEZFILlF3GHipox7Fa7cDrbFRO5aYefrVK6/LGgXjXUR2A4avNRIBJ
E7glxgw460n6YCZZaKF/Hl7Z5kKKsKAObtg4BLktUxLFN3U0hM80whf+3Fp4
qzgYzs/DPAeuENbvXp6Nupln5lLOlKYq4OB9d/2h/PbM0S6hV/5aOHQcYHHY
xAzAyUAh/lqlKKDKR0oCpNMFqjMCFVG2k+elxpMZjh60tVrD50cZ9jUqA2Qq
mgJf4/tIHED3pLakMThXDTkVYxS5oRCXJnJI4qfVnbo1v/dAiv3Zg+HGe2D9
/+gE8fQWXIEcukZ81ji+bqEixuTp10hG3WVqs+2HSZluVPwMU6ovszHifby2
rU1eXuS322hKMyDk1M1a/u/9kK2qHVPumqr2oBYrB5h2Q/I3G2K7SaYS7+8J
Mu7uwKrMK8iJMqUBlwrFnQlitISW9tztzGA6wdhDQvoDxNdnUAY2YCCfhWwj
kb3BKK4i4QxMBI4NuELWzjYeRLx9oII22dYIZz70PNfrZ74bWg9SQ0RqsTYi
pnEjR91H9Ciyb8ds4Tl5xJn/V4u5UcVuscyNmBD37cRTWUfIfVPAhJl6a4Di
ngcGmgfFzRy2oLeL/ib8Tmy+Mp7Ube4KdREV6rEyu+JdkPwH7B9J3dhNHvxX
osLCtihJm5MDrdysSi7mehTmaANnZruu3KMzk7Wy1s74cahohked7HPoDCO9
9zPTQDrxv5BwOTs6rdSijqufHfsURAEYMi2vTc8/NwDt9wb/Vpz0B6otznip
LK+40zGBPJQiHas1RJIiwgLk4T6+0Xzb5JiBLZM4hmr72KLW7SPZe5yh5Wgz
jqFYCUQ6HnNhRXBiYLhdQ+jFdMBys4eb5meWdkjG4RbxQBABSRvpoeMqkRkg
1i1PmC3J/zNqGjvQ0Gq7LX6QM3BeulSkWH+R2+HcOBSljfEDaLFnJQ6SEgwv
2x3vQKbxWyy7J8OcHy87s0fUJibVqXjJ+ZORqYmrYfxYCUTEkrTbtoko8L8D
OdpxYgzmXXMGx5qiua9KlML44AFtjh1RyykM++/ds9Yb9nWqKTycegdCIaO1
LDDpXiSyLLbZccaoqD/59pty9d3kL+u1zZ0racYJGymjEsLQq4x574gDF34+
1kLwr2dAqLllNYIHaS2XT+Pmz4HHIwuq5V/rclDlIJ1OKt5HLw/mktHqohUv
Q7FTx3rd3Kz0JhSTq/RPuRV5E4coAhXy9GrTBSOxVu9uD5O2dUYyv6n1TTZ6
XWDxVsOp5kFK4dMX36bwfXJNCqatZJaX8tj06zmdAnEcLXDVzTtZztzauodd
Hf4JBu64nWvS5Q34uTgDh8QcGidzb2VoG/jovQeeNjee/KE/mcalgPSj7TGA
u3bhkyQTzS1GCKdiv3LAWt+JELMZ9ljEGSfBUUUds7dJljio/UPUTQvPfXXU
T7eAvfUDrx0Log7gpUUJUek1cAGgV2mkEfRr2MW/EUy6fakroi+BLoe+pkXk
+Ec4fvBHgW8UL/T4QD+SbjuQCxSNrqPlbSNAPykIQVs/SSh/QRwkkm52L9Ol
gWWJ+8JZbwa+shfReAk3cDrXNXjhWJg73JXftYuDiFhaj+2YpI/9fgBNEa9P
wJj/T/DTDpUuNxe6jvvAFXGFusTp4QrrGp1HdmHxiQONdBSCfuH1qWlIUEYR
LVFJ2F6omsG+iZt9DXMGLOkCmhbK2ih0Ny8tn3Hoh1UbnlFXOZrqyMK8DJtA
PDM1GgMrQh68gsarQJibT1yVKp1/YVAg/DCHdlnRrmUye2sf05gY2kAh4xXp
H5m+Eew29a9R6ntUT/rntodBwAZwcSl6WKSzp9/YQmOUuMLcqX9l/fouKwb6
k2IeN5IrOTE5ZoHFvOPSnK3kpPcM/sjB3W4DeP/ZRtfoXG/npWoTtDAjfyGk
C5Zmc+4d5YOJPrdUfRcJPOOeiOml+ykPJBKTiInj2KDIDw1Pc6rALByhLzJq
3LwrSmTxV3hvIGFnJ/apOsfhmP0XHIChuqN4EMvpmvM72VgkTHdj/EEekr0B
eiUbyY4YrD8HjVF0ZbvVLQbYSWcmOf/Bb7LK3gmYRweDjta8J195GFskZkNO
X971fygpV+T7VXN4uUCXT8YBFTQlEOsTgVH99IvU4BZzygW+BJK5N/MAU1Tb
EUi028KFzE/MXu8A3Z62tMX/jOBVf2KeubZUJALV9SlEZFQQMfvnX1DOjg25
KAy/Gfm+jtK7590fAlDvuqYDQ2UjD+xfSdW9ZtdofSLeIJyAC+Rr582sI6li
l+Om1EobnSrZVn/bFzAhyUgaaKMVv4DELwe4J/suhc2F3moYtzxgqOibrfU1
nFnNFBER/DCA/UkVXdSNPm3YvVceJxHfmWrSWwfsJsWiTkI5QVRQqkWV9NjP
h6iVsXKGOpxXffUI8VydJf+B4CDwuwo8BlJ/NQYaUkYrPJNIRHpNUKwYzFgC
iNCQd+zmCjhgJlOqY8yyt+RfSwnRtEZamtPMxA0D/HA+kD4OEVG7bR1/Hp1H
AqoMLB+ega5qaxAeYqxvrA/62kLQFXqs5E2aTef63KsQ9+FQlIIy5swIUIqs
JHmIYG+zCurUoKQHWhk2NmqYz/CAfX/xfZdEBl66D98FNfV+KCabz7KTSx0z
Yx2MikcTSitruO7SLE6FL9P8oBj7ZHJEGIc68i1Y1cGLQyKBOKEp8eUam0Vn
sf782o8KL+z5Wmd3i68cctNw00oNwuK42Vt5x4s2es0zwz7uDvvERm1jXz/r
kmdiEUzE0yzAyDK80ydavuH/REDyKQlK3HtlNYsbxehBG4hI4MY5UqQaYfRi
1V+c7UVcqv41Ch2XraXKHHTpkOwniJ5T2Wp/D0Yp6BxwxaEQWS8fsGqyLpGK
p0P0aWqOhWTWJNW/tI42GNmJnN0OzRecIsoZqfp7Rru5cDvgDMa0wy9STcw/
0MTUZA4APq4cZn7KL9UcVmyeHvA3FWWUsnQ7oZb+ek1etaPrfWsT6GPCn3x5
hLvfj8wpC0WHgqVtduqiIwptetCI3msy6DC/DOos8oRtb1GK63Ca4Fj3YMeK
by5/GwDgeCGqiYivKf4FCAfZbSZOv4/HcBO3jrZ2nS19Nvaa2t81fojw0AU0
rNZ+qCYI8TQVhls6WveQPrgX1nfsm4q5blnKePc8GcZqL7lS8YTEFCzUKNFb
HsfD4jpnLOhX8zRNU/iS/l9OIVzA5Uy4JESHzDQ24f3axWXv+BI8OYrf1ZdM
0JF7zw7vHTEOG8gAJWdEBHG3Rla4onloUkjlq52S+IAaZfkzi2WhB9OTOaK1
+P+MI/D3L6rAUI4sAjmkhhUXPOW9n294PsGxAVqhmC2v3MLLPZPAe25Erjh1
YyijM72B+0JDGI9HIJi9zvj8r4IemDb5oclMyKv1rQI1Lse458GIYmQNEN1J
UwNcbaUbbRFGM6m+m7ZfNPL/mOC5/glvtBGIwLQ++GEIWvzufmhWarO5aeyh
ClmmhaNmDRu3UTm21+9PSySVAmWZ54nDAErkqwWIFeS8cnmdCfS6r52nYs1V
mAAgRySlDDFuUld3Hu21sjtN2kM6TlhrXY+bOO4py0yPzPqcN1k22qGIcLgL
LPQVuCD301o9wCv2tsoTvIL+fizUcCMIKSFu5ZQW2q+L7/GFnagakpKkhp6V
JGmHOCLP0ywR8jBhztVC8icQQCxBYsStxse/xzun9a+gC0uK9CeXb0C11O9Z
EveyjA4bO8iPG5VgMTh7NwqLqd62rFNUd7QOr/JdVeoVHehEv8cTa7k3srDo
3hLNs+kYbYMXIBd2Kq++qsSzc8EN3PHW5grF2ZqHNo8t8KhQu817eLKbsZHm
ymoU+r9Zp/GGdZJs36VAhG+6uNWUjICjc9VSnCSC8PzkeLLTsccYFyvv3a6x
uOQr5+Vw/DvUwpuA6e3mK5h/3wfbPoiPOjqHV0X3Ly1txeKd/ciDjSaoCEDT
ZuKxYgnGuIFG89gavV8vCTiux0Hh98755vhJ3m0JI41732pzDeNzjtJbzi2J
fzUSJviSxvhNJNXU1BxrrwcUspiT7aBaAmOkfepPltrUXea/JECpsBEJr0P8
zuCT0Ec+RNlytbA3jMtl12zl6iDxXR7hRJLyQTQ7d7Xsotshf0zVUhlqgcqE
B0PZN8zQ3NhjuzvKJ8CmYpGhKqkm+L6PKDIgbj7X7Q/5R1E2o6g5DwEbkoEI
PQ37AlKq3IyzMOk/9eZCxkJh9yzBsP7vucC6gR1vPOLKVd8vKpXCM0nZmzR4
f23cqJUZSXgHL1zEh/NPIJhNR4hcTo6AfiLztwynXZqkl5nfeeULvxp1WlB1
GeM8+zwkwqT6BkqwvP6RsTplksyvNl5NfoXJ4dsXDBB3OzVkFuSUyVLQFoCv
eMI3Ia9EyrEesh2YClwsvjPXykH4TUUIEPe6obxl8OyTZMkj1hR7AhnfuG3L
EUT+iBBMRxz+vUT/tOhSTgvdCHSXKMxjbmPTGaXCJNQjDnjlGz+f9LOJpQMz
YB6lVyr9NeAHlaoUO7ybzgro8UKWadDPgbNMTxI5i9WERcwGLUw3jAAic0Iy
ZxUmLyOZXsZcB+C2sxdSDXyrXu7kvEw2Rrb917WVMKmx3yvE/oMXnTKXFpP5
ThrNY4zRY9qk7nCjLVCTMA1ILiFPOgZgtzkkc2Zo9LbU4Ztl61xjhm6Ospxt
6WgqOfqOJKkYAvZDmMJ/bdvM/UB63mGxGL8wn0TKOHlB/xlCZXw8NdqojETB
jfbFVXdkTRB2ZpF49uM6UQpaXhHhZz57JqER4Ew1RPctv3KOWqZPtmb40NO9
9MZTUn0uMFNUuCeBVrXNfy+Hktzx5QtWbVbMCqAwCQi2Gft0VxjgCRMNxX1c
/FDQir8O4YwJRNkxcdzMq3yAmOK70JU8yhsNAq3rwkfjqMRLBdEuW2gFcYaM
L+7si1zVaYxIhOA9douku1VIYCUznsbD48L2ea2/xxxwCJ96zb6BSnSiz4XN
sviPgwNPjufZRZ3C8LGVPN3w59q1Lyor8VSbxFNNSd0/93WZZpqb4uh4f65a
a3zhgwRSsVTXa74Jg2ZgkNOXFMBjPuF0eYbYNlaNDJgMz2XH1ARKlkhqxG8/
mrHnf/iVA3x2jRGMRkc+fpnXRvPkhPKYjFy4diAaRq5Uf75Yvz93w4cs1CQk
86XJ0VJFmY0olystRt9s5kYEovqaFPUHKeHd07hTtqixK4XzeFY1Udwwk554
1ny5hK0iyhguHUSiCfAKrX6Z7Nkj0cy2SpLg40zLb3za/cd1JuKre8fzcmH1
ZT3iHMuP09xO8uQ6QqUDd5dSycfz67vfScjb0ZgmTqbY2kVjodRzpL9lzkDl
Y2Q4WtI2wpUi9tN+hLeoJcT0czpYx//+cmmHDMRpHEXlNyAo76N3i4By/Axf
AEm4JkgFeIMFLjXiEux+c2nhxUeva783Fhp8vvo/XQYKfFuhwMKQ8wR6RM6M
tqiW4akvPuLL9pXn+OTOunmU7GWBT06DRXM5H335tNdiE/cfOXfPJ/uhjJ8r
3GqE1eZHQeEQ61V7NIYERQQz/O5PqL8gSIF7Qaiu1UUmP04knvICc5sT9hhR
WTsGPtSP30oPcCZ3pmKcao6xD9CaiBpMqP0rdd6C+nH2p5AqJPPDoXa2uK6e
eIn7HBtsuCM3U7Dgz+qO8tGzlQXO6dPuzhhjhg01ruwdkqoiREgbEdTKwvKM
SXgm3nX7760zgmIgl8ydDGloyjrQRyDrilNsmzC51TZ1Kl+QVSP7oXJ+goFh
A8xRmaKDFx4ZVVaWL31Ad4QZlGSMitmsl4i8rdy24cjxZi2yc8LxoJRJyVDw
Euw0yBsm/tlfITHNdFtO+5ynqepNnOteWFcTOwx+9Wbx1zDeTOP+NMse/00U
tLAXedL0YajA2OBBw4qEnXiW9pvugxSDh4v7SMuoTkd73OV9FEyIvTXBopM5
l0Dv8lDX99gHCkSeIZZ6lYOGG/ptZgkQXE7/0C4OnvM/kUkd/0kgbXjiV6Yf
G58NfwVUGnIyASsMhSZo8UYCl8ChjCx/kM8sRKFd/EYoEvqfPjjuxmkJOKx4
uv6UJZKExRLp3/b+/LiByMdP2uSYDuGkZ6rKRE/OqjOaoZWv+LS+rFTFORLc
jHqdy8Y89d+1MyXXlg6Br5xSb6LMIhpoUXV4C6vhLGq34SEJytl8CX5huP1A
182nhzhThXPtIAik9MEjlPlz2ehD1EYkjQFFAyYbmoi4aw1qSwLibxvEyDcd
TXwvz/4/qFwfY/x8tMQMQrYdsJzOn7QWwPTVt6Wj2gIDtGfCaDlZWaJapmam
xxm2lhRdTdYLca9OzkqlHZPRBFWuf1W7Wj23iYbiCKLLM6VVG/63CCsJs6ns
XBsABK1AL8G7Dpr1gUzUjjVXsLCyWZ0unDSeH2oljyct1FwIdKb5JgPfCDk0
LeU51P/pVyB6g0w2zD9j17CE1em6GT0okzlojY4palNrAlApmGrbHrPyylkB
294WvZ4w7zsXoXQ8GyD1K0xmg2tNKBn6qPxViCQq6whPFEp84Ljj2HOybYSQ
MgxPZObENUmYUdCHsEG4lB1PisevdjWsqNuVkOIBYjW9ML9vhnG0lE39tZav
GJaD0+ER9LHb1h/psWeGz4BdsHuo4UBEn9JA+YM92MyRpvxCRMixEDzOHsBU
Jgclkhflx5MjuFxxKiAsZ0hIq7kA3T8cXKGH/yYcfcnlcBavMdziPveMG527
ncq4WMm195SazaE0bbb/1zsIXnjyuOGqKhk02DKDyGY4vwjO4TyHP3dWWDOM
+yCRQZlhIYEhkvjx6bwn5uL8xmR+tJOAMzeaE/gnBxcuKAkrsq10l+YWEm6D
z4HPzH8nzZDu60jsF48jB9n3nKO0YfgL5CeQv/OUETx65I6x5PYqGB/G17a8
PSr9Yk80rbi/3MM4UAapaAoehFQNoohc7B/rHXW+iP2+myF2m+vJtsXgubzQ
zLSwwsRQKeWuvTmI07y/Zn9fsdAOjgsA7PeGVOKSBVd3Z7zRe3tYCQCGvIO+
rbYb6xqOKBKvr7U4LA1mbIsy4v63l+dmlQe80lzfCgy2GeZ0Ccn1w2WhIIUg
OsnywdNO9stipgBW+94ODfAEuRe86xHOZP6BmblLdSreSyiuXn6dVC/39E2H
TVCihRLBqBIlCi63dvZq0ex7wgptF2Ag+bDwXekXcJK4hnR8U9Oclf9n8qKi
HwJIu4bxvoH7onXiLnJVPMDiZ1cdCRGrGmiFGKhkJWDxo0aPYsKQxnhO8SEM
nVlTG9es+S/uCPvDpqKJossycd40ZDKQl0FG4uoadYruoxvTZLEEc8LxDXEc
sp9cDk8lH/FZgMUQuQCH0vMK+VocGIibYPcA/csBfnOtmMeIYt4z9sS7Lzt6
ki5gApmN63yqjn8tW0LqHAyCLEjaQFudpwXjUDKt0KcSsOojtUhvDfanReSc
54bvelcv5Dqh/Uie1/oxEKMV9vEKPMI2pacqzLpYdv2sPApGWoDf+G/baecl
RnOHz/kgad8FY/cQW/NQlGZMaFPP0IVuX3WZ6DwJBvHliNo3TKPv6PpPoM1V
16ffBxLDwHuCLiEKy9pjIpExAJj6YjJVDqjevIiZWtxdGT4ApSfyPrNSjrWy
NeQZfxBk5P+W4RuygiQ+DqlpayMFkO1wrzqTCufDz4wAgBCSHbFdn2P4cQ7W
DyhtawuVwkgIDCXP0RbX1gbxz57IWffJz634QtwfCDdnLXkn40bPBml/XCW5
VB9IfB5jl073hRvoERpMHHl7WiEJ4MWfbDWiwuHH7FYJodawGWiUXPwnoh/W
MiA+nwTP15wHy73cMpWCYW18m6h7I7BWq1+wDfis52GCnf0Csosi3VkuPpda
HCf79HEx/hvAL/lI534D0zdnFpQz5zkSIwIOa9LeDlPuyatvA2KHA+foT0vE
p2KYsUK31y7BZpoNZxDEdaNlOZYofqTQEzMVOkM3q6j1u7Tuv4Iz8iBoYs7G
E+eFT5BbHERi86enPb+rqjOuEO4SEOnJcpAqluYSVGR3CQEBHOvgbuvcxvsX
GLbLbBhCGBAYNlP1I8ZdGFX5DPxnvS/fVU0sVmbbdDJMIsrBn1kb2gR3zHhJ
JWLSwSJ+2NenbbNpo8Q2Po91f4PzxFd2zGVj1FdPRGv6lZ+S4KY4UYGwZ/B2
knjp3Ab6G1HvMqIy2i3VVkKxuxr+T/y+yhUT9CV6hjV1hcTYVKkAcd+ozVwT
4EahyX7o9jzw9Rf3v605YFcQ+AvpymEeLtRxqqDL6Gt0BX3EfeH/bNUxEpsn
/a73yBzkb8Mssq45+LcSzLJzVv75a+s9nkzXcb3s62XavPQTpuGPnGpmTLJf
l9S1uqUbXB3n5AlRHiyZsXcwWqlmQod2+y1WT5LCasF/W7kXsa/qvvRDWq4K
soVOFwvKjBKvwXcNn+o0FMSHRyUrhHlO9Ga2GturRoOI9eah4kGcDKfdoz1A
3PX/JW9eRkeWSz0chgG1bWq3tooY/dOV0ywTtsI+o7ScYEN2iRZMJz4NySg7
q9D0gSG6CEOYIKvuhD6AWEQWqOGXwj4j/6aLs130mGRkWuUD1KpPEImYF2/6
AkPsChN/t0pxAMiB/vbBU6o21u1NNFD4BcTMuxx0Z2so1pTqu0fvDwOSuNZf
t7nT8xRszM2bF4XK7n/LFnEEDtyrFf/6Q9twH5wdssceGwQ6SkcfEg4CbSV3
eVnKmmykb5N4s7Shd96uyK7MYO3GexXtu42S4KNxKYlI0JuB5lrJyd9Zq48Y
wtWoo9bbI+AL7hjWrbjUbKNdyN0kCqPvsClAftDjCViK4Nc6HwZe9tfxGn3c
9ZyiIW8YfYszYWQG6zmKBfdPx3C1MpiguxSduL2lfZAznuVzW0rNnjMD+3au
NlsFnwG+D6Z1qmicwlrp5ASeNPwM3i+vJItlBSnRdWsywebCTJKjLwwc1X2R
JNTYD6CTx2gv9xPxcKqcO5TaWD5rBpyk1jHSuA9YDfDanpT09dBsywDwAeoQ
m6ZKl6QUvf9sySiBlbclwKqtBEkeumrKl1zwu5/nXLfsbwB9vas9MHw3BXq8
HR5QI9exnPYwpKSMAdyDVCrwMKtIPMgecK27EGbU85BguusRC6/6vs8UO1Ga
K13HVmqhZLSmaMgsvVnc5DsuMEWzuCfLVkdeEA1GRMzrk6z5iUvAxISvbkTf
7lQ3mbIGbvyMlbudEA1QfsTRW34DG1GY76erX3Ei+A2+bJx3P1qCdDV89r8m
7KHfDzYpvgoJLablt7RrJ7whTlSUYNKXZZs2gebbr2AEhFlO+AZPdcxzGPq5
lQkUur+mOWz2Gvp5+7UH4GVuAlmjMlXx99vMkuNVFTjvmAiwt8/xzInf49XF
80A+cr3F57SjC6Hs+2OlfJBo0cZPxMqHdN5oen/+Hv8uLCU+exojcpNYT8rn
WmAjO/sCq2P8nxZJw4sM+2tOQayvKKAaqJteoF2YBmVYoDStPQ2uokd0WrQl
UYdXkEmrWvqpwoLYneVrdGpC4MK8iyMd1TTTwplwwmmtJodcT9dWfYID4+jd
wX1wyQbhFn8AtGaiykdX9aazJdQM0+XegS5AUB6byVnY2TLlIEpGKZp1QUG5
YZIhlo5W+luGaQeURkx+tvGF3GxBHZlkBwqj6ctaPEHJio4wvudmPVN6zvEp
YBciJCCzvebLWDrhYvk7dlGIypbuW7A0kxrXR/8+w4eLWnBoggYr6EKn1G+I
ivVUakk+MmhQpgjGwU81utgPbIPjsA15lUansWn/LQ4Eq+65l+LEjpzKppww
0WaecFrqk2YCT1NQ4pu2+E+8Yn0SA/Fwk73DsFWjFPXY7sw3doqK/wvYKsAH
Yp1kHq3D7ranMVqm5l5BGzIvwSaYcfUfgg6jqAbh6d0o9qxJzoV+p8BytFgK
VqcqrdNgVbfHfxDbIEQSZHpB4booyWmFuL+8MWwquxsKDPWQHHWauljNK/tv
TVykerA6w0RWKxsK5qHFSBW56kPNEf2u+VcefXk3qzy33D/TarLslMIQw1Ql
w+F6aAnDcFJPnmj9YG3UC6vBFRHp7t/hiD4bX5KP4nW+dlV4U+9/CsXIc+18
vUNRuZGVR55iG8QFogPgyThkbKcHiYamp4p5XGQwUfoxKDTNKJB1NM/j7Ust
sISC6UuNiMxQ3uLjjkCQX4XMLkwQ2RCNo800fLH+w+eBK10LWF++n/PavIRv
mn4xNyBrQw1W3nsCHvA6plHipQ7ky7U1myc/sTuPP8OdElqCPJuBEJAubl8d
JLDYiGM/WdHX2kUsFr7N9QPkRUWfVr1BT9fFzuIs3dTjAfDp2aKQAZ5Uvi66
2VJdA41FGj+ZeoARXo6G2HRwoqD91WMrZe6v0ZDli7lTfY7i9w2Tz1uSWTca
ZbZau2pqbLw3Utp9rjoTewnoaRP1+fBGUntB9I4rt8+CyKBjag8qxmOPLV8b
BToSQTY/m1VtMDFbaK/Lsd7jQIbfc4t+bgEP/vfuymRh4sWstFxpFzYK/Um8
SGny1IDvulegNTHd7FAP2tfmxD44kBT67o9BEMhxbMHn06eEWB3+X1o+/cM8
xRe9DKYLkRRjPbiJefRd93zUEWMRtqV3Q+wbU25VJJxJ+/3uKH0uFiknjUHB
WSgN6mZByYAGlA7WIlisWM9TdwAhr+D/i6FX/78TJ049+XlPSG8YDu2ChCjD
gOUy6JTw/7tMfNY3S8yRnZREpvp4n2eB5nGl9SmrDu9Fbo2GoG/PLodvGdue
ye0d2eMvSL/ZFFOzu+kiVALZdjMObR9ZXdm/Y5YhE7GDgnKG8FZ6iJDDGPbN
C5CZ+SlKMnnq4KOnoiqd9XK6AAZ1aI/hxyzII/YIWY0yoTtwDFqioDWRwbMq
w3RUoJcfWrDrBOqY94XuWZVyPJ5qajo2NopoAX2wLDUa/vaYadLkyyIFvO9M
3IHEGz0FGWYP7i128MVZSnhVKv4gZTeQ40bYla7fOFZUAVVWRL0dRlv3JHM8
ChREnh5ttTxLS1eZx4rwCqljk8kNjz1eNZGbg2EzpbxxarnFmL8Y3NVYtCB1
6WtnQ3t5tIjXZIvVsNpnVQG3wfB6YYhaqOHAxpOZNDlpsj+UiJ1ufO4F1v6I
RDgAPZ3h9sRbMr3UX6XjiQhY5yCfd6lYKoyLb4wXKb2iYyJRmndyKJYQ/VbB
CpvOeklOcJBovRQwh2sYDOLQ08FSR/OtT6V4p3saDcvQ3fM2rxLRJT4NhxM4
kWMTId7VuM+iMJ71oECmNpW2dx+d7GghNtNhHxx1JGsdnwqUNgd/ySbJZ3b2
+B3lJlarE017GFzCPq+Ha1+ueFNhi7HopCrZypGddK5S3OWHzATB85LzC3uv
USxOnDcYhVGAypg2aEW7SIpl3Oy3+ioglbgvr+YG+dFXrm5miRMuIWbV3s+0
RzE/GNn0Q18XhQ46KOUZQJK2+A80/+rP3I3lZo9DCVgK1CPEC8zuHcc3NGIb
2Sd2R4+QfhmcFbBcicDFNHimXK+6gWGkDd2hK56kNkLG/i1gjjiEpHXdIp/b
YCs4G3wFpC2lAHfdKerF9V5Gcy+8G5eu0Js/ZMIwySYvxnU=

`pragma protect end_protected
