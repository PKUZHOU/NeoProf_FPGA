// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
zuv2KNCclOZvmBWDuBvnKFLRHTB/8KNl/zCjRLK7icb6cc4bbG2gDuepg/6vM7cosysA4AbahPoW
2ScxwJsVy1ZTDfgxmyA/3gVVQpb7xo9IVznZkfQucdaqKElx4usFT3UQQILdkCBKn8zxM1CINUTB
qyqms8Cnmqv1WbhjbmmQBHK6Km5EucFcTfIPOKY5GwjplxvWDZNiaM0Yzdd4YkRaUqYfYVVEEG1o
xIDsDmdv6t+EgEwVHa/nhmo3MwtLDsMWUzn5kg+X4sPjWRwOpLat2RKFuUVbFNdWfO7HPiPW53Cr
INrI8tCLa5B12YbNDRLd55SkEwfuVVTMyJdsAw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 10560)
W4GUB/AEc/clryhXBABwxwCKwYGVPldJJhBt6sQQYRGNDWL0qLA3KnXzji/HRKwtw+v/il58YLVl
jzNxvloH4i7DZDxgAGDVCQLs3XHFp+8idUx9+dorV4timEtdg35MSL2sTB/QrzzRjhhNy1QB81qT
BSBypTrsAe73E87IH+Nlu0NoARvZem2vJsEPb7sKxcfR3tpqpRq0LnUIKKnfrUYbw/hsc298bAAj
pnwNbL8wzbFNhLaPQDLfYKXpRgoWC8RJuH1sxp3nkmaogD9fo4eaJkwyHUCeM4RGqKkwb5wpnivd
LXKldXOcUcrVK94tFehaqkDOC9QAdI4Ln4zTH10IDjQvkw0i4J+MS+JZIfxbaNRgJwT4NK4u2S6b
5OZjoEg26Z4ozT2G8xyCjm53w0VdQXUEakSeOyeKh7CTvo+m41NHCque3dAlRr5qajDOMbuSt7qx
HZ/P+4XgGfF+t4PwFFSo+7H3hNDAbodaispUPp4Dv35mu1zRgrOEp157UlfsABq+ucRokd7C0i40
ThE2DgDw9Ae+30PjHLkIgyB33DSkxV9tAfjG/Htjh6aEGnsYOr7iUhRO9G7GUW80JMeQ9jDoGugS
nj0d2XrStkbBdlcc7ZL03Q4nKVOP5R7KE9ZnnPM3Ujf76BHvrWXrGuN5rUXUmKw9C5UPHxS/yTtv
LqoB/X5Edo4nfJn9LORXdz8APsAJ8c4ekxjseSSdp97MuKjBvWUrJJOM+hcgk0qpN0u08+dgh90p
B40BMC3c2+7HG96Nsuf9APsitLs6Bp38p58Q41Lxrthao3Fi7+HhP/ac4EDlSd58Shp7AGO8QiSQ
iCea2QolABpIlPW+znUlebSZH68tetCxMcM2Q8fCy4I8eE3tK9lLsmfCkdIjU7dnhgvsjx+mYYmo
X91eZc5PdD4c1wXzhbhGbIiA7xOdIXYDttD1Iddi+GmGyzXUPo5gw7L2lL9Nt2qUcliY+uEWBs6j
PIz2QFoY0dzSQO2YEDKqGNG48G7Vta3F6S7z0D95SD7aIdfYnomWDdXwFQ+fyb12g1OqowlUvPvW
Whd5VH2j65+oYT6CsM8Ombk9nv72Uxu7s99wjtpkjVTeO1rW+gcWm+tN8b10LAvG9WKaEk0zsdnH
B4C1Vy033uzENgQp6BcZnQH06+m5PSTZ/lEzT93+m0Hx4Ta9mcfBjk0j1ekmPu1HTUVHcHNBDHDJ
Trpi8+YpuDOFkidQH5nOiH9UKqutluA6t8aWbJ9PPDvcHIBiFkSRWzJp6FXy9CMadqX4NSQP+WW7
G5xzytTnstJMXGp6fzQn+54uZmJhEnDaR/dOtk4vXYK0ICnNJW5LUaRbd/IpAHao8VDa0eGGneWL
yCpJyRydrhukeKqK0GuuBT0iqippFUxuXFIkKRQhuHes4x5J1YvQGBSx4P7DuLqNMfOkTueQvz1b
Xbnva67lfbdvUj4V7vMpMpqR9Pq2vUTlf0x9klCEzTMUz2FQOd9M/SDccYD5doCtosH+qWSYcVPd
bjeExyGroN0oyZ9kZ2AAihn61zpRkGfB2csYJUHK0p4Jc4sYPwPFFgeJI1wV9/D3gWwB8U9QPr1h
dFanLLgjBF15MJewYsw1mJeBqQ5oAC77Fs68ENJfHGbFCIGej+g+2Jug4hAvbk1AUcy8Jm0mdyXr
+j6PmcUahFGKge43JZZLfUJ+bkEfuHtY4DNOpIE1e8KskZnvLFioxtDxsNm2OBeFeytKPm3dd1BA
nVSgPu9SrM+7SUz/4uvxQjNAQgGEUWbJb6wLvO6cbiwE3Px91oc1z/1Cz/iARzGQDuOvRTJobXuc
O0H1Jw3RAJn/KTkwjz7FdrtRBmff+/6NUsnYeDMeAafnaYQjZjxfsPj8ySanCmiO0CNjBVbFjk8e
8H2LDTiS2Y4f9L+iETccbclwWqc/oZdmY4IQHrynqCkNneRxG9wGmlOBrKsXz1ZQ/O5poSOoeQWO
uc7h5chfoAOeMEI9SMf30eoH+IvPa6BccIK4CDhXByJbehuxI1Mo1ozxDnIB/UW9lN7NoB3xMT5P
8YTMLxVk8phOtJpV9hXlS61Du4YNCDOhTDmTvUv4d2sVuCsnNpCvHGghQnLiltgwvmDagtNEmHhD
1wuWDJ+Lo3/KTUjawFiM0m1oE0O9jUCDV/6HQSFdmkVoXl8iAyd0CWEH10CVvQvKq7lxHiKbak/e
Gqjen4RdHHpKf7Wp6wPCRdD3cTdRc0OrbSV20qDjxF/WNHfCxv5zI1A0DdO2wnvLr+c3BoSV7Y9q
w0nWSFbqg9vCnlHSjUGDF89s24Pp/9Qo4lg/55JSor8708k2rCUhOE5KB69x/kOFb3CM+oxEodZR
z34Tx0+noDK3WO9hU590648/3GSPssrLuvAKL1Y3YFQ0srF4HX1llA+R8lQ/LQ3Ku3fyIH1NfMjI
nnYPVoHIigjiwBMGc/8yFirLAWkumCdr9MYKIBefvY+2W+XY7S4JRrf9Sj1TWacdDlNUzz09FbmH
Slk/BHAKjE5ZuR3tLs18KIt1kstVzeesKaHTflUfwecUQca64j35vZXrwOMRYn4V/tjK2DDPCOkI
EVxuj7LfZIMGpEXHHV9HirCaCietVJZatxH8mgwuHlsudQz6RLkxVqXU1lxmf06bri7ZqFC39l6S
MRxXrHkjrYzj/oALeOeBQvEldPhgCFmgvLuMp31xJhbK6fkkj+HQ9y8sgQphaiLthnrxkSo+AkGN
KrXhkpccpZyyMRD7RBsp1lONeQxeDhMukv/nt7poDjckNnY+MG/b+lE0hQyKB2v/RwD70Nj40xhz
TjTuI+/iP2cmM4xjBBHGTqEBvi/qhv87J74qTrNgWb/zWvfqYSio2zV/WmLeSftBvBZOqGI4h0I9
e3DrPVcY6un98SHExUe9ocdc+mIZeP/E+/Re5iEN/h3hleE7ADVIwxB4Ck0X+TjUlQTtyrToq8A3
cQHRCwJD2w9tDFjg93XyA6uAyLZNgZECCQ+FwbgiavUx3jbx4bP3HvFi9yhNLyQr2+A7BGzya6Fu
50/jsSPK2Mfo0ehhfVM8hm5dfzkNX0ysXuWA2WpaL8BRA9evkgvKFziHZdSL04Ho6/9/CxImNEy2
nlwhda5G6ADk9yiM8QBXg3uDg1BCmqafbNB3Ny7YH1KYNn5zmlf/cIOD+ECFfeUHn/JCk4NazEHl
mDsODoTA5ljbiBNNe7wURlJ4h/VI8rf75RxlcPWauDlE9jsTmfOf6WDgpWWyEzjBsa6GUHNK8LUD
gBshsuA5HEI7K0clks6rIXg+kCilw2rDIeLXkvETsZkC3ii2bZFn3bS1+pgPZbk7hHetWj4M/pIo
UZuMyZgLSo0r4OkSStmVRc1v959F9tnB5gmlfqYSC7+tnd+IqRnjoD9+aNVnAGMi3jowLxk9yZLM
EMOuCj/nQe8JwFH2+K27mN8KnQdDI0E85LOBfIFEQToGDa7hQnXj9XVPUL0pdqIvQjGT9/xmRQhp
4ZcJSJVJjYi3e9QAGQ7ZCZ86HdmQ9Cz2n3su2i7vm/5vyu2j54fgEHvTLWkcCglcyoegIRlrpKLR
i/TaFcnx3qMnLsDQOU9twilRaswxgFBZOxaM+RI8usKlOUiKC4KYKtXtdFAg6Ec7cpRsIGlk5T6c
1gv3rIWk6ktpKbeobS+dAwaGnx8JcuNl7t9N8ryi4BwTOEUxoGLH/xpUWNp/dcUcKy53bpa7E5ko
fdwKgKSpFJRXfUa7qQ+oY2l6XbFVZWJHK5Rq5+ptPJ5HekzdL+ddQ7aDFv1BKVX1/bS+L7Z+HZu2
91gTVDQIPV0TJ/v1HloHrg51WytBFoiUSwX4NJn3QiGxbWSe3YlQMXUuLmlK9IPcyIHw6G2/HS7M
t8GqxQSTsPjz5E7CWr+X+/SpNkVgba8PR67fzDfyQOCmYZoyE2InRCWb35SMDodIsXjgnjGb430L
Okmnp4Qxe86bHRple/yG0QhOLhe8h4sLIsnmb2KeENXcdN8sqw0OkDuJfzvnBM9CMma3UwzJYpsY
/+I4rVeNnBcUNqvmnwvOZHTgMOyjti1OXH+HJZjefHj+1unqBfZKlWj7svLEqIhWdYK9f129xvRI
ia8nz/s2g8dlApqYBGf8MJWPtF6YHtm1SuWJOglM4xwO5apArgBCoLKpGrqU5znkdcfHTWAZaoQo
iwGO2D9glKWI3E5ouJmcEnTHZOig1FAmtk+lmdgYIknnKLyt5V7Twe2Q2/thq/ve9iKeuxYEBHbo
p6rUF7HCPkNeUkSp2vQjMv6JbsdhNTMZGqPETICs1EQj12BLz5vH6zpzm7APd8pUmNa3W794shD6
109nvfwolU/F+x6NuBG4Cxx8zDQenCIbf+4F8zx666jr3Dto30rNyQcXEoZYI0xFNquf57xNfWdt
IuaYwcc8hIYOFG+lbqcne20Ush19YhY1VQ5VVVYuZ4KwvoARk0Hm+uqhh8qeXSnM3qO637uMH4ZP
rbuOUrtxBJbUCREM3TtMaTZT2Rc+pjdk5QxvtYdqzLc68MOObVeO/pRQoBX47vv60shb+4f6typU
p39mserr2eq3H5po1X9M9voFPsU6MLbtS4Lrd6DtZpBo5Wd/RD0OJN1GT77Q2kkphc/QT/5AAjTb
aUOdPonc93UGVecgbVcNCZ5cd/7kmo0PCiKzwOxkTREzYbx4cvxxu9BqIvv9w8RcdsfcQ34dJpzf
PDYIRmb9qc9gSDNglYds3fKanBXSZTY/aegqc0Fw6nrDZr2aN4kXv6VoVNw5tQrmblxqEFDMRYpX
LIwlpAVdD97QKf5syQfjOzNuh38uI8Yv1IGzfWI1jTA+4+BTKUzqMmM7WzU9yIRDIzqFkdlG40k2
ptBL+kCHZZIVAkQqTQo+TSlAtlYj/vlc06ie23d3PtwFFTjN+5UVSCZxILaoS7CfwoRHYLeJ9HIw
scEwn3SPuO+m2qvPw7flXAVWMUZoyd7aTtrlzvHR0lgpthpdW9X2uldLoyu18r4AH/zkTJ61e4Xt
Te/O5Vfl3o9c3JPRRl1UV6ykzmHz286bzM/it3FNpQDlm6PJKcni1JZ1/5iWvmTw9T8YeFARlo1/
MFg+PAxoSwEKhYwM6DflusoJneJ+Ehj7AvyVu5cCAJOGKdG8gIupSvIPePrBTe147oEAARsA34Eb
J+g4TNxNBc1W+52Imgsxqn7ivh9h5vsKd2oPHw0d7shc4a4+cLYQegyZAe/eLloQOuMbt9amksye
Bdz/wV3yPCPJuqt2tNIt74wgD9LPQuhjjjDpVPlHEkn8ka2z4bF4pNGBe01QVh1JEwI7Y2d2iYJl
d4RWv3YQVyYWn/puOUKeOve5bZpQV86KR5Gw/ltlG2WVhBgwHO5Uvi0SHCTbpnsS/DT85JO2AbzY
mGzRtgZC3PXQ4jfFj9QENHHeSVOPTSXoY0vpI9knzsXzeE5QYIHt7UHkLYd5UfGNzS719CapV0rY
OOEK883IbgpGZd1crjV/6aFktl8szliZUpkKodyJHXxbHB7f7D50n4svsv5Z/CCO3P1+xXiOpEN5
U3d/umGvlFAVUClEgiY4hdabSNdNihR+nXhaA1RNzcx0rgVSRVpl3/34Vc9y98HH5QVvmfGYW04a
RKRA0rH44iOR6U9qIcoiGtFh4xnXW1B9U5DtCosnqpw2ofblR4/2t2gRS62aID6dA1APAD2iFcks
3rkHEqneLUSUJlpG1QcbFOorgLQ4BFIiDlzJkcmVrHi5dP6nLfTFQmOrNRB99/JmRnoPFkT4156s
kUoUsgdGh73j2ot+xokzmXfwPzTWrmB2uQx31kcvSLyN7SIVk2Jimws8q0HVoiREyy6aOy5LAcg/
7v5DmvLpfep7WIwL87Mn7xWxEuA71V/SHW3weSUdfwJD3o57oXD70tuX82zwHP9DRJerM7/PzEzY
j0CiJdHaUIRKv2X18yBkuRwS8oeMaI20S2gmIYU0Jhg8sg/RK9Xi+1s+vHKrCAwGkX+YVpmsK3ed
Tb3gUNfXZ78TKDQImOO5VjMQwzBA6zqqb4N9D43d0JDNFetLGccueaTTjWOsSePQ4+SC4kJ8fO+l
3tUSeToHgGd1R/hk7PZXAFs2XqXRfOHCOE43J4lltWA7ryd5Ge1TyjdcJyGE/jG1jIq6dZ2Mydj3
47LwNwJ7uWAxuYbHdmcNP5hjL4/4Knrsba1jXaWGCVBNZBEfQM1QRz3i/ZSdEoxv8NLGE5iHa+y+
CPcpflYPT1mkOzu7zxs56bbzoZAjfawtALfLuw+okSdJDIL5dq1Dy5xID/ChKfkK6+jgWgy+r05o
US6seJ6yA3KvnasYBD/xMPDgA2g3b9ARg3WRsh9FlW9uX9O7nxyvJoj4C6h82kQvonCn9iFqI6zK
CMkEoQ7E910EuKgpTsWHtGuwkjMWyI97CsWyVTeXUFjQG6T+Gr4VO5VSHjCCVYHCEU4JSle4VwCI
SqZqnvf+ORsyN42aQxXSWhZI4Iy6/maimPfIghaL2bynOjwVXL5TRVhSmXcj4A5nItTVRHeKAkn2
QZrYedWsDeSN/YBuUX7LMmhEC4zXipBTDRanivY5+pXQhGdPcvXhzWob/FuzSz6UplfcQwkzm9nC
OisGw4kbJY8pa2GoTWfEGtnLkMEl/pzi+YTOA5LnR5vN+0/Xd4evzzqxOyeJBgki+QbE8PzEEMbI
kGN1Qln8ohkc2YOsoNKO2oizvH+/p9f8gybewCvJ+NLn+WEOyBElqnuRsDLhT/Q0vl6585jrZMpV
rhAqlkHrKeNAhbggEuT9csLKhiuoDEHw/F70Xh28nmfrqdg5v+g+J8ARPMHjNSPmn12vK208u3me
e9OYkN1hfy493n112sPaxuulzr4mHqAKpmJGbxZRZ0vb73cmu7it9sEzz88oxgTO89nhA3PULhng
r490yU68TTfzF/yW1j4SybBwnvnr+nIe2IKoiK50uZxPrJQ1yuhKSe3F+1HkzXr/nWg2JYIazp6B
TzOOz3s7hr2rTJRVE1MQ6Fjfa5Uv4Y0PhD2Pen4j8kNWoQEtJ07EeFkBC3SNPDOec7BkQpBeoSbp
wWmdHkNXe/OXwMWo96izi+zV+QvjD+74JutNTp1jGWW1CpieSytn+kpT/u2YhatGYJRbLq7Xhbzl
braUxZt+s6B4qyXXM/FKJZ3QIjjY3eNzPUn/ehLtGT7YQPRj/xZ1sN0PxxDkQXokY3SQeCsmHdqn
2DqVbLrDMP8LLMwyzW+5mJEqFRX8SHnBw7+XPDWe373WA278MfMTsoef3Eqfht2Vxwi5LYFTQIce
G3asSnV18W7SNzONA4Lr7A1kP9sqqppmgUGQWyKg3Ke5MZ18hQwcqU6G+1l+l4f8P+ikwF+cGbK0
XrKLWGavlqP0WvgSJbbfJEkeyqgUaM7GCuHVnD4yH7ZXGYa0x2xC2+NOTr/fVCGYL7kzA0BOUj2w
1KtP3LrhcNOsrR8KQd6bcmx4dZolf3QgHW75s/1ZEfkSz+MVrBFQt++zKIUeMBmCsx+seNhblSrO
OIRy6gf6dITzDgMVFCPUM53FZkb6gjUiOI6hjiYs7yPQEIB+JHxnmP0ZOcwdV+o4XuWAV/CSjN74
BoawGyjQbadHIx2MSVnrUfQArY81LU6XZYkFZUzvYqzJUD49TQbPHsP1kxQvWKywYfECN5lxp/G/
FV4hWaLs6zh1lkUzrIphIwD6VeQgdqalDCwyts0tNlGbXUUdF2ybLfbrqpRXy5oAIMKWzFjQXnfV
+COwe8AjEJNU2/UW2cohbg5hDeIbPgR3qqDWH6gpks1Qf2AD6whfX89DTrqJ4m3yxTn72Rlb7VHS
4KzMjF/WUpbTlCIvMZFu1HNm30sH6hZS7UmTgsdiPwMu0fcVqCsugcN01g/u2urM+A1Lklso5y1V
p5aPOwY0MrieZ5Yfg13FU+bxtabKRD7POODYTk8N/Ixtc2XBIcICqXYK6Qkpq0gwSHs8Tx8TCKas
R1O1UUT85KfYORrHcZgyoW0gc6COM3hoI5RC/aIRYdlJpjGreKjS4ytKMeapVMJkQvZGa3f50aCi
Q8+I2qYdS/Id7Cp/g2LIE/tIeZtR+YJsv56hHXE3v+xjFSHfwqCTG0BoIvptutUxhgpWekgiQOkp
EQ1xkcLEMZoKyHVS+rEOPkK+Ip2F3uFVmhuVYMY5Zy+ReCU2t3OSdhJvo2+OGOauNOAiSJv2C6g6
NijbszmH/B5Z1yLvsupARlr8frdhSYpkgIfw0sFbkLms09Y9At47ufzEQ5PV4UC8qdiRB3Dwb85q
yKqXIqI83Q2c2UhGJi+Fpd58LzBDJaFCLPGTCzxNQid1FF8Dr5YUz6QPdpxPHEPZ1b2EjwLPTdsb
LEKdGStaEx7YPKhPKtqjhst5VqjfksmAODW3EXt4ZLVnHFqOrvwAOYLRRZDT6FKrdZ1RqENi6Y4S
MUvtCNIdj5PhSm67HZKI8EtRagGVkUEepXj8tNR/T6rdu8NzNbMl233Zc43ei+cITApHd5MgkrQK
WxOV9vSzF6jHL3UaEtYAhrRdL95P/FsByspQ/vT9lP7VhZEvOvt/tAaE+u2TGF4mmQRUC3/ge+8+
s4r+90iEKS2u2RlK1f8g4NQ6KSAOvP0G0HliAc9vR3dmFVHvWjZ5szD1JmGZw14tgnG7V48GKbnZ
Lm0GW89QQmRJNEuEPZhDCyavHImvXx8J4zvz4ELr/AWzyv2oGnuwE1eQXl5Mq0520Fc9jTjyPYGF
txI7GL4GXtZW5M4H0+vhtN3QyaA1QPqrAUsLYZFR4vzEVztxvNV/9aX1UEklwuiPwXrsnRyaPkN3
U95XMxQjCRBiiUROGAFeFUsWO4G/KSZNTarc8YveRQrRAPIIWyCMEeduKFr7sKfSvxoIr+8G59ee
NRIBtoEfmxRI11xBOvqQJ+KOtFzwWnqRCCdrb4AQ0L9aMuGhyHucJ6JI4PzI+voYHMyiWnyr70Ua
fPhv86ReidimDxt9zbz8CCKERFbTaSJTyV56YIPMs0I1B9QtSfoe5Orp6SdErBpg0bMEmG13J946
LhnQ4fkNfqNMHIGeu1bRXh6CxsohGnuFQpJxjpRyYqU66zzns+tJ7E0B/s8LtRGMaAADmg3GfoNu
adf/ebou8+a97HWr1/8noZCXhiwXV7qyqqVsPUuc9VoiXmkkfBsvwPctcKODWrDpyDd3+in3Y+0N
U//xzV1/KSNdFahBkbyHvGvP6apKtJnLHkkHIX6yKo7HgfVaVZVaJLSrTd6FyTTpMKUt4Ff1mYuU
htqy+dzCO3eUjKcnIzk7FcbN+91DSp3kMVE5JFzr66tfsrRDndyTGlM1GRXotsumQOZPMYryRzTA
v1aS7QF/f+NB3TyUZQi83uTRvA3vOIHlDzl6JHneqVR71PmoHJArQk8hw1xVa+Wfelv2dcV4e8pu
3iwJgTxucryTxcAXNeSrOB3rXQuoghNFeRLwhzCZB93yXk2jawB4RZNcImRqaGLFj9poMFR/RkIM
T/4c0gNmmFA9vktDVfLE+VMb0N4gnEagWrHb1hvy1cDVWs+piqUnHrvxtKxPwo3JeHTtW6MZNlfB
RzukwNcFswsXVWGtn1mTdMH67uweJtXN6XhU8KIReUiCVvjFqhg9c/z4zlGa/ojxR42I0vAM+zRN
vRKysXoGUma3+pIT5d2JuC9YWe26EK+T1Gr7dh5mOamY5Y48jlg23QRqLqeGWRApPEmG78c8WOM+
K3Zqyr2yz0xP7yuxIivXEBWtYDmE81GIjY9FTqRB4SAEpbm2Plh3QwBsxyD80Mh+jApCJFL3Gj5T
bDRjim4IDtGLbkheCiUzM6UywQp6egUa2y1QlTxeIgPBYNYoxO6WF7R0tOMqeulV3Ln/AIdv4DgH
t/fOyNJcexM4tRRCjpqnd8OXWhpzRqdj1dA954peqa2iWuor4vXyMBmARVgt4B4BSqK6i4r86IHx
zdcodxJ1iAmbgv2luqqoIlrYnqLeLbDp9h3w/1VbnfhrOBnnC870BZMrSQs2V1DxdQv+m7PecijN
DP9YC+aWaJmPmXkaEv3f9DeRFIY/76iTHjCr0erA/O0vXwAUcvT0UZlBnTKAEfNsIJLCG972idhS
IfWQDtaoOjNT5AlAFr805QPVna2CrQJ7/PWjORlApDV5SIV/3VdrIef3o0Km8K/CsmmqJ23ILd1u
/4QOCP9D0TxiRK5xoGNeu8V0UB4V9czN2Szhjza+P8cRKCgABo+zOnTqoT2b9+hwllNaPmnaovKy
7ILwOGYPip5GvbMInUeuyH/n5ZNC8876LADsMRBGqSYFeBMMJaTzRs0XHKON0NNIgty5aQ0u9cCm
tvSwlYEDGjLNGDKE0mk37B4mcR7POjaBzGwybwlmmBBsyPcsNerbnlEe9F8wKw0KUhzBSI48x32J
+LQGzqmSvdnNQJ1WTiT8nEYmVkf8PFTl8z0p5NczO3d6CVu326SUsC7dtw2ELPaMXzyZvhAMaaIs
VkdZKxRqVcfkbHsEjL72uQfU0zlvhLxDEOjf4tbNmSKXmQ162gCT/fr9WZJIgXSg/XENcrzjkzz9
vCapEllN0nKU1kvBnK1ODsN1hCibvr/2YTx4+YJDxSFjo8hgIFjuYlTDb7FwdZJWV8kmnMsHdQs+
0aqscLJJwcUKd4o7Wl1o+sUIwOSWqW0rEbebPvL9roSu/66MtKXao1imqVJgSN+WvSnH66gxlxOs
JEgCiWEXY7xQxrpqNw6uuSGv3emhuhQYNYE2G+VzrI+5tvzbkWZz05MqY13mLTnAr9x0zBXazroQ
bQ1Dpdcao4bifEHIVHWBXBy4W0dq7zx/jasP/6/MsKeLLSEMTnLLC6Ppi/7CPmzNj7ABSYbEg3de
0LG8KkLDEoy79oUMvVqtmh+CXDTa8dTaB+eff9Qx1nzQA4kWnjwH93NzIlPUO0nuL7ThqR05EECG
1reMqyLrgrubmC0qM7QICmBAVdrb9OVpRp+YeCfkk2tIiaqFUTg9G0YUs41MS9GR1ADD3cs4MwDz
51+Fp1Eg3I8h6IhzSLj4H9iE2kYdp/b64/oLsYN411TQjtigkAqZfTSP5OQii5nuQqMmc4mnWPxH
Jlv11/Hemdx8a+vaP7aA8+2p28kJysOcFatr3AKzCSTmm2RLR02HAwKxPhfoyw508tNNFZYbuRR4
NKs+BxvnfxvHjRiKgK9mbL1FVowU0k68LP696Gm33QWcqCfB98tC56o6A/3DMZ3306K56SqMyFNE
ViHWr4jZdZ75OImjxalafwD/nnDWZGY6iDRBgh9rDJQdpw/zHEcjNok+eWi6Pb6qzug3oSAQ5Rlo
2Af6gqp6V6fHNfMLgP7qdqXrSwnDZfY7Kfp2vMFGLVFfjvb7Ir38vZIBluJDd6c1fQ+RWPY/sVlD
+wKK1f431kN24b5gMHAkLtceFXMX8DnEDKxWO9sU/2sdYjHsOH/pk14t2fEHOVs1qKDQqrJgT+GF
fwxSObP7HnimjI7bsMGvV6w8QdFIXstqdWglfWgd+BiSk4GhK6nCcDcI5RiVNHeAjLkBdokzy8OZ
7758n1QyaLQvbISv0yo1HMv8jc45+nX7JGJ9CQ071wauy1yJyjxU9qYCkzoOKZgTyabX4/LkWf0Q
40PwOZiwxZqN90GXzOw0jp+gAsrRt6g4xzvgdOI7dnMXUwkEvDKWQBqc2D125aDoVB3xzfkG3Epn
FvYX3ru0GCgaXx2k2/R+GVZBuBUQ6v7R6gmzSxZerz2m5ARHV9tz93VxegPP5pYMV3LlrHqEoQBx
cHX/Thnw1i9C7HcF7J5YhHP1YRm5YU7BAphejyK+dnfRFOMS0jN4zNLCOrMEMaW2Ypnzx1TLhXuw
sg9TKf7OhnD0IOWB7jwIDnOCT0rQpd5bkRkrWz80jPx4/j+oiW1N1XWbusUxnRaE08zN7HyFqBIQ
6xDgJoE4mBeB3+LYeuhV9c1G0Go8++AeTwA3i4muwwszHUCa6B8m+SzYYNxvyOFaOnBkNlu81cDh
2hs6rJzFg3Bq4RQunGEASK51BGTn/kVP/udDvhMuDj1uDIqALv9wV28B0+chwskEqDHJftt9d5Z/
mi5NDLM7qeGsiJE5SAWKup+4R8h6iYbXLgu/++j7t6TopHabV/wI5S6Ceba07CAARGs99z2SdwAc
EkDXwyUoBGOr2vOukEMxxzomxpv0DqtOBFDZi5MksDak8DNi6oPDvci+xwXr5PKmXV2bUAznjL0d
BOt2o62rvHfce9bWsBmmFoIKWO35q67enl/CI7xJKZTr4P69mjCGBRFoSn/TEiKEQauPMwPI5+o7
DPGsO7Odp9KCCg3Im7ZO6YW5EqAlMMiMSqDLinnTsk34p/6KdMKtOdy5fzR515NmwvHETX0ySoLJ
gZIRrjSHxOTNaLSi0vqjUkw+LOJS5+EpwTRsFrESNmNl8VWhYCcbYLRRMDk9dqfP+fWFgjmXb4RK
7k9amc2V7TI5/JtTkX1Rrs8t8TM2NoDncOAkAbGcktXjAcskGeJZePPO6QII6r362OywJfQ88QRP
YtO1t4/BOEhRlVFWNpKUpQ06A37dfDE76vQ5XI1EL2c0lBj//plZoxaY+ruQAcBFhx46qG7cbUAx
32OIzlK5CWxcXTmske9DC5boTNRxrKOxSxFsLG+0XnqFEYws8wSGRnttA+4ZbNCgfl4gF6h25xTW
amxSa6VnhqTipmld2cWcu1kLCCiZ11Oa5XLtpNgLbTDFu66PcvvjBV47Deel5HNkuljdtnKD4bP9
NXVx52FIIdu2+waKdayp0RIIySHvoUE9UjSg1rsDDRRbxFOCh52f3N6sxUf2jRXTzVTPLQxwLVD4
SOCauYF0Xw0Ut21xlQoFyoOiCqg5cRJP+pfav9Vg3oH2af4Wzjcl3q2qa3u32hvcFPhbToMbd+Dy
XR4AS3ZavgvxA6bova9taXqMixCWVDipqq2DWZRyVK09oEo8Xs1oQRcD4i4yGAmZi/93BobJeY26
Bpx2jj8FyFKp2DZG3RcWC2dPfAS3Pp+2CNgTF2pdU6N+iEPmj27/QxtjIA/KxPm9z5dB52QHsJjH
mOOVo0pwslJz9ff6tgoBrjJs/lx2tnQLrBd4BGVeXZE0vB3xV0emmG4YwnV6qR2vz+ImIiBtsxF3
YOZhWDvASriRaLOTOZjKvGOCZX6buQEQ7VN7FMYU/MdWE74s4lQN8/V07XLExAFWIM9o3T2dMjws
FYEa3zjikh8nCWSvA5HK+rE6qOydLYidv+89VQ3y6DfpIidjTmwGeB6vVQ0jnEdhDYnS/iU8xJUz
0C/QsEpdXKuivW7jX9RUpFo/350W/ZuqTSIPxIg3y5w9dVn3pyea31P9l642JISBbpWWCxGYwEY6
8AZgLhL5TcBDjY5cq/gCQguJvHeoMW8xwgvLo08ly52o8uBmxawNaAQQ6xt8dqmJq/rad4zMr26/
msW8eHqBjz0b7hdfO/s3EOITJ4O7NjwgbMDHnILxtzAjVJFwaMSOVGkzBTK5Ph2RZ4+yKnAPcLFD
R7OfHOZ3gwMVyrzEfYmXn0n+3X58oF1YmkD6Tc3B/xbYSY6/1zBBfu8ZgZiWhV0CmtZDtTFbOVx7
l/IhtXZxvAvidIHCRZzCQekGgnUx2iUDMYO5PmZzSZiy0zb4EzmklcMpFQwmQZb0CJKjg24YmDc0
T1BQCC+0Ux/4pijPe40jB05B/4HGi6ujquDx2Dorxdj128yCt15+8/VkHY7WvferbleoHiRww8or
ZYMGde+RLjiLWc+viwJ/lv7xBUaAtvZ57sjoK/vxidDZyeOetTvqxR45lt0nmBxWTGwDayc/CbvY
cZ8B+O24e86gBmDrDLpdV9ds+6RXfPQCAWvMROOyRmDiQDZ2oO2GHqDEioZYj00BQOXdf0Hwp5Vk
mJ7+xQ0FM/mMWNBacAtxm/S3SpEaCKw3EZWF57fqljWFsxrT4t/1HqwT3co86KrHT7+y4q3jmB8W
RdD8ZhewIppwXijAW/ZxMVGyMAJGMYwDsulfRaZZEjqlNycXJoVRPFKxw0j1bX+0Y6yf/bW7uzsD
8LbTgIz+NohzREc514Ku
`pragma protect end_protected
