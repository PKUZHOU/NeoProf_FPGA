// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
R9orTAAjMgBm7cTrDZCh3T5olWAra/kn2uB8tcKx1YZYyqmnugwqV/xUlznVOAvGFRKMkRmStXfw
HdvHkndhXFcMIzVBcllol+v+uscDaPasfi3IleOHwHhWWiBBzJLyFH1Bf1dgHmylU9bfS7PUF4sQ
whkin04xPhRIWzFvSVfep/4XgmZTIJ5imtcmu9J0iklwVDRuYACI10fANZqiGad7mjXnv11aqeu0
v70EyoqSSX/QjN6SP2Q5TkPVMzlZwrrNDUPBCG7CWJTJZZCwJ8eJyBdP4UoNUZTqTqxyDZR4lM5H
w7oyZPpax1GIqrB5gpSSbkCRJ21gJbTvgGJa+Q==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 81456)
iYjDGVeP12qhrfUEqaBbxBbPVFiChnNndE9COCOp2Dnx3You0Hfid88RkGAzYjaUPVASuatAWVck
vyRrgPWhfTg9lGPL4pCm9VBEhI0AtooBZ0pUy9PQElkApUYTg2EcjNoKVbUek2q4o92D016F9hph
QZBnQn0IJv2m7pXr5OkIVaLzeJHhd1uJeBDCeBVGdTVff9PnxoN9O9hPLJcHR8RyiCrJJo+cBZ77
tUKJtJ/OVa84zD8atrgRluyHmwTcFkCIfHULUCpnj31e2by6a421a67BADGVewhZit7rQSLkByn0
2ztLYNgNYE0oNelv/ACWuUfhmByyi2dZ/HhgLneUrG1M1jhGAmGY7OaDXsEH5to0eSqp5EqJUon2
wj25XdPUEi+fMjs5yNrIhNkbP7gcIV+af6P6yZqg1qZ8tGho/jAfxlEV09+CVGUKAdeuTEdiNYf7
RRl3xXeK++blhHHZ3W5+wg0irdUXZLLV7TofchoqZlJU6z5bXeK4YiFMBejC0+lB28u8lC0kjhkb
fZLwh1vV9gGAKfdo2gtNO7q77aBDT+OOxgc5pqzNWLsWFB5FoOI9+GpEK+0QLPi2ofl6StrRmPCC
bORmXM1Co/RalzsQR8EGHnLGzRRj54wHFHDixLQCi1TOYBdCD3BPNWqsdUXF9YR/CqFQYvsj7k0s
JWB8vetoHj6FTFmSGBfByDj6yzvvdfsbWfFoO1C+Sn2D09ZAubk1SaIEgR4JKTfXfCG4cxWLOTgo
bvvjKQfJsqLJtD8rhXVBTwbmnMZdH0Ujkx+dRKSovG72QKH7SSAQA6g5Y5zIT6mpVSFSUvdcE0hF
pJxQLHo22l328AOomaGjNU/Kuwx7FL+Qbxij/ptjvHIJMF3/CuAPx9W/Hgk+KxffhSaTn0Tb0BeW
6sT0/WxTAXGsMaVE1QAYOtaIWB/9yNtTMx8pflP9Q1R0XTdsqSbFLzpXOZx1Qvg567uD9/wBpisn
QYMlSBdrEQy/qpcA1MviSU/USE95UYEpDwxmzboKE0l4rz1nJyHw4S9LQWdjMVQvAkF9h0+W8Xlo
ii03diH1tLZVE6CfJ+rku1BPZAEL6TenDj5ltVOTnN6P6uT5ItXDRu/1pRM3FMAaiEaBw4pegXz2
Ide2tPiLnS6pNNh5FYwA3uhYbAGVAwJ4A/jAvLNiRxplhHGe00n66o7eseJksa2tu2TeqzZEphNy
gWGUuUPgrxyOSA8yJhpLy55AIwpPY6DYzq6x18XQQZ/v7yyqnVYkUMZqoEXJ+ZMdTlFWgnyDpSLb
gbtN6AuAMOGTk9xVReK12wEypFDb3/4QI+Oe3Ds1y5BET3sclfLHOmgsXbXmNyJHpRWjfzPI+7K9
AHqw4MNV3F5vsC9aCycywrMZQWMbRbUbOghtgduxXJNoneOUp79rOkDRzUNOqjumA7tA5C2hpEgR
rGtfUqKvt8wDxDoo88kqFqdXDpJInTCOQ9tRi/ZEKaH6GfqR/dsj1gaoGsWIHb/gV4ZVBb5Q6RGx
Cb1ot5AgVUKNw24P5YpnZ8lz438+mRstFzhXrggEU9TS2b7zffzp0CmKAZdd1MrIYdwUTNXJ44Gc
2EnS+mTaHwbiIMYsMuhbOWRQwLhLk635muDm2mYk784lCBb9NM2agy+afDk+EalGi+eDs3YJlU89
mqOmuW2GuXBNwt7s2bEL1WICGBIBx7udtmVdyLQU+b4LRVGiaBKBbFhWkG3x+1fTdUX12m4t2oAd
WAI0PKLuJZOoe7rbTkSCNErpRPn35gRmxAndF4pYs2SrJhzjmg+7OTXbzXiARZkLu4QX8v8aFygl
PHNBQ2EIoO2I8OadV4CVCiwW8hnJxyb/+92Gi63J8lv3PcpMDlXwGYjtFZq6dQNhkQRo+XL59XDh
my8uf+y5GPsJ5oDjUUIQGUQiVLNAB57AVLcGbdDQZk+C1+A41pjPynJUj2c7mMl0b2t0TwrEQKEj
Wqm/S9SGgEB9xynu275W6Sci2AfnI5a/Wxto4Mfggr8Fnr0VDmXoir0tRhhz9SlMzQwLwkxVTRwL
ztH/6NAoATVtjsRMnrIOTp7FsHq9WMuY59Yx2oGEKs8W8Ij6J+ru0+0cJiWE6utf/6fllD42RSZR
pIvBot/00HHwP8qqcAIW1UKoSYuSsYMB1lINqCKHVV/+pJWNNSN3Z8kxiiuXVT+1TqVfPk4RtTK0
yZBYtpfjSVFLPsAsRYS2rvpehNlemMe/j7T6zozrrXyMF2ZocyaDg++fqetKTXDwgkBummcOip/M
tncQ62dH4ynqgjvffuQXLwmBiQWmge2bWytwsCGmr6s64GtHV4QUYs4sJeI1OtmrWbwhMI++2hPK
uDLZwSph4isOms845kRqkEbu7W4b6gQ1tmYQyMusXcbXBHQgdu1MEFPqytCVR4qjamZCpN9NVwuA
B5/ix/73BlNCbAWMCM3Vqushyn8hpiCMGiA0oDTDXohgaKfY/nKEc+lm3+7zPo8UisNyv6bdWJUr
HQ+iA4ChUon522pShDNPaGcu81t/E1qyj7In9ZwOaH8HNdcTM5P8QxRICj55/VJ82IIj4e2MDgtP
ekow7rodzvzKjxkm1H4CwnHHbfwsCxgO0O0Pzx3mCxqB0z+2kX4Jy1b5CgBHQ7oaNtlf9bE37F3T
nw1Om2rl76CunqrQIt7S6nIrs86Xr6xbwtdXQsvm+3PgaV0/QYvAqXKfkvHEOmAaUfvkfH8Q02ZL
+Vudw9lZGNFmSKu2WoFU5FXssFo8vLedz6Y+9Fr2jSUVPJ1HhKPyczq1YJs7zdzzbhaDSwxzuNHO
azN+kFU3ouBu26ui7fYgPoZzXXEKEy4VqYlCv6ddxSyik/NlAcJmZ1pvfrU6ZgPNTUG604rcbXYF
T1m/kP+eOZwCKDgGRSp40N8uG/BkWioCvTajiBK8kNC1Zrk+F5ZOq46E8AwpTbd6yFF+Hgn5/zlO
j3IqmQ+DtBwUkXUm2eCxmtZH3x2AAeJaLCaiN1s+CUqCI82gghvEIl6TQrrYz+4ZVDhnjIDaubOQ
K2vr7S31bbfSRYhvZPs1dIBuGJ5EUIz+J5YnbwVCCYHXkIANwpSObgbwsckdL54eujeeTEOry6Vb
m8p8Qit9wJ1NbsT8UnTlM3rtjQD7lSPJBYDqBdT+6LhtdhP+qjbaXBBQV82jPiVCEBBguhApq1kU
zwXzI36IpoJibKo1BZRN/C043xWTITOoyzqWEiVp5kqNX5EPsqW62VGtxjCXb3yCp3QI3hEK1BJR
0nOj6U3yKPGgMSwl82FVtvCCfn/cNxbjfBx4DI1EmplIevfi+yWaLH7QigTrHSnVv8hmBjvGX2Ic
xWQA8MblrF8UUFxcKNb0JU1nwpsDyEao2RX56F9iAcHYkxRUkS3cVTHtOnjN7rFqiBXtM9pv8rym
7dv8wAgYi9/IFTHBTb3i8Vwg53ShHgHCqlb30IyhSKOZR7ia4bWbcxuNeuqXJXLw5KnOctQLgG6u
abZzHLF1iBfcGbPAyZZVn9IgPwdWKplyV4dnEM3YkvSwjdOjLIhL6hUQgnKzUGhfjog1qKfv70Lg
vyl0MJvMoekc/dyA+eZ1zQxNALfRRPiA9kbvB3DlmA8NfYnAUFrg3tz3RDNhec815VncOFPQ/U00
olyTbnaOiSeu2CadoLuSd8OBJ76TmCBrPjOGLJvWEOfurJdU00qoTTfVsZm9LWvSVSSND4Yu9BBa
uKYaFOH3KYdWaydb2FIAW/Ib2G5MtUp3yjydV4g4FB8SRMrX5K9WEKyRGfWJdM6AfdV4wsucuEzw
gKqk8GqwTvt443lqHSqPtLwaq3vfLdzVJdYUZaIOAm0UgHviZQqdnF3lNSz81HDhQ/EwMkc4pP4O
BLgmkoKZYV09qmezlG/MIAL/oASrsB3lt9qwAu1p3pQonyqDWS+tTDykDNgbEDiAC5yzF14tbECg
YusYyi9LXOtdzcm1pnXBo4rgYtjTSmanbi8C9HRu4O1iDFB3H1voZdoHMNTcq+dNCaUd1mi9zHD8
8/wg82kCq+IgxcV4RV7b+uu9gchl2rmFbd6So/4G72EEG622dctlidV85raHW6LiL/0vyZkI9yhO
6atWbcy+sJkgs2BcWlzWEHOJBNMHVcjUj7of9yLm08G61T1G4i/MEU5R0CI+MGYHgDqnIi3V0rVY
R54wfTZbPfFcE6ufkJior+BXKfMxe4FnoJh2zD4UdDmUZZEXMzbudlJtgED9xeIJ+LDXh/JTevon
xw5ZACBhFTaApU1etuUtc+pnZUZ9Skak0/QkUhud/0tXWlZ89K3mXDxEmAAUX1x3+mKK7eYI97pE
K7reKsSnsj2MsVIqaICKLrld/niuVMWdTipkc0eJKSBnV3EiRtdfIl15yjD27rbZzNMSHZ+M3e2Q
FEVn91M+YdcgsT9TcN/zwpUJ2x866oes3iqDlz4Uq5C+eLS6u/95R0YugJJgaAX3W0TmlJ1tOta9
NT1VXvNbshQcx8rb94prtAmzSgP/0KULhvC3No3D+8zyzDLE7RR+ohtFgTuIRq0ye/2HmIle9Aj0
KGUYNKi6RoUQn0dYkR9XAveYpJVFY1VDmEVzCF3lohD8ncGq983wlYnO2c5SneHf57X9z18quPSy
THQhGWTRUQjWKXZL2XG9eviij9CqhTyIMCsIKuyir1T47GJ9mi761kbAGWcjscleDzqxEGP8+DFV
357khZ6XjdxjcIabx/gnqI+1CiRFS+laXruh+GZUYqb4XA0RII4Ki6V/u8PqO14+OoOCOBrcBar+
LxzNbKHSov2N5Fm+3bNSo0glRVxAYt2liL5NDH0LqK3fy3+UBn/RUgQgq4MilvhOK8zmvDkXM/ZZ
IElG8j3x842G1X5MGmqjahnSyRBYpnzONqqW8Q47VyRgmrbkyp8lvjdFUiGpl1W1UaZi9/9btLrI
AgzXHlvCRUT+jwyJFVclAQh62fMwxI+N5636YbtL+TEpg+t3KJd3CVL4Aeiicv84uEK9S5mAM5Ow
6RFTm7KmqmLS5EvUcCFao1GRvDyMFHxadphSbCBWap8JG2T3e7xlzY/Jmwxc7oWgDcBvH1uCDDJD
wGUnPl5KMjWjF2ldSHQJ/QvebVqHHzYOOZIitiuY78d4m30rS7rXFFm2zYumeb+zWzR8EHfiuf5J
NjJ6p4hQttCdFiwd2vEYuhTweFvCwSUuQwGLakFyW+1UUXT9QXndtaHM1Bx6ItBhiAqpyZ07H1S8
Y7VsQJLmfMcjaZWsXNjCBM4Fwjy3+R/vPG2YpmS1lKl2Hb4EvSAYS35ngcz+wvWIqiiiB26If9AN
H3iYc2m2Tl9xt1/SIibsirS/piaHbNYJwHzBUfI6LpvfuinJiI2H9iJAOa43O6K4UdaYVrl3qmZG
RMDo7i7bBu7Lhq0v6JpBbWyXz3G9cFw1238gEntzRsG4sc0zVFYgGuQ+Hs55J+rAWD4if57kMq6g
Na8FRWkaJWg+dI0E8NTIqistkkY9DtbP+FIPCjoXivUW74WRutMO7+BI24LHSf3qqc7GaERtlNbW
pi/0OuDb2MWNiQGSfu7s+H72raxvGUW1KeluaFCZR3XXWUv88PbHnQEYLQVVhu9FPfrJEz65wHeA
86DXVV2kx59NraSkKK9saDA7wamw9zkQdCWRGKb2h7T2EWNiPOIPeW6G2D8Z0z9LAAmUw6sAHIX0
oPFjFXH1W2l5VCehJud2zIRIaN5lIRYVKiBCznycvVBBUMBkoikywuzZAAKwmSgnPEZ2dgioQi3P
9Y5HsMF5qs/7GGRC2Bdp5cejY8D7aM1XZua+1kBKquOOLHXQpVo8KQqotggTplf1iBYllZohK00J
HJNHT7IuglbKZDXoKqGbMVHsjEhXT1n9A+4ZwT75ki1UmlpfzXmaNHPpkwCpTk/UTRJsSu8Y56pU
OqaAiTUNQdcYlVTnfwWnZY3IsL/eczMIP2BCLzgccI2rstIkJLEvWTaxPKffeYMDTPLSQo0QxJOY
JZmxB1N/xqIAbm7FcInjAD/KqYAYwSEF2GTPqk2KkqVQF20OfXuV/uMXuxyNZjwBFM+jPXEIMmj2
hWjieKlt9A3zrQun5m+8BfNyuXDGfC12dWIpTaJmqF/tqYaW0XUvbirTZhLjbmr9WOiWOUmYf8Eo
oPAlKRmzNDjz7PAaltW40K+BMYlGdV2GH/uiavYiGg3oZZDJIwVEpLWh9VL3ECkLZL0mH4o9xbmx
LNiUNeFHKvAXCP5KY7AYVCUXopZXv1HtvW0qw+CHnO1kWF6BTdiQgYw28IVCQbwJNX6MRv0ouYiI
2w4OrrAcPXTeDqlrIty+VnfmGm9660DbEfqrKpzyi98X71kdCzUqsXFdol3ChreMAja0cnAKpKtL
dToRFoX9nwsAG+d37ssjEiroI7zgrtIfdfz+whZUIPq7uGvaLSKK6fGxQ5t2Tyz8XdCQ+S5RuHm/
oqfGtYbxWPvtheGAK9ozBeoLRbE/o2lf6mIboYJSS34MaCrAyfpcQ/9b90oaJSdMrdQSz4n7Hku+
OGFmetyuGrbYyXQd116WyMuJ+g4vVwodjmNUwEgOJk8I8ARgib3t938wEovtwvRKZxTtJgSh4A6O
cVef+LxMsGzqUFadZSek5m+D/SKNYzqCVyAILsJXgYAH+AGU9ESgPKq72Af83pAao6gi7iyBSBdP
u6GZIEeEUIvX8Rf0T8+77rz1A16iRVoXR2b+r+eXAohSg/vRpbt/aZiUgy8o7bFzwzPatvuYygYY
ViT6nPH5zPCSV9OvKr2RjW9LVfVGZJZVuU2/joc4TEENGyOi4PeW0sd85UutGkH3CpsVoz832AYz
3BxS3nu99TEWL7o7K9TM/TvNsC5h8DLt6xSBVxXNVpH5IHJRF8ffso2nAnBLTeDsAY97N/VIvVVT
KpATZrPK9bY1MOPNYXk7+15HcMXa5f7yY1l+co4i4At6vQoDL7HFX7txAW/BKQK47dEZhLE5fVHj
ZAkApA89TG4R3w/pr9UjkHs+OkkmJAzv7i8PkLk2LPfqMdJ4yf1maGvHi5QJO2g4FEPLxRl/Z5Sh
nSDMDP3/5A6bTRvjrUdXC83iEprldwmKdbKVGd8f7m/xWufAwpaM+EAXpQUrmcQjWbyP8IgXSsVi
hcELdljaemW1oL9vi0vPwHP+kQ+/NPdNOs8XbZGpu6hfN9xzIfxlx5ATYiqeAtciJL+Nk7oCn9nH
G5GB62581V4Fe2C8irfWJZYWf8LB0m1QyfzYJEYIHT43eCh84UuX3aLldFCefqI8BEz417RD2zH/
dkhibcCrlUleLbtD5+nGW1Ehs4lkeRHM2upJtwW0cxBVd6Qc8VTOqUXNZOUftvIzACHmmjer80MY
a4YwUoHdWWawDAZdcNCOiqRLiEXfzk+kJg+LVhWCtaUUVDDa0z4Vm8G0Jj1MSmX1yhDYfCoi878A
wZ4lX9VQ0zoDmrqM1Da6NyXCUCPNeGoAG9mcx+q6HI1S4pC3qiy8fklThnr9wfzn0N/+WHMQHVdp
6QQXfaAWRZoJRa0XofqMUTDKECK3O05LnV6VCCsPQmnq/B1m3n7t6YZnxM1I3x7Smtk4LSaD7LrK
dzEFDipj4s2MNC6ssCPskG2x1JoNBYYqlM2e1/hVsjfRF/AUKSdOUYAU6EsGKKqI8ZT/2yw/jIDE
k+g/hWR8tkM0lZvSfksH52j1bsUi8QhTcnYSR9O2iYAKisOhq3ugSuK7UIqQ5AxvzSsf9Cq52XzC
F49gcG4hHXtK4AE8MB4bFv8g7K/YsInLR/yKYyn+OCbJeP8KLnEuqAKqUEQjlfhCLl0Ey5vS1kXH
XSKa7+aFdnYS14b4j858YocO4GT7zw5rB2N8ZJR1+7awSBgAN0QB77+E4QyQfPaehOPvgm04+/b5
ZMU4neXnt4JOsM5O5EfXV0RA+aiBBui18yYE0IFvz02vvFoFTTDdxTSzBM+D+581Or47zBfY4cpC
rt287katyrUmRYZNQ30S3FxU/5M13ztEvY9rxw8wikROv0sGbP5/Z+5Hb/f7/GxhDkZRl9t66h2o
Z481F3ZzdpdXuhnibPYQS5Ak8DCZbRm0XqVQ2Q+DZ4xGG8k1ow7oKBT6pc3QrP85Z+uES4fokDpf
57CPr5RrxubCbfALn1+Y7x5mWJXC26U42qisI0DnAwwYbmdkB44E2wdoM+yyRsW2JZ9xR33xTgBd
cnPTiPPnh5WiMPciESEWRPAQeFy7D862wuVLueURB/MXXPHeVs9hD6tDkOTxJLDC+UApGpA8TfvV
AZro67uOke+f2eLH3POyyvJX8K4uguJyNhJ4Pm0jEBuNC84TOa65Xmi9/Uap9e+Idx0mmFpUJdfp
9++Z1Dssfe02NR19XHZZ93yScnhELpy+eZvUO7l3W80EDnE3EolsftJ/CcCa5DaEcjAd60LAVp/U
ghaIIigvgAv4Yi+t5zxj1wp0GJena+z2jKqd71lTXkiHjt4KKuNxJbW/31PcNDUGaPBhKoEztJmX
DIiR2N4OxvaQBBcMJ2NSt4mLTqacroQgdnDkJ3KIjZ5V9DQX357PEOLct/S3/rl8dmaKWx695XnY
rhs1P5OrhqkuXocDtI+ZeabRPHcKVIKGx7USyL2pf5F8C5wQnYc6R4WFiCV42s8Wek4rsqVG9Ri7
oQznyDcRLbf/hAY1LIBxU4S8CGQ3UrmVFEk9WSpZltlC2tJ/mJdzdzYvLUheMVC6iumKqlukyHV+
a97h06++0AJ5VKYsIuSgVca6Sd+lALDSM074DnrY3BfRGc7N/nHP5hUiVbYsA/0Ekh1lK9KVbB4k
ZaXUZKcccdpft8nyS7xqzl3pV9+YmwsM0mETyJRfeU8ZJJAEGIEEttpBODFxg/HKzbbSCIPcgWn5
m49c7ZXLQB6u7MTnYWOOnvFQYudRBIWGsMZZrBBixPts54C0VzoMNhIv6HZAFKbHNws1N0+NKmhx
hC6AozNgbkMGgsMEaRlllRyIfq0mr5oU56KzjQtT6R7SgdGEjlAR0GPFUc+yaLJlgL+8QSTW38su
f80maCJRbniMYc4obwbhpr5wck10/9o1jr4MUrteey+7oqYX476qho9X9ee8P709qcEwPCa0UiK+
NOZ2aXsm8Ae53CYXaBjNPqTbIEDUu26ghYRtjRx3b45ICs/xarmdn/yFxngDfZYEnOOwUDq2zhg7
RjjjkVA6MhGqZAjyX64huY2dW6XFBSXwc4aBtLM5zhIVuh8eqvfRn4YtZUkNrnOaGFsKDbCPpU1l
EuekaJBOCJxXw53fo31pCv/ZvzlNx6M0Sd2slzKqhkZMkr22eScZsS/9URgVtltlSfleQ+h5q1Da
bKtvf4jePtBtItLbXfdeTdiwyX8I+Eq5EM9wzKw89aQwrarl+iaDJbDD0+r6iyegevlmeQheP4iU
179ujBuEtDhZ+CgYCIU58e4HC9cLtoOxjmUcPdIsAD6IrJF7x5tsGl+Ui/j6weey6MXnketTny48
tYvIRJeDLvhPQ/zHnqydmf7FvGRdP3nS4Zw6aDomT9w/ddKbj55RrV+/2XQHCgy4nMd1PYwXSWv2
i2apfGVw084XHZd2Icbcxb4AzEr6dSSRDROURASxfJE0hOMGBNevlZcnejVQbUCLi97OZ4ryvYha
0/3IJaHJnOR2jKQTx3MDvCHL/3ZHXw5kiEugLZRXjrX7/qLiCh9Q2mLCfRVmHtpgIS0F3AuVd5e/
qnE0EEN566i4EeVcd8iMWwLtuRho7+EtvTnX+fZO7YZw8NA3JvM2rYWbBW1SnICTStN6vZAMXuO/
qOC2M+rvQjXS0jikgG5dy7g5UliX9F4YncUdb32VpwKG/70u9+F00dSvw9OWJm+Ax3Z2E7LT7Y0Y
1Sqky+7Q5Yi1ytekm+iuPdc6XtPvp45JzKZm1jo0WNHwYkYJ7ma6xxWdjG9+k/s4uuIgwDKY7sk2
pmMWlkXS8++Ly/eHD599Xqm7Qay1hvXs/7AXNLriqzi7mKuF43puDFQAIsd4wCveT90KkvPxUxFr
nSwoH6q+7Klm76yLGCD12w9sGoWlCGbbqCqY0IhnWTJEgqIkpj2JogdBr5NFTsIGqXJo0DDeNa1V
fwBWOg3IZpiT2sacQBbIpfulv0PtDl373t12a0ovsyXsHRfri60brOVTivSXcRdnxUXb31dHCXI7
xxoQYYtpgx9yfquL/SNP9+ZXvG+fFYw7M6gXgVBKsVXTgF57MBYYHWixlVPkmss+Mo3aW96Y7oQw
TkVzQWNw15pOslO1uX/iw/FtMJfKLnShsMNYViFEBIRcs5wOuNyq7Z76UBx4y0suF94kgYfUHpoz
LxGHg0gsQgpuFXY7/B5Me2OYSmxvWz9MVO8cnDisrjV+Wo2LvspDQXiD/KYgsFHXCHJQk8IOkuoY
6vOuBXNYWNblQeiJHG1op4dHB5xYgeQe83mVmkX+y/9wZLuhC1k9ocwuwq0oMABppjfRmat3OGFr
/xL0GV+/RVEAw4Am3aiP04XvhqktIEjwaj6Q1fp1hbo8G6jwC6OG1J61F0fBEhFiWsx1S1AcVEdt
LSYOwUTqsGKSdEn2PE5iaOADQHi7yi2Yr1xtBxMKcjcBCJMYgM0BWZoDSCrFwmYH4C+vM5ojZar8
4kIrOvUyBD+8vVlta0TExgh8h7gNkECA0NOqS+Pv729F2oex+V25ysSLPWLtmjYNMcammnFIBOVe
MPPPflaX33/khRqNecE7aAEhXDaCB/t+Mj0tXxrKgB31D+DqDhXcJ+9o23VGaxGVFkGQnYbpOdGE
kPV+BnP9rzywfvq4xWnilremuFSa4Wp81rEuGgT/7XPr3jtmFxY30BXnyyLdihNi/j9lgnJMPLXU
tjkvODXVdIr4QqnBR6OFuTjCQhJC80Dv3LbK0Ad9yvjGfJ3I4uNQEnHhjrQi2L0mCZh1zCG8OLbW
fPziyVxScikBZ7NGcebLRFMDVyq7Ee1hgha5P3YhN22RKepLV61CaweEkk+wX8BpLefO190/2nTh
ovuhTksqGHkv7O+yRtFh26cEg+TtvWr5h1gRmN+u9P1FQvV2RMeHS783GWc0Xsd+XtGVR+z5VQWE
sjcmrHjavTDDiXit0l0rmbaKDStIL2hmI+LAuMOidaOhTh+8W2JXzV18Z1Z0kEkd7mH+odMsGgAI
TBS0TuEYbqSMVZmxCA9sPVOqQg19uhQvG+m15kqbBBi5zXMaY2gGNP38jjUrbBsg5cIMDvl/Aq0w
vJVTxjc1uUXHG16CQj2BSvtVik7hhZGNz2H714+qtBVGHNYprNlHbKGA1PFoAl1m6LdFq22oKl5N
ei5kVG63CpjieMBCoexfWfD7KEuyddoaRwmGJZ5RisKOpgc6yq4RDGmP+J1vl6RiRKyfPwFUAJDm
vVPsNRF2IqpbTlC8WI7Oiie6VO/7rvc1fdkP1BtjJfhJ3rX8AJkHE2NhONA9fiQWvltlQFsZoOMY
OG3OyYqWig0QiSBFRS8Ooz1sutQl0ZNbQcridGtA5mnQYhAsbGHonJApS5omeKU7fpfrQD67nl+7
DWu7dHE/83naCxS/Rp/dboME9eKezm4AEvN7RBlWGcRRkzp5PiiqhNx5DeZXreohbAB9tII0ya25
sX0E/5t8Q0QPgwR0ROCNKkSx8a+m7nsPKtHJAaZ/x5pfW0okyUAzI6T0RIU/7ClzB66XUNeArgHJ
AzGArRTnhWUiBFJuDoq9uT3pQOpT+tUFGgHYLE1N2Ac2l+o3wm7A+KiOoO5DKKc9SqDrG0t3vhho
RF+vIr6ZG65bZTD6e4nNRWR42ax7G0UwrfSPEY6++Gd3zwZF83MEHxdB3kfUG98sbU/r2t/uok10
zcgpjkF3alC1Tvqv/V/U34JrCo7E0dirS9Git11xsw/Tl7nazNlOHHV5G1OV9UtLf2REXNFtDhYL
p5WAKiGJr9vW6XmsrxCrZd8Ek9o8aNQ9k9PQYzE/McrexaQZaWbF22mGiDGNkbw4NOrXmrTeB3mU
bYD7c5SbgQKa3p3cfSVhxNyCpnj/cwz+j2kjExUsTYvHDuS0ZCm5EStaPC0zynWMvkunIdadxLNz
lia4AQ3L6Kbeh4Qz9r2Vcp7NeLo7E8M3zVk8VqFu16zv+y/hrGqX1UnUN1J2cvcnmZPDStI8iX9h
OE9pWLZz1yKM8vu5Lqv+PYd7t9Ge18GvwvZva8j4eMWTS4c1yLeD7BBNDf1oYnnoFNep4cFFqWJz
UHxTPzjCeKSKqsa9eW2k3YN84QsxroUUZKZ50fTEJcqRF/zXSzYCr9IL5c8RpbYeRnCsNxk1BowA
cPWmMt79b0lEIwqiVQxztxf7Nl9+VunWpCmpdPZO89IAjepyJ5aL53FWeeCs8nasr8DectORiPx7
2J/7er+FaGDX8IQN7FocQVjf5PI/C17G9oJyD7bseH1JM+TpE+VqEFdaH3ArI9Ae8h92GCyuaqzc
GStx3AlLpQs/KQchO0g5vs+K1MUx1WANSTlpTxQeKVeJHb2z6ux4nCcB+238Z0DksTrOSNr+EPA3
RLgDBO0JGSDngzhzeEvF0x6Y/z/365RnNjqQ9QZidSC6Gz9T8653wTbkSfpQufDFfYvWxmP5wKl2
x2jMhRM87ma6Hz/IjnPZxI1b3syXt1XcAvhiCNEV+jmIEO7yE8adZt/wepfx/QDFWG+0wbpCiKHM
SEqq8qSujondN3LthTm9YrD8MnetwHUPbi7glSSWKXtusYV1q3Ztz5Rqwwfhv7bsT0iv18SFig3K
er8KoVWiauQkte66OLAOnf4LPpTTWEK0FiM8EimYaQSvx1G/drEMmX3lUybBYV1KJXTrQBkmY03q
FlKj8eSrs1TCzdFLM2FW5+BmpDi21pAEem+owiaESqiTyHT1ccBrsfqOTx5tlxQYFX/tjzKbybah
KBrIyGRkjY3YGku8ZSbgCWCNitNZtz81XQFtcbXZY5UvpN6ugHPXqsBeMRiSsFbuc9xHGjposzyU
2DEgM6gEQwpQHD14yFQr8RO58dhzulAahVuOgTXbGQuibyd6UBNQhDZ5LtOPGYMTZNmHm0tpve/l
00q4xiCC3Rr7YH9tmI3B4bWFszWfeWY3Yzree+rdI9qhyo2FNLibgMjXkDgMB9+mm8ZqTxdSngZw
JwdpQAYoNpAhJ1X95O92RcPCoQDlCCNs5QlC8a5/xYZoECJDHHaC+hE0V1h7qC/waaxnK8s2cL9A
KunSTW434XDMOrUJzEHiaFZuxv/7Gwn7MjQ2qMG6uJI72E8dura1sYTf0GOrM9llSmqUuFfzgqsk
/ALfbbcFt8tzU/fCYnk8MGX1G/WDtm49STzVLPmI/xIJJgIze7+sxOqEBF1HGJZbo7slM0kH1mn7
3vD7O3PfsGmtQtVzpVK6IZsScnBjR55k6Rnyx1Ujq7o/7Bx62S9Mlh/3xGLrZnVUIXCfa8XonbMx
BfR8L4JkTWSVkmNfbDuhJOo2nsR5GjxGLpnPXaohm46sWqM1OPbduePikDVwPpeRUW7LmMC9lrLd
0Ve2GuHpln3AOQIykUsPouxWFEoPuYY/hBP3IqRZXiBbl4djA1gaekgJzOrQTr+Dn8tteVMkkyt2
wUZ7R73tNYpOy1iOkTDwMDN7qBBxwNakia/SWJLvns9KEqjRokWT3VePnHjI5S2Zp0aZxyXzJHo8
8Zl1jnRRI7+x/xQBI8ViwjJ4ufdfGUtiGQlKZOBAkefKk3QuS6XWnrXdffUBpaT1A5tdhKXT2fNf
+YtekWwdpxjn20KPc1YfgMlMScJHYcPZ9EGEeemotvU8d/G0z/HpePKTas/wi2jnBjzlIZ4/xhB8
n1agpPuQn0h/AjErjWXmNOfoXdZI88npiC4fmEf+6e6JBiABXsklFB0RIUuyFdd8Kyjhws9CRFRR
iX7H6VfdoxfSWwHyPj7u8/OpvxmJIJexy7cW+M/4xMlcVZ4iTx7Rm/W+QUaf0KBThgXgEOudnMhB
UBWlAdynQL8SXwWVXEj08Uil9l+UsVrK2xqRbAnm+CbD6k4XeB5CcOlrAX4GX8vwTIhBEhjkclM1
SSiz1cSnwYRRtwIe9//43Mss59bJ375RHuvbzDcHckRkbVlAr7AEJZOoGopVRCOs7+vAb3CW3lju
2KirCxk+vwGlxCxzDIaSWneqwDZ5lbUmC1vjBtU9bVRsya8HfENBaq4JHjI2FOxScJKJBYAIN9Dw
1raZZvYS7L69/7Ky45ajNkCtkzFLZLqvJMWmmIhpMBWfFyWaNdpejKnc4UT/o22FFm8JE4G6TJwe
z1k9I9JfFwrpWZ70vfq0z5TWaxqD1szxugsdxirTssoTljP2XHkxLy4QjSdXhEbK8t7sTOVXDIsj
0dWHEx2cJ5sr4Ndwrz8K24ObRK5hPEXNHpXTJlXB3Ckrui0+ArK9vCQMhheMwRhWifwYhRVWjhtM
L9xokFfnn4mTM8cUrGKIAOE/BKoYKPWpC1znNLcJg7NvZvu5L+UCGLpUISGZv+5uKjcDKquUiW17
9fRJL9rWa63DkEOqMfjlWNDN1BZ3t438iXmIKF/wVfFYlw5uO1NBsbwbptbtzgZBwi1/8a9MgavC
ngK2aWKojSLCdLLeL4z+puOg0SF2yqXfhLpx5g2f9Uc6VaiLKbi9ZmgjJTior+uuqUw9gXuIUnjF
2888U/E/tRiUPJcpqwk2eOOvl3Wr/bJUKPLdsHKff5XyiVFE2sMPZlgjUjXbleOjcHY/B8tgtzcK
TpciOpdtlMHnHgXRkZxh/frm30rjxaoKeIjEr9Iw0FNFEBwGpd9xZg/7ztsonVjLpzZXwaG9cKob
yYPXBG3PUAWJyUel7PJtFwx42Qqpv47MjcdTh7WVAT2z2FfYFKfvHsgzLraDVuto6Ho/tBIEvURT
i7j+g+SRJZpjLlA4wfaRHoQ9x1smLiPbdXEWPmhbtTlr4Skn/V4QweQ1FXs4QxIrMeBBSyqr13Ja
m248GlX7u3mPrMKI0J4VoYJYvv/On4GJvcHP8L0bh6MPQ2NBsNQc4zjyJuQmn014r5aY/vCWu+kf
Y2cBSy7utPodDvv+UbBSs7not9w+Me4PAc0YcyHzoWbMexfe28seZN5GfbugVpkd+Kp+vR4G8aAT
zGHCMfoQuC+sAj6A0ioUHgzj8YlHPkPrFLABAtBqSNVD5TjqqXpuatrlLt6LABkozQidtj7jr1Bn
jSoeN+WPp8onw/+n6bL/lJRN/9m/R5IOTKTAcQtdK4NIGDKl21iJWfa98wigsNY5rdwNdSoNZs5L
wPzHRsESJWkRN80DXBvwSEKEcmSTqJCeJ65VoAOjzDhgcHIonbQE8KnfULvd3Pug2AdwOKtF6jT7
Lc5AXmbm0b3/LQLGmrfl+jSmSbMX6X9tp9RR9YkpmSikfDD14QUcdhjTTIP7DhTCbR4TMc03EFOx
22vlMnHooC7WK8ysUiNXj5VSn5DkQLBhnCIS9aoynsqH/rvW6tt8mpzXA3T8intGxMKkeNgrrxxm
v8yCXUnt9b+Gl2vf0QJ8aUiWHfWenEeMSPVBbfnu0XElN/gjZHB+bs9H4E+0XAu+Mpfw8nGuAttN
iPvjp5BtvwNc7o1VJw7yoSP4/LK4o9k5ymNGn4lqP5YEp6aHV+5yLeV4SPGdnan5IZerA4hUy5vC
Suz69wGuPh/b28XbtliJ4+tk5uOyJxash9CjdvJjeN93GtOO5HpLfCYFNyFaKD1zbOAfLgve52sH
DBzTT/M+dh273j1fOsE0mBYFBxTiYQyBn4LiAR2rjFNp0AthqHoHdpRj87PEnKPWBuaylYOblzV+
13IhQLwNtXDa93i3RqlaakGnf1cROZz0RtNjoY/+CMDvAjA0og9JBuwsY6EGRKqOmnM4zAZPhXAk
m167tm22YIq6OFd34e+lkIrqdfCVi6aVqpAnt9Brhng/zT/1Fyg40Clx/+ccQKktNlI1Oa5pH50b
/B3x3y2wa8W2C4HS+Wf3PSBBC4jhxlnSChN1oD9VT5/hXskRVSCgFD7t0b9+QbjuhaZI8N83U9dN
3spCnoCyy9d8fIgUBNGdnGbiwc5jkxMWDiCtr96O7x9zaESgqNkrvCRdb0Bc6Eq1VwYdk8mJpbZr
HB2+hs5SA6gY8WdMfAYxBAUpbtzELpEDoa+M9Wtk6wlPd1ryb9z5GhfT5If/0Z7pxDDVwQ2Si6M5
D6nxV1tk+3wjpFZbdEilJWiMKeInoO2VNPx9+DW9NUI+V6H8KfBy6m3yekODWY7Ph/03u290wpk2
/U2xeEJVhJuAF/VGAQ++Pjm4ydG9L+SNDRZ9QYhaOWIkIvTgUymZ+9xfdrsEtuYHG1c9jHH0Tysq
LfFjQqumAxABreqyAkHvfZpsOPHnvQf5XcehkKIv4VuvKp4xM7QewdzqlOyVHYcFheItbZN6ezzv
ubEahh+GXQas4bYJUQghQ4hKvopqsvnYRg1Tq+XLkgEi5f1xjCAMDWilIFBQxVMT67q0lfDS8jEw
KLjly6ZIzwpfpaL2Kuk2pg9OCcRRYd0+kBXsil+s/4VzqgVzVl6aCJ7joIYMqffdCtAM2mUufLxz
l4+UT0zpyb/D96UdaAvbEFVlVi5hCRuZZZJxGSlOfnwi0kqjy/DJMCVyjWhuoABa0E/o1S9jvdzJ
rA4g8a+etMnSCJHEn4yi1AF85pWUl/2VpIFUt7JhNPbiDMvnrbqUfBCNUc/HOy5SqEZIe37HuVPL
60jROes25/99IYPiArIMhBaOZrKysFXhPiNh5SrnH/nx5+qrITrOeNL85vX1DesXA7EI+ICVkmzV
O3RR+AWWFMKDUY5qQgYfBIN7nMdZ0fEHsy3CYuEIt3mLs2kkC3Z0b2Z8B5XDuQB9iGjSpGua9q6V
Ba/78Gyl9WCnnpw6FKC7PVGhQ8rB303wEyr/IcYbAvyU5q06tD6fGdkuQubR1H+Myl0ckHvvDuS5
RHhNgA8rcz8QVXYf1Uyp4QWXyULBO9gFEBYXJq8iY0XCsSLKv7Pxifh5Prq+9/cOupN3ydghb4e2
T6ltSK1/8tjFUn1r+cgVti22qfYhMyKok8ZM0NCqWZvmFySYTOMxE/fAaulODlblKiJXhSe745f4
entA4S0k2TL0UibskB5i5w9WJkBBBVBXPb86xcrD+G5CbQBkUvMv1+dc39nSqtHgkEv7zvAk/CIv
dX5b1libtBD9gyzVrCOH436zPMAYWAMcVqqz/TCt5DOmHHTkhWSiLtkl9I9wUAZxkSKfrqe2LCHD
KZjZyxjVYNIZTZ3eLU6Z58DUv3u7oU0WtzMpUm4Bahtd0vUPQUwwG3R839Y2VAUKS4v8eMmUsXlj
yVr9xy5cdWKknetaD0FeN/TJ9jmWS1IwkFfNvzqT5M5H7uSxVYG5Vxg2Wjkkl/vJdLcWO72JGNxS
iJb0D/wkLRKrxUibPou8+T87aTa6jYOWWrj/o9aMHGSY/glLQ7RfCZhQGyIu6eTuDY7gdDh3oxq3
7HYL1zO7D4a/tQfzHkNGQos1G7hyYAfoBG17mM5ml5XFX6TypNVxvdimuvkR39rl5T9fHlHOHbS8
yWul48GCjZFR5IoAZ3YL0rdatBT9L1YxjnFCoyeHJIVHdK8DgYC4Z0KRcQiyBIFFTnfiiVWPOOhf
cFTXssLJDTGaMwPj+eMTp5kv1yhiDgOa9EfI+jg9b1kWlKUKh24KHJcdN6DGa/MiZfud4qnr7Ckk
eiercFDsmuQNtm5zMdgj/mF+fpKSeHk/gK5HEfZ+eoboQMhigRYaNO5qgbz5PDfiDm7JE5wa2DFp
qhCGtJmw6vv1s3+XXQ9po4qlmdQJpxwmnlR06rMRqBD+X+ZIfYSL/mk+uCz69h5d8wLRpa0oAPGB
osCnShVOMzARoZOTbyNzxFWRrN9JShy7VN5FlMqUgctz7WrOQojtYz/N3lc2J6zWDCVKtR+1mlZV
iz1WBZTKJ0xLXQlyAFREi2IKhxOz/sc1VDRUbeDkO4JtWenz6WZ8FkysoptGAMZbTHojR6dfL052
3eE8ITUojnDOlYr6j1ta04RbO9kwBkgQW64V+Yw6qj5GGNw0Y1ggt3uyucE/ytw0h+NM4mSw8Cfr
YQOCWYWXaxD9yu2TtEVKwXJN1DnVTjiVVE9bYrIRbmSxEejmmcVzVaqx4PGdVra9Id8owaL332Fp
kWYkDTPo+5lvEkRmcMBEi8/MAW4BIZbCCFzFK0RT+23MqEnJlEol/Y+WBqpKHjExiIYj9hqSndYG
t6a+txd5zq7tWKuMPcuT5b2pR47UOAf8VBEUi5RhcB8igPAApnlfzIIutmtjtchRHf+Lat77YDWs
ZCiTvWdw7ni4Tu5JrI13rosA8If/P9BX4NXV5yqaLrPmoTTJtRyEOkBX1d+SDoyyYvH/RucIxWxZ
mJUvZ1hhs0Sl+IY5Hwc6nkZMwmQNeiXtgQJFvPb8utqrgsUYTUA/dbKf9vBvflsJIYnQtvjOnGoJ
H5/vMG+rQGAKbawkoQu9oBbUgyyv5UvH9kLdpSMRDx9peQxscL/98IvmvMIHRcmGusAS/RJcUaeU
l9UokCdGAIHCs1gY0UfVkiKlP97V6T6sKss34lvtQ7x/dIwNlB6QWE64ggvxZb4EcxHyclHxiQRB
EC/KtjlnpxvPCb6hAXlwzDHTB0zGHoUdASyqTJdpku4FZgcme+9Mo+TU2gfOQJWM7FrUJKMLfhW2
l6VMhxl6S358jRfPcsUxQCkR/V2rulGvqu6O/PYShmS4ZaIJs6kXTsJQFNQJCUXuABgSkOK++akY
4NeUy0uRO/aOYl44aUI90hvh23rlSySRjr5dmb51Bp6YtJvEPAVcBtNKvgSEwTtnsjcB+l7cWucq
O5rUCJnDFh8VDB6MW0ZaLzi/+vPSThXDC6KZS7guUdZCXzX8nMDyB2i/lXBpCnhSQcltA0SK9piI
heYRPhJVk+gWBf3QLZ8ywmaurTjORu5SdoEvJBph+oybAdG7y1rRcQSFGGn+BnuTp9mv09Kledg1
RNbzrrG1yJIKg3hYQHaH9aAX3pSVMIfe1O2zcEmHLPBIs2jpaxcpnEuId1lfnN3IaqSGgkgYjQkd
qIc3Upi0iQiC8H9+W1IVmAs4y9s1taDQR9UMExukvTe8GcHc+Bfr6eaZXSwf3BqChsd6QMscMyjI
QlYZ5dNg+K3ksLlb1usexPtLaM8AVuemUyr27jE7avJacctdbsu/eOkw75zmm6EO5UYfWe3IN69D
6fs0KK6EQI14IXD8Rgq/49ajVgTp45JMpj1HFlgg9O+ByjB+ENGi7lV5LPPcvNW9ZaRxe+FN70Th
jhBddF62HBRdXxDrNH/TRX9oXRen2icPMTIpcL1iSG8HtXO2kZvNf11dlvJhvC53p1j5gTPs9Ke6
KwJEvIXBvP6rSGOUUTD0mpmF+BFYXfp1IWAMv6NvGXOgQ/X4Gl42hGXVSaFHKQG35N89Kz4YHDEc
adpmiSyZlOZ8u4ZQMZ835/+h626QDOaOZnzt77WEqleUwPUDIcai7349fa1ANYMNyaOZ4j/mTjfR
eQ+K95LqV1O1GSt25SB9AOgRvwYlTUStOrbfs+85KgDh1IPdwBptUc8J6jAkE142as8SgEz4Cqat
dUqSSCMLHcp/OBeVG2sikPdTnz4hD7MI8pV1bJvc7tK3RSp5ircJCMV/PuBRIbm9TEoA2pYrjVoD
0oC1qQMxOsBYybU0F3MthNgnpeEzHcu6uHox1VUU6BRqXCX1W4xF7LN3ik/sEBzPFttMd8+moUX0
iQZmBhp56fZwl2wd1d8wIfp1sys2TveTYJevWRLrWJyHkqLUQmYX/J1hiUKg6esxfpjBtcpx6rUr
nABR6lf3D6kB87z/8xJbvemPzfWULpS5ph7Ikr1t7ic+Va1cBXFfEu/51d4rq/iWijjTJcJBa7k4
dClDNCGPqZQhECJI31HAcTtku5sVQ2i9VW3SwZX3g5v0fZ5dzuEaDO0JgwuFuMMFF4OuhzYHzrJa
Y8zIiHKPZtOq8XanhnLAn5SWQXFNpFdnJv8PEPPF88xMZV8THLWi8A5ZTb0l/O2OM/gRRAJogWR5
ErP67pK6OUp2TaJXoS/y2onRTGrXtYkXQiBQ1/qL/WseGeaGDx9uH1KNPstXsuRctgmoq+Ii2wNw
BJxnDW9VNCdpd0rT41YasoQWDI03WE45KGrlwIvslTzPE920SYsMd+be/beUFAeuOCNONvbUw5Mw
v6og54TYPK3po/2XipItYfUMpydzWwV7C2YEE9RfyHBmIIlAx2kANj8xtRLAgN3NL0cVOogIe6+0
/TTfFKh4ES40yqK90gbBttLErzkJoL6KcrDebwpyn57V0R8BbjA+gZmO7wB6jWWIPglr+UPlzoQ9
iPZkQTYKVEgbe8Mkj5jO7jsZUu4QAztOeJjCvuy+xIAs3MIIDe9Exa0ORfWqgy2StTrCaHlktQe5
05VnmduER8WQN/broSdKfGYs4u2xCaf+N1ah6ZLFNG5S1KDUtDb2W7hrkNB/UzWzqZ1NoNDBvIEZ
K+lbR9AzqQTie5Z2tFrGYx0sZ+JhLDkYBeZ/KQ6wJpiFETEoXqiFur/hgbXxhWtVr0ysoT/qW7zd
CC9BUI2QhAQIzATjrgWf5v9arTe0uQhShtUZxuIAOUSVWf77YJu10S4FpuEh9mZIxlzTSfhCC1h6
zLO7Se2Rd7GRIBlz5Xu/1L21TzOHMt1P+Ise5itgxXHFygDiI1aK0pXjNSoBScoDZ5LpQwNcNr68
AmwcSJzaYuZjt+rJqOGg975rChVqM66FLHIFUVYus0LikteOKBql/XoZ1y6psL0BdUB66caqceEh
beCVHJNk+C8as9S+aa/ClGS8K9pvBBO8OgJKcT99ZEUUSf0wK7jsZ7+sQkWFzg5iA81YsTtfshTn
nPOxdyxd3utCplIJVxf4pgwkiR/S1cwTEy3Yu0oBqQ3XHHmbjOWtfUx4BWD+DFEVFgVdn51EfXqg
BQv68cO8Y2T/I2jkqp6XgWc3O1qgRa3e4XDsYxVNYFyi3XWts1wCpAYvTQcbmmKnjqiIrtnTTcr2
v4qmIC5Nuadfvh7rxbF8bwqPV9FUedHYKxsFoY5SnlIMAOlr4eFDxVAHX8cvfzAboAp7G1McES1P
JZNa9oxNl9uXcOX25uWIA+vwz0mtDBIZBklh5jHti+8efUzgUhnxt9U7PJ67amPBj302hWcW8MEk
4DOwQcD4YRMMKJocKYy1Uy8SSFbKcTIdafqtRUlNxHNOo8IKcA6L4GN37fjgwI0jddd0XB0o9uzl
/ng/WlI51bqJx123Ki44t8O0I+OgW75CHwelOiblG22i8tLyARVUcmolMakM3DYweVatwPS+o4kY
pJoiPtKH8syiWGtyVJM/yh3090qKqlwjakI1pKDU+ZgGIey5UPXxYjbplYNVTqj/IlnD7X/KHy57
2owdWbi+CphGC64rB+c6Mv6KvQgbnft14IcNRM3rdCkyGECbcSGJUMEM1EbMQsiuPjDqEn1xcZL3
T+di3VB9nzfhnmD7x9Fk41Ya0aoPcXFIlMdZVCBZS9YFhC8yttQy850H4SlGHbMg67rTKsd9cMJ9
bwFMgGLebbmxq9PfEAr5tCfmqmrdpevnJhlJgjT4ImbDSoWF3TIyEE2PAqLVEd+pht+yy28BvakJ
5kHeBC/BDjw/PRL/LCfOUg+urL1w32g6GMYeTpLrB+U9MOg+jgk1gMut1E29nk0WNJK1WaNKyegm
LDi7KcnoomDmmH8EMeBH0ugYSQelx7DTXHUKwaHK6mXCC5uU/LQkDHMDpQ8utaTkTZZ1QEUu+uuB
/96H791hUiAIxc6oSoaiYf8M7TsyUGYKXS7MRcNL3BcQg+qLFiAhN7C39cYBzODOj9etgk9wT0+u
c2wobuQgW8iPXgbMQCyTf3DZrU3+WcuXrdtUWFAvbY+8SmvQz+HogCLYRUeVeBhpGoWlrO+aD0yR
BenvSvGC2ePGidRrDH7FnNj9w0pP6vyylwNoYP4o5AEf7IojQJ4yVH3X8HNsgnkriqNdTZVJJ/5L
EjnfAY3PMgGnNuI4vnCWIaDVoYzHPyy/E/S92wuvL6YrB0/0e0Xl2zJJDfj6WpwaPwtfEEViNzcm
ZU3obP0ObOuakX3fWKHCHHDEZD5lHah9jZEW79Vrp1RCOzXcyJWmsMbqx6BA1hjJcOUsEcnxYkCx
Gi/Xa3ij1AMJKEnaePpR4L5K7skKkqwdv4Q3R8rnT0WIUW5UM/Q6Oe2Tpfx7GKP1ZKNZOZpuyljE
coTfCBKchSFQDaKoQo1eJz7fYqo5HQLs3xRQULSn4+GxjXvLTa2VE6C6bopkLNKpPrhb5XxLKwtQ
5uuChYCrfSuYviGgKOS++EJyTHREZJxsqcsRWnZZocOVwvE2a3JALAB50UIc+F2WbHS/cuoxoSwZ
8HqV5m+23hpq0B0Co5QEyu3YA4aeLmAXvDd2dEKGhgaqT7mB0XSY3Lgk09kU4HJZ1Ljr9OgGzEDb
+/8+zjLsIdRJNq2Sef4sklMUoG7olkobscD94wejKDYI40NwdaR7foxt97sTwyEOGdRKF2Qu0/V6
m0AHj0XAZd7Usg0lBXLs/hiY/GLdYpCOacA2TRddhbytCpW8togJOzJ1x+wt3HChg7A+VaE0vFUo
EeJjEH3uXuosznCqxxmKPNzGhL+PA8XN8RgvJZ+1yVM1xEBtDXlIS29NSKZWlcND7sZ6wnvDaO5y
QQjwq+IcIzhJwx+77r/o9BrgVpisiTOfRMLSf8SU9G3uejAFqqsmQAIUd5GwTMCDKsiz709ToMy/
XfaOZLj+LKgTg0JnOZodH6qXxB4/vwIGWbcdsvDB2IWs0XpwkSwVZ6lAEjXXv/s+6TzgBiwRDKbC
hamhzn18GPBJsNjuU59L9lUjXkl3ZVpdgtIH/SSfIIZc2xLMT8xRn7KlFTZqydbDbpa2W4bSz07S
s+JfrVhEF+cMKyjHi5fv8syqCzaqrdptx6UDATmDd40Sfj4KqjZ3VIQOD4kKVP6c4sZ1SrWrhHhm
rPpFxfp5ISIqiG4RUnB/2fTxUt7SgLWcGu3D2cBmE1+vk7HZyuLLp/AWlwyErfrF+CvCnvEjLet8
lxu6juqNQITc/inpS1pfT2E8ZxTDIBWkcWpFv1JyKt79Cd1zi+A0T0N4faWcGQE0tzgsZDXQQZh6
dZR1txUlISAFBO7UelLeuQxpZYmly1k1g+LNb23GTbVvBdRZtQZfNx39hrXKkCArudnViSGbJfL2
FKitViQKC6po0I2Fmal1/pnMC6f9LYTPolpGm2PGVcSIL/4eDyZDmvn4ZKV7HmrGWfZx6RJAoSJo
6pXi5XMHq3NZ0ls7PWSeZrVfeisJYmcJoq+TNZ63rLDAjpQuiASMbz0UKGh8Af3uAyPxtseVC1GK
akDJaLH/jFMC8Ni1XKgSXn5jRHR5OTnBl9DxbsIVMdCu/4puVjMa+WyKOzz+OH3GKrcfEG2GhyN3
lq4sfXNdVB+Lu+9wwDF5rrZ/BMBrDf5qFnJCdp9v7cXoxZtI+hK9DIuaGx5dkZeyuGXELHKRmfP+
i5erjXCRyZYDJQfOhoH5ppWBxZ2uG5I3+c9iusl5FdZV7nsf7ITu/qIMmSmGS1DWfFmFFecf4HjB
8Z2tmi9daxV1V/pmI8FaVRwY02h0dZ9Gi1epq4kyN2Hp1fFHuRfAw/YoQNfYr3j5VGayQgU8i908
OLPO7un6X5rfwo3ys1HTXDU2nOKYvObZ08VL13wnFkiP/Dn0OU26KcCQjCnUn8eaOQGCBuJ3QSZR
qo+7vthEpa0T85MACc0ixAgTm4IMXO0VbijhTQtqxx2Tvl0dZYiL7anIEtKQM7vnRkuHrVZZG7sg
WWSksUhSt3igzwHt3QtAaG9xc/N3182TRv9p12SmL1ZHPJDiFUWAjlpUYfg8e5sAQ/b5161T8fcH
gdDvsh022U9I1s1c1cGS53CtEqxtEJPrB/Nv49vOYc1RHENmsuxNBq0bHqYNZ7blBPhYEw1Oz8MM
NXZSXCqez4yXwjWu/ULLkShk1h31sNIAHQtJpv0lgiRI9PmZ/LI70eY26UQE7aV7PEtRvitpXVWV
vXyPjuhf4x2MJQzpodx6t3oBw+jVFkHG+n90t5FtYR9bTWGiLa85PtuVIcjc0o/ecD9QvK4bT5yf
sO3qi1ZyNqLsQr+XfLWUH2zeom3bghKmou5l9Cv3HjLlKDSfGDbOCM36/9xlCCYdz1DKq+yTVmc8
rshAyW2TKLKCe3sAsfGhiDSIRtezlkmk8qAtgzmXJxLjApvehtDtK3CdO7XMWBFwjBv6O6GJQ4kz
7CtEG7dZJ2+JPxD2Pw8b3YWSvRcOIZPdVNSbat81YKgbrFH1L3LJrSlMoBz6VbLY+PI96Ghynge8
tiH7hUcd0tQ16C/Ox1WnBVAEBiYxsPGiS2BSB9n+1aV9uBdwPuYyW0phpQvApDyfoOjMKp2N2dLP
tE6QkcfBwJBOWJtosZjUyBO8FfmaliOkIQzAntjpegE7xKazFxBqrZJac4H6nTteQYRapy7rftpV
bZWoyNLcJlTkHr28wJ5UUYbeIS3n0/HguekIvuT2bWjwOeC7Vckw8m1pHzaMy18SooQEOD/UguQP
g8fSzJAIdxMtk+nnu73x6+bQtaF/0cAFtqLJjCm9DhHqccFVUtug6dMZh7HfanlSEmpQSWE/03C8
XP0NBQaLvw/NVPb8TEpywLdQdayeubEJR+CbBmcqScs1d9LQmuTp/is59ND9zS5OaOs0eC7Ay0sI
GVG8r7iJEOAOPepL5h3/mvbYBR6GBsvhj4Qtd5VD2OfvAwnOkq/TPTtBuS8ELgqA6CyCnPr4O7B0
c52TzMMjJCWsaJpgv9IAI1NzYRh9mYOh4XUCzefPkcFb1RYGNI2TVP9rAX+QniyzL2SDAyp7Vbq/
BaracEEwifyrEqQIwqFxPu4n0nkXDaon0KB15NWX+I9Lxq77d4hszA0YIjU5XFY1zeT54RKd8zzB
SCYNZdBR+om5acCtMvOzHQWO/DLQo3xKj/E/GCBSvD+BLhA+LCpb0Mh/VD5KcSceadaaFKdCwq2+
+VQHCaw/RiUjt5cNpfEhX0tEA66mnPg7JKBFjkGjw685dC6WNs13nw7lbRPnhvgdj9UbZfHpWVz7
1Mi/LhlOVk5KfmZlq6ZHQ4oQ7yzyJkDUFsb0mj1OQ6CWN0EaO9Bv0DvMH8PJGuD7i1u/BryMAVYl
R+qcafeRKmwhlT8wkH7f4W1EKVNd8rqmiEbJgqGU9XYq52TzywNrGfPizFSZLeduqC0XwHIJnkvo
UrTJIE2+twqnzcGhuebz5UNOlSZrWJgUOyMCFlvTgiYx7Lv4Of6KffGlls3Xs4F6KHFXE+aKmUWH
JUKyMgrbonFTzT2tEcMNNaXfCIaOmJaY33IZl1Lioh6wrm8POSvcpZuwg8z+6b6nyZFMHSwMXurF
g1gKXzBjZMil3agFu9j4gddlZD0ocMAPRO30rDN8Yy5JHw7IEoXmG9DmX/gKx9kYXzMQyndc4yh9
Ej5H+Tk5Ed5rZLL/JluakyHP21IFFKVhWKqRQggXHBvuDCDzx7lifpYcIn+CmGgMkK/D8RfCTNW+
UPIEgIHe7E5CtXVJPgSgdNuqUNKuE7LR5mF/+rvVEJJdsSl/rkwHhoQdkrkD9Ov/aR726LbQiASG
SphBTyU9mZpOQa+vwTQvGk/Jzb+IwMLs4dEq5UBnNuU8OuJvey9xTgOLTpzJKmesaewvKoVY48MF
ldhViidrtcd3eMqZE4qqVmLamSWhoiN7FG6AUNnjs+jYzf/weKkd6m6JpGTSBW12fdJzeJY94Mrc
MPdQt3sGuWU133Y7qJ8oWSCGvlWVOIzPks1AET+iYEjI/XG9ZQzgVzgRr0xi7Z6PFeBc+mMt5zjy
mhK4u6tAv6++QKAm+qovOj4j9r/aoucxRmilFKkAIOa8zjjfjy56QY02pbzDSIaUmNqbEtbR3Jac
7uE0lf1kXVOu6s6UjoewciuNcAOOyAmvTOuQ7NeQ3DQuPxOsHXozqFmAJpYGLE3ZlsKmLpUopS6m
TsSOxHAPRN/3tdu3t4NIN4/q+b1qLxWXZ7cQ4ngc2NGoD+N1/QQHG2lqO/SBSXsOgPSkMdhN4PPh
EKG0biaPkHGLfJUNqvFe+fXkQAkqgAdFbpj5kxBH/2pHtluykJEw/7gNEqERNUvOwfX7wyHiaF+u
phb63Ga4DUmMomMbqzgEPL3KZFLisdHAtgd73f4Dn94DSKl5Wst2mNf1zPhNgaxWn3WAAoCr2u+E
gNYaK3yntEyS77aGKCR/j3gMmirWEy8IyQWi3w3zx/H68SPtyODeOqWRLVEd19dbMDKa24HXC3gt
dbgXcSpJwSGfx5vdDlI7c12Qy1lhLz7aS3kL23eKP86YZoZbJf04D7wZZCeqhunrd3cdnPgW00td
cCm2tAdFQ0m2gqCB31OW4HwxZMWdh1mEUEAHC2PHdu4m28licOdraDshk1iwepTTqrJ1bIoAE+kl
5E5z/MGD3V5kNJld0/JXvQOJf1ytmm5pWAq30TSI5RdJY94d8SjS6fCJSTkL/Du3T6Q63mZT8PtZ
X4K8+i1JtnD8I0iNao/BRUgg7SGnN95G/yYfIBnYhlPDSLeVOnc77Mku9sUTUGp9dm4EOb8qYJrv
wcUsCCs2Cujrr0p4nDSeFezH7U2iWWtyLlrI2tLX6iCDYeUpkXXmp7FXu3bS2lUuBJ/zhFCsh46k
FzhN8oBamdJCXF6ikYzU3H3IFdTjhEvffgQLfhRVL+Rqk/nMw3UeJqy/1dnsyPZ8PVP8sxMzQg4i
7B4Ta8SkQ7V6C8tezUJk2YalDCgKKpyN9S2JrQc9PMsCfqdEunq10VvPB4dlELCE07PbHV4cJAJ7
VnEclMLvKN/tUKIKjAT1ycnYX5a4jbGzZI6cTeq3HUzv3oyPKx9D/NY8BLByEAwf3zRrzE8S331/
CkrcVbb01FkXD4BbM1bdhrXERe6C4IV48/PWwM4I5sXyUsqS/rZbh9MHqp36w1pTKOv3RuQ+IYxz
Ce9qTT9UHhyPWbLlhSC6066ITfSDwujVQ/rCrK6tV3hsUqLvu03XVc735k1kTyQNQI/mdFVV7TdN
LuAht1s7MSCs5nDWyFOJAdY/sZFqWHl7Poec9T4loAsHN2XFwvRNHThUCLmd76RL9zAmuPkgB3pS
sQn+maWINDksE5EShSroru3XlI+4vi00aASYqSPSwraxbGi8w7h+mtkUi0mB7fV7m0CAz1UzUUle
DpW58yREElstBNZzOcomd05ml/CEYYHneuW8VVRLMDYJ/tr3GGcvAdwfhLNVtcPefpgf2nl4jLNf
nCJL+8thI/tERsM1b62y55QS3kmOiFkBaMZfNECysaUlhtDKRMpeZLCf4q4hlwpDuuD4E0+1cBM2
lQ+oY0V3p88VyD+UAympR3JixRgJHkion6ZYG/aj6VDruSojqGEd1cpw+0d31G6rQYGHp6yIsAyL
C+yGi4aJLJS9NdcmiBgctuylu1Mf56lgbYhn8DqqL/lra0OeWkI1lTrja+Qr0FRvP/BXem2OMMBI
sSWJv6Bany6UhBvquToxsToC9BMSLJ9N5BUlaETiSB0Y5EmeUz9kyqzbpnbNVHh+KSGXnLw26q4A
qihBRfLxgyqhZlDFhr7SschO916enKMe4WVHf0s8CnEfY+9WNFdDYc/t10/W6r5GmhwLmiLpsrSt
QQujaEyzWuhOL8BoHhAZP1g/owS5x1Cwx79HkMnbdneGGDkIONbeqiirzfvmBcrOy5RvHYW1ruLj
eUwiPXEWUDPu+4tc74Pke4+woLEtJj4fREIRAMRtgdPrHBh7nPv91sY+Jphv/r/Lm+Cz1bTeP+QY
chYHXR3Ll+eCO4SjSsmAKiDj+YQ8RF3UrAI/nk8E56MWD79Eyzti5v4Osl6Ry0aOeukTm0E4fwmL
tB4tVEoTSEC3mduoYNUTJXPEFqboNvCC6cv1aF4rc3rGBzI6xM7LSqtbnWoalGy4X4O8uISgCSrx
zYxTDpAcZ5CeRzondonJmiprEQWIa387KYpLS/Mo/nLnSLt8WK2mPhPjSskcWQVsRukYydcDY41c
4FjoRikWlVp7k6GJHXAWMqKx3eC8UH5Jd+EUZGBmohkcR7h7utyn7EqLc3K+LjLMUipl18O6Jis4
kZbBtVfviCx2Jh5vzkzU8RAhrCEBcEYTRkjr2Cc+k7NNh5DIjCacqxbtGESRpNaNBytst2m1/nKE
To14koQGR7CVWvhQCo2sia94WIBTHP05l3BEutJo4/N1+kspJssNXR3CwIT7mKGswYW/rQiqJtow
KTENQSyBkkaxJ8HgSPgnfK4ixtmA1pa+wSMHZ2oeUkHParJlAff5pPw0toV1wvCDZJs+dvfOdwKS
hTdAXKd4+vUKQhTasnbSAv66PXBKzokraySJ5AZUOUELXSICZ90W/015IeBPkc/GUjnGGYhXfhau
BjfpoV9QfIcxWhG2kbB+hvjM1/4kmGIbbBVGBrXTzfZIa5GJnu0Dl10oEW3J1REZfQIk5CBe+QDO
a2LrHM0H6nXit9eTy3W89LcANi74CcSDhD81iQbqe0MDY70mJJxF+jz4+V0lS55x8OjKdATk7XxJ
U9/HylAVnLydu6lzC7zYZmWkrJTyTPFz8O9AHxji83lOdrhTeV4ePbmRG1AMOZtdwShjY2PunfLa
ZiN6UJx78oHsc8kyyYSSDLqj18fqQZ/ogY3waYL1N/hjmZfv0rpgPjKFKgyQ1Rrj184BfiwR3kZS
s+YDITs3EPEDt3t1RMprPkUF6LHyT1lxO8fErABsDIoBebmC1w36rWM0YzGRyaqbBvMwBtqCDdwf
I1gHfz1+6a5YwETECMw+YHvc3oNJMmtO7M7NblKwZh+J3VgXezYGd7F1P9ezEJwP+aEem1zHkOsX
Iah0xnoS3imBic3S31u5jJIlyh/Xs2Nqo5qFHNWgcgO9qOqLfUEbv6KiRCJqXxa21N6Z/oaN8R3Q
Y/C7YRY4k6EUCbP0LAlBmM3bocThT+JnbN1hL/zJ3RalghZi4mjopvhofoMGmjOOt7JsmggkPtmb
9xO/AqBKTdmVXEqY8q1tk0QDhl5No69dCZhTdfdvirgCZi5ZK7DwURbyhiMmOKoe/i4SE18yal4Z
eFWuzfni/7BFVEMtC8G+XY4p60GIAl8vdROgvXnV7MdShoCJLYeELUvZVq5pTat92EcRWpVA9eYy
prdfEKDiL3fEu++UVOs7UOSu95wiN+jxsqYDGzxmmXVgyp0rm6JFpZWwfVFRWiqb0TwkkZBixa5s
0ntAs+HV9XWrQPQkHuTiSvP/2eqDOe28slrQAqLHn0BS2DXTZbQkeV9kVwcaC4WpLUAznmKtD+Fr
sv2EDjZIrVCygF3SytixowAHM+LIqdoG7xqPlpAy6hjwRIjSHyoSQeZHYBw5gBrtRVzHtiLzajWv
0Ih3kaLGRYuMzbqrxVgwu4WaZf5VAOefN471kivYvT6S46NRf1+eQESKgxcx6I5B00iCOulwxkQB
6wo6giu3d4/AaaW3BLQvefqlK7OBZkRgyknszGDtkHVJbLrGDUcaQ5Et2kRvJpDdokby6+23k13p
gC4SibWGxDmGGpk4w7xWOKhc1EuuQ+SwaOZPsodnL0wkK3OGp1JGllhTSj4T1iLs1KWzoAghG1/I
71Re82wwGVDgyKNs8zaTb5d5smKz441aRZX4xfSGqxzDhTdcIvxerSCig6zRWbyaHtrpYS8Pwf/I
r1/r/Fnk1TemWGtH5mgyx/6LHTc/+QiGKAq7hCfD3aR0U0jR/eFqva5ETOB61W8nOW4sYo9HYMdu
d2l9TA8fvDuluXfraIGVw1EQdivBHFyPRvy2g5ZK8LoWcBKkY/N+04QBg5il5qdeFiPdIZvmvpRl
UnymeK5enh0QWWEiWGQsuDVhCisa5NVGB6ttc7rp+iTMKXfPX66Be8+2pV9iuPFOu9ElRgvg+3eJ
GnvY/3h8ltEzms5wfpTBvQTAh+Mbou88Ds1vsQZ2W88cLlBu++d0k/jS3is0vXz/sTg92mU+e7lu
1dFGlFm3yfxA6nAbU7ZyGjp3/9W9To371yt39vLOPF17x2HuZih8AmuWWJiberJdJ7B8X1mbcTsW
3+c7sKLFKJiKE0xMJHhmLsFdA7cD6E0CDZ3uAUoc6xdfrAuh9dFAh0dOxSwCoF7T52rdPXcZLJbj
FiomZyc15RxCB6n9LrhmGIPV3HwEw3hUAHGNQcuq/bZ02+taAwbaKYLYmt7ILYOWsHl5sspRmPt9
inTa/cBJXO026cZMq3FRAA0Qjca3q6jrkyp8ZJU+krtKAcYw1D0X895Ao9mcOfHsx0eTUJQoQKNa
fmB2o8XnhQOcG/5EzuImpsxN9DvUo83Uv1b9vV4vtDFPEEH9kXkU/wQ4QKyjMQfk5OPRk5iLbHUd
HbEm/YAjOhtR7FutGC38sQlsaX9lSm9GBZVJt8tKphvkC95tGPC7UOeldb7ESuBviMjRbfPtfeZH
TdZBVX2mnabJunWaWFEHQHOiNYZD3r7CEoKkupf7HguPugsh/LHyGIAcVEZGbZCetTwWO9+HxPMO
mCHxsYKsyEumc0T/43UCP9SVRTPNxT9FLNpdG0kjzfPKpDh2+BtVkxmVj7e3ofT2+mJckxweWYH6
6Zz06NBD7AMK4q7V0zoKdbLl8r+7VLa3K7/xGtu9YE8Cavimm7Q62kDkV8CBEXokBmdNZVSOcyg/
88dhgfp1CoCTaLcnf0b9u5tiEVHI4l+0WMB0xtQ0XmxLN0dv4ubj/Qj9vuoWcm4UvFME5sHUbQOw
oh/i5uIq59PlUabahN/XU+Yz0hKOYMmZhC/y1jDrgOZTxRCbUXFUoAf39UE6bFjngOmzEFuqU8q9
vlrq1Yn6ePpxieywWpkDD+44cwxpPxj1W4whMmkGeFVIgkMdNSq+L6imxEl1gH+pmcqiqq3m1Jgv
0Qqfcls/EQKkSIpWvndoLlQMDbQSTfxMjLgCh07dJPczRUAwUzdG263LGayE7JUjG02E+JQ1+vOo
39tvPSDLVmg7DfsEj+oTp5UIBaDIxLED4tF/iaQgGwyHBHmH8IRHoGkAQxOtKHwsmfeAkelllmhK
A90Sec2Jl6jwlE2Go8+yEQBvKVxNp4aJBNRxMzjcGSy3lUDji5nV71cSJBB3VinMyz9S8KILVLG0
rGj51/VPWBrzIrWY3UrDKHVxzsaJogbFLCJTMuetGJ1s8hvg1wbjhKvU8aCGsNkgevG2ptQv/TuX
V2QyK/2n0aSjUg7aI6dRvz+rO8i9sDVuVgIi8Dzo2qYdRoaV0OQQE2FWTH7+p7bSTnKttj/XMzk5
BphkJwtvmSSp0WoysUlCeP89f1yL6tMYbqoYn3lirSi/xcMSVFQFAK8ePAB/BlXyEWOjZ311ijcn
mAupbYhZ/kCfl7tAKdRsO6QxMEUt/UeAs+0hoLUd8h1JgfAOrY1P0JQnruBS7kBTl5Hz1EO1x/4w
ryT6LhlD9CHZmhLTQR+EGN+Zz+IVyrIUQqA1lHV/2fdchgrKpLknnqgVnHJRhXK3nP2VO9dJRLUD
jwH5+jj+SsgvlBmj0A7Nbn+QeSSV+IaywP8wlC222wRWXdmdddxTT81AZwObjgVt/1r68KNQOsp+
m1hmEM8YPCspL8rV+m/4co1UjxffqCnAjPx5Ai5eIV7pA6yLEJ050k0nw4uhUVXS/ukoanxeqzP5
DHdwwHkNvvvKZd7+oWF1xXM/oPZtBmA923/IGsohAdeutJ7JAZfyWpu7cLTRuuwvY//tqOhJKJ82
6z9+PBEFGd9DYXHxHXrnizg2ErBsCU+2op8l+vSY7Z4l1KFztXQxkGdzLx8WNwDBIsaHNG/TeY0q
o6q1NiBQdtho4oP3fW7MROJx5dtDg8wBVfTfyoCJ1IuiirFkwLcUdhH0siffZ/r47DjF0KgnV73I
MbDJmc7zGFvfAa3ZGue57O9C5HWGSe/zbjSMPT6dqOq1yGBXbU4DmBZyjKjqBTxZsSq5uo6f0miS
3dZw2kyAENYltCERDqBh4yrGjPo54oTrDAa4s+E872nSy8TfudITbnxyUvYUIlm4R9KKPMta/SA4
7sF0LsyQTtyn+f1uQc/zq8DdnmfWX8Pzwjg98gs2uhyBHz/7SYt5kPhxAmbGiRcjdLJ9+wHdR71V
BZNf2TSlzDOEJDdKX8G2hq5Oo27K4GVoUZbF+Cvs1ekC2iDgReKQLeNmZbfzj+SX40cPy5YAgBCl
IzHqZrgyt8vfZHT2HEbSiE/zhmUyjhsVuRQlC910p39hOPMndVvaL45AzzanR3NUZhbJJXvWHO7k
bq9g3arWeHyblT196aJEXPg0l+MykzN8PKdgKDJDpop50hQn+r8TZCxPCACyjZgPTJxNQDqfyFMg
i4A7SElJQzS0b6koPIpRQL5KOmQuujWma6wQ/wuVKLQX7U6PPDR1eiklNz07NFSVsaJiR/PluCAI
va4cmW52YKbpO4TCkzDZS00xOd3+09HGLQfX3PpCPNdlYzCK8/HpPoBinhnzeHIylHM2wjvF5KX4
N3CFJdF5iSZ40CO6pf6xpQOR9qafGEmGM+KE6/0eEqCvoY7mPbs+Se75OV6fWJ+J6YXriCb2zCzz
4Ewo8P6F95zVlZo+SNCvQAEPyKY8mWTyuBShoQvmZ+b+utNdfJNEhmFEaeJSRXwG6mWjIxqVhEBH
fUiT4lCEOT/Nls3Ilt7V9WV00Zpff6GP4R6SPZm9/1Qa1Jaj9RhBqNWdMviftuLjyhZqVcRtrqwX
UWdfQQp5JeLxdu7n3gefkHymgLS8mnEdCQYxpiPP8RFVEvIDLm7G7qMb56J8+qiQY+XrD69kOPb8
43R/LFMzP3gcroCnq5CMcU7yMdVsjk46QL1ezgv4vTZTdCBEPtj+RYpyBX5wceKkSw1cXZU4Mx2K
QwDgwxbSOReGWW4oEHmbW12EobaHbmwzAeUK0Cu1Mw1MMQICd+TO6e7aiYey/Hhkn256qwLvb40P
blMUHnyt5ihwHOwaqUpC5wmDjGiKIk6EtqGSe5rxTS71oFxl3l2oTa/9Bsn8gNZGiGf2/ZU6DJ6F
Ble7hxKeFrxRaExjHve0phR1Xz+yS/CUn+HZqhCYGRNTjUo2+hGzJr0wGwEaGsRcKNViYnapEsNd
mMvojim9O1YN7XID41HBqM4O+1iljX/aoHEbcHA38V0Ulnyq6w03CHszO1FAyIqxHGoBlfNrUndC
75ctlC2p3ZTS6sC7QbqgI0j/tpWDPOMeS58qJ+8m+oMCcWKYhVnTE8xQ62GaIoSkiRSNRU8Ot9w7
F5ENNJ+2jpxdZ4e7K506K6KQ3Cypx2Y+c/F98cvEDqM9iuIqORKJ36SehN2apFe4ivldeAiIPGfg
bLpXufKvyvAmPdE6Mgeyl6FTzi1STPadhLIZBmHYJ8B9watkurSLwjjdmGAKRTuHxYiDppd6Lj2+
2ctnJZW/vDc22oo414Jn9u7CeaWFrIIIvIRTkAei7zVHgZzEbirAh+Q4In4CA0a9xwyhiwz3tbBk
UFBudSBOHNUDQXAMKdXwLChWXEoXRJ2tA0JtU3aoYDXyCiiuX/MQnFvdrfH+a4B2YpDy/Y9yd+GU
TVFp6FcSRZEKi+bO10Bs1hDC1MA3GqrBGSyrO+0Az9Y5FBrFl8+jGXXJ7SC1kjxPiVihHlbrPJPJ
KyJ5QqSs2vlrTp4HGK5uJvVbgpMzDX9jnCKyUCy+r8aHRFnQhl90q2cwZ5JuIlQZm8DmuceRVTOm
s5y3b4lxUERDqBSuWBvhs0zyXo3BpGAPuR27iKv60Nun/ew+dg6+brz9WyVfIKNk9M3nwkcCzYGb
lKUiHJmVuTGLcpD3ZDyhN2k7O48IL8zy187xvqnguYR2ilUCRxdRa2DoKSQyvBU7EmbfViBh79WB
6kyDhuc9QZWqxX4mgK781VZjyFkvqb475UXSZwwOJ5e9fWLVgyeNrc+OZN4m4N8ejjtRIE5H0MMx
AGjEx0/sRyxwJFC9vTtmh3/Z95CuYTFi3Bsi7QUdHcwjXw76v5iu6aDylIBkAcronzvrAvwr8I/S
xUbUdP7X8a0qrpDjgaH1UQXv+gX63MVJLCK8ROTWh+GRUBQexDUFL1Oirqgoi3JhxhpN5SxEHlzp
PkQCGAwTpC7hBWG40XgSvLEYEN5CsS/G9TgYhe5Yel37nq7lfiK/DUaR+1Oqw2Jgsfn7VfeygC4A
b4ZkiMXgqw1W7QxE2u8RyS5x/gcGv9ctc6KRYopyPHz5wvBN1uAtJPo3H47riBZlIHd8XPFmpO/w
Bsg1ub/oXXYzg/BooKBv6eVuHX3+3VFO04VTKcH2ZIfah8kMOofC0pZvTn2IJgP88InCoJ+Rroft
LNRL44rE6daIHhHNe2CsOutOWDSWtlw95qyBrHUoAo2UmOAa74oeqheqlPfKXkOJBnV8exE86ugI
1fbDa2waYiedzG40/U+Q4d5v89oJhkhQcFsJ3+zStFt2QQ/tzuhKlf8XkQZ3fw1JgcWGIMJUELlr
y47OtHkpLOzAYrKE3oBvWsCp9Cs+1wQYQX1eg8ox9dSgq1wg21vyFO7ezIs/Gn3ng/DQU91AS2Z8
v6YSiQU6HoAtX5TXS3cq0eHrHQqnJKRrTv+iwyEAq7Ug2QrT5G75NhKrt0wr+P7ZShq+IpdegNnH
qRh7HnkWLimoT1Lq09v+yW/ZBopUywoFWcgS6ztf7AbTnlDh5g9u8H2/URsJaAGL4N3YLH+1/vkz
+U7uWBT8wSN5OMEF+Whfiigk125RMyE1U52+biaYky8SS8mUntCIZ6emgqP1/xA5LR9COgGsxDg0
brk5N2XhbdYPCSpF0As7o2SJFdKXuPZNfITtKeOXRLicTWMEnWzr00ZHPI9u7M5yQwFQNfaVdpQy
oDXaGYXLtt7jFc231ERA1dB0mET2YsxiIfrhhI8myQr9S2dPXBDC7qwjeYirJegg9Gixv9matlZy
LuJE3boNosb9ClXpp8GBDtg8zDJGv+ERqe0j8lyClVubEi0ZEIM2syOi0gveHK5d40LJUyqKTbt8
HqS33Qz6jS8EhrUa1rTgZC+LYf3HLqB+/Gm+nH2q6Uml64kBe6Or2MtR+5QX3O7GbTAYrdVAjjyy
2F1bYbAF6v295hsA6d94J1UknbbKgWndxStccg5JYUvN4EohSpP9KU91R1LBfJpae4qItj0nCoz3
BRpgHanrd7rsLfQgE8D4V42qgbR6e9ILg1g8IV2uMQfxjcdYNorw13tMuMG8J147GVtTAL9Yn5gD
PMnm4WmKy9p11w6vg/+PdLl7J4+rhwrFCQCRs7C/Ulzwosyw+Ja3qQfUOtQk4ECRA7lW0WZynD/p
QQ2hs2+HvwF7zV8/99bEEjd2Nkoj64xJpeg19AtrN3XEjXfUaCbJcvzvH7BERystskdxebdoDZAr
ULZFS2IegLbha6gfbjZEFQDh3B+EV7yzdtXSxs5ZjmPyidrBI+fnIHO6XoJaZ9xeXTs/ax0yRCOC
buAUReTRINoaso00EOHRHaQ947gfdYHcLErugkzJDZEtByFc0P5MCPHx9XwKfOOeDgbDC+pA0b5G
ejqvKAHD/h80H88qLGG6i+66IKdwqHeNNY9pyccMP+PRV/Z9rDvyFsOeZEZmwvgsB7g+wsR2GTdf
bac8u0id644ENTf5hrNHjdjL5hB4+bEAbe490xgO5FTsJohMEZ/tUYKr3uSC9vW9QHBxOBUAge9O
pQNQezVNIZ5SoHL7oK+sgKtvEGViT4qfiMu1EpPdA1GnbrkbNCKlmBAM/YA4c5M9DCRxursL66Qg
4W2isdM/JxulARwjlQqCqlv6KxvfWySVD5E3k3LZT7x+iwe4irJJyNKX017DZd215lWxglMWRrd4
9/7zQvRmJ+Bo15IXANMo4W7lmTEvzvQ6WVT7v7Jy8dcsBaz7vzWN2DACcJF5FMF+6nr7JvPFtplc
e3Q1U1EQ+o6OGy/aKX6kqi/J6ZtGmlHutWScNGcWTdtzSVrc6YKuGW/e5pOYRcPRqKZd1gYdbq+y
0czCvqygjgV8pxtyYWrXulpsl5EIvOxDSD//o6H1vDZLEF6EV1XmX7NsRHZTmUm3r0AE62c5DEz4
zg6WLs8x5TBw+uqy5+X/QdubNhR9LDaSTSNdV9jc4J/YdofyXeupB6FVzYVLVU6qtSu568a2LC4j
ndyn6BJDgcNeYrIlzdONkZ3Tqhk4TbOAvipDC4yXko6z4ro2HaPKq3Ty0BJFOvu+Tkjl8Vyi33Os
atxDd4bS2ugj3kc38vgNJivhfoY5lLonE2MD5gGDxZvxboQiRjbEIGi7TZlapxLUynaMnTBKs5AJ
3uEZ0QFnhbKbPzOMp0VnaZ6C/ebkcp24J94dcMfqXwd+AItjAJOYSPeaRfure9V+wzHU8SdnC0zu
uzJWqnRXQOux1BK5SOApXK79DqHqpPID1PP/a3u0j642kAC7xWu2Gzcps/psFybCxGgjye+juoli
42gnXbfDMdQtZIS4u3ZaOQCBoQE6+ky2lndfN7hrzfzFmGsnIsHzqwuetZM+WIGdJH3pbO3qBSkC
DJy3AC0LnoBNpFsf+ZhgXi67bOuyGkPG+L2YGi3tmJ2uJi62mfrQezieJaRi64ZE/leRRDM34Ao3
NGy+EU5WkRPmRZg5i4FC5rPwuYT0w85S/BWWuabr7hlixW5vuXVMNz0i2e9X+VHMzj/Zb5PWvI8s
gdTnkI4gP/f0x0YtIcjo5tFT2qZdrJ6l4veRRautFk0DvzhKcbB2IaykRlao8Aosfr1e7/ovz9pP
YCEF1wdkliSdEsMyzvyApOTlXDsGpfRAJHghiIqVjZbdyswok+wsmPUqHv5Ym7VuVhEWEjMwxB23
EbRhnz/yoyIP4K+c3DenKqMvgP1QwPckezdpt/e/6EcZfGqoAhyVe6wiIjiw+hI3xLKocFE2XptP
9djDdC8RFvAmAWX1wRdfLi2BLtRAhQCB+B2226EeMfkLCJ56Qr5/LncL/8/S2y5/Atd7uyEZbGT6
OEA8O+MKYewvqUQWe684NoKNOZuXwTr9Rh189EkruliEDYvgNLGzIMQSUux+jGa1zgfcpB0hLS+p
R4H6YYe9ea5bUEgQKx+20nb6pVhoOEk2RampY1+BmyAa33nFiL2uLWI6W8rH6Gvd1ygWe+d6PY7K
EntMJ1BpgUe+9v/MEgu1yQBsXdJ7xgyuSjcajvarj/eRdQrlAzQlTGNUpF3pWTZIvkVB5HcBWN9M
pAWO4Rk67QkYIXm+ohg+h35J3hVj/dN14GzcppW9HyyXMewF936Mn8hQYnupq0j3Knzn2UaGlq1/
ceZHTvJfIklbEi4jMQ5/NlWZYipjehmUW8hGUWd8eAkGXb5ekUOj3B4h+0jHRML4lsstf+pi31GR
z6PidTzCHFC99OZ6ZzEUwtKOyx5LMvk9aYYgvW3t5seMglDkCNp8KDFUtlFh8Hg/I26xFhyCwf2u
eX1j2PVjBgF0atvZGed+QlH+vwjG5qTow/xP8y6qlUAhCKZxRKOQFIW/44S6UCDErVHc6FSS6T+/
ppy89kmzV/U25WQ9fXqCEjFEi9oNsyoyUf+O6sE5MBx1L1JYDMpp3bX9Vb8U0Z/8h4r4LQcQCEZO
XlQgG0jms6ke/flf4E9hxvnQktN40hho4dJrRMTX3wdOEeHkRY24BSCOZ83I1pMYfbKSdsr+Lgph
YPmYN9XXMlVS5KS8ByY5OqnN2j2BLtJkQCdvyWrLHBqTZ2f/KXDJnP+njEK8gSW76wnPmwTDfTJs
kVsvAkpFw3vU0GexXEU7t4VZrCYPtYM2kHkoS3fOt9P4h8pBLGdSLUAZwh1fnP2pMs+MvmTxMUAH
gsADlA8oldaXEOnOcklQIUBgM0+xnq/cfFOPhqUrMJVuuvC3/VnhO6yQ5hlx4dFzhjzyFRdvTyJP
qnqIDgv4OCQNnbJQRmwy8dh7IRjMf6zaNFVVxnJkvvrILdxhudLsuKWgzATv9JkjCNnRHTh4XtgO
nn0VvgsMFoCn1oE5rTCtjSL/hbdgcqLT2XySQdowRc7DbTSpLphX91dlv/R8I5b9zmcxWinUwWkD
fNXwyYyg1O+u4sumDcFzXwedi74uHDKxSMTxFEh23M+tQ79qyyIcB5K0bRxF2UAGAg9wAVcNDDK5
lcnHMLLXI5z1n8XT301XI4LVz/IgacuyehPOAQ9rNUEzP37F5TrMB36SavD4d1S68I2nJj7DdEot
A/U7oj0r6tVcXpWbSkBhkrVFrBHhJNoK5oGqpkG/b+HgZLFNY1aYYdIPLsEUpNHUNe8inS1HPx6E
N8W9jBLrLGzj/iVcN1DzkcOYdlamTTCvcHbjjh+TzqZ0A/2cEYL2KDYjukForIouSxwwqqpjl7nV
AtP+ioaGtpBqAGLJqv4fcMDyUqBVUZPTeRS/1SaBHVXJFOL5+CXeVoYhn+rT4L5cng8KNFBACUza
UoXCRNIAZ+zp8wuacfOZBKSs3c23uXbXHjNjrU56itOZsIedc1QcygqtZWVeDnqwcUN0TPVcpj78
TAlDwUibfmagNXdPZgY9/Ac/CA5jndAsYpE/mLOS1cIVu/MsrekQ0R8/x+7MocY3/m15f7HyLpGZ
cZWsGTqOOI2n8c20Hv6exop1OBPtlb1iV2tcGslCFk8cVVS8Ci7wOx7xcShLlV4bmasEJgsaluER
t6lQZixNC0Jk4wEhfMIlTZzGcgP5a26ml/ARAsaY2UmhJ+kd8UtibMXzZEZcC2fDI11gcaGfNm24
zOitld3/POQDWOenTcftmT05vqoP/HOiyAyQtx1DV+urw8sUI+rx3OKkCpyzuhx7FhCtiUm1nFaK
jvMqoF7ik4KGhIZqB+HI7Pnpz68BLZIeoEnnktScO+vuacfcve5kzKGnUFMdAT4woaKul3SLoxoT
Duv8dOiVuu5sF7IdiUQAPOsqZleW6xbGKWR39JVTO9mqv+qer62WRXYtDDjQFjxJudtPstKDsMyP
cb38Hi9NUhqTeGm2AN4dzt7FvRbNGx0YALy5jLSVjzSxwdNbP24VFnt3GB7i9K3KOAgQtmULlWXC
/m02bh3P7AQV2aNWBQPM7bztq7P4jNyo60639bSs5ZccT6DqpVe6BP8H7VUHXauRNF0236/cD9a+
BhyGMjrqJX+oRqsF2sEKIopGiOCGip2zZqsF4IE8c2ZK5AzlHeatpmcUl5CVFS6Cwt6z+GzTUAkZ
JqaNzxtzVQCc4aX1OR7bueyQ3NAkYPDhfSOP52GRrYSMOgszvshuUqVi/awbCA43CX7GZXlq5H5F
HZFBvXtPygXuZ3Kjj+LxRqWUNmr5RMKVQkL68afmImf5myJ2xeIWdvrs6rr/lbfDKBKaosPjlOhD
6SL9rFYMACk52EiGdfdlTUtKnrNiiRPDFDZqq0iZOvV07PCiqYAgQEJ2/sYQzHCpe2fTNNo99BK3
PbVZdZLFSH/pE42cTgym3CzR2sv12Rwx4PcgoJS5ugNEdx5AhlH30nb1K5JqCnHiYzBsiFsv49bk
Rg88hqO1ZFhgKkwfIxqCiz0jFDtNakOD6UFr0mN69UvzdTG+UwWBQeUOGf8GUD970XQQvdaRkRO4
xeqTvLoYvBMchNj8JvGOFyZUsY9W648jATonDTaQIPvvEW/Pif+HtM+vkgRCxVcJOifHD9vqwNeu
zJEu9cl7qVuyLAKaYRPVEusLd8Jg81p3gKQBubnICdkkSY1IBQjKHVmAZiPrz0jE3pZQuAll+ZgE
WrYdGaMgApUtMPH1BpGCbV7e05NywNtuEnY4dpTxm0vB8dQ59pdpZYAdD2dvFWv8uPFpiC8YwM/W
QIWyHDLg8X5gDEMTcEiLqD8hyxgWK7q0aE/nUO5CkBcC0JgFItuXmSSPFj83xAOItj0Am2/VnLpR
8FDiLd7UB4uRzb4Y3w7VB1eLg96GRZk2nYTPtPnGbJRrIZKO4DPF2PaON+A/81YF9wJ3MENudf0j
kZSxsKK8b4bTDXLawTeA/O6+DnEmRd5/Qp4kmX4a7b8yxV0DdrzffpObxnQQVMgqg+1QgKzTsQjV
N6UV9lEJodHZWjr8c19JRwXYNtWtIe4Vr8psTt1Dms3WuuR9gvPbIaWIjzW8L1x+cUNrMjAS+NdG
E/Scb8BHp9lP7onwJps0GSzPnBLUnKPiUEKqrUIpwaxcNo1QIgN8BLL23vlGj8XyAJIERRkJuczI
eXQX59NeODgOGDRT6fQPC0TpSQd0OSwQqIVqRoZM9cuvcceb+PSJxMmnF/Mty6nev+ri/NsOmNjS
2sx89tFHMeyPikrPVYx/R8/fSFcF9vgoqvGfUPbE/vYAiOJ/wqL5DCWXVZ+fjQbgoQ9gbQaMlg0I
Cab5PC2se8gGA7OBZiHJ5ckR+6a1xvTxWF5HJJrewlBsaMMr0WfW0dOOJbUZZtbEwMujB8IYdjUM
fjhP53fJMsayVE9ajqZW2jRW2MBpR+omNNqUGa3Qf0x7tS5Cn3bkteiWqmRtCJUs+mSbUSAh9mmA
6aEexguomq9LuvYnXVIHlnUfZuPXXSFzCViLG9g0Z7xmHjxj3F5mg74FSh9enlhwC+/hamrK2itn
3bte7FupFsogxWKZjz7TuYJUm1eAYncMXYTvCI/1R55KyU7H4ajrRnVm1Y3KrADF8HIOqHkfImjB
rvDyXjZtvHv0ZCcDOzU29bLklXp+/LVJu5FTH3yRrS8NsDj6v36XE3hPQxNSnAHK6aZf3nnn5mHD
Cj0QDiJrvcZMz3Hi9/2+Mz0Z5hDM521NAo7DlZGcHipmgL++pem4gG5e2ZP46uZjz+K3h5Si8Hbt
TR/h07oq8Sp3P0wEjDURJUK5rYAAZ7xBDv8GCfz0CgQiAlb7+8NCo5jM4bxkHA8yqcPLuTqOek3u
A1l65TUiKbGdtizHW+WBqT/vFkEMI7c97ctrxiMczzXHeg6eUlvot1a4rg4MZXb9nc9xs1ELwdNO
nW8Uag1ytTIKZAkPYsGA0ozGRwPHsXJKaQOiIUKkvjN5pRu4wCGSA4+VCcZ5Oe0wYZMTD2Q4yIWc
4HucLj58Mf6B2JfX7flaMizmFyQIeWNex0S1IgOs6rM1zgF74AW6iyADBto0B+A7XbkHtAa1TM5V
kfleURs2q0cel0KAhrtpog8tvJbhcliJXH100QRhHzJHOMQySsxz6GgbQhpKZgX1hAIwh9pqYzB/
IHSYx88HgigMDzEZuuASsSTeVtysZaezmy+Nu246pNO27tbV9BlxKtBs/p605ohxET1iX4I+8MGH
6jrpAF3n2jIPuz1IGXKuvX8IyKRrMxYE/jxI7q2F0lueMK9GnLIEISqnJX5aynFm6shqMryhKOKW
8ePzIewQSkhArtuVPujWNvH7hLrYq00ilAsydC919QVTvlqkt99lsPG/eX9qF3bFY6GBK84BI6I9
1QKs9bqrkHCQqsnC/iHJn89vxAAby0wydjluYtb4DGqmvjwVMd6LLmqJXFG/FCKY6ZfXtovgTtI7
8G7TanF9i5JhSYss0hs0Pj6XGxNFK2fKdnp2n2JrPaJed+CmHX4aXVdHQOC2XkoF0KWzfVCzFPPz
bm2rWchT3D4jKYZmIPJcNhjZnDHYToI7j0AkfCZPbu7kdKA3pBvUSsPNl0frwfuwm978beKt6egi
OFb3QSANURaUgT15nV2TdPS94C/uHypZ3Mu+82FAIjsl6ogfzF1u0qdXdTsGyGswWKGlxuBKhNPF
NGaZuNQycHKbMuQbL5XDkt825HWLd4qepHdRDx/wgUjF1inPr54jka6lEAk6Wls0qjEByRI9UUb4
uWmVs4I4hLdFWxrXJsHoGzT+IA0ZSrdcjqpjyXzGFIjzLl69KuWZH1yj3w56zZ9CfqFz4ptXH6Is
nVXeFpdp/yUOczaU0/jY4jYP3E7cIddNDXhYqZgH27u+BQNWv9R0Ay8zFmBegtuYggHnM81KXN26
m34LdZsK1SuiFMiFOcAKtbjoEOH2f87Uffu4N3UJ8L+qpVPHHJceCrFnCsv3OW76vtZTAkTwIA1g
l11Qcl1H7cXEN7cIAm0ThfNgs5W66hRwIX2D5RrkJL12/kQExcnGVTI404aMIAOoq5E+eGXf01RF
yRd4Qjen1MDsKHG9pFPgyC/o7UOoTN8+emtqcI4BgasI9H170fifNQjsxR9oNtYpoXYjaqKN69yu
GfaWmrw8PyW2zMBEed7BFzCg3nbZLPwUS9om8yAZoocZfZs9P6/W+P7g2vsYy0B9lV3h5ShjkPgO
gghLO3b3UXanr/XOA2N5GIMn1ifR+FechhxoeILqzJwVkwaoyVtzIjnSLELYOGsAAsOV2N2EbZ6G
imqIdBo8Tghu1PaEYnT7CqFLXoVzQQW+mSpfIf6JAyP+ft08xfVeEaPf9FkzPI3UmJq8x0LeM2DP
6ksk1WgNoM78p1ATLYnX5o29axPg+plkoWtdfD6QSXfKoBumUn8r6tGzQtu95EyMkr5yVaCh29jb
/Xa8xKNmRT6ZpB1cciEUiHyePvbXDkyD6GG2P00CwWnVWFG1JRy1MgrY3Mm7O00xcZTDtfBc3xDg
4gOVDTHSvpjMh26ZjbuCzbLToyi5JlO9Es7qAaj6P8QT2Y7hY+9FFO1qSRPLSxDuAeGCPGT4aBde
80Fd8iCttg5zNC6s1haTAY9R2JT9jN/OdvF58Y/lXdfUygdEfDggYyUar7xar1ykK6a9YLOqXSXM
rz3LSyZrJ2OHqRydzMCx8ere3KCYDQv38NMJP6ltifQlfMLd3u4Gbp1WorJYHJW3cjFTE0EJpKcn
xay8e4SZaiCzQAgMFUThvIExpZWx90q1xJLrb/ySO4jFHB+/n08tMRnMacjCd8Y+w4ZY9YhUpQ8+
h69p1rzRuFtWY/UHBWJJbrS+eyZSUXq+TycxSNZC+Oj7oA18kJlapi7aBQn62LZ5+yJ2pcB7lUin
TlnfZ71SdAurWcoQAZb+7G0A3Ws/JuuZEY5QgmILKQ4pmqGQfCTlDY73lYNVKqcrr+8qWSuPHp/U
9fT+quhuB1LMVrev+ArcFnPrgH73iIFFk/g97L1MtwhkIxsv9SC70Vo7QlHYpXw4wZ/dYLcv308a
GG9hQaw6IZbyD0gtbyUPa363AN1QL/tZr156lJVEfdmx2v+UPWShtMqB17GRHILfOLTVKD91eseY
6h1lA5cnl+vJXgdPWPQxYl8C3ItGJbWkPfWCazcdZHgaH3LsYaBswKWSI4v88E+Dekd8B6HzZP90
QnI61X+wjr9Yk30M7KZjd8P3N9dBJOscze3juy7WzEwbCRr+C64VnSX1hhKlICnFwILELQUy5eNU
kkGeuwoDvzy2DQWsrfzHwY738nxaZsBNPYERB1UePdpHrh22nEUJ7s+yUrLuBR4WF9mHUEd+zWsj
SqDhJpIN5Uy2bx+ylQv3w3PZLqNVb39mzBbXjWsW9c6MVAeurSFJlWo+wtv9F5KDkAUTZC1cAVAj
fpWYjqjSTsSEcRkMZj4dY6P+oIeb1hHViSk7YNtXb7hF/mD5M5rFlJE9yhQSRqmco3o/rHdhHEQ6
8gU0Bx+wAsY2jpZEEAvCQsK1mH0i688N4ywJmeTn9akyR68Z65lwDnCt/GVtRlnDRSuB7VZFh4cg
PJBAOkuv9Hslz6wZQcbCwX+Np4ZrqNbcCvuRTvvWZ6hBQSdjERACWeRUnARgPDdn2QnXvV+cVnps
jXIbZz2ditBgmz6h2KEw+KkTe/UYQM+rxnQdDVQHEBYvAOsHIVB0Fp3Cx0YYfDlV7s6S8Ozent/0
MY+X8ER7+W6WS8OWjm8lVolRi2/YB///hu64ladm/vd9oLOXRTPeCbbQnt6BGI/g2KpHyE2KT754
sL4QIaOIJhTzIHsESaeUYyvBM/strY1b52i/otG5xXl+L4f5bBz7NmebbqEt/ldJGeNa8V1dafJe
EMrqZ/iLx3KVBh3rnvJquXhrI0TSvfzjdOYzs7vozJ46jb6P8ZK6VlduNHve8ffkW5I3obJwaHgo
FZEFNB6gb8c2oADFepQpDf6uRjMzSnGvcvXzjhgB5AorxmWm+5Pd7FIeC6lz3mszQZV8zKAnwXjn
dKl326i0dv8tEF4MuxL9Nt+a3Tgr6KkhOtJu5ccTHn4sZJZRa6T08b3X51mhQEox290AC53XnhUU
PrDnRDZl8CK2kF4QCbEQduSHlU30qu9gNOVH9o/S3TEkf9WW7W8Ou657oLGiJ1ioX2Ij0fFTCJfb
iTOF5fbDqFrDIbrWLRgYuPw4II5HRh6ddC1rTQ2lktGunewG/6Hpt3lXyZwvrOeWQf6NgTGeIXog
9KCZxUqU4OzuesuGySsO8Vy61AwI1If6FDJQDoSoC1JLmtIJyIVoKQrpRjQ4RXZfV+Gr6u9nE+7P
M08hBvqYs71SFS/3hATQ41hafas3NfcoHBaQYsIB5MaYyfPoxKw5ccf88CkPE7MUbLjVl9FmgK84
Nx3u7G8RrO3mIb8uh8+jVPPFAsLVf4h8ZJSPKoabLtz91HZHDTkj6WTBwhUNJFwuM0+RJmpWOF7A
1UMcivfaLvsU5NGFQBG95JriAgUpxfscu9qoCWk5TtNhvYBE36ASBK7HCmnNyd3jzQ0e5bOfeZ+w
5vT8BUCsPN1t/CsDBfff/v8J/YjoZo1UaOAvmEnv9deZPi7cqOlVpb6aQrTbGP/ZG1OibAG9CEyJ
w9I2SvY1aZ0015S0GrperzWDK4RdkhRFkFWW9XwY2n0vwRUy7YVN1BGkiJ/UymiufPXIeTW9JMJt
AAl70QMSw2nFAEqlUy+UrSofwWC5LC1b3G1DU7CAWsjccuCYvS8Jdyxjcm70bfI9PQvExZUs8BA0
Bnfy7/+WmkHup42ZEBAn9BGBL6FVbXxSHrRGtpJaCFo8c6secBceiTeQuUg2uF9su7sCDPgeJCQi
mNZUX649mkZcJrE/dn9HpEH57YwyI8RFXOAvc/okGY96UzlX5TVjPL2BVSvaWwwLiwime5gNIkex
jo4neE1RjZaXBLVlmu2dPnsdXgDND9IiaO3Qj41deGMf++oqqd2bs4mFrzz9Q6Cp6S/Kj3TqmCyw
pLqh4YON7DwFF82B2JaxyUS7YLnaUWu+KDYVEdH+X9NNQu/UNJFkxHvVB1snteDpuVFsJamybNn9
XEDvlQSBOLSSBwCJSXbRvdRM2dGs0zyhufV1XuJ5GrEWP3LNPZnxeh45xCMMdt9IC+zddyOYf0ga
hlO/0rsiJee5b75e4lC9eN/75qCsd0H0ecYv52nEOiF1+60PcDz26XOEikYRJ1Ly0oGjHk8JAJRA
it+3qGLitlVJ1zFxm3OpXoP9Gja/RXXYntrLcsBJsicy8wqFFkf1bIcpv5cr0NSDdFoEhqJ546HR
W/XhxJJHBL2RuhLOcjNOeJpCUVkUwnQQtbGu97ZApCBbsjQet4glcfmoEhsDRfwhBnvb9tRNOGHd
K+0XAxz6UFSIRIQhtoDCcPEik/tTGX3nsAXoHgTEoJ6bii/Bjo6syWuKTTwj4aAKhq3aOzah9eyq
bAYMI+UBn3hqJMVxVA7xZhk5y/+YI13BK22rIz2ADZP0ZxYTookiT0yczlnvVKnCgYCLp3wzkP0G
Jvwd1T0HvzFZrVauwG0AMM1AI/dyI4iOOC0PnjSj/nV1mB9Itl2LKdtxrzm9BAlhwt9zEAJkIGVI
EcT5PLmyO29PlRMuVOJg+dlc/ng0xDpyN2GdRF2gEsF0w9/DhKEGzXTh4FfVolVkH4rRmI46QG1q
J1qSyqP/8aP1yO1FdVyRkRWsTz1w7ofGzgU8n8SZhpfzxny5VWLmYUknRYDhT4+GE7o2jwiIrwu/
C5+snI+3KlOa44hcpPAPcL8qmZhuNylXyfkEs+bEXJ0zCtbvOscDMT2TXH1J33bk0cK3X7nu/PXW
vgwes1ImdGOzc9lYT899Mf467EVd0snBmhnFqA3NM2Ir5dCLQWd1VLjt7CChKJLn2ZFz9WCUuOZb
Qx3l1172zfs+I/n9d29HgieenoLalNUVrcgQ/raMMkOb0wIzzTIoh2HVmHa4QDZ9Co3QRumrsiko
LKweQPNnsFWdNo0rsQikoeG5kEaBEtw5aQ78274xVR4xkmw+/zvOOI0bew1oIQxeSzphCUB6HpmG
LGR+sHnvkqDZXCdKyBXRhugGAPgiuDEm63F/hBg1f1SgpETSw+vqnGnMicfuhdM+EBaD2HdS4pTL
3Mq0DKOUvuAu/l+mQuXp7klHW3hi0+3enluOMX2OUdRNIjBSX6c+X91vDDRNdFieGh/it92l3Aej
T9nEnaNGWVnpq4akSI3nYrVXKA/FvrOgtVVU6lpcB4DB+fZiRP0Soijg7N+l4T0YzmPVxfkTntry
J61wUDsX7WvJ2R0hF+/Lg4ooGIkpL1ZZmFRFipFNlg0HZV2qT98EXW+qxrBEYCo0dET0oHZlYLeS
v3ATmEpaCQydorPSehOzIf/oETRME8Sni93LLfMboBU3JqBeq/cFbLW+QGbQkIBl1/tvOa1Xxl9v
HadVdOUitH6qYG7yRhvm6nwuFa+EbdTLKyp6itHxXj6bt95MVusLvMb5Cmuw8EVniRkEaBkhzCgi
/CptE6X0J/r6xVdgLCOcWpePwiYB0JUJgJuyizZuei8eNlenkOrIk7ZwR5dRYPQ5JBWMFzxz2i/l
7PJeJZ4LAC4O/+zqyqBfJ1Wp8GsE6kWPUXrm5Avl9efQoeCqx2m1ppHy4Ki7Z3pkXklJ+C/Tjo80
rBed5KrVchQNfJZOnVRjNVexXpzozkW+rjHCoKEuW6Hown7spfIrTNQLtEwrWBKnGBs/dS4zIvaS
HPRXlwopb+tjJl25dFzUwlgOOw7F1Mud43iDtQF9cybESfxnIEIwtxhPbExyBAqsldOPWbQuW/mT
Z4bx720mGCK7jeu3ftXOOqRbnFvHNBmXOLfEBWtinfZc+570Vt3bXYHWMiJVVqQ6iCz3PSUHp28Y
KhH8HdaVdIgJDCiodJGi0bqfcC7Xgfw17QYQWvGqsSdkE86TmJABiaGza6WveUQIY7AfmdHR2SK9
jlhEzOWD9gcWuB7OH9n2DBFxFgyEAW/8STiSPUJ5KKsWphSuAN8K+lhf6fl1UPkL3hSD+LKezKCc
bYMJeJ3+mwZ8PaGdABoeJdVBMdp6TeNy4m3EKA/tmv51taxgJPqkAdrIbWp8XNBd2E2LUBS9IknZ
lMIH9Uo1IeBy7Dha+66nEV2WbLIgwfYIypr/5IVe1LJaqdjqf6rlwrV/PsXtMNDFTwBnx/7LQL9K
fZh3GSMv7YM6wmluToqG7hCWcMHq7WzX5yRWR2gTqeAn/P4rVdNMaVNSazESqWKRRqFckWDLkONO
RbXJrafd7kH5Q/gMuLACMdgFTsVsQPM+vs3Wc0e57YHrwQQ5hdDvEIkTYArHeid15vayKy3diT7G
uHKkgGHocflFJLn/9m0zQ04TRkGfGXcjxPVszIkUVn6H7iWJjdEeZFTFGBMtDIj5TD/DGNsAUELt
e2X5bLxXr5a0FMJnSPkr9H854tMbIJW46Jc78VcOXnpgRTAlWdGk0GgXLjR2XcU/eDBKeJM7zwmG
aehdIpmx1zhS27ztZGV7+GGXk28G0TR79tU96FowRE2r6EqzLirBn2SSK4PPt9rAK4CXQFV9N3nW
ViV7W71PceLGT8mCFWIAbgW5eBJlezrsW3fVBKNcTktUg1KOZV2ERdqyVGrA2S/LJXXzEPMhAg11
TZabIXeK2jOM5p9M4dk9G8IkDhSB7hXXgs97k8Y1Plq63EoeSdSZvVa1+NuOlqDe5G5MSQRPn6Sh
prDtSOUyy6ktjac739HG+C7x6BqpP/7MeZLh60pFgqxPXiHB+azzgcXV9NAEyspSIjPzKxdFI6/m
C5Rp13GbQiNIJZ8iKB2phhiPfue990qD6raTujU7N4rILFD+9ZSrteLle/z/lK3YHn8bttQn0w3+
1542LvXrAH/jlR/trZyTOoP+5l2K0Je+OIej1GBf98MIWeYq6JJea26CYDmWZQjRPEGgH4NJnzss
PL8qUryOIJ1n/2pf+a9lp9uOIKA3LsBr/s02K9wjQgEJDRTNiWeTGZRLerzWjCa/9SbAUIZdNt8X
zf9S14BIEnM3nf5LPCelgC2XVNPOshWHDuHyI4aRytpJNHBkA8xvTRysbYEgXRzOXXpXu07vH0OZ
F33gVDCfVDlTjDR5OFO4flbm018vnOpn57DEePx31Ei8OgnPrqCvHbbintFIsPJMFchbAX/vUdgc
QMgQPibjOsBRmkF6kwZRl19O5kzwHqo3c08nDZ1T7nZEh+n1sxx4vcfyqbERwdLzYpO9n1ZtrEMf
HIHT1aLjfFz7xTImMbNmQ8muSM1fCibSkEP7NJDubnvoCtHSWn2K8Jm/7t/qMFIUknnsf0S9zQuP
/xAW7oa0bTTXJVGflCQZl5Rc1kNFIXIItJ6zfMrPCygdKArz1cE4a+UkDt+BNzR0H4VZ6PH+sh/y
Eqo0S/jK2rczS7A4JyRcOiVt/tuZ16e3ffmTKpiLMumKCarKZitLDaO/Kr6WSBOReqc5nsfPYXcc
bk01Wxt0Q+6n+YNCKMnegF88Khl+Dsy2YQ1+H5OdC+HlmgZOcDEJipkWRxeqzV6tCJeC/v0W774G
tsuZ5avG4GQ5cQOs29A61EGsP6XdOUX0rOKAn1IZwAd9kidXUenVO3gWriDGgra404ZQxKGhk/hX
5KEQDVX0XseWstChoAVaJlaX8rEL16YhuLrCUnWOt5LYfzu6WHhy6XfRILx3PQLk6NZO6fC5J4G0
ZxSOWYm1Lr9va6ounQ+JQ3/otQ66B6wGVEouR1LK/x4O3sI79L2gMwiFtPlPsktdYQtur9QlGj5a
VDlhqq0ej77D5b3BQvU+HpXwsVVyJho9nMK1bEBrHvmsH48sjqByJX7KU98WiR9xfRFkFbBigrDL
yeK+aZl2GyY+vNR1/p2lQWjzFjfQjc7EJKjz6Rtw4M4OVLPi/92EC2/v24aHBkh6T5FxJJ4G7HP1
Wt2VjuH72ucdtz60GFvXgppPIPhrnVk58e9JX0YPFZR+wUPo/xlLzzHnR0d8MV/intK40hXA6Gvj
8K8QBR8m1I1kddN9JSdKJLG9NvWGNsrQ2ReBqcrwJPIctN3cqQbIg+1Dolc/yeG3DXJ9h3F4B7+a
Nj6KEgWi2PldWaYrw3IUlH3Kgy9/SWTLZxYQO2UdW1VjS4VXzZ8odskZtjD+u/cBXsccAkGCRmNl
0/kC6MmiZMLL/GD95fCrh4xWBcX71Ut/iO//C/Qlqj5aU0skjAUMIn5DFXV9DpQOWx7P1wi6YsAS
e30o0AT7JUzID+Pk8Ol7CWmtc9w7Ks/qXFei6uA7qLPMEeDYK4/bXhqdXM09lTOqqmyhUspE3qE9
fwhQC/OMnarN1jia3zvrDaeSfOgksXXnAaaOB2/XhSq4GPe2n6hHm94FDhaZIhUStFfQav7ZVOJt
VkgGzwNiN+nrCYnVUxlRe9GP83ygipBLKZATLQUW94QldbFUSVPukzHLTEOeoUW6g2sLC7z8jVEy
SZ8AZ4jItVnkwG5YNYJwLBrU1d25Dw8sGa/GAIvbm5Vum/EIcRqNOMm0NRPKRTtSk4nLB6kSY+Yr
51bWhI/AZmf8cO0Ii9ZFm/ycA0trqCPgu/IT5Bc24wSzMkqOxGbj3jiK0VaE6SbNl/3svuUWRdsI
0TjrEKX/apbc+u/livJ7yv7Kgm6ARxms1UqVtOc9MQtcEAWHJiTaurnA+CGEMtdMtpD62E9xAkp0
NAkTmiKY0Gvb8FeBWvaNOvHbQJpAkoI5BKgF5NEs3rwxE+6+XQphlwxnPoOfCaxTevf7Jk9adM9h
6MCFcwBMdJx6GpKnjEAzQI5O2oWLwsehq4hEWjpS6qcYKqCWv5t5FtHS+fZyVdj7ZbqGGnMd/OUy
YZ6kzWF86zqcL7NDXphASijJBbTlN3XuEf7VqS20acni7PBHRXwyFwAwGen7M+E/bD2t8W6qqfzm
vLR9TliSmNvKJCl+jzSIXYS4KLY8MKW03A13SU0ZotASY8sTmQFIzqwwtQU7Grs33iPTj7hhjfp1
rEnSFSQW3ysHfNQy4pcgIj5XO5J2gbAFawh6+gpF2PHnz0CBwDptpRAejzSse3EGpZXHXF2QEtu3
C5zvp5rGJHSDxXhsahcZ2+IsdmuWkC9f2/8EIJe4JZr0H96MRhyiz4hD8g8wt1/IKDZAI/tmUXg1
YYY4+gbqghbsHLp8VN+b6PW87rPeN/Oj1eE4k0EKI6rt+W7ldVVAf0YmVPkSikPfOK953Wnyl2Gx
HY5YYlQaUfwM+sa3xw6/Fm1/EU8HKxjg+SQaWUVpE96wjjwIKtpHpWicBApuRDA/Hh7wy3lPXwQy
n2mliB2B4Xt+8jpB/GzwK5S3wccGnHs/1OUxa9wOSho2XzW+9QGwtdvbMAQFWn5mzw4eW3HGhzRz
E+N7LfaQCuDj1x3MfaVBsamQRfAYAFfSS8RTpax/m3VSdXcdiUW9RfZWpKAymCwx0VN+k88HS/sQ
vGFCfZkwCvHlwEpLmgIv+BssJuje4tMbNVhx8UB4O/mLJt0w3N+B+Z+LKi/KuCA0Yd8B0FvCaHov
pS+njg6QsoEsg5ozLlln8LxNcSNtWZ37DIQTfjEXsuXvki1uiZ1fTVA2zs2gqp6rLwdrParWs3Hb
Yzm+uxTBbYCBEZvCDT4offtSv/66OvMxfEkY0tirqSfdi9cOTjFlbvrjl8VgNOs3mkhaiK7nEirU
GWgn0zt/0WnP8kHoiNEmDzBx9Fvo6PCi1YNgu3kUBIzTQJWZ3Gxmg73M5b1t2QxdPIfNjpbRwLja
vc4467lLAb60aFQO8XkYE41Q2P/1+MlJH3MUGv31ghDQzna+qod8CAC39slItyZ1Oqc1gX7MLASq
wPEkX84BWyyFt0aIyYiJovgre1OjSf2JrJu8nKT6k//sVdsEBQqt8qaOWGCcbKdwGEIdUND/EO0U
Ls4BqHVtF9UiIjnNxaFqyf9aGmB0DMfxWKDxlfLp1r8Iz/HULz7dxr8rxJLnvZ74nPOmBuhBIY4H
04NP/15BMxU2msXQYEALbEK6oZmVELovT7GmY5qEYnxz3OttAsOCJfQoTb1BbLwjjZtSHJPQ1RQe
Hndbwxw3oTrl1jq5BmfEb0DmlJP8ISFDbWzEeK8YJoJBKcstibN77heIIAakPmuBPdGeV9QKJwiM
awmbigdoqyaQrAgPLTvC/BYDWF9L16ZcSsLXYekvVGLrwKHlcT7Xx1aQgVOSyud2ahauDkf+VXzz
6qPseTUN/AUihltC1f5MRnl/GAd2YlQ0WQNjUM4pZG4y7cITcQuuIJv0u4ejfiw66kqoI7g5/DIJ
GuTTXE+e8hvta03VjNf/A+8G17JELJvIBpRjaEsQ7w4xYcHBUNyr8GSltYwshmPQj+Vuxm3JoXmo
2/eiXRpLxzL4cicVvHL+iVeFI3ARzqdnnWG9adcJyBeN7fzxKnKSRD3k4iq2OTKfvNWZzmLpgLiu
B1PZDe3ebbDPxbsJ5YGfSR88A/xkbna82H62hiR4diyCgLkSvMbx1sZPuqKKa1BtnHNxXSkyCoLX
DjFNHtrR+deOGY7w+VUnGzt5wVATZ/+/DmjXNHX6yocmUG8jsJxMiJ7jkBxwtlBIKaXJ8q4Yrlfx
P7bYT5j+nUSpoiHUkqbEI5TWrmlipFnKsMtJRpuqblbkaYYQck1JOGmqLwAUHeQcPIieRpCe4Cpe
mSya48/lEIUTJLef/4lbr3UmIfZ4UaSgJxJif7LPVG7iZUJcLKECTRQezAyHT8K+QxhLltuqwBLB
Fu1e7T1V1RqJ7niqeD6F5goKmVmZljAMOwvIs7jBGlmgibbfLPiC7oeSt6NSE1QaAX6MC/OKVi92
0kBlPhcUqAs4qvkt2QrALDki7kT0oMPbh8B+TGo9anKT0dZCy4kurr4/k2uKqGUw6GKhhO/Fd8SC
l5zDHeN/eM5CSAHu7aWrCERMGc+dVAtmc/k4+2PzNv6Waz/sOIqmzB+k58hIJZYjzCZUZMR7eRej
4XZQx/8aCcOpUs3TffmokdPslw5AffIyZO6dUp3ZAQeP7YElaIPT7A6XjSvFAE4Ow6WPLMb0dMsL
kThWgJGl9NknbG5m0Oft9U9kyZa5+PfC8drz0+bAQ+oXD4eIX3gFsbonmCPp87ue3k/Afa4Plpor
BDSoNBmky2LaIv8RfjAdlEDvQehuTNcVretiNB/lrk7MPU2PflIYj9NZY96ks2iD8vjeKuhvmRR+
RaUa8cAdkn1yT/oMY34mYrWtAr4kBBLsqmT9Z742D3OKSWA7ZmN0s2RtdfuGsOHvgT6QvjaqOkl9
DbSVl2yBoP1S72cgdUanU2BtNcDnBdwsCSTU5il1/ORh2Qu+klgYupiVwLSD0KA+BKH3SVA6pGT7
nD1z2slM5BlfoSyNR/mk8An3LPJiGukRzL1HKvoRd+2d73PkAcypnYesNitkBW3PflVC+6zS48Zw
GgNtvzN6q1Dkd9wSGLfLM8RmxAp6zZZXGzWuhenmDRzbrI05jZ4KfTjBZXiN36TvP7rwVWssK2ao
jj2CzKhIdE9rQwgcea2m5+QiY6xw8CVMb3yIM/kdJDjSvJ6ySj/WVf8ZjHxX9jNHn4Pd0vtumuGZ
f4hFo5EStzYJEz6ighOvtBHY6wj5kQDyPpcUSDFvFUjMymVEQJNHp2goAuZUt2I38988RUI4Ypz4
K2iVvnbAiW6rRLpyftddiIPuuWZHiqHdoFf+fuuCTRQqApJLt9R8H4yFDmzRqnEIDr22Y9EgEDwQ
K0U4iMpWNc73vjFJ1IMzLBXjsLXiGSMBpy/NRq8DofKqaTlOFahcJdh9UCG/PA2C/VuVlOeH1Fzv
GVo/Gl3xHEkCLjbe+R3GcnEEOBeVRvYtpTibkS1/ZCP7ha+zyTCEH9rxwdd1q8RoL+H34QHZujg4
iflxvajXaNVaGd+ai9pDHYZ+5DzUwPTdqVBueL/9F5IiUyv9pbxcfTPPl/z2Ar7h8pbUKOHPlM1c
2gjDuu0u3FkTv7BiW06l+eI8k/b4PeZ29NeYiI5iBJsEb6Yryplk7/3BxMVqh7cRuvybVPQpMkwV
AvPP0YyPsTHue8/8FeWvDltL9gqix/7Ap40CUSitIQ2cYEJH+XzuhaOqJp/eOZnr+JbKI/Gaq7XO
G8aH1eb7/UUDJ1xhGaZjQabAKXoxOb+jSBkEpJ5RUfqKs52EuNPrE6AA0l6/SFsCoE2n+NFrXRTv
tmo3+ddb7K6bb6md5zp4/QP2Sbb8MyBTNA8+WVFM7ebJyz9C3phlvNtbHUhKyJAPx6bXdOXaoypD
cIr0AHir35Wp85mGDtMG8duRd1+5CRX4WfBrZpFMqJb1B4Z+ULNEBBqP43Uv8PZYDJGP9rshdGBW
Tx/rDgqdShpdCtwMxIC/A+N2w0MVqjjbHlwK6pRhdFaVoZkpMYn0BbxXS7vhqOWS5FN5qZjJLqeT
YhN3oJbJ8CRhmWwvLDkDi4QZNpgEXNU23CyEHMo8LvVgPxcjaMG6p/6wBJ9Vp8be3Gxze0IiokMJ
Agp9eH+mWOXNs5iBFijJ+UVhtvIZqLsxwrQVWEFwHRESQ0GvFF6GZQLDjm6zykCMNYaLum1lqpqf
sCF+MSOjroxLNWmV8h+hL+1Ae0qVhc3lTbv5ZlFrRhh8hft2+mO5Vwo6MlaZeGIx41YUAapTFLRq
GQ15CtuIzdd/pAbMIT+Z3PPnay6MsQNULJvzDf2AvToNmrndbccxzO3LGMXFEQAgdIadlLtkjFB8
i6vNuEh4DopMgH7b7lzFPSLc81HMJTAi8jERHSqMIoK7tW1MKCSEO9V+RaGkhg8q5ngH06BJ/3Op
We9LLSvFRqo0pZGL7KjAbj2I8IwXepAddtl+SMiFUTFG9DmvqqZK0TQ4W4llJF01bLeN70iVTTC8
0tGnsnzBqiDys5oD66gvtxLPTCaAafetJaEg7KphHsokG5+WjTqxad/L7xXoZIfZrCBWn2sJsPwv
lGhwWra2rSwtRhlsTQl2wqVnbpVdYmTTLGpcJjRumIIcJf/Y8LnJ9dGpJmLd0Lo8hpIOSjRXS7yl
b+HRDkoxFUfWThkIUU4oLsXiGu7CRKmQ1frkxPin8TKXX/tDM3SFv0rTiArPKZuSsjIrGGSIWZdO
W4bGsImqh1YVHVs4EGv/5I+ryYF5igfBL4bOtKSwmteJlwpgwoqXpcg4plAqZAQor6aPMLWuVv1U
Q4P61BoOBVbZbZMafn4pwHzvCL8BMVYuwjiM1msiXmCbAFwfxR/qFFVmswUVOqTuv0WiOEAor7S1
BWUz7p8A5xKW4GmwDra69CDIu7W9J3l3nVYNh4FzGPdUMc7fFuDRqF7mSN/VATskGHs3eAMj3SmX
Fz6htL5m+zg2NER8hThLjodr0dcJYyFkKNvwK4vJiprxGnmKTlYU9W/xB70ZDAggofrLGnJ3NLnf
Q0Ca4phPs6HX2bd9lqP76k5VNPXAr5kwL02gdjhNYqY2T/LmTuT3icOqS2v+wPAGn2MS2PdKXK9a
dDUuOB8AzJcY7ThNTQN5VkJztFI18+l7ch4ZloMwjneREImHtTL9GlIcPUPY4qRp5DRhjKFH513g
AzGFl+isVYQQJLU38OKJb74IZUfRbB/G008bSQhlIHWzhX9V3AZtL1/oyYTx2sTJxTPXNlVbzIUr
vT5SzS6JwDBjT7cq1mgJbfyKsu/9grbj1UIwaQR+zA5Ufw8QiufSAbsulfi2ULrYYMEzLfwfjzOk
kJNOqpmPvNT1j0y9V1X5gIBxBqTMXKY1D/fb9o/byFxwhl+nf6yUzECsXYc9s7FrE+Kh3hX0QrB0
Ckk1RkCDf8g9PWoDFU3pFMWWaAPKGhYfgp0MMv0vRRRDoD8o05XD48PeAh5cdxZ+UwBLPO6KqDur
pwfZn+L+Y6AtUMKhRaZSM2TOqiziQNZ6ZMiUo1zth7dJ1n9znIVIuoslWeHX6zRB3pVQ0KNjzkTZ
LhaajqKb6IpAUogAJ48tt2j7iJlhfHc9QUPdmuq6VeUmoxddNmWm0V9bibOCGGHvzpRzxQS9uKla
NqSjmATuEJhtwXu95IViIDiJHHWE0sVCfiglF3QDA48ON/Y71XzG9RjydKRkXyeVeAXLhGJJjL7H
6rWJkd7M8IlhLrf+IZTNHXlDIxFjRFfspPZze+Gw/UqTp8JEDueu7a+qGbZ5XC+uPxUVsPPXappT
j/Bf8gChNzebAzRNS2xJAsRjT1+BByM1aUbXmT1N80mgBOC80CJZ56LxFADHwhgaFMFOWtN+svFD
2NeC8bNM5qeqfjkwUVP3Ra0xwZJE1ggp9GNBrkpzjw/C6nqJSlIwrY4OMtsP9+TZvK8sSz2xM7bV
OTZO9q/qUGl0ZJEN7F7Ougm+PzJ///hG8Z8Q6KQMVps11C3V+G7qEppP8aHs3lzkP3j1j8J7HnMs
pw1Jodj5kyGtfKM7AAHFgrJHI18N1WlR5UEQvuAsXtE/6spbKVm/L2kttOVe6jynsCUYQ4Utwuwk
ixsEow8K8Ohogt1zHg0l5vyHmc/AXJrgk2JgLWR+FlIuF27MYADHLMrLPA1dSyxNQBd9JBvqVi93
CFt2StG+nkceymeJtXAa/xCiCZmV4CB2rFnG4GYcFCYs41mu64mjlrC5gUe15O2ZrN73rzOeNIZq
VjVapZBc1hvOFWv+27TUmPIyb29GFix1+jlqAgSV5LgPmeDGJ4/s4Qqds8FItv2NZfIJOQjS3k3K
NyzLAfSaT4hOx3qdxFwQFz+YTnQQKvo+LwBMD//Ce0wk1t+gVQYXAmeWE+0Ca6YyraeC2vVftAt6
8OiwUxBYV2ONwc1idQFcY0E85uXqu+X8wC/OV9LwMr0vQKMTzuUiFaHMpMWkcgdvH+J//zt0H3M4
lnTzPf/Dl9EKDlUGE4Ks3lm+o+yBb0Wh3TQQxSX3SOAirkL1ZsqS/1CO2HA87Jd7bInFv+W/OJtf
YlwHM9N6RocKE6SWSM9Fk0oRqUvY4Q0tREG5wgdspEaFqLBrIIHQRuC8runyKdylZBgi05NwVQo7
8lfLjZOqPvBrg40lPP2op/DaMIO8uliWHJsUDbjO6UgJc2KJP9/Ex8UdcnIVLkXkTVgOIYCslnCw
KC8lDdmMCvwZnz+UgitETCgo0vZBo4cOoyoIG0Eb64ndK2kzuZkTWteJ+J12LWtSg1vUb1kbJOGx
SJuIQtgDY6FI3T3wnbSuulOY2if+85Qfm/geIg7rUE/eSG6IOPrp1CVuMVOhcNiImiig24WmWZ9c
Hc1/O6hdEgn2hCnBxQOVxQn08ClzIy+Qq+c0ByPjQ8lYJ7jXGfR48ojumR6YVLSZRqDrwXBtJ711
/Fr/AP3OAWlCmzjc5oMOl5lJ2OMya161Ddgss8f83QdGs0+dqjuCOrTdf8Bd5FHf3/mdll5ow+FI
1nuqKquncQQR39rKWNsmw0LTy5fieKouYFSmFCvlAuXNwGbaL9yZnXXyz1XxZlnY+An93qautJ78
5QtyVY+bG7pOhSG3Ia3IGX/wsKlmGF4nfm7R2u3hUn14GLJ4FB029cT8Gg3P5nbQXUJCsnYtFMRy
D6eSSCkMzDxxvS9MJNum5plmCYF9qBheliOeoptYYuUZuFgrQPUHVyR4g+cM8xsFgn+161afzPeH
hGHBnzhwHaLK5gHtAEsM34PWmKip/RVDx9VZUnmSSa4cl8wJoayK8jJ57wCOtubiBu+w7p9+NJnb
hrDJE9hy4lGa89n+TP0WeNvrJPdav5IUaRWTcBu/kMjPARZpOy04g6XSFkKKr975kwE3MJktsewu
o6Qkc2orjfDYLE4Y5rSdqPg2NhEWd7fm7/NVdZB6Utl43Bt1FYeejkJHcOhwMaFW5oo8LSad1wik
6qWiErh+1ZgTsLdXKiKFRVZlamURzIPy8ErlIq475qx2qX2vxD+TTCcvnBHJ8KGG5oxlVhovlMpg
L7r3/bakpv567i72k+LtO4DocNt0g/MOYdGQWlP/um/HrXEiDM3V4FdLTsO3RN4TAk7xxjFXsVVT
DBhfnZNlGC9f6qWpIQEgRTgQmLaI0lBt025Wy4sNY32SrVPvNvr6+UY1d5c85ck64EHlWOBUHaFW
8TMK2pOzCU5YRXbSUqaw6/2Wf2FNMoDHQpfCQliyGvOmBKxx0YU2fhI2hQV63Zjj4pJQmhi+BYrm
nWa0hkezpNqSXmHcVcHxw4VF58hSqzBYurBy4Sz0srCTzs7UDwUS8zgfvlbyXlaBqjmdMfXTeXkD
YXkfhAANXi+dXziU3zQtdhBWd7ABSQfiqzV6URZ65wx+juT47z0TnDJFHJJEcrw1cuMl+4NSGs8F
UjCwl8FkYNZyAA4T01xVgJDgNwoztzTErRLtBBSyL2I+AjwsyJHYN5FHFAGJcNFaXpR9cjPldMC/
X0xZ5nJ1bO4+1Woj/YYv4Ec6oKQOk1Lw7w+24JWqpxl/dqn8QqHFZ/sb6YXcuPGGW/jz5Lg5MWd2
txc4Vu8Z4N9mE31RaORbv8zGlCJnPYGxvrPR+OwArokz5kt+5ZWA2WasY+PYZTiJPXBe+ixLYZjz
zzCr7bKHotTRSszWm4Ub3aWy553Xxl6+/rtS0xBFrQEUi5yQUrIt4D5fZi8Y2TNQNpavjC72Ckex
KSTalErkNEF4WU70GqUZdhFWtQlEZHlHDeUbAjEWHJ/HF4ys1JHGVJeSr0NIzGrWK2xO4hvyE0jn
PGplPve7aWf3dYiUVTe3wBM7WCAWY0RPE2PiDdn8VosFCtRCPwQc9bcvSBybtutEPFPMy8sWGcgi
s3mE8chesJjan5okhjhEdJCfOl4038OobXYqUjCtv6nq4/2IkyZsKGjeKI1YgKU5q5M/9NjFLHsE
AoCHkgNIJ7POf42TugdQuAoz0e7q0mC8/oBhJViIBBa0XKGyqdaM18jK/HeHgQTCJYeLE/zB0MgF
/fEdMHm0qEgHWe1FlJX1wt4fb2Sxb5bPbuD1rdsxqTstsJSU9nhDLWlxJI1OpPKHIE5MIoT164Z4
Lwp+vwU02Gjo4m7JTVfRWwXlUTDv27VVs03sNPodGrWAWh5tkwgCPG9I/9Hww/+y+V31/4a6/IpH
Iyj6wNZI49S9BlKczWcfHpv3+9UAmcVOJpr+wxub0S38c2JHVhxlZMqXGgiICAHXhakOX/PHOqzI
bElp8vjd1SW1SD72yp8hDPv2akea1k6PeEJgCA9ADjRGGjatqdfVZ3t2FVIPCJBTKMtz2H7sKsGg
y63kVmjNfFh3R0PKqJnstUV/ldZdNaTE0NM1p0UiDzX6qiFmhmcpiCxqIcgDPm2rd/Xb1EpDvBOW
jGyZ37C2RkYRhmsLcCjCH5+fY3itNVVwhDb8j8CFq1Gbv0aJ4ndALvj0pF5Uz/Fo0RHjmMBE94NP
Od3zmlOzOkITi8nzhopOzx4JQ5lPMR+L0kshAMCjl9CbZufdn5q8jMW8kkR/IDDxz7UAIWET8K9u
HzY/wC9tJrJw+u3P/H2gV8WKsNWkL4E/V5EyPTpK/g/rN2APt/x9LfNdzCNGZqmkJXWylWf33ch1
y1LlF2mFPdhEnWjePmUmDYNI9vZPPjxDxrX5lkz5scrVYO4v8tQw6uyb6B+4chQMxVmdgrEqgPpg
YyJe1BJ4DvkTfxjVPyo4nDXepqE0jgahkp8GOdjv4T1OWB7hbLlOn2dSW+Ffk6dyeiEzOCK7aJ5C
EqXj7Ne3tG0QKHEttUy8+h57KE0IxVo6LMM39P0TNSbRzAqvF8Ux9I3SlrmtLJYg3D8IRuucU6UP
KXHS7TqveTRygSkL8t+hIoIQ80LtgRorPSDWMbpF1Nm288RNYFQGKxTzfzsHjq6MzrCoPJtU8RHa
Nc0wTsmf0MME4PBb5aFevsktCChR+FNJvwT993O9Ta53W4PgYXYoO1lLcY3tCDp2Wi6KBQ4ZjSS9
RdozcuQtJ20//LwXRCpQo39gnZKHrPzZaYcjNrvFcYvpzLu0oXtYqsZtB3RC5D5h/0mn+7oNkQWY
lpjzVxHTRoyBkKnn2SWTbP8+0H4oGw97Z1vGVhOn2HUvElEeSeOYIdq26McIuWz4ZzchfNoB0Y4a
ww4m3Kg34JYgiZ78bmPUZ0jXtijK7Lt2MqXdfz1YoxiUSQEQ1YMZkOaJTRf+X1Q2LGPek2PUzKge
DWsiezAm8+BUgGxGumwXnUZT9UUHQCxPIIpvT4rXV1r8MQffvPYTXBOr37z859sJm721CXb6/XBi
5HXMd7MqoaC8y0AE1Bk72rgnnnmiPKIMu3i2h0fsyPEvgtg1Iht7ZhZYqo+bKlvZEN2T4cOk9FJQ
l+1leMcT3OQxFYJJCzm4jIGVvX6u3dv1m5v3tE3EMfzgsPmmxnFBYTNBZNiSQgNItqKHJlGbhuZc
oScF/msaYGM6TGm9ZzHR3ac2tP+oXgubbF1/fjpShk6Uu0yvjLvzNliXfLsaeB11iU4gBQxmTTsW
ThKqFUt4W8ArJxb/KchG2f7Z8J9rEzQ3k0z3pYgW3oHRZNLkwrYvsKZbGlI5V2GKi8s1ARmWkIcC
ocvdSTeV2fkI1h4EULXBM3/XXGCWiSNoljepUfW7qsg7Btd5u1FluF6ploTG00vf9XfkfZvkmOgO
uSnYjXYeHix8ZopHJUtsNdDV5SHrdIyxlI+R2y9A+6gcn9GaFj1KJ2aXF3zhT4QECo5GWE7rXEpI
ZxaSrebEFBR4XBPtRkZbV9u2dQzjIbEm4fuPus2FTGhdKO2hpXGFNscqKLJinUvqV6t9ZcHSE99X
akUbaqFx5TXAkLITQdklZ+n4Z3BiVLEOiNih+7tCi9Cj9/GuvXEj6QDkwuOQY9rrRc0ZGJMj47gq
cRJ2uHAfX1XCOym0l0binyK44ETG3Q3AiNYZCMuP3JRMNsx/qmeLBR6qgNXG9HWMCGE6kigYrr8p
xotFbfTJ5v+J8lE/fmkVo8L+rebt1KGdt1RnwdWTXakC+brz3i2Rv7wcVRVkgbAWaHDSB0HxX6ld
F/WiJ/FDkmxCsoyca4RMvJuO+BPAPDpePk6QCH3qW+DMlbEMuj9GhFgZPpAPIEnDi0HxObBMzJoQ
tlOH2FA7tMmz8uPQlkH6kBk257Lw19Uy1GnlQhrQL3nWwhV/xAZtQKdwOeuoqQX4cZu1XKQlS3Lg
cFbR98ROT/VyrNeQduncp/1SwpPLu4JpBI7k4wPASSyFPL/7jp0NOQ5gE5m6Utn5Yf1YP7eDR4Zl
cUaYLJqHwGYAGGdptSIxAG/c0wGIOpxxTNNTeiHHpt8Tdr1SXIzLgPAyqa4UHEQJ/tFPvjHgH8XH
gSuL//TMTsFY5C/18lATNutyXFjaef8gH9Oc7vhLb85ov3E1kKY/ho9oCVi5uWcWOz0fgitzVLnS
JXRZLmEv8Vu76loTpW82ODHNgse52BfkV+oF+3hoWr1gJHXIZUvzysHHyoKxRsC3aR3y7Wsyxc31
mxUqW3xf4bvSosN5hSLWYjgf7k7w11Z4Fy+IGC+fdih+PdB5u95FFS143kstPYxfyT6b7JbcT67G
K6F3qrbsp7kjTgB+G8bEHot/ri72RHivtqQfGehTzOYvZBF/qepy3OcdkzRe6eBW3NJCg8Tf+z9E
2dLZV/5+0wTXLLVaPbXWRFpeO5+JaXji6c+K2n1s5QGi9wHs6po2RVSbCFtBqxiDIz7WJGM+7V8B
LKb2AxBok1eloThrY1PyFIxePgSZLRI9yZsAktJlJXM5pjBSI1gCW5usbwix8olPXXty7hA/f9va
tCwMrTskbwtn9MpW29Psz6VppkveKMgWVV1gRW+YbhkU5OMOwFcoBfZsVbc0vUwQG5wHdnJVUlhe
MAgtXEHSCvMlbeL/7eZSndhttyN2o3IkpiT0+pk04dnKmd6WGCh7aaDAtlAAuCJD/JZF3vkeBNwq
TFVebQiylwXTLOdYnE3kW8qNmeSFjziWJ+oogYKwjbRXNVyyxqIVOG/PDPabMJ9N1dQKi1eamugl
s+AEt2RLq+EQm9pP5klnzm6quqpObqEriaCnipF7XVeaQEz9WtwLNaebmNidYWENOdEnsdGLZhRJ
3AigB1yuqz9ir8mkHrvG9lbmWwAALhdCMDQms8FNAPF/X3cAJPEXZGMRUsGvSIWk+U2bF753+BX/
Yot45xQ0p7J8hhzKz4kZgSxjmbQWY1Ma2iwtfjrhP6xAKnxhP+eoQFnyRiJWeDX2fGJeNb3ortNK
bHxepElDKZUwjjczhvAsVlh+FSSOpkU/O0UpKEsg7tdA83VJ5eLWOpN34IGiBv54GlZGC/g9mH2v
ZMQxMsiQnQQagI0NFJaFEpPlZzcAOp+TzsZDnkEyUUMJdeB34neKsJPGdhAmKclQKUjA+JpX6Ps6
Ig/oSqwz1rlIFuYhPmn9jA0xOZuk1n66J/0gq8TsHII+BKt1jqNDpqNMcbAAdyaWc+5LyvYVLWWz
qTMHxpCN1hr4WQ6IIZ1tUeYxZx20PqrLNPX1juRJwN4GUnEzwtAtgnKhGuv5kw8brmp8j7OYEQxI
uq2kX/c5broyPlzq+Tl5uUc84WMZwGVxrY84TEHFYWYWQ695N+Ze7tl2ZHUT0uLgApb1FFlthwVV
GfZBwG2t2YQ2Z6COE0blTlthTrcBDXKXk8kl9F3jpsuRWtIhBedDjqbBrAoEM9gxGlqQHao0rdDk
nggODyaZiQ1PWO6Gbnm4nevvvZCDpr/8dxvrBA+4wohhvQZsr/pHhzthZj0M6QUCaZYX16gMSAOD
xwfB2NFgSxAedkAOtt6D98TlnEWHB/Ru39MM74Y3DwzI5RTwiggqlcSQ1rFZ95Xz24+/zWBL10cg
+uyDwW1fl7FcHENGGr6svza3cESlhVIWrYE0nJ05LsHVRVrrqNqU2XdbZmAzB3l8MWklHphNfrJb
NSZyJ6mq/jXtJ+R+Embt8wte17PWfiy7fz/X28sNbdwSUrXdkdmHsZAkzY86Dhvc+IWet0C2opV1
iyPkF8HYNNU84x2JhBmQB9ykK1K+LxvBBDAcVUkJdm+Rzt9ddt40zGSV8hb8weZjVZMv+GZXNHL+
SMP1ihOcYwZZl93dRnyQ2kAL4Ltj8Gi+PHeVnC8JQrCGDauL8PZADPVxfmtpDqftAVlX7MqAo3r2
vHMeasqnqPPbfGYOE2MoVBmOazQ9/x3kZOtg/yiVbxf6/pWoNld75MJVh3ICw+8HfMGiQDk0xYUM
siMoibjKlXXMPQvRj6XIrSul79/uDHHvTZfA1MoZJxIkLcXbOV3KzzSVBq40wuVfUGolWs1KEK/v
I1RELkAl8AmbMd3fM13+7PrPbw4e1Ru6/TqGDhHQfHaJSDS9kIG7pw5OtFzDZt5dKV/kEsvxR+En
L2XGA5NGdR7JdXd0SNu36ITPGIoPE1wbZYIrXb9wpyc+xxfOLMMrjknYTaToDmEaC36j8DZ/+4Ol
2ICjeliBc54uvTPIp+T2joDfzjaFjNVMAV6dMQXhjllTLeX++TgoO7ZCfBqqdKdtkbp4BaQqvszH
N3NJevv+HOWhJ6S3Yn2WsQqhYOsYmVUDpj3E1a4KpWB1Nt+wVP3K5r1ZUB+Kne7aWmHJ1BpEQlw7
UDrls1u3+1qwpry641pMQheXwxg+g6Z1l8QIq3jqJBAiUaqfF6YFjuk1cA98+beDp3wHojx5SnBy
Gp/W6tl7Z21+mZh03jil2BSPyZR1gkPJTdGAKCA+3wY6p2PY8VAHxojoiosDYnHWbZnBwsQHa4q/
uCMaJ+wJwf4xw7ddA1I2sirDbfCmSo5nnzPXvXg6/zBkVb/ZvtMicJ2BTTDdL0AlOIGz8m7yh6Bk
J5LR5jWphlboH4xQVb12g6wP8aA6zIWOe0pbk68sinlBA86jYLtHUXkOGhGGVutm1d5/Tpu6v6YA
73BHjTAdgF4L0YEeb0h55qN1Ahdbkz/44MytBzfgvL2WncuViKkXZV0Wqi9SCRmPI3WmfOucICeJ
TIqFlG+gpEEFqzTr74OsvEGuevNcOptczl1P/oxZR+yRfP7MVOXpdHK3H8hETrsVJTFaJq6VGoLy
8ZVEXIsxR2GCUSlyjGIwGYspP4PEh3LYSGttmarOsQiFbQ7nUuF34lNW+DFygMiukevqoeIJ05R6
5pDSiAfdYQN0Bx4l7J81cJ4QpPsswtnKbqibHj6KkdZ0zvWC9EpEVL8A5t1MEdVRtsn0IfI1EeGV
PmUMar3GREMS+Humcm3bjEG1WoTaTZ/yAuBMUuZdCIx62r2jCbR/P0OWEdE5D8tSVjTJFz5Up2Ih
2KxX+dbaQHXLTZXwnTEQv4xCgVHf20udB7vxZJ5pFfuXWvLqAjUQdxYHGN19rfmKA1AI5CituW/E
iW3cF+2Cx15a+dmZFtGGl+y9uk70GKEHNzkxNrIchRYPqGPvXg2FrFgkjisz+DtNp75TeiuVTMdM
9oW8J64QJHdlhnNHtR4B4OagTgDLQivdZqXLv3wmi04va0qhsJLrbXylhPGNwFfIJayoiSUaIhsD
jWBTI/lrHpBZ8CDJnBG1796iRXsLQ/KVtEFDuAJ/ev6A/ofQjhKe04ownmiphl6GTp9VyiEt/aH+
Cr3RqyTLw3alaj32wGEsA77pZ0Kz+N/FBe5DX1Vs65PI+REtS72LLo8V/Hz2c21eX8MFW3Te92WD
dWlpb88jFG4HY9wmsf5/WwGcg2hrfqPdGK4gyNUTzFX2vAdth8O90MPWnHtkddmbdYHlV4SiQK5V
qrgxv5jfQEP04EzblTCS+NvL9/lmrDqmCJfBfym1cOeTm4fQ3wdO6qllIZn9uO6Avdgx41qhcy1X
tStBpF+EORB9PCLa0Skt4b7gpXsSqhMeZluAxuVt+r1CJO6XU39FgeP+XP+RJyxpKkZk6wbx3Mk8
sZrTDCh8tnaFZOcPGyyHhU/gWz6nf+j9GRrkXvDfwZ9q1XRHrD8DPwtmg9s9q6eOcPIbeXokfmr8
MR4b3CCRzXsZ4r+emRz3I9EI9jm2DPv18jIrwsMJHr+D+zt5+Hpcsh650yo8qfDOlIMhG1w92Wro
wuDOUtjJ6+nAXgut/AlUUWxdSIKXpcpa+qRmLtC/jveIIK1Un35HoIkUv2taiS7XyrGSZhr7nQg/
yp3udao6L9ZEbDSbcEtH/KheX9/yLkJfV0bUpx81SnXrJOxRMhxf2LrLrEDlqULnXpBPTA8w1auy
FKnig78xL78WVUtWXmQdu6zK/D+7ipxOCNCYlzlvDyEs7czFMa2jlHHGZOzbbP7X6PErwjtpLhfX
Q6HNrCz9nuc28yW9u5+v6AS/j8f9W+JgecEkiuLdQKp7+gqr3FORRseZYFmLhv9Fs8tjnBE8/5FT
hNMu1b+TYnxLLDH/85IDhJCSWo/L+QW7EA2PFgDsS+kyux1WEc01EAg33xExxi3vqmHJl5DXXulw
NWMNrbe7s3tgUpOFqPbxNAVPfBAFynaVYHtOOAqUNeF81dpDdidTUSR+uzsaX3jSzIonmC1DkF/l
4dGg1yNnxRRWFDHQJUpX0ULJ37ZC6ur/4bMkPVAjIqxjd5I0ZvOrL0NrlvsY8sqFGoWkEPvKHcRh
j+Ah8jCi6OYs2P+NaZ9tsJzJa935E1YFAtvtq5OpfBY0zakfGZGo9xiGP3/SjwvDZqYWGxVc9X0F
VHfVPNJI2QCIBVHAm8sUxIZYZdAdSUE2xdh0JCoQ9XB+yQL2YsCZpuavLNEmHqJz8NB5Hck7kYQR
q6Mxe23wA2iV0vpbFydy27NcrVGK1bO/u0NwuN3dTJCQr/csUFyWviayzMkStaXKBsAV8tq4hu9K
cy34qAE4Q7YF/BnqDerDT0v44LJn2VlQ+7Wte9YtoHbPSEugJos6BKWWVyVcZ76lF6qAcgLxnfJ3
TPqP/nDl5TD+pJZ/k2a6CbgeeYiB4AKsIWxtyd6sA5A01eJ/2QO0dhlKe+R21DAYdYf0u41hVjsh
ggFdX6RuMTX7mvA5uuCOu2PJXsaHruPD3/dU8mV85NuMJbKDSLNzwcEZkJwHj4CWSiNl3Z6txWgN
entgk3/j5MchoStuKAwPYQmBHv214rH54bjGKDnicicnAw0GPOkty5hs4er3qpaEbpE2rzeczhWZ
BGuSqDUzxWrAVHJzq/ulZzwTIBglN4TjrloP3q7fSrUQAcleDiWxLVB7RIw8V/utVTwFpzEO6RKX
wzYiacvLqrvtODlX/1rxybb6hn3tuxR8+iMFD5btzCrHNWdgBx7jgbFJ/i99EibZicTrf87obpQg
i1vZwygOBwqOMCGV79rDi8Dltm25mb9WJLDyR8YT8Q6dGMDVunIYeyHl6iUKDYC4tmHjsasLBOTj
5hO+qQmqXYnzJdm3Ochn5rLbQaWYV9jsbgd2KqeLIth5XVmFdVOvc9lxoqPpdxzL17s/o7vA3Yrw
Mhz8Junw+uelmJXI9OUJYxMlZIt0aI4/RxYSUE4an1/5afju4rZr2cae9Y6WDGcpm2q0hIGClI9a
r9uXm9jtK+HN/iBwwZsp7HpRMsXOLSoeOaL5N1vQDmeViNnucyQSbJNHOgi7Lbiv36enLqFtyT+p
ALrrtXUNMC5UhjHbiwKMQcHcTb15FCffBbYuBRgYiGz93flLv7CRr1HrHm8LhzbhgSqYSsvIUgPi
Bn7gl7BFZ8dDtMSK9gNJLWWQF6h4rHcaDpj/wL3mCpacongPEjyaDSkC9HETcPYQndpHwbg6jhKJ
kwPH6iWxXGyAmWOYY13DWftu0IcIc8WTlhX5VFPfZET263evcpTZYA+Gu6PUJv0shz98t6sp4T3t
GtKmFASpEOr/vHEs5nN5BL4K9ust5BWEVBRbtAXZzYkSBvfHnv8nb0gXp1QmoeX6RfOEMQpq0v0Z
N83foHM3h1Tza7ZL92CQ1XzGoW/qYzSNcOs2k7O/2w5Ozr653ierodt5vogEvqRNZYVqrsJnHjQx
CuJfUXQ82W5cLQIf0oKJhIYPxrmkINMOF9brEhA0pQOagyasgyCpo1uGT3EFvxHAtEeqVpR5GXFY
bFTBlUDY8Ep1zOY3/RlzsqB31bJ3lJyKZdPnobAO7YGrJN9JlhFRpPjJ++md+XIcAx7p3RL1g+6M
RADwa57iOikCF7d2+jnSs0Xh9UedCeRvQBGpPfDBarWQ5DHMsBGruoCW8y7yvCS2uCS4Lo2dqbxF
vyA4bBP0XRWsm40/cYpWs6b6DtPt8K5/LvloqZfkv087MoK2+1amMGMJsIG3C6Rrcew4CMO/JOUA
ML3QnaMOZ8/Mn6LJwWcZB+/ZfeCXnKlueQbA6qA+wLL3jOxoJLtZUcbcYl4gV5MQQf/U7Sm1rzbu
14FQSouWhpm5M0VKcabD2scTQiSMnWut9NN2XgrHQHRpmo0y0qZZky9AzIYUl3/hGFaJM0yGssX9
/Q2UfH9MIHEGRVBHBZPgeFUJDs7TraiLPIOzYnOP3VQ7IC+0DSLk0Iz22aFaRgI7yDafjXikuI+H
jX3RAzvEfVzr0MwTwEh2SidyRRonvWESwqCehtcUIxA+9sfYcOkqqlsHMQCwNqkNAVUWY2b+2Qoh
POD6QKeE2W/o8E7QW/Zo2nfPDXfwD0XNntfUp+wwqSd0PGNC/GZ5tEMt4kRoYCG/PY/Nw4aqghsU
Q4B4RiRjOyvJuU5F0Sl/fTIzJJ6805IoEPnyfaRPTV9u5LenGNPzyx28HkHLgbRWOPryf3MZ8buR
ge/XQdBL9Wm9IIMi9eKZta7dm8kWlA9iHCgGxcDtb5w+daraP5Pm+slyXOeKSuYmxWhOWT6CG0Vv
k1hfH0NQ0zZv0NFBsQhbdAmvJ8vCt06/mV+mNhuS0Kkjg0tsqyBIzEDUGyCgDzQUwZIj1O1/qbfn
uvb7byrxqkDOThcgFlSpBKpPXkQ4ICaRcKRoN1x572DG0qOD+Bgzohxz1t9skqqGf7PMKAb9N+Rp
fPCypowLjssxjz+BOyDW9abpmN3jqsBJaJyLUYlerQ+xWdFf5ZBQoS3k4HDiQ2mJFBYgMYEpZu8K
KTzwsR6NIC98/CZJqP+kK+hTVcR5xuXmjUyf+1jQLy95rA/VpsnwPP9/0YUzopYj0Cz31YHa/hVN
X3zF3O23sbMZpOJa5UpVAaQX8Da5nAwGH1KBVXOgFKo7xJneHdMOHoj6IFQtnLk5LrLkqvyLeXwM
ZxdoFvkCY8NBNj8wT691NGZZ/cOOe7Hi5JaWDG8PqtWhOsEXKZ8y4nK23I8vQJR6fMWEMwooKtUe
EcM4enarhHu+YE9bx+255Ul+2YWK4A1oOpZ+BOnsoXoHz/9VPexKLLSIUacAtxud3RvqF2XotTYF
+lZESKieHzBUanbRUb8SIBTA584yZqmuuwvNb7dWlo257TldLbSPCik9NQ+7bx8TJgC+cPkUKIf8
IDyU9V++s4T1qljB0/lZ55ESkR2sVWd9H745XOitmgJeio2LLXwpE3MmHez8EUA2V6/Kvai7z2Z5
qK2/D+UAEibpwekXC4qD4eecp19LAqz9V8EKw+4W0jzouhBwyNia2fm5bvYFIBMbH2I/l8gwn1uA
uYMThRUCJiA5yxV87fOvNf3tt/lkft0uZpqjTk3lLEoYJmtbIyUm3hJH0K+14V0+AJpNayVUx/Zg
C9MHIZ3IxjJSdMDhRIcvtTk1kH6G8ZJFXEixxPHHI7wskvJBZlFZ9ITpJVEM9hy6xDah7MtC+zTf
AnSpRBdmzuQ70hp8UFLUqH3wJcD0qfv4jfzUal31KU7ncp44FVLi8KKYsIbmhnZaK7b7F4LDmG6e
TiSF83ynQbuqoRa6iiKqE+2+fTgB0YDkglq20pZcUgWMwv1R/VKW/sBk7zGA7oLKTS5JU6Xhpmgw
37zzn/5fvV/mshi3JmsSJgfMYX3nzVTvvekh1PfmtMX7ifyH12a8mFlrV4vTFts9Q6jfl+decCUG
oho4iOUVT2BEnZ9PwfqM6hd8Wh0WCrQ44v4ONslbjM+AHFQfM2vy0ssxNrdsNsMkEzeVOzE2vLZ0
kxO2zj46DLISgpcFTUMSRWFXpdxEuM6IVDcM5o3svtZ0G/abEe5ZMfUsxQSMCBPurYbovABu98Um
dAHZ5i2RYKDljfkmdP8u2/XDaBVrcEWBISshrpgUObJjtA3kGASnovypSx+7hA/THpv4V5UpcuoK
RTqzAqhm721W8gcMdruDoyZtz97Np/1jJkOb4/CxD9LrSDO1rycugQFZuLO0beUx5X42zy9Pfa1/
IPAEclHrz7hIjv9FwSxYrbHhjCzWRD2b/8ad+IssRpM9X/5XLM4NVHAHogPatGJ0/zGhNETFu42Y
f/Ngrn+k6YjcMMVFIWztWfuDJPKBuHE7vR+7i+Y8cUBhrXk7IGHi0bhU4EesHSyvQXGnFSvnqW8R
7FxqQUprOhv+sIl71wSImIoa4crKS4oNjqWHUaOfLWhvKNpLmxJlaxIZo8Ilz7CIffE3WI2LA6hw
Co080AyXbyuIem0GWoZ3xZKxBshfQX9At7zP1n99cAYn2zdTSB0EreudfYscVfpAEFePAL4sFczZ
NlOrMOQy/PYF6EQwvP9X9ydZQFzQtnkMc6SUPZ7TC4s24wS4nRzlnTqtXkSegGB6im6cGOyWKFcA
deD2gSSkJ3H1QUas0zkNsG3h15VYQTAETCIzu2EqLJL+2ubha/rMzQf/tftFCgmLzVcVwHEKXayS
lRIN/XGmLvPNeb4o1v9eJnjzB0EX4lwAwx/IRRMTYbdIVy7UJfVOWZlQAw8haSNhhz8rQYIOUUF6
zIpSBg625vbtmfPvaaZkMxX/CPutuGEt0C5lscse3qBXooviDfdCLXLMFJjaqbXg0pQZpq6w6KOU
85f2enmkNcQalIa8mMwUCb6+dmL/y6ENhNbFZu9cIEgpt9A1qiyVuY/6J/sxwkKN/ee6U1F1wGYG
3kT2gh6KLICgBXgs84i1U3U/136fODFjEcPIkeJWK0HvcsDr+zO1yS8vRrS7anPc+AOLoQeXvybW
94HOCYx6tTbhE/vU7bLYWyl2Owq7lSrqm+DNFxaiBT7spkhFwxSlXT9s1JIMuwYiAVIBcwhtHLYO
mj/xsQMk/Nu97z+vB+BXEhC4TxGB2hAmR5JyJ4fCLjSPSvJjp4JAVVBumoXBjV3HS1vfSWfGdesa
jTAZc59NdzcXHKLyw27Mp/7m3CeJf33KI8A9aUR9FC7qvq3MPyjwuiRlRF13S2K3D3iQjHal+3Me
eX5BqZqh9Pkt17WRVF0zf30pHdTeh1cYQruLfiwbgqRFtpzjtV504Yj8hffVfmcGzJbCnuBq/jQF
vXhLKzccnTdusBNR0XTtqe8/e+np44iTTs6YkIwti+k3BF10kNrmW+NSySqGT6ju72PelllLc8kt
jyLGxgtSkT9vuufQaZ03xiPj11IwJvbg+Vqu3GgxTOYUvtqQ/L6a+FTIkrE4LavGG3248/Fiehap
jiuHBN5kRp0bR10TmotitZB1iEr3g9V98mTTvjdUTIibS/5RuruMxsF6k9iDCuUOhWTFgNzlzzmv
VzDYJCMIn6Te+NATBB5t6w84MPLPbZ0z1nPmUIog4/MGQE2tC+gXzZrmt0e9XBfqFRFGpXDxsJxF
+Ddo7DF+Utjn5QS5bBXboNvpAsZH+XhMEsO/do8bLjAAEOA5ORV77JbAnUgcI+Dsy6xLib81MfWl
5eEM6lspIgSK8bcmZR3liTwBsOKkZ2iUDzL/pDppKPct2+HTI8JVoqmyh4g7baNKU/mruRBtnlvb
4ZKJ3I5VF9/Qs+QS4LnPPZk22z6BYyBZjZQfFsNuIgzbPkv3S7dfMYQt5WHuwuRLI8H6nAqY6XY+
EgqpOMqOcD41W31vS9T2NijsS6K+EDg/0EVmZ3L4b+sFw0hQ1FCjuMzvrU0p92UCw3InSWeo1xFO
JefFlqjEr9LtJCZEg3+DSfrzSelbDMByF9q3K5NalyZ6ZKTrn08fMKlifLIKo6RxBTqix/LoyJOK
13wR8cU1zx+bBE9vl7oF+N2S9ehGeQHcs0FW0JRakvxX4UAU/qvd7RK43Zl9bwJSClE1GY3HYdgu
xglT95PtYXp9AyvXeqqwpXjXa5oaMtDldpYWfNuooROIsdu8rrRqcyUnsvp2KtvsO2dUu7Cgk0uN
yNihbCAqVY9HHhHFLxV1LpXeoOEENeFeSIPFn6tlPFenjofz1x0iIJsLCABe1Pn8TDNLOZKRJ2xf
tyomNSgYK1dSRkC0BH2PI/6YzZTMldZ/GFZ3SGTk3RSLHb1t9QFLZ9HdCxsVsnP6Hffufgb/I3Hw
WrnbrETxflHPyr1q+BmAEt8UABCgU3a7T2oBFqK5D8VQc+sZDPbDCpubsH7mCVGPiZ1HcPkDoJSc
QhjSmJ31HKv0zLOaB6zVhWI38cVrvrWs/uZGaNYI1me/J4doxGXjRaMhltWeRtF2y9+/5AOd4UmC
laYBehWQ0BSmbIOZfA2LkqILJq+n8KplZ3wIvES4Y1EyeCC5o0qFAySg/KOyhRuMV40oMz7eXy+V
VUeHux3YBGRl0nlUwVNPKpxh+cQurPYLrLvtRFpeYixCz2bk6xZ1YE+dLevwfQzJQb7qXnMY9G0y
Js0DsT99wMM/2T18pjh7o9An3NlMy/Cqy/+lhkuGcrZcXuyZf5lBUVFO2sSx5/YBQvKeTN2UHmcy
D40g0G8VCDb4ktcmaYJmYsjK5e+SPUMMS4p57F3vC06IAkhzl3NjZISuZ3PPKrUDmnPMvadgukbe
Sxi9Ghq0ISih+Wg+lYsDjRRdIK8A4HNCCuSq2jZPUo/rLjPUQ46ne3lSrrsXb5LOA5u0ySQFawKg
AkQkmfBGCDIOeP/SKBNIGgfnKW6xefSPzW/O6pmmPyO80jOthEbi24J2Dd+ivgqyC9wTHKaoYv+3
TMjPPM1d2/HXzdRN2scgGQzj0iFPmHm0VOsxsWUBkddd4O+1Fd9wYzWs5HbfFLbRFOxJdsoUidCO
b3H0Ec2bN7Rvn6AfIasjNwAOgPo/GHEJOxvwlMhKKl2YeOL1wMQvJZXA8/SFC+/iCs+/SxgChIZz
/Z0RjdS1Tw1DOPQog2VHyT92tUQ9QugMJxAzRk08eKjq0+nLqYCpgS1rDwTc74V3p/h5qmeyxWTM
rFHWfeOflrVL0nIKphyrRpwu2a0S5djMcwPgtGztM3keXP3s8JCohj8PE9NO71nyA/eQCXBD+ZTZ
vs+SeYBeNa18ZerEOksZbGqX41LKldjM2ejdXGyNa3sGAZbwNjDKc2cTbztPas8rexeXjGSMe34Y
xKVLq3OUWaiVy5dslFj/gK0ymnZKyxBtmhOdFAGcAcJ0Sh8NSuKnpr478hskueTf6YLgynISJP4t
s232r6oPIUg/Tj0RFpTe4rmSCanHrF9K5qMwlqhbFAWGLSZPcdjvMXtd80cKxyoFAGMVFYweIHeD
7SKopjFEXiTA2d0X5+UYX///KPNoemSLcXS3t+ZB/pct0K/+CAdCDy4bjb45ojhZUs2Zxz2q4sm+
Dz7FQ+aMYyhoPgRB8OeuyB1qLwH7G9lhjF9GbxqcMo4VwOpk6oB6MbN4WCB1spSm1dalINdN82Jm
hWl5cFtU3FAjhpFo9ye21MrFTaQrwa9URKCmPxwGLSLGBnUPEiLoZA9QU9H32hIPvxrdYPJ/42ps
EVtXm3fpPppWEcuXnZpc/yxheL+mXzTX2Z/7z0Aa0utgj/94tqm9gpC6kS+5j5dsjuL//bnC6G0+
LxGkJqRJ6o1A4F6C69J2o1xGvT2+cPQK3T/UGqgH6+/7gsbW1N57yD4d0ghcFvzAo9SgZqA4PH2i
7UxnML0oFKEv8s/Y0bmnLe8uFzzcZ7V4sXImRWGowKj7FF6WUnsmNxGiH35rqH/+P47MBGYbYiPi
M72zihUF0xe8JP00syUwZUHU3HYYrmHSdkDTQBqDYoPybutVH8+4ezar/uxRP9je0f3hnV2vOxfz
2aQieiWbVeUxVH6uFH2/OdYCuOobrr8cSVx30QLNRSHT9T+dEy0TZ0AizacD7vrXi/vksG+8HrtQ
/a57mGaIX+5ic/u3voi6SowffgLtlrv08yNoOOOd9zLd52GTyv5ysYrICl4P7pTsnHo665hfC5vK
uEPdxoIF9QhAqLX9BlwOA0F+NfEdikfGbHRQZr2IZ54RVeGf4z28t/Ipewc6ZcaQxjbUxAGZYZmV
In9p2bWR/DkfIprqwkXQuXZ+v2fBePNX8/+v0JgaXgmPgR8udQ+aH/r4WlKfR+aIFaaTvFF3jz06
se1gvbPkomcc5vUsvgL7VICMp4LLJbWhCTu4kcmS4P/XsqtzuhZxgUM1BE8H16y2CncBQU0Em6iJ
Mkl7u47zrfq9qljTb6xaUpRtQ8+05wtyH1IGiC1iGnbUNPT5AeJTt6Usm/z3FnBnIUWRvj3HZXWf
lzykG6ZyirCJChOAQfE9I56f3y1yjilJxviez3zJGrFSuN10bSCtUA0YPD28ZW+djcA8WnPH22T1
LiTklezAZJhJXsO5dETQZTRoEDryP23YM+AQKx9Fh8BdcfBK+pXABy63Uub+4bD3GMWccaTMr0yS
Q6CW/QvxnYUx3VMRGN1/htuOPUphL+1mbr9M4zSYdmFmZUJyJDrydW4BuuUSjaRz0PCFw0X2h43a
vvlf6eeecQcAoXnoGe4Ab4FO6JlIeAgZtrRSd2nxZVM9PSAlAUY9lYMUdeadHtqyqIzyYkBOuvSg
4O409lXq8fpIUSEQvUNnoaIdA7BOxI/Ukp+lgRaEV++O0umtKYV0F1IPUfy40fET1ZRFej5I+f4L
0Sctp/Xsc0OSLgtOjp8p62P/py5E/U0FUPkeWlOqNB5gPf09geiBJUhYpdg4n/uTrAUGlj1gqe+R
YDRVzd4CaTlclTpx6EVYoJEQBDAcZFFMeiIMut6nVUNFaLTHnYxUcDj+KmiK2tm15ywZvH1FYgbr
2At+Xcm1Hl/U4cEplyBjpbctpN5S1HlfKMhTKoiEcOqhgOUMaFgTwZ3hmPas4LBAqWz2DrPMq2UQ
72tBLIYDbRroapTHLe+OKFJDQwEB8FvUkebefkIy6lh7hcNAgnO5M1/MJJ1MlIyFVDevt2tYOWWB
82rvbiZ7GOot82jZmiIu+4rvdD0OCY6IqUN65b8a2CJjR4vPZmEOtfEtF3W43sHAuEfxiKzhQQvn
ZMw7gjIs4PAhlifHpveErZ5RzjLxqnH8+20iKj6l11Wzhyiefo5XkjjfAd8FZQVDLTN7ojHPbjlj
iV8ag3fRrTWHchKnvwMPwphJzdUvm/ht9v3+IEE0AVEmm9cBYhNwZaaPRl8H5SmaTwTNGdjZ3MEe
xSrtB49NoZdso1HNZoI7Wk+ZO+x71TWk5hC+dFiAwviR9uE179rI47mEPl1lUA67N2werk1SSGN9
c116DHqZqNilPpECR/5r68LMArUHuao9wKKEPp5s01k2l4+lL3f6H15e1V82Q8jXZGDcne3K53O/
Us/pFlKNbiIjvAjRn0Mtq06NW/GTvcQuyrgvL6NNyNTnr6nS8GzbA3CTp+WThuwSUFIndh1CL4+L
gfi40LbkpPZVXdvdQAuyTZEOUxvFCFZW9AiFHJfEPx7A2FArEBdSezUyMmgsRNcICd2YipfkegNc
241bxNtW0NCIwLL54vldw3xzKMp1LQLqe9ZXO21gdwXaYVrk8OmTLubkLFzLIoaoBjlfoy0ANGDJ
L327B59xujkrHjRUCcAHtMXPAPQh7PRKy4Qiz6LvjFi0U8A/PJCFe/WqhIwMfPQ0xZowtLOl/DEh
JkGTC8cNGZEO7UMo1X5MbwMObWhtyk4Zy6Rnr1dSTym1sIGzRaSpNSGtPYqkdd3/OQ99SK0x0CLt
DQaGrOkN5Y1GlNnAP/0YHTJcr84kngPw92P7xxVzMkprX3KbbS0Uiz8IqpqAPwZ6wt1WNkEf5mle
rvqaQeszRUIsTXRGjTnMA8t8CCCXIY8UIWsjJvkGVE1tMcw2zI0M865WPIWS581QRAPwnuMcH4+Q
6oObNLhsxvkiZk9JpJMWU6BVJUyNHW/4e+V7ywIoRg8kwzcHMh8g+Py5FQxZ5YhYxP8oeV2yt6gr
pPKFMFcUS3tLCPtiWmDAP+86uI4LTFjbwitcHk6o44x/fTxPDFTadTcV35WpXhamUd4oZ7YxfgBB
pg3OhH2wyj/DWdN2KlOw5L9Mdn1VgczVx15WMfa1QGPt0fPzAXiNc+JHynU5kwSZxxenAosM3To1
Rn2OrNTq3GBTxBPkd71xBAMySdX1VokChqsSACdtBXrl2hkIfrS7u68VtLgP9r5cUj6v/Oe6SLCp
SYuaDcQBOA4Dse1ZpEjBamIryg/vuIuFgGrlbK+iFz7B8eJDC6+jcQ1dDUKllKeY2EbNioFdLcHh
eOizYi5EP+ub2I6nD3YcIRe5t93G67RlYVdaceOVU8X4kgTA+xMBXN5Yw48frAXdPsRC841Nbt88
PAYgfpm4psZQ841g8QjFu6HEYnayvN1g5TUSZAk8LQtp1AKBIrUSih0I1sPGlRmatMDSpicSKrHW
coZKu7EethhrMHdqEclnZiEIbLBRXgIsaiHEZB07GaJcr4CZKRnoAWQzfv5GiorPEAZzWHKq+rG+
VaXEZeyDxjdxkrotWvHaiUidrUPLs3MdRu19bQ6tHI927ap2W7u0esUjDb8f2Lds32Qj2sQdcSs/
O/YDELkR+5Iol90//PJgaCo5Kcg/EU2PP1gPOcqgwm1r0dnhpB334XwndZroe8jD5CCE3MkAgJBP
VUyTjl19WR8AxWD2Bub1tNsMZFqj0s4f6c8+mmg1WCzx8udRlpzqvkXQIs7T2zO6n4bHHDEhvhme
ewrC/rL+B6nCparHp6eNVjn0+3sqaZiAU4Q8kEtg5cjAusbG3QbrItmKXPTWPCz4DFUz1229MwZC
LR3Yybvq5tge2oit2ShfcHCkcoqJdFB352fWNblcJW2OXq0IUfWmZg3WzWLmm4q0ykJKE7k3+Nvu
BVl/NXwoWNlFMsYMk8UJCNUe/gB1QtLvvVb6hZDq4EVZa8AE2Hf4iTd+CrPafcvxZamlIxdh8/Qc
iPcaGKJpvLhwKYnwjr3o/VdaFe/Hn9n6oc4jiG+rW0X/pdepGfzTyoBjFM5JWYBLDsSNIDmmTPp5
XJzIdHaJgs0vHd/fBpaLbUHpl+Fbku8daDtKV57AtpBvG2UwWF/QeBH2j7Sp4kt74xIGP5vgfYYF
I8jnh0pjVCaxWyNuFCjJnTflfcyLeweMgKkCtYCEdPnX6a7cC1NJHxGSeDwi6JEu1RKIM1RVFYlD
EYW0292Nf93eTx19KY8PTQh0xXCJMUn4zaQiqevvoSOWuK+uc8g0Nx+JC/Au8MEzpAoZa0mjIYyj
U9Q5MQ8nVPm9DMLBdPSce5CgGFx8zUmuJ5fJYDCouf4tJx90M7pHX3BtrtQmxaPTVAla2HGIbmwf
Ru8n7hYMor5FIWZnpu6KSxL9O2C/kuztzmJqJEGUpJQLPJzDAWfDz1yBOgIQWjm6NyuVUUXYwvir
1YNjzkm2F7AOfIODAkWzHvl3t83KtLbuM2+5W0aG7bFf+/yec1SYYFms3IHp5mnmOYqiXcHbcj6n
Ea4H4NQOhixqIX/te2UwZ62RyJMuxEL5Xqd1QqAZy7AE5/SZ/MfwcmKJIgffUrhnIo8YJe9H+ol4
BjJHixkkl+hlsVYwf8Esji38MXaL7FMcYEZKdZ9ebokY2gV6sMwMQ39lyt6ObR8L5FoDgXHeX1LD
AZFkIQZMvRRnT0nkN2TcKFD5Me1ydMDpVR59Vk5mfFkn16mMbX5oY3/djEm0DNhofPjd/5PzMvzz
xjxmtEFVcuurTjnZrmhVwR9DfnH4SkQSEBrNONYw+vPHz0mOjMzdecI5AcZfXZB0BfT4n5Y5KEBl
aGahjvZGeie3p45boaI0O4H9GBSfSrxfJXzs4/1JLslRuBnWqXbTX74DxkarlbzuSjOpSjrnQuuv
Al6bwPj1V2owduzX8ZynTqudcCOoPvc/qLr88hkLE3F25MmWJBlgSmRMqA6uMnGhXb4pMf0fV3QL
Zx5/Vor3Aji7HvFWC8WRWqisTx7jtlGBvyuXCWqRofmR9V4IPlAyinSuVvkLXW53PFrToWsD3JVg
VUF/MO9ZbkzpHqWdIicDIQ5GkEcS9jG72qNUdxrl3yqQUZ+2aCtSQICWDWFOTDMGHm8LGlGPQSxC
STCT4Twuu3EaeHqZF7oB4QRgcfOrT5GfI6VddDFwlPnQhZzRXPSLsMyAGFeZDkJn5Y6abb+kKsmg
YG5dITkzH8XTO3G8DVk5hPMlEdwHFMhqCggFqQq68J9NoFTNs8rk9VOGqj6w4ykbs5MWEi/oalk8
QG+0m7KoLlrQ+7Qnmc+6c+2eJLzO06NWXYlCsUnn7u8op9jArrZVzT7353aDWpmMsmnRTQHwoGx1
c/Wd9zjVnW6wc/aEJJNrujEbugw1EdB668JgKOXolsSfJBq8L2HdMO6/ZgCTTMpOElIPlfhu/5VT
+/G3v+noJgCJDayYxMm2CfRDLVn6KVgX4FDDbEltdIB1s6AMvFf5srF55f047XlyyV0MHFI5mfLw
MlPrVEh5arWJPc+UsHLUYCTs+JDLOE5FbCGCi0PX12KJrL3wHS9EOoYDTissmwQgekAzF/Qlnfvi
J0TFaQK6XYZHBddBhKlpVXtNIMeWyi8hby6bSUTL+aPp3glbvGRyCAdUAQ0DcFCWABwVR1PI5azg
L/TuSFRFuGxogSToWqDnZiDYcVb1p55WJJVAKy1jdhsZEDli9eyUfEmkwA2Q9/t2YwcDt/N0rf74
aZPw8F7uK9bOfTzrbXZldppio1iVCRKa9AOvtP3Y8vSgagZBAgJEFrANwURaZWU84GeQdPXmWG3q
M0WwfVkVo9mMuZf6A49xzGBN6LNDyM2ECLMmaHC3v59KPO9FIeTCpCEX3emdYLKA6fFc7Lpr3hme
dSrrObynnQoP8SRuzejm0jESKM3teWa1v8/ITRnz01wbI4VIOsCt6/+W+d8gDO6DrINh+HEVGIzZ
X+1AKg6hmdMXTBxiq6wxibXVFc1NeaLe/DXeykccenmQwuOKLzuvu+dU5dZ+08ppUiB7wFYQ8Tce
NMuz2eN7SGXm61GzILxH4H5jtDx3xl7i6wD0IlxpBY0UrRKXpPC2FQNgdd48yoXegbn76d6nQm9A
ubAOrFBhfAJ3FsqfHQ7l6cHcsurYlAvYyQ2kNs2+/XHMDlsJDnfAljkgYRYfYdRhBv2a9L/sNLf4
kM1GSJZz70K3ar3JrVsWccMDPZ4Cuho2jmBJkQWkLL1TjWZlNiN/vucXR/T8S6HdRvhfkGiUvjhg
y605yUjOmRQuMscNXprxyxeP6EzinrEDr+M/QUyCmBQzPwKQs/I4bnQTy2Dor/PdtJNdqUOKyn/8
ZV8LGtIsE1lGsaQC/b0QOVLgeT3SlLq8gQysFhDJOzxQLRR8+h9C+1zhN0ZINjTG7WUIx/1rhdYj
BzR4COjsCvUQGpVLYGo/Do+WXhNeY6syPNFY0Ylf1xumOKg4ubU5hPiGG5lVaib37SvBjIB5OGrw
2aZ3+yThgbi0qzOgcGvnASMJYuFxlgEjqix5q0t3AfqDvhVdS7prNSvuZ7yKVU2bxuFYYBnTZX00
AWJprnUg750q4p7hEy50vlM5T0t17YY+9HrMLrbsQJGCK73fpZRWvdvKA/VHMVvKX7AAcUeOXf/7
BScgEj3jQccZ4x+NIB7zTBBf9Jb0e/uNVlBkEcqjttCNKtlmZHAYL5iL2xLhQGZKBYPX+5YMUnRf
JwCMpyT1Y91VEyLi5o6l1zq9JZXQI13ZA0YsA4yissPQVv5iJruh1hJ2x9YyB+nbGxJuY8DbjaF+
CW02QXTowB+r/h0ZJIGaofREI8Vl7udnQi4cMD94+Qp2dOWQ+3gt6QDa16U60aqpVTn1F4Si7cF9
0nO3quhyIF/T60oIJKPKY6lreYymkJ5EraU3R962YVg+oMB9eJArS5nFN4S+aZPnTb/Gdf186CfL
cwSrXwM4VrkvW9ILKjafTe2ZdXy5lkKC05H8vxJbDw9CdqIflqVifHzt0KJT+mKAfksLmi0YJd8T
0p7IFdAgMegXB5cIsCiyveqxLwNedW/CaQZ+J4mmHnkt1njJBmLBhBTl+9bdI8NzDCqRTYe48SHh
htY+tZPvrvSS4tezrONujqAANPfa1WXUw026XuPJqxVO426oWeT/qEy6r24M5oEZXXJGlB4kxNJR
Aol8+nCBwQZPOBI1FhDFQauR7oDjH/486EF8ykzOi9KrTtCRjjhNwsjAQO9xBgqvJkaImgWbfJHl
PGGr/5x12sADs5N+3nxM6roHHtOSkzOfGhHYIEdBCxS7ikuNf4dLB7i+coR+LNpuGB8hAh0Ze8x4
eWmrH3zhCNUQzTQD7P/EBwEr67+UlAp+BROc351ePsOEwjibUNBY3qiuJD1jOwHzsuKFuq7J4rn8
ZMJGYS+V9AobyDV++edzHWDS8RaSc1gjEvpYGgYMCASk8fnFYZzGf8xDAP8E1n7wYBRI9I5ohnEK
wRo7pzeSXr0v/XsQwLDPxIjR1bsqqU2P6+AI5ANswCjlelFuH+bgALdiVR4ukSbFYLKVqFfxg/2L
Su5GlPTaMCRLAU9bIrjgIShuWuF94FRQLp4Jq7Q4e80/Cv53BlddBsZ632Y3LXCQdZdBWVrw2Tt6
0Kk71OFnR8Q9uQqSLVLEYKyfPbxKAkdKYUW6bmkQLRElb3jM+JI+PAZHfh2cFlFKd8Q+WC2Q4xba
mam5IatQmcvYF+f6UuHqfQX46AF48itHKItp7PDwH+TdQlkFD4y3247YOiIMQHUrZkIwYtJ/uutk
+zIrMMa3GNoF50vuYnL8Mwhl48+XVeQq+twGQCf6LKog1BV0NA39bYo3gnlu4hn4FRxnjPPyYnJE
fsvRSBLKYCPsnITsOOK+zcSAK/7ho6SRCWXwchZUoPLmhWjJYP1SkAQXYwgwgEMMYGUQ5QOf/MZe
C7xsn5V0YihSY5Pp/MtoKjPzsrK51aEVkpr84lQi3WSWpFKcIWQ6Y3mDTg7qX6pgxGifd5gNxw5W
biFndQGt+KQY6DW5v87x2Df0aqVmMXJC/DmuXsV+Yuxot5XfTis1e+HRMwNcmQRXZh3IkoQM4vQB
nRkAXKP+s504Mul6OgKH+RoYz2ud13219EfbqQnQs4CCbpNw8drrCLZL53iTBxh9uuahJWJ7rayt
eigMaBN82b7QQLkUUFnttf44yRhrR56VwVqTdrkptcALqSlMvf/VdbvpBxFrhibCk8eti/lM7D8w
R7RYBZjX+QJuOPJ0gZiOQbkMiuv5tzQaCwI0FW0FqVRoQnatVzMKumpExawBeMWzCRnob8hCeR9o
0EJxxhEbnI1h9wCUewoeKSgVvprcu91uHV4prN69sP1E+XpAQpZqYrLaB55FuXfwDVE/tU0xjqHO
xDSUmbuBsSXH45Apx4Ey55Ll6d3AncOoyMIKAOO9+SgF0HL73RiNBUlQ0l+c2PufXTZ5p8j6W0iL
B3hM1FsjfOGZCjjYql1+7dhxPtY5XFEtYGBB2T7v7bR1VfHyfKnid3eutjnOcsv4ls3wFxrnDgg6
P9Ip5T68sVxTrmvoaTQ5/JEYQXjgNA5TPcAzKjYCuzononYzQsAnZE8bx38kVjYCJhVzLrGUHZFD
hBZ9C2zGSFjAkT+ZlzbnR+RDwxef2pQPFDYxwfgWkOlsatQPjIUw2ALRSd3/shzsDRPDFpg0A1g7
AgPLSxHNgk1+teGKG7gEVolqtBz9dffbj1RFPdADK7w7P0j4C+aOYxEPzaMGWFiIGNwVJAvtAaxn
am4jJjJN9A8HQD2oOXiv0KGJGkQkqu2vGQx9rOTJRj6mU73rq8YUekAJjvfya5bbSl+Vk3cAAi7v
jDvyTAPu0LDsjOHLYs4Q7nGXEidRCE8+PkqpxOfQ6gWWX8flEY/V4CCwqSXKSrwM5A059EaEwxs0
lxw07s47i9wS7i5wCmCY4jROcFz2dz2a+zD/AxzfUN6xC2wlXLBlgN9HZEQWcW9JlLpWvyu+Ydxb
Xl/d+yfaElAaRsSJysDb+QfkMnFOSFIVafP2WMuS6NIqucxJAxmvI3vb76xoGTuw4vlBdBZPLja7
qyBRKlQTirDUgxz+xsXAmNNBCWNk9ngukeIEoa4EaIOpeMpGXpEynhQ1Ll5mMi5m/sqk7lKf+oEA
fZ2RdRLlPXcEKu5MFvs39A68zHaEzOyGQTplVnVW10KFT/yVwaphJrJXxklPnpkkJcfnLfCBYNZa
C0pcWvUiaqDzROlXMWxySLwYRTKQ+zmpIP8LMaKzaOi47qNNIrGBEjX/iwl8xtBdcoLIV3WkxBgx
JqgfEPvzBHmEziKC73oAoaNE0udhvd8KgVJDg2Y0bUD3GpXV5n/v4s++2u9b71rYyGiHLobQLzdK
UG1UI6V0Re+AapgpZBLAPZmGBaGNfB4Tc5qlGErUQs0FeO60r/qBY5SKj/YVKJEAikTaratXCPI4
36HFRtiRAJ1vnsgrW4pONTmYqj/fxIEMvXBNqhmTfpzbyLUX3/M+cAa5HQIZdOI+HP/Asgf8ow+W
5GQHdMETLuGCz/aJjzrOAlKhPZPgu7uBWR12FwGcidCQitLOAh5V4Aopk85waouLSScunBO0q2Gp
caJBOplcUS8sIPNArzvnjM5khNVMXZJ1s9xo3SVuLGAL2fsX2QlnpSu+lOKBRIKVFlcFGKYPPk8f
hTlHNkodsKhXNqBfJankqbKlLeXPGK6VVb9PpUbD30at7YkKhgf8p+kDoGLupp5zfrJ7XbSABABd
y29uk6PT2g0hg9PAeNdPk+47oDI/JcTmp8sCqIBTzKHcxIMXfcgNeidU4bownoqnpD+I1ptqSht1
xpbAIMDhcqAtbIAx00TRVidttsDk/rZZftRFGMGUUGrc6qXvabASYz3MQBi5iBY+Ni7HXUCqVjKv
t3T3PjY7iG5gY9U0AEX7wDnBH/4Gz0nxhLGQumubqrDIrOO5qnCyjOy9CfnA6gnADOH90ogliIP/
+lnWlsi+7wFhLgxONVRIsQOcw+rsKUVa4JMiMin4TgwEgoFHFK2G4liy3D/kTYNU+LvSRKNWomij
GGMtcQDqKtTg0Tcfto2Sf+TEQSob84CE9oclIQR1tNpn30WldtyGkFrqaPR0hGM2HdF0Gg1oGLBa
cxVnqkRiovD5MumQNtdGBca7ZsVKueqb3IOJt0/ZPzuDJHJieAqm41EWh5wzVCx0sGzy+krllFIc
b0Su63ZJyYhE4OGih5Bp7Y5v4X92rmKETJDb2C4UMr6aUQZR986XfmCRwaR1l2Q+q5545XLeIce+
7/75L8mY3Zt6qIivyAieAdI6uLxpqtYoFhLEvfvTgOSRKLeMQbEDzgUJTDjyTVa5VrPHZfY+pN+H
pq/me9R1rNxp48va8ntxOfmndgKycfRAud8l5pPepitKKcJG/Xxyc8lkDiSn4DV5mMvMfx01cupY
wkUlGfSuw1Czmd2r4L50eTNN5Mnn0bFjZ1znrCvRn95RVeVKY/yn/InoG9WPLafUXRoLGXFYBp98
ZRgOaAV519WZBVzA7JVCCxnDGyYthEEPwzAl/AVLjPOpPP1o2xyptCqCQqb7drA0uDfDbDYsC/kj
XpLZceG+BnWW2t4uhjfMb9aCVTgm0zuZT8ZNeEDnnpV4l+GV5hq5gOGwBpd/ZCo0pwZwufGybBCU
SXaSBih0w19e1Pz5blDP5BEd2MVqdj8OCVSzEeEfoJOi9BGzoCAF2rRj+juyopT7zmTx+LX7YUmm
RpToGQTO2BEzTYICCrpct9d+lK0hcZQdzINCJcI5eAb/4L0+D4ofhKF9kqJSDzZLow2TVLS0TDCG
vwyyHGXvOyrEX0VwDgHvw2RE2ouDIxSzRdxmDVME3/gG85gyQYDPpVQ9w/SxGCKyNkM96UNOUFKB
2vjFjFIOIyG7sQbqU/rhpSlMDfaRjRsJ7NG8GIHHyW6r2OXtGUDxhSh2C6mEBWotXPSf/6mH5zZ/
UMDiT2/Ogr3dl96jFTMXr5uZuNOmEFJAECxSb5+bXKKTxAl7mWEeJpk7q3mMJ/tWjS3QuCTfZQPV
D9Gco6HkNuuq8xSeuCCvnD+lxUuNLv+d/uioRcigRO3Bq563XJdwOCngRsQQ7TnMt9NUrasDsz4i
dlu5oY7UMXZpNmrHF6iUk3nHhmamfEaWP0yU4mwPsD1PazO6TKxSxaAhbACBSglRm0PsW8/Cvubh
0kD3g6hi+9Yzp645k5Cqcp91w9neMqEZHUtb3M2kUX0FbKEfI3N1mWssjP4iJStquSCEsQtSgEor
B8R8wjOM1DNryTZCcBFHoM17vvQlHrMkieNtGhpoN9sWIP9z36tWCpdBsW/hEtps5y6jAYBR9MmB
xYAIVKdUvQWrq7Iw84L/HUHMnOr1MFoUs7oo5QV+vZOfTSYbyS4+g+JE28F/MJC8X65wkk5/kRlc
RqkJrFxscpwRocfSyKi8PYro30udUjDCW5tHEwC0UXLymHckOlf8rwuw1k8mNEJpHY3k0waeDBPC
OnpktvZUlhA84SFeRhGJGW0V0tHTdtGSx2wWsC2vx3rzjv2X5Ct1kedORkTgiFhdoXOgFjaAjv6F
4b+k4qSKTYDeU/0Y7vogzwbuVPEQkf5I5Yb98CdPN/xK9q2ZDi4Sx98hME4ovv141C1/vIqsBl6U
96ly0xiZSEow0qyiCZPeWs/fzZAoK1WwmhFtyOEO3WKS7+9oRq8tVi3ONt8JHfP8qVyNgElh0Ld4
0VkuheIUIw+8dBkMOo9wwA9TYs6Q3rt+uQJ+ug8DhfXQ8DcGVBwNagYuzFIneUOe/CzWCait6Djd
jEUhqjjbGrlDjVO05M0FBMGu8p7WjlbJlG8HGatm4qD4RQqGaTwsI1a+XiLIhnPMqRCezYwJ89kH
BEv9opi4AalOl/8+hR65XlGU9DXFcGWAg8xverMfpADwKRLbhuOgcCgXC7DsGCVPfJ8i+vkprOzI
WiJpAdlkwi9WPBGS0kGhngXHZvfl4VSb2FghH8y0EpVw+ouSTUelWBq4nmBCs544BkKZ8TYrtN4U
raE9oUBaEVvoHfRldnbcxafmRwkRCIaldX+KyrWBaYlT2ZlxLYouKPBAKaRVhkx8uc2pxAQbl9Qg
pxW4FOjB7pirclujJWY4YSyotsL5tSqTFyUSYiiUTzsqpDK2/EB68dKgyiMkVGOitwWs6S9Luorc
xZmnPoDYY4XVhMQtdEsEQ4RZBfUubAtcbDX8TxeEslTpfobzrwm/j0d/Wa/2ijcYvNryXDTKPsp7
0OfKsAcCNs8/ZI+Bz2HIxhxTQTWCABDamDuJhSA1hg0dK/6vt9fxp39HFCl9qAvvUwD3S1AQ9UXV
k1sf+PdfGm3vfqTrAzdXT76d0Venmu2t7HovViHuTf2Bh8S+k7EFql9b+JS9Z390W+BRHfu4v5lx
4jbgA1hONrs53l2jWWpI2eXhJYY1S1ak7d+aVCcbT+cPI+6Lz2xMbijeQtthImc6ZndbM1PHDVT8
jVHLCLnmP8ogRQijwARdimsfeJEZDqdVZyOvs+uW77W3l2iaYamcRHJv4sXPyGJY03+JcBUp2ciz
+fiaQAqNZACVKpbRlGrhEbbFDSp3Aa+YqrGVuu7UDBpT3L4bPbrP2pqhbHllztQ3U0wQgDEKhsJP
wGSxLqwRxb48J3gjp5v+rtrJ2Ppckb9UEMnOhbU0ENBqg2pLoYcF/Og0Q6MlA78VlC3KmUUX4hei
AJnEurktlBLSa5ZYc2Ltzgl30JC2cK3Oy1JR5ywljVjkKiOeNFwdRFVfqQSXFz1XYJmM+dKQr+gk
WuuIPuwsCaIuD45WiVEISESF90LdUR/Rm0NUAWKEBW3a1eZ5D9ITE+0DdrUNylYREGgOCp3/6QcJ
VqpbXn2WObVRCATXOJggJNUzV6tf5q5XCRtjqK+PSONK7Ci5J+tTyWcejVYN6Q4G8URDffNYDwvG
WGoww1gaIlWxCYPfAYZLhGA4JtABvESdyOzYkid83/RSw8g4ODtQS7iT0GRvaKezLuYqMYzpBulY
8YkvtU10xOX5ybjwx+M7/qkkGct5Bi72PNHkTmAGAViy4uoOsG5D8WeTCc7OL4GtwJmfN1aBbfJU
zr9KZHnIn0pC2QX88P17M1etRxz/vlJ+BuFtz/hcalh35ieaMUdN/7DZq44FwsMkCs4WzqXoLcpR
LiwcUoMDl8dVifAbNMiwoXQdAXx/Wet/YUOmJ55pJqV68+m+cuT56EaPvBQWaMk0I/A3/v3Ahf37
4aQm8aa5dyLi6EFfFVIef2cay/mJHI/gqf3FvtnAaOJAUrbQt2wXzcHixzSlVFJsrTT8cEEBdy9g
6XwhOmMnAisoThMB3A42V371jF+l5a1mzhuTkoLNqCUi+LLLpZwA8qMHVNgKhHzmdLyyLUVY1jPY
EEAL8QqxxM2o0tVjxrn60IST8MezJm8YTuNc7jrsApbbRqRpPfU5yIR/VVL1L80MOHt51kiNj1wN
cHtumRqNT+5luNVzBKIwNGAlkp4HsJEsYavD5Iy2H6NKFbhqPMgyROgUwEOhNXtgpxyeMsG8Cix/
dSj20rC5y2VL9dCimB3UBAgxbeDLWonDklOG9zSJnhkArW4Xp3d26qR4eRm5U2LuiFNCiC8Q17MQ
hWOO0eMgtwUAt52VcU7Lq/5x4u2rzGOL+kQnEUciaJkFOv+9ZP+B9gvsVcwhkr9M/vo/igUniLHn
4G2YHI5UOijkCC9M4c9tgdGeu8fApZ6fDzAYVNOidMfdY4wVGjqrc12L/wshBW1ZbAnADhjvFCGH
Dyqp5BKTu3Vw3Mg13NYqPbCcr56FxeEXsFo/wuIawIe0Tlk96ZJ1LGAJ1tdlKAEvPnRfqVsI3UGR
61ou/C3vi0ZZRPgWqTLa9ljFmwEnMBLpC+rcRjgVTzbAbCPN1hXNGYhl7FIA084nPkZpsENYDR6X
K8tZvUkMkj5tbZXFuG8DfCce/4+thxZM46NQ7gmIKUKwhRJLGxvo2SkqjeZ8ZkQe0I+gC6ReoVZf
//P89d92Q+6lR/OCWgHuiJI8noUYOiM5a3IRApDu2sJagIHOWVCkHLZexhvlD14YLWkLt0Y52dMk
+UR3ftp/l5OAeqi4UPK2hDMYP0LdjEbC8UTInnADDxbd2k2GlqtIY9VxOAZmEX9sTi+ExC97DVLq
+qOJoS2WHup7Pip0kuAR9nKL1nn2bq68dRoEQistgmMxnjpTvwOhJM+l+GBoUus/mZHEhpfN0F8k
+phAySuKL57/TZJI0HYk1K4/R2+8s/SDKfody3pwaJ4Q3uag5OMRUaUJT6FL7sTIEbrfl4TiZ6PG
RNKUu3vcjHwfyjQ5VLCaJXQuRiMDypcl8T4zGIhki8nqE7ZPn5oaHg/zeUUTIx8rUbta1GDcKv7h
S7gF2S9/7eE8+ykDR/Qr3jg3auar0TqG+xWtzo6kaPv6tb/nmf3Vs5ujAzHCpCrVrR8nlE1r2SHh
OGaTIjyPVXC+vk7M8VHf4LbERK8xU1GnThRl50PFlUTNs83i9f7DRV19RPYwQnjr96PR6M59xYOR
AFwARqw4gBmxjqT56/baAUn/yPM1ulq5cmdvMb5OxXZoR4KlCf2lImkXhZk49yqPxj+3K+6oxzeU
KjpEZQycsh/3BfPNkFzTPoKj6D9Bq6eHqRgecN0A3znwuKMQcgXh3H3cWMB1VjRkZ3BhEJtN/t84
2VdXjHu4kRlCfnPLYM7uHo2FV1FqzDGwUmdv90mWJjlTwivt5KTxJDsBptxHiAjo2TBQjjLcxAKp
npGQfEXNfOsOSfsUnDLnSKeV9nAWcVbGrpYLVzCKwZXtH0muq8WjO+JRC6mMEaxigL4oH03XVgH5
6xe7q1N2i2oGBqhJEwVdBRk7jLgAxmmXAMbQiyYuxxfn6Bpk18duwDgtQMRpNUluDSHG6PQCsKp/
PgXg5oozQ3SN+6coUIu0UaFfmJ4FatD/FCMXoNzLoZ/fmItfPEsvyGd+cnC+ou4EUtGXLra2n1xz
u4xCTsGPPq45tdL6+zlqJdav862D5xnJ5oZvhprIXNdp9QCmLd/nZlbfHF9/rFgj+tqsoFRdHoU+
HVvi4kN1R9YBPN+2v4gaXkYEga8fzgM13rpNmjsaJ22OM9bqcLeepm7PMzE1BGwDizv+18pR8j9Y
PUTiFVl7UUkA+tHpaiQV1oCjSH93Wr0YHp6Zoct+o0cwcJnrAUpflgN2XJShAd66gNEzR3R6Cua/
EWLc0z6uaZ9rkrB45NI/T08p+9mlcJsBo/TJLPjpe/EnQeTtR25ElHbhn2P+6eGpr8ucF/yoOKsY
06Yw6h/ka7cWtrdFtNsIfWlXaGocsQqVnQycEQtFi8KrOjeNWwp4MJV8gv7A7+2uNTT9tW29Z1iz
8sw3XXF37B+ATHMVke6+pFBoswBX0RYLgGUg+BS0dvE8d6ZVDWfidbduS6aWDlA8mhSNw3sYAgjZ
KyfrWPdxsDDBl9YqQnmB5h8Ygz5eunLQfcWpv9IO0m12wNhWUWiv9MyZ5l7G2y8axBbkBmYhRG3L
pp9Mjzp5N70kCDB7j01jwfHl9szuARGGOm1GGowkYhjnLEA1ZN4UJUSoKLnLtWjAEYx+y9S6Wa4d
8hOiC8VzfbW8RphcBKxyWJTo+B0BrEtOUE/dw7my1hDj3cXihRnNN58T+YLNkiLsfZB/ckuS88aW
KUGPIau/aHMK4S+t4hoapoo5nVWVBWPcnNQc5eYKhQbUDpZUwSGalQPrLOwn0t77+fTiq829YtiY
AnbQPhJUuvCwKdDAdlbH6IB4OnS3gGH4+k1Lq0hCA6590G+X1anwA2qIL7cLPaaD+SO3T+Z1pbxu
mFohJ5+62tvPhO4QMEQWRo1LDdK4Lq49kPv+7PvF6ZYlkxA040fFLU9gFcJAUdjs91HYIn9UdYCF
WT4kwFq8ap1uUjeXMEZxJSbJRdKP1hnQoL7hejLaLDKjdqfm8WFU2M/+UP8bUo63x+q9dZ3i2L/9
NTPVl5hOMQxUNU5PiBaakzd2rE7d3N9kH53Hbc3uq0y/ItM0WEhTJikxRydsJUm0rO55DBJDENBY
jsdDHl9FzZ8vYFoAOpa9pzcNn/WI4iTEhyE2rWVywJgEofQ6UGo+8BYHQBjH9HcpYc4Nm1Rn0Ehh
sApbAfCnj11dfocsKwX6g1HbqrQe7+reRDf4w36HJl2yJlUJ65ooOky5MMFXcjqKnhOwZiG3Xkhh
grpI2itXibauGVJvFEgOPb93K67CT2rAwhcpaCWtltzQ4Q+JeBbjI3MV95Zf2K7q9HfYkdKZ8Xzc
c/B+h6db9S+2JSsBA1Bc502akad7IQO43NQyjG7wsP6ZgEs3JJIAfwObN2sVDnQBDtC5wdts4RtN
LajHxO0+pS+sQDrBuD2s1XFoN0m0isjCXR6NDUPH0xppjIxJEbgO0bIDH4a2QRuKPuNAKEM2b5fh
Dp2kH+kP6CTK/0pstQYpZlTLUH/IkpBqH8/SUZBuu/dNZRLOHG+KXVG2PeD/d1aPkuGa7hQCtZ4e
qg2rKziRt4QH+mZskGyJ9aDqw2slpmFWNOJpN8T+0SouVDaJI3IxuZi9GdhSirpQ1MySFAFgqvCS
cvzXsqx/pVHg5X0meYwhSFDeRmh95wyPwxph82vKkHtf2lxebr7T7mqF7+M4/XeSstN1WCB1WAWW
MaqsIt8qdOXIIEi7GnelFmlvyRC/sqWBahlrzQksbdgsbxW5clypD5GuHXcpL/dUQRRewXV32NKa
0EfSS2/5QmqdNb1RxaAOOHI13j3CNtyCFqprh/KFSaxd6FuRabtrwB9lT+9JEBT7nRJWIl3emw1o
8tuxdob6kHely3YO1FuTw6JxIfGEPsaKxO0u28ZmQrCbQ4cAzbqQ56IijPxJ8OMPX8EcuQfpI56P
dkorBy/JcSaW9Dxg3GsJhf4Mqqp+p78rMLRalwcl8jkj4FSATfFb5HZn88qeDgjXyqSWFBOf930o
hHDUxSmi7VmlKt23W9X3IXiZd9aWirL+DE/K/TgXoZ+8JC3nYmFonot8PMOGd8qGpNh5f7Us3Ku2
NkZ8LdZMIzJDNaBtdxoQ+bB8NKiiyrf4aAkmBzhU6xxzudeaQUy4QVbLKk1EEc0+r6TNmdmw7FAM
yjvzRZ/hKYYg8yveHucPyxOFz7gz7KlWHEnx6BIgCARkZavvS7P+VtQgXj4ciASbG/9Y2oBFPUtU
huXUHGI+6iKyUE3L1z0grOCDhmN5YAhQWkeoZ8WF2kPjwK+x8i6ZqTnOccOo53OpZujL3+13tzQ8
jeUBtirBpR+6e+GPYmIoJjz3Fpa56ypuNnZ6NarAtX6ewAQwsn108+w7foL6EgJrPmJW0omhZ1d/
o3ccXUuQNk2yDHfezGBrEP7n9q7tFyNSJSkMRj3BFeKzi9gKWGGsfZq38+X8KpApggih3L0yDg+8
4AiYTWNnxWW8+jk92S1iJryz6qYjYbiKW0IqNIPcRdjjNcIDew/UJw8VghkWgEQuRzxj81P0ZKVR
1NyXIDml5qmYcZuPSYlbjxWV/bJzEPoKHmzGdrhik3ap8RNAC38FA/uUtPA45tCN7MmjFObCkz5g
BIeW+mM/IZrvDPK7j7flmUCO9rp5muCrnA1kjpRo49ahWK7AW+AAztuz4g1x5tm1JTUrWU+rJOA6
mKRML9OBDY4UkF8rR5t+YHVOUuv/xzxedd/clkPXEwPxaKbTo+Qdhor4tAOe1heI8i+2C9vbJBwC
EtRQI+gfSdjKphMH3FWGVT1WBQSX0xk3XvpYxbE3yOiI07G4wBGeb258zV5CUsToRcs2Skx7UNvI
uSvxbkDp1psWJ1EfmkTaueSJ6Nw0BkqdNRusp8NSfrjMTotjoomNYhm1CsycRZbXnpi9qGD5ZQFO
BnI8dwakJfJSJaHU9fgNgRaUbPU0l6kQfq4xaFH9rJISg7sXGDgpm7HBz2ltmTPvSi1YOQXNcnXo
3Qa+RRwfCUAiKkxEOW4rfMDNY4i3k/Ts7DNFmHz5Uvn3QSnziMEPDOR86feMy+INeXbYC/cOrfr/
KR5moHwbmEDK/XPtbwrURngfYR2ip4zxjRHE2CCruKGj+eeszyOvwbADerEtAzNGKGhwbcHBPuS1
3Nz2rRixHdZLFyKgWZzpiib5NK+/fGUb22Ev1A5bja6huof8QZqLRfSKMulRta02IBmqaexQAzHm
JERgB0nAVxKHj8EVXtj4m0zZw7vbkaNDAE497GOnkYJuf8HC4oPlo6/r6vroD4V5cGphuw801Pe6
FAp4Es3s6RhFIOK0jIPPtO5+xhMyHDbzjwDe4uZNwoe7oiKa7Ta2dN2LZIOMXT0zPhwuENlfAPce
OWwlNKUo3eMeuds8E0JftIKt+TAD1h73FDei0DqQaumWYYRWHNuPlG1S8I2Pu0toS9sUFU3l2dE/
Tv2dqDe25jRB7la26fzugq0qGzKJSdN6dMKGtADZgmEIJVhgjKvJCue/6WRF1w8YiDvboZgHQEx0
DcbbciN6m1ZjQH+sb70e4+WquFwNyNjLG68EEsQA38a6JNi8avmVtHfGHe+WXfEWJLKPuvVcvd7f
IiHPrJl4JgwtcgMfJJwxoPPrImx5DT6hxKQinUDLPJj0bXYlz4UhhC3CtZ6xJU5PRohjqHLYjc5P
HUMK9VygfJyWjTyW1xay8xzUSdmwRhR42syl/65fZYxi1hjwPt4iAMYuuBuV+EJ7WLjXzHimwDMA
t9/9xX6EtzcIARexSQGt78Fl1a/VwcenDyjhlPLdvhoDDdZKlwPFGxSPJca1Wme2uGgOBiGQdjqZ
dFas0LE066NHYDJM3BeRqR1Tw1wtWGuiVz+QvSep8/hZ95Oh9Jvqr+Knr0AUncNRCsWGT+aZSOLy
6e3wgo8bWDF8OjMKrJpysYelY9SaOKREn5iiBZ4laDLV18p4WfYFdbHf00oZ6Viv4OwcR69nxL7g
qdQYZiFTyez+DfaeeKp5ejbO963ot6BkqNBfbKE+5tCPxWHANgisfUQcH24qiD7O2hB5OfkD0zv5
VjLmLDye/v8wtGRIvGWCW3P0zzPyjRSwS6pMzTjYA3VNyzIvthlFeGCcxBQFpTlgp8zAWungTt/Y
pXK4jhjTp4qVH5EMF7Qns5w2e69K8OCStL+VLZbZaYheGO4MhNKnBYTKkO6IgRfhDWu4kRpVBNwA
Q8s2p6BqPbI4wCRahQfRSK1ojfV6qS3hF+R1GNjH/L/TVBL2bfUBzh/2bf25JU+BcPU02zWZEi/i
1TEA57OEr/UwGQmycYnhVZ3DozVPqg1QxFSJkuvJWVjYbKvHbpWcySIxfkCrqrndG8hdp9911tn1
U434UIpBrwsBDX6/j6jU9MrFZkTu9LpIdP52CTaiWb2bu9uqbC1CrQz99SGe6Ahv1KN/923DVER1
s/AtWE0A5PlAksg7iTmQLQ71THBVUPpWeGYv0yYYEciCtLUtl5lPeE07OeqtiYBakzkZ4BEDF325
1T6qutxknwldOpO06t1Ap8JathIAcUJfMrcgcSJT68Mq2pkJ4fcggqW+/lMTciKxWgr4PrsJD7dI
SA4OaEL38wenNBAQ9wa0uOs7ViLWpRJqMWhOVSec/sLV9zi7QBbJR5Ba1+2B+SJwVmZNUEttlvbt
NnGSjrEeeI615OQ7mHH1zn1fWkV/ImWZm06quDZOvXWV7p45nMO4LxhokFMpLfgFH29M8deg2Vk0
qnK1+fGOwKsqa8IH3srX57BEwhd1BqI5c4DvzUjzkv7edeZMGS3JOrKkBlBYcLQ/02R0Jo34271M
lckRhKkteJaV6uP2qnbwrWtmzbl0hEJ2OLdoQvGhXzFvz/qBi+zX2wZSeZUzgd3IDUzLdtCDQomO
cIWv9JVGnHTQrmIkDIzb9GUoet4kcIIyRkZkrdTMzAnSIT1eJEMF3lyaiRNF/aGnEpMmvtF+vhdm
AD7PdGxV+L1L2egVXcuHBFjAPMQYWS6hSXJsrhyiLR3Lmi8WMz+m+Hp0cWeUu+St9sYUfkl7riqT
CZ8TCFi1yIBSf24AB5a0ZlkeZHGjzAXcLd69L8Um50fzdqy5k/8ZHNdNFbJRB5DRDNELDf3Mt1Wc
O5J4xiihuAOKXZNozDpBH1BFp/nNvrH9Yaj0GhAJ/cvvOssjDuawBecbNBXdh2D5rTh2Vfso3Y0f
eZmbplSPcCdYEZjraV/e5NlQrHmbhAf9Uw3vqfz6Ct+T/Ipi+BFkPPKKvqfoWKZexIJ8PTYVXUWr
9D7wa+lEgOJgGsHnsdqY3R+KLsdoNwd5WGS9towReTFAjtHHRQGklq/j3v0E3Lip5hwPdyWL3IO4
Zk+jhD98m+VFpkaGYKfgO2jqOFDe7wFBzAaQAi5n+VNdpQNcgYChE9H66DRn/WyxcHLZi9BalTIb
mae/0us6Ydt7cU/i1v4Y48TQ3g6rkFb8XhORCW7ucDHRCdlC8FyRoYfC3dQvK5GBx2vjQZuRbI+p
PVDl9Uv0i6FJVYNHteCtToYiwhGuKyEyJDYRu8jjf46RBmGubPN6wTbQsijkQbMEvf7LjoTOyipB
F3m4dtMAds/G6y/HQ2rH3k+MmsJs0dTION/yQUASJib2aked3CYWMS/63w7J7EDHZPjjXwUmRnzN
MtWYkf3G+/3TCxphVa6Zra7X9ksJLLmS/kq/l0WiG8/Wd9oefN0hk+NcjNxr0cNYonPhus+LkuZl
VJM3JD3qYrdgR5z5qzAPXCiQTtke8PRZQBoJPqrT/8TLAxb5wpCVFBlyHzb3TRcHFCMw8DqsgEuu
wIhHzbilOHR8snrVk2KkhgUjV3+/AXCmPxi1Pfo8ZYFRVIBipQc0qmE5q/MpTDb4YRzvq2odREKD
g3ebelzlOuzzp00JnzL8iXW5ZikUOdZ+g6Rv266Lym/gSoSjgWOXgjYpF79hYR4GRdCLqlRgXk5x
GArqtSdHP73Ae8xGTlys0ZNcCGy0zsvdw34HFDgwGk+QZmzXzERruSp7Php301pczNsZT6YoX4hd
G9htTEBAIVrwnFzvvhHOMevtyVfWuemUMcHzxFvhnZ+GMeDd2qQfG0PaAcI4Gi/g1ITKTOmkMD/n
JOM+5Z7xi/b6vDNbrEHt4+AEJbF1oEt0Vrd7+PVo2Tu/V7TzG0yRqXVSZR25KQQrLe525mDEOsXp
fiWW/sqPsc+s7rpMhEDSIjUpZRiSGCNBdfvq7EX6qXDc72kxI8Pz4FkiAvJjaKnf6pPwtRJdEpL8
uc/YIiJ+FNoMxF7FETx5D6Z4hcukbUPJP+VMx1P9hR9sVPoN+NTv1C6xe9t+R/Kf72j9jGg43DNf
FB0zfJqPWm3rEYJ+9ss7Sa0kneW5ReEnri5LP5uKB37jjJ7kf7X4tsjwSwe84FL/nLr3SBDUaaHP
4yvfz3RD7EPl/CkN8ijHLMyJVsyovjEbWGf+dPrMDLX9e3gmVyVM5PJjtA6unm7HKpcC1FohmRqW
kbp1PRjh4hT7bH5NdDcdRr0Ci0evvo/XQBJ2CzNXvhfCMFhdbdiRSHBfUops8azPJ7umwYK4R595
IDACI4Muy+EZtsrLkokHN1fXlvAUsbs06x4wu0Jir9QQuOM1Pb5eNQ/Tt+4/Hc0ymohA1nHL+oym
OfIrCOEX8pc64MhgqTm3XFChryQvYfbh3F25wpyhsnvbINa0+YRY+nFwVqwRgKo4fRS2oL7pc3ty
4jx99gAlwurR4UaC5Iw/zFBHDthDUwkcn3x0w+Cx/ML+citZJboE2qwN9D9QQEfhT2agiUh6ZdtC
2vK4xViuF2CmNbcIwiLjyJnofZAtPQ0XI8vSYmIcVOiJcGatqNhKSrWxp8jhDrQ2dVMfbf0mst8E
S3pNcAXVpc1MxF0eKQA0sv9P2DPpYoSetZgz6HoUg7l5m7O0h0fwTXRAT/Xg+Pk7qb1z7ULiOiGo
AhCXeQlmCcs3C2mY7t5rlKUGHbLyiIooipMWAuw/hotknQXk/PVjYPY5J/JmK2agjTxtfAeyfJUs
ISOXVrYwzfWki63kgFVxPrgqTMnDrjL5UEjD8fnFDvMmNPUyD5lng0WrwFkPW8o6pOvTsqHfGlc8
VSjevEdFERDtMpvsX1ECKQYMJAgVgd1JW7+6WGq1Le32mhhWnN3t4O9QjBf/qdp1EM3Kf0Pr/Lvm
9Q1zp3dxizzbzpYcNFbwOcQGVGmOdte9vJl6F9lTZiijlh7wnxQEvtghDfs/N9tPDgY02gD5my07
C0jTLaeBsehMuu/WI5RvEJVH9f+6Jo01BREtmk9WayOQDq2BrSYNfMflSNwV5sYltmHNBzkI438B
SC4I91XTlGZVIWhJTnTWBVd/F3x65E95IqfQCntYgE8QPQywgRNMhybdonaWAkgmyZ8cJjt/gn98
GGiXgkeLTIXPbou98qXFQSWpe8XXJZb0KfKuaE/gocMKg1dRMsnhYyUu/FJgnZzv4qVVb6lvbccu
3Vslv4/MTVp3D38NMqE6vXMz1agOZ61D/sUm8ovAnZ7xS+mZ1uKAJE+tFFmfDUIcLyO2gDnvWji/
E3XbYLScQj4UGB9sXfEyLpZKeZmKBMxxlUvQZyg8JzaKF6AsmyHEOy02coeX/jxwPZsX05x3gvsK
GHeXAkfOT9awdYfHW0rdNFBaoRLmBbeMVgarQriiQPXxl/kK8B5xY3DYRYr6SjKMqhgesUgCuDep
vJQX8yigctKIaAjKN+McHrP4GvPxWmxe1ssLL/b+Or9/dNiHo/3mdiXdUIFB/VGtCeCnA48M5i6t
OeE2Ot/CpQm9M+xG/ypgqa+tlm/7HfPWZQLMIIL8XURE0J7Ooy5/0widu1lv6JWs5viduqSEvqGm
ZGWGpm1tOEff4NYvupFgk6dwcLCmJ1H6X4A7lwzhKFtDjUOL7lW8nUjSVGFAjycioBkubt9mR0zt
Df6Ym9q6c8weead0apgHtennjEWXEbA+wKlcdE6zPKqfZO80Hdnqh2Da7EFgsJ0IBzriar3mVLDi
Zvy+4yaGNsMMXZiWUF08QWpA5zKGR5WP8suVkSqAE28MFEPAi51rUEPXoKiuCnA1JrZOCH+H0f9h
P3iFCQvPbW0JkSzSTo61YBiIVaAusVu0+ihzwtpBjMXon9NpEwI31choqzlmyz9FfyGRy9seFHZC
U8YUTKtm9bcFcRzAO9wmY2t02eSERu3PYXOccas2VkC18IcLr3M/H57m/oTX/v9mku9hw5iCEAFK
PY68Buz5Zz3cEvI/Uy0um0/H+hWKeFvcVVyfaD9sJqkY/3zncGufGbF0xxh3aqSZXkmnGj9Rq/yv
5Tn7BLZZpLdtKfbTzVXox8REas9mcB0Fda7cv7j3oa6TvPnvawwpv3YmlNU6/T3rQksNflYHt7n0
2lIzuSG19jf620iAyKRAl89JJBp+aVWoHTIggvSIFLt6LbCKQCUfNMn3X2TYszaPOkhs4sesJQri
QQSui5WMvjHzeG3323u44PZ9gKaXbOSFxi89twO9XaDGOeFJRhfootnb9KEl45ysQyBYdlLL2eYo
L9w3hFI39O8XJbzWTKxyOCdUXqq7vZI1HgJ0Xno+qvKWkBS+ab6WkqkV69g7W2chtDmocAdJ7yZC
Aa2b3dwE24qeongFP3aUEkgdvMjMBoFXjNTJviYJFS0Axg7N4czAAuVxZihTcX7zL+Xiliqgmd18
mZpCS+3PwPXUWVqcO0lPIt0RsH+EgibYoN+L4ICYhWKRauK6nXwNpj25AFDescDwaS2httQDMFMN
a6IRC4ztm6zl5Dsd/AhptQ2k5lzvMfZp3SoyVTGw2IhbnhnkLc0+8cbQANCylfnTI6Mub/W8KwBg
5uDUVrdeOmv8l63J8lKgxjCZF05QrpeCEwZDXYUT1jWkyUfVgpnkifAqYSllGL1qPUyck23LN+jh
zu0IxGsvBGi9Rf2gz8h5fiJwNv4qV+iv3CWBcIda8K/RoKO3UPKaM4Iwhlk2QH0xfh/dLs5gbU/X
nCZ75hazKG2D04x+V8E67AEMmjTjacJiCn2OiLNORoPfa8W+VwpDPkfT5PTM3JPuHvXoSV5snOYL
h3edlAF6QHMVKMyVNN909n/ujcOKue1vmGgrSJVC02zkWFQ1ha+dDp9RgrO/CgaJl22BV0HI+Eql
GyWhKPCECl18Gdb4QiK0XTN4cPriI5ZnWojdsaqOxFv4a1aqpRG/POPTJedqHkO/b3cKnmRIWzp9
Pf0wVvavOzSXGVlMINKWPDprKZNDbpAqUSxCqFk5BxQF50DCVHs8DsCA7HeHyYdXHS435PoTKT35
NPpUq9uatycCcVzKzATrR3M7vQk6LS9z8mon8a46tdM8exhJSYlrtRQUbtA2I5VCcryV+i7xKHx4
1XZrAJ2l9DFOZuSiegggADnxz7y0ww52fVCd7f6M0/InKok2evRMDzPVXGiNQGFXrOBEEj6VBjIb
zGenL26jWHGWWsgtY0hgBMdVa/UKExR68H6OQE9HETBeSNz9y+NGJnKtTMmwdskPc6x0ipbmg7Z6
YR6W6lT9QjggjR+Uv5SjTUktUTSYvHcwwTRr1vLSTGzDVrtZn6JrBgT4Lax0IeC4/s4jseOdK++v
y6yvCHRKTdDtXpqkr8JYnpV9KAPubouhshMG4Fb8h8gQKY0kGAfb7tu0sOaPdZudqtfcRKzc9OJL
PIDXv3Hs3mZaYz1auqzQmkdFVbQIrZYVK/t0Y/VAtpSdwaF+ff9BI1j68YGj/Z4dmokIhjWIDoyx
WH2OVlgu5NHpaF9xF1qzS3NhAIHqWtfWs6JSxTb8iYKNU8aBzyra0k4UFg7XRJakpdZkiNraokq9
VAIMfKgwltQ7BOeeZ/rImH/i1ltoO8/6RebYHtMa35ggmqGwW4h5+j/iH7joggj4t3m4SygRB2gd
MQN7GTq+Pk6EyO/B4WdR/jRU1/DqE/2BS+t0c4KrTqclyc3z0yiZI9uQe9Vn6PGTlZ9XH6dtAeCG
FC7F7DVZMiRlRjTAZ8bHG78AJXgAxz+UXPKPqA3OyXRNKYORClN7Pqgr5JeFqymtM/MjhsIM6jAH
SZKSxoEZhSaWCflX1tkLfBy1LmKDcFk7cCXNV1kXPspMYASN+0MeDmGzsB8h4CaeYNLEuJ3alxGR
5QgARPjw3yJMcbdCIF4vT61hAo+m9GVEANj4PYLi5Tol/Hc0JjZ31s7G+AhtT0NnhZAGQ8P8NYmQ
yIywxqqQl6Q4XIi092CNfLOmHDpHIYv6BqbOKGHkgRRXan6AkxsRKRzC+KtCXJFXi7ZD5e/on+FU
3czeZUIekoYF0yGJtqeoquXIA/9LjGfy64G2YGOZOXO4bQt26ficANxPNFUWWPFBwPWn6C5KRjcN
xSBCWwfSWAouJJ+L3udO4sWkbHqdEW2JlJmLvcLnM8/8+BdP9FtaGshZGT9NV/HbIdBrd/7w3p+T
oOXmm6wRGtUDlSEUXl5bJQ1/em0HD9dmzphrGA6FUDXHHdLPUSbxrYkn7KdXtGLZ8Ya0PV6n6LEd
2YDLSDHJrMW6Tsj9jRcRPJDN0raJ509yXBd4+10opHlo5ZNFSsdthyH2pmSrI2MlNQKS49jVVblk
R1njrS1kVIUxRfWCbIwRC6PLiPwfmmriI6NBV6woicINJ1ql6I7IjmBrVzn80ul/Zmr4vaRjd0WM
UA5OTpRoeQF0RoAhzfgkJ6XgUTu0MN8NJ+L9G/rNuQcqRCpgjWN8vC4Vdgiy5Cnl2V9mI4CmZUhE
/OLK6mKn5API67WSTISLXG4m0voyF9C40wq6Ugw+MZ5zJDDX/Q6APDbWKf4PYmqYgNCzcEOITNmW
Uw9DPiY9iWBXAI5vn2fqAfEXaZhSU/XW/EF66g6bxNVa9A5me3S77fy3icHIq6F9CyW/SNNx6b6a
5foyJlbcvZsoL5b7xr81oG6PWo9t3xabL86YkMy6A5Y8NWSMz/mGQSyzW1l5xnC035h39XNJzirr
gfA6CXmQtgW3kzQCxqSewMM2lA2fGYhVWZZ4kywzVfvZbAuMC/8BK3/LC3cAKHSK9ybzKl3qij//
67K9+yzqKN3sR0fKeNh6Dw2vAiv8zG13LkCkJG8BTLhz0DH0ysAEJY7C3lBhw7CHQRC50avWamKL
DVCXYzRaTtS73hLE/L5leCEIc+6S/vhP1HK1O+CVqw9EzUW81SatO0bdDpXKSjxVDgIFzfFBuiKn
8Ljy/x6YhtR/6o66IOo0A62MjF2J4yS5EDWj+x0QeDV/ENBh7m72Kb1P9ExqyEaDEY6jtr0a4vr3
UjJujHdPwMoCkzgr108RmAzYOoJjoqpQrM3GSWE1tLSNYKTuwYuddMvauM8vEYkQPxxaboMAmvGM
5qkuqnTunE4z0qNR+9wRGRk/FnugL3PYYi4NfyWxEiZFolPbMGqEQ7c9ktufx49Rr+KXcVvsYeUk
L5d8y+TGo4qRN7OuPubvmCDG1DPYBGyQ4lnNdinpnlHszhFBKDel1cYujgo05NPtbaTrj7wXuAnJ
BPcW66eT3Dw249b9IJrBMaouK852OgmnkIZjS43IFq1YSRiMBom+ipRcOujZi5zdKO9/PpEE9JZt
RVkYr2lC5FODxQiGqp6Q4A3N2pvNM5nNTKG9TpefzhTe30dJn6yu6WGzhUnZp+SIAfGmcoyCKJJj
P+fGUzW3QypoD8gH/0+okBAUqNI6D6v8CyWa/cfYaOmQmZ1XCFjcU/DwR/BaUeYvaJ/mjKz3yLmr
+HbfSmHlqLPiq1Xj+UXjaXh+y7APvUYSh+SlW4eEolwxvXSchMauNEh7XSsN3C9hnf7ltcaoLvLE
hfSfUDfCwLXB+0o4+qwZ+HDoiPE/DJw/MBJ+uFkfHse5x3rPBjBr8xVRMfJ5rJEYfFGRG5xGVpao
A4ChBjg8w6dXQizs0Jh+foVXOPc4AWWB8ETUyA9hvKN8U/wM8TwaxiC3zMb/zPy+h/vuQJNyc/m0
jpCv4fPRvVRoKZoxfJzLzAYiLBl2H1ObDdiJSaXnnOrBOHSznasmLsMPIEklL1OLTd0scRlzSqpP
B8dAxvH0L3eLpajG3cXm8hU0J2pYaW3JdYyP27T5GfGLqIx9fkxDv3Lsyrinytfb05A0Sbc57/Dj
yVKroaP6PlANkyPSYVTvCTYygDJkwHcOEaXa+tjizFw7ZU3x2O7OPo8pugwxa/h54CRlRbHB/B1k
wiXa57YlZ1VRaMGZb6nh1/GaHN85MSE1rQ4DuKe9a2dnicO2T4kCse6EQO+mmrdI9itEwI8uI8nQ
/KLnR/t6FaUztrtTgk5ZgbEgODFzZXC+8VN5tr+UK5KcjhdYGC68Z1kwg4eUJ2Q+E2BlN9oiSqHW
CbzTCNqv8ByFJdhZKptPaMPKvl63sU7dKqpJXtmMO/inygtXdMXohA7qnhixbq9wZRv+vT4H4keA
DGa8JN4FmEYpunmo+Vq86xKI2N66dzTc18DCijQh24McfHckT5WgSujUvVCzC79Mg4sHUDJWKugz
U+yaUhgBVmlqU8DTBcFh3ZxU3tr6Ynl4cCC5Qfhmzzjhlh8iGTjuOMxVr8L94X2XBFNsXCNwbnNV
dhmPOxhdhrJLPk7cqYLlXmmoz37M8H7U9sYJbXV+18sSdH9TjlmLcT0MW5GuOQsKvJspmfNSGCCh
4t4mdwJMd3GiFs1VshI6ZJT0kxObzU0drZAmfn9+mdx5mOYyI31y9e6cjz3EXOz3sRoqRop/h2b2
jlkcf6W49c/GgCifqWOsxeD7XQESMU2uhY4uqj78ALi5UhSnpqOGiLm8jw4n/WrqdwK/zHwO9jDi
bVahtT3e7POxlXBEUxE2XJW5XE5T8SX7V1vzuRr/PVOz+JdRuzmvdKoBPVHtoaDmTW6E+brSKueN
MHpRs71zP6MUgC+UW9Xp4/WWGtkjptM6teSdgYoQ70CTbGHgRCHKS74su2Jo6yYq3Qh4ioE4srZd
1DnVnn2Ts5/LeTwjkHk05bfrnIvAVhlpcV0ZZVmPbMewGLbyQM5sdE9wpZjedxkf1EUHAVGOPCk0
ooOECz2pLIdd8IKVSdFqWi6b8LkW3W2xJ/q1sRAFe8iUdeP4HLfyL2+TcG41xNBQogico3RXsKhW
C103oR9Zm2kSe2KF/AODG0/JhAmYeRW3tmXzDIFme6ugmqzxrHjesTiierKMiveQHTsquOsqLaSj
insXPrNfaVaEIYBM57DRa6TJ+StGuiBxFYoau4VfEL0CNzgNTxNcXzrfhS8eVzohzvrcQA3BrCAx
zU6IFg1+mS1qu8subtdUu0K7pNI5FNKVtTVCGR/E6SJ+UQf7ArYhZbFTkVI9p0O84zweRZIXkj41
1c2nsRZ/xnDVcNk+CxBl+RDgAH4ZYnBi3UBHTglx31Cj76vLtF1z7ek8v69ijiiH4WpFXRHErFMK
6CxHd456vZhJn0Kfs/AbZI0RBK+k6486y9qQ0zT32GZ+HIE3ghXr2SsCX3FuBHqBCKLO5xZbDk1S
dWDLv45yQexYSG0RFbizcjm2FzgUDVRu9qcBKpGyyc+KOloCG6sEr0qABm4hGBKuWZXOBYeVPree
3sxe9Cj4jBJJBoGEoyZDVscs6Ktf2ubZ/kpoJ0GRLigXiCHaw16OiAA4TX3qXjohwMzKobszcQll
E8QjbsmhOPXY0sUV02Gz5dwyIYdhzgS7R5Ke9WvSz4vvKOrTjkPiNsOwVNibzBT4StH1buKgc64r
2nPtNfA3Xglq648jZepcEUsUZGpuOqRsvViYy5pVh5tyoCD6uIA4Rp/SRrRQyMXcUPUhgfLrq3RI
r4Zdv+JrScwYKsaNmfqe7gTNYyAQI+odWbYfmsIWvdsbXbCUT1Iy7aqaNxOc7bM9dvOe96p+X+Kr
e+uwGri61h0ayVWzDmTpHbfXAbHUmX0NNm3KqfUZXatYp7a1kb5eb+OQ78pyqVXCA2wcXbcISgOp
53RVG+2LiAhmi1N6nr6mh3FzQU2dzxYPk1XqTjoZ4xfp6EvHD7bFw+COHg2RzBE8pFnjJvVMn8LE
cxe2zpBbPm3g1jT1SolKAHbElZtpZh+i3Ss/ljRob20DF4s/BqmtgVqTL2Gk8MmPUyHFMpnw2QAa
OYb9u7tDfN/W4L2ga/GFv35i1Qyt+GiTH6i2JqH0fLW8M4+5hrYBxI5ScsYN3bQCOxGRgtK+TwW3
71aSSJgYh00oI2dNtmNzV/XeA0SLPKknIIe2O9u/h1ioZhKI9G42oyJe+F122u/MDyn8sEd3m3jy
CCo0DkyaQPV7fqfmyMuYEi7OOCcO/IJKkTRiv3Ov8ivR0xWVCV6x3Kshdr21ahPEM7hcvW+IfHJp
mDlrlzxFW9brZ2h+Y9foq5t/ZrDRm8tzyuXPXzaxka3f+bYDuR9XVX6Ieaz2kiq3p57n3XiGYF6M
2enIaG8ktXTKxTuV0MyLOdVUHAywfgy3KfL791PnUDwQgT4KUQNOqehONGJTxLAf8PqsCH2x6QKx
FmuAa/DWSh8z1nrelEiD5+0EqWDB9K3CWdEHHeiUQGDwyjYHGpCfHhiOnTR7a3QX6E/UXKPhimu2
WWu6L4id6+OMomrCVq2NEfn2Po2VvYC2zL1YOIk4O/w68GPJvF/5/w1Q9hBODgpUb+ZLp6mzlKMx
cM++wyYV9Bm1MhKsxbykdBbEZS1wrEG0PZ7ls+8nLnsGlEMf3z/vtMtUosjGbVGzzh9LWpZx3yfl
NdwAf37YPFydfvfPcvnwRtijAQDJ19l+Idlv0GcSmKs9da09cF2D2Uj9crYR2ADB6wJSPHLzVtxq
jRlVJ5H4QznUyiLNz66zvPsJ8Adpr+xg3Klw315VeLlVCyo+QYtpDOz2pDo+u3rP7pBbtRaOdI4/
XkzuvRhG92U1vLuJ5qMkV0cAQrDZqs+SnW+T+n0qMPlAf5APIFmucFW2pUGAwBzlPJP24chG1Y6c
fXtjsVaeqpOHXuhCbBuwnMWUfq25FaJyrXFEKTEqD1/kdvQ4+Vn8/AFyOeeYvSRVpV/TUXMoP0Ho
oBlaTC9s6MZ27i/5TsGos5pNEtpw2RfdkxwNLX+6LcT5lrniY6BTfxf0ZSErB3ZVvEA14BZ5T4rA
kyh1Lb9UoI3Pq/MlzV5NVu0b3pQvnqVWkESfFSE1IiX4l7m2athSmPVUC0A/q1Q78ZW+Y/OCPFk8
YxlH7rgv/257H5tnXPQxAv3BMlj2Y41aBHpmyEnZA3ErSRmNhA1GxIOve5vNuOkQdy68KBS3NRq0
FJ9umV8PIgd5qdr4C/m0dKNk0/t8vzkqJRFfhgN3ODZpJ2/4KNvVQOnuGDfdBKbHV9t4IDv0Vcla
S+YriNaednLvGqAcbJh1bVmMrTSywefgk+Yxf9g9kXr8MLRWUFkcQ+SS8WSvYWZF5kq8XFMyHwRN
N5PYQJkmlzY3rHHV8+PwNGLdcuttj/7nuJRUHdP+l2Pwfx/VW+nONgaQRBs+XewOyAAZAF1LoK/R
Xj2qhAZP8yTD2ZhoSC1UTGTGCo0e3x4OSDSG16Hob2nyitTpETrN0AQ8ZMD6ZmhyRTJiC5ayHCjt
mVLR1+EDDK015pPssoC/4/4Vzvuflymtr4O6njyulcw9cMWnANTWUM4YBhH59gG0A/erziV18ZUv
PafWBjIcQ9MdxGEj52YsFmvocyS4oT1zaHpE3iIhYzqU70ywgHcPPJ5WN64nR/h6UhnmSvxByrPW
InTg/KXLUCGfCM2ITzytFdKfAnbL19LvNMVl4b8HMwPsw7CDrAsCgaHPZnxsy4iHKB7bmqTO5CwZ
hkP/hplBDcoumWqpn016UI8kxkcPMkuKxL3njTKPlQH58u8YL6VnADtLN12DJ3g3kW2m0bXJtVDa
go40b7ZHgo4ymmUPJndFFbnwe0EGfObbgRoutfqYho6iXaiKrlD3BAF0LK9tuA9H6bxI6oFJY2Ni
Oou/Ev64jG9JYe27SK3lHX68Ia9ZFNUOp+o44pYkngy/+bEy8WPnhcENa/Ae//Nl0y3TNA1jgs8+
yV6o3Yy2VH/U/YXbziorwLhAdxz3Buo0K7xTvRgGxFnUmOo2MCp/TkuDrA2DDUr9yhP3rUwJxbYu
RgYQlW/M4ASNzYIvL0t/IH4nberbrZZKtAeRAFVR6kVCDhmq6abEvrippvMGU6W44c3/5yX0xIsP
aHuA6+tW5P9tTsaPA53rl+X0JSY4E0EMOtA9MTfQ/XVx5i8qmY932mDVMmUpN07GVwOw/Bf2eTrT
36dd3Hhy4DMGXssEixyC3iGJrwoXlURngGOlSVDXLdgos5xbtcFq9bveighz1d2zIdD3K4BuZFLK
PcJEr4HhdvHy6q6vBV8YhuNWe/m5VHFhuL/FLkgGtGZ82y7CYHzPXNd9vpHVPqpoZbEHOFfZ58zR
+XE59OlnF8PhY1aA8hUm+s1fK0OIiZ4Gd769gVJlG0StwsHxX+kwCBRuNm9oY7gVNmjDfonWRywA
iLeCY76IrRpfi1VxaVETPp2jlhzWJhSxWv9sn+tSOn+0luz4d79Ao9bVL94P+mg36KiR054aokeo
rx0bUdchOtUgJUZlNClzCZ/Wz+IHa/cTUny1wCv4Z6y68mQ+tCGZj+qe2ijceJAFmbT1klyuTQ1X
uYwVx+W4im9yVj6JJ7I0pch+sZkOqMv4IHQOQRkjOPsfqtOCmTNqXznxDB4Eaj21gqLnxCXD3ibh
5pIi1rMavxmtCIgDgZEfA+emTZKDzk3pfZHq4+TjsTUjBV3k1bMR78UJaPI+udIsGF1swro1jkJg
RsSioRURSVpcPAM+LiAjqBnGx+imwYkhqxRbw93Q7YLL4zN3WhnqEPdFjmDRI3zyJ8ejfi/kjqMW
VyjKM6n1mr4f661IzWJcqK2TaZMicV0gb2pVhxKN9mFtI0Yu3L7Em8Lb2vxcS2xYiw3V1STeBq5z
/fs7DYl/WXa7ftySjNEGt5qE6KfiTxd8C/KNa2Tn5+iZDYCB8ukq8ei4XBqN9FE/eFIDraAIdPg4
reCCIWuVKCyxV5ESkPIY9PkEoE/OcPN6wnH/aL+rcKrUyhbC/Zlqem1zEvdg3Yfkvwi0bIOTvSn9
iFOm1qMb/qMvwHtR8h7OCZITz2BPOYk9cIXRsfA+RORbQaWG1efo+ypRN/kZCk7g3Z4nrNy4C/2N
NTNtC/qTQWrH9pIN7k37TYxL3rnNE6rV+vTgHnE0rWWUtyVdLZmCrz3Uq2+8rSHZcrQ4PHJBrdLv
aSlqL4JnwHsZv4JAjQdU/3ufPKaW9oP8wpqHXsLNSClOC3YcOJJk8XnL9qTmjdf/1BzjYoIhNAHE
FXyQbjbwXlLbwlWVfCxUBu2Mo8W05GNLv3KBcXGrWV2iMi/U6WXmfEvdT99UsZ7y7NaCemFFZ8T1
J47csk9QwTKl85j6oTDDE0BAEFbOaul/C6jlzv72vcAi0bDkNlamnJMyEN3eYs0Qi3GVomuHkQDt
FOkXamC7r8vil7fKwF1JaTrVgoqzFiAcy7JPcmdUu1a2782KjS28fl3+Sa3upCo0Jyyza8Q9CxzB
cMHzqQQu915OG5ZDwacVuyamQLIGAVH5qem8W4C3sUDXLte2g+zz8xLIAtzdTp418PlzOD425/wR
TUAb5mH+xcFCLR8+sUbFWJ/NMyz8DM04gg5u1hjett5OqfrRpz3gcPI3xslw3NOy/YaS7wjJ9mEY
LPLaav2mVMUcSIXwJ3t4RmDEgJudUz27lfUlfP8+NZjRWVsJYzD12iatq5kQtWVWLyw8btiPNhp/
o01zK/sZwD+ALf0AlsThkq91y5Ivh+aOhPh0mFLg0DsHb6RNhFY9J32hRXNmDEK0u/sAhsrpQnqh
hmZZG7dIKefbdbyAtoRZAZnlD/j3aGuzF22IK/tjCeDexYJRQ9+r4HlUToIERaOUJi+mqvzUzt3x
sri24tr8XJsg5zqYlqw8FCrq6Y6eI3pp+cGFz+i6PapO1vUZ8YcE5ZEYlB7CmJPp0aHIpyZF745S
dz4j2fA4+YTer+6IyT/oNVE3LcjPSFV92ZZ7IJ+R6h1R48bc6Hzno4hCELVAyNxsJPYPCMpFjWqN
8PZgTJutKG86VSze+QxkaP6iKBILiPeVHQ9KPnDLBEnDd0vf37s6kr5eIgLtOvphF9DaTkuy02NH
6czjzaffb5/O8st0dEio0+i8iD3gtUy7q2opxNrrNktDuOJvpbG5RWdlcBUiiRGQI8Uss/DhnTtw
u8NJj5uBc5ePBcx6l6EJgsYNX44l2v7lxmhXf0Wkyk07Iv9Et4QxAkMttpxC9ldWH4ZlJ+iqJYB/
OOZQ9cSbX0R8rTxGg/G1Fkt1qbA55oZfHHJdpUUxjJ7q8ZvhJ/pVd9kRn8kQ4akJcD0kZx+QAfRr
c6Okg48dDwfHx25Inr/ToCbiJ+eP7v+4o/QvLz2hM9KCun2GZY5fprmKG7w1oCB4DU/UszMGMAsg
gqkMkwevlqCliVrCzArLEtAcsOReD9aQoYr0rGdHxgK+e7HYy2QwPGsmVXyigBQdZITpObD0iATM
tajJBp4j/Gw7HOPXDQwL4XeVgvGZAVU6bbYe6Eanwg9hy48geBILmVdRIL3NzITQeNudeogcR3FQ
HTf3Zzf/aRCtIqgCZaaF/q9VThnq2mxaYmH/Idu35K4YU9xmuZO4enAfXufkIMm/QoPlFB6gKO6d
vJpHV8TOh6iLfq+Kl8L+VHtb8zdwnMmee+pshYZ/p+GDqkN80mDv7Tc7WLZzOiLHJRKAvtxLylUr
zuXdOlPWAk6Ke2eKaQzvM4Z+CCHQddz6ZP/ksI+TFV8Yh/K+Yue+FNP+r20cT/yNBpgpaqM8silz
J2RMW9ynPJwd2VPCwf+F1N+Q/RcYoCbnaWRk8UZIF1dhn3trZ3Dic6InV1+KGDQ7pGsn+mv85gA2
ALxUwftVPayid/nar8SNwBP6NPcpQhzPUnQsXu4edgveZyEALV8ZGACKo+Oh1VB+qQX+EgAgn09u
PMuxCR1xHBY5TVnYvJ53+TUY78lKkoxG/A5m3Xm/reJAFCFXXnPoYAf8rKzPC6ohUlWl1EPa57V+
TB7Eob6s3RCFzTx8QlI4mP8ZhpPXSLKrA8LN+g3RFe+qZvXpYuA0D+g+QJbfFvCm/9i6bohwMJ25
Fy8sMu49/wbhqMa3f+S8APKO/xZqxC8+M4U+wDcxHplbCA5wWU7JRPzbds+rRkg8Z4pP1tx6RfDk
0Xe5+ZaHrMyNYSiqpsQZJNZCqtmLCfLuRCUdNmanWkOKfw+iyn9LDqYLs77wC7aZ+a20AMYMycDk
a70d9ECj6cV0gli2veBuFICeEPDh7SyRV9ioQfi+wZ3Rmq0zDGtLsVCiBOxREkCap3+VOUuxvXfv
rGmdCK4cq5UCpGNQ8vemEvEETjIPhWxcy3Gk3cfD+H8bgOWrUCUqQXzNhvSBhxHQoxuROKVDt9HA
IRxLL4h950ZsiCD2ODgn35Ij9+VjNlhWYHCxRLVJY4ZJ0Kn355ZwbBvF1oZHpxJ2tv3Kr9cUhozF
IpctRiF+DiOxtwZ5fB892QZKQ58pnuOgJBdBd18yQfBMLqsmib/oRtEU5lJDCgXa2iDeSOuQQqe9
JDNC7++2Q4I184BLnp+mmPXEk33n20E6vfsiLaRKXxwexZGouexMkOGVUnGBPPcUjA+Jaokpt1GC
9n6PXw04hRU/VWTttHKn2AxR+flbVBB0RI6POkCKPEcaC4rzNuC8qNGh37+MVi0L2KD0z9V9s1Rn
L9lQrEwBrkPPLTvSD+fi06jdFfPfNnnk0HD20dTYCIrjOgCv+0nXaORrlVZP6YODxFga/er0tmKd
eG7Cus5AJ1PPsotW+nhKkFViHTWJWIj2hAiY42zAHZp78WKp/gM8w8yExRtdWaJN4fZ+sp2YccLJ
X5tt6XNXMoE4kcaL4/56uPPYDm4LeIvOqEjqarLtf5F2xo7rAsuCnNgRZCTwhj7SULwbk3rQRzfj
UJGjZwfuLu9tsVaoHus/6ChfVr5J7lRQiEilUdddv6DinyKx0GRoWkTrVDI4cjzDrOB0vuQHipSa
B+Pw1YbQdB8UFbqrOMvk22k8CZmjnSL1s8gocoI3Du60S7NxXeK7fljCdCjk8XQkLmb18V8Qaw8r
wlMYLoT3dbGHDIfrXV0WkPgyWrRKLkpnbd2PZVpGHHI1fnR4CduK8VBFeOt/XYcq01LB0//GT/qR
aJajlfQvgBBvj1bt1If8ZDysQZWyymHWV6oa7d+u3Us3odJWtR/KKUOrDFsmcJ9Tzr1MLRybhpJc
0L65BMSqI4XoSlrV2bWpvv+DmCJaTJm1m63o+NbmSrkf8F2NKivsnj52X2JFVfFANnZ3Wl74bbFA
D75EUl5cuJXp2i/N4LOIUC91NmDkSNS9CVq4uTUbWTMkhNcwRjWtOIJRlD7HMtQfU1bWR3NNHeP9
8mQDCU+zM/hulanB3AHl07Su24G934b4e8+bHBZkun6WU8hwpg6b/u/FDMghCDB1NQ3FdytarWP0
kIBtdEue8odhMFCV9GHXkClghl7ibJWJTfu1LPGqtyp8HctxszUXAKXET2GYktWqLlNoxbcqlE9g
cmTnA7J8cJ7nteOXxvFmtRWtKjH5WiS0NDWT1u0v8UWaud6fu19k6N/SUZpKB2DEb0IGAJApi+IU
28rRo8nE8mwDN6rQUqb033FkeaOWjLhf8ZqFD+aJrV0bAU+MV72DF4SoiYyUnhSwHJkw2WR+vVtK
6eK8kfPGxtoprwra1eWiKv4gHEq4/Hwj2lQA4+iOoo776kKfOTX5uNwGt0NL3U/zRE8YHizjCICS
UYdQvgsqqpvRElNVcE94OSsc8HefvkpTM0Xa7jP5SDGRwATlGp6gdUh2G4O1/IW3HMzrYTHo3ZfF
DFHfoH+Qtt+GgEbnYXb5r7FsSlx0F0xaBrSGyerQgMT9ZaBGDzRBp5fTXMCI2VGYyV2HJ0bZ/YWc
6Vc6+k8mxGtz1xmUCJAO32q+yrQDaweh/QiXLyWbh2DYIv9yWb0N+LCTZ1SP5CLnB5X3nLeTOA8e
sziDAwuf26kGCb1Z7URJE3thGO836Ala4Xv/IvaOljSOvnLqHqqZ97VgDt1KovUSz/loMnPxn0vl
uU3fg0/jzgvmtSoWJg0Mw6F/k1d02lIbttyHBHZoQPknuF0dKR7Rvv4TVZDkq97SWuif9Ar+zz7I
ehrTBaCSXw8ySQh/7U9zFmHP1IIqe0//TI3IzGLhzggV4IXABIHbqFBPZGymc4OABwyHJOxkLcat
lQxjAmSjdIdmBfcT+nfzn8hax5f8Yu9ePLwSFxey0iDKPFWc0a8h8dXVGNZhIvFZbew6u1FZfApp
Qq0oko7g9wcyZ5JmxUrL8ecapUUzopriE2+qZjBHKJvBOYaWDucSlt9bP+SCRp34SyMG9VcTMHEs
hCp9B0N6grHNMRU18SHfgZhMIbmSjcOa7CxvMv2bZ+gkcBbyJe08Al923AWiL+mCP0aAQaBgeXUR
Yn4VRV6BXfhCSNv32lksD6xErnT5CbzRYfF9OfyMFFByKKbNndjKeMfeva6V1hr9O3uQrBisMKxQ
D1un4YH95VdIa6b1/vP7Q9WcQjzanq3gZMXWuXugLGL4h1WQtFNw0S3/6Ccbhi2Rzv8KLD/xCqOf
ZaaKGoWjexS/tWASpfK/dAgPT7seG/DiAyGRYFR286eA1rIL3pQXYserFFW1amNYSKq4WBqhYEn5
lcDMM+/Mh7kZfl8ysC9pMD/aGDthWz8LlX1jEFVsRSpSIqmsssXazkq7yitQ+O8vecoFsSH1aI71
IQCA4CQ8izlTGVjuPU2nelQzAcS+bpWoXp6gdx0w4d7cQfxxHDUOMHKPugcHg2JR/BX6mlD7zOOa
L5blfiAeQBUjmusiTeLtFfaj4iKtnJPRRt8r+tzZjPVlkecvWUyeKM3bllSbu/U9avlBByPaCaYJ
q1jh/aTMQAn9iuf1WDVRl+Woy7JivYsRio9/wqlzr6qqDx85JlVVwoJcEzQszc45G0kfD4TnTNyY
7awwuhmJjmqYN2dSX8AnUrZWLmj34Oi1SonnBIAGL39qoFDDA2iQop4A0CteGWcvXSu0vTgF9//P
thxxUHrMMvSzEhrz9QJyYppeh3NA4OS/3biGEImp+xGQnb3X2gQDJWA7Qt1TSgdGPNPoFdCpJS9x
tweU+vRUCPOYtDf6RTrKJNFD0Oz9xFww38Y5d8g3Yb5YLk7joo4egpCwkbenIO/4w9kcS7Ht2kri
MeFsuuQiWDiaCCW7opNBKbzsUrJD157iRaniV3g9bCUDtXcuQlHNo9bjQlT8CpMA6Se12szRqm3T
crHscbbSmPBCsV1qld1nxHmijX4NYouhX70ic0GyEySWPQYcBQG6+/QwgwGjU0OhdxATVF4WJUpN
2ZT/vedSVXwyXJZbGVcykvw0DOLaievHx9eq0QhM6SzekyGguwy0FAXZcEfLRQi6I8vk6MvH5Rnc
/RQM
`pragma protect end_protected
