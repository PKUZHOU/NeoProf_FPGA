// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
qPipx9hJ8SjmhanrWwftKLUl/ZLhs+kEYYLuA5aagW6dDqdbl/acOTeW6/Tbnwri
aYT7rm0FzAMSItGFEo31jQsGxyqDBQPo5aUV0dEXEp+0urAy3MYqEVw5u5MKEmcA
nyiAynCMGhNkE/jXN+jDVoV/Hm+EjjmiXelOrkLuJEg=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 8496 )
`pragma protect data_block
d73Rf8uzcCXGe9KGbuMJNy+yifcNI9AR5hfj7H2XLNu45oQNi69IFuca1C6zs+rS
EyZfp9SYmqVQjXVyACFYzJgWGpWd4/PVsjGKGjXxIYrTKDw7Fjtnog/FiEQezjWl
X74GMdWV8M9SNGdn14wn1QakCPIIVdTZH/c2MFqTk3htQa6QV0/AwTGC3LsBKBx/
+97OczYx4FtLYnFld4Upg+MthveucvuipuwcP+1s35KVqwuYNOjLdB3fB7OHVHGU
6YZLKJSXM0RY2YMIX9J38ZiXyNtXctFqltAUgoSTLO2fEpXEXN5clnLHOXxrvLuT
wCBI0zt62KpZ5cIYxQZ4jbfAEv2eTdTSGeu4LB4yGrr37YVPJ8t1CzClIN6foueo
vcmzJOzYp+XRm+XVht3s8XDKaR2EGeml3m/E6Ji8PaAX2WGwOTI+qrVfvpwv5X6+
XUsC1nucr5rgrd9vja9hIivsn3QQRQ0btlnqOCAOu+u0ilsOrV6lLmSbNfZYLcXJ
h0Jnz0i7hpVhpA7ZffJw0IQTMHZk08oqySSz7Z0ivxvz309EPdHyTRC3NQ6a8dg+
HRj2J/32MGNTAEPrYsUdXUwU66PRJmbU5yTifVpB9fftSBZyMXkD29bbXQUKjKAj
Jr23YErPiY0ruq4mNOn/I5GB4Zh2komVPNz6GjJs4Gjw0OIwL6RMCIuW67Bu/SXP
qg49rMoVvRnaiGefinNnT2FEyBudRKTZ9OVQuHh+R8qjsT2FuqPlY0lwkjqEcKwj
ApDWuupP1Yj+1FYdaFV4NoHElga5leV/qU7BsZalrL1qlRP2PBXTlCd1KZ7jKM7M
A+dGDc0mvjnMPArzl8Ij0Ihzg/gGLbpFTjLKis35Uw0QE/DhlbA0iwQ2rrzCNWyP
QyOTHtcrTU8SAa3NQtbz9fBzg5o5AF0Kq9XDALR7cBFJDDxKo5byMrd1iXv6NYyS
e+dePbN82yF1DQUlF7Gfmju11WtirkMLYewGjwWzI1xhtw7cgGo3rnmBiaS28EbH
VE6YAV1m2zfdWS7D6DeRhGVveCTda4CdLxJGi/UBzPtcy+W5KRtE+afkFLb6BZw8
emuj1uzIffQShsr17BBNYzszau+hXkKh48ouXlvo+wqUaJWe02CxSRB+jdT+qtNj
D+Bw6BS9UPbsNnWDBHNuOJoCpoJZY1jFA7W0j4Sm7qNoJPjmqXQMsJRJBCzB4MFx
fKyWuq1tr+EZhnPkDLhuLzaAUCM7s+MF6r44T+vW0GjgLLmtcFAd53LF7MxFatEZ
AMg2O6XbGbfBPPI7Rj0e4uvV2L0u8rQRcLz6AW1HaFDmqbmUvShwG2xDJOoHd5eU
KR/TdMK3cMpjj2fzy2otFvf4aCl2gW+Cv1wAyxkgp8f9o3EoHmApf/yZeTVMWQlm
OW0KhdbdqJ9IKNA29sOn0++5tA1rIITeF5PJMxDnjweLUWA2N5/H6WIZQ3Rr4jEG
/pRIQ2jkbdK0EWle1SSdqFAeFlvEfGs09subp7hnMYPS0l1AQ905KgRjG1q3LpGC
6CO+xOYwl+3RHQ0OJOvtZQxV4bq5O0nYJu77Ci4Zof6BudnJ6kSFliSPw/s+BEmm
hPgq6jZz3YlwyJmiKiCvdv1dVfvWN7KD4D5GZlvGcGguHzySqYNRgTMZPDNVkPo3
RmBroV2YZmjB4eiNFoyQuvvI24E1SntEEGLYIAyHojNU5DcvtjcN/Ypoz01WWolU
KGlaCesh3uzKKb/UlxAISZSi8/bUn8JQ4Jw1tSVEjstZjih4MJhiR5lXi2XzMPMn
88tSQ58KvCizBAiGDvhWg5bR49BEgnaGDMB34r5NzW0hiPMduBCGci3yPhGfcuJw
TCpSlipOE1ipJ3B8neJUyrMSsXoRPXMupsC1KZKAZYVsbYioh+NKaLzvVyBbqdgq
q2Tk5YloeW1uhcIaGOCnWULb4UkJlXc3n2ff91bTrlXyaHykDOQYsbNc8ZIvIqja
yPHY+4GWBHQF41TCpOw8CO6hzE4ytZehsuuHOzFTAD3KduTWqUIH/EbDmmZ7LHIQ
wij4YCtu5XL3sxTDlj0449etEel5mUmsISJTBxk5bIJwrw5awzAuuMEDXWgMavI/
ZL/fhV3js/Inym4EEiS7FgdCc/CqvHzeOnCTlKKpXPazbRLNNas+ehOZj5XMIXGB
+6OoH8VAfRK/y9z6MVXybFdgm5Fr5nxs91RaQcFpncqGxJGS+lyJxbNKnj2clajT
Xaa9Pl0efhRifXXYMfDHK+I8QsTdQBjjqNCcwCr5x1oJupZB6BWZu/CUwGciyENI
oKElLD13VdJOVZ2lOGdrqVG/4k6w7Ym1pxk02Tbe4DyiMOo/KgpVI4ku2T80RF3n
FINPbgYomscBDG2moZGrcZZyKdRBhZqNSISufo0gQXuKCRL7cnQVHgparGHV6w7M
qSPr5ksQn5xJ1JUxu0/GQjYlCZLBYVyZNekoYe36S/kvF2gHOLSbN0/g4GtpPN4k
H8KoSZfKpcUoMFHLcA0/40gaZUZ4ysnuLD/QD3svO15h2JMiRNiE67Q9rhmDzJGS
Ei/WyuLgh3WrkoWEsvTsQn9Z71QZ7i5Vh5gEdgH4e25MrKoFJV/VhBDKrlzkBFlS
akojd3hzozpxw0Nn3ufpYR19VgaV5T4Os1JYRmyLXuPHVROP3ojuWXVAGisBYioL
YjnMgfYbAJuJmmgSpDZKAbkfAoYbMs1yT19kpoXjdUxisZ8zbO1DFX2Q91LSIBch
sKOdG/9M/gZ4qTkxgWYuYPSOwqx0zVPKgjMGAWKAzs/2gWhvB1pkoCYxKGqGN4Sk
xwQfM86Au6c5lD4OylQ57TpzylZEc546ymyRUf+hOOr8U7STqlyN3rtmewK7nEA0
P4zLImWOOLewNNpxwMX38o0Fk+Tdum6IQxUWn9pdpiGteOSZH6o1Wc83teSWyWby
Orm9AtN/Bzq0XgSgkjUAUL4zyA0wvpd5b6nv37yGqOWMLkHb+sYTupEk8QrbxQ0C
d5/BG+rMOg7QHOitfSEWk1p8YYC1cLeCXbfaSY4fG+DAANOC6BDxIDHCIPwvyFGW
gMeQ5z8D/NxeV8DSaG6ZQJCHDZQfVA6147jljq7NqR+Q31UUI1/jv9n6LW3Vot0e
7yYMktLAl1xBsMiTJf4A33iw9DywlVRvHd3Ce+OCsKwOH+j85qrqLfUPhkDIpOOR
xo7mC1kElpsOo1A9O3xlGhDMyTkeawaa5PRIo1tH5Yst72Zr6ew6a6rfq/vmaUsb
OSTP28V2qeGfuy1x5FmCsRN+hcNuHyONt4NjUeYnKJZdQ8FrdgvelMIGnWy4WKJq
sHKzUwT9eG6gvHfVVrP2AYCXi7WF+FidTp4Q9npXw8id/nf/wqT6e9oBRbckWcqk
xoxEOu1cH7GvE50K0RsvL+cOrfZyFddkArl+bIe38CnV8Quv6kAOQgcGGQ/L00CS
woy9zKSX1Lu86e1dPc6vxkCr1OnScOjisk7wOUgbXgMWZiQccSYMkponaxF5UNoB
SYS5vCN7Fe8VhMsbPK2kg03Y/XoVqfFu6VQgqK3tSLUeRmMgMwmzX/cKHC1NQOjs
1Sw4ZebebPL1+vBIIZuHmhL4wclWUyF2fNmzDZotGNVzIHIGujOLPXxd4MY1aAme
DRTK95szNqF/7mwuFVgbYyw33Xnu+B4C4VQyXBLlpM4GZwcWkbvm8LQElcJvje7A
RAlSGL0vrnKJl3FmqzDEWmA7zpb58f1ZD4yqd+9W6qQCH6LR+H7taio5gnWslK5Z
stykDeWPMqqALTxRQsconfEp5Ky2jA5VFzeA+ewXWDIAG08jcQ0NlYy9PXhy7Nin
9SRMw2F523kHPtPke/AxIkR0dpm2aNPyDsPmuLXy39fyxuUYrLgMWgDLVUrdNsvD
NJ0GxnuDyll2lsZFn+4hmwUZBdPU0Is2P4/r/QhyB44ixwUzYAXpGI+EX2pE9J1/
uKRI47NbaE9yTAIYueIfSd1GL5VEynYRKmgJcPBJorO0pWYPTOaDU3dMeDoLWJmm
n+G3s/s+ypMCij92h0zg0UL+0+OKJcCH2QplpPKb3BY78sMJ88Sdklg1VxRQQm1L
mG6yN36Va5VpYxioWFOnLITRXZR0PtGsx57LEoI/7V6W4a4G+O0u65fgZKdWiz95
U5O0/yZXoYI4oTcsvNNbzRLL9bLckNba9OYFfrre0CmSRVGDTpn8YKk6W1/vo2ko
97tr9AXh7XmIbit5aH/iTfdulzXgtwsm3FkSV8O5FMdzuTt1yWVIqbL1Ty6Mq/s+
kcfvY4jMPvaUOK5d1K/1giRb8YW80LwS/MYjbpDpNq9pbSNOvJtZe2crC/vAKYK4
dNOfDdKWgyWdAq+xRELLz0/UCUAv/mqafOHNZRYeC0TPtD/Z32xxOpyvV+YMMEKy
t1fWEV5BEtUBUZ4TNB59wD2wYw4DqfcF7tHw+5dFVrvZSq/L0ozRR+wGNDltik4g
IR6Zs8d21QKwir2tLkp2lwcQxrFByR3xoHTmHXQ/VcM2IAj40L8wCOPf1DX+OwTY
GyAxTQ2kUfGKQsWeT5VPyuhqDQXyTF6uVEXzW6CYT18iQk9lwHePuOHCCuJkI0me
myWUZh/hqK+ZKDxZqnKQEWtbRuC9B7qaKSWv7Di1k4ZHZb3HJTjp2nHstDfPCV2O
TAzrVofypVqIB4AIljowf/ehAa0FO6Bpw3IFaw2zP9VlzLio4KeFz9g4jurJfscK
KslnRTvNn0kJG2sUc2JiZXEiwr+zknSFME3KvWPUeCUa1fm1wE186Y/ZOz88H/GC
yrnI9HDFoh3Hl+MKDoJtG09AzO8nnaITJvDJEDdHtzVWaBLTyCagmZPEnznU7gPa
DZh/RwfkT5yiyPOLIvtJv/g/PV7T1Pk2NJpddVaaFsrsYAZyxfPK3EREHvwNX/nv
RDYCTSG2pDnobo5l5ftfSA9sGEJ4pXQvmuHP6Q4sDF9+QYsm9RY5zErhv0ADz0iO
9kDdvsQSGZLqIzevC/d5Ua8ckxThOxqN3vrxqagryOESW6xQuOazPy07WrnxOUbN
n0Dgx//5A5UF0gLk+zdr2Epx+SF6Z8M7XWiHy+VGJHtimMvicQytcUGdcVabQzNJ
E6stKa9wOJ6IIJqIcLvZgBtGpD2IJi6FUHIfOBAVxqBnjUhswvoKdKQQyKkgOqGO
W4jHQOfhcKsGYsvTnSI+pLDwpuEPvtq2ko/fAEtaDrNQ+1ajRv6TX1IjHTDRqvED
5bfFfnM/Fd3D5femC9Oaocxxlv+DPL0nhBt0PCVNf+KF5guZlBAc32t1ZftW+BM8
uon6dNgkXNuwLAuoKMJ2eHYVLE9/tSE8gj//R/NUlT64sA2sLGvlKsADGZnEC5ja
mOMzt8A4OIIeRwXSRu9lNg3j21C8TOwpKifpuF1ZnmmQqVw7TXtG6vc1uVMLdWHl
fZl5ZxqNnK0/1hWhgJXdJYmVIs8O7q2cRUK0CzWkAg7hwhqXidv4atvMKYU48dqD
QObKPzFEU3q74PyyVTHheZSbnxZfXJE6zlS+qtUaJ3rtuG4p7HBERgbQEN4ZU3v8
7/x6iBpCOk08HW9JWvE2/56+mgITE8xHN4fVRpvmeT+49Tfa+hNbnIYB9r7PPQvR
lX9kJnVKFx/juASM+sS2vFoIKMMghr/Om98mPjgXv6i03qqDjcYl9wZrRRln9p4K
xFS9Mj9g8XPHoxVjGewYEMAv/RO+GrVBLvSFL2/NK8TglGcVr71y8BxE/0q4j7nq
FsQZrx/aYKTCObAiPy0Gj+hXsfMW/6kGlVIjy+vo3BhTMScgEctgLVsr4Q1TZzRo
rhYDZzfkyl6z2fhD9GbkmEcLZgOFsuAV4SR7nd/slE3TU2Nc83DF0kvd2eGcOuR3
bHdpQp9zWMVPViqKvRET8uEgAh55b9tvGQ972lQCoz6HfytW7s7J+W+xMPMoA/mM
ne9ZwsqN44YOnuIvtgGAh3Ti3jOkNGFR186CAVAnugASI4d0FJrW9eLOpF/+huVi
zPoGQtdvWdZ4/PNk+mmmZPwT8zZm3v2WBiNmeEjYwmZ8VMZ9zlcaMp7LWzjpoDS2
XUpZ21+a4i55nN4gqjh/a6hNTQxfYk1vDZwCgJJssVK9dIE0GlF1CGvKjLUAGNVL
py5/msYie9guE5ub0qArnzRvtP/VYa7PH1N1QE2iI3kUeJN4wuhAmPi19oRAj5GC
lsp/HuXTuGh8coiAADbw01edGONHydUfpZC8F0LMPHuRpDp7JMvxfzNdNKbi6uOP
qNLYdrqGEEszfwJJKOXt/rS+6lX5pGx/PY9PVvl9rqz/UUpmTtpTjJifLqV9Op7H
Jgr1DjzrIyZCIFLT2iLQIs8Kumaw97iuwC/z36Myo7K/EsQENxhNUBOzWwOLMG4L
DDuuE8W2a3uF7XtEOJc4/b/SNv2GASJMQReqWeTnDP++HJZrW3Pa9250AmWduAzO
CIyQv4YMakKyze3sO5LSNr8819B8Nt9E2XY7Cwdi++4vnBecD4EzOAHnyk+MQzyg
6kUkkwar5qtADbAL4orLjvDgJ2wvQ9/pT2k8qCUdLku3V7jraPntlqboUM4FgrLk
5sPtA3Gp7u6VccRjrs+77QDdQuR+6q4h2kupufiBYlXjpI6ybwCwxXdAQCodBdW/
kxtsiTV77bNm+k9UYkWWbMdrYZ+KZzKnOQqDGM1XEzs3PmBXxthkQph+qtBNue69
HjjJjcQHuEQZbcZNqrDj1eVxInWw7IaAMaPZ5gPHxW9V5Y4PNLt+N0ZS4Yx7f10R
qLRCtrhJbnUX8aT+qMgUl+VNAYLrAe/RSh4h+mhj3Q3EgO1W6RSwqVpRabTyyUOL
Up5NkRl8j7pm68uTMnj+Wy9mK6FPzHvmpNiAkKsRMocMEV48yLTu7beKya8fKDHI
vbmV36IJGTxhj6vuJpfuE2OcN0iafC40l4YV5HDpgbAjq92PeiqNpgKe/Vm/EBL6
BJCZMpV5pXBV5h91Yaiez6SU4d+paObTlZWKSHjWVQ+GUFFPVifuu9mFpCr+BtId
6g1OJpZmWY9syOnOFdPy/RRtC4/V3G6N9KUnN3f1+L/kKzCLVwkV2LRH+Ra7xznV
9EnqSXCv61w3XRirHCr5c2eFuO54MGb5qAbUvQiAxBXptsgUj2zwL25TbHQAuZeB
LEvXRqcwMInsIoxJzc7gjVWV3zP15I7572CAWVTfpHj2qYNOmc0rnP39aPzwjTwL
YS8oQksp9SxzDYdl/enAs/rxrSJc+yVg59BXfgjYOtoSyP0mBt2AslHMkODDnppC
sQrE959jnqL1Sh5mGuzoK3luuIyonFDlK2L1tEvJDwxBgGmQ7dSXlsMecBuX71gB
or5nRGSe47YUkCnwN/5PW49sketSmafk9GK5CBZDVtXDrtjSnArH7olUB5HyR5r+
CzYB7a+vTF2kq+Jfp9wv9LThQX6rw/tdCSlF4RUIX0Z++kYYBPHYAmbguQoVrI7b
FZqdaw1gqu9GXlKv9neliK9fxOCarWUCpUJJogEQNVl1V9Rm42ZgzFhNA+7R6Btl
Bzz5BhV9rC2MYGTpGWoHvMKdKj8B60jhOyG8EiQSwvMs13n6/XGuNAXga5lk30YV
mrU4kPP1itWIOuj9XSJRTdQknTNPLSFiwDDAkPbsL+lQ4TgDrJXB3z7qU57yK54j
6GJo/XInj+NC/79X5/Fns0USK17SEriGIPi8zXJ1ARLOKQEt3V0W6xMtecE1b8MF
sWeipoZDAYt6bQDA1HUKncttWWp5QX5w/Pp2r7oI0vfPhqz6nZTSndSIBX9bpZ4D
5uZkxrxpEuVJH9aDUbZdtYuqpIVxjlJ4k1VAz/LuhqiN5A+8ZrTzTxDciba+5PSZ
kvB4AY7NTMAnkjkwjCVqr+ru9U/qjBr+LYTRDbBd8tSFAPyZW0lWRN499/kC+vG0
F6PRwr/TjTSO4TkqWtBZHco2/JwtxF16UxUO66lz254+Qq4ot9ag+ALolHGKDT4W
dZq+4sg9x4DSppyB0jbZEgXcyBbMH1vQan/IFqVTSUVPqeNbMQi7C40rTta83EyM
BmjofvJwSuTHfIp0s1PTUh1qLe0NCYvRsI8+a5kDWa8j6FmydHjRqQgAK4yuQU9Y
Jvz+W6iJxADBg0sgo1zz0p62Gk7jHtVwHerOqFY1tbiiQBg7MvMJRugqPiu99JU3
6Mg9huYN2FJB/5FU/ll7DEHL7VtmNV+X4c6IlXV8PHhBpgXyn6TS682rzZbix6p8
N+QhG86I/YMX3a8qYWPSF5KPVb0MvLs5tmExMj5VDfyM3CiD/QXNsiFqJpP0OhE3
VJR4ffUg06p1KyQpPAuEttVYoLfQB5WXUVg5bq6dKfnMaVaHbHbs/TQce5OKI50p
2X/e95nc9khEdcNZyvKYobH1MhFf6SV+8aESBGtZseTIm36MTSzjIbg802T8SCI5
5N3Y4AEtKULM1qmBFp4QZcEYumr/zw4FbpnzDwMDCPS7TEK2IChtrxT+2cY4j1Li
0NXh+8Z8zAcGT4Zrg6VR2YDvhsvxFBeZNpO35CxsqV2IwWfrgVOw/ko3SSPwmnh9
M/sL8SucTJXxzdobpP2Tr0n2xMsou33iH/F7hYEjfpMm0V5PuXyarxQlnHu97FOC
KY8IYDX7Cx63TvFhU9OkEzLf3d2OYz/jDDMk7BgeZ0Qq7n4Q5ESNM8kdPJ3EdcwU
bqzrGlsEkXDalUUScPt93i6+Hrg/5YdouNI2tHriJcLlX/ROIqtIm5FcJf1wjv2T
9SeUAC7O/LUU6LMvxPsVl8fiyNxbLReYXeJJpzy/b6b3TyRmSUTHwP2mhm3UC24/
XTtfX3/az15JlgqYDJ8Ck7v8ACUXBSc7hAh8grWgPtCWUzw+oH2XQmyo2x1Jci6k
YzPgO2U9ZkCheKonThpcCVI7a+IxWOYTDd2zQspkmgt1Bs7PGgsTRTjeJBok9t0L
2eHuYLflFNcrJdwtoLajEJl7zfeZyJ4tYpylWEpS3/WjzHzUzR0UZq8Xhg/qEYwi
AcefqXOnw0pmyNFZcbfPCxLH4kHFrLnFB1WrVM4lO8pRwwenkaIZSagNKnXW18Jl
+FrdNyFXF4rIDfJzi9GN0LtaK6WBvE6rLZYpF0xNSwiPh54aDPRSP9UejbxAOuU1
y9jTPiDrQYbJauDkXFOsSW9tdhaiRiG3k/N3Thj9YmlyATxRqP3KypJVrsIY+gpk
WCjEWfWytxRZ6NJHPBtn7Md1iJXbBDW4not/FY3W/ORu9ygNv1l1LD5t9kohBr6B
5iUbABeSoqPDEypp+JECyVEheeVuUmWHVtReAClWeV9r9oy6MkNSdOmW2D2N2wyr
Ox2pKtqY6ZrDUDM+oJztokm664LeKM/zTTnFjkTk46FRvDUu2m/DaE6+jc2eXI3Q
NG4RRJyWiyPJOrBUmDwy6mAsoxy7SSEusdQ/9BbCXwJnLpQX0YWnVObFy1Fp7tm0
wMcip/lGwMhlOcxBRIo9JA1WfREzCWv2QGKw8D2LmF/XnPrnhySFv0dnPXBHujOT
H7qEj37Fv2r4ZOJHXYinhTvt0R9QocAmsqWOE91kyQcSqnjr843cOCJMXd5aAq4Y
5JW99bwTInyy1hyzsBa+qnZ38C45rASUVKup6dacxYqhZL7PXZuENQZyrc08K9ds
BEoh3nHhzaKU+XvAwgj/3r4b/qjaWoannpjIyYf7OW2IusGp5HSDL9XHnhQF4kRq
qlR0igXJX+lQH+0IiFTz5i2S+zXgw+SYSn4SiSsdn86U0RZf8aSWkgAK17M+zPnv
0ZFMAJNJTnAvRPXMtdTtV6BiEmbetI+AFBB9LsKKpJWcCrpQ2SbNHUfCB4NDkXOb
EqBrAfwHpIybWGgvb1Khhyd4STpn0nuYSV2roSbDWu1CWZ4uNgbcXS7G0D6Q+/Ud
Pf0UULjp+5opGCY1ISj9OIs6iBGvXHsKfXAUA4g8BlodXnVa4KG4jLValdqXpyj4
VaBQOlmQwlRhJ/m8YmYyEyRkve7gid6V26ZqvkIjIRWeUDoq1Rs6gEdlgoOwKU2C
XbpAlhToJaBL1VV9MhgdaMZFxWb+CqQszrJzdBuOPffyuLhYvkYmXzRaW3OrTjwH
w0FbJYyjAiptUvlMW/pRtUp2nekZY6o9FNkekVPp1pKXRQCSEjlVyBKAicUJjeDA
JEPJJao3TWdwpLrDIOitTjKrFpopcySPFR328TFLqgO3999ldd9/ymygXUNzT84e
NWoId3jQUAGv6beFoX6rkhvXTiE4uc85MlfOiybEsxKRuJqU2O8OT3yLRF972Qr1
18z6VqM5Ijo51xL2jg56FVj1NdlaoLL517Q3z8q0QUVZyoI43RYrzSsPvhNOekh+
/SCRmqMa6Udd5uFtKcYHXlVPKjR60wKWTcDMo13sKVQspx2+rioPOWap1ycYmFgv
ECNSJk7Q8SSpbntFzCDjmhFAf6cvLUUH+cDNolWw0b++4hm0k9+DSpLCXtZ2a0cn
DfYD/flgTY6m9M1Uw8zA/MtxU254EfK746VxG9v+F2nvGKzDMyAZ8VpFQnXZD+/4
lEdJ0GCEpahzB0Flvx8Fr96CHgRNqux4r17rp4xIxP6XOkmED5nnjZCA/JWXGES7
4OPBpDXj0Ld6eL1Jkwr2WKiGh0HvOMoScAoFhKN3HuNYlc7xme5EijNyxkA+krjq
bpp3POd1nKcbAovifjeLaFUrHNn8egEXCLmRgceSzKJCOc/WWnzVWeZQgTHyLJQB
i/R9P+hbHW3DIrF/ZHdBy2jNX2hErQNfGdF0CgTU+Ujn6yCOziF5ELf+16nIkhiK
IWnWgKT26YQCwaIG2pRS5Dnh0xVhvK1T2b+mSYFPrcmMu3M7L7+IYc5Aoj2fbh/y
zZ92t1Gxb7JHHlH1m3ISIXauwzOAxRYIqXgHTrCd8xveTnDFYiPiMR3oCocwnqCN
Bb0aEAMNC8g/Ip/Mqz1DVqrpnqh2mTwLrglH8yYK4fWsCdSaQ9FtvicOOkmEBdr/
9ZPDrWboFrKaehKerZtixWof+WhkVK4xhDJEaZAMB/atQjl+ODSkbeLL1yvs4Pb0
0is6WMNLd4XPgDPIhqae8yKP14wCDVswsZGWs+Yg7NB0P3XQyoRHN9jkYVPbIF7V
KE+o+RlQjsHy1cTvojHxbOD/BtCQTo2WT014pI4/DI4Ozd/AR4U7xmKz98FSZppr
LbNQjeUKxTFr8xEKo/DoldJw/ekfadZBrNoQiDbSGIHM8F17Qs0ymQ3nxOLkNFf4
aKgyUn+Cz6Z6yLmKcUhBIe01NrERzGHk0KwHREWI7W0CeOLDDlASKC1xWL8VXcxB

`pragma protect end_protected
