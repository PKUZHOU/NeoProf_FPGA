`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
CV+5TBLsDr+oPqTNs1wKCYPMvqvEc1OSkwACmexSL/Vn7ZcvRuovcB1trPpqQjgn
XVeBJ8XFaB3TWQWwHA9mCUGdzdvVo8m+gHqQB9xSWS5gQwuNIpE2edJ0y5fPbIw9
i1FkpdyG4NAGpGhAo5KUxKiGaNt500ubuMsP0G+H6Ks=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 5552), data_block
4Fi2i9n7g91HWU3Eu8nnaLudc18/1pd9Pq7Dfdm3v2BtxCbzqi8dalEIXTmRms4f
SKoRBo2cmn+JBMdH3QDBCIbJzX8nN5B1sg2l9StglrAQ7RGOr+YkdtH22YsT3JV7
KEbVbhAZe8mqZ9mmMqFnQNYf8bsdqx6BuiXr3PfYfq+3N5YB/8T3RBjGe9nVZDqV
n1esofw0vlsdxDROpujrV6H3MqV70lYyjK1YawqzUvAeCVF01wY3IGDyPtWHRSYr
C4FbBKRvsbeyqKY0DjZsF22yp/87+6Soua6bru4B23J0xfe9YdCU1JurSTdCIVr2
2Xi8gavJAeowv8wTD7axt8SXeu2B7E8hH1ct374gdMPUz4whg/ep6gSDyht0iIzL
ZqdyuggL+7fZMMXLx5U0UQAwstqRFjBYZrcXR+FPafI8UpXGFRGwbPqCj4Z/xJdf
vEdD37n3VXXDDAQJ7Ul4jCZ1wPUaR3ntfp0S5NUK8JGdKC1B3FaEKW2wwjIKXItq
zqedhH5hXwc5iGRKZGW9C6NOEjwwjWS/aJo2ZJ4bI7+755CpU+BRF01Dq/6LLqI9
jVWh+WjUu7N0Ft2CZnU58ytFwpR5IhdrcqvZadVOW/T3vKx1f/zJlDenVIa0evoo
4pBq9RcmO3VEoi4gPGfX1zvnSioFXSFkLrmEe4Dcd4IdKyNZi80PDZpAStu4UyMo
oV3MWsdpb1ouDZGPpC6tK4Plg5Zb67SWgY+LYJeT8JijDNHeuj170ccJC4WpUlqi
uqndklrrGiByzHloNknHitNtuOZFgJH7CvcwOP3fC5wTdaL5Gq9jU8PoczcHgQWD
JDQ0xmpimHot6R8ywLkZ9+nfugsSUVOKGH0H54RnrP+LmZVYAeJCuOXNLhYpZwij
xsHzQd4YgUv+OQ9aza4qqm89YMLf3Z6UgbDyruD0fryC3qLcQ5hrCpt2GM2Lrxpr
okK7+ufzpR9ke3mlMNFD8/H5ACVN4zDrKXJda6NjDJuj2PPsbcRZRp0QA3A9PiEf
ezeZwxmbTlbfhi5NVgitumR8ZxVauEKGkNpboRZU1q9KD7M3ocHS8NE4wV3wmG9T
KXWz7nl2quUyt9/vqmdrx7SgPBGeqqZz3ysNtFGw37PsEvVfuvl/gzx3oU8rkh6/
MyW60nsi1QHFzwrR0VYw/YKZJMz9X3TdT6VIFHNQYyelauuSmCF9WHZm5CLWvE9R
UBLZixO/fwydQrZ3nIFQmdr4wNzsSB8o8HOXBTkAa9LYPpnnCiYGmnHap9rK2fRf
zMAv4+SOBFd1+ydQ0J55S+GZggTPFzLrCbTcAMoWqyjqjMJ5qV5q5mMLQnU0AFNz
MgVk6JVpLGW5J+b6Y/MSgs00PRPup2lsQHM/d+AZdBppMjyuSb9HAp8IwXTyQG1M
uVckRy/AXjFnVYocy9Ne9inbDQcDAuv3XYCi6oOR7NU3tG0tMjUoZYfUBsqOAITS
ScbPbz+HKJciXE86p/KZ0786Rmvgd5eXMcHlRZw+mWqMO+wUju3bXjHUEfUgya/8
+m9zCwwRSRmA8BzzE8c/tcMeOeC4oAAaTO7YLgWya5sj3sLyEbY1fbQfffClx+Wm
VAV4TrB3y5gVUXcFA4uZwPPiT4TOeuQaJiTvSwq9fhL8ivAsJlHtl5HAsh4Ib1P4
14wmvi9dXyDDk/rnFCqz+s35P3hV4/C7TUca4pqtP5mLjGRmIxM+ob3UnxesBK7m
wvZHwoqZQhsEl9rm2ZhngoIMuMzO/Rr+cpFsMUPeYYYVGZIOjDC8a2xIWSGLwsNx
rx3Ajce3HqFxgAtP8KYXJx4EQoPv1JyqQ0qIV/kvl6xTFJYPOo99glBqYKY1yE8L
BFib4u6eIPvBUlKSsCjh2ocwY9+a+kxReKuKjiutcPBqLTIJacdQf3+yjI+LFFKr
iPUePvgmhCVcOUXh1Hv+RTXy5Tb8TVWulPmHE01PxMEsZXRW79f1KU1D2PxRU3Ly
gvlszDjKspJMYMTlF+5JtVAQqRGXlmH5UKreTSGU/PDPu79dqdsVPMFNoM0B0+T9
3iecOejzUglyqf/34u+IvVwbiYu8dOCHFaBO3cxM5rtY+VWa2f0fkqdjvpxjbjxk
3FWbbHDpi9U7qlW60p/4ixoyhTTurbLp0sCRjD3iaTYEdtBYNvJFawZD+x6tzpY/
saDVK0mbfsOafVnyV9CInUTCVl+VKM/TRsRd7j/44KDOuCikYkF+w4p5/yVwewc3
Gzm/6129uDWruWaN5/Bki6BSwJO2r7VuiXnHgLsyPdHsiZ5DRUIk0J/HGNplX06D
ZT+UqX6DHx1TIY2pIpqmU5RDMMpR0UDReB/JavwaqBQsTe7W2ftsE8vb8zCtFN2w
ntnTyQDHRIu9UPx2zbAAFj/1R9zVKGvMrnY1BPdfh8L/hkzx4kjknoHQpvwQg4oU
0GDUoN2fvkdwCP2NkwnnlwXqP2tKVoOl9hi+JiSZJWRqLWmOydqs/b5xmo04U1vc
G2bO2bEZHy5FFJb/tffwDiaLJPp1ay14SyFIYCyXj3diGfM9o1Te4NyJZASlimYr
yKjv7dQmqMyboHsjUZrSq1zK1LUlR4Ckvazmqxalh+p9EThuuvmVURaKfzEl1fG1
O4gqcN95tYnaKMT4DPkoyV1sSxvyAY751iSMo+OAp9TliuHS+CrybUjHyK/mSFfy
ENwP+HGOgiHUQYEX4etvZtqrTao9c53IVr2XsAYtbri/1P1wCnyZhnng4ANxfTHc
plWIFtDOhRI6l4xNKKokomCusV//ngojnb64l3gzkl/SRPqGNYoKceCWevU0EXfu
i1+PlnPVjesHouHuflTpCOAIXjQZ3/pDd2IQbGWM5zVeVsugqTgmO3/VVwIQdlO+
+kSm5sDhuPQFed7w45UoOtAySFuNXm7Z4jM/njzkt2V0G+lbjHfEmQquyIuULdXA
fZk4Q2lrqxSwJoCxZmeey1tRe+YjYhJesiY6cMLHe1jf9sYW5EyIfdApR6b9RPGJ
4kAUncCxtrZpsPsjpuQUNdAD468tKxdR65v42YvBD1HUt+FRQgDNIQlvBmxZQ9Sh
jK2trCmvXiCJip6ZY0eiOycjp9E0cTrBbwOBuCg/dSMWdrA35m3CMOpb2ZqxWPCk
agQPheKsnbVfIMgyY+xYCvlo5fnN2O2rYQiSfgY5lP8o+jgBivmjREuhf80TTRAy
v2qG1ki2vhHfZjhE81ILD91mmjM/k8wBb0B6Vo5MH1g1ncpTDbB7WbIbzNufH9Qu
sb4Y5BH60Lzndt5IlkkPdAmYkO9D7bfLDVbKnxoui8PuV6jjdlr/Il74dwH+Lkrd
kXDUw1jDRn/2A+N9NMycJK29ffxuWFqZB23b/SdhR3OGtuU7nhxuu6gDIx/MHbli
/s+cb5g66Bk27d9jMdalTeoSbW7hT34NjvBxQVK9FM42H9O6s1vQdrxXeuabGQsg
MEr481DaydlCA6IOXT2oagr5/aiHZTBCkLovOuJ8Z25oIBYiNSC7yElMf79AFnqW
2g0QfCKrUHXn6XoZPAf/wk0jg+Otp3GzvOojgroROTJlrd8Dr/VBo0p1lxnQiobi
vvSzA4OIX/SJk2OGz6usVb5ovCkQFo4GlYRHmympMBnUrNIZktwOszUCidhkHiIm
RrZ6dJjMt9rKMvaO6TsaZ0WrNv/u56Qiq8LbHa7dfDnvOWAw3DgDe7d0TSqIztEI
+MOk1oKN5vQpkaP+GG1USMeOK5IejEETad1lMbfmnuJMDoD4QYxjdGzm7W35vs56
zm1oMcUmnJyMkfj50AeThLmJndw0oROoRSL8+n0XoClY+ObEG9tAtDUMqbXFMw4F
NwHEBevq8q3kPNn0leBlqe5OGxDqw3Hlxq3rVfGQ/KFyq8qotgqgMnyQC+OAN5Ds
Aqb4NKrgF2yXFFO6mlI1YTBaxGyP9QKyRaVteYHb1fBiuBrpXRmkK+HeA2x3R1Yy
sM4mMcpsChS/zPtc3JUnFP/DVzPGTtFIRFlKY8WwycFdkBZl9d8hxQlCBvM95/6n
rpdpj01A62P+CZ/f8z/mCKwsK32jbd7JyX4qfO7sakwg9/xW0VQ6aVCe71EFoNti
hvjnXMvD6D/snVdDvYKG+LSleve3Cs10Ry5IpvUfwLaq7m5tH4+VJRtoQjrQfMLg
0zS0Ffhr/EcGajvw+iHnDLF7WouHLt4RciwrbE5pxKL4gkgqytpGYU9G9CAL8Vh7
9b4hgC6XOzRszvHyEgGgbgCa30dBWnP349GQuJtaoc5lfTuWv8uAvNl0WQBk6AEE
+Tk+ydcSpCSnVLh+7nPbXrNX0OvKL1jZnuQrBycY1lk6o1C3r0QhN6L6M9gQJfc4
mpbLMMZjXChRCMta4aYR9AzTLAs2bOa24m6sXcxQAOtrSmyg/xE5QlpvjYYxVpYU
6DijQaR1Ac2p9FmxtNbzpbZc5A64LO6c/5G54xkNw48tllt22sHUl20A8xYmP560
pPQx3LFYnaIiMNEdfx4uY203kfhMPNjFvHwkiZde7FEkDFDDFCTKNxBE018O5jA4
tYQoWWleYtpUeEMJsX0UDHKEoF1NnSyNchlHuUzmtEx80AXRLTAYOEqFqe0ZC+Xh
UFX+rM0nho6hqhq7V276mBa4HsweaQ0YpN9r5H/gS8zkcoVnfi9A7RApQd4YQODO
JwLh826kb2rYcF2rElZiJhxlALIlJBkDD0+e9BItDGqKrgW3f5VTi5fTEvTlJjK0
Oh8AulsYJ+rD7xw9IelwTdH2TokkjUE4MkAAF2IWqlkS4TWI5MpYz33FTkDryB0N
WVyKSdMsEaRN3BNBKibvSOpNuA30gdyr0ClIlTBB1/hjXI2cjn/bfJmozCu+t8dr
x1GHDKlKQdEMpOHCX8EXdwBhxBZtF4D8hHIc98Kb/wKu6EKEzgK/UC5w6ODQ5Ixn
XmNPk+03lb6WBXSrdPVPYybS/p75JoWNePhDpdfGAKGD+WrSlOS1F61TARmQsu/7
mJFAOaCuWSthQZb3D7FnpfwaprP73j72udQzZeh7uiFAHBFigJs7c9Y7KwFxQ9rV
PRdrI7XAFFbd8Xg+XPs+ewm77m4H2IsfS4bq3lSqGUgjv35h2kH+YSNw7YJMd6Qx
gw5a0clRNcfiNGJ9gRZGwCpcQhDWHu0pxSVR0JJEma37WofkC0/L7Vce+m+TtcaR
jMGiB2m/yVLUqRMtuKc9OHWfmUYgt05XABnJa0hQhqPK6SgsjGNBRJUq80nDjaKC
OZkzmCiitsNZkLoFu2NXLWCCRuUTM9l0pkAIkUBo/J8fqc+HmwMAs2hkl91FXvKd
3RAK7nke0rOGvfKEQqNFmiaR8TXBgxuv1Zd4JDEiNrCahOHKFOXAkna15KLqgbNz
ubLlDpZBNuIofd3GcZnwj75PgkhLvLMzYgJOQVagOH7ODCwP21F2zEchRXcHxvCq
3mzBCXB0vMLSv8sgY4A87Gi5qigX70HMtDcTOSa+oG16gPdOXl2l9ymHG3UuE1Ho
DyAStHh2gnW3GlCzLcLUNpDLlN5xmyqngpBzg15r3brNStbMoqTfdv6NuWI+EB3Q
jqu87Mm/1z5MtvH1dTTz9AAaNuCvGCBNGFQB9luMs86stgRUYwFBP3mlrOUKT9D2
pvukuJqHRL9UM/Bvwc48yWwSyfboCssoFbtozlO+gbgc2HW6ifnQn7eUdyRWP6sw
R6BSGUMHOsFIXw1xp9USVnumt/ETIEIGnsyT4Geb8hU6c3iJxNvK6vLW7ttYaMeK
AlxLgaW0eqZB/sSBmuId2h2SHtKQ15KBvEswMhtkIw7Mrqq8g+lKCdAzX91daAJG
qq1ipJ8d/Oky29Lk21bg4jxgyk48hnS9bPS75CvXKt2GDE3n02wncGNv1YYh6QJ+
99/TcaOLyitUQ9dNOK4MBmyEOGzNeLNPDLNcMRCMVtEOmShXHPHsK4Btw+jF2dld
qF5fTYiz7WCHI/ijwYaw+mRPpIWO0tFz9j5L/ce3nrQXBtq/LMPmKcByIqY4Ek+r
EZD6YHW1fKZ5+NaayI2RPvgKgAb/23o8NbUwzJVmMrYrGBNfIewgLzTngy0HBn2G
xn/TRQ5Q8cJ2gRoiltWxD2X27Qe98FaU5qi3t/pEBte3MT3A73xa4hFMVJfu/JNB
CGghF6PTVti77thnf8RGTmTl0AHzgoDSpQnVYPY0L8VRL93boNApcg3opKrSjd3Q
hcOkCBWHfIHkQtw7t/eg36zveTuWUuj1ymtdhqmhMtQD1QRN1iCwN2EoL66BiasR
jjQ88Jegq6+NM2+tFmNyG02qhs0PaU/1jTXcKzMW0MkgupwoFVgcAxEUapnase7D
Dha5x8ZgUTLMX8x0P0yNC8147VJsFW1GlEWG6JsbMFhA/s1EQa0pt0ls3Ye2XUxt
og4AJInnJOsoJ65gmAKw1NuFKzsY7qMJS5YNkoa7XRh8j0O5UlwZFYWoigwQjYrJ
kY0KphwSZtBLD75xac0gDxTR4Ggr0Wji02jhYn37ltB40O8GTdy2OojGhGI+44Z5
oVIwL1pOuPELNOfJh/etRQM+R90TjVk1M1vP3+vIgzQlSRU51zijctxpXhB30phx
BrNKLFJwOZeHeoctOc/VXsMM4JCmozB6gYA4WZJeoqWsyMgbq4OY+na5n4lU9Jp1
TkLzE/uD5nG9iS4808xe1QQF6/qspUSqJc8Gsb+Of9qQsefg0IXvR2i2EpxTPEbj
8XJnGHomNuP31XgYcMfcL5Q0eSDfKSwBqvv1oeZTrIBsb1jDZD2ruJeP5c0iwaaf
EWMaLMoJ3EoCANjlwyR2rTzohMkAKwXP6eGgXwsOzf1Az2lGbeJd5c3/mFBNyyGx
XFgj4awsV0+5v1y7rEdVg+z4oyP6aW3L1VszJLyzO7lPnoShPNAtjhQVy0+Y9cML
OZajnLV88cfODb31PBOZ6wz1Tu3OBQZkztseaMQBI8JVKKE6MO5Ae6FAGCf7o635
3NQr+3VTkoTNGr7e8WDrrun0qMvdR2mjDgYWxlcZip9QgG20wztNofVGN0vJ3z9L
DOHwmfsEaloL6agFHEVeZVaXfjQpSd/WfC4XbYBjwXwYJGqnS56+eILl+4iezDaE
8qw/HusKMA5bfNBqDt3nQX7olTOYWVDFGeKper4OL5V561NyQ8Lh6EmruyEvTAah
acKI+I+Lw63QGzY/a/0mEJV3sa1XqJa9T6sN2wNmNyXTypnK+A34VP4BglVtmFO4
VpiTmr0EMiRHQHE/VomGzHMenUGSPJHvo6grRD6goJCRuEhe3HefJirit44dj8vX
CpMbx8KUPPwwyedrc2nOsIKfMEy3+YMGFt+LZ7El/8S3k45LlUYqqjmu5N/BpNAP
Vc1P6lbBoKjCDpwDvZ5Qwopj0I0rhF0uFDUUquAIKH0=
`pragma protect end_protected
