// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
NSwymJPXiIq79OacBhthWh0O91WAUZ4MsKvEru8VbeGQnO3tkdGrzw4Atgky
nPXzOD0Y0evIOTzh+ojxfW1pByNG773bkIdbjCOX/o5iZrc3NwgCy7iuLT7Q
LR9BvINlvykgRU/i0lKq5/GuT2OzNvtoChfMyrQUkSfwhP4nLail5kt8GWcg
yYbISDaLIIEbogUb+2JjfTZok4OfKLmiWmBwoV5icRcywyvDXpkSMmXoSaqo
ZT2x+WqhounY+2YEzkGWvLcqezfjMwQFnK2VHFKP9M1+C0HK+xqOt6gAl5zO
YmiqQAd9HWcIM3ecbBwiQd3xmML4OkgOOhA3x2nx9Q==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
SCmjp6KdWFQyHwwfcUDsUNScSHu1TRe1Q6THtEqHuRwqnz5R09066n5AwlFz
QG+j7kKxrWN2oBPYHUq5NW9K1OsnWBQj9pZKSRUGk1bjREyAhj2tE24VGUVP
MkRB3rCF+S0j4DDKz9sGNLYfboxRy5Yx/9FfwSL+eFpfM7iqHxwkpfGp5GKv
L0+junJzPbNph8MotS7f2YMkuIS5KGUh4/XoTBld2BsXg3QuWQvLQgOPnGqL
cvdFMzidQuA7GAzbg79Fv8k2eq6a4c+i/Aa7u0lgNBYLShsYBfDmEBqW8N5k
wv1Uk2eeo5kemHSBYVQOXSU27/+CHeO9GUsRY5+0Dw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
edGPZmXjN79UptIsqUlTjlE+YpQXwfrEtTYiUfWjozG+nzC6ADC7nKD+//Ft
bZ6cTSGNQh9cHbWVrTIFiDfq5ombwVRRzzIBVtlumr1fFb2jjOQnefmLVae/
dV6csb3ip/hgsMhxMeTEOUKy1eT33AZaxnJ4HUj9prb71FhmRn3zSqC2Xn7L
O8TjBcUu5suKyr3ZCJ0kH2DVUT35uvao/uIpdZscSJBRtQ9lhS2L6SxFnFxw
I/pmWaNIFQtzRW11KIaX9ke5mcenoEzkDVBhvuo3FeKUVJe3pPeH6impwZOk
nPye6OoJu4gXKvhxwwEACMf96hueqUrWlqWuQJUl8A==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Q2XK3cddf0+/J78WujhEUK2haGIszimuMYVgtNBx8gKOvTTaDdMeuANVTz2g
aPBGkmEaE6qP8MTli26h28FvdifjutWoz2c3sbwpuYsjrYkYrML22iGprw1h
yyuMuiE/1Opv/lKXDOtB/j3TcwXQ+0i7kHbUXaoBJXqCYFmQtlQ=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
WGb7wdJZvQrphAYsJCZQu+/yfbPbjH43IyRJ2IMgcPbBIjS1rt+nzNIimi87
/5Rbrk7yMPBsJGDx8wTMe+KVHlqmJ+aYjyYoSM0+NN1embY7t41sdtiH/LOO
Hji5gJyVCAJ9Y8bxKVjKmNxa8Ac3ITTFCaXYEslQsk9twC+eHClXy9miOda4
KVyAWsNtZd2nJwxTVWAJ6Ini48zIpDDtUFi8F9v1pEHKTS+e6SCxm0Bu9ZP6
iaF7vRQ2CKUDHfWu2Sposnzl96idKf3BAoPDutaaYcv6Mb/TNHgpg2AczIU1
ILWgK53450L+L7nNCxzeNeCF1mDF1KnTAYEjXx5yN1yCkmZOnP7eJaIq4Ag9
m1ZI+uBuENklenh80y0PYVRgaS546Xs98vNcWKcPTR6TzJI74xjdJO4hZR3Q
qSBCEV6POm2iKeMFcGclQo23AWbQl+HONXezGUpjLdiAc4jWitnc0HoU4pV3
aLZTwiY1LWEJZ2/7emX99QXSnwYCbaqm


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
PB2WhJ2bmlB3Jv+eGN0elGb/ilyHks6sgg6UzNKbfDvIzpC8+2NOOFbxu3VB
t7UHKz2ZQf6HaAVNoCgInePo7wZVmWK6raSfmgBmixtpuyUJPaStc+7W7PqU
r6nE8hcsxWsJyFrk1KbSIODt2tI9um2HSMMKDk86+bk738byq6Y=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Ogtg9i86O89DvE9VBpfLgNMtJhec/HmtzcBXz/UFI3N3IRUtM4fpPMaAN3M0
NE84AcwGwOsMju0aBfGa3Cbe6IWj1d5EdP/OtME9JzwH3A77gl6wjdp8vc70
MIyzbIvXbS2hQDaOBdke05CE4yAyMOii7j0bGy6j+aaLoY+UVMI=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 31216)
`pragma protect data_block
D/Gwke5sW2FJkmSdicP0/SodTi03prhWZnH0sTyh5kyTh7rV7TmfBfoJKPP3
K6HhYYR6iuHTLsgrrTniigmhoiR1m0gDVtISlQjtKNxtP0JihcTubqoqShSN
zjUztsWnLQluHeEgUdppVLCHDC/MYLVu4NxP0HN7cDLLrz2WgQPT+JRWa5BW
AzUOs0Ypzvrr8zxGIuYSkNwSPpnRjB+zvZmtxl1oJFKhgOpijqyu0JCza3Mc
iM9xB/Nxd7Wydz8Gea4ZZPod0q8vOax94oE9T2g2PrtJa7stT5xzQnInPSnn
5CAsHhvzV/7wSRpeEjuvN2NSYq2dJHfyT8RvVs0jb0sAP1tv5nL34QhhoU3I
xicWYu6M79L3+x/YdTEQcicK0SEcIoHCjx6FY5QV8d+rgRCCi1qMhiBM/Bd2
ZvurhBZDlF9qmrw2+eApL01bvlKb6ZOHDMNq6ipWN45i6bNGU/GfxK6h8k0n
4q60x4It9ER3tzZq0EuFTIPpsU8gPyasp3UgY1+gRXD0IhRQ5klrvdZPujZE
RArQJlhz7EMq1G5YCCDmC59ISmV8vIH46iSmgN3pLVbn2YDIfwxOC8+fzHPT
bcF3FlID2ixCbhNAl/cnmnC3o8JKGiXZh5dtSyime5P6O5V2viPEN84eRxYm
HnfgFiQsyoEG0ZzGqsJPNkZitU3JDkW/mkVa943RhZ3ue41OecPpRzbJl8IH
4Z30Evz3Yxmdq6nH/N4Mw6GnZxj/8QisITovzdleDAO2gd8D6KUxtG6GGxyx
Dz4thjxz7NjLxtBJckdafQThHp8CP4OwcQbfA0ZREYbeU62zMCd5hBossQ+C
nJMp1fIDP4HiLMW7GsVU/MYejsLwtegHugJji0yHzsPDPCx3qt3KR+YOwJZN
i8XMVOMzzU2D8OkPysuPEc/SF3lLUqZ5BmqhXbgHIN9V4ELzxDXoMn7P8rtl
jkzanq6RJDpT0mzvtmPbVFu0QDGnjreKc7u8WmSlBeXSCET4Q0jimt4bu09u
Ue2Ium/O9MjHabA1332pFBRyOKavkc4YcNES9vE1wxw4MDjgovIZgerykVbY
WNZy4J+P124LxgFTrV5jd8SHjvczjCDPLA/wpJLJhCcDFu7Vm2+lz59+9VJR
s8xKfNX5fIzYGaxRTyWQ6UJold+H+BMszCmPTxJnFvq7c4M8frqRqTLbjWYt
HnYOAhy15GBLZKuQ151fjzBssKWHGhWDHq6H41NQyLQP+DX52l0nTSHmA6Oa
uqMlsVulL6eaur8HgVKwYvmcdJe1pBJJmtxyuFPATyGPtiBKfH+l5mAruz9u
MthNwIAy3LxaNw6VU/QRj4e+aS+vs0apmUdKySfqIA7T9am4sGsYhBAPfCCi
/ABCIybRd4wgyy087KSKwmMDXPCBUVHpHr6v4Rv7Un2osQv69ZdMIk0IVrDF
/BR2+wwlbGwHwoaDAP8KgGSMlnBjjChLJJ3QdsIBdLiQjG+lRAaTc9Fmf15Q
otfCQLf870FkiX8kgLGy4R+l1pP2G4BUeiXbyLvyVJ17aJToABlW79eg98bC
jMQ7U15/FPirQxsWBuCQiR7GbvvX+ZRCcyPqPM5j1774mXMm1emApKQWKYXu
L16Sx/4bVGT7wk/K2DN72ks5lXNWyafuchyTzQ1qaniHxC7F7/jxTK/A8HOX
dEGSl3IwUClRRMmpeA9C2A5MuvsK3jbG2zMlEbOWAlgle4eA1q+jD7L5JoP+
u56xgiwIW3uK0OFud5Qib6jBnGG16P1L50LbC8yYXM9Vvv7JqvJhCAjIZLIU
0AyoF5OkuVmgIJLtfQ41VFqCWBzdCVac9/sde/50zAufTHfNP56b5R1+XM0W
BHzqkbnDRUD3m0Balx+PTdtrYvjvNjt9DSXQ5KMqQAUpXGT9Oi4Z7qPsUXk4
o/Itk4lwA0DwYg3vVywoA3+4PdDCSQtgCx/ucGb5byKXXUh2wzr7vv228+IK
lrXXGrTx9fsRCxInkIN4ZyiJ6nNLFTAzoayuIRYsu/ZJWsFXRr7C9VWLgvhh
5pplEMm2UeANf17/InwqkLoJ5TSuPkrIGZXqQqqWuQUboIMMs1BJk5Tro4/4
6Bj9hMhvy2pPUm7chwjYMWak5GXyttcVUbMPqh3U9gpgxLoaCRQ1egKwXHwH
Mth8IANzhd8at37TVyuUblRpThDSNRZZ0Fwu6YJzqwEM13b6v2su3771Dz22
1vXkwd1MFrtPgAgPg3IHdtb3d63/8IYBBl7RlRm8APKqolX6v6OvmvDS5Fgo
+6Wd7eNdKoXjirM5vFT8VtAsucKbXo2D1ADoPfxcJ1gf6aMjS/xxbyZUfghQ
/VztrqpaQP80KIzfPXhZuEXoP2Fp4Lb8PmJveTSLUYqQHy4mCqv07mnVEpEy
uMFpPrQnByyNoZzAiDKB0VV4yNvDBUgAJmH4AVBtLrCi+UivV3G75jmWAA+f
2wWJC/w6o4dTLVub4UkLmg6MCgcNNtl6GoaBvSc/aTY+b0B5ZkHnBjbmBipS
frJV0pLQh4s7VOAEzxeIxbxSHdskWPHi3Z9C1jsFwH8VS0Dp0NTPDG7htiUh
KxmnbErXez3sDGpb1UwhiFpRVMHBqGdZ/FQw681IJOcRALDzK/iAfSB32nXf
ZrynfxLc2KZu/dzp3fb8IphUf2RNLGCaMFrrUoQsA5ZCvrbR3bp3t8eMqY8b
Rt09cvoz1b4VsShsmAJ1h65zoWfCYCAmOryhyqeC4VZJOqezynji7gmfp/og
3eQENcUPAnSZ6OC1Lbxi3gpIkS9CuOB3hQ9Lqj0YdgrSyCdprqFxiJ++fLyR
AWkCoQpGVrPd4IjL9CMsOw7CHy2+WPJE7ua5r3VhzHTrjduGvjImsAYv+R0a
OmQ0EPz/g6LPzsPGvKB4MY9hnaEXfHk8diWJscqJsWyItK+9M1Wl+lGmZj2g
9dCeHIeUBPmGebPGstT8vblv4O/f0MNKBQLrPzZt2V4cRdAU0DNzxzUIXDWa
fG69aAH+jm84Ec9rcz79bV8+j7CsHMgNNMnr1AX3Fg0cuHteeceWrXj/5O1K
QYoTkCs5QqUxUqdpbMMMV186GIChi+yffoAlWG16BbeeLsk6T5soPsZ4sq12
Jqbj6Dh/Bsvbh1scqmZjMqxVWL45kEn7nzr7DH8rxcqiC9RDbb0T17uGCYjI
3PbWssBrO5MwVN5+pCt1Y7ZWXsX4IwWZ6tgTBjAMmEhYh1+3GeeaP02xablq
p8Oo1CR2EE9Yf6cizwgjVzek7r7kOPDoe4Ab1kdaz1K5rc2eczcIcebHGzcj
fR/ff1OqWyYoJHykYovzyZoHa3SGk8IgdhebNyh5iZ1cg1/M2BevAxaoMGPB
HFJuQN/YMmmKKJvCFBbNqALWboT7mvCfWqQqGfyB5v8InkmKBV5osbWIAkSx
VywMzyZdjbvgAEIdEsz9udyIxXsl046GkrgAX7ymdeGe51yfYP2Ono3CoFj/
Qbj2xWe54oi2dprLMV3agRJge56KDeZJPOR5ODnX6DeakYxBmTVZcnsImn/g
sy1hm+8ggWbnEiUarw0Lbb+ZyslU+8u1uSmDSf7Vx5UCL9ilMcNCUlA0/pYg
BoDFhDiYuXNjqPpAdtg3j+lr9NrDXHyZZcwnWbcOMjqlJ7f7MCpr7C7/XbRK
6IymxuXNWYt2YSC4Zmy0elL63WpYoZ4PuZu40DKAvt/FkWyh2xrzBKi5e5VF
qApU1jVowAtszldbBCxdJhX05SONJ7j9xGB6b1TGU69Xwki1KxO73To4ffZ6
XmqB1bydSzbJapv/+rvkMMSQhDVJjxfipRsYaK+EhN7HkfU87L+msHWCypli
goBN9u0kEVKlY0SbcfSIMZotrFqvNnyOYleaVK6B6r14+Q+8epDC5HezynPS
oqRmhw0LeB8eOPVM11j2SvNrEak0CtRM0+6RVqMVhkDKGFvirIu24UDX0tpI
mywmbyqlRuW7vqOj8ZmixmuD6F9MM5h5QM94K1pstVtgSN9vVdZAA9Lu82ph
hERqG04l34HpNa6dYseOnwEfNzoiR6z5p1mZOYWs399tV0LP5whziUVPisw0
MCRqWs3XMMswdwoBQXMv83aLhpEPV0DStJCbm4DQhZ1Etwq4B9pIyZmQu6yO
j2qcYYLZVIqsFC3X0mEoVZtqcAhDncgVVLXlxZCQUYnOe4mFTtbhTDWn8SvB
1E7pRHr97LtfDveSrs6tu7nREEk3IwwTkPjH2oggkd2u8fgb5CL5rUC3/s1m
ad9ZVtp7pCn2QyWL2DnMP7SKWE/o1zwVukwirEDXn5sQDxAnUjALxxwhv6tF
txxhu1NWahQOFoBVk4ebrW/avoAOnW8gEUdHxeS6u+HFM/9t1fhBqMoXBpcl
07V6GUcC8l2S6lcvsKs/K3oovpN3d4+17qe0kgU+R4Y7qpEGLG06/kAjBM2y
0e55M9xhkE79FJeRPmgK7fURkiSOIxXDqTMYaKlTNZx7HbX6e3FDqeQn0wjD
z1pzoEb5SqJP4AY85t7/2q1MwXtnhETI4k1TKewCuSvb6T/lsG3SXzDsJ3yP
LdX54OIOdr55gg4/ak9FVz5cGUmMt3VPd5+czsdbGzwjZGOJBPDlILM79xTA
pN2++jc07sJTzrvm1n0hIcHaWEvTMeDradXVlKOX4z00nHlDyosF10El1Kny
QNrrXYZT2UICi4SH/rX2JJqXtx6a06pUjLkQi1xCj95gr1V7WwcUmr4qyBKF
Lost4iUVXqhaWOJR7bvS7U5bJqmQGtT5UgffrxHWLFoTERGwvvpXuoH3T7je
6bSHlpc5pJvDz20VYEK41zUA3GaPec8z24aLEfKp+FYurwfjlSj2sxy0u4ip
XgXy10btRXsW+l/jj40VX0O2rB5KVqTGtkGp+suA/58/su1AukZEpnIdyov6
T6gZi0prjp/5goBn8Tm1iS0feJOFh2YLrWyfpNGYqrI46ank0f3fS/T4OvRF
sbFby94x90vqfhVX7MyXJEtQ5zNYdSyuEr+nj98kDouXvmuIC+3+4nIottbT
F6p7vf/hQgNmClOH9n+87+wKcG5vAx0zy1C62OTVScdNUvg6bK4boufaduJe
gTiKoVU5NArtzxRzoqb8+F45MiILjX3QmRh0Qi9tWSrG87kj2n9pSTp+8t0Z
gyvY1I0PvGMuQRoLg1yhDAZmYI2/8l1F0i2lYafYEeSmMp7mbj+sZr0iboVE
jduzp2RiwQe2qKRGrPG+83TDh8rBGPRFSPWiWCQJR4oXpnV8dZK7ux03Xy3y
0vSkY4c+CN8a/sPf6GVGG+P/+8oqHoOzanfBISFFa0ldQjdmQvTlpC6WjZf9
ac3ad3kk+24OHEuajQLEzYxTcg7CHV6fCNRrh2RrjacEa3t0eZp67PsZrPrG
F2ACKqDljhp2rzFdCXxIusHAPFZvN2DUdsaCS6aGTeT93gHUSIaKijURYDGe
/9pOjW9e8x52Ave6LuT1vXp9QP4tv04knUSZ6DkRMDV9BLFIySD4iCIormgM
wbcYNK3+lDBIopnVDFvF6Xjp2PfYOL5VF6box0ByzrExkVIHK6pYDE9IJb6J
qm8nICrfvofVVIEPw0Jefu/nWfGb/Xe7+UptJqBhXzLRuFNImd6lp/qx8TAb
tWTgh6DtYYxXnn0a/M0k2gbz9frmK9gw/R9BPbKk/M/ulEBI8XZ0/+dDnely
mAfQ5IHZY2FasM+fogttYsahxTmpKr+BlSSiORI8RvpzgCjHK5R1+y6fNjqg
2r8gQ0uR/YdyLit25mzovdb0UWpwsYIydLqEYi1h719TWYF8bDl28Gg3AsR8
j9wWPaf++CPUJsohGsBX9GxkDV5gJewM1F4+MTgcd2RWpvIfpJqgNMelEbI3
sRKZ8FoEUlXHvbe7eav5NwNRaYKcjkB0bH10eCT2czE99UMUUJbo+Fi8NA0e
nnHX/isjyrmO6QzUP6/tUhym5NF2xjxxsUSfNknQ8ma2uMHoTAOcqeFgsqhP
BDzSCzZjItDiHNgk26KleYxOih86xFjt9b7Wkra++S8v/g7CN8Pm/MpbfpI/
wQdSzLBnYI4Fs3nsk/XhUhQe/gY/SVhOAhlpXVNIiEN0pqeNhau0l1WGVygd
pHlSb2jBkymuI9xSl4OqnfQoEihPqpn8KSBpA+IFEElsU1nSzzfFlgWG+4Vh
IGmi7q3CCDnmJUepmQrk8V2ZTwrb53QcvJvaIUVpUHjQJRi5ANwWxKt0pZlO
6WxloU79nSloFYmflU1SyVnx4REbcptSvVluCILfU2tYTNX8t1YnGRcbjOsL
FW0UYNo7MyEEiA+jdVknHnyqPuQlz6afkU8x+3TQLpDus0lOIQ3uPceFG/gX
w7FHhKbPpgPEN3dkwvTWNF+BH7dAtuyQ1OeUkT5nzvzrWDwhEWZkb8p0SWqx
2R6xQwVEfsvFVONTyLESz+ivuD0sE6PEEvfLZZWYrc0I2VJnPCvFmEj9l6aP
Gw83GWH7nZsMcj1I9upsmrl3uk8HDYJAgebzaILO7J8P7cn+XdS56sBw3Fhz
CjuuBr8kQWahGsYpYyJV51bPszA6XmvVDfPqYInH6qYIWXwvuX+VgL2j1BNs
ZFSPuzQ0tliXNoXElU6tl7iMA2KztddU5ZATljJpU74EgGvYsQngFsM+vsEn
0rgqFfFgAVFB0yBt17YArzU+IyDBAtFsNQ8yXdVZNqC1dR+DLDqja3byELgM
NwB6idP3M162FtVJO6TQmNP4w3pCkRcW7w8sYZGVrD45KIab+razqjjf2kl5
jhT+EhEsXIzxAzrB71g2u0ZXNeWcKs95Jk7vIy1pac2tv7933/umTpYeJJL2
5wcdDm074OnkM7hBaaoxA6IQ0ZRvjcadq7A6NaOs9f5hQgm1+enE1efMNx2w
3UzpZ68N3XHEX3+DI5rOb25nKAb4ej6e2r/gIiziqo0m9M3Qt7sJY09yE5Zv
1WAQnFVaC3HjTiyoqJBzaZP4GYnyG9jM7DebfrRUhtEQXyAxDJ56/d6dbDld
20mba/b6huPxc2AFQRM70zRyFYQPpky71rJIZOAROvXpNFrfDjN9moRvSIbB
cjASZlCk0VB2FM3nVgG7BtZw7eNOKFft3629fjISuRsyfkengHvGj0jdYq8N
Rr0WgFbvtXOXEh3hfRIn4Wad2lIZkudXbtQhDrT/tIGRehBiHarhmQj6gm59
+WLTFa4MHPHzfpfZ9B/o4ro0gPfU6DK5g3bbI1JrpBVIOxwSbLPwv5C2wD3X
f7ywguhVNpCLRZJFgCetW/pprp1ytHa+SAwCIRl0q9RNQccpHaTAS7hF5Mzh
LVwucOiFhRCGX9Ioct5RNVnpjunKpyFNMqMx7EFIQBRflo9CRxXE2ax/Qdlj
tAOoUrEPcePrquOItV5a4l9qTfZVh1I8BHD2K5AkuuuFJc3LffjZxLC1rGvL
urLKdS4LLX1a5Wy96tfa7OdjJhA3+ig3PYNCaD0saPayMia+GW2K/lPsF2fF
/dAJqmFI2h8HD+D+e1pTJnU+0Yr0odhewKdB6xhem2t46Q0TEn+5bzcSCsse
2NQb2Hk1/hq6Z0nKnKXxThZF+vqW+UVIa7rycal4yrQctXR+IchwpMNLiD1Z
LW3MNGNKPsER2lJXO7O+uCHBQ2mwFKAFpHy3gCwU9/7/AF7Ew2dXsCrhfsY5
UDlsnDyRVqf7ImjezG4VFxw+Le79TRC77aJKlwdo1ni5+wBg6vkegXTDpejX
7zO4LF7XNJYp55znaKdSxRUF5cRzbLTSWNqvGmivKo2YyzLl7pesruhkYND6
V0jEwneaA7eEVOObFFFRFAIub+5zHdaVx10Thmfwl3labxfgUBoVNf4WPmxK
Tv1yRovW+Xq4/vgc4d8X17IUFtBzklbpaU9rQ+dj2o+UX47fcERLk8QSbLiD
8bOoAdM6pRGzMHQ5N9XBJgRMDUfcpAzuc4yGwIP1JD57Awxvarqxy0DxEB3/
Cibp9qh9EATfVRWzBFxK2008kN31aqBcvhMOflOvrr+lcBe/1zPFC8G+w0lE
w6MgYMq21bAOiRY7P5pADV9oAgbG8kO8NWSd6bknyU6F6+SEvd8WD4yT/PYd
XvKNwZhgXckG01frGz70agZel4eJz9rUfJsY5M+Bgri6j7S4gg7W79HYB2r0
u+X8vnpEQ7J/tkxt8636gQT48PluDTsTf0tSc9LxXULYz2RUMBBHBfSUKSfN
G8tA6Jym7hZTI5fyXcw2/VhRcSVNAOz/e2mr6lDB/KckOc7BOvqMYASLWRJ6
3+I0IK7WPoM0+bbPKRjDOGQm0E6/Wo9U/SwCHOHWM5eL3IoUqqXBN6kDMO11
kxychDWgRlP7c/H2J5lz2i2uRkoBI3fT6kCBp6ySnXAsR9wz+tvNuF86SEdt
uPqYxcuICWOy8xXu9H/ZWPyg8sfub1BDvq8n7ZTI9Fsrls0yYfj2P2UskSAc
KbZSNYsPLQOG12usZtSUeMy/wq+e2Ttm66azgsS3ZrMFuOBh9k4CG+KC2uHW
vsS+m+m/CBudbmEVk6r7aZvlxaQxkLe4+uhn164iSCBXTPTP3p0MiUXbwgdb
csyiQ+6csM7xLGp5b6MYf3bIk3TPyoOAOL8I2MFnRtYiWIgLfr2bZvYF9M7m
Z4+tY932qHy1PWeeMuiV78UaxoIS+3bF4+PWBBCEaBzaLKjIjQZmCcyJAg7D
uZryclBsGLmG6zluzpMSfM/guUdf2rXzzQ3sSZRKpm0Dz4D9U43LL1YBKMZb
3hoyIfyOEEe+VCfcn9BwDcoS9CXnUGWFGEwKN3zIiRuX+gMkptBElqC/3rJr
hPa610FaEYE98LDbiE/Pkfn5O5P/6ib5xhCMiVJWE/VXebJW9C4Cm6xsU2jP
XA1N0Q+gWwvQAH2hnGLtRpgmjJ7mR5BPsgAB0zsuWVHAQw3P8pY4sAeyX/IO
7FnLz4Pgsm1yLJw/rLf+2PHCShgYwNYT65ijQ3Yiztrvtc5M86j5i3mRi1wc
bcd4OnqQki4Qge7UKeRNQTN6McNO+85OHvNeKlFxbr4/8dGXSEWgsYBGyN5n
NXH6sqB5tAbY9l02+xMhAokH4e4WZ9mPiUXfYWCmb4UvKBgsmXO+DsNCwM5U
okZ38IZWI3eZsnFELR6OTPlf4O3my/AA87gtsqrVeSpSSdngt7tYL1SyxTUT
FIW2dMP45TnyQsujz40t8lquhQpR6/76kkUj1NWvIg3gFMZNpimpykugZzUI
EceaZM4Etcb8kYswf2kIK3QpUcoh2+5fOKUwUNgb44eeXStQLf/sfbz20cYI
S/BhJkMfmrpLrcZaFRYdtH9P/msrLc2bm1ECwDMpwSLKSCLKL/RBtYXpvIth
PoGCAsLjgRmiSwrXhK3/BcIuKIWvOhYpPvSVFgif6fYWmbK20NYIP2EHcGBG
iL8CGHnUYeKyVUUhmOn8DJyrpWRaVbs0opEDFJ2QQPkhEo04l3GUcXJUnjp1
zdpY0PjnVAatEABRN/BxkEQ58QfDKQLvUGwWtAzimYfUmnuLHHYLS9WISDwE
2WhpA3l77jFzYsjipa/J9u+ok+PJnGS+igQJt7AN7H3V1V5ZC49NsQK85tRG
JJfxMNpNzwkH1UhApWpD6eIxrljExnMZSUjbEdGecoFLJygPB/9wXsgZ9WEc
Ie6MeJIt+76yGyb2B417Y1F+Lb5/J7eh4EjqN68T9vcf4zrqwkXQULLDGhdW
aHn1qWiYnUtg0iHYwqxVcBLhQgWjngpZXaGdmoBBnxYNwy9h0Sj3jwrCRETO
iAdV4SsTKOp0i48VnS+ZgtbzwsdkHeSdQgGbWKYLwniM35RZgBwXYFmT7n5C
J3RxfQCfIMUVHCJah36rWrQocCH74qNEweBHpPgII9nqhRaC/Xlsj+z0TdXL
kU5H8gNNfkqSTjH13qmjHeZ03bg1XXo1vEZLv8CpxZWCdDpWtjYFLM4llJQZ
UFwpnokrS54stbalsv3KHDgpjnvxr/QSCor1A0b7koDSpYUhB9yKqDv/yFe/
SCGpFFiObwxun7gyTu4N0f+zOusWc9P1DZwKGIG3ryQeySzrEh/E1ll89f8Z
BfslnIfB1KkqddWCFgGhwl4XMJ56/i/tE5PGdMh7p8vqERZFkZ84Xmkft4bP
k2u+03NHUnykHDdvszVSb007juxpdJf/eA7AozAUHCGqlg+L9rO5R02NRECv
UIo2IkBncBywdll5v7SPWfoH8XKvm/6hnXewAvmykokOd75o+asTQADQ2gvI
+nWu9UZhnJrguzfQkldh4tOtdr4btGm4q/swGoRd+L9/zGRYPasIH5IDPhHh
ogpsx1ZKPFMpnEukTOdRtu7lrJXhbDAUPbvJVvySVH20LX/Zv53MgOhEoqcV
QvQSFQCFD/DU58NVPdL1jUNCFZJIKUlqpDiWnQzfoBH2Swbu+asSlTGgwJhN
rjdrLlUeNs1jc/s0yH6KQ4jvCKDkyklARB8hAc6IehQOT7kCCgh7rhW67uWB
hdW657LHnaCuCb0qBlzIfj1qYCW/EQ9cDkuKb0bg7tjCvi9ruj/1Fl2yPiRi
lhXzHQsqNuhKa4Hd7GytyMtTxX1qil1WVvupYgR2VV4TAOhAojsC23aB6Q33
SZoO2c84BUn4M2FOxQv4zC0XDvNMQYxUs6wADLoQCH0BqxhV69K2hQa42Pf4
LqemPVHeWm3hgeLlBJ0ykWTzOrVKfJjMkMBiBbgexqYhEsLzyhiZYFKm8gQn
zcFeoClUVC5TDFzP31puzmFs08SyX2ceAO0ik4b/4nZYLUYNBxgnRcY/5IMh
nq0Tn/KueK0nFEBOHgptP5rPV7RVXRD6kd0q0isziVWybJld+0wHkgSN/Beu
KKpb7uqIXjqKaUG9QYH7ppLF4NxNNrbbZbK27SJ/kRrbuCm57qmK6sjdjjc6
5LM3QYYBvaz4i4AoMA+GpTAo2yRrsUKoKNI4ob9A8D7tOIydI+kuwwIj2TkB
hedh9X2TluOTMNUkrBGXUh82VLT3PnOy9jHOiYZggcfXgA5wGQpenSE9uDsR
m33KgWg5Y3QbDSH2clOT2JFjPZSHzGV+rs2K+wammTvxnYK2Twl3+nPhXPln
MewxRj8OTnvWUNu0ng+fxr1lGCVXwsU+mpM9pnyIy4FbtXudJkxekXQL34xY
MoWugusn6/VaW33e8iKAZ1g1GHvabFC2CdT46EobmisS0moECuVdMy7wIztk
HamANbQmJ8V/Evt1iiN+YwQzDZmB3E19SaM+QJuznX4czlWep4c2VEnn1EQ4
F0x4+NLR1AF7V4Nc59s70fv+eMpYgiCuJt4ei3OH3xd6/anqyop6Uxf75kIj
zdWKOYxzZWU5ZTSUJhCUo2UAf8hfkJP9BudpQ6+FBLj7TCRMkbMKD7YhVIUN
soabRW9FC2K60MSKFMPn4pnMzzePp57ImWUyFrsrG/HV9g2HUYQHZJwP8mCx
SjCtHFiLRSU4RnleoQf9gTk3yLcyNJmC0KYRTIsOhgeE/1jCxdok7R4+FAlD
dZLc+IEzsJXczQ1lSyZfwQ9mswVE6enVhQDG2lTyQ/N6v5xG8Ou98fTdKr0U
kuv7Afo0ZAVEgOoBxzwFmYjqOfsSI8T38gf0lPdVDtXfg+CjByEIl1B8Z+zA
cQTZz02d1X3RE3e07Hjz75pVGnuBZL3MCenrKF+yqnLblxg3ufD+xJoxonv0
I/cNJKBL0AsN6hCySx0awo05Tmb7mVPZopLuhgMebPyl8RQJtLYOFQKo/cB/
/9u3+W4EinBy3FYe83hDLwDDvmqIR4rW8s6xARVX6fmERvy3bP4loLS2ZElY
hZfGJKrmwDoRDsmfyBeZbM1GUC3d6itzujVi0c91VsvsViGxx9GrkHpFdMTz
a7h25Y22bB/al5Hwl3rzxC7SDVc/Qwuu8TklNGMqZ6NLXTGDJabsyxkww21I
TdRi3120Ph4wtp2bCK8In0zvpqwCApQAuIjKbYpPvY9UoeKHcOMiFtYr64r8
88aDxx50pUjIklPcX9p5Hyx6Fm3xkb+Z+CW60967OB69HpqB7em763jNqSKH
+DaizK7opeFNDOvSLr9pN/oZbDNjMTZoSyBYXP+KGdgCQ2hS4pyZwbrHKwQV
0rb3TLq8bhEcJ067w64HaX8sHTERL4AGJg35E5aWJJnHjwQf8t2SJQ1AskTS
4yr86ru0yfcbXgoO7FA6swS0NI7ehJZ3ezS5unSToSi+bf7hhKkRAUW4NDkm
Yr5trsG9G+HKwvKrVTbGuv7tg/V/yTlpr3UQ/jlne5+0gu5x/BhgoNWZCjYQ
wwIU6BCCNDz/UMfM/hTRiS0wI6NRyWs0/qPGt8uQaAM6pkqirGYCl5QXbCFR
s878Gg8p0wuWjCF41HcClU5jv0ndZbz3stcg0nY9OSJMZEOrUyE9ZinJivn7
qi9sWubpoKmGyDH9DYplQEZPmtSVaHEmmWjpRHVlmMjb3YSbxxV7rwYAQaEv
zV6qtW6NZiyqiEL+p/0FyKYyUrUA8fbB029PKD+t2NDYpJPY+Eo2paRr5/mX
H3XJKulF6cwSStmjoxhtI7cIn7MPo1/1PMws/fiPpoKK4qnqqV6Ks66WU/li
JpuIenG8PTz0uC6z6ycQptfhVCZeMRRZWOX+P7dKPJf+xPJ6/yEMXBMSh27m
neGJNIcaHwJr2BC19IiFjBZONQlcSYGJZrNUXHhRq7aLh4o5XET/g/jAwi5a
oyA/utRuEgm76uFOt5t2Lr6lSjm2vj51PXSEeewaXR1HLFAolOAGG8rrWkJz
LfYV6ZouP+outk32cuW8K2F8bTFZGNBSchmt9L54zn786vZR/EsrYfH2IfmY
MFtbafIqlz+W0pH7mnJuZLCd1ccBdiongQ0Vg//VfydFtA2rWqYcP6m5wrj8
CBiRR1Y4i7TJzkzhDoYRMNQnc2znppH1xxgbDqlJtpEp93aNM3zTW4f++vJq
r/MLsUv0HNTUuni5ooTxFNs8C885iMxwbSwnfXvADUElrAFpA+hwYjkm6FFk
cJlrj2NRAb5e3Jf5oxIvUliL1MpmrSIzviFqI/nyGpPEcB0YD6BIKiCjjwYP
hHXpsY3pwQtwULamKUzcQJ0QRdgzjJFVjEjR0ehzzFAAZO9Fp7CwpilnmScT
zvUw/Vu2CWpTfaD0NNsDLj0EH0wuXPxDwX8azxBNbnMa2mb6hzWK9BeimSNe
1k2xwDl8/wWw0R3ISE81hRCin9C3UOLKdLQQnQjJWmWs7paPX8IcXQ0aOGP5
yC/koVs3YOhAg78s0IHlsoAdxS3I8VhIjgHQg44T8obYAPPJ9GApPxS8bBHP
O7y3Kwd42LFN3aa+/ngU7Ge3iZ4t9+yILD9VMOKqkJpNPOlVsOSkwSQxg1EK
pqkFvrjtEvqlPAFl2/C6eWnn77GXG1ZA5DeawOnPSu/QJiQC7kkiTlQmNE1h
2+lfQSTODe21++L0Sx/ly5iguwwxJYJgpX9U8cO2/82ureJ9XGW4mygBwHmT
sRwllOQNBHQmD80Xv0cVzxxGwc/WYlkxOFrcWDUiCx3ilnv6E3nCLOwt2uYp
r3dW9vZgfDZ4Q8n+7R3HMHJMrRDbRGYFQFFZdI5aQ6F1W53U+zn8t4J4YnnM
KzycFUJ00rCnu63fMvIbn0C/KQu3CnrxSjJ5WmNqv4iDIa6+cB/PSv4F5D1t
Ew/4E5G9nrtUT3Aafcd+M8tTr71RtVvg3ubnQtEbD/sUWd16Rn7bO/oR4NbL
cL3awVHIURy50m7KHYP8UHAcyaCeSespAnK8scJoyRTd7fUK2lKTZObJs+JY
W7nIvVC/EPXCKZ/yS0O2iePjWzlQvz557Hy90sTyR8wLOUd37Ef6UPnwbdkg
IIxptcqekZ3YDDlibQS2LNNge9xtgf/LWFHwfdME+MOaWKUTi8050Xl1Ce0C
1o5pM4Z12Zfe/jx+CmPCkAeycbxHF0ILOlO2kRaJqXfoQCcW6jfZqvmrQofD
zXH3UN6aIlft6VmKKuhNQ9EyUqdhekcer6JAfVVVoyJ8Oc1Y9VZOgoDF2WKZ
ni+j7KWb2ipVdE7eD4uf34Ysd9/vGwzdvKZuuNK7DS4ye3/S8oGvbDWGfNMF
k4zkkCpTvscWo5tdYV0UAbMBG3VLr4ugGjiUKH+TDRLWSuPAoPqa2IfLltCL
+LTRaEgN1nGNsip2BaE15Q3imQ4khrGm4/X0QI0ZFZjj50rd7WLop5il5CRK
tRaUyNWkuozhcnBSA3wp0NSMZX9u2E8km+Ba5ezP7DQiB9flzdOalfe7motc
x8nmxFMiT1HCO3o1Qh/iyh2vhZFzaRNfwtqSQWA/nLlTeFt3VAgo6+gyTgTk
nF8ycDYYaxvdgoAYeFnfnn4AfILqI2sWYGOekPCQuzsy4wxfKnJuPPOr5xwl
qTKkdQVUXW3Rfh17p1TJ8eXyBSbJCqzfcY48+f6TR3KbzbIdhf4CLoRn3/i2
Ev+qfcZO3uX+MmkFK+oVi9SA7EU5aHTpG0yO0fFYOH4KtyGO88lUZ3Q8QEyu
ruVsreOAuL7eNx7Zu3T7tKpRbseN9jjoSi6w5qpPH8xqmEXMBURcE/mtUZiJ
Y7ZtWrm2EUUKXaaqNN0a9ZP4rFp1cDW4v50MWdKkCbTRPveFVsAE2QLo/zCo
NvKLwlNuJaFfVWkhMx1NaiNnjjrwW+Qetqj2XP292dWEDVIbdpW2PhYnNGCA
Tg8IP0fbIKbS3LNvzC0Xkkp05R5mmxbjxNuYs/4bn57RRdrAmuCJUUY0J74g
S4Tnp/xKoQysMyaIfdzMDEk6PnptaG3/VSDLGcIhWd/Zf4A/yH+Ap2RkJa44
5Jb/MpAlIifJOYfjVWO+vD1PgY75aPgie9337fZQpNfVjmlHcd0FZwpShIK1
CQ07B6UoyOy4VsXI7fDNVcjlo82EMXopReHdGi8m8P0fWKfXm+p1/g43712P
v+XQ3OaE78eup9yS4w4IHXjCOZ46jgg/TxI4BEAklfIevmDlKZ6BBuc0AXS5
UrfBziAGl9inhrfl36w2o0WhiN+hvnjbcDbTns15CpYedQ4lYo8KZkdTTgzm
IwRxQ/Rzidm58jwRGspWggIcS9ZikZcrQWouk9tKaWVsOgpNUvFSK2iJGscR
qwoR3S8gNima6uLZozNL+QO6+PD3lmgT5cYb1jetXJtTIbZwRKQlzYF4fcVh
NmlTMeRpyxySn8N/Nd1ddYrj/uOpzmiVL3fhn55CkMANY9wBtiZtD5LEaWWZ
xlEj9J0J4Hsea2QzaT5UtPVbjpO/tFkuMDIpiNzQKQm1rh2uQyD5VYHeDLfg
9J4wH0nTj6yT3HhdQLGRivX+U1FS8OweIuswGqGgDYeE2zdmb9CjNJ4OfH2E
/TafA/W/FJX2f+evT/9xPmCVQ84nuojkBptlxKAFoRGRynHfCRiPvdcNeBwL
Vczq1XvcBNeMbJ+2AyxnS4VeUqT7ELCHl/vrz0FpR6oX5+23sHJqHG9OY7jG
S0atMDo4kv2wBnpkUUGahEAwB17te+xEvaClIXibKYiaqO6J5679AkoFym0H
SakAqUyho3YwHw6RpOCkVv9/7xZw5LnbpkuJzj78VVsbnCrPf+uYAEPEIdFA
e5dVNYtWaQZSsWiS1+EJP5VR9TxvvjxIaktJgDb8nIhtwAilRld62ZCWhGn5
yAnb7qSw5GQjqxKF/7qOiHLL5FZZoZNgJTnALThQ7ZEUMrR+f1gzYHVDls8o
kePKsbG5yQjUPzbyPZyOyd8hXsuhvL1weouvFRyh2pVDJq+M60UmvdD91FVc
sBWtz4Ykyl72mnJzHdfkDlbfbDFFC2cDhy27szehTGG6o+S0bmIdN9/zwhm5
aq80r2hwlc9W3ShPmlhaUUvec6VUKlqvV/UjqR9mZOgDPQ3BCplnQytJ2R+U
ThIYZaDYPkHPYHCTwtUj9v6ReJq5QcrYkcJK36zNmnOfjebChmWR29sRJ0PD
KK80WQuwCZ/pg97sdn6arhxxi7+dPQk+QVEZNU43ZlWzim5hjmk00vNM8d9s
gGu/R4yh/AC6gyiiS2hflFl5K8ORNGMIb6QjGV05WvszwO0gdqntqMPwsyfH
VTbyeAT8cZSSaPhyne2onsWGsfc2FAdRTIS+ZS9IZ6Q0Qmyk29DcPAipmKSS
YDgxQ6duXkls4FpB/Y2GmQBVQKmIf+8QWv4jA645haJpaSj912UpCbSdB6he
qtRVVM506zteIdARh8X666jt2Jb9QKgqhOO8dvS11tfgOaeNXUHb4Uhgerhs
/GI9kOogq4AZtqaM6CUi613oDo/SS1m6V3hUi3OlVDmrDMtPHmhVeWiIu9K2
UttLDSoc1ANdHPn5uCCw7sazWrzy1c4Y9rLAcMdNh8NYpiFXiczN17C6ZciX
zAeVE9frAc6o+n2n19/fCByS63FINsppmIld5AgB1SHUasodRdX+G8lWHlOQ
5r/jf1lySOZHWqyMwU2x/w7YNt/6dwFA97JHiapvrEFyN2gqHop6/kGWjL0p
7LjoCxdK/VPR/2XC/BGIXMpIKSOA6W7PXQOZqLX1IyscJbFpN352NCb5m80D
ecBFogI/cEtTRXR8IBuFoAy/2g1tHsWV4dbkDP6DVtoQmAmm0aVfEXYGyiyv
EDnPOf2Ag+3rmadLgqip+6S/s6KH6eEUNyGB/T+osFSYLe4q4+RYwSoWSUmd
XlqTxijTgstuvje7UQ+hiLPvlVoL8GsMZtjCnsohVn/cMjjYAfRpvjTKFI5f
83j/XKQUVfx9sNqykwPNJrOwUoCmXWljWOUHSnwFdrc2Ei2x9KummqS7jEsE
YZeKF+CVXNNtydU80kTKjNFo2sam9N7NkNNmf6r22Rd16Ibn1PYc8z1boe5y
pgfGLpqr4+zYDQr7YRlg6JbCjz4i4Gadkrz2xI+nq9YK//6eOKqQfrnDqy6V
YkkqrYoID2Y4s0uR12l5H5kEhsuWUX3x6PjbCNG4kp9qSUAAb8+6Rl//aZBn
JO4liI9t231G7VJwLp5Aoxt17WotTlmsV8pBoC/Mf9KBYu7qcbnaRyHX9eh5
M9E0ZDsKvuOkptpgeTu6KKNqco3kuY9mprT4WN3pO48E5A7LFQzHIHzdhf3K
ds/qBZkLSRPIsBJqyJMZr4mWrFhw/7kHYGotYdJ+aLrFGlhC8FbFe8gYWmc0
69WSWiuto16j5Lkz3nqXit2YGR/MtBS+CAbZvZX1qBxV6mF3v7dwn33TBV9q
yepW5w5HHS3UxDVRAqYR0TXsWGuCOn4JQVA2tjW5lLF82WiNrOGfSVn0rz6F
llVeVSIuK3RF8h8MhomKJi0XH+gWGuQeOtuR82uoaA4JitChoWXxABW1OrQY
a8hU1Gn4rO6L8Mv/YTTkBaZR+cuUjYOjBlOGtEYxRN3KraMsDfK9IDFqiz9Q
5tLbsZhFpY2lF4hti28ZGkuScoxtlIGL5fUxyftcFZnYZ+/208IAikXera80
fxt1Hj1jAd/82WryQ7sQKEvFWXcFvEliXTnFm+lmHUTNdw1V0C4+ituEm0Gb
nA6skmjf5/543oBasUfqtKwbuA7oQXpBm/CnNsqkAGOrJ97Z42sAfvnaScs8
n8rO+wbCO0nu1kv/TeEq8ZWPsjb6KOZA7HY+iQZLjinEHmB/soyJKT/5I46q
yxQukdHhYF4OrpmmiTcWMmTS78vymtEgsUtzhxhk4sEKbtLm8rb+0FBRk1Sn
rpcAegW/xiXQ76OlfLGj6+YFvGh6yJ9FATVQWKEUYlFmYH4dXnlkjliJowZS
QmkhE8IavXFLOWykimXI4Xb8tUkHODpi//zaUDBLn1FTGePLeHPN2BkaxrJG
Q953Z7QnDN58Je5L1Vu37qP54Oakb7haDn9yzfmy917AsiDNnmlhxkN6Mkr+
GudATpI3KnQ91iz38xu0JDEXHOFtIAsdMoKAX95vo0sRsPzvwDkeOF6QZyvL
v291L1jzQsHJvDIdV8LGwypJ3fjqPPR0J45E18IClLRVWhFSmNf7pyhrSs1J
PmtXXLp15Y7bcng12GWHbCWemxwF/Dm9sHStXRDSd969JMvUv+pBpCPSGKUI
Q7Da6+0sku/SJshUEIgkdTQMcPUXzII9PsRTjw8uGAR7uR6R6aS3mk6PZs8B
ERCO+B9SCSL/YR+XhEDleGvCkMDBVHUeKKq+HTYFclr82+PrpFzO2AFhw/+z
aas+All9ht8q9SkZRgRy/8OLiABGUriY0VTAq2nFDcp2ZBARBvl+YwWHVBNR
bEUbpAv7Tvfj25t/K1dOi83zG/aWYZYgP6YZmX//dxwu1ZqBmWlXiR7leBvF
oK9UPE7B70l9RmskPCqc6REeLbUV3nMwW2dJH0DEPrkvTsYlyAdxHP+kDPLi
C/qRe5K03/RQ4MW/b2zNSIsYsnjtJ/d5sobgaS/u6nAkEMJAkruOTMU7um2j
LSv1We80qWGos8UMgr3f9H2vyytb5H80a7x0hVpJksmmsgtqIogavKpdGqCF
+1cojC3ithamD8ZWcOEIGtSbjNs496JNBOVe9S0gkN+g7+/iRe1CReRbYUyj
E5oYKHtdC2gB75jeGP+lh3yo3Xt1mc9WmvJYgFp7NEm3AYMVz5lOIh1UEHrb
aRH+rKGCSeteAbxlw281qDoZDt939BfltycY0ELfmpFbu4YO1B98p56E3Qyf
OwuUnVLx/p3qAbpjCtlVC5jQOaxnjEIv3buqImILOMupKiN7qS3lDnB704Wd
tQWkERrsnGQwYoArAfkfQImNT5dASIPznTfOxlR+l7rxpeDniPFsxFltJelI
W75DFsoA74B5EvLWgMdNAb6oL+QcRFnKLEIXx1n1/FBphICn1eRpFXFvZfsp
7Bvia836gXbDiGdJiZX5KYiktmZ4Ubp5O7muRYTIYD3OqkCCghf1Vdc5S34D
EON9JNV3COQ8DlJRGMOhFIwV8E4xrfezLykPaRyTCeYyXAR0cJOhew2T8JfW
owgzauMeNjBIChxU/rdCwf8De3/Pf4u6ZyTvzmwaFMDJW+X+aVhM70/FJpUU
F528nJgrxRnriBfyMzehcZhSK0fnoK3pxW4x+EjepiRuT3oRIL3j2YEGqRrx
JAY0eY/6irQNf9R+HQ3Ke5rlz9xO8VoJ57crsiIPn/uU+cscgM2phYS8l4nr
XPTroi5mKFwRaMdu/qH2QFH8HKyEqwypFArBhTEF32jACh/504mFctf2ZKvj
SIByzUv+3i+WCY/aSuzUsnZ/WmWKDQGDOI6RXISrGrZMZlyOlUv+vCayRN93
qO3zATCCYR0FBbH8O6Irjed8iUxPzjwaesuDls5WVflVbRqAov7ZvmEdVeFB
TazRkqTZ7/2niW6T7KpwwqKdtO0pfd0F/X9Q0jwN1jVI8jGJAJColKQY24JE
lfcE/Opz3hvT8MukkUREsGE3odm5BRp5P6u+LsM4vyKVtA0DphRDQ9dTjxcc
/dOjzgHUVym/NMzoc67/dgXQ8hfNcAXR68HRumnPLv4Ty3If1eD7+zG7Ekw4
Twy0dxDLh0qXWi6pmtmuE3Zcwp9+HRqr6zAMwHjruSzkxn4GzGk+r4t2iof3
9JmMZUQ6XurXmEVDMkecoYTf9dnmF73L5NvbiYvaf2G9U3r/M4U1CIika3xY
PzB0GWnV8hRXByO6XbFpt/V1jrvtPk9+DGPDw5a0/6VzYNZu5El/cgxH7q9y
FL0dxtqyY5n9ZGiz1Pgc324P/yqNiFRjkKd9IjiEbDRC9aYjtqiLYhdBdbrQ
8Y6rJoiuGTMREdLvLZYd58eDcx3gIdx/0CWKht2fdZF/94gsg/Q/Hg9z1NFW
/ekChQTrjBnqXpeMa2utU09FU0K55pt1pJofBnKxRGT6vIDtx72U6eJlcLsy
H4KfSbQH07RMlD3gCdFEtdXuqOAuRpCbSl76cDXIc3w7yvF5CXNU6iFQgAnW
RVjfWvFNrcbcQvCH9sv8mr7LBKIrSs5zqytpviKfV8OCUjYClp7ZGnyttMkY
fQ9mdnbuC71/hwGd6xbR52Jj/DVTB9t4uvU1QdJYhWa+C4649BTuMX2FmOfp
KFEukJk3N+i35iTXCZzcfa7mIEYK80Vco/A9T2wXax7DSQbYvRqvuzKqTwEa
K6m0ccuJzD6uIdhHnzzpwZZNVlqg+SvRJJfZ8E1Fs9l0k/5px/cothKrvtSh
fzm/+0O3CRJQAm51SgkSW7ujbgc9KCE/D5epNmJqiGXaxb6ui1aNTIdTtjF7
L5uVfyN6mDM8M8+AqbiblaKMyt0zFcQT/6qow0uXLn3KUnwFbaoA0hWCym//
lJYnt+b99Vkfqizhxy1zLDYfHyxklamUJCLiomGiDom2fj2Ie8Gm0iaSVE3Y
8/60+1IEEFTFoMQJi2FulPRtO7D/EbUStR7IhgkW+TjBCDiTRo3lhEe0NAde
3PAfc/4ux1YbR7636gftRl/+QTxL7FRovn7ZhLbiY9znFIKl9FSrSqKEnLLT
9xHKqA/EiBD7uIr+hSODqAzB7BrbkrFgpyzLzKZIacQcfb6MWiKcDmQ1+JP2
+pbh3PPo2XNyrg1nt/BGkF55hP9/+wrj7jmKeoWr85AeNx6moVfEdmVwq5sI
hZEGDlIvZFwQ6H9XGI4plwxu0ZGC+T6SZHvE2bxBiWuyDWKG66hl0Ok6W/iH
E9smQZ6HKUgpLdhaHETSNqKLIqQoJLlKMla+C7v7R9J7EqNxWDaUpMTY4k3e
IaJeTkz52TShfN9YLDQLY4KyMk69ZjaRYAW526f3yCI3jr7JrmQ5RaHSlFU+
aYPE0KzaEIXyxvdKUjSu4anDC3gJnhJoc6wgJ0Iy5Ybu58PKUfeWmwPZfO+k
26XK6sNciXjs72sKIkZUsGibQv78uAdyA/xeHLaCyIzA97iegMl4kD3gpelA
D0mEbz60K+0TnZDJh/cleylUH+dXwmBeaIOYXf/o2KHWEzkjW9ElW/EpyLex
ydxMuaJchK5uwG2GS8vsMfmirDrV+zJw93hImKvtT8oOX0Jk7eKfLgXbJw2p
NVhM7hE97Y8XsI+3IbnEB3REqbt6lG5ssRxY9oyHf6qA1xBN/KhV2mkdtKaI
ANtl7/qKf1jt+zVzN848XULx9OB0R9QDpk6TaHTN2qBQjZcPnPEH36BLlkig
0y0nkyyGCA4e/vPd+riwDhXa7FiocvkTUzr5VQqGobPqxQnyv6RG49SM21lZ
1OWHy7c63TMAErNNQXxiSoVLnGuYorVrCHt03yVht8B9XqcBXtEfaxnyGjoY
9s8Dwm+APDlLWB/j10I3RWp3O7Z+GI+bHxV3Ti+pupcGhcL0fXgVv3XXtzkS
iBHGK9yXeKv51X7K5Yka9S3tzHqO76zfGj6mq94KvRY75Q0UMxDx1wkLw8Bu
2gPLzYMWQtM3BoP5SGRRrvI7561v7B/g4FmpJTxsKdovJ4lLUIQsh407LEn/
/U97CqQ636tVOwH15PjkUJUUuINeqWJE3/E4CDa446+qnpAC1N5x4gEOfK1J
uPmkfC852A1Sw18daTbBoRM0hul8Tcb9NDEhLn72kDWiz21ZEZ/fK9OVERcH
hyKgxKsv/3w4n66zqJ62W+y3jlDITdXGFsKdDQlzhsqcN/lR94Dgkon6tOTe
J7x9f1tzTBDfnPHmFUOHyDr9o44ETVSG3sa4DpGoZBFVreRwdk6xCu130+Ux
9o4gYckqd71qvg4F8n3FuV/tQOdrHP3SpZzlmMum7T/sQBbI/L2+zXPof0Gz
h9OJTrruSm0l8EEtXIAkIMjvCGTkJ/CwC0m7GCMB3IPex/v5g1PcTi9kMSXC
EYJIEycMbh7cQ3IQ0a3EWCzGGhCdXcP0EPAwr03ydnaiikc58tK6zLPgFvyW
Rx0Ve+XOVyZMvFx75PpZZ+Yak0WrEDguv3Z+eN+R2ltqA+Yb1SOlypN6dydV
k1NVz9ICnTnCGui3MP2YC9jeA9fF3FAKYJ6g5RJfBX67QHJcJkDLOlse9tb7
vaEhpyA7wINyxA8IWB8kTa+WakJkEwWM8s/1wK5Sa9niKkkyVyxHJawt0PCk
/EJTA5G0rTEQ+F34w9IAgBXWnEkzxguC8D2B7Q7aecbLRaHcD/NGA0Ot8uU7
Ap268zSgqHUXQAfDamZKFCj+PkzXmIaskwHaV/rc1gP+EgXCCcei3bN+TwSE
vXsr4x5nShgGnI5of4txuOMF4zpvwIYBIblVHSM0EJwWGBBsFYRyzhbx+t8Q
lGsomF9qCwot5E4AX83kncR1oomYhM15MnN2HdKHUHutjJS0AeAUbAnfq8Tk
er9V1S0ijEZG4ej3cLiWnNay0qj1bHaVnnuj0mUBEid6kxOlS7/UnzNmxo2J
BUcD058dKSRTCqCtFMvuhtZfEZWxnpju12iJjy0cqfsjFwKZusdQVYivvihE
vS1hZoY8CuieLBMsDzO+RUyvldPtXQD7J/vknayGhYRdzcrpqQPZRzy1bSC+
Qh309LBU5eyCe+KFy6UISPm9aDuft4nOLmUXOBpJIGxNp65qcF1ODStONC7N
udJWYsKsnJMalkfJsVqba4p6iUL7UUSH0p3h+LBVFh9+6oWcEoLm/zWf+Mvr
RKC1JsLJ6tIKgHeFtGgVeyNkdJLm5vuJX6CP+1W1i2inHdsLz2wQQSzPhxhW
XpgqPnlomf//S0lZkxheWubYJqgF8evmgAfoLFM0u6b7tF1qAUrRb6Cyk0gV
uT//r1mFkMUw9StoLssnaJ42nz6mnNWYlSeDsAc4l6kHqmV+EBfnz/w30bdA
DxXQNrQgcKxNV55s5q9dJZepIWXQEez/ymXRBckVSrkWsUZP/aVh8tyO/b1o
tkqnVbTuMWVMItl9WdScoBEKboEpQipX5ibB1te025Ap9xDROhyfrp85zPdB
Ma/jJMYQd5fmSGNgi1yomSdjbgKsFfRk6wzlrTMzbjhfSqzDV9ciVyE8VQ8K
iBPSaHAM4SKPizodGGdnOGMEORozv66EbukY/pq7uTGzx6LIxLg584whyJuW
t3GAxFBmKMskcUIU9emfaBHnbc4STAOlEl+M6JqDQ9gLye7H6/A5PmibNngh
pztVne7XBXErfl4J2ysLF9XxxqLjFE2ygPfQSizjHUoyb7snh8eKNzJHXTUU
gdfJxbll4JlRa7nVCv19I2v645szxiS/EE2QOjF3SANEeZdkHxsCUH8+gFoL
vhRCFjMlldkELLTYKU++odp0OLDZi1jilD0ecDbSd/tzAqT8bANZtaC0AXpB
RCMXFiRFldcHZKOCxbqfH8tOiT25ADOJNLXrOKcD4ZqBmrVZoL5OJ8MdzGzZ
ATPUl62tkbQw8YGLMcgC0GddpDzBetbi8F6xl2D6MXnergXEmGZrSP/yHgTS
1YYUxw0teoaiXwQ1zhHTCHKov1sTHn2KnXGBNl0YrIikOHNTEVzImr/HrO73
yMIuvtH3WqI8VEd7Q9J9nrOY/EP0Zjn5qKstVJtvVKTvfpDNEsLkpmp5BW8w
hqXs/92UBaxq8hGYcu5fzurb/qOhcHG76tdekzI5IgJnQC7tnnu/epqA4WtE
FydpUAeLAA98fbpNiDyoQlHkoC0H38khwu/wlXW/B+zXnVHfAjwhBpiqPYyO
JNO/8U9Iz5F7Noq1rAuaMbzBPJI+6zdC5Zzz9ssKNEV5EngscrEn/YN9nQoK
YRKykMNvph3u9YcMsqXuvoLnnZkivgDWyGbrhSK/5c9bL2+7Pi2QpVXXZY6J
67J7J5gQtCnIZ8nEGD3/HXBEm3kL1ln6mii3gq7Trfb7cu5D8j1DYUFl/Jrv
Fw1eg5CNFP5D2Tki601FN8JO5K9rKEzTiswJLJz32XedNnUAwmJUFBDSjBu0
Ob8NgyErhIVFqhH5AulT+7P4hPut9EFJXOAgcI2VHK/3xQ9F+USXK9rn47yO
5Mw9hKIcVrHrJiDaxcVat/8FbnvLW0gx8y+1JOpWy1dPazVdcRXn2lYI3G7T
hlP3x/52iZiaKErLbDiAyIi5VII40QuQnboZSOTreprfYCxnMoI2qAbEiQei
/jzzRSpYxr3LdAcypJjc/KEVEKw2M4iKoRFuhx5hR4o2ASlbx8W4tI0INPSp
0PLytA/7qhXvIMuExiHbKVRGzocdeDLs/IY53AaHraNYXAapzngTkDQYPnlj
KwwJWr+lN8drx09hdRvfw8j9ZyJJKD/fMzOYTGKbtd9IEZyHL49McO4qtiwO
R2hsE7gmO7ZtrxBucGxjLkCdy7+CjEKobkKXQ5u1rm6yQyXaf+GWCB/Dq/2F
AlbHtT0u0Bswx8LS76f3Kv3MZQwI5IX/bGAkuVSOKYlRvZdexmHVlTqnRIrs
4wZeczBZfZ3wQOkDNDdzc4FO4dosVpTeiTYCWKOG4hVM1wvgM88Qz7/XcsUM
Ubr7u9XZcWYwxoA/kaYpzELB2+SMQCi+KZpjG5FB+DxiTRSlRlJWgBvxZleY
cQ5+CfygUH0CkTfXq2XXB7p+XJipbUAVGGg48WmmNyeK8AhZ5N0d+2Qpl/iw
Ph4WnW3nEv+95Tevx1VAVYHieRJPcg+8njaDXaH2JbLa9iqUQE5w14B2Ik3d
Orz3Gmzjg5O2BmWcAzGKZzNsG5QHrRI8usRAsHuEouX1X49AI/H2YDs/DRpQ
4C10PbZqGNImMMj8G5HFSXVD8a/U2xT/yol5E9OGpIc1+rMoX7qqgkLwmchL
NURqKPtsslQqNcNErbjQOrikwDd1J+WFyqW9xDf1N6iF7iIaOIjcAio817G3
I3b5qA65R/tuU4FwYus48mmvvgWQs7sslI27tilXuf23a6mpTMgP11bZZJzc
iQOQ1goz4oUM+CcJY4nMG4jr2u5CO+W2LvQSoYYoXRndJSlfcC7k+IeT052v
BxB5v+tTdLyMc3uMuyy9j366mwdeONchbTKE5pQ7O5tvZ0M/zHR69wKS447+
nFPlCOASj/xqUVccNUBepKHjxAtdNVoP17gKAhF2Jzs6vvJ0rvReTmKBE4KY
K192OYDnpB4czMQiCVWnTLM3Q9y1qSs167S2ZY2lF9fALeNetLO1GG6r9KBS
G9jkXiRbOX3cehB3Wy8YY95hM5PrLrMXN3QN0hWnQdGzmjrBvmtTDSUnpZuO
743HN9Gofx5rwEgggyXEH3zPY7Tmwp10eelGTUZeRMKjsJKCIEs4rjeevJyp
G9kpx0M0F9X8HdBA+EEyZDoTZEhMEWbU96aiLnltJV0z0AO+JwAqZYE6xghR
+KQ6v+4WJbZNy7+kXyFCrX1fENS0nVMy4ezTQw6MIAoZbBi23hyHts5vcdCb
nOwwY3EwA6FlQ/zH6GQJgG+OYncW0sdQVgbnseONXeqo+ZS6Jdpe48p6AkAm
A0MuLD5H/g5dNsNcKJxame4PzAlfhuDbR8LG9UQXKFyBywWpkE3jWIXnvPuu
sDIHVwxQ+Apfwja8N5SAQNj+dWPbgFDykfLxViq0lTbvB2ySC0a6f3+DXee9
RPrH00wwYsm+6F4LQkAWsqdJDlW9aqXB4jsbZttyC+YyQG+PGgqIxUCS3isq
iNOW4v7FF+mVlQIffbicGcNH5BmU+7xZ8TXfjnHg7mbsgk5h4XcG9By71LGg
1XqN4ppeT3pTTfAHu6aifETBjHAZWFoaqqyrR49kcYpTZ0ehydx/Xr4mmBkI
W/k8rtV1aV0qh4iNQk2kU++k+rtnyBg32cu5nmmF3kGwNxU7BjxIdpBmtfU5
nGeFD0mHbnj0ujJKqGuugMdAkuq2zWCIinYOScUwfb2ITslh2qxuqiCKgawB
kPzoTThOp1WiLfacO7HUSoR5y3TvwSpxp68yuSkBtap3PpeROLIDKFS1QeCB
TSHWcasS1TebMqG/9cD04rRSFxgjiQm6KZALWPVFFyNaOhw/3x7O8I0R3xVJ
SmBZvW65YlZyA8YXNgNRVcAynocNPljcrrSS7HP75wlQb7Y8sN+c9U/s90T+
vh/XSb95KKV8ONmiQMPXaupSdHTzzz8K2fV9M6qNMiVr08eiyaIe5y7zdEdd
HKyeTMnyDfEKVqsP6r5yGj7FmWWygXbtOiOGF3swYA/2MTRHsMv0Uv0wyvcd
NQ+pZQnBCwqNVUIW1MynKFSdGaaX03KVrGuKRg+Le3iAX7v7G7XAWKnqU49+
/aL25c/TU111yYUWrnaXjHZa+R1vS6l90HS+zpc9Db5RXoicySphav5efTIQ
KAIhlAXPApGBkQxqH+GrAoeyTFlD26KMennr/tEBtqtUh06AdOoGr2SsrWWc
ttwLPAkHxe9TP5+ZITFwO5CK/jhmwBlBlSSv/Rxpdcl/Xd3JxO/Knt3Oy37p
YYIKvKc9fSx5FJMaAwLoIn+504XKlprN0KdbdiV14zrf3Lk7umC89P2Z4Cr/
phHsaHdwm4/OkhRMBSBg50uGPDkNkVIF1aNOz15s5+TcWtDj9WHDiqgYqHsr
Mvi1vpMHjbzbM4QAUG8qINfFIL1IQL0TO3S6mHB9ILiShSpRs54LZzEigoNb
xQlodLAToLkLyIkakxFt+SwrcgTVxjmq8T9yvCZMAr3dWkK0l4D07wbf8XtY
GQTFsV0VIbzpqeyLVZ3gpcp6S95/OoMgaDGtJZeI1ov2ai/jVjFUPrG9rJaI
UgNP6goaYp9z5bWfiR2IP2JZAxf7u0fuNaMhv/eMaVbgunaZ374vUxkJTwBG
8TMl2MhyJZlStwDugTJWB8oDtydyZftPkNLg0RrKQjeiJlABIMG0NJYJJYVT
rsGA4dWxHkiyjaMsJ/vopfhszNhtEREsS2IwN5wyvGEzoYyC4eHAppiDJGWt
yE2Oq9T4eLdYOWPGh0PTXhTAq8dVQzggDDy9+5ncWnrlh1cBceksrMYSRVrV
UQIjs+LmGmNHxSB90TxMXecIYrVTNPnKrHM4Gw8BhknFIzfwkfAQ3jaZLPh1
S592nh+NXJKg596XayF6jg90TOWjr3x5HKKFkGmUzBQkmV01co60pSkWDRJU
5KX3RIz59MMgSWYKT/16fs4xnbDXMmfHXZ23sAiwSDSUU/wNiCLr/QL7vx07
c+lla0JARDs3kUxifYdB3xinNaSdPV9IbXOhwrRDMbl8hYRiu87740q6lN1G
NFAHDYR4evnXOcBK9kjCWbPt4xlfvgwFlKsV1LG0VsA2Szidm01zE/V6t/MS
ghOn6MHkqUJp7t7HjyoUwzOSJ32foOnjo0eHChf2O+BzGh3dsDFxtF6xXHcF
h3UP2AiuRLK0kh5/quxN2iy8Y0dPFgf9zTS3l3KPjF5MRRRRdQ7Vadvut2bn
k409cv6oAGRf746OkUBw6mruGplvpWaP01SC4Mceff5LSbIzao7dIxJUCJaN
4X/ObJKiEGIcqksVZgkRQdnE/g+j9CGzHaZIdpxWdQw2h12mmjKR6A9/SwE4
xK7JEmw5cHN6XBv15NdCbqrcK2dwH4JRysZfTKUV25kUV5z8e52pKSdAfbbr
gXDoRWo1/V8x9Qa/6FczoEoDYQPIxegUOD4a4XKFOpmOGFM0CD42eqNlWABa
3q1IulqCJNvYbcckxEhTJzmeQwF/0NeGXUujAvws7n3vjrVg6cBoDAi3XtqP
SHSGkAoa5d1XnLdgIg3vBw295uPf6/WJDsoJO96EVpoNvNjZPMpkcNBA3k4a
QxcT55+s3/C9sHdoTT3rp0NPdAY0E1uxM+Shr4m2HzT32KU/GkF7f0YLypTk
+Nj+U2iyQmYJud9CO2iie+eIK4mIZKVwtswdFm6KXFG3+p6rr2d+4iNaYOcx
1pJYRbt8hYXU1HCmVW+ovAbXNOhKgs1a8qnNNWzQwfyy7VZToK15SGBz7s5B
0yetQSMEnaPyHZ5uMibFK/D1DnaXauVzxUm54axmXAQHHa1ccsk0jwpfm9qq
eNIV+SLCfoFqs0fXJZokOSs5HW/hqKDAPivKFFmjSEuokNdjULeK5F27anAW
BwNyxsL392l4TU/3qQmrqfDRT6rGHgdix5rgpI5bmUSTRZnb10UavrrcRxlm
Kdo7EqDVf4PC17wEgp0Qmb7wcyDwBjCtsc0DscsqriXbk5nTLGIOxFASAvOg
GmLIpeSJE0mmWj6BRB+HD23wM9MiJ6Yf31sPMAUuDryOJl/UWv/1UXHKCpj0
JwDqMU9FkQb/X6/8nf9km+QVuCA7r7g2qFZc4LyRrLT0yxsEAhOYTnjCGQIm
SeBiSpZsBIyd5iONChC9VQno5LCLcfdNnlz2Lxogl+lwd244Iz//70BWbkuQ
Kkn5z9J9h7gRG67AWNk4vqs34CrLf8hnxakgj4fkSkYBj2o0n+HCv44PR0Zi
sxn41M09+h90KcOaJWaArdDUcL5GGwJ18cUNV6i2Mpm56/ti5mXiBU9+/1xo
PrIBnNV2f5V52+Utr61J956U4DQz3bGAf7yn/5WUClhCq1Pm+oFu3a9ugO9O
vjT5e7kJf55n64rrUe0sLVA5241wtGaC6HgtsX7QzGNWJtEvIKFObUE8QYNz
PqiIAhHKYl8LvSbIN/JDMaiTuwdk2wPS3COdIaqrJDAI0VM739uhjPEoaMn4
Uzni+6I2CD/EirMy45cISLuWSSdabTNdm4p4XA5mtusuItFCWP9lGQgD0Rtr
wdPgVRv6YwOiMdcesY4MyxqXabbJXS3op5xH9ZpZCRySI9jI9N1GZItXo1+o
TQkPsFiQdG9wiuMhwNCr9W0Rfdh2ae9yShFK9QSGa7lPEhB8KZlj9XhvPau2
nKXxQE2TL5Pmy2g+O3jjazzTtpXGqectRl8Y/3W4wKZ1EUnvAWVeJBigOwUW
ydwaTZulCzBnC8e/mgO53++8Xn0fe8sXZXiA8dxXuy0Q8//BK8ucaAYg6LxB
JfkI5ogoNdIwh98HCXRaJEwIl8O8pGvnGjKB1XxJvkaTNE888acpotZo7+7R
QWjG0XlXCHSPI1bYhHMkoGgcIyukQpwRsLDU2Hfd+D36B+6UGH7dLIKeFAOa
je7+9zV2nCuMcdoO/N4Yo525uK0HAyZJ0T8SoWULYmv/GJugK7h00lNmYh1+
VKRCmqzKgRm3r4j8Unrzi1yhsnaHsqvys6B3aF80MO8AdhJNWtQrB+/1g8sd
SrI6UrmmAZ8OJSTaGbxHGh5Qe4SxJvn+UKz1iY8DlO/x/JerZ195NMy/Wa7u
QOj8VAsIUjvuhiOAdytthSDsUA3O+ww1a9yNP8OxRiHeK62kDOA+AW4qcgON
HqVeStL/7gWb+QYFdDzvhjQ+OSaypOkv+bQfAmEGubLyDPevMCXFTqPxtAJ2
RbAfzIdyHhtPFb/ThbgEE/xqOc0Os3r825T3byCRMG8fejHY6vRUo+25HYMp
XvKFtKAu/oa611+/75ktl7QXHFGpUmodJPCD6iRzURzo7DYFDmSuO7zk68nb
yKRxM1f59pMO9k3eAxUx+YYrCP5dZHlz1HgQ6dueIOoMEyXYk9WW3mVvK5XB
8VefalvuAdAn+SYdnyR6IxCNB6jcpV2DkpGcUfewHtmAiq2+fG+L0NfEzVEx
UBPPhSzjLS2mHyK2qmjLDKkxSj1RX0KcTOLMYUZmYuxp4FAkj//jpd7fqPwp
JNBKKhn306CDkft1Dlog8et4xvvL8vKtfCGdDY2WR9GzaM6aUIBTofddyeTL
2WS2idVsQ+q1h255Ltbgqa8vA9UAM3smSOgLQ4+UefNTfFcvBKMURVw3UTgV
f+RA8S4ZZaToYVfSs1s4bS77YZk3qraNmpQ2oGIpEewL4meFIbElIP/gLpK2
IAMPj802ukgM4ZBwQyhQE0aruXHBGHhp+F2xATVu97WmEJQtql4hntGMRo3B
u7PeqRDL2qKaAES05H1NgTKZurlTEaskgSIrlLDlWEPlNbcnh6IedfLkIYB/
WH/cuSa3Xul6OIbGNje5iTzdbJMHN/kADhB7kA7TSitPuzacdXaiXaiafc0N
utjaaRHi6gZZ+l5Xm9tPqQwfkb9YW7/nWyMS0bz3EgR+d4mSN/81g0L36SfI
gX9WdxN5SIKtt1/on05uECIYMgv7844BNysJV8I6c6QaKn02b/iBXwkfZ+oG
Wwe+0qrd6pCMgh43e4BYDf6SLhVORlwvHd+aeJ0wPjv1AiFnyFH8jW7wu2Wn
5WfUePe9M6Ixz+4BUPXfDda9FkXhmeCrwJxXWHivsrUubDJa2ds+qwd9ZWqG
3egsK1qFpqw81PG88Sac0rn0tdzjsMP+7QwKMc3drkEnGM5jblyds+X1odfE
/cq1lCw6LWgELJS3dO7y2kDN00Wh+NhvH1A5MDMyN9+iPWmh3AsF4z6n4IqI
ssJwnBiFFMm5tPZz6ViBeSHtw5wLewbKVDHFmNB9JmNRK/xeJvIJoD8jU2Sh
LvFE1Zbf7jiYiCczvH5DCEZ9GkbPBMMCVncxmDIxvbC3J+pQawJz7ooVUYBy
N4euqaernMby/P1bJO/8VYYK5l8wdg073pBGL35Ovzx4GQf5RPadouw5cGN4
12k0ztMXeDmUANXKaKNEjSPaBFYl/adx7RuZTne9WwaS1ikc/ayA+Q2Vnuii
up2yNAKrBTcTZJRiOp0acaKcdzWNGRKBfRbDSlCdxj8cYf+gA5w3U2diuIIE
usT4P2VAwaE+j352IDwj+fHzL9qxM67fGSl5XuNrgkRbIsI4Jal9Ma6nMF1W
1YBeRZa22b1avP/SZQBajX5FsUMKV7xdueq2EcbA/eBuEj7QXICbrRU9wpzw
vDSt0v5FN4hAlSWkgoohoUF9ZNiWuKkdMnKNUOCLCCzzD3bujGZfMK52GRQ6
SSkWTeKnRVcukukz0cd+55K2IpGdtTdcjG8A5/Yp9BQ2Ltr6ySQi0Omh0xKr
/Cpv8/Qx8sOH3NNf+1eI40IntpTpsy8xrYE30HtcSAmxyzWhTWibLXJr3xc/
eBrIojSZwMn7j91Et+GOHn17oJJqq2trPScXimQgb4ukkknZw3o5FinalxCQ
08n9ypZjbfuhkQ7ZFvxaakfokqZIJl6rQNXjxOFCn4OtIr8pGezWUFFCDIYH
XYePlMvV4rB78HQs6PdO+CVANghWW5Y51ykf+anbhPjJGjz9FLCkzHshqPlO
jXRigOLXv+lzdmvcgu/a98QN8xJkCY84+S1fmHd64Txd7sbsDfhA6hjt4p5f
QbGlDs0tks0Fqh1cgF83d/igmzNU1O4fjCv/kPHNlKe/Mq1R1Bj6ff8XrssQ
jl2Wvdp1UozBhSJwnqTj8ouDmNY0Dv0bmqx0+D+AKvnf2lMNpaVeaGfHLSLB
9BV3jJHiHvdBOKNl46WvgadfMM6AKGt8MNwzhLMYdLCgYhA9Vrs2+NxbLsHm
uFSedsmALWA4XRbflbXmdEq6wAPfGhkyx7I8ihMKF9Bbff196YK3z3dK4VSz
QCME+9IRtXxtXgr2iFJTI3uS9h950DpjJt/Eke36CncqBUxKE2omR7V4ZFTA
TAG9g2lNqGjmZnKA6IuKdmQpMrbVTr9oiRJqqYX8TglEvmGPzqlrWdGC03Qx
qbVaQwLLNsTgkwP64Nqmvd32i/xAaYEGbJZLCX5N9rTsB9tpOnH7NFc0MLHC
0aT9lb4P3aL9dmnXwAFmqhnsvAUCdqJw0uRSlBc+rVvPdospwoz03yY+MvFy
xNeql2hxlcToiEiAv5RVtpmeez0sVwaN3wTpebxdrHtOS3yTIMTCMgTXHWBn
L2/AFDukyBYun+xsNPNUDLMg7MDT0YkeWLBFmbTg1jaK8KcwPYNoaTmK7Kjg
zVp/saJf3AdDk7ywT7ti+SAbn7GkAe2sj9r7HhdxQLV23paMoPwIGGHAdzDw
UppIigPhj7M6SZBOfDiGOBWOhbOwCmObhFlAbEZlsdqyLEixclIe8E7KsVvC
GD//BYrx1ue5kLXPkvOHB6yBQaoebquLrmD2v8bzHxvQxwMw4puFUEqZTOw2
sa/zl7wIRnSRzP8X40+OMnyoRAu1fOjD/lTG2gi2atneLbgsZ+JfMNWZVukM
4pwAHWilMD8izc34jbM0GrCzEXZJjpGGyNyRosvtG+WTB6v9E5a9zA1z5qNn
/IT0WaulKQ7x3oRdRYeCAOmyUADqeryuUKPFrkOd/8jPfuu4zWl+IduAKJuz
bb0d56an5NYcmYPqx0RA72uBulNETvf83xnuvSG0LXdieeEAGJHQLR/WFIRy
6IWdeFKBc0QGyZxoDSgt0Oa1k+VEwg44dMdL4SVKmzIiZ0Pzryb2H73eLtGD
Veyy+TP35P1Srb53Iqs70uwHjC/Uj6OwFETo4RDOuG8+aM4VgEQqGUWKQ3Gb
XCR+U+Aw1mMcinYG1xHMgUxnH+lqBx+OaMxX4iYRiDLStmBG1xJPdwei5qbd
aUAs+n3ZfuU2XwmkI42Sl4tXcaeIxmivIG4W/Cm7FS8VQLIxR6nQNRNcoA30
xvaxoCdO3sGI/pZXDrdSlmqZgH8Y6BS6Lj9N6VfwD4gH8KEx8ScJ87LcIUmz
D5Qa5Vbv+Gy2vVolb91ACl+trJ5KBAZEuS6Nwkb2OrpZH8BDZVCA9rq+tBY1
3pAwrDWDQiB/kHEii4xUyCc0Dn6sf/33mKmHvB/SjP1SneKjycEzLkWzbrH5
e3sNCdfgYWK9F++I9z8AOCQQCe5Myffvk7Mt6nNuiGeU+/dh3HcUsGOpdkcZ
5accjz5te8L8kjfSvJlAbjK/S44WfHTA+O38lL6DC+aLG8EMZ0fjOvWb8z1n
EAcKMmLEy6yqLLeDctnSuCm6Xc656644fgYyts/TcOTXzTt3BRPz4N42h0rd
lgWgHmKWdjQiyDFbQVUNTcxk+qeTMLCeUpjGGSV9hp9L+k+iQQnNYj8W3GM2
yUraNS++9GXol1pdODCD9vK65mR9LV2pcDFJjy/VQ5tRLGMoEC0jpaLK49IG
7JUZhB3oPSEFqlQ4kYf61fdIbUViC+W3XEKd7FBg8gUcXmvytndKmp1RKoDa
QE6zXLNEXahe0m6DFrMWPCwRSEQHJloizYbGOyKDwKjpJkuV/i4bDOm73B7e
S2X0LjjfzsoTNsxE5cqaVKhrP22+Padwy47VWjC3gZ33pXrZg9cZ82c9nbh0
4xvLcp++Wiz83A/wmThi/wcMoyqjJJ+Gz9eB6cZbiN4xquNx8f/r5dd2a+cM
Cie7zoB7gXVGULr3h5SNRjtD72eKa8caiaMfeYTBpxNUVe0GWffXHUMmk81p
rNGw9mjXJOmaZHunFr46GrQmMa917JrSuBcLLjyXmgOlePyN2dVVTqzwx6uN
aNP77Jwu7ciNTPvDr2RhWsfNGlUXhzH/wWFK2F/YalYj+YMM7SRuYd+3Sfc5
ZwS8p2RD7F123lVIN81HJhwFqPsqINJiwKCj+cpMzt4VxT8Xi29/OFo4k6d5
Cib+oG0PArB3LnepeYbdFLES7aPi0pQXbT+Djab5ibdMPTGz1/vtP5kV3fEJ
/VtFSbfiS2mPYHTLJaTll84AHbBxs/fnvq4UOA55eBftK7nILLcE4zmK7/fM
AkfMYMIeSabbxOO8OOGe0tsLG8EXd1zMPSdq0i8VBowsJtbBG5C8RoaT8aFH
fM4nSY5NWW3gUL5VoTldrIZqGDAXUEHW3/0qd6K43Y1wPi5FRkDVgutQEdd6
L94MlYYhj3NIN7esA7VCC7oE2HGDHZeRz3clwIGa/K5QfGPpyxGwH/U+7aE9
ebEeEhUJgobzAW+zodgWmZqt4YmVtGNvOECZDixER7yxTEjSIVZJhYCWGEIt
sh+yoQiP4/ZHU1+wJITNAvn43tFENJBLEEkApMKrw2Aqlyy7fHIghZYtLIpS
4yngImF5SuAoztnU2mZWox43RI7UvYsg2ynY82qE01QmaIhHCZtpX7bB33xv
zHSPYXCxdXZKAnQz1/F6hxz+fqRwcSyRNxIaXLCOIiQhMLvSKTkY3XxEYCWC
fS84h26mgFhNSWzSea55oj7EGuzH940/47l69gGpy6MfLEHPeRzdyUY/GJWH
Mx3sQC6RmrXebMFq4gJ1Wrksx4MHZvWZjFehVkhxcrm61O4dO31CUHkrj3R6
u8e4mcXcvY1Ynqlo478kAMH3ZBS3SIwJ9WbVp4IMiZRzRxyFEBYXdNcuw9jW
FqIe2ok+9duAuuTcuUhfMAzmKi2zquHphYuhjkAudAY9FbO3Oj6iiciA0jDp
AvHgS22Dk1Aq2WBTKP2zkmPE0K+zqZZ+ZlSsfbos3bu3WFLeXdXIy4tghNX8
LXsq74I5fjT3ppBpcK3q3pu0bpSvtM2Abt8ZhfSDsTn5lcV7ykC22z9MIpiK
5+zlxu23edt/mGw+FcD6tjwO9Q+bTdujG0G3kzuF83g3eDDRdZQx2fpVQkBI
6x+JbT+XcK7reNA99+2tJz2H7rCVKrjSYcAabTewitTLU3GNJQOmqdq3TBxP
AqlctPX2yJUtQJqqTb562qkZUIwI3BQwfxYTXySUbbiCT8/2WQSju+FjMPf2
0HqQ+Vx3rp+I2LuQNxIemCkOBbk1u6qanOigV1SBaxPxaNX35QQVF6dyUz4y
kF7k8HVvzVkU4/d0Dddg/FBQOmA4VEF3Oimw7H7D7TUEnL2RIcSbicolWR5s
10rjkjyDmlW89HtJDEs2zHcy0fIrX47sIoInWPls1UIYTqF/iFMQeYmAVzNY
Hx9AP7rWbZNuAlHvyoKdNDhlBfLXqe+2sKhnMyNlWjqzK/G7MP7go9oeLbHZ
AvStx8ai+VsJCmbj9BKCbYpCblcGEGqbwt6Q0jN6j4DvNScZjDO6h+6pwlrS
ijqk/m68HxobRcDyJZNe4pL63BC9BBY6tg/kezt1FN4KSmocYXICrWLwBMWN
C39kJHESR+CWfgKs9qpp8dxNJ+x8TlrhJU0NqIg3FuCja3tidWLjeW04H7cj
wPOXrFTK1iVqEpAe1kIVlc5TM11XZwZBsdm66KETK4AP1c9l2Lf42Eae5JgA
sDuPgLqNNDjxqbct5aIoS+ED5RZ6n3sBTByzcMrRtmn0LPLVX6ybOMHOC9cw
JzarkEtMYnnMR6e69iAKRuikqYxKpQAiRwIqxhrMhlyxE48G6qXaAq/Vhbhk
O+qthjt+0f+vltlJcQSaHpluLciEmexvnqJ2iHbm5Ik5kL33Squzl5rtFXlI
k1mlRLgT0fo5ySS2PoH8TWfZ5w3H60DIYYH/iz/nVvqU17/eq3Wf8qHRzKxv
6KGTwD4gew9DKzsgZnGGsZ4ELKjJSWfNieM6bVO9ITbeeIn/sjAfe4HW9+2Q
y86K8l8cXz2sFzF2FeHfX31bGWa1pyCZVm1l2Ts3zOGuj1ItQgl6knQ2FQNP
4LcgBml5ax9GUEE1H3A6jKxPuOxiAFmsAscoh65fsSL032gZhbkVcAyc1cIR
xig1g5cP2kvAgbLvkXZdihFp/Xbfok12OSs2GSg9Xi2n4zY5WxTF3yRR/MAl
IrtHqd3PgAgm7Qn9TEyjS13qZOJPPf1pNvabLd2DSTWyGh2r2SAfZiBwVHLD
37wcVTawtMYWcDaMi3i1STMoy60J/YegRCJlUXaNQ+rQ+hRrAbbOOnG1qm4J
DZKoEtV3oCFcnvMzu4WUKRgy6DsP/AOwcc9nE5+Aqlh2ignUGExCoKbuFfcx
U4XeDr0IpWuY/4biwgJ/JLfWpTxmX9N4zbaI87knO5VufwKM05TX/gB/gYkq
mpVjbtSgQANDox37JmwEG4g3Zo40aFgMDvzcOp4O2rCiSp1UW0djo90y8Uzf
G1ZiNP47nHNR1wOYgF5veYa2fnTGemKy4Gwdbs7jaO4pTAXJ5vc8QkOuw5oo
AajjAEy7lkPJ02pK5wK8ebDpxEVGnUTvMhyH/qxO2hqlzEYPW8suxIBC9yJ1
3JcMGVUoLX+XzURtqyV9CW55gjp4/8r/SIwCCBvMNCixcnYprrghrPcvEwDV
hy6vi3wkQJRTyo0smon63AEMELzoETgTBx18Z6iynqy4oKUSU5SRIhRsiNrG
JedVfE0Sy2dAalrekJcYuHvRTejJXL9aHoNCcQ43fNF+EBN194E3pMZ4vJa3
7jGmbruZGsvuuS4kdZKKHVSz9BPjlHfGqEsguwEQbOvAeYIFQOLnbwk4nba7
afEp+zKYhXj5djSWu2iuQBkyt/fOEQf61B5YMxBRznFn02JPgzAMSpQSuxL+
RGC+sEt7Lb68A1YpQimQj553Tum9OtLoZcxFCEJsKuK9JYsO+wLUTfqWIK3+
hRriD+tfrcmk/tjzh9n7/acc9bqnVYEcRi/RniPVb3yYxdaMs5/7Px1GzKwg
8uStKdquqNjzg0tJgsv5qZyuXIVbQWFjSJVYy3CX0EswUKyiyLZ5O65y8oOe
X0aVkQlWPn91mHJvXpzhEGNPMn6UexDGXLP3Ug3Fk5z9rTkvQd86LiSHtqiP
OFADR8X/wzOzDp8Ts1eOjqRUMEEj9lduD3zp83puY3Gi516ubAGV3766hIPE
nu+iDtKgRqxM2lM8jlTRGhcD39eSdp/8THgaTMaP3NS3gHNC2iHwQYUa1fVi
lcs5Vnzk/W8EXSK3oSj/lBUdsoBEa+9uX1ezIcSQHJegvq0tZMGHvbSwi5qL
TXSfV6GUo+wMWc9uMqDBc2RKr+CVeVYRN7n/km/ECNCn6zyjjK1BjyzLFF1Q
PsJHvXCwLtZaXQsKOGAh8pW3HPXy7uHoIc5SFu8Gk+GwGx35oP5lxNMVrV7c
m7FQ3O7GATREc0AwJ576JUoDIE44mnMIpji/iBeQOMazOTSU8Q2z80oG/7bn
XwVebCvQj3RaXE1tc4IwxJn1hU7uSHUCvoep+BmvPlnHHyB1rjEBdbgHRLyN
8i6269FvmpoXComIuJ8LWzk4dZ/cGmtNoA5/oC8cyyqpm7n0z3gAPHvwF4Ju
kU7i82q4j0kFx5CO6R1e4d9BV1pGc3JAws9dZIJfJhW0eJDEB/FJpZBIBMEK
9t9j3JXSPgV3KDjxLI7h+rLipCkcRpM4Zwsw/uWREm4I4VSoncmDjvKkXlXs
kipPPjTFv2gb960Y/H3UHhvqjo2Mz1aO1jP5ynkFiwos+uzTrsRqCazr6Nru
H/vcA8oEWdfxcVhgWXz6s7XQwrI+Xf6wwX0yPFo8j/6fYHovIZyZMumZOoJs
PdZznJxtVTHuqntRIE8dW3KtDgDvgY7aZYgnGdyaMyrnkxk6jZ/prf4tmTzT
aX6A2Qi+lEwmOIDvHACpvR/Whv5IhRhOpOsagGxR9a/qu0RViGxqgXzgl8vA
3Xjc36EsxSNc6YZLJJ91WAAMxPqIjpLqjz0WoL33TzxMPVK5wCZvBlvU2+bL
v/bLgJUeUTjW3a6Xvdv85RAJKnKdYFlWjX2TRG3jFv92l2WKl2rR81sxPeA9
014lH+oP+JA80Xsy3pUm/ZBBNVZ4v1Dox0/FffqCxsvb1MB9hv+9yFn1oKRA
H5vd/wwRoeXSbXY2Fj3RnUFSWWb9j43Lf4NLzseOUQkgjZFcNB6NLqJ3HSp9
dtT6ZmvuFNvENH2AlAkcHfsMLkkgOgEij8MBwA4hyeMlSwBU8/p5tU6ZKKI5
EFKSM7N/2AnlGHl+J5+6EgSU9icuLZ4wjq3ubA0UzpB5O8dQBNyB8/4VydUg
1a+023331pDDQHEGZB7xKH7odG9NEZS1QoJJ+guA6nF15tBaM1TK4KCGLSom
6q6nc4NiemDMjCgIm79ZYTvgGMfGTYyYxt0LZ2LPAzdQ3AH5hbJXPpJYxTik
N5roADQOTS2eRGdts2ZimJAAaXsbq6v+Gk5ajLnu4CjcBirM2cXb9b+G5RkI
dwJKTKSKMBH5kRflmU9Qb2fCK0APhQsz2dFGCKAx5LVQndjl3ZR98sWPo0HI
ARY8ZGN3PrYXGoG+HPfy5ZLZKdYXRG0he88Q3XzS98k9ST9V0qY9UByUVBsR
aQQtS1NNzkUmLSeTM7CuczmYDEXxNeLfXSvs7pkeqYm7MRzUNd03VdU/JUmC
wF7ys7nc892eBRDtUHYBHUsHBho257HOCUwJ2LF8jrMTqB6JJP5J7zKQ+Er/
5GonR3HiB1ZPORlA3U1sDl1JsKYZ3jvoGpO7el7v1EiMVHl+5gRMKhCadXMm
fEcbHi5EfwyZLZ3c1QAuw9d3ITyN6QscfpR+m3X8ypetmvhTOb1t/Iw/ChOo
bIIIOrWcB1RrN5SPo+tojiVfVoEwnuAayLjZFGeRot6907mkUn0C68IdTz3W
8mDYVqQsFrXkRoYGrRgYrTqFUkIPlSbgePp2DjiGBHYtsjKVBnmo1u4tZe0C
5fx+xbqD7zl3c18tWxBTKH+lz+ir0S/sX6my3u/HgVi/iOResv4+aKbA3aFe
86qF76CCXhbiSvcRqRB1hm6tcFQn4VKzcZ2loCjgP2scZqpiAVpnvdmIibnc
6wHBRryabuvl81bLJl/pPiOes8pjNxNi8Bg73DIu0DYuApTflCyFyB5ZDZFw
qTrCJ3BfroOY/hwJ5h9j360kABaMPF5nSGgxwMCHeia3k2TLDw8T8iXc8h2x
qI5mQKHQhtpFSf0tUiSpciKlW+Zs5nl0AUNI0/gATfD+VDiQdwEgH6UrFCAO
Jn7KdPnKKBgsEvwm10F9LEksMX1ns0OmMoIVpbreIvE6DlOUEBA9NoxedCxN
1fDZbcglRb+6sV8j62gse8AW/bSOZ8hgADOku5Dw/GjEtfS7BG6bJIuZjCqU
qpUxvDl+A70upxmATF9lWGcFzrTU3A8Fh7Av1x5+Rm6RgKrVxS8iUoAywbOD
P770h47oKV/Afw9EffkvFFwELK864WPkfQ6Q4DxmGYFTEOtZ062/6bKlyCXc
B8Y8eGRcYnJcRyB6fHYgDB3+0QMMmDrjhGJENOf6FVpUBd1VrkJAOZ6nc6UP
ngd0YSauEnrfP/Y5WzPzX/IuDJRke8GnB56oA1cWiFze4mdje1vuLShy1/I+
Qu7y7MeBKAM/eDr2iFcZIWdYXvtEyi+KxrsBa96UMyFiX+vmfkas4Zs2vE6N
inoas6M8ulHe300Jogakw7INXi8XbmwHvTd4m7k9++SH5zxFTnqEUlbSDDyn
UU7wq9WAP77swE41HFq0kH6/fJZmgtNzDBkPe5DyY9hOfFwhWSBS6mlKsQtk
7Ed1grn5tldha+nZjRhKh768hqs9G/WX0HBfvf6b1JjoACz3Vv+A6WC7Il28
AcKyO0p7eH3nUvInvteromedNWbq+75AUAzW1H3n9/me58ZohFsKQmZBT5Nj
8gXI5kM077c7EpURMm82bJSRkA4+IneXoe5ck6RxXRlyl3anKxR3gZOwU52n
C7G4V0J2UOy13MT+FaxFmShDd56tYbngBCFjszCiaNmKgRgETRf+WE4a4O3M
8TLWvJYKHIw4SMo1JS80NlZvJs6D3e26vPPF7DrE58dgo8c7D4EgMBguBCKq
o76D796cztry4VKtA3pmSPSl5v+vTIr78BDwxPTUKhlRfvRNNuCLxWXN/eyC
OqQ2F7gUdDLbG7YBjCbU48SqHf578x+vmK+RefrRPzVJetU7625NQtQwdDyH
A9QpoYxL7QfRGiE7QiKCy+X04br7aoUwQmNmBXDIxRJRiErqHOzh+LeloyuL
PZ5OW20cd4dXAz3gKalIafBU1hvDGxFfyvYH0YJeiRL/Dm9tDQ1fB9RWB0B1
RdMYXTV7KjmmGlJph6pR8zVt6/usgnBgbPXtfDJHUehtT3DiVNBZhZxv54eg
b9twb34EE4C0nNfiz+gnYdjfcKAwt7Hi1KhF8fD0OjDXaPxxGUNh0GOD/KIS
DAL/j/wdTpHpVwiEvln1RkWAQLsIBdUlsqqPQ24EW4e85s7K1ZLcAPH481i7
a4sx0rbm4u54JFifFIpcht4+nst59wLd5i9wxvc4U6Nn/WG4ds/QsMtVu5jL
U2DL/EfAv2kvxBft8HA80/gqu0b1gS7nbezarCx/T6Cwb1bYwg7/VQMKpdkt
DXTpS4K9r2Jtg+YkSx2sbhKKoJ40c5MT6RlLAU7gvBvJbAIkSSMiYQdsYkO1
kInlizOZUk1ANU64EOd9OZ7UbE1fESswANxVGvkHYTSg9XTn38jvAMswRuer
TZhhrt0rT0lLxVpTgUa1xi5pP44voHkVXidoOrQDugKF21PRBl6KjNx6b1ai
FXFB4zv5j3xJ5EQYAEiZ87iwy5Kk50vISGLOgxU3faRSDbiOEmwOIcnNOiji
zYEERxD75jJX5jmrHoJ0qzdXgL4RR5j5qzmjjqcEQ9nnUHrCLht0o9rARcmM
6fWf/+FsaYsUGb1hLLV2BIvMu4bnGtCFZUHXfgSfSTRvA9KtTz964YbqNRWX
DrxbBAEBh5IZ4qlGmY04YYF9W2XIykVCEKk0w1giapCor5EfYKDOHAOisxHw
g6Gyi9ffC8qg++FHyzql0JLzvuiSkPzOzOXzeuoV1GtmpCuKsOSG0drrSpfk
CBdA9DXPIZ+QO3BRtrvTbYpJi6a346s8JWSVND+u6l/seLfHPoy0nnYLsgpF
BSV5hSjAAtLeoaCZfyB6sy4Q2cXb83TUKstJacu03b/f/Td3aR1vYNPPwj3O
tXWOjOVP5PUwrfdaGst3V9Fp61nWvSTfVhtA6VfstjcdNpc/EMvgGMyogc7j
IfSFJGer2vdUqiy8hFVDyB0FuzjSfXc65fvy3KIBiu+O8PXEqf00SgiPo/as
xbOHu5vuvzxwm0hCeqfL69B0P0v4EXVOE1y41YO4qdRs/tI/rOcG/SL/uvCW
vv5oAOXSh2FlE3aJHU4Y8iIDyuxZlY+AQmbwsoEbELEamgZGRYn7A8cu1QKF
ATNFUrwbMnt268bJbokGa/EsTlfco+VopfgMelYeD1tL8QWfk2VkVQcw3GPv
lWrIjS40u4eVVyfPtFDD9GmB7iujlHrlN0KTW1+u10qzURQEPaknjfdN5sCM
bVfIDqVfDQp27kzX1TDZm9pRG0izGZeVq8uOnxvlNU48wY2yZQs9erybbz9L
vYXZ9utyYpzUapvTmVPhTikpyy1WQrRoI6K1kwDl3cwNsvbvrDD8GDTk8GrE
/FYtWxcAob8mevPNoQ6DxlCfDQR+k9Xltpf00X4OQe22uAtVf/WNN7P5k+xs
vug/ikFIw2vPTphk8bWtImKC1xfE969XAF+FQo2o2VNhOmu7xAVKJEtJaz1U
FuDPo8FZpYwwlyJQzWsvUn+wf5ayjxwlPlQUOk+sVQDY6LDn2gerdwa1HKHF
/myFRrLvgvcA46USF41V+lhe95Hd2z7aJvgtpG1vIgt8/0awyPmu1pgbUDhj
J8PLOG0LQbpIjML3e0nJlxPoKtoCoXnG16MJVOTQ2Eqp4OfzQVBoiuOfySfA
L7cg/2WV0n3avmGOxlh66+sRSxdmM9cF+nJ43haaspLJOsdYOS2hqj1BDowN
Eokjg/K+pOzk0SPHZnHbHloAxoR1IGRa+TZl7o+oBQ7H+3ABw1l2J8BOj6Q1
oEI2jK3ftsP2jNYEYF28gn5A5fnrxkzY/rxD8BVo9FYQ9lschFqCG+5Pnd4j
tOHSgnp8QHhFiaeoRzx7uqCkKxBoUVNRbtrv9cOGb5knRsaViVLgqW45ixIk
vX1ivz3dens7Hdk+XGyJ6DxzSeO7rbxQynXDildpDZP+zmwMgkDj7ZIY4DdB
yBIUMnrdDRE90Hl2hLt60y9VmnQ6wJGx7xwSh9keLxfA1ZANXpkDUu1oScHe
Ije7U2lLiE1PKu8I6sGBjiwd6catAyRboiD2PKJPlQ==

`pragma protect end_protected
