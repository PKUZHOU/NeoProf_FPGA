`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
D4cNTH2vkcXT08p8qcKOy1fA7kZ/ApteWU2W3UyNRqjAFDVzijypLQuabvAs7THv
YyHAR+m85Vaxl1e/UDR6P2cwMqO8fPlWnTRLZfZ2huhcgPUx5zDMtD6JUF2VMc/O
bO/9PnVM5UWHeG2g/WXT+kNJ6awR8Oh28ABWhQU+NYQ=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 13088), data_block
dWIr79KYdV2K1YMVYXxjzATkPzqluzMNWc7edGY64bz+zyU0c+HZ1fwzv0qqtv4+
4W4JJdQ0pq6EnDJs+LqlfarYnB/IBjnPlfc8c/9HhIz43F67+/WUDDa+dJ7VIn1b
iSKKmlksiQK45k0+uGO5H8lGTGMh/Xb8yhF63wMeOCPnhdyCDXJrBqnRU2b47Tz/
slXf5KLsOLHB3s5wv0qWrAgjg+XunKgdOk6ENrMxLrp77IkoEPtXunC2w9yHPgLv
BMJy+EneY/LKkTHXmQwtbM9QifC0xSfNN8Dls2H8PSOzg85hUDiUlt7KyXWhKFTI
8up2xCHUUkxRm/NmToGMJ6iYnCQUhv4d0TIwOwXd36kfzsajVEg/FjuFyFcX1PSW
VrT8oC71KKpmTiH0yXNJJuRlXh1LULTUA+It3f/qMHUgK/49LhZ7tY2b9GLzL0PU
MzKqBn5jCDgwGOVTngarCFe/8RQVbjLdr7J9faihAg9fqDN2Hwm1Rw7RpqvDbU+u
VfOqGqcgQlK5itoz5Ofy3GLceIAALqCc5AohQk7saWW9WpwmrFbBrPGLJFobKZZK
mswsOUi5sE0rAJk/MgqFZIg/hUpujMhlxI+g0RWj/WBcT7+hXXsfPRptyPB2xxX3
nq8jvrAyag7SHsonvbIZvzBUbc3mKsnqg27WAQ12zGvsM5gbTbuLVJL7vYxRZRb7
0iuCfhzVE/59pLDXZqNAgVg6fYHIUkNtetb6q4jtKOfk7d6GptR68JhVflyPD19c
meGHDvbLyjLpnHdL9/U4ncLhrDGd8EE7wa2pAtRkYugkOVUXaWVFtLU1KOutSQHS
4lwXq4lWX1QkOg8cgglwalEf7QtEUVY4pBHtjaRJvNH0bf6++e4LFMVZIfFJ/Xz7
itob4Gr7VF+Sq5hzNEozJhMjmQRej2tMKjAq6DrDrHMvoEqpoJbzsPMJ/b701m9a
F36B/hlZ+c2ONdv1jioszDhCt4vkfxK5+qHKbGSJNQzY9zeIPkPvzmpSsib4MBne
7/RaJg1T0YKk5PV7CV6TcUUGZitVi15pwtNellT0rFrrQuxTzjiiSqrvUfay2eUc
NekyQJj2Cb1SbWf5C3+zTcKz3epo5M4ceA0qhHHzIBS9bciUZHyYUoK0XE4oeX0u
UAccpOVq0fJTqsEE/eDOYAb6UP3F+S0JoxFmT2aqrkIYv0Mowu0hBWLwYtf1h59V
YV2Oz8VZR31QvTt2hJGJgilt0y1hygMBXSaZctzQyEpTfPWmZ87l9uLImjOBLVZi
WX76BV2DVWln8mGczbC5Mv6461ppqEMbNF8JxrRyhHtt41TYV8iI5QD/xX1aayjI
TU15NC+hPo3yrG4v6MSrCl5xXRUNLgRTM+Mqzx927pesjKNBXcmkU5M/Oz2/425N
Iav0iSJCSocQNRBlEzvWSHyP1POyumTjxw0Og6njlm4uby4arqa8ixPEfeoQmBHE
LdUft2n4gtN6IvjtbWE9mBiY08UJi5WU+Mc/A+ckbDZjnUz3KsTgxx43P+6//fXJ
nmQHHvEP8ruAVTHmBROS+WR/w/V/bMo1jscpZ0nYo2j6iTMnILajKEvQhG3inbyn
vDlkB5HE6JoYuW7O6hd73Kz7zXme25ppz80XSUqrSTLVvwwWs9ZqhGHw0BvXlVZ2
O+5+VN21xm7k1q8CUSmMwrGv+INsrwF7zR3aOOp4SISoHmVfm/YgXY7OMNDsH45s
C6VgnfcFcMIhVRlgeT0bmcgNP0zAD3QntUpNpUPFqflg/QtY2+U8xPvmbcD1tS7m
b8nKSkjevKYgQZe0ukeIEqMQvyn9ZFTG0nHqLy+AQjpiz1DcfVUdNJIJNiRfSd6K
K7BqTsnFWUyirjFXEP5lea4PbnugadnQbl5oDegztjJTTTqvStPmzjZvYXT9w9UZ
MTGL+0H4PFBCir4MsCLzZmMXYakULN09WMAqb8SBfuo+qr0bDUaIxyiG1USavwJR
VN+PwtoJCiynv/9uroRFVYJB85CDrzbx1mAnUrx6hQfrkBcfP/ekM7o6S5/YpK9t
KkuDcDAw8w7lABPYb7MGyaqG6lc5/Yv1F92/8vjzg7K3NjYnwS5nASI5LKmdNh4L
9WeHlIh/is7WZ1LYSOIuvkzcmSO2nzhZDGJy4bTntsfZsztTO37nKIOcw52LYaW0
bu83I9bA++EWoo5F28zni8UhLvLPpRSr/r5qBJmhtw4w9PaJdEyJWzTU00TXZB26
2Yn0Sf8IE9en9nPICEv6q3I1Fhv9BjlLGyCghGJE9uuujm2afBv26Gyr2K+QHAdq
UsLWVsI7MSUkzC2uUuvU/YDwfFcowqVDWl/3+VHX6puoqdW8RSkPjH89FjeRV5mR
YBRPUt8FiXhdTkAE+d9UHFVnjRePGCi+IbQPBL1Am/0mJs1lsZSGr4le1uC9FVGz
ONfOlS+nNNK+cz3YHi0A3ukYiqhVxdZfUjmSp61VgJdfJJRHz8fbc/8gdkfVDa4r
4Xgg5BZ/LmFSvyVM7LCiKI6kP/YMBaMVNFc8W9RTmIO37j7LWZ5l24fM8LGYyh2u
7G4i86NDSxobo0+FBEXsMgFbHiBvqDEXO08cb6ZzaTF7AB6wtr7mNxIECx+h9O+x
L8XdONtcf60hYg0GqOhIkHLaoWmxUI1wJrncPLEZLjqXaiGHH1SLcK/htG+9Kzgn
IHeREiAIgDrSLj4W0jEXt5x/F2RmbtyZEkWP1P+lLvRL64fUxxXRLSj/bX0HLAJg
RWSNI0tbUYLIWSE6MGQdvffLwbD4883WYQieMaw3xHGDkwYKd5+guNtThpodXzLR
m03NCvMbKr4lJj54JMFEI9wGZ31wo6aKTWdLsVf5pajg6clPIMZCvuuBhJlb4pyd
zgkoIiU4iaNi2Wj9Orr1qGp8sSXwnk32j3OvOErm+tHDmyJ98KDZmpwPOg7HX/R5
xhsFKkVfvhfYe642H8O5JVN9uRZ87eLNXdyYk2IoEIdo1rwrqrV+LRMwGTa0bdlv
NWNARHA1ozj8jtgtTOumXfAm4LgbMvz6SwqGI8g17CcJYR64EcteAIzYjdsbvux6
nXOea5fHK5yOIy7nuqe60hlEnl+o0Oncm7GH88Vr/Yudu4OF7pU4BAm/X/w/vF8+
OiPCKfjegZsJpbmlslYnIQuqGPwH/J5+6VFVz8dTjdh4D+aquPbuLlJzJDp7tPHy
VQ/ZemwN6Y/Ffr06DAhg0rJF6/ZNZJHTlO7SqspZi68sJnpwW89OEhu9JwmaQ/oa
xdf5V53wOQa4pdxiQqC3Z+VzWvqJIY8vcXGymPH8Re534OZ06e7w652Gr8HOwXtH
49L+KkVJYpA40Ctx9u2LUZ8x2/xrBlGRg5wcR9czwWdJAKF7xVeR/4/d/8V4dCO0
WCYPSfaMBw+CmNuN0fPhO9AIwpOICN613TI9FDckEGEq15Tz+tKL0Vy4uK2s2x0s
6bKBwQAbXNt3NDrSLt8ZXzGx8AsJJLS9T+JUHIi7jydSfH3jHUrhdDj9r3OKcIc5
YLS7qSfwmX2Z176VMro1hi8Ia84uSKWftkB86n5zP05VTkzr1GoA2SR9gvG8MLwx
DY2YvZBwERcIcvovNYiZ2qEq0pbzmVlxLt91dZU6i4xSpt6mBNQY3l9YN97FLnRY
IIh76VQZi2ezgJPmepZkoiefgS7MTP/HChrN06CUvIfuMIXDrNovHYpMtRvHbD2l
SJo6hEM7JnmQzZ3K7N67KiHWmNJKBQtWD14cV6RzE7Golas90fwGzIbRBoXaNyfW
vmU58NFGYPCLgXbU0FnaTewrYL+mm1fO8Bsxw+O120iXee6qbsYth6EEs5iWeZXc
RSALZ3xVvaLilhUsXIX0axbFIpQ3IwNItOWZ+YQWr/FnLAaRZscCMsbqirkJGp7S
zJWGIadqHQX+9jeIFRJcT8X8jPUf+OfZbvq+JJEP89kr9vQRhmTbxc/9Xte0BPJB
O3H4BEHlSH0TJMWcvmDfS865l8/ctSLa7Ekc0OebUfNIrNwS/HIKsMYl9TKUy+pb
+Qe7Q8G04ZwEOPyCfQMDO91cRtK2DmYl+X5BY0sqpHBBKCqdd87Z9VNJmg/YHu5r
vQ1kJZsxfmrWU12kx2rG1+0hLh9wVl1zj6T9FsMukHgYXup1PlMKbOIuQPp05yUW
fWMGeAg9CIja3ha2aeZ+Akmv93IWsoUCxwe8FZ2KYhVpj55F/EhSvLpkkROjquyM
RHhUqDaWGB8vLUr6KLQwFWxQRfzjTY5WaNSuHTLUOv2kwQqgpL2ujveARy6bw7AF
X4SF/XxDK0h0NCjtw5Pv21ygTIENd36JVco8GyOu0qcQfBQxlNCSMxKOMMpPHO9c
By5b1Nn7WgSVeTS91H2LP3O+pUE8qt7wugXNSE8smO58QDIPhTJkaYopXkFg5WV1
rckuVIBz8C6rjPP/wO3676husziuUNF8piSjPG7yBhnTRO0gDSHXeMLpcFjGOMhs
9V16P/8UXvJCv2VxjrgHAPcGWRftQFVMw0fegDLxlze5QHKGD5w5mH1aGvBxpVv0
PoN97fQ9Kc++JkjF5t/j/qQMP77dQBuot4PlC9MyVewyOncxyJim2+XnHjWG0r+O
HbpC9pXxIWdTA8ROA/ydYyHOO+i9SkX6LgFcRuwYbiQunQQe+/HwXdcD8OpGwsSi
o5TvqRTSKevhuKpArucjF1NTyOejBlrZ5fs8PoUBfil65/B2yd+9pGQlUOUAc2Xt
4PBzpGiXVCvoUNx8l0Bt6HwObz6iCwS85tOY54gmzgB0B+6wj/LfcQCSNSwUNtf2
pO3mjSji5JmF6MoI3ZDEwyaMz8875S0jq3QZmTHVazlTYzushUHypGsLDxmI7asK
NuVW7zsdvFSrwyrSJE6RDfpfpOrXLWj0oLSP6z334Lf6uQRT5Eylcsi1ZYNOHuIW
YFd5Iql9iF6w3E1l0WVnOL9ir4WoV3fF80+GJieCcTWbrFXOCfPRyvmgIbG4L2Nd
I4T9H3Bg5X18JExmqlhr6WanafB6BxXFHqCObbADtPlbpilgI/RhZluF9qI4ytUO
OL7ByNzp7tLs5R0HkHFEYYLYjOsdhX44DHKzF30rwvVT3vdInzde9KA2KDJzVQBr
31VhNf4cJBmfbjLhQw/i+ito8Llhw6f8Sv48sutWMaSkVk+JLnjvEX8Nmxkhw5vV
p6jSZBHbASk+JjzXA6M0UvdWn0MSlxNINSdkD1esZ0VQqZbOTMVI+hym+Wc+QYHL
2gT0kjUR+Q6aRVV0ERw+ZF+mzpT4lZGzUrNWSHksxsl5E8xsz8PRnWh3jUpzFz0F
gpk6sEPK/uD15gvuqO5UmnG7ODinYhOrz3g76cCf8eeWQX71kKDksJtWppRkwEkg
bbfDjW3pPVJ6UJpXrkRb0AV9wx4H306jJhfh26qzPOQ84KMYi73CldMvMQeL8bM1
R+ywWk20326igRnIcOQ461sg/1Lbgr0Iv1Nf1rZlEo4f7oqZlUQbwAiQz/h+qGzL
jgjcpmiLqcsJ95TWDFknaSUtWGDntGxIO825VDSzJKhTf/ayxA/EldZA98QtzEn0
NNPJRQZsuBN2OGGvC5Fv2dwp6LKCsvG83MIN+Y5gLAMKPhVSvDplHRW5tl+zoD8W
eGjiQjps2o+K/XmJLzoUFVtkIUCZHGHY7cwVCPIGyFKxx8UxjgOjPey9NP7am3y2
/1B+mwwOMoLdbCmww95hxpKj8u25n1+ced0G6LUCefQhKn4IZ/csH3YuxT9nyEqN
0O5QdWT4U4mE+neArwZbBm23nuqLivQ31WlGSLe6MpLvnrt3h8p3hTkyC3C+Sbf6
BE11TDUqv1CqMYgpxMkAXWu2FNX2Q8uz/L7lcg+jJfnLTJLgOuVJqxA00V38Tbfa
YLiy8rGUlUG3o1jjcPv5/VpFnjUaiW6LnsR/IDKRfmiXYfDgGW4urgA2JJ7Ow+uR
NUnMWWEXk7M4kKIaIxsUJ/XMQwWRpQA8WTvRUBoH7nfg0+ZAyBSmXcEK59nkeE2D
ziczJLnpG5vAJZmg+91l1JTzAtBVrzQp//I4pZEIGFegAOHbheR8TTpZDLZgowYD
uvZoIBQm+iSsWzfJf/0W+SeRE0nYIwpWMQLLMdz5l9h5d5qsVFDOEh0HyLKIVhju
YVSJr3cENUd8J4vmZUgRMSC6tXXCtclw2cPmMia+AISIPkhAXXh/8XiTp1jzYeX9
KU8zAf46yRiyWbVZGVu58upupnUtBq498tiNXXF2i7+P9k5RHHlXvPA+smngJ2nQ
bH1GZUs7r6AfI6pPP9k8LX+lqNFsYPrY/V5OZh6ic2RfZ/9hY4bRSdpHoewgCqAO
c5VjpaFDNzVvk70N3FxlKxttsg2FTI1yLCZH7U6SFqu6qu9zmQvcx7QXcwMkpqTo
9o9XglFoDSP3qLG86+FkT0q5fmdsd6iaD+FIp0WA/XrYveC/b4e8fD0ZQEb30W/d
I0mFVyg7dm286YHC8LjlaprT+03eChRlMUlUr9OZkvFc1+u1KKER1GSKfJuWo2Td
Ke/HawvcwP1WAR8bTQmnYT8XDl1L9hYGHJByXVpnkEpSYyAmwQ9Jc/7dvOazftz7
KYM90FlCgzblKMl2ks0ifFV/BR89RfCN51rp7GEJeHzp5itz0TfClgotl84nI5YZ
w2+EbkMHz3Wx96Y4ZcmocAvVlrvvapmvgODag3XVGUJ4xHCyd2V1XpzZeypDyVpc
kGp+HuvVq3fKcgAhQ2xptAZ/8BkLVstocfzQDsVojIJRVq4OVnwaqzyG2Fxz51du
gbOBp6hlMh3f/TIXs1AKSCCnkzAgUJJMsbEpedjOJFCfD98JzHEl3gS820f5KRzK
hyolFIiwEpmZ4yeuM+U6zq89hQC8xL90L0vvPvjHs5g5JjLLQcpu2kyrdmYkU3Gq
vhv83dbiWi4GEQT5Uxpo23HPGqJ5MsPDSyPilkkZc0ZGAsuKQTKKcTnD0pHrmhdU
VgYoVjUmkejY1q2q4/IIaF3Dtae8ejgHnq5zvRqF4FnoGYefths0weqsW31SBLw+
MwIyjJdfnMUbSzIYORoT7D37RXj8dCZzifkwObUpw6NR+R+bB5aUC3b7ix9UBPEV
6eCiIGszIhRaj4bl5ZKB72LCrsOHBnuJJHKCgbESwv0PjQjOjqsHGqJv9PQfjpI3
RMNxaHWVllOkd7xh7Kw/9yQHmkrHXtjnHK+vVtGrNc60G5p+XRL0nsFQ36F9gSiY
BkdrsQ4Q+PznLd/vfiD3Kuz2nEFiqX2JDo5NPKzbMaKCTVMWoJybQ1wB1dRkPghH
6sLHJ2wtzpGU3CgGhPI3l00orS/h1xL6qNh6ZQQ/Abv3iRrgzCNZiYkvt4eZpQWQ
dZ7x4ktqjHsGT5QLs7ohcDaewyg4Ty7d8tmv4bq0w8VwZfCNco2v0SJk6VITVT/I
+QHyLNGsb3HN2flxgvsPFqUM6rzdl9jtVMK/370dhSiIVp4Eo8qvAJ2oWHKL8IBE
iZco5tdvLj2RRUa44LHEyZfJ7IqGMVCKJC4VCc4XdBIwKWfz6cu9LHrbVreTJtVk
6CWjTKPtIqYEO17n7cY2TVJXVpc6OgKmUn1xltar98lNNQXxIDr/CEnVmxYiRXil
cOnGK/s0d0gPLC7DjdkkjMwqSqvsL06ZwOnwYGiOisGFfw0VEzCbFm+8x1YuONtT
nh9ivuND0UUnHNBRB3GA1I2rcPnlLXYAoxc38N3W3SHL1fVtCU/g6/erZ/+/1QP6
auLZljqUXk7JY0WmIBElt9Ds55X2Ke8ZfFcxRXDCz9HhdJTg3DcrXMka1w+FP5kl
eS/yx1sTW+VzP0tXsXLvpGQObPj1q6USzt5jZuIrgrIUHccjXrcUMKBtC/qXpuAR
4y30zecptKE8T3ACrnDcWPzgpMVLJa81y/VD5KU0FRE4HjWreXFE3Vfb9ygtMkgP
+kCPNlSWQjmliEIrPdTYbJIJjipWNWGY/SIzc2aareGzrWI7hH4mQCG3XKqj9ePC
tw4DqGERoCyrAy1yU4kfZi/C1vU/S3xU4kq9lWa0zoRJ0LG/MLwPR3qJ75o4pWvk
02n3Lx4tOX7LEXIGvAxuOioZVxi92bMW94I2kVKzjjf3QHV04OiJcEAI4JgynGHg
iVKDv5eDrEKqQ+F+RFEwBceszZg9WcMgSZ7EahY957hmaU6br6OZxA9vUP6hlQSa
P9stCwuw8BKqquKyfw2Xiyb3fF97HnHxbs5O3gLP3fn4vJnvVDl9ZA++wA3fe2ss
Q3xgEIWwnfXNOHBr2Cdp9MEmwht+BsPVMuJKlGE5zRvyC8vZI5Pa/MVBOPWCvL82
RxKFDhS7ZVifJxWuGzdR2nk0/IjP5+WVqzLp0KfDKff6173SLAGBch06J8/LQiG+
lLpJFRwrx/dI2n58KjZLFK4XSdW2LtXKvmcTTfB6ketIKF7rexm3ro791gNkPNLX
V1lyZDYW9Ei8uF5WvmHPyndVYhOhe4yiiLw4ZFF1ueqcov1JbTF1m0+YfSHy+5df
oeIce0UM5RA/YP95lKcgl33v3tv9e6o/bBxPRAX64tqwYT7XkpFIlzKtlg/6KzLO
/yixOyEDOFDzI1XRKIAsA2v30V8PSZPSizuyMJ3qro877x6YLch38K+h3Z5Rzt0I
FweBeiaIvk/SDdD0lPv82lY4c7FPG/a8heTh23FP1T5Dmax3cfT+1jocsw0Y9/hB
aaYEqkiMKcE+306k1q6L0F8IsLt71yp5DJHhVutnRIldgHp8u44GN7epXuEWUQjJ
Ig59ge1QKz0IpE1psYEhVR9BLUS/5gJeAoVUOdrPRouMdkLUn3eJ6Pv7eD2L78Cz
lUMKlj0SRhcTB2Xrpd2qMs1tcea95RuafoMipM2pF7XOqiB0V0Xn3X/Q3hdnIEg2
hiJk2qb2Z/Y5+rNdXMbkqkmH4GIPIblyprmAU4ceYdX1wqHyJog56mIpaA6awriG
qJExC9V+IXIm5bCr+itPA2CtS7zuY51mmmDe2no4g6g9jyaGZcxigo2hvD7REAKp
zf5j3H/2F8yyNq4ocK6CqHXQwIAtXFDdsKoaZYZR1z2vYbQIyL29b/0MHCbm3pO2
tLDPWa/TBT0QtQXIIbj/uK89lLdH3Y2MQza/W9J8HTLtYd2PA+UXsweASki/lROK
AtJGPk2Frt7RvJFisheih3DCwdKl3moC8iUR2liLq/bFABgOspo4BHuIoMkblOpu
hymIcTtwqBjmFDPGGcJAicont11qiwRfMEvTBaTT2bdSjyixly1I+pSIAYd/iNLQ
66hhvDrX2l5QMnclYXhMvOqiaGdE8J/bclgc/uCaNhOwGmFG9S/1ouei+SWi5N7r
NUqT1Grw0lWZkXgOTv7N6FlYdst0oaWo7wQG5AuGgm1RG0sLrx4FzzZaQtzMa0Hl
Z8Nt/4GCJ3BC4kT8bYRV4TPFbcsnMfl/YzbkbPIl4J+sGAuHwIurov3Wqq1K1TLO
3sw/ghhttsqYn6/oRs3wxs4H8CwGIvtymTpU8UsE+pEgEoKaotF1ZTB7eGk6m5eQ
Jj5RAbOtaerw1mxL+0FxBQa9wziWztBNOr/yDcQkyUkKU7/7aT3dZGSZr89LYhwh
ZHWMpFjrxU/0lg4Se2hZB4A3+67U3DxPF8ciThpoIN9mZ7Un1I3sNwIdszsJyA8i
jTTmm5Pj3fV0LRpxujTUL5LJWozn1m7Owc9inwGjIcdTIXKtylE7SrPc2Rl14U25
d/Nn4XgRFIl3rTNaJD1V5qXi5Iv7TzDlk5HSxrQdIpyZeZcEM6dfpZBKv0BrsnLM
EeqftRpVN/Wibf+vpn1hggp2ZxkqUOnYAKQ2Mx8RTEIO2xTQgA8JVFRho1w9q8aB
LYZfbBJ/XfFa5NIYlas4aZ76UjbBG2AC0JFA6Cmxe/abxybqTNrBCVrt6b8lyeRT
gAOVWXe/FYxs0GD9e7d/UQDLqY75jwUUwlADV9DhltOe0C93NqeVkHD0t5x2bszO
4qKGZFWjF/caFLNxIn2wbTARB2KakTmQIZR8TD2xVWGuKqcHnOzDa45yOY0FcLwE
B27d6kWdkNJnoHiuR8UVpiIt8AyBHXWvSuKkUc2+vnyw1tiHKGS4RVHbjQDS9DPb
Q5BEfMzBOXYvqebY9BM4qcobwaptXtk8Bj/rX5kSvhjEI1/jR5kFLTXAPEPUwFjt
CX3H4y2rCq/Ze5wiBAyJqijhRbubDH7DucaHanwXEWHJhsGqzkXnz2lLqzG1VB8+
4tr0wGGq1dRu4cx1CnNUAfyN5CAVo8+3aslOSV726tJPSbEBo2SKqFtl2fS5P93I
P2Z2OUgSRvLCvogTPrglEgGyMIMPczZsX3Emouv4Xqj4uQAfpI4fSvvBEZBQAMTS
a2ChdnaJQOzgshZxtoIzJChzNrFLPW6QqOaA6rFe3DNh4XJXHcWKDD4DLAsAqtWP
zm3GIKon2RzbzBR5nrFAtFEdbq1fSSO/EaofnNNV47qR40ykg7aAeODUv7AeJBeW
SedbrZSukCQJIiqw7wrKgEwyvXafd6IPxQ45q/LDrdcal8ZOrXVgNfsqcH7gIOUr
CriljC9jmuCztyfcHEKKIty9XSbkoGP3K1baZkIXujqSYVjEby3+vn9po8AiY9EQ
xN/L4x58fjzYbMqvdocptiaS5A9BN2HVlG5ze3zlWGlB6aOh4IYF5hxL4b1RHFyi
dR+sSWOEDBnKoiynQrAEL7ksUuIike52hXriqsuMEKtEdqc9kkY4PWPZk8m/Sf81
TSYEEwXxvRWsuzY+aQwB+iwFh/107mq8ZihorMsVffJ5Xc3oDaM8AG1kZI1sYLWB
h2mrIwaB7fGzYMOrjz0s5pXn+CeojiP7S02ihegX90jn1aB6r/E0g0l6JOPHDnES
vxYBx2DmtgkQb4ak2ubUt5bBEh6RXmbHpKoZC9qjFjIthtetbQOqWbZBToscamWa
70iFwvlSUP2kD2HsRhmI88rLivkQ+2HSrr27JsuALMQiwA/W3DjyaYUBjMyicJqo
xt/jngs3w4Ee+gShE//bZa8BiB1Kk0RrB2z/4cNewMPhwqmTOhxP+ZlREEE1uF0K
/3h/BLS/0uSTUPIfGpiikMWKlIBc1l7V0uPgMETjnEfRtKY926edDRWjt+uS+3hy
dtyzI2DRB2IlZGwr3cDka/BFU/R4kO2lZTM6qybeCN9waBrZiK85QtSxcCbxy2Gf
gMJ0rUL4beFFaCMf/VbMu1WTSNYvd65tnSqfNauysBpt1uDQm1DGcgGC72SyxcfQ
kG1GrmSZMobvWtX/6sFeFr301SZHrEbPb+PMXVGzjiyRaaLyfD0vY28HxRHdpgU5
e4jKn4QglZjURnRJxrC9Sr4YL6mmnwKbTazBFdc3lGfS112J0KZysDJEEYFC3/XL
aQhY1UdbSO+PVlpGKvslIjOmw8Yj4tzCQxIiPUrtSGoiliSi+8c/NQc7ws7n0DFg
ovNyFi4u6g8sbGPxlEWtE11hOuiOT+f06c0ivPI/Tn0FLMLLbf1gs8neH+tULjvH
3amipZ8S/nRqm9XCM40vLhPAg0c0A54elHaPAyDCMa/VmRGc9N9WZjYxwPPpgXxw
VS6W7aUnVNtGM5pslqPtLGSwfIJncyZfbFjVnCa+kSOAqA3sccg5B/sOi+yghRKC
ejztXtgryjvDZcEgZ87S/AwKBb8iBgXUOqg1LiHtxSEZDrV3yjo+PUB58uk2TgFi
UDKM4662LFMX8BTJdUejUKQ8pQdVGnZqQ+rrrUl7ceCIgsKN/O1IvePQ9iyhEKHP
TbKp60zvrySqS0j7VuWQ7NHYhXIzW6G3wlhDN99Jkt8fscWdQZDHF4qgIGyI9eWx
klrwCkLYsRC1LhkW215BxmriJzUm1lXXsvKD0cgYSfamzwFpUjnXT8AGl/+TJtsr
F0U1OeDg1pymcNYjqUSFHS+W7SL0xgrNEhPUgiZ/6fZGmBsofrMibj99T4nI0by8
ZefmXzaoDWYe0r4CdHBaqS2T/p7ZsCZjjqRD+BSzq1zVdeA1z3ZSQWed4mJJi8or
K7e/OslAknoJRTcwP0q91hFjq/o2o/nu4EEeBYb+jlGau2uwfhKjWeW5B0ubgmQU
fHqhGRnFrf+VuuIRu98NXhOmr/KXSU/cJsF/H0ffgWvvL1SaP2RtlSK0tXVAQD6d
GRrPLM/g0wXYaZD6MJGLEszs//y1NCs5gNDs0/OlSkTumo8e9OEHg004414fnAzW
6Wd/TlcfCJ72NMzSFd3t2yoEia2Oifz697awvachpYVYI9z1XldQnmTEZdUhjnEK
EQ4qpZGjfMF/D0pCadrQqwotIY7iyq8DMzJp6gfv4Cww1YhSwpuUjGvW5tmCXWwI
9sj57V3fUFlQNs4Dbzkx1ni/uAv6tUg3fcvwSnefcVQO4XU5RB21AiH3DlIEc9Tg
qVPNNTFA6QSj/lJyqmnBatPCztKtFXJXwhSh3fLJrdg3wUndX1f39sEPusNWOzS2
L8ufNEx3CmBtOabQudx7pOZEA53TQaFCNS5HLdGMVjpDfvZr340Q89Sy0m1VURZA
Q8Jbnv5jv2oRrBcTgy//rPANCpyg38xv+BkWpPd6Qwq/nznSCGwMmpVKeOE+4PxN
OggjPwyMYKsCW2GGh5IMRNpOc1c1cP1jTH90T3L9gYvTebOnSu9qCKMf5eb27JTJ
L4nptQQYVecWkfwey15c7TCTSVds9Klls/GDvS8uYQeH5MDQUpg8Tal9qDtY+bQ8
fGcNvmhLDQlJMlP74ndFMxan4q9//JTwEtT8iZKTJc4Wd2twMcX2zatTZhMXU/xl
LQhrbTWAByjhW1SLdhHk9kZrbomE2yIHh8JSSGbgiWZB2fgmhm/VPpPJpBK2DHaz
mdDyVirK9FoVnclAsZRRPdnxt2zQ9sFPuc+mpkiMvixMFdQwJmtuY6tzqK9HTrR2
UMjzDxVm2+ezox7d8nH29XfMpthdJcxSAF9Pc8hM2eau63+JNTjZhTjpEA7zTEwp
ewfgAaKRNz270Qfhz3vDcE9OVVTA1pCuLs9Ap3GWFGc1ohz+DJLJTqtY6a3eoTRt
ekU+abLMYTAOs7ju8DQdlvdYH7J3+lM49z8fbvTsNBo2UuCZosa7ShGzC2SRbbdz
9tc5cFKTvgG36eHADlPNnNf6mc0K/qX+lvZOxbem8j0mORcpYMFG5cYPrz9GL5so
SAOWqKS9NXDr05QrDO7saA+/sXCVPqKoHKWXh93F5MQWxhUWNKjnfwGRxKuUhwUn
7MHjToqS+IxHhaJUokrxFfjKo07BZQQTL3wFFUadSgqzxLVPmTBq3GWoGFZxmG0Y
KwxgmhLWv+jVKEZ/FqFPfJ4cTh2ro4Pd7E8D/8/UxHjkP0BhSEgQ1LPF+Njm1qiP
lYBv7Sa7OjBr137PTjq0gLrIQ9X3A0WYsAP/jGPgm6U5nKtwNB01CKIYsoTlrRka
zv4iu20+FfLBooiZFr6vEVmnpcyWC5VnMchKs0LhKWKmuhqgVBSU6V4Cb5xmAcdv
QiYMAeokWi8SPUee0lKxDYxb3SyqxY8dulAtAwcE6GTJsYjvj0j8UD2JBZoYQ1SN
7NvnMlUGAnGB5sl/Vn9CbhMqKS4YjTTDUfyWLVPhbWs9e6qTrqWWSnmmhcbVfc2h
5FPhvXMioaEr47oDDEVd0S1Bc+QaWhGYNSRPW0yC1XAuGaCLIYpAZyVFlFYtdl5L
6ah+mVBezTMZS1Ez6on1V+ZGhjtpTEaBrTK0Gnl4T4rjEc9eToDOoBT3MlX6xKLg
mDDkYbT0Am6a5n4zmIJ0FjBOjXUw/bBrq3fcgtEdYYv++t1AkrMQi/s5SF+ObGmF
g1J466bz72MRQdqtax1ZOdwi3NYNVqNMPzlXcVtN3W3UQZD2Z7X76oSRCcdd/M4q
EYUkYZZnfJ+VYfBWZ0oB74lXooRt5Enny5j+KiOL6Uo+Muu4s+lZnU5CCP//iIqM
LpLL08RGgu860LNbirYPnPh66jpi2JgtUkGvBsIr8ygkCH6s0d6pEd9P3ZJOnp1J
5n1pB0q03mtVwZkm95NCf/LxJbGan7jI+5m6HuKecmYq+3u8ytr7fG/4gpAizJyx
2vdsKmuhk3dHzcAnvnl+HRJyFQ2ejTPjmJI1ufX39Y9TQT11KXwDHWvwWVNEtoeP
lWJ0G8nDWLXIPtG4Gf54luulkImn7E+U0TfNdRHfO78ZVf4ajPjHMvYk2F79ZmUt
13/sBUSrEDjnTjY8+og2Nfj0tpZtjsOJKvy2nXtzW/IUzQ3qGccA01eP7lCbWA/s
heitnUpMef7tt4f9nmPHHV403l4n8nH7PaJkYd2pZ+oWTDQZ9/rSOgxIXMj15SQy
S2OhMb/Qg89Hoier/KdtaTIGPCty4AJA4iw3cH7RUvyLf9v3SNHDeaJhReZC8b5+
ySACMyz71HNL/MBiHmbERh7WU/lx/MCibSnwjIm2Q51umHGyajYkeO/T7nsVxv2p
4O6wuOIc7u9tOXATJcmX6+B8GH7RVXH6a18J3QvJllcB45/NC7LtgzcS74SZUfsW
dPmh+muaU6UJCadrkAL8Jq6tiDNz8UkNg3X7x0RKZKEF0oh7Bgx09Hc2X60X+1GB
oAmofpKM3/rUpAt7YTfUadT5T/vCzBjpdNuK9gNHx9uQfQ/fkgCokZVtM4+7dIGK
Wl5qVubBVq2lvUB3/jKlyHISzM1mX8ztMUFqoAHR75jA6nECV22J6BFabKk23S6d
yqM+BL4723Hne/d59fG4csEhu4zTeJpa7ueQ5x66nh1y/sMD2vtrLZzXP/HfS57K
0dMo+xyWUfnSC/J3yms4+/FfgK02cBtWYZHcwPZsmgPiEzF5s4U9xBfsl/bfW7FP
JlYuy/i4Bb7KQImgKH4IRMhgIivRVo55pbeMpYr2xSqNzozqyDKutVy746m2B3/q
MEPVkcs6mkFyHBbobT/4i0sZWzVdxxtu0AxnHLCxam1uz2T3ccatPcrFUBW/jGLV
uT+U4eiYbsg6Eh/oKvbg0Xqk89O7UHP3GGM8ihN1+fIrdv5yJDPSXvTwPdUT8QSb
Nr4vFjb8FbkPqR5/AOL9fA8ArDZax14dPAdHW4tdgYGx4doRTH9AgXkpcScwYSTH
OAjSqmtC+FykaEXWKPVWaiCTW7iHxuSlDRSO9M2ea6OwompgMzpX9pU40A+xFTyE
oLmnsUKjnpF+0DNJk/5Gi37KJowSSicLypK2KCRb5OA8OS0yleksHmKRMZb8k2Oz
80YTbHRXl3kcJMlf60Ll2mv9bOAddsUUaTswTljSb0hJH3HM4QYWqVcD3qDo5Uym
ip6QrqZRmaKLdcCJF/h5uH7LzzoACXDihcyd/b5Y4eSgcSmpz25oeaUgxEP6F/4n
GOuLFnyah4NOuQoE0fryy+DtPi5I2mZSjpSUAHOjVzAa3MQtt+/PdAWyXSH8it6G
K6EXrSRiqiOJRT3Nl/klrnOUs6rBZcriWJ/rcsKa3YRWVKgnCZ4nkgfmpyq3u5ra
7VUOAHbahEu992HN11avVUc1+NcrxU3BZ153fnWI0+EGh6YsMMtijxpyZWi7GnuE
8kWaqsG+pTPUwv2QBCV3BZ6pX9e3kBtv+VZDtzB/RAWqlDdX5bGgrY4Y2zU6Arcu
M06I3iisTNl/v4W9R/XTLSVk+t7ueez2EGkW25HNlcTo0NMNH3WDB0PyGo/ERegA
0efzLqpHDy3a5kYkeic+U+diWG9+bsAOkT0Ee712w2Rig6oFyrl3aNZqb9Vwdw8k
2POd59uXr4p58/rur9HMFE7sbfp3dJ1QqWhyTwY74q/iUV1k4apK+glG+jR9bTb8
MpfRwKnC3apHH6/GjGzvQl6odb0fHGiY+5ybG0iM0K9QXvz3IyAJpCC51JRlBU9P
T0qsftPsANogDT5Kc+wHOUJpCLJ9jWHnssLBUVbR9H8M53f2fjwJg5FApfEWY/W8
B2rj6s+O+bdXPedSwdCGEKDPt+Qzh43ZQ6x5WBzmZnczoyMWXCAZ4mgvbaenThWT
onP5HAOgvzDo62U0i/JCZ5dkyqLwV500mUrkuOedUYyBUbBaRGUMBn0q/scNY/KX
5OS/FNw5AVA0+L34mlR7OfXla86ZO2NoS5F2sO73QhJQzqhpQvXQBTFjbm0DcjvI
kMC07wkSsAVQlN9tc4bvqi5jhFK50H94VgCU5bwn6XBYSUjUyBkXeD4eUJxnVoO4
KOE3azrWDcmJhdBXy5BeY+eCmVvIlCeheW1XExP4RkCSghsAElnLq0+1rj/qbAuy
+5pULSCgZmKCbx8FSmd2L4G3HXHC3XtjUJhgrEkKHf9vDx8TwrZ6EYMjyuPguJ2c
kRr3unEPDhGsQwzixm3XzWE6NEzM3XTsaB4BbX9SDnmzvzFIg3OmxaOi58xQgE9k
dL+a3tv98gw7m0Y+L6N/DNZ9rgrc8zJ2m7puw+ci6MO1v1aWg5pBzYyEYyXZm/5P
A0eoZ7XvSb93z+NLmGXNvV5cQw0uA2rBJfm8T6PJ+mUl7Eary6K8tW4jVUFLZlge
227Ufhsw6BUQ+VJ8Uxt4kPkfxQm8Rz+utXu/YAGCcQTR3QzEAeWABhplxSVKntfq
5e/zWdPHd7I7Y6x4V2ZlEp8ynSOGdXY/VeZ5NMxkU8tNfHHVTBdJ57QaAqvcu9Rf
EeDtYsjq+dwp0/ewlsnzgMgJBslM5xgF6KRu8PqNRuXnkdVwzNaA/S3Whl5ekUhQ
zfe3lO+TMtatDUdCIg6PdM76/ivE8Wab9KdDWsgg+P/3imHHlHjN0euRpO9D0xDs
+coXL99V54+wGppxwkssb3bAURQx3qI/NTlHyNW4HxoagM3U2RZktWXgcEmWHmgo
9S36GTDBHIbLcFwCE7rklsxSyq4NrBIRfeepGPjvjJrsXhh5lgrZyV52/DABAVy7
XdCi0dGYr+tcQ+Qbmrmwld2Z+CfmwNGHXNZAls7VG3BIA2OQlsiIR9EZWrjCFuul
9I7yCJq1ik0/7fmUODrFvIrhTsC5Z3RbqU/tpCV65uQVFePTH0/YgQjKJIePor/H
CAX1QQp+Ht3Tq95hVeL+bTglQj3Z1QD+2AVqqoHqZbFwYuKqSKxV8DRQ93b4jFQn
YjbYKuBjhixyj1yJwLUUPw281CsTlpAVA8vQVzHDlL2HBqTqQQC3c9o92ieEaTrd
aaf0eQfXKuR85jSWnRh7SYC3GIN4BGIic+EXrC9qCWeuAfgS+nyn3VlLiVr1a+hJ
3S3ZVLbIQhdoarjKeJssm09FMxev1U30XvTmAqDupYVXaaAvyffZSjFzmJFZUM5o
/Vvqntf1ADi4PxuOQl+Y8uCUXKTU8BcyUrkQYXJzNjez/u2qTc+vt5w4Ge32fUAu
SB+KJted1qPlFgXXIHr0rTH/8vYBdaZ9eWyWqSA9d6XDawfkD7mZ8NJszyWZpiiU
MHVvjcZ7wAMwUS9VCK++MwetgvOO+Uydn8OlLle+dlM=
`pragma protect end_protected
