`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
P/BXVLGcQ1fv+YrpM4tJp9Y+opty2t6oA7+ceBPzr38edEBf9AdwkhnAQFG+Qyw3
vI7FP599JYwvIErKPWMUrrgoUIIeNr0g2cbUVKd5EC7tIM1LnZG6UTd++x5zoSII
DK2+kGjcXR6Tvs3b0tkhfA0HtwS4oqhoACuv+RXikL8=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 26576), data_block
46RNXSKlTCe8ksqu+pEUQvsr/YfXICKbtQIC5dUZykcG9/w02qniDss/ZQWMmuJ0
cnRwlS9QMB8f0wkL6nO+Fa5+4WAfu0hEmQYaoDmPfuOQCGawlrd8cA26f+0UtGrN
/pulEHgoEo9/C0H7gSCMxoJlda3GFvpoKMc/lQ0B31wvGCxx9w4iIo6lG0lBkYT/
vBGYnqvMK2VASOOrY5Q9RiA0gbZpL0XZu2+Zm8Q2GtbxyNyhKeSv6XdOtTOfbzzn
xnl0ZAJQuUHHTaPEdM2XYIyxIgkLduYNtO6yrfKWVgRn2C6YHRU+pHSZV2w5ZIDT
2I4wsm5WgYFrL/Ebm4Vbb4TQBRwAYdRV/XXeTtsTRKFVhr0n3jsV3MRxSd2TeRT8
O6ZTpJAbSeubXnPx73n7xB6LEF6jsHSWx5nG+Qe6mUnarWIxZpXyxulXP+Nhw3Gv
lLeMR/syn6b8HN6l81IKPq7gKVAWejU4mKw3iS8n3Tvy0BX8me5PCg8qJAnRGiQT
kBd53zPig3jTBpNOYqrARmB2x+Re+F2LVq5aP3kyp5GFc6QSc9LrBuBMvFFWXqa9
8xYFuXjvl8K3X3hyoWrUDLt2eYe47lfgayfjOqz3etFiQWpsDTIf4XLvNzq1i8M7
tJiGI2HhG8TzOlW0zwUnYAFUvyANBd71laqgT0VFDitrtLlVvq8jeGmSWc8eKJrl
wen4funQOxOiyn5ouJlBlFL+S4V2LKrDbhqgFDMbu2a55Roy4P/TpythcB/72lId
AgleIkm3vFaLHjSYjyy4Le85t6U3wG+Kh/PjVM7dMpd0Lk3peEaiRC2AM8LEFvAu
hIY0/MC4JaBhtxKgaQ2guAO/VU5xNzui+SS1p9kT3fR4viNkPpfziGgZSit4kfIP
ha1FBNaVPXsF55oZoQoxw6OXymZDNUAt6yojaPPVOI6Wdx+42on0R3V3aAvPtOql
2Ikx1+g8RM1t1QZmyux9vIxl6SNl/21X/XMdoOWaZAhl06G2WZQu7WJggwAe5GcF
4kvKbKTmkcq+bV1Wj0Xi1lq8BE8yPgD8RQT4t0KGhAzX3lqQzKiwBaOF46fvkhLB
6+y9RryEDuwedgs3Akte2I1lLP2OzYaLr+hdrY+FCiDR66nU2/f6d1fZKPJZ3Eud
PiZ2YSm8WNa12mc00VVTM7m2IuVEqm9S5TDA+bJ5vyq8k7Jft3CdFZZWgEmfGFcs
+mfAJfBk1o5/AaYXmmFYVWEONs1vNkD1zMpKZ8nxtEa0tr0yi1ckr9OYtNlciQx/
KPsHF3N+nprrlcAOdZwmwdnGNMWKIougN8OGuXV5be3JQzn6x7zc7YlUVnPq3wHg
y0d/EkMzCWV/Svx6XLW99h100MGdaDSeIj2YKmEJp59+OQIKZsw8I2O3BvXvrpS/
E+RILvXkRjHAjvvdfY2X1eP1as4dU7EuQjMIN3FaxRDR8+MfTygBfV+iCKKV8Aws
hLS95EEMSYEs5Z2Xf54m6SYC7wNzORQFqXzwDOnPGhPNdTlyTI3UA1y9V52QzNkg
CEbjEcxe7cUBPeDooKEgcy9NuAbF038K8KeaU62+T+GSnYsa4e4bzkD9R1Prn55t
r3TU9tZKpanzZW7C/w6stEM3xIqsrAVCaT33YE/UFFckeqDUeVGwA2IAm1VpGPhg
FBluueG2/VyuuvkrYZctw9isv2zZqT7K8w/gjs8jrR5G/wnvtuHPPIq2KK36YRMn
BQqn98O4syXEfszYWuNg2b/0dz1U2l6mYejI5Z/3Y8SLrGDZtpP8bZtIdOe3tYBo
9Sp7ZT8Y2O9uCGvqVlD8O+F5Pgf8o9mqnqtPGgjReCNoJvLqoxgp56yPU6YI8ppb
RzFmcw147Ws4odI86aHl8EB/IRAvsVyEddEw5xXTC6X+VSB1z7u1CFMcRC9G0BnF
WP93RRw1+Ovt5jiEbKP5gb3oJLL8Q90rm2y/wiTRoOWY1ip1sZS5WlkfzQJwcjQP
PkYrUlChbbL2tlnfhfeqgkgWItWz5CCk2biPfmmEY/o/e03xXN2/vpBEC9EDtymE
WdHTLuishk8pQNwrWgPMDRTCiIngONbb65qoZ5figpArZ9aPT9rjdRAzBCAU/Nex
twk0i64Ph51ntbyrlJqF+ZBXjp+SAFFBeln6SD32reCN1JprrqEJILarmjVqLV3Q
IGyIS0kbOk/jg7FYDwyb6cuH+xHn3S/9MNrkv3mPBCSLp3zKJ8IPf1wSGWokKnrx
JZAJc2Ay0q3DH+Kg+wwwSUef9VljMl35oDR2LgcSW2PyToArVMBd/fe6Yp6Tpg5m
GvgIntH+u8Tbo1NsDYtEigR8AnW1Ac0EOJCrIZ/C9oFlGgNB8OF03YR1ycIuvcsX
311R1+592PfefiKUntxTK43Z12XO+8mvbO/FYFOWFWr4/SnNeufiN/6TyJzYLRG6
C3dGVO/BQHADPNe3t4b5n+kMvr3jO7ujWplbMzznNaWDycnuzsFDn04we138enrc
mv+3SJ3fdTTm0TSHQXtmh6RFT/DL1GfGCaVHXGSH/uClKAT0LlnQ5nm5/0SKdS3K
2Pazle1BDTMbwjQYx1Vm8ULtK2By/+lEcAiX++FW1+piwgTxjd17Px1xQbpAZDb5
2wgGwfWl1j+0SC2IXbEEg3ee3rSFU8TEMhRXONgEE8RA1zbgStRm69OA6ZMAkN7x
iWYVAR/EOh88GWYImWUURfZkAeNiQ6qqnuRgTHCxkA1TPaOWZkOapLtwyd0O7I5c
sCxAv9Ktv3KxWy9rykFcmQ1R0bUByilp80PERqXaD7q/wixrUOslXf0PxCRKW5ds
LzMkvA1J4kGHxsRIVR+Lje9aXuWY1KwMJgajGj2ekL+9tXQBpHGuZngIZQgHraXe
IG0v+nFQTbNa16yzSP9JBHwyDqzTToQRB/037Yz+/P7drKfWquLlGT0MRpjJQZ/1
D5sQcNREcRHNq/gUj2cGNYC/zeN7rkHUK2Ur5I2bhOGCTlDECEodPUANO4MRGHc9
OZ05xAihdicxCarm0+/ASLwto4+NFF8jSo4dJvAWxGOcgDNRd2z2CD113eD8tiBG
MVgiiv3QtkWnEPOnwGogeIj8sfgTutRgySHIlbaxbTYnlIRRkYklKpDQUECpHsXu
fIONQkF8wWrlKuzL12B8h5Eybsp4JqUYhU3nu9xf9ARAhr2PHVkttI8XgIj1fGsy
XPEC7MDLCeDkafWiNP5YqhmzWKb3wKgD4NLNDhFrX96oGrfyqTwky3ezgUnpTwib
XAdKxl/PSLFAc75uDHRhEhzVrv6MaoKUJ06idJQMUd9kcTgOICiekfzFCtT3YDdi
UmhKFslSXDDwDiljsdiE35awQAsVHlNe8LgY8ZUMSY854kJ5JnzYgqh7fBjItoPi
Ef3tDfYUAAlejxVAeu7uvJahN81EVCde3xLCW7Tai6j3T7WX+stb7kdBKe6t7yzU
AvJzqBuP4/kZ3D2zG71iG7rNhkFqQpaK3TLKYGzpttdiKN15TXuQIu6QV5itoR1H
M4Oqdq1no8mrCp8EoizZc1hXp3bY2gDkHXgMvP4GxSxCI87fpQSqdRt2hKjTcHRI
wa1C9R9d2h+k5xM00I3msZWdKDR4tD9mrTKmFyIQgMQe7zggKLNrDe3Wc6/vzveA
pqQ4o1qtSC/rgZfjc4H7hhmKoOtNHXoMaSzSVeEtJIrm/ZhCOV9lLtG5uj6YbiH1
Dwdm9Au10D9SQPbntjODhlQkzO0qwIk9iqCBcUMUvmgvyLwfXxCkAFPZG7Gucwpz
kl09reik4v59eEKUSGOvBZYBm+5pd9PyGLELN/zRy+BAx2zOJHYA2s3IiSSiyD3I
CkJDp1M04U8kIt3jGP1XZoLEzFfAQ7/JFI53FQu0GkFLXdHDGclsynDyFY0ox5O5
PI5S0vn1Y8iJadqlOYwjDCDCFINLpVXlZ5ObADMPVJHRqsMKREVq68U56g/7x7Me
5HDYqLP8QJL01960nqOWA8ujMk6PyOr70E+KWxrYouaSJ6ZTItAc2SSYw77oh28d
DU9xS/egit8vJKdze0G5zQH4YI3JRL/XPW3g+6xS3/G0TP9mdgmowtq5pr/oip+X
F9Z09PCm3EJktjy8RBRgeJq0M2ff7Eb57IGdxPeonv4B/WNTtBDtjl6nPQVFwb0I
2W2AvFvF570bzsk5v4kEQmnMmHbX4m8SgPEkbcsGSAGv5/PVAoDL2YayA2BjRvTh
IFfokdK+0qDAg0TBuCGegjtuC40qmny1nF26VUs+ikVbWQTBr2B9y9YZETqTF23v
Z33DTwE9n9rZmIwUl1tB698V8L6qzxLJa2W2P3MlQwIQTET8qGhucIw7s31QP4hk
+eQVCDxjM0Jgntg5n5a7yHvRoQzJq4wG6/ZFy5SJ8GtF+SJ1Pjz7iPKQTkovpRSs
z4gXqen5ia0SDPyHnHw7Bgj1Yb/k+7vsxHv5uKMfZKexuLD6MfDqqzGSFUcA5t89
DR+P1LpSPzoC21BMyh4CUtdYhXefq3pib62mXPWuEBNqDmfIcG2xOqd103+77HdK
OuH/8nVtmrHSmLzgTbWsNAkrjDmsLW/4CUrO2cwOHOBoENswV+ioh71QUIPWh3+W
wTcquEXBvdoYMvZrDBfP3OCgDvYMV8dPA2+NPgldUJ/4yp8z6tEiEj8E3N0Zm8GU
xLmA0ZgheI3Zjv7rYgfXZDTz1FQi+qxEyzEBnRS6GQCJjq8M2V0yuaDFuP2ZZLXF
sUpDde/enzP30FjXwNeS25RjR+5W1wJLZzCz1CQlI3sBIYVOMO3PTr197WjmJr9T
dGP1SsIpC8szqCjNZKkfzI9ALCYRNVv0FkFGzTiYv8N197IsXDgiaiIov0TYtk5c
cCMKZG6wbjTk0pQNVjIZ8FhCijPHoVVVlE36Qdi7vSMzLcspufH8ouCYLesbLeQ4
nnpDbXn4wG1D0GVEAaYUXdjpreFjPip4Fcp4ZvyziNnlp0nhCydxvoLrXdI2n7UB
JVSsgDUgY090Er0rXsFeK6L+xDji+RNr7KQg4WaW3FQxnL8I/sTfXLuC9+qFeVQV
zq7Q27tL2cY+KiVKam+LqzPQ0PQQJZ2xWKi735FvbitgRRUtTzrKLdXTxOsYpSDh
b7qP0D1liHcP9nHAzzeescn86rZ88hEQkSxwp9ub91Y0TFmokEl3uLh+GMCxQ/vq
FM3DaR4gCafi0FOc8gIRP/8jxxJLspCexuZRtAHWzPQs+QZuzowvY5y6dgk+x3Oi
OV93H7MUOebzs4Myk4ixacalDAhFXbmnP0W8GJTCebxo/Uu9STIBmlshJxe1orH2
ScQeCihFK9C+sI2j+4j1TdCvnkcKOiC9FOBlKVPcdKrxsKmY2retfCn/tz6vpV5v
3KHiS0G1noyQ4AKUxjae2wyoGs5GaEDMyNFvsbY5cHMVq/WW5a8CI1KDRNPnj0Jb
ajR0V2PW39sX3ZDshhgoEymTwFO96kRmaUzhO/hDTh+2neEa40QPYFafmS3swS/u
8VPqRy7Dm+uAukjUx20mSVh+87obnZEbfCHMZWrNCIm4U91JMjlNlF+LbshcA8a4
9RtGmZXPAdkMyGIFeHpLc9vo7F9xnzv9AtxkogDos9PlCA0FEB5Zqur6BrvcV40i
zAxelioVg6uiJV5hyjdEEZrUCEUAXPrrB6lyXihE8s2itOrH1kWOTiEuaBQ4AckN
ECg4Y5L7FNTb4jAZzIhDeN9DltI9Mg2FC/TJI/7EV5voaZs6nnzocJGGDc1OxugI
mzHNd52tLWnR6LE6np3ybu1y+PeQR9rP2vp1mRtvnG1uQ3pPEANxMqF1rdWGOoVy
BqmS9gEsW/47oLXeoA/fNRkNIVP6JfLqg1fnCoWVdGArJbuABUKO7slTIr0/1oI9
ZwfQnU2YWdQ8Ud8bvpMn5FRm93pF+lZzitlnkWveoOYx+2ysCLgrHEUUEBlhsad2
RIpSg6oiYO45fJcNfgTXR8QLEFwO7cD7M5uEnGN+pPGMcrZPh/3ibVVA+IxrZNKq
jVzElKVST/QRR9WBenRB+gJgmJlJponn77ElP+fzaVP73qaZy2I0reFTlHtonrkz
DkvRwRtmHRDCjwBMJI/Ixir+KfPKAA9Hdv/vVmVwHnyUbbckFSoQCLFs+CjaCUyb
xQPd9VX2q+Gy6s01SMpq0tPaZ3uEHqtMuaVKs+4uWGS0Y8cvsuRySfsevUu4ZwRR
c7rVTy196oKiY4e8VGWrwnmUk/LeH+9uKnGx7DH4fcYlXBH8C0baM/nh9pPfCJL3
ECOe7TpTwq0XeHbJXaBcy5OXTEClxNPBspVR67FXPn2maf0XmlVOsgLnsbw/KRUL
F+UaM00/lwUcdcbcHwQ3Gv2aom9u8AKWm5EnREeRWdT1GcGPPNHKCbr/kEt9QGE+
uEzxRXFF9A39gM/jbQNIGNVc7vX4V+t7rsF6saKWjUSzHH4blA/qMTj0kagj54qe
LGb0lI9aJkRNZ1Dz1rh8DHGOWVzu/4wVRyue/tNMAo6tunkQti7cBESt3mgpdE0M
bVV3OLn7HaeWplkY+p/wVk2jjvb3ajMYc3bCFaspKM5VpHdSyuzkcPpp68dwuKkq
MTi24Kg4Sq92xihnehH1cX5B+nRAJYjW/dq9LeaLOAumEUW5gHVZ6N9TWGHaB4ZZ
lkB8WLVqqWE90XH2NcuopsFVgNV53JlCuErB7PNNIbBplnd0OPAYLUhIsIMDEy//
PIQt3JGLMssDuS2f27ukK6jN4NGdFu8B2l5+Rey0GpGkCmnrHaQfrNtKBsHP5+k8
Y6v5u66vbyZXoPdyGNfWhS8N0cJDDcqkh64hvYYzffF0IRnIXES9pV21KPsdv2W8
xgZMyFkxfyj7FCmfc/NiiusRRfk0SYgCjAzrToYfB5Yc1uhX3adgA9Mxk/G445Na
SmTWZuiZKS97HoZ0HQi9M50aKlf6YwZ9rRwpSVqvPmVwM2yu/p5uD+UpA4ewWy6u
kd1uN6ZEie4g9iozQMzZrTt4l38PQUBuF3zdt2e8wmQZv/KdFajfrd6sivwcHNsq
FJ2sbHhpIei3AkBfCvoUvfItx8t9HQDdEF7mPqrC4E1v9zDM7Z/+0VkvUfLmRKTf
EIOWfVGv4FCILrcr7WpmY9r8JQ95GSqk6deZC9ocsAPKKIdgYomcVhXG7jY//It/
kKlSKBjRiz5FtjEXaaB0ZkmVuancY6buc/NQwDgbhN0XjPtbfMTCfIhf7x8MaAja
jtP2FlMx39SFlmW93edjohhTfo7dgRLXrPrDNPJePVHm5d1qFjoq7hqAi0S558u/
UMICmcAANddBZELgnUBq2u6JhFneUPfdowS4/VGauNDVDlCVWbEseJVfKFv1l9H3
LxE+2p31J5gnELtxGATk3Yzh4d7EKUjarw9dFA4zzDg8qP2pk9cTIVEjCRtjeF3h
xhBDEott0pyywj4N67fAcaX7dHmnc/tm6RX6Z8WFF0Z8HR7dlKjVixJlNIJjcCrW
fNL2azdKa32jbJtPmuYAIUOBxTozEPY7vz1KUKyFxHYrlSY98V88H+oXYAmpUjHE
02RiBYnqX2EcQmfq9qqFZmpp+SAfLu/lG75ePucCDd7BMS9qHlLtiUTpZKh+zdb1
2CrOF6p8wDTyEtqKiPknZ1SyEtWUmgPsVSOVbGEsZzpYCxV9+sr2ZvvRris0w1H0
x12k7Ek1XdYiL9dy6p7WltIGtOG4vYXFXxOBMreBG9R+AO/MjpHllWVpP9ndQXUd
lyvKhfZsZgq6MHBeO8lF4MeeoiPwsVCAEE0QrdO+htsZXjcqif2mMWHyqzsuBT0g
dk7FtSFveLIl4zf2Pp5ovJZCEzegpoTGSrfGTOnVY8p+dfLaLfXPHiL5cQxrXXlt
911xc08V7l3dJRUVOyibaIAHjtv9dzksC6w+/AnJiPC8grrzmJVslyasrsbrg/TK
C9tJS+AtXRjVXyJz/kLDk87l882Dja3BbpG25yPJhoWG+yZmYsbChbSc+ViN+FW0
ocRS124nhg2kxHPWYs45sDy61wo0pjrBDgDFQoPHZ6bMmp+IjQN9Knb3G880W3pH
3fXaRK5jFG1OuS3y+HJTrrOgGiIs3BdUeWmLQMyiUu0Juh1Obtvk7iXWC0guqZqd
HQVVhIDuKvujIxEcQSIdAuFLC9ah5pCeaFd2/DWrzSSRxux3c4oU+1p6VvEBVb0m
Gpp9Vhxu1srIpfPQSugu8exOYLxmsYIj6iULV4AuqD8N8U+N8gItSleZKiLb23Uk
Gb8X47yWmJ+Puo4bx54gSZN8wqOPXPd8xO6DT9I8R6IKIJK+nJTYgWkoGDQFIFEn
qKawkIewoWMIt1/cSlX0EKNGOdZEcjoQVz0Hq9Lb5ZrpW0STHUOmMJVBW40Gmh3Q
TT+6cDZTeWUZlU6STLuCCTqfCJbYDoUfSh/cEvwwhqs1ea+VZdpy9/f5YOWh/gaJ
eMmHFC2g+yg5prZuKgqiHCZ1Ochc6M70bHUvPQnA24E175zQMwyG5vvzd7E/+Zsh
nMNec6yB6MXxmRpoAb/WRXhRmhIqc9UTVpl4uxkAM3APIc5M8AOcPZhg4AOwc6Uv
zTeYeI8HF3QHh4hcXnibySTT22GjP0Cga5x3iBniGCU9+dGy97SfFOFKOkpe/4tk
C64bUrihL96uqNlRdTAT0KcbFY9oE+AZvNfxct/UU9AoKIrndYZ6R/7AMJzA2MdP
UaOj4yKLvhR1QeCToZvktXXGCxg95Zr2lZbA8qt9VsLl+yXhx+QoGXOeXie/FJy0
jkcpmsOryZ0FaGOHj0vxUP6khRNEGwfumKx/4kWUKO8dfFa5zEfO/35/fc1guxpp
1r62jiOmuy9iTlN10NcbPHzTxKdaSy8fx4ZYGoI3xGmtR47eX5o9lc8R6jllLvXq
74/Ip87KAuFmYkkm3/aHrnlgUgbsPRt5u5vs+xYEsehpInxBbaMWcU27Wl4RI4Yh
lCajKjDJMHbvO1tdCnBvevohUW6O/DeP37CWWx4gGrYnkWHOh+H01WtHXyTbC6J8
aQSl8ol8AcRtnt6EUOdw+Xhq0znsG3Jj6vAJ4df3TwoWJaxebscEbd5k30SaUDqU
J0mNcChUkSvcDFGtNmuLn2RIKBbJ4J/9A/d9lANInlNp77lq7cwzYMGseRcnQsnq
10cSXtxopnID4IvXMI9fA4RnY1+OJLMkbB4Z8zwd/7rkn0GpiacBc7FDQ0ocgY+6
Zm69WRr7D+o1Yvy4Uf7F92062BuW96CvzXJm45ib7ypcGKrWetG4cDq0my9RhUxY
2sGOZCL8+quueJf6n3J1bkbJeVY6FTHCJWPfJMn1g8wiEL0/TiAW6Yvu+UhU7VjL
y0jnVFz4RNV54yL5W9RLlMo8NENV8BzTs9Cbt0jK3un90TekOboaO+O2PMphprW8
m3L6gE3ZZQNxb6oMwHeXO6z4tyKtPYVfQu99qD3Q1JzzvbFkV/lcXwX5pEOh9pNm
UeYRh84nScm6zGU+HfSo+xjo+sgsShYAlJIcqB1muqK527jBWROdGGqhMauaUu1P
zH2R28BdIEBg0R6eBoqjIsbOS5GAEXVRCeodICGSSC/2bogrlfK6DaPKiz/k+sdl
9jUXg/fqJUNBp8qVeTzD2rH6+IKwG3otGKnpokYv+aPqAgiCsm8+lRO86RK1LcU4
nFwwA2z+vzheAZ1f6DrNI11DGruHvlcVIH9dSVTzGJshENHmpPZk7htxM7PIGOg5
N4hZJoAkGPAR+bQKx7N3CnChn3rWzA2QnhogBR45sU7CLc9pbWRZDzj8+UStDuut
UghayKvjgscWoYNgyrF5PC/g/hPf9kE0JBsYbllg/rzd8MYERCofcJep0xaI5Bhg
5gRX0bxlU2ayX6MiPwtwrw58RNvBb2Y42kiv4Ah3abzHpzrnZoRebEMj0KlGgF6Q
K+jVuw3mF+ALQ7taxAJ7I5G9zyjIE4m1uSJdlPjA/7DlROOfysNNdc9I0H7XKzOe
PdH2B4G+TrgKneF/8fGy4TKVR/J2T2xpKgDhyceR7Y0BeUkThbXQw2AlqYzAgP/L
OOwjbaniUsxSokIxEWLItB0bkbgFYDXrCemLTns+VXh7tK/rmZ3E3WR/mxWLiFUl
5sIIgY0arOtkTHmHiBGULwCYZtwOl+698QOJkE82VOq0OBgcwOK8avQQdIG6uFff
MKahMAFwv7Nc3ApQsF0owKiezIZv76GtF4o/3813YyV9wAeqAOS46FZMFuOMc8Ku
YK9AJxr3p2Z2PcEXAF+OB3VTJ4j7goyQoX+q4v/lXPM10qiKwgHmdX3eKdAcqPqb
dEQNrI8XZdtd80M3RBDJMBZ0XkKH1MkKdqKgKrGfuqIUlQzRMe9n8fBsQR6339/+
RLfk0K0GQs3eWfgS0jajss93Nuxd2PrZvSs0na4xJSuunC3OvagzAx+/i/TFppbg
27apYEG4mY82YPC3X52jbrYpnspJowXAhkMg7KZpeMT7sryRV7iVEvyPO876Vtut
++kIDJDzazffu2ncIvLJRRRvlpQtmEtsL5OMYyt4ZIKcp5M8ak6VFveqKmelxUA7
K3M9veqaEuE0vgGsqpAeROeu+lkLE094qmEHhiHl8AYVV/u3XUKM8OVCffOg7wWX
h1HpPMhBrBUPR+4JzFG8OsRIqB/X1tj1FjKeoiW2Rqd4rp63p0Zm8nPtD0pWb6u2
RkJ3ulvr0jjg4LS9+nGw9v850O4IvpgT4mTOMPBI4VpvknOr6nx1vjSsvA7zqe5t
j7+hwQvWv1A0NbFcQWUMX3brZAfJm9YRrZpBaz6KmSwk9mXpkc6oRv0E6yRd9Igw
7CJz9ibr6BzmKSYK9ztbe2IvsTcvydzs2dpa9IirVTh0Kijqn2dOSqws+lWr4V0f
jbnGaVkWuoFJwLm90bJtOaKB7d6mjPQGxdC0ON+wyaCJhmNQskTDktSIe1ZlKLIZ
iw5ck98ppGykKzBDmh/i+FO0EnbiFVM0ufGx+AXlt8zlGeptHuteZ6c6xbXf7YFI
0CIhxN293G0imrTJSU+UH3tpWVzPqfUOZp8XD25lOkclf8IpHH5oZpgVj8PvaZOi
eL/zVB6IHGAxUd8fvT2YwLuQ7GqhnC7MBQdAYxRayXt/iLUgIHvtwXxmfkCaLEzL
omsw3htyuu8tj3qg/heZPbhhkSqsjR4ezCFUoWT97dcnheOrQqmA9fFBEPJylAoC
53Vaa6SVpOpXsDIR9qOo3MRweB2LyTQxdrXjk/S2IuHW+9pvUt3WAPrkTk6oKePv
xd1VvcNG+9aro3ZW6RmycWYP/ozGrxBa0NA4kFKqybpKq9Pq4iibsePcRlQP0vVJ
C3htDnfd3OpL9ujwqSEew08Fn7+BqIRKP++Eo9yUI9H+MR7X8LnWO6e6rg3pU55M
DJs6yrz3X3M10AV8nNmcxr7Jc0M0cYgUraYq6z0BZmxeCDqrVV8iRZjFCHrpez64
qJQBjBo/kt5woSdnkK4WVr9Z/5/5xZ7FC3xsWdC4OEqxJJ69KIJA7La8dYCCR2Km
A1+Nue8fNsN4w+S0Cu9MmW3RVFx5ceWv1rM2Y6/kOf7byk/m62u2J/O8Pee9py4y
IY+dmqUGBy7G6mljQ7mUIa7sfd/0WbXGxbJjlzZVc22HLQT4N0ZZq/kscqt2fGW7
q8g+eHcy98yHWj+Hb3Zw1qtpCfz/MG+VKeVSDQ4+Q73N6p6Wo2GN6zuN9VOr+8oy
aaimW+UoksoAbvYO9lSC08ImEDtUeCGkddJaxLBkRrn7mLtPJ6c0Vd2he8hgUTA8
wpIIBdQ1eO8bc3uEuq/yimGnc0MxlUobud2h0AFEi7P2axPpfAzdotMt/kaf2YTJ
S4sRHPXQ/kdHxlywblCmNffQeZri8sI6pb96TrMhhsl9S8pNFyfNdp351JgCQC+F
DGm25AtgqZkGRVDZ5lg5uK+D5dJhVr15RR5mGXBxDtFngW+C7vO92AB4JBeuCftX
5GYySqOZ8n/WjaEq6INgh7hnMUbFwcBAORbCyOGXjxyOHTggfrUVY4Rpi33hKw/X
bCkEOzbz700D6LZQmx8IirenP0YaN6kSrdKu5hwcPuVfafoPbdesU+TBoqueFGAZ
zmn6G426pURHjEa5z/z83QPuOZzVOCl3auBjT9QqbYS/UcN5WFYYMDrQC1m9ssfR
rt/BSKDEeofpd4IqJ87F9bAGD4N/4/JX1CUjXoBjyCK7l5RgiZK7hgjVA0ZNyK+c
dpjTNs0vTvggnYmCb2HCSZbQE847qLy4zuR5JGXWZmFtvznEa+wXYUa7dR77o60k
6IB6qqOY0yLWUGlqh+/e5h5B/kpfCDK5ftfii7HqwRMMsAekyvRqplrH8Y3Yx+Rf
OKw4xTh6y1rgPZzaUmE/zp20VRDm+fUc0OzyFkjxYeyMY/xVmZRQCgSyOuqo24un
wTHxHRQkAzvwVBcYVCCOjIoaNVmwqlxcdPIvVvGpeFur5tRvVIzGy1bFOLpMHlYa
JSZimlMEbCjLEse/rG+iuoMhGHPg38wRIMqsHDK11gbgLYTPxHXiEKdc1aouM/uT
Fsrpt+caKBtieAeRyVczXH5lNMwN0lwEXEkWOYOV91HPK86GVqIFcXuCX0fmruhv
zO6YbvnugetNYkeIN/xNQ16N/87W+cjp+ousZ3Bx+yVjOp3dRgTVU1RX4KVhPjpH
4pvkAZ1PWX1/Ho3pvEqGswKJHA65s8JA2EnMaPWYtay4VkFin5HDT2Ky8HmfA3qy
6XrgTUYOFBEoP1A3WbHCWBFBxrCjTRsEVFLb4a4KeFNA4kHPSYBeVakHEzrCfcUv
ywkLaMWu96yEmai1qGeN/GXaGKsIWX64NsJhJ6aVB0pWD45iJ/yTSQpROQanBuVi
miHEWv5CpQ+wcXMgopo+SKgsf/ITuScfzJ4CQrk60i9wxaFlliospBNBbg39zyA2
LT0R8xnMLscajGtXua8L7RWwIpwYmq9X5w3OS4+ZNInzqmGjmWaQumBbVwb6MVjc
sDl5exl7Bc2g1Wi9XfhQ2fHqltrCkDP8NiegB+DHeKm7E2tEgz0xM+PhVmLZ/mv/
/XAiSelEsblCYlRo/hdjYUefYhNDXEhDA0MtUz5v9XZ/S4QrRsXFzVz5XFTsDviF
aS1qF392dgaoEW5SgVju6ANbPLUCIM9Z8CRSyg7wlak8hZPv/mkQbBd5oL70aYm7
8tt42XDHdND8odESuI5E1PlWqNK9/HfNCNvj81szk5lMQsiwuUVaWzipiLCQjbGE
Uq7cDUJb8etlj9POviCxnCCnfps3GtC0Wkdz0XnQgxHIcMyvWDF8uADKW7RLtpA/
QSQLdzIvhWCvz1IrNeiG2vlUwwazVhdvv59KE/UWrsduZ5Kb+0ju1j29GTs0xskk
zuko8gWkNCkg0nWVgAzYBnuoKRw4gLLVgs+5Y3jPHiKHhUj0EtY6MAaZdRUtkxTh
6zCkrECdqW0yzvRGYi0X0QHY7ESsWV71IvYzUIhQ51342JYEp0RWgeCGh8s8kscZ
W4cn4eK7yJnq0xt1dOrOL6ga3T5dQ2uIRUyXlNV+FJEDcSkVVliSqGQmhUBaEdVv
aD8JFEK87n91RtwVR+pVz/TDGqU9ZgRRS3+Jm6GJNK5VZtFiBwTNIIaj3fMXIq2d
p7NH59LZEanTuexg+oaKVcIcJHkzlor1N6nmzJ/QaVPV4Imro7iaSS/uGdb3NbGf
RcFeOF3pJOoqxczLIcQlBENU+IK9dKU7lZuAvV4RVa1yt9eX8dEphZL2+RQXDU+u
bVF7S6JOePDuOI+Pu4N/DCAGDYsNQZrCH0huAiL4D+dEGq2AETQgYLVIvwgBaG/L
BCSYPww8nhkenS2Cr3jKdI6owq+n82gkwieo6pQK7lYJa1t1s+G67IuK5InFn9Su
ks6dw03qSivRzW1hODY0DLC6eFDK5hTPxRdOvCUQdjQSz7T8oX6idXfjJGdKji2y
dUW3Qnteb75h2v/7PHEOSktv7bb20yGcHgpwEFPi/sO4fbhpN5WQ2KaCZpP7s2YN
g34zpoKCDzbFavnEi3S240+vzqtet+NI7JS4whaeF6vqF7DI8qtxieym7/SWj1n8
XiCVA2T/k/iAmy9hiDd3pEZDpMuDpEDzbmr4t2VOkz/0BQJQJumGroA47E6Wv+5l
WC90PwpsvfnQOxyYRAyBIi0xtP93WQBsyElx+BvD8RUZf9Rdv2gBhJiwu5EQisHK
faQyrFhHT0D5ZDfusYSWR8mEPLuWz0vaOj1WfTLvRpWQfyV8ZIyPC1zDoMNRd5WS
SZU9OTWHq82L0cYfljrOju5ajr+4TeeXqVEWFtgtzaYXyS484QTRbmbrGISMBCJe
+OU6Fu8mfOoEBACTXl19+mEj4+AfEIDcI/QvnN++seuEDTn1TRv3dCdS4YCudNjC
RaXySazjf/ZJ1NC2sU3pqwiF1NCNKKS647jv2YR1KDNNrZckYTw2qrwPl8WRZNWQ
1o21nuE683n8fbmiys0uR5bcpMjHcDk1Xthpe9lm6NOMB2X0QfbaNxBl7Rn+2VPE
SlVyVrgrhDD5QvI6uT/kAzNtKcmrvvcK62oaAJfrVkrDO18iNAiDt+JEU4OmTFjb
LQSUxdL/wTuGW+KB/zOD/kBSgdiGBmr43Svt+69/FajqxIoA1CeVZF2LewPfMB3A
Jv9qTqxG+CUGLNs7VPz08dRqVSNWtIGltMQ8po27ugz9IT5gtbU0cZSpnxiYDuHi
9SMozEKVD3rU+tLawTGnuTMK+SptqdTtRXraHqiFYJOrnIBZ/mXTKtlTyb3LaGTn
ZVK9K1qKwZ+0PFA1lXSHIDEDgmM/NtNEYAlC7kYmWWoLroJspJaYVW3l6gMdxU6f
wFekSAPZM/B076aWvT0HrNH4vquMLnkkg24V8+meoT2w+OSDgPDACZTX4MaA6V9K
Aw2tn/yG/387bgy6u5hFlVg6iLRFLAza40Zsrkzndz7wjEoe1wk6N3xQv4l3Vrf9
sCf0hXpBxpPnUFYX8+r16ySd0t9hSpK8D0wIxQNRXiatsVHZA8mfz79Y79q0lRjB
kxY40YBQzzm/r4J+AzhYeXE6s194uF+FFBv4GjGICBP2lPl2vsdN8IfIe2OHy76Z
PeNlGqJMGaL9he3kOTiSKGm0gPqJ233dfAyUEkhkURHoi6Hi06IAipwl0imXpYf5
3zqHLaZKge9baRQfeBE9sPustPRh7Mbs2JmHl4Eh/zJjmR3yQyYKfOhc9s7Nfqov
r0+UZF7YYwGSZEgjFYwmv0wz9tYtpS/RBwwVbNmv5zl/k5xr+ERtfM3NvYOc7Pns
MoBybmY8PL0MxrBmlzdbSn6mlM6yJN1LEaZsGV2ts6TbIllDs2qJMZEpkuT7jwuP
0CL1jiGaHLeS0DPjEhvWSuJ08ObuXPptC5IB2Mdli6MJbQE70u55s/+zhtKSpTMH
jOKcq0HPGJk9wqoSaxmDJIrlROncHmpOR0s9QGrlPakjnyMHSScsptgDXrttZg0i
xOZjoLE4sIn+Q882Ru+rqviXPoZoVcMLZGtiDrGaIp9Z34DgZZlYdEZ9A1qzsPhE
LhyaBqdNC71CCO5Kveilw7sh6ln0HC4b2AmYRpTAUjuCW+tCNViwbTKG56I0hq5T
5KZZSPZs1ByXUcuFFXwp9ijpuCylNSmC3f6oJP1312d0r4jqNRZakVKqHFKwijLN
puyOn0D387MOqtUA//uyQD8aL3CZNdqNNCiyvyf20YO9OHt5DTvKT59YiyjCm2Eh
ZqiaLcnZPYjmc3rEijFcKFA+H//XvKbHTLIoD5v/GSLUdC0ssNpQkkPnWhhFbgDH
byPiUZ+sxD99ivo87AMp67coLsQntTtGsdf9jD7OL4USUwY55vUTvOs9fvTULtV9
UyXxSqSOd7Zbl8+BxjTx/BGjjs9eSqOT1UdSvx1vPbqcv6Xjgrs3DMQrxAgEVrAR
geAaII9pMARp1okaTZtzvn+FVQZxnUuDwo7QRQ5Ka7HhbO+nBz7IRL2cSiVbfdGT
JRTm4g/UJZ/Zpx3yNtuREZ4Z4vfLzWZS+96E7hV7tp9fg1oDz8BcOirzsdjEFPNv
Dp6Nt/y0QeK7gvvqIWP/XnMj+I4BxKDOSx/F6qT8tEOH/v/g8MFWmS2LB893ciA8
h78Ts7XVZYQR8xlEX6szlJaNvxmZlHKwKQla7PpPOczTxme9WzMHwvHtZIMslPd/
0NS/N1+nnvdaD+a/wawCcNBkZcZQmwCPqMEI5tudu91RPLJX3jbz6/sI4Oi/G95P
IHB1B6IMw0elFEKV81L/gKcHcM0R3ebPVZJVT0Ya1v/XrCNAOjUBpHUu1PVCXjTq
Gs9iNJyhUXinDtYc7sPdTPZ6FqS6/NkzJy9J3Qst9wxVeSSaOjD+yDNTjQG/hNcz
PdT2bhXZwJbiCd7/QioGbnLc9yNkoRmrxeeyscn9cIoFqajxnd53kgzJpOqqQc3E
yCdrTF/UCdptVJKnnJzWtlVSTsQt96KvqfIf6B08o5j2aoW7cjGbzMlX1wdsV+q0
iuqc1smCFEyKLg+3ACKLJNPVy7IlBszzro59jQQ3oKdJ/D0jBa3iE1Xj+UkObCNx
PAmBAFwyCrzledUe0yzWXe3Gq9qhcUIWYjZ3aN5txbiYw/s0lSsShOzDocnYRgA4
SxmssG1IDLTOYgru2PC9Q5xcI/uvu9FG9SgwZxd2/+qVc91RvdnMF2hac/lZYCiS
CPfyvPTJ99TPjq/hUoyK0SjaOBxa/dc2Wa64zBOOufV4PpJK+O6fOU7gm5yio5oT
LxwU6ibYviJqqEKaVJtEJZQVmReqekIEMyaE+woNq8Q83zD87gwb9dEc/EwEc15R
J3D5gRKYEwQbiObDvlL4oORFj3o5opVSBoA4gctCkywe5ODr+eeFpC8NxIWc14zg
zr6B66plcxNJyOnpbIThFl2pZmqzYBXLbu1xHANd8zYKXTb6BQbvzg6m45QVam7P
za464Duru4G+PtbnWC08TCimTAF65jHruOzQCvxldnKjStkQctxVkU/Tv9jEb6gf
HwXMD5NzgPV6eevPWZymnYUSAyrYMp3aU4LQgeJTljwO1an94IRtfxeWXKlyht28
CbkxvJZFL2VT8+jbKonc3Tf8vDazlZng4YhACy2mAZ68ULrWu26o+DdVDw0Q4APW
pa5nbCiqwUVbLvQ6CwD7ucnzJMefxfMCEL/6nCrMvUhfYF5koazmt81EHjb6L1Vj
10hdwFraHOlG3iTQdrQNsZ1MPi5cdhpgbBS4FUHPs03BtbP97ZoO74bxDK7wbl5Q
aCgtHEwqcMFdgqoh0Tg7BUEzc2p1ygs0UByeJDGi9VbGKYhh2PnHFRhicKSZWCGs
Pi5Uo3qgYxEYTIGfgd14Dsz5Go47kbv7Vp8uSZRv803SmVoG4nyx7ma/CU/A6rM7
Vq5T+HPUz3N4g6wlbM6xId9wuHikEuKLihJoAVNccWDM+JKgAUf/r+JMlOBA5LLa
tfWEnOwZ2ru6Xhm2jhEpxNAOqAgkUv/w9qL4o/6A66USlYsjrFXn3pzyHNof+jpV
AtAa6qNkMAUFrZjM3Zz7M4ytC0XYaofcaJ49hnkchDbn8psa31gqmbw3jMUWJG2q
LgGaLlYTKTTPLNsO7WGuydk5JqFWGc9ONpNyKQDKWOlxHS6wtzqg1H/4LW5k739l
b6BnwUEDZBhsKqDCCDkTKEH8bZQNc375rDKvdmSXYBp/UxnNkNjUfuFiBpgK6TrS
xV48vztpwscZTLbz50x4mQnzzxs8Jz3ZqKaQdGP31UhYaJqGLn15ei50IsmpjUFn
jaiY0iicJIMSpe/FaiFbhUJnfC5r8PqfkWxVthy6XTCLoP7Eccjtst2Og2rcxKnW
Gv/XjTXPHuZs5J5xvpsYdExQJ61yYkYUzzAHj/r2GJFK0aaxHNMIOOI4glsWNP4v
J9HrrLF2ykR7UWFeKVXR47srDdS5YfI8epq3JJPjKSLlktJjobMdBGKSTU6ZTI/i
MwO4FudcSjpbgJnt8jiTShif3AaFLadaUOJE6KSF5DhSLmGxN6YOeu7ZVMvVkDhR
VM4qz65lM8peZmU1kGetl6r10lY5jXZlMQ2TI6vMedrp/vbr5q7RgQ6zw1QrTJmB
SvH8k1EUPKLzewE6kpuf2viCBIpadF95yyRtCY59mfh2hs+lGAsEe3EeCV5HdJEh
u8utMiFgA7lJT4qeAq1txFKpuzy63b9tptC9d59scPEtzPQKunU0FS75HIIA6J11
ii6Z1R25Pf/LnYTutnx4UV2odNJc9N720KkcVmh0Z0+7DKscCg3WfmV1D4O1zcSp
KZVHcRzb84T3+UaQ8mUY6I3ltJP/b2FSSCecH1+qBrQIeTiRwHq7DQFRf+JsA7mP
G/FRYd4DRjv56gbA1uC/nuxnucwpdJH+4irAv70sX3MxRzERsZy2s+fdoqkB1AXE
ATYruPU3siyeqtSWKOLfZ7XIc1AGcIEFUl0p3Cw7xjWCArjCiAHeBD0JKQIagmCe
jqouWU+UquzTLaNAk70pczURAYQH+LUtNd/+cYfvaI+MWItOrUYJoTgA2TaNCTFK
a2STTD7iTZi6Sy64iTUjWqLQ+vAH2bCQpbyfHkcBZ62b2NkVm9W1sGPWlD+tBojd
QGvMhjrA34TTGiJTlfF5GNWygzojV2qd4YeSJxCdF3qP6Omr86doM9HFocY4jvlR
nlOqMKXVF3WYyCFpv6dmr1hafHRTEg0pTY5I3/986W20BV8gKJWhSirdiNlots2q
LfnEklNCHjK1HwSSwJq677bIzcIXNJiUxnplHWqQGvWZcMJVrMyertW1iFFMX8oL
K0/OZo64dKySbOltAu1btG1/tvrys++uyhmx92phEJnOx9UaQ5FrcVxJiGwCn38p
rzSM9zZ1xnJshwJSotzxTTKlc+XshGm4+abyUM7QtTwQqANULzU5lWyDfofOmOpS
p9HkFGsqCM5RiHmqDfCXtousYDY7mnIdG1JozVg1AeM0tBn/y7ukj3yiOxahMcHU
ncVRQv7W6vLHxrLrvSkclvuZmazTOTeBl+AwHwt4AbRy0xe3NuyelOnyiFSqtbKh
Lox7R2yM6ylyw/Wnsv71F8dCypB6QefoaljN+o6QAtVAyFXYqeU2JyqYrJCSKOoy
2Z1WE4JjvRB/oyy/RmCbEO2uwoHEQP9XWCW1kqtwoS4IcTuNpyEXJdRgnSjBnJGa
o3KwzO4fo+CQ27x6O4WuU1T4+tEaV77wMOUnqwE3IHWJY9zFczjfsICytP6b2JC/
OPuM+Rqwzuom6JGBHXhjF2vDprIjwoh86fURPArCjvWWGn+HRaZJ9uAcv9i60Bbc
4mM5j3ftQYIMIpXGdnhLmg0cMvDnVYYB3Dt+LXwFnshYWADFgUV4fDbrIo6NomHu
psSDq1d34PbgGw6iNRgHemwAJwdC54j6KY6ONLHBYvOmEgolRdl3WuSd00HTZ45A
KF6m/Qk6NwUSEBa0tvnnd3ArT2ZzWE3y8iANjnzTtMRKx/edVWp4mU0wBrUHxHo2
plSMn+jQITxhHbEGWMncSiPDiFC3aQ10zcNYrVufzqIjvE7FJDk0dNA+5dtQzfcj
+aKaFdDud5OAc32jANa2sv/gajB9A1sSi+2AQi3LfAlT6pD4n6ajNP50YtdXBaWK
mdoSHp7xpNCQ1wg7cyqPRc3liGefqiYQMltJf3mM29sU3zfoVBPJrsmNBEfweGl8
hR5XQBA35FxecdNvwgoNPabnZfGq9U/g8XzGtzF878nE0SGnt6+cTNIj9QeC6rOp
MxsHQhLdUMrUc3Fj6HCPh9CBGjyXwABhZLy6bMjOhCZhaoyfbVHZQX5LMI6P4hIB
jIVv2zJqK6Ku7njVnbjf57xqpXnMV7wOsMMldGecDs50L9sKcz7x8KwDcXvpvfjA
5MhkthK9sOKBvwFlU5Xra2JsXC6ggP7fqxHv3XByVae14bZad41yWu59uFlbX3eg
5oWZQC/7xuFDR1hsXAqGBwdGP0/oFI9aIddMms6dD7Dyr/pEjx4BvbsbXG+RiTm4
rceGz4Uc1rpYfPVXV15i77pk1LeUonHNo44gVmS+45SKvUERaIBpg70q1/iixbpj
pjIFhIaMSIehcxZbMQmpFyscRyATdDFa8zEg2FOtn5H2Xh4CkGaglgcA3+m81Hkw
2oixz0Y7TPSQXvM+zkpaeS838RMa/ufDXz/j1YVUiI4hnqOVdtJk34KjwysRM+Lx
d2VOCsiuhErLvTmr/cQzAE3ttEOI0cIn9hA/wukG3q6ICGuC/8mqpLX/d6CDrCK5
FBBGzqIwAH+7d6oHe1/GumDJCJe89OHn9WvjB9elQBwEyHw8+bLXv+6DUK4o2qrL
cmQLGE/2iooXeG4NlnnleKeldqT8h+RE2CishQqIJDnBiVbC/L5vXHZ/wreWY0Vz
IGfRgvlpw903VzMfvQS/iQRHajFuEE0pPd0vE5cKD9muPw/3hP4HidVH5JDZ9+F9
Y9DUySpKu8P+av9k6xHLkpuKD096z0LtZEAOGN+cL0xSlBxZ4T3Q+tEvfuCAxcEc
aDFTWh9B95DRtZmuX4C/zimy+aIY7vXwfTgZdD5PKDmGqayvnSs0QFTOJgqjYuLK
eKXzR7HRTBZyTcd7FfMMfOz8IlHmxGp88EIKMokS+GVgnZa/qMu1KdB+FAIJlc2G
uiXdwaoK447xMSvntJL0frhkAclwg5fZJgI4TQAno42fIeF0jpdSTt6E6kkG9r8F
P9JhMl1S3mIaGYLkQaswuk84GVc8sLE+3N14poo4duQgBL0ZwaoY7pP+h6k0Jefx
5yGsiFko76auk5LQENW9aXFZQDl/bIMbU3/BlsLkpQl5wms1XkDb4+/fr1oPQLLl
3hthkevgz/vOFpEs/yo3WwkI7DO8ebe8ohFYsBnzw+4JNKUz1kaYQunpRRXFEtwJ
ep8bJZPVhhm8Y0kd85ojd9KeIzKA9Co8yw1P0K2mo+XCTiLBwqptZlas9jrMXct7
+2RHGhWbMyMwRY/AvUYPpNza+Tpbe4xRa+ad89iuS77oU/n2SgqT48h6CBY3s6EO
lJq6KAqVI9rM9nse/kBCQk1A8OoGAnpJBlD6vvOxPHKOgN1D9b24GElxqMyxD7sW
3vbktosdnKIII8tqvSBTRzKytSQzjidGaU6toAYtzDu3h5TWECiIG27cmZcJzOUR
7+QkpX0tl+/w9H2YROaNIEdsc9dTshckBJP/aPtUGdI6ruzSbOritHS9JAkesID+
wx4Y7Vd6iYhz9GfDW5ik2Kn+r5U9rQaFfX5SNWPwQGBxn3RUkdDyPYZITTiT24ag
thr5nIzO59b9l74/MRCMZ/HeHx+IPUAb/mx8IaoeLXG/jgZZnxc0PukjGkV55rLX
iC00ansob6qMHNvwbgNkOJIpEhANkFGdOhfsTkx2mBBH9FT1fD3EueDgYi42bmQr
iyFWbu6/s9HUlrU90RtAGXnuMHwuBdFafMxhlk9z+TsZzpod3IcvY3PjUkSYQW1Y
k0p3v/hRg8h7Wh97CIFyMqpNBrNQFomtz7u+3CawGKciSaSaW9xOQ8E0z3+tZwH1
VmCXs+riLpOEoD3/PhmS1oAV+ilqvzh+x/iRIn1e6bwXF7kApA3P2OkUzrBV4yww
gJCQ/Q2wWGWHaRA393BKJS7HCElGU8LqEU9R+uLqK4Cbp4suCWPLiAZyXb2Hoehn
jnRaKy3DEY+FPVF775AYzs7hzQuDOkW1yv8qF87EVqoLvNd7nrUx6bsMunTdq4na
0PvmjWo3d5x5p5/94N6FhEL6LQYiEWxo+XdB8/g/afMFvTdlNvpOvPuMLNg/q8G5
2n21EpR5Hj/slAKu2A9CPJbW9097Jyr7XTBkxPt46p65gYTPxX48H12IQK9GPNu2
8ZVOQIKV7mI3nYhvzWa2+cLrTQENdjquVrQ3G6DBkldSnzJF49MwxbvywHeb6Cpl
YeEHewiRaly4r1O1BNA6bkTtFnwLfyTLdJ1Y3227TUeTg4D1i7IBsNQ60lKRB0dh
lI/mOIwuWE0s4ZukmGlAa3geGt96tc1G4ygyi1jDdJXn5pbW7ftqMRYlGiBdHxfm
LqTBnbf6TMKQvdNI8CxBhV25B6z1PT7Rm0YHuRbLhz0oiDjvIHX2628MJ1Nd00e8
T+tfOh86fVO9EgWIDXMJBYrF5SUp7AHOqb84GK4Vltn+20BY57H/ZgT4lZcU/6ci
hzBOAW2iO1Avfv71DusLTqQzl59i2ZZu7ehcxw5jZ3oRtFnsYD2D8eWsBMEJ1Qla
Ysh/qX5E+u2Vy9KQ4cXZIG+1Nxo4veVTcDOodHCJQgsXvYKd/3zoYM78//8Epv11
UJH/zNlP5njHk5x4evQlJefWynA5dIYEZyQZ/f/QgVDw6aM/gRmbLQ8uiJWq1iC+
6bNRyorbEPLK2Sx140+nQ1R1y6WGffx7aiWUMV3cCMIsk4EE6c/sxuWaRThJCeHu
kgrVVmbUDntRsuWJ+Utn4S2bXcwVIYlr7VbtYCYsTqJDIOGG0K8nVHB+m9/MrhjJ
cb2Mt0wCUffvWh04KXFNACNuvt7HTRWxNFNKTFRmbNKvwND+/pmbfbdKN5fr5bUf
KmgVsnNfMOzQ+Kq3U+UU8bxWuYJZB3Do9Tsgsi1uPLn4IO7AE+MZ2KdOEY88ndhB
Bhlyr8ZoE6JhjSqGEmqKO1Q3yo3usRPQjAknrf0F1+cSvFkK+e7n53z1IPNt68jz
ycmi3QGBbT2/Gy8wJE1mPT5V7uwButH6n5tGb0AyvJn9mAZ+W6ORIrkw3zTMRQPO
QNJmd9fH3URYrDQMNpS99Co6hvhYX6zu6Ww/Kj3IgS4Ey+1hbJrS0+8x12kqL6L5
t6lFzyq0CuQu0zlux/2Q+yvyu0C63y5x0hS6tHxw53LVI6aygSq2y87nKlduidzu
MSDwL8JPnVdCyN6ImTdMswIhANAhKj/Ep8V/KZ7HCh1cPmLSjJ9wQFDvRRg4BHo2
8lIG+cPXo4N4Ub9n8w5KBOpWfTJQ0IBOPjCXp0xiw3WdkPu9TB4Pq5A81W9Heeup
9Pd1hRNn+vDcMFcsFiGcbzPRDlMt9dlTEHncG9M/bpEnWY1YzM+VwOK4JhzkeVdm
J3Jeq+13S2ohB2pVw+XgsA1XhDeXP2RalFcF13Xg328DKLkCsW4pKQkRpEKr+Apl
n1bHp9EtA74yjGoZrixk1BAmIg6wg6J8mQFCvOqRzyDCaEizF0TalBjT6URIp22N
lWld8LniTJTPNjX2LQf5yKZJt17TZY9lrPHt1f6GlEc3XpCds+sZb09/TwmurE11
Jp5Ha5hOBDzctVGg+wHmcF/mMUiJyOnXUs03MPfqUhUvrME7NrGtoG5PP7uH34xv
uSlVCPva+ZZgJ1s3kUNI/Vxzf89CM9GzrYpwte167g2ZgkHDHjNpNSMu9GqwJgla
Hjk97X26WxT2JC3XXrvk80yELx+pqWjrT8ERhmmnUoIwJXr0G0PfhVXWnjxGqGgy
At8VuDxkxfVQ2i01JsNxC0cQMcerimgCfIetpENRu6UeHsfF1haPg3Ywricmwx55
s++crXum6In4HQLHmBezxOqJ3kX7L9S1yj72S97idb1WeS4vRLauwocWjiqat+ZD
AuJH73xITr72HsSugZZvjnKm3ZRMP5BS1gcGz2DxJ7mTZ5Uzju63ij9+wlN9MEUA
GUJeIEKDvFCpeObL09cBWGXXH+rWppCG9+u6YMMTuNKFZbRBOVvNCUcPar60V9Xr
nRi3cpNZPEoIzgXRbBL5C0dvTIaZnQeYWGXbQrYVlquOaXEfOEE9vMNxFT7YfO/t
zdFgzWyXmyr/CbxENJJOiBAnJcSz9fDVQbds+7qBvy6IW8sNGrjrYmJsHwIkAdNa
WCPp+IGSHBmwtjsO6UVtbowbQUurECMZbRD0BMMjMWNvTFPKpFccbpLkmYYpfu2H
BuQYEiOOOClOK5DQ/RIiHHwMjAhPvjHljS7177215XF2PiZFPYXubDdzi9rJOFxC
Yx6RTDozb6Eu5BiZNJUQXclhKqiL9li9RNIODjeTNkD/t3WQqbiqF4GrIx4bEriP
QSSGZjoBOYSa0dHZvPjIxMxzKizxo8uOLy4LRub5XPnXz0igwikWCxlTcGAoZyPL
cTpOskKuN3c2p2YD/rfuerdZ74LiH/OG92Pf3tUv45SoXS7ak68qOchZper3IxB+
0fBhFhzGtMEAKzNsqoFvVjU1WaSonQPIA+IEeqTpHbUzOeLBPabXBBSk5gd0VvC5
n/s5qcEIj0H9xcw62cgnrAnXsVS0CryXAQ0rpOFO7DrHN2VW3zxakzJyTcH9jeQN
1Sr+quh3Tm6B7umFJs3XOt2RI3huHXmq1mESWggncqtkY8dxQb0t75usYvIF3gBy
A8C8lISh0goDUZ9mYT0EPgaBWAyHS27zBEYXUjHe7m3ZMl8GYmtcoGlW1b1X1vMu
hvONqosUfbjZEePSoa3f6ODU7sM+YoPIsLekzdyzulosqDLOInLXbR31c3ObCX4q
GG4NeU3fFkR0aXcAU4vK8DypgC23o4zy8OcWTiZmZ/+Z363aHPk5LPc+dhAeFySU
fXGNOT1ibLmEKRubIcrnslZdLpESq9S/2TvFkBJaKPoyhx8cBGZ8QVCJfNZxSdm+
Kh3xHqHJ2UW/cdDQaqf9dBofM5+a3r5+0+w0HLB9yelc3rkv/phnRSx1hoxuxWb/
iS4YYUhzOwuxUPZ8XMwLAehT9ZzRbRPx4rIxR/2VfNpDy52hzPd2/VdSuYSpF8Pv
O+qb8xx7LLgMLAdRqOTJbVQPD2gaCmJ2S8Hf9klLANz5wyy5JIfNJlUuu1G7xmJ3
aXNsIMegwx0L79wzuN8FP31LgcWLxi/J2zHNqM4F9Pc9TWHtYRj8c27ByDBiRPHi
tDlfAtxk1Cm8MdQovzB0rNFefxq0ek0xVs2gZHm2xaekEANV/91eodzFVQhjIr40
NnhSua+wKr0wif74XsElCN196Set6863vg4DHqmGV4zD5KnCQRss0GflTTUgTyHY
hjLjq9cuRD3NvZ+W/FxvmxB6ehArj6f9RWs5D9c4WV6RBuSFtD2Pp/2ZoaTb2qvf
WDx79BU/Ik/WkBmHSwVPwSWMEd7NU9sLaWolGUG/BG6vcfNcDXBG6lNWacChUDH3
oJFLJassg85AYWmB432s4OYgHGJibigjBVnu+0Re+3zXTnVedrCxMMEiTgEe+eo7
2lBUmSX/Dsy7nAy9tvuOA+4ZvjoJyid45wPDFG2As+hmasaDEGZyKWq9K6oqvkWT
Aa+xaTh6jL9j5SUkL0tmcZXCkpaAGCQeHkdbVXKtov1jN7BERpggsoQngyvId33I
6xhSGPfbt1j+skpy8DoGrvFnALpXsMbz1d1pNH9ggDyn6EkqbzGNwEq1cWpBHtpp
PHP3n+uKDmFEv4UGN69iTik7f5p8UgeX4KGV1NDcX8ajueUjCE8jYDyMq7sXbf5W
acXwk+DSyPQ6MV7KpvWyswj7nWiZMkKbsfvlIjnC7CF/cpHqNOSiur++RkfqdWIG
pWqNtytVKatBuPilqX0IcBCdQiTe7/XtC4wRxFcOf+aU3voTMd5H9FX45UQMOceC
T8L/89OV1XWCQtn1MQd9W0SoprPqtaQX+a7AolMoymP6I5QzFZaAjTy6swoWdK9V
e/6sJbYi+Aj/NN0UUt/G0rvOGMo3ygkVQA8Cv0O9AGuT0d9sn5e5EEmm/1pwV/bK
ttcoqxbChJDBGBsPXqeUpKPVBKPu7CAAATff8g9F3YjBmG84XYE5zJlVFNy5Pnjn
h7ST80afKwRh7Pt4ghOYDEwz/H4AEos7tOTwr6a/KHG8VyWd8EPM9BV6bRiWgPYH
NXiL50THMj5+ny7qW/Odon1E/viJHq5DLdnOU0cnFqhHWMARmdNctgo8gYa2oc0s
9K35EscewTH4HCvTt5U1Uw+Omwx8Plf4M+8MMlvYcrQMKPXGEQShb/3CTAb+V3iL
hocboBbjWAZI9ApLFVONkeMj7h4RYuBvr4mQHfxQpH5QXXqTDDtYjbzNVCa7+O0H
AqwXw9v6jHGK8piyTwhV4P19I/3gnnBX2qzApb+z0B/t3zaXd4sZgVzl7FUmfVX5
mwbHMPiFAN5eMsfzQ0PInXa6m5Lrir5UrCjSDHYR254M6lEMhdHpBjzC7nTISFzn
qcpWcMf5tu9CQNJpX9UXsLormJ9Nukk3u1anAi4p2ZPCtfuLmAetCL31WUOVulWT
3hZ84VBR++8M4yRo/MZ+uIux6O5EU8ydP+Pqsqh2mtEtSvnoiLGKTAlfz2b5k++E
OfkkQ9RRmodbGOunhPyQUEVdlRtW8IbB4csjZBDj5VJxfngyGCmg38urXsKi5CEi
AzDrfm3n94FfUjRcS13quSI71hJD9HvsgSqrlvyV2dbyIERRBc+U7FbCrk5vdc/l
/fvLF1kA4Wh7YzdO6qP1yPxKM2NGd7A8JlL5FspRLGMXaLlwzVtLUQ/rt25MDTW6
ZoGgB7x1CelRxiBwxcZNCeV0dK2wHt7p+xyY4ADXYg9W2PJakIo5qvNvXZeAnTAU
kzQrhi7+kB+npNlwaRBifohBCShuQsscZmQrXu1Ow0O/jyGKNPyvY/mvrM5LIN13
am1usn/j9vHq67AvSpdedKBTqlgmH1OO8/GFj6v5mmIg4tvx5eEqBvLHN4poS9sx
oHfHmbGySxbUfMdN3ClbD7d775k/6wxceVWqxLzS/1HiSyi9FvuB+uklexw0k/Ah
Pv2xuLHsqdTBwHdpgos69j+yzJ/Q5NEJZw9G1Sy+6PaEe7BzoWlo+2IMC3+rdybt
MLz4emJ70m54TnOI9XCP5B3ZvLitLMIsuHsG3TZVeo1XZLRd9WF6g27haUao5ghu
l1s3LPgez1VF6KGjOq83gqQKVkv/QWKPTQlFlIx4dwVxL6FGMYaFGMp+D1PoNUGt
6yrsp3FL6qiaWfMvUB1jtjJgXE2ZcvMujiwiShTrQl8KwnWKgdzX5oi0eSeXIVAE
vSFXYqgCvWOMDErIM16RRYJH06BwnTdsbVcOKlXE/J/DQZNFCJcI4RkX1B8qmy5O
3Puptf1QGNQCYikW4oAtWrQgYk2vocQCxotnBSBlj3e+ai148HsCkqeeplYZ6GHR
BC0bQurld6zvNpNXrHMZs/gLSf3evUoIkBr9abBhb1xAt2lEzR2CS8KxlbtwGhGg
2TV8CKXtdXDUX4gGQk++mJfDpOG4/MRdgMro6NpApbDTDtyQyIPbXKQNbBrXJs9U
ZhvQ2+spNuxuY/bRDrDu+t8CTclYKhXJavSgFCiQcXl3gcV4mz2dJML8IpUl3fz4
MFARevG4mJmPC6QJU5aDqhVgOfcBbECyeWW+fiZ9Xs1+tkx7r/ivGNXgWaJIeOZR
dzTjwGKu6wXKbFX/mcSegt2ogGuzOniHIh2+2USi/Khrqe7nN24xoJmr4UdHqchf
2PtINbqqQMoWqeOjKpB53GpkZjRUiGC250triZY2q8K21UC6zJ2ao0XgL1YhGsQM
IQ7wX74KHkTHAa8vYRu/snyaukuWvXyy1t480PFeyz4yoyjFZ5sSMc7yBvc6sPwQ
pfZ3StB0KNV3zhgRoAGI3DlsP1mPMVS/vaekEcUzipLARgsZr2Xt5qRa+KNCpMp/
+SBmsIc4f86uX093AYJA2NiHhNwsbDlPm83fqUGLd4Ytu6Kieu84h/OAdjcmBz03
q8JLn0F4GK9Jdh9W6m1ctdpHmWR6p8g7WrBt8XkfhQQjcJtfWCOnOIjkXUcvSxaw
7Sikk8chdiUtfm8mHprNp7rXzLhRS5HDB5W417n9KjI3lfwH6yGHOjC+ef2VAgNA
vL48b3nrQFLFpxAXNXQerBU1Bt5Hr14fD5Q+0s4jAI5gLRW1J+mk19RnyZnh+AVi
7FyBH7RBhOawTujlnTwHfIYu4lra9qcXz/7IJeOzUXXdG2E9J+27iNB9+y2I53al
wWMYlwhv7WkHWDsopxJpLY5KBHgMBz1mo9Ww2Hz9cK3S9cDgDRUUMDiTA6NHm/dx
4mZ6144Q8aUxaTjrBoKGl8QV1s5pF4of81TZNs+fPwI1K0s3lK56H8M3srTPZv43
VGMJ7mHMNrCu+UtDp5kXtzIOCmvu4F7h6V8mRmL8ubIuH/GPDoJwzKCWsSPJkeF+
L9tXDMvpFogSeyT41W0AIiyLQ2w70ZNUuJ8IOAzGVqAzKJvv6EKmBKDVNyg8MltF
uswPR6QxFKyof9qGM7FOWr0+UHjWjitWuM371lEnaPIjAq7Dq4AKgLZsokLa4WQ0
I/WpEBjIjDWt5ol+Mlj82HQQxYGSQ06JtpRCEm2FUIRbPmEqzLd1vhQVl7us+9h1
Yp50wrR1JzgpI6X0ISnPeDl+lirnF8HcZiymveUf9GGGrDIRZx2jpWxkEMyeQcN0
zsEEqQeKZv/+gB5uXbhWtMzXWJi2Ba7R1tlFwQGKtbmjKnmMYbmQ2EtrKvtlq4Xt
kebYntrOSy5pvrpy5ARlijVsmqSSFm40dnheFjJTix7mG4ze2AJdxeYWKGGxHovt
Jtu4WVkOJ6HrfDNBz974v2TEM51zg3biiVnxg2ENE9xaQ2dppjBOLE3+fwH4MIww
HG65S4aBmvGMA35VpD0KjolspIxl1+hK2givnHrW6oNRRX7gs0e53rTV99SvCZlk
naGgkFIOkfQSllKk5z+AxOrkQvFQ+C3H0wyfFZSt/0JJ5w9oFuFoj1p7JE94wy/k
xUpQqq8E23Hm+N6JO95ujSSC5v5RksveQM4JbbpMSHzJE2A/sw6VrPkAz/gqrjcH
HlyhoR0E5/bXcOIy9jFDgrfEuO527IHKW0ErALJ3hXyhVQqm2a/CqqgqLFnz+vc/
Qv8Y+7ZpXsv6qwBo6aqcRe6RUQcOC/YSvBAPjhB4VbzFoXNPtJURNG193e3fVgNs
i41CTmlDCnxf1QTIxfCIXHEfYoaEMm6dXSwbI/VBN8Rw/i5ggPCZPZhpQZdsOucy
bP9mkjkyjgg0Zltrhrw22Sc7mHQdQkGw06W8d032e6yK++awKd14ABcIpsMZNuEF
SjsTbcqNGqhT2njoZB+a4zhArGHbPX/MzBvLRr51XyLpT5XZLE5o4lzOcJO6vEU0
phl7NY87nQeZLYHYECkCuyQuWOns8N+ApdUEXY4IgucKEE6l5UPnvD1N8tNxcLy/
/wZVbWQgFSfn45VBL5uYLXM8mxAydW09aqtwdmcXw+acfA2STVtj3YOhAmAlzGwO
qObLH9mcJqTkuwmeClY1H12KatKeEm2oDgGRUWnBfjMm0xrPxyhIrTlrkco+BEs4
B8cBR9i3ZyMDzoeSvlpuix71m0sYgdtqmlVfnB2NizcIRF8utZxlz1GGE0eIFosi
uGGPEQN/Jo1DA5K+l/Z730BsXrnhUVixjA+qzsqPArWcXPrg5wDcBXaqII8E487c
fSuzTG4odSUOhuvQGt1/nFYW4/0FHzweO4Bxuno/BnkSveJXvY0ALJ6yR3BX0abx
SkxsOYxVuIk2eg6Fs3NFB4SV/hkgaagnXX7/3rr0MiZYMDlxofSatNXPuRtVdC9s
L8mpRnINFwfeHtpdjvdQ0uE9XxzqXvqpcWafZnYhMNaaGGLeLFDgZ3+WOukdT8OB
pVF1J8qUBA4LDDRS+ECvxEuJtUrOosJkLKb48Zx3KZEI+jRBcnSJtpvi4MJJRnnA
3qRl3oYkEGXc2rl+4diuRpUf1lPhxpFpmXzYEKxIySynQDe9jhu+ExMduhHiOz9m
hghiEcEuM8MoBRKLpxIP/QOBUvXM4nnRTN13awCdVQNxBVBxa5ZhiuDSBgxnqPMO
mO0TLKRGT5PVis/DxpQp/KcXvIV0Hjxoj2RG+/2wN7tsf3GKTetNMar6NQbLmV4t
/T3uTaPheEWxMkhXBGomKHcWQQoMvnBGoKp3EKu09veqI3HRzAPwP/26bxZ/Be3+
IFPfaMVyyF6fvTl4yzuxHzVKiEYRLjwvix0TTPt7MqOTQ2UL2pnAR7POKq4AURBn
j4f50gnGOBu4FfMJf0Nn5DxE6efNEad8GIBPjtd9JrAIya0lFs6WSmJX2Q2Rpl1h
CHycRbJhyzzoJKI8durOdetY0btip+ca9cfhkwJtfGXtIwp/K7Od6cab04dcTB2+
r8GkOE4vqikjne06CV3g91PJY0SfXV5iA8inTThQhdaTb964ICMGuMUIoboJBLZf
3vADBUcuOs2OGfg6uwkczL4v0vuM1m4k++cVrvtGqKA3KxeqKGfCzbqP/otYxA/S
vPA4EpeYNCkPOpMgDUoZQX1HaCaBg90LqL06nMYK89FzCbOwCXX4c3AtkAJAzjaU
zJwgDer5HjjYuop0SQCm9A5S3MNOp3KUNJz0iMZ+KMPCcrr0f4L8wksircwIRDiq
nD8BDSzd9xLDv3dLyawvoizOl962mSQvYKy17v2V6yzl/6aIMhGFhzbaym0qSYIf
TUFbjCftnAQYCvoKtB3qfUs4Vzoskqcta4yA9oiRIXRSVwDlsHpr5VSyhJP0GcL0
MwXlSaDgW/ern1AnEBROGHHSWRotb0uifPv/IBvF6hHQeaKtrU2bbdcjD0SEq2OL
4IR+taowbQ8SieimDIQeVoamu8/+aVyPVlF/OBi8SZ96m83i2qe2ZVjmrg6NFwHD
0QNl5DsVYF3nhW44fxeAUbSyyF1CoaaCR8lVVFsC4xQ48auLXuW6RDulwqxjIgX9
aZeV1Q4bYpJBRLUx+o+1CMYrvezH5ra/fOuNOD/yBpFznl67YmioX50HKfznMEPh
YSaG7gulvGr1q4sHEPHooSMSFHGKMsjUU8zfZEXVPDTf5bjx1bw19ZBxSamekQDH
aQ6J1uGVMulSAEgRxaO8+xCNhAYAyLmFWd7nbq2W2inrEevQl5wv97jgB97QCLrB
Om3hHVjJT+KysBrKsjfb8+ctCIeXhC0mvsA87DeIi0W/HM48a7fubHbSBIR4uls4
tGqdi5K6QGGNlNLM4rLVGpUamP9h2xBgqaK20Rt74e37r7OPN41iYxF2Lc+boQUo
aSH5aUhy9/z8Nxi2vZhgzXJ1tK8/zZs6vkNMAYNoKZ77VBoLlkWvdsDhYvBWFcvd
zupey3Y7bqs54lQrTT82yWoxVWTIu/BecZL6JHLYzKrp1BHCAleVeV9ZhdOwBS1u
RMMgBfQWZqIzLd6EkIyhhx9phCUOkYdLpJx8tkUu/oRT1Qk3otjjiLpShBFIQ1He
b+DiBTucBbBapQSSEmGLb1MEEBdkSOyNSLhsdlVKswgcmoMNQkpVnPOLHLeOBdJi
RGfAgn++qAJbcbFfFJLuTqCaKhlJEPUs7spmDW4CaJaqI5um8CWheoRhzcLy70FI
IYO+ZnTSFwuC8Zg/wR5iQ1h9ji3/znIKVAPdF9AkeGFYznMpXmeBF1HpEkRfFx6Q
Aovn97HELj/gd9DfmJ7umq9vfS/y1n0lfAtjtQ3purmOWojaj17tVH7gn1Bk2hDi
I1Uff5sz5IgH4P4PZxE984aU/y75ieqpRB6cchENv5vqvf1jwi6iabK0x+GRTpoC
AStIEbgGpi2zvov862eV1vSp9GCbP27lodwmMLdLQTQNq9kx1l6Ks+cTonb245vv
SsOHbS96q7nH5UhWn0H86vUb+EBHBrv5EHw2jmJqoOeulIUrHS/qZ+8VbqZKfTa4
GxLsgp34YqjTLR7wcj9Udz2TGa0x0gQYBz6m0JWf4mjbjpGmQfwWIkCynaRcKVRE
Qz6rMVPKqn/T9IFOEiG9cEHTYkfamFG/6zIIYjKWKD8kA5dBXxDTe1Vfbn+LyhQU
P5XTtcoqJBaoHuR3k8pgEshxLrD0Hvj4c85fqUOiv1BT8Ox7Y+kV1LON3h6dkCgb
VVQl3+GWrfwjIezAbYsG/zUOz48AFsdee0dbCsiD0EppV7V92ZIaqrmCwBkJ/61f
xx81Sy5J5lYj4tJAITfh7nNJ8lq1pyvGi+o/FA3jHGhnMx5H5f1R4GFlI1Mhb7JL
D8EIosgleqt3QTF/V34aBuyx5blLpGD/5hiho3hJcxLKZ/gQ7R22KqEmrH6ccGSn
01sssGOa4YX35NwRmJTtmXPWeaQM25UuOjkI25mM2iGxM/0N0aSkPih0mE20CVxQ
b5EDkkgS19Npqn+Rrdakc89vrqkrtgH1w85Ipb7J93Bz4O7kS/LAcE2rpDYAkjwB
anORxiILLlp8S2E6ZXP/ztRBcxl+UnKvyA7Y0uQIYdE0RE6yrknwyxUCy1KKEq+O
W5UzC7qRbfTowYPvXbgCRwf2l5x/99PesrzfJLU3DvBB3D0VaaTKjINQy4v+zg/w
R1OWCzZb9bvF9UWXu0V20FcCDNURglYW52q9q/cq5FnX2bhFxU6lMvtCv/VwHQtX
e6CP2DO9mYRTiXuCPngO3XXilaZhvzRQA0V8vAat8CSr2Y92KspGsZBdMMCfsVHc
HDpTnM2JMtKdp22kkz4XPuk6Juw3FiKENvszPSQIMNz7+jI6iSZyrK8c9UN2rHRc
Vfg6kZZCtCTC3UsE0aOrxoxc5u/e0b8NkQwIy8MhizsldrchY965P7kgzQ25b5SD
BNSr6ozOPZmtTjerGt+vDuW6f4IDTKFNFW55P0ToVCAQx8NIgjj98p3noSc6JDB0
zHjY9nrPLEtwnQW/eawfklzndDcxA0LOuKKtE0zCpA6ZfwD1ytqyHoivn028w6kS
wUq5fh99U1YHdOoXGetOiDMMUsYfSe4hizbpYE6kQmwnTM6HEPdoNQ6LP0ODoEa6
aY2tDyJSiNPb0c0/5bEsNmbILEeuulTlO/bBzvScTvkXw7/Uzpez+/+h8j++Whdn
l7i8kH6iLojZTdG3lXyIwWf4QERc9u33i1tZP5rAimRvTOW5DuQxmxLbrq7qvuOu
4aJOcZIlRq2inqQDi96HmQUvtSz35sdV1uIQq/O6/9DShhOyQrwJuglksoor0kuu
7yy0rg1SKYgf/pJXHwUCHuZ0KEhz3cRSZYJrw4zetYM7HrcsWhLb5TMhYYzJ/KDF
uu8kPmHxPUNRPWyEC+JVVnaGP2WSsRIFf0kIn+YwjOqZvIQrEFSXOEBm6YLF05l2
ZXEJYwK/7f+NcAg+jXNrluBlCFC42sCO0y0CD23GDRjwwCN+xN8fL8HcK7s4ypeI
OSBiQb9FeY3hhg9Ze7PisYhgHk4CpSiutjb8V2nyTLWLsyS/gF0syzMNQ0/AOHw0
k4c8nSEI/vA+r8+hKJkxF8nnTjWCzUmuAXq4kWzC1V3oFZ2hxCy4T0LMGMzchCaN
6ZiwYqU1Nol+OQjJ/42/ZbEbAKTTiGD+aoxJbDms+z1Cl9JEtr9grqOy6gn6dzNp
5SpMOl8xrc143UdXb2VChyl88qvyh1iIcRjbgy7dSmOoEzvMEZ6z3UOjL61Annw6
JDE9FGTXReGllwTHFkGSMcEwuo9G77Z1kZnVWDwaS1bA1OGn0Jv4y5VGfpDClGT3
6s1wsB1so8bzUXZTaT4GhTVnG5cTdRdavSVY3x7pmIGs88fSJIVWpWbd5f7OgvQZ
PvyISxBus2nO2iVSC5tXoa3oZ9Z684GA4VAevXOh4T8DxEI6Fomrui9WTBZTesuh
Q0EVN2+8SZziyOPTEapkOPp8NbRXbjrlZIDRQKshK3IL2Rc8RYYS9QvZ1wx9EzCb
sgb1FNIspbNsO1nLFRqMlxWQ2MpfJs29cnIGf91xFIT5IvNQf0LNsUkgz9gJdtI+
X8X4xAt8ifQwNPTxRHOGDY+ifqHRnsdsMoGRFfVMEw1ZbhAzChrgFcS4Qvwjdg6E
8mPUPAqRnpBRW8NYJuQL4SQZI+oVgEHolFv4exmb42keCKPgeEazLGuBDR3jGnuF
m2FoOiqNoU6H0L4DpPB5yDaLorLZAPk4HfZwco8ZrLFOIG2UE5px7Bxi4q068quK
jNeblmaG3Rf0MlBMe/sDb31H7xMhq7BC71T0tJP1jPS8juD8N1d0ETUCDx0alte+
kJqRQ2JXDIgRSBo+pYgoNyN8Us86zVzeTheSTzwm/WkIExjiXHmPTXNP/WO/6kcX
qzx3+KI7upr3Y6kVpQfIHAOX2qPdGZ/ULX5eq0sGuQLmUicmWFe7WLu/1IVF2ZTH
FR56UWG4ZSf+D2bj/IZP9QxKNXIhglBoXgZ7QC6kVP2nJS5W5/sDGngT/Mw3Fy4b
3RNc6GvmmhqNKTC0OrNRUeJvCtELQfD8iMLGfHDIxAcv6KHtaI8Z6QGdxyPcoJgg
wn1sIY0PBfgJEDp39b+QsUcWUoqkx4Paqze7lYlBWW9kAlGcU7Y40y3LwowF2jqH
oXpQXJ8M06nqtIi9ZQakjqS4Ba0kbdguSc882YWYntB0WwOwhwWfKnGZW6QlO6dq
kQtc46KBOY1/ryL/2Za0A+zTTFpBjL6b7Hniji+4NmAHnMRsIoy40K/2H7sK6Icz
45ps1POflC/HBj6KdgAiBoT+E2BSuLoopL0tqIGBFhHuNfoxqCxcC2WHa4gaJc1M
k8Rf4Xk7PdI9P9M1At5fffsBZjE2+KOBzriQ9PBZeEwW4+TBCNEhgUwmCLNvgvDP
3EIuZRt4LQ7Svsbh1bJ1CLZIBLdk2qjvd2RsZUD3OQWw8IeqfukbveiDNsMp3PVr
h0nkC1Vh4W8pQHaU0NxWCEjtOlmwqsxdqZfIRfhq1XBy2nFqz1tveZpXq3y5O7Nl
tCZS5ExTRdUjtGK7nGzuZyNzOrD6buUB8/QygaxkectNCY0a+aSm6IHjKEWHd19f
Sp2Rc4UhPBwHF4digu0qdYVcX9MZ35EFsmIf6AJ5ePg+LzVwhq7Y2cIZEtt6Vcri
7rFHuYN4JQVCcEfJDEOdSERzULYRJNN+Dv+YaZ2idoUHBvCQGTpm6itC6t33z9s0
aojZkT4+/sCT6CMG7N/k0CG9PPzy0J5Iws3DIfu79pP/avJUS5+VWfwy4t4rGcZ2
64lAGHq66NGJwBdLoHTrrEpzoFcevQaOsz0+U9B7wYGW9Zq/U3JS09a1ppd/B5xT
4rYfx51ZnroBgfoEMnh6R+37zCwLGl+IuvIrEX+pbZeNtzVII5Y8CWA3wTXZO4A/
3h4IoPjszMqvmbxk/mgvOMuRemBygbV5W2plENnNRh7yEHY4/VG7LIQb4Vefc7br
xZDM6MvQQYwPQ7qccppaVT5GP+fFjfGW/Wn2Qs9eFo5rgDXArwVNSvgi0gdbZml5
Kt6VjKcsxKLOnk3DqCi1WEE3l9Slaofo4xaeTs68CtfhSWMNXKa3lzCwxlvjySbe
i61ZGUQ6Dud+5Wtq4X9EbjCZ+PVdtj2ce6zoMSx3kuDwkqWlmk6MA6PkLD7Mh/s3
ZImgIha0jXbZmZKVlLMjfCpKMp6k5SJBEFQEA42nyhwD31fD3GDM5wU0w+b1cdl/
2OmpoMwehhNo7Zg1cvolNUGibhFW64yKDIE2xvh651s=
`pragma protect end_protected
