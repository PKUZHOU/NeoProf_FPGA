`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
XYaW58K0l3Reqwg6i/bfa338QMZJ8JChr/vluuYPLbmzXqWYl8vqWWS1CTpWQcbd
SFRLxz2cVI5V46G2RNkRpq7WvAiP633S4EP+yx/2abGUJNiFXzaUHu9/sE76V/w1
I3/rVrYdwMySOkwc10WiPCHecku+eGcy5wYA+lkNWKA=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 15568), data_block
Bfl7SSCbY0gVHVYqhYVmH4cifGSIi78rYK1taQfCEUNv+3R5rcxKL+j4Md/ZSPVu
0TuyoGqK1Sjl2oGKIm38Ll7f8OQpIP3addhaxGkhfPgH0qM4lUbXue1v2MvwSwpk
yA5UGsPuFOhD7P5Rf5mnzfhyF+gZ0/v7vA/ywN6RVbyJ83t6HTkJN98yCBF5l41r
Ubg56VwCmAsLR9fI60wWRT8qsioMLoxYu2v3dixAiHtcOEG8pQey37hSvYAgNw8Q
LRZWJW24Cn+40F2fbwmR1E4eQjj8elR9dgh0np187s3YKhyGlsM92OfMb73eAvAD
CcCLdNja0MBQtk9VNbljdF+6YJeOaAN8s2FwH99JWR7mECPmU9KJZyJ95IRthazV
NEYwAmaLAkxqMZiiu79DOy57jDh7Zt9nxFwBgZ3G8bma1DnMc+Vj24E43jprMts/
2vlqsBS/Pth4uJbt/yjW7plolsGk9SSqlXDBOFHj6srLseUr+PAcnaOvJkVSQoZz
+Y6w9f/XudNoFL+AIHPz/8asSr9s0eATkGc0hPUXxCufxWO6GGEQB6nuTooK3hP/
RMhssicZ/gF3t7BdajFFVIVQjPC/w0ElJZzekjRfSgn2nOCOut/1ttdpLq+1V94u
s3+WRCkc74dZjT5zDD1acqE0WxJiUKgi0QCvvEps0n/wfkW+IpeCwR29jXLKPMYo
TiQFi2Kbn9ea4cHD2+jGxXfkszJQc4J1FV62yp9WZBPEb/GRVCMTvU2euCvz+f3R
D7P1Twa0WLPScLjUQ8MwVX3Pepv+DBsntqSLr0ouyFeeVemgK21r75POJToPO9Jm
EpHkt9aT6gl2go8070rGQfKtUfEIRTMhy/1oj+4FIe1IC1oYS/veLA0xT+D26AQX
gwd1OjbEwm503Rnvixd0k8OuQ+QIthOYV4CUhqENBxLosNwcQiDNMUXAJvqbaUqD
MRGTXClDBTG0+yZ4JgQw8bxfqWBxpQNnjMGSAtZihHmg3EMvCPMclW0giJK2xYyP
LnAKkWNn3nUFjVUNtBQgB9UJWaQON6Acm/rOpX+Hx9ah4rZw37X/PVyirfZPOKZB
vLE7Ta9MuyVRB2SC/gYgigD+wzocevMQte5GpqSORoyPvic4EDB3Rx7JkHT39G8g
BRZWRBMpVmVQ2aC6PVkuIk0gGL9cmGdCqfsE9dbRMw33dbPWQgN0lw3/BU263n3o
onYI7E/6t/gBFjDZrex636YQBD0aVck7RzMSaTLF454sctxyYM9W4A4qL7T9saOw
0cAwQbyOBTE1KxJXdt62kcYSmBtA8xjIJjj7VVASdzEQHusPPqpKHvOHP5BDS/Zk
nu1x6ZEcBuZJLqBdBAoXB/BUGQyR75p14WK9u724DLPcUeW2sfAQV1FfGEN6nhA7
Kg6RrLQRQ/LUSrx+LXCGeRwCkCevffv1t7LcVVTWVGN6zLbAsAxHJn/7QYlJZ4/f
XfUe3Q8i89sctty3+X0/EzitfLGHLUidYzQTON03Ic8ApsKQKXMy7wyl4Tdfsegp
gO5kvRY0eMhFaKoF58LISSTMAk75JRx1JP29waqJ0yuZhDxH1QA1/dmfMwK2TAfI
lGZ4NvRKusL8ktDSi7J7FJvjIg09/LIoBJrjS1tjgytLrWrm2wv7XG7RNuVCf4OP
2XRqbb9cieK8EHKCmz6Gk3ztKNminc1K5CgcOVwjqBaOAKSS3n02Mcpnw+4HFZYV
/6nhdG1PMYrJoTXciC44OLvCrF1XtvBOnP5sNRBbJodepN1+6zZJFkw4GzSGmmbe
oSp92EwV5s2r0LSHWoNWsThE+WQm6TpTu2tk/MOEOcOBJlOSrslMc3v+rY/fj1Cc
Cu1PEVNxrjXfoG+ZxwbzdQ5opyJbUMSGotld2yh143M8pCMtp/n5yQSOK3atmcV+
Oz4e4y7mQwrd9bjpSBUPSmO8QVIKV1L5/cTXL4+pHTqh0jG09SCyAm1NSY/Jb0UJ
0j7kcJnzSIZuH1Ss9RzaMrRr5+OMNnu9O3JfMGfPzUVJV8y80qG8r5dzxByw1aWS
VBbpSBGto8RQJXdBpr2TME/ZDOPWU6mMXWqnRC+IlUv29pLe+NTJwdE0070XLndq
05l7iesFA6vSTGa6lEMtwFR05Jeo8uL0EmGn4SJ72MOzLsw6uR9aLDvQ26NPz/2+
fCDW1VXOt7RoB0u7RQIQhsyirl+zdqFP0EkcN+2yR4FrEesispBxoXFkrHbzW9P3
Fc+Bk0CEOAr/xKJMwBEeP7wGisL7EZXvNjpGEX22oeGonRREfKpZkovGu3CU7OdN
dahwyWfbWAHN94pElRxNi86wwhKpaibHUb0LVFFg081npYc5JAhsaB8C46Kyarqd
McNp9LFWYJQ3p4Jq6bagil5sfeRD4X0tZ7LYWMk+q5mKfRHqUnnkDYg6yYaizZPU
6WK4+fMWKHmAeF/3CSNPTS+i4ZUBKxI1kBoteG4LCvJ5ytbu+qOWLibmtx+Bls+a
UkoShFBrrMcq2nTd4zpG84DqpKI3QjPOzs67vJ9/7IgQWrKeeYvT0lnvG2WrPoM3
YrZdOpZFR9Mau8qCanTO0KPymeNDOOiqpMmi9yS5IQqeZADAwkvtyNhSVgJV6o1U
UHLacpZVVYP74Kng8jvootMfsadgakVFBIC/3qCNVA/EP01EYi9bkJL/AaK7wy0n
SK/qvgDnXhiRyKXs9orKMoRX5dljeuvZ2v3r7QNX3yt/URUK03vFFaa7K2YLDiBQ
XhzxiEOBBW5q+97ojgniBtCEenGrhqLJjBbkgKCAJn/VawvGylapzLEIF4IRU1Jp
Ek3OJIhQhimHwceTk5TSWMqVbpU24DHlr1owvGLZOIMYEq+4zxMcHWZpBDmxlYA7
9UFxVHsdA7QGayNULeT5vAr0+2h9x5RHqQ0Sc5TMSwg/a4KHOU+YOfjj1xbrk64g
HPa9Ec4iAvWNrRaWerZ+gKk4TAaeZ8DPpUHga4YIE87P4zotE3On2g6kK2N0bXM3
sJOh050PFOkLpj7EjFtcNy+de/mHGeshpBxDPSgMXOHj6/bFpjvtXwnpzjsjC/Mw
DEGxH40TbY6OeMvq2m00oSui3w0eclWCGpFHPplp/khfsycV4hAx/z8+LXwYNFC4
RuTVH+crMH90R3Q5/0hdI+EBrjFRpkNZKnXG9Ne5MT1/9lB6p89kt7iNqappZG13
U8pqEfY9AyPcBe4d0CEuwg5GyhWK8KicsrMTMsJvfBx6RmhwCAa1EHkB91spJXiC
BBldopj6uXuhP5PzeInp250FG5Sydkf3jL1r6YS7ENeN4dzTnmpvAXQ1vIN7lKJr
l1L/44ggXhLUPi6jsHuiOU5OFJZ5/cjH75uVJSST2BRs5/r4nr9YGRelBK+hO9Vx
/QYMTsBl3vDAWjVfgszAzvmjmuvqqdRyutdetfzwJiCYUAyEA8AyahEz2eBz3Uuw
HQ+zErAfhqXHXuFYETuS9lnphznfH9M/6bu4AdVu2uui//gaYad2WjXcDpCKqydf
OllICmexT+ubTnW64qW+xbak8uN7qTkU2FO8FgscgBUhYKYA4pBuq0/c+N6qFJIF
+qDD4PtZeqzOO/+rmct8r/QPgtjRKQzN/6WXmvL/MjmlaMvxwgmyayMfU3Xj2ou6
Du9A8CbynTlSyniYKzFGquoKJWxBwizaTHXY98KalFtr2w66KyHUZ8346P+O0Qhd
UQ36HIEJR47wTxjfRBR63D7lnpSOFIBtibZcLIfEUaR++lDAFJJNIjNZhO0mTVfu
2Ps1tSrYiGSlA1wRJowmAzd9+Qx3EE3CmjRALWCrS6a+xAVrME+MpXztXKKgJhik
62xKpMDHk8aooZTFBAE1rpRa3PXMW35wGW1TEad9u8Xbu+ki46I/81ztV9Z14+2w
moW84fI2CV9BErKzglkcGSoI3OAUDHRQyZjQjEmUaDfMYx4M6KwLROhw/qEKJFAA
LNA9vXvLYX0LiW0Pgem2FTvZ79xRQ/0kMPV3cjitUIlm3nficlNhok94g/F1rgNF
TsLoG+mIkkWOpBjk2ikTs1CrbnJiAbwfgQ9JyqwjHB8QKAyORCbKx637YBYu4GNO
/s6MH9N7omvjrhvfIFJWY/I+iwZ7R1KF+8D2K4DUDai4NPiorKgULJYLc9RX0VCM
Z+iF4W9150dvmFhdwgEETl+ONkfDEiyzQU9vMddDfc4vRXtgqnrItFiJjWxz10fT
eaA1BDrOsgKP4Wgtn5E6RBuWveZa1cn76kYs6BDLGujnxZuoqQRBovqoobf8/8tt
zvnCQbdtju/Dx8YMyWfp5Y4LPfV0vPYIjB6XEBiCxbunvaaRrH7PQEcAjMit6Lfb
pdE+BzCrN3WZFxJEXZ6hU+bou6foi7/Fq/BzSvEYAiav+oeZQcl3zRpPxqUfdHJA
SN3ahiDMKz09FuznFQ1fn8rf9A1pinY+z83yEjQb19eLdpcpNh3NEwzjUm+r/CZe
k3+EO8U9HnUGeVAbce6CNkzfCebzbG8if3LbStGlDAZT87FAVFEiOpypCiuzwZAM
erU/ld9Rh5Uw6UMmE03dO3+ainBTD18/ZrxhMQPy/J+l9T2OOSe6IvAAHKsVl3p7
QSdllXKcEiNA6svjubxhGhuvoZc13EXZmpIO+OdQyNQqqilCK+X1hNJk+Eqvhp9y
o6KgN6osEMJphfrYFsBcYutrz2vuf2wGAA8TJVeMSc5iAbs7zc8fN1np4/tCr+xX
a7ajHWW/yIVYCV06fz9wLstsDqrRCU6FHLp6PBLxjXUyAJSQrsVLM+rpiD4olubM
WvOoCMIddI0vtcJe4nsJfcxr6+n3KECD8/7cdlGdbHemMY3zr/KbgFaDWcxl1xqN
mGcxHbZlGLdbyGOIpZ0HLmD/rrTbBBSollsONWq9qbt2JA9IZF0GFQIv3kQ4sjDm
C6YnrVb5IAGvUNGD/iD9Q+iefCdGKaDnuMIPfc4BoXin8Lb9lRV2/zw9r6tfTLhD
icbmJs3e/FzRh91FFUYSoYDtglstrApMc+W7g31Xlw2B5r3OoaIoEHzzsSTp5nhZ
3Svoh35MbGP1v2KIIxUL/myNmZ1DYjYL7OZSsmS+pDnfi0LThG5wUGXIEX6VTOIi
diiarY5eOOwaawl8sXJpn+ErmZBB8J8Neiyi20LPe9Oskdk25zeEyVoCEW2ARYQU
niG5Wod07CQC+QVNoUDwdZdNg6xvUxRuRMzsiTM08B57y+E42xj/ctBAGVfDCoVB
N08Bb8KvTBW+PlvnwgttH8PuxLoKZJIHk5zJ8UFW6JdAVadaL8rd+yJhx+C7W/4F
HAc7bUB4zxG3OBlubIYxGZTblatAaoMjacfJYtFgW7C5vM0tFPIEHWBQoOAEAJvC
btg6wAl9cUBc6NX64ZegIS5iCxRgIazaXZs83t3IMTKt6lvqVnqX15Q4dChFS5mX
mCmfXEhXJ3j8OcDPmBUfJ+EKIWdF9DmEQEsv5nuZniPhAmdm7YhatQ4ge4V89f/U
+3xXGFnLUSFwmZJs5ickKJtTb7O0TtD6qQgWlOW9E3dFTjIbDKLvhVm14HfOG+1e
Rmm9K11DJ4qm5Aqi40q1ndnCajD+eOaj75aRqKS6IpbkDXEDvP2XRbtw+212emad
ukK2czeMpijctIb7ov62+iEZvpFT4ggLuiPT9y3vWSlWHKFG2qDo6q7zfktc7ORO
mRNOfhJQHynAtHGB3f+EQPVwrkd6abzlJ2AiTWPAtvmmS2WeXSO7IMO6VKYk96AG
A5nf0IFzqnR1KFvDMWb39SrFbJ2q5HQl7rApzLQ3Phv7+xKVfrQYVXJ0INSGxC8o
uH7i7jqqXXsJ5BA5HzZPQmCPUzhj/CW9KPqTu/yCoOm3qHxAyhCMMwWLDQVjMLzs
W9UF27CtzTdDgOJLBoDufjmV7deHAJN7dCAWH5ZXzKcb4aA/9s9eF0y9iG2ELwY6
cm8JBfQjgoRXmCQSbXqChGGd0aQvuI9Yy3+1YtJCNk18rKDX374uRb+nrE8GIgUK
ndxBSM2K2rULwBKcmLRQkzEZfRaXusKjj7xGoGNaspYPiovmHSOxt6tipWmZAt/l
gKSo3TVFiChOiYxmzN1gV2m+ZvVQNGL6gibQ5m/2MD+Bi7VF8lU62ml9LOPVXh78
pXrO8whoHQ+Baym/jmqIOVlV6BVenxNTQZvRmEnRwOtmfrPUxAHsZQpD2LNCkI6/
cdSL27A/RKjiGduEG1i6YEoVlTf46kEUrfhfiFjBz5UreXGSlWTIkePrgDkrxi/g
zhotKFmTPMDF7kvDKR7baBO3fDrEbNEUCiiCtWR1RBEHG5Ibx+CL+5ClriyXs7g/
AvGgMgUprsfWUklwbP8GKAwhzZhqJb8YtXvpFEJ1VFj8rro9tTdFLFAwqzBsXnzZ
hQRIkb4GAqkyKQVMTglS4XiHbKCFLXc/asNZFVLlNggT+H42lj092w9BqIt7qQXg
HvaiX8XEO7Z9vriwAnnPNz/Enla9iRqcT0ooO/NR0HLNcZJK3XT9dpfhC9KBYARF
joxmUTnRrIB/vDYcYN51eX1s76alr80Q/fg5f8oCl7ywpWvlemnaYjpXI5p7S0iv
FRtYs+1zQuFZzl1OiM1zQ5SREjxLnmVjfug0o2oZrzz9KKZ1uCn3D5AFeckZLjXt
Yi/cQAlVxcXh5nxlBjtZwpRRpziZHm/7lvvaR2N9qOwsB2F0+WJlD/txFNYHm2lM
UZczf5sPUS1XjudaNacLo95JAGolcLO05y7dh+E5jWaP1CE55q0jRRmGihq3rjMs
gEQaeXTviNN3ngY6WV3CQm7Pgin2qBwOK9a666pIQtKxkyp8XfCj9JDn4Kk/H2P3
mJZya9B3/xH7WSnZzfNF8KAX0dB8HQYJGpTEsY6p/9xP4dXX9eKQxNhyNecH23yo
gkJtJ6Umok/EBUnnr6r7fx5YFlK0HbaYFUBiIK4RxYcuHP4j/pJmB4QNmjHmhp3Q
JuvPDKas0qKEZohM+dO/0v7L/gzV4Ngys5NpQVrA/JUWXaMRLPyBY30Ka9QELdSO
BMkR0BvMXzAFA+agCkQeTDQSEXlmvCoK1k+gnIq3+kB7umjI0cCRGjHkWm2ma4cU
FWMgdfcnZiPeLC9AqHTxkQf3JTnfWAZVGTAD1WxYuBTuhxkaD4r/ys7BFrhFjOzX
TRReK+1XbkJr4lwxetjP4Whhw9vBXQNrEduniPJCK93++xPb1qleVQIJlNRw7AlN
iCS1ji+Qx3XK6se7oI4WTfsq/dCjyHGMH/ff0v3k+xEaY2ft4aJAlQCWSiQW1QEB
yvRE7Z8gj6hTvhRkD9eq+Rlm5+naYuZkNJtwgIuzd22YEUt8u3n58b0zAzNZdEpo
a7mKkGmzTre7BsNpXhS5H4mxanhW13Y7pjX6hIAkl0yr5sZuJljQixEkElyD9EUw
KBaAV70wOunuVuRc3FcxzxJAB+5yG+vF6iqvzzkMziNRMXg2dfUyMN/Xjrj9CvrJ
kgxKsGz6mUqjflOiEsI2M99Yvd4Jzkj7zRXF6FEy5sSrmkkK16IgxOuyFsL8vWxe
VVoGoVC1hofybJUyGHhhMWGMWViKx/9yoM4Vglt8Ddx67eVruyL1winZTagIFPaX
/emIIQl1R8D96f2cWwLM1kjeoMIYcxnLk770iodVir3lHbFOZQjGnSca+9bKDnBE
zt19lbTafh6Z58GGTDswUFR5NTiEN3wjzo+yu91H/t8FmxdS+aYglnpbKJDe2H8W
whJ5KIDIIlfU+9fwJa6Dc2CEV90mjri91IRC85S0G0x/XG2JBboYelO2txbVgX+0
OxqdDtZhzrkNg9YtkWwOahYqYsqSzr/wtkR14kqo5RjPt3kVBOneQG7Wo0FIHyDy
YVShTXaDw/7d7hjSD7Xe2kiw/ZjosKsTZ/6NZNckm2t7hh6EwTL6Msv1Qp/tJihg
SdupABjiQnEe7MmWV+DdN9zCXpa+za/7O0PMO43QEPmuIJlqBCS6Y1PE5142bYv7
CMo0zy3J+mWzYkOfTRK64a0L0/zfiQ8ABm/hazAAIJctyL5AF9j6l6S69Hy7BvaC
dN3S63lPoTwIdpDzt3nz3aFOB5mHydU+0hKz3UEL40r7cJIkRsEHucitaEa24yxT
zR8m3JxU/DU6hZpsLMRTEQfJaWmJnuTUmiB152tSZCnOIKRJSotVstZ+vAnXF68g
GTnFIXLIjWjaoKTn9ysqJjHRQuH1nRdUyGw6dGLFVgldx5bHwx+DuiUaBwzcQ27w
KxvLFV+iY9T7xCAlR9kPQYeH/5G7G7jJ3uR9VY9RcglmcakFFnR1JK/TO91lgBak
iQRC+sqid6seCHJDmC4sQ7OyF5j7kAGuuUN4+QpYJtZ+hn07S7iwYtiw5p5cZEZU
QiL0+cGae54Kc/OgnqT75hVOmDY8MHHG1X8ZH+KhAIlLYnTMvpH2LQgL/BSWJzmE
JOgwQWibf6FJXrUa1Zrq1pzMCL8Zbi62jwGrDj5qGYKmVG+cW9URRzIpHqeP0RDT
fOLreaaFOPUfu3YzVIFrQHKlSkKYJ94+lXWGSesCjL8yJYU14a4gixSnQLn8lHdR
m/vkrGowwbK51VM7Ht3DyzN4cx7d7uu98LAL73kpMIuKgjeur+UPpzWKXEjvp7I0
hsOr/LmXk0eFyHpCySjhlDLyOMmdTQiu4HR1vtp6i0ycfx5o2CJWw/1GlBO3qtMM
4sNG73aZggnZ1tLb3C9jxcgHUK6wKGQULGMZkVoXXj4nndd3w052AIoKoAp93Q/5
VhZu1DGnX6j3tX/ABUvzuBsKiZ+CYgm4xp+uXfmLVwuKo0Iqf04o0T45xbz5rRdG
BboBQZ+9qrJjtAsXnwq39vxrNpaksB/RqFoPn2AlgWs1eFTiWWPKTbYxaU6SlAdh
N5HYYtsqfVM1ZbsTmJjFT3aXvgw99CZbutjueZVOze/tQTtSsAdnMbjeVkNEjrBM
6mKx6ESXXzusz2bkARdIDdrb5By0rHWnlXx0r748kIaljk0YmGkNjYibPwhui4+T
xDOAK2Lg67JKenf12zffiAjXi7qVa5kXr8XNC3H7vt4s5lqRz2AaXQ0hBwffkiBa
i3DW8/bgRJFGppHyKMAQEh8h1KfvuGxU6QoK01PWJmngx5raaoH5bwFssWeFVUN6
AYH2es1lke4ZKdo2ZxOl4napiAzRHNrYHY09KOAAKfkTe56b0Yz85AiAERtZWQc+
y97+hqKHdY1WPHLha1f/bMlQMS7B5/iU41M0XubIxLm2GfHbO8YE9Qvpo62oikxj
ks24fQwk39wQuUoB/dzezQJDAGPFQcb4XVBt6WyY2V81Ibm/XXSwizA0dznJvKdX
svstGCt4vpjuCZMnpwXFn59fpBy54W/kWTyGEWt13BTi4a0akSykLhfIna+PkHdn
OejrhY7yEp4MIvearnJRp6BArFDbNgO69yWFjZaPOn/BXFD7RtsuyPcZmaaGC9IO
P+jSKu0YpFulNaucg2l92K88srlLUZQ11gwetkOLNAtvegnogRGl/cnUGy890+28
ZZjImGCCNqcbi4LiES1MP4Qm++RMjxXc1IAP2UAjuveLhRSnZKEUer4Ns67azrbU
wC2WJlHqnvudaeihXWUMeCWqq8gZ3DOXXFbyOtuK5FTJUhoVx3LL0qqLyBfC7nS6
Mtj0O9RtIvo7xj/kMw9L8d2V3l9EsjuUWolk2zDvRcNQkha0zHkz0OZUq4qICreg
ZcBoFHY1lYDRxd+5NYaWHdsEOU4oeoUGKEleUnQrMxpLYgooQHMA9aM9nUh7DFs9
onun24AUcHxlRQqsSbOHVySoqcMC1sCOKjY0XDI0zpEepdZWFUenuGh+BcqdG/Vu
0HTMv3uPpmF58jbSjcx3O5T8C2oC24aY/PDa1WSM0oceQecDIeFdvRTtui0nn2fP
RvmyD+Zg4QN4EReeaXxJzObU9M/HE1+oQoZI8PUv19QXU+E/wqzbUiMJAd7EP4Pt
TnaZjMZB6xDqw4hqyFTTV40OXppj+hik6i/UrfZjM4IOo/JeWbKo5/ZK6LE7SQxt
dVQ+c0cMR7I15S61kYC+F7iyLCSwVQx9LxOa3LNOd7x/Pq6bQAFLBvbbqbc5bxYc
1CQ2vCBQEofjg589zFZQ192xXhMAEU0/TYnALrxV7N6S8+SruPiPj0luaEF463od
fiU8vfWZQqFxpQGOJ1maU2udOG3Ax+DUsNVWXO2ik4iBYDM9ZQZUh2TMdJnbVyJK
o6hICWsw4g6KpLAPMA3t1+UOYiOAa2QfYRw65giIwerq2P/OBiDIyUe4MJY8LxB2
ECsJowdK5mdSrtx2TPiWJJdzaybvNVlg8MUW4sf4lzGyeNLRG4gMhMshcHrLND8X
PyaHt5ypAgvLRTGQcx8u+/bHc2qe24sk6kk1q6QkndoX+58PqU3FX9dSrtDY2j/7
9SDcDNW/QLI4SvmB+1xbGVNQ57IjUogf9G6NKHw6V/M8TgFcjRsC2+PBK7ESPhtd
lXYMgpAar2Czw6/kl21IuDerUSToCTYa2QwO9Ssgbpss5DWo1rmq8GDKTlayEA5Q
hztH0UVS3eilPhPmbewHEVNIKp9gRP+IP9nJb1OybclL/z6tqCSPoMDWg9IwJIY8
0ML0qnk/sdZQ6qpOT0OAAbvuNJyfHS7kfj+kSW3jJkA35apdJ242HTtebmC9mTbt
T6VqQr8t8Avv5Bm3YgjjOgXKj5VFP7jYMZBolCunW2mitWfm8tChvIRIaI6ld/Gj
/7UqtuOAjiVkq6qbC/K4y2MJomAq+BTHB9NHfnS9KdBRLImOaO/0CH5oPcGsAFUW
tSOK+Paxle92ugRKZ9oZE/7CXWzxEEZSRHu98fCvEJx9hX/Uf1vSsns1UdYGkN3q
OEWSG1P+aOt9E+mECfi84GdGnVkqXt/peQ5yDHVi2dsz6NqMUH/NRURZDb500B2b
or5AOLkObjKZaemjYLEYNG0JvAIBY6zrUXhj8VIBYoYyrPbaU8yeruek5sCK7qEV
1L57CnsAGo5nZcyJwLgk5Jxl1+wTR2xshD6bsPJnjQr5T/KRN2MFNSyweE47B6IC
UxP39H5+zfI+oNMCV+rT2L0iEKhKr1KHK0NjYCm1AkjGsJ2ce8Jg0iQ+iofGDHbT
y/Bh6+MHrAjdZbOZbBVX0NrRsEMyMwlEaG6UbYvKqovCfr4raNBCE1ngajwPrYii
yHZJlvOnRKjxi+1I9zRFWKulDz+1ZbTy3whtUfP7vlWJ6TJBLMQn30+zDTF3WhZf
C/OMM+CA9Vfc/MK+B9IXybW67AhoTa8IaaM8U9eZFUMZAqioOrYCNDPGhH2eHGPv
kXTdBhuqu3S+NZJSlKAQD3PUXlAODRbzbcCy4CiCRyurhOcJ92fgJlahfDi3RvND
L6WDemnn+iYwnBeU4fESR5SG/ptOdGbglmiaXeJRTFANpN4lv8UmLK97Ou5z6PoU
FGnqV5mv3hezy9UMbhnCGGLR5XchjN2JEn2XkOuuUXgM6YAH1cde0etDlEOIp5fM
2WsiTB7lfr5dBSyjCCaVL++Z9i5fDCnkyp24AzjCZa+We+FlTULVeLhCkPBzPiGM
S9Sx8jEPJV5BcDtCz+N34fsmjp0HYCxDEFHzDd92O6kfG55eOf9+zsXt1Wl2jDqU
Ly9ggLmbwfKNvK2t2D8RU6lmh23abYiKLcb2g78HscN8KB41CDRGf9Jz2h5pY567
EBDvJnKI159b2FOxbgxfYZ7i0pHJLsPQ8xOlx1L4j6VxWrhSgyMd0R04BkKkI7Wl
F9IR0LXEWdhVtZPN40iUGkfMjU7B5Bgit9mTmmVf+KJMPUQ3D1c3uY5PCBwf1lGc
NOTX0egLkLQB/4nu9AJCnKDiC3K+QNStxlAAqUTyHHLJQ+BBgEERObfLmj0FfidR
EBwrw8ogwZdAbiemhVuO2OsPYh+Z8oZvr5XOtxW74ntZ4rQfKumIalUbF3TO/MYn
MNqX33l5ik3z/6pvedoYPnGjoAs/V360YaFCGGSg1FyeNJli5vpTyydXUsbZybqW
P40/wzY4IGxBJ9aneQwKxN6lkFZ1VRtAoNHRyhLlUAM4oI1oKrJkBNfT1Lh5GJoZ
RRXT1KPu6uJTudMv8xtWWGhKIO392Y+mIGFR/RbtiPh85H53kW8kK4bKdoxjaxd0
AjA2pHzw4U1j0XFSzCvunW/Eq2M+a2cKYHxXzavP6x9nvtpPV4Q3yi64HYSdBdZh
HFsbGSWz+GtfT9Mi4vlzrtuT8Ukq7fzw6yQ8MNX8SsGeTqqRhmCWDhkNqm4riuL1
aVQjs+2JxaDOeq97EPsV7BKeGXKUbpeOM+DdVmpJN46dtBErFK6eeFu8JIV+w+62
fVGP+9b/1/yQQpeP8x+aKwnJkS9RbTlpfezl9r69cHZjuABTCx5JMKF9Dk7rCMj9
EaVCoh4M5GZOpsK1VYBTOZ45ueb94uudsrEsaUMqRqH8twTnU0fty5159Z50NXYz
zCl8b4/iclem/z16CsXj0xy40i2HnLjQr8JdW7GyyQFxiAUjblH/AzCO+1SU24hm
456Alf6flAv8Oww9u4fse1HEVZuTcfcrpp3S5K0wco5IgbGNZqRb1abj799gefHq
FI6Ml+usql96ZFYKvz4AdrB1XA6GowXx8MyVDSeUE57UlVdAQtbWKAsvVxddRbUR
RRaDnNPXdAamUDkm5Qk3tX18bLSZeSuriZ8IXVuGYx0u5u3zRp2+70Gd92AiwiU9
XjXwdSPZFg4BkYu/dlQvNI337V+W01wLqzJ5SZhxBN1HWEJLcwz4+etK2Sa0FTSg
SWW/6BvpHDR+tapR8wgINGWCzX5S+JgT2w/jGurUpXs89fmlbJfHHhkvNkLfrhfQ
In6opRv+L1jbc/saxt3Y0EYduqAzMlAInqAES/WoYokTRFWqzE48Ob363HT+AMOf
uJd+hisWE1wUnxmwlN2qtUMmtRMYEV1nhwpAARKfLqHPR7frcluBQCy5iHbUn9q4
5Z9za2GDcWTsfFkepV+ovP0fHM4UAkerPFenF1HvVSEk9hntiQhAHeLmAyAXrL03
dUakqGqBUQQjMT11aDkc0rZlZ2guHAcgDNYr0e/4+eVBm3Lel7TDrwqm6gxknWUt
A0FALbI1CcG1GnwXx1lBaxR024cp2rTJhxqk4c9CJgYdV5wnifo3FVIs/pMZ8JBs
DGHuxl9dNzgMeHbaqyCctgM0p4DCI+to+qdEKQCZxL8XXT6TPiAENWLnkbeJyW6M
Dj5ErxEMyFwLhMAGWxk/EeaPqPV3i4UejMocjMQJG5tqe/JirQBjzLpzojl09T/1
gM1iYP6o/Hu/i1v15tkSTG3BR7VzsmNXg7zzavLamRfegjmRIfRCfeQRoiNPG0hd
lsjH+4rQewKMorvL/gqTQGkwS2Jn6NJCztpSw663zajdgwMo5uvczigR63Vns6m8
5FTaQeJJv2DflYO0zWlyklTP5IXFH2bwFr23yyv07FV3xS1L8zzKDjPgLkK7PqyJ
LlGPgvNz469vfin1z33syx5KzHnEeLEbNKUjZm6+HTEI+gNnxreZT3Cx6lwOfwMN
Xcoj2hgB5Zw/1glWSA+YxMoIcZfZ4vyH6CtqBfo4DUUboXV+QP8kera9LAxBtsjJ
8+y1GMfHRZO0+qLZQnwSOcE4GJ3NMB05qwhCCmTeaW8T2Qiu4JGBtpUyKejLIFZb
/F8oxmi1l7R6Eaj2V8WRkQ+uLQj2YwERzO1evDMI763CIxLhBrBlZVygnlalHG1c
UgzGQbQ6k7rg3f7CCVpKAC6XU9dGrvVCCfeDfwcAsUeiszzSXngv/jMe+94icFZw
/E8XvkF71wF5f993yayuVPb5l4RiX81g1uN6+N1mzJYpKSNlRPmDVjE9COD4K8Tf
J9scQloE4Oj/XJqj0j5aHdY3DUK/W3EINuzV3uv+z4Pvh5GkMq4QzTDPKgxtBq/m
T+5PdY2eFgoMx/OaJq1yO5XTK36MwhebnvnziOoI8W9y/xz6OGdJ+lXm/9VQsAok
znotP4cwWjpFtx+otlIWlbUKuM7j8XGaxPfurY2LhnH1DF4DwSVTsj1fVIjoOwR2
jGZYtuf3mjBKorqnopBrJeDgOa3akJseOYag6JfyfFqxVA7m+3n3NUcfFYId2uKk
V7ONY6sWQE1ayxcTCN5+wJq9lXdpcSSMprvLWOvW91J9OkgC7YgoupsEl10sGzVR
PQq1KCjGdHtqAThEFtYcfO6mBnNDPqDDLSiWs8eDowmhTs4IKFbvs9BaK3KRPm1V
pRgdEOt7r5P+l8boGoIPZK1nIhP2ZrMtd1k+44/hgfh/zpcK31UDdyJxMsgqOAFm
ite9BsxXh2x51UqUI+1va2W0xBM2LZjH9IpRPcNHH9VhJuvYmLApWVybcqlgshOp
USTP6t/V7VThPRqx8LrLULatua78QcU5m9q4D95JTfLfT00qoiEgdqYmnk1Mk+g3
WKO/KNP/UDDk01p8P7MSTRFNFeaiK3ZOQ7lDlYqNAuWfv2/UEyWwBv89Fc2Sqm/i
2pJMpq60SnZK2UilawBAPd1jWhsNJUeh8WIVMehgeDtaEAEYwTCym6h8AJRUiist
MSb4FddeF0wZcq063ZCQjrQdLBedz5K/w+xN4QQUJnJWVSz/kbV3wBTHVI+81aLO
eQ8BRqSMFVKHe98pGpAt31Jp9vxkKLUn8XghViqN+PkHxwwGt0E8h6fr6yK7FNLl
vZjNh3enKu+rqceQ3teVCnOplAyDMUSV3KjQLxGOd+faTLCkjRGIoX3mMSw5JIAG
7vdxRlG21+TbmgLTYvPEwa5JahRgeyfjFyi/uQKlFVV+eE/uAChbgOC8vo5z7JzY
V6IyVJernC8zc8GMKz9MOI4v8k5fdH0v4g0GCWSt9qZEFD55+uvzRCbr3heB3hSw
EyTTXXJ4gahRBOYIaImOAULI1UyXW8v79uwLkS36C71Re4oi3EsNvSaapKG1oUQS
bhqb5+tSIeQVYpc8OMaVPOkw7QvLpblR4EwwyFs2rM7YSATzlwKAcdCf+30qpvlz
FI+DvHOZwAOPoaOdD2zUMZSIGkAv8FdBXPhj1JgEM8IxWsWRdG9eDs5F+10AcnJh
MYLA62YfpKBV/CC+fhpZnqYBxxw+pNAq4YZ+mD96n5kAnMRRkbhumoS/1pkbqs5F
xhm+G6Vq6YPfQwzV00dc5Y66Y+gjz6Hek7CBW90x2VcE0KaOJBkjDW/1fdWGtYA/
Flb4rWdnolrRsa5PZIKBCB6NOHMKnH35kx6ERi9g5L3QT17EGe64+Q1kzUV6fKwU
1pOjcO2bzFa7lHC9EziUbrKHKQervOa2sGuQwiakFSGiG6Nh4SCeBqJ4eq4+kbVK
F2jIlR8JGhfu+RwGrTJRg3r4R5yeUP94PM+tMyXIFHZeIwlvJvF1LKnPgKYNZY4L
8/ygHhD+9LkM5x8KDUBXuhGIEXvTsq4ScrYara8TbDmgGTBr1dP0k6gyift9NRxu
gyTOKw3yVMATzp/uJfQQd3MGiKn3ldKkPC+br6ABjS1dLQPGhpdKGTqn+1M0kT0c
cc9DQvF4JBDfr0+e4WlpPtOszXIx9kZg3ML9j2eYt5EXn7juuJD+NClD+F6Bk2xl
cpU3iz4opzJEitA94c/9KPCCVuKtZB4VbgbL5dCxTJvylGP7LZ/3LQD3Wk1HlPc+
qEtPUPfG0FLyCCAsbbr8ASVAXdXkMmi2wTpQOW3m02KUxPFj9j12RkS4la1H9/W0
7AF+0297Gs6G366Rf47DmIceU4WJD6pWADiBfDli9vJv1FumaVh83YEySo5nVZHU
UbrUUA4etY78SsBWNlMHeyyjVwTD3cgUvN9k2gKstB/kvvPfeyG2RYPvxtGUlN8A
ZD6BkIYypG5WRdMcFUURAi8sEVwSb5PcV6PuqJg8GKqhCpGJUU3TKM+9+3Adj0EH
H+CjttkZLFd5cAhTuBQpQygOkshA+Gi43MRK0l/bY6dDcPzcp7y5qls9zMyfdu/H
Td/tzVeTzn5sKld+ydTkX4ikQ4ope8pc7Q0Y6ilRWB8eQ1rIWGszgfLxMZncYSq8
nq42WWhteJ++SsY+m3G80VS3wMf6TcUP0GNJC4qPAD7Y4s0Y/aZ93/OFZxZ2BAWd
FiKrUtR0lizV/coV6Xy8Ya1PI7fHXV/yAK5bKOS42szAmAIZVBOuowULFmnFMTm7
2Zb59b/zzo2QWZ9AVoow1kbjCF2D6WAFMrSOS92j8qx99/PKFIDU9P9XGkgSobu+
7AaO5b4q0jQHYs0LouzusvNGB6EiYJK0jQToPnKH0TWguaOiCSJxDVAPYAJWa2aI
GMDIKw7iG5eT9PVvCsDKfpanLWmpKM6jb25pmleJk6QZ2kM7vnzYy6n78zh1/KBU
sUlSdXXhk0IZEC+CnegNPZ7oFzptlanSdjiXgi6KKEbaCw93s40XrfOaej1sehF9
MLbnIc0wRZ4lCq0tPd75O7WToL+29/pl8oJeQuclZdCPr8bqRVfB3RPxryrBOk6b
C3G850uui2QTpp+vnM8Kx3Y3QputMpUWsJvzaiE6hR6HwPnIXXiCpbz9m6jaDsJw
1NqY4sXTwXCjND656r/73bo2Ojq5+X0yDiR33QYA75FS8DocO8SK9pFwzMNpFWjy
ROa3o2PwgT7CBtO+3Z3T9AoBrovZbD8JQGQd5Cv9JlEcfFDDAdRJ3owm7oRPElcL
qui4BfRHRdJkXE49NVRygT8dP/x5o1ZMBt0ixnrAcdKwK/X7K5J90D5ilfDQB/mH
BuBAtLAe/1UkM/G8Pti5QHdmi6bwGsemRsZ3f788sH/9YHZFerjTa9G+dnisG9Ws
Bmh9kfsuo5v+v8GRLeUVCHdpLrgcDNe91mTiNc/gXNNtLZBk1NWtxCqWuMK+Zt/5
qF06mkuH9VZ6E4xZ3xv99BfS6fg0n98HDoiM2OpXTsf7LMY9qPpq44FNn6w4LqTP
MPSI8QgxsTUgjLS4cSxN0j924n9yfqpZAAHvcJxfCaNBxpH6xRCl/fufvM8y7pYN
11TVGkGqBvQ2iz723HHApbzR2O4Rt6/pXzv+KJQCfSEs3/1WmQBpMiV/gjcAGVPs
00jMGv4NLoF1iq1zo0Bt9Vi1xc/LfB5omABB9y7sEsn8K1T53CYIsfnWDajNFYzT
WwxrLJu8F13CwqvIccYNk7+ndLC5n8IPXj+8C0QOO4xBzBS5KwjeWLKph9tKvRar
qBLP9XleBnuK+7gPW5d0ISSx+NdzYismaPoOr7/LvbZPjEPstNRHxlWME6fOXjUx
PouY6WmiJk84M6m/eN14zpGrN74hzMg/fmz0uqJfWNMVQlPFGAqcijhiCck5/Fiw
kdCXHD8cemzkrjjcGXQgyvufESyp/9GwW9+DaoofQ7gI0oDWizdfxKOgIeYDtxhk
zl7gLc67BkE9p2LxYIZTJNYBdvuKyrxklUT2Wd02LJjnZCrJIanWthP8CHlHn9iu
gfbxn63Q74EVJX4celjb1YjVX4Iop1WJebx5gxPhDNasypqApMNBWVkudIFEcGcH
VUjDL/YHBbvjDMKTQ14qWRL5zzMAexNwFfMP6vPktE41ligjDbbBSaHIpnGB0UUF
a2RxVXcHtUkHmk8pLGsBev1A7IEVM2sp5fMs0fAlvTmKAnO9KgcnZbidXs+9qmDm
+bvtd94sZgt//Lm7bCsfk/qM+ysO+ho26jNAnSoY/hDpwdzyuF1ZUJzq1umoQz4d
VTiTnWNJF1WfRlCZMV7DNAHWjyfoq3p1q6DZjEBre5fjQJUkoYAvMWYzISRBnJwC
KU7CflPrbQ0IaZeP7XcwZDZwHSx8FZa+sgaN3u0hHPoh5RHSLTMYZHHaXVB6gyd7
NfuT2PbOkmbJfCwkJO3AMmHKhXZw4TiP1IvvWSojWO0sZoUtfUCg41mM9krldw92
fZvgkPF+peiVtbSUy3z5iPp6luvJhnaGv33XauhaviWhOdNlo4n2HDC2PyWJvncl
e795VoRQr4DfkUHWRe6AOqEouYXvpNGkkBzuXZ1THe5c32+YcavbC6AytcrubNTG
T2kZ8Za5dpg8BXonq8MMMHzg+RNvQ1SImIjfrCqc8gFR/YACU5zF8mllLZPT2eng
wi35fyIdnGrarxenfgwc1mDqnnwxCu675GB+g6xK45yX+RRfeOQdk4ID6tHJ/8wf
IEjt/BHfsourwq288v0/Mfer5wIxWbv0/QcGw5CdGg+99UFF6LVkk48VXappIe2z
5eBYcQd8l1UQ3cxyek2FDNRfGc2tGYyHBpynX/r1r1DcDlGmPMitwOYek0osst/W
ZMtJrQevBcglA89gkYe/xoZENAF66FuBEZRQ60pa7gon5NIidUU3OaP3HrcCF0gj
tapJ2nnUk7YlgJU2SJsX8D9UT34DJy9wCcdkfQ0K0WE/UKG/ACE2gWYY+be+55nu
ZmOQw78udZ9K4i8qcIjo6j3r8/dBzQKFmVH/5yI4QJdPGfzroEVWa6G8Q9/0bcZO
LHKsG0xQnYhbNQrGs8xPv2J+I1sebg8Nk2RsT3HKD3NOawSag6aCAv9xGVNZw8cz
3Wk8uNJ8qRpPvjoNXdYAxAptseq1T7aJ9Kbm9P3V+ZjZEiIFwkuX9nubOvcHVO8Y
nYwK/qD479l9bWF7cNwFITZpEh8bPMD94y4dZF7++eqGCdrIUABvZiUBsh0a9j/V
ri7bPS0+6Ne2ABCT9Xi3vZb2xhhngBZ3DfFCjol5lEFc+Wax0OWS+2oSaussZ8Xh
F7DWwfErWACc8xKYVaWUnbasNxqyEBzOk9Q3Nc9YFHjdpmvoaOmZ0+QCxz16Rq6H
SPK1ZU0mpqfuiKpeUQaBqTxCqX7w/xkx+kTof6HDrdjM3dsKq3DaZk36jPtEHHzO
YZIl3g09jNKpQvkC2YiKrRTrkzCussSRdiT6glo/8YmCf5/QUOTSQVQYaaiZnFrt
O+uOgmQKZCv8A8mVpL1qVePCrCYCPS5b/43shVZz4bcsYR2pL+6GJFo7wuUhZIvL
cw3RphC0KUa/BYu8/VB5XDKDVmxweNmNbuvAhjIM588CKxnw96qw1vBgmF72yF7V
X9RsZCrQjuwDemViDeX0a2gW/PIquL9IU8rI0kzYxYN43SRjYR8g2d38YuxdyuYU
xxHyt5izx4u+BSCMfC4EGmzzjHETyfOPW8MjOhI5LRFAlwsEfejYcFCoDdkbJGHh
Z3IKqYIzz8J3ehnfolMffn8KisBswQYQWA8Yf4M9GUoyPr0rryzUTYH8olVFHjJX
sgvWm9Sjmj8cEXgWBs4jicLsnAkYb6Fdl8pN3vGaAhtmX5Vu9V9S3FNVi0qk/YYq
GcH5hEFkfPU248LHainHpk4+bI5IPW3T5KiF68zIY0wwpOHbKZnctHW/AyGzq+BT
RTqxSuHJ+LhpD2WPnciVg8dyGTfKahMSMiBUMP1qNrCsLa3Ue7fU014A/gdLhMOG
NBbtjkuaadeDuQB791zUsUq9YGbJVyzQ4KsnvBRJ/boe3cUZW9LHI1GW+x/nx+71
EWRYI4C0Pa09oNvFm8Eip/QQOYIJ4GnPtwMlsTzbeSZ9Z4RFd7SJJNFCWNvlTaM+
I/GwRsK4krxup9oJRwtuc8Bv/qL0YPcF2MuZ5nyGfRn+S8MJBNlQxTdNT5tVeieg
9LMwy6+oanhkLEvsK/Y2aRDo6m3Mci1bvK4Pk23eQxcqXTgjwLEnsLF7FFUMHxgc
ydH3VpCjWhBc52DhBnyifaNNhO+DoI/DRlMEYORv0Jww3vsSQbEGWmtoEHu+h83f
CZNDwEaVHiVVJ6LaRLULSPuIz50p28JPNrYu4LVF3/TmAOKeGQfQtSR8rQBIyP8u
/WpoYnLHgi2yjqGyZp+U4Vrs6vuyLfbLxIO9sfECcFOKQISDQgh61Iy9tAJnH/7e
lvY0hTOLrf95w8IVh+u3c5BIx0M+zJN3MVd3P3nB8NwbmaMppqGj+uFB5xgFSIqV
vs9q0HDUEa8TGuoS6xcc8S75ZYZ6ut2zaIGgVfz+K2vTwBm0RtKkUu97h96o6lC4
beTsSG7vK5xGMyL5pAqceGhF1Z7oUpSh+h+k9eVgWR1t4KjwsRGzURQT1xiwngqJ
VJqYZDWlotB+WdqZiGt+WvUuTHFV44ZB03KGTSvzbAPmdA4d0nDFalzZe3T1qyW8
JLOe4TM42TDYFBNb7GouYZBgFtg8GCNXIeMMdrKITy0GT4WYD6enR4BuVEICiyX8
tUeuvGQ0Q5vbcLi8lSkZZaKYBVMk6WHJ9HwWteVw0TX7fIrjw92Yuc+DArFFyhUm
/ndQxNhnMl6XZYuUrJ91g4rfUrX6uQGBRpd7Y8YI26IAX/EUk5eJUbtDPkBtYHBU
BRrVitDc0UPsuN7Yb/KhCMt0TTJmI679VlwftDfuC8YbEqi2q5cxI532ErbFFdC2
8mCfYuhHINazIr2KcAjc8aHg18Mm+RjHWJyE6GDUVbfyEVpyU+tLYIuuQjuqVfqx
9rjmuj1+XV1xXdh1Z6mO+IApMl+zruKlIws4knhVJSV06LCNk3mEeFaG+Jc2B/i2
oiFZE3lkeWV1Ek1EnJdYxAfNlMWO2i74yN0/XVFu3Nm+zQiLtIo2yOUgQIyobucB
d4QX5IGbtbZUheBQ1vRg/MdEH8niuP7s7/qw77L8Tz0nYjEyjTZMDuFEajEzOIwL
6GbHpZ9QIvUeW+cpXkajQBvqNEXd8VF12pY5GD/RRI0nFSmaCga/B0cV+qIb8T06
TNQHjR9oqPKkBuvVb+H1pg==
`pragma protect end_protected
