// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
QfURIXO39VgVV3zXLb+B0Ha05bWpx1XYO/2uQbahYA1h1mAGKE6cCyjpdvH6pVbk
0qsC+ckoGoEPqvRQ/tUgi4n271i942isGs6+8am50c0WHdVxitHFuCAch8kSDHOa
A8JO/lfJs8Crr8BC8LHjoxr4bGjLrx5C6xKAdbcyfRk=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 67280 )
`pragma protect data_block
wtPK6dXcK4DNpEF8O2emTis6mmhT+/xZov+T3NerwpG1L7ysoBb2dJhL3bMZwu6+
5QraghgVXfllDrH04ai72rNxmWHDGnuDjWWqnJ9aKk20EweCTyPwdwYGVcTu1p5s
bOShZ9I5WwWa30tPoXRgHyFODEwFRe2nrGN7yFP1RySvuAhLiRSIsmpVO8QWiwJT
K6BXb54NZ+7X9iEEzLLAlTuTwPy0rK2bL2/dW9OAjk55uunV1//KMb/fhy0C7G5/
cj0bgSzP98g0MLH0yzgsrkJ/XJByf8tJyEZXRpHHkI9yoPxI4w/jcR3MQTJF7cCH
6dtNZOn5iLLFBZFPEM9/d0MkuL8gO2xUU2sx3PTqdhwAgr6kHNSEI1I5ceJY0342
o3D0OVRnqrQg5fNeaXV6i5I7axCYUURD61OZhNeaYp3x0ONg6Qz7x5KiTY+NBZ0D
xgo4jaSwSXobztavLAHfYX1IYbQ28RYBkRrYAm2UfvVbDPCxEXiAIzGiMLmNZBov
8A8fPBW8DcydSz72R4uI3KaIZkF+RBViKKPKuRQ8zPKUqocB8+GJ89K/TUmW+Lwj
Zi1Y8SRyWR4NzowR2D3InKp5u16dFGTh8Qbssgxt/EorLXmS/FN1m4uJPF2OxgRR
pLsgBvIzpgdjWWAQzCyv6tB8gO1mAk0NtnxzC+HkJXlSaseDMVdEhB/71JNZOJfT
tNdqShREH6XVZHmmYFcUSnRZzeMGVoBpUQUXzUYwyCwHXGYUUfX3E/2c9QziYQMU
S0CeflUniDkK8GvYLLVl+fCYilVUC9C9tBhAz92wjW/qbG1r/+hbHIZYzVtxyKHB
AWkHXEjKJ6qTQDbqNUlw9e8Mb3Y20y0I/8fTShuMFhJ8hkcEJFC2/8NZEcU+uS8f
DjlFom4KgE/d7hpOlQInITTbO0HzGzqZTbI+7hbQKvjo5wBWBlEzT9egR3TQ6i0d
vO1ilPjHXsT3D6Hs44lc08YoHodsuLphYZ6QPsVhnbcN/9bRTvqqvyfXFepNJiE/
R/X0yzwv2x7OPT2Fu5SyKzw2tZYbmU8NF1b0knYXwavcjAwOXMX4IF6d8UtdJT2N
L+FBo/gV7aq78FHZi9B6y8EJ5w5T9V666nMkxRq6y9qkdvK3MuEZyAwIj+E0itcz
GygTw4Lq+oVX2DjdlaxJWSvgiqjRdVPc527hhorvZnz5X4GJCtkmjL7dz8/psT0U
0v1TZN84sKzW69XiCrc+YANOVCgO8FauA3cDIKz4tSwtZJDnkgqfK7dyRXf9jgia
rFzssJ3HKqYP82ocRfk260VhQMvbrUbJZ9vRK5r6fSe1PGnJEsGjsP87G5YO6/6a
ATcxrQbwlBht80YTklU5AgRu6MleFHOOF6B5Fvp7Ugx+LqwA0zrbJ0UO7l4MfDp4
czT00VZWjQF9dKBW42YlRvAEQJEbpvwLxV6QOmEQw4EvliEFAIOG6MtjewCMr3ou
2UHswhuladdUaZGnr3Loi0QAhaBZIHgkkK0VsjXyyfo3FsnOpcoLstcTbRc89Vhm
AJlwXdM84gSnJM6IBr5GCJnydGRqD2jo9g5+GXfQvaxMCckcBznoglAVeQzfutIE
wtWvlWVyBVSSirSNoeRVzV2lZhz0L77Hy8vWsgjKeHn4/sChQ5CV8mM39qDyP/dE
Etm1afg0BPwus5Tm1BIhFEhFh1HUhtf3Mk3Alpw9dtUFKu18Afkf6xvv8c26A4aT
yBluY08a/eiLl1+gJRzNCbDE79Cc/MxeCUbNjyuJPnXjHjqGRqaJM6I/inUacfv5
j9xcX2GD1PPnXQpq3q8cZjKpXqPe5mMyXjNT7BisZbh+kH+oanR2ojNILSSIO67c
QVzkLlCt365X3qWfFaRKnrv7eRdbX35LoBnyrwa+UCBz15h2brTP0Sqbqk7BL6RV
Sqp+N+XZ+clTRVvBsWitOVeM0B7h5w6axq9pC2oAwjsTBqR5L8nSKpT+MHCEef5K
DHOc0o0iCrnURu+bUqH3tdkyPZFPC8oHXVJyfSnR46Gb8s05Sbz7J0aPNHVD113k
5EP/eYGu6qdRCiZnZeuwDrkSuXIxuca8en+XYQMTG6VS0FVi0+SFmB6HkbJPmtfi
2Ncx10+72SxYyyHF2zNFncxnz772saJNS9EcXek8CZahLr/wZdIyhAEkzukoxLI3
YzqYhOxdQGcRXWMsnQjVA0R7lHJNhabst9R/xNrcMbRx9Zo8NonErSnGS+mUXE/7
85qz4+OTXmQpylJx9+OwxlFTQVcmgOjLf0nbqwHaUT7YKe3Oik0bwHpFaLWSBYwS
60RP+AeFrCwvThqucbAmROqi/8SSgKyFk5OuDqmuzOZBtwsikYv0rQVTRpuh0sVM
8WoDzG8sUeBORMBSoIZOt1YSUHjwXNGLddpfX6pt0lWSDFXu9X9o3jAad6NQQTW2
LradaevfZTnVln2fbkbaHAojjSVrOPOWwhQK9hY3CE6g0Ttv54LnPfv4Jntql3Fg
/gV9lBZTKfiwvn/thwm/Cq1vST80E9mfyFTHv8TAfv7FAYZApbGo1H9m6Dq5qToT
0ffxf+xpCuk8QKWkn3H1tv2hr/exsD+3PSFrhwqTXfdnO8WPlKn1VaHrkZYyMduo
QOHhBr0954jokzl6/mSk3tfBAxQwUhZlQNFtuV7n3/0FwaZuzwx/PvYGqeKKysgE
voh4r2oXDRc4M5od3K2+9nFzwA/VuVmdC/pQuWugjxx6OetdWfJoxjhVhkthnNt3
WoAbu92Ju2oA07pYH+c8G+cfj9ps+AmVys4w7T60MG1u3PXF7ibgJSAMBXLBUCeo
XxcQrR+elM1otGuQ8ZdpNBPGbuODV7+EYPlbMX1Z/x0kaND5xyN66FX4WYAlAq01
AeCJJcyuXw1FXTtryCeVxHjoCXbi+WKgzj/OifMlpVbgS3RnsojkyVHLauiW9Q8L
JRb5WpyHAnXD4vgOXR+EHyTkAy0eN06wT88ej67ZsGnheAllAn/RMkbIznJHE8LM
xm8auiWPS/DB8QOV98ChPCGC96kWSUp/JKRSllMiaAKLqDEInZRRekPATQG8YY8q
p4WISD63dgbVNtJegS9DocKbRPWnYBciwErIvh0m+n8FDvPIkMbDgkbfdciOZgPn
iGcMYgwrU9QglZ1uPXkM6FxNSrLNq/4fBc9+Obu3CpEK4GvbQ5eWrRAdE9lOmxJR
s0i+tIWcaYX5wGlBRg7gohib7i41ZQXLDYHn7Ow7qnxCn6olCeIpumQB/A5NhsMq
p6lMb5r6tDYnGbymM/7xF4nXIlNSLCh83pf/f2J5hy8LZRJt5vX8npW3uQjW1GHq
djd/sVj2qw8xY2JQN8ZuYNVDT2XlMMULlF4d9KJNni+7O2lQR1ZRhMUiiWHfqPXS
gjHWF6TXS9Nic/l6DLUrNf8WW0chEGaYUB+PDsq6jfUXWsAS8JkgnGwZ9I47g0OV
D2oGQ785bfeDTA0JldSGvAbaocXhwQ5KjC4ECa6UWWA2LlB8dYB1znVkgEEVgBJ0
cd2e07BxyIAkHIJvjtSsfqn5xuPkvnHoIgX4RmiW7KPNMkvZbJuIEvN6A7bNK7js
trJfzsP2o97vutwxyq53ZMT06HN8SZ4RchTeSlyF64E+Myq0E6Rt8VIlOqIz0j2F
7zZ10mzCNxjQ2Ab6w0Yst9jzMXLRVlzWtTLLXWyN47hphyE0WlkeMRxLEdM2b4jP
m1UKHYxt2z9/JGrhFWQhnvHTGD+oCdHuC8Nkr/C+lJ/bRwDwwSXpE5SGZfy2L1t2
1AhUX2TUrFLPh41xal8tzRIj/rlou+Uq1/839K8r2ipYEjrum0BlscOd83tuBMt6
J5FIXwENTC7x15t3MD8XYijvq5IxDpXZRnc3DTMWfD3JpHtpzMhCRcel+iY5aDe4
IJ/A8Nw2zVCNO/3/Lz191vOK1TP7iQWQztaP7lP7KxWCXeWUl/Mjh1mXjV2Exsfd
DSNgOQdLJvCTBsZ46Q54Q+eUjy274XUmapisC5QzcDc+0FlbswKlHZkBg0yrHON6
QveHLR2xQVGu/MFLTFWIBV/G5KUgHdM/0lgEOjvvK4zJC6bbaaUYJdwVbUf5iObr
8FR0AjROUGOIEy8/M2IRoT3Mq89xrTooA8uRZAuSaf/xjWzwvRmuaGQbQSiNRfqu
ueGR6Xl1z8CWe3J/E02qbVURDdLq7wxFUHaprSJsWLOB0IgOBnvdz8B4j1UbDd3g
1iHu2SC4Ns0qL67WY5Hsc1+xs7nkdYE320NEuEnhvaj+153TvzX4TNLo3oH2nHQ3
CazHuP7wxrVzBBz00YImJDNtZSLhj3X2NTU/pEaNJpctP8Cbt7sKN+xXHO1vMqEr
wJZMVpPqIVe95vHdJCYdL3j7H1MyjvOpjHiBSVLX+2cXnasC6lk6dqvHwwSV61B8
pOSwN4M2l4wtbibblY9JdjagY50wJlyjhNga9wv+86zkFaX8y/cBb6w2fB5LU4N6
b083Qz2VN3mUXAUevy498N5zcMio1iseIhOoxBMU3ML76iYlEAtzGUhVyUZBtYFL
7jlMSbTGCC2sIqXi3KbqscwMHEB6w4YS7OSpFNGGmfDDP5nT79GfuUD7jKf4zJsP
uHI3Ugof4U1NsaKUO741VmCsxNYdKO8Eqoirb1IRJ+wuWlhXM96oZsxqr0sRsfSR
ihCM143DJQO1KWSZ9ub06Xq/n6bSj22zTUsFGrjoa9ILyzbrM7YbqLe3XcJ9raAr
eDb856rcHSYiTcg+dbVyPUBCXbpqzYo9pXiG2IXgsX52EEPoPB5Hc0YbLBRFSLrq
UBq4PHYTmGGKcdXp9VhXTU2IgthGHJScQaeqxJIeMf/sCY4f3D17xNSytZCZsDu0
5juODzf1BkCNKQvrQSwy817eFp0BO4J5bhxah0rUH1pLwDllkSG9kq+5OWJcEkTo
N0oLJvs0kAzM2bOGzyDBxQ9wNx/uy/6CY98+Bp342K2dAYVkF6emKdOHoJuVNafE
t6fFCYG7udpWiHNVZz0pJMTgVKExcnRTKo1FvhB9ExdMcrruMHQusOg033L7i4wU
7YUIO2Ecc4AkJkzx3uXwxUGqz05gNUPgEP+TGMFs7tP457ypGgAc2y1fKWecSEYv
NC06iiFFy4HISi5KqwV8JM5UNXzMIX0U440cHqPzGqH1tEz96gRaJwAcxLgMHe8h
MXAbzGmwVIUN+REqeTwaSc7fBByZFwZiydMVNt+CLelz68CPPWRmnFezp4+62D/Z
m0Wk02tNwbeZmchfsk4gPxy2HQVXxJ3X2ndTremgSqhWF6iNK621S1UndQvvWV9J
Qt/TUv4tYm1O64VCOWmhAD/NoYEZC4+oHCCHU6gDRRHEEHMCxQjC1TnvkrUQ2vVE
K/4/BWLEP3GRwSpANDP6BMiuwP3PAQT0fyIxCLIVONRDoeaP+jCHeBohrwWrcCan
EQHscd9lUOvQsO13dOukq/V2nn7J5GnwOwHw+jKBaZaKDm6DSC02+eQaS5SG8js0
m0dPC2ppYOZ1idOqFyM1BZ92pRnW0JVrBgvN2iJKEL35yt7APGTEp3pxGkFkpDsI
QXrx7qVfFit888I5m9zG5ayaJoOWM1jQOHq8MILFm8cS9ibcRdGobtgJM/7fxcwG
xTuxP7Yj6IazPqmdcw/QOEjzA8tSmAwgH2+u+M8hGB3kbafbDQtiFMmk9+jS7r36
LxVycxv/ChxEHLTKd8MuVYyBmsWg93///tELflK1RiS3xOcVtF5/u8uxTmXdHpcG
xqyU6+Z23Yqb5Jfh9FmbO2KAOSWOkGy2KJ3enUUSXqvJwzGuNd1s/Ysc3uCAdNjc
DV+PWB5UgONm6bI+9RfUxwNpCU+LHl+66in22qd4SPddECuuVl+6xwmcbQD7IiE1
BkEbn3p1NieqHdj573K/y3pNP1gFbqe2PINwCoamOEJ9ZLZPa+ZTUVgo2jRL4ysQ
vuLB7OwdA7TQxRkKp8O8qUPKh2W5NMFygwroBklFn2q3DwfejyJ46OmMILiiZW63
TKMfnMBaNoi5l4xsjOT9Rjrlz9SqXv8krFHfSpwvf3EDwA0JzW9V+EzctR7JYn8R
uTCT6ilNkf0gz8x0pBecRYcUSesR5zm4qogB6s9slL872H0igl1gzxJypTrhvRoO
X+0sfu1MNeJHURMi/I4B4hbaf525qBYaF0YtVB0zOHgHa9dQMrP2MyDPDgbdYASi
DCMwyRxGM2UCNu6Pu06Sb6QKki9EU8ljQ/TgF7N7M9lo87Nw0yN93mxTQL/dA8wW
YjVs6U0vH0iVWnERuHL9RiijRqCFBgLMKIjIiE2aAVtXtl1DzLkfqPuRJCw7krQc
hVkFCtjYRq/I9qlYLlwrtOEqjSRIZYblriIh2NtLPlJPnsVHXU4fR+j8E0/xjWkR
MJCCtCuyhhYo0ugmlZS0+i3llqGJDEzYZe5X1lgG1ssGHraMYAN6J+ZeBC6pJVYe
rJkmT6kAixtZA4TcUtwvxu/8Fo2FQtkh4ZZZB2XjlAcg8VQ1N8ebaKz9exsQwLqy
EapWfcKHT4On2vkz1dqZJBE5/IXeKVLwbe1Ih/qEOFyXqCCMoWvmaAG810zkrP9z
v46ktV1GH26/YIDfOWDAaKD69s1JRC+8AJvp0sDKBDP8RNYHoTjLZdQ/FsHJR9Eu
0mu87yNOkoUol63/gMcI6uEF2V6qRyoDO36cNx5zFLu60Ihrczi3wW0NAltuiOUt
cuOc6DMp6y0nKt3HXOnXc0dgbUx/FzlL3LImbPuI5vlA/dZMdZSQNpfDuAYqWxWe
p9XAbvy1fJc+JwA9Tsm/K8p9VuXLY2IfVUwTjACbRZL5Fm3XpiNKW0fsUvzVghvl
O425qdPqFO0gxNj8+V4YlK6FBPiXGir62FEE8ClU7pCDIkBJUIt3fN5l5yr7uL6A
i3plJJlLSiZ+OI6BPPjl8g58dg8tGEhvYUF33S1RcLshiUah1STW5q2eUIyK4E9S
kEpLtpspqVgHX0nmK2Vsd6kTKmO6r3Bs+fZx/mvxaoTp46Tu7Rny4gr1zGBTaWQH
kG6C0ZMDvM62C/S3mz7L7eraqjz1vPx0XbquVuV3D/40FH9DWZXGLKasiGWY31UR
5KNG2poLAumlriA6BLSsUu0go5OSfJvB5NGZzJ7Htv5amn697IrwhJUHqzNthXaK
S7x3H0nWO63iWKGLJluQaLIse/Mjavva+CxWBnGdoCMYjCZvyhFXD1XkOW9vxWco
ZmF9qbJ+nucBykvBivChNe3nEIVrRtMYH1FkJ7vZPCekt1cFTmCjGG7sLLI/z5TS
NmG7lSLMC437eHY1UXd60V/tiu6ZZ/PgyG5xnEkixrTWrD1xwLFateTsNmK4A5/D
nnQdI6PxXNxqyVYLt7+WTClv9nvu3l4LBfHd77qqTIu4AWNLHp92Df9mSOt/wTSm
We3QXht+mir/+tyIQ7vF4O3VZe7QeE2exzahUndaI3Khk8A4JGUsZRsEB51oJKTc
D1l986hC30CC6+N/cVOvEThiPF8BnhozXtjaNVsLDtuOE2OSvcVl0cwvA9ee+553
OfSbj5hS+aSleGIs6u/2r+gZYWtckhu5V+wjtN8O66N5Jgwwob1b4qp788zaLHOe
cPWU0ZtFANdYsytyXpGIRVgqzDLjiJwwh7fuq460Wym2YJ1ig0IkAJYfzVcgx24s
BqjrYm2CIGQ2jAhYLVHljgFyZ98gY5boQPYJbRg1HB2Z4QZck92bVNozJWprCRI9
oOziYWxHWZY9qlwvOl81LBs6EbzX3a7bh5QtGtna8b2q8E6kBDM+VQ9/OumJ85Ky
l0OLpcXVbvJsk00GroXnzvualYGrh4gJTyVtDaTeGC6BlfiOmXh4X6CwoeqoEwu7
ay0jBTCOJrnifB0fTo4JcfgsW/QA0uEz99ZP0NnEIibYoeyyEq9bJJW8KbhJ2Ux+
//y/sz6V32jTWAKRLYgiF4xCDTSYkJD7OeASSrq3chueYFftwSMPe4GFYhTGGMpC
EdbjX+Av+VDSqG7VsrwpY8N5hmSMsgwjCt8+Cczb/kSHf7A36+3NWs61fE1m/y6Y
Nmzj2qbxD6Ir8ZmRs/ejQz1NE+NQGdPhF1S4aZzIm4qKN4K4zTlFPbeFCAc22CIW
T2HcXdAqIDDaeLnGQ7U1xVu8n4j0ITb7ugUQoeK8mkJ1KTGTVcLcYNDfOD0t8Ejz
UTLB82Pywe6lxo2xes0uEX8SQVq61CwDmgH/b8lori7BFEz8RP6+iY6KgNFi89q8
NTuRfg/wsgcrnJCMfMKoJD0RcVUJF5sVujNv7D8/lXFG88AboqoPQOEKJnUWiV4v
v9SwmPhVZf1nZa+YU9Q/vQ0vAntZ6GDq5rNmMBuFutQ054LbYLGWYig4LKm6Tgd/
szc3nqIym5DdXso57PBx+zA8JhVYQYacP+AEwrnsCiR9xzsg+2IC51S1La5ladTP
laVUp0eVOTx1Xxe8JFN5VaQ+meZXyvbkMS5dko/KUlcLV0k4mJHtS/pWdO5B/c0K
GeGbTtyckAdLl4I4KrWYUaZnVBTGJhKdtyhAHMLoUJYEx+O01xsGGa47JM/2G4IJ
16psj5hrhbD0FnTBNHhGg21HLYnawye+Y2oIsJgALrntMb6vJq1vFLcinNBCPWVA
EkF/XqqNu8gA9JVoTsqUvHQlkLdSGJN7spQoA9qWjKUNr8j5IVbC6iagkrcTVUF3
v1gYO5jr/c8zHcKce7g2+bZ+aF3ta1okUqF9reZlqmn2Ccm6Z81cdU1UqgqZX16C
1xTrqbyq8tvSrx8uv5eHLSlyZlIzN/y/Asyjd6D25c5XtSG2r//PUsyPA+A/QTTF
FLjuyemNMfoTsRpWB5O2XJpxZ+Z8GopFRLqZ8IXQIc+K4uylm/c63amnXcWTaIpX
V/VS5FgDHzYOy+1ZHrV3WyZCHq9NTQ3Cjj96lUvDa22bFLu8DXV2it+x5O/yN6G7
YMGrJKuVjDiWtUqn/4kPrpR+wgkIwgimoNtUvM10+GsQk89ZiGPmRkQwxdgwRNm2
TclU+ShvF3Kfv62zJ+HSP6mvbQI0WqSh20dY586F3fHZ06QSSJVGsTNnTjf1+MC5
cmxUJvu8ycmHlt+CD6tdtVucOQ4DXadCZFkvaPsIsByxHGanfcM1Eii8/J/OJeV5
wMT2S+JZaIVE/2pTZXHzuoitTQMDk+SIm6KTS/OxZPDRtuE9TNFmQd38E+khcAik
tqs90TZLTjoR23fe9Rt+t6gbDsaxFSVjDdgWYlyBB8K1VUPMbCLpK0nue4PBEZ4q
XRHeel7Hqxf74+abN2Srj3bGk42Tkvayag7T0XGiZzPKNCr9xmlTN4UJ6eK5n0Kf
/pXjhbOUwwMBP5qh9dNDRFMzRmipyF7OO9Efr+BNV1fy30MmzuxphhP7BQbjeaMl
vjqtCl4ypJL1pYlbT6sPvZSkgCPveeX79qdDx9bA5skmYl2HRECcl/EozRcNpNje
X6x0jbvImToQqgts4xs8C3PBGrv5baiH/J4TXCa2BAERuLjQ7YBkn5Vlg1vE/tT/
DtaiNeHOgY+ibuoJTZI+xrGI8Lbshj5xssxkWt0n044HveQRxehtQWp9mhiX3LfQ
ruTS5cVCOG8Wxg7QsnaoQ8/c2VHOBmFm+N3Acf3iskVLCeif2ZWiMWsfhBl0m+Yu
/Q31c3//ZRPViPhg2VWcFAzBimee//LZTDFsOo3x5KKLlvAiAqUGik2xdSW5b/cQ
3yefIMo3Bl06lonn7SIQAjtLoIfumu3I4THLtJ8y3vufmRH/3KCm6xg5uE0KvrfA
xD39pH9xNBodNP06iOjiAUuJhGJmrlOXjH75+s86CJa/Wy0tnMoNaNfpf0pViwPD
yEHQQ4x+Rd0LmaOnxi8BycadlJnFXtyS1YswSLXBak3Ib98+vw0s9utpYvEkUD0u
NFM64K/TNSJZXKdYjL2OJuPLMF/VwQSqURcoRi7b6armIyJwlOhHrGkQl6kU09Ts
ItvfgVGODKVPj67wLewvMWYKO7MmgGGMa5l8Xm4Da0edaLuUYOaBU5WZiv0swAKp
W/c+7h5wO1d3M1PJDkFVIwthJtumJTXJi+bSunfuOIJpvR3AYEbakMGDWjcH+5at
edidzxBdmblsivcRLndLP1dPKOfNfFpgjInroLI7+RZ8Qzu1wi3ny0Mryq5lS4J0
/8/eTfL9Pv4yGjXnoPqE1+9Ng59lbqKOj4Z5JKnGq1l41JsJQEFw9LDeFGQlT+6E
RISCvsNJeKHO03xiM2UTKIcRuOWAFbkxfaogulQIohHU0RmjVKMmNHa5I2/uQrwC
+R12mLtis1YTjdsQmhO2sAJnVmAMIJYJy6Iz9GaNdrManZbj9hO0wBnfiQFQjuqj
dqNw9L/AX8V2V8Ofsxyr5hho2V8YAcuFIu1PI+qH45S3px6gHJGr44FQ3uYZd5wB
aRsh9GJuHY4BIuPgTmZETPUwK1q95ZoqFo052TRE/+LfH4hhF+OdJ2GENh4s7kSy
kwSr+yaQigSIdxZjVNoCCcrHYsVf8bNHpFn30n+4IVh1oLH3v120rgVpGC0EkqRq
+VHAXnuOEwDW62f3C7VQIZhqpGi0++1EfQ+NqSbxcjpQr75OBBUwE+r8rTGde/P/
wD1u3HWG1FL9byHnGOMDCpviG0VrjrVvJcpsp0+MMCYjNFabFPtDWG5Btx2/eB2j
Q9G1u1XjeeNBJejU1jICIs05MQExRwR4jfXmlskmcWeVmVLCt1jsBde+h890c4bx
yk/vTXFoOjjue3r7LEubtPcWhJtGZMdjXNm4KwVinv9u4w2krb9e2PKZRdeZAL+8
inrcgFwMjZMKIhC31vFxnBteUNPXcYDwiVCZO4i0DcEIOP7AcnBFqKehZvta6eMr
syHrN3HzMIz8b76qqkoqeT177IYmOclEDSng5bhjXrpLFMWMSdNuwDBh8M47vCa8
SsIO9xZBwAEW8znka33MnZiTpIMBft7rTAickj7rpdNsQZYT+6IQm4+JAKXwXizb
omD0Aaw/b8X8hTSMzBoSzR8dy/0SI17qRMVQnGi/mA840g9wYEY6tb8pskwjZRkp
7gE2/ImseEmtGjXPNlZZ2hT0pqFNXgcm7K/wB/BEgf6JElCmO+N2xf2g81SvGgh1
bgTyeUMIg3yXui3NVLjLygfT7GDzCFVDfM5WwT1zzGAGBtVfYRfsY2qyyzk/DReL
RiXZu1BNm8OEa2y/UO4Q7GXF2lezfcZt2d1LBS6akt5E9QhvJiu8MCqXl+Xr5Cro
WdH/1QLaXgp+nSeAHhjbPneypzItweulgtN3rBI45v6+GV3VDAvmyThHcJPLsQnt
arj+wzhhHe+k/Qlznu77CJbNV5+SSE+AuISQB+AkPBTIabfpSYyE+c7Kc4mANfwk
W42ecBgQLTEdtj80eSr2P+aUXbECNmcwIuNnd23P9ftKOhb/Vvh8mDX3GtMduV9y
IkcUkkjvz+1IwqXECewBvk4n5jYQzHQBxLt2hCcpppeaG+4tZKICk4Flowor4qKb
gYn90+GqcZBw0BS7XVgFcQ9fB8HnKiqXbg9osGXhs6blt72qzPYRExBY8fWsJhFn
Fj6E13Qw/h6Tmt9+OrRoUxEDS29PFJNmTlDI58RK/kobJXO9cYTjUyj7v2RxjNz9
GseQ8S+HjkF/4oTrQxTatKKl/bQZMS7UC/99IzGQb9olcjeIoa+yX4P1q5g5HbAs
BeHe2VEDs0yesCSQz7u3fsd9XiHZowTwRtRAvV+uA4nsunP2RV3LnkbHk/MENU8C
c37D1eX3J4OFqaDgB0Cfc/tCQVLQLv1LOOnwRWzgu/0/a+txrj17NZ5IYLqp4pxd
MHzrssm6MyxmKWlHHgV5RIrvR1p5waOEIL0b3Ia3Sij4mIfert8GkQWhaEnibiEp
ptN9E1Vto/VDV67sEi73XcPbMcIYy1BswXRMxmxpmW8iVlnXL1833W4xKDGAW9jv
pR1Hk5A4xKDGdJt60MCxcU1lPs/7wKhuuJCBD0jpKGdACCafiJZHe22/HH2oLFwV
7+9Q6yCj4OEBtng0mj+BmghzEKv80cmIbjH4t0rCEOLuxKmJkg4k1kG/+uYOzYTU
pWkW5gDpgEjPmsOes/jtZuwsZlvMSoJBspoDH70vxF49glZWYxTintPRFOI37K5m
pQ8hpxiuWf/ri58YXrdC3jMdPKOHuELISPXf4vECZf6StFDgczhdSuRtYKUbKPU1
djAXGpokctxd0Zf8xBy9pe7O6Ohqz+xmuPOG5jVn14cEH3C4ixoy1Am+pmQHIngK
aAhPVeUxfIvgDT4WTXRoxHWfPM6upiMB89kYoA3WijJPoyPt03H/DGhsKQw1LkiM
c5+ZVQoZsRtRZlOxQSgMp9vGOw855S5Ev1GjwU4IQiY+xO/5L5kGonmbjI3JDOAn
zRFRzn1RwZ43yi9T+HzIcDtZPdiXHVqaRM4LVXxxNURME3naMMIFnVUGLM5gefZP
15MH6o7k2xQdY9Ogb5NTU/snggPRKLfSiT+TDmJg/uhVlTXlLRB4W/1jtOUuaw8/
FdXyKu/M1BwTei2b2uccOKcd8OMLPVItoTUKw2VYkLatN6UKxymfLVzZ4+5ScA06
LYwazEwRKDDwro0WHp72pdEzWLfPGbfxm4gcDpOXRQl2z/7ORmBjJEcJzops8WF4
xHw2LoOXFDdCJexbYFPoVzxpZ4kdjvymyQFcUUnBQ9EyW2XsoYSJl1VvKyJDs0cv
XxfY1Zj3yPpebCSCzff1nTiApdMyBZMrqBHdebH1eXl90hsp5md33oMsHvd6BC/s
nyKZhhH79rgRfLp11UgyPBQKIi4c+4e8EidUAqMFX4U/4wO2/E5qJWB960+4dQ0X
NPH9ctS4LOu5qP3xypPBkptkmL6EkIxhw6UHwC2m2vkxhlzkQFH8pAmcj/yPS/mm
Dbw4UM84WK+H8NKI7ZpqwUL259H6ERqJMo8ZHT3Q7O7BeVGieitxQaLDQYLicDt3
9IEeYS3Xwxb9p84Q5i6DAzkuk9DvD46e8gvA0QDq9T8WE00hUWwTWjC3t4SDDF9F
scq8XAQ/mzs6WebV0OBdtNgRGSE+pLX0Ug2z57+uX9URPWV9WKuQ0Z1wrnlhXUPx
epGdYDqM78obtAW7MRl6Tyt+c3t0psKRYS8cBt0pDj0yivDJx0J4Z5+EFKZtJY3R
V9d6a9JMbVfYcv+eHfAR6NCrfVEVcxHj3cxhDp6rewFbfboLPF212wXkMKlQK4G9
RfIrORBoUJSwYspYGwu0mrM4c6s1lCMETMWDVrko+IiImnNZimM9exv4OGMeAF4j
LpD9E3bQCBk2TmR3sVPxgV+hdUaQ5OEv6p0Z/ERPXoOfKZx+04kEwBvLnREiCnq1
ezlFl6md2ZIMOlEmjg0+T/gS2sFW7kepDJ8Agj617PtqQ+dkJyJFKsQIIrCWD/1w
BtGQg7Idwfc82tZ2MXXWTwKIhsWOBzpwPB3K0O8XAMY78+QSBDotK2x29fJV3UlE
cZMDEeU7K/Q057x4yJ+Fhv79op2Wsm3B011Oz0RBfoqPgpYQAxxsMW9IKpUiBrcv
VldJPY7iij2LlQE//eYRwoXb09xGLvgZlLHkF33cJIhShHwoQGlkqahemEtHFGHC
HBEm9oGrq3Dwn68lBkIa1C30LS+kbtcKna+p6Q4/tBrmw36RWjDbJJTl+VT0BwPJ
wxywRj2tN9Dks6ZVPbhhyiNeBiAB4h02hqANSwrUdjSc8skJIch3ZPP+A2fmd+si
ZgAz/8FJzvt9I3Y1rT0wITBh+TFXMqIQKIEPpfITI57R933tiAFrbii9ipDvkVYW
XIH0BT4Ggc7jkt7PGylwibEyQCy6Aj7WDaHGjs6tBoSGvT7bTG1UfAIYtFD0XPLG
fAijKxgsQdKeZdDyhRu9417U6r2ql+0UOx90tUgU+RepDJdwQOHPa9PicPe74xrR
2sjEeePIwP/JqDq0b9zdY+yf5SdSGvc0rRW6oKiTAv7kw29KDvqzyyNwCZhol0Bl
LvMCAMkiQHudsZbw//jHhp8TtuD06QEKQK2AEoO3IWZIZMZNaf3Dvz0B6lv/Xjpl
IBXlcGKyhRPjlP7k26FqjnJxdGcxwKeVdcZ/ePLRKeN/KZ0UYBG+bRPV1tVF/GZ6
Mf5ZbRM4HIDrb6AInDcluT0BofiEWRmLE14gICgDU/QYyQGd9hET6tZUM4N6Hkja
Hx6tx8N7jpcahbAZsYEWlXf98xFznUfHv0LqsDjhD5iN87/5LDtAdwMC8YyuzpjT
T26o7sERDBTHHpQgsjM7FSc0ss0thNC/fMsaB/pO5d/BXj/GIr3FakHHAsxmtKEQ
hdWfsf4JL4DeTcoKlqomtEF8ahZ9Ks3Q535YTJtvRdMVvqWtsA0achpXGbv+Yj9S
tlZpI/izN6gkq5lYdYAWD27A1Ttfzk+fXTGv4mtxfq4X91Lkj9AhFkSz61EQi/WN
Ru7o64VbiCROsuYf9n9K4mPmGhDPI/Hq5exxcWx0+nv7XaRUwZcjzulWlh2fKReV
7WMd9Chmw/Ju7BIaYMYP7G+s9CYpdTBhB2k7cw7DVQnm5++UUAhFEYlpvSAxqsSJ
27J1T7wlpV/N48AAXaWg+rzdAxvZGjoGL7lp4r6XjRQ1rSveG+COFv0dg8VIhLHB
DdSE1sqZLfMkFDDf7SlKLSVSM2Bh+rPWbGByQxYj2mRtc0feXgS1LEBOa4MAzE0T
hvBQs+9KpWFd/fH7aP92JP8R2iIBQ0CwFzjIc2eidfRi54iVUXygIIq3of4vseFW
kvcipElMxGwJCS/TjSMes5r4N8LNZix6CDgISYHdXQUi60peJrxib3ny5UCaU5nt
LlnWJUpwF/YQ0sCCSwWZ93AURhc2ivZw8aPaMiNk28WcMjASaW655IXbkWsmGh+Z
N1aQDMrlbPHIgW2xTsU8T20G1VQjBbFwxHyV4HNRU9sawyoCeGGVJjzNtKEyGay3
tzjAjUX3BNbhMJ2iNyLojowx2UfZ017YzuARBaxRbn5aX7blG9GwD9qQMe55ivzF
UrHsdORU1QED08nbikIBL3zKk0ghnV9M/nu7w4YdQi30Ycyp5vuTaWCsYbj9FmdM
fWoCnNiFbsHnhr+ASpHbPPFmQlh5xzlVWRMDMUxe5IY4LAC5UzjOoiw4N+FP/tDk
yJ2yLS92h9oBylrR48fRs9rU69WJA0nLTDfRgRUNTvcg7cqoYFyv4pgs3YGZBp2K
6CmTPLKM4gP4aCyvyhh//ZlK+RrNVUCK6UQvBKM2a4uZ0qAcdpMUzmrmI/EtH3ax
yoStF6+ox8CDQpmJukwAWGQQriJAcL5JBu9l6Uhq7anI7a5nl5Hv+0lUDevwWd8C
87eFX+1l2oKiQ4Q1hWVfjBNjwgWG+9c8NHDP8d5LKyz/eQuYIjWpvXdW0g1CYV4+
MCAnB/kZAskrfi0sJW5RlriTx0pvb0Sg8Pi0kHxf4UQq2PEffKOsf230L02Rs46E
HdM10kLBuWNo5EPuqPCBYLt/jsB40nS4TRWZtkqRIJe+z1xbqN9l1fbynWrt6oCW
G5FL9zFlAsCjXEcTk66n9p75Bw+va7OURJsEIxU0DkqpwzmfVVHzOXnDzTZt9hqW
iGBUbM7f3ss6ZynbxAnqFBekrckKhtAhEZMIQmljFFpQNzOiib92QvS8YzR2Onmm
Cq8l8H2NEF10KVS7cpkpp5oq6qhG+Iyei0+H+3Jjlq5gk8qiJ+oUgC4qJ24II5rm
LANFKT0Nu5aHekCvoyvfZRUaLC5Zl1+e865e7M5NzEC4ALGYDKp1jX42Fegn6tLd
gnZ8Z5JoD+e3zCi/YX5idw45lfTYyjssCUwjkTvMCre4esOVb0KhFJ+4/Ws1Wfw0
6QttU+ZqJ9Q+j6zqoSopbD6eqEvLd7vx/sRqFGPIGK82CJWjM6P8pxfH/lLgQK5x
KeEo2oStxX9y8ZjG7gOEs2MxOhoLolRraji7A6wMMAhjTMCqUpJE2psswIQIH9MT
br37lfF0SnV3WI4kU+jSDcfqZjxMcjIaZKQG7oKnqAg/zWPGfBHAbnFLooC0r2U+
qT0a2UVTVPz+TWjN9fvcfEpxQtbUCqgYJCFlEg14W5C9Pb9hFiAWtyePtH/P1wtH
ZLJhNOvoFnVQgSqlau3HUg1skjluBDAJUa+PAFeQ58AKL9Pqu9/ALMwVS5hOHRWC
uDt8Uqnz6CRHOmpK8HKdz5Q/ewy6Ckwa5K0T6h+TfGJktW0Cu7GPugnOE8WcNNmz
9sAMHgxITdASRPCVL7JvwLJUkfQ940hSkn35hNjdgU0PBmBvU2+BNzbb394bwAbD
U5O40po/7Q33aaYkGsqXXWS7OewvjWk3pRwwYWDHaayY+fINwkidR7ebBAvZU5AU
1GJsH0Gag2sOLMqm6e6pymxWfjq6uMYfypCuD/C1nohd74yac530boHT4SgM7x0F
BDH55uz1a2Xm9xTAcD6wmvCAf091QJJJk58IubXq+Bw0R8F85A5J+R0FDttP7cVi
9KIVe7jbP+NMTgPPujRB6fVxRClOqivWbDsh7MigXewwYekchewLxo06YTl0wIFJ
NpaiK3ZnpjsTqXO9iJC5AoMMok6rhYnaaIuEoPvgj6GRRWeU0btAcTxMSVGt0sVV
/4maUR7me4H1AyxAMuVTEkXs/Db1csLsJdSpdSXpVyW/Uee+XKVqjt40FonAFxUM
ph3+gxwIMPuaaTmQgHBEX6EUhBm+NMWCUa2M8xdNqoOkd8KdmYx5EXB5Fc05R8AB
9i/sZbBDXYS1V101hzHc1/0tSGDWHPsk08FeVCkQbgEuCPNo6qsNdmmz2rxd4we6
CCbyvjg844eB+Bn94x/5v2PbfOvCE5LxtDAD4IuikeBh94o9i0wrecN67GMtCUU+
9lpVwTp94PO8bAHL604a/qcBg/BzjdYItOm87LvNHzDeKBmL6+R13yp1xk/ui29r
osjztsZKtG/Gez9riCaLLkgNlJW22YLMvE9DGj6ODC5x3Odkb81OZYV8LUcrq785
yCErofp0r1ndlpvtbl2vVLep2a8umk2YbOf1io1vBiAs6jokHzbv+n4O1L+i67aw
ADnnK/kbm3oNG0iGLCvkk8jX713J8CiKPqVztyrMh9UPFnJ77LrWLZl3NijWC/lo
JtvqHpP+2OAv4ak66FvUhDWkTs9stxS/YCanYfrqg8KXmSoK8qLYaZ5JIsxsNeR7
s9/CqMWoLSfQTW+itn0u8V8JkeNxiJwCmRjHVFCTYTitygonU42Ysfx7hpmGMFpG
p/PCB5Amp4uTcl29LP6Z6ntQocilgq9HADyQ5p+F55gBkaAhH7LJuO1uVBKEcPcp
x4Bs+0wDnQifhU2acRNfFpI69uPXX/cYR9vUXtfd7ZzpEaSL7ATbcn+nMdGhhUQm
H50Nc9oVmG1rnkUkCTC/cTMLKQb79Iv45wzUIOnRkYi3wG8uCjYFlEhsCDYAD0Pc
8W3ZdlLuzZCGhTPtHQgg8IKVqLzNiWB80rrLJQYEqrO+etrQ7PNfliT1urrW5E2E
yTkLHFFab/8ZQV590Zi78CY4b5FmaBKv0ci8B9M1h0ITzIyVmpJutLcs0wD2n1Bf
5l/ZeTwqH5iPRtdz15vfGc6tQ2TkzYUNjvO7KT7LRwi9lc9TTFf2y967w1ICoYPr
USVPCw0Ao2vHHMa7vGJnck+nM/qxoExFi+trBaVl9h5gQlR5pMKVYrbX39kH3Xfr
Ox9Mof2YWdNw1pwy5uA04F9enTZDQ7FWJEnd9CTnuT5ERpON4Jt+i9cHFDipGYjV
F1URc3gYNqUomIMwW1XBoVYUmVZkXgZzpOwpHFg+Yt0/qb9y4B1HVlsN4/eNq8NS
6WYAgioEZ55FTYBkLpli3cliNXoh8BGK3h3uIBy7Sy79p7Bm3BCmdnDAD22eU0J5
xURYheGqbubRgHYNze2mGDrEPSUrLiJlk/vv87aXqgLDOusgsiWrzTgxi6Ab85pK
a8CSY81UuaXsSCuq11lEEsNbYy8amZe1jBoWDFXFuoOFWdyQI99w6VWKIrzJ1V4P
lPjmbVf4yqh5t1DPo7CIgITEqmogXELVs+itqbmX+NvQ3Troxzpd7OOOMqWsjdsY
ucEjxAf4kpCPNoNjObS3Et8I6o+9DINLiYlPKKciEgNmCQYrWkIrYhPQoK+Tq212
Yxf372i8eYX0R8de93CQfArPJDibxKrQk7ODMDcDJj5wvOPI06+P0w2AhXSFIv3W
D8UJGCB8g9RJZib4NzfgvLcQKF4xDpIgxctl+DBSJECXiDU6DuSSvJVFtB/cQ02g
+TG+Q8ch9Mmc9ltNoiW8AZBs31T6ULZi4MN06ys9Kfm0KN1q53bV99a1JPG2BwPR
a1Fj9wKSnGbxelSFy3aiN8v9TEufYAwVv6wR4EPJlgi1LZZw7fiRnwJQh9QGJ2Vi
2lmUCq7o5yG54XzTVuNgeN23sPLNYXju0BfAJ5J8LZ374zo0oNZbv9qGkVGIRQHL
RMPQlQdELmCnaZ57S0misWXdEBWfBBdgUxujaNSIpVT7gL0/aZnh9AIIkQtaqJ0J
1p/z2ObSP0DSvsSGRPelcWK3eXI5aMWWJFbenOagSMOfLYGHSFxbk7QLoK/54BP6
VmkG5mpwfT5iP6pumFweihr61Be6qpQEGwULIMUwIWKQSOPQlQ0ciPpGRXjNWPbR
3d5FlUb1Ki52g+Jtb8nzZDuSVxbAlcN/RdN5P6IN6ztwUlZmuJ68AnxFtBb8YO/8
GDcoss6Xh+1RSojocnrlngWl1iww5aXHhE73dFwDOqv4yTVZxCwptux7PmZJ+PlL
HLtR/VnnO12dA4wKdJC6xnM7aMEJPQM1C2l9s/9oUeBGsAdBuXM91pZmr0k1OCfg
0tJtSwXgHSYGx2FFibKND82KRbKrZtx08VZ/7AnzOfD8OiMriEyqsAzKq2HMnHr+
IqVTkOLPZJELSUnPZ6vBpUP0x/NgqKXHdiNlDUsVjunAaMKz57UMsqUv64rORUVh
uHEXXTUASg/KuAYdUJwxOJDFmjDzc0EWwXttJNNS3BNVGiVMIfUs4Fnb0C3Y1PQG
TK7Vczxkv7SxtxFKKtlu87Yb/MLxf2z/F2XRSZRJD162JHB2HzMSWiARlTEnXiCh
O3Cwr8YZX/YyViRZFjNohUsA06VTWhbpDnoUGuumML93v62ADJQAd4Wf39kD504U
Eah9ASqR0bkXB86kT3LdE2bWzY451aKP18oaY2jPHqO9stAAoQ3q+Wvzibe+HBhv
OoC/PbLzGcZltZdp1mLubbkHaMGA9Ufq3D9deZWLfV3zUJzReOFNViYDLnkOaklB
CDK50/7oCEjZrGRAu1acFLn7CT7Uod2BzOJE6bQoSjZa21jPq76kfIl4YEc4PCtT
ZHxVRJDu2VfDOMyYN/hR8XAOowHmH7w/s6FfbzheSl5nF2hUSJ4eoElPOVlyvkcR
Ldex2MStRD29ii+qWMsLU6F+cP+YbmwVUAHO0FXYsECGbawr+DG1BqSGyhepBWLW
obR8HA/3pd6XXSqP3Kt1GSbgEzHhaK/bgbYUNXX9e1vsK6OCRv1fjOOefymTD4OD
Z7CGvd+8TS4zjBhpbk7uSXN54LQoA/+Z7yvOR+yAQ664Zxk7ikyMnK4D9lXEg43M
QYDVzs+rbk76xCb8QtBwZGQDcFoE0ChIAXa+LAVBQsTvICoP8bh1i4JmncxJlPa0
pkz5wjyZ9kvbqLUjCtr5QIK2wZppbpuV44Vi/ZvCba6xddw1tfJjKJTSSmAlVY1n
fn9COUJAE55rK/AbhFiZVpzPXtGK0bjMB3ea0Z8M9J2Ook5qwVQ/JQnHwDtPtMSx
/kieh9/uFDL3EMzBxoYjyLcbS9C/5q3hy3Qy6mWeTZKsG8hvMEwYXYypzqeg1Ukv
NWcAd9i8xDFfTFMRvcrpa6UOysXpX8zEHwoHMynDlcZHr2dVWC+GGQQQiWXnd9sv
kY2ZWmn/8t+/qQIUg5tZerii/Zh3AuUukaiWWKw2ELFKF/hI6EvcD15YyRudUgl1
9wimcChtcQffU0ZtpcUA9zfWqHChcaqBxjvEn0UksLFCF/IWuaLiZgNmFTp6v8tJ
n48hMLkjy5wCXDtF+uNcSBFl7spltu1L1v2Lc9xqoDZDBB9rQTqRDLp0AmBonWiI
/zJmKK/aYoU+5QUkb+DrZsprmHycLAZicf/OB4YiCq0hwOUuVfFrthDwX/XiiqaD
LUdjzHpfZ0dcWreWFxzYPY7UUohZGgE4RNZIvjQCCY+ZcRI5FDD9hPDtnph/40Xg
6qvvKYc6qfGLy1zdITntvpduhf7UaRzW5PomorvnwRPnXw3Mtk4PtA1ydY1Jkg63
C8lCS8r4nEvIW1aIKKnypQEo+2wu5CpiZY0Svi14+2W7fnXlW9aHW4HDvnmaWT/7
VxMhHNij3Ignk84JQXPh5Vhd+B+vlXYutWT0AB7BfT71rFxGP2sntB4+fdW2ZJhh
4JZeBybBP2SVQ2mYIFlnjmu5dAMHXe/16uE7zcOxg1gMo7C34ixeoNddrFFJbxLC
92DvUQY7H0JDkA+xRVl3AF/OIrmdB++knoCR9iqk/k1ikmVvIixOOOubEVGd+M+J
xmSGUQcNFQ7keR+AAI5lTsNSv/DPjWoiiLl1eCtUPk/kBuNP7Wgf4pPAUOjdAbtY
tp/cI3z815G9q8oyBzK873mkdmmS4a932vnbRM4UZ1NhS2I0FS9wm8tdImzMsBIm
nANEaUR9yBZMFn4XnTTMV0GJJJkzsEqZSMjpjeLPx1TqajSVTEYEVxpfcepTZmjD
QIcMiP6JUocFuf7ZLeYaBhoExgbTv3Ue0Rp5e3blmUdvEtN4szOEjGzJ2RJAt+bk
Q2KSU33ShwOjSyUf4lXeX3gF8E1YvPAa7LZ+X+aZCiAadu4dN9zN1CKS2cog1e1D
QKgfRBNfXEilNMO0yoojGQczTVVryGnXvQvwwuQF8AlP/YT37xtaioMjl+7GuJ4U
D1aLzQA7F1O/cPkclfBtJqs8IJ5AcBSAkfxpbyUNNr5UfB5g2SdXSFmqzJ8bReNU
pWPs4zDzWM3iE1mR5mRNteVKf9Qk/ft8OwiuYBUlG5koL7mX6DAeEAUSFHW74lpa
6tzQDI5y39I9690aWfLBVaaOsmVnKp6Im2fhgE1iTRsVcfw+Y5exdSrD5VZDeTFh
iD71TqAjJGdJkUEqoKQFBzlIIaZH9Sel7L6Gh7lZg7VFPqCn8zxmOxcvoTg0lVRe
kfJGf0QKEr2JjRXJXfZDSZR0+DwV3ljKgp6ZRK0L3Pf6qytZhv7HegB2osN8gQsh
BwOVT5ata6Z+uchaymrwrSuBv0mErxYagnADrpyYpJImq8Pb0O0+84tWPk8oUSMe
0OsQOAIroe7tj7opmRUfw9Nbzgr2bppRdlLdZNi/HH5jC9L9SoEEL8GKY8XXVrRV
SdcuoaWMgBoLitoaYt5u2jOK9mv7GBBaebgMsMgt3ti7aJzjlt0CD792YrwPQrbg
vKmCjvjSu5/ClK584rHC1o9bmIcG92Zoo2J39umrh5q2cBBgc4V02SawQ4dQIiY1
TYDoSizosfBucwGRuiM+1lHSEFncAwpaXQkeyvuZSbfMxDo2apYCI1MO0DVk1P+t
7JHCwKxm3dA/0Qz8G4RXxbSJWrftc6DKuV0Pcuo1cJ/JbKxAysySMnZLnVleeX42
XECgtmpWLAhYzZNbGH+Q01bsQHKjXWKI29zHty0YGHO1W2g9tgKV/W2ar+Lke0jc
1s0RbC2CIv51rBX50NeS+w5wwGlJ4j8bx1IKUKC0scP76e9wD2Hm+/UfBRsPDdxq
kBuAjjffG/jyXdSyqtG/2XiokjlLtUwNeVTVW+cUBX8h3FECyXOZwqxUNZa7IaLg
NnkSjw/ovwgGuougGc3qkGw0jQkSFcwmUyvek9WoOAkt6vGPbvNFK4qg+Z5L3ibE
Plg+m6hvMMme9S+UJGKPpbqXJGwtp9jIPVQo4VLbN8ImeVtmQjBLtMBy+X+NIAhD
BZJ/tZJGwU1tgj1pv27kUVlVuqsR5eavJKlcQ+QWyi/6WSO+RvYtumlHec5GQSed
9kgcMB3lz14Ns14aHXPDPSXFplxyn6xz+KpbTdCeLuArjUadrXcltQ9GKAmUSJ83
KU7iIodaTMhbApwJy+Vgmmx9n/n8pYq8GI34KufvdNGlBhMFf00chWyLfI07OiKI
SiVek/mP/9j3O/TjiZo2Xh+AsMeEF5MSvSDPCakE61cCm/MpcVU5/Q/E8FQrF4aR
xBc2pshV9qZ3iJOpek9FzvBOxVKQehBlmK96HPIdRc8dxtjpuh7QqVjPeJochqs3
x7Y3QGfHPgJQ6gt/0u2j0DZxH7F3v/cWLmgO8WYOzvsaZT8KzLutiiL5Nv6ciJIT
xK5rbGm+zhk3qfhrjWsTpr1WNxEF0dj9jvuKOdgY74cey7NdZpgHforrLJL5/Qkm
gC13wSYLGv9TUi5X8AxR44ytjP2BAPbTjGx0dudi16+z6D2jb5Hi4cGE+JmHK350
8is/Smwz20GrmsHRLKOAM8i50vcHXqAlID+0Wd4OOaEpu4auQOnXgRQ3iUkmb9nL
XuNC8E8/dYozwdUsxtQRX7EG1U1DJPVCQF5pN3z8AZ4Txlqka1bbrPw5xJ7l0CeU
9qIL4+2rITPwxlK4Waudw5X41B/cJFIPoyvIntdYYGxEur8qb1Rv6gbDKMwBHCQG
vV3DxKX4tIUeSgv7KZDlTbTMwaupbminzqzXOBkFJX6R7qsO+fgSmspmH0b2R4YN
0/4FXEN+DWd6H0hOyBL2S6V+zUcXAgzeXgchebOhxE9muuX5FsoXL9uDHMQWwya3
MT3ZdfPEIR7M0DNuxxcy+rzyFk6lIB/yxi74R9IbxpooyF2KCtXnYO9GDLryzkZO
Fwgs6zZt2NneQ6xxC4wUhuLX8tCO5e8Pe7Fpq12/USYIQo5JJt/bTxfDakNz1g7f
b8iNK0jMwr+U9ucHx00CALMMhDnKgYYj7TKXPjuh1wz88taM+JcQ5prV3tdIgeQW
Pk4fiY/+3re3lfH+COENxJlnS7L9oqGiOVmaUI2ozzEcbyV9eJWaNHoedLRtZSdG
HUgHyYCKlcfzkb2fMhV5Vhu2+/k/j6hcHHZwkNiuUtpFiz87ZL3igd1Vw9S4ZkYy
wF5X3th2OYoNjTozwfV094YAy9Z7MAuK1KmKV16q8v9xLltpZ8mA1ULUP9/TkkF5
KKxZ7/qM2POsMpbVMBEBMivRsHc23hOvlWdwyKUfkERhnJTYsk0/Nk3G8l9DkVLg
yWJgxh8xIalX6wXoyWzGBzzQnWaS5Zy22FElT9EUPoTZF8RaJ8WS0Iowd3qEkt++
Ddhqx3RVAO6cCQ43yY0kN2Imuh44YFj7QRaqsZBxoEFZfTiJYDPsyjSCKe43Lznb
qUJJabMVxB2ZTJ4CqqpYgyurlP/YVM9Two0AQV4jRGOuse/PNuK/R88fxdrjoEsg
4axNPhVDuh2MKBE8kPa/DetYKXTZBWE5icIoOLl99C6s2bakIjThcqC0PRRbkSh9
7wsRwNjy6LgbCamrsYBbv/+dUc+zYMz8OCBc1evfxAkUsqNorUhBVVmblJAN0HmI
TQ6UC1DwXVfV5C8wLTW/4LqahMiAi+JMzmBwxhZDrMifdh0bcyXhsACFYRRkY9JM
sqrVXxrq6ttNHAZ0UxhR3RxX9p51e432fLEyMlgV8weGpYYq8DxoRqA8B0t3uMoF
abs7hIHBNsW0OtJ9V1uaUvuIGjUA16IvEQQ1L9qzya/EuacpRtD+Zlgdt+zwhOuR
ZMMzPy0N0S0YWwd0SPP3u7DQQyMQjMLg/zIUpDkx7gqZogYN0NyaFcUgjt0jLj8z
Z80ccQtxNlfOjaWjGGVDxEdjoEqMdDU2p7q5X1zmQDAXIhZ6rVYAt0M4W2q45/zK
BLz+W8plD4pwFDu4pRwKK5fPbzuLoKujnwNl39mYDeMwi6N3BBIjHsb7/M0Ky0ai
6w/G+uhFQD0VoQ2H/U+HGNokw8Vn9cJPU+Y8un+kYAL9lEmEXTcw3wr88ZDIgo9+
d3FkdNJVZxL9lgVGkUqym2eMIuaFc8hr22lYN+ym10u8G6ZVbIgdp9kQKQd2ZP64
lNSPWVjQSJNHEFsznDKpVnzzR4yIhsnTne1o2rlovIJfezguFAzbHKRBNhS6EPYv
v0a3jRzCaCAJNsZDBQvXfAgAb3n1NxUOn81K2OxHM+S5cR8VfjSaNwC5x+sZPIii
I/+TQrQ1oLIRK78NoDiMeKUoCmhoV/9i+hOrO6LqBU8+DJlij4pJvnWc5Ro0xSri
iZI7rc1A6Vg3lg/eEeTftHc6NyRa/9JmvUhHVu2GjNPEeHvkI3EWCjwaNHVCILti
ldmrwtmCKFdNFJylQiuKISvh/bq6B9q2lGSsyA6HI4C2MRhmr5tasbXlB3Nwt8W1
Xx4WlGzGmiJYrO9pAJQJd35zvWC0Ep2nZ28zrtL4vHrIv6mFEeehcLdZ+Ab/G1ZT
+OXGAwduCnJwu9jE1ywFLEaA1f1DbnjUZLOmydqhJ/GB3CHeMlkjTUkaUeVcvkfx
j/M3hAsUbvMSEFB+NHOunv6eOBicTeKioQJyTIwbaoC6muUVrh9qVLE701eZNYUI
/jqna949gkHOvtfaJuBX0gSNEhBHdeikLX4i4XHllerPz5IIa6I8Xhedg5+0EG9n
mbX9/C6ou1Z4wJACKp9h5W0tIw/ZHDXrLBJHKfF0id+DIz4oC0ID4NTNlIxKGuya
As8jK8NxeBE5oEQo+B889JbHXH5fSl3ttjOQGcduTd+Z1yHw2SqdQNGUGDMvnxyF
SXNAySMHMMqZcOhnHhoxPue/Nojz/cQQAZbo4br6KxwQH7yhjs6PKT1XRclUYLND
Ly+FLbELwfXkcFLa8OlJtShfJ80iYXch5CgSlItU41KAwm9x0Q4mDljqdMBMTxM1
vUN9LOFTMoBuJeQxAYy5akUJbFYeMhlE1hTWuu84Dtnk2sVevjgkT2NfBdUu6mCd
FNj2khUd/FlGvisGD52r+vp+xQXgbb52sT+nRpPxua+DeZMK7yPf9qTOmHr2u4cO
HjEPPmbDumDAUHCqxgm+lStVF6y1MYU3DUvhHrWtMO2SoCHQwKK1vJqUw0J+tCIW
FfmDGa5PAQq1+jnExGL0LWOJNLy7s1+QKRhmdIn8Sfl09pxFAq5gJg1uRNS8UAuV
EyW91RdLGXJoIHCvcileBDc4nyBFB/sBt/W5q0AbsXi4qybkG1RJ7dqhDcsn1fcN
T/3J3CKUrvpvqzbf67UG+hQjc4t2qvIwEAIxQheHxjuFEpIBpAMzrP2TtM5dbDsW
nZRGgjHAHDNY3OIJDfArDo8h57k/2kewORpXx4VvHrwJN1b1lk4Rig0U6CjajuS5
uBuQkLE4eEZMoYNVY1Tch0W+e94knz/Zmm8+uiGc6u3nPAoi7CaNrDcSw9uoSyoH
G34tBIknok3bYRnE8QKgRIfJSvgZtyQ3WssgwKiP/Z4nAjGPQC8hcQEXhk7uUcqx
Z1U6RTIED+/Xskcu20oqrKY/2DMJS9Ppf95Nyg6zfVqfpekf5LBG7MOvOmih3HPU
JFKULJiJcXpLwZqkmM8USx5Ig+Yr/0u/wXS6ggU/5ebcUDY2f29K6KKmJoTs0cQW
+Osn3DpDtJHEWDTIomlo4/YZ6C/Rx6V03Qs3UxyjGFZ34oiXT/V/iHRQIQTZgKC9
U4yY8/sOQse0uhb5avqQ2CcoMkJjB1jxIB5Lj9/KJMOWsbMgU8B5U2MQyrqOVHWL
d07z2k/QQOsFkTEVaAhDJLQloLwQLBtXY6KqGTM6C92slkv7Ff29JNX+9VJ8Oh+a
vhS6wCfqXtwweuBJCCTBBeNMmGjcnBDbN3EXwr8IJrT9U5NhpWb+l33FibzqaXJA
Zvx8fW3G76huqRlgNs/aLW+CIaR4qHfL7WtYtjY3rmJ2wJU34P7MQAkY3YkAj2Mc
ubXG+GCA7WO4JaMYGLoHWTEmCtxdJGFAu7KxkPiVQM7v0/ZOQERZSugSdnfma2mX
FAflZJrOSLyZXXodk1nr3Xth5gCH9AEOQDIQAtRYyolS20rPqkJgxQP3jn1w4G/1
b8yKp2ascrNx4UTvRlKDtF0nukdeBTZJezp4f4YQH6xl19O1V87GudNM7a1OaSRA
kp2wmGd9yppm6RRZ7eL/VNg2KKVqg4PuHKZW/e1pcPOo3SexPBz1zJpFSYdiFaIB
aKOkmV9mNOGygQMUIqqmohgB1rQ0eS9/tBkchYgeeS/pxS2QIB6g/IlqJ+57dOrz
x5g9ixHRvgvJNRDjsVAaelpw0B0qVSB9tTG9ZLt6gE65XileDuMKC/DBb67AN+R4
RbtJSjepsjbFc4TJAswIbp3mfaustkLAKd1zeiVXgVa+nHUWyF0Pcdzx+Od1xuEV
461n+DexT6FYumzOteAQe84XiQ3zBW/MRc+aGxvmJLDWcaFW5AG7lTicrt6mqJU2
+uaZQ+s0wirlS8wdi4VgxvLaNg1PbN3/pEJvk2Tidq4a+OSmsUA3Mk0I15kiJFa0
YCDPVw+V+5IbCtkCSrTSf3430nhwswFqG80ENSLn6x80oFiXGosbF1PqDHfxEHFC
yY/wiuIWeAqFuIlXQU+ZcT8CC6dz18bKExeG9zoh/9wHkpkGLT53by/uEHw6LvsX
iC4B8c3ce6yj8nbFxx5gVK0dHYWWRYHyIjUxYq107SqDaXB7mriewm5tSsy0bKFC
g0d44NIKc9UQQK3FAguIRg9pXbn0PgajD+0Zx6pQBylnGQA4eeYgyvi0wdtNz//c
SKCX0PT/Sl2GhgTgGGTWBKiT+KXq1ZuoFL633bbHTUxmqEARySmwkg3hDfIhJ0lA
MnpX/il99W/gpJX1DGk3/7+DJgI00wLgMkvvbw6cc7Ww6e1Ju5kB6boTIkN2U6ct
snXanIJNXLRPSqr6lxObaMJtEZhGhhMchLXKKmiQIYZet7MOdYsM6YrXhKUvmdrL
JjPDNLZIJPYXZT1NC6IEOlxqBXVYsIu054btHjMixJmT9QLJR3MHFVLV0bv8t3BL
X1p97Zav96zAAhEjstEG1SpibqN+cMCsddl0kvkHntNzmuTHcT/9digwCA6cJGbz
rWV6nwonLwtwglVIPAVp0eQNBz1IHnHZRqPBLWbOChrY6s/qh6dj9sIHP60v3xWn
UA0P2F+cRyHLUEve9ubDEQlKRi0uO2guzEYplhYUYdpjeOjgPig8aja0IAAX+KXr
3IL2S+tvv15yEWEOrg0NKT6J+Rx6evMD/lVhwW8OYHE2xbBn9eJYbOGO9locr/VQ
FnlyZLmUmQ/qx1VRDd/trgM14r+FhV0eGu+8SbuaLwBFa6Ne99G8Swht8GdU33Nj
P7Wy1hzgAvszcE0+NZziweMHEInrCoI/fixoeFiELM7cTg26WCpAPXeh88f/UEp/
SAX9QIRjDG85pCOjiVPzJeJkFPve61Gw/X2SKZiVfItN+IXvCN2wnnEjA0IL89fu
oCoD7nxEcJ4kR+60FZ0Y0xTS4vZfifofRX7SamhYkwyEjsaL8gVKPEJIV2vNvEa+
4TwJWjSyavMJC/t53wmzAqhWtprYZGg3hjBkdeeDp6aNAJdNYhXGyQc+cfH12+2q
G+uzORXKh7f6Rrp1z/5mOk16eCarmw2rnc9K0ZBlNo6fUZoFmi2/Pm7bhNXI4lLv
jBzAXbEEjI98EXZiUrR4ft8YXEjSIJ8L3yMcneI7LkY7q0gZThVCago2pPZMIlej
gGsn0p8bBr32z29eLzjrpDv0n80Bk9p+fysMaFakHaZ4SJ8lvnUcE1jFBXO1d0rD
/hiKhUPc3MNG+s5PvFD7CsobYNfecUKaOsAyyVBPVSQM+T2MbR/YPHrJ6PzW1CaB
xeikM5Eyl5g6elWXio/2Eu6vO57xHUqVHQrlrIWekAL167dxD9izjChNR0LMZpnW
OEZ/Tq0MabBgYLltK8rEcwd5k+TItwtcjP21WFNidzajc8W6sQrQmL7Z5bIoiiRN
c7CI6mznM2Ox4SvKmxAvk0gez6c4dvzBz20evm4AdTcC0rHQmkXtgmB4jycyJjle
E2uX868wKxXmqUCc03ujsENCdlEnBFRxcmRRJsGYLCW6GKM93RHH0jL0y+auX04E
1ltmB5q3xKzWeh1/DkQmfCD9qAazawobPWgx2otXFcNwvhviADNbsiCTzWGtmAhY
ywZB+mPLZjzGCflBnuOdkoVA7wq16G8Ec923QWVOUBVLJ3hvyj3WQiE/LOtj7cGa
+kVOok4vTLluIkIDh0rEJCT6ZIlFTuiXtD5WUm4f6jmYEe4J8n0FPcy389n4EXh7
OwMXNbqU2nDyBNxe0gYE8auv2StGI1N6LXoUpCYrYq7bX4//UGUKffpcl5D5HT+e
NVYpRYWZGN0c7My2RF3H/ay61fFTTXU6eq9Xpe5fDCtAdd+OHc+vBuKGqnNa30kg
dEQicntLhtKQnQ/fU6eBU18qWgSVLjToFMRjlypzbRSBwGD16xF2fkXbCf5qyfVM
NFph05oURiTakIsQ9fXS4t3mWbFTjfPV4QRee2D+zEYHLyHYMhyAGQPnw4lkG/KM
gL95fhfquGR7JVu5IgAmpoXe9KkB+FFlrzyjfSWrgAW6Ua1f7h0+ivj+bePGx2Rq
lXmKDqBSDCogetNtXqKVrfZuYz4nDRZXfloogK4iFC+rgoHvsRdCXM5L52vxs/cw
PqYWsei409IgIoI5kcg8UIbaYKS6hZbceEYtr1OnN81ahJb0M+N3vsclhci33PhV
KQV91R047MrDQzsfdIUgJ7HdKsK8PyG5i2rNaPiw76x6IhcDUGw1XcqIl0OnMvXJ
MWQb9mbwb2D1QDSEAq79EZqXtr/Vqa9nAwxIeBHuWvws2Nnnw6p95KiDY83OzSeZ
40DiDIQrIJcdMBGS5aDvAaW8VgRtsKOsIOHg/hTedSdBqga9QE2e2s17+sPxXdO8
NZX1tuRr07z+XAc7AWNDiUvQiFhpQKF86uKL72wXmW45MdrhoLtCNicMyeEL70Qn
r3vUVN1tZ+raFTg+BlktIQ37ZpcbWqF7b6m0VaZPMUCep//KlZx42emkUMczq7MB
LN322OBLPnH5ciHTft45O1Na/q5ECvAalbwpq4O0bSMgwWYqesEVSAnjuWop9rgj
OLDOf8xmS9BMY64J2pQBMdslGrKHk4JFTfJFgVv7pPAS9hNroMB7wJ/6kBgURjbO
5589PDpDp7E3EOSfdskFiCPqUpm+Ir8HLWG/TxJddkMHdFxzktj16Extkr4YZjyP
NkDK2tomNZ1JkHNgjPVWlixE6Li8brNk4/uq/GkWOn8DM1wB5jzM4YsxZm414chO
hOq3E11SIwMaZSwTgy4xWgg3EMHEEQ3ElqK4AF3mDcf5/foD1jd82614u4Klh4qt
pkp+MlFeqKIx+LGPdPmaEBFHdDpX1qNWUab0tF12xdnYE+f+Q1mFa37dygGBm3ri
m751jKPqu2Piw6TZntUnNEM5FDOGSUORr3k2UvNXwJQJScb/yoSW8BbBeu60mGGZ
4XX3oIY6yCHJ+fytM9C4/3/YokU5podtSkMagbCIUMt8cuxxLkVRY/wDkxToC1xo
jlJnWD0ie96bDtlO9kTFVIqm7zA8gRvhGXLPSMQhirLot13N1Mn7g201gLLNFlWo
27rv7D01vG4sGtcBI8EpIhXlRVWgr4jH0suWQuwNp8lJXD8UtMdSKj0LiDWEIkfr
jI9gUCt+YSYOnMUqisYHhLQIVuvdnkRgEofaKzFNt7mRLT0Wvn27HEZzLjQwVupo
LDvO27Y4wqRVqC/f0OUkNJOq5trL0a9GEB2Ku2uV0IpXi8xVLvPfSJd/CUAv/ex8
luLKX4Wsr25JfUWhNGp6H3uU4kpMNi+My4hDk8b5+VajPtNXZX5sFXXRF7ZKEmhw
SRzgty6GDa9AoGyWRL9WMf1+li+PqaRe6G7OoVkInYj4fst/RVxPdEI80ZnRJp6w
3/iLKM5iTUMLnGuDUkceXrz6j0NBDmArkZdo3ncbP2Ny2GyOy+TbulaV5z/S/0S+
l3+u8MEvgQ7c+Yn7csu6Qjej0gc1YygoYtBLcswqT37jMn0UVgoQTQGooNrlLhND
bJRCx/hzJJGRdUjNbbLKhvqIogWuxUJ9tm90c+fA5FcbHZXQLWxvNO00+B0akUQM
tl8yEchp8c+6C0t/DTkQgJXjp+hleIzTgGn4fUc5hU2SEo/L402atyXY7LUyifsn
qZL4oGhcepXoSTuVRsNJY5EwBkN80B7+f/nKstobe7/pqX5m0YeCWklToa6BJDI6
UJ4jlFYOqJvNTNMdKKJPOnl8oPK1PCDxuAS3Q1q2A8SG1++p8nL5uTN9x3Bxd8xv
WBtqucWju28GiDj+5PpW7rzbiclutcx8xO41jrPnVW5P+6IwPLKnK82oxC2qz8Th
TeWJ9CODrcNXwVO5eImNh331e/8eOvWecHggxn3jCHRsivQLiSDgLtIxnq80zBAt
GSpeuxE64WIKQ/HBnbfdzPQw4uy4Uc8go4QiiSkcSA0UPGdTRP85BO11Xast6sf2
eFPIQv0IzdUBKcWJNkmCW8s76BdTbFXfxgSaJkmC+EcE0JpiXOUTMgbZAbV6HOAU
9OPiZnZTqPJ37xwX9l8UGf5p6A+Ydg4D1bFDGAY78ZyONa1vxWizwY5OIR4SmKCf
4vGt8T0vsA9mvC0izq9QrpltJX/gn66r+TrukHMNWalLd4JOmPKo6J3+0hOLGDMF
mIQU493GubSFBVhuN9dRfq0TltfAoPx2suuebwJpQKELhB4j5355ZyHyD5xyzOrZ
ly/exLdKHHu1S5RjZW+sPsGXU9wL/5yS3QawL0dD9T/TpK+HirMsvfg3fn/zMwEI
NNNLUEKClsUSxEylREqL6k89VxcTmmbilzzXRPIfg+82l6HI73A4CmbtAzdxAIIe
wI+Jhs1gulu/JjWxC9AZkilk8TK+ilqcgAM+rQMBbQQB3EeOjVMJsIhR1lH+b3DM
h37VU/83iVQtsL3m2QKJkaOVRv0aStsFgoUByhlMubtSear2KPA185NYxuv7BbWz
P87u+LvFGbCMvQ5xowbBKvRfHnuN0zNMjcHQ7u0TSXBDldfZzPBJDcNeGYhvc+4H
L1e3or81Sjdqp9VwfvIJmG+6PqxW58xQWhriaNLGIzQWVGQ0bbfqRkPu/ZrHZk51
3odDildswbkH7kQdVPH5udjOR24W2FDQnrwxauDn6wmA/sDDftiPP30eaKqsbv7i
CMA9SyhzVhp64glVet741s661N/teE2AXoQeoPgY/7m9rLv81mWOAN2yFD3kFNCo
7Uehmw8nbQiiknCUMor0H8854MjYwe/tjfm+996CQ075IksHoXUokGDMUYd2fofN
sKmCpAtEupFreLACpuT0b68yKXdkVm3nkGzDX221E0Fq6riR97xKBmLnTdwZmAnM
UDM4Jh6SMGxMHb26HW88GwubBcajfkGKDuIXVXeCZotrHCUSvEOGWzKTzC6MLecs
isx3UGfS6+/+EJf0+x4rdBkH4UgoVIO1VpXFB9Nk5fBSmoRLCD+ch6YTdLhDwhH8
PBEL6z74Z+s3IR99c/1yJ3YL6vWC5bkZ7q7witldB8P5Y+DxzEMpeOA1IahAZr13
Q4tOr51+1iNm95HEcK5/YrzDXuM/Q/7nkuC1n8CoaiMswv99yz6Nha2OKywpjxAn
6Bzh4N/mT+FAZ/qYCHUJImwHpT3P6V8o+zYUCqnFIjpokkbkV/2BgSs16q6bwB42
clLlBbt8bZETnSZlg48qMEviDWPq1THOjnfyE6mVNjuSszOHPgnxG4B2ZzZEBDPG
1T7SuPO4sMB5fbcWGcNjgYQxQqFhECO5siS2Zm00cDQkYkbwR4EYJuLksQtLB8mf
KjiWErniVpEku4udouaMBG3/Z4WU7JCDkz/D4TTEhZSFsjJ2f3ZKezxgGvv4iIQc
cfVMdgJE9+3qWpB+IsuubdfHOvL9vy9Eh9LMD0eYwKFOVxj8+gRkLn45dR3bSEz1
X3HxKVXiREXh1HuklrkSMzS79lowXd++mGfhv5oOF0447lCOmUgnP9SP0TXFAG9B
qN+rbHwMtCdGlJTbKDmF58XRxS8D+xpxemuEsCJhsV4buiJhOKCNn2bmU/xmqoFi
cURv8Njg8RUmIRKPitIDf8o0RMNYg7l8vnggA3E3yEK1/uk1MtOH1cAH686J2Fd6
VhLyYOUF0VBZXjEZ2RTYJDlx5sWh0frV6RH+MdL5c9haZDyMHZE2aDrMsWzqioB/
CU4LN3xeqeVq6W4+H3xzMo4eFwqi5cNc5o9CRt/V+1LOhVStzsaowr87MxdB+R7b
QHkSftFFlo6HMtjV09vR0im+ezXGQH4JaLskyM+LW8YX7NTnItHTR3zeCIDuGmtB
c3MhCB/TVmN33A+Zw5/gsexvhEcPkNod/DDdTFzGtjQPSwuNaRjSx7jHvgNbsYSt
3fzHrGc0FTK4gu4ESLPkIHtphl4J/J4gA3nkospvdStj3yiwzA1etR28xa5PPuWy
u3cXIQxOqkl7n/176sSZjMEhciFLcy6D174ehpgbfSi4k+ctkFLb19AVUy4xjjil
mO6z6CsZ0I/cgkfEX/B6spgjIj6i36vIiRdi43IwjSQFe9/f6GnlS9jvH0RbSRsB
jMBf64wVWqHc+R4MjSQGf3xAgmvqHcOSQvQehoy2XeO504Eh3GANKvuGqhGtXaEM
SEbOGh4JImEU3AKSpfVve9dlBypr7AFq2Q4Ad4V5qnvoFFY5YDh7y8kMFNFML1ec
tYWfFIv3cqAXvGEC3rBaAcMwatwMWXX4ZgdwVLEn1NGqhREdkhlVHN7qu8IJ3Ipw
Bcpgx6wk1jc4IlT+fSt3jM1XL8T6td9q22PaGJifePct2rQgLJ8lgIRsUru7FCMG
lZAK+hs/DrTn8dHxjf7bXSt1iYtNMrT9lLM5wEkaJdvwCof6xL1vhbkL4yA1kyAk
dPri8NlbUz+VnQXaC9yBSPdhIIFUEpA7I8CwSJpadxQfRv0ZKHpVgDRpumNYTq5G
kAbz+KiPyBiGwcMTms3+CiwHreFdmaq4b6cFFuTbeFGlG/jIjfFcKs2egKAuQb6v
vJatYrH3Pf8qvCNblSDZCuRA2cXJ+wCD7KXbJTtTwNymHqO/D3T/D/dbIcIQzcUf
D1k7A2H00HKF3zm9Z1f7cUmTs/uQ6IfQdYVi6YG/rjHzMN/Iu5iwvH1Ni+BirJEU
iOXMMaqMigUuaa2JuXsCGt4vyrhdLz7LdrB+oZoLEEiTwn4+VDS54DGj/uX0Q8QT
okESLrvTEBc4kuQGFZf/+YPdh2hAEzi4EZOEGHaiCC0MvwD7sL1ZBktGD/6wr4H0
klFAe7BwgOi/b+I9mypPB9VWEYScAoVbX3e380JijoNM2spLCxPqrp/hq5Ag/17D
O+fWkAYuVDtSHopojIHRihUeW8YzKJnc0WG+DTwglk4OlleTXhF2sIzU8VykrUka
8G+yk6Ir6K0a9vWnwWLb4SLDZYIQZO1Y46VIvZQbnWThbVjdCRQ9RyhDwo+DlZxe
pk5O3cKmjUhs+Nk+MJcyqVeUB+9zAeVP2tezTO1SO6i0T+bXaHu8z1KWQLz2gWlr
P4VgAA62jEWnSexqr8XuENsxIuzS4ZR18RPotiL/3gt1VO476hqKCfGrChMAPTuU
hPi/qtrpxXQs7lS/moyPQkDHXHRa+XhsING0W6TCsWR3+bWEjbf9XroQMlcA973G
9Im2U3WQbBiBeQoZjs/kwpxy9USoJi2aghpo4oZEmmoCiC1af+5RKhE6D6DefVtw
UU6wUfeyBton75kWLEW4RTdaFSuDUWBmLCU2CwA7Qcsr8+sps0hEWo1hF+9tYNxn
pzdP2tJRcsfBLvwZKIV4NpBR/RJPhuhbX1FtXbrJO+YtFhszqaDk5Lrj6N9122NP
qfyZ9+64VMP+nnic/Eur1Fnda+us24dTr5MAh6f6BelJEk8k4ZL/gS4u32Ge9tas
T+tlutTCmUH25dsun7/Ry2iRtP4d0Oni+SohwR2pbABybsW2pHoLKw1+oemRTkyc
hGcgAgmo6SapdIUg7GRFQvvRnh0tWzZ9cpBdGrNaMRMVrAgIocBb2Sepvx5wFwRH
jbEqpJlc2T3o42d7Gsj1F5XYh/jPmd2KekcsSRl8jkaqWRLloKX4TZ3MoXGU4fUS
6lr5yo6IrovimMwiB7NKmjQVM70YEdVAnKbSNi3eXm6jS6eQ5BvbPwmETW5WyQdI
RuUHq4ol3HYyDVxpUjL/KQAM4j8UNyiMZVlL0WbACpEXZ4e63BcToPpWZ1GXTFnI
zcyOdHAWShRBXdvg0gz5gS6sjkn9tYILxOsduqxFT3qF5J8Q46UE3ED98XmTdlYH
jQlZJSfjMfm42fDh+tFaVDpGzpkzJK1+H3Zz48RjiIMsEADdpwoBWLWYTwcAox1J
NLUE5+DVz8tukfoBmduvm8mIL2sWAwh+gJmwN9Cp3tRI3MhSEAwH140uRS+bH9Gh
72aY+wS/mkvXDm5T//qL+wlR53L3vTjv9B9SUMuVluNC+aV5JHleG/nU/q5EuPuy
AMrHwmsonq0MznDtkBPwJz2JvLnNfyNmMhaG1Q4WEugvj79D/rk0FDNJeN4FIa78
GIaFMa6LBTYF2Gv6yIY4pTXkaUPDgy1dmQgtf1I0MKlopY0i/Vz0D/KFSgik+ruj
fYfvm+sHMHzP91oWApkQbe8hPGWxY0UPWzigrpMK5GYKWShgcXErZEceSYFWHyub
HB65Spvg6iiaKqFlCN7o4UaRSiMbeDv4p/99hL2oyfx422+AuvOFp342Fz3Tg5tX
PCKLIgtfZ2SSlLWBJsOCuLnvElzM2bfa526S62MrJiuwzMMivcbhGYp2ZSdq52+I
NBv8RDz6NOSDu7gcHG055BTsk9ihlUvX0ye56+zvKwrH6p6IAZd+nYR+mQU+JOBZ
j+DeAuDy7sP2RV8E4GnRNm31UKY4ZRG7R1cFm1tO1OjA2Yq/B+Ppwf7jtVa8bZeY
4i6dzSGXP1JDTGHNDURYb6qHDJPehrXWdSuqfIPI2kSAoBG2OLyaHDKY6iaITkyc
+V38kOl8vdC+yNUC0I00aAg0W5sAO9PQYE0vvapFSNsmpBJknMkIWq7XnlZCIWb4
uOW7FAqrzOUG4V/bkcnBZmR87Xa53kh7vFjAfb01YKtSWzhSTWgXTRM7XYwyqWHi
EPkeDLxFiHUYXtNBSbFao3GtUxpyQTi/pBZ3WYlr1E1W4WXRyeYWRjDrbcktXvRR
PIbxGmM2ESj2RexaV27ZYV8fxmC7p9dccp8mBIhxsGhWwUq/IuCLdS5m537tSfwc
JwY6mxX/K+P1K3HylZ80rSbfHM2KLiK7hfUOzBwyDeBnMjpUB8K/Gb+nFKibZ+zH
w+ikNVHHRUyeSCeCKyzgeVSPwDasH+RLkIs032ucdz48/K+O/nSRTQpZS6G+Io0+
ZdDxZDBaBzwjpQC17PYSL1ChBIKe3tPQjJl36hGSY7J3xtDUwM7xi9HAS9Xr9Bqg
KG8lEIsSdjusIyqTv07wirY3pfJNpP0nFIuCW4sH0ZTYFduvF0q8HR3gH90APCZQ
Mdy3deixWatxIZV4UufXpb4Eci1r4xgDVN/usooRSQ3dCLuVjqIvdcf1ZZSzHHFK
r6KPf0G1azGZHOGkaDqKmStsaEwd0h86hM5uRh+iIISvdYxbTUvNhCAqOTSqlzCe
FstYy0fsVDuIYCa4mXwG3uk7yrlsDs9CI2nh+m4UW/QsSWOMFyBM3H8HsWM81QTY
wLiRwTHrr9OKJ/x9spT5gwSknTCg0L9fIImkAy5hfANTNgLqQ+YzKqHt7swKKdFD
rtDVyifcNrdb9MY9YvtHx3mGZtnmIjxJ0yFtmvcrFJqOSGAn4Solm6ch0RJtWS1O
4dH6hoDuhHB/SRcbaQE36/Lo+siz+WQeVooM8h2c6SlMYp9yXifE4szpaNcxFq14
3oXDTyFfITYhLUGkZHY18y3FYZaY6OxcAzutBsOHbdBv4sVRXb2wW4kdHJx7mM1K
OiSG2xhM4ff3de9OnKz/Qoduowj56ik3oV4t/bGVxJTwVE/DD1ZqV/3dtN4nyzI6
l1IizrL8hIoQdUCu+c71Yj1qCGScgdIo2vGr7VbHHCG5eHGOUf5Amdpm7N8zVrfW
qu7bBOAKVN46ApeCpR1p07GE51EGg9FH7hlrMcFxV0CR+Ob+XBwFCZu8iAuKnitV
eAlUPhM8nTA+f6TAnQACe1tjPZRXf5LvFA19UbBulGHkLmrS3SWKXJGh4BPRF73R
5UKjzwD6+3MbCWj1gBXNKxUr02iILJbUQLjO1MSjfFb8pugfyvTP9rQBHP+h6Dz4
fi1VLjrE8NJmMd2gDgS3vMHc7pizwB4WjyD4HRN0d5IgWqpYhaLoxqlirylwfnbD
ePDLJUe0dIjNvc8sWbeU6WDwcZLn177RX/C+X84VXOMua33TuRDfYn8x/tL9/8C5
dYHSQD5CjrP2r/OxrSq6BDA/tSDQCqVE79mQwBpciM+8w0acr15ZklvQ7OQzGEBn
VxRHsNxM34m9WLIRf5fRR8OB+JNF3eqxPl6JiJPjtX31/K6+R6T2+o1iA+bnmk7G
3q3p64hsFP4Hgd4JCphhRJoYdL5Iz/0AcJTzGg9Vi8Bm6pyn/sl7NiTyVHOf1PGe
6tK0OHMwkGijkfMaLPRYpgOTu9jf01ULhCqj8SmwaJRKD8XUL8t3gBMXXnPbbj6Y
G9Swcrz9Fj1AXZUfn9UgyK2c2nuG9sDzPphRfzCSYuTptNDJjOs0ymssTRPRR0uE
fWwKyssiqOP6DW1kxinxO99IWvrjdwEtk6Fa03/N6u8lb/NBi7jol9F+7tGq2Qut
nrm/rH1DsP6ja/fd4XpaC4G/3kTYqWKFXAhIPqLaI+i0w8EbIBMquUTFxfugHCbo
kPpj2FdQEpDOaybnvPF6SCNAM6Zw7v4+8d9nba9m5EjLAXW0HBcEftYu9JMWLfZQ
d1yKa6vPAtXLjQEcq1FvjPzLOLysOt8ApbhgRXR+YmCnKDSJZ0ccZsVH2ADsLb9T
Dyzji4/p9LwPWcSPSYcf8fK77mOnHHXLh+9030f1KFSzGKnhMrfOUFrxJlIo0aQI
GJYef3QA3jnSEjvBTca80+IEH6IhM2i7QOdgQB97gmT4Ndcbjg6f2uLA/LSfyYH8
F/Cywu879HfUf8UOQ2PXHeUyfEd4Y6xmgXbdO2B2auFg0bfC6tQxOrC8OOuD6e50
RAEF1JfZf5sAZ4744WgtIbIONMRAc19oiXtP8yJV7vmZRPF+LNut3xjW1RfqydqV
P1VOkfZxVTjLGeroL20Lo9Gs8Qlyi1jqMuvk5nTDnWEjMA8rMloN1sKVQnKOTMHE
2RwTRjpQPgw3uHdF6nPMp0JnNd4EREuVD6IHW+BS35qyrUvrmXz/4LeftSJNBREn
Ue2OPity6BWSt15vrfKSLTHztkjXjWGS2iQ/ammpnsrF1QWdVb2qqLIa79a4K4qW
oO+Gxg8wSprMWhmhuzwvoOXNnR5XDZXiLuXEsJJeBd3nDcta03PAqTMXlCH3FK7B
XS3ptPehkKUU9JsQuZli+5njHBtyt6k3jWZ9YSK+u5qyQkdOFGk4l5FHNCdMubNf
h3FcUZYH/JtCNWTMeuiwof/0vWNoYhM0J57GdfvwgGgMOy761UYomlYh1wAkpOJR
SafV4FxrVQhb9PN9Aqv+Ui5SbwtFHc69qf+YMXT5CzL2BC3JI/Oi2I4X84+EWC0H
8vVud9YvoONyNBcde19f5PCKj1SeQHgh3p9Ha8Ba9qAORHs4R+XCWb6zVbzkMAcb
W3W949T25oBqu/rQkXtW7f3jQHQDkRNrU2nG42QibLwVW6TVfuVyIUegoRQIy2e0
3/qevbRgXJ50LbgvxaFt6F1a4rohrKVpKr9cGk9NxMQlC/EzZd28VgpMcNo1Ed7t
mtDPRZUM3utwGDiJ17OmBXRwrge+1xN/Ey1syJicafx8m1e3zSEWzmI1Hex/cBNX
ZbeZ0sgOe/NqGe8n5n82EesKRnHcNZuMuTXu3VsA/pafl0lVX6r1YXcXlc1o/GY5
X1FDKLCqBptQnTrPWawRVah3mJxZa+Ol6EMoDVp01SFi2oKawNa5cJqIFC6uysWD
rhs2PwtPz6apPc2jJld6Yj79Ljy598KY4fFTJgUW4gCe9Cj0okqPfuswS86zIFWN
fNs8uq/tFOZn50QCd8Slei77x5WAbLUaNFnM/PiVEDk9G0UVSjW/wiMrnvJ3wqzT
DxiVFJbiwpovApnb5cjN3Bd1Y1er3z5YwS1jyQaMxTQuL/F5jCYBmgm7IOt4y8oA
v0kKSU8hu0KM0RX5+jDCqAhLRT+knvS38QaheMou2vfOIAGIrmVaq60W66dtvQ6e
ct4bDRIHL71iABj3Fh0WFg2xZ/jLFOg+rCz56zW1zrmgxT9JTRtS3mJ0x4DEzvxK
rtoGdKBVkof/jTllqdLSPahl5kPTProuBznfOVgfsFU5KO6owSjxyxcWsRjyEudo
Ql1dOGEoHm/kSXoP8R6Kb3fgUJkd68O4p51HSyxaC9aeNHD/O6c6PkQaWAn1n/bF
GjhNm8O20gGiEVu87KUet6erIoY8QuwSuY5fEpNFcky3AnyfH1CYZasNHRQ7gcbU
V7MKBto22XNCXmQWARLVOcYcGEC2xngILIzWJc4ShsjkgTMnm92jQLjK0hdgy3mA
Zc9On9Rc3hlp5XFJAC/gWkLUyDubl6dKsFoHi98Yg65O0I0QtusFwwniS0Ueet6/
Dm7LQsbRFh34dHLeYOm1xeRilxGFC5MNFXjW88XJK72PQGysfQYRqUMRk1w3u7gR
N86uTNx9yrQH17RrBblIjrlceqU5ArllzEsjx4mltIz4oIgv4DPvzca8aOnod/69
pF0WmSVhtCuyeIHpO+n+nrHz56SXOzKeKOH1JXKvFRs/jHkKJ4+41nR/3xfkGc+4
icVLMMhbvM+lNZFviVzT4+8F/yOkL1PN9KvE5aemBgxzaSYnaY/gljeztB3gQOxh
hcRMkMYZng5YwRGwyoNEs1DvfnbGmDL+zHXFhhofa76pwoQudCr971iEC8AQqsvr
OpZKumqDjQUiZR+umaxu6sa0Rlm479N3V48ae++aWvEsxJys2Ffp7IYs440sgiW2
+uxQJmoXZTDGyKp7ywtKAGXb9dhslC5H/NNz9of50yWCxmmaLZMD4WCmTDm3+jLY
puKA6rZ2JA8dD8C9o1bxoAszwJSvhnwi9VMOqq+cdCb1Cf5DOGSuK70CiaYegIYE
fZYhQ6L+evDwd0cb0GtFMx3zr3bfHrsbopVufsLRpaBx0q9w+SINsRQNh/gIK6Nq
yt5uW00a6vJSL8S5vRkzZrxXNb1jzP4YK6uF7Zv+x9rXucCwfiSc2QC+4pW03sAH
F/IM610o6Oz6xdMV7axMfLNZHZj8SkZEXsXlapQbDnSfCM9uWCRG6+HJ7zJ6Eiku
WVyOJO7UHMDKx1k+UdGoR4PfFTcvs0ZQ2M2djg2+2TE46g6u+XBgCOJJEk6ZzkL4
dthJnXPleYIlzZMMp4AXSmjcGw3D6tBba5ChszznQdnAuzl+oGRoKFV2WdrvsDhM
o94eFmG1Niv/+31cJ4V6E5IGx3pAsHE4+zXgnWEHvozvaLgy3d8laSRMaxCAvjjj
UceuO/VAhNctHJAk/8CgCpsDFsdhHmVDrBux9rjsAFoJYqEdX/EcRdeZAavofgRu
wLd2Q2IwypTdNDC8o/UkX4ZlrCnPF6OmTE3n7XAhkZ0mkUhVWGvWmr30Sa+PAWnH
0vZxVDSizMT/nuWNfT8T+xe+pWosYekNlOvk28ZsneoD2Icvwi9RAR5yuQIfROhb
K/Nd3DHOj1dMq7t8j+Ena36P9tJT+xaEy+oEpPeUo+KZB/5y1r/fSpX+WjpPtDOz
+6mo5PVbhOTqN9nXAhaWUgwjdNZxzWmVqGBz3/OYZ963/oYkEGxICKyMB1D08f7b
84s0aV2m3SbJv4lU7u9p7z5fLBSsRCcHCTFi0Zkb63KUpVwVnagV1Lzp6MXAPMhq
u8r1KzZEz7PlN3tZ7RAo3KqUiW0y7CMrM/cbN2rl8tyM7ZLyzYyvV5A3n5iZXaY+
GjbE52HpjuTwaTmWGczmB1r7b/rmveGq7eoyqn0wOL2uS200aMgWKQ7cvvcTlTcX
uOx68ojb67YdY+0UvfpJ5d7gwumhCWZzU//ru7AsxL8FaZCPsTA3tP1BVdeBTYuM
uKTgZjEXmaOIBZeuc5M29hOq9rDVyYIGQ/2VrRDLmpSNG8FWFIq/PTK9ovb4lZAx
64U8L3Hh390xg1xHs2XI2N7dZww9JQRm8bxx+MwlZTosL0yzbYYzqxyx6mgirkJA
UjjcGQRnk8UWBy/NAENJYRbl2XZl49korWEaXDcLeBeGtUbDweavNc4kmH3FdQ/d
8Wf5WUhng8Ddd10yDd56RZx5WZ4XRjv/X1/uOLBfeDmcba4lRITVvQPMtKCbpQCF
5OSC484gHTdxKTXvQGt4mLXGCwI7Ekhm4BvaO5V3NPKolpjF1iLAw8IY5ZnODdq6
96HDht1BgA/ilUfZg7INnJQ1ZH3YzXNmhF6U6OFtO44q2BAFT1Iu8h15BogiH/qV
QpbnHGmYOh+awNI3sFqYH1Pcq7DcrkDbtYsW/e8B8mjirD9oQCgKU/a9/tVbLUwx
JOYGcqPh0fa+mz5TDsHQi4G2Lhd0qHg4JED0kGzUY3NPLf6o2pMI+kgFgxnWAtAI
giYTyCKB7qyzFvaj0cnAf+sNi8GSMP3dNxaarTj4pS5kB6LQ1tsr1vS3aYZH4IBt
oBdvmBqnuHr7C3p6QTtp4buCqE54ep9cx4drjbSwrwSzdWN1tWVZglT9xI/THXey
iDyWSlewWtPl4kSSSlHQTrZRGSdRRb8mXywL44iy14nzH11H5HgMydFfEF6K2Jn2
kAO03QTyUzPOpXD/R04WD3yFfaw1y+3mrwHSHy6vRecTEN+ASorqhFpqz0Kfm1ar
PH8QxAL+PlPBL3bSjKVBizePDpaD48D2gelRwXOAwehOzR9IRVZrYC0+Qq2Tpleh
6qqB0QHU6BK4woPUQaXpH0vqJRZ2/QweSk3NUAb3zk+lZ3SEoMRlES2K0f2tseNH
M7i5/m3Ld+Fs6xaJNvGZ00zaqJo3UsWX1nphOxlWQtonXwIa4fTZlJbMaaGzLT/8
2fJ/qpMozuuTigp0oFoqzJ4+IWU/F66Qj6ve0iOvaoJWvM1k08E2GgnP/mQXgnTH
SeXI5zi5z4Ubpo7uVBiUcSEckMciDsDAsgR/xzPvfoab2Qt7OCzNnAsPAY07HCaR
AaMSUFpqVBjPwdppB/0XNQvqiW4iMD/WViJOQ00POoUZ7euF34EkryebbTeEZeZv
fx97rUS263D4a4GAat2J+caEea/+vRw5SkooEBaR5vdxfyugo58XCOeupSykgz0G
TuklppxsTnPtc/bi0TURgn2/OBmYf/B5m/C3BeTxZvx1Q20U2xT6AtqogkVz6+Il
eIqm/IUz77/hY7LUheMxwvKNGUmx9qb49gIjbJXfV7tMFcrZm7KBOAicndeDp9i8
eGNM9Ln3bSEfCp72onijPgXOY6kwB/RPghSQ0pU/rgxGuQdSGHcXyBSkO19542cD
CHIBJ6wZqpGgUCjICN1PfsNU18Y/K8aWuHCisp5uKhbqTQDyS3vmih6OwxXy4lqb
DOY3cxZUrVSNymEFay8iZRc7Q0qtsqr1E5GgM8zr/4qlBBTOUBSU8Y47grHpM5y0
maau2yWTgh/mUlawFjeB6mMUEfgqh4mTnYFOutHCrGRlcWphtAa4AZQm5a02G79U
IXfbLEIVs8LKFnAhZdfNLDDIbx4kAbtUWdXzkGJ5nBuxzG1Rg/9obqDCi6o01HuM
tvFNA9wn5AJ+9JtLjEEPPbHyGei1AhffYQBUusZn4WnByOxKwbAt7SqPsxctA15+
nI4bQPn5LvRn1fTBXzUQjDiMWtYBXBvR9lVmE7ZBwUnlh187saxYNrRMKQ+OKdyI
2hvFx2Bzc7IYbEYfHSzSK6mc5fT7qzahpTp7TTLNSlSPXubvOqKA2srgalUImHTy
+dc6LijdCPpNefI66AAP8A1ctfeeS2Tte/kbedHQ0CSBya3MiIepdt+64XtF9qyV
Iwh78oJpOUfIDmsi+p8ysepcanqcqex1BdXLhkaQIEoaWppxlh4NNiq4gFSah1iY
yqsQiiar5Bsk2svoOlfpeVWFrb8TodIrS/SdvwDMj3wX2Us1dlLvKZcnBdiQC5i0
oxCCc1wqKhYofWbEgYzp4zI1Sf6WUPMXBv2FtEJdvxXWfk50SUNiPgCyid3s9UiS
dDdcAbqyV48Fjy+lsT4aiZpSDKsOeY2pSFWIbf3TgnU8fJGfkNQ7rN5AboEzSTfV
Vka3PCcq/KpPZfONw9Um3IGGjbZ9+5xSJ3miAOHYUrI6an2ouz5MJH6nyZeBvpHL
gYvHxP8nmrHuqJnMmSXNK4OSiJ7YQ7aNot8jLAALWGS1WOn/d31IvyT8EkzioKT7
msyyXgQCSu53y9ulmMRzP2/x2MOfd9XNLTCTL7QxanDyyDy27w019IlhJtg8I7bY
UVxQ5jv54Q30cmP3Dn3SFXd4bh+p6FTkLPUK6b0UfDlH8yriiDPMDZ/uBc2YSN3t
C4QhpW9GfRN4pBc+FEz2TXvUdm5kHnIvzrfw9hqEfhsHlsFTDuzxeEGP+YAD8awp
kvUUVL/qdeUWRQ+X2K1kwz7YZBFP82XEx0czAqnumrYUwTQXMcALIcOqBFYG/n2v
k43rdLHcIuSbjcdQI93JRnSATqxOsBp+83dXr1gQAmoORg+jkwN657lAVA+6UFH2
58fVo5efX0Oz6/hNSgzsWo2QQdZIoU7WZ77eUMPON32noXMD7719j+Tts7Nd3lxN
dh0tC8Zpaj9bGcbproZp3dNi1RkXI9jwJPKOQy0VHLZnHyJMWpTTPKpwCAGpyA/C
8V36H+eZKLYzvu5jC/CqyTLDZNroQx/nWcgvj6HZhdcADlZC+9L9fYu+pmzK2k+z
yx6XhOzcCARc0Csw8FkkOIYivOTSN2KOlpHdPgsq+t+k3o03ncCRUsqCXU43MARM
d219i2adlv+XINMxWsoy55HLZQ4F5gOOUdOi6Pq1iGXH23Pzodx8LFqHxcXLjhrY
kVzwGuyCC2+do6Pn704LG7/FsV/ROZweg+FzDRT8OKV8VCIxYATJAK4Hl8ixFFgm
TgEyem5qpk31Sv8fpA3q9UT4g8xu1obOWhd+rCJtSyEubcJJMN1atjMnf07EgMrk
2Rak8d0e4naizmSLfUU6fPXF3kkkI19Nw66rminRo8OeXGF41nC9VIMPQHFflEDC
OOn3v/GFR4QA7OuvM8iqZhwsqXrgLIBikhh+4cIbPdx1lQMEYfowXkkIwGy11R4p
u4cx+ZC5gLmWVRjVb/IzK3YtV5ixSqkpJrBirs+Rjalhp8bU+iQofPPSny3c6lSA
oA0mhqUCvKXTk+PrToZoGCe/CHpNSYMYXkv5GFPmDUfqKmynWI0PnGsYqSqKcVl4
2H1n3EED8d2C5BDwx49XDT4CJ/atHxJCdhQsOvbpwKoOVTqICsTZB8nZe/K2YAxH
gp/qqwc7pEAk4s03tTbpolOUI4AX6Ck4FhH0x594NngNzzXVbzFqnsq51sGTtRYq
BOfVWaBPk77O14Tk1Rkhsmj3fO5icx7QjJ9ZImryvl52oLAHsdZv80FA/LdiRzZr
rBY+uPpexDd2r9MYU5w0azy+XxX4ckr/WUD/3XkC8tZYmUiDMToTpC5pdb6Yb4py
+v17PL0jiq1n+RhcwHNxdSNvgPkpIo1FRzkvwF0ie6lKZtPVq0quAmnXurLdJM5k
D7Ut2GEAMbRJ7LFGl1DRJd1jqIohGPSAzA+ZZFHcjj2iba8WEyUv+zlQKWr2uzf0
s7flpxfNMKSEaVNLEVibPCg3HXTyGgtFWGd4cAQ+bQVE99dmWx9ocu6Si4nORdlh
cR3vrd1hGv6UsIcuc7m901n3SwZNYzgvj+kKlP47TvsgAHocO2uHl2ZQADnvEW2Y
ck9AB8iiCqvcd+T0aVZWujKJkAHvY4j3zqoywh+8RI13ecUBLuwwwckcuYbL7a41
QjivNhkzTkFBd2GMGYh5pM54x0v6wkIDZD52xx2gxMR1vmMgusirzpOzdRp1ind2
/JeETvlXD2j6prhVnn8ypej13DJ1nDlABjJ5VGS8eoAUbl3bxXgyg9Y3UA3sitwR
y0JzP6LDRP7R3nRnKO1iZA/dcm4WSk/TafEXdaEN9qzFOfCzJmXdQZiD4TqrUncq
6p8E9uZsyzh3K7VxoXPgCWSg7WUcl9LYbINyP42DyQTZ4IIeu4/V2/m3VeUaLuTa
8EP6gLlKiYwE+Hm6xR/gb58azQYRhOxgYSYP2mbkac48odmWGseTETet1XD/9ui4
vNtipT/3YOnOIL607bh6nc5dv6Nc28w2gRBHp+enJ1VJcYWfxAov+4nQq+wmLr9E
5Jt/5eaCSb3onLLwB8/kOVuUuz14Cf/WSH9rbQ3IuozlfYmmcj/mDG86a4bPrAIL
dnZ+/9FIe7P1cjJ3j1ohJKJ+8Sfx9CkMe94z3k9mPmzINmfyvwKS/lokSZ1SIOB8
RP0QJGQmnWooC1FW4aHaA47U2ycTh89yLK9jjS6TWOLvA50B5w5xY/khlfhQDfcM
LEqlcnROQEgr20X9SJs9Welkl7ESrMi2H13WbM+olxi89vc+0Qj4Fw4Hfs52eibo
ESqtvpmRlivOTTyCWd/CoF/cODpsfxpgMdjCt01wuWiyGmo4DoG7hWUu+7fWsLjL
6nj9pieXuUaJbgXYq4EW2BcbNYAYzmcxyKV8NWjFXGigVJdse8aNtDF8bMq/6jmv
PlxDIq8qghnAa+dUEXq1M3B5Zac/QmHQOL/fNbb6wj6Zu7qoaCX85uOh21hy3spU
ByTPKFKkozzi1ANlIdYZublZBONGO0duvHgad4Gs+FOxoWXGDO5mC4FxHteQPjwH
+R1AKpQgxZOMzYZZeAPDXYMzdKV/t2hRGgHh3ejVdRZPiCwqIfl/MX2lSsD1uluA
ONugzfzU0Vwpu1eVPZ0tZaLdMEY9qT0OYi56UydwIrGPK52V2K1fQ0LAaLc2bEOW
NWGNpPK3+ohZjUxRcITEzat6JeOJ7+KVyOteyaQM7LfCzj50dxZdzHp3QkxB1TsO
pZBV8jKjeY2C9ln86ZLacCOgH+8lpqwMmoLWs1EmXHbRp3rwE3IKuPgRQWRX1Z74
hfxM+xyQPt+HPjxa/R5RePMgxRrpPvBf1Kp3ericGlgVrbQ+hugaaDdBS5eJmK6k
ftwngZCsKq58kPCL5kM3Xoj7JlJoPNLSsFgjwQiZjZL2lB8vAs9zkf5Fvj7yiBCl
eidcOTRTVNGYmH0BJ8tO8fk8NfiWcM6P7XDZvbL9SM9+cMbYKZ9glLHVlV8otNxO
yttfXhRU4ZIVQpheZa/O9EMtan33dgWYz0AX+zomuqcgJNMW9KM5yiL2QQjqgT0y
UMM1bHq86ATVsDU5oFtjd/S4bPwOmfnr/ccYIbw7a07hAjM3mLorgYOKr7SB7us3
3SGKaZYvewx4WI+5R4PUT9+z7dIWMWZxTx25JCWS0GU1Hly7Qqe1Kok7qvva1+ZG
BRGYIcWUwrAu9SzK5eZCIPAt3tD2Zlf8TuVRspysVJjfSy+57v9uQhJEhdkWFz9y
4FKKNbIiaMM1/KClBIQnMIjKUCKNohELsSPmAZ2IdgqGqmwBP1tKlHbnvEsA/i3h
XZBpECuAMWPMnNrKa7o2LMh9pkO1IKM9gvo+w3JJlhaFckStH7bHzqkfwF0Kucnf
SOTQ6FOyi3t88cel16WAo+m9fuGKVbHSk1A1O3k0Ph9pEod+gpRbp6BkAn179odz
YCLiejXk70Hy6mCx7ChgrUjzjj0hRDTFbKrtHB2xWCW+7MbPvKsDmaSohwJnSpRC
hIPpe8uRNtM7GpTL6ZOUcVwbViNJQ+T4LM5bUq4P3DzNwTPu1KtrNMD+iR8iznWS
pvu0+pm+B5YtRdfeo8waPOFdqEbG0sMqZXOLhNIrszMKYGTYbQsnDPOnGsu06tGH
7mQRKAPI2tRpnrpO3nGUyW4ARIVv7aaY9x+LAik7m841QzMDC8pV2x6nzG69wVl0
sQYH6Wb8PBSOSqTgPRqNJgbMmjQ8I1BHmjMp/PHUPEAT8A8x8W9maWWlFKzEGl9o
LzYmbQNc1HyaEmPAsFq8E86ZvRf7+iUhDMzdH6uMe9FdxEQDRnszc8fdIhBd4GpF
bkl8WsZ7SlLClNnYoHO5PeKGKd4yxkcMs4+k2cAk1+P1HueTAmelIeQHEcrWEk+R
G02TE3Mr+OIcKnEFG3rA13cxpjrltqQvHxw5grdENHRZxkM+r8ep1Odkcxsjqp7W
MdbEO4oONRni4rRYcjfejFHYngbhwQ5wMod75DZ3yDBQTuhoSKtksNXB3WTqmYWi
7f5hPKw7YoQm7aT2Zy8YIpkEvrHDXrgkmZT3TSN/BnI9M9czZOcrX8l9pFsXBhM2
3Epu7hNbKLKvYiB+QbXU+GYnuwADUeTmqJ2dAkiJfboRR8FTanFmxA69NYRZf5oP
m3xCNaf8kZyUGheBSjhemAGcRE51nELbXp0/ND/euBv5/DUqnxdQnvc7fo8Qw7wY
FroB9eDBIvBPFu4P5TKyuqCTI1bLFIr/gLJJoLWVnU7JlWzTeISRkFV6BXsvua7D
sLxarNWxVtO7DCyXtoIVtsoDIZ/iWSrKtQC2/MozxjL/9qQHrUpkPsSfFw2coo4G
Z3nTE1dNrlumCYsDm6zlDCrySfqeINNRAcVmvJoXPdeCxL78A+h+i9GnKzVCW5yd
jVfM6PgF81RGGhWePXVSl4nkGnY+xCMetXam9I4dybE3sNTOBM0/GGXK+pWmfFu+
yI+THnQIgZPhSIyGl6Je72YW3C4CfrmH6vcMbt8o32vaXQkL3LDGlTPHtdQLCnQa
jzm5fDiqMYMYzYX8ncZpPFPuCn0Xlp1y2vE9zOBGsfgaGgPpqlXomUMbz0PWoo/p
fBGeCQUYsknaCfp/qGBGQcswCQEcXPLdrFUwULcah6NFtf1rSJQ9dEatJpCK9Lp1
ZrzUaqF+x4OjChHMQgweGoFhNfDoRr8ceSH1InIEQmvlnvbAiq/x8XUUOgZH/xib
73v4znApnLAIuyWCBilupBrs4Zt9TVn9c2p8oYFaaVg3kNQcrmbrZiv/mg4rGoqr
bPwgQeFwaZlBU0nAsEzaQkVkX1XQvnIWnfrgavUeByI9sWTG6frF8s5A4r0EqjuN
c7i2QT7kW4RKAweAuHrZSKjUXVxPF6vryqdXf3C7Xp+F3iWcDmfVBsqwZfGXW2W5
OgiQUHa7o6/AzOAHhvds0W+bnTw/pYCtpHZyB6cCUbl7RDCAucDANNOYuv5kUIsL
7IYM1WK1CGb3LB9riuG+YNP9SCcy9hfEMf8e93VrBh+BJmemKkUjw60FufDAvbdf
OjWT37I/IuVaNgW1UDwCilNmnHJH544KEgtAPGKC9vplRDYus1TU7XecJVo1t15Z
TnW/7C+YkH+rlbt0Iwt+Krzc4dITUK99VSKRPOz8eT6cDRHzHiiq0+PBaEtegyy0
0KKgTgdEWWqZaVZB9z0m1M2PXX78JOc9LN0vKXpTSdE4JGw1jOHgt67HY7vzLZGd
xx6taum5HgKzDwNtgWS9NzDTg4B7ybCAM5EW1pNsZs7OMr5aC+ILXfm6lGexb7wp
0MZt42VINDbf3tQBgBQS766toR706H3bcC4VDx0gm1807R8KcoHHhmskbnp3gfBE
nep00KZ9VZXBS//JM4ZikzFqx4to4LUWVpJubhZ+imwHVFgyUGDSudronn0QqnFr
3Z8zcds1UCzF+6TcMsvr78SFSLG6mT5LUeCcOUbNPj3cnP5aqdXGBS9A/CviNVg5
hu7JhQEddVNbSOfg6JkTgFb+VdO5DQ/HuQBCDq4JJNLxx00vi4hnBjifslV9zLNM
FlfDvprYpV/bxRi8GijZ3NlV7tJSJZFGVJJIsIsb7Fa7ojtENc/WOJC4iEWVDhMq
rzyajsJAasUk/yAe5r1R6AtF2SNTOPQVvOEjfIOT36UJXvAnbFl/k6ih6V6EHDvE
H2Zz4kHBLqlYWX3MRZxwRzseCMTiQZm8Xy4BZTg3UooVL5TZY4DKZlGr9/gLJh+m
spdE10yM/XOr6L2QAByk7r5KZOUga/kuomtzdMgJ7sQdnYTO7l7Nx5R6rtJWFHtl
1Hq1unqkbT6rVGORvXYCNu0lBgnTca+3NnY9ovuNKw4YD6OIe0L71t9k/ku1dUm4
jnR5Ci3/C7hdTXYkNkJxEUrP1/fKRRnN0DYvmz0ZI+tjP9Wl916opQrvxVVQ3793
DzJ9k98i9sqwwzDk/iZwBrsGVR8Vy7VDIVE88hH3cOc1JaiIbG+Kf67yjsqF/GRB
2tAy5OJKz3aE/DE6FmJqLtPeK8slP4R85aB1m7NeZ6+VFJWQSwmt6tUjFvx/vItc
GTmEZRiwsoXXlMFjD6+Q8igw1cL0/wRdcU/4SXrR4nCBTEVMdUdEK/lV9hy9SoQj
zUXB4GnoyRRpAWzx5UvfREFzwCt0mdXzNurbqLj+HGjClsFoqQeWU3hSjgHTjfzL
dkO/u7R8dzTFCri8VC7a36yRQV4f9bGH4bYAGD+gmyAh7e5hD0UMdRabE3vA0Zvk
kMSwScLkYlOdeqCvg2079j1+uVlfm3v7ZEPNSiG9xmTao490P/exr6iXXJFx9x3Z
+YTcPb01MN6DE+AVe2oJWavnr6Vx+ig/44p7gZIrwUUsYMY2MQ/5gMH67F4EyHA7
ly4UxF027cqKtN+qgYddDVZyPbHifC3SKWzWfQaVYkqZlPjSvYEkPw/IVD5szbeM
TkX/tF13psewsLzQNC/Gl45hZ0UwNiQc6eewTthjmDHykKGFtWr7KtHP7BM27jyU
/vfENmoJFo/ueoY91rVRB4MtUdlo8b9boLjciHPsQMYqaGpsGg897yKSP+PSMp3T
8oBWsRKTjp8uBhzzog+OboiGO8kMRMtgXB4yQ5kNAOupTywo24kkmbXZK9b7eXgC
rbORCwJrDgb17RV3hv0luvybLatCHM1DWHL+Xih3+e1XNknLLZfatyA37/uHWOZD
YSDAA1WS+71Jg2QZpxOAslOtCZqQOsXLHsI+kW5CBlpCqTSvoTtb51uR0AAwPrVu
oHXcQnYXN8brOK0ngyV8Pw6oi2dqmgviiJsN4ryUlwUeGzvf2LTdZP2AfhgAA5XM
NiLIG7OyuINCVNZTUufcgoajKomNSHVgIONZ32eZiTnLFpEN7wl7Bu+Y7/WxYBok
xEyROJFmVHdJ8sLYtOVqwdNSVYZlRMNpFWzcBvVkj6xQ9+qh1JGBLvVEZpmua5KW
sz53i2Ti1vCG0Rs4ABugmKBYcw6MoErR5oST9L7lRGtRCftW5L58tGO3uKxvU1mj
NnU4Z7MgMtTzlWGKJ+qJ01PWLrgVSXDdFOEq3rAoheHVWlUM9q7qjZvOG/WPvpNL
bXt/szOqFOzpPjvQK8ZAiVWr7dy5e1cauBDbWmcPUpqVGQOQ1XJgUoVmSMeAExxZ
6+j2b+W2wkMhR7fxgbVYUdUjHu3/8rBmNKndnWTHdxcuupFIlS27G2koJ0ATy3M5
3Zt0figQ6+jjZmfaF4uTCEv+fD7SDf9TQoIxNwebcJVr2gKI0Q9kvBhFmQwQUSmJ
RCMHFFSs1jIXBvvMsN4BHYzBUcYwC3kbyHjZQ0zqjBjo6g6N1aZqWSAtQhuSi14Z
gKJXL79YEX3X1DTSd2OXqZWN8yHwvHDOL2LKZ3AW86Xwi/wUQiXe/L6mlzeHL8F9
mrU3lI6Bnyb/prby9Uq9FBDoeQcELJJ8X/ilny2qxiDiBpbxF4fecvJWslC2ClZC
DHKNH0pRNnOjea3fUflmyj7y2nU/KXqX2zg888zChmflj4O5xGao202P0dHtlaHO
CWl03baRziJy/lrpGKCBI6HR1rDm0gi0jLQ6ah7sbjU1M9TfabzmbtUbJ3t4GlAd
W1YPuxtGnYvzpdl118bTWQha8Ulvezkdrrq1kwEfA2L3zm/4RnfzhGuV/0gQOsrS
fe4BVRGZKoSfvyVVjnQLXRFaGVMrfBud3SSRSAGbzQ3uik2z5uSUfYuzKtdePlmP
IHVJuAJEQeIOq442mJLrfHHTI9XlAMaYe18TBG0b5A6tAPeTtckWfqFyH0YR2IU3
l4kzfMAWlFYti7zPhQtOrxGDAyerx6eERBeVY/WIwMaEbsNkHEXvSNt6FyTPBe4T
D5wDPifsS+0Wq7TQ3ob0JF9on++P1vckKW0nP9J0qu+sQut4rhhQwUbeR0MW7Je+
UnNzg0mLRVoXhGckYZ5YqWYXYsJv1hA6w4lQ5jn9sCG8FM8otr3bab8yqG2qVtEr
Nc5tsb3IcP4iYhprK2i5RS22Q+ft2PphGU9RJf/wuwXA91HNu7Xu7PTyV94WIR6t
Mzozbqy7Rv/akwkSRqffAB1CkA/MBltJ479Txp59FoepCL5YdN/dJMiMwAopcpID
GbZANUIKKW8k6DI0LazSrSqqH5cYj9m/NTthmoxnT/isR3Y1W7NFOx1kf5WAg8VR
SKbUzY/UQYyAViNa+vlEb1BOCI8qhkvEA6RVcY9GYdVR+/ZHpLUInfVToJljkgF8
bpRrCXW5erUMI9eEaIgjuEiFFJ0IODNybcIRV5H9dWXhmXw+6T2AeN49J2u6f1Cu
BTCM+3nSlW7oVUIgUuoMERc+48GcgK4NFtw/E97f7pheb/5PKsdF+cMkdvtUL8KX
oouEmBSLCD7eDDgkS16pTKutDZDvQvmEK2LR/J3xUPG/8Ih2jfsWapcCh6XEmv5T
RLMFxeB2sFbIP5TjNVdS5ip25lUALsP8mstMClR6NcgfISefcStDygaz4YCPsX7+
ubmT+DAujWVjuI5Efxwlb0iMn1zrSEfwNsjwi7urUo18wTMpsrn4GscINdm7CuMB
hYg6AKybLIbXpG6D04llEL/Fa09Ww4iGbMai3xTPm4CQhq6RJStwdQBYhgIoKpDB
QUfmJYdh0388drsPCKzRrqkgm7/6vNkqhJ9WzED8WCJCQ7ThXkByN7Vxm1wLMd8u
pJfBwa4Ot16FVqQDvI6YqtqV81nXeXQU1ihKvMwpslofnZstcYnMbDfL5vmGKZ7X
S7gP8v8bkGEoq/njE1sGjguyAcZ7UzBAs5+8//1am/LSNEjFVskk5zcnNu/cYJyA
mGSQZTfcsVfJrsAtrshZ0MGn/FQwMevoldjMa0Y63XygJXEUYvPeVYEMg1R9vLPf
7PvCCh0gCesol0JVM6oPxPsPbq7VOMK9lUkC3Wi0tmN1/SBHAbq6BcyZ6uKfuagg
lJWuKWDFHeN9XRCyJrdpDeaVNMV7Dq8hpEKfe7lqSiBb3RZfbiPyEt9rnorfqb5R
nk7kETXrzD+0vQF0rn7Jo9GADopRELVJucPdoptE5BoA8EQ3mQHY+1SlnTo3Van7
bDxmiyahjT9Xo2Ire2CKmsMizvmUKgb2uyoih2xHzjgTWpS51/YHDI7kq+TXjvV5
1b1yEBeTkOEwZTW4rTMO2gfHHDbbjtIbCPeYNJ4kNsFyeIPaQrx3r2zPrtsuldJq
Gw3HCoAFmX/u6PF/8TyTTP7qIFxFqFVqEBakL+iSK5cLTS01jG87OtuYYwqgBSKV
BMT9dEZGfg4h570QAdU+dVtL744gP52LFMpuApNgQsqULqaK0gcyKwuOPLaAZTaa
h3yWYXFyT1GCiuEgnybDiWUF54CKae60Hce1BE37G+w5w7TBuaLBOG873Jlml0K8
BIjivMSmaLo62hWUdUCplfZ4rpv2Xheyof6ogbTEkUDcUEpO+Fj52lTfj5c1se5Y
0vdVb0og6hMn8Qxc7LaQC6Pp2swbQdHk51n3gcZ4d/mJcGBCjWeEOV/+PALtoxQA
ubFBuhwlsz4D4wGYuCBba8inw92u/MtnaLWRz0KAY/JzZP97K0sKYLCZI6fjyJOS
JHbwOf6iDOwgddQIZL/YYYmjuTSXr6bIR/krQPgKOZW2RvSKshL/FiKu+TeZfVVI
ffY9Rr7jazPlrPZz6M7UCjkk7U47+2+wS63mNPLcWKLqIVYXmS1FRzMcftfhYcF+
gQKBRYm6syuUXLnfYmy+dcoN74T4cx4cZwN8MBTndSdIbaurrpP03h6X+6n9P0nY
fkB3CDJwHO73Jpu32bkBhk+2KNOqpGN4bjhFMmgxD4hh6yYFCY6C6pie0R+ikoMZ
dBX+3Z6qGrTn4QGEa6SDWgJ1LQztBIwRiPGDINhiwTKqOdejNuiooI/COURNlS70
HiVHJ+KasYrSMDIJ+9U1JbqFtD5j5h+B5EihkXI7F7mkRYM19mtLqsjdPs4dx2aT
kmKdW/0eib1p40e1dObR6+AorF2zjqplWu03UVdJhsS/3HCxDzgj/wgyPmHAPzKB
phbrWKpB/YWH+WoR8ZMoUOHc2kHdK3J7auvbAnRBReZKspHwinlDS1L0prqpBKhu
AnV4C7GSLIGXnwATGI7tk4klAEt79yN/H8CT3RJA8+IOwi0yoBcyeiqswiLETnFb
ixOdHjY+tq0cqCmGXv//mUdQtkrN7LMfKLCNFsLqyTWfi0ljrQclETKgoDWRGSiz
B32wG+1lPFVKt4RXUPYlOIJt0I5BA4UOogqce8KZYDYxU33x8fZUycN+VJwd3ipp
n5ZaNug4EKZFkk2/ijL58NR3LnRLB5STiFUY2sFny7d6h+eJzIHZYRtWjEFw2A3/
Fn+K1DpZKA+KMA5eFCIwMFq0DWy5QinHPnD2kdVDU/34MyW2uh6XS5pTPOIXcr9Y
DQluXgi4Qo171xuN+PLq1I9IX6JAIptTZPzx0Siq3MxxNv9X4oC4BvSI9Lqc48dm
iop3pmMELdPPAvCRwXNYT4k3Ar/40ofuuOgDsPPGzesA8Q1fIqcF/1FvnE8unvzq
ghCt3wu3LzVN68fzChHyN8j0ye2XHoFoDPTYMRtPH2uhD2XHOJOIfhaY9tVtd3Ud
OSletgPm7X2pXuQiGnLsdHrxhVJfWm36nwlqe15wbh+zgzAvh2H8eYpu+nyJHSmx
Se9LmwLSi4te3cHmRnEL9b7FoV/eDFKhnA1UfxXm4HwMx2lqEaiNrqcHwLB3Ma5k
gr250DTAwcQf8miV1i8OKVXcqTTGtle07uAXYnNuJ/2nmHTIovOFhHVtCwsKaQr3
4SZcLPFp5n/Tjp7PeJ9drC01MkEvPojRvtEyMtpA6zHnBcX59IsyP1nsj/kJq7zd
lTsHgbCQosBO0py+TYn6tViB/Iwfn3c48Nw5ByF4ZLDgq51+AAV3zaccn/m8at6R
MhEdDHjHFU0d8M2GnJGyMx4Lv+dpY3zOTdIIx7BE8X78HG05zny0HSwJXhkn6iQs
XW7/phE8XT7uvIIbNc7+7S7Avbw/v56pYXYxLuDEViHocbO8znW5YG6gioDLNrrG
zORNYIq9Uf7NViG6OlX7ljoiWAmVFmlpZjv2TdrTkD0wXY49itFESYhTFhBfEQQB
pF2lvRUhtZxGjYoQX4iXjxpJvK/+xA3YnPzlP6W0KkenKECYlPhjnBNVq8qBLVuC
e4sP2JoeHqyW4nygfgBsmTKtYjpKTl6idI7Ek2yfkVSlM+Kakq1+0WBsYqoHr0KJ
1DTy01axLfGg065T/aw61jkAQfUDSFW8urUJ7ZkgZRgTNA9k/y3E7bFkMzH/6GAA
pmXJfjFwjL/wlVHetufK4iL1rFe2C2gdt0Hr4KayXHr8MlKSkeZozs8of8q+c3KW
E3RcRWkHV240hOS3nfiWqY5HvpBl8y3q8nuGBMe0UDM9iRxbo87MbzRaQLaNhol+
/M39Pa/IcCP01JwKtjLGgnFeyoOsBSjD7s1ZcKykJRSRRiFX+za7xuRaQzU7xvEg
YiMZOwymjj34M0kVpPfw6JmCPuyCRDCaQni34EiVM/5ZWpfSfJ2rTgQjPj2RGbV1
B4XYP6avbswvnkClIRNOxfhoVyPnlcENw2cfZHOI5sSf3ekKyDEtB6rCliwmmwdj
bF5Ng8dt0SEFC8F++PBQ50bmPDYyIhvGyp34LA9cs50J5oNKTf47djOrs1Fzb7av
pBsZMLl6BtGi7Y4EIB+UKKVTw2utC1znnHzzZIgpEpexLADEQv/p7UG1+t4jTUFz
fiUT2riVVArkC0haxRTsLtxeK95HRT+lTlCYjsmbJHLE8cKb0Sgv7XIirdp5Tsj7
L92c3c5HcusXKeI2PIBv67aqAFmH3uniFUPzrGNWc59xIcgeVHOd/tq41uqSm7uh
m8Ur5HudDOHDA/AJJxytVdr9b8qYVsf+V+fsY7locpWi8Ot/4tOQcEPi79ZhC4d8
zx0Eud5BFqHYO0wSaBbMJrMqQqcdkXmKMghAL8UZpC7QK2OVXsqugW1mZNhtWrA6
k6/5OdLOvBRcU8G2DR+IVw89iYsWhsLKeR/kfqj/pL4gOjQswnwl4dWta9Ib8Unk
rKqpOdeBRE8qw7XC8huQrffnFkNqgHJdjcyVVmdpPpPrIzuXCE/ZErUrMegT/Y5M
1Qy7UQhn5UyCt7WEoL+Ps50FMD8wDuMKcetzFFzay8q7yEGJD7p7AFqc0XizxPdE
XwNmxKxUfisUrqiVHlZ6DE/srDojZQlh0m/XUsf3zPOKvkhhVo3Sj0epf54+13pD
i2qiwPPnBslyTlTHT9u4MI028lrN+u8LivLCnDNZTJHWtL+iYCcrOT9/1CC/xyb+
oB5bmFp5JIHgdLb3gUAn24p3eA/bhGmTeXy8gnEkndraqndcH5qmn8ktmhE/nfSB
4r8NUodN143QUBTLO1jArIE7yVy+0qEBD6p3SRMnD1v3wl8EOfs9d2AvYtPZsV5Z
HTZPpMg20NoCDEetw0glQsCKavGEN9XarOXp7YAGxabVTkf7J+jpm8pDvsiUsb26
jtRSjuHDOfumTKrQwJkHg4yMRndnLHxTohrwoNiuBIfi+H/4wyAPlONwAwqct+0A
aC0CYAoJbUN7X/q0d9a0XBNqc8qEwdvTom+eGGvceB5GMc5Ii2PaN6IQvhutHfzG
OBVyBt225KgPDMg5rf/MZUBS6PmApqqI7aXy0HMqmgxRwTBCp2UuJukQ+q8qcfHm
wE1/tA4IeQA41VJSy1TXQdO72BHSyg9a3uesuZHu+7zLFH9g05HkQ1OCmnKcpf+H
Gf7Noo3XAEQV3aBO03nIFQEO7BWSH2eBq8WI+AaNfUdlPgpIhPxR3bWk9m4IYWne
UR4jqTYWxHt7ZzFqCsY3BeCyG9vYa49pKC8i5Az+rkz5UKGdVUSZjyeOIH0CTUqE
1v1gJrLlhhGPcT7h2czpt/jKtUNGmOgQ8A93OLmWP8SMWJF6dhAzdz4vdmAMjuiW
VShAYdPHEDk6SHLIfB2TpxdaxZ6Ddug8ft8CPtsdEHeLCOER4yMpLpAbHK5hnswJ
N/b08Z+YrTJjALHTq/J508HTZyHSR7xeo0QUkqutFLOgFezieMU4JEI1F+ROg8Oi
3JOj5AeYN6eqpdmM1gxx5kzX386X9uEbJWYH6tXdW/CAHpP1TuGMh0zzPecKLQN3
VOzQnungXDAf9iDPOJYq8BFe8BWyDDeaX7sjd53iP9OPdr8qjEKoMOMgP22TKwuF
cJIl3swjVq0eKaF7emvUhpiy1u7wWGlwmvjGbULmJUAxNfd0nsd8el3XgN8Ut9h8
2XSpNjD2co3y/SW0v4iQm54P9HBnsY45Ybhd9+PCA2hcBrx0zFj6okdlEMKS7Qpq
viE/T5GjwqOxQGvniHke13vV/UOrn1aDHOFlKPPT7dnB07GgxnsWaeev7PfJnif9
8IfS4p5tqZEWz++ma+vuEVozz7jWtN5N29nyJoevjBiyiTgcc5CE8do4Nv3f8Mfp
VLnhQhGEP07dGIVxJJ1zl33drCn9vFSQjDTrxq6oS3iWdh+vp9NFstmV87hfEEMB
DC6NgIInfqJ7jNuJ7FfhsrVkbqcQ+Z/PIVzp8eRob/M+nVguU3d99OJAU4VP0BEZ
6+39k92P1hW0hx/4I4v2AfHohmdM/cvkyYOILQLN+4bPeDdrqETdJslQHUPlvG1/
tqvZo8UX41I/Kx+kd2awft9fY2llCu2tCPHs3w0daEqygmOzsKkYIcUrDJ5NK0AY
KF0RoDw/Xi0w4k5I3WLsjR6Qwc+955hBGTOb3I/6xpZgFH84LuaWff4giVHah26X
HimroIGKVURp5pQS7XTSFZ4ujSFP3+8igSZXxHkw+HRAMoNtXQGhPE4wbi93TdMT
b32VnBRv714XZ4FJDCOdWk+3U1+RvM/V4Nx8jRqRbicRHl44Xhjf+ryTnlNItJc0
PynimoDU8sIPn04TD1lfz77/J0j3UXGnBktM5NrMXn1r34FWnxa/4ytgFDNEgxS6
7ylh7WVpkTZhTwSDiCRKUTnFi0Ce5QRTKmG2gjCV2Tc2hHjnUUNWLusjIxdBYhrX
yDuBnz88zArOLLXmfsYXLjbuuuGgO8vLqIQdE3f2yB4+HjjDc8fV1JRovUWENZ+Y
ik0D9azBj0gIrUXjox8O7cCXRXQIfXyl6Wr1XfFBU/tcO8UpiNhf7UlbFio8FsC/
WNDnWlUZY9kKEiY7Kj8HZIAYbkicxDcw/+09nGTLx8SMaWY3wO65VlGhGZM4MlfE
oYVmgdrGFJaXUeBN+Gjyzml00id99/tALBghlCBKdyjEBgLGHqBxhkyK1V/SBkqs
/z/FJLaBs2nGUJUP/YSpEJKHzYU1oV8X9fnDP84iOK2zJAuHQ+myavx4fMqVV4rg
pnpzTwk1pCJ9SkDavtzK6h13T3rsqIBRGmLKl+4SdAo+oYUnCrliwYZjVIad2nKy
1in4sIA1jf6+5PIx0oiYV/xchZyxzzCUtzSpad3GGifwkBkZh2vLBrlEfE1PucZW
sQ7gAhgkqNJBBo/gGLIJOtygItjDsz00vFc4OtKEipwsZ7gd7bJxeNKzut8Y3QMx
UrZoTAf0HhlxvyZUo9RPQ3/hBrLkDgJn18SUGRfJ+xtUfuUNj+itwq+ny43jF00J
gErG5GXWnJ03dfqrSFGn+nxS/+8todhTGsa5Ddpo346jsIcVG+hklzz4BcuUXS1u
y0e73bBL3Jl5adaTQn+mBSQ8ZAdsf5L9ah8x4xQuRUxu5Fv3pY0G0C6UPpt0N8PL
IgTyDk8af0CZqUK5eC6Gqm7mCKLuRyXB6dRGcmKULVlLfwj+mQuNh4Z1hBB3rTt9
zp28kviOjw0Zy1IF+jXsriwCONZO4KHkY8gbz47xyKCg6DiUjdYvrhBpZk/fYw9j
TLTmUJS2vKMrRSXeee448xo9nGmuZXfp3hr3JiTSR9iDNQccW8bIM3nqpyEP3Nd5
Gdw2p8AXvJpN9EvfXSjJIk5vRiBEZMXTjA+C8Jcmba/xFRHXeNjntAYrzkTkEV1j
UzdtCZp+vKfQS6ZxCZ7+B1CzrNAI2WRem5sPQkObs/JCI4b4MA7k7xJyElYVpyKx
PebCTB8G50DdQNylB/VsC5S6hthBqTRklI0F0oUUEcnz7IVaUn8q9MYQxN6ATLI7
YEp9wYFe9UDt5/h0vNKLsrW92UrlTbsR+BdKnoEn1gr9o+qLCi7v+OIywV+WRDs/
acUXUuWYlfQotiumNBlUum0WIhpa5iCxN83rlINtQ9h6RvesX6Qp8OPT8ImSgRpX
wAxnQ/n7dsaR9Vm3KkDiQ/INTSfGZDpaDayFJkNOA3R/t8g6UYQzPqwtNN8WhWJP
zvHxDWGUU8A9P2+oaTrDbBSh7Vvqcv+YM0CY1Fx961pJvXpQaXXXfaDDuuvB9s3k
Zk4I3J6XrP2Mv4+7P9jEMISmPj8jVzxyvizRh93OtyLEq13EqrX+qzj3bjBEDhan
qKL1J0ZB1WkgGcMXiUsJUZV30buBcffr3Ut7xqzEtrYq5Gg0M/5hlWN+dNCTNnXp
hVDB+1TzkmMGfUPxtrtEzMKIb1PLdhPIWRC/6AX/RCccNSa4ZKH+yDtdNwfWQZVt
VSuEYgPOn+Qohf0uaXCQ0EVmOoeMtBua8Zwd1oeQU7X6biDhjIBOQberGOrRV3Gk
JEJp/CHLLDskcvXnYbSq+zk9Vn0Rvp4UpNDByj9Hr246c2/D+j0w2d2+92q/sKLz
nWUp+a+rcCWmCwDSRm0pLwF0EvIJyOddTe+kztIxbWsZCFM/A3VAJmT5/ZFQtPHs
Wo4VI6/UPb/9xh/GkSEIU2Yghb4JlaKjSgZn2vMSOQxyvESlpIHvF0iJND1eO0Xb
0K9gOfttpikzQm4ZZy+qA7Ed8oYV9WBRs/944CCZsbfF+6yVPguFXifCQHoZLn2G
rsuoCd3DWQex6tiHkc0GS5mPdo8FNjUz2qeY9QZi7ES3nTt/jE7jdzfbqPl4DyUh
YgS9YsXRFiMJYnXA4WySb7jZvh9If1svhpAXKMh+ZTAWgLi3JftlCEH4l/b3fhAX
WSPWCFtwrWfSRtReKeTjQsEY1jBsf7+nVG/0T4PjCMKsqjyMD/xzwi8h6rEBHRLQ
q1FQGWSl9JdZZIVl1HwFxKQRNgZzaP3ay1E1YHPriwXDT9aeK6YDbptTJsEmmjQy
gdh4aLBAsaU90rlmWxYeRqjaYtgEVFCI6su26i1lxg34XXp8u8IjYBat1BawMScf
wgE4bl8v7R/Abqqtr2YVBZZPYk/cCCvrLaDPkIpz9FMF6SP8UAzcA7BiOHFuVFFQ
uL3RnzZTUNINyaKmBbM2dWqt6wHlszktBo8CRYmPAsGyRepHJ66QeYzaMogC31JB
/S+zAYnEPmdXpePFpvQZuaQnHxm4irnRcEA5ax29ci7Yp3NhvksPd09ADjlIBvd0
pMbrNkfK0zcP8KvchFmJUhVquL8tAyLZVr7QSNDiVlPPEkDZ3T+NBUu/bqtBAcZi
Ine8UjudWyRKnOtv2fmFV/8nSvW8d5ZfZ7+vEAJdY/UNsCps/I6AB1RRBRQFjVpS
Y4iB81BV/MNASAzgHA8R3WKOCXvaaHkDhLI7ihApZjUc9/vylyP0PTIO5rF7Q8Vo
Nvg0SR2s+xS1ytTLGtaGSGoVauU4LwvcSqcuXNmqpIXhF9EOXJSM9LPHw0bJsLau
hVx9BxBkH9kwvJP1ryD6H501CzphAiZucZ/v/JTv2z0rNUp+jpXflYHWOsVOqSko
l8pB66+wlZOEvKOq2DY1hZmJ17b5puwjyyD6w7y5kIZPrSaVbCEaRiFNaIYYKzb5
wxoGYKy5buMZmSOs/5dZfZ7+GwiyQGr/2NMDExwKoXtxKMTD+qXSVzyQaJTrM5tR
Vn87Qr5z055LD3zTGFi0rBAvayV+ratNnIEEc1K1aC+oep7CcgETF0KwlaXBn3zX
SrBlDjoBajau90hY4l1f45D8SLsJpTMOLYbF9j0MFj9reNkCO5lxMpSew16DmYw0
rYktixV53vyEBC+TVm1Z1V4mu9ghAxNhqULI8Ueg2R71bQ4ODBa1W2QKNQ0S435e
KJHIanX+GucvnfHVAU3JyrNo+hkXPS5EgwLXSYOqHQhFnOLWANhiYUQ2IQNDnTQp
1dhxoiOCBRf46NNRg8SCHe3T7X6o60otJ16QorCmwfrsjOXjkWNIGlI6MsQFxpmI
WsMceuNyPH0mIWjcHafCrb3tneCuKrZW50t6UgSxMSjUZYoFGFE6Q1IEfxHJtrRj
zMfk+3JC4aX6gsyMlmzeuNhbwJho2dcWj5ngVHw+iBBeJCiDsbk1D6FvJOgBwi9+
wG3Aqj+Ie4j6Zht1bpGYh1SVwz71ww9jJYG/aNTkICq1Q0x6g3RVwNC4AgPPaJQ4
fLygs/o4XQYOwqPTUhiNQxNJnK2PsHjiyUJNXKA+Up3Db9dMkBsipBQZcIQKNNL6
6mHdkzoZM+41qeyqbUTlUboz7VuCfqcZ+wRF4EYmP1GIXc+yln5rlNL2ppB0caBZ
vz82p4F2a20iD6KCKAS3laBFVFJOaF6rpMNVGUlBr809lMtQUp5WH8wQ2NWxfTiW
Wml5eYHusSRySdUffYmbBOgzlvPLjeq5DmJ4evXy/7JA70ixXY/9+GsLvXOIaSyU
HuacR5hyCN2uqMPHKdwYEd7dVJjQ0q4ssA+klSbHL+Dm4SMEZ/4ChBYNpQu77uoc
s76VrXZjwTTz+tJbtfL+Bo3Yhp35XW0IG20BnVqOZ6wg4hHD0UGL/rUIFRiK62p5
Qt0uA/PEcHO0wvrcx5/XNg3kCYR3PMOVRAIkLF1Z23vf45JJAw5hVoHvtj/swXXz
/F1d7T2OLVfeJpEDnvQv/lqpzrXO1VBuArSx50NRw8+AFPXPONREotnsIdpWvRB1
KeqEEnZuzd900UvdAtMtg3gD5cUyiilb8WXAELXEYG1IANLhuHHY5I2TEJfY4aWI
Pbke9+vHe3UT0FOedcydS31TyChcfJz+Kb4CFFCNoVK9JuCclcEAvwHVGxYBPuw7
2gT7HETlEEdx9XKMnJnk+oU0Es/fFEb7JpJREzbZVWW9m/A6NWvuRJ+pV5gpdKBa
yCkPF+ikUNECQZ1yeKtcfgRYu10vXzZnj/vMLw9QKM48mkECWg5d1e1XiyFUdMvt
ZbdxL1eI87txR3rNTo64XP+edbdnJfE29zvk41ugKvz5AH8M73ABG00+gsVYi+Ay
eI3goh40Xb6B4tbm4DgHlaf81UuB5KpGyVnO0yNipFpo93sFgEpRV7f3VXU8/65d
BuHv7pwtmNtpKnxmEaVw6L1jtYwWwYirEJrugLdPp2jjHfGMX27urPXCUt2e/b4z
/sKW2EmNhtbf1b8q6WrmtUaLP/5Tsfu4MYWiKI4a9z7rBwSE08gUZnbXkwrTu6J/
dQ0reSFrZpE3cfSTsO7LJjRMIn/9fymOrY3Hj+553J5dOgQJqvLsBveBTeeAWVJE
XmzqF59Jc4T2Zlu2Fm9lhdvTfejvQ/QD1eIuAArB245oq3N5IvhCfjD31igQAwXa
PPsty4pd1nMvIW/SoOuVTubeqNyf6ClPG41SSjwPtJB+flF4UE/xCQSU4typcwlZ
4Jcbf8JXuG62lV9mPAjYI0zGNDobN+ZSYXHM+Sugeoi52zy1zeaaoFqZOaNMsq53
ACIzzoCpi7AGcIOyHwRFxU4q5Xuv5zdsQT/k4954sxGjo2XYdtD4JZbtADMZwtdm
0SH4NJwdIe/9ExCQ6srYFYat8ZRiGhhii6iC7axogAARxEqjUO59OcwmIOKpKBGS
tECtoMJlZXW7ahfG0JDy/nVYLJAcuW0bqQTk3cdnW0mZygcj3CEVHg+ZfFqCEpf0
I/rJ7Aj9X+TN3OcK6/JeyOQehCvEATy6rviAPsoADIv2i7AqcyKz0SVwqg0cFUx6
uOblegVSDcEt+FKyd40oMl5rowYeC1Iw/CvU8UeCIiCebZrac+WzSEn7th23NFZO
kCOXWJ44XGfY8L79d/ZzUIcaN09zws80yr85qzCRCgodjXgXFFCKQqKa05clgnlP
nJxE9GBCf5N85r1T2eiwI+EDu7a10vsZbXFaZJ25VNV91eQaue/OkV4z9tsPrvX+
UoDF6jjBT9oPJ9xAUWztDjH2l8E4RswKMSDojGq/eknQdlCXNlxbMuhBuxq8DAi8
LuB86VdRF/yOdVSu9ySHpi6mWUeG+wrQoxTKfnOtMsCUi3XxMGnO6SrGmWV0/vLy
XujS951mILB5UIK2o+W6SKNtyClnf3ue8aphoXg4G6815Rq92wlpsOPnJV1/tRzi
75J2adUS4dUOrH8pOtq62JVcLUoLtNqwzC2cTqZT8sn6kXcK5JbPIoQVnYlDUj4+
C7TVppF+xgjDBg7GbujXJ03naI4TxpXRGILNLAMREcl8XcFSBHKa9qM7nxwSpMVi
WvLRNEURIKTcHg78HmsymqZjL1Vbb01zlnTBdo5USc+8cFS0gEuDMWMCj0pxLiLJ
DLfrAa9U3iDMJDRNmUgbhs6z40gY62k8ky2u+cKg/O8wrf/AUg9VjywXdZjmLtRf
ys8k7UGnyeIsDj9620YfdSJw5NXwZWpP9GBz/47ZOm16DtkF3qRcykCqnthLfuwQ
3F247HZ7lLsVjf57y8QheZ4TTJLN5zT7p1a46aRiHzs0zg38/m0SXDjU5Bks/UcY
gsaldpT+ZMNptNmOrPF0nqdjyZh2rkAKc/DuvF5cO1bnHkMbp5p3Kdn2042RAW9l
t/5EEq43EWf/wmCfvAlGUz8miiF1KvHOvgIz6/U6Vh1PMJc4UY1p4nPg1Zn9s9oG
ZvrpNzpKWDKgFn3R4xF7eZWOfj4hHv9ZBtKXZiscxOV7+8DurDeLCIh0jxOdoC89
xnn//bvIBgMB1Xf1b29oTU1B8JIckBtD89bmAhzBUhN99A9ZPKKRtRz1kVj6hDnf
rvq1KXo5MFhM1NDLPaRQb2//ApGDFavgVBC//3aD46T9ZFMweE8anLb/Qxw5hpfQ
5xQ3SQ83NlL+AFoaXGKzwm7KW+p+Spk2hq27ySzS0QgeGOmYB9U2fmlApNM9lRZ/
EVFID/4FQ8DaMtRCsv6MeX1CEIYCnrRRwmMzf3WXokkKaRMqD2ogP59QcAwsfuOY
ZF3i9Znt9800bnqO+y8uYmsTTIJU9je0cAkLG9XDHuNC1uUb1i+A97Ug96mwnkeL
4BqkEGhxizyL8Tpf0BF3/827Wtf5gfuHJrZglGEHMnXeCEdIuMziHNJL1X01jPig
RNDbtGju4DoECtEUb4/nmMVBNJrsAkj7/hneQyLZKkZ8EVwYUGPoenfGQaocLUkp
ZN8xcDBXvybJYE1SzN1HLodqrIzq+uTWH2P+s86jY5dXzBhM+Ch+bVvFOsB0+Lde
cR/ageTyX4juQF9DiPW/r7jztd8kjnp1/iRIJQpeLsoXK6m6AAyfLz4Ll10C804f
7rOp56llm1dspxfd+r0T++WMV5pw90IB8vb6bby3FdTR+yrMsX5YC520rS1cVVFw
EeBqcHqIjCc3Mzf1gkW04Uj/tX1Yc05jwjkKwooNd9zZpciOQ4kOOwB8+ZFnVw3A
MG5FOSsVm9/2s6DCDQVljiDBCMgePlwYADl2plgCyUxRDqdUEwB68xTkSsxRYpJp
0FBNw0xhZBqyii51unrwA2aNc/3aS0Oc46fdCFh1ugq7P1a7yL85jMqlH6XoF8HY
HdkD/+u77KPfaTQQPzF5J/F3s2dek9r3wLsbYtcXc4zGDNhAfO2DciBFt28yoMQR
kPVKR26RIZM/z+Y+YCSfNReZVFeKl7VsTfIc63MRDt1vUC1GrAE71zgT7ka2EBWs
BBBuoAUHzwP2VSbJLONHNTdbs2lrNc79OMAjlETnfBGDyXjk2SC1HjVE/GmAVs5q
K0UlbBveuFR6R2mpkFQIIE8Z+UF4aEK7EF2z/Lt68775l1S10ipcW5NxQUbPEz7B
9qokPegCjVhJxBaEdI7SuZ7wZ0jNeAtUcuuiplER2vQdzecS6Fy9so28efr1ZeVB
WJtxlIbuQOP0O+0JBXi9hX/YIGCdKxwYcDccuTGhkZfkeY1LL0lQIpIVJ9hCj9nR
ipAv4D/jbI9Lm3qcs/hYvZWUB2NdqebOeXa0zP8mZC4ebsn/ibU7tb3OMOSqCtTq
/wxJ1Va6ZwkqVHgNiYBufax6BA/d/wJr2If3q1wCehWDTn6Pgfy8TwtnE9jPTdpv
VRytcJWG3nFmPsE8JouWbSnI6S3B9wP/OP04r3HmCYkx7r0vMFqKASXJngJ14FBu
3WxaUctA+Fh1hbRBgbOD5pD/ldV1Aq5Mz4Epzqolhj9FOGb7FHlwhnhIM26US99R
a/B6Ux+97fG9X1JWB0bEQIjwy+TMgAWAvgGVALBUQ+kZGA6QxM0x+WabOviQ4Dwy
TxhC2fX/SEUjYwE0uET+wOzlRhrfGFWPzsQPnkRZv4YGsVeSkORo+vtRzbimCI6U
isWdI9ILEF/S54AmNK69Ii9Fx5P5bPFZ6BMoUe388IuDD9kdSQKDEGqTjiPeeI2M
t//32th1zKe+FYRD868TxNueahVWwMDdUtzuPoaUiROifrYfbpioshparJGd6LmT
Y24gNraQS0D2HJIw9ciji4iSBCyU6mM2qSP1vP+C6nAM0tlYSnwxGwTsKAC78rpy
ihax8Fc9fFhcZEFebvluaSoC8UvOZwY3HllOkh0QYMvGm5o4cHv2PXXAPaftWKbu
K70etGAOZdh/DYDZETWeVc6Ge68IjmdlIbgTg21ovibWbU3IoeVcDlMnL6VRlRZ/
TR3Pv9BUHwVYY7942n2RNgZ0E4K80cZDYxBrMlU/Es55Qs+EAvc584SPi+ExWnQz
+PZHc1vQlHfaSxi57Gx4VtQa3pTK2yT9+yE1aGbRArvRRW4QoFI7TEsYaQc0lHil
oX6Cm4wulrKKcgovuBUw98vq6ZQYK3CeDk0Ybaa1vIyGlilpGyKcquP5MrSrRafJ
JDwBCEjFdNrrisY6+7U9R1ELa79mJUZsWT1WazMeUGserW1Cknyts9m3p7TWm2lb
b+DJ5CWTWXSvonyyEyqFk6RB5FZXxxOwp9UPcAXbKwg0WSMR8RH7OZHyfIRa+1/4
hjWKO9yIubRHazkXC3WyEgOjRxzFE8aLLGMkVOjsAMk7ttLy93arD+dZ489+mnB3
YMOPmyHJBL14mBYeL+/zngCQsDe3Bs6rtTxiUdcOojm/OJMVhMAG8TAKaKbvB7e4
jPGfubbEf0/UStVcbCX7+MU0NHxGAPL5gS6nl5ul2EHl7QxwZ9992XQ04mY/2aUz
MgZJt81FnZfVvbX/ziT6DSD7Caza05K8GDci5wQ4ol6kh7FWhy3R0+8WOxRVUMVQ
Ijlr1OthmdES3HknMfAZur7JCWbiGRyJ4qgp5vG5Uiaf78YV6i4vFt7FJKBAv1W8
QqC9fmdXivpv4lDsJb1jyKlwUaE/ul+OValyP7UIAdrc53HuMzER4xzH1gul4I00
T4fcxMAW6CkDOVlgSGtTZljLWJRlsDtVsTcN4yBedqiD+CY9E861RqO9IvILemuy
+vP8orrmYvO3nE3Wv6sYnJSWwR19GekVzwV3UsDBYLT5Y82Z13+oAZtglZtQ5dOc
YR1Bjyws5njxQu3NBq4+8/pCxazUnG0rSW3AKBjT95MpIgPAnKsstM1WJUoUtIR8
T/yzS6nsQ2K8Z1pe1Xl/EaymBcIzu226+W73IrdXv1sqSdI8a9snXVwOZuCrFqGH
YfnIJ7+zqw7DUOYXVdwJF1U8pB8aAxsvucYUeJLrWarKBKtPs5PaSCsUZQmopdT/
Z5RkDHpk0OQS1PwI9lo2k6OaJ5aKCBS4JHjt62HfMR9He1INEmE6EfpNv1hW6yTH
rCrbfpPBnDqT8wUWy1cFMw5jFAILhWEmzGSquSeixQPfnRHZjQJFy4GQk5NIU0f4
MtDDtp+SAHCiKGcfaoMxRtUOySA+5VY3kfOPc3lhAXf9rNoNOat1DslgT4UmfhwS
PhhmGrIRlM2RxwYMaBOW3od+pXJKuF+n/4FVwsAsAUfOahyzTuz2rDXRDFarrM/2
2BMRKf4GZRyO19CBWhPD2G3hIQYPv8n3rGBYn2U0kazPSXJZnMmDOcVUDGBMbg8G
aw6KcrZ8z7xyW02+fHZw/Qev2ENIlMfRjO1q6EkgpAUv2cOtee8R0oFqekG+cpV9
/d/ot3hEp2GiLIP8L60e7XT/CxH0Jf6bGo7AfBotiGon5DOT8nnZTF9MOW8/VBIM
wuC/EnRsCa7d8d29Ke01L7AYjpdigR7fLosDXMw/d7pJT3uWQ/G4w2eDrfx28Mlz
l/J6cE7xHYlJkWcfI1gZOnlQJMlArgiTnAvZjTwRjsHpqZTNNgBk34L8aJ2EMMo4
DON7UxDcTVd0QhHk0md9ldjzfLC3jsm/j5htY2LLq5CbOwY4U04aNouIVnLro5xW
sQPYYhu/G68I5oNdh+pNG7sGCoRnC8cwtNvdJIRTIDYSE57pk/qcPWRJ03h980eA
akuFBZLvO/OS8Mb9P/aXg7DtNQjGj+Nr9raDzXwlMautnuPPRAaQMhIeI4+RM2+M
P7WiWhCw6VU+CTkkrii1urjoZ9eZH61T4Q/gye9nZoCIyzv1+bEYB4NVkaS3ow/L
6GOYtQS050acilo0HaCBN8MzZber1MFStQIqfdV7A6Z9kDMmzrMGsZWFCM/vLrf2
wGNexKEgaKPTuHyxvWp0A73VGA/8vCbUc/XlAFRUCVvrWJyDVTa3PjEYnhNSs1XK
OmvhIPrUyoY4IeLhHmseO54sa2u0LT/jZyejsJhhfGD4NvmqqoPLkO0dB1bkaeQO
g7HmsNSLJmO1Yz2HwrHh4XKn61L0pIeGo6iQRJyvi+XFqo7T6tYFRb3dW14fbbz+
4qZGzyu/wVv2CUqBjVY79m6EOPmS/huc/pApuZLWuaWlME1swlX1aY5aojWtVKV4
FxPcn+Blekw00Vu7G8mp0Ache5GEtOJIPU5TiqpNkNstaFwk4VfRT76l0EUujZrJ
AyUebXWZgSn33KxFWrWcMpZJQxY3nYsxtRHJDjJdnD8s8QZ/eI3R+b6lb1bq/GWJ
Sz6O+05mxu4prsc7Fep1mwqbVfmoI64jyFoAijXDfaTPmE97H+Nk78c0eh2X41IH
BQx1SrxvM1BMWp//WLB0G6abRXHyUt+pB7N8ttHcBrJdqFZy08tQ10ScbTxjP5+e
damCGHhpW+EOCoj/vofDRsb9tJvTxVGIId8diuJcSs6WBOqwV2gNLU3cbY38FV8Q
zr3JMsemknoAbJ/cHpDsT5zSIUf/SgPTXI4GyfEDRoBU5Z5AQhhZgtc+uh2M4tcm
rStjjT6PBEwWmsYoQuoEIkddw3k5xaPRW2lpOqiwNItEnDwmGRxuFbW4hyOCerhm
Ycf17NRwba568cgWdHp0woCDBsU1A8vxLkuYTqqFHWxjg8iH84lMC8SKh9hSUo9h
vaPDToYUk+DaE8CNDbpZ8xamRyqzNnikunQ0MOEaTpSVB/z4RR3TRuhsjPnLYSgL
g7ZYl2hFdg38xWsPJb5HdJkpzfLsJi0ovzj9SbufS4qViht4PAtdQ+DiLJiJCiHX
e6ujJEB61PYyrp1DqihXAcf8UvRomgN5kAH0yWzDgTN1GZXIXpjALqm0gBd0PCan
NgaiawtHEdJGbp4LOvtRXtJekH96TBzfQqsWjPHKVUvzo335iFBVnVZjzIEO8V8k
WVxE0TgWIvG5C79hBKRiHCvD32+J/L2rg5at1gS9NCOoEyvi+Kpc80/B2mGS7ScB
Ysgw5Xh/Qf8Z7TySM7PHNEpT+enESstsireO0RY0N/AFbCDZWVgwsWDhw0lsz/hW
V/x+Q5xrNJ93OP8wU40A04jO4mfIonr3rLOluPUfSNnl6kL6WYc+WBMjl5MOGJ0S
qyHldCRMbNfMethW1hXTPbO12dBRB2m9eezDN6778jUE5cY0Dv0WfvLTgGWhXlMS
t5GMhd2MgYD59IMk0qD5WalP/x6ud8Jn6i94aHCtGRGRffdIByjlpCRYsbIQmSOd
70eRcVkZu+jK3gKpEbks6U/WZI/U/GsI0vWKNgHMwMXetR2ObrmvB1UCpEEk1PDn
5FbSmEBEydtv+EbBHHJEJ7oYigrkuDCnPHQ45vM4iCsgqwGMe7V9ah4Et6tx3Kjc
O0ENcbtP2+mieT0rjVr1ciIW78h7efHOz7ucEIQ427DgncogdSMNeOUhyPme3u4s
Ce9RHgHEAgC7Uw+VXqhDWVVfXa4+MzTc/KB8GGvCCYecV8oNC0TvWyUeBXI/Mlot
Kz10EpCCKfF0DMN8p0+D2pH4or2rYexXBwcSSFsg7Ny1EdGBbK6iNmgKdrHejpr1
4c7J7eztQa4zxs7Yk5/vToszXbvVKdKiqQ6VUoNqUtSSWAvdl2Q+lziQmy53dGc7
naACj1LMDX4/Zr4i0rTJISKkxQ2Oc40350WV0rD7WbPJIzPkcxeP2u8sXukkoJfK
2NF7enAG0Nk2F+mCe+RvIN83/9RQjPrH/pTxZilBJUz1+XpDjzhVZCwnI2O06zd+
ODxw6AXJsoTHdUxKrZ8EbM1GMVkFwGUg2YvQ1+8Ur9PNwG117EuKSEZfiOAzgGVC
YZSBBxCBLIu8aHhNhY2de2zEnOH/m5R4WO4Kd0XWY+nffv9lBXNXK8iZyWJuKKCR
uMcn6hiSrbeyR96BHs8Re+qjnQFSMNqdaroPGGobzxS95A/Z9ZKwQ+Il16HsDKOE
p92rAUr0dSNab0TyMW0ujdOPOzyZadqcUbNJOzW/f63jF/LSgJ0Kd+ybKc3L3HbI
3rpjZNoHb5PaX9KrU285S7J6P4gThqb10+WIDipDYKBaerWphJtv9v3xHqPZAyc7
yf7ub/gb28WqBaNFuK7o1We11vPR5AD4/KSmeB5H5jLiglON/Radz3KmtDSF2VJW
c3KbWMjnyHajTwumW0ka+q7UKmsjMacQwF5jliCeKE+cckw4MwUs4MM2vdD+GCVk
bjfY7hIY+edFBfFHKT+pm3zNSIQ/edfXJcV4RvbM/OsfyREbuxOeLgP0qXI6euGb
sMSkTyK3njin5SgCZ8A3bG5elr22V9s9594bi/FPQwfyhZ+glQHGAxQkCyUiBcyF
/WCK6x8F3OZ0AIGv9E7DpiFjiIko/AwiFJ7WammemSaJ0TYqStZecknw0U6jlw4B
Ny3spChSTKjRB5Mha+PGdvmjGm1xiMPOP5UikQw/b2brWX1hbY7I6jf8XFPZ4M6g
lPCaZUSk7I75jMN4KdlUpWtyGIyiAvXNCd7UymP33d4DgEbTivYCDHYEZdml1GJw
I8dZFSffe12/8wkBdt0SB+q859B5FPVDS6anJ8I21SM0a/N0HTpOn2sAjvZfvOgx
kPlcd4zHJu/ZtcBxUNGqIKRkYbD5tN3Brk3B29Gxzke31B3kZjou492VNcwXjImb
YfAU0veM0CJNNmlqnuiGyAjKeRLytUKfozeLIAxiSRKGMNvas2zd8PbuwFJ8uWyG
Vlly9qwL+l7LwFjkLkJyQVy6H70iQAzz2snwx+EHfQ7Y1U4Yyr4FsYcDzj6GjBV+
GUcHOtHg/ZKiKp17/In4KXMVDHJc53fPpodiLJxeQAR+8mbamJARwwtSOxuO6THT
CzU145bfQrmnlzgwL67EcVfhhtBTLtf3f7UrMStl7T5TBBOwa0+jHwBvhYZU5167
RxuNValJkDjKDPSwYBC61VmyzR9Ycqq2smhJ7Hd19TMh3uJITIWf3X59QQ/tqhm2
TJU+TcJkH9q4Bzdy3ChizzzZ6w1uB3BFWtuLINQXEbOpJVlzQnOGge9ovpu5W3bA
hWmhTpNzRSiC9X1Xt4s2vgP+SkiapIpP/ItWnlKiDzOxnVz/nQLij+5mzcg8Qp3J
JUXegEMMdRmC6g179IRkq6mi3/Bqnm0zx74xn9DG+t46SswFP9Y09RXhYeRbl51/
auv5stQCoqEaS14p/y07jmprm8QZXRNKu8j+wUQEsB1Rwzora0w6jTTC+IgRg+56
3Nqsaon1odJM0Bt7j7BKBJlKq7v9uOUyplTnwUGMTzZnRWLAzkPAeM+ay2LPyP6z
JkLUNmK4MFDvN3Trw/nZePXy37Wf6iYYrxgakA+qJaRs9oDQfgntb2H0UXTajiHx
dWjUWCXUdSibEygU7CKGfTQhyEX2mcAHeyWH2bli3JijRESGbzTL3TdN0XhKqswH
TcIqe8CTd5T76lJowL0Dnz/KogSta2EJB2YjgGMFZehRPn4kul5zPiuEVkN+qP/l
AcAN3/S6PH525oQKWh9EXNJBIX/gnKGKLhxZ1rRJ/vIwPsdqBBQmEt1RZ5BDwRIt
6Jfzb1qJjGzcMn4CbE4L6pdjOtWF/WJWAWQBsQLcAgpI7X5TNX+ZW9ASFm40iBl9
QF8PQKfvppHSseuUCEzJ/W3ejotthScHm7x78b8oTTr1LEoFR0rGTs3BNHzuCWMu
YZyc7WrrFWWYzPQn3l7LiCH7VV5fBYUr10gBfm2STbYOhZXToE/2VU3uGUd05MrG
bMlJVNGMC0dAlHWpY/9bGUm9dO8Qa5JWK28mjDzDkiRptXW8mCW3U20s0zM7k8wZ
LCXpQrfhkG5e92f5qpAO3/P8efKDNonSaJ2a9Hs0rpwYdIncyNjpXINaj5+BjJ2M
f+jJTOlgoI+1q42R1BC657hImg/4K+iHBSPSgeWpszPDCrnCUN+5FO+Re27Sj1H+
sOpGHpYJG8rEcjeFld+fvK12wJ4FVWRhm4Y3f+1DjvJIN7bpJXzo2aECBgHPfsji
TcuD0DKwVEPxoOe8g7G3S0jHAXUq9SGOaNSTILvOHdJ0hd0AqNemRUhPYE761rpP
YRnrDJZtgeA0/K8PKZlGvlIpl1E9jt7Wqr3B/E4WEv+elGOT4lFbyYFogimWqI/j
oBcHjM8qtu8Ai8iW/EXQeAfuTCNgrLgcjpCpvdaWGsoe9swgDTSh/9YK086/o7Jn
TYd4B7Qe29J3oZ6ljuWnAHnGvlH4u5t/SnXfSAONS2Km+XkPDkR1Ge7usOL2j6mq
f3lHckW4EnNgC+MZ3V2VtaGHvlbvfpozhOPZI5Bwv8FTUuS7SCPojnd9hLJEBGoa
PSOmhw8DSwM2tC1QjlmRFgR/AqhRWGx5EByKacsZr8JBMvwMUlFUItiwJN37UHn6
8GGVc49zSEsFEpFaBky0EcVCCkVB44PD8C3/7RN3W1XyUf4MpbesVvbKYqLtiTAk
VX+NgUo9G/PGErnsTDNEQIqGWxDFqW/tuEULwWiJZb62Glr78K8Tv34M0Q6dFlAI
WYnz2vgIwPwoUcbO3QIN2R1nnvoqYB7oTo+7ZUxIZyvEZGFSX0wOfhWBztKB8Eot
1h0Nzyiqdh49phVBxxysUhY50M8PTG4Wjr7LElvdL7ltWMZOjDXPNXoir2/ptj71
QuL+SErGVi9l5pOT+E4DYonuEDgReQOkc5kSdc4mLYoJcUM1JGbs5FxSPo6klExi
C8nT4z7kwBBZBDMBaXaoVN8+3oIQKiuYYViP9/8etNi/uLNEm5L6lHRBy4FIER89
D9eAbA8Dnqvel/oFt6oln+2t8NBMb0jzWeYz7fYIFBgnjVzEOJBQepCcj7CCyVeg
QL5NBODoTwizxw9+pOYl6m1il3OHRNQKrEOVz0f3aH9QFB0YxAXDjAKcGiRWI1rD
D2mi4j4TAiMc4catA5L5gGvOfdimdnAot1XWoR2YqROeEdyyYVHm4ZnMoNazEl+1
cGew40QuAymxYly2HJyaa3qbssS63gyNULdbE6pFQTSScWbq/SixJIxbL1AxefPH
bRO+zJOw/Z/CGnJKcJxjMCcVculMI5xlAD113ZbGyzTeGeZOAOQb40WvZ5ROhpQq
TgKGhJr8mixeznBdOjIObOFjrlC7/HSJ6Qfb9YlU5PVUNWZkRkSnwDXK7/wZAfv7
UDiMrdR0z6K9NMZog0ySuRrmJuXtflYgJ6ua1r/9z11iHkQ1ClDMdJjZ3WwYdhJ4
sT5Uno3JJDajjLjpALo6W0HWZceRMpGgvmdLmq3FLhTeKsMO+3Whl5NmicEyKtcc
th8+2dozlUO/S9kPbzX8A8p6fS/uC6iMqSnJHTa9YelWyWN50/7DYNJ2n3BkS/eu
yK8RdRgsqMnlvdfsh3fnGz+Bod2M87zsB3akSypNL5nG9ONK4DAu+YA+8aUPVuat
tzmWJR3fc8Q87Pm3Z9ZPb1WbvkVPS6DMfNUO5EOqG0CTbIFWhmZlF0CAll4CHcKF
q6qfjnBbFQGo3EKyIGdEvlnRBaem72N3JPM08vy4nGNZU4ntjxltaetAZYgNbcWi
AMF5uTYqRnB5hELKWPdE6dE5qjF55qydbQxTZTm+9P0x9GQ1x4r4HCrLXyq7Lxcv
ihPsHTC02RJidC9Pwju5+ROaaOnUG0wI9qwrGiwpVAxZHmXEWUr/pbOqygj+KD1X
KD7KWj4N1qPFSvmDickw1/YXSmrvjEfZG5adHbILtuU5Rd8Ji7aZNIKt8IsZDRR3
g0ojdPNZOw/k9gznTEQofCUYr8WJvxIORD0ou6+kNvnB8NfzQhZeAr51k4ZZbuLs
LRQkBojJplvD3HyVYuIbzTwcDQuN5F1F9eCIbhjlft0k3z0IqmX43pikT4GDhd+x
D73Nmvj5lzwbsvfy3X5ZYK7F1b5pL4lXACJSlxGkEQEDaDwwuIpvb+LYj/diqjuJ
qSuKdZTwBEfIDF0pk78AtCzEN1ykkE/4pSdLypVE6OdhIWAGLBCuehJx79oP2s8G
LdJ6kuKvCHFeF3SjoaZwTL3fkh6ff2q1q2D05jbVI7Z6LBAYxLhUih3sMlvLOB/Z
nXCDsji7uYzEcibqQp4qBVfFS2yclwocYMYYmFDnsFYUPAXwVyXMH8ZLtMcFn15t
DfqhQ9NagCDgDfDDJIG4NSIn8tASCJGo7356taXmtl1WpoGH+gdneZv9oJ8OMlhZ
sRwBW9dRC+o+079SImubgdyZArIYJxFRz2o+2Vpm4X1sF8RAXkegwPP56AsaQ48Q
DuXO0BBOEcpn9th6PTcK1CXAQgMgHXUDouIIlANDXG9AlAjG3fv4YfUCoLqjHNVZ
3b4/Aay91woB4d5dR88qKh6VJb1PKvGWs+evyP8C10Lm9FMMdEpqrS8CiwLp+kYA
JqqwZdlNslUQn5JmPv3wlcZuS0bXiP+1sqvDCdaRhhpm3PHQI2Jpu87bviJzOJkv
7WeN/yqJbHz+htK7+O/Qc98SwSfChudkemWXlEwbOYiWRm3qRwGNj7YnT/V9F9VT
zAiZVWd6DDYJ9/y0oLrwJFfUICmmGQGRithpaazuxe2HFXw45Hq8uD1OSZymrhD+
nGjmDH6X03Ms2Fg1nNz21YK2gxu5yY3ntxpNcKCvc22y2kzdlNM4Fnyf4JkWxC1w
K6r0bmTPv83y5U0aQB/Z+n50/ucYzRyz5ftw8Nxm5oUfCoId+Z+owPTahheIEWfj
zotEk+XkgLkJOjfS1szXqb5E40cI63farz4cHGeGqPpXRN9CY5hXtItcx0riJiTu
6dM10E7J/ScuhrbNSPCqqG2Q9G6uRLLPBzrnKZMlTTEVK6y59aU6p5FarzARe6/7
sI4AXYqx7rLO/Pg8t2cv2YPwVFPj+fk2eYm/6raH9GnrPRY48+rkV7mZncGW0ZXR
mN3l5mOzDGRHGsebAX6gWspobysAou9jClTJWDkdxRLoLi3NdT57/L26BV4iEXcY
+0MM3FUU8YSUFjoHa23igNOj7utG/FZ6x3BHcpSK0qK7MASsu12DsMtC4Z+XAQQG
4uud4s169bo8IWPJIYv/wJ17+tOZJtISRTqmrCaGCX5zWjjB/JuZMOpp8xT78Ayh
If/G+ETjdmxQL2jyIZG7nXZ9KPxmXZocVbD1cwZHH2h6NhtGVH0BGnWmkaRqfkOy
naUzm1eadVfOhHDmJL1m8Xx5PjVtYbtjwRucmNsl5UFDDXCXQWhR5xux0m144Ey1
STJqtsYEti6gs2L9Ij04sQVi/HIBGob/FPO3H6s5tf47MXT9yw+jzFkaQS+5Dvp1
AaKbsL9+9kZXovbXLDI4FM75c+u0h18gNJ8v6ZoanJDjCt+giza5r9/OKXCunRfg
jhzYaLYxK8sHzb+xtHaZycMjcsU8nI4BXp5SutrNuKzoNI323RNmcufWg+syeDu+
6+gw7Xa4Sbn80tQpfIz6qVTnb8uFEuLnn44ncY8mo6Y3pP9G+GbfzWHtD2P5ugOe
VhsYo18ZUZgnEBC1ajSN4RF/Gbn22rfFzLnllbUE7OmA93allfFYk/4Yl8N2Wre1
bhrH28TltBIEY5MD5HYkKiUcImoHkZ++I7DU5PyqXPl0/dF7zVPn50Q/H33CZ8ZZ
OF1EoHe4rFV/TQ4xnmtmmJQ1ZsOAsf43ejAsVw2+QmDgB3gBylftAOc67fSW8yA1
UqbesqKYYfzPNCZYqkd4s4+IWsQzITn9yhD+g/fwflui+SFUJRaJR5F+eR0KIb9u
fo6zaxDlo6UgTujxGTkr8PLfRJqHZcLzPCCkL9klj6PSmc2qsltW74uSkUu2dQia
cQGSLbXBVrCZzsAZiyL+CJtH3M2j5MgtHAvu7dyt/G7eX6Dl53gjfva4U/xGnTxD
vnq7AQON99nBBssEd3XiJl4KRf6b0K+zgOfH+f8Oi58TjlGALnBbLAq6If+9H8B0
pkpkemqJLz6W54egyovvACn1khs3p9TvGpy/2Gph42DGxlOS+CaFsVxWkErTbLHu
Wuou9Z0lMXsewR19OrSbitwzd0t2ulsEuqzu33+NgskES41jqvLIvszhYls9z8BJ
7qcyohtliShEC+rBUzDCgz8/Y0p78j6DGp1hhQpmWFlT8he+RracfEy+w12GXFf4
7J+Z8PBlLten7De/MNbV40gkKQ8XGbEcWRN48gq8Vc4rERFUrAe4GDFxx0wt9JqQ
JE0vRin5+2tPrO27SSzxnIBHK/S758l0CWJ8q20Uqk5NKMlyqP5TqdXRCFhEKjdz
PJTyeFA1IUhTfLaGD43M5r7fB5WFKW3X7trijf494RiaQ+qPvLMjJw+zOzbxH8xU
hi6bGVQnlPfq2n6+FbgKxZMiHAqdnUABysutdCSal/NbvIvXI8+xmaqnqlvv/mXI
BRdZC2d37+5LhRacSY2gdqSEbFvSrLIixMN1td/4sbtIoTbiGi5ckd8wRsBpr0FJ
f41VpKHryUOlOJR0DCYwNhUsglzsE2iW4lAPJ6q1guSML8KGTZreuBsm0XseZl70
aDQMNymeyrfbRwaHS9gE0mE0YfhqISMZSIp1I40dvR9ZscWK2cZswlbeu2UhJZsm
CcmdVvIqPBy3Pn3cdUHJGEZjdNISmBcUsnTg8xhE4E3/6Rl2Er5qPFp2RueN6h1g
sWc9aCwyQdwuqS5puLJ55spF/jyBXUJtSKXu8ZWSK6MmlJ7wNYF5PzqKX9GEvFF/
bLlRnXvkqg+ycbWjHiZU9jI5mhdH/j6Za4PY2/8SPE6fQsJru66FpkGTSZ9Hl+NR
Xyn7Djuq2d72LZbRaUq8xSMt6WwAOw1cEZiO2DNz8Yih7yWRjUfNpurQv1BJgB+C
lgZQuZyTbWlvyPCZIyifNLgTbc1c+KlkyKjI3nSAA1xBinfe9HBSe0UIaZ7YKLU7
Br2MpTFxq76nQCQBcmwG9/2z7NMKy818OOPYMxrSI4MeXEdWf0xbBBJddit/RrZ8
xcaXzNKJrS80J5pSiMChYiEm6mte9hm+SnG69I40WWJALXivtULdtsl2eyOwWbxS
o1dvxV6gn1TfK1IKJhShN0eqN0Dtox5Ey4y8+masoYi95tHNxt6SZ13GUuNtXP8C
3xMejBz78PYju4D4/honAzy09Lg0sWqMbFeB2dGVdQW6cHCpHWE7SQC+o7Tpy5/7
uUbrpvG6r2iiKsMy3pskZKlW+2yeHlre/+qlvMkh8Q8M4jHLlooffDt9lFCK01CK
VLRCw5c/2npOL/TIWisgWzow6ezmBncyyXF8YE2GdyA+amLJKvBmJ+v3k7s9nIWG
+NvlgCDA/kyAIAvd7Qi5N46kd4rLxlRJg2AvKSrxp5RK0Nue/Rm5GJzElQmPfG9O
bCl6jdR3L7hhq3G7BtyQO/foqC5q8JERP7IOhwa3ZIsgBpvHolVDcDnli1RbqlxK
zqIRtblSgxyNdD9fy+1QU1gIUbRYDQRIpSMLlwQcpmNr8EpK6akZ5BXDC6wlPNcp
UPbfR4aagwea4M2liCEXHJ8Jix33QQpFQKRhmJb/zdWe+tioWK+4Mf/QQONviXcH
jvU9HeiLCtpdRWI//2QmgewG8rP4g2vWBSWyRVVKSdztc6JMI4TCgZd0WNhMp6Je
DVcYPn7A9Vm7Aydpn6TWUZcrd7LVw2RnzDr/osybaThN7Xnd55cZGwzDSw5GExux
C5ZrcY8Pr0oNJl3i7evM+XSrnBVHMzg/YERPHag9M61Ud+XsCBI5F7QDQeOdowXF
phKXLQDTJYb1vHb+uwgES192J4BDWBkufbYJL4qhvXKJG56aszXvfIM3rbZMpY+5
l2qfBMo1v8EnnQusWUJA5xSRc0jeSxvBd7thJ9bdjNrGE4U57nI9F2uLeGin+5HY
U6Rr2kh8LLkFjgqgUsarCWVk+p718Wsjr+Ew+u4tGdIpkM9ybxo6YtAdMaDCwix0
b82yQ4MTCdnLZ6e8m1NlHPFKoU/bU3VPoASrP8mGRvEQW2YfpCbb7kaw4cIMWa6T
vYNjtU7Znf0O//6r1dbmIGasa+SmldYLKNTedlHyCTl31NJQNAbmxtPcD3UHAXgb
jZApVjNfvKOz2a05CHXwc6jrf8FZmu5zVBH79d+xjTClQSclvwtHD5yBZe8uzDjZ
+5zALC8Zu9eIEi2zLOQzISuvRYWtB1aUfO5mlfBks1SoEhrgupZAtQ8PzXgxPuYu
CCL2MBtk80giFBKjS3a/Ff4V9dUOwHEaA1TrL9YPUW0OPYdc13RmUE+t/Ny9H4PX
BhYzs98or4XVYugp+W6uNhsuUIYSj6Na27MTujb3cpc/sgU1KO4YLo5NKZsSXXmL
M6RFIEEc/q+Lc4ro9ia02VQjnE8KV9qYxy5SrHvDAQK8PGiyFs3UMCH4M94xVT80
MzHngUCY3me9rKAUayhucY9nzAyUW6fVFCCSbGa/dKhaa5QFqWArRToiZS+/a5/0
9jBSdSnAJLacEXam6tHmNE1wf2qm4lx7FSaTxnZ+fpTraHKGbW8rxzK6beYdv0SM
2T/fvWIpjzSls21zjcHIc/nFsU8lf/tMhGVjwdhenC6JIIoTxRkt+2Is5gkghA+F
qeoH9wmrq3yyETyHhFQ23lN0GPCTaOnNT9bLIzfalSyQjFBPMtkZtFEYRe/M2s9u
OrEL4Ph7ECwJ/Qa2+bo8DZzDxO13VXPFtfUeHuhGr+aOYd768BOfo1VlYW7VlklZ
0dkS1qJxW2zIJIgbCiC/7/hk0kXXlGvFLLGNJibNeN6JLWshrerKnXmG7lHvmTbu
He/DnrlYZe86MHLScQOuJX3z0YEPusWBmn0vdAYbodlGrqbh/lXm/PCixtT/Yg/5
cpZfLSelwjLJXqIDy31Zk13FOnIss1kSavu6lDI49tKEr8llKwmGW6s62nA9pD8V
+xahxz80jRWzoDHhzApBigWY4qFFujdZYt5dCAQzpUZ0aT3m0D3nXf1Dak9qa0wx
sTDyDCPL4ollIoAxqfYFCeAm2W38Pmq0plszM4dxkt7gFMJE2jsaCgnSm0sikaU0
U18mLj60d5mbgPWCwJctXO1tjg6FmZ0prcZosjfQoa6EF11lNCh4pqglUjEkQV/y
xGcNEmKW74yzuWqUfHSRwvAVmFpUI8HCAOmd5Qds/QGYzYXRO99QcKBoeZUVR3wL
3cQV7u311y9lvPGNBnLKC+6hg4FM6Zn6JSNNT8eH2Kdo33yPdDNAJAyF2Ieh2hv/
56FW2hcyZ5kJwIVMapzDndazLfnZsoxmw15CStMobUsE31vYXAi4UQdEmCglc6+c
EsMVUIGszDXuwRBFSbTx8pXfrN4NzAVbDk5hnUtQhRHJNVzBrD1s9xdyvR0ojSGh
nbzhHR5acLUfoauIi6fx/iHJ3gCstY9ooL4N/ihl4uMKZOpTrjJOiAn7cC1Ygoq8
2mRJC5RTZaHAAnnjMbojlTo4zYia0i2NFOQ7653ENJwNY/RG0jXMC9IJO4UxooBB
YLbJ6CLrPK83uEZLefhIrs9/V5bs6LztWOrQdnR/bxOouaxL9V2n2DfRTWd9ePYQ
S9V0DdkAckFZhK6AXZxc4tMXyqd348ouiTo89E98rkAgJK6j3qaVOl5jSIv96wnu
sGWxAfbVTLoWHBGbo5xU4WoPP5CW0wTgh/xB5Kim3IIm0eaolIfwZMuRqHaXrdYl
zVrWArKgkFqoeVl0FmYpOF5T8mA9nAOpNzcNqY/bV0vSPdGrTm3gQzijlPaHXXRU
f1G3k+HiNwiR7+G//Z2oTMEQ0K5sujtfkkW9OFZ82Wb6IAmKpSYdYXDMR00CZXlZ
HH4HoKSkCk2B0BNhqgSPxTdG2ge3HiN27fX9xHOfY1OMJ0m2SsK5Od4+IE04JwNu
GNODBAveI5X+3xNJFM58teECzFVXzzPqx8PIW/4yJsmBfpHY0PuVGG8pSQUfeT9D
03dSab0kWFjyixVDydcpLH7J7ogtVVOzMHiAEGObD+8x+1AWr9Rk/8q5GT0BFaG2
AhNCDhpWaLqGbjhEzwIhQNU6SP5FSxw9o/xf9kjpL71RzIN/xStgtu8x7ZJSS4Wg
tSwkXzpubYA02My2bnsi4tuYZI6NvSDycmFGKUCWbGAt18mTQnDw0Lmg7x2NomwN
jb43+j4ybAQLQC68QJPw5UOSywe19B52JDgrI4N1m9105+yi0jWdCAHitENivWGd
DebH7oZqXjk1pbSb8R+Pf96OjEAnB16SWj5IP37z9QUP4mH3YEUN4i++Or1ylcU6
5xZip2FpK60CRYRGD7oC1qpOL0Zzg6RQEYuGrrsmiLXN9NxAjU/lHpk8FFXYinK2
vej4twLlFCCzlgWYyGBSyF9Oaet82AsG2TQxvDk+O0yhlz6GvYniQggmqprL+Ilu
iX/hB5vDnxdW1zlDGD2clpR4NYOohdabQIUQVTELMQST7xBNnRHEQVpFTjJLtUIQ
bhw1MbD/X3hTOPHweUDRegZZDLF9a+bjL3CIbwbEW6HiUmxtTiVEe405Lhz1He9/
l7q+/XG5jsvt09cUixTQZfcNFhQuMKJ458S+6u/QEERqX/5ZOMbnF1y79OfSId7u
4d5a2pW+klKXy4kNJzFtkRgM1nJKR1IZBCW0jPneNn3U25TdPX3DHdmJDF0aEXTi
UYpsm5OZCNW1StZ9BouWZ5FFcoN+EbiNJaCcQdO1/KN4ZpX4M+SVbr1A7DfeJuz1
dytIttMgORJBLsVRrcSqNxhuDI/N8/lytxdqFfABU8VS2x8iOtT6yfz5xJ2yy1I+
Q8TaeTyBQM58QKML4pYeq4NK608VOY5hAzFdkwRrkTgkuyjfb7Z8i4OISRdJPT4L
cWwVF3FoPXTVLJndZ7B7MZJQu1GRyp3gqzp1vWnjfwW58ueZDEbwdScN3+HKdoaS
skpJFGPf277nhgGVh+aCaJjrJFwRZH3gDL0aBSxMPqFYNCZvb99Td7qISF8kY61G
Q0NirJqTojJE0Xtg1VRobhTI1zZ6tjFGFqsSBtuC8UhLehFo4RPjkSVbAU3WMZCN
0zRy2DLKBSe6jVx9tKlZOgoVdoEl/Lwk/lB44Cu8PtrYmMohZBvgbF/l03KW3UqN
Fpou7NaTKnspUC8wOhstjs1scfrdvVhBcCfXp3M0Zhavn3+uwuL445QX24YK663L
gjBf3HkveY2nueck+8UKIRhwiHnZOUR99xud8v82z1phWkeM3Gxcoezj8ESoM4ex
vhLCh99I1Tbwzif26NFhx7Vk3jA7Kve+howChe3LGRG0vCkm/F6IkVzaeQy2uuqA
iyz9lIFl5yv4nqLrlkDHTels/I+bPGLdEqslyGUGZvf7iwxdodYynmGYP3tCN7SE
iqV+Y+V6ifrOKCv6XiH8SO/wdvkxDqJn0kddqHuwIqocr3WvxsyuPl0gH36SBeNt
PxPQziE5m61jZF1qQQoWaCl2hnsI5EE4Tllrks2KCeViW1PUo5ib2r4xX7zfGmEc
2fVzZxOSB2MJ6Y6X+zPKC4/Dc/Apu0h0MMStIZZ+fHSMPvNi/2asKzuscM9mPJ8T
dmdOCFkFbRM4HQYEMrepkniXRM6ncRy7ujVU4XI1AdBxuyMeUcrMO/twQh2wHQ6u
uTdu7LlhOT8XrSpmDs4CtFW+xd63t+1aClM6KR7vnsOXwoRcCXoPfS/sjd0u7dPa
u5iVLgKn6RtLsvL4BSmIqC+5TPGdf2/QiV8dY+kw1/+3dxdtNzg1umiFuki8kjvh
XF2jOe29E8Pz2ZNnNQ7Xna4hiuXyso85nC3OGdI5V9OaecS5ZkfdIlQZ9asMlVHy
XXnLA/h0mMRodHzgofjBR1TYTPhix6N5iEWjJ4jI3fW8SvtGHJ/Tww45sHaa2DlE
m3N2UdgjbM/8QJhI55z+/Jd9izcJ7OqVL0QfC/J6oAnabiKFa2ox6MMXwVqGFk9A
oOYY8Savwz3iJebb859BaaCvtzJBpF1asytajRR7OAH3MU8JOcssdHC722fEW1DZ
vmDkQB2TFGLTNjNkxPEs0l3pnAi346qOEgLsel8071bMDYU9J/1yvpIq+HF5PZR1
16KkppRa09hNFRZhuqmOQnk8FHTuXuYWd1oHBwrHetqCBqdvjbJqcD2ATZJFJWz2
dDviqxI/MONigyF7kzJYlfkBQQ4vnoSZHQ1878jYTk95KGPG9WsvxxI1cOY/uOSw
MtaHJbL4uK0ObjvZKqFp/7/fY3cvsLijUXBMaxe+DNIZSUgjvV2Y2npdRCI1n49l
p1UDuvBPsfGAXcoyKzgKy8Y34maSBCywANc/Z0tYM8m+TwH+Ze5yx6gDZpNghujF
z+gmWLodcewf4hnXwPGpfp75LNpEfZP/jtGOy5oUMtcsP4EA9dNq8P/Ei10q7D2T
0VfHlKEqnhNCYnpZ1Qchgstx0dmf2Oz1/b9ZgX2OfTmPEiJRzi4e1ABsD89OnOmC
Wwgt+Frt48bkpylrFOlO1gUnBg2TNOuWEQZTHsBRdqq0pxYnfmW4wEeE74wpLZue
qDGskwJeOe1a1mlJD64FbAodHZGT0qBoxATgo+N9xm3MEcNEdgDJ8V4LHWHLqHIm
l9PKT67HuTuQkiOaSTMvjf1IQyGugjFhCqdlGqQ4zqzVLCy6XBzVz78MHRvCAsWo
Bh4wqu5bBP8wD2/22/BGhXhCceo8Q9bCh5dC+jAqhiMGPuzlm7EP/f6yKy17LfBX
VK1puKVS352V9yDHu/03RnZMHVbZmRLVWDiRPInWVrf4k+EUbE8esMzFj4EQyNd4
rplSRrj9NYOwO0h14es9Qon0BPWW3jtfpEroWJUJ6wE4kyTk82Rv1pV/3N+76ddV
wqV7zjGajK7AasecmRBiP0dpeNPTLOstGDjuEPlyHxGpOZN2qjdXs7w5MmwGskk8
bcyi3XwHVZtWhvsOP0F70aJx81VDFzSTyP16U/xe1Cn3MmJppjzxOi9GtaCxk7vJ
saf++UmYSEjip7tJZ6ED5sX+pUUa/yvFW1qMPqqHyeEodlv7tjLPbN3LlxBOvMni
S5voy8M5sViOdGdBQFoJuFlmtfk7ELVMvXKokfilS0vsdGCiiEITiVa8pty2isAP
QyiDHRQ9Rb0DJ1Bto4fXEJXC74e3eJgCHWbaFLXD/SJ+SDbt8lEjPntE9Ud3qQP8
kMMA36mCtUUWUrCPw71UXYI36F4ovZzl935TzWtws+RbqO5IJrJZopQ1Zwt68ZWR
no2YnWnE6UN8yMJsDgLu6LiSlBeY+xXqxN6eV8M6/MyF2Jco/mZchO6SwE7B938k
eO6aO6pNwIlydyh54l33GdaIvmZiF8MdaAGIUrg7lEUD51S7C4dny/LEo6UvGKIv
50gUW8eSGH2MOC3w0Jn9YqconN1kaF4UhkNiDMsuk59aVHJFhjSz1zlOL4HDmehw
15m9oTKKnbiB7vtRrDWYuW2lXT+xsza8s6l/VPosoDbX/y0dYeZ9nbIzeV7VIYfM
ySrToY8kvrR3AA/llLfPwrhu6DOfffSj6psRsWKzaAiysaOkV8MK2Xn9CSwoVFNj
ceq1/J6eph680rfrRAuX7D7iDdge6oEpBmMnIofAA8MByGmhXuexFDbfcVGnlEnM
Sqiyr8L7CB8zf+iG/JxFB72JkB8g4aTL8lP3kqiMBK1UmZX7rPJ/D7bYDVlAtrTF
1cld4kSFzNvvay+bDUMoviy1mlyJ3Qsq0/DB31/rPokRCN0cn8YABLRbqmYRBbhu
Lc7ZRYxAsbuaIc5F4h6NwT+hGgkeh8FaB+ZQuXQjbl2E7vGGJykWARU0uRBEudY8
tO/Rw5GZz5tbiU+CGnuKUOUbcrRuhaZ5ibNRoctKyg8BXWbbLWYEquJr7tKJtBA6
ILIVyKhJHqUWmwDO1P5ToNCJiPEOK5017sOfb64DkZMnFf8azOgLzoNgJlGNhf7W
tyD1UnZ9fHwjvcKcKP3aG2MmJySxoWyd/tF2jlKagaspq24nVEOky0mcEHOOQHBy
rt5VTL8Q0mxFFGh+dV7d2+QgJy6TCAAYEVO9pC9x9h/4qvqsqjJNj9409Qo2nbRq
hZWnTvPa5t7+JVLIYDMknkfSPoOZ9wTlgZJTmpWQDQVwoXPS975O6Nm5LMuKFRpE
SqSub9b3BnzdcUa/vVOm1MicPczZUWmfW8TlUsrzmQo0ua0VcQFO7clej0JnsHAh
zCowALTr/K8CoGIB9IykIOhJMWm8AlrGvhp+UL7gzDd2SZugQrj4IdL1E9EAf2uR
VWn9ig/kzmd3V1dj3By0bgCfXz2OAjDT97J1ZUqA2vb0E8lthmJ0vxb3JSiIhIWh
3VIhU6ezbozdbHZyJuUAwgmXsqZCWKoRLWSwHsyOMGI18xbU1wombQ9Q/3+2fvrx
PpAoqb9l+TrO2h0C/unCEDFR5x1nWORsFS+xtCO/chpXmEUWar8LztiFp5qd9nhW
Igut5EuxmvkwEmST2qUIK+mVWHNfgsxNf277INCFHavbrdKIUE8OFtG+PGqSm8eT
KQaMfuUrDvzkmoedk29n+qWgEDwy9y4t6/qvv3kY8JIZAghsX5uVIFnR3eCNfQsL
roXt2lGpOYIy5kFwdBYDBgWO/zrgFzsbVQCe1ER0p9WHPmVzN7G7wXHRlp1201wS
q3zWXYLJrxuRcxPucJcD/8DO096XsSN31IWpDzaiMvEYHn+NMQNZB6hhyUHo8Tlc
s6olpRWTT9ODh5lbxZoPGQ/xgzvHi6OTWXW3rtZEvkspJs6JCp/904TEe++QFvqY
AifEYOjgatRczuRZzDbwp02qEw2+ZwhMJrTzg2TOFiP/bBLntrYgxw7XS3pwgiY8
Ue8FSSURz97dIMzYQFMou23/tG602LGEbeyTsZUONb628BFWCAkHrW86p2xFMK01
2lwMBtpLwC/1fbmp7ARGDekOu+otG+HSpZwT5Fi1fBKCfbwHm4x3p1AYYkAGcKDW
lL9Uk5IdDXBOe3igHw8ocCWEHFjn2HDlHAXLgnWYIkob/CHH8Aqbgf7qpzYauE0E
uhRjQQYPE3CDYtM7sB+VYKLru0bcL4yYDtBr8jKptXgE+0ekBHZuQx08o+8yyJ9P
V2yKHNgB7m27BP4Aav12+lpbMKBtgv+5wyAFaqiNH0Xe0bQ8qBMPs344uDuWU86w
Kf+QUceAmLi1v3unxTdROZNWsDKrwdCNJYS8Ty1y4R3UeqsR1S0ecWluv5Zomtoc
dsd2MeevlWxOy51Dm4+VfYeWt+TQ36IZKbOU9bKCooTMdgCtxeP0oLjNueG7bo81
MKFX9gd1hmIeIeNV6d8HwgqYy/PJWgr/QGFxlXCGJ3j302lSIROKtKVjgj0QTBNt
gPrVN8jJtk6bV7L/uvmr5h4RCI4r5Bu4nhMWSQmfXz28ou+9+DMOZL0PYA/mUx3P
8EC9c9zx9D6E0CjxLmDFFM0V7hS/5cAlOGPqwxN28ayJR6oWEdKaes0BmAQWzb5G
5DW631suTMcKu9QI17xV+nzxBK/+eWHetUbxInxTtWzzFfQocQf8gdzXA5stbNDJ
+e7DmvP+yfkirYUc1qe6A8BDDsWL9IeMvCHvOrSkU/nOc317rHp0AEloxTSLq7bZ
4IdDdXCLLjFgi8PdNJ77tNTzqz9tzTW4AsXHVmZlbpcswoH8rsNw5c1tK6UUp4ht
2O3pKECATG0BC93DupF8tz7Rq7ufApYkMjkA3BgVoRHhZmgcAoTY+mcrrXDxcDZX
9tHA2tEY2AEo6hs9fu4vYkpL8jmLW5wScjAHVtGzypoCBj1F99TtqZHm+NBFvE3V
1o1928SvrVzq0bP52+ZKTdVkWQGtr5hHR5nBQGu3kzLN7K1WethxAjJAb6Zx1+uo
Evysyg33gSoHkYFjvXC7MKf0dDs/lKfFrHcDRhrLLBYh875WERYkvnvYO6OX+yXj
mLWsIP8Hqr1uA3fC+QNvrcQxjOW6yOEDlKzTCvne6fM6WLGxY/dQBhbVf2c4MBQX
IoDY8ZZhTrDAodaNZOEyVQAGs5mDBC73XX6d12qhmjeCdvw+YwDgPZ8/6Vqqv4fO
WWpYQQKlzK0gX6qZb/O0wvt3s9byP/GSA9Nhzr9fEIB7LSbLAcf87jjWAvJ743Df
vz71CuGo+OA10Y45XLT6kJkgYB+eRC9OHRK9ylJHEvh8Digmt+1SCZfTG3jnW6zD
rKJAWRPpfNkyDXMzZAtIOXE6gJ7AKRhKjEbaz2XxgVVrO6MImRzo/U6Dn+feSFpb
jgTF/LeWd1TnnTejqQTiOatuhOyLlvs5xqY94EO0cLjGDpSvsHtCsB/O+/ZZ4t6n
z6xlLubk4idttQz0upH5QhsfVPwDT0cco3KW1522kEe2X3J3wwZWnDODYgvEHaKB
yU6t76ddewCq7u2yNAFk0kImTyeESgZ4P/CcYATvWkkLQyVjueGJdVPzAjagZYir
ihGZn111a3XJQrY2zEcPzAikjuTUrAdkaXRAgPNnUyWideF5NyOgv1QG0lwdvKsk
LlX3FLZKBt6V5o83hhofYbgun9MSz7anR7e1qU+OlBpy1LZExmEiETGRJf6wYpTS
dzpBAQ/tNME8ACXO0nG82NL+g3LJqdgUFsOBSZc5mBUG4hQwaee2hJOhe3nNF9IM
r/IdTSLbuyznxxYvXCasYr7CDzcqRNbmEeEKnlPqyAG439ZWuXY7fWg/wloHtqt+
p/pC4Sj9bPBD8B5In0t+IXb/KdBTsvujtFErTBuLOEI4Gy+eBLg5gCifTNMP36UT
BfntXJ5F1dh2OlHjSBNh08v0PED7qXNf80KihvGVVfXtTk6MjDU3HIk+EFN815V7
AmfOKOwlfJ6KpOWxtbX6/h/HhHnuDKDaAufsvLCrczTEwpGR3AczJq0fO8y5DR4U
pvtj0c3fQFq2ltJU8ubKCFBnSxBZXwIjXukuAvXx8+aMlks+hwk0n5ZiB0P0uhMH
IU022lDucER2n8WOzatBLCHyllUKCwxqEH3Hfa7CYMTr3PIc2lG5t4FPxQrkBuNS
mpgBqhiB/W7QE2Amko8DqYYdBJOrYnM+bLCyNFxbSRVBBdK1h9AmOoafqxAc/UaB
Ko4Pe85jPv7OSk7Ze9pxpFS4MY80+fwYVf/tz2CQnzfKv23jMy9GK+hZPVjQWosN
tw66m+n85NZ5xhzWirjzISJOlSJBDnqq8Ukc+FSFtSqsB+un5dCs9yAHpwZlv74X
YSo2lT49vbg+BuHAtILKXInnE5nfBDkSU8J+iIR+6e5Icfa6iQw9jSj55w658P7e
UwhMBASSk3rGoxY7PkQDVgZCwHoyUGw/FSE+oBeqWEPrR+7rjvu7/lIo5Uqw8Zub
qSM7xUVdsZFrVi6TxydT/HX2gJmP6qzW+jQB/vOl4KcA+lffq3rWKmXIlp8G8OAB
YGehn+CRxyJCD2OxO8Qk97/SqzlwXdXyqkN9wdB1yERwf0EyuVXwAygyIkgw50qx
sabnluxLsu2N8U3MFrwOeCLztiipEPgAXxKfVEyH8isGUn7CEtEQt1wTQjO6figp
xqIIEcWDqI2A9HRE93UeW9YjTm8bByxOP6a9jMNLXxgVMyLo9jbV/KeugsupTFoQ
BXLPFrRglqnRqNSYna9Oa5hsqyZpZ90lGgRbIw5mSYCKDvTD/gIPWeppFfWlVw1M
kxZNbg3FH8acN6NFplSf5RCOc2h57szDBj4TZD2lUtTzFqwZeFETIQOoZUias7e6
Pj8qWRO3bZqMKYC273EOpjvpXZzb6H65MrWjKIS7Py0OFHXyjLPVEBh7EiKWVqWj
SB+4N1wJ5LXcl3jGBHeIF0TcUMr9p2CTdpuuD5APjZsbyJPcFSu4H+7r8nyOFWLI
FpX5/IvnLixS33lGAPCc7BKPCJo1itFWz6TlxNT3KDflUnXFmhrgrXlwdsaN3V4k
OiFp+HvQ41shQ0lNKessvR16qGTr/m6GTszzFlC4A2Y7VVc17CqZy6lrBs3FXaYD
yjU5Ti+LJ8vTtpM/uzyXhNoeVqWCLWrzo7N2UKqQalMMcfBg8NtLAUpNCbdzqh3s
En1iiDyTad579Tn0VMd2fFFkECGWZankDFOCHn2EwP1JxsLPVZN9l6D6/gshF6F/
n0Zv5FgBcwqxb569qide7loloH9s4ge3x1n2gTNXoIC6p+VGSXxRJsmjbNDxRBVU
VVuif1H30sSswT7GXI2cx4PG3IJuHJ8pqWIdRi04rbBw3Fgi+USXDQ39azWTNYPl
mC26OHoeCdPDcd+2qumqcTT99HIsQzfRQ8it+tSl5KKx4Yz99Ad4PsWImUOCVXC3
tqKdsam+tGibknVN2GxclY2dBUou/ky+u3393/dWhE0DQUxcUjX7oAhbvs7NMDCJ
Igmr06GvbCsPMRKAWqJr9857pW0kEWu9acbzaOSo4qn/3RoyTuUrN+MYy4OegWYq
QkslcdApfTUJMRCVLPSTRuMhaZ5Zlnkja2L2qvGCdmT3cyMIUJik6seFIXstSN3C
slz4+et2BqtSGNCt1whIYVvSfR/62P8GAXta+1hMyCjKlPFhG7x4qQAqtQw7PEtC
t1M8gdntHSycCp6ukWGpK85NJZ087hS9Rl0abrfbA2W/1+kn4Z9BzCk/GtG0sPdw
aw1qpTs4C3wQVJie7+oYzi+AzogfJxfh95mYVqqGBH1GeD0gbQh6vYXEze+nijby
cfkutH002KlhDrQX2zg6XACTX9nmOr9q5Ct8DkjEUYFv1dXt3XSIN5UZoL7LpYMA
DvolAlTC2WWrta9hK/ujpP87Eo7whXwxTRW6QWniXW2gMa8mYhOJ+l5bA6XlGw+/
MqWRM1IvFcoAMzd+wXyJqqAQF+fow7767bV+ESPS/OatAYTPLiACA0UUxomqOJ4x
A59j02wXTPy23k7qnt/eJKBx18lVnMt0NVuKS17oAQxQpWpQJsdD0fbX+7nQepaS
ZhSs+mttZvZ64TzIz6oXfa7W1bV4virCjo7krOQwQTsEqHuFbgEr32VRU9+nzzjw
G2EboDtioWBGNhjsX6dZuk0N09gQduStX16AZwDg/49fO8gbMpGoByqpI8C7sp8u
1o2jzIirbYTdHpFhg9jRcE8/nNx9lo72V0OuxLdrVY/mQW7FU0FabkDGbXLWX4w+
prvWGvTgmcY6sM/9IO4/qhbHQJDISmbaswWlVFBI/NOSLuwufMX+TzAzXa27i5Ha
hKfMSjNlrIkA9QeRkhhWtDFlE8DGU+jSvV+1Wb3ikiRj6QFCS8zjt6jAcPDsQv0U
4wsPklpBDc6o5YuyjM0lB6TeL0r7zfMicITWWNReFzUtwmdycJdb6B0fiKUA10qh
g4C3OD7fq+3F7pNUawU9rzn3N0dbyfe36ayyP2KFKH0x/D6j4jLgblV4eDpWBIKE
rpGrqoD+6s4dnQ+cSPiQFp5v/21HcJLIdUTuojwcubl3gX1fxSRTHIKSszFneev9
tTKGsGHETaesbXY9WWUye3fpFbhQ6pTmal7gIgJVXNh7ykA/duBp5f7WZWoYDhsB
2q7Wqyaw+uqa1kcq6Mk/0cpPefIc+r9SDb0oE7Bd8tkwD2aBsUbNfjsd2vaMtHrW
OcArSIMr2dxI8XYr78SpI0/8BK6a5Z6SxbQdiG4sSNoKzTlHhjpCxACSIS7r144c
uXwU9PSRtTfiGKBdr2pX6Wt1E9AXXxOqTMrNvdpo4XFaCYizI/ZE6p9N6UOK8J00
vO7ZBujcGqc/Jx2rQNXqSJoQmO4g3UGop4rRRW0e2VttpGtsS5GYqZ9/dMTOsXuU
yHVtMc0qldPkVZIom5dDjIaaQWxaMi70WHPAEcukdRqmHo7JwW/CcF7gh8p76+AK
Rf68TsH8WugyB0dHIGmnaT/m5wr+l2uUYBQpwV9cs5fqGAFNTUYrFSYM81F251NA
hUq4MeDcSBOYN8JQ+fVNrkGTMwJyObI47XhAQlcWHu6myEIKx8Mq5f45KIxmTmYC
lYcO6gTTaKka0vZpxdMsC8iuwG7AlnmLzPOhaiDooPtrsxul0rZRRok08XLEp7UA
TdrPF/Mg8G5XqGNZW6QYFy++Gvsg28uA7Pjm/TIridAk3xSngq67nDgKGMZBA3Dh
8LfutIw3ohdO/Z+3gBrEdUNTdwKU5PIfX7lkibeZsiumsIVpj6jlsq06u+AfIprW
W0VCCT/jKj5ajdzZPZAnDYopJST3PCLuWxtlQZ6+ToqFIh/ETqMzPgwP+TOj3Hbv
mdKM3HkyOYx9C6Wt9qMdkENyh9e+kz9X56mORW3Tm3n+udtgyxGEStQkpyrMiuN8
l3+/Ea/Vo2ONZ/C3O7cok1y0nXaaSenwEO0mHHMPE/fmInRaMs5GgjuuihU5OEkn
4wni//MEg3pSfBNdcnDEUPhYNFdLXj7TKjpJLkcuGiG2hhV7KWe4K/wat2YTiSxa
YvlCtZuZLQy2xJmF00MFnTzrtKJDRDBz0VqJMLQZiI7VtNcV7KhbH9WwhcIvtlvP
PsnHKUZpfPW2YfNRk2DcAPqC9oIXQLB+Qhb7O34omwGzjbeEiRTvPqUFX7zBouXF
rJJ8HWoidOuNlIdIT0+EYETD72dyU0Coz+J7VojzjmgOaOs9s2jsvleAsDTPNhiw
+GZdbcaAQZAr5/y4alCbAhKwYXWkrZLYrTYfaBtKs6ADuPdg/x+9RPVdlsc+1IO2
KJhb3rHg5j9r69lSlcsGe/oXn35x7KTMFdmCvGiJYje9YS5mVAaV+kbf2ASSbYzn
HlPuMQQwvhC971TzYqs7kJ+tU3D6rVvWFXXbSlmqEz9+813IQqwRzlGJqaWPs/GT
KygckuoH6p32RSfdQiTG2Xc6tK73yfScQNoE+cdXqY1KqyoicDe1N4U/Zc4xRR9b
4RPXopj8QkPfxZBj69kNPRIGxKerVEK9FxjoUbauYU8o0IrrJDoYQX5tTWFtHyEE
zLxNNNYxcoAjpF+RIYYVEpflLy8bqlfK5pyDKuhKbzDXt/uB+Y9kVE8iXtBoit32
UJg0bt8LTcU09l1uYTcilD2bYgghRXv/KtIT3LHxbFcqKRhxoW04Bgz+CzKqH6R6
mmAEETZTrMpY83FzEbYpAobXgmXv1HBCKIv4MU/XwdOIiyShBfH3wtHiTvFkpGyC
7LThc/x55478CQbggeCO4EmB46jMTYjW2mUjHpLx+CFUgDmFKsKyJQLcW73rkS6T
TzYcrg43OS+KRm3ckx9Ao4irVal3CoE8ZapBOZTDv5s8Mjx7hziVLk5VadY8KZfz
ajUAJgiSOYk0N1Fn5BGXPLM8tHp06PtZEwkxbeMW3kLNkGjtNLz4cvsWmbvM6LgK
X48xQ3ydEcddRD7kJ3RFpSl79L4rXQNKS+FSIdMrx7pTm36cV+a1KevblcXzLTXm
cVgmqrzymumqEKAVSHSJpa+UvxU/gzN2Q07MVivHYYo=

`pragma protect end_protected
