// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
iLo1u72lr5ZdHIbfG9bOdIKm4aGJPblsGaPqpzZSc1bHKfivDw5ofpZ7jo74y65BHHHPvZCbuD+E
T9+yXRM5yiE2bbA54OXcClPYYPHTLS3lFVzpupcfygNCBunNA4iN26rx4aznIUlKMwg+w11C+8Na
6e3AFFIqMfbxTZzWzUbw/g2OD3RW6xE+RQjAXFrQMHJcE4AwM/mo09xahsZo6yz4yoVyfh5uALaj
q/kOeswX4V6kWk73RiyXTmF+iw+k/9fo11NuO+C65G4/1ogW/5PCf6hH7SCz7A+ZHv5aKeGpmbp1
QKjojmOO1391oxK/O9rLj/VXo7xTNjznTc5wHg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 31408)
t8VZmKmpZBQBEm9LERo+Eys5H3p19qlg3oZP9esE6uUXBMq3xMfProVMEMdRf5Tz4C5rzpSBLJJ3
ONdVlTxCjkxV6XQAtUQJPBmK0123dRERctz9SL2wUM11lcMLNYdm62fL1l+WOq1eYFrX/66XD7Mb
QUEmPtZtzZJLYtha1TgsBJ/ZriLfilDmqQRXVeI56o6rDH7byQy+716W86U16pWxq+7CTJFGfbuT
/zczeM1qThvExu79lC+7tdXHt0yvVQO+BNN1hzJ5AcPGH4YH1sgSqqBAZ7jm4/mgJPBuvWiLvPrO
Y8wl0nnvVcPhAKMcF3fg7Esh37nk+3gF/tXnTt/WnAAmW/KZakcCC2flyV8a5sze2/Q6Y6E4eeJG
qYeCvg8/n/up6JOZEg0Fu3ukP+of5XHFz092n1mo1IvqLcVpYJvKLNKPmGCMjZ/JiYEeBqyNibry
7juNFkxmnop9HLjmTTSPGQwcMD1ZpjKI0EmL43xxlkWSyYLuZwWihS2ovwxL5ZjbdNfwJPdAMBV/
pDegyuKDR14cPIAnPPdtvuPLqnpvJsf82Z7hrDW5HWeTV7b6qTiYInrmeB6ttm23DfR8MbKb+/86
PFplnsCCV9sGPxKuFw8PYHQrxWzo9tOF/ptRCkQ6REBI6lsfW0OldfwSKngxc3iYAekHLjOuyNfU
wFz7xuTYDnP+1K+syI3yl1dtb6gKB5AA3DqKtTsIhtOplofDfaCPj0Ys3xhsbodWQFxdZ4u1zfr+
cyXxM00oBvxqwxeZdzWwSCELl0BxJa4iPSX7E4Yf3okzAQmBtDY99EZAggpoufHzAR1AjkqaulsO
uaN/TqigwgYgQSb4j/RWREK2BzriJmKRkP69xh0CwzOB0xF8hPrYULiExeqHHam331chjak9tuKJ
DeUC/jAJAzUuvcbbfpyjnBhSkxwN/xcX0FIbKTKcIoqMDLyM0vgyDVlRj2XiZfXc+P1hXjwdx2nL
0le+WosJl9LtX8L03Qn5WPCDQ9yap9M2Ph6co9StuRG91Sos6MethhAVcEbAqXPSGfW9lTRBeKqb
NJMwsz4KF/1Mmd8FIE7H5Dfrw+ln/KEcgvEqvb39nX6pjjpowA0CGVwnPpmSTktOzxG2ZPKewZUR
B211wbJF1GRULk8DesRBigzGyY+moaOujAXv5Jgmh6LTe6mN2FE9e/bs0idMJFgp+MQQVw4Oll59
2wx6x/HMIZWqJcN7/Me1ls7DsAoIXg3agM8zrJIuEGtxfgNLIcbCNKz/1YQViR8sT8lAlkUbZGD9
rYyY+I2/6zKsVhDyF2xY/ZPiiyEfB6OA2FjngLx6AiJPPZGN9P4tPqyql828nAgXzMFzl+csPril
fDRbn5Y+yJRsR0zoyhmZYGJhX/WzBG9TNS6EumZ6ckmaiGYtZD77fSp7A9Pyw4NwduSMqTQpwCNf
l6oQxSOpdFCrQTC0kUxGwLN+PS/HHzcxzTIQslMYLtcEgpdK62U0mYOBrZPzrrpAdquVevvCDh91
b1Ro0BNq04vE12Edog7qW9wu/7WMSp8egBnEVtjZrn6dp/eBPenwUE49prL8SpN1BpZutJdMHLgt
5kURXKPAmOdhunxXgPo8asKZMV+cp6PKCez25q01v/1SojsWBb5mqrLJUtCtix99sf+yMIoNaoeJ
rOaAR8xEeFoj/hQGHRRp50Z/TG7N7W0YoS/SNujw6F4abeYkpqaI94RqBa03CKaYonIoZOy319bN
HN/N2w5aCy+WNuSeOOJZgYfhWkxFgGmy7d5O5tq3ZKUkWXlaOx9soljbsKpdEHHGGI01fSVsjWeV
TynbvnxX1otMBAqvPhrH4YXXMIJ99c6LbHXUMCr1Ae9Srv81lAxh844sTIsgSXaPOELWEfbHkMr5
SikBwDygHmCL2wnQ7pyqt1OXLcnDl2qUOwuoU7l4Ojlv1kr+w3Ij8VOQbwhLOa4cy1N/hOB1nFz9
4vHOr65QE7kHKKThTeEoZCNLWvw1pPhluuJzuQ1an8wQ79PsPgrIQ2tV4tylaPNRxI/2fyajxzrA
zU+KU3TZbOrTso6fyN090K0FybwNZ1mGwj/IW9Mk0E5WbWCPekxKXeG7TpcbKfJxPI0C6gThv9re
zlG/IR0mogPWqWX3b1zNuixs/b55Xms31HxPJl8cb0g38UnTWAlWt00tAEcctHx03XWNgK51ytR8
+dt7I65Wa3RDW9GdZStocLUe9DblecAZB1lFt008wTEGe0+nv8xqp9la5vqqHmhkqc6Tc6Mgpn0b
89cQwIFuMw3QR3EKZyn9wVu89tt4G/ZqBO6+D18WGX9vHSKaNeFdy7rEBbo/BOnGzDYEG87ciAjj
MrviZBV3OLUWdIjSUSOwIcOvXzcwCI89N3Aqy6guuNjdUNL9gGcL3IgZB9AXIIb9LTG66MxkmpCt
j5PscNHxm8NFZFKeEWcIA/7RKq9C0UmZ2EGnn55kqbASpm343k2tJ0COdrBs2/QkUyaUP7/ODTLZ
aqFRUVO0ry9U789oH54xWYxVQ220JqBfct9y8E6EWTidV4CEmmsczyP0tUZhK7wF4Cm99TKf2XDn
W4XmdmFjf2c06BS0nrlTiJS6Bxc6i+wG2lw3wIykoj9Z1aYrlZpZ7nGT1OCPLkK8+uJSDqlN2PB7
kFKeBoNRdLe8jLXcj9Lku//cRN+lHXqvHwn5uMqIgRVd6L62B4u4MOX3qyE/X0ZlrsBfWDloVIBs
9Oycy2/VDvSSzytsAkEbsX8Mi5STmK2hfzbWMo8Xhobi7ZUZjd6Jy+cY26H/ckRbr7FfofAATkxU
wOHyf/NfgKTqTdfITc9f6r0RyytoSlilqZv57OV9hW52wi9mHdVg6QwPBT2e+GJub1/xRSEltcei
nO+k41VvBEBp+AYNjQrl4u+JCGt7v15I+n0SyCwDzBQgLJrsjXM0Rjkkb99PK+oH8rAWDtHVB9GO
qtXHdQ7pU9j2SqToef09BqDfnas4GR+YYYxLWL3gidvw2dQsSRXl76OuflAn+FOhgOMZedL3kRFj
9C+thMx+DKvmGRyoCt0g1G5zlpaCy/8gShXNX41D+ejcZ9b5OHZbIYoh4qV2RBPackXzQhN4L9YA
nOu2/YPDokqUJ/Bj+B+Am1AT9fwJgP2+cnk7paRRu8P1blE4yFijb71Mn8hLSEf094oY8llUP32K
UNrdMMIJ6x+Fe+eKbY4UMh/BSVfIh0ExjnbP8XzXMmw7Y2G8dE4EK4jPgAfeHHQiOE0e4jR9iemA
GqSXbj17G2bFrCbRxqijOf+HMVXB1OkFI/lhNW0Zx+G9PZJRW3PUdofLAd+Ybvs4LMj6I9lde1OH
XYsHvRUa8FIJg0VdufWAaB0/RN6wTXp4XZ01KlaIpmPGLOLNyytBS9Ff8GgaLCO4XHYkH3zDOFD2
1oUPWBX6/RrNTzOPkNHC7FD7l/ntE2H40J19c+1s/NiFQ7bcNXpGw5RzF0rNZKtV7D8KYzYUfCoV
n74ftA8Bg38VzBAzFhK0cIOzJNNC3J20YCdQ3i7XyCtBpPDybOqQJhfRr9fZdQvD9H4jpA/YAhkH
MtG0wUPljGjgGI/+zUWeg8oo2D9fYH++XS+oCG2vxxhrTwl0S3eB0A0RFoTP+0mSMmHSQe55ITEU
8YFkvXle6PIAxhrLdVW+nXkpeBYSF4+hcY3OiVrzeEQkOsoUIsj5yvZth8kKf14TnQfNULyO/sF8
qZUhC4i9/7AZX6pLYXjbjOYfVQKiUWSJwfQ2d8hjSTntfsxhgNpXNvPVnm6gJ+GJnd4lkSG9pddt
PPW+26pTStOAix05k/MyjOJxk3rflR2fHinrS1phY2HCBfl0WdJyg+KKtGY6H6InPum2LTNWzLVP
uCfb1K3a5W57dujHKGZTQY31Y6PyWffIqEcx3G1CYk0AhOO8robMnuj7IL5EcXHOh+tIKaKlRcr6
gf6S/2cHlXDQ+jsrE+xsN9IFfJ7a+7IfEriOmDvDJ9DgjazVBf82Hm2BCVSZ6alfWjLUqRjod7Zc
MS5iIqoAyaIJH/93jkt212hRQTXcSufLgA1o2UnO3lgWYGp42/F1vBgX9wZLPvhshA0vpJJoj8NH
tWAT9AM8xoJVYLYS3tTpDxwacTPK7adw0BTa1HD8KdCrgbSos5VDK4n5ue8o59b6ZQdNVgWP691P
nzhWWBUltrldSY9JsH0H4WcHOF5g2g59nPunDtyToYXpHmgfYO8cKS9qKbvPXaTHElcC7PM4V7W+
LWUkxm002YCSuHttr+ugEWez90YoNs4fsPozqYsoGbhtPffUAe6MqU6E9d7HVcZsbiQ8otEQt/VL
ggfYBo76fwjloZuRgLyNLJuZCQYMBaqz7Q0FFcSvrDqI7FanTu1hm9jmBk7WSnH+gk7tRfMkGS2d
oXQ+jI5KZDRWqjtNO+hHirDj0mACgNs1zlIRKmPuHVIo5jTcGwcAm6dTT1YEiQnhY9oG4imMrJqk
D4qn90bwa0WzzwG9MRvMZlc5xpHmNrkugwXzqW/bpQI9nkpi0hgt+dMBvt56jqY/szHEOtcGigog
k3mzJJaLSvUrmS2Wn5095VIBbXuZSfu7XGhWiz9EyPi+BK5aj/PWASk20q650Puff4fV0R1VaPBM
KbLvg0+vqteoUQHGsdXnssh1OhoC4adBHBAoHB3xynaLJQHSRqlFxqxFg4ybYptat0ZifjrrCN/F
W7Jj9d1nQWMhjgp2y/DeWXFGf7JvUVhY/KTW5l/NHmfaCuWMJsbULxO7rb6UxJscvVCVRWxhpmYx
jSWv7J8IKQwehxokkvBfNoPHsE7UdFMG0zNaliPtG2FB2tvGttBqZ5BVCYym25aHk5fwWLrct49g
OKKbi0xJGFzlVm5BvB1JmHsYcIFi43+RV06hgxrkQKdbuvgo7om0/R8o4wl+xaFObgGSnDoY4q80
tWhQ2KLBkvrF3zJ1JT3v59/jmLvouyBSJDWQERTP/EENZZ6EyA2IB9dNLoYlMkdAXr+jdCc2MtLA
a9IdhidjnEfIyKmkVaGw8DDoNcnu9CFwj4m6hRRxPIQFkAc4qVMyg/o+tipKc7jP/gIA23fZQthk
nOPjWliz3jFNEkZvuyrdE14591A9PrlOkmaw7ZeEIfqVYue40pGEVLeWMXGmG4drXANX3AstG0xi
PTtPvQNkGFVdYAUgb1OAK9Gu3otTszy0A3Jgky6s4HPNJxdAouFFxrbAAsMbYlIR1jhlV4tt8v6Y
bkmzd6N3PcE7/J3pauXssLl6QYjQNgwOqUJj/JjGYsWO/7kXQksfOLlDyOhoxFuIw5RBRL3G2qAH
ct8tvitJiQdwsR/1lro5hHmfX1JPEm6hLKfEPFNGuqhdhsp5w2CXmOmpMbRXPi3J/UsyuaLYBW2O
/gKyTYQgOfagrBUIFxFIvVYiFaOqcHYN1/ZuJoaoS/6Av/fuLobV1DNcrVcZsjuzAQdvE+HfX3nf
0ZPOWDRACWtpnCsdmXvROiMP+QbiQOGL3SfSRFwLoC26h0tyxo3JhjsdeKDXgzScYhFsBtGbkR4R
g9JeWx6V1S0+iQ9Rs3omvHNzQCmMLyM6RHl3KusGulJkWL1LpAp1wth8uDTp2MVPYP8hVWvKjW3p
SYUSR6Qm17SbkwgriIhGMTIcXaCrJog3KOu18hB95ZppQbrq6rE+uYYJIEVJjfW+GL5eHbCXkRKF
ifOQQwxOZg5niMbYNWi2y1F7nrEWJWZ+35cBZzY+erNIfGAqi73okHFD981YF+qk4do/uDlJbx8Y
p4+KL2+UfQz6TD080uoQR5w6UIA8DWuEse+FRJLvazSlVs5wOox4zCtjih+cd62Ca6Y9puykM2mh
zyQ7yc2lTuykbHHmR3hf47LxNrH88+lyWfh3j2jGaIPVcAVoiI1peHNRnp12Nd9Uop5LO76dnp8t
6gHE5mvYWX+TrrLz/g+jxKolaD2Nqe9g0IINMdzDWunQODhnTvcBpAcymRQrKWbVwfTjCjwZq1XS
96/pwcwl5/IdX5TIIPohpAxSws8+1pgx5m1Ux1Ypicgy4CB3vZ9t+mWDlpJaBIKZDyIQtzOEFToa
9XPI8r7q/mZSQRPrfQrlKKxzI41CWH8IvnqzhO0qanmeZZjAelnVp4wtp5JBvrKtqquL8tHBbDll
mcRKgilSziacLTHBvIOWTgn8CmiU5eiS6bhWiOkAQR4UrRhMEl5f9FxQe4+oZao7K0K5gqc8Kt3s
grkRkq3Aj3lmoDTqyih5DokiPjKGxN26RrNfeG7xIZB4914D3Mynek5lQglHgWKym0IBF97dHsKd
ngQ51p117aqh/XW0IWrOjYnDEeU2axnApEuTdk12yy2gBS3Pc3tiO/MFhLbsYHFkIDEG++4GYUeA
Q9uIcTqfAUFrTA9PZxH4iO4tzFFT7vY37V9hcMEFNPPzLrpiEKJobUAhblMwIEC5+8vaW1J0v1uw
/SB7GtsjSBDueZfKx8tNO0q0pbMWKWPzWuBM4sA51oepViHGRoAiRx1SYLbGh/9D6+bZoa5mm/Ag
9vjE6Pqvx8Yr0A9Lj/QE6J5UH+xK+g4nu4a0LyhwC6gVO7ZmtXU2X7aGTrNvwdfy3coduBc5rAA4
Zdko8A8J2ogQzekVagPovV8hULGCf5ktttVxZkJXTnHb4wMoU78cm75W4BFUW28gJqukLedB/bvl
GRk9WiaeXWdWfYbvcMARTqKmhnIhI4AtC6yWZNunHOJnDofBpvmm7rMVTsU3iznGwozqcE12LC+l
B/hvw9lFuzUMt4mcPCmM2X6gMo4mvdBOTVYS7oNzU0LU43CEzFXbav7svFB21bz8tpLdati1Bw0G
eNKOO6l8ci8DKPbCWbtUW8Fz16gFJ/eNhgVPf1nduc67DeW6U7U05YRYTlQI+babrVTJ2NtO45jB
nzZV9SzapPxOA/ZaUj49VtrvWOvYIIOPiqbOtiMosx3lASNffa3EGTBAlfFtNowxIdrRBKCZya36
ghy16WI2dktx/yrIjh5rQ8cXO5NxK8zGSEr7yviND1JuwnnIlrxQSgTyHBcTGmb+I0+J19EBBaLn
uQgBzUJMGhvAxmeej+2rPOcy5bEtT9z2O2c05t9KqAGmHNgbd/9KncLE5QEv1IdZgB+DRLZEMkCJ
a/FkX5qbnA4II9u6uXHkpMFaqHX41V6fgWYB3uw/ok9FpGsISCd0wrkkp0f36zRPh/XI3KKcDJ32
/vgSl6J+F7TVLobuhGGCIoCpDQNuIrK4Zs5QqgjOAXFQbmSTXKSoGPX+RiA1872GS/OC2AtryCdr
7mW6s4hq1X5iUN8iTP7D4KoN0Gg8XVdjIJBo5MpcERo0HQ59lfjnizNS4Nk8hUTc626q4qp6UPh1
nu620GtBnrA4707gYK36FwJOnX6OVZJXSaw9Xfrsj8IFn3RbJ7AofAF4nVRQn5kTalHF5/DTmsIF
8nnbWVoSYFpFRi4yB/Fv4PnANcHWlnSV+x/xwPmUt1LUT5NpARul8MJ/WidkkjjItIBC6izDC8ke
R4L81oaGFir2hQKMd6+29eQnLHN8Njfw/puUi8BLEHp1HE+wxcdi/fsgH8odmsf4lT8ThbIAwtgl
PYes6e0aOP6i4btKDeCZu6cNiXt5kMcjUnyWWS1p2uzx8vYBnZR1zrMClwa9Qz7uWkKGq2jUXFLt
OiVTHMcdUFDHglHtXGVF5kQzBvVwDq8mfZDUc/3//lFu3Fa5/R+oXz480ZWcZjW9OLtlcytrpWmD
jVpummNggDscf9wpos9u7mPv4QEI0QtCkXCKwYxkyuFkvYTDkRBw3LjMbP3Szbicbe9wbw1vNOW8
Uy4DkWSuvaFiZm/qEGNciSSyOKNs6blcMXNrgAYxsdeEqUdLO/cYnsKdoFU3at+EpLToeUn/uPxs
qKLkjXkpnyl0omucZTccjSyW+SkCr9HlMmlBIyA/0jv1o1FAXRxdkwXHAS1Sj4XcsPxuiAWnlCe2
rCNeIGV/v0ddyK45vc0Ek1h7QoQ6YSERab4sFTCkDh2yfkiFkkih2YuPnsI1/q9sR1kRNNGoJZzi
Mocmu1G6prUDUcjV1I7q7bAIM/Srg+ogZJpmDgAR650cocKhH82ZGTXkGoZEAGtUYHbExe2XpVhf
K0TkoZkt1ZeliPpV8DvB7UFqqE0Batci/jJBma1wD0OaD8Xu/Oo785qUDZHUPi/uI4ECklnU8RXw
9DoqvrjFo1nU2TnGkeL5A8I8eWSL9xICSy9w0DgFd7e5v9bVuavsyNGbkcAV9oINKspRWpY2E91o
uNuQhQb3YjSUqNCEo5VC5pEvSkbCr27TpY7BpjpvCNW8/VECGqxj0L6VnbnR9Y3qAKgD4gJl8S9I
9ZlADbQFFbhWPpYICHFIqVRHM3M37F8H6vUeRqdXn7we9RyvWaYkrH3WC4AS/A5vIKoyuiy1twcR
3rQncNDy2t/QeADeiVWdwcQrRklzT0L9+qrg+RWer+2ilyYqEWhWKQeTbsQsZy2zg5RK7LzKFW29
GK3tkqrHFRzMi/SfDE+UzYoTBX90NCI3tUX+buGeS71j9BJmERVb8YG4+FW44DqlT0HIV+8mSXxA
zqd0PWVlN4m9D8znbQZ2/6nmFxABomD6kpGLLK1RK2iTvfzyH4U7cYevhEq1C3Gzdni+hxupmVS2
yiOPOcwT6eJnT21Wd8xVxqx8wCAjzMCtCdqQWuulHICr6x/WjnSt6ww6N81mYMfNssEsMhqIr/Eb
EDu/KtxMN4MkvH9Rp8navXJHaAWlj6IRuoqIcfPALHZrtNthoewbT+HClfIcCVA3efyBNkxDt99v
GHFI069vJfL5XalgSUMYKmAVoqaov4LSbKX9SwosHbceXu5/G38mkTL3knxR0ET6rH+FqnwnsB/s
bIKMQ7+ScfMuqNR3U/21kJWkyuPkFSitPuEnVLZ8kNxm16dNScIuM0uLzzcwKGZh4UhVaViZz/JD
zmOLyoJ0Nza/0AATizwkQHY1+2GTtPh3UBCaqX7Ysx78HwNrxAVH+KX6yBOg2rintYX/cGXsdjSG
dZ8ooKQwArEvLTbptRwETkP+Vk1OG/dJ+Gu3Of5ISg+Sthtf7mf+ifnP3fkPI3/WDhdGevpda5Tx
oEEGmaJF6jQSwAmKe+bBB+sslMjG2sMcZlfgd3X3J9IEOlZ0viJ/FNGtYuzp+5hRbBLJp4bACd+x
PlEpoP/viTTEBUKG/Isg2W5mtiH53SzAp5u9UBGHhSlGZVXk9+dCzKCR4ilSNJOVOvA82UNU38FH
t1hLrafQdXftZlgFcQdN8saltPwZ+CHhhSsPTdCfUHhvbxcqRx2UZySAWkKANZ+Y5xouCpriOfo4
poC8TZnhKirctUUvxCAmkAARHNpVljPhxO/4jld8eq/9GIh55J+LMB3AMwDqSeO+iZYcAlCcQjDV
p5lll7nc+GwEVVgy6sRWLCV+Zn/WozkRNIh+Lw+lutEuXOqiY/1PWcfNdJ2AUj9MxTnJ/Vs+RkDb
qmLOurmYuEvxKGs2zOA6nbdGKqzv/gehQS8i+2DTp39uJPn8Vvb8PCzheGhnv93WBBrQb2ZRSbfT
I+tM8iO1dfXNw75gERsEmHz4NmbR5l1qck5wqot8Cn2oa+I3Lzfcl+GhVSSVSykyKLRh0ARVTNV5
PjCfAmuxS+0lztF1RrJW4DhQp1hysw75s/SF4cmkauoUQ1ObhCwXe4HbOr6lPEMSYCePtqs2Zhpq
4B4kXzppeo/zP5NMl2mgRALDpn54c6+x5BF4yRz4M8E+o7EfENthYImJCSS1fbOcwTIWM950XS7+
9xl/UxYfqnDnuy3kOyaiFdz3DwlHfveoRTsXPh1nh5Td1ipeySmWg5EDdWRQfaB66mIUpLZxvGi0
m9GWneDWHFLEWXLeX8x9/0GSMlmydKbA4yTi0fmmIgaGXMtC3ucwUT9Tn1mJ0gwZ4n9N7gmvTpO7
ZhVzqRtSuipXGCfR6jrtMXtnXAF8nidm3btX5Il1l9rrvjUdov/QqXPj8OUM0uMI+nv1o3tb+23I
QnpjluDUEwWKxGAOxUyk9t7bQh7fdSorD126wUAo7zfCblBS6MirqvproiqhYP28IZll+DskY13t
yddUwPyJw7W1DLLsaQ7R07N1UI3R8e1wvThK4bbUGTXJqGvQTb6FJljlpVqHbChOvydb45tKUm5o
eeS6JLYasuMoibf6LACO77qmaMeGDKjhgcHdQ8H90J8aPRl6pKlUMOSwC4fMRlkZ5IpqkWS0WQ+B
Ecsp/aNdA0M+8E4vtJiD4xmzzUSM8rlPVY3LYBxlWZqE6xrwdQIdk8wibMUiEf+RwnQ4FefpSEKK
V7ZvOZuTgS1XnE+KoH9p5qDo7/oK8ZWCpuHv7XR03AlV/mT155dHU5BmaYzfzeKlaZiINX+oOsEf
JcutDj8HbofYoQdb6W5+yy+1KPx51dVyrgW2Qtuk1B7oKPbkQG1muy5qrNBw8OiZpeMIbyCHldkv
jAlBHijq4eKOjrZXl5hTcPFCD1Z+u1unguRIQtBXxDMt5i4PzAqlyODNsSIRwc8rqlkT3gN00jBm
+/DpH3MD3+020g42X5Qs3dPHMiE+axR6G1YW9DY+qIximBUz6jX8womGR2scVfB9md+HMZ6GHmt5
tmnkI0jZirFmy4h3lK6+HGaE14YJ5WVAGvk24rXr9ygmomCcOq+wlNtnTp7gyTBEIfdrQfPDDyWo
gZJI2OSqvSl15gMzmSm8PFBKsfm4UWy90ePcZ8CBZFMs32o5/kQNY0+4tq1Z26F0SfI7R9QX/deH
UFiGljYL8RL/wumBSjVdlweFMD7Ro0+sx7Io4BPvWzdWJyZLZw7tYTheBOjbcXj9vIIYDyWdsQP/
6EIXgl8V+SLylPiN6H8fSLSjQ5m2vx8L8eKVZphuNHx4siXIGt7tTZo7FGdRLHufUUcXXWygOgtP
ZhRjhTudUleUtaTpbza5wKCNowIgZXSFVK/427fyaYgzYB8dXRBYlzvWQn86f4180fKfo3kDcFuF
mIJZPq6flf+0gpywBTLGP9pzfzIRfis35hJ5Sgbqg9p4qoGOY0gyhT9ff88/4i0Nb41WDz9IHD/Q
QpQ8MnhHfFzw7cMc6SwbxbLeeZNTz1ArCd377wXKKT1jC4US3MEN2ZUPXpMPa9yoV6o4GHMNv3Jh
D5k0WU0a2aOjgoro6S07B6nd9bLD+s1Vuap2bSuFCXkD0dP1BZlCTiPrGhOlxU5aeuBvmuM+hW6h
lEpdL/rUFJa3sOM51bq8KDHtK6yC2+JaS0vCImup2MLKqcF7ZNWwuJkeTfcBfAjw73h3BQGw5q2I
3Y1n0t4Qyq3NzFF0+K+ruEbB4ZATGhP2XN8R4Xvj1zxkpfRyeWHFCtXeSkLINGALlRGPBILQm1x+
hZDlmXoUDYJ7c4XZG+R70WKPCEr/AHgcTr5fHXax/0zkxUoUjdKjfjlsB13Ku+e7xizyg9lpvSgo
5WClSuLDHLwzrVbVz1tBppERPUQu7wEj+JXNMqEP0v5pGmMA78zXVFEViAg6zW3mRrRn+P9LTuUe
55V3DMem8gzi7yC/oz4SmARZEIaoR9BUgQriNMxnOZQFIkePFlYQ/F4BWh68AuXDCZTJBHaUobQ+
DLpx6tm9pTJomCjyexqeG4bhiHHy3VkuGvuL2N8D2WeM27kM3Mb+DVy4wTulYWo1Ewpi8IcUFztd
24a07FXqvxlOEgRNiS6Dw8Dyz/s+EegcXb8InUH6krtKZHhiuButt0oy8yt/URO1HMMmMZ6i+tEO
ijjDxiBb+K81wrhx8dZZZ8cwS7p++NpzQIJj2CdfeaBz148cLWRngknfZ298UELTtUTcv5IrkyOh
P/fiHT7Cq0PkBExm9pmsENPuBf0XbVrla/NxKZCXgCxwJDmr3vElMP10LLEpIqwgg2YjF7AwX/Hv
GfqUJsIO394iHyEy5IIQm5Q1zg/Pdw8NhmXZn1RuKjQGb6Sc2k8Rzd8HLwcw7KeszeLyEeR8MH4t
a+qwuIdY8WsYFX7oMPJ2qa2rmi+N99AQJZLJdkvFhTuB1heQMJxvQhfOEmArUsmbQZ3S3HZ5TzFw
2TQcjU6e4m0xxyZtAxFFBLHJl9aEc61PqAhtsn3dL7VgjSLJ8EgRC030jM6jU56B3LR5YXBdUIDB
LYBRnnEe+wBi0N0NQqydKJfhS6Sya/KevpZMHRdOrPhnbWPrHLHjnXLF6ZJ1h2W02ilRfQKGA1Op
09PSs5IZnBSeiEiJG+rFIzXzqNUUaQSSJ0vCCb04R63P/RdJqOZAAStMPTnGsQawMZRI/Cbypl99
OywH1CrrkE+73153hmmNjCtmmL2pPF6egk7T/X56WxZ0y/lH0Z0ze7QQcJgY50LrZaA0C4x2bXd9
CH7khaR+rJkHTO7W5WAA99fkK69X94xfAwPeT76wm9JYtSdYkv8EVSxIJK17s2UeG0bIQC+J1paP
eEBkaQgCFp6/yzeG3d0cIJB3l4mrqKxZNhdsT2MUYFTwxEKgrMn8PCB8Oz9IXsdG/ceciYANJnP5
j9NOe6uUKkIKMHCQ7K8/nxTJ0ACBtP6bF3j1/A+/09pzOOoCwDWhNn30sNcYJtehWuH3HeAnYeF9
iTYdMqA/ujqAut78/wkpnd/0/kfYxrRpx8dODQNgFx5b8YovI8XHIupI3l4/E9c4ZiBc5DvlrKex
rl4btWEFyj5dnmlGnUA3mbVWD3Cmzpcz6nED6jbfvQrQSUC4uiXPHMS4evX1LoNqpdOjSzEfHLpQ
I1zVr/tsQr+RY2GlFEkaw/BzlRIAQMkYmeX5Sa/pyvHwsGCWYtruXUmHoeXyo3mylD7r87xan9Eq
BTXwEfMbb5mmKjIh7nDqfegBsiRrL3evNZL+oJCxzUpFEQyIbXMxy7ZqVP10dYLbcC4s668AxZLR
b77AcdbrTQGPJoJ9mivxlBIp3UqaFiPUjO++IZaea4u+usgFQ5ijyqGj7OsfLGU2qAvs7Sg83xNk
+ShzztBwGY0XgD4JUd/1VYrRVkSuTyLpGUQld2gT+kQM3AjB24UQczLp5emxO4V7CqqwJdqzS9ND
DBADWiRhaC+L8v7tTAB0j8QhKdZY7ltqJm4DsMsTWYkxkNQdOaTGZhd2Bii055+mblvt30QCzRoM
+4+sEi8IOtSgcPMJgMBQJ3xeQ5x29d+ck5MQcBTPL96KGMFzueCrVcEkSwKWQmdEaNck1jjiaXgq
BmSd3Ur0u/OGmVf0cHBVr8Kk6oRzMKKShnioqJnNzD/O/ei6p+ZvypSqsO6wLvWCDoNBzP7Jamzh
jeZ6O7Yxd8gzQYg8cdwnPY3JAGK6dVQhTRQX7RDHOoOs/ZS/vfN5ZEdFRDL27ZEctAcfqbM32QTu
oXkFYYpN/wopM+o4FVrqiSIjsdQLFlha5XI/m8Zs8CjjM2gpg0I63H1Gh1T0Br449Hg5QrtDSo3J
4UnRrQPo+VzdoMPM6yDPxZiMEwzQHuzP0fvTNSRcpuFqtEBTuylI0bnnUfkFnoqmqJ5sgIaBzyDX
C/xyCvr6UgMRxuh7CXazPS123ppeMj5CMEKs2mNqTH+B8HXsGCpPypYPGcQAX//tHQ/CiGYKU90v
0ESArzty3nLtadOMAvx+mQsnCfj/JeqttezaDwppAZ5uxeR7RMJvxTStwqJxv9SRP/GMLoNJmbOB
1vvqvDLctNaRE4+ISkHFMh91YXcaBlb7/EeT96yVc2O4agFFrVH9T1UHyPazBnj0PVYJ4+0dq38p
aheFs5xiuEFs47TaqDh6pYWMmmEpu7Ds1zalFmZEmMSoEdYf7kLJWIAaExUGNLn6PQE+Rqnc+Yzw
JW31ZK0ODymCY2vti5eyL2rsgvV+W/HJJUfp0CtWSP7myQUSM16le22O2tQwLqAL44AHXPghIpz4
lQu6E9ow9KmAKEg2Gto2o4v0c1aQx+f99ANTauQx/OAZlmm9qbAb+dxecOdZenaDsfGzJmpSyKKe
f3aNgzGlD4dBG8PU9wRwQkb8Yy5JW6M3c992Je80kdfE3s+caO5SuZ7uRn4IuSVN+vIPi8Ol4BuN
m0AYSdoZrdRi7B9GowMi/+iWm96biMhWt7Jt62N3nYEn/Sn3lxI6acxpv+Xc2YA93iSYoK374mE5
XRkO9Z7vGpVFp7StT/ri9R+wb1nWguhMx3Y5r4zm4e9tfowL5rwOPKy+e6x/9Kl1Ck4Dq/JQs78R
L5W5F4koutuKfuinX9/ankbDm8GZPYcUoO9P8idJugv/hyN7igabDXuMbzvtJOLn+TpQrIRoo81L
tpQzrVSNgMUjhx/b5LcezCn3vF32gagw6wghjiCQX+NuTrFYyOOsvpqfBRxIO6bRqc8CTx7z2C8O
9+Z3nEof9rp7vH2kLtMM29Vs0vWvH37EAbRsWZfQTSbcbrtbAVmAuRAN5OAX/o0pQIJZTDX9CFhJ
f5+jGPBOk1eVD69yD/95aIwBMudHbBvOIKmqN+X322kecb/Mh+pCD/8IR0uWkfy7pOAqUVsX03bx
d8siX7qC3g5U5XQlB0RmGD+j9fJ6uTRgb1vzrPtk1dhyC98r4VJ7Y4bwM1w2anAx6C9gFGGUxmZW
9tz9+w7pmUmQ61vwqxzIMSyFV7k31UVQZFwgYzC6RAqgJ9cgDjmZe0tn80riEIjFc4tShAz+s7TK
XeF3VPojGxqfd+aT0IYVycNxGBSrws/kfLMOunJqu3EYrKZ/uI9jFh4fEEUolr5yHwOnSQ6fecxS
PrhpS9JbXLFMCPGc4JcEY3b6L7DCVczHjJTUE5/dPwgHQyBaFnvtEVtz7zsrJ82Yc6WCgdm4RYWK
fRQ2eneuqTjbD2dHCDJz13iwNMQtms0RUUureYxcimRNrZBlcdMM2WL+e0A9wzXZL4qOIsUiHoch
buQTDpx5MQkHhbxW7NWrCLrw+JgSg95JILfBXEh0E4P99hkgERpzGKxDhmWjFJdC2xZFR4rQBT3U
qdS9vds393Zmh0mws0MCAhslzBGrJ3c3/srBth8F8XP6MC2mHPS6XMQuWT6PLrekC7LG5Lgesiua
vV4BLC9Cz3rXfGL7AsAr837TlF4vgs7TZOYTzL0xep+nWEf4AFdeVkMAvPFqGSryuRfJWCDUOuM0
ZdPlrqFXmqmwWHM2I4pNWLHrvABq72N+j6EhpY7+CsI5uxnowkdKRKQMuYZgAOuv4oVgVg0SA740
LrERnFHmtUbkJN9vl6MapOxmmaCRGo+2CfwM7mUUGSx9WeGsojhzT4OzGpzdIkheOK8NUKO6/iu/
7uyESbMCZGc4R8r3c9VyF71JIJ9YcY+AiOldUbTewtAf64eZQI4KcqZqYCNhWyh4Kv8T7ecNKo9j
kSs7D5sLvuRAC1jKfrvIgFXRBfxLO8p20hyZnDEnHCyaBZrblL/cnyV//auzlGinDwNyvpzt01UT
LCZJUvwgnRCu9NJQiVxr8NHgho0TZ+0bkTKv1chUhW+Uo+ryWTKZMdcrH+UTIlhG2k1lvPfze+pV
se7ZqFAz5BngdcDj52N+j0RYTWnDL/fukEmxmFWxXNHEA9KQAIi7k554PAuFrEnwhIH8GLbEkUT8
eE1O+7671OTDDZmxjeHDVKlREvRljSUvCjmtkS9MB25PQR31IiZH/HhXtF68USFf/nMyspwh09Q5
QM4rZBtArzt13VbZGoliJFca18CZsX6qaoUqyFJFZVZAw+7gmne+ffVQqrA3838dxSck7GESXBmw
IcUAl3mPngS93jFBFW4P5QH6hfIxjKmZJDHSC2aTImFL8Ky7xHgqniGSr6XQcOb2uP/kCeHVMekW
k5hVdFdj9j1VtIoWIhlgWAMiYgNAIyCzTBF00F17lDGM9DpcjRruUcUhzdrIHWOalldWQMqn6QVJ
zLYirWredIS8o0ipHQ4CPxaNdimpDMCzjEgtWcmnanksLJKkEhaAHeHHFZuVMQvI+Z72VTzRcEC1
zXjQY6Y5LhJz/RBBmHjcCnbQR+RJCO5l7kL1BJb9OFZLjGvbdWBSp+HXL8HtOfjRxQRNti/sxT2H
dsSzKEJZEW6OshV/lVstFydAulxihda4VSCwpAgISZF1cg7b6SU/grs3GswdLSDPjfG5HXY0F0aL
FMEtEuGkSmsC8bsr/PSJHqvkgDc2zNdoqHvXVe2SnC3Wid9v8uwtvmKVqbFj+8KSSXf7ENor4dJ0
vnTZUWXPbz4YHtCpDU71ldMsYHZkCUwF6yirkaGZCy7IP7q6uACHdCbTt9fcFA3ht6GviaNtUvrT
+WXcMdsmEwEbdunpXDrSRtUi+i2P8HZIlUM8wjAI2w7HdYmEYDig0RuEbdH85jJ/WLh126ViWeXG
8LMssDaOZ4ZH7a5ui2X7TWmERBXCW3tJQJOIPh0sqdARfqhwDThx/Wvlk0P8+KY+XvLpOuNClmDr
h3XeOAzZdRHLQQz4aE43qlTsuFXlvVyQaAE4AfluCMCBl70ZvLQNaQRa/DsRMF7HQZsyQMfanHF3
gkNNbL8stgdrMZyPdTIQVhu6zFM2qRAtpA9+x07DkFxLCAlU/K6kXGHUZv4sjC8nKkatjVLaJH8T
PbgzPr2RpTCLKJUzgyAZ5Ow3moAXYF4zThRZpdonN2V4TPFsaEMJQN/iauuVEU6WxOOJSweS8Sr0
dbLGzrLLo4cTXvk19vKzvKiklj8QtDIqKHh/xURhZ6/QGc6/yHOFkHN45Iqn8bHEej0JbEgLgNcW
YQjYPy6VRcx/f6SAAF5n9N7NIIe0vDsDMWXdYtnYN4+LY7/JKzAOXiN48mRw5NxuWRCyGoZt7xm5
DakeVjcLQeQ0IQ3o9NFOMlXnRCh2ASzWTzcNn69UFokWOih7o8WzEHLLyxpIreMmtKufgODP3AKL
yOb5LympQ4uQVJuh5hs/5fEo7l2Dwrc7Yw7xZz4YXG+4pu4FTGhvEPmsOegTWzamvBoE7lpqZAvz
D78xCJcarWjhIhyGbNKVCOhY/EGpXdwbQdqZqxI5DiPPOHp/wkXJIMXdWDn8/uCM/iRR6PFBbVzk
uL5MepzG6tsZv1VPFOlrKt6NXzNLe9xt5IuKgZP0gWoWg6ALR/zXCWUetf+345r0FNlc8J0WHnYU
NXfFJz8i9HOYZk99qkvD/Fd7cuxgxiLhfBQhmWzAoCYBwbctB5RP24eQRUidWI3YhxM+/WZ6eJGt
+DQb8t0cs0iTM6dZTJ3voegrj9VZjg3ThVmvtFVHj8F10KUi0AC3M5zjzoa8HpxuxWW43LdK+He7
dB/93+rHSxq4/bRcZz7MDTTmibdUZCacsrukC34a3WpbNNXv2RSiW4uBv5ACMrHzdU3aj+hW2QOc
fEJs4YKRIRkQhF+YvObnKb06ZP+vErVtXeEhMpBXBD4sgiWZym/C/+TlGVR20tQP3V5r3ovltEOG
41wUWTj9T/J17eSnHEISf2paZM3dRT4+iYo1P2/vPVQzrOYE57qEbQ6rBlJTaf9xrPlnkmIa7nKP
jqDbfdegvstIuQlMaA6WluwA1EMxYnwm+1EZUefseHV43X71eDtknnebLXcbvjsoiANtN0jehOtw
+qR/tGqFBy4xrdF+J9vICmkHCRk5AGTUIUAqsDWbFiyprDeNUK5NtOlLfpuhDLPzCpzB2vMAhgal
m3LfXnUH9KXTS41nfbQ/2SceE5e8SolK00RuNaHhf29JN7dIxeitjU5dQEdIifWIoFTNC/55jq7Z
ipZlcU58jgk3WhZ9kzwRx1tl/fidlLDlpINaboPT4C3mpaKDsGWB2I08u3gmI9cWj59QZM4SCa+B
Kh5px6E/JuzR/5s5m+PtXO9VnTdidhqTIxwMn2bEjaXhx1lCzSYbpODBp6pcyzRGZyoiVPKP18ms
G9zAI+vUoerOMMFy1qup9dtk6ZQnA4Ig9Y8c9510p88WUQ3Ha12pHYxfJp2SvuHsu8sh7YsCUBLc
A8+Hzf+SFab13jeH3X+iw5ZiipoO/5KpWuYDu9qi+Da0lSv+YPiOBBSIfmElHVvV0CTBUqiKfWiS
NYpSkJSb6UdVDntGF0QXtNlHNezBEytzabkTzr8+957xvacBZKrQ2TwUscby//DITU8+ztIUIrnF
QfxfHZe3VFcdg9s2DIyCAhTXZHutCKgDlKgN0zucEtdlKyXTbFlkKJbaTfLcwoqFos09H8/u/yTF
61INkNJ+ZB7yl6eD/ZEJgIxu+GR7z6vBBuuckC5u0UXRpjZchDaGEArFU7olBQl/tBTb5lsg7k2O
gspmkXZ935OzO624uu3ID8/eFAzjajvS0AEvV0AMcwpU/+lPGGcUmgQRt5/mfjehn5DLi5YTAfd5
aKlIm+JE4aQC+YGI7BcI32GV8Tz/Z2KUul3Yxs1WrVfSDKzlh4l+P6+qgInUwdJgbqnOqFOaNZSC
O9cSpq+1Ke6bfhOHZr+GV4ww4T09AJW5X8PdqDDK0QDQwYn5+zT81hVzfAej+to4ncbOh9fspZnR
tyB8zHEaxwZZ5O9MNTr2VmYfxCAHKIOU6830UEKiFsclqwIhif+42RTsAfp9HBVm/u2MYkUwq4ZR
o73QsnuyHal3AGsrN9K6JcglgaWt2y/CpIdV4eMahDzhbtrM5w2DD2PzETvEB4w6509OtGAtBQ97
YYW5qmf6FuD2DIBTzrK1G949VS4HbQ3JnPWtStAHI03TrBFARuMXWRDlxzUuxXWjmrorf5OeC6Ch
w2rWsEvoqLdb/PUIyL1t3HRYwesqtRDQNpfAsiMwrHiKxTp718wVspQ4fxmr0HT5OyPJQiLTjOpb
gaAVD5lowyq8pqixEj9MftBQkVpDSJiUNQfVIbx80w8QSjrGtjtZ0Y6OwvnrXGqypKK0W5Iv+o5v
16iqf12zt2s2gdbqbvjz6A3wyL/ocKvVPDM9L4Wx7sJyKQqsMSAoZb7Yf44SSJwkRA65iymDZthg
hyiopqmjxFz0+FBNLpUI/r3hLUwlE5r1B+fDzqlSgWdyG7uWkGq97aZ+NGdI1qdXq1EKLMj15FKP
Y7uZaFC6dqNkGSHUXNMpmhG/sOycQo21s2ijK88mJwNUR64uRehumEN32XrJh002XMFYIZgpzBrz
xNu6a6VljOiyUrefTpQKaSU8MxyQM0aV2NmvjxlZUfLsotvYQejfHe826cjX/LwFRnMgfG68TxWn
KXNxeZMoiXo/NL1je3b8zuhZBAd9ZWUkUTNhX21qV8Ia/O5QtpUwLPfmQxKDhEgQGPQfwF3Nhm8m
AgghRLTHNl70DnWP/dsCSgw0UFD/EJ5tPKbqAONUfZI6QAT12lb8YrEsekw4y5LK+wnqpoUcRfHo
Iw3CvPLs8BGxGyN0ZeTruf4tvheQBteRdaJEk2WdeJUSU8ILLdnHG3SnDu6uW7ml52kjUpugo05i
LX2VVSJVZD0dbrNXlk7Fn18cZLlg6xsuqGRSD0mnEvS+bbAtR/izTnTKqyfTbj149pu3cLxxoikg
JcS/TJS6DrQ6mk+z/qJOAirjLyNZiBbVpSaqZNbS11oCvzAP+0UfLDBfuocnyw9yBdQKQDPUFFry
eLOnndKL5h1SoeMEGYjeMZ3hxklwMqQvwvUvhxzN2brphH9j6zQkfM2Z/IfCvPW63vhUZZ8VRXFc
r+DbvylHxL99dRlgmuARRtgPQpNvZP1Gebn79jAjgzwkp5aEQzpZCH8ORhV9hRSlGNxWtgO8El5y
k76x3diCOcnUglK3VQiBhiGtCtguu3lb27XUvw/TEK3wFjPFLQXiDvDKXmaxpdq5DzOSPuzRoQJI
pALxUm0pqtPDVxe4cEK3cN1gClXOW/xvZK1aCVkimeDZgezY+wVdPUy80ID0SQoc6dWNVVuG6lrV
oGDnPVt8kuDoK8v0MlDPj4tTEhhe0Mmp4D5O5XqoCmkHKozopSYXXOySmJmZV3CNWvlGj9Dzfegl
78OPQP/SKkhSJySkfmxnKIy50wnPl9muoBL+O0jbhYMj80XzwLLylac60i0At6fYYuJ4BAUW1SLk
epOhOFZFKtjNz2NTNvbQn89wY5y9nxcx7UQ3qDUyXi1V2euyVrbiACf5n15EcTUM4O1AoBbEWsog
7I9L3/yowUXFtV8YYzwfVRehkZaU23X8RxDia6jCUYQmKqQ29Sf1XuODIiHzQcQJ572BMIZSjXAW
uhGQDgj5+aC5dQ0BIl6i47dKi/zK0d2CRO0VvPuAvHcjDBbbPoOjLJL/7wjyC8UqZIQ1Ao5AQTER
y+mdBhv+jJLa0mquRqtr+QBBaPZNQogL/HLhEJ1Wzzii7U5543fPcnyZ1NbbwYgPVoroGhdyymZB
WFlpJOSc2dtF+7tsuyZc45jMqiKNueMwYQn3rJ2wuZoZChuJAxXKHTQhoo5LA5l883FHvTOKVaaq
tJvZM/53gwSVkEEpC7Tl+uEDa66DcEf7Ac22ofenKBBP9zvz00c0tVY7PwVtpIet4YK3gtzKEIpd
C1v8NleqxuaebPb+uP142OzgkDwUfhtzgjjmShymYAEh2WrqKGEJAv6z2zdaBX1YV5EJe2atuPHl
3/kyIH1yLBY4ZdHk1ZUTB+I3QXR3VkQv3DZDWETUJWyi3y7VWDCH+/8qVULizr5QiTw0PVYieW33
wRoFm4Ws7YQP0UQXE9r3Tew2/KssCtRQZBm2sNunF0WiiV3Wjte/Gi/NIuEhWWijPN/ZQc7JB8ir
xW58L0ldz/9dJkvfT4kcTjylclXDrzw53B1GWhxw2h5jF824Ctlm72Nn6dYthxCR/kbDnYyzVY3+
vCUIZyVKKBkivLLngpvX6/8mFyCeEAjuEj4PWmXt2l2xbQny1qZa3PDTjpzYyYBzUA6EhCxozn2t
dND84eJf1+x/+UAc7JAC+VBDx1M4uxYup1/+lLq+CvNuT83DvY1pdwNutawhBW9EOXyHAr+5wY6B
Z901fM8zNepnzP/1AaTkIIc1y8ZMg+Fbch4FQLfAoIVxL45jRDVXQGyHetIzTeqJWaa53UVLZsXH
5svsOzvOklGphOdMKhAJnabirw3NeTP0oa/SQjFLlGQLSRhsoHRS9Bstr65mWCi+IJPn7/D9Ojt1
WFzNPz7dkd9brWPlYhZ9F2613qU9pXC1m/Thlyvmkq682g296hf9VfUaRrl0UEBdfVUEF1TZvMoH
Z1TWn6znepp9/LmsxMhOBl8vXlg7GhGGUV4RAi9h8RAx/fkm6CeTGZnVbWGyYFKAgPxzdlcyuTow
JmldaS3p3sjo3uWFeVHliUBwN3tbxTa9VGoT2KX34aj7pG9nRQ8kW+tz29EjwUaUuKZFKru5qVX8
WfEYikgEmEWSnReSa4R81s2NE59BTCWF4OaLQvzjK9bs17HEBS3lOPXQnnAA/EpL3j45WT2/Uwwp
Dqe5Qgq1Vchty4pNOsIr4ssWOZKiTjiCc1KpkQMYwTRkvADfJfNyeGXAdBnUWbgXYPyYCyHxpEtU
LJ59moAsbJBeTv86wcUfOoonOTAk7vcsA4l6aOuGwPs5VTwLEk1yFqnGed+ucyMXSmUVCKPe58Xa
obrz1U2l0DQ7M3GWmPqOLNke4s88iFsOLdxkEVkIxjtPrFCVyPcymw0RYAy4bG783g9RRbGgdiMq
oWob5EceV5s51jU+foXD08n9ev4BQ4alrQ8Zo9UIfAv4JA4cJj3b8zC2YxA84PIDiNFjE4H7jd0S
fASekKGdfn2IcEF+goG/q/YD81p5gIjL2geSUzD8shx+ZnSYHyiuUcZxPZInZk5B02ScEHG3aSu5
BZdVovB16zhaU8xmTHTxYNZkbrqa585DCrQoTeTPDWMx8T53kB8fwoPOmJyicvp6QLHILqXndw9A
Aj1x61/ree+97kp7ZsVUFpCgM0eKG809LdUmdZSsPmJPtf2FFBrcWclY1N63PPKf72NFFhLKI/me
J0lRHlgE1CjceZemCBDTch0eob5a+es20sIrA5iChW7hgAZmn1xhK3SsiqWYoQX5wVYChZDHhnBP
Jh+4ej/rkQ3aUjk2sRgt8JQpSyT51S3tfufYVtWQM58Ojy/JqvWMTtRVQCoDoirlcxHGsfQxPLGN
vja+I9JwdBTcYgdrg5bHQlznKFltO21Jmx0Q1RiN0StGvsYeL+BtL/7TxFX4+83BAJMCU6Tlb3qU
qr8oEkR7S2UwA/hdm7DxCHJgmfje5Sj3ppKKtI4AJx6Gm2mszuCHIitRRteHHdduCyfjGs3nuphC
CxagRaJPJhTU6HrjRCUrpFUBwRCZQvoWjCAT58n3Udk/aZJBqfG6ahZ8iLZTjR6eqpG9nmikpAv8
qiduGl3v2lMcsisoqnJQuuFsFbygOhjCxH/3V5sTQPEUYeTnCcqwcpOPr9bRs/SkgDtQFOSXXmFK
Y4IjQWxla/BbxaYeSFt2QKHNHQGMeMJvYG56VTt7QeulNPQFKQv7uhdoyL7JJfy9RGCv1tqCspzO
i03NMaJ/9QP2yAtWfH+m854/vywvXjbDoQyR3ML77jCdnV4cxrWVSdm8/aFynEW6rJMDydgw927W
gtlegQrAmra3m0Qq9n/D2WezAjMafw6IcXl41SX2e0STfLyXs6cGmqTjcMPueYppu1KlUIspbg3y
l9CWtUrCki9LiuQgqUZMaJ5yHKbRUTeCQe1OMXcfdJE2Vp2nb3N4o19R+4j/lnh0mJiay9MrrZH/
+VXro85ErbnLRgnkot1vnmlJMGXuOBMjScLpiEm3dqxrB6PAUVw4DHgse6RpAQja2nyrR5+b1M3k
BQjjki83XdivyHXWI/38QH+4NasFYTkbB3qZZT6oE0XPQvBd502sWaB6K7AEDxxvqXjlhNBrvD7w
TUbdLSHNcZSU4zaPeKzHoJ9b3uZpbve+n24Bv2mGPxL3ep6uuE/fH8K6PpLU1ydAq1gJ0KnMiqwj
LVDHvFWJFcR8HjjsUXdQn03MVDKG5RVQyOvKSP459ZLkS1hz/mZvAJ5mj2J/qSQNNes2LE1i14UB
XONFuYcgd/h85aSULZ3T9/KyyyQwAZE+sHpLx9im2J1VvQt7PvFV6FAnC8a+6bLEmOelA+pBEdzO
8aBgbLz9h71kfvR5yPoyfIgGm0Y30P+uG/5VNNvnV3IYlpFCAnIQfKnrVPynBNI4jAEASuIMncK0
9mtkPyVgS7JfbeUCMpGR7LVBjf31eAAsfdTyplG1FYIJnAI2PWaU8HmTGxJHcEEnfb0QNGb88cW3
iZEPRRDH50gbT6boa2oRmK71dHF0mtUG7DHmyKY74mtkydi8oKV39vIzTo1jnaUAoyIXLiiB3Qa+
mVjaFuwYbQOTdt0qP3JbRoS+xoZZAvJUcr4MJOBzq0Y+uwHcVwjAYuh3+TuWsvA+152xoDgA5fp8
8/MHyH1L8uuVjVCDilgUAT9mx3iICi9mae1yuvo/TYY7AHpTK6XULdUQL+RSVAiOuEDuI5iVWCI2
EjtOMxiykjzy45KYNGYji4eag2iNj63PQ4AV5VT+LVVBbYfzscMStJeIZEaMRakMwHKjso2l4oRS
ljWMGe2fu7q88m2b6IUWU4byTxvZ7XPN9t8u1Kft4LvwruelC73zZRuD0bYD88ZOKi2uqt2V78PK
Va6nAJUxlLvGmwmadc/sKrvNhgVVPzhLPjr2Re79Kemt9t73kWOsegUut4KeAS0TzRIvNDNUDrzA
tpf0htGispl4tlGBfUG+8kQZA9c8fnSPoiLoPeb7c02HT8SOPKXIK/TyQ1uqxM/Z+55zzlMdwdSq
pN6W1UUovOmn3/GQo+QbbZ9DpbLgJWnH7bojCMpKMweGq9XuT8D6SLpnRYzXN2T+L8ECmWf3TWWr
pMp0KMv1UNOJ+KQR3x9dj3Wmo7RiDo1kBqS9IdYe6mZ6pPOBx6C34+9wbzjQ/gEOPbjFzzjdCZv8
ywo1oT8Djwpwfv4LiMRPxHHHAdxYKzDe2tcYhTKCGbeyMKJ5VudVg4ebIIEFUdSXYo/j3ttZVLjV
4k/94u6IsyTapE0XP+45cHzo/qVuUaIEC/Y/DzM5aA9rrGQ9CMPvvUC0cEPku707MTBWxn0wRuHt
CYQH9gmXnVFNSJXKnBj3bodI8GOoPwx9cDCbogPDypaqgcCuy2xpzl7ZxYAvXcrIfkqo2zyiBtLP
z8gWOCexWlKKckXL1fdKpARLrgopiG1wY9DNmyZpts6u/AKs+k4ap1/BC9iiVNRyJz3A2BEhZJNV
60nC590DzAa0owbqy45gwsXOWP2ikXSXx8Xp8Dl67hz8PLZS8VPo+y69FpVPSpOjtLUIUsQpm2B9
xKhWTqGwC0UO0syDeowV1TdL/iT4mnsGYr+0/Yb96GfKxE1DKrYxbxyYyCMdu/UvUGmduLbEZ0eK
ieFdsuSFgLeny/vAtfrkQPOOcEudJajwqxCr1s0KE4sst3NImWy2EyGCutj9z1LtfbM5wxcwFa2J
CjEihpnki+XKapoqqvnXn/1XAIfFMn7P+IGRa9VUn4BYSAMz6pMBofP+S9I8SkPYcAgShw0Mj3Fr
qh0FWu29qjxK3ziv3xdOunJyGstUQIXVINJSRaQIdaKLd7JSh6u0Yt3UFwWI8he6dGlJbRW0bXNC
0z6qU0fE0l500AJEkeFKikKrpBFvkswwyK0pbTGm5qienO8DlueWqGLX8l7Rdo5yZc+/JwQ8zCBK
xA8sM4d4yrsDU6Sizke4rcyxFL7orKBrpYJM6lvGUFx6jXkXaRmZsXW9Wv6s0ZHYtJfRpt1mGM+z
WbUg7EAaWf3NsGQ1+QzZ6k8awyvJH45QxfaZCVEdCoIckKsAUymh8MwN8Ye/OYBiqWCAc+9KBjiN
AWy7gvx9fa1we5vsjmE112Bz4r6Uu79RUXe9Mt5Cz1AJIbzjcVOO+EzkXt5sGYUgZTj7t0LdagVT
f7NfdoOtK1MrAYW8qEUhTMCkETZGxVMOBbJStCsv/ubJnt6d6s/2MCWxvUAKoQ9LoIKHDhjaDg0N
25gCVpEI8/BcNnMhVp1VThvdhoymaen/49W9bYT5+RrCe7PPmQ82ipox95DjRZPAR0qwcqyPwbsw
GPrCTyFrF7F2A2zB/QYybmnlPRPDQIpo8kLDw+X1ACeoIetpxiBoRU+LfxRR+fjs8r2PdchiIkL0
6CDJwJAbFHAp120Hewuh4njvQxWaS05MI0PKZuie2EVsr+omj8d/fP5Zg3mN0p7EcJEls3+zfRJG
f7Ky/PsH/UlHZiKjux9xMeodVqTsrXzJDynWwUh6gAgjNloLESzAIby7WkrhCbhWJqGnMU/irN0y
5OaxoLmjSfdVW0MrDnJjICpykqgHiJES1mTn55Wu0eht9Ple7XVQKzIaDPsHc1vUi34WYBR8cSaM
BdnLv9ye40n8lOgxnOtHcs19RNbasqiAOQRGfgRyQ7S4Q2Kt/ES3eX03bZvnd6fCjO3y7hYp0EWW
CJIFNlL3V3ov2bdQXBHBBc2fl1955hEq2tYzAG4cusyOg9F7OhSIEQ4w2GrNnb8Cu2VnVI+1CLSF
CR7HleqMp3fTC6frV5X+YRi9NLXUtbk1hqV2ml4Ko+58CX3lP1ck+7XZrDCLaoHXDCOKZIh3NvNe
mnYzblcvrGEMX5ouemdFFDDfefbHLEZIk6GrvQpgbpPee+K5xE2tfTKI0SW9cKKSu30SXwIAz4GH
pDgDM+4lIvv7RAQWsKGLacdK3SFCrwBsS30mr8K7ABkyT29xY0ISo4EfpdID42n+GhC7krq3Drnk
CqhASNHn1gfg02cA+57sYv14M/Cl56TveijtH5SkS0uTmqOXHLHNtTwBPkEasazRoNDM4Dj6A3qO
uYehVdHujYLSZYjavu0LKF0XCrqHaJTkHqxZAr8u5NU1V8EuRZtwRUwzs5hKWe9O6KuuhgAVlsyZ
XVENmzYpQyn1xvqZaAjjvG3B1nGpgrnne25rni9XHWtghXlfWfZ5a6UBU+V09mv968108Nh31j9i
GcnZabeYFZFTllqYyG6iyzowG6ExeBaukpyMGgXP+JEDa9n430sb7oOaJONqfKsYSvoo+lNvnzs0
HYUDrKssDAk3v9p20+eTGxmxjKmfIaKSL+22cGK7qsyQWWYRVyrUtNcRDcrJx1/Y6G6JrQ37DEN2
9tI0WDULueqMJ4qqfaSZ9d9Ro1HSLXwPS4ou1yRSu3VUP4mIUGloOiZMSJsZRvuOcs69k5bdSB68
T0KQqHmxWyk21RDVdpZmIXRC9dv87O2+R2hdC0TgIDkOtm/hGWYNDk66BiuuKC8d22A/FzlFBZ8P
ooxUU+GyEyppcWHfOqrcHTwcfSvlUmeI9vl9PCzVCBcAJv9ii61+4tkFGE0iOYoS3MTv2JuWbROW
F3xOSwtkGEGBAXihLlEJ4kBhaWSq5g36uD91Xd/xVTOkiYF3L04VlteUw1P3WZVc4gWmXmEM3ABv
jK30W5vVtUKeq0Uk2wz5Z6wBfF6MTyJ9I35caq/44tmaDPDpdY8hvelaJonhazBCu6TcBP+d3HuJ
vya1fc0BFrn5zYseCnorXK26ILYjWhyyuqOzHkZK4/tStmDZANuBIBwlvBZRTGnQ44xp33Qbb+Kx
t3B3FGHU/gDHkUJRYK551TT9NVvk5iPXHUJqnkVaDg2BLcPIrq7Gr5PDMp4rTsOGQ7MukirNqxJT
ZppNoxnlaa20b0c5IqS3iOYXUN3oxBfJI/ps61RA7PiBkkSWEc4It9xEzzXaAfJSPA0vqf6UvXb9
U+vZe4+5IytZH/spvk/oYRotQ8FdLttMmHYrpPz4Ak75NSv/oeQwvL7UKwNxp3fLoiqWoM0MVNN6
NbI1nQ4CCuIGV0LwCjDcNrN+dGW18DZFbc2S4BfaH4Y4Q1BNyyMQYj66ry48xjIIm2PO2FfHkBbO
UXc9txV0Yr+Z1zLIHMBfHGZZeutwRjt8nXW7W1qOtqyi/8oCvDI030+RdXtQorPzGppr8T+Rlx3K
9CJkJZRf7FrPQv3vZF2UPgr8RblrU1aD66ccRLnqxRsHmYx2kP2XusJWmwF164pl8mQOho4uwkw+
fz4Q6tX00d4m4d+/iHsorQPpvGrg+jrcWK4JPijVYYXhOp1MCQHYJ9FINbqsEanhpQy6VdgoxIpE
TcFa+ODMcKJjOlsp7ZniGdOZwNScKR3c8LCs44Mus6RHWUJv3BD7Wi/AErQg22M5ziLVYbR8m+Or
pBOLw16AKUoGi4BVSpvspMLM1+8XFHte9jVX8ZqEMxKL6GiI6vzziCVZdrImXTQ6LltdBUarUVkn
s8IujL4rBF3o8LZmqnmtS/Aop1XHfdha/JHBXlf3WH1ADHFDmNWndAMKzWkje8ouWx8FG7FNz0xX
EiX7daOyjI8KrMYEV5cdmZbhmhjMnAB67aPvXl8i/V+gxUsjAvihP9ig5OcuQRk/N6DzKdrlLZ+1
KMJSQFeP/ym4kDhz3hrXk14nYG/G0Tlt3inw7DRMp3aGl+mjxalhZgAnDhHbg4mlKy9WjEl+gM2+
hUPpz8l+8xSRJKKOanlQ8Tr5zn7vbU1jGTG+8R1C9KBARMeYg3aZU58GXSBnH4M08I+40uEcf4Nm
aQ1+k+ZJhDahlBEXbH4obpXXQYCvszMuT5ObITI5Fq+MfE2k2WX73qk/VgHsErHlXMHNKyJp4DHf
lcQkTJL8mUJ5biSGYi2ZoH62uVj2Wtkl3h7fW+xIH67gKjAPKyap+fdiKxIVa7CVY6CPfM4DkW3Q
ak6EkFo/qP+vPom4wh8C1CFBtqhd34eoXqYs3+dkj+0VrFxGGv1GeBQUtyBqkfgw8h1adOyzBx/K
a0lo+pgjWhBJGICs2tkmquE8tZon16wJ5kXBSVKw33CcvP1DuEObFZVjjdyDnGdIi42mWiz4Sref
w9yspmJlaNqk5B3Qkv5FNeDEueaag+fU4KQPB+bLdV4OOIpf95zUefIyUSXIKhvDnsNI87Y1Eym7
FdWzTY58LUxFZCiJuQUevZEgI79oS4qFBNU+d/5xnaTRZgLnD5bgJDEzKewDfgyDdzoXEtVho95U
R1TLx/oZw+fG0L8m5AzvijIVoWpfCubN3xTgFjWn15aa8z0L2c7H87RT9gi3Z2orrp4ACH4575MN
+3X3KTi8HS5Rd9jtBs78EdOfVit8f5s/vWYNHwqNPcK6vcsbG/IpYtmAKoo/suH3JUuNQeABrE8Z
UqzTM5I1xG0hpnnJieCpCoQ1PttNCckRDDNEdhhOqyd92ilS4PMVOry3AD4ZoTKdAxmROoK+VRFy
LaSB0eTyYLPK+Du39+8llAV8jt82/gOiW6gmg/Naau9ZJdrOGBWB/g3AUDC7pEWcRVMabLIPK8T9
hefNKyQOjtp7mkd33x8jXLpDAanEWmgutszTG0d0V3F8LP8ke+GjYbeY9QGI4ShTroJ2EAtRIt/d
deYoVCdSDsLcSsx4FcZGr58+x2fakeyEj5UkN2UhygyNp3L326T0f285wngpNrmctw+iDrRqVrvh
qpo5PuulTtx1o7WGPbnyucRTEA+2+AnqdPNXrpIfEAJX6XouqI3w0vgwazQcI1SVQi8/r3VU1Ob0
eKv1zaOT5FpaqA4a/gUrw8lei2zEvyq4t40f+IlrkcKPohTVKfYPOvEJTKf6IoAZkJ5uMUfASZsU
hMnDn70/m8B0vbzcyhYJQNewhPd4MVBJCFefm5BqMRMaNXNOemCnAYMXarAZupwQnLEeqDSCbGbN
XN7zmeanZdJwvfnWrdgBm3Aw3t6gXduLgGgMV5hiDiMVdBIbSartCtMrCW0h+PIe17aR5r67Zdte
In/bO0a3t2kXVu/2Ns6XA+B/UIgyzb55+zJCH+KRAYXx7JUJ2riy5DSBX1gdyuYimJe/nJXr9ZDk
D2zj/9djhTkHF+BcfOcgTMxep+54JXeQb2I3ufznRxLt1a5Uf8kOysjzpKl3GgKWZeQSWAbnHiM+
bD/LhEh0BsJVLWquOk0L1/2muaP0sspGto+EJJ01aPKVt7vY/S6kRMyDkbmUTGY7cHSfE58GpTwy
Ju+IA9PNLvx9foPqSw6hSSdWyQNbEnuZJbCll9bKoff9EAoTbOhgn/jmXWGsQxYewzFmuFaYW51z
2idGfiztrE6BjkVD6urlfpl4Rfg2jdK+uaAICYKNtGvb54g7J7sq1wllyuIje4OeDZ1ATXB6IBkh
XxGIVgpNShW7nsJPefZ2H9plOdN4hwpqVfnR2rR3T/6sSu+23sr+PJhOHjbXlv6OV1ZnCzzH0KCN
hJgglt5Ap4/xOBuvDQLvD2vum/lqMQP6ONPJeDWOdFERtL7bZ13OcgEcJioRkk0PT84He6fG/RUb
wGkRWG5/I7eMfM8pcRjjGjvIodGZgi7h2Adf3ZuXsXSEPxjO1QycIaKA6+DnUg5CtRNvKeS8X6WN
sIOPxgDLxAN1DKBR65H/2Nasfzx+a6eBb3ylbz/0qK+H/3sQ/V99pu7ktyb0M4SEKR11BmJ7NCoz
yclJ0UzeVOYZi4ot242vXff9bOQfUJHHckOvjAc7QMrnjIc7ek7f2aCctXyQ9TbZFPAgKg+3iW/H
t27n2s+tPw6Yb2iSZMLabRTQgBpS0trGQYQSBeWvSGQZOUqLDvRY0lORSeRcOsiq08dDAvO8zxfk
+cK8c7+nq8GjMP4CoTgHKl5lQuA/FocJmtktw43jC+DsmEDpI+SA+O2IEf91b9PDPR7pbu2LvZSu
CSdGZsIChZTtpYD7Sif5Csfh0NcU9wEbdT65Cvai7vWH8g6zs8ZAJw5c6eR/ZjEO5lvfM3feRtqp
mCJdJYW/KgX/BeRCdoCNGCedCg3+gkTxN/c+6iO34yGQJJp/khxcyy/ob5TXj2C57cLUkrUtH97q
KUWPL4iXdxuIydtFJPf7z69SJQSYfB0ICuQksHy1EekS0IiJ1LQsAzC9CGnePuiINYCBUu6Tj1YI
mg4Ow5POWwQUwRmePZWVMS5k5+Y2ES2AmFrDeriO1Y8fpmD4IfakvcuFUBeUbdYVh4s6DIuOOq1l
b1Yiz0Kq7+ZmLSKC+t0v6Y436Vl5vDYvdOnickrDutygRs2eDjamW61/kfKaLAyPQds16pxtBLXY
WqxYrs/EMZoMwsAd5vxj1i2mi87U6ovyQIuyDMocpjFs7jl859VhtbsIXSewVrWWE7FXsLKC5Lun
rANxgeVLAVpwzJxCUEENrkWMXcKJovxSZicdZFByn2EH2PoM76axtSS8Ehs3cdLs9ldC/WYFlC3j
gsQhCroK1BS+oqahj0aGPKdY3Vj0qdobCda/n+zU8dHnpKToUu1G2IwjvyvJfk+fL/enm08GJsh1
ZtMbZNauqWN9hFtfTvI3i4pb7k8t+q8ZOvRRyZPYNJHHDc8JgOLczSDsG1fKHKmg1m9RhlIbUzvP
uyj9U1Kj+810Pj8PdU7MMA2fTLrwJlE5NkcyJLcVaJGn79Q//rbNYUYB77yqzRvmf9ZH0+2iIc/G
ga/7Pt8B5qu+N1tA1A7gwKWrrX5aMwl10aWj1scZgNC02fndDWA6FJ7lz86F38Wc49pgT+IhnQJ7
8IJYUHLJ5Lfq8RFj6U5M1ltbUNcxCBik1b5CCeIA7k75kGy9Gv9N1gA596e2hRj6MrAVrXHLtCqA
6PZ6b4pqs56ere47NMs+SXRnQOrjAdKlFIqp/81O6t1Goseh2J168qVSKsvUpeA5zF6ugP962cI+
1dpRp7hVkDkugls8o8h9wUVbH8J2CXtiKJeKtpKAnukXNSpH1QX6tGSFgR6oCgi9gWppoqQq2NF5
3jyFyjuqZNqYoyLsLn/OyOZILReXKJgRZMgV15Z08pXQcaJ4ka2PhDD4q33mxdxWMSoH3vZ3HWOe
1qrNPh4x1l7T0GFEqg0m+68+zw/0zn8qzXYDSidhTkqxwSAIGqKyWZR0jDH1leIoAjVkV39tQ8Od
Wajq4v7Lr3u7GlYK7RvoDyaKzH6EzPf9EJG8tTguCCkOwK/GCsNKAQWdWNd/AHybo5LDetTpYHto
dYBSTvspF6xCN/63HhO1GwUtB7lAf994ndMHm4IppLf75VOksdUtyuMfo0fmRSFKHMW0raop9WBg
ndh5DCDyqRUXkHAfTAwquE85BYM24hPmL020ypluOFCJ8M/wk2lcNIJSVTXa0LY6G5MktFivupu3
tcspsBY6KdKH2MGMUL/4bCvJiw1rHvdDBVDkgnEglPOy137B7yOhF1iHEL2Zo6HkBInq+PILSkwc
zhpRKY91Ww9jY3ped9491bFZ7uZYa4sb0hcWMkk+6WhDa7pd/TSCVjyZ/JlQEy0OAi8gWrRPPxcy
LErU+wwzOdgG7tRpKpdoNVq+AWfwheBXA0itcjecSY7VeVHNcTgy+MYXVpExOsNF7mALrA0626bO
3/C/20+3nnm6pIsg9DdW6Cm5uLAI9BvckGOpjXkJaDjvIlr8R1J2wo/xgnERPzdLVEpxyp+oTNbY
Q8NYpipn4crktzUtA3yOqKRe9CO87S1TqwcB4YHhHMuu1wCXA07gDSnb9W9yuFlybsQYz/AJdahL
cq/Km2SjexbNKfhpZ5NCMWwWx2p8WJV1Mr9szcuV4nYr3L4Oc/+O9nj8T3HM+GCERxemVD/nK/UK
huulFVADuY/feR3wqURDGpu1zLfrPtaK7OMk0KJ7ogiLmZVXBFu6uaIM/NLFaSj8YTIbkwbxqoZj
ar4fhD+RasqZAws/7csJ+U2uetrCR1J0tMiGwknPPqy+2eS2vvEjeKj4ke5JVmt0WbOmORCAJvY4
6GLKDNE2we30A+qTNWcdZfIDy8ssoOCu35qo7zjsN2/ksZAsYWC38+hdzAbeP2m1mX3jeCStX8q+
e+eRwUo0YzkgQi6o/5CFBcD1NkmFIzoedwaxy+UX23d+HG0Urw7pDr9IgVmK0/DOKr5Io2oZrXeF
ytf+OwhDGLPSJEM3CLI6heHjnFjf91Jko8KLiB8F9zzyL2FlW0OtlxpofJOQt1INMXt5caJHxjAz
VVFzgE1R+GqIKibaSIjaKE5seeDdvFsHN2D2ehrk6sh4IHfz0PH3cRtyYaQBjftxA2WwxiQDWtuy
Gc0ThBlGFEjACjBf6IlX1ex0WDUhMuIySqeP5jciWwtIObyw76ICL136S9kFpws6tJcio8aW7S7V
WhIa+XYOO/RU5JAts553x4IX0ZnWwC23Ts13cysHC11XLVz/NgKPgE9sDOzm8TNr8fGvlecyZgeI
4DrD8lDyIC+n+/FOHc3fvbOp6D5YjVDZZKsBcbcuxhtVg6KpRgXMhBZJpdIKoft0K8drDmOB/g4Q
Mltq3wT0hLK6tKQ+BjLbA+DevJCphXBCqYfG5XVOtbkIoKytR/pEtjeVa+RrGLXzUSavh0lobzEZ
cvI+20mreMDJLsCk6PqhDbfe1GYxV9FyLg2hA1bMjxWn9H4iYOwqaVyQQPVaWOq9YT1MrnZnTz64
w5K7/H9OVHDNhC9k2WgJA2OotbvKxJclYCF3luGhyuHV52GVWi34gkvUYiUsMkCGsQfEz1VoZkzK
idJd5aCAznl+TNjdEo925oIuU+U1XOs73frRoPMLmokRdD4/LvvfUU6jcZgsSe5fTs091KNtKeno
KH01LuHcTheX37LB+2y0t6tk6IRych8WdCiU/hjvAHSH6hEFL52oOF/qZE3zJ2iltn2Bs2ywiU6V
niKsZNOTwEv8C0ItJANumP10epVEc6LvJPV1sEUcHwQAfGScHiYHXOnbPrV+O7NrATjFAavavcNW
PHP0DOaDlIzM/6fbt2ofPs6rfD4zmupV0W/zIsWc9MX+IN/Xyb5K2iirS2JTIC5HbqZ9n9aj83hV
omeQXRb++hHeEs+jNdQcWWcvo6ao7S0Th6ygfHwDXAyUTUjy/ct9ow8uPxGvGe82AKWX3/ySSBFx
0dMJ8V0iZqO1HEezYyXpq/bQnpGeN+lY6pnmb2MIH/hVyCNoA2VPs5sg5kYxCl2CDPWtut2Ab4qO
OzRfpsfmEjKARX/TJz53ojV+fhwCE3mnMUQOeSrR/lbGS9Xc+lH+IYpxxg7ypw6wQz21n1u+umNk
/vyWNYkncEQmjA+i1MfwZ8/VYl/nU6oWrOv+d8j/WlqU67zcqy++xGc384YNfWcBTjxciB2V4qjR
codzHHQf9Z0hLkxzyJLw8J4VPYFkqtZKO7NifWVOoEB/cbjdCeqZeErwLJ6UhqbJxTpwAl5rY338
a2r8Q6MC/huB5ZGIfkJpc32J2MDRzoLuFMdYgvh6LEOIH1yJATF12AzVo7Ds+Q+/cUkutoGdQYbh
EjUXzBit1vxw/Dw4SjV5uXc1idYUbQvyNhNw9tk15y6to/z+6zPJiCRK76KB3P10QXOGyoXhBctD
Y+MBx9gf/ay18MhDpULn7J+ABK4aH38/9c9E0OVz7gO/QnzAa9w3f7RmyZc3bKmUqKve3us3tdz3
RYfjEao1F2QwD7tbGQc2raFtOqyJCgeuKdwD1d2Dn0iqprk77NOwYNUrBIxzVirbQgPXYPdOC3hy
JNT/tG/E1L9VphNMu+sC5232Jp57VjgrMRsePobniF5jRjH8KbT7E/wRlSXZYPCja0SHBvj91+vl
u01IXGxY238NZ1VTC1KhQkVET9JG1/uKejdL4oohQETKBsi/0iX5PgWK2wsvEKgXcMvikJyNfMDu
89rDZpNKAs+DS/i2VwtCLhjtIh0hF3fL0jxI8EeUlv3Nk7KrgnsdpDpmrVgrQdAYi4VC5PeoHArM
zx914DP47twlqQx1nXAVnuxUzQX1IjapMGX36hzk7HN5/Gs0iuVFYjFFJ1cmKOLheTNP060NHiQH
fdMFWF4OkC9n2fK9XvQZMpUD+GKJ3m9GZFAJzLxTVN0LMib/I43y41psLbdH8z+4NLfF+Z1THamo
0G5XcB+WdHb1YKaAlmMdWxcB34mhDBQxlNGVd+WKdQzPxb/Ho4xo8sIKvcknpsCbTml6ali56MJz
zcHAdDcPMeWFOLEaIAJOx8Z5gPJttOP5b+q9smwa0n6UcIRJ5CnTmQKU5FkjXsEKXQphFtDa9xYz
elNJ+Hdq5kcAr02f9rPSWpm+2MrxPn7ouRm+PZ5nLu5iMN8O/ndKDMVvvEsrvt1AyhxFYHEORE/4
R+RkDidECYw+HEOp0f8FtRY8jMJjr14J35+oj2xGpJW20DzGbnBUlBGorMWMwaqXmybdXdFOPJK2
OCvF9AeTO+XBsD6DnhueJQNT6f1yS1OCRpte2Q+fHiUkP8VyYPAyUrIretwmjb4KR/KHYi7lBH7l
QWvVEbFf6Vvsq6dGhFvEvwnU+v9BLk/ynjM90EUmLyyKkmSd4RRGycjbkgy5IjBSBbfMYSNtwSUL
9p5wqco1CGION7RA8dOTkrPMs3JhA9QITyBTSt8ZLXNFLPdjxdrjNPeuhO/GVAnfHlnEhRfRPu39
3RVMiFi3fam+XVV5bUkoRZMq9rZ9s9JG+tRarCH2kHRWYSyKzHqTxS/ejn3PK4sGLF+eIal3aMdT
2qZXTcu+99Ak/sdocPvYfhf1O05MtJpqMqm+GGAMkQAcGmjCahihkdV/yr9XeFWKT+eUkl320lm1
omMl2N26vZyxgjftyG71wmORy4/8vtxiWPW3pHAhr1Rsv242C3gfq3w4aqbNJNaMftQqEWKUFLLu
kwhOS++GFIadlrWMg6SrEcO5hutZP5ylzBiK0Az3qCT7P4j/W9KwMvijXomSiq2NSEgC01FS9FZt
QaflLZjwXruBrWD6HBSPxyE2ZMInCLHHb8FbcfhQEbTn68sHpR9vcQg1K5UWFoHHzlxceid6h9Bz
Us0CsmUWS52LxoRs7i4NM5OaPSS+tstR9zEzDqWkHTgQjNqa1w6YN/0J47DTt47Z2UaXd1NJZ5Pu
K9SEUGWm6Gt+LuaHxKBE5FqQ89h6N2OCFp/q8RL00pqTNm/3BsNVf89SvmhiEKtmTaF46cxKnWSn
V4ss8jSjF3weqMoLszuASCAFfAx4hNXKssQPtMD42uvSgy6T/esADXwTyvcHmsVn4TGcFISuR2f/
3rrD+2fzWmOC2I7RXwN8Cpi1MNPGcEKetQo6JK72tdBYBxmo5Rp9SQYX8WFjFnA5WJLom9R9VbTF
NgYmHnwvXRNXb9W/NDbcdcY2/DCY7Q6/rnQgDZBwJOHVWJDaajnev3AGnR8obtoGGSB0iIikgdDR
hNMtHzl7eTslVeJuV29Yp42M4wCM6EKCZT2KwDI3OJHHNRomPyPdSQYJUNOjRqL+3TG4xTQjksTX
KFMyACBguMUPjZfIyEG04LTnTascUo2HWJIRtiIL+tGOhTrjIlFsqSKr2cPyL7Fkttaluu+cUb0V
VVjx2YJUCPGIOPLoPU+Gu51/8cpAxNdA7ScnKggcAw/RyKrkTzhaDF8HJ+tdNAgtXdrMoz4sFlZI
HuVkBVKvUP2NWx/wb/NPmFA919VGZQzyLzsE3zvWdaC4qrwiLAzkBTnob0vn6aysumH8xNQptiuk
axzfwCq4N1vD25i2PjOMS8iKeyVCuVGAyG7qgUcsP0UGWWSa8NLQa6S+x6bEBEcFUl6ek78HP04O
eGy0KdYTd17Dc6wl6Ht4a3ATqbtwswc8d6zl4sLvQSWA4hTputTxFA9chkG5tb/QLvSh3hFnw85s
X2F+r/MtCAr3DCOYVYzO3PKV3xNi9p1cHzcCRMmPyvDmGjBobvqka0yMeJpEmC2ndYsUHYVplkaL
Uuql8MffiGPI8dO24zzTc6YJbgB2qyxpXoikNrkGLIk/86qEA1h3LFPAXLQjc5cqZsbNwWClMoeL
/ICG2vbhMHMWBQ6GTGIu0U2goOPwMbN6dW4qpaarniCL/T3IjQfNkwS0fQmdg2jLpnCnHnu0KPSr
o9FV6hSJPJAgXDtfWVKRm7/3+p6iTaPvPLDFzNlBhaSfZmHrbyM5oqchbLKPGj8sIUL0zL6LPCvD
fILd9Aw7AtueBhxA31wUsYJKVBWs67PTNA8NPM4pPecBlNYlwqRn5lqizQWvBhA4iHZqzd/nbNlm
IwzPmBh86GwSrBHLHagj1/nn5Ue0zwDsdVNCS4wTjZ9GSDsS8V/NA9EQ3JwjH9W71bqvcjS3eCnv
qM0lK4CL1YOH7PJZWLT2USxuwdSWtUquAFKoYxEfV1lZaQVqEM/XnqS+MWNhaNYcUyla2kiSUk/B
Pwg54AZ6fBGp6vUtElYFP1FdbmYk3LS24gm8cLCHW7pVZQmYpT11MBnTNG5D5Wjkgv4o5+r9Jpe/
h8HGo3TzvRoapUVxVM7GFNaSNuE5D1syYPX53qrTJbcmJ93wRtIh2S0mJYOiuXPB3bHg9elK0ecg
CszNXuVwvrDXVBzcBc98FkADJhvPmBDojW5/HYLqamHtR4Fwm3mwftpq5bMBo/t3zqY3Uuijl72d
JQgTr25F+dJMlgBYjWpFE/Uglbnp13Tw9kWX0v/+sTTskXpwpkadd7g1wYIyEEV76olJ5552hFlZ
0mlWOxtJZQRZ/x0QJ6PUuh/NCr1yayFahdb4mBC9SLArf5Eo2so3d/Pb9dNfLWB5gvOzEiEATs6p
2/qOfAu2gyhMZTdSCW68RYJV1MNCGnK6MiB55qMOCNazuQulIPS+sMco1TH3AsLeH6gBitDjsTid
svlko8nuCNsRQPZPqTIXDmpPnSMlIxDRvVuDrkcwZ15WJ/0Vme4f3ZCiDb47/PB94/T92e+4/Gbl
p4KpB4S0ZFNExOjI7ZdfO8H6z0FigL//ZkKBikF4ehHzzQRE3d4fSr4f2vwrxBsphxLgs6NnTKX3
91SrDhMoag3mQYSK7wRyZ/iRGpL7JoDnC15D1QE2rRWMc0D+SEhz7lh+A8YwkBw/757LKvyx2KNR
kwlouguKarbWoGbMgmZ/X0KU9fwaGIhTeDzalOqA1b2Tm0jEZTZBJLRvpP5H0uKAHgty71AaS+m4
6xDvi3i3+5FJi14QAHvwuII2Lg9iAmmn+tP2OyTHwFWC/5Ya8sXuBnVMx1bwRbz/rLj6bPLczOpu
fjSsd/TVqriBObI9/aNJLc80PUD1gviS7RUVPtwD0z7AMOK0sQ/TgrCa8w2giKrdWl2Rei1golUU
mlGnbHaVQfetBOXTjCwwSBU06cQz9Q50LgEcYdcjT9x4lWw25Q/UIe9OPyKn5HRpSCrfJlbBlnxC
3QXre29dfG23JSVBJqfKZUkf3Vl7v9iDmc26leCCny4yqRn3BYrD81onE7rBmiw/2CRhV1caU2iL
+eSNIHXZgEyRFZ1Hk8QaJ47aDys3RFYbLl+eiCHFuvxO/E7TuDZLr8MJO4ZSNzHxnh/pHm9DeNFY
C8ky+5/l/LcevZm5s1dVpQ20pFpLm4Pa+fCSlo4hs1S2c95UFjs1TuvOml38ql08y9etpCPBrGSO
ZFiFSJ3YMEb7pqirV95fpBLndnykOSK3h7RjsrITxSQks9Pbrcagx5N/tcVsqwR04LnR1VT+uNMd
8UdR88iGhswbDMLSS8c7AqUHgPpPqiEP/6Bj+OrsNadD4x9DkLJKFMBMm1n7IE2b4BoaUTE9KWzU
bP9phaMXGsf8LhO0ugD8twxldLkZnkhLLkS4awza6ppCnN5vxBBAvIJdhoRC4bcyFkm7P9nhyXZl
itxBLJBdaSP7+njrQND8kUiarlAdWxxmCGoUqVg/AyZpRVZj6nqLwdW6ohcJlOlD9ZKASDgkCLui
OFYFjyfai6MHhYpYu4xVC0bjlRYzvWEGumryeDrhDkZulrYWrP+JncOky1T/EpQ9tvAcYX/g3YfX
JF/pxmAENHRSP3KgNvtmdu5LFsylA9CbzqcXFG6bMfubKkWLkb/SCaXE0AlLqldM0oXNTTTIMMUk
zB07oZG+HaieIZ0j8UCQrK4pt+q5aeUwZJvu5Ri66Xc3ddSAVEmT8A/bnLWtVbuTMJbAHcjLPWNf
3k3MSh59m42ZO3P1E00775fpKigqBYWBN2fwE4Jd8z49h5qA2bIgPHZIy4uiamCtTMEW990F3Z6V
MuDOsaQisk5CmiXD3bm7by0TLvMhjG51016mMfuSjpUGISen4NQgMWYhnsid+RapxiOTBEoUgn30
D3Gy4etp+qvuxK0M5LrunsKTsZ9xqv4rhCq5L2wVU3l7eKebIuPx0YiyXxc+rj5p7jqwf3Nt8qOO
7oq+wKj2H3yh5VV+5/lqHcFjlCX5oGpBPCxpILThk9v4OYa4gOKolC/AuG7R6bs6qp5Q/adwObIT
0u5Y/o4wEqX/J1VQNpGz1PH8iSUuGrCw1KaNRuqBYmvNklDG5J437ezQJMYRBWPnbJf+yh8TWAVI
66UHdab8atGX1/R0kRklB4+Laia1gQuz9GrBr/Wq+ghjlfLxrzzYNMhl8dwUxJJ/JD0XsXXwUgje
RPROt61aPsPTOmGqFmAeR37U7WqSGWpzxXeHVBpQIEaOntqJ7cOyRpn3SDszWNSiOM1Qafh0v5jx
s99i5MO1TWnIadxE/AZOlht7LW6oBE2TYX+MeKaFwXjAOSfs46RSy1RRWG+QQ03QzyjsUGiFf+v2
70zGrerrj7DprisJ/efD4ZR5InS3Qu/1ZC00VRtTfAyMfiNhAiXlfAptUXmoESBBZw1it7qHhtcg
Co7g9a8nWV4l6xgxOAnQMX3BLQrxug6JnyHxDAEKXHTq/NPmT3HHECui48UPRSbzoSnxpKjjlnta
oAmqdKiBZOUQQ01gklbPzE7K2OVzpXz8SDpZDHGp4XICnQOnMq026PWc0CeGVNvl1tLdByLopxZv
5ISUYJP73CmAZgjmkewcjRdhrNsfGXRz3WCgr5XqbYSIGLYFOIQRFwtUnll4qfKjVYSsYUh204/P
ksZS9jgmwZ5nG90S+ut4Tlxu4LhQJ60rUJ+L8EyvOSTJ5Y7PbDnZRvEBlSqLLGiNfrCbyW8WJu/i
9eBZFTZ1/H+LH37A1MulEwnZPhZRj24GJ0KvLU58oFKWJ4K1bs0ihtiU/of4nLuN5RpoDYN0WOJF
swDqvUX9kpXY5/UxIoOYadfp0EDJW/6L9BaFDmcaDWS4jxkaE122WqkM5Ji3iFV02kcYKuu92A9j
ispOfGhIevw4QWlabgCruF4xFQmSFet6amgCBXFWiDrvkAsa0wJ12hXz4daX8r7IKIe+FVTHpHOO
uTZ4JmNyivqbNy1uaJNf88RkeN4mHeDobFnrgy5+gG1uYjthLZZy/iHj+Mpj5RNfc0ZsUm/jHYyP
A4i9nNNcv0sWFVJqkTOqlTsZWm/kOMA9bTzQJAZ7VwOnuMTlHV/GtDubyPTFz/8iwkP+f4//QyXR
bDX1A3qGrTiSI/x2zdCnRXNpfEPdCE+gQrLh76Fp+vP7VQVccuo02ajIz/TKx5a+q1EJrz2CSmcC
U4ISgS/MH4iIdus9wADO2FpTiv3HZ2xr9I8B0z2t3NzKFJuddoI/9U3OYnFIqM1YxNCY89VkM3sm
mt78kPaOFPj0V2bNE8AB7GxO8gW4uCZ70hHWiVByb/AL2vSYAWVp9T9tf5tdX/ult25kzuWV2DAi
wu6wkJVxBdQtX/BfsyN3syxjwP0SeNEYboX/woVyTrFaC6s4jmCeh49CkOjMRLTZ9kNCs5m7/F6s
txv6SwefH33wHUAIm1IU7RL69H7s7McCTWt3qW5wMQLYaHvN9r2gWmVmjnFflo4UOkdiQUSreJno
x1Q8+f9+C/elr0ZO2lhbwTMiog37tv46H7Cw1Dl26+Z8m8LWViRwgN01Gu5Hsnh6HIsOg+gguAsX
jNOcWhIvUK6Lin/ARuUyOaOvMKEuvuOIZQxhOaGVlZvuc+6/Teg+EtVVagbNFqg8uAqk9ofkyZ3K
iczDyeipnXLn8UJvyYjYh8ftDCwon5Xi9kiT1LEIcspEr/0jFbt7pebfGNU1ky+rqzVNUSH8BPKI
Jep9J4xtm1igLO0FOvQ7hIZupwbXLSfeoO+xmR5B2zbkMpDDo/TyKLyCq8Az0duX0WbJk9x/quZ6
GiarOh/1xR2X+orIxFzbAcmxybl2Es5N+wyQni2OlBcKk+r+SZGX/KwWjhp6Kqiqtm0bzTCvl57p
shx7qIuf3cnmeFhNc4pSUUgr1bVCyGNmcAVTR3CU77ac6eiy61bQlDdakN2OQKrPnZT6FWooGzzI
not9lrPLQSbmd0aP+gmBty0PQJfVkHh9r557vtkll9nAWPrgLL379B5HJJU8eYo298NALQTVqVnM
HHXyjBrehKJl+BSC3C5W733n3VD4+fvmZu63Uv9bTQbYubxcJwjuqgEC17xZAmIBHlluOEosZxFm
PH30H3i7twp+V20SaMCkoiF12eWL4IJKrEnaxLZ2B7disPMtIxTcPWq6HaGM1cGmhZ47Vwt3xS+W
26oSG5ozchcANkCIFR90wmYR7Uv35V2BJuoihpC0Sq6A9v/gbL7yk7W0urKn+QQAqr7PMI77qdzU
aArZt0jRaoZ8/enhMDMH0ubX7Xi9bF64l2k0Rg2+jNt7YqaVLSQpMM1l2APbx87yR7bGevLBGzbO
/UD6dM7rRHZ8YDuQcOQa33Cxa684uXohHK+nKBqxZuhk5bFWu/IdSaXEfHMNs1aH1MiHYczDcKd1
qOB/sDkj0NBB/u/GqGlxh/NLqcrmbBfakx9FRmSjvpGsImEBRgy78B0i5y7YFaIqMEWnj4xXP0mz
+emAKT7zngI+vPFnMVVF1NVefUe2hqETQN7lX09hCjBKdt7FoAjmAdf0b67vcQPeLuB+5URw7Y/6
Ty33zvFLB4xwyUlMMot3IXOWIaykk21wDIWSxS7FdYjkNdjGNFn8OmTmu796QfnNt5M03rrRqpui
saGdzyumTUBgs1Za3AdtOCaABSbvLQasGrRQ1SXwEniloZ88PoWmfvKBv5I7bT2C3kO7IEDa8WRP
qId5OdscrHKaBx2KbfI9RPyZRdX/bBCYaF18fsCwNLm0fPwBRuFC+Pqb7GqftdK2O1SAz03QrG9M
HKhI8NH1EQtnRS9n3LYf9s0CRJcyg3D6UY4LPyW96AaQcIZesELj51RuYFKwZmAabkH5oV5PhdnA
YUmTGt2h54+zgg5NYhpG79NkrQJfRrrlOntd2J2Ep0A7LSgBenukGo1wasU2iw+k2D3WYcxiQDyK
yaPUxyJypXJaMEcRoaAHWK9XeoUFCLcStETFNUgvp35PsuZPYOqIhS9Z8EabsSDqZOE/d72REmXo
DYxfNo045XqEB97iijlk7KZhzuH+rZHw2pce8iUDyX1Hjl7HpXbTx8DDZwtiHoNHo9K2egiWYiWa
osOpyKtx+gvT2Be9eDJJ3WZjuqPZp5Xwhvf1WSbtYanJvfNLHT8YS+pVxuiGvVPO7odbM7Tjjmjk
wlTv242s4ZkoDPIahPlxI6eupT5XWPlVcFCaFGf4Z7lDpdEZZzwUBESSLwiF+6SRqw9zq8BRgM7B
PiJ3X6jSytoGnuvJOnbp6vINJgr25H/ZvoBR+Fi1v9071b1iIa0LLddCAsevUVJJ921+9CygYcQq
GEBR2l68q25LnCzoBdd1fna85N4/pa/XdKWAcaRgMZ79djJ7NI1xVVuvlA1+7Oi3bLO8FSshJyBW
qY4wRCuKQRQtPiFSxk+bnAUWe73uX/9ico+4KJ8jgx9HsIErAJ6A/yIdLb21J8NPKy6puk4gFP+A
PeDkynxd5whSSO/aPq/AQVOMg1an7J3Ejrcks+vi4hM+IRwqR901bTXD5joM7F/k/6AuLbtRwbNQ
+YazvkmTCO86F/qtGDp0PfEM8DtbhTU2R8zyNEGaEJQfAzawN4Mpb8O55YvN6f9L+hiybORK1sHx
Ksoz/IBSeLNAS1amoVo/FFj3N4Mk2pKYxsWI6GNra2wVZ1iaxAhJySHqP5HR39G4h5dmPCHGhL6h
pA9N/uB6CCEmm8iRzKrRZxIWRpOL7BHujm4n0YU91+4LgxgZT+Io85tN9sWB38Ntp5+FiGYVUOqZ
tg==
`pragma protect end_protected
