// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
E3y+V2loj1lOEH+bypN7lGpMPTQuK1baQ2Yn4HAo/5oDWZfF7MslMIe/iueC
POecBUd3rbcHe6BTZspHLLOghiU4nLu+N+hDgofG2FawRKGDFLUngzijq8WR
x9HJ6SVObXxD1c3GivxcL0TLYeSntcUfUpDrumCgiRJpTYxnZFua4S8/Hs36
aQV/u+x7AKYNJPsM3/cszEiV+P6n0nkJHecdlc9NydQ1arTEd+/w+cCb+pw/
r9cgdGVWb46zfCB+NgeWc0DOFzUkAP5ot328AHTqETaSCr94AS+s74Xq/GGl
2gxSka9iId/ma7AxK6Vir1rkeRLABAsFn9e0bWCmiQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
nok3YAtmGv2PPJmzP0Xdjh94ccuChIXcSpQ+MnG2S8NOO7PYCOgQOujNxC4P
G29Or472f6bJH8NueQOoy+FRRrB8xRDNTzn9QeNsD4VJzCQ5H6Iql1Kqu9ao
veBbtnq6de+2BsGMUXI29grbiGRBdpy37ozYAiylF/rAcKq0coovBE6zuGwd
BhhaAk3akxZgjVyGRXH3/ufS8rM+vnIMIDFqH4XxDIEoS12sNTXxSQSsJ7Ft
HmRdy89Q25kvomaDqkEgTI9UWnhcIyKODq99c2lFM+z13paueVnDVz4hta6z
2/6e5lbm4HsPXg4//yiwyPNkKFxF8c8R/KP7+WeSTg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
pqpkDW84RtEpUeAv1L4IUyJPutfDDFN0IMM+YWJN19+LzRkZbreduAGbZJcP
T3HU3Kj1X8MLGf1hBELeOFXeh4lbypzq+GK61Cf6u2WyT+jx/8VJ3vdqTErx
/EsNTHB9syB7P2UwT75x/Sn0Ne3MMCHpg1OysxJTlUk6zou9dkeWRqEOF6ea
Pn32YAVNeOBxZWFKkZAe1/rkyN7CUb/QzAN9P3KEoKtSt0Q2MJ5Og6EqUNip
zQlzMnmOpNirl4pj8oDnYP5NJVPuxtQVgzH66eRxkLDq1gS0FMvOtv/q7Rto
vFWzVaQG/+NeevRMyadk+JixIM/koIQDFPElmWiTFw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
J5iMpN2/D5xFHK+p+OdNt7PrZJDir1ZUMRASHwtRPVtNpZYU3EepfS5c2+qi
88nb5aOQ0JTiV9lqxYtqDNctEGESRDM5W3Z/lCr33mpMiQPj7izcD9pUvSr3
grU+CGOs2URIAh7PsDPQ+unhHzZFAfndray+0iO6HRHhj6OVcUk=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
awCRSNHhsTL0/xdg2VagxNYQMKnY8a3eqXlvUCBC4UIaVEck7LXCsoPxvZdP
deg0XeKhqkHr1TUQjeQt69rsECjFiF6C+7UfvwVRdl5os33B5dg00SMuF2zo
z+1uQPuqsGyhH7nnbogzCw3Dk6uVoPn3EnxKDww/7QMEQIOymkaq4pM4BNr1
hXOS6WGOuSuL0Z3+XG2j5lSxsQ83Hvl6kxn/Y89B4h5rPSSSzdRSmGntR4ul
k11u2lpBQM6cX9PvtVsqnnPRabLGtEqph+bos2z5QaM+x06Oz23lco2KsEcM
hqgnE2m1tm2nxn14OOCRtcl6mETq0IY2GKjP8c12Hz+upD0sgSv//Zlmjmcx
vS7dxqWzyw3XUgUBU3lq5/16QC1tvhF6FSjrMVxIMKhuvmRTsH4w+MPdgrVk
q4Sw2Uf75PwqbFSzXl2nuQOH5f/LX8IRAlvhwONgYRz9f0Ap8bJa3MWCi9k8
p5cqHR3JtBog3fDkpVSXe9g2UIohAIJ7


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
iTrMZ+ohok5x2/Op2QLJmToCi7UhTi/lWMwlbflZt09LcIT5pYqqD3fZFo1H
1+Jsm9oeQDiY4C1bTLRSrjlAcBupRFi3aE7aAJd8UBxfcgd/dFH0KoQUYeVQ
sXLpztgKmn5xGWMZd6L8w6CR6q1Wj91klRa3lk0JI9Mzc7KWsrM=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
XNsBqFyq0qRY02yWfo6KrUVLXXKdLVGjJ2/ffkMmkIraVr6Hd+17fWxkd8yR
R/9pEqAj79YFcNgc6xEjUorpWxdpIMHvrf0Yl96l1V3GCSgY+uazy/7scThD
uAqdlXbVdKFVhZtqZosJDRVPNiYtPaRzwholXp9bUAuj86oUlhE=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 9008)
`pragma protect data_block
Ow4dAx7o/geE62pj/2ECJnGwS3hnPBD3wNjylVKsL1TtgXr06Tl11Aal5GYZ
m9XJlBrIlgPwVhYPT9VGCW+j+PluJp3L0LNLiBK78vjNNqWts+qaI/pv3bHj
O71uEFKZmF1n5/CLyOuul8UsWPFNTzlf911RvHtX5NG/QDyYesnwk6Ov++cN
CNZAd2P0fh1ZJVdcoBAyzhBpHC7WFs8lXGl+Tj4MtcPz041L9FbDiLn7av0e
Cf5H9dF85oQ3r3Sl7zGwOs3gMEwRpfBOVrys5Z3enUFRsvOOfvf0GRmRwvmP
+rYdo0S6cs4DhA9HMBqToWURBND/hqXE8mxl7QtXwCeZNptEYMTQiWhiMRVc
4I0jqGB1V3+FKxT9LFEroXCHT2jWEvj/mhHDMrfgnI5/sjXaLbsAC9OBwyzu
UKkJd/cNVGvLdUDGsaiATm9aTWzZ4PkDa5ayF8jwFTQpMl5m7N3Zy27CyA7p
pA2ppZITAxzDDfyX80Flu7zc2zwYu0U9WfZ7cnjMdWr9/u3yynBfpJU4BsmN
VCtBLS2rnslnOLF5bXyna2yRQQTwayF3A4V8fo8epFjq7NEMc0w18QXdgNwB
9Un7InsEJlBkwHDI0nAls+GzJJ5vcKBBrAUpH+s/CrwHxe0OCCl4XOzaiC59
2FIPHSrOJfmabczkXP8JM1MxbzYVJF/EQnShcVsz2fAuxUD4GgIcWnR5jHLm
1HsTsBQq/VaMrbDVNCLKaTvj2N/q0EENG3YOW7glon9Y36bbbzJ7QFJ9HdaS
WQq3J9qT2C5vRZzTDXF7kn5u2xIE5qx+V1ZgxcdXIB83CeE+5/YSI1w0UfO9
oV1DvF3RPVXpxvHJ320nRT+i0ruONlyTHTyc/R8AnJm+iFzN1oscWq1IdBP5
usNmDXBkIMHGC5P4yI6A43e4QPokjY/iFY+MiIwW+wz10+VW4IQrtC6P8IFf
BKRjJ8XEL9hTyJop/C3wmj8bH2RZ5FIX2hLUfeTflmTlWTS0dvksmij60nn6
7I8uJYH9l9N+bB87N06SpFKaaeubqHwwpo19ueIG+XmmRgUTgTTLMuw0UbTZ
occN/ic4FR5rMt9WqrXkCrndx1crB1T7OP1Yd6m8+UYGD1X5haL9DHlIoU2L
c4fiHwTr+Y0zVLoBPz+ZL+9NJMOnqtnDDsb0omASE0AgNmis8D/uzwyCV9UJ
/RX/2d2nPN++w9GteBd0RFfOf5HnVj+VNnt94giLSea1+IBVp729UXRTMRrP
EiKgQyxVx4a3BjSEj1RLY/i6Jg/tJpl1Eb0zZq2pP+Amdf7Jsry3X/nFngi+
/nAkWXEpxwWjczXU3NgNieS83mf7wcCrosm4N13Ec13T6Ym9F1Xy6QuOrSbY
rOK3HUsBmN5LfTvJlsKXHx2sq95G4amn89pzSzmFhrsX7e7A3R9DSDCXBU5q
KM86iMot+47tG9OpjXuqiRNQRJiIy4RpUhXIjsuYBvFGSLamnUEbtLP1RcmK
DOV8rxeMRyqTSnWzGQIVHvaxxliLWx8zvW2aKN73YEWToZx4x4eHTQlPbfVq
ZRUB6XuDNNCOm1JPDa02hsX+nbe9hOfGv/rLDW1giBk1e7lxx0COezUZgo0b
LYc0nyVup6gJURAUY9C99Q1Bl1kdc8Aiz5gec0Dwc5FM/P4VWIRG57wu5DIq
4iYlcyh+56wlp3kV87gbMkwPBC5mtK6LxRrQd5E1uUpE+VBm4f7XU4VNX3eF
TRvCpULspd/Wy5KsrjK4jrlqKt1qQo+xdhN3wHQ4E2FyOiq05mlFw20ota48
i/LWDqAiFl2/X5MOxR/Cg4jv/HrfQxN+Zk13DE6hTkXN6b+K8/U8J41MzPci
C/1e5sGJVu+9k088H2yAmq27c1mEthd9aoDGljEyeqyl35u/LWWZQPS2AHMx
hcnRqbR+G2mzKXLzqQBWKXFDhy5dZ6BjqipoQG3IBKHlfsGgYvkK4xo0imAs
2Aj/GOUqlD1zEfc/vt95v2Exx6k+LBU6VjGp2Y4E9HCSY6Q9pUV637NaypSt
WYk+G+heyYdsZ3GT0+sYF+ZZ4j26hdLWNVScprZCVyPCk8ctVC+zwdAWncB7
7PhC5ujdXkbvsINppce6Cr3adfEIEP+u53lXyEeKBMfU6710lFEUe5j9na9J
fYbJ1zGZIUT78it5/m9rfQXVHDbG8B5ZNPmUYTsf4wgRlB58ccgZEEN8Ejsy
MpZhvaE45ludfZhXaT/cBNoqHJSTpbhAqScKkJhiYYLDLJST7qvxxZV87qu0
XyhDszi/sdf+uFi+sDpKMYxijqAGJClbJracsNXj7VucDZjuyarYkPzHWSj8
lKQMvXFstnOGkObZw6LLWYiWjtjUJMsChDYVHZSpy1QnEjI+RfCLsnhj56rH
Chne3NU4cxEyEesXD4BbKoRuXClVdgUMw1VGxkJ+jw+vMb0qAip5G5zyRyg6
6PKm8X1NmWgtEihEEyRf5MgfhIxKxRVpY7me/J4AZ78j9GhuYwmM93pNB6UP
x6winKAjTMnSY126KRxpPN5IsOOzYLkMJEYnR7Mo9/W0Bdb+ZCDtsBe1uUdk
wiipsmyIzJUOObWBxZCxQCTtnOzX4aCi8jy/brUwzf+hJ+Nesf7EsJcmpxhh
DkSl7pSJrddKsnOpdwUft0CnX9fKH6gxnCWWjy3uhoQxrdX9D3Y84B7uO81E
R3IDG3ox0KCnGrd5yjWypUP/5eR2sw00qLud4YZjvDV1Az/kRObM9TkH4D49
D9+5tNRjKhxyJiDMc83wJqaJDCohA/K3Kgrijd+QP85vhEWFxSXNHJ1YmlUq
3QIoB/mbuJC0v2qqUni8lrLI94C2XS7VyuKPnx7BkPmO8oFixVWN+IoXaDZ6
0UtrnwBgipdn/GcIFqfV6tIa2X7xP6GTQ7E3wcK21C/0p2QHmos22hU1iUdZ
EgEK3XYxdNomO1ocMEHQ+K75lF0m099kjDASx+UKVAeUjvNrIzYAo9wT0zJ3
vewzrP73jdKliSYha2dnbHMah/55RU8MHC6MwrFLZTnF1vRB8SkJ56BHvTuX
wW+umJ+duBRprcKJl018nbvQu3nv3z+VVRo04K1ppTfsHdwbKz4JfJCx0l1B
ErvdMBl+ylW7Qf7BVhBFCIREBhgsyMe2rdlM20Cp8Qkh7E0T+qvsr73dNk1B
HGNBgsVPLJAbWusIfFj/CJXfvsUamaR7h6PmNNs/vyyWDlVOyc0wTO0E1ZaO
wzA8MVxGQwLBvXluuHv7QfrKZCwBc57/988qAJ2Vzml/Flovo6x7ZJdg7bhh
Cu+B9HauGXBmNRDrALmkVyFxAAVkGPrS9p9ZZyeeqHQ577sYOLTeKQ7Lx4+O
B+gxCA87qAcJf+3TPBNSvyKd+fWV17nQuayCiuC3X9Y8V912ZK3tLBl1YBe4
MzL2PD7UlSHw6QaH1XTliO8Lvo33UgUGe8xNganIUHnKTXYsRh8Yk2dl/ii0
klO29aCDW7kQkl4hnTMYXCvNKMtnm8RZo4CdNYtaBi5m0KFzQbyFYXULS+Ed
2+jyqAJKUUCYhgK+f/LOFpOag3xzEY78/7Ku+sKDwGsT3569xRLYTMXPtreN
4dk41izdrf69pF11X56P1u3r75ealM10QOnamuwx2A3HNIhrT+/yGnbb82mN
zc8Hk3AA7HGcLL8FPtQ1ljgK35F3f+lmTeb4Q7oYtPPiGPlwnc41DfuzSLzJ
AKOs6MlBj9kfZm/TpbMskMwc1N7K/ElBkrkFQ72fZBViNypUyXR+0fA4I2gg
wzRDjLKxIN61s+gp6jbaH5M1gED8KD4xphFz8zR35vMnZUpAlcrzoEydCpAa
0iKtrIbJ7OUEMuQlpVpsUbz1NkStoJ0/QKKvw8olVEcaV92VXU64cgUugGkf
S1xeNYbjvgx9JP/L0p/s9KmHHX5MTbsGYEjpIGoUtYVYdS4DO9/hTkJ9ivt1
3LS8CBA/CmWkDXWtvx5ufGRDf44qvKTr2xS0/zxe6rlq8U7CUIzxO5R6DV3i
jF0GjRKGDV/BKC/evEjp0l2px16d2JeP2lphuG4vy7mTKYH7JMkHU56Y6T3K
Qf28bfvkQP+orSOOb2hiS8AID+koKdNy8EcdWZx1Gq5I+1YzuaLI3RxtrfEK
qpy/5jd2xSPttg92Fn/R+F1HpIpCXIptYQQKMN7ov3bqvm7af4Mn946KaFbq
MlPk9xO0Fi/zlVq9Wlk6RHw2M+rlrgMSiuCb6zgH8v4LdWzrpChnigVMy8/3
4hYTvSd/l9aKmEM9xAf5ttK9D0bIGTdj7RgDAp2Uyo5dgdhgUbIHTQs30u+E
sS3nkn/jw1ZRRyKMi2ahpgtjKsdGmGuHIK+x0aCv+yORYmHKtPcgaXjPCMBX
FZdBWpS+NPvEJrRAI2jgb7k7wdFm30Z+knAOveaUIxY5KZB1a7EahQpGp0bJ
JSwD57V1jTaul7R8P0DMgQzqwgQbjP5/7F0Bvjkg8T5614Rg8CDXQPTWnzb2
4nAsvrb82IsNLZCUXnrP9/Fwp7//9hk/6h/y7mjoiBqFP3Dck7Gf++cYTNIe
Hipyi5J2x65Wab/6W4ci++C3mIWcl9H2JYMDr+jNSOFOxFXBHjZ1LLKHzgsK
QRB0MF4Qka7JzJeqyXp2lvV1et8KkYP41XJ319FP1UYpbxGxwEti/Fscr5U6
nRf39ruevzjBMOEvAf/kCLk1S3xil1UyX4h33G2NPwsrNPbpI0E0rN4O5QKi
xvWiLC8V9r7Bgr141RZWIzqW1sfGxiU1z4KJNRfp1sYLWy2dQXqEk0loi26q
2jGDqGjLol7hKoTUQUwUkQjHsuCTIiPB/7F0+UTe5T+bZUa8TpT/DLdklv+b
xNQw0xOjtxrGiob8bs/K6cYphGjEzuXsafGFBf2QGzK7Au0lDlF9IXQUqHZf
yGLfSI15mwqc/rY9Zj4ZqQKXeggHruG37NW+zMJSOO0U9l+X1Z2dKnzZbhmn
oJcYYb+CcLUw3qxfwosxV25jkCDC5NUi404rheTycGipFu/MqCyHz4jtswDt
IgWTVdAeQM8Ncbq1V/R/GwMRdK+eTFgkrvXcWqcKZMOpOFN7465+N8mVVC1o
0GpDkUjgyT8pCjo6sU49NVOHg596X6wj99G4qbx1oDrxhzS8O3lEN4K17O5l
0OSyUnE1Jll4dxPvFPKKQ94ZvB9bKkxLbKIlsVlMwimdcQC0r8kgKLQqIqHu
u4iaLz3qUlSK+NjXBaBjQ8i60xBoatQkdATsiIFaDwoJ1KuxVE3Pj1TRlMkL
KaE6oAWePC79stsqUv99xkfoxHDLlN8ruufGrYr7Rsq+gOr0FN7eKkz8CydN
bSOoOjiU0LSYUzkA+OvTvKI2Y+38kiZWoHcb8Kcdk9g8uxwrL6+3uJeJxwtX
8fxP3T+T95b6RtkfT9TGLqSPoO37/v5InfVOiZWA1C96YaEy11A7TzjK37A5
AK4GdkcD/tcfh0Sapy8TU6NZYqlaI1t5V3pWgqyp9SwU6JfUJKAyZpPv8xT/
/EIdRvW/w1s74ULrzGYzb/Y/LB1jb5HkloT9qFsNT7q2KxgsIcnhBDlCyiRY
+nx9FJ2TEhsA455ekJnGVxeYDNEFbPe+PJUs3rIwGxcVWFOeIj2apbZJtx8j
cdHEGwJSuksvaJRVNFRsSKnY+brrHIpnAHB8p3HvojZ+vBNIgTAK6gmJC1/2
wytRtLS6l/EOcLmcpDfuLiMaNosT7D5WkdhbxonvSDlFy764iU9lVA6cgUEs
jvOWI11PsR3/EhJrviG6qZc4w/fR6Oq4hVxclSjpRM3+2kaNnjjnlLjyZRhZ
qNbvr4MpKxZmkThT2tmeuZMKq0/JrNJP5bBE9mbIXfkJVViCRN/QuEzCIBnd
9K/kQaGDedEwulRMSPSBIZ03nSBrfE/pHpWskmQYd/r6bIj1zfTQ9i0TCvN8
fnNNV7xp4L9g4UsKOjCcEx/yXmDo/Le7FcdoWyWlAQxD4bXfa5tvqROKVTsO
u9qIi8q2vzRpeTYV7cVogtdjaf4kEN9nrmK/DacYhlTbLHwt17aBgQkZPXhP
poa1De0RCtTkZfK3HQAfJbWO1p5xfNQbZYR4dkh/exptaVTgknQm6ZFohXs1
aFnMEdxRhrGAgR89LbX/uSfnGLb0kQdModTg5CHQq5WhvNy81v2vOZJGRTrL
4a19JqGNEcgtps09uNJPVm+9Y5c0M+nEoF6z1CcqO32f3bimtfn3f49TEEDl
NOS2hPI1kBRiRK+gTV3NALdZVhOvWsGjSXCYeW5jswwgcFOh7+5FK/6aVaEv
JMaRGP2ChcYfDW8a1DuD5H4nFZDwMhpOf/zDfu0GGX2T/rP+uS/sonXs4Tra
lhmH2m4iNHTh3h4vqim6XLabaATsRZGsB8iJWrgeQ7j/EFsioMKeVUImoZtU
kDAVVuY+mrhbViM5kLLVm9n/lZNv3x//8h5N6GgA6Y2n9GrRvt/Tl+EWxN/9
Ujb+y36YO4F6WXZkc9sZ0Fxvw9831xx5zjfLSktCiURTpQexANSR+99JYuOq
0kXWOS1XAVT47JfnM+H4+PNhNNY4Kg/q6B3L9SA9LCJZ/EXeGIQwXG08GInr
+l1L6sE35ZAQz49jz0oCI/5FNa6QwClG0R0v89z1pgFmClj6JJfafXjk6fZa
7+LyP8O6UoQYLwowXGdvOY0DmZjvM6V7/KhtsX8ZECoWUFYthKqfQBM5prxq
jzxHJ02aiLSEgm4xaOSFdOq4Ta/4SMjkjxcd/vEfMFWznL1HsdEly3YS5nK1
BTukD9OVOkB+Wou9G0kSDbRO84Dno9i1VIJqCt8FGY+Y6YSE3Y1XnbyaPWob
Y3qUaPPiTNs4piODy9g7qc/MtkuL6kOz9R8YtK43yE0/He55L8b2pF+P/8Ay
lxr8VvQyx7dxzs+zsbpoLfdf+C3H+m3XrKtyEOJpEp8TZSVPAH0mOnpDdF2+
/sERYMy187etaz/2BVe4J623EtIPa2H9uLICLdy4HgwQ08UjXRocxu1+GeGi
MdcIMXwHQ0nmgaw8iHDoky8FaPo6xkQgIoqSvFkNT7rtUXKOqoIdThUEb6eG
lsnMtz58iAkbgNfwwOKa+iczu7+lgFc7KhvrLJdvtzbMJsuVm+deIaWVbmRe
VXHmVtHqsrmo3A0Ibpo9X63B8jZ5UyB/GsElbIhja1CaaF1ZzgWB0Ab/yI9Z
Pl/jz9Ua9Yx8WHoo9rY7d7AoI5Vep3Lwcdt2VlZa+OrU3kT1XzCyB+lFTYmG
OIR3viRz4SNsH1eYT4gPcDvfVNd2atlRn8Q9lKrKachqLqdsR0OTOEPTnEaS
sjQCKQHVWO6pesQ53WGrfTTaK9Z6W0EG17mzNWROYpYvng4SLwEaDAYeXU0Q
CcsjCZ1RKTA0uUObTNJaXZ6Ja+tDt/qrwZbByStBRcgOX+6JgKgz/vtwaULp
0Meuy1VRnnnbjbjH2+82a0v6NfkMZnpYi8JvE0nm+N3+txOQMICorEhgeQTI
IMrAfl/qEoK+ZnrSIb7t3lnYtOhbZGxzYZ0dB+B03Y9wz5j7PEYIw9d4n9H3
ISDMCBFo33Be+z/bLfLR32cgBKCD0zO52efRoYFgySh4PY9hIDngWgen85Jl
+C/cO4Up/WD3jAKYuUqSoIV2pZKgo/ayufNSyxyi9VEj1UpWEOAT0uK+tYqx
l0pDrw/jWKOMnsX7RAXlPIBlyuw5tDXb/rgjDzEG8EWiJgenBDEDAPo+BRMs
b1pO6eCoP1cXWaJGbPMuR3ujomeagzX9V3JaUyAgjVl2QQtXC6J7FFG0Z1CH
jB05Rdn4pf5feS21ALtwTI4v186sQ7tyjESrSe8yZx2ia26dUo4FFsZITd1y
xkHapVIIL0mJCQV8U4VWi16+X3S0iagtFS66BsKXRkNpVv88npoawtwGq5pj
PxzswIOX9gK4yl+2SaBssaSRZ3g2wb03Y5VkG4mAw230Lxb29wJi51JCVqN6
XY0ezAbd0YSxyzQh9qSLsQTrhpsH0s8XNWhgW7ZtBCkh6bbRWmc0zLzPE3U2
mJ+1PSu1Ox67DpHXZJCMyeeHnnqYDb1ubRTOeWuzxgaWvW4ojAlo5arKlfim
8fbxuzMKJey/uybM8/sMJcWJmpKTpIVPJmCs2y5p3sDAHQFnsxwxylK4LKTc
4+uRW05aLPyxM4bmkDFj66KftQ0f54YJ12fPSU1uBiq0uoftqbqAMyYZBRiG
TdFrOEeY98k6LfEFfWoJ5aJVKLxS4HwykKYuzgFx/PcSPEvsAScr9eGxfFjI
MDOMlztO47681jZVPwREUCQcXQWuEdc75cNSMdEV55VU5B7jEF6rItYiBDuR
uMTLEN21MCKi0c7/mQGTsjKNV7aIq19HMDk8iEKcHROL+dtnP9sNZaAhcdjg
s30GfS3lEhq0/LZQ/vn4BtHerK471NMOmel+3dGMaiKVunrkj7bs/3u+bSIg
CeBbth06jRnhWF7XkMvJ87/xdCykC3cqNfdhb3QRsTwuYaK/rlWAfHmFcg4n
/VN1nsqsY8dwhwJ8Fck1QeFJDtSZVenei22sJSa6BMF/YmRLpJymwRo1ih50
WXckjNQw2MYuWVGibEN1ZERYQ6IlYfS1PbrLniWdGVx4Cc+hmQi4sreLgZSg
GV7c8r05M55wJ2/yofX83uVkFmq49PoFFUlr2Heyu3kiPRhcAqTLiuzHeO9X
3p0CyUwntPPALG2I+YyicE5RH3KJL1/Vi3Y36UZx1hoLZ0S1mBeXG5P+AxIz
d7EruLXA3DEl/8ByiMIYlChiiGzm2jj+t2pxagAfQ4BF0Hnmh+fW7lh4/e0d
ze2Pm8gDy4kR264+kHiSm5oo9IkjFs5CmPHsBqHYqd0whZVpNfobm3HzBBia
Md/4h1sfwWf20mkaGW5sE6aaLxg09LyDtqoVQOdUAlatIfsRqIobJxUeVo9F
fz8oYhmy0eXs+T58jlQyV0a10lohqeW6rnUCYvm2eS1W91+YV4s/VaEI1W9n
MFVexZ8U6+Qku/iVeeXgkwL0vvA7+Y0NkM/UhxiRV07u9NzQFu739T33Kpwg
rWeiUKhIUH2myhJ2J7Yy2kBGjkTWqwlpGMYhZd31OCPF5xSFl1m7DK7VX9HS
hRC5apeYQxvyq6a/yULYDZjXFMjVr0Uz2cgj1JDBeJ9eYd/ShKrFifUW7TlX
OSTQmmaoljVHHcrqWz2NPQbrro42Udm6nPb3lbNxCr5fa7WgxYTikxedzPL7
liIROF2ZMOMiid4902uxY5wNbryU+2gh2BxyfcepFnNFn7ujwoWkyWEy327u
kYVo47ThKH+gQhN+7tfvFUnUrZ/RQ1HJUBy8YiSnWWhWZAiBLDlne6QB6IdG
FGbeNvpa6q8YQGnZdtPQH/E8ZRPxuqpOi3vTTZUNKd8R+2IlHt7pXxy8gopF
CUi31RVUle9BUnS6W3nJhIuuQCBZQMsw5cmgkHPXvrqR3aQhRacam8kkapgx
aEvDxvlBDlOXPyXVP5dRckkqVXb3/jMPVOvMYJrtdAdLgvYLLS5eoblq5ASY
spVn2e08od14QL3j/G+5fjSvnloyZ2MKTs/evu1NA9KFIo+6KA1rNg0G9zKS
rqvpp4KS4DGxRzDgGrG+y37LMvtgBjO4BQZLR1PeTSUe56VaFjFUFIsZ8FI3
2yG6Y5zIkJpaB/cyQG99DjPi6jpnQjRl3xCgiYDHOc42PoZRRG/opOcoJt8M
ZjVrTwBUl6XTEzb0eo1q7iHkwLKwNUnOaO77MC7P6Bi0J6vlJAJNf82ey5Ja
IsYjgldsVfAJKQpm7/hVyOKlpYhvex3ehYa7a7K58yFAeD6H0Obkjh5JpdCE
FHLjgtOYemZBt0ELIE5Be/FO6/rl33VwLNRURMSEAl2x178mhGdAKLEjimb5
vJ5SzbTGfH6w5WWNgXy1W3CKFbYirGFn4zStf1YPj/ljvmOklaeShxxmAh24
k6GdyrZB/0CLUshTd9HBHZAlAGjkFjeHSZDT/4opyKdXHCBVGztZQHVdkXYy
EDWw1XFiXQabMFI/9M9DIt2MyqTf5Kxi9JthEuJ3/LblppJl4XoJv6GXgVeL
9c2xmU/46IV3h5cvVokde8NJ2wenKAkaOWEdYvx/+mMF+aVgQVIpLx2418F3
+f82AeMdctH5/3PsCbsqgxWN1MqEJEXdhgANylcrFVSeJLRYo5oj1sxG7b5D
sIXluk54g2PwwEL8LdflewJot2DH+0NabT/Ppt7J7gBCVWsyvmhE6SOmHeBU
pDN+dmM3Sm2wY0YGm1nKtjRY/82qI3ZD82zHFpcN6j385Z+yWNkZCWt92hT0
QHwbFth3xUboKDH1gzAAgcLxwxpLZGgg4FI375qqDD3X0+Dan4lwmwXnK12k
8mSM7HjDiPFFEZ+PzpSbAHlbGEYiACyLv/CDrtEU/yyj+NveierehHdkC9xM
68iA+GfQa2bgGjueNNf/PaipIaaxaE6oBgtOgLdIwbGWpV21utTOjqSRRrWC
nTw0AyuB749sQPCvElm2qWN+GUoiMHpyvRFM8q+6GkOPt1TrkC3/TZ7oCn+C
hMblQm3OtHF75W0FaTPvGAE1iZI7KjIJt/diBy8xLrimvyFtHmZuzx0WTCt0
yDM7DTTd6CVvzT4eaeplkxczA48M7C9mRbAxshhC58hs87y20pCvdg/Nyb9u
ZCgL+qDrfiUMnHyt/h3DlucXyRP7Fdm2meveB6EgFHBzxpWx/JuTC0twlFMT
Edj/GyDNQPIUTydUP3WCFuoWB4MIYDV+6NYGYG+1jf0VvzmS9XdO/lGzDZpp
PWLZyAi0J3U5MuQOU/h1hH58v9qboBI0jEUIZXo99cmQ3ZrYNlDTb5pewlvc
RWLHjuqtNldM/Pq4I/qwE9uDOBDo6SK3vQ1RYVOGz0MbGH2lqLUXjns+QU2T
1jqE9MJDFNnWnB/9wMLCS74n/w181F4mDkLups6V3d+18D598S63nFff5f7j
ieNC28QXdP2MW/W0Xb6tpKedh6HENDEdmisFhVhPT58nyIF93hGTDqM+GDsT
Am3ffJ3A5CZimdgbrEsJ7BNH4Hx9udbKhD0AOeq+JSjRwsdTxyrcdajaE+Iz
bCZDVo4PjZnolLOmjgp5iqSYzCIc7LrfPzcYK5S3qfSn+n7dQHYymQBnidks
sfHpEGS6C2GWiKl6np9AcETmPkAG/rA5XVbi+6OfN27UZzMlVDjZvsG8wblA
39/xGHV/SKrXO/AGaB23AvU/uNnIYdYi2jG9JUgzYQtLRvwwc9JgvEVLY996
OS0iWj47nh8tMMbn1JVP7JUHa91AM5ByFbrLx5+wU7cssAMZSjKCcGbjm34/
CJbGiQ3q/eAQiIGoPGRlxWcI4iRfZ1eQ9lOqgGQpM2bAA/0wE3+bk1gUFSDt
YsuPYmSt/PnceRsrjVP2gQDT3+oU4QK7CAtIfLl+X3SIpjak+t/LtTnPuc+8
Anmwi43IJuRZxWNub0+gEZuYVF/fk9okT7lH9SWey5x8i25dCfPIvyPoaU0G
R3m5XokhLSH9auFa5F77+UVR5GsIkwSZXrL0NNnbNxSTmsfr5R7vxBNbqPXU
DunBMFWOTyRzih6A0yf7C7PVHE/Hz20x9HqMYhmS00H5VvAUiZTiyZKQWJwq
vwc8zffMr0EgAmWlP5JPrqiNVMsuyourm25G60v551IQixKeeIWWOEX9KfaN
hR5dr6CEEHphS3BZcRtrJ4WBz3GM5Pr3wxoDe2Q02WQITk4BIrvnfqRpBojs
gVjM5Ow2pIM36Bo0sUon4BTTyZ653FkG3UfedjMH2VblcYJ0i2QWL7ILQQRU
CKQUYMBbP4uB3j2/2KWyA1yuj2TV8OZMuj4X5OGUVZOlzNgd+XW3fqQb+BDb
CddhCEsgAYfWE/R/I0Bawk8FrSlaGSTockdlGdSNvdYSeg27Zu9dm0W4FUx4
kXiQ6UBQoGhMKStHe7uK/EkFkePIeCoEaKXDZBduwDxgAllNe6J+hACzuCl+
bO7vILGNDNc=

`pragma protect end_protected
