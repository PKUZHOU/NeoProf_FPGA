// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
TIgY77YpLYlRxT3tRhoE15/Ppu9cJ2zAicuxUIyIpvxkQyep92mIK4EZWBO5juu1
lUN2hJykFrP9TjZlJch9Y3lwk+9hPkh6xZAFTfelsqlcIVfx4hb747gmj0pizr8c
vxp+CURfg4jLq9C3pmXCEmbKYA77sWb4xnoJcYUXlLw=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 44848 )
`pragma protect data_block
dAecJTDLxPtp+QHeAcV3WzFIM3eecsD5+8tH7zQYihtTwoNZGHhVP0VYWBDPlIfM
Gx416VwK0DrohAuO0/fvSgxS9o2dLRWoEP/TTKUJTSaVOp12TbqS0p5aLT27BqKJ
uVrAev03IOktAR1F50LPNDaMZOM7VuW0utn1wGAZ8eHYoFmpCkS6gpLcHtcZpgFq
xLCC03AJv50xOC6k/+5gZ5vqdpGLPjitN++uKnjSjeTj7nqUB0s6O4nptoHU4AX7
xpX2Yb1mS7tDPWgSb7b1G6fZWJWZp0LfVuv3bxyuIevk6Uq0JnF3hYBmnAoaqEiD
4lpNbORlFUmj8xpgyDadS4olEzQwSKft7ISH5ULO1F1W3Ndt8ikorH4/de0zncie
+IWB8s2W2mREac/RDc5rH0upwW28eTAks73Z/mdbxJwhK8soNmR3NYZ3TCkZdW3k
6iCH7X7Brr44LrJ2k8HsacT9XS3qsUqc2Kh5rzki0b0/klcpmp7s301ngkz16A3j
oStRWbXz2KDwIU+90vnQwfnL4MH8IWPMZUCpEPVLbK/oWsGgrugF7UQOl070gUnW
m9b2Kg9L1QJxX9rUcZyc8dJ87BEOJdwx32+UcLa539rjSm6g/hVBKoeSyynAlGYc
OMLTQCY6LY/KrI/Ncg9UsipXsFKotBKtpQpN4xPBOayvOfoamKOHLv27zjy8I+ZA
TYJo4l1wFBnZyUY17PeheZD9pM3f2JgtcvOEINRstTX6024GaM2pQhnQ6WKhdJL3
HUHGYsWDaqNAycW3zgKCDaqogsEZ8u2hb0myIlDK2UBpQZhcwGcxw6fnOvEsm9De
/WjvNhpoQ3bgO3pLQzC20AOoiHAqJ5tap3wYZKgQAyBsiLS4FtnCdwEJOT9DL4de
dSOs9qA58gJmaNdgrYxCqx4sZ47wHdb3mFP031W2JCVXKY5xiPIoDzO1XF6c+BQD
6ZhSefHzs3a50zeUv8DCIC17YKac+7m0hPtmek5mqit6jFZ5c64mDZAD0o3w2MjK
aa/7DYSHIoz85GYt3yv3xGnq2Wufm4CyuOUelsEwhdjU/qQGFnyjX4wDYWggySmq
PFbDR70KUOYPCH3FppxmhnBOibr9CxyXIOKoKPFZ46C0jR4oc7x0ASEvQbYlcdOF
yaSTi5oShQru5CI0m7p3V1mydiabP2zUiR5YNVHtCF9eLrhtxJvG6jKizz28Fph9
XjT5/RPXGTn87hRam5RBr87Pi/CdtSLY1Ur2ly7hb/gxJwNllcRgthmPFq3Ufcml
iOiX6a+KBXwT1jKK4uYyAMBMooSFzMRaqm2HTZ48ID8iN41NwZM8buXZEPlWIreD
AcZkwo0J/PdH9bhIIE6DHXn84M7+auemxXtBDsftQfCog0NKmUeRUoHKktP2oMbx
r1eO1xsDsVF/VjiZAudoYk9gC2VPXqkv2Ef9PeXgKDdVC2oJGemtAfEz/dHL6ZmG
JJhgUUHJ60HphzlnHzu+gNeWt+VKlEGGl9lSRT0B3tIVEnHeQVpvd3u0aGLK2jVM
N15Bx1k6LJ5gyVxcOjQzH/ankkQPghf8xbtuSo3pgCsis0v0EO5p0uvr0pRfQPwK
YVMeYqIC/NjtM+JV1PYk8ANmaKAft5y/AKcuNxW7uPiJ0ff5CO7MO0fMbD1qJdNC
f9qfJoBTu0sPPj8RSFRBeE6ZnhINjTdx+MQOs9S27174X6VzlEXn0IvGH7Htw5KV
4FpDL6/O4voM19r/lTwv9cMv+F1v1QDaxHbR29Axbsuk4jMOlCvrPGCrALzEQZv1
v11/EH9aepkeJh6cQ+jifjXcVqGbAfZcm/3eHvVSj6Y17Rk33bxoawWsJ1g5Uxe7
+clfN/mlI8+A2gX69akGBM9giE47MEKwuEcgROgCMlTq6Lfmy3DtLc4rOIn30IM8
g//mtT2a9JeGh/C1mCpmdKN6WG/zhsJif6t8g/ZdHTOlAC970tbSf4E7jdOjilic
l9O2u5fzE9sd/oXvW+yQDAjK/X75JM8pzI9RSVrXh+QEH5BRbD50+QrIhuK8c6Io
8edKr0OPl+wHAVlKetWB3hV+k6IoU65HQ3pXlfDp3qN1yH+Lru5yurEXt5mX+/yn
42cq9aJD4/7pon5z0r0gtobeLKb11GDIc1KIG3ZNQVmHIrdxE34cyyxE0gqxu1+R
9WzG+ML/Q5UNVy30YznPN9KvKhFfurPHYFZZPPQDXC5hrUyc1P/l0aCcRtSCMR8B
cytoZ9naXI3bGn3XCG1OgTCenIWcG1jxtTRHSnmbmzL+4lgUJ7nKAcUGSSqalPRt
PGIUt7Kd0CPL+f3TE6TbLkWEuXhmlBonrK8mR2eZnBPKPKqYs6DHwKLGbmKPyUku
2smylViaXf1mCcmAvnyun/+WiLjSxKdT6Nf5Hw+bRAbSDnZuj0kZionkAmv9UEFK
fTWbn/C1ex84UMmIcXema2HgQYZ++ZWWAYTfDc7ern3wBBLra+zHrpieL1gYl+P6
NkeYn5pCoiLilU88pNrlxkXP5N560/8VD9IR2BWq2s8gF/kBmXXQrUy8L5RDGQLh
s6UA/AQEut3DyuAEKYnC1PWqT/XjWMkkp0ju6DB13Sa2vUTt96ozKlznyHp9/sl3
/B4ZC/bgCLsPemaBp79QlVlg0zd1O9cThP2/DNWaWIJ/y2LEYlSg2iYEzA5If/mw
o5qTGj11rBfIK7bbrBSmVRmGLlZwTXHD2bNWAgGftZIZsMRHs+KOGtMjPZ9lFU0B
pU4+Js52NCjPNUF29OQJJMuLR7LA5mSWRVbMww/+GcaFN9ZcMofpzV808G/5mFiH
Mxcz/MaEiimf8it8fRvUntsp09pw/QIOuGC5T9HOfdC097OKWWhVqqw8nDBCMUTU
LzoL2gZ4XlwDKP7o4mitIxuoge8buyScOBOhM5styLTJZ5DgMQ1D7yGtTkZWJIjg
f8kMlF7/NzVabISOcRm/pUqv/xWxIIt8XR1MePUCvsAgiVBrTeKfeYVq3qVMakax
7LlHMifOBzyUMKDL/IrDSnLxxYUNGFMMT4pndujqntDB0p1AK6SEw+/5N+zM4k/m
iiUpJaZugmp1BAFChMZPRSjAyBbFiMpuv49S9/AUCX2ku6+3TocpY1ImBZRttAOR
c71WU6sk/38K3Csr2PXOfRxRebwKbBQlX7ODd6NA884Z8w2V0HgTAdTSY/YE94RL
GkAes1IAXM9yyR1JLE006yK6qcuYCi57C4NS/B/UR+nhns8UKDPdbI+LhIMjLovC
q7Yu6J3Rcfj+asg6LvqxEYcp/Qf+IfcoVnRv1U8+yO/EVQ9p5DaKIkabmGHQkKIR
5c+4RTE+tDAHWz2m2x1W9Ur1qh5Bf7WFBcuhB5nbrvesAGsf6TeeBlVSorpZdAYY
5T8nTtbIC70IGufCCqfIRT3X5gWLnf/R1AczqXvWJKnxWEIshCtnV8CIR13Rl1Bb
g8pR/2Vfacr1LYePbNajPgSA/r3eHz4684m9ISdol724ZELiRPCo+A1vIgqKJjzi
hgr44fOE+oNRAjnSsn2wQXX4TXxWC8gfxrsVlCY3HFZsvRKhHWnMdI7owAlbDqGu
4Q9boKVfI3joFP9OQN5JUjQ3AT1Kv9OrXRaj19LRYchv0nY93FuZkusvYZA0qgQv
feYvN7gNDqIoabW3EBLUOz0gOTGd6QsKVYyyGD2z2AaJI1WfCB0NXn8eedPYkJx9
6utA4Gd5SmOA1ZQ443PGXQLiyDNn8SCfTogeL99C8RsE9A9pYrWt+YYlnh0ApP/d
b1HyYSYZw/XuKrXpMs61MDoR2Gcdn5lJYukwbYYEKQnzj5wYn9/HtMTE6qRwh0jZ
h8nETk4K0nFl/JdqalX0jw4+Hhlt64NhhxqRsHulXAyiqdo0Nb3YVmMbiag1FtFB
+oY+Lp0IgxVz1mDv8CumnJBMq5Pf/Y8G7Eu3SEJxwm4zXLSJesEjqw8PBsSvEZ7S
+lljRywoeUGEUyorchoIobNU7XjIH+1+B23Co5NJKtWKJYf80D6F6At0EQ2AXpbV
dkt/TXaRehMAQL3SqhdeZhPj14mqnzPB9CyS1C5+6Rth6Es5DlpM9As22lXfuHoc
q3jz1O8pMlL6cwTIwUpBy2NCY4gaD//uiMV0GHzVX/19aoeoxOqdzMVEyMYMMEw+
FOMsv8r9TDpyBsdpZt3ZJWR2WckW2zJn38kfN2Fh0M/E+Kkce1mp7yzHJsa8z/6A
WitfABxdWo+Z4D+qome4ZroXOowV9CazhRdyoInDpr5o6PFgADLa6ezcqMo1OuCM
c/ZAQ9HWZVU2zO0DS9UgCSdB2zR6YFjAW39yu2kHXTPfO2S7ERk8x2Y9Z9r65sAj
7SJHFjb6c61OaOexjUUY+jaOHbmFfPaOauUubNNatO+QGqNg2zf0jK3vW2ikflli
9vPqFf7E+cMezv3pgXUmUXPDFSG/p3yVFaS0nK+9XvhUicwFFtBif/FW8Q3OS8C4
IeLit8ZLb/b/v8bdtPZiQZyZEJ1buRP1MFCI1JFk+vYuZWDbbixh5NQZnC88jXT4
f1lCxLG2hhdJbg8rKh0yv52wakhJ6231yPAhVAuD/QoCej4JauWf97vQ1bJJgXqg
KD9oq2V03PmrPx0ssFGtW6YIsrbgXGRMsH54cMXyXobHvm7WFZCYlPfUCmZzkj4U
T2mn8G03/RqPspd822IIrFmQeS9AinYUlhkxlAWyhso7pPORfKLLnWna8m3OYVcL
THa1/scQcQtJLHWQzn8d5xPgxLPbE4KbDQZPe1NuZAcV8zhiCRMM+wZklxLgArre
QIMdM9UHHxI/9HrK/df8Z7Xdkwu7fiwC9FAAn3PgbFgzmR5S4xlWFSS3fCI9WS7a
hn6h/qfHywX7ZaxkO1p98LXwdRO391cRhiQ8ALlemd21Mf1ztKYs6JY94v0WgSI6
CMXjjrUOm1sa7hxUptPg0SZOCEw0iJklcBej6NVhCC0LWBD4GD9cS99vk4eqJFG3
ruy8hWx4hL6+kfy+yxGi9BsbPcqJZ7Un1HuuPXOHYqYX9Poek1f5MQx0CRxkBw7C
FEqOifhXYMaYEqiCfcWqDMRVeVUDGWSzEz1ONaoGKtMe12Q+HlHDQDfTiu5N8pFo
tH7n7QvNTOf9Wq8lTyBUTcybGIASzzQc5YWzm8ku9BNvbUQ+ndyGnU8PoomXY7aK
pTRmUd2HW+3HIngjZ2xkQoa0z4y8tqQ4t4aacIJE9+eYjR9heNkmj/HGq5SsMKex
+d5YbrAvaFFshLKAkcrKwBgsjzSB/++1Ljq1vbKqMlzU+NfnPls3zphTX9cBc7cU
4RP+oxXlSHOzQG58ei/C97Q9VuDc6qZ+LsPixslipsAMVc04WvpgnDTzt8NHugow
wgXB/nZKgcVPuosG5E0pESihX6QmNoLqIyvtY7DEMk0cuCCq8/CEZE6JDDRUsVJr
oguMhsz8nZQlOG/iro33PrpqvQP95xXPQgyUDqClm8N7vpYRI8OFFKxx3r0gbw36
2XNcv+CzcHeKLtS+UXwhR2FyxsS+X9bKm5cQfNs1W1e5bWQGVmIdgddl7pll6sgQ
jnl7Nd7t5fayIwnXkDG8b2+qL/VyAXK5HWBBxvFST/qGBNU6glHYbPylYGQlMt34
c9NQ21I6iHF9r0/OEBdR1cHks9DgSE/AUAVhDaaCzZADH2yd/u2NjAs9zqhEAH7K
jSI94PwT3SPMNTFV0/PFUpZSxF1KmsPV4Nw4DPFjzvo6sRX7WQGcy59Zd3IN2rWC
5M/EIHyKOOoDYkJ6MiUK8iH57CUlghKNt5egTTZok59dYh7fiYqmblqfcb4UhbJU
Ncs7r7ZqMrBzLgWtX3WSgHQ7oflU3dqkhRLH3K8RHMrTGZEsYAoeGXNp2NME9mdS
kk9X1dGXWJz/thav0Iz/PbEa8NZarXQRvWaurkBVa4SMMmrAIMtrRT+RQxAiQiYy
3ixAq/uCmyp18orxuZqmy2wJbvzxhx5nRJDsFBoFGzJA6oRU2ryL3RWgbDuU8Rc1
ODsnsQyiWbtUKPnpUgZWs1tiez7yrDybHWPWs8bTvXWusC4Hh16APZvXhKpyc/Xt
DncH0NNgy28EMbKeJOS1ufT26RKcRZ837i+RdqGyswxEvmgre73wdMHl2F3XbAR9
IdyhkB7DtHUO6/Fdi1WGNmH9rSmwbsOj+kpYTCThIOGIVjZDYh1NR1r2pyxC8YYU
UDZ8pvvw/jVHQ0yahqDf3sXQ+lClmsTNCyPZAsyQg3elmyN7lBOWFYq9gp54N4ED
9gp+tHFblRy9iZ/V6lxGoP3V8207w7hwerOo2wce3cjPsQJ4Xda8MeZfZo9wODAg
U0wBud3eSSlxo000cOLM/2lPHSma9Og2N1lvkFxeFv+e079QisZtyS65DSqpUu2B
jAEJxXe9q3Qq/ELW24RNRUW1mrLSAFi/ovXvO5ajpjCgJa/S9gJwLMlkYjatq+I3
ahiw9RbaHZ2aQtuMWeZindsOPZaiP0KfF+6t4waYUhDXaLVK+yR5PCgrqbmoZ4Ry
9H+jYVRxGJQ7alQfSSrc1vsNi6udaksS4oTwOr7Hc3KCb6vQZz9uN3v/zllLrZRa
G79JJY7O/0+wluCJEm6narB5Rcu2Kc6ycD+8eJFIsxmsUHKSOmeGmyd5kDl4KiXL
Crtaz4hgO1EthGmZ+lTq4SxrA/Nu84JIqIaxqNvBRFXwV81IN31fbUVwrSIyXcrY
fTv0IWGjk1jlmsjA4NnRa8IkSlZFWNGgVeiGOHUEZ2PVLua0DQot5Nlmxae1l51l
j0OU3/qmYtOJRVILh52w8OEKK9sZJEIUODbOPDWgxUPDsxCdvZjvA/mKmkkM1XL0
PEO1l5xj7hKLytdASrp02GagCUYQZO7PeFr3yhNoZYknlNZ3xZeAFpmWB75cm6oP
jPX1ntVnMr431NbDJNXg43zGA02xry3V0aAFh/hXu/cHiG/vUMbcPmcaxkKtAbCB
X6eyELkcHza0Zy39Uhpj8sQHls+I47uXc5jNnlZuTMuo1AkiHeJL1KJBY4zkTnaR
PZ3oVbcYXFxvY1AO9/IHy3HLFR5DctyyrQW2SPEXAn6XEDlu3kCoY58r93uHrli8
YR5NEmLBCRLjpL5UWWCSoRIj13HqbDsiSc+4suobezH9oaxkmVtUPEolYAil8gQ0
Cd3seKt3KgQsWsFZsZnHby+/14c0D6xMwim+RgiZxlt9j72rlNBX4+ZSjoQ3DmOF
Y1hcANIFCjWd9ik7O/qIYj43bqP5a+Edfy4PA/gfs7MJb4chBElW42qLSaIqFeFi
Xiq8CL9xK5VOCINpM1d7dAnFEoWujUQXOB1La55AirbavwxKq/BYz3OsDaO+NM4W
OIVvaXztawX96Z+ckStmeZLeYaahZLqJAlR5wOV7OHfc9R5yKHIo1lI9herBpSwa
4xrapfacSXcX2LET865cTCb2cTNCTh7LxubaX0U+6+B8tV8kfGi4QMaxRn4DiLJ4
Oq+AQAleAn8kp1hNphyo5gw91RJXpw4w2HrgAP3bMN7/5pPah+nL3G1+rY2XpZ6M
gRtLy4KOGa6nOWsdVdfnt4YSlG2vW6ozDCIHzCicvoSwM3xSAFI1ieBpwfagERWb
mHe69RoMRrckV63GMogmd5zhS03dcefb2hUPLVrEkJCYhET1q+p0xN63rzxYKbR+
cVOHZ48hBmqHvHuTrsyPexke5UYZP0OlEaHgCnynDGGf0y7UnNHZoiQYSJIh/sRu
8znB5MSeQuXg4tVyLm8I88OBVccZ0I8dDuXA9e97zHK2Q9ColXTa9p4oXSuGfbmd
WRwcT5lf+pAcxbn2Nj6/lDXevaNly39aGts9i+rkGI7UkdSQlk4vx9GrfaUkhAjE
l6YzZ7tgVWEGvNpj5pW1XuxsL945s8WbjtLpOLxIFzAJY60jF2cyb3gS4I88W2WH
70dc7F9PhHSyatAA5TjphqJH0dutzaP5nRiDWvSXXv88qntp/h7JaQpAWiBrNBzg
9Ga9zGruuzCW22LNp/r9Z0Kohh7kGqknaMN/UYGhiJMkwXrkcDS+1ebSp33S0Yew
Qc9ysmR36ZbgUy7YzaWyLJhm/PSpK3AGRt/nk8xX6XQLs0v4BXX4ltE7orqF7VZk
8CbqFwXvk1vwhzbgzSofdqLhzhCqUQqlA5KsdUVTvlvHyLP7a2XTuvhsuNAgKolg
+jZlLAA0zJyPf/ruSMwVIKMPPe+MS3Omgqf2A532YzGqFoOcF0sJP4F2jc+ktj0f
U5JbxIFh8ky8ahiioAxTyvKrWuXjpuY2MKe+vYMfAZj90kOx0fQD0lxAzaLqF6lh
zeUTyrdOVhxiYfV5Q1LohNrG2hdED3NggmAiV2OHBrFPwC93E8YwcxHStSdtWHT3
YDDupBj3476ILdmY0+YdcV/QRo7wWl62CWBGwdestbdcKWhS3THzlX+STFHg9Z7J
se9Cx1nVctAqb7o5W8v+G0GB9qyw+kIQMBTzNHPSa13Mt/qVX8VwzxhiOhj+VXkd
KN5rBkgYHG6IResIXmcsSEhcFqVMXeU1jW8dF7iIursF3dbYebiZcuiOb+6DF6zZ
BS58TRQ1/240nH/f+2JRaIIozTA8uOhvcSYcvJDqBl30dRWMQK5+bHvJeFx9bQH2
V0jyfep4H6mVDDMcb7c8KBCu0FX8kOndfi7zx32/F9npWIVSe8vz1o7gm7L6ge0b
aqYMPOZncLKxdRCIDp3FL6pgb+0FwB1u2egis9LHb8Gfba/iISN1kA69IqkntayJ
632ZQ2BHWT1sVOEIvJ6vbr41kCto3W8/Esc1ifpi1r3yY2hEwI9LCtjXvRX1SvhJ
WyNbmjKXXKu89jZmXCNmXxi1HWlK9hZe8bLBQuSUXjV1/Ow/A+MmnUq563ouJU5R
imuUb60TDcbW1+Y0bt82ZzRVkuAuuLXOjYmJYU/Ty4OVshmMedg6maawYoqbuype
wKGTAYzbDSIZM57epOvF3/bGHAGbvjxjLYa2IOFmw3GwXV9y7Pu96qGlMHrc4HYs
aClQip2gU8JWQOUtcIIHpSr+qsm7suXyuaqdAo8WNwRnI2wStK3z8SJZ+UvD+qis
47VXMgXeS8Lo2C8safviWOeHs7O0wq/FTeyCbfSApiA3cp7XwHgt4NUXlInpxaWC
LONAEiA6CpRc2rVd41dRBnb79O2oMxk61XQg/QQV14WzmLtjfR/A6XV7hjbYCbsa
wqcoMjTArns4owNb+ORhGlar+TYP4DeDAGOxx2AqFTphbpr3GQoMXQ5jnblrP0io
0pHlZwMM09i8KbEa9urCPeKcZ95zjmiJp8vbG8qbBTrgSG2cVY+L8Uke502v6RP5
Yogu2kOZe+EhonbFfZQZ/vfqkiWW8SU3Io3i2ELisKmUkYoOi1OpIfl9Z9UyBnz3
kIeUL+mbKAkmygPhsDl//uBTlNax3qbfzTUQCtHs5HZHq3cvYEyrh3NllTOLdk8B
3aPkPThyD95ooqTDxGvtK01mm5H5T6fWJy0FD2FTMEhhvT0fEnxyw01SQMQC45ir
H1ATGt0D67Ho9UDeUxTPk0MNPa8bySR04rsxzBHNLJxLtQIXwbk2MFKT512Ig3EG
0GZCW59UbU8JghMPCOWt5VEudXEZRW/1PlEXSKgaBvu7U/0C1Tm3dSGelbvd66VK
KJJrYUYKHTaoSSnYv+m7QUDJO4z4ndBwyHFpUT5ETMlL2dg1MGx8IMqwEmj/q/15
aZxCP+M6MKd+ySKoOEfExgHeXcFlm5B6mUfqJdHc2Eu3pJz5g+JTfL8sb0jJy+z5
E6RpcRYquaQRfUQoDDprMiuCWdDUWSIidocHsxB+hLNmo6+41XOTbqOp1gNBN2Q3
w5BGM0shqotcf1kgKm2vNFYA6uDWNZrWr7XzvYDVb09lrfVfrijezVNGOF/DuoFj
nl4AbQhNK25FvTnfwKtR/OlqvCTHr8rZLSNJNN1L/dad+3s00JejYyPeqsW9Yv0u
JltNEDVlDm2b7axafthsAx0JYQwtJ/x9yo1WuwaEzuyqpP87c3VHYtQ2IzfY/yeL
DyNRusslU6oK8+w5L07JroGD8gyMmlx7B2lBGOjzG9fay8ZQF8rl1mhfTG2MqRM4
cbBGlPkWokfvcqUXx9cvi+DyB9t5rLkXBPyFoD+s5N1jh6hfB1UFSvistBvhTU8b
YPgw2un8ZKNCRMiC9b1RVzcWk6/qdpfjEC+6c+7toOmo7iyqrutWiWLO6QS9ciDL
1ka/454VJLSxV5LPHoA7zTFE1leSworDo3JwtY40epjML5ICXjSaoMD74qh/XNuH
zqibAFJFFGmxx/ETeLNNPh1fiQvWoYdoHNfZRKVGCIc/fVKHQzATIRTQyX3ojn9v
jS0QkHJeAxr5bmTaYiysunZYKRmL3ZKCeA7tEDCwDIdpiVJlgX7buhJScQq71wuk
Jft+wPfepddceWfDJyezPuvqrmo9MvJMED00WkW+GWol3J0opWYzeb86gxvCkGtk
do51d+1oPgDhwMCyJ4bFxB9PzgIjmmAuR0Dnp1XKJ6KODZJPbQxTiWlo3irfoHBB
xaIEc6aGHGjL7v+5NV+VB5plL8Sa2dDGkutUnAMWP+KiTJIQkFfD9/djS1kPhjgg
biKCtr6crquEqTPGFFCajivEn77UFQdUzaiQ8RCGdTUeQY20aLGuFkoD/amIMrR0
azKEMMQHNAPFY1vsRaOojx/0wMQPBOlrI+QQEhYk0q6z8At4Ux+1MGxLkhDP7I/8
TPjY8xoFcPtr3Wbyt22hsftz3jcyF7IhzyrtySPS7q3BI5fJNRdz+DYEC4RbT/Qc
xzrgcZhWI2ZloceVj+Xk0Xpp1Eer7Wj/4TU3DDKH+DgGg+ZFQlSFFCOBzOQL8Rkd
/5WGEV7EHl/YwsAAy74MPttfMpsIy5Q09omhRU0FusiuxIrsB7JBwehrC8xPvjS8
u3aUtUbL62PpPfmTQiNJ1ZrPGHZIl/4NRZEvFlZNILLZUgErbA01Gn460QDqYiaZ
Jh7Rn/9BSRc7fNnQcjgAexQ4lxn12vgk9DQJGYmTKR9ZC2oTzkTWkV1x7ccAjyj2
UXUrWmN5xXM2JsrFjy/5GonS1SOh7KUnszR4zL7g9rBbpvfhuvwuPXX5ViSmJ3Nt
OOMI047K1jftOAQpOP4FIexk5uFO4yAGf83lW94jjZ30i4YUzD6D+glmxJ8WEEO8
uUIa1SGtB5j6tCoIF3mszx+dVLq6ut8Umx/EBtcC7NxvKwE/h1Il2QL+h+wDAD83
GtLjXeMMngYkL8Q6bCxCqoe3qbELhwfCLgIGWiUQeonnvgUffrQgg1B6n3lhIV+8
gvGznW8sRq0Z6nYVIE72E9IkTyPwTtLrl2LqULdgCpUSxKQa7oHCWsyODAoggq5W
QBPgrLoyrGSis90Zdxkmo0vPZ3LRi3Q9ro8+CfQLDZ+jiv15k1L7JvtcuIQXJbum
+mck9uqqmnZUtY2NsSvvdhrYn7Cl93SHvBGPsTMNQ30l0fskt912njD32j7/gXr6
ZIZZtwwxEaQhk9IAvzqPdtMuceyWyLhWz+0/KY35Yo8dJWiTN+DAe7p+rgOk/V2J
TKlbnJRypk5j0lF34gPcRQMGLL3yFfBZU8R/75+V+yQWgNPp8KqJu/1meSTsZYnX
zdPguAn2AG8oWR9Hzo2diD4u/wQcAvO8B6TyE2N09bffIgQ96imOIsgTHLx0WAms
5LPD9gKrKj1tTcmggp9SIEI0OnKE/AUaDQXoiRvKDy1rqoYjl4Z8VCKDvtau8Tpu
wFVrbeRARuHQPq6ndVv6gvTuKrH6Q7618MMp1eSDZyqtC3ZJ3vaIMm+S+S1T3h7O
+htZMd2eUel64/uGHkpcigRiol1/fmPST+dUHVbBH0it1CYiiaA5cSOEBEps2+HW
WIHp7G7rDhCcodyCcE8o+qdu0yQzDy/L252FRIbMokbNqQqJ0eaw+A1bFbr9BrlC
OqbmkD1gyFwsFIeh82Ah3Y7am7v522hICLoxOMrjEx+NsXpl11rUfHL1IHWsk+TS
SZasmrjiYRzGAoJRhNFxi4rRhcueh3xNGJCPplw4yGhltI9UDaRUuLZBGh0VRuHd
/vRx0s8rzx0BE16JXncLGAx/pYujM0ckh2xi+AVhXGjNXZyWwOutFow9lma4oeem
Qylbq3KIQhA++l7xngYKVOfysndZ5MRbFJ8yea52jzU+Rnp3XcPenph1ukpwCRVk
ammcOvONb/ObU/2YV72bOzuQxCZhplmahe7wAdGCWKrL0O6dilvFnKUeRgF+C1f1
aUG8qPWPAnmlGfiaM1rE8F4kHV99L9XkdsxLNiJZUTmk6NyQakp0+R5iKzYFlu2Y
8iOdJYEaNGwchU50wCOkzhQpByPKJ+KNdYDu6uzxsWNJvo+EdQ+Q/DMKGdSdSNyk
PHRf/U71uwLTYt4oa7VhN0yxfj/TOyq67EA2OVF5YnKMco9UK7WHHuSgZr589qsP
VZQsPXhZNZ0yD3dqv9wQLiuOFCdHb0/0ElnY2twPebTfHl9XDswTJS6bMR0HYVd8
Mh7XnhM7nQRJPXEoi09LH27WaZFDePnHyRc66kXPO/pUA2cVkBb3tYW4qyOAvm/3
faa7v8y6PmaQ2uQJWitBtwohSZ2LhZ3ZNdF3dRk/YgBSG3GD6C/XKMOOEabxY1NN
QA+BFdzekD6+02wlgbhcasaopOtYSJzSWVcedmYp3Sx9Bctpa/eV+btOTHs72Uy2
cmWtATYK5P2bmV8Hf67YkXHdEpFgAU/figHNnuAeRiCCeIQc4PUQ9kZN6fmAPGur
q9YkojFizAJuMnZad8dQPB8xdrSLZMeL8hmB6H7scQy8j/h165HFeYW5dkb6e8BT
e2U4xiCvtkTJFaaglgwv7sQgSzfODWC8+LTk4+Q1MqmGiObDJqVhJk4tuvCwtFfk
FXm6spGjZcJWU5QjIylh6+VuhZ4fAvChrINaNpeOz+XqgezZVjTTgNYEjcS1qKsj
2AyurI1QWoCtUfQu95tSFOEePyzAc5mTpbL/ADvyqdmFJVjVXivMMzLnw2OU7aG5
QUqz6EBi6jUbNf+8CgYx1ZhjdcIWiF4rcLWy8Ve7EFyYz6qsEFKAvS5PoYdpaBg0
9dY5P0GBYkHK7k6UScdpLwfYrl36jJtjvWQzJDc8PyHXxQM9YB9r6yKUhaLj5FE/
HUazeugXCBBwiQ/c94S5wnEl37YAFzz5sa1baqI0kp+lPwj1vbeRHljqMQ8BZNWJ
ZmV+i9ARychy2UYBPgvimSTrCTyGQIHPqpNDwu1E4w1i4BWs36NEtuiw4qHdc2KQ
g5ETsPAqey6MdPvVFji7yBqCcDWpZzzFFoSMsxpqZ2EKUY07JlhkPaiBh2Mjf8SR
4hfwQX2fWEjn1oclFyvVh8rMoSC6xt88IjhW8axF+47O9bWeavEJJEqPpGZrMhv3
BdFlxjSM0GShTQiD6XtqCks5B/IAFL/68AxqU8YlJUl/Iy+/18NOSD6SEF1NPUrv
6u+eLWQWMEd7l5+Pehv7In5ffjWmzaxIJV864Dlp5v8hp6CaMTRCtc1g9juFfnva
NIMHWLcpiMdQEmtKCMKn6itqrqGbGIBSpjU5vOYdTEKy2DR4gtyTqGnVxXxZrxSC
RWXtQGJvYJ+nfJfw16Bw/i1s5bSIP/oKQdvZ5Ix598a8bYW0thvNR//rnAl4KNOQ
V1LSazyb9CCeDqeUhwQVMaHwLk1lPaZfTPP5NT70REUjr0wOBQWgQQamDTiVkBIe
e4OxGh4wxKo6Q8kwsDr0grIuq1PnHIpe39ivif1q//VIN1L1BEvNOmzFddG0aOYJ
CDs1V1O9ahLWNcHKwmM/EV8DwwsVr3P3p9CeoDRis8JpyZfY5KF+gh/BrTAvwoxn
iLru8NrJjDnV/3W68a6i/7gI/IWRoYih0JAIg5qFBQ9rKeFiR7NwVMJk9Rm2uPHx
HTZ09EkFgPlC9LjvJFPxFHQ/cju8DFm8H5+QWMxERpILk2JrsxZUvNJv+wm/9MI/
j3Ci/LWJhWlcisCZKBeMCPu9PM+fyhfMdndn5oHFVhQ6jqYo3npkxstgPoNBIsMc
laPpub6EMALBIKYDhrcR39tzMYt3RnTCWdcw8tSAdhdFj6osejRoEI3fT7G9kR6I
Oa+uQEQvSOlSgmhW+X8SOr/Jv8nuKYXTCoRCwYWyhMeHrCs4xRtaOhnqfefxmtyR
MH3SBTsRLB0Vgc+V5jb/o7hiXgpNzBPJ44H63laSn68zsy9aDKpdzPff/uuqVzlg
do1pTW5m3lGfekzsmy/xw2o4ScTSPxvB0slS9/pdqbS+W8RKlclLKBjDEPk19bwg
H/M/0cD95wzckxlZoXOWcbC/KNycUCnA4Us7yJRsXqgjSGs0e3gmM7i9z5OuI6n2
BIy57ObONkz2MZNEgRgf112KT/HfhhSYqOjf0fbrQN50Nh563BN60VqxjxzHSC0G
c2FxI/VgbsATqHcYz//RDJ42Dwjzx+4bi9FOwm0DW+M+5t+H86PUR9HJ6RsIU54l
WRoVF92zrF7ptSMp/28qnyIfmzv4gkbt8c7L/uX61dBBA6hU7XjT1WkNU+F4to1R
3tQhQTyCr2vNNGQmqEj7oPqK0cW6F8prRAJvS+Wb6FZmhcDEiSkO7i8sQ+0Q3Zx4
BSsPCcaL8JZQ9agOTflMc87WfoC26J6WVlQyP5yqxzi5lWh5XHrDOixeouTNck0m
+aLLm67o5gUBU9SS5Omuoy+XbCGfQgotnQmXfw9deCRFp4B42H6LljZzBSRPds/M
FXJswaM7V0/J1AhN84vfV87nWz1L8iLysmVz5pYjK9F/4CQ7LFveHVlSLYky4s7q
7h9DM8GkymVcSf3hbJozWyktL8Ti0XP7q0GOEI4wObHRkpit+zZs/5Otpz0ZiMbw
8tco/AgcSs03wKLt1KMQldvGMBj+aCW2egXH6cBG7l85T7opJoVxG3qePIxOhOzQ
mQdjbM/KK/PaBq1EO05oUrCs4rUalqPfWoqA8iFVO0AWp7FcQ+LHBTAgTIv/pN1W
6qGrTeE0ov1OkdZaWAYIq1TQbFXlbHGjSU4kl9orLWB3ZWYCsObbHpG10VLJW8/M
M867BKlOuZqaP0KtGefx/3EJyOZoTtppHSJs7gcYfYBzF0pv39+DFAn3EKwSwEHH
rfS7m1RMfCGp2G5/a7C7EOyWxGeWk6aXcIn6PmKBded+K62U37OrvZeqKl/Eg7JV
wJbr9gHrcOTT8SNOTNCfDn6cD021grL384j8PRPA/m2mnHTciHjmV4AEQbAWJ4Ps
fsX1j/PTnGC/jTQhRHHTKQ7rx91AqRdAEf7LbbyAG0BCelBh6VGFpVUn3izPOUZg
cwgC5q4A5UWGhPeoGhGFN++Ngm1dq9tP7UyfJyGijyeF3ll45MHYa2Lma/mhAm3D
3oud0Y/VN4cl7rCcQt9g54hTayJDqqGtLgC3U923CD9fE5yCO5C3n1TybDFtx5HK
Zy/vsDB/j8gdTYNgNJp0FXCZrXQhRblHpPKPR2ihyXhRZM6w3qwKAhBFOZWbZ2Sm
n5/yt5ZBITlrfMyp0UKoUGWiwSB/eih+vlGKuQovFm/G4gXsu9dOWwmiXnXUpGlx
h7wY3tFQEfmRl41F6S6b5I/XfuP+7wh1lqSvISITgXovaXjvmykseTt+vY/BLlyi
FaxIUKtgqTq5wVn+2l6rVq4HUbDeyOrADWoP6pdHtcJobLZ9bLMBAQoNRXoZJAuI
8OJ1yBkXs/nHOsC/j4CVuGYpSfIMggoUCHOo3F2lUK2/IFiXv8NGTvhml5vs4G9q
vxSiza7EUq+L5oqCrC6qsozuY3iGFqii2xM9jjvPkR1cbEI/ZcuN3KVIOyiB/exy
c0e7Bq4fQVzr/9+id/iaW+VP6l0FJWxDKi37Ogo/lbJagU3UJfPM/WuWmfvOr53a
ODb7WqbwJBHoNZ7u/WzK7M5ebBntsV5hk3zzrbqqBRlAXQ4aBwH4ypKZwuJBLEHT
Mj3ilgztNbulOJLU8mOjyLL2hOHNQuH7Ew67FYNrk+NkBNxGgMcTzxXZ+djlHr5I
WvGlsNz3XsOnYmtwrUUBAK2JT1NpcyAuotnwCyIylu2L9+ef+UnMWdKYCcZVIN+Y
ysMC9fEA/AjNiYk7t3o/3qYiCtOrg+2u2pSdYAqvacOxpK/jnp3M7HJi/gODnb4z
q9vOXBLdi+k2KdljpCdcoDfJgFA4aeJ3Kfttwfi5pGE8MLnpMQSLVpg9hZlNXcxT
zkH4SQaub4ruaeMwOPr3CPJMfSu33Gq5sqSSUx8GxrGtqkig8ChZ0mU6HXTF48Gc
ZAp088sasAarzyo71ol6IiOQInqumY7Y4IMWSCKd4XayLjaxhtdAlh4NomEEJ3K7
aY0JNewhyloU4YacX22xCM3yg+Ob/0xx2e2eLtUk0b3QCI5Iz+iUEstNToWqTw1o
8AU0PSeWSRYpcYpo+02W/tlCgIaDGdFosAkI2c/S/R9S0UXLSA3Nc8zn9eNj3EnD
JoUnUQ1FjXrEb/FWkjgie+Ntjfup0Oazw6FUmEdsSsB3KhGSGO5nT6hGTakTvgER
GQz408+i50h0Lt/t2V0rsv+Lu4xhX8HXe1YewPS0IXeGveDvnSdMV1UOze5vsOm1
4PkfPJXOwlJy2xwy3jtwTSzTwz5pv62zyfKBfoYXW6W6+eeLyHPwx355zaOVtbGs
1lkBYNy9Ff5D9i+61XKJjvls3YGI3bfQd6jmnfwAUYfUTV+QzkVYJld70bJ7LHBX
T/WhlksA0IyP+to2xgGGikkKLKccxSjRg/0wvGzBZqFgkgJd3vuZpBc6TILt/JpY
HLo66Ho+VwqN6/9DQviDVyzJLltgKxt9eFnKqeapO/cfflrBC5zZwU6Zs5GTV9jR
Qt6JAvxFB9Dn6lvGy7/EgsZrLliOEvmJCew6yYpxBTnGnIzBOfngopLqSnfjHFkm
1maKx5tuq1elKzuhEPcrE+Rf+cIKIV1WiUKLhenM9y/F4l8VtIhJASBToURPz2+f
ootm+qt90yOaAbzXREAZYyGoxqd7FZMjUMqDuPe8hT9KVcZ26uKZwgTFoEb7eDZv
/prVhRvDhoBZ8tqk+in0D7QzXtH3poIXx3IQKvM7UCy3N7ZZJj2N36NjFyWWfdEE
s3TAll0I3yc2e678b/TwKXlX4Nyh3jE8eI1+rSZBWNGuJ5uWILWAYCCAKTsRzq3/
YW1+N6voZ0NGFrQIUxfdV59+C4vqOqSXvPZSnXJDlsaeXW3kHJHJkZafSiQvQJyV
TJ3G8S7MiqCIF30yUB1AVyWc+erp6b/Aot2QGFifv8bh5Dv2ojtXq53DtJwyuROC
NNVxRfimOqwrDlmqNTMR+ehU4hb9YnAPbqkpFsEVZu5P1x3R7DWvHr6ItqGVZ5ow
lqVxVEKVNxzLZLWPdkaFFvgZcnQhJEJelKvFqAut1HmQ2FfmnMlaDlmJb00pNVrk
OpbesogcRwVcdix8fR4GEbVmHkrWniN2D7YH7KCqxe8/CY1R5vMVjl8pxSQMHT/Z
EzS/d1OyTdqzp9ZFz8qjrWtiCwottuzDdL6379STX0K14xcw+pa96tFmtPsp/LDZ
pNaaeaC5HVwEouPCvaPkbpL73TW4O7x6exbfZ3sAXDiBC27bMYIeFqJd45d2NSDI
aVabCTLWOerrnU645WcwIUhtkBdJmvWr8/BmVgtUyLt/MMTQVeNQtjQhPqm1SNLS
XOKEc/Y0MTF/59OlHlBAPasSJBwAqgUsyCLIDOmUhX3iRL5gRFv/L1mtoUBXqg1q
LSzFqBwo8fLIhe7ya7kBgjtVf81ZItBk84bxi4NpEwMFvBgbI8QP4kVIIhcsONeE
vFIxgFS6KT0zvnuDZ57qgtcCK+hIN78ReIty3apySTy3cncNbmxZpMj8bc1+RJSm
ZZxZAfswGEMfGGZEfv2Djr4pDmfejlpyXdVDOzkh8slG1lBjhzW7RPUpI2WuwLoN
S/1Vfm3I46tG2nTRxtyPqFhjllgpA0n1qIvDaJLt6shQ13ht2t/ZFnCAQG40TFKv
5liE4K0ustCvO4JXoKznjmkTP9znXIrpyMiKgUI6h3R91zMATi2sE022vu0MzWql
z53p8cEmjruDjL6hueu/ZZgNcTZ8nrjWRzyzUetnlF4NUFITrd9EtcvMqiN7oPX1
ve+B0kEBE9Iub8+JyI07uSFs51i7LYOfEK+W76AeE7zLlA9VcYwZDhv6ncF6VUQh
o1HhXfrkHbtSKhQp4qqvlV5f0oOj5B5VHi/OwvtJ+OJ8EAct4C8MB7URrFTeAZCF
y/e4/2Q4WKW5goph5UjVaygnePIoM/j1Nf61F3iy6K3oyjyEOwUzD5pqa+79ji2C
W0BjflgsT28SOCDN+s5F8mj1uY56h9cIa4foM/mgyri19HU5GP8anYmfcNv/PI71
xuDgCBGtV8PWiivQfAT140RnE019G5NBnFIObmkqrOfUNpAT83u/fkrUmBU0nFLp
BmJyzp8aVZ4xuLvL8YoFPgfhTSxMobZPmD2Mx8jjoYvey8qxpKF68CV00O6NOFB2
hKq7PHjyr67trkPp4o8GbonZWWFkoJeNyWRarNwwMdkwEhAGH8TzG/FtgU1GP5UT
IxcSg0pD5Ejt6mm5vo18SpNmkElm/1gmGEjPF4c4kEellecWqxFqJrtLjGgESCAA
VibSRaa2255PEsZ9UYXj16hSHvJkfWl7z86gpyazvdZkhcO4NWruE5jqVwrIPIbR
ZepOEX0+FtBBXka7VK3qhReBoW+74iWwZV49bX0j5Isyqy+CXd6P5mneQRS5VWno
54ZlzgKmnnrvB20IF5PvjC3GyKozdN0bw1jaLSbxBXw0IV2z4TL0LU3YrIXW1Vu0
tARXOhqSGRWREcGcbYgSAVJxRVMbbLlcdEx4l0nLjZxctRv1oLeKhDV6flIVZFGH
0h2gTtJPsWuxpJwAg51R7FL89VLTqTm09Y/HgBHAJTXJh2fhLA8lroM4WUGJHduf
nNwLW0RMSa/JO0jttCz5u60dkB08CqsJL00hloJko5C/AWnFHuBbRO2wS0RvWKwE
fgZifdGnLbfk7IDVFXWoVl5kUG+yoiEXBjuYAHgJ+ZCQSg6+tnuKvCoG5FXm2zTD
KnRMLe6RhOtVnbPo1hxMpgdPZ7ctuKqCzB3AQmYnKEJUR3GbL5yfolaYreKGss2C
4psSec7Zut4t+hLT7sUIl7xUqHktgx8wCvGUUJk9b2rIreVZMYYnQYfJ+sLLfF8M
48XbmfLy4RJIl74mYTyR0uNjBZ123rHOSqdo75vXoIdCHlj7Wyzvo4Fb+ajJcKM+
Y9Q3i7bifyMPWJTrzKMgBV3wMIoRaiYrRmE/DoBBk0zAUs4MbNmBxhQdhY1lB3QA
kUaA2KlIXvQa5Vp6UxhglWtrGeJ45e0q5ghfdRO/GNuk+P3oSKEpbM2hBfqimKnh
5vY+FLv/yZObOaD10AnduUh35f0AMdKjFOfasyCnq5ERB2NJQS+7p+b7LVZwfQIO
0s9Xbdg6wdQ03hXVhs58LIWcbZP71dShNbqUKcF8SEzGDC6MPhs5mMlLw9+zhPTi
rgPFAbQ189pw+ACybiiX6jkeYz59pSbW7XIFwR+3WhBnF2Ve/LniVUdImptExQNh
COzp/d45KxxULNNkU9ZKe0sI07akj8EmViwqFtTNYw9joHUtMVPh2qduTahUcbHJ
D2RydLvzT6QP6MqlSt7hv39AsCcd/rjC3/z6o6YOuolgwKvYoqDK2pkZ1kKHc5nR
O8gZ2w7STSHGTubxLbNYv8G3e4W6Rh97pb6/ogT7niWDmJ6kIxltQYeImLHJQjtM
vbGIMa0eFEyMVf5Dfl6CzyiK7ewU5CYXlz5JhCQU1REqiQ0n1J7yPUQKqfFVSIji
VyaAqcbXHkqFs3vCchy0jMkd/c3SkVLtGmCrpzIFG8Be8wI3/ddV+Vy3mpr4Jvfp
/kraik8vHF3Ehl5Od1JvgNHfZ1FFVVVReryNoGSqzdIYA1s0w0AZc8UTkLx5ibFz
XELFdJH8HjYl8rpQQ/RzdJxvdwtTCtOXEzg1Br9Sd+dcIbSrl/CVM8a3mDM/WRQL
e9OpXkwYWywboTKO65GPhqLesb2kSGsMvFH9sFJUco0jVKbaCpirc2nOS7ajAwqB
tGzWhkQrWn0ehlnxh00rUm5GvwUQ8JfD5R0YmjXgpWmnKOlgLZtNncG7T95U4rCL
+RMqalQyv2/h5XX8APeaxETjOMFWSpkss0uqVwBCVYvK8mUcZwWOzTbsCpH27qht
Dks0lFyAJGm3jVOVpsQRcyDE37TktN1bc0/lSzaSgTUqrm9CL8jva+jCERtXnjlx
9W1sPbRnK21IlyXDvTJChQZL5eQrMI6grTEiudPQHW3X3JBmslCcE8Gp+ArRuGIV
aUhelqGuwbcGvzMc6OazEMImy+Cu9nE8dvlhp8iDqE03TZ/JQGaSeB/kvV/Ezbmd
Yghb3LrrwsaEfUe/v8LsiJsJVM21dmlabUmaI4oqgGbxSv325WI93a2IVVmSe2cA
wldvOWifYHIhDUqqGEtsAxmq9mTHGbfwA/EhmcaWXJq9hliaAm9/dU4Nl0IQa4Ui
+ggLcm8yQOi4eILLhJdxYz0YCgS/BL+HORbn/IWV0UqhO9NqeHsbPDmXhVcZQZ2N
r7BFQw8sIIYAFLfz5rMuqwdPUUBa1Cfig+ITGSXDUaZ0M6AWSOb5AxbJMJKgk1lM
NawiiHOK9JLbR/0K7i+EYkoZ0rn43RBlq64+MKQJD+XPtOmIYoTM6T9EjhWii9z4
dn2UaucSCbcRv8NCkILaW7OHINBWdII73EHpPkV3Z8ZQm2P0f4ZHFrEZErkPjOrR
1l91J7TlcevrqhR9P18lTSg2+fs5oLwhieUgGWySPCuXX9M9Ua1yqxD/Wz17AHuN
4uanXFcyvONbJZbEoTGN6SVPPLoEij0jtTJarIDY0L11jZ37FvOMpMuma3aT17rC
8IpHXs3lEHh1mIY1G3SkfdTj/LEkBOgZ1VyZZnvw0wxF4jz0Secnn+n+U+/aWyi7
tf9i8tg5Du2/b6c+sd7SnOsZeKcOUF70++2tQgpKumdztZnr07phw+8pLqq36wrQ
bRgItrV/4GZdAZdVjpSVRF55xWL06PWXNVxHJ7dRJuEyO2a3EUNo+rlU+ZOfb4VI
P5FQHBkiztTZJ7+VALOInBK69zSEa5m2Ms9UF4avYjXD90QNM0UZW7vqmCkw58uh
nZTJRugqxs/EL8abe8b1+5pRvRAQ4A+Xl43vZnB2J/eYdKqcbh+KIFBqzSkGyye6
wvJWbGCsdBvkCczqviEoCe4eTZojHSThJQlCOGqcecnE99/hD7F05kCCeoifGDPP
SBzEVFzwKrY0DHqUAGM+fkAzF6fxZO3cEtNEfKWumDaozeKBHPT+CxYZ7QJ0QLoC
k8ls7vU1k9KvoyO6nqfJ+DI9FqrLSqbzYz7WJcP20cv+qvmqS5E+hs/+JF7uB1fm
eIXFyjRD/DVIh8BZ5VaoHna/x2HgMoKMOyNlRgXWgpdU4NyFrkaeExRgdRc4Gk1B
zR/qmSRsaRHRwIxuwwfEn9qkHkBeokg0NeMS53dVFOArDcEY7XGFmoC5jkXEmzux
3ewJ9duk+yyKXcqJO5WU1Ddel4J7ykRVK7I55Jwommd7Z/61OKtLc4zH0wMLkMNO
ImynkIDEuziJkJvSVDIUMr8MLvnE5a2BDh9AJB8ZY7SsihX8BLFM+1TiFrfhL9Pj
hLIrvJzypmV04UPD+fmlaVuCpYlviIyPI2HH3gwTSUJs30nW1SMQ3zAn7Q5/P6rR
d3bxWGY++FMjOPnir2+IAaOYwZ4WP6GZV030Guz2WqkTmSQIv20wnGz8az5mhgTJ
vNOnfe0ntg/QhdMIzbF0Z8vJsJT0RcNrCHYlZx24q/jL1syofN4URfZK2jMLtuq1
U1GyAtkfb3/cSqHip51fjkk6WDHL1cEilKHNsfphnQ82UA2lOAKACFpMIRJDwjij
eYspEheqdfEWhly/WfzOmawWnnEnrOzDZLz3TlMCYy56W0A1zQj75jiO4mo5Zn/t
nOblGKm31v2HCsjrOAbG8aEwlD+vMskaKbz5NCTk3nqrc5kOrU4q/0xMMgRdHyD+
OeRle6vMfT1dNgnZFEEfo+V2LZU3Cd2jAEHpdR0vMUvyHZObQWb1C4ZnrVgNdrkG
7hS79o6uQ9AYHuKUrnYwApYBlIhFa4Rj8abjguvT14ckp8+qz0xBeiFZTeWagD6g
TItgcKSCh4pazNLKGQeN5gs1QxyQeWr/IQtNJ9B7xkz/Hup3pbsA/IfZAqv3GGmX
yfJL3ZN1UkYKVDQIGyOJK3oH8O9aEzk5NI6ro1nD3+58c3ECOrZCa7zwVxT7led8
vjaLv49ktYKU/zN0E2Pw8/zjJwV1/Zt8yp18+25P4Ktv1qM2TBFhZBfHH7WZvCEE
UnkV2mZCvlfpKf7j//LhsS3Vp3+6R60tb5Y3sIWorfbFc/7DNa4GyGmw2aeC6ALi
PWAbyXHa50PjCSHXddbC27KMOeEb53gdVm3jBkl5mPC7rjbVejx7Ln6G6mZfDALD
3ouxergzNHbNtm/cDJgp7QMmY6s1NYh/xp5CJiUDwchGHRLNti64fdsR3c0sM6aH
ok5r/pgM/GloxKINfnUQdFTyPUC+mrsgQZfgx6GZREQihGNZ6HrHNZ1x/EUbS4SE
ETrpT1EleR7m0YcwDnWam/sSn6+fSRrbQN/VK2QWVoQyecpY/miYN/o6KUsEel2V
cTI4SCMSdPDZksdVwOlmSIa8a/zPqm6wQtTJTFHILW/O7of0oUmU9Y7UII9j7kc6
EhRY21puTGiA9ODgH18AV1sOBn26keuzVbb3rkuoI9YSHvPUCyTrkrLjQ6XupzgI
WfF4bL1RS1wdpEh9nH71TAHEsBJHjSXAbWvxY8RtgkIFNFcUeg/4nnRKUIdyCJg+
PweEu13cCI/Uwr0T08guF+Negvp8RWyYNWX6ZAPLH1qhShzrM24ibGBCi358XY+f
PvXkODVMF9QTcnHWkW2wrkax8fRCkKH3RVpmAc9DmDfz0M7SZEZfnjqfCjTphsND
pDD46vQ5tzpgcYSkQWM8u4xbRbee2iw5aeDQr/jo2oUKWs3wiwPC2xcNxryCIHkE
cJWREYOSkKAkdH+Ueuf7rrdgRCWayBZb6vOg5zgnFL2xX5m+XTCJe+bKClsy+Zu0
CgIPQvpuk2L1zgZVlLnOg5657diJnX8/bEOl/HMNndjPMZcyz1muzRK/L7MAzth4
6qI+KXog0jAiCD9aySGBesyI9pjqKQfyn++lqWV3gQkvCPG7dxZzlWGd2QcOnHIh
HmFjuU1KNEpxS/MmbrPlhBBdPRX6MnL3OfKKLjDYCPe38QWHarZQM7VEW4iSa0Pp
cAvwZ/w3xbP8tOr3uk4Q+6zs4H9O7MUHHfD1q5DKBWJEbxKsFhKn0+XA62+ZYavl
ggYBd3QNb5bUdM/Nm+fzSAt0fCJj1WHPAIAv5iSHpWn4glbPtoe8rVD1StZ7bN3I
TG7g8m6TMW7c7GODPM8CUO5S3flsx+eP+yuR2Np9A/EpLehvlJwZeCC34RxPHJLc
rYdy58rdJw3vy5YOrCdH5omky5Btf/82B6vPouewWYh9Fl3T1qo6wEwOGFy585id
zB2TY1/6DdtK5Dmf9XCA52BtfNJN2KkFxWyJD42LlC80LTOiNQl9fmZgU1Bx/+Dz
qMcL9PgBMZvscmDMcsLWF3kxZLS4IP7htX/6oz9KpuRnaIVvZkWlACzOKvRuHPdq
tYv6zxQUFJjQnjZx5g1uQeWTF56v9SnzAM1nlzfNJAkz68zdG+Rezm9wa0RDRV1E
MxtCXSVwwPArY4ZcpgAcYsT/SGuEDZ2oBaKaiz9uIgFxBxLvz0NQyTszPvxn9XDA
SRsEYoOVheooLxr8ljkdpLFsDKQq5Z/qF5BAZczppJZCnElLA+FSNshrsH80nXDU
TIOez9I46wOj/6JWNHOc2ooEWkI5apJ6/RUIRvowZv/sBUFtqaPt8TieD++vjnws
wZpl96qtIZVC5RsltAGtA74luVaniN9UIYXYtX/ODiug7PVuGz7bs369Cb0fqAWG
E2g/vWTNenYsX8tQbKtuUoUVcaN0u6s8AcLDc/TrccB01qN8nOVIpkVRay5rv3nX
+kYsmquqIEcwB7ohfchLPWWvNABeqG0kHPC+8h7sRM0LJJUSKxdhBYuhSmphAhvY
7xyXC3NmgpWnmasdpJpKjYBZXuKm2gveCBu19aUa7RZQuCVm9A2+lZvvCBQQiZQ9
yaLXIkes22m1bRdanZQfoP9zk7WV4g0SboaN8G07oEFM++3HwdxaeEdwihCjbREw
WUlFvzL+V4LjP9BWyIJ3Rhjvm4dbSzhGtLHKDeVdaHobupX9u3uVKg9g6Ks6v3Dt
zW8b3nDmdhZNv4z+FVK0wyk243xq9lY9M4fNtZf1QNHT02l9bV+/ImQjnbX4Uv8f
iUWCn/42twcTh082CbxuLTkTUloMwtE14LjIqA5do69sIrhlHu/DMN4RyLGEJa1O
9wgCo/Sg6svYDMPvTXGE3CuEsGcocFYsNZdSA21W7eQddoZrJDMsIdc+IHjyffdF
0kEwRR3wtfSfTBFq2yBwW222DZw1UMOjP2JxvM4UCmwH8xaG5dO3O4gfa07Ww5yt
o6XDI3m0sc2UOTg4b78PqUH/jGpJ6LPtsPBNPoAKltzyCZoPwNttg4zngRR0NSBe
LaWuoXUg+skxLlvTbhZbHLxbhjXGy6MzDf6gy+cZvNUGxeKAhry1VsaJs3irBFNs
LSAf9CLoIPVyN4VfiWfbU1sYUsPg3YQFPM47g3OnCHJuw7tbN/phGGREJuNme8TP
CTsiOVlZ/n9iiUmGAbQT4l2tSnbaHTITVlpdQQgEmZb/LT1EfZ/JHLt3phf+aVTe
KKbQ7hE9RX96UlnOLSrwqWqYtkmzDEGpu5WO4JzmCQ44gfjQ0OzMLLuN/9lQ16NK
SHxe38tGmgZmLUhnKB3qDbHX+2AfEhKNBsFZQg1VjlK0kNsTB7XDdJoIPT38OXQL
AoYerCRSwbpfRenyOkeMcDNL8nNHB8QChmfPquu9oW/C8AsG4UpcHGu5zBi+Qb7f
e3TfbwkgiDyvv6E3f207nJoVjpo1+OzOj92eCWq45bE3h4CdGak70uXs3gWudE6U
QwHhZYKevA4CcIdC/IRNiRgvn4Oc6YKatQZHWOKl/dvYUQMqVijlQIdE2kXrOyqC
UUOt6Uqbv5JWhxJ4q3wKWKs4HRZEg/Odsam46B1kM2jNWne3y06UFaRIs8mhIV42
d6ihQuBlVraF+CerJXn7K4AbEeOU7dC/7IHW7aFzY84MqYvOWSYcQwVz1x+GTZ6k
FnTsJpF6LCNxfdUHLx/EIwL6IIHvouGO6kjuDeKr578kobxRAN0gfW8kK0lTwe5y
NrbNG31ZPRUdPJ711w1DTudyeTZDBZrPdMc/vzRofZoyBxBgxKT273DFXc+bLVR0
xjYqh22bG1SwrsPLwYH+IzRhvBS68v67z5dn0z2OHJ18VjKAIcrkn6PazrD+9ucT
dYNWU3vqJK+GWv4+qnrkN3e1h71MK5QS3VcQdSIcYSnWf2ZwSeLHhnec5O6ZJvx7
g3R2qoR7tr4fEXE/cLvEpBbYKhEA7PP2wMEgvZCvvBcdIvpru6iGDkEtzQi9BBy4
kYXKk8lKtUde4H1y/swPBDp+62ppMycTpTXt0SgoDN8D2bFfvZbGCzLSRzkU0n0L
2n/4Z9qjchbUOETDSGe3aogBdV6KKi9QtRWEfzts/LVi8dswSz9jU5cYDyAGM4si
/nTlbkaOd0qqmDqrKImTVjeKPDR8P4gqGvKzRqkZU57prB8LdNXHcn3w7esunAyx
Apm1gmCV9rfSPQ1F4puuIZrMAWuvTjCunQ13q785vYHGQrQZYshtW91pmbOfyX7c
//3WrVzW3p1RS3zoc5Rq4UB+TfOycANYr3LxSFojnl75IMUeRxqEhT39eRunLAPZ
lCBc2T2xEiBVYRi5VKeOlt8YY8udiDUCxvTS8Xf8Xpd5ll1T0ebZDDqZoZrjj+Y5
By9DMNwcvV3c3qtT+Y4kjMWR8/Szz50Ys0OS/gnDEDA/FzgVLeTTB+smaEMyleRH
zSegRjYlbpHruXiBiNqBhcyBSnxZF3tMOzON1J1acIbzIcZSrSUQvb8bB8mbkriv
5ly3FxoP6FhCkqVLaoYsazpUY4C3csI6nIWjyT/I+Dty+FjvHGyucSuwr4Q1lfAd
OfaSQkGk2JrzvraowqtGPwGCfLKUjQcYDmNFfFm2w7aTnhe2Z3bRHRDau86YdjHU
JKgfP4Q3lJ5optSXQnAKyrTJzhS2PIbz7ZW/tZkz7nMwh8SScdJXG/KObVASQkum
tKHP0rK0/Aj+jf/3wZazsEhV3bcKli9F2XU5HmzezNYZnn9EjlvKAUYSb/4/ReFy
tdbq4I5Ux5S0Q5ibpKxHiSM2V8BmmeJozL+zugM2BZaM4o/N0khxxr1rJTGoYpoC
WdaGkUwrE5kCRJTncvA+l5QRAScfBptmqi0Y7i6zc2gmMxarSMtze2kKN9Sfcs/s
CXHEL9ycx5YaQzfWnL37LGKg0wgDb7jobBk216jDPk26GzO1CKaAoNBiTx9P2BMc
VmJ0uDf4RskIS1OwbwiORTZYH2QB+74HFWd4P4+scUbzlhV06XNjjGO+PWGbQAnH
OUoXp0ZQ80b5DO0XRJwORgreyWMrNb9RYI9jhqvZW46jOQ28sPzMhx0n5RC5NJRG
5DrLxIZX5RasKLoLIaAoFvzTIjqINdlnPhM1wXC0dHn5ANJYlo6wPHQbKUfA0qNk
r9CqLi1YcED6gr+GZ91DBOws5y+rIKqYxLYqePjMlqtiZR8TtD1FBSmCKnz+IPO6
9ETNyRlCx5ib+h6og23QgcmDIdIRo64o6BgT8C5uKMARiOXjqzlkoqBWNSumRdBg
0ZRCQHrsaqzPXSU0HdQ5xNk+3FKssol/n4lbbfOxxfZqVaZDYhEh/Q9owM8WdxZB
X4sPiX70/L7PtC3M6mv1a2K1vCd3MYFvv3balXzpp8WzkBt/VIc99fx6unoEa2Af
Pbe2NFN9uX7tonsBQ3xg5SMFK5z1oBPcc53Gd9Jb83WJSCCK3O1Ld5j0DSNf2avG
22sb5duSbQ+oJOwSJ8gVwu1j8KX7XxwBIpiaA1cf+kWBIr1h5pGN9FCQbCVXrMqA
drWKB3rZBnROvHLJNwbY0rimGJ6ZPcE7BqHccfHM63dCGZD/a7cFAfubG2k6eUNb
sE9kWSrMwhEkW5BOJYJmMkHq+FgaVkbakZB6VOEKv0Ids+hKkX7S/Y6roSTOixaT
bNLtP/rQX4F7mhsMOFsoKSeaj4bAfPyt7Vugy0VuhiqMOtpO57pXDcoBk2/zye3R
xX/c88kchnozrLJMv5t6wDMpjDjPi70k+fiw9+03z0lxMFGKfIMejnzxeWztvurA
d9xxZtUJU1uwiHqOU/SgsbX6qe0G5BHjCk3COGXtaJvWSH1pb4cGWsPlbWsEZwMJ
S6gu2wLXRKa21d8xdG+Vq1KtgYsf64Qja+N5KDN1yRbJBqARKUaeW5kUFetqS9kU
zd7AWlUrSSQQ4t9PqvFE4oqVtAd76FHnBCLFlU1Pa8ji8TVxfvNMVFa12hLYkptL
MPXUlfHTn+BmtAqgfqzjCiA+mApnx+XocR8GmaoJHpzEWP6JA/dnDJTm15+Cj1Om
BFPf7E/FXSKxcGLDL3CH3UAXt9q0vDftXgrxFY3+I9LLqP0Pu2Tn1/oAxU4GMxTn
bWCz1EIpQ5IyLuU5nMZmWJwaJRp/gooVxNKst0xu6KUxsAIUy7OW7uyejP7okGo8
jLil9osvfeIOK6SaofveWPsE7Y83GDz6iV9OVef4BLpqdQn7Ytnk/edKSAt8ynkm
QAnDI3yan0Cc/9O55gw7GvKxlCePMfUMSrtguh5Hr5t0JFg0ngpxCZGvHkNYvGGr
TjOHe+5qBRaGSfaeHllIQONuuzOnPO4zcTIO3rg7NvNTUClSHTyYjXoNi8twWSgS
Og5WVW8xNbcaX53oJ5qYJy7rN1JktzLMF/4yRqguXdD6r1p5kHt//Seu+nzgu0gf
/yBlcdsDCxxZk769zL1P0L6XYgziZdX4lD8a7WmAjQ02QO0X1u3W2RquK3dr9K/n
DTREDvpqZKRyKNbzIObkuf7Ms8I8GnWFBkgYaV/o8kaSXOef1/qT3sZPzkbEQdpY
xDT79Az/AY3ccnQtOLmWM2Kmr4vAiv8JcEV0uvuW7LZT4mQTBYrcYyTV7QA9eqxB
Ehuu8IDidI8a9JCA4oG7ZVDw/4DO5z6tTiLCAB+Vpdw4hF/YRVKkCydf32dieLq1
iEaPP6aIx6Vvj1oCeuvh741A3FI5DTmzp9wdE7Cxx3KY4AAELL+0rOX56NJGnX31
RGFtBa3vqXDMihFoqKdPFIOW374CoKZZWPAZDnSJi63BdN6/x7Iky23SPOX1c/oy
uyTq22jnI8O/ppBBmpaZdVPvKMOVZdKI7jHzl/MUu+jhO9PkBNCqQ6IHERUCjhbA
KSOUMOfLJN8VrdsdT2BFjz52/2TJznRsI/H6PKUSEc3E44iY0eROc4rNpCCDw3CL
cSfgfOUuOA/30eb5WZ6DTflyA0pbbhdayG/7158zmT7ltA9cXkxREVlXfwfJqNIG
fcaMwwABraWvlEUYuqeCU8FzFYQN9EbhNBBrmqyx+/x0MxohkGQJ35zzp1aFu4x2
qPPc9JK0Lf535bmu5QUnNCZvf+7NMlSNkIk0/nI2/Ojt9Qy1oCbf0NsiaA2IXpIl
ppLbnqnBWKqIcnY2xDY3JB5hTTzJjmGUGHqNi9Om55EU5dDjcUWgka2D5sZ1V91e
YWsGX3CYSrEu/OLeQilcprPKUUL70pEBsft9p4KSUGh+RAd5oQWDd7cDZbgqKtPX
EhWpanOza8061eFjuJmVXqSRZV+IhEYzMwrq1woQbXqFBsCt/W4xwk967ETiOolV
3gz5gRo5IIyAlCPQifL0cfG4Yq9yDLKbGstFQY9U8G2FHQoS9jiFEpqFybYWcaTq
BNgNAeu3SHZLsR/SRj/7HNyAyNyGaDRmsMZCK0telsOUOAdHYSeejQcXidGIcmry
bCNhWsregSGg+hSf3K3vFLLlXnLTMjF6oW3krqQNlnvBJ7tL/7dmoJJ/cv/on7qT
cbFGadZXRglLwkLIMsU9FGCmSMO3W/EhhWFC0XHABP07nCOBx8VWjBag5SOxHaqj
PSrOUhYPeA4oCzRj9jtqX0rmlw5hufxV9Z+obvVDjSoh0OQSbnHYuzAZqvKn5dem
LGpWiDSfXyt0tbJO1L7BwMlYi3Ty/i7E1nCWXF2hQPBzWiq7egUhQkNJhSTov7Lt
dvIKmpSdI1KCfgVQbRvh/EJzRp66B4vQ3vYkiq2oXA59HeEBIet+a04fOeZUXcgf
ITvO4uCMhgMUZBqscGRfhAckl+wFpArZAWG5Jk5JcscVG4DIQ1GI7awci2foyhYe
rOUy3Dd/etM2wIOJXkqXQ8AhAU3tzAV6dDN2Bk1UXbg2FJ/kWj7+8aH4pAfnuvgC
KUuBYlLFL7XZN2rvQeI3GMsa+as328doIPKvcb2YJioR/PkMYaIC6/Dg2rqCD6pt
MNlYXsrTW9meyQA/68CrlFgYqo4boYWtlKcWMVNoa2LfBAvRPkfN0VXbB0so3sha
oZXbK/HzX9eBXpL8x0HEXSLkBnwe5oaVf7DcLkZ/M8aujs+f/eF+nHjVfLsFgpLg
7ejfi4u69X6hbb9CeFFELOpAf6HuaM5k0SI+dRQ15zTUYJ1DdbZn7Heq5gwSE6mj
C+/LNjgNpVoOfVRAeu3OqwAnQ4NBdUkuuyaf1eBu1A/GxTyxLFVleQzmPrL1BXRO
QwnQ12aB4s+BkYbHc7/MnOBvq5kZQP088R1iZBPuA3F+LYB2IYIXfJGpwsy8BzHT
1AtrHAyNgDGbEJb/QK3xyJJVaWRAz5mh5aVRWdFCfvNoJqXYWKKC1tjDlLJMlXVC
+QzqgvfPDHRAjUXjcMZtKrArRyjh5gYenek6ZVx6R0VcSM2DDNo/Nc4SbYbueIMW
iH2oJOknfR7ZmfPfdreZYB5PiK7urowjIhZjdBGqAW96LWwrSzGBMRwHX9+HFmiu
EB88/2MJe96KqZXCwZW4bHUU74BOxt4Nf08ybk0xVfa3Qa8MCtCsVAvRCaFsyoxd
cEoe9zv+tELotu6QPhEpc/kzuaAY8ZcdInuG5T8fkNpnkyBReIuA1DJuvj+F8Jhp
Pdpw5/ZrRil2UMTCio2jiZcg6IuWQWiG2OvB0k4C+G9uojvTourlihXcVqMq6lEo
fS6Qb/bkXA0xJ1nIRcrVvS4T2wZqlV3AEdA72gKevlBYb/w4Isk+PnIyoQxPRhD3
+ATjF9n1OZ3tXM5Bij4cQNE+GdekY5gcLlui47mIRMSC+a/fOqhyzRFvpxdeMed3
0Ln3OFqZ/0KKskNTcwmYANxZ3k6HK551iOCQ1rzzElt2hM8lOKWUwI2f3OKfyOQB
rsnbmBJX3O4UTRV4LNbPaui492nEYnkyP/kAHB8i97EzPZhoNFbj97EwRg8+Azqy
fVWmzH2teFSb9e7gwvlI377XqxdiIlSM2aV0wc4GP8hZ6BkO3CkoWm0gRSjCBNCU
7w8aVIWzvOXFQ6yciVsyhn4yzBzEsUSRTUTNrowOpAG4sLxq2ZouwICiPNxXDbwR
gcnuWBdcuPim8L/IK/nI03RLkIORsvx+ADBsrGx8V4egrA3iQfDZIghG7tRTdoKU
43fGmaxI6i+loObKTwwiaMUALG36qX2nAbm6lpFiktdwj03JwuRBJb/tJ0PVRfQf
vdwChUAhdZnHxPrHsq65aw6qP3p7gTBTgwi0ioBxt1CdqjTGvYXFS5A1h8hfKuh5
ZaWpAb0K33G4TgLyEXOOCJnWX7DACR9bZ+7UOwhL94OAMXjo8qhTOi1m1P59RZfh
+O305CZMVyfafG9i1CbiPzvDmjQoasp7QGVuzaXOdZjVdviSfdNXEoE7KVKmNCO4
OjIftZA0v4GoMGh5g6TD4A2iVuMnkAfsZNWo6N2WU9pWxrwA1Oi8CuHQ4q22voeV
lYT0rkzyFUKOMvj/69/2eVQTgcnfks1qF99OxvDFRKlSYXl/a4d1akU7CKN1BeR/
yXLt/QeRSmjVi2EXD3vaULfsqyvMP+CH/4OCE1dE+Lw/n8N4B0wbgtm1U7Qqjlpz
2GhsYqO/ulJgAuDBc5EWln/bcKbLNjVLC498+F8dVmNTiicdlYAL2aQ8TVaJiZLG
elBzC6zvu5D30fKvRKCTWWtADwKWL2dP1XvIc1dEJ8Y0uTWVUamv8t2vQwo7geT4
yycEB9XrAesBlBgHSXdI0WVVhiltQ2GaDZtX4cVRihUJX0Ikt7mpCc06sb4AQcsJ
R2xg8pPtYpdHVxuULqCSy+L757WH2wigII9iWTQPZIu7TMqix95jb1zMnn0cuhzi
38UaOjQyDnvTTjt5rIqCQQ+eI3D0qMc6304yx8Eoc+29ezaa2dvIWo7j3brzgC6K
4JNrB7e5aNe5cnC2+6db+u1vGXNqgXimY+tVIPtkelEzpxRGoeugUmUdeTX4OJ3r
NQ4dYyHk5Hz5zFz0rY0fdVvt0BuJX/cs+IFMlC3keDAoFEDoSyCwDi1gpR7lAmt2
V4c278+HvYkAgzHQ8v3UM6YwSbn3/9iaGgMCmUIk1r0fV8wTGg9NKJ9+pmTGd55X
OEkzu2Ir2sbXNRqjj2WkzCoGUTLwDAmrjCtDVDLCzvqmocnSq5C8gpPbBuYND/OB
0UVeuDwIbQID9K8v/3tQys+rtWhXRAaam+IL6LBDDO8TFPzj98uxUdRdUW/6uijm
vKpTGg5EiixO08ROhcGin91mLtWxCqSL6a+S1vu278++NGVLq2wKWqqyMwFo/aTO
c4ghuI2T4X9frj7HxCoTlk2O92RCnjuEqE1fZGuaOIhPdY/8KftHLRu+sBngEDMt
GN9cdJznqZuN8AjHYmQoZpxfzNMMZK9kCbYrMurnZUzs38mAUO44K+o9mSmLSNjG
KhmSEOcLXcRiGP7rLNp5msDjwd1pFVC5Rsq/v/dQJmTr7BOhPhDRZ9bdOF9OpwU1
8SxtoMYF3VDt+viBG3uHtlZEiFJIJH4UOhK5YbDnk8uHAXg77WLpMHijVPQ5jojQ
k3Alvibuw75b+e4+Rplwm/r+8+bveyJn0Aea6opTS5+Rw6ALtfrSYJLYYg+GwPJ+
DztwXRrUSEG1YKNSI9t+NaQmE70IdZootB/Uos2RaRSgD8EBFINDMMTtmEjNUEPm
F7aM88gk2ZK5bZwwvleBq5ZYQGFNmv36og3lhAbRXUQgAAqKK1pAJK5D1/CH0JYI
cIdLNO59sybKDBAPDtsILyvTaAH/iiwFv4tLkUnbKLQXIqFLYoVcZvHIfC7sQsVv
ozQayAS7+9slHbWXMPMjocfXcIbNBger3m02zolgORZcs3AfZcxDu92gS5Zi6Rp1
kHAQ9mUYk6VmS9iPx/7HW4I07599TKrj0MUj4kNKzYEDVpD/CjApJm6AajCldum9
+LixEmahIwsOeFwj0qKdPmphMMpjKtGeNN+qspe/FFh/5bsRisfu80fTcnp5GGmq
HBXtoGtVRZdmkNpFGUjoZcSKPPmtMjZrDMXpebKefijbMH2EuSuKgAv8k0E8epGP
ZXb7kZj+kNiUmuLzMDZ5jC92IXwMehBpRNw7pfHcjeC8Uo+NZ2+XWq7PWlgUPGby
IzHmFCZkzR7ULhYEzZqXgXFitTue+biIJH6qUWGKp7S8zYEFNeuSsDkMP2eMVPjc
HwXveCBFFWeWf70EGBA1uhGmQLXKsaRgKyUfNLTBHeasV7nxJ6ZIoZHXBiO8F6QI
qcVCgQf2Ui9GiroHoH3DHFOdKuw+i1dL/lRJJ5e4vYkI7TUh0wriVSdtzUXgdo/f
shdjOrGhJsCPYQ3erBCpaYk86KZtvhlTHu02vptw6TvPeQvSGz0TtR/IT4syRH1N
31e2odVrpkf5VO6ppa0zWjHHJ4iAM2HFXdKaybwQEwcLlt1PReAFsPehzXV1rlAl
4szThE7uVk8RmIiO+APGYS+bUCoFkEvuKtkcvEIm1lQfPOWNAGckRKqSN1b5YaUr
Zkyhs5Vaz6LVxubdqrfMeRZZTgLbabmmAnAHweHaIshNG09uqo3U8ieNCu7V/m7J
4tpj7yPl6dSyMNHsj05HIjrssEJQFoZ/qu4A9YcziQh7fypQUNd7tNhZ6/vBIKg5
fmAosYyfnjPdAQErCrxE3BPcWFCmpQ0yXDe5yFMgBs9zixnz9SBAngiYAHFG0H7X
195XMY0ChPdm5cTl4ImdIQOVZwfGWOPtV0K0SoCNs3xrl6R5HLMaXKVcn0IlEI6j
kzaoHiI0jVDUd7MD8GWc5jQiKITHf8jeG/aJXoik+5aAL3ooYO2trQ+e4N6qDoRu
GkpcU991IGimAACCj/eJOvxa/vwZdmJYleqYmI+YxN72Cvti0ccv4yZFI1GUO/sD
IvOsaAGnCDsy8Upw64ILcdvARNGFcD73fHDVDpjLJuNgxfxyRo92uc+VObG7fiJa
vegd/RXAVjga1eYcz5IoCyHgEXhNhfSPEcUizp5y6yQ5Fd/RBBwyxdOlwXCJhhyH
0Tpf9W1yvXXSiYomEoYIP1m/REQmejRTnLb5CmWFc3hDG3vgXonV+DTTwtY98UHH
9Ym5RLtGHqZ4T70xXgrDuuKWoQd4ug3LXU23A1uCyPa9x/1ml9zRgMYBudGFhMP+
iYII+5PSCV5va0RItsdCSi+KP+C7s0N+TcRP++esTuJDSRVPjljRjeUF4KbKaR1W
PCT8Gp87Snfoyr6Curl3XFg/bw7OuTnfG8p0ZNhYgQqkC5dKmYLncO7XXj0b7TTg
FFV0lJdpEHZ8o3hxDdMUlPz10A27B6SDYFipjal49PPjq5IJaSlYT5JqKKwO/4OA
zTWJtAGxdYJR659l3SvkhwO5cgExDNxJKuzX2zjMgUo67lhq/f3lnvFZK4MxoLBF
G1+n3AxPx31IjDoXVoGYJWJYSS1oPe22/18HHpHFcxL73Wt7X66NPjCwP9FOop9l
Jm0TW6MbNcgfGILHGltF8HSqWEAGP2kssS5qNtRi1Q4cZfsc2vJqgoeBsj20+Z1T
DoyY9WnugUNiKkZMxRh+PEDXm7/rKGuSKT0Pu+X1lF93s+sGxf+6FjZ/ZerqUKXS
pl8MwJflj1PFlFNPHeIFmgCLkH9Nt1ySv7heMn3cB2POpiiQyjOB6pdv3Iou+R+l
SPoG3daaqQrisMs/CuFKNmgftboNPL/8M0GAEl8GWhOeI/8MkkI+xNNiCNcmN/2q
yuuC8hz7mDCjRtD+kJwcaB8XCxEVMPbfPRu2WzumOE66qguCC9a2cgYt//loEiBH
Z+ppU2z+0IaiNOpAeyKSWT3w9ub3UPUMA9nFrW5QQjth5S8+LHs9d3ZaZ7ubY76/
uLdInHj5A9nGJWVR7NXyTVjF19WpndmYnHdnMzGDl7UCYvoy1Giu9tXs47FIUkjK
1y7aw7qbq4vBUhslHiLZWkNnc8AK2woitfxiG71TW9mE+ME8aG9DcFO/jP/mRzzx
B0NpNC2RK+5eJu7FlQS8Qe+swDtouYgEQzPrybAzIzcz7dDUGowpJEctqk+70fnf
qLiWLsG+YrH6yIVmq7TW6V0IUXZZa135Gm3ubJfTymJYsDPdLBW6Y/sppolR9dLB
Gq+BKBK0r9juDSvVmKaXGSPMwMuv4S9jgTegV177IX06Kel7GyKaw+d3tgnydoPH
tD8o5O46E9gFTU09fpDPeWe/N8hHrq3cTRD2keYoAzHuAYUr/6VuJaNF8hM0JPT0
Lj95Hxlll8Fr2YKHXiilny4padan5BUGyl+KFdqmyMgHQiQv+MmPJrzdH08uV8eo
2Vxp9cANMJ8ic6sJSvOjVrFwvaOeU/LRhvkCuRa/LFExoHrL2p42AwVwfBfo0PWn
BqIc6YwEXIDA7vOuE5ExE5UHwa+g3vUqOsGslFj/+9jIjXdc4g5Ou8EpD/l7ltni
vw2nB9/FKQ2EuUJXFxffJ8CCviXLP4paQC1vOJTKm31LltdUP2xDEd+dH/Qd91XV
xhyGzvietj9IX2jVr5tQ/xgafSPmQLmlA7/ItvWB8WM1Oeg3wq5kIrlgOtUZB0Wz
nuQh2vXzq0Mm8bkVOD/lni9uGuJXCzlt5aIirzR/iDhDCBpoTeDMfwRNKG93oszK
tdgEIs0QubFpoHTXvbwiVdbagVUCpjIuYozHwv8HrzDS7jAdYpiJCF00Hi6WYhAO
lwTLvZl5ni8tpiFFrO1eeRkDUKK/u9xmTYBPAC3YF8SKvXQGdlthyz2MNGRisn6m
OqtPUosk4ojx2TaHyIWiOIBpo+qt3mQ6hfd/SiR+3qtUykiJq+tDVOOrPtjJIBW6
ImsAvdY4zdf9YlmLaxa2IEC+L+2jsPGGvype1IuZXK4wjcjRAiHJCwQ+SgA5UPL9
HgzhtcKy7uAjEJGoQmhHIHzMjoZXXOBPd8j6v4I61nXU+Qtw8zrf3o7R7qnw2nHU
hP5GOkC/aJW4uZnzPm2d/kxhXOZ9YmNV9CLyWzkCCDk9VIMczdlhZDYwR77Yr4u5
PB5KCwsnRRStquIQcQNCdeL+JpVn0p3iXTdYhr/MS4Hx3FdfAPtAvVUR9sgu3nFR
gb72RKh4t79y/G4We19j3C0z9nDRBDNk6dWprIRGkebjGDyNkz0aCxy5gtmf3e6i
dNH6xwGZapy3FKxcqFR6XL9lCt7esMHp59HNhDrR1uNgkn5QhDO7yPee2r36eN1W
hqKCFlsZghzADelkh+T/oR+kuDvUJ9VdEa9Pd6W2w1V+3RjtJTKQN9rkwC6lzfiE
6mscVPmC8PvtrwRMSOU0U2iMBYgkoeMsrJiDQr9PV/XpSrj4LkWEI0fQtQhfWV7b
4YuigeNbLJQCGIDEJETYmQ4kRerRdZcBRn6RGmD0rriyzveDKsyP1/BfBUz5tTVA
L96NR0Zwcc1NEXFPfexWFGebNrAVnPz9ztEKmxqn8itXh1daKycStvPffwYKqJUp
3Gj+fuWAqXNNhaFApHauNwNLMs89nLZflNCNuAq1PEQw5GlFIMRY1+4dnCQQafF6
n4nm9pFKIy8j9HiVJMgvzFmBvEdArhcphyrlGilquYs+B1CtpC3GY9rG2/QUIeCA
XgVqCCGFUXeQXNJVnH0eeIO1f/O0l3vmw7SYkHoa5z5bu/2UO28unfJpChAayG2x
w8ZT9Nr8P2V9GuHp5tUM2Twgzn6aO8PlRTEkBkLF1rKs1EIcbbDjJd0ExcZbX8mG
+9Z8i3rzaZGfUFj9Igj0othhV/KGBl90ugpAadYkx6JwcGxZKD/CEkek206zvs3H
0Ilkb4cEl5bxyqL37av5nCkQvDuOrNB0RczhChRVuwzsc1Vzrg/PcRQYEK7Roba+
ZIyuWC8VVt9waUKq4+8Jqc9MqokMaDnqe0+9UxlZk/FTuGYahDUohYYNJWwzYCKm
AiilV4yIeRVEyXoLPHw721vQXQus4UoL5MAGZvQIH/fRSQBcqI2+lrJNwMRnOf9Z
T4BInyUaikeoFxna8J01S+3ps1jT4Yi42ErxvyjKy+oZUBH0XvKdoC2wNTp5biwx
sGbna5Oz49n83g7tXgpW/lD/1Ccj3UzGWjTG8v//nOGMxoc0ihKXdRHY16vR25vC
jjZOSzikooq4OkVm4Af4alIkerQFcTSMVkYwaM43wHjYEjKb5zyoSIsXlGzz3WvV
SCjRJSnAAg4n4jQ68TYOqP36DFYheWGubi+uqjnP5iA/EIOhQUiQMefAXGAJi/vJ
TRTR/+iqdJAYSIitOGxMax+Cnz/04ZtWJvOTBFHXVs+0YQ+T/NOYgmyn2MOpxzNQ
gn+idRLcDWgT6y4Rj+YOf6cvTu0Y+cDzZLttQZ7cuGJ5myibMeE0XAGFrl2L+bQf
qX95CBXu6qhPH26W2SsfK8FxCV8pVfAU+PC252tWe2fE8XmeTw0p5XgIJZ2kWD5c
b+W5gTr9zXGCDoPEwjFzN0av+Om2oiTTu542wxWPUH1GhzWYvmHZxehxwDwMwCMy
XK0Umyscbkvedc7AfEfSxiUCJWpB0ayMwMcGLlIHEZXK0BZF12uIEXyzmk/8Tjyj
pben2i+kbqOMfn4OEwySHLII+C8PqGgMcV58c0HJFr/ZLzNoHEBbowhkBlCsElK7
4uAP7BtL7A5U7eabMcTueUxMuMPU01bzooXQUoWuytObGG5WDTGkjsfVP8flIwJs
0Pvh3fBRJrxew2mGjeFPFvumZ++7YL8D0vD/xRUFz3Zj4/emxE+yAG+UpJiNVpWy
g3Y49n3PrS3gnJ+NslcIMXP/iZuHHb8/3h33k7OywzPS5zC552vcIwZAvsl+Wali
FsTmxkrxH8EotkXWTiqajxTKwXGsIbHPREreDFWoLCKMYpw63vYARuSbSzyxodOx
mg94EJ4NLPzTZUGDLz5a8EX9DsXnlV2bZQ4863YUiTtPcV+YX0gISXiEAhXgENKU
bgNoeAsNoUdF/nCTl610kCiLcvBSNpez3ucRpBzDwM8/JJqFFiMDCf4s6khJCZQT
t2061pvX5IaJ2jFQvFF/rtMa6DLNOCQEd2a9PRycBJC45DCF5zw4lnoI5iAltB3D
CakBOA0uOqScgmoFqzeMXdmz//T1v0pZf0bbCUdhYcDPXh42XoxiULy4zC5/8Jt9
tKRpznqPn7KkXlDSTa/aLwZjCWokpvSmTMzGGEWBfjGAj52nMjiXEDq57R29s/21
85ZzEnDPuO1hSg3dLaDjw4EBGva2Vt01t0Zt7v+PdDfLoZDN9Ix0vX1qK01NZRVO
Fz1YZyokpt6sP+uENf1IjUjsjtuRYjhz0FQwdDDkM2L99gTZp7RucsrvUS9HKiW2
1HeqSt4J7CnnAHWqXBrXT977aFAjsdYb0lH1yQ9YiC6jMp6/z6RrgdFhBAdgkG/C
lRJGL1hKI0g1Ar0/rv8b8if2ufmq5/uSQxXLQW+FkaoKCf12B+JqczcjFo32IRJe
L/lV8E5CfxQBlEzF/95nsQ3x9E2frARx38UUAFvFLx4C0IVj87uPbSfAybtobfpN
35hwXpOPvhhcm+u5HE6uNzQu9eYGFrR23DWOyo82ucakKIc1vfg1Bjl2TYFoXHDJ
uiLKKwhrYN/ltdg0lGYe0oib66I+O9MS2+6XHY/aszuYxTm0+6LSHtQhBPJ0MmPU
IoHTrG4ZOX+AoW4QYt1NKhYbouo0Z7lQ8qHK62P4OA3kpNHusd14B0n+pV/RZahF
2AfhBxhlR0LJu2LDLzVCHI5ug2GQ5y9W/Ikv0wR7yH6IfD69JVvmaOJpzA4yNSiM
5LliwxkfMXD1ciWNpdv1gW9ZXynQaqQ0zs+p2bcN6nHl82JIdBR8PqN1yNcRsxSq
EIL+UydDMQ1Kt/wZTMXhpwa/sHeY6jEmEET/iY0imH3buKu+toZAsVgOU6uYTRiR
slaeECbNdQeLm4TF9ZAf/WhbP27HTB7pkjEWmab4NtWo75r/YhV6F7GOCV/jv7dD
VrKpHzWuNOad9bo5RaO3IGFN+ha3zoR+DdMUf/TZZc6FSxNut81LLCea9hsR/kVV
Hr62HN2xiW7RPkQbmfCPa7tS0urJxupXIXGcGL02sgneSTkiEKckFn4KbvfGUVxv
fiz/MXFZSVEEaS+/84e55DtkS4KhH0lfjKH+8cg0ATt0gG2ulMxXKCXD5NmxC+1D
ZinshTMCD2xjlBWve8pSk8NkqWhWHnk9tV8Y2rOdh1lAacbAFdHqTxvtXMpMJDbX
P/1kWyWTSbmIo+E2o1ak9B/SL38enbDVZmoBMcol6D7/U0DznEhSHH0OEHRVWFlf
htg7a55BAZ0AgIOg/3ItM6SuCp2t3J3e8XTpXJjuHBovgOPqI+8UniTwDv+GRKfH
Ta7IQ4PyF1ubErYMS2o/dz7gxm+OBrGSb+b+9O5dg2ZPrgS9+VuLvfMBUUuDFzr8
z58uOnqGqOB0mzfr/ZmiutEFQfFHoGkBC3bv1rXUXjCnMeSr9/Y3p2e1EZsgPq5e
bNKbpFHfcfHnsPZ2PPaAXIgbNhbMwPOaTAzCHralwJEnQmp1Kb5SKM6sVss3BoQq
TfaKQaJktztEx6hdDOYx4U6Ml52tQMPLS160Ci/kYAbKmDp8m1LotalpWReFM24g
Ues6rBN4Lq3JbZLAvVS5CEZavBqllLOw0oJcPS/IWvbcWXu4zQ9FRzNTcYk2FAv/
eLxLFGSvD7/govZV0CygMeuREcnT4R8MT5tuvr51NaTlb45881S/UzHic/ZmOsvr
xHLOyRYUOILqkzXPtXFTb94pJG9Jh8Mz8d2N1fvEMyWNKkmf+r3FriBnQYmv3TUY
wmBKYHj3fngUkhA0UMWnEXrqSMMsjNnUQnVCzvU8eAj5piXTSvVevhYOa6tH+DUx
YaDiV13hPGr3D2b3RofSZ+/H8QwlXHJomSCptp5v+46GgD90ONTgLnvs0KlKqYJf
Tfu34K+xZV/60CI8X7rvlCdFbCr1/JAXCVj88KRDGB6Pf183ZXnDE7682j8UkgTh
i4AsgAEaqQsuWJ0BsI8JB2FEK7Jj3KI2LjFaNdtxU2K7eEtrC/R74gJuVEJxT3RM
ZeBbuD7DVZumkfQ3JGwViTrXzpxeHQTUOfHh4/hOl8TTW18+xH/eUIoK0oiYY/ar
sM2SWc4SRRFTI4TvIP7Rce4js3iwKLmNHDhf4UoseIoGzTm8CXBis0fftZPwxfSo
H702nZ6J+7AWDz3xnX0t36Z0qgD1PsEk3vJXnkQ8JPQ2LiKBZerWl/MHNgsJzF5F
y5unn+/sX9nCllUQQnBy/qtGRDy4FSl4/wAj9wug/Lfhq/8lsunB2BAiEOeogzsL
CLc8nd6mnRMcIkrUim2VxakgIXYSlVRYQ/Ej1dQ2WFmdSl10umMFKVXzDd/5CmHZ
W3Wfgu7paITbM7vFv8OZ5wFzENb1uE0lnPitgr3Es8pvpYP4QEV69U/RF7SEsmYI
IVd2ykEO7LUVgHn2mQQQTNMRG+wzx4LWz4Sx/EQnzG4+GHFgRD2AkIeO0KlX9q1n
Ua3dha0Guglt9MtgWftjfowcbmA8XFLpTUMPFuaHKhT5nwZ3IINJnE1pg+rHTdzD
ny1TGC5a+ndimrerC+iohqBIpWuvXAD2QgTBtb7uTfyQJTuNTnhfWWMcDeyfql2h
ObsWvBLrBPUSD4o8eQVdFeeBhJWzmPIGTPQKj0aNVUtpirap2l0ZOkh5kLHZv9wc
IEkvyC36BspkJOAxvY5yO0pquIsS53/3QN2ZYMN8vPxfRAtLwiQ2Hjh/TRDG10Tm
upuX4V22BB3NnfcVj9v71CDQK3s3ZhEafxjWBo0TMbjyii9G0bvv9S080Mo0HnU8
DKp8FZLj8BdwnqLEUtt/Ru47YC0VzMUxSRe0c/N0Vzsxhb87pt11UA8tO9M5kgWQ
scxgqeVe1wMN96IDQeoqYUtUqJAvEbOGXR0Xqb0VYzwhjzg8LTVG+znSbPyRvvBB
UY1CIkwRmDgKjbt1mk6gW49rUcfiq3cVnCPRYLmKnqJ1u36JoEWX6ffaEcyYMM3S
u+5tpwaW2B4FeJxoAdTJgBxstHlDpXEbCdQrRV1/lySlespRkIbcbE19Tg3nJr3d
pJj40Rsg1cGUhoI5FZwIGAkBYSwKLmJDKCXLh727gYv7Lf+WzXxeom/c2NGNvoba
wwqVbgHaE/cPJo4DpWN9rc+NN7jAoCvFyQxi0YsxiBJV8cbBsoY3w7ZG0l8I3HzY
LvxmbMoLBoGXxC/S2EL3BWxQ+vUJcMQ/RPExTv3UMvErZU3MEmYkH4GQMSXcuQNC
cLvR4rccdqgx4me2BtIFbgfAS1eNJwh11lqJJrNNv3/uXR1o9gVYz9yLWAZo88SN
qZ2CeMMSSimzWjXuOXY7bfcGbfVjCz7YoJAGq4IvevfKXpJQWrG4VT+K+e89yofJ
MVEpoW16CKX0/l6vbP3/NEaqwhB9HbvYZXRG3sogRRHyrjIyOdfNLz/F0ZdSApjN
vjRSp8oEuKexsxoHt0UgIx5kXnqEo5Ph3bbFxkZdiRSdDzFPWNbE7cWH3Qxxka+d
TLJyk3hDX5D2U///TDUhSeVqWWLN8vDYr4rT7132W1xQgYJ72LebGCF2ROEhBhTf
ZBWKou3nDRX3XRC1mQ1n7UTuawJlJnsa3LWTGHPAuct8bSYZDJwEngY/rXBuT0VE
PSZcDUAyzWqLa/6ud3i7b9Ol6Q0uwyQP7r16ntyRm7fUKt1xxZICLHS6eMzvWybR
EZRpT+rAXzhEI73uIutMKRFrZFdhVdSNt+Gk691rxnbt4f6mYYPREPwyNh6+NCMi
8ApbnwZFr2SjuSpbIUQGXERLmRUA4UeeZXyEEvO1qMsyFm0As0v+YP8nIEvpm91F
FjotxDGQmdJ0dt3CfSTOVUbV7cHpmD5x9qVpt9W++zxRyYny4aYU925VDwfEsSEC
3JOWH0gH1AWnUmupsHU/R/apW/JfB/JuSNNWePrrbNUxoHXZ+GohjVaYSb1xRgcs
rk7l9feH6w00LjCoQfGk+ogVYuQNNloc1GWGahCmT/Ja7QPjO2PM2wNs0pOQLsUo
Q0Sv3HERAiAPuVrZ89bIzERvJwvkHU0mRnDhNYCLyDZIvv+5bxkfFZQmUQYsZJ/N
1V0mev2tAMTI0tTzkfRK6refe0s98TKjyDmTEBd5ocFQyUMf8rMwMhKJCp0AL2EZ
yvNA5brGvEWuHS863CEzlt2+e8uuK0SKgNCFTq68hQRAnvzjWfJ+83b3c6in4FUt
YIMoJMAtZoyoTzqv3I/cCRrj9wjfEuQ+d6aibbmBFVt6nZg2pxIjiKo541+RBlto
DBthEwK0alkphJGvh/+azyNSIsRi8fcr/Vt/E2+hx55b8kLgnzp6nqIdG6nlDDDM
P5gF6cH1AusNBn3SW9eoWfq0kRbs8riC+w64EP8dYmtti68MQzHyGkHzjOcweeFz
8CwdEXNBbk0vkd5frFApTUNwYBF0Jf+Nk8WtaoEsdQ++TdnlqztKd5LCG+I0PPnl
FRH40kSEDPj2+u084Lf66gMJzfn+kFihGTuWcybDCHZXKCYpTAWN+jk33VCRtTjf
3WVjJk4Gcvq5F+QUja/cu0Od0XoBwe/i30ZKdoRJDqw+AhNAVRoOgOFjTlUUz3Ps
h3fRcGLYaP0TyY5a1M2Ojuci3G82JefLlm2lz+8UbCC8HzkJx+D82+nPShfk90E9
G6dX/QCgqiI/wCj9YlL/pcYhBueU+ZTtmXgqPbdCRBfHZqPmBnOsr+TNsnMRMTze
9GRQs5szZltnW3JhvezVAXjWUvvLB0G+2uE2cTp2rzgwx6ELSY8q/X7+UWGRRFVh
23r6TSIa/VN75+ZBbETgPPFFXxuTwOc8PUZFzkVtAsG1grbxpVXU5OeuJAFJh50Z
8UkAvW39As60voq9A7ztPKwbwcK8VsDHT+FA2WZfV1iFQdkKl+0PkdOKzAq8BkV8
NKaPZDv06AFNdKBheszwcjTxbcskj8BWFvlLrbLLyqzHlE46LZbzWwVbV729YEwQ
Qbq1dYWw7YJwPDnBsnt/pkImLFae8QDU6bH/4hMDdnVasfFNYbGHKanbHRtloRz4
mSmzxIc3MTPmwXyVgO7PKSeHDfvCQmbi4YOECsi77XuawbmOeMu1cXRMs7qxOsef
7JN4s834rALmmTzQHZWEQyaFXDoJsMtMXIS8IdxJGBLtSPZj7qdMhTDdx0SA1+wv
ZIF+eFN7R54+F/CzXb/PiLFJLAkoeMgjwjj3XxEYuEYwCL2LLM9qCd2/tECl0mB7
J/NmdZ+cgeeFL1m1uUE5sERs8Mr9Q8PZ7c7AH9YsCzbLA7Nn/LVkdyN8FMadb7Sc
IbLr2Dq7re18huG/8rbDFIr9i/ULcJ7u1HlL7Wp24SpB5JT9RKTKprg0khdy7SnF
6vgClHSDiBZd/KbgjxZP2ZbxmJ/1LdfqCewhSn8x4tOPi96knjmfvk9z7qs3rrGo
wdGqy81yKY/G9oclSPGW1bqFY7FSHja4fYTJxXZD+vCEEbe5dVWboECHp/QmO8Mv
eniSxaRx+VSPxvGAC3nDJsys0pXtIwirVtDMELZbf+RRyySTgpDwNp0xSHwA0Z8u
zzF/Y4yp5edm98he1cU0TX7119of7nO1o5U1iRaYaQvJfzKidl5dR6cYB5CEysoa
WchjFXdfMNr5GQkxUAGIzvqcFTH0ln7ufgt4psA3ipXRweXP6cjmNU5M6ZuI9VV9
sX8GbXACb6ZadcD17TnaXkWZlbsCbZnHZDVdOs+GlhAb65MjHe6qshks1xzEXbfe
+MXGITMyIqUC0UTKw3X4cyIHvfDikwZrJ0dFpi43nb1bWMxwEbVVLBWu/Iz4uD5K
aLJhi5uTfvieY6gPdzoLEnml7/LtUjNBQ6GBQUqyKJLxcWT/72ZPOtMPyIUnQr96
y/W8rwFnP6tVvb0BrzwImB3NJ6F7O+DquiMBIH+G6roEP12r/fyePRJ+q35HR646
Hy6GhSVkAiQfXCB7ohiEiBGHWP7NdnKo0PtR0OSSPHY7qZSv/RoGE0flBMeOmN+Z
h/0yc78F1LxTxbxckGaMJt25gxDMLT90mYKMUifepO1+wLHT0nhMeAyASTcfEttb
6pFLH5XLjU5tU+hhSn3BewC8ATAmbA0abhGlGBCNWh55MMkiF16cDZsqIq2qyWke
amoKxe9ejc+18AQB7JZTr7bkJZI/wbRGFwZhW+qiYNgSmQKI+rSznxqoBMsNiRHZ
G9uYontb9Kqa2nuWeeeuD1HNvITNrm450Qcc+4e6MnIbGucntmB/0JBWmVkU33kO
ZfW5N8kv3O/mC74JNTbzSUew4SodVn8pAAKwFI8LsYVXia9nV7vzMI7HDG7TA41b
OH79XaKhA6XZTZ23R2lQs3mpVqMVD5YcCdol9ZNZxyxkbianyDTehbWofeEtG6T8
QwgYcLRWZ9yEI2sasK/a3MsPoc5ThSWIGr3CpBTz0BwWv/KGLK6T+oDjZcOB2XlE
u/+tWTLTrMW5oMlYIuTevT+4wbBEMoVhGF0JZy/Hk2PtUlCRRomhTILc9KXkAEOK
QcMAGRuoVzJU04pzOQ89VqSAhTA7LrD2bH2Ld/XZqcUOpCpdeZ/tEJxj/mo7jixV
kpgWDGRy07Ojou8MYh+dAvBoGyMdaWWijr/DVq14lkvqHL0o99rwhoJwLZTdzF/T
kY117cbM/XOCGdUQlZbF+bTv8iA5gQDHqy4GKbMw/SBhtZcbLd2a+luPCMQThJor
nQMNdyjuOgk5/bCtjEXsvFfVqC3SejRwRb/bdg+7iiVXCg3xd+mBxcJmAFgEaEFv
haVsUq3Cj0mroVSZ7DGzudhvHWqdiVOx5CkwwUGT0xKQKETEGBPMlPWGyZ1Jtxwh
6z0X4gXolh7tah3StUbwhep+8MhfD3XCmu3r2SLNedmK1lcS97xhFQP3wa2nlsyH
feGQvjBT5Klu5vqZUZwGqG5Yw7BMw8QhsraOXiCUJKkkFE7XHNM1EEFSnJdzg0g+
BKHhSO/J6koGkcaP1oVxEVAhq+vAeuAi3u+HK9iIssBSZYVpw73Ne+oD07EubtZg
zQpCNFB9okwEQ89cWaRsgdtglxEvO8Myxv+1I8J5s55nFUaTSlSfP3Ujsq1WFN8W
3v9iJ3PkWV0r4qqaPpguODZtRpHDsGSUy6QDeVanpKxzYGPRX5gSr2ASv1rcDs03
FT5x65MfwKiCZLY1iRmWajCiavFneIV1FKGqHXgXsVYnSb7r6bheY9HM95VgxFDB
Tq7ZEM/yXIIV7bLO/LCtT/1jA+WpiG911LITSS3WGe74gOknZi/OaLLvlLYD+3+f
i/mGP48fstQih0FJI49ou0NCms1OiJ7AUgn4U5hVxkS4fVqptlXa1bdkc35kRmUh
ZpcHdzli0UnPuX8G2sxCkVUg/qRiwyHKDPKpzO79z4/FdFo6/c8aY1rnoFlGtVpK
JCwLWSBuhkzWu/lUn+gFM0q8VoG5+7UxPL5vfO42FqJKpNg0V2fWIFFNX22yd5hi
3Mf6DHkJZT7lhK0KVrowN+ZJ/UbvE6L7i5hKy1rKEL3BXsqjzU3pqx+R+iltFPKl
oJ2t4nuTIIC0fN8j1HCmocpdF225UOqFSQokG/guY6O+NSaSge/HAYrhyx1kMJHz
VpIT1st022/4Yqema5ueRXhtVV7ZLDcRt6Pe1LFcTeSQ4Tyb9WfqSH9b1FYZh7nf
NZx4PTx42hZMhq4eSifoV27Co2Q8ONI3DU5UqsfTzdGlvESa2R5UL1QjiyoqAgoJ
/1vO6fguk0DSP09zZQNJNb7RYiembHDL1awtMEvQUN4GkIdyvnkOA25fXvVj1wpk
BkyBl7pEuIM3Ozvq/SDKxpHO7vziMq2k6tuUdIqiww74TtAIRzhAX+C8NcgF8vn7
uLmETzBDgphCZOkpYe4p1udbIvujslbRA6ThYFMJpNKE/hyIx/VNRzukraQLkcBI
SdkvWkeDbok8IzhtzmfWMugbIMeP5OfQXfxn15iBFrQayZolG1yHUGQmDgbwipFo
vFO7xk2QoBFFtP++8KsYV/VNBJkYH7E/h+0rODP4MbGCia8rnR/+Zqnx4u7hPwXT
HJ1tsGZa9/dRLT+00NCv59eEPkOf1CZRZbzqPv/J79bt/d+jJRc29wLy8qiS7BUO
JHTJxhu2pkMcSXkWJQ6YWFzmlmDZXujaePasVbzjA3awDtQdWeoeFB4QhSxCzJ0z
T1iRCKpEjs2/Z8D9bA8BZbEBTrtngmzebjFPNw3j1c+RzFMOafFUJKhPsRSm2/eV
QLLUSCOI+xvFX6ZEKcSMcztq0dL/hEfieRcgoEMPPagut70P9lhpvApq5P1ulZZK
HeDccucSqaVK3foYGtUd1FNJlSps2EMax6xOFBoag0DwCT4rm6jT1ErLkMDW9Nol
ht7zDGqZ45EBj5TT6dstW3SocJ8p7Zvk9NGKOMNjCvbT6Ye6HnjVpZMjYQeHJyeZ
YvQKlM5QJ/iR3S2YxM4thJPGJi2IA939swB+XNQacCgRXaKF8zvEEh9Wpp1yHbkb
x3xa1/pSPPbIoT/YG2qyrt2OFyJKctxTsk2hZ0IW9LNid2Wkp9AQJ0McFsOU9aVc
cYh31W1wvxYKYHcLv2gNUnnJ8InL7PRmVlSOmUOsx5OjfoF8PW218ttCUzG5n+LT
TtTXv4+CD7A41osR17lITI6eZI8e+B/YLzU48D57zZ72Sve/+t5giPMUmb0ywws5
LFpHKK99eeOABy1O0ykyxOHHNG28UuE+/qDxnD5+T+1RDyHNX+7+zYiceYI4n6Wr
N0Eb8jeg4VLcKbtlevHjW0WIw+TxWCltnJKmlkUgb2gogCtOo7vfRp2r7lMe18W6
jJ3RtsVbC9Q6AwgjUNnsETUYge+7R1QM+e2uBz+nIPIBZO+x1MCioI0V+nnyafAj
9Qj3URU4891doUbkbdrU93VyjEMCw49EOQUBesWOEvy676fIpUxEX8YiT7Nh9X3k
sRA3QfKM8oU8vq3rYWEF89Z7BPZJKn4uegjsGYxCN42U+Vz8Vaq20sLwJ45r6C1U
PBq2KYbSnw+I2lWdgCgFLcI6snu16mmkZtFx8JTd3yCv52wwGMvwB0cF0hnZLeEn
MxaHGcP4qZ2qoLy0gyX1l8fkyve9SgwuCNYuQM/zwxud5Z1sz5hYM7no2uLmtTiK
0MeE8B0en5kAnrrRlZKbTBBIQqISrR3R7XpqH9DH4Yi5oRRGyfRlC+N7XgnR2Vaj
Sy58t6i0Bt2qx8ffKbqwtO0Rx+AGGNQXdAHisrv+v58Mba1Gdsl4UwQWBokzocHB
yiq8PZcSt2D+jVuZrvn7sJVecICeAbnQKQ/vorSlxFYpnj/vdDC0lvZWN3b/GqjP
2GgDLmkSsiIlXOkeDeJBtVfMkyWvX1ViXzjLsX+FQNY+jZL/3Xl9zPS9yA8Ae170
T6rZ26pZ5Kv83dlI2xak/ProfZ/DeWnBNYPqlvbJ8dOrbNbxPNzCGMcE9R3Q0rUK
y8BEx1DOO7y25t/XkrwKp8BgqEnlzgWfPxo7X64K0Z1mBkgv4stQHVxcU74DGUe/
uYAqOh6CjGXvhNq2nvR4JsydO2a1AKuseg+y0YtV/Vn3c2EilaYqlcSp91W8J5uc
Ry0YVS7Cio0qMKM6gfgXV/v5697gvOQIGPwRuGEb5+NP9DO52FySvYXUQsSiaOKT
unqM8OA0tb9Q9YRVapL4Ta2N4ofMbJEi8xsxjt757IkGtjmtkesq5ZKUDadz52gE
mk+J60G+16swFuN+oO4H0kja8GCrCka2/FsgTOD7DwzRdZc4ZkByYRbECrbrOQ7M
6OxVAyrIBzm05gEUz9/3OklhjYPC/oXqzgPWG4mkoje3enDulV64fuiGAXUk4ipx
KHwhCb7oUh+gLwCvoO9BHwA/fhFiKk8df+Uf7ly8E6tiJjmsCen+tYRBkqIbDBk0
nw1cuqiqzZ4oHXrQd46yFtb/87SqdqYUl+ZMg8f2wqS90rC3scJ1F5BEb4E2VpOw
xzgVMIWPi0PwEnquXDCvg0duzTRk0s/hIgj0HzMuBftrQ8c1a6ltxAF63vzDjDYF
VIOvkCaGVpdlkIyhw85YRr8i2btbSMaWqZVSUEJhw23EqwAD5Q7vhRPaVBXpSM9N
KJjfPxbr4pCTgmJEx3XP6O9159iWYl7S7bJ8AOb7XI+QNG1pZVjuDiu9uEFAjEMz
5K1Y2y2eb8WhIcFWiy3I9I1kL80m5wxmHITGoXCGrB60Oy6qs/l6KFbyr/RG8Hif
scgu3K+Jahf9/OyCDj5/3zrBFT/cn5hCJnlRKSxKZk86CLsv6vYl385iJbOU8gJm
IOvwXieX7vylxdklW/chkKxvWT/senKhth7oWYqqjyqPv3GjoBcPa63eaY5YzMz1
0zIOzMH69oHWZ7DJZJic4IBALaGgsBUrjOg0D+LzrDyDsHjvIRsRohkvaO+dz85W
k+LmfZCjDk0YcXPALPGol9TwhiCthQX//VtYICZYahTo8FUSmQLUw2lxdx+hawjZ
g3x+hKGm0rpR5lubiHIQXjFJUbpDATDO9zTr8vTag1DapBRCmUn8PsFNH2knVKbu
cDJFKshY8vH8km5g0/DFXGPJt/ijr+yj7fEPzBqkiE7N1pfWbg5y8wR8lfDI7+WM
m+9aQaUc6jR5bkJuVeB7Nh9IzaCIrbaDB1QHxdqVi0wT+pmVFoF5R3IV/0HnbE0K
OhvxSnpYOhhsmfCJ7FS16vMzLIgdVvBWgv55ugYPHgcoPi0CSd2eTAbU7GM0O0Jk
+X6axw9FFMvD5Oocca6fJjJyL4neLrFHj6g4hGaB98ex91ogQ1m160l7ueysX9Hb
zreqxZdvNhjI6qB4Y1NAVQFxmkR63FilfEq+HtdnBlHn6Q9ILJkNA1LD0SVDES0x
aBvkiy/dakurGTYIvIzJGpzZnAQonXgrbU/KXhPskrA7DNcM8RU59DbDN4FucbN9
9VNWKM1a8RjLvH72D/qL83O5bSuF0tfnkWXN6LarsBtnKwqyFiIE/roY7bT7ML55
+hRnXldXwtau/hPxCpfla0gMct5/sbybynHbhEtBdyhP3GgWOYyjzSLta39ypzeE
OeVLq4V5G+JfBv8Tqr2aQ94P3+oBkJ2jX1hCjE6bED0CQYj9mhfVblP1IZXtIwF4
9xiJTOjqzaHZJ3GNYROr21oEVOkumUOz6q700HtIjG1Msdphwb24gpSPfgGJZkhz
QYKbnEwBruhAd+IAH0TP0MWwfmMip4zMzzIupKLBF9jvEb9CZfjoxEX37q9jFfJI
jq0VjnoIueupvAwx/clHKaxFwD89cee7rB3zBS7joyktk/Ldqjiu8c1J9mxAQinn
m1nkEVRDKvUCcm/lPsnnCzq1ouoQ7Bx1QBfbnfER0h52O02pb2YKfuUfnLRB0V4U
38fK4EXrwaW4RLIZY2+K98OvVbIPERKL968ThP3DRLNKdBnExmfnWiPFzLzQC5Zb
Oj3hLQ8ZS8GKf0P5TW87M0xTdnjgbvO896UePpJ1iidFKNr7UlTCyh/5z0OCOh/x
41c6HjDi9RNcPIGhSlqIjgbrElaCgmrl2PJGwUBFKWUVB2AGd3AePOktOAaNtszT
ZMNN9ovKN8Mk76xjB9kHfkQWaqDVjXYqKtDPjnSGHG337zLRhx74lJPxrCmCYHSt
IqUHYnVn8E6fNA4ewD1q+664B00VCKNRhKPtcS8BZUjd7tYFKoc22uKlBidw9FOh
I9bd1v3FdRABwi2oCX+z++Ji0ChN9wgjULP8J+alfpYH+0elw8WL7dAi0WPAG+us
6CRwPUMwrxxhY+lqcccn/Mxc26+H24VOqmUT54fDNcOxR1NqoXwWEvMLOrzOUKPG
Fm7RspvBXOrEcOyE9GAgTzDi4s0kV40kEIQW2nkxSFrSOsMeP5RXbynpf+Rh4Cn0
NUR4LjnmgJPaTqlLdgmBJrZy/PqsON+VUnoDhx35RKdTcSVIjgSOyyio4PzJ61LX
gV30eXgN8qcohQsAaKIKWQgqs82Cg10A9yO+N3g0iFJ08RqGPN0jJQyWmKobZfgF
NYBymmMoCS9mGdTTK3CCoPRZQzpR8YQNIiZlA0cpGiykp+AOcFRLyMgW6WCtRnXx
G2lANxKvPTRF5xDUHoWH5BtxUO3lZ7sSdfy/OF+QTvdGCG+LlRfiZByUNh9EaYhZ
NCJi377DEP1MSZGiiKWewshbsEApvvwCT9ANn9uvTsQppQ+6cRVItChr2sYkldWl
gen40ApmEktagoDdGTwy2ZfxSiSNGSOAs63pi7UC9QEnvMlGNHG9CqQF/Du7Yg24
W9ICmrv9U1sKa1gVmBvAA+OVk0yqpbFfFMQy3FYHqQS+E3S5hoWL7H0FroXE0ZxJ
/a55s0xhAkQFLXa4pRe7gX/MopqdtNt/TCpyWpUUWz7y+cuK+IaobLM6SdCZNSA/
0xOzMl5PtYz3MXjmyAJ1GJ35CrtfvYxPQZ34I2bsnVTi0frarg59dmNkjYprMj/G
QYtQ52lMGM7Zll8bQy5IoZqsOtlp7wv76KmC29ki7aKGUKdg4apAYccdUAnM8E0P
6vW1vtC6OqrEVLGgwV/veVW6BDLr1aVisH6wZM5M5ty5uDCj4wRqknxac2zJP0St
Kqc2+MHplqKWf75/7w8lHbAVO0HjFptUBMjCnbLMjPL+sx0VkwYX9pgRdgg3zW3M
h7jEbg77LLkBM4mqbM3awlcgyK34C1yyeVPMTBvsZOsCq2sQLEpypBfZ5jAG4AaJ
R2H92xHtBDzSwISKvxPHSUl70k5tHlxaP4PTLMkqHI8OZcf3dCtAjbA+sJPr6TDq
kXF+NInc2/5NVU3ZXiBgqvAY1LBPH2gtVRVndc1O2Tj1SeiEujC+hl142cYh8dbA
GKo36n+olJX7lshgh3GNL3RIBc2LfFj3RyXhioEBhWf/sNU11mn9lSfXIzlchZxc
hcNMwBrqB3vNLW4Ttlkmg+cI+feJtApVcpfKzlYZGd0/xoP9e2997YA1803lHbRM
hnqttf7Ece2cxDg3sy0JxQyc5SJI14/5T9+jbRmWM1F7qESvCZnWuFeousV8qcej
WfM+yacSl1j5bFVusyUZjldVepDrXr6Nan2wSub9h/u51EwxqvS0nX2lfydA2GtB
Iju6dj1dpDv1FmICZ3P0jwH1RmoYfh9GwfIJTo7Y2lvDzPO7fXD4bJKktRLEBpyH
yn/9+Sb8bWkMy5AGUkwyP9xSQl6CWLP2WpmRdXvvtdZNhSn+x2Tw9VBBIjQqdLPh
j426QXa6SwcDktgzBT0rCzsaiggkrh6EwHuNC0iKqiOzgSmknegtQNdZxjlY2ORY
3vJg3PVJZFjHKfJcv+K9oahxvgKCsGS88WI1HbAlwncuw33/Qf/ytkT3nyrdXmSS
8NMlE7REXzXHDOnbNBBidN0yDCHVFyNpDCNW8n4XDNvFNsOvSNavTFildvMFRRgS
kSs4m2OwiE7ZHx7yQgnBfMKFi269LOsI537uwl4KrWti12S+XC2EjyHW+qBZHesN
jdHxJ3JZN1aBmrEL2ZiqZ4J1ALm5xHrEVlTjy4fGEncUqvebuabdedE782DbGtGH
JtFFmZ7gLrHDCI0YDq4LheWHHEHTT06HKIm0izL9mPKcKkpcdUhONQ9voSZtiOTO
T79ej9OjsQyIGN+uWaklogeiAWV2Ix1dzLwkvHnGBboAJ7NnAc3erhKgWeOsWB2Z
B7C4Mzg3GpasFJGHXf+qcFUhYvsPzA9agYyFQEBOHrca9brVtv2J9TvDZvmXwWq4
kZvLqfTFGuqsqz0T1jns2XmLKFslsdloIt2sVoyp0d8z5f1JVxVKkdR7HgoMgDQs
dM6V5Ar2423iKbnELmprdLteZggTKoeJH0B1Yq4oWNvE50knvaV5GbjxoEi9tjzL
4MF+AVmqtBJ/B9EiXnF4GoXZuaKdd2Ifnm7+oRdXajtIaxklnIwaqzk51PSy5Unf
PMjML6mNXK5rzqKyikexRLwTrzIedJhpfhVEnMmo+PnlpsZ2lMLxzhvHHkrTy94B
pqAfNLdu2vQZdQk/5gHgD1gtOSydxQb3ls9pCMDuROrgVrAsCTaQJ3NF5jefY/SN
2cFpibtLy3BJBrPN1vSYGy8eRg4w+o0u7cDKLDCzSH1njgw3k/Qw6TVBzSSOeMGy
ryZY8iuIdIWcNlsTEran9aNztXaxXE9Hk4EJHadBtPYIlpzxFIoHHIa2hrfnsOq2
9WMgqKOqYKe6UjOvCLmtCEkcP/zszxvJAv1tVwy7AHGuAXocxn3ofP4sUjNXp0Gi
pXjpe250UD+Zv7QQr7FqlyxpoTzuYp26id47gs3CrTeAiLUc94QwmYI2VVQb/EnM
TP1Mi5ZWA15M/VOEKdx+9Np4n6mICZZiviLhYWdbA/rRgoq5py30Zxztvn6pzVt3
xyIiZkv8tSF+nRos+ENNbhBB57k2Yi/uv4oHqHc/FaLr15O2HE1ovsdhXbSduc8t
rbrmPZ+oX02fyrXcDql71YIUUOaH1dAUjOH1c0IYZk7TqnATPRiZOH+TdoL3iKsm
MRNgGc5suvmjmdxdLXX1GSCCMGMozlveIHLZlpKQkIezoHEb/HU2N2rGugJRe5B/
iiEjr/HJ72DjHnooe3U1jjHCTQ5Hv73tBNBR4TrnzLrDl0rkLt481iidHw3H9WZv
wSL/XHm7Lf81dqIuhZ5keNBxpCkOpwFkTTdNBgrxL5icOpYnYfUqwSof78O5YyEe
KeG7Qy2aRZprkQKK0MkMli9fBT1JGbv4TnZODeVQC0yk3zfLnp2UOmIYf6IAI+xj
5G/YZW1SqQm6+rRNELBk5aBBxnn7rpER5ea1bFM1js084547OHXQgvshxS51fLAe
t2qwn+J5SruOOMzxTtKOq4v3wMXkzsKxTrfx9EDqee4Z3XbKkzPSf7x/j5ZWwnPI
qgtIod6MUMrOKvBuTUDTTfsiM3Mz2BlOfkKMVe6qs9kjJ36DnZCdVkr5TVBZFjE7
5yzwc8mgGmWwgCpaH2BZRqIvZ4B/zILjXG4fEdGALHinmmFAGczXuNE4SVwxxqcd
NNhXeJg5p8g0rSRYczjQRLwjzO2xC5Yz3NF+Cag/w2iDfgL2LN4Q7Cxfp8crVb3p
MeVytoBwsiGRaw9HgrMHJUUm5LmqX2xqOWXgkvcMb7sOSm9Ij/+m/gPi34fYSWvp
UM5wx6Z5onScV7IK2OjsLUrS5zf9kjKFZ6XDN5bAzqrVQA/syLUGFo12ZFtL+tJR
FHVbdld01QUlk24uwbBgE+jJL6riWvcJ87qJAVKuQyPclaKqd3b5x/+hQV2DCOs7
hiCwTBVIvkN0zceKIx7gsSrAj2B5rXgo72vMwbuSh5e9U8hjR/mVP5ieVkg4R8v/
EJlZPw+OcNr12nP4swefXYS9PZLYoc4e921jvAUb5D+3G6p9rRjal3ZHms1DHPY4
dj/oc00H7e0MwrER18psfRVQo/vJG0cluuyxWMruNXCqYyV6c9SN6mETZvbKaR+p
cxo7GSqQp4UBk/UK1CulLp/6tDgIQWNDcpxKAfbMK0wm9/6c+I2igfw6Cf1dwpCM
YToPOywVJqa+CDh6KcJoagzca/mwTCVKa2BW528oCQeMzhZ5vjEVx8wjSzoP/+kl
WRvQoJoO6b16QFa+TIw5bWzHojTp257D2XDXU3EIRrF1Qq1ATjcXiptmdxPXOtOo
0whfm/dQUL6xclQ/On8V8ZOPHfTE3WNwxj+wd0arRFOo0aqzZKgHoo5QotORgfE0
6kkg8F5/tjHBMKmdNMjmIdtmfCvQwT4OC6WRaUqA+Gi82RyD9034ipBu0Bhm0sxr
YzCcFywvnYEXAjGa5SY0gYZm97rPKRLiUpHq+hiIxrod6atjkzAFY47319gefI/w
iHGxbrWGpoSTYtZTHpMlFlbUZpHP5D6x3TKI+k3lwJekNlVmkoiApyM9H83CZsLu
wMH8CkJ61KWUGb/cq6+sNha0ZTf71H5R0WEpylZ5HAJBV1G3DkaZD5KOMcXt9Ith
KudaRTWP2BCAoAh+pHIoCE/FxGmi5lLCX2EMNvlNSmX2HlVlQs/LDfTCkbYH9TIO
a5o3JGl5D7MYpNBcMDtAW6xide+le1ucO+R0eaDkKdXjKYv2cjWJAo29IZZSuDfW
t+8+CX/UPX4Ry9t/IzkHM+yYTHEQMJZOoXTQZYCRG2ZUx9xqgu9YGe0mWeJn0RvM
cpv66xS2SG6XdmYRC6AumHNjUTGnqn3XgvPLkqSs8FtgybuHS5pe1/VI2oiuYk+W
VqZu3L/GOyz5qZoDo19Oq6SaPws30gBY+LuFQP2L/UrXxYmtypE5t7WUeVx+9B29
qO1dVwdaiPduixNLYsFxMJbaIS32IprtjGbnqnHV0X4I9ahLgjrU0BJ6rn1abNNK
ftbX4PlStELOnVdaCgN0ki48x3SqCHATx/WKZ0fNZaG95h4jvOxKVgg8AAIErib5
guvW5RPdYtiDvae9JeN99naG2GYX/dYLYcvzBXBc7UV7VvVRJSlJiOOE9muyGrqW
LnwbmVptvFakZt//aO5ArzxNiHUyIFxR45398c6dXgJxNv3zFE/v0HbyQW/ugZ/i
qDpiKsS1jueRPfQ7ivHDFVroMFtFHoXnlxijdx0xdGern2vDEDbtnzDVzDwPuuQ9
bQ/S91f+zYlnxyfnDVHUjk+Nj/9c9k2eafmObKXedf/DOXzCDtMGERCiy6gWFIlq
MEIU4sOFcIc1tUi6oR+XZZNFXIJeLF3nOtZ9+FAi+SmS3lXZ9LkcAgArbNKyypNq
m3UIlSmdW4Rw/UcGiY4N1blysKw5NYPf/QrkWi5/rhySVwixRFEOvm+JDa8xiwtD
CgnjmjdcNWXODt5BGUY47Tw95YLq9XVDOIttae10aO7cY3JTu8eQ+KmXE3l+fNlq
o2kOm902YEZyB3Pn6I69JZ8u/WyOabCQxaP9mUssRhiVWFyrl86UF8brf9OonfXb
Z8qoIEnaYEDHkIES+1G03HsMyjG3MeSA9ZmuSyotGyt8rSuB/wem6nMAMlZo4ZsK
MQ++hWHLtnL45Oa1WlK4FjEKkOglz2vRbiv1h5jmD11HMmxSB/34K8sTnVmTkH9L
H+TGnqYkSffBn2GDmRUgJENXQbDqRSgUyQv1Vfc2J0mbtiPL35vbomirrIXRHfoy
77H9cRyEqd4unaHy4G2YY6SrzBDIMNRAPhT6d9B/VFmMVyTO6JqKecYwE20B7uq8
40fUYB7w2F9643N3kA0EaoW3qGkxPvav9RFu6PfGXQEtnNj+0VIDtSf1Cz20ni7E
k8d2msXbmJkncxK15oESywfQFyfemJ7fls9Q5o+44Z5bTiluY1s0QtfYA67wd1j0
hmocLGEE7O0w+MnbMfRyWDQlwXxSFLa8SpMnK57P4Um8r1tiyHfg4wmFe8M8wiz7
IPtCWgLKzP55y6KuVRsJXrDfBwk3SUy1DI6GC1dtnziqqj/PrFjPvZ27mDdCKgby
FAA9KbbH12ksdVVEGikAbB7aYkmDc1/C8FixSsYMzeZ+pFROwHRtHjQCPBw+hqbk
y6s9BL2pYUVT7SuOSTeF2bHBf/l6GnjPsJMFu/FEcrVcJlPPdW3QjzAwBLwhnZCu
T/FKa6S9i9ySwWObPiHxKmZuScY/2HABpA4j935BNsmdNNXP82rzsGhE0rqIAjDN
/mBhoa5ZjyzPhIZ2LeQKFybtJaybzxlB50nmALOXY35EUIi5ZxxxOWbfBG9CfBCk
pZJ0Nc357FkKjXecaysbAnfs2Bhh7aSofgsKk0EvBcYebxemJKr3IEkj2FP0b3sE
Tc5JfY2t+8P6uYS1bcPjFjCXFy5MxI5fSnFZKP/khlS6FKI21afvPSEVdOeiqf12
rpdyNXLfMcFzYX3gKy8SoOMb59eNpQLbTYQ/OM3kXUrs1PCa3aLaO0P3SaoLWnHw
K73Is4wOPiiJNkCEsVmgAx+QTcBmVEo8glsIIoQ4absO4lNEDmDCUyv0hIgl4Ahb
Et5NnBCvGhX5PsdFksST1sSDt6ukENtfDD1VYWFhSaT9lpDDjJ1A6sKrBtDuiz7e
6y0zCY/kmSPXAAMGo0tFcg1QiZIu46wT5XyLTnjc8wek64z6mIkMc1KW9jxuRBB9
oiYaN/oolwXpd0MC/ReS8UOZywcjVY1giJpBrqZrdDhGAq9TA30GhM656x6lLlap
QwZcLht0+ln9Vp7KLQLsQjqDQv/jtRlH91EMqbbsXKSnfLUMmY11H2kfKM06+nk7
p3hT41eZj2h83gQGSzTfM0smlZsw9D7c569ycSCM9qfMCr+hF7LOSzuCrhQub3fh
P2e3nlZC0L1CTxHtlV4Xja9ipHvGrIoyN+bGSOaaDo7vwHZEeZtSOddNxGWacSRn
S0bF3xUQPf0Pz8LPDlLrSIVlfR596QA7MHPsHLN+G5wi2kacxRH1Z7+VyyQhRsxO
3Fm0Cb53FjSBXviRvgka5g2aHIjH93PLIauA/1Wwk8sDAbod3NKl7+J9jkCvQC8J
mUr44G2D8IN0Nwy5EbMFgx8J1ehG/7TbXEBUjjQsELQr4wcn63UZRaFU/LrLklyN
RZHE681fjvKVw1C2ZbVK7MVbg8Wrazyv9aw8ZudnC00gZ/bHiUWSCByjV20tt6Nl
PGb2B94PN0QXDvvfSDw0JK8cUxK24GJ7yK8NpZWqSp4FNCgMInk2T2eQcV1IigjF
343m0lHTtmC5MS6dYJO9440Tdm4RrtQjaNzYsSSAUXeM56ZI4x7w1mdJ2hYKlUT3
B/hCrfgU9lHe7pzjMXlndmrDRzYwSGthHBeDtMw2Ji1jRPhc4jknqoLf3Sv6wZHK
dB6brGdhwRGS6AOfjtg8L1wwKGDya03PxVtui0tkc8/2BPKTyxNoq7GxGcrQMz6q
7wRUtLahx3IJDpBTWdlW40X2oCp17nVgP/dqRj1jl9zuMApf0g9NIrofTFtZDJrT
xDdMKhsSq3+BR84foNcbWwER9tUN3aRo3U5T+pA8E79t0mXRwDAf1YdjJQ/sGxiy
4KK9V7NkvupFwUBbvlZRKi969rjnH5Zk3tMQ24vLY8yENFMCcqjBKmMuKkdDmfNx
1lBTozcDIH88p7DkO9TXr/tTMz+yJdI7M3KcNDx5FY9teOem54pkrlNWchJByas8
9IYt/HhSZ85y4H6gMO2g+qWobvkoDIbQTZWyUP7mkYvkPsR8No/ntl4DztbLH2Pr
WI85Yi5bkQ5Jrtp7uPK45XLeVPoO/j69pbksRvPg4T300OD+S6jj0gTQJyffSXnB
1dJlo9B0k4c+zPiQ6vvEkYwhdA0rG8Bm1QxfalTV21DN3Yjg0tSC3qGG0pK9qD47
Hhh19UCrbe932ti9lwuAozvrMGVD64eufF4J0IavGuW7dIbxqCsEb/KXNZOax4q6
HRHSy4SfUHLVTIbhgpmFrJDYnwV/PRv0BigS/LIVkbV97GFdlcj9pKMVCzneNZpP
UI9phvJrplNVgEToZyEK7WYFJlKIPN1pqmjDJxjlu4tfBnJpQ1YNUwCbmGs3bU7Y
vccrErn/EYcO6YRVtUX2sVg4gdJC3dbr3QmZCDL5eN/pxLKwFDLnKBgihb8S3rwe
TiY4tDFgGzJ2dLk4CpME9eIduNOwyMUgBTOqUADGfXTKz4UxldL2DRAECjjqRs4g
uvUm0e0MB49xvZjzrmSYS2vhXM7AXxKGTI7HFB4qpjfQ/DsuBgI7ok2tQDcQnQ6u
hFII1ZhXR4OsG328Qj+Eu+hf62OvHUqLYXpFEUOrkPryAUSwELhMYrhSdtUZfzZ4
ljepCpMmZH9bQfgSn3lQLfAqWOzlBOsw8E05ZQfdAtNDjq6n/2qp3Y2bX7COGNzP
KG2wfaeqXDZgNwJea1UuvbmkoXSbMgxTeN8MRdJFTS5PNUVTu6GPRUbnbxRECVun
eG6xVTnYe/XlRZnrlkbPD1phJthaAqXKmxdUypKBCehtbLLZ8Vk9HPawrqNdW7oh
6Rn3IVRIUuBh0JLJ5vijYNw61Gohq2LmBEB8xoT975YFLKrqbIyVJ41rT2PfpdRE
yDtxGWvnKibfxBE3zkO0zENlcyyIh8+jpfZVE2CQGoANK7R7C0Dhb7dEtBrjl+6v
58k7FC0Q5jD4khB3aqdRvaSM1eNkCpdpeu51k6lFGRc7imTd5vsvRRGwmToKwPp7
PYO2pGpZ1QI3FCwREkZHcZwu/sHV6naLJPAFafszHmrNv+KexXdcS/3ZjqlkSziI
1yMpmztV7ZwsstpRbDXJ0FcRQlrDhnxG0gLxXffLydWb2+rfuamFmX/iKbBJxMJe
dYb+Z4ofUGMu1LCnMuAktlmMMO4rQ35qwGrGGk7oQpIIUeYQTon35bsIIPji9xXl
oq0sQn5M0DSKdeMh1Qr43ZQC/mqCKt9yJcxNaBJ9VWRNIZkQCECZpTldC6YX4UuB
ccgxC8GTmCMbmpKLL0VUTkXapyxLUzTPkyDp7ET6On+i9MmpU0FaJ0tzdKpe7hD1
TroP5nSSieYjmnkbU+Lwzhh7A57z3Q0x6wsfndAv8SwQx+h3rwR/FUzrQ2qk+DV7
Y9DIBTK0ZfweIAc7JQSP5OgOOb/HL3mkL4dygMf3Te4m1hjT0dlTc3Kn7dnZsObh
BiTdnhX600uFLzlS1sft90dVXbczWf9fIGntv4G/vMATEObaw+MmiHhaimAruXfx
bGW9J/TeITA3caEjF5oxbmEkwCfsuDbs3zgjfQkH2YU99mY5Lun3qIWQETdnW5Nr
qnqUBzWfnXVKbjGcVhBnMoX/pSL8BwQutyiOJLtlGy8GCKPUp4+s97OVy69UJkL3
thv90lyhNK+5AgRnuQ2b7etRLTnwIAbb3wQOZEuwoYsPGTA/eNqYAobxbLEuFMyt
Am80Vq/6KM6C26vsxeMxDy+dH9/WbpJd7XW83UCCSEG2gUNcZHzS4MTPYT2mZ20Z
zoX4ClFHSPEDtdIIJ3PMEC3//OKtHyq6JGunUyUIn6Xc1MvmhxVWUWt0qXxyTiaS
xZ6FE30QrPHxRtSt66idppgg9HextmUHfH9csOIqisjnU5XhZI6HMwPt3/5rRolJ
bbzC4P/6g5gYdCyg/qGO6kBi0Ach7cYjN6geldZI+MhNXw6v8WYI5BcdhV9V487z
dxYerJP7C9qswc+90Q0yUIwW1+OEqn8FhSim0q71TGQBLRC9KN5UnxcKm9gDM2ej
N23YVjCCbh2DkMKMR1v9YYJSOScGW/SqpoDmVyJpaQ6iwGGaFoy90VCChAyTQcYQ
KQ5mz4bQBDJnlmWL82h1Jf50HNPJngIboxG50OqlFZaPRMUdes4r72dhYa0qN394
UgDpoh4FaNAtfRrFzRgBcX1we96Fn2Akw9ixW/ejIw6LgFVluB8GrIFjihdsSQE2
VW559/YA/bPT2wzjdnqwIVFgu/I8Awb8+064fIcYksnhLmZmISR8u1B31D66lGU8
Xzn1OQtGx3ZR48h6elQ7GvK0axSNf3NV/tmvMI2Tr22f6PCHgySrySG6JVgIRzE1
09LcT2lvk9AuYgUbltYvZ3u34rLpRUEkSeG3QYGg+6ZxAtq1zPFVii/SMsVW+hO9
Do/FAbBViqMtflrSSHAT7R52mRU1XpKvtFcDsDQ42ess03hZeWIad7dgV4SSQM7b
LZYlPLxcJxibvsYAOAxIUA1Pbm/TtHw9HA2JKvP9Hl1Q+6JP3CE5KV8fPOAMZD19
qddWNFjpMXR/IjiHWvLXfydOR9s8RDS8VAR/F+FXeVZOHgInS1+jYUStvZWYE9oV
C/lGxy6lLxhs0q/LfS7TH2WtcqMxqtETkjijSrR0kMOzcKk61tVy570/n9d+ORNc
OIwgVl2tiMgFlTalYyM5GeVlj5MEor/81ZMBY6XJV/Pgq41m551EpIFc589FvA4X
zXC/FECISmv54xEYKCeXQ7dFxHAaS9dQBL5aYZfT1H6pCsO7uoTWtfq4zSz1As+v
3zJvRlZwNZZ5LquYnuDD2FKXOQZcvTeo2zwX5i9wsu/DiZzP5LVCmjJBBgP87q3T
SmXGxqgUjRAxoyAcXlH4+9MK8V4lUWYqEVk3kore7GlzuCsa2h/S7JO9vRiaDZAn
roY2pOopmoxBKjzubbe+KQ==

`pragma protect end_protected
