// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Pz8WfIJRwZr7PNzkaJch1qrPR0wZnA6bPJnjuhbFN2SxRrZql2WgMBn8EEIz
PzEv6/+a34b71UZLnoyAuKDKua0RYmQit7x7LN7udlPyLGUuCez3hmeo9ag1
c/0ySZzkFEuJy4DydTE9N21d3iGa0dg+b4aXLoHyYnnYd3e5gfyr2KC9CZ1i
6e5zmZuGGbl5zbFlKbQBaZJpc5pHM0vCie5YRIUFjZhsN2tgA6GWO4sBMwMT
K6cmgrMPmQhkA4xXZoc10gr6htspVANQx5970iDEmnOz6t38xg7UOU2q56Ww
1fGQIhEsRnYi9JU9jvnAJ830oPNTBvwItsZSxE9LQw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
qC9NxV8eZxEbUWyIYPCqz9qBJv+FHctj/4tABei4Nh6Xpq/ryquXN0o47jfV
qhp9z8dhCt3819fD0pTarktb4nlM7GGm28K6BDrd1sU1dTgkasCDpYxgkh0X
c4sP7w3X940DHqDBMxfO3ETRme3PfqzcD+qYaafvbvrnjEU/KiSGH5SZZwcT
0DGLo+I3IQC6KZ5rOtqt8iAsbJsSaWQKpHPn13abm7GMM4AbL7dcRVjcn0cw
cwgSYfMtyAi16QkrUnmU0SZE+vVXwFU/xwnst/HFfs1fZVND2UkvGhf2uSu1
h2T56TByyoxULqYej+SexrdjnozxC0NHV3GRvQjb0A==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
My+hdH0mhmUAfdc+ApeQLOto/VS3OuXrgvTeGxvV/42g6icd++nNpe3M4XKq
e4aFyHph1Eme9j9eeW+TXyScD/qnSCD4djBZAnA+harbEmnh1mRzG8oCPkvu
n3GE4cxuuo1+A2MYk7aRFXxT73mBrzemYsP+1tEY1KCd0ymxQChpEiUkpxoL
kf1ghn1y8JN2BK748l0E7/WQajxIDLuaSczd4Ga8MQOF9ShFK6haR9u+7yDU
bSRbivvoLkP57RzSZyhTAhSZr49yT6wV5jtqAKIeCZNjPBSe5I+WlN07Hq17
pNy6rISXxVB+40igI7BanC6SUzTn1Nx4XD8b1RIqZw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
BN/bQiESEobFfdqSKV0LvTAvny/U+t5PmYou0eZicP4M5F2O47YktngngXyb
3nRT8O2DaHS4nQWoT2pMlApx5SiIc+45HXroAu4gVxY9Hl9mULcfp7nAli4p
V6MTLYhZ0gk7J2P2FCYD29rCsIJ7yljrllwBhDw7lGCmi1VWug4=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
pjqoNYf9QJVIg1OrdBgP6Mpa3XT8VA6qnRGZ+Fxle0o6vjIJs9LqOKwCOq7v
ETsl1GyytXN4TIk1vu1l2L3RIA7EC3ULPSRDIdDVFpZ0L29kCmW7NoQG6Nsm
NVx8/Qv9wGFGXYBUpxMcNF4x4s70i42SCRDkwtBJUg6ANobxKwqVIQU9vcyz
x9L82KXv5VFRPnzV0ej64+3VrtVmE6lqwAUYg1Xt8f177RVCHVpOI10oYRjl
miL0xxXzTIdBjvxI3srIgy1NpY2aW4vXHacKf+MJrBWxw81n4I7KQ5OvDWLF
RK9xn7ROXzGqgTIuXuDTjBr6iwS6I4OG0tiGJ1CCyRGkLHzhNiRtoO1I05/U
zwA4ay0XDSnzRPFT5NfHwkQK8UxkeIDZ2L1ohgBXu19B4LaGcR8R+W9Af5+Z
0sEMieLxgKPEviGDwoT0rKS8VA1lp8Bswm3gTJKGfPeMmoE06tC7k6TRfNbY
eO9MqXpap4XkrNh4S0/XblPY6H1X4TCU


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
sZTUfcfL3Xo0RY1ApWlB/aWWJ4st76JXTKavWErJAluOaVQfcgHWkbkpZET3
1lXOPFVIzGV0/EK8jIyr+g0BfCAZKQ8v2GM2D0NguQy3uR1ShSqGCtv/UPQ1
0mW7LJHDJ1In4BMnUUtd1ARfO1Ix9gJITylrNOA6pbUvYUANEJI=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
hkMIX9DY87sVgpLTSEbrdzxMmGF/0luaNZBbSJZedQVb46WT1PqUC6OT+QTh
tjrePgkO1Y95AFD33H5YmCDNaNyzg545gDwDjjxc544tqUyAbk4sMNbLTsK/
6PwGdgWQ8FCZs8bjKlPbi3srE0L+VX6YENStWTSL08x/aSdPtAQ=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 80544)
`pragma protect data_block
ShKSBJiQFlnobHKEMAZr0IBLoMY+S5K44CjlhaDBIaif7hWOaBUhxswWp2Gz
NkTQ0w0Pn1GUo2Jt7tWxSAAVpiXwVAPKG9tOHYcrzHtDjJg+uSV0kNrhyecK
fMbKEWxqobEqQTSFPibirWZpAegQA0D/0MVNdHPSKQnKQ3cF1rfT4LFVHwXU
aagHdB6EBnVjmdT1zVn2s0IiRii0OvIVy9ROxOhrpq4BIs/uZn8uhIDhf/Yd
Uael5z5pkBHy20Dtf3iUO33ylMtLwESB35SkgmouQujrpkk73u87lbYIvK02
8tP3krptaeqO/VDBqXcuziWsz3PdkxdbM3/vhJeoaNvG8t5c3gt0QXXHL7Zd
6dG0RNrqaTKLuRIEbz4kay7p/NLOyXrdTjf/mpuBN4oVT9PEv0475LdlsqAI
iq9PZQl7UNmIfgpVP+Y7bUEq33mwnaEuF6OKlvsmN2UCRVNFMz2Gja0hpILq
KifPbS5IL3DO77calQE/rJNYGgyhuP1kGpNiJUjGQKrq2AscInWcd+gowHAt
APhS33fGMNVeNVhkdsqLEo/6kPzjd78fXtDpyQcD/yn68LD6UXS/OEV1lTfb
EYiAnMcysVB+3TJUjkM65xTyRylYG2vAILZ948YFhbyIm6Ym995t5p+lUGaA
D2vA14gZ5GCtbw1yB68Ha0OkuD2YeC8dtu6bkDCamiuoGepvi/j3VhmttZ5h
jjLo7PF/zx40EZaco3K39AZzMilsqcnfU9hBpcYuAJZhL/oEpK1T6qG+XX88
6m0JGAByKXg9IkjY3s110tdC0JfTiA5ChOshO6LdAlNQE5+8PIyesjG/Ybe9
7BSMLj8xaqtB+hmSHfeSzA3tvilnSB6RHBVV8MCZrlD395UgHSJcHBqDhhe7
Ln9fK/lvSMzOSaYIXrK0AjC8YfdXXdo+cqAGtMCH7rnHPnoscNujhlUMViai
fh/0Sm4/9PujWfzrdjPwcxWtJ8VO4bhdB+sYsbigx6SizG7BKX1DPa5Y22fs
JGSWmm+SIxnkZgyy8To0LCGCnWM6zWcUA6Y5T7ZsiLcRRWqgaSSsLL/uVEQq
s2uCrgXvA4ALavvdn/JTAU0BeZvlgsXFA1k7y77L/cdXBwsCxVnCHGg2ZI90
L2LrxjbuXMVQ99jOLOpmiLsB6sVtKcetJMy9HNemxI39Ovj8z3Xsvq8l288o
P/Z6pr2fhCg7nnmynEBpwKK7fb6ODZJMWnnfJqu1NyuW0lzjfseNlQxfi4ae
TEF0MhXQLagIox0aEmdCVpdVVbtITZ6J/eZ383JfLzxEDdhPxIAvxIv6MWy+
UOvePIqNf+zQp72hxsz2isOSuHLmxexNl/ra9z70HBQQPFeUKUbZyyto+BI6
bjbm4tGoHW/9LIYiNW3YP5hnVr5kvSxX7bip7Bgdf2ySyUAdCoYwPlVFzor5
3+LTFmvskN7whniLzjNWsnsE0rAyOI52Q489JqTqhDjsxzc4mh3Isr4h2WHh
NkB2APoTTIe8R705/OgyNH5qoR+HFdhStAHNItd1gGp0BVfXspNnYf7+Q7gV
LxiuOWC0gpJ/WC/iCyL13ymFbQ+ipT2M/TxBTUv95gUo+KG9zHo9itVOeUqh
XxvDZNf8/77X0QcT4v2ExE2VpAMLH/NfAiOXXk9TkUwjtEOUNU/vEE4tdPNs
CW27eTtxYKdaiGnI4pKZhwtqgUaewMujCLvrB9sDnl+ObV6FBaNRqZ/ybS5A
dbG2Pb1EzogOqxrxpIZuRs4TJwlMYg2xSdp6+12BI6ZKluo/yoQ22Rj8sXmf
NZFBWV6ooiqi3bGNX2xeMa0pT9ZFe9KEokOJc5Ksx3LPnPZmdJgPSL/4JYaC
6Wrm9yo1PmHNvgVTy24QscTuWCAAMLBTTXqyUu9xJ4PLPkNBkwAS6J8XBmlt
s2r8lpYS6eA8ktqcNrev1PzHZy72yinu36scpRG6nIGxQuW8JXVDw3Zuo0Ms
anB0AOgEV98sKAK5uSiY+XNr00dUaijZi+s+5D3DedfXY6NPKK+b3tjYLqDv
5sNd0ZSSrEICG/nj8nZpST3I1+z1j/X/u4YyKvA8nV9zgQLu8VVI2FqaCmTG
mln8vYG5g/0gzAzIGLtrD0FhGxyJU5y8vrk+PfbbmwELpjRwkGFVjVst1Pkg
KI8/G/t3u9vzTLRPcs2ZoCCaek0K1RQoOI0IPK42qM3bkLPjjKahzlBqak0f
rHTj5g1hLYlCZY6Cj6ShMo/CwnN2WcQFGvIdFAYN1TAvbrDOCvXU4/sTFIkY
JRPZDh4fes5Hm/VbPOs6wjC8SnBiAAXWhRmhC1hZlwYcQyQ84WYzcHs0Cx/w
hlXOPE4ZRY2ocz+Feq4m0BfA9aWRREOAAT24/f6WAUCp5rujmofClr2GArMv
FEwh4BwU2+sdPoLXRdZeo6OMPRbqMaCDsylh82IZIyh5zUwrV3Mv27hdEvx5
KsSSw1rXN9AR1iqnZhmvJ8PqHGO7GsA9kVLUAbOr6PjdgGJ6PG3dx0XDRn30
gvkTqnSIM6xvjdxdHWUO5czzZkxjkOREmyzvytr9+YZCX+m5rkMT0jwiQai8
Xgc0iP4cd3n+pOPhAgB8Z5zRzwCtabTqWPq0ng1XrBpStqNxcoHzBc+gOd6K
WtDVG0Yn26rSBxZTPpNnim/BsbDaLrmMJPcYAW5EijBuR9onH73gRW9aczSk
gW1vHOK2V4R0ZNNSSYn2c1nAo15tMJhwe5gujvlCUZzDUHAjikT+07jkb0Xn
/HMHg0WvwEUfz22P0/xtEXsBSLj4l4s+aUSkXdOcLPcXYiIpC2cI7BmWfvLC
5aVTjNkmk/AY4aX58e/n36m0kz2YJoAlJgv4ifYsiwfDyP4b4qBnD3jeMDGK
HnK/Lmjl7HRuauODyzdm1f+R+Tyg4Q2zaiFigDxrjjq/YHfMph32dwqLSem5
eOI9Y5JvcA1rrdSKqDanirgWvzQ0tYp3hX6/8jkblBcx8RLpsG/2FbsH4mk9
JGZ4k6ZgOh7cnugYrP7OldFOf+WIrpCRobcFaPzWJarOPiGSaH0qpC0alhnc
CKOhChWVXMB3c1f7X4hpbRmOKZE+AuPjojZkanoR0FaSWxspBhkZdlE/aGbC
1kkpjEE0ySXfKRLZE4bI0sOiTwMxlaLvlu45VUZZkMAMzYddaY1/DCV2Fqd+
BeJXhTiXRrUIddfAc/FQeUUoMvwgSEtEYs3bsPAmIigp21FM9epemv5Rzlk3
gXZ/g2a6oJgpuXktp68eMfS4/ehlt0ZtVaqjF4CQPjHotXS9/m644RHUR3OO
Ix/9LbCA+ZjS+PTTAckzDNIij0ARGna+RTkCbMWmZhpIULJlBKCu+XNmA1K+
OtA9AsG2RafXOhFUNoWrrZn6ZfDTOQmXl2NBOSD4GKPELfsPtJ8p9wQ8LJNE
JN88hyIBypKg0+hRZicabXB7XgZNw1Mr5SCw5+xEOnzGoqlAdgxfE1XSw7kQ
jLsnNEMUmnvchRiDrGWOMEfVAlH3XzqpLWrKOAyAcsPTbFQJOiunLH0Kqeoa
4DvcVtNRo23BRU7VO9f7cCny4NV//Fvch4lk7Js6aCo8Cb3IkwD6CCQZlRXB
H4zE6uiR8r+LmuzTjnW8cGgNM2eCR7+TbG/a1y8ft/hhxbybEuWTY19oOj4c
5KgzorcFDBDcW53u8sU2p4eaFzjv99idhXSmDirk6tK42Y2yW6f1vcQ3KYk1
KnsYfSRNn3pR+3+epIWp938913tC3mcSn/tIJALFsa8JBhITLGmEKtVktR4P
fJFzkZXNG+CWscx7c4VkcGEzLYzX3p0JiC2hkrjKOCU1TZ1dAOCy6dYOlldq
igiStFAa4eVNlKM/xfG6REkdR8omSspTJhs/TEHxDMrVtXDt7S5ZHffpEUAG
pgm7/y3rZSIZwRGOSc3tBUU2pFcfXt8rfBbqZOZltDPyMCJBbG9Yx1fmsPeg
PmR7GI8xd4BnN2dj1DPDjoBWVpFpDigGlfjv7LPx/NZcXDDbUlLvkXZz6/kF
kwSKsfPPHRILoQqcGkSTTUGU6wDbLzbNClaVP3NUCDn5gEgGaNzaJam/+/KJ
N6nbDJV9R3pkmaEcGlomxsg3ZpsDa0a3t4PV4iuo5ClgT3NFUbWhcAqKueAL
4UKp+abD/oyvcjwIrsxHtYygaWr2vYA1TYij7JQNAruJIQTVLcRxLhQhkJtH
8gspG6pWQwj+NsrnivpA4dQddpOh8LkI2t0JLbRxdng1kpaYOzo5XD3ay434
OoyDeXtWuTG1aGGQgsVWyJiXo2qu2tiU1OvBXWQRuYUmPDryVVXg7DCCWt3D
ZUS9Il6nYJdV5wqA6FIbJzcZmDBhmIAZrl+2qp3EmpwSWTwbFjoD5MfpEveF
8muOXVgMg+i39lKz3fQ6ZHzXWif+vrxIrtuOTwrvJF3evweanf3o279xHFxm
RaDXTjDm7NX6hypOmV5i8pDenO8DgRwMOHtKXKRyt4lIf74uJxt+bBOGEHt2
XobuyYkMXt0haRGiQHl0rXw1l6DUWZmmLRvZ2vzx1U286do/r7Y/UbEN9OmB
0ZR+8npGS38CRDjImeBQRtlVsU70X3lHq1IDQnibQKaiNXYlMabozFFQTQwY
vnHQaw27KtbD8Jy/6+S/T12ZyRCE0fp9PYum41gjaYXZp+1hPdWT8Wx8N1ii
R2apUmmHJ7wEsC5p8LFPTCPWr1OlkZfEx2ADw8tGP0uSA3dhWkKUWPUhyVqw
bclrMqtAu+1YKulCgiYYPywRYZuvw/2IingQQpx2iJAC+FT+pz0lwWXyeYSp
iUPt1FKs2oOYJeHHe62It4y2VsSAHRgeABfKFoceTyxJvpHNG+MC5LnGc4ap
XCqWVxIgbSd/i7dtAZUe2Uz5sJQt7XgDfAeiLK2Dff0jZJExpnHyFYXy7Gc2
kclX/6YVu4YtWrzyBd410/yWQCNGwCH2WWC6mVMPkwCOvaJgqXlOyYUVfepx
Y7qg4xx/MqdqGo/4EDNdHgWVcg62vAfKUO+0ufSIXTxOvifE54iID3nbGf3n
LKOGRE7+jZRgTX6Ecefb+I/LIHO8HFhos0WeRe8BpTxNo8HcAMn5YjGx8Ykx
fara7+bvKk7hEdl0hWVF4dBgVJUdoxTMHgi64wGLd5egAs3oVw5o91jHemac
ypTB081J1KqzwONno59NGoS12h6qJ1Jg6hEWjd5ZghxGJoHYC+ngIj1CJ5Zc
OVNotq010/e/Pjp1AxUt1el+NFusS3sF17Crfyj4CkrmnEtjp6zjKgeVTNtV
XNaSknlRgcYiZ9pKa4A40lhr3FIS7CD4MDWUWIBVg2kCP+oytD9+9Hf++EGp
OKpBDNSgry6DDdJwkceRvpR8dcK9RvxcYbjvMBfzgFD5/MIi1/56No3RgAFh
IenGYZXJ5hBYq4rUX/hkS1q4RpH7WW8UDzizlfuM1z4xfMhoMUplZ3qoh+a9
o0KVETyuvLspNkSYkep919zcG9higNHk0aiw3Y7znvMwQzFiLIgewiDN6hwP
9tHO7864s0ZzjtYDdnQ+LVP+jSTNnqh+lUibiePv2VTNoFmv+yWB6Tsky00S
soUY2FCIL0dhBoTx4iZohSUX+ElykpC+fpcBIEDgY6R6eBKFLz2tqfEJ+4Go
0dhjK8/POrwJ9mbRZDHFeSRGn1lwnNo7p+uXCcCyN9C4D6YJ3+T61dKWw6Wn
hPMqsR/YSThbcVWX/MTnhjI9XH2LMhmKF2m5VWylc624Z87oia7btTDOw4dD
NF4kGPANgzNms6ZNdwSG+mL3dgmrojVtQfdHX/6CuWkWFFFGRCOOG+qwra0p
8Wu3v9+Wga55lal8rskTImiNEuErWUOJiOddvYDxr4HyS3kl5/O2yMjvz9lA
FpUf0R9o0EqPHA52s4CNmXqEOsDUydRro/6W5JDybo8I8wbCen8J+FPcTEcc
H0cpYfrkpPVgIs+/sff2sh4U9+aTTgmAoETD394gTNCw95y12CQlhR0NL+iv
LwXcbFj3CbjSaldSl0pWSFQXkn2RrOCMLJzi6FKG887QGCj7n1q9wydiOPNu
M6/83OkhmoUmtnwLNO9nVocVkzJ7h0AE/6SYILdlU7zabqL4AhU5fB6h31H0
FfsZ4J7y+W1f9vpMSFxZv1ZqC5KXs4VDSXYnL3rLaBxzx35oHI3NU+EaJa6a
Q/E9Lw5ogRYIBmBFvBGlhK9yPvdf1c5LKDxgcIH0FXsgUGuq+z+i56y+Uvp8
92YrIY6EA3g4ztviAi/jKx+aVDoOdVDXcVhD5RmiHclxq8oOqZMSOF7O6dsV
f5gtJCcLHs+9BOgbaKUEDuZ5/9e1Lz9IkAlsXe4pLDHp7RGlxFsIAC4AgqRV
DYrMm/7ohIEUWmcTRvAAX6trYU50RjB6v+v61qyV09yOyKNSGwtKAfWtxcm0
MJfgQkKH6pnXBX6frxB8u7/XXdfG9l31cMTlRNfPICfL4Lf1l4m2y71gtpF/
s43rB409MQzY87XLUb4jBAuEJrFHZAZiyNAzSv0UXvezo3BzoOIzoH0lh/0v
ygN5O71kSYPVS+TxyPdyFaTtiedkl6QSBACC4t6ZTH5lGsKFVNvyooUuYYRB
88mZo+NNt3zq/3GHQW7yYJXneytO3ppRoKhebSSFBuRkRCDur1nyF03CrTna
vc2QuFI10CGdWCDqUszVyHopmBua3bxOufi6DdCA0ydiuorS+jHDbmSTynBV
dPK0hOXvi45mnrhRzHVTOUB81XRJfrCc5O5ms3ti3axljY6y6+vcwM9U8kcY
Q134IcvBQQkB1iiF8NTpcQxmlo36sgFgfDr+10F85P5z3RSJIWFWPyMiVblC
mF5rbNV4JGXBQkwL92ZyK6ITmvNL/UKKdPBhWxdj6gDZOb8mhBiNnJPePxsH
nOmbqnKiSlqZEdf9w4bN1UNnkHJ2fitF7ISkvDsSJ0fQGm+1QJZ/SWhyBtbY
bB4wjkCflRsTPGYBMRC3KcKawp+8S6v5rbRCfKbqzL40CDKKrUEoJNnIZjut
9kUoszBUJcJ4I7P9Iwl9f46V9+stpIz572aj80FRkbcLPuwNUBb1/fBWb8Qq
liriY+pyWMXHs37BkNNpxolUg9m5y4tCJmgH2YvVdJbliC8aR95Ai3Ckr11i
9SBsxv/6KnDp5voFTKdSiwunDDbtSuoJwEU0nmrg7ybBMCUC5SqL2IGSIUQG
v8GzI2Yjte2bUWl6pxRlpObCGgM2RTILVBB1NriIF73WkWx797aLHFVO8mqd
Qwzl9GXWQsddUIg+v4V2B5k5CvXzzqmQ09TZMjGNgDjbvPVYQB+7tZ3/Tkwd
8DHhSST44hUaG7UmLCDsNYVNxG9G2TZdfcKtcDOv3KeW50n/CB0IWmuxCpYg
X5itlTEE4yDqKB8UvZV8Y5LRCdoigsSjN1lbd8PaScdTkSdhX2xB5aJju0G8
5OubzxZR+GKrliyJpTDryufmx3Z3FmoqfAcIomsTdEVW1uhRt315hEkgb6kt
xnyNKlowAybbo4bqg0/yI3LEg65fxRODBr7b3MqkU2iNATHMlgvCYAJ9y4lB
Xk8eN7LPgUHRmlJsOBjpcB2ixnhBn7gSAmc3jB6iX2W6UAKyDYPnhn2U6jAx
LeBj7YpMZ0LoHm9BDn0MZzEQB6mM1+nmo0TrlwcfoKA0UjS3XTvAq9SusGZ6
IW6FQ23zmisbnY/7iGCbkjgzSTVq+7bkMnt3XMlbweG7tzpBkidR+VMZy5uA
M70mL40z2Ks8FzgEcI/aqNLPq4pjarqi/rybZPt6CFyu2/JbXzrXbnqg+tOe
9D6EMJctTAuwl8nAhX5PLEUPKdUZqouZOfwN9+PKJ3UDpXFyZpFKI8EQ/T8w
HPT5CZ+FpHWAB4yb+QL10FWB0iyn4kKozUDZvgmaRpaj2d8QC7tuF4JcH9DS
Vh26MJKOmnQLpn7fGZjjOMyPiUbowX6grISSyXIHykDVEu508weEz718sWsv
WL0t6GxuuEnqLSAnSeU5z+qmwn1EhjeOgoqpuNKNQ/PwF+QTZBtQcZ3MxMbZ
nXGrTXJ04sZ7gPpAG68h5ycRNqOZpqSRqZ5d4UeL4KdwRYzHmEch1/VCbb2c
sl0WAGLefHwwFm5g16n3V2rIpyr9r6DNW6zjRgefqbASapSYfYhZtazaDOPB
aIy/+WsrdPNSCKa0lXArQebtAXnNu6EVUNUbl9pjOMBojc1KN7qbhIEGQNnA
z8xaCKYJcYdxG/WXPmpWJmaR9m243J3Ihpj4mn5zQ2kXyvV+S+GjN0F8D3ow
awPRe8pLpVOJfXORoBlQ8UPWSOPAkFm6S09A+JIwAgStO5fsr6TfVrtZ+4Mw
yxq696IYr3y+xEKxEK985bxZ6e56JCqTPShMvQrQoUDl2YeToKbOD+4jwSjo
sI1yMPDX0vbwE8P4untvppVHoLEtpcmmIXd3+HMIbopoczYYOuYwsuRFEUb7
D05EQh9nMWTmuqvYAu65RJdvpOBifKwN8zyvhjMp/JVAtPD0l/0fsY68XJ7q
lNloHJMRna84QEexHp/k6dSUYSA2hYxe0avqwdNsnWlPUIM0HsEQN9FpZDJu
l3ToX5VOfcFZKqkY0keBj9/UIZAn8XttkiMWBzYl9TaIuw4oV/+FGwP+Ozi+
TpoCu58138O0dqmzUMVKYrfgbWMI1oL5P3GJDGGYvTKoHzGd15AFnsjqLjnU
55eAmL61lnpeD1wQ9Kfzi40kZYHNRQGHUTcrWdVw3HGdh+xwTI/gWrSpiitT
6CgWy1VrXYEMNflWnx3C/TBlov/biHO3f3ZM1zt5249S4KMVxJRE0sEBn8TU
XXbkq/mojH4f35GXQfP/ACQo0c0nQoIEqYmEKYjwifaa2AN1IIttfBQc5LmF
f1WrAlolnzpZxNbQdWWFq2kDN1oOA9S/RdbroAYkbjJSOYIit3w/LELC+kgv
Neres6OI4Jtzvt1z0cReQwz3LG+lHVXd3v2CPbDe0dscS4NQ5ObMt8Wgq3K+
lfceTjG87fmF9w9HRT2/Kg2KO8CtCMRKUPNLAhJuHLHF4kj6v1FoMTM52t4E
fH3WPkw0+y3P4Bj2aRf8NBb4Nx54/VurK51Qxq6bnBRrdvC+6KFDpaAhtqAN
87pIWEEScE9wurRHhGXycVi5Kq/7KUJTy1AO0fGGkhRyKjy9qdCOQJ5te9A8
tKgJc3d5huGvNPfTP0Uehu7rBG5CQjIQJhN1nBjy8gwJACU0wNJpTDN79lVE
LQMQYLT4ocM9I36smvDaf5jhaOyXZo0juiNWkGHclpsj2vAX7SHjBoUJvgP+
POAfKYEWOR6Spq4+EVYp4OTfPZUtHppxXlUZhgMlgbM/eTWbonvENzXEQhpa
4zlFrS56v7U0D8WikW+438XrzK4v1K3HfOF/al9FE+agoVq6Vi4dRrOPBI9A
IQDNG1a8/aKkxa+GVZwt9xvyGlTnvbrM99bhzMGmoZt73QzobUyGxBYdcWin
X6PxwEj4YpEuT1jLDr3MkE2ZAWazGghkeeEIhHfq/9zFNZtDxjSmgqVZ+hBn
bgjiNyxrEcbhpX7VdAI5RASy7/avqb02PWS8eurN5bEinlGEqBr+SSRHw+vS
VhOPK4PUa6766pQ8G9VEu2s6bFamYsLtbSpvD/G8d/nokB760Uz5S7cQyDR0
NI7eg0a/Jue9vMVd5G7dufnup15Dw/KRrKArzZ8iO6JC8hrEY7wlLFYlDepI
CrPmuNCOSRhusYSMbuIsBODEFOxPSRlklt2X2zywZJJVbrIBu0v+xTdl6emf
GVqC7uU5hwPYnmGAVWLDo0hWQhb5etJ7Sd+FBUTbq5WqNN1HGahd8ztJL5Mr
tF+cXDOsbyATlCIrW0O80x8uj70Xde1E+mqr3dxCRcNsQrffS23kuiNbfuvg
/ToqHRR5cv6hq3SR/xcDRN8ScaGC5q7quSscYpsZzC4XbOk/xkeQXW/9fRCk
46mJKqLM5IbUMcmJOEFj+TQd4sbg8nQ3YfGrKgiOnuH29iR5Bd9VF9dCUjNR
SjgKvFF+HuWedmv50qSmG266mnG34cd3E/3YrRpj9QZhWVB6Aco0KiL54DxD
Q26Buoqz72/g5CkJc6nuV8/28xG1WnW0yo+zuPoEWx55UdytSBpquX7ZjBEG
odjihRThzZb/aLVaJetU7NQqntZ3RDQYYUTZtb0EinX081cEXJXQv+pM0IRt
ulvkGgWSQY1LdlYur9U2AZyoeFEoAXV5uWM/K2TyKzgBv90h0bMEjCC/8ZQq
5rMfIwzD42wJreNiUghkV9qawIS9XOHlH6tUglfLNpnh61hRv02XaKZduKTH
rWdQTbGbSsOx0C4kMSM7uXCdnPLrV4l63N2EHUFFqd79fRhupxoccw8stZvV
za4pUOnbsafYGae/Fz/U9G1fyIOEwO+8B6Ae9rjvLjddKHV1M0eae3G1TETN
A89CKs5UYG6ycm7ARt7F9JmZUd0zqULRoHTZ9laPxIjF7BahzGZWun2i8xsy
41zC3HthG2+o80IZ+s35qGQ/IWHZAajlxS/TNH09g/JH7lQWUIfTye5eRaBR
b0tn6QZhmzO3HP0+7dAsTAHZQwZPneZaXe7SssG9nepK5gKbFR0M6yudZRth
xd5+l9EJGajIy/68FaLpojEoybjh430tLrt9G8dWq22Jj61RGv5pOlSxZRiE
kt/KaAKCNNpP5TQMxaFk1G0pk+YpDSEAkMCJUgzZFYM4TD0GIzMf/V61MxZo
feRW6Q6F5UpZlQ1aTBth+TeDePVIMPbNmd0cn3udYEAZXwmBa9Afus7dMEr8
7TN5QhWfhqW8zvfnZ9yM/qF3MAgf/tYtUz5OBs+pnw8lS30CZoJAHNX5fRan
Ub7szgSRutE5KC9/f9i6sl7JuBx++cs1o49dXzwPkMCOgIfjHg++wJFuII1N
ZmVVoIWhZ6NNpKJ1pGKsdRVzHI8cOk/iTK0LpOHmhs5qPThePH+4B8JoX1ed
ghsIeNRtq7gsTmcEdMbmwpcV6Q5wFQbYbbUUUv7Nn1fT0RgWtm6Ntici61t5
AMHd1r/A9oCi8caLtglxTJ88wnHAa5t20PxIygULeTz261cZaj1iHlaOA1k6
dXfXPDzESHNRLgG+TnpxPzxYdy5/TdAyOf8rJaZtKfQzz8B2ZsQoYkLXc2kt
0HVB+UDlBamw9fOthPgu7XJcSW6bZWRNUpZrpGKPlem7wiZbWWU0xjNAUBAI
w4gHvwKYlv27SHgu3XPufeIUHJiBUIIfn7N0mQ5j6SP8LGJcFG3YvgATP9GV
Z80C2e7SHmiijZahwi/0+UguK1NVYUN8XRkrcWP91QVkJXNfjSVJNNXhLqCr
upelvB3wQfqMPHxhPZ57sxg1pdhSw8k+BUAdzwpLNvy2HiBV8v8OHb4kprj9
CKKYc2+1HUg1MdPxU18N/nFKjVWrxUqW2uljZzBajcdgyf6/r5QEEEFBH0Oc
MFrlMtB55kHEzwUHu74WEf2TQ9XOOEa7EYm69prX4c24UJyyWcAL2IriU5qr
+ZQnyca+dQxagce+EasGgh4owHQVv5LNkfCTj+6RrG2kULC5pbPT5d9WWaYl
j+Vl0q50rn1gckYT/+8Dj6kLbP0WnmYywLyyIhCHLxi67Tq7kaRo/ay+k1Ty
uiDl0KNvgjVQGiF5Iz2qgDcxTHTIfhgwr+qzmlpgEfp+hhU94CYeOQPeHcKP
ro4pH5ozCzdJu45b9lzDHC8GkL+tDUZZpTvwQsQKKA6wRvWeZKIr7wnpcMwd
CByh5cwhafmf1pXsHqHt+TbxlwKGJDZoFuoIKcQn5FGDJBR4EmGRbEfZ/5yC
idFYTSZNHsn8vbIpkQNFcT0IPxddMCPXJdf0c5bLpAMFpX7+RFUihQJnz+g1
zFVL+eyJAnuMv1sEhClWntlohN2P4jk6S/ebEkGoVAeLit5RgSqT8E39XBqP
Q1xP1on5Qu+9viBBRwEU3706vWdsT4h3FaI8GZj7dWEJER4rHPb0q6oqNkiZ
OdTwFTHG3BUNKLiYguQuoUn7GQZ49ovErQdJYZcjfIfMjNTuqO2CdBcsIfwp
WNHkKOzcQw++kckp70jVwiaNahWg979UVTL6YTGI6VD0RFBH5IxI33tx4Qs9
0AK/Q7m+xWzHcdm45BpwLHFwN6AkC+LBE1SvYOWb/yibxtSjpKrVcSCINPr+
y3BFRjFDvyRGVZbX6+zeCyKlWu7nwGT/uo9+Pfptik87YnNDVFJCAhpO+VU1
gINl5j2zRXVnFJUgC32vshk/9r7NRNvXzJ7745cmtzwOubwJIlcg7aVgEspB
34U7Jyt6YTdmr7Y3q/bRFUc7l2cRYozpqZMPwXOysJbKvW88cbKc3dEUDA7b
slVM/3cZov8m4Is1rZBE5gTyc52z5NCiykH/pAgrn72+5mlw5CW2PKZxjLWr
y2E3Iyf81arueqydmRfyul2oA5dUUWDCxNLzAMZls2sxF3XuY+paQb0qZuD8
kaq/1XLZFJVmkxi5ect4FRkjh2MGbxzZRSE3by7FebTtAl2Al/f++GJv8hhV
w/gEcHcMym/54QBraBoogi0/MiMecQnUwzrkJypwLt0MViwtwNwX9RojuZY0
FFrIu5M/tBUy/XL278h7rzJBP6u8NI41scvVBhgfMy53AiU8zgRfVdsmus0y
3eETcTda4KiFah0P1PJ/9frsFyRzvUqVb37wnrt6/gmugtWpgkkTzS6gpHUT
6fnbf27MqOOSCcQ6JcD/sgpL7BZ88YchU1mUMURLH1cEFIkyfoGEaGMKeDRP
sRsGepTXCtXUkpV4HSwj0SFgWeBQa11ZvbwlX8Y4ZkIYiFRTyPzZbEh1NXbT
KKua0uewVbtNe0wl0/KLm5u8r0kWUi2BTgHier0SJq+MHTWyqt4lHIuKPiCv
Ft+jTiD5m9z6Vfz05ukoJvwX+6YrJWgsP7pUYI5604AOz+0lH98UDEUd1jsE
WH0caNncR377+NfHDHhYk3QqHV8OEvho1am/4ZcY8WPM3E/cvZTwzt3Hdsds
4qy9qnfEcwA4w+Cmi0jyf+fcpHlRy/YFJ4mE4uBaMohyVaIWna12izsGjN+X
O6RnK9SaZqQBrA+pkoQWbU4wqOVn9s2ENd4BthsHSdig2s10X+u+DDuvT7Vi
IGFGlkzR0H0z7d+8xxI4fLpV8YPB+Wm89BqKkeAOi+gkFYWOjlx4WmXFi9b/
UxLl1t36VePHEzL7JhrfUCCjist/KhGIDRJE1izevP6eBSpP3mByRfR+DL84
8UFnNayyvTerfWYDACDgCanEaiK4LczKPixGCeb4l59gkiOUhghJN8MHFE0c
erTX5p76e+IWEwPEL3NRr3ihRAYknNPcXtfrjeq7Ny2ZvXIUQk+R081NRTgf
wOPi2OELddaqYMQoAW6Uc0OUJwXLfob3NAdM8SE218ZdEd5JkT+YKhH15aMG
6/F3UIQLUo543h+nwO/rZGEQwDkwC68KuLuqucdi+/JNL1b9xey9EFECA9lr
z6tANSjZabtmC46khywSTCYvLlC46w3vNYp4NQ4cJuLrIjijgqdEfcPaVKpM
Z9DJ/U3UJRutmngy+4TGLmVVzQ+J95Y61uDRnsycwpo+9hTjD9v5TmsImSPq
O6j49nJlOi2UaGA0C9C0TZRF3mj4X7Rhqi6rdLBkToh6Q9XRVt9OB91FOxbC
6ZLnerm/xa7lMPoI6Dn0jrCE4AEoIri9PJgELqF5zSWPAB3jx3RbtXq1pqkW
jwhZB+64l3vHQ2TI+a6aZ3/iV6qwm8YZzji3YeSqv+SLOE8EHd/QE4uOLYFA
sSxHZWiHPU8sKz5uHOoLewU/fK7eSItZyhz1DwpsCebz243viVohcYpK2+bu
nKneynP3ExHl0/ud6lJqUffQQw26eOQ7Hk8G62Eng7XzjsbMZDuuqEAe+Ox7
remlvwYthIOgmnUsc/vb8QhzomR7WKhcbfC7j3L5V9JmIK5A0lkK2CcvI3h5
Lycc/pUz5kMrMTfmq4ihSST+8vdgbUnDZk9X6VVfhyMJB4wX9/ROH7IvmQcF
A8NrGOcY8rp6g2gBFqlW+wcrGrnbDwXzA28K0Lxgoi6YtaUm/y9tG/jYlFR9
BJlcXKpfWcr5eHafiRpWGAe9PJeBi3fh0yqhrowakDbBqbyd0v5Wu5nnvLuZ
c7EQ0gE+kCekxN9PKqm/9/5ht6NeEHq9tjDQPTeS+1fJiq6luhYaDTq63Aae
48a/LwzVyw+1jGGsEC12u5+vT1CSIFzviH5Bc18QNnfKqK+g1OOid/oTf6fO
R+1wXDEkqwimV9a4LrW9H/KcTKhFR5406qsIZcVPfAJNgJ8IAvCEO/0Gq0Gi
/NX8+4H80ALjqAMDNail0eZnu7rl0jQC8fyDt51DadVeoe0aJ+qi0hBOvaoe
hQdjUjHmGN1NTvLnG0tHclLYmbhRGNPaJ+BenbjG/Z6mHyJnIuu8l/R0lEUv
A7gQnrm5Jlc9KHRcpQX5lpyFDkfZVmV8p8M4w/EszlmHcu1FUpVBhEgTNcCx
VunRT2GzJXrxwRUuX/xDC57TyrE+32Dz5431nSCHUSj0c64IFuqAiN/UIrIP
wdQOBAjufu/WONX9hFT+oLsRKVE/k+Wpk+r7GfgUjDaogyBt30XyuM109uTD
+l20xJo3e1Pe4FhJJ5PwMMyXUjcZUDW/uBtdrATUxyGXjerBqDMHCPTTNAh/
QEWpsn9Ke69Q1GvEsCSKAY+bpEs37f5Sw6RRb24UuK96QbXZBUK4zj5g2Jlt
qMMVYQnwakXwcSUMAnBfaUxKXNwMFBqNEVIFYdnJ0J9m2E+IlnlMC8Ns4MJt
sWReakYlbSjcXDdtASI63SLNvRQsrhJyIMVwYtssEx/szIClZ6xrxgSaWsBh
Xz2d+x62is2sqUxZBX9D6UjQrvZKA1drN6EoU2P1JHu+aWlp8NA/0qdya0gn
JEl54YTZkHBPo8POhfh0qnZC0vPtQacGBbnM/5ISaa6ifPyC0NKfFS6e5aKX
M5sI7wfjRF9DV4RrP5ClcAAKss0aExw/w36C1rmaNb3/4u7erq7pL7zw6ylT
12JxrNO/tiZh/ZP95Tlisnj6d7OetL5twp/yqPT1/skZa9SsUF3QvH9TGkuO
zpdlTNGmerEkpouI8GoWw8pPVg1oJ1pWcdgBrL0SviGCZEyDuAQ4vjE8uMEj
Tiq7k1Ohx6xBkTt3TRm57M/G2E4O1ezGbnaqeBIhP1frKnO+k1nvOX3a34Wq
Pp/fQWK2Cl7Bif4xQfKXBK8VObTUI1b8XC6wSqX93v9iRZjTUfLhn2iryvCJ
p0aBe4+Wq8+wA62T2nh3xU/hwKXOHzACIO0jIy+r4ejK9ag07uMQXqxl+lRC
8dnQ8H5++0gpI7hRNkDo23rBZM2BL4AuXtuL4JEJBubwuaN417i9BEnMNHpj
pcsFDZKqN3dEzzEJZ/QqH3SLWB0XiQT6GbQ7F5QBwoUvdtYWMJCNVY5KPWUw
CCExfqELjAZq+olgojcr+f4yhZExWreRMos4GU1NilOgAfdujWKtJyGj2EIm
4VGc2YJsFWwxawpk9zzE5N6LG4JQE7IItgQ69k0fzUSrb+HmIWBNzw+Jr8bT
IsBTggxfLTzJD/BkRPBKHHvs8QuiyoQVSolhdKG3cqMs6tT2VyJ87zmC+qdL
sc4iPCdVnz/cWgQnIbNgIUGrUIbmW4K4GtVdXwfwTobQjieVFtbmv5YS3Lyk
bJg6f78Xc+SUC0nm9RUY6jeUi3icyvcrpXkhdDnRRmn2REsFhOf8WqPyGLXg
MnMjA4vmIjIe79AV50y+mlbq4CACvk5KpaN0OjmJmaUA3++N53Pfea6ON6Wk
fsVV5plS26aJq80esYz7lmhBunZwpVTyy7feWvH5aKl42EWCOKqQfzztVvYc
vIeqX/JZ3feQ/XzNZ9IRMMRYdUej/m1uKIfrEM5nt590XUQPPn+Z4/0v3/pm
8XD3bQVg3jgWZcJJj/9dcYhcEiYg/65JbehGMjZaEmNDXCw/iCLZG/FzDfC+
xmbGDuZmyzZHrNA30qFi3w8my94Nu6nPWFSTv6y/qen1mmnBRmdPlYoCujiV
INn4KnEIiCaE4mg8Mv7Aw487Iuf8TKuZvDCmMomWJhrbnmkgFbBRlnlntcYj
X9jlJY82mZ+fYDD6PF+M3x6SPUBBxah0rNHwLeeLT7hp958rn/W9x5DA1aPj
Js2aVIkcKIYuJ/3J43vi18v2bkF21DUQPxCw2xicEqROlmavqRi7bgc66ohJ
kpXwFIlgMh3V143JRz1x0GRX9y1//yoSqFiocm/RyM6D4yT5xjVCpO4SVW19
9+/hZKvwfloOS4jfDH4pl5KUaFOphSnxx0/Efa3GW7jnE63U4KENdfp1NBAZ
6LdV0O0bV+y8Ql5nqkGYSrq2IIhA1h4QhCfTw/Lz8/sfFJzbV/3Qg3Uz3PpU
qnbRRjhv+eOvgHUSnj9ovZzDX/h+ea59MwzYVvaij9aaviWvZAaBPxawQWeO
uEDhAS4vD7/IxuwsIaVFRhxM4x2hO1HCI9b8P0UzVn/IAXxwvkCstyVoVTiB
+DrS0sevL/AJJLAbelINFy2pEVPZXN+Z/uMBVPAAlB+Y44S9ZM2Q2jQ99XD+
EgBFfh0NgdVAcYhgm5dFXyqkIoS+5U9/eWGWyJZcnW6U1UAclu8kBY5lSMT0
4aFyrA3IhGMNUXeNkulyi6IVq3qK9tySAiK51axcfM82nbflBeQgVX9dvO7Y
BuFaTbmDvZd94GbuZnFVqbnTxI45VjkwqLjZAD4d531Lpta+j2Qm3N5YHg+6
etH21Mw+4AfjMaNuuBJaSpLkdEjXrEl8NQ2cgSsmQ6qIuJq4IhRm+3seoAeK
NJo/tj4BkrSHO3mODR9SQbpqVZ4sj2/98FgiDgpzqPHEO52ne2foekA+BauN
48883+DOlxjCPKYQyBmTeD0A2Tn3WR7AtmCJzvXcqyeipZ2UAjk1Xr72emJt
JYA79mqMtri6KNZv9QXytJyJbLlWMYsbm5AOeud1SZzyw1zW/Mx4fkgh3Ixm
2bnLNc0m2HN+zu6pYVNTFEab326NHo1gFqgExzwevQ87Ov6RxPFQp93us6dU
NdT/WtakOMNpndmI4rl/Q6n2REvvFnwlTbFRkFfirQwTTAb+u+p3mt4FafKj
hohH0CNCBukqUsmcmfUYvJ2EemHRiBJCfNAbcdaov89xBkZtwbyUn47dmPAU
84PI1zndZXC1HePhyv6w0+PFnAeHaYZfpPc/sUNCmyCaUfKPfdbsLOTxz0+D
xrjJ162Qrl4tBbzgbdJNd4SMjJAFKxAde/N2CEl9WQJTkQFO0q8XkOo+Tg8d
x6NZt1+eWTF3TLwt99h+cIfEy2ERttRaWSf6QbzPCdsTJC+U1b+vsPk+cJ8q
3bvylV1RTB5HmuNjRDK1ZYfwi4L/TjnIaAN3TUBUIJlpcHOvDrxtg/6PcVWq
CoV88Q4d11cKlsAYCf/XPZTNm/mnPtW7eFAfiZd7JLga4mnkDxo67RQoQAv5
zMw0kc8f1+eLtpXtXPF2p87kAs2rwmZowmC64nmqZjAvMwUh1hqN7ypmYNrv
zNfL5ZVTP+Jca57yNqlmillTpya1Iw0PRT51f4Ng6mzm+LksCczixSkGNe/Y
hgqYcrZefsREAK3I8JIDARR4i5vLPfyzIXJ4nECsRBMDZjVf8ptf8ctLrVO0
7js9MJ2+dENiwAntZjgYQPxpwCeBDeq70zNNazcosOFqZCiOu1pEVr8X6yi8
U6JV1xyWbECtg5zorKmlgbw6Lgli19ICptfTO2mKWZb4jUCj8Wh/ycizQSBs
ErqKbixYACmHj9W5k99QT88lTGvWSWJgu18LKa75jQWAeWfsxuUnM7ZRGWqq
FmufFhQ66cW27YJS7GwXWsKLpsymXOOEZ7C3rIzem5lJtkY65rQTySJ10zlM
cqf5aJCHgtItVWujcFbQSZXY0Ydqw9bzgP/SCLmdJkCGhJxWRjdiOC8nJzvl
XPm9WCh+1Qv8i7L60UCHO+o0GjcPwaaA/FO1qtOvdHDdwFrlbsgWvK9F71oZ
juTEcTsM8x/QkXXPTm3LVnU4pH7MrBR9ZFeNwSviP1zcj3p1jV1v7VwDr1Zh
su6NPdvBEWyl0MLOuLZs1DrfRkb0uHWD9UJJXTCxQdvB3iMOcWE1y5PW941m
unzJN5gDOKpg34thTJi1uLvFFfmtGWtTViKYyFivgPhGYGYoIOEZ5/ayxeLO
BVLvolxE0jTCJUKpU/uiAzezUu9U54hN1UzSc1pOflzLLVViNhLN9qeglBHC
ZlDPAjssVnhAgoVT66hKqRs2LT60d8RkWVa+bps4dHy39CMJy1j8/HTHgzZK
WAD6/t05+1cCXBvqsqTQ/inTp3NEtPPmD25BBPbSsPWUUthGdsljj/IbJlfg
pPeMu4qUoTKrZHKemL5hMi6lnFuzUe9UTBw38Uo8wuflZXewLou1pqOgtdeJ
3uV3+AixviAnGRgoz3GIF6dz09oXIGynabUtun8nczT6Rvocou4hHb4Q8cYA
qGOzFU0rEhNH1xAY6a/8YyIWlcYc5gu8QCzOJWO73onfHNe1+fru75MceecF
RgsKFu1TKY7+xOp70i/jZtd6IyD1OkUEV5pK020AA1VKuJBCCwI+JlOOsSUz
oTCdxEk5AkyYC7SfxcrQr8xvGr93rJl7ZoIu1yMZRthW0N58I3rgukvJ4CjN
lsCAO+wvsxLk9JpcerZiDXavbOpvXG7PRXKFmrzLdk7ZHJd4LytD3lP8yMTy
setVBETUtCwjBdpt35wOVNU18ClgzGPAe15OxFPFGTgAmPNzm0venTQH97bz
JKis5HgISt7/uyOXty5fpu7sPthfIkOWoOM2Ny3S5QDHZxQeJRM2DyPwQST+
xxV2WQLgf1y2G7n28nk2kgtuGpTLOnfcqiYdVhpfp+3PgjQ2K78NY9rkIYEG
W6Ls6xjoyCH25ozsmNw+8GHwWZcesdM406Npm8RvjB4mCGeOrxSTw1khBe8+
2hvqlGDjCPIgqgEvA36uc7fwjeqKJoMiB/mDYEH9lXIL9VzlJ0NtQxYlun2U
FkwEKwFEUeXoDl+GW19zUfKDVFH3bJw0OY7y2tMloSpnEBoUPDsr6Ey6IabY
7P0RScaCPdURlzFFUAxoteeeBafLzeMrVAmuknPaur62b0BXa6WzAWBUGErT
wizKKuVPUg5LSUtkrzY08AVm0ksF6FhCCMbGQqnm3lQkHIrc+vddDYLBAeOm
CK0ebBr8KH0353fuaknaG1LzYXJuTalCklMHaYnN/k772S263ZTa04K43jNp
k+wBj76U+dFBEWddav32VJg6t+iRfB7Oc+z3V8T7kKZJx1Wfxvz4jzSMUzLI
TJfUiFYmkgWdEbXFvxRZxRu+EaSC3Tf52vHAB72B0pjKr+7bz5nsHbvRXZVs
ZOeNkcszzR+vT87v3RcZhVZWO2KHpm2yER1dhJSSqopHOgLM7r9iImmgAjpY
BNzXp6gG0v2FK45AyCSZY1hppBSu8d/VQWMNQtFS1IEgPAWBuD678vy4SeZP
l8FUAk+otuEqdGHC5Mk9/KIuI8BPd1Un7ms/ZHKwBWHWKxel8ucDdy8xeTq6
qQ5Dnu/TZtg3NLfAaffWPPTJAlpcMTM0mQJj854ebA9m8T0XdoM1kRa4OCet
AP7pAlRf6Xmbsy6Th7BSKBWKwEyqyYH74FKwGTd3vLhGH8pcdXdfEfITfWAI
bb7me4enUkfOx/d48p321QMSsxk+w/XcRmy0Ii3Uh8QmvfouyXH87zEpuNq5
8F6QEsnjb5gJMlsb1bwPwvUl+K77OuhWHLufsM0BBXD+bgRzLXVTxjqZ5Dou
C8w/vBI5knQR3Pp7lSbAUo7vry5rGuPQYq946Lfb0YsBzfB3KUtyewSfSFnw
6dW7Z5cLXUyv89yQNDgk21Hs98ATGTr0Tvg3FYApeU7vmS2CsiDdbnrPS3tm
UHEVJriO6zQqqJVGSCH+S2wnUkl6S0rLDagPfe5aUdDVaxRHlXZh7pkY3nPp
WUVzKHuv9UARlPjHYz+/HI5RsSsBs4tDr5K8K1t3WRyjHUfykZb87zZH4rrs
Qn4aIzHr1a8duT9xUV8cFSfhY/4BlHidlwtbnxYD1nS/GdAOf5J5/Qmbmef9
bryZ1+ZICivTUQnWRJI4i+mLonLLo0MsSqVzh8SOlcZXokEo/alWwzeumEE3
p4U1d3lPEJosMzUsHFfGPIU4rGgbbH7U+xz2avX2ukkEodncIrZoVZE8tDAa
lpZls8MKykYM+U0e9df7OHz3e8NzXyuvXZSU3EEzkZCPjzUtrHEKvMfc38ck
+bOo8a9Bqsmq8GECVc57qDe6UrB7BLuXLdCKDvGmjW+r2GEChs5e/FZsr7/3
ENKbrdtgwKQegPmlrRGM1vXfTXyGWgynbOwT7BOrrjjhVvfKue+LSTuhfd1w
DlKOLsXjcsxrgbnn8TR72YtpdOShfJXaDEMmJEkMN+8pigV7riQJtVPUobkL
2ddrFQ0bsu4iOvGZOrPmOw5DQoqZrSNYR1lUAfpG2ocBlo7obpdNZCeqGy2q
Kx7XuFDE+PdJCfjV1HHgajItW4PEBxvNYvjpaclyircPz6aarzh/xds4DxdM
mHSJn89yT/x97/weqPq0yebHDFlqftOUkRP/6+hICa98qHYdQKD05wTC7GQh
PwURFlFz437YeiiEiliw4gSWSronTjZ+c4L251tlO0qvW7YfDG1PlKjMOQ91
I1A3iHF/Facb2Lbq9dtilToeRBtbhOYheJml0vgAoK0YP72joZ+51LjYZZgZ
ZhRH7mQ8+7fT4oYbIRwCOAxROc3v1C54qvHt6N/PX9MFH7kQTe6zUadkJGq6
P8/PHluFQXpyTuNc4e61gHaMuEMBwrbokgdtUSNbFNNmPTXU2F9iz5uqrEsO
j0A8doxewF3aHaQkFjF3R/JJLp2Fgzg34CisuMTv6Iyg09r95TJTCfS+Tl2Z
I1TekX1WynuK/Xgq53KRtryyB58pEmRxXYnb87uCTX3/aAKesx2mXGSCKXbb
PIUyozsnvHednWyWiuiRnhO/sJJN/N9j4SYz5eJMu4qdUdGeoAmCj9vRjeEN
rvXUzZBDVowtgJCuLLJHYUrP3P13qWvlxdqxEaq1z4UTokUeUNhCzcGLbFmT
1BrbWalK8s36jZ9vXpl198yQ6Ufqb9rezlTiYR2wFHPyRYOXz9rUsoow+5kp
tta4sZeveabZJD7hfmlA3pkJvcBWpwp6qTD8uL2Y3H8pyb7ktkHXRWH+mdFo
QcDTynJmuCDr/qeQIlQT7Qmfi5nHS4zNTy5ugjJxfd8R7G9wa+yaCec+SA8o
i1RdDdMQR6x01itHJdW4+iulusC0WusoZZX1kdA4gfjtTZXxxRpi4aSyJPhZ
09F9qU3FYDKG4xaJ6umAX8dGYV85yU91mX/WJD+3hi1YVdJS2vXvXYho327N
rpT/bove7i9n/iTx6uVoOouNm/Zox/duw/OBAmpUPvEe2AuPlADBzBRfI0Qp
5lCdYxSlOjxctVM2lHnH3vlPY9eSU4XrpHOvYG2AqlmrAgRHyX5sVjEh9F26
x2mDZtwtMiwmXBd64XzOtxvkahdL6X4yaZULyQejH5WQOZYa4BuSJEmCFUp2
u2oLrMGw7L6zrHFH+vjIE9fomG0zpjdv6wDVlVFjkd7/cJrNS0FyrPAWtn5e
DbODwGsXC9Fm/VgMtfvt5Tb1CgPU/rTWRANBa/MbEJU4m6zncMBx4BkTHfJx
cuf/6HC8/e54+suY60g74AziU7GQELsvXI90Gd8OzponHrZ65PJzliN6rTSh
l7B3dymv17c7ta5APiffAPGsAg7+IxVBQPQHQOo5moW6zT7RNObihM6R1FkL
3qMOYn5z3aBwmZRypHZ+GFm74WW0ht2doVvLIQwHxVmyoFXmSv5RwVmYe0Zi
3wxyU0g3DkG6fp0yqXBp+8yTQ1A54lpZkfRvyM8R3pA0F95gZyizQtzF0exQ
r8dfGJXgH4NgZmLFWOsSEuL35Cq7jQB5rtECdsMDgBouJc9cjEh5+FA6AULm
fyvSLqMnkoY2wy4hu+nDyZeuiZJeBUVcuN8uVnMrxR9eIlx1DTB4fEvKQi3y
oq8BrY8lIdlz+u2ROXX6A00l0Wnnk8oKiQxpwIJWT4YPl4E0LIj0MB4iUvSF
vPud/ENrAooVg5ESMTZXIIuJIkNYCwr52MLgTxLP4FzVM2CTgKcqH8WyVs7l
Sz2e/HazBF29QSaHLKpq4bIjEMEgUVrvhV/jxqF/QdXeO1DWyUNBLxzYFFQa
VnXH+4CiHLdWNjH8X79rsObpO79VlExfxXUoCw4hCzQOCdmQXqQM2nKUUugG
iK10iJe+wrEi5po1DdE46ZZVNC8rBbziDCertwxmn0ASXIDWpj1ls94mdSw1
lKEaAIRSJUajtPyN1bLmK+lmg11jlH81C1+JvmRtXEjcMmdigQmGspvOnc6D
3swEeqPF1mWdYAAsml1hooKomA3qyPP+mvVZzKbhA/838pRya7daPcM6gRWt
1+2+j3nAHSuVf6x3saZb+Zu30ZdMhtBTwi2FDjQj9lJR9d+acd1Y+baqzLWP
O/Mlz4TNySIajD/d4W3+N1F3ChO45uJE9Ryp5I44oKqnwcNRi7EllztirH8p
fo6OYtMOr8o+QQgO5koMV1rocPtzUlsfmW7rbmeVYofru0T7m4NuPMvGDt8Z
YkatgFG0PQgCOCsm9ofdZPMI+WtQ6wfxs3+Hd/iGqnoVQLQ6xWD0liuJm7Nf
X7c1qnVMSDecRrktCu9Hny2CQHDGb01vA4qfw+CX1wbQ2lDJPrL4n1/K/vZX
hRfqmsaRXcb3Tf+tdZ5s7X7JejIlRq6DI7qVN7zkxvsRDr8y8gSsLVXnQdJN
jDbC33O2kqR2sfPtw33ZzXqUHLDUTggr0LoT0Nq3sSPnIz0chhUD4Sbt04ah
p3WQitdYr3Z9ViDjAtV7cTemS/rE2rjZGxogAA1boDx+EZuqt96ovqLNC52I
w4VXczY2GDZxPGT+/Cy1qOg5jN/7ou5wd+FuPOBP2OTJEvMeQp28E99LM3X0
X0ANDiTzRHbkmTHuflzrXWW4oTeAlzD4+UokWVURrdtj0GMnPPg/xs3KYziQ
dl+nVyhe2GJAyfB1j8ypHUgrsoswZeOVuACsxyjGnCHqqt2G8wywZLrEGRWN
p4zWmTv+z7FU7QWOFcWaZe6MOn+cxCSFvpADb3zyiDEUn920ydy7QTQUdKF/
UM4XRpqjSlJ/pIjZlDL2btqeAUPdhEyqdR9tTwL2r94zSRwYCr+/csF0ZZzt
u4mBhZTSECgMtwR9xpyx93O0vHfRzJcwxmE8w+fZeExved0EyEtSU/atJFAH
3njIPTVtCjLqmRQ8ryL0kVSIsgYcE7Cjek0OajjBDdDa8OeJlRQ0Ls8QuyVH
JBhMBCgnvM2YIwdbu2jhszeyzEy2GIK/fNtdXntZ7+BWASai5urHVvvH2d1c
FQ3WySgjHVN5X4zs90P9u1p+tsw2oXnTNSzZwzDOIY2r2AlWso6iXsnGXT02
ONrIZnADCzD7yVAimLlKIhaqKXshA7vICJ5PiorNuRrj1Tidc4vdYP4h0vva
oUOQZ8tDrdZQpGuNO2EMuaxQ0nZLi6kRf5NVF4jDnNI3WnedD5+tieczx5iH
A3CIS4/u/dPlIT0vDvBKyPQiRaF/hc24NGD9oq1ki50HvIXzcd9xltxEYJ4x
nXlOw8YbRjYDHIprzYbWdPhus2+xbEC+GpEc6YBNzmQm64i9IOyLF9yV+cX+
uHZvrng8mfDtJ4yMp0HULhQsYBHfZOXtu5Lt5OYKOIgYWkV1OyObvbU/nAc6
pY3JfTnyXnGIBhUtheAxNrnR9j18HMShzDdvKkHl1G1/FZ9VQ+Q+eJOcyjqq
csv1EP/r9IxHXmM/GSbBA5+5WE/fzmKkvBpQaNO0A3RqZoJeVbEnHaARWfZ1
qYX1yFuG/JnlfusbWQnyF24xPGxtCRuglANuVBQLsl710B8LWC+8+NBjClga
dcdnBb6yRAaiN7tiytLGjLQY7irTZGs9wWUxOF7mjbhqP2j4IA4yB74AxTi8
CY0VS6b+fGFUWPvZVGdZSks6b5WDpd0Nk4WmCzRLyZZsJrsbqrnxqCPt1BE+
Me2czFuKXmLutQtWc3osRnm9dwPEEeUfH/9NpII7wtCEWBZ2QPl0m11HRuc1
R2Jd6JPkJ7gGMZEcif3gL6PrY/y/K/TjFk86Slw+0yxD+8qGmG54K6Se3vBZ
hIHf3qP+l6DcPkvH5mlAgYsRitI+ciHGpCssqsph4Dw/0VxU8ACXWS0V1KxC
rWsF/1IguLm4Jdqesblpq8d82/exeUQppV0bw4ikwDQcNLllQgjnHfmIgJiE
Ob6aUSeUD0BRMUbWaR9ciIsr8HkOFl5Eau1nOABmtoq+t/pWfGShuqmfqSOv
RhNjoRuGJi8rXEhr0n5dwipqTSCh3MW5AYsev2buXsTuWHyz5Z0b+2DA8QX0
D466r3Ww5dl7mYxA3RJSWUlrzkUtcylkBHnCwCwPCXmzeofDvZYs47HX65Kw
aLCatGnRWQiLxtw3q8jEfyrGEku34FDIHBp+MQZiqI8dy1j06IYz1iHK6SKZ
jkk8r0+kHqeDIqickbPdjNj6Rl4sQvEQkB7q0436gNtR6xUG59mkEahmU+rb
7+SQGMFzsqtZ/TpttyFAf3a7qrcgkAMsof8g8nqR60lXUTsrVDAHNONhTPav
SRVKm2mh7R8FSJ/FKpAjyqgGU8AfOv3eAYrex0qbc5Wnv1lyc7LbX06pa8CM
FdQWl9ZITE3D+9Vplxcs9h6eO2GCFn11UxnMIHpb8HhgcId6Brigb9Seqy1f
I4Z9m4WKTq7Gt4Dzo9OOSMSM2R2R+PAAHYQF4o2qaWt5reS95bvPtd3jjx55
q6AuSLqMkxZwvRmu3AX6yc2auoBY1C/8kBNsiZgR0T+apc98VksZ4HbcuzdJ
eOPhXJwz339qJU89tTzd3rePN+GGw9KqEKpUuB0yEE8tGN3J2ztDHsfiZuM0
WwrM3usvE4WR2L8uuhPsrdtqo3raXkXIbDYFMZ5kZ7Ra1vqg3f9qojuTuthD
/hxFEa5kvmoKINWgrX237/bsh4CHbOzfSviF6P7n9mMKxwPHQhLcdaeytKLZ
3M1Q5ZMbBDQ+VQx+gXr2Eo6f1U7d9T+NnRmKR/llxmvxIh8vwWEfaqSXdUfb
oLC386uR2Qkx+hh0pZq3oE0K980hx0FJFI/e3k4g3sHwchIjynI2E58MgADf
gFVXUD+VdI0epdfCWBZSAY5Reuwu1eLYSamgiaQFe45d59Edb/+0BYpXvDxd
3pSc7kFb6BPJy10xWfLgGnz2h68XQacpCjRvszqgK+S9+aZ6qfaOtRv4IxEX
WmKNtk3LAMFUfZxNvwK37LqU7TUV8bTe8+/cXK/vRX+bAVNNX4uFXOQlTR6p
yDgC+bD9wT2s61w73pAVCHf692mDBc4jcM0tDFp35nhmSsaRqWWzFi+MB45v
7oXdTwPtmCYlzSWOfFWPUdKc5tM5HF12pJ2rW8wUyA/hIK5mvPjDuIRZIZuX
d5qBcky9/p9xXXdoV8v2LHBKHtlBMLcbvl2mFBpcv8aVhBEZR5UHcsCA7SJi
KS+iohbwa/FLTjPniCnTk9jDId627dHgz6kMBXzSEcw26OoWJpVgPbVHOlN3
FJYORPyWgdalAN+PdaRFfmc1vLZtVjqmdAT9LZH6BhmXMKIxLHl7J+dtgTy4
MzB1+tkejjn34230hQiF8ptiqb0RRrb8r/b14KDSuzex8+QQPij1LxUyUlGG
0wDxGfEN1lzA9Lc6sCVUKh4fxdnjBfyeHBUL9mevKiFr52wWFf/li5i2qHsB
mw6s/dYWyPsc4E3zGwa3UUUG6g9tyfSJdZs5+BoLYHoEPY//VZ2v8fGAJE2f
9BSjUh8OAvcWrdkluVr1jcatBPSQ+5Uu5Tn2gcjDWCd8FZ0wUQ5pbRSQG7o4
Yf/MxGzMdSbnxc0bMG87F8tan97MChJRl/4YCOZjd4hmpuFEZ1fg7vA6PJYL
MajOxqHicUEjvVh8yGQ19CYTKiY/HGcLXib3uirWAGjQcaZ7Y5TbYsOzR+yO
bggmMPE8RJknWtQ9av3syUdfA20YV5K5NCLqSHU4hhbngyDPcsy62FKZmBuZ
oLX8vid/dnoSRMzPEoweseFjB8Wb7D1yVDnRRsHooH17KT0JVZK0uhCRbR9O
CV/h0COanY1NFwCynGvT/w7kWa6GT39i0aFf2nmwxZDKexPc9VoadlCQe5Ns
rrXPfHWSEZrGcoNOdF8raeamRvP5PQknQ7yffA0BCOyq1NuvrOj8/J6o88O3
ZZhmeOknq/HOivQfy+j4TiAMy/4OEKJ5Q+Rom9l1FkfJw4ZrXcw+cbpKTP0x
q+TThrtJldtIH4QGBfL8iXovchHpLNrEdbcPRE6dSyUW3dWmHVN71dASI5sI
tkrXHNGllH4BV0+gaTWlxUMccbhuGnT0E7jk0QcYAtFVNWLwRYpusUhLOzFH
QqO59/Ns1vhb5DQmEaSniZHM2lvvOil3IinkVkna3BM7FTRgXD6TvwEqmrhb
yjrDtm/UaqSYoEYpEI4352HPr6g5dQTjtlUYpPnA9KWPDsQBVK/BqKjPjo7V
LQhIdKiBUdxElS9S+PuZRp4IpqEv4AHBFtxPxzLtGkLg8zhQpmnNS9aIVbkj
bQO9y2qEggoOKGXqa8ENf3so6QEHysr61PIeCbaRwRctXiM6uxSQHlySuqIa
uIxLNFJSJHPveOaxWIiJCkMNvOiIq7meKVQj3FSxLpZE6I+8Q6lNsZDSb0Qg
dC+MLjpq4T9+aJWSI1szydJHsfCq5qTWR+Fz/TmyFsjuCBLAE7EowPxWJgpF
osT6yJNTXUW/OrIiGswjqNXuDfZmMMOBZwj0JZN9Po/pb6kxoAYumDzEPhTU
JasMDj+yMRmfb3YtNKTt8g2UFn0eOK3KuuQxuFki2ISzz0v88lerC7hXIX2i
IIxWaPFgs1LdlAubSWcsyQB9vnuQGvXlbghnkK7FFQ2wVSDK1VaLYSPjFQs5
1LKbkmpbVKKNaV9I3PHsd1JECw12AUc7YADPVueEOMT4H5odWSBL1Z/s8cg9
tbC5OzpAZpqFioa/peh+upsIN1qQ46dWmcVJLpVHwSAnEFTMtUb9j8aaRgdO
MB8u8XdAYsbuXeHGzaW6EzzqLFqKBX4W83tTNxApeO18WC8ZLr7S++Y9wIL5
pxa9t9Mhu8QUjwNQsbRkmEN03XZbYhl3WX3qN2XGeceHb759DVakyW5EZRw5
j4VLzUpLllIbBS/XkuWeuzc5shxNDHg0xq6/SSHT+WHnR+Z+XAD6H/tKd4A3
/jxut1zvD6Hl2WvpUWqL+rDmbnHUgY128cHtoSopkCWCF4aSkgTgGlQE4UIj
UkNjg/tdFKaRfrVK+e2kvq072i/MQE7w3C1HWwwgBo5q2C6wjObAmqiYt/je
erAGlXytC28ZYCnRlxbaS6c9/l+V/blG/kDfHaLkRYB+Rv3jbYH2aAR9TDzJ
OoAkA0Q6I/PDl4SPWXTxBzX2TWeQr3aYiaGYXfSoIRHl904vCx0JNn3/qW1T
OX4Y/Nwd5+xaz+DgNDrJNkER+5Q+5EEDXvj7OUaNCI5pbm7m4jkRzY8MwCGr
zg1VarfaZR2gT0tpIRtJdyh2HHczabqq7ZrmUypvJ9rfQDJu2SzWs9dv687J
lSZOWb7tgF0CCrb58gaYh6jzhK8XG7KJ4AfnYvfC+a9I3qiie6hDsNzi6I4S
ZxlX+Cbje7sOhPEwIsqkHIkan9xxoalcFuIQcwia3shAa+oBMNnv7wRbWzR1
WXSS1Jiu945ZrBryrV7r9ixVlYtlvVxBPzlfSDJRxsKSKQAWj4CZvC40U+ML
Qj6ynSoPEanaLJOX4h7DygLWGs7sTwXC8kvlgzETuxk3bAcWG6TUh19gEnJn
YzSsjQOH5fInHNoGWZRSjp7cxV8LY1sXg3RiTbXGAOY1aROLhhEu6S+5BkRp
Y1NljpHTxrYVfNBWbcmXPfLrdIBFD8sz0hpjor/2Ttr/uN+sOdbLiQPLVSb6
s8eYUVcUeINVFQ+ceXCvjn4TT/r8O/emI6z1nt1ONLDshhWdA5HzHGb5hAqN
2ggOzt8PY+HwU+7XZCInAzsSgTpubXGV/eUYwgmBpd9X6tqlh7/6/cPZXEp2
/mdExFIGApTXk7yVFP1b7EjCcHBhBDhld4X8vKxMaODLez/jcqA6O96hP9pY
K3DriHPeNfMVmE+cKtw4BE7G9N8vH1uc6WEG4hc5b++jxWRrOXBShIb3oPUW
OQWgHYhIF3NX4jOltx9jarVSa8l7G7WZ5JRdUK5gzYseSxg8/uW9+h1iDQ1V
VLzbrtJ6LDMVNDF0osjne6889IPG9dOpa0tI5XfW4DYzxdcEuMxxevINpo8F
zdsklJDsS4XB+EOUmL+shXaD+154OHqb+2TK2sZ1DYaoIgbbxUQuZJ0+6W5w
0ASJSlMawEBDuYkzgXlz3B3/BFVr6X11Q8dBru2HNy3pUbt2CiDaHCAsbrK1
XMR+zJbYcsOwWRzOVdzwVjJ1GF4uldlh1aAawTJimEi+OH7otuyG+Tcdjpm8
+hhQZU6s6DpuOiVPHPT6KgdkjTacMHJ6kNMDOoBvwqoehG8lZn/qPs/FF/L/
iyu03jy1iu71Vd83BNtJcJRs7yXYgoijjvjzVRESr6x4CVFB9sJ2SXpKnTfH
kR991R0Wlf6tZ9IoSShXeXEYIL3mVU5FxtRg5rU9mWlWgf2E9yLvhjUggYlM
wXK+BMfQ/9+vX6+Obp4O0B0qYge8ECggHLb/uEJMKKEReBG5+nfe+VO+681Q
fqhfD8CcOLbJs7PhY9F5NYhaUZ2qQ938j1djSBewB9ftcpBe7TmAUGR35RKx
rRkNx+vwc+OZ6RV5htMvOS0uziyoQmNzK9B2Vwqs7CfoB85ZKUJLCrEbWQqk
XAFOEZVQCzf3MbEVGynLpS0PRnLJmvF7uS53F3mX28GEG0co+2HG585aHzFQ
3wr33wP1l3EwV5V3JcHJGP+Ijb/l8DIHfiPBxG3dv2SXXilCSRkPW2jnVAYr
nMGASXtUxPFbii2+EFYCgCd+lAzJkRf2pOXfoE58eZsBZEzuk0A9NMXCI6F5
Qn0AfS6soH7EjlIuoqoTbAnY3bB4zzcqE0eygiX+bMvb1HavY7GtFc0kXUjm
U7FDPWnPwb9VQgOCjmf8HUowUMn4emu5vh1G/J4R+oPuuwac67JRdByW8FOa
rnsav+koXESWlQHv0ABHgHfQCIueTBaSMxBj6yJkwXYgYdT0JS9VmY3VMgsO
YtgaX97aIzpFEa7NrMAvfqE+OeAiuxke/bHooZdyy9EVzpY6vHDIOnwGhMWZ
Zlu4sFAzDf86uNIMglL3s3qnPlYxaI2qBgPcX4R7L6sN7X+zKVAIamY/iWS+
vmay2UDXfCW3XUZBey/byA8cOq1TBzNBUzZWwArDQ28q4wXfGKkNczDGBLaG
mPls8YOZ3EMTeTtEKwUrTUIURitfXApBxMSpkzkR7ac3DjxZui1VT+IOycXx
4miZvm56TztUlMUkvmox7XV0XhI5LCWU5kSsXS9mDEe51lgJ5Eai4Wyesa8Y
QicU4QijfjF/3DGzN858kYUslrADMf5oHYXAU4ol4z/eM0H5DGhT1bl8R6Z3
t0hgXQvxzitDXi0vX7DuksEdWBMgGXFKKWR5bT4rXzGc3ACY73cxPUOIG8wg
FQGBvqeW598rKD/IjR5zQapgjJTByvXqAcD0X8hfAJlpIrRbqXBpXssRkXQc
yIQkTJq1dsIRpDwG+EU6eoY43mze+hGKgPGTw6Ak3e8+fM54xEmeGWdaSMqk
E26m3+OrCXUUINgXVRdhzaGGyTEY8RHB6qeLciIMrKHeEXxef5qCPPjTK6j6
rwDTwCcKseyEVwtW3E61Mw/nkO5wZLiAnPIqfz1rathLMdX3jXfuXc9QQugm
gGpZ6c8nZattNXb7MSbZEQaItx2cSPdAQalkz3Rjru98yFxM+IYzx0AoGPVX
zLlJJdDFFcX2Pn2hyF80/EgQa6Xe1zwIok7lNmw9AGSqLmPgoQm1VNqv5ANu
qKDdCcejv5l1eQv4NDVA4KGxJoBcUyXZfu8QzpymWbqGI6spPfwQRTdJA8PH
SJ2eweAmNBtIq55H8U3etiaAdSweaewPGQvF4cVFj+LdkCM/3H7++5zhdxka
jXh41ArAE5vI8+/4L6DtkSz5xNqZ2JqvRcoH/icepAYKyJIi7jSKR4KM3VEV
7F7lt1sEuLie6kIgBd6Te+Bp7w0SysdradJiuK1Jih1b4p/pLn3fvUiMbWHs
3GYNAlUPbk8FMGajLhb2l5PIY63BH/+wIMvul97dxNckJ4DTdU/KasTEkc67
r5rCQFsqE1rZ7wXPYPmtvwyeHNQMQs6XIlYpZjsDH8AbCATxHgEutO6sZtNz
qbmhAGcHWtwuZv/lzRCBw5foVMeOly/aFTIoqH+3xHLQgbqPCMDeuE8sQEGy
8Mpg7B2TpP7YP4yHt6n6MWAITfpCJTcd5ZuutqSYImm7kntUjzEiMAMe3lDE
dRx5hENiDJ3D4g5yVAckgandXqTbbnixAYd89+9bCu5UXX24SyRdQdXnAjuo
sEGMEev8jx4uKl4Ef6nBzfYbfCS36qNzIhGwlFYev4RmZPkx/0c8Egw9Kxh9
yH/9aGe3M7xGVhXWPMmbw6OQkZ33Trjxo5GiIhEN99UJa5LjH2tzHxLxartd
0xovni32pOqLezjOqbLl4pdLhIMvPGmHJAifJVQVC51P6A1jheYR2W1binJy
DPw1rXRwoNa1qdBC/VJHcARC1V0qC+cQ6kdDiyVVofzTkwvgQM+OV+cogID7
cjenyy1Bw1hofvdweULTxXuH9gYZt4x9UKdiIkruNf6a8qQ//o8adrjddyEl
dzVi8TDVVcPoLHFpkWDOw4tNBemGO3lhJ+NK/7rPoR0CdNErMQQJ5ErUfHTi
0VAQh5Aqt/a+Y3ISYUZw/5LFLFq5MWjdX3j5t/VijyT33Av0t0YPMraZy6kC
kZahqUjfy69z/CUsOwmdKQsC0KApwxrexrbKQhHWfSLVGD35i95pYOyOqt3D
iGJqK/rADOASU80VrzeKPlq4PfyyYaollBFEr9/KmPKi8RS4h6rR4WV1FqVS
nIAfZL0heVlIh9fB+SYnLJ6upaHefh90lLCeGN+TBdMSwj5TkP+X9AbZeraB
InDdaeMmEBcCVWRaIZo50ecLIVkaqCI0jdSmSZ5GDpNnZ56Kb3F09Bd3Hsxc
m4xNDktYJfzpin/ctfPhvqsareDbXTOK12ps0L9xiv/VgdPMg8rbUIvbvfk/
qyLumhnJGcpVKHlhhYHcBd9AW9Xrqp9TfbOcYxiri0RK4HdB3Tvh8pGIngI3
pGduy/dNGakxzngKgxRpQeOIoV328NFdV7eogcfIfB9nu64i4ngMqYtlhpHA
O3eriaqftGBBu+93k9DGiVSmkkJ/hHsosKhCH82yx3q65drSjEaugmo6O9CT
YW/kmIcBxi+aAO2YRNv6/D6ppHeqt6DVN/LUPJXDmwMKcskBbjddOzqCHs91
Xj6dMOuZ8zmNox0ggMe0Fk85MzPuvLDKNxGN0Y5mSB/f/iZHblfpPNMoQGtH
6SWPGEq8NyydHuNMVvjQjOlYMW3rL+/YQecv7dH/nohubdwgRj0mu2m+dfa9
Trn39kQ9siTD2GKz+8ici9txEnG4P4uJq3WTYez/PlA9BUHzBNMPRJnU2W5W
8q51r8by0BKVlRiXu6MnUe+/xj4sZ/D0vVIH329xQCKzESr4YKFVWalvIXXq
npDgM6DVE+mchLVXmJNYCei3YVRgvo4gjOsQ3UBIo8CeoNXwR9XH1ZxWHNjd
HEVS4AM7WCKlpbuvylFLpv0J+1kzlVrx5PLof9NSCdIwAQoUTHTeVr4a8Eaq
w6NvBbcTE73xkWVLocE5tf/kSeLqpYkFFk3i5znAsIOybFSSgsgCwrL4bMHv
y1heKiVeowulgVoppsaYs4KOGNCjYXueQkrfPvJ0rJnjwsxhkgQx3NBq26wC
2shQIwfPY0xDQZp5lpLbp5QRzpSDWeLbiSc4RA4ungkRQNZoHD+RRu2bVp+2
J/N/27ffxr0f6M+mHZ9RCv11BiomLIUz/AeqZuUYuq7mbH4uMlHnM62oZgd8
kCx5Ted5ZnJtScIoUgN/ZSIcfaXOVXo2603y9tNCi7TBJbMyOSUAUPEyR2R0
dS5VSAQGVYV++wtIUat9Uv4ZDihNb/ykZgMYRo8nvPtEztEtO4gQL1KA4KFM
Rs2omPusMEfMZP9yEQ9FAtQmAoYzchYXagiV7tnJRZmFG2BUA/uumhQUdP8N
BqUi6SJSiHE6zwIB+XkvE0cUYGsSlxg+TRWLvkTovns9mie0WbvdhKSRdm2D
z2ZRe3ztOpyZmXbUWPMkR6/QP+G/o9b2pXn+C6zUnQidw/3MlouxgAIWh8JU
9Y6mrbebOjXA00HEkkWCSmNgy5uFY7VM68JZKejC7hYPFMXgqE7SRrtDX0/u
euyXxxjr4hZVKFSR3q5gJ2soOC3THFLUlGyKabjeM8QA9KSZ2nikg5+xjWDR
fExt0N9Lg4I5aqjsMxpLormAewR3fsV3ycDSuOpnUiIKd2ZIB0H2I+vCjb8P
3q/8a44C3W6NKe60nioAH+zZb+DxYUihPmE0G4+D5iPEH/TrVYogEn0Rwcii
nIiYuTPb2KSS7KYgHQda4mlv4hynjJlYu61s94Bn79fKwCer8tLtbnKIq+FR
VMPOdrxHHQ0hfilBOk/2axvlqNwtopo3rYApPlt+cmggM3+YuiLnAP4pRcg2
dwbUAMg5wjDZF5qFvXyVnz1LdWg3hiLiOtdukY5NTZzzDSZ77uikeeAig812
IEa9tDTQeOSDuI358nk3Cs0JL7PcV2Y+F7GojjRypzR2H4H2crrONhreTemZ
3yACoCLq2h1fFoXv0WySWp/0gVKhy5FPXygKJ6tEoXcLP5TaxvZ6l5zxoF9E
bJO8n/89J8tfEoGx8Rf40HSrnB7gArz8GP90UBlXTH0NcCzHLKYXPCTw1EJs
sUkTB55qp+FElscMUw8QBbjlEo734EdUQr6UsWuNmfn7HZq1WuB6oR4j3RoD
DxaCctZaZiWDqW4b2tnY3i+hq/CrnUZMDFEEvqSd6yzUN3fZRXujLEdMSPEp
EL7QauNNbNXiWr+Vxcct2hziu23zu+jkZPP5wPx1I1YDPqa8erLTnf+z5gkJ
GIQQD7tCcoBfYClWXnWlaxLUJBgjcfZuZlugofxPr6uO1Kv1wZoQA8noz2jR
uH6b7+Dw73SUBOSOV2X3BGAZzOtVLtHw98dk841pKAtNNgQqvc2y8k+HPoD0
B5NBizVZRixfBSHgNtwZz/PUiUN8ziVl4uJuYJ3TVdczVBeuLg/zI5CHnvsN
cFt5UMi6oXFG2ew2YusWtjXA82DZd1UcmH1nkqgZZzmsESsAibRMiutQE/zj
GkUbhQqUwIKB3UG1Y+75G3CZmdfSWfFPXVLMm54clW+6u2kg6js8KkwC0ZSU
x8RIv79tXAhlihWgh8q8kPHUfhwxGDWx08TXzvKPNLbvoMDPKsVKQflklQNr
Jt0VL6nnak20ZiEx5W8X2II6DWI0Xti8AvvmGJACDvGBYNOgW5aDhEr58+1F
aC6ZRBHpWm10QQ9w4qo5hsR5bJnqmw2vqfD1qOd6oMh7ONqO3rDiLZqWhTzi
QPtY4k2FPl3J9jNfi/5qaOq7I5AYuvsUD1w/dwwPiF9Mk7RUrBJgsjGPx8oK
97LM/vcrXiZSXINAKAXUHdfBaSeAmGPWmq9exkk/1zLw9F/uuxgs8G9iGBPC
aqrtJouYK803JPNuVRc8KYZmco7U0XMJAg10vy2FnDR9JYliska4Hs5131Fs
pcGxiVV7z0IttOshq0BJrf/30KA7HqkdzQW+l61AX87HASWQKUY2kNW3gzic
rYPwpaNLsLk3LZGXWyx/EXXlZu8QAff7xo5qeTHiUA/iqoob1X1pd5+AMJ1A
DUQi1X0cwkA4YjL2u5YCSAY273FIGwVdSob3LrMZW/3R8Y6Q9JmN0lix+3jk
m7LCXpFOp7aBHVBL6DANNnJX9v7uosXNhzAfq7CXEz3u5sUbuBiPzWPI2Mvv
i8W/4SqCym8M/jvFs8hNpaVG1UebucUdQmooXJAyWgZlLj4JXtzs+WS+4TF1
LlNe6BJVUyxcDa2J+5d0Spu+1ALyIIinFTdbsxgpdgi9enFPqGfjg6ewoQRO
0htiYQegPts2HwDx2NkNIW1RePhcpvFglD2N9VCBjSIt7Tetfu/aFekcPldS
i54bLoc+juInXN83/zHS9NbDkqTDI15zi86QXqR+vsWhWAS4qkVNOmHDNWzv
ngm2/6o/BTLEywZg8wHKhdSayVAmJnkREmDlALwURR0RNERXb/JdTlVp1pBO
rkbbh7jyvqboW6ZDBRJRaEmSOthABH97RZiB3M4KoKR5VGFSuqiXvmFg4IUG
fdXT+ZmbMpQHQv2pvil47ALMkJX4owutv0nAyZi05q2efbh+FPHfi6wNFcXH
iwkcNRcSsedAD3G6yVehDSZraWfm/a5r9s8c/5kUpYsLySVUk7ggozcYIuvw
DolTBFw0glVVA8fEaIGNJN8asSMV2eNwZpadcPoFszqzbUutMMxl7RFsDnbN
Txhz/jZcfupuiP/fT1cdExONzLSdMSCdj1FE3Tn9AV8PFF8zumDgBuYZE/2C
1lGM31FsjXV+wbQqyYqSHiZLfIp1ead4oiYf38VwEs+Q7bH7hmDUEQqfRXnW
bpu1HEhY32Bu8LdEsPB0C89n+C8YVlEHBMpsWJ6l5PQP9LlEoMEfKBUB4CZS
lRoh32UW7/GAa92pQTiBSCC3/KGsbUz1uh7EuxpSYf5fdMPl6+PGpMWsERNa
ZNpAx1fEwWCXVP9qdHQ9uOKWVzZC30TOrpRGQstsC9IqnNk3D8odiHO6sams
vNszVebyv4+HXjWN2fjU8qrGY78KAwS5sXukbtFRbXlZksEFdsE1pH7rjBDV
xzOj34sz+zFCTr14aVJ82b2vDqMBSW5jRX8Sla+n8+hyKCHPIFZb277+lsdm
AMD+OG9m9JOIGB9sE55G679KFzbkjKD7ZKzx/z5RIpqA7mZUhjygqW+e12pq
6GSq/2VahOTwydyEafMrDa4LIUV9olsiAO32v8Xn1nhYVkUxs2E7RAMoLX2I
/EAt/1NtbtEvH8dXrEBc24uI2Np5JIZEZgL5IhaPCjsb9PYDt4cHzWEZY6eQ
eFaBMp14Zlx60lnRmKsW4OrTsG4ld2zjpv+xbnV0J/LLDE1gzeJobNv3JQCw
0ehAFv1t2UziF6FA4t/nN4XAFweiQoyXRdoSf2oSvpe7ZuRJhwmReLl1xcci
vvpFqRma+9Qbor9ZwKIzDnGROa81lj8lGl85z+maVLmRJLu4NS1L3XhyVCS+
TLIVDTzgMDFrvUPPnnZDFD6ZtXVUliMvnh74wNHeoUfjduMJrVny4iFFGJ7+
vTtirJ5aWfCcyuidNvcWD1AB1hgWgXJNSDOKYVlQawTu1y8JWfGTt1jfW54F
93BDeZMVBD7rPuIuswmwR4Dgc4QylMwPNyYcNxgpWRU5RMk5K4rhxhPVXQkB
Y9J5B0QSNVC1IIiiJyDEW1oPb196tE4DtWHK24yhdhEec36ugSJclFtSpQ0p
rCEQRLC9Rn7Ts41Yrg02WnNw6JotD6bHu5+MpfD8V3q1Mh+JxNduHHKdDQcH
ArjW52i3ivwOC4nL31dUpHfs41esZ2OHSvme7FRCvvLN2wh68hgZsHn97fqV
SU2LNHY8OedxER2d6TISBR07Fz+ikeHma0hL9SlQ9X+bqMC1nNCoq8O6rc1d
UCYfGkfRJJLuu4DZ+qkTLl7dlIFC7wa/94A3+lwmyMXm8ohkTsVRVTTbMx59
yO/2o33U9MhfZ8Rw2sr/qltDrpT+YxQkbV4r+depO+5CDjp1/jVDNzo79iWb
XN5qRuEwGNN1Zrq4lmM65lfoOtNJzL5AY3OLSuvk1Yf06UjiCh7mHLLYTBVK
qC15mZ0tK+t8NjYKZnhY4uefB2V+BnZ3b17xAvYmdIwMxL4xDuTiKYWrETeb
q0XEG/GWfR1Zk6CMF6F+T1/SoVl9vHMjVnN+YJiVPXVnoOuzFRkn6RdhoA1D
FGHvurW6EEgvTatiZPA9QOFSGPBkbI9Gima05NUTCKy8wtMgmJS54V2N2KPI
Ml9I7ACwncWwpWFa4eTynzHd95DLrbtmCeMObygF8pU+HxPb6+M/EwJO7W8e
HlL3oOOqhtmh+FAg7bWtpS0h8zpo9AyCLZIuA7GY9jwr17dCETrf2aeaaRxT
CttHvt0RjT8xABF9KyRAkb9JNy/7EB7OoJiKHWubULACsowCWnH9T/GgG7IY
UN0j0eNhMRHe6V37nIOKrlytg0I0yoo75OAtXKp9/cq/7QWkhFUaQOvMtd9X
ffwTyKQxEP6PLn3EacBRY0tI9R4bFHe1IODVa4zYkd2SYEaFBJR0aG1P0tbW
bXram1wrF2R9GrNeIT491OHvIvtvIZbsk4+TWTMuq+XRIZmf6LSA6e9C2Eep
iCkMWlvxYaBuTtTxmm1l/Iva6JUixRIeHpvCM0H/VwVVPUoWNCgUYuIlavFR
vHlB4+90Tcq6aohHqMxAgF+J8zPYONqrTb1w3zko3frT/ZaAUuete6GpFDou
0l2b6rL1KThbzRloeuEnq1J3nJF1+5Nkm3VaTSwbkyZvR99jCDjShRNWy+BV
qsIyaCNF7ork7AKsl2Mz86j6EGFGLz7lAoJU1Vo+0o84ovscwK9m8ZbvHE/x
NZIo+qfyYdfOvGmrZOUMhtCyLtEFa4FkzJjpCX3TYC2sGSYmBULRZaZ1ZLlg
m20PrwP0uO/EludN7nfaMYS2MsKT0XUJdjq/cmVWlHcRUwe5i3QMxCpewFJF
lV3dy6AEDt9mRgkstfQxWn1g4POFkwzKUkWTp/85BTNrfcEX609EMx6qezmu
Nv9onE/cJhmSuXLMEPC6pegMQI4Tum+LSM9nuy06vVd6YBUZVtfUtAy4S2Dm
8ewOmPZYxL4mkDgkqV0Q47Csj7L03ajv3KgHiJsMoh1yGMtPF2b4KTRryWeT
bwPGw6tvARhuEV208JQ9mLhgQtLb+kApatxS8JvcMyMIMhpvtBVLViMeZIC6
KCJ2oMF4u2DUtN0uH2UoIFPqC7xEevOIHQu9jTPOyAGyN4RygA/Gl1dgFEXS
TZ7zlXtIrTHX8Mfa1L1WMzAJqMhCibCXtvW3jSVPL/Sgr1mR6612Gx9fqZxl
Mu875OLlvu1STwfEWFpucR0yoTwlLgJH2kw8HBc2+pIbdAp86KfBESOD+Q8v
u7vr5pjH0Loh0AZdikn6S2Ez6W7ZDLfa8rBQl+RtsQMwl4KpiiK9S0+KMUxL
ds2WZHSXEOILfdPElcVV9poJZHgA6cuwlWLI+xm6OomWOyK2BHp33OXYacGR
mqz3MvzGFnmdD+Yi4jclSXAjJwzruighF75Yj92f0UqFIpr6veZnC6idqBF+
TwdmeZkmJ++CZmcMD94nzhQGHfLA/cElDeyqZihxPe7SXd22QwCwI4dAAkWn
3m0oKOT/988fDM16yGd/ni7+kyO8CQSCCTFKQCRP02J1Jfye1vqs3knRcYPo
7ZD/07frLGyiwshjLSXxS5YJqm+Om79pAUtQ3jEs4rR6aKCiZE+yIwQQoKqe
W6Wd2i8pFh2fBF89BcCVBfcj8DS0CDVpyp00zy6tA3RE/67oI1+nqnzcgM+J
rxaCWPsIFL9eSV1l924MdPGecrjxcd8ypy42a1mrHT71TRjlbORh1IohTG0z
Da+0avhD2mI25QHEMfQW7KnfkXoST5PM+ebZ40EvKVTCFFYsOgn0yRAXEtdK
YXXB6+UsQAGQ7TbSi1ZNK0D2RrisBmEGMmxyOE4wcZELI+15mbCceP3qH4dE
vBmHdrTVBusUk49Tf7K3vwMP7j7im9bWJtph4RWTI9SYkJ+uP7SdBUZK0VqQ
zbrktqkUUAUPczMX5ez3kqdXov0nqGRDXmmLWIaKtyXkChl8FUsQrHj7o4IU
g3dWv5rT8hGFq5JwjTwQfM8Yz+LLJYq+Wc2DjJMq/YqFL1Mw/WeH0vUTMt8a
JQV4U8WzTcAgS7uDiUt7f0mntVAigI5+5++PQf2nkWkMvrj2oGpK0RMt77l6
VVaUx5cUwLLwltiJFY7iDIbo/4xSgaWO9g+HhcDNhHT7MlfmEcrmJQEH4t+h
VzzmHEYZKpjuuEmLouRXKYXfReFk4oeWs5sIIyOocvpOArkyK/GojF+mbjFP
D78PJUho6d3gHAde968G9Od547W80FZzm5ddAOyONto2qi9688uTMJOulVW4
dzflCL5KXwX9oagYkzv/WUMwHTasn4+fditHz+2LOqp5wJwavjrdvVu72mlg
CKLotOhPdwcD70TF+OgEkKskITQU8C72uRADlsNWEnLaXSvyy1k/w+EErmJX
HTTm1kb53orvKfm1Glgy5ttV2IzjUT4gImnf0o3a4uxeEK+uJF97Zj4VDUHN
SJCwixl5fdVordXIZzY5IOrddwpbdHrj/gu8kSHNWehx99M6gWTTQWdezpPO
pvPbQ4tu4u85j+gHmnTB3ytqKn1Puw89Y/a/jehfOG09wtWtTY5HKqaFwpnz
haXdLZNUgI/3gjRHv4aTY9k7bn3b8mAF+bi2avFFkPTG/e66rzPG0zEVu9jd
swkoQaiG4OWpT9nYuy6pOdyHNJhH8LV07g/49D3vQJ1r3FqStLTcKHmY09cs
5re7hmk/qMOvxGU5Odzr5Tmkkc6eyDtoKzza5isqwrl6WaKGmeVKvt7YdT7p
0aTtsMtjJEUFw2N8fD2DTWM4wLcA69GL0tFI3gd2ynCGl99eAc3WSMTezXAD
L+dj/Hy+Q953dT+Z6Oc9H664IZEPQn2m/omA7eC8IBztHhJA+nVdg57u/tWN
QxOoTbW6Y6iy7C5GLuV3/5LeWMVWnAJjAVJrwX7GAGokCmCuoC373eOYak/s
Zr2LMK7X0kB+vXfE76keJdhjvU2FSW6bG4E4jr5C7/GrndoqDLTLIurqbyCt
Ahq8fa/lfWAtonEw8f7fBYY8iDhT4oRKV7hQrH9BF+ZYREzDPPGt7NBg/JOS
/GAnHjmd88HXvCJBoSrijaOteDSUIIg2ocF5ROIb0FDTq9smwJpF8mAgJcxz
4ifi267RCLi297Z/wwCdlMr4/9pdxDKvboTwFUa+vcV0Pd6ooXYjN143mJsL
vRqZqWrdYLtfrjaxI09tP2MFxZjAvAgRMHVRCqWTDH40FixK9aOZppFlPgcx
inh7sezsfe+akcL8NmQWFtKBBLslMzCohGAVZtufWYU2x0pH5zS681AqYdrl
XpC3xu7G5DQUB6b4P0zzSUCChUqUemIneNn0tHck/0xEbucKH3ieL8FENQBC
K6b7XSoUzmg8kzWeIbPm5QbjOG63Hb88aT8eLI06jYmsXzl9cxXk+Ir7OP3y
1dxBrMOUxEwM6s/OCGLTuFhAarXp0MhAWYhVqBic/zB2epBDod784l+ixWdw
Ue8LyS8sTNBeu7GMFFF2qkBLt25/OZXekMrxhsf2FR66z8NlMvUGF2k6b9hy
txgBSBhvA8UnFzbftmo5I6Vrh1xD8L3cuz39FG49ZxQ4dmr7dJd5VyRpNQJS
IW7RjOPJgsJdUYoQujubvj80uhXm3T+X6kHRbeDFoNfEbjdbfII+yfe66VCL
xftMMC4S3/th9CeievYCdVXMLJL632PbFip3PPQyJRgQW18wKwHHn72s6jBo
yI/Ncj37amnr3i6wR29zOzRzF33WYyzp/ukQADmDhAp4Ka2OZQNnPBXhf2kE
S+0zNHu+tRfn6Ajhp00QeO03lt20T5AiB4aGm5tctgoZ0MBSjcotlPp1wyBK
nXwamHJJGJVyjbANO9wvhxPrDxI93kqPNJElRwReEb+tcRtR5g8MUzcQ0z8t
/uPEEJTZhPS9pw3/WW8g6kHbUeJfx6yVQzZPtJiqoQ4waKTrN9CFL/0RsBpL
XmbZGjETnoon+KW7SxRe8ewdgPo3EbB//HuJRtFcER4MAzVFU2XsYGAJbVw0
OB2NY1xIww76fI3f3BeUw79JHFmnS2f9RpHkYw5y5ndaYwLJESFwlrqgLkq9
qt/8mCzuBSwcvZKo1xbtwX26197Fd2Y/yaf9bQb8qDZad1wicRQfufyKjyTo
eQKKnxPJvavaAF1L4Wi9mBD9wlLaPKWuSrO62S/k6tUSNUlrdKPlYUsrDeij
y5UBE2+uhiT9YFSYIZQvqwWre/zpwFn0U8SdYPJF7msGiVdACGvegG6m6aB7
RKPq8qoizO0Ln1vkm5El9dlz7HXSE82hm5TW1qkvkNK1srs6ADB182Oe3kZh
c1/7Zq/tzXrQOGYSZrkb3umFUtDjSt69guL45307QsUaMLOL/OHOyDDsP9hh
5eBQ5umjhGtTzjlFiSCtj2TIKarNSYns1nDnMQlznS70FCyy0Ui1FWfU6pEv
pxe0mXS1Hhpg8pzFuDp3LSn8Fpyzm6sGUkFFroyBQfs3Z46f7BBNI10cSixl
RW/+yHcvFcX7UOCEq4ESv/FaVNJnIV2VQWzd6nQYe9EgVVbC8Y7FPUSDjjTM
KgZmQ4rrIek2/ehL/icZAC/IkncmWbuGJdD0dGQ6vRcFBm9pNkneht/fKZOq
eitDV9fBo/AKKHCEDGyifj+h7OoJVmE8acNZ9jqTa3lIHQpmeUfTOopVdG51
rmsuNsfSYcoAWfiiv/ERtX/Hi0PXfliVaLuY3t1bsmPiwJjm05B+tewKGVzo
sFCDBVR8n9XmoH8EEIw9q85bnwEgjcHkxO4bv9OnTR3kF1Eksa3VwFjkpJfl
uRxx9xPs6J7iN6F0AyZ+GGOWSEBuQ5CmMzWKPARyo10IWMD/KrfK5LUqffwp
sECpnoha5N7eYl+VzJoOFaQG89Yp5INzrpkFNm3YFSm0zXO89yvdj2YRljF8
Ij7VDac+oS0PxnSbnByhsIYqSuhIxZOE9rmL5JkRPMra+LWDXG+1iDs0aeHG
aP3vJuBogWFeMO31naJ8Kxh7RZy58U9YCYw5OiKRjOz5g2lf3EfSfR+wmgiI
JVT0QCkNklm8uTDIC1NsNRmHDGFLNYV6NPouZ3zEj0HBebuCtZ0taC2V8yRS
GLbguiMSU2Xv5yDe47JEKkYTkbu4DP1xWBNgtgKsmf9oamKlWxg5ndsunlB0
BbcghGvgmcfGBgfnhnVuEZvHw2xRfVAfelJKM/eSP9UuEHBWpWMZ5qybILGU
AJ/N1pkga4FEEdtHV6jl2dtUCaXNSQhesfCpMToXlQ6Q+/3aHXWMXOVxHCAF
2vpx24G0upQTlXrdb98CIJ/EwLuzuTnXjPvYNnmuV6dGnlrujtwHI4qIUCSL
/toUdIuoIrfY99Bhe5SbsuBr49hu7PnsR5HFNtn9AmX1l5HAsn4mab/TOXPJ
A2A2DdNOqVmB4RZXQtUxjoyMmUiZn2h0cw2IrxRl1V0cZZCnaBD5PQaJVp5q
colCB7KySRXnexU09m3p0ytFvZ+H+tQhYHelw8eJ/7RKMjYJOAtEk5xczKao
TcvUZp5VfUr5Lxa5AQJhU/DfUDxdh6Y+uGin58BtSls3mqTGfSB2lDnjvI9r
mNJ5tzH671DOq8GFtwx0ejIb7D/96AaAilwNiCvgm0bVOM0szwKNz74CFLF5
F4peZ00jLnQ7h5wrrU7DLVRC6V/Anh2QcLQsjMyO5PHUVlMqs3S+Fcvtl3WU
8U1Qh7OM8qJS/CHsT4i7xTJrhLacewMm8q5aV+6i/LR32r0AoP5Gb3iUL3gn
GWPFpM0hvl/9dFC7RvwEsZ/sIpwHwQo5LXM31In/nyCQCZ/zAmGLBhCDjBcz
5TkcynhuA444x5rMiRTZOGWUNu8qnwL84La+SD3haHW/XOWWTCm6ZftcwbvW
WlqCJvG/eAzPTZQof/cGb0hYI8ktJQNNMk0qVkIOCzvgWkX8u4HKmbR87ZPD
4JWtNv39o/r3N24zmzugZ1QAtJ1DFqOLtK2dHmWfyYQrbQunq/vDs1SWi+Jd
SywqF6BhFU7Cy8lZBwnjDAbmRnkctH4jdXXiA19i0zUZYFXGWcCMtskr2P8A
VwOlyYjijxQ0c1njJhVhmbfxGmKKEzj98WbQmPJNn6lWYDzZWiOwZGQq9YvA
RzKILub8PDct2ze38+nrzuNxyjYfU26knZxzdlp1YpjTh221gsbZWNLZKre1
yARUn0xGQRbK0dfZmdXP8L8P8+/RAuoMbgZ3QIz0Rshm74rht3BbQ9W999kH
N1KQ+p9EGJ/3wpYEX1Cg70Bs7n4z9e2a5RY4uvkcS2Z/FENeDv+T6BipmiO3
Ta1pV1d8GwW0DjWEGE3Wk/+h1r+y31prInyk3MMSZIxSoeEr6qQZTcmdqydX
uvIH5/jgFhgmW89d3ZsJENtbEcmM9DX7Ay5CstmUoZeHn+oZMHiUcA/Za+se
912SiDhPeV/ihVyEjkaZ6PCAFpshhgkAw7cjimP5Qc3FvCdHdWyU/G2tfVik
6mmzxvnl1NWxmDuPTWrRwBF99BppbBrTGIBCCf1PD7WZxESM7rFnEql6pdTZ
0vnhGJTdyXMKkQnZPPIVS9jMHyOgXZs35j95ljO1IdhAl00qWN6AGiV7eQt5
QqtEW/e2AP6K5XwRhs+zUFJk5FSIvkNNZ+zs1W+B1f93y7prhmXXDx4wSqoJ
hxGqAfpLrHxaL6l96QK+dizNRlxKaR3GAgR6nHcTabHU8xg83C2TYEmER2Y2
JHyYb7fnEqY2MEW0iuXXJ8mT8hbkrvgXdoCRrwFrKv6YVt0lbMQfdFrvv3xX
gh2IO+aZRqXDUmnxr/ObP9zYXUvibFytmucZt+xVLQeAMKrif7UAInDydWEA
/0AMVmwVMYOI9XFdTf9isEs6yyEcH1bTBHA8jlgFLjcwrV6AbB1plhXln64e
lBZ+SA87mbRVCjR/aKhxjPtjpcAaAtep41ue8USi10sNYpzxmRSRZ2JJWgKJ
A4V7y4+xFvGTNI+wCXtHQUtWWHhXoSb0+3icIcm0O7P5xH4fYUi3J4PvaahK
Aa8V9+mhQmdC3NKA4Hoph6yjbqy4lu4eY9RxjJ57lnp2O4pS3EhlVsR/8yg2
DOTXG74sMRNoZdkncaYTUtvv0hQvzH8AJkfDXWZrw5bzz8CachKLXibvs6cG
UzubgR6nx04dUezAoeA4XSD71X09hzkp+yjLIa7AMV5FfRsWyc1wcxHkGC++
iqN7SedfyqkgU4r5n65hHHwb8KRqv10ycJna2kcqgHp4jMxmewBoUFjBm1bj
roZZNWql6XjqdlJXHATxwn7I1Rn2lXomFk0jtknVvXpiFfe7xz0uMRjJQaH2
C7BD1sVKFCzEeBVrvNGv0NlR3p/pg/cfSrdkv4TXt3XOJSGDW0o7rk8E+ftQ
dwwj/7ldODaFh+ArUL1dZtpGWJQIYw/h7mPN9XnsdwDXGt6EIj3isqn1YXjS
UMofUrlYJGZZ4j6yPLP7VSwrhyr4aA1ETmZH4i9d0mHjCbyvzXf9LyUKSnAs
xOtRSOaUOUxBh8VzZt/VCNDZkjFN+tlnEuaP/oqNw1rCsLjmxXGwVxNq0JoD
ZhYfesHyUrWF9Ivo81knLmVql9P9pylfaaemUGu6uAPYsAIf3e8/dG58agbK
n6ldGvHjfN+nfeAbLTAkcleRrdK/lF0UBa4Pd83QzPcxi8BC1/v96t2RMyZ5
m5nPOhpTx5WJz6NCmjTDuUX5/CuXxzC0hny9i1lt7xHkBkuHG/moLu28M+KF
x6uqn1OUotGzttqEg/0Eduj0tj9rdRxGe7HTAYwW6znD+dq88JhzzoeB2DM3
BKA7wxMBTLBnJUDl7yBagED0bKv9lfZit0aMJe3bBiWUjk1RQQiCxO76czy4
yeqqHn8ns9vZ54o8Hbf0z2Jc1GSxkMWM4l/0UM6Gj7Ma+4Uawq7WeZq7ZN7m
KhZLcX+5N5U5qZ6L7RssrPwdr43Gw7JavhHqGwF9M18gjKtE8aIwjrmX7kPh
qspYLnISsmwfMDwYnWILwqwiW/rs5YXxuAyPfd0O0w0xUt77j31Bg1ytriuB
zVoRhDpvLjwXKZYxdcL+03vXx3kV5UGBVkqVbR6Fvc9H4SOokG9F04PO4Cvk
yOh+v2Nl9xjo5HaHpeorLMg0KB63ANWAteL94mlTNqoKtWekeRMzWNoYUOri
K2F9RsJ1mUeYp30oiIuavE5VvfkYYJUlikh3/F8veKS1tQhnXj3F5O+2QjhV
N9PysGZ9xmHb3KDnLJtVOy0aFDaOj5o4+O061haSDREe2O8LgbJuqsjzAH9L
Y6DeYmsFAZK7teCMJYC88ANx69MhJf1BbBaDdb0Thp0SlW9JMlrmJUPtbZHY
yj+KOUxUB/8QPczXhzAC7QcBUOp8yY8mgkAT976qxXA6tel313WSmiqEM182
0bOyFLQEwq0rRLT60Ijf6Ok9X63gUVmK/eI1xhFvpWMwchaBzRdsPs/Foqcq
a8CzL8h9h4F+P+olkZDKtb7jfhmpfDIShJLKi2LrpXNDd3YxvJJ9xGu+47oZ
TGt6y9AczUT30q2MgoYOLnk9dszpme8S9f4RW5O9aXH9t+NmRPRjd3184QCJ
8+AWTE4/dr931kErtmZy1+XNh4OeBCCI+n37wyme1bOnq42vEMgzbFrhjEUr
s8v3TRDylxrAu83EA9csEd2DN4dK6Le163jhUCyiOHqttOCDMEGFTWxy4nfR
KA3KE2zCEfWh8tiSLN/ecx7++tLdN1fJWo/aeAd2T3pMEUBXukSg1lkM0Omj
5b/qoL8aw3qOC/3NXCku8fuZG2xqOYE53IqbVmadD6H6I1jQBkkJGYMV9OH0
iUDVxF++EyNHO+OrH9SokHDxPe/tnmKyYPqUrCNOjFELAx8WjtBDz2StAe9F
kSpK1s6ZeD8/LkX4/OFb07n90rA3kg/4J2UGeh3JMpSupULxaeNVEo4ONYAC
+5rAb+iHJF2DEPZ+AG1+CnywJmJ7r1aRKzKJqLZzzIfLqao/Sj6DcpU3Pju6
g/qSwRorwE3vuLmJqXsm1r8H1qXS3fRSu5/Mi+wk1iClPmKAFTZ44cbNxj+q
2QL9TVIr3Kgze3DElCXssFx3BcV7NXkXaidg7P1KadmgBOFP4RXshv9fDS5/
bjLId8DpPI+c8JCmrPPrj1AytkBfu5HRZF4fqhl5FDp6rPiSTG62WGy1R2Nl
HTrJoweWTDI4m3CfPmUzycgb1sCZqHQavieXCtZxb42Et/iwUe+D2cIZ1Zru
rfkTJYCkAc+OMpZ4RVQEE3zUiUvsq2aWA/4FV67+iukXLDHYMGC4ZYqHpHk8
2rn4yoHXEQgTYfmFVnYPpCFVMScor2NPKYw9t/ZqNbEKsGNdjbbKuA1iay8X
oSvuttK9zPKy1heymO+kifmUehS9X+185lB4QYLzol82Y4nChSAOoRiZxb0x
AjfYhRatAimGarcd6Ztx9F+bDe/Mim6gW5vzUDlE4iygeuwf6EoCXkm0vLnt
Ju5879vrNVWOWkJOCuylrcgYVsaZJuVnIx91XZguBvvgOltbTytCKFxyUOrS
A6OMjLyAhs3bsKtPZO8BEJIWODYPzp8GCxJw41d4h6MxkD4hz4pc9ejIcTt9
ZHP2la6ursmZp2guIuNi6eCshrBkweRyfCpjUHxzfKva6OJpjPUeJdMEWQtX
gZcff/LN8gFPGXeCcx5YW0tgX8NxhBGpmjyBFnqo3uAki1Kbi5ZzDc3vgGzf
6TYPyXlv9UtGZmk/LjhvQrVd0EeRGHhu501Q/hhxDpbN1Gqtch6mDCAEim6Z
+dJ1TYz4DJGzRsjxFgzBTshB0HSoRcqyJu5j6UUVN6Nqp/qC8fnOvBga4thV
tTuvoX0bBle3zWduDGyZGAQgZjUYsPIgM9dP37y1nBE0wOaQqf53YMwAA+g5
MJ9o5ODTgNrKN7ciYIyhPU33CuTARk8MEKVuW00I1PsWa9IViDf8U5p3yUAJ
95y+q+kZW+aKJ89hwp3Q6PjXY2nDvTSOCJ7vkGqGhYs/jZDwxm0ANDGNKYrm
7D3kSZzQti3PDT92QPE4l83bibm3980n7lDpySrBHVu5wrjy1vx0V07GTbmi
s6gPsC0dEB+uAMy/utU8pXGTJeeahT9JGYq3WNjJljKpHXfvvutPESFmr/vw
0Ns3ifRQEtLcznEPdhbtugm3WivWiIaarbJOgVsWFWcWEBiGeL+wCAiHXpAN
e/Ao2x1B3ZGMRfi6socpntzf9FZCIFi22NgiJBrn+j1/vLe4sO3zp37WLZX1
quhf24jnqz5KilVmZd558+LNu0Qgw5mDErJlmzNWzHGws5Q5ztZmJ4TZsnyr
nXhL2gD0gaigKT9feQouytSH4ctL3szWvTEzYSEEI6nNSdFLpQjui5ACUbX6
jH1Dd85tHFPImlKt7u4Qz8CSRGmeMce2tZ9taAoqHIPHj9HfUUf1n9IPOVJi
OR/Suzps3lF3ipJ3VZMGXWoX6uSIfY96azIIhO8D/Vv6/TrNQgia8LPpCXF9
Xw5JqgizjkVMf2QCZWWTPZhmj3XlGuYWhWXK/YnMP6VBQvxpPGjcJJlpMTdu
pbXCTaT0QxNFFNPae9drIngOi8hF/Z0RuPUixwU2bG0u58pPu3OEhY0a/TTp
Rd4MswrELgRVzS0cSxboUbLFrTfEC2GXw9H0xb2FVEEFVUAW2pUvanpSyqwO
a1+XKcgOce8uA/f0ItvDAboWDmbFhx070hEPFVjS0gpc3DZ8Z386nbh4+ho1
Zv3Dz5vM7lJPPhvi0hy3AQibrWbWH7kVuRPQXScfL+zL3atcdqPrUclUMHXu
9W4HLt6PTKgEJ4AqPWFiG2e6NEwd3OnrwcEdjwnl5h9s3YWK3+GbqUZ1SHEo
muA+NrkG6dyU2xrEY8wfA4zR5b4LBYW/he5qb7jvYpXa2ZstlkS0+AVrPpki
jHlI/GzXN4OGBz+ozQYweU33ctV6svuTvMndOS4gZwVFUDwKP2UQ3qlWednk
pRsoZO5Otg0joIrb2R0lSmttgCZbQopdXGvrfp+5hmiNnbGsiAd+6vEvfPsr
e+EnJmKVoa0YnMUX+mtEdTusLW+cuVaToKdWGXyiXxR8uGphtmIFI298nlB0
59CiHe/Yjdi7acfbphQYR4wZ0ODcEo87LAMisB/VVLK7pbk4RMnTYB38GAVW
WQ4PRWnMHs5d94XuFXiqAzem1XlUMIsOK7u5OUfkwTqfENtge5Brwkuf7eqt
0cQ2W4m33da7CCBKXqMKh2YnJlXi9r13HQHtgxnC9k4d5c5Y3jtvMc8PtKPO
e36UFXQpgSXo5bzZ/0QQbvCZzefOD5PHbdScp3wR+PRMvCP/wpJYxjw8tJD/
Ym9uavuTEChnJfHpyZPjawkV+Jy53qUh4INJ1Gp/6hnrA2AkS3jBUYLOiSCu
ilOk5pMqRFV1zkm/XVxFk7+DTx/EA4wV5ipaQW3SyBmR8fmz7DMcMgJxe7/a
HMijL2ykglJU0xySIDLWoJlpayBOqefO6tuzoc3o+wG1yNf2XyXpWZlro25O
18kCz5EBubUqrrV5GpRVT2/VxAzdCvp6sWbXvPCMZpKb2KWUvUiIqY4Ccl1h
kHfbWjd4NFus5qsZz6LVn3dzDu7UFEcLIWnNNfd40fz4WZ0F5FUyOQ3SLYm0
FylbM67Ygt6c94MqZ9wKmv7YEtarRW0wggmmuYiud4u3c/4zIzNr+nNh4sLI
00Ngui38UQbevkKi6wYOwwLVloa60mYzzleBhQ9d3Ctq8h1FFg4VWf8n16eu
RKbVeWLy7dh/rWn8RYLgbrP3DwOAt7ezECcF+ubvDG3e1fEEw2ECoeMxqeV6
w0ZzIwkLPA3T2LlnWSBPulgLmF2zyAwQDxFYdmnWp627kiQizM+J6utCgrLM
z3PGnTeLtfFTdkibZkfPiAj+bGukMnTsNttVu9w3KgAZIytKAenBs7U36KNr
6TzVR8jdnPbMsOxHiIxqU7kHuUTZlMxMelEXeeP4fMiE+BbmzIRwEmncH8NA
klW/zqjEn2em7gHSLniUmVkntf1khPsx9I4LcTox2f9IGpXi3Q/b4e4IFdbc
QgJrFRR6Rg0koeBfFAG5bB7i7eK54dDx32JY8ZpKlnVe8677ULptZLXHoqgY
hUmHLFIwxsHesf4x47KijfdYhZPZPI2v6RGUTqXGF8OsvZJERnt1NkZuKdYX
lMRLBjJ0kHlPX6lsNZYcxeSrurBuepkJbu6u3i+mPzxXrPKbMPDIUpbxFanh
I9YrXvo8hLH9+s5X1b52Ay5XO5IE4NFA158AcWvSEynLVzFfYkc/21L2g7bf
BGNnjFSN4I7/eonK3W1EKA5r/NO0nZPIdaFzhIX3NMekPqfQYMDSJF+OoqvO
nEUON+xwhOBpE92wGY3wtHDWwJ4vVzmpozurNsbglH9A21qyG6GJe3rqCJub
8OTS9CDTcuQq9p+4bsScHuRCKD7xqN37tJXQSmUlZiWcNET8Xcufmg2JjkIY
V4Ndr9XcEFxcOMrpURx5HcT2qJXzaRFZxNDuWCGOCMrCIo80pvslBfTuLu4O
pKM7qcvOBEPG3ZSzTbTGMokkp0Mz5wWcdJJLDIAh8QPxpyc3KLspQtYf/kge
A5bjrBf5TtW+rGqkLkojo6S1Zzz/fRwA7UhmVKE61nBWHtFvX41/d0Gm87LF
WCz6piIKbgpaJPnP+dD7m0m3RpRl21f3+cUUo5h0PZnLp0yOPY6ONRJXb/PT
AOlZtUzsCx3yyUDa9deMHlpsV3gnVeEaKHjm6QtNd/1Q0NbJESp56jetzAq5
AVka3AHc/AdJxBdjbrTY3DZ9VcdeMLUDnib7KKxIqxM6MCGALz3ngBq3Ge8r
OBY/j4mI6BG/AMheNfnkebbX4QSmXKxu92mW7DmrtpLOlhKKUomsxjgd3rHR
0cCWugRK3fBF40nN6Hk2jlBCbmi/EIglA0fz8OTTYgMr6wdMGkRTkD36rlld
/NyXouQZCbIwEhdzCnffDiXCrBlOPf09wyI8Y+BqGdcmXtM4YoyShsueZ65a
pdZu5MW/EeMtAgY+miESg3BE9mVmCwQF1r0rKU1WdrDWX15KWlDUSXVsro/d
/EKQQsMopXgwUTumDGr3CCXL9v9rV7IMJe+QRu/cvXAd1e6tJUd0Fw9PTWrb
MHpq3TUKcVwLhkfe7D3q9i5Qo/fNuAb/FRz17KX2ocIN6weMEzazdq42g7Gn
h9F1UeEVW8VyVQsubQK2v6pF+5DodMxF8qs/sP8JayexnZsx2AnuJqbBLMgg
8ONoIeqqTV60VjiIMlrU4X2PaihmdMucp0T1bnCIo8+rEn5JKsRg0J59SryS
m9IoNs891my3JKOToxL3VelOyjZtfSll27iEbFFN1haNh/D4Jmb4OTL/8mOz
7cFsqFw6v6oR3GT0YPKx0bNLfeS655kOE1yJ9ew7XZoOXLWrNk5ElP+bZOSt
h+ixJoq+8z/iDsFyrsc6PUPU8yj10SegZz2w/zNplpKcCwbOxEVAsK0tOgO2
WhnZtevTm4dVEAy8gh7R4sSX37HJqz8YoFN45UibYpHEZTs2S+RQ9YMFqUgY
R40KMOBLaI3/ILf0G6s1CRRwEQQk+kyYFncCTSiwSUyMogIWT6oJcWUCQazG
lrmgRFibqDEVZjcHvWV8XgWbLiTiPgrH6rcsb4Y2OXkZHx6M8DJ2Ka7MDVgm
MC9tXJwC1N5Z2hU+465sPTuJYdjzhwbbYzvebhwdyekpeArwPQeKyhxXzxb1
xPAY6y/lzUcFf5QbkqO3vNfnpEonTcWodqQjzOHdGD6Lw5o4kxcXBOrIOn39
IlR9i5GnsSIt2WOJGgXpkGjnp/Y+Xsh0fc/Mp3FSGF8uMPc4TcTE2X7t7GMf
YX3AndZ9YZrXCK4VBxLicXsAB6HKfO4MYWRZlTdgRkK4Kr6whHpI4MJCncxV
BXiI7Tougo+VIIan++s3PCXeNARq7rA9lV59OhsUM19j8jqou2JzhG5JoU28
GZUtUQ7zE4qcm29meGdGAVMcGDGWHVV7Da0u++xD6mqq7cYcdILIPLa/AjWG
NTr5J62RPZRVaij+MQo6TLF7SNoyGK69q04hGtq/WaAuQJfrlmEkOBnO3G0u
Ez2Ymh4XoY3qM+Ef+cvLOJT8kL+RO2xglMImRce0ycShPhrAAp6MqTjDEH4b
lftC3YbqP8dyNjc+tGBKtQynh7y2Drq9xpdpBc7LUCwl0+Z/d6LB8PJTXQx/
Wl+9CYxCyHTpAnXOkYnz2tlV+K3jqtyKZji5h1DuxdfWq2LHra9gIK/1WLAh
K40ROk4mFGaNAaqvi46yvX+ys5OEczZmZvNbgBNkMbjV2lQQpkkAVpwOIg/h
EIzwcXow4md1xbPxDpF8gcIlaymIrrSKqQUeQYfZOR0A807YvPp10NSVgNdQ
pQg8l6B/CDAbflQkc0O5OauIhQEuDFrlCLJ1CAtZC1c8AMxafBGNFNQNTO4S
8cvg+wGGYFU46Jmtb22ZJ0bNZLnJuxJzfWFjtnyHwI/cL/RRJBCXy2+qXR6A
29Z6niVnvhsNeEUbHt8zmcT/xttpnuY+8SZ0L/n0kb/7QqRBZpgrieMctn3P
8/c19isxWX9ri1GiGK3cMTW9GQ6JLbN41+qc/LJisrLX20apM56e/+UvdPXc
G9BvluXBj6p59y48SPG6aovG/salGQFxTGWOl648Znxv9s4XV4GvAu5ojrEK
gtaoATfFvpFQZbk1pPelAGPJbH2xzevwnNutnMfnH+KXWT5ZJj42LbSo9U+1
bfsiNMaLSi5p2Nuqj2r3RNR9hGoAOdT7gSiOi1KsDFe8kfeNQPEh/nXKZxPp
E8qu9z2FG3gPfer9DnqTM+TBZuSVwgxPdD2Sq9id+jbmZXAvTUKWsySQOhpC
KfX3/8Z+cHtpRW3ePcQZEEpgc207RYFk1stk82MRZMmTeEfN1YTUYaoqFSyr
WPpn0ffKqpc923HvrOv7B6Bzwy2zmn/Yq/KoEgVGKBguinOTmxi4R4va5Maa
xRmdPBiYr3GC4xVVNKgX52ciSX3R13kTAsczZZcDZcjpwcFrhZxIcR4dFM7R
1SjOgeaHsawN6AqJfuvObYtfSer47pM6JD6MS+oBUoCoHg2RAxnupEue/xhE
LekohoAyNAe+6gmjP9RzfevN0EHsjh212B24mrQNYBXliyVxGkkvauz5tLyM
6EJkc+L9r4MkigN8lz+i1ngq4usaBkB9boZQIA4+ZcHBxf6+cbjlrDb1kHcW
BCCcDXwNU/tNJGR5YEkVKfjaEhKDl2SLVt+8mNFlF63tBJQ4gGTJrk8tPvpU
x8ETP3r00YOMbh15zLXZZ5Y+G69ZhcxR4PzO2qfLNMHElWUqMdA8/FYuAr2c
we7FuN/o+y8OiazPcNtupbtKKnFW+sxLg1dQKO+Po6VZ5wIpoeWdZB8wPfTa
apfTbcYwXLaW5wF7eBTIjPE9iwkcaU9939DawoGC1W8HShT615/OrXQfGfBd
Vo8bjRgrsQrUYqUylBqU9v3PyyvFDMbc8bk9VIXXUKGu8EQjkS5R+HSEbihV
zQBeETvDxErZLq8z+TfbwrV3VCe1KqZjur8ZTteYQtFQ34K5nCvj0zkU87rq
6taYwIlUG51Kz7WH6giPSEP5/mC5GMAQbJH7Hy4g6tPUCsUn3OVjAqlw02Id
n66gouqnMaSwlKTpHtM941D3+juBwah6Yy9vRaA/bRRvBBHoXgdV9XSj0kvG
LjIVJHFYWzs/STFSbcu5y6qVOXDq01mBdgrTYMPPmsc0aLn8hrT6uvPfClYu
GmbIItt3IArQfy9WeO6DbPfu6hYWjh9CK5zpoLL99q2+vJrSMfv7eWwItfrv
nfYbr9FiM7lvOHe56Z7uGdbi3EfUQW/mooz9vk115m+Cd4Dlee1LL9RVurf6
lW60u577NJxf7t7QPs/FCCRpz3WKjSN64eTChoVffoqKOFUGeJyeJuIgNByM
DA8jU14Bk2/BKFArxZAqo5tmu6hcEQRso/grQnsSO3zlTdeilBYbbiwGpgjA
uEYKMUAy2aRSCthElqoh/3dlJtMUblB2GVwBayXFsHVlOSfRYTPLT7+5Ucq5
V+GgoC2G4+qW7VYVMhKsNNw8OoFfFOfP3zOkIj6M8KZcmNAw7BfCKyiAb54g
dflETaSaqKd9WH2LK3tFYSYpLHKpWvmI32YXQ3FE9ozzElAZFZyfv3qZfk2a
dV1keW/hRAIjC6j/+wacRdClAskUwjqmZDRlLn6xP1WQXjCqYMqje0s4hITv
GKN8wihZabBClCnygu6EyyBHrv7LDr3Aqqq7GJRc7sQgX3n6on51vXD4e9fZ
2qhvbKroHnPEd1mZGC7kABoxMpnXgDBE9ITw9bszjarceEaiZbyneOt2IciG
JXLAt9IVzr136Ht07mLxH15hWYD1MEC9RMqZPBKWtxhp7YNoFUAASGU1GMtv
mjg51DbSXXMD3gFHeVK4ieNXx0KhfpRwez3mgebnoZvLC6two3MGK9XbnjBz
jwjhIAvYaFmAWpX7+2ApyIZ/V+OFJ3XBuYyDnV5qrOExviuj9IqVVECcojvQ
yS4o/7xtzYptBGZIcsVhAPvVjaMaroPxKGjJUxxfFUR0O4XSYfBCyL6Adm6s
8xh18MsROC8aecwNfT+f5YYiM5H1QMgoouyY81jKD75eit0cVQ3OiyL5T7R3
RkL1RWEreRFkeMxdiExF6PNQ0QVMpE3ws0qyglVa6kiwYoKwANf1xoJ8PsYQ
8BbmzSrMnDYSDwAEfKMEqxJIJcNx/dWi+RIbQ1LLu+un45l33znGFyoj0UKp
qHxqpJvHNmBeemwJ5wmEy2HYEgvKtCzTGIxjb/SvUZp8vOotpomcth7qP4DV
FWI2tnIJzn1d3NPXbA85lhTLs4yYfSGP3dY2/21KfL0xoZBBhZWCTJ2DpMIc
1pRkjOtwQs+0Rt4rLkysinDCv15Pdf0PBYFHcQdApqn23+Phow/AckDLUE0y
tu2gRMUB5tLe2YmiuQk2NJBykidq6M9eo1bt3gcUL8YpyA3591EuNOnuADjz
cuUYPD66ENj66n195XyCYlGel7UNyp03gjMu8yUxu5mkXc6CEopjpiWXsM3/
WbGMWfo445ncw21QPu4BkR3lVO1XHxP36JJH5j1CKtlh/B55cDTaE8R2mDIT
cFJmQRcfrpZFcZxBHgX+YolYeaqw817Mb969ZRDAOdjAKVsR1SNKPbg4q0Ch
KES1Xw9RN3TGV4bDY4P3KsOMXNc7TMjW54LpWbxebzdZfDXeosZNwPVWVB4D
XyYBbPEyZhVkvtw2OXu6R26kxdPiizq8Crr3mgINUDLfKFkLe39hXGtjTBpg
ecfXam3QdUJuowF6DVVZ6/X/B5nFRMoCn5ynEt/RGSHEJPtAD37kloo8kVTw
HDNXNQANLZRGyCIYOwKfE9cPO699l37IQlCRzxodxAjK/GyNU2FErPdBt84z
NqNNU5upTH/CunkFiOwljl5gce5UM77+KOPcAAZLVjSTl3VbvGIqqg7qAjhQ
AIFzn6rLmq/gh9IFtUBi8eGzRRI7vEfdQ+1yuB3uwPbj5726OXyBastlkkDN
8kKvKaYDuxWgDqT/+p6vEAA1Z0Rvq1IxYT2q7jPjzfk7pabZ0sOcZU7pG8lk
qE1h3Eeo3COzSxL/Y5nzk2IW8jDu9VZWuc3B5v3S3kh0Ou/ebr0jyQnNZrOY
+OL/UrSNraL12awOfKgfYcVCjeBQwRmmiSRfem4A4Q3YAbpv0D7cv4qZuPAL
jJcgCgoS3vtQ1jb6c1zbhRGYSZAjdCj9caHvkSj7b+Eyz4pngOrKwk4VHIcr
OQp7MIyx2faqG5QcTDisqp9/LTWVTUFbR8RGmXkTe5X1q6cHmZ1yzN7+ANTi
HGi/893tukGYModMpxgElC86xU9HcLsrd/6seNbX9OScdYH332fjrh2CFLkm
AnCfX5mHvXmSz9zfpm9kikdNL+JqYfHeouoVVshQ0cz/WgAqONTKcBuqPslf
iIHpDxq4eEcJ2XTyYPLxg/TjJPK66kYCg9U7euzDSCouRYbavkXn3y05d7kb
SA2mz1kNuTufPnCvXv7sxF8l9nBow5SmSHqpLrcWChNc67nrNRTSyxQFEYY6
U6VtpsB84Bu64xUH+5BoXoD1x9/FYlJfjlxyIr5fDYejZKrAwC4rhemW3+NK
UprYMKKdAeHFntK1KKUfGl2LU8+i8dzNiavbF0OKbmQC20z8g6OH3pL8tMMr
/fR2SbUp0EUbsoBfy6InZxAyTTOvHClwtQzl6BPJFyydIZ6Xg45wjd63OmFZ
OSiFSL0U/2T22HsDpiRvIzu40up6Zv/g2VDBpLf6f0f5k0iTgDenTzdL6kAu
Il6HlUO4GEGsOVuWQBFRjZWivuXTaqYSvfopkyqHJjYV80o0w0266McGOJOK
t9WyQXEQzBeSGxw9eCOw1IZANyl520MdZfegRVhXGYYbqj6tOFHDneLWlRy8
P24cxO+qB4yfUevi2at1hegcc1aSMSGuQwRr97BMCUlWtChBBr+JQ7n1JhR8
V1vntXsyGW7v+qbaLjL8dXe301E8i3yakxIhHEcjCuuw0s5SiXWAR05F3p8H
kbADZhGDCZecqYNLfBMi6h3iyz/5FfSKIOyPT5318d4rKaqFIiZ+FlPoWDwH
kiml4Wt/FrZhxtakwTwHrdFMJNsJvdUqIBnUv9bFdIEJQ52zQIq6ln2huNVx
U8hcfDkupugyco+SybC8s9i+1gKCE6DdCXzdx173q4WROx5E6nyJs4MQWvBQ
7BeCRTOEsB/jdkz/RZfJ50IcselO6yOJOmMhE0W6ZxwNjBqB3YDgU6sLX69y
V7JhlxVNbzmlzoSbH7FGsHA0DwvykVpL1vLJTZktfxomvTQ4s2YycpCqpAdz
qQix2L3OJCy8QATm+BVHw8NokVvQ1qnwV9ATv3uJ23yI8VQoX0uNiv2180P0
yl473RMsUyvADyCnls95yDE+XdHkQ/h27N6MrpUDyIydxu+AA/hJptqI8iml
ohf8gtyFV7IjkbYbCU36AbIsy2WWKK9/Px/vyN8g9NADuiuSqybuuoQcaYXy
pZce562j2eKbxHkXuGK5a/LhA2PnfDm6aphidUUOqFyDx00s5exv/bsXi0E1
x6/pa8ivM5N5NSFJfDL3ICvkXeuXBfp8gGoE/3b9eMSKCIq+OSRaz/or07KK
nwlNfVX78w8Y11uuloCWBB1g2s5V5qJYbcr9Ktejx0F1A2klRkX29jQdPrQJ
1BJ9wUoZtRZ0JVIaARgNVhHTja/tOSAzInDd9rjRKq1/sIigE7+KNMbDZNqN
f9xxhCF4EGB80O+gfCQULa0Gw/J/KIFRj+yKI+17ICvrrFa6as6ZguuSxVuJ
GomiFFLtH4YLZ7Es+62KUtfB85EKI7/JNPMz4MaVQQPCdH/UFlIZBe5QksDg
hK6rlIYF2hIWFcsQughVGreFFTb665cAwDUeqk+UXxHn9mkeyaIGXYa1z6gm
dXz1S6mesIhW1V7+UEV28e50q/NODFAFduv1RDIXc09ozSnqRpA6kC9kOGDC
SwPJ8esus/GodGtyYOG2CPY04eB0Wo87WslF1TsqZpCaakKPDfGsrzk5uRf4
nE9nc1KTCF8OinW4kif3F1DakuHNK/OOROVj2LnRMXHE1pfzYGqoWejCmIMe
LcQ+9g6rkbKYfJQPKQNRzIYQMhB/Vfkly1XMEIFDi3lqjwELk52RQdYAvXZI
JJj5NiNGTRUdEAGJNFsh7ZX1YxGhDYltHOard/OP1f6CxBaY1QsOVpsC97fL
D0/R9s8PZrBBrrGEZC5xq1YfYLYYRNqVzI2E+puVH8L7vonWDheWpVzQn/1g
MFV4RYTn2KGrzBQgbl38YYqyyH3ItMv4pciwycBovKDJw60z0kIiH2L5u0Co
f2CesN2RQKYudwOGJWi5IfgaMpTzpFkhYA9Xrof8wvGXpkqQYUHoJC49T6E2
+LJFNF320aMrSF0nLmvG+0I4ThAsXb8Mq6WwQzARBe0l1mLe8OQxr01Y2aGU
EN/eac7+RJR0TUAE+/WuqYTXAH+5pCxjRl8MVTh2tv89uxoFqI93qy6HT75B
otJvxKbdHr8bxZw5EhENzL+5IsKS+Ay/NFLMgbLhHy7Bor8M97690BGAgLjD
GbHSNyVdxMTQOsegxOUCHE6nC1HDdQJnvajtGgJ9xRrvAAPxTQVoA5ihYbjb
AfDCWM8oQMEB+D5JLiJXalxT8MrR9dYrQtipIb3JRzGb1jIYQKgsH8JD4+ge
sqxUd9J8zy+voZMe/7QSXwyFyKOc5jiQQUQHCHYyNG4XQfEhKH9D5PrqFVD2
OlHal8VHuUDhm01tjqzjVl6adq91v8CIEKTgfsHmwQ5qsjUdo+0jyNJYssbB
j/NHaN4/3y1TqvP2aevHEqzNwabr+0h/GlX5nZG6MzSAnTWbSj5GRiQYYUoj
1HxZZeQeDe+mlx2aFGt3MKaYUMCd7kiCci9YW4ksczq4zVE54EPMt5JVZlng
GirtR8Yz8V/OWodb6D/+55FMRYOf3up7fwAVesojuN8/QlpZ01835f9/cw2T
DdIO97h01i3Lb7NsEdmlfKRX/OTB1epKKcTHTiSC3giIA4DvISy8pRfnSYdx
1NCtn+SM8uqCkit2l7uIN2hE0Xq4ULV0PKrkBOJQ1AgOaEo7P1+IuDV5ufZJ
gnAZzJDiB3xy87LwQOndNuQk/0UJvNUlI63829anv08+YA9KgzpQVA1519ri
5X565omjEstvoDffXDwvuZ5uJoceNcKMD3RMxhNVNaWKO1DnUFGGaogF6hZJ
kgvTExL4pWEtsaaXQ6TQr20PXwbgU7sUQpNbTtmOSvSXw3brNv17J34RvHZe
oT5l+KIGMisaqEx8ySM46wDI7LuHr9ie1pKkq33OpEC+3p22gcsJOSOBX2AF
Won6FcBIIc5vubB/8jMhIOyHxRDaQpphszxPe89DZJbhrk2xtORU24aH/Amj
+UgF3jLY+UjXUZdr19kICiDvoW412GsD3bSp4dqoMjjuMcgX9XppOlpNCMC9
hl+5o59SlepOcBpi7IrTqIJHBAfaOr9s6BW8TnRwWrZX18O4DC158E2fm1JH
crVcpK+T5Meu4lsOGXiQ1u0skyfd141AoeLoDjslXEvEwlM4bb43ff2HfRnk
unAfzxzSQH0Gf/k8waJhI76YWphMXNPSg2K5oQ4ZmkvATjLV/67zEpxlzCmM
+zz4OnLdDyeLud3f6f8OyxFd9hP9WIsXqR3XjXTbdS5WXOvIgoHwB9pbczSW
ovLbKxv1fIt23s44S5fpzafvUVgvi2uqUjk1YxivlL+reA0WxLT7UGPhfc3a
jBA4xudaUfKUI6NXWeH7t1I7RqXHEpmsL2Q36yDLsCh88b9/6c0xP8T4Z5MS
332rW950yxckWj5wkKgSN4QSKPLvcVJAhMrK6avpO6dObjTnDyrYowP+lGDR
uYLhCTHpuhqU04PMGiMP33tZlfi/a/kJ2b82HRjiqgLHaZV7/nmMa9T8muks
gtg8fnLlLR5IcUkl0eix10zb13fQl3JqeYI87JVy6WNDch4w4ZlBOj/UK/mD
ljyTe14Oc2W3el+PXB9VW51N+/bkkBJWMKa9UaoVGnVNxurbOphs5JVkWpf1
6Cb7Y8eVF6Cfu5wc14jYG4GCIASZpdNR09pyKlZVuyT/vW0EVJGBm2CaXnlS
GGrZUI7i8fQBOI+EaHzDO+B8NXNi4HjSnNPIgc5pdAPd2/0hXqBp5t8pnkI0
6Ur2VeEZOvjYfwv4QorIQbs895GIvmpPpjvtePoxly4alXhhTDO0FqQl+B+m
efPpHOBAWHPIDSZZfyspGybJ+aY/GKY6dAdVGJ5PFm4G6GEFYMoETwMYqcax
rH27se5tyrNAEd5NxrxhlckzyKmb9y2zDDo6QL9nTvrQhRfDxq9Zdhh6BJzO
0EJcBjZsPqjSQQQKF73lCLqtuSePqoK4eqtT8xt6xWx7tOP4wuBlGDNtdt7X
rtb9ZU6rn0J/+1jwwbA/9/lmm/WvCdYWIx8IFGO+gZH0aPVHeE4g3hxJpCTD
e8WWtACG4K2dJuICnrTzXAJikw3jbAilhJTYQn20H0jwPcQRR2To7+buk3ir
Uu9Ag89SQJC4o/ehFsoVokBiyN9JJiMjuSmkvXerN7bledNN5/111CW2p30S
eg+ufQZijoKs4lUUsHJMlhfcaLNvM17AcX4jMhXmdp5S/lu7Gr25q7OCufxr
zwJC+a4GREPDfTcyN8SCswrSSEnNiuBWwChG1FjjCjo2qlWc5nbg6pW79Qkf
hJt5fJV0ogR+oDv5kbT8CRaXE4Ob/grPuLN2ib4uXwLGKexGZXLOD+YTVTFR
XmjVmtdlWCUWnZx1aPByBW8ry3BVTMKuq/auo3MV58tvZ2uvDHcPuctCl6RR
Q2b9mS77F8QxDHLLl5NB0uty8DR6ARAmCK3ByuLPkpmPJuajR4wJPSH8KJYQ
OnbFzY8RDHW5M9X59KyJxO6lFhLMVMOAb+8GX3KUjVcp+KaG/HmqhFNcxBOi
sVm/uSxIHtSOqtsnqPFtOASyOmfzoBj4HxOViF0VoqiamkZaky/9pzrOxOGm
8VG9/9Y07HfD8fcPwlji65V/EMjFAfRIoGMBJgLxBJ9E8e8cVCJG8jXu3OsY
8HSx5DkMxWFlaHYRmXQhpVln0kPAxIn92sdHfPitvIFv2PwAvIsjGUO5zwmW
GGX6Om505caHO/1Jfxpu1osiQS+MNLnwpRssgWHlHDJTnUDCgmPxjXebl1uh
r1aTayFngZLBxKJvLIUagx3A8+e2f85tm5iWFL0eQEy1hBFTiKKpruTWqLdR
j0v3WJdamD9ctaPpTTdCn0f4g+SbFeylMTjGkxtc6+M1WoubAsAXn2bFvoPx
Fvna8NvZF8QIwHPzs0PTdqG5tEvG/f01/zIa7BPqXDdOKHiM3GSrheHTCwVq
tM6e89z4GsxkIfb2DOXW8V7d6P4k7pVgWtY+auy1cKKTHZXAZPUhhYr+GzrA
S/jA+ryWClKnIxmoyUV13AfOBHo7vs7vLEeCqLYuik8CYali82JQFlAsJtrv
GB9n9cqkFOwAa3co/H9+ktKH6vAJjO57UO9b2z9p2ZkZIsnomVCtDL4GOwPf
M+tKcW70FRVd6iNAse6tA/bDvU10RPF9qfuvKvYlVbBKEmB415X5KdTN/PyJ
4J4IhWQSjFK/bapdi7gb53Hp/3ib+easrNJd/dJ5WcXeerpkXklrNxf9MIdC
vtDjKg45za0nDYtUZfVN6bVBtDQtO2uKwy2IAmnEZ6y0LRDpNVrPhIUKxfJF
KzgKqGT8tvgJgJEpsSLWyaKz3CAeL4AbyXfPvNhvNrC9EFKjlQ3RFT1gSAYq
tTr+tYMr5TAXQeUGt2D4ZSGimR1CFU5VcpvvgAuMa7i6e0VqBw7LXwPC4Pwx
Meii+aAz+v/f5MWOqaW7QNx9TgUTSIrinsrlIb3jsig75SacE+Wi4mObLKD7
Qgz4/GB1HeT1v4ua66JQ6qCthlIz2VuDzNggnq5pRfXCq9kEsYbdAM28Ryuy
jFK1aKPap5DcuTp66GK9lyYxeJAy/uV4N1gdrX5B97b5mXylKRvSb1FifjMQ
Qxdd3uiJROSgpjzKsSaqNo6h2lHQUSDs0+e8TY4YubJwI7WKardmxV0g2nev
wRZ9K3jXgbXMXnYmqK62Xphb8wD93SAA18RAFjSUNMExmtgXazLYDdhIPP0w
5dcjNqKAVrimbOoykQUPvjYUrslx03UsSFjAFqL/F/QMudQRVAkMWoM2/PtM
VAMrhudpGVdyEK970tOEDlR0XjtrdbOCjB5qW5SYjKaWtOi6MmlodJwyqHxM
bcrCf6Czo6ZzoInfF7VLf53pnAA22xmQxK4I/8taYtOBkRfEmz8jF/baNRT9
/STZUqp3Uit5victR/vonlC/buk+iD2q6Wr7E8zosY9CCtvqbmkzaFkVTLG1
nTSjR2cvKlzA+tsEs4cUmNzvvjnxE7o0g1r1eSmp+ve+eFSYKukFzqFYzLhB
HCjoP3OYjVoHSVuv2zO+P0r507X2kHLCpF650OCvX60d8XShjE2E5993V8Oj
hCHIiFz9OQhleexoxM4v9hyeU9U8Acpn4Gh0puNpKKIojechsld/9osA7SLL
ohlHeUH0qLftfYilujDE9w8TAKFVKIHoTVVE9gjpBC2z6o5pKGOeSNKFW9ZR
1xC+ZnP9LilqgV7gmaSaPR0m0wPNe7sei7oCqQyudmND1RmkYqa/HHJZuqZy
RlK2yL+eH7evXpQT8l2lW2cnFFDy7hkws/sh6Xf3sudzmapgR2k8L2txN/+1
Y06MwTGnO54YzLw9Lj8v1Jj84DPOz5WGeV4HbdZDeb7qnITJHpk8X1vvPxDo
f6XMN5bpfGE+UDNUq2FKDQ5zTwgg+coi+XIWpVf2bxsopSQj2/rU6bfjgTu5
HpUrpQQTXAqIHK3Z3gxXfChpwFQ4rNW2J/uxBcMRvTwHbqFBoUfKEmYVvYPs
bNGvkG0oWrvxzKXMLWjmaO/izdQVfLv2ezx4+wqoVmWDo1HYsRm57MQh2AAi
sp6YvcEx37JRu4ozx+vb3qZBgqrZE89e57T/Z0Ki69D2wSRAFXlz9xxgU9Nh
RKgF8G8hXOmKqfoVscG6EnFitns37MOiUzDMcsY6/9E9ozOGV24x25AOy56V
fz+PTXRhylO+5UsdkbxN08IC2Timo5j6voAF24YPwXNeuAb2Be0C/rTOfI/x
OhLXs5nNSygWRIHLj6MWstePp5mUiaHnNcGJmzOg7kCtnjX4DY/E/srId5Bu
HIBnsE5vYCM+0A4errCFHu4hBLFlg+HSp817SuW15RruKtGaGNB6OsQJdEAE
nr4H4siND0/3krE6ACPT6ImLioHi0sohCohecjgIAfVdUprBrGRbpATtT8LT
2fIp9wbwQQzS3QzLkJX51Gu6RRQ2obm5qs3m+AMdM6HWXZiT2Z6kRnxBeW8R
ALmqoFOQb01XSugUISBNpZ+4hCsKVKL/dqpJEImVJTj4CvNISP+xqx2DT08e
DP/48X+5MDQOKMXnCnxmdeIa07zmYbE8WhdgTol0qbpjp/Qv9tMDXFdSj4zE
bYwXkeZkX6bomrTIVVwyK7KopkN4G+Mjq+jIAhRmRRVczCY3VgM93kJyrGyJ
7Qqao4NGYkW8dcupUfDMe+HauLdH1zRO+rco1JIrg6Rrh1Wr3TVJ/dOqIf1f
bfhDozlPH2imZfZmi8dSRTiyvVXU06/hGLSSpNx8r+s+4CISJHeMwQoQqhg8
S319r+ljc1xR4SHJgxKo08B9xR1Cxw0dGROi2C5uwSswOaG6Ecv2EXPEmagZ
OyKdzVg0JagFv7rpNjA1omOlGvdKA84Rj060o8wM91jJLNtqjnZkNqY1hHnq
O5lOtN+u594NMW0aLoQnrvnKY2lxX4fFdMffkUtEnBO/ev0jSPdp+L3MenBH
+O+rN3WP6JzI01EWPKIBCN+5bLqLu4BnmOvL//plvOuDdBB2Pgkckv0QyX10
AAvoOPz29ALkO7W+MsL3WAfaxNqF8OMJ1u64aDNRbllsteBXTYQv2VjJMOaM
VY6CE5jrkPeDs6fmqsKG00IOLU2ouXCouvjGsVwRiVeIpyJLZlPwPw2+haj1
JKRpr2lRSGhfY7GGdMHGAIvzX80MEkymNdAg+Ed/pSJpSM0TPv2fD+fyUD4F
9fMAkE1GFAngO0U8cFxM+2reXzw2e0tlp/VKId0OPNBFiaeRYb0qpVt9B9bO
wT6X5ooz5vmpEIYo9dmFHO4URQ+sZWfcKx2AJumNvXUY7W6DhWyvl+lXBBxI
PmgZLEGYr6oE4bPP6f+QMBu7okjSLFltucyWJmLaX3cE16IH03O9fHYCouI7
08Zk7g/t/U1nlLPaeU38bs/ypMyqsRLXPqofeYKTwWJKOlfqOIdXytjxJRPK
v7Q23OK74YGoU3pgWYGb9RAci3BXocgOoj6ii84WLekEUIBBvKbWR3Sv7Bvb
c5SbB2LHBa8vUlyGwzR7Z8LyUMO4m26K4S2Q1PsoekCU+fsjOj7X04UxxNCi
Ug6Ns0dPZZi22bhm/nP8jy1tetdpV1IRW6iEM8yA4DpOkNo4vMw4drmkEzOg
/aKacMOjFTqJ1vPV2J5pEy3jzwST5vTGcc/ejD9pKDrdDmDcIGRr/OuC2UbS
RPXfQBq/u/xnGYZ3OYKTKyMvW+z2caGNttsHCSl6elkomZLjb1Z6iSASbdj5
fQx5Vo8xIuJwh+m/KZCsyL3TYJkTwJVIatu22g/TXW/1wbIkPd8sPCxWZDrG
nji32ddR593iXLimfSb2y8u5TrRncY/uhtQz86tlFnCtL3Zf/2fVFPAdzPWg
vZlBSIUrh2if0ky0GzH3mTbTYJHgQnmf7QNmYak6RXPc1fwUXewvvUHjJ06N
oGKJ8geTRlUz9URPW1ifsDlVUWzwqlYRMBshUTyN/YN9U7sernkXnzI9J6PR
NuSC4E/wVRncHOANZ3kUISq91Sn7mkUXfEy27QaPS6993Woi1AfdgKVcmVDn
psQKRpTdwvE51ADsh+kH0+NrZe0gRtB1hQDx3RjG58GoTU7Eqg2ti3fndHOh
zcQL6b6s6Udo1QZQeyEo2WqJKH6DfWmnMo+ew2Lhdc5OPdTAab+GF8aFRCxH
PhQhRoxi9GF3ioZhCiW0q3YqkSIUhTsmOHdhAIidtNO5vcz/xWX1qveU2j+t
5GQ+zep5dj+kgoqFGWak1irTyU0c3EKLl/q0t2cWnN2w4WK74b/4ve6DOTmM
IH/jEOrXRHbKVCdmdEcPTN6cZS78EbFrX/Hoc/QMGCeOLJtZaptB4DZ4WUeU
ftyiYGgB9d5rpd7ZqkDGzY+Zv/OSSoyeOoqkf1bEnm3uT1XSalVLmLQG6fl4
SenjrIapKkDYVaP4fiTYb691IUt5sH7YTiCef8nOb1MLTlsNLSZeqRI2AVgH
MDAcc0brMgj5s5W44xirIrlrz6wFk8HUQX3o9R589DScKIZm12GKbs16xBVG
7xMO3re2B74sttaL0n6kTl8uiyWQTIKqCr5ZffMBM23SC6oqMoyXDA25i4jA
Eou296tM2CPIGESvlvQ/1+aN+zdluO7zqHZ3DC5/kaf/PNV1uakwa4m3PjfZ
zy1gOO8Ufy9G1TamN5lNqXLh7PUlLFskqgfUDZV3MMkfC26ht885ShJbgu4D
7iA8jtQ6LVI5XEYuMzUrLYHglRkDkEhTEX3RuJvdzXSt7GXSxam0DFB2XPfu
9XzJmcznOEeVnPVjsjQRyvdu86IC5tLMgGC0h4RdEp9qqRDW1oOBBRF1kvWV
jh4/jlrCpqq3QDs6pght5f7UVrqKq3dVt+2gavlGo1XloctGYkp+71/CSXHO
5r5OmPKFmjvLjCjyNur+d7GEGHnYzzpFWtKXXF5/9rlhT4nqOFZsZ5/t/5hv
f7M9S/I5JgQL3vf1C4J/9O3svf7SE5lCmUFJdBgFj39RK572aS27aQ2JAAMb
bjEw9iFnhcfG9gQGqg+95oCTI5/ur+3gZAaO4qjDQvhTkHp9PG94CcI8hNaq
v33eI1gglanDl1qR8YReHYo4SmVs6Gbw9yUm8xr9yOiWA4IKMZ9JjciYM410
lIXb8vH23riY9TN3A3Czn8fEJAroBXIWNxqHX7vUgGgwqAvHydFhUyk3e/0K
zKr0GIJR5xsgSmYNWDzjCwf0lR8ZI30kj71XOf5TAS1ZpTq2Z/KTkmge8KTe
2eKcbw7VE5pFspF5IYpgJYME2DqTJanswXC3As5LDmyNYoO+Q3bUPI1h0Bmp
BQXCK6FnEvnxhNbBdONH/0WnVEuelUp2leNe4FJ0S6dguuFHhK1uRi4LLQf4
o66xk8q4JkBvJrNbiezocH4I3u7P21LGckhvP1vBDJnPPbMxPPo1M/j1qSSZ
/B5/WYk14C/iYQk1Dt59AgCMTsJs9muaPvoNVnE/xNomXcdJdhkCjMThfhaV
FG4FXUNQlwpb6N6GwqnK/k4PzN+yo1KmgylGkelQgG2UXF7cPuf04HNyXfCV
6rTipk3nh+lHIeE3GofyfssYaXOtEvdTXDpSZYWbm/c6ylhDQBMWO/VP9FT6
133am0YtlHxHDBy5AVFcbL1TjQV68Sa0UHJpSxZ3t2zZa8UkI9pjDRzbGglU
x9FiSA1NaDB5yPCYHxUAYfBt8JpWVLg2pCml37865BcfuuV0nMChT6JWs39U
NKvu73wzKE/7tLYKQlF/PA0hri+COtbwKDex6e+v8KZ8wMk+E59mPnjSbW4+
i687sSLhLBwO583W2ExenCQ7XTtCPWS+swvDgaWDKml4sDRpTYPRetKorMgy
F6ny12Je0wiOBoPkfLUzXuAWuB6P3DVldaEKhHVyrajsdIH71mKxEnwyaO8G
ZpY9Yu+2TjcEu2zprfu3w2NwCwqDUa51jkkTi8D/8VzTa72KRTiBhnY6eI1u
laCqKxXTF13NdbPCfeKmABnJ6FV7Yo6pXI6IIhx3xacoDh9ya9NUwkiS6qcw
n1D/8cc3PapxTIliUeXBAAXjkWcXkWmtjJcvbRjU0ZAUY29NZ+701uuHte1s
jqcFiRrnnPakPtn5Zvok6jSt2A7NmCieTzugHcjYA0mINUdJWAze5f0FKG/O
43/vcRbXRsK5ZY7x+w6CdMwsvMO81rx2oj+NfGSlfYaKsyFsJ4vWImksfipl
37mu0LqxPSPGs/GFUjs6/1phismsIbgjvmDDMWNW0gbUWnDMkbc5NT5tucBB
NWmNcYSNZTGFUghAKa38jsvJVeRoxe1zmt6F9xDDMHPw/teCS3v6Jd56u6Lf
wT5yxHtxsD0Mn9OD6s2eigMBbSFftgh7g4yBnU13qWmKOhAVVvAswnwtadBt
GdufHOr80G/GALg1NVNlbQFb2QKMfw7WLECaFrThXWdA10j6fx8PQSCwSj1a
+BLWYQRdAAumYwxIreS2c0ePaPO1L+3aVJVxV4fhlIQ/q4Vn94YkvZkvFPE5
xoDZkT9BLGrzPJC7jRwmgIB6OqoeNkjAP71kf4Wnf9t3tprMvLv58S8DvyY/
1QbZ1lKR0BMIABCzXT1UYqdFJf+OZfqVLrFqw6iSGjRaen6CfI6idOfrEeoJ
f1UolwJps7FhvKHzn2PD5AqZVdp2oJ93YPUUyNh0953usDvHyzRDVDcTgN7O
TQZxGsZrak+QUGkY1NCUWS6ZCDl8oKhtuysm5Ualz8Cfh0tGZ0M2GfXSGpOZ
JD8afQKO9RCShYpzrkNbY7gbZCcK3SJDkm4wQ2SZKLmQfhFt4o3/Ur6VFRp6
By8b1NWJQEwS3VF+ftzuO8j6Gms2eL2lpvTWAknbBU9rs9gd4fLeuLCkX6Zv
kVvARsv2XhptL1P05IOmedb0i0epWVugCy5hTy28QrqXe2rbMCJpkui7jOZE
eXg16+Z9DPpez6TCjvoX6Q6TCLe5p4EvzMwhXZ1m0BFTV6HdDPIXcdMRTZYx
qEz7jzYgose2s5OosM5bNVcXCn3qC7QQSzdOAywYRWTQfpV7k3VVSNzUuA2a
T9QwvMWG9dwGxJtMNMGzLkz6MwUAkWqqYFfqkTugU7oqEk8dLb/sXb3DESCz
znh0jdMJxiYKzqB5OTVr+YaGm04DPktdoqx8SJO9vzUWJT70mTe/t46647Fe
XIkvak3tHh0i1xovZFUVtyHEZNdT9tS81TkcJU0OpkLYK74RmxAolTc3hMU+
4ypbaT4LI+U1RBNJTuie3a8midjqtt5dsx/QR9j6MiMym+aDTiNLZlwSleo1
R6vbMv4ukTc4J3LV7wzxAgxHf5mI6YMqcqg7XGDzofj6B3qrVNI1TGPeok0t
0omGmL2gSCSOTl5AgBAF8B+H0Y6dOx7nWGZqZEUv1tBJG5rLsYJ60o2f0m88
f87+E/AWXT/xszvVzsJ8cmdYDOONB96vVaWhaWO/BHmXkY2ybHBWrpetlXJe
H/4j2IZjKPjrXMBGLIoXW6yaCLhpA3UOHhE5Ek0zwdaZu7OidRYvZIeXNpRj
JxC73c86OYC6xthBUrPkoncgo7qAueUypNj4LrlrA7Q1fmBCkaNEnqEYlqbZ
CazF251nEu2QHQa8EStY5R6ntkAWM/HfOxOC3fJf4fxi2Lv4Gl5uDZ3mQL7Q
ZrESnTm2ZK8cA02Yi7sLmgKGMa2En5F1kQZbLtcoYrBH9JkVpwU7iJ+bAdji
LIwO+yGKiHi07VE30LvJ0OV874hPJIy/0HS4RWoTA/mzish36Qvenmd6JWwG
8wvRChCD5fIOudAow/NNsZBJw47u4KHQ/AxtfArPU+UEhvmzRHOGeykQwdFY
Xl6cUdS1YBBaQWbH+SlVawsjyKdzDf7/lc+5B2cdLX7uj2QI6AwEU4agTfvv
PXRYyZm2Bu4XYbdn9c9riBfoG3zQiDshpaV4n0UPhal4/sCv5XiTqH4Wa5JW
navPDCffDOk0/x6ChnzozDajbnbMVhM1EqnaedMTMTlG6LPyxBmSwT163cUW
r6Hl9JoPszIHiuTygXgiIX4E29WLVTa0x32jAqsOA56zQwEjCnvHX5JzLmQA
o2K/ml2To3HkLHPL8a+60+kBJlkJXg7gaL1S4LIli4xaRJM12MNfYW0IOZDx
0FkrrZaFkRRrlKQOCfiajOq0LnXx5XI00/iczqY5f9VjPZ88D0ybjHl1e+IT
+WIM2hEyccXU2dzqI8QNcWrd1gB8l0cfqtBfsJOg2I0PlKFAfeRzDPbIU/lJ
vs42NGWq8xJExsrVEfdGIbl3x2kjY9LfknyLlkg7W3lbV8kTacN6LrGwx47p
twlN+wW5NqqpyJPjaNCffvBptC/Zy3VOc9M6WC6Of2iGPfZmSm6LUjLV38Ym
vJjgudVDQCMUxBSYZIgnQA9qeX2WO0DXT+ocd6xwf/SH/RQY6DN9+Eu9GOUX
CHYjYHg5armUK+Zu994DZunOruht7cJEJZ4+K2938CynAZyqOLfLfGEuU/Of
eMsWZgmWV9krVISlB2UG1NikLh0GY31WNnc9IUAiFqNH4+BUQXu5e77S2KI6
qtjPlYL0Zj2e1NOxHWJBxyRUwbWC5pwKib3RSdEbrSKdCHUpYgZt/hAEn0kT
DfxeYtuLDVppjcGXK9wq9C1zUdOjY+ruqo3eh9qtAvLFEIvzrEFSFJLg8VmG
IXMhDd/ibCNyTP980CMNToMwAZDBsZFtN4ggGJd74IlpmrhNjNVBxiM7hSbd
z3P31Je1x2vWU24/CaR0q+yb/8LHczE3oGirqWw5kldBO3DOg63iDDSdcLDy
WNKeO31Jq9E8DsdtkCH8b66mBNbeok/wSHZORKdWOu1zNqUtV777p1Z/Wwxp
mE1I0/x7ZI+smANbBGaLTvpRmS1crWc4Yfsts0q+grKEIzxC27QL2DtYqm80
q00/5HPXNqUMakVbHgp7jxLUS6m9D0h3swE0goeSfkbjbdvY6KsVnmA0emaz
dayQZsM4BxqCAht/soXQjg32IL1CV0V2MWH8q5JO75C7k912+If0a8jmGkVo
SRfWqFDyOg4qKuDrFt0LRiNFoy6JwJ9xgbNdWV1oGPzJv0Fnmw8ed9dZLsTs
ODVt4IdRNlVDVvuPDI6dvPSDN5AJM0LTnXLG5elqK5Ug/Ep28AhqkM+bsDU2
otkWIBPspVLACqlECrrOVBF4EYqzEbGEVCNHTzW9e+P9g0UF2vcg+83/kgro
PsQri70fQp9JEtzQXGNnO+cX0LdL71ebR7aiz6vX/8F0dnbObFs72StzIR5A
PP7+MLLj5XxRCMAoVXxFtv/IvAKuT1Pi4gDxDl7Jvm9wvGDPDM1fGqctGQW9
MVaaVl9dZ+ZdWcz4DNBN1Qfy7RiVIJqmZn1fOcSiwnxY62NL72ihdKvqiJWM
6TNWSLYOrS95FXNAQqVtbShRyuHgp0TzqbgMK3xIog8UauJ1hubgpf9xznaA
T+bI504KQWL8uPLYZN1SXCjjLNeIsWqCLJS2ifV46GKmN8uenOPvc/w8usU+
u0VUxYZ7TNWMfKVCi+5TTzIvON09wWZb+rK2JLQTX+nGVK6Ii3hDTbYnFBQT
sgX3Mv0Q8Dfn4uvGLgYOSvZYZrQni8JG4XyByVlOAm7cUtOh3v5qNx3W3zcK
fq8wTIJPTwKmeXgY9lubgiIH9Ti6sUWc4t+AEJO7WgAqeEYbeT2WPgcg5S+Y
kgUxYlMTGPIGSOt9KaSFE/pNojqYvyiuBEMGIZe7Burj/n0NUdEXGJMJP52e
gbMMM3mgKZHCEkY1Vjs1vkwBnUvl/IrQXcc6KDWgs7/4mf0gNhE8LejVjoXc
XIuMk4d8xc1cCR+/SHUDNA6adCpOH4R13+lLHGfPXG/QF5AwHssMmWZSMWpq
JwA96O3KT9aBlHCVhUMzh+7yvuBTz3t2h1Q8Vkbidrnl2OA/mhe7WvJwXZl7
Knzu08Sdh4Aig+ifMiFVnyrn719T+ow6Z0QdX/rWNcWTtjlq/7mft4NMgn5q
38CJ39le6Hs8XzS4ZR8vkMv+s2nTogsJtX2PVwXdA13hSCt7muws9nRMc08a
p4PG2mBbc1OKgFT1DdwUKk5ni1h/S2BjY+omFyMF14fItEfJwkzB5rL/Mtb7
agnjgsQILE2DyVlLH4Ics7+8/jPC4iKVGMgClcJZtxabX/6SMJWpmoZ0mmU7
6tMjKE2aqrNI3ef6aWODYtpntqGtf3+Iqz9XyuBAGpGaUfBZ42jqfD16M2mo
VDXO9N/oFNh54/RDp9dIIJIHY/L/0nFA06tI3Di+xOEK4DBu0tg2xRgm4KH6
VHWvCXieYysKd9NT1V8hs7wKNPyTGP9pCFlOMCigsxpgcNzUVmKTQz0AAGuK
k5gNDNgIIBNUcoxDG55Go070kFo3HEnJfT6j7dkeS2WGycC1aNiBjSze1iPs
zsMbRS6bs0jRYS7iJLc0bJA8LZbHFZL0ztDpxI5fc+ju9WueB1GVw8Ainigx
S8BPNv0TyQVBSfIsPunwXaNkqXhYfdFa2DPV901/LgQwMArsse798V7+dWI3
3LqjY6+3R7jzH3QyFSG00Zpzh2bIuP691Efxp5upb4wmwDEm2knz9KvF3AC7
MagOSWDMTdBpz4kbH3Hp0X7VFTuF1Lxd5t3cyM+TMCCCKKR6xCVyJszvEcox
nrsvW8HVgtOhZ5Nz+22qm5TF2EmtKbI8FuO2/V7U6Hv1X10mKMhOh3xyOQQr
uHcsI6v4X55p90hm9A7ooApagDvjKjKNSwIkM6+yRc6fEjWwSejWQURHeLKs
GYprY+GTWtJOxZnX/JZ0YbQIw0AD79RRw/ajzwVrtYSpC1bwqz4zZQQbbkf7
umCg/4n1hqzg2KtUziW0CUlKrtpBczOottUX7HPViTDHf22oJsN43OhPgQxJ
Iu+TGZ2AGiKJ1QgTgwc9czwLnVQciAXnDZ7TQTuyNGc5pyLGL0hgjs4oY/DS
7qH4TnBhBCD3RqDWA/b9k7uEQQq05t1bx+1U+1jfLhU7jOVpbfC4rjkx1JLL
+yLxIA1wXV6/ziiYuUv/MahpvbW8bWhyPxU1WRoNlNrK+xgN+AgdvTvgr1NO
Ce1+IJLajO74kMHKqfA4FLcHeZNheg7qvDd9pXm2m261ne8SK5W2jTiFxNpw
N80jiLR3pLHlcUaLa6MPviCqEfjMNfhAlqEmBwfX7yjfKtF4ooNoC6uxGnje
KKnza/SdQZeVV7o2A3VA/8oou2A8jH3QgoWFraUdL0sEqGlihN1n8nxVjPKB
dTKcT/bjZAseAsobHPthBVY8vVAduWMNFfa2nvVllFNYW4xNgY+JkgAKR55x
BnxbNTdla/wyjVsP8q0S93msHmWlEw81TnWWoz9PCG+ApYvS4o++YIybbtrI
UTboMRAGks/u098DgdKivpaQnqxYcFA4M3YN8UyO6yuPaRTj4kM7WBg4wfXj
sSpvx2+He3Do6fl2erLo3iWnXGQECcUasfAsFeXS94eqfWLOIdqBCXnidVhK
cXJdP+BSPsootYOyCKZky39t4Args3KJFGXFdOWi5mJcoLFqdduSF4apnNG5
HnBCL8S2iiM0QVsAhR9q90iQMwAeqNE2Btu2AYD8W4cARhYrRK+m1xQYIZ+x
8MRjzItjU/2k6atQhorNE/kWpVc1//dDT2eRpA9RELgOTnn9+q//I2VhjiGz
gDa6LJdQS82C60b3CQ9AmY8fNaY3QI1QjrbneCYV/JVVZGZLtPH2+ZNoSsCX
tvs1Bk56u9jQEsk9khaauTluZlcB3B42X/6F+TP0C7V9DGj3nEKktintWFCp
EJ1XxBlJJw36HSry88UzG+TPMHZV7XvmufyO1bjXKib8cmFvinZr7Rlddp9R
l7FZ+OvALlmPFAZgtcmzn9YCtOWkDjVgFcHp+ueIJvl6RZucxAmaWh6ttVbk
Iscud7PQ8Y43mmBSPLWGoFZQqBziAALQoCEqNIIMR1XgYo7LqkpYBhUox80P
WyKUgE4uihdipSe3JyrbDnFCl8SPLcBw1oD9BxbOaJ1R/1mD7sftquWXgIZ0
QGlK3J51G7gk+lzJv0EmHPbarPg59Ros2KXcW4KdfLvwX38gwaBMXL7uJpVg
KLgB2H7uIqTIchcNSGY8p42vU22dQ1G3revVNYFsVLPcX2aYKztTrScghQ/m
cgBx0rCdqNDbN6XC2Rtfn8ROnb9modn/va3FzzAeMRh5ak7V/BiESrmRjbhA
Y3ZDtTJ5QkhHTnxSDnILF6z3vHGN6J58Sgp9TrVOywa12FXgc+TFsq6s0Lhj
nA8+uu4OqmUDzBTV/FyP+A6nIQmS6CEAYXE6SodQay14q6ejxvyHbB/JpLLZ
y7nq8Yn6GmMZPc/h59rOtjjF/gMzzePWdmgktAeKgjbPCUPBxHvb2Nmfv5L6
b7H0peUtPM0VRftXUahH0owGwVIBgtAWqww1eqSI5R05hxKzTw5+ZQ8MP0Hl
ohB6ZLG7Ir+qtudvJxWfEnvCiLJQRsR2i19F3q0BTC+8b/M1U0o2hGcuq3X7
5rryh59izaMd0KNxa5I9FCdrsWCZUHWsFUB6G3HcmKPa4UVlyKE6iW9awqSr
MomYOSPFF1oO+k8FTMEvmGYinV8j/hhNR3LTO+hP1747ZODJPdmVjg2q+xIG
FU4iRO4tGxggmJe3oZenI6E3ohMsjQ29//NZLYViKoXwFldBZtYNU9SXxYq6
JatMHwjGuxJy1N8idTO9Tlie73OsutQ11TQ8cW07wC2XQPTcWOIz6istYOHp
zcTZkT+MnWTDgSVQyyI7kKPfrSGnmh2t8gYTz95i7nTQjwF9khaIf6kODLnK
YmlZwjrkkGK1QYLf2gHiEpc8BqoTtbbX77DKE/lwnPr6C8xl+vkoenqR5zM+
ImB/keAFVhkVaFJEMi/1KHCPsWCk+KpztwmdZtipmx6bsRk196ZOVXblAqhi
+7VSF8IUTf/ZZTRvzscXP6oKkTFB7F2w4iKY1U5yREyMuCyYYZEjKDqX5tAc
QYmtYsjiwECu+GAkq9dSDqnhmpTPCYCYNNPcIRaAjP6VaGior9YwF3YqwTJa
N+cG1AGibr6YdluUm05jUu+OZPxXHnW+GPY4VIvwQSRe3tnDD9sda6MAVDJt
XtH7/TK2INuEZyMKMTn7PKMRn2zNQFzbGqU/sDj1UHALkJDxSlTINKAp2/bg
/Yalveu6OjcdW4WO2PeOfx/CFE/1mHNGbSGXQA9yTrGEayHFWt8o5T2XqFVn
q41B94yuQdG+uGaaZj1PGtMu3XFhSEjtTA1pdEV7w0PCGmwykaAIn9pd9Dh5
z9VDYzThcR2gJbeMc4gO3zujmIK72u3ELsDzJMdurX7jn05g8q5zIabwurMM
4VgeqfbAH0DeEH/OnDx7hLJBHge+Tlvt/55S8zRAvkVYtOgoeo6ZBVDTQiod
k2cNfXNs0yjM93nf4KAflB17bu0Xz2/aVnR0mlCVXlVOohOiW6Brzr+apVt8
Lu+p3eNmr7j+Qtvs+Fcej7RJ1NieBSDRsty4sdTd4R0dEqxopnWSfLxyYJRA
bn6UgNxg17Jw5pKsIgB1DWLcKk+LIfZwzWrzZs632es9kpRWfN1TXKseWt8n
yrzffMBTCAAiaKzoySDSFx6v42renh26UcAYXU6HCSaVDUjLhJBg6pJ6HzQD
nB6gBEO6pyH6aw6GMvsJgF9i7eNmzOC/HUQw61azPHV5XqUzWg/QKAHKZBBB
l25GXHlrDS0U/4z5CgTkShY+hBbWsq3z/kuYSNalQ4P3TTqvJbGQwbL/lShK
tZHMuy5HJ7MqcS6tggJ64dI36HzWMzkky6sbiSSvTHSyaJq58b9yTAWm+FlH
XJTnY85XcFw56AoefjyKivNV2XFb5tR8nvJCqS5MEo4orqt7eRREoXbAjxDy
buqg7H4J+KPC+hqhRP3ShJHMAefBCshgp6fvCZHVkWW+Xa9CdRf8E9nPfnPV
XYuweVX9YnwtIBB82cxXVA6WEd/ae+QTB7fKB7hw4yZt/H46HIORY2wqt5G0
r13rQdwlUZeTUWWmoUWyipw7whhkmZA8IuMQEmWQVGByv4WiJbgYExw+//ME
icl2fePsXqir6nxy30q78HyeYUKcoPWn/Cfwgoc9fhNrHcEmemWCRUt2Kww5
pOMv+JmuFC4ngEVv+p9Gn/P1EhQruf74LVqV0SdiFxcPoVlqLPS9dHMM8naJ
lAHYTXToBTugIUdJjUIk71bywf8/ItF09Eyie925xqyZ8mYlLzVkJ5U3zO3t
PdWt8tFQs2JugF5N6gDiuWaEliL4qXMN5J138NheUV5VAiD5hFSyuRtQBees
Mlyv3bAj+m+GJuFQxdVVrewW74vyYA07i4+p0Ban0NTUL8L2HLksJL9gdbQC
PLg4h407Gwa1mpcLaffQsK+YzmSUVZBIiwZZLLofaV3ajrGinuqiMtDqyJy3
R6JdTaeedw1oms3g+gzmU4BcquvTSgzDy+mqME6HZg69fSZwaOhrRZQKzo7R
DjM/YOBEXOd06vIwYb9msh6BFIIdzvY521hy8jpJ6hWcFfUC7WYs4iq0gBBH
KqReSiGc6hOrcywKAhD+NInGIXf1JOurxRMBtKhiwBakS158eaFyr9pfPZpa
KFSbyrpEEgw8thKZfLZ5+GfHMZxPNUUQ0d+zJkO4P1Mh6Ec2tBRCs+veRM2M
3YjO+ZHY0frRaU4GsfebKqMRTAg5mwNXrHBbZfVJiJSV+4MEQ+0SShv8Y+rN
F1mPfVwQOe+cK2pVFNIpEq0DHDA7+UhFmkC08A2ITlgHW+rOmL6s2eWv3MbF
EgjQtF96oEC116nMD5TsiKu+ooE9kx/XLty1wiHwiwMpjeA3I24FWhZVFHU5
rn0gwYTAhUBobTFvF5GLoS+JB3fu9zoy/YsSq3U3q58qCTSG+JiOrhBj3q7F
z90fWOowC/nU3uEXrYS11JxDvq9CHpCk3GSxqndRHBE1dDweH1A4z3IsAXhO
9CZzHeYzkX8fO7qeXtIQ2Vf3cULxAyKXEek4WgmcuzFvvPKbvJXcHxYtS9KA
t+hQxOZrCmt/Acy8pBcbwPI/rn6XXcIzmguwr/9TVNxx5XPcqEzs5tGw48kE
nW1RaojhQd+ZOSJIGFAQON+9quV6WDtGpTdH7mT4cO0tLMNzAyUatCvIZ0r6
vPNf5C4Txnp3ebzjlj6BejwIwKLCIe5ihyRfhUk4gq0eCHRzdzbBmFwc3tZ/
pd7eXUMDwczLnCHS4KwhlgY955cTX2U8H6uYggldf1nkvoG6talJPOnl7rhP
eZ4FVX65hXuxfIyWqd2il2GL91DQINgJHXchlzRDYy8enyZFlfHo6VLBuaBj
3VoXV7PwnZ4mqG5caAr4n90VB4oMTCSv/4l4CH3fZMT3LyHl2FBdRikV/Ur4
k4Jo+UL6yeV2eT7f+W4Ha2Atv9ZROOdSTPco5kf5uFcbxBsIovwePW03RnnT
qc49n2xj9VWHDq4J1MQfT8LcG+DYnB/O9T7YoN2IVdSABBvap0QMnziq21/T
tI95U8KTukk01ZjxEQixaWTBeXzsb5Mbahq+2m8K87iYyt3oxmMHzpOLSOj3
jNNj9Pjl2ZwitcDObfBhMvNCr3PHps1mJNwOXQc3Azldw+kozbpV+I9O3G8q
sNm9v5b+Fs+L+Nk4I8zEsjnwolL3+8+439OcLd9Nkv3iR5Dpnie8qssotSNo
IYh7gw8z3lnKgRmS/M5nz+ZZMeymOpTTSK6RX3II1SOtJjQa1r+tSIsnpUXm
BRxcgbxKKk2GOcTMQquEbldvhPhsEg3F29cRZsiuoteMFK7W3RwDoXj1CQFd
Jnt1hLxHw9wGd7GTm8eOG6yD5ky9EWosTZ1m/1HB2THAsvLM0JLkCtrL3yjs
NmxpSWvysxZUNd282s0m8l3JKeHYCJ79+jTsLbDPRTN1cmMRuCYlimBEnDI/
78I7CYzOlb7UpgYK1q75PC58k7BOeYeoSuzipFj7Rx13h0R+LuLsXJrAbGSu
2mNTU+I6fsGpud6+rqiXIFsz8j07+z5vRYWzv7kpxR97wpvHclk0f9ebcmHP
5TMqHXmsEWjdrlOcRtPQJpCwgHXCx28cVUAoDURSIt5oAYDZTbIvqzikjVPP
IDySrPnobxAE2WaMwd+zIswM9XH7W/Pyuqq+Jg2xQB7FBzs2YSZol/tjL/ZS
jOx/LJCED30NoSvMwjI+Afeeb0fWl98orxC+6nRRRoqbe4sxfV02+Kb+7g0D
Ij/AfqFFz/T0nDMPhuA09OCtQxZUA2Zln1gGlpp66rP28WfaEGn6P6xDArdQ
UmLEZMyTL7FPFtJsCtju7lJpfIC0BTOdqTNLTbeoW2woK5S9TVjTX57R5ttE
yfIkAsQ8QwopE10HV82/f/N/1OCzNfj/0J12oQ6GZM+dTKRaVUHA/LAk90Hk
re6MXBqGb5A+49oCbkynZCBZqZEWW1tnpZ0eKEVttjQk+8Of9YUcCDF5bgxI
ESQtuTDjq6M4dFOqK07O3EHCswkVumorQt2UdJbNMvlXfRIhuOb+gkkXu7Uu
OwAOyKpZj+6NpzMS9eP5pzzOzGQANGsQol7bRqWPB1CYFA7z1ZlP3x0NKOIC
G+WnXkZmPcka0QnIHc7h7uucF6cM1MvqLEXdI9EExrfeh8+x0bTCJF3nqiPR
P8AFyP8Nt6Y1Se8ls+YmV84Sm5toPl3XiviKEGtwv+I77q2szMFAILWMeVQD
Y6c2/pUkEsrEYmduYoL1zG/cw0N4u3DwkmhXD7EKuAWc3QhKjfNUrDefq2Zv
5OpwCrLAp/iREAtMTrUmO54RWT/HpGRIGzDPDcoM2ZBRNoIJSp1LR8xlTO1T
5lOV70sdIuzw1rkLtGcWZdc7C3y3OcIbPv3ksNFT0Dn07IGaXlyoci81xQvm
BEgx89DOR2sr2yHXB87h3dEeK83ZZ1PVMDGU409YEPxgHicVM3qc6W3CSloh
4j36Is70Io29N20pQS6VnXbKh/mObqc103tlMv3TbWPjzjaY5DKAaNkiiEOT
LZfvdewIw8uhK2Sy4avjy/9AUy6/xFjjlAcxZKIxxqFzz9tg/+5EhL6s6rS9
/bP5aJNW1rkd4EPjIcGjzjrigDCrz+yXcn9wuLG/o0rC/GRkq0pV/SMoK0F8
gr/bNiEvjDhIX9MpILIiKy9YjQ4p008vSDri/MnSsB+R8mISkcfjKSx2dT5a
st3LPrml2qWPWeb6DPfhNe7YqMT7lAWswP/vzFy9k9+zlNGwEri49m9ovFwI
7naIO/MCRqSA/oJT9jPv4SkLZIwTIrsQbrytkoA1g+tV6zTeT6alEKgGzomi
p2/SFnbpZsRVdP24Gl47fbC1p5/nri7HrcfkbTOBbUXRlWOk98mr9X6JRU0/
HztuIyCZzAcRJi3/L8Lzds2/iPTm5WB2oXOHhN/0Tn4nast2aQl+e28YNst7
zqJ12EkmzGE0ITot+HnPjtVVWw+8NdCiSqHP7Xa1s5GuecvSRqyk+nVRG64o
vBHNhm+yqFQhxn4gXnLkwkCLH6DZi5sFu4lVg+4qghaPsWYUxXfiQb5NuZHS
v6CPn61b3MPcqB8KImXpdmPgpqYjCxTGQBkh4bXRD10qtp/z3NyCQFvM504c
SQKEiTSXu91M/xmlXzJo+SJInSApmAhwMjc6bCJHR8rW3wOqTNOknrvatraG
vpCBA3b9sEpxJ9zsl3fVBUNocQOrUGf9uLHOR1x5V9BD5pGYfd2aZ3AGe0oH
OqVt0q3KkQLne7p1PmYG6oiS+/RfmYc0LAcddqLd/kgev4iegeRBgf3QZula
RkHh0/z9liSYJ1piY/dellyd1d/A9NMQ6Bm1tV0dPrk5kLlZT6LK+Onj2qu3
suahlm5nCfAYZOkQOputLqoiUWYkq330JzOjdGRrZkJ7IbV6QMRAMjigFt9E
/yAkbdtDX9q1YMoi4hz30avAuYgtq4+yx0BenG1NytGHKYV2QBphK6KrUx5N
kH9uu+sf47dx4pTvGq/i/+RQkYjU70Mfur7sMCTsgShOK1uOS3lBWRtyODHC
nUgKR1ssexqjaL1iESBUoCgxHgScHgOJ1B3QfSts64ho7a0c/HK5hiXT19Ql
W+nYGbmb+GyLG+9/Caod1dZ2xsO/h7kSiYV/RXi6rsivdNn+nGn1ftPDEnSr
15w6dKsAaGvY0q07OXXPcFQA4OFXfQUJ+vZe4fFl8yDTf05fZDQihDNT5h6P
/F182PUmmnq1TZsXshAaRrraa/0rxTQP3sgULXpOQYhvzjNO2WOJBZF0HVEM
eAeGRCwx+NIFdhDy7gG9d6EnSPtVPFuvpfooaZTPT1kkG1qfTaU5LWzmIBAh
C2mXvThqYqp+s833O6vBXUACXwvBlIBnmz5v1+91meJoeavP9SH2LbHBWhCw
3hAvK6tuNdfitSRG+2mjWy1He5H96ee8vSe1WCkvY1n20I91O/tqbds1ECZW
tu1sGqp5Ks67uqx6kndt0dCE/8yYvZmt8N8qowtfWcLhUtta0xPQxIF96KUw
wBYyA+k/KZhLw2xZpjMhwTDhSXMN/M5x3RgILm3Q2qRnANFrlnO44EZ+gLN9
oWpRLgtTOhLY+j2aJeJk7TZ8omOXMUQ96xP43XHA5Qc22C21F0wIY6/CtlkD
TMGxLFybaRfYtAPbzwzEJpcz40FtABOcBtBr9M9dYNsBFe5pHtseBI5//Xd6
A6Sq+Eo+gap4jSZluxYBbgyqYOfTkE5MMk8KGnMvE9xGtIegMo+2ZqL76Bsc
6mzfpHI0RPXEdu6ccjve69wYxNj0fNeiSGUJ+uyTTyxkGTifSAPtRPRloNyR
v8SsgN968Qvw2UyvItomQ7gy7RkaZ0dEfgfXzN7ijL4F3nbN33UJzilmrD2R
R1W1RLIwbF7S22wLdstq6dS8mevUrFkvxjQMmn3x5ayZG2W+l49xDQy/My5j
F3J1YN9nFrxsMGh5SUxs0pW5bw8AB5/Zq5keIElAKyjLxh8jRHgsFL1AretB
O5v8UzaAvmmHWgmp7MKQfO6C/ZEPKZqxvhgRKNK4Zwun1s6p8iTgbgGs19vS
rrQuGDi46q84zqeAK4A93vgK655O9llxQ99+5RbJFzQpdG9A5TfeyU8dIZNN
jsspG14tVJwgUaYbTUtsQuxuuECTQy284J3v+TLm5GvKqYOan2DsEgodrtJ/
1ODH+ZCDesDlHB1xQSJq3ZuC+xlwX0w0lpuNo7S3wY3l/vo7M7/x6074I42u
yJ4/ZW4MgLuaQ/W22kXZojIabRIgk9kvozsc/Nb3GO9R5EjwcSIs+QUseD5v
lrd6UvyfLi7BGu9pfCQRUdxaa58rBuCtwSY3U/fWVxQtwEapJclKKEMZ9Wet
WJJpuk6KNaGDc86sBWZFY64n5pmI2cD7BtZJz2PhtGasBtg2/JwpyBFJNc0m
nPNOTdXwv2W6ytcmTzDZyQH2/ioKm4isol29C5PIGrf78/HJ2M7DxOP/p2zG
YU8b+DcNBZX6ZM9mH81kSiH4c2Izs68brPKATnlapE1FTprUZxlFjxInZhtC
wS5kcX0vNG3nFHxI5mzO5g3xWuEL4QU8a54Ipac3P3FtWWYoIFQ2yDwxFd34
8cWNDxfOt/nmHocXq9fHA+ekPEbPFqZQlY0aka+VrF1lL1KLFkMz//DLie5j
PmJ/LyGjWSBG6H9nEneZCik5VpwR8zhVmS/NPGsm2sLOxQ7jomsn0t+Y/n8j
6i0cfuDl1K/jcrPKv55mcIKPMF1X7bemhH6JIDMfIfrBrbwPjumcbI5AJtQN
QO9/l+/0qEpkiobvEDxzt7zwRrxX+CBtNwixlVCIkYnx0bPFWCMd0XokspBh
qf6dJN+g2J92lNplRdpYDbGkI3TL2q5OsBrqL6vcl/HCx6Ze/QpBf8C3Oh6E
c8Omf3C1AkjM1kdeTxfBd8TfTFcxld36xrdkpjSiPkYNFSkgYmfonJgl1LRS
TemyqfM+Ug2WvBsx/N+rCfEIfvbgJZ/Rb0OEVOWxBh5UJrMQH3b2VQyn7RR7
34ChRp0uaqWE39G/0w6gUfQy2UUBIfuAmSV9LtbJSjEw8FGp8BSgCgNV34ZG
MMFnKVFvHJh+k/Df1R8UOtedMmYjxGfZpkEfqSjsE1QuWzgfGi3KE+x+0Cy5
uHBjp42JHHuAtN4DI+PVN3hYMVPHux0lzguBOF7J5IfdvaxDvG+Eoacp1NCJ
/sw7BKB4N515uJt5Rjyz6mcswHWjHn145aHkj4UbylZTmcnAO7XPP+FUl12H
7iOnXGw3Mrzbu+t4zXFO0u1EOL0YDdjBgX9NE1Mj2azn90FB3mVe2RQ+3NcS
XkwQzABB0AX2m/LQll5QQLXg34Un13V42jkJsktfqw31c5ANBenWcvWz6FjC
SeN5oz3sFylFSNc/NbYbcGoYkRhzCL9U4Z5yuRD4uYcyJ9S3OAVvB260Mwf4
VwlxCdJTL1beMa+GvqBHXcMpjA6TRAkJs9YKofUmCSdre3poU7VpXkHNkmAc
WGODjqIlc2Ng1QcXAUK95OxEVTxbGJ/Lrgm7XdDDCaBbKWM/MVe+On6tA5cu
Ef/WxgY1bCfsW3uIVjbEXVJTXRmlSE87gdBM9L+w6+HSQIOq6kbe8dKvFROs
maMfwwQWHTMatraKw/LzkljPaD2GshmycqKmgQuJZeVozV0mXggL21NSNHHY
ExAufb3NJeXuez1jBWD6ObCnk6CrOu79HSAndTtYshKt5QMbvayc56HEwe4p
lmk+AEyUP3ZghVNZmvdoBSGR4bgVsBlvom7ri03MZRhA60mXc97VnFMEC9jR
pZbfeJ6qs6mrsLJN6Bj2mCLR9cyiAscm+gUSvjltwoxZ3lLLE1RWELbLL8oK
s3uC+UZXB9oEFNxqVPAcnc6ukD388HummUquFvb5O5+Wvd1/PCfkGB7cyp/m
AXE2N+Cl/z3KwWo4EGgfo/Qy0SLbIEeUeUoM9L68oL+Ag1RYqgXOri9qtAnA
U6olEjVpS72glNXGywlqGZl83aY08dbAG3kL/jsWJg8KU3kH+7Fj5FsvyA+f
pXpxfaR8j5lmelBt/jkByxIhoM6AivCsv72UkfP839UvcFRKyCLVwEGdm88J
AG5PoXBLS8gXmGJgYgPwALOjDgzbS/KxwkVmap5rUnxRaO5ArGtsie6bCh9o
on3mTBgtPzbpalGhQ5Gclb47t/UPHkCplCtIo86OaqVlr9Xyt5agUd4rHdHA
EWLDWZctJMA5yL0dkSahB//ccAiCVQjFQVPbFsZFrzbspVh9Jc2b0F/MK0GS
p6ulK/VWwM7uOCMUeZuE6l5jHVX5evKC0FOnO96IlHZylLR46ljDBknXdFpj
f052KxY6eophXKaX2itDMsXdO65Q4DlmPAN0T4kob07TlyWLhLWFrN3F3MSq
TV4T4oGkB2J/tC/MDEZGNoWnRSDSHQCVReu1tCGSf6dYU0ZcPfMN+trXgeXV
TqObdZO7u11F7zMZuqhekV0kMy5tRim+m6c/dDaARv8uM94G2O1kx4WpFwem
5hl5CQBaR06JsmvT2AfhM90hxXUi5HC2HOjqClUWyL4iax9GdpWd9z8wQ/Q/
zcOVSLUhepLuKgUdId4V0AZf0L7xyXrea5uP7dgOKW78ogZQvfFdUpATjoGk
RB7cxOSt/pfShx7vuyhvFKKEC8j/VGXc8M7iLMxVjfDE8mORvcvmiKHC0k91
cpaePLxDlaWbfgMPd153ultpZcVvWRdfjhgeF+oNRfOu74ILkXMI970/o/eq
LCNxrxgmR5f9p+LS0qFFzFdZpk3f4Z0cjbmTevOAlL9oT6pQjqEnHAkxEz3X
GBOQPFFGYl/uILEC9tZYfGoeP6XvKxOdXx1APwxnvQ2nqOKh6OlUrTU/r3MZ
1r+NQNgPIZIjqTx/LssbREHzMnRtB4YJDhl5jWdGIh8QlcFdcOmekxMrAf8M
w0pfSAWCTqemiRfTJLc6ctS693yt75I6ygI0zca5Y89OwuNLqqP76IY1jvkA
HyYn3jlFkTPPXoEiZk//t53OJ4KRgKyXihVfCOBSCcD7psQ2eKCEh2Q972Lx
7uaVHV0xwAMZQ2tJHllt/L3uWKxhvQ+kcvEim3hGAU2ytm5wFD0WK7z4rsrc
0Ij/u64UkFcMKKA1a9JzExBHsZgr7abj2GWW4ty3uplh5CZp2N6VyG3IX20A
FczsUorbxwP4aIfycxD+uWO0RdhHjbSFO4/2HkA6EZhA2Vt1vx5S0dGKxr97
cOmJJcBC3XowHTUTzZ/APQHSKWzeY/7ex6mz3jfFp/1Q6sdm3MTCfNcH4jdX
06FG9LAw1JVg3LDXuf76CSPKPRxQ2bzELNzYdS2LYlViUxdNkNTeVoXnGS+5
dQFAWRKevPQKrE6dYOn6pwNXQa57hSdJ0JaPkVpzV7/qGGPDWwB4Ua+MnKzo
1iNtkPD210YYm4NfKpUSGfm2bdyOFopBrwvworHiPUwfcfasoz4EMgM+ssd9
EwkV3zSwzh/BLeo8iMXdUZskocITAAiFE+SDklhXRFYe1OBvfD0xUKrzTEn/
wtigLVbdpP7M3umpKGnP8CitxkkHqBVCxlcWd4Za9S3Sm8kL5aqArzNeiHLw
64cgncDRLCA47tk1q29qZ1cuwZ08ZevsayHZ7O7Ex/vrBuZYtiKpY/FEYVP7
2q4akabmxoUVy+v9OJ1E8kmxb6+AOMhldGdukFUkLpw/3y3ayT5liryAb1bX
zvijiFtPFDtr54nQu3qhSvY3PBC2S5gGXtlmdpHqlnDN43AE4OOz/QE/sVST
fdLUfINK2xxbCJ5l5r2YpINKHxhOPZrkCrEv/jQwfHf5ZroHff4QQM7fvDCr
mi3ENE8EdhZzsVSY7+e47mnlvjvP8J4PxCWUi39G0nzkPn1n4eg/h9M+THuz
xivxIgX98btZuW8aj5hcTXoFC/TmnCxohbsHV0nUsex40MzYK36kW9xmKZR9
Wu/K19b0Wru6dl+dRsguS17NDnoXPGatCLnfd3ay0m+ApZRLViMCzado5890
TRrmkKYqjqHuRqS1U35+OFiM3qcs2R2go/kkcGJ3z4c5eB7pVpZfFprXnlN7
/rFqsN7EXbOkpVxra70VjNT4WEVJo3d36TBDpBP3VvNuIKHQkiJGlzK2moSj
bNmDQc9geRZkFptSp75eLvSG09ZyvxQceA+QQqjdJfxEg3D9+DKSvqV/hlMO
9r5HjzT9igVwJAKMKWil3Gn3bViphLMookVr+dyUF9385tpaugporwYD+dHv
wZbum0qW5Z2ADqdzZz9ykG8PjVNDoBgxD5Tkol6+ejPzbkQheOfrl9kxFaKu
iosUebP3KlWD18E1vcE/yFbGSPrfBLT3VO2ko1uL6Lz9L2Mhmfkda21+05cr
Gt7Kyl0Q9WH2JTo92g0+1du80XD87Nf1k89fuG7kqS6ScXlwfeaBRur9pr7X
eU4Pd8Sy7OLJV0gy0JpL5GGNlJ09R0z3yjVXkHCRsbRrxdGfN/mKTV0FWZ0S
oZsksh0pAEBkIB6Klu8+0/G3fJgHMKkaquahwvnfi6mzr05mX51JjXO15hAv
VJRx5e+20/C+EgC2H7jWoaT39bSyMKGRI8ft+4TNubtOGH+s8CVTSkbdFV2z
lDhr8uMBnsUktd5n+NvGEW1QQ2jyMHqE08T4DzNKePzsdW1pww5tDBShw/y7
T0o/ZKMEgnqA8TCDbTlvydgVdpuw55SF49xdaqCgK8x7QumSjFQI4hXDoHHw
fnDIwpYJhr2Xiz4x+BdycyTWBKratZBnoloPo8upemNHusFoA/Vx06tluAwE
sXfvRHURVPZeMwTw4JIfGjGeIBaxw1XqwsmeAI61xMBOt96xSF5l0yN8mxuB
ANW7BLnpNyWFMbCD7RTsh6LGvD768l0nyvp74T/0blt6Kkw3XXuThOryLRwQ
J/zszTrX7/8Cpo8coAEnpk+9XLjmvgQEKjDZO1jB063NBHjc+0HuELWJvvm0
/ilkw+0c3KACTKS2TUoCC0UcBBkHarYh/j5iI9kLOPrKSC+CKC7jNOTza/WS
p07t3K9BOIsYej79EJLbpn+SW4jwZOBAvyCsEo9k1O0zzuUwM0DXq2VGsGO2
EY4disat5gbc6GcL6v+4a/DEh+G2AQh+RcCQT7HPVs/FdTeJhGgWTrExzDXi
4274lizb5VaIwdB5XwKvwCPcWVtDGZJZEd7R4Qa1nRgjSMMTshrhXoONZsyM
bPopGdXDkyNTDrPxWwL1zZabyGKlc4hxrHSjNio7a65n3r7c7vHiQtGYTGEk
SW/CgeOH/a7p98e4QMBVmIj8uKN84kZVTlIPYKzTeGtnzWK8p0N3xny4IKM9
bPvIfoHHeqXUapx14sSiBjEA3Jgv9IxwD99Y6flIX1RLNTfLcFhT9e3LBfDR
DoThyBEN/fivsY5r0q6R0yI641knGkE77H69vuEc9GfN4fdf2/7LKuTemwad
IDDgPyv9G/nkK6qYwriIWw8UNs7wu1p4RM8+bWTNLQHsYoCTp94mt3dnGCVU
juV+KIbYShJmt+RMQRUu2+MdDM8ph9mW2OOqxmwwwrlTyoqDtEYfOds9rpbm
pSmVNnYGkljdVsdrbWrH3dDHUpROvWS33K2alywzs6K4xUSa4X26PAP4HGnb
/qz59YAHhbjeTkE0INfTj7mjV5ZJG/yMJS8tNihTBAmQuEYDSfwLC4sgFY9y
PvznLgdU0sX8/fnRf+obIOVwkqTuiTH7f1W2jq3LjEMMZ0MSFWLV7V9fT5Lp
CYq8AkJDAuBlsQ2BBveIQTriMdTRmEmMXnr+vhjD8sxgB/Sg0wt/IfVxCYqZ
OxFlTweVm62wDYXZLrngnw+6qyo7BXWxl6b/hHG5190pNN4GhHnIuiuyj9AW
xOO7QybjX4CFL9Xl/W9U7BCbSQQYYX6P2Xxjrpn378GW9GM7EsCiyRPmnd9o
yN5LzTpyUosbfJsU/9bHcDuNqdeR0hYof6qYlIyGO9uABSbu4jayKWZ0ZWjJ
0J/zYtswogbm1FfofHBaN6ybP6qvUSyrXDPKGFiOwdmHLOITxh/qDCS9Jf/J
TwPKK4qfIXlalgN4JtkQmTaDw0yygcSF/lCLuLow1iFlF9llqm4r/a2vvOQQ
S9iIvhc5CScgxgzmMQ5y7AyYwm3nZKoCuGIx3Mc34MlRDRtAiubGh8e6I9qC
NH03eojykcmW29BKOYIWjCVx4Nrp6YTHs67qtcpwZDlH1sJ2WpxlBnVwImqq
rK4qIqmh4uQBdbX+6dNK6LvRyfmePc+kznTeIPcxEmRqNqr7Ud75AvLmeGtW
KDVkl7Jnl58FsfQwhI30EzuzMflLniJVi675Ps+WiqqZdCoOzGaAdgvIbFwY
v/8vfj0va8Viel87q3wL8XmD3ZVGskJfa2PUne83gbj+S5CKw2O8LYviTA7b
9eH+R99lzt32x4yZ/IsULt9bhvL8ILyW2eTE8B7XfQd8hSb+V3N1GIY/cCUO
V1TRTid6dRq5N6rBZCAN9or0X6w81Amr+eUU/n9eujLiJCOTIMgLB+L3OLNr
bfeCnl60CL2Hp5JNdqW+bW+h3e4cxzyB6ldK9IUC1qbvg/BWUDQ5zeMBThJu
j2MCfhZW8qukqOEd0eLp+S+ch2IjRWLIwIbQnPXEIBj3xnIVl3cuMEC6KofS
tHp/xcuPdE+0qRh90JKYxbc2xAdLoRTISTbXH7ltN7wHjfEcH/NzDqtWZu8Z
RIkxngZZYcx/eX9pNjFBa+vCeNe3Jkj5s5XYEe2/Y73NQqrmtJGcaBItOvd5
8YN0yIL7mki245005JDIloChZAeoBioFvAVgn/h0GkGT+lSLC6CMrnWn0EQC
xqeqqDEbLaFvirbz8Z+OxtDPgKUVrHFXAnkjZ1aKNJ4DJXH9b52UhpWqOqds
4mnUpieFynyaa/v68W0+/0B75/VgDUet8jnjPLOIyUaY270gnHmG8lECWgd4
/P2MCApDijGkWk+fcEHIWq258ycFKJsq2SmKTl124iEkiQNqBsr6Q3uVNOan
RqAz2rVdi9kxyFLHDdXp7eB1Wy2iA6X186Vq9p5J6vp/hEsNt99mkTQJjOy/
utUR7mRKqYKn+z0kx7CIG2UjCzTBVtiUQv8tpeNEud5IyhwU2YRmnVAHmxkr
pooYNYCgNkI8B/W5VlwofxZze1xNexvcIhdIjV5FBXisN6RcB+Y00enqre9a
J+KtpJXDZVHsaVWJM6V5eetNP+zauiByU0iMYA1S6DewB8as4s9YhMWH6dU9
JzAV1cM0M4GIcxUXF+JdmrMkBLiXlSOSPO+JW5F1VOtpeZQFABrf7BNFvmxm
Ae5v73UcDhm2Hbl7dJ1yxiRpux6BfWwB/Xv5N6QXNvYeFX3Ff+9SWk984n64
Mz7CXF/smvBhL8WYeP0n0G1t1COwA/3iUNKRCPkoMMZbxJ2Z6TOXKE8yKKqW
yt3Wx7T2l4NWRvsZI48LroyU+iAFh9RtBACgTigx3ivEP08SDyxUuOeyqBPt
rrKXmbIDxzsAA2CKYb2MpbjYuOn3mHQ2QFMipLoAyc4ND4fmjP91/T2jpj1K
5h1E31XXg8OBiAAAAQZ43taUqTS/LdZpEhxnVjM8L0WNN37O0iJWAxhbBzfD
QyTa4z6E36PEQrqjmLqTZNca8AcIpJJxFa+ZQOY19nXLHBt4LEFV3Er+yagf
9Tk/kaJP/OhNd+izUXHzgGR9uop5Z3JiMUQfqjmUtU7KyR4obukv8ZHIpWZ9
VmP79c/6foBjh7zK5wrytEMLyGL3kgiI8pKbw1QZh9RFaVMI6zm/b1ImO0hr
M5hU2+dCDbbx3kjqHuvzPPGsawmxeYOmGRaGA9G/5pL77GJSeTp1/b1FG1CY
PJuQqv6slUcz3Lj+odYpcmUEIfoPbEOYncexqH2dA0bnDiwM+TeVWgM3kYZW
BfShaHRwub7sFq1jHcva6wTYnsYn+ViaQIGySO3R7glywk+TST0frnhq8pc0
n+F2pJANmpAwH3KdLPqa91aHURtkVHyIUqLBXcX1lKDgGwZ3TwYGdd6R1oDO
HXBjt0zcTFEZXClMa/m/Goxsw/AiZ5TRmAkkSVMAH5GSvE639FaSIewxJhlM
3BSCpN+9TCkG1JVsdBAPcsRa55YK2RTHX9wZI0jS75pSuKgfnV93KbfSuZAT
R7uS2aAbLICPCDWi5C7xSJo7cUjY0mhbLFdaZROs7U/D5pHZNRYoVNacLmR3
cZAJRgJNu8XpB5U5P4BAQZFWWoEAChHv0CvwoxaGbOQq5jxPWsAypy9wT7FD
tv7kh/qeHXekGJEUk9gqhb5CeglRRM/YCaGMdUF8DJMsOUbwMj6+5EJSWJ+R
PAVKq9nyFS4AkQrGDuJ6GUbVthudbFDceK6tQW4k5w9tQuPASqDzPmd7Mcsc
dOCQeG/D7ANimoQVViK2+9ZstEI9T76mnTzQI6kpZObOd397T9lGF9l1+5+F
6uO5vfGSjrlP+RI3Fo6E0yAFlHmyyQQab36+nbqJEe0Sy7sSabTUVOn2RDCj
j45azZrwRAhK/9Ff2SYBG6k9zVSKLVsRMws/QRvzUW9twdfpyJM5d18Vf8e2
dcwgEDOCBZh8ICeKw8bzWgfoMPaEfbnWqHXqwtE7ylmwDJUY+W2eh0T8IAkS
NwpPD1H3MJvN6gGJ2tjfzJnnoTOhM+eKg0LXujPtSrdqac4IQAFMuJQ1LDaS
MUvxAe3OuZ0yA58PgbREhdeWiPEmkx34MEmecx/4B5EJ4h9Rl8S31z06I+RA
3FwTGxdta/4FUdhGELD7EBxzMni3GGn7XeEiGEbcFqTfrhimue23SeblcyBo
MflTIODxd4vLe9Y1OmDzlPgNj0od4INkKhIz8m60gVLUDs2BWJVIEH0dpSq+
UE6liFEN195JzhbLYcz7OCszj7l3EySgAuLcFHIb/sb4huVR12tB1smiH/El
LjGBgaHa3bYWh4xTIAdJ6y4hc+VzpeK8V2B+S32R92UWrawo3ZKKB/3hfQAP
y1K7C5b1W+wtwYA+bBAAed8TAenjlQp8Nb6+NaPCIHv5w/zpZVy+q2/bvEQ5
juv3wdjZEJOnkhBXyGNlMo8zvErjhRP4TUW8PiSPwZxhiyucSTnqUsIStlxe
CThUW14RfAvEsPQj6VVGfTg4iC1KdV1OhRy978Wd50+cVzCHmZdDcm7pcRqZ
Nen5XpRdCXa6A8qWWyzuwaaVobX0EHWE9aeWbAx6QWkLNZsH5m9PgxzkW8X7
Gn+0u0Kln8HeYVzJFQ/GH6lf4cv/yeAVkDjwZ0WuDwA8Ngp45sEjFQOzgm1s
YQs6+jkLy/aeobjUIsAx+3zrTxsBCY2TSqP/VchgQ9zdmvdlnqWHtq8a3+Rr
r26/RYULlpLExoOlx6sKDkPhbR6bTFvINEusxd0rKByb3yMek87VceD2IvNH
4ahskovs3s6lU9nai4YH0Lwhil+iSYmU4j/yEcclR2dDrozWr51I9v4GLB4N
zA5QmDCxAoIrzZYx5YogWM8dGDkX+5G0zFu6iznbhUjuTJfRLWdtxEzhtVUg
O7pGQLNcPz0hcrr5qqL6kUk91fyzNneB2UVi1wMJwgziNzxgsDpcex9qfw8l
2IoLt59mBw/G+wJd2GF0RV8xVGey/JZXau4dYYVrrv20eEdUKQyEDguWiqxB
mpM+hjMZFMZx+A6hw2wRZ+dsu6LDnOLIVg9zIyiywwRWwcFT7BgdlJnw4zmv
BMkJ9ehks4HD9vwC3nTbttJUSe1znYMlV9mJ9HlZWVO8OjFivL6c2pFvTqQt
19PP59JRqfTowT/dQznqXK5PWKAPehpgECfLA/SO+4MPVCtrQL5UYNpooXTM
DrEyscKEBmIJjoNMB8xrNdsT1IMy2F8JN6uv8OtSOvr6Go9f3nBEyuID13eV
Y78G2fSI+z7gVg+l+Qk7aKfAaoOxNQev/wxZLK/KXboKJpyqQ1D73jvJcgj1
/nNNA94ek4AnT9+U4foi52ElkTtMnai4gE4rMTHFhQ9jfQktp70FAmjebR/8
C/2qGVwlYDXcjJ7Splh2DaJjC6c2RGte8NhN6Ej8QlsH8wVER2XPxsWQmdlC
IpkIoecWSk1vymeqGIKtCmwg7EVfe/2f0LWasa+wVSb4cpU79F1Ug9/UYK1N
5GxdiKi0clqV9l0W9b7uH4BEX5m+CfpMkqMBpSEKQf+d41CwsMep2+5FgpHu
lg7spKb3KHo3Mnp7mJN+ZK6H1HOYdjd+IMisEqvL+nyfpBeoFfTja2c6Ci67
oH6nSHQWV/Y/EiOHa5IBejCCLrAk8TTNCkLHUd/H4S9PLunUkR7My4kuEdD7
VCoKVYbSH00noR7HF9yYvWWbvNJncBEbPdAT7oSpJ5+/0SJaN85zVaaU0LRR
hW7GJ17VR9UNIjv5vI8s3uYjqloFDFmIfUVgxwCbh0ZsGkugLTD/Uz85Y3Y6
fpj4Fy6e1iI6LNMEgR6jAyi2WtGRP5SeXeCASOYtJ20CaDDtZtMSAU/CfO09
7BIW53v6rcEwDjKjw/xbYWRqksNSAYUeu7kw7iwvaf1qhaBH11flaGL4ganO
odfwxFppKPkoyz9Y/4pJyAySv0WdFwdty7/y3TcarlPTkgy/K+/+iv61Zi5V
tsZ5GXq8FA0MnqQIUwJBS3LAdJdIMFI+9AvC4QANmWamDssiump4qnY6pHu4
B+qHfreF5Ff0r8XFR6AsHXUuzzAhymIts4pJPhbKZoCPOVtlAs/k8RK2i8BV
GMqYpdzUM6ZAyZuPmYAVtvbGHl8x7xUQ6jc8ybkIiOdo62S8wfqJOdNcxCJC
NITaMIzu8wU+GY8pBXUDZ9++dV4lFkD3U22XhWfKvJjtKNTl73vOjqfAp0oP
9h8WMhm1eITW8kBSQ7ciNc7xcmnHUx2dxBgKuyW2Y8lkNe/q+iMpXYp3mc1/
fblYrb4TkzS2aOFgbhE/IpO1+lLcjngwvL/Wwx4ajzSCqfC+yQjh7/AGlNQu
3EkbgWyWpW2/y2M2d380/ozLAN3xrLSuai/cScSwY2ZpdFgQQ2XD4WWUfHmh
QnaSbsePJcRgFOkEBQ6HoF3g90MzzsVHqiMlcifjqt44ljxAzyulurGojPkV
gi8onK+KTzV5piHsG16kLH2Qt0WoQzFGw1wGz4PlylaYd+nlmPU8fa0A+lJR
stDkb55bbTelkZ55nn7PXpW9MlMa5hxRXleFk93rhjWs7/4/ej2Qj49yyGL1
E6W1fr2cAGVFBxSwLciPXY5B8OK9ac6Nouizx96qUUBIWGlvFyN8MXj4Gvy+
R3alBL3ftJDvWVZYT1BrqUII5+9SOQA7tTDd8ck96V7BmZ/WYwgfqvUCBEmd
X0NXC7Av84LjnIz4CvY1x+99ewv1f1HLXsqSmtiNio6IXei7/LrdiRtOBO5o
opXdF7dEF/ygt4vcvBlmqpeeyT7JfQ6CY8gfiP+akCoGcYNo53hnhY3Iyw/P
myFN346Znj3DjPacOd8v8U13UB5oHy5hDDFPV5O/J5lgEcrPfem42B8sphoA
Jl9e7/ZBm8HRzgDubjpNsOhrFrOtoSkmY2qBLUClrTehTlwSnNwnnIWmVJoi
SrHGYbYLqwNk7gYwy6CbwneQYiJG2NEtlywsoeLScNDMPDbY8lW6rmzF7Q/R
mvgVrVi+LoCkwBm5ZDyPQKgd0/i16r1EyQSqtbUdi/LbeBMrZzDZvBpkzOFy
9K7ck2eO7v99DGr3eQj/NboEhNIIjc2xtaxjFHXzRLKm2Znp0+9TyYtSkW11
zRY4JYJtgF5ZOMmObyFBxSq2EjxiMCMrZ11LCOGe4ZoCa0ionBN7uWAe813t
lEf/WGGhh09TrKX4kL6GbNqhAJX9VhUyE7y8PcX2i83BfAS8YvTrOJlAu+HP
MgqNsAw4m7Y/bnN1SUEbk4gHIJTrrtev2aD+V2iZnfzKeRo57gE9iyBm0Ur5
tC+V+gL+bbMQrwvEEhX4bGEM6aNtsj53RmhKlbxAWn96QbydWwBFt80pAL4f
LSMta26z9hkZT2kJ9B9tRabHPlAMqsEJkde8+sQpEGZnSS9w5eM9WExiQjDS
+4A1hsPMnpVKsUVpCnXDspERLx1YTybC6aD99g5fXKsC79pWnuNPJFoylOnw
NA7CYquRKR6ji++UMVuEmfT7DZE54ma4hzxEPFpSIR1xBkmxe27mDmo7PASp
LWDn612mUJ+qQBtwh3wYDbXLaqctwTFLeA871qV3mSuupiNqJ53daNhGU3QB
lqO9tjLiystSBeVqNC9zbur6DLm3/kNMayu5axcmSX7HqMhXty10zT05YHd8
BDVUPDaDomZGlJJwODaEVF9L2b+3DKWjK+UKPORkhvVVDvWoqA9QZ2wQI7rb
9VIMUNqwUHQDnwxMHDFPaMs6AiqKSGKwFHp0aNkpfjq3XT2G+oj7+qAXPOhM
iaZHN8KZVSMntzDGuXMwK/fxLSC28b89ih8JVM3Ig6ysC3qi61l+oS5lsuum
VKGiMBPcSb1ADSYuBpCwinbvawIxBxqsRWrHAQbYL9TYena8wCZn8RPM7TZZ
Hnc3fYbxNeUjnai9OoYPsjnomAthu7tMrk1G10jSgtr21jdd7K2k1rQSXG5M
H9/FcRn1Qduwx/da3O8r0ZdORdKIXqUYqh20bYxRgFwMtdgo6mFotisGMBBo
DxeTitF2njy5CRqd/jWziy3vXZcPXXzcrdisSYyhBfxr42gEbDH7T/1dpZ8G
hU5aPb2ihACoYyitZZNAagkJP+4SJFIWiSZWL/jm0QUlYdq0lNPEkAakh0c7
BUrFL8wWGd/ClWbAfJno00GtEyAa1tVJBAmbO2U3wNBufjOTWdPks/CiHqc9
H/Hjn0SWsmY7ZZ3bk20c7Udi+NwOmgtW6pm8iu01boRuu5+HPIIF/1MLk4cv
StJLrnL0DymalnVl3E1VmZxSKVcYuscAxEBbzfwbW6Xw8qZRaoHZBKOKmVFo
V8BgrbuM0H5U8bTY8w+wD9kE/4+8Vjx9/VdrXO+CX0mnfW4xnU0xQ1knMj3M
vuH4eXRmhQ69GI0r+jNfrD3y7M8U1BZuvfm7GU/H9IUGlV0LBUDEAMfRMjNu
bUHgntw9qJBOtfA3cBfYY67DO9jpZvi5HZMTZB/x8UZhMhm0YG9rmrLTaCZN
lDflbM7s2YOQnEmuaOjlwwuWnIpRgs7MwB2V7F1r35lgwJEjdg00cYLbxd4x
EPAYrS1SAWrC8sQKmLLLBVutRasaqvlHEm4ETtYy8Fa8Uawq2FF97PcmfwDa
kVUmoYcDFWkCgNguMJ1YTmtO+gPx1DBS/gMPTE2+iVSSSaEt1OKW0MRi8I02
lRz72PTkT+xlB/uA1jlU5SrM12hN4qX4ykorTe5ulIG0FNrJMlIUx+uWCeAq
SBMvuMksIvmBwsd7F1k3pyTe2awRP4zWgPRzYSyY/9pnv/taDgXtJz/wNEay
0y1kLph/i/FPtONgnJfoy3ueiAqbWLsKGTZUXfWmLE8tq0w9Tf8paTKgnOt0
r2Pqpo5OjvmM24J7aSKp/txpWCimun8+tWKPrepfBYYo90GYTliENIy+GOXZ
0xZO7hgXwyI0Xv7kChj5GO8STtNAZTVxQOH9ooLze2zeJG6ehOsE6hn7oOcL
IvS9JhL4sy5dsmFWk3jlG+aBX1s7H3pCLba2aFEoVNlzLFIC0EUjIQkAE8RU
QMnLDiZHkgDpuCaRMbWM+R7h6shUg5S8MEvisRc6pGsKH4eQeoRgtLYnLSt/
JIAZxRmjc6GPOn1E1h94OQXEtqc5S4pzDWHdwVm2WfTsNSmH1z9LVxyKAGVL
HxT49stbOb26m1R0xxjRckVE993eu36BWr6eYg93Ru4S8sd3ueJSLEB5JGpq
3yiGaLH02mbsXSZxMobreSB49Cr23YgAcL0QeQ/XFaq8qHSca9MQZuTKndBJ
daiznu8UlQo/S9meo1x2s6NnYIS/xE+ZGKsrEfQBX6gYlqs0yVsBHZnRc0F6
XHKobEqf0++g2KiAbi8qcIgMd18PK6/SpK5QyfT2OLZc+4InUdaVUhVQ7yo1
Y4rB4/FpdOxAN8u7njwQPg4I3Go5hqBo0MkxnQnAcmagf1FM7SmvSWncZwRv
1dqjq3cxsdP5W73LnviZ2EegSWYamV6q6r7JHNE9o6czxIqmZBLiWo490/SX
me7WhH5jlfeOwB8+GM/a9cgzUdVsf3sKPfzt5fVvl3dLUA7rIrDreE2mq4sf
HcfoawAZOyuaONDTUTzs/XZOmwspPsmQIcwrKxImY90b3tefitYqSgz7r1uq
RKlLlKnFmRwKkNq2mLOdWGMoPsRbgkVxC1l+3ePtLGKgpPEOAo4nAPmLGOsk
tmuDyGpTDZhaX1jlezMxotWQaDPcBOC/IqlclpPhbxxUYp7KOrHWJGsm2vUA
jtGucyrXVBTwrifuQ3/pe0A8chVqVPW1IFq0NIFSLXZLDK4Ld/GZzzhljm4B
qFz97zpAb9TJMn9DnpUqyPEEICbRNXaG51/oSzRoeM7RTzAF5gL0vFyQGSMf
cJ5zJf3hyezi74TSfLKBVuYmgs95wW9cIxHbcP35rK1lbz1PzEbjTdBF1bSb
7eahX+KRSbE63aSbcHynv2Ji2NjpgT7NlVQQi+bp5uyH+RrRc8B0dMxxJHQe
0/Ho6lFhzC7euOX4egb/HCd3DVWZnUmlLmXb3yL/ZQ7oz83Nwd6KKeqE/7Dc
1Z/uMBAomPsCPdzmbB/fANC2qqAyWiYc/2ilpHrAOM0CA0Kh77BL73ExMsrw
KbU33pI1fi5j7gYHwxTJyhqdS64G7NnIqau+uXLoTi4Pl3OUK++7u7CWJv8g
m82OdCPWwAmRjpZlC6Y95dNUEcdJgMPuLUZg0+kja78sT6/JQNxReNXE42bN
EKPJE7aWUt6GwALmbhvn1SOKtrYLYYMiiMXVCRVDS2k/678YbdupKnluVWAC
VMvqX21UqglzNTi6oAFyoLURKKQ0fizW0FHnWkbeNLv22hpga91evEXTAoHz
EJAdEcQXCEOYR8PmGvxyWe/XDMUkJUcm9ZvGQj2aWHfmjsvAihocyunJ8Yz1
bn16iXFTnbeoRXf4rKTjIcRDBHOroeZjyahTkz4dQMdfAxQAtePJHH/YDYwV
Y5qC6HN/l8USHZJmchehDUf9WVlZbnobMRiX2tsBt1wAHZbSPwcoSmRSqAnN
jcwzsDowDuYrQ+eAPeIn1+OsvQarxEo/2WoRJsgKxqLEGzhf3P9JieAQii6/
hV90d9YOd2vJUapxtrtTf+hg4D8/03zOl1v7m5BM0757RBJKvLTaHXFOTELB
zZZyUgi5B1Xb1++oGRbYM7fP5n5f22H93iavqKl0JvxRirLX/X3owv5x/M6e
GcJ+CosOAsQnDYpriFu7xM8j90ywdw0k3O7FpbYhmSl1U8mzsE8LdLnannlf
s4jbXYLic9DdsszFCPkauGfMY9WvIOlq+BUeOYFO9w6mWXZuE2CTUuNjqefk
nsSMM1n5baXEf/t6KPD8qZBi+JS8r6LIexSkNd4knTcuANQg5y6nvCUWf/GK
oP7ulhy/g5gEwa3pcgAja1nxR0CNE11XlRNlQF2IME3soV/TNi+uA5eCFtha
elWnONkFXD0HW4dpZeD42/Iguy0yWmBSPc0Z6isJigenuEuZMTJr4h0PxqY+
O8neIdbBMQHWXUVTOztXZXvF7DTzBYBY0IzY5phzkOYZ24CEgRLkSHoH8CBV
na+asxcxu/aAttz89orVRI++Qru3vXsKCI5m5xBvVyA69EoR4248ek3AyjJV
C7KMQPBfa8n9kf0mtsH+ehQ4IcLLHxU4Tr1NN1xz829t6YFeRhhG8eWZISCh
jP4/vemzwwY+1Yrq3rYvYAbn1o7D3OzdVVo3pLvluktlQvLMf9mPV6SFp2Cd
NEDh4KVHW7OvxjQCCFltY+Agg8zNnXTgK56cT80b3pi9PcVtjSzU1lWMyyww
8XRC0B/yEUPOppLnutWZIeXtXDJh/pt3Mca1JbYP2IgylnTDliPDtOVtSz87
66OpxDqAmdBbtmqzpVCemUQWdIeZnipUSSDAcTg2FtEb6Z02bW4VuowPOQcq
jbU23vTNEsd6aM5WxEVRIx9ufzggOsIjjzW8s6hpA3c1uRjadaQ3DcpObwjt
sPkwrwAIdgpMgKbol5Ayk7xpB7MI/KXcFPPILx3TD/ZCK3aiPoZkMbH3oKCI
6rzNVaqw+64GwD9uPzFwJD2sVvBme7DcS+PlSUcCxvVvAzg334Qvoh1Wj3qG
uhHx8q9rYA62u5MVQKSjbrY2AP7K/nez82tySBHEl0XRccf+GM+I59DhhdTR
SflNVms79FPpqG3lPXjXbUTNeD0G1ZyTdr0XbykAF+7cse37gpIqL83q4NJi
ju/rr2RjUtaFNMEZ65PJ1MHY+nWBt18zSUXdiwlZ1NCEwFvjMICR79dNr9f0
nytquy488G6MtggkILFB35qEV7fnLUfwro9PAr9681+29Lp47BdGdepQHbXL
VLsluZjMjPjcZtQPM+hMrJexW3p0KZ7vZi7eBENwJ2emhE3Et7VGgtYg/k6I
00xvkRJGYFHxJ6fuxctFCl5W+R86DZAOM475eO5CBPJddUjzwU2+IhU0D7T8
r9GauPOCs7aXThH6INqH1NbL6SkN6gKMgwRMXQ7qENifpef9rP1TR5fitRfB
dJZs3bYTcPL9oPTd/988KJmyJUX5elEHNDg7zJOtcyZLtlGYV/5PD9Gh6fgw
8xWXk3RmSLxezW4aSDNCRHJDJUlHTlkZoX4y1Cb+2RpWD57YYYpKEnxyG231
bmdK+2bqi6HWfIniZfjc0St2aY+84OzbFzUFlo7CROhqfohztlCjCjmGAWaH
a0jiLPtntqGppIGOGN3Hn3lzyMoKcXwFSYf/2pl4w6wRmwCaFXN4rYzcxTFf
wB+6SfsprLV7HAIt7cMMeLCtkZ/frn8JcZaTck/GAU7z27rtWavRCxP6VDUr
iQcblpaJVCY9151z2l0ujSi3Pe1+ndskrBE3h0zltT9j0VnPg43mEYbtpfG4
ND0rvdf3JgUiY76nT+qi747jWYebYxbw/Ln3BYf8mhJ3hv0r9wJ/fWxfLVHm
uAnYy5RYVPFbJfuYCrUuW1f579Xl/jpaTbafnBUlU0JxUlDVyrmRMsjogxp3
YkHJ/qWvfG0jPS/U2/I2lLKsAKIu8iSGPdUvNQd3AN7IfCBwaho002X4nMyZ
ij8T20DFBcQW8Lz8e3eHw9g9oEG6sL5bCTPJ9nhrpOiceFbpA1KOkCMPUrkf
tB0yG401WfHTM+O8CnW6zqSFZz70pTx5N0crPnBYv7QRLIloSxrlZlQIKL8P
i2FecDY4dXuZN2Nr0vSlzLHt4hCKdRXNjiJL+6skRnQQ+e/u0GRsdkS5bYtB
cVDDGWS6Zn9aKBALLIT36X0RBOBgvwDwKt6nxACVuc2QGDI4gMKoa+f1/qF7
B/2u6hhHZKHjPoFL/wfqzMzjKdRd4XUjoMB6bc+hSK0Xscy4N75pu1Eb0kIZ
ujYIkb0P49BBomGISApX7GL2kSpudzZjy8MpNMGiHMw8k8PfajKTevvFICUw
f1KBDrIUPcXqMs2ObayDNSOVt5TXDkazXSI0U884ik8e65NkZgYOw0MdVP6s
JuAu7hCa+wW4xnie6cTrXjegOzL4QnkPirvk4py6RMB0TwnY9/dUSvsRvqs4
/GR668i8NK3Zb4Ve+JTaRbuSvGE9LVVt1dUHgtKU2KnSsgB4XgoPpWYEadAj
R3ornxsYEg71oQvxBlRz0YnXbDev6KF4lkk3mif44m/Fd91qiiKK9hoDgtA1
vEXthjKpB3N2bXPkTBmAl3+E2vzzGgJkkUK3/eMARN/iBfrvUH/mki4BUJEu
UVPaqksgjRm4ktqnTVRg0sBe8CDd/i47Un5cqbicYDQsFZ+Dj9Nn7CkU7qyf
KKL+3W8tTL8AitMKudl2n8nrE7VgEvlYFqq5P79/w2N/6HNwwVmWPyRpUGQ3
wmCxi+LKUOdMyb99L4GYGyte1zfeDnh68V+Jm8pWzGKqH2rGNK5CbwOUDSF2
mU6gdZzXWPgwaQKo33UtYLPxLepphNEoS3cQe4ofzCio8LCrrk2oCiDx7aLT
xLvys/5uanBTT7coQ3sC5y2xI9xaVVucZBZnJp7Qc5VJ1TmHDXfqcOsrcuZI
+Mbc4X2j/GHmYDW95CO0dLHjzGsgBkPT9mHO7vZMqPH2xk98X3umLHPfzb0e
7kurqPH/58Zho+M26aFzB2CdOSWTOPofHMM9F+xFj7OV1Kckk/iwGgDSkm3P
Mk6d1FocyYCicoCNnOMMZ5/unjMXXmUMBuRfXZfolAIERUne2t9tktUqclFn
svGOQZRMJaG0cXDbwb4kbRoIhIpdR8kLxdqHaNUG8p05fObr13AnXH9CWmx7
1qcWxn1ht57hVB2KcjKbKKASmK1N07XU7fKYGxn21Fi7KxXFL60d2wM0qiA3
ON02SdgAu4j2W8BXuslC5UgNq5RGr7n0KCTzfnyQ0oQEbwQyGeZS3KJHP6iN
hisNzIHFsbTu+XqOpIMfcrCtUP6OwF+OySDKQ466N0hHS19qW4954+ICZmnm
gH0Va06CbTZcvmX7LM8iPj7wbQ3JOeWqlIjaQbUiu2Vn7kfv9Nd2NyRf8edm
2nRcLB+N3zGFJS/5AepTrILcLpsQXQSg8pJ5UBdux0EMs4KtKl5cxrUuAXkW
/WfAGCzUlhXVRV9z90vhuppe78xSCjVBbBN1LNkplmwDZNtl8HYxqWppuHki
KZt+OIbsmuFIhF6KkGC0L+MQYsbdii9ytK5lwuIoOGsj0Eb/FSSfQx/CIo1Q
e02EPUx2xQmxoL8Zzz3vZ+NGBBRYANP3jLnH2fh/oBo3YF1sx1oWjpiLnaoO
T8/G6W47u9Ugru4XxtrfONcBYS6NhTPtybJrTJyBMNNnF4uxPN3JRVJgpZcD
nN4dKx/XE4bEYN4oifWJ1DxxFrpxz5PZyQAzOzcQCJeZ8nyKbL+XaQm7SC8s
N7BR7fDSoYnu2y4xLczEMCz/cFPJJLrvxj5ym896ORrCST5iTbi1KtE+jgnw
EINp3NFRBAc+c/XWJ+RcdieMd/g4f9zeld5vtZkr9dI/HWajJSw3HZoiaBJa
dA/DZi8inmJDoc6WCh+cT7yNQmD7tMREegK34Yas3ewb2d9C1bIv0qrYV9m2
ao8LRTqRf+AeC7qjK/G5m7aLWXYw4a/24j3ADQlq9YeYIQhUtj51ewJdx4fs
fe+lrq+xFTzqstrxQBr+QeXG4LnGgu8iltkHlDECdp7RI9/fkUtsYh8v8Nel
lLnL1+0IJppD4go4HEH+MI2EKQR84ouVHh1T6RNEjecQY7HXACovX7heVVkj
358r1oetllMxtXRvY9XLqsXUsvKCf825mC8R4iFqkP9WpjknAov9foJLx6pi
/gwEQJIFtorTDWYjUWPK2mVt1P3IchW1nfJjrouEHvdiLP/7PD5F1rndyKEO
pgfO2PvnPhe3xSFGTN+WnSbaFTUSFwl2p7IwGPcbtA5lCLRkobf650CU7v7K
L5m4bBR9dTRHiwEAyk1N5VOamfDEV8HBuUDY254m2SxZhT7XI9Kp7Vnr9p8X
fu7zG4T04ML8i+mZKbJBRvY+K7FLrPeQhwVzUQWc/5+1kAXMTdgZB+f0zDSt
URyYeJwEKbqcR0ZWw6ITuQRbsmFy0m05fKDG7KKOaCrmTYFae+ondBOObpBv
7zaPVoY0XiZVRIH2dtQD1QvrZzq0W6XXxECRF2clbyswLIymFok4fAl+L2/a
+o7mbTixdr0B5zKOetXls4XBx8epmvuE6V9Jw7gbVpHliMbUtiAX6QOJnaRo
bjOlReDBghk0lI2k0CRSdVoB7mo7aNKwy1vt68oKWsbHl4WvpzGOoC33Udor
4lhieoWFvDWn3KElEt1WYp+doK9rokDnciEh/X48BaxS4RCcgOmriHLhNHxf
1FGSoYzDDjuc8AsM03BgE5K+7p60cyTQs2Jv1r98DE/1wjgrG2P68aEXDPEd
njOE8iWkS9ViwrGgkxDIRNudsC7cEMZ5YB0EfEC184h8l9aHhg+NNC9ZCfoA
GQXprLqmAREhh/M4c6fvA3TXbbJYiODuee2e96uNjntf7uUYiXr1gdwQyv76
wOI+NKIVDfCe0Mviuw3PMuQRN+4Wdyj2vPJ5CMNNY5fMGgHxwlQwMTZSPG/z
5aP8qLEl7fnztpr6GonxNBtU3CGp8VvfZ95w9JXrtqin2DDFgmGWh01TS9IC
yDTZvEu7yFAJDtrIhpcMx0CqBASCQl1VRfgk9vq6FskyIF9AZqkokmq6GNqs
THtHlIGHlHApekUt+v45VZP8uWWsSm36KPnLlH+CVOEEooWonX3B+qmrV4qk
piIj+95GCoaOg14JRYWVddcWNN1AkOpzxrmvBxUVoUDf8n92B7JcA72mW5BL
yZ+Tac4s+Nje2AiCJVsxp8hVleXBt8jgjeDVKq6fKz1BVmbK/ciaIkjm7WTe
JN+uUo2K4bYq7OeaGDt0EANSCPYKgoH99t/FovDRexmTY9slqxnQt607iO71
btEMMExbWr951jAaNG7cmp07lxXw0PKpfHnm36L5nd7Je9Y73vwK8eahtOzm
16TI7oglm8mzx4Dpisn9WnKHN0yvuFxunDhY/boMlNj7rTgj1PiJBE+oac8H
q2GXZ4kfJJCpQMJjrR5vAK2sz+nPaoggaipT+EfEXBDaKj32wTnPWhrYGuyC
FpJZy7a1vsmfsrAuz0539wBnWmC5Avy0EHKNqcKNuK4yXykDDsjk5QSX9c4g
ut4jxwBlhhmvrwyH/Dfe/ydbcRpf3gbNyJe77RNXqS52eHVcnj/low2jekpC
1/IUI2DK970UGhqAMl4Bn4nHmp/klSIFY4aik3GtxsHG36sxZko/BFGk5f7H
GpEPf9zFUtH4Ta/tfp54kwRNRlYpaRltGNyd3R73VjQx/D4ybfRGBFOe4kT3
2HqoHi+0LJOVfj5Nc3y+uoQAPWpxWIFegeEZwhb5KdWYq0sgtBJ/IDya36It
tjmRJyFVfTS8rYV2MmnMGIj6h0f6ca7j4yeYF1Rtq92lkZfk8TFI2SsINFc/
aW5YWs80KZWW0MZXYdmcCv6MPXIG4JDkSUqEybsCjqjvEi77i0B9X1cwl6YM
QiBLxFd9eByZit8+o6E7pzEvbfZ5PKWHqhGjEfKc0g5D19U23bT6BtxPeSXC
CVhKzlvw1+uR61bnhKlrpd7QD3O7rgVUXMWWbqsaqlAnGUSyqr7imWpcidfF
9dQ09L2uQxY4L/PidlAs/2HZlPlm784W1ohIul3hE5vowe10B0C6jCt1f01n
el580fnYY8b8i6lTZXKZ4xE01Guv/k+SmYYVWB46N7iFxCuAgC70nLF8jsKy
d0wPAh5oHzu3tlT2EaU5tOq69ydmGGmX39qvqIL9SGNXacHtz95fUv70ukQ2
RgFo4UQ4eXsxlKDsAu4xwXd68LAysfH4K4AkaijABK5eDYhWwoQSs7en7qLS
q2cwEOdacIzRMl3/eUH7EDB+RYX8neI3J2/nRw+MO2odcFk1ErDyC2VhOFfa
yRx2kxNbcHLvsY6PenfA/COWI3B7FUAtGhgfVs9zJRdi2u7piPT/jVZG6FBj
KJOpOSSwBSrn0X36pw+S7zLsXzYQI4i7jKFOpO/r0t4iH4aM34OzxAM/Alnw
mPkocwL5c2DnwQOgjvJbuU8Nt+WNA7EDz2kwTyHMGiyOfPmmV/EI8qwHEy92
O9GaMDEyinA9D80Awv0hUCDVkNDooUK0PBPKE7JU32lZXBTCPGLXKzkZEehx
r0Ltm+UTz+N7pi5iItrZz5wF+1oXFscYh3M5CPgUPyv9MMTuTaLFujSCaecn
oDO0Sr//fBV9BSLS/CyEfo/yGnQgAx7i1ZdAYcgC1D9rBYXm9K5cBUTtJdS0
o7rBE+kq8v8UZo/gcpFAMXz6IOGkzzAoOo22ttsw6SDnnnQ7xkZ6nMjHgEtS
cSSUtEF58NcFjWJJ8XkenYTeuab5JGOJuPabQQPNBlJ59jb33yGm58iRkzoI
1wXBAzXherSSXTSUGdjsUWMvSo7TsFzS0sLS+cAI0XhVdmdhPtW7UKZOqLvl
wO9liwaLEjL7/fr+CMUlsElX7lxwFSDF1A1og1i0LiXKv18oIUVhIu6tbdmX
aoS2FcNNZ3kMz1wct05okKCLhIayNhjyN65LiEXUH0t7pJ86Wo0t73cKvE+e
vCxIo8i4C8G1/mTRhAC9e2HPtYnN/3DTbTVFhdY0rATN/UhF0eSoRZVtuD5E
sJMVDZoNsI6+n0RShgV/KKE3VrGGDiI9kc8c9BpAIga5bQ7kut6/DBEn2jMv
N4fc1P8q4BVluOWYWPvABubPcuoBFmXTuoyiJ4StYveEQ/tNiop1mWe5aPUu
4uzZD5hwAMG6N3+H0OSGi0tec0DQlaaaKIqig9pyz+Gp88vDzroLUo2KLC9S
TnovdWyCr/iycLHhvVDchubhXMX3xAGT7oe+32vcag1Hmado6rcY1treSrwJ
zAhlDaKBhscUsF1S6XfkI+aaAvbrvCwBBPgJo7H+o8FJ9LFTa3aQOxdzI2oM
qNK2FGBeBXnf4gnxa0U5qI+RMRjC13FBgQxsiEPjTXf+QHOm/oj0tezkfDSy
mLZ0ntIkI4+NTHoIZpVlCAS8g0aPdWtMCx2iOKAD/QNfo/6IgDMTXGIYdAwV
mmpIqzyIgGmo+PayPcSkkOBMgciDYp5+m4AbKqhYoNxEOgurDvpT54oFOAOR
EIZFUe6/yKpPLUMGfx0xc9z4lvjtukzJAS81Gl4FNJ58lWCk5mtVcpJEofpo
gM7l8q0O1uETswfRA8xi91j7xz9x8qVlXdpfAn88WJTFE0I5YL6vaxbnd/ak
1gDORXam0cBP0vEjGc637C941XqQ5TtHCFjWrxFIsw4OH0pGKknEwaOu7hqw
WqQVKwvBIU6Ktc5u3AHm45kR8fKjNXZ+aWTqosR+aT7OYvtt6wf48vmNkt+u
lUVwsz96kCDk2J+i4Ju6MKzBwfBexL4lEMlJnaYeNGprhjGqFSxtxzWbOuKY
Veb5EmGn0TtvMu6ASfsEC8l6pMPSVG+KzJ17qpP+T39pE9+qkJiTM9BuKlem
jU6AyP7w+AuL2OqHTqhSf80eRI/3dC00S4k/q5jU49jGbB21izGGXG05lOh4
EvFqwLF95ECVcUJ/BgzNaDsrI35OxgII9LY4CmNE4dTQWM+mCFNMyK8S2DLJ
4/RO7MkdPa2M9C54EbzJnOFe2Gx1eDmULIgM/7DhAg2tF0BPW+zSM3zxZ17i
1Sh9eaeOrEfRueDZZrXiSSh0ilM6dWBNRs3W+RS97LeRPKJyxcGM+C0FPlDe
2XFqH5UZa8TP8Wwtbm/x948P73OhdYZnsZgxCXmK39jS46YDXGf+SqgkhtTc
SOyf15WQWGEsn3vkM+T6aYLnHkkTUTTX9ZcMN46zw7Xa9MEH+2ovCKpP15Vt
Y/HvXCYuOpyRo8h5dIeZMb3MooumvS0+TTINcsmlY90FIClioGG7f6R294tH
Wl3+x1k+cdIFYpuioo8EVoVp1khFBP7dUoJQAAwhEdgEDRMwtIl7GySC05JE
dNmdaKop12T64XtDY3arNrUCM070z1YRV5bBBDS4VhqVyUoRTbsDfo+KU0QL
hUOIiz9f8qZ2ri7Af8G0s01iV5HE7iTpTYO0w/I/bUBQbcmxPgvy6JNY/UQ/
8AJJSpegFIZ7sKpQ73Ut0w9wDd37rGBvHgqyfb1W6Vlg7/m8vxQ/vuH/l+U+
3gvsplQJ9btGCQDPt8fIlpIK+m8rm2hfdrKdYVPaFxjPG1PKG+DTO3opEubk
wXaFX6Pv5Si9JZkNjVkF0j/Wr4jIKS2SI+veFWPJPQLHaILrG2RbiYTEpGOw
ksDNCPGgDNguEgKvE3KXJ0RAMnDpXjawpyWwixfojzMkD3qf8Ni2L7zMYu6E
r8cNGQDIrhYqrRDpAxk3PX5vc90h5bhtlf2SFhbHv9IWPscFDmlaoSI2ns3Y
smIUqti72DGSf+ATKEZKG37v8lVNo3YpRFRnNgm7xKqoJgkoqOnkwEN9ub3h
UNVGxB0DSQUWlA3jGLHZS5+unGL/vFjzpCTEn4M3mkg4lDuqaF2oEip6GnLN
uvENpQQdkTQXXFlI1n1aJuD1gcYG7sdNGT7Ufneys2WcbXlJ4WNivoMlnrxC
dY3lGYiWm7KLoNECsfNkOdb5I9fkCjqMlq6yexB5c/liDFS+Uc6BrsH5thIz
4iDDLg53456iUWty90HxYxAGVucTaavayXbpFW9xoxkqlPtBpaWjfKTeqC2E
4EORDV4+OGZyxCCFbsd6wCeTcWgDQmjsuM79AOZC1nXzQhnT6QR1/dwybKef
Qse2U/GOayZtIigMXi3lI3k3XHtR789Xq3DMQAAEhOlKkIcvX4Wk5N0k4ryz
rd2GBfywgUd8YvbW9gl3HdZ9IPg0BNwCHKnxykP4Syk2HcX9CThHtgEafEto
hoA/60T6lRGlBKlzUW1LPYEbQDuP648ub5HyWZCyWMm0B9Q7DM1yhYf4EPS8
rxvmZf0TiVoFOZnFU9fRKVb6mMASkhRUoLerd/Gna1/2O24c1mMZgHLHnmNL
0xdD8nL4Hw7Y/QcbWJwDMK/GezvTLpzHt3bmhd5SqOsEq40HdYD2lowdVSei
oLq7lHmA85zrPULoc8b86PVf2j8e6zeQsZxMGmqn1f6lWOP84E6JjZMbC9jt
f6ySOMM4Sm6yI6SNwCpO0M9+iacup7CYNQj/9oARQ2j08sX4RhQqC4OHXkp3
rqsdCWwzZsz9YoizzFJcHoMhem2WMYPRB07Ahe/TC9NdOQNwjIkRE5y42ggz
bjvlJpuSfG/AimOaMeZVlKWE7BgpZH26psjE7iFi1vFMb4iR6f/f9ukt8I0s
qCM2Xqz1o2eyTmeoy5gxTrMBD6gQIgvLIULOhfHOEwe+K501VfzqpSj0zylF
aN1Ip7nb30kOgijKsLL60q1KU/lXbpWKn8C4GWoDDndAIOhLGZ6w2c1w1Uj7
v+uC47TETBaHbD3nLKP1WN0mfXNGbAqBAvKKlioSQUN6XgAkw4tPKjER/eG6
GwpCABDDpkvd3kdDUuCVIH6QnuYd9uDqXwAyVoLpiPTKZxAOtR0ja95KWXuO
phogR0zspVAL02/jHoFpaMoAPVvXlmhmSxgNEUHQLoJpcNXo54pNCP5Gb76f
hggcgrwPW76TaH/cBTEgN1tsHsaqhunOUAH62Y4TeAxpxG06Nvi8N/7NqFoS
T6Wi0JnljTXZaK2V040D6k8YZN/YP2BFr/fwzoF14DROuaZheoxh5pSesdfX
gyq+QIRNiOBMbf2+XENZ6qox3UQ4/+T7+EEC8Z7pBU9dhZ5I+XYr62jktIuU
ym7I2+NpoMLWsS/tfz+5/GxKv+00PZmVgQYHDldZoT3R9bMO0U08P5g/K7mW
qT6jLvTaY6IOYVl4DYgGpn/F0T8Z56h1J1lE0bXzN79RStRwPkMRy3HoeVkw
rnSbl1ix2JxGdoIuoIZRRfWoT8QoVBK7kWkjE3Ik+fkyoPhemqjec37uULJF
cZfjckDtp5q74ioPMMZj4dJ3MAyTVD8laqVBByVPz6NA5UALXOMnhSVsu9FH
+6Z0Y4S0DKpSNTzTqGrqH1blhCdihU5TQnx7g/ZzwV8vGXMiyahxGAZP0Plz
sggTEg3OOgsWkjYbvNKjMhHYWqcOdFmY0ow0Zab2aZ7RTtAnp0K4CjmSi935
e1QqeSo+IXAyTILzVoviTmESn/HNV9L7UGzUaOX2EpWeDXc5Oscjk3ID9HL8
gSIQ+B5vQ/n2D11HoZQrA5w4JT1ufo7S+oeKwp77c/Cmze6Gnkyy8DjHY8lj
y16y57Rel9U1eQP7CKV6+IM+H2vb4r/9MfcqdosWJJ7VYq7ZwK2BkbgAHoDG
R5CwNmyHIup5Z8ucQ1MxvY0q9n/LgQD7unbjX5IlLgfrmHAg/KZxHy6M7OLC
W9GusALpwdbPT3jWkq5427ZMqPe6tsbJhK4uxzwCe6qAj3VrPT7Eb+dd7sib
ZFUbcSXGOIPSuRXkd+BLpkgQI7nJ8u1eD3nlxK1eIsxIFOZw7faSwqNg17ul
S7rH26gjqNr2OtqRSUQfVmH1I9BzyNYSr/YfU7Fm6Zp0JgMikS7iOft1IVpS
1VzYJJpfGPMOp1SunMLpye01m5kAJG76OcYTI64kEVKg7gKYI5Du9HNzhS53
ROO/UpT3welGlK3Xo4a5r8qLJfVhKm/1RBiX4wbrmX8mLdY8gkpbx0FCChIQ
dWSfByXHZtOti0xixuTGVsmrvU/t1SXX38OLukcBPqI+WVq6I7kcXUgoihlv
moTDD0PmoWQM1saNsWiuYSjhLkUV7baC0ypRF5fSmogMKnZNQMIu1bXDO458
Wk60pGmM/OsAYDSKszLU2Jb3AfqMCmSoqUsNFa3u4kJNtGvKXm9fZ+hb4C+j
UqTKVcBkarDNMsrekylgn/whe5AUj8TIYufjwn7w6zMTxQZWSUjQ/HS+RFje
VIFtr3rp/r7XnjmSyQ6y6ULHHoNP19vpXatx9UkG3fOnpPyauHgTaJeUEzoz
5HhdzGBeCsomXSZNzejFZTCapgXpfKJi+2qlSil9O1XKrCxNK3q4L/Zy5qxg
OwYWK1FJze+XnEMqK9nHCb8HBPemGeQEAGr+FfzSR0qjDtstQuWlmFNzQJhO
AkBxkwEx0EnDxsfUqyOIi49c1nk6RU5GoLXjzEPp0dCdtRujXRv7jDyxY6g4
4TVLgbTiQ0shFPkjF6kWWdNJH5d5gpiVenpJhpcgaVIoDMU6pgEfenrOzeh6
9S1c7aOMxA304UBAkVut9TqkFTTP4kl/cKK83Nnv6ihnv0iInksZsBd4wc4b
B52ZAL2hrb68VDLacuZcMZoKy9K3WNubs/s7ygPmNVR0vnBe1BjWUWjKFWA3
ar2N7x0k9EOf3QxiceY10a2xnoxPXZGGnQgWu0HyVnB372TRpN/1bSpcf+8b
BRMMkdlnb//ON0CMTChmdgzEazeTbEpRXWZlDfiOf05YpkDXkMZgJq4m/Zhe
B4rJJpCJ7qv7NFjfhvlE6r4TYj7IqM7vDl1dofJBVaYHkitLAwbGEwDatxBr
VoocoaOPOFztj5Hq5g2R6LfYw6nmMI21PcUuVE24h3JW4AXb3CZ/NTKAmP5A
VUGvfapIqilAOTz7q6IhM3p6DMMwwyVG99IR34oTfZJ3Kx6m/T6Nsc5hVleE
8EBn3TEHNFN/3b4vEjWX7KY9BUuZmJ12elHoNvHkmSErZjPXbFRRPQv29Gch
F4+OKWgymDJE/kl/jD8ht/fbTmn08UtgT8SYbAIAIqByQneKJyLs2uEvTkfs
1/GT4LLakI5mvPz2j8QoaT3XTCBx6L7khWwh+BuhKRfWRy+EsTOi9+wlhqKM
M8DdomP0mqTuX7/1LGgpwYgFZ25zzeWs8ZKLlZOsD3MsrW+Zo1aH6aJyLe+G
fC/9HyIprqwYO+NAe3LVoXSo4fiI8rIXczUkxIOC78f1gt3umQpj6MMsXbbx
4G9en+xh9xPaRZp8VE4JUXUxL459Zryc9g11OpKqs9LjbD3o5vjPhFddHvsv
DDvyy7DcgdUNLi5bUjyNtC72A7+a3fMQ96l99j//uBlMBySgp+3ORfuC3XV1
aZEFjMYMQZwpWNN8brSfMOwQzIVRSt1HXul5nNuLKWt+bu9lb8sjrADt4/Jj
UfVgcTHJXqFMPKfTfT0UbuWDHy3TaiP26k8L7L/NgyntwAvpUfQb4JfBNY2/
MRejgxpfyhqK558hqOiSl//avVV3EB2r6177g6UwJdVlvQWy2DKI2ooJM4xY
jLy8YlzZ/jZpjgoS0B/Au0CWLVDyGTIFn+79GBaneUJhLosvG7K9MbrZW9U5
5/T4zc3kNpqd3xTVjiGn+z4xuUVHiLz/xp/1oPuRpKNuNv+iRnACrGg4pjpc
DrTBCjM3r35IFSFdlEYzlVYP6dJhV1HfArm9NklF2UvrZDfTEUpn1gkWU4/c
BMxUDCGHtS/W+Kr70j0vc4aB6Mx/G2gbK1aEC3nQnEGVhzXe6nqTxW1K+JDb
MynHK8AUiPJm9c2CAS7lWKwwEQDFVNA3WvslM/1ixZybmvtxST6wVP4Ih9dT
adMfK33WcFVljaddO3SQCB5aziqqsSIwVP1xm2ccxGUGyLNPonQUGJv/tY+U
wx1LXty+f6voKUS718hyBRNeA4+x3WLSEb1uNMKuvBWzylLVVBeVe7J5dh0G
rkIpuAR5Ge60xen/3rwNWzAH38G9Y0Vfx2GtVkFbbBbuIQu+U8UsIEsePHQm
yZafqOeOL1d3XrufjhNlqsHMtQAMEPZ45yBMAS7oMSG60FFMtQDgAmb0sj2d
dDQN81Rnq/CWgFRfWiZwVa819StJeYx4JE3oakdhjLptWUvgA3tWkvxs4cgC
P5DzOcK/e9kNBT61jVPT+d2hTxRDi+5f6CXma0uEwfVHpMQ9DB385yd6Di16
fK7PS4aIofGKltm6BaNiEEuYDx9bC/wZ4vamfM5nw/XO789shIPN1l0S3EOO
FJsEGY3wcD9Fk6jxNTZ/sV7UVtId18ANaLBBqniomPYM8ZDYFex8vCFO0MxE
7qAjQpeipEHP8GtrSfavbzuVFILwrgpR9ZBYvmbqLwpPrxWoRO7+wE5AcdCw
WgQgcR5w4jrjWQG59/fMlV5/6wdstGbVSbVRoC1spBzTgZgXTdrJKqb7kxGA
OcNdQDIQ4t7bqwkEz9qouzCQDA3VNu9mWLWPlI2AJhyJv4dUWV0woP2GZP+F
sZUKPiuYgE6gVu43rK6pQLjGo+7J1roRFK5qZidEAuMbhd9iU/eRRfpKwfap
68AQ4kexdZYLsnLCCDVMnNSgl7Zp9m0F9Hk7yThENxGC9C9gFfsSq/ws8tBs
tAdOxSygMJokfvcZ+xqrIa4HK1+pIpzq0WW5Omw0g4LO7dxmB8O9RFwaC8k6
Sz6O4J8W1xTnpsPVmdaMpLaYW2s/vLr1juh6ij/mKvsWfHCvY8sd0Y1bBeug
JSLU1mEfUOZyPqf3AEWmim+ZtGPf5h64z4PIQpAp/+/BLoL3XnvHA6j/tbK6
KkkUREzZ01PsyAK2kjZaGrxICmJZAQHuSxEI/Z3iVkrG8ysWMpTcfc3ov5OK
YQDWWizQ4LNtOska9K+sudRLM3ZD2s9b/uUiteaOpnd1kyWbt08cUfWwwDCA
rmhcdnkgGiBFSy4/KfBAe04QFNZ2kRvCX46FIaUsYjuWYYOJ/xN0p2IMHYtj
LDElk6qdKVbcXdvJAMk44Sz0YzkBu/kgLQfh6U5NXpmZGb0fLiyanPrSp2ss
ojWrrfPL4G+IagmOeLpsbSjZGVy7JYEKYSB0t44cpt8Sna/RxRFjFJq3vY3w
bnVBRnnGuaK+JIA2nCw7d4jOQSbAFmWRgmVR7o1qn4lABWPQOXpJKCNelPi2
zoWt6yB4oqoeJ64QZZ0gZVQ+Z51Mrtyk/UaMlxzHvNHNdEZaYdS7UFEUK6eN
fdLGEDmYt6Ml1Jp9Y9WbUAFbVmf4J3aHMgaRY/9v2xE+Tph7UYu8

`pragma protect end_protected
