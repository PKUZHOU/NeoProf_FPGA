// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
MnCtu54bAHmu9uIUoZhYa/7F7/Uld+6hoUih8sE7ghzw1hjV6vaS7d7s0XNe
uQVi9UN8E0yCcMzSuT6msLK+o9wJXofiDDeYW4RJ9L6gMipP6ENh8IVjdYQC
VUoKBEF/h/qhpQOjtr92A/J8GPUejv/SfpGK6f5jV87IAKxzCp+8CsMMxx1E
BBIv2JC9JQ5SE57Av9IGSIcT62bsnQRsWojQRiPYvGwp1y4QxirvUCxg7irZ
vUrEZO8v6m09o5bqes4GlbblQ0sUgdL3DccgcORFxolE6TQzcE4AT5sRSQfI
bsD1rNjyD/2Q76hIgeYg9x840fhI2aMbTUE6gnHOUQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
iuLc4T8T+uY4+Z1oFXGyodnOF0gtTk4raUTDgkWsh+dDqhP5ey4sB3BJ1mxi
w2WOw/nr7/SP9HnHAiR9HJL97oHZjIAYnS1UmpS3MpJrgoRz8TvvX8wPjT++
0FkMpiSMI/sCcjLyVq4crK39Z21jcqXafMog7puv5zgi3VW6ioJDjEySRhML
By9gZdNZ8HgozGK9vD3De5BTTIvaLMwA58IBEgI3w3o2/Iow2fQVruCzljiF
M7sHqzgjvuWcu2lzjmqIteTgielFPBZoAg+0F5qzLZks0FVmBKKtZiNky/l8
yhZxCY9rS25tobR8VZyJCFviuLYnKGNh8K7vituJ4Q==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
D/rXTZORsZzdmyph+2jfrULZkRUStuM490oQo7w7UduugSIgo1AR0gn8qoOh
vza9vY0R2i5TBgMhhiPP0ICDMmBXIesIM5Jziqn70quguKNAHBZsWmklu8wu
PqJOIZiakaZuyB+qc70Wvjz0JRQ8/rhum1+Ur3fLws6+bhL3o6s/c6tPILOH
LQniqSIyfZB8X6EpQgXFOMLIdy0E8UPRuLpSJvsNC3GHG1m1rPcpFS9s9TFA
UV9Rp881D5tGUlCvQ3IDsTtHxYjxlmybWxhBTGo1qgJqDARBaqBwVPOGScoH
lG1QK94uZks33gDb15b7DVjz921WH5nt3ohV8RIMxw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
bb13kELIFRBf1PanzklguqqHRs0FCWedEB8+p18GBoK4u+wIPXWYi1PyIgEI
QVp3MqQcXV2BKhBXjTtL08Fl4qRRMkjF5f/3deJ12QLgDygFqU9G5ebsRPIc
yA7TnXZmv1Li4RWdZCQpy5r1qtSeRKvD31QiZLYf6I+Q4jKjzkA=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
F78AT6evgWH3qFoILWcSZpNVF0mnQz4qq/Fn2E8WDLjuSt2up6J2aO3aDf4c
lUK9MbMlA/fi25j9GeUJLS6ShColW3rJgO4jiCrkE0xrDzInJXo/PGmvgS7m
FVEtnKRKHIQc58kpaZx4yLuR5KV/Nuq8trKEqaM878ZTxjVtb6IzA1WV3F/Z
cZef63qpNzhXJhbK0fC+iVqUq/mQdh44eJMZuhBeAj6JU4v5Rilye9Wf6TFU
cwjuuXaguczOuPF7mcz3z0iCc1dRjqROcW8HRafmfu3ED8dZCpMhyunNI+dr
+0Zv1IjT90XIK/4rNs6cpfZq054lasFdnZbOKBGehF7LR90XR4PSzEfkz+od
BO1PXD11Vulh9YDbodYokV8usZl5wj+Sr7GRdDZ5utfxJWeZwOAHFeVr4rHe
fkb18202wAvdrstoYfxwi+wWsCBb/4Jxdk2fNFhDFN9I5G9/H05D0CE7HSUo
6PhWWF1p1x5BVEP8CCxQ52+UCS4yLYSJ


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
sglM5FdprvWsY+OUE+H5EL+eT4jTcIvqS/r7fJF+nYiw4BMgYY1X6nErfqV4
ZyXYx8bHFK1QtrJ1/adrWx0mift7Vf9EOEDb16yam5YARthZlVLecu8BYgji
c2544WUKHNINmGs9+NJvLApw2FG87kjr6tK22iOGU4h3LUl/RS4=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
GjvnDlzuXfawrohK6pRomRdVqdlEDKovsdkcRZY8iMUijs0S0bKNBkTscyp/
MH9eaKcUgnzwfWnSaMMCBaOEbE+Tfdrtvadq1VBYNA8iyiQdzP8XZIEC63YO
kogwiQRpkDn3ZKzw93jR3//kUybrppTmxUeowA2TUfyiIpve5Ug=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 15568)
`pragma protect data_block
3RQuthh+OjA3WxaT73cSYQGb2VihDCCuVKDTfoBsY4zYfDPvFk2aRvumsRIv
5XiBi4vRmP1AnzyTADnOXAfgOjphPsa2dysMvstHk5tHdWbEJ/cHTtu8gk8z
TGNcDEWVlnUFHwxdUN1abIIBrTa2Vh0MZ2bw0VbCknqfjv/n7Fx2DaGVK7Hn
pg8mR/C3YUne4Fn6GWTg/YBF5/mQZRpe4Bz3hyxrS0lSHkTUN2bS0zDaAp6j
h/IlynHMSf2DZFPI1a4bkuBGzMdBvDuOR5es9t3LIxfW/mg2rPCmtXg7dREp
yUz/MftgWB++gCOh6AIT5ZRqrnH0pCAByjpwXej+tOdCgZYcDX0Bgso1ApKc
tE7mtc6xPN7FsI56M5LUb+cLRhE2E7oct/6f2J+l5J7omc6eHpFVvRpjkCA9
p14IFbqjM73hjosRT5uFVWPVd/4RZBRxaRfAmiZ2qQhqbK1F9b3R3CAu0Sg0
BwYp8sE0xRXb5P0pQsFF/cbh/8ZR5ZwuM648hjoHL0r/FipSNkWydQTeoEUl
+Dhp4JWKCx0f8fr05f2d0dXOjs+zMuxn0iTulRw9pLrg8XMXyn7PayovvxN+
bcNXLXufGuZoYorjGtu20rJcR64qoAHL42SC32Q19VC6FfnT4t0vRPSefoEt
CfRPNXmg6hdqT3EofC2T4Zu1YQiPdIg68a4PvJdSEJvA6ud7EU+Yg+oC9CRk
XwrSXj2IHlTVHmYUBs2fPYddqoe7uoNy9BgmOOYBYC/G8VUYxFRFDuxqiRDr
bveofuqH79S/qobAugMkX7laOBki8ha0Y7+RaCDxN9bGiRlI5VomS2Xu/hqJ
Poyc0A52CrQe/NpLp70QWlMHFoSBptpX7KcnhhNHtGXTEDKKKTGL29kmqsRh
tFDgAvC35HwkDzPPrn+j4iv64rkcpcKHF8Yaat4fKInP9cYPzcaudPVCLfme
qW4J2kQpfkHulTK38Y0VOZqmbXleZm7pp4dxzDtCQ2gj9K96/7mIw1Q2AkTK
j3w4PqNQ9TXfu971nN32UrDs6MYQlbDb/foJlEihawBB6HJpiZ2+Dxq3aCSf
T2KU3nIVqdCKVo+aNI7DoVmOoADJINFClSa6AeZdOYOwD1fRR8rIJP0Qpk28
hJwxeQCBVrn3r43wQ5eM81pUkVEiELFBSZ44S3k/CfY3wC7KKV/lw3bpBA9E
9f2ChMdEVx//9o/QCaYhs0v/b6gNLbiLHaR3pAKCYeoxnCjtsw0S8H2ndWOm
MCzZZps7rghN0zBTMEGuH+yk3mR6FEN6jPIHURU1GbttTaxUpHc/LPyBYIpK
SLGIwLPPUyIbBXHKhRTA58uh1adUzAQD5z2HXJujC5QySZ0xXsfrXtQq9ZmW
CnRr/u0guqaW8No1rPI9EzHAUF2boZ+Wh4Ql2u+FO0L336vBeZKyDKlh7NpS
8pND1t6GElIfVMSsVej9fKdCHn01aPqCRpCWpe9ChvMGdIWG0qGhFVrJtVs4
+lzvoj8eeKm1Nn9DgRdLjJbjzsq25yI0skbtafXQU4wL5aM+nBrsOnohBPvO
GyL5PjyPkKbVDLcB1tGRlBn2OwnSVyJweDa3940lSB1qZM4SaPCVHy0Khrx/
N2HZ3yNTHXQda7Smh6hPzQUnj02xlxibQhQm5w5gZnJ3S/doxUFXJYlSLpH8
nEyQobWe34YxYKFi6vJX4fOe346hYUX/QBxLmdjAFbtrk+GM6qqJCkojud1x
wRzqJ5xEu9Xo1+d9VPpAs4L3XmvaKAcyfGzq/1LCXgBV4VC39sjx8GWPqM1W
K9HFlrbgURDyP3d+/WFWUxTlmhIRh1VMW+Nc+JzKdG5e+Ob3wqko0Ha18NUZ
RNkRP1WmmPlTR+bkhzuEDD0MjkbXRyHvtHYLAcy3/hpAGUap6r9CYbq5lhuI
kSGE/XoAX9Q3Wn3xZFpNYqN/04NYZnEO5/PeTDX9laD4A7IY2DVcq0o4OTeR
b4nOtG5ESZUMj0D4I2R51mXK+a6kjsfOjySbLcExwJxXgGUKO++bXjCod91t
UBPlcRXCKz9cdZyiXqiJSgyHU3o0kYL/q3Q2T4z+IbPDBFuOAa8T5jCm8DCL
FtABiJafLPqUjs3L6zdW/klmwDIEySlt0G9SSn5nJMz96zVI4JrLTpTkkTYr
877QSr5e55nrYVeMgNlITVLvRHIbc8ze7NZGPo7myYYzpQr1NEaz1lTB+sPP
NhAnW0fiQ+vCubMU5nV+6S+uPb4sgcpxzlfdePzcR4uGTP2oCH3skoRNRU8h
r//VbC028YJWjzHfusgsxw3SN94SnzYXpvXnphz45mrNORTxgrP2Zsxev82B
TG1//Y38uW1WWbS2tZgbUuSVvmHkn+CzlMMIBxgNvuNEhC4PT7Lir/n/JKLr
i4FYjN8io1mOMR1kszXY4R4ltLEPAb0SjlZqPZDq5SHIzF0vjf6nq+XYGxmf
G0G08IkpAZqC0X36LZbSlmz/n014PVUonyUXFbwzXzmc0+Hh4WSRVFS/4hCC
WROu/oBPqhi6z5MOMPnMA/pMV3sQ8fPLtfnRv8MxuME9iW9uCXEhEpKKkcL7
QZe/zXOY2r+7gzeLdQjUpmzgL1mG73hdf+RNhnw353DTXE6MjncCmHE0mLto
i8JmvDOlndfNpuf47GKbGC/vGw6RB5/H/90p3tiyR0QC0GWpCzdaKfvwS6H6
UEdd2JiHgmSlpqtIN/HOziJIwHbHMo3YhrNUo4iennPSUtwQOq2enKWjDjNk
2X+E+2ZY4CcMDUaN9jsWfroC/ieT0JTcv3YK+iIQ/Y3pc+nX9P+yOM0sl5NS
a/pLGP8n2rHjjL/Oyjea95qvPxNlW3nIPZXOwXsC7w6nuj/eL0OXu5O/Mw8G
QT+1o/beKP5RH/4OjX3vnNjLqT5GCOXMkezcTisriwDc8oenbZTNkDQFnaWN
VkSLzbQDiUlB1zT76EWyKFQfZc41yoiz2zLne1wdZwnab7PL/QGhh96IQHA/
jLkopqAHR2/SvjnP7otdZ/Ro7GMa/+mDsndhUV53lGzAtyUJZLG+CJjjTJus
BvPZzsmsbNK6nzezCTze2dw3v+a1qNJZxQBnpskERVbeVLwHtf4OZkrmTTN2
t+5oLOEIz2e8dwAnPzTgz5WI2rBHyjdFm2HdjcZSDAx4fJe7Ryg1D1qh5QxP
gg6Dw/zlSnwk0MXsjw6OetxffGKUlI2jjuTwk9hyjZ7vPcEiScJ6veQKBBSP
y1gqQ4xqDUb4RKYaFaJ4cDr8AE30Rddr6522SJ89nM80xm64twZRKO4aOdso
QHXwcy6YRwQBk6WjDnlJsC5fdxIy72vVM4KkykJezqMvEHHyseXByhw34oy/
k1P3A+TTk6af0MemKDfw4Wl4pit5wTfydeBYUGcClRYfgXCYEEBGJCWVlGA3
FJHnoWR1BL867eX8do5GsTvC0TOWNJN938PZrvA9CaQ1xBZQooqa++HJMVyC
F9itPIPkNr3k6k+lY1lPXUgiKNPEq75gNOHUuRe1ZiFZh3+BWgFc4waMjjEj
1d6l6Cfz9nWS12RtjqGYkrEZy9Tmx60KPKyXkEXFbRkLUaGdVLTo85FL1TSS
KeFoL9fwgAjP50x5+KVxAhPIU8v583qAEUG15W+4VKrJOI6Kza9mXj+DwY35
7/Q+yRALyEFRSYozROEbPmPRTnxZCtVe69aisPNDPkQfHzXQJwat7RR4lATk
1Aj/tnt0KHnv2ki0nUGfgoVNjveMiy+SQHsG8u1Iv7Isreaz7c3v3A2dnCog
4ryAWmwdV0O7uJSaaD0+X/j9sVVOL7hSUilgSOf6MNBs/6I/3poGLbL4fe1P
Mxdlj3EIwH7J9GMdJbDIPcxegPi+bONbk0/972PhhbCbYbgL0OTKC4+jjgXX
+9IJU0U7tv/JaqIVQuHAF/CmHCs0ESeSLk/+Lg7tmEkLOI4+iXbFvqLUJWP4
bxD2ynNvA3cFSdS71Nr2P8WZ95F57GA8C5bGezlQQJC0kYW7KSlzBN4iHYVu
zIbHCOoB3jV9sCnncojJx3tvGvJtpj6Sb/Wxt75KsQSM6dTN6HWTz+GD5IF+
kFBCVyiLdxUZvOpUunqY16WQE1nCD/N9V2KPbXjIDvGDw5LyEbeoDIjkWjxL
Exvp6YfvO7pFE+gq4WYJEUGQiD20ITOg725b6iobotY0F+l7Tu8ZAKeIK1Ra
CcA4WzWJbq8EXcTwJNwci1rSG3mwtoZkR1ROTuI9bVFOANiRJthQMtduhFJ6
3qojIlKK1IwnrCFUKpbovDL9D2oiF1LNICAVzKHHX6DW29kUEvvol3z57oeS
QsDo6E6KH1UZTHv9X+UwEX83kQkEauE8cr/UwaKG3NV7EwS6whyCdx5F6LN7
tZRazY/ZehpS+2HKaUR4e17o7UZJhQ2M17Lh6MvtagJw1g1ug/qGaMPebivp
DOkaaHHev3TOQBoNqNzVZhYleTTbTAW34+y433TosHjbQytL6rWRg9H/Upid
IbXUL3EQ9nL2m1j0VgQqR+16CWxDZ3PWeyhOqqihi7Y8JNfJW4THDkL4R/e2
MDpLzl/AAiMNWacvEw/Zhx3GfZRz3KNxhd//iAp5dbcS4+rL0BEZgkC7q+bz
yi2YfD4WRDDqS1shypQVRtwLsgHt9sZuOgRM9nNcmQZ7VgHhAHptaQPQLbLO
ah/E6ZZ7NWaU/MhIOEt11DZR4XPHwNWTcZ7nTwVUOf2fCstR5BYdehe2SAf2
iVpRQjz/184QTgd3EXtES9lHlYmOhTxEakdgRakLkCme7Y2S+YVOIv7Aijpq
aT4qTclntWDsMOuVuZNRW5IzKbBi223y9DuQNatd61DcCPC/SbgTwA/1MC44
qdX4Y0xW/PzSJDFokqrujy9HvVhvJnNuPTgLo+teAsf6viFja7SdzVLQMweB
yHQs1xqpgn1ciMGsotLP/JAmC6atGn7MczncUp8Sq5fTNvHHs8ZHnjAhFwrb
Zd2E89+q6DEsZGsczybuDTCyVtGqaPWx5/EaBxj8KBT4XWOcd9y9x5pxrez3
n5BvscCkpCv5qtBM6VurrABHWWTqWlcF2u6u+JaHvRXGolGFVdMANC2juHG9
QAyur5TKUnfrs6AXNaXR1M2hjYyml08hM8SK5DjeU1vphkigfr2kc6lDZbRC
37eyitenT7gGMk4EYz9xae4Z3o2AsLyGc5Bfn8o1ZpO8VWdbThJMGnt3njm6
Ho+zdSDTaP9mgNjgW8+tCZwUbnMBvpXBB+uGMb+pHbZ/s6V3C9beqFVVYGaz
J98j72SJanZanlnEwGHDAm+HOKAG0/htO9fIfHJ0FBI3KWLfp31DiJ42ZSqG
HqQSxiwu+LqnR0pcwDzePvgFHu7XaotCjoNbFG5KGLmKL3REre1PP5KOVJBd
VMmMd71IUujXYrtzwFReIrHupjlVGDfsYfjmCzXwGSm0dP3nL3HbMg3W6Gyi
Ty/gLXHIVWmb282WW3fbruS44egwc1vORNidQdfHweTvtq1GPO+PWICCU2oJ
Gy9DlnnADMK8iqVf6fqKkxXtr6kQVDtw+HQdIhboJeLlWlVlizcOzkynLRuk
o+rVQ2YhYQC0AMqNRuVvp+HzQoFUsW/v/1MKCzXMjJi56btZDAZCNHs1T8x/
CJUY0viJd080fXHZZWO4LLaJ5/rh2XjVaZRsR41PhzhIi7uYKpgvAo+/jMrk
pxsRucviO3wyB+5UxmHaxaY7CxTmb4kj6zTIhiukBkvmCC8Eg8L7grO4gDZg
9RP6f61/Jmt5uiLNlyp5aAqldyY+ZMn+Zv/vgNGkqxn7q9auZr6icGUa4zzc
LG/FS3I6aEZN8tx0PNI9PhA0+1XN8apVc+xauqr/cmkCUQkHfwtGSG2qT2JH
U+boByQLZKFakt6gtTeCylyMEc2JzhwQ4KMlZJl3NROh49pPTcJcwLgIDuVM
aRX1tRQqTMgEIHPi7zGQz8TEsFT861KYSsMCNW0ocmUFM3ipVIS53fZl2Lv5
meWzSQ/7vzBpO4bTJpnw4+grPAv4pD5n9o5FAVEZ3wUWlQ1irtGK3wOp6NbY
PAezSrb57FhN/109fBphOmwl4fRFo69vJlXB8JgCFV5aVBQvgb5mSBYlNUBg
BKUv6C40H5V4ldtKfsaB18fxvmpStPnsrTUdNnuJXMNUnuKq2SbUYApYDoRy
H9ZHLM2ZFGL5CPTfcCcqlOVGzbgMLLoKgTO+MB03ZmFo4d6a1lSTLYQKOph2
T1tKcUc/iv31hMzHiaEe341E2MEpDvCGpE+d1AyiNOUgK92Heo8QjeLnjrBg
lqeHWNvsl9dBaPj2+Z9BqR6A8kOd5x4MT8sPKMAD/T4nzK21JmYO2sjZmDCm
mMXWA298oNxzWp98Kq6LZ5q+8jxkqnaCAKoZs5LAiHTHqxLq0qxYQky+BgtA
n/Hjdcp/qpWvzCRPJRBw26ZbeclvQChTP7vk9PIO9Yk8JqZ7eaPNW/VXeMRx
5opEtmevd98wDd8PsnylvF5SJvgdRz06UjctT67LJPn8jx51IU8ysW74VWGJ
UwB9ZCJxavywogsVe+wRuulPzH3Bz93AJ9rt8Yr6vHcl1yiavnXHmPil9qr/
T8AW5JSCvy+4iv3ydLNzRuH6B21brUXjzXqUgQ1pGPLI7iWrpKZ3fvo/XcEi
s4oeFOorx2C1tzDdX5I/dtkWyMdZXm7NYzKaenZRd9leB0PcdJvlWz/C+igW
eDnrwbQkqZLZuNu3d7wwBkEC3BPHEyRqsUDLhu6zu7GMoBvKOCWpkRNu8Xnf
7zzbxmHAoWxiLIYfx2vmliepZwgS0A+igLuVXmwE9FEYUejT1f1vDXD34yh4
kcd42fv95RXV66UGflWiwqGRIe94uVBRpxWJmmLiYo8l/fiqVEkZWTOwS+sr
uG4QLVFnZ8IU4dPgUj5/XhqA4QmC52K6RtScUZWJkXBeKjq9nuqzBjEGLPgW
2C842Utp0oc1o7+yHM3DQuX+Mt1Nzny36vFLQAf62ibLt9fdmUwL/QFqykWG
/A2IU0ZxX292sHRYZv2/tvPXNv6Rv5THA5zJvt2Iv9STYMR+zcYIxhP1azfN
OMekIhX2ssvDGFziEL+DeMB3A8rKzccPigWZbBU/XP0fSoJfhsWZXmBNWPpn
JrSxIqDwacPdpzx91ZvWUKYGGMitlxMV3heVvHAvA3/M0W/7EV1Jee8reQ/U
CGAp0680ztcZgAzFNPB9Vh5PW2K1jM3kLXk1/IGLmjmavlDETFd+JaKm+L+S
7KW56oPZ90IRoE1fBogZa+m76Hkcb0TKrLNcxWYTcD1Jlz69PpUUYNzCFKem
7sykKM1wSjUlhJl7UgWefnrx/WIC+8Qk0dIHcmNAh4Gl7FgviBi49eX7FYUm
sXIcy5fM99L4NMczqPrik3/SGHJIwvhYEWl9IxEkhXih2FPTFdncC3RAXksn
FKQ2quipfAmGxrBEKjM2SdXLTWAVnsPPwIT5FqLrppuwchHO5obVGRw5xNNl
WpJypO89LfQs0WE54XcRMDunozPuW5DZBnM8iSizkeZkZJpzyl3VbDAuAXdi
+dZ2c/81cimj7g934YbbWfJTBTnA58HMC5B1bHllCHp1C4gwgHLWucvsf5A3
HGvX9U/iDk1m3r9+Zo4flrgp+Bqz2EBhN7w2Q6DFTauGhmzjxsWPCnNK3zMB
kAFpo5VCCMdObA5FSIOZwPix9kxuJOA+wUg3i2yHkS76DgQXdUqtU1iyzwRq
zNca9cxWqFWfhhXEZoBodFrKGDoF8eqyAKJs1IpX5WPgzNxy2UKqjGEs1h16
m/hq7HAKvGqWl7IBefmhULvNSxJxEzDpu/ENaB4LtgmDvCIZcEtx0X4YMa+2
I/+SCHZHy10elziwewBz2hlvBZ+souNI/gPY+/0NDX+GZuPVh/8HVBFdORZk
YD3RvV9u44NdRemhZcbFpy6u9OhUv5xATh0r4fn7XW29TaSTvaSaPiVP9xwM
zDqj6+DbUJEZzBy24Snmd24ZlVvi5lQzJwDSKiadtmk8sr9bxe/xEuT2nM32
hD8S4cOtqIoaJu4jwnUzQkgAbpmiu7HND5R5/7KF+yHOxhlNbypxOoaHueI2
OEidQ6U0ACljA/mE14zk2O5mLrT4+FnO/vthrwaOTw1NEVLlWGMtJxn+IWVM
SP6goY3yp9noyWrLGfBeHuhZAL5LRsHj/aD9N/1RFZPDtk3BNJtT21NE9sxl
tTie4Mxwb6BcEZpOzTfgth98ZMJ5bsUCXqdp/XmzS6s5JK6HrMXk8AwRTHLH
9qvnvmrz1ovIKpYyOtuB+WSFsc+0htS8F/DKywqJNj5XwGlecAjKEeX7yNFO
HhmQNLn7TOeDLYm1Mq9FJX4eSAtEr0SjlnTylY0EytPWkll60/jZ8WE9IXn5
Vs8fru+qAYO7vglkHryrOA5wYydsEde8BukZhE7YmEWp4J8EukpnytQnA5+b
LxfCfTQOycUjMeNRa/z+eYwP+gdwixsrKWNW9LT2FaKMZyzOhw1+32sGPbre
i/CccS86YIPA6fkhxNdP1co0rnSMhEyel12NV7DR5llsJws0uIofypaFI9jQ
LUALYXYkji65YfuwgWm6W1gJAdlFxTqx44Lw3wD/s7Dcc1zIrRb3M2UUFD5/
89S0O8TEKmQu9i7r/0ZtQBQJ1mVql7Y5jtV1WUYEoZOdtYP8fMYBa/A1f2gP
osi1jmUFasaDmcf3mbhsq46QpJMos/yuSV3enBDqdjB4D7jij545UeEd6Ehg
Ni+UaXKJ4/jL8TojoCvJVHiNom5RwwFPiXAO3i/qCdphlNjqYqsvasse92sJ
a0H0k+3qIlxJvtzwlhpmiRscab8fMFFd8uqscgCQOAJqcx5lac95A8iJAx+G
5lxz6rJPvYU+klVK1qIsX6Iqb2zr3XcAYJgn25SVu2m9Iskv7Cuk16Jl9Lu8
y+TkchYY8fixWOw3u8yG02Scb0F5ZVt0z2LoVlTCZeyoeMn782yC97taKyz7
acaVBZw17lAeI66Oa6ekSSnyfugopOwczJdQlFOvHEuGT81ZJEyFYk7hul8R
958LJPai8sEnaPgTk4OTkErd+9W5L9zRkzyFQwdTXVbLzLxwJYky9H4hPRWi
jf9Q7Apf1Jxg0qh/6FUmOK/5IgzaiMvaumqB9cw1eeY5l2JcoVoV1ZTlB5ho
E830wjv01st+eAg4T6PQeotZCEZqlEJKMePvcOEOVwgBFb/NKOc8/OZ7kMyU
H6F3C24J3VRmTSx/3DBTY5rXOTku4Ww+DJT680HMb9hfDY0ojCNzWxFkI9oy
QF8d3HOL5wbIXEnXf6eKSm3QKj67EU/23zvXO8cxUQwzIWDGf3bE1oTX5rpy
K5GUOSrPX5ZuQXlb3p4mOAGBCVtP99WqX+K+xKxQH7dykb9XbRS1lHShILau
YGZPj5qc/qzuMKeLjmtXt1imx5KGUFToFwIn4BZ/JU3RnPlD3TLdHLjOBgte
ixMaonYPrd+wrTTOBKW3iJWK24E5bV/CFA2CxSQT2v9jyKpQRMek06juqg4G
wD/TnAYGRAlVyhloPDswUCUbrKp9gvtzc/APGdqcF2wr3oy3foj81xVIEbJ/
TVONgLdrsyi/Z/mMaL969R7P1a4kWyVC0psp4zZ2ipSo38yi3wwBjtlWVArr
IbQr5fX5wuDd438sUviGj42creMyn9dzE4XNxGHfvvVWCA3t6ywHAae0o9wG
Ell0LuAS4z3kPOhHAHfPHi/OCMPAIzD6ytjtM9lGl8J38VfZvO2c+ktF67ud
OAQv8t+/cJ1qSM9Io7aJXwKFXziwcWUb0WULiPZtFzZgYjO5kvjnCHZaK1OK
7GCg1wj8TrP5asewsWo0edZOdvsuQTNiHmoeSRq8+46PLWIxijhXo+k9m/js
fDbwZvpOHviQKERDwPzi4qSU4KH2L2G+fP3UEPmtbpxBHiUZjjdSG9DKG7ek
2NPGcAuPELzbpJJ+R4APFqDe2uA55XClfjmedKav2aK/bhYCYVn0Lp/6mSAo
BI71lbZDG9gwTaCGEasQREabM1hHqDjVbb8TLI/PUO9ZsShEuRkwvqgn2UrM
9j4eY+3gu4WWDS4CE35/6jKTdAHPllKAWfCHPEVryZ7hloK+7aggSkurInhr
f9Aiz/zgTHTFg7r+FjGd8LLvOn2mfjMTSAMhWLDT8FCWuPrGR1AtJx25WG9t
yT0gi2/KhC+Nj9OYB2HYrcXMV9vEjErwtIkK0pEdF/K41LL2LdOA+OQaCDkU
A9L5l8qvNThaXNbJXgzy8J9VKK7jmbw7/CTjqfuVsWD6slqwx3Kod7hmd1sh
dSVS6Gpsar1+3719I7AOw6wjuZsCKlzY15dGVMuZc9SUV1O2bm+w+jg8Xyar
Lk4gMcYB+E+6tv4D/H4eoqW2MR7DxDA1JQL7AKZLHBSIPImi++d83TM3HckF
sKMNUNrS1Kic7UNg85O45Dh1xurGRXGhJ06ZPDtpGAXp1xafEsXikVpfabje
OwXUcAiafV6+RJq4gi88kgfcidpotxfLJK0VoPoSTOmMXuRcg+IMFPgJdHn1
ToXTDCLJ6vYLde7avwUzLdfYqxZkk1Cj4gc+vNaeD6rVnhfxNoiInCO5vPVX
gUmH6XKUo/S6GVDmS+BIIdkS1eLf343/vDZgbUrB78luPQWpQ9GlVg5pXnef
As/qD/lhxzvhCddK5E8A28dnjE1NgpKPMB+ONgwdwl+1qb/6w120B5ok8d0D
iPIM0dE2qDSk3sR2GSa6fhVOcX2BiAJCet3AE1vU2rfE0NO6LvjJMiwKXj9n
mcKqWohfktJ0hcMl4Pf2XDnwWYE+k5WM3GDVB6hfEB+r7Hpt4ppXThrkPznh
C8qTiqX80WQmi/OidsyWWihRekmC3IbbAci4dui/IMj4Tx+HknU35fR2lFK1
UuJlh7D2VcKH/nmWXKbmvq4PLRET9OnT5j8FI4oKGR486yvvnsCydhtYnwvO
ohPOI9KaZP2WaD3u79kQiPk0TyrmuxAqslgio00R5b/lE09fMUMhhof2Rxv+
nLTg8KZ8JJJzGXrGCaSzjy3mFA03ICUD7T6dLOq9kSRShAYn4JJXwqI4Un/o
LX6/r+DP4/6mk3lXelOVZyfphkzMmYDXtZJCXPeFRRRrdyHIzXeTMW9MA+Wh
bNyqkJYrH4TUiOXYhEmmAdyKSf4s7zeUtE5GEHzTwF/YtY0CdO44UYQvSsUE
7g+7pjRfcP2Kt0l+k37s4OYQsjbFmgL7opsZhvFYmooekDNfQ2PcJ+ssdDho
/YRNM01i8Tya2U5v3EC6SqV9KHQe7/vJL1yaUJdtwHi+Mtg1YgfJ9s1mXAt3
zJkv8mJIBQcRyOsMJD7NjJw7mDwflQAX2JmKbiXDoT1ycbdva18JiBqNJlMc
hMZag2IzaGDaMBaOVUUeCZbwAVNOrZ8O5oT9ELS++zRek7XPAHsOPltSHhzw
RnEvN8LJvqI7Deps/MWWQ9dO30RqDH7O27O7ofp3xVIMeC4RCUn7uG8272dL
5NY2FnSd0OnYePXsIuA0i/u6O9vXOcIdyK6vQEKMilJSmZjnNRwHnbBidwJ3
hRm4LOyE/4VG4RKz83tJgsQk6iODCFBFyRzeF3NsTiwO6pzFD3FH2qBHTSIE
mOpIjqnC3ViG7uTVQGsEl+DHL11JBIsnv27TI0fRASi3WfOjDHVL+kgxrwDe
Vpw2LzkzJGIqTbgj8YRpTAwKmOTAgiwKpxdKlThT2wkYMdPKWJenyjOC5zQa
+ILEKBc7WrFLdjnv4IxFoNansLP9OeOGd3ydoXyDRlV0SwYmrFwl9caHREz4
uVjUZag15+oU21o9gXXGgUgx2vPiiUsMrUMKD1uxpaBRMuEPIgvDPbe+/h0e
NtY97GbesfiXhtCFms4ZqErPrebIpPvVdUqjDPBFRSYLgPFactE268ogIUKl
h4Z7VJ3RfZtDiOslKgF0kKQJEt5Y0/buXi4dC7CXKt+P/N7oxLIhMq/7dR3R
Wh/oBhOgAsbpfaMLeU1YrYFodEEX3e1NaSid5f3qmpD5sSYGjycf26Ta2upH
vF36O+gV1dkewTmaOJInEpHQHeKfJQ//0x9ssgVYhgTooM69hqhOnk+iaBJg
vv8EHhATHlcJj5NZVLli0N4LOD+bAJUmeHDj0qM2HIMEpA/FfLmo5EV4BbRC
n/aX+1ReZHDb9Y+Gn0hFrnIBDiqHTxzJ4xIP2ZQ7+7kVvrEuDuXC8nDGVoYr
YgPigrlwakVgLI+iucrljvxRu8aH4lqBjWmt0c1k6H6a93kERKMLwfWDK0jH
vyhRtf1hpEmGdNtXS5SQrdwqdFGaXtOqAh2vdZ6JhgbfSF0hx+eCmrIiD4o4
omqQuuVioBPKpERuvmk+kGp9eHi6Qiec6fJBv4O/YpqcMuFJ8ZVEm/CqAt3V
K21tlSJ4x15ldehokR39auXU4tOLGVz/xjIZhcOFZSu70gFxMr9TS+0khxNW
MkHdgUEANKLb+i11IumWn1lJER9LIIZ9kGeATpeH9qTwU+ZuuRUg6tJPBGHX
8g+9GRGY5OIWsA1cciQqmRf8Rg36vkdTejeDxPgtQZ2FPxxKHHQorzhvCtW0
zZljMoh/6K1vUZhDyNZxjQdsYkU4kp3BOvNRgRnON4f1eytUX8dSrmYumvV9
Cwum2a6Xp3vsWdQHnOBp3Ylsw4hhP9/T+kFFXaooJtnRF1iZjss8fuOpZK40
i2RW5EValBW3a72jma+ebEpSQpF6Sx5661gR2ATpDSNLNq/ca7yNAsgemA2z
9b/dJHXNnWyEkfibRBVxTboOPn7pBwkzZ//bg3Lcl0yvmsGdt9W96G/Fv32I
HkI8cZhEs6K+GyJ1TDkogQD+vDTipmtNccJkbyg5W+YsJuYXsuGtL3ET6sXF
UXH/psundzVPaEgI4Fn0JYuPQm3+YeKBbT9IOKAEESIqT2qzlhpvrBQEDiBw
ULHQyVidfvBXQsm9YwKNKdlBHgbSUrzJphWA2xvGHJCwvSSozi46mUipbV8R
E8tFEYmP+ALwwjdonqId5S3uN8DbQe9NtRVesjT0Rm3wYz4bbq2UrfiISAOb
CvmpM+zpaqdqa3ioSe4uh7pEiARi1TjCHHH7wR4WAKB60EqLya6v34U9q6s/
vMrpPjvTZMGrlWAm84B10cvbxkWSDpRQ/Ry7H886+VYuqqUyXfh+IrAyI6Q0
YoE9RdOoBNfC/tuKg1rt0z/w7mM6wU/UiPjSArV/rmxYY+a5OJPfFqlcOO8V
82hh2ZYsoLQyeeZsbu+kLW9+27XVBx8oxYmfLqOkzfuYYbWHZrz5AR4Vsjt9
TJK9ZvXCVPpOYDFes8tprdHDCTu962G0NtfErdb51Ns5XBjBUdjo45VFI10e
mArAjJ+GiO2JPTkmB+EZWXjgtntfVjqbqfd3//WCMpIbCGsAL/CDLolfJXrQ
s9ywpihFcz4LuzbmHeTnv3IMhnL/gcUnsmbRdJi1wi3B1XtLHNZ/gkZPriNi
hlf4qrJK4cIq1BFJyXA0lxGpKFQjQ+xkNTP8NpASL6hqVN11QRFJsyB9RZJx
fSIFJEkyUrHGsbYzc8Wh63qwE1+bqoghrFo1wOle7Sxnt0QdfYxGQaFlJDec
uvfPsgrgPMciyvJ7bCNSjtvnGRPOi1wvHO1d7moWUdx9DLp/anXwOwCMd5eT
gcxVyhB2INpZJ8kSvN4kYFC91LIjp9BzdIIZab2XKKJHPlP5XumSBChhYlXz
ZHkzVoOMtTVtqYGzhk+YEHg9F/OHMYezNS0FMDmkAIueFpzOL3LEAPTAoZ7e
e+Z/TuWiWbHMJiYurqxVce+GgsTjuneT+RSLDZANnAGgiaCiTDxbRK6G7Fwb
WMJXxVK/kiJD53nwvOF+at9Szjr8kQYK+xSzs866jY01Sa0/YPNOA8d3ph4K
hFS5pGF4BzyusddcpVkdOtHmjqKDhjp/sn0KaKknIHlLy1C9ygVXPfK/Q1bn
FoPl4zoIqYhFqb3gwbEz/EtgDy3kPk7mXYiaDT76z/oaDDFKTnSSaxB/8NjG
KSrTA5ETC2P6aTMwOLIS8F05sN3jsOZHcOa80j1i7IuaXUj9uExHwXyywXQZ
aiZ0IQZR5KZHfY7Gil5pXtRCK7yMyBqyoA/3GZGfENEKTVYPrzXqzZfZkHDg
CKt0wIGulOHNP+BPR3OTXFj9w9EtMuXEczBg890AbF54nF4DkuoVtYHWcCwl
u6AoZ1U4rbvJDXRQCaartSLca6//Jo0EIi3Urvdo10IfTDQ7uNMGd9EpfeZr
oRitn7wotP8VcxhJY0pdUvGhxeg4kA8mAGouObGk7lxFR0PH/+SqReDHaD9e
JHHJ6SYnxdSxmxvaNaI0nvCCsTKntsmODZYN0alyPZWmDoa276pR9EkBIM80
FqEHaZy1dAhwr9H9L/LsJeddwOl4T5iKbMCd+UtQZciZx4Btw6I+ywNlQGW4
ksHf7q4Zu4Zn1Cz5h2klTCZ1Sly2uL4Jnb5uRhUeaAfqXUzmMCjtZjlRbrxR
mvO0r62HdwG/jZWrACDcLF/QJH9Qe57gqYxkBX+NRUmUIAuvau1yLjoVW/Jf
nVWsMMKlPdp2zZ7uC3XeYcxISPuwep/UOwhZ2jtP0ssFfXXSy7Dd/wBC0trH
YqzsyjcvrNefadSqWuiZTIRwPdPyjebe8wfRocK02JwQkv7fwNLlGyjBWwAG
gpGdSJ6LsAE/RZ0CIo/QOJbKVgJ61Ne48fVTddFrwzzQ0MLeCryVPW+dRGwb
SLMD0XndwcGfOdWonja9efk8fNKy3aXpZXg8CQHFhImKGdbpWBpwzeoi/+tM
SAMBpHLNPVchHPHhLT82lDjmSxHP0lMmz6m/wIQExTxEtBmCBqbsisEp7AHo
krl+IcRJqg2yTf2DtTFwKFPI0QoQcMFjWZu9rWWXwhIZsKvoJQw+BFAhxhxY
4a+/u6sY7qTS6L74nLozroKqSrVSbJ2cZ0Vj4RxMtlodotBTRl3QW96hUnG6
YEhFElBLZ8O/+Nv6LGRuadvMlwNFA/iy8z0fN34S1/+QJx4pl+IRgYcQQPZO
AjfkpJg7v9ujybs4m0dEboLLgn7SFE2aFYZJbIN6BzWD7vvW1Ydu76lwcGbE
Uq6LTF1nDnfJDLok6X2AzwVETuw9UQQdEhxcAS2KsRKG8Wo7rcPo1YUHhM+q
OYmPXi8rUx6rRdIPqjw2Z84avQUZ6xvOikcz3ihOhUohY1+qBXKpiVCjH3pm
qG7+bGeIaD2+cDtuwFS1uDfXvHyFVVTZoj08QMz3Hs3Rkl8EKzGZnUTYFq0s
6ktKuEThmZ3cIwtB/BnE8uZbaELA7S671DYRrxiMxrfadh/J7CVnadx3uR5R
Vo0fj5OOhWClJOw81GXhxbkw1s8yGuEGY4vVMEbtSdYFAd8JstormMhz4Vki
vHjvNtBjzs7H5/Idh9zR+6lhiLs5vDD/F5shlsOdz9Vv0wtigGqWCfUvK0Hd
w57SA721quvyVKtVytHZy81O9LHXG047T1/MdVUG9kfLFMMoY2BKhvnOEgYq
RrUpXQx2ScFwCPP2ZhxCwmRvwLTxsB9X9YcNu6ldEn+fjIn554VW3udw6cj5
Ie1WWrHauCTARqUkMQWdUG00c0E2NKFSUMmd8jh2fifrvV9b1K1AgLRHkebl
bLmyE3MmNnhM3fheoTcXFO+OSwnkYSKB7I87os/l0dnt2XBVzLXz/6fLvD9o
6MPzruoiR6vax1ltvRBu/d4exWZ2h2dmHST7Z/Y+y1MEz67PdOD1q/BkbBKw
XktMcoUt2gxapPIhhas8Pz6MnPo23HTRYPV0UkBUhakN8gzv/OnBH5caHDc2
xNG5Y2012lzzMpFEOBXMS1sT79R+Y8AN+U2GIJxpUZgPYRoztgmwozwL8j+6
juQAICbBWR8TyPhGvnCGqQwQEBwtHOpccP+KYnqjoLtCU8uScN6HJpbcyzB8
2b30uOC6rX31lA01ILNArPpx0R89ebMB1vYcAXBFyKsZndoh8Mq5w2U2BUi0
UAz+l+5Zu5vT8OJYHGKuIovS1/PbxJ2AknFA/SXzHh8lyz5qeoOmXtECxO4b
FFdkqNQv57mOBoR3+KedJS5Q1mxMRKn9WmtvHbNmeLfyP5bIpOW501q+LfVY
ba59ymxsNWxQ9Dc6WxDS+pDNn9q/HX75Nw1sM02XtdFV9QuvxEbwnIC+d3Np
1ksfXmsP3khiajLborS1JKrWfc4oiKWScTB+aEAkV1l+ZsRFue/Omv1Grl+2
5veInZEYYZ/p1azEkdeF8roe4kGw8Ci4wFW+Wt4/KGvYqoxD7Gqn0909lcmp
Xuts8UBn0Op+hnHKHwEL2goJi5bneIkavua9imDk9OklYaNZfmZPtJQkTLSk
negy219hhvhodAwQdrwotx3aZU69pdv2nxDoaXD99EGFYmMGuQNNAu6qLSjW
u6mS0yqhJqHVb7NCXmE0T6zzhUtSBSr284U1pp4O1/2ILM+D17Su+0nSDOqN
jB9jEkORcG95usJNlYbzR+rybwobPpKEdxv7DIVn320s67h6TMRslWbG2DZe
x+2pcQbRf+4BAByb7DObrsFjyV9GSeVRZrLZhOSkBVHoPOgSboBqlA65EM12
TTNsKFfl9R0IjW5KAfYjnH4bl+ReOuhlKFl/IMnW6H3tREyXlu2xX9s182RN
6Q70XDhrE8LVWYIcpmgnH6MRXjq9MVAb+JnvLVA7DDvM9ZvshlWjeeWETqk4
/q9ib7T0rvSr8U9Wb/ubJf5qLuxTuSg22JURrIn/fWQvrBh7JBnOV1kQElXx
Y9cIwk4LRK5Lzrphi7TmqhQgYvxA1TTSDWMDtcQbHOf9SAmv+ScYSkaO2ihm
1qCRkCD1v91/GR+T5MBZIgnQrX+hARmuNauiT7jwA2U4ZkBDAgmt+XKUuTty
24oXBx4oMXJ6Qt5VIj59EdYpFwnWf03zeyBQcTfLZhqUv1RdPpCPaoUpV/Ba
r8yCHUSgp8lJZAH2pRMg7+azQLnf0rHx4mZpqH/Sphb9tlwYEaOG8lHVuK93
q6XtwytUs3+HiD61enEqLQPJlytWKuDCNk9yD9aORRm1uV+Br5vksDHfcYTR
+E1HJKeWz+8NDmvZwuWuKTbHiu9zFjHSdhdPuVfRtVujBzE25vQpDYFtEBL1
gT71aXyC4vS7PzCUfj7R4JG5UTj2shrIJDw/sH8O7Xzv2lkEl+VK1V2KJSxI
5rocMMjR6i5atDBf5dK5n6YqYraPP1oHQ0kGvIcFx8eSsn4tNZCYHlHX9R+i
EGnbYVaW3sVHiQDPk8QHfQZ42orrGqCnVkHk4H74hZaEHJBfpFVB4hnQcw0w
tK538g8RJ4rHTAYGiIk/HLftmazPsbRYr2CMdAednVi+PHh3iE6zQxpMI+nL
Cwuh+YfkGF9txMB4AWj3taWuG072vrSRE2OLwV7zqktOOP9DPSY5VNOGsY5L
UAzsT1h9OMpCICr25NidW85cBcmyxlmJysZ7sXhVcJHIYdzAVWo9PztFHXJi
zMN2yzS6B3xRZmOOpZTAkDNTt56Q6FbwjyOyRLKn8Lnxeiii4De5ihi3bRW5
yZuFbuCeRa874jY49Zd3sHiZ/M+57NeHGWG1zeDTpsfUyHvzXkV6pK1RkrNj
knxeFX7OIRNFBsY0ed52VGPGZPc44ezXbPpoirs+IK6r2jtp65hKBEHjWlVW
nCjoEDG+15wmRS4CWPkh/VZgq4pvTiWjRKMMmgpIUHNoOsAO1RVsGPy+ytxp
b9WZUplidmedQ2+1zHdcSkzlzTVcWyBVUMhJC9qPLnlJ3Dllo2/LU0Y2IBYW
SzlYVXrHlNbe0Uj3I2IDGX7Sm/SgudkHwMiCb4d7JErZTx850bpHZgM5lh+3
CthJmYw/femxrB7k/4BFKGkDSd6F1n7r7oF/Tp31ZQcyi73KKpdqLU8czZ+d
/wW4mqX5Br5EPmH4q3UYqPY6zpJ/cPIqcCyTpKRIhLXLuwhZCZIQV0XBu8LZ
kQ1DSntjYZx0zsNjXuRn0YYquA+EMqm9bvfKlEhMA6atgcj1qwQTlWRJFWeI
9G3Dfbz1YE2LBkA9ovf4aIF9PYSloKmZ1MQ4zSnG+Beer8p1LByxFKd3zdBQ
Gw3j8K0auf1kOapWo1rpdg4v8WAAv6ximka2YfON356SdbCA4pby158XY71Y
MVlQ3RonSmGQ6RRJ5FDvTb3H66765FEMzopjT84AYZAouDQwvxriCrWAY8D/
NpJN7Jm/NIsqSJGIMO/Rd01ZWtDeyZdSQY8azsd1g2eFcCQQkgB+KtlHXqo7
szhFlqw+YHOL+L8pZ9L+NFEpzRU2fw629kddviq9Deq+2SBFK5p0XoU8E3YD
eco1//YfLqNCQO1NzE6s2jDCrkQ3DP39W+CWkaZezqcJ2jnQ3u/h8IRSAPBi
T4N1EZ1xrDWpxl18062D9SS/Y87L9q8LY+V7xib2cELMKwFnIq9aJp1ok5QL
FzocZPM57pmlSlqpyHye6XU45JDeXWf2z6oH5CEUXLqs0uNdqWOFw+MZlLMi
JnrWNl1X4CMnsvhhOlavAyHquRBPxSk1al+rbrYSOphqP1fjw4bqDde5lDdf
aCKCIPZvVfi+cKjw+zdGWrkeW6Wo8uqkkzhzrzK5cTKHgMIm4dyEiAsHe4pr
uKALdihy9jBpLXJqZNq3P8PpBlCQYaPWAs92BNeOYqlawg+KyRxa91ZNFOKI
xWFqHBqL6LJwr6SLwNYwLrnyCn6ii8fLCnnZiHqPHQ0dErMDOXC+p4yazBWh
yjYZKbS4w+UVimeMiBzkfJo96WcpGzxHA4fPAo8xvxTK8aVsSX7kyA6awv+G
dRUz8wsmtXzrsT8IIEW5xvMIY2bRKL8djSy7Yxjwp+Jkdt1wfKBHQbUoHNhM
kShwKqm+FiZ/bjo0XmsXnUYNz//Q1b6cx0DMLK1FKX4tr0YA4Kw6OCke2rJG
li7iUXWp6HAehTZNmzPArJiGpMU/oKRcGxwMwD99Dpr9jOQjSxZ7AZVoeZX1
vQcrMxoKRZQvlKMYi49tpwGbqQE5OeS0uCqEcMFFIU1dNxO32acSelH2Gayg
lEdruUIaceAh92FlC7jndXLm4Rd5O/9q/GZ63mjyCm9pCYH3cXgVARDlBmJm
kzDznjMC8hHDxwQSI5j5mOinRSgbajS4DdvF/PMdebQJ/1NlASgHueoSavfF
AJlPlEq0ezc/J+nVNn0fZxM6gMe+g5RNa4D1KYjl9VzxDZzdXAoqOdJwlbSL
Wd6UbbO21lA20zNtZgn0kop1CUF+tyVPJqJbe2X8QGcYI5DyMpGWTZTYKewS
8h9Mv25uJ8Z//f/OEkUF9k6k2tKgv1hxg9kIjQ3F7MVWvg/tuPWMTx3csNdx
8lrc65kgOaTkB3ndgogLmSdtQDsse3Dn9Jz+GfaR8iwzPbborisaHtLbjEnG
fMJv2cB2otMnCkpAvChd9/e782Uft/X3Br00PEw+wfWEgqhrpAqv4UaEe37x
S8cDBzSkxvNNrFbtGx6AFfZ75mKIkhQmfU6ipa29AiXHSo3itiyISq/rfkiK
5HEhMIOjahldMNk+rRy4eqk7B54uNZwWuqs4GEEs8+Jg5vtCRoZxxnYpw0dB
oymF2Kh2aFEsOyOA5mTUhp6Ugzb7x2gI5vAelNZadTcTp+g2/+iZoo7HSRcl
Y/3HKEJ7lqBU0p7LL2QH2KhtufC2x8ASdgRqTzxFJC29ywwZhWhb8T9LNZuZ
EoWdotx+XnTMl3xMqulqn9Inlv1Lw9HHiQ2OhkE9/i8f3RmrBwtUBQxVOLY0
n32itwKh5OwfmlzPYrjDvdTsPmOm2XFVqdoYDOoaeND6SU22XIxfxxuu1csN
kPh7ShIG8jUKTBV7b+BMqlGbCmmJfn22aloKH0kNB1t9jYPaauy5MdO+Aq7M
mLdYWYhMu37NMXaPN+mbUKs8vMwA8s0pld9dfw0H/kTEI85DwhSfEazCjy5W
JWUDtlFK93JHe2xqJkt/nSVdQwGgyR0Ka/mgRWWe7fhqaA0D1XxU/oLkPYof
V9Wj7OryDJ+f+MDsvgn0E+82eHAbnlAc9wZvRBaL7amZtHUs/a3ZCompjiC9
gbCFikYG3az8UC8OiPfyYSv1VsMf94pKzM9g6ANTGMM8lSDBdTmdTgXdOTgq
VqLclutUa6PHUoz9QZMxqRLNayQUtPfqgZFa6f9fjtyZ50gG7OZ41OrmyJEs
TVQwniFdTV5P+e/sot9mv8qpW9bDfEsSpO5f71IkOruBVzQzSlbGQrNCiqrL
bQ+JYqlDjDrIh5hnsjIlLw0P/SMvAeHGS9WGCUWx3gC/BLqaFs97WE7VvRXJ
LGpagGI13Ks/ju5MzYRbdYSzAKZNpmUJ1JHpoDScS+LI2RiOMMHG6BbZX2Dm
mYu3Xxv3xp1vYv+qyFqCPTuXeO3z/vbo9AEwz3hrnXqnAUuGXJGZw5skNgo1
0c888TiLvYeyMTklh7flAuju89ze0B3D4Z1q3pgUZ4MWEPV6R5OdZnpFsPbc
7CBGkj88Y3QvLMvfLjocfwqs9T41I0NK5M9MbV6X8kk/dupIWhaDUfUorvWg
bWfu2+m1cnUfDfSd145Fn3BsnDXug/7BExOswipSS/E57sHLTKnCgtTNKlLZ
YDJk10NSNqN+HbsfXkB/QNnCS3RuLl9ZaEthXr3eEpTaZb52EjFEA02GX+3L
Rm0LjNHLL5NwrYJ52B2nQNpuOMvsaEvkTN5war3vCVtcYKy1m8UK2Da78w==

`pragma protect end_protected
