// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
1wz+EYgYPa3Fxpcj6U0UvVhNYx+EN7JS6MGKQ4MXvlMzqUXBcRhFdIAuLviNAUE9VAmnYNxjHtWZ
XGkDtWkRC9qnEvO0JI4uScIvx//plZzoShavzKO2NiZ55/lKKOfEZfNcuVdu3PjGeZF9IQsexY9m
GzshOFyCrKlLjmpzMq3t+cnqIXoINildq0WAQAC0YBXP7eDUWcl6Dp/NIXLXqmjC2+KbXb02oJeT
AdabnThd0W6UZQSzklgnGYc3rq4Qi322h0UkMheowK60DjffXzw/YIW6P3uIfzFW4Q0qaniBztR0
UrO/bOirrac6VfgnI0RhJcuqY+Q7R1Ihrz9oxA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 11120)
44p+WSnHzb3QsVhKu/ocu1UZ2Yk9hLrPvigdcOJnYB73c5WCpbEWD0X2WhRF4aKDjPSMN2EHaUVc
mW09fq/augLnljZifQoAjEpl1jrAboabkV4V1tEbPNMbXeYeKTEL1tI36VD0Rsd+KqCECejJkShn
bjAXEHs/0tbHY2CiwTIuaFc7zFlTSOCGq6bwnnfqWR43CwrDkaj4iJmFg1+qzmGg9faf7qD7b2XD
8PQFTaM0D/l2fEtsDFUV34WaFw3Oj0kdTRKsvTp/l1T+887AULbOr8QNobEoD7JyUjb74hUOtJ8J
jVuaSh03qLcSWU41tBGw0Bp3aRBgrO2YNmjItTgDJengEBc3Krj3O1wwfPt12MSYRv4fZpldVUtP
09PU7vsMYSbwAsrIpWqGXmmCNrtjrrW6/HU1OKacyW9QNzLA4m/FljnjIk/7mIMapBG0kq5A2C0a
BoNxXLzy6PZdHvIpGCOeyL4YcF4isqinR6B3CyHjLm4RVMoLOAiTcDtkxT+RaiCMQTaq3OH/pCy9
tq2TEi3pZqA+uTfewo55hnvaaIIS44VMSj8dx1akyIsTSXS50cb3h2vPW4IRvyTCyPjLcbZ/YHwe
McMBXXBuVP2zXhB5w+gUfeG1y7Bstviq9gwitcnyF30xP7AJEn5IaZNFEdYwErjbc20qW9NqY0Ot
i+KV/YKzDc7JHL3w17SsP9ahbjC0jkU7R13jMJ6A/XZkOfEhL3KUGO8h0sRBXZhj5iLL4jWq271C
iZ5WwDvbL2BElGExR4+ENhzz3Kx7z3ZEY6EtawnktWM2Pevbd/xCZCJ3UcDdj6hemmGM+L18Ja6t
Hc1xQAvQEHmtpTwpnhU0xWsHzaKWeMszgVkeW+aU4+QBcx+waRSnPnLyXmlIz98/PyJ5mBxvhryx
VHLFpB3B45MP7QIJHjp1YjcpYoAV5iR4DMsdMs6hy10uQGy4Zjb4z+d57W4vYHPAp5h0JTi1VFVI
mtpW417WRJgcBvCDm981+Iqv535aQUtBteOrFe9xzbTQ6GZljO8F3ckVkSKWmCfiRlxHRTngLfOg
YFy0TBORaqob6E+zQ9HxaD39Bp3pKM7tgalXIC3CbEmrjkNIhyXgARmwAp814fgY089lWLuDaYg5
BYEipVYj11gWGvi7KxbENkV9HHGShZzYQJlkzT06tomqkwBPQ6DkRKZiNDeT4BUb3oYiLnwsEvgD
AXxT/6FdS9b+UwtM5U6aGmcs5nnT/MW0kq8X087lxnODK5kreBKW6ECV9rqWH3E9cuQ8CxEKpbpJ
w4KaxMyM+YhNFb7y99H9dDM/E2rYYKD6b81MBavgQCVxorkkLBPkPxAZPjn+Cjn+Rhh9TzZsq4eM
1i3c+8QmOs6pcZVTEYIjVT2eLJJPIwVLRuJgjOeN3l97p0MSljzwplVtYHWcHWoPgXhTQmWs0J5X
8Z/1kUxIzeeQNeDGI+IMtj8rsVNC3HY/4Q+QX/8SacZrnDTOD3XObLnT5zKZZ6FyP+nnp5w1P9Kh
whBg8/vwcGLDMgv3uVDff5e9llZXHceo92WOqKpjf2A+c6y9GbmkqLlfGGxLfjyFVUJeaaY/xNH+
mvUt0bnE3yNtodlkhuz5mSc9KpNhh/2yWF88yOejN1Eol43x1eJrDvhnKuhMB6GKdPENVHoBe8+a
idR77yX0zUiPLA9Nxyr+UiBa8DzSi3knVjJqf2m7RBQj6XEsBeok0TZTDqUp2tvfCWYNdQR1SJ2s
cK8g16mFgv132A4aMLVo+Szc3i1J8bhmhe4bZvhrjHSVdonXL6Kp0I3+y/O6TzCuWbVtZ06dOi9d
+nQZjL8xsfKfM/Cj3Kw9TO7/bp/muP59vsSUFrASVTFRu7fiKBouhZifUU0YuuTgtFHDbFSalo3p
b9FHV3m4thJIkRq24UfSIajDojdYcQg9BKW0O2PYjNp7YWKhn573pzeQmg1/kKb8yHMC1QewaxW1
8LoQgEP+bURP8vxm6YjB0O1rxdCpxP+Mz5zinjrmraVNHvabjoA/J7CRi8YRjRdvDExGL0aO0QSn
SLz+wHyEq5DsdopyVcCPK00uENCf4t0vwS2VA5WqpRXMTkOFGOUK5tpJWGkrWkdhiyFfOIIlJva0
KH9HcycRgWV5KpNN4ZImeG2wixacfU4G5vKsWhwhy5xhd69548kyf0sMItpLbl7tGOowsIyO4MMT
qcmsPeoOm1ijWVnyc2VpdaHjjd5i2zxjP6QjsYLULVXN5BwgpqFTRLeKlTK/dNRYoQmyAfl/zBPK
oonMp8ueIGviP5KiJfMudeKHnFXojBNQJaq7B+D9m+2wqx7/kCV4iRpdRuEig487RxaOUqJO0jaG
iZ6Ob7mQKme8kCltU2i/TXmTnGoJQz026TssiOP8urCA6Gzofe4t3Ad4pF6OfJ31NErzet802GBm
nbIQKf65wpE1bO2RTkWWWSFzTVf43/NSoSflzES6Lgu5O0HZyyBtC5vJ/DJCBsN3s/RokwmJXdXu
rQ5du7yakUnvrjvFwWkMEeRmuTqCI6GfTLG6sb+sKDqoEN6ltsaIkFAZW0lnkQdQ82GHXXEzhDz7
7Ikoq9dNo3hiidDC/w+TbNQS+8f9E5neMv5t0vS+Zw+LNV1HvZdeghgVYd/Ro5SL/IwUTcMngGvY
sW/T91NWPwrDG55AGg0Putu4aAz6x7wchwnVht7U5ROlLGpXLydhi40BbAlcR9dDWOPBrYFR2ToL
Mvam3ZLlpvrzfMbeskAL5JnmP5Grb7nKyW+U5orpuSg63aeP6aG0lIvVqvFFmYiHTzHnmFc2gLXb
My/6Alju6qerjubmYECTE9H6dCX7GHwU2vZoNx42p4lsuPtGe6hExa9RQg2R3+h7/dNmebNqO7PY
swXpvv01JiDz+zUJiyYK8tkP3aaZi6HgskPiYHI4WaXLXa1fdtKmFHff7f3DTDrW6kqU0NHbc+tL
1C+ZPYW17TJ/DifQ7cYeRnWjLwInKpVjUI4mjkwm5YRkcYlm+uwzr3pbDledmOwdD5eW6A3qpaoe
DDRyYz7Xk/sFbi3pFvyHaiGgwiBysk4E5WmCIn4uR95ar6aGaazmt3l1NxxxLkoGkqvdfyKf6F7C
N6nTzZjpZAHQQjKYUJ6yJp0YobZMF7j3rhqjA9QMBgcW8jYDc8GQr+RT+bBs8McFbaK6tIezoqYY
bC53GycXOsFdrTlqBz5VZm00xFlwbMkV7P3smmXbesqLJldbbAS2SVKWdBCXwx+3sLghJiXwOcZ4
NKRIyVa1WLd+aLpssljlr+lGbKBXOW5wHYxb5H+0zJYxxEyP/fgrYMgdgYIM2slOFtg6mpKa28nE
2AjAH49GQJ4tBwlKVoL0qfww9oArC+P8CND0XmrvUtRoz3U8TRoDyzDQi0/kHNHOZpsCo6Jekaw1
WUXq1Sv7tVwFOfy7BbKjxDMaLEStr5ELZ4WWoZQkUPLpfFXdUkIRq7h12pZGsLx6dWSuBLgBBa6Y
j+VH6+YBTFfdfTc1trFDK1krbbO5I5kMKIFLWABfOioF5vLm9s1taZ4TfS4HcR/Pu34Cnkrt2M1Z
c1++jZPGsXkA8c79a9pmdXUePuUM3jY4HhgUMP2DV9bTT7JHi6wEZ+O43txoXIvRkpAMEvwlDau2
PU7T6+PW2M+PlRQpPsasLwkfyJ2G6cu44gn80UO5sWqjHsmUxHcxlEMa1GZii89xFqHvJIzLSbIa
+71tK8YzV8mUEcxe+NG6vOjbBG++2bg/ymWhDt3GZcgdK7p4a/azjsaq5PA7BJLxdDMlhWdI9X4v
WjRIgVsUVxRNwlUH/rETGDB/mXPvMs6EZWKD3D3yE881TgLyz2HQD8518vGocY7442jEa44967Lz
qJrCVyCxA1llVq+Bza1ZDjAXxxG157uTgS9iN01ZNnszUAVTHuWHInhE1Jqp+Aq8eEhJEK6wytQ/
SyJNyZ2t0B7FkTiuLggRQGaBTIm0GB9MuNFBK+mc1DwY3DQKItKyRapRU/ZJSeCQ8AIujr2UTxhp
2PmRoyPdZ234x+0xXThHM8DuFko/CZ4n9O2JbINWAJDFCnVnw0mBmmRk7Vte5D7hANV8ARJcqqym
jYt/E1lNKaHQC3RwSJZhWJ9a6qitrHyIkORfYRb3d7dcac9rFiiROmZr4+lLMfmNHuEk0ZQDtEnw
9lQHRXU0iZ0VlrUnZtKmTpQMH0Y7exiXe7+HspnvQ3gJmJiE2Vdi7oxpwkYj/sbHd3Js3YAN1uve
YsrVH7BQfoN5lowuPeX3l/x7VWdp6IL8FNUhZJPrbU2iI6Wgz2I6B1WEwlUBYTXWokDAmCfO/F7m
UaVAgY8YCUyYkoyq12cyaMmIK3lll4cE82K03+jKk7cdCJcWiZzrbQV2HFqx69q8K1WmeUAIRlf1
BQ6AbMq+2uqXyYy1PzHOCECRr+oa5lzEHSlBay8/yw0YnRlP/DWeS1JBXVPABDFJrkcQHfgGleJd
AAmEufz6XpJ0drU0R2/QyNsVkTfAiAtgwlBFoQLtssyusS01GjNduHS27TRd0bCxeFH4kl0Bc1Jc
I7lLmuqga22zcNdIo9a2eMso+ksQ7e/KUcT02t9ylR3XYvXkWtLU2RxNOSqOh/MNYge5/TWwPcNe
AvCoaTn4I3ePnyZkvNhOwPN/GInjAkgw1uucMle8fYUBDivxiYDWtYZQnjl5VC/gD53iNerK9nMJ
+UG8oC72Uihkhw4HzRswI92GXCVNK5dwwILi9mlX348RRcDn+m2yZeWZ5YzeL3+bvvURMTFWFW4S
zC5zGqcKKhXCyowzgczKaer1O+K15jSsWcxG3oiYKNEDObd1M9yaSGeHbo1/DbXCqK5LbU4YCZ6+
6S+ahMixU2j0qIz44Qtj8xbggz2N+lnWLNA8yt67WqiB9c4eMZkHGiZ2RNiVICPpP2qzRZrXc6fQ
wknwpmQQBf8WONbiXlNlYSiQdkLa2tMWqwwfIszYN4vZPVL946SjKSr7O3vDk4FiLtOiH+Au9EHP
s+8KQp2JlZTcHoTV30LVWtCnYU0La3MAPRdUQU5fRyKAg/3dkQAIXG7yXyNQ2HYbkKs9PiGG21MU
X4AuWWmiY+TWCIm0lw23zks3aGU+8JMq1jdFEN6ayEdDbjGf+eDL93KhNZLnnDrxndXH+N5OQZ/P
Q9TJWG3TMcc2iWXlMSLT489pM8lr6zwyM2N9gtInIqqOD3FjhxdWNyp/3+YMUZiUS44ltkWVF+VG
n0hhYM3vRaEV33IIMnY16vpZJIPQSHzqUczUTXHfJIDRDaUWcAoeI8yb9d/DF1cPRnT/7cgPSEqo
5mWPTWtVSWzJ12CKy3zBgMpnvQqFPf56ix+pUNt9qeAPfHXbkuID24ygs23pzENGYbI5vZVAco7b
x+Q4hvoac/Lc6Kqq7Su2Zw+hXgiZBh0fu3YjvCr0/MTtXit1fAU7NmQDzEhHcwMz3k4dnENk2JKK
enwxTBxAZLqL2mJznEE50J4yk4Auzra7iMfi5agVZAvHUg7/fYMsj23NAz8MLE583eZuMjNTbgsq
c0mC7qEdxlDMY0g6Y1dZ1sFMXRY6QQeMc2LodWQufwwuBlGt4XvJE6l1AqFJKLeD0FE6m0k2pE+S
71Dv7ywInbmAQxbs4LSuSMSlEQ0Qef5xBpTnpPCw9oZbbVihn+9s3OrTPuG3vZtT6BgRbz61hvZy
kPLHq0d8LxWrnDL8hCEug00N4LyILRVHII1G4ngF3Q+9fX3OFbOO67MLiemdohVvcXhN/8MzenrF
bjlw6Q51nMrrrWy7M5gaQd2iyDF9M/5mxgJUnGVGaj0SWMvHXJlG9/LQS3MnFeatfzN0q1+MrLbx
fj/g9vsdbjXMXcJ8bQtSFdm993QY0sVxJWloXpUohVL2gxMoHq3YKallcEMVeR5ZOdv8WMIur3Yi
5wrOuiPg2ybCXLh7aBIpuxQTktdPou6JDEJkHJFnHzgBV6ks0vMuQaTslStnNOqF55mwzAsjFC78
J31F5i/AgANccrArMLe+wJlkDMU2BIE7czZCiVcJGCAbrTqY+x/qgiB8T3PXYBjpDPxB9za9DK8u
toEOKu0dArjmCZkqji+HySGNd5ilgAywAPEsgYEpqV9nWZCMD7vYPXTvP3zrTLjAswyJDtwiV8eL
BH//h04TaeXCyatfYmQq32XWNEozshpeoeToVmfSkIlH4xCzytWPnVWtPpyU6CTQI1G5Yp9unGNn
ypjK/PfwOmNSfIJZ0xPnDrsGWIt+5j7oQjQU6CU6DrYknjS+/OPl/3kznbjnMePrWr5zh7oAXbgF
5mAJFTqjhzHQq6902y48jZCAGyfkX/UkJjqqQjHRPS8Lg36UFXd4uG9VNhIXSgNYPPcFG+x/weJP
c+3AtWGgee8Y09zahKSm1I1E0ml7OUtT2I3050s58qXLpPGYQVRnxazedSYclA+/gt+hgrBx/IUh
FjNWyAPsuqGm38dMFN2n4Yoio9VUj7qTfk0mpdoeSt0O1Q660E+iojC8iwT86/QUQPE2Vx9CPYtt
XXWjahFoRCZEi63SsJwE7t+X+9ODbUd4Z9HdW+VHIqKJfLNEWwM4lmggxZypjO514OuKlH9Uy1bZ
eEmE3e2WpYzU4hYYNqhNABoqiMwbwKhrRzhGW4NB9obnF7ZwfDY1ZSYGqfq5rIJUJmBulwg43NIT
D+vjvRUf24VPznLa1jH5qT9AME1jl8uTz+EEJSOvS6aZGjIS31kipJiLwVRt28jQz6ooZqStzno+
4jDXMEY9fwH55+tgMOSIvZPmbLUSUIWzB6PoVSg/+QzK2zx1GWJnKe+0M+d2VosL3rAteYsR6kxt
k8GguYoREIuC8OQToP2GnEHdYlhGTQIgX0mp40hDN6gA3Ts0pZEcwzjwf70JcY6QFpDPQGj1HRwy
YRiReG3CggwtVwzRxx281F0iymR7L2zuf8O4HdKot/b4FglETZT1Ek//s1KQEp17FeXEMUrU2mlh
2i+aJQUYJWtjqrGsubOTZW9p0aoMscgBj/fJjo4iMdKU3ua10PYstPhjHox1UQlyEaEE0/cHc1Sk
Kvu7VZ7EyiTZX5xBlyMvkLh1s5CFES8+ZQUPUQQ450w9Ot2L3ECEJK4NVqHSzaYF2B0EOrtV2wBu
g8muOFy5K0vkWST3N+qU9afk2+JLbnQZ2gK5RbUbv04FxDahl6HUg6rj98Z6MIzB0v9tKSVE0twN
Ob1HibG/dUV7M6PH9Y1H8XEUYRw3EYbzEpv4tFPObunUc2YgZUR/SqVgm90aJd9upvG6PwnHWeUj
HPexmBuURd/sxw5FrXZ7kBOET/Emp9TyvEm9qSZdg49E7Wn1L8yZmM3B0yBtVJ66QqnglBrbjkuR
6Uv1X3K5hiNbdRoVekbw0ciBipCwMPNyxObsQ5zNce77exuAU8PP1lCT/vlOKZcgUNOgKVoZHwVo
WxVIyaC48AHd6yhGsEu9ERM1itbvKBJKKhWlH62OuM72s9ivEPvi3Z5k7c5y4BnAR/Jle54Ct8pg
ElNY7qBwDTmBmXqnOt6l9qFkIF19Dd5iduo+KJ0EDaWGhdYkb94wqrEMe3IiQAlZD1Fitnv94XB5
Rq6GWwMvyIqv0oOcziu/ZN0EFNa8n3tnk/gGtyUSaNvcKrpXt7Df5sASOg5w9luq7X/2Hq+6CqUq
z+Td4wgPsLeAXueqfR5whfQhFEFSuFGkSW9rMeRkoyrxQ4c4vkH4ssyisds/5TuT+Tc6+uStHhBt
K+Xm6+7PmCRssU3iEwAaF/879IXz5/Topzw271rDSFAyBIms+jJ9QWq8nnSafRne9hLX6tdiBPbu
1f9uwnNNPjRF4Kg+ncTN+CKKjIUJlnSCE3IOxVw4AtBUE/E4DMAwOtdMByaD8GL8p3jS2lMfb3VQ
HYfsJRN61AwF08go7WLY10TWe73Bc819QVrAmI4Qt5H6RUjL4JAL1/6xBca+b8D5qX5qc/GDqkrH
N5Grd90Nimp/xr9h9VUyohSrLbrquiYjzZkTtXIVUaEactVDGAuQWbTZXjQLys2VcFqqYLdo/APO
6+zF5tEhuDNKUAV9+yVemcFNrKomduTSzO7jOp/hiSv0GGMiPvAw1ncPqEva++XI3JXt7t0T/EsI
dzfZ6Ws388PIh+SbDcvcZdRmHUU1Ugt9U05C45empsUFbb0EmQGQZxzqoDB1ar4a7rGq+cBtqok9
AVgT4FUCxpTxhnq/qPX1+w1yl8OVpqWhHD4GTlPSrQ3iybf9FIydstIGKNBI+IDe0QB7B0chdwUR
RJNiEOyLq4cm0R4l2gnQqTqr3Ant8y3pUP5iWw+N4rLP/3USgX1SSPJYP4TECqimXFLrMvGOBhDz
MFNTnyYch/liVi8+dk1suiE4LJX1dFWdMkfFtk9qCXAIGt8e/WWKCeuFsFoq6kmz38kvr0+HkiY7
CK5KZgfOiu0I/nX99L0fiJEdR5s/JRrCpDcUCtilUrXZwaOb8p4gvXNlBcPn/DBtVeY2eM3pa7vI
6aOJHwSSHNVhs3TOIdiiPFPdbkdanABHovqzHYggmJHMUhk+6BKRBx8o5w7Jbbk805dg5ydlvfRq
EpO6d80ma5c0hZU+h/a5VhYaGlrYm3ZhWOj9KLMdzNyd0lzON9n4CbpSsaOIKzSc3CfHBrjAcGsZ
/FIjcZ1U5CUlHw3AFigzVvyfjkWAsmiNnr8nNyYyVdCV1V5FMr2XW0rnBnXgoC+VxkvPFAZrrNzu
L1NRsKy1fkL1fTbPYNDno4yO49uXIVKG4UkJlRtCoSWyqj8Du4bqbE4EkNlur2GZ4HgQdwhQmVqB
k8PcMOaDFDT/xhoNvEKtVRe9pBaR7zmiT4tKasVuRo/Usis3cas14CX2EDOQYOznZ3lQGKxMH+St
v0uCjt+nXO+Mv6wC4x24IooZM6aRdIi2EHskaRVgwdZIfJppTcEb3gpsm45ENOiizusmOP8TXHki
bOpr6K2XZKBo81qyHwFJwbXsCSIiLdvJBH7B424FwIayJ3Ny+i4thLKIV2vF9KPAARFgwCXjwO4r
/TVVquZoDjYetaQ6ZR7mBWOWioNkHTJYVPfbcyI8+ZlFlmSKgugS5GHTsxzDEn1QO8W8br522MSD
b9ROgclmGuj4jZZEAdIeacRTPUgduL0PpwnYFTo4qWGCg/HX/hnuhteI+MvtrGWA+zU8jET2rc1P
QheDfzgA+9CKpdviDgrMEFicERRHb8VTMT3h+sza67chgcI2xn5EuAoe+9Mwd7VIYi4uBzvGz7zP
Bs8JNN7qdI5aSmIdMcVp6AaFggbxV5RBcnYm7sPR5ciWNsohnVDeLwxV7KEIrd3LsF3QkbG/6B0w
/LqDMKrEnCM9N6xUYPTh6liCgbbh1Ebe8ZrcsmLXxKbkxt03wqDEcL3+Xg0z9oKTos0wycaIwdM9
i6lUJGA6Y1uzM302Rt5gF2nJP88kIX3vZ/011Zx7HEpwPKeltsWJN4go8iP7tmeXtGEodISE9wRK
5HEsx405zwjejF2PW9ZCfALahhNr++EwsdzcHPzYfE5ewi6hcKZYUYMYZuJ5IasTDBB3ZxvWEZ/s
uDVR81MstanJSHOEz8jFevMDSnAbCZefGoV6/CWRLG0JmXN5OZr1PTlmyoquJ9IRFhYX3K80nGaY
CuMNX13gehGEcVKmBzloPw9bpRQoEIUwLwC2eRIQGMcLoAfqFI8Jnyd2HL5TnTzCbT3Dw8cKs6+1
/rRn9cHO7n4ZtSPj0GQOO3pnyyY9Rs4Y5i3B45jxdfRSovslcq08HaDbjUyKCADov0vjmEMwy5LM
W0RlvZqnHxUZTB45+O3DNseDXxRcp5ghA8jZirRLxEp3WL4zp8wOpz2Ay5YE9Eel/V2gykM2xiGQ
sHe4/Kmr8y6FwFCAzLis7cAY71FbQM30M8ftF2+PvhQ1VLRZZ0XiYgHPFQplbsJ8YjQ0jgRgycYn
9+PS4fqqGFrvOFq/bWTPM49lLG+fZNfTrmSsnnpRcpk30VVjOiwAhun4kv7JKirs4o/gIAAcHcvZ
pm731bmogfoseX5rB2ikROjA5zv1RY7Tia6e4Yz0jbATNUxB9WXzRwH7uijnsFtqUsClqtu7AQDW
7Ma+Snw2MsNLXERBVJbqeKZIwGMtj70va9WirwFolb4OouFgZn/KAlggZ5/XS1vD6slzkhEyQwne
/6yNwmY1nC9ciQH6fA48/WCikOj0Bq8ogvXMVeHV9560wgLRH3rYDbJGnNODbWS023LXCDh4/X51
qXJsDBQ0uFmm8WlETOVUK0plBfFc4LM9jb5CERBqBB4C6fn37zC9zR+CK/mG4Z7zkGQQNEYamUIZ
6PT3AIkaa0soaoWXhCB2pWENrAL3604QMLGUw/O6yuF+py7tFMlZs7J339bEHjZ+z8Jgacejg4ih
QJLjnxc+OsDee/uQfelQdsJkHFB8O8myqCdyqPvtoh+x/rirZQFfT4NUvTeG8U/BVD5idMauvF0b
ctyA5XGdBHBRBcUimaRYqM1Sn8d7fklOsMiA+dIuP5vPDL1xZ3vAzvXrIfwIBrkdZXKY4ndxgafY
eyEH22tpBOAm8BtPbcnkL0M79r0GPfqIKkjZzXjfvqf5kvaEcMo4LBlIDcnpFEjSq19op64mfqRE
BENLrGWUaLVgn7zFOl89zUrVi/0cvYpWuSDolAbNPyEeOp20tv9mAxICVLuVxYujNLN3NVL/bSls
oEB/YDuHvoUiB36jI20+UTyurrhvwlKuO42S4ZEAfBWX2975ZJw2P2M1aUUCGW+KUTYdqD3kuUlD
kY4f6AXNbusZM/gYGBHjoBk8aOKJ6ElvNWqbAfwJqSc5ODxA1Hb3jXQ0w+8KvgYWSHBx/VU6n34v
pLE/BhPH339KYlXwjLY/+y1BPy+FTDXRWrqN6DrLhmtEcf6nNlIAN8blRS7qG52oBK3rFH9dG97h
es+Faycn02XYU8KKaF2iHEtKYYcmkKALrzQahHawgMK1vNK473YsYQTJeHhUxb9qc4isL3eZP5tQ
N0NSWPv8uM0Ix7KLEBlaprZVJsQ6+wbs3rFtU78T75vHzzmsGcwX2fLfSz2TnFEyR4gKlh93MJOI
zDWSwTV2M463XnKqfezzNEyxTCrlhUpGjlbWRpdoC3okf+jw4ZFazxWXCmruB2s57MPMHw/r5ALS
CUpK5STdFrd1NfU+n73vvzp6PAtAIiF6qpbHAwFCwBCrT12DrDITgDmQJ7QC8xxM34hYkftnY5St
iHwfHADur8KbzvtPcEJ7yRRq5jKCTxFDReLPyZKEmfa8x4u0p6ouND6F+18y6cM8Ko0lThqAuhZI
ApmpvSaGXtGxwRO4XBPlNkafiAjc26KA7R4D0dAjdwV2gm3MlL6yLsSg/ZbJtQduay0sFg80muz7
F6rf5+cyl6LvIMC+y1coZcP1b0IjwqEHNkb+FZlcH7z2/KVl9GsubtPBkRDEMhCAi63L0cdIPoXI
9Sl304LhVP8Q9gt57cKL1C2OIUxZxOfDrM79I9Ptz3ZftLNS2S/gbprxpA+FultNH3JrPxSHJusS
3Vtj2QBUuCfuLhG/e3BAmbxnVSgI/7po2tRCcgVRivr7TV4JkQ4FsEs2nTDnKZPsbM8Ea1Ua2rYF
LrR50KubRf7ZmZhB9gTXwqTrPeMNYAlcvrotzlm48zqMD74e8d2IhEnj6uCx+FTq+cFhYclQJj9J
8XfgvGiSnn6L1/y4h6M1Rcfobjgcd9cWjDeHioZ0BMe2FpEaCEGC0VxdUfvGFpiyidvSJKsyNAIB
EawT4EahpWLWjn7FhaoMvqOM4NuVvaliMn/lzoZxKzCi98JzbWkUoH0qotw30bxFA96n8eixCB57
DqGM2heiV3X4gPE0l9ZClksEOQuCN/lrhYkN1B1rU6f3YEdsCoF/HNolMkftEH10jpTvTIshl4q+
BvZLaSJfj6cMLgDz702Hq5jlpJdSjurk9on+kJpYtVThUT1uKq7JFeTySPRKUJqY/rQTo3c/XJ55
WCwKArAEqWtb+6l8tzTtITMb5yfxTKZuXhF3K7CiCtqMVZ3H2QuN2pUtqEp+HY6jYotW8CSW3lEy
xPdmNNjCb49WLOknAt2TTncitPEtvnLy1KACfA1YPC0XUW08PL3YWiGZO1WKgKgoTfHavcJDpm7+
rSITvCBN+y3hUe/HwioVnmHZwS/5letIOTxWSujKhmA4fbKhVaNS860R6vpko6eTjfItU/X61dBe
rH1TxZ61vxMrBdzpvbRNZZ8fqJxDMDMPFyWsX4N8Tr1rTDvVDkwnOxz8WXFdGsk/QRZaQJgJvXtE
nshsABrue53TWlhqTC9L8LB6tN9JQmg4JrdeJ4Y+/Sw06AEdNhG7hzspQJwZSNX1qozpte6CRQvW
e7ESfJtYCoA9z9q34izyNSDDLzGVjVYdyFq2PbvzePypnj440NjEkGCIIL6ZW7rFhB16Focuxdt9
1OIsbcZSEwnLts0M3/nXm5SIphUXsE/DuVgJni9R1OJ8pcjHPNM//CCHe0TC6pnyjoxWHV49leqW
9NHTJaX1wxHha7NS2rhkFBc/LfDdK4iLog5nBYNbvNCPW/UlIAFzsFaNpUWaYVrLoAaivKNTqTXa
M1THvf2O50jiS+zG8PemRDAHBLjdu7u9TMnlE8y054za8t+07CIoUMkNbF/uLb0ZTgu3IPxo0WB5
pFRziNeoOIL/ILE+1+7b+FMtZ90GxcHkKdRb4EcGBBRWKWRT2w/fbWyCvs92UyPZu2ZTQCyx82CS
0SdV6PXdhbMK5sFR6VfUS8mdOBbbPedm3JdWNj5Bgd2ecT2g0cVqoFLu2uROxIfpiUb93KVFy3lW
jRAOlELG9XrF1oMMQ4JZTRMnlAKoGyGfy1V+pWEXtzXCIBGPxmd6dzYNt4oUxjW5mturkf2qXf3u
kINRwPqtlea9slLlPULjRX7bePjFECR0pAa6CLr3UXFFGJWtuSypQXG4iuLOOKZVQwzHClOrHQH+
EPDHypIB2MqJ8/K5NK1msKiSTm9W04QneGYjo+VB2zBP+SNx2KfwarLcyQ8N6FL9IO3N7XdJxU3Q
/3fSZAb6ZbjPeq/nNDS9Pe+b9qoZa6Zr0FJVnlRDvkvTBZWV030o2PvzxWwqpR9uqws6qKTgf91t
G4LwopjFwuAsRoB49dlGKreq+ceHW4SsL09XtQRtWIJeJJXu3Ce+HK9a63XWIdaMA3cmt/z4iWqG
qsF+S5eS3VD5tIWwrulPBIym6lJN9YUL3xz6ssNQn0bJ91NcY6fhucrjoDsMx/UvtNgCExux9daX
GRe3dXQ0uIF/7pvX8r0jR6VcIAEUwKDe+Wss8+ra5LyHvnmt/eK8aX3nJtXriqLASQrYwgVtrgdE
yQRuqby3BkAGfu78E8LVVDu0Zoaj/poth3WcBM5WYIDIibjo76rUB/Y/zfNsIju6s7Ixc8aOC6cJ
ZLvBBvxz2KownmeNNe+PLTOJmmEcExT5BdVEIQ4xOKOZeVVfRYT9aJxstHmH3wUneBxyCeLFEm7H
sPQitEpzrTD4oFbBZGJK/u9tVmbKk1qkYMaJsoVXL12Iq6F2nWQVsoFKC2QGUZG33lBsujYYAVbE
mb67uGRs84Uara06Mf3o+HXXsb15ig+ZQ1tmNCvgvKsObvwR5BHVZvr/nbl1n8xEVWgvuDmPvmGQ
ah/lyaWCORc9ekjgtiHMK/rMcSJFIvlUQalIuZ5ea4jZ2UNxbjKmZNO6JT6nEdTczM3IYMp6d+9f
yMs8xTKNIA7vXguSTMDqPHtVcA+h9RlBJ22ls58g1KX2+zuhYTY/tAEqrwsi5o0e4Y8iGWKhhZKT
FdHSCuLbjMNYezGcs0w1RnUwtBEoTi5D4eq92eDpqVpGOWvpLG6sjE30e5y8T/399UybRdXVdT/8
q/MzDC1W5cG34H9m/OhOBdjFalYNYTQQUeFpgTx5zgPGtfDEqoBu00G5MM9+pytd5Pcj0m7HIEOZ
iBmGZsKjSEAx2TwqheLtTNzLnHdOI0IHuFwUmxH3zAY5/CrE8Xg9+IYdBaULLEyiIJIr3J0NDgjR
FAdLMS2eYoaJCPK2bQIPx3W0W6KxFsY81hhxMjXt+h5mlnsGwlYpARIjSPBHwyzClVqeryuJZYy2
N7vol/YFynFfPSx7WihUpZC4WJXlAQ7T9z9hiqA18gZKIMuOvj5n36lhRI7eZM/DilJRyM/QpwE7
h9RWg7/4BbXfQ7EDAMBRicaOdakyxUhp/wwBjwxq/rA57B8Sb6aBZ7zClyFMnibgoCs2+z1pAPBM
UsRkeSabrkTPyNHLAlGnIULwEZnzDz17YaetF84Xtqd1M5dWapSQNs9zbLW32BnVKPKBesrEuVa1
JehogujfiGRhFvDGyL0TlIGjbwSEaaDlu1cskwMC0y+kA7cz9StSp7zXgoCpzwehj+WUiTaCagFy
BDPTtqlYAv7HteyQjL6784mS/jB5JL17FBnAyIz2keLUGcpXEkGHt09jieV/hfRpRyG9VCsHOrCp
RQv3ioYYlmxJ75q4s3MIuo5bo8LYpNDJSkweZRqybvuXROM/1lWPWVvmZ9rGe19mZmFFYDTMM8dJ
SuhRplRMdAmJMmE3uaZWR/nwK0/wO1Di38gJzVX2704lzlYvPnnQwHbUwT+jE2ExQVI4oG8lBR3/
SW1bMCmbuFh3PdhmYFPChVcisW3TX14q/j+uDRdC+/hrbzkfJiyk/UY3pb8CEJgGGzddgVWBdaBT
ubhkUcHUW8S0Z4oZ103KQBqnqeNgsWGOf2/2NBGrEUV4slvdO1EmVgF1qNuNBOqZO2tE2jSVJAYY
z9Xwsts=
`pragma protect end_protected
