`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
eSwsFA+ELS4xIZGdQ9QGimY+OxwJIP/LkfVXlrImmHGmJFPx5t8mTxNur4eLihm9
TBLELzrceHT6W/Id6F40HrjeUi03OKwLk89+PZrgFSFvdWgdDvEKY49AG/mDb+7h
tdLJBDk6Dv4rLiFcF9Trgw+qBK2vjYtEEqLe6M6GRR0=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 6768), data_block
RdbSqNVLeu/DldWA0DMbQuxveqE2g0CE4sKCZolXxIDaq1WwSTi+Q1I2NrTzAQtJ
OzCAPpbIOhMSq0oarfJ/3GYblZHfxaWdndThAlzzgi33wXKS5dA+cpcTE55p+jo6
TZGzexn8tDzCUunc4VelyMzG4enlKwyMPX9FS/s3236Vs8fuivtKyHHMHv+FE45/
WP9NHcRVwzJvlGRkifFjjygT9mby35FQYiTHsUEKuJyNZ5kQ+uAQbxWKt/UC6D3q
OkAwsdfnBETiWYHq/NYHKFeZPDyYYxP35t2fxWENc3W8Hzj/xKRjWe74va5F62dp
kZI3woSwJt21pKx6tOjxWytRDqAdUHiGOFRVgnDOLs3mtDj8Mh+IT+dfe5HVOfVZ
bnlkPQkMqqNrIpPJFl3MEUqjNWvPeJlQR9hm3SCjMeYKZfy5vtc7+t7Xaddwecu8
Z6OX+PMB3/h6z6stRX6hSWn4U3p+HGbIJ0DxgtUlBQcP4nlkfL9tLHrbIfnq9zXw
S7fxcIpg8/BpG0Dt2T5Xpdc9ln+B4kpbqhdJBjqmOt8hwzbOB6sPD1y6/qGhT7/J
+CIV5k041bCbBW4EX4fc8LYd3K0s3442LX+M+wsyvz7rd6kTDDUUnaO5pzzwBCPI
1D1p3/xlzVgfviFK85hxGQql5K8iqfS72kG5tTWjgrNJC0ggNk/OThAxKJebBG0j
0b5HaiOi5EHq1lAILMPJXzvMpI/PwPc2kwtOEbkNA+4b+DjQEiMSlLynbcajy+sS
IxpnpfY5zuZMZG2GInaE2ibB2xvBZGTcj4t9GThQKldyuEw+TSvcS5KhUn+Znabg
3mEDcWAOzU5E1UxcUlfmlpy6JnsxRAXRevP/vIJffTtTHMSXp9yrHZd92b2xnUlw
4++Ksnk209VpIkPeeXNxbivKpcKYge055tzmTK3rnr+RBjMBq+4exKE52E6B3LYA
qIwr81fw2NECLhvTm64lb9kEHK5D1k0PBKIGRcDZjXu5wTMi7GugdKjp8/dZZAYi
Lx6lIUjK+ETt+jSQ61F4AgaxBUtC/2EuSU1ADVMSbDbe9OcTyNcyttDgJHUWwssX
GIxQQNlWS/wOPXlUmm+WTMnDnAudmpTL1IWYI1hR8pN4BwIy9riivzEpP0H91A2W
lWM0FSySo0+dXnK1q0yq4iM1qBupzGp0fak3URVRv24lH2hK/RBwKlLPXOWuVpfl
er1Gxm8NkEtcxQ9+Wnr8xksrfT+6Sh9Jqr8gEmJ3Ps2oyIrdBPAZ/zr0NlB7ceZO
8lNZatWDqhYIh8aK0YUl41N84Pbb+KABipw/eP7xfn0oEqkN4NlOn/vxi7qERPZl
WidN+9BI8UylUs58NSzKKnQKBhydqDz6F2zwe87FgKmOPOVCBJJZ9n22v4a9DWm4
W9+YxFvj39rgxKit6xXbvhwmWbxJ9Fjyn9V726/boXEDwrbKctAo5mWdfxwZHPaa
XeCkUTI/E8m6Yfd2Af7yRTnumcUdY8gLzRx/v0yZLSfSw8mw98F4VYb25gXjdONo
futstMZQsnHiDF6ZHeJSdYyCqAD8Hffvkv829aShhTgoZ8jHklwJZAsASBX8mjhl
JTK7s7uzNnanjz8sav+MGaMxxVtzh/Dkx9GjeZQuhG5ikS30q+RKP2NMeUCjgUFe
eyxn+oVkMtth0BiiZvCHrwY/OHCaqUQfKdd+6PF8LimpE2Id24121UUoBIIF2Bff
ReGBf+RWVVayZRruS1VrpysgIgaUXRzGBDqhwkqPi6wmF+7/Rs2+0s6JN+rBtcCr
gOaxFP4DxT0tNGqHJyqKOMGlgpVlJxU+0LH1sRnSPWyw3nNsZQLNUZFtJViWzW8a
FOh35eXW0xlccoowXQMoCQiwOZqp681lJDwQHeHu+uMcHCjSZyS1AXaZvk5grCCo
VUFxnqeLoweQpY+qs6//7GRE90V4qjEzqeZOr4yRpTAiMw7uk89XQ1kcBbzg0ipb
v9Gapr+LGdHm30g1AnwsIUKwdB6XTU4TKGU3S2KTqon5eKh71RoKg1xOCs3R1qqG
xzkLuYiLTYtcR8Er1JkLIe0/ir5ui1u73s+3d6tP9zsqpDmLL2MzqrvzSrrYfSeR
If/6/P2zOT1R9FKq+L9q3T2rmNPxmZ+ZTJawi7WoNTxWrb4le+m6eGvE5NKJgNPX
Bpbv2Rm2GI0bonI442XKWm5iuSssA5x+KaxHaB4TGe/g2IldIryt/X97meZAF5xJ
QNLi3KIsrI3pvbi52UAT74sYCd9fWK/QsAB6bHatC1y7XZLv9CzfXfVoXrsoVtXD
+o3fww534QadbBq+4bZeeRQ0pXBXPrWAziD7MrPLpVJLzAFH27mnYbEU8N9vdh76
kpeXEp3TV20M4mZOwTKWSYXUSnNTnzOFbvuahyGKKKCEn+PxhSKjPUv9g0L2TVzI
+lDz0Bebl/a7SDVBE5j7FbUA2AR/JZSkl1xgsKwXIK4+Pw45Lsh7HKx2kZQhgPQW
oGdA9nnpUZ1sn1tUMfKPeuT8M7ZoCpxDMR8p6K8j9+PLNJBleRHBkxdH5nmht2oc
5ATo5Ywt26r7bHQZRUoTSoGQXYVAZgBmhfVqVJ02Tl8ZuSTwHT8OrgAVSVKmv9dj
+IMCUTZ/c5NgmzocComI+mSoi7ePx9WRIfFDX0Tg6w5E7AL60RVupedF86NeqXVg
FYQ5vfq5sgG4cql4huFVcxzWA8+a/3+g8ZMpF0kRr36he4dsG0vZ4nJVC3WeTluE
m12WFVHZ4bl6d9c2V3YfAvdxatPM4hTBgAw2+bkHYRFfioBeMOpG8cOgowXTMb+I
P5vj22AGKe6RDFsED7U8jTikcFR2t3abfAuNzyBCVcE3mWyeshC25jrZqr1JUM+7
A9AxH64S29AgTAaV99Mz1pJApHkTjdJQ2boFwrVK0J3lUwJZ0yeJvb4ooJVuvfRn
P0njsTMla584qgdzfeYtpthx8jsenZ6vdHwI6wMiyMoo7Z9KRdflnkpE0h4Ui7C9
rWhsjfMc4rZxx6aNtUmXSqztrkxL5EuazJW2xHUnOYRe8VO5UbZ5YR60JxmmLHeC
PkVL6+f8+ABZmqq2P0odn/3m0YXVZzk3YFQy3AdWQuM69tew+g4vwWviNDCfnDaV
afKLKNE6ShgN5gqnJQ83l+0tE1y7HWrtOeIw9IezpukpxJHLwzresTQcxMpH5BZD
naj7qvp7+okfdyRUZ1K9zd6aq+QWwQrIz/BkkUAoYGd/qSerirKED5kvEPUqp7jK
6GLlsaaV/hdqhbJ22Bm4PEG3YyhIjQNsDEVlp0zZOKjfYIwwF04z5MPVwtZw6YCY
4s9H7lOiMu86shsxqQTKwJT9W3jiw0TB4DGs4LKNY/oaH6fZJPqBPey9YO9Bu/Ox
+hhNmFumYH9NMIvYEwA8uqZHV2D2PHx3GC4L3zlaDPEslimQ+qPkxSgaXAa6j+6Z
VAb0kQYmJNd7V4ImrXzww1Jyh+C6HC5a4beY/HtFckJEPRY6ntxvLovR8zuTJ0G/
AzvnVUmnbTXN6vk+hiQIdX/kSRvbJDhzAchosj3yhrWJK4lAAOYQj3kgNQSr6MZC
qVrMFtFzUzBSkO48kG5+i/FLLuDMcaHsQ82nIq5CQ77oIdPLfzKk2zVOqk/7TX8C
V11XeOOc92hbmq7aMts7kfDplKvza2uZp90N02HXdGFFqN/Rc1o/HlKsgWsyHLPc
6JPRhGePLwcHBr61n76UPWzuA9bEF5uod+9MRl43gaQm6x63Md6hFsUextNt7+pD
S2XDdj9D8QDrcVNvSAB5MX8jDxkbSNidVTWrMn/jFwLt+MsAWKr9QesEygWI/jHh
X7tqzhzicO8x/y4hD9EfYxBODuDL4lIvh0d2xRtjhpql/3kJZ9PIzCKwepaA5iqy
v/ukhgVkOWWfH4W3sabdZTno2/IRXTWCGwFn/SghPSaW4etXeihjcQB9B5E7m4LB
ZcFUJRr5DL5BcquSpi7w5FUEDQgctJvw+Esq89IJ2+A3wlOozgD5/mcMtQahbUvF
HFG/MBZ6/9qY1diZvwEZtvtzxrM2pEFdvRdaXMj8OdVsnYYOdJp0eTD9SAcFxsn7
l/9eGHyp9fInwiOuGnPPEVuBvknJoBV6QVdFWys/Mmlw7MoIrNh9j+qoTjWMH8gG
BuvEWE4Z5T0o0sv8MrDEhvhHapvE7JH+Xoy+RHFBzG32M8KKkRHbo2htFx7Kt4zv
m4EgbWpmdRHsuYMFnGVAMv9FjPh7MYMd3BtJZiKU3ucomdLcp2sCXAdSujXA3XFB
7lCRWDa/yrsaP4KxNHqwkCJNUsfz8JvuIdaA6xY/QPg6PRCIyjZxPzyhbCzOefrr
bxSvJmwwcI5SHD6qf4SzHzaXKoQvTG1oDZkP/lnVCQumcJnODsXViG/ZLviDUguU
D6rln5WPeVsBAc4+xgFaduCybzNTtPjdeAsK+F+4+50dG44mwHvW7Ra6n7e2Pa49
beeh1hp9n1xLbozWqFX+PvGAADxN0OzLh5huvaaK9/vE1Ft5BI4PBaK4qHY+u1fm
jEO9fAGFB3fiwfojBgS9V/Ay28ynvBNcBDkGmwdwHzsz7/iwDPeBrMBlhxbvFuTZ
tlLmvC55/Q0XlnOhrwGLJd3Fn8+Qyms59j+XFRIAcIzXcxHVOv9rsDfU7uAOnZGV
UvfmVVEI0O1aBWSDrhDCIXuHIVHsO8PBwtDYZDryzv4JkwWqEWnHX87vkxB4Dk1u
wNoHZAVSfNUxqG5DjuUI4twHoPD3wszJY4ILU8YFq8uAb88W2kM1DSJ3K5dIsZb6
JsKNntl+c8TEknx7jr9GxwhL/4hAfIGwESa9NZuIKqviCER9VaRrSTpruV7gzlVs
hyvCQ0KLJ9DKkGVdKsDVlvVp5mVPEd3WKbO5EDFLi1By4C/AITGVnhScPpmjjtdg
oStnZ9ofF8nUgDWZtfEAjWxQ8SDcLCjgJviHAqfbUmBFLC+X/s8Wn2SSNKzV0hTm
vrYvLMr8CMpa68p19PkwlEHMlWJqQY4T7XT9ppwKE37ZMbOQ/vy/on8Lavy4B1t/
qoSvST9g7JYAq7G487RWKVfoIC9mVtiHf+BumvSkvOWWPNu9aIgErNeuLU8IB1/3
/xz6ISmyP7TEFetQKZbfKrIiimoPCRkKceXN3R2BX05Vyc3vVNNgF8ODdslhSkP+
JYgPOBPhSx6J5EwuS75DOvdolyCBqlnA+ey10tHcOycgooxGA3CUlaGg6uHlThSu
klMs4hLrdI6q9utED1keBS78W2WRbZ1bqI3XUb6mh9e/4B5Rz9KFs81NymCeRnY4
G47C3k6Tj5szHSMl9Z7usKkcB0/bwYQJcdHODi3uDAfe0LRc66+yBYH4uwaL/M1q
zH51JwzOLJAmYbE0SRkCaZ88KjtCf9dtiBj1x8RFC/BonCtYYmXcSsKQ42DArhZd
WZWDBzyo6KGdWhNNoZykgr4PtooLKd8Mx4H9kBnt3RsjZvFsAv8AL3OduUr3oFck
Yd+dVrojVmdiJq+RG3zjmeJiJzojUXJqy9nZX6z0JZ62Txardb4P76o0rQdqZ9f9
/X6hk/1Xz8MrwTsIbim50YMUS+3CZcAr0OuvuaXw3rZKMbxkqu56HYc4R1629fnZ
B4ZzXNjLYj2AF7bgXurh1MAwB+lJyLtpPP90SORoupwZ7Vl7wu8gFIVzT041O+ff
N8D7SJIPHz+62fVEooqgyAdUsZQ4tUX2xLrOWsm4v0H7wlguSpieCSVA+zEQ5B4n
3S806ZPPJAFuij/2yBm4cCR0cfnA6va0TjM0KJ6MnPI1R2q59eEETSzXuMHhO0rD
CuxCo5mjTEhryM31E+UcrO9JZstrKm03ALZQ77VL8WaISsxWlD8wyl522KkTH9Bn
xZ7hxopROGAkFRncx/+QoNjtFACxNWcE+bXgdxgkIIgmiSgkHxW9rrb+b10tiIbz
rjJ1L5NtzHlFC/Wmxoc0Y0tdsRFl6UjvTauNiD+6eBNphl4nNPil832yCA7lfypv
pK2PKy4OPpdgZYFHrLbNZn10kNGMRkYPBoMaDP9sRqFNFBGcJDTB7BxkkRkiu2vN
IXjvXV1fdje1ymx5KiMJVVUeU/Uo4lGM5tgQ09JYpYjk9oP/rIL5pn8Cc1+vt4u7
MONs+Hn6KbO6XYfBtUQPdIFUKrXdMfmGKgslkUH9FSe+Aq7XYE6R1vkuYxa5G9PS
i1Rc0sqjqlLFU4U+kH9I0Wt368mNAiUXgEf4Q9pek4Lbl0TaXngv/M2Bc3f6qi1f
+Z3HHcFseJTdeJ2qbk+EDKiSNtF7DH2atikPFeMoKXL+Bc6PgUTOGpJ1onz08kFA
dsG6Hx2aZJfPbaHPn3WxE/y1dvmScXp1/wbfXbIPYAlcqE5+JhJb2GKIR2HMSVOI
O01rK74LPBTsWx9zNpEAMvUEc7rWeaelJcNa/B7tqmyZbZdJ82e3Bm3tjd7f6M62
0XlB0LsnvyPIvmD2x2mn9kCYW9tOtQQmxlg7AI+KlX4v4erB4oQFH/2ISJ3lOywF
wStJYXsq4sERK6FnjwM4MIJ45opbcTJbev34ADdEBnM08Rme8kfo6NS4f/C6N+gz
rngblUeMw0UfTtZFpar4MTwVg0RmE3aYB1qcp6+aKFtwsPrxUJyyJc4KGL0O78IC
Kpr+/WZ3vHnxY4zjXSEndgb1Zu63jiI312pPfQjE6DIo1mG4A7rxYmB5FSg3BnF4
93giCFg2tRYEDYA1U24vFye6reKX3RT3MaHhidz5ZTTL519rtVfwq5wJSF0h9TyO
JsgFsqigDf3MPPv43KkSKqYgJAeLTwUkc2cI2x1H7Pmmo+JnTPfelW1+aiArtfMw
v4nImWKmFLmL5+j4vDuIi6hU5rTf66L1HDlY29hwaYHM4ZX3HbKlLq5TDFg09kyP
eWvHalbECePMZEAev+ESw/T3UjP457dvmM587mIb1hI9JStIzsWFqz6T2rfVF5ZP
PAeVCDo+qbzxBKMGOd90KQr8u4y4ISVjjjPedUx09S6sLs0v4LAvlcSlsznHznb0
pu01fZRHDMi05+Oi9bQTHcDP+XJVzGq+GJsjZ0Vudx6KtN9luiBeNtsDLRUtiBCe
EV24Uy7mL6NbN+fdCrBO0OOr5jL/7/yfhsjzLJ9Gyz6FlRpJ07WWl8ib58cA9VF6
lcKnDC04NTybM0pDWKB4RRML7CmEH/wT24/uAqA14s3ngnUlYXcMc3oArGbk+KAZ
zlciez69pPAOdh1ygwrjbnxDUboRhTSqIGtfibBXLqe/xIT5fYfb83X3gAS3gY5M
65aAU6mKQFz13bWh5NijjJHaZ878TBFhZvSpmBvaVYxI9x5ZIQLxwbAmxPdwrZm7
aJnd3rqxGiNeMAtfAYHzho6AhbeJIQ66ULIpoeTP70bWW1+wiw1i/vYbyGyMol8b
r2ikCfALxiCMSrKUm6VF8wOddwiXz78iTURgxPk5+l/k7AxyEIQcFpkV5X/xhkTE
B1lTh+KxcT/kNjZs6dC2gA3CbQDsMIPelu4cQCPxf1LtcAdrdAwOAQmmknvx3eQR
4QOgNcDRwhGE63yU1dV1EVm7bwen6n7O4EzHT4GPJNovSbF2f9tbf3gi7jlGWSLl
rToQONpQJOXRr1ou/eIg9eL8/JZRkuun2D4fkOup4biQ5hmx23VPCXzOo2WctHcM
R2PFqbT80C2Wic20Jh3QTQvWofmhRDBTFmfLIFtPjVpqSPHFbHGpF+3EwLmXulMX
cfNeYG3O5UcBo71PtGsTcM06H8wb1JKjlFitUM9iPr3c5SWYdfgUqJuXyZQYgTNQ
Sue9DJN9dxgrBMo4nxvg7wm0yGSZJP5pi6v5CUuceR1aLbk/dNv5oS4Cc/h6KNpy
p8oT8wwCJxSIK4agQUSfwmmMU7IZtwV/PHJLnnvYAB6sQJEHNaKxVKIPo6A8GeRz
hoyNShoFNINP50t5ROiQ7fMjHgqM5hl78DICh0DR8Bol5eNXuiduHhYgVe/7xood
VeGZkRomXeFzybGfqSAH72jflKX6CjEd6sLpLpYvjuKSfCDqObp3AlkmaEZ1Tc2g
/FSPP8/4o1C+9SEzm1gt/YOFZTv5koYH/M/zsLcGjHY6t60RO4DNZIbuAFIvFVJ+
uTFfDMdMFOlqAFH4N54kDwZEAqauvqURIzYOjfGlHK9KCQwsQnVCnniDrc3M7OI7
Im7e2Bd8o1ct3ne0cG8S9UOeIXoihGxlUPJO1ZT31fZrzjXE6GPTblfxfKP03ytF
NYGULr5kDU49BWlooa6zgHCDR41/Lgh6qAYJsiD8indklSTz+5Imp6UIsbtq7dMO
DQBGdJ+IsACxC/FqKWT5ddg4jkE57KyBFSgFsiJGQICVsubwFky41NMl8Yeo3Tje
4QkgQ7S8wj2qgw4voNIuk/HV/eXLSeSE4Kx+MIOAnWc7KicsNpvEaMloIPvBGGCg
v3AoVQsq/xyGv3joZ1ZAB98Oq3hASSGNLb/iaKsrij4ZvlmxioFP/fhb2xgG/LCP
8MKZc4U7DmrjkpmCCNMH5Ujj2hOPfuSmFq+gH9xmOw3qIh0hKocrydV/E7HHE5P2
6aSZ5/+Z1/8bUcikt1MZ2LsKHmYxqE7LPrR6h59W491wn68BF4DTmq4fIr8QcL5v
/hpnWZmP/rSslUxM8H0qm/r+ec9cFHYZThifsRMWsqGbBiQAVlm8PxQRA60VfgAZ
XzVHhgDTfKV2i7270/vIMnzmQNZrd5e56Rfs8mhdNeM01tSD0+sV8g2nG6m/JIHo
bdr2lV/w+i13NzhsKINI2WXVC8Rc/d5oXUC4c88vD4Uv2U3HGI939bnyiFN05auX
fQqVyYHpgzyO6rR5w3ahnpE4JSdPon5TVOBGRdSOvO7qAT873P2CAVuWiZZTuCi4
iDbP1+moK/sUi7mfkF2uxY+2EopLGnNaeLGvFBw2LkKonhLd8zjaq4YB//jtNRWD
4Re9uIfsXQet8zC8pSA6OR63rPb9qyzARrJi9PnF1Bxg8jwIFZlsfGOLC60ey6l1
`pragma protect end_protected
