// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
tHt2TbmW/3QJ1A5Fn4XwnZdpGMZVf0ZuWifxG4V2lu3ZIaqX8c8fw0SYNs19
IziwwoKu7w1jLtoGDZQYXhKTthSizP44QuOhOT+u0rnEpyq3US5NjbSIRFNo
N6Gt5FEHAarNuxSmffZCM7x1bwz/nXWzb/SYKfZ6cDCVK9+yHRyCEwg+SA8O
4Yy2LO7utZwAUBNihUjtIeyPtzFLHGCNE4df9rN08Z/0SKDki2iEeS9RDX6r
z99dkPujw+c7H0sVBJF6kiRjmTqSYFRDEbDaXm7PpPGbRTi3ZLykmwq2f9NH
ppZg/WCHBCLGtJnu83rK+MIAEu8zaFFcJD38Wf+svg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
M1Nj7I/ZZeDywWt72Zu5fEREXbGenZiER76Qs50jM6rJbE4KVsx3Tux2dfuT
gBk8PskLUsqlloJ0pPGSAQbhPy5olKV4feDYDWLcqp4TzaZRiH5ehAmfHm0A
gZMbv5DBKf6jRlLFEjNYDi3P91fLQcDwjkKVbuwFs/MQLfUPRTvr59BgBRzg
mhrN7U2e9ScHrlwNn2IUU3lEsIol9/a8em8icwbnTpSlN4tIjKQkroepjEen
RnbUHESZET9t+NHtWfAHdNnwX8a/eNDtxMsd27UOD7eE5VqeLGUlTludi6Lj
r/e7RXSiB1FoXC/JibwzestDKyW/PjAq2iCg3Q1/MA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
O5YKXL4t2EbNRH48HG+ibtaBQSSTb6+HQJUZUEPs+81k97n+kFfU1nT9A1af
iNFUYp1GtTflFnwwKfFVcYc86UzNAbhEBKSozOCh+w63JYjaeLUps4WKsgMd
RS0LCp1RMxneQOyq3fquaVfT7mE5iW+r7jENGTLzxTDg4z8poe8eU2bafdN1
70BQQnj3IfUadS4qZcJJNhKcFwBszgIwZOnFT5nwx2gojgkxtmZfhubdESc5
yVYDvw+1U+ct5BuW0Dw6zFtX6KVVVTJ35G50iTj5eb1DKKtpMRRcaLrt3Q6H
cgm1ECJqc82rtglxeovqS2hKgUAs7S3hbzoWeerjKA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
FPwoEl0cuLMruJkoaVQvGzGaj07h4xPm3uXemuRbG3/lioAIV0PtX9zeHPhn
qtFA9UtTM6mj6Xtk44T3YvogajfSFjoEdHq+0qX6A/dt/fi7WIsbKO209ba3
I70jAvroFN/4E4x9MpUenRIiGEofHEJYra5BeQYUXFiTgT5/9Ys=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
yawfaIMLIvqDwF7bFRfb9f2LXgkt32F7J5IXh5ixCOdUmx84MES5IkrgzQv/
5U2+xEObeegFH6kjzxNx5+SyZGbXHyb3ceTvCo+SKyWH7p2PpRFrjUb9auqC
ZSflLoCY9GtASxmsbtqjCG8xpDnb92iyt+kpyx4nQ+yIqXkEJ88JpSFcVMiS
jCe0rcMmHVaheC9yJoO4bviA1bIvXpAm06AfGiwR9pVU8pJ3OMKgrlxDePcP
tOFp5WzgJGlTQd14iMPqj1zf55RbOKSDG5ZAsTrPvYOod+HRR/4RGmOt1hoq
Jjr+fRkJ1H3moLXbqn80XwZF8eGUUyTxMpI7kVsZAyBGKivlpE9MPwRcpusY
KxCGyPTfe49bRbKkJ1t+sFp7LvI2WO+NdKb/FFiXsMCPctor5h03eP7qx3r4
40gUcWnb6OSBTLoE52l3zJwZzYUD5zBku1DVhcysOaPwPYfeAaLWa0YmDm6L
gaqFPJ95vodCm0JqicXpmSR38Sgkbs6q


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
fXHP+DWU1uqAM2KdSK04lnd4IcVf2+uCVnX8pFDLiRfgEIw3e0Vred1UmniU
0fnz9nvum1BNfGPVhdBcJbjkYfnPXvJU6h4Q8FQ9TcufIUWGXcRCiOEDd2CV
ywf7FznQZG2WblI8Om7o94+dj8SWALhsyJs5sIsz/inxdghfyok=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
BE54nGvQm6hg+fcpkndo4gE3IuYqYoQcLf7oTAp4aFV1NhGvBwmwNZ0/eLtD
OYQu55oyhz3jfBnPxpEyPzaPl+S4kif9ms31T2pwXpClIYPiyBoQVHgAZazF
M3oLpE4DXSMvNQnLXGwcxjch4q3ItYBV34ktdTpWK9TVJokLTq8=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 42320)
`pragma protect data_block
TAPrnCx3m7DI06KPGkVdqOdjkBx42EBoVgLhzy6WADlkZZPEyfCLKEW5ziqP
CocqBAgSXyDQxccq8JcvPkq+0c7AxAiKDKcjpPjOod2bRgBsHVEdz8dksBBo
v1E6y/m8vA3LIu739a6F15I1qhpfochg4e2a0RoFAzSL4b9IuVGlzXe4wp4f
csg50v7+J8Ki88Md/+wILZUHv6jyitPF2g7sedPM739ZjI6GPFjsyHwUseAo
Mv+ygdU57FasUkkeEuxDbSvr+Ui5cCH4KjIaExAh9Zrv0RQLO/nNciBffJuG
0OygeFlmc0KPMR/6k93gXCuupcxLjYKjY1z/UUi6LdN90QBtMZ96ZMdu53Pq
BtFw4KfgQY+ndDJQvN/3gCbOo/SV7QmCt1slrxQ79jGYXGNBzv8zd4dbwDLA
+aH/rcKU+odUKXG/GH3YlQL4hZmwSDdFzvicHB6KjsRP7oopaKDArUBvc7yy
Fa1gz6ezC1pK1qtRr/ZpWq+Exftc3FXwzG/a8I+Uny2XlABTllLkKScNK7wi
0kkrSKunBwH8ZtdpxgsEjqiaSBECaCfslJxrrVFhmOyC7/EA8mxh8qoqtibu
Em2tWW/dXvAE1PVuQoviWe15Vpvr52K8T8rk/wC5n+cB8ZrhIKNNlSWG+U6A
9fwIO0U37upJOZXZGmZE0N+CDyhpEw2euQwIjlGO6F84Yi0p7gPaSUFSwkh9
M67LfjnOq5Mi2sjNMuw46DtdhCmmNX8uZwF/b56Qys/LAl+bjhPv9FDiFdpe
t0omPkMezikU5X2dudTS+vHBoFfpqkYIv8odDTAp3fbyxv5ZHQ7UVZkZ8uLM
RNlL0i7ZMBnY0F7ULU5JOIJsz7k3zy+3g4Xhf1C8JqKd4hYZ++28FXfhascU
DhhzqJkDMJGqEaIGAIcUTEsZ2fwJD6MFTaCsyeRNsN1Sm/Kq/Qv7dMg34SQ+
mM5wzFDGvBzBfDqz2SjYrhzXcRShj4/udyOg7wO95TArm1XL5dvBXrhooGYu
GJHya2zb99ZpcGm6/42vn8REYFs61BSgdB0Htubl4o80seZpXec39dYjJIvc
VH+SHDuxLCEY0K6QojDnQyXxw1q/VYoSbDutlS5vjDrHpEqxdzz+MOoSz+pn
FowagifSyMO3wWQ1LCcbJX1HbslW5XlweED+JEtFtg9iiYBJYCw2ufQkPNAs
snLzcpReR298sRizsoaRwExfuYk3p2YsZCMTWd3opDvUB+ZNaPoNX/JesI1s
ZMUhSrOPddjwCgFW1dTPqCbTRLq5fnyQ9wNX1phgxPCN6eaqwhq9rxYP9vf8
LGtW8D7e3E84mzMgA6fuGBP6A+Lmn22pmrsmbFAxut20QP+Lg6Px84iJ1DQ+
cKhPRbm6Ha8/z39E0SDfTf7s+kn+R2zFj+QpxN6RDoJ8h/vKR1NBtVtBDJbY
/TmxxGnthG2cjkCmjsin1n99o93Hxx8ZAWzM2+dRCSDelpIDYciZWU65yzld
y6HNkDbDC0mtK6PX90QkpPyvqN0IeMmQZv+pNYzqK+1DvvbZq44MG6q4ZpSV
SRcCjMUb29YZ+NBfkoe2p15ZL2k+E2yo8jMVhhTzVi+XwVRPu5jQrlq1Eim8
4ha9F81QRNTcu89YHufWecAPK+6hykIv0ec72Fwr6DjtGjbHEfbq3J95murR
QZ00LbduAEvPYhA9STwPqseDBEyGeWvHerAIHv6I5yhU68gd7k7/QTCFwJQy
jFhY63h37v7VmU4pOlP+LSutihRkUelQLOk/ReoRQ/1deDXqT0pNp5UF0mDy
4eEGfK1xGidVA8lHQvcsEQsfPtYjRynnoryvUO+MgWCYOPLAkNK/Rqkkvcqh
3VeaWND56eM/mEOukTdyOH5OimMlGAoI/gjpgMEF+4VFGhYk7LCL8W582IwH
12BuaXFr6beEMUsuujv1c41giyldgBD86nX+o3uypKT0BsLzTNN6zKtKFXFN
Dg30ilvsZHg0JUR3bGJJp+o9uioP4jN+0oQxnQ5Bl3Tw+XGamANNoVJHXvMj
l28eu8Ke7hXK5QWigNDe32G/qrhv//f4W0CP6ihyyOdeXYIHv8ONHbIs9/w4
efZ0LTTDp6Xyxg8v3WXQwkl6ZDxokUXEu3U/zmJe0J+CacR6ISi+ozRa2XSV
w6Utje6Ez4iWg3mJhIQVAewlyr3fimbT47mte161EyXS9/6IQPKXONk8qJbl
drZ8wNdyn1iSW72ElW4haGgaELiv7OUFs7pPqt217eOLCdXyzR1u0wQsXHec
jK2RIeBUiZdIFnVZz18aLkkvnBmHgstoOimm6543Qn1irgBePiJeKyezSEY1
vVs9SKT+uwbzzXRuHtJEV6yjl69pze/JNbQaFNPhWoCZjsgel5K2JzPv/UTw
KtIeZ6yydDVV+QR8TvehN+BH3qMmyQq7un4LIk73G/CmFYeqkNICvtUa7Osx
gbbTDFCr0x4XnZ8z3KdnXwqMKnonkL/6gyAH4QWSZYddx4agzB+hk3Sgo2YV
ZtnfYuGSbx8qtai/tnXKTmNwDsaJnfePqADeU8btrZWH9Qc0azLBelBPHRaQ
xemcQrzTBQ7ubqR9/EyG4bP0wl1s5JU4H6hEpZcxXRJ9UQV0Dn1rA2dTWmkH
K1ervk2FOFtYSzLDu7KEFwwn92SIG1xtzGCZ2dTUqC6rJ/+4DO49eiqyNv5q
5YLxeiXufrHNH1FKZiiQ8fSbuK8oZBCIBs9sClDYsTkPJQDsF/EuaDOAXqI0
1/rNQxVsZfCHUWJ3u0ep6XbmXmM9m426pJQytcaZCXw8KOfsl62hOPnHtXiD
UjsHW8tUjH9KK8/mUsar+tnfUNnglzmwcqqRS+4HHbfZ2aPInCsU1z8b6stT
vsYiO7GYfoGaPvh7i0el/CAiyrO0SwR3qc7JEqTGa2SvAnP2Rw9215iT1M+d
tozy8xf85Iip4cRA1gB+DKz4txkgQ4eFvKUmRnfAI42yBiQWM7wCVlojE0Or
Ro7Gi38kfR/7HDkuISCQhuYVZKaJwvwjf+TZ7A/7HvHgK1NWVDxDa/AoERIA
c7s/ZYhNAIHoYawdsfFGp2+3eWy1HznMUROUPgJyyfc40l0+vJIoHSkto9kg
vdJCMUP4Supi9Mnr5wtZSwdbjLes1t806ZoFVI6PqUqUEyddh3yd2ibrqXXN
v6VgSB41iKrFXpYvHWusyJecsM8w/AIRZnWRB+eF+j2oMYAk4hmAJi8DXU8l
kdi2yg+98BPAPgYlMO6gD+4kPYo71w9M1UsKGq1WmvpJs1wTdOvW9Il1oUHA
zcchvzh91ThRDN1Tz1C9ZFyzOUh40ADAoP8855zmHyf1LAn7W2/eCvnQMnR/
frWLT1Cmw1L8sMWjZ83dCKrshBKUD3Qj/Tz314lMI+7CP1BAS/TiGVUHsJBI
Kq8mfoMwnM0SB4UNEJFGxvHZ1ERVO82Lb9jFGnqAVof6UG33YJxp0bxAviVl
UPaLiB8Y7MRbueCEfhCQ64nvcqbPobgXiIKIxeu/y6Q0uHvvbxxWGMEj8wDc
XE1iJhhKWfbg1wkIcZ7joYvBJk36vKgLzc/R9kmdRXGppjvIPBmxVmxZPSKu
qO7+L7Ofo/qs5wYLmP2KMuoyVn58FPHPP+9qcBX92dzWSLlMJrcAZ94jIzbA
lZYOInUY8zQe4RLfiDJYB6bFYRIvF85OsSa8jOv4ggvazK3Dub0G5OcMDnJj
K8tHrYU3xY0n7+4p5Qtb2dcyqV0scHGkhV4olUj5Lg3juIqHuTrke4ayKLg/
aSj8Iqc3f/0pLMbKZcqLfUS37KyH5A7LFFyNpzmM074ubNSBfZLGwFtwuZIh
GR6nt82V0AShdfkcLW4xV9lxYFdsOaCJOxRNEuPcSkOX5DlOB0yMtgh6Z+lr
RxuUcdbb3mgCqXwM7fJVp54lu1nAIrjXFf7e9V4HoOgllgVQbgWPfH+6X1cb
IQE2m6S+6+YyQUd0m6yhE0jLhN8RiVaCv3soWIiBLVjXuilN1Ne46s5yJlFH
z1DLcFuuhEqsZ3yNjGlrXwA2BCAyL7EDOld/JUiHnv8+DAUzUYl9RNV9f1rf
LOdUnWRLOFJnY9Q1yVulYzq+JlFZRD3oHZYpPm8HILCG1e071sjJYvxZ0JUg
5V9aUquYJKSKQ8ic82mCi5LQdX/x9gGgMD2AvA+iI/Zx3vIOvUV4BWpNuemQ
gO8wuYC34zB8ueMGGrDNWKj/sQ2I/M4JwiB2n+Cy9TcdkenSp/pLETvX/+3e
X/R+Y4/jNjUfMN2m9TFxvUZZtgPDWpxx9JeW7k4S0frDIbRf6O2lLubjgkwl
oy9ftXn7MXeqsDdlV6Alf4VdzHevf2FP7xvSvUfTORn2bJDSsk1ZihrSRoJX
9XR/ea58k2mPDqhc3wxJVPNONaF4y8DchnxFBL+eIb4jsrujRf3mrbBiJ2Ub
Slum2GaKijdKnrrpNH/eqnrdL+XXdNEU2S9F8OtAdvLQBp+OkQdiiPwJTwQw
vqL6RYykujC2aNlYlbJ10xgrStqa7detE32+fbs+Jmj79PC8NmZ+iixJuuOP
osFyTWn/lzjluJiouTaDSwDszQ+resHvH7stx570NKF1JBZ/v5kof1MJtJ2l
rw5Uxo8rVOTQr5MhzkyvKpgEOcFS91fyrQHIsX32wSgUW+H+Jc6XqdghbmX3
Tkagfiu7vTw4vRo7aq7Fml4/x8zTp9nkWHt5RVdkV4Ln45OU8yjgjawH4t5o
Y+ggoKDUIJFO5KPY7Hm8Hebw5taiAYulWJVVwjfUq3vO0UTUA038utJLlNp2
Og+9Vei7gVH7kg3TQpusqN+9JyYRJHiXMCWh4qXMcWWGjMCx4VsdLG+FfSC0
W0KTKCX+6W1YNvpveZWo8J3/taVYCGxkdFlyzAWuAwPhrlGoAokgDi4p1fBL
bmsbGMCQUAcuxylWo6Rx8UyqWqrINK3wDFgIBAjTzTglKDeGP6vZvdSDJuFo
TDaI2/4bf09v+Z22jxf+/w+tK1mJ2Nl7QS7rrq5B0AZ+y9tNEMCRP0oDh1s7
YFKKT8gR7rudsJ1jT6NsO4+AzJ8e3x1Qq8ObIxLLF4rQ/OmClIZ/yv7BkhtR
dOxT7VSOcO7SaOyMdTDfcRPKMKpC0dIGP71ev3L4Ofw8yqRuLAmXSMxvFOKk
0KuB4GslrtlEmG6IZgQyMo1RPBU9xJBJ69kC8iEbEKesZeFFqKbZPID1Q5tK
qR2jnA0Azq+cjWZjItg1jpNdk7kVf8eNTkg/eJTCohX3dOLY6tkUnbBrJDaB
kXPOZ5zoaTM6EFBfzXwUoRsS86otMOCr5exy4DpFJO/U6+Z7Si1QBAcxPTFY
L718L8ksUDgVODleCLG6l3lq7VtiuYuAyaTeePou2+X/JCfMNDAi9no00IeU
DWB5yv3nwQ8GBUvbg9+/PvVBMXrac18x3vKDUZcptZy22FTErZUR2/WPMkJU
qyKekQ8Q/sZQ+96IX0ur78w8WACXhC74aW7U7AceWmHxQHsEW2wjM/34Mfdi
O/LYTsVVfVbvOImkmNtT/eRV9S+dZfsXlbeQNDfBRC8OKYZDCW9hSPhIOmTU
1JycbllhhPY2yex6/VaCvRXNxS6q7VBR3kEoh8a9C6XXtHRJ4JkWAOTmyeFo
TZtI3jHJ+0pG475jUZ5TVWH2d/bton5wMGJjd1D9guLya3vqWv2A5hxzjfcN
2bSriMmjPS84lFCAfQ+5+fX+bTs8zCSRqT/7aMu1kdgMogqMvcjv/p2yGiFj
kn9nRQFYfOjaCYsvjMUxcmTsggyIDh74WmSosZc6SLAHdt7X2wmNV5SYk8WV
fjWyIYwc6iApAai7Labz3Ghtj1/2LH/1f2+viUnZ831ayoYMeez3IpOPYnpW
WnDBcKTyFjnetFMuOpthS9HkI4oE+nUaIRdXPRslkyzOZRtkahC0+pn+B42A
xkhPz/024TPsoWx1MJZCQ2O/KLo7+P0scGHyhoyKW+W68VIOd0rz1mA9qZXx
IgFdRrVw5/wbDg/gA9B1lmww7eOSyL39qy3kYNzFYhwpmFdykHskm2yn5k2W
GNtHF13T7ckz5uHn9beAz1/BK+a8Ap1rAEuyXG06RQSzNQdJho2/dFWu8WDv
MP0KCrDuWANO7uKeOV3uFmihQ837zGygsu+D5/gPD6xGWQZerd2+36REaZHA
n9mKMBQtebZUWczz8QNMSvEc8Ovbt0hCR+qt+LNef/kidZi3ZitwquqZeqsy
IU7dv4dO5XdHe7zgXXcZLQ1YFvxyNWrUyUrlOK89y+5AKU5EZTaFD4/jrmeK
1pvcIBL6oO8J4+uh8kgvrWYQCWpfppI+EsBWFYSJiXubgDvEyNUhm/Q9O11K
Xa3MkLMjH1887BdxFpS+dNks2qH8+YGkgPLXbXy5pafgD2EFzE9XcnpTU7Hr
mw0E/ozOCUsgZx9Y75LHYMhcNB+vot2jkg6PqYh4ImYvrjy5U3NDK8tr4m6j
uJAIPQshjW+suOG8okhFkCy+6Q53X1FmGs596QLJW2NBqdtNjIfemTGhSGIq
wy7v/WIWs0kBqKlu+PGWwIc/oMJuGmVc/TF4Urw53+P1t/nnpD1Z6MmBPPns
ByWXbZj4E4eIpaerb7b9f/gbS3RBHxa6b/BkyRvCiL6J7GNj00RTum7VTydX
75oKl+j3wmWqvCCFKD9AOyHy0wIGSSzatT2ag11ov75yCsI2rU2mWUYiJwxg
onU0chUK41z6n4BVIUm/KntLX1PsTsiKlURvfGyVeR3+Y7yM96diFpndx9U1
En0vemVfyJCp+gxn1vXe/X5ORqKdSeQBZ84F76ae2cHXgEdj+/2TOHNNhbJ6
RK2+Mxe7F/UYU3ayu98JFvPbjfNK9Rxh9yzJjo+TUxIFJIeE/4sZUwIBlvaN
Bn/67K0iKxVXRihDNO2RXQzzyIiudvYRhr4rKuMf88ve/lEiOJa8WmQrvwQs
2PqWZnYd9Q6JzCPl3N+i+xMeG6ZQIaoaMwdWghox4H2FhSoji/y80Fm8OitS
/GwHiRimyrjHi7bh7Ah50n/VVaD7PPSQw6SE7+bPEtCXrHYfezPLUyld2ic7
6o/NSMISavkLVa+SBpNFWKhovszL61cx2mZoQUlqcaOF9lKjfZ07xf3WRHif
zarMIpvNggFZurqTG2PjPCxBxas9UZTG1hhDzv5OQfKHFwgtEieU/19hWfAD
DhWO8irfHAfJgtnxWk8xW9kLMLPUiCLzSAPGifZ6Polr4dCfk4Tu5Iggs404
sI/a7/xb8GY+kd0IetBfGZ1EhHDN5hFpN/n5tzcrIxAygZpzr7kE1mi9VGf3
bqKbkMoYyRfLiwAE5EXMxY1Q09v3qR7dfeHZV3j4192mCQhM77Nt1EzSSC6I
5Xo6q2XWnuEjpLcxK7BMfTrpcS+kNw9PrTq9njUgSJ2Gyk/6CAjr/NLB8MK2
0A2o9leBKdVO4oUlfbiUVV/W4b+AQv5IQtiaXNuOw2e2s8IHTHXPFLLTXNHM
zsd5SdUDH/zoAcYBXXyEsXGV2aQG+w2ayiV9dDf7D8l82UgUXvCVoDxXU1L/
X4ktFRtF7dJMltdNfEV+cBvRLEOTBxT5hsaImrcG6MEuk12ysF8kTYdBXIzV
0vUcNQeCmo06K0nb6QYJ/Q88kJnJR8Kn5VGjtciWZcfub6jWDFxaXGN38x+1
gJTOD4LXfq6tWOr8jz+dTUfBGgZKDar/TYJb2wzVu3pVSwNZ5Xr68D1ZZ37K
nra8O/f/ODfH84NCWTAeCE8tI2WqG0yVIEkQZnIIK/0qjXFDJteLfEKsoUEs
vihiSpCyAL0OW0CvpWDAdA1NnysjQM+oMRJ9+94oW7nmq853BV6n4LaHxMqw
UBZfKN1K7Etp9ehYE6Jf/QrpEyytaIbfMYBZBL1fcUTwMi8z4Pquq8XMfekV
xXqLDyc07mxBuyftrNviAAKK0QlOmgteSZf13vagd0SAkMN0IeDIq6erAZPA
UQjSg5PysPJw8vDuiIOJ6i8OXAlj4BestzWveen6sPU1P3kEKb/riMsMliTd
4u9wRkpimwLWq/Kfk5pZxgnRZQ7zd39naEfSOvsGO/e/qGwsbIwCionDAeCo
AQj9AFQ22lPwdDTgdlQ4fyK5Z56Ia+yIUhPznZbB+Nk9eNC3N+TYOyIsLQAC
mc1SHQNmwygTFbGqOJKsYIbZGwmXTZoLh5RPz91wcqoxtmnuiGikGIOUAU0l
q/Ai2jAVJFzh4siaVVc86feBF6N4FkWUBnntK2s3pq6A/4c8Epe6/G93FkBr
IWmiGzwmwtk1tGL8Whlt3bjWPYx5zc+3sTRUPpEN+Oy0xcOlYl9QAtsZx/4D
t9kmy602OO8cJGSEIUnES8mpK0Bzx11mwj0KN46vrVsXxL91Zqmjzx8YTyBl
MJlveIPjCxNH9yrZIyz9B1mavOFuFiG3mDFQpWsmwztKvuxzL7gLng0yaNoD
mxGtd4cLkErTClVTvfDEzG++Il3yLrnGcf0E5qbyjX+I5TofR/50BWToHWX2
XVSj1jOlC+0LK/sU9iPdWphy4N7N6PzkpnJ4wZSrw9M+7v7WBx/VOtX3cjW4
0ICVJ/9+p53ZJqLy5gxUx5nMTIM80aanwxINRt34r1HP1mcsRZ4ERUj1GqNh
A6WFUpQvIeZnmKhkiAFGugs4qdCS2JW4/XFyZfov/SKFcVoiUzC1Hdvq4CZ2
Y/zrZ2iC4tc+S1nveMmXG1TEi9YQyLqMVU09GQ9gCSg+1073wJ9dUIq5mkdA
7SOwcxaAfSm8ROVMRrKs+EXKDsv1gnGY+xJXgAmuSP95ya0ipfG1CJpj1k/O
vDI9ukovxXXfYoh7G2SzoNNCsbP9/g9CvrNjkY2Oz9M+f4WEJSBsipg8otJ+
TV6pyyKaTqxZT6V329i/OCzv8GxuoThuFxrpetJD6J4M7ob3UTefhClTNM41
34mV++4/7OtHIqkgyxfsu1DzT8YE7ffA+i5G7mTcXK9CRNxaFnGDGMgj7iFC
o1gv3/G2FpsLa01Hmt9TsQkfetG1UtEdlUiEXNYooO+YY2KBBY0SphIvRqpW
EZp6dVLGVh+A07Lyt7GuCj6PL+IQuhr797lmBe56ei41RSxmI2382YyfNT9+
RRXsVuKr9BRHRRtKRWbUAznuMfysRzrKMqrCv5wvEufsuvBKtmjw7UPUY2ca
6SKBOgeaShhrFtPc52/ZLDl2qlN7agNg2dPWG+4VMuvTMqWCm3Dy6vh3cufJ
XoFVAOWo/iExewTP80Dft2xAzjxpopym5F8xjFE4Ly57WbuXLRBV8oaeRAPl
bVPvC5VFX16yFeUblzilkvjR8hhuEP4nv7plL1C2Hsl/kPZh4VWZr5q5pRz3
mlgfmgu/KpmbMg5c9kNSqn9qHrifVc7nI3CEa+B26jm0/+zQvAVL8gjYWMoX
5j7jdsF2TnhU9/1DEdjogY1sUHyy6wJH0GLpNxhqUBNu0mbC1ab7TmU7wRgj
UX3wd48nAF4ERFum+oD5rexPAjguS5ij9+CPe1Qx/PNmG/vd/0DaAAHiG6/R
eaK6KsbWVz16MWOl+EnaSA4aTGFQLvTsZouWSXcygn4ROfKSrFfNuRyMA6Hu
TeqgpcDW70E4+u2BqFbgfpCTPQTAM+lgXaZ31BdnQBZMGQFixOZNvCBCxgSh
YGxvP/Bc75reOgNwFvSbI7DFYFoLC4CEd8gr0JXk558IMrjaAVTnxePmOEvW
9O/cWBkuAqZl7eq6S00QHrJ4ZjMJ/zdBz74Xz9pmMGdSGLbtv8vjMe4qpJBo
zp6Z9OYeZ1tkWPx9A+vqu1HVD5zb2OcIsV/Pr4guBomc79k1QhPSWSeqw1zb
jloUrHlkW5KSe1SuuUZ2ffCRuaWCwZqYIQm5tp095ed2NJt/Ci8s4969+y9z
a8OM2NPBHGfkBK0UlGzgBf+YoL5Keh3fYyEERvA5uI36CrIbGuYRujq8N5Qc
qe6UNNZeR9SVZtCVvVmp00KnzMsjQZqastRljp+Qv1QWFyJN+twg6t2o9KWd
UTgaHa53I80PCmJmrp7uPZlkhEv9iqr8wMhRUE4CJV8exyX3GljZnUyoqiKQ
G9Avq7lW64jCdDCMflA79UPpxbkklkayg60PCyHSTt78denWZM3Zp/YF6rhU
zZEYaTz/3+6GlCS8ViZEbVne2y3HrUGP7H9xEyofY98HSaFO9w1IAFEkXHtQ
sDOp9A8dNco7ls5scKPR2F2lcbJy4nDi9IVtBTp6TMBIrytut+1Qwc96Y4VU
s2tw1tnWn2hNclE/JeFBr3IFDYD25u9rtdn24Lk4g7RBvXE91f26khuo/JPO
nEKXJUx8uPZ4/A+IfF+4zB2VNxrtN3aqdleKHPSLW52Sd2pYQXfMjsCEsSfP
DI0WsaaO2kwLoLD6FGv4uelocT+J0GlPn7EbIIAtEQpMOfwDxoY9w3Pa6e4Q
mXL0fVng5bU1G+V8eOV3TTc3Cz/NEkoKeRRWVBQLu8P2DRfBH3/l+p1VXnnx
BbWKs0KKLO/ndXL9zsyX7pyJU5RxYvTfbcRUDrIroqR3x/ouabzdgkFzr+zA
7Lki9G/34r6LlJaHm51SzIelKgC4eAIDV8T6Vcg+eDy5nFXXttKjxOAChOVc
ogJOo2ujDSf9EkW/fdSJ2tOHb2aFtxtm3v13PwJ/nEIuGerYD+uJHkuI3tud
rk+6wrHDWrHSCVO7ERJDT3WmfhMuJNsKkzhtLFlDYh2HZQbd3UgvbMTL5Uka
kPaCPdrJeIHq34E+Qd9zVCBxk6tcgpe6rB3vxkmhrTZrKfzuV7OccJg3UD1g
Q8NqEgavbqUR6WjCgb6Wrug3lH0dTkAGg2Kq4KSSXLkhNtXYSjvGH2tNrA1W
LnHHMhc2SiHk1Iz+7OKyp+BN6kigN4bfm/4bZPsR88gen8zVF42Ziu7bFpOj
2mnDxYzuGoQwkN8mO7ZV82/+19bruGk9XctjC7C2uv7aSpMKnzPbOO9XewDV
y96Da/kxKCwJ6ohzI5kLDGS6jDpZdG/R9Bk93N5ZaUWpqpI3VobhGPiBIvCf
sg1cvS1GUbrCA0+T9tRX8O07eW05TsBfZ8XQ2RSIoQW7Hx2NO2xYT5APCQhj
TfZuxKREFaf+zsTaHd/qtLRnhLmA8TxZmiS8shNE9AzEED8L434Rfh3rOoRr
vP/AEsFKjTRdEnivwB3JpwrP9umh4THs1NWUf0/emaVyIHTd/zzWWNF0dkjS
PiIEbg4XaeGLWgXjIaP2FPFs/WQHaTokMUPlit3PtskZtH/MOg4t/VqTFUzg
UpeDKhBxv7256jKc/s1n+TuXr0mAXMKz89hhiYXhTG0GcrI2noiiHWersG1l
cbYtUhTKwgnKL9SPFb//9E0UsgwSZEgtJb4k1Kz5Cmmi8QYsZ0WSD8i00zeS
dRZy69zmDRAWYheJN8ZAFL17r9BVlpNh8nj1Wz8wc9HiyMZxtPskiCJIfvwP
wStdGOj6wgJBNatJ3V1t3KQfPGovWg4mAzAdBH8CKQMwg68TnsNNSAMwgWlT
6m9IPOR3SbpW+9XnFDL0Fl1WKeIoyazILWwSIIRXmGmVGgFqLwEvOISmuwoh
SJ5r4vfTcmVA0YquSlcjHjaKghD5BCd5Gt97A8rWtj0f4zfv/rXXVZCG6Mfn
8k10BnB6C1yCIoRKJ2Rs6w1ngS9DF7YAXtONFoWP2+i1+alUKdVD8WBCnkh0
FPH6fmRPHEXN1U4CV9rgGMoAX5GaeikOy5N0Evdi4B3CVF8Cb89ZrNye/LGA
13ayRCk0N1SEwY72PoH45SQXuOYrzaYnL6LyY8cNcu6xk3qEC1y5MXfEhj8W
i/oc6gjznLJmX5G7I3czI5JBYa7Q6g2JopNMUNI9qJSm8fh4WVi7G+1pfTMq
Y55ojzktgMvXjvV5jDKdpM0YCFkFSpQLPVIDaUqYWWQQtRTj1/QxLLMN+1rD
hfApKMvS/bUJMDuQE5TaMAlHj09fGsIV3+ncWAXk4ycvb82B8U6flUdcCQDu
nE8/0IrzSnvcXi7g7QAab/APfjltZPrLVsnT4zeN0WW/5ualc9kA8nyV1q7U
P/hBS/EAVNUaW6jPeCOl2AbRieJdcwRFe26oNqzvjgBJpBZUQsvkb6DfN3S9
Xgoz1Y7Cadb/0qJjp13gSIdVLP0qL2C84FGT9QcVvJ7FKagi35N/V1VTBFMy
3iSK8DxhRBW9YmU42N34Y2tjOkomHRzMquyRqybSNKGmwi+CsWI++Z3oODq3
7SrVdOjyIVHNvtk8r95+oH2jMurta/I2fMAkGc0diDeBSOqMcbg6GfiJZSh2
oOdSpgB2JKLioya1n18TWEqnmLxpRMOTS5cmR+j6JBVdMmZbg15ePSgtmTIR
id5UMwEJfvlzME/XyQXexwzOGiibOk7P1kqFvtb/jj+DpjfqYU1gatRBSpyl
s1zBxZ5o/o/p3qgKSA7tT6m8Ci5x0sc4ZVJbtr+2uRZ3Wb+8izMS/iXgv2vZ
yAnpzT/SlVZNaNLR1gY+mSTyCAaE2DNnuicvZuXLksXfAgrf9AShcIeEe2Tr
V6Aa+XTSAJR5FrrVSP9dXPLX2nwlGZS+XHK0ZIijnyAVsCK4yq2BUKw+0i+R
NFIOCt0G+7iVfZdVK8WYHGtbXF3/AqowqSR+2MsAWv+BwNTZdN74iRlCa93u
2tCk4xS0yYYJlXiUxctl/RFRY2PtXaJRs7yT20s8PBTVGSJ4+GG+QuXbjYOe
nlXNF3l/1UFA/LAsVnWafnYKcjVDqwQtsE4rAPEAonjkUjvbrEdl+xVpodWF
2XhcXi+q/RFL+7XmvvPfhM460hAQbWklvrSjaTlikJ/EfiHpilfTU1qwl+eZ
A3lEXssnJKIVyOJHBYV8hvM1lWTvylQm1HjnsxihOEew9k53+6VxHrC6e51k
CPRO4hoPO92lpMTugPBDdh/uxLhJc/FNXFX1Q+nRjEgqbTHUf8J09+NZ6+pX
c1+ZpT9YLcnVPDwoZ8fhBrF/hTVygaMQHP3J6AUM/b+oiON4+v/x/gZmptmZ
Qhqa+i+A02y6wohOMVJDzniwUiXzXeq8+rcx3J07nijiSXmwNJNbZNEqHZbJ
gVuIzOLDY8bjBH6ShjxJpgRFC7qfZXloM6SFnl3HLDeCBIEKax0ct87nTcjK
DSYq7221gKhX97Dfk39YDEPrPfIEpbLtfD29m7BsZuSP8pnLb6uIqZ2ffB0X
lvT+5uzAuf7rhd0l/aTQXG9jC23qclkZCkecC+Ca0iteyuNtQeCFk86VRL4M
0q1vuuYOSjaujaD6RuhdBA2j4+FvcroXskH+RJkkKkLYgY+aTPhEC0mCmE9n
qefpT8rPPwEVPlkOw8AKJ4wh85Y7eJ+6TSKo0bp4/42uo39piZ5rTpWSUvkk
jpo9mDQBMSub/5mRIm7ssRfWjE3IPlOkprVx1RlEp+XD/qDatUpt+2vlkyQf
VE1Qi3fHJUQFGMjgOPCEUoy94ONe6Jo8CWSIIMqWSIeFYcoVJMQhxEhagIUN
PRxzHhjO/ikxIc+5ALe2Z5cEu6TgIsmkY30EQ/+BmEXXqFmIQmiFo3f9FD3A
yXJz3gbVcNaqAMXuQv5K1hH8isD3sFB+hWT5jstesMWi6RoElNthHccjgoab
Hz6ndeEfEmy0l2iuDcUlJKj+V4l7xNDS0wooRDVKR+70RK1Y7bH2lOIzfqHI
t6KgMvNC6eemfC2wS6defhKuL8uXDBI0Lb1NXyedCK6iTyWcCiWB3hwSPSeT
PgB2qRmA+7vzs7YSWZFUUnXwepPr1QwsAe1eaDJ+4Zn/tDDQ7xXtnvUgNPIE
L7CGm66I0h0vaB/6vbg+Nkknt63tUPBPVaqQbQDFupMz7ivbTy2vv5Ktjs5W
mtprMH3P9wxWXXOaihBpaFHTEMRCrUqURvW3v0HQs+S3polqEyJ427ypRaLr
RcpVXy94Ky6nZxWQkEsZZ0A/vu8HjR4jhVaY4RzVorPXr+3WoM496QyEAMvg
F7zk/A9WmF34DbtCCQw6f6NfIgZBpSZfUvAXd3m/k008gtwBqE2G28SFivYu
isY94hfenHp7QMT8i8iNWSohPUM5nn4X1UsUds3HxL3KJW1wA4McLTcgeQVN
yn85d0aB7rmKnCH5Mu0/j03/8mvY9iuiSa/XRJnJ6SUb5FWRX7clIMCWY0HD
ZBzNN3h4m5C4egzME9gm+3u+EWIBaTzr30+ExYbzGAMHws4HawwXOv5MjgrR
ESrN0KUPmc5Ylo0Qex/7QYG7M7QeNiv+Bl2QwJP2oaz/hO+IP1jfzlDfeeAu
mtPKXqlaOKgp1+wjYgUPZRmnebNI4Q549akIGqgLFEXh9O8KquooO/+aCa7O
AAdn1RsqVVELopzsV8pUm0Iiqzy6dT74RdtxAH60Tets8+N50mOXyS5tCPyc
aF4gRFKZ7fFdku+dYFSXO302lBM+Dtwm4kxrKv3ySQnUX7LstPpraP6ZYdZz
ukwvegEv/Z6Jl1006fWg8XlZwDfsFg38kOB0D36F0y0ROCsgzixYxkbn8fMP
mFtm+xsQuucXcLy3LDfbkoArrzzid8GaVho6wTg09NCcFhXaVD96Mm+ojv0B
Q+UJy5bdZIqEov7y8gL6cngCm0kjsrk/+qSj+ngEYT993w0OlwW13Iiy64Nj
/wGZ35Kv6f8yJ5SH6QppEVS2t6PSCFXAX5SiuU/H117DLuZbhi4im4JwralD
0b/RTDJbQqT8NLjR1idbmXdVKinSFWl+TXBW/8nPedqco37rcbJFZkR4dLhH
hnZofmkC703MU5DZij25+/L6zhmavpXX+nyMNrFPQ0NksZdN1LEmffk09TcZ
7hBEBZEeqvPyg1Z6FiErOewSxzwHvGJxL9FqzDE3oIIJZq/WvGuxqX3NUj3S
NhRzdGh/jjvCkSKKxEH17TI2BLMgToySHxWO6/79oORFc13BOF5QbthOQvX6
eMC4gZQjSI6B1fyMUb43CqvqKdMjKhOEcs/nUUidt1WlInIO3itrla+pVh4h
xDQDeTXAT56rTpRXniD4DN6YwmPVny7qtKOkypWp9WjNfwZyP3C1QHxdNAFc
JnCmgNCzicun2Lul4GtdB9+zcNRnGXCT3fsctuQUaMD2ACDoLCCl2Ze+PZjt
phBzBVpax2W9xiGJYtDAo0U88gUAqiRjzmueSuU0wp3iCT1l4KU+KDykfwBa
65erDd9PB3aXL89U2kmhxP/YpnyTGD4zhS3ndiqiul/936VVJOaxxvmFc8a1
7nQ+C965wTZDOn93RWkS8z+8EaGDFTtli+pcSsDA6tjDaRJ32zEwk6QU37XO
VBZQnvC8eHzXTJZY7v4V5Lni5oaMKOiUZzQY/I7iVBqriHqzR51pYv5EXG4t
5v4AVDbvHCh2soBrbs+Dup7wLYslNzg5TGWEdnFgT9/itqWi1SKCvTgBDQ6+
IEc4ftuFRfAaJ7HkZibSaZnVX70a84aPCIv0SEmt9pPQjdU/GSKi2QXsJZig
GVURCRZAFMR8HdJJlWWj+CGjP0BTLV3g+hdIxAnHGlTVPdJQGeXlW4W+Rgil
lbBp7C6qEykK+O0aGoHe704jFA1IixeLG2yWFj/JxpHVYIj5S09sjY0S+VbZ
jrFwPmfs4uiX75Jzkim5PYxzJsxGa1TRGdCT+QiKA4ztp0PYc3U7ClJrETtY
qLPVlci8ZndDx4c/SXyOhmzoLccdhXepNoFOC9eVjnnL1szhSNdrBxM8vup3
g2DmFhhVVX315GrOpRj7QrmhnTIycDQXPjDTpDfem0nPiW/eviGqbdhJnCDi
Bo4LQZrt0VXAQJFWsw9rFffo0wSA5OAS8VV4XB33iUVSGpCUK5skfLFtFxto
F4BwSyhyAcmDJquev5AjQ4uv1fILmaIPYJeI+9kltP2dio9EavvfXFioq/c+
mVneZgmSSwCww+Tyk4HSrFgj/jGrH8liHRLOr07LLDk25f9xq5lQ/fHrBBwJ
l44lsbzZbOu7IfYHGsf2VDQ1fBUxfCAe4RUKQNOo1A3rjdPNW47bOo9G4Dqc
F/xB2YlnRJjXhedR1CFLFJ8d92iDlQL9PJJNvxJPVLeOB2XHWNW1AvWvC3yj
zp/aNrGnsUF/ySDJyOgsdHyO/SpBBzD/wFmF6xKC8VEVtnHfZDdh1oBhhrLT
qx4pfvzPsbyAnwCrkhDzgrv6CKfli8b565Tp9jcDYe2Y84dGZKUXC0RP9MW+
++T/stOPseArvT4Y1v6BZyCeCGNgg6tXdephLWE/EyCS5gE9t31ICElUXRXp
B8I654vQNG20lFWzfkyC7mrpnn7Ccv+CCoUQ5zGCg8hoi0H88h4i5dYzpXht
S7eXF8minGY+AL4JwnqAvFWIRd/pcOujWdwiajixwEaI4245lI/g/FVgGkQZ
+wuEjhmAG3h8mtTyZ1yZ61GgLI8z2tMWmXSQ3v05ze3iG7R4NuFM3ZhhkQK5
ECPVxC/RFK4CAP0xiGBPDSi7gyltRgR7pJLt9oLCVSjltMwQoIMKrtOJbuHk
VNv0Yo4F8MiYOA5Pyaz+BI6XtIknkEG/cj6FARnhduyFd3dgBNpsrbUFFLvZ
YRnAJ4NCezO/QLVCyggCJermhsuKYDbQjFQ2nzGFwPejenVk8y5fqttu2jJz
Q0TOPcd8K5KnMRT9gXm1hPngSXQVQVqsPm/vz6EpN44Owj34w3OB9IpDR/y2
EDEiujbWnrRv4Ls/m8PoJU4qrNcDc26HqJS4AbWYZBNG/oq143BkFmFu9s1N
TlGLZYdf7vY+TZA7oJtc9v/w5ujQjSxGp5vGXJQG/+WbM+5+oatlOsttAIkk
YnhkQzfKXUMTA6TpF2WbdO5DWv2HGRPk5cfkx/v4HZ0PzJOPRRC6AhsQmwkf
tpBm7ecng5cD5CuXsJX891uQXIUrouk+2J3LnznUvaex7OP5USveTVqyYYqi
Qg6vYRYYcJ9UAr2+kHjV3uOw33Y/ImQ/khNoDPHkKTFe7v/XaFXtH14PaekW
bsWFGL5yqmv1oV5IrgBwG7LV3XodBrzNl4nc4j1Q1d4u3fVgBtzZIZHQzS86
8UYaVGevhPtjk44BFQpj4JBXnBjbp34sSNCixpbxkR8vB1ByhRYUY6PpSLiH
XRIgv3soCCsZOo5nHUgiKlLOfhDgbcn76ONh+wFWLGk+8Wzsqv7H9Hmny3zj
57xCrcRmY4C3IhOMxth6WLPrCmyEdOY1uE7BZUPMKOnQjpxy18xVezQSYk0n
WijsdtxgjFGDFrVALkFEPTWJVeWF6EuKMVhcp4ynquEqHb1t0+05XVQ0SIwL
aAGPdr0+tmcIVJV7zcs8B+Ydlx+jpdPogAjk99IsN2aGWDguiD6tMVV9XchW
UAzese9xBGNXDkyxmOP0ccAhUC2mXb4cfzfwBFaWrw0Wqwa7pZDAXPAUU5Tz
wtr0/HSX/95vZQYObEmcAfclN2p5HLRu7oPQ3yC+DqvQn8BuaRzzm48OttnQ
61DwoYgRSc8Hgy8eG5hMI5TFDPgAMsf8BfWWDybZwU6bCCl3BQpDeiDOKlv1
HTAT5VzWdsWw9GWw9B61/pqjh8OUxoPYabk8tJpF3UNTS1ThM3VEuFkmW/z8
iTFNKOzIY29SucvBvWSC4Mo6lkmNuf5Zp+yZGW2EH2MX2yHVUQYrbYeLdj3G
MYyE4lVsB0e8JM8FdK8H4hX3GMY23ESqj5JWuVy72pzLtp1XgGX3I8q+RBXx
+M+D5sZoRBFDdI6YyIC7ftLTrdu0GdabMyxD7OO4zX9ZYLfxWeQSR7EK9v5v
h43qL/Lt49canHi/Xtjd7ol4lIV5f+RdxMTC9G+7vFBlZd2VPTa4ll3CRvTb
uRavJPb4hanaqkLJcq+8OMBiZLQQ45q3m9Em+D0zMr0ZOMvU44ecbIrrDMLu
ZXUu3kJcvrEOsuYw4J8sH8ZYZEHiJ+YZqP/ZfdbosU+NeKW51oFNEWzHbRih
Yu8a5yJcF9wxg09iqihX5PvWYHiZp1w1DbAdYbwD6FOawNSV0NQAtjfssEt4
qdLUD3Ie/5t3VHdE1PvxmbYZAugN0vdky4Ygfm2Ku9mMNVYVmZy7WICjLXCy
JhO+l6BQgDI2ozS3jh0DJ+Xth0Ys5JNVfmCL9WG2YppQRAX9LIigkt2cFouD
uoyS0Uu+4Gsa+aauzZXD/C7sc05ZW0ZgIh5abjltgjmv655ETBKm9snRLzgS
dWzFQ7feRrn81BajC2waY3v6SWFzXjKhj/nhqjo3ESZK5UCFZ5mdsMtzwG3n
+tq3lJeGlXJRQKREqiTeo5wwmzp8WMlJhvvpJxQlZYL6KnfO7W1oz+Ngc9ZV
QdobE9zntmO0IRO8Yla+n66K6ovCYL34k8VoBzNHhf70rLw3cvt98rkXgDxv
ULBjkcR4xTSIsIJgRGKJTHcTOnpE+3bf8GIBfCtMdffbE03UIsSsSvbmzsMl
HNusKBy0ov2YzKLfLxzBVHQD1BSc5qhxrd5JRhbtDY8lkwXyK2cpyG9ttzmN
UNiNJnegHpDtFTvnsowV5gLsJIwat7jqyogrl+MfaBY3kUMRnSLWlW85xK37
Cjwkn8p8mNEUxuNwQ8n6e1NokGOrhCCPvjs4YVTPPHDc9qvbgPloEYPMD7JD
/pHlwJ5KRqjMuqYxuzlyE8cw2sI5iRj+GZrwPuwtABcnPjgmbRUVQ2iWdzT8
iCzYWttDNkNHU6LDDnbswKkBnnu0YzhIehK6+Q4jsUykixKvNPZS3ocxSdNX
rcAqTNjDGR19AKBCDoM0jWeWj5dgMTzbMMS2iu/MVsEcipRU0a4jost+p0jC
Nu65CtM/aD+yEvbReB3eERZRGXGvNHXJiXq8ovHX5ZPMp5UOq9dALhJwf1gb
u+xhfAThFIZ7UvJFVuI9mKVwZM2uOk+JSheceiJ99cEaEoBKDzC+kTvyHJcz
JPV6pXI1jFnD1tZz4sSlxpNEjz0/SKT94Ixoa+U2mj9iT7+XL4iX8fpI+5n/
+nZ7hF1hBcZHrgtYzgusl0pro4M/Xn2N7zsgRyLF6WnaYWpieahP0ornp2ap
IZHPdu3pQrCOK69AJxaoTvDHi5yhjQ68V8fUBbKtD8l+cAy25W9109XnKzN1
En8wPx3wTaO07uhdNAYwwchFR1v1uWMJo9xwkjZ8HGWAC818HD3kP5hbMQiD
5vR2rp9rx6wOEHjvAgUW/MnVTAWVDXn4XdLV4C36CROK7Ljb6b31uotHdbN5
ph+qI0/+d/YstYNvrjAxRppHZ+MxyI5QRC703i9tqhhZ4l9Yx30gZd51fN7O
6WKyxWUH1/ut9zj+yl9r1TtFgGdR+WOxOehMWl7Edvx3gu84dGJ6DpNJP1+G
VkChjD2nZtyj0cDu/Qp6bKz0y5RM+LBuzU8n9+QsozX4LwhGwl2pSyS+H7Cb
mntl3O92E+j+6sHvkqThmfrJcPhTr71u1jkTYYHllE1o1So+NooC/lw94NzR
+WcxNMdWIkF+Nk+L7BR9ivGFvxLq5cWbeR8xWx+V/C9aXkpBneNZUwXiTRuC
F4E9OSbxqM4sA6eKXIzObMI8bRYcc0vfuJjx24WOcsBD07LiFE8mlGg0zKI5
33o8aSRJ1v7kYjQfGqUwhdBolGKq/iVKl9sSTOqg7bhX3r533SB+o9q7U4Jp
oA1FSWhTT1dVQnm3P6vTi4vHGv+HWkNVlmueTOu+wGYljHZkCXM/fAxFKKsG
hBPg4dGiGan0jBCK+22cm2qzc3TcDnSnBRq/cZ0W9oSIbMUabG6DHISSvWvu
UZh+v0uCq4t40t9W8meEErB42Q2GHg36KV9e0vZnyueZ4lcrB1RA7GceUgG8
KOi5HjQUIxvOazAFHZGGTI/wQkENd8YP8GeBXjmRKDYgLosDyToXsJdo7PfD
YK3ym741XNxezii35RuIDtwCW1a8bMxdkFQuKVsU201HxfbVjLMnwNQd/LGJ
Pu26z/Y1kwx5Ex7kWEoMQNxgZfZPfs6HlyACyF/e/tOYgmd1onjqc4HOlRDZ
E9pYirVIfPK8JnXNAiAl8jITEkCLBJSdq5H/uwLxI9JhljgYaEeYzeTwzr3f
mLrJy2PMcUhS+rdx+DnjtL0gNAYVJgwPsNTU523dz9pCpeV4o2hFzi/srCZX
EXF5/fSjXUmacV73DN8j0d/v4A1J0UCElYbEqAObQv0QrBPevfJAztpZdVxO
pDeAkR2P//ELJA2g5VcFMU92WIxOO+p2hifSK/Spg/ZGLBqdkKqAPMQr01EJ
4uulXgwbTokDJ25vaSPTXOIuuJp8fiJDgWF6fxFFOI/J3uO4/4UnEvmA36Xn
BF311HqFQQYQVCvwcvzHHaf5Swj9sA/uo25SEOWo9DXHRNyC6BuY04iLGqqs
bKpj9jt1ZlfqimFTa61MCVXrfLMa3ja0dvfr+RsmuwznehkX92WEqqrJxDmu
NiQX5PcfIqd2qU8npnAbjr9xhnqa9NzGe/3zYX43anCSE4b3M72qB7+k6dZR
49EOh8Zwe2z/CnzqWchb7pydFRsxJpJj552iOboBi+y4MzeoGgV9gmhQJSHO
CSFQKZqXHtE0eYWG4cQO+GRaLyyKLlqyfVwYlq+jLMY723mqECQZVNL4I8m/
HzGrWbVRBHlbTb4qGQomCXE4vjoNa5jDFVvu8SEVw8DQWgXsotu7zsywErjs
IlPzy3TSl3qsYG0+zbuMGJV0eUETBmiwpNamJYJxXL+JaIhWRcIHKoKV/So9
41pKCkRXJkcv7VigOKiRW6B5meC9j90u9Cy6zNcwHETwf3RYF9Y6qICSMChd
OLgFR0trIbXr427HFP4ZgW8oIjgWJL+lw/hYGG5yxIYvbU2wltaU5l8WT8iQ
mdG2aXQdybBdIwd2EJAGTeEaUm235WxekjM1rqu6QZAMbR43uKQKCI2bcMN9
dvpqLlhuddqBXlRkgGaxlhwCotB4AAQ6qh7BDwUqagCre+FAAvk0wnutirqS
+mdPLv2z39+W7a/GWiwfJWiyxzFKU5jNHneg+PIkdCJsOHlZoE42rzA3UaBW
TR5NxA+Uj1NZfwdG4l6nBSgDEWDgdNvsDxmn15AMjNHxwy42namEV1u39Of2
0wZykkNPbM+nDWrJIXGR64C313waMkM21I64NL21n63RrJt/n8dAO5eh68cs
+S/m1+/cW3VGFEx78DQwC7A3SSWuV+SzpDrG7YhQ/YVwT+PPbUFPC1UkTMiO
wbwbfUeqlIrI1Qq5peQxCa91dL61OxRL8sO9whVf3qeEz2UjxwYCJZLT4WkE
zSM9MUFk/dwR/Lnx7yJ0a4riDN2aadDadk8fH+Fne3jz+V/lqsjGlw2T1cwD
aPG+5SGSbViOp2PGHAmyazJIagAGW5nMNu2ptT+gKX51Uey6e1ZwwCykUycW
WLF7SBU2yKcvNfNB6htkZQCNx+5X2TrPS5JhlG8kZ8GozPRH/0mkEFioJR6d
allilmwLPo1/2Q3U3hM+wI6P8olkJ7wtJF9Tc+SarJPKp2cgon3qb5QlgUPW
Borpl14qkkoj8d0L7YeJ/LKStdjA23KmG6ZC7xnrRySMl8jSNZd1fzjub90F
8ANJdk6aaVqeFqm9UsAEfBcakveDaav1wsnen2FCmzeHwwiO9k3QbS/IbrR8
cNbXJbhjoQv64rX+7mOlFwgyt0zfennNvClDnyGCKLroxg0vIMP+bgvw0h39
qGI1T0sXCWwj3nJ1+jGl9VU8GgWneHiaFCG03o3Hz9+bmlULmG6fxcI7obgn
SvHZkw+odApOdybFxtJm1ZIbwi6ZVr21/RA3EoeK34P8vDMH25kcoWbSTcII
ryl4WjZmsotg+Twk0Yd2xnI+CWc0yQ/lOe4enuBrmAUtT5sPCioMFB6y7H8m
YX/LsZlQekAgWnEMG9H+QVOauoOwQkyK3vQpSrI1Jf0hP3HhhZQd/N9jrb1D
pC2h7VcqO8m19MQD8BqG88+zZap8MdEMU8izx3G+cTbIUL9j2U0xjytwXoP1
fl9GsN1ZxE3+L16Gtnxg3amhIuAl43CXwiGc7WELG+S0CXrgCB+zMcOdY1ds
JKcflZnhwbjes2TCGm1yiXZtBdhwcv3O7KqwyXu1L/mvXjLyJWzoolwrSKlX
1SlPPAirA1FutTjIfVabKd3p8eQcLzUSCdrnF6ZxonwQ0+rWrj+abjpt9r/W
4FzXBXvfUHZSZiVxn+S7vjR5jHKUFyTj/Wccfl2tNCgyFL9xOgrqiXta5TIC
Xb3eyFdA2npIazqcG7sAyz6/ObO0MStLGM9UHDRmkbxIytp/DSIK9OxfE6Tk
Ph0x/ceEDZBzsFVfokVaTEcDOgmRFx/lX8DadL2cd9vfqZEDo12XObMuikG+
2RrggEWL7JOZ2mCPGqlyM58OM9hCqxSOel/u+XQaj2SMPvVI2HprStIsT+RF
Gm+e+I2n2WBw0NUnK3HPH1ZqGOZMKeDl0PrWq/FDu61tXClri6CUobHhBayS
bvimR+GA2Ry+L9wnmDxnT+RzMiGSgZEtV+KJHxznBOXFFAIjOzvYPX34Yy+d
fU82P6eIcNPX1WlbjqhxsBdGEOAmIZckFteLxU0i59tsecL+SEV4AlUD+Znp
ZaFYkx0jrNPaFnRN2ywUYYMYVPalfl06yqXf9Zn841F3kc+YdLa+15h5FOfh
SL9iS32dBW8EM8hfqub3qPFQ7IZg7Rpvo75fSTkgfI+QwgN3mRr1Tu+V+E7Q
9FWr1tNPEhDUKC6JpRH4CqylTUKFSW4oZTmRc36wy1Zje8PUlPeQc5wc2eBh
qmSzmYW7Yk4ZWj08ZUs9D1HcAnA48hYtUkgnaSquamU6k88YMFPBK7XOWGX9
Kl2CWaCZiNYtS170pfLeG2u9TA8ZdqIGR6P0XYNQEhJD6QP9uH1yACDX4/Xw
7zCyGeHt191mXUacG2LTanZf1JKNFYCdctgPNbQfpNKGvdxQmYPhGGTffiSS
TunL4OmIfYS5qhz6FeEZbz5Fctp7rR4UKnGxWJzwfGVOWLAmm5s7CcGLbIav
//E2Hro4rAk8/l8EvKIQxE2aeRyd/2+jKIsgdp+6S1pWAlYfHBDrFO/aP+l2
fvSRfDhRL1MiOm9fzR6fLrbUTwzaKRGrb+b+Dlcvq2X/Xs8sOWcXr/2/S5lm
aTuAQ8zC8fXveMkthmgInOk2a/Ztg32Y5mrTYBJgytIq2h3CA9kn4S5yH4e8
64hBVpvJymUO1v1tW1u7UxrwUfziA6c6k/Jzeb97g0e8c78/f0saQOY6TUZ8
gVKx/qdU9kjv9+QZFIlX2NUQ9uYnHw0w1tS2T1fEpBFadtRFpTfC7sHtkRIi
nrThAa0zJ8TM1Uj/971at7aackmk99z3eZhDK/VxTAnttsgkrakIN+lm38z/
3pZURoTL6CCeY76Tdd2tu6BJelcBbehMIwQtKY3f10jyQo1ikvvl4rH+ZFMg
H13BXgsZtPiXg8Dg1j/sKV/8ez2f3+vnXmhJpu7Tmw1mJ5w7LouB+fa+LoS7
N+/ZsI+nq3W1Z1wNh3IboLAJjyPbgVTmBP4/LvPBusEOFseegGMfeb5hCsiy
xned1dSoyxAwNGCJjvqkMlQ+fcH0DY+Rvxd55JnvU3VZm62KUkHZRXQpwogO
8yip2QhZn3SQs+qNpUqY5nE+j2gbWoPXKCBeoSnrsYqzJXfXGMKhYaSx3xrT
zXrpQZVesJDvpVxsNHCRpG4wSJEamcnnGlEOINtvWjKWxTiFl0rcN3YSGb/V
26sCXB2TQCVTB7y5ufGgBBkTQwQR9G08eFbDFk4nOVP2eHcrgNesTCyvEvMw
MPsh7iNnHe8bJZVxeUR+tZ8Wu7BCKW2klbKmfcMOVtePqipX5fJ6D+t2t7wV
3wpqq5TqSmUkClCwGbyvQHwTTfbY+z1r4BEBUZ1NLaGfC4FO8r7PoGX7/gyS
PDH5PWS5U340bZzUPruD84vZvOGBienLEOxfCTc9LP6lvVDhGWUaVG71c/Rh
RIl0XDvjQcjpnw3IZ9K5blnSOmnhZynPrLHyBlT1R9mTaOGMA1EYgVkGWd/t
2EKV0VFTp8O37YY5Ek7j7WE4yfwAJ9JTW6eyjvxOhH+SxkAj7/NPwZfomlCf
CFJwIAWDEJ38+pYacPfJuNEb7FC/1LDUY/KnH+HoAKEovNsNBc8Jc5VdlR38
rC3TgNgtXSz0HGuDxyFc5P/zbQW4xYYbRIQWmebQkNVYr+m4e8/dX1+5irhP
bVqSdkrWEmyayUmo7jtDqSf6s7XVXBJzAdKOPlhhwsLFNeHFvzLmNNzPKamG
dUY/8w6E+Gk4eG94khjFIEN6mmppa4ene9N0PDm1d01BYwV2m4utwyFAotPz
iYkYJSN+RPCcDhsA0bi9bhZeH4WutAWmdprav0DttMtpSScCRxhkqIEt3PhT
fFL11ream2d9E8Zlqxcg2ZqHTYRKBMyccQvXZTZT2gk4GCEX/2u2tr9/Hjap
Y/QvRQ5POb0SudMMjXWLqwd2tqu7LQcN8Av9vev8HSEBbnTkJO7k9+4LgTeT
YARheAvhQ7k8iq8BPHd+4UpUwdcV/JFh0Uctf/MfLh7J0KjJbWiC0PN3/Tnk
KDhzkBC/VctvUPHXj28WuYpa7sMXtgoqw6lzzGMc1pbrLnv9DCuU/jjeohLw
V16kdjcQPGSdADOEkkKc47WCQLK5HjtxZmb/5hVrJnq9LQ6nGG06Je3vm7YE
+66pz4bQWLBafJWlgs+7EH4GCcY1Fis7Daa64vSS3CncLtu4NNFOwa7PHLTy
kmQmOTPaNn17Puw8mZzG3JUkhbLEd3COw4cEByNaHVkwq3sHkvXL6ysfEteJ
WXwqNen7l2cDKLv1JTz/uRZxGY/pE08gpe8Xxx//Z70FvCABK23nESu7UaPk
f3FLDNu2z2FwwI3Vy1lZbYl4hhzJtMpEmj3D2aaUAPcAv1/YzQIAne6a+t5V
oBBISI0E84Ui5lk2olCIDF6Bdxc2TWJFLK2ipEou3uVXNKTRjC7EJK1nUl8W
6o19ywOE6+nQjeOAwrG4MF8NGWfIJGntnXlW5evWBzRxJtH4JKMfPkL1VOnT
MobwB5imKz9p4lHL+ygQ6Fh8JbZDcTa7dL3rXVEmNoUI2vRCpyK0Go+IysRv
W9XvMMNSmQ6PjT+tdzZZEJDObziP8uS/hVOANa+1cMbqRUUR22G+rcMEilC8
6ajGo2wYFAENVEAoAdjqoewKo3kT8qnUrXxwUhybqjHXGlEVhxl9LTR/UjpD
cUJU4A3HAwvGwcL0UK5glbu9kOvXXQAcWanIcw7mWzAOduJxFBa9mJBT6oFq
HQcLQciKfHxUdCWlv6y5M40yB585IAcXSCp5jLqUBTvoKJthnDVXd/gMnWmk
32zbBXTZg/wjb/n1fbs/UbYJFDGHFH5gbMyYaO5vpf1OTCPpd42XM+709J61
9o7CZjr1h3DOdJxC7t/hyCwCDGp0vEtdAlFxW9uSJkVeUOuWkmOxNJSlLfxn
5e0+1KGoI77++J9ilyCEDSUrf7hyqcDW6u9/bXRlUtdIWOEmopQIPVoDwJRn
JOJB+T4i/S2hj5puA5FehGzYrtfTxSsXMv4QbejSmQ4ddqhZC4n/v4aTpNJF
fxq+J0jSybBwaP4B+5dIIQPmumjs05cyH15aikjgO/MNcoVBZF3c4Tm5NJWB
VcP3YWIWvMw29q2YskzeEmgPw2PYT+cgnjt6+XEySKu4hubuM6xP44iSK3FY
50XOD5mZh5ZweUaLbkPMACvknUEQfnda3XbBNkr98b3fWd230XgKnOfJg2PZ
zKBruFD19wMSkQx49e12J0xNCKJ+pfmHpyyNGv2TPyUJ2TFRrKVGuJGoM5h4
V/XnE/pGPTKdCHJLIvWjGjvCWJGf/HnNFjTeiWLxVBH8Q8bk13VP7hxMzRhR
99NBWDSz14CwyhdNVSBxBCxRjwS0b/TisbPBmVdUuUHBfKmH26prpiw2lsPb
8oe5K95ENvuZCF2jCjZpJFtwLOxL9G8FC2nuqW+lqzWobC956FET6NghqG8I
o6MwV7/IelAGwhz4/artx46zLF0JD14OX1BzTyvsSEMBoQa9id5ofcsCx4Ye
emoTGjOt1XGWMvAFwDYKEKF7toHYE9bL6jDkp4uWJPlHwsFwKZEC6BsRu3r3
OOqASZBJphLytq8wQbS1zsyYWWhMiaJxTfqf7y8tvLiGQA8fyq9m4nz7156d
rQEsHYdOUv5EiwCNwoO1twPePtq4mBCDYf5UnCfZyN29YB5chC2d5FJvgTBA
iTrQmO83Ww/7BgqRuD7rVpsKFuTN37A4p0lsrL5mM2wWpsgPJb8KHtR3MuLA
DGM+cJKkOQmaD7n0gtGboNIrk4A6B2nzI4dLaBYgDaQB3lu038QKQXT/eQ2G
pdInyeqwCDL34GbiM5Kb6X6Sc1uQtyfWsufIH70AeLZ0eRFIJ5XPBtCnts7z
EpM9gf0P1xxh487XmPbwV09fj+aqe4wkdFON9NLwN+PXpgfmL8m+LDlX38aN
O5voFt9I1nlmtME1Y4vND638qpsdxU5YiHWV6Dj8KmFC9D5u+NmciivclJFY
3K3Lr9k/5VRMERtqRWh/VzIb2MyMx0Ncf+WjTfDJFeQNvfI+TUgrDSJIp9d9
XVa4TVog33uimUxun8RAOzJ2nAGX430zBi0I9IVpIQ6JHagq6GiQc82kqugz
lkavaKp1bEbkezhzFo4BJoGNVCH4CoCu5v1KSk+WBPDYyqqvX7AFti+WxObA
9sqenjKI/vqqBKFCUev7XV2vSt2xr7z0bl3XVSrDT4hCBlLvAKYr06PFHtcF
7AMjhWslqgg7Of4LRc4WG0ibPZwJdQtv4Jyp47TopvsHzxcW9GVWdAr5PyIy
u0rfH22eoxGP259n588cbQSWppw8Ff2SkTIMisoYUg3wT0QDF+assYorFiZf
1ZMe0BtZqNE8LUfuZ6rRjkgxXsoPR1Iba5NY8NiE5qXU1GcnY0ozJKIlZE5O
mTch8CQ+AKy5bRvaarXZeBMt5/gmtbO+MDuTlQhF2ioqsiOJj4hlk5alw74D
PfDBsb/iDC1UMPGnT6TBf4uyJdXLGQixvO7UAC8qX0YrxEmxV3P1Gdw2J92g
Ttd9LSzoCnHjbF4ZipQ1syy7cuuFFNvXJbEW9z0hrX9b7hViM2u73g6FqXsU
NgTwvgyZ9DUN03t46TyDIDS5lAIt9XmVgf0kYqECtz6/JArXTQQnzMkhqJ3i
ipTkKhYOqBHM+WvhMKVxOwMmdLPOrqZ4kQpso3124huUds2dd/VL8eyGsUpi
FGc7dgNa77zBldQ6nfJxGfARfVM0u6hemPe+aPK9ful3sGp6qPWY56Bs85G4
HIyZg/CyQ865izrWCLYriySY44lRx6vK4iWTfWCSPOVQ4rO2ihERZw1dwXbU
EUdSyPR40NyGDJTgi0ag8UlPFrImVzMEQqg2ozjgid1fkAe+UNDbHXXLAt2b
vu02ae3bAn0yb+B3+yUnqM+VeXxyFvdgbpt2wDZaFkPcNFwP2npaHnaQ3L6w
lVd6KSmnlk8d8GlzCzw59QpyRoND+wN7wR6zObOkEUOM/dqD5o1TEpXH3Dqk
F/Uzw/gIUpodYOHkfuXrK8XSU32H09SxYajGZ2nT3uUe/W7Vbr3ejYO0sCsA
JpLJX8ANjiYR6LF6imBz8115iQRcVwg6QUtbxNzGM7JOpUB8VrbUpZ5+Xqd+
5nYNJ7FIMwL1FL0ioc7D9SQSU5/nUqVVca0D0gcG1IskDUGfqAUJUbKEEF3Y
Aa+xunaAKv1iOXPNMfSP4oYIOHTf00W87tejTmhwWzl7gDYjelxu7I+3O8YO
KKWVVKYf/WB0eeeZYncOsymObjMro6hQYq6aneGWYc38Xo2ZJB/aSEULeXPJ
SGEeOVlj5XR1tW7g5qILFV12GnNgO84YCZkwmpfWqFgEPgAdsYnx0WAuiYnk
N/nJ8HJy1vHdh4lNzgFgkduFBknQhoTt/JOrQrss7pkhs9iVP+v2yPEXckPu
tA50D5dXhfL+xtSOj7D0xZW8eRPE3NMZG1AZQfIdO/zwajiLZ7rNAGFJz54l
D7jWTA3Jz4+w1pzYpsBY3BYGAcx2ADW64rUVrw4zl7GZUWl3CG+gVhTcH62R
yyjAY16VhTfUfUzeaCTWXF2A2FcAug7Gzs2wRAukBHC4jPqzQp2jF0KQmXWf
dW31EZGEmPtMFP2ULjBFF3QQpv/OvVK1XSAAJMVGNavyJX+0npgwrOiVGiXJ
Xa5SDE/yFsOjDMr3cxJsH4m7WOOM2/hl4WVZmphGuw9hCCHnYUcw/alFHjI2
nsiwhZd0o9w5t0IyuhKuj6qYaIU0f6gAXn9dGsZJBAnon/zm66EJxLvdHEUb
SIS0VZtLUWtyQeU3NrlFBmFTYYs9brNVTRLYW12mqlL0R43PF81eUBboI8CE
zipfoQeEeoUKmAJCtY2dSOuUD+2wcmulNWT6SWSupuq+jpKx1W5m872atJP6
0eeawFfBZpNOiR6wXLKpKz7/VXIIqXp9R0Pc01ZWl5XTJLmqfBVtLYhMVhzO
zfjOwWcrLWgVyWFJ0Wu+pfyDgt6LtDT1CGiaYzJGWnvU7Pi3b5j6UdjwVIFd
/HGjqen5R8nYYArbkFC8nRgMqEquaX+buaohwjPBjWfjJxU8pPvj/o8jJ1H3
pWD4NA1H3X4fN/DiN/veuuEMrTl+29/KfF40cpwVZDb3eFcansAyU/1BoTXX
D3+3w45SvUBO/wzs1/6+B9FBgGORdNTkjqDlYz5rlPMLjAL/yoHa+LgXEYHW
27gjIB9hgVWw3q1LxeVXJhShv/jy2Ac0df8HoibwwqyHQqPnr0UPQ5AJoUkL
vVcFjSl50YhxLB5dKjWssivkfepQbj6wskDDySw0BusG+QKbSGJExrKbP5GY
Nrbl38A+BQr3cyI802nKm6TJLVnxd+7X5xA9C1LcsnMjuLLf9Z0wKJl1j3r6
u+ZkydhDLLe2ra9yqFi4/HSGUwJF8SZLG5/BTjVrysDCcPcNrpFecJgohR9C
/zO5YqLWz6UGsa5XOxpSajfrbe3usETqnP8qo7WexExLrPWv7J5Ggq2mwBrG
4FD3999Mm9qzQ4t5P7gzRexD29hl+dQmWLjR61sIUZSq0ibrQ99qEOSHnn/2
hVAFczljsuBiHpWTIv30AWzpHYe1MnhfHJyoYxXW0HZvokmSZ08PFtzQWoKB
xcaDUa+Eg2SLx6vnpQ9IF7K8gpuaHIIDVpd5Jyo0Rv9RDmkoCrTyhyQeC6M1
UnQs12eHx2I6rQN2fGyhzubuXoYeBstuijdHkCtcnL8EHp08mrxhJ14i9jnY
Xt3sMXhzYzfW7IWwSoDzJiBGZzfrdzEcOsHJ6X8Xw1TtZn6xSfDO9T8KHjHc
WDzRS11NEJkdqFgG3LeNujEiARMDg5G0teobv7SWLKnZavSOFAJCPpJKXuer
maMU6i1jUAkrtWyphykByfjkXqiyBpaNUeLIQrVZGjn9NRkNKj7ekZqGeosE
t8o4+DkLc7K7yxQLZ5zCD/2jlwZkSqkLBT7NzsxoGegVNzlvB4xRn3CPbKnZ
iWPfMs0ASfmFOKsPImQywjHXxjivN+fjxyhgdNUYzr8gJ9yjFBxbzNokzalk
F/o1RYNyU/E8527sc8/5i4OhcgbfwaR2jXz24qfaNdpgJxYpVL5tcOBTUv4U
PH1ie8bMrR2+xe+zR0rEtrdDmCBD/2w3VcRP7rETHIpL0P9clTRj6ITmsMXi
cDHWlJmGQKRMvtGFBSheeYvb0wrU+WvG8VP/FRPFfGVXGhdi4SqXV/3jrzDm
Q0FMhJkDt258a/3ZOHUOt4JhgEEUFp+4PDq1SrNcPJJ2yWQY5QlVYuDgADpR
xKr6jee9196o85HUUGi75Rw8jSapsfAJVEzGabyTpiJdaQh3ocx77SJiJS9k
i5Q7R53PcNGT5SAF1j0KhlJgESldGI4Ae1Q9amD/tD7ryeUDOkwdoyBVhJmU
vqorA8JtvtkQuJ2kIwQIYZct5gzqtThhgyb/sXic1jGos184ydCmpLDrFeT/
n20m1+f9e1WWMBtoyeWsLv51DC+Df682lxbiBue8VT8GQueHrsoj/O2Oy7OQ
z4EdEKWk6+AWVWMkBTvxjy9lDQCeKwzXP1cUaoaBO8C4fMsUP7Whvg7ClohG
NY07av+Uqtn8Kj4ZDuBcs5X8Ms5VNa4tQ3/jKWFs5Osrojk+DifNL8zkxp0+
ehjiqqvdEor0hGWiqBqVEF2vW+u8HZs3JJAKInfz9hYQy9AQXprVKEZ69/ek
iBI5/vUZl+9hZObK9TzoHC0KyexzBJg2pd62Kol2akWI7ThLwa5OXBLhwq83
D/9PS1waf9uTt+nw4GARlblWVwMd/bYvE6IfpNTo+C9PeyPJuCJEmRgRY1ku
gk8MWAwfJ9CeLKnIcBWkD1VO5FuefczT34LX7LHqOiwTvSfuEv0Tby/mqTVD
WhToRWQYfb6jnZZ6HP9hLeYxlT5XpSQU0u0gYTI4als7HcPgYT479zxZOSR7
1FNIT5JmmWBmml+r2QhdUb516x1E5tWQf1RjIpTuzEOxtoGsjqXb5+iafdTV
DtkGQY1VAsSywz2P5/k5jZcZQC5zYts8Untc50zcELCvQJqT5zAx2WmQfkEM
pI+VEZrIAIf4bQ0kedASXW38aNq0yawp3w+j6VA+njPGi21wcGwuySAmEhaR
B53N13VSEbG/QSTzbGlyqu2KVZXAz+Iq2xva4IHEu1RT7WtEOiz5Bfttd18e
+/mAHNy3IZ9r2MMPwZelpXeSV8KR96M46iIczs+LfD/X+vAYX/znd/dBKQo1
WfKiB7s+kJywIxpJcBsJT0qOfrkBOpwjnLWCy3RHRRPRoPIJfGtE7QuJVz43
vc2YJffmJ7WExeXI15ErJtrztSqEcrvn7307V2qhK042uZgflBn5ciy63Swv
9YXvRMSTgYK4mANxrBl8xctX0IQnvzSf8eF1T/TvU3kAu5ZtG9QvzZg2bdSr
tv4Swga5s+uFg7jSrBitMh2nXYFxB6xC3Y4CeuLV27JaQNfAUMtbU35M2fer
R2mGnlS0nPxsVzm8YX/hHcTdYH9gIZ4Bcx8In05TMqKh9JGRqGoTf/ofeRii
VMTNQjb60gK01Mym0j2iQNQQuu89S/SbCWXxRRjTiM78Z0O7JELj5X4hRAwP
rlLr7C1Jl0Zkkt/PYulyvg+RwAbv0oUlK2sIHhYcuk/nCGHBe3wA6YCG+7Oc
yowNf9r/jAr4pAyqQoCVQbeh+X8gx+g5HwDLG8DFhjEKSzixyzustQnsSRTd
DiM5EuaerpEpl0qQJRO9/IPO8X09nApfeILTo5B84dlom/66mDXyT0/+7jga
S5wv3/Yz2SIBGkxF1Bp7RFMbro6Gj3itrYYgqpN14xz/okNC9BrtLbITW9lL
e+L+WuczwnrmvqNNTtXU1Nk69maxv0wbKEpq4+gy3v/OFnsbknX9559Gf4iq
AApW0wu/UzTiu1OcX8oUdnuIR9nWvcsjJdJmD8mAhPDggKMapbtxVOrWLJW5
0xsSOlRqTHKUDvSarQWjTXjl7BeF6DFkNXPtQ/BU6nvBHmn4RSx491dZQAcN
5Bg+sGaULVgmR/yv85WTrE1ogVcnkFLnGhiJ9Gay0IZP9oBK5/VwkCrDVXoX
or94HGNESOgH8wYmgUu2AyfvCdPrNXFB2GVSkFzxgKU5QWEc8CqkxhDlBYho
5yg2ogQ45giEEwywepSXvgAiRk83K1+Fed6HjkSgof4YShiMaZU9mRA6GGey
gAKlkhSlTN7m9zCHOOH1XjDvE9cKpPHRbyEIrZaEVbFoZQmvve85C1KKvX05
Nzti4MpagUo/Io3YN26GVArstLLdS9aBZfBT59+PtTerQwF71rmiI/4dUI0d
vv58AHi4DUbSM9iXKg1CtdDZxyeSVRgW9y2HjtNhEAbKTbj1Lck2JnnpLSq0
249Axq6yXG0MzoO8oYih5026UVQtWOLlAy61EUfgHfdQkHym1JabVuvlFEwm
gUMALfqJ0iyxkqwUTPhK72UNafJpazLvv5393cGMYzadds+1U5t8vGrpaJwr
1iA5Lb3dKgvosZV1epP0lsMBobqtRJWBZo4vFcwKR1Eb0Jn5waRwta27RuSv
VOVjPiCoAlqTcdo7u4GROb2zslNbi3097K2sNxNc1Y5ZV90ygrVgz1FmyR46
TAw1WqBZpcTwbJE+arIMoj/iFQy5qJbbBMRHRCfT2xNvVhIs9mZXJdSvyoGJ
amNgLzzcEXfMc8ytYrV4AtMxdR1HdZu6X4S7WAmzUe2cuVT4aR7bI9NUZcD5
9aW1bYOt0+AphjDmOa6J7wTm41/vSpyd8D5s7kKgNMuvSwXzbEEXAf3KMNvM
2Cg7Y50rjLynTn6B2WoHySJkgCDIuhWR1e1owbqTDzv7h/P8eO6YnBZFI0cA
yV3Qo5Ucd/t7lQhLkSgWSIWkGSHJmdJEbhjbnSR97tNOV60GcUY919ZPiE7i
HZvItg6rvveRYpiJ5aDnQBn5VJyaGDgXX4RXJ7CyDaHnjQOUEYCIG9W11PqN
+RtBgTYnN/62gtVCxjL3yr96n5lA6CtApnVdQoTqr6XpxW/EN2yjYUk4N96G
v4rR8ajV0bPRw7wGK+gqrwNbANImDZIUWkANAIptG/rH+m+SliA4UEhv66ml
4OIzja+gH2Itx4AU88mjoZyp5ozpH1jmMoRiveB+i8CcDoWY8xZgLU7izkI6
xHPzxpYuqITmusB8MsmlfclIMW4cCBWwsOfn7Cilbqdxm1s2e501Kc7cfsbv
Qq86oxRisGj/qBDESlt4JpR58kEtKfMu2AS+l4Ny5ywzEyK2GA9nex+EMzZB
C87DRsHaw1lxvHwb2WbdU135ACyi8e3UeTOQ1r04enD1jkRw1xoizXU4TPMR
0QECzqYriHzbCLo2FGq/K9cWs8eJIoN3yn2OHED7hKulD+HXpFz1j8M3bVub
UpDMEWFBwfQhpXdu/myEQOK+So5FXVuIaExdFMA7HG8Hb5SM82cHrVe6wZhM
og+tLM1pxPsMzxKHQad+wbppW6AGq/GNMQZk6Fue4ofz9uie8230XOGhAjVz
SYb3a9J8Ogcf83MEEgEH/8gJ0nIVNQicb9RASkTMDCGLStKjDj1B3HUgeZI3
QO6bblghnb20M07H2gKWL3aQ8DoRaPy3efOdc0Lh6RhrV5a+4gqs6Sv+10DU
Zy4awVA6IUw0EoIOcPYYQTjLq2oPDrrHh1+9+Dgh9RWy09U1xnbq9wKov6hi
JSw9wxH45r4EgqejZNluVoBDMJUwTAAGwdgcp++/jTHSlVFHkJk4BaMNeu9q
IqtFthVnnLHi/bD/MoupJX/PmhkQhOLjrUsjdORNLOGUESoBUDL7KUcxK3xc
wSz99v682bArCrt8h6a+VNL/YnHYX03NS6tOXN/X3Gn5WbhFRk+ci/KRqNUb
fWSYityNgGxCxcYacX2/R6d+jfmRUv+EU1qQG0TRRzJ6yZ3p5U9TmDx45O08
CfrGTk5spX10E72ti3UWwktiI7FmaM1Hrtld2gI9BZ9WuL8ynVu+Ndq6WTX+
+ML6swLNf7V57dF5ZLbiiNE9mwsTWn5XceJu5hSqlt5VVZJb/kAoomzx+JPM
knOEO0koNOSuWVnaGND6zR02uzq8f3DugMAJEH9z90M7pl8ULNUMpKRRwbrY
rmkpujT4X9osyZMju9tIHxum4eNZhHgW9vNAyLKGbIzoZah/IC1H5h+7+WFj
iOpQlWpsJ9AcwmXjgfMm9m1QhxnhlhnpS8Ht4tmN7klSuWJMSds4sdomRcSv
cBbastHFfoIG0gxDD4gC4LKKNAt2wBUVEY8ApZjtnrNgHoWkEbTNeVry76Ew
3ifHukeEFgVFV8ETgS6HlxxJRBw3VTINQVJzT6yiSj48a9f8f60SXv8InwWw
kWUpk7HuFTnOfxG6Y92X18H3K2fLa5rJ0VNx/9HgXFKGw+91mcrlRftvf2up
Wek2EFsUGWCUGoEpPNJye7/BU3hFyPh73y1cUxKULggTIV+eotAI8VeOq2yP
SjNxRcZH7OcCzWbvgdYpEeLLntEPDjylL0kD4z+QLInb08ewavpWb+hs5fgt
hHcXHFduQ9hfUFmQlaM20zRkzOAdoiZAhTaxh4xGjhE1EqeKeBxipuzRMMxk
XQvqFoLG5dePfmv0RaNk6p/gHTUirehxcKbF0Ztx8o9qo0EqnLoJLk2AfzzY
5KbH8hY5YNbnhSe35VXsczqf8Q0QHQPLkUI+rSC5zAIS9OPF1vITIhQJL5zM
JSBhQ8an9VMW0epgS2Z/S3ckQM1S79NN0uE0hKR6aOwz8cz9GydKVkBPS8UQ
MN+TZ9EuhdppRvMTz75AkMPAR+vU/IwUE9Hr8AoNGigiiT+AgwWNjRRcU7xt
mkc0F6Lr1B5bBbXHmEoj/yDOr9cfg2Y0JzphjQFxoIf8iCp6t6uhIttSoh5o
T7NJsU2luRhtbuXvKeP/ozhXdKrNoZFDv8xiwGjcwX77/ZySxTJm+C9Q53Iq
1vEn7VakhqEswZdvw3diMqhcsuU5eVYT/xebKYcpbZGQ1SzElhQUJADBx7cm
ncEQcSzDQHiG4lriN/ARpByWokXYSkM31Tuv8H8zQ3IFoL6w3GYVehMXs67y
JIqP+JtRIKrSOjGO3b4aphMbqd+IKZ91BnYrDCapC+/JMwsjMrcbcsjBpruX
i1J0Y2YvF2+cMimWKKk/4mstd0J5VUdBGikRomqwacAi3wo2aNsEuMXYEWOQ
yF4VeldbkF21Ttg7Uolbor07RErrcXvoWN1Cs71MCxmZnBrWyIKUQ8I9a/KM
OW9onWumxDcyu995z8NdbPZzuqseezNXRGRw/ntqPPCcSxscV9N6R/XeCiq7
lxO/nG8PFW9jc9u6ZGW+Co8vFUTrV5PHHyJaC/VkI6nxBSM8FwSfXUS83h9U
rmPWRiBzoIA1dFy27ZiKDxdT87HTKxKSy4CYFR0/u3gy5NBhqaHmOdNKlQL9
lXyiB0YeblgcciiRtfzyShUlPvaoFS/YTf6Ix13MqNJevBF3rUqabOkL5n3T
UshlpGEW6po3ddbF3teLudqMkw68YUHqA6bmNCkexDqt+LQchkSQnB1mQGu3
yspxBEsezwUeg0SIICakaRirRF22SJm3+CWiab7H7mb0SY3WGLv2Az1W3L3B
KiBn/cPS3OFwE29ZvMGqrAMi9OWm2MYoFVWIuk04r5adyy3GIzbPDNB8RzWf
cA8Lk+xhYH7FKGDLEb9iISHuF7SHeJVIdLVJHXVVzUt5ezeibLXLDmZR2aMu
HNQ33E51dUvd/ug40rp4XrGOxI2vo2k7kB22Piq+kLxG6OI5KVzYUNyzx9Jn
IncdrS6+fVSV6oo6AuIps+vf3Pell3spuvTubWC/LP3lOC1A6tBNyJFzLUCx
Y7FlfpVnJpOTVO5PF27UGPzYOntIKhV1rUnn1QmsV+c1Wxfu6vqE0i70tpj1
3n6a/Y43Sjn7hnRLt5X8nsW+nAEX3aBR+7VSdMYdcouGKlF7550r5wKurw06
lUxwVacVIhkxMXHC+tqgR3HaeEtS6278my3FpiljLCW5nYGISTfyJBeZ2b7m
uz0xi9O0NHj4SvHHjKRDBBA61rTxpLzeUOQU2iKWlBG+KXneeHhrh7D+MjwO
S6lVZFPwz8cTrkxWoWzEMgfWdwO4dkSzKigGFSCZEkJR9ZhwgyLMtzLYTkcL
DId7JAujoAgha3Un3GQozcxNswSkieekC4i9V1tliT2eIQGzIlHzEOorz3Og
Utal1uDjnJhnpdjrRurYRndqwP8tUUCFfdtNyfqE9yzZFP2qf3qKDjPZ0HRy
+CE3v/zXgo7xP2ctdScYNNdZnV6dnJg6vfmqX6sN8c3ZNcfr+Egm7nobP1kh
nZgt0RJdef/UwUbPFYZkHguIAVTsGn/nkx5KJMkBS1jup/JXiuIxXlzzbMyF
M5mHXT0F69+OvEc1WtB6eorCth+zrs99NCf59D6kJUjeyYGT9NEFRY2Hurm9
L0zDK5cRb+Nyop9SOOtXrEspk3em1ZiF7vi++Wbc95TvbcKz4QDMTmVMStCq
6wc8wWPSjwIm8wzjqTvQ7XllBPDCX9M/ePItbPKqs2GYIx/wt5Z9wpFk8v+Z
R5loeghyP4SMR3MpoZX5wx4ko25riO7JfegU2nXIVSrneq4XwF5TrcKMjKHI
kbCdYhmCWvu2rEoe2sPaIq4O9HNt7JsWImxtqsD7vFb8TCyVUhe4pHDVxEMq
lzN3TJTgmxENAj4drvMHmgjAXcFjkBrfQucL91FuHrJN/rfy957zdop86y2h
M7cYjGFaFm7aS6I/2POUJrLbK8D30E/6D0DGmYbkl4ujQQqOJ9/cbSofJQ9W
Ha9UoWFX8ACvXnFYdvRTi83p44j9NNo69e7SkiPlxp4mObFSwSFiNZp4oSYU
yA55de8hzGFTgmnGCKiord5Me568mJ5vdIPezMnghOwmvr86D0mQI7N3b7An
70DZGXGYODwcI49usOquIkA7NY0LIr5JJSgTQoHY1UiBgJCHYZkRkHBkpqdc
18SJk8WLgxuoerEfpKqV1OPCKZ/6dnzZBpPICBQaQDbx7cxqDI+itZlNaNVx
5gEYLX4gz7CXBuJiby/oCbaJESsQI55RLdKrHX0B3UFChQ1mDqTqCeZzRhkV
UOMfIjtIkjunt5T0JDJ42lrFvEyTU5tYYKstKpNT3ZST5uF789G/zqzHFcYz
lmlDWUziTsXV1H9Ws1fQxyKrhXgqUIpQH6ZO9o9rzMWxXOpBKeGExq8fpLHm
vdP+6b27MlgY5UX9iO7HGzjFS+ng69GQYH9jr/pFzc9FAu67rXZox2zLzyp4
W/aR1chOEhQXt62tOxfL7jbGwhr1uOz6Gx5pU+y+ogFChz/IX8YIh1dIbcNq
cChjitu1W8JUOV27BPhUoxe+jdi1eSP3uPZesUEDqHSVnyD3oelCyWoet4sJ
8Qb8peBGpRkkPZlGOaUE2cgLwh9x2RGDCGRHrX5yvM3kDZIYRIPxtUo4YXCx
4Dpp2am6/Gc8BxpTI+2Kw+c4fhcICPxNHuODNTw38gx74jeLXGq7jSYPz1lK
4peSJgqUVMbnkNN1tYx9IQvA+EKo5OCxvkC1RsA5BttZuWFDxTKMAWhzv4Uv
ghPnP3fuQ7IERtZkNJYHpJV/GX91Kg0eD4NoROvm+Ug+ma9mX927lfU9lQLL
dzZgA/63dovHQymOzr+HodlGN+tMh5V+HqTkwKHU5oAb7/ObAOI7qSgjhME3
Sb8/ywZazuSq2tU/NN2eXPIWBKQQANWwa9DisrTQETRaqlA6tUyEAgLgRSWF
vF5Mz3XFMuFtHMqvoFd1n9ruklJ+gjfegTcmBzKEw5OazOSCYX9PhX6QtOvq
rNLPej0eWg7w85We/0GbxMKZUumw4VHDZfsA8Dft1dQNStGHE2HbSCFeyjtk
CMaLUnZs8AlEuL61imUKaVUiIrZtMO9AOeNdJlUHmwb4GwgICe8TRwTzFX+X
VJ1RWB+dRbRPhYgM8VHGRpva+kBV4MxR2mTJFUTPEDpJ/lD0It0dCOxkzYLH
e+9uM4en/RAWZCzHkRIVY4Zf384d3mpldTayGFMGqVVdwspss7FVVyNJ1tL0
s6epeNJl/LhQYZJ4kUTNa7qhDcrrssppecImTUc3985JWSXkUfdBDdhh+Mes
fpzvCJZ7wJn5Sp+9jwE9gpUY2nYoR6d98EL8xd5Ihf8gx40NPhK3bGnnzL4q
0yE5FzT31isnVZvif+F0mLawJFF3mQElG+aT/LOyUaQSrBhhSNek9sahsbkq
5mAUlbTg4ruIaVNp+yQbm96d0wGwooPKDLwmc1cvrRjoHcKBPxxiEFuSOJ9y
vpgfdPBS+0jfK0uqWzaa5lLcYAMwUZRqsqA8wSFdChSVoOCXOcIK6N9mnYGT
KEx/1hPN+ILIBQ9kN7DhEAeIlG7bS+sfAsibJCmJw3sTYSJX7ABR5ppgAWHk
zYoiyIt5ivjVwwNiKFm1RJg8NnYReHnkrMvDu6s3xd2Sg609yickfyHuz4za
RABfu3o3EgTlHvoN1Q2MtYyxRaBW4D5s24VqPBSHPsZHdyZ9fu4T6a6EFAGk
fJNEMwbHBReXFyQFIOIQrqKOo7xf/cJotDT6E2Ex1iNvpJfpdbti+xO/NJb5
qxatL6rfXiWuvIxWbbfyjl17CNXh9KdvMRqwd0s2sL/iM0I+rHMTzskes7jD
vIQtCPOCU6q7WizLmoRaIfNnZJnXVnmEJYXwv7B17BU/BjSWQfXYPdUzMwdo
zXpj2h6TxxABTrf2bY2xMLGqmXgQTV2+h0X2PyNN1MvtNNeqzap+leG1n+GG
Sqle+TVjZXPK2i/pBaGT4MAeXY8/TysKFVUlUv8Eou0AVUTiEfbbwtBK/DhL
lsIDF7IYxStrvZHUJQgbgzkKvgEB9TSsxw0p2TNq7uZxzC3Z9D+oZV9bUfQq
3FYVOrSSgKDIfuedEH9J2VYXVQplqmix3P30PTsFkjYxb7Wte6BN+yHFlMGr
M8YXgfqiCwwGl0jGl/JjFAjyjlcPKfAOjXns+wM/eyPMcPepKp6DMI6pJs+z
mFXntZ+a/kLfEfbih0OcIE7v8pEFzD/bXvB+hUVfflwnf8OZFcA+OP3dNL/w
OdtMoYQBOZWeZayHVkuzqobqL1v4ZZ7YCCvaA4esq8+FQVoescAYuR21B8I6
Gu9XD/FYVgMmz+ckpA83hb8wbS+sntWp2zMhA2CaZJ9w2YiNbiNxe8RD7+y4
uB5869NqotanHj8QaAL2rRAvS5Z+tYkOMM4gakoYxLl/NMd8t7T3zAhSRHsM
LKWM3yREQzSh1/Ldbek66ZwFmBtfC8WeivdVDnQ37lb8wMfccYlwy+YPMnUd
HkBAETGzseNT7NwvKfnOoYyYfMal0WWbz069hWPp2jMSq+JyJyHieAO8t2h0
d8ICM45DINv1kp+BfxPFkArXPH8/W2iRcl3fk4a5brq846CVrg0LCv/JpiC/
Vs1J2/E78xjSmlPBnUN45mSufsNI/NNCqVo80MwXkKLSe5+1Ic34O6vgOCr2
OXbiOt9Vem9yiBuqXjJDBKk04akj355crcFpb58UYvSenZueGuYOTjtiq4qH
C0jdsEor4VFOaEmsasumjkla7xEedGmsUFGNXianxibfCAOhh9n51KKbaWh4
pE13rotI5opJAjgt+85yA7dO4CUY7DQMfWHq/QapyRJHYpHrS5yBwXqm6mGV
qvIVf711DD+BHyJMUV/gYWLqA2omH1OSMhm9mnANB+WF2oYG0uuZ3Y2+gS97
QO0motQFaAm+xnwC9mp3yOjBwNikv7D7wW7Cw0XHDAcWjso0u9lyPRZFbswR
LzZ3O7jmfJVvUu0V/gqhM8niTtEGs5ULLNFyhAXMTx6VgL3kcqrxxLAXFzwh
aMh3aP4Q/eRFlb0AuqFEIVio2lvmzQijiupevxaZMZkrO8ZhnRgxSxQ+5nzR
Spi4Ffxp9ysWykRBuuLaDkRVtD9P++f9lJ7gS6Avh/O1FB+wyzIAfVf8e1Pr
y6O6EBNItn0+zPr4ojUVYMSI9y0kpPf8aV6BBY2xJZ25x21Fo5WuWoqIrN44
lEvojw/mDznvfGc9YhKE4yy4Q7VjK9oYebggkUDPTxo50uecrjqJ8EYM9yC0
uaBq1F4B8aFDmuXrbLZLu2cU0pEssbA0tMjEbzTe+bPruIxDTqXvDqcOguIi
hwaBIqrNpQ/RcX/tmgDGtm7lXL1mM4DPYYWn1fJl+gat44y3CMxlgeQmpZtm
5q5521ctKoapexul1uUDszHE8eK7HHgvS74INYe4/1x5VMb/WEcKQ/H7+Ojh
SN15myBnjfEPP/29Hh/cpeksRFhIKG0Z15qVw6hC/SAfzFIg1fGpJIpXo4Wm
+l36BJaP2MvYjWoRy/BF1VLwg7fJzaFcAfFKSkW9Q+4Hpjt5c857OgxGBWDc
c2RrOi76ZrxGVQJ1AZ4odkMTDSz1Jheo3bAYEz1Fis2LXMIvQCNIahUTXPNw
Y/D6neeyD9BLPv9oUbxD2Ib+FtUbH4I9fLHc9H/R/hpXoGbFwxO483TiOu7F
9lr9Lbey+zJArzgDCObpYoB7KV7KzlQ0zULWG3UP1RTpkyAJrN9il7UmTBWE
El3/8x2arilYttWWGA9UeVMfW+ceYKmmj3PJRR3gG7XqYJ+V/FKlb1AOYEH+
m+5qIeecMpag3BaipdtuCrx20T8A4xVxyFoW42ZGmMXnRNiyFLX6Pv34Vgp4
gwPVpdf491itQBK5cd+rNO1kGY0MgRg6JrVAvpsa1vZb4JMAGdJUrMZyuQW3
5hD228eRvk2pD8aVBoA+w4sLZu+EHQ+Z8w/qM/5quWkW75ATEaxASd5ECn/j
lm8063DrqrOyKQTeAQdeu40As8jNkWlp0dHCy/Kk1R1cC6Yj2sHLJSFBENVi
kqNewR1TGxdySvAj3ova5EqMRl8bD/6InXFUh0Ea16qLhb2WLqYK98brfIin
IE4PSfi/b++7jR6zlVnlmR+/J2mjE5p47xuu9EvwaflDcxgbp/WLNcXs7J/l
QB5vAvjn8ogpGao+528qlCBBEAYQDWVDuNjEAkGjtX/fO5JZX/T3tP26sI9F
vghO7E73/5fd0/kYJzAFSEMbmef7pQEWS42DJPFGIrlgLAcCg/e5nd5t6lI1
J3I25g/aTF4ScCrkFHDTXPHVyiZDXH1dTnFZ0ZQVkpZa8GceSltj5IoXfl0D
SFZQMVFxQoyqyCLNbDQoW6TArzMrsOXzu/mUm/sSKHTntVyHHsZ2mqKdC87s
MiH1ZypJH2HU8ZEX0GxdEu46T9xx4wyiJ5o1OyxDa1Bm5uxQrDn5y6PpDYnr
L5g2wYkCtANvNymbLIvzgHI9SEuT/pqkFbJz0MyTfK+xdgI+YnrfyPRlKNgw
Hxj5LfyRH1JHmhiCrRTd5xYAOU/7D3aoRiahlgbnanVvoMYrMVdU6hsCW6DN
4NlSpZ9uiniPFGlQBq7vMf2bS81xcZL8S6i15fiY81TvVF9org0xttqcc7Gz
UgXw48CtDM9koPsQay1NmBi2GsTQDo7XwR0XOsfctr8cQxAnYOv2Fy8Ntcs8
M9dtfykTBnNu60aE/7iM/x4Z9QgO5B8/I9h6tUqusi7qs0FoRuEnK4ZmWrHu
earKsmgdVJHUADjFtcf25YOOR9oIKhG+DZi5cx9KpAC3kwH4wGXLv1PUcC4o
lMJrzQO83++WScE8zeJ+LCazPGudGA8WlXB7WX9iR5hEhc8XlfLwee998t3I
gijzNG2ADpIDrcz7zaZxz6QY4EKGrGIRPnrhyP4oqiiJ2Ge9Ossa/Vo+upho
XZ8s+HcaTLXWB+Xhw/XGtFA5bsDOPkA5JNKNOYlDAqo6SxsfXAmKco7x56Pw
TX3aQx1oj5yzgFhq7Sg1PZkVG6wDHRldMWz8X6P+Dr75X5GvWM5bNGYaxXHl
KN3p3Yi3/JMoboQr0Xtx7MHBYLz3MH3ZNIgk82GXB3tOsvOit0aun9pnWpDP
oYVTWodqLYOHR3/Z9TTvtT+qnf1C6RMhBx1gfsViTyzz5nrJqkStOTWWC1Gr
3hGl/mJ6gYbz1hwnOFO8K1MO3MuONb8OHh1xTVWUwYN2uAXjyvSt8MBzAZkw
IZZC1O+Ne0Y2LeWx3YfUqYRto/p0GfuJV400JDOpuHth+My30ldYbLjJaSuv
J8ryJlIrwMiklfDVIywqmmgLQJ6pJ4zp4YChfZpxboeZHaXqcntFTaKEvmcJ
DXpz9vIoYBusqQ2nt820x6CR78zcrlWxYXgDmoDqbA4tbijE8c/kaVoiuu8A
dz3uHBlcUD32I6BIUzADXs+/wvleGym9U64WGwf7qlFOQQcgqC+6Z65skWKc
kgg0BXDU6fX9Tm/0XjplYAiRm8GvSYe0FGpIV2Rc+FioB/osu4TWwDk9AnpN
04o+RaWltWJl1Rgjvl1qK8fJGhkfL+ZiagHglpoF5Yev97KJJjFPi8DJKHW7
wCAj8MpZNRUXVavPVdn4+BowiIDlko0pxtRk2pEzGHm1QJ6Py9NTaAfIP3O6
qqKEAaQ+wATiPV8uW2a3D5e66ASa2cWpNAOUn/w0+9rLuBxqUasP1GOWCmvU
FawkLg1FozC1d12Q3uoUPrhUYGFEeVVGk9yMUlPCajK+ujC8u/OmUtXQ+T66
gvWliXK2sjnpr/vbZ8FgMdXhYD+h5AY2RqIwOoPKiXhzj7K+9mFT7WPmzSDm
1Ad669hOP8ciwgy9ka6yRzu+2BHyFrk4qDo0kDmZEyY51SdRfLViTliNaV1v
JlqYf86xIBBj7xlYCBPk5hbx6wsRtrMmjE940XQ+kBXreC20wMLdhiQHoG28
B0LHDhKYxSmjI3RDXp2eQEZI4yCJntrq/tJWaJg9AAXoaXXAo23P+rbjWfmZ
kcLH3F+piRCPoglk7sNDxUr2ZPaQu9tYJIcoakbUHjGb2tOk7OmMMfF7jek8
KtYsjYVOT5vRrMiIZVw7NW5OFZL+1ZyZAVfety8LBBC3czkg7SEP1YlAvvfT
VF09qoASuLBXXBl1UGcISwk2Fn9ERZKyQe/OuUsGnfE6UX8NDdtu3PlsamqX
QXAN7JFbUJfIaAurDcyYq+nh52YQe6Iy9GzPoccjXCCZoqlK1e5EsX9n/aOY
TbLLwoWWQajRitfdke8NjLcqInItw6WYJHaPzqHLqVXCSRqGFlDltZe7Th/m
/bUyKDTMxtO2h51sNFIepzeOOXEef/LFc0CMU5LvLLz/bjU1qf3B4365vQ5i
lZZCIQACZIBJrzgNZslzmg5Koon2ALzcmdjv2vdMuSpqQ8J8SbDSwSbmtPii
MCUEXR8tDY9H0da6jj2QGRxP2l8ZHybe0a1d9VgcFSGh9D2UDE9PP3KzhlrB
BCrlbD2WH8yvkW9yM/eZ8/fwt7AniAwPFK6gNlsFSvykGC6dPVsEMxRb05WR
zr83A7fhhJYYGw731gXEJDzVXbCrBtr74m43rBfJnAYhATffwhw2PxmSzpwj
ucEhBXBRVZc/kmoNlwoSdUeYj/7G2DxOToSfngGZTpLw4LWRxiK1glHPN26u
0B3N+GscqFwBOsXplfbojYXRIpMQ3TU0GwxFUQZzdtuAcbT7ZjEZBkAsy+MN
pWRlVPQ7DcVstkJWWBMIpYmkg6TDWTV1seiuvOaMVmjqpRZM+umcEOKGzfOE
4RHTxtL422bNGCx7eG9aAIuMNRXByjCpUM1JqumbzyAAR1uRdZddx5o0tfXL
w9mkCDj0pggvL3BFTDaTiljyr2Gr4AKvyTms2BcRbBgxQxbggcm212QctTTp
iyrrXJ/PQXo2cECAOi/mqSqgoV+I/I81Xhgq3XUR21iVIrCdaNG0Lfe2AgV+
abg2WO2OwXeD136K+2Pqt7wGLOEzzX9drPb9D3JzSBkrR6w0hcIN50Gn9iJp
uzR1F77jrSocjMY8t8H3zvXBBygnqvBuNj9n+ABCA5hb18xlJDjWQulwqvDI
epQU5iTKuyjspbc9HW2An1OwnnYhPxKIf/dmjpVGUjZpZv/ZS+CpAP91oDKy
IAmVEs3EQL4pN6ryzjRnj9GPHRAq6lKKJS+7fpUZoeT0pFK4cdoDkb4ITDrx
yOnrxv0MCA+IEnkja6BDDcmjwra6h8Tmp6viHsmGU56M8KUzqm1Vn2ISTLtZ
k5qSDewDOMwkqfvvRONUE1e1A0UN8bPHluvRwghv05zyTFqfmZ6e4ek11ETI
pE8OBz10gxPGlLr01ulBNUwTI3erFDflLLTAAWh1i/sfLDZJTsO9sNFKcQEK
28b9/RcWWKAEenvtK9hJVsjzPzU2YIDvY978lpPoHKusCyOfcnmAmf0//S5K
l9MBLe8sntiMGObEYfw90g2GDPMoL3Te4g3P46B+5diEgBjFDRn2JeFdeKS4
eKCR0MfwgIbj1hi2jqnLA8G/C95dUwi0q+lWpWNtcTe9qtPJniL84cqe4be+
b4tHtjf35PoQwoWVnbCxBsJCGxMNBGzp6902oLgen2uh8QlVer1ird7Az/1V
g5Omf0ibq3OQEt6A57Xf+EzbYL/PiynWt7uRNr5P8ahkVmdqq+KK+uyutvx9
q7SLEMQS81WI9b26c0TFBxH1nWXTmySS9vc11V6H7vscruNk5hOLb1a8Ptft
dIqQllJ2xC+Rax9H9z7A3NZkaKqIX/s1qzrKaWQHNEfsohGMcqtugJYKDq+1
0h7/JABfgYgSkzornnS/Qm2v0NzfqUqkpKT5Oue+NrORHX74g7fNcPsbSsIv
0pY9ALekjkhlXMSXrCZzxCZil1h8fUE6m21KRIcv0uQG0mYA7A+SvxO2w+55
GD7onQRIJKbe9iDWHrKWsp0OTzYOuidld0Pdw4nL2rIabc4MAgrHRX0nmndE
KzWoLHFU8DTF/pDoW9RTsQ+CI/Z0kxAvNNm7iMR7uFQ24bqcknMWpOEgwLf2
lKk+m3NMhG3zzqtj1MzO5AZUUiSWZ/R0mBMuoUqOwMFMVMIypnymN0tnVdlg
purVJxiTDslASpMyf00OrkhGkaBuqghpju9Cqzh0Q9n/Hky7jzR06iHKkdkg
lI+2PSpRdQQC6v6r6Urf/t73nVbwnchchJLyakwpErqNfCu2Tn472JC5+Qoj
rI0Jh3fYKtS6c5iMb1YNMymV7z1b1jBex46lEmadR4uGvXytnszL+tQSW8HN
sJdAykjgxFhgwcVF5+2HWsBnTyzbA72L8kQ0lGXHbLghM/MAWzVy1Tk4qfON
wcDlvl18npe8dTYv9UszQDw1YQ6fT9Oab4+HVL3PeCnSXWwKDjmoR+F8UPNg
6IAvcE4wfFDQzejozA2zv12Id8DyGxY0RDcTO5JPT0FlV2Y6HKD8x6dFxd5x
+G2alWKlIXe+Dg6oj5R+JSD8/7JaD1SVtE33uYhNU8UFl4Ahg5IVRTxY7CZT
A4V8NbxAVr3i25d3gcQ2YcQrzng2PwinEy3sEdSeTZOaQlP5YI/4jgkgy7Qi
0C0B/nptsY8wBS96KMhB3VHwgdQseF3BX/xeo1IbWTewlqa2Gr9r1Kdu+rw3
5U79vxPMVig9/RvYnsu9U8CjbEnrDZVCRMwfi5v26Qu3hy2cv5vtYGTgkm2z
JOMulRaSg6celiHuxD7pUfyIjhP4nMWk4c51ucTu7WnLwgKeMuoWSl+jQiz6
L3KzRtfqeH5m/08jbU8yvmAhxnAC9c/eETT69YQvx96A2UtyC2jjBf17zGOR
muwhsEFQPhAoXV2rlIFp9KC9PRLbRfp0dHYZK0U+0xc/G4mZSK6WP4giTFqA
Sv8qFszuAfj05iuuHUgoQyxMU1baLcmAZ46NoRtAXUHFh5GWhJgIgwY7445N
nQUjh+gNbHm4SjAYfjKZK6732SvCkteIj1X05fZou/AiuZxQr7r3QsvzMIaX
u612mCInuep7aJIZX3Kf4PG878aNp4vqbtXfW2ghknhekHULftVxAU0a3npo
AlgFjxGDJRdyFGDMWhJ70+lsTUY+okOy8aN54DR+o1Egp5m4JXzKIOrMFpm5
EiZo3n33A1WlsAc6BNe1fhhtlzKJW89zOT/cGJkqM8DM3ecROCd3TyztOJLy
zAk5lSIf6VV+j7lk34/QuHDLI2GwTR73RuVamJ0mB7f8f0pluE3Xa67yc8rF
dQdMGQd6TTj6NpFrby71njbZol6kv5SoePXqBeerjSyOQrl83bYuAUAx5GAA
/I3Yn1vneHmaPRfs2mICrnBZNti/+KrhfOy+Dd99a1F8RMAtPRepUbPa44ot
w+R+48naCqHr8VcGsZdWy7ipdxYaLQ3wl5kaXcPch+p4XcIJVBq0MViwH4Rf
tWKnBnCWoT7qoRLeRZqpmehHL/4ZSIj54CCooZDCajVIGUP11EZLBVSG6DWn
YrRM3x46ZXsgM03M5uA2cRRgiEZDLVpb3mv/lOBvCgkEexQPeYNYOILtJJUv
Gqw6nbL8YQVtCC6oGE+FBiEGE82PkPoV5w03EF4F4UtTII7fTm8oLZNs6hNH
sthBhOAkZxdoJyN1JyoAxfz9bgj9BH/c/VMxCUWkn9R1GqmP3q9D1ZL6pX1k
RoeU68BsAEQVV4Yun9U2HJMwjNRTbPrzAVYDHVQ0tAKA10XEo2QuckZ2LGfn
6GwfWxd0JOLTFC99tAdI6rGbiPnyYsmZtbQt4xDiMDFD0D0pxnTUNZp1NioR
i76bxIDaFAly3lpElIt2QUkJIMmkWWpvJGicB1UAzi3yNnGCNRfbDRgkTxyZ
OTm39FWe/EvryrxZDwa0qqULy15x/ZUbhz4Pt7eEmH16e62bSXmGtpkhQqtz
WKzzmCdXBp3ecNX97ggVddUQ3BQv5n7hm2CrqA7+fy7A3v8AHg2mN9AnxL8I
tQPkl6H5ywuBuiJAAX+eFArVhIkrhlXu2ujvHb93hfwehi0alBnRrHDvzzmR
DqR5efU2pLk7kCErMSchiNt2JMcWurH73FDX9FxveMdXJE1by9RQLCLethgt
tV81Jv+h9OKf1w8+S8rTP9F3dVi6OP9PCvqU1mkPp8mSd8oFHi2OiOyrJ4CO
d2rmh4GC6X3rDd03oboqfemowEO9rw61YoC3gaCJ/aF0/aInIo5nmIKbJpe9
lqdZ82dP2nyHV2rHVDgzzPWHurCs2sczwBUc4FTvlCiPBlwLJnFOhryLyqT8
Ac4FsmvBzmBsrcCIDbsjjlJpFhXIm/vzG2nrSSupENH5G3GniEbjuJJjjxxf
Xd9D85IXQGJWBDtYIEi3I7ZbJtb8ylrAa+BdVeAVbetQoATkc4+mC/Xkmx0y
KGAvMlLP8ZbnTeRTXvl3S9bGjgABKykH4O9CjRmsilsQuQ3qLd+1drUvhBuN
JYckq/XWTLv0YLI9939ZvvcbWnAPJcqlUbs66vFWpPcvSBu7rEQ0eDQUOm4a
1WZohO2NlF4VZqjYexM/FI5GEKGVRNGaDB6wi2dBA70sKgzEGyocS1xq1aPw
KV+lg8YiEDB0AdXxy8+I6fbdbJ17s5wdtGkG1k72lfaRhmteT0D8IkMnlHmd
vtDvcz99lS1bvNVcNtiYrE9PSXImmYrqTRueuoRu433eiCsAsbAlF/U5s2nS
o6gjtiTi67pGhxLX5ekxXrm3ptFfW9FjqCBtMxQTY2VSrbJDpEpz6d5D5xIS
GZ7yu5URg+80cGsnJDeqHfPEy31VA0ld9sD+imZ3tryxOa4uEspq421luNyj
27ttDk8jAw5loDB23WVrkuZluOzLG4QOur3eyFOb0JIpmfyeG7XV0pgO4STk
EfXmAPnUazKHYJONOFaXPPyseYQqr65/8o6oN4YRXIqg/Crnc0ddXS9GL3B5
Mwlml6/+Vhoo7oz86BUMzK2mBi5ygo9SBqE3FcRGS+ltxK6Up+oM2EeyPq+i
vysBP6pGqYErLFyHWYN4dUCcFQU+wl4x2azhD+C/WTnEMTGXM8b++82uTDmy
VL8PTvERdQJ3dHTDtEW4sae4gq7vR+BA4qFK476sOz4Jmd5IAzMGnJ/BxTzi
cmyRDodPW3vUn3Md6no6stL13rLYXwyT7EYR6Y+hiPaI6DctrTEBmnuq+ydB
b5s0ocKElr250lBRWHLisqHfDQSamtBq1MEFSe65UZSfaOaS/Mppb/tA6+9F
fcrV5bWrT9VJrGBybqNAEcDccJdfvzSHDg1C6mZ+lWIW+c17mnvh4+go3xoG
hK/M0bKJlxurkAm9I7dHWJuAzIQI+ORb/bSNmXrd3DA9gXrmz3BUILm3hYLy
DgbAFvR1t6wZiBOvfZ8525GSl3dwTPVsT3UecDFuDI9LHX1pLpX64RmGlnCO
N1zWSFVfcSn2JVFDwQZNPGTY2v0o0/fCVcLZ6DWh4rAw/bM00ytdRGEcloYe
oh2MjpDmqNuJCzKi1wUV0Jk7NefOnSB6NjAT0pYzR59VDu37UG74FJ23uQ15
tlU82DFX+jtHwvS+aSAoMYi+nZ0IBWpaHrqAFvBBUUBgT/ZbAndMqH5wih5u
75Q/RFzUm4VZyL2++E1ngJFnkeuGW2aoxh0iqOjExcAwgwe24gEMCmQ3kd3X
Gt9J8cQ7duD9SHx0P+Agd+WsSx5u8TO77Foz6cxjSrbYXFyOdQrVI7KnKn2c
hA/Bx7tcUmF7OiklnyNBplKqXjvP+sSS5emdHCL6cSNLIcQtSPo08zUJmIWj
4X+WBpaN1xp3lbgxal1J/RQt6G67piYVNlwIcYVsPzFOPiUF5VYi/B8fCTvV
f7sxEPrQOwVbdGPm8syoS8l9humigzg7eKmSsLscW0HJ/0ezE+co1LGVR2wq
4Ujy298axCOkPoNP0eiKWTniXnXcSQA1mdDYqvn2ZdR/eVsGUoELaO/w2Qsv
WIfMv2nZTeXfZXAkDfHvTKXiAbdL9N7g2d3oFiQc3CpvtYvkRloAiqEPuWx5
EVRv6eeW6aQJAJ4ikp7P5ykgq/wYyHwNbjceBchCEnRPbDEV+5Wo3DqOI79F
OXQB501RNkhGaiAYOTDBysbG9lGa5jacikHB+btMGDRYcd9OnjMTbxW0AxZB
DpZ14ZdlOKLay8UiM99MmgmhjElF6B7ynF0H7S7Zp9VOeL/HOINzRZcHYxQ/
fI5YFw52KqukOluojb78TNKIMg81RSnTO9h0HAOhVqKRDk3haA9OGuiR02cp
n6Sj1VnQkrV14+4TjZvX1EbtMlK/Gg5z/iB9gqaeNvuScuXJ8v5eK2XObjKc
Fg0LBH6DrxbEuHysAEhZxhmy0KirPvpkIS1Obe/H4hbP7oo6HaheeruHiqet
kXbG7IwZ0LwRSz8YBRRMA/Wz0MRGR4TXT5EBol0TvOd9fMeQaWEfeY2Ka5Ug
C2V2Vcy4Kya+fWiM3yxQJ6e01vYwlh2ao+bCI1QTiZt0s/Qr0x8zglfjPBc4
MKuRw7FpfHMYh7ryPGP2EoSX8tCe1pYqFXTUAVEHNTZDYyh2g34P6nUn9mTO
mow9KIVg+qsKi0PJKV928MO/HAqchiTiiGrDSmWhfznJ42+PbE0uElbPFOO/
M3GuDOyo2LK+wnfzfiObN9ASztIcsbKm2Utq3tn2Y1yU6k3URVVJn0iZNvo9
tP/em01Oo6b8U+iZAPQ7z6jA3mLa15evD9D+eabLEkgapUy6+ZYueRFiZ0nc
rhWCkUecbODlyvBm5aLZSvpLSLHgujYmwXfCrX+fXxos90GmOvJ8WPGf5MhL
zQVPBc6zFVCqvivEB1u+XvY2QN+2CvNP4W0XR+HtLgj0YgigjHJiUBzlDG//
+2nHbm9ySnrk0NUIKZjtGI1wHr+TO6oVytimeQU7RQkXMMTOsmaket8zOwA4
wd/O5UeCFdufejVUipnZTx7flr6QC42v1TgzM2+WqaAhG8bMjUsUvahzUDD+
zq0d8ZFShtOzIHYRziv1Ds93QOpc8BjXHgWnSEV2w+Nx+oCIVtFXK1/N12Xi
zTM4nF9+0HRpCSupbF/1JdSYbgz0jum+pk/zvgiwnFKSLJNvnYiEutKvlBHq
puO1ecDyDjLlZgzv0DweAC1dqPYToUM1DoXiV65wtgRhxc9aAIgCLbFItG3t
yY3VRmOpNilhnkw5iMxbijYQTodNBXO51keJnTiva1QwtRs/8Di74YSAIIv9
CJlKZysxLpkIClaiSx82npXhH5dHxCyBBM2Y8KFyojAiEcpknulQvZWmWLiY
4gs5arlm+9K3+1Kz8Kdwt9RZXFx/XdpVFUxFCnksCoc47Q0w38B+8zqJWpbV
VAkplqNTGibLTJAZHvkVb4QmJ5pH3hsp5yIjoff4e1wA5yf6nFf0+TvmcLtM
vUu0X7SdSwnuhEovb/QcGuxQ3sKp+4j9keOWd5bmoxrLDU5vaNKi7hiHAliG
pB4o7JG/H7H4LGhteHnSUuznCIdp85lGbre0wQOmhh0oGya2ANUm+EXAz1Z0
aSV710fKXLhfAxd7IvPE11ZJ24uQEoCcFvQMF64XYltr+N7V7Of7t/AJC/sb
07YsPzzVPK8GWNkUNCBNEsJS21GhWEX6bmhBgSahb8tSGvQ7FXeXpGPCgLt7
rPinf0+E++fWZtuw71agIm7LCEbd8rHIsHH5aIZoI3WzgEIyLZ51boUp7zsI
r9zXVrXFaBFL86ION5zLVNw/uKrdvCjFp/XPGCXIvqjys5e2ESjuu9AYk9i6
i6nWrFpB4a7TLLXLjaB7GycXa3MVcaunl+h8uLUrTYHlMjY2dUNgDk6UQLHz
uPL9uc05aqdAilyqH7a8zrqEh503Bfd+rT1WKxAvQPPd+OyPBb4m2YJyukaI
uSNnNFtCtgLC/iVVAChcRMekoxC0BCj3OOWGs2YJWIRZEgNfcdXRulfRAneU
gxVP5+beWGlNXXqf7KDiDRUX913DyAXFfwnX5Q3S8gI1Bdr3DPy4w5aJDVPE
9r1U8C/j6URruavEvxcTYMx+dOIoDsdbemKSPxMOtivy8rH0GcBOkBCyzMjU
A3BQ/IknaUWo/hf9ngC0VllOMqEq8/mNJRS7+I8dYalyzDImqhIxOxXza8Mt
M4qrKBbplxD765DCBRCwcfEptqsSYZyVq/CtjmrjCdaMo9Pd9xxuhV1pxBbw
Zi9bt+6vAnp7W5mL4TAfESYdnxoSfWXBDR66PPIS+Fs1EiHFFHsNDUNbAbRP
o3aWQqcZpM/l8mI4XSaOYD5CxVSHJrwF5ngDgBHXeXY4XFviEum3jkXSctqM
rYVRjBNAPTKKa9IFxjp6XRoGOKOPYEK9+ksDm876EogLaYUz8jtdVZWOdU5Z
dy8TQE10to0BmehyAPkUcpJXWpQnySlk38RvuNJ7qPJ9OAp6arsVUcU85VCk
ksCXLsAWDhKpqMnq7r1iEbtRq0BJSk/iMmRVyG2g7SiwQODvDTrjkThZ28s1
pjh+Hvhs2o6sU14r+pDqTlRxUWMB257gGuIZomoy4ucP1Zqht8RcLQw85qNK
LqvVCtcJrlYw8xWaa66qud2lRWsmEUzSvEEPIlW5WM5lAkwPQq8V9E5RuckE
YCfLziRS9X2Cs3pHQczqP8txQ9j4uoxFBntqaVhrXB2f66vwZj/AYAemZuXR
RVOwvvKEMsQq3rjow7kCe508xlpehLEOT8G2tl9o4EBTMxRSrdQsuFivT+rw
wA3u669kc3y9o18Mhl2NqbIg0lU+3PHrXYZAtjuIj6YQn+qby5C679zISCSB
iOo9hwHK+Me8pmvK4/06tu3XOxJQo54GV3fNTVadJINcB4B1ochhaBgpO/Wz
xj0fQnhbEzt9epKJPBtbKzCSTkZRWi2ZiZigJpRx8lpbSIP+qhyfRTzIGIBA
3R8EP78mxc9qQAFd+S862wavsqlwcUy7cSN9wYNolZE50ANSyEtm/Kl70pch
EM+I2E25R8SWbu1CeeGh+zdk+KXJT54bIAw9V+S06zwWaIUSYfjjidY1KkBp
Z3WVDqI8zYZbr5rFa7hyaKNnauyxa8vq8OVquExr+KcFW2aTGCMUzEus3IXY
M8cvkcNNMDAUcryUyjicI9HDWF7d6jHrqJs/7ioB3NHbX0epHg8K0YttAXuw
4a1VCkCRN2P3YnIY/Fb8an++fPngFpqUAYcbBoKKrEPvKncpMYvR/cpr7z6t
Eu1VKZFk5ad71fw5aMGnwU0O1KC0qg7SHUVLDiCZSy38n8ZUoXb5ShsiQPwG
8o6gW6yMhr7SDi8EMD+TA8cIr5j/9Bl3+oAqvRL1gUwjwAX/iK56S+XHbgmh
DOJl3MBZt4L62quASi8nKVqrJ9S/Ot6RbDuyxMgho2KmxiQBOygWkN2IMI/r
SdJuBqdl3K87kVpo+7wnpk0p/BasfPl47zFNmECf/kz9egM9hx/d7sqQrSVU
tr4NQPL4SJbGm673nntmT4SBL5AYX3I95zDPJx7Ck+v8miTepV1J1+c6dCZM
zFP7wUP+A1fzzsxAocYA8qE5MsW8CAuRwtkFxf5Ea6+wzt2qasLbmUIiUI8L
we0tWd4nmXxT9lxeN2PBnF5aDmESwI3Rc7tGSk1iOMbpALwYY6mgJxUfO8Pk
Zwf58P6maSig4os9Hl8p2Or4TTl7Hj/TtjYslwMeEfuBoB5D1l5dSShs+k0f
K1z7caLs3pvGBYr+xfMi9oS52jzAWTHSKWJ7qWUKB5flT6rDh4p5aXst5aff
IVZvxloh7cs5eZrWTBqOaj65+3I4DOrl1oTTkP6GSXvEKOgTjtUcNw1WUQ6c
+ovz5i9g3M6COhbxNAnQ2jp1CKMpd6shDUOI6lE+QhUkM3uOYF7vkzgcj2tR
j/NqRQYuAhnSzGMMO5rdkYBC2t2JxMifkpaQRTAyAGXx9rV6h1cUP8CFjAjo
pwZI4/e3rSfF7V9JVGNDP+wfYLLoEc0sg1FMHj4XSInASbrWrrC2mni7SQQz
7PRJxJaZ5jJFRKoNkwnCYRl95ExsgLd7rnZsCo4FhqHmG3KyLpTiPmR5itk4
aiMyXw8pRpDc622SEyzkmgiIqdwOwkFterTcVH8LB1PrWmRRopxMo+Rybs4h
ipz1DbC2eD3W0k0+pX5PhIvVRtaS8rLRHETBUleHon7N4Nh4VbQ+1lW4peXq
GUnY0PLKx3PzfLk6FTX/GGDjxvPAoW1x0+W83wiZTPXXwFL6lPxNQeWjjOwt
epZ9dtQfg2f57ek4T4bGzyS8JvBpTq/GAmP4gnY0AW7o7Wx0LdrtfkqhKLHc
Cs5TYAIp5ihOtfTnRCO3ugQ4XVJoVfTR19hgMqx88Pum6FlO2Y3nsCa7SdPb
7b2pPcJvK+4j/vkhHn5keF3aoGvmoIg8RMTKg5Bjvhxqy7WRPCxJga8FeDve
hoXCs+V2sbGnoRpEZg5/2UB3FXuja3xBiiujvV++4fgBhkTUdyS+GPq7GM+Z
1dInCHQL/Z+GMsBSAfoyZGkFETWvCsU6J87Qu7D3vdE7PEzA+iUM5kt0jKvB
Pz+iHFAgqIF1Nr5rvGHxlCXKWvb0Y2kXxe7tW+7ZStul2j0mNur74XZL2Baa
rAocisAE3hiWMnxvJRWNqLUkSfnj99r0BalUgKRuvkEywR6qbkZbLUcEHf9s
e04y7oSl07/vOt0JpLVi3GEqZMHBq/NBr3iPhWKdz7YE2R/43zvPzfHydG0V
MsUX4EbCSJztlR7tyuCeYJWuTWJNXtDF79nbx6W+nSQPfwWytgYDi8W42jza
fUMJdIe4J61DFIKA9nWek3m97IL9+V1ukkloSiGqrukX1Xr+lDVU2g+d2xwp
LUjYNWF9a5umOSN8/pQD1MyhzbLU89jLo+141NTpkNFly9I+D6ggpZx0W+eL
II/TibE6MQrzAsZLBho130Ru+JhZeO380BByrQT7BBD7/zjKWt0zkCzGm53Y
KLiIku9lRvDMIuFXiJg5VVydejyO3pV+bJZ1THYv/hEW4h0oepLBUckcXfc4
pCFfJ6QmCnfOVblpUsaYITvS35eMURACvst6MhLIXvkf1L7MPGqi/2mOMug1
DUBm9fkvwv/egKKipmj5of45WnjFOVVoR1zRbvdRThIIkia6j2QfdENmvqfd
6IuN7eRycsjp96O7maRKOzgTsP32+aiOAuUsZM/9ehbf5wIEPRu7CC0n/RL4
xMoaIt+mE2GaUNT96RCoz/cUTFSRvusdlgluYs2Aa9mUbSdYKOX1BmleW2lz
8lUDrOXrqFazjQzSoNFzSjWHZRya1GV2MNJA4nawUf2kOgYqJ24YuK/cZe7c
R5QWWfIKOdgWUsy/Z+/aNMkNLITy5F4x3dSxezz5OJuQkhuHeF375TkRmko3
SkT/J+PwvKmBzRP0ID9Uvi+VlU1YJPv/DfakZKWHtaa1w5QWDKkn/mLRTwXn
B4ZnsFQuz2g1saWHw1sktK59n62hAWcFoq6x8ZIoah0xS5ovibPuYzmjh8bB
JRv8vrHdRVCvxw582u1pDcKVJ0fdoRyyKiEwjOVc5SYqIjAV/Kk7aW614cE/
EISm4jGa0hMdVG6Jgx5e3ZAuI98wNu/8zzE0WanCdGRneiR5DzEfYwHx4Lhb
ybXwEyI9K8QDUbn20iCM/VQHo9WBf2UBH/qYy9HkPqci0CtYekAaGqD+PAYK
NIP3xYX+fwIaOBqWai6o29R5/1Xq3ZD0oGNoblcbRFHJBvZaaEo4vOm9S1I3
CMtWNpT+LZ6i6x81MXm+MA4LccVXEYytNMeUjCL7tNOpmgPP8bQ7xejVkZDT
a1OGDS+vsgf505MHvSMT9XMs0rea9niwV0he2SoDwYsLLveT3GvelHqX0p2u
9MTiUY8ZjTYYssKQc8gxTwtLLhAnGHZ3yFHvx51Tt8hOYFWKfI1P8MRPd/4O
sDrSjR4ywg6GlaPr3zJ+Ha0l8nJ4166rWizebYOojUsGgLAMNixiHq2HuJnS
FIbt0kLcfn67OWwexG7sbyFmecjqFbdAsaBmusT2Xl2XFgoVCzuZG+B8ekl5
MvEjE3NjYJmbzuACtte0m0N9Qok6QRbo1kVYHwbvTleraMORjCvb+G8yDHAv
yRQJyBshcrkwkiyNFnhpRZVB78+fJhmh+EFYLR4QZIW6mRmhHBEqZhJ0HZJH
T4IG2qLhNtj3S5uvpBX+F+hPunRorPjs4LTwAHz9qUiPsRPvehVpgKbwIwBL
LvCNfXtOwdezsqA+NNWhpOhEVnmUZbj975906XzgFJIN18ESfttvNiqXuPos
syvKkhgd+8rJ3dOfEM2mpRJiwVC8F963uKEfRnWtKSqICUdGVsqsoRrgJD9O
1fV3UGPkmAY/DgrafvzO3VpgSi15/ecadzvGSrywyfK+No95nRsyMZjWJXkR
OMUtFer2MvqtaLeTzkrlBU29l5GWt2pcCchMgwwJBGxBW5iw6pQ9H7dkmqWp
HNPV1k7uw7EdAPSE5glORDMjWOHnY4fi5CzPF6+xw2DuiBBon0ImJg2lqcZr
azKYtF4kyo05Mywh5tO6QIo3VfTu30/Z/4alAaK3MOtrRXJZ1vahELd15zOg
UI5x/sAhQ2VtEtNzM4J14zYCZiytZ6rEgZoh8xZLbMGcYTYXBmcQbaaxQnUS
4Dysos9js7V1wGMi57gOf6gqbAgKSqQHwofrA4rwfGGcqC5PXkOhZbK16yNu
OTKNXXaCf/D1uyu9auV1282sht3qZIqKRdWDpRsko5czex0G1++pd9Br5DtO
GbUhULx0ZyrFfZdBNXpNGiyu1+Rkr62Lxg1Ki6lBya8MzhwLkwRTvokCk+Ng
WU0IGb2eOdWFLVpA0lRGBEj15doWCJUxXfQN0IQGbXNnz8YbuzSsWuYl4keN
Xbsvfpgqlem+ctvxZRhoR2fPzup5HU08g7+C5xCQ2osty+MXC4zmo2rejQ6M
MjCuOvZ8FaQKuKeGHmXo4npoCfqG7WkuwLyffVmNjCqNA9xNjs9BTBjBVXc7
9XK1YkDZnlWGu/CWifxSH/DY3644o7qk/drzH2YcmPpyYOm+PfDxLrQV7nez
MkCCnhAFkW81ohpgM9FIwWbEgdca2cas2iQnBkcue0SFaPiMVeBau9V9YkFv
zjHZRJL4jonS82j//zIFaNWs2GyEmEizWx5AxJMzdMw9ifTJ2K6acJSOS3/j
iv62fUTFnvLTO4GCUcxq7gNZQh36imoesO39P95kQ3muNuOH1Fder7yaK8Jm
R6vQB2nYrgQwTgO9LvGVXHRuu0Ab5+NJTciFb/qRGWrzoq5vvRKFic5b494/
imaco41+4SJOVsyi0ue54+E+1Wyup8CiuQAoW/CPiFTRaj0+05e/cFIaA/s7
d/IyEu5zx93VNun7ZrguFGKYoSEXwWDqAj/U5tBv70gUwfLcD2BcBeqYimP4
0g5rc8eB3Mw9lZIbQ0BSAm+DsKj2L2abW6sNOKFBP+bgBuBEghgapnf0CD1+
DKFeZ50TslcNZ59QzD1Pb8t3WFoKuc+eKxSWChIh88t6jWkFT+kugM2lF/Hr
jlkflfgKmcmQRCpLt0+CkgEXYkLxERDSZg//B3liZxnd6WZ/tu9yFvg2jSLN
r1S4pln4kFai40pNECV56ugvwz9Cf7QuGsZZ/fNKJtjM4TIbhIIo31T9XE1Q
fv3ez2qfElWStyQb9K9ibjSp6lfy7f1uI2VMjamXoSqBsZ6CrgGaSfjC2EFr
+nzghLYrvhODhOA76P5H5GBqDCKcdiWDITu/JRWltAq360QS2MvQettwLe2a
uJjkKmtR/4T9Qf2LVxsIjy4EKl3df3Sal1JW6WXHKgG6cPNEiiNVNklVErwK
O3opr0O4bTeUOW1dcjjPk1A/Jo8CJl9syvgeddNvgPQ7OqRfkKE77/lpceMS
BMR6rNt6Jb5pBrY18HkzqfMl+wTpnvqcTiYfUpMgGHLK+6fMTfJLCoknHLxM
vI7E/gi7Llzsqm6OKRtF5Jkfd0dgD8V8N3aAAS4BwG+lG9zoj/1pJswqY+x2
5DySbTobDUB84MZZqfZiwNMycfI=

`pragma protect end_protected
