// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
sspW59tcYe5aPN1Hn2HHSUrh3vWfvk6YnK2JmV3o2azG1le4s2NZIxOXqL9SQMtV
ndFFbNEHKuMPc3UwiIQOI+Epiq1JlxMb3ETEGxyXWE8n4XmIPd7ME29GnfKy1peg
PuXMHnpcXNswcxy8tPGmyoCGT12NLh77JPQImZOUkLM=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 10272 )
`pragma protect data_block
gy17Gg0WqY2jDgdknn9bqV0rKZhS1PMXHE5EEPXDonx36niCpyrUeyUKANdz2Hj8
pfijRhBsrDrFEvpIAAk5Ih4yzifsslKBp59MvFjleO8ilP9g1ptU03VX4EtT1pi+
0GMl3tIylaSLn2uhY17fDirsmjGg6vwiE2XlKwmRV8dfXDi38+REOS5ZMjmf4qht
m2wYo/0Y4NlPMGflfKtQj4SlWpPCC0EJdeXDG08U3IkNo5pWhc0hqxGk/jyAZ46G
DlWWboasbWEesUa7eU0QnOGuvpMLTG0EJa83TZpjKCnFYsxJaif0cKBkAi6WthOC
rlzGIXP+krC9Ie+NP4rD3bO5FwmZPSVCjOBsW+psBicZyG4G5onGN6SFXSZYlqHx
qyVDegwcQatO7Qqz1Ytezrj00HkiKYV2trBKSbciPBeUKeOyieVRAaODR/1YdDGd
ANcvWwNIhdQOk0FzWP6QMKfYgxXuruWhV8PQV5S6jBMzMvgtNj0XVJp1ZoBT/pGM
2FlAC+bOkCc2VQRNAJSIDQ8qxKeSmX3k2HOJ2RaPj1n+z1QqBXAQHRShmeB03vs9
o+ZIKb5rdIVbJkwXUmPZHXCapL/bYp8PgOhnPkZF821Qb0jSeK4JfGQGbTQiKkT+
cmznmg9ahjW8Q9d1nmNkQHCIWIabKpMIjrIFFJZ7xV7+vchoUwh72CHKwluGnMxM
T7mTqXjtMj4VkjLhiv3yKG5RJtVj7pYpWzX7dGPHYcmBGV+WxB4x7XceXmmwBh6x
ljtaTr/mIbRwiUyL/L7BIzGg38YL8P/s3LEQU3pcKWm316wF82WQAvVpbk++mT1F
HaD+z6xYYLcHnYbdIgnnNT/ADy7aKlVeJZCo+E90sjUs3DngY/weN3OxIj1i59eu
L/Cb1UIhmG1pV2KAeDWQfynFXkYa0tEwX2vZk0C00jbVNUlCBu43ixAZA9p7ZAky
+mF/2icjl96LP4NBUXZq03fMU4dCKNSo5LD2DzJPdjUsHOols907K3m7ulyPCT9r
3V3XSKcmUPY/XZQy+7Wc2m/sQb5/JNqxIlhZAgnLyw6mI6Rb8apRMxFctra+aNoY
Tfd3fUMLQN7tFZejxgDwzp5SPHcgQbVT36Opxad326r61IpaOl2q0lkU9Kgp46IR
Fx71qTXcQvzLPCQOKSsVVaS5SaGRFapceo7E8S4afDVNnmL+DMddzrN/YlNiMCua
FK4NcOQP7JsYMj0zw7htumYPqfaJ1a0TSF+y6+9tntNX/VV1o2O3BKn4NJ06TRo0
f9Oun4reGVq2dsIJOUrVXtCEWRgTPuvT/dLCOGZ6BW6xQt2gnzQ0bdHJjEYRRdBM
kmg6ECUJsCnyrYHuKFiv0z5uNLKBItwZaUv2D31u6y3uzW0Au0S85elzGVDBd8OA
IFSYnaOhmI/3EKhUwCVf4fYrpoTSCu00crYh2/Vt9xntIYuaK8exYRaMqryvI30G
9dwOQaxg7E4Dt0KBFwsN/4l6/UtxrL7fwspINtVC8Fa24QrMMaMD2RTdskQXiC/4
z48Gl9z0Um8kv9DofdkOznNk24lFYTJpQ3LxsFbJmPzRHl6xz2OPlazK8WyrcexB
WH6ZwFSpZSmStoWfp0/ToEXUbxpAB+LJQp8QdQpd5QCDDW5B6eTpzMlpp4RzZtWR
opwsNSvRhqDdmglQoRPqqSScEUJ4IPR7/jXjeLj4ZuX/fndeRXxp+e3PVVY3a2RF
bNcAo6f04lzphWXvm5n/W0VPdR5ieISdwK1NIpiicJMUTwaE8mA+IBdL+HFZwXSO
WsPtXOZ9JowMLYeli+zdcyrHbLNVxh7JVKgvwrMlpkxMByPYA8rZQK2CvBlCnYu8
cPqx6xmyDGsrNdJnow/oW9aSeIGLyeeCrxavMsxjBRvw//l6iSooMjRcmVG0h/dV
1osU24CfsUG4w5vLr5nCxpr6DokbeT5FxVkkmdg2gLVhUJXzZYPulJYdhc3woSvJ
SVJLsMmO6lCdgX+FYHuNO2bDHcxHPMhMvkrEZGYHGx64m/HoIeg1U2qLRqntEP67
wbTrrsk/HDzikcUWlNRWOqyBDWomDuwIchHrmT0BL0yK3PK2mxNy3W3UVNG4DFrz
vRK1hxwaIFz/Upq0nvJzfKNwxn/lRxmgJSJg7zEgSreo7sLE7QCt9PpFgirXCWkN
Ehmy8jdXl+J2g06dVLcgab+jKWjAl00ptc7iDhWQ/XVYcTwzvOQvchO/Njneb5x3
EzHM2oTU6pEnwrWR0Hr373iu9+w2grprRZgK/s9FDBSNt0VmQGyUGrNbHCyBnU/D
l7Qw9hYQ3J1NyoEVleJ6uR37LhXEbVwynXzAQA26G0uM7lzup0NYuvPTf9WhoL8d
wCwzw0aqMT0Mq3vMYIPOcInx6bQJNWBDNI8TbUJn9tdpnmfPtfFCKiTOO+GK8qiW
K/3U0XL6LT4cnRir+YkHveQY1OkTVHaUc8+6JRvCuoP/cKzO11ThlurZRNHxo4Q1
tv5i2vi9g1IYVqEEY3G0REyGPgpHol6dZm7a60fu+VtyzqJojd+XvQKsSuZYO/pz
U8NQB6o1oQVh3kVVjV/EzbnlgslRorc6gHfx4UPAkQC6EZg2iyr3bhWI4pozlxdU
5E/C0eL/9IqXjakImJlSEWGu/KGMQuLj4CN7O8AjsJxC//a1bg9yQkX5nBMUzIn/
7P5OWACumiMUzGOrzQ+xTS3681bbgeLYhfIm65rIKjXusoQXdvPc0YCeacRmHenF
3w+0/gUxwFa2E+Fq48IzBqv1MdlJ9GLhfBl2haCGh3/VgeEkt5XeVFiQhwD1uGjf
xY6cdf1AA3cfvoXuJr5CvoszN8ap0Dz5deUIRxp9C6/AjWgRKw0L8catRkH5WJVC
FO4y3uEGnQ76pxnJjbuflBVKr1xBnGTNRPuaoVWR9zYNMfXX2SWAw750XVPHT6lh
pLywGGUjPgP21ZaqBxp/psBw2eSCQdCx8stXeUPg+VKH1l1zbZ1LuLLzGU6rJ2wO
GAdrguvlTWUHIaNLQwhW8uwGa6uUUMISnjRLagMC/ZZQnhahoMnG7yPk5/ZQmHDf
YgTkTPI0YHNCz/JpjqFqD11SOWdLSR7Mrn4vTxko84lgCTi0rwU/40TDJvqLYX36
gS+IWs+xdtqKt7C2+LYmJDj1MUPXK+NRXu1bXzIGP7W4g3Wx5p3M9edglNQ1KuuB
j58+UrvGLEED69kQwCH/o7h8fNNchVF6nrTktWBaFqWvHeqxT1QNAgs8zG7ccWa1
1DaTWYGr3Qzd5GMoDnkuDJW3cSkjeos2mZYcJvTA0tLbiVLygj0wCPyu9/+5h+aF
z47H8nLb+8n71NDFPzRnmKNrarWNz7W0xA7rbKgR2xP92P4l1D9ueInb+lAzc7Kr
CXxhxthVLkdQ7ZxY7AbteniLLJ2CgtmfNqB2QjHHD+QHZezXin7p7n8CfLEDglmz
kdrfWKsb7Z8au0tOrMFG6fsIkVKY4o/sko/emra0ivJK8kHJ9mGd9ZHdlUriwk1h
cEgrqng3mzW+StncvOryTuCpw2wR63L61Y90qAEdaQmwcpYKmvtk5o7lhwt1woma
KPy7KK5TDG7BGTJXa2goCLjRuWC0u4mDGGW9qSUz0GTGy0BepsJMARtIriDtkkOh
8yT1I3YwyPGHwoXsI/VtwK/aHgzhhAUkTxskIemT8n6b4NPZOscw8sZPqRTsYbjC
OkBSpnqCgWBeOvCPa2bAKtmuxT70MX0J4NY7/+tc5X08nTp13n5Xdcrn2EitrBA8
u/1FoSytr9WOQP7T7AUoUrvDzG4VXSoistGqhtYJb09HzfEv+EE9M7PxMBAB2rQy
bPX+MaRPgAZL77X7DTWmOkjEL4yXTmsSMgx5Ut02zJ3DkZ3xL00arfVg4GCt2Yup
V1crjeIt+GZghrXlmHTW9J8zNi2dVbiNpSyc7PuQkHBdV9UmdcZcqIOLWGQo1eQ9
LdnxZH3U0VCxP6U7rBDgf7jVxAbmwteymzqcEBaox8DPFrQc33bNRm1Du9qOC1fz
4GFkxrn7AEhJirNwj3WirJtQOxMWKzVe/JrkBe9/zfrHx/R35sVv7jBbkuZ5ZO9k
UOqSqWOCkhjrp/X+fRe7aakD4ENcoQ0mz9cosUOPe4epspNH6m4pY8LQTIAeqoah
XhahTsHK5kkzi6LCWruAVfnfGHGwfeBr1LHt6Ks46JMZ6N88YDgdsF7M35srGQ7Z
0KAAKJkLvXzfI3Zpy0uNKMuJdZqgVa5X1U27JEaQL1wlMHkiSFjFuu6NMEwuUZTX
2dCC60fyYxyi+6v7DsjS0441lhWXH0pJkFUAgspV370T9DAkRhBWFRO4bVLlesgq
lbkMDsqT/BtzCrC65EwubqVsyrjZ/BopjyukNU4aEyhkSoG+QgbAGN2mhIaZxfah
0EPb67L5fO6ZLajlyzhYbmHaqzP8TMMs/TQfzPoVAoSr/L+xxDf/t086fTjs9XyC
hn8Pw+ImflROjgqBhHlGgAdBOkV1plJ5jsyceEFwvvUhe00qjcHeGSrRZ445zEUt
WIhoqFWkkcaCCSwtPkSg0sbYKlLkv+cz2ZcsLZt7OqNfGfO5dtuEZuUQlU+Lc8wA
u54v4hXgrz0cUfXYVaqr0pFh7c4w0eukBpyMnazE7Jma9AvsUFMi5pIoNA0BjHNW
Jk89RRM051QtFA4aNwmQsaKlIEKyt3j87ZCovZvIqfgNFKdECMruXLPzX0VMnLsz
ig+c5AzP45HZP6AvlruwUfoyD2W5BhQrENOCTzYAma1Z2+Kcg/DiD9GrQtJFjsE3
hxGyhOeMy1Yh6Pdsnamyd5cVbx5JX9TJhdPh/QCPeXECfjXCjjXRewzfCl9zZvr1
UffQPGsksNjg1rrO1ZXML+dJFwkhpENd4RPgD7d260cWP7wjfust/ThbQGzb4zVp
XXfrUnb6sENTUEvjMmgSUF8b7V48ndDKEb67Ndg3XZV5i9rOVW36lbIF0oc/ixvr
ahgrpBwbkfILUq0RqzavrGlRArNnMYIUzEE6bpezf3tPIMGVczzmnkH7R2iyc/Lp
x6lXOEVPcuN8T3crE5lZhmQfXZdQC7gQDJqLsYP91bblNJmbxhuZWuvnAR7pLEJq
+rWNcRrnYMHMvKwtf/gYfCv001By4oqpeEBf1iJcMaRay+UCvD+4bIq4ivKZOTdP
x/iu/0c+9MojIcQWeE3Ht+5A+PiGP4LeWMEwFssWB6Irj9lWtLSRi2xrzfy8vZqm
zIU766vEKXPaF0wjQT7YVLXwfXT/VwKUp2saaWbVQFju0NXDDSoKf33RvFYEUbhX
eLXBt/GsmBkI2o8elZmLIpYM7gkwZLf42WzmBWJnHHad8d0DEIUAax+4BbFHN073
q9qPNC/iC3VR25F7vDsTTj3VaayEPK5TN9LY6xHHWkMC+EEo5rSQXb31pSHJd4aT
t9fWFU6HGX5l6b6C/JeFibSZef8yQPwepFeGBHN2th222XNuYxUioNak+zpmqQBp
18UZhkMvyEH5jQMotD6AfChaxkr8QF8gZG3n69SbnhWT2Hi057iAexOE2xvToSxT
Dx9wenRj8at+j1k7H/cR6dTdGqmpromSFoNicmpiTnCvFX7c7j2jENzl+wcmzhkE
vgfL1L05JlMcICjW74oNQGH1JJ2UDELLue374uSIK5/qa6dFMNzlCG9yQKAyWMsg
YLrM/7FUl5CRkOInvk5xBr9qOIokI4oxkiSQOMgzGPXgXKC2Qieh2F7DtyNTxclU
d7BNjz3NLDyx9n9BvkIUDWxfRmkVFwgGB8cwaA4qrlrTeEpWsok/ufJhTMWvnCKq
nTmEKjO0oZElXZ1BJzhA+4BTeJnaawMmCrAlh3kCRR8B0nAuWTlnIaHF6I1ClpMn
4bH+ALdlI1ib+DCY8ClmL7E/yE5ECDpzrRonhymQ81+a+qMqDJgsXYCi5h2Shjlx
2kYr+VECbLZY0mZuelw2a+X+ajKpsu1tRB2qsd8qGae9COIqWij8lWX2Pw70mK7z
oMTS3FslWKQN04UjLstnoOBbZwl+TZpxZKZJamj58U2bZzPe9xrxmGrXCxF3m3Ez
fXGfw1E/DnyAKL5E/qmZoy/CHmmd18rj2jDLtWVHDyhJUTKPn3O0hz5x4lVJqzCT
Hacb6d1ZbixFATBAemZP/Jxpu8A9tXj0utQ5itu5MEBLFdGpoRIbTgWfbWhSAIjP
RVVEewzzoXzdy3Jbc/Zxks04y1S9xE3iELV250mdhnYHo2VVMhZyWE509XvX2Jbm
vN8gerGWOy7MBesxEGVoBV/pjtQJQrIEpuknKB2qqZi25+cNyObPG8OsHvLwQSOW
R3fXRpwsqmsIWSrLwgwqXPKiWeoKnKRk46ggKpn3VlAaIIz5m94OrSywU4OvlY9E
wZ5s1gqmNfHfEqtOWtCEQ8T2HLWkow3uqfsR111Rx1PhljUyQXr9Qf6nybrmAuXu
b7bnn9cN4Y6uiP4i301Cb2rHI7BpTgJ4U3b1i27VhKVdx0xTBnV0tODh9Q3mjSUv
z0Od1Pme7s6xF6U4SP/qIRN0k0tgiRZj39b4gSEt6OeQJkl/wLEua0RcumeVrETt
tLfLC/PEBGsaTal/Xmf6BUv6thSo1k7uRRZ1PXDwrASa3Gix5PAWVD769jBT3BLW
k3JyVWZjW8bE/e7eOROOj6h/bb4wr+wQ/wRA3PDyPDuh8h2Xn9s7q8ex1Sg2XQMP
z/LIrUa2qQrpBJjZ7tfwfOHXt09oCZsnh/1RWl58Jk8Idnn/Msh5uC2FKtGA2jyj
pke3ZtetWI0IHWHjOqy6iG/SectDzHynnLufIXWzY9pyPp6T7BpP7X27/G7yMEA0
44jfNV0Mk04XOBPsx7D/ek6lvxHbOl03cnCFF4qwomkUu5tvlwYGGS9Oi518TCL/
E/ml4Bu9jCpF531M6K4Tm2ExP/6qVoSBbdzKnkR+JB+8r1iIzRyD8raTibKpCbVS
G71k7EYC4UoGGVWiAbQBgJ8lp7dtakPcZ5M89zfbJAjSzLuvl2NqP3iNLG5V5/qD
XtyQxdwmbgzbB48BIKbCrKmdJdr8sziNKWZQaJ0IWWewK7Jgau9P69HAtTKy0gT8
sROe59xoOQZb0lEhBHu/huWsypufEJVPZkjnSg9iqi1m5S0l1K4UD/ucQs/gZSLx
mJNNiGTA+J5V5FQYdr/iPQSiC+ur4aCmnyUaUnkbCtvckBNZ/9ER43KbadsZ/5V4
VXodludjb9XN1wvd1lOvwKgHbgl8W+G2BoiZ8TK70jDXQ3kFLlzeW3lhxzQvB86O
S62uhpFF/4eJcGrkrxLlYMlqrunJC7MAL5wieX0fVUL7tqrGFVphieY+LnS/RkMr
KPq7TVyQm/gHrgJTSDDhDtTD2/9IWonbnKBEuF1MR1MMhR2MHuMaBe16G8i38mY/
Ld9oXiXc1hSZfyTIAto3ZuNu3HK84hPlwyWYxNoblpFEoq6vhLYSWm59ENzah+uh
LAwlG+dThzqMxzcSVDTpUkXKBWTcXSFPHLKM4/fiWBYl0Xg68+lQcMRKW5bjsdAC
6g49BgiwbeRJPlezbq3ulfxLTvqrYPNeIHvPk+xc4VzZYYk5ht/JHWN/IX+ASDzZ
ZFU4zusdMdBPH/gBKWAYy4BAMDXyXoGiURlJ4PZ2kXJXiozwcA07rufd3eN10Dhe
s2Kaf3hZs+5yA/TNfLHDldIqkuHdhw1MGmfqi8LZi/d6FECK6kl92suYMh0/sIq5
EQxLtuItPjf4oBzYtUR0vrQxSJopTpn2qf8dvy7e7woDXMF1NjCAFR/fnoPNezHt
JCA/2S/pZyY2ZQHlPh9aXIe1h1tWLEWDNXDgkfMRA0L3LnMrAJg9cuRub/y8Byjm
MldlU6RiFiFAPjlB97tnEWozcXplOUv38aG+X1XaU4YrV1Ks/1PaesgyyBk3ifMV
q1d3QRVFYKPu6Rq0mvdLYrdH2X/S/bNRy6LJDfwMeyPKcrQEclAeMLdx3COCSbjv
UB2TyM58L1zuV+VjyM91y11vqVU2f0LAYLfnBnL5veV3eg82ciGs4EQmEMHv66Mv
gs/w43F0o1i38+f2arDdkvV6F/udLbA4sN/PPMsV/OeE91PGgCcK0kYAc1OdbmUD
XXk7qlSaOpFXEzEOXaOVT09oB40Jh8CkD/eTsT+Q+ll9KUmQzGRr8Qk4YpnQY8By
CSKxceie9Y3N5RX7Oi3SwkH0r3MM/efnHBW3Vv2cPd0kD8N+D78+0f+xYZdH6cio
5QiV6ilp9YViV/ScHmFLdNDBCbb8yX5+W+0/dUrOm3mV1xnnND901qW7piW0ldZN
6f21af0I8lUzhNbG0jwyLvqd2vTZBXVd0i4P1uMb9vPAPssesdpuIzQtBx4jBvvT
AzYfajlxXlSzBnNtN/7E/Wku/O0xAOj10IA2rAkHrvNsu2G9vAjt3mepX4bF7LCz
+/mfMfUoFzO5MaA6pHM35uyybbDauYbWC2fG4GIMWAan5iPJL5BCf4tbnYjTDCVu
HFGRS3XdH4UF9fJf/JfFtjcjdPh4TpEjwaDGgJ8HInq2iSQ1Ke6uQ42dthrNS8a8
jgLD0v+1Jv82Z2DK8diOybKDOasSkU2feNi0KLHcz+uuAPOfsA/7Cowm8SNzCl/6
A3mzrchMmS1kE9xbfE8UUSj+C+1W7fy4T7uSA7fTUGGha9XdmWsCooDN39sgSAVU
cHDfVQFd/EY5l9GILbrdx/qzfID5++MsNlUbZfdWP72P1etSp9gReVWWgtiUbaTY
z/vS2Ghh9erdzhM8KesG58RwwLvIk2xieAL65A1nj/hnDr7h5aixu6YeY4Q+KBEy
YVYJlDRc+X7jI94sYT2qn69SrjCnupemBZpYzKPEbueuick08BNDx6EFYozcq6cD
zrYEEnSRVcCtM7SLtW0pkYEgneAZPeaLbhO/zIpH5iYBmxVeJcemIRWS0oy1dS7o
/MzSJkIITfaO6WQIyEXGwp2Bi3I2zmXgeWev9kiwWqIREgPtNKWWEWzqLXl0CvLx
uG2nUCHM+6ue1KQqD/oGhFTI80tU3x7fgXJKU+kdX+0BZLXpBnpIDjtHKmDchshi
UnOH4g34OiavCXO4/1M0pw/G3EHMSSJTQAwk4Ty+CEErf3bovfXWyvWFkQZsv5JI
vXqZ0XBB6X1XXgnkHf82Ivs7jK6N9o5n/84NJKdXk1xE8dTSFPzCRuevEiilXPbs
xD2zRjCsq48Kos2hq5VKRQgNJJ/9ZZSN0YTHwfdjjyHNul5ZxSGzoyVMJH2qK24d
dR+R+d7uDCxrl8kXsuFM4n1XYQWmm44j3RSNJyr5xzDDHYLd+4vDr4SLq/QUusw8
Rm6abrfG9YvuR/mb96Va5jBcbDEHfYzUE4FLuitrYydSpWvr9FikYPdi1WrFbdjA
u9syhLR0E5/kT8zR6kI7EdJYuvizhs+mPV+1qtqYMRzC6eFbAZSy2CiSgXlQQsFs
nUYcbZFA6fEFCF6ENtF9I0TxckUkOSxnDDJ+xG12BVVdaBi0a8L1DIwulS0qldwq
rkXmciSmxiOYlvTsOGTmpM4H0YsZ8uY/L60RUzqfUW0h+l8TcGIYywGRSVO7DQ6F
bgEYSGULsLG6BygV7kCzS/hAOkw4VIMXhf4HPAcXjMrZTIz2NijNeywo50wihJgQ
CDqEfVx0pKXelZqmyOyWGjc/So2g0oKcUgCyPM5OdGDtpM83zhV9OTCkuLFSwRxG
C+ZO8+YO5XkkvBLZBXl+ml2o0nAxWSFy3XOgYWfaJRj9WweHXI2bBn+Tjpoy9Y9/
/MWoaN2eMTRaNX4FW7n76SMO+cQXU7GxaWSbx/qpUqwpu8gH+pCqhabfCwWRxbM7
lPiarHsn4MCZEyob+l9gA9D7mweGf9TKgR5Lfg2JhK7sq1i6Y1jNyYtPNUTmy99+
f1PCn5JJsXBxSnx0j06VYCmy+9l8XUUIeNII2N9WPyoJFBNqEPMpvlETfcrY2n+c
jOINRs7w9l1GAu6cyiUMveZQ8ryCQYu0bodCFq0uHH07w1J83ZuPrjKV2MQ6ZjyL
N+aWMro3tx+pY4c9yvVV51+fQCgi4ih7BTzim54WYt3ej3NkY/fLIZIa18+FbfDf
gi/i/ry3P5wPluvk3jyPi6BrQnBqR1KjNFcxa/6abFWxaQJWQqa76+eOjS0dkkCn
NflXftzA9mKCPYG4bbSA0HKcLmWHsaNZ3VZijtV+ZmaPUrJvkbDfVYmsLmUzxmY5
PF4FcV4WerTCL+pehDcBaOX1Bwm8cT0tnAdUptQTTdmUFpaYrLTlcPnBm4hJ0K1/
A6zBq+nTpH+nS3pU8gme81VRqH6vlW9rCBXDQv6avnH+WebVJh1UrYGZO/udKmKc
LL6ngx54t3Lk1qV9DLnVk+WRlmWX3dZ2HiFdKuztseqPBoMa377jt8i0qwe5yrQy
20TOGm9nQu2vIBmVoTqqP/ZFJ3ZdeEsZR8NBWSQsmIOpPzTt1IqHdafMNCc7O/FY
Nn94iPYIjTHY/o6bT9ifHotmVfhkrvQgUACcHx+MTWahOK6pwW/Xkah2iAoxfllC
0nfJg+QV3VYQW6TxlyYtt0yRiWKzdhbMncg9gLXbinwFjKOcYRacT4meQOQ4gMcd
14ki3DcvxkACeJMzgcG8wW5+VhgwX1RfsBgLzIMSOECdOEoa9OArDmG7BNhxDCFv
1rddIUH6tEA8l9tx8k0ypUHSwCIQr5iHTNyakHT2lWsMvcG8azWuHg9TRXtzbbJF
ETj/hWLXQqdBeWwbxJ9sNAbKwOw3G3Xi5PUoPq95Qf6WvF76aF8whRIVefIxxlvi
EhCFibP0BWELP3rKx73Kq07iMkV5zdtqkUGyXYzEpoNC5PUZ/vYoUI+izHsDaosl
TB2vjI2hKxpSw6Kg8uN766o5v7MjjSH+pAc8A87n874hycrbD1D/MuHx6K1A3ezp
0yzeSyQbixQPpdXyOKkWZ4Q8R1IuSlKA8TQls0PBL9meTFyHAINpCG9mkznhPgEe
/YydERnwSYukGoPHZEOFMQNar0zjm1PZuleIJ4jpekFUzajAfjSqeUpvCD1UuF+R
0OM6/yZf6S4+x5BGevnEmU9eqd0nC8fXuWSqiHl+aU/VUg5g3Bry12QSCqXmqmsG
lS0iPsA73/vpgdE4K6qiCmhXdlxxP2HEw4D8buT0TBa9QLDnh+PR3zBg/0CuOKb0
KxOkI9UWEYvHBsIN0uUS5IzMPg/JGh4mrxF08jgIKEsWVCr6JpGKgjUaB8LFMdIU
7pmD20CiEWf0doIZ+TIC9U5Ke+7BIKjlieTpbBq6BQHwBnagGc8C5RL5zefjdFpg
n2Xa3AU8qP4TgpKzs0XKgBXrlOT61I90UTuTVvKqzYkuH++XVomusj10LpaHQTpl
STRD9H3XPerSwZ8BKrILDu+EMO1c93oHisL31jguJVE7MS9enjzmDT9WWtXBYCEX
2UMT3xjENOKgxJbmbGIgOEcCv7EzcPZd1E+yOaY529P6782ME20g8CWMNdIA72TZ
Qatfs5GHxmVH6/fgZM7w760HFROrhD2DT4TfDWILCibgP33MBROgpaHnGZbiEC7O
klL9Pc7hueHssL6dtbVnhVi3a/Jop61/beBF5m+Uwj6Ww9PmdY2SOFKcA20to+Sn
F0LXSbtLiq8YbkaQYtvAJfUtRuWA1MdC5eVSH84HB4w6PyKNUFVYmRcXFjGP0hvh
gUlbuDR9M+O34QiL16tRUrSa6PtWekzu1p/c6q0u11jyq1YdaZ2dWLp6CWfOXUtK
fkDLaRlRH/2tLYu6cPb2qtKX5iVY1i5EwGHfSpGNxVr6XAjEqprLWxxztC039LLL
mrkEM0nB9hwBUENCJuA4e/zOWJmZ29SMEZcLo5nTYcj4cHq0qF4JMDszFpBqAWdO
xuQQeLovW9cv8Db6XO7VQC6OAbInsFqA78uPXxsag43zHUmfUZejDzlsyrY8GXyQ
QHAe4xPriYtWW/ktYFunscaiBsfWj2+FoR/PwsGoShYCCni9MIrUbPvDq/99Muv/
Z0ib/5eKgsnxTD356APgBhQGrpRdvhhK7MqN2Bxf98INNH5ZBItFHgZBD92SFZ4/
j9xxLQ8RzKxL7Vq1UrvlP5jzlIhzw/dBHQfQdZzJVqd3qL5SNyqP1IgKQwA7rEja
JK258avjIXpozTUL9oyJWXqrRh8jwBqkVgJE/npDy6hWIXahj+ZBYLd5a9/kY/3c
ib2V4z1hcMQBkFiCxC2DrF/3Xsw9AGt7+qOSKgv9Qcl9qsNX3hzQ+jxAXgYFn9zo
jopFdRaeLM23KsLs2KF4AJXr4XolzIbBcPZrlGQrmVRVsbgpcaohTucQlmQc+QOQ
Wh2at6uP0wMSAnOabjWPeiWEx0vnOX0pBUAAPNOnOV/O4u3+CtOdE8zreCjBIEbA
5XgAStPr87kViPQmorN7HVrPUVP4afVOV470KlmTB+41pbtYuxFldBghNIh14HjB
hlIy0Yy54rcXJYlDX7sMkSOxoK+Sg8h7IkGlTv5wBcjsmWzXlxfyqDqIykk/eZN5
keywEPFsinB96m8MN1DMcDCbzG7MkiCgtYjNvVPI1bkilpDiB5qG82CsW0hwIzbD
3Ml/z5RnjGmJDqLXCAyzKDbEUUu71VikGEj+D/N9b5OjaZ4UBJ/7V8XJoWGm7iHl
d7rffFXvNei+8ZTDr81os7d4ezqe7kVLdxUQqlhtTKJS9EGaxIx1QJgG9D+YsixU
yiEwlRfQTXNXwNQvSLtSRIPGyzT50udjqMLGtx/GRlCvIaUiesmfOO6RzrkWHcBM
q/MYdJeckRlmbHFAsK8BsqYbFlzpij+2qDJFlqIaozr9UWPiNXm3OxjLBj8qSjgd
rO1t6mVYt3Xjn44fameEEwwBeqo/eHKokrvVHoVNErVPk65ctH1wEmW36oIcR6SX
SqZgl6u7QOB4jw3ApvYGJ2o1xdlN+iM+w0HUbwLJJ4MTJpnWrpXGu9ci9eidnpC4
b0ODQjwOdZbuwi060egWEOU2LKWZtLK6FLMF/oGWmA/TR2EEWgeo4lBhio6ctljL
z5SDMuvUpzLFUX6JixyyCJ9Hgn6eouFyBmiCKaIUobJlOiqcNL2VGLTHeUj/U287
OAda4GEVJ9WEOnnUX3UmdvEQhyExqk+6uIxyBrNSWI9+JaziaF3zT/NpFN3qs1N0
admC1KYuWDBy7Cexrnzxqu3cLt68dHcMYfYs637grZTY12triQPaWtZcfKSN+B3j
j1bhVvPXUPgPSsHQdpsM7/Wpv/lh/24fSrajUbo9eFMYnK9apm/2bJc/6XAyxlb9
V6f041pu4Lgt2ZvrcIWaNKXZYQgpDpLN7BH0yrEH/sZO+tqGWkEniqMFZ7vhEeb/
VmoUksR96sY2RtXx1Llr8MNZ4VkrB3fFBTAJmapo6uk6oY1Oq4/rXkdYcOBo7dLF
B6t3E+BZMjHzuyvNxdoieqkbqM5q2zGwTKwygO3zZmsj3GFKQIzaTDzJm0Pewzmd
GaFpmpC1RnPpiwO77ebbbhhONuZAf97I7N6R/84/BNpRklglpZjAuEcwrpTwEWNK
zPeF0QaxVwW2GeTiaz3amxQLjJN+rHfj1uWcTncAB7Dv4p7XgiFaNZ6Z8zJ1o79V
eMztZ5W5DWrf5LzFzePMefLpVP6IbQSvD6mQtGbEpbpUspt70c92ZY1wkm5GA4ZZ

`pragma protect end_protected
