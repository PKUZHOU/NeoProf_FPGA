// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
hGu5l824n5as2RyoU85w2exRqX0Y6HGmfMHwID5gweorIKfeavGtzZo6GGhQ
BsVVYwu7Ot1B1lS8nhD3dwWdn3i8zfHkCqeXeLiwXwxUnVJ5wkjjKi82p1sd
dUFU44Y+vAtOF0AlCb0CXUTsJ1GSKSeNVphck5OZ5GRc+YUbI4Mi6BsA6Xhg
Cdff+9apO3ZOoeMW4VV1IWoeQ3jWBdMv+ao/E0K5kY9rN8RwVquq/HIXe4+N
YzIJ5qNJ69eadfvr38iplvacmj5z3KN+nZFwhjHaPEk4BEbW78//VFR9EUm1
EvL28cWtyDP/r7PIqnnG8Mz5o7E4zG1WrptP+kcvGA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
AZJMj4t1NHc/M75u46jXjTnGs3mny9ylijKQy+2tDrq0POJoGD2YOBGsNq0H
3cXeW088ra6v9g8aFLPNEqblDrpZUmn+AZrbiQPAlNw5RMywZhfM3WxrIV5y
X5Lc07wmN9gKKdOIBTrGg91+LMZcLXNKcRPKupmn/T53vIOSsxspHAH4qd/e
2jO96EdVGLGHLJlqTvzcqBO9gGSJmCNjv0jmN1fqS3Jwb7mRhco3TofFzG/e
WHDO0UNtDAQoJOtIOP5gA9/IiPGrO37Q9HOzYxYvtDLjMUKAD2in5PkceNiP
HOklQQuGOU3W2b9ayPqaZ+Re+d6slEuQVz2sWl69UQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
P2M9itg9tVxXjbdH1MABjOcY2k7UlnhL2o34UeX2th4/2TT/42We1GlCve+c
sZUSo1JyVzGLuu4FrN5w/Z8SsdyuflQnAlrKugsrsFDOWDPx+V4GbSKl9Xix
51XvyxP7n+tYvC8Qb1RCoVHwUYWChgvpr8tCSK3ZrLMA8VBbIcwXf+Kz8/sl
gd7s/BSsksp5MkSk1WstfshkR5Lt17iOAX+bexTusGn5iTLLEGiO+F/mVkT/
Zp+A+poLJcj/DcPaa8C8E+wS0+kkOpzr2p5ZlxhAMIostcdrbGJ5E+WW6ase
JtlaDcYRjewwzcf4VJhJ6Z8eDwVhiHo0ZwqRG/UEuQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
KjE/jot6OUDXFEg1deU4Q8za29m9aTVDC09NCoG9AB2W2VD7BbAJs0HYhny+
gellgckPlJ6sg6Ia4KoZA4y5rdySgfEm3hRgPyFOYUbbFyd/MGdbn+qcAxw0
rKcRFR0lPyj0al4bCWRHWMSXflCFPfaBTxmCmonQDt+ShYP9+WI=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
X8Itnb7fvcnYXTFv8vZtDWnhQoYxQYER+44b059/AxTa0yxI148SNNciglFZ
gSVVUnJUI+ZbsZbandIGd62TLPspr86up1DFGv3arPwzpshx6NH3XVdbHXgE
yxGpQiooH7EctkNwr7LZNAQDJIxO6A5g+cZyA7BgvrWmPL7fjVfZNIXcbn/L
LlQqRuQ9HKHf8C+sUYFhBRDMoeA6XFVmFIUjHQJ3k9RqDtMCLAprjKTsKX+x
xlKwr/sqIoFSZwHikMvfHk4scOA8Vz6y1hheK+ACQQpnolTdEmyg02UjMGHE
h2SVkG52Y105OnS7DTFs3iSSzqU3ypVTG2arcAgJ9Th8t/+3tYAiQf1nsGYi
mF4jzDphgT7Leh8Erplz6Mye4MBvVp/iILTvPZDwDBI/ONK+HVi5JqKUjg2W
CzOXj8xQrZ8lZbRMk/5MkgevlIx3M5mpJqvS5fL4/T9wfKu6HlLuwFa1dJPr
hGMysDzuLr1UdEIJ5ZC/jISPl1DN6Sz6


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ThBjRteL1S5jklm2JAugbLCDUYqje7BJOncKsI/EDVxGdZEZ0YG60erPXmzm
0v+OQsJxYFV8BCNb1s2yhtsj9lLgCA7t8i1KZ5nAMlZV5yvzj9TP2s3HRvrR
eUn/KQ5cTiiQ6SIN6/p9y1hONKIclpTma5+uqKU5v3W6rSOVUqk=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
fhRalrsWnu0oUp4ICdlSQQy2o25VgAgq5oIRslLEwIBnGq3GsdsTbDzjYpgP
LIKiwU54ZD/HGPeFd5Cbtxu7NEqK7toOxQ/KlJXg8SYbkIA9PmtYIoqI75TZ
2FGRzm2CbuOvin0RvvFHKchEajj3av4CRH8QNDr0RvCfDW/7QB0=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 55840)
`pragma protect data_block
z3mOdfHP6tS7Mm6H5pOVeRdlsvozOkqocGhJjOo1mknP6yo7x4S9/pHXkL7h
8cnj0K+DY90tc+X7EXs4tdykoek5lt/2M4DokUqc41zq/abEngeZtiX4k/pq
7unbNCRvw6hShQzbONCNFp//BO9dhxHWksFmeRFXrxRwMvf1U6bYgEHasXjb
oUeKGUet1pOBD3eiSCBdXnwEevJXNkbn/CIIShsrFBdMU7gjiUs2uOMn/JNn
ct2ikkSC9Bip6MPt16NIb2f9vGVECnIzhwljJhI4oEPAtE1fvfzzOnFXkR5H
ECrnJZr0KiSC4Jmnj8mLgCc7qqYX/N1+TkKdicWvVb3ho9g29uwX4uv5wW70
DpM24neFaRnjNx5SjtBZbI9Q+Li6Cbye2MS4NBZcM761sFB3x4fEFoofLrY4
kHpEWDWnF5COx1WL/8BUeBZNdqSYamr+ICPK7TlLn4YwQoUEq4cpRp8fWhCU
F6CtGnz+lDNvKubM52RoLEUpNf2Lp5aT4/fiEhk2wpWKb78V/sPbB4JfCIMf
uGH5r9wPhYpV2I/+gT6r/my1xsZb9YKl+NHE5ZILAyCeSR4aUND3BndGHUCI
FCKVVUVcqBlYsC5HEIrsVnRvEXhVizMBwlVJT7dfPv1eHgn70NmJe6hN7rlj
2pWrOqmixrLdXlQloS3HU5+xUupGvD7uc+f+Tl5PYMLDC4yKLKia6rHJwLIu
Yd+UOy+Or+NPnNNWzxHc6uVKZrJckt3rKx6jLAzTf0vkNTxdWTlAFcd+MOzW
m0RvYlHQDKc3XMtzO/50V4COJL9k8TDhh0Ofc+V87QB8JHpYAqcAxdAKj2TL
Av8lvCX9k/LDkXUeR56HN7XUM577nr8nkT0T1eVye6DnTIHwFwwNWam//hUO
DxRRfEGi58oYiffuczjdIOB20Ycd9L81Rzfu0tXnivGJeSX9o5SnQz8e4F66
JHZi/1VpnZASW+4RB1YJwa+DzCzwck1hHyUCqBRRXtNxc7NEmOdF6qzjhNxK
bmI3SnMJbT2uwF6g2Kxq4zHTujNzko0O9W6U2t9Gr6R5eqbZ4Mi2DpgykCbc
vBp5YxuVnEdZs94I3f2SDud4x/8zCiLqnDnFr2rgfVDSB6zEmvQuTg4Sbwzf
PlimBtdF4lyra2S8yTDuDwDVDo19Tm08dzKL7rmtk28Ep+z0EkEbBV5B12pJ
zrflBewFf5Y0PNRgqt5UMu/D54kdsNwXfDVMFfAyY5+RRV917nbOGXFwLhMG
yEWJHqQ5JIqEsniuT+LF9YlLygD2CSTIpEaSCwXapWwJxf5PHKqYCsTpGSvP
405hfqdR1uEqgMmCbr2h5MLT0y8FMBA60PdOopjCBrA2lNOqBz37IFsiB59q
Hb/d18rKJsoCQBCxnTm2vTVZx+MPt2vvToROtXr0+qJigtEFlT3MdwRictuz
mZiEpsQLgbFffYexGdWIIp3y1QYFiedgLgQafPJwrxXFyWclQHTEdNUkotJ+
lJRssaVPiwhj4suNdgVOjtADrpMHKOYZERqhchDF8wzmX+7EcQaeTQgY+FiN
RUMa/l40LDgkDj+0hKLUORd17y0NCzl5pt/cJPwxoIBMrX2QekHUorf/UpGx
DxtEINwXPiK2L0kPCBZPW1UyO9prdjRsIbnV80ZJgt6hUnhwDOyETukW2GRP
baNvjdn+viIHHPb9xlFIT2UHVAJQy5mV0APucet7YP5tyM+PHm+m1Kz1oFT9
e8SHmuwatFs9bpGhiUmtrCk8XLDgKAFn5uvu3PBlWRGgtNo96UkVvM1zZhOX
dCLewkz0+ASqe5WNP3K/djCiZjg3xxOf0tMrJeWh/6P+wuoJlg/DXkGTn8tG
1lZa0PgFkKYCwOyN46RXpxsrbyxGVPABjIKQLxzmg+lrbKCJZIvVyoxz43lE
Lr/qGCxDPdDW/Rp2OkIePrgxf8715IsLsWrzpZ3BXUahKpdqOLSQtTcm0u7i
TH2aVOkLyv7MS1vEv3v1Qs6tZiz0SBrx5ip2xHSc+Pm/SAXBOxwTcPY8XXdL
359m3xb0O7L7wf+AOJeDxyCwh3f3cGyUGrCsVUJ39IMLwqjFpdex6zFiKeJH
h9jWD94L95zhbDuB0riuq7A7Vz4PXC+XR67Teuqj8eaEHYDWgZU217sszb6S
ysko9ScOl3tHDDB/R4NmYShEfzxxJ6If9b37rCrgulGsFjtOABADcIigrRxU
TkphgNbT1tc5K2fc1pyxNsXZypEmbgIST+nak5q1lBoXRPraYZePCX51fdm3
bL88G3DkCkeSC8ggaQV76B9+yu3yBB808ZgLEh5CK/0RRCYBM3iwc+swaFJk
+Fx/pn6lqxVLbxZBD3WFj3NdpAYeAmo2VxlNyTdiF7/+aNsg0gV4AHod00gZ
xvIqwUXArniF784CLj05y2o5lJL73uNCjql0b283XP7VtwHV6Gj2ipVJfkj1
1ydlgEwzbyl1FFWsjvdwr+tQ6VBUEaAQ6dtFuAGyhiBvu3NmB+Exhm8WteOp
4F8nyqP3gL9ikdK9XoYEee0taa3Ma/8Zyu/ZtlIrH3qbXAVypDagLR2HdHpD
5BQijDsXKm9Pf0plgwv5y99+R2C2HGub8rY4SuJyBfhyMNU6+e/HTH0TS4Ss
QXtaJijzwn+4HKRcjZQJeueaI8dNb5oY7T8pSwhgoOW4LkeU404EvakTkpDI
bbyU7f/f/bkQ6cJJGvkosvluAuZK7/9blhCwjwELE7d9KqR6xeDIht+UXhFZ
K5gqx8XqE6v77fDekQ6j88LJ9Qsi04XBwFrcnFUJbtbdrUgZuksnXKJ3sbns
A8fu41bl2jn7VPCJ8pWajslz39s0PhYWmeEky2qcUi8ZvZFHYD0vryv1RJyI
SiH2SVdEDGWK/WUBNs8nhlrnS1SKrEPJtcmLs0Pr4fTBAYKSZkrfbYLsIM72
SAcJ6ZgoLBdR79unrenWYP/7YuvNW9VPy/qOAnEH/mHXNR/MWxmU/pkNwZy2
UNJRDRWNvJedyOwK/b058vywaRN/EUF8CqbGpWxsNqLKs/KFKyJmSxP+msCR
2gOyE7lD+Lt2iBZtwWH9npz0fLjRPrjowemhSVHmaIKS/QZAtsIrhJSYbksO
WrQrJ34ScMgV7FZJS7yOZzK6ZigtFw6T7JGovLxMkvYhqzxtutBLVmXC9Pad
nV/aICpGKj7ckSirM0UKW0jqFk+l+cb7Vhk4uYYwRhuDiPZyHOkIwiMab6nK
jJmvW0xUb368oFqT+cmExmCyCHDbVUs2vysEWIFxP56pDyVVumjhMxkkmwFW
IB3kZytQjxxmXu90BcTiIM4scFtAe1jO2AO7f1uHgzksHKvNrJmqiP5Zqq6a
966fe1zOyrn9oybD3rtpIrAujEHrdU+BeaHtgRA6k5g0ToGHMIYbLFZc033A
cGvltAfHfNYNc0FT6kFRdSj52c08H6TmJ4hGHFSnPFI7hQFjnhpgJeMGqk49
yRWkuXPUdSpCXVOVBhcX+MrHlEelKkIe0qsZoUZq3ZDybCyyWHZEwgPQYWci
gNp4zgQLFm6gtxa03SgAnhh8lEFCVEGytey1ic9iB16xrdHoIxyfGG3IyryD
oq6LqAWAvhCoegiWHZDTHJsVf7Lr5tRQ1Fz2AkL7N0K1ZfVacWUDusdecBDi
JJS+Z7NDdHSarzvOPiQzYhZjukrT9AlzZJPQf4ppK7pbU5qgsI5YFMvloXgT
wisnSggimKjE2NRuah46VgZndJR3UZC+Gk9Uw+eevwWlTeHBkoR7TxsF5mOZ
tEGlq+l5BuRlT74kd0nI8LI9s9YnIcpVfPHqsO5DtvfsIxaTh8rFiGcdv6Gr
GmDt2V2rEWQNqtTqkROF3gJklNd1ozfe8UAS4UzuRnOjugeUfOTyDK5CUvXM
RTdXsRk7T1QbUBwoFNjgjKc5tmAuczNgv8DVbYIFOiJWhqv1alOdfzKmYE8W
vw6VOGLg49FkgNy1oUyTQsGBgqFdDU+RV3h4EuUxdzdGIl0gCk6DSKYY7E5I
o2GEHTfZAITwfH3H9ElhGFU3MDP5LuKEipcDJYuQOWpCiQIU2G7KLcgSbkCx
kqfTbknubVxVXyq9vE2U25TQMijHtNrMsVWXrkE8+mxze8VphKhd4IYbNFjo
clwdAxybTnahgFnyq6IOHhfHcfz557JFLJZtT2MlLY9Tm6ijePxfnfFmPi7L
tknaVJqecmx2nJeV79ZTaXq/M/8q3QgWWzNjNZK9djKVmeUAzxgs2o+X93Bl
Ry40TXHJBXdRyq9xX9zUdZE88jIgEOV2gnStSqJOuuhmSGJbn815F9AjNjeD
5Y1kfPchyVY/ZgQKkd4sazdcBU+tdStcJYVt3jtCMjs2AQrrLl6p2ZVVBBAl
SjnH+ePnZgB8l3J4fGKfXJ5RxUsuzsaJ45i9xi4u9L9nJSzDIxrwQNhvHNzm
7z5uIiqZ++QNKUnFsbw3z5SMC1/R31+g0HbiYT47DnYIYXIS31fDgWJoC4gX
ufHBK0w3mVdWKW+tCmCriIf85oK6tC5Tc0SCWgtoDelTln43NVDfo67PZjdY
g2X+KA5MGbrmK47KH0H0QgkWzKEJ7Qv6K6x11hYjY2iw4y6V5ZGrqBfavbst
j1nFVYSwhh76sVGb0W3yt1+b5kI9VH/ltF4gNOi401fGYHc0dWQimpIU+aK1
vPlU55uWFGR3Er0LMb2KarBOEtsFOnUUSEp91msWiIV7XsAuXab7+ZIYMuZx
WIjHMerL7fbb6bgwj1Il/eJn6mwm+ctbBhYDu9Gdqa51wiFr5XrIbufqNu47
2MrDrOiFVefU2mrgbIC0vAG2N9Sk2WQzdJT/I7oFcAb0yMT2IhKxST2oeYNq
6var+OkCAfbgTq+7lisQpuoSW9XHTlV1lXwrscj++j941wsDVZh8zTNYOdsU
k9rxYjNlGh9XJBq9LIaY7NxsPbFs6LwWNSYpwpWAbF8giU4r7OFNTy3blbMS
zG3TwHuknIwpzbdZhEuxk8AobxwSJsQkuXcSQtVG+jWsCb8nW9g8Bu7ygdEp
7bCMCoHJ2wK7//25qbx0fRtS0eZJqlo9xW8fl+x39k6Hd25DYEuUxUBGp7Ik
hE4UzEw7oVZrAV+kZYHQvQAVYbU00whDPu/Fn/dAyYnNSFjatEJovQLwC4hb
BK2JhWNCeMql0SJrOxCZW22pBEWq+jHBTh+/fCoPiaZ36HdsQJXH5Yxp1CCp
tymXcIWrTaW9GrNfBAZ6SuuG9exlVYa/cfDA58w6bfYNwkmUWC/oF9GkY1nM
aFYqyNxAgJB4KBXMWULIWBxFBZFzzhRIVQJct+nVio/qxqv2wqBftlmJtRzD
dPU2YTthKH5L3ugcgwgw4QExXI++N9Ve0uTs41DNlm46BPmsnIw5RVZ1msfh
Av3/LNsFVcZmUTw/twnNypE0MY2IfSC9mUVTVfXOwJCOepk7P+t0Am2komtC
XpRp4SsWKhPlAAAji1OVKcY9NV8AMomkGDNLKlb/dOZwfksioWSzsCVNAnVA
o3m8lYMjoekCisHSVqsgSdaLwhOFG0DUsuAlmtiFdIBoauqNSRgLJhgSpxgh
q2rcngaxJbjd9sY7qVc171Rl7WMJPoNOB1LeItRP0IxJvqMaI98fAA1faO/K
lX4nLiZcLJzBy1NDZ55ycvKPgFCpL6lPMkJJ6GesSknEI4unZ7EQPJoLJfiC
2+pXZfWGnCC6F8kzR5ksiMnGfGBIrVJzhJ02oU8SgkMW9Qe2kXdE1sZ6uFeB
9jWBFlSZzypkuaf7Bd8Hx6SzOK5n/EtHtvUimhvmUvNge7796W3v/oHomzPq
lbLqT9y99R/XhoiW3ZrTk1nhpNbz05VlCotN6kYpdKltzi7R4H53r+U/sdI4
2E2GZkYr75mcc+ReeR4D8M6ii89TR1H4DMT8+f7jYUncXKO42+CP+ZBss3ri
KNQvtoxDo1vkb2zf0KwV51ejES/5L220bUjxWsadLaUKZ1GfeZADvYWBkMIC
Opv2I5RADbXj4zqvYL2GETTu4auCcTsbfYgZ7rt9y+T7D8ZoxXJpMa9XO0gr
aqD4l4u3zmtFbYE4M6466IpRAhyEt+PY80wYObfzTfK5BQMhvBbXwLxxpMbs
cFRA3uVIf4on8KAMJX4EjuWBSeEhCBUJ+9uzzILpzDVbAUs0HZNu8rBCPIsO
bkUy8djlmiQ1ybT5oIR4hfHwdPb01EoGow1ZztYlpPmFrZvxrdQPT62Kt0nr
vXYC1coqWPuzR7NIU9N4Qy04exbhBLfZMbuIf9sb6zDp1VzGGcXOphFIIr+z
N1tEqYHC/TOB4lyjmDx+iSWndG8RGfBBt/uAHUVj6WefzOxwAmQAYdDCA1Qw
3T7SHqbZmoDZQKvZmpsMsxSuVp5nPywrxYFOjovWkTh4WUx0IMM0UEsyZCvd
PQI5DqUvjEnmp8JdHHWHexfAbHCF3E2VEnWKVhRQil5PjoHSMRj8xi23MYpL
Yr1dATy4VuN4xzBmN7iOMPwuTTlvH2YQe4dH5lWaH+d3YlcO/Zjy+Q3vdLCp
A8B6B9LKDVnxZlU9zwOPtf8AJhT1Aa83Zh//rzcKs6HAbbFZDZrBc85NWmju
vETTTf0CQQ+hPi9JpNZuvcFFXjXLuBMmRUHmjArKDq5mmrNiwsNucPTJkG53
EmfYjYewkwsL17Z5T+s/ucy0HBPuQWVfTnnBT4IAIz4/ubSI+NFdKP3Vng7j
aModatNXOdROuGpeG58DbB9vBLpYurb9/Q8I+uSAQiwdGJVAiYkvweBifiP8
5iimkhQuydXnjYPkO/wCHP/4NPgbl54kZ+nX4zmHoxft96m0vsUPw5XoZ1oM
gOEJ3D1f/e7/xdJiXnmEeniFjqxAO36Z26ri+1q+iob9GK5zaoueKsWAz7KK
nlN4Q+D+3d36EZzdo7RByc9oKKCcBMYLzTZF5wD14TeGbLAAqYilFwJkFhas
B2gZyWQw4XGhddS2Bhl7sreKGUnYAQL30v9VhpwH9oIAk+pkpgvFaGy1aObz
3b4qmpW9gYufv+lpqG20txMcai6Sm+t7nB7aIRUjd+eHiIt+N6EpN6/SyFx8
ZVTp3KQb2yV/vPS0x8pcbQxi+TAemY4zmI66Tdr0n6thZTUFkN8nezv5f+sE
/zxgWOP2GJSlcNhA0/OHGiCL7BGoo4bKLYcRjHR0HdXGh6V9BBxzgO8aV4aq
SNp76FqivVXDi3q/NJZyMW8xiB1ABEBhtBoVqzV8+XcnzEa2FneyhZx501tp
DEyJ6wsd7z4XAkZf+ohsUs/8cejfXrSvvBvCRNoSM0KYtoqbq7LYo9i4z6H7
T3oI34Q5gEIJLtRjxc+VtOJEIC/4ok8hixgrIjwnrBTuuLREV4ud8cTDvf0t
HmgYIoMBiGUiEdsKH6tbWmx6DkKzYSl/c7M2+sIhJe0Meh5yUGepsJ3p6xql
QAe0FhqqMbDKBrRi+2q2WQkyalvBwgMMEmawm6EbQUYKOzw/uq3kabHSxoVS
KVh6zc41+NEKqosmQCeIQ/8yFOUiGa2W/T59VopG/3XiNc1YcnRg1PTRpm27
blTuLgNUKTszIvnft1jnzHca1SoB6TZuuEPfXLGs+yXn8QrslbcZopJbN17O
iXkLUwX6+Og/xyqRRJwNKl03BFybPABsEjiyf8eVCOwJSuw+GJwqybm2djhp
N0624XRa7KkPL8BSQBLdBfxA5/vkl6AuNTIOIW7pGsYyASYu9Kwf0YlPO4Uo
DGvcqhVxWFYeRUDxsMzhQn1A0a5kqr4cUKks00Ltv2qcN6amWucUsp44Js42
fLGmHRsXZeWldZ+JO++99J6hQYfikwYCjRJGzU+kqN4yqidRBlwcVl1dcbJQ
WtdcWbZVyvSs9aPQh/HMAE/pBLl6WelGqNCmbSbnopyQGyNtVr9XvVuCVDhD
mmaDsCHtFb0Nntvx7A4KCm0enKtr8YBAL0eZChseu4zgPJrJmfnO8p1pSqNR
By9qK9UUHHBr55CST41Gs8FwGN3bRoVXXmNil/q3lfx2cAHBeZe3/JUqrZz+
JCUNkOmaR+4+M/vBIynf8x8DDEcGPlkgmAoid/qEVjS3BgapTPyy1l2JoAlO
8pASgCT5U3bOEAD9FLMemOrC5IP4cRjoBlJJPqqX0fJl7uICgqRzCi41napJ
7kW7z+DZtqGl5EvAFbxJahdwiSOL7knMg7XYcCVAH8uCjINFAY9/rlJcL90D
yHbd06IIkh9yj/HB6mmoomGCb9BvOKAyBK9njfktC5umQkV48ZETsvFpJJuJ
Vf8TzVvBJcM+0IWKNz8jtrkd3IF5jXVe2jJ75R4zKrG/W2K9EISQZBIngeUa
BObBVe/pJfVEeGCFe/c/n9Nos1Duhwmwh+pXgV1yIzxXmih4dPz+Nt2ubGeM
qD7mQaTh+xg+oOg+l7mE6p3UT331imvFZNhvrBw1r8VU6vQkUbnpYOhcyI33
QOUsc+Ckaes4fPiiO4HCW04fpY4+2L8j/I6CDm6mAqXsy5pamBsISaEZWwat
FmnjkK2sFQ3eFkTBcPHDX1Ngco87UN7DhfPDTRmHOGn2ttb18tAtLlvYIEx1
ULPlqyX+QM/o+yRjeIqERv7BayztVQYz1QRkIuZGWZTiQXI/tWA++BPIPWjl
2NPvT/FCPu4Hib7FgFxWetkW6m/1w7LqLedMmV/c1sSNyTWSmSXZT2mr/gCm
AANeVOvD3Wi/32HR8CUC4bDpuiYYu+jlXAFUrss/2P8BQCxd2cV++sy8u0IW
xId7LBpqbVWv/4I1e/IEk4L6stAYoaPGqYa3UU0cHmRDFobj0Oo1E/k5UPI6
hTzyw5bv16Igtt6TX42n7JPu5f5uJ9ucPmWybatTYH7MKY2g5xZ71U5dnfmm
JsIZnaXbh7KFwaDIfQeMBmJM6xbR9gfBX6ZLGBoZChd2kAGpKlW3R+1IwDQ9
/r6Da037sIXqbhZR5IDT05grKP8a0LEYQtGTXnFtxuDV3GPYKyiwijEDxwBP
igbpn72RFN0KL71skC3WjNPrdgpbYjbAwr4B+MCe/tQAvxYujX2An4xcznCM
sh3FXX45mPfSnbl0PoJ2qin/VpF4Yi2T+UJZspyPwnFD0kj1zrv9+IzjbnT4
+47Q9OGQItvM4OgiiDfo0x3bKxFuY5fpzdAX3tmtCx1isvde0GLb4cpXRL09
5DJvUQyq7pwZB91LS2Cv11zEZfAwIQgdJhIjSZYdrPCJ6ubTYSep7AuNEU7i
TTim/561MdE/+qOr52FKXETur0NXOiLK1Sz7Sv+twSBaP++/ah0SvpzHJry7
G8PzYzTaRVagIIERLCm1ikjyDIFNqanvfXFFMRkPUt6BHuydOQYeOBAYIkDj
isvJKl6K8z+G0EfqXZka86Qyr7A+mFXN5fbUG6+Qby9uOFdmctTtOLPV6x08
F3YabYRFMLdOdusske3dlV7oDMNw1jgBIQ1Vc6920NA0swS5rCapHAwKk5Cp
RVs+Gb7h+ltWgJhu5fwhtOWLZrS/ZWqiEsp90n7kEVY4AbGDfMm4s/WAN68A
jqz3h2LUcQDmwZUdAUXer+QdI6IMN0ebVG9Rzu3bl3QdXNg4xkmg8NtCHlQS
/7FMixkMPK5wE7Ey71gnQqhxGs3yLIDNr8P7xrcjiVMBFD8EUwSuNSfppPiE
Is/CYOEFym6cafbCzE840SX3uaaWypa9tl8MMVVbg6Oy6WSySdxXU4nAU3JU
Pq3qyZvoTpHkU0FDyRRCf1ZOUVpDSmxwfnQlEOiV9Dtg30GuxHke6hJ1TKir
sCCdZ5peqj1/WTzD/J1970t7VHQkAYoHBcrPbVp/di9Fn5HRiwXpCxeeZHka
Ate5Iuujv3Ac6YqGn+7fnlJ/za8IOSefmPuFbyPUzWeoQyxB2ooflVzA1u/I
9GsOALilsRrHz8nuCzqyl/4CMK+JgG2mIbfSE4V80yv7Ho0yMS/kmSpe0DGl
M/LQOqYBUJuZnfvs3+JgAHAjN1Xo8rIwcxPaRu9LPRORPpPT/Jy3v2SM1CJP
okmr+fob1+E4GojkGAyB5FVB/FFkMe3Co64FcwPey45fweWaE/x+r+qkZ3YD
LZbFpFPWHdsPsbmeHlW7d8ZS2DTgoRz+/y1fxrkJ/q/3OSDHmD33EkMBSCR+
pmcR1B6aKf/XJp+NopILE0x1AjZFWl/1I5L85kpHfwvvp1P1934BkSYNVG3l
zcvtPuhaGmJCRqOnymUaXIpU1Z65j1CMPkGrcKBcPEUPTDsQNlzRjcdq8f4w
EKVSCFFbrBix5Ww+VqhzdzZKeQjUQYbKr2GsZcafpI16AwAJuNX3bbW+Pixt
Ex7nYQOKkFNJIwoucM0JoGaHNwSjcKJ65KowBr564gdmljOuER8B1Moftmbu
vbrvYZec5MSGbZ8B6nrJaNKCocnEXbYrMosc3rs0saz8ECN+xP1W0jzOtode
MW0tPSdx1PL8oJkqP9DoT5WGc7aNJZfDaS/RMnJ0rR9W0qSPlhf9yFG3IM+R
IZtxB8sTBkem9+rwMGB6Zvkl4PTVcuVrSWurnPbVGjkXHVTRyu+1ICvxM/2t
80+eQ8CWZBAE7pRJ4KGHGMoIOYwxSVwmIKrXc7ghz3WBMesSFBuVaWUnYaOE
P6+ALbaDUQafE7AqmNz8XL5Er8PgJDCE7IPVBfHDsvRpv46bgtVnaTeAEPoA
1TqK1SA3g2S1DCfp5CwXw0I6C2HY+E3aMOcxmD0FHpT6mjl99xEoAJWqWQ9Q
eZrQdew19r9mGWQHRLkHqcR/Yrt2Yo0QrZKZRkICmAb/O44ja+KFFEYOTS7J
Uvbk8pMLSLdEKR8j9fDFgTrhpJFbfMbLf+jZRd6szFxdwp96AeQTOTjFTQr6
EDPQR4AXnsh1gZQLXP3oWaeNgxyMS0VtURBhU6Y3ykGtMh9zt4qn/LsASG+Q
59oiBtwenZ/ekB70vPEBDANW9iXucuiH+vJ84BkaTSia2qhnYRt/sLoVD7QM
8j9PvvRGpCZ7w0vy1rF8pdI8PqQcbCuVQyYTt8bXjVTCvjkKsIvso2vlkQct
8e7RiszFVPPdv8KFYqHH1tvfAxiiFtruEElxvrMmBd+7hkiYUp3EigqP1n1f
sut/daU3vL8gUynfuTy/S/PhgMq85bmF/m6frGUYmaaFtAstxVb2iN9JgBF5
rsWTa1AmIh5U/UMAskNVqBTCEPzU9pXAI0BliOTd9pg+gvcreao1BPdcQ0lp
Wx5DMU+ENcq1nkPXpkn9FpBmG+V2dw1bFnxMFDIuy7NZng08ytmbAk0aKSc5
VFVzsFapQNuL/PyzClQMl2Sc616ok3HOut3QSAv2NMewr4cuMj+ji5nnjdS0
rrp8LHLL/D29KWOGa9+FrYmgeGqoXbT8X8dG5B7pQz3syxkLEzkyOdom46qc
qe7EpJMsjEbtFW+CWmbEiHmUgW9nGSDWC2vJwFM+JJ5E2reQZFFbCTXqtCSQ
iuCU0TWfZL/4FdHEB8/bl8W0R1ZSIbxQq9W5jCTMW/GfuYjSrm0/fS8msFw/
T1q62hAY611t0w8wk18E4KrG+Rzjg/9BA7zJCOnP0vvGfIGHR64H5QD1e73f
TOSlhxGtMx5IeWPsTD8Ei/Xb2VOXudPeCzSsUi35JCA4IkamREW7NOnV5NUp
H3Zk+DZNZvp0KRwgrXRiiTpbhp5zNYm3NVFDU/WX8aq2fKX4YOKs9B1/h0FU
lLpxkirSMKJ/zfg9jrApXaTyVdBXLDETJatZklfVLFsSl/1v6hbjDV4hYOJG
NW9XDMSYW+U6HQEZxxGzkluAhruTSizXf6NEwQtFcdZMOEscckyEP2wFhfRM
c8lKSKQ+fYbJ2amqpSgge0D5GP9LdyK3xUtiobUbSy1wdRYz0FeIaq7iqz5G
pogiSXKWsKn4WWjBZjJTfYPtfbJyeL38b2F3YK57FNPILxeR/nAWXsiYKz63
7xry9w/T7BgGZ6uzq6PGERdNp3SGxZGO2mDzbvGBsdxR/5P+B7ycCt1kbSa5
3Jl7AtClCerdqS4FAcyEQVJsP1LYSM2hHEuwXXlFh5iQYko953ZgWT9Y7P8r
jBMMSaV7lH8XKfGQT01MXtsPyB638lpSK1x+GP6K7Rv6R3uzWSLg8VpGLQws
sK4QLxYTD4aTuUIwkcTuZrEkfanRbA+qyCwc+x/cwNr8ZwQcJP17p9Ip9DAw
LeycElvA01aokxdSlFJnkDY11vKtpHyixST75dXek/yAdy/Jkyff52IWqCS5
C5QupJ+Y/fPKvkKmTeETRuR0/uWivf30Y4bbcMCtyv0RGagzuSWdPZWAUCNR
v3/ZUlSTvzHWnq0WU0h2uHrG+Be3g8fV2zgk2pgElNSkjNEyLIyTuuPtquD2
FqR4tBrDfUKKyApcMDgadcR9EhkHF88lRSRbvsbb5lZTDbeb6suHKq6p8JeG
hYtgUejdGIn6bWxr4HgiCOdmKZqomivmfC4LeJDXKLpma1uvI4ZFMX8usY2W
KTEe4ej+n4PKKfE8mRsogUrVSbeXrEOXoAcn0iGZ6tpo9eHEMUhtJ4KdJz3u
qPN3DzprzezfOZlUan0ifa4mFU2aSbUYgH67VRbXwBxePAfnHjhlVrbZ1uZl
UpSII1BvGLGj2Z9RYdjLS3P+MyooMorcgnP7ihg9FCvQyCy7pCQnJvhLd705
g870pCmhAN7YJkDE8EobzF1dzi/SmgHpCySWTTXUw6ZBdBkQuHqnk6H+JqXN
3YZND7KDrSMtaWSADkKBUcI62j04Wc3pmWRnjAWFyDDhhbDpSa1sSuyD2c/h
bQZXoFJ6yNwx66YSvP2+rstIDQB7If8FsYAc6EyjE2AilQL4FVISpNDyBK2z
dOF0fHKl2R030qQBRXmaVCyMVNH1M95oa6S7bU9uBEXOkScnFxmG3V7FYzcX
B1w4OEDn/9hPH7YePcPogt+v80GIN7MR52AZNb/Aq0nGBPkufuoLJqwzyBRf
IbWzcKdC+T5IIZJX7obk6j8pUYb75BRZZPRhE0y8SXXQmzvBQGyaoyrogCN2
AatQGreXlUQ1C9ZMg0YAvECe0jR9TTFDcCTUAhJziZZARnlHBGHKvA9ke2zJ
XDd4h5Ah+WlpfL88OCfxv25RCwvrRyMPP7y8UOVbTgaLaNQi/DZLB28ybRTT
c212r65j5PdXdLVHMY2wgxssFNbYQ857cR76K5oKvtzCmE9tqCRiVHK66zYJ
qNW9guoL+gYgbAF+W9MloLvHYwthzDdAXZOOyZ9H3enOAlmDni9pTx+YFQ+A
m62dg5LWoidj1h/cfbWyTMFk8+GYwDYkVNCvAvyH5cQqcw7W272ReXPXTgmb
6AYvrL3eYAFCnQS+BoBSNrmkmP2ODYhTuownvO5C9oO+FRMf1/hNi52OsG1L
GSbGW0lraJ7+HwKbU6Xqjwycnz3imGwwWjWoADXjBIcnbAZSgWCnlyT8jZLw
8Nn+x1bShBsRd67sm72wZEoTJc1fhW/CO2R72GMQVhPRYjinADG2krEiUVy/
AeJpspDTZjF6PMcCm1hSIZu3Va0zQ3Imyvf/p2CBkZpyLu+L+DlrZ/QCA3Jy
Vd+DbxLI9JC57pwQwKJdOgnNeFbFZ7yGzvDDByhMj1H3QookncWTfysV6Imr
9VZ6D9UDyBwWF4G59XyW1ukcS2kWA9KBBztg65AG9wf4Qt1Asx22zx6eCOOe
9xMEqejk8fR2HxhFWGPJSxNDn4Kqfu0w2xhXWvDoz3zHoNUlZy6KJtr5qTqm
RiwSxUJGH9E3brJMheBw5pEZL7F+tsk37fXkv2jLGS99Vq01pl05cQAV2/EX
+CulbC+zNeLtm/OOPxAQPRimqCyjmNaPROP8ae+395mblnyoJpBFE2bDZoqE
33D7aDybxAj6sQ0WdQ091MSg+zwnSW5ofaa4BmPYK/1iQIC0bFUdUc1AeXZu
6toQFzjZqqnFKbxMD3XculC9DWxFJaQKHDPp39ZJE265PLuEZp0RRw77Bvmm
PUg3QJExFe7iX1LVas0u7r/iBOl2/FPNm1e2egCCyPKIDEu8e/Cem738wYVh
kMvkL5MyMiLWUtzvX1XmWkAxa6khQu+5YFPtKbbfGPMpI2UmJklwpEA2OYcn
t9u0qBm33Do1FATAJuIWTEDJe1sgqV4u28P2szBBTG04+VFsnQ2eyBOytjdo
WOShQfnLc2FYrcNMZN82UmpPg5G8vVIw9RiA+B6PPqKlyhoGFQsagO47HwVv
O9T50FIkNMQHGkPue1NNDGCTiNB20vwZXpWAKnWDwyy8pV6DLTpXgQKNhL9C
udaGGobJk1MD1x5Xg6cUeqeaV0xFfpcCeRbaChCN0y4wO0jFY7r4GPrJRdf5
Ovr9++i0J7t6TyKe00r6EmxBT+fJmlcemECieEOugMH376I9iVzJXZJTNPzQ
kLoylmi8vjzRV9owAmXsRrxMZo6rNurpGbFi8zTz7VH7FUt93dKm/2JYzuJm
6HLH8gvp8oSTw0djZaxHCX5BoXvElJtE/4LvhACOUMinFKjD1Ll9i3MaPMFT
p9GH8ZvImBJo78Hc797Pz8BU2OAxgnReLQIQVa3Xuy5A5jlwUaugpL2iISJb
1CU73oCgtppG5lhPq8lbGXMQdpaFitGN0sadHiJUwtsgfB3lEP6zHgYPdHWK
GFoxda6g24nOyinMYWkgRVRWEZuDyhy2StMu3zjaePyfi6h/WTi3ewiRhc1v
GNWDgRvlq4jwe2m6fhW9XEYjJjMt/9ufQ9HPD8grbsBF7PZ2PHkEcz7oEPn/
FUSSay58yYyEMS7yenpMgakclm/NM9EAR2kRknEA5LV7SczglRrETHyHQgfA
v4pDPPMxTPZwYyS6nbcptlR+hcULdIcvFEY2g/0vyhlGLKLeI5w2ojnT3h8S
b2UCsGe6lS2gC14yjlUJSw9HE6VgNkxCuxeS5A6cUyvtUnS+0e7cviPZga7I
+DyfbYimd7GbGofwXa4JBR6LST6BKh9sYUYjF9xpCpWphi9yOxKKyGRfmU7i
6wPh8jrlPvlSCpwl5Scdw/nZGMqIvx2Ihov/2ZpI0SZbvlwtFaz6zRz38zG0
lP1zAetQqObt/NqEZVWt6b2RaW/cgHp9WiSmGAt1pQvzsdno229/G2ZNdCs2
0X+AeFU1DZ2WKh410pE/5CYkGzGhV8JqoAA4uKdAb8uJCUsEI5Kkthc/ilTB
AZfnI1Qn9iJvXi+ztpYqzIRcAVkWTjDZDxdbwK32fy4mDR/5+kM6DqYcF1DU
d8eaitQ1q6b+HRnTaMVewVVOLRE3lm+T/sjkxHUdGgZIFDhcqmx3YxGPfWtR
Ity98fl7P5MtDm8s6sNJynEoCCJ5cfSaO2rJKtL30kfRqvjYI41AP87E26fK
Rk3YIT3JbjUo+EzSHqJghCvfe9l7ZkJkha5NaSIOH+ygBvmRTl4H+3YA0Z0u
5Rk/ZnRUwzg4Mhr2Ivf+lBbAuDsZUujNO+OLREfUlWjiqADfk0epteM73zrX
TdZwX3XlAgSmxcydsk22Al+2Xld6jrcdy5yqj2cUW775b1AeK6E2DE5OALVQ
T4sjVazPAgUJOc3WuOIvkxwTBuZD1krbZF+ISAmo8YncTbQ8w9SHmaVlr7kb
TnqGhNMnvwU7itFkIlv3d/qziXxISxSsKSInos2LGWuWbV5jrPjSpwMas94T
ZJVdXGeFYYcRbHemGCr6zE+yPpoyappt5NK+ri0BYnLJHnKd78ShtO1oUi+K
Gy0RtOFMxCqsUn8sdCNNHtVoB1wdWFFoIucV7DZ+K5ACXq4MztXaxPWw2O1H
Kv7mdKCcHmsLu/1gRRWFOk54nk0jnlkqRWa3awJlcA9sGHtWHvEAYXHTsttr
6SZ1hspayumyJAO98HnHfbSC05bG1GCCrcbBX+//AT6kr+Vtat3ls2Q2ZOWa
AtT/ODBA8vTkapx2C6LS0uSHAnTwLTPQ9MkBoVFwSTxWNlaplCOVEojTuCaS
IRB5cIhq/JSxnkeHXXssOSFWx4fAs55romHIVDk6LDdKoNRmBcbXj+SbpTva
n2VJbOkk4IOGFaMpXWwKdh1NZ78L+LMAWrq5ebEK/TNX2hedm4l+7K3KUHdt
/RG5qSwfyc7n62P6+1Yz7+lGjeCqIdGUUjPzjwreH7GuP9HqfRnwNAG26nWD
PqJJuMYou8UeCNL8Al6Rxs5If1V3RgHKGkZXs+tdyO7x98EwHtLhkIVmN9se
2aFx/1sp0E+KWhZb35fsEgbTpoPo8xXnwCf+8PD+3rGRzpCIhNDvr9Nhj48n
bjtKeBZKvBTkxlvpixTp44LjdaZXgXoEuE2texzgNwQUDxXEz71ufG5QFtUh
qxs1h1cbmEjik+6kFq1kyrQeuzUmsiU7v44sRnHMWcxjQW1wer6KSwUZlUY3
mKrI+6N0BUhZOPbNnNq1ARdMNXBGYb7UhnJMpaYp/K6gjWuSrZulWI7uEwmL
bCCLhLFQwhxSx5wqCmhDNW01NnYvqY4LJv8g8xChAtLEfvrOk37suJVtkDNL
3QeEjS77+6IKRJqEehMC5VnYwb4IY7QK+0+YDM8Eys5bW/ufFqDFp/If4lWO
xvEbp+c4gckl2ki1EzXkMQyMj38r98YyvjRie9SLInfUMnYfh05tXJCfuFjT
0dx8xwDHLZvuNPuyMi1k0O0zhyCAwl3za4PM7noy1fLKFO25Q4kajj7+8xrJ
tiTb1TD+75rE+ORuz5ymy9zvVv9pzb3q3ckLNss8ulSqs+IkihESiOUuVp0e
Ylq6AJ1B5JaGromicmtm93a6DuBO5wqi8QXolF+1dOqwEnrJlWsKsbOHywG/
tnYpBqurxCdcZ0M6ARcA03AAc8ptzXkVbwqruHAR7CkdehjXLa/oEhxi/sh/
/ecEaWeuyLk/dby34+Rhsicd1QKyQm+23nkDOZtz5Dts2uJ6D/+nZoNmWzvl
02bIIslkeVlnucStojNFdn+5OQeHxRj55bAlrQhJ0GSzsWVB5TaPgGmaWdxG
VC958G0nqkEEZE/EScnuT3XaYx8gI6jKSHJfHq5TF7cM/tMoNVlqUa/nr91V
/GLbJU1rmEInWe2tIJW5QAQvuBg4L+Hro6AvYbV3gqpyPH15tpFiPB9Yfpw+
s/dhwfBLobGr29P6oCYCHNlDHSky8odTzLODDxLbhXFVm4sYNDRVgNlMHob0
XIkqA0xE0QNwRaQt2vIydP+frRApHywGro2+iNDs4LpMqPj1dkLOpvZM514G
mL3tduDzfQ5MzMtauSNIcpvoRrzrsIeIF7sRoAGkVvV2gbNbNb8iuKq+fYfa
UEjGmLLMUvQ9OZY48h2y7+hVOmU01WfPRbv0RxX61kuaajUOo6W7X6Vf75/V
aTMcUETzj35QZnkMoDc1AFqPMAu8Ur+31CGbfSvaj6XCli3x1N4q7UN/oQZJ
kZrCgfKb5SsSVgUNEGSqLePAYBhQSmE2AgdG4jx02OuLhIlQHRXZY3IsF5ZL
sTbhvAlGlQHvIoPI69mo2HLoEyx4Iy+BUyrnMom+KhGqmsFHQ2mVOfkhR3EL
B+aSRLqA95fs1o8SQXWNmWZzgO1QlUvXB/NoLkUMKsPrdlVDu3fc8zXb+IqM
kJCwieM+5EbT9ceIosVcKmhAicV5CXoEaOYAeHwANFLmBReQ6MPMtb/Jc9o7
B3Xk5zLjmUVOsFwl7fqBDHXeeb8etfK/kVDSPIjbPyBU5ssHPSahnKHiftaX
Shsxej2PzSv5fkFLRYs3jfJ7AhPAVVmaETg7iSekFqSppj8/o953lMMnxzPc
vUeLoQgFg05MSPeNRnXm2vxdjGxNIoSl7BHbVRZgfvs74+DrldRkS3CcEonP
20gOhoRdra4kjeQ9dG0YrPc4lwLLpwXI09Cg5IxCAqfW/xYATwKXrgF6bSD7
ySTmo/eeCYoeFo9rMlpSbwjh/QAmtbuS/QYwlXgZSfMchDxZXCMpt31FYFML
q9HPNx1eggqEe4KyPVrLqH0gjwCEgUkih9I54UQTymbjnp024X/0kt4A4jDV
03YgWoONP9bQz2IVHwcH7XVeA/ODz4InFzjzG7kceE2R2nEcghIDhPIYZaxi
Vu1ioFxcc7lJIMOQA+6Qhy9W6it8HvQqfetbX0UE6u+WCOCXUO9Z90tfqRpe
pu8uL0/kEvxeTsO0JoHMWe/F1hO4CJi+m1r9YdtP1JEXT+hzCcXtUA99ntD7
Gw26swbKsoqP9HQ5kg4vanLovuSGY/ErH3CgRd5qi0qy47QeWl0kp3PEC9No
X8mFAKsfgJ/HPuhVVHkMb7Whel0kbQCy2B4M3HyeyYpW6bXH4VndNGP26xzM
pcVxV9d+bfKh29QqmT9uF35wS/kkXnX46UN7ErkWNiwLh/0Y7aQU00Gsqzvq
7FkP+Du8ILc6u55//9ID6OCqQgtLIuRUKvT4PGc+n6sb02FgQ87SIpigzXHF
Z2BPEM4mU2r5skEvSSGu18jffZwaIfTSUw4g+Nryz/FI1tkzEKGVK/o1JbMV
lhoOTEBYKdC9aAo20QPJdip1qoeg+aFRGe0G1QxoTWRAMSKcAdPfobXTYQWG
xk4dgixgZKHuyHAqqDo/y4/9qjX+FXZ32r3mrLdtsSPn+OESkDGAf36AxZiu
PHmOpzRfJTsrjA3BG8pO5YXQAdc5ZcjKftMcIa5upW1+auEi+tnSMqxjXCHb
aIFDzGw+ji/6rhjpAQiL4Dbu/jh79JrqRArWgGorfxMQxlAad9gDt6eH/kJ1
+hJk/ZRAnCs745ut8Lyv+xTTbdYQuB7f4rLQyeC0DmAVHztJV5tAeOKTxRr7
BNqEhVw9Lh4eI+37YNonPhAnSD+Nkd+auY3t5vxIB7fUJBqcp9RaysMblObO
eBmP+aohOTsElDD+Tkmc+teML+1hoNfloHj1jWnSCtdn0PO6KgQWRNKPjpge
Ly0rrU1UWc3xuRlySTi0n51tIr+7A4dzD4RwnkcUoFEovUwO9Swuq8le9ZEV
1UAnbNr/ccNfKBlmVI1Q1q0M7+Dl2H990xtdKQV3sDm4AcK5p0ZGJ36TFt19
3lM29bTc1rARwxT7wsrs52ws4oyGSmYrq0tf0aWpeNlu1wbgfV9QDTINNH7C
9tHE12jjZft6EC7Zh7TqtIpn1q9Jz6sVWifWs0DAPus3GEpfAovMByLXEXJy
k+3y1cz/G7IJSMLZQ8n2Eg3rmsjsnPQbPB55DK1WBO8tZ7LsUr4/79a4XdfV
9rANESXGw+eBBRPf0JitFeaGuWC17Zaef2KbR4wUkgWrqW+Dt0b/jn92fVMQ
PEI2DTTRELs5fXunJ1SOfnaFT4mS0QySwn9jvru26K2RArczoQODf5x24j+K
rg7Ro01QP+tCXM2rfQUd83z2ad0Of0lbjqh2EzgpVhu9xqDY6m1RZeUQfGKA
s0zIaJa7PS3oOXKmro59rLO/uTSXnG9Eslecu34R9uS94yOTL+nLj4XhjoWM
sXLC0gTamBPaGmHuIJzajUW8e7bhQzX6NNa1MXnWr5el9F9J+w95BPMHN4wF
Q5IbOhZnbVm5+IVFsu3D/qkX5b1YhODEH/6MNocl2RZMb1HDNxNwb6lHTbN6
+hdY/aDCZ0fX43A3dPw0zP5+e3NDFzclOw9HYrzJD5abktj0tnxd/VE5KUI8
YVXtpShm8REJUqxg3y7oOn3YccpBwhwZ+ELrLtzHJATjjJlV6e/sf/KEpiAD
wwPvcFFBMXXYaXgCNFDYuh+jnX7xpTIHMuRsFhCHv2ip1hs0ylfSU/Cu5RGH
vNHTD5mrniJBvn99NnqBlZePVeUqyJBPGuu0GFZAIbfo4bIKBZ5+mXqnGf2W
n4Sb39Gy4NDWi/r1NLtPo8knsP3E8PUuNj4yZ4twiTTQ9RucOd/Ye9fBI3DN
t9sv3XsAWIsRMZjZ821Kr3meVgBM2rt0/j8pOWlf4H6ASGAymLs1HIKxpFz/
WFdqGer67RzmAIWx1xQOw/GWV3HBgEIyiLUTgEOAr8sjzFQ4tcL0kYbZTl5T
79N/5hZ20w4daFhScu4Ke74BqqveCTgJU4w+08/75aYQ7gg+FDC9ZLuvZcMO
BcJBWKQCk/trCE9+tOsvyPfskCCB5tgPoVgouYDR2wRqZxDcJrmI9Ugme/Q1
a9oYSejv1m5HrikRYTHE1z84ujLqDUJ0LBS9/KgCnlmUBAMoxufSUCPwMbgO
PpChc3ZEqyzju0E/T6NxBxIjA08NuIXyIFjCXrhj9D0X3OlwwXJFuOUsDd5e
VNdZo8Av/WSOezRTngFsRj76zDhlffIRT4oAYYRXQTc9fKSW5jJLXykOKD7Z
3ar/6r8Gsw0hEWvFQvTEy/w4WJ8skSAj7pFkcm6jjktdjWDcmjpn66b43UC3
kU0hnFnS8txyT4hGTrbAWQO/TRl4H/WfUbKeXn63ewQs/6t1XJy0nwEnuRnw
FNU80RsK/sxW6mneC8Rp6qkM+lRhl5o6Y6kcgmjDWyPNP2L/Hi2eglJDS8SO
bAzwoMRfsZj325J9tIBe0z3dz7wMMkPHtjoHH4kxxaskSa4cmb4k4TttrXNo
zG+cVsBJmWUkE/4CQj3Wha7lw5Xql7fbFiXAON7sXfW7Y0yMZ5UJlsiVDcaG
FG+jkJsWBSktIOWwqqZr8MUyRhiu8K3lsY3nwx7FdkPiz0cf4hsy+ogT3E74
epuAZOILV0LtHDe6FhCDu9g6ALDJCUQj+msxU9+6CdOTWySvSKxkgkbD5G89
DuenON3n16ZWMXn2TDlA8B0I6y1ANwpHqr6spUSpJdpgROVDE6z7dlI8RlzU
vIc4BDulcoN+/b1RfrQ+F/l8IgyaRrw3rzRLsR6DBhve/XmB7bvfOj+W2wTm
7d8z+97gNHxAcaK4iWLC90NWZytUGLkJqbNqnI9OlXn9ocGupCoOvsfr5XW+
6HNTuI8R6eiM/3Y/zM1tggrMZCZWnWaIBkNSdmePhzEEkeQG1G6tvou7vbb1
DxgQdgw2I12b0/mAlfIlxNXYQJr6/v+zyzrvYPnGFgmpDJiuvxPaHsudlRde
O5LlKUBr5H0MZvHFUGDWm1s/waDbBVGknGomYauBKLl23nRg4ANpTtbWQ2Bw
KVX2imtx7duprB1Dw0s0hDjrVc/hD6CS8bMXFB/7IsiRuNa4s1qliBCJdDBB
4+3eDG7/KItqWZYwiBunCByjAA4nhMV1phtP1cAwLGoztiexnp+bTEZm8Y0T
uEUhlFbCW9bU1nqe6nA00eTXw9bPF+aKPPMQjZaZ2fnqri1WHLUy5rQ4VNSE
UoQOWNbsT4QprN+rJNy5M1imiRBdCy9RMjNqtQ6vWrIgcKCdN51NSRvyuffY
PfGa/QTgGgSYXsaF9U+WDTpy7PiXUlqQuo9qYh/7VfUdlIvad7eJxADcv933
n1yHSI9XgJ1G9yQ9Yv/v5RoCfceJ7SM8Ff2Vu3SODk6s4ZI3y+KAz2PF+fnV
6pr+Kufw7v7OHiNOVg3VszUgMmtQajR7hKLnYF2Pi4p2Y9GzCEY0WXqkjZct
vhh0t+jeqJkRhi3lpau/jpCaY74nIBuPkhvjrPPAByHbFdre1+YM1rH69Gb1
fnSe5K+ki6bX4SvgHUpEMmYoFJaSmh0CJzYMgYM6htvjsUVJylTEt/rvqqA5
bnEZe9X5b621PDDXmW0lh31gQlAsoBa4JGRbFr6TayzuzrdmkXmJthd7Kceg
lE+jLdbQx5eV3uphho/0WaEiLUIKMoECJbXgQ3wyqmublqJWTLA8vmjLxXoI
tnBtTUcMgtskunkza3yUPqICSO46cA3WqsHGa8XbyMCga3eMhPyVMnekYC63
ij4WTsb2w8WH5Xry+VaRzzLnkFDoxoGcH/wOIf9FnXr8CjLohYVAqV+t2LN/
J4BJnI1h/2eG9vKcvz4IthVbC3hxVSel65MYybS+IHLJqIHbX361ti7MOTHj
tzJIpuasZhgK1Dc8EPk2yMljTVuVayH/bvqyHDsU3O9DM2REk3BuskfFbc3i
vlJoAJQiuIs190MD2e2gcj9/Lc3zH+IwsMuGnlcezzIT4zfgrWXJFDy3MRQ7
aQPOO+ddHP5kfXdrZmXdOH3+pqmPrS+nwC3RoE1L4+TuZ5Rbi/Np8ulKJyP0
2k1aqOt7ICFiVFS5iyyEDvwooX0qLNuMskD1XHwzmtM5LSD1ivhDTH0g4ZAz
2zXdf5FtA6I4cdaGsvaeQXBRhU8Fh2yqV/dYfHqmElCHAFlWC8ON1DmQJ/ZD
Nq9RSJrQazMKmfTJ2Z8JTDwLhsRtZxRyZYWjF/IDXbv7vVUzg2L7nWgioybp
9qGggrqoXSUSCFxARw4R09whI1RLBIHXUaq4YFA1IIX/Ml9WTk+ysPGW4LoO
rKuze9WW6svzO4lEHd3h/42JD5xc4k8/5G/jWlKp74O7C4IpJam3raIlnw0E
NEFL8Khw6myQEpC5Fv8mZoBg5vcFXa3eTemrQXJiGA106ETLpSps9xI846vu
aq5liPArUJ5Ld3RK5+chkv0UgMPX4o/1F+FCMFs+jk9dEUgZBokX4QJkU5oh
SFg6SxVqTs763gCVKtrIak0nKzoc2Ls0YosN8QIee5hJs19Zkd/ezN0UJaCF
i+0hOjFmCEm9oiqwk/PlAcPqmUjAZf/0jwMqEEnSZfxI0Ri1QI/F/raHqj67
WMXs5nbl4+Y4pMl/kDXOwLlHD07M6H2kpR3Ave03Qxej+wkuMY+rs0QkAn7i
c88hQK7QjfCjZNEY2Rfz+YttLMOFnAFk6jNwRe9xdnIINft95IQSZGfLwnO2
vSypfENh8cTy0eWx981Q8qL9c+1lOkCTk138Un/yVW1hpDLkLduJ3fQSw/wZ
hGferUeAzSnh83yV8Yp1WkBN3r4IH3cI4AiQ7qom+CeYvOeFY0/UU0YM4G0H
a5nb9+Vv/yRjfIEtFYn2tlVt3bgqlFD4rNzDTDHSrxfERFPNQ8NWlRktR7A/
5FMq3Q/t4CJfUt88ACUuM5O8kxAA2Ow0NUGaWddwUI7UDw4bKL+kb5kqQ5Xh
Mc1wgNsnmikYXZqLbgk7WnmOyGWo4VPR/cxEo2Ic14xmqkiQIUHNMa8QPYg7
nA0dSuQvq8hxA3sUZjJqN9aNpNZ0LOcEOK6LX5Gz6TIEodIjeXbH8BSB/GKe
d9g6Krhj1N4PRxU+jNKqSA/Xw0H+hyzjRHpjWAxwCRL2gdKfihVFAJzjVjL2
tS0tZIUn7/H9DfRQSluzPrrm+byKWk/HmZgfqkakY2VyCyHY7JuUTN9hCZ7W
0VFgPU9+ZDhz5LfviPDKq4cAd/nlv9xuiZjAYJGcsnOLtamgOl+jjhOFQZCd
3q6xLBJ+dj9X0fZhM+AQvN53OkQinxORqeZptV9F4hEODq8CQcJBuKvUlY7J
77TahIcv0B5O4aUSq9rH5tBUPaE+rtgjXBPrUNujkLWAxniym8X833+4XFNy
1EcwYjKF9imma/8UGlSEke0sSLQeeXh1SjELnOUohoYy2IiYMBBoBI1DGZJZ
7Cpuif2D783JLsY2B8mlJKF2rD8Z1uMrADVOl2S7NdO8zp43bxI++4NutSsM
WpDyTMLW1Uc11CgEkflJmIBPRXKZ6B+SqqOsEGhG8asOS4r4bTspI9xHviRv
2TPS+mrPPgwbNI8XpV4yQ5Q3gPG0O5nMbrd+XpnnvgZa7A9yBjnKe4hQq+WC
UsLm56oDtwT90vLZN+W9iPHF6+37IUcEB3o416BCzYUpaiMjCjJ7jooQv0w0
1hsUVmJ3iba3CUcmI77udw/yQ0+NuIrRUDCd/b02RPIp4F4JC3b+oK2b4bzn
HqueoAtzaQk9bj7e6zvxDfPO66HijytYJobhfO0D5Jyfl4Ku8RnSRdheaRJm
VVDgIdhRUC0Tx7K5L0MSMOr9oSSDoYTUAD2/13htgk0jA6K+TVIR9ALwXote
LLHUSMPuCKYtDUfQorcRorUHTcTGEO1D4iZwumwZySRd3jKGdYr4TdqnL7rw
r+Xnz2s3a2PlCgZDFl1hMJMlzSHW7XpCl4ufOuCgJ1vsmm12QrqsBealC+oX
ojf9ZOX4LC+kzKRuy5VZLXTypgMzMod7od3kjVTxoRSIyejGgmz2/aVgyhWI
mZvixjB3s+euEyeR7pNP4ktIcgcM0lg7O9VLaEU+9QJYA8tbts50gyXwbj3D
X5KRMr08myVwzx99mMCC+rvPP5//AxOutCLzTVDDrV8Xl2OYFFHDwAZ4rBWi
58RmuxRA3uC0IMDjbivDiH+rdttJgZelGes36evbP6TTK/PzHKVL2oD67BfJ
M7jsdcQcJyOpiGzH8EA+txyRKsasKgbd0FL65h2jbMSZ1PoH9Oh7VJV+24Ts
EijmMYkLH9AZw2KYxXr+1LnGn3b/JhQ0w5W47Yb/r7CaVX6UgA/DEhQLD/Rw
LPgoOJbzepxL8jJMKrMZVSSkiSJ2GBBISPGnNnxG9RoGMKByWvcyQpm8tc81
xG+x3lB02eMGt1VEZtAc36TD1Ky9VXcDm1bRIFZ3UXaahD0+6HN9Sj6uyTrR
8VP+SIuhyYPIOecHofbQqM+skxSoRIKBx6yTQ96ErZ3oZmWyz1VbWYuNJXEf
mDbO5jxWVtQWL0iONFhCBMNFR03hU0sGV8xKFvEa0dGSP57IkrbCIYjXoPK+
YfoSx+wjBEzLWb9ju+R7xcEHKwWBjjMr5q855vPcC0hOIb9b0zaSXYloIMCc
4lhHuymCLsczYFtCL9FrCpzzX1nOrORyL3JH4IjIJPY20o5l54W/d/81ql+V
d/Mk3FPDjpE/1nauFnB7oBeMQBjibnnP/wH+2gZK8080Yx8D5ugjUofbO8Ht
NmKEBs/Ycw1MWYMaHXFaOhkbw1iAZDJ/92ZCRYLO8u6wK7vRbtCFC94pSzSW
vtszCuGNFxlPpsx01twPoC2lih/YPeoEXquqCeh1R8WEYJEP/3TjgudgxwZV
NM3FulZ100Z0fA5A/7hA0ls1+Qx3nXrRV1IPMLG4dfXdibkh5zpdzl09N68c
ft56dHC+LT/j6O6x3AMtbdEG0lQtoU+phzQlbzq50k3liP3QQHb2xOHK008W
xhQ/mQ9rgw0h2aEXy/mQSz76bvpe+oCN5/AU6VuIvgtrFcHisHB0yN+14P2E
CrFAoZMr9aeKiM82mrO4thDvvx1b/meyunQdQfo93ggGXdS49l2JM9VZ8P4l
pbaIQaeOYS2Az8HS7pXPUt6oUVEm0T/fjYltMMZXIarDNpNqIszW6/HYMVjF
AgsdfXdApw+FIZn1qG/myxg5nQ4Hiv/Dyu7G4uLvoV1aQRWyxFvl+QyswMz4
DjdyFevHx4TCvqoMhqwhlIO187EhraNlBva5hPfc2jnot3H8S1pFfCFRe5Yl
3cM8kJkYqahrwaulJRhRjhftq7xjDPQtCKeZKRstj3vKS/6CbJSHAaP2QBP6
8ZdKEJ+G3//CmO1OjEfJQ+LLgOWz+lgUNMX11hLbJkS+eIQE2IlJ+P8R27R7
GSYnp24zIb337Aiq9QrICHigDFbcOvhIEQqJsLYS3DyS3cQxk6lGLLapxOWM
zhKh7uf9KOLjF1g7q2mKtwpJ69qCfO42pU50SFipJAkQUqKrCT688yAX6RoQ
jfgabtJki1E4kS457L/NDIo6pxzEokS6DryvHYzGULF6wu+ajjWeO4GgvjKm
IeIR+OfZVpyYLpjsfJw+ZzNQ8VY79qNlXsilS5K7XGcgTE6Pu0eJKzlEUuRb
U3bTS3l/3u1zdHaa3O8EMfusOi1oWcsZMXNiY1DLDDDH9n0XOXNhU1i5glAN
V6oeGbuL7ZVgkDVbaskIxMpnvRPYC7kT7E2NCtCinvq52pveFpOujBgFJhIS
w+ZNkJ7mRK+0mc+4OSyAJJGxxtvqu5xot+lenby2jNa/JNhaHAMmQm5NBLw9
VMn/bXmSA3rNezrfoInEnmjPrLJ/+OSt9AbnRKRsiKycEqw9PIJUJiy2OFR6
gXynindBinvWravMTd4YG3CT6FaPOtwbgJtXLwQFMAv9tDKIQuE5hNaY/LWY
qPdfbENUAbWUAjBFp6URaf3219xLGwd093UI0U6n/J8whuOQL+DwBHlf8fIG
6RQx1iHJukbqkRbDQSWch3bm1rogdcSwjV/Njlu1aUkah1XgTKa1iORg9GEz
zaOADCIpi0M+WMXLwxQtlY6ee/16AatqdzXmjT1Ij194CwujSHp8LwPDoByT
VMSsg8EwlQ7JLrmcm/f6bO9bGXFrwVfBOwnphBnuS9i5b+8DzdH13Bq1gzED
o7Y6gu0/+QjWI72DSCuGUSpSo2vEVZ1bc9o5eNp5+rooZAi9EONqCcJO5/TW
ek0hCFZnTcyBMVsHIZjhlXzdgHPTsj9nr993JzL1Z2DpVxCaTGZ0X52shEeD
dcvbX+G2SWeWR39e1DrNuTyRshS+Viz6LAVMZcHYqw+92jwklxKAqwCXN+eZ
kMLcuQ6TBa81hdu0+KlJkTbNqbfj2RvJuhm+BXVYqunb7wfR3uhRVKBHNOOy
pOpmIsm7XJPoxmPs4KETAvNkEYDtNJGsujKMtI0AZAAOMjSRCGEbcn0+SKux
OcsQt4w92JLE5D+PVDQcXV+9AZkcdwcQdybWt6N+nrcu1dmOJO6LZIpJW/dg
baqKV/DI/AmBE93+fDCh2RCsXKanUD+sqpjS5hOcrgFNyWCq2DkH6Orlv/On
k1xsFM0fOLBqUpz3WlQTRbc0l0J/XQqHKWCRe4aWE24s4X9uo2DGLkXxjsHf
KOIwcsmGchf5oTwm174llfFYp/aVAJ55i1Zq8c9a9QowMTqUx6q16fDVFwL0
CBfq3WuM+cfl92+1tOUlkSngZtUY60UK2+V2sQWNeLn0+/sksQfnKK2T4XcI
t9avKGWjyleXoDqdAkPDVLoE3/kooZ4CsvUbnknqY8MI5XfZPJKCW6TCAanX
wOyo6UIgYQBhCDlFqKH4GBXrHY8W31ITRxtAtYHEnk4QandHXFjNq7PQEiOQ
vRNQI9FpmxMKREBny3nW0giDTY23ccVXnIMql80/DE47ZyZSG/q0D2HzPku7
XhqqS1DaoTSz5Xo2VDjIwrOCIrjKFrsRGbeq87R041lzwvP4Ly4Zyof5TYOi
iN8sCUXbM+veHLDrrWopoQExSe2UYiHQC6/IS8QNwDtbfAeFQ0JvHytzyl4p
9O1TOwY3TyKN7XesEIdgU3Wh3UtDZ5v9EuLY0iyD85RtsgE+M6TX28NdhiVL
woCfcc4MieAd9qIVr4Z6VulGZfuOaK9tZr9eLeuzp1vvQAap0vwgZgk0JPCZ
g8UzRlYOb7WBQl62KL7b9+5MDD/+PpqNSqhEKdqg0o65GFrsyOhd2nan0maG
YAFagY7TWiR2VMNspIaFhAum6Jzhdm/CXu0v2SX8Ui69ccpID4EnZVehESfd
+A4j1EIYvB9F94mqe8Du+SP3Xxm4fxw6An5nJttew2/j66KGcrluzGjRFpT/
+k5TNwUMHd5bgcsJwWfLUykLq2fv/Is0hLsoPxaQAsffAZ8Jig5mjqi94FfO
rPx9bY+7FkEUVQX+M7DjBWGYUgDwJjxoOl0mdtQmtOFDqszS2kNZrqQKXIuF
3gUQEQzWyPbNcV5E4+lFYE9FaRl+65iSugJ60FVbHoZfse3fMolv3BykEsv+
pwYllerCzM5C2Y28+sdwwEs3qvjVE1r292XF6k6bIIcXSs8o7xIg//eBVuq9
yqgt7mxQaAMh5tUq4djI47uNR/b/BxjxF96jadGYi2Jza9P+1c+ioDWb2M3i
P1TNBWZkMYDY+6GsQGM1VNrHhG/eCHpUFZDeDjQwhaINBbkspcs1+u28eBys
bVwnljcW/VV+eOCniZZRCtC4kXeyfwJVZtrKdhjTmhJ28m77KcSxxImTm1pG
FI5g7vdLHeb6ytfjFPMZkUsyW8wnIw+kDNH2tXqB52QBO3FX+nD5tHQ8yug+
7M2mj+DIropH44vmp31JHrrB0Xgp99mKIz8uahDh7562wB/+8PDEJRyQrjyo
TGET4t87nQF3WngmuV6vg4a2yuWRIpANXMHe+0ujF2B4Y9yCsrmZNF9gT/v7
p4/vcHBIR52xB+h9WFml6Cnzji3Dhmwr3Oyi547+e7lt24ONYubiLFzZ7NJt
wPn8vZMuKaRi3F1ZdsbwiZIamlv7MtckIvq6LyDrjUAlc1aCkr5sDON91GNk
r1mJ3kBNUF17i5jnqYauXla68Qxgl4ExeVSysApPu5COYF4tSUYW9E1D7UkF
2k3xBSNQ0IlGxrGMLwwpctU4ticp9Smkn/1+DwAEbd9ZW83wPaJi2irplidj
hjSRxNSsUySmebKLxTVEUdeQ+hftn1Us7TCEwhKte21qx9TMlkBikPMngdma
m5o5UJKtjEMuSCEpjq1kUyhHh+zRrRD+iwA0h0QqMH2nmgkvD2NMzwmnysf3
7NH2O7AMgKlJFYbs4jpvQAwRDaNJ/buPHgYJxsxyP79nHGaQJXqoIDnxbz83
jlfLxANjuh1yZcS4/MP6smEvE2qSwJ1YfFVDwtGCCpWOHNKs3KJRQ0PF/7Gr
CEJNyFw2DrRVVccQUp+hHVqIsZcLiqRzAJHjSmTsNT9c1vrqZAwnzITKFs5M
jCFmlwOTaEKoNYGF6LYpRDXHdfpMirYRBqMj1oSXYFCLbKLZ4iheH2D5C3OS
3TaI5/tZo6RszbcCaBrFhkCq+KK7htj8yWhrrbmu/0D1YPlF7HuyN8firmqF
Rh2re8e/O70Ce8Ggrpd6oJG1ilCcVfreBY4ewJ1zCe0oBNaqBBF4kPmQNRea
OeAwgC6ggVFnd8Fpt71ir9u13iFavqSOZQNiXL0qvxS0M+/aqyGucqt/G8UP
3g+aCE+kk8UHyuja7+2ACa1ExG5xspJTLgGcKO22OW17ssvF3iJCixoHFeCz
rw/cMwXkOR06puH2WYyIN5L4pVvFlHJG3mcO+bIUz1uMLVV1w30OOe/9uyVk
YJOnnj+6o8s3Y+dSpnguneZExYWRijXv8uxYauzVQcyzId5GsllkjYAfNYob
rIcxIQtOD1S7NAEPVzw3/g7uK4lgf+2VC+xBa70rTnWEfKU6DnI2Kq4u2ulk
Rr6tgo/A5I8u0FKxqTkjVbtJ6BBN3yXZCPY6kPBBgpDaWWibwIGB32pdgb0l
RyLfltS7Q8PvufLhgOfEp7Jd/ix4izmbgAEsupUV8wwGjdKWlamsr8bWM6D/
3yPMQ/zTebgctVNihQ2lx0vPscAbwGs2a519d3sO0YdzdTRW4F4A+qOV/9fC
ePovv2wDkAhWNqF9cumILR0LEiXzkKF7OAAdzFM0BFBqj19RhBSTG2ZIC+lg
4aiMEdNBgLdddHs6V7z7owzzaWC60OjZXQ1izKEhq3aqDmzAzWivx/G6wQvN
zWE9VJc/Ao4wypoV/VTl4gu0yl7Zi9RvX+GjqQs3AjDY3OAE5xbU3k5RJ3Dl
i/+MbjMFyKqXfU7bodV6kM5EDVctvvsXmsl1Sfr4kRVk2aPi1CyY0z/aXmfx
0T5yVifvTCi4jyzKftNVLokbwQHO/ISYzpzpg7Qndzho3yDjGvnpxtnHO/dO
YLCnOFimPXZvxNcXpmQp+7b/qZ/8P+4PaJ8pV/zagKKipLp3Se1zKuxGH8XW
At2xAeYoewDEgpqVvH8PQ39PcFBKlBCPZXcY9GRo1o28fW67SVPlFZe7bjU6
O2TQpvvGB/t+r1OC6YYVyJZZW369a+kd/mDCNKoEWO5zo92qkQRENl1xNxxe
zayVPMC0QMOoTbsC+J9KTqFU8LhLhGTlmaattkrydzUNXeWSOYIiA7jNeobH
1gmSxQQA274Z+R9z4D6qrwfZYcB+pSxHcMP7Ej8g+dG8J+Wmn+Pu03mX3KUp
dXwnZ0rbLn34KGEZe7cqU0tXl+XKAFAhwQzhIgCbvLOxSCv0GHQGuMkkNwn0
QkixKDM6ickbMFnVLOR0ONNF0tKzB3LCOWhkWGhz3/U5a//PubnZY2me4aDp
4mfRHf0uLciGzQvavGKCdNE/V14f8NdeISa0QfLcQdGzKdMYjVDbzfWzF+d7
afl8NUojfFnn9z86y0vvhrkS2m2I/L82DXiEqrIlAUv+Qrqssv4D3OydsdGZ
bKAm6VvprI1HXS0FsvQsMc48yBggFOcys9w4MFAcahW8ueRtDCsv4AdqKSM1
FbqDkRmQmmLoyQtY24DoMQHYqxjnLC+EUC+zK76xqFy2E/u3vFrgiffm8FLz
UT/sKJKyWC5etf9pspEqfNXSsn24JWPi3WsJafCSTJz3JyGyb4zSCzvCCNc5
+2/Sz2M/wtvkvLbTdoLyBtJNPZdGpCalcaM3wvlwDLPvuEhv99kR67YxmJRd
wbR6t1rNgEYkuF03/s0GMKDCed+UXJnDoIpzKaGOyL82w8yIFrjRzjRrfHf0
DBQCrtRvtl5Ucozke+gc8KG2AbIwICAMZZMh+hBIRu0fH4Dpvj60XXoQqpxW
0n3FO6YqCldizPElhNeMQQSfxfcXP/JMB4nlojZZgvVjrwEdSYJbbtnRX8JH
I/ZsZKbIzgGwe/7itEdK+oLQUo47yJ2tPvfmwyzoLRANKsFSSjIacQKhMfSj
wALF2W60yCcUNyHwrxMHbQQsNexYPtrr3pcXjH1uGMzujzRclejVxbTdjuz/
Q3HLU6MDN4JSxKd7Aanwjatpi4LnHvnlCvi3zcYURB6o5lB1k8fL3F19zEGC
O6PsHfIbbLkJRssV04gIAWlbHL1DgE2/NeOFpzIsURVEwENwDoVGsOwdcfjS
bJpbXweg27LZCYql4g00LO6CnoCncdH5DDjQiiXbmvtFPymrD+86B4/VotJN
bayzIMG+mlbCKqXH7FyohPxGw06tOCTJHn0ZBINNTaqR9QV+gYvZdm2oDZY9
2NzrmGoc7JwxyBLbhpvh/OWOlZlpewq473gvZAjPPiM6LQ5Wv0EGxEytCz5A
zfr/W2Bz1eEvkcKgEIY40uoSxGfcAsXW8xr2KE7zGFm8cfm6GFJaJQ/tl5Kw
Qrr1wV6F/Yu/Q6F36r51iG3BV/cOE3dkyVbZjQewHFF2SUhdorW5NoPyDHTG
QLHYIHtHJXLKru1KzYf4ywhEGcacXpIaJnZfG8/HfZzlP9MS8cRTpC68FSuX
9iOnedhLIj7NoCS/YO3FVHngjVJumtO/adlPABGmgzLeanKuARjbtogmRhIf
YY5S7LmPzV37SU3b5SdGhMGeL77mk57krewDc1DHw+utZEPezyDKd98pxljS
7EpirDGxLpTkUee3pVV5X8O1+OPt5V85PNoEmP3Pns6apFYJLueIfPfW91kc
3vKflt7HY9hECs/6MCDEtfa5e9BU3B4HlxBLK6YLbLJLAIhrYX1+3k+8tlEI
MP0Wr758j/Lc281uXh7q1p8YiQtJX/t70z9ZxM8rgwpcNiyURX+nxnk2VEF1
I6hGBPisuYFqG7lo9lpQgoLqCUGTbSnI+Zrv6sVGPN0n+YiABbi8ic7wDf8U
sIIabruA44toc9yRwYIVxJ/8QYVabmO+88S6bKq5ucZSQDF2ezg0L0zRGn59
3dxDsFNWc7h9SIT4knXczNNIFQlxDkTMjoCUhl5IjIDzWRFSlo+OJuWPAisL
rhp5APCRefSHj9BnjTti1ie05TkMSc8sk1Ln+YD0tcayADS2OZjWxZkVVnOY
uFLDebrL/pWevConl6rB0H5cigzlOG86ccSUzV+/RbDNglgNKkZTwCgK1NyJ
WOt8j3PdF5p0afkn+k1/4d2xD2R62XHJHzHpAEs2Tv8X3IP/q4FfXHTu7fXu
afpFFu6Kj2AQcaBM/LqGOVj062OVfmIVQceeRFTfCrzpsvHf7lwLq+Y8i1Jx
53pFEHuzIxPN7S0Yt3HkCIJ7XYvnwX6su37RplKyUcSOrrXnKPSbidpWTj/c
wrltMCqIiUk9ANyIuGlbTP2JZx7Qacgo1DFJXD/MO8SaxEl71vOX0m0WsvQR
+AZTZJXNLR+AbzW4lFOxPf95VVGU6XVROUwMbWoTr/HYNZSfLnWFFtPSrBwZ
hg7IUVBcJg9O7x3DtR84GDmwyFgs0WuFJTiIuPPXOIM9VRjSTSWMaVcEH4hd
o4XTO/DcGZMms5XUQ7N7OqIcxaCb2x7H/utpUj/sIGOLxJkTqI6f9TiVspK9
V5O/uTVtHaSKJbLgZPKRaHjH8xYbQdJ/BKy/uplUHFNpAGajwxgI9DyPcSby
NnHVx4tn4IShUdq5G6OhZByvrrqRYf+kbTlsE9uVHKjls+VD6ntRTuN88oI1
/ZfIfnzIS2B/UX2sl+BeZSkqzfGCIz+F8TPyC3xSN/xSjGCbdzMMDV3zjLUa
/2e4cu5KvskWLh+NZZpEFEdS//TmP5GlCwokADub1W0gUw/GxC9fG5qYHY73
opLLAT8DT8JLWR5UNgi9k3TW+HExPVOV5OZ7/VfoUIeBruKOgtynrk1jZQNe
SxBel8v360Iexr2TTt+lc9DZudwj4L/EBeQ3zn4jFU9rxgiP/2+IFJhhBbwQ
B3+NChecGkkSxNAIC9cArv2kCiFnyZ9W3UmKXkPXNhRpArczesCyJgQ1LkYG
E5uM077I217NNfsThNNGRvYw1zrPl82xRF1Wl7QPGY2cVO/kLDeVdlxA9t/F
AnkBWazmQBJBSfcT0HbT3SMuo98RkVpvy6KFpokSY+HE9eKeoh6dMoRLIr8v
T7OJ6kPmZV7nbQa4eAd6BqT/tLxlfNPe7lOdm7YwL8c3/kps+TZ3GKUZeoYR
NBBmWDOEGaqMWFgFuqhMx18G+nvKlID1Coy80KsoY/OT/3GvMhzHWXn8HnuA
HUr3SaKbowT+wESr+CO3xzE3uZ1iyidS5vx6PIemye7Dz/NnNt6vEBnV60Or
Zgxx2uPtoVp2jQZVduTjVUij4/NsS50f5aJ4JOcdbBjPu0cwc3nnNUYBCMiD
kDAJLO7khXpbaHzJTmJOEPvJYj5Z2YQsYy+no6lT3b1Fj5fldSmb/eYKLqjK
Yb4I6JdGBmfD+rsWIa6OEEs06yn7wM0Ge7hjzMiQDl4iZyi46fB587tBh3bi
S8nohgJ99xFdNcjiGVAD9KCxJu352Asd7RZEnvax2P/WP9nLll6y6UdNFGiI
IFyzhQme00q4X8yn63GsP7zdhAJblOv97AGZcqTrdD5XYIfHZnE7OglrtFhr
Mdros7OjXoAvbjSKybjWmlgUrQ7al/CA5Z167UW3JF0pTXw2V0JlGEuaQGxT
YTRsLxec603K2+TrM/82/+/OUc5qTR+BBTmbD2X7qJVvYxi0vmI/a7nvj58t
gRzV7NxQcyllfzSXP1WyZV8nEqoWPvGVJZa1uS5YCIFbdsk63uVr7E5TbZ3J
LaybDfUYZBdZiQH4+S5YUDdiDGlZGOJhMvSpTvEKYTg00aIipDGkaEbllR0l
NM6KzsGtuAUj8WxK0b5VM2yimmfJaJNw6A2KGuQs53WtfYbnYzsf/AYwNOzT
bTPBvH41Ef+43sIjfbFCgvOLfzyWwcKLpAMs3kl5pVZGSTC228mtqtoUlZbl
9hRZDdi4HNYtixSVdXkIeQexzV1YKQ6MADHVXF+Sy7s2wfpZppGpq+P4HJjM
PjcAiD1Yzpi2U4Gi4SBgxNCtVUvOBEqc4CP0bXADveNHxZY8DMnU8SzBPI0B
QkUhw+jpxQiNSJdzoCXTSt+xl4c/95VyEdzMXH/7BMX+JRmeejIaamEOoD/t
Ykk4TQHJhQb6Z1NtgiD39vKaMbd+5uq+DDNpO5yh0ENYgvKezL0tYvZv8Gms
y3sVSbu1pZ9WwPTaItHjjboIICLwgpPzbphX7XQYpqLhf3oRhjJ4OClxLZIG
aYL3RO7aq51oyP79GWKGd68LlCs/TdRiFn0NJzCTtJa0UA/OXqAoNpOhi1uP
KcLiXDFK1dSmM+RT3r9W1ulw/HxSWRxOVtnZWiupQc7NRSBojVjJXjsNKjpF
SNNND4ktEfmQmizRtEvuBw1Yr6cvUnryJIboYCH2hIVBBJCoRH+KAMcsyUsa
xficm45qTkVYBf2PK1YF6sW9sIoCmcb6jJI5RcAHCJ2Moj2/ceL9oEO5mZZZ
hIpQnnr+0IPvhcIRpg7hiizDj7hzCL4KVqnl31FpVxDSFu7cVi+f/B2PMo4u
xhpztU/QkOXasSZFVYCKhsq2drr23hmarA7ksRHMfphuiffdE7lca1b3bbKO
IrPyzsYA2i+EYGFPy6f4fB4THmHXzHopyjEcek0wnXL2uj3BxE7oho2Cjsk6
T7m2fysV8iHnK3FwI5Ieh2C8GzcRu0DMz+WZj4JOLXbMw0xQgcUFmDcPcsEt
liJohfOcohsq2eKGVspIn/SZzsIhuf8l60MdRgqpr1V0Q+G4jvZvCWQ8Imfo
ZD3n1PRYcMpaODAVRNWKBSxLCx/To6+DoK59N9TblAQlnF+77XrtIQDq8yzI
FiiWSvChZDqjOMcW/8Fo8m8nHYxaQhX6mPG8mjfRZbt0rU8rvxrI6QsPlSlF
Hw5P1jobUsqT6uUaTOSlZgFBdakHMBa4nII7qLlgdB0O5Qh4V1ygP8WNirG6
PzV63VQL0ikYZxmZDe+9HDkqXCX7wqMBXfv6iid2Ls5EMxxiq9mxIELk9+u/
WePPDkPgSWC5+tJBIB59NZkv/Hyfi3EHVwgjVRdQQa/kVus6qbYoja0VrnI5
kajA8BEce05rRbkt3t7lJk+q5/wFSEkrCmnSQWmUt1xuGvx5MOL94lLOuet7
cfb0m3ARKjWhSw3ioUkKmW0paaiNDkTloyJxBe2VhHLEQmw/M0PNSzGiijSd
Z92Q8i2DZvDD81OB8q9nyw2WL5VieP6yOPN/KLhRosWE3tBilSinpe/KOhOL
P2PcxDl5e/veEIGmbzTMMW/TvaDz5ZhM2mPeczAcX5G3B9XiggiamDqcLqZu
NzUZRrs8FmKMTZg0kqoVNFY3vOJyscziEG5cL7QPGxMnnxokxnG+9CqikQBl
aD4gqLe62HkLvrLr7Co0cZoEyoVoDjIZntrEjJozJD2d+pA08soRK1wXieI3
7suMAdNxBP/earUJw+w2bvehL1J+8tDL8gY7B5M/iEKdKLCvR/CLZFOQBBfI
Fmb4ynHkyGWYOFM887iRhwso0HAodH7v1zzZ2v2C4TgLPUGi17hhdzgZM+Su
9eWGn8MbEfbINiibuP+1+085233vz/6V2ApD03+QtB+KgaUk4qfIPzyL+oCj
kT73DHcQgZny8RBUCLClSVNyIuperZLBGNQfxxyB5q2ZkmUqNsN6MQdNDx9e
dxHKWOmsujrxRZwKlx/PGSGUhfc/AFD9+tmIOG1nKC11mSGnt118WekIsQkb
pK5micUh1Lbh6etFn6BQlx8lPhccCBpOks4OUHvmb2ON/y4fni5C3Nui5uJU
JyHRJnP+6TVZZaYlW1gR9+sSvbo2GzNDZiEsFTBWbcedzDZcIQi4f8YH0xyH
irYQdiylubudQvqsn7X9QTKRJTNcr96ipgIwrseROP9pzOvfLU8tzfO1YiWm
cowzowgl9vHlbOMoIZ/dSxQefpe6MKNIgf1oI0qDSrl2hRcRES2ERYrirxHD
FvNvSVJaGFurmZrK890js645/9IYTEUD763oRkNWXovPzypCdnq4gBkGzgl9
0TqKsVU9F7DUFbtkcHnIr8h+lWHuWkonMS7NnHEcveWA8DQYP3hILvGJpvAB
F1aei1uGx3rOmKfbrgUKXaDHzcbG5C6Cr708ne3MKhTMDshyePuMMKUSF1ES
1pf93obQHdnkHBQtioWsjq6c6kjYEx67/Yqn5qew4hAj5KW+MwW+tljsWXnx
MmjYrp2X8SXMrh7JdYiF1JT82qdkFnkXtd/NpqvpJanWkUD8IXm7/g01Yuiy
Ad5tiaezG/zggWf7G77cAIaKe4Ek8dTKAfVo6mCezUjGIavkkhtwUo72AAeW
wPTRWGxBEUQcPnYgS14Xo0nQSlGjTnqwRAesQvagRxucEl/2/wQsdBzQQLxV
K/m9t7fu7MBQPoE9uYIJcZCUYfp/VSPx7GQqBoqTnNycETD1Ldsi8mrgTnPu
axx+SMgvhQ2lk1wt8C1WR3O+ottaR8B/hTkpedoY9q6WhFw5WZEeV8buhuPt
LNsrzyOeQJc3dt4XDO2hwm6Lknr/R0DrEgerjl6LqyUNvJ6ibnfs6jjKfDvP
/TM6y+CmcvlRc6sMzQNvyRhD/rNfCC7g4OB/6wltuxo799OSCEgLagm8kG3s
9gp/4OL4sqYH5JC4PB/AjZT21vis5irtw0TTKM4EE7s9mWF1cveBNsT/jNUp
g1RN8yE9/tNBdAdmFksKRaNB5BcIvH8jwLfugVIELjtQF7bXGfApar5Nbke6
T9zZ7IF6y2rQ/EmAqQYs5uhe3pSIlM5wbpE7XiTLalvnDNRgZeJIlSN8CNdd
BGqOXPZRnIpRw0/+nts4RQTW3X3kl4PUEZIZnNx+TM2fzV/0k9OMfkZDzOc1
upbXBMITWxBVolQK1Y1+q6yHeK/Y+tagYqrt+y8NpMIfuIJ0eH5wC/UCKhkt
ajpdioQJ70VK5DifGm5extbQj5kMyuiHScOcbs0Kem/r2o+oc51jq54YoMHU
R82/QfpuEihIyZ/VFk3UTVSWQrjJ+0zmNJHJA6ESmCpmhBFpLkQoRIRbWy0W
+SwwEGOIxTOsws0MqSJahJSv9IJpDJE+97b9zLdwYz3n5dmyjwJgAk1UsH0u
QuBORxzOI1vVatb4ScY5UHGSrCQIBtADFBrMRule2ANcZJ7TSEGXNoPvhNpt
6P9DXm3bCkM4/HxEvFEw3z3HIECFaE//dj01nEPTSo5ODrZ5bHTUxJNLGL1k
cxmvlARULUfDLEOf+n16nMQtmap9NS4ubeY4Kd38bErx43+2dhiUbgueuEjj
T5Jj2D9IDigZWLtUmt+1rrkxj1W0vwYjdvovif9diUgbc5aHaLMJF4RDtVyD
3QsgvYK2/JP5SPFsb9SRqNOXT3mqvH8Cg0C98F5irwSzyMs5Lj76xYKffUe9
iFIrYML8OGz8pO8sKG63JI5NmqcRAbeFCbacv40fjmIRteroC9RRGk/EBZ9K
AAKLBfU9onBvjdqC1PX91w98eQuR1ISLDWuWajzfMjQCVlpq+IEO3buoZFS0
WlIsg/2wbcoHgmcyIhvkK9hbVHMbPXgNQ8XkRN0OrOXTNhDrYY4g7OQ5oqkK
6YNfiPa9rIoQ7HHy+y5PVjWUDMNbToQrVxvab24ZY09qEn9BmTvWwOXqX/hG
yW1ao77WqqeOeA0vZr80FlBOg6X4PTegRkVW4RTzIibw2os+oqgG/fsSNnsU
DMv8HbGFLCXUslonWPI3sqJS2Zp5Lr26qHHMVL1b+xE+cQ2JVs9KgmMqdqa1
/S30Jd7Xv4CZjoFNsGif6fGdsx5AOMYowSg0raeTPW7kv/4Qf9zDuOpK35O/
z4rZ3EmcMHAMpI14yxKelQ73U3GP3QRmfx9jTpvSBuUQJYmrpqt0OE1oLvTm
PXX3tVcE8rr5/uhitUkX6UEkwt4Lrt/11HHeu3TGXAJNnXnjHEj5dLRu2IGP
PMSMVw2RmUv3444rLwW9RSQ5t6zmEPZt0UOSaXvzGesLOwCtjkdv24Q0KA0G
LkWxPezfTbITPTpWaKEHr1x0dIUlrPmuLaxfA+PxiQlvpzYG15QrSkKgdHCE
actCTRkwPQHZhRzqTwr4sltnX49Xdyalv2K+Kvj/Q1LwTfX/gQJhOtWXlbum
qImUfKGtF6wBlO0/bv0BYxrJtvpcGElqeHlGWBQMw/LVgSJEjEPvMGe01t0n
G/b9YkV/FvhVk9qdfLQMaXBiwQ4XCr8P6yak89OP1Qtv6x9KapTTMUQaighK
cCbAfxtrQL0M3KZqM476+3OWyeBiPbSgJk41FFZQJDaEavGp5lwjVlEosQrc
nvgG8W90eDOog8bpUPZeyug8f4j4QcunTtVTgf3J4JpMEwWLD1ZaW3wNnaV5
Obo1Sg1g/cXfsUnoPAUQ6Nc2M7qWOcpUPveRAqlHLgl4jd9d2DK9nDRLViZi
V6jwwmgln2hVkbR8EvVjiUn9uLnh2+TUKfZIjgCPr+Lb/zkZZ1qBtrz3MmSb
Anae7yQav2Mn23T1xcC4VivnZdwx1kJ5oXlKRjdolcdumBVww1WshylhK+fe
dwjIvyo9vR/sF1/bX+WbTeHg+6ccaqNgvmol6RoSzEgJH2VYomLydhS4PwvX
wdK+cSpOzks3Np7EN6Az+mKQu1rAA6DQBxMHyQDCKotqYc9imMcUjkk1qKdR
GbKIVFL2KTUfBq0g4rJhd63eHvX2m3kQvBsBf2y7TzpuHYW4nycDkXpsT30X
olsYkDP6UPj15ZMP89BvMVysfRCD9IVmdA+MHFRmGPY/kH83r0h4sbSskGkw
0sBRIvGwRGPSTItylOF6XPjYBRoOprM4Ag+LtBQyI4FIssXKzSXyG2duJe8H
SIMGp/JerOL9gHJtlvt6uvHrmFJc/TPJnH7VOmpD7K426Y6YFq4wky1n+57p
/Y9txxKqBkj7iy0odjq0oGKDwNlKYOpXljHELfqWoTCFexxb5vzJ4Xt03CaY
UEI9PGdFT2pkfxstZ+kEePkauzDc9bM5+/0HBc+4y8duF9GhOWgQkvHS80DV
gh/kfu8zLGTIC54Xi/wtZ6Tpnico4S49rb6JOhy8p5QeEtrg7L0YB5NNxZDG
MVwX85VIFppL2R3JWeC6POE2ZQbMZadzWiH907x4kunwFaw8ffBBEm5WAzes
S/s/h16hjpGM4PQ6/mhnYwMcxbW6UbI88IBWW37U2UR2RXst+WHt2i8AvrFd
U8So11WTe5NHF+3vqQG91zAKJ3lhBLvdIpTXLfZ+ieEJ+zABh5KwnC2ndXCE
U57QRqDe09nRSyrNdsYUGW7pte2Ef2N5LYuX0P/vz2HB6tMyw2UxnwsGzdg/
nRxv5955pez2gFHWxxD6Td/CcyFPM2S6o1mZtVkNDi2drxPRsIWcx1A9HA8v
TCHY7vUylq3qvrkmzRUXIUwGEsGoHpv1dvAfjPNfg5IysETT9V1Pm/Bp4nn2
pZMK5c0aOm4EGaRYMX7qR3ZTOkRC7JLb4h+0fnGdjreQ1iegoaWB/9ofV+oD
sl0UyuJZhsltZ8niNHuwMl+GUL1kkw7gKMcNGmzjWR2a3e7veXYR/igS52hc
/8cVgT8V+MvVtG5c1bwKHgttmw5XGkB1CnSXnmwd2C3L8kHdTzftZU0cqPjg
09ePhFKvxMF6rH/os1RTVjaaq18hoPzXgW3r57S1R2E0qDyzJLEM1ANgEwpQ
Vr72sVzHdRNdJnC0kzOqh4ebxvbsOl0k5kG3q/3t2ORla2KXT0MqwVsct7eC
UFROar4Giun2xDB1r6j/JJt4kBo0lqoHEeeqhtfM4jLmCBnP2O/Y8nua77ul
AGuB/hAWitjWQJjZtGQIcSuy8crviTdsdXw8AUj4vp8e8iiEFrqGe4o3MLaY
rvpXaJSO/wPYShIPRujCW9Aw+lNipMj69rTYYIV4M89KydRxGzZa55gnGo6J
jmqBRvJLZmEwPZdvPccXtL8P0rdygZ+Hmuw10Ap+8iWAVbGsOyyNoa3RjTMP
bR6D9X44gxDeAWAowhoFk8JV9UI2bvJ4na5JLUuCHalYx45NReVWLvEVxlHl
IUvpJrxih+0+TPOT5hiyqfykvmd4rulUIn/GdlNnsXNLbTxKJfK3A3lMaXd5
zdwRd7g023qgoTAPO2TABlz7AvwNZB/e+9y5qbLNkxvMfqD5kbtTgT3UNFN/
vaWeJb75C/VRGe4Xx+ZK/leQm2Ms8DHRE4UxQqOKFkWB4McneRXEtjG+iwRC
Cu0LjHxHZzKyyTcaeMXcOaEhpSSYUbaVAUdQoj4OEOWStphD1j1k0PHrHSs4
/DhpOkEZGgeolwqRjbBn2DvwIToFwE3amGa0JD63bLz+VCrVsF/ElDO2606G
wxKcMO5QxsL3ORxSeF0rAhogcaEdrbvnEb+lv8/w+qdBEQe9GPXsDq+pgWME
Yfq4gJfQENLEwFj8k/qvfpZJQ9JGPgWXpssa+yTjaz4C041D5TUlm4LVGIz3
OX1LzdHyx9bUNgLLiftVrg2Xto8ZfUIQV61EwmEc7Y1ZVZUJN33kIJ0Ov52s
iBpeB4Y+ZxA0ggrBy+KOhqMWtwWzgDtLogARxUEe9FmOeY/tBSyqiFzZx8Zl
DK6ZmDHsgDgKSRalyi6IWQfhKeV8V+EGb4nB5OaGJPoVx1U15baQ29v51LC2
T6IFA0d44btaHwsCTdbKdZx6TfPYBVZfvzHUL0hI+HFI3UwH+esC8GihfNgy
t9GjecjU6p93hXKzyBfD5T0Td9tEKJRsp/KxzuXK7tg9qTAF894LamsmeCEZ
YQvO5V7JeT05VK2hCN/co0B7Lm2vJ/EEE6m7/TWJkGdsnxiCOyv8MG0+mS5b
PMws5CXVuIyNxb21ACqLEVaJlyXoff3LyVz6EgHtDmizrpVopN50wRJP5/Aq
Tk5lKfwKozXs6Gr/P0lpGIOgZuIHQOMsCXnykvc5SlQMJneYCYdHt/jfhEiO
RA412i1bhJULZibF/SZbPm76aFJcw7h9bT4Lb3MRTIYNsoNee3st4MYLjCGx
7AtxkQf0Bk3QAiCMDfs5vM5RukSw765igdKBZgk6l0K8qfh5sX48Lu/2jrq3
AAMt/HKCCauBwVuOitY/RBMOTeiXXfOqQ/fpEcGtaltS2KhgnwSo681cMqBZ
PxaCe6LoSgNNcuBUGYvVtcUuN22zuzQcnwJ5CaJfHlUVYSeyoT9fSF2YFegS
GHciP4uAiAL9tl+A9BUnl+Tmpy+VyT+2O8bHgjVLO3LzWt3EbW06XoQ4OROf
9iuqp58eVGZd/FOkkFgL/NdOON/ty4K7iHs1qjqeH0/NSatUhsCkxposDkO1
dU930iZZ2UIWJFoai0wBd2JOSJGpKjdeCGk3wZ2+mmFrES7jzfqV7/j83inu
3iAW7qiSDMwitshl4of38waBknhVuZjefsaoz8RdOWRXDGyWmlDwHE2OAyw+
3IS9ABoD1VVMnyVeN8L6tO6uStXZbISnf+I4uv7KjZ71zXGB5+ecXsKgRypw
WWTuZCNmEeeFvUfuF2j6WN1OHdp5n1/OEf49nzgJSC4t1NnfSapeDuHQMeCw
osikWZ44oQowxBwYKQpybGgFuUR9qcJNo45XTrh++KU+fdnAPHHn+xeTd2kX
AG+dpJdpuPXhQi620I8Re5Z5c6w+9dCeVBMpPKTpl69TiS44/+IbUyzlVw7e
eX52ZLfjzayjRNqAmfJP7kZ48blN702FN/fM3H3FL4ZvaNTuK/zISdBVf7hM
InHMei+mTF/lJd5kTYbAIAl7ywv5rdvvaUIfR3kpEeSX9hbq0w4jLfO+bZpb
qO9wGDc3sfQe9Jrepx1W2Rroo2dglwYkELd1wddpzTN3gZpYHwstimaHzRFr
u+FFPvW4WfNA6wsMJnXlFdyrbEzIimdr7X4sh+DUenT9ydfQm2JeYS2dgbDN
fymopSxv64WGJeF5SyoVG5j8iRl426z8EurzSSrnYWBzVGhrMdY6n3FDO50h
IEM8UJP/pnjdWOBWLGadkFm5dF3AMDYXK3UJopEobp5yaJrVY9x2FwezFXrr
rluIYhs2XI1NQ65jmGX6wS7OoPtDZBoSsvhw12o/S2bo0KQQp/Mg7nTeI+N1
oArxgXHkFd1kOPpjikfDMqpSDXOrta/PNpYQ74RrpTdJjczYxdR+kxe7f+GW
dBzEdRqgbUW3tbA/G1Ww6MTUw2YQCbZ0GyiGvjB5qxoQ3ccGolD4yV8aeONe
4zRybzKbU4mZuqnK52MNm0ea43mdshD+Zs56QQhspp8lM5e89EfzwU8KxWsj
anYByt2ECW1wbEfW1AfpnboQeXZdQO59AT/2GXz4UivYeK9qXO8ZvZqCtoB7
C9YwFuqvig9GD/CdOEbm9fAZoB5POkR0D42jcOVZUghEDKB9G74M6v485i9h
C7m+cyAcwMk05mCJSt2+Xs+DlCNMBFBiz4tY8A5pqYhyUZ+sA4icX6qu8XlS
4Yi+e+p3WMEINH8R0KuHySN1JF6/zqA9RFXXDGTP6h7xlAz6TCXf4SStLc1X
ZvHJJ+nPS+oxgoDJY2AqNd+lTkLnhoG3Tg4+r3zGYc/zMRE0kMkY4WX4iGFG
VR9B4L5Ep0Ab7Z8q/2ApZQDPBVuEnzb1w/3QsxIIft5FxJnPwI62OHBEyL3f
K2Ua7rSjVCEj3Ta2uRFeL8x33jEcGzgYo2lh3Py0VdXpCODiescreZgJkALe
wXcPvWnKqJMaZuOENgj3rcdLGc+7r5egNPCk2EbYyIZFziX6rIWEfhi3Ba2G
TXwqqW+MTrj8YtbQt9XUXDPrkGTKpVEqH3bxzjbjrE/UK3s5SR/YBP7mo2IE
r4CAKL0Xg/AaiH/dvw0nhP4wYDtejcS1Fy11ZjJ81pRPfRBpRgRsOEIP7YPG
ctBpcg5IV9lSrGygBJ8CCiyZV3LYk7TNT+pore08wTqsbXgFfU4e6A3aykzO
hP5/zyD8fWTqhxI9OAA63JB0IErWs78NXjAYtGkF9oJOktltO13Zzu3fjJ16
sbC2VawH2mUeYwVZB+6QqgIZfD0zZFHeSde1tXp0nDmaxYt6u0j+lMGQ1qjQ
h+NZzSeg9MPNse8JDFjI+pP/YUNDa66UsVdj8s7/quUHU+IZW+xUIyPbpxW5
aEsNwmUE1VsDqfxdJMzMp+OgbtFe5iHVoSmJg7KVnA9t4cTANQl6MbRZNeJl
y0TgB9Xmk/6pblHB5/JcQu09tk9nFyDhjdiLFx0KUQ2Lh+bg6/FI/TCvochg
z9OpKvU2+A2kNZqDKdU/uCwvE8TxRTwXxTXlhMcL/9fvZLxAomZRp81fwA7E
imWHABtXFwKG4cV8QHldnpi5u+ji0oCK2jt3dENh05/kFlfMUKQZbehNdPKP
RVGJ2shFX5BDoiDOOtu/BR44yGBE3pjJ60Dzs07mWdQv0DLjc2NSQdx0FBIY
NyXhC1AkxjxNvTGIqicOcbymprfcSI1WEA9TMvkD1MbrrSL6DZCSN/DhFLqF
J1kPccitHDTdOgJya+Tqir5XBM0jgwtSpWj9qr0VJQnZyiUwCGpdzqi06Bjf
StmxB9I+xqWJBMmJZ0kmBqc3ufZ2x9QzE4sK0QlXH/I1URi8ssf8qllVOKX8
1wiz/uUkiWFW7mGtJxX8gx7MxnILyf0p87rhnxTb0DCGjsLnXM3fIUJ9QZDe
fxlqxSPNjaVUR0+SrlijqtFexmHjiW2o4f6lvQ+Bgf67ArWdec2fvsU7HGCb
xkVPH3UY2cyPyDponra4LjLx/dqyKiMcExTlPq2Un8l08nfpveZxBg1M/5Wn
o841cLaXUMKEePRpWK4EBsfHNOqcfo5e8Lv3SNQsK+EZwe+w5RH3xRa9KbZh
i6tIAul7fzCLO/4wGIaxcolHDm1nS7cViS5lESsU3k1DikvMDpKqhH+J0mxC
mK/97WBvGo5HzJs+jKzX681wPr79/Bk8ATa33Fs6T3P3A3eRjv2/2MT2iM0+
FuFDmq9BRq4Wb37UPrUXRY/Kc+tqiOwdlj+sUu7k81a3OaVyu7aNPJ6W1GI/
VO29pht6vM0khLtJva0KfceroACeQe9dw5M0u4d/08xhSCqzXnNIGYopdHVm
g96etAcb5tE4bj3JVlGASfrBACBzpFVonpyy9pZ+D7f8HSgUNpJ3ZZcET4wU
qaghUm1KPUB2m9GJ3RpFKPWJsQJRsgQc9IUVvyrJvcJozvABbyPdIzX/UNyW
FLtoLeeLrT1FAM9f+c/Xdhmvh9ZgZj4ME0st3ALG2gIvk3MOnyq32rbEJ97E
ivGkosmTyrG5yGiuQa43kVC55lIHDZsCcZ1CfnOpyd2W48skKLfN+oGeb70a
M71BeisSs6DWB5z7Mqmy/6Dd6d16o7BSNoOPrbXwb/K0sZojDe1EV3hB/WDk
4+5ztTTef793FGGAGPPFg7NC1VYXfOPaXpPH58yFiTj2j6ZFAxXf1+tLhvad
ABo0ijgqHht4OKroR1OdDpEJOqbNO+DgfZT2a/uRUxKG52MuTeFUoKl2mt2W
ManIWmnUjvOLUItldWNh20XFNuaySoQox9/UXRkjf608hojvn6xiU7Qn7eQ/
zmRdPjK4edGgi1oKQIAxZYjPy8z+Mx3gzI+bVg+dc5cEsibIUk7mzqSpsnYY
6hJP35gX59dLPe8V9l8FESvys8h30Ap9sa+WWwDouN05GM4WQy8Q2IV2r6Xz
1T0akv6bf5MtQX6Cu5GLD7ttAK1yNIFx4pE4bZuehdRfaYDnvqkU2cg6188A
kve9GlUPxab5IZK21FDW5J4Q76XeWZL66aHZmFGyZyFCKwu2NT8cuMI+sQ6L
2aCfZ6SArjcmHCSEkZjOPF91MfzAOvgoiod/eI1nNSNrZmGD0+w2+LtUDJGh
vOVNn6ahAUrIiwulvpWfj4nPYsFBEmFbHJRQlT3N0wB2RdCXeNuy395QYrs2
GBEAC6IG+veIjWUVgmDPVoMyQgF8W4Z9OVf3ZBjY4BVES2KRFcSaAAzJQBl+
Qz/clgrJXNjFRVFMilsR+f6Cr7OAkqTd94SfsRS5NihbvDgfeJ6mbsp5GBPV
NDPJwHofD+LCm+sSdz+wJNcuCNA92keApM62VTnY1GqXQPsi0l0u7FdzqOy4
7Tt/LSLyWIl6+FX7HNg/7L0Jky/Pr886djpYRpZNSQhMwQUHaHl3PlNvpkek
yBs0fMbNv31qSK/54jEAj7JFL0pGaqLMo5FtuW+7h6xFYZfbl+pfPImwUIsL
L0AwkeFVQ3BEkbv2DJ1eKuzGg/iqb02D1tj1i/ghyvj2xeNcukwEkm3gpk+d
nb6M33TFJSI7J9t36txfieLm+MRKf7ToL/ESSCiiPE3d6/5qi2eVYzIg9MTx
gsMGaDIbnUWgw5g5fAzrqA2EMsIBFOT857pUvS5TrFjBNxy+2bAgUw66Zfoa
74BMpDcVXEsDp1kTtPip9erKrHBLkTD/rQqKnM6mlXYwcwyLP2UfFmCkq8/1
XqpPhMYbrxT9+TT8GdEA6fOR11Abx/GpczZMjTHfZd/vpRaRA/saqNBC+HRn
zDza9KR4PE3lyaXMSwBiqLr+QFv/15zP0qPSwWxfEd1lFQCIX2kvLrBG38/g
SXI7bwCaZ5qMT/h8F6LHCndFmEQGC6LPOqxPV5yziprSRXF/KksSicbnkMVa
BPr7ZV+UqL1xC4SKnrxi0SmoWRWB1RQBCPDzV+0r2E/j3kH2VLftxjeU9Ssa
GbX8NOlo2Kl17bHF/qw6Jduy9ashp/FwXBYIwyR+Pub0LyIf/l8Zzh/BZOF8
oez8L+vDcA3PVCCzlYLjnjZT/R27XY7S4NO7iC6rJwWEoI7DbRWlkb26MxPs
L3xoMMHV2yj8Rls2unTAuijfwQEyje622uY4YDijwJ1v1MttQOfoqLB0eyeV
aKplJVP2YYvoHG0j5e6xYNXqkIgheuu+dMedP+6CW5WjzprRzCivagacyxf3
UWVYurNPXdO8GxR17N5QYe7lRPk9mUV1YvUDdzTmiKeXPJdf2gD59pX7dPqm
iN+mHaCcYKmq0f2QKBtysRM71QHblIH5U6RlKfRFkfByOxaZ6m+SWnXWbCd2
BrLV/yNkcvY6IizsYXY6bY8cfCrakVSEgGCJEPbZmHIlRfVxQ50uqXwfNQ3e
B/o3KZ0l/ryesqIUGnFSoGVRzgd3jOBt2k06WEE5dYK6aHt3JvHYySY6zCqR
Fl491gfXJpioipWclvuZtnqNJj3O3X4UZuQn61ojihcjLio5QId6yclGS8IA
XujOq87UKWIILB7lltYkYCBpmry7DgeJy0aBxXbyp1UxJjcO3Ok+wOvhcLuM
5YrnV7pN3LVs7eiBGL3+mQMaw/3R+IvvybxphofaQvTo59cb717AlH0QVTQd
U+CofIif4MbqWJl/C0aZTrMyJvpCqgjPaMHi9H17Vn0zYnPy0tICVkT5dio4
jPr+Ba7L1fGd7KIod8zgfNN75KJO4uEpS8Z/guL1n7PnjwG2diZPBB/jeVyM
Ucw5uCCvnCuI70+IaLsqWSvc93qrW3fpX+lsqQLiNk+yTzKhz2cwRBo9biVB
dTUXUQXd5q9lrrjF1oiMepGTsYsVdNZTHBOwdi1TJ/OWyZ+uD1D0jDuYX1Wy
18VTDwt6gdO4dtgIduKG5Vc6sENCDDJdGXcjc6r8ugkRJabLwYke5+CJufGV
GtV09cVQpiVEEHtYyyRI5cso9Iroy/iFscjT9YjgTWb0YqezKn/7Zc+w+MpW
nK4KbXlOKAYdWAgkj5leRDJMF5tr0MvyN9tdkovGxs8e8RE7Ax7sSWQ6tB83
zSUT0UQk4Yq8AcBpHHYdW4zV+sQ0T5E0hBM8aPuvyi2ZLPHwiGGnCwAwo3cA
6VWgGkdFMopnAHV7d/MP1HKvvnZw3szZv9QJJfyZCjXkp5s5outpkpIC3pR9
3jiA7cNkCNuHEVHlJ6+cNx+URTka1ewGcClrZBbRVYH3EszdP3wpq/lZjS79
NgGBKPgGzb35uchs3eXhwUir2awZQfXkPyP7S2Mr8HPejNhlg3Gy8EIvCi/i
UGf1Pu6Tk0/rW025DGfgai2vhaw3i0cQd9HXGTok6m42DO96Cdct9EAZo0Rl
nwLBNBHxr3+6h6cmuCxsYcOAFu0FUADQ2KriK5V19bzkZHkYxeUa8eZzkS6Z
x5+c0wF3VaNaiUBKF3AJKaV0pVzprOT9Q6cKCr4ihfaVs6bSy+1HvySErgoF
K4qAjxDgU+pOV2XykjzGYrZYSSomZX6JXESNpk5e88cbmTwrI8lptqzqprJv
oCaYEp8jRIB6iYt30b6DYALsm9vl4Ml7tdDtxu93DwBZLE7bSkv9D8mxbUZO
ib/FELjZd5okDQnajpCa0aRe/DE8fcsmEy3zz1PaOrEcHyQvYX/eTVoKcPLf
tl+NqfPkGMMu1v0iTz+0HRWRG6db2MdBFpfv0DSJxfY5VlNGW5lsa9fUA5J+
dhqDnqpdWwwf4BJzJBU0oqzPDS+8OTW7EnsmqOClNuhLHqkRcebmOcDHkRZF
X5iN2CBfZAiertxm8HofE71FpM3Ua0d0jEJA9PRIzjwE8oh4Ro1ymBlQ6aWD
hPB31jJJBX1WRGrU/qg1c6dUHuvbXb8uFLjauV8AWx5EEtbVRkDbb36PbU5j
I9yl09OBB4ywUhRfqe6OdDmuANA9xUOjpRrenYso3jsdZKwI35LOlnFvCQmI
x+yTszkFiJb0rDk+4tBxJmE42YosPwEoYOaW2o8+2E4EYyZ1qPzBJzpmV9GB
ld53Ag6siDuD0NtwlVarw5s3hUwY0s6/9Gh0LgoalZ5f7Gs9SOs0Memov5Rf
ZMu91Aikb55Lz0yJH8N9EOV7HLJAFLXDObalXIiv4ntfG1nKyzEDFjZtBUGO
hoob1q6tGfE3pPmhckBkfRAuRlux0QmmTxUxrfUxX2USBJZECHwMW2u2uB7i
bBAzwclzzYP3fjptsb1Xv4iBdeWbFStMnNQhdCorFdvSH112uWY5DG1rk+aB
sPkqexMoqjzjqKxEQi/zJ5yofGi2noQlrtzqXarESZUC8rg0ODI/xh3yKncV
9/eV7fCtKo7QRKttBk0CB4Qt7Tvxq21mnrCEKyQ7cDuwoC/cywoOmzMRp1hV
dpeSith+ptVfi5dhTubCDa2YmmOszNuBDZ7FoMR8kSBVojI3omG3ox07A1cz
3G9DzTv4FUGfEF6Hl/PYA53Hu8UHE67KpoxyDwMUBjdUy8FS8VdqQl3i6han
BAwN6InNhpOI2v2iNvFH6h8ceFsnd0hKeogaTlUdVmJZfm34wEYbRyQVVBSs
sYbfeijXT63y5AnUT2BD5Yv3UCIBn61pI2nfNHV+Sfq8LTWNyioF8UqHCSdO
Iv+FNqdN+wUDuuwmdZk4vfnfgJWGdgk/bD4qCx39hm5cFmHapwPyCFGDz7Rx
JuVQKJoe5utipa+2B4yH258EMYwtJCOcpXlAUhZI9+ogwCl6P+6uIh1gYZ8e
rNN9DObbfdttM98miUHJjXTvkhKYqP2AabRipl5n1+y8mMC9xzYBAsJ/YiEL
hfzLE95jUMSBVT17KBwSt+ZMXGy/SO/aJdJLcEeiMzoEZ2PnTYjvw/8Y5RIG
HSvcLc51Ja6HlUqyGtbe9X/wwc48k9Wf/2myHXMhoKW/4c0EIzGbTDe3G6et
bw84GkX9Ls0QXOzXsz3YWf/6DA1wlEvWda30RvYwVLbdmNX/+w14dx2gbysb
SX6hF6Ca2kZhbDs5fAdFmn37WffqOLr6QTOL9Meldu4CQHrRXeYTuSZiUun9
bx/JIjWueJ+pndPPaVInWZNUlIodfvYzoSt5ZZsIQH8JV9k1RprIx/o8X9UH
ZE3HHuhiRjSIFjKE822J/5OLw2e4maAGg5cHQshgBiXPywagE/dcZc0/w9Sj
SKUMZjyFxIYOV2MTkXVtFKeRxSQ+rYzVB/XqGgm5YL6tAqRgYlHwPVGrNdTf
SbcXGgL3Xjcb35vin7g4x92WNLMyu0Me7hsyaeKWJv+MNgsdiqMx8943SX25
n/z+Knf/9HCE9oZEO7jRsvK1Di1+yQIHqQsrEfEfRX16veYHranjVXIZcMy7
lrO1lbx1UG8B5OExvvy/yoO+/fdk8ATasOc6kwLZYCh8b3ZiQ/nJnrpaNcXC
uISQRRtoYKr0LSQGA1gnp44PqW0UU0apZsbhxkjQCVCgcamzCjTbR2ALrRkA
0zX7n8PhF818x2eqRGtZDPZZ3qwzZB0YLtA91IZPZ8Tu5wBULd9PHL8Aw0vJ
qiAV+TgT16mJHsIVtXbT2MCr6gQtHVr3iIS9eGr3uR2XldVyX/RlAARFBeLo
o8aKWRuGFxbbnA11s5LTdv7v7pEbDQ+VnOY02N8ONJgOkZ1CnOSXs6Y8dMZe
RYoejcC3CiX/mm+N2r4q5lh+sME20CTrvyhuDBliupXn6SLll6rxwMnQ676H
uq3qLWxoSvBZxf14jtTw8x7fYl14J5kAVh8RGj0AvZ93ptbHufEErZETU7Ru
CwfHx0/s/D+qfkVUY1wK7t2V7yZSI08TqqI0kYMv28/aptO/a6lRnTWVjmiy
3/3FnaJd+DJaQhPWBVygqy58pPN2LWYcua5rqqvB8Te5YS6/x0wcMfVPBKIY
Xcx5WuhVmjB9FRNY7cZhBJaxYfY+rLkGLSZHwIzD+DBjBnEf4Soh3kp+T+kf
+aGBAL1lXH4Xh1xzuafx99mI2OBbI6f+4h0a2SbPesBgJdYPly5gmjs2ZNcy
E9TVBWuCv0+zfB7bIzKL7Uqnrl2PRuNg93vI0y9O/+2w707SQ/HkDpV12Mya
ulukhUsXqjBHoIkaQgLFImV59u1Wmb9vw+GkpwEwRLHLSAyv0HnIcYCYXey3
7ZHt6JHuE/9/hgN7irWJxome6947bB1ONymxIrE3fKwX8srQeyRQ9D8neOdl
sIh71QZxXaXKnR0lMrwjTT0p25esRdiCCCB/9JVW9IrKN9QFo4nebtixjwAq
l0JZ+WMg4JyRV1FzIbg9Yz13OQQwoG7cH7Dtai0b6W+ynP8xsIpb9xq44hxc
4Js5UWLTxUzbYKA7Se6nxTi3tj4wjUlfM8fMBgeRjKUby398gmqWVeDlajOV
mEeSW5nSVo/xoibSVUFzGGgwK5/b3rOgBAySZdAlT8vf+JqqLhpeYj3sIvKw
R+OtLtS3Id+0J0Kq+YlrD7CU7RmmSi7G5ObLSQrhrlkzdrmFjVpb9cPKpwo8
LF96m9wPbEZOfOn4zNyIToaRohUHx4n2QqPtID0Vu2dm8deUt7BKaBPpNdfd
Kiwyqnb/QndLpF05djo1ST+aTZ/T+vmfME75J2ven3XV4bPN3CjHaWYeZ5w/
6EZkE1wW1J+CdQ/qVB8R+6mZboO77aIdY4Wf4vHD+kLr5MVWOYarM74aBSCy
kwTmKwZo4d2uz8d/CXqN74hZM8Rap1SVHV3UXrm0YQWSDSonmTDaAIqBy8Pd
/CXltiUEvdCPVVfY2ZVa9vBzz3ZSYAi3mkTWKxFDL0SMLORdcXdPPE7X9dmQ
yT0M8DtFu6Zg1e6ak4szGu3JMmNd2RArMwdeIvsAxaKcbKpJVSXvoNuDEkUO
yzXtLaIBm7ZOe/BvjMSbTsWy/0EmL5m1ncDwDMZpioTwJsPyko7FZX853dqB
AOp2PedYPJxyTxfv08jSEGdCoa9IKFdmuMuHwu6/5AzWM5pwLlURsY9dcpqp
yd4WhTn4BzhDNt6rt7xQM52TrQewycFdsVqvvccAS62K5RVm50bwp3tm6k1r
lsN/qzBT+Dr1jHNSWzT/mbIcxZACfpbAT5oGSdymuMHtSvj4tiyHG8AqogtH
LGEygeOqg+ylytFIlBXF8jGegEqjLGs7GzbhqbGS80F3ysCm4igA1BfFoyJN
igYDwMZ1NWjR1uqa62Cq/fkZreEjzqP3CcatgmT3mb9fySoWI2AA/dq9Kzv5
JYSWwBerTrnRR2B3h00LR4z/tpDV8CM5QKr9tiMfanVY5BAhsppJ0FoiXSrl
9tdZVgtGQ1I038p2+NOf8E/ZiXhwOUM+hacjFfYSiWfqp7IskAKl9af/i84L
5xswgvgIJQD6aW8SqoNv+T6CjoAP+EwPDcMQX7czaH5l0ohLialsPHAdgmfj
KgOsks5ivj6I3hdlvRV44Ddug91QNJPcAuYpE33B+2iWzZUNmqHiE17GK071
RtmTpyEulPvwL61EMEhbMpOCgyDGdimfxz7LHdaqQ5Z8IVd5t28Q32b1B2Rs
jhkfUF41BIlQ2or7Jh1FwUIVZUZzzuFmy0Acxweq0iKWt/6dJb8WNQNgy3QO
dF9Rx39M3FMeHRQnHGJcBN1Cq3hQ9II4J6KV7tirlpZ/7uaHLBWTjnwODBmx
0htBVkNDJa/u736sZI/g27XFcP/dAYFsV4DAc5nwPWZasueKyIbtRWZO3fXU
019pcT1d5Wsged6PyHx3iy4e93QNO0aYwuXE2SvWU0+0Kf63ml1+Wu49n3JL
htxzWnnJlPpwO9EjowcFi5pcBU+U1J9fizsdurWP9t1N21KhfeM3sNIgo1e6
822hqw1mDMWqKALq9dY3BicvCdzFytJdVYosFpomgwF27OwWnbeiNOUnLXbq
XPD14IiMqveGt8zzzbZAu1RqyljuWhazYMSz9ZC+K62nuSlvWTNdXiVfM4Ea
4dPT0eaEzs+nsrqW6/y5mnxX4V2NRWpv+tAGRThqHl6rPXgB/RVTXDiF6BTh
tlsUadqEgEyMPwZp/Qtp+v5m/XwP5x/lv0eQtfGuM4oVdRrLtFipAlmKiKCb
8ZY2X8LS1ugVYOQFo76NtwfAD7KYXeBvIlKsFlSs5qXkochQK5xvAkqAyqo4
YJCU0Y99CC5TOljIODi8Z00dPYSeCskx4Y/PePv6PdMmnUTR31sXJ601mTAv
BYm68kWnjQ+ZXKS7DNJ++Dd37iBS98izaz2YFfaNFQMQY/4/HYQpi+SPqJdV
AXAJ7fuMfYXKfMShYABXqXpiAym/QB7xijKkRUHIF3b+zXYDldyqSj5h4359
hFK4voCkOXCqZf8N3ypnKfYhBaR8RNUa+BC9tGLAHmU9BzuP56nBv0XLEdtP
Zy0CDxM+tZmR/d4wbXCkEkbfzAJ4nplE/mVhSSA5F5YoCseXNQsAGb3Hu+JX
xPTUR/eR3sjKN0k/UTLjA3tu7C+Nf28CHJR0+ATYDjl3C/JjaSVJkrxJlMvd
8mAsTaaW5yM+wyGJF3at7cnR1vGONUQbB3ZcXmXv6T9KN7bbtO1j+7qTjR5r
6wKGYltpuqqLjk9kgLQKxmNjRRx2bajQYauBfhfoD0phOIzr7h++gc7Lumhq
ZViwh0awGPb2WBrFO0W0iElNzDO3DtkwGsZ7iFvryariD7b8GEvE9Fs8S/lb
l+oo6xGF7OP9lpMiHlg81Se933PAjZnfGB84lDyn6P9je2IcFdUS0lD2+vBZ
uuQmq6WbaZxB6ZegHPpP/8OqgYJvP1hKSR7qJ9yMWSsah0a5Gslb/FFqdC2A
3/VktpSSdCNNZ16Z4PR3hYXS9eOX2fra6cLZUitSZww4mBur9iONAl4VuafB
myX1zRoH2clhYowGdVodt+YSXtqryBPDL2i/ynZnLY1L7j7ml6oLxraKSZ4J
V+sIsAgbGncaAN/SIW45i6XKv8gXH/aMrnDR975crz76Bq47tR9xbCsapA5/
hsFIyq8ZcM7SuC5D2DA4HU9zWb6OueI/N/+d747mwFV740PTTbUlAAuTzz+C
ReRaj/S1WNiRY8MRP1Az35fjvB/PwBr2V0V1abP3M28l1ky6gfzCbzghpQds
H3me8xvHjTKghznVt3i7lnxtfRR0T1DBUSpSsCdASp9v1yd2YftanIWGxPCN
DtPczaeOP2kVWegJlYxJ8niT6r3FWHUi2ulRMgEvo+K4rRM1s2SYlS5u8JoF
LGD3lcijEU8/xr4zDNGndAhqqElGTd6GWkaFIy59RWyGoRAD+w7/c+vuc5UF
9Q7JC8FWmaE6QKMuMgSuFbJUO5B+KcEwSGkCIBkgk3J3RJS3qNG0dP/bCYTD
ugMVrDDk/4RSjg8XUS7mBO//lXOZMMwMueCWnvQsAo97N3FtQas2uQchDHD5
TMFUHA9bK6ws8blXb9uNY6AiUiLfOmk4DDtB/kJmrYzaFMRMXSzvypdRgnGJ
qE0nFEclE5r7cgGqFi3U5+gW84BqC+Y3n+DU2OLiEdWRF23+Rsz/P/X8hhgh
VzhgHF8DIY1CXtQPKKyzNIc54bRDn5xZt8ULerROKQQcvjhvBZU2zBw/17Qa
gdYVeVsozHLzLbTWDas4PI6x2Of4iG7aJ3ZsRKJ5NJ7AH0u6SxHW509o/Bhk
L3OV5yAYzFMVtkY6HisC0YAgI6XfAhNaqzF7gzeph5dlRzt8t3XIrv7MdgDm
N6GBAuj14Kf+byskvosEn0LAgq66xwmtPkYWwD3YujnsG4akxKP8qfhR3r9w
4Yy901yb2gYhSNrpKvdnDta4Uh+G2b2IHwcBn5Pd8S0WwWguPxvgRoV7jm/G
1QrUO2q6z4AJOb9ArPZLLCnAUCk8ZiPVP79Tz7dYBZmL2LVPkps725TXQKBb
1oMDp0yUM/Jw+AP+qdPKjJeskDCxfiD4Cc+YmhRbx4UpXcw9ALwZnBcr0nWn
7/LBFOO1M+lcdIXdYR3yjlOUciED4UX747yDocORRniXFyPLAfUkk9pBCSgS
TH4b+dMDJuarDWAbN7Hm4PnAkdCQxM89tP4NMfZ/wi4vaMeO/FvtAwqrHt5m
qK9ZjlWelHZVtLugWWoW4OOEugyaAcqDLmMpEnsJfi7Iv0+GqL0ZhvsqGVuj
0RN2Sk61lwdZL0JClsIyjBvYeEKblMwFaDe+cLTvruHd+UDBGmGT7aOIJnNE
PvStAAoqN2D/B/zm/IxHOk4gKjLjtjVG055ad2rmdVAJhYuhHRntqTyBhPC5
W7cP5ggk9XCg3Ddct8d4vTFEylD+B5p0ZbUjpHEtvQ3pLLNHPHFEVRqNGZec
ALCWvwfjHZfJ7ki63cWOWGNS51qQ2PGWzsO8XWUokTzjg5VV5mrOyY8fZgY1
nbL7S+n6H29Edp+tG9Au+W3jLePK5LcBTqwL+ndKHqKRjuFmhECf3T9hyBqx
LnK2PlY9MMNy7VnemKkF+HznaZ5JN40INvj/xq5GJ9Yczw95Dun22HBtc8+7
2NeMMHCDTHDYH/8GCXOPIeQOuEjlzBB3/9qgPtXDXINpDdVp25uohyRgYdrI
N/yiu+TIi08NGTmCAGGc8/ejGh8o+vaxjGn/MjQqtJXmUcmj/yDLzDBuCXwR
ekVKEajWTVTbEFaJUEqJ2C14KTwIr566JZtT/4hauSZkJhLsAm9tbiRxxx0V
HLR6uy+SWZM11YgJ+FQyvgM/KXDCgCLhA4kdJM98lz8BXKKXdYuHwV7BfGHU
HSvSQ+/jik2CI5jlCV+jb2TobdkokBpJUMfg1JsrvEPt4N+FeWtvwd4hRJe5
RayaZQCQpLlEXzLhbPDYg4+Vx2L7uIwNcIrLDLKKAU57yuKJbgNnS29B1vNH
0baz9w8ATAlhYLfRCwm+BulyZqbcH7ps3jLbE7IXg89qHHIOwAWL8prXi3Y7
P7+J6u387Z3k4kIsQTB4lBjW8D4+ZFE8TEprY2LVF3vsZU6Y6E6iCyzzb1q1
OptmHTi2Vu7RX0f3BjsYb87bpQEaM4RvQ+skBu6PitxciONfzT3SOc2x88/D
IfNecPS65FG6I64E32W0XnKsf6rniDXJFUndOVUpF3P4fntTLsI7LUe4T2qD
/eELg5Ugh+NpuDBlDozj56gZ/WdQvR+TEBYvBElijj6HS7mEmkW+hevF5WGu
ztifjdzeMLwJNFLwHteLmHQqLFldXi37y9b7t0MIRmFPY3yvY6QQdUKFipou
i3k7U95VUu5aUboWu1qseaxvwrNX7mySzbFB2KHZPJ6Z1Z93+wsqQC+ZKS69
u8OmA7wUHvx+U8qiO86cc6pWUA7fqNgxu4865UUGGUEXlfUBlRMDFO7hc3Jc
0whnde0Z+uIALiPI88velEwEJxF69shghEHXkRF6BbFCD6kvElyBbkwbHSOB
nzJ5LUc4t1ca/3sVmm3mB3INr25fuHi1l/ovWfWuYlcYNZkn7FOfn2hnfvkJ
Z0mhnTTbYMRfGFc4jKeVovGjDdx017dVAGuddEFuJy/Ty4ivG2IiDVK/CjPO
x1meJzYWJzod8g/zbV32SwgiwFUM0blSgaymjl6wn/O4AaVy4M3Zs+2ahusR
E80XgSaPAwKLV9I0CNg0+jgqaQCjLugzMW+8k90Z9C7PffXjesX0NEoNC+yq
fnpzClyYFr+WlLL99U/jWL10PegenNI+6/v5YyZk0rECKniSdzD2rJ/pY2Sf
xWEMfl2eyaJ8tHlvh1aAcn5jAogIJVbaQOiXFdwmZeavY0NIEWAinTjWDMNL
IbOJS7HlUkJQI4mNJgbYT/Nj30ZtmzSmPYMdt2jM/oR2NyTV1HDci2WmLlwe
H2HTpBfy3R9+IaX/rj25GMslJSyhiI/dLdmQKa0PYGSRTk+MvoE8kjfdKHRO
y9+i62pUOsinbEZaUCgG8Ww9EwSvKR7DVVXAxCRNsmni1+ipaGFTzJX1HYRu
K6JRG3vYwYeXF8seilwHlhsEw7MmhrXRUE78ishT8xitvhDW+CrmpJD5Iaf3
Yk8t+QpBWEv9SnAvyzyW5F2wcCqt2q7qyiNOmunDrLu/ZP3xBmkybF1/3cJl
iyu4rKe2PjFvk6HAjPmJWhWgnPilx6gxdpsaRbKruXOV/cSGx5VDpaYom5Ib
DH3YSrSaa/uxBoejQYp0E5NH6ygmC1czjw7uwfLa6aVjDUGJ45jb6sEKwvm7
xz9WA674rHVfLEBJ0Z/u17SEK/7I7wvKWrs9iEo7SBoXJDC5yc3T4eRLBYZE
RX2KJYKvtQ9e4H0rACmsR1QYdzNrx8IPhUawrpuiRs4lN16P3YoOaLZEzXe+
DlQw/tmpWQnO71KmJHUTxwScqJfCMaBFoiVvNUMxx3IU9isJs3D268g51NHn
lBD4N8RQ4IHV26s+kOsz5SVvZA1gkENQDd+zFcZPPE5oJZuTdigr7v50nsP4
eOlHQ7apA+UQGc1Tn3SDIQy9Nfh8C8fc973KxJwjjMX7q9SIqoacoZqrUr6R
1O7KqHTqpDK7aNY/eV97QqsFXLE7796CDVSqztx9BvHmIXx+7t5Kq92cAINb
O2+DZJyojSHOCF8zaRu4YPXcroTA4YZBd4sbFN4gbvxaot1P3NhSj8X6W5Gm
PuP03vPay3CLnJvKLXl81xo3kTw39OS3dXiSP5qIyNF4tP8dDMNlQs19s1Sw
MMofIIiUNy8vTSG98hyn0l3BIBMYorUlrqWBfaat0m1xZGNtQcxssZ1AOZ0T
kG1CZp7EYyFyq+g4bn73gkjg14qSUokZNW0/H1OFtPkCE4Yu8SllmPXJ9VzC
WFTPdb3FGL/XH6NEW+93jgrQ0zC041O6nHr55HEG46YW0rfq25LSGC05ZVW/
qBHtos5SZHf0FstMY5e2psGOdivNLDsLTiWqTO8ftlZaUvNc4UebH1+55wFG
kTbwvop4gdDbHgPW1d/MrRYNZl9XMULkTUewi1YxkdC/Q33M9lwvYHyJSoZV
QSYsJ2ysZPJUPlCB1PilvWXaNPqKFsiUt5uzPG0cRphIS2tRu6WJJgy/Dd39
qa30VU3jmP2QZt0/AekCSXnkABE/fSuM9QOQ0nc/pZY/H0D3yM+R1buikjui
YEnzokAydEQx3/IOLhyiMpZGarLWDGWUQcLa1IJlNYylANS0350cKfDjhcRR
M1JcrUgXNDsA1WkyVTRma8talr7AtDYtkoDnBFMIdcR0hitlRTCgU7uVCTYb
E3ZhCt1abr276euMlCB298iIs2UcrPMwvdcWqFyR9/w3z+8rkXVCnYV84SQP
BVFF9pxKfSIG1yZ2co720z9Hk1YXqiPj56Mp3WbzLYFPKDyEzktHq1aKs/ym
H27vIBPrbjl66P9nkUJbtxVFZIdJhKLX6BRjb33EUeYn+pMhxSO0naHuWohI
juiV96yQGplB83kt+iz51lkKOoNLN43NNXZzKRP9oYwR/1HcJY/Hk2ngV70P
cINPryaSY9pSB5/N0QR0fqZnV/6jmq2telOuEt6Htv0OaglZUUq+My4SgzH3
N1zYBAqL7D+8dL8SaVJbeAAbWynEB0n0Q4Lab46Tn5YQJCXHZvKiNfXlhcAQ
VansGGfT05v6X3LSkQAk6ug0ddK4UjNNb45cVSdbBRMCOkXpG8kYsmK8Qpud
pMOvvrvDApdMyc9MoDGdP8MJKKJTAueownW+jNLx7bCOIgEBoYw+NNCjFTg2
6Ad12qPXSJNa+E3CknizA7vkqatC5NCvBBLY4zcWG3lhuVKwA9DjFqn2Fvkw
vuq8P3Cxs2og/TKrFxv4YB8Ic3X6dQw+n8QSX6hORnskoQCzoc5PPpBUOMYc
ZVccR0cJno1Mbm005Zq5ZX0HqlpUaqEVgAbmMpy9jJ8bGrASRjtNE4Qymq5z
zIvDzelzUnANT9Lcm6WkdF3MsxALS+qBjt9X9umBYP5Aut1827mwoPsrbEEj
99Njal1JTP+zWhkYjStqT6xf12ETvqBgLPyVNwUqpMZSwDzVh3r6AXnO4ean
VxwIwjVP0DC4hi9/4NBNcpiZt8pb9SV4tKXzFXUMsyV+TyhnmQGcvR86ld/0
oyI5OXuItTDGEXl7a4bIyw07f7yIpq4Y+mvw0pdcqJaykomVeIYcAenr4i5p
HOySxZbjXXl/O0k8cFeVplx1ZEcfd1/7p9ygkTcZPGlJkSsI0sOa2KjNRR8C
f6MzjU4q/QkFvRG2gP923I51DYjkLsSSgngm9Us/JEb1oDB07iR12eLjlA2Z
M1zWA0WipNFrT5RfSXedVBzJIS1/LcngqWirQ2it84Tz+dy9lD4HhFs+JTAU
5C/GRBezNdBh3+ia8apGaAUgswPStuwqzLST9h8JUqou/8L6J2OUtoZdE7qG
LhE1HMFPPbkvI+IDbafegXfsFIXCZkdSchR+xIzvPcOqH0JxAA9Y4SzrM8V9
rrK/qm/z0MYjrK723/gfR4bh2MRdvG23G7NNi2bd6zCYn/qONX5gU9TP/nxn
Ej9WzQegxC3nro8hOBOd1ID4UhePNApZL9gyiY0407S3jS0JjEaGYi6q3M+p
UUNPjMxFe/ywgP6icU/XS7H/EaK1iKWlFKfBWNbNaDzxz+NrnSkQmEONHvJZ
qXgYdY7mzeESgqEfKsJR84gYDDPdeK+56O0rGaIOtCWJyTAqgA+N6+Mgxgq0
TlBgEDUyhT+u62QyiPiXboa40sgWMDK8KFJkU4oO3rQeQ2GD/O5/Xj0noKri
WD8ktBiw47sFV8RTjlDqAflMyeb9nmTaL5wLvlW7B8JkQG+nhFFzU+oaIhxz
sCljwPFLIfDLoB1+zOJAbhiddAqR5G0lH3Swbkg27XX0kBWEopehAM6Ij1KN
1JPDFkeQ/it7QfulKLcRGC7EqogjLa2u8wmnRbFFZGsolI0MZksz5ZPi9koF
sWlMfgDlJgHiKXJuAGzExBVu3Mw9XDnFZVDEs+Y8Ghme2n86QtHe5blliQpT
SQnnTQpQpUu9iALz5m5QqE5vZS1ke3IsQX5vSK2JPXRj7szkURWhU/ESI5qZ
YjdxYrbvhCIMftyu/l5IWalT/zdQbJHFmAq/s9heWeL5bL3bxKwSKBRbckc5
DQhd1GU/MMDr+r5f1wA+KOea/B2nTscgc41qJHIGyxMDYqmEQI6GbrCnfCap
xtIjOY+V6ZI/6IBy2tlG3c3YUD83f9AmfCpMVGOz5H3aFvTFZjSum49Bcuu4
tdOki7nSrKL1RxoTdogxq5TWxfkqvuDyp6rMgfKQiOhmRBVbPWdW5fPwq1rd
L0O+V+13ZCmnQOYwLraw24GAzon4taTI3EQqavDZSBaPelrTaKkgKBhOYGwQ
TS0mMAFlURRxxSvKYClaxBmYbRJmZwc62Y3Z5eURpeH2SgHrin3HF24BP6Xn
hgxwkuur7utukzix7IjrfW9kDD4AXYxCJvPUcZuGycMtsUKGiibU+1iqO1/N
ymY+rNEwJ4uWs142kVQDpBFnCxrvYXuRBb0bVnsohUO0XUnjWF/FyG602u76
IBftrT3l7XEzGHwO8c6eRZkSInEiaHdGD0Gcd+9R/mKP/PuaU0PGLKSY1ejv
gwkNBT72jt7wDplKdHZVscAN3dOQYQodix692nZaPSrdJRK41QIz9hO7V83a
lM2TDQbsBdWkeOBHUjWdEWPHi3W2CMy57mPwVnWhrpriV4Qp/uA1N9Krxi74
f/p/PYa/IFMkoECKy+/zj+sRy5az1fdHjVSVnBD2Y2I34v0gzo/iu8d82KFr
bfXTpJ8d9hJHjnTW+8fQJOqWkBFKv1L3/Mlu7oI6Acgw9+2aRKjFMkELLs1u
VKPFFUpd+x0rxdLUsNDFiy8lL6HiRqGFF+CSSyibi7fnAJoaYctFgQmqH5vi
LUOr3qCvqQDH7ZzZcW9f5j1vn0tuxYo53MSwb5/aCHvTx9MrvM/74OUHuCRp
yBGMERCOc0tyn4K2Z4dKFpP7S9itYpIy4j6NPHH6iO5WzzPqb6DfkXPgdzRg
2EOYIzx1WXuK7OqH6NZEj82ts5yAtl9CvPSX70Ha0w7g4bVEH2lveXRzp0bh
DwTZxaiqeTbHX77JoLy0tKCwqFcjNrMuDVkwxe3cOsyiyq9PPhX2xTsfnslj
0yIG1sjFst/47HtfDTrubP3kUbfM03LguIxzOoKrf3O1Oxc+RWsBYMtllphY
4N7Qon/PhY9GpYubJn+Wgw3GK3dAq37zEROmDwdVgWbddzPdNXEwdtrwmAK4
3b2jrFQ8KwRcWNgklKifhRYvBdoW5+4W0RyRUGmvMKj1Jcieb4KCfMihjHGy
PEKE4hEcwZ4IXmcV65XpOAwB3H+7Ts7ArGjF+t7DYh8nllCrzEbmcdJLsYgU
nXtRlH9uEqEOumrgq439DZtKD6hF7uS6i2E2feNKkOnKl6tUuxjBECark4Yr
t1CGsfl55RAEdT5QSL0yBgItx6R2q4LKRTZdLLpF1JVPKkiVtMkeo+LaISHs
PsZDXLxoLvL1A3D0xlRhxrgM3bBgFyagNusruoCcUA9EYmJ0KRg5Yaf6aZ+3
vmRGYEFGmD4KPI8/QckEIQFo0ucZuzBNDg3lU6mz6CXrztrIIQjfuaLTllv3
KkaF0Pne/nhOukLQ31lbFGqCKpNzxe0GJ14HLLXsr80V7FnDDCgCQ4680OPq
5xughhzOKu6eejGADtkuuC2Ec+pwmbIvbT3KZJCfpJW5ZKeFbUcS2S3cRmHz
urdJJGwMHZh393DJIrH4n3R0jqg1Ufk9nSc76vKTWoy9juUlT7iErmjTsoHQ
o71bgYvgY2CBT8J1tplaz0KZgKr302I8TRVPPITv4eCO55bsHkspek/OZOOt
yRKkg5ECWK0V08FJE1y48xYDLeMURX6fhgN8DL2ffChqHJoukGQCFKxQoflA
z4dKFvcgJHTWKH1W8YhPVvGRLLLpRFKMIuZxjSeBmIOJy73vGtwvMOc8y22Y
EiJ3nK3/bIgu1Vn03srY1FvTXnMdi7eFtNGzHJD7saEw7cHQrsO6xwPyTc59
nb3cSFFfQ37PDUcGwUNudwhXtISXNusm5X1GsEO3wzICzKuSfVV/GfgXjxm7
X7R2maRKLQDsfscNrFTKfU/737RGi/rHW86oWCKErE9NBZwhjNXdeRxaPtt2
Beq1VmiyFiSm6ktqgoN+aMVtNrOYBdwR3w3jG5Zh7bwwVKs3iEl98QBf1Y63
6ofnBatZqvUeiLRY6+ndoMNlcVxnv4YaNep37iKsc36JsMJRkiFJDNBDtDRl
H83amQ4XaI0TXlueQnLpQph/poVZUrB7LELT/YE0vCR/vphppsfwCvsiFfYD
ypgb8HmlYqYsuhCzw/Nmzjo1OrOlOabQtuVDur93Txnm0sHQfxYmEj+4EwPu
8K6uNf4j9aEtC71xS9ZP9XL8yLBOxfXcjwjDEM9iAFRaB/hWc1rbdCPgqjzL
75vM0VL2JoZZHx23loscZkmb6JKiCclM8OrGSbeunIFeCpA7NyPyk9LAsBWu
tKAaV8T5GKBsqyfz1wwrNOj4hx0VD6kVO8rSAJ3Xyaj57Eqy2YG6cwNcDWQH
y9TnOVbQYBFj09XeWjpin4EIck7/cM9xIpobF4PxgHIqZPk4w9ETntyfP7n6
WKLnEwE4vjINrDhIGM2MBrg5GHTrqnE/8XpLa4J6eh1F91i6/Fj57tqAN+1q
Ut7RGxN6ORpPpr7kr+XwRonca0XpD2/+50bfKPn6kgkf/BbZNjRp2fiAMY9p
czqMVOXjVlGiJqEG+kpvr0yY8JydTKUWFdy4ZqByrD8Q2n4Lh7Uw3ebJhdLR
FFZcHlV25ScUO/1TzjHw7r6pIsG86h70Iu/O4e6FdOgRq/cdeYCp/R9VeDSH
G74u1/OoD85ctkKtVg1g0MLsGeTb7N/ynPJpJ7M1GEVLgQXwRCAwd/geOrge
lcm2DxU427YosNNR/dJwXgtPc0hTL+77iAAGVXAm2NG6aQXQ6Ba7oUNKMs4I
BMqs+14+NBS/xcRHs3knqRaLsLK7HJaiGWRlq+9htjczsDhbi99KenWEDiyY
w7zK29L36AI3PtINr4UDWRzqYFud19Tu6BoaUmX4qcLtuqromfyQ4VCLfhkD
2SqXYIsu8Auk4Wlv4K9Oxathyz9icSDC/fTAF8yLqA6Y4ddWWuvzcWsUei0v
ZiJG/8gGoVl7zjMNXT7W0WD2aJAKu9rC5Hx6dWPclBbt5oXCT/57EL9s4seP
O8rW3FsMPsvNPkp9FGmZbUIgQGubbh6ZUSObrY43VWltrp+VtDZ5010yRtK0
1/DX5iYxu+MO489aAFLlFdIwoVuodnTu+dpcmjykDYP6+XbIMMr1KkdeIH8r
hXyKhkF/rsvg/6WXEmqHiUJbUXCOHLwRtEjdSayaYLAcuexcWfB7Ifm1+q3d
mTy4BP2nVw9UmwuRbJGJosYICI8PJLwH3D7vIhYXTBblM78kzPg1/b9O1BRy
yswd4UrsvN3HLeIsOjVZAbZ9uAafGuf+YzNCA2AW/eez7EfUreyyCNtb4V6K
a6yjWSFiXZjDX0aj9p3iwm7fs2lE0zENPWEmNk2NO5VvTxkf4EzEWCklPdkJ
Ph+lSloYbFByYRStjxI4/XFI0O69gkhe/ewBVxiWpldfecVtHcKfUKOXZ1xu
TLJEZ4+/pgNRAuSaZGOy6U+AJqSwEg/LCxTwVrT4W38dvNweX/7BcckYYXwn
xfKwXy0PjcWoXi7an6I0vmUf1MJzIEw7cUdKt1Gj77HsbjiNVLXFQQByREGd
sGGNa1BM3hW6tc86H7N6Bd9dES2a3w4uQe0pFEgzOcknzV7KwPjPm5LwDLLp
HIyrmLteJJExI+Mef573KxsarbrZUWJHx/rXql3JAlYJVTGm4l0+aoB6u0HA
ZHe/mOTKzg43AW+o9cA5wa+5NZ9dmHjh5Ul+4v46H0W03E5gQSYQrTC/stSi
woTfDtdm2TjjEX0XktQeegmS0gEAiWiwUuxRXC1vqz/D3S8Rs9kuxD/rsXs5
WqNc0PF9JTNCXs4RYS13wEpHI6qY3PvWlHdnvAKH7pIwI1nUajRiBZnCvSvO
47HMl9SzqdMhlPb/RhYPWyFmxV+cwXRHDYxFn5TGcRh2UTOIE/HQn8tApEdA
QeFM/3+4TtP7JmT+JBAMIzdYoRPSCOhOVAGD4+eNRjwz6EWx2PQuu0zWH2+Q
CvVVaVDIgw4eC1QBVqeaiYeHD3f3kXCCAAcYDm8IDfB7gsv/z0ozpATk5Xq5
UGUbAlP85Pa9jzvSSqv4Za/ThMF7kDz+mMzO5rWbStl/rDRFHXQfs3UAU1T6
99oqEJ1PRFb963ksa0MymcG3hzuS/70TR3pvNWwoeGzOYtJ7wU/QKO9nNeD+
iay22Egb+FfshzeknH2dkr4akycKu2KciwQ9xfWcHchjrKQ87DxTBYd6epsv
+J+CM+2NgtAYtF1s/omQvWAfq5TSqYlebofBuy2RiKCgsseohn3e2051B9j7
O9DsL8UwI1DI1HqY+cSrm1C1hyF4NDFi3F574m6CE8nUonMr6nAiARAthF5q
rXCkNnM79AxCLaQbOumB57aSfv8KhwhHeSI+6zRIZegIg05VwnTvL68bxDtr
i4xMpy2LS8gjyEQYXBWOns4dlxMsMFHlwU6VDjl/t5k/4hsffbswGmm9ZVWM
uHsJ/PIH6MeEmv+IPcSs44G+lf69yGEZSQ3/SVPmdIQmfbrymyPNG93tLZSD
MvnbvUknBPDSmgfxh3a9JqlQMbH4rST8avd9XZPCDS9ibooMXBqlsbvteJC4
ZKSIT6OrjrG+oVk8vFBmCSoTwApHovZi/9GG50NbNnPn/2HjSEoseWnX+i5c
9z+DIDsMS0MhwTQ3YtZP+gBbpkEPfdeq0F6i9dVO9+lzrvayW7x9l/jMsNGp
bjIFSNv+JC8L8iSZu+8xmICkV020Q4Gc1pu/Y1mpMQUgLwIQ+fGuUYmkf1C/
EYTrKkBDCASEL6hNmWWIdpEdXGAcTZtJvkbxbuwz25qK7uMeSXPKqhf0q63V
EXvpXXwmLO/TyTRcHnq4xRjG7cCQLIrZSuQgDaTgDuESDFksCo+k/Obe7MZy
U9yTHsfIpaxu4GEaZILhZaDgvqw6swZwOBQUuENrfZxnMC5lk3c9PRPSuwdw
dzz0xvZyySRGfOoLxdbPnJM3+301EgNS7USXoPmq9V3hwHlqnOI0QNsVzR4T
ittams0EPRTK5U1ShRVtniPX8bKrUh+tkRHrRELBq/Ybr0QAHvsr2Sbz2dYt
D2t0Yfe6oCOkXqWi+lGfQ57WRHsP/7ekjwnLODYNzh64sfVyQpMA4GS/4z04
a7GDdSnuDtmKkgbm1SQCKg7y11TTXY91RC05MJyUrTIbZlITSC9xONlnILGm
HGBtC25gMqEfmxyOndZx11TVp9lJNqyGs6HBThPDoaeEr/z2dD1BEYvZIYce
f9ypPIR8Lusl/0ryYtsvvaYbx+lriS0+vDpxUurnd8/OPz6UNQrdGFGu6fWr
pm339VhB9yIUHrTa5rflr3Hbs+4EE5fdLS420KiAHMomaGTrZkhlxt1S35qD
71fDp9/aPeLRWfVLlldb78A/qCCpCXfR+vOlIVdOSjEkM+sT2oiW0AEBvBVP
avv5OPszF1mQJ8Gq/DhEInZHNlVBv9cYLByKnVHo9qs+Pvc+R/KUDTCKhzmf
tRaLGzh69HPOAEn4Wci7dxYDO1MjIE8pY8Htb4mYpRU9BL/Dg5BtF5HEpP7B
DqobBQsPRrb0sdpKD7/gYf45nlGL3kt1d8iCNUw2gp3rMz4lMm1HlW0ifI25
ErLbx+V/qTtzzwLAqYD2WvOENdWwQ2HGqyyzlQeAplPi8UQQpfnq5uVPDvE2
ZGrdEkcNHR40V7x2ww0uXy8DeVAYZel3+zTRMk/3oA6HeQwW5oc17GKkpj3u
AyXVZeLdA9Xryl+RbQWfniVvGztFbUxHhTPszo3OEVK5/XlAqTLULCKG1A9I
V8xqHkrL8QSuq4VcA5B0FWWTXRy0ZOXW0B0fUhgf01xYzmeE4+WOqCfpfJpo
nhMRqc84fp73hJw1FNna2dW/MOhrKYVRRCHAhlOXsJxHQzBjj+IJgm7ymkG6
sPkLC/zqradcTAC/oyxnYbVadSvvb6bZpo4HnmU1j/yBXS+srxRzXHdq8zTF
8fozUYvQlC9CxO/EOMnws4FRqqN1zqa5oC22x1/oVsWmz9UYJ/o/YEHlG/pF
R9d3w0L5v0faUK/+9sApd4Nlm2QwgnZXQI71O9E05VmJelrq2/tMLYAOCo5P
gtCcA74HV9DFNs3geKTjQw8F29wgmT+6I4+cNbWyj9Mf3bDjQslFUd7HSL/K
CLf2v+Hgs/WQY4LMV3veTA2i7KFoaeLra6yhPysLnrsrZtmh6+2KE77sYrsp
GlPpI6HCoA0T1rYeSHX7dHJpAVqZQMR1NAHItx4E3xV6TEznIY9AtBU8G99/
VRNinn/qHmQ+277wPIk9E0qnjpOtcdMNvYjkd4drfM2RT+Iub59CifC+fJad
6rLGvlVxQrRdmqdl/xdzhk7y97NjnOvOu2/7bQPxjdS33nFKDmqpYykD4lIZ
yGINEgf4KXiXtsAnQPFrR2gbBJzMoKH/vdi+zoTFDmzQAoYIPQbxh/YCuHWT
AIQ38BpbGV2FN2JkjF4chANGqKRvxe1kYNn9w6R1NjJzmlNYzqkU60DzCypy
dqTl4uSErYXjRpmyqDSm1UJNA0ACikAsopQPve5l1qD/fWIkllSkVWSSpSXC
NaBJy5P03h0e7fR69KHFxd7I7aSC8IwN8EGKSTcWhiWzp9lDjPJ5uC4SEXyr
tP4MBn+FYyt0CWe4DVKnVZQ55F32tedohXCN7JjDL/c5xGHTS/ViGo3MKiVX
4hGnfBRdTmDKXDcni88J44o2+Gndd0oszLDsWwHUc1/bac4fzt3jLknpWm54
p1iwZGzcwdQLrbSp5JWOXjJc/cSa78t3YWqk4yxUS+kmYs2QRoetowLV57Gy
Z/QuMckC4XYKR4r/3dMBvqBon9SDT4z0AEYC/EXoq9nLJ4ZjRbfkjFLWnncl
00JpELQqzU1lx3kTRoCQWkdiY3wWbbem+NCFAKI/U4p5uNfh1Go4XO+5B+sh
/RSsD0xdPOcmDV0/iefYZgWOZTRnu7CB7DkfnLs2vPVL5Vr6NuR2nAOF87QR
xB071bCeL9v8wF6dvZiSjNfecXUaZTyLm/GKiBy6A1k2koRUyEeMNbmTT6K5
7Bf6sufbh8+iSawPpeNuy9C5JapG2LkyFPwNt5xLCHk/F03y/M+Yu7s/cJYQ
y+TMdAPsX1Lwn/qAJN4Sa+m77HmK+q++Mz8MYIxw81C9RROdJETRylHb4QHC
dbvbt00m8eHETP5jaki46HPjt6sG5YlDt6oxQTqsXTvGbvRDD3gGI5v38k/u
rpJYdkXkSOcZaFnTjlSq4Si3s1iTvVfjudrIJGCkICwV04e9Y7UdPa6THvPa
fB+Sa8H12uqZINT2nzvo0vF3wswPnOqqMf30gaMtAZlYGDTWLqyvxzwMd2eP
nZIA8Nhn8kx9vIMwMNjkcfU/YMdwOalPm9yDqyY04YfkShizopht/qjoqXbt
iHK5QoRnkZFQOppTmzU8kBhoWbE5dfnkkZBlD4nJrqQtdZNHrFq42nOYDIgw
knMhcBrfLQu7zpyFNKCHW7PLWS/jfTBICvEVqkoeKy46hd1TTplSDO9KDjko
6Nn+61gNYMApy5nHtNT9XZ3iVxxomWgix9je/6B16ArMFCBmbl2zwCnpORcr
8jSfC0FK2izA785CQSUyixxfBa7O14rD4rERE/nhEC3r6FT5+ila1UWZDXk5
JyRTnx2AuAzNqsndcH0RwTWWZPUjtPObomMaMNrMUXrwoWuaVybDFKU9IjUn
rM27RowoO3mp4v4x4XCStJe9lO4MvyRBzsHbvr/1PBRkZMmWBEf2v5Jg2Yq8
Dhgdrrad3w2iuk5HOsuBw4ZG4z4U9eoLZCJpAgwrAnteOEssfK5uqogRq236
FTY8wc8oKlDSRVaYIF2b+6NfVHZIEEjKHM1+8V6nZKMkFqIGsAh5PndVuG67
PP1KS7GXHkJGj6FlE9csolepTs/3bXys9+Q5YzBMPYamA/nhXPy+rEMsdUVy
KTQu46qjJt+U+fGEWgLAZsDPB7dRYo2Ssvr3lyWGqyUprK5H9cLUhgB8iRaJ
bR3jg8+ejUJvRwGND5H5RCLsJhsA16B7ovLj2/O0qvHwWB1+GecXuR+SpUnb
NBWQwC8fSKsm5CQIaMfBmhpg7QU4b0FnT5s0kSBV6qW9UIJAp/U7t7d1gZMU
/YvvaQ0mUE+pIYp1Bd3etTmM6qlG+yAbTxwc5dZK0QkKSBMwFink1bbRcZ1M
+30etN//kdtZiQKewmUHUVIsc1V0WB0bvfvWHXhFUFwsXLbhCQhmPkujBX/I
h7vTm6LIauVEj1fcz02l/7l+SWwr62QHSwpyN/1cFC8kDXiwV5KIfXSUg94F
WrHB7GpkWiNRK+HQlleWigKFB3O+4eB63oZZfQMy6S0vqjxa+hMQZIkIkDOA
EDoHYej3nvVLePaTrXMqtkSQjKTY30lugWb9vJ3e2Od3mPekWkkFEY1cH8KN
lagM/yfSZuWKb5cJDl8h6EGh7R2j7YbwS4fFqnLYgPE6nHU/wjthNFag6YZK
01GAkLSzSXTs6YcheaD+zfSIaW+dun8ERAoMDKoigXX/JWEBWPNiZygQiDeL
5h16wdyALMIpXHiy+Nt+R6wAKOY2hTQBcKGwhzycMTjoHMQ0nr6L4mhcOEcg
WFEJGJGT3HKNjFDHzBaWqmHR9RWlwrRQdIvW5Cwg00yrGYsNZVyqx8OZ2og6
E/IC1qAC6+Cwm0toAdeugXMI0npZdDRDgMiX6AHPgUYdA1BQeJPiV8SN2zMQ
QmKdJXmaBuehSAZxXXzalDEVtc1iimtNf+9PXlpCZ5ljCGcihKiRNRKTWhzO
u7VYFrmx4jERsDx/zYyIrjgM2zUOYRvKl3RJor/WGnIlQ9adk4bRB974hZ+f
qDs97JjrulMmhH2cNY6NgtrhsXbHIRD4nGZQIFPC1K98gQbnhbLRcpu6qCnI
CSVepJx/XtnIeHWuij8AGPZJX8tCUT+5XeQtSjQ/3XbK1ve2G7Bl/9dBhuM2
p/SvJ+Qpw9Me4OEBLxFL78x0R9t6ObDuxnO8/cJ2WER3kS3SGlfDPcih9ZVZ
Getc+mFxTRoyNAj0U3gTU/v8fhSV9puwsSgpz8IQhaQGiFdGKYrm7vlHn9zI
ULOse+2elYgnVAVABKFaqsgCZJf63uAIOXaimfb6i3WSYjm9fLebEDxbYp3X
JzWT9kOSZcrnZ0T0gSY3H03iC5t1cGdkH4AowzHGKGc+lokW8sM1FiazBZBt
QiC6tHl2DrHtZOrsTZhEx072r0kRSNauJfCLt5qCdPGSXkLm7/AXpUOv7iea
X/ebli06Bv9YB+tRceVcTDp8mXPF0Ne5WZmeBfiNVsJupfUj/ZYiVWWQIfrs
eqEi2sGvGPeQQomArC316CQz7OAMhnctJ7G07vcnz0WOAltgl2/PX+XzXE/c
DuZ+dYHW3nDT/lfjpEIfNrvRtBwuAjpmh0r77ipLv7us0zR75+HjIQMPbkZD
qwFuMhfr02/DU/HtUbnYtgrSsFqqDhewfQiU8J6ieW3YJTI/CFR1+Ujc9YgI
pIoyrqCwmrrYCkiz+qHbpi/mNVQG58T4j/QgXQspUHI5JcMp3ilQxA52ggQD
6HX9nzPDye4JIBZij3vuweghzFMKbIrdCL+CYBh35PHBX/oVeRCfXjx/0EwN
dwddYyxor+ef7bS0AUnJPGKbCb4BpqcjzyO2DdWGXyWA7QhfxLCSLnN5J5D/
8Okl4RTi09mBee6HmqQxsTmauPRepZYA8VGfftDnF71DDO0s54KVzIo7a+5V
OPPFeu7k7uTeQkvdYRO6haEGFJe1vet26G8Z3vDL2dvuWukzan+US2Yj9nEr
zOhnWrVXhs6Fp9Trw6C5R9PwR6hjsueZMEF5GshZpqBkWE9BS5lciapZiawT
SWzIuU/TMW5b5eLaymKw61h6mX+J0oJxbInpPMDegjMScOjFwhr5maxC7jA0
W7Xk8OB62/141Y/ib+GAJ39ejm0P3RWGAsMe+PgPLjOdvtxtbGY/cSV9gh78
FXNuJp7jVOUH6XP44A9fZs6VTlMvknyD3qzy/a6Vw9a87gmaK1+tC3N0t3rp
XLeVjmd7VHiG9JRKq0g2zidPKn4flA4SekcwH3tvWjEXJm4JAIBsql2ILNQp
c+Gh2Fd22UMXndBpE/QNgddiskYfDSFGXEdsv4chwHe/emhrivjmcsAuurAl
3ul2wPwDHHpN7T2oL36whqEfwoDHTjKQHuAFuIGqywjwRFtg7ljXSbgXn0ph
0Hp6szzQLeV/J1kEnuih5rYK3Poy7giX4zn1K3SWgYJSJnNebnlh8PYrm1Ub
uGQfKe+uwviMJt6pt5kCtQrFCBJunvSkzljPhcwd69i2ftbZnsrT+iRqWFcp
tTGybV+Evb2gig8FC1GywNuCTjFwe0fBxvraUUEhUWExfWWhsinsAP56cXVv
AlrJ9bSRjN2bH0+sRocXdtIoMvfEd3ZnSpkktW1dNUd0qV2MnH4COp7j7Ylu
eQGzsKqNs4B0t64/+5ZU4zSV0jzAQs+RYBya9mMWiKfMwhL+8NOrK9TVSWZh
D55WQSUzGPJcK6n2vzn0wF0IdQ79Mkz5GsI31FKS5iyQrc6wo3y5wYNztvoT
HX6S1oJaTo7YmWwgLOEcRdZ475ceZ5JBb5rRkkLOFryn3wZ32KkOvq7aVZjq
Pa5Op9ZhT7SHiyMiFhKzFVpUmyKNIo1B8DkaFxj5w8MeCwrxQvfsYc1ISC8V
b9iTI1mUwy0VUhFvwNW83GQWDuWRghD+nltWGnxYwySKpDD0DfrD3tVUW2Dn
r37ksIvIp31+bZs9rD7kG4rv+WaVP0I+ObGmrHrG319ZJAHpmsBw1Xm4DmNN
6yilIVzzW8bVtceH3bYdR82/ozFZokijhLS+WJviCtRMnsymHYoHttmShYAU
k1ltosyA74Qg0BEJRnoRGdpZ5YDIrp3eaAAgaMyeu+a4mY4kOf9eCOAf2ZcG
93++vkypUGwbPNgFgqcQU+XdEi3mrqegHFo/SsY3Sti3mOroVoK16woo8pt9
oaqA33A+xtfj1Tb7hEIjqCYcfp67jgQuVHvdpgDcILqTUjuMDSgUyeCd7DNO
9UQlbZxi/23wrCsdd3pB121MYYIjTchFmjS0GoXqpeZhDfkvzNq+IiVvQqfm
WSHL/3MEap4wRzkdArahOPWadDB0FsJxDifmwAYGrgaiaCZS8UPAAbsVahUd
O5yNsV87vBUFG+1T0TD+cXxAqCgQaKYlw4aNdbXjAqpF7Bcz6MuO5C8jkhUJ
rNpddqL1LKs5BuuhOQ/sdFojOn82dqktiD6gGozmSUoFeKLL15YGYj0Oxe9H
IIOtUFJ6S7nkRcmLDLL33NNLyuPx4OCQJHD9ip6TJTQfxS6Et+Yf/mQwvKxs
19x5VMOovN1aDyAUAXOIf2nmCQso8pbs9mfZ0GrneN6UGsqR39FeNILgKV+n
XLm7vfpv1/JIP25HLsuKjIKIweEHLMJ1nHwzbmZzMh+ig54ftKEWq2iReYGw
0asBl5RYxjDvByxe/6Cb3NksOPyRZTG3WWgPuYqus1TwhR5UDmCgHO2aesdS
/axv2vWf0W/95VMS0CQnaFEJZWH0K09wGBPQqLY7JM25ebJ0bzeE+VtvnP6E
ns+otHEl8zlT36F3wsCm2oXIWgq13QhGXasA1cAexNfHKvsZH9W9l2F/tH4R
1vCy8ntWGV9CxTK+2sITELDVqwmDk/LYw5aoCv+3Owk6/2qY/6ZFTC9svWjZ
gWpZbstCXpl5UpmeevnIdOvL2W+VnftyaADhx8thvUd9u5WN3d55xXqtqw7D
XO3YcVdc7k4Pq28XOaUDublk39/eVWZWTW9Dl1I16B/EPF1E6ZwPpyVtYco+
1MHsaLaT/k5P4gNutLEoKo2sl2s3WxFw5lk67KkbzdAGztueiRcSSYz+wpXj
sL5iyya7nJHGMr/mPu/GJN3gdJZpB6RYtqt4tx04MniL30GdaCM++a8MAwe4
kVqTFVklsdiGWkv4bU2F6xuk4CjVVzezn9RHWh9RxJFgO9E0Ag51DmjC3Pl0
iwvghXra0yQZrVusPWk+NDB/hiV2qZVpByq/sj6jMExVB8iE3k6QIs8Wp4PP
YV/SuFxSFr3YVqmqrvc1NCkvqalFBMzgsmz5oywxI6OawQoQdJteAw6io3Lq
lmInTP5sAJ6rsZtN4Y0U8w7tIvyx8lvCaOyOMR8JIdhKH167cmIwX/n4Cyrs
cou1YZ+6/hzf0D8MWdrqUbFdb/rpNi8238dRKulZokul6Gc6mwiLmixlzLM7
7YzYaiYRGJjq5k+nlgigsDIyo/gWQUcFR/KM4jcs6Yg4OX0X+vAG2d0k09wC
buM2o+UvGZSoHex0pSFERA+YJhhrCYjk+gAD7cArH67bQnZnmqpeS4GB42Ib
SCTPAh6pY9Jh4LFM0ZulCUWFiI1aWJ0r+QtwvbXomqOCb3LMDLo9Qv3Mx925
0y7bNPsZvWrvo+o4wm0YTbYfTNWG8UliMZv+KTm+wJKDeDp+Vy+/IcRjdDpa
QS756vogTiD9Z9UCepN2NRmyGHK/61Zp+j/7/QD6CGbe1ccKftsBXvbC88sL
kKllZUy1pH54UfYq6f0hHI+KfiHSP1G8Qmufi670liQTSSZRSCec3O3COZEV
ZyDhTgslNJpW6OiYQkSMPJafHe/cwejtmrLfmY6QqJYgybjwy6p9nmXZFF9O
ppsTJ5JDxXyYkYmg2eayTLEsMxFp1dyp3uknqkA3l9rWIc0hJCGba9daPQKx
i7I+z/hpEC0oY7XHe/CXdIUQKGGAAjhuGD/E5qAO5eS5KC7fBKJBJ/FDFLKC
m022eteVHvRM9McAXooSZAZWhMsvV4RPjmpe/X4d2QsX1TtpFrVUhyq4i3+K
xaz/fGDSuZax/ZZLCPBT/qrGXb4TGV+yQaBcDaSGOpPNOAn1cBdq8QB6G9nx
6YkbPi083SVbvkbIIQWTPDfkG/VpWn6jb6JYh6qREeupGgwgI5XYtUqjnTei
betAU0gK6Ur6rtsNnpJQUiy1KgnP8r5yzGgqsFsG0cQhGHi69QktK0D/4vCf
mwdcIRhk1zmHgmD15uhUikd76defVxQFIyv3sORfWxdSKM/rcpsPMmlR315N
Wa7QiVwlGmhK9EaI6MTSDZGuMdqRgvvXUn8P05vyqrquHZcvvtYa8x41EQU+
Pc0nnOHWEzhsa4yeB17PVzqCzikU5+ccONZWj1W2UmCveKefW0j99Lru74W/
vTujiMEtd6ShYEle8u9r2Ja6k+vVrODh+1bThutBeq7vKSY31B4NOWusYHxx
ucNCulpSw8DofiM0SZFKaQ/7zqNzbKE+R/GvXOau1sNkQ8D4eeUCtRRns6gJ
tRyGLco/6P+A/fiEdYB5uRbBuKcIJZAr/oCUTA0/Ogoa9yLoXbwJvtWrGf6y
p4X3yVy2izA59E5aRLDCfESehzauWZadg4/8h2Vr5cpcWyuR2+Zi1zzMRElF
16v1BvNT0hILhQoEJw4gOxdFHRs6QdDx9KG0B351sR/W7fsJvJGe99tOhhHC
SZm1lDi1q+KCMAkeVwD8flUN3iMJZt9BkM9BE6H3MANLRD7Ieh1sc407z1f8
24r0+BNjMC4ZWo6Q4XIiKEFmMQq+uMns37t3OapoGzd/3ire2BsAxT0JxW2e
8XwwcpLTS1g1yWRmB9ra026RYU6meExVck7OQbj6QyIGG1JJxqbAZB9XNcR4
vq++H6xs9sZPqphRKjKoUxpAF3u+NUby4hveNuycQ3h0Xl5XMiz2RnmtX56M
oOSgkfknHskRFF/MtHWct5t+8c9mzGVP5+ekNW5RjyTnOrb3sa7bfY5XYpgP
0XiztcAFFZVX8Cl04xT0LeHWFqRwpbyMoZXeZSJifaFnOR886spwjv3tu8ZQ
ObQI1vgcY+EEle+6228WfZwfGQP8cPRg3kEW3AKo7YcnBiRw9kMMeOts31jS
ze2eAnefaN0/6rpmda22RAzqOpgC0CinPCuEhgdK8xnQ/GJ5jJWoBU4ag7Yl
dgnMsuv6AF/aVx8h8+QtN6dQMtDptkB1YKRiGu5YdttF6+B1TmMvDjn3iUfD
HN05wy0REfNIyS0BnGGcErTHuZM6nvX0Ar3G4ZPHEPOQbd7t1ckuWMbZ1hqG
KImfq5oIpobVWKAZACPFzzo9Q/26bFLIYIZK8AMzLxqT92ZdwK4uvmIVT1YQ
+NKuldIxUYKrMAsCQbx3aJlzPt/RZq5T/C1YDJ6Tedbhous11cxOrxUm5kBy
h11hVwouyWELFeG/ccUaHQ9Ba6DpO0eH/vVxVxnD+482fEEDr6sKt7VkvGdT
SAUH6YIC8jErI+53/3+uawlE5ldw0AXcSLAsAbyeNYMEirtaOQelg6VGKnNT
GJsztr8izuM9Wn9oRrbydYQ+bY082WrVP+y7wswPEQFERa2vDYS868VLvsKL
LZF/haPAM63EKeW+mbjX1dZQ8WhbK4sABeC2UZ7CKLyOozCx6yMmuhKsKZ9q
neKjaVB84cT6qVE6vrH5S4NeorMD3hiPAl4XFTPQZY7ve87RtePjrO4D+x13
S6neEiqsCwGbhMmGkrxfDkK1kUfVi3C44FG7bBAmU4tSxoON2vHdvb92v51a
hpTAhrO93JbL+4nNjwdvezk8aKGW/6Hoq94gHJZjmK7tWi2vZA0zjy8Gzvx9
Bm2PfcYkpUs73tdv9Cvs1DcY9ic4J2RXxcAFyYXkb9ANtoMK1umWZ+vRm3rw
zAcUVrFOwOH7qVwYt+FNIgJxCs3OlrvsPimd603oroSrFnECnsqbXG7Uz7kP
zxRwnmIeBlo/pUSEQwmabmwz67vRplX979H3VEI0k97qpvDewvrQaoi00e2P
KBZB4CF16u4dqL4oA9vGnUVjBxrN6JjCaE7kf5L/9GIQxLwxPy2vADUP7fei
DWXiqOLzDyys8oeuutqwpR+MXWSDud4DFw2dlaQ1ffpByHp/7SAyzSAdvZB6
e6AINBVNXg+h7Nqf2/2BsRvOyzvKKPxTSsR/WDngo/oZ//Aqi/gntnYXAe0t
1MMvxm2m56m1O9sOB9IgVnjnEv0XLCpZeZe1KA7uhgU+fVVktf6xy2pd37cr
RH4dpig6sw62WZ2F97dThC0qlTbEpKUxp5m3lZ4G6cQw4Hf0Qy6Pmb+eWZeo
PCs8HNDiEnHEPsO0UZ/U/i5Nlyt58pKLY8Q+B5ok07mJHPc2sMBDARGza1ub
wVkXvmkyScgAoYyjJsqI8N/rfavfPOyJlJyAd0DZQD7XRbgMukXQ/rkqHCsj
HgyfFWZOg5P2Krx7yrhj/bLDhvknCQXNZzOfQ8e6noZqsB4bDVTDKjWnJLfo
LuKnf7b91ghRtTt3IYBqQ7PnV4pU5ouFxUISbmvEUKhuynltvo9xQOe5T8q6
9eke7h64oWFKkaIyMb6lfLSOA8Y9e2DNmlNTRGdn0N5rPTTaP7uyqKnWH416
+ytb7+oun3rIuJ3jUlosdvd1UsfGXsRb07hns9mZCV60mPwJOMTL4SFrYupa
OrOnxT0uzQFl3zpBiqajFMZlu20zii5NTKe6WYeqmZkoD2RAH4l/YA05U3ZT
djRa/3hegFlZ99/t7rApjhTESndI335kkvgJOg3QiIRaBcKByEVI2pD59rFF
TdRLzPepNqBMYvNT9ugbMejHTkTOkY+wQTD7ieDONLImRBonrXNtLT+N0YbS
9Yc6V1jT8FXxjUDcE1NXf+T15D4rOa1SrwJBdGj1Lo4bEGpz2ykhmB4KPhF/
w8U/2ZAzDlOVxBY8HibLGNsJfNefEffkae9U3CM0ieKy4PFBaSMLOwTUGg/E
IcMCjAsQa0pS0mO4yhZZQCdbyCWYHLeZ/0848XlqeCNqYugvKfynyLUcK9QQ
ndjAqt6UMhve0ziYs7SQOHRVqhZFaD5V+taV+zKwv67szA0o1fOzI/uE7Vvp
h680iIS6aOKhrRspqZd9b4WjQYuvyjZqJ8c6spktvNSAdvdKocyuR2Z2LzXN
Rrj326vANfwhCxsbeKDafyK1WSkq+wg3A/Z4frfvBHeQI0uLeKI7L34Q+Vdn
MPP1j5omtpldAEAl+qmlH7BRt60KH0GMlaHdCDrp4B26GyxNTZsVwQ==

`pragma protect end_protected
