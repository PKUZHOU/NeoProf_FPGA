// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
TwizZyjanOg+yoiaDatEG2ENo4D7aYIOptqXe5WL4UeXKFAdYB+5/W6IKuIBkGi8
LaH5ZDugYLA+/JTWjIHwxktgQxZQOq5J4fjY0K7Gow22IS6ooVmetc0SYR+5f1uZ
Yo2dfPrd9+9IzJyTSNVOD8tOEfpINlfgWiMeWv0873FruEp+1OX/vw==
//pragma protect end_key_block
//pragma protect digest_block
kt419o/eZGWKr9lC6X2Wltl1fyA=
//pragma protect end_digest_block
//pragma protect data_block
Mf/cFv4ikDZgzxBh+60UzdJxh++eSijBm27IoUl3DLRfYJ1LWbYy0kwXwdKqxtM6
Y7voXTn125nQ8/YWsoQ31DfQUQzLJ7WePaWGHJOcb3gdSb6A5g6Bibt8tyYKawOr
RMyK/tB8FMgk7DVQOcpo0n+WpDWoISnK1NNW37aM7nlmZX1oDKVi+1AHtz3BBQCZ
SajStw9IpvNkYVYKVrXuRBkm9hs7OKiLA/aEJqnuqqBS3k9sdTr8SO6bJfdZ1GLz
Bd1d8inhpj7uZJ6n8osXbEzUnl8VTvw13qYoCUFsD+Jdxv3bFIrs5cTD9HCHfPtv
kE+1/8AHe1pquK7RN0uLvAbHwna0sFYduUm9FqvGseiXzjtIgaY1mFIQBXn635+X
1yEpyXR/AS1cG2+IB+/crYCvf3BaJBtT7VJeFI0DTjuuckPwSXuYwmZYdqW775Sy
T5WmdfFuTs83vgpFu/g5CdOZDulUAoSLv+a3C4/sy7CUClatBMaDuol5F7sJm77p
AapQ6NY7Al/NlXw31psKIcNKqsH4mXJuXMOiHzyh934NigzLJgsRnDDmQeEnxLpU
XnrBqcliZpg/qSSLtK1xF8VkwD1ntPUBSXUQDQsLbFYbUn1Sq8yyg/m4l3VPa3tm
AQBnyS5AGnyrlupo/N0fT17f1r4VYBcZN84UdGTQ08/YV/1S9Ceu+i7mfSE0PRkx
pwr0EFmd8bzwjlMVpvplQPrvzV+R7LeRTekLO1mG42p5yaE7Q8cmxrp2OjujLerl
eW7CQXPP1jDQGje85PQHtywmgE9gfaaFGcLn6sPiJbZbhkw+X0eHGqT+nm9trAU1
W63Aa+Pm0K+9QwD/tGcEIWNG3OCE/uG8XEyNKuixqIuRHai23QoSZMCVLqs34Izk
9Qyp6uBy+dbUNiub0mGdFsrGKQ6jc97aMCSKLbfT8L63dxpWVxjUGYEJqsLCe6R0
PW0xSsEyBzERQYE2Z8DTiuy2UcH3AhFO1sO0Q7wqQJjt6jzKJNPgfJn0Drb/7A0s
Iz5akp9R5PcGOCGjsrv3O4ORu95ME5/xL+3MeuaXeGuIrgVbQt4GKfyRfH3Bapb4
Gikxa1NjmLPMNKvFDpXs9losgr2pzzmaYCCl3TXnYIXMIq1kFRD2pQom1y6bCgzM
oRYJ2tL117TECwM6/KtNmIdUUPn9dIl8QAmkGoOR/fHcgBE9In0wDlbQVNuou6CA
C91s8/3PpwLFapRLgQGujOjLtez5k/ztspjHKJ+SMgbxACzYQrbZWnTXkrAiS4Ny
5zoebC1LT9kjLwciVGol6m3VZCXtwQ2xhUgLNwOzitXXEigYjXtkt5gJ4bLvwBCd
NQjvDRNeFGEsUjEMOUqroOiIU4+bmgjsyTmaxt0uE8ahNEMvBQ3vpgB7Z3miNmYc
JkQF4/K59ZLW1VdqtTwpUr3O7NjeuDPWUoB5Gv2NGeWokv9XDTJaJ+MbFxOUGWig
GK5dEkoAYwgBqvs6Em6hKye0FL6fTrUb+zYEFRcoeZAq8Xjg/clRivki0fXQWEvo
peNHD9VmNn7kshKjJlQEGqwe3qm6NJ/h6V7wl1J+VzPiGBARooGoitaNyTgAgaoN
1Nm86aFVfr8EDazHG6pck16R/sgHyPg4VXuYUKs9JAaOdxL5iAvMc/YX5pZpsZVg
SH+xSy26sxzASeWMnTliW/gjLMY3K8TYqMpT7lFmnVzyB8+0Me2RW7CZjifVpLxa
Ry+9mNY3ou5eKQxGDY4GnZb9wHvLh1Ed2b1457Xvs/ZIcVzBIh8jU2gT1zeHbxd7
opkA03YIQ6lH77N5aLDCaAK5Fyd3NJ3rAPAqmDlTEF4cCP+gduoSL5/vLmIu54Vs
1KU3ScyC4qbuOC+Ft1BWjzCFTCxIk0GWWMrsp0px/DWho8wAXlVDMbo+585a64Ni
0iW9aEzbD0XOHFr89owY6ERDtkYr2x/tLfjwt8IOnWzIL61oW4qfmogCgugUKQfp
/cf3OSm4nbD7qFXoutt7I/psUWKdITBLbDtuTrUJE8IHtaBe4h6fyJhg5aXLIoLW
eJ8lpACW68gIzCNEFCuuHZasMDnDPeQAjIP8UFvyvcPiFpCEEl5H1AXKMylNkqlS
aOY1f9tOV9Vr7/SV2LoLG9WFt/KFyt2aDlQ7D+lgDliHVHIZzn7aQjHvvXoBWeEo
eGAb4gQy9vUKbgiVE5OO7M4LMMUjzBEyT5RAhXfxfBCVhDdkNTB90QYNCzFT/OLf
7fOqXH/ULYvxeq6CDAXc/kmnixqO7xKYRYmI5Jn43vlw6xMslcYrslsCqGSaLjXC
L7KaFqwlghMd31UVvycyptP6hJUUUsLo7NMTknx/rRaTQ1r7KEzy9r8lsciuM8/p
+OsVxhKkhRKmbY4FFfdvq9+XhJ6V07rwoHTwrSPntvWBniDJyx0wwHoIsVMAeIlT
ZUvJMu3CdKNizKFZ2oGXTuhaMw8wRdb4faIhkUc3J1l6I8YTAmPkC5o8pRQeAKo6
pKKoVjDzeLwo4/MRw00MErLn/k8uJhuA6pyWut0Olhrd0s8zyngJkWGCVIMMndkC
pB1VPVACV/KKw2rRGHCraSfpfGQvtdXynDVzkYU68ErNXmRcW7FgaH76oM/XNj6+
6ZGj/WnjV7pEekPVQwfXPjOo5C28c8NAgbjTrUcsR+D/OXIpB+jm9e8ag3A03exH
pk6C4nukqgkE3couVV0EAVXIFhgV3vACpDh2nPNfi7oIb++YmhpjTJ6ea9CUeB1Z
uvt2g1JOY0HUU5WBmDoX6+Wdu4cFcUUK3YOOPG4C0xINYDh0CZQB35EumRE6fG2R
gERC3awJJgYvQ00RI3Z5cjdYPatVETpASn2FjRVNmlWRnPYw/7SvYQeDfEG0ShlO
vpudPhCRlwtq3WO/Hto7eudvHKQ2sLtpHSN3QVpF7LANE/prUsvoj+HuApPqjEk1
JPAPnc62qwoORH1u+Q2FRwmAE0o4hkUwOW7l9e55W3MA+qBk8fUHRavq339ONjAb
7h+tWLu5eIYEANYHK6nEzYBEwtKoOUfayaCm3JpsxI4t1z7dJU7olrLgVQLKnmIb
qM0aW+GvCqEYS3VK91IdmieX8gh9sV1PSPsOBhJS8tvgYCbWI8WKQQJdDuLSx+Vz
bcpnujjEoHX9beeDiKjHmRP4NFHxQpl0amj+da7z/eLdOZlYFIGo2uZzn3bMx/9w
KtdtEZ56v1NzpwsJQ8DI2nzBBhrYCjFbgGgWIFRmOQQHvW8DYCD29T5emQuVxzgP
wqHAyhUC47f8Ki8134cm07S4Nb2gwV0dbBRb5Cj1gmBsQhUNidkkarbFdtje+RJf
nZOwy1hz+AfhXsLZtkCQdt4F42LfDcShZmJWZk2bsJv3Ux5h0fHvdG8ldycbMKlU
4qH2AsNbVN54kg5EhozncHztg94yQS8s3TPXG9szmiQaFfKQxvMjvniBbQ/IQGdh
MxtbFAeiSdj2fIL3+8Nw145OhqXMO+bPBEdMScJ8di5DTG89wWGN9AlLlC+i/ifU
c5PaPCBNNmIUjLglaZf7adYCfQfv7e3eFVaZhmns1x6YqTfGo/pDmjXarl2js7ot
jOPua+XbIWJG6Pa+L4phiOztT38/vHcq/gzsPrF5y93HtEm0frnlA3qOB3c4Lh60
hlMzHUaaLpn+enmwVifKsZvy2I4jkeNFtpR2IldxcEXfN/ggfX2y2Qif5mknjipj
n6aH6xNcqpgcrEInb3pcGmH/6dC3jiSNVK1FKrGeCiwrp/bGwsZOuIqT01VL8fT9
aMs0rfJEo68Zdeo+NLyMpZJSdKHYEIbqsaPlm1+HMagLsgRM50MVnN2eG3gW5qno
slnidjauKLAxbSuc85OEtQsQtmjU0Fjyg/uYT9gT99DmveKlavGnZ0wqGMdvPiTy
7ybpjDagLdpbwudQfwGjz8iA/QgBOXDYWizT4PR1HeJmFwME99kLp1XYoHoZoqej
ENkRkmSrUv9g2VETknQo7dYCJM52cuntnzLmL90MOmwUluTzY9L2/q3tLjJBq7dT
BpEx+/rAjDpqIdBu3mGirRTXabMrrbBm2OQFfTEV1BfbUkfaQhWudtdWUbFsg5IA
AmIb2xiOTfDzCRWe7mejyFvMQ4PRrKGNgNWqJgLxok03BVF9Klk+2SeiUH00jSl8
xjR9Fbx6EJy2G5lQyGW6A8CYh6pL/gTrraOpU66EoXy+f2oB7YA2wVecTiHNRheR
kGc1/BMYfaYhnZBjKJt+e+P/Sv6D+iCIv+ux/b/lfHI+tl2tbMivnEVEsshl4lM+
6rDjyt8Z0v8ITUoPueSbXlUrD9fB2ZOOOOaG+dNkDw589lTnilpuMSmK4YSDymRm
Vg0T8xdcaRNE03O5v8KLOUKsbVpJLocCpKBbp6yWwzbNtec+8QVHTmm0Uk+2NaFR
R6vetPLce+MKJXXnEwZiM8leoL2rbmUFfMrFbHTCKseU+W7RgHI2IiFmC2GQZwZ7
QY6MxQiy9OSX/G14fTahtY7m5Khjy4htkJ9mq2/Q1jJQrDQo99f0qEOjmq9b0nLj
AEd+tz660OWz69HX7s8/aXg8ninEE3HAYmJo7S/Gviqd4GAWgEz1UqtElF5Q1a4K
e5gKZeoHlUbh9rWT2C8NbY0E+lVP81btjTmTUlmSfsewxBjvelnTMPQkiagyqZDl
AMD02gWzWxipbSdpKTigiiTREGOZmGU9XU9xPSrBRFVWo3ScLQJK2JdnofL7J8fm
TruzQbSB/bxak7pc3PgOUPsGRX7JPMs1hTZRRZvT6pA1mJlSvVUXiJ0xu68M+XeC
uWSW/uRsDQIY/UwrGgT1HgRv1gTmOqvxbkDi8Ql/+w6fml6FEXMqonQxu/6p6SoQ
pBAiBExErw1U+FSnF3/LxBH3+CxsuY2b6MK8jwculmDvkaeUb5YNIsdMvlsJmo/N
wIuq39T672CLpJ6PC+y3ozr5gAZ8p2hq+pS9YnzKLJg2gmeY0QGsvDQEi9TqUKX/
TIdkAB85pPCYuTfI173cUCvXabcspYU4ZkjhzMcwJ4gaJueVwwUV+zkgQGudHrt5
Ts3QNDBYutQhRBFahevXh8tUop8he/1UcjVkr0Sme6X6+uGABXSstmhkaWvr4S0U
N9wxFM+SqnTyBBMOsTaAYBjIdhmUQHGanIzSh+d++xPzAk9kJUgHAwycTr7cCekR
J+SvhiaH9QbyWIMciqZTFueCSJlu4uNXnufi27xlHlvDEtM0kl9QHBEz35L76dnb
lze+DvIgArPZfW4T0JAPWmWKI66pb0tkWgB6fAsyJBKav9Ho7LIpTveRLKd01nqc
m16Zd2seU354YLbXWOF1s+bVqbvAoCUKVxPdJ+qD73w1/OHcyGDR2InRDpmM2BTM
Twxys8IQdeYKxaiTq1/edYRQ5OJifgwLWoaqFCuKAyZoBNpHkeSbE0omJc/om9JS
wBvJuZQx7fZrWYcqPdPxRTAE7ZfGuEYm0thbY7B+amIct7AmEwt36HaHxvWKw2pX
aOY2po2BWh5R/CHdGVXd+dNwh2ZPM1s/Np2pIagzE2FZaKbbH9zRAnrCyD6KFfdf
sXJ+9gUZGK8DJ9DC4fULng5Zins5aTXufFttUVI7+d7u6/kBvBI6xeJV71ljTjRn
Fk800GCe15xi+w0RBmeKoyQ+kM5Yw57GgRt6uniWMai0AD0nKBgkj+jtD3+fjJOu
eEztCmGJuKHadmDP/fKSSEErYgmtHu+z30PWweK9OzvINAcQLyjCp/r0H8XsGvz+
P1k3A1Egz9KuxWEWGvgIwvE8m/kBt977IKnOuZFg5xIeZf2t4cceioMCfSb+9zuI
RvjNZejbHFgKZy4G5bP/aooHhT7CDRVreXQc75dLEfTXGlE/24QSLlUg/T7RfjS4
Ku/p6JFPfhGPQaeXkr424TS2/PJEOL6EekdjKeOSOinKmiEd7GvP1n8buDcgbqYF
pcaF6FtNKbk/lkPxQIJCjNrYicw9VLfFc0EzDShgX5JuP3/nlwy4UHEn8mdb4KqN
sR7QjWmG5GHwqEqo5DYhw7pFDlk9GIog+HFXuMJ8b5qT83Io/4/2mfIusxUJaWYM
78o8PNuVdQtBqePLcGuiUoyhHouh9HywcUfSqDg9tnVjpOa9ziGTfGpSzdvQIEHn
jGTLQ6TCDm4RSMaFNEzNwFn2OkCot/YNwXFlEcXXre1yZx5sQsKzgRWxD5jI3gtK
WKtv2UyIL/gXdph1cVwSFJ2Cc6bcPb6mok1xkHBGt4Owry7Qc8L7+0dp4Gh/IGnO
XobFHsTJu6MGkvK9yZj8tW9bCNhW4t6+gXSVryVChwcbnEZaPYPgO6Vb4HOHRzIq
QF+m3b/reP78w8hmqqdpPopL8X/KTOp3gb5+s26CQJqjLZHOjGOstnKVZIQCpS5/
tuzdkB+j6rGYm0urn5xHpsEEWfd99X61+MqUVKjmrZrQDMPoxP5L+tr9rUTFRki1
oRZ0Vlz3K2Gcwp1+FuxHxF+q6N0JAYWmQcrsF2LhDaBpNKsNeRWlbuq60rb1HDkH
DiPZj29u29xPF4V6J3MRY9l4Dhq+FBPweskUui7JEqY8rprKzEjDmJ6niwRca9K7
wSLHMH9qPjqNrwKqTTD+vKjNJMb9eoWcRyo4o1mQQadIJ3mCUHMacvV4whV6ef29
dMGPziqmxOb6kdW7L5U/F0Xott5HazL8v4dhd/yvPXcNZ0UkCRlcAJDT63bWxP3E
e8L+QCAKY8BBq5pWbqDHLJmAzPO+vUht+18/ZS9Uw/JRN3hx81S10GGm/5y5hJL8
bGZoQXN2RvheWCQ5fo0pYMu9f0q8T54vP0EVJQZ2Rc5mPqf4VU3+v3Doh+mqS1lP
u45Nvv0fWBIIDmyfnr5JqHB0V0ACbUPg2Tr3ANSg2KQCWzw602DmMGUjtFuLzBLT
JMJ+VRduvo/GvafUqHEsZZJ/Z/W6SknaApCNEy9chM7Peao66cGtTbAUp3IeVU+7
c8T8yNmjyd4BY0s6Q7e18rzuWWS+UuvfPs9t6eTOCy7tnfWokiy9zXAQS7POaOKD
bCbOydtr4n5bp3JYLBQUJtzQkqIoFS+UGGxMdjQoMqvN18xWWx0XkoWiunf4gu/0
x5gge8UM3283f4ihwWrztQ38etMgt1b3eiUBSgJtKe7I1S6aiTr9bJMn3fnZ/FgN
LRNc+KNGFw/15ZB0xj/RZHdjhI/hDpzQHzOFxxk8Exe/HKgmdxySwJuPI084qwiA
3OCO9nMsYFXHG+Hy+jneAR6xV6e5ZBnP5XZMbIcAK7zr7yvIobLhiwWOCEGNkF60
vH8eoizJS8Jls6dJbsAqUD6nHp90hn9Fxu3NNYjDF0y+75eUIjyZaOcNNwMLP9tB
0v2NJwSiDThrUtKb1h8NNGuw1sksRzcDUHu9t5E0lwLS1FJRL1DbYPu3rPMSi/wg
vCkItnYse3QO3Y+nYWf96yKOd0ZxUJLtgBy6VtYU88E5i09Be2WubMNsD2YFPg7m
3P+G9zx+HxG7BSjcRzJ6tO8X3e8iwYpHDrBPNpuk1eMbpv91sVU2cNwb7tsoDxlI
ledVGjFnY9FOEediHVcPAhA7Ym/QSNT9SxZhe4mEdwXM5YO6yV+FLS+eebF1Rbcm
NcQjhCqzoDynPpt38okUIsK1LQmKoG8wLWDIrpzXsxoeDPOgMa6xyzrngQXX0SMO
UacbiFGwNFlfdDq2TkB/0W4kBIqvrIuu5vacEilpMGtlKGrwfikFmJyacsvnwR4L
UokllugHwJEkcyE7qf7cvV3sMf4Rc5oibG4Iu1RPg8k5Ue0AhfOfwGpZf/JRfTWa
J/xvUksS32SsqwTlHQ1/OzeDRDEQ1XqhfZ5EOVhnnZWUtJP/4Fq4999syiEntyHK
8uA/Xx+4DXvDPy88dLMOYLl6SuA3/TrzDojvSqWpjUOeJw/kjyWnQ6k/Fi5YQl8z
4ozwa+Kc8SYUgtfDHEX5u56yc76haGnVjMK8E0JCd20PzJHJqlZ9b+waUWHFo+FW
s0K8VsFouzkqX55qgso62NkAvChyecwiccww9iN2RtlrLd2qgDmdD46aVlznhqH2
JgCx/F1x0dGQSZH4bUk3RRxPeUfG65IDk6t9cW+JQ6Eh9Rmz80exUHZaC+bc9MJk
Qd60jZw6Mk9aHBLpqvdCDB0w+7DQwCdQ2x74AXuhW+JLJblM3iXLS4rB4J3cY76F
ugOHu2vrJVqwib8a9tl0e35ywY19Uepbfh39pRq/xqFMkLS/KzpAkgsaAfYY+9RU
LBsbWPWcHJKumjXDHGMwofIrTWt25SYPLEdeb3jsEQc88Goeg8+Qkz2+3oNsSgaN
aWY//ClaByKO+L2VMVZl8R6912I4/q6pP/tuQ0RqZT1Vqo0v02zdZV2vwFsv6bv5
ZXF6P8+khX4wmvktfr/FMXOzjurET2TQ3kiS9bjMb9DAdi60AkL/SrpFNu+Tk1HH
GcDh4KtZeX2LyuZTVO1aiunWKavkKj5X2TZqNKFKoWq9eZH05k8LCL4s7oj0okas
LJ4EpS9judNm/miBwfHXfK9XeQ5PbBp93HcxwglJwwkwMCRiCksPnESivystEuBm
tgtWyntjYfwSOigNU2w5N5gsZm2IoyOtKOzf4aTpDnJA7HIcYJ9X8xBAjcMjrxGv
7DzpTVVewCXFRPcHaOdI2ER9WewM0cNEUkuM0QWHxvrvv8ykPbFcNUm1nIWy8ua0
9LTHeGAdIHjWhaxF2ZUOCYL7jnFgvxSC/DpaTrtQ2AKrfYLNZik20D9/0eSx2v54
3PsHlqkul9bebyQLgN+Q/aUQI+Znuo70XclbaV/CzpUrWbQ8d2rHr7NzSnhSHm7+
X0908YEB5q+wG//fw+vQCvDt7+RqrMxRDRoPh/pg0rF4KlT0iMNzkwoCZwhJ3urR
bwmL/ytxFM1eIAJ+y2dkkjfh8f2FUic8Ds9tvmoeYFFEFMxvReJDxTjjW/Yat24p
G8LtUL7lz2A2oEfo7NogiNBld7jSl7IGrwGUVVcvg51geSBMjJtd1yUkAjW9LBtw
Xj7QFQjK5+ugqjXKOTcBBEJu0IjzxGNzNvnR1OQaBaHCG1k3OzngteHsVmmStkjP
Cu8Q6hRRdlczmujrow+BJhNIrcmVdm1/D3tjGi3XHiHcSLoi4YdR6773G20YM4t7
YRIKCvUVhk7FPJ61bXXgsLgntwuVnRH1ArLxEFWMpJhDKWUd3oaIZxBQgRMUCYMk
4xMtLRSw+5KO1AhpSx7p5UajbEoDynpmxqxVn6IA3Z6cY0bytBcYw9M+xWY/t1J0
GJkvi7arhkom4Xa8JAF8RgYoGLOGW8BnYDaI7wqoECptHhkCqcSa05dBENWU+gaw
cvQOBQG6rd0MeAq4pHrpj/pJRoXcjSNakpalW/12/DlKSF4XVmK7TMM14EUR0y3d
waRYX701tADd6K7prH3Fp4Jkt9nTClvoOw3MKbzrXFR93MlDUkmz3jEbWd86HpKC
kNVm0Pte/70nKc3ExqIC0VOk1MloveyG7TKj8I/YuF6uj8N+V57GLBAdZgFfKNsC
a0qNzIqma41quwJ03AeyKNd1wonAw295agYwR1E8AyS1ZSQTz6FHktMJaJ3jkvjp
sqxcN4aNix3eRlrYs+bnP9GggGPx9FOtFjJ2osOIvvqFysFVC+lD7zHmPjCIMGB7
ThNa8ch9w5z8w3W6PCky3LPV8efkbLeHDGqq4niPFaQhUkAg0wBVHRd92kM9DrDp
4MGeCHWIDOWNmx7rXpYWPGFHtPA8hRjhFxQQC+Gz0mGMlbx8d0eI/hF2RTNR2us2
6iVIuUKXCNo4hHCP6qMKgM1tcrSwqylQtEn5X24qhTfoq8ATZb9bzfxlRLqLbnQR
DAKjLrcv0s+jGt2wiODyvvElmlMtpz5SRdUnSb81iRj8vxytsO17ZX8Yi6ovEj4M
ffIKffiLlfAD5of/iw3o9HRX+2jieb15Z5KYskttnFvhFIZvY+RhztKWb2tKFDJ7
SzcSejL8b222q7n9uyCMi+BmkOAG174cnsFh0sQ983EQ82qvsrEu81vTvPc38cPS
wce0R83yoihynnnHtTVcix7dmI4jZ+xRrtDwu9KxHlUa8jCWOKCKYgiDX1dAaj4Z
9omZ20UpJemAoPIi5LKHCwQdmMEaNqpMExaJaWeYmRlq4ZjWZKa2zifXgv1WC92V
o1n5TlJ+zt2tZcTv6JuEb2MqNhvecTE37Os2kvrhYGyZeC3FawOsEqFD+tye/FoE
ktC7N3XxTwI/jwfdI8UXgM2+NZMhRfzIT22RezYqNDT0PntCIns/LRq0Tdttfj+i
GyLwQbrO6wdQm8MWSBIR9/AGznSnyHct1AwqVQ0LnbfV2nmeFlG0BZDFUgHajUGd
91uu7L8qpTxRiQit9h9AHcZqUUmWM6RRkOZGpsUahJNprAnqxnsyVDG1To73gzb7
NI2TkyzA8uT5vNF0DHi+DdkEHdHt3PgzF7N6XNKmzJuUIfq6gYI33T6BmpN1KEoG
THk1rLOypxcPmg2YpnBwUmef8MpBjbykL3iyOkptRsL20svdeHu0vq9QCtX1Ab5d
PYb74y8FsEQXtNHlRyMIP9RzUSPzdoCUSZWRkL9BTrC13CkEFr5w7mE9ourhb8WW
nyBmYwvoXhre+42sqxJHaGtBTOKNwxKCVdRQslKtVCOOPH99Def1+XW0nHLaq9zx
4S/86rGCf7IxzOZPBDZ61Mb/1mlzP6pl3RlBg/637TFzi/8OYr4RnWUOLdExmeAn
b2PilBq9JS1KJJoy/S8GmXHVfGpl32uTbVQhVIbS7gCs2eZiY2Pg3WgrPwpnQV2x
ETxHTfGHQPI+YY71zX3YhwFuT87OCdn6o8G/RFPZhvv8GURbFSNZqvzGUQWRR1sj
4mBgx9XwfZNb8Gza6M6vSin1doGofIQJ4LY9YBWdPcjR0e6TlfxTzwQ7fyaQ7Zvr
KsN+sKWseHgx3WWfweqABvLrfg/xDRWhzmcQox6DBLfhfe9EY6ou/ftFS9B5pMFG
SQQ3oGmwpN/aX/IoWSOYgqri5w8Qb1eNOkvLfbgVdcF0DSnGy68EnLxbMNdkH282
x0rccviw6x+09zUiV0TKGG8v2gL6Ow9njf8AxdXsqKQJB4mzjEKcb2xvfn6ItyW5
67KSFLzh8mmVIo8on4hBauMMULWfHFmKksUe3EjMQo/gIGrum1xBRWcuSinIsB8A
hyHg9gIkTZi/IdLtqeC/DHN5r4r49R7Yub7qornlnDY2Nee45Ybv6jl2i/ACjJBb
lRmHtcc4usUkp4s0lN0SlHgaazg0rGD+9IGu4ZOBq34xbPjnM5Zfnk7667pAtGhQ
IuMVYzwBcSS7plqb9AFA0fb0nPaeL3ci/nihCxYWRYP3WjAlDuWtcOF3UIqr9CPj
3Lcqg7gSw3Hch4zpx4XeKQwOQ35fLxK1vMGo0yH9U8KHbUefliFHzy11EPLgjG9a
6g2BCicDpqFCHUPLGDPQUkVaDl5AkT3btwXDIYXnHsOLIyqJr7GRjYEcYaX8GYDE
FrzeHN4e6rRLm2aTm8SDHuFX/ZQE5IriXvBci5j7cL/RkQN/CN/EmFZ1VIxzapWJ
0YkmkobpMTiYFbLXZDqZpPHobxBSnaoxhFIato/vdn+/CGubHKnHGRI9ErqxMzvp
0xj0s4QqRnq7zqZKYlZJIbgDF2nJKVvg6yu0jpXUxTv+uVciB/ajF+Ob2NZ8EqSx
URbGBcWKYTK79khNd2Uu7W9fI8XNcrA+AjukczcgPyKLDme8j8TWnwcweX0I77oM
97gFVGtyWK1/wmxGBBebJzteUTETYyxXCnZ3lJ5FuoKDUJPURoGgAu/sQ3n8n8bb
t8BmHhBIX9vf9kRijzSHu8y7WMmt7RzN5LwCSaXN5Q1dWtiN/PsjppufuCGld8AA
DTo0ryFmx3YRMG23mjYthn88xfwqd6FqMTUfddyeRv0pEZKm8I++QvA2NtCyjDQq
8yTs01VF6FqXVYmwOc/5xeoQhWRFjZ/J7Mo/ATrjlqRfV3XSYWoYZgXL3hW+nrnM
5jHbqANAkhAz8LH7ntYsGHUNKvCqIWtqArL7APaX0uCxKhH/IUg/vL6BZn9B/4Ys
CQXBAmxHEpqZ3o/Z79v/WiopDfHka/eH71FU/xD/uiov+Sh+7Pi3jjrduVBO4jo3
+qxbN5FKhzP+n0xVhpUKGjhVwmAla3rUxXs+jONIhuxyFG1hI/rGrToY7EF67x5/
Rm9KY4laG0EuZ8s9b2/R821JbNH+6pUeBS7HuL9WKnVGruCZC50FUaQ791gg9WfF
TLG8rhPJ65yP23zoLxQgsiU2VNaCMthsmA/mVtu/oFlNsukFNqJbRv4y5ojBAN9Z
MurCIe3ViosRpw5lZ83BhjdtNvk1jA0YNyQ2SAFi+l6IpkZztnuRHWxg7EN+Zoto
oXtdMhzyNPD+E1kjlKdqr0Ouvdomdf2ocQ2+YeUBP9s3+TE0H7tlFjwCXjhBlzyy
fFBgbeQnfWjjV+RJoUvAG1c4WE5y9HDq54k3yAMzQJhZ+iG7SuW8b44ePK2X419W
oOSQYjRcuVaxowJCJRFOdu/o2tetEOrAaU6U7SPP9di5Xy5wp8GGLIfjey7wtwHL
FDtM3z4H2tuX4JmSk7GUlDg7Qr9EF7TG7AVLINJmX5fUMfiQIEWsAUBavQ7Cl4HK
zOtvkrBSkpSzKyxL75wY2UHhrgPVHpKsUro/ZEsb/EVFu1NP41vs9QMwEl8PLAbL
HDqYtVnd9iOEKQhj5xvVmJKaZN5R4tBFSI/y05K2SOr6chOqNsOG7JI5k6QN5gfL
dD8z4Mw9Cd6HW2CvQr6QJmlxf+Z9iXjIS8W5rH5twmwW81cMrdqpx1tJQQB6J4Gz
6+CTKNpszqflAl+gtsQQAWCwtZd/KHFOo7fEjqa2o3xf3v3rZOJjYDXECQwDcjGN
kFIGAL07RySn21umAM3WigkTfMhW3SmnpqoxRYpCJkWAPRCsy+ojeSbikTOwWyIh
KCy/n4fuwqq9kVP4qvEQuaS3kMHHNQm/BU/xHoME0Si0ChPXZAnRSP81XL6lG3vB
gv9MLxoB2DLkd66gKfKSdRndiD3X8IueCTFqkkdvaf/FMTbR8C3NQYH5fGr17sbS
1KxLXcbi68eKaJLRBT4TC5alMQquGoOXxWvG/eSIdZMTAvoC5LYTKeQOpEw/qpcG
VUhgbef1lVNZQcELlX6OeKntaoyQ0iAM8vnDPr+Kr9YilwP3veEe9Txi6wTAipFj
sZ2lO+C7y7J90tcM0TLcsd6QA8s2cdTtGMyvXJaXMi0FPp9GNASrEY32/auDkAMe
AUQkAMv2eruaYruk++DlHpH6AifJ0m+/mq0RMI0HzY/1tMZ87Cy4HanBCYsBnVCF
k82znErQ898Ezkkma3D8IFnUBLq1515OBdwojEHkF6yMM3dYpE5JPZiHsrtZoqlu
FoacAB/OT+jb8KA4kJROwl+3gb+SRYr9GaYujleze3BiF46ZkDGAlKyVwkbdY7hZ
KmkawUc7pUuIbr3FMGU7xde1pd/UH4D50/rvQIp745yFnOJ1MxcvtkIDjTDzTnEn
vlC3hgjNwLF3c3Lxb4zlC2kQ0Jc/NR5vwoE7cTz062Os9WcTl6CVXtqlmVtQXAFr
1LIvyDYApj9ieaWoqRs41Cy4/mQcEWv7V3ngI31CY/xQb++qca5hdJsG7ozliH95
OrDlRzd59RAD3BW2Wttrqt230cfcWP5HFIvrBlP6etfn95pWboAPRNLz7f7gYv6K
Wr0PtE2Mt7D56Z3HAipKf3bOwcO076lVFUi09d6POA3F0bYV/Orwvjuj6kngppYY
I8CbQ6DvqnBQrzx/N0jp6yKdR8MRQ/aixZrSNrLSKA9Busxtg9dG3mK7ArZg5HS+
c6txub+piqQV8xahdMIwcihzzNa182SuHYx990jxOo8ZsLSfqveV8rpbSBA1KrR+
ZRVGCxAwQGUbjMEariAjDPeAkB3buVmGyem7yvBXT8Q1E0oe5V7HCIJWwPTWDotX
BBT0uQ/+i6cS0Y5KIJ9Rg7AeobkIYOngJ0qp6dzHsAyuTwTPqEAw96uWkaGMpRHg
ej8XFTU+2ZC72qHdY/9alRMvs95VHhZpNTmtK/gaFJtHbT4T9B+VpEapLe64oU0M
lLBt9NMghITXTYKxxtwNeCuIVbE8XDZEf4SyurPvURJ2lUlFdP69NvqOz9xzygYL
+DkzalmTLWmkCof4BMEUDApWMouUAAemdhMYjRNcfsSF+viiVqBCStcNchsOZJLN
Kf2McDG8NiyYImsda5R3Ld0a4ZrgkSY/qFDkd/1MFxxSOHCRd6w0ScrYTNoIakmv
0kRFXXy7+miv8EFdUb28+Qpl/PEG1nWhu/zWzkDHJuII2snO6qXEjKDDkrl9i4Fi
h0v21JmBAa0MSwNIdIK8wrm+42hOIqvwHt5jc9/o6kIjYb/7ciR2gjjzkvMpmWK/
rzq7oJ2L44bb+CByjkZE9FDLtA3kJ9w5wM6MYd05o0ohsgZLMIPdk+YR6YuE2qom
Ggl1A//oVIrA742zEYMChiJZzYgmlc6IN1Hz8Z53l4Nu6kH8X3pTUYJ1EzK1A/xu
H9EGFXE8L7F2nmR6VCB0XODAvZSE612LwH9JTUx3spPEMQuM+UA7aisTsPh+NZAD
70ZGwR/Kv9bAPb3Sup4ckduVuBNZakveuc2bfMySg5QmHboi9rlg2zmYCG4X+fC8
kQ4viIqpra2VOz13EN5cAV5f1jL/z7RD86lbXHh+G6OzBvgjDXc5T2e37i+scYIW
HCGbJuRbGRh9YyeA94ylRPpDOFvu3xUUMEWFGMmZTU1hqlQxEM+V82UeiJVxwRFu
LasparDJpvu1gAmzjAxF8qcVIrScgKv+1KcTeP06pDr8GebDkj1KUTUOC8ltLxfO
sB0gtqIuDJLwM2LJCdoLAbAucdlmiImTtaGNUKlTOZzyoaYQBsEPxAFDlYwfNs9l
ma85XiwJ9A82x9j3bcFkIXuAimFqZtTne5Ayvtruz9MtIB1Z5/dh5Ih7LSRAyHN0
eCIxdnstKs4wrTHgIgtf5NcqM2OfGDp2cOFhqMvZnPvq+kcio0N8/4A6QHlSteWt
GAXrOVB1/4PpZiq90dLXytGYBKOf1u9sKOHypNN5kDbw9kol4aUTGjMUcRQORxW7
NVgxPcC3Ft6DoehhHvA45qSKk1hQe0KSZmClm/FIy05gSPde6iHr8UG3+o4aPlc0
2UTJBqRtxKvxFlj5FGdBRG1sO/3mXFpDXfww0buSuUpWkPB4sTtgNqFcggTiJ3kv
zmxZIMTwro9+Eii23L61JdjfoPgIyOubKKEDwiGX09tWlcrS3AiqMhP1DZkfbr7F
Z3Jlr337hSG6H7/4maGq4awqr2nXzv4yfy87NckM3ncPXt32X0fEHKawUF+AeI63
1UGuJMJF4d+Ul4y/Z/m7yJIDhsxmE2K682PFZftV4Q2dJprH5zRJI77ysb+0sEMK
Y9sZv+NMVnYv9QrJUUucNKQaFGCYe+8eRnMJLHKyKZCAFmy7xh9fswnKVK60zD2+
esMVlNl+i65UmpHI4WYjgOlyRl7+3sTYRlAnG5K+4DiWXePYvbqChjHYM3T7Tpor
pVhCUrnxHqcoVjQtW5pm+QOqmsO1FT7jDuu05NM27kzSPE7YF/kBzp0aZ40Pp7V+
uN1Q2n4ZkUFn9Aj60viuTBXBtzYDT1UCBvOiJJG3elwKylUqaIBSadMxZ9xMbDU3
vfXNd5OpGY8rYPCPainptSb83Ygcx88jBLhBMdprI5O3tprOs4GmqoobKKPu9ljw
7Qg9Z+G428A9MaizZsh3jUxlpwXDski5fKwujfEIbvwM5z5i6tcVGgGokIf8HfMw
Rfo593BcNb1IxPf5Ia06yitTjDcAFgSSUJHNrf4FO1mZNuOWsRkjkJLF+7iSrAwK
9De7zeyKGhmwl8ifNHDSfypREHwPQblbYmikdRNZ5Klc6rMgjnO3Yox7KCiBQUVn
xANxSluDY/o3tFXFwsFl07zRuvujPaxRku3glBvaFsLhw9uQLKznBeNZAZtwrI7C
AsdbD10CR7W6+YvWnDy/KNDMKpwwFwUPTEFczmAgrdvqqRbvIFeS6JJbt5nSXEcg
L7Vj3d4g+oOyjKQoaTkl3GmrgTKQNqPhsQP01haK9BXypFWksoOiOqjhMZl3VpWG
BocFFCfdGzaQYNJKX6xNrfpMjbs6/L/4JlBr7gV9v/DJQEPrH6OgHlYUGQMd4NRn
CwQRGuFVqQXbqHsW/CZLNK2kdyZVvyXdGo6H4UVYlQnbI2lpapr10pfG2QVCBgUE
m5vbJ8gkgLfixiZNFkdZb1sLfrtQk2u6c5CKNTWjFKradM+MDcuB4MeFoQkf6Umo
FeDGJ/M8FqINEBZ62oeWJHVeKAvbuTcM1DQN57aI1BMSJEG7PODLpVf5BqcHGDkC
ItWq3tqICIuHVU0EyhAnNblA4QViZ6ewtNHnYiAqMkKv2PhfCoK5uYLnXfWfMIkm
RQRQ3ogkw9VVPhEewdVnOGcGRIXiDSzBtaOTVgWhNSFHRH7QJ7Q8WEss5CO1BnW9
3FYU4OI0C2SpzvWolaMuvgblZHIP2I/5UxQWc3IfJF14Eektm0WuHd1eW+R1Tdho
baYsqhh75mReVqSak3Wfkkyqcqy/iaqH387hKIxdFXZpwIHNb0a8wqcWYmjaWzHd
zvyVHWI4JVslmPixpMIlSKdYxXvyI7llRMaApmJ/ihPD/o/QvSXFLlQyAEcHwC2j
QAPygeJBBEfjhBxWxponWaQxjxS4qL5onw6L+s83d70zm8e4ZqMtfK1AkziNp/2g
vGCei3fQ8vZci6vA9LYM+xQTDwtN6PgH7VgFyaCpf8Kvff3Q54BHMh3dlUuh6EPP
TuR9L/UIqSaF+XItIDmE1id6nHNmcfaAysuslKHqyUgKhcjUbCr4Tfu4a4baGfEH
5f0n7TEFONSX4DE7ZqL9h8WVsQjAvF6kV7F65N4MttikdgZ7q3QTmCUKMVLwpmJX
3FIlcAq/SaEp0hiQlx+nsOxpBGSh3dKboxV4xuzOWXnwalbxLvnFbyf/vsjhUguX
nlitNIt7IxfCFp7xdVRmK4ygspJnn6328Z/TLJ/IkgdIAAIHHoPHN/0UL3+AvrMh
JAjHUHrtnh/LKs9dkH817PsSjBCym514G9bHmLo+1iUHdyciVEjeYF9bcy1q6zXY
QD0Y2m19x9fCFGK7+iYU8JxNPzoLgIVCOtW73tFFEMWeFYljeXArEKjsCfxiyf0z
XKZDerRUF5doC3/yshVVZX7KbjTZNjmMzXzrdiSDQG5qsuDhBMGU9wJ8Qo7aj0gd
Oau7YUfi6At+smesoH/0FZOAoLqUbuV6bmmflYmSlNXPLsH+BbRscgg42AQ3VZ5g
+fVofWnUgIWkMWsrCyf0qqyiKPVM0oxCuOgwsQKu38ZMo0q1eA8wsfVjK5BLxp9K
o978bZ8kkLXEW0XJbp1yh/CbprR82kOGBblpblLehEVXBAmp1Q0DLisOBEK2b0bX
5Wt259+BJZJslokzALd6MdH2rtMGhk0LsYpW2tZM9mCcVeBU+p6G6P8drOvw5JYJ
IWUfPIRmVm2ZhNJKUwaSuBirv8QKcbfeqqR8+EsXl9KdSmALlezxqrX+Hu6So9WC
Ifcn2qdV7cLaZiyAQRPE5ilo3btM7LTA5JWXXY89i5Zs8sizXF+C9Dq5bxawJHy0
fQFSuYqoG0iHHXbxMlNAGUcKpEhQvR2+ix2xJfLYHWX4IGFjRwvy3Wt0FZQ3f/Mc
mnoVdiFqHVTbMAbvIqH6pXbIhp8B8KKw3Z58hfiZyVs6/qdrwFj/yZorcXDDE0ZT
35CfT6bMLpg+B/WAbPeMB98cSu+zBDyGAA6bgk/MQVueH+mVt9HMUhHhI1omuD9Y
hnTI/RY935J3WLOqto73aXh58b+W8R+egTsheWneH7fYZpy7q5Mw+81HPqqD2MKl
6iClsYjnfIVR/34/1AJ6HqieFrk6GLmKjEEKYVphEZUQHFSaaSMYlfwwMZNUPhjH
D4iBlEhNpjzjfy1MW8OJFms5mIDNPaxf/GBumdS65NVvcFZWE7NSQL230z7BhD4w
94pAQWuxWe3dXHcYNO6iPXglDQRxzLSyl/lTRreEMa7QuwCvLOPaVbDvzef4PI0R
CbGzfcMdYNMqHTxK9UDc4pBQXw08eCbR8LpIIBUuljgfCM0KIotPy0UqEnvUnc2F
COM2ycm/iLEPaBj+FdJDYlVGImhdCXpW9vyJsgdkMaUy8VNBWLbhsIUhxKPDyXvN
Xfe9g8g1g0Itu81tiFpdrrUyb9OVcjOHZkd2iWrohUC7vn5ujiwZoijKTI1Mx64x
mZGVPlcqAvJaqqPIQkF5H78qlLaMxdd4L71PG3VCvL9r0zO9muIMlsR/ZAV9fhIR
0vSTlGsTihktDRkslWjLgBFVzThkOIgFoCBi2Ezr5LqyBlkTAiMiV+j7BRcPxWRs
4+Ftp6A7LWDARjOOO8826Ja26lh/EkZnz4lg3JY6Sg2PoIYRB1IfI1dQq3+rY5/a
zGJpq44JHMtXUJzrXDGYovmOLq7ndmU39sNYiDlNgKlswmgT1+NtnU4XTIRxuyzr
xRj5eh73ljojnz64ttNLPuW3pOWItauoqul7t+W7JJSQdFJ1fkBtcO/EAXqudeWO
VWv0NZtXXbzqOpE72taDn2ieW8mW4LocgTkcqd36udQWC/RYmXcWYKNv4HaHhxHe
ouHSWLs1+4tmtjnvGDPh1cloNKS/ye3V5F3GqIrWhD2lc+OJKTxBQTUc0/yyA500
quPqxAPeDzSOiFPEZi4cArYs6Xzg0VKxsfZX2xjnC8sdNioeLkMit+b02xGiryDv
b9LWR+j2AuUkvZhhFLii+Re6bR4nYXmuitkQBrIcxiUVx8nbzkJ+tKN+G3/o/2q0
ExBNb8m4/DO9rUmJxe9tRNhDaUA1z9FLGbvoaOyZ8ShdF7CovdoTn6jFAgBLs0OT
ROvmg/I+JoFUcCA2+m0MqWsQwCSp2k0hH7OH6uKiJgJAoq4oVrwPihN4KOF+NleA
XzXKnt5zbD+Bel6dgRr54tb3S5qBXk3+rLlWreHc4SRS9QusFQCUWKJntedpcR1D
LtXrx21BNL5TblnySUo57G7Mdux7aVWweqxjZBBQt4JmaQdxD3PQBg5wKhPrKltD
RazvPRuyUWIX+lIEdfHB8b8bWOtlXbmr+albSW+TDVaRrQQpV4bFI1fsYTCJ+aEQ
+OjFAwkHT/C9qj+JCh+wUmPmJ8fpLqKI7AYjYiKef1ne5e9GNWORBs4pd0xDZeUi
oQ6/GKVm6/I4zORIkXWCbcqRrgdSJDOOeh8RArjPIeG+erzZMinRAT2m9Lz7D6Fb
t2hMeIl9keIhC3si23Liz5x+m5ubJSvUR/VEwyD2ac4zcY/t4ZO4nC4vugoof4su
LmtClfacAN9Trpla+BmFH/ohRLf02SO3TAlO4IIe1An8MYmX017oJeksu4tG/fs1
EFemd1RXhLRjpUfyISFZHEhwT3v2E3mv+oXgr45YRG1FFUOg8H3/1LFDC6WFAtmI
RPREX85EETM6ydGVt/M4TBkurPzXlLcQPTS0kBvFKtaTiR9DcBXsTMmEaf6O1jgK
2eGgx/VGyCw3QulYyXMf41BVrZvknDROpqUDMj0yYl4wcZqrfjPGYHkn24YlpYKm
MCDh6zfsdUiaUKibyqFRLDOjCtwOihmZz21KLSYlNObsB+RS8kMpQP2T7vB1sDig
Q9EeeW78/loLPVpLtNNk8DvnvMqBZJIEqJOS4XYvtIaBbBZe0OcsytPqC60ejie6
Lqzoh0NvXpuo0uQ1hzzxfMNt3cO+TRXaKOx1uamD6epBYLJ0XvP8m80BaRGKcDAf
FveC1P6wBy0LkewoS9ZcjNsRhT4phil3ri3cBFd7I31IenEaqp+Byv1lpxvkVTKL
4PzE5WH4xgseSzK0UxnhiaSaf/SoMDrpJD6A4UhlCQyN6u4Wc2UgAFYmd+36X47A
wsbn6ejXCsQlGzisJjavC7rjLd4gVuPYad7fY0jlQXasQR5Bj0eW1kw8WVKC+KK7
20A3amILHhdcOA4veF9muEjX6O9n+hakIguRNF6A1iAkEwLaTVETbjRDgNhsJxj/
QW7YhbH9ARKND2Jn3sX/l16EM4IeUnqaeZyDlPOJ62Higb4oP+E0uJEgnu0y4AOd
rA3p1fYHkBHKhUDKwkHFYn0IyQ9FK+HmtGUWSzgOExtFJ8foCP61soXGBcWlfpbT
jYNT+KWjL5+M5osX1sZ3BWoW94UDjbFMmMao3QvspdVZ7Dg4M9NnH/2ONYqwHZWl
0Af6fjEov3p1QxseSJbd/WyHyMuRAryEVlTn3SE58DxByIH80jdnSI2n/ZiEUyom
yUaLsHvDdZuIskcoG3+qJcxjIbxuwALjXU9jcFVeWZVgW304UbkC4Ojw6xz1RqPL
dxTCqcFqI9PFd+v/+AJWN9UOfMkm7xyAQhywhhw5lcdc+DMo81ZY8HEfBU3auLdZ
2eQ3yRpHCE81ewSF1jMgQV20BNCiuerUUxwHX2xLG5DY0vgoX+YIN+tBsLsyX4mn
O1WthbsMeXy3neSwVdvDPKu4w4UiiMUqqdVT2DCfZf2TCzhuBaPGbrli00qyWtgl
UeL461iIsCH6ubXJ6WZ0RU8zwEUjymTRdUylBSBhTolm0k3Z3WaIAxlvUix7v1mE
ma/PxLt4PwWCTWCfYO0YyFeucrOajltuovDZTBq4fq4S3K2IZi6sLqfXXCgVk5dI
p1+3zpda/O7mVWsH5U0mE93djYG3j8L5EtfCPnN6fKBNRAoWDk3cMKMV9bHnHxxB
f4zXe6nN+zIL9Ek9dl38b8bThLVOSCXLnJJkrm6uEJTK6N2zG6rvmR1aJ7vdWocY
JERQrDkQhWJ+l8+AruASYA==
//pragma protect end_data_block
//pragma protect digest_block
u/pDl9RV0jcsHoJ+sQqlnKpZ1LA=
//pragma protect end_digest_block
//pragma protect end_protected
