// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
0K/PsuqqzeKqbFbysjjwBtHHRLopEmc8tCGskq/9u691UDXHHWdKJ2kajLerx3L2
PeX5BapZa3pcUIHQArwbnbBOB73GPD/i0anYSk7NYUEMT4P/FnTpb0ajcNs844qA
Xb0kt1JgtW6L8TBuCOX754mOqXwL2OcdMeV9Nozvz8nIqXTa8H6J5A==
//pragma protect end_key_block
//pragma protect digest_block
oHGB5KSIlfGlXysqmJ5Ct8cMhoA=
//pragma protect end_digest_block
//pragma protect data_block
0YvGcBP/annjllZ4V9FeNdfdsWKUOEgEZ0b10VJikOwr6czM5Ahp0ssYHGltWguE
NokZzWt+lFUKR7s1jzh+vI6YmsqBM9slggaM362qiVYz75/zNQl56iVWfkttwx8R
pxBfyFPZN6E71HqmzBi0tdtpcSBQx6cD8U8kq7SGsc8XOOSqA3pGDkxFw9HVYx5U
Pp5w3c2FJ7s06TY27Megyz/xzv0FXb8lUPyr50g+oXJURi2n54gJCjp4Tu14hnwh
iTdWNEw0ppw+12ZneqIITVBIX7DnVIdSnmB8MGGQZmxPEGos/g1uepEvEZFeFKyP
3mcwLluCCJJTWxPSEyYhWNJrrq7YFus5rOT9WyagnVGb5m2VR1oXrsEqcYoetvDq
wkmV81v/vqJnbWatx3AdDMNxsISRWQurpzaFNYZL0iq0tawN5ufF481oAGFnmbK/
tH43YE6sNBbBotI7Mo8KWZExabQQMYW7g9yltWgU7BK8bAEqsQkrMnT+q4ZzNAcg
ZMtpw1O6mKVdwQqHXZaHpWRNHdYruKjjMYzY/TIN+Oj1oH49V5M/6/VHGjZphlxE
fyp+IvrCD0X7zsthJPQPDINTFEpUYt+/uZ+rbrherBaGIQ55VcqubZnq74upejwI
5AOfD9fhoBXe3k/a800tYvWeBDkbVxIeMXAZEPAXbitotZkFZYR0PDfmMgb45zSM
DuKtLjAjBB5zOgcy2mMb6GDkfnt3B8cmVREcwK+VF11EzaheOjiyLsdsTquYrs3U
UDRLsO1jixmHETFJ7xVtcQ7Jv/Jghspmezib8g9OrPJCsZEb/iM0G7nfgA2g9qSk
P/HUwKsxkSbKfIPYyB/6FW070jRwWy/vy1uI5xz6Ss02bKxzm3AIK24WoTlQ4bX8
moYylD/j7/wBMYuuk4tjU2nJk5U60MxNJ7sJB5l1Jel+nJ0uCd1vc41tJr3xT05J
gkHwOD+BgO/CWdynrhP6GEuvQHor/uGVwNnXoh3J8efB5sk8GervWzBMUlKgqD73
icWFys8UHIFo2FeK+I5p9DsPEQC3ajYN4D3Oh1/lrcpSWiYu9AP228jQw+nHnGw/
0XAN0MopJ34gS5Gnf0cQXW8nqSAPhrEMREHguSNcU/HbLWYJhDP32dk0YvWBpDPF
JUnARTPWhHgJv+Fkhe42498qYeI3riXpjRL+Y3Q1rE/GMD7sh8EDys1DHkL4S+NB
o81zOqD3bQWNdnpdj1PCk0u/k1jwM79bh9OFF6K+1u5+uvEiynSfy4uk+jvgIr/F
riyxOzl6+B8SeZcrcotJtfvEH/Z4QkI6PABnzuxnHpRW7ALT+MoZ7UDcUhI9aFpo
U4nQkrjyjTlPqXI3LPKL8Ss5T2aOfhE+Te0PoWwye0j26pfoLXvHCu6v/yQwnKQA
c8vjL8Gc5JgChkDoajXQ3teK2rPRTAYJsdtGQ5FDaFxUDl8+0wHUuvhPdw6BZyDV
63rR33n9wXc/YFdk3jWyNZ3s98JCqceav60PcMDD2Qj7h88PCxzxyjciwEc5TqH9
AxAVSGw7g+Muxvbnmufjds/7bdg3iL4OFT1k2vphB8J8JaGaE9+/rmcGiLQD2+dR
PIs3RljfPGiDT3gIlnJCwwpDzeDeGewtu7vuxEh34CtZAQSHquViprLw3g/9O9au
bXdvCZ8sXpkf0b23VsxPh/mg2lXbl1iDDqf3BvL8yNa6qZOrM+zGUxUftj3AZVaJ
yUeTdMc4AgKxOjsseCB45TqPpt1ddiHY8fii8rph+T6lQ7C2r59Vn3wK0giA2sgb
bBACxewx0oMIcjFvYFGpRR8FsFlwyJPekEulKxZojy4QwgE2OMr7lJgfiYW3zLbm
a+6CNATcwnGFShokYhT4koSPXbbYU8Tdcmib6AwQgHpi/ZmxxtRPWr5wjx3IVR34
yO1t9IqLSCCyW57hCv+9rpbcXFmvtGMIeX9q6J193AaOMsWq//fw4eu4nsQW+UFQ
Y0d36CItbRNrSy/6RdfLnW1jem8mVN0HD417QrulzUqZz1Rw4gCC4H70G1vjAQE7
hTJJh7oGveSJZPWF/7SJ31EgZkMEKAGhmai5GF2RI8GvJXX6Rn+LjAc4vdxkn5Ga
nHCDTE0L125dioPH0z31w4iXeOCR7QGTqcvXRdCU6A0N3CskLn5Q7Stz7b7WThM5
xesCFNbErd+gN7tJJprNeBTNLL+cCZvcHB69v2XIJivfUNFnxfdPnml6r5Z7sD25
idYJc8EW22WhI52Z5xmx0+OdHrlqYyPL/e9U2mY0MEDs9xOiNJn5pYfQnj6hUMqD
yxaaUcAuyCyG/W+t9Ph6a4YA+qslF0VKpnw5R5JOCZxZ6a++40ekhUCUFyc7oj56
zf604H+7Wnh65LBkb4DtBKm6hWJ+JsYM9mqBIpSLOAkBASH8cDnFfxZUiQIAe9hQ
G/ki2oJ1SkhL9mUMoio8c9EoUOjtcTVMweSYuntUB5jRRuMrl274QsMl/QSGnlmc
4VrnqsDVcujRUFXnESujIzOKsaJgHX9/yPAetV2yCvwIkNPEG0mwuqYIFnMHrEhT
oEt6Tk1t5sfqeNPnQi3MRWKhOd8n32T3DqjvLk2r4r7I3P3k/32kmfJB1VvLJcDr
CIXkffln2KiAV7zrtCLo1DwVmYG8e3/I1fXX5+QoFqWE5a41Cx3wR5I2cTwt838I
irsD8s5XnkIwetMuQbmxccynlrQpJE+kfb8BVR4TIqCrrYoKditxTQHxhKXmEwIO
iCqECwR+s9OjArvw9U2Cz5IMVL9SYARqA4czCXtBqpoSQjsk7AqhdH2ZxpZIjeuM
mRmSV8qhW7zcT0FpdcNplGA28O70wmH0vzj59vD3ui90+rCQ5FucMe10y6tc7BKy
zcrz1XZl30/Q03ZX6UFNcSThlqK3l/e1ZcWtscucS3McO2w0+N+iqjXuMWr6jOpA
vgzu03Ok1ILNZoQtrxGHJ1GkVwGUq1J7u7V1NJTPskn4lQg8y4fsSjSjtI1s6l0y
7lvQ95CqS6fb8nZj28Ea4lVKHOk24jUYAch2tTys6YShC1127WkZCyfHTJziWpSg
4v8mbDyECxNa20R9lev3+qyHubqfAe0kyy2Gz6JLYShBy4QweER5UhuyGQwEyfgM
ehDq//zDzXM2xgCS24m+w7/p8w0eDjPVmX9M+EeIrO0GFqlf7TxYmjy8JyKpA4N8
ajjFidl7jWO1uk6r8d/ehGYkZLJtwUgxGYe3hTLaCLLYdeRUWPNQQQvuYUyvvYNo
4VAbukCnY4jg64LihgEzd+QMIbHriQfEf16uWcv33xMpC5qHlq1fsLOV+9dFRu5L
fklRaH1dKl264oaB7EzxluFLalFdf/8bSQ3rGNHlBz4rUgyZ6RPXBZotVJ1KTSkb
a4xHREytz5WDXAD9IfmYiBlkoMBg60IsMSR2z2+8BmWJ11QblBolCJPMGSig4LXO
FE+ZFrjLAa/JVJXn7q7OwLKg3h3kvsKt2CanXjxhz3q2Efi5Ggw2oSPtERmNTYLC
T7eNsJQzfw0poOusxdRIdT7EKNdQ9Mrt6BPTC2V7kSGol0kK5tbX+KfMvVxMHj+O
NjBBkeW5krqewwV/eRC5bFmlUJuqU0Z5cdruWc6wtn4cRuV/BclUUIuGmf6aLXz0
eO0egQ6l8luMAUz84ZnCAK8Gu69GAy2d5731Mecn+TAV4Lixj0X4TfLvpVOBLmQd
iFcsmg77H9OdLE06KWSeWsSBFikQ+BzpEmMyTIKprfT0e/DK1euqpbklGSZ+D8Ru
1/QdhoTeUcu9+l6P9KFcQMf2ifPmPeTs+VkvqCNQPq69Op9ufx/RoR9bkm2Y04w+
JdHqUOTx0DRUkkGx5gxsjJIJczJoq5+TkPgWmRKGc0RlHYZLuuO6WYCye+hat2iA
DWEZhsz3bU7oHozx+UFkiwBU70lQDmOVM+vYBDBZreurmRPnXESF+faN626lkDK2
WPzUrl3jonyxAudeLcbBq8umPYm8jxXgp4jeJ21Lh/0+qTEgkHoOquXBzShlmTzc
rDXk7JslOoECy6cLM2L/gBziuwas+9ZM/77OmKAOcwggY8TIBUK0ZTQ7KRRASCRh
Fg/YlWfn7qw+79qH3hqw0aEDfelR4TIN5mEqQynVoN7OpGyDwqZL92fQiID0s9wl
wLOV+mGhY/MCX8xWVPcJOvqTpRPFfhWNo2kBKRF77AkXthG9A97ohU5vBN8YY5DO
4HVI8H0k+bWxJUYLi4xQkAOLAI+fBni10ASo8I3VI6HWOuyEf/1xZIVlqk+wCyYy
0C4zOx17/fMQJjyb7So1dwaqQ90cZ1dnRpmgVeILGOWAUreg4xDqOv5hjHaDnTzv
jBoh01SkqzNp7IN7VbVTvgOTVpKOEd0ikyaC7Wed36Ny0rVed84vNa8IWq+MKzqw
w1TejZn7FmqSEW/fZ7XVMgwr2V9PJlPTcs9epHDBEx0R7HZz0Jgim3N221ZiUl80
YY2emaOWV36W5W3nfqoNtSEJrV15I8FqO/dcSuHK8XTL2D2w+XTAS6a+NhxpWmJf
RyWurfmAjhdn7dvV+X70myZpY75hoH1PeUgzn71ZM89u5P1lzapiNV9OcsPBrl8J
HDPwTvo+kGHUqShunFkio5XhDjCpNQpncURs0RIsIi9nanoNa+gmVVTbvBFWM+Vo
VR5uU0WBGAfKBtH23C+/cF+PoyB7VJdWK4dy+adFGGVplK95WrWAZAb2+FMnecRR
LoYh5pD7mATf1OHbHm1IFMzfU7+RWnvjKuyj+8CuA0W3s/M4vHLVsOo2S5fbroFc
JaP5VLeVISszg2gQOfDbdlcXAlt4/3b7dYsJGPpKtyK6bkJNFKGHSZAtzp/bpMQX
S3KAxtF7e+mTK0npKjfNDvIgoQKP8Qfv6QU7Hl/Kec5MI0QdAIgt0cglbBgCJskx
V1iyokH92VBpY0X2vHMxk8m8ls8jsI8mfmXUyWJt4eA4Arh2puPRlWv42T2/f2FN
kU2edhv6BoyqERIGqzuwN2vJpTLVktGRsOLP/rf2Rrs56MRoJxCdDR/TuQjj3yWp
IbHZ0+VNN9shIDe2HL9AkQNnixNgxuXh83tZ1JPDbIBoAmMI8DaD5Jkz0QRNEYMG
Aki8c0gMfb3711JZA9fKJbuUUbki42zMi0djIQU//6jVwkAbcjdrWQlnhyyi4iwk
NgoSN5IEXSIGkxsbHuXboS3RfhzbyyeemBPuBcN2nUbCV/bxGScIDZ4ivfQyGvQ6
akHXwRbMZw8PdWvkF4HI07l2oiUF2nNDVgX5xrvDhv1+PpA7hYeaM6iWcDnv+OoB
iLt1+KA3GxAAmiXVPCVyolLm5hJoIyQFtMF1r3iYpFz2RkTOZEUNdpE91Nnk/yRI
JCCbYsIjGcv4+sW/J7WgSgsSoLUq+2r9qUEWff2yEmDOvJDbGnjAgx8pECsSScNv
rR/PJhk6PayitM2z660VSFjFCYo4X8PtNwCiJjWbyVOoZDGUFxdB2nXaIe7nmXg5
zUXjKagFiMCsYjvWbSALAHAYgRD4OWUV25r8kIBvBvK4JOx3DXiUMpN3JRpP+EnF
XWcOKcAETO7GiRPV6EKRnwpo+/J6odG8e7zUUz8OjrtlaUq9FOFK99347OqFf8TQ
3LDDB6Ui1zU+pqUnSf5q08hsI0q5D1NZhkaUY4JbaQIregR3ZqzbELM2FFFpb5RH
4gF/X3WdJ+mCJUid7CiUhrofiW5wqEx0OkPtgTAq1yJiRw073JswN+wJdsoYktF6
19Q0Lm8obel76oDWDe4dDbFVkh0MZtfHCmZUVWXN76aywBQHonFNIPzxOB1mCH8r
65fezOchEBxrhUX8yC6TFNLWNmCoiYsVFe0PJuOk+HGQG4AesmmucGT/wF7LACSl
1lgGjMIMRIxZFWKBN2/0wqOXfaJrLX7VoO7iXD3bVKzwbwrBua5QEvzrmpB3elbg
trsOahHKtB4ilGsKNiX7nzid/TVcWoqLbHjFCqafLhPiuN8pi8r5evUVnOJFpD+C
eAXvVpc4W3H+ydaGm4BdlsHewWOpnQnaJGvnj5b6GPUMMz+S35KbJZVZyoW14MtQ
/DC5C1liToTMxS9znTe6D17zSgijZ5MBmiUgKPMH/lvvtTCxg0MTld3VF4ejvp1I
rE576hO+v4fK07pufsofbYwVy2ErfZKJn3qkAf4dF6Gf5H08wjW2UlVAQHq0xWMS
e+X5tiZemlP0IEBAUj6F/LJbSLVuRhhjLuEXGcfL81ylX8xD/DYyNpa0y0EZs2TM
clyAlJy39yMJUEMqQkCsjPW8el8XwAy+3FnP462rQn5wjVktS4DADRnvihGkd/Oz
/7tqzV72gUjQzxeZJaXjdqEXi6M1PaPvh58jnT8H9lJoU7T+KilZMqpBrpHhddqX
o7j/vdpPiaDsTRIRcWgmlAOHB832rrx/ak9KX9Vk9kEtzRzU3z4BoVflC6+aF7pl
m4hACJI2R0uOsKfBTqd4p866gtsx5crz1iIxV7dFMiY/zd968ecTrc30TyFLyMo9
4jiucKQq6QVfXkLLE8gRyzUhu4xz2Dqp5RL94DYIBJRH0rpTWAUI4kVRcdfAp41+
GliTNxiKKbuo0D3B77r/OhLzmg3LS5n9lsMJWTNyMi6Gm7wz6Gvn1c+9dCqatiXH
OrX1MwcztK2cKsERzSRhtg/GRvKynvLJtRmkp/Ny+aWAlsq2+3mMIyEzqUjVpzTY
PESyq5NLV+NCvmbbxBCoG7plLSuNStnTQoi3lVrwxZ1EsltQM5qBiTHjVhALJ0TR
ORP7qplk5pYPsynrCNDecLOiH1XzvP/CmHUlkEcj/ZBFVoLnT63aUba7JOYo/5Qt
XilzQNQnV3DWegIDjFQ10epq6cFFOVU1gS5p02V5cpaRXvJbLnC1MpqJE1M21rPx
dD8GI+W0F1GbNzr0aXSH8+AIcskQuYE26DXXJgUnCaUPZI2zByOrYkMzqWhdMZpg
/BlhvQJn4Dy0hSHLKufXb3m+0sbxibAXvmQM2iiNh+U3Sb+oyRrLmBdwDwWWhe3H
sBmCDV6y3IVx/8at6iDp+H/Ua1zVHWZVOZeVqbKQpoowtLBAC0D3HauOj33eD7vu
qLRSMEtPnjTX4N1uc+wQQXWd6cAzTf5djNHgajwVPFuvkdrTPqNpTNT/ZiJvAbYd
IKWetHIHmlXh0diyvEC5edv3mrSjIzgqi7UTnu2n8de0vYTcWDSE7jsaudYSafiZ
xk6xj0oswwNsWUNNAlaSd730kBRsouSTlALep6NyVo7ze8ZWIVhldDh09+OiERSb
jKRzLm2lu42vyA1+/ybqq8q6HOicp0W2gwvaRni6cJzjeRXHv8Y3ZdBbowgsx2ZO
+clz8pQc091sc2If+ih2czf4AQ/E5pf9+SiXcjHej3NGmYO1fBJDWhfUtV86jw9M
k4o9BI0Zuf62hPT4nV8AfdKtaWGv6pPbaPg3FrlpzOF+3lyimXihl0UGi4pvSvWM
z1YdDIIdBgRTxpr9umI9ZlyvUF3rxS+9VB+4MXeLlH+Gyw6DyWNZRgFs5nB74zQf
X6Ph44RANnKT4Yo11WIMknwT/Jd4CKTbGq2GLtbixbFda0RxN6WU8IqOWB269RAT
Uc6avC6KF2+kX0lU6g1yHbRTjFf2vqciuejacHJLDDJWDHdEsAdFPEsLV1BhI9pJ
2LS9+qIW6GTki6E/PjewjJFaM2ATutdDdcgYme2Jr6uLfPO/v7/xAX9aS5t0eRmQ
kU/AoomMVQUokLEllUNMrcDQavWf39R7O5UQBoWZuQ/AmSj8CpvO4wxLaJ3ke0rh
J4GjbBEoRdg2MB9xs/QaILzS8Ndqf8yCpS9lb7yGBuhrV+OnYwPpm7d/S/3UcjL2
qO9cSAsl+VTR/klwutFck6jwli4BPC2tGlt3rtkqDLB1+aVMuBt9UI7fRFlq6bmx
L/3mbrWj6z8pXf+JnTdFYP+4hpzrGZc/KnEOrfLAFLXQGjCMRTJcsp0UOfmUQgxc
QswnLzCDJgHiDGWzHj8euS+LIxQnRDkgLL1bqUFKH7d4HSlc56GioPOoKVHGEUs/
NeZjjOepu5mp6lB1mJy8e3QqsxmJ+kik29bdljjxKZEbzkQcyNLpyI2r3peHLxwa
EzvUHA53Fgp5KGT3Sok2mTh5XPL1oBv9REFZAGhodklJCIBpJVkgBkrny+1HX4YL
kzQR5xo6t/1EysXoPQdzPnUGwSvFlL1QwaqwFUIxCNN17gHCTyJKRVMrhJcz5h82
ITIfsoPuAKYlzfZ4ykDw4r9sWCv5ttnsBzKTZo2X+ewPYVf/UNj/JEKws0WIXtoX
HDWOm9O8iCd84NSbDfaj903/SFtcROGAuWfmcLr5k1RmLYVukc1JJSqA3x0ILlk8
NtevQEpa/Wq3to3CMN20Ua1Kxx5DMo0/UkzZsEVMzRtRLDFPAxFb3Ne59Thky3iz
CQzE30hmI0zRolTufXmVNcPo9q4pBlmLYQay+9xJYW/BeMMQWef/hM5Dq7TkMqVT
G+cl6b8RGxghYh6g1NIEMxS/pGRHuehpe8xCuZii9pTiSfHwKXL0tYke9xrdUFr8
WxefHdsgkbL729YY2DS21MmBva03aJvREsTdZPq3qePf1opyhMtNzvwvJ5L9qjEw
qrh/Tk7ANF0czHjXAR5HGqboGQLtj2TxZ+M0qEXyGJwv0QOwOftymLDPx1ByZfUa
BBKcta26jjoD8UnaUYckoBZmRLO2It2BM1bGZMhPFW/HMz5jHR+HgPQSQ1XPNxnp
pAyC7wdGjgrRZLAYmc8uv4lpgEWC2Rlhimtci/9MrEckuFlLTmviG5o6OPyNFEra
B8DFafe4IqFa2/tH0VZRfrRtBU16NHe7Qko0pUXX7BcDGcNgDtPa82qG7/YPCPGQ
3+L1W/dfshpz+wQX6411qwqZtbqxa+YQtvmwFZX2TvryiQULH02pUBQwhKZXPRak
QLkOf+Ne2WjgCNkKzVBlk0qtxDzdbhNHdYVjP7/hl403Ah+r+TyA+PIvhCnRYwDb
1W0tmLQciZYBkvPxIl8wUhqtmi0kDwmBIsSKmFykHTtmsvgk1Y+u4kpFvZJB3Lwx
hX2eV+iUhMBVyhO5nwGnUAKTCR6KKKBLvJzAi44l/aIVINUaOWve9znCRqFvTJG3
r9QiwMGfk0wiolG1BU3LvUy4w3lJCnsck8LnIdz7mDXL7cfg2yepusJOcmPQjhhp
9tits8kvoarx/eJwlBfem6XgEIYiuC8+6JJ4yetnWzac2VXXg01rfP1Xi37Suwcw
wkRKYnF1xFKILzftapw8ooAvDrUxqovgvkqDFVucky0VUg9eTFii4sQNFTdVlqOP
hnLxpSbG8wzRYE5Us3ntKPKpH1WBKWI3FvAbNbDBNJI2EaL/0aIY7LHETwiRHq6A
F1z7Cgd7Ie9+qFVuSHlgmXw4gFEw70AFwVfaK16jcTMiM/PuDwP40hTCojwgTXEy
wzKaR7loB1Mx9Ni379S4ggtHz7V3Ildkgjzo6epNyb2h9M8KQDVG6a35rPXf9Ezx
2efT8TII9CM1vlQy5C+qiGb4llsytcmOetjh8dCwYMFznWX7hNiCqDDV4YudOSTu
qCCV5MmciY1DU4drn1PJMn1N0b0zTQoE/KP+e0sYaxiwgYKe4Y//UOwJJL6yEDhW
EyxwMj7f0G7dDa+NftX4lx4i1q5aKpMVV2NHu6vq5u8+rvrDc7Z6Po1jpHekNp5h
COPSTVX8fGH+QN2bfRR4xLPh40OZL4Cuw/M+6vJO3nA+ZZZazcpA0gw7n7j7ufBy
okxybuyEOsKlBewoFN2iHUESpON1+42O1IeF1sSq/ok7q579ZdjMmJpxPH3hW0V3
A26w/9nKiJYT/l5p+ymWUj4Dv2h6pY+dHC7YR+ONtk4Uv8CihkCNldKiu8/y65ju
mkzXKhaWonyzkRU3MrMWOzTbysns05Hor1nYCn/b4Cu3oXhvSGcF7ssUz3q2ytz8
5aGn6bMgfT2TgVccz2QyMuTU6xt53MhjS8PE3xHM+N2RSiqtdANS/rrBXyp9iDsn
kgeXbUAqnh2kFy3WRoDLqup1JVYG8+wQK3AIAJsEP/j1Dl7VsyVPfMjTqexGI4RT
953JwEamP9Fbfrpnc5cYeG9a1nNYTe6X7w/duzcGom8OqgNVOUjTfaCIL0bl7DHg
IVk/aSb/uxY4969ZrfcSquQBuiRvb1nJ6A1GPzBfpzo8UEM6kkf1uYwpaHW1Fafx
VQTWwH3GSIqqnHgq82sxKvssEyWXhS2GqyVGe449KO7Nixis0vDlOvfLHapKp5ff
ye1cLfS/qrK/Kphy3kDbul9ndMstAPe4HK31FUZmJSGQfLcTGHhG9YqMLKwlYD1k
ugnwupOfZZVKoh4T6/jdv/98jMEQgNJ0naVQhxgShJgWpgimSlPMtdxngVngxvbo
7yTc72fyIXGIZq+WYUpYlX/k65/1uogxGCHdfv9+8rCSrM37Go4ifzgziiY9C6uN
C+PTWlXBSonQJYj20ogNBXIMbWSnwGUzk/hqsAidhIOFOdIyThCMxqycO44RVevO
EjaWcUy5zTRQSxb2khDUMXlOYKTuTqZ//8sTClNBvicsZLQnZpDbJKSv5zSAT8Sh
jtCjdAZW7UL9SZyOXyPhAYfS2uLbVKmay6AHgX7DMmDiSlekccuuv48ROfElz2f4
TFGGigZYhSx3LlBtoUfGUgjU51E3m8oEnjI84WZLGqX9ASsVoiKJ5BV2KshIGrkh
357QcwK+QuZNNQ9jbU7ecM2deHrehT0hRuwiLv1wqYOoVPtzqOwIYVNZSY9rRSpO
dc0JfO/+2qDSemG+/8GzG2WnukGC7S8dhIKXwyuoJyf7nibmzFi9S0CG+kkNcVyY
gG85mHKjAieByrjH914Ihuu7SqiUCYzP8eieZ8K2j7XOAW+BaGZ1C84WMVoOUn8e
l4M1QQfaUXP731rM9KVg2qKv4XDZy0wUDNjQczM3quQZfBh9MjWh17RCVySEUmRs
4idKikus1M3JCxJD/fkFST3kaEbzzqmtG9H+NOF36k4iJG2K4Rylb1jw9nhr5xNb
t6m/8IUVepzqPo1m6hf9NMOiAjQe8bRvSeRbzmLh9wN+91ofDbj7zxg1wiAUfygb
S9Fg1B+K3rWBYwHWB24iYXMmjvQmSpp/jtZ2K4YTvJVWv1w7PN0ZBrd8K27El1OX
ZoVUZ1OYIJ31nijtZRe42LJLFkcpxhK6GIp2SbQ2HWN3rrCM35EYZvjAXT7B9rI0
8kfKWnfFgSDPOfMf1odJiLBUWnA6avN+i4ryCUSyPBwuWgQBJLJs9rzH21R5wbJc
MvHSNlqDOxNMVwpDA7Amo823sukXywsxNJ5GJPV8CIt0nrNxJ5nwAb0JscaQ34za
p4OZ/q4vnM8uisvb2U6Jior9BETW/kZ642fdYf+L+Sxw2v4DemkcZ0kqkLpE3sBW
0JS1brJ5N67JoocG1GCUGelr2sLweq8+itiUW+Ax/zD9xLnuklRpSNvxkjyFRq2o
ZcILPiZ6O/gs0Hj/gmumHyyuAZdKR3T8R0iGDQnk2g6H4kE3HyUYZmNRmhQOlJmq
8iS+R0OXawgVheL5wMF/ssbggyJms6gZyPov3SRzIhUJkBT7es/OsaVU5GimDXD3
X5fOOUx481igsmdsSGJiUfMc0HTrcqo4zaPLtOB8d340v/m/wDnCJ+JZPvwFVL7d
/bOCTsm6vhAdAez6W71GHEEEb4UcOaLn8c6hQBxvCQEE3EiDA4EETSwqbI8RfmoM
Zlywc+5DVm1TTtrJlYajhR6Ckt5Bt2doWP8niUSw15aPpN7oBHRmUOrkziA7aOUP
W1furgxlH1vjatDB68+/TMbzIx8vE5dFccSHeiLPCeGIRAIgpU0QeJjX8UBNj5oI
Y4heJPxjq22YLHnd1BJnVk3aV2difX9fW52LcKmR6M5zO6YIX4PVJM5Y24jgBoot
2fgXAeqbvaQfZ1GDjNsQQ9VaoAP0tFrVKN92FgxtskxOvILAdNQx3zv1+XbnXfgr
NvjVv0VlPcu/Sar5H5HeZpq0mDOyUIaStCXKkfa63S41Q+L2E9c6iK52b3VmnjAu
oBwo330kYUGZ1yRdAWs5lb6Pm6yUxJfmATYzKrvlqWXZuqPR7C32XlyB2YcpOdox
V8pFITTiDPXnESesAcNPkpKN1wODKUOym0gP2zHjtL+rhG9ChoPac1qvX1bxmLON
6fBdzzFT3lmy3nqbsd8Uwkof0ewAfD9CUTN0zx0euLVcWcNRWk3mRKgLuUx8x3Ky
hBSm1z6ou8re5bbs6O0YP7ioC4QfEYmOc9oipW9fxZJH4EFX1+HgK4OuqMeW9NLx
bk5/DUZxNuczwgBYvmXTVqS7kCpNR7Bnp9bVF2rbpb+kzFtf+v7d0/L5AdQtM7PE
3BubaYFmGajSqwWn5/aZCdnIwJXUKTFvkh74rW18k/KRndtl/4ajrK79b7Z85SfL
z8nJhNRoRN340jPc7hBjZRjkH6btAheHlaZFJh6N+WROkfX4mhfXD9/l5Vtq0YFn
RuF8iY/s+PZ+K23akl7yziTFbcCHzcS7j8AoEkRUdDOeizARifgwjAOpz3mcuekb
2X7x0LKHVtfTO6HirHAT5mnXWXbqKuJUoRPLcvT6tBKC6Pu4rHXx75KafVvBl0ad
QZOSnsKSc8ul2xWtKPJAazb6vxMthy9P1dFJVedvpiHmqEfMmzTKY0leMNXeo8Ui
Gxxh25bBmWNP8pEpk8hDAVIe0LPVVGZHO6y8j3JQKREE3JfbTpcOtxJrtAaU/fw3
039vsJ78vAaA6tH2FscAr+59rRzOy1NPiNuuhmV9bbBQ2iR1oLlB3PKXG6pSBS0h
qn1OwZmZnbfjsXQSMrIYdpBFihUYn+J2B/qVm+o4CAHRrA+U1LdtMoyJEwid8OIx
78KCgv20SEwuDASGvRBgt2M4csjiMsOM5ya8pqPrf10W+XqtnHUZaCLDSbndWh/+
go5r6ITzQ46xz1j5h+OeL1E/YMNcas4pBub2Isw8DDIbec5KXCDm7ZAshokYsz8x
k6xOuOkPklihHK1VzipqroRFuNxupXFq5820XcooJmmnvNZ9f4SfRFU6BwFRlxt0
XEqzPiiP8rrxxAv/2gxbmuJvAMy4wVGLiRHsEVuHd4WwC0SX0adZfeMA34WA89e7
3LUs5qI4erF3SsxCByQ3J69lQYcKx6YbGg9wl5PdonowDxH86zOAcpJ7rQqg/4N3
3/hFKKzQwTTaRpcofKq1hFSzyCP9pNQyOvcWMu5QBgghuLSJY8boMRbfokCQ42rQ
IahZ94/9hxowCJtJfRfIUl4DQAtl0vIqIriBqPtSwIVuuqSVJAJKmSbxSzyB997M
nnEaZEtZZf77Xuct/NBJZ6aPggdYTZCirOrMYZkD06C62JGgmaAlJ7CXu7ySFHN6
pcU1Z8dDxZbtuMHt2qbHqGWAJNVKup24nOWQLa7QEVtzeICJffjECJp7E0qTUNjL
PqEKHGkFxx3iSR/CNILuPG7F7QblSe7oeZRHeCpVvi4qREqsj7AaR8eJbqb3MxC/
igwDCV62Ojjxvm8jjEQer55bLfXAbeP45fML+tpM9NA+SNL+AGW4EsglhiI1G616

//pragma protect end_data_block
//pragma protect digest_block
96JeidHzfwMu6tfsPjwr9bpBjwc=
//pragma protect end_digest_block
//pragma protect end_protected
