// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
0IrCba8VF5SYMgM2xCpcBWmdpmidwrx1ZNkOzLGv3h5sCOkDlaosMNLWv2br
EpLzsK46zSTagYkjwWdY4OBejf/b0XZ8NBk/fXfhH7ydgoFzCNg+akBRAhrc
lq8kWie5X8JHSCZygZQ89c5tnXWd71vlFk0YmVcMtAO96Jmgfx6fcY+ycdZl
/Gu2OnGFlJI0A4XAKIXv7KRCYxY+LJ+tOyX4eGm/9L3z2B+9sHi4AWFrOFO8
GNStfZqfDrc0vogFdNrfHlGZT/vvPrTxSNXHBPIpNAQz/C7T0oWkVWZwKDQ9
sLgYAe1K/drPzyS4tdwPpfnUggJUHeK+eLoXzziIVw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
e+x8YtqTLLCtWCPQ3X2cMgAHZ7RKRLH+wklqa+zK1ygbrACuhzM41NjngdVo
47QnbaMXzUzWoXweMt+Y/J4aQqw2MVMf61/aeQy4v/fQcN4Ty39dBRr8S1pm
fbKv6ahWeYE87RzatEQ0X3OWDSTG6cCCApGQH8wbJXWBocQ6gt6ynJXPZMd2
LE/fhm2a2033yUmaLXdOJd8zVyHlujgrnaBTTEQttgycSTjNtD49gEyF3GN6
xx9IpdBRI6c8GayLwOllx6Jw/3/Sw8gcnM1ELnJ9np7VeTMpNQGROx6StriD
mT4TE7JZYkMgfo5uBmhx3adxUsZqYN0iyqr4Ro2FZA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
HPir97YLhXrKGVf7PDfx44fg8RNNw4A/KwRlWUKgbCn10HrtqECaCQUa1IhM
ET6bbm3lQ7ibxwrfBuMqvuSziN8R3P2BjhcK5VCA9zLrbs/MaXexjJV+XH86
RXiezHWHQMyjrAAqjWvvyo2iBHTlu01ITV/P+mC3BxE5s9uIu/nh43vRCe8f
7UGgRzQqaY7sUqbg/lnev1kXvnUtI16fIXVsGKN9zu++M/glumHeiUB5zXUb
NI4q6qqepAkWROKbeNIB/rsLwg3NUvgF56/tgu+hqEdtWaGvHoqjFiifUA11
nEqAzFe11R0OGbVGGbzlhgufXSOxOUOVO1ycF8CqAA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
p1JKCR5USnmf5h/m8S0UZ5VRUSCchKTY8Q9r5GgcDz1/Uvr/y4p4XLlC7h0e
fMoeZO6KENDjfAgBukVRGK5aAZc4DW3JQryVtTbLvhOPAZ7WX/a5UuGOAOil
FmFp65i4kVljoDNTq0TY9Gi3wiUNmO7nO6AqyN/ROvp4p/ZPSGw=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
toeWurpvVvajhQCY5O+aOAWKrRkMl2ZlGiwclTg0lhvfzKwUXZRt2gfB2wHL
Ax/fSSmwRBC3DPVRRGIjV/Z4wCNFWLkgcFnVPf3nrJLa6ecPZli9nMnNuGW+
g2Gnf8Hv+GqX9cqvOeTCFyB+vhNoPN983pTrpW+nuD8S9Zmd7T/57BuDhRcv
NI1VsFCQUfYBajrTlk1FaNGEmnbX/GWQ3/KeU/6XYpOZkKmsOm1i6e0dt0uJ
nmJPZrQbhrKvdMvaelEIKmtnsd2ilTTxhs9KaBXvFcMxgduw3EkneOFDaXXU
pa10th+SkdujLee9Zzi9yXS6V/e1NWjBRsz6wlktgOenxcVHtMi/nG4E4Ur0
xEuYtUDenrFXhRXOQ7I58ZHcYxLo47f0/s/Dbx2BpLTTPShIYSMjYHqTVygM
4z23aC7oqhoD8iJbYsmJSQRnvaWHTHnkjNiQRUWxu8TgvxxdJjb4BFFlP3rn
HgjTM+hsWE2kOhtVVLEVsX1KEKKwNwq4


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
rgLH4AgRSM55Bxtzpt54buJG+eS6ZNphXiYmgA9VLmF0Ve5TgREbaTRt1lBQ
DvlAWfnek6Tiby5sQxc6YqXYznozO7+RWX4fbjfp3bGUv+v+EB8CvNjsD4i+
SmvsDrJL9BLw0NVjSjPBmvgrszhbevbDkkQENbktu6qQ99dMfg8=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
EjvJxLZZwfWAEH2k1pbz3NnkGJqjW3d5V3Z3hnqfO/Bygfppq1v4gDuEoclY
xoIrAbReF02kalh7JwY15h+t9uMPoemWF40heHbCSKB1uLygHwjzVp103xvL
u9CGvEeSHgPMFUf4abTXOgC7aLhbvug45QbebPYcNok6nE6qJnU=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 28720)
`pragma protect data_block
zVhk1BYiEgZr3a3cmQBQguPwUh0tQL5quGOBzKMHLHKbyb0HjeamLJrijflG
tTLHdXdKS4jXpcsGg8HR2LRVQyFPBaAQJSnOM9TX65qFfKCHsiWpzSm+B9tF
RtKoeHCyTiFIUbVFrrQiAx6uGBOmTLzekip7x8rwkLoFfOdj56t4+i9Qx4Kb
y5h6XOmqYUZC8iOAqkwA3dXNUcmj41nyCWss+DKSF8gSeiAaCA16VcHq1HaH
SH77JvEpAK+dOyTJDXwtlk7QFPmyW0fs0A2yVnTkz3BHPIVmZypyHVeKhL1J
zLrLhZV7ERdJjUl2GtGVG6FryMOVX4q5qVHpNIS3uenXOmsKp0An6gOg/FWY
BDrKo/XSKYz1yHuH4jPzV4yB3YcppmUDg0rAC/E4M+L7TnLxRCNO0PiaSPMO
cpXBzJjDmGWj3nMzXw4DlpZ0eX7XsPwhQ1eF/s+uApgDgTZi86OAAxdFsnrf
AWl0p6FlAXJOGEs6nmaCVtS0Fr8q2YIzEW2goZ7qfSOeLnYO2FMlmlqF/0Xz
Mbj0DnIh5xcp7xql/4dbWv4yvmLOIAqA00MJQkLf7mKYhqWHPNg7hXF9klxV
lVps8yFQJ9bRd3OjrFatJ98zhWn48nj5NCe45R40+I5l+Z5Tj/VVt9Dg0PV6
BMhXdCqx4Z/iIkiYqkU/BhLzDirxIAAcnMj2Tnzc7eNm2wpz5zXcW6QNY8DF
yLxAg/1ltbthV7uTHlIRhpkDl5I+zm057uogb+sRQmlWqRhItSAmSZuirDS8
m2HFTSKqm+mIFsNLydvRMFZc+2/5jjp0OXSvTNDY1iYy7qHdvlx1qJCcmAi7
Z/BTU0+GJ5Jcuu5l0lLym7ncs/gIUzmp66V1YjK0pJfGW0dUKbeCtD5/wT6d
WlMtWUKEUUvEMuX4uj8G9XBE9snrOkWVZougdGJlkNNMWDvYYbgK6xgdWMae
+yARithSM0OW81BFsh11dvjdjF2SrVlKcMfvSjC/tMB9oJlpBk69qJ0QxIqh
PTJrZjTc1kBsDDHamgulmgeN/TSYYCNArzxTtwLb8Sdd0ZRzZ+xuzTmQ66Er
gEuf4B2Z/xf7FpzDafPNrMu2lBkglSqzERYRly4QRXAJXPni8WUZ2AOp/fUg
kj4dlxT01EY41hVLT/Kq7vCyz0S4kKMtr+pBpgg1UFJ/q4H+Vhy9eiSOLwpD
exrlzAzdw4qDcv9/fFwGvT68S/4O5FKzyXoIu0kSQwPPb9pgGn7ddGQU0KtP
UYO6JXtt95VQilNi9crJkcqlKwIAszJ0A2aucebLb+7LDCl2jb+af+t7vmjl
0HuhONaEodNPh4A60dHqhdDRvdNnKvStzdUDi1wgOgOLT6gwtTWu2tXjQpBc
B2zlHYsrSCtlouCbktx8afLlpICBqfNaiGqCp6dk0+YOjc2AHCjXJfMfeZu4
JrMlNBxPNP5lphbcOdD22fCzP3NHgeqCWe9OwUE+rri9rxY+T/mR4TFLI6hD
QM6tCut5bAzE7iyhusH3NFNubOFm49Y/4t+e6wlOHj405o2TKB+0flRSSzSA
odUYziFaxHBjfWQ1ySyIV5yeCX2tqvRI4CloKn8jRccu1cMW5lM3kVg+tbts
BcCjz9mAhOzxeJVOynNpnT3k0U6a4A6mPaj2W4xjcRHtjCcDEaJ2esv39+Tb
GiVylcogxTjes5f3bnQBGL5NxouDyJcIwNwAnYhXWb+nXhjGkaNeE5XwCDZd
XrYDXxxNKqAiCH2T7TIo/LthKBMsnh8lOF6qySKgLckDoK9JHBObrTTuPXqy
QOIQrJzMpoZAx+suSe3PcTjzAClDq893lh0ygVVr8bCnTcsZ8d0nUe8EI/aZ
ouZOXPfJPfpaLQyBFvVjIBnos1HbfdnZvlYS6Sch9HlClT8xS6JK9Djml/2L
M+7PC5AAuECvsOujQAEDalPRGNJ6SL/qt5/eT61dy7gt5PtOP7poxcd6CSEn
6NAOrIOXalUspOQi8HDtepSXXex1S8pCUekqBfA8BlG+eSJEanY6aYczCVqA
90+ba0zUUkzMEJ4c+QgIOgy7TBNvlunzCxilqFz+2sD3RHeOk5tlEusPgnIZ
wKAAQTajBeZNnm2g8nzMmzmPg5m9HO0v9/id6gpKoLG5m42Vam/J19oTiwbN
iKbdxHvnMy/VQw/9RFq17z/NwU8ef4t5BzEujcZ5FVWSYfVchWviIp2t0VWC
knzOecv4OIRk8/t+96/1ND0k4ljpoM0KWAGTW6LQc09CUuHtX2vKyUEYyvgT
mHoWLsEyfmn0+cu6QZNMif2fBvwC95dBkVyL3Oayx/Lpep4GMqxiHJ19Qv7r
DQ8wVm84PIjI3yX1WjTVP1zGj7YcPLzKuSUwvox633WePGAN1ZA93NG67iiy
pJTWusjZ1I8uTeOo8ESgmHASQoD0hAv0qIR7VG/2mY9YGMzNE14Bo+tvZYr3
23uZNFrS+4nfuJp1qBFUaKkpl5sYNG2tiJUQE2Ymb+ewByNsubub2tJHthd8
GinL5RboxXIp+B2O8rFUw7JTaoTbpyrLgWKa7icA3FLz4Lbnvp4UM6kkePgb
nfRsLRYfQSXa68zEcrOWZQJTSY44e656tSJEmZx3ni8/7rNzE6L4gc+wgDSo
Bx/495y/y64zcRfNGaTRls2/BiR99EeINpaXFzDQjiv+WGwNASe48Z/+QC55
flun1/mvIBP+jPZZebb+teuIM8yp1e7+QgGHKxNDVw9ClQyzNXF1fAHuRvDk
ogZ0iAqk3fVm7JSji0NxVuP4uvWQx5vMYw62r5DA6ujyoruovI/nlWYHh+rU
vRtMAmL++Ch0qfixqPf9HMItQioWYsqOBNuXwzxzhScNyj1aB5kKUNflrTdz
qYGLGTm0jQ5kubdSztUCLq0GgK0LFiIolVpsG/w5YSZfGGGeL7c6qsFOIRXd
ty6LEzzZO4mdwXuvDcrH8UaWzV+vaGs+FhXDBbG6RT2T2FaMXsMaTj/E41Lq
yaG3RVXk+uJrRfSFH+0Lk1T7OIRQn9qH583t4atrKavYN+f/8PrHKnOyq8Xd
hYsAlcIwx4luxgEKqCMFS+89ZobEynmvuXzYegPsXxx5+4vKFhpt1zYFvZFY
vv6YZVXHmDq+r6VGT5AqnGttxNbvpgjwKJ69KAdwACsJrLs+WVMrasp0qty7
TOnBZ/cwy0D1FSDRozYaw4p/NUB94f3fOXAvvTGt+d52JfcauP7jxzxIbgsv
M9v1RkZLxKZCHVvf3zqigbhdFueDLiA69TxwW3gtwN/15bpiD/lKq4ti58VS
Z1iCX2dLGJBEt/y0JX3bGiSeAHGlwBCgIwZ0z0+U+VJ4dw7dlHCV6NugW9PH
JL217yyskYHXMkUo0l5O/uFTIcESX03byAHz3xnmi6C9x+hlukcAAfj/O879
JEJvP/rDqqnl2uuu9yj0A3ggachYc3gBZgds7fC1EeDZBrWcEgTqlj5xTzBY
XfYVedkbvqeLcZc6J0wGYxyRGv81KOZxqL75jHQRKxoc3pNGHe7ilpzaCjHa
jiq3W85TrVgkURu9Hjhyc7T/94EijnjSYE56JkZbb7OvSWM6FvqN6BOufngD
IK4/OqQhQbrP8S1P2W0AcLCoKpPuIvqEdL4YYR33GNBMAvaNxLm2g+SmC1ja
bqF9izLzIwrM0/27o+gQGaTBWCn4HYmlFTVe9v68LX0k0z/AyZH0bzHKu6Ta
5Ly2XoGYcGXit2l3oCuXmJHPHrSMx5Lpgpru3Z6QMOd4tQQddZ77kx0xvFyl
962iIPT6NwQbCAprPv78hIBgTNhV02EZoLwq7Ypxho8h/K1k0A5026pi06n9
VB91wkVVv8hJqN6I0ZZXE5lTH+B3O+tyPMDG55KoiH2+kGRMZUfDhdPvuXzm
jgPx3AvBRgfwBFUeZPycG3Hea/ay/CqzaQ0bSZWgi3d3eyMKf4w6okGcwhXN
2ErZKNKAatPvkjujLvsWq5wljZn+jx42dK6Lpy0266Kgw/4PwXvo6uUGjKof
BbDawrftBZO44wUPhDN+y6X02lttkvUw/7xkgL77Sjy+w/knowk45K81EqED
4lw8wu/Fv1DjZJj80acOrmdw4OJJAyYvEWWkhPZX0sBJ4zKiN1/AfA8wGZAu
jJe7TpNv4uTdZfu9OBcA8KvllCEvwFIh1wcEiMPFXUeigt5Ik8k8NulQwYGX
8A/8XeRZK4h2Vkc18xmBCzGtLtCQ+BPQWUl+0nYWrsyNv6r22gkzA+yk140X
IX1aLFTAyW0Hq882gMdfBTYTRxFmAcUNT/xvQG2KTkOrXbtdM5nq29gqept5
zQZ5GWW6xSm2HLOV4oefQZIwW9xNNXlZNArHjBJ/UP+96UPI41ZLZ/iqL8rn
xZdfPn1CtqvlDFkFhGoeOS9/cWFfN9sEjYQe0JFQbc8LpVDRwLX6600DMpFQ
qECj5QFxeHELE1oj/Wm2FjoWVvCxILqXRcCBHXP1VwTMBVZ+uZJuNh4JmWmD
SnVj5D21fCOBSHnFQYOav41byEhlHVlzyHkR1N1ZGDDTuYs2LfKaTV4M8jfs
RtgbcqEpOcxc4L2DbYRDTV+ED7n40yWmpqQnxuJahy75deCMLIGNlOg79ABF
xJGLtuaqVsWRePcn+VSiBMNgqxCEn9X6nGYXSX+dT//5jjyIV4V5VhH6WPgI
eRJsyXBPO11R4hPPSYYvEe+J+/CNsHduZTjNOk2FFqrNV64WnCuRBrNZvDMg
jwTcpasgaFD3slzqLveuH54Ljd/kWPKvYoOEsfwd8nSrWjovfWZIZcH27P7S
5BdSY75cqq+MoBy92+0JtPhjfDvxyFot/Ym0Q5Hi1wYkDzOqL9yUxciNV/9n
D/RPh/GHm6ytVK4688OJCsc2nBlzhHfvicXC3iPxnegdD1/0LQTbG5s+3Axo
iPC3Ljt1ESqF7frX4HvaTMClq2ZGAXi3H8okSKGqgoZ0k7HZKM2cHMp67gYR
ZFhffukX7vGAc8BwwIslFgNckupyUlgEax2E0tmtOIcPF8yQ4Iz107LWXZEV
aPAnqLxjRx/vlBwNtumYaQqOCZ0+L39LyWGuQ9lND7ZEaaw11w9G3f25a1hY
AUPCvRlDMMbTLmmy2FEsvf4Midqd8ah8PLl8ZrzHofSA0GtTtIMh0GG2FHxg
tToXLOb6KthDxtmRIGegegtkQ0vHTcue7Fjdet5mgQZSwdmkB9mLVAgwZpWH
jXCMi2cnvISAe9PnbdkGnVhdmv8GUkUZNg0aPdiKExnxkyiER23ugABE12M0
a1/lfQc+gubKibxKmY445x1Ct9EL6/FQBMoH+kCwLDlTvpjNN+Fpxu8ub22C
EdRXNkAv78ILh3TeYrvWwHF0WzyJkmDcM5p12kV5tGRuCrmAjBv91+zmPZhb
di7GHh7ROuBQCNRzWHevjKrZ/ZRm5t9nCQ1kvnVfjdCPq+pI0qL5gvIKCRAL
oB3GwroZqhoYY2hGRIBHwYU9QBB9QT06Dobuxj+5HOpEVMYpkNuYjk0e9mr0
IyuTL87uUGH/fyBCW16RXSfNcR9umaUdbJqEyk0wiSO0ppgKE/bHO7zPyDjb
zZUpACw1FhB5b7ntYFm3LBiwJcWjXlrSeJhs5gWC9vkWtYRcqPnfPfqGzfcY
DlN0XG2rH3tzTuGQqY3KAJGRW2Rq6Q2JbwrIPEauT7Km1rZDbT9YRWy7SJD+
4El2zUGx1XBI5bBNUHx9n1G8ht9LoTfZB/97UfqCrDS1uG50rXB0axb112lZ
R8u7opX0yuG6zQ3W+KdVIXwSEZ+I/mcQRlmFECGPdYdCs+e3bojkuuQT98Lc
U9OGbs4qeKs90IXZoV1eSEBugcr55rU1MLkPhprcZl1xLQwMFLjWzFWwCFCx
tRCm94WTwEKWeysiCVvwkd1lHK72GeL/ZW7qcFuwICLSYPaBwFOgT6Z0NG5/
EKm8Rd3SnA2Lxr/LFTA7CcYAad8DoE7BN0CFUZ7NjZOTJABG2bLDaUMxyKeO
uQ1YpLLA/+rWBz3emYvVrmTORHHwL4JeuSFeRXpF+Kuke/zKeNnmLU7JMgVn
27BdH8tM9GXL/bvSKiAbfgcsozPoEC+LvwmNQtCS5DCLMho02XushEs9X7VH
+ljndbmVkMAeG5aSZQnlJPfibWEokR7WZi9WMlvH4l+Tm3/lCgS3bbIFHQwO
3Q6vPLSJzAUjHtTpnVuXturR8W1x6tT5xAq99uyPH4Brj60qtvPtBY6a7UVX
SFZh2qzmdSb67gp78oBoaSInT42yPQRhXC1XxmcL61TzGDXy3rLMGh3csu54
+OOI+7zeaopikh33izHPy4Ox+890MVAnlrmLg8/bUO/wmAWxrMV49+3/lrb6
Xr2Fakjmps9msciY0nBXaOXAPy1nUbqg/g37EqHI1BNoRpD+WXvXsq1eI5az
PmDiKbwsQc9zyRd9jNraiMiiyQhtNLLCKYlG1d/mvaI3+WmeBHRNDRQGhv+K
NmnfGGFgnIa0HOvtORtboN91z3AiNXLrEaOqszGMcD81QX0ZqgvTrfv+NH5c
pLNZg87ij2Er4WObkVEDObbQ8/eDPjSyOqyx6CK94s7zMeASIKq+7CJ5cbKN
hR1oFpsPouRpEvBUYrKGv0OT4oR63dzFJWBrjna70+W+60S89DR+zuNRDdZS
k7DRr/oSQzf5rt3RuyOsuhGrTVw3ZFVhRLATK12m8TBDPehirvi5VieGjhH3
4nTLP3N3xWYLSG736WORLOSRxM/VNUboXLeOYgUrsYZdIJfYhuOR8AYKCngY
HzzvEbzq0NBHtnkfPximo8/xnS40QGrakjTH2VVOSnMPzRG3L8q4vog+jbZM
Zo20E9TTAVA4S2XGgBVS27jpIju2W/VLeJnpd+Wds/+IOqlD4+DOS9mvI3JA
pXEzLsQq/W/2c+m92GhJ3HCFs7cvnzI8150xza2ReAJG9vUHFY6T2BkhAElQ
K8CDuqL7yRDzk8Kr5QhlT5cRQbFiU1f5FoduHPP3rQ+fCjAb0aclzrEo4g1t
sGNLpaHvbkwb/i41LkDUThM2S5J1KZqAHMagdPSTWXK0N9b2HBbyZYbHm2ut
Nsd2ohxCHOngZQRdAc3pvZ60GiKEZIDwDLE0A+SivishW+iClIUeuOAoV/nl
SRtMLNrtICOZ48IqH1NhCijgleAnFC1zLGqcnJFOcUK5gY0BJtZ10tqLOIcH
1GxqRElg+xb8CyW3RPdfyO0GQIT8Jw761rIEMJdZj4GvEk6hmZ7jt/0Xrd9n
0HHSrLwm/GUuaEiq5nvn1/cirn/ayZgCH24slTSW4arG88xoMwsA38Bc7xWZ
GQ4glAl7iLOLFbBkKg1pmF9hP7LpYFD4YexNlSLD+Uh6EbFFluNJrCUnAFTj
ledD4hOSHDG2Y4qkllp0zalgHzDYgT5UNvGtHt054hZWV2pjyMxIBAzQV2Yp
Cadca1Q7MZtzlm4AV+vKzghpxit4iWGLimXakzg65XmsWeBY4ORlfsk4Wuup
U2+3vi+Zoawaff6d7hwgpN6PpVRhCNnLqz3jPfIeeISmPg49LnyPnrUw7Rd+
CokHkblYvUBz6eRxc23fhpwTa8s0GuxjJWpBwNb8lkzh4hdkeDOMbbDod7Rx
TrYk7Dmo1dshAYNrdqXNSU354ImJqZtuYfc6c0AnNiu0RHO5aJW/bGMXZS08
ytOIgWmccqAp9j0Rjljv+mmLUU8GLA77SZ4RX5MUlUd1RElCaowJXkal5G7u
R/eq3/2vx4/n9AZT3+SKVIS/H0POPvJtKcsWIQuqaGRl2XS7UGJl8meoAfzU
MhBDsFiFP+8JPFayyyQ0LiK3vS4PtP6FwgYhF86HYFYxtBTHLg1bkGEprDXg
pzqGUzuj8fykjLx1g7vGz3HFj5nNeofQ3YwMkuxOiTmKukaQurliJYFk0ug5
2YfjqnVizIRYLxo5loCJ/swOGHvo6u9IIHsrIzwI0GeWPYF06Sw+fLw2IMGD
dRKkXs0g1j/pP0cAWAgUwtor12kqnK/QsGRuL4Aozmezy99BDAGyYWiQlkan
bb+3YCq4rOpPNv9lO3y4luL/kbB6uKHjkdwYp8Ni/B6Uo2ahuwmBw/YaiyXt
zBbV6HmGd/UTdxwbf00HZ8+L3U1NjI7OoibDsaqH9czh9XHHCv+f7BxdVrh+
fgQToyq6Gm28z8XymsTgdnn284LPiNrZ+UvddLbh6MvFGTBWf5/9peIpCKS4
KOOprnDG9Or6X0n8/5de5m6ir/sZsw5OdOjFgpT3153YnfTTRiA/+tWzd3g0
RSoZnP0RxXHl9vk4jN03iqKGBmZ7d7dXKwjjmtMZhTfDteoIvlwjNat5n41q
mHWZusargreSXaFZGgPw+0p3nC4QVuEgh8PEaQ6GzdwcURSkrCcncgqbdR83
1OAMxkYjHiGJXnbOwzziyZMP9/WWSuFyuMlQ8sNhp8r6TkVU7Yuz3RY1MCOf
VBdRk/r3HGgIDASeaNztGpw7rOl6NiImUOfQPvVaSXjwYI39z19bdRxKFWBD
Hu+4PSUhaXEAtzr37lYwyv1Y9tmwvjoCSMR9pDxBRa/UFWw8B/PzodJx7f1+
q2QpXVeoePQQaEWavX3VGPVhZtV7v3VND9nc09XTRBJibHiwPsr3aBnO0GEF
Ai2QRz9K0fYubkORGs1CC/msk7RJKVKsKwp52X53lcZC06cOJWSX0UwkGlzp
cuxX+8mGvrPA52PWLR5f1TSZ9sprUUDM5lNNSvswu0RYHcwnskrO0zVrKTka
dV+PLjDSZgGz79yv7N/OmOFSh0TvHvjUePcIp4ri3mO1lc53CWeKcG0MIFOb
nHt/zaqxrHfF654S9LkMOhjUSmweiFZOdg9s4Y7aRDRCoo+yYM6HpaycAW8/
2t38yPKjd+WWjUDmMIJOpnlnImQdzHbF79uCivTGH/f4hsO877U1vFOiuWdT
JMrQTQBex1egeRJ3NYMk1kBBrl9/b3HtqDzM2hu6ksusTistetaGrj3OgHtP
nYeWwNO+NTT+moWcHP4Qu2CUBOmre9JopErcwkY9s2sNF+0IVraWL/qskvDG
S+OVxtOAj4EZwt5OCllWMQI+L4U5cYgd7bezGiaSGPv4i0AjWlkUqXPyi/gT
lo/hvKK5ZHuZBAfQJKNqJuc6V+/so+DeVfPOBoqKegQqIU9ivMXFKdePD/fk
iZzyDTQDVF8b1ZCtonvY/8N1aJtyj8h1SVAWsnj1ZZQ0H4uSx7FjAKwBLb7O
eVZtSkLQyLI8eat8i3kZYw1TtkWzN6Akr5PSRhsXqnTMGkjO+eRgzT89bsO6
ZyrUNNXKoTlVcZq11jgvIVVaTz8l0/+0odUwgoOSO61H8JxvrPmozXyY6gk2
eeG7noidYwDHYp+n3dZEPUfjgpIAr8Mp8IYwbuuU+IdqTXY8X4NHToLj0czX
puyQSw4pCAHYm9/ML8zD5h7PcukcD3tpx/WEgLiTIu6KIfGvxTPmEOHTChHX
QjEKkanwC0a7X4YqqLEu8GpqYciWpEH8Y91G3907qijnQG+ttgn4Cz6ONFw1
umjjeNcyUf2mcKaZd6q8FvLqnyXsunGz+P1bdvA8X02e0x4ts7/Cg92XtQUx
whHOM6fZJlC1c9ocwCUSw9ANr2IcuNHjw2pLyZ2tQxngYBP6KQvhMjwk2Apa
okkN1RcnS+c7ez72Mp0WVWa3rfvVK8aTEZ0CvGTRx2WNWyuVYt3cusK3u3i9
0bQduecBVu3ZJlQIZAp3iWwfknSwmbTGUIMMGz3d8OdxdtI5WnR30dh4CDuq
03cxbxQwG/OoqWZwRBkuMoUSEoSyGFpBV+wutMYMOZkQgLLPR57LVwr1xGCy
+ptg+PBZH09buDC78wSg2BdVup9DDVCfiuOoP5cOs6qeZDsg80f1tgq6w5yE
GCzkYPjWthhHi0iCQdpIhpsyrOmCV6xjbcS1BB2Zr61H4Amuqv2nwxWnRsWy
keLGSoAeRdktvJK/zeTjqx5XyqC4XwVDXqn1CB+yO5v/sNuaFUdcfRWX2FXG
2twfzEGwc05G5XwbLTgWMdsgS797GBv95jVfQu/dzcA4bGCUoqA98Rh19u3W
9OEylMTbV4Umq87pQJXyfzy8GpfF7CIwX/Lz3mtwn4Z8aMund/ngh0i/odqQ
8CBvCHrK8IVYYy3FYKi3U1sdbdmrVmUZgdZxrENsqHhO71ai+8dqcgdu8mBK
LaHyH9b9IV0+qGOo/MuvmUq+sapNKc1UZMNEutix33Hmw4ixzrlAYaeaJxHA
JekU6Vdj11DeAb3BCfLxkjDyIukVJn0+LqrnhhkbN64G88Ix4T+Mxs4rTZKo
2P7nt5FwfkqUiWMNxujIP+kRF/OhlMIGueFiug1WGNIvbwLe55eBdMlb2tm0
uKjYwmJ+rB5GBYaBnqwQ1HmrEU4ZWQp40l+z4CV9jjNqWHo/x2BbaFksCqu6
v9Fm4xvSsnrdwEDJmY3+BVchwR4lG52wBvi7fv3YTJRCNNc+qzsuq3ks1/O7
zehL3y6hs9vp872/SVeGan1TBXgaNs433KGtEljCwxb7X/4TKbL2vBKsqIIf
A30MtN3uGwzGx+JvD8Rc935Oux+WlHKmppm2Nhu6v1gJpoyFkZHNM6GgBgXw
XYD2rfli/KivzXUaLc2KgBPX67hlsRQpVuqBw/KJ1adHAU3ID7o0R+XarU0k
U7N7YvUI+REFgU0TlfzwS7bS9GCpHzFasGGgGv1S48JGRJxz8+wdEjlwEb0r
OyRBJlskCT2miZg5SemGa1E+FFddHdoRrqbVUALaxgp+iEDYyrQmLrTcqtOX
Xr4b0TJ+9LZX37NpoBD00ARUYWhgSBDi+5JUhGSjvQy+YC5XeZCV8S1jHS7y
bmFkCLlkJr+TfGilBU8slIGaySUmY7ywceaBHwPLlLImG8JACvrhm/39IPK8
JHJRpgGOUH5FZcur9djRSwG62aBW/bz6MOqv9z2zDjeSIVYcEqBIB2miOpoG
5jqLamYkC3v4tFTGWbhatGGRMVk1YbZkfd7UqaXpYhJurWbUTXlwBw77+CMV
lHgnt1pdul/mVnToycYIzoggL1PMwAY5smKxYfW2JLzaC8esP+n1z2ko96w4
LQYyqsTT6WHRjRKz13u6NUuz3xoca2FI4wSfO6JqOOuWuKS+UuL9OCnueuFp
Beoz6xV4iptEMdmNaq7o4T37l70fzWHVJPwvqPP0/qHeel2rCvepC4y7Ag4l
7invGUD5WqNM4QPa0VyacslYBMiiflMvdYHf5tWXJYn3pX+ImCxVECHNCwrP
+xea6qYr+Ytk5D8n9SDIIlQTl4RKjlr3heNWBt1VjH4wT7rOgYBPZnfJALHD
BTDMp8VqvXzroE5RCjUhsI5MuG04bENNP5uC4049n4QPg7AvZIlK++47IXWT
T/FIota6zu+7Z4XuiM+OISnNsoqPy1nhN2YlAleBfuDXDDUGiKijaBLrhwWc
ZjVhwAfH3N0FEc3QwJ0OU6qS/mFTJNI1w1rVuxnit3qqTVLwrXWVN5NcYXWm
R7lU8etr4Z0/pxqVcsDj1ddkP1nsShPY9gQUZmqJ+7PBzOq4JUDskPy09mYd
VR3T8hJhUBduLkP9vsk/Xk1XCLRW0YKFY20HaTcSLqcfeLbplwLq3ILVQrwU
ph9fMq0aqUzT2eF50GFEBi63OFLhHpbDQvM/PzN/EpFnECYwumDljdnnUd/5
WqzLx5XvPIBN14BY4ilOBPffC/DJ+Zuo6gZWsG1xLf/vtbzhV5GGzjN0RIdC
C0etFSYWlKmUA7p2PsymmKWoqKD5/zWjzVt5SfdwwyMJ4KXfcfyxnkGQ8AhN
oPXWYi0W8dX0ZcWTx2em8vzhhx4MahgrYdFFt8i3nnzSmDKx6fnAOObWM+ZG
wRk3wao9m5NUZ8l0Yr7Nt+rWLlohwS1wTHSbCZcdNdg7O5Xjy9vMWv2DSk0Y
LbODRg6aEed8kXdV1VGdAm5d7Od+XtNArcKnM89v6HtWSOqGIYrvsf/dGHGd
lUkxHglaqK4X9FJb2gPOn3INSJo2IbgasLy6lzBMJL3FwtIRVee4QSs+jGjc
7VDHxAnANUyeoliolbTAcrUyv8jRe3UPIUYYGqDJCVl45HmDKva/t7qApaQN
YQ9MFZASrV7gFA/09K+JMqnkNX/MU/TYjzpp8oFuK7VBdwm0WncuEoXZ0EeF
9NgNMFvDmKqdvcpJY6Zp1GZdPZzHlvBaT9RT7MiHOpWbYHd5U9gwDvVcrGPz
IrqWn9UflBge01k/uOGSVwKdUlr3fzKP7dB3SvS60TEt692pOCBxKyyYX66A
sTXJKHJQ/DGbQfbuT5/kqMN3iA8yNvO9837akPXIzJmNUG91slnp6iaFB5T+
JaWhBFl7uhXDUjDkgvemz1+qrSiKimHaPw5NF2bYfsB8fo43FM9GDev08fdn
CEYue12Uj8pwV1Nes4LTLgJmQgAawbiSd2bWv/sg6Pa6iKtvjasojuzEnUXR
yzmuP8ievt3+F2M+YPLLbAV5ELMqYidQ12x4VKxP4H4C8QPgWfS6mgLEkfOC
iIZ+BoBCxbWhU8ttweFMCUibR5vkmj732l6j1Ciu+Tg0+LApj+59fSrNbiaO
JqpwSbDBPHclr0HtnHx5BcQ3tOuFOqaKzgie1HolhWXFoTBKPebRMNaGAjdo
OQ7I7PPwI9ahuT10NvMnkWR2OqIQ5sZLtH4gxsr5u3ZXXiMSOuUliQ3pxQGr
kFHY1gqPjNh7LOOB8rjg6lsVKsAXd4FuYnqakzeDevEqG3Tsk2TlLkdFcyEX
C3+gAI1jDIbygpgSetveqX9jZzk+IBvbWu+yu9D1pWl1WRM/oKe2Jjl2zJDs
/BZAUtVX/B1+J5qmdPmPiAOvJY783vvetuzFepIY++3zVM7XiRLAn4HfaMxx
VJ1ixHlCsU2ueKxQ4Cji3R6IhtLJtyr9E5/UUutfzVj0sAVzp82IDlt74uoo
2qFzMJKabRDSxl/nknGKUVw7orgYKNUKDXgqr1He/X5fFEjzUIwnwn6mMEyi
dwZEoDBSCPtl80oaNjR1rQZ+46zv0BWvGst27rCPuuWa5Lsst/+Z5FuaLf7h
RMT32lSI3qKQawhDcPI+hlopi8sqrmCyE8YHWyOvmMwwxJVnWA8GDGLZ44vq
A34t0mVN/sSNQsWUbEqOzgfKXtncU5YrLewIVIh/p+rtviqSI4MQbOmTg4rf
tN7UPU3uqCKsfgftUjPK9lYSO6Z5GWOoDMxKLitV1L4ei0t4OvGqpmGjpvU6
GBIwTnEXOSKxAaBQ3yBEbCw+D3/caDhA0o0kagPI6yVCuNFxcJtxm1Wa4gC1
2pwb6jJyn6E0zhPx/E0XK199hVwupjFHda2BjYLv78Jp5NHtFcosyFL4Z1Mt
gniiuOaLNmI82sGK8Q2TZ6bSK57Wm7Niq1yHzkaG9Ovf006C/8Q9/aEMCOZ/
1x5qe7CM87NEj4IX7Otj58uPkgpsqnVOFtGdFWFggDEPmf66jH9qLIWeCblB
+wVkTbgSTDD2RWmQkXOdpFeHk3o5C9A/yNLxh6e+yM5K+6orYmtNlV+S8S1u
PCzGJvPZEy/MsLfxygyZ0CrCEbLomJmuwIwMIa+OBoUQDplKnQzjANOBQFG2
rrsk8dGyMSN1WbWNPoGByEhWwwFmgZltRRNCFmt7v5RVX8JMwX7t1KhcAAxm
45rkyWURTEPxF3yGPf/WFESb2FPYSrX1kMspy0ZqPxpgOPjTYtQT0LNcrl5N
SFcEpQAG77Lgxm+M40lkqZ7MPGVYQ3Tmp6SLmQrX8Ogf57zBGnj6lwojXMuF
6L8rGu4dnDR/VvfwoHZAbRTI0yHneVxMbg9A/rPWp0LrJL4vymbSLc67aXNu
xgA1O3glnYJ4LNYpG6RdciwEGhlFkE09ILW06DiJod/BiP8XnJ0Q6XQhxn0O
9OoqE/t3Ia+YG7QcGxUezsbSWngOwBiaS714PU09Sn7H7id/EznfeAO0iDCw
PqC/tY2IaDnyDMxLUxgL7mksfS6LZSYrDsezEqYkf7e6QTwreeeG/fkaHTCf
JYG5+E2X/m6q0VvbELS5sovsgIOOUDc9sVnk1JsRkRScqTWy69vdyBpZet0K
9XqsGa2+XQmMjyvijleEp1cidNzxHr1OHSL3Z5Lb/u84lpRztucTzFn0RCmZ
wOloOBqSNQlAK3V667LUXOZEHHUss2yErjtb/HR0IzLicE58L3kT0ypwUib9
EmiH14tYNuoCkQlLedtw0iuMUVpXwKxy+JNPiYP7qe8bndvLiGEpghTTaGos
zmzMKKEeD+esdo828CCDvMa/tDK4KS/twIZa52W86KzZrBLYFwbvJ23m46ua
7stwNktmOr/XfzMY8gjZ3WH1li8BZZZmOk85wz+dBkotk/UM7yfc+wS3E8i/
MaDIh/QmAVrPSkPmD1FvIFF/tw2+TjtVRL4wlb5dNdvvVFkfvbMhTQV7YCfm
Xj1Gljl6SzKFVG1c46cswzXj2w2kBdO2mwSfyDWkRqUX2mkiExt3TJ/IpN4v
8KOYjl4OSr67AApc25EVpAdw6bRk0ke/AWdf+mpoMKjuj1/PyyJp+PkkCrbF
qz3xPiJ2JBi9JUmAy78nX7D9rhTiNirxjgsoUHHpV128eYO2f+tntOhtFeJw
L5PB2zyl+RDysC5boXCBo+zNym5ZriV2MC3McezUCO4t42fhJobNJcAhx7je
vaFCUyshSY4qFkMtlexAxzb79i3ue3IT0w11r5hEKvUKfz1GjSC6QD8bUBIt
Z3L2Y2OU9DBdBEUogEepLenBoVRxwH7ry5KdH07EjBtt4vG6oa4nF9FePwmZ
9DopSIiRQ9Zqlql8oImBMRk+UTlLDMxo/g0myXj84BViYo6MyA32cWS8MTmW
VnAAA7AnVkTLNGZTCdWEJctskjuRx2A0XZ0DcrPBp1cBQv+7+wu78CB20vTI
TGIWOYFtnrxkNOOAQtqLTfsptUStEhR5vDC7M0RFSusNn7EBCLmXFZM0m0Fc
EUfl67QG12FMbvmkhLrZv7QtN/r3BhM8vRq/oz7TySOYsshpRcXenun1Jay0
+kfWOsWgAi2eGuxZI8UGIOAHrwnnd47gbkap/cAUR4WpyJ1cU7Xx/u7Zbb1W
D/3vL6DzG81icIhpEkohOY6BqlZyiX+UyEFdQC9wOj7rud2YFVSxuFRrvXsx
woKhrAa516tG/KDOt186o/cZdqEM5IPs+chX/bcV17EWQe6p4AhHLOAgzmY6
Tft7qIaEU+fCvf/5D6k0QouFglde5dxYb5uykFOxtDolLKVZ4lEYxwfxM31o
2vItkYor5C947PVB33Ux5NFGZcL7eFiCEir3h4fHks6XVP3SPWOs2eKfJTI+
/h18e9VZ5DbqdCi23KCTQxt6aoXcQII22buLomwZwjOb9tKwe2Ikaqt0eIBY
jqGAmu0x37DtJQzzhAxb90iiV5pZEFgid+zr3SLlbbNMEOn8/T/m0f+W8Eho
RxekDdz8cEyvOJ/+IbYJL/Y2iw7AQSwHbrwVgDsJgP/8bMIymYHjVgdOOy5y
c72cFQFrIlgLdZIqKD0oSmLiyLzusY32hjRnPF4xEUezG6K8kaLog4gwakEW
BJpMOXiR2p0NSmMnM/rKIQ92GC52FKtahg4VVAuouVJbTnSiou1mua2BFC9Y
kPu0ceSm5ke7tnY7DVau0GEgijBZ1iwVdrjc+W9E+UnJDAWpT4/XhV3bELER
6FYaMm26LvbVQ8XBD1Yur6V6TMT3ifkciVY3uXyw1b2NvHO8XoOm1RbAp+Mo
y0Fs2qBXMKzK0qBZYqGMNp3HOA4cwttHHIbEmsCl3TxnS8dITbaJA4FoaRT3
bFtNepnlcxORyF9IXL/fSZGi6GmhG3qspSHEzDbF1mkbBHx5drupH238TSv8
/K+ibwFYYOXY50PJ1+iC/jPqICsK6z4rTe8+/yd1YKq7o67rnjioU2Eavuul
8xdidRe09hccu9BXdNsLwRI2pVUlKls57YrlsSb7aMN0SzocbnQFWGxK3aup
X5KupEQjNXLG7jUbo7jDFt2rjmhBPfBQPxTjk0nIP29+vw5/X62qJAkwGjUm
pt1Cpq9LIqAMIn9ibqtonABLHDLJc5j4UwfSWrAjb7Ewm8q4I6xnYEyeIL4v
7tN3HeE8MsgUcDsVi7DFQcFhdUyTsGMXRbqGzIPEMgpI+xo0pk68vBNBRnqn
QsQqg04DKXdCilnlQQ30e20Um2Q8/un0v2NREBnLqCGCzsr6EwM2GTktVj5V
dp/N0Uu+lczuONMkG8UW13F3cSgyzQd2ws1lqB7Z/jHYpub77I20ZxT2qvi2
aZchagKRKlisxEfNoSDCXEB1Ft6176uHAIIRXE7VkRndwEjGNcrX3N/KFCz5
hIUYvK3u+x5jAI4Nq9qnHODaLoMxyKjI3I1DNgoNpdxkQtjA8t2BR1kPdLkH
yZ6JAT3pkJjwbvWy8RBM/Ol3LshECFClteNW0xXO5wN80c2HWXyDPx9H2/Qh
2bhlSIGTWnvTPs3WYxdIk0WKAYyDA6mJVmZ7yaq/As9lp5HdbEdErKR01fxD
EAFLN1bPxkiwYt6IUSHuf2U6FYSXYiYdKfI5XmBWvbk5ebZ3FdaSdIaEFrbC
3XP3HcVRIVj8tIGNSBy3VMt8D4W18tmcyI6J3Rr7JADQ/mYPCQ60mS2sztLT
fNZG42mp/WzH8LqAZCQuv/6eeNtQmph1tvRsXWRmkGf4bTn2Ypz59yOxdkGP
WZkw/aI8HlGkLRX9U9/2KPMlp3gF9Lm29UvdNPxofGw0fe0LoDB1+lfMlfex
YmGTgyHtQjuWrSpbwohlq5m/cejj0kSqO6KC6L2IBBD4pZ8Cx0qdHf+ixnob
QOQc3kpyK8T+iajHKrA1EfeAAnZw+7qSU68VIlWk3q1NJNiBgwykj2GG6Vk8
uEurtdoagVGZmDp6BsE383SGsQEuk9YWEAyMP4DQWnnlqV/jC4ZfDLZfX/kQ
4VI1KtjenokCtri5TzGPu9nj7tOIVMyELrMFKFrbZMl/M7qewpXRODyaVHif
BB0lhYSCScvRfNU5ZYHJnN6WAlgAm2tUgvdbVFh+hsNsrQMg3OVozDFpfAjI
FXQIMEjElUtR3A7hAEEztefgJaV/iauZ7v3mprtNcMOMOXyiW00QjUOSjhar
vbXyUSOuD8bvTiS7iLkVXjc1cafNF5qXVW0o/w4cnUv/mZ4oWdxoHHCsk2qS
K8mK2yav8mSY042cjCe1ZPy6E7nspt6wKBaKmpo2AIQ9E4/3MrZksw3M7Be8
6ICpzX3p67yN3ymTOcMOJcAVl3Yv8Cvd7fZVTdPYh34HFbqkxd0GRgmy3H0P
cHn0qUupQu8ZpF3cGGNjEGKNr/Ft2+DGeitwKTA8Wm5ZGY9Pb0Di1+xIx16I
zZtJ6f9Q5vfYU13TeR8f3ouEAWehi+U8iq5iIbJLkz6BTNA8R9feB35JRddo
V/uezmPpnDsp60nrhFhqBdB1XVeMUgybJscX1puI1De+V9aOLMHYVrnn9Bvo
CdDNBy7KtP/cByYMbCPqCluejQn8hCwk1kTFJFcj9CF8mi6BVS4FQaQ6zRIQ
L0DZ7/K7Yn9M1y7h0WA7oUT7Rx/l+vItJr/MYMO/sqkjWKYFkZZgtjwMJsgp
9WhO0vnqHLs+hcAvs3NpvdE16UzWEw6mKr3Yz1P3Mh5cufRfTD08VdFpsfRr
LhXrN6T3zAfcavqgRyVHtIduq0LP7a6fGxF0nvU+M4bp9ojOr/KP5OcYNxPy
3dzhTy9iM9ahEhXRPmyllVS2N+qOzSkwcNyqtPT6nqgC2l3yFPdBaNnsgF2O
upTrmgvAedBdYPstoU9FSiMugrW677nbBlFr8RcPrnOoSM3xhehh0pJduHr0
TEAisehVuFU1QU4LLeW8yyTzRdsOEVVC5+t/+9/MbMycaVh37//8hI3NHZQj
sZZcD1yaGDknYB5Qwwv/YGPUyBItWotTKorMUk+JVlq4e4lQPWh+RxwJjk8K
N9qWNLzrOeZ8VIbBtRYc0bFf3VVWFRKdaf/WmbtqvOMoryjvvNOgdLDXDOTE
SxXia0COEXk46xBJlqK3g+ho87RngUYKE38qPdJRkh4A4dXKHkFtR7XqESj4
S6RklyZlo3CfGRCIDK53Y6qMyjx/dwoSHdVq6I0sy0nbGx5iiH9/zv7Qngvp
E+JvuTRS61FBkHwWK6I1eDPgo96eM5KW/Enb3VVojINGA2aJvBggo5WAbwLt
eMJmlRqF870D5LxxxQtD8d37JqvAP4VcZ3GzpJWMfE6rVjKNEFrQ/rhfShXG
jtCwxaujkN7yR84r0HRSiLkk2pIETJ2qas9itxRiHWv+yCBb5NjSuxlqBofH
y2HR4TWh7XUq4ai3tCBUYkwS+X86I3tWcDpC/6LvpcFmryzRj5RfyXh7AyuK
MsfpYAdTjWgeHwuOH2o0NuzXHFbVmEeNheccsmJabaJC/OjeIop37ktl4OTN
u4KF7pq2P8DLdipZrtTCCshGJ2ulo6qEfVVOkTlAuLvjT+8BI3jcogQrv/G2
jlplSk0EkWU64w8YN7v7O3snSKLlFbctJZrnocvjoKW3JOYfOjnKlV4eZkTc
7S54HVih9cyQyMs79i9U4vuksDOXBEPkRFeKZ2E9xsHw94vX3mCm1daSCtiR
I2KET58Zf4iEtFzaGpdNPi0WPb8G2qx0PSo0/r66hO/qL1+uWWBh2b+33iTK
GyFWhQsQTQ5/18Yq7cXdaLzwauAg+8PFFdR8fXIRGuXUre+xUHEpvMohXOKY
Kl6AliLWAcbVoq2GK8+AnNDK3i2MMbWrvBqlJ25GHEAMAVxCVOAj+yso7Xf7
S3jMMCgLy5i2+QeCC/l8Ru5Ie1+oUUMksvFiRbdBpdfQQDsYi3RZd2LxitNZ
M71pefw0DddiQ75AsUzieEoJUqukzBEfBJM25r/ofhVelnI7ReO5NurNU2y/
DsdgF1Vvpx0s3eNA+3LYZVwKAgranKZyEvV4x7N36q0tnVcOebckTK1KH7+8
BqdL5D7jx4LevzJ/QEMnUIG7WblszBCcg5LZje9g+rYUteHa4ZrWkZbCfaYI
BO3aZWal/0LYxIcWYpJHVsg/l+KjB7gH9aqHK4VdzYIIyS1sOLle9dkLQh/L
PtMcgnn5Hk/EwyOMqLTLbVzyN3KeiCN1y2m4j/pMJyxn4eLAUthtSvC52k12
MOjZ89CDJttZ0hO7o0/5r+O7dTdQyrcIsLvvaVQVcdeXS7W9Yd4IfFTI16mN
mVI+CHon6yKUYhx7jbi4f+cIk8fqb6zUdgiPnu9/1uGYhK4FLOfJmUOlPM1Y
bPBIvcT4mm6wTuDWqX3HFYBVr8RKJY8qyR6rlJYzy+D3bNB/VSh1IIcOu5gi
NwyL0TbioyKAqCbAwZBGXhBNi1RMjw5kWzb6BaUxaZn7BElBqOMRKRxoIFO7
qfE09q25/Y/fqM8dWaFilGml4Dftuk6ZiNOwHWPtdmjjgPSjkugb+tZxKYHn
IzKx5tDtahc7JBJZ69JkO/vmYVjkNfRVxFfqN9oKoJ0Ii6fJvSO8Hpi52pH7
4OumfMDANq295hLPh6x4G8dD89hQ2ITrsP5qkPJ7qFbvEbGqZRZusn/2UIs1
ZlkO3gNcS4IpRCYzCavIi9ibTOcFsighzQaLtd4YeRfwsTt0VCfeRIQOxdaP
RHisWH4H4BOoFhOeXJNdhsWt5t6ymAB8CQIREB3zgUgOEfVywVgUaNbnQQdq
qZMYv+F24UGm+lPdpFVbKfvjs46wt2Sj6LVneC6OnzOyu51Ar5z8SvKToBa2
O2omcQElMxMRhufOGLKlgwziN9Yz1g1Y4Qk2A49mMPI/55K8QPFcOT9YCSyC
mu/z+AkLQFgZU5+fauhMKGhrVYJSHF2XxcHaLPoLxQbDMzAtYyXBaiTOEIhe
8LEVNFhJguvv9uZP2d5PL6CV+QflbfFQNhdRutE0AhZInz9p3xTEq6gnatPo
j4oHUZ9A1kNAPSQs7VWPTuzX2qABNcn92PWnwjcebzHn6ZrqRyf4C3c22Fb+
nZGlQQmZUiR8Fd8W+Mar6IcknkahbSWGN1hwiIbYwIKJW2qM8SKzPR/oHT5U
Y9zvHfRdtM47eYNIWkmiwkrj9pB/9yFMjtZrw4TWQCDsECkgpyQPO2VDsaco
qBm0fYeouVOH7c4NgD0GmO4YhqIs05MOSmeNADP+H/PDc3VZI419uLkwjxh5
orRIXDDN/3McBnjINcwatg50dq6f+YgWclygrzJXuZlNWnq0ZAC0WIQyW1DB
aXUJ5XHwWQzZwTO7FFIIIVLJ03LZ08W4l4eukZu+vbjeHS7+5iGWil5LtCTK
RUbxxGtxYG2BpCOno3lNpt3nQHZhPkawjhuwzvy3GBt4454xB1z78grXgpoq
FfLvgdtqUHTxNIK9sq2seSQDsBIJjodidW6R0+pXXBdF7vvlZGBJ5u2lRMl+
JePm9vycXN89UxzLIqi/NyZJAKehGWHFDT0sPz+00iSP82vGex1o5AMfmc5j
fIbzQwyZvhh1M5F5eRfRr8qkqp4Xw1FmZrHQwzDtpm9M8QjTfxPROrk6nvUO
WvI4Mflh8+3TVZhUfed1AaVPR7qSvrh9ykAO69ejTa/WiULKlrqOpSSKDwi3
7O7xu2Mn11K9BnsPolHGJju9GSN4kYm/AqC+cIWrNnVM0dXhnN99CEuSR+rN
kmmNyCy2KBTKMmmw0EdOORBhdiy+xIxjJUkYxHt7Yx4OW7wJ4dA35LmgINOZ
HgQSZk0UrLBknvuTqdTi3UvSCzJ/V7HHRrCkDT30JZ/LMDhpHe3ysBPKaiZs
DU75M/THrocDVclqvBvJJTElTG8UyIkZF2/ztfLBTOQf47FGhI+WWTCgtNvA
iveJVsgYdug+5J6CuWFaiMLawAHHPWETJlFhtJBwkXOlQxrb3pR2nV5zInc/
kTpPFWWw/E3QMiHhEhcQ6K/vcdBC2i5mxBviJcDqx6D/eKO98Wh5oVW0wcoC
Pc9lCSAyhY/3D7xfvYYuX1Dn2RmqGWqUif70rbYJhcD9UONOGPfH8ogaLcZ4
XICZKYlPqNLT4L04z2wwRyhlv5XZF7JBjaKsOTtv1wRHTe+VeecSNq3Kwupq
hQdUX9IkszRBdh54QITOW8TRcOxVTc3LPivE7G74kcp7MKPi/xokH8gY0Fc4
6ze9MaPJtjRCnC6e5w52S3NuFDABxJQAgHR9jAbeS5XFzPsUeiMdPOssOZss
Izb3g9Mq87bekGVQJyn7q3/XPkL3bdgQgHjkOd3U4GCzeG3/iQV8+nH5qMgj
7MJCSVbNruNKU+eodzqw9N53W4foLbfBnww9jM8CnMqqDlYuaM9i1ZGmLjmw
hR/beSHdr0l9+rYnqW1Yj4b1COlMBe2PJKRW2NeNz3Wiz7M8oXbfwBH/idEx
Bh4UkuM0cYugYqWO3DeMK13DWKiYr4IHNn500pooFZkHjUT8UKr0To1fBFM7
4fp8nm6ekWaycIpPmt97UEMokPlzTEw+XVeZuK6viuXtgO43ZxiAAAPnuf5o
1ImCxOX6DEcnBdEMJSaVkL5ZOggdrV1K4FzBv/MfhzpeYiHqeuUSqO8ZulKB
4GSNWvjMx5hsdKfXbsydxDxogn8kliaNXGTwV907IBPCUi7b8jDJQv/kBtE4
nbbd1dM9gpzVEtubfiTjh/7tfuBJVJgsUyqKSE4R7358sBbi/KkvKzBtQqDM
P8ikFKPuj+4ITNLb1QO7PEB9D36eG8mtQOBpZmZbji7u0wIbebbTMA6xELud
MSW3wsRIiXkYprxJx8jP/Tmtb9cOsvLApmrgjmR+KBe3ZdY7R13ThfefDEef
QaqBO962zcqLtPSJEB36SRbAVVkE8l003Gs9IxWGRxXBJGtuICG+yudrkxP+
8AxlcoJROJAewpvMnDe8ohcfBEPvB1yKUhoPJiGqXbvTZ9Z3q/XEOE5rWHjz
aBejY2yXoeXnEBisYtKkR0jpvdEcFs7nLs9bXDHpswG1afDBmUHzXWl7mwSN
h1OFv2nWU9ogluPsNOvbEG7bQe+J5IW9jEuFGbXrISUWfJ2cC8iJZcfMXKFI
JQ2tYxMWijnp4O1QqeQaqQrY2ghSQLaEcd+XV/QLxr/rP41wHR9szOR29STm
2lgcbp5d1+cNc1gaaECkwjaRcM5hBW2NwNezMWht3731z+M7ULiX4M0XVbtI
ONYYplyahdqqr9YSThhgH1jkNj4lWukBI7Af3SHfAjYAxxkJEsQl5mF0B7cX
Q9e/zQ+j9Of6vZ8Eh0k2AvY/lICtk/MRXtVJUCU+JNd2QORlV9q1ADCj5lS3
fNXWUacjLVXtUME1ebaqnDieU+fp95UyaovDkzME84BBnw86i5O+e68zYKrJ
ibjWny7t6HHDnpCedHSqGWp1UPLcKlbsG6yHF/WgiIp7oSG7pUNgmcoXNDEp
FJ0aRT6dyrEwndMwrnD9qDpyUq8RWhhN+Alh4WbURUDPzSEY+X3eaMagylMj
TlN9fnIOWJ2n1ujHMydzQZDCSFnR58H/BgUXALoLA2hD6Rv778nnaLbhiM+n
jxABXFgjAOhNtl9aRBci53YSsRwTJjeYoiiEQ5J+ccD5ExcVJCx2mDaoCeoK
z5ih/9ynAeegdo+CjEFCsMFgtea1X1ACaDpNoQc4V2XRG7balJbTVk5XVewG
17duNFc4nAlrIDi61NYrbpzwfzioqv+5OF0uI9FDUzWkw2tgnKrRL3jR+nNc
AMULKo9+spZRWaIFMY+i3VBr/EdQclWe62PjQm4G66O1yv/2JTiOwxTbgdKp
p/S4hibdhfhsuqZBBsl5kY+H+BrmhEAoEdSwLDh5VZl1z1hw5lUqUDyScEeN
hNUru+3z7oQeT4Gkmv2snr21YVS3Bsk+FffziTxNmjQdPfKQNkkd7sx3T1VI
5ZrfeXsFibL+dQ3JLAb2ZARCNo41Hodusi/eQ+i8T4elQKZf0aG077OLpt48
uT9ZbhJj0QZU/ySHBpARmFOdUFKqGU9TDaiIcmX4aRt3nZs08hQVsMu8Ce01
81kcx0YgizrgPwQdVfPz/wWlf+s2JsjGyaRloEuUgMxu08a25QSc5jvE19kk
T5Khj3Wiae0mmQmzn0lzjby6uU9fuYatOeWd7wRsWWeMh+UO2LGc7yW9abJZ
UrwhvZcOatQZ0M8dTZbXs1Ykhu6y9kHq+nqeIfdzSAFa8auug3SGeTeC2tRr
FT6R3GGRW5wbCMbXpSg3f9t8zPnwPl3rkv7cK0271RbjSBehl0NilPivDQl8
X+imSnTn4vtHoqwNqZM3nqPAwdlmeXS6uGBgdF3iyL1EDPWF9xvwFX3Wxfoe
YoMusd3xBoQ3jbDRLR8wD3/zNGEmn1x0pZZBeNp5dIQ+K/bAdNEuqnQAK8xS
cOn0Y8LwbDSgFekHLwe0eH4mwRE0JTlrxWBfBusL4U5oU8/L5dL2Dj26chrH
c1O/u1DRI57aiaFH4rh8Eml5v4NNQkqHmdIQCbE3ogTvg4x883LqgZTfKSOx
hCqOzN+7r7qjBwAeOOtQzqnc9fl9RazwUun9JBacgl48t7fyFBVtVGSTsgqg
yikljjj65VmFBqHqURGyorz5W0yJt8+tNrwtql3ai8HaIHRDegv2xrRl/qTb
fDvotpYz1Mnji3GDs1P4I09tyVm7nt/CAHqaRCKz5Ytir5ilAvJvcWnQpBLn
Mww8Qwng5pb+jxEBZblGTOTKB17dn6cw0zdUOXD+avIakfwa+GCpXTGuoSDq
RstnD9J44q7O1eES3jfP3Pl7ffMf0TwogRhm5UeCMjwShhgu+ZZu4f6LDJVm
xqMG3VGiK2KneahGSB53GhZrEa6hysO/lWOOZxTxebiSZ9AqVllWhlwcqmOj
VaFkJY61Mha4x2HGYiEBAMDmC7eIiGCFs4Yz2CHqMUjdygtf3730ebcF7RAE
pYH2eiMzA4jwQPbK4xf5KFU4ip/8MDnp4iO6cSjuuLCAyMBPgNnLwS7JtaN4
ZtqTtlK/Rzc/Dk8W96w0u+/TnvrkV1NFbgnTOEj/k8VYQUoQ8hNFA4M6pfkh
FpPeNCTLe+ucsrca5NNnlWKJfEAbwj+wRM22IiDj9t0q7c+e3apCfgF1B4bx
yGFp9sfTSIfNVpCN262HcO1esH3YIoD6eos8Ip2TndHn+EFzPer68AyDyZQ6
BKHJp0Sb2hkkBN1dLALwCsqLsNGuK/Sxda6AaiLFwBHlw7EkDgG1lm01AOzA
Dur1I8b+nG5F8zTeffTsKP4uUvP2kM7VwwrzdrLrhfBpvXWgC3Br+1duVExL
pSFIgyeZWy2n+Pe+/1FWXukdtR5Bh4vBekEtuouE3/YGAu+Nt5+YSJugrjD9
OElcTfsv/zOP3y96q+xELAQdSQTEZkL8c8rF1utNkvEy+CXBM6k6ejJNsqte
UMfuziYLvtTGTOW0SgrPJiS9oaxoLoNjY4xrkbm4Hj6Q/PRCNio/f//7wh0P
yd0xeNNMCzAiqbV0qAOBw2us2LW4a59RSpOurcsFmi/Ob77nvQf1Mwxo1w0Y
jeUiKPOsvaB7y1dfzP2FI8sb0L684F5UtZKv9395CHq0sKFn+VCrkrzoh+Ft
dDosh69RTwape9iWQlxl7spp2hXvoCQbhB6LlnmFG27cI02TMdsY5s10DGhN
WbisTLcOH3j7FpotPY500QW3wxTwyzEPasVwUwWZVMvI4xnb3asMsH4osG99
enmZKxX7C9vx9umrx/4fupkAXQiXLDsmu8YMd1Kukiz+0r8sKViuU35vklxd
EiEm4GRri/JQNiyppYvZCCaUZppsuJlziyIM9LudEe9enE9SlPVFm3d8nnGD
mCxwHeuKUaWfkAJCei7ht9jVHcfuDWltATSErtSdjVhDoYcX+cxQzBrkY7bo
mEZOtcddXBAUL7gi7WErhjFrP6LudwpNnvhJl1LrGM0rNanCMH+tFDdXP7dg
dKzOPW5CuDtqFk5RS6BMUUqii1KOxV8XcfghbWlJO69rNe9CvZU0bluesSnE
/2k3vtAFEuWHI97jdvNFrKoXszbxQL1OYMuWcjyEqlUKUob9kBFhfCXfikvv
JTMqjBqzSsI1J00MUvjFqS8eUYGuAQzuzjp0WR4UVfm28oDlr3cc6/BBuBhi
7z9vi8xx602C/e3/dhdZEtfCNWdW+JWOcFH6zCLPIwhDpMhetwdc/qdWV46Y
EEYBgf9ff4RXcFQgl4WDGom/uGzbk89OHbkWTwM+bjM0sa7+SQBMkYYU7fk0
CJPD4F686y4uKi2gBwQL8IcfDFNeN6f2/M1vSvLGra3B8nOjRLvX0fhonc0i
U8MZYRqd594cHPrT/KNfcNGd6fPvYWolDkRc41fGqq9FXYYLPJGR8So653Po
R+II1JztXcJhL8YTE7LeX/HDEK7yJ4ofVX4byncJC0QgadW9LVy2QMyUSHf7
fw2yGKUMwkCIVCMlvZtgLHtjUdymBz8ukxugFOOmlV2ItDGxmS/TQpO699Uz
A2Kb+CjzNEiZ5zk0OcXLxiqqjyEYeeWKGXGVACeemCRTNpay5Qwx4uC8+3VN
F8mwoJH891rfjQc+7UW7r7uzJdoanKsZLgT8V1iVAdrqwN18ME0MeFmdnamH
kLlJXRdpKyPETMmGW6PfZLCAV3jQVN4EqjqNGn8cvmSbtFj56U0Ebq6+snWT
QFR8WFkgG5TfyDFP9YP2MmX1yuHfNSnUxWvL9oFhzc0p+BRBOn11lzRXHkw9
3vHvQ0TZ/Ir+OVsFFLR01Fy/Z24iN62fsOgsnEvcNLUbDSMc85bg87yoXx08
f8yzlyizhSF6NSyBMWvxmiCpLylbLuw2dC5bxOs9UKjhMiYtA5hcfS5YUywz
A3FzSW/SuLTe7VxNkOv1PkqclNANLamMlMtWQzT7OBVj4z4ytkiRingrUZFh
H1FkPX1eUVE8tyryPNnByRL/myBujT0Ip26bWra/+Aw1ududXOd7vJoyv2PN
NtHOp7Ap7aLoOH+zeeTrze2NNz94J1gA/LqzeRXxGTDllOTlfr8vtp/gR9xr
1EWsRn4naR8jfCQ2oOWHLza/CLLYQgjTkOJci9cM36S2zsnSw3a8hlyFHMkq
DnvQyNpkU/GnTq/tyFv9mrF+eHjNZSAgzURwi9QSSlqxciVgiLWNp0Hhw8dh
vTQIJhUFOi+PLSeLjTgzde9zdKYvbMUc+EYPoixxBScG0MJsEm82C38EcdPV
wRxtsz2VPfnGfWDwLAp1Mn219J6K5E6ssJl+oLufO6PjdclMduWaCcS2IV0l
35jCZ8zSfWaMOesOnN+Ab17hnlkzo1Azp3IDhXP8ZGHprKwyIc6fEFBdqI5v
l+8CUodj8N5sTaA5dfaBDS2e+DYC99Tc4bKU8TVwWYWZTVz3OFNJ/vyGtz5P
DDYaZLo+Jc8aYlAydm0zZzHo7aG77Xmv3sr3oSBSQEFM/9ZFe4/N0ptNn+R8
d8GFQFYJ4qHXUirLBlz08aJ5isf9F7UULWJ7YSXP5DAagTtRKET/ZzWzEhAB
rUyKJ/OHCK2v0mnk4KmdNXCwaVYhLTPP3FV16VqzQnfHaKRf31jQF7KhsTX1
lBSQ4Fl1Qi3iiol5vs6cdhH8y0sLM3hFV+KQAB7kqfuaMgN1ZofrBVxuM05t
VRgfDJQCrcUja/sr7K2vU07t1fZC9XWfZg7JLECfYYcI6nFMR/2D9Vjnk/Yp
kWA1/bvhq6f95NB0Nv0p2n4wlsbK/ATlwW9bh/BMMDY7cSGQJmCQFhfCYoww
Y3s1bxA1q8GbMZSZAR2mz/BlajD58C4/AImJNxmJUjeqqYooRl330pKUtw05
u3QpjPhYFAfpKj7OS9P2bW6WJmaiAecSeGZkXr65AInYQxw4G0Jjba4MeT7A
wUnjO4bUVnLPXoTuYvSYR57UrsHOUEpGGVpRNFH4Fo629zSs/FO1kPLgMuTO
IjZgBi/vxif9mlJHhNvpkPNUOH0DNtMLFpBqOkcqYEVAMuKCNFvAjv77xQls
Nbed6XlmmpliEhkPF9AiENOEZmFejEOCCnqfrJisPMV3tvjMbVgTLuSdVdcf
37QlmXm990yhIn8yp8ti1TQhJhdX8QrPKzm8Q/7lr90LfJlsIc35uFathSqh
QAXCoR6ZSWH7BB7DMvFBVc1VhwRhnrDjD14Im+yQH/qvYf9aLCUyjthrfzDi
nUoNUXQxNQNTcLQcN8OYog0g0rrNmiLPDdHStNwdWL5jWLUKclXGVp5CgUm8
VaFiJ9LXo6DjwVaGde9j1v60iyYwq8yw/uYmwE+IcZZq/Eux5lKGtvBT8dft
mPxJyVk3N2GJ/nJWaa0qRS4/akicsAqTj57emhvQzsFFBbRoIzWfpY0b/qa1
3dGI3pAtXXzQg+HwwGk16wj0e23p+EVzIH7hx8HSTlgx/wHGEmSJAXMSdiFl
r9aFqmdFJniI+2yJVnQhs3llS8PGSNdPOSJlmWw5lH+whjNS9Giz9qqVmWyO
DR/TZsGG2mz3hzKth4qX6TSSJl0fkd3bWY2+QYZtOOtye7eIo6JHAr9iDdKW
PrhoRGCO0b97swG6x82xW67Jm/Jg+jiK5LFe+ZFGQh1TyEJlJi0j7NgQihE/
Ovz8en3i3QxUsjJU1PTFxV029cuALECiOFskRrhBDXnFqfeaq58tWaL/k5RC
8b248vFhnXbxYoz94Oru9iSrRIyWCY/cbfAsT2Oe3dPeLUOVPMvf0JFFFmbv
z3rk64o1jwzigD7XoCGOK1oXP/kioO2i+ceipj/NEPxqyoR+ifsecxv/Dz90
DMJy1QwhqSQq86GCLV9ihHuo6ulpuHCEBrdh0qDz9YvKadu1aXkdcrJtPhkq
N8I5GKcVp5jV98fvR1kUr17fI6XfrvNNTKrhiIf3PCA88dElm5IrZ0byeGYD
nO1Pxm/ZPdEMkwPVCIus8134DEV1AUU6skFOKA/8J4ubZwwVsmSOwm1v2KvO
R2hNO9HgpqIkDjysTJfCYlsOnuK1W9AogwL2FthitsW4kcLKncgFzoYfhPlK
onAu6ta3i7CfWmKH1bUepLMUVCSppWOM0h5NRUDLFuH8xr6sUCNg38l77I27
P58/KvfUaw/CeZryHs+ehhCMVYZzTHgT9eaFmP9KhfPeaPYE1xFOcQpX6ZVU
iWspWz7wX2fJmVbTWTB7Dts55uSR8R+0DaK5eo8oCqOvUc+TcaNzS2BLbExb
dCNYMEwCUT1VrgEw/UST0W7hrp3XnShJMV8jyFBY6Snmm9JO2cwZr5F4VcJy
bl5G4wA+LfwQ9kq2Qs4ES1nvxT32T8/P1+fs3D7WJpuW4iENdCpBpZSatWnh
eDbEnhRtD72gSPvHyzDLIuOtMAGMHPrNoFex84RKHXcp4AJzkgxLtstTsBOg
g0EbXeXfTUJDXZI2QSV3v4DEANaRMPLZOFfhtdKVhq/ys6M7qwOlQNRxTz/3
KHGJMllZRajz2CZnoxkjiIeFGs2BaTfwHEmLHdei7QKgZI+GGnGJEQeNidvo
PW1mbtXNWcSGNF2nOlq32tbxfjFiGEgbCwUdsSoynnbVZw7ivenE3GuK4Bfv
bVJAy5oziqAhELNixYwkbg+9Fz8WlggvsRH7WFEU2IHacWj6xbVz894QXXqc
Y0zm06+cOIvni/AgV50wuVuhxKy5yaxMsUwwMOswhgkTrOM+jncJh3lz28A8
SdyYJFr8LlELsiQYsSlpJ29dgd8RNpjbBUkQ+CwXWWifcdfSTnkNtT6QiViL
dRs9y62OAg0Lf3bP33/YbJS07IkNrWSzOr+Lc9HPQuy9/28coZ/DfUkMSs3j
rNM81XeSpVJVFFjolr7NwXxJd2yc6Oh2wrz+/cKkTCYqSoSxWVXb9PYFnN8/
0N8MXJcVofg8M9W7mrH7USrcUc2lZmDwWJ/t/MKG329t9FM4qGpsWhfA2prX
Euc6J8YMcSZl3jSPFa14u328+enA6b0507nNP8v/fv4NgjFnQe4WOgXRuMLR
i+vI2fFJVUkiy5GDH33ZgDGyxQgzjRs/4M4CjkOTSLHHkmhwXxt4ucrS4yhZ
M4urYqX12jjakgI/RC3OggTIIN16g9qw88DyghqTTLg0e0eHf8rjRd28Zvyz
hvmEhVlYWGgocOuheCa73zDxeuXoCOFzw/mNBOuD5o5PcYbY9NEQyM8JNb6f
Ffciq9IjnQkrbsh7q302NCgUI2fePHiDK6SUDlzhu877FfzXWkiiG+MABUiz
2Im/EDyp6svEVlDZyUa1ZhB/tFM8FZbBrqh8VnBHrqTwyhCgkkzSeRGimcFq
PuknUKVkro09rKAsnkyzsca6YY70raa3n4Q+YsNO5hIUVapOUWt0vZDzWktL
lHi9GWIjhzxFjGBwqxsPY+TxUkLuSDmO7k6aP6MvIOJkoLkn6QCV1ZZFlRtP
03D5f3zgtO3KgNfBUaoYFefV9FsBnb+zw7KQ41/J10R2GIbhJ1htfLihM1t0
M23Dxu2FyvJkpfDymxP96IpeNAi2tTxDLVDkmyAlZHwa+HgaOh7Hq+q39UXL
vUE8TycTN6npqGC+l88baUH3olm1KrPFrqe5EV5Rpksj8C3wvFBhjZQdNCXI
lwrwuG9RsC+Pqx9BwRbB6l+cpRCa2Dg/VLgDHqsBhgtUwbX24lhj1QFIkbY5
o7ZaP5bBUCcm+IffLEWWogTMOMnbjsNaTXS96fNtpN/PzgMjbpTkrjm10y4q
EvpXC0Hmtmls3GsvBFAl7bdti69mT1UaT7lp0mI6AaL9NU2Eio/bVeyCFPae
BIwdRW9pJkHOMo4GPn+eaXWSCJ3QiFrdhTWM+YgJftdD0nlYsTtkLFrK26Ui
9BL+wE3/yWcNZdsO8kOQwvDAJe29tlX6p/SYyq/YPyAilZuvEEnfsCmzN5HL
TPOz9Hp5vCmNCo9Db0c03u/r1MIv/3Jb5DnGBcKXxdIenszuptMWucADq3pT
vleZvCCxeYWkh02RYhgesljB9ZrqhjQQUSLLEaP5zlMSS52YYsK1f+wmLNSi
LvfvZBIFwYaFvbU8McnMln+KZJ92P0Ad6PsvQ0UfeccDe7886SDfVTX4ZTK9
UhoGz5fZuEAy2i7lJ8Sms7pxT4kVgz4csTC489yAE4ptutEdg+fZaXln7i/e
z2FHmVJRtqMFHV1002rEpHQavLSRVk8YDYaTabpwZO1YQ4GqmKlglTId1qKS
umlsgqvR9Re2JTerXreY1aU3KztPWOpnn3ewEWXvbuDqttC+aZUfASUSxToW
fNyTIoGRD4Nt8hlDJwqF7CL2GCuWCr3aO+52y0mV4bSVLqnilwrl5a7nNg0B
nF4Lx0YMdpfkY086fiA2nnhINaUdTTu0kIuPsJdJQ66SWJjqKyhrSYJb2vV/
C5DAHF+sovOP8cIIn3IahSwd5b6ptgWixavvv7FdYTV5ebbGxI6u8fMYoR/5
QAhrg+GcAIsSztUBgiLN6xBTgxKtxY6DgvGwVa4u3McsLH0UOr3Rw1/p8/o8
WHSobFnKg0/KwiHIftFXXWyaGC0YUDRpxbqxsTGBYoIU5ANb60RZ1fS3TtmQ
gaXT9Dg4z1lwGnigSQ3e+qaw5iRUTrL6NhQWUMc1hVptvCZuB4shrxReA4cB
XoG2VHEd0PKcnvfSTnatQGarSiEIsWx8EaNavOSHtjhM8dE9s8Frhvu/B0RQ
RvPycjkJxp7/i9NwS0+5TCdDZYPa3HSjJOCZHbFIJt7geyt+s+6KXHp7AxqP
XLj92UMtEmn6vf/gLvw3zCs0/fxnXJAss0+rwR5aiFPwvDjKJIu3Uovhja//
tqR3yTWeb4wRJJWBW6PkYv64+rM/dubxGimDFnLqYLe0YHCxR2tueX/jSN7M
27FiPZYPAr9/6waLgKHga9NwyDBAzhJowCpbTyO+lzI0ldAxXi41WeU7yd89
1uVnUU2E11v/KAR9FYYRa/UrcrFJ78S9N9f0VP3c4MHzuEwquSQo4OZoQ81B
OzgqT0d9zg92gSJdpFUqMZqU7sAzHG2yY5BX7R+BCoHj8xYSwum6X8yqjDKS
/J1ZGTPmck/0XRX3qQHcpVE3q7uqw2oTr1G6lbyllCUAioSvaolwSvHPe3bS
YavTDKkVcxJQ9vv6S3XEFIhE6VjPGrKD1TezH3INP0CWtGPpbTvCwXNqzZxI
CjJbnI7p/MyAq/wx+feYt+rVBgHCL7P+ZSz+B1iG+rFW9Kh5cwFZVpf4hE1S
tQafScljzS31VvG1QHNS7yobP2HkF2SQeCJGHIdJ/BJdylMrcii075vXLDrg
CfuUOjB4yjLY3kkmHFA4nn5M/sU+YHGLdQ+DpME8D/XVQAZPJVSzBqbpf20o
jHKquti3xGDufVVmOsjuXkYN8rrwNtSVkbmU8l1DGLEpOu4SAwo1IuM4kTBy
PsqWVtfQAz7aT58aqgTZ1CsysfhD/Do/5lU9bzg49Ec8sp/kiRjNSjLe/daM
c9kO9iBVYNiY6VU0GjQxe2zq6ImIKPWg9NUgyFw0N7vh5qYZMEeiSfbtZWHK
VIPkbxLQQCDWOKqZIBYhBodzZnfEFksa+KIRju+z/e9MqmJzbvrMsxLlV4M+
BNE/MsO8vktjAgJdZ1Ew5N23jFqWrf2EktBiAGdGBfKcD/wQQ+bLyUuWBUR+
tELG+LK7uzJ2HM7Iw8N+JLKrpj2AUG/xc6bD6K/wrf3DldbZ8BUBkMTvsoqH
TC53DyucxhYI0xSj70sKbMnaiFh8HWh98oxLY0zaoPI7gX0rHKvB++H6FNbj
nvh1lqy/smRX7u9GB97cZWrp/1pdNwArIvDi4TB4w6HFjnZNqQxDIjAZI+LY
pX2/IcDfytHn3/xMhWMEBWTRO0dWR6rgXaDu3ZRmX/wf08AiHMqQu9saNaCe
2SPgS7EbnO6XXtrn8jCr6fJvEWPiWUvamt8JOusa3vg+MbhrvB6gpP3Rjky3
1uAHtXXSJ2xfHpUwbCKtnqJN4IFiWTsgjcwaR+iZrFMJ1dZWC24CVSTtfrVY
d809k91A5/C7LzL10la9VF9lNNF7ZxJDY2FLRij2NVUTY9bHmG0BgO9634U4
+BEpcVCGBsGk0i8GRNzWclFXTMfFxljOm0pIaYMnoPBJRqzRf461uTTcPXLm
LceCUJTha9OFexKQW1JhQjGZJLFsKFcRYLdiWGPhrDgczJen4U2I3NVuGlqE
zSvvu37BFtbT6YuWk3rqPSbFe6eBtcFzVPP0quOKl2YVT9+ZTv0LgMCzRS10
o86N2APEGj3A/5ea2iHVJEYga4/HaWNwe8oZHRMUJj4Q73dRb8EfCh/HDxZ9
Ur17jF2OO9zbUnT6ILA656JyapD7+jrTQvVnjKQbzSWemvQOTaDwNOLXv+AH
WKvZvOxd/abH0ibqi//18CklQwAjGPFMPKlpNo6M698l+ryhkPloy+nNbRnw
wX6IkmWU5uEz2YbXw4H1uvdMETXIyo4OTiIN50TZFwmLcA/IKVA/O1LbRpH+
gaCsRBk840nZdS7vdQa4KiamthzilOwkQas/2A9ZGgGZPXH7fJWTsMpg+YTJ
aoVr06w/app69b2WFQwZFRZZoTWIul+Si7e19pjVyBWczzKuWGKY49IffiTi
2RAPM7ZBHu4LOkNzw6S0gSiz1DMl77yrYbq1N/jWAJ3bqETN03jcK3jjlAzs
JEZ18sgg7G5s8Wv8VgEwGnlIEL9oQH8DfU/pz2z1y/D2TPygIFvnHAxVnBkm
FZK8Zn/emEch2GXpbwydxUGG9ASCzQnDBIRi+FtaiqlJ5EHd+X7pptu0tRLZ
dKzWnIJo1pFjlpXk2QMMz96dJslC0U1/krNtvISi9xK6cb8iH6ON4Hy8IG1i
/RhAHkCkVUCOMqfcamqvUQ40ZIFvmwd/KWCqpJ2bQ+hcU1kK04KX69x7dO7q
Hfl54oGWiwOjvrP6TU/7ucgCjjy1YBPeeCLWOvVFAOwcqET9nZNHesa0+B9g
emsMwJTf3JUrLPdEAM8F1vg6r8vnKd8SUpQs1u9ciLw9OECzRa6ayd+ol/Mx
0RPhEuo4bCsw/BmxEMP86ML3wmkVxMJM48thrm9wObb/QGGA5m/ZG+U1Cnda
Xjc4nW+7Efjd3PKWxEQI9CkONgsUr8CgQGhMx1+QU9cxjmwltIT+mHEs6Rk2
ZEgW8RPVxOG1kqRy5wc5Q0VN2pEfeZyzDWmVRQC7roMeKtpFmsA4N3dSumSB
3784FqQ5D44oi9Tw7nW4I3vK31XmSBUn8U9vCpGkXm5/yka3+gDGUqpwAO2N
MklUrg3+FOCVR3JZoNW7S0N/gZW2qvxH0zxsLamnBf0crSeS6qv98dDCggZp
z0VWe4bDV/tBasMSNRRBCZsdqkUgPnDAqDN3S+sMrj6uxbHXeOJQAshJUUrX
GuyiK6i9rl0bw3EvJf7Ep8e+AyPlivrC52RgnNRozrGAWd9qkBt/gw/jZ0ZL
uiG4NJOfgEWCS9Q5E20mx1Dr0oMxpH5E6q6mZsqiPGVMs4gdhOCGJ5PN7L0K
7MA+seWOYaqd6dnr/e4NLXklAlOIMtBnhH57uxfwZmHu+NgtnWVeTO8No9my
q6aTRfBJrQyGNkR5+ia15YRP41cUrVe6BLRmYvY2xPWCKIQNqmojii/60BQw
NUdfpwdKqEEFTgIESzmR1zY68CQyTMhrenmg3uT09FbyhDQpica+IM2OxX75
OBuXiRg3hISgd0H/tmqT8IAeB+jdWrCqEtpObgMMW6fvWIWF5RP3HEiNTqz4
/jpRIZK1Vzf/6dDfrYMoCBp5IB+URFL0uvzuiVrTBlt8fbZtbkn0nO2U00Cq
3UR2g+gOhJYR+OouDoqxgfh9g0zEuO7CiMdqb2XgdUAQksPRN7F2ACy8dQj8
gVe2yZkpUpQFsPmVyJPgPzPiVOXSBe0tWirczS34DVCEf5IFifJ2zYk+XWBG
EQ+89o6urOu509IbK9/4oBUK6+b07cURc2kvnAqdIxiA4yGX4mXhbHY3iFOv
xfrdKlqEoy7SN0BjUSeL2SmduOV8OD2DV3/nslUp+HwZH9EGKQuagf2F2XrV
Zq7nkD5wIPN56snhi5SYtz+hyjFwiWJ0zUL2LxzFDKYh26garyE3v5YC8HBg
07BqZTBFkKVctsHJ/1Qh5Yj/dfhPuFDU4o0sBFMmT3e2d3SCGDldmBjO07MN
P74fqn+XM2EMp6KsEpJ0AgJYL1zERr2UV1dWHhIFByI2hjEXZ45QGBocrxAx
NFjbYK2XeO3xm3EcCLSvUMMHyRMcHJcNtmdnT0/x7LR2GQAm8NuCZTjDX7PG
Aq7Ldq5jyGhMAB+FZW5JKDt4+XRFN5UzLiCaBoTYc8VFy/F9+EZ931+Wpiam
dVK6p0zhhHC/0MRIImaCa5iU5vyVs4xFpQ/TVxwD507NP5tbrZgYIkqmU4+X
1qgHQLc4ZRj4dIIc6diN00EggGXvk8j1LUxm0YA0JIbm5HqU8sIurWIw0UXp
wOKwsw3dOeNQv6ei9LXE7fCANgIQqBMPirKMqhFVyoD7E24YHrzhoKs2jHoK
MBgP+LrqmTT1aDhT+2GML7Io0kQ50GyzVGgfXBus+qePE+oljIPVUkM8dFj0
aovjRwbwPBQsBm/ZfbJWRfmfw9gW++kAEVuwUx3tOEZCjTQ7XneJomgII7qf
8aEN3dmXmrHAvT1v0Ya5Lq+TzIHYXJlfPoG62B3RQ8+2XAiEDcxerpLv/Obg
vXTvV2IVItDxshKARC67szxjltHqNQHR2oPgX0p8x5mA29xmFSdH8uHO1qvB
9jgP/tlblILLm0ufKQ/61O28KocMMM08IdnGmvR4vQej7YN1cEKhn/20YunR
gNdqpoW2Z5SeN3bf6+/8RECLkQ1rMu7dq92u2XNxBeP5Cr29Rt3MHUSDxP5/
LSJK1Vh3aySlTlV0NMbQMxuAPuH5jK346stCKsawKV8fgD/4wq+E1vGsoOVM
CjwFCnDwPk9OPnUUkfhQL18j9HpsBqwUho2SnbDRc7sNktqIK6zmDTB7sACS
mOFmVNqh+2ed7pR0Bw5NWp5fCpA003COslGEa96R8pqeAXXJNkaU0i3yEdU8
ZLK/ANGI2UAzcTaE4HAtpYoF0TGZxgyaxaF4M15dv9t81xzNOLKWfn5Zc8Ri
JuDG1g1l6X0N//YjVr6tbP5SJk+IR8liITm3rC0XQWp0kIE+uchcuhwNaxmd
h3sVeMPqpntHc4Xff3zWYRgkw21/+2dDPrk3oKOxteSmASOF0atqK1g72MON
fydr9eEKf3eC+PyB6BgLZ9Q6d9WsSpFaEaJ7jCXvN9mXO/qQ4/SuwzseoI3r
Siu/k6pbnoYmS9WsuxLMgTR9YYjAo4okgqOzdZHXBDWftVvpL7Zue1DTYQME
jmPB48polIEo0xKXBBq7+AQkmLyxPsLoCmML8JUZXDiW9xlh+sX88sOkaCQq
OrFgdoQME8n/2Sq9GqmFN0DPj9FGkbDrSV5kzMJGPPk6QfrwISuszeGJJIJ7
xAnm/TIIbzAraK7Sq20lk8uWaApDvAgdZRt9rSOuGwU94/nnMmD2oChzSYr9
FFSBRF85lsGHJGc/V7Q8S59Qv79kcBD0gsb0AM+b3hTxzWOMV1ioKISi3nJx
huBCPVLHdE9WhbS44wm41OUgQY103msHk0eJB9iCwJTdrENL8G4FYSn9Mc5e
jdGM/kom1cosE6IOUvoBBt1qrqKluQc0DIkix4DQ1cJe8tE63VYC/tLnyDzX
d8sa2I2OoqYeq7OmyNOu26Bpll4Vs3CbSIhPSWAZin8fxsjpAv/T3eHEFWrP
sOg3M6vXfUZtDGlZQgdfQVZThVGCNeWIMCYkabcI0W/9fh0hNbt5+24wvzuf
3d4F5L4wCRLgnekzRkZKwlGY/fMUoDAF0795AA3LYBhPBqoFTQnI1WpUparo
5Q9cM6cf2p9NhCfSiydO/Ylj8PQlnd1bxFfCrRRbEro7RJUoVtwVVEjV9aFx
ZMgvNNMOextA1VR5hxtvw1TV4S+xK+KRXe+bb4jyFiGT76XuCm/r4/Nebegv
w0lN5+Z2hIKfL6HWm+mx5xzPR2080DNq562U+RZodPbr788h5qotlgWsnAip
Q9P9xQ5IXLTnIPta+x+Xa3ubmQ6UiJQbEa436WJP8kcmw1C2YHV1Dvg9h5gg
RxJSliURnA5nK/diYtYlUR7QM8kuxnWdUIiyjq90fQBFLxiaSA+yyskE3gwr
Kni86A3Q/BlrpE0wl8ZvT2MjJaShNUJTYqx9IKsPMaKH855A3539n9uUqjzw
65zWq1MJphSE5iQBEty2IB8MbeXlpI0viRtEMR2ddjE6+OhUzyVRmBaWfqaV
XhLE0+6bSJ4GYZ1akouvNTnl5g07dDsudKlJUWXooqd1yd/Z+FV6F9MnlLHv
fVKZy91qH/Ib74LnSVa2+q7f4XMWvzFI8OizwhLK8ipZ625WOuVSHG9ALJkB
3G0JyptvSDiui0rRPRrIvCfjoE4a9fA4I06HWKNg1UsaKGSyVcBH2twhCwh/
i8nt4zjdfUoVZz4RcLNDAM8HndtqxhtWS/BLqZ7Xx6EK7BvDEM1D6K6P930B
TL7iEMUnCToQPvgZHQ+wuXwsHHlizrMpwU9XiBO7brXJ/mXdAQYmkGcFvqPh
1G+wnPDzZrzJfJOrHdGhBxN0ObQjygbYoDnjZfMILiNEyJgk5owsKCCDr556
hYVM8jSRy8jz9wwj+WFJAwVU1f+PLYiPb62md57+7rV7iettdFB72dJl/wYl
x0681YL4jtv/1mjQ9nZZznWQy3/hTCp9AgOmVMO0qgp1jlZHXnDvwqPnDEjJ
p/xSN1sW22aG4M2FlSAoxiiIXz1nkYtA1cb615GNaLJGBxJuUeGyt1/LvFbc
Og3Bct8OlWWITS5uHcVqQIPK9aP5K4DzIltUWOVuvDkLKhTAgHoY8O7lQOTt
ztmk7IuYbDsOoLsGGgTLOtOqgVSjynHieQF0+ExWT5G8PkOrPU0JqxggKJgd
j8/4Pdz6R1qiEwNJLX2sNmDwUXZ1xNKEd17W9te4f5lEXuCwtrkx/KW7KltV
ySG0uyy3IZWPFl32Ff/1QBiZcrgItJHF+vLwIpHwdUYXIwndpJE9ohFHLwih
EMwaA7bNtvBAJ5TFhkGi6MGZkcFq6zwWpiCL0/ZnVRAztW3MvtCR8ZY/3ic/
+PfOeL3Ffc+vNOt3oLVF3oBJBogWPKI5iK+1K82GS7Vjyjh38BtnvFYx8R3B
SMx87qzEvQCJ0vz/rRjYNY3ml9z+zKcDz6M2rd0ilKQ6fp/J8NpgV7TXpI7q
wHPMvzgqwxt6v3kWIPII2w3qXl7rWi3Fc1fw0iU7MaCRQO5kP/FwX7+xI3sJ
47B8vuZgpYvTPq8YXYAdGyFavZwrCzzuA4jSRIO0SyhIgOaOR94dT3rndpQ6
M6ehqJ+RR+4fInoFVzobNFXW2kKurMIuHbHLVo30BEdUMJGfDKVACnNHj28c
xlEGaHpSgSilZeWe+UySubxAeUthoyBJzxLCl8tEJIxMrxDs/JR++kUynK+5
uKa5Tz/W9LG8ndXqwUpo4+Op6WPd2ZzYfSSVp4RZRrpEnqfTKbwundfTwSLa
nqo853rhP4A5n34dlytClQikfqtHEInwTZqNHJkaCPw0Na913ryZmcEiRDn1
C/RMiCNj/FBAKejmR0Mg4vnKsJfw04ROQLo+biVO61GCr8fTURzG/MrY6q4K
XBqK1DSA3CbhjHjDpIzQZBiRtXzMuVfaBIlaADdTZeFurbLV6RGj8n8UZU7D
GC4bm67jpv6t1PoqxdL6wiKIr0mHdQpjaX72DnPKBHixKJsGyCB3j2IQ7DeE
kiSQopwhSLtxByM4tYrj28/PIH1YwThkaBiNW4NVsuuGWeSrXOUfVmkqb7eD
FUt1hiopKYYTeUlBuVG0UNOu5wj81hIshu73GQz2WzeYQmLBrPGYW5znTh66
DkgUkgsf/8BDBUUfwf8L0gmYesXrJAWLHagkpIwr3+YemTtk5JpbOrVQ5/3b
6LINo5WYLw9TKtwjm7sOr80LtY3sHABqSYgR8mLUFGL+2fNqtB6dMHcRWpga
2ebOSkkZ8GFiyrU/bDWvkTzLhAd4NS8t7usFC4UEiXJdlpfZuR/6xspfiIjL
BABZDdLnB5Z5shDjnFsKMt6hcRppGi0Zo0a4LIQ1b0HPiulkuoTPYuy0qQ3j
3sWUZIFpRdHVsPaEJCwi+DCnmseUb61qR0ObriwTVerJTh1KzOna292aaOk1
ln6Be4Zk8iBUFuVW40FjJ/xaEhcbonhCaP+lmXVwpwPP1TaWrVIxYFvnuJh/
oE8KnNsActhWbQ==

`pragma protect end_protected
