// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
KriAg7N0rs261wYcad7jJWuXfzSa8AP4mRiQl33pjKLhAioI3VAIdFnrQEAy
2mvR12a35bjsJxMO+Sn/ODcPqWcRGT8vkg2w75V1UpqzHM28U1aVLKMtmmVu
BkDmEc7k5Kp92oM2WKQbG7TiOGBHxF/xDkSWXhX96tDxjF+GXRt/tRwkm8qm
gi0KHJ9ch2g7UkZNNa3Jr8XCTIGSVIIfzBCD7DuzuMQC+8LO3dr8Ulj38pP8
yRz1a3jd+7Rx3YHb5CtV1DHeYazB87qZVLdToBz4x5n/t/tpyHCszWN2Rw/b
19iD0p37CCOpkbcOugzqIYe2RtZq0FJ6LEOZxnMRHw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
bB+I8Jx5Ez9tTbHF2ldamN2ZGy1JaT8sAY75rSNy1wOgqy4iCK0M1rUtRoKZ
S3BFKCdkOIF7nXRhrRmUBAOyM/2wjagBizWu1hYlo20Tmp5NgomTFVPBfWrM
ObHnYDT9ErOsQzPauFMw8wrpu6jBw5sh2+xe2eCVdR3cxNUXd/ftpyTSoenl
niF1SPxfI/b7R8iHF7bl7UAw0/zCjTYgWld9jQhN/heh7BMTx6d+2nB7/1fO
EJGF+CWMkoboPQcKMZ79PYcqBB0y5J9m6y5dnWm4HgLPz0el98JGEp/HAqTw
yj/up35kI7bMvSFnOi+tYC77wT1GI5dXXgDtWmfF4A==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
flSshUjqNts2/PuXVImYFJ+SQOUoZiqwd0yQjBjCGvErDs745a5f92KKIivz
Ox3w+bJnHmFi5EyM6ySKsI6atqlLHua0Zv9pmb/eW8uOiHhY9LBoDUIsMz/6
7xME4IdN1bv4vaNxe7Goeq28kk61BmnNHSLIZbYlc/uRLxQkn2AT6IOVZg3p
Fp7KvqtDM/kQiV0tbgFmlvB2V8AXm2ZRrTzq0qd7VreFeNVj9jL433Uh15F7
dRF5iTzWnv1xW32bWWriF4UuU3MBrHNF1DxMDjnnFhMsNTpoHdGMkaF5f5uv
mldXpq6oUpD2lMXGqMc+VfVoJ9S5uWR45f0StXtRhQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
qcbTMoETxQ0O+WAsUP6Na9JZd8u+29GYNmfsVgTtbD0f/sujEB72bmuGDCE2
rkjkrc2Lf4gr+Oozd8OQJX+6KyW5HGTIsTezcn2E7ttdVA1QAq/SCvgGaYYo
IJYLYZa7ENWkOR9wKUBPyaREklE7QwZPmlaZVhUN+RM+g14AodQ=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
CPcRsJDjAqc1wuyLYiG9zcatBYFTZnyXfYBpD5Apq/Jsqejg68nmpbrf5YN8
w/pIyLFYb0Q5dktfGL8gJMtMn0Ll5soz2iKMQpg0DQNwX0WLlfMGXk3y280o
pdtcXZyicTPw99bqenzVckuKXiiK5oIUOUzWToty/XA9/Gx3EWoZtKmwHzYy
3yJdKVL5070BcMViwb5kOjaB5Wnv7NPGxZBYHyyWCMQEMCXz+jDJmPVSP6/K
N0gaNuof89hnb2+y6B6kOcOmU/ysn/+JsnGky7HEMNMZCpi4Tg2Tebub1Z42
3s04TH+aPipOyMSx7Bwb3NFL8EuLm4ebONdLRrN/ytKVmDxF1eADkBnH47C0
GLYr48lvXcH2QyUclesoHwEdeSEDNhk7pdKyO7nm5DHks3sz6sRYlJzGa83w
KPcx8iN45TK9yqF8olEQv0wopTuFdKmY4+GhE/3D2Iz8ZjaKiig1U4+0qDzo
eSXqjkAuP9idWYWxsOBjlrMs9KYuGEec


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
aoN18BL+kKRbzUTbMV8tBcc+Qx6nh2+teldSPXAIRLd9Xo1dnzB+zAsZi0H5
aEo9wR1AvQOpmOYp0PP07zV+XYVjsoExJtvMMc01LEOjKJjFXfT7ZIH/G3xd
D73CdMZ2Q7Vo8ZgnAp1we6tUxcO7OPfDpsZY6Js2CTVy8wyL7gc=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
bMpiP62+Mso7EHl/owT+W0RvNNhjnPt/8N6Vrs6xN7FxMp1NGQ2vuhQelbkh
/IdPZnlmeNQW0kq3Ca+PjKyDrHHXAOHsrARnhy8FgiMeKbGs22Dp5cf1fD0/
EN2PgAJ9mtEgcou1bl+Wr1YRoUlQDKWUFuq+0HqrmxZHfz8ZLv4=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 10768)
`pragma protect data_block
tBPs5RrVbAhPQsqJM/hhXIC5C8r0Kq/NkpPvsyAJig0dzYhvv3nq6GOnUjDi
MttM/WardBpFjx8LN+RF4ICUQbT8ERKHkBsuTHeNffjbfYHVBfeKm24Z+7NS
f559PxiaLIM4izPpbjf3SluiCrNcPwEfGq/1dAMmWDYsNQI6vuu0AF6qnmpO
ymkEd0TZkN7vBrpRC6rEdrPaxGTkLkbGyCFwL4x0Q5lS5Uu2BvoJaDBfBOhQ
rJoOPQbGiX8M79Emw/wNBCdiKlVdoTskQ44EB/8Y2+GIVJj6eh0UCgRY+jgE
Gk5av51uJ74Bv1ZC5uEHlsk2FU1Bd2AiM/W9sGa0Yumzc6WCrOmi1+o3TxgV
uGFfirQqSbnDEXPQdtInxOcFGyW+YJtCVCKF8U+Gi5K6vPCmmCEz9WsW6n3h
L7obgYbd5n2Q38vLTq6elM/nmdjjuDSgFIicMTlFy1eQbHiGVTfAJ8PXlEuw
awmfzHTjwuztB7fWibc1KCYmEcFtHoWf+SXcgmqV7ggSBnnHeHu7bdVCEBJz
CJZFjTD/lZAgMACmhT0qwNR/ISTd5geo70rHM3t05ycKXPh3h58Kn4W48fP5
5BCMsX0FrNGXkddi9u1BEEZevVXAA6Yzi4Lwn9wYppznXQRu6XQlY8L+SMKr
h4ImvqaxvfUEM+tfjCgHIcmHpt6qvi2y37BgFCaSEYiyIqQpxXVOwZs9cxmb
QHHSMn6l0Y9WdtGmqVItze9gM7IinWuoQ3h+VNqWgkfF9ASGT2uC5NfoCAz4
rxsU94PBiMQ50nTC/GRQb7BGRtaSOP7p8N1Dp1Z/VxqF/3gDMlfEtWC8Z0zG
IVjF/Z7jw8ngbwLLaIRq8/Q7Idenbyoy3UIb9EKAA32QtoIepTo395RCEnVt
5pqhpBzDRtyZByHblQ/VrATrU3fn4hDE7cgX27m2sQuV90jQvHdfsQXlSsgj
uJASdp8hpCo4T4C83/+xDvAaxafoiqQhbquFsG0fjNyFX/erhpTd2ROB0e75
C3JOhhAdgVvaYj5qITIgKcBY/Sz5lTTYS156RBTvVjm4PjydMu/BtQZc83T0
DfxeDtF1aSHCaOEfQw/WStMuo/nB9VJKhkBmKgIjzrsPFE31GRyUDVBcG2TF
zDYVivkCbdvtnpQNnPL7ngLnr0OAc8+IqNfGfp4RbEx6MALjSt0cp9JcC413
nuF1DrZDaYbT5xVFUo+Co0bmwGGQeJ/9gSRtwmwXDccCf4xgMmE77JYbqG5L
OTvgI2URKcfEozp5V3IVLj1Ze6doRKvXP2uaby4D8UTV0bW5akRa+IV8iSOA
bTvROqbaCap6RZov8J7kiJyZIVGeEFZVW9HQOjGxrGr1bcDOYwEC1uPRjBy5
qjCWXifLcY8xY0PyThaLXqD7N8aEb+R2NAYJR+Q4WY76xcySHpuFF+YQjSvj
ZvE1E/GMAGLLAQIg7fMTkirfRkt4tWbCflscZX6N4km4s84LPlpUwRdoxZmC
9O++E1V8tYnDIZbq6Q6THXtr7iJjEjjyV3ng/VbAPm3WEVvY15+b0h58XnoZ
1HkuIt8c9RSoFWnxozhsOjuT6eKd5lZWpsAHvKPkXEP/TCuLwVn6vTfhbLNq
jToIE8Cwo2OAFbMhylUIDqelUkML32+4lmnDm2qTimfPLVMIrCu/Utt+YNCI
zOiVEQoGu7XGuUxo6aufTmcthEJr4GJeOfgZNDfqqgkJssbge/wkue5eJqJ7
HlOU3T8rcy+KB4DcAOg3nrdSDLsFWqAA4eOAU7dgxDnBb7GhEcxWNjohJzs+
g9UWFHJZOi/iabCCoXnHltQ+aP6F1VAQRVUVzknz3C96Dev/jgJbiHM+KlaS
NTLGPQZ3RJjc9mDybf5iSBUCVuPA9y07l8z3OvddvbGCZoHmmPW/hVSWgFrx
8AGl0KUPHTioTGk/16GMMak7Mwh0f8VkEN4kN0cRAdSTw5Pfr1UmoiAG3E1M
bGe9nz6+tDgevmqT2CkyL2PFZGVFAIEv/thA7h6HiSd2rfPE61lUnLysyzyt
8c83uSv9Fl15TY5NJJMxGw+mMCKV7Gnur3hT8Ci0eqCLmXI99SunFKEl3EcD
0kvOTb8mPORXSIhFnVOK6UctEQNrGLjmz5flIlSNZGkGClRn15Gg3eVTdIqJ
4BgWTR/Qy35JTm/EaerXJdkHplhTy2XRqVV6wOfoHNBsKjAgsvDc//nUbMOQ
/KYj7CVYT098zRdB2ILY/gZ9T3i3FTKJuZBFkHi+Q2oWOWFOz6haMU1gmeRu
1BO+zeVK+2qPwH5mkwuJ0x6BWGHgCXqWu8UXpz2l93rS97DL1aqpaLoZzZVO
YPl9lntd8SkHR/Uoo3OGtBjIQVs41w8DeZDjdx2kLlqnj0VvY+KJz+A5b//s
oS/Eb31SNvUcdWGS467H7Xck6AYKmB7bGGOFt2wSJoXrvJBef2JmfiHOvgkh
9wN9nLx2dCktqQ1PiVFtoKt/l7bq/JhGKJdArTgvJr748U0OWXDJQWFigojY
2YGAECpORwwBhk66eIyf5/egiemZpKzEukKzl/NJdnhuVUBRywGsUqWLvbJy
Es02yu7Gz5nMNR1414Lm4HXf3bVZwm2IVqI1zkbBXZ2SfOIezbWXuguxRU8+
5M6pzGD1qJQGSpCzMnbWsgGbN4ioTmD3uhLDnclcGpP94fJ6PDzslFR0l8Sh
aZspn7zSfXAxfvU64oQx4tWLEIt6bGVRRx4gt+MnoEaHKbDM7MyGT50d2nwu
G/pc+gBt5KB+XzhBTsKlra1BToDB7cp+aDJjF4fD55RTsklu0lnrPLKOqcbG
d3CkjT0EWfZ6hsuK6NDZz2MbubuAY6dWAKrWF0c/TtMMAyoxGjBYnS6GkLDG
hG67fim4gnUS77FppQJWo6TqCTPT1dpiFzjerxo/QW0PYPM8oo5S8k2v0smo
4bedHZnyTNTMbqDIx9pvWGndKJF1X3mu2oDjNaDWm9X7DG2GSbOk8XZmgs1p
VmntOdaF1rZdWnyb8aC3AX4bfd9/7rESmzbxTDa3XyKSvQSh64OwiKd+LUge
t3wES8fQnOYdoytiDkA0b2+sF3K/mzk3yFdzEpl1TbK3WNBIMLmexVuEkxPd
ssZXbRynH8Givqbh85QXqtiqPxz+QfVmqeKnx28093rkXhIbIzdD8hglPmfV
2CAZsA7ADh1k4GTi16+CIqgSjPMhMGNHW0+3YVmbJUcSV9i4RyRGGQDw2yJ8
uaHdTum1Yk6Myks2QUnB+kLhRaorpOYcVfV1A0ujec/BvmoZW3o44GqcwtPg
+QUuoRuhLtRzP1lwuCYRzFo2aX0g3LBFGbjR16DD/ebhss92H9n0uud4eOWg
So0Dds5l77KMOVD4URKbqjVsFiVd4jwekYxaxBH22PveAsdRc13QR7yMV7N7
aOKjKlgureJpmUs4Bamh8cxeB16zhaKixaxKputAjId7yKR5mF59u8RaOz5C
Y5qIz6cslw703xjiYR+RuvYHtqR8i6gsXjqV8qjwPszMONpEyBHZPRy2GKx4
RGzvQSLTBrFQhykO5Wjql2UnBsTQv65fZqzRiievtMaPcYl1EzD+J3P84jVP
BRkmCIip2TLmo1IDrqANBJfm7W6l3hsVrUH8WBCQWFyN1A7r68FwjP/Nu74E
2zaDfwiX9Kuriucdt+wHGzEHFbdjZm+w2c+u9XkdNGupIeKveH9T0WNZIRLz
V64DXmB5p8l6XM+Uun+tzF+fwsV5Myu1Qz76JPpKkIjxSr0u2x1cBlAkTyWY
5G+YzWR6jibwcU4ZVpK9dPO4peS3UghMe/yAEM26FRl69aPYJv6OxkcTn3s4
cWJXxPc2HeaK6NgzWeR0usJuFR6HzndmsDziRmiaWK542wcnHQf++OZ2qLcu
zD83e/dOqgtuSxejJAErjSN2rCPDAbEXCPuTew7juiPibXnq8Hd05kCcIuu/
NBSTbuiH5dkWm0VV91VpCUth2N+gmdHZwoQMy6MMP7xeLkGs9txcdKeMJhBm
H7R8TEQxWzsnIHgnoE31a2vBcLvhJvqS6FjvyCQSgouV4SPQIseVcpeqETG9
bq4BWGCunmgoOU+GpjpOPFzR2m6bVIfX026ECk+Yaw3qTTdrRb6dsN/mm82O
EpkLHBoTejsOJFEQdN6X58DdZMCqpE0KIhu0H2Y2G58yY5LIoPpn5DOSBDtz
bW23aCNo2mQJr3zf3VoVeUl4+2qmDlI4yfQs8SSbTFE+osHuLvyR4i0oMtoc
LhjxdP33JmVx7V0FulNotWhPZZOkzU1IIDpc9cjGM9+9RRFFRMeLRJHxrkwu
tZUZmkBTtXH6vvvN4mXpIazOdvtlALk2xlyWfejBoCg1/MoCdjTUOexOWb+2
yfrELjQPZnVoiYHwtDpUtXfVIapTsLc17ejJNVAaXWe9s98z4UpiRaevJulq
+DWVOuAPH/5ZbUTA+O9Guy//zvZEEO0c0vKyr3qJ00ujmmvTqgDHjR5v2LZ7
6U1hfGxBqeKCYj4ObPvLix06ukkes0jTYkU53vlVexlrdN4cb3lzuQhIyfWx
2DOE4P5GuiCFwKn09MLhDWI1ZCXQfwXriM6GgUBt+Mo6OR/+KVQdUTK4I0jR
zH5L0Es7BHfgIoCA9FAdgUt+v0/HjTTeFJJzOTUVSnIQaVJTOVroAB/SHGX5
UVzz4k232YH78FAHd/sQItfZjBO0mjVfQPnBLKPUUyxuHzcRWBZZPPhRbBv3
OoIJT7A9jJKryo+eVcdysojAIL/XumSCtb1l1dAaOD4Vu0Br1PMqFKeUVnzG
/CM+36yVCaigK8JMzp28a8gGGEI5MApnPbRSoSgMVtqHRcDdutbbRD1Q8kqj
Ofa9SQIbVpL5GqXhpLzDU9ZtQDSDt0klbhS3tQFj/vzxqjTd0iZm2Ta92bxM
hLtHbW5YyCosnoNu9VNy9x80PGXImMzWuROkJciOnIU/5JXjzL+UMvpT+FgU
Now8V8rXissECU+oquz2BPIQgeef/Q7VPOtcju129YbzRur32g8SqJ3NdCdY
upx+aanoRzQFd7RX+fswgFWgfr5S3/RyP+mT8aQPWBxdFJidLbxbzuKf/Zda
G8UYlgKbX38AxApnLwvuUdqPrHbA8BAmSOm3ihnvUK1GGa/fCbVONLcaFQse
5qOuc9whqcON5sfuFlgZ14y5llinxAi+HdW1dFqdfjyCWP9LIhEoHoutJ+Am
Qi4SvH4dZ1zh1kVx1C1lzimqcFyFS1ly/PetTZj/N17+DO99ERXWTTBEJwJn
cFEErPDBn0s6iNevPDDmhfFBe9gRttpW4TNP3IMAkKbM8mrH4XKA0t10DaMr
UGXI4uf3pmfKZqNxO4/jbPRyP/o1Xttaj8AeTUGWSn3nWPpr4CeUqhKMBF9t
xWrRMFxsiZe+ffBsyz8l/xvu4OSd7QnsOQV9IANXTO1BHSffUkNwgDmP+2Sh
QRTE70Kd+5w5n2AaifuJk8QCfXf3Fue43wKXM1BRN6ttRnuEIsSoazn1GyyL
vnS9nsmqXlNLtWkfH9UyExDH5s12ESsCVJyXrF1KJB7re90HKqKAGtImm3CS
8q0/kfX6gkrb04sEHrIxGWxsnf/DgWO9pUAhT7WTpcjlw6GpkEaUbNj4KZo3
AaItO1MZDh/yWuoP42zuMb/tIfs3St+zoUcdtEVbmNEU1cy8EFUb4Ajgv6oR
Os1fRDpU0sfSh/Aq6/8cprUNaAkWaIDqmiKIGJMZiMuvyNIxVMLTJES1vQvD
T/b63FLq/pLBv9SjJfulw7bXc8eIPlK4ELq8S7eUyqaahnQdPYWoIGy2g3+F
i/hHR0IDtEEnoNIuDfRTuZgpD01YtV7wrXwqIuMDeN/hbJww5n3dPIP9hKHH
nQqkNFZ8d17ZnEcjQdEMfJy534BXv6RabloZueHJ6movI3Ep3e+hgPjXDB4D
/IO9BKDiQzobJddn/X8HW8ckzMaAdcYY4blPdxrkagmwIn+b183TrvhHXBlR
psJie7UCGZCBf5h6IBV6DfPkXJ77rpG3QPp0vEuCAXvm/4lEXJClBy/JoRs1
b7UHYTILd+WjDTBSjxZTL/DOiGTnufFujVt8u28WZont9phQ/eZLZxSSzJvh
I+oJfCi4M1oNUE914XwBlxYqFGy9lLYbnkqnP9+oyp0oNW2IZerd+20jtmcf
ufkzTNA0LgqCHfcQL1yBKTTqvwj5yoxG+Mmy0AVQU+0vUfkc9jIieJqadodF
E8+49qm6ORyiyj7aXbmdnXhShN83zBld239HHXFoqgXzGSPJ3F85FOGz+j1K
JurqtnPvCOVvHh1bK/oeGU0STMn6upLblRo1TB9/3ehdwe4hLSKyVdtcskEB
rTEjSe8MBTF6bOnlnl1WroBuzZiNlbL0B8E8AIbB+guncJdPfGyRj0u0Qq4i
7c3l2vLOw0kLrpzupcO8bSYP6PsQpjQXmDQkFftYX1a7vnY4ZY4QcsKm/brw
gDYA/k9Qb8NM8LfIRKRqTTxZcruVz+X/KTZ4+hHEg1hU81Cjs4OT8hqBLyLg
4f6ViyS9HwNHYhlJ5XFimefRjYGmQ/hyOlG0DnnOs/8EINynHa3bKXIcmjKN
+oiWew0nr/YGSXZiikV5Y+nZTr6+Fx+8o5HqzqdBKjTuGokatwjcA5nh4huh
0Fs8oxSnw7WJdhsVUnmmLtJFeiDu3mbLSycYKHPqII8d1WaXQKBC3x7pegZ1
FI8VmoDw/9fnQZX8J9zkqEzZXtkb0QgEZBJgujVACMkEoV6Hvmqht95sRipp
flM75qFDhpE0H0ufL9uaAoqrHj7dJEzmVS+FDVr9Av0KvBYc2+HxA03LCkZ+
7mfTddsu2df5vaaVtBmumGgPXkpIwfsdZKAI7KRyfyX+AwkSCCL20dHpMEXs
NIWVZcn3rR6GgAYcH1cR16qhSpxG03EqiRqEHdOrKYhAWX8G/5OwEmKcSDfT
mBrPj6zT6O2OwLVTO56ciP+XJXl8Wbj2wHLTENDZNtWm735PPmiX+KNtFRui
Uk3BfmFOEzlUqz/0uzkKa7LCoOCP7Wa3mJRpE8QmuQJQsM/JRnu61yT7H1uH
D9z98hQlZ3oLzezYXgH4RuVDkVt8OErXgwdkKql7dg1OEJ3Ti8KttdX2y+3z
52/nlLdh4h6Vbqxqllkry/awfgnOetdNMIj6a32OQyEc2O6Nrxl+CMf/ijF4
T5VqmvAVlT12f1hn1oE43QRVaqH+4MkaC5eBuSsA/7A6Ed2yamYx4auI0fpB
hPsF6yUiXryLSXWs4JjuZBgwXEmusOPP1aWuClZNWeonRp+2NeSwoawIrSsl
HWMHXoU1LgNVXQSiS+IV7WrFV0NBvdEOmFd2M3e/LFM1qYckGx4slEMCi3ig
LyEkW6c0pcWFuopmTjgz084i6yTMiC0XTs/FWtJ11ivB41lMeV0m05FTRG6k
xwFg6f80omSFCEKbhl6c6XmNhDuEXcKxJJoq4orQtc21AUmWq+RpGJhSZrAv
fR4L2732ennfqKlZTkTKJX7muORsklan+cUMvYLAEbZuJzva2rrC38tuoogz
TJeJAIdZY3mQ77oA7bXx1Hq9rHoKcUlcwZ1RZ3i6pG0ckz1z30WMDbLSDy8W
J3Koq7gjO+6rZbIIcCMT8vptOKvq9VIWARzHFODzfp5qV92Q41y4DCBvCmwD
LCA87zjQaiZ3EKM/o6RvPNkdkBmkXWQBDskMUzipePmVkuBkBBzMgoDnG/NN
/62tTErKSxW2GCiSGkv2U437tL7wkgVgmNqtrymXWTTu6GJz9p3xa5/8FrUC
cZb0H0zpC+48K4x5FbxSC4hPfQ/pEwWb6l0akLlXFXlvsP9b+9n0OPGdQFzh
tkXXluHJRqXt9797FAgThzYWF4gCa0c50wDPqHA27HbBjdjVcX8NJyCNJRkc
jrUqi7nzcJUvV4C33eS1ZJmfdrm22c3IYsg0Lvna7aAvACZCTgud+dgOmyCH
Oqaa8EnRg6X5KemKMWZikA5Nc9bR9FcLtbEUD5Y/otUK15lofAVc3LPPB7CY
Q3yEGrysDREmEgF1qsNiCbXZhu0Ii38yUgkpXhgp2I+rDi6HHNozPUd9fVS3
ZRFJifSLlrZ9nj+AQ74NOpfZz7w2Bdi/nBBn+pR8fDh5FceUU95AF6Y4EXTx
4v0GUhAnxLcQxw7uyk13vEtwig7phcQ3KM5W82MKra8nN5fanAOretucFW35
Ur1YRzUfLgNHfnPPnblkG9/9D0fEoanqeuMLyd233jkRWwOFJ447tg6nNKlr
6D3qSInZRmgngAEyYyjXQWdXWlhfOYrnL3JZmi8pqoESmT7zt1mi+o2wdvED
QfubIWrQzL1rD0lxC5LzABCqXqyUZ16U31QjmydqMGQZuF09k8azzMFprHbn
7njg1IJGijg52k2RSOyT5/9Za1Bz4C6eTk/Tdmqk1o8VR6tv9O+lsE3l+Eum
aZrRge4zuI0SfDch7P9/UWlVhTH6L2x5xlZkrZnjW1xqeBi0s+nVMlv1L0y4
qUduVaEqqgjSXHJtoVulLBiVOTLDwW2jT2RKr5VgSi+YFn/2s2fhnnm+hG1h
kPxJUSmak8efmVWKs9du9ayyyPKislBT+rhGsu/jeTuUybTLeveeEy9WxD9y
DkEDZlb8JSBW3lZxcZTrEdQ+PuRHSOEJDANS/IyqCp4L/yw9uL/awkxkxyno
09qcDCmtfgIYW5c7R8vfTZRi3K58foFuPegHLG6vPhhLbGIV6pJzkqqN8GEi
T6NNlZlWdrvOhrN8Nxl3RmyOSDKc6rxUAkcHV2t7Yh7VPrQDyXQLcoA0Vyn4
APLM9rH1jNaJHY0mouaiJ+DGUGsL2HkbQpyTUrH2ZIPHiGIj2RVAqnSnEXJc
yLx3Yjdp9Awg95IxuDCnm3JKK8NXZw8odLTWl2Ea1QnDSpvOtseQL8UQ173l
8cS8XqSGx8VQWqyh3EQ7AvX2Dn52psuzOeQdU4jpaLnq5UNqkihPWrZL2pHb
4SEqso6BiPy8MwPcnrCDGqPuWM/FsblRpbJK+u9eEuCudN9YtvDFISMBu30P
svnzKdreASypSpdcklPDU4UgN11X9sdB4sedsYN0C2fxmZWj1FsAZFxSttta
4XP3m8P1Za3WxwauZBppEwF7QLMTxGbayoFVWoS8N2Ai+a3BHOoeTP2T41ft
wklA9X8BbnY79soMU37LV/y2AZJ9g7UZ9EFU+oF1dzR65JwJCnMTdYWWAMdg
HCPILtn5VRmjRC3B8g/Tc0J4jBVfwqGjX+EMtkRdeJkHXhn6AD2d1ZBMwzou
OzIV4IlhFkJFciRQG/0EbbNxS3no1V3HifdthntT2gDA9dCnEasgwc0NmOjI
hmqztOVzOKuu1frKaaaDq0mdqpjzhpbfVQQMTAEmIUnwpGXAGsM+MBTEnzHJ
5SpOGAbWHA4xW7lWF7JN4rAhmWSl1zNkFtyx+JvDfDrQb8T1JOmsVkSZtu6F
B3ljqRCdS5QBiBDLMIMo1s35SOFx0clcTuhfq4HUOY3vpd+FihNMwzhhPDuH
rB8QyNWkhwRt+lgPcfYGDd9jtLbLY+SWBqTDwrolnW4i9KYXBpF5kvSgptph
IVb06knig2PSSNabeTJc8dmnDRODAvzsLFPNn4w0ggUx9tMTRyMHA4Fb3u3Q
CWMjzQcMXeT6frSAkybrZTN6nbtq6bU6XJwzjQHE9Lm20gNglwR68tHx2qnN
zVV8Eq9XndmZibJ3NIW2gddr+pXWSULAgV/AWdDm6JxqYDAyiOS04SnCMdVw
rLSwVPPRG6L8AGKE7qtmXObH7XN/hOmzYnG828tAxvZhuEZmWIvJ1PiPy5Ui
VOzIOcn9+m2KedglkE9fnRDsgbG00MPnKfTuZLn+LsfPvdVjo3pgNduAONvd
OZDQDNTEvAcvWqIy8HCLAuptk1YHdQ2lzchycvXekp9vLhJhvWdDchxoCXDt
Tv7YDvZnAiYVEfRfn0aHNZn/zd0VGRMdHJL1GJFNFZezq0D2Bq6hlNB7inn+
lCQmvjJCO5YRB6AeN9D1v0QgdQSmR6X9IRnHk7L899SA4GqYD7AsTaKsYU0c
7IhuXhyGulzxsho9KHFdSwhWkyq1f/Au3l0dNL3RP4WbeK7y1N4pJTMO0DNT
ydpNHWQ11aKkGalnQfGxTdRQtKCHram4+jz7IE+FzmQwOqUZCVrXyU68S5+V
yoPn6fvaysIJeWOyeFRkjr3RYdZlxdoImvGawPvDeWm4rgBvNNbYvc9j37pV
mbTK6Aoam20JPSFJDzo1T6Wkzbu+x4fBz0cVWbNtiFnVW2RiIQEgQcs4LCYG
WREAqHWLqTciZxqPUFGxusQVd4o5p+dNRbp/lFzP9T0oqXrnrNkQBfZENp+l
1sRsAGVS2JDLGPFIplhmwi1rcrRlFjFWMVqFsrmd30mjFddsNP+RLTigVXwo
eawwNYTYwmIu7Va6GxB3U7+oJioRGQbhx0DdOKis3w4p5XuUmJAFuV+eCjfT
VT4yJTNUgDSZ2bqHjiz3lGD/C/l9LLvKMK3E2P2cmOzJe7/VwiOx02quwzpK
l2UdOT5b8PurFqxTg2jDUAhG3S/XXFiMVOhZUC6CD/Cb6dv25Tu6xQZw5MGl
H4XzVpNpCU8R2H4xnv/gmSPLwXgVZUHzapIKx9nrYBKRjuns133vnnKXmT9a
eiRNi9ty9p52ziq31t03wi3mb8UpyNN4UNqktoeaGCWp/yfqafyMRumZB86g
8JQ37T1AwnaMwuu3FK6f1ldlMpT9cC6Xi39DxLIrU8++eXjIvWOR39Velzp2
eS606KdY3thSZmFOCpW8xzPnEXGBqT4aGnjOmev6RjF6tLNeXWz1grwHBgct
h4OrwC4DhlIf8r1xagkFbYnjU8tWBbYCHXoDXo1ElDK7XQpSsJ9JWWdlj6al
EiECFZt+9E3LON8dXEblpubHC+d88vJHQZ+wBp0C+jFhvRyHxbDK5EwAmyBj
ulcwnzGH2uckyHDEO6U2pVHnbcpOfeHp1aoXYAEH2vCWRPhzxgtLHtIHTSB/
rh3XmCg4L7XN/gPq8sNUc0uet7NM4ygp4+S5+rJwPsCqbENhxKdcCreNaxHx
jcDzjMPyjZXLLxFNs0LQ30ILFVRyEQzJdKeYP+sepH0qSRwf285UNBj70s5w
7FujMA7H8VvO8xnlPwvseOSGLghigkQPT+Y+XiOrUlblz4CMw4IdubUcHuo4
1HOS/1aOz2/Xsh3MKohYyY46HtkmbQ6sAEktRnzA8v6Zb7U1dzVh7+ptjh+q
xq0TV7E5kGDlQsryUPMUiXbyiPvtIjOSoY5yrtyHQD9HALBpqt36FfSX+8am
TCWsYNGhiSmzmlZBr/8VtwHrCOQt44mzhV3cE8kSGant//M1zcRKIrUBVpxm
lCqDxYhk1A4W/Q89SIu6SEu5OYUitRD1NurCbU0jq0Xp+EISpqflnOvA5KvJ
GFhAM5T5tUn5avhCxRq0vIBqv2Xw8kMKlIVNb781pPnYF6docmNo580/CuWc
Dh2mqYQVDBCVR7timEc5uRHie16Upq2ko9xzGjPE91uYbjfJeCF/VM7ZSTY/
+wVl2q6svotH3rKre8czHRkHV68focF2qahowJnT3td03wIJhFARY5X2/tkK
XTBPHuaR+NXBJSNEYAUjxw448v37ByLt37gnb64+1scN+YaVmLL6+EUdALpd
2u9tTW1afpbSzyYVyYj7G+4d6dC3OLW8+OC8KllJHSMoQ10//ia4jAkaH54V
w4zzrQWd6dfZTrcvLkIHdM/CSBCHq2Iwl24jM1bVIVgKI2cngdoMddShNvXF
c16ma56Qzp64+3ZxL24+KjGclCObNJrSZNsAI0ZvCxXuMYK0R1GIxNk3k2Op
OD292s21m2kbGDaR+nlO4zC4iEC6h3Rsr8UF2SoP0WrReyKyZgQ7nVkLiN60
YBDBJnuQKSVKs4rmUDbOVx5Vrr5VmHUqtcGOW6UI1UkjOQdCMEvxLJxVQw59
VhV24nUyRuAnkmcC2Fh+rOx6Lx29Koo6LklJTJRWTkWecTsgMbgXc36safC4
aRxOIqrllNzHMt+UjVEOvSc2Ykno8qP7mM1khDWvpKtJLazEe6/F5WGbom1J
BphFIg5UjnGFcbmOq1Mo62EIBDvX2FT5gf2jTjyv4xEWgJk4hiAL2dZX9q8d
SXvfB32o4DdqS8/qXlQGRa7HsG79pSkZvqSoLAXUHQ/wUM69QanmSxylZI7D
d7JwWtQMHM034aUr8uOWl9guOMKv0Ir2ggozlYlcqSrcQo9fm4VgqnoF2ULt
uEgNqKCy5bIMPpZh6stBKig9pTmAR+cawfaiFKUWS71VjDX53DImrlco3Y/K
okylnuXOWwO1ZYbfqTHtGGOH2e+jaQalxgHe6l7AxWKpz8eJBK28bU/5EHLj
G8wvkXPqKdHSKT6uLUVMyA0c/QnYQznEfGXu9xDR2TkrSn6BgY8HeSwUs+/H
cKNlWeww3WcTowKXArhUT4D5var1+p6KQBo+hAFkItu6tdEedKSzMyLvXF7y
Evzyv3jkX+GhOqGQ/1vteztZkTzKDsnBWgtNJ8TlRHZuJ2wz2SxuAszeLGci
yuxV21kb/7BlF8q+GSE2YATqOMf19LTDcZVCQBsoQV8ve2pSz6xujYzQ+qb2
DxGViZp3KXuu9vWv20/aNMxfw9KYaTu29KJCNNyvpAKN/NkqRqfoZdiiRsXM
C1iAmZDyCgkYuomq+O6C9VgnPVvvNNLk69zh/F4vGO6RCgtprSB0QZdlGcNC
Cg2P5xZBJpC+bhNWg64sWLCfiwisOAfZaULpkYYBIN4Kl8BqotygJ1uWYEyP
BKH682JzjafiWsAywfw9MD3EOFZGRSxqKFbly3yl/1CTCrNSr4WVkukVM8oE
SL2YnEtME6TW4Bu3v7/zfy5V0iqko4uz/xF4cx6ItQlbp1I9iD8OQLTdde25
gqaawWOPMTLnJUj4swpdZL1ivJm9zH4yvjXCp59IZXIhsPZOl21LxQFCH+Ot
l7vQboYKZmwz9CX1eiFSoCsXIqu8asVPDhyy2EVJcGWqtNoRgP6b79r4HrIL
PBJY15xlkJVAfHd95lkgGRmNq80fGi1VUMoZjpOmUlHg61j2q+G0alWoSlb9
EiNGv/EsVDXMq58d+6jkUo3XuM+dc07YxexdcYtiHsHSAF1lr8Ssi6Bx8v61
SfH2NRX6nksvdxPHlIiC4fZSB7t/LRA2okV6IkzJlK6o9ePKkOVAJOY7dMMk
WI1Bzzc/zEEGExTZItbvN5NSezzZBBAkC8setcjk8y8Tj+ghp+btnaXuQKjp
jmrNAu7CqZTMK+rSAGSJe1WMSjWSPr90pbnlfWYsL40p/eK4Ut+ljYmVr43X
EECJwPyURW602k1TxclryrDbMKPlAY6bF1DhKC4wy7sR5Mf7EC+u7pnyr3ok
QuvmcNc53ure092NuQy1EiTGg7Zw16PmQ87/4ZYzLcPUjmFkHuskGCi494zc
OEAxnScUme41+ZLoYmSe26hy71AmdmjDSZqOdgDVUHG6KjDNJOviv+xZTQpT
rSpbXo4ieEClsvxm3fZhX+7k4kv4rx3KJxM8M3an4z5gx8MoudB+IJdowS01
LCCr9saKqi4myFxWu3Or7eRpneaV/LNMUlLa/6wtsZ6QA5cNbvA3Ai1WabD2
JrEB+StzEDiLu7PnOISCMr+lIygkCGayPR8bfFHfYRlqUXqMzOu+xmzFRcvt
1zsushDtIvpghjCg5mIkAE0jcXmQwmYlpFx/pNUg6juYRXmoZE9Y1sETnEGJ
P9jIhsIhOccWPTj/tCQLoN7wunE6Kwu1JRBwpgCaHsWSycjpGLwFAEa2c1c2
gGb1cHDKPcsZGt8QRT1jVkMy6TwfYFxWuSTW9V7OEZqx2ESbiBa5mvXjUpOG
9bc46OXJ5s0to1YxuWZ9lOXTtICiFc+Ka/rE4tYttwqY6bzw+WoIvgtd2RtY
CQbv3tUtZjmeefl3bWYja/N/PlCM7XjCwJgEOFHrSaGFdMHX41t+NMSY1UD+
N+9kPoqeif3S4ycGWC436uz6nu6v6/Dl94dGwwDkjuhWX6SHI64fIstB+zdP
pM/FaWZxMYbypopHpCLy5h7OXvMSax9fVIP2nuYKz1CGfVjvo3oS8jghTint
cgaN1IoRyPkZdV0id7kQIlDRgOqxUsDHob8wwbesKJ/2ML4vhEFLQhASsayG
zHa+N+VcPeEs3Y0gsey9k+PzOR2uehsJPwfshJAjLTg4NQC3CmJW4LMhO7m1
C163EQp3t7+IqB3hwArw6gTslp6I6IlPtGUgcWqxEpr05obPDHdg5wbT34hb
iJwQv/in/3A9VcjaEg==

`pragma protect end_protected
