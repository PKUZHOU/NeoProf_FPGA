`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
X5H88AfRnIIElsVI0/fPEu9agDCDaKtO2zAWR71GgRggndPcld2LyzO/1eBYhZwx
dJHZ7rpox3V0S3X5tkd6KO66giN0YFd1ew78QvonZqDtedQkw6LkcJoeUe5e9L2o
M/cdNt7qZYMfTnI862YzdH720guOhh9tl3AGiDartGY=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 9616), data_block
Us0LEdrYgCjYvWJS9KMCGkJguzvrcgo+ik0Z+NqSbARwqolC1uym3AZC/txWB9M0
qA/x45sNaPBaaNC5EwLD8GhLCAVJZdmN12CmgB0dMQW/BVvp0g7RJJL9QJ9hA3mT
5N++R4Ui3VCzPsu+gh5bQlnwpYf/6pWLZBG14JZta0pcdRpJxNyLBmjCke6ZoAig
T0Rj4G/H7Ghw5V+4YIIffz4vUVKqv+qcvyY5/d9Ydate//1LS8isJWMXJc2iPiD3
8DUnQj+aTpwt/OFgMuNF/T0mPDIh6Z8+Olq/1XKc619s8HSNRidq62p4cnwsk0if
6BVPNj+Bskw976zJv55RdC4RfMK6mNwotHIAH+jpErnpuRotU2zyOnJJopTzN2u4
ZtiXt2zr7ovJY59VT4eE/J/1fUQACJ2bYo7/o3lvyXgvszkEWQQoDitxX2UoWQyG
u2veua5h7/Om3DiQD/az2ZDqMViplxuLGs+tIJDRcM1Cix+9uwLuV844h1xV8F6J
7QX1QiEo/Af81E2ZmlMol1dQvoNixbQZdZg1nutF53Xj4DA45AuvK1F5320qnGSk
SyqAQ4EQWxbUqh0jLdoBm9pjaCE8lJT5KJzVRrL5rgWWB9tgK44EOha1q0m4Bbb4
CK0WDf2/S3gVpFaXwss2vCc3Fx4fwxhTNWYR8YZxzaoTB5e2vA4xUQoLijwdpw8C
gfKwfnoz2K/tj40pLX79Oet/AHzUOZQyyGpks9sxUd+gjo45U53n4OeQ0amnRNCH
nC/7E19l3C1RBEcVz28CvJ1A+qfJeUtfOHZXYUH21UrH3RWua/FgpR2jcwoEdpRX
k1ASlop9foHiYYA8kRIlE1/73QkuzfGFEn0OINZV5Ptatk8x6PD/ktx0nZ6istUd
oqPhFvI0OPiJP/LJxQkiyZUEAfs+aZfMwb/kIaCsCU1S7pgUicGKQhdbpAYGUW/m
BFzck1tfOdZu52ribFTphc5D6U17Zf/w2bA64Ul3YSiqpnIIwwMoeibtZq1A6OvU
nRacHu08zXvOPo7RzIYRbsPG//cqQBbqQmB8MNjZx8S9DLnL17wBC9ZLFNC2k08y
fTTFmrq5Qj1vZJh0Ul1M5bg9gSJ+K21RSWg4xhUM7ZSkc52XeFvHi+xpk40lRCXG
3V0/TQ3n5RtAGmPlxjOFULca30Za7Kuwro3nxZcTM5eNX0Z4SmAvkf+J6YvBKS1Z
p5+9FWfiCFRNdRLfi+aYh+f/bjxmXnwscCLQ89FOA9QvP2GPqXbL4ejpMWrlcu+K
NCwWS94WsuupU/XVY/vs+fUEkNtFakxQ544BIuGcQyIDpo0fqovoEjKPLXYM8FI3
WaqZFntu1yUzG9SaXlB+XxJEWwCl2oOsz4XngTTY3ENN4smw4YG9zqD6rVO/FrMs
07ZB+iF32myRrFUuamgU9Pfx7y0pkFPHdOM2y1RdUyxVKUOMbCtZTv30NOAnFErh
3aBmM6NLdLmBw45voDsHBQ/k6IU3ICIcJEXOIYKK+4y5aTgkxvqyLI9zihEMZD3w
fHIp9mHlQN1YKTIptyFNiqKGxCLI0yrzFd+bGNrQM0LgwoMNxWZShBmpw8/ALdcg
7I1rupQa6UZYLnlSvmYr4BjllffGlWZOeX/585VlaQuy22YNot0hIrBzSdxephXP
w/uAYRIXGFWMe4OrC2hBqHAmxhBCOB6oi7gxAC7BkdGk6wj1Df3sprkrVVq0pDzo
12yeG+ssaHos4u5Z53sdxiVL/xDa+CjS6SfalEcHd5IcMOcq8j9P7vbmxSsU3irX
sZsBVUwSsmDStexJqAPypRjFmWeCV0UAWFgCEC+T7r7/fU002/xqUalegp9UQVCB
+NMaXnE7KOB/4kePWZZWfVijwm1gstYS5j4L6Ev3EzLolLu3Hi1Hm46tSTCrw+Wr
KNdlRSW+Lg9BsE7BxLOYfzpPw+9RgCp6+skrHVapfGIbFdqzo7mNYFy3EpXXz+zI
ypWWQIiF6WSs4dUq/UEIio7J+oS3vw64zhScCKm7Cls9BbNoJqCHAhOAx9aq0ikE
3qnHnGNvOK8rb9Pazjsqnl9yR35kjws+Yq6X0un3yHGW5mD091b4nEIt//Selnoz
DZyaKJxbuT3GGyh0IrFHizXqaPE1VqniFgchw0oXe6PKdGGFyc3wzUYTcbdD/H+2
ICB3SOK4O9yN39tj2EomxR6tNERGXOyAZ/X8OWDgyMMaVydSA2c1KIEaKfwws1BL
WSSkN8U5G3F0e9RQDsqZFzqa79JEV97xp2BAVVG+jtLO1ncXYA+TA88CDot4/f3u
fdkbEeALSEocQ6JmsrUiN6hF2U/2Bdq/vegWzEUFgmBpST5JRW+muq/xkChizy+4
/0e9bID7jbnPg15IrC4A3mhjDEBLD6n2r31qw6hjPaN3YlORWUa/WDukoLDKPYtl
X0982ROMI+LTErkzTeCGZY5hWzcgSiNaRQQQ1h4hhmp1rVJ/Ynh26+EoDxNMpnar
6pCFSjxD0gge2NK9iqrD0VVQT69DOlmoXTJqsORiOcf+QWajlOL3Uxd6u9nD3f8b
/uZHgD9YKfL+063jfGabSrHe/XSlMnGRlv4P6l3JrXyDVJyRGyJm5n0Mrnz2ifag
0Bws/t5CQLxapqr1sxZGemqKNalINZRql7X5f6Mh/WocTuUrV9oXRf0qx8NhNiot
9hbluW/+6WIuh0T5TmM5d2ShWkQUYK/Ury/CJIPi9qjRmW1UojjleGgINhTN0lVh
v/+MFuYymA42xPtGEsv8P0j/FRzz/dO26DSPlu/fMXaV2QKE6Uu2EbFOovOStPqC
9kvxjCX0/xbqWDeJDhOl7Y8upeW7cqc7+SPGy9Buon9kZ+Z5w3dEOfWDik4Ot0QN
TuPsRVH8Jh9Z/mm94wYdX7HDXHn7k6gvqBLD2cjpDOEK7t4gBdKOUMSMCnH217YA
9hbPb6Glzu5+TLYeRGNP+Q04V+dRO/YcSWpBO0IAdhz3tVuZ0/8jtjlYLDzYJvL2
UHDamDAcaPlZzyBO+/NXU6nnmMjKvJNLDXmsYHyPDCwTbcbWDuNohkOJeWWcULje
x6NjhSpZ2WxGxQtA3yjLLXDIcH6g6CRVmYZdxBs5eV8PP1j/ttQIr8FW5VpA2WJq
g0Hw7+u5wTrLKa3grEG+q45yMKIytorAYKQrNpwerAncXERo1viFNxU775s/F2/C
1FXW4xpU2buJR3MHkeLAjJytQQo1+na1dZQQm8AblU3TwPi3MFacBS0fA18rrFeF
LFFjEUiTxwtssJQ2TkhY0WEF3q+OtM36qwaiB8eSN+07aj8/5WUpsQfH/ChZQC4z
VOJa9r64Dayzq8tw3CyeetwXRg/OtItwY3LeQKLR6Z68E65v8KGQJMT3iu3t+7zw
ASF2hvlJTu9d5JWeSWLRl/QHxDPK0DyyFvawSaRKUZ0HAThpt/rx7WI+UXGd0CA8
8+W8ArAVcywGDND+7AcPtUsZUjU8ZLTgx+3AVqw+6R+gurd3Nx4QD0HARDcteDKH
qKozNm0bwZYIbRLrSMbcrEwrGGu+n/ahxsbm+5Ue1Nn1juY9ULT+HIj3HUCFgkFx
d3H6KiZU5BDoFIdPz+8pHSNACzlWzEexEmfJVb9FYg1SB1zB2W2eYnTpAKxGZb01
MzTDWogK02UzWQpvS+qFxM16TbM26xQW8mJQH2qVVYtlL5Ael8sNpfhmvGuq/oSE
MLIhWSpN2KdTQ+9MgX4GD95sOkHpxbIsFviKEUIf0aycMuIveomypLggEHNr4mn8
lLbzfGQ8PYQXdqYxnCizTpno4rZ3Itel9EObBz7AUQOXjNf/UTzqByRVAeWNYVYS
YAQtv5IC/IPFM9RqtUGmMcPb7Ck1CjFLxoXhGnnLchRnLLHvd65vNH03Lgcz0n3V
OhTatX0SJ93lftKUHAEUEpzx3fBdK5SpSsXjtovYi/B6vLh0joJzEkeuriJlrJd1
xcg9/2zTDDvcb0ofC1hIdbj9v5PT/fgIlQGIO5VDpQdPOoL8IU0W6WHd6mfBOfe/
PHLlqeXuo8TqEcyjqsGYsDbS7P5EFOYwukb7IqKByvcP9wVd8kxWZxNTPiA6z2FL
PFTl5Bbo2WNsSmHzB/lsrpw3x1a2mNJBdVGj8kwNlX8X6gJbQl17ZKuB1Rk8wtKm
NvOAwnkXmuW5E2JU+oQu8Lwozorz2JWtjkuh0aAvnqUOTt9tSK2Zrnsu12GyniLi
8pUPSBcM8qgUWJXjWgxdkAmj2nbGr+uQBnGPt2Y+zTnELH4cGvPYuVzomKBdMZYQ
uFFLcSV+k/YMP7xZTeM3cQKJGNT4WSkQ899MiJANP8cT8cVL0IYodWy3U2tEmoUY
+aCwXHUeeZuZr79llfOUW3xa6FDCyyh4nANGeuKdNlMR9dGY7LABoG1IwaP2yZp3
aG7g6fpC3aeViWF0sQ9JghOBug7l0GmwFvPIhcXy28ivvJ9f6d5MHVqCpfZLLHd4
WutPBV+1mHp/I2x0WSCq6dV28fe7/O1CbljcrhAN017x9h/LJUgyRP6J/UHSQqgY
HqhLOvk+eYvleRz27qF6LPpGDqHH+5KFuUm2xNqBBhA8XgnEU21DkJTu8tsppUsS
tBfKXLWSu+32/aXeza5KwZq4LZ1XaNsKJ7c6FUlXeyDOVJnhLEP9Sr9zCzgLIiZM
Bl77Vxy4yZxP3/U6xXBK/OimG+T1aW9MJdd4VY+UpaKTDY12fpTPcdavStn7EH0y
y/JwBN2SxoHFSsuggOPC8+mL/c6dFIbNCjAk9Kuv+swq6JiFdlsW2qmBKcEKls0V
EHEadciDsa5X4tQ4LEYekcdv80TYLnjsGcmFzkgvyKkpgyXIlEXHMHzPclmy19bC
qmUHtqJwQkqE7YLhHAao6joqMndA31K3UrOjzJjRw7kbreEq2YHj5WsIhC7ZCafZ
m7vJU1M12Deua9VI/aHVwcOtixKnyCxslEfrHIXBI6UTjgRiYjBzbaOlC/V81TxA
BWQXMcqk7LOMHjPmJxwL8Y/HdMZ19RoDdOPXK3KayBhHOYBAhDTo4tRYfw9fAwNh
8jbGOli9JQc5iny9VRiP+VPQsuWOUxw/eamPCBLsHfwwP3vKq+B+YsRLKcf9Quwr
BHfudrh0yrO7oj+TQjiO2Z0xZekn3OUPW4j/ppA/X7YdeLWMZn94eQtwGny3kEWL
cDvYaSdvi9AP/GC1qdq5ShQTvBYcnoJfbnjUoAoohrWue3FNFAokJ9wNUHBPTJV2
Lr/46z2GFSJMrwyRaQN/GrI8MCRK+Ml+KlYisyHzur9YWdJjGH0gql1DQd4Eg8tj
RclNJM8FZGuwL8VbAHvdA6Xogf3KbmVXnU9qFPueZ53LnnuL9zlXu67poBZZjDOn
cwvrAAOa50iYS14ygjKaCks0SkxX8Km/DkkkeOOCkh19YsdWmTdI8pdnSgrukwrn
BxvkhHt89AcYhlN6yXsbahchv+kb/nO2ftjlrESGasE9vo+mW2kyPC7US8siU34x
wejvuZ1k6gr8v3iTkHUimud6OypSl/zWyD0aEZuh5loJH0Q8q7ZDyjZFvJ4Hs+Ej
UXIPrAunI0JEYnR6nGB6HVTdGqf+9KDkRhj1RUi6rKgP+7f64OkCXDBALBeuoz2k
ijvBCVsl1N56xcwzWsCHXAgh5L+Al7gpTWoGsXBLAJL97e2cSy1yiB3uNVUB7R+P
RgB4oq0MJ9ggra5EJ485sfqaybVE+ZORj5vwgWxlhUgUHx5b1nagEZ65DosA9lRc
jyWPWVI5KzaMIJx7VWUXO/HIujbDhnHfk8VVl+R0kVhrMSh+pQgUxEuXcifvd9Bb
UFJcXfRnI6veLvLxBUZsOOLWkOu6yoTE3cc8caz00tWr/A1AzMHOnNOmgGqA8OE3
4uIjKuknPNnQrX7BqWgCrdhxoZ/kCLbKdf8IPQlf36xmvPqvJiKLmUl+QX/EjYri
ztocEpVRlVzrdYyzclMeBV9loj2Ghv8fZI8VEf0sCVgah+ldmMFtY7Oi39X1bMV5
7eEdq2fCzxPK5+dIlZyqm69cdUjURhnpgKplXaSDNdhpSYak6jKsUaFGen8PMJq6
OldQyJyjrAFGA2tDwkFnqUcecfpeGYAsm27tWQT7buhiVn+Dbep6eShEwF9Rzt9P
EUKEyzWW24L0aVcB8BNmU0zbH1zVYfutLNUC/eMT1jrz27RMo2Zy93dwbMqMWZCc
7uD7xkmWvwO9Rgut/qlElr+XlSC/f4wp7VjM4jjfSp63JbLEgqOoHHXDbH1Li43q
NIPEgJn5nL8W9q2lAFy63/TNv1R5dq75oa4itdN/hyOIK8HUl4GgNhVR4YxxqDCl
4PwG1o6REJBVMcdeiDRPDSuNsxW2LBaXz6SB46kGQoNJ6h2wfn8078MprFRszVKI
33bgDWhSetCsjyyiZ4F8jTM4HT8o+TggOaQIpQWw4yAcrdj/OXaIF7PJ7ejFD37o
4qwO9TuaokbnTEJvozWIUvQk5h6K6zbuD6f7dnRuGwa/OlH4h9kQUb5IM7txkX7H
GjlQWTqxWsA8jm2gmksiVkyUA9unTBqzgRObSkCDQ1z4BF6uFx5g0ynkqoFDztuY
DhSB1IYnJoUd4G86i1aOG5gPZTPJO638mHtnZ2+yMjhMFnkH66gZCTFb0qgffiti
/SC5FopPzg5Ee88G/2yZxN4IH2jTWIGlsCaUvzgg6SZumyFckSgx36qPT+OEQZ+K
f5NuAvbefBDEl0BptocmNTfxpf0/LPwPL86u82wpoonwODx2LvNJXSxbVT/akA4u
iBm9knvawgf/iW4yWK1PnapSAwF8ucLql/vQvt9vYup2VDf0dhhnvQS9gvDVaedu
9Zg5rhpY7bOYQDBHLzvM11cqknssQxX+jBZGVUeNFdp3gIJINEChG9DR3y3mgJ21
ZQkJTOnwEOmqrc5q2c2Xk8RPdPHvQJ+uhQy2hREE418nHHkIGP6n5IglXDnGcnkl
8P57L7hu6SanfmGsD6G2sZbyY+5L+nMzONEKFZk6scP0nBZ3p8ooRW3q6Qg+xXI1
lzExFA65h/hsbuQyB2m20LwcLje/g2kR3Vnu839Qkb6Lszs9zk1QF7uO5dqvH/Y5
W3m55tOF712CHWI/XyOrFkxKfRn5qMiVrazVDibYSiWcFnkLZWJ63N2dOwbZxPEU
aTdWadpMRIcXigKBQKUCf2SXkihtLuo/o9745zPvryXPNqON17TWvdFyFgZtk16V
94QEFLYfzKQWaAWpi3JNb3Q+68AMar7UGzNS2rUzBMiz36TcYWdQvSMki1k3MbCD
Fw2x8yjtWDDT0Yb4mkspeqm7k7wmksPC74Gqn35oj0H3MdkNJXbdiFp+jSOpHSFs
Gmav8qn3/P3e4xLhj8d6r8grGAaEXTWI/YwEJXT+z8xi8f1Ps7udYpPODr85A2cw
GQse/C8aL5dJ+UgFQgZecNcaR33KRNGecwGLoE05ZmIohWmR4WDwRPlccLA7i9aO
peIBPlDUMV61frYtG1Xmxj9kO84i09Dpb/2b8rXnxUGoUJv4ZAs1NlfK2QzjAMoM
hrpJQ9z0iTAX+XEbxefYZjz5XMZnMNTev8OuqRKXa1NN/MsQU1GmNRoHr9zvdU2o
706lBSf5tDTpY6RB3+SFnbfNIdTdn/DoVPPjAL/elKHey7Uehi530x6mC/5NGGqd
4gw5smvNmCRVRddpJQGUXZcG9+pehiQHdlf3OmFs38N3g5W8Po3Z15RdrcaLrJ7L
E9X6tewBcjSMJ2tq9ccZwbuOSW8d/x4tbdR8uKNE7+iuXOWGdoTTnQe8NAHGp2en
EVJ6o2r6L1byLJaDHmmN2yZcbKNt9ybDOynKBoe3r434pTh1Wn9y9665iV+pU1wI
xkCDXmFYjdwCfOndsUhQTjgTv07KIK5gjx3b5afPd4tBAKmfBX5lTfcekynvTnBi
l4P8SP/rhIG/tbtwGOuFtZ3CH/E9MAxmGT5cOBidY6pBUsOZT5uSanGegjVLau17
Fh1rv64prkrw+A6Nu/uHppqEO2Va4EZmJGPytm0vH3jJc1zR/8QQ4AhCGPVYhp88
s+XzDZtwwOJNhtLs6QXICkiV9lBjOvCj9RklIAGRV7WkALmmpMdilLQXO7N2L18w
9J8wb4FBGhC4jT8ODTQVSi5TQJrXHrrLdCEyU7I0Me2u9e+KPQSOdjR7qrkjb1/U
Y1b90Euk0t/i3wJBmMOJ7fG/d9mA+bhu9unk0oGichYWh3SFDSTl49OBOb13zuY4
a1cQoTZ8sAwVrcHfo3fPr3PS8hkDqaook4C8jMXFbvRT/lC289PvDhHRYHoMP1De
MxsI59B/oBcODrb+1G6iArI6jeSGZdFtURiC2a0YQkNb6/mwIM3H9YbqOcbXJ2S/
o79+ZQdpy0bomCnK7TYEBmLbcu2ZxtQJ+uzCpkpiwhdF1XJtKlg3/2dRdycYXjd/
lXlWU6J2/yg4y7uqhNPnmuXyb5rCapAs5WpzSS6PTpEAUbBoRzfbL0qYkgkCXOwz
ohr2uLFCGgW10kdppBh71EDQfR03fK2M672T6Ysd3WkCDa3RgSpeoiQQg2zlx0Z1
Nlg6Su7e0HS6nXTU2fyeRIYMaUaKwk+VdmOOvg1x6iUNYovcdAfbwXvZZyDF9Kgx
TOOJvgYCC4oVSCzlF/8wEwM2aLQASpdjvKEpPj+337psOTwS2/WiFHPS7sug2pCv
9Eceg3bjj0E92rsA3AYDGwOTO0hdDyusB+w25lKdcbxd59KN76bdQ9sMAxn1pQDa
P5+cDZYhKqiD7JaW9MP+W1fHSjsvh7nb3DncbNxNjOOfS1ePG6bFOm6IQAWh+rem
aNggtnlYIEVoFu2xRr8b7eCk7mYC7HIQEej/354FO4ZLLFJsVr0/VLOAizYw66kr
uIbscQQ8pB8m+R23hQv11g+gJmI0/0EjJQdctGWa6WQnCBHgCRcw228iQZbm4Ef9
QNJ4ps4EjISBpfUT0JYrUSoHvFt0hMbvGuQwOJsPWMecd8k2yh2tgvT6GOAH+Ute
F0QC/4ZjeOMgBcthePzy3+Y/oTzXeeO6UR+ikmbQXhitzc8f0LmA6gEBCr5Q3q7u
iz9kgQ+U16lgFTAZAE0GizYK95lwG9s1rKfMLaNVrWP6vB6lQGcPe+hd4ZvqJenz
3I01DNhflimRhzEur+ftv8xZqwruNPJkzQ6jB5omz1Zg80j6CV5tvDwnZ+efSB9G
krn0r1dOJakbjD7f4VjkQfNQfMQjClehbLJgoVxAmaj02LAM1ZKw9vLalc6wWALk
PuMaztkyUFHf57QgPEz0tpSvsGOaBDS8nh7UyepUQpqT6VK4vNK957J6wE8TDUi5
z9vT0gkybGpxHGJBTmocNaxjt7FQasiuory5zASRFv1y7RrmV3nAm4Kfe8Gdm/QH
ZbpXDfq9S3sSPmHOQlunGJDcBaDgnVvi2H2QRZ1YKzbEoG05FvfuZyLZqug/dPzV
BJ1aKBPHC+8kOdoDvdJAujiuy2rlRk0slTVjm8/lFbUQafRoXCFnw6QPcoayLB3u
Hl2BuUJQV+iwmUcWVCqSqgsc7/iPzjdNu76Eo8VdAXkDA1qyeNbI/23F2Q1c2bfP
haG5SbIt4ptAUDpoflsv7BNgyAhXE0jt/p5MWkN0+Y4nc0RKlBVHeXXmKn4+CuKD
dscU9ubv8XxesA+G75hoIgHD3mTVEQ4vxs2Eq7PHKBAmgtt/C1/ghBNVRiWrq0nT
OidFWN4VyGpfnGPq3R4VcQeWtGoBxH41sb9W1Gc8S8daP4n5u2l0lZCK/lKIgqEM
epugIhkHELD+JFYPuI6rlcNXlJgORLcHsaRAt+CpCQpT/5Y77AM8sU6VyY83uKvF
jpbdW9gJof8oviSK5OTJzUppXfQ62kbC9kLCVJhvZ392PionqEfIC5h2KpMpjGHK
CujD+Ivu028l4HNfvVOT0IGA6lfKvtv595NAVksEclYgJao2DLbTY6T/MuDw8uEa
NzjW/ju5SShIe0TlZ1PSvrpFgvYRfpprm3b2kH4+v997PKOU3zEhgPWRF6E+YY1R
Hq2WE21MQ9MfkMAvxZVhUYCjlIpgD9C8JqYc5Ze1b1WGRaPVhfiuZZaI0YBwFw/h
lMTjm07NYtn6MjsuJzZLFOuT7zyUFhHm49B411nOSOP+KQyFneTCiECwMjlqpHwW
rZNCTxsLv4vJkfO31gzJ2OI6LKzCgAXZ55TUjj7UnmjTBspkNHYzM/83c+oRx8R0
iljRxjIWzrWB0lo9pExlegeO4tzaGkSrxMRSVQPcKOAQRYEo1Ekk9SR3AvC2Suzu
2XAi3i5yjSPG1kMPnyyEQQe7xdkxpPsT5nA/yF95Ypc6t+I2LFKmt/wWnkwpxN2L
UONpKPmQzYu4Qw0//TX4crFsnmkTqv0HJVc9IvOjmFZeV7v9Xi6MRGI9YJoymBUk
er4A7XmhYUySJujN/nQKtn6S248WMyZCA+T3iBfF/quU7f6awZVBQSUBnmcXOvA6
0OXMy/vbhDgbDp/GfBenf9zXivTMmbi2s0puWAd0R1qgom0K7BBqpL2GJSKa/+pe
hsNGciLDRR19Qx6NlWhvaKPDuV4St62+iuSc7r/kIO1pWrUKgNQtFat3r5w7JQ1y
1orE7aqy8bsylHUMRbVcTpgrAjGf5lANJdHTC1PmdN8FicYU2cZn8QEtWwKZaJ0W
KJaiWCpTC5r05ELmLZ1B+QiF6LqCYKBpMqRmD8Wy2hswQHqo7xeyPwNm/UwzFiOf
emWp0uzJG1I2tPSLes59O2huA7LEGHgo64BNvorG0qGK16eukgeJm3qjUDi6MJjC
92i1eo6NCnD6BwbSl6KJTAIMyK7sM7kE3bFHyl4R608p3C7OHqRB5iCT5kS4WT3a
GIvzbwoxorwPXpC58H+IGwTaRwRkcGH1mRmqWkyDBSQ9XprS5ePMN1TnkQRc1p1B
RgK77E8rU95G9lDcmnrznWGzmpFH+QhIe5h+27KuECp44CP1dd4RSCyv84Cahtii
SSwz+eVwEJDqnjxyyoWfjWXDG3JN0+enoAFPADVQ2/4bVLKxwUFGQbxCSUSoPsfY
GKr7ht99K+67MaSyDHuYibjfmR7JxwQw8yz46QbdACDggxPkFqGdcsqtDFZ/Mzat
X6jdqWo98DxA9pqtIppeBCGwjwJtR13Q5ZIA1dgGobqMsyPap+V2hjOatZJNsY/A
9gpa3pQWR6DevPH1fuyn3MjzOrM5XHVfzqW8V+ISKaYKlzC/1fFG03nh6CAnW+ql
feV2V7AsMIlL2xV7OB0Fx298M6E2hE19hCazB+vSqqJ7XUBmHpzB9zNCzZ2Y0bTr
quxCXmh4Re3JbZqvqDHNuZ++LthxeccCt2+XiW8jHKe+DjSnJwlrcXZt3vqAsbQG
gO8mRvuk9JbC3L3lDFRcpLBzUkuM9Oxwqz09khhJCgnQ3voJ6nec1lDMT9OhjsBL
02Vd0ZWtujP89Jk1JxfVMHe4wqvK5YYoy+tmWSiKYO2wir5yeXSUbc1/jehkvzeS
ZDGiG+po4OKy0en7oP88vISCGKZ1TaPSBwwJ07b/FwN/CACYZKVJz9eebS8KRHNn
eXC4De0JFu4YciKZd2WoeJOJIArq7JIYGSLshQnaqKcSgpGha0lEcY8KtwScSudn
dTeTFKLeHfmJ19uUoO8trLV0c5JFwMlnAdg1CCgW2vpqydDbjy6Mm9N6vP09/4s2
i/uM4zINhRtHryprHkryrQc45YSOojAMdp+1MY3yrG4n0W75peu7YKB2hds46tFk
wTDD+DcNbq3ixkpOfSv+wFJwlU/b0W1M+V9h16kjWQNjbkRm25brP4CNLRYbGYEb
2e7yyn2i+2i4TJ1vCQkJv7ZKxIWowaXjgFrjXUpJgzkvfvfB/bj0JPaw1P6iH8FQ
xkQu6kttzVIZgUhxXQkBhx1G+9aNu377mpDM+xljSNldCPupWC9xZLo/duiA1CTv
ZT/itGeZYENpnfQBfYn1LEQ+YZdjIdDsbYchLRJCg661VFBl9rD7SQXQyx45ono7
4JLC85TZAnV6PXhzfXBy4Qr6DQt8TR6SBxvk3sEN6mCp6aKoCFpbYSPpeYrWP0jQ
t1MAv7VqTCvmHRy/Tg3nDFV8yU2929spHc7wQjbNB30z3Ss54H49XtsBXHpNTctx
MU9q/P3toUeNe0iLe8LecwNGYyKJ5pCWF62IhrTDUOb8fsp/pBFoWinrEy+V/ed2
EEf5Gtc/uyLR8OS8rLtBivQuzK73RVV+G2gjQCR8/wjT1MZv1fdU0N+34bshThvE
YHUTUVJE1iBW6CG51EA1freb0kZ8p/EjQS3KsjshGHeYdRDqzAU0Edj75+4mHngU
4Iy1Xv69lCnmTv4bDTWOPmHBsF4t1kJjw8Ug9Bti/5ewUjvfsyzBxf6BWxYZEo9i
YrNh5y3HSnXBxzC4jVQ9WOKSDKXJA7BF4IlHQyIVOwYSqyqcQqWL2Wsxi/bJ+Qfl
r4eF5fyQgF31LTaAMurPbDzWj0RDzZEedXy64qiNWooXWOb6SptHiQ4x3FjXuzWd
NoZOqyTfZLhCDqUrWpzmcpggf9S4QX70DeD83rDg7iOH1Qk8q3m4h57MOCaOjlHv
nN7xdBJsUG9MnZNzuiJPDxZpLHhwrgFIu0NF/5wLVvpeolUBWNh7GVHg91zsDMsa
jbRwuur1DsRxRu8rAkDFpu5LD3BqjwHQP4Z8UuCfCtzOS0Svl70P8xpIf5P3FUCD
CSFwPy/atvWcArNJrB5UtlhwDw4s/JHHH24aC03nOQ35axjRnuwKBhK4wS1xRub7
uGHSwIqtA4LyTKPwXVitXA==
`pragma protect end_protected
