// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
CKA9Mv7wD0pgw2MYVJNX2ReaUWn0ANccfrciwgOxkllwMxzju7I85Adf0Fc2lfpT
i93s7hx+7PlSqzohN+EdNhYiNrvWT2FWeXTrcgRKLftkuikO0uQMhv/y0A8a45Rd
1n8Bgzecrirsrrv+rwyJxBlR0KmkfNNq9i8hK/KlgkI=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 4448 )
`pragma protect data_block
ZlNUyeHPkvUels65bpR7Iu6TFUQnwdeA8uJF7BEx3vl89LK1rVFOeXh7h3N1O+xb
TcKGXefAq4iWQ7FTTZqArDLRRq5/hbso6SxOEw8ciKKqLJloGlWP2Ve3Dx1lm+Jv
n5Ua0GerefSQ+eKJKUBhCNX+dl7e3JXviPyP8uTcR9gjlgCgHMtEpTDxpdrPU+TF
bCeBfIBOXDpW5Y1A9x1CuRBGrC2X+oYPWROaWagUxxiyBHEPZi4ZoWARTm6IxB1H
FEUGtmF1xxLAwbGaDRtiw9JNrV6sloyHmcDkFl/JAUFeIXpUqPcjuhgze1dynlki
HxRhlk+lvroA0zdoR6OODmy+1hsQNXMz/qj3OrYPl3CPq7MZgJFVGUADQrC55seE
GpdsOgpwxs+F3WrR+UjDdCg/RpGnsVyB8RE7klVAFUkStkYkIBYA5gi821bhxwCI
8faN4+uhCoqUDDUlh1qs8BJH2Ztu25xNwIsz65ITH8nny7XIXDDDY0QTLqHpotZR
TN8zAYukDf8nng6skIgjN7wkOrhSUcRVmHsEteaV7DCLgKAhigVhtH10xFiN/KnQ
WjNPuDpwumgV3LoMjGMZ5+x2RrxKk/0CXuhYIY+a5K+CVMmlYP8u0L6AZQbS7vhJ
lGYZJxBihoGkBYab0oaAphMsJzFMIiF10665yN0fi5GaPHcmTNHXZE+g1pA5FJ68
nOV2zrJiNfGZhoXjlPpWji9oeUCZgJHMDB/Rak80O+d69CfkcnoRF3LeTmxy895/
m6EnTEVHa4RY+fdXEal0drgV4IBPj9j4pbrn17vlw0KkVg/kG/Q8ujBi8F39e6ML
Dq8hGS2NCDVBG8GW5m4djvEo1H+kz7FkoUz4sWzKaAZC6Ys4MgwkWAzDAZobm2E3
/2+na4TWP1P+WNv/YYLSNp/JumX5pp1wgTtvPcnrkM6nkVhdtk3dqBYayq+UyclQ
FdD+bA8huaaOy+UyD966mKlhQ5I3BB9zjStHpYZOk2PDowuceG27LjDOTZJijmBe
bMXJieuA/FF76nMMm+spEGPwGrF0SNE+ywi/lT81g82yzNJzOuljiETIeVn+F8XT
rW3Zhwobk+0i1V9HtqqHkj8casWHmQHOKoCkxDfNq+S3solHd9wmsNyRmJ0Csj9N
DeHtq9mNsfvOTFDQI++E6muQb27GDbWtxIq6Ytx1XTwvRUBV6O1PenumBJpwB0de
oojV72ZJaB8IXnRanK2K/s+oiwTrrGtVxuSP3ykEQsaKg2tdqXnr9ckOH0APw90W
SFPAXdqAlGsTfBMa96F9ta9y0CyuQItGA9fr40YCui4XD3Hjw82RV1UPVEQSh37p
dSPZCKOstB1zmSXqcFd8y5RFan3Qdk99PT+7Tpk2m/OMeIWhoVWik8eDuTZSv2C6
dGXk9/ED0bZ9zqEdgJmwBebcpJMNwYsl+8g8lCfL4Fxu3Ni7j/cASo7dqDuPYd/M
Pex4hGqyvi/FYo8oN7TB6+IUmdBbBHnVVWYEwO3Ly7k4OOzxF7QIH6hqr3NhPChc
8P29VFoUsQW+OD2heRlo5NPyko/s9oJCYielIAv+IfJ1aWP/3/ErusT7+usNTVUi
MvlU2Mcog5u0joDSkCwc4M+LHm8viLzRbDX9p/3WZjELX+xJ/+i43OP0kFrGooH1
wb61ysI79tM9C3piBVcycftGMvoATiNJGxMu67Sr5M6cEG5Em4rv0/+dHCbXGuUh
WKMVIz2H3OVqix3l46xdRw5OKTrezNNjwDfWn1e9+ywXie6AGAs7zKnDix83MKkD
GZIoi37MJl0yoau1jBbHFQmNZ4yX2C6rjkloKpk9N6IfeGFowFX5owasyp75iYd1
rBx+ApjX1KqRZzbWgh94Fx1ShORKa43jwi7GWkW5z9AlNzgO41Fc+fAbewA7S+HS
JrQ6GWdKfXin2zfTx6pUwD/hIc8IM0X3/CMxoR18LaRSGcbMtyzhnbSA2L+MFjCG
bgyxLzwDN0kXYnPD9w4OI6BjIut8TcseT7ycyNvFTs5qiQ9PBXKX7LtSqOWkQHmF
TGZgc0rTW7axhmLOVDZRJ5G7T8sePsQB2EtgSPMj0OGjtCL/ySqP6w/gkdmHLqSv
wNC2js6yS14JuDr15VLnqVmzdMSJgI3TYXLvBaGT3jX7uWyUl9XwXDALvCN34OwA
JKKMxPPdJwsN3mQOHjQXIUPl/USGVThKLekxcxm4SvODLUWsaoSDe1kAb6NJdBsM
49qLkuxfaFrsBJ82bYJzMPDPVrsJOGUQ3Vzx9uWM4ZaJP0z3zCC6CaFp2IrK8DHL
VrbrXRO75a+/MWhcJhNFjTA5gQleD3/O6TvpGyDcQOX0u5UT9Aa6QY4V6PT9Qv61
hvou9+2nMQk4OvheG7ldwA2CjGVH8CcpRS4IlWrgQFzy/bAOoM+Qvu6X+R/2vdb/
BBBBvZgEHSxmAucCtwXDM0eW6wSyn1B0kTWOrQd2inMwoUFfRWnXFFdEreedKFUk
FKeD3B27nz2Ry/P1IgZ2NfewKHL63CAmiLKTJEM9Wuseva8X5FGFojEJiBepA1vd
evCsJWW6zXgivLXYf6e7ySQV/js+U0RxgQ7pudc3Fw4CFs/Ssg02jQC59YXgvuwp
H/UEqlDzvJXgbko4OqYhS3iruNfExRJWIsNV+Oq5O2KDNTxJlMp2lT19lC3LkZTY
3jNulKxo0mkeRweAMCF01Yqu+OYFGO3bATOZitFl48BYc4uklbmr6+NW7KM07D/y
erjZOvWv2MkAQNNmpYB1fV9m55wEW/Fct3HopA27yg94gm/ExDG+RaD1ddfmCBfG
192ku/2e35HGSvDan8soL8R43nwNVdOd72JOzAXGfyYHzy4BC2sgeuGr3mJDZaUP
cNJktJOg0UVZhBdFYMzYRoY+2X3Xh/kR5Ux6An0eJ8o0jN5Gxz5q6WOtLuSiSRJa
6Q8SfFOwtegTNZmLgCZJyUOG4KWFaVqXnmlbQ4pQB5r+ybEq5eI0SiVmQ/U+2Etl
qnLuPunKO0zuTcmEPqfBcgYBPEsYMK+IzjFZ0wCjK8sMjKgXsqiTxpBfaiVukCHq
2Ci0lxL9uQONEGnX6/py8/9XSBrYwLHSRn8K0XFCjJSYM/+IVvoNtkzb2GyOmtMG
eQBFz6+Q36bw+g3uwPl8irFh94H6f9A2/xu6VsK+rcBl3upSHmsUYsfGjk9uqHkd
quUg9In35fFPr/ELtuDZk8DkdJSsnEdLM+jIBVLQdNfjJcMflSGuPM1hRZKb3/lW
J3ZlYY2+Ft9RoJOb0YkfdOzkDdBKE4garSH3WEPXx2n6OOQcdBx4oDD2/65zTuiK
V1KNboC14IkqbDPQSYowYjDIA6u0WwnUnwuB8ftDXhvud9zVEdJ9a7vDSKG4Wfzb
GGmS7CrAcpm6HTZumEzsCRHVPwJ21jfCk6ZxdM9dW5KeZrWveUdj7Qq95jeqFWhz
usKBz/k0mDsyo0IjVRv1WoQ8PzMyARJAa1sCO9V0L1nqCqEqICk9efBLxGuyeknP
3wzCtyFQeGPvtLAkruf7gv2otiR15CzluDNPY3E1gJYAKLMdCnJDz1iXPH43K4iQ
URAyaWwRDgFsF/b6xg9c/5U7c6tFdlfLZS8PERjugDuJrKtCG1j4PrSnGDDpOMWj
JbNcqwDRLmZJna+p74fDWng2zw+8mYw3zoNFRQcizF7PDvjXh853MS54C+tOypdU
OlSsNBIkGBF+I9zOYdvYdaV/sUuemNoqcmjB3ByJbKQy6VePsilx3IzMzdcvVIup
BvUFx/P9CNEx1ITbCThl3C2zA0xW3dwjjo6jhvRAl4YqRJMHiVbmrceNrYMmWOdi
jtc5NGXTJlegOJorOcmDMuKEbagPcI3z5+t7uQMLoNNvznI/no/MmnFiEvzMDxFY
wPDoHgvqCM7nTtdsvqn+pgemcqlS5rAHtlO1rnvnvYl75DcDaMynixEkL/ru1TFh
i9fyeWe4t3BB9ilAHWG+rFO3JQ/JXZ/hFwCTX8RDtSUjbQkFxdlL+JEiZXeMaB6q
qPG5efOuLCPNNqSII8pUp7fBRrT7AyB+1/ivgDSbaO00ZM13qlWohlly1AIbaSA9
s8vASxsDbm7YnvnTD7JbDt8lt1qoqfz9byrUcXtVXYMhNmR8qVUck29BeDMn7XYd
4GDeMboTJXpN3jgFHYBS7GtbGlnt0DVPhXjjau6SUqjTCmuG7FJGfLJNyJM5slt+
iNJiAIIgVC6ZvgKEgZ1ttfFkwcSaxAoEjdH+c+ZP3rG46w8VTlr2y8lEKLX/KNgI
l1YXsLljEO09vv9yfoVv0/bRHgYjEG6fJMxIVF/vhE4zN2zOxUL6OA+bnS7kwogW
h/wIG6cZahURnQz70PSLHjaLyaWCR4/67CFeiRfIyOsEst853+VEuhnFW05B2hA7
H5iqLBWjSukTfM7/L6ZRma2qMsZOPZunHKP2x/gVs+qCqSLzoKt1DVimbdHVZRxW
L3zUCVyodi3sXhtdFl4Lnvo4usKTkkZl2Oo9VAaTjZ29Kpcg28flHjVeelSHfuMM
juX6RD+Ok8Hj1hE0/TiNEfmxlL6g9OUJju4hYqY+EVWDOzYQLgEOb+XQEOfxmPtR
qv1YWuL7WkvXFH9XctYcrQybY5eo0axHRxaqQk+FXi69nIF7MB9GHMR1G+Af5+Xv
NJarrtqby2IBpTp8gyYCiC9uULGnLk1XHOSmjSMSG7kdhis69b9qOpncncW45Khp
FxUgVPYnKt50RNyqvT7iqq39j3PwARU37Cx+lrJaJUxPJ9fwlaq2kdpoGhzp0gzn
Xlj/kCLzAJSIn1i5MgYkgWXNjV2srI0xrIiAJ85TB9022P70mTUCfcideEQUzFoV
JxMoQc/OPC9RG5DPBk9mvRenOT3i74DVLYkLTnn2vXUioPYmz5IaTHG93pAxqDrh
vv14jYpTGWp5NGuX3qUOUCkcFdBtiEaXHTyMliYrmtvBEjfwAwBIP1aS9vtpEgel
kWjfGQojOv13tR8qsW7J0bzuZpKHLNhC3pEed/tl/ugetMdZBa3NkM30bMLcQI/I
a5kyhSuDoyJ6Jb0uWgCWCvGy0dD+DCaNoV4sNJ5Xd0II1IwwyEaIByTHLVykahW6
ubZGf8ijBBzzjDon26HJC//RqiLzomP+XGlyXya1VQz8UuPJhoparvZty3hE/sXa
Twq7C/cmqGUYTHfSOsXK0eGaPRinjjCHAs8AoToAttqxSXUlquXPi/Yj1CJTarge
XzEJJhGjexD+YR+tV8VTVRg5DXCsMJiFv2M0NVf9IZaPQ0xAdBPFW42wVn4N9Pgs
WXf7qZm9n/ljzYievP/EFd3yVtmVJxA+YHWXQ4QBwjEcyZmgmcr29OaHU2g/dKts
FXXX92Smhq6i5VSP548k2wiXeDpDJ/iR0Ngdfg50QW3v191S5TI+rzQoZsCnNXAE
aUVtrrM0Jzcgb6xe7Ts5fNLQRCtUzyzwEmoYv6p5KURIvcwimTh2XmB/Z25UvU4A
i+MlIOPZ1JGWbdJ2GH4anr2H5UfKQrTJgVjncD6PvlntzdSr3Mj7tzx5UrwAb/cM
9H5bNM0XkdINZQ8nPzvRbJAZbyD5EuFUiCry+3D7l06Cq85UaCanD0P3whXbkOcO
ekraYIQISQp5QxrlI50FZKwGGkgb36gfkTei/lZP6aAOaexo2bLOzADSUSwDA0ev
SFpspGdMQSidwjlj7qHouEAawzVZjYxv+hQjQ8qAa/uHilZkl8j7hIBW7XvInKI3
8wTsj69I06DiiV7El5WXkwr6up5hGVusfJRgxqqbhsulTgi6+PrE3O8jDZyIDMxx
3JkDW5F6Dg4XcZe0Gb7coBe/O9zVHY58CUes99ErmrjeSq0gwTHMEXCCzFpoByPz
TbIhP5q25unacoqeGi3Hi1GQ8v5w6tiplmjV5YWy6yY=

`pragma protect end_protected
