// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
vlT/zIBGbHilZy+gcdVGuaoMw/5Hpdx5N/GaW8EaUSd80iVl74cWvzA5BxTH0oCVOsRlCInrrw/P
GW8KypNXt5gVKN9yWxRWBuEhhM6LcaOQbpvVP7JDqRRhVktc69z29zzMSbw2nQTA4Nzv3XtCylag
6PnjzKCYoBr9hOTuECu0HQC4rUceXatEo1tnAdB0zwPG2RpkrHRlXNd9x/KAtCAHIjbJ7SNsWeA8
k/44b7NiU7492UPXUDAKNkcI6MbUgst2juTEli8gETK3xc46O/GuLZcKX29rseaTxQS+XR6xnu4e
RFTR6ACvbD/Gv4V0gSuVHHFyJGg3scuMBXh+Dg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 10512)
QAJ1ygpR3xg2UffrK3tCg0JXB0l5M/jltdQT8vX9/JvAENcJTyFCw9D1S48MNcH9MpKRHbTFG+dA
hoyRwghY54n3mr6K0w/FtUuJSvcKzbXFgeFjWLGbEeO7e4VVDvvmKVENnjf04vX4ycv3NY8COB2k
ILjGFem4X9QmHel/t/h3Sm5SpIN7BPG3c7i9UANo66mODcBB1GkJfGZlXZ5lFVj9MM9FwlErricl
oQgbQJdar8GMV4wa0dxLU+G8uQjFod2ATNSAT9cOwJE5Z1eYWwpJzUPNytUoArfVhtXiuPFb7LLV
s67cYcPtnc8T8XOyxgPSr6LQi8G2tI4/1KS4HgbeMVVBSy5IAomeim1qq2uGhgbIHQQD/onwODFU
skwfoqq29CuZXK5nyzQuibqSCEIQPLQnGj5yoX77B8aRwjIsATkLE0o1VP0zYvWP+R5M6pErbJnx
qu7eFY7cTBTPihTTS1CuxWrPn4d+0p/tBfmvJjlmjYcnB7gMcem6EcWqdkv4fc8FUEDAKndDyiSz
jmxnBJmmVRGL+jAZe4kXMtUHeiUttmPj06kAg24UtmF46QNkpoknK5wUNq29++Y4hwiVsS4z2/nq
d5IRfKSRZoKNCbb0Cm8FFRCTCh4lUlQ8Eq84N9KcrMVnEfIeNC4YxfZsuXEqHq9QVloT3/jX/eSJ
IKreGPSlzwvMqkP1iK0YjQqeVjjaONMbDK/fMnwVFKnDjbaGDTRVyMCdnx4z3oaw0MX7bvydV723
Efwrq9Tv6OskiRlQ0UeyyIYOsdx/Uk5BdSnD4BYk2/fFdpR23bSV72AAGV8MlHkpvEZcKK7p/Srl
tKmKsxIFZomv3UqZvqXezM+ZBu2eEA/MtzXGDKFNAAAapMKsjsl4DzNkzLbIZUoKAV8KIP+4Nz+d
u/vSLFFZl2uhgUsAZ4UO3fX3hySa0S30ukMkTdzAAsLyGOGuQXrYmdvm3/daqfV5ym0zyHKu7o1G
fcOe7mFJfHyyuHgeSSrJdXqTy/If29yl6KmejyyyFxE5FZPeIkJLFlhc3TLCnhvXE5WBFTvOCiQu
iTPkXPwg4d16EbLEa/5X/qIulNXMVVuHIzCi+RppgUIeFE6Lx2LTb3hfXd5gY4vBMvDI4y2MqL4U
FSThqI4En+bgxciYe0DmAEZ0LCDi3sMYPm654kv6CcF3IG2VhTtjxFgIgdEYt7r2roRxISWpJ2vV
RJO8vHj1wSqN4cgH1zvejT2d1pVuknf0ATzJwK3y7yvkPDysoEjX5cLioGGXwscT9a1DSVyd6GRN
ioiLd9Y8mx8nbVWQbSIk3asewuVrenMtIr7mHjZfyZs7klDrEWysCPC0OUjtOQLtk1Luodvb/936
zqV+a/QLkJUH3zP2ZSYDnZ6f8yl+sNbwAvYGUeXjEEWMjBAxyiI1JDNPQApdOE2wzI9zDg5d5+j+
CSrIqQM9DQO+sfdGbNOiXzyzw/Mi8eRSJBgkWpTPOI8WNqc7W8XvB7lX5KbHci+k7CD8EVuiqHeZ
sh7zDXRFMyQz0RtjyqKjI5Vy9NFUsAaxPaHBzQgac0sIF6YsiiIwaadFAQ5P41XcSMsb+THkBOpY
Th4xSwEPDI3LUF4+My6qscbRnwHgCyfXcWSPxgbk1+n3noenNR3U+gt3ZoNHnLGw+iPyA/aBOhru
tjyVV+bX0Sp1Ls24S2EZtfqN/ITMN7oc0gGOzGj7zRQTGMH1BIEsw5vkPkGVHBx2gA5MOo8tqeaT
e2ggNn47aaRuHhYiyqTYVbSoYqYHV1Rs484CcdxUurmplb5+CBLKqQn1iLsvvHOrMAEgUEvUeJ3S
Y8K3rTrA5Opfl4QJTWADCLS3FYeRzbaFHjzuf58sZ16k7qE8crYn4DwoY2wVitIAIA57NqVZggM9
JmDJDZQ6Es7MkPeim05GQqAewzUkWhFJZFBJCAnqaIrKHVNSVNbHWwfVwr46kNiLHnyQ62H1zfbE
BSshRVbNUOlvYyTEysD5GKpsfOtZFWPxL9rwWI7n3CgsVxqQ18nDMzRKffGLDRlXdwpUIOjKc+bg
2bULR+4KRQJesymYL8Z8NOmJaO47mFbjP+lgX2B0PI6XcsBFkcLvqYrS5mf1Rt6NXWRm/Evo7RQf
OZ0vp21kNHF2x43DDSAKejNgo3KnQvmo7x4UkgSpmdZNVbLi7gMso+aGRdHaxiy/vY0qNCRD7+p6
gAvpoiM6h4cOuFH8kVh6W+T9pSahLq+Tu9+KRnAeQlQT1kHW9bavd9BefEEhjiA532l7O82R00EQ
WiVHREw2qB3EgoKBJ7bs4Mm3Ti6aun7ruRqWsBMM3sLVnJa2MoDj54ud3xzjqFj9XpMmMMXSjLd5
1ByL8x/JLjcT9wojW0gefa3bSQyLw6nPnGq7l17tWQa0H5Z9ZtpBOFaoNboPlpmwGpsEH+sGDMK/
VIWhoNIXKfna029G23iMhpo0yX9r01zxrhsEx6qIdL1b2UozhjVh8BqsrkQO7+v5wGrhS/hfqYJF
x46W96CThts5gVrlSLy+mNlnjkI0Bjsu/GfFMzIYq12lz150U/KkJJcegHuwvayf2qtZ8EgKKo8I
Y6ZUX+STvusowaV/2VpPUgiQBuPE1VNs40ns4p2+2aXlUjnjJVhOPRc6ppybiYmRQB3fNfnGXwpl
K2+GC5lAetrR35KDcVDZn11lWgoSEc2P5RYW0vWemIQadh494WmQOlM3Z3zCuqRr5I/PsPFqhtmo
vrKBUMnv9DmPiucLZDe2dMh5qFW0g6t8p74b6zs7EQxJdng+tiXjJaa6lvNeBfv4KWDcJF9ybCr6
ZjnCdfMF8vOdnWgSkhThvTPUTWnMzg+9ZtTMbyPdI6GHYnPlPFQS/0OdKQXVym8IQJEvfvbafRgS
SiZzGQZsmjWoQevu1cmrXRsDuv6RBDgzJrcEsEundce3G/gI9nM6qNbxnMODLL5YBmvJ9MkYQ2MG
2xrau1cmnS2XCi7BL0lATgdgR9CyRHOwmc/TKs185+BF+po31KRUGB5GtPcVS7tpHdpukyLov9B5
nXkkNubwI9rSqA2iUrRofdVab/tKEW1Ke39pW8rPMuO4tQeJqbX8fVhTC8PlfAcyXpf4Oe8IYnJj
c65PXbjH1iAPmTJx53g2XGkug2NTtsfg3LHXDsQy0pbeMPwDDF57oICkQe9+TqmXnljeYphH9jz+
s1cb3WiyJagW7p5EXJlfNTbrv3KBF2Eze6rkxZcwiY3Mkdef1mi9aIpcuHzf7kUMnFXa/I9EZNii
CPa8ONLORlK3Ul4AKV0/5Q68MD6HTCBHHTqtZFDwwQirNIH09f5PurWXVWVabbs++j7uHjBefUqg
boVlJ0/4G+VRkFkDzLzPxK+n2wXyJMLvUd8SJ3w8d3+Wo4Q1QtnxTV7Pjfqa4UeGLKmuiC3WCIp9
v3zUO6a1qA9ZdAzSmNgTewvyCg1aoTE0wEvNGv49B6baDlRfWeZEkXmn3uEDM7SQK+/f0mYrDNaf
gqo3m9SIj2r+nSUO1bJZIdoPtImcERvI2tLO+Y1HB6iXOdMC93/DVn+O13P0ceOgjg5wKdLJvx1j
XPqZO/R7hnBpRrNfuNzKjbWiOY1UOuOw1ek/aiNVmdrYEzTe6YP/qicr98AEM+P1+4VuthulzMRT
LBEEaXPJjwyR6aWwtjLfm0I4BA+0+a7RmQPrI9CpKdD4t3QbvlZ2AAdPpJgQmTavRRl0uRbxuqoo
XjurWySlyBTF83SExGaEm/DgMxWjf8ddJGnYD86dxYOlfbIe4OO69qfVfM60jFj9LlsoWxJFdEmT
+3GkebIW5FYJKnr7cygkN/gLVVaPLAJkeHJY3TRNII+THG/Z0X2GCvdo869RUGXeKZYsWsJZUdar
P3JDovm8ob+sV33c/Mj9b8EPcubd4GNDt6qnvF/gSMLhwxw8uXk94livAvUEgXXuT/C66aQhLMDy
vZmZErz7CN1eafulp2JJ9uqAWMTisYaxMH/M8UMpR7W+hX9L81BZqF030mRR+sWaZ/+TZab0Rykc
2pr3tq66HcKBndMGyCzVI+98XcW2Jt/UGzyrwSzNUSu809SQopSY+JgwXCAbcpjne0sPhhPoFqQX
E5lA/ZQUYKeMjVamRFsfpEVNQDBPzUw8TakOdWGRX/9Ff7cPRfqpXEsmP3TntUD/vI6ABvPCr5iw
gD865JZu9MnsrXD0XWAL7lUuT7po6SH3QI8W27iAcUnCpJP4TGhD9FrrQELtVtQj9V+0tngKf548
q8sm5kPLiM4cBuQj+jxSuyJMKpfGDpsmQ8TNKUuCyrOVvB6LiT+z1+1aIZVO8o53l0GpqAJxY6L2
nA2kIajPEfKgDRQWOgSg3HnES72ZDOPsGCfoIOfxd46AspRa2XHODLAI9eXMMOgtgpWwbDpP2YSz
kT1v1b3dgnWMgVj8NndULUOhfeO8A2tkHEvDGTgVv8deQUeutuvkSeaHcHcKOk/hwOHv2UBWo6mW
7/19epBkYozRoMxzqSMGLqxXzazXP/padw0aFKjcV+aaAvjGXPHq7hHb75UsgFxWESrPr8K9mYeX
kY+LXkatgpJYeDtS66M/Chxyz8s/pFW2VOY6sUOLQ3Bm1PcTrh5WWpIK/wJxly6JC8pFNbUz2exm
w6y479dFb2m1WJCSkZzM8FY1zxWgWyoczs1kdX11WEcGVPmRlC+byIOPMY7fnV2GTLsD9f35/kAN
jnscpffbrD3TB6rlLaNH30abkBf2wRvig0pqSGf1ipapGdz//dUdJnMapZyBHOcQWnpyb3WhEkkf
a8Xj3rSBWbdd2/E8TDAv+YVAyYx1Yy43ABTsn3Jb669ixcOtrpsYlbSb2DYBGHlgjVTPdcuuau4n
DuMVgc7rPdo8qPhXb4LYpPwp7gQUu48jySqCxakk/+8WGes6LoCzPddJOFln5Tn9gxJDcorpzkbK
1JkeKqKYwLaxT2ypulCSdEa69OLdOsWpRraCNzQrivsFCRZHt/TU05JReqjcAClzVsK+TUFNhdCZ
vzYpm649w9PXWoSGiBZOd+DUMU+qksAt9BKDxaCOwH2wuERxcPp46eM/VCIAJVEF65FYEZEsPXD2
Z8B8BICeNUdfe2F0WkhNHuZkDdPBmjJttlPz0GJOCpjhxybq9d3ibJl2pb+8HsOdjVTHhC0pCj3z
XRkFyXcBx+WVhI5u/OsZCg6FWFNlUBNtoKdfHXZfgd/cJY9ni8vWp9XeWVKBb5DFUEqcgFdDjGAx
90SVT5AuDsEm0GPgQRpYrjScGIT4hNxljh0fNecwfuhr05myqkp3gwTRjpkNBlwbrE9v4l1gSfT/
mmJ1D0OzOaVhZZQXKvMWZPo9xl9PfiIXIomi67IBp5px4coXIysHtJnDhzLHQxe+osQ0zDy23r02
x7E6Y+hMIPOdidUVzAb7uxZnNB7axycANPTSJG5yyaGNmdBb+qWICRBUi+ofvw3EfmN9ZlnvSS/6
NqesSpg5WXJ7sXZETrX9pXzQkCcjFjsykc2rDlO/B4ygYcg0FcYVbmSpSzrzMJ5dGZKofFKAsVaz
D81GMVrTpNP2KWGqmSe08g4is97jFmadS4GvFRFRMIsaE6mSEVs/93XRe8SMgru1t54bVRZGOJss
uw27qyM+7w4CmpD7arJa5t4M+XzwWis256drYcB3dS6kKZip2I4Fv/4X52lo1GsRZ3Ym6TfOQU+b
j1Ve55mTFYp5m9lO+HAeee93aTxkth8EmxH576VELLYStIqwwl6G96EpBh5OL5b5FDeIZJ6LxUBo
RKm5pFe77zDGjOMOh5Zb2Mr7aniCyLTQs2gzFKkDY7zT5KSu836xposXs5nhmJ52FHcQs9zbWb10
84ErMx0slmkKDFiToxvtzDD3wELWCGIUm8xJAi6klaJtg2235P8tmEpxUfhtslr0v0dGNKuwc8cC
w5Tj0cboF09CwhW+B4IVTiR/zIXKnBDOr/W/gyB4vXFQay8SV11riFIfn77TcMKXUlNSdEco6WoC
4fQ3FMoBDBoR8f6LrJtKfsK24jy3l/8W5wnpK+cOLe9E57twZo1tFJkywzGbjNilCEZJJo+1WrgD
CmKv4fRamlnLs7qxC/pFaJfy7jYjboJw7OQW/hfIYsHvvxt0WUsDiwor2GRtz5NeP1jpTWQ5vq+2
4Foe5xRr6L3RYALhGqP47Uf5QkgOF9rxG2Chy0vJYcohEJPb/NJ0rqbxyG7Vg3lUTFkTqlZNtVDm
P3QN4H68AbgF7HTYJSgF0d9nfE00s66/Z3EtHUrI0ExurRe6+6tKrQf44HBm+aG/DIsU9G6eQhzA
PBbUae8xfcXdNHXViiLSGjsWWsVvVYq2UsVUUE6hFobmD2Q14Xt5YQEX1+ipbsqdoZgp489J3WRh
et8zlUHjbLlrNbIhMeWEV4nZ00/9Ksv5OUz/0cn6H+FAuc3W3VR5ieU0ERTcNF0b1+5cnMwboyPs
EN10bajewoi3Tc2UyR1fcH0RTknESSSjXBbiC5lREm1B6HhCQxRy5LgRhK7nxOjo9/I/g8I2Opt8
svjpmm0tcH1gt84ImZ5KQBwoD2+WUJK0g1CXmtT5OSse8c+dyyXTzhjTq2F8r4+ygCW9xmivvuz9
idMyC5W91a0B+jYQxD5mA6h2+cvAWHzlivKTuk7oyBGrpIAnJPmox53DtUVwZPfgQ7rKcx1H3fft
hObxeWymjE9CmmGNMcsRgBZwQ85y0XMYwl5v2pKcVIO/TJyCm1HBokxBy31pwmS0JqlkhVqHm9J6
FamLajY3EmZK6AANRl9TJRhHapa8JzLFZLCCw66ohMmAg5V4Mhi+20Lcqfqh2NMVTPBhPen7hrV9
85RnVhlPL0+H7QBaF6tYO3DE70owWyL3AhFG9ixfOjyWQ+9GsG7qsQgPc4AWD5jtoGJBuSU5qXlh
JGNGLpeysa1oaVW0SRkVFB0Hjil92JIPaEMWRQ4nTLNGxjNIrMUgThrKCX4k+7HHr0QomKL6ocSF
5/mkdBxuhxuCKIjuF0gwweZ2gITpzjAyhdat3KCNJQCr+fAv6Rfpp8hQ1mjKKYO36dUQZbPqrWbB
TklDYeoETFuT/QlZ/WSlM6CzH4AGuil8VvrQ1TFXMzhXWqFvAj73TNXrJ2P031rfMOWvUZwSxzJq
y2s+D5kbZl6bPRRYTEo75u9PpISAAgBjSnkztjEpRVUFUG2JGFkiJ3Db0Aa37zKasHsgPwcCWzD9
VUlNpccmcO7/owN4gvh9wCKhYWZElmLjXMUAd0MrS9L5ktDNLDqluHM2YWTpQNhfJne6o8WFPj95
RV5kWT081vJhCKfmZ8snt9uPqRK83ys3zsqYwQXmo+F8hJX6GgwAjNK17OXdKRNB+A7EVHeaCxs5
c6Di+I/TMKlUXfVmOmS7Bst2y7MqyjuavVg/VOWMTrDDbgpS9QlC2xkMLuQrzRxAoNMlvgyzpS6n
hOXc/LXtBgd3HEH0IDjzKUZ+0+GbYFbHM0XfOFqeAtobOM60QzTqn+kAkLYn1k4ns+1+gDOK8Hxt
LWNRx3tJYeG8kx3TiVY9wT8b3q+PuUtFkLWCIdZ438y2Yc/1tFPDFCkM+pjSQMSQgEccmXgJW12k
mHpGExL9HWzXvWZ4hHBVmoitK0Gy9YS2YmsCdBpoihkv4oeC/s8tk7F5owZKey4e8bsIzXG9xO7Z
PJ7g4Y1Fdt8QMGKZqd1P/0kMhiQakbTxZZj7P+0o3HR05AkWv5WKn3dYesBKja4oWyTBgfOM0svQ
Mm8IYO/f6FixKnor+fwVoKEsriyw51WCoqwZ0sr3akXJ5i+rKnt0wp/lnqKkLmRqLp2BftiwdiT6
GAtduMlMBI7EMP29CV2djYE1kTqOpGLT4MtbKY7UCQQRfvkYrAwzP8wEJDk59r2hgJUjR6yL7wLl
CXhMGOc2IdJQZqXup+xmljZf8Yy7clCRF2FfkNvGDJwpRX2MlHxy/ehjUyusjYctZsHnwbFmK99s
TFo/P/e3ST4PizgvgmZbOanIn6kk5/XearUJHfUfrm7raoGlVzuBjXbiCLeCXzbKlAdw6dciwc34
2DbgYDjzp7Pmy5LYQ3WEDKudtWdRZ+vbbYpUO7XtmyVS+nopINZbWvEp36GykJT016ryN0ijCCDI
31zr4gE0osd4vHORpk8DaTHhfys1EaI3XADMWZXbWh4bItF/snhyeYPT/d/8A4sa3OWqVvpoV6tz
LRh7RwEFrr8qRNFnfLVn+m1LncI6vxrCmU4BNOz+rvy2zkvFZc+FQFVHgUzJcFg1IT+DqJePxe1p
u1h+OJk7zy7SylqjjIJ1rdP2f68DEefR9aBIn9bSNf8B01YpmK8iQJu5CJXOSdCYNFzdPEHnaJu9
iGMJn/AIYzeHLzDapkB419Uvc4v24nb6LXJ/CFw/4EMtiAeibNpUczGF/uCOxZpW7xsRe7ZMXwc3
+kYrMhthtmPiNKFc/YmPkaHjEfoEXkKjIB9RpmUu03vLJJwv0wBtBQjWbc9UoAE6DjYR9wpnOpQG
ldjVgbxKH8YC2vrpBvqn2qvxSCOwAV+abn6RGVVbn1c3t4Oxu8WRyFVCj6k+Y3nxzZVJ9oWlxsYW
lOM/VfjbZMCOniLL5Dg2YuVd3osuoLQjnKQlxhb0gBuCnI940AO7Xnmj4+GIqvWvqB3JCO59Dymb
9eUKXyKpxYc+52SvepxsjZkQ/iR4HkVoTiwRA087NIgLy54pLRzODFY6XKtSmoGQAAyQiJMchReg
IvjPbqg62xXISe1EEe3kkf9B+EbdzsSa65qqpmSIlJqmjLClEe2I11JKWJ9W9K8pVke+mgCmrl5g
h65Zzx07X2jK3gNPxUtyS0gkIlxGQgWocpPCLxNRSCvwIRRNVGzB7OkFDvTy0ygGX/v6jm+FHoZj
dJ15TkdE7Vt/KFmqQV2Im4u8zsMP4F8mgOKBRuTixD2nZv9uUzv28PT+jkcUtifplqqun0hIBawy
g4r7qWAAHUi1KmaICpVpl2KcQjeVUJpzlt0Dsp6qecprEZH0jwMynbD4asXhhEL3yW7F3uGkHQip
+GG6ijYV+1Jv2CKEAVaIkdl2Vi1L+44NcYG2Uc90l5lq5i/Udn7LN8+apcKDIZGnt85HjX4cHQGy
G1zAsqD9h6Co2YyL7rMBBXk/qUh6ut1VChuxQpk1dhfvbZOnchxiUlFcY+F+qC+E1lSHdRS+HrlM
djdwt0vf8iSaEZCBY4r+kCLQAJppfo7YduV1mMZTKPv2rXGsBtju1jicB7TppCpy1/gOiiuCwJpB
imfonSSib0LOW6nYdSVNZsRilUBpcriEmisY9Bs8yDGA9dpcvuuzae+E5kjm6+U06lapgIHazKh3
4Kgx8jXRbpajeXbe+HpywOumfwYJVX1uvWIOxEhY/JzdKBjMei+901FQS25C+CguGhUQGayXfSm1
0Jr9jWRdycfU3KPEpdCT9S+V/L4VxBFzbmpUFKUpVUinRskYX+pRLUlvzqZW7bU9/0oVQAOiZ7yc
ulbAv6YjZR6IHneNLXxAygJtU9dADQhYUGnFpfknM+C0tS6wjiqq8GKsvh2bsBwkVg+KkfEK3eLi
F0zqwEfKQo+NfVBt8mjXruGtfHLz9hKpkZ4vom2BHbMYgDi8vee+aJWPSHSDLRnGxnsSuvS1Prhh
RXSd3yP0o09yeUeiATERZ27pS+EVKsOMawPkE/6Sm6TBe420WYmyoszRlIY5gGTEKjYFBQTLJL4v
Oa8cBoEHTiTbRVj630z3tHiqrN69LslrcKFKGuoY5T6qEBJl/w60U1n4I+vnLGi487wKdrwdCoOG
7f/MECSfy16Fr6fepgWzOLX4FRywovmgq1LKe+1Y9cjAh7pdt/Ne7YNwFHvRcBgGAguK9roKas76
8MNj5HHho86+G2GXvT9kOPCrpqW1iqbi90ASvKsbLZ1YIVJ231AyORRo72Sakv3eIn148Y7raIIS
qE09YJFBAjRiFa7gs8V9Sa9AA0oOm8B6nFfq6ObxLCC6pxrNRcay/v2Y1rKLTAF0T1jceVzvVBaC
tZYm8c3JY9MxAcntH2R+EjM0JW9Ffj5GH7QIVS6oaFwQirmUGEl5c0ZOHdk6SynxRZLgy++L8+Gu
yD3ab3ZgBZ1G9GucHZLsSor7VSUJc5L16yrA+Ru3h7UtuSYzmQ0oiNwS0crxCt+B8+nWN3tvkcFw
J7qqNcIs7sjv8BtMr3yDclMpRYtBeE+TyWJQaNJ2SFsanSBOuveXfCyBdA2Io/pGYZY7efbaFIrQ
UAOkn5/Oi4ZVdhY5UzUqr+WO57ZiOsgqp9vBOw3l9L5mCJNJc30HdTj1wiSGSFEEMw0k0Fps8A/P
2F68dx9AZYAnm2+KXBL9ZT19Q97vQGZDvPgbncAiAXB0rc+YCU0/eBISrXEfvgxkPVvdTX4l6MAE
48vhSEVwLYso5SRyn/68YhTvFFGhIxjNyioCesdzPgoH7dZpe+ssbgNv5BZ56sXcEgje1PafyPBd
aQDnNtUTbBysSRkLalpCnoNkduwKn039DpXf5tqQIxVzWQZVSeHgMF1s6JFFpbNnRS243D99ZCh3
HB9Rlu2ItXIOG/fRXatLGslUkxm9T4uYt8H7KBiS7wp/ExvRNxsy/Oo7qwH6aBCqfzhCDNoalxVR
rep3ZpgG2Pkr/PztBqDwhaDQmfRN/3GAll2R7D2+1w3e8OXe1YoxkK8Hgc3vPa1ArjzhLQ8Hm6gx
K/BlTve+VdCduhtP+IGm+APsriube9DA4z3qI88W+NPZy2dwQ5q8FdwkvC/dqPWplB2XoD99laIN
vxbWqImbgrV8+XGrvvFgAjB//wD4fls/VrRUplTU/Al3bekcO2TxUVu9yoo7zRkpRFlq0FQPjZDU
Z6JGlLKvmhinnsSNv/xa8mhDa9NEtujooeqT9nR5KE4IQSMw09Taya77/0+WXmjxmi8DZ/MEyC7Z
VvNaZNaq+qR62sy57eBYYdJ3bwoEeRS1EAqPAv/4NUt7VXcP1CI5qSeQS7EQv+U/r+x8cv2NCI+E
gAaLTQ6Y6UVmgUTeaGT2LCRofHgQNmz+CEXUCzGGQeGsTwgd0gsHwEKe/NlwYk0libO22b2BT6oI
gbzZpVv44vfJuHmNJeyq6QzQVoAMxCyQpYnzL88CCbDsqKieGYsAbHRjqR1J6ABG5IuWqff2G83Y
eC3TnNOm8Rx9Y9oSnFIzIzKkOcFocfiBj6CxohxhaTt8lOp6zlHx3RUim0SU0u1vpFyHes52HSDN
t4/PKkt/N5HHmhUKeilknqwEZh+Ltf+vFIxXEcycxlC9z2S3PQhkgoeebfw9HoFr2jbI2VILYyXE
9NqvKsDdVRItQnX/VqrOMS8f+Y/reaWfHL7AjH+Sf3CqrVXFIPVIJBi3NEVNvqUJOfvE7y3MEsKx
Br05t7N8WxZQYnpKm/1XFGh7x9x5zKjIQYDQACDzHH1kBiprGZwuhLetn+FA+39/zP6Wwk/nBOiw
Hv8e5bej1uiYZ2JvpNfYiigTr+JDyLCXCLvBvxp0PGtvL/+OlKWQpMBN70jHF7lkzsEuIizdfSbN
p00jdk2fCQsLTO3BkFZu1/gpPQmFz3KLzT0hQqvKw7S2wKTOnu4foX7tA2U/rloxHrhrooQitKfM
zD5uIdQHhY/xHxHYRhrfQK2b6Mxp6O85njrTgGB9sOD1e3X8qsuLRYyzumQkufTwy1VoP8cUCFbe
MzOfyQjAVU2xI6HWMVRe0ub9kvjoilGQkWV/GYaOVZMw3cKTTu8usv5BsG7gI6OZRSaefSSCk5/o
PCmDYjJmQgk5H65RGlA49OrGIOp1x2BeM1WkNJ7IHv/09xyoAWP8FeuJeDIDOAQAKfYLl5tP8ZlG
A50ZVgQfUiYkP7qywQzwR8QqQBhg8u19tbxu4lBurhb7vAF9lUGkNM2G51418vlKRjk/URofL04S
FC8XLTCReYpzT21PFnbWN76viicX8ekuGfOd4mPHMKYXfjm6nyvJZsNrbKP9RlYlYh7CWyGd9GdC
PWj8QFfa+mnN2XJ6tjTGC3QHeMZiOvWrGXpNEBsDgQeqMkm/yQ7dSJw7e6sDegB/EBpFlsnkO7NB
ut4/jQBUmxITAMEPqt2Se5WoS9gOFfJ9rAk4Gb7+X7hPOY1fCY4t2NTu1G+NniWUBrNTc0J0bQRI
Lp9lgVAaYJegNr/AuNMpXJ27DKd9SJBg3iur04v4ztwfofwlfCbDxSFAQfPhYP/i54yz60QhA90o
tQzK16OGo5xFlO9HXfwm8gKBWRikDmnAkJ4ko00aAZGrVL9DVDhVbehEe30GvDOTmEj+umcjzMEb
nhywgEk2HIIv+/sLIXTz/JmcLJ/bBlu/1Nrl67O+99jd5cN/ulW8t5nehZ1j0yWetyCxj3uIgqnO
0K7R842F6AvGj4tbrHBq3imhwTNiq1KhBjA8BS1feM1pu+MwcRtH1rrTCap6+YDLr+B5f9QDXKQA
8g+Xdfvh/cjEQdZh4gQLskFjvCFyjsDtiRMG8jpkrqz/WU2F+g2zE/uSqeKozaYrQWjac9R1S5t5
U9i1b0/MIarWXbDeW6D7eMQYlVoda5WI4Sl1be0CWTqUe2sVX4bC8xwo3ibo684ryWyldHwiK0sm
uEpoEhSUmhiWHu1GtopIdJkFe4v5m4pK1AigWZ/tJduY13UpwM07CzhnOEFVNJIsXC+DxAoleztv
ju9UCMleYjcH6jevodXSXkQlQlTLAIIn/B/JLZkIvwoHahqf/G93QhQPxUiNrNdM/9Yq97o26vhB
jtjYTtbmdrvmsKww58uFDVmN24R4G1uDzFGN0ZiFDuiHOSzkCnkqOPZ66WtrtnxA/bWRZ56o1guE
RlTe7dHGvScuprCmKGK+cEjwyNaXwBMFnGBbHRIUtgSDE02a6E44pUdouoIm87rrx0KpBJJNZwsw
ddZMIzH2G676lHz+OuozwoBOgwA3Rl4nKxOasnNQtIMTxbgss6gDIUEiV7O8HvBw4ysNHCg9DNMM
Hutxb2dyk89uoniZviLTdi5Gyv+2DXDdmZOC3uoD8nkcRRp0XDGFfX6WD4rbhe8ipOUKdXAmk6ue
JZH9EHvfj9Uivv+Y/XlTEH70NdS5MmBOFa7gcGIFageLHjTwZH51uflyA+vEH9S6WLXRE/J48V+k
Xb56OBI02OlzJJjdfdiHYdozz4tf3JUPlTbYMQe44gNtzTtPIPNSKYzO/0b2Wf8sQTvkONfWAg4o
3p7G4P4kMQYUBLyuj3ZkI6P82+zwIaabYOk+v1QHcdWNpVBNcWlSS+/OAoIFn6kJHGuKqFU9oUB8
by5NZvlZk1+h5GKLy6x8Z3bEr5W7m/ljYf2O2X4mphbbYhbKBFMqldvhoU/Zrvy7pLmgHdJgSRk3
iPCut4RQ/SvOHcnAixCTWvPsLgpnQIeuUPIhkv2lDkSWiRttlYCMbH9xe3XOQvyRLN5NvVXB5gPw
UWflyGFD+x2p+xi/okbhFAsPSMWPBLFcI4g2/dbqeKCr1EPbGNFTuSgJTPVsrf2jTGqTnVJf8X/j
ubGLemBA7P40/WF2Iy7wu02YDQwy4ol7Gf1jei4ee54SGMLF5x8fVms8STjSRfxOSTJ/dXccA8Oj
z2t30j8CS2aE8PMeHmdmLCEIhHNwA2/SvKB5sCnGWg4oIIclpF2otIwP3VyZWPn3hJhmVI8JujLB
OnyhI9nWSMeNsShMeL3jPV+PblPT/tqfD8wc6e5DR0xZz1SfqSZZdwxckrqzhwXa5QrlUmaqKGtG
fOZ5IWeN/5+WY0U8lA8BmNdGhXZvVuQ9j6ZJa7nZfE5cnDPvQIaDeDv+TzNwnXWsaAi3+ZTXKCS9
+XFlF1KdZw4DJ+UQCpPElPGIdXUX183DMovMs8LBekYfaugcPSlSP+O6BRTVwj2P5Imh3msyGgRz
m0PsgY++BPu5HG5eUXk1+t5ECb2VELiJeQUL4Tq71Icm0gWqy219fAMFRP9QaEozdCtLW1jJxe5X
elnvbr+lLypx57Zy/i7BD1Cg2YoeQHyr
`pragma protect end_protected
