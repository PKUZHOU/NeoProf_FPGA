// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
H8bAV2i0mV0yyskSKkptLfONeu4VPGA30+cgK6yUYyewqPXKWxzOYvRVOcLBQsIL
Cgsy1QruTSAXkgsS2qIVBRG6Lma+UfS83RVDSOqKiPGGiXNpYHW4190Il0enBbwK
fw+eOLH8z4EsFJwwV+FKlCiDcH+YCB0JhI9n9hDM4tXxRWEzi03f+g==
//pragma protect end_key_block
//pragma protect digest_block
EMlLy37/CSl2kRs9NsRakv7eZ6w=
//pragma protect end_digest_block
//pragma protect data_block
rZ5DfIWhw1AC9p+NLnLITKEWQCHm8exQl5m/wtCD1Ay5EaMjsOrYwISwQ/b++gT8
YXnLzDBvFyLCdZq3Tw1bhHyfMy+hGqjT8ElHQ7HgsE845usvTkOFzFLlZtaaF6g6
xDZhxZ5WuWAvhZGKkUjvAxt+z0tIe9iTRe/M8dtwO4r6sg2YnaOUwEw/rC2JAY2W
x6Men/gn/ecgKjkGi6ufvpB9eFwhJLA9/hGO7lbuhz07Xb3bS0I57mRIYExrHM04
y7pSvdECH7m3m3nBTZJ4k9uTSNjXBp3yzFJgczKISmTkJ0G9ojkLETBgI+EIEMpC
vKjOAMIcDp7dCAVTSUqQkKc31fdRE4Wru3QcpHBczC7MMakQbIsmTFBHxJGMffDs
tPSPNwChBSZLC4NYQdedqCxLAtLjIAxac7Y7TYet+uGshNW6AaX/qSmP8FM2u3JN
ZVfhA3BPENZvsme6It/GcNpvpOpqfisRnDCxwdjS095LN7UFYu+5w4TlndTpE8lV
7alYVzxpg09/jWaERJcFJIu35gJ+C4Gw6mb56V3lEYdhkRBOsfDHK1HBzVSZNfAe
hq48a49yROGNCWJo66dJpb/293KwUyZ4KlsNOrvV9KoBcvJ3jJuxbGAULneP1sX3
oowEN1fr1jPe2LOqiPqyLt9vBSaxhfLc+HGnaMD/Z3ZFl79O7Bko1JfAcqsVMbhl
/cjGk6UlDpxYMFjXOXoN1mNMtdpBtfeZcLlsof/WbZRnxNVfmM47u2NBLPIGoEVP
56wOwWpt7AFT72AVVCm1ejDi78AWOfrXHhrP6v5eifYrLR6ue81dxOyLPImIFIQ+
XmCxuMTlnnzGcjhCXygE/HR5akwZDwsyLFHM2ruectj/BjIRFO4b984+QqhulRAp
Kg33zGAHmdAtkKTiju3IgnCDAHkoB350h7ltqGzUudI8krnN9Rezhwok+50CEfRW
RB73PaG6dF4dYybSJhcILHlwnnEttX6Rlvz9kGFBoPt1lzZj1nUVAJeFrljI4exS
AuSaDcvItYtw0tq7GWDtGD3S+2PaanZ3yQlqEiSrwrkNOMLZXr8bWX9qEZ7b7UGS
PpHs66WcO7vP/CrG+RrF7DX5Qx74ptFFmKGBfVsfQMGzwt9bDx1OtCXP6xfuHHUl
5/GFgUsVDSVOMnj/UHUn5tEM3OTPQHnrdgpXOpQJu4klrnWvqVqaS40BaIeHhDYL
zh/OtXwed8tAgaKQbBLqYgutSQsZd77jDgWLOJkkG9CzjFmqGswyEnir0OGvyxxb
g8p0YtZUPjmx2riPq53KEBtm2I8GoFVKqr5sF5rHKZ3T8SsXX+JGIam9DN1HCPFG
zRhb8e55p2tXpJOq/hgQZJQRDIpJ1CH05YvaibdSrwV8jJsY6xK30OteCzIUxTm7
ucz164A36Q+C4h6cQIc1EAOxaTL3MkbZ4NF5N63CNobJAnfYHkrhS3MiURaUua3M
tgEtuddhXsar/Qt2i/s5Vuqybs7/q7DSQZ00UXrgxpp/5IrSnS3xVJ8X7flnbdJc
Tiusi1CwBYugh+43ibHUqcL9bDdk60tBoOZYzRGcx2tS+sqL/EjewO3ZkuoBxK+j
kC2K7d0s+Kg17nRo80LLZKlQR7tRBIA8UOibXkto5d+hxk9hKLh3KS0WHT4IGzsz
MGVIH+bHFrEeyeGef8wmlZENoSOs4Er7J4qjpeNhq1YdrLWl000FLIW3OBr22EsW
NuzK2uggOV8pJjQE2l16zsZ8mp5CMgaGTRMyqIe+LQK68h0jpmAupCE5lqNMyZqy
zN6vJOfOy87G25SvcA3RGKS52pS7dPig6sQxrXqgKThdb+581EZLtOa0D0zt92PE
PE3W5sCZjScy0H1DcVmtXkRz0Hyt9P9j38fBg3Ho+40Oo7GZtd7SFcf1aJb5KPGV
/JqEZoDvrz1jX13Fp7T5J0PEHrRdFRkesYv0txgEciHnw/gBiycfcjrajb9RrnQ3
k+SthK8tLXt0MJ5apOlWco4wpg3QCpctPN3VZ6C3VcM7p32vjyViT7l2GOwVIDIj
AVT1CA5a9TiC1ww7He/4+06yNNFD6HPU6HoVuL8mkLa5MFb+gVWD+R7Z7ezUsdw7
0hw9IpaWe47Z9o5EeTyO900/7sZAJ0R1wrCe9hGWTxIaE1oLTb390nRacn2NwGgK
pk0McMQ/zxW8Bth71b2dM+ZkhOKl3yip8fy/Nhbd4O29Gnr3Me8SPgTK03YfXNXR
dblun9aTRtfADQ1Btlk4lYxumCN+7vS8jAfp1Lc6IMgdgcmzeAUAKxuNB3NiQ41o
ryU5A8btAUZTGoaExenBbgT423UqN1Inf/WyOqmvHG/tbL0X9skHeg/9TmIT7Xlg
au138EBmHpI0Ogq46ryenn+UkDGniQxL1oyBZQYKMIhKJCGN7jup23OVyLoshmz8
cWLpi3ggNZi/41CMXlpyGT7/cyfpsUMvfX+S7IHVWpsvalHQ5meWTTdn+nKhTU2K
b/fWpivjbkLrhoBGrSSEGQa1CgXEztJCZirE/4t5+t/F0zgdX2b6k8VuwoNNkGnj
w2kgnNLNyXVORSS8e5+M0A2wWB6a72K7kLQQYOIxUDvfuabamCZtM+S4FJXHRuaM
c9aM54l4DUzR1ZAlzJLSyft2aCTW4hhxYEXh5Oh7mRKoElnscmGQewGcEzv/f5A5
brgDAWrPM5mvlJPWHo01QJbDFC1FuI5ZqaqHpEOOQMFCZW+5DK3NLk7Im5RcMyVI
mSVoth63VmnqIYFKCM4CQDyG7W1DwFqPuG3H6C9thbUSov5bZBzFE8WBE+J9XpHz
doXOGCdJMZTPKWTDB+ZgrTeMFtcCywY06MZx6jVUmESvdVsvg2DCqRmNlWXhKpDU
AxNDUixns/NQj6rSiYpBGBTbDZ7lEbQ+1PzTKDgS93eathpj+KKcWZgB/SiRj36I
uRUA/yj3fqnTEQOKNdSqtjtmmx8iLurDSEgtLy9uTOiro/4sghAlG+Jr75nbvuN4
cZjXmOW9/Cf2Nu6QBgyG+ZKhJ0aS8nVLEfjogo4j0ZsWt3+9QCKqbXhtoX2LG7OK
5WJraZSvY4jr8XafRrzcj8rYTFPyBi7e0+K5rztwGwNW/z5lRDLkBxXU18FT3/1n
uXMm6UBYDknL56xuUHHHDqMseUliATuA2MVinW50LZipxTkfRPZ+pQZz+P+uhMO9
uhuTladMAcP3hHP1ZpGBivz025jnaJFtA0yKWfFGlnH4uMgqaFfnQoxrvd78H+mU
VSaTZlfsGp05dhbEgSS6GXskGEy5Q4M/cXmH5KXtooutq7TTfAarry5nBOEiGDKA
YjKWRDy5OOcyKIeL7GuIgPolZbpgb2kuyoSq5PCqyZSLt99qXLgYlC8RGMqipS/Z
JwiTgBn8s9gYFAybnROdXPg/t0VlXDBm7izCcP/6VLxL64qQBcWKW+c3P05mq8LM
zY7uTxD+yRobPsWktNT9qIwmxMJg9tEVcUI/bJDilsb+qySXue+r53RwOiJDY+HK
wKVXGPCOkLAhdww4CRA5UCpVGaeFsbu4CgALtkAA/DTmKLBK7WriXDLZhJc+NxoI
jFxMU52f7ooO8t9OUwPmqpBg/EDBwhoC/0yQi30PRfaKGhmnbtR2N1PPqXKmC/Jh
1oqniriPuBX806VxHBYB5a6b5IXRQrFtTURUPniH5LZBG0ywehucJJrHJANrajwi
FygPn3RNEKwX+dwufiYYj6DEkqS7M/EKlVCXR7uA/o3x68jKFpEVX5djz+FLXXVf
/ztOmT35RRUtVjCurUMaiwIg1ocSdt2ExhT/fQtea19rbaMCbmA8M0b7+jq4mRPT
jxNvCWPcMb/uGCZtIsv0Uq7/G/+5vLNXpOsTt4eqDq2uPmTdKQHXxs+yA5MvVr1w
koym1nNazkzvb0xWq016tGzffYOqnDdM220u6Mg/lVdHxi3QB06mVcNzvfIDFGvu
lco31RmqONFXpTdP0NK3f6poP9WXhQwzjC3zZHtiqopooSg1LD/jtGvb5lJLYKmF
5oAMMUzBxFdiwBmlRAKSztmRxEZYeI9I/7aEP9Q4POQwP5Z25Mz8swDliCon0ZxR
fz9N/aaiVN3k8ouYG5/WyAPm/kmqalx1XFLr2q08QXXeMbgsMXNvSZB0fFqTAjyS
6Ucfhe2AvIKWb0USsE0DwcLZzw2x+jQBBq7ZARRDvI+0YWaRp5L977W0f8WQxPUa
WVDjblrgJmATf5zsyFliXOrHixhk6f5SPtEQLgJ3gRcR6FJgBs7e1rUT87HMJRmZ
nptGIIsra3N0qZxkRej+xnlOrUkhwbG7jlJse2K+QIvnWYH8tJMkucfYtAfBrzVZ
a7iXl7TzIO+F71/kM7qE6N2btx3yB3uLXKuN3ga8ApBEaOXkxIP6en/RXqlsYwNX
d0H7yMAwaelRiTVeTdLQiKs1stx9DGJ1aTd7EaLgzpXB7QJzoz6J/qpWdJvyBsUT
Ly/N63Rpfy39i/ZKTqo8Lwgtnsu/FvWrQC8sS9DICW7ZvaugOfO8g4RJVsBwapKj
qFk2/XWKuJWucFLm00/vHNFeAAmdI/C5+y2dbWfsGxY0RX1SxST8qt0Qabm/6qL1
aQUkTHalFuU4xNyEBaUga7O9xFr9Gj1u5f4JzI7Wa45oRCZ5dRsGJiEW8y3oBPmG
BeODpqQNXKpuV03DoOFCB9SG810QbdNpbbJn/i642A0Ww/Zwi35Oaojkn2/H4kMz
dAtXC07L2NK+BpyS+OeKLH9Su29792ZnqcRlpKImLyRL92LGGoJ2ITynexyoTv8b
3WYgpWKtROLpar0lC1x51RudVi9teuVuviNDtOXWn8x9OZIZVJVWCeK2VbwO+wqB
Yn382n+Di3s9L/Hug1Q1Htz8mYIp4o/YYLxHel2YCbbQBRrcm1n0k5uXUgVeJtu4
7Tz+Zcl8pQweITp4Q8MT9bbgK+SKa6vFLa7NF45VWZcunFXvPIjXBSuGP1JqWd8J
KTOajPoZaZ8kbvOOXuBmBUrwrwMgdSiETzvYClfsjGUPIHnR9CWR+hoRSA036pWU
YC7dM1oQJSWRbCSNVDnu5ewlAXQN+6zB8G/Axp7HTvztvkCP4IrDwYr1CjFGdqux
xZBY4ZV92P1OJO+/1tu5TI/MibR3ite27bAmsKDydGdtK9VzOyhFp9LszVGFN5r1
OLexULhkjRqJbDqIgCjRIZtU33UIows8IZttnAcGzIqZzsh58zKqkJ1s+uEeEALu
ITgwlG8pTz9XuSa1Q+pLsLX1MJkT/UnOw1wiz/np/0NqxzNe0Z6chMtWowga/oYu
oOGDBGYfj2dI+MlahTqUWHrLUd1gmWuwdAbZ7aqd3CGqeVUw68B2ZEHW9aPhpxM9
Ey+1vSxtLhb7xTaMKrMYKoNVoGbkwaq0DzW0mHfYawRbFAtC91qKcJJlWmK3jSfM
q7/n5QRvNznl4M89rR5pELTLkbsfJuvKKY0aQGLJMPYbGP1qZf6hKF8GVnVeB7Yf
IPfhlL1N7ZmP2CpfmZsDgh+OXG1x8+9raCjNlbtLsMkbflCK37jnmsaV+m9Yl5T5
JeYbnku9bULQV1d1oNH5Kwfx5opirckE0RIwyh3rAu02+Ci4bWrbT19CIQH1Fu9+
VzRCi57jkllFjZptXuFjQX08T9TNFHm43M0+jkxQK29IHJHAN6/T8mVTrWr5Q/cl
u899KQn9dBX8R+Ynd764PkYKAepmi6/lkGv85e7aQvAduuJlnG7hWL2cTgYvNtCL
7j3fAwwo9tMxoKKb2VAxbzvr+17XShMal8E/KQs1El7/d1wZBh3W7/pKoYLGXo6o
Tklx2ZlFBX6tqmYw5Q/x5EUHGkLj6zwOQkMaLTws3t/2TRwyDnI0SUbAlgxyc5Te
X2aG9+RxUz5Z1+zSQ+/JVEbPuYAogwpq68HG1zS04TKT8Sz7z2DglueDt8nUCrKx
ntdCP5KdiLOPdtyK793tAfnbCMXTHyo5nXg0TEg3JaQkRg1iIkSpb8jvgiy3XwXM
NrpLdEnZz8JEKGh+detE3MUtpO5kQ9MZG0FS8iKRisah+Y9FvgOq4YpzCP53n56/
lubksLf1nAd4U9VjlJlDwB0190bRFl+ZtKFLdwEUsWAa6m3SjrLo3icIG+/mkODt
5aH9atapD66Yibuj70ghPO0YZ3RbIsLW5Lv6MkOkXZFY8GPwV7m21VhS8F+4DCFX
3QNNR6gZovxLUdNB6aue7Jftg8FRnepQQTntyf2bJS9satfNSzUw7tqkwf8V2/Fp
8XN1naEZHc7D16ukhD/1huW4sQASCBqW8t1ZUwcAf5vd8MNh5QVU9bFPYwLf1UR4
ByFqxuWmMfXYtKTX3bTCPB+njpFzAAmvlRfJbFpxYmTXJKL1K700iWD2ub916YMe
DnANDHhTXwjg+2U+EStL094yip0cHTXxSwjKXod2iNBhix8Cn8/VBSilKxzwjMdQ
EZinXFS08t4E0E4EBQBmuRxAHSqk8vlnsnuf+c2TgwG65iXH0VC8e109kQt/UgT+
UYH06JJRy1J5ADjsT0ZO6nJ9jKwZX2LjEYpwsLJfeH9kPqIgEzTdpYmgddG0hFax
M7wEurDXusau2dRO2UhyursXW34A6/7pSxmqkiOsy2/PCXU4xQSq78LarMZaQQHP
6Z5g8OHh8S20wLO+6H/V9Jy1Mx6UK2geL3Lw9CAaigu4hOwFor5mAHn1i8pa79CW
DJEorP+6XvnR9Sq7uTVzmZsnCX9rz1UFykaCPeA9BYENIszgvFCH0c8cES3CeHvk
ropISr294FIrFGpZJ+ZA3tL+s4ITe0Qx9Mc+5y2V0/XKdtraazNnVPBkhQ0CuX8e
d9iMo8WWflcaFDz8tb2nfQq7wnlDI+bxLgy0seGNoOO+LwNuKSB6lrNDP6bv1sem
wAq8tvzVGiByQ8gvWkPWCjZJu82KnN+cq1DzWNMqRzMS4P2vMTJh5PhZI2jnaAum
MbqYY+JdmpvWY298WwMSGI7NOw8dkl/zPHcomHh6Gl+EQm56VeNdcfRxEIDPD8Yn
+wrZ08nbDuk2ORGZGLHxlRMS/2nkpsY0QmmxwiBAgMO4HhXvP1hBUO3eboluOW+B
5Fq158ECMcYGiPq9giIs6Uelc9q+yqK2Ez1X4HRJAX9+sk04EGXhjST69gClpd0E
EtYQ2AXw+6h3zEGZ1Aw1dFr28JPMBZwvB6GqlgF72W4ndfoIWts5xniHdSJ3Yz8t
Ke2Yfltang6ybz+pKm9nu8bKbwF/yH8kZpCinRH0khe1gyQ8icTKZhxnK1QZ5G7P
pidCM/8E8P6Xmg1Nms9bafOPYARquTLugXVTZ5z/tSzjhnOkZUgVsCk5/BxdXy4W
WXrcJN1SJ7Sen2iP2xFh2cFbUNJmj98O9JJd+ou1gxRhQOWqqxFjBRMe4s++2t+k
vUJJIpOnX4a/0E9vKn1tj1xiSMFhT+69RlObM5C9D7xVC2sALt/twUfkD9IAGKIZ
3xRVdkHECD1AdMqn2dAJIKJYBxtCWDX91mMvDNcWhR8WjeohD6kAHbADb2kC1nfg
GerKIh2kamd1CVX+27Ub+sFbjF8Wa7kBY9fAqnotrvkct5lKyVLiNF50xDZfJgwY
iWBTLVmvXPIP8JsemNE93fcxmila0RM30fCJm7km7NdVwYpjcDu5EwBo+1N2sRPN
9JFBhujpOmkGl49XYoHhGlV7rbDAH0s5kmQUvN6ict+SObDf4TWbLnpuJjovcGNu
dmqpqlmgI/9C+4+jag1GrFskQ1ILKYgggxvmC+91pB4zyjNu7D5qn9kr+4AuPHT5
ZJ6KHiwKxKCmz3LcJQY9nVF3lnME7td/Wzh2qSj4VVkUAR+wZC9sCXOOeKKBs2H2
SroXIsqCbOwke0fJ/J5NXSaUUFaBA6l5aCKl8MZNw5H4l8XcnqCSNOsIrD4/y0FZ
F0Yc25FYu4a+wG55yzQs4Kq371IhPMXa8qKFSNNUbWkl2okCiRU5DMd88OiYpqQd
FGUbms9FtVNpsF8XLDnp8yJNy54xmhc/ZufcstHuMyKN1W8OVbgmBD9qxeHy0IbD
aCl2z1ifTcVstb/hPM/LomWUKFl3nZIxvt5fZ8y1Ksgy0yttTr9+swqS5NtPsGpG
H+tm2wZVsk0yxWgOzJom5ZdEdr+BJpjd+KUnzH+fC6Ip1r/L4qqPDH6qOmtFY7sf
t2rDTuOrbEjmWWaW6hKLHQIEmiewap/2BbbTmsCoom4m8l4BroCdr2iX8ZmptJgs
t5Xh/7rlEaTurkCjWL6De868rUU/W8Yp0FuHlv2oeLYws60SbpbuyQuNwZBekzsl
ZJ7rRexgVNW3YFhF3NiX3+wWwS8WHfnS+qAP+VeJMX4MXR+zfMqvMgvR8J/7zA3B
zmrj25aZztd1OuxQbMSVnq2hg2Qw9jGFIOhu2IEqD13wlDVizRUxo21hjBAf0lLK
uLzblXyE27iMIT4P8B2orR9POXOTajldY4UPMWpmU87IcoGOdfbDfZdR78IuAg1s
+LvL3h8hvkoBsb6Pnxg1/CtJTZYfH8fD01ANtO6YejTl2VPpjLk7EiCF8TEpY0rp
2GNKVHmXeZp37Ev/sUJms2Q2JNTS/fJ3s8OgXOesG3GUyvhCxqtXMjLhg5szLhsG
qiG58NFcIoCG4NFWHcbeeLphBEd+b/GgEmm+S4p1vq5/SXIK+38Ts/tOK/mr1sKy
ZScACzwvPDZ3n10sm6beF3xK2MwkOnxGNVKp1crZCu9t10pQrW4ymsG6PBc4n9Fw
0dE6kJJh0A4nZorfmpeYOVzguvUHMmU/u8sveHJ0kGC1OYU2RhxPE9PO/lWFeWoV
YyzmlpCyQGKp/jK5cMi69kGkNjOI05AGDC+FxUS6glQz8MMICh0AuBJAsIDfWkuZ
80p3D/ebCsEG4NOqr7h9O/itqd1sS+jywQsFnAT5iQmzOTo0s6YPB45ATuF/gM1L
V1U8ZBFLztMFiqPmweg+ZYwj8slngHyVtFNu/ReLoq4umxdXRkSPurCFrHDWBY9E
msldwGwuvxqMZltDebmmws74owqqgdoNVLckz+iIdonWxmXaVUOijjYAvbieO4NO
WNZSiMNgs1gZRx9aP5qr987LZPm1Me3o0aWWnSIkxhGOGvSPbeRgQFiIGmET7O7W
O2pSpy6QSotVTtK7PUuOWssr1G0/s8PVUongVetazjPEyBOznSgvdPSkcrfYNH4S
AVOHoOpaosHQo2Yb14pQKIKeVmS4fedtitImgicx/Ys/e0RpcgD/y2MdevxxMckA
1WjW2BdxV7r19Gh/5Efs9Ua5srL7R8mkf0OIbqbVWb94UF1V7K/87M4Ke9Kjqlt7
qaB9uDCPEYgj3hGZRpQfqva2ild9gxR5xO6WVlW7rwnGdHDU4vaqydfXTOJURdpB
kRFeuRzqVOhZeddt2IVxYAHEJuZCXMR8Ml9YC+7rImrF2roqQpkHFwPBEbP3Qg4O
D/F4WBPGBQMVkRjwky4PMcdGp3m70Z9ptQFbEDE0irnL5RcK6lm2zLSQD6rgQJiZ
Jx+NaBpSKitMxFAinVGAB6xeymFOzl33suFKQWjBeCZYy7x9p5d3D8pMek7JAmVj
HCxidvqWwvoO/myHrJXCF8XlDiwGY4zjJ3xr14n8QA1Cs1siLnD74RS2LpoWz3PJ
xAhEoXcYVgiohohSug1+KVML4chd0+LtR6yQo26t5mazV2aIAu2r5ND5Lbukasv7
cIWuraATbUwNmz29T74zUr+8PN2zEk4hWcx72Z0oy5Nzjdpqkto60yhtLQQNEj7X
xCx4Mrf67o8JhF94FJFxZ4rEtXjQzJbFbOdrgNsHmfdjjlIS0SSFU4vteGws+xjD
XoFb4URXjMpouE0/l7sVTWI/tnUiGC+mkpKJhhPc5d2I7bhm90Be74VgtjmgMrNa
pWcKavB7LI9wsiq6QfIBQ+DRIoxCj1RfI5kLwZUnoX2y2vrCG1ETKWBoi0xMVPLK
b9DZ/+8BawUWlG7rjdqDnZ/12ODbBcKBXonCuhjY+mvRGdhijQMFBkOLqJf12+J0
IGIYxvzQndzTzvIBQ557V6k6+xnMN3DRXSGnXN5k6qm/AJgwnGVX8hLVdMBOVY/1
yZC84ILUhj/1yob+sPHKkcWVWupROBqJyYiJ5FoYfg3fiUpN4hlEwE6qjl6rUlOL
1FAix7+wdZiz+ubyK5iXjzgQy0VRA/VoXikwFk+nn8JX7SivNfo9bJ7sKSpssewW
ElVG1RcrEuWc70XPdH5+EVIaK1mBp6Q0AZmM1sBnzQiXvjMG7ufQi2ehLQ9FofZ7
+YQ1wwoixl6vLK3P4ANbnb7iKW0CfWfaF0kyjd73Hfd6uG0z+It3FhTFI4z0dk+F
8exxAq/lacAt4OsCsmvT58/PIO384iWx9P98UaPh4H8/sh+FW+S1dYsg7eRspwYX
WED/lGyX2AckpmmkCdZgBTDcUNuzG+FReKOkQ+mDTBsKV/CLWKv1XUC3QoGFgNkf
dwMH5gcOHXaqrjBw6xgt7gdk9JNfFNSzQvUBp+DAsiGMr7NwMAiVg7GbpMu2OETb
4ixdotSILGCWGcdMc1sEskNoCn5GcwJC7gJnMBxEJ+SR/4z/SVxA7yhiE26kP2RO
kLx5FXPizITHLfktmed6zj+UYUbSa3EDextNZX/niJ6Ji2D13DYBp4IXFGKn2NJY
5HamQGgax5EopfMniJ/5po/EtTlRgbHR9xB7x7kOwlQAEtFAcEeaW5VS3JVXmZRK
KDokWHtZVWNpQ5C8rNQewJUcofTTebdHQjuNGkAdJ0YyAoNWuMjzdUehbIRFG+FF
pq6CM5pAeOnqLMj/4rXKFGoL9wBUCkasaZIvIdeVYa1DtbRM1VZT7B9eaEMhsCbG
yH9CzTPQ8kHfXV8IxN4duoSmSIY9q6qJG10Tr1PWtH8nQRmeEp5wzyK0VECslpyd
D/TxMcxCGq3XWRyvZWgcRBnZRd/zgwCAQ8//b7qZgyFphDyazAAe+qSINC9EQgwj
Rhe2YcqhEjPE3paKq5GdRNza1+edEyWoiUj/hKaW6oq4f6tx1jNM9J3DH+4YZbE/
/x6sqnG3U64EaUxpEDh9ThIEreO6x5omWgjtUno7ca93rB6m58zOsqkvC8Lz3vDt
VMVbY65jukzI/PyKLZeC5bUlG68FYaAbcx3YUo1+NpKO9WN3kvYzSKXdBB4rJO5w
vY7IzCEVXSI/R92BKriGn8ja2R/A4Ow62LQ62SXFTU42LQn64w7r/rQwkPyv2irQ
KeNNNDFUs2phz+B7jxh+ZUIpC6995HCMwcJ9/HC75FLE0JeeG2+ofNzkQH+XWn73
dVudYPUHtIFT3nWQh8DgXhmsWhYyEs6mhWwYN72hQGOKJ3eIEPF+/Wwp+3SNc0qp
IeTanIcE7ArRT6HjKR5k8jsC3tKgZQYa9W2wQ67SYWAxIy+UEnp11Tot3kiKf20B
/b1rj5HTWUcXqQz5um9stuHkfL481hzNFukyNreEWUS9xjQ3kdcxEihSHnmohRuL
ywhqrc2KOxYm5OARw5gQhM0W4Q6nIHKIJF3AjZFc4Ffrzg/93kyYIj5V8bDKfnBq
oGNYZmrYkJvIGD50SQNpXWXYocGPjahRCcZu8c1hj2o=
//pragma protect end_data_block
//pragma protect digest_block
vYs21+lxIgNgNIq7jKrsdy+aqCI=
//pragma protect end_digest_block
//pragma protect end_protected
