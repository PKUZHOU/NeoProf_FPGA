// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
bcy0CEJLy6a406yN1FLM7jexZ6JjPCylWVtq38QKBkqgfAEDGkSNr1mefm7Z
JcjCU+ks3c0E2Gaw4GhN0AkFfkZBabw9ytLY7c9xIxyBgX7zRacCYJ1ZlYma
WUGymBA0ZHuE3ht5Q56Kn6sFmNH6GDNz5Z6FFQVlIxnkDo5c9c0QTbXigF4j
8O/MjU3Ra0jXfzHXwHbh/JflkM10KFKKBwTLeAPk28EOoBFL7UQCjlpB9OFC
PF9ztaaWw0anoLnzyuBV/TPp8ZQfqNRznx+cbtbIJaYQlZ47WLDIXymtYS6u
CGNsMPn1CVBNg/jS9N/U9CprhcSymZ61mX9cP+j3qQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
EqZ631DzenqzFs+M8J+fX3uyqACurN6bjZ6056M4OWHt3ePLUJjlvMC2OE+E
Qt8Geu8/0wrenPafjwEy57Fq0DcES1qJ765E30J/rSuV20zRe06JY4siLUPy
molsnShQA2kgpXhBqZIIlezWRYrpUCrto+Yx0BenQOkMnxn4iQKNfgdRdYGt
moI6IsxV3VvyguuQItTC4vTlm16h0/bmNSq6yoO27sAYRd10h2lyUAb/puj0
Xj5GXvj3wB8RPEAAJonzZG1Ga8UUfO9t82Dk6H4FkaOD80HtaTEq2s5SvvCT
DH9pd/dQlXGvqPw4VQAnezgp4KGwIeNOjOsdab0pIQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
kXM/LeJSRxZxRDa00RBJoTLoEm17FG8KR7tnow4xLmohR6rWnX/lLhr0DA98
5F8GZ8EKexkk4od9r9PoYz0Wkx77eFxo8+q4+QLT1YSsM3kF5gx1vMeAfxR+
MMjGi1TbDjU26aSWfHKa0c8rNMYRvW4Or9fJOXYTfBUKE0diEuAbO3wBSl+1
E/UK9mZfU6IxljIBZLhRnV0QFNQeSDz/IB3aeHCZe5ZTcKNXysPb/aTotnsw
2P/xYAyb1z4xi7ULMgdgolJF9Z6YObK/wq99vLhdO1k+vOgX/k8mTLl8efEr
ncP/cPrc1oAsYUfZbJmvLAnROFww2BWBtVZ1t8gtBA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
TjXLPp2RWDkls+JkAJ5hycn4xqFajaHI0RWWwX2PJ5e8vDoeCrq8eAUNd8xA
WjvY9Tyq4sHMbwmAsqtdly8elyn0lOT5GuLm//4k4SAO1UVvieyhC7AmQ3J5
eSAZFZXB5C9QmVCoBHqZbG922thHyvlAjnxSXl4dOm9RZQYYgF8=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
a20sT0Llg9umRIjJXtvCWbB/HsfNDC/gBQ0OzqI2BfcLfpzJmv31WpMpk/dA
x4e2k+tfVv6uwV5qRVVysSOzBFSLLz6iWsmNRPCju/VYRjKsTOlevoabP7Eo
opQxWVzQ26WTXymCZFqbTKYZDcJcSDHZsd2p4FFaMYcvnQxtDHZ7SmHD9XSY
n2FdkdJrfr5oGWFyHSr+uncAJE0TSRSZvHWy2BhxrwycBGSRp142JGbxwqsu
RAGp7O1A+P3Y/iLFvU5YYpldxEe4O7+Jplxun9LnNiTsQjGbSBWH+hJsFsm8
Djr3esfRRPnNwvbtBnF9aIq6QpltjVmlhGtBpXmYS5ajDXEw2vTHYV1Iddp9
0BI7OBPmAg+TJoE800JXCuNMvGDwykJ8s3FxdiSy9kV5ImB8x3Jcc/DeKW7f
GuwIRimSJ0E+eEqn6woJ8IBRqHRKEwNieJPYxc+HnNASEEDSrg72+0pv6FgK
AJ4vbn4fAOsWGZ2cgcVEoDwnnLd8wN6I


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ZAh6enX+h72rBUn2SxJkXdRNtWTtybk4z/WMC6L5Dyx8Uv1gZ8H+4AMCIusj
1/zsY91TJQTROJlytw+3mUVxhkRk8mQuNx/O6HoxH81pbmZOwQcA+qS+JT9v
yC4nD4kNJfaig+zLJyTGOogATUQl44Z3BfJDdIXlcAPYXcWABV8=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Ct/GKqcQxg5RXxeq18FJWgIYBXk3u+U7g4qjOdYgbIFrf3YfYcrakqFyTcO3
me/4ZaOt2fFnKp73bABkTZC/S0eCZSkwgZ13QTj53fkC4XWaRm0dN0anKj55
ERidoC7asLFoLmhapukuwhpd4/agS8ckXH11tBnu7FzhGl9KGUk=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 7056)
`pragma protect data_block
FYJoi8dGVcboFovV3Je6/voy22WRfOu1fAv0ey2n1HuGMQwEKfkcbnntTUA0
hlAnDUEB+FSf8bqNC18X966LR3IPR8eRlWs19SXDWrOh8dzBsLQFvbQipiog
TLJGBu9jLWhNXGNdTDmyRI19SeRsB89DWQA9ykhzWIABg5Z8aw2LJtlx4+og
32j373LtJ7NKQqEmbNHMD4qQkpKdGyFuPJVgSE/C8M5yEna9cAmom/DaqjDs
2F+uhMQTtiNM1m4V6GfaXCS0x2uKHojZS3Glj3nccJIp7ZZvcVJ1A9HhdJSn
1hVQjlQWCSuY1YSJZ0si6qOwCQqjETjpdeT5cAdjsqkRimjD9zZTp2p6M0GH
/DLp5RCPYPJKPLEXQ+m7irSERoJioH/iJQcKwcG6qvi6Kic/72oKvVEyC2/2
ZwhFYEFgIdLyqARMhBrzVj/+fon8LiYX3ul6MEHHzgTH7F3tyPB1iOA9u7HR
vFaayQYIhndCdfqnwsKA24s2kHyTNgib4p7sc4xi8OWw55R5ytysw+Wv0Nkm
tnJeMUGGNWkShGsmWY6YA/uUSn5sjkfxWka1C8kdPb80/FHDPTgnl80UHbw0
arx3q98Feg0zPnE54Gl40iJ1LnGz27onqbNDnDj0wBASZtws2lnUmGafaatl
/Hd2mX7/qj5oiKXJ0k1gw9FqF4ZcEf0DwctWKkm14ARlKhLMkHFTYN9o8bt8
PlvyMpPbJOLIqOlaPeYdZXfiCI/Dagi18ktGyz2vYhaXyWvHolYEEn2i6+Fe
kdxQ3le6Llx3FC3XoxfkJ9rvUKmEIUUSyrSwSfLS7InIp1z4k5m7K3aPDMJh
Be8KnhhmavaT0/XT07ZaVTi+75NZYIx6eDkT/uYnvsuX6oZ8yjo321svchgx
yMAeiF4YwHYi6kcdJWllfanq0GhjcB1wGUGtLCVYI3tZL014iGBPsZnUTGcI
qBXYj3rVditD7k82IEmDzPWivqiHndsAonQfyHnW5WHaZEl8Vvsbm/GwMGlH
XKLuWd2p4OowJwrkFK6c0tAu9IjeeMupDnGy/NxX+h2Lp7c4IbQNdrtFscys
/TI72R1YMEuPLbXkZjPUc7aI050CobQ+TMakxbJtVjnfiXeYMVv28hoQnK8/
Z6AZ5SMp3YquZtxYYh35ekJTqzkCNlpVvAfelwH8EuG4TYTxNPeXvnjwvRUa
FAuJX/vrDr1Fw7v8wyDha2xqSslRr5AEpVh90vQvMzHLAoAEB8MjupOde2Dp
YTGN84CzgCmxHHvhl1e93aB0kKSZCNhPeYYQoAutQFCWgVk6v+CHqn/blzfT
Ih+SR7fbO/zgv+FuGCMHCinfJ/BFNlYJxDmBo1Abi0+VQkuaQPfVG8S55+U6
niphU9xC7FWywFbfXNruZj12udVXDIhihwweeo70DCC/zDjXCzszSz+JUK+J
XnbLkX6QXiLMBEzkyD6MajK4k7G73T1gnKJnWDEayoEtO2a8MsO//uynNvWN
1n9NzRTYbxCClGceyIKnhDDkPVOJ7L5Rg43u1DJBr1a94esUNprBZgeyq3pe
TAxt7DeQE1f1q5OXiMRxxqyCBJF+oyPen7DmYyt/SYZ127+7PNJdGEjR+2QH
tGeXPta8y68a6Q6ShCoG3hqSonO3eEPvnafcLdHpe02yxI4O0HfS0PclMiN+
RpkYhM87FbRL3sLVs0OYtXd54RdRMWuGRYBrEvuIqYyUA96DAmnD0I1g+Ixh
w/EY1BuWMenrZ/ynenpo7xndDhYRH+9VfIehPdnj36TfG/VhsT5D0FF2Iplj
dSJgHzdbc4gxMJhRcx6TSVwWKAmgaYfHXN5wvCTxk7O4MB4A3tLbjuXkudLA
5Evzy7752A/tt/JwgtQXfzA6i4ORquWYlfKNF+N1iuPI/QS0WlJbSpiafvrn
34IPONlFfZjhE8X7rtNpKcKXkz43VV6JNYCT1bwSU8dAn98YOPuEbKNVJbRI
4zDuX4kIj8epIh2nUyj6GPcE8dqLlcg+QKYS9tBBWcLvtSTaSL8cyuJkQxss
RvwwYBE6wjoH9nQgP+MJjEBSalUGFiWnVw4IP5j+AonrKQUcKXPjMmeRUBpV
0AUtrBgnDUo4NszV9hVrT/B/5BwQdkI1GcE/IYMkGZg2mTfq08Hz1UddpSdA
IeIwzqgr2OtVcVaKsMy4Siw4T2PowoGnKEHK8twTZ4RI+jjKet4UgNkxz8dO
jocliC7rO8Cg+J/6BuTeDxhy5kRjJpCGNczzsE5q5b85oSRYxD1iWEo67IvX
DUWZT/2a7RdtDS2Kfw0sirAwIC3tT2aBSBUV9IDciXdMi48GV1DSiheV6Yn1
NlCrBQN4S1f9nbtc+PybFnaXFgoe1lAqz9PbDURyaL8gV2iIJuHOI5Q2e4s+
z3uMH+rDX0p4DG9Wy27jUq3KoD8bE7jMq+jCGse833UCRrZ+Rk3/vFT3B8h4
KZl4BErWcg/p+7UYGzfb9C/gzPjXsHS7/JmMMDxoCCzzr7fJke+POxwHtGNg
DGhHiFM8hvK9/aAslXtkgMJgYSZcOwT4udRsb6mygd35fkGiCGxaoEtVnzCr
r37fLmUA1QClXQ5oGNcb+QV7cOJsjlwMNYtpspJvkRjuLsxD2y2fhVvMc8os
84W7vfRQKKKdRZER+cVQnufojDB34qpwy4+kXiCGge95dCgRR3eu2HUye6fw
soAt9EKIZzoNGJ+hceBvBeDnOFJJ5lMfkoCOYBEIaOwyV5WKfdZgoLu9guju
YatClyP56x3izLfjUvYiiGBY1z0VKGORXUzNLz6k6/8H5zRfXetHemPoc4nZ
R+U3AC4Wm6H4NrYgOozndgM79c9rQXRX/RaGP816fQeGGVPFdOFKbN4aNIjh
/bJNTt9sZk7ufLlMO5N9OJGr675CgWri46DuP5PTJomiQp0WUORC436ny93/
S+FKxmEi9X0lzOIZOcm5mSFitEhuwcWcqzEi8SYJUahMBIR5bChvXBlJN/Rz
QqpkvEP58wYai7peWDcP5GsmLOoYMwevvFqhCxBLjge3oI/8dUGzIt6EW9Rt
QCTJiiFGFqxphXXPD1TfamQza2EIK5iwYhGNyLH7hRhN75O7xJ9VyoQTPYPY
IRsYv7nNsNbskH336rCTfntgvovm6SilhkodB9G0RATMGcwJVY97n1yvYJEt
wldyiY/a0Zkn/Fy9rxN//wROvkSYP68MzvXV7ysZgkZpUP2auWopYAFsOQC5
KHv9gxahTCCy/f86Ay/7cnwgHRNzyneS1bqBzrWvlEvnnZmESrP7NbvyQKQ6
6prupnpZfX8IktMtsxUp1SibWmI6jUnojsTfzKEB062PsyPQLRQv0zzrB9bJ
pY3uNWKXxBt9OYcFWZoL0niSGhOnLB5R4+3ETvM5RLCsVogCAKeEtCnxfTHE
L6BLRST+PftXaWuKRCqGDYXvtqtrL9GYLAa0zAiP0zRYa3nwJviUyvZv+AeC
wxjc/XwTu3sRraIvICZXZnh/YKkQL1f9tzN3pA2hSSBn4cVULkIlZ7XhFzWz
7cRi3ad52gDAqZhGIokgK/obmktNnitl3brvYbcEoUQfNfiAEbyDFJzkzcI2
JLit7DF6y2xkTVsXD8TG3E/9k//IxJySzgG9Tnvifn0FNxfywJ0cB30iWsZA
BCupdzEyChpI25t+vJFVPrKjb1bgRVSwbLBMC/aUymURMQqNuZ7yC2kezImj
0x0FuE5HrfloodnjPPhdeO7C0JXdO4Bv5GFS6ma+1fxo1PbWrzSFLI8nYi8r
SX5jkrySFBlyr2M/trtzFWhnM5RIKHAR30O48hpY743u9fnL29TVuzvC8w6L
LdqLe2M3RKXKMo4jOn4xZziLQiSSCPMO1xV/1VnVofw6YPed49UAFgHSgeJF
y32/bZkrS1v6/Ply+mGLCrGBfMh1APO/h7MhANSqqCnpNwo6kbDJ2nq9T8dA
U/jmbo1T84+jeIAPRuCFVwvZvNMPS5tvkwIv+5PqHOTBMsGHQkAxvVsiGmCP
2CW0u1bysYeSaqLkBWmm5d7yGnNHiWUfo5vCbc9q8+Ef32Or04X+hn6+z0gt
01+XPsTiOuIKhi3+VtyCwBntBkklzZ8gjeHwwmo7m/jHK074Yvlb6vfDm1bf
EbRBUrbSpY+rDAAHpoA6vcgUaY5ltn86A0C01kW+wvtInJXPOXGEOG6BpMbW
YsVd9591b/V/x2aStcYOE5XqntXYEKM1VGm0+YxEixHmS6CQmZpI+OgdQxB5
B6z71XcZpkHXK4tWOXd6XJRj9IXYrWNBAvb7s8uAXU/0+KwJ+Pb1pkgMBGFt
1rvLRZD2buxigvgm3eyIfXf3slX/psLpfE0qE6cvDT3anAANjzS5Dz0/uVdA
BgxkOXxoGev6ZrPQOUjMt/BkkBNzhh5VjPaFVBrePNUhUv0qlGTQd+eSsagn
RHrQLRLb/MrKQCpNNWGzAZ83hz+Bs4kapYkMrGJrPuSP7AfRsHY3862NfuPy
S1uKpmIOH1iEESX9a/aF91gxe4uTFZ7G88T0wSldZ8qxoAbwO8mwxf3ft9Er
Q0aen4OTTZud2CYBdRAv4HFNEE3XrS62UVurPOJrGnl4mY4iHzwnSm/vNGAG
xqiiwumh7Ig6d1yjlPmJLfa38u0wk0HzBsrZK4/m2CAl8Ykp4iHnWMQRyS5+
VIJyRGSEEROI4+js4ZymvR23om1Xb9w7lJz7hH8D3mlXvisWzQtZdbAlzMGN
QCLSRqMycecKKlhnoH99+H024g+6gu5yPDwx6uaiABX6FS2x+G3bQj+wSl3w
Bfho99SEjU3ZMdHewSdhC9yu/ZzrERCMViKLMwVNZEelM9h77iQKf9MPOZfZ
bKccLJYXVNNQI17cGNCi+1XUE+pDRgfeMrRlAOgroLu3iF4GtlPk2BL0K1Vk
sqkEWUMUYvJw2rAn2WDvR9iD9NHC7/cvTzjf3PRW9uRqyusvWRTvtOsqJpen
lnmhZ4rkrC/q1ovvHrekIA1fOLPITKW7WxhmUFRK2rKLh46CNZxj5nHikA3V
dNMcX6HFL6GR2vTZfDlOph1P+5EfLdWBpgWIpf/HKJMZD5HFAEn8yIdlGjTa
DyEXJLeHroXL6oUEkygj6JImFLkLC8goREkHKRABRBOPjl5uYWSovKFhjol5
xlwbbca6P5QuiFbpnurX8BrnSufjnK2lDCAf3UxJwJO/qldQs2ELehQeOosL
v98WSfmo5WCKuU5W5+cinCBW/Umorf4hWw8MQ2w4ZBGAYg/POnsBKpWmqe24
lmByIhD0G3FNm1cA0wjo43ZnVS2NVUqGm1z/HIpPaf44vcoN0qE3GBvYutPH
Bz5cZLIBJFlP1ldyrmpnjDFlFXB4SwMMfwkXVkqZ0VfN+O6kr5aw0LpE3W2t
rYssfymXmNIz9ezra5ODFwk+hJXnXuq7OvK/qbi5AFDEhdZEPj+fGTUmSwL5
r2FeRTYXRI9LTupIxFLHSKz+I0T/JC6IN4Od4elbjXypYHT7ru0ucDSHcPy9
fWybxxPxBTmOT052NtUcoR0WSlY512RkN2PFLbeGMYJjZSRuRDN5GMHInYbB
d5IQAPcS4mjkZktiA7mvc5AjX+SC3lf0gpYii03KET1kLrvT7+vujFzfk+br
qrbZBGqi4SwZ+dag+aDXWkNoPcrcVU+sNeLXzF9ipfGhQOkBERL4GY+crikv
oFiBUhHEJPLanJvPTLYoLYy2YMnVvGWbfGenT6/fM1ALxCZrkC3jWEUkJNc5
txSIvg6gHLqwPo7kLwumsTuUbu/aXD7Uhb1BURcWiMXmJI4WT3nBEpIuQLse
VMAsNrY95f8PeX5FJBcIYQ/Ja5gDS1NlXElDFer8G5B5IBKjgDzetP/upcJg
fjUnWus4afhO5Az1GD2FHv8Lwn1CBkl2PdO3SU2rYSrCyuyFq9o4Gmnho3iN
OQjeOpsk2IEu+2X40ihOibidtKQMS0JU/VPQJLKAXdNknLcNTp5Q994kkHdw
JfJ3iKsDOPvp/sGOeRp2RnHYGIgifaYyQToIjv/Y/dCw55NKitKXO4j5cj/m
H0ine1PuIGon1yZhDFqxwNC0flEN3UEBur25GBU06+BOJb7aKkM0jWtp+bJf
GNgTRURPZGTJtSl/Kw43UGksxh33rz6jHr1UF4tjvqPz/TOYYUcJMBEztdZG
CzKWnXGGG+oaks85JMbHill7KuYeZR1/TbgWSI1NXT5CsXBsqlzVmM86F0A0
BWZ0LVI2VJGxWCI19941q3R/3cY5kF1+0fP35xAICRRyqBDvACMSuSuCQ0/n
wk23Dj8mXhdSJi+JZwPOYefxaE/kO47865fv8pTY4hT3/WN6R9A7kBvEsWCi
c/idOtNxoe22hDqS34lxIS5Uw/lR0+oDNYySp6JVIZfEbm7fzGflIlkFyqVL
fr41GeIqV2TigROKfSrImzVIueSzqYoYj7wsbjchoVfb0XwNjBezV3Nc9Chv
KbDbef0xl/HYddAf/eWKX2d+JkAq0XL1QXHEMZFWo/0GtW3wnShC0kIOSE7P
NcV7nLxr0W8iAasuD8tmZ0F0XqFqrOw1OyrV0k0YgOD7w9glAD0ElFW5PqOb
x9QmZaTT3OsEivV5yapJl8e15S0d/4JTdOydJXhYBgKCCoKZrntLjTWf0CCf
n5kZnFL4zHX/RwwP9qyCxYJbpYzTxyVE9OB5x66L5JT88oNvYcLvYZvn//sI
8AKxIw9vkfbDvLY0Fum4U6Q3WtYlxVU6uSanuC/mHSLN9R4t1gDJucBfDmBb
GAi3Lmn/uU6ebPrhSPNRmQZC6d2rlr1BxRHrS4H+lCSh1Co7IjOPEArNaFP8
IJzrS1fKBgewSaAyYGqElcXPVp8D6ANF4hq04w93eXSOhzNNv5uNCSxpjF0C
H7nYBJZThOy1yxH2b4H7UhoXBoIoInLIZPM45T6jNbvJ4HYbz6QQUjCS8y/b
Nz4mTL0tQjlkDDU++9qd2hgiAr4m84T+8kplSA1kPI7Uk2L3EzZX3DLrlb0A
O06hD1mcCqKil5xY5q3BgF21r/6s/1KVeU+z+vym/f9smXa7jur28fNgv8FT
6VX/ZjL7ETmY4abUvaqoLx5vJkPcmHS0JzoQ0j8bXYoveOOSwkQXcjbMiuH6
NwaJSllICpStHjsHEQTmdBlYrSrGB4ld8Gdc2cSsY54gFu3XXB8YFO4ZnhgA
DGgFfgwCPk5WR8Wgk7r6yeGvki/omEK0j7td5ba2DzUv+QmLwgop9xe/t+ne
r8/mZPAaywzS5mTef6Uw5idlRVzc+Z1/t4fOAQE9FIcxvsiL1nnGVwkoRI/+
ni/CRxKw6ZSKBn6B6mkQBXEuDuCAcHfcFEorCuaguffZMXBotX11N11YY2mi
TTH7XIAxOf322JeCeHQ8TaO998DNwZU4beN+x9Kx+hbscSds1SnNpMg5XwLw
OsAVLUew6ORl5Zc0DsaQOvo9Z023jE7D8+zD0jsHUGo62tKMVF16VhDa3hrh
sHJ3owdNU4bQbcBmVmB9N8mOjirP4WoDIrGtc5j/c44szjFxbu/dasknS7l+
EgczuSm11vV/mz8A4gS+ZfioFqWeszdJQxEEr/KK3Reqc+ioG68JW81iSFsW
J6BhlRLclE1HVH/9rxQyZ2mrvMCX26Tpfm7wl6gbqC/3/rkWwuG0WCXnHAyS
PZJJ5M1LXjV0trfy5hexlSgcrVRFY1xEzVs+TwfzPcCh/kTswqzT2K2uWs3h
BCZD1rWUB9VTwegS4JWCkJ8G4cRIG6/F8Lw0mhcKmnM6lAUzBRXRLAWXC33L
Px+LE/8W+TN/0V4kVKFsklAiK+Zlc3oTFBCNbr9FpCi2XGvpNcUzn6TGn7u+
/jKesHyui5jInmWs5aQuDulG3NeTcbnRcUX6qlPnvVAmp1plHi3p6F9uT+hC
PtvlkYOZFXSkdMl+IHD10paY+oocPEliqWCeDNfy2E+ellMC4xJcUo+Vn1Qo
VnYIqvdRCPwazOS0Z6KgZujVQCUuaqp24Yb+CRU3yeONFpikpkXCtmH2L62X
p4Zn17wbAywsqH69QtX71Ft26eHYuIZVkbp91Di+QctuaVi8BXZ8+m141Ziq
DjXLRWqWhhSPyaWu471pX8V3IajjJLhFdtTkKnYtdIliL2pUyHp7AC8bQBN/
pBkSd+fZihIIDXv9HqLelWhdRzwirbHzgXcXdOuO3v6Odbt/4nVqahWmn+Bp
Y9CsTAteh5RMcO2Dui3iKh93JyfMP4HGHSv+4xr3Mh1VUrZUGM6efm7fJpUR
rkci0vtxDNrgPC6yI9KrzTSZqv97NYFREIsaP1fouB0ncXeBU8tkl9V5d4dv
IMXkJO4TPkIAeuQlVHvOTD2KH281ijbaM5ZyJE01NCLtMcktaITNX8fKKx6S
Yv6HDEQXqeqWs8x1C8s6D2uT98VXpEKTvISBFkiGoeKEYjmZ1hAJREa3rjik
K3MeyO5nUckQ6qa6krBJgoDucJsPzs1jDvLD4JcDLKIoJZGGI40M+0EwBh2a
WwH8QslfqVEm0KtnSXccwM6zoAHwb+8NSDXC8AxbQ+ESinggAzSvXALgxMfS
YqLhv3ODvP9QdBDotyNZr2nevSOiGdS2pH7jwZe4GO7ANjawQHLQYFNMq4eB
Z48AQ6//NgIWeFzNPndd9tvEXbrxGgLsAbu4GFxRkzmLWgARXwTq3UpIyypc
doSCvdvRjxFFK39XyYP/ELS6Qpz7L3HPE0gOLBBdWs9MXjyMLNzl/PL+oKD3
fgvEIzxawKq6113HsMj7dNCf7jXL30MlLrkLxhkel3RWMGJxAtQBO43ZiegC
2c22keSfm5oVj1aBvrg7pfjeiQXLTbwLDd4L89kavVdtGybtyi4hP53EE8RK
+wR1wc/MhL1zENcCmywKjZHLgUZMjNQr/3owrrQgbL2D4lJaaSea6S/6KZSs
Zx0l1VYF6W3xlWCo+TYHKDnM02AsCOtpqmypjoyDAU/Dltf530sMOAiI6icN
IYXGz3SMVgU2Yn7S2RyxyNZSXaigoZsn9LDe8Nk8Lctgu6txpilhE/wtt0kL
qDpiwNEe5HqoX+BrXqh4YUtgsW11Vl3T4OC4lI/jv8DG7WoBSTbF02U+4r6Y
qj0Z8OgEhLB+vxBVnjTB1QtcLg8dQEjngrxmXvv/FsM5t9YF8jlgw3v8yYy6
LGGqRBMUzKyxYa4ohq8au3LChH7albBIAVloY8hwodQzWh4q4vtOui+sVuxB
sowVt4zttOsqiPoum+Diy9SCYSqnPfRPeiwo9E25kpnJK3ZGVoa5vMrQlwuh
dGMm6OHmhqa69XGWX/mphaNu43IXJzSEekQ8HZDUgb4goi7WvTuO0zlupzrK
gDZJ5a6/93HVjV+nhvQ1z9YfPozw85EQwFiJaa5dUbJimn80

`pragma protect end_protected
