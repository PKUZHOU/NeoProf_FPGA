// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
GiDWsfPnfJYZqYjPlwhrCP8PoEUcd8XsCqNGCXuexJT1M9kFc7iScuGBabLJ
Bg4tdAksZypxzQbqCqhV6Smak7eJC41Y3cnCtXw5GerOY9d7buS/koGz2JTr
w0A0gnKlGjYbqL+Apb1wp3CiwdUUglDcScMGAUypd6iATAdzAxYtdEDIOX/F
EnbweW6Gnx0MVRszo+Kkm3Ej8nVei2UZ29qbPcHQNkkUNQzjSNLp6VuBYeP7
0iNL8Fjq2XGDgIgrvqHk7R35Q/jH1G7N8KsWbyV0J4gYHL+ZAJE9m93Dqw6W
7pgspIUbRnVG6H2dLJkQge9WjnxVYjVcpb9ZklJ5/Q==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
kNndIDvpMTszItblgKvCJdkS3kZV+qOPQCAncMjNatby9cw6hwmEPX6CbDEC
cl3s+q8mKdNKzCb5ihK3fVxIzh7kZ3K25kOSbPHsouV6w1Q//rtgB/Sic1+K
DK5E8yW8GtVTTkYo2UkPaVhvpRtKvbUjLFf6X/FWO2OLnh1J5N52yJbTUEdl
5K3P1ulNV0qoGVPZLzOLzpMDqpYkglLavlqEOlMregVHJrZHrnItLNa6asoT
8OzqH6gIqdrtaHHhHWz06b4EWJNZpw+hzXEXPcGJZMR76NuMTJeI6WJPJWn3
REq/rqhQ7m7XrUynfYQHW6OwfObQgE8UGYF6U3X8xQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ppkBSubOYsQna/5WUs0B8+qD95fWUIOLGHz17DjtmFnU8DXtq3ukL4bE6rnK
Md0hnywe6eoWoL0x5e02vN6a+RFdVGgEbfF6r1ZdPhoMQlJxpLQ750fTSQR6
aAoJGdegns+9AD59ojjh3Md/DVqlh3XdakbMSBe0Rl6LTJxBuGguzmRa4+KI
DOceKv2HRoAxxGrMpwlXCU+uE5kwrQXCV6GxDIXDsFWVEw8d5Szg+jvT7A9B
wMPfNeNsLO1Nhzu+rcgqrBiKoY2FBklRXS/b3fpwfrnD2xpu2+hfPCrk7f9W
0mvk4VEisREVqVqU1P+TUzp6jW2rLhCPv+Bsy8c4WQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
UWgfUglHHDnVHEiIcriI0+5nx9rfX3nUFJXGqLgBkmnk2RabSB5PjwaPVEKu
/BQVffpn7bFanLYc7dnWTCajttrUkeeKzHescNYxX26T0N6OIWqCCUqRoxQW
mc4S78CaB7ekxvyMogLmXOmEhPi1cKoGF/FCgnSIRWxxBLqPVSo=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
dnIfcgzuXRYPri2Bf+dK+l9AnRMEW+QSEruQgEvuqmv3ccxO1RuUE5wh3SMQ
EOAD10DQIEZmk2d1UD4AfU7+4mvptSjz9idtOS5rLhg4vTlrqKgBQJctD6+T
JIBPspjmNt/WYJ1+UufSP3Cn0b53pM4MvOKPFY/YzQd1RbnubCU0XTzEHlxS
nkMSB76C4n3qDv1kQlRE7aUUF7yXkwQi4Vk5zpxwPgmvObywSfn6OcUQHJfy
WDfd7pQenHqrW3iW5Qe3aNgjfbqovy8OU+sNWASGwcKugHcDSbriSUBNayS2
mbc6nYscJtnyrbwo1ctPGC0DxADEed6pVX0iEj5q55JVXY6XFK/4gRY3ZaCg
NT8A+a3D3nS5UDr4cOlXWmU6lF/X4LgesDULcFmCzUaV191lngYQrZ+vtgi/
fb4CA6WvXctJxe2dQxSqzR0guspClqIZ7HqDIkTpwxmi8TlmY6ZK4Mj028wu
8rZHhNTYSe15nhzeR0nMNSq1vXeW/CU8


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
LYqtkolv3tTU+6zKvPEzx+QEGRTAa2aMlHJ+2UWJe9JWctmgq4WYLXPenTjY
QEFwCsaXl2gwjkbF42r6Zc4Z4ZSKZpkh8Sbc49l+8y4hXgeOuJjI0BRX7PYP
5AvG1w0Qr8r2wuF6fLiWvkMaxy270oPaM/9vlHpb5TOZJ2ToAGI=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Ti7zqIWbmld2h1Te70nDsTB1NM9/PU/yXTu0bdYxdDJtzJT8xyklMVyCv4in
PsMgoLQkuMbsYcxcI0fQ3h5wUQv78ZJpRf+In3kT50Xj1xcE9T9BbL3X/ZSB
7h87zVEEpWE0OgUrCEQ8XYSw8kPtgSVqUIUudd4M/Md2vNdHgOQ=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 3568)
`pragma protect data_block
yESjud1SiBvaSg2ICUlg+YZejQIWguYcOZ+LhumB5rOWwdRncngTXKgGI8gm
crvwzKlSTC6GmLBRMQJYWvOfzWO8DsXzjBysDJfeXf1sKul9u23i0eMbRWUb
IDZZbHwR4i7WhHW2Aw6KKxjsxd3HwE6xSmkIkZHy5pszSvxQMUQYKbOeZzme
yNrjTyBkqejCQz/5Jve2DJvxUVvU4G4zq1rJ7sKYYZ6cHPUgrXBLAkSFIr2N
yG+hX6BVBzOqjzkfohe5FeBNPYuAOVSOcswarRCx0BBHisOuoIAU4vql+FFW
0ocC2ezOW6SkcMQSK044h8RL2Pd1f8AkRZaiGCunCXAUQ252F8rE987UAmll
SQROR4v/AmHSJGUze/qwQT1Y+N+wWl9ioYqtQYtvGu+Jx+RPFgNmd0BLGBMP
kcyJ0z8nHLCNjvOEafjYKdiYsTqdG595u9nVHEHaJtjIuvh4nohtxGr2XOP9
Noyhth8fnxmmCBHga0VrUh+US2hyyoYId2pwFhqmXCCcRf8ljkrP3KSuFeDV
AOyAlc/LG8/Qr6Xu4l+axJxLon1Cr+M7y26TG6giq8SayQ065ZgVPlkc3X2Q
jSGQHCoW5EL/VOmzKr569zzfwQ3d34Jssv/mbjl+dHQzWB6YIN3iG0sDDwGF
8m4FM4Ju7/0JA5e2KdBxL7or1k+uqsCAx6Ql0FSI+aaGpVgjpTKz2fXBurZk
wHFTD0ol/gxEUnhzlW7U7NbwHvVI+5CUVcc3J8mhHDuUYJAJi1jVWvHgK7Nk
OfWYRxz54blmk87PBNwp5xUBQoNXIXynSbJiyUmucEVEBes3qBJLrrZHMvvL
AizdGWB3GCJlpqJ2Vxcz5N+CScbHgJA4KR8qZr9pZ4SH5xytgkHHiOUAW2q0
62T24+z443EQuEmILEKT0URwcXOJhXsi7u6/Umv4zrGZNLTnS23QChxiICPK
LpVi89x5pOnWMxvOq7XplX6LadEEqy0RzW4PRMhvwbqx9nd3oMHo+rGU/Fcu
N5m8BJom2yyQZJKeCMhbBZya1Ajw4Op4ySamU+4e8xLbf/H/vGsJvI+G2N7D
jymqWacvnQCT8PJfa/Vr7eZ8srvXZnTcc6n52y5RLzzh0sTl+dfu/jA8iKEG
mPGZk3hzY962ymaWr9cBJT9F3e78pPTg9RTJtaO7AvZvAtOYRkVXtobElQYl
nuOlRBwzI21lL2ZyHl6sl20EIMxddnx1pCf5/lUiV21OF/Y/zmFeK+UynWfu
U8qYwwSfv66Wl9HvIJGXrUq6iZ162C7ug8ZAOsD9LeN3VI5GfuXlwu0VA0nI
WWvSYL7U0hEjnwbQhOBF2rGGy+LKI+elE6m09bUaybdqDjSLdlZdAXscqd9t
l57np15HVGcAHyom6Rn8/CcjU/Zx8ohqZQ/Q7TZWsmiPSQ50Wh4FxOVaqsXn
x67S4aP4MS+Y6ZH9ZlhCz5Ey2LoeDxc+DffOSeA6iFDdUh61SeU9zH/y9w2z
/BwbRr0LdpCK9F0+kGyS7bDRZ069p59+vtIZVeTs0Dk+y5mGMd6xR+QRmnFo
WADzaUk2vj1QjnfsmyX18VDRSCgCfSl27YQT8Irg396RBhO1aWzho9xz0oyC
8aq9cH7O+85rqylDW6tBNolCADp588lvq+9uvsyLsnqmhpQrvVmV+QnxwpFt
cHkm2frkdrtsQO+tRBu1dz3L+xtWv7f0rR38GVF+66ClYDX7Du6/lmrX53Um
L+hrbUdmcRRJadjwVq6SW2xmGdazOemkCLuzuCx7/t2nvC4YKTjtgBgFkDPn
3DLYgQEPDoPmfyJQ4VtGXgd6Sikeol0Isp5JqPS5wHj6Sd/udLXP72S3MlNC
BtBd2+rYZ8gnkVZGGLeotSRCQjh57YCVOn3l82Eh/RNMX/MQ4uTYwl2DA+1o
dZc53mFaGs1m4R4v5r6ZZKWIjykHeA5LV0bdxbhF8X5+DkFwj05qg8vn8qb+
MaZ/OyzAJfLyw5M3/IMDAN5yZlHgC8Y0HLQYkjvAXS/yVcvpdWskFA6lAXRm
DfYNSXU6sDMrkPoJ44K/Aapn5vo0FOMQdtYjDHXunc8B6CYYJARqywaMu2wj
u9fy3KhJh6tx2Q4cyi8+Mo3zrUY7Y5qdbsySFFx6LzWPwxQnhtmI9dPBA3aV
xaiG6q8vcqcd6jlB/d4p6qjtnnrjSDQ3oz9J1NNKB+nBdHOEuXsaO5ZdkxNl
vCdeoFMggT96Wdh3YHQvJvl7zq9ulaQgHU5w1pzzi4L+ENuLWiCJ7dN3WrKx
yw9R+pwytgbxbn81MIx7cmihLBOKbP16qIxLxE6kSeM24QqBTU5zNggWWUiK
VkbfzTiMh7v/IThYK2p0LktOOwNDuQgeK7CoaUaNgQ30P4h1VR2CZAJgUf0R
REzPqzE6CWPiH7oJ3nfabT9iaQTQ1zQTEdr4eJiUYS0RaWRoY0zFHxv6TwbV
gWihpajD9bLjDb23b+DgFIEuxlWvT8ZTiXWOs9Hx/88iQrbaoF4tyVFw5Yj8
lMBdjycHZAAcZNSqzQl9VvRiPUQR3vmMhDTAJpYB76MA66g/szI7hjqkgtxn
YZnI5du4WqpONNxJshm8DMuHGcPi1p83WuRKq8WphV2uPX5s8fcSnZTCCuh7
JG/h+yH7FJ9a7wjPymQn/yjbWld/1uhA6agvyNfP6OxOGeo7Q11mqyjVaMVJ
3eEiYdPRTR6QBTN9u7Tt57eFdLoxf/z6iDqliq3alBfStad1A7/3kg30Ntge
MKvDZUa3wb9v996qlqK0L9mlOkrwmAfVeD7GWJegqIQ1tRIDtw99/iGUSKru
vcng/52xe7MjJwTJfjoTLgT+nTAzoXs9W6R4e/5XEm9p6Q5I5GutHdVogbzl
3KE4CEDfLa0OaT7UjUxEE9ggEq0DqjMIlWpAzmXLeWkvUczz/zNFjLbAqJb6
e0yix6Rszu+zPUR8sdgzFR0YwZ+UAf1+ye8HXikpL39PBRtJTfvvxOvyfpKO
1n+tre/ioyqBdE6R/TmaOOeOzOqOp3Ml7fN/BKJOCSRurTQVv2A5Hp34knps
4ykZk9cvBVZyNEnjGOw1UyS4D4C3L3ZO3CWe0ujwSmrHqMTnvrsgCb2WNEV+
h5Y5oMjYSHov3CKczQzr0RpTcyTf0/QUZkmUSM8nkwa29KZzL/KkeTrE++uB
Fhs8ckov0PR7MizL7O3axlwDSfPRKP+q8Gsewj9pmCL/7jC2zgNy31zLwSjH
/S1wWGsPGO/rntmj72DQ/3s5I7+/g45Kn89CQpBGr6Z3oQIYJimlnzDw3Owj
DD7zn0W8Wd58h2FPZlCh0xgAmdWYbLRAlvLAByxCbosILl/YSiUj2CTqMVVf
5yhE0P7NlX5BkC7SrRvADtciQphmvMDyt05L3AUJcVHoR+XyZtG76xFs+Q6D
6NNhCOZhai+LR+hmDcKUv390B6NaYxFHZ5wjWY/eqJKzt2kn6RNdCI6IiL2O
85exgvY5E5UyOhEWlYoCJvabgTl0DmttRcknVV33k2rQDYhKFhszfg91u+37
2KdK1cSkBwAg5D1LqoyUFo/raTq49xFLVnzlJTRvMNXFnEyw4wlghuQPCvbf
CszIPDQiXbYCzgWVWbhofbMnsXPGdwQiaMmO6RRkKgGhKD8Q0eJJG3Y8MDZg
11aySPWTxScknROKv8xcuVZHqV3XrFWuWZJwgy67tMnCVYLPAhJAU4gofmTs
CO7y2av+qhvzMhFzvoBKO4SHFEVLLuqaL50Gat0RD77NSuqyxxkqn46NkXWs
WuHNGFlC/42Q9AyiCXRYA6OYoasAicqtLVTvM+1LyVsvMrdK7ya1bB8TRNBZ
FBXX/ttJ2EZPAalG8LU7Qdos4M+j7zf08eTGAAE3336mKsM0vh7RIJ+QPq98
Qp8nUvSF4UA5EjmlBRM54P9s2EBtH56HEN3JhENvZj34gupPByQkM9uKAPii
R66AMs8nBmRQ2RIVq+KovC8TElL0ysGOt7HGs8qkedOhoN0k136sO/GKPRWb
gGWSmN8pZhLWz4rh2VDRFRa1gfok4gGAyBZz79Ju+o6a4kD/0v0m3ZFcFpTx
DQGq2rfjbt8CNmNRIGEEwqRBqblwcZ8UIyB5QlhGIoYqyGusBM0bEXD9YJRv
s+k3Rn1msyq4t2p/0aPoSG4Di4ycccEdPEZaZ4GOuHQT5IWpKdRrTYsPZiJw
XwPdnb3yn68uIfr6ZOEGOkaK04VbyuYCJKtEQ+t1FdJDcjlGmGwqzUWdroiz
aGIjyMiXw0Qn83Fv+uvKrrgxftwDUVMZoxRSZCUwqT3+anASMrYneXNI5M4q
KemSldlRU88rz/5/K5yYzUlmS09CbGpL1vfwR1dYFD9AH93b1r5zlsbtYIO1
pkM3n3/TYf4F/bkvqOF6Od/rOxVR9wcXT6p5fRjY24DNQC/wyGTcbasvCJs9
nmxYucU+4ndenLyQUfKPI/5o6uc6/nqOcZuDprzElRQdXr3NGekpT5dNy5ZO
ICSV5pYEvi+xg+Hz4HnL7YOptWfrr73FH6HKXnkUuNs2ExlhAvYPndyVTkBN
wjGhJRgA803M6XO8r5fzpzimOQsiO/XOYQVKTTtzvD+M602XU5i2h0SRKPhE
5crhYnOa/RfRyK4H4aOylEQZfukXmXSQnJUDsbw2Usi1tYGMgTsGpw2zIAw3
Klo7zZTQ04VHvhTeIFVBmUoLNgbDi2l3LvJUDjl1ZdwRKXSi/n1V+nV+Zn35
zQzRB5/pvwawWXg9Jg==

`pragma protect end_protected
