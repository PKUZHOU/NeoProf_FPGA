// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
CrHVaMgIA1iJC39qDaVga4yCPB+ThgIAXYKzCg9ocO+/qMne0tyU8aGEVdcqhbOH
xD+59uWbDAGzReyfnKiscm3IsaKbP1mOjmo92ThI3Xp6tfcV+0BPN3NOgoDBT8KT
8gW5oY5jTp8yvG1VPhQhyod/BcrZ0sWkjHso+5CT2m0=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 217824 )
`pragma protect data_block
oBUAL59ss0OqOe426gI08E+PV8TxQJQLfnIlkXiIq8Kutqar728HwtFNN/dbArly
VhYEYsdgNEuVdzbkL2ROWKPtrhsTnEEHrVdHZLlnEJnPI1t3mXB7HT+ZSCk4VIMr
GWYVbhRbrahcHK0SjP0y9c9+fpmuJ2CXrTMhiSaWUhVEFrXrWuZkLjf4uKXUJutn
2xlEgcnLPMsoC/VwshfuDzqSf3I6g9RB3k7+oO24HrSuHtEZbH6+/ShTxBtQFinI
FTrqwZ/1XTnQdcIBmJBY7YqXUJ38MiPEKd17PNdbMzIUjAuK+6fzefVyZqCogdxV
vsYzFy6YUrr0uIKQ2ri/pNTau9Q7HmdVuMIBNqREWuO0cr7nmrqch3KmXklihhu1
OQJLgPM+16vLGVzFvmjRXN1xnjItnd0EPlQpOxmWB7gNDQXQYX+DP8clEQ7C2j8j
52lICjXu78DvXiWebL4JcHxz5Rt1TrJKydD8VjOl642Ytmu+fCQuc15nmm+2Qgzz
y5n054LOsebRmXEH7hnG/wBNK0ow5dJtBL0I7D286h6aJ4JzBo3zGH5hVslVuCIx
nmnbnhD1JWLquJexoWNRHeUB5Acn5tv8B9VILk8JBhQlpnsati4UC3du/7fFnH8G
Ce5NGJveXi42PCgMqye2vlki6iVnAgEyU9I7ywQT4sYnMemuntUD+AZZ3HM1klqd
nVTKdFNAQ5uKRTOPDDX2LU5O6b+YEK9YBeeiXyWea89f5UZ6gKFFzyIMOjdA0tco
BmSLAhyPkAQfA9/KoaJQXouhdYE3n5aBYGcekFF5NRWJDTyrfufq3LxHiZ2ewhtE
CRmXdHqL1RJXt5qj39kHdv2spr0SumoLr6fzRFx38md99sVDWj+3FYuWPSIHjgPH
+dyC6aTO2cTR78Jhwwc6TKYb2+k8aWxnLp3I3OMN8LQAyiM4nEkXmHpL3OLrk6h1
F/CluzgKYWz1dX/XoIKlRKE7uqzFNXImssq2UX3d30MD5M6z5MWif5PRqKj7ZB/c
Ynzk3AJjGLYZyosEO71iFVPg8coZ1FYDju7HYtPPMQJeB24r6B8Tcq5JndS7FpMC
Ng4KZelz1Psgpamoq+C43DfFyt2KPtvMadyomJE5k3cXJX8XQxdvBo3P6lRwWxnK
GgzJxTLjmLD3XA7vFnW4EiwGZ+qSwAM+GLI1CmzzdMIegBwG6/6xTbpjlPel4UnK
LH43StMUZdk+md32BK7HSr8aAbdVb1XnvuGYvUiCiAZIkACy8Wc81b6L4Rb73pys
COlnhUyKwnsaP8IIbhg7pzg8YX5yAoOxIZOivKVXZFDN7sUJPuYF83fVBIFr1eDq
dOzb+mhi/Lfj9xkJ7Mldo1hhmsAD54uDQ3+h4yWBl4i1PZIdSVYjouQkvblPXISk
bZLJ6hGO295kvhmtwUQat0YT04qLsHiYyuNMBpgOUgSXsoYRSygPhTHaF3RD0Qhi
UajdC5h7eyMWft1AiTRcgMFodlsRBV/AA81EveexH7JgpChmo8erc9Er7R9QRT6D
UcLsD9vWTMW/w6S2oo1g4vafD/VncRHAi4iR0yQ6PAsPojksi8nAr1CSMhmr2nm6
Kx14RaMY+Kj5l9NkAexA+tekgLd/ME408hlS4w978sUrlullfxW9FhMBhrP2cUAU
p1jyJlK1BAc1wt3Daqb2bSDVSXQZgegIcBq0RXEakiOQHoaQkBRGJB++OUwOYnTm
jznGhdPBz+SXhiPl4FMFYwX2cww84CvsfGMjzQPnjnGxfgGEqtxJ7D4wotRhvcdu
RqPCyTKnmtKOvho+oJPzmuraQITPZ7a4zoopZGufJRqhoUJ1l1dJ1SUzTr6Z65CP
uJYYI2MOOt3wNpQzdwJJb5twRC0a3civcJLMZ9AozyRAaM1n45oHhRfotT85r+N0
cIrDPJKjCpIJyEgRg5zpY/xnfwkZAAGxn9QWbhjxE9RecQtBydSSMWPFFOw/7cOr
n7K6yL7OavbEjeW6b6PBh0EFVAyz/n+yuUm+nlUOL+nLhJttUJ7GbWiPC7tj2gNE
ebHeh0sns4mbO/O6cy6aP3dwxu8SFb909i1Yfq1wxrb03cacjdH3o3hQjDR+6+GW
Pe8cRO6F9k2vZtR/nz+udInwzHXQuS046Pqr0Cwh0u6spIj+CHl47S7ry5fwKaAa
YV+dduCfWvFK3fJIHBjnye18ZsIXs3PN66zjUg65mGny88AzydsengqMk+/MEE1j
nkMgwHBHxoO6k2PvNPP4gnddujZJVEPCXFPaB4h6o93hkz1VZRrVFogkJPCCTIx2
jIUCaF/3mBy9eWok8G8c/FqA/igpw9NkoNqkQACpJ6Oe0DLcye5N1vV8pgq8Wq1D
VNygC3oqt/vn6kQzfWtFXoQyVi15AgQVHM7yX1XGJ9DScgDV39gVcAutbFimUQWy
4hEQMJPxl4Hg63w0KlGRSnwh7EVvjy7rPFwhgKAM7tvz2XAkGDnVPDd3Q7VwhFNr
niIJlINLdrUZlSxCueQWmqiRFCE5KnWq44UetTRx1+kxFslMY6H/gHqG2smvieu0
ARpseF3b79SyVHgyb/rPSxwSMEz+kvK2F2QMOz6c6kLX7N/qG7ijCm8mqbAZQzlD
Qe73dxQnZF1YwdPCv/K8z43Ees+JXra/SLoTZcir/w0AryEMbhkiI+svGo0+WCWA
95B0QX3zdufdp8I7bOHNt3rRpPHQWogmTlr8zLSthvq9o7VRfVLN8YYT+k+ZFv88
9AINdsxbb3bOr7OIE/6Q6HHwgrQ5jdEv0jTdIamGm9+Qs7dKg04F/62G0BQdSplh
nS8UugFwVc+eBrASCaulaFFHicinfl0azNJAv1rNM1UiXa+WEF0fSk2RFYS4n+bc
W3GEd+m0EJp+9tULwhLXmgIR0wf/6uwFr+E+hflyCDHybteR6UhZMluAvgn6wvxi
YqfACp5IPV+153XjK67NpZVuRYaqft/YShdxiOA3+xftv2vR/qBTZs3dO3E8b2EX
YrntBqlrCLnT8Vb5c3z0F0l+3fTsw/E6DjI4k95OtqV9P0Uv/thqQ1CixTQmgo6E
oM6km5uneGsQmxnx8kjYcoX4edLo4WzRlQ2m37Acj3F5YK5NHSrqm1hBBrdjqXYg
7NMEPsLtTcBmp6AxrKl8C9lVfagyHk9g7V+5JjBLSyZUIXnVN/SnJmX+YWNgZh6n
TSusxnHFUJf+m6n0h+NDToHviPS/HPbb97AAbqfBxqEI6NVUyrTgpW2uCOaPXxex
1mQCDcv2yuthzKe1YrKiBaMvseQIbGw1fEHqUU56bNnuyg0kFysEnUXoPSdhV0JT
+cNiCpiRhWbp3zQMpeGfKthoslEYJhNvsAsHEzg1FyEEmExHC7y2DU57T3JI2PXr
g1Mx2gWugATRekdsSsCPRtiCoTKaM4bCXnq+aiYEHTVdZccuXb2UwghEXLUlgT9J
hMPPq5U+ylkhNZDY3Jf2hXQBANd42LU2x/0EGiw5FCo2WwA14Bl34XYO+UpeLioe
At0T9xLEum4t80Ioxh5RSlgjhBfRyO1Je/yLs2VTrVfivV6hHTSwRFYqtBPYVKxZ
xk5n8b9hUnvusIToDOhaOhE4hhofs/uhNctNqGaR5YYBVPs78f0fhgATQ0izqkoM
dKnWRWa5PaUEgR872tvboueWo/X3VpwsnNOC7/mempyxxomBM/ARz5jXdVuUOz1O
380VM5sS15noc0mKxhC0UVNsy3BsyaFE9H9o3aT4LJ5lrfA7bAQKFDtyybHCToT3
hZXFGHuNcY6MYd4QtQkG/HRxFCOalXJ9hanNdw0L9iq5Gf7yGkZc5JIOvss4V859
kjQLT2pBUxsHdoAR6+pEJVbk6eCUm05Y/1e2CYXZpFZeP4H0wEqbF19XR6kBZVhQ
Z+SGAh+vHypF4Pwpv6l9/SCketLC7m4pcQFvlRYRusPWalc5jOay+HYQZv5f1oYt
Ip47ab9SfhyoJiOgLNru0rHO+TjhUeOEv1acuBA/AczN88cThRkgPoWIf4DcHRzK
/+8aYETmeKox2Yxy6S4WjL64bCJBg3FcDx4tJsR0oYH87zDUhLy8k30ooefegr5e
jQ3D9r5+cyo0eDyEtaOeV9vnYq9hRMR9jjEMQUeTTvGaU+hF+ReBxqcSyApZPKqO
GlLJM5HZgDKrK8B9jVj8t5Li6gBl7cUOfryfBmkxTp1LJOvaT7y8wMmz5bVtO+ve
K9CzcB6UxSnm1Cw3u3vB5iq3a/mfjaGUv7l20gRujWiKXV9IG+GYtzpnDA9hsZLy
1daS2mbbEn+/Jg+RB6B2wPPlV1FORqtntJQEl4DDhqMhxZiLpaIoCjP7NTTmbHpk
NwWe/DTSZqr0gDUslnfDTXRxaDiBmanSWcrCP1ZbjvFIyUV2YW6rUJ3T5VkZjBk8
Eo2dBwf3wxFnqFKkR0RGfzZou9GM46Z0uiRlqbJyi7jjLkfh61dvAxOIjP+9a6BM
0yM4tHzdGxLZ6mAecTjzSYNA+GjqEXank1vQSgDIRHOiY6i6jLVHJfJayeGVnWUy
Sm4Zo+5GGDPxD+vdmy+uNIYW2tArVQ/Xmf21H7FXlj+GRf5tJa+uoRGY7/dtkGIQ
GYx9n7CDfaUR8lT1hPyC+BRcp7UtxQJpvJNHvYsLtnzH+X6NK63DAUKKkwy+f6r4
tcF/8TTq1F4bv+HkEr8jsxaxJiFc6XTbR1DTIy7BSjyozXDuf4WfWtH8njgJE6mU
/488i0WADG4KNXSU5DzKR1FiJi7zijmZxC7NaEnDHHE7odkVoinPc9AlH/5BHg1K
wVtRilK4zzqWHFddjhJqk6q++W1RJf83vJtHHH48K3fIcYjV+JW3v2tRbYr00uqf
8jlIecWg//nP47DzA9bw6zV7amfqPK9o1cnMzphvoCE1Md//W+86o+28cOtGYysp
OwqzIfSoRJBTCXxXpB7vHmCK9AWxRYHBwPWnBFUxrVqxqpIF8BGGI9kf/DXACRh4
NbQtFHd3ZESkhZ18WJnft3AdjhuKmYg2NdaFcERAkSMoN/r5PbVi4Gf9Gy/03Mkn
hzA/8fIDPv4jNBctijq3mhsddZLkDrEoENgZOQesbPv2mJ9oWJza9b+ZpvJP2tfm
ZcwZX/31p1eOMsqJm2xio1XAb2JBWFzqOOR9xDUBeuN5xqXZCP7aMTRo0HFBvsVJ
dEvqS9bHrC0uV0Ac6y8YhuEjuz42JjlXOZKj47rW2oJnNslWUly6Ory8tUA8IHDN
IUh5iupN+58WF8sx8Sa1zAbqs55TNBOHUQmYw4CSIOKNg3pDPL7cVD2HF0WwdWTO
MNZGq54pyq1Qf/osOUIc/QnWugE39zmiv8l5lghyILc845mlEjUwVLm7xIbVgOJA
/a0PGNdo2NLu1Mb0cPOw6F/2Lreq6fdvB/KlyT9Ne8YXwPqHXphYnzlS8rNwkxpG
XSkxWL7WatCzULitgz4n051bDHH+MZGQcw5NnR+KA45sKdMaN2ZlaDx2BtyS9Ia+
oeRjlnMo/UdmxJFXsEyMw0QyNg00lTWAhf0hwXWUXsNeIRBwroE+r5WlVteMSqO6
B42oms9GZRIxn5ph1cZTK3klYTGHLVcsCxT1apkVZHcGJrnmJ5Qe+I6HhQwT4ITq
eG1cd9Gn3aolaaTecjTIAw8dH7sYQoglzVncS+3bHG6G8/okv6R3N3m2YnaEAHm9
PHk5oS07ezfBZB8v4X0g0OjflhZa8vh4/cAZLPugCtIu3TSS6JNIs5sf56/sngc1
g3CDnB/YIkFoO1gbalGAD98HEHU3QCCkje/P/GD6fBTx+bpw8qW++8b1aBH/Spo6
/KUZc2sBujTzfDDmVNeBDCvGWzWRaCZjkEVeUT4c2pSg4hyVZi1/Dul3X/EK4Nau
fmOv+7xjQ6MluwYY/7IMDTBUUi7eLdrys1ZQmvYayY5CJVuvRjdqRnu4/K4zVwwe
hh5HcqZBsdL+JzFhXuHhMLl8RcxleKxTP9KBjpKxGkrXrYgrVqR4ZuDRcYhQWyBu
p72QgUO8XRUD2IrOFhJMsUjSi+cFZGF+wZ0jx5C34mFRG5Fl9oP6l7Ibi9vZQRv7
NQlm6Ks+38F6eHKJlXm4NRbc0Lf26MDwXG+gmF1H6vyN+XapCeCcakj03N626YnT
os0lSX06W52CJf/15pWOyXiOdeAstEuoRGg6oHz5XZZGZCnl1brHp4s6dACxVAj0
B4HiqpRi7yfvQkAokQmHSMXP0FTfbZdnAkOg37e2Psfso2MeIVXW50HnIlCoeWbP
bUtHZ2ZFk03SEl6oF5iaX2nt/nw4GLJF1AwmytKXRsfNfE1y3bl77YlZQ+hlra3U
Hsz94/MBeX29SBKocCCAGQj32ZetVwp3zVnleUS1WNsoTjt+SX/2WPWCirBO86K7
qbd21c4Rdwraz5tokG3l0JTRdmykPPe35MktaYMvyNpMWzSwGdEomb+4daFmh7mR
QDaRLSCaqOkL+i3HNVU6m3zVurZmGqmrYQR6nuK8Xy8V1iT0A4EG3T5SjBKIrExX
Wk6LwB1pT5N4wNvXCygDbFY8kUjcIpP+SGgbJD/LTJ0z2/qntTrRBax1KwIEetRy
bjRNTDmydvKn6KVS3ERoZhvKfxYZ4oiSBNDrbTZLZdXd06B6v3C8A6E4awyr0AUL
ZqdeUWgITrChPXOJxS0hAQ4MHXbYIKXb3svoX2YqIYeXUgQqED6F3sE9KQgQXhGU
tU++uIkPEKf/ptH0kDNY7fRaxmnXpW8hWh+QrVEFXMHQqUxnqEv/hOgIeshcnnnO
mQ5r2700OwzkIXk6V4aN0C0yq2b3pcS+aZvfHsawlZJwZYNyePzI5FHxMCAGR/F8
79Ny7wGgLb/mBG8/hIJrcxYPmyWqWQBcPCkTq+/2gQqjt0w3PmgzcYr+kj0aZg/j
BqUvh3etYKVghwojFtqVDspg3QP3id+hWcmVkUzcUVLlxeQbIX5L48F+WLhH98i+
Bi0reyOIUlY2o+oi4f0DZZywAEuPzbdRB7ioPACnLfiysKgtT9jxpxGV12PI6mAy
Zmzt2rI+YUqbKaLa/cbAmESHACheqAlqW8cX2W9Ty6yBe5kr4w8NnMVYuZ9yZeYI
raQhRnBoPhQ+0RM1JX7ePabwRrGIJ5x3/zw8YeQH6sUxFwWC/p3z0/I/pzbk+gWF
OR2yf+NMTaFsncim0nReb0yXKeO9zAWxqyn++waNtNvKrgxatbqoRaPXQRmQU5qw
X4JoLYEUQ3+BIDkz1g6sdaZRqzFdW7GcN39jV68vDSZyhXe2ebGmB+9HdvzvaFWX
u3A9oZCgv5GLkrzxr5RJqXy8DwMRXxWadSZ5wNXVL63Jah+Ro6WwnCGpvq1G/XzD
Q0r9XhBxOCvBFmMJ+DHg7bxQxygDMRCoyfpi6ryoWEOazg9Go3S54b+8eF/ZXvHs
2km8gbayceATBKIitzQLr6cd3mRFR3hDAvP2t3ecd2qLuygaJ1fi8BBLTzxp22xx
d5PjK0F/SOMNSbFkjux0RWD0i6K3pSSuIH5Z5bLBS2KQBYd7yO8T4PhByXnhUUu5
T7y+EZVkF7WzJ5FyM9WsFcE5agAj+0/uW0vWRs7UZe6AZ/VgHIYSmNnHNQhnijWh
cXo3iUMNO2d6zmf9jxnX37tFe6Q8Q7I1eeXTbwSmAt+6A7ipPZTljvkVRQxdhU0R
61/a3AaUmEI61upijzqxDshHA0Y+GE7GSZGHuepZDCkS7Kt9GFtX4xs+EpxOelbU
y5EMEwDbzdHWcySO36KYaV2UxX65asz9qSyzcZuDPcV6mpGql3S/y0wfvbPBgfv6
8HG2+UCIoHDqaDNIgbNhojTnyQ+UY3r0zkDa/9nQnwkQLSLF4XS0WIBhHjV5ItJ/
CEAZzY8sQfWuM8Fi4D/rSh41hUU3Leod9FW5C5+dFxS6CXjPAo4ZXaR934tjz4Sb
U6454h8rs2SrSK/Bzj8SuC9G3qcAarRup1Z1MR5hCuQpb9U3piEOhyavVzaAI43V
4TnWqT1g3YXlS7+bDugEuN3QUPOP0K4OLbDEcXVPVHpjs5IwcvBSBH33Msu/7Rtv
Ge5lHe0KliHnzM13tsGU7QWrnLYFJNp7r/oBkseSrIudojgMspcg1KSIkYTRbvPA
sX2u6W9PoUzrAa7fjvB78dTAD5L6VwAo7VYwk7860qxztC2Zn4TKQOyze59FZ7cp
P0EtWn3tntRsIBfgJFTkc/2WujfwK/ZvpJZ6wRLTBBH6wnMkWPotq544gyMNrWI6
Rs4qHJBnLWgRLQ6VD2TQfe91U3Y+A6E7k3blEIcw+pbUpxjrml3qfoAdSgMWwL/U
/qKFXrfq4lVZjPQX1+9Ncy4GlZlJYalBWroP7Nmkj0hEklH8CmGum0vdoxUkXeSL
/ZiJV4AK8iHFVO+B1w2YeziGnNqKcCf/hEArnBsTkCZFds9rec0jq4p4ETCBiEkI
rk3OWz/Tl7TiSLXqWGJgc8ZMwl8VVHjnAeU2OSKdbpeTeZWFpmun8Z2LcGby3x/E
eDq0vQnIG4iGqEN0YCizRQZy0SsHLOktPK8YBmOqQx/NwBOqs9BGYvbWxZ5v9LGy
6MbjifYu2ohkVlNufxGnulZcWSlSJ5nm6s5yjVUhpPgGz5W9NDKOxsHdJFjqGRVS
3pszz0WboomuG/UwSYK+PbcfZkNnad8rKyXB2lJP6hxOj4prQOYesOo99MCZKJPe
deOFmObJAceTGm2GhUmjO3KNYcGogyOwkSrs2QLWyoXGjbnV8drih1HK/BoAmEpX
b+sPxk0tPSyNqfRmPR/jCTB3ut9AlSuqT9aCbOZfk6vyWSCbXbtmh1sWP4ib2E2n
K1ZAPutCnX5m/xbVUiITCvS40UO0nNhUZtaa6nRi2Am2lobR2jqk0YUdFWgMnCeg
meWmUQpC7ngzQdO8WbdG0RuyNJ74pVYBwGxUm2JD5nHSX/A01SmqcF3OdJWZgyCL
c0930JXJNit4b7uJOP/pAlve4kUG/zNLRVblcYCIiHbYXvd1WdofeayRo/ocbJAW
qPnQ1SWpZO6FDAoqt7qVDHb+T3oDk6Q6zsDSePfY8EwMspycEvSrPU7eYjEYJSJP
Z4X0N1RDiXmhJcLs4CeszPDPlxxBYCZLXHwlbsZh+wGiF+ooNZSnujsELxsQKKtG
qQJKNvw5KIZwxE/8RV+RutMuRuPRPCxqUsAQw3oY9a0o5k9zOBt27X0s8RiR1R0k
ARNKqBn7hW/hADMmF2O2U3HDeofsmliYsnPDWIOylSZJYgXlGNWfNUJjC1eUaKr4
4RT4arc7WnIRlp5+jzAC+fIG6UfzUf/waHV/BCLW9Nbl5FNZz0vrgU6Mvm98NGgq
ayclYqVswQOsQIRxYvA4+1XWJ1fwqNivGLwQ/Pas9sA4hKWS85tWW87kt4T9tRFl
Ya3Lxct487VE5+A4HiIz+Pypw0BHc8w085Q+6eW/Tx4Veeu69L4LS3Uj2BMxLjbu
WeGPG4tXjwSQcqNS8b32g93bZwK0J28eeGalEV+T6M2wpeM10TbHgo0wxbIRSAzg
HoBJVgnLT9JrHH/RoozVBnHxmEy1hIyWsnWzNVWq4bc63PhobHH0jj0ak+rjhDTD
nbf9mkYWV+ffJ5gZV1JEn1aOpvRc1P2X1Sbx3/dDB3UGrjV0zhqC7PoJYYKPWiR3
S2F0rwymeGHLL3BxQJmUuiwUTRrxtGm4JSLi0fRSDJO8uAqKUBpBb30F08eOORxR
7Nr73t/fqwzGvjfuJXDaS4G7y0UTLNUhETngaaHQhHQcWO+Xyko6GV4rlBPQABdv
RKvj24Tl83SkcjfKsR6Cupt1yl6CzqlZYERiVY3UfKiebk7lnqlbaMOf6eLY+Vc6
pFflLFfrq0GG7GJxeLmBXE/nh6IcWirJHhiVmI20EnnlIS35c9WfA3s//h/mjwz9
H22yWAW9fUdRqGAL3Fwnx06Y+BUKYTAH4MEEsoJBto5/WLz/6TaA6jWsIyLmsQ3S
dw2PT7qxET6GmF6tfuv5DDieTFTnqNvxPQsb35vRtF2/AFEWT7cg+bdSTcNtPCAJ
hIE0x7ngjwjHw25O6ddHptIHMbweLt7ms562GPLHPLfHEHvtGpmFZrKmRRsMmcG6
LGCEQJ/fWoZIj46tmWjMH+8DR02MTj21h0j6p9JF912tbWsyy2aJobOauYrpbsH/
/vF8fRIV0Xn9QjssDtW5iCPhp5Gz4FTAeL2/8xOzGHegm780IJJ7ALH8nEKB96/h
62Na6c64qAg4Z8iD4BgHIFclIL6JMFHvtc//o++8s43+1gVWikxaJqPYA5/zX532
peno4qBB2oiYUxO7l9xGJypwlQnhuJ4kcPYJvvC3GtSMy7J8DezDlu2SCKy60RyK
RfS5Hvus418HsQZsPny9jckAcfrZSh4tY2dVrvIew+OnwyLUEvCrKa0mkzOYfQAI
MvvdvWwyEGsmMWRLWMhC7O7nSD+EVgPdfIm34qGUWZ2en/3j2n9zDzc94QzX7fIR
SYj9p05Eci94uKz/KZJcW/x4Gw5AoJKq90HEvLbzt3y/HQ+erCsDVBg2/lAAyRUh
CnWZG19wk/kK1HFthOa2sEVdmw5it8b9H8AMR3Ed+ZFY4OZyHKUNDL4FtAvxdSWf
7cTKHFDtQ5dVY9elSenQWsrnaaQVH3HhVpXnQvV3WqB3Nxf9+aHSb1981c0Sibdw
OcQRNWtyViKHxf5E12hevNHdG95za72WHftd7be5DgNyNeCA+L2VHOpWQCBZtEDE
SgM0DYSKM3m9mP8F0TRnIO/f082NZFmaMVquaxGr+W5YdnBzNTD4QMhQxru44YL3
3NcrR2BVb/R3UkY3ywIxaIItjasvlItYW+S5U6ItoPF37bHhjIKyCV4mbJQjFGT2
w1unysOjncMrRrT4TPNOX4UC/9huplotUVIVvvxCvTC8u0CIE/KFII5nvAhMS3Ft
NEyCjfIo3g4+OrTR0e5Yqo2cMAnORvfrHimGhT82XGK490VMmy9BV6gzrmQM5Cn0
W81dmWlq+m79mP1yG+slJJFm2+gscWXLgyPp7r6+thGe5YNSJKYr1Gn4L0XB0Fe3
k0PtyBWNIdg5g8ywldT7RPwslkaibiPNh9dNkdVL1+j9aWdYtPJZMlH3PSpSbn2C
T3b4SKZAKwGhUykIn0atPNtsZvU8fDuhg0A6NbzMe2a6A+oSIouXchKlpikAQRuf
Ybxj4sHIsIOSjN4UPnXDLrrhQOm6LpcCfc3d0H423XjffKd7WiQfvs4hAYhtJ2LK
K7qNrc94iN1t5iU1J9iNdvU2GliMLH31FpwaaLXeUr0YaKsosfHu7KLlnR//x4ec
OGSGvNScHGEa+I95SPuXSCe/scczNKxHxygy6SbgEYbJ26HNwkAka/lVvFvSofUX
s+Hbr0Ucs7RlUV3tPH3nrDMJVWUkrKwOYRwM62hCgaCVu9FC6zzFgH6cD7sQmif/
k/C4aG8RVPBMZkL2LmcAPMMVmqlWnbWaix/tuEmr/tdmJep7jbNhzjQTVBQVui6b
h8E1gJJv7EIEetAwdwcuZd6BQsw81155tX38E++I+Zg62rYeEaGAX17MFc/Qx4ha
DyMGtezNJ1UYqxaid5h6a2/ETeqxaG9k6daEMMOthnyplnQXM/iO6XMHZioFmDhO
ddzGwlNSFCWVHs05UnyPRj4/nv2Ib592WyGIU7FRMcBpMzGFtFdSvKhmRx4NLli1
1GrNNF68W+vIE+l6YVaysvljdL24/f6L02QXoKzyZMV2bhtHFmanjLJ/+MjRRNID
ldiFZ1g2ZoqkghvCbPCotxduzYZzi20ZuarzPZv909Ir0VsXScTiiQtGHqOT2+hp
yldvQxN/lQoVMWFyuMIn0EZOyYgrP3DMB3pAuJORqEsK8tMTcbc/JJP0+rzLSezu
3L7s+zxljNTIJipDoHk1tFV2bZYr9zY0GSTZhD2M74OOCVnj1Tzc/Khv27D4YLt+
9YJmFyRZc3yJqejg5yBUiYIj43IbgkcKJ0YReMSfemUzgt27c3N6l5eqJdOlkEuD
yh5bxwlpDpcdeZ89Mn1GbH0H1fv74XvcfeyNbcc4XWIkmncN1pM0MK8LbkzxCrcd
S/rz71Z5IU7Dp9b3b7Y/WxPf1HJE+Ck3YX1LVLa0rRMhpXDfRY7P31uSGcONzkVi
Zq2BZkJ77ez3NVsgQ9iKHsiPZsN0sBh7W94I+Fvot+ck2rDxbebqdlyTviKQFdJ6
5HTHMdkXtMINJjQK/3yzUZsoLI2WsVD/BfdzPqNpAgjBF05gpN6/i+9RegDZGc3y
Bq0iZXCJndXTnOenQGlkbQT8b8xbarOwRFUa1FlIN3E/begShLsrc6rsLg27jp19
LlHtCqqiqEXeM9blM7InSRYRIyBRgmS0MkTu7syK3dW4j2eAwKuDcjrRGUV13e7g
WSfOxbp3ukuLyohLuaIjYOpguc9Yy/HFrmevOQrVhlG/gRcK56FGmItAjIPRTIvk
5rt/A2PbmPHJA8UkCvqxahPMzReExJdChnkmO0/dT2YA/2p5m8h98XjSyCH0Bl56
9qnYyXx2ZmjhTsbeahNPNDw55v94gFyDU3hbA9VPQCMaI1Fy6tV9w1WU/NVjS52g
Q/kR/foxBTyXHiPlsWis+atq9GyjFSzHID1+Nof/mEOA0jWQgW9IKtNITkclelao
W8QMsUBbddl+ZMLXOquUgr13wdyiYn3msBxesBBHyUbFOBJdW1QH3OlkPmwpLwDS
O5rqeL9mJyoCQoQxRgrk2+jEarFY30C8MQ0zOj9u9TpEz9f/zTXASXjv+UNeROoe
eFgEi+vCfr5iBXR8SFEUsD5u+nVbVhqXV2EMuKbtWAyAfPbJjmzyyUadFZcvZhvc
l0515XVMYxz5eK/n7RSacl2cEkb0VPmfObl4RqUtxFTs2+VTr2di7wVU0ac1fxyd
zm5mKDjOCKn4+1Rb1jaN2h1ST+TFv/jW8OAXqC3nMPschp5bBe749JdXHrqAPSKk
biv2th+pUq5cI+9QKA3/31GYIiNbsuvzjiORO+7ymtQucTdk/O8waug8B38hVKaQ
Q5OcD5zmR+vnsCdHT08ORw2ymRvZlBBCIDinQUTxu3lCQ33a8lFTBEJ9PTN4exFK
Hx5M+TlVABrf1SwJA5ViTersvlnLMocS8HFfkCU8vGCLa0yddFin6nPMnUzE7/VV
CSJ5tWx5HkQrLEFK/OmyV5Z7KhhziqVy4P7Txz9AqVxU09qYLPz1+psZmctXL4ku
ZCqWmqQWi8xRfgIyPL+AtEweAOTFgpRLSn+9uIJGaABDduq16DKodJhIABLJKNi4
KEIIWpFFA/RHUBVijn5TEOZDxgKMctNXzIdvU2D6xnR4qqWYNGTxaHCrANG5ZbhS
FzgUIyOVh0Rb55jTabLrfHH4Vjq3p0htOF7rNZi+7IqU/8vMcn4dQUMufCif81gk
t6QdJafUeNZLnfwiA0kn92Cdcz+uOuvl5mbcXz3Vr3DuZBYBYEYJCGoL6el2S8ib
1/q4xgliBcyAp9RDVHiWU1syHMuWE2FZxU2Q3Vg1bOKK6c4nKgQtluuoBATEqv2L
AmOdVHxZr0Oa4lYA81aE7pdW6/2Djq9A0nDYFZucAZTshnBvU79iY/HzHNCc5w2Q
aFuCI40v2j0uwh6z4S4kFuYlUg7nmcWZA0aNBfG1v8kvlNlnrzXBq8AcfI7oKg+0
96YEFvMCk3BxbBSTMHhPAboXDfL5LCCThJ3RefkGW7q6EsAqEYEqzigeq9FUs9T/
sGjz9WpZi2rWR45ap48loAUIUTG7uun7Dzm2wY6UEtiph6LsLgGwOUIbeKsJ+yiz
u76tenEKSQbE971sloE3Fx3z8mxaFJKMlr+D3cji5Opjl3sIOoCca+IvPypgGd1F
8wZ/lwQz1NRfD3rjYVYCUsTtnGT5bW869QNcOxz4cgzXF+wrVoYQIG4ugsXHsiuV
RKc/y3JYwRrAyBOHLo/hY8wSVbPp4gaoU4YxBviGTXgwTQWdWyaZqmDw0QOZYLfj
RGw0HDDHgGEOywWuMQCVoqubHt29/HOO3fd5lIpR4dc/aiA8km8em5VRMjhGlzwJ
7RB4p4cy5sbhDgShGS5w6zmWdo7zZNLdQcljud58UdykJ2KIi8P+7HHTZVU+QwaT
1kI/EJRJ4Tpd5Qoi7nNGhOBn1hn6XmATbUwSvIWbRsfoe5nywrwzVcXdIALyj7h4
zYMTbaQ8Kl1lX+kBA0gRuQuQHbJ2vZb6pq0xaCcKaMxEr96UdDQphCHxiqi0K6rY
Qf+JVr9HO5cHhvbDHOvf/aOGr8xEfQcSgJU2jIRELmGikH/96BFsVZch/1ycno3L
9pTeVqyJbOYQeLn/d37u4nLDO2YjMDy3wQoHgwkup3UGSVNRHkqAUMcwEGxlxdnQ
FtfdM/e+/pf0H+9j9AOFfE9AhyAChqQl6L0mEF5cHTVg/F7F9b3u1HfnBgXJ0J1s
No7drS80WASAbqkGT4vA/rqJ1DuvEHNzc/4wAQlsUA8hCXd+yn25z4X+6H5zML3A
G6XauidPsSyt84pP7nc/AtqjIWqZJ2/OMLTA+Igz1zkroN+09wvDHdEMcvxm7+hv
GvN/BheQp3wRvCEUkrhU4iw/Sicd+3WDlZUWigIZEMn4GavqtM1WohMGi8ijLDd9
o4i0VO28vGZe6ghHV6JrTwgV/Ex6iRfVm2kh54FpHFCmbqc9Ro558AQZeonk5o/w
Gw1ERPGSre79HkyTwJo35elJpru9hwSWsASnCGTJM++hZ9NG6cMF2HT8GNMwkuko
uPB1C/iu4oFGyAJo+1nExs9Y1EH5YO46m+BMq9W8AUfFV3Yu/YGJJDy6nCE5MOTu
IlWUFuxyHZLAJn3UrLYyxg/gHJRCEWRKIHacx3aWBtYjH8rHXvoNLZiZNCfOyQWZ
z0YUXVhcpyXdJcI9KkHc6XTlYctEdldIkOg4MFriv8V0G4hI+WnWjJeAlEt4QQK3
MgcY+BAZ8Uo1lqCk1GjC3DtW94SCHxD1G3M191eO96vPr/uHU6/xffrH/ucmo4vj
G3W6kgzoZMGNDy85rLk/enx3dDqmGs4wfAkf6zQ48Wb2mu3iYQj9bvh0qHz2UGhF
G/uBKlnNyaiz4LNm+FswoX/fq3w5V217qhYAGH2dGaqn9gPsZxiUO3PE+BwNF7Fc
DFDXU1EdLlkHDqXC13ht8UCwgZ4SrPloRTAMi3+Z+JvzJBj/wVm5Og/fbjb8+PTa
nrRw1dEpXiGpNOvbBoNbHtu1RzXwx8lQGkcJ6cCv3Xnm8vJ67AvL0eHiNkKe7wAF
SlFSICxkKo/Zl+YQ7/cUOqUgHePUQJEOWHpcOdQK6k+xwQs1ZJVwumLpptPXLTAm
KmCLyPQvx33sHbnvJbLYBQvoRY90p78IboA+7wiIzYw4vTQjvhcyHOc6rL9zeVK6
YM5Z4v9312wTOZ86SzpRIQ3EVF1GoKJj6oEZEuEdosaYmy3S+gtkg1ro6mufblpT
DLCUEr1P4idUGWjKUDv2cz4edJfdATmJTCMP2K9qcG4X/Xt1ME93FhnWfFJ76IrF
K9XBp2U9YPStZKDartEYAo3OTG7WGLPZzITcZd2qyczPdLnJzQvQrYacPeLCGpkC
enIbBOSDYChDd1KzFOaxp6378DaPLVR9DrUjx4nA6KU8eyFK4wdC6QPD7qXG4lfq
CFbpMmFj92R/DyaETmZ075OqBBEewK7Cvo0hhoD0UZaKEoyqAPi+87jDtaCsZg2k
c8/5lqnYQawn198Qn6GgXJs7h0WC0r+XFo+omWNoMsleHU3scVT6Ge5zXvlGdGt2
OUF1d5CvSkchJmmlGs6YmR8aMrR9E+1nsunGTmk7vtkJTqtwMu+ZK+vSgGYNuk5o
eIzQQq+0Hkp4myIrV7+flii5NQZ3NqHsNrzl6BuvZO9VeSeIb5qpUJ80K8a3DQyX
Xe7xKZNfbymBgC2cyTM9u6IT90m1exJtR40PESyDY6ZFWiLjxHWZFNhGoz09ajOm
XmwIKYDWbsScgcnqn6j0eoVe02jFo89EqiTZGZta2VQe7QGNP+FenSOraNOIISHP
qMP50bRu7fUGfoGXpCxn9tztfZ06qUE7Qyi2SOXmd//5E55tEA8fTe1yxDpH2jvo
n4kmvQbRelqc3wOO81v7WCKf89XoAzHzJDWV9M9nDJRkxJCIUA0uOIdgAt+KSNDt
nZ3gPAvmIm18P4L5he5s6MZteyfSDRHeXhjqkkZ7r7uopudfYUInYJfe8ivjvmJ0
+eBbcPxhlvtdO/u36z5lwKRK1AFpKUiIy97490t5AT/VTLTB9fvfTet+uvbSSyhm
wIr+3mLFeCd/GInh4I1S6FEsoxwI6igiPV0NjOLb6V//qHsq4EBPZXNQARUv1oi3
7m65ZvETWgBgLB57NkrBbCq6ec22AoAgodZ8EtzS6NfiM1bV/1OUZnbuAEMdynae
HJU6sFySTSkgft1YfMP2tjQaynvdwCVuL9iUwGNZYRAGzZmyNurkgBMLcGLqQjQE
dTTObVNZ+1Sciy0R6f3Z2wIxHx51uEkdx9RPsQH0UsZAdgBTf1tQn55UD4FdpKSz
3vpOTyIanykk6gmyB+7VimzleBdJMeordNu6FFTW+EZa9UD15/AGTspeIXmyJvCf
dbNbdCV7qB7hF7Mw6EN32XRYReUHYYKnwONYqiE0Z9YnpjhuhKYmBzStm/vvzbgx
rr89AVwrsil1WqIm2iC2SZDQ2TMhhZJgYgzWGPUF8fktuAAspTsMR+xkfeFXDc4k
vm9+ncNApBm/Aln9R0K4XH925Ubb7NSAy1ewWtfo4faIgbSI88U69ncRxUoxI1/I
wyuInultjBz/2Rk4fQGsWRMEYtxinOEjlwN345xbpbAU2mYCNuTxBiGP1U3ehh41
gDok8E+P815cFIGU0HiLTowe7pBoo6EqvyN5RIy/Y4KrVwm7JqMg6BvbkOjt95Go
bSElAmxPOqeKFXu6tKYCS9bA22sy7zToCsJc3veWddCwdFLBbWYCclsKSTvn4WPV
AwD1WCI0K0IezqGjoanOkECPgPykqTb3eN5llFpfXQHi8Xy9uxydCq2LYwI1HvMK
MttI0HNIKbxIJb6n1OYXc4gUKsBIdiscU4sz/m585pQSP7GCVxRNgX9En3BSCPIv
cC/KYgZyhAffQjREXzp2PDSZVCIq6ZM19nPH8LEE3aG6SPC66iMBb7jQbNsn4wU/
CHwYWe/IFLC9nAYGv6uJHPxEFINTwtL8wJl5aT8+FRMmZLmoVMAViqA/fl+BDYOR
ZxPRpwU1NTFmQB9GvvufijrDR8OpTPTEjFFWjPno7cIInw6grbkeM+QtFjoa1f0I
cVPegQobCuHZC92x/99yRchdECRDgRAtelw5ZOP3k2Uwd1YGTUyEFs5ue+3nshN9
n7crahy0nYXJ3g3LPZMNhpqK9binUyTqB+/KNamFXmoQtYX201CXI4A72/OxNVr5
2RSix0ipr0hQQz0dM9wYHM0/+G0TDOhiXHAFLp9nJggHehWhbwGxBQeJCJr+cxUs
NctmFpMIinz3vm542hiDEuCX4bZ32BQ6eitsUGdwn1Od4F1onbjwYSSxChaPAybr
Xt7W3RQ/kED2iXbH/ezPlJzsW2dlPHMr1HgrVn1OdgWIkqbCdLHbp6+3PTjy6bEW
t+jvzLqD9RYxMfHPlblZ/me8Ac+iJrYPHciVz+vjdk54SSsxHmOCH9kmzM00rO4S
qTuRjklI5Zte0AdWk7/ag9zHvQ9IrU4rRo8hiGQX5tA6wPL0mJETu7BZwQ3c/enE
vQBVSjq16jvlmjaG49qOlrWwxXqbqwZje7WDlc9YOmv2Xvtp1oiQ8lJIgvSUUO+3
AphXs3l4FrrPdpyuQd+63vQvwc8V7cqfLd2Jp5NhTOHlQ5mX1npFeZQZcWyeJNgv
GuMlk8xwrXJFKxgxJpIvJY4H+LV6zOK0asZNYcFjPLhHzlfMFxYQDGd24Pjyg6mp
+l1rgr0bCe+VyFW3CNe4NR4+hTvx/dhhEmJ4GGEcaP2gFokUR5lKXYA/hwIXUxF2
jj6VnSuxcY7RXyn41pe7+Z/IMJbHpufFMh1NjTxV+VPg8OM/4ovcccGxVkn5578s
qHdUHr4YqMMCA2bXVMfXfR2N5QVsR6BYUXrFClS8pZr53DR5xiRfJu92Pi8uhfKl
5/OnLtVZ3BHiadRnhANXefSe5gz1CbRzJFEKIlRllBv4MXfMK04d31J7i9DQelas
Pz8PT8LjFePKBUwekXWsA2cBtlnT6hjn80JJSfg9kfVdHA4W0fiV5cpcFWcgvQaq
WkvummMWeNe2DsTdbdxC33/BHSE7HdIWSsKitiChW/Q4ppJrKoZnvdjokSpJ9AMi
ki2u5SoZJb10N4diMfGxwj6R15x4wOfCviwRS0wmZm24487nQozUpgkpysMP28Y9
gdGcIX93Z4T3xMivhgA6SkkayEiM2+CKeYs7eX1dc0VyASkDJYT9uATaBP5Bpvi5
EPF4jDDw9jvOenYUmrje9PE03iVD52qY6ostJc9qtWa2XObavraiHtuh2AbGdUxG
5zaReHskZIRNeYvVmRCQuxAnONPwqJWDjwOeQq+pNuBE6JsBDxH05HllqIbguCrx
VHNLLJyy+ZhnJV8sWqxGd002fJKFg31wDCJcgwRsmKAsFoCqIwwTwWSRiNon6ljR
v90USK7nuqzip5pATD2l3Qw3l0w0h7rRgGTWQZvSlFEQWxzGiqYmDHpWAXYgf6gR
n4DWmuqcyOCu7Rtwy+papDsJ9HUzm80J3ZY2MrrHEWhwJ3UoNgAwbGVDu56qjQta
I7maAS353MDwvRTY4t3EXscNK63OxjLASescJLFUnyhvgIxudHGcDShujTLAVjwn
fIevdDzSqB2BrmbPKykjQ2ggCApIHxWJr2KjDewp2DNfPVdDU9/pX5gLN6oAKA2p
cD1UGzbLuTLBJE30euLue/wV6PFoD85vRS0eD7VPzmibtOHYCxnvcDgZj0obyzYQ
Ka3uoZekj6xy/zcwgAEZvk70WOwNkbbCeZRuNQVgkzoLfhH3jxi63tKzMaxYuMkN
RfmlMhnQZkXMfedvBaomRY3mHzLajK2XRcvauA2TfcCkMzUad+AjyejaNYPerxEe
U1ADQhXm11JHqLZtg0UIge98RUY0P0pb8ApgRvOnA2lpNha2eqUrQtja5dd3P59F
oimLD+RBvYgH2emKlz4xNcnX4Z58HDh8/kxn6vajud+1f6Gxd+fiHyNp3dIporjK
eIwCirtRvdsN3vyoE7OdCRvZjLMk/Cg50MNuvcHJc4WSDEUhaNBf/o7G4BEZgprI
EF5PkBqqJJJKvdpkReU0IxLqw2hGW7/O10tqcSvbGCylAMO/T5vDFdmckYJeG3oW
xsyhmXX0fFctUxkw2LWgtx00EaZuDvHRwOiF6blk507uk2dHq3mlXs2o1He1pvGi
lojdnEtMDTdn8dpbQuPKanhvYSz9/Qym6SY5w26tt4vv4MFuB6iwZjX7b+3OGTFJ
fh/N1Aj6fmDep8y3XlGARbInOTZZyhE/poEMKV/Goi9mFSc+cCpskPe12ZmDgIef
kVRsU3kPpYxJB7UgcU0s3DwmpNjGeyztFWKFH0pjeZFrXrE05J9LbSNte+Tsr6vC
T9rFsjuNpA1SFgouth+7YHgelO9T4t61c95OLR0gjkDSmgxj+pcihBAGoCn6cOy0
6vZdKlhxXgfWsj/yDlXcM3MHjYyHJu0vyEHT6J4WOqX79LBPr4/2Ig8GP6yxK6nQ
KFCtAzUaciDm70ZKT1upvA1HT7K3jGjDRx4/tyc6bJe5gAx3yCDNuljx4zX1+FTN
yFQVKSGL7ndCscun5hcxWdG65A6buDLX3NRksappVLghOkDXRy894E/xdIjX+PxU
PtkmdK/J2ICaEpG1dtMk6TWApnDJNMIJuM1WVdClNV7YuCo9WoMhYfN2r1XMZFWF
BpJovlLDRHZyoB4qHZyKLqgCI/CZzG/mfVi6RGGtUinXeAXuELHg7yfhnYtSiCGt
qmXVUjCzgVwrb6Mq2IS2p/1ziZc7mMG/RHpGfhGFhVu6rTRk84J/fqOGnAxWq2VL
6RW68zKipOS2p2Ofb7oDNWmaT/8OZujQUCziAOodo3qPJScQgTTZg5kP61ZMvQ1n
FfmtFPNCsq1GMRMAHoEAv++6UTQE3yZtRO1IaUzCDB/dx+AnQfxic5m8zQ5RvDsg
LQTjIZXUT5NTEE0lz4t17IIZIfHXyhuatQlsGioqn3RH2Of5cNli6HeuENapZrTQ
P8RGT2nuXvwVJvDK4q36vHQowZdQBzqOeufCeGGK0xjMd1RBjncFjt/qvQw3csTT
P0xIgs1LQs0dUSBOpHwIzdVtgsLMz2uVO6xnaA3eWYebPjU66UEBJgFLjx2xNxNn
HOAz5gYQVbT5r3OZ/6zleQ01CCExoFP87h9sCBqPaUoXFYYQVSoLpw0KnQL25YUc
Z8TWgWn0o9Fwp1+D5LVnovvbMrvqY0+ew5mhXUL2jPodjHk+EK9zCWGAz56t6JPb
qNdL5kilvAPlYEY/QHhS/ZvIT5+opuItcyogd9gBiETHMt5z3J3O25ligUP3gPHA
h8z5h/HC5eK0wiFpoqNTh1t4GdaOj7UISjTePm1TqK+Wyzu8Lq0/RGiXiCe6Hpya
S6IWPL8LkyMFPNf5TRyuomePFKCB+eNRg0qBl4haFy+nT+qGEJpgijwBEvKG+EWQ
N/UNYU0UvfeXE7NKtEWWSqCKcFrc+wevKGnEzmPgi61ZZCz/gj1H8hOscyztEAWo
XoSsbZeI3b4xNxmUilSA8hl/mKX4R/vw0R8YQ7ge9kNXxEThumhDhpeMf+bBGFxd
tnS6ku97iagEYQTAa0oGGkitk8nc6fvEB2oKDg3NWwKL6n2dkcaNMZUFkcAfu2uK
WlPkJdtvOkVKeO0AnHUadkT9bc8hPQvelsDDjsmnUr6+0UxR2+H/9ua5GHwbVGT6
/2FOSfIhGamBTIkYfTmp952PivWoiT/HVuGxm18b/TOIzG2Ot7/YE/0ZqPfigz6F
sTIYkxU2VCPRQUAUGDlBSGb4NCGulMNrKlw6Zr8wmC+QfcpSZOlsNEEhl3Nwpd53
4jQhPZxVLcGvGF0a4ysZHp2dz3u8BRf5C37a7XJoczeiLCEwYgsliXHEdIBCDk97
TE8a/yemclwRntiwpiD8yIBxvQ7yDfSmbOZd9X8ifb22NPzfjxbxVDjIq9AIef4R
xHN0c9ocusjx0NgBBXtHNiJ/+4Jv3rZLeH4OwwfDV+BjXtvFDjYtOp5X86XLthHX
Q6f2XPyxgxgC7XB/raXQdD6S2j954PoefPYn57iibkiMygrYAhkq2pu49Iq3zsU5
jI7KdmvzsvDERUhrKKor1w68SHMeUjiWoG8Mh53lj2okj/JlK43yaG5va34nEyGX
hXbXtSo7XooayLf5e442js8+Rmtn91JC1rz6A2V1+3UgAwqALeiGNEWEWBNFk/cz
WWM5TuJGLpTeE9SK3B9m3kCFa4Weo4U5lv5qESH7G5W+pI0z+8WlxuyN2fBmGv4s
oRaJsRuMTFINTnIpqZEZIWUYlE2ptWFGKPkAT4UpRzOlTgtNnP2UvD/sDmF13CgA
GRbQWaltRdod0KmX0/+DLsHM/ox2BocuenStVqSVF/JjFvN3xrAf4NdIZrPdNyIj
HKkdyeDrtpk6AK2iki3b/953EN+pYDKNeV+rsHvEfInQnliF1JrOA7AkXqmOLw/P
/yCF271Er5UM8Vrars2wXF/lx2jw6rr2ODPTfGDp68eFVPIYXVAJnWFBQCz44u7h
Sn+/x2Is92C6L3CXq5chELTb/lM4RV8mNPXlPPklGiuQhX+4mviPX0oNuUvC4hcg
pXG63bcdB6EorUl7iROKTDK4qPwSzSVc5E9A20ln+uqNL/w5S6aW9bL/MUIzkR6D
VKhjSC/o4A+ohKFoT5pbB5+3dTSP+rof9Cl3PbxK85/99Piyhyxd4n7FYOCzfVOO
YNm2Yj3xl9DqGGZ5AU3CW9x/AvsRvRvv0zsFdGHVawua63IyOfdazt/ahampK28Z
YHy2krnmkvG8/2ffZN1lqb7yxj+QKYlFUhhkvDbPv+yfOSDqrZ2AalDwXSbk0UiZ
XNaSPU2HfmV+mraw79z334hrDZqEoDcVMf9W/CG30dAAU7lj+CDL4XthylMv2Jqb
5XNRbKgbmiLjFUIqtmXpKvdyWL9CKkZRo0+usp1yOl498FoZEmnXer1tXwXUWrRT
BKngZ4nxzNaCYyms5b9k+8LyJO2HvgBvsi74tZ57iKNR+wEzjHn+EgJHrKKk313Z
JpzLXJqT0qEV2HjbGcOvKEkyq+iv1Php/iwchllMw/XkPqNZeczz2RFwo5Dzg8K0
itVtW0h7eEy5nhVPnmNaz9ZZF3KPBgOOvy8W65V/kwpYVimH+cqlxcIrd4vtUCRw
p5pJhGMfVUqqdaW2C7nOFvt0padLu3ghMRArjUoSz0i3BzVkGv26pqxaW9wvRUaE
R6e95DuoaHV7PwJsN3Uoi4Hk0le7ddO6nP+SLQiLJYmcfGOZMY3Do02yg3D11uM+
y3TZ1mCbq/nwsHNrZ15woclbY3n7OjlEB13av9BMV/XfqeZuZlQKgrsHuzqBSvVd
tOCXyXPvZihoz9TIxxskBgA1pt45IiSh9Xt0O5G6gyXQeZq81nLynApB1YZi7zjY
Is6xzuYpLcd8W8Q5LWepiBcOlx4sJHma7fhaAwCWT57xxhq6Z+bg2h4I51L+/uY9
kMjVg3Y0QkD8aWP55mhiBh6atMPNjlQe9sv4Ht5Lf5oxSIu6T/abEqT8piZC4rNr
FLoDYLdcB6jCzsqE7Q5f7kWhCE28bzuICklpHfW//jYOBAtbdYgj6N5tCdK83Uya
wWm4QR7XRbbtApbqDpfSbxDCdXpLdIRsVPzyrfJF0roAScs+d4zpL19ODkfWV+x0
kSL2I+UrMOPj19mSsBrG04kyaFiwPNeuLB3mWZ02fQk9GSIRgp8toWGKiUHFICwZ
swkE+CUyTZpz4smRgCYUlubo8jK8fgqPPLY1huCz6RLBDdUgePeqVmDnkV7iKwyZ
wvzQ0IsdX1QItmAsDXkTOmDd/bdibMpt9ByH0WOnCXTZLhM89CBbHnE22TvcdIXO
tpDajGEJdaNR9+Hyfv9sMGBfBw88Mu0V7d6MHMgbNtaG9F9ThbkF5T5Sp83SAoSR
uZ/AqBL2lhf53NbAFglbMreaZ1yvfeJ2FXn223hMO8s6/hpZninbaDAN5sji0FDB
q4HPXFCvIW0XscjT47qsrLarMgHN3o1h2Ybx1UWc+BeGw/4qqdPFxgh0D97FZ6n2
Zkikl4FUvL90dBphiuMq67YZt6SYHV9stH7RjYjrZeR5izN1WMUBNkhsTsTarEZD
TI+pKWPtgr4kIfQYqNTy/jz66DAnDvlNFdk7Ojy0SiK9MZCjllA2/NEtGVV6GNTx
j3lZAr9exyR1ATXdNe8r86ug7tvKuja0BDdxS/7/HMmoB2FrWIpBHrLGSiys9Z5/
nzU7ViVT+a/CNMq8+/Jdn4qgykBf295xJo9JcMfRXTHn1X/HI+sNq0lqCFfoP4Wb
aPQMiDduNJg7h690J/H1SuGf8CvteflJ/rHqlAcJDZIVMchPmlTHLrUpaOsCpBsO
DqHENDPUYHX3BHzaW4y2QuOgfHKd70eMhG/Uf1ejiNGMgDlDzEgbjZpfcMWwWFeA
aTZ4YecSvG47dtO5OBGQT7Kn1GtPcGwNTeHr9JL9NOw+NiE2ONbXTd5WCM+5EwUs
l9NghTE6lyxKCzRaGdAtGdWYGsoBFyJ0noqWx8d0859MRrKB8F6s72yj6w1hObhB
8y+zW9yQtfykKyFCvkUqcRYF1cUy6Gpcf3WpFzVwjObBe6gtzYhhGrMMxmQ1nYNM
F2iw5jnngLTJXBZY0ogIwnKRh8Ybtoho3UqWPcCM9zk2h9RCklPnLEyh3ty5H0Mg
lrMFfPuxDNyPIU09Ad3K6Fv/ZwPpnyRtvvMujf2B82NfT+FGDGRyLdp+vQS6dlJ4
t8jTcTsiHD3cjnDHC6DhVBAO6owgtJ8du+OoKYSwapehMEZDot5zDL4w8wMTsNFj
GZG/yCsJBfreOOMdMUavElsXlagGrmBzIEiPC0ETvQs1etmu0+ZBOc3qv0BKuyts
Z+i0VcJuB3niGWoPawFcs4d8kvFcrxf0dq6rkuYheFE4Q6483QHTGdKFk7voX8qZ
nYiqXLRCNMcUT4RYHKEYsM0LRD13W9OhMXxRUsa0bAlEICa4ofaV7k3c0ZXPawnx
bi/hCwziBF0dc1cwhjmcoR2X/fO2EueyNKOiY2PRKAwR1N6ZWgv2d95zdZyrqMY8
C59aw4yrTgya2XJlH08g7QPgFUxZfIYzEw19tskW4Cf8i26aj6Y7fv3m3gqgg4Tw
ng+RhhYS/iPHnlYwKP+iMg6yGDzDpoI9GPIPA7w09XgvV7d8g1XY8CCXUd7trDD5
+RVR0gN8Cwsb4MAxNmidYdJV7EhPFYP3Cbee05lHanb35IMB81WZ1Sjx9NFFmvlZ
BLodWrZugEVXW2DwPK2m+33OaGvoZNPEeOgZZSkIbNjF0ql/OGpvRbGL3UzDaABK
tlZWhecrrNzworJdGtAqfZ9ZYyLOdVy7wGiZx9ElChHa/5dtOSXC19bMyZldDk44
jFmgTEzrIFLbthJWenCBW1VL/mSDcisQ0hwWF935GUzaSMjYfhAwE5mFTT58A9Kc
jyJGWUS80oRHyTzpTL4goQGGnVlwI8/zrZOOLegkRiDr3SIfiV+5I3O+NOApzGHw
iohMtFoNJ27k5yB/oCutmmNdKjHMzk32pQgWBE4nZ2wMxnk0w7NYy2/+nwcV1Y5Y
JUnTlxNNB+KLsRnq3sdjDXG/eaQhwMGOJHp1ey82857WG5ZnjTV2oNKuBFY7MAMS
RNcgJWYILD3idhPks/7EhoNpBvWjr4jbN37G7BjXfzzHYHp8M2+j+zVW7FJ3mrPt
Nz+MIp7pmjACmkNVrzEQZw45pk9xvn8H1AhHs290sGILWbvBVfAJ6JIW5sU48LT2
dJAWInkcQZ+B829EJU2Ce537ZQKolva9TBA5wkg0YRW5KIKtjf6VX8lpm8/MYoV7
ncTlRMeuMfuTLkFEFufVScTivzaAT1uMFD2z1PTPx+0AN2SFk3Y4VI2Gwbp+Cref
fA0p/YkvR0X69FJWJPXazhXXt1pFfKlGUg6Iew5XCsE1qCWqDUB97ghBWW28YAhR
ObLJeYhHyGFGRW52F/pQ8TKjzDvLifyHyVx1uKbKYtgdYA8Vr5+8lMzuI8YUpm10
IFZYJ32GZ/u27W4LhISRSA/qoJkca2ioYmW+HIfCiE5O1w9T3o5ujj9WINgJfUO5
FDcgTYJlX+zj2JzmjwglswhGibtmlodpfR1qqUINENZJnEwFeyfhbdyjeRxMkKOY
6MNPrbii1uolCWHmwCf+TlOw4jiTzxEMV0fTYnuoo9fqOpNhhlqghBWz0oAsSlFf
e1FsC3d8s4px95eAZ22xqspIpgrJDU+cBlilxk/EvhnUsg9NaqHqcU2f6YMwcPIY
pmUoS5mD/cdcB8VXpltEEOGApZZpsPULV8Z83e2jAtmr3hG8BEuAuY2eEBbOmmib
9bApf4i1nTUHu482nAoI6HISPr3niSdP9WuXYTeadOqJD8fo4sdZw2HbYfCUWMG6
JuKc0yApJ7/dtcyP5e3MlclFrSQrWN+LHsDPtpO6lTBGFB3APuEplh6fE+TxlcQ7
UYTQy3fNTDCKexA7h+3pxEfv/RocuPLQjbMi/xZTWgg4asA/z8VQF6ETB+2PhDe9
K9G5wU2XmOeQe/fORNvTw488d36LRFFaDczohPtqEMIe5gng82dyCg+wB1puc8Cw
1SZDE+fWtH/QgZpyCbFiuw4hz6QUIiDWzKBaJBQd94tiSGj1utwcoCgjSxTl+ADm
9dSdkPvQWNrHtSqQNFXItXu/Pf2uI9TEKTUD+jmu3RVqiVEUEpLIGyC/Y+ik80Sx
Ink0XN8k15qAeGs/OggSn+KzH12B0flk71+HoffKV2Wu4cPf8BEdwIBE/bPGS+eY
KCOGqFhrGkUf5L01iqPdwE60fXEYVbuP+0yauGe8Q33drEPcnmJ0vM/2xHgkwPsp
boALEMJNcT/gnJCdnIIo+XStvRC7CuciEXOH/1yo7Dte4qL0x2m6sWe1qVpkn/FW
+BlLXd1/uyl+9quuQdr+/+jb8r73a4UCsiVR/zalAhQdXeWP4FQ+v9iQHJ5Zyweg
ck5DXf3ha/7kEbHPv0IDGYJY5Zn7GT8cGrDhjyPMe2JCapd1pb1L4pj3ybeJSvWP
H/jFWXVBBbvDGUR4SZzzejfAWyDyrvV5skIPfbY7X0fUNGGlYBwyXWqK/eoEvQo9
aiYhq9Dfj+bk7CAphsw9uNFRu4JBCd8XUDjKADeVJBUuwLdD8VJHwjaGUrVvLs0G
1dwrlpyiLk0JVbxWQjGUj0WFjWlGNrrKN6Xy277Op46r9nTjtbCoMMsEEysk7dYs
zuBouB0gYPT+MiX8dxHWqZ0/3BLTuEEelhkkRoyGs8RFY+NZ4VLUAu63aq+AOBTa
wneNIU5xaiyqOlVg0OEEJJ8pVk98qb66objRbR9stbYmUmEEq9EkE8jZv/9zgemG
FDIQxKvHRvMNar8gYBTqWbXVdZn/WCFSSIhy4yvzuEViqnF6N2fy+CkhnJXKl74B
ChYx51Q+yFlE5dLBxphw9M91dg5tvmo26WQwp5pYyHA8NUR+L+VClXFg/QLv0mg8
wI7gkcF0GddDYiIYD1aOkPUOwZOEMNp6KCsjmQovq6MLhnigUC2lqW6RJdL+rq4b
WeJSv6LElzmMlHbUZmEdinkued+4g5kDIMMm/UJ99Cc5qFaEZRoLcCFwxnpWllj1
QqxVSk4FoSXQ2r1uD70aHBICdvNkTV+7qtbpjWMYgA3a8YFOpnRjMzmggn+CcZwi
jMYT3bD01IYliRKPvMFISM++abmtJOfdhxDjLUYIk0Ivea3Okk9888vHQkhvSKOH
Shl6XnYlS0WkCx/UT3SidHERJnoUFrmFPcUelheJDp36SwpKaPt0Oi2XxwQFmMtT
PWuKtiQce+0VPlG8DAUpmUmnFELY8tke5nmOFsrd850Y/OgeZyOvgdVYHzfVBT6r
0E5w2OIeDqHEFCS3jWa6WuiCyDMPUkDAk7dlZ/g5i9Yp/sPG6Hzlv/gGAGIYd+q5
T8lvYbb4BpNcwZUAesF8XOeztpvYODnU08IihEpGhPCpvUlTW0AHIQ4aqJK6jT95
LpHBq0J22L7PuNkja6BiJOraMsLk9z2jrMA9jA48ahc0o4RelhbseSr6/gzXruWl
WOx9P/iInE61IfCtYdVA2uALlE/Ia0A3csgD3sTh+lOyiszOJbt4MzA1k52MPQ1E
YXtFh/9ULwMpGW36R4dYp6IVVSfiF4ONGLigtqdYADz8Dc3Ekzo8VTve1sX/h3ti
F3y3rj9JxjL0pG9Z/w0qS1a8LZLC2/dmkQxmyY4rdUaE6KyIDrPpgy8DvgoE9DEq
ODnIw/ushPQV3mOO699YaVVTwOj8gm3tR/1de87o1+arsXkP4pQkk3dgRO8vltaa
4mA6InL/GzX/MORbolfG1jFCJu2MHTEfZkHJ5ukldJ82mKqqX1NHLf/G6h2rymRU
tBqzxuX0wt4pgb8F5pr9jg/7DHn4Tnw5z0W5rfA+0E/zDdNFGNYDB8dee+VDVTnw
+Z7jel4D7pzPO5CDNJsPeTJcIBvxUjowJDT2vaX/SPc7k4UyRmWS3BD5rbwMlflo
F+RpjBPBxH16noYdl4bMbbSeJG+XhYas/3CwQyGYbK9oHt2HRdJt34dGVe1Teih9
oq3vmaOfF1Lc+y9HYrvlVtCQae7Qxw3oduOVXWyAvnAj1lRKfjpzAKPIgGUIybd4
loZhwddJjLcZf49S9WFtu8hzriogiOUO+le4uaivOES/dJFqkxMTj7RadJIFVia0
n3FlH4lEBnQN49gUlOFnsH49l90rMkcTu8VqZJ4ETSfnKj4AAGmVRS4i2Z6JdJs7
gMGalnnqIzh8XVM4xTgrzZbq07BiiTzSex/lGgUY6rYlvRpbJFnUy27/+lf8C3lU
VMHf5is2KV+d5xFu5kpsb/Mi/3LYj7nQY9eKI6/m2HbmqlIqGfz8399OX7EIGAEJ
y9dqXG+sPFdJ933FkHl3a3XbOzTxoTxm/DCw6ZbnxQUJRaEwQRBFyTTwLKo4NLmO
AUntIayqDfkyFC93ZKklGSFarbBVM+IYo5xjjpsQGw39U56eF7yqkFhSxzkximFP
rjwCSFGuEAmJO8f0mp+kivkPhjsEmXv6ViowD2LCvoSbtE0SG4DFaTo0fjWo1hLf
DxZRwe/dgMcAzRnlO536lwX4NtF5kqPwlr0ItFHZrsCRq8pOaATMH6rI8zr7zaEB
EGqDfKjEUcbM3ofvarVejQl42IyJ8bHS5ecpyfCqu2qDEGBtP0SErM0zdK3eyCxm
rR9ftD8M09Xnzn5XXQAHI4V0BXXAYE8v3dO4shRENGd1BxT7Y/LHokSwXsO8XJlR
bs8CMP0DQ7gSzbGHU8p/m/58ebWIs2FVVYLiIjzpLrye1Eh25ky8vJfgsV9ownrc
t1yaO7lPuHzRThLcF1RXE23+jx7grU3b3UPLYK5wKCKD/LNjgiCA0Y6GexwESvdx
bB3n0jIrkYIkWv15YEYjx1LbL8IJcukf79RsjAeyy9lMBvv58PJhlCLjD10GXq60
E87UhwbtQaRqPRi7SmyO8OXAd20vKgfZQCY26Oqn2N9mfCz0yd5dB9g1JtZi7tEr
p2e4mMIYncwlY1uKfuVIPbHVQo+pX8YsSgo+4iG7OcWoYaGD3mvbyCJTSMCwehQ9
ggU88qE/3CznnGoeWo7iard+HEaRgrfxS21LoCIrd9eY7Tm3U4t8LcTSWrMZpfyb
AZvvoAp/4/lckNSTmBiC+7uJPkQEtolj0Ww79aGNkYM3difkZqPbciQJ1+R83dbz
RYceNz+yDC0LdFJzT8hxIF01TBusZJ5akaifcdzuYZeNVG6FWORXEbgu4owOvZdC
EA09BzJDULy0inT5jhsFTSxa+TUwNyRFuDHRHOXRu+87pkDa/IBG9LHDDHf1R4Lw
OV1W0RLvpCKD0+2z2cdXkDy9E9HcGEhYM9jlw22pf3XFNv70WrXa++EfKUQMwOhG
f0Dbf+PeNeeZ9Z+BJlMBdkibsXipHrlHCGF46LpBKbPgrs0cQsamusd7yU8nS0U/
dfc4sxYpLTcYsEBr2UsIv8rw7vqOTNHVFJ939yJcvo9jvwJQ6agQCbVNXAGgDLno
a2w22LjYlr8zr/+jLAlE7nx7cNcysG8Q25cEEfvWOtmghM67PALxQSRDLg4gxUpe
EEyxFwtXAcIyBdJGMIUpV/WlpFPwa+snIgK9bceWvMuTAUPF6UifANzlw0xZs6oE
T8911vT1O2YM5Q9StlO7XTq6TPj1XGnsqGk9bwyeCUYtW8f4ddFpe2YHMjFg//vm
9L496LKR6+fe3OgWzop6iwGN1YKTjbE8yEfCtZp/PNMEhRh6yj/CDIywQgn21P7d
vFB4KDqwTL0yulcePM587A5b139P8hxG8SIhdUAlEbdwesP6J2EyaYDW7NnDNidc
QBj2C7xPOg2mzwHYrgmzDJVl8egzexkHzuohEh/MMUcH8aIWKTAUUlLhWKFHmQ6m
Mjawcxz95Khq2jdeAdIWt2wQefu80TpK5jwLtAm0eVThSF350RABnqmc84K6jQva
5UxLSSJndN0RhILyTdbwi1CpgdWnugfm5r+ZDnB3R9AmN/00OGB9seM7EN19hrqa
sHBsZHCdeyT+CQ7ol9VWo6PMXPwP3XXogjbS4xuKbkJOqhFbjDKQGrTUTEzZwUA1
CCa2ylIfD7x2rtHGa4t3MWcfObgtLqgMLO+T4h1B5Ovll4KkMt6ahLiBJ0zaT7Mu
mXgjR4qjzoCxJo4j1SgkRzewN2uprOJWI1asWGBQL9yimNh/HA8+bhYHsohN/0fG
gBrGQ890aQG6Fg1fAy7Gn44jMDoymajq2AuEiXQ4D3/dWZAA7hAXQh+Opw/OG5Gt
Y+aZdj1yUChYT2lEsdKA0wjXH250p1ODPBF9Cxo8s4mJBlgYPC7u0OMWfwEdYCMs
qE4ZjFR77MwM2i97/PXDl/YwUWOJTnaQn+lvW88NDJNKCIF/nZHZ+4hk/G8/2Vmd
mZogWd2SIhMiu8DmfjKc7LlXkw74Ybv3bDvQajDHcFFyk/PUnqtsOLJRn4cqup7L
8abay/cyELs++/rxhvrw5woSSYsrz91ozre0DA2QNfXKXz/vtadsdxT53f/gCXhV
DVLvFZ5eRYFzw6HmmGZJb0e/TmOwpBLjnYQIJyzGadQ0J3NoAct9A/k8ZwMJGQT0
bERPrBIxFeVREJyfq/UfpUuVYUhlAzbv/VzX6VkhQE7IYXmxAn/OgYQHBvfd7IyL
nZ2KcJE1+5HlfunjOP+vGWkhk1GWLgRwTxjBapRKiISLVyDuQnA1sTlF2/dFjsHT
wj8klIXFsTq20etxH0je5WN2STmcpT4a5YHp5kp0mN7mdjbURLnwP+4k9bn+Qh+Q
g0BMk4cBsGtA1yAIEaHqTuvJU4QMv+IEcu75MtFMDzeYAa5YigFiadzxCj5Nqocl
td+EStpksuLwnNQVUm/QIu4+BOVzPC3qPSWFL7q1HrpdY81ZEw1Y0rpyjtPHOpLu
jdObiIagkkIK79l2Ye6Q0yThya1fna1m0n8jB6YkhbrYs5oqOY/JaFd/uAcAc8Cq
Tl8H2kFs6Z7nlTBsoBTCJcy1NJRNoXIcGZs+RdHzEFxQgDDZBwbajBszPZoMAYz6
xYFzo4UEo+9BU9jaBJ+3mnTsVXhZJdrWDcEGz1MawrTs44oHFYw8xsiN/olfJByw
iIyaJQckQlqX3ii6ccwbJuve5Spf4bM6qbtkFvcGvEDVO1MAXxXrV3p2nnjFv6uv
nvkWq9YEzChCe1rMTbUhVb9NWEJDWs9zVfAbiUHtT/AVF/fuiLMJdAG3TeGP5U+k
L1arzH+ExUfSBdj20jWj8lkxANskrCqY0mTRCodC3rwbQGq+fEpoh6EEiPSsEnB5
Hmw7pCj2ARYs2yxpMAR2WABrbYB/BygwAbr9amh5PQME8F8gdn6R5U38HFLl4IQG
z4OUpt5K1OjJkRNvTiAH0f5W2+9ev7+OrqnI0/WMUS4fATaPVnfaAA3HbeOlOf2+
y9GdsG+VpdQOWgnPuf0rgij+n+/z97savrkgF0GUU36MlmIil0yPVJZCxNBFC1Zd
ro6mSL0hEK4dQZfA4STxzY9wBwh1tvmBKFKVFrYm/jtZptwworARatrFmF3J0YvD
3bWXEyDMK+7bKiNIya3zP4weoGCxZqanbC9ifjFh2rrdMJKmFjo2OqDU5tyA26Pl
XfrtI/6tg04SdETxCj4p/lz9IqeOoW/QAbtCKtqaCek1FKo9xl9l6PSAVu1fXqJP
VgPmWEKEckOAahaj6b2LMsZqhHHza4brjM62QAzMU326gxyXjmMBH1/OZunB8Ylo
W2VvaCLAZk+a7Tb5f1/Qw++0T+G7frmbQtm6ez+CUtO+R+P31w206vT1i/FzQsAO
opJa2hQ5yazK3dDZpOQOcedzHETcfXlqfnY7CyC7CstsR6kC2uGn1oshTcqoClYS
E84i46CDqKCWt03yoTMQNI0D4vPHQPMC09TAK4DDeFLIfx5INpm+kCzs0dqGPBL7
QMW3gSGa4yiiVoztjNIR5JZBUxwjEdzu7wP0QltQpJvF9oGRXdPSyEpaaMgjyUHo
IfJc0eVYXwdo7UEjS6MAud25c+ZuHQ7HP+E5nJ7hNF+bZcZCNAi7ujHWtacFOX4d
8G3Im0SPuLmzuCjPFBzWnFgN+CEc9ksuKdRlWxH0EYGpYwFcxbqORYdiaOJo/fP+
SX1xJAYyhy6+U5nDJZbvE/dz8rkomgmoTg+taI3f8dtF8nFFLI6JXSE8MkKrzZpl
aH8nSlOQN7w5dK8s+Quh+MG44fXOlFNfODpl8I6iyOieAiSk9zXSvpoJE2kOSdDL
hKn5Oj6ka9sD35zj8j5ks0WEz9J7bitCUyGy7xXfZs7o/uuhPMMU+MNJb+Ld/tgb
7vvskuFLWzoPxp5Mz4mWzn/cIsW1TXQcZ2I5k2L2wVf8dpz/M3B0RbU3iXAZ5XBS
wssxvLL5GePE5/rZ4q7OEWadpBxuIcEizEpADTtKsChz13zdKksZbLQIPBiCfbv/
DqBKZuieBkCVugAwDmYnbiSIxDd4NU81SVpHecrrNw2hWwO3IJnGO5x2GiR9dmbN
qFggd62guigGxPbMm8jAAk1TzuHg6zpIE3mV7hQi11RZgzy8sUErGRvPgeEcpKNZ
3nq1eHkJOWhNHN3Sjf0hIQKlqlU+X5ULFdZW3JBSRSRF0W6C/b2umAyNNWi5kPsV
UB7fW9k2vPWHOCpLpYnRZFtxrPtE66gyX7hvGxNORUat1IAVaHq+xdyJ1L5aFtst
/oAD50Y2K5ohVQkIIy6Tv5iOZ6hkCN3F4atP9LDxQSWHHCcH3hg/0fgYnn2ATx2k
o4WWRb/4kWexiqwNRKSBt3HDH43Jy/SYfPwU5pKPvZ5z0BtrpTeTHXEIi9xlO8+l
HzMebloNfcegIwMvXXjlBgEfZBBVj3OcMl0qCMZnli0Gq3S9D0lD4jgzK5qwKD8a
bCVieP396F6GoZHDOY6HHIvnKFJ5t0ME8ulf3SX2WxzIvzU2/ixhjenPrMJ9K8DE
Aat1V13TkFdFl9JPiv3EQ0uqPoeDDRuJnzQUce8ZimXJ1JIsJFgdvw+Bi054/RM7
2gXIcD/BPa7gvNSZSxbAaLpMHza1Bq15ZLx9EVkCiVjcc4lRyTC8+2uYWfLqUlbj
Cxe8yscHM+hjj9XVIzAwL5Dde8hLJFQgbYzsSZ+FiJO1yX8nSyj8SAkc+mWIkVca
Po+/aYbLWxwWkIMD4r8uAw4Y4ThgXCqctuSWXQFR1CuK2pRlp4w1l6qedbsQerDj
riPRjMFvRqhaZMdpdDpG6PCm/Iglj5y1hxuT2tNUBMC233ASX9gvSF/zZveiarrW
sq+nq+YSDQa0ad4B8ZlWKUtImzcjEkdqpbrUgoT99PRAEdMEwv5SHTrRW3fVJS3B
i3eOog4fTptPMXYDM5vsdtSiZs0uphNOSq1r/34CdOQsJYDN0yT75Zn3fQ+e7oif
T02RGfVcs/UlWXzmqz3UpKvvKRRitQZ6kF9eo/pSuOvuDlMay+cE/csq3Iditrzp
7K6RGn7d9yOkqKhhxq3P4nJ1fBO+fIG/zICEZUAcgW+ZpW+TNVNliHhjEMfVm1tV
czBVmUFG2yxVtGFBLP6ZcL6ftcQxU0AWyEFWARZEuvEuiF8yZ60oRGFpL4k6Jr9c
lnEiQXvhsC3lOwbou0FL06+GPiXAXshYFD3OhrDxV8uldlYMKQBwsLFEOLoKhLfN
QojEPOfOsjS8TMktcvo8ZkYzD7U+IGaOIldpksYB74stBzqwoDARuL4u4SPrHzmX
ViTA5/a/QuecoogYVMEz4hewQ0h0udnEJPLrx11bbEPhEGw4uE5ouhyOLxXyBD5D
DeCb7LgMCvS4uvNvk798Uwn8Ixn+c3Gv4vIEGfJ17ytFSpNRbPLJZxKFfOgyfa+8
js6D21R/BAw/PgDGMuztPnGCcN7ADOWWSInBh/LiCtc90LsgH21haPjs5z8UBKTQ
OoEPAYszt0AUzaB5AL2FAA9bPfPsZJ9fhQbkDEoF9RMEt2wPXP+af3UCWfM++VWx
Dw4Y+GCzsYwY4hdU24zWOKu4dYIzx7uR8IWdbX7Tu17F218ul+u3jCoYCVi9PX/T
Zo1xhD7uphmFxoT/VjT0vHiboeFkWdHFlwDywjhQ29aDMiN45JFMEDoCiCHc5OJt
zoTX5jVlIKF1Tr9Tap1GUou+a5nbSsZDHSEqP4EwBNlCMVpOFEmb3lgzucOlESuE
Q8ARxN+4jZxPdT0ZVe7XPIgrQtydd+AV/9nUHZLjU6SSwX1vQqKwuG3Tz2zMZybw
Goyujnxi4dthEq4XPcl5TMVm6cOgZTVsvrfxPZIDjaibRS+RstK7oeN9u1CKGl/5
c4UX2hTy5n+dD28CvBrGxw8PQJp9M4H7toUC0E8kWlgdofiRpwkL0WPNSl6GwwSc
CF1Uy4b1TaG+1PqYAqN8hluO02Eia2DtW3TwSqjvYHKPDL5PbmCIw2sqpn7ZWpIg
i5h2ULZUVvhvHOyQSmONbXzePnpHGxubA+60AazQl4KdV956gAkpgxKq+blgMbFP
gc8FrOq7Bmykzs9lGbYtqB0YDG3D2haK3GzSj5wlD/aqq/UkTwUi8Y0qmzi09sVJ
W/wI0+ZuxlOXfJ8xhqB3/c4mKwcqd4V/PRhCB9aIQJ3JMez9nWAZA8TrbeSwrtKy
GjRtnQgSbc3ZquXSuGRTChFDBZdvxp0QzldK0kjDQKENAqCtin6/fcKg7qxUuzSa
6pLtWjh24gH/Pj43UF9f1GHPbmw/+HnYWJ1hxY9W8KmdO3aX7kxwLMTEiQ+FKHc1
rp4ZK2Cx0yopUb7RBKH30rjR4SeI9n5k8PHh/FSVTykCuChsf7o5gmgqj5NnIW5m
o5O+fh6mk2UoNTWx1n3egVx+s3FOYNzo1WVHmE6v3Pz3zONTyAEUx7m2tCkOTVf+
h1b/OKMqTsF1/vymdl9ohru1fLLuwE0xSJsbEH4g8BRlbFAMdGkZhujyAEjsBguh
4lSuCwbwEmnnHtV2f9Gw5AsEalNDamFkZCXvknN7oWcGkDd7Y+PzUbwHClqJRhH8
0Ia87z93PT+9GptMrjLCAgcFX34O6BD3NrJtSnnSmJik9uF6RISs/Mb2NKSzfG44
GTMrD82ujdFaNHJGhhtoP+Lga89V6pHRMFGMTlAFTyHs4AUOd2O9U8Uymm3CKzAl
pBI4EDBT8Gu3kwkXzz9IbQ4UrbSCWzH7cuD0jg10jZ4lMHg9pVh79SiRghSVxJ4o
O8FqdZqUG7fT/wgC9bDzR6PiWga5TGNUQ96ah3y5TGHDjglMVn1mBdPCoGNpc+1+
T+7IWwRlpasmr10JR1sUUuOKyD3DTK7qKXLhAKT5xrMF4lS8S7N9PnmYbMGJLo4D
dfFrUZw5SNWDxwU604YAs0ylTCqEXnWAgG6GI8kJlmHnhZN+p6qw7yVrkCzeFlCJ
ippb3nqOiKSTjZKqtJQL87qgqYcueJJerKSjXTdvYesPIafisgufIAomTfrXQWfb
1gvuYUOkwNwDG6C9Gelu3q80foMp8znhLpsMhVVkqXvNqQoYvUHDJUXlxjLKKDUp
luxpwMc77BQ50aUgHtWROpmwmGQ3OeLId1OwaGEWDA0D9V7+eypxhUZyVhPjzsjn
9srrF4WIE9ySvEHmD2tu+l7IclseHRgHWNsAOvDSjnUkH0SwN1a4Nr7QvwyRlsJ1
2wUs2NyW8fS3ydfcax5STE0JXgqhUpcSwz5MOvJ9h/y4Gt0163dmUuNTOrq/9Ivj
qMHrZKphOfVGCBktL0c1pO7phKaCV3Hj+GsVgx3XBTyj3CNMvnELJVSz8Sd6YCnh
Is3GVCsSRsjkFsPRHJ/z6az1Uou72tCwYehV9O9/vLXy1riSZoOFyQ8QOYxA27x7
mEaCzG2nCUWlH96pxsx9un6ztE4gxRhk119w15pIC5SUG8FSVNakWnundmttA/5N
vRBFQDQln3beq3kfmp0lArM01e56T0qyvIhKJXiJK2sNR//O2GMZGNE6U/BhoQYi
rs7BfSjxAekFeYf9HTam4K4VB0XqM9oCtTrcs+znQTykccOH8ug59KkF8RtNsdNV
uEJQDLgn5Pn1zexUeHEX/hhOK6xhfA+YK4UFJFZ/9MqhtBVqrvxvFE2UD/SMToo/
mWFcY5ekmp7CkkMV3u2aN1xRlG/fTqq5Jy9Ju+s5zGGq1TjDg3HO+lfNeJc8JLww
Oo0J1d2WjMjHjcVXfx7Thvsu+9UzCEGd1yxlC9B9wkg0RUA62srTyv1YkJFfxX/a
//Igd/KR/koKuLCFF8kG8/ivXejrnNF6+wCqbSw/VdxH5vsA6mDU4cZIQChZse3W
LXgou+dItFQt+bsvHUKVOATMjazim8/5hO41bri13zEfQlGUYEZL2Kcj5RDnl9+D
oSiMrYRiRHaWPt1AKYN+/n4E10dDsbuOlO9eLBmK/4HVL5DXQ5W7lAkocPZrchni
HgxoAvGQ1apuiGl4e44I6mh63vsI+sC11M8g/QgJ9i5z/3Lt9kQG8NWy8vA7apEl
1GN2+fdjBGueO954yqcs4pGeYcQ/arJG4vOCMVvq5g0mnEiDIjRq0nDBuizG+YQ7
LprJKkb+ZR3Q3cS3VLeS9TwYaUHOdOXDXpbtQf+AhlyF0h+irfXJDkRVH6haMV/k
/flHTLayzroXfrrYEBBWt2XMwVFE4sGIFZfjETeUUknekQQ5sP2NrS1mEKZnGpao
JyA+jZp+TlKOI21SD1E30CzU75MPa2AELjPJ8dkIWW7zUfUApL+5MgCNKQ/7Aiwq
40anEYXPpMq+EQf/brIoA+3eR3uwVZMjOgwlKWcvO0H6hJ59903Dk18+GTN2YyG3
E6zCmqEGPTwKKJkQb01dja0NaVdk/1Fhd8lRiPMp7FBGX+PdXNjHxPwTALx01N9X
qG7eanjEzqWlxTHi0Bab2/fag92YxKokUS42SRv1gMsvpXBiDpUVgZQmbGBXjEIf
Q0PMQvDkYXksV6mNHN87hLBPB0jrtKViWYHTDH0P+BXGXe3gcfRJbUoHsvbQ1mi0
WXVOMVWO8DzlTZmGcx1bnB7GJBUDrrIbZj4w7BypQ49W+3qKVcxv/2vXR025V8CI
CePjDRN7E+r+U4blCc52aVKQJCG5iC10+VMREUzFSfdjGzuX610DbShrPFANfq6V
/NubVIruLO7gf+Lx2My1s8UR3hde/74JfG7OpCwFIvHsdVDFNDTRM/1JbSs+le7H
PmU1teQMfwb7eKQyD7l/DPC/NlahN6/Cp1cZ/lWS4OIn3EuQRt272zenyAXyAftk
m2usTs2MEsy6dT1ahP3i9NS0e6QbTGWzpo+vOWtto5sVA8XHEiLel8GF0IzFvId0
vtCcZea1cJ5a+mxPGFMWBVvZRs1Ekgs7TZTR+Qi2Yo5CWEH/Y41ZRpmJQiAE7wti
27C2XfvKs85sdf2S01yvqRbwiT5Isq0tlhW/rPbEKl45XSwjWSAXBQKYldzcpoy3
p8mek05uGlq5farqjnL3VDVmmmBcTZ/bjBP9R+GrZaJyl3bWbrI4WEp7DUOPzyKl
MhEZKgzfT4tVageHTWkNi66Xr738/SRnr+yLpvSHdj6ffoaGw3gA77WlzIFFkfJS
FWmj1zJU6tdmwotdPpXEs2yFm3kecvPY9nvUzGbTNidzbKe0dzg9Pu0HKMMDScuH
JrKUPE7DOwXZH4HHCpBUdIPNhIuz1eHOl9mpu7FNr0oJftBHb1TlBhT/bOOqpX9k
oZ7rlg2IZa9HTWFRPueGkMy8rUCw+7iqAQmVHbFngQ6MHUKfzSMnQ57AgDvQFKSs
T4MoGmCY2tevvBr6ge/XHltBpmuJF1O4vQj9Mfv1CGuJo+pEATB8/e4vaUF2jSlO
VNZYmK+XVNT+aXvCTvfwMtWU1ucqM7EHu3Yr2n1HoApT6MHhcYqVAZEVhWYVZyJC
RCcp2lem0DahIbkvnChDy7jRPBzS6BVU5nJutYN452GwqytzTZdDtvQ3WrO+PJxe
6uePEwmrenHYoTANarRAx/uSfzVn6T6V/fiZyNtG6CDE/1feZd6knsofFrntpxlc
6j+mzs7NFH4XraUPVdLprDUIVlEEOQvSIYitIcv3c+5CsmV/A85oEAAISwQp9QlC
iB9ye4+I2jfY4TxrM+PIns7y+JIR04178NnezOZlebKoQZC9z53cf+YuEGwFGYCI
qJ6KsZBHx1CcpaaZmNu0Bav/By1ObE9feC+gY/vJloAVXbO4F5rwAuOmI9vpPZ+I
zz3Gz/cC29jZJAAAQV6P/yIDzG7DYefDebFPD/p6RT1nowXhYzX94jNh+2tQduJl
tZVgfcZ6ErlnGTc9S4WqDegR2gGEGHo2ydIg13qolJhd7wSvo9/dz2ordmgBr0tr
j0KEHDwwr+eIl/RFLRWGVrw+5jc9APKK3rgj0FefwXtDTJTUZYH7OG01T9o4XSLu
Y2y59N0BKKVn8kIIs07UOh+eDwtGnDSzwkpzltyi53o59mkVTFoI9SkjMQ3yAheo
B+OHRIkrU+hQkNWOxwShHPGWeD0VoLmK/dPWZVLXGLc5t4v9m8+zxOdW4JmUXb5B
tCIGEmIDCq29zOL0h8BmJNriF31Lm0DrzmqzcQNBW82BQUTFQyAKwkKpFFuosL5f
l2+6qiIaZLv/VF16Iw2FOrTbpECzGCKG5s/suABXBUp9RFVc5B77zq1I4YSZ58mD
zDCH6WQ/0JqDUauVrkw3rFM2c/SncKWF3AXnMPHUIocKQzKf8BzJ3A7zG1RZDA/C
vSskdivtFXpkFcFb2D4IplHM/n6sdqydeHUrBT/LyEgz8GxmAV+roIy2x5TBmb22
TxVvSrx5CMi8KrbWBxAWyXyCI4UOEdG+CQocIDG6KrVAUEq1E965gOAN4r0ucyS3
4FIbQ/z7FWL1HXrUNoTutNrKfNXVrePbEOenkgVFg/dypBbRKP62QhSJ0q8ZwpK2
qzUesy1tuJr2NgnAlROy9ZyiIgHkAddduMEcr0dx2j5GHUkVlEBnaFf2pVFzEly5
BhcNwoK8in/CdBsuelVuo+pOikSB1mI6S4aid9MCqj41vb3eHTaU7TFHL0i3WO5C
+x2rfPmJXabzcdHWJ0rCrfhl1zM2gA+UxVQSx9fSllTIr+OtkwObxEMLPAFar1nd
Vn3kg1JxyL6dOXrhlscRJs3V5kRAd27Vi8F5GQgpY/xEPDLayHbmYQXzuB3KDhGd
s6A0F1/O99ZSyF06UMTiqY0qcOFnTHfjfuZDfOJPGrfPg8PqB8m2RXK++vH6YKwn
mXrNq/Ijuoh76MpQ/HJadwduIxeEA0E5w5XGv4PLLz4RAuRBpHzw6V959lFylWxt
ViVD5+kX87SF42/XeFBDHgazGdihkNQPsJ2/UU8HF1g065t83IF5B6a0ctzxG6ZT
Hxwrcy692O0n2rdYMTVaUVg9/SewSTqgXWE62WkHURvyZ7/wK9s2Ev+OSZudNRcp
jh5Ku0o5m6jQlDhSCRBu33cteeQrcKKDwVJO4WXKO04yGbCyBETlKEOK1yNJt8F/
WNMrVrwKE0ueop1qFG/wA4D+ceYXgQyHqwwpn8YHIOn+t5T9W75vEINsubo3MNPq
8AYH+8ZVPOpB4VYct8MG/KRp7o372KNn8c1D4cEhSL8NIdwmvDqlKWklDfhk9xCA
DPNHQw2rSdxz+HCuj7TYZ7KlWzC7DqdofSvfOAQB/gKnSgtvXnzeXV4VDPYyYG7r
HxhlZ4MqJVBPTjtDo75u9evlPpywJb0qOkvikFtLvh8Wp/aWC8hf5ZxdT0kT7/0/
15UQXCDVR4bddrNw7fP6hnTQQP08CLqIk8BnZdRaIHbZ8tFujDIvPsTT+pbzAi+N
DoCRdVcTAvXQvE/NJi6uJUH0FcKH8AeB6BQPLPHy4IoMsRN9sGZ9bm5a56WW2z0s
WPfwkWvPKJfFJZTbadpv1+xGmUV207hMU4Qi2xWtGI7DPakdIQPV3eprvX2d7F7F
QbdwoEEiFv8Xa6+JkNizQgox4HPlxdwybt5uFP4pfw1Vm2oXLveuA810AqJxsDJd
V/vahKriduYMXf3BebWL0FSOF4SWWuPIBfr+/tgXNNVv3TYVagV1SCdC0pHmh7IQ
xIW+27I2xeToGSqp21Bhvkg1FhiZ/uIXPoOov8Z5k8pwV/f0KURL8VrJux4BwgmW
b2bUqCDesGeNmoYQWtUQPc3tev11eld9kbxhm8SO0yoxZTOF9G7xMuHsWU5J0Vp5
RGVxfurxzaGbDgw5f5JIeR0SIzDKTmTZoq/7mnkM8JWq4T065NVggwoj/XHbUCnO
UO7eXzjoZy6pw7tPQUnyu7QbscZQDcbE0X6BGWVcI4Rwwol10C4bE/N4F2FdW+5K
apIatZLp1Eq9bJ10QzP2oOQo34oEGWyZHvZwnOdUFg4ydIuBhdJKgJgGom4Wr7Ow
WH0eMo0ylocv/J3cot/m83rad+jjcJXDOb2AXRbUHXIhJoCBnEGnxCex8OAwEj+q
ryojMNUPFz3LpphWgSghVo8aXYHPVpiihwJs83DD/Rqptwtw69dVvjlwMcq2GjOo
wQ3BnhgQRZJ241XIFMmsXOEjJW1sALTeWmLlwen6phh0OskESLbmH5hKNYRdRBSp
/JjmeaDj6c2BAuQnkX7cZptEGj0Jh13O7Nk/K7UdruYnqqxQOMlF77U+09CT+JC9
U0QHyUJVWr1HQXodVpieHC/GHba/ssN3/ep9S/zyBsf18iHDk2Qcg+wNO/xWPRN4
01BjMRnd4+HWowT0K0hbqTPdBANpX5KAXFVLr8ivSKs7WDiSOxLVOT+HkcSnhoQE
m3G497JGzcOzqsKQhmTep3VUiUr1ZROji6OcadKeWK7o+4EkG7byGm4pbCgw3mch
fg6BdljOV2JCMtt4/vs1KmcALfDu/P1rxdKTHaQsK2aWhOqm7ssVcyIleueHfHJ1
3bqw0/CJ2mS3yG3MwoS1TCPiuQso9pnVRZOIoRYJCpvVR9GrrcCUfjH4qBS7orRC
otDzLF9A5ZQLcqRiPQ/im3bDRnGnZ5nUC2/HDaCHLAmcah3BYYA8nALEBZQvasWS
sAAtSlPJQt+EDyV92xKYOqnbnVc59C4a95ysZ8wcWJQCMEdB1kWlxolhdcRYrViv
dwvTCAi/polaQ0AvFWkmJfmL1K/wzehwGpxABvpCax7z5VMkxTQd72w1bSGSOHU6
O6H9ho4rXuQgIVaEbiXf4Dnkb+IsyoZ5LR5YgoSYOAcKba/Eye2PuvGM/+h391OD
OxxmqM+EPBxOcHV+JPd5PNA0bE7OJYlOr1bpwlZmJjWwhy8T+dI2un38ee7MfiTZ
ftdgKmGw4nOoWnHSjrfz6cTlq/eU6k0goMGoB6Q1VoTUFajUrBT+BziNkt0LVEq1
jTmWavXcTDeWjcphgZPB8WjRNiSF7uOqhe6wc732VG5gad6Iwi1zSK+hqJXR5gJ0
WqoqC/x0uSHjj+PBNA7acmcXyqWl66P5TlHzi0ygTWerqpfRGobahqR48mFpMrby
53+3eWI/bCeaqfMVTL3ktL40slRHpACmhws1ylG2k/QPs5V7K5ARUDi2TzLoiAVN
vVKnhUF6Xg//ujK/F3YAF1WeBEcw8C5SkSDmobUgfychf0oqPfWBea6zcpQRPZNu
bLqwjpKfNuyJgtJ21c6tt2sPflNAN2mzZgqaLUBm6vf45y/KL5SEANwPecaZ/pnm
oAPf4dhtQn3ZKGA/bGdLRvYENBys7gLNl39gqQ5R1T9ayPnv2UKHuGDy3Z+wV3NC
EXyYA5yytBKshSB9AnE2k4htfuoDX/im1uLDwMb5Q7V60LfUksgk/+zgHEAiDTD+
Tb2NAnbosU3l7oGHWqp93g6/Hu966ofnd8QavBZRM30RlkHB4u6hNg58wOi6V1+9
dY83utKYZjshOCdx03XJGXUjyPCvjT5fG9n0aQLIexa/VMRFGY4iKYcXS/LHVfza
rFiFkdiw6Bq/y6ALOHGwjGJj3HMXdhXTmZ3f/hXH49BKEvYCYCH/ZEq9Kv6+UJSr
lcBUVigJWDRAI/1qrJgh/1NaSUzR25ns/sqTGGjBg8pskxUBvLyhhlKn8jeQMZwe
92fhMNtX9HE4NFclyAJ+y6EqZ96yDN1KT/SnzgkCI5njpOp7FrxJ8QekSHy29zZK
8gE6pkdr4jG/QRyferlL/wtiMh5G92fOzf3Gy+QHjM7xJh5zQ2I+G2b0usMDkUkz
yT/2IjdWUyn/MCcGQQPy9XWRZuH1Nt3z49Fyqu0hI2FFkg/A9e6IEmZT66PoI8AV
vRugBhtPNoHripdpzDcdgVi78IO+14VSvk85uZPG1uZ9yx51+mWiijmOiVQAVvtA
MaZAw0JW5ptr6WkvV7rE6NPyzp+0vXRgX/tvwsfedL+uxEcJNkY+RFC2r39KV3FW
4aEykbFs+Gk6cq3Hd+PEXurA4tL5PlT9aleXLW91nN7JdaUFr2OOO9bezU6edRQ7
ByjsqkoE3LWO7DOG93wb0RlL0MZHiRlconLMxdp/OtmNcrmgNlvvvCHuHcl05tgO
CZ9B/VP1Zs4LLbkLDiHQel8pOAG323kvGNT/mzj6vuv75t43JhqPn85uWIg7Tqn3
Kek8rZfwwtEnuSJ5SJN5ZEVNtzjMyemq3s5JXw5XsDnOnulTcQhEJanBpHXtHvh6
k1pN/VHF3eJG/8Q7KVjobAdK52Lyrn033ANtbyTljtvXb+PeCHrKgu/YgG/A39/A
13KBy+v0mABBphHa0o8xBQbZRXf1zmJCMl30BaB2wveDQkmjg7d1x9iI1LXcAOhR
QeblvGk3x2Tt17mvVkxR1P20kr15u+CiyGMQ6R+g87crr27/vHaeM8mo9W54haeu
s2yA3H+7MNrstLROoaJuEWY0SIdTYBT6sCMtKdMXFwtU7LfC3Tkwr7ecuk+H4FIX
z3OiU5Ezi4CqowhYEpn7sOA3GtrsYUc61yUVuTa16oWmv7InWPp854+gpgxMlZ+A
O3EdxKnWpcjbAx4yOOb8togJyeZUDt1OxfhUKZcjMY+cKLMUBq37uUFpbrloAeH9
EqW44SEzbYI8/sgoA++vyrLxz9Xj0R9aKfz+NVImiBXCn4DZGHWGI7SM0nW89Liw
OrHPCirjD+7zIa/x/u6ofEQIAgxoLCw8oqhxKy3vGhMW1ODlQq3NtYdVlsk/fM98
pfCRcSLRp4pi/8Ei2EysnS0p/knsVWqzpyKAdmB6PnlAKyuCnB3PslBKnisj7NnN
xxoEmXu+kVoXgjChOZufiKs/w/OMQApC2xJrvlrWpNs6xOGHTpaEfmRwA1DnkoPr
8jKYNXljCrxPHx8+pseyYqu+MPuYw+cwhTZT7mkodoTxI2Snk0XnCduKZhM5IVcC
mE070SERjSWHTg9QE+4j5ZfKEkWSsrrfUGyOHfDqUFcYvUjmrh68IyZ4xz4g1HUq
fBSMrl94GSgqr/JaK2UaE5XgeLCCVo159J+DO4wjtXzr+rHtyTxMx2VFfHsa4/0Q
nqrd4j8KIt5WDC0ll+WmAqjehjLSqAOPqypiqv68CE6jG6se5V/+Kf33vg0yNpir
N9Gz7zdcZVBZ+16vAe6GMDR30nefvhnC1Z5z8V7fXB/XsHFHWYZDBT0+sCmzoeVP
dMNL+GWua7CNrMpvdX4xA+keyiG1H3gTqJGc/TT6tml/RAHVa1eku7XN2U76SiX/
zaz9tfzFcg2DufKh8/IUKgBOcOun7V4HcTNFFhfAU6Np47ycpXiGHW0IjZhPGwgY
+s0oRp+LdhjDJkVjeCrvz03p/nlR/2yufB0WHl/nIVumCHjoqF52juGCzLHALw5J
4OhyLVlE6FBslI3tIDmyBRAI6vCwKzO59BaA4cI4ci9gmcycPSWs6fd+RfsGiIDm
hFOnktFgfIBPXlZG6CjlPpqiZG1dSsU/AOFD7XgyJUNS4Zl/S+rTevnrzaUWIj+E
EzPVLampy0cqR6idlIkNLmperrh24glEyP/OCP6ab3OxAmwTbod8EvwNZpYUp5V5
db/k7ZrEYHpxYpSA9pp/+JetXi91dU6Ml98qHSflBHRXsf4fBfWc4xSU3AJkNm9h
+8HhQMocy4etOypdBe8fzusKM1caY8v+k5p6M2OcIgCQCXwjm+38r84DAJ7uxQwL
AEcVCi2LspGk1684RCEgPPDhGtGVqC4+bC0wF1wPijnqGYXsB1awZHLMralaCEgL
fQdKOWatSICpdrHRTtzkDiD0bk/fW1DO4LwTYZnHl9SWpF81ZtK9q99Ym2615wni
wvBiS1SWFi6N1Noh0BD+n1K/iLgLWAA+3sGOUaq5TrSqZQQnZ3l9GceQ+hP8J2kk
mj9Brw7/j8vVVNHKJl4PWiEhS5nx8+ljzhRvH6GtdL2ZHwtycQdaZHKZGBF7Rpuq
aQwIMXlNlVS/y2yORX9ORfn8fDIRD3IH3VCcBxR8bAUSsgJMXQLykRdIF5he27DO
Wie+Q2Hpq/1BB6z873QJJjovZeHJniupB212ZkfysFSgiacz85gOeAZ0of6K8Kg3
sgb5HvEkhfc6bOgrWfEAOHj80PVwynGuYNQSnDL22YvIMCfS1agfjbLwHejllKT6
Q72O5tTX9/HWH8unCWK3Tq63JuUGmNrvj9QisCFYncTpCl5Vtu2OVWj27mb2awiA
3rrDhHWzCV59Xjb0UgYhv06xE60TR4y39ROVFXO99yNCBrFgq1ULM0Pd73oxMfpm
1IJ9VAhHq4dDLdjXsHmevRN8r4teoeBS9NjFN6WQKgf2oIhr6QJumQVTymiIucR2
Oj3Vcvex1t7Jnjni+QOj9ohDVRogRL+5+YYZ+4fPyhHirfhYSboITycSybzzEts4
LP6Wp/4dLR7JLO3oQJJAx1pdYIkXgvur0fa1E1N06OHf+jd4bSiC37ZHNxgIBYrY
PM4o2XuxJuMXldADsrG/VPGlxAgU0XGyvim9hIukGZ1A4ESn8vAXnFQshgtG0e+f
QcXXOczz4G9Vn0I+o5bV671qIZrADmlOirMCXNtbiBs/PSHQif1lD+IJBtjm2VsB
Ev/ApXmVxaNx2+JsDE0ZqD8NpgZ1on7MzMilvJzSr1g6pp+Q4y72wOCkQ4OC7Qf6
mh3yzZ3ONdGa8QD+8I5akF+MaCZYLVkJvbcCPrtUUsZ748Mc9ME2wGtLuM0YsRVT
yXb3GFh58OLRSqk4Gz9pFxz7m36bgSyZLg4ucPtaKmCpm0Os2MaT0+SU7kmK8HTa
Iqoo0hfya5troEC8rCW7FHTruIN9y56yYCfT1pMO6HBqnotrU44I9N5tPnjoYThD
BntuIrzk2iRaA3TPbFIxBwVwzEJFkwy756s8UBiRk7DSV9qbKskLGDol1LAdA/NB
jM7ai7Hb6u2+T7/f6V95I4WxbU9uC/OvRf7ltsVgE9drUQFRHZ5lj9HDiX0eopOo
0HJTLxTfCc5nCfjV7SHyi/JkSLtLBCzig/Xrzmfuk0I/FjUFsoTpE5pfRSHiHOol
17GR1aLE0dMmL5lFVvGesw6yoqS5LWSXLkQIBwyXAHczeIRV5pLLEcpoKlMazXyq
IyjVmbcG3u9c4D3ZDcRlxWZbMCFOUG1XtK4l/A1KtkipeiBC040AKeRMwwJbCfkG
ozIBjhpxaZB17a1GJ9llGugHtxMFT5bgD6gE6WDXdFTTUGqR+zox3LKVn3hU71P0
t1aDmdwIpfZIr4nRHDz5jJNZ3QqSbQXJCdKXEo0ddbGnYmMJCQabPmeSc94WvNrm
UScDwTDKSe/BAMoGQ5NNMNWzBNryR51QOwWHIwS90jMwGdGF/rG21QpQbu0T3BvT
M8SuOSpUlv2oXJCO+iUsNhsi1Jpv/EIsDQIdtcdE+U+WZDYD24V4yeX3a0uzGITt
CFAJ1OxxK2eQSjvTLkwoR8mBa1oYO/a1fZSWf76+yVkgPZl/K2kCbD99oM07ae5F
LQg3s5JDePdMmjjdjXne1L3hP6tgA0HUHsHFEzfOLcixieJQ7fA94qsqXyXxp/xg
kyRuyFldYX1i+q21fyso+HvTsLkHO+HMZ2OM0iP2ufJySngC+F7GM+6bhbRAYRF+
WKGiJy2MgAnoixQwnDGZYth0ynBjwohXbx+VGorsVKEf0VWwhKwOeWL/BkTmNq9/
qO//XVptsiLFgguy1VUuhjAj0RFONtsPnZUrtfeNMTpv5Wmec+9ikw3KEj6dJan6
AoJUSsFMxpPrVIXId4heHZtmI7gGflN92FuFHfLTAIXFjS5wMmxAy7e0yqYwKn9T
XuBPdSZmFjCCOJ1RtW0jPaQD7vDHSHsCZOGSpFtuRV+++MmR8lu84sdGl1sgkrTe
ESlqDR5TDZiehlQCOImHNK7MYqo5Hvrt30CG0gWNrQa9CNxbFQBN3O2l2X4NHeCY
1+DQCoa254ox95Hc1G1h9quXQxMx5yhplK9lfvFvh5svblA7pwqUuoBqETrh1+sQ
/041cRzTw4ZD8feh4UpVUJmU9wzj7Xv24A6tJsAzd1PEVaRIYii/31eBwmoq/L9b
k2pYoWygwJVc1g7/BJHLftA0oiu1ZVH3Z1FU0bMxz5NHJTj0i+zkogJfO7agt7zr
Gx1V2vO1+ur+u9eb17a/tJyVgl+1y2v0nyrPn6D3KxguXCQaZWTXVjMK27ZdjWMz
Jy2MaWxAJ40ctzJFTW/Z/u0/+b/TPRFkxCJybKIzumzUd5UU1aIvKmshzYaeUZrE
xmZ6rUKAVtEJEcLezd+DJiXOIYVknoxwv0RbrTpJ1zCwM3DlYebKdGiFl0imPYBJ
VM1b/0iJfF391/i73O7hqKEpiWMKRBIWtb6DmlMtjO/RkqZmtsl6HCW03sxQbbsB
Y9piwEaSG8kM/WgFGktSbSGCx7Eyw/s09duKlp0CpbOU2kyZvYNvAicrjSQ3RMZs
aba0bHgH9KtM9mkkXP6da7Qu8eaDcbdXcvPNviSOpLbnCvEBmHX9YyuHS6f7Wdt7
h5hTgwT3TX5KfCwUdRU+oSw7yBsdntT3gebPX6umLBRNeD4UEtZdhLAuKhE4Phm8
r5dbGWqQ/xbOSxqZwc4qQ4blu5Cu0FASe0Qfcn7XfhqhmPXsWFnUvwAaGrbwDvj2
eU0h7sxNNjbdtKN7/ezdX1SKiNsGuwO71NAHIpzarxEbOBj+8KQEGZe++ppRvH66
ummlon/928qt9wQ2CN8E8dRsqDwfTSbJdwKcmH0NQQPSsbHkm6HZYiwPxQJ+UowC
CrP/OE1N3l13Bbg8NPrAIo+MZ4RPr3fnRfkyaC52qAAPo7B3a+zTNn439Gs4eSiM
HXVzau3YYfyzOLCc7x8IZuz2byikgIg1pl5dPRZqWNEbL4i0C265WUaQqLu9sszQ
H5gq0yADf0oME9I2OXEn1CiSLuLDX7Maex7vXXNPakXefvJqdXgRwBpskUJKQHcr
rfiLF5Jl28HtEQmIKFpHBCY96ssLrpfNOXqCUgQ4a1my8WkhzCehxzakYwYXeEgn
VSkdxCf3JUYJNW0NBDRsefmPzgeLrebieh/9kKXGDbCG27huNUgaGhciZVS9Qavv
rg+WeO1oIMkJwd539LuIoTuSoCT83+ftyiRa61mKWsxOM5Dn+SGwdub0KUiJJbEZ
58nincddJkvpY379aZXAD2kEdp6UzGiLWvqH8iiEd9q9ro4e6FkWh5RVCgrvZ1zR
5gd2yRLjKjcKZIOkoH49dM4hJCpSiN1rmCpzVSATjmhxkkx/TF4SiIPn48YNNTCM
zOBzPIMckkHGs+hVR4xEMWOSk55WCZS3P6Y3z5ZVJTRM8xOjp+IRxRg1/sRNKVjX
PW4mjaUPzCUVx6cyPNcjS5YckByyWKCa/eDl/a1JVyzKfMubyLSbzJV4UxYSharZ
l6jj158QQC54nyubD0q54nviNjw3litP56ekOLXaS1+N+obJF+X7eGO+mIsUXfU+
ykHMmVo7fT9cg5+aGBVq67pzkC7DptyR3P2QJqn4Tp6UB/XwxHOrvrJevxfH2s8+
5RV+n4cX9pOBHnq28LH7ZpLbQl2m7OEsfFFSqXx/AE8UFkujayh7xKDn7fAsxxfO
LZBZmYunu5441VYwiHGeOtbKBmxOoKgyYQ5V3b1Kr99OY77vrkpjIxGggtlMJmH6
oVphKIRXTGgn1ep5AwjMeqdJ9UdClxe15zxOusP+xM/DGzkjpnIqEc4ksrp5b7qd
D5lC0CRv3NyK/ue+NY/pHi4vMO+RmZ0Rgo2lCRpu59PrPXv7qSBOzdpM8eAI1uuZ
VzfBHHLhA8jLppDr5w/0R+rs2dzmvGNK9zIpClMYb8yhS8ClgRlNjiGAx9/4wVqn
FEZ8dr+WMQs8Jciwr4VXNpsISGkV9gEj14vch32qSA0CkqNrjaQh9k77Rrw/jE7l
jZX6h0EEdomlCqFFDUU5RS/uspMimnG1KgyK0161bXbhwTQBExiAzGQR61PC0M6r
TZnekerXKEpx2SgiV3Gq/YuhcegmL0ePufoV0OdLD1uW8/S4L9F/cyp0OsXpSywB
q/oKCJh0vAK0pdVxy6Fdabsb2/DBi07mo6GXGbRYSinJKqxeYwAo/68aMNIA0OuE
29YzM8BYojXW8l59QA2nV0/RlQ5ag63iK1ePi1rLGRLCbq5N4JUkZWXEwEumPmJW
qfLp8K3ux605l/R/cMSCDFx01apiAfj3BRTSusVrtVyEJY7pgwcFa89zTGgdcu9C
+5hH2E0oo+f6+/xF4itLCp5opbVojVGxSuNpzKYdARbVZcnHrT3NQQ8Gyp49CY01
PI5m/1LX137rTRzQN1W9EvROMH9JKrLY5TbAwpjkSDJjYmsNR8t9OfCG08vlb0Eb
UxJe075h+EY6vS2OeB9C4rS2WsF9RZLPXCK675rzDkZnzAx+uCqvDmWQcd5EgoIB
S/biOowUe8f7AtgjZO2NxhpcuuVGBGT8SpVPdQfqpX7UkxUoeK4VDiNED5yJQ41j
QiKeOtkjb9V6ptQsaS4PZ9y41NGSEOpG2TuEFjQJ34zKtbcmDrEJVSCtNV922jTK
X0b8cdxGyJq70kg6HxPFNgjXLAFZf1ImSW12cEdbIb4t9Xzw76ORTMmpLcWQguo0
+xzcJRHrqc8FTrz7Zw0q9Ptd0LjorLT2kb88Jro8Yb2y48gtUQoQRz8kkgA547mk
GTIx3vgPotAI1GcCip/kJzJDkgacmWCCA6gnCYwDIFw8KgvoR/sOHYeffHuVwrBg
ZmGBsIOTs9ui9ahE4579w1y64YqfF8xXBNm25ogcXm35hfcWgF2RKrOmuSdtQLRy
VkQ+5h4JjM/0f0PSneQKjdoaqjvCBUP3EKvYsY2hjKqX+vKbVEuU+gqIc23bgdlE
Jac4c57tB5ijgrI3UcRNQvFLV2eomujvWr58NYplgChTjOIUldoeNTun61K6cKT/
TKLHGejs+d2h8KJKuvTt1bImth//8dw+demEprcacRUaV63eNqG/UFolYK1LZlj1
kBp1HAQIqlOYThCIfiV3kFIeLSZq72dis/6DkwAoqz3/twMNHDE8lKwDGleMhLQs
gO7Q6njcP0+8shLcvwEYQQWibP7elc6QWNdrXNClezmNBvYjy+gr9icyFLZXC45E
ulVJQXUmwNefqZyv0WIs6ytAoOBp/9vnvZcC/QbYLClCPWcLhW12xqTiPB6YJcNG
kKACz9g+nNygJeQfT5OR9xN0Vcqo9PYmtbbKyosas5GUjfYj+Bf/GVBSCPs/mFOW
WwzlfLQnDebB0ltKwV1p/Nn9eSwjmEk7ydzwccLlT0pDURUdstmawdi9ZRRWmaQv
bSlEUcLEFVmUaYzMA5//4KmVTyf4+dlf0vQHbLlvL1LtVt6jI866d2gTT6YN+y5z
zH+JRdRt4OkFY8fJJP7Ebt6bhEja0NJmFbrkrbMJOD2VYHKT9MsVO7vO+/KL65u5
48uAfiadFkSHDGsz5PtquL6b2cFcUU1JH+T1zgY9RMjRv/XTZA5t+bwVXZWxapCd
bHtlygNTkCmIONUyJpoxKeSfyn1tnOXhWzA58c/+s/sYDPCIbN/qweAHGZ7wmAqH
VBkyFy9fWSCQaaiOzyQ4/H4f56Ewy0cETbsQfjk8IWxvPPSqO8BmpJmg6R/pgjBt
YSZkX60JDR7Y0NZfCSwQEeua5gU1+kLaWOXge4QPoCBTSQCNnzGstgEmVAB8nx8n
/IC5UYghCIC6dXbjK8i+qJI0bjxmW9tvAGxQIM5g7oPEtOG94bUVKb+iauMAY4Ww
TjCql/djMEAL9+okqhdGGmIRSdnwpPDpeZ+6snk+MfEGWHSwyRHYa/uMzUwGIrww
ZBODU7rrJeMKEdfQo7osvNN9dIHVhQO9XM2TsNpUBg2GW8YHZPNZVzyK1pJ+2ajy
APOhDGsNjjY/KgLyj//k1kC/Cq7XLg+e+Voe42FPzqKT1zoj4gybG5tMm8CyV2Yg
NnNIw83BmlGNveU00tjSGH7cQ1Y0UY9Hr3iogwxCWt8HrkN60/7oPatLlSLVsEip
Q6FmvB4LvElJuc7+BZzJxZm4WseQip77CBddNxuNNJR8dB/mHy4VKM5nrd50QXYR
CDHGE1mbsjgDkCdAdjhc9Oyk7ttaVkcpHUh9L3o+Mz82hpqjszLDkS1NsFzTH/J0
b15joM4n3ZQQRT7duA2acuoevxPCiPavA+GBws0UaxIkEAqnaAmtewSOGY5J7yrk
RHUHJfpo981TYoL0eKdZeesro3pMjsRVnbUjxZfmVR/vYDUOOmBABCTOsZQxbORH
DX0HI4R1Sv/SdzRQryv7WbsXpCZDQhoOr/6Zu5A5ehuO1rLwp4VlMpO4GHTs3Q8t
F5gDyw7+IFHLDQZH4AwO24HXC1oOWFf0yuBF5HPAUg7/jRGcGcnMH/CGW5u1r8BB
JTQBMfHRp8gdivX/faSd+BpqxVXwtdkVGq4At8a2SI4vgx5Yzqd5xqNVDNZVQBZ8
/wXLCLqjPIyidjf4YWQFU381wFzlivOEXwVIlMbYygYlZnHuyZrIcZc0LyWZDkSI
0k/JmErK14bly1vWQTRM20NIMsh7WiTiWZzEmdBwBZCQJWH1tuVAKgn4vF/5MXSr
WTXGHwzkS8gGwURdqv8uGKpIFjr3kO7k/lNwUPMaPOont71UIqEMpPtkr+aYzKZZ
/PYl5ojI+JkGQwrxhNqR0uhcWhOvKLKOedYZpr4qdmD1Gv3pK6wetPftC+lFz/I4
0ZnQZZQ1PAej3bFph0WDOBglrUCRz7bhEI+u5blqu/Qr61JuovXQwAwe7+XCnoUw
2YEBYzr+BYRALVKnHpRbRTpVdctjYFAFbnK0f5D7jhhAo2gshoxXihfKaf0rc2wl
hdHE3mp+LGcnjJo6dj17LhQlN1YpmhinJLOwsrV0BG37oBAIOitOIgUfJQD7oCqE
xySaYcuU3rRa2E/PEme3a7unoRQI8nkNyRhzwfVUnfyOdoEmWgew0KaFzkpO5Py9
r8Mr+yAzagpp3E08bEbN2Jk8ehDitPAF55n2ngwtJkDVGA9x6RgKkHZ9XACF4pxV
R3BFn/i8f3cSZ80JiE9g//plRMN0N77GuOk/c/lP4Md62edYxCtyNsmPCx2jHt3Q
BR4VviBiWdNOIzu1kAJ1p3S6f+rL6j46QRusRQWTjYR9ikjAwyLxJ6BvkVafYNfQ
VhCrQUA7gBT3c90t/MPIG4A9uFqcNusKMz9eyt/FSRFDasf7DxnG3ImAd5YkLdCL
L3hIc8F0WM0d2t7uGgmqsyC9KMKgrr//cI1zzSh54Thqouu3kHsPOvalFdyVCISk
tJ2bFt7h1/cDwEz+S4U3KaTDKEvFcTImFzDT95rdjuunHxgP7mQj/DYzDdsQ9C/A
5zDTOCR9A6qek40Npqb5rXit13wDAHfWHx4e3uyNwp1oNh39g5amehMYMClEQ43D
2wX2PhCkhxmMsJ994anWW6sX+8kI56R3iNCgZRf3D4mMtpMbTpx5Zkq4LsXcZb/z
78M5wVy0dFcXaB43jBmovwVhW0TuGCQV3ai/LNPbBQLiQFXyixN5Ns4m/jujH+MC
xcMnzG+pHP6ZAQVuG8ANTDGlAaEpXOXQiDzbnuIW4UZm/PpDn+IK8qgcf1a7hqzx
KXV2k2cU/ldm61o+D6/AqcHRVpr7DMtB0qugzqtPAQv9lv9mDbYwMc3wAVg1dVaU
xRLDrmNmSJR2QRtSom8L9flf0qdeJj+g48W3ZVTD6Gf/k6x9c+Au4I1akiWExENK
D6e7h6FMI8/FE+ULbCjufZzU7UxBuo8LaabpRcYA6+BwMbZEyM3q/N/g2jUedNIF
LSq2ug37fv2a2YkVqlv3f9tqLuNHvViVTcMUkJdZ2Pf4/szA7YwLAmPxlJdH2O9Q
WrE8yhBYHeDo487EKflcm5q66gSt96CTClfORbATfV8cdyH0EFymfgnNVZdJ4Jen
lt8pHufYihY6p+N4LYtfx607PMvfxmLB5INDdBtz4ejDr8x6nn+TbbZr2MNUyO8/
JrQ2Oymd6zjUpGuwv2c898YJ8dK/CivPSdz5H2Q04D3Jryg0dCJwZlmc3QveXz/r
Xty/7TyUigmHRZhUOAGhnQynUnjnpyuGrZUNb9yv8Hc4RX0aLt0pqoGPO+uMpHcj
5Tl+jFAN/DISsYJ9cJqN0lXiehBxk54hhT0fgyQZnr1DksfbhXBAh8/dkmfT++7k
TUofwshrp5gDIKjj9g7mtyO1Hklc5FolrEZsYu4GFUmpOBNIQBxgl0lv0PKWYBtR
Vi2X3GURfcA2vxaiAlaO6EeLKbaE94O5N0WKpSm4BrMrZ0cOgvj9W53HDhIMN0pD
XkBHH6hEKnDpYWSm5S3hrn8qHMXFo8Cy/i5E12KSXMKcxSAjSzH6cTHLqc6m1cA/
wv0TGj/gvr8dw0KiF9i8VXcrbxxXbFhdp/+KdcbsQeUdp//+BllWEQc0aAQuIHRw
ye77W1tDp2aY4GqVSargq5YY6qZ9IGB6wc4Qy5NzYFcpK73CUdhsrPWgqj8mEN+X
pcmG3MQVVW3qVn9EdwT6NyK79CA6NlmXnnhebsJi4yMJj0LbmjjOpEKbqx7v0vCF
w7gOce/w/TAh2Qz7Urpk9XS38YNOkaRVRzU8CnlyoPBfHb2JiTVDWHGIcaq0I5QX
59efS5h/aQgBLNpxFMIN+MMwKPJgw9FK3iwbB+ETWKa/66kkJz40k8P9trDuQc/D
sO92OChLW8mQe5B4CrrI+qAqmi9S3ZIDYF9o8UzjlhAjuDgveJJRHlx9zJwStbFq
JsrJ9b5YoiCv6Ud2a5LTy5HwDLnyDdTEQeXBnrb/Efaq5Fz6H4U7uG21358CW3PR
wPusTNHJKMsr0QmWupw/hz3HYCysS1kJx7GEpCS2h4UxZc0V7kl//faIUL2NzlnU
9TZRfdwGQlNk0FSXkyuBlhN8fbF7Rp4pt0k+LwplIYVSh+3aRqBy0gB9ceEC4OO6
tMKSxT7omMSWH3TRESeGvK+dASSitVLqmsHd+Y6pBcjG5v7BgaSkEEcC0xzMFPcl
8cUil5kXSNtF11Sce87ji6vq1UtRniMa1iazdT/Da1rUnE+Qexh+JDC0bbBiAh6K
xPuRVbn4sQMsu9y4P5fqBgS/KE/e+C+FhH+LwX/197KUNdff9KTqbY7zvlgk/2fL
htraCVsNvh+zJYT3LlRJEUwQIEixayJ+XISZWIAb3MQNvvx6t+Y/MhnPzWT4nohI
W2xIrGZvvdqukhFrlx6LeTWqvK9cpZ1EcpMIxPrwJ0BnliMKgQOP/NXoT6IlBjVA
LA+c6GTSw47glQ0hs2IdGqatBcd0CH5RHktUp39h3lHKbIs9VpFegka16ZsEIaRn
lcpJkI7/nL30vGjeTn2SRd9fGc6F99tNL2XwH7HjOAGFXTG7d/M0Ir+Ax2Wnz1hC
BLRGF10KufcGFqHcejQAR7Fu+R/GrYNGQRm/WAAcoWzqy+o1Li4tA2CDeDOTx5UW
PXfpqN/h5kFrGfMbGMbURRCABlwL/KaCPLAYA+VT5b7AFu9eZsMnJzm7F6rRRd+H
u1Fj5AgPqU6zbB1u1fhl3ee/dlBEBzOPyiVXO/cnhw5LHcoMLxefFW4E57yfM/fo
Z83+igqkP5Fbn1wAC9q1Rs6pmXSl9i2xZj30geWK369aLE25yK9W6TGdhdTrvSo8
UOWZnaYrqFQ1K30+FaeQsLhzNNrjt/FPvPy3jBdrJiPe6WaAbfiWJ465vHU2ILKM
c901NHjCHgmi4/kE/2ZuKCI28OXGg60wppoPSIAI2UPJ8MG3R3LxydoJc20W08f+
riLrp2OM3HrV24xbZJY86wYIgS2rXmltS9cgq3mRg1I/kJpDm8GoAntJsbVzX/+H
X9av2DjIIIBw62Xu/Jjx42nTd9fx8E6l0FgY7zOOK1FCWWFHEcQUUJiIa/tuUvqc
+bbf2HSW4a5M35RUcWFsWex+el01Ha7fwzU3CfCntotOcM2upy6mHQUS6Yui9MKj
VJ0O8t/zifFSJNX0ec4gDHXJAzWesAw9qpy4SEBfxsW5CI23rrpQXjSh6cYHYWuP
u9F2eIECs72qrhm6WO9URkO8kgidWCKMqSSocO2+KUzsa84MSb/PreURAZes+4Ak
0IS/li6VT+EeRNLTNhWnPNYR9AGwWxOYFacnsFJAdS9xkJGrMA1LQz/HRr/g8xKJ
HqSukHZprNmaVWqxHEv8U3XruTPm1pK+J+1w1st/DPQHTxhz69/JeJ/ayzHBGujI
ZRQXKCkII7gpcz/zNOVInhwhyjJCG8gOBIqvvtlQlrAdrFBpEDThTohDIOrdnE3N
OPrt1PveBiGTOIQ6axt12SWnzvyltlXQjr87fKsvU56eiqtVDQ3Kp13o0TgWp/EK
MlkecUgDxCpDyB8m3Ej2wzFKu0hVAhfjfFFduK6yRWHtW4C0UkV1SN40ceIVzF8C
gk6HsIxpUwMEPl7eem1koxoFXWImcKvrQvcb8BY/rdKr+kAvcRYuRTkwCSkoarnW
dHytf3kgEAGlc7zquVTp1yYNtMyBGdTiTy0M3ymK9dvn7QcX9XS2iE8l1eswsG5l
I++Yt0eI0qKSH/91F+E4KIhU8IwfkqxzsXWFdih2Lj0uOcPtee3a33xvS1wvueR6
dQegCX+j7CrlrCdd2/7jHoK2/8eZuACdZeYf0l9c+P0j94BwOw7Kzt834lTXxSQq
spKhhVIjLH7qeVCggyo09MQLbLe8WNoe2jYyxmu3QsvhF4vjDLK+cA13Ei58QpYN
pPNjjI87vjpn0YzvkzrCT6Wu2Wrqw72QA0HFBr8DuNiotrUgl1lGubR6UFV+siOy
eCOvIhGFsfUEHrMJRVlPIVvFepZYFkEaOw/TvOZ6aG11KyEfnR1ITPZuYJNS/JQZ
/uUxdwg4TAZBHbmoN+6+xMpitMWibFnZ/4E20oDGv3eueU3aH5iXNulhCXf2Swsx
wvfLUPjl8GrpjPVkjUrvYtQmBn/ZwD8n7IMuoKm+0V6IxhD/KHCKUoCrStRT5yfv
2K99iWtyaPfnKokCumjqW56wBavxG2CGUv8lvqmpNKAsmXMm52USe1aE+rtJZ1Uk
R/xN3nJeZn9SBlFSUhFE23zaiZBMM+hRNoLlrdnlyxkbsgOgGRysMJxJnJ1h7EG7
+1VXACUTuV8sTDZsbxzn1Lkpal/WIgR2DjggxAL4aYqfUlVrh9Iuih/Y1KOjle4Z
sGkcGczTeZd+IPFhUTfTvKjxZW1RYQWA8ZM7jo4apNafG7818YBbrs6J0cYi0j7X
bwnDSUBy6B8CruyBh1ttRI9VloEtAhsfVNf7SN9QnSxV+yV4/8riE8UzbKU0u9R3
81dPJZvQSnMxzHPUp5w7uXbTPol7L2zIusWPX1kzjOb2nZLA4XI20L6xdi4URwcR
d9cvL7vB6mnqJnrymR49iQc+7rbSQ3dAlDoZUFXWpB/0T+ZY2XG/+SaC2uYAMqV5
RZXFuFowQI14gcwWWa2dBT2olIGZ5QsZ3s1MWfRkWD5muQEe8AoogWUfAfyGSgs+
z9KGZnZrEaT1XCAywtKNoueyfFH790xIY8KehQ7HMFmK5UAdE8ShPYYeUp52pf1m
JhJqTXn/gjwXHgT6w8r3b84w+NwY1SaG7Zc/J1gUd+6P18eXP2vrXJCCl3Qtg0H1
1+79/9UVWGuT7Ajhpkrk9PUfFslVrL7EqiwtkyMcm6mZXJ27npJNVRujgUKrQj8h
bXBsfQZLFZQdMbmt71UZcakvhRZFr/wv4FmY8bVj8N42uRMiV20oevqR6KZt0iBo
ASBS5XBbX7/jfRiPRp5N5smZUlBwD72TTFdnFcn5etpMmWziKUV6SpJfyvCDOQ0v
NqmFNuicQKB39d2UHqGB9eemkpJopBfr36TZ9W0QzewCrawLOgomCZu1hzGUU18+
6WL4DZe6hfecuVTMIDoA7mK/S/PjE3Et7VpShKqu1oqs6sYHO7hwvKV/T8LSStbm
0GNApKrTggb2IsKBPNA6S9TxaALp5n2wPfgsuOYma4lZjuS/xdXwhCArkioFfEfC
jQMaXFwyg+seamtE66ZMmxFO9FXpbA3XKb3ZTrfyq6eWgCdgUkfxoer0KSoqATxh
tL3XpfCmtW95ImcFzyhnFHDZaurlnxPBxJupHLvzQbHZf3e/0k5n/9FLSjZ+2fYU
UmGOEtj5nqF+jWjxaEG6f/i33KnLvoFMOMRRJsjBPn0wVSn+ukH616Y4GHVChXhE
8+vR7PAQ0uPONuXZ+u7TprRWudRo1GGGGomCiYe5r26QpeX9fU2zdEBIuudE1B7A
wYt4MlV/PpP3u1pKTPYoWAKpFFUUspSVyVX7X8sMs1oAh0jI6SinYngsFT0RB5RZ
x8qx+kF9gs/Dkm1sAi4WOaydOZGwJGInAyWY83TXqWDatC1Cmm/z/1ahKq7thjST
xw0sRD4VOa4S5XKmtjCDHkUnK9RhWJtPee+jB3TGuZgMoUNyJObLo3IkK8cPbEdC
JAmF9vJtRiLDzCMjgUpgeoLdqkVijkMOKHliAnU1vSet9ItKcUDAJbmdaOOz/jsB
qcdV8TErQN0RcUUa/YTz3M/giuZLgEfXgM65z5I2lTaHypnWK/FuRAVEHpCj7YYK
7mX7osV2L33dfoD12KNkcgnNn/Mqk0W9Kx9nmCYDmP2nStuDsOjT4U6gGrucf3LA
Gnf9fqbd7udd3lHGIN4gkmvRDrxsaFdXa15LQ4epew4RN/kAb8Ioshps6sDGAIGe
dX9srRs0e4Gr/g3tOuYxXKwXEB8FmgnDtWdqCI5xwdSRV2vm7NYCHW/TPyI4ejy8
mfsldEVTtJQTfMGPfX8J4arCp8pofEQTzjw+sTaL4Ev9xRsa7mVOe4nrYU42tl+E
slXvEiEfYPxQLLAVnSDHo+4ir3PP8sXf6nZtpIR8sAhex3JXe3cwqNTsYevmh5Ub
g2MXVnSW22rZDbtzSdX25msTOoiE6fplLFh7nI0ynGFdbmQ/vERfTFF5MQ+Vb0oI
ZNjmZmcb25aHXMPRvRlRJGnXtY8f1wr4M34HbrOIwkNLRYB4WmJxzRkCR7IdcWNA
2YC6iRZ6RPBd7W12paX6rzqk1xdTt/MS+kkUtVHLkLJHikuizuiz8WiK4dMd3rN+
K0BuuLwYHcG9RP7grsZ2hd9bCe4Hi0Mp2r0ipXvlyZocQvXT/IMGFc3uHJDAtQJx
a2UeqdIwRbskyRUf7tPeW1CPN6OL+R7e6cfFMQK+cxZzaRQGxYU3Y51SVRsQIY+b
UCndCEnRzbw7GhsUrWeB33WabtkK5t3/y/8S4p5mukxdMLZQMg79Q4tgk8279c54
SK3LQqq2unQFioGOi4MPz8fB2LyxBs6DNPyB8K+ctNGRy3NvyT0d9CswCSUMm6jv
vRjv9RiAOR74vj8ihdOtC+/vdj0X1pjmn3uaudQTjNS+J0mJJ8bXTmQawoY0zgKq
xpwk9Ae0cY3phFuEjO8Ow6O6hf4UPrfCd7JMkmsLuFLou9KnbkjRmNzYSQDP/gLI
G9YhR2YFWhs6okyyCd1GZpStiV0U3eOvQuh8QqllBY0qZvwf+yNBQIJhl/nMGm90
AlLAE8+OATWkaNL7LpMiPLVKneB9/fPXIVCmVMxQY9P8/mo/ZkdhqPA6hzUF3wK0
M/wJtwY939Qn2r3Wdh6r56GL5irvUTmlWHOyzS8QdWQhyUYvTaZFx7vPXitO1F7+
1NavHJfsI2A51b2MGxoX3QQhN/i2zcHn33MYrzphdUxvwKA7U5tMag8hjrdsxP0s
MocxdL0/NdZ/qnXwGxLA5+KS+Me6BYl0qmgei5D1Y4Wzo86Z9nU65bCf8cgn6urb
3DNnXizSN6DqFnVoWkZaKdkDUBemjGAHXkn94LeXoOXg7Pms+1QXRq9MLV7VisVb
AN60Kgt1XLtf4ePM3txC4lBnewxLL5xgSEhRdd5RvVp/SlhcZ0Yjrg7t/u+BtUPx
b4BvicdEKaaluU7krxZpqe14wWVrK7aTwmUa4ax8p/QvsybzOPm+aKe9pffy3GLl
YeYuMp9fskRMODk6tfzAqlQv+ARE5owJE3zhBf8jg+rDa6gfTzc+vO2htP4xUiEU
02SATcZaSmGWzurzrwN5exNNqOgVfyL8iwJ+OJWG4biUFV1hlI/DWgXfN1ctQ7Om
0muMyiuuIpmJY3/3dbFNDUSwUEjIN2MhiFwNqYH8xldWFweN/wG/TdkRVPLANkE6
4lf6XnrdJj9mofhB9fjN/f62BJxsK4Q6eEFNl4UJ4YJGHTiXgX2cTAYbjzbTJl/Z
8ltvZuNxeLMRm8DXW/0i5hZSm5xLS+7Y+Y5LJad5NAK1NnXNOg1nN3W0a+HYtRl1
3tmLqBkObQUrkGNeBF18zyRlF/Lk0jxS6uguXjQoH80X67qKyZfR1Ytl1K/dRkrc
C/edLNPuFLBzwEV5ACofFHML8JDGsYw7ilDVzFCaCkUl8wCgTKJQdxvVC3wutr8v
Z6Gv5pYvakPKM871IG6r65x0LmiAom/15bN26ZDjBRA8BVI5tlfqdAxmQpp5MDzE
W91XUO9QLvciKtxCUHf8/sOQSC+6ZsgVpLJn/sQtvm/VjfhuJFm7xc2yXTSl6VBi
lXuFv7llaZwpUoTD3cmA0ZiH+Jqyn9uJogUr3N47ItEnHLxRWiA/6uprdKqwnvv7
eXLxOiTxwhokiznSEhN5N2BD83DrE5tJjsdgkE+ou4tllhwyU3+S+5EENayiLT6w
c0hr2AYgumkKmR07d1gNn3aB+0Qc5LdYagzQrVgPO28okPlr0cK5duurRTtGL6Hv
I6VVsKZ0Da6C4aE84WPnRAlRvCDpeK4Jsl2Oh6xc/mxFGiV7KpZL5QsMe0NZzjlF
jx3o7ISxzB4aH+aMjxX5zAUjBkQy2Xps28xGURDaP0gWF96kf27/P50pgC7s/qdS
25bG3BxYBU8kpoa3DrqBeLlLTm5E5fm5Iy4PDozoxkU3jVdC09GH4wHlyUdd81o0
1w2jOUVKjjp5YNyqvWO5UFQ1RNX6UM/NaYbpoXCVA4dwH3zCKQq7npUgYqGxKaJa
LBZmcHhbroCKuelNh8vb1fJFSPK2daDBYdFp/WuuIEzvWMUrWJP5pw//SVtBF+W3
Veto1mnLxYropTcVNOug1hcYWBcXVaW1Y3CEDKT2O4PLctMCTCI3c1SXm8JkgJRT
MoibrQ1VPrpAeFIluchCXlP6G51gLWOh4uGMVdq5B7DCde9tNLI+lHnUmVSazPqX
zcFh2OQwB9o2hE7Cq2j1eelYYWece0XSM7bIGIuEFKcJlTeEPBdapeNGOiuv4prS
N01SZtbx8OYc7NVYkmD4tiO3zrWRF0eb5IafmtGPeToDGGuCa4Ai5vA0GsqZME95
q8QmFo7/5TxUKdlBKeEDtbPum1S1Bt0mDSbdSxvdl1uNu6QgLu3tpgVXF/PlaBeq
zoWfLg9hO4wKGVE2E/rTN0FrjICMbXBqJPVnZdQmq+95QGGkYkdzk7O9/g/wJb58
z8Z9X/0fgJbrimWhUsFRb0nNuUBwYqFc3MVONFO3pzii9WI4CTsmGM0PHohsbcsS
J39IEaZQbzZ4vPe4/AAHE4+z/bhdXmLOoumRtB0kQGzLYbm/O/bPibpvdPocN2fj
BBqwz85dm/bax0LI62MDk7GOxn90e9Vzm9mDpJ0uGTQqNYoR1MuIC/2nRJDlg5V0
5Nb6creimKRwwc5oNsc7Rnj0JKIdhwv+PX9jParRa/zwyPhXjf69OZjChLnL8eAK
dSOSeI9w3d3EG1dWoEI1XedCRpVooeGGrnOi5PxKtMTaAAuJ1Ezb2T+1IO4HWRt7
L4IU9r2qT4UvjOsiYWaMatTsXISPTgwta3EiAUDGWMYd7aPvflFtseP208cW3Dnu
AKwzqF44nO9ywrEejzjBoD6913Mtcz9NWt6KQqA16KHt3o1dURM5VCLEVdWfYYTS
j1bSSFX6yUatC2KJYlkp6D9ltnF37GNypGncaDrkTxOlnuKr02gysYsE3cQVX1FJ
4QhvMJBHCzAdawaEuXmB/6D64UuyekXGmevxnzhQfdGJUaB9MxLcHC9zI+LQ4n/y
MaNsa7CrOibyp7M/JDl81BOFT+lMkRehWym1XGfjKPNvwZe4akPodVZAA5YG/6wZ
ZbqHiFa5gI56JZsm4ilDpzv3uhvW+QaQ+FCMbx4ufMx7gmLfEZc9SvuwU1Rof28K
lwfutc/z5Ysy8C+R5EmQd96YpGPk8GkalQEI9KXEnq8nQGEAjbCoJwYcv/fVLUis
Q0+LgilpNrarZT7eukJ9aqG7i2VHpoM/NDqWMFIXhvK60vU+5Mvo5Sa6A5j1Nqwx
+Z10eGYAolDy8XOYi4kBNhTmxKun1/b09PpqUhdo8b6lao3DWF7pKoZ7Rc6PlPq4
Di4yKhwfG032KOXOtKD9MJCWHPf60miMm3p679O8+UtCUQvSomXnvARfBqK/fWSO
dx4i1VwMki4tfUjPNnde0TeaTk5FXSMBkLkD2sngGuD4E0nKzr6dbH7Qn32/xtVe
yjL2+s9Knyxll+MDdcXalJeAFZPEJAWi9OjZlaVZr/TBoNnd8ihTEEXyb0nzFQMG
xRvxvYj3ZJ9zN2jToozfiIlGTKqFFJGlI5bjsJiw9F2LP8LTGp0I0QQKFWJeytLd
eTiv2K//abi+Napj+fvD+mz743c/STn8fvmam4/PGlppEGp/I7vWppzUvgg9P4o9
CfWhQ/1f029cOkXZTMDMQiL+lm/jiE4YRLyV6NuxRUA1/MHIoWCn0UFc3QTFNZ82
X+oiNV0M0+63I1qQx0afBov0TyPSdjKq9JLk/bk66qp+iWJvx2LChHwHu20Yps7L
WXTs0JDntXegUYFb4JAXRgOYsiCoa3hodtsp+veWCUChLIM5U/N2pC1gAwJ4r4EE
a+W71Z8u7Yc4X8SbnP0vBi4m5p9prdYSOB68FL766seBJRuq/aDMl34bzFL7oadJ
5/HZajkZEOfgP/7FA5p3JXaCHKYl3qUgi70FOTFqCH9oX9id/4Ba3LKrx8COAYo+
N7VJvGkJJGsvNa5Qx6EMVfHNdPWkRBJTrQl64xKPA2yO63uiNZqvOg+T+WgEWav1
kqmS2fUMK0DNvRmmGBZ1zzUYBO19C8cilbB78/by/EpKy8KYEy/HQchkFtd1oAWu
GjeORKb49usuhva6KvLh50IZpQ9cc2xZUQveP1thJTFMvIvuYfMb7OKNCGgezuKe
atH8j1SMeAwBMl2ILJ8Coz96xufbh+UW0Z6jlaFQ6dHySClMHgaJWj4G9NV6vG/+
r8j7IYVMdwGMN+81+zJkQvWzmxhrboc9DvpuBJAx5uBGzv7GOlFhUxbZ3vmFptrN
90qQBx4nwNBQbClau9nLMRyIlyi+1ht1osFiKeKFffTSKstBZ2tMpdhDfDloCLb9
cFix6oErfSFaD3DgJfDWAktEP1vFFtia0P03q2hZYJouIwuNCH4zOSagLIWo1D73
hhroki1ELDNhyXXJvjCke8wUJ3YdbKEL+bex4vAiKL1XzWb6tmn29dssxOirVtAv
A1vbEUpXfCcE7gkynWDMz2wewe0K3X/UfpzI98IB7sbw9iSo34CdsQwBRkivNqEZ
wj37ib7A40o15jLLrfewmcIstOp4eUdjDJAHrQZZE9aX8W8m8BqcT+6IvPbPa3Ky
ybPmMY63BHfuB68pqXDauWqVzNEN00N3oelAgx91mbDBdQ/a0uI3bowo7F6rtYKY
ZWr/g1iInWMN7aTKw9TpyO9/jwWbku0HjqPhXMzlV8FCk8xAVlZAW7t29pTIVfNp
cKIyiTxZyG7VPuu3k/XR9VvnWbuPjy/tNQTIs/SqyCvMV9Y7Ew4n7vAz31QY7LMB
D4nx0DDu8AdMoWdkW5+rIY7RXNikapVf2oXNvjbz9w95jOZheRX0joWyBabUmcVX
265FFpdcTw++LKyFzF2+MumVdEou5RLGaPkJAEqSPVEbl0Tl3lK6fOCHiflkCUnW
QdpFxCumaWODe8Gc9rkqpp7rgRLmBnizkZmzJLUMC5eFgHnrXgd390EAVwSVTqfF
OgVChVMlX+CIJsVd2uZrXBGbD70aUCLAXfS9wpWWr3GR/5Sn8vXQhqWmyxPlnVk0
8jfKmFyz4QS1Oh+rri8cutzlJvZGIAPkpicJaXzX/ScQQn0Atk/rQMk8EbCI7yWc
ftPvciYkrBuLtPmaD3eOknaGLUAcw5ueTUblmnf/x7CB72//nIMgpBPH4ayBib5V
9RY2K/g4ZOxz+2bPO4ktvbiWPoG0QFXzziw9cG4ZM6aHpF5/j2km/0JyDikbh5Xs
iU1N4LFIqeSYz4/vx36IEOkNXxbLyM+3SQYYjQFgJf++LT6AtS6K3dQtzKbrw4qK
XnAqkrq3AtvLaNEe73uq6qB8o92O1TAeLBfmJOAlylFAUwUAqzuho7C+1MhmMQiE
FW8O+LQNd/Z7j7AmhIgPM6Pbcg9+6WIwKHl+6epTEj+q1mdnOBDEutWTukDgPA35
fRi9rYjNO63wRkzIiOQ+BOIn+lqM+/9BRd/IXI1GeF9o3ad7UKeyGu4rVPR+mVur
p10gf24JdIlPucVHgkGZit4xmEgCmtafAwejBoctzp/K/HbTQ5ZAJQ2BbHpKrn0T
yLzXxNa89/3JEY9L1PWS6FWe/pFTXu2Zh1xDxANEN0WMQtmEDVp4EXKs8aQ00JU8
1fFSzVgNKk66+aN7dgXGNa0E5c2a9v2d63zU7ksCUTkA6lussP0eRy0Z1orW1xjz
d7b1tWPqVAu19Rl16nIGi5kNMOt6Bg+jZilmEDTXXu7QpahNSfSOgSbGXOTAN3Xm
6QUz845/ztM9UbapNkwKOZsYu/aTZRh1MzCq4T8hgrEjDINa+UvUZ7oMwoDpcAdK
PpcOPG+UHI6jiBbnE/HCCfhTt33/33Ie54b5GTwYLIw37K2x3cvVV0/01u9H5vw2
Ggg+QGujevlIDMbZl6hryI+oPjBAIW2DEo2ZvUWFFPUiANVUzUXp3U4UsjU9Sp5J
og877W9sMSKS3FDSkZrdd6Y23x1dSdiV0VGdSTMz43DaoDiM0yCZ5VGMeOj7BQdj
wMYki+w4uEsYiwsHPH/CN82C2oul8G+LLQSwvkgFnNNGb4L1Q0NeQul0Bc2XKHHe
ogDa0XUmeNYtInjqMsEKmuOa/J30vwqRVUBDDMYa3UmTUftcqtOfOevFGxrDDJK2
ZOjJ9O36VPwggOHxI2Lg1vQhXiitcdnMn5QMDF/CU3weH9MqRI6j2jN0Osmrds/u
mT7+fkwdZjq/KvN4ycbZZmiaMlYWk87p4yqs2xyHOtb+IxhDXXMz0K4WwCvJjVxf
0WD6Rzs94nJpUFPhe2Sai34iPUxidMyt+1AhJ1F4B4s0qlUpu/GhqYgwm/IRKVxK
vppBhqTZXrxOu8YpDtPvs2UBePxR0df+7ihbPSXOK7gyZopTcdt2+5H+aO9O7oBM
R9nXqLa9JQsd0X4Je17OdoAY8MI5oMeBAaUTeJd4HTnMoOw6GBMAXyXLVoaVLpH0
L2cZ1UCY6/jtxr72P0YbM/jAJ5ydJak2dZ1L36Wz69SIWfCe8TLRQ2CRs00N7nkJ
Xp9YuBVwaSP5ATCmDKc+pu3dTu6cG9Ekvafj/YVr6r3J0z0WuJVle3xp5bu1t+sT
39vT/DhicbkoIh14FLRN17+yOx69yYdt4oYhaWwgJzy1CyKudxqxz/+DwijyguoK
ojmAo2+TDJhkLL62pBh6IZeHn1fv4rm4hDEAZBoeFqTN4cGOOLxgKBRAN64Q6W1+
rxoqMV/5gPqcA/munBJkg3ygVnHwS/DYFc/bIBSCd9g+RgfnFItQk5eRInJMg1rO
AZuaWZX/o1tw+sq/TZ7Vpz8oaLLMBXJMz9uWqLQDrjK6/4oIwMgEtkefzLWTO/2A
dATs7bv1LYXA7TCZOE13jWIhQM4m8eHduo5P7eoq6t5OyAExa6R9uU2B1sgZ5nRB
V2sb1FnpmEm3jq6mXlf/CCkV19XruAHRH01bS4VDf4+V3evD9F2Yrji9PhY/LWO+
lXCn7rtYNIna8r2d7wmOmHuOMDlLuJAZshzZRpQnZUZEoBkveB0Nmg410yxKRanu
G6R1i87Lq9b19vLJlz+VRgbIwjrMoRyJt/FiTwNiardk5ht63vIXz/mzOYIN0Uyx
LtSDlXUzhUU/ZyLoF0NnMY3X+oqnP6vnlCzE5vQjLb7GE7i+m6NgGnPhHODsUCYV
fBqEQmAed5OtA3f2RUbzqaLg5zuqQ6fmhOYmlm5zN67J9vLu51kvrnIFKaoN975P
+Yj3e7TR+rBopqtwy6wUQ70LVyeBbzD5REP5/8mCTGnDys4PedR3ta+yKRKPcKD7
NmWbaKa7fYyJTZq0oAXLW1mTQNe/3Eg9znFE2kdEyLXjMRCh5Iu6+snJjnVaG72i
UIlp9jkoHfuxLG0LeX2qne2wbMqOJRSmpS0cCenJPNUM2EVOdSeEzox51XgosmR8
EBf7I5cQVWZp0hx/+B3jZJ0xC5RdCFr2CtgwSg5J0a9PEbkzNrki0Q1bbOFn1v7H
KRPMoTe1IbF1g9fpYc0EVPaBF1COrbouCTTRianmcijnNhtQrzgGHpOOxiKET/e9
+wuQve2hsWzb8a0G2zKu5H0K0dDW0kcZne6V2zEQvjrL9nd8v2uwWIfYzCfss2II
OQ1m+pfh8zVXQEldPGVWxn3LQmq0XIzoy0CVcpdgkc+StsG8AkJRb4Yp8r3uKjfb
4zxnDaNTUWzlDIxhVWaNSRUymPIbtI2FtgyypwN5mvyFowDPbwrKCBocSJkBTsNJ
ljPMovfUu9Uk15G4ByNRHq0e20DSAHks7z53f+nwrgPHyBIsfhf6zdzw4TSPjJy8
9bKPp2lK+ltA89FnpnnQbVOJM91LsqtGZVqz5fGhiPowQyzc4jlb79DiYQDLmsFQ
FGZ6xmvEkOHlcYzjDk+38z5FNM5hLW2xeOhoc59ZBSbCFpjgstCqwgqJrjDerP1Y
zFxi1C5Z7zdIjMAsMRmxe37YxaZcIf6CsArQyEQrBtoHfqHg2HLIjVJyJGBu1Mhe
zrh0nzyy2pb4XokxWRD2BUPNsvdAg21NSHwd5pXAD244MEQHbBe8Z81Vl/jRP6T6
I1XYPHYK8pJX860PVqWm6Uz0uOvnRwBzm/1c5rb/t1Mo9uWGHZCSTc6Ugakuax+1
h5qzZZICjLNs8tPMwe6ia1X3Azas3EnNpZGBjxQ30sjwk5gqNSjLcP9YL0jx6y0k
i1gZ4WPnh7Bibf1x77Oqbe4wFi3P+jBUpU2obm4omKmZ8lQf98RUtdGDAJJKtaZO
EdPF0eqTCZaqTvgJs1ZpM9K2/vU9yC6uLYnCDTTeV6SQykDN4VbrpJfHU84g0x7e
gBYw9msP4v/8fezGCVuyrVMe86ae8ZbRXu5dH4HVpHU6PfxhYjBqeQsZ81RX0h3g
r857Pb5m1vdhZfb9vVXoccf4kpW5P9SiEvUwGCmXehi1yQNH6VQsHvlRYE/eeltT
uRlqOzaDkuxrTofmOngm2RLHY8WgQjRPU4WM02wKlDx60Qtw/ysrtmSljE+kU4ze
Br1UobCjasylFcHNTtatfOmf/s/pFDVUak3pX/bK9vZi4NWhZLuZRuPKyuoAqbX7
HdHYMS0G8Pw6lx6LCaXWW7Y0bUTCSDXFL+Ux6H5OEcmGRv2VOTlhKjCH2d4Vo1Ks
bRrjaGqc2gUWhwuyKMVIpY/fPsrsoTYLGMUJumjMrP1umTNajSBXeEk0/w2DJGES
3UCLE+LItbA0RXmhIn4JiesY/V9vtmxZl6dEg3p/FWQRqCfXn7AFQml6aVNMRKvT
IH1/gTFkpER1fM9qBinb3Q7Rok74NBy1CLLx4JZYKc6LA0NJpbpmUTBj7DargtHE
FZjFa0Khq3boWJSMPBJYfwvfl+a2reoeGbPPLiI4oD8hPbzd+AKITn/snz1H3UUl
+1JMdSNLHQj0cV2NoYq0N8D8bifYRyrqKYu4bIC13fkVX2GIxVbFu6djy2xb6MxL
wybM5RkPAiY5X8FkNBUZ5lto4RPTLfKZK9lJ3wkRo7CEm+accYQNBchxl9b+idEO
YhdA4U/vxx2rqaFBD+FPN9JQXN5MnFNvNCr62sh7qlyV73PpvG+Pj1UGzxgk6TQf
iDIJNdZTfAZ0AwaxKiaUs4aehmLMfh8/FG6+kKCG+fzFZ+/O3TbxBtAaixUb6r0L
/WQXFOdG/OQElHYdzwqVtEdgXyfNlOgIxkQX53OZIxDzJMQA212nqltfz1YYhUYV
xyz02lanI8S+Gb66xkgA1SA3RDcyj131ja+ls+gCcbkcLKDUoExtD0SnOGVfBn8C
sC8+X+voVPTYvLbghiM7/abEq+SF8Jn9zLspNSRy1GYohknND6y3MoxVHlVmFp6G
w3+rIcDDs+4peaodWOfeY0OePj9UzYO29YFC3Z0cJjcRJrxuJ7fSiVL5ZRpXF/LH
7iVBuQT3sisZhdJUbt2itx6elZ29d6fJOXet/jUZOtuRUORiGAxW2nV5pK8iJxqx
mVmXI4SlcuPT44baqr+Dk1/VMPYrcLXcDZA0SHdzJWndjUDivsnytxy/9NEuUX5i
0QmstHXRKns2ypFiqRcdM3uJ+17Lcv38te6F6XmkjNzFP0dNDyh4u6wdHIoaOr5r
yiLSXhxxIeZ/0D5H9tdU4TIV7P5aIDFyEYIgUAAKcqO7FB0hTpZfIeR9TaCMmVLT
qlTs8lwKaiPWWkRaavsqv5Ini5M91LV6zidk2p8RuHJFin8P1ul+XAa/0rlOv4cP
EbY+7XK2//of8oWKTGTkOpJSSNZDOTPWi15McM/BOd9oa0q3Ncpvm0o7b62GD6Ve
GM9IrtuvWYY9Qlq8p2E/M8u0Iswcr7WjMIOvya6Xo8TIvXH6F6qGYKKZyVQOcUQn
Ba5eVLDXc/auQL9s7GbUjlxMc2DRptdZTQ1TusHOqCfabe5UcIiqNH2w96UzBNWg
zk6P6sJ32i4p4pX921M2dCPvrN1t+7rQ+Hp3aqWiuC6/bLmXxhEwvy2pMosMxdm0
qvvW+N6hK4+JcPxIgYp7H/LuZpxQB58p2Soz856vTWgP2DH8LBFrbzqhmtNKsQtS
9/Hh+FDaTWDZO4Y1ygNvOMsTLy8Egabqd3+N6SVaMZj4JKsfZnUl8Filai8ApHVQ
2fqoI/f4YtaMjGpGIz0NtN6+Kt4HofswuC5CzMZ7R9DchjAT6Z7r+7psTeZwgcvk
dfeidX8QCOY3iA90YrHu4NcdgpPm5hcaYJdGZaT3e1OUAnDAC4QdwQ+RDlEf9zIS
OUkcPRTORyY4ZSJxOV2VYnXJkYvYQEQh6eBbQLRj7GO63oJuUeAs7s6l2brD1le1
5eHsESVgoY8w/e5NRDe3afYdTvsrF8YLazdL9ZKvOCz7OBtwx74gy9JDAqMDoBIV
wE0p6nmPeSue6Yv5Ojc0r6kLL7Dn3MRqm2JPeahWMGqVo0Rm1WayVbPx+h7GKskf
Ud8v+77aNxHLK5h58spQsutkERiFbVkU7LmSpzbyzdYZ2Di7bKQPAUpHA6joX+z+
1GalwcM7zdcKMKTqpRQxwT8GlEWi8Lt4lxEQNPF8MsQILy7FAU0H02giXyBT26sM
1LNSLbLU/XnWOANzDM6d0iS5wRWKC5s5/gcjcc0YDyXrEW6F4aNerZyQLa6mAwKJ
ybj2EWwOLz//DjTrahJlgWrWh+Mr40cA6kdlrTBzLg626iOATEjQrpvac952GVcI
IWDzs6qUYmFo7XliYKLORHlnqPjMKnKLqNj62tGAXLGgNChDQrX7fwNx5d4C6AtA
uim5pRyQU0+j1e3v7pSxnqSDugMMxMfXohEXnEkqtK4wML5wzhI6rI4ncW86Uadm
OOCtj2nhkDFQ1xB8SQWJ6+ARViOqdCizcsf0OSY9wWZsYwGMe/6rwclDhwxPYdhW
kqtAGxo/dtKOGunUk2SkLUWGI4jeL2sG/tbk1Rqpd+4nHufiVm8L8c4jWr5E44xc
PZJobx7ZQ1UQWbpduSKbSayKrrutlncDnKvrgUMUtOFMGVG13dLYhStc8tZkJj6x
3faXfKO8KT5IJVojweTYrwsrRW52luBgnnpTQHztyDIVYH1MhNDXG5MOBQ/Y63Rp
qlt3fVORV1KhWDdYRq42agmNyGyZxw2v5cjCxuteWWWjVd934ASbzLKVpvglOMpl
L7OQjS3UM9O5fNDgm7mTiVYmEkz8EZKkkc5ytGlIltmredcmZXsx+QMVRIhzs0Zt
Wz+nKJ3aitBCaNvfSqNPyVeHvX3a1GxNwDfWqungqObKTsoiCy+bUtH9uKD7sS4m
gk55Gfrlm7DHvrwJXM+Dkc0Ttwpd+5w5g7iQb4ekwVy6uQ687M8fUo+lrrqNoBix
Ulk7Gh5g4i6eqDAU7YCFTU/EFbcdPKEzR9NkOxezv16qPjfab1luLxbepqiEreje
gjLmz+MdeYj71e7r7sq+pAqps8mtDX0NhY7vQahI7zDlEAreX8aDOP1UtboI3ZJ4
T9j7btVInv4PxZ04I8qfOs/H6Bqg8NvIuSLZe3wvod4MuuXbVsHua4U7I+hVddXN
c1k6CRLe+JEhnKugsVUI3WHCIjSOcDy353kTOV7jOICq1qQ3anwclHHLZuRltkgy
rnJ5fjNSZ9GTztlKiNsJVmBrK7kFx4SaQcWitVAcnBE2iUg4mSSeqC0EAhgXh1JF
vjtswohGq/a102lRsyprHji5yZ+flWH7YCjotAI/8hxHfYKPczMJfihbwXsiq5jx
NtTQVRNoNVtE52VtAleMquTyb55tf++n4YLnxO1vGhwzrQ/w3rI7MjlsWNOassPZ
mc3vjefZ13LpUMHaSHopf+LX6k1ph1jLwWZlSSJFo3mFa3mTypZa0bk4+aS2djRn
YwB3ERDSf6REnTAzi7bJSk3MIUfqD123uWMXQqXhZWl8aqhhTgD8yiaDIe81xsDy
RLLG6x15svdxy4yzn3HF6LuTQdyNfdfl5q3GkJwMfaedK7OAPDHITIMLxDBNerfi
AAzFQ//JbFi1av18Mm3mSKX5ABIrh0W0BgUNtr57Wkrt/JTPEj3EQvndiEQwl4iq
YOxJ3dqDu/vXpVNU2TlM19fWSc0mNO26KWHMGKup6DCYDxzSVXnvGDG4CXrxkoud
6mx/IBxLVWodMTzBLWgLdtAi4S2GOzkeSDd0EEK3dKm9ejnW5fuHqe5R7UsP3ckU
GNkw/Rh1nZNXA/H9P8hicjPa8jlDQ45G8tzxMKLsojamGaHvw1ymp30tffwGajKd
Bh05G9qxBfHcDceoqePspP+T6uPUCvlmzf40l5KHHrdAb/z62h8AAYDRSRUyUZ1e
CHfBFM1GB4cpZy4NwcAWc+CqlYCSGFLw7l06EeFpOrHahphlBufMfIDMToIuCYi7
2Dd77nXP4C2SQu8mPBHEn+V/24h39P82nPRitABAsmVzC+vDCrM5AJEqPZX8CPrP
Qcm99vBwFSuZTyhjpiVdac67Np65Wz9N8vuVUTOyvdfRt0F9Y4jtbbrxr2YDhfnK
lurrDVWNmpIVx5lDeBkAkqm5JZHKC0RasN9zZt4L0w3L7hbdo7D3IqocxaeTu5bq
prO2LkQDcuwgyQzantP6imp/pi33dbJNaRns82Je7aD8k2EK6D8V7G0WyFtusxsW
9VUIpcrPbo+Jm5HKcnFRp+Tj+0ywaAWZHztrAwiwuBVihD3zI53J0f/YeEed25yv
yWFRAFnhQ7maohGuubq5modn7NRjXL6GRw+YDg1DKYHH1ZbVZBFZ1zZnDLgvyVoL
yAsAm4uaeYDVIvWVhk7Zt4Rt4H0r8vpknBV/OTIVJVvjOHDfm3cMIAy0zbSq9QG8
+jgmhyJ4aADqYjnO84vJ+DLSv9F8foHgUuTEt/i+11F803VP2T9BlPs5uD4+oFlQ
Kb1oYXsJSPE2JxQ6Wj6nQ4pyDHsL9m/TJvcdqLkasa3hFMXUG2A4MB9q8ChjkCC5
LIwLErTysqYXYpLdSHlI8q+aU9Nzunwsf5b8QF+iiEoZTJtNQsyL9cxBgWWfE6Al
kuKaLWfOouPUaSKmA99KAOqQ1kng8cisiR2ccJ2Afu19mj/UmmTAxXxs++ebxlz8
LOPhmiQTCzpOmbqEUBkIhQBIZmvRkr0sjPv/LB1WdGjVh6nPn4wdZliED0keFmBo
4HWR+Fnxe/xZ/dTk23o7iQprnPOkEOrD7t/5c+ikjyz+Hj02qRTXUyFQcx8sFHhz
y5W8/vjymZYOzgbiy4unSOYl5QPpQuHkPxJ6dEEIW8D11V5m150chs3LJ/n8bpn2
7TkWR3ZPlzL7HKzCU0lbWdsPeX/rdAOHzONSobwDqGVcbW4zX/amtW26kY5IkgFD
eK6Xb20rNa5dVMu4Cm7B7WkrAtNXcLorOIoPdwtaKeRogWNNWEtuprFhW66Hr0JZ
rcVFb1raROWQ1AP07PWl2CgImIEyLUxz5WGM/+68esk3/rgDZtjmZ7Lm9lo+K/XQ
jDYm3TsJ9ItnhjKPJYWQWZ89VvfUqdnEYlISLZBl3Oyyg6cgHGvJjkmT1wZgdB9q
KCqpu5yAOBl5mV6WgcC6lsY+Yz4k9dBwWmL05Q9xD+2v6Ot5NxuRzuVqk+2KL0Dr
hVZl2gFggUiEEJVlvYUr0rq81fyMZ5/SEhWtRnQwHUel+e+7HjCJKST2GqezRkuT
lI/4GRQve5qw4hw4+2q9L7WzLv01UPjtoOioV/SY+OE5tgwKlZp4TQFjPhlxVlXv
0WPgPWTPGotMkE8rTVm+m61R/R67FzqqaeiTkphkyS2MLzk7ojrRC+UORIiYMDl5
6tBHDiKPajM332OUhnIB62lbtFZdgvVBFrsmlMSwvuI15YRrAr5KicW5JZ0yUmf6
yZQQCsg/02dFyAGgLB1dd6LcotOA9v4mbI6g1jRA/KKlSB0U5WwHS+ODOM0vg95b
NoEEM/HhOPgsGS9SRxVj3sD1sG1yXwyrjphv+kneW/7cr6YBL/PsaV4xYBflxp7U
4Fx3Jj8gRCK7jSkN5VfVZ6dqEdaT8CMOFwCEcUyNORk1lZh8ImbIchEm3tq2wbEA
Auvh+83PbzpdMulUQGPmfgqDK4OizY3+eE61EV7zv1lggMVelFObPvpulnmQ8/p0
8Cmx7+aQDo795cSWZIQARhjISOhyXEkklNuVizZttqBVVg3YeSZungWF1k11IM0f
28iRtMOSADe1sCPaEyvazDu9q4+T7w4TUROGZIQkdAc66HxUaMZJ+CHvnU9QuqEQ
C24T7h32yPc7QG7DBaIGwx/5Nvot0zPjkQB1DN7S0uj6uyGKSu9E10XRUM5EoEN6
KmD8opYkNhVLa8mrjQzZtJPbipIHQjwcyP+11CI1JvjBVlwam492Aqt8dkCYxELC
6uiU2/eP7BO5TYuvAZyDu/kIVaRt/O6ejrybTjPkwwQfLuCCTu9LStNUy5ng4q6X
pbfyIXq7EoKIxvk9J5+GLEzMYHJCApnkw2FawM88fxkIXyRGI8Ch/4iL3DSVxJfV
6n8mFDs0li3OHxcUqp1ljoCoa3bOcKvaCgPw5MrxbYEL+m1hWRdf8tVXsOcwuGnJ
XDJoFaUB6xB5UaZqGX9r1jS6oFJhDAHBngucgW5x1Y6ISefQ+sFHDNiT2u59vtai
hLKIeTys/C20mFZlee55ndaIHwy8ltQvt1JpDAaGfYJjUfCg/18c1IfnqmVPCKx2
SuO9FeTSmAfYHK+RsE+GiRjjgfwccjzEfVo1OT7bR/SlfVqcT+qQxXxyA8xOoJAC
wh/lE9ubvr4UjXsFTn62kqj0ed8PaB5kV6XQ4XJk1L5rrOuaEtUnw3bPlVB+WZx5
3hqrXKq/c9Tb2BN0WiS+YvYJX4DqNwNM7KNPLdm1y9Snoly+O5xfKhCSvNrONcL4
yMewzpMJbbFxWatYwV0JZvN/TQXw7tPce2lZpZGJA7KtIhKjG2au5REk3QibCGpd
uE+MNjW3DtUX1a9MfqC5NDl3l5zufV4MArJrv5DSa6NRkjtZeOErBa5QKeKNNY1J
4pGDLPPy3kvqXWDdMtGlATZGZb5HpqszFlH+hhMhQ3gkA/8zSynvPIJGyfxOi9k7
FSCSiW1YUNqRBtGNqLtdvBaVKWDhr32drD8aHq4m5BuODwPtYonv6o0uoEk1T2sl
Do+KgtQymXm3HoVyaazCt1SMGRkTL11CwAbN4FSQmLxKsnNuoAeIcj5JgEQMbOEF
cgUSuo9/OXutuHkop2KBxxQBe6Cz4nrvVFChtTrcV7K5ACHwdOXp2DFYKv0u4ZVW
X8OqIBL9ise+W1KxkiIeMa41X0BrthQYzKzR0gtyjQ0zx3GyjajjvZQRdwW7/vV/
O3CKvH4LtIJA719gBrTQYQUtDEc0NF9APpvimyvDvW/dWFbZXH7exMJrPhNjTiWz
I3/nqnAFaw+K/g7CwnPqte7VPCAY0Ht4tSVO8fjeTUK9xEGQ7wk6HiOkOKqza9UL
y/z57whLTPs28huFQhhJOS1WXSJeMx6StB4axNJfzpEwQAi8opjzV0Do/FofcjKr
T6ZUnDHdNnKNqJtoUFbeVHtL1HNQnWPwJ9PHh7ZYz4tUs/pnhgyLklzvgRg9j5Gq
aiXL8hPH3K31dnreZICuJZyb4Lye63NBEAPGZAK9H/5+3wfbDpSutMgybabaPgnN
Ory45Apeq+LqQVUCQyTAz2rVvrpFCqpMxthouBVAH8Fli1YVPkgSWHPeucYr777K
tGdTJVSCu0O9imWhpiLLhrL9ZjEHCYUdC03M/RdVNqau2t88ZXcWCu7ZHXrZaKwZ
G3ljvI90dImU1slnY8r4d3LMzykVTTmW/mUtXH9bgvPG+PdMdjaTaiKrqHfELrs6
Xv1+6FHXf0TucGV5ddlnya2ptQBHMQAtgwE2aOaKHvjQPUl1jBN35ZZCJVqNckxS
Pv0QvDWR0WUfREd/+YFBbCwi47fafirxmdvpAg3OGbSFZcudOJvuWb75e5dtJaa4
0bDZOrflHISryTIHW0yG3A91quuEwBYdU+RSgcME+Mv4f2T92sTauPHhibPeVcNn
j+In1i3YlhE1jJWLlGFWZKHSqdASl58KeemyhOhJkutGoc/cb0Q1cfpi45RlYt46
QZtOzhwnJKMzY/mVOt62pcRQvC5szXaV7T65xypPdmSgJA2euoIRmFebl7nz39j+
DZ1frHNrE4IMesKsyzHRub7lQT7nGV0XdQuoAT3wIhSVa6fUQzhShYlKvJV+SM9S
+6NjrJXlCg/Lz5T5Ym9STeJlLhkyiEzUlS/PIWlLUCG63wwrSXH5zunMEkPvocIz
hFLJ6jeciFKglUMc2I5LpMLlCfKZ/yoo1tZvjZqnl+fAIaljjnCDqm7ZD6tU2dsv
z2J1kxhYk4zuoSDEWWFXddIfEg8T1qGnsrC1zJuqaMeCLe2La8I4rjCzUqU2qY+b
5S8EHqjTpnO5WA87AkXDq90gMow3K2sYNOT3+5qa/hYaMxI2j02PbcT0N7Z/FnaI
7Ll1dqD3dYfn2I8OlXHrP7A3evOXGomIiBjM8Cl9rGXmA6peydgrgc53nWHdZudA
rB+uIVtytpzH1aslQfXJxHTqINVBAncttAuE/QneVgvMwrXHgxff2VkIxzMHoCBY
hS8ngotTLoyCBobd9RlsWs4n9hHE+ICYBlvvHfSRfOGOo7SlEPWncVTTGmCwUqeF
up+R2ou0epTETql6ggjRfytHsirml8bFELoEzw81Fk7+somr9/1sDvWgenwkdfAL
lF/Kb6qHPjFWDZb2jL/3O2YaOaWq7M16F45Bam+G85HUzyUUjDc4bhftFwW76E2+
Y5MvJhc70c2mSzSOFuno7Vrje8Pv91DhRpAsK7aDjzqWfcir+TiqkDpm7JQaNVXC
JERYKiwWlRjBZm+fBj70wBW9yOLQONMQH/qGjbkWwAZOuWHi66afNmKvyGfz+/vE
XEjtUszdKwOhsjiFN3ZUxsttfDRcs6u91EYOmRaABnKXQmAcVu60NCwAJeq4L8bv
T5mU3U1K3gMNCbdoZGLS8GmwVQIkfOBG7Jb3JNeDntbJmyFN/Zk/WllKZEE2bUzB
ROZpthUx0/+YOKct2KhNSMZsCsSgKfe5PnOEtM//oxjuuqKmYbyN9hVkXbihhxTn
DvkeS2M130beklZi7YuQVtFV6Tp9aH8I3KUcA+AUtQSDOTf/ANW36jRpv+kePsi1
BuN4Vmp1/mNI77ilR2LLBDkVEkULeo0LEMvcPcK0VuanfNSyKGaayg/ywbOgfMlV
AxAuBNYnNsmEakPo1s95562UjuSeS7W4wpN4aZhg/bIMbPcw+ucDuFZcbSq/FTGf
pZIcIDFrpoRc0dWO04cZr01hjCjH6pPutXOqFWPyPYO4VUOUFjCJqB6Gk3h4EhLd
7ruNgKjDkRSHmI7sWDzAy8jn1zg2nZPpOodPNCpNp7So4OrzNg0I9bxVJRSnABL+
/O6Hd1n5joPe6lRd0Kic4BJAUHx7KqsopLnrrw9rGkekpoTrsXd94MBr8ZxjONpl
sKJC3dWx0wC2E+ZOoNBoPH87BlySftaN0xPNhx2X8MvxSTUFnHblvoq0GYH4mi3C
eLKeaiVgaz/dJksTVgT5ah7GJFV5gpJWaFXSnO+kYkFeRrSYtIwbJFR2Av9xdW0d
3KgnQTbfsJqAB019BMCF5pvaXlT46vBfpRpMAUTTvRKCjJ1e4/ubVsUr5+8HQa9V
LcO+OhmiB/6puOze8HQgqP9wni10bIXxUQncNQWrlInqbvkvYFjZHLH5RJ2eAbQL
lZF44EnOTIPy0BLm39nTD1ECjb4aHTQwPbmjZarQNYBkEvAIohLzJBhjeoyClB9U
DNeknMIF2iqo9m/ZO1aGdYWgIQ2LAimMd3OgBSZ7QnqiqJuggsbPz7MMYCLVvrFg
6jsVcvxy6ECf5Zdxmpt8cPDKHq1l40Q/IxHmJC9z//SupEggqzEDx6CIfqrDEW7d
dpQJ5ujTci8M9KIxrktFbIO3dZjsxHcCuTxQ3QCUsbsGg4EfTeosKMPQ7Lq9nsf7
BR3X2BrVt4ZaD93orKc20rsoOMXxCvUPtL0/HSKKvzaoPBNwWxk1OkrHD+sHlCCU
QnuQNkvNOhBZQ34zQX5UoKNGet0seglj7E4HzOn8AuMzZselAZAd3Y3Ggz4YaNnm
6FxMQkDMvyDTOdWTGbdGcBlm4YMMK630fyylncWtzpF1dDwahmomUgK07wJaJrpr
EkrQ+vuV7yDgaLMIxeabFPC3zGFPlrdxTLg0CvDVuPytS9Aox5c7wF31aTGtPTm5
H1170VzpT2vQcGU92LydgOeU2VhtYCOfmeVazCHEzZHEb0WLNCV1vE2Idf/5n9OT
fQaLOmUo5iS9akJjNljC0kunI5HOs3o04NfAbcYDkr6mm97yKM69sj2mrXZX2q0/
yMd0113k0f31fHcPLdkhaPSTF/9JED/8wIV05zmpFtlvTu3Fd9LW4JUfRONm0Yti
o1ayNkO44HOGZ2oDZmuDuC3lBALt41hZfMmdMPSAArKuGj18g3ZFDlVoGpPzIZlj
QhNrVUsLfOPjGzxeMlannVWnJkCIlkP7XDGgcn+6kdppjtn4THjpzxr67JRY36op
VyDJgbkh/3VK3rAJ+9MGjMFKPQLEPJL+lQ2QujyV/7XYMnXJbmkv+PqKP7C+rbbe
HCTbcOhApZDr6r/a330HS3luwxqVBAaGsqiVECMYg8L0Y/zrwxUJNzRP+M78WsUE
kR1vx6QSWmzQlFdpEHjYfdIjcVzyBvibfvpzU6r37AUK+hgYPQMNAWRoUm2tV9gX
hDCfzUzE0TXJnvTPXnmBLCjKc+FXpY+NSEUShFDA741NgAU3PgSi1dLonzxz/Itn
baTPHU/CKz/h//bf/KMYq3YiQPUXb0KTafJ7l0XoeDdfqYr1ox46k5LOX559QfkF
ydMaI7Oc4fEYREA2NKNNaGymBPIDgXQWJl1hQS/AbnIbyvY82r2C0sLQukDoPUXX
3IYD7QH03zEJ85osSeTSGl7XzDO17QE2rUpULNq3HnQryMrg2qubqVAlALJIgg0c
2BHAFje0XNiOkd1nfJsqyQpM5jd7FM6vz2vRYr7SpfQNjAaGipgzrNXayv/w5n9T
tlswD8RWhBs7ePscrHD1k2Y5Wu7yRFXXqI+wnx+3A/jI4UetQjj84dVvKqcDty0Q
Q6N+ujjJkuJNIBjvFDAA3lNOqubaWDq/qr3Y/gCatZpz1OtOx4jSeoU9y4LZG8Q0
nl5FybOc0yHMrNVWnVYThbk0FQg3FJTmvtbwAYyk8aoDANo2OJfZSBNnTb4bdopm
UquWm/LRxe73g+6ZvlDylbrTa9OlE1SKSZ0KP/Fjgi2jLM+Q/zpkbjKGbLlRez0w
HuoSorOuL/K0DJdKEN/rdMYKHkluvqTMedXtsh2NAULnNYUk3PjJ28kg0ka0a45C
ZrHZCYfsZ7ZPRb+4DYIgW6IhliQX6NDquZ7luR2vwi2ODr9DH8Vv0VBa5oxF0KvJ
cpgL1GQtCl7A6bwv7RRKSLPzzbSlB4YOzT6DHJ6WGj5apkuzhlnD/OgToKOq7OXD
ipJXabTs+s+2JA+L5s6X1z2xKP9Y73JJxo4yoSB+A1zIop0lCJpPTC5VepmrSKv2
qepx1teUuWFLylojhWyIgOFWukEy3CUC/w1V2raVPY70xkSQDc2lj4ypaA2oFSyn
ri6RSXtjERMFh6mgsN6uBVxWy1ygS5+fV7pVQ9u2vXbeASwxsq3lX2lHVxxn07U9
J9aH5Iyjlr9yNzWgxmezzpOKkjFZ43KJNGojCTevIrs/Kf83/AuwS6oOTEipol+U
VkdS+ArnOp55O7vWtmYMCLoMXl7BtTW+5kWl4YYQUpVMSiquTgERg+VGkr0zObxU
aisek9sNMq3HyNuZcQgwNa+vnr9VdsbU8js8YfSU03tXs+zLsBvIgzo01eZLiLmf
IY0ILBdmyP/UlT234MBMy0Xohle+cpcINQfKas2/nUuhncfHBssSoq3DsVM4RBTC
MkjjCabKWC4Oy/SYxjac6l3qDYaj/1dzTCOsh0D0y73qEtY//8gDzLoxM9HuiDXI
vO1btqRXzC2/CmRMuZ87ifoh16BSfTkuBfIAQe/Kji+xUBnsFTc38cuXVYidsye4
J+HKFSQIdg0B+JPNvwWsvRB9R7WTDVf0CtK3IsXFGOkiN9gaZj/YICLLpQflI4cc
qbW/XZ0qCNvIkA4XEHBwLhQ24A1NhMgB+LdIzWik2MRAVnlVAH8iewHe8PoW/D4v
aoElHmQ1AbpiedeO+5JyOKxML/Re0wArTNiXHOPV829p2+1FhN/XN7ad+4CUTPgV
53iccyVfZoQirjZTjpxOtZZl4+B/LXuX5quZIxUw0zfPN/H3piq6NJWaKzbvdtDa
wIks1xSmiDQN0BsdL/aBJOnVAQe5M7/xPtelsEGFSaR1zSZPz5IaP3fPgpB4KdDG
9wdiQeCUEgPuABGkkOGxu2w/RdqpcczqgbKLRjMZFjB15GunyUf6NtUaupK2eDNK
Ns/1VD1SeQI13JI5FALgzBcED7+p6LkppjfjaXehms4biSCkkjZdCMuA8h4DDw3W
rWVCGuL+JadPy27CF9Cam8w8MFMbms7xpxRes59n5m/XqPcEVw2FarO2VkB7rRNx
oHiWVtNyIsqBH40xzw1j0+VWEizMAVZqktspiPfh/w9nc1dtqsew22QfEs7LvEQI
YQgEXJAE7pzT7W9/fxfMItytCxJ6SUknCqV1Z/Og1MSC7O2QYbjRYChjgw6bPbYf
XhM2S8xlvd+KprD8Fg8ino5NJ1ihbL16G7reeA8zJDcMjgS9i7dPUkwf2XNBqR17
6jqa++wi4xL0OfXA2GF99FetnkNSKbDA9SJRdMpL0ZiISMRK9nS1O2FKawOjjRoH
6LQrAj3VDAeBr4S+u9Le0fZ1XW0OBpRtk/ExMdbJoppZbWcOO2sAgr7Axw3eFMZI
iLSvx0ISDI0fP1tuwRivW0DKsmFhkgb22mSmHGDfeGrWPnqM3ftOzBvHqzgS/ste
Wt7lLgHq+pJQFhNK46OHZLoZPtb+CPMqn18dNaH+2nHC84uZIjV6GpbzS2WeMkCt
EKFrFaISM47ihKIX0vRU8pN3TuQYpsy7hCFNbFlRx9a2JCv2Kfo9NfU2tnJfd54W
kr5+qOA7RkMw/qFaM6Wf/yQRwgadFvMgq36ZJe9riJI84KLZ0JRTCP50o3kPtrLy
YR0vt1i5g6StYVwcHaiv940xSqi5+QM6KAjdIn8675Rkp8kdCD5e00si55AeRMM/
rKZxCS0r9Ed5hiPgpox86mnyLvmSx+nk5Ba/RYoD9UnLaF3N0vPyANcwZg7M2ob6
+x3iZZGmglzU29VlQKDIVLhFJGjuF2soL4mHP3kdBst/nwVUDXoLBB/uXvMP4QvS
dXi685M47T7y1Muv+Ba07aoqz+3QaDD/Nh4lX00ebK1c2r3g/90vRqRnRJfx5H34
nUNz6dlT5c3v+/oJz21xMxzrZ+MgjyQTawk5VBdHUZ2Y0UZyfruS7h4HhqzrgbAj
J+If8NRwdcUVYFuD6efxxix/REJ1I5tB6ypGuimS/oSiqZhqPS7cfDzgwiWDoHMe
zCqyCNlEaH27RBsz/3MygdYNsvrdK6LXQEUrxHw0fGrpVY4WkpmN/F7AWjISHlH3
k9hw0gSsNrlIsvaOEtMjr9krc1WAWoddvMi/OdvcwvnooMFkxC5TOvciPOEPVa9b
MgVX/q3NUW2Npy91Tl9D8GWmHY7ST1QMKFTyxXH+h/VIE3Hs4i6XJ5k/sh29yE/T
LuTy+fqD62SrH7Z4jhdNzClm4kV6S0Y29PBUjjbwYmWqT50+RvukUFOsFk5zDJFU
GHmuhxIGBlWXcXiI3I/YSJEu0sJtJ9mm3YV8zPOGp5UNz3jbsOEMJJ/TcTtXKPa+
LJihHVUBGjQioaS1giOpuA4/G6A7o12Z4+4vDDcIIYh0t2MCOnOwWftr7fcyizex
p45GNrZXV2mU/4C+DmN2qWjyV2IdyuY6aNEeBNd9E4hSAgLY7AX+LsVFva8c+jeE
A4N6LwiwwvkQD/TdjB0tNrsOgp+3uz7H3CPgWmahzxJi5OSgMQ2mi4yfLAbGDTqA
sXP6aG0+w9FClA/y9pbuMHQ5aATZlHkcY4AWhzI1oa02JGMJnmEQOssWjiseRMw5
+T7SrcuOnWuWe7CCQwufN+vcuUOJGMvGkfaeympABBlcfXh8mn7iF6eu45+cT+hr
Smu+eL0MwJ4bNiqXeHBO0KhJ3EIhJo1DUjqfFZpvXJRFwf0LDNs6G5jEc4PCj7Sn
1nuR43lFZwO6WXU6ODPjwKzbpVGwcQsn9T1ayTUShgwPZ7/SM3u32B8z+pFFvggV
i0BU3NQCYJyfT5wtTxfifdLT/AmaF5iUmb49/sCK4eTeUH9KXH4eTCPOh3hwS8f4
9Srl3wxlWlnooGtZ67ipTbjZ6ZxWuJhae8nSaCWHVKPeLOiJSgv5Fo29Zb592sIL
Kdskorl8Kkg9mAPzVxeR3RHMTiI/RNpV+6X+mDIVHc5ibhFUgVvTihIBOaRKSnLQ
01rLCAGiJnFuSkYtI87j14loYZ2zlIFqUkjWReGBTicflpDclgHs8lq/osVLoA0P
pIbOzBfeNYWKhveMw+oF9psdG7rLdUEAAuCjGRM12+sC1epbrpiGSL6IKbONCtAh
76gsDzLxWMazdMnEgzVzwJKltdwfBenOOt1fPaJ+cQXU8DRFQ2oOZKPYOpyJTwss
KaQ9gnaI/qQxWvd4oRXBYnifTj1QXXBpcvTUz5xMFGFt1VNfH3S1Wk/U4BgTcFR8
u0qKkcW7h55sijhrE5xcsSjmFrhIsg2Em2rtsvew6o8hj9IYYlIq7N0Tohs41goe
4tlI3cm0KiT8deofGqsGT9617r/3XUo4muDjl6rd5sm/w8nN3cCZoQe9S16usC0O
QMhsOoJrFEyczIITLeDyvaCLhnjKDu8Wx6iU9n8uSZoOOvVS+0N/zqF3p5OTGmom
yxkfLsjbB9A+KPCt3RvOjQnM5Ivsde7ShR6crZ8jt9uKpXOSXcN2FnihmGYVgzm+
YMoFUs2iM10Ij0qaZmDI54x+bo6w/gQIaykyoHtk450ULPWSlo6c+psJHlOBDS0e
HVwvu7bwMa991MyxiVXvBh6i0eQhS5OcpFNH9plOLU1CzFJUjdy9XDb1sDovIY/U
4R94Rjr/iP2Bht2C8sRafp2+RxBfqRKUTAHb/PmrlQVdhBwnqn2SFRpEgqEU9Bn/
ff7WxHIs322SM27xt7EjjpfB6hJYMUnTfg51BXUTe2NTho7Snw4+rUOoQaDqOVaI
EK5eMkTqQm0tQstecTiZqpXXiEyk/3HiDcDs0qfOZ9ohWR+MorkvP3YMQ81uo7uw
hcL1S6EuQcf5+9P0OvyhXbAWEF5Sm+I8vEQlp57lNzpDcEaegcuXazro1e7jBYJ0
B+lBsIKJd3QRNXImPJjF1LeJ4igKnDJJlcuDi9KyvYR3NnZrbhbfIkDYlP7WDfqD
jhmNAXG9zDVr/uG/m2i0XaqaOTPjwV4F74isRhD0U4UbHJOgj3owDLxLY49KV+sO
2y6Y6olsm27utkgiwalfzKkm1r5BnafrHbQTjqF+MMsDTUFyTLkEACPpKtGCcHMD
5rcmodLlBZVoC+KOEL+xM+RnjlAjwQBUHMHILOsBtqL/J+sxpumRPtcesss1ODXI
OKfrMq3XwQQgUVYSDTMbQEIkwZGK1tbg625q07dDz8Ezk8x+sQ+QXNeqZsdHFMHB
3YKKe5FFO0mEstVgKN9s90r1gsoHjQAlYgYX9773pWE7T1NsOq7+n7vIsttREXHG
1RLPKBbVM0wdjqZxEJPqEbBau+QTeTkLkjVl1AEpL6y8nRjuhGysFwgwiM5hKG06
RtWwXDF1UZ/u+QWhVqDaceSIeN5K0x8O3xjAwNGKoyLnugcj6fOis5AtYFoGbkXD
FLE8xrtkQ+EkU+18kJduFXnntDoJDFB5w8mYbgkXGR+qkkIMhqVEoR1PEQzS/2LQ
77WzL9FELcrWz5B+5cI7T7nHidgNc09A+hIbO0tzT/1bLiGjPjZ+YWvuFw6Jg6J7
uz7Yjyov8XcBLXJbV3MvROnJyMBmqmv6mdDWOs0w7LVcw+e5T2FpAMufL1PfNyNo
ADjvf1vnlHBBVy2JdQcjLoLKt+0ERUlbRIhj4iCQdDOBTijGkdu94156CAPcAjVb
yxiE03yFZD+tBY3F2+WYlnWGRRUJVy7ZhfOXaHhkXHlqGnnBMFQliwLyGm7+xZ6G
ffqOgzF+h9Ta4oLbfl3HjhjKnmJ9g+1h7NUBd7d37U8DYsZ/Prxy8e9tyhxWK9/V
MbhNpSYloq6IqGisXxdDLo0P9mDoAZqtW06rqoM+q3DpK8VqWI6L8J3DJT8wJ28N
bM4pHZTsymKEzs73v4qGcLBJQzVK9spL+CR6ZqqrpuZm1pY7XONMDmKeFNsYce1e
bVJCqSs+M6asmerH94lQE2BCP0eqH4QdRBzbSF+7k5DqW4lrckFWI3HVBnP01utJ
AFadtBvuDZ2/9OnCrXYgtY9Ilvqm1P9wDnOHx1DgaUr6UHEVGDSI9HTyeir9p4pu
gPamSf14R9Ax1Zi/8KeMszvJF1lvDZT2b4IG10x+nOgsb7fpPNBcwnCd2H0xlJDy
fW/EtCZbzaCOWNnVi3J+Cl8sztcuEwdB2hhFQiZqvcIFM+QhPzQ31LfXgtfW48UW
iMurecHJPl8Yf+fFVVJPlfXu5EkNMGoY7KuvW+tlYqB6eFOqYQmrvbrG07QKLTtw
vCnxINSy7+MzzMYrMGCpJ+yaj4mLYX5qv8BlHhvTK/hSJHozHMe58Y7dSV/GVkwq
LoDu6w1oK5tGMBXzLzydDXWGA+dHquvnSF6IIjz6gBztSwDdV/C1XnpQ3LXQsbDs
9uT3OIEypIcRqK9Gxd91QnkZOOmQP/sFLhjL7K7LGxa8UlQf/PNzLn3//ntmnd8W
7ftQu3m624hrhNunCGMrRQwn61dIP39JXxYL1SDPfjra7IpITo8V9FdINxTCdgKV
ITE4jGb5pOfWqFY7T1lsBj8IxLoA2gr0GbdpsJWqhttlJVof0zQyE1X/NIbrVu8f
+jxAKV3l3exNKWo6yIZmRfa8EVhnXj0dp58e3lZed/GSV+FJD2EDLr4X8xiiquvF
c7f8s6q3ArsiIB82iKzTtv9ZnAJ+eqNGV3abtmU8FbJf/iEppIX6kVs+aegJYWqN
gkKfazDPxwIK2wdgWti2FJzt1ECafHMAHBgz+UECPr3gk+q5OUZVgD+a4Ha3cKYr
pMaz3GQz7b2ZUPGb7NESDIZQmyJ/Cfua+1XTe5dFS7tg89b98zIDOR26ETkG58q1
21fSkPlCzfyb0PZDP27gWGgXBHURZbf8AV7IxbIRm7RBIW2bMWQ7pkkKG1fvpOEL
Cdu+BBPuHQ3YE03IZMFyVfjXdrv5wgRDhV8JxuVjEBgm6AhtpVxxuvrpqtAsPecD
KEOjtcCe5z29uyD+/367yDAu+g4soax6qut9GdozrUcL6OMdERBduFoMukO0Qgkd
6cxNT9Yk86CsKOqgggDAHCmOXO+Oh+8akIsQW9dBCzISzm60UayWqEeYc1vlMImX
UwpQttoNhDEMTPpQT55e28CnBxJ0r0KPekF5ULDlfxPbrv2twP9yCpSsJWqVb/Xx
eMiDDFh8yAOc87C5McV0ItjGDBYjpT3ROqkUt6gb27ObEms1G42vpgbjdFAN+lUp
BuqcZwqOrLRCfmnorTx4JNYt0tg8weubfJbdm0wWkcUNsS4bPIUxqptligqV4ihu
5+e33j3o+eEPX+wVd3inq6JYA7tIZHbL8hN8iuRULZsSGnS6/Uyl+rY9kd71C7pt
LmwvG/wNYMg8NTrDCrZcuUmDfz0Q1NjfdPUBTGVsgSxcJES45iKtkz+R+nkff2fz
yusmFk5nrAKOj9rZNQVMHlbKGRX0KT3nLXsyXc1g4PESA1dItKB12uvTPdg7OYeA
zmJPRbdV6EQujgqWvSqx0k/0OU7RfB2I8NcOKPUuT5q5BudWAYyEuse48vFFIZbI
XTGZkANCy9GuvGU0QVwK2RZFu39AFBbAKXmy8rO7XajcO/vKYBKwIuBMc1CDlGHt
ROwhUpvrhPT7/RckD3ZAElVcIqTgUaIPCJ407SHyX7z8a3k/ZorWWB7Z/20O4/Hu
2Cj/D1e1BssJkvl/Fj+jTeRLBhRi3FDX7dlCJgnbDOT68Aqqp9S/xBYnTiZJUeCL
CJ0wlaRrXzdT0yXaiNMu0b6Wiwn/aAWCQXKNl5+rzwL5PQzCDqml/pMXJC3Z+BVE
NvaEQyLKNMAmml4apKBzFFakfg6FadJiAaFBYxFunbBBasNpNdsELLI/ONLsLzdJ
ZGMrub3O+ARqfM8LmzCy7NYVSHK5sUGv5w+iz2J28JMg/i6T9G1rjpn2XffPkW/6
wtJs3L+YvDyfk7YD7jjvCeBJITYlKdDG4Hu5PVxJQrNFAmoWvfkT//n0VUNHV8xS
dILrlOjuzMjsFWGSvtzze4SguMp2CLgcF5lLGEZLOagxExFd4PXj7kAtGdXG5d1d
5lu2p95BeCagR08ZEAsFIVTEiKIoc+hxmGPnmUlJ+/f7nctoGUGZZ32i+PdRuxny
vgMgQfa4FEHq1qjYmrRCbE8JDUEyDcN6tS7ltUD2KyQWlVT64syr2QOLhQKS/Qn+
5L98tXwyoGZqVcfZzdRJnU6kUb4FPK68n/RR5u/CbDCngn2b694VYZsb1QnVbHfG
xdZTtKaxFqbYYxSvCUr35o0PZfB4ClXWb/QzVEZFse3v1i74EOVZP5e9Lr1HmRyj
HBoYpautCtbmzl3aLoPmwmkJe+zgM0Ict73r0UcJmkSaYYIb8n6LadCnjo7HkXTb
Koe2hnx/7e/sVxtZc6+OfgWlbQgLORvXDuzQtoUltJtpCLvAN3kRpfDhxPl3Ht5S
1/IPMV+sjbmnNOvv0eZP77GfFhk2I6W4GVkzvv/TjlPjMDie8v6iJNhQsOj5/Psd
L8i/yOUw82E2GVYsQka8swMYOK8esdBjdn27Ls6CUMQoxdZD1dS65AElLfGU62Ux
F9lpe8vM5wnuBkDFFxLhTOici7ryCf+yQbQs1fPm1s0th3Gh4qZ9t7LfNJRP65cn
bql6TL0djFg8/JnyIgCOS0jYZ3d0CdnYRBYjOflytd8NPihr2tSboZMrtWvRRZKf
g0+sOT+7qpWhON0uWSzy/qswqu9h5sqtd8tLlGJSN6wZx1y2WZ8BHXExbZWltz+o
UbbX55X5mKVDPa9aTg3svvj/ccCvTehVGsZuzJvSNWZIAisxnO66MMjdxzkJxdaD
GL0FI8tiCMLW8rps45JEkupP/CewRkRD27XWS9/o+auUOpJEme/iXtJcAcWTZ25g
n8hHtHRWWpmTixWtnpxPsGjIFop5o9s206/xGZWowGujrixdUIYxEHsU12fYYQ1L
Fs0q3sfe+5DQ95OW7NrkMGK4XkT+sbNAc9dhCz5lZzoj9FsWKQAcSaPlr5lhVbDA
LCf08UF1dSjxO+Y9BHvOwIoUhG4r8s+lZLBkT9OmFIZp4+zNPThEdvWJpKp0mGwd
xwYjz7v4dQ20vJRnxBC3BbW6ZNLYN0IpvmT8jYfdJTRItwpp4CG6wa6ZQJWnfUei
G7fqdawO3k+0px+NOeQWADYwdthmbpbZDIszEm6lQfF+xD7+Mr8ziqYDemrmHO5K
q3UTxNVEz5N5mS+mbrb4tLmE1TAKDw7KFPbhUkALLXcJaA4996LKCpazlAbC32Zm
nF6UOWWvKmU/qcxbwTJS038aSHLB5Olw05xh/AS2rovSslILr/lJvatykDY92oKe
HEwe3WtWNTBDdOiRR8p5ZMkiGcQQOS/mPL9UhCyZvDwFr48jp28vNGX8wn61KTq0
PY1hU5QcJ6m84OiOikJJB6nedPq5IZz/UDXO6eMEhAYF93EmXAW0da56x2Dbo67+
dH3redmqM7SU2W6d1lMwMHvlKrLwGFUaSxIksCbc4y7WEStfpQ20i4PCbYUlbqMA
qLeJrSYBmnVPf6m7ciOW29GucjYw9pb8Rndhr3C1gfbIFLuNvn4lVHOIlD6gCvTn
xWTzsAkPqWNk2Wk1OtGWpxhItPXSdOqMkuq9W2b91gVDpVx+2qJ31DH3ktgsTxa0
lZ8r600taBF8JGNzAlymOv+eykTp9ekkyggwsJsqQajRJY/zGWp2qxNFEK150vAc
vlYrnqizXL3mY1AC4x/R/cvEfEwODfdRIxLw2wyHg8YE/pFOxgTTnVR5hGFe6eeg
rpJ654N5VyndBz5OUynjzfRn3mqS1bnpDIMlpMjfpHJyoBmWSVP/7wJ/5NBqDvUs
0jV498VhkvUkBWM9+FKvETRnZ3JOPxhiHAZwvRwucutpX8OOkGgIonDXSRZuHF2Q
Lh4OcdyZDxBt1dkHQ2fyn0h4dJNgICkIkcq6a/Uv5kIncVZiKD1251e+GflNRfkS
j5lvyZnKJoNhAUU2Exeaksb/2JJFXQmQgXNb2vyRet6AMwsO8ZWX7xtziSgcJwtV
+e94C0oKNDMy6oGXUnaPty2QRkkgULQDdWAihSjYW3QPPMsDkBdHXXqHZnEmnvp1
PJ8kwfOfhbswWjJ96PEBxJ7u+GMEZYTx7taQ4I/J1fehcl0Mh/9Dw6J0Fq0xUxwm
OjqQGObxwq51wIKFHC3lzhLzNRUkrkg5Npu7nyX2D0+whfvOQVxIcx8YFNnhR9yZ
+4C63a+jV6tWXxpUr/bx/uUsD4ZFMQyXEhcYhgZV8eqYQJ6dvfjRQxTlrCKV7yyN
Pal84P+zvUK/Qu2B5EWgOW9OOJwwL5DeYrc4Dz8DTIEtSsOtWEX96ke2CNINp+ma
hk7EHZUmfve/6+ilkIjxsYDAn+o8NxpWC84ddWePuv2Ac+kuYDqu2nxnPfLmdLQw
e+98eOhB3gyJz5eljO2e894szx2OMeWUhKXbRu6HSzgQjZZt2zpeZ4ZUM2uGSyWL
RcTkUinDCxvQeooWpihs+dp/O1i7NagJHLVeQrNzGH6bhObDKrYRJUMXSVxys6Jv
WwBdPfBp7/qjlkzgdvON7+s8OB5+kpaphAxvGHLYDfo14Xgl6rLGvRONtSHLZu3m
JiVTu8Om9zi6pFDyGW4WFwyhYb07poCN8U2M0aGB3XE3wd1l+dHridw3ifLANYjy
eWtjOtlvkt4PDE/Mu/g7apoxbG+g6GXzqyk1nSNMtVNWhL1uey3fBmxJSA7Mctcf
s8kx/80VnfA/chwAZzSylESfz/pU+Hj0V155I507s34gNXE8Bt8fTiQ57OJhCix6
WbGYUDl/vEt2LMDxULmwiItlO8bCi/l5BCGoEx+C15RWxKZZMYx5iyGbZw8w1XZd
CJVioxZwHszvECcYwbD7tI863AzYGIgvpIMsDms9mIY4IPVSOv1bKxDpueVQCVZJ
VWHXyg/0vPVorRIVQ5NTNKpLj1e1K+KYiJiw65XTo4k7EoK2Wxy/38h+eoY+koLH
vTptHKgJRLSsmv6Eoh9upjXgEtwMy6GaT9IS+qiN4JUqk1BM8skKUGByE/nuS86a
gcoj2yFhOBlJR6PH51pS6SdBL0pkq4IONcneOCZM1XMlxLkiuZU304agZy7Sy7RU
51pTQzF5h9KP30qQF8QGLErmg+eac0JTcHbld7NnNAGyNvHZl//eG0RPmFnyKOA/
Wpd1BbgFRhCTl//ixPbiTd7aHFcNLuVVNYFVBNxhMBiNwkGrFepQSxRJAjas+POl
LL0aPRkeC0WLnuxA1HSy+Ernv2PFlxc5In+uptBt7L/fFzPl+0xGk1feqL69S7h4
O9N6ybg9trbxR+xQB8F2ELgT3wcQRAf3okpyDsY5Csg6VOpstb6Lb8peHnJXhCwl
4PWVOg7PgrmR3qRL/VPo3HhvHsVwYv1oBfPEZZPSOnsoYQENdx5Birzn4ozYndKp
lhkpDqKJCf7f6alu6ZF8dvbGtAInsVY/CzvT3+6vYsBfxKp5jFDTaEsy/ZBmC2LO
kwIjNcnuNT/jKRQRnrhn1QqkVEwV6aUXf38kBL2r8B4ylX5jpwyHQcX/FMZoNrer
JXJdZmh3i1PvhvYJlGJNHRnGS+kr+br3wwCY4pfX2MGk5TUhK9ushi3ZpUsjLI/x
sFD0P0LLhHjqbMuJKUFm2G4NGfqy+dA2mAtGR96nIfZQDW7Wnn94Zlo7lvJejT7c
VemRr29jj55auXa9Zim74pJKHFfO9T7bAh+aFVJEYXyVBZS4RXsO1HtX0tAuKGJ9
nf09I/QdQgb3Y6KMjpFiCWyhyh2dGrzZ4le5qyOTfT/9zYzFcVCic89dLk9GZMFE
87Nju4MBvJPHaIJFi/y8HeR2VSQf1P2DJnMG8Uo22pvDMsjSoymxdVSVHhD3aBQt
PhgJMNyavGdR98saSBRKMQpMgsqfhkcLKvlP+UwDshnWaF/mAGJ64pv+8gs+HpCg
l1o5574bv4jwgCa4FexZgpiqLcJwMDr+Xgu0cBYKq4+ociERAizeVARJ3iBHzY8A
82gGs6VysCdOa5loO+jO3WbUJ9xh1bAcyGKRkP2tKZVvlAH1vMG1d0sEDd6WtCxm
2m8kKCjVtiRUt64vXdZzDouTCTsrg2RBZsejs1NrOIoATVh413GsUoPSZsWztusg
n4DghDpjPo4u/PGWHfAgxiHRTC/pOvyfucUhXW/tCQyDgvRach6MOBKIAWX5xSlX
j7OLFKK7AoRd9Hk/49BxaIw0OO3IGn0tWVjoXD13Y4E5d8Vd1tosjaHtZast+Dhy
FfpGgwoHGcIVNg+JaQq0NQDESuxK3eqA0yy0nrXO/8jC07cma05ZXlcNqSxYZTUR
2zt83zOm6yoJ0eEV+MDb/hYhGoaHBzofqokXQnauosB0Mlw/GHIi/u1Qirfsf9nT
PbPhlPu2mU4m3jrS4oPIKyCV+roFKmc96Ort2ylbPdLtefoXFldlSMWXARcCMxu2
ghINFG/4ZVujiibd19TiYM05ER9765jcMURKjOXmyC6TibfTPCakd/fIWr+UxKj0
vpINBgHEFjXfyyPtOEPC7ttgegzZIMK1bNiqwRVCSBwBsgyt9HTpDWC10tnIgO3W
iSNPIMSRmvX4cKPb75qUICkLQSGJsT/SNbFhlgQpCj60zxeHsywd3YYM0itVwgav
ldA8EKSBh24TYaO4QWqPGDe/oNtM6r2PLmz/vN97PnBV8rVqM/BxFCA+6iyKnli9
68RNNjtLo6VGFNW/wU+vwNj/Xx2Rz0MsrXYQSsvVDf+RbRr0G4go26BDGXj5/hJ2
jYJd66ogd5/oDNbfW0vksUCTywLFpNTTiG73k+usqInTXdN3o72xyknc6qhZDYbL
/cPJAzGeDGr/zZ4HXRJu4ZPQKexFLmItG2NAeplmttdP+cJk+xsd9L/U3R75106j
UW30qzeUXBz5Nw0U4O2nDzeuc/Wwxxw85cNJpXMm7mYFt+86SDzYCQkHjP54gJUF
y1wIKokM4iY7rqHl9bqjuKJ+h6fOyBKBungQNgKQ/55jQkT4ptpHcfblP0OlFqwg
UPzQA2zcMchXz9LORubzOWFtHkH08CjCykcbQfr14DUOpRdnWGIzfZ80vhLe6/uJ
r2WAPjO832LKS7+Q6SngHr0C/Ou3vg0lzBBtG3+Zbl9GDkY8eB7jnQuVfmPcWgIY
QlzG7pmK6roT7vhDIALrwWb8nh7GfdPxDb7EBDypIAGl0MGTXalvvjHAztemkvRC
ynCOV1E5qMvHO2OLG1JpintFVPA/TQV8VJSPfA94LSyJL6NVjoe2MSU6k7Qd6lCt
anBSimugTh4QVTZ5HddUwHkE2WKZrS5rdMPku9h4EOqyk0yW9aQa5H8qNvW230hC
quWLrp3IhJ+f6uFpD50UNTN8/0Bnz2V/wH3qu1fgFY1QerKDND8sWIzYUnEG5DK2
NasK0iMaoFsHOlccF79w/KetuV0s6knYhGPaJxhzlMh2f+ZuzM+qPLfIV1ECCFrL
CR0P8Mtf+G+QMtuY2A9KSrCtJ+5hPQ4oNfiKT0Uc5bzQuQn+E8DTMFj0mpq8C8ew
JMwJ3A89zXNj3XzoC60YAOxTVBzfDi7YhZ6xV2mO1i/nsrkXdVoHo2V1xNTL2uTr
LF70xeoO4+rjmDJzQhQoWfV4ZrCJKyZkPK7oRWoWGiUt7lktleNL6it9cu4vhCxf
C3uk6NARFbezdC4feTQcqgCIrzX7fTfTb+eNHDGSyqki50i2VT7pDDXxEccXenRU
vRdly681U2GYCJ2dhRjLE9rjii18ZqRdHnLdG8Aaxp9CYOsuuLyHGNE6TMfAq2DR
MUxtCGr3TeZf6LmxGaLSw4e1Nqnl9SUUWHKDB3EuCsheVpnuLZzNZDkdPqrlIonZ
u7rsgVcTkNuFEfKhbY8XOUNnW07Nj303g1ReCgLDHrVvH2U9+LwdBZ8fJ4yBY7US
7xBPHFQRCZPOuRtjP5OVU6jkHKFYjkzWhSsrTIT5idhktH/FpVIPL7cjXBAzb6Xa
9AAm2OMydRpuEiEZ/H0RpR3gxTL+LwgagfKQxtX14dtebdRoD3ySLxG+xW67dIFB
1fqsirowNbo29faaQ5UEhtNw7KUOJgiFmiNRFPJJmhIAZCKKQEsuqKHyYbG/gWjn
k/UZXuVAA1vr3VGx6cUQhnsMV4/yrXeV5uSXn3TP4JQz6EeW+agaCG4yXjUNwQCv
ao7WqxKcadqefMdzmmFpNo2Vk45uUrx4sBO/09Yn17UmTWniy17VZ6+cWXnonQHy
Me21ajODervaG1niL+Cg77zWh0Dg69vHBa22gtW1kmtadP/oeCiIUZ6jqbUyL2hi
9Y0oz1Tj645lwaYoLSKb0/4hfaRefbjp1mHOtrgUOky5vK3EZslWOSbUnwtsQjZM
THFMdROIpAigXk4fiJK7Vuo5xRqfUwLuGr63vv/yFAXBwH5La/StT13fpS1W5q6w
rQ+Wol23ErwEf+JN/9NX2b+bCmspe53V8ufHV/hZfhFeTRFEQDEVAE65jWVMIIfi
eKszTDwG8Gx3ulvHoD/k6bXN1C4/EgJsP8dkCRkE5zlZTdREA67CjIfh5wXUfw8e
N7b9DNmLdnKZSbR3dOKDKlHm9xxgpuFZPq82XC6F1r8z+ZkMDeLb2guFUjIPhOjg
WPyQdeTm34AcURVsGti4lPc4dZ877cjFDTzJPQoqP99rCayhSf6OhssYjPO04DOh
8TEzzB6mEgePbLvWrmqENDIOO60Q6Esi5aGGchmINuGbYAVtVFlWTXEpygVR9w34
CjOWFeXkaeDFrUHk2Fix9w4MUYC+AgYc5qFrDCi7OrPt88JnFU5YUNVpXXs53uUT
+yShHN4ZG80arV7chy6AdWuUBQEa4EA+2Mhmq6Y0YfUCE4TRw/9L3be4gb9anYRJ
NDFcrK5LXhUbzdIZNjJ8dVjWS+Souzx21bu3odLNYlU8J+cf1UYjhvW7xAXSNKfo
TgJ7dLEkKvWAa9+xpvagsc+EpJJQIZgDrpbYwTpBONvplP0SzJwivCcdKKHoXrST
iS7uuQqewWWnInD+JtZ/mNV78sZK+zxyfgWR3EMK18Mx72+EhTahz6OQdJwOZNAV
ftLS9Vv5LVbnnGv0wwVF0o3eXx0LMme9qovMzM6Cky5z6VMGuuuhUtL5WmWjbYif
f/Sbkkwtwz6Mf76/oiJOs9d1yxPoPAao3iSTVpv/VFmYDkvITMGoJEqD/xmO3ZUo
4fvHSQx1LXUtasL2WwCD6fRqCk2EIJCU2qrgsOBn8rbkRX4qIv3D3L+vRmIZL2HL
15pRImsXU8IdR2cE25lm9lGC8gBPUC33blvnr8olry7c6ad144saFGvkXuXV/DLB
uI9KrO1U0k5Ov9sqjyshAjEC7Cu97p5ZqMDGdYZ981lRSDzFdU4BycXyOhLHo+Ic
dLwfQnAeRdLbhyzkb0p3PDvkEOx2xquulsEZ8kb3gI91cqloeFtWhR1Ld4cZIJsC
ztuTXO3/QZN3Xjuzzdj3SyXNwyFh+ergzdfqaFZF4d586OmKgCCMIYNGjyNfT/ti
Rr8Asd6y/+h9ivqQrDdeImzpxdesZbNkoWe5EOOLKVYn2sbdOcCKiocdOJ08RlzP
GgY565/wq1Huh1YUuqK6thGVRofdg8/hRo8Q17wQmQ9+aYXLvIjnEXECYk3w58IE
i4DTnlwO5RKnxWXMvqlv2AW9WblhQwbzuYx7HaufKKJr9zpunwv/Ai3WYpYWcuAu
zMSu4B3lIcqDUBc46Pwb9p73WkIY+vP0T/G3OMxdjSSpaFQuWdNv1mr8pkSHvMMD
hU4KT7/cck/QN2BOfyapeM5IJ/BlqIb6dSHrKYbgCB4sfq/1eiktb+tunRdtMp8Z
tHptwCnxmMGc+YqhSstv8BdTEtuhmvadBX41etRd6V4nE13gHWrWx0Mec3/SQuMg
KvswdEcoIz+4W3wb1HL1JrE+mZO1GRKS+JVCuhesznAK1Z8kVX18B+r8CdOIa0LD
ibE5k76UZ8Pgey45qB5ahqfpmk2JNHOp7urtKE3UNrheaQXNTG/s+wivaYlAO2Sl
NF+kJw6lXoBXIbXUNaXLncPdfKxi88Y43T61eZXmFzebHlL/7rC0ZT3H8JdZytBS
p4JCykxVJMFPX1DofG3ya6I34A99Z477o6HyBnzX3LI5w3rxZ/3sGxxMw2kb/LSt
lZM7Dx/sVlkch3ZQrm2XazzN33MbAMAUhmm6T6Ahzvv2rjOoYkNNtMQ2DjxR6YcS
P+c5g1Dpv4xd5l1szGXAK6vHkKRzZdLNyRX89XTxKD8SiMNZnnJyo6PDYcJRrw7/
iaIBLHk/UBaFybC0CqbgZtdPEZuEqt0cloTlZmp6I2nqMJ3oneaccENpvvysboN5
5gkrWDP7WA+fYQQRy6YaeZ61+R0pjuhhDwF+7uDx89rqQCU5DMfpCEL1zztdXRfg
33wrzbJTMYTTI9h6ONWHwUaYVh3Fwj5uuD5FsQzDiwmJz+Wd2x9byFyvHKwmURhG
o1xsNiaYgizn2EoHp9pUmgjmGqj+LTW748i69IyFE/eFiUBKG1wSKDOvjOynPLra
PV2LePJmGlTA872zaJOquJsgn40xX6cn0kzNwO5d+CGa4yDho77aFV7GJg4tP+RE
rOxUEbmdmJLZd5HlMV0W5a1RBk/WGmBgfiaXkDS8Z2vdQrfKHxJEEoKZq4zMZ16l
FL/1gnES4UBNy11/XJONGxx1YXJN+H3wQ6JpJ2T1rp2Xw3zF5quLMmFwge/NSo4t
itRTkfOeGHu8ga99PBZBlCmMvJNc/6EHGXEVjfSbvgSrP7vTfsa6Slmaa50rlnPv
t4AqoW/+0df05jp09WCc50D/hv+PHVtwyQdYw7mpHPL5vkxiQSQVVfAmeaY3kAeY
Wu/x+yiT2EDjM7MaIghzDBms4rDlKwTOpe20W6Wm+nhZ/DS04XIGpVZk5CoYv480
ymyu1A5GzU63tAyZYl3sP/MLFLSpdJJ7wQlA9KsmLEdI4d7JLt0zaQ2Ay9doME1n
B2K/4E5UfCYmmqkBfLCldD2pU4o0H1H19oknB0Nc1Atws1D8IObtXDtGWXhVUXaA
L+9iDRGvGKPJUUv7okQw8bBae5e0KLWfiKLk/9hsCmP5jijK3lR2kYcZ8SCtSliB
RLz4a9HBT2x7ux4eUE/W11Cnws/4Xi1Cz+D5wGnAR1LTyl/XXR+GOHRRO7u1njgF
yw7kjDO6a7fojWalEv+xd42vloJ5gK1+3Omn9zATn6AQljLlmAyfYTt6aB0F6u1w
27694xV0YP2pTgM+5/7SEQnfv2lwL+e2J08aIZp0IUS+QWFTQmN7ocf/5QG/JaVr
Ic9gt6GIAx4ygpyWXQxh9qx8edNZSrBryYlGkQi9+Gs+F8LAaBcDbfbg7uq+HpOX
LKDW4QmlwtNbRGlY6ihxAWps3IAfmMXUScmCfxkpt/KE02eZ+zZjY12RBVK+5bgz
lHBHd1B/07J3Z8jZK8X2vhMosAP99abXZ6zO71qUwJzGnCIjsfrlTNN+NOIJ14/J
eA2ze+zHosFLBVbyebgFF2OPVq5LNXgvDY47fQYqIk9RKZy+TuJUyAQ/drLLVn87
ICuqwiChMhIRMRhiIefS7zUDgQ+II2ykcQfeGQrHfCuxb+qEpZzLs1v5fhN+B0PX
l/BZzyCqwqX8dbjX0sZl/AQG13JVSxmVZRn/Q4F9Ke9nHOg3RLZPlJb9XoHJdoM2
/hYz+uZOBRrO1mkLB7xXDfzuX3ksYVjpVA73dhMyweRdfpsTGqILujZj9j5mavV3
RoxfcnoVU0Bh/WMRSt6hZaJCy9Kyd+Z/euQApWa59FBojE5xNWio+rnhHgzAwBNG
UJxJCEP15BoMPlR310/0jXWWsu5f75aLlnypM+G5X3hfmWvIMZhBd7kgIfFM4TeV
F7nFmdjoqS6adp4zI1iRSuy9TfvnM9iUxxiDm6vi6t3eFUxP/WQzxeCi+ZPkHhJr
/PS3THewyQGmqj/HGNdj5Wb9my3cvDTuWNFNHtmkW7ktqrhYxtzUA86EFL2FhjuQ
mXV0/q3XarQ4BTMlbNLeUgJi6svdruXnGsGQddLReDNgSSNtU5CFmc/BKBdSMq20
JIsc4SFvghOHmsBPBg5EaCIZXhgzPXzjq5SNO2VBiNUn8kzlaxZQOCbwQRv/aYt9
THhwDUZ7kzelBHgokjHaMkcJMzLoT05B9YvsKPIh+ALD033BhvyoCFPuAzYQzXiA
vAwkax7e7KLTeuyHeEjr7JJrsiO3O0BUXcGJJ8WbWGJi78HerZ6O0kmlegv4BEWB
IQqtSaE3IsNNG7v1M0aaNp2dZBWVxKhZTT6DEQwfdcBjgWungqVK0IXzPzD4KR98
Rb6wgjxRdD63rQYUGUEBSale/zKSjjnCtRX3fgMaVW4Y9XlPhP/7CoXw92ieH3ng
3tW3QSXwxwcyb4lXliFQBGk6W7I1sUJJDJK++9IVr67apGmla4KSa5AKcla+VgB4
/dRfAJY1IPNtiORMzzfU3cyVR5WPO325DobGElhV1ygEY46gq5XY0GZPeMqUSGdu
GWFIx4j17l5/M0AgwQz241ZCscU1BwJTJYqIPO0Qm76BGL+VAF5+mEaCFsISzvzQ
kZdpruJjlP/6InIoWoB3Jh/WQ3pjKhE+ULabN7pntw5TYkY78AlYpOck2IWr/85g
cb4Ds6aZAcvyeOqjUkjRRn1NI9kO5eWT2g4+zeMyrxhApM+0Dz8ZLYlkWF/jXZeH
/8flT4IoFY0c2VU6kj9Z9LX42a3wfnwS9pdM02d4bwhgi61foqcuYufjiTkAp4Nq
KUfrswVTdg0L8/oV420owBsyMMAfnjSrfk4C/FIZcyXrKdiGMTd7m6+ZEEyNh08c
ePaabTWuL2hNe3IVfyIQqz5Klo8TcUfjMVTSsEqkhoWDi93BSvilFnYzlD49K0uw
uZFlV2uwjjIULmlN9MusajmzYkNK7ZYEY9CuUqdEA865XCuX8I1hr8j+thTrxI6G
b+C/nvMI/u3i5vRsGhVjwBC6VsR5CmtHR9S0s01EZDmF7j9hENpptJ9k+3zHUPEI
pkMUbsCvTCbIWh31FWNR0rsRM2Mb1mjd9dMu3e7Qi2mSt+Y9sCYPtO/gJI1XDdzO
Yfsc0cHtC8cmsDNsUs8B+SoOrGwnyE5NBhoOF2MA3PZ0YaVfMCbm6y78jBmPXNZ2
uK9cg5rvplLvKcOg1bTI+sE1bK7oLiVGoUPYGN7BlW2TyGKJMmjrtvehr2CPP3QK
lFZzlx0EEHno9SIVdNCXoKfu81ENIrioXyMTcdDG3eUhHHmOOo4J+eB1lOJDU6LX
Moj3kK/ssoFDP/DTTyfROMTorNAqatPbfiZWu7cTps/5Vl3SN9Ya5LA7FdqQEeoZ
y8kdgtcfKcpV9MnDOiNN4DBDrcnAFq3zCJTAckonVA3sUMekp3ZfX69FcY+wqllI
40iye14rmqitiNuU0vYiQP0Wf/Ix9hOJ8IfmPxKeocgYBX2EtWIhji98Lt6+biXv
O4pdrUv0ebRiPHmZzH7BoXLGnnzUom/57KZch0TU7wdLZgfE7Tc/OPWpnsb0Fizy
CazI0nwR7mPscOhBASPrWFiDdFTiwqptBZL6XOlc6BLUTj1D7UoMpaGRphNKjuKa
BEQhi4yCRX+CwgO9aQkepSYv5ZsQcu/mN2Bei3WaQB94xsmuY/BXC5cW6piOkJnb
ktczNanlH4G55sCkP3iYyxdPXrdLgeTUZnF8H7TmwNpTgOR6BI1FghPi4sjVkgYo
4v7CQU+y4HnRn5CC35kvGUXNwG2TeJ7i+6vkDQx3JQZxR03C0dm/8dmQiMKqaHmh
5tS86q4UyuW+4x0OJRlbDQypnhbS3j3HQLTr0WB2dS93aVr2ubf4auwa+lI5Hv13
tduKmaXC+1F+khaWnXD19m/THgkRvYSVTH0SS1qa3uTkDyM6gCyCJ/PmokkStbDH
BahmwPktETG4M/gVVgrL33gVGLjrGQWdep7qaO+kgQGtOgsTkpP527aF00W0V1e8
KkxzpbUVa13d2La/P10ezQLj0953J/2/B1NpEUaQYwF3gVOdVCNa49G7v9tqVXY8
CDvDL12CLETptEjZTdSxgS8rgjGvmo/cNyZQBCWhLqlnyalmWGPOp4D4GFiE4egS
4tRPVDmVOjUJqnH6Old0wvUedx4gknVBPI2RU3M0q7+OFlHWdxJk2+3963Rf1DC/
ljr1HBz/W0kOpvBSdWmVO3lL27r2yrl8StyyhGdrHgVhXnIqxjXvcPbdDds2EV9Z
VBWCee7EudMxx8t56amHdiaUk6sLqoyz/p4ad3l4ibNdvMHqB/k0kw4dUiTn4yhs
F6s1TpRP3yuvngiFN0rGz9DC94DxSX5pdNci/o2Y7WM3sFUhRYaTs58IigeEEFcD
q5lbQjqjRFwoD3nNcvk2bgHs/V0WLUbcOv/6nQ7hCIXgyjyfuT/gS6MHU5nN+NKZ
t9Jp7EYt/tDQ36C6A5h5F7R1tuiZ2CgIxAh5atp184EylCXFmsjOcicQDh0R2sAG
xcpJT/oNbeNJFYuchWlkN8tq2UXXYViWtnBkuR03ryCWJS7ldnraO7vJzr/hKJYA
ow3mf9i1bam4xdaBxoc1a2gcleoVTJN3dhGIZzzCcK4oUyqEza/tqq/hBMrN914w
49J4tjJs6AGnNZrMt7aQH1P4qe4iEZVou8mUlLXhqHs1YNq88Anltm7qk07ZPaEY
iI+uUakK8iH9J1VOruHU+vZpM3HAd4ECf+BtXp5S6TrQw3V0TocaU3OQF327rcTf
S8ZQ50y0l2GtIWDqc0CjvcdsQ1PvVMQcUa86uQg8UvSY2jcVifxHYdx7H2Ls65B/
uo3cY3I5PAHkbHCOcFwuS3xHSghRQAA8hz7ySeTjmGpGLntPwBmJOnJ/SUOjv/1L
7FFAvk4gE+jf4bHPlwV8vpaXFpAxvYf0W9kaRFdne2eZY8QgH4eFfaDkRxjbbnWH
/yWbE1GTaQFVIFatZ8NMEaA4j5V1EAd+1DOa6pZ9btM+tl12bfhRJi0ixOy4MS/m
CxwvzFHc7+0XdxCIpsd+aYgxMrLxTil9v7Sz8BxEdAZl/oTKXT6aO6ExH7kICxWN
W2991yGzj0bvrJievvSo9gzDP8vHQ7CBlncHKWsjciIbPiptJpvJCrbFHJkwmZlI
826gpy5SR5s/YWJzCJZL0oBppOpq733Zc4PArTmRwQxzn2jryNeU4Km25UJGTRfl
hR7tKNj0l2f5/X3O2tCHUGHaVDTUx/XpMptCcRRmjjKW3gG2vpmNS1FOHBbOkafN
qW0Zf5OvEoHlgpc/dU5o2Vhxf41EUmyAEBbdiIrblr5wLy2MgY3aMps3cimEqWLt
B1QgTfzBMob+JMd7SIX/3dghf/LdjhkJDhezoOEepBVzm0JrjtOvdOkzxPV9yR24
DEXGiYl/BB8UOPaaQUx6KGf2UbLgeu4JjhyBhvRf+S0kDzjuxavcyeqNv6grPENM
siLQSWO0pzw7gqhKJW/jK5FrNJUAlp1G60SHofx4BssB4L8jfSEI49V+nTYig/Ft
sAIBacUUsH0ZsOsCUmc3FK8K5xJTVVz7XbkAotSEqzNc68459oxuzHwtKGUSSREv
Riid2+kzvtH0LGnuxunaQH1k19TZEpBEAWsb17N6CFY7SWcPUmF7ljWn5OZubuWH
qBSNet1npswgIjZa681FFo1xuCSwH0XQCNCW4jsjbSKize0hklzvkbKWkHGkrxt4
qK6OGdoBpyeIJeCqA0jfVpc4wmi1B43g0XnDKpOIyWc8c8J9hrQii8N70Wj9bdfy
5YataOXLJjzsZ5U84fOnAK4LxsjgjS8qpXDtuxSJ9ZnMW2aDMguob5Ua9oT/B/ky
L275FkO09426WXVPyr8vqeUn6PDzlYBm7+B6oglbaJATJM3WtQfDYNeuwKIkNGhR
wqUB3IUy1VOextAsyx3eXznKBZ/pQzoWoWj37vga+hSYWj3z+tnfROk5qVXtSj55
WE2TPJi/6e8VXTID968WW0OVP9rAbB9dJqYrhPTT+nxM7N4+EzOTFzZjgG3Oy/t1
/YMl535FAN6ue/vKfuWSNu7wJWusB5OS1y20V05bmp8k5W7+5VPYbdSvT1VoW4AL
BOULbMHgF04ElLff4ItKxRGNjSziRF81kG4hsYSH5i/je5eR7MWLuPGNfjUAMYvm
cFz6iXH5iDCp3myQPktDTHM1Loezt/RTAbjzzqvofjeOXK4UfKSXBaGKEVeh0/b2
pXwha5e01hwz7h+zwEnmc3uID0rGDKQ0yavhuOVH5zcUHHM+gM9N2sEbUAYL4BK3
uTmCPhMDDeIGO15XcvsY5uSTRoJiDsgA/rWrhDIpDninMGfbiEayWkc6cCu6VctE
zcKFCTll5lwY/qZswQviSuSupLOqbUumt3m4HN0ZAtr51djCUPetaIkYj1K329ph
ZpBVFMrUwCgm0qMwX5nQt38DTqpJtorNjPIbmyASrwdEL1Qiz57gnqX37mIPWyQi
OwJwXdDNRl2/9mhDpyjrc1TERUq9II2VUG6P9Vt0LLHmjIbp0o+Abs4vPyR6uGM+
ZfomjfkylX3stJ+P4sD4eM+OdTRXNts2Qr948mc8NDhhSfWBuSuT58uvooWHmC0f
6lAZcsC+v8FfmmQ4QLvV+rEHUy8aEVJCRpXh0tXMvP74Ej4iipvrXwV0HHM86i83
Ud2TbeBjB3KQ05RaALTdBXpvoQDe956/xvX034dObZxXm8NFVVeHG1aJY/Q45M2E
NQvvKoaEwLgoWfaPICSebT/C2vNE+gAQRreSo20AvyU9qjokM+7xyIAiIBUnXT2V
IZh/Mw2AqaTRsEvJDA8g9F0BLePU4h9K5W5SMkcSL2S7GbeBWzfyQlC+FCaI9Z0s
kXXyMgdVzCGM3hZzxE4193f5waY/m84bCAOmwkYp2wYIs0oJH61XBf9C9b2K7uI2
dbqS98DZ4gimLLK/2uG+oxEBWdcMSJPxa6Z6gY72T0Qgme5MgxdkVDVdjFEAn1v6
xfrLauvLkt+R6K+nhaml/vJFAXmt3fU3fMt60emGhe5iQ/8w6hdogtluqOyIgOjY
+UM1VN5DJ3bUB7RQ5ghR4Jqk+qSNnD8FDG/ne1yEBp+Gli0uAyDYjAi9FFg/bR0F
9a9R9tT/DkpWn60Q8WsoMip3RJbhtjE/gQx5Haui093uHZB1LPIrJetUluo/Z/Me
M36Fav3ylo1qDDgcVX/KDFwAyIrRbX+aBj44x4Kg3ZefFkNGyeAKRYAmWpbmsIxK
nK6dCjdk8Gj/gU1+OBllVfGgSml0aPpzjydx/TBm807yvq474T08oC22XbTzLZSn
9QmWCmS/tOzqjPtonhkjnhcQJ33bVr8J4MfBqdtAt2KB2gd5DQdB1i4a3Bwhl+ni
p8hYU/u7UE12ji1fJvmFevm1zlBmHmp0DOYA/59u1SwDUnkcKz5ds6oTQGXdaoQD
cdJLixKYB6gQceXrM22ucHltvhfkdjpz2EBlHSa/KZ/jHES453AfujTHf1EvWTrV
KufnousjeA6FTAeKcLdgHya/od+GOiYX5RQSuzY5Tl3y9lethL6iC0KbYEerKej6
yinih7qMbVeKXZwv3CyikTNGebyBE9LkkgCqQWggX0aP6QOLvG5oNNuF+tarH3Tb
7DyQyVD2Pqojbq2I+tckB29f7rvwNNtoUZQ8Pj87UwfCPn3gYgj6Mp9aSBz2/evZ
lU9Y/wQXzDMEy3bUPRn888Cpb3Qyyf1NyP3XvjEYmfRGGRMBlwdDyDHC8pastQxZ
OZOujFSbdaxyvw5rZKzJ/+3D9U29bCM8LB1Qc6urH9qd9A+KMgFFdtXbWufGOn4C
bUNnophi2qh7+49hsYQwIqxz1uUO0nrqKpXt0/uM8wXT39+x2tlC1zKAO8KDdzPk
vB38HZY2Nc67T8JATSvAohvKbs/R5AmoWE0D1k78OltHRPQQdSczgm7+drq/wrRu
GXSg9UCjIVGGmMciRe9pmveX91QjzH2pWE+by7/CsXKiUd5jSZk51V7ND4PPJIoT
F9nUM0jGmnze9vAC9MUf4DYhygjkUbBiretDz1fu6BePZqc0x/IrbFD6EYAT0cry
EMpY4Ydkhv8mheR7tc3x6JikoMjxhJllkzT36lwqKAjk2viYv1JCr/dgCMEgeqwV
gJf/RGj5Vigryu/JkBShYr7ztGzSY1tHW1QRGzGm8UFes8VRCHewTJVgLv26FRHB
PrEbfkwsHoN4aUVXh1bwrL87U+j5SuaHDg8uOsbQabXvHooTL2xkzuF8Pt1UUqJ+
r4SB89uOf9aMq+6PLgTOUe8VbYlQWn9NakMS+VDhT1zdGzV5a5nBKy3VzXDngCj8
hkPwbX4i4Zxhb5tkM3iGXm5NY9MNoa7GnxA/orEYWoWjjICxCb/zaKoiulz7tDbP
fjwfL55HomYa6NGe1nep7uHiPRfaV4r5YTavqre5woyKS8hdflKeoyIzCHQWUmLV
o9A3aTsjDOq8Oj352UChqtPar4Jqbin8UW73P9vUQoOoReKXruXnag4UMFaYf2Qr
xIhWnxOZltW6LgnTfVyMEBvp83cFLlB730o0wmI1CFrDICqQCF5Eas9NFiPwUtv7
dTipxq9f+xEHtsqneyo2jcAd8RxhpijEEepsnddiZqDUCvVHNLxTbXew2RPggJOj
Vk/AtV6Wkui6YQLmi1/nOPJxR50VV9lHe/iJibQDpt+NYc+TNyEkwBGFgzm2F1xK
iQhH66dux09W8ee4x2RDR2D2BEIvqabCntktL8PqCGEWDjw9is/dhX7aalScqgox
z456epdUnhFmRQVB60spruKYZVRAp1dJuBmD3thuVXOVrI3i5JK8eapnWTXeRMJz
5yAk7IC18j6eLCdYGeDoChptg1GkjxFk170FMcUjid9pIDbmvARn69h4uS9Frfyw
sULa/5pg5vkXcOh9icI+Vjo7Gniu6m4gQV3i+/TXbSM3vHKxeutZHk89OgF5VO1/
vM6r0e4KHUaViEZRexOFPf1Yxd6i6o3CD4UNyKjPrSmN1y/LtX6W8/bSLXIV1//a
SiHmcYc5u0VGbojhzbVuv5VcTPJGod/qoCD/gSV3OViAQLLH5JYWfeAerI7s97Xq
+oqwhIo/p4aGlpp4sk9z2KWJd1cXXPDqoQd1eJHjVVTUieQWTXtHb0sPL/nz1oH5
J+9KnfAa3jbgAzzBufR1ZSgTPv8HJBW5XGkPtyRcQV930f/ApL3eqoDXzKWNsHh1
dRskSY5FwfQXAfQyx8lM5nNGLtCZdTrbMlamqCvYJJXLEJvUWQTv2RHUMRTx93GN
JMEi5nnMR6xdjg4Eq4/samQuPr2JAcqp4Mwji5wImFuD8TvFV8/cIPhv9My4eGh5
L85fP/YPq+CKSK/oFHbr69GSQXmNjmLPW6WD36QWNEYlaVWakDE0cxvgCW62RVZs
qYWn6x9wfCFSl8tv+qZTQbjzsh85Zxi+fKZG6hCPyf0DDEa3cTvODmqELP7Sz6d3
07mkMKRVH8f1Sl+9nbDQlPndAJMX3hYX3r3zIR0Hk2qTjqagfoVB/b7tV27dQBUy
9R+d1SXNQQvxLdp3lo1TDaRqPxNY7BGIlY3ISBmzDP3UcjznKByOu44R2hZquKQC
lj9XA+GS6Fr7D/m8wJA2u6Wu5e6Dc+clTUXPI3QOf7FoZcTmUs292im8LTnT1u0m
SCPMefR6CY8obls4yW6tnjEeVgiKdw8PyEHv/nL+v0rev5czLWBmtC/xsYXK72tQ
j3Cjh8+P1YzQsf7SEarLXKdw9KoYFLJMSt2KDQpwrNBwtHNwq70jAJdLTIbsff5X
0DdZQFKBno3LlwySUPbG0fEwSdLFj1VWbG9e/qU4n3na1JM1/3SSFblgxDigpuMB
6XM8T6uMgIvv819zMS+ddv9QIwP4T6EgEIzzhDZVHEovMqRwgDK+d/V6A7vj9y/T
6TKxsOyQCbfhfsCTP52LtNLE5D/JKzpinofGqUNI8KXF/1dXWy1uJEzpnEhBGoL/
6z7ciLZZ9M5dX7dztMBCMpDb4H2YTn8trCGXLL13RbI2eEYltzp124lmXe71IOLJ
qYP5+00ZDrnGk0O8WI0Svk4cHKIBBpARO5nxvSAvNLhf81dvfpFkEvg+3mU4aWmX
GlWljObwTRVfgCpTSpn6wjT4Ea4Ogi6RAstxmHSUIM/+NRnoPtzwWn9RGnkHomRu
LBCME4ww9eT1uWcel01r0BRb2nv1kVJ0WKx2H6+L+cUSa1p31zFu5+W5ygu33wSf
foH1VyqgIMt7dFJ+qXFMRwYuZNaSF/1fqRDUi/wqkd63qSGoFUjgNdLbzuMUrl8H
OgCwfaPiLcfXkSsA0MB9GsqGxhqUP6g2QbQRpMYLmOuEW1VjTZnKkhvR3lR7ohnn
fDs8cVzyaGxCK4hh/yzLcXGbEcyyqH37ZjNC5vLJtFE5XYbbxr7q1aTNRjks7Eb9
58iCzGpvHCeEaf4lb0pNtRc5/hm4yPF87TuUVOHIUnWQSPjJeTb78zICD9KLinLg
De5x3icC1FYvsWk48GvD4qQVhvTCFUsNYed3F1AWyTDY+u79HO4wEiHINopc1ika
3GPWtnHyptZnKvCG0V6eMbrtoSuFBTf9FhxfYRGqfDi8qwGpZQwWNQfkwBlIq0ga
QlwTOJPKM8DMoitHZTlJrr34rJGJqhf0X03xaQHTbch0QiVB8i09iT8VqMTt0T2s
1lR5AKYF12vkTD53+LpOwFxZ5s8LDmuNdDRPA7h1u0m9lxzbS+y1rX8XjrKndIZ4
BT8BeRR2ZOwmKqAQL9T1uukQ92NLVobaF1AILyLcG0PgcecKBD6gPUisZvT5E6qc
KeFdpSICUjAl4IPqv8pl+tnGFr7p0SgnzQJGj4/qaBW3bi0/g4vNdOL+AhjWRQyt
PLHWUFcc8Ari84QB/5nuv30FP29SVmeWkBe8tqnlXi+XhiYuoVI1oWLe13s/QQYl
wSGa9V+37zsH5gJNezYR3OgUKn7puT9yMnTBKUQoOD3MPoPB37lyO0aIpZYYDwe/
dn5kuGqi6McuiatMLa8J+MmIje3Scxh39MqqK5zxSK20TYpSZkTQTOox09YlP9il
smU+z/aPw3CkVtkxaBxH06txiVKtpJiJAxICHTUVJglWAYajCUYYATKQiyJ/cQlY
5Z8gTTaSomr8YrrWrzZYMP97u8jCwvnzcadpCof7IJq0NvBv+ALQhbTlZtgM+CzL
FmjoPPlKoPAMXAPn67IbZUxJhsChkGp7uAdZrBvBvtz2lIiLEXP9nmE2kbYIzPUZ
vmyLznT6CSO3zyGbBaRP7qmG+hJIhD9E3H5PlCt1ai6t1Hz7wDSzPzc3HrWsWrPX
9HP1EdVm4EBO9mtxjfc68DUKUsjO3fN1MzZm2IWj6USnDkVKeiD90WIT6W/QHdi8
Rt5JXxfRix9HH/fo0C5dsG/2MLfUNfckIze4tkhjxT7PoFpEuaH600bTSgqW69ei
Zp6NvxNWIlQ/sCBADs3/vQVlY4NrHHJSfJjlpx72M5L5uOnVnaCNX8vGiUPBWhBx
0kDSVFNdXJ44udzgIULW9MzeDtnL5/0oqZWMZyIcrOHWacWmvlJo6qXsCM+/EacX
W8emnBLj0Bx03nh1/tThjx1HhGGN1ihGrlxfVywoL05mPAlLwePwg1FBK/4HwT9Q
0B5LJO+pP6rtmPGC9dgmxZB80A9/ih69Qx3+AID1JhpvWlxHZ1f9/3pVfAL3xot0
MFbL+1kgDufFxSJstBINxI9eNNrZ5IAnzrGrA7ivlhyZ/BHv0EHnO+XkwHYsLkhM
m2IMBhJVn5Kh8c3BgRvmKP7dkuPDbRcp0lara6abiBLdeZEuNMwI1zzA7Gsu+NYZ
s0LvWA7ReCzsE/HViJo9cyHa8kLweox7iSlkPR6k5/o9v9lOm4J1zwSO4wSx6Gi3
a1GY02Idkp0rJlNy0AXJLhCaIkQfMfeNjFdbLS9F8l5nCpYN1zeJwawF9lGPzVaX
v61SjpOm9d2hu9268fZNqXLZDx2DCJPghR3GzKpYr1ZYmW7IHulNEHxSGCjvMqtK
XqslPWHCH82hIdVRSbzEYg5Wo459Wu4sYXV+gLpK4rudhqXjKdR+fTmTVj0B/ZZm
JwzdyX9MRXJx0VbKWK5cJHTE1dS8M/WS72TKIrs8LYnHHW+i8EnUXogM4FFl1YTC
9yurQnUFHAmNLHY9rSOUGFT5/lPoJjSmOO/RIjn+vHVl9JbonLqDstRms/J33f+g
4AHrQmwq1a32cgO3CgDckRMt5c/y10tFR1ZHDcQqHti/taOaqwXLevwEu5nidepQ
1+F1I0ezIV9NMN7zJn6QfpDh1UUKnLEICjY16Tli+gBg6LN/ZBFIbN9YBdNs1EdR
RxbZ0KYvz/y+wgiRJ9RpDAbawgdLSfk+SDBjKFPxf1g6cTQlWSI79DEHiec0obYy
yY/l48RpqOQ1pxou2fXGf5lVTw2Xb3GYLuZjwkArpCtrGQMvYeHYO9dTjroANc5f
GesnRifEJJtU7WmzPosHOYizng7NQMvMC8QoKyG0axZt74CLCBpgIaZfQxYl5Z2k
nuGrCf1N7eDp/kjRh9rf71sdXldCYbuErzOLLxTitCpZPRXZ0ZtHPZd9MPOsPzFQ
rxcmNsvfp9qA2tgcLlEYu0/2yVJEWO7bFJS7Enkh0MAgF5oTrPxlW7o3G2s7UZ1+
0gBTXN/5JRf4+ox+gPcMsqleqRDjGTjrORh+SB655SqNFSxI2ocMBft2dl8QxxQD
BNqSHpr0ZC9Z2NNvTj3wpJiiay1YY2NX6BOrtsLnIOUSpmtPyJmC5rVqPRCgGAI1
+YUht5LjIWwSsv7fX7YDc2SdhAtTAJ/2rg8NBQ9clzew3T0APtOE1FdZ1uzwFLgc
PoEYxD1gwg5/eX27hkqW0aB8k5JSKPkM/T+mRBcIxUgoXKLXmabe3cv6mml3T9qR
VlmYRp6TN1QDkxPn4slROEYH2cFFHLSWSyvXSq7gxx/e8wOd2sCwpW9HTCPPb6ny
duhhtoVvzPtq1lKnoL8g0YAGG7Yz/g/Vf2w5aHrjXzIJCG2Ir7nQdXn2OP/4yh8p
XZje4dhLOL2Ww3Nkrsv5HqLnUcSl9GRdio7acm7bYT2UoQ8Dfku1kCXwmYyxNQ2U
3dtxLsDety26udFfnMhcbFUf3hvQ4UCFyl39DwcrWpya5gk9UAueJrcJMuzlJDgt
YUSgA7hcFuuQeAOUNTINAcwOq9cn9JHX4dLQV12Ixlmv3hXTeIQCJCmbFhb8m+fW
iK5FMFJqmPlPifEckRKiHBguc9ATrH+M0CArG1VvgQxBFv3rB0hloEEVt689m5Bi
B4toBKR2fGaBNY8cCBfN+7VZma+P2IAXkI2372ka5QrD6QN2NgOalaJT0+zQ/Ln6
gAMu3qfceUaI+AUZYUMw/hfkj2zumO91Y9SudI9FK7K31kE5LUQbhFQH1k2ISxJQ
y79huJ+/2921X5sHmqjLnPMP5c6BQp9B3SuCHhtZu+7CZIRZeqEHy/CgyaaA5wot
9CBQ3SMtWck5kj0eLeD/Ngoo/Hq2PGIPP54Jq+4waUsF/9vgETgsMzCR7oj1cH7v
wUlTOC92ftwkNPPVzJhxFBEjz5B41GnnSWZp1BFEtge6gG0HjyvIrTTqYZRR5ZO1
T6BaReb12oWLpEf/lwM2zaY4/LREokj7wBkLdyGBLIGD+axMK/O6qa0p5P0E7iJH
NgUp1Jbn3dVTEI8foDslvZ+PMZxRfeCKMMY4LIN/m9uPVOkdHRuPXi9Eu/M0NDUl
mtYpkg6h/vZFxwx97QjKPk47XUyuVt0HwVagYTVD6t3EudS2kpCGY2z1nK2YPsKy
9zkH59ePcmw4j+zYYDE41uuUNyw/z7ipm2RFb0wSJtXQoeqoSy0kxkLsn5HjNRXx
Px8RcBMTZhNNnWb44nS8GCGPGnIWJq3ZJu9llXkcRWTF2P+y85AEgHadFv+YTkVs
XwjpRvRo8zsoAUe+wjnfG0PO360UEPjsI9459+4sl9z6ZERyU9WdbcvzqRsf2840
+xhyVz25cg55sFU9xQrl/zQ7rcZ6Bj3VsA1WV5PrAzaEKoESLvRLVxkXYOO1EVgV
KI5/eYBbwG343qDl1ShwlEJxOSZqXo5NHTMTNHC8NeT+j4J3OAjJG3IrUy4stvUu
kb0KMo9E3iy+WWnyvPqIZlU2yR0XG+xJGae25KesS2EQGNkdE0lWsE8bhSa01T9F
rxyDgrKSqTCWGuE4MndedKw+quVgxDjXQuuN2rudtDZm+WbKc5C/f90GEMVT97iH
Fs1LvOq2b0Bm4QDz3KhFLOND8OLrz2OleXROnnkNLSwm43NX/dc1+u3FASnlDasH
8CqRahe73M8iVtYKnfI7Auf1NeZWFLvT+uGoEzUh91lEKQ76mrXUDjzB5XBy5q8B
iLq/y+oE15g+uqpUw10uxx+8Zs25gNUFJusNSQtv212o6eDG/IfRtaR7UMim62DH
Tv5lbbmljCvbYWlOs9UZPufZRc4xCROZB3BzZqu3/plDClPCrgcFR5YFaS9ov+3A
BSyNI9HrGpG8rOgl9Vg16ujK1taMWiyVL8JUcb2oVSWvc614YHG1imq5//S/lLHE
l7QDY02/UjiNd5SZai6LNyRrl//35Tar2xIlV9jK4xfM0WHqjxY5PPY5dIHlpbxK
aFPc3b8JTywbrgfD4SXAg8Wv+Qn+4IUQZWvlmmbcKZc+f/EOiBZpQ8lME/dc2Xwz
8rMPn5wTu0k0gZGMp2EHf28XbTs9loFt5FxzNVlEqy76ElxeDF87gr7lWre1SnYV
i94tceHutU+NIRn53140Nn9M1iON37+yKW+A2+eAdcVf9AVf0Y8+RjKhE/SL6tlm
j/rbR2XoSl8QlBc0tBO1JmA/BUzlnsbSwti67PxYSqLqDJAWhZ5ooTLhGMVzi76w
zDS7FjLr3p/98e6kEU1lmxUtXckF3pIKxFYteMDJx+f9BHFjVtoB9uoYQRDR2jGX
7yhuQoH/uuVhQ7PZ0s0Zt0d+mBRp9X00SLKgY3lSwgy1pTZsU5crnvbWLZJxaa7U
xV+ph2tZmYzG3lxkTi1NgBgsDlnsviRf9zlLqOEPlYo8x7eXJ9HRwciPLZ9jXnWz
y8DoAKo+ZFoIJ4N07bT0L+Gj1hvkC1eviaTdBlOSQEJ1Rj6FMRnl223vSRaFdMH9
RNtYcYCJMKFtunbmieTNtWKdkLYW09beZgjSZNC07bJ7Vqgim7G0Y+useRMR4cED
Lhb77lKQJPyFlQyQZIvLAfd6Pe2592k/E8OKUbY0CROo5timnlwARiVfhEe2Solf
HlE5v98H+vYLWPEeeygFEmwDpGXxddh7Qi2FalOuJqRw04CV0qFhkZYpMmtBpwS+
71s/4lKXt2XzHhn5GbRKTARM+B2r5VDYbIJA6r52rZlR8033twoXhBX+Ym8Hn9/3
WuzhnUX9uCCiJpPhtNl01IxZAwSFycrczFjpb0DtBK4AwpWD/BilHSEivwdkSxpQ
aXOtdVbeTCM9xnpUgcIpeDy+4yNNs9FEZqMjRh/J+yuI/EQu38SmLGItysJdIeQd
0aPerOHuJ38K6EHnsxHRslI6MpT2/Zc7ghB5ARwE5gcHBTZcFOjJwUvo+snpBngi
b1RRT10d2/UDyh2cDB5DgECDUtEXZ2hVVfMAynGZIK24pjJxGBvmmdqyte0nshzv
LtM042FAd/SnJykIRyMshpC7yH9w/Xn/nA09keub5ovP5IY29xpmfUD8Npq6FEyQ
3NHhEfihN6U6PMjyLr9OGakVJ8iGrNYM7NmHdNkBNxgd77v370UWS+zVT2Khs0XS
DhfqTYSW8g19A2JxYKaTMWwWGkEPXE9DqwDA9BT+s6TOgYdH6/A04d94yygFwGMJ
bhN9jV8sJZnPJG697OMOam3BaIG9OZetoE/aUFGEF2b+35QwYiCuRuKJ6GOSNPwD
8A8rCOwaGIn8PPuXHpG+jONuj/03p+lf1Uxpd44P37FG0e/lp+j8R5dyyVzb2r08
ogjwTzBGhSG3GojF72L7OkqrD0snkM1+gOyhKBFreXZY/glaHrvSnVCOh6Sf/H7e
u66LKyk2kP54s/6tyPAP7Vo9MqNVzvBVFPEEmPucTgfWIon2pTbZMFdVeFcj8mfO
2vTUSHwAOYIjAvMY8RZ8SyFEZwvS7X49hwX5bcl3rKQQZCqOc7fCHrBzpGlGNdSR
BOn4e2iOjEGtzlmgxrq6BsgsOp58qZrIOZQ5HnbKRXanXA2salmdyDAwxOwtuXve
bUWRxX5UTa8jDmk9Y0oLHMPVDmwFcQ43yM6gZubWbX6hD3We5bb8ztH0uaSGHK6J
I85YlebLc+8MHakYQLwS9I2roIIqqsXPn+JjtNXNgd9cpLcI/+om0YX13Iyz/378
yEU0vxhgWHJ2LMDPMGDg1dA3fAVDI5jAnMLTnG/aluz6qqWa1zXw2d1K1/9h6IDS
eWC397OrNNSUSzv7MmydJopVT6+ON21YgN+jaZzeDns2pq8NJG1szSgJT7f4QICF
pZ6ihqjCmm4Oaght5zsN6SIJAuYU1Q3rqCC+2DFzI8QJ/WX/iBJzL4d7JmtrtR4Q
EgocaYSy809P8TlQVDVXb0WrMg6O8Zrl0x+O+fOkccB98E3DFiHqYRTK7DKBbPTm
Gvzjs2nA4I0QDauwLFtvpJGyUpAHoHIbrvwW/BceezvP7IQYvXY0aHmECZlHaHbu
2vhaUipOTYvlh6CzEsgqfaJTpVMiS+6bziHd9A3j1Gv1Y+uy8DjP0RdG+6WbdJhi
MFxRyXpzTopR7vX7ZS6yEUjxw422MF4T3gq4f456KNrAH7k52wX8PbJVvGv3Ay2Z
9JRkFKYQyXlACuEmyrF45/IJg/ffzM4AxiBdXZcxq82oV5a7fiOz9BfJPdPx8DDU
EIt31pSrBpd77Nz84ZV14ISbhsGDzN1Ya3PRNX2+80im0aPqyLZU7XJc5rbR5MaU
BhshB/I1k2GRjlCGrZw9C3gtMcZsVR9yEDq9WaUeQ+H2uuTIdx/WfQK6j6ojlMpg
uLMN+r1Pfp2kmVOLNhvK2ee7z3Lqcwh0UEiRrIYhoNvUSmUAuUB/yxH0RBJXZl+2
CHzxxyS4KhR36khooiEmSeLnTO47LeT8ZKFpRLnVJZm1GS3NLxUehv4z8S8dpa3o
NYQPu1nYNjj0ZQjAOUKrdgKi2lVMfLuzkeuNpM0oU0ZDKcBJf1m4Ou8seWA/LZPW
wuPzudUmIY/oi4aclr2UPYM0cdtVXCnMlKzuGC/9rrT8qyVfb2BZHdXgHwV188QK
83ZvQP2VsOy0xAYvqeteLzk3yufvIXOlNZFodY5qkOXIQTNE1Nv4qqdolqqM2NH3
Ci9JYFi71pHOgKtI0bnvUMIyUF7ub38IEkGedGqyPcKmkqSgvlYorzZa6+QVfo76
sYRa3TwUc9T0E2IzQaTnYVKIG3//wN9gFRcsYZcLicBo8ZcpHFOrw5planvq3Rfc
qzCtvY44MECQGIgDlrRgI64N7u2536twC/gnY4aHs5WLbqjBefTa49TwW07Ie8I9
JcoSDe5hwJ/nY9T3vrcOgoaMGNFPZvYrKYf09hC/hkE7uDGc0DicnhxRHXA8mm17
bCuI9ni9oea0ABAip/oTrhqlpsrk8h+T74eWRPk+bjXXHWJFZl6Je0CFtBsGekCO
4Xeprc39GWAGyC+3Nljoz+N4tRY4DceL5voL+poGBH/83K4na/IdqjZ9hhWE0KFL
2fy+/w8i42X8NI7Ld7mMLrVK1YpcpqiNUXCgYvhP7FZOaYG6KZo5UavRFS0uzM/s
rwj7U3Y/r+HKgFcZcPWutq7va0GXAy+Mxn38Oi7FxtRkBMkicq6RlevH6rt5eck8
JYuta/iZKWp48erEDHbGEsyRwIococKC8LkvZlAbXAbY3bBg8F8JTAXhO1sLjZ21
fiVPjoG4dofk6Fi+dZnueKuQeG8PX7DZ2Td9tiTi8ga7+IzCvO2ekrHZjoMWaUzO
M2ww0H3wkk5ni4CP1Ql2yQMe6grk2/2+Fd5t3FDZ1laW4dRK8LTy8BnHWP3yOagn
C6myUG5LqubtUELccir07A40A66TzkdANJRgFYMqKB0J76y8+qft9ZgzBN3PH6qd
0/elPf7h4lRVxcFY5gmJ7yyQ8YIJ8rlKHr17gZ5Bn8nsB9O6aS84RBuGcd1f/mbQ
9tr3ta9jNOrXWAN6gfdIuf9SlV0IPIMqMtr9P9oLcLHb1QNm0vj09JQmo/sSkgnV
WhWbCtJQbwDHKpi6hBuc8nMkMiiKaRrQggGN61Bk7FwknJUimeObrw68U5mxB4NR
n8UTUepxz1/rjIBRAn3oy1n+lwoJ6zU+yY5CgCId8bLpZd3QrheEtHNZwpESSLi/
3B5i26aXPxSpkElky3pZcuBW2py5cRtydnFn3rvtLCrsOUh2GgTBVBn4g8j6OF8E
FTbfyzNawZUZDoswRIO1mU+6XH/kopv2kXnUJuGNdZ191r3Uafslf9kP+fWPc3i/
B+sUjcRB8FjrJIBYT/NX+6zL9GEYU5Sv/Qk91QAcZyU5sgrRqfN0/SZmmCqUOTNw
F5LimCH6fnHnxT9WyzrNpO0A9+u1wYnU/J0f5ou0387l5nTO3jAoVeqWUPArQZwN
5hEXj/Ec5/JifWj3qCRImB4n0kngklgeClR7CSQlU7u4tj8SOrq6LAIi4zawPBuI
riZ+zeO3cWIPb+dwGuXukHtcLbZa/VGovFU0metTqYz5xhL9YoXi/l15G4cYshPb
gK0aTMR0FKxmwSDTTxwICOCR5+KfAf81sCeXgijTCcHQ+Pz4AltjyyFFDcchah0S
KZKGRfbBGfZOKt9Cr5MTl5z932Kkxwq3x5Fh6ALzYknR244dYtcEdJfD3un0q7MN
zKA7wam1CX6ySYMF1HCTFmKVUXpqfXnGbmCCNpESgwcvHkDi5mtFbK8RuVFteP1n
ZbBzhjcWqITYrn+//lHgs8lGCGcLcLZhVRzyPmJR5GW8y1U/ElnaubEYaH6hscPE
EcanEI61+TYxZr2ZvLiQucpKgiwNoPs2x+VacLX1cfJ6hVBdvDHYxSzylM+QBu3C
hzOSvZ1zlVnAnEvT36mFNmOXxBNpzvk0MEZxQ9bN5nGQGoteIE3AvJvjPA7Onzac
PKwTZvMRTNIpvC5whri7f+oDZW030pKsF7Rv6d1Eu/GsWhj3si5cYbaWorlA+Owm
j1lf5JKR+peSbmO6Jb0XXxYEbIxxu5fJS8S9NVCyzWVUAlK/9N12/z+2yir+bUKa
yazkc9xmNVmTM4wPsoXx5Vyu6b+f3gfgZ2nBRuvUF4wp8un0lauAjNjcHSndo3tu
uM7GV0ZtFVzfmmjusQpq3tVsaQPRe3+T3mYhNEATJv7Mt2ACtu1iyy4krpS/+4QK
5xjvE0wGR0Th58+CyVTR0sihfhlsiRAL3Pq5V83rMJP4zbnK8rHaUXTjD6BtWfc2
w+eRTrVukBHI2y9UY71KaLeXLdvQYWXMD6VJFwzJpoyLLgcaQYLST+J76pVnjJoC
J7FPwPjjDO98IUK5Jf8diXzj5wpqSlzByHzUdKBnPs2m3XNxdCj/+274Z3JLdSux
hebW4beX3dSuGS7jZ0yDvL5OmtJFwn9FJZnL5AHkpQYWhUv43Udq+GafqKjG5fSI
UY9PHvmFBWLt9NCKYUlzp8pb5woT3r3IulS5nvobnOQsO25ORCvVwoTdTFQ5DEx4
wiIKkkpPjDupS127it+ov2isqun3xfrdjAQBmoe2+attTzY63k2MWfOjMuYNVB9r
VymRRbxg8TTqXXmZmS6xlVvBTW6iuH1XhKNoTJbxJz4hmt8nFr6hJhgcdnmQLjTr
wnXUKNqeFoN28e7fmyxcLdAuy4fa3i29FOA968OpuGiDM3Xx+KdKiGE1GDB8WZW7
c/51u2Vow7y6f+oiTOBaK+8iur9amI1xIsjXU3P6pAnAvbIHUI+o+gvCzOQk9PYm
UKsPh46gC8VQR210mZ9DNGmEMrSQ3FJIKGAwsZ0jkhfR/jh4aAguU6xxBmE9szE8
ff3zzDK8vYuql6Sotgb50J3i2Whcc0jG4qERBetU7NaW6daGXD/UdR8PrxsEQryh
nRgykbLLjDA9O0AndJ/aav3br8i2TlaxI/V6QrfzlQQIE76GV1X5GqhaeyCPVMyt
H72V+gL9/ejkb/5bOb4Lj61NFw6CvdxoFjyL9kR7snxLYn0BvR6S2qpJuB85qrsP
Rhobq6vEDJ2crnzSkmgABx6EHETl8eohNBVw802WDirhGblD1CX5hOrcEAUQzfUV
Y9OLPyZLksa4n6ZbmMtpZJ6azWiKLsERf9e9U5ZOBQwWBNgsWFDrTnWUBzDG75rN
UCDfQGpQbgQwtjTpGaHx5igepkzuVq2EQzaiXYZC6kZv8uIh+/S1k9KsNfcRiPK4
w3mOyWpvtTJCmP4hfeelhi7I9oF0ovMJ+qZoxBYGIKR4D3reAA9Y7h/C88bn3fmI
OaAmTo1nSc1T7ySi6Bke4oRVjWBtw9ToGQ75lWXYb+XCn5HN0pHN/24tn9yrqQDj
LLhgXYKXZrIOfa5xyUF9heSZbCGsTDFilUo/c5MiwVkcP+CDG8KH176c5bBqsWKe
daVH6qn0EleIcNLOMobWf9LfVKjMzv+ExL9fBHUyd5K+wtWJzO1pIca6Ee1FFG/+
Q6YTq6M+klxbDf4LLTW2fGZlV+6MUmmrzpZ9ymmf127mrE5WZbgNpc9X83q6ITmb
xmMwxU0kPJyOx9h4CivnihL0qtv9+mModDFgH2OUZhcJb++RojoZ14o2bhcZ7jm5
B4fJNeefJZ+ZG0iujfByayWOviPvZAq5mHVNRNA4fFXBb9jyljI2PAvuNqZytrm0
E7qbeOpXfAscTZT9sw9JWIf2kXS0IDYBBUEnJrPBYNp2Hh4c4Qg5iL578BBhG6OO
FB2ZpUSj15t2eJK0FSjCsd86J43stVL4TlzGb3eOIPjG77bs2/DNxvtrWKBy4NLH
RF/sj08sJPPyd/P8XAYXOkvRsUbwA4xL3akLUbDQ0d5tthMNCVFfCMrYwGdRCRc1
UsL/qwK1F31N4KOAFrdVc/EmMNOAquLbP24Dj4Sl64HnYPYilJltDPhuFA2gmvHo
dM55373ogkjQYT51IsQ8H/endJ274xacQrv5ufr6FVCQ9c/C83gSVPEYH720B3OQ
GMEbnVUSw++K4BasaLw42l5wArMIsRn8WUSIYHE7hwA+SKSETIH5tuYa5ZYvpjPm
QSCre0gxbp/TuS62FISMXWINJjo/+GacNNp20StJx3lnp9SQ29H2qknrDH6xTYMk
sgwY2HQciNLzY2wuJHa59TLoAZWrP3+Dn6vcZBuGQ1vJs3TNYkBxsHY8pruri8Uc
mpRJ/Gf+dznOFFUd7LTuxLmWv7PMqV3P54rfy9nvFw1OfR8wgBeqmncKzCBxenX2
Uf1bjLLQYLkDrH4w+8CjGfd9IRhbDpbXwD6WHr3uf2LsxEAcNFzq8TVXJDlTPear
DU8Em6hqLotVJ1jxOxyJFw7+WjyGDXrbQdCyHo2CCbq7yHAX5PeojAMfiq+9FRpT
4Bpa8jObLhf1l1/8FrrXZ1frslSpWQ9qvpNyY5dxYBbBNBixVRUIAjr3m4jFuF9R
dKUFCOLAKVuM5+FqpfZ2IJc1vothP0oPLX5ZyghMz+uU41jV+tsdkuByoNDVUCH6
UsGuL0OCaVhhe/BapFbUaGtlTQyUe1bKOIlkQakhVYghh8ikaRBYNwJl5oZLAhQ6
n6km3FyVHp9fJI144APdHbXK34KZLghFWPVhsfkT+GRiM6nlZ7DFqTN20MWCC//n
vvqIIXXqUpBnOXXPXRJZR+jeTNidn2g1lHraOk4T+5XOkeG1TYRYIUadafNqQdEN
Au6vPskO65wt0NVh49+8TTu653KZDcN9xqs8rjVGF/qqMNKabePv4qQckkXh7JR1
KmneA+T7ziNznzCagr7Nrxq2M1n221X4BRrTx0IwQDSp5H6C8B0T6/jmPPfRYL3L
WNtBdnfMRPWSP9d50h7INA48A6t3T+mWRzENNtqm28QlJUK9fgr+yp2eAcu3jOEl
XQuZk6iJS5MI9bTsfvFtPTEJezAMab8MFoPgUWQtNvDCp1OsXL/wQlzZfiV9jcOB
Smo+XWS17E9L/BtyWF4OKnOH00uFgOvqevWlgyEIh3KZuyjvbjjVCMYA9/UWnMOY
aFTR8/jlT/oE0lc7seIMLp2A0UyiGDg6YdMDkPfOnTbyh0R13kpqOLOOxKsyvW2a
ZS5kxoim+3lmEP2pEUQtuxTsee37mr+osa95pO4uPd8VONf07NocdbJj9zjymuOy
YM/zNh0dMe8adx6/unR7VqO0cnPI2vWT6CtIlkf/SUr2dfUxP4Dofkugn/7baEat
KRH5pODy+P4o9xLmkBDAFBKo84KB1Yj9tbFKibWz+KsEtzzgKZxrZnfn2O/sHwll
ZMtnyhIf3u8NpOwza+e2KEcKKhIdjsk0ZYtrVq6RXK3RUf1S5WryGZR2FYA/sMhu
U39Hg/C6D7bzR692gVJp9rSJuGds0nlTPlgwf5UEnU72/4SsaAz/t/oezyQiosq0
NFHqbyenfsEEgSoiorY8MC8nV1dRLlIBYJ15QhaXwIqeNEhgrG3lj/9jGbUiADBC
LhfjYsdodBvezdmnV6DXB2pE58165s9/k+ACXAofijJLMTHd1arr5DZ6H4gFlspa
GxBbNh5MqoERYlpjY2kAp9Q8r0sXckWvfzlvrNL0RS+/LEnNFOmNov1fs/6J937V
VBU7V5GgM+OJaFrxvDN6LNZm9+JSazYqsFGRS5EUvV1SqfepvOk6rkhXRVk75fHK
qn3OVwp0EYwYM3TVjLS1PadaUTPXGAsNRYrbJNttSuZQxaWcDmwvjEMH4JNBsZTG
K4noJBsfiOpAtc9PTOTT45PUDu3orL4CCwB0tkOniUuO59fKH7BGIyOC3ssIBVQE
EDpbOEoP/I3xgoYuXZRXH4NCHdMSI+083jPaMwohNoBZUinzxyEXC+iN2Wx/udvW
7umBOSljAwGcS4vafYyMgSKZI6NIoySZsS2nMNSN3jM7WdVy+Sr2ZbnvFm8sIyiR
7gtfh3XQG3T656iRmA765NnanRphlMKM0iVrRKmSqkrO15UZ5pQgBjSySvevv3FQ
WNXR6qVA6GauRtBULmDMMlQnG7uSpkG+Cp2AaJH5z/9gb8WkyJYWebEDPF/u480q
Da1+/4JScq04vMVtbIiTWa/lbv3k1OQ/jz9NCO7aLCgaGVjM/GcmfQf2Ud8E6W7P
hYL1VcBNl3wNSgnAmVqpwZoOtljyu/pULntLSvJaulGUNkvSVOdexBZuNf3SSAaH
RdXhJcmw6WHo+1WSkKf1xYU3Vx0PpQ3GkLAXrpA5KoqYm1v4NhZ7GfnQNoaeMjJ/
QWWsFz/y/bLjFbRKRSEq+d5W/4WdbeUbKkgB0M7U2UnVJZrwT5a32Dh3KJ+vH6aZ
3+it+sxjyG6yOt+EIF/xvi0fkG4WqDf3PZTQviGqkLL05x92X89o2IcFzQDN+pY3
4BdHzTqR78J9DRlJYbMXX/0TpVESRu5MsHP1FuyKKr5EtIIhSEXQBnNcqinTEQq6
TKiukMgbzERDC/PGqM/HAnUgKhMlqwqdxHAoN1qx8D6JEdYVmoU1y41VuxyATpjo
wnwqXFQy0N0aoEu+68p03X7Id0uqLXdm1Hmpg8slW9ujkZrK6tUTlpQ2jb6eTIsi
DQQ9G2lIZyaaNys8u0GGhzn+vnp/Y3hGxp2VjI0SDw3qBsCQLgXX6K1zCLHFHqm6
/obPu1tm8GTg5qFdxeUzM6LSr5n8vwaeInkSIIbEyfIQVRsFVQxlJVUx5P++j/VW
clt5qHJoincf0l5p3W9SmNG1n4tRQ1/AR7TPFJQhVQ4Vofam8m+RGJApClwkz1zo
xyFeBgXT/MR76SeNfCfGaTpNeiBgtvZQhNXOKi424LzO2Oa55lIEpyKaJa1JzjCV
sh3xq4dRDkH1XDGSJvBMnwpagvqEczcmlXuS5cmy/InIdMiZ2Ff7rGOTXRXl75ih
M+f2FfcJb7RsEYrR/zYAlfFt6qEMu4WwgTkkJ4oI4ltbC1z11xlKGYlWLM8sUIpd
2X82fnAlfZX0EvQaHZLtmptmBfKSxdr9rVSuvtaVN/4ZK2KKgTWzqWNOI8Qr4CCo
3wylWusuWhPPSnEwsTPD2wLGUc9rza9Oy1K4y0FprfZSlvMGY3fOF5DQLSS6Bmy8
ZyBhH9lcrTc/oMw6tXAC6KRlGljaPr7GQo8dWIGZCT1M9v/yUP9J2p+KwFNYYCHO
JxwxKDbk+sL0nG9n/SgGH8oCUsPQFs9qZ0JhOOkVAm/W7hCr3fYhONMov/UjcojZ
Prem7Gyut/olTi5c52sufq9g72id7CBQOwcNBKRSqV0XTUPWmNj5YER/jDOSZ6n8
f3iv1SNXNQCCkUTV1rlKR+L2RdCSSPJDRivNd/U7rAU4KcWAES8b76YiKKskyi4B
TaX8yqPDEIL27O0PSKwEqJBFDhOlogjRd81SyduosN7K3aH+9Tw9CIcIbB4SzytT
hbXr9xIh48V+LJ4J2Y7HbIgPdID3heL8QdjfrLxx5zgJsiONUUGAxuzk5PRpNO3S
nell0VuqzQSdQB8FdNgVvVv/Q8L3Cd/l/SZM7rCQtJGL1HVoCwDpC/GiOy7sGohw
UThztDv4qIJexp02An1zUUCTDGQRsgjgNlH2qEWNrRXUmdMqfMKlnC/yC7qXY7K6
lHM4DrjIbYXnPJVbIo/GZVqMZ/3niv4CFq0ARRQ3YYWpPK2ePrbOdXzGjGZOVJnk
VieV1SwlVg3pfm36A445msK+nHCRuwimJ67VH+9LA98iiam7SLHjuFdEFWh+81iG
A7rUGnZfcseoPkFoGcmMnKoyqgZWYSA4ac3jjV6gtRras30eAMqaE66trGJ0R/OQ
masPHCXkAQqqQKv7oK4d4Qrc4HvWkDsVMHpibdxe4IAe8gVRsnqJgaMQnfHNqZb5
sX1AQQuLZ/4xXuJBq6yP058a/5SAdxlJTXr27Zuu8EJKf5KXQ8UI7Tg1EmP/NWhM
cEV9hkJNSg5BKZYSbLl0n0mkO4JxiKwJrDEfgUZuBvhFrIrIZRPSBYs0FW1yMJ0u
48C3B/i2N++3FAyTyNxJk97AGeHBhhAnK/5jrtxpDwiuYeaXNmLZyCf/IvMAg9xZ
wVmg+q8H8avEFP4Rnw+Si6bsKuW4FGYlCryYg/yFAH59+QIpLl0bIGIJ+wskjG/P
TLvAnkL6FLKUOXiyBnwnmuTx+Ic/IOZD6wE4k3hiB9sFvL+DDNN3SGByZWVLy4o8
60UyJd6w9C880FyhaYytWz0961Kwe/aOhj1sSiuSgGO+2gvbSr8YpcK0RtsEYFv+
LzugdhqAwyiE7py575dTSnLv709xUx2Np10ygXZHnUpKzkOtvdN52UeeyZkhQEBs
oTjYoELWwLRakBmvdOrSKW7Kf1vRLjHeAvZFlPsMdZ56ZBifwLTuBbXfmVM28ttY
0Dtt0eUj9QxZCeAPnUZwqzJlp+JLW4KzVi9YawQMHDw4jfOTPQvjZPdFrA4NXca6
YAVmNB/kgK09O1SPMOJtl1H8Urgw7LWLPuiP7bffzYhei66L2hInUgXyKV+ie1a5
Y5rhUM88QJvtPTgBlcAOOsbis3h9gSv3J+aZmwRH+mOtwtk0ZPl95GxZX2ji18+h
kjvugv8z2etJHjq6JH7zcz64Kpcr31A82oUWXjHmvNwfRBuUUtsBrNBpQ6KAeG/w
WzodLB2Qx+TVuD68e1l2YLIee2aVgKV6YHEa1BV5bSGvw9d0s6IOzPeP1yDqBqT+
zWD5gDlGmcHB66Pj/HiQ/yLpqc4cUDTn/Fku3brmqYTDcpsrMhhvLE65eojdSWPb
aRU8X905gLRG8ln3g9xFeej+aavLgP+9IzrVLEMzHPYyVipacjH+BEZuiUFos9yg
yExPaP6zMjvB9NXoN0/gEPohQsfUyea7oT5+dL3HxRgJWb+RtrBvVDbS71zbiAcg
I7rqXfoM8RpobNCU17nd+ZjjA8L6vPmq3jsZUczMJ9bwERlIQgtfNJyOERVa1rwx
EY50g87Qzc+v3AsO+NBG6s1/rd1sLD8vfxmrYfitXRxzQNkAO7Aq+rlsiOofMRFi
GQVo0kWV6u3H/vyegu3Etb5KIT4RdAklvepEhVW3uQgLJLMHhuYnpIve/rbWD3+V
59W/48++nxhVizsHxkcgzByH8PWdjBpvpbR7IcyduLTwxOg+9bUOkkzYT/e6C1ew
bRiacqufSu+uxuOlNxIhp9E3Xd4SZyr/olZAHN18elYyJH9Vfj5y1YkgoKRIdXPd
wBTfXPyR9nVDDqI18XU//Oid92tD1NP7Wx4231XU+ccaW7Cmyy6xj1wyuTOjUfeL
ujvLmwN2akaVQ9ANPkFCXlytgevpqEcU6uAeRlBZYWAOX/g4mYLvp5G2IgS9sszR
6BXEDWB/dJ3/WxWCGsonwN/i2ZMxt+ZqbBeKQIi9Im8Z0XOc2RD+Eb6AUWfPSrmA
53A/q+G0EkUOhX+Kl6STLJ1oBEv8O/XnwuaxOn3Ic0hG8pVabepQRvATitQQcxES
zb6S3TwGKQzBFCJ1SHBR1RRs1U0SqJcQJ+22XAhGVxv+43eeDai3xKJtHacBWUrD
wIxwb6yKj80jLqWVixuTp3yGiuFDPettYNg/B7u4uV6rigPl/TpoiCIo0gJaiOB8
fm81kO/owxI8WWP1reKDeTbKhRtp4p66ZUStoX1dHp8VCrQ2orpLst/Ne29Qylav
+Pl13kcYIvjF4w2HFmAdD9r65PYRU0abTqCKQMyeTASLtsvU57sEVqOFraRiIAPo
lrB0ieJFxPoKFzUtL+wlm7qyhzEDUbT5pDj8G90Dc+hswBacIvGkZawKycQ2nt45
wIWzPZwGYB4VV4/DpSWIWH+fOMm6j4Z5qyrERe2Yh40b8CqY0VXEaI+uAgTha+Z3
djDWIoWYWhLpyc2SQPhe9NUI30cGrhVyabBk3VEWdSTY0prp9ZhqlEs0iGeuAoa3
7qe1jVS+Cf/DK6yPPLhPYwSRqmfBo4qxvkCmDidVZUcqdSQFDhLcUm8uFjfMmMpI
rmEBjZfH5Vl0uXuIZwIQvBPU5Wih7td5KW0ybyUkmxYxAwwZ0yuWaN9f1RXTvApz
UG7aLtc2cqP+MfWAT00qkPnFfgxJm1lhVdINPWOZMMwusAOUSwUh8lys4ZXw2G4w
RrmSwZo/VMzNk61Ocx1gvSbizHwVRwUL2VSBwGhIntahgZ7cHW7P3FXKBLK+XdH1
pBeXbcVMDmZpjGMlryEFO9i9reKfeJtrYsHHKfuvyNBGGYi+8iRNMgUJuWXDHljO
hAgSEeSO4gqCRe2K5aoqSyHADulw43f2C/qllQm7fqLlmVQJsQGKu9nuvp7vqH0p
ERXcKm5Dulp2/U2C6MKG3Yn/j+KY/0MGsozLmRI8s7F4OSyEXdS3ovCPmIYk5cfV
l8xepHk+yb9BPbQATGvG+Jmdglpi9uCl41BVvSVLhnHKjywhDzQi6AEzuI7jqU4Q
3X8ESMUoqafw+BGd7Y2r+dyUKQhgpDQSzWZIjxRTDnmwMoYre0KhGcQkMlSlq9ZY
q9DN5qOiBJmpGYRc9BVF+oJC28lrIyZlVX0bYj8jYwLfjdzmZ4z8PWmCQvODofzf
0Mv6CCHQa24tqqtJAjeDxVUftbPpJGjAyhifTRjXpxfaTV81WmKoaTsJL8UHI8YH
mVRL6gvzX8IozP93PNFvg/ICPW0eNw5RTDUTV3r/uUVSgJ/maWypbtkra/XS+swM
BG41KJ0nKtStCLXtDHav6aOh1QLVqzKTjfchbxS/IhaRhjbarO0CAgs0hqSUMT4P
BQhizrVb7lFkTebE1HU2DwVUo1eyYUOxwmjX4iNIsdJp63t+hBkyCjby+SnggVM1
Ds5oQlf/v+Tu7TCNCdQUTi7LZhnaXBoctiINP81fSVDzhdM4vU6v7eWdQWc60Rbv
yW8Cuhcv4K6Ar1M4B13kjV9yYjNMCwYfFh/nZYAx6HnZuT9rRdNORaxvBU7CowQC
JyV9iwnVQkiQ+nr63l/lPGR3jVCiY3jOU2mxDQBH5S0/VTxL8FlaTwoyddtaz2zf
5TAHfcbxEH/Y/IkfKrhntCeuTMoeTQblw0FZgI9FQ7s1pKtdHErcFGeVeO9zpLtc
uAQrubTahL6U20Ougwvqm/tSaR87IdJZPF3j1+YUZ2FB0+jfyeGLoKwRvm+E1hhZ
jNydyf60HiVc83hPEDBWYZi6cRTjfVcOWtds3eOem4kI0zUs/kv7ZjDiN6RmpLY9
Xq6by+teyadr21k+zCkWefKfv1/jF4Y+HSSrM2cUlFVLKwez8qgg+WU9/88bEMMu
Y6rmOwJusXWcHd1CfRDocz/TbUxKxChSFwCWsHSunVePUYGMpAC2Np5QcGlAqtED
3Usl6Y5tTdl0NwIcaaTD5d5AnhmSYChQfJ3xw+A/rVLSI3GyxKt2o/xwcBmBCkGL
4oYTZ1ZPXCMAfTX7of6enD/hFPFIUQseuLtZP0TLe0Pe71/NS9w+r4dpRo2JBeuy
T5YoClqgadbTNk/8XVrzT32Z7OQr6OrGYXCIJgby4pYteyWRPvr/BEGk6h4Trh42
iKcLUdj0ZiNRxFwk0wrv04XROQRq9m7/l9kUS34rn4ukIM/ibrpoCdsxCar3yYNl
yGKzHeLxOWNpBc2/VDRKtdCrqswmTFDicmjV7Wr+LgCLlAIRXRsPA4UOVfjIH7TK
O7o2yUlJ3AG3zIeqw/pmTpGJExsyLCd96OKBB0uwCDXUZjDCth+l7B74HTB2AIYp
WWB7jrYP8fDMbFrIVHZWT0MLclq8aWepvIw8O7hrlx6o0M/JxPf+yFe0w8S7OfXK
APJW4NPUq2z18a1s3xGG7x6uCMPM+ZG6HTPIGr5agh4wSWlKub/yRRIS5Y8A4irB
idO1X2p7Q4grahEUHQ6NPDL/HDyrQ9rb5TCyxIq0ahthA3lwT4zqpzjQFRfIwycf
I3KcFgoR0hxkOtnt8ZTcVz184mhO1QAfW/PaPgZCvTt+La9X+JMHIONfgR02Q5hB
K5BAyZzUxHWa0SShNKckAmMQIUkio4qzRqTOco8S78jSxg39hJTQvn2GYaqZSGh8
TuIcurkw/2HfXg5/Q52oNVibqWsqlzyYFjv4/Xh0hdHzajWwppIMMXhZTcc73n1w
inPjbo4S+J04RoVFddeMoJneezOF6xoGEDzs2VKmb4aAjAYepdA6Pfozy0wvjg6N
wJHSGz5V9Szq1pSQLtX71AsYk7BJMyQ24EjAGoLNIWHQROqwBbIUeb3U0uuO8dGJ
KMnn+lIji7PEhyCDg0QXjg9Mvo90q0dYvDV854KUyWKtlSxTWRIfBK+ugx4jeoMo
CFUjWzOC3al2N7AeYXVtdYW2VC5nPcfoO2MrnrNUyUdm1IEHdrbDO+o+adDa29Oi
pFeVhG8Wobo2FeKN2fmp92NIS738l1S0AzwC4PO8kJEvJptc/URLgv8US/HaAKqC
P45ot2fB9db4QLiRkrfkhQN7F7Tk/s6S8LWodphA42R8q2zRyvxP9GKOH5TBxnJy
CbI4tiL0rLZTk4vy9PHsgYwuKA6tW8TSOl+Qcufm7HfCoUwBjr8xjBMJ7CkTNKhD
UQyXSI2wMnLpVg3oIvHQTFd/BID454TSgSykev5ol9f8jzuJoD0LKKKYelxX5z49
RZknEpycItc6qTT1QhGNhPUIXcMpxDMHr/tSGr/UUuJEjqCtBK/vUxSlvuiZW8Ft
wEWvS0nIIhZAdtEy7PvOF5EU0PPJt5xuy9yeqanEgPEUHO0p9bxVkaMu2+sqTHl1
Wb8b0C715/FjAzHhCjhOSWQ9RM37sKdzcxXC0llabXDNJ9cp+FDGgG1C2cOdVuRE
sAjexRwm8Qf0jems9M0uOLl4s3EQH0F1aaPlwxmx2SLMJwt37QWuSyqmiGvnVXEo
JCDXqfQkJv8GsvbdxmYLCx0WhyayoOv7D7Z3K8vh0FVHxlhjDlH9qADJawtnWjN6
HM0fCx9aM9jv+FnPv5247Ug/aXjOyIAlWWEp18ZgOOmpxwFlt3gQVGn33H9olXVn
9FK4Qdz0hzTcFPXM0wLE/UZnVGySKN7rjx9YoVu8ffih+UZUVFfDCOqdKwloGRZD
Ds0ytB6QylDadEO82KCVy7KcbAjK9Hmgn+lrjqhUj+JB+mHU3AmLfrGSomeIsmVa
1i5qZg/Zl7sBpUeHoSmn26IVD1seqZBhzJoJ6F3Rekf1D27KF0b1Q5ME3oSlnHJg
wgLkK0FDcVkC3NepKfOpUqqQfIKbjchqV1MDoQBxSv7zKJ/sdwfYFJFNGkOPFIK2
nejprKTD3k5QdrrhvOAq0X22in2wN1tLBxgHFnxCjZpSRvfIeZy86+CYWgHji9Lt
HkLtsRXUsdgKhGJBi5bQ0qe8YBUOEig9l9qyRbmbl7+8xMlwA+DxqT92EvlOPp6P
WDmNc9UGs7hQ+J08kgprp2OorJYQEFhcXZwZ0hGXe0uqVX4As1jzz2etN5hkF1CV
lrIGDlhgrVX8oZ72673OQbrOCDix/ms/SGREQxXqs9RWPeYBW/2KQDmZ9rjiZicK
Q43Ax9E1UVFrfpcpTIz//isiim89QYhjCUR+RHEc2vslb275l7wvsSC5L+45oj0p
D5oh9RVE3MrzvkguT0/6mKVCwg8akBRIBLjGVEyyuy06wP1n3GGC/2vC1evx9Bkw
PBmHldbwsAliYhzgHimhCTPAeb4K+h3O7Zt5SeKoBbu2gBt68IEeVQvnfSOsKCqJ
IrvuuD5zdA40bhXWAjdm8oUWJ1xUa1S1aID2VPKKZ4M0lFFYJikXBGp0iR/HDma/
A2b3+MJRjZcZSxxp9JyjXRAqfbX2gA2+goGjg9xu4z/h2vzI9fEhNBdgJtImWsWj
v8QCgQoUsebpz8Aus5AM9GzOFTQWlSPxk/6j5rOzh3CJp+insPB69a7N3EAuGmXJ
M1/jSrFdZnGbsK4LCdjw4prS1zaunfwIKGRir80bBOab0KYicV6PTBb08A7Gg57h
Bs81XX8o0hNo9pcJ5GlwedVoFB4prvcziKIYYYmz1Aq2h54+4usXXtPm/FoNONp/
wfU+Iowp0+EEjhycPEOfINumELfBK+KngSwldijCziO8je1v3rNjbu6vAxT6c9LU
tHaw6WoMv9J6u5GzZWLk2fO6dzoyKfYD4lSFI0iVGLLS2bhvi5rdvg1FlTnbdBEn
tAcfJ/uFg2HszxubbXI662ziDMeLyN7+PHjQ0QkuMfzAi/sQrB/eBFV0oCBoZgOV
Py1OPd/6xKWjEi88mETQunYOJRk4WPH5FHSi+1HdcvXofbuX2sHo1iVmPEw2E6Si
ZbvW54h/OVr6tLU3PXBNxK0hLbumxF0dnTqPiL9D+vCNBfuxBFuvx5G9DkVAj+w5
iMqnKyZ02tWUdF8PxJwHdtAtpg2aQ+CnkWOE/xEcRHq8IWYUehwixlx/YKvWITp+
AUpJEkWCXZ2kgEfZEzOCOXF4xW1ugynJ8vkY5PRlrbzxXWlreDs6U70KAYpfhK6r
E/BEj4JKH83vlGlsZx9+zqFr3vFgpE5PPuLVy4O3Y/AMMpNz3gYp0EbimC01dpS8
tdPhoa1oYYsWktHJn77mRGnXMXQWDDUJ2L4gYcNgjLQEwNWxVKi0xGVvI+HP+ylR
SOCqjVT8AqCgSSbOVZFWJqkO1zYHtO4KInDw2x9cBy9bh9Va00B1w2YNK2hUEYIp
AUFDW5bRjjtMkcvboT039e2kboDrzYPQ1H+ogUh0sRjKTWanWP7voqOO/5HaW1pI
WUBv/3eNwPWKEDpvckdSWcXIi7GRxGUBwdnTLLQsZjEo+cbxskjaF4pwmo6aKTCF
JVzgO2J8YKQ8sSnlmDl6P6qXAOrIQ2kckQxOveFjgjBwGSQgsKeWy5BbwXANQ9gK
kUquStv0rGDE2mqINNhoQBkK2Hv3oJDvZzyvEwyGZc3Vd9YKbhDUXHQvgNSscCAb
L52u6wAX/xCbn5ouLnSrAc2I5VSEyn3QUpkOAzq/X9gqIoqyse247ns7vOpCzWvT
KtcL5x9NHafkFCnejikpp/s2sY8/5lNe9SCwdpRtxiCJ7WMlBNgpTE/PI/bDz0iJ
bpxiSCZKiKUWCbPo7C0/+Muz1dQ8pDFT0f4s2roC7fFF4If3H4XxsabMbx1vFH2Q
XurU7GRnrYPZebLRoBXhAC6Mcqz250bxqF43aieUnt6v75CPZI/88SDRA+wRktf9
KtHMwqjG3Uatqg8v2L7qHYuQsZMURZUTsxs+ESUFVLhlsxzHsgGglEtjVYEf3XRQ
4/sdMs3h/FBQlW/u7DzmJFvVPbRrn1iGG53D381F30hX0M/v6wU8NApW6f5wzAmD
aurulen7uvYE4MjXCollgZNUGKlUIMB45Qpwb9Xs7gYIDylsQ8vthegZ5+XEJZea
4IKYcMQMnNT/yEHVtJJjk64B4NaeMuTbEq5crTAjrs/rp7MMq05vXWSPcos++RWu
3mewYm2BePtHAIQe6EyPNVq3mUNDqGzgmYEI4+lbkSgv1FtNYn7VZIeCDFQoo5SF
5m+Zpu3ERm0k+M8Tn5EK9jg17fsefQ4cRvQWSRhqpmV3zPmNMGG2E+mZmfldgpEu
35zWaik07T0VeRmmY39POLSDJQ4uL77Ds/oPslb6zvbX7aedVUdfpFFHdE5VzyD5
xV81d37s9KPDGlARR/7tl/Yt+ysWWZIctPGtgcdskhORTkXSwSlrnS78eV1ldg+3
6lVGpOt3DwPygui3LNgBf/XYpylmhWivTkCH96hz8qWNHdzWoQ844Z+hpJD2Ssgo
GEkdgtzi3AXHW8P9NhvHskf5JwAvhMKN16/sypOEvSfr74qM5xGnR3c4sizs6iO6
ScLnZohZ9doGT2zDA4WKvZ4bTZtxGwvujJNhh295O4IynnQj86aPwLeTL8OrkQH5
zyopuZqJNI0WRZ4UxmNtvdYBg3YZ/CRcPPO6Q2/Y/DIhgV86xUga9n7jK6AtUugY
UkCjc8IZj/imBJSPR8oNQYufwVoCIXLWbgpaFG3uDPSQB4R+AuTVcnPwSzCzhQnE
s/4MC9JbLIyVw7MnU4Sg6fT183/9fVD5sIZyNoq/8wLFjB8PtC0nThLnWRfF/1e8
hD5wZv2YM8SJIkCuax+Eb45bLSWHN6Ufr2IN0EryC3TP/jKrdr0l95J+ZZIENlNq
6tn7sXqk3feZJcgAHuEnMzhBbJ4Pe+BRj1TI6E+rV6HKHAgjvz89MjdRnljtfIIX
dBamDs0SKMyNgZssFLoX/4ZJeaM+D6WRkUhm8qQAnnJAGWcUxcyHPq1krxnbownf
eot4i+PujcJDtVe9k4XplKXzKZgMJoTAL08hoUdl9XdddfWS6q6vlMburFzRA3kU
TwQjw/vv7do0iRT2cgjXxBsnph9mZL2CmWoQhh2XlU5FAVvE9/iVN596yj+2KaIC
6J86A4R0HGyOmOCf5YXgRWMe1UnzPAKRUWRt7+JYHFj7BTBQ12zLmm1Q4pV9HdtP
3ufK2VukOaOZru1cKL8Iwm7va8nJH0AWG4eXhh7COyHwVYnNAfX5331hL06fzUe7
SGPE4ogOuH8MUnvikt5FvPA2NpPolzTrdFvSsiuLfIZudfIn8XuuKli0QSZonxkA
choZ/Cy8zFdNMfDlV4k8Mf0EkUJ99ts0x5QkR5gVhHxYNN67IoLCe2085X9iTMww
CFxyLki5kAotacNiVAIXm5gKjMczzF4LnBiGFHaC5NEBE+xbmlYSRSwlL+7eYRZd
X76VVjdj69WaZybTzGbVKeHmiMKDp37sp96pLBHBdu4Ww0Vg/p25Og28dB7u3NGJ
g1HgFQXpSsbo+JZ/IIAEbvC25B8rBEB9bxuzbDcZQk2F+YzpldoR+w5JHAkFobAG
18E5euVQgvbARxP6ITEp0qisfLGG1ZqI+uW9mcK0n3Z3YruifKVLz9E0g55lvDng
OeHY5NqsuXMV4Prtq+/aEC5QVdh/bQeDFToC+/wx65Z0QkfBaaE0/wUVVvVEqyKt
uxbheWQSZoBHyPpoqLdV1V5BA7Vq9SIZxNtQ1YvKVA7pNJiR88StmfDqoC7AfNUw
6LPJQXm6s4jbAo4sZagabdhtliLaqheQ6ry291/H0+USiRMZb+zXCAdlRxBs/rdP
hVY/Tg88j4N2+knILEqoLf3wvWZjb9GwrJBZCq+f6JJnF4taRHl4HH5sAJoc0AYW
iGGPyv/rM7kDsy3uaw+9LjtQgsRa4ADXpaYO/0X8ERThCtiRm/w3g3k9e17gCmN1
oPQ59AkRM3vfNEiyAr3fGu/06stPpCekEhrt6fIoEcPY3zt4XfMtHKqJao2tqwjo
QwpYbXodRZwkYchxLNadofaIwUgxIaHiaO4LvpXrDZRlGCDhvXgUYiWt3W0193aK
Vasp6qtZ3r8kAA+TE1Ltuw1qFlyFR6rha8Y2lnQLlUxAdE0LZkepp+kKCmmyX2PC
neEaJG3ryNdOUVgAGExNgbKrRNr86/B0sGScbrBT+ZV0A8PTIdnSoNmixxVoRTdp
SQXE6ybYCtepmjp5zUsRCFJWV7C4TjJiXtRz85oXy3kGnQnw4jtqxJHAEtTctDnB
kdWvEaH0RevRowObdsBczuh+rop08Z9pZ0vhJjgYkJJ8epnIvK+9g4+eH1iAHm5y
pso6zNAxPvbOdsRVYQYGgw2OkHyooYa64GqllziMw2R45bLp9m7Qht1PRS99l67K
+ww5SmB05A6kwCspchlSY4Hqr1kCphfd3uSMRcp/nw2l7eYYyRRnJljaZeHtB/CB
U9G4rOfF3m0WP1WOvbUFsqRYw5Ngmd0Sz5hwJerLYuC2ucYsXJz38rXjyYS8jskG
0/ms7RjN6hwN5RzyLD37gk7gGI0GImKYhSkhyb7V7rcBhV/WZ44dl26fWZY2LlyJ
W2qREpy/1SFFvAgh1dYbUSHM+qwgHcEAIXn/B/hel6sHebPLbNEcVyQ5VICASj6K
VYFS4m5lPrperT/o+CyVzG5qBANC5VrM/l4jWvWLYecK7yYMPfY7F9g9dO5uoZSF
AMI7NhyBRvxXS51MhB5/fPJ9XJ/T1msnU/GJt4bj+cablYuUvzZnFJfZpkdkhHoH
Aq7Uvr6Qr2JG+hJ5OCsnVl8F/w9IyhkF+H9+NzpjLtywTZ5G2h7Yni9l9Mmxn6Vz
ocfwwgevypeKOnCdefNJudq8QY9MX0IbBPEPJ+F2bV2GCliZq21Gk7vy0et2Ujp6
bviT3HDVFtbPoDBQyb0NUvyaJkgH+BwwLDenr1Fafx9U4zzzXb/ngs1ThtxVTRlC
kwTxMFFFekanFDd3B+qzv5S3W86lTkW3qJfVEqpsUHgEKo7FQPx4YtUbIhnEe89s
9Vkm9wz9k/eOwHVQaX+ZHZL/eCstH1GI0ZLiX7sFUoSfKMmOAQjYtpcjDOy818zc
SRHwCznXd1ljFk+znVeDKN9y0OtzR3EPU5/0mE5LRCp+7zNHE43/1IV7qkUQClm7
nm3c07xLNCAtC/HfBz78G/f7XS071m3N5v8ae9gv5Bf8u2iYPTTj/4USNAzmkoG1
2Bc6q8oG95SpQVnXjlwGT77+3j/hZSE0Sqbb9Lpsh1ru4xclItKkQn/0xp2R7B4J
3bfZnFa8N0axqtPu0Le5aPRf8zbVuOb1PYUbV8HzrVBthxGJYpcA+VZIvJNcETd/
lGrzNMSXN1bG6AqdU8dHiqXA3fvbfszk22JjtvvIBNOpQVan7Em++eClpzR3U+9L
/JGvsbqY24bywsU3gSU9OYzz5+WgG/ZJxp0js9TweKSn/NUf2pLFunj234/n8hI1
b6WwyTrzyhK9aIUP7ewJ3VDzie3GvzPCVjIf5beNYyu1Fhang1enVwdBlshX6Dki
wp1e//kc5hTacZDfHCxs5XESTxl//Y59kOpXj3lYI5yAPCTdUD9k2WP8jujWSmA1
e2UNAhHNWTt2lVb5JX0BN2IbThBVUu0V/Ud/W01qaG4DLY+FKpMOU/u0pCxrcIcN
Wt0qAclHJJYUWfCqlgdEBZfJEuawV7Z6sCeANzCwhaO1rLtmb7vOv4UnDVfxS5H4
WskAHHroLH13VjVcJWGUZzZN4X8LZx5qxxqI2uCCDE/UvaadXk5IUAQhsaclDnWy
9LQ7+JMX4PXFI8tmtAQXys4MqpJEtd5awknK0naqtjso12sjP2mo+sClU5I8kDaz
xJBnyUIebLKulvTV9HeDmotFwaVtY/+cr0pnVgRbhAz9pU+TmI5Nj21kMQm9qUGU
wc/dCClaXAy4MIc/mUWuG5ZvLyishVeoQiCNfuwRe7DyyvYyI5oOMKwLawpY/Tr5
b+gLGDMBq1exlleQVetDoOh/1RxVHFJKxoZO4u5SOoWYBbz+Y1/Ux3iHtj6wflMR
aW3V9usY2trCLX2z/NodmV6erI904ehuoQY+8teSUlvW0yXinvknf6t8FwwVHy+T
ZLBG3eHASqcFI+YcRpmqJ9cSwb/ssx1wVN+BYaGkoatbznrV18RduDgtwQkM4+BW
iWeCChOn0hAJZPM/fX5tuhIhZmm+H2ZdzqDjN3iOOpKgtAf41dllnVCFcAxZNzG3
Ifa+HASeuuDo0T/IcQfGNKR9xEL9kgTNPmVK06Uv7okmuswMSxkhrtOMqfeYNJpB
8Zd+NUnDPTrbCmCt0acwKsjWqCrJpBtSNthXT9ryBCHujPq8iujyHincOXnmWWy0
oD7D+X+jwxFe8AkJfSnYEYJaf0H9/MKP6y+O5CSkvHZbfmcQLCVLzRfkeuEWldVO
ym5hf/9VgdxN34OlzXBgRH3n6BSz7iunrHKYwKHei6mD4FxCHy2YXWuOcdv63Rbs
cc4Qr4afyE3XYHWrfwoZG3pDti7b960Qg0jaqls9jqmFTBIgFlWwpOdhS2m85nTQ
oBKl451By2XacoxhcGMIYd/fZgr9T6fsf9qDL631ZlweirJzz+akMaqzNn52l8B6
tQmpzIF/5RQ7nM28IQl8oz9/8f1M2gNHYEqF+s39B5LahsnoICSGYYeY7GnY5zwD
4nT1eLvkuKe9WZrkDA2Otyu5mEYA2dTnlKBXkZJ8IW5Pg8MGwmwwEWpP4p5xgF1w
5qjUTWc8F58R4hx17mjxDIVS/3OCYUuzCZiv/a6yXh2YEHrV1hnOHks5xYabjL4h
e8y/li21PkmzzahMWhRtlArRVOJLXqwV+SKtM2YGHpulFNGovo30o+ILIpg3rHg3
HzvLg9bbvq85VLpSvJbtY3rwquf8Ud8eHNX5bIBamAWoOVqnAO0EDuRIodLm+NUD
QLQUeVyS/3FrIG+o/HrmgwodDuRKnQ1YipA1nqS82AGVmx0boOC82adxqntTd852
rL8LZbGoAEK2VUJ44/Et+K6kRH+KpFUn7S1b+GXSjnVMteufq5mebIpZ5NtiGiVY
Wcfc7ZJQWUQl3I2QdYAqL5bm1SKEaMLBWV9loiU/68vZ8t9EVbe7aFXSAXgEe3wT
UZU+SNEL608D/gufNYepCY0l2gBoUarmZQeQ5EjoDnRiUWHebMBUWF0QjBszDJHi
KutvUC6IqZWTpUbFhMiMdV/9FCQ7KMDWmRfP+0yyaewXQnssFh/dPhJmobV9nqKA
n+lbsm2icKJ5EYeNHlEwCLFcc3HM0/9YwAwAfIdTemD0tOe96LvN4EZvXMwRyFC9
Jh03g+uSgbGMpOanuDmpM5uWhZsfb7hZFEF9bdbI98QfHap4nac29zZd+tS4t6Ew
Qw/GWdiJfSCMva4VaJzdh1qIjCfMBjHHpOSqz3N/TrviiXokSMN67jDt/mOLku3y
cHX9t7nEW9KC/ia2SpKNCUMYxgMv2K3+1UHEnff5H36pFZbStVr0B1KW0B1sGcoi
6T0mXh4QLg6oiJaU6DPPQSiKbHmreNXtMOlnh8VR2Z5hHEXP8fmc0ljgoYSiy+oS
Xj75R69/4FlJzT8aIEBvh7rf7bkI3MRPmZfMb70D4H/HsgRUzuW3kU2+HHy6FERc
UkQu6cbKO20dMAugc5pQjhg0rsgT2mwGxMa/WhjT5svUox72Z1d/BKBDtm3JRwDo
nFUy/+s7IATCtkXFA+t8192T59UavnM1P03rmhLeCrgqYUIHM/Y0uuAoMz4XqdRH
oCiEjtZm0fWzEhRe+JJYr9lGyVeyPu+k3q23Uv4wqHZ6N5oACHJ0jze2m54R7FaG
1R4xTb4mAj0TRnjdg2j6tyy2gM+9h5r6m3QKS0rdGDb1ZV5U7iDYVNQX1OjaFlbf
jJ1gjL3h/tVPDp4TEzI2gO6cs/xLjXE8fP9APGBeCtzlXWsgqtVXpB5clwthVOn0
Livmm2r1fBIIEfOUcaDh7C0Nd+2k3IZ7LB/6VkZOR78gTsyD6wy8O89O81YNqLA6
IwyKFCHsnjvA5rw7kTdXYddGpiXjYWuXUlsH/AdsMsiK+QnXwypNKGO+tbJ+nDNy
QQZ3d9Njw1xb/68ZCT1uvjhepnvgAdQEGzH2irFGDxPm54bTxn4kv8lxk14auWIE
nQTL9M0VsIFzSHyo89fuSMihiEhM9EEaR2Y0KDBMrOfQnYnTQAAVT8rvHIpk4F1z
fqt/j0TBsauhh7FJUYqGwAsqCD1KJFx2B9p/oUjS2Z6SEt07P2up+ToSAkteHW7/
6iMI3ZdOngjc3kMwrvJjnh0n5xzLp6DMQmqo5RCSZz3fQXjl5HA42hsVqMn4BwES
kQeAQFe4eBYuChOE+3pIoXvYa4tlgSB36HbYAtdw7Xx9pfE/bHVltyaxfaR2QD6Y
KV4mFmKTLAfUOdbPOcTywvz4p4bPtYU79m5plpQai3NsGxqnzikwviyeZkn6CmXd
lo/o3K0jIM+2Ty6OwG4MNWjhfC37hG07c7ZuV3AO2WceNEHdC1OYgwPEfgZfoE+f
W+3IHLE1XgdfDStqVCuwjgt34BT4AvbT+1Ft+EfJEvYoBW9rAwPVyJxO+hMB5jJI
KkPn2bWDsWtu6Z9UzDT4YZFvpsaojBbp0+klaKERIEkJnJdn8ONV82ZSxibNey74
jSAjEYIY6xjKtT9o/Vy6YGhBKpzCMATer+Cqjobg96G+uLhUG1jhTJqndux+QIcK
iGveYk22fwTZckgHHxQu+eAvgIVckx30+hO3ChH+cVhQgSH3o9E+wM8D6Bzv0voL
zLxku5zA5Wg/w+oamEc5PYUX6sZ3dCGUi1ImlP59tuJ3Z882ZpIli5sr/n28TX+r
k152X2cZVzCO+ZklYo95/b4xy4UyQuKDGNDbCUJHQ1aGURaTXqzBJG2sEDHwuPoe
FOFRtkb380ewJlQ0EzI6XHGt4T+pPa1v6Xv2RmO805qlhw4EpPOh0C76r4NhOZuD
YTadjT/AsK/9LXEC25DVPViaP8JWy/dbbvRPNWsxh8zMhv9OSs127s+RE6Cxod4c
dID6k9a5JDOBG0wi5wc/6LmyvQ854hKQHOcojkW3789GE9DuOGSJo/qF+dUIdlEs
TpNy2Vy6zYvDWOyoG6nsyklpl3D6wYRxAYPVUMqFL3EJDJKzCpYCdGRfrIFZ4bQx
Jj2X6BS5dZwCcRH3egRDtBfaZOtmJ3S3y4f3bX8o+mFbUBN5aj5Y/qTuClyXzCVE
VY+v+lho3YT+7YIbG/lWrALEgvJvIUGd8gsn0R+YVc/X8ZFoVFWumdsB8hR5eITq
iIx2hUM6mM6lz/gYA4MGpRscwwh/VXnDLf4O3I69tt4eONuZ/nsS5zhIkALKYP6C
3EgCjnPTENCWUEahNPMFOtdGQ+0okykxLN91NIwbghgOQx0AoaGzVajuqJfUepqx
AsefE3abyew5FLDpnZT6yx//e7Ioydt7ml9J6L2/WVIbP07jZMtDOMNG9uhS61Yt
4bATAtKibU8QVKNVSktiiJDQKQMe9J3rn/JQY8AD4TLt+44bHhpLHayQRuJg4MXl
+t9OQeCS7zRkgmFiI/XuyCTBvSKroZHmwXha7PNGXOhKlhiB80lk1V3mldEmlUe7
Zyrqtzks846CUgvM5xszGqv+7zoeMR447NbZ4EK/lPpwqtlVCuIvGGehK1AmTYSy
C1QXyIKlZDRAvaAEfF2hqA5jII0moLicIvhdAzYGLmDGAi8rdRZP11R5/npu7tPE
3nijx35dmQT11CmGdh+92ASF+PjOWr7pxhMrpfaQ1MbpNLcwH3hxn00coHeaHqEV
DEVWZzYt2RZGw11B32eqfeSMA8rtDqwhFmB9t5rcYV4cubFAIu5sYGCvaBdxcRk9
qn4j3mr5sMAf3pzUhFN2xo8+tEcdbaKaDlfmxEHz5T8EboZ++thR71PmGPVuLbf9
06rPFD+pTlG6NHh442YpOa4xLb7yG9tkbFNAWJ8stWcFbHayMLOzP5aZLJ3PPvqS
y/2Y7UTEfWcTvt50aSpv51k4Y3XjO9Q2kJyHd2A+QIv3DZsIjvrt3REBKFPeddtT
bcy1d/Nr8IYDJgUeOUKOIupcai5RH5VeGdtGwdkphi7g8Zgz0yVXq4yAGNf3Qmtz
zsoP44/iNaw2LDwtgCkoC7rFqMO6QHD6kDNb52QnznXXA8zdni+injcoZLj9NTuS
SgVMG042o13Y0WXfjGfZsn6G1QzkydDpXWI6Lxe1XSS3dOCHc4zyKlDhnZHyV8KV
4qUkN5HPf8FGtTfZyR3u5l5LsEpSt/JzYx3HooUjHtAfvWHF/LAc/FDx3eyP8O5/
EwGow68q2XmPfO/H4nOV5cOrC/ghZbGvVMSi3mGl4bafVuEg/trUBjPtgWryPpJT
dfvXbieXrfJMEVaHkjlUkrqcg/1HFqY4ZW2uIuajTRAw3BvyCVUNu5aqLCXGGd1G
C4jx7Qf90Bit3COKAyQlQfC2Mxy6+FJcsox29hPJipt4eRhXmK0r680JBeG3W6kE
4kWvXC1Jr8v5EYxYH/N7Ny0p3tkgGNd8jAeTD73EniRvcDtENW4g0TjIg6zUfFxr
nvWHejZTtRragTcBW6vdFgb921Btf0u9UNGNsoJRnp0QLy6L0Bns9xzzoo21l7ZQ
0/xKoWpuUiluPtHufZncVGBNNZeG5eNGd7zmyOvnWBU8ur/peUMihWjgrkbFdAnL
+xlvACTlyMotQnX9dDf/4+eoUPyIypx2/Dsqg18wTmhrzNt7jMBWKJXLUCKR4sYE
eciYPH8ZUmNzZOCczM3fRzIUhvWb29glHP9drBN9FQKzuMRNeqZt+0WClTtGlInn
a5Zqu3RdDWoiC14/X4QCNprTv9zt3Na5JnfgBObicmfv0OCr+D/e1sqndIeCtnDy
NhRi1U1zzay9KHesog9ELlSff4Wz2FsUIrba29str4xqOvyh/P/namjatG3eL5kz
enmFHtQBWeE221BW4rVUNko1cVCOE1dfw9hAYlHqJBzXWMNODK4ophWn8AwX8uHJ
m26c3XM7s+5rcBuxb7p5ZlqyRScO/lG2BmMSLi6W2rpyRO4KYxdvrOlWyp+hixPb
Ppx7Z2FYzXwuASeXHWUCV2utlbyUNEjZnaMPbbIzOHVF5qln5a5+DiHR0Isltgjk
tg5QBzFxS95IOtVrcmUZEAsl8VK7HtYrU2JYzK4rD0U/D+6yk2yzpUfVZEY1GqXe
006QdoRlvAD4gtN/owQSvFdi0Vg+fJ8MdnyFAXFhOBHX4TU7yXpNsOla5OhbflF5
3uZfTTOjrBaEKdK0+tNvezMsWJBiEFPevd9mkRdx2eAUV1sxfUTDra093A6pXcXa
ZiAqVzhKzGma+uavgyJUuredeJhB/Qs5H5CuwaCZ9HzOj9Iqh7WZSPBVUd+PP6kV
P3gpW3dQYUi5ws/ZqF89C7+P0vO9AkPEbKW7/bvj6PrNqctAr7o+cry2W2JdpH3u
kFzePhjKR7tQkQr7Zrm8MSjoIjndc324z2YoKWg/wwBU5K2qbAQV96JHTjhDefvW
KdMdyr9GfzSfqq5RPD4LbWw3J0M4VYHzr61yvjQzz8W4BYStOYPbL3zl5f3Dq3Hv
rS2EDhlClEFr40ggvf5hRbDaZv58Ol9qL4n8PStrFrSB/VrmBG1iO+a9l5Ke4UKB
qFB6T183gLQA6Ic+KSiioghUvhXwRAPs2q3462hS+Cs2tUnpr85d50cyhgTROoVC
op0omk/r2oViKtYo6bCgL7HsZr+KhuIeI8dHh93vSNdpIDlP7Pv8piY56Kah4OJg
Qfcl+DLohfCsN/3lliyFWS8VUa2lqW9lWnEzzWbfRr1oW0NLQgO7JhEqsMNvOAvk
u4EvBt9qxD5NcundxQThHp7Y4tsZqpvwI+dkDQj93XkMEO8mIG4+F6So3PlAjpMJ
Qbicxo4+gRsNZTH3Z/lK4NJLC7N5srZgEa5KFAIkYMa2R6l0Sw18qc9bDqXa6b8p
VVCQQchRKvKxaxk2StrBpfn4Z/FR2Zdo0ulFfR6XnGNxfmSSR4po7at3lIIihdy/
HLqftAEOBtQL8sar4MRtFEFqr5fEfY822jCA85CaqJOL7wKVBxPsRf5VYP9eOQNu
XMUIQie0Vdg4OPXHYgJXz0a2yqBXAObLOEkYAPVmCXEQFywZ4+z/udv8OwnWGY4x
egVY3Az2CC4M6Y408mkl+HDqCPIV9h66ZM0ogaBZW66E++7T0kQFnD0TQTvhDck4
LTqTxTPfRdwtQCMIXv8tK8SRXQFoEng8212pYDotZOsufGDQVu9x0fFITO540KS8
WbL3R9vtpWwNCi7tNBrbsQXEaMzeAUFmkvc9z9+K8FffGThsjnn6eOU/Qz07qLcI
yOkeZy8QqvMS3EU7w+uOTy81rzXG6SHDf2+ZHFHQh5eT+Jfd26OUIva/IhWqWuHZ
a5OcSQQQAZZjO20SRGfiwJElaoNCgmlIfFxe0lhElez6fsikeaPd7r7o3Br2acMc
35wdn3p99hNGDnPmi9L80K57vW+RLqHjYibylhZijEGjdONtY9OYfrgZupy6kZaO
tI5PubCe9darSvaM93frKxpyhJqEF40jdGTq4j0kxi1k/Ju2gR5iZWqLKvuqw8P9
x73CvNdkZGrMnbaQg00uWW4aH78KsAjWlsgbkYfC23HraLb3Xad+7i2rZJfgPWYX
eRl/6iFKoKAasEjybNmfEu5lqqKLy5ZGp5QIJE8siOMdb14K42Mz+HUg8hGezZwX
Nrz/e3IkY3lxzJYyIK1qhVN8Cg0GdZtQSBMHDYzRrjWPMXbUNtHtkdvJyhWG+B6q
pMO+8mQtC8IVL+z1OXqmU5najty6dCPNjITFSouo09j4iBSVnT8vFb2vdH8x61uB
JNtT8kj28ZDreVEKCW93jGA3d0MVcFbfGbZ6Gc11ULZyFNaseHMREwG/MHZFgLG4
9FBs4fl4FpliMyMJpYRdmUC9/bywROURtNoeIPYA2nH/kZUnIpVC5RD2GIw74T/P
1/0WNekicGUhjd4mR1G6lypncWG0OOYp7U/WdjT91LMnhnyGKVuRgzi7erWVYPOA
v/Ojny2tq++LgB/BClr/LTNgvevL3fW+9ScvM6BqwDvD1swrOVTTMgzutKtxEc4X
1BkheBls+dzWsCZPClrrcLpVF8NhOHH57SydNWCxavp6SfN6495gUqKFkD9eWHAp
mqTmWJu5ED2B4YXMVFiURT+VvSXqcCjisAYKIWWIDx2rYnnwOWmi4uF9rq3ecI1t
NS18+cwNNAG2ltmdzAoCjTF91ODhJiQz145ubZJLZnr9vz9IEO/WBkxD7Q/00b6U
ePxp03YYcTu3dYK1HJFHteCSxMEiAJ2IJgqr2QrX/02tIgsflkehwgCikOaavb21
rZ0Ki6O57hPgHbf+as/n01V3xID4f5xeyw+mewMyF/r/wBD+X0ZDTI7rsJBTcGdi
70R1ZSXfO4tL9oS08FeL/oNpJfYZuws/+CwWlaofrFDzARlP6T3yeYkr8TmbABvE
qZ9jWEov8QVVyueY55t/QVkmbU/Q3cfIXC1duTlbCcQ22ICJ0500NRSQKt7j/krl
qHUHOvjnwD4IdKFaiV6eFR4Icc1IpRf/DPEvVJ7SPMLZvXD9YOHpqgpp9yLjjwKG
TLWaViyq6oKEyW78YJZEXWo88tKqdLV9Q93z6nRoL4K5yl/qlnTZXOSNkzPkrgHZ
kyPdt72rIUJDDWTXLEinlyNHVWajHxhcKqoWPQoCWtBKShkV9tDqrrjwBwCwzjE3
AjQNshROGozpfoJiyd5J5XTwjmNBVcw9yfq3BzrJi39jVwBg75Ul3/KNXHO6VNTE
uwAcUyrcUCy433LUpPSl4RpgtDc52ejS1bmYQSMcMrFQazvVi+9I/gLM4LbFBvQH
Doq3qIJ8Enx3HIjsNvvgXVCfhloVGxQGcge81385tqnxqLsvAW68gvAvKpDjrPl7
Vdhghwo+oqHA4sPT5BvZ7RJifodtZkYXWft0NNWPA2cnYm+0x/6S9nnTccweQ0D6
hwLlpV7zf12TtfO16YNkeKYYjDC5T2mwBK9zIVrgleoF0+3qjaXzvKgCLl65r91Y
tvn2+A4Ez2W05Fu07NFpvydSXCpXwwLSzk9e4k5gSgVB8EjLg4nDX66kgRhB00Mc
Z/wSi0pLzsnVKs8CVApnYWr3RKazGoSnx8TOZ0g/batvFbin9OoB5cuTv8cZtxX/
thCsO9prAgwh2RW1OaJB2qYzrPlBsjyZEDQdqCdU4Jz+W+eK8a4/+G3MddoRrf0k
PFL5Qfe4xz9gkcN9z106Sy0yogmk2VEj/T9N4r15tv9B0KsIV37tSYuxRPAhhAIf
cgLG68NmUPNrfZ81iBnO0Sipsh49GeMviGzNR8z8pmcsVCHJM4ZKXZEl7aUlKke2
feTxBMGH8OleIPwRUfYHrmU6vjAqeCQcFY5weXmTsMgdwbVm4q9xvvz/ZaipXtgt
lW9FlAuHmSqBknX4Z0kjJHHL+VwFudTv3DIqxsW7oyyboJsvDAOcerqUb2cSPDMR
mAlG2W7OfFfBMjjafHX92CVLt4HihfAZ6gEuQd9iyWeNQY5rO4fDtgikC1w+TmWe
8fwLFwW+tvxKgNc9to72ERRF3in3MFQjwt1RWptnp5YKCjbZCH5oJ7peTInSC3wn
mf7qA4N0Ynopq8TbOiK1gQ9PAwvStVBAdfFHHA0rna5u2o6bd8HJwi6weBMMqBTo
aWd+D2c5wb5o6yXS2HYfd4lCoVpAMN7XYh3Y5my85c0n7IuQgyEoCh0SIjmTJkFI
3qHcS2xoEbYpowsVFqQTfdqC2a1Oz08StR7Aw7K0MZmZQ4pFGyuB5vj5QTigYUEI
98Qasi3xayibZ1eUwu8N4uk6sdiZtOggV8Mg3BGpsFePNq8B1Z1T06mfB2SczBxY
42Da8xRJJFszw/7n8byrdM0XvJE3XA23J3T1LCBFf3VcnDIccjzHwmKtfNiu08zN
N3lRkqzW04kXoZlmC6TrYJEa/AbaxoIvkDA7WMAv4JlN/HSkLdMFU1F3HxgjKNuu
ZPhWt0LnR9MpI5KP5dhfPKgnu9ElCOPGWlWQ/6XX8M7g3JBZdnC5HVrjHi8OeKhR
jXIf8FNVmuPlAJu0y4/0cE4GUsO1cmk5IUekUJwRzPvO1is4LsZS9RLPqlG1VyyQ
wDrpjDD68O0m5VglHV6iW5dfMDWRWeq0n0BCMQlYO0/vExEEeWTC/YKfWkcntkqn
OCKAjSMzW82xoJG9jTTAiaPBIu0XHMhculu/ZwcOYVX3ICjJXQKUxITqId0z8ZSa
2Ys5GIRQjctdvi2TU7xkqBIdgQhueETnjAvGROtJVwzgFvuKpNB5shnZFdhtC95B
qGwlQ/GoH6sjcDkTVwxewsUHZ3kx2hRb6L973QmFl11DRr8Se96tGe1/XeYVIXkT
RP6E6EivduYVri7DvwjD23PeRHMN/Pzq0pid8IVkgoO1QiZ0vTYKWe8thV1e/AGb
j1zFmENhu2FsnN/akTbfRWIHp+MjWDR+d4VZm0SU7cRT0+QI/t18+3yPEGKNlxN3
I00HkdQlt6N5zqS9HD8BOvXYA0CEqbMPmtzP1AmlF4kxSaCDO2wmMUfZs8G8Lo2b
HZfitY+nvmDlRGePYM0ckIVLVB7ngJV8DcXPt4o+10+1XMUWrRQ7CaDupbEkZmoE
x7ryjSScpPdA4bRWmaK4qK/pVwGVRtxt62AjX9dUC9H2lr6qdaT36g1S+ltMJYw0
MhdB3KwCMl9BBLmJ0JxjufQm8tJnmXMHjSOSfyx+cEJd9bpndUTMmdDgMgOkSIr8
R+udDm9DJChiUGogcqW7tmq0ZN96eocl3e3BQ6LM4rqVWVANGZ06eBkb6MkRA/uK
CrohDudHfwpZEGDRfsNIijmSfrZqIc9XiHO5heramtiJ8J0HQTJyQBf9U4NT0Mge
Uo1Y00TIVVXdk7d4QP6bZmw8JuMwBj0Zhxh45pgUF3Ez6U4idjLYBzhNh3kHZB0a
Vik5/lGQHhyqjFINfBCyKGdjI1r+1pt7KjSvY5//o6ixhYhmKS9q8kDlXq/HqpUG
DemUf2sJOH0EKtzT0QpeCg82FZEF33G+HfT0V6xRoU5f9f8VHMFeH52bW+0S0jbj
CAUJTV9qETI1iPDbbE+5iVvywOI/ZCTVmOjJ0i0fSlo1+KUgl+w3WicBQEafYtW8
3gmKRfsz2YG6I/1VwO3PaUTXBJ6GBQX9wcGfEyReu5rlEuaDwo9x6vvqHxXr+5Gt
BBagx03wHwfRlyjk5XJjD0VeBV5VjYmyLTOqSwozhCH5/OjggPYg+r3xbn1c9ci7
dxsUTXhImBW2lNrEvCyKWUYQ3oCSvx1/IbjhOZ/IbTn1K16FMXI82dXulHQh+xtf
L6zDWYKKNDn0RfoR83F6VISLooFP6hmvfOXVZHUKeLy3UYx4ecKctQvV+6O19xoA
x2+2dpt5LC1tQJMDQZkwzjoACxj6yIdniDgxsxCv6DJbbEmshuwHPWF5LeKNe8zh
UhYPEsMq80v8umlvyLB7fuCaQ99BcUzVueRNAzaH3NUSve8OWQx8+HE9DzCyA9c1
2usVNxcP0hvql6yIfINSf29NDY7qM49b3C9QCoVhnXWPIq0od6rXYIWFCHjRTNlo
GSE2RgielBcoyxnCy91jihNSESzeV0tCiNUgbDpMBQ1yUamTraBZoFxPb4fs42IX
CeNvIazDJXgNZcMjIFRg8kxvU822fQjTmQIf4nRufqvlZmOKX7Kou+e9T0/mTyHb
BYEKPe+RYEqSqotnW/MMI+hMNF2hwT2N59oG3q3mX1+U8E7KTnEte98JQApyPB/J
ZaMAgBBOL11vFq2+sgghXG4VpdfBQzalsID69uP30lh6IdnJf73aoMe3JEgVPdJ5
FVRg/WPFn5eGy4BNG4At8osL45rXck13qWoVytsNUYcGpriQ3Cl5DurjtwF6G90K
nuLhEXdPT12RNZ7HmSZ6P+SBFcLPRV+P+adrynGZ3Pj2NYAQHivYEiXk5LdiQdrj
7Kdsl5CP46y8QBAV3SvTyyBFtE2lU3SBtp5Igu/4YL8ShT8BFoi6AOBgKFzOaPyz
eLA1mQbUb8uM5whga1+9uBqnHV3RY2qTh8X8FYyoR8/l+MEoZ0b/SCs63MWMnr77
fEvenxefn5z038exYVka10pAPMVvjoVnHG6fzzAkp8MQ7qcmHG709K2YT+LN4BvQ
9qwVjEs56s6ZJIn+c3JfKGlNHiqdtHeeXFQax0izcrt2alDV6j5fvv2LZ2+2zsfj
LFKJfWF/QNfTwzmYh7p0nX4EMiYqSzaWg1XmrVEh1DC8h4EewT0Mi1gJCLF3UnIO
zKcblSBT6/YlKvvjt/ldtIU8wnabezhp8aY+mKRYJiin5kJwf0VhoK8XIUpD2HF9
jooQEiIf/yw1aYWKUEsTk8pKY7Rq0eCVMARLnrwwpQlHObDBZhhEY6cTLb47U8Hr
tncUweuDkCQ4QRluR0AaGyLgT4Gf6OF6CHeZK3IWXICaAR7tgbTagCtJltILM7g3
THvqRYCvhO/GhlgCHOFcbA4xoKFLBWNueHpPNFWEMNatJneSCXrW7Fmp1Y/ZicvR
mzphF2Ww2rTzEdgwNvcXhj8t89qw3iBo6CCObiEsBA1EzEC+PCOK5STiiTKLKwkF
XCO4HcEF/cdU/a4NG3H8l6XZjWeQVlSEcUT0TMsnJ/r357OsEbyVtm7KeLcRONRF
smWZq6zUy3CKwgo8daFH/E7cqiAGHAYiqkQXJutLU0UiESIKAzMIKIGJX5Ei+Du5
cP5DvMZ/Ci4mLhoy0LJY4oT3BWgemaZfm+ka6Ue77XLVD+oQSdK3XwZ5ad8/ExVa
72yEoEZn7vKW43LImchzit14cei5GM2a1Rpax3VkLoCvuQYBKXOjJqX3wmXlMe/F
HcQ4Yx8NsM+KTW61pY0hhKUbBXqD6RsRjco8K3m62QXoR0jDNdzwAYjnSTijX4AQ
MaAeb3WNyf5QyySkv9vwfBlUsumz5Wbmtyqa1UvEOGPInz7p2JMo/qMN7Un44uTH
Dbhum2IfNlZn7kh+nCO6W2n04tZ7GhITXdREAVYqVqgDFcHivoGgCHKQIAS3ufHJ
R1qDDJVUFkdCjL0QfvPB4HnCL92W5wzJe/9ncKSt/iKTJ2uM6ramb2VVCPteisbx
wrMPht9Y16Zq4A47ysChhYGIt1YwU3mjN/uWmqbEN4thPs9JFTTvB7BrQTfYR2VW
z+2ewYrxadm1pZ0YEKgPA+BSdHVh26fMZY4QMu/mmiG0PrxZi7d+ht7lknjcIuMd
7mjZTwTLLmU2bK5w5BOTqej5OEPN0+A6JKYFlCe4Yh7vZ2udP5VxLTE0cMkdplOj
Sv5GBekFVVoNmyhIku0sNaEemRSStJ71XV0VILh/P2FAKYnd1tB3uRtVVebDcOT8
vT0cE0DgGDLqBeVpMSVjIu7XhJnzpXpWyW5Bx+ZA8Qa4N6j+DHt7WIvFhNiERP76
YjMh2qAQz2eNuZhaksVFz6cJOk2iok6oUT2JG7Aw10jaWr0bFMwPRBrWhIv5wsPm
UALVCFtWeTqNRVp6dLPL7gsJJ0yvM5eRMZ2+/ZS6zQQ/uxkaGIBDNqqGEbVBkmy6
83CuQ99o9n8275ItyYuYCpitRWI8nH+A/7Wzy+SyiwPW0TBrjbQQZuKf5GUUsHg/
94TgC4g9s7Pttgcp7iXK7YT7kaUXC0K9yVgkpc2oiX4i6qYenPTwEIMwZ8EuTdZg
0ntUA3IcgbSi208QLUL7Lvl5ZDlH/tRF8Gxdavp3C7l+cT6Ox6ytdgUn4sYNdQGC
l9nATElmU1yNZDePoacISwmjK/GkAj8UlFQXW6NI+9MmrQEEOyIk/HBos79I4TWa
OnXHrDhedB6UQM5xpzj7jxuMTShjOcKRy/hhh6Ih1kR20Vb2vw7d01gsJZQRRoLw
NChMMu2biZdugMWW2bLP1BXVdKWDaSOMgnRW576mGaoueTieqUxCF/y2ydxviIMs
e1j0z+NnUAOMwIj4JKERahpVUzibLpmp4HosNSbEozPPsHVVNlZ90yGaGaujy2Ph
ux1rh1aaV2MegjvYqsxx9xUZx8OPd9VSGE3owexUTt/QOa0rZatfoDmcOkOJzHgr
VRI4dyVSuw2DpyaPvOBlYuy2lW4dYvVBoUHLEMLYg0Z37p6Tl7lyV9quj/LHHt5w
UKsuHnE3EyaYInGnhtl7Ofon3mc4KKsJW31GEZdXUpcAScVoEAwYrZyv7oDM9v5u
5b/JAuBGDme0445T1fFT/P1R9+NpxM1KtaORQrgCtl5vQqcgCyyW6c0hAA9Tzr6r
n+63/0bK7Xpz+SORDF8mdS/eqNal7yybqevSkqSN56CcCe5261qgMNIUoehjpW46
j9j8B7F71vXxHqrvqHJi31vBCs0rYA5c1MjnZbn4nsGN5KGTBvvXSpz0Zwjm7qoG
7wCx7JaS93IU64sT3hvSQrxHhOLUtUMxN5M+4icvZKD5idsORge9hCWQPIMteglb
4cADIi5gCV3wXaEgxtN+RwThxxp1gb0zgvn48o7TL+sbfYu++VhdfEB+KCedzxWS
bo6mEtJnyUM3ptrx+8enXMYvI3PbpX0K1MZ7u7lwlBbGWRFND4niW9blbJGoIk3x
BHGqw/feSFOz+BpOVe1mjWLzGwSiw4VkETe2aZluuz/cJrqfU7tH4uQPJi/a8qGy
wKv2So1Qllq+900YfN2rP5ZIxdtxgcRdiObz2OI7VnMHlWEOCNozrD6j+BEXA0uN
Q6t3LSYaBGw+JsNQ5cfEEuF9boiIiGZCnjuoEUGJLYivgvrpluNPFnMgCweuWcJF
L9S+0rwQqKsPu1tkO7u82nVnAHC2d+nEhv5d1zjJiBrFs6EFrW+VYWZTjk6v2hRF
/ax3e7NKkhd4Qyx1wkJFN7GU9/cu4D/6qpAjUSgXapkUU+f6k9k7+zqmDUN5iwFf
3shoyapUfRaVikO6Mb5XSVAnzyzacOgiz7uksSiv08SNR3df+ZZ0iJSPv6gGygbd
sPcttkGXM6bpnK2uCoX9YBUIK7+z7MqRUVvQKxSa2751Zewj7AUnuB7nVyVZOknu
dTETSzrcrDTUNi4FH+Zlew++0xwuiJenADQMWKzucj8a5GmUtyFaDUpYqWISWEL+
8V6sE9xMrID81tsFLp7X04owTh0qsze2+yr7SPiPudDYeEzrXpOiqn+P5YEhHz9s
rm0vUqKwXvAJC+xZc23tIwJ4/5Gkz+RysKOYr8H15Uvng//xzBxh9ok8ktu3zc3s
FNs/V7jdRUMg6jeieQaNBzYf/QBdIFhVrVr+JCfNjZqtAOkD4ksxwCl0WGvQk3XE
4mb2S0vnf1Z+4pXg1I/k4KLaI7tM2rVx3c8qqqlM3k9yB05FZBHaZeRQQUrhj/Rn
+rHNEMLlDG5uThkgS7ppKDTTcAjhfW1fJdRiJStOvCZJ7I21kTwUq3AORrY7MoYj
HnmrGiGHf1qOUrrRw5E2EhEYGz0s7O4QY5RxdsqhaCpElkHoWUtmfxEvnt8/JxZR
rNFruPsMUs3aPco2Vr2YoP/aSbuOENdRq60yz+YyeOP7Ip7WZPJK8HRp1NJceW3i
Km/5ATotv8lvQp9NNV+KlpRgBhT1R2oES95mQYSCfLwXpeHLyWcDNz56JNSjTbmt
R73PTQDxZmWTzy7Mh0f3oqC95+68pLEdbpieBU1qb6eT/K4Anxw6tTo9rfj8+JPr
7SBMGlDynsENKmd+5eDNztr8i3QKxI7tw0rAr4WDwMx2Emg9+qHRfcEtTR3e6fAa
qwy6V1xoPHzm/197uuQUBjuqeGNQCAUykHaiijsnfPE5jwMLtvo1lOft7KG9T1d9
VeA0AndIlavOVOgVFwf3d4NXl8c0E6ptBANeY2axTbedlR/KafsXa87KId/hizNT
7f6IvlprdXuAwgjvZEul8GBdk07vyuTF/1FGDXe/sPlDNnP+p9EfwPJ7TuPyGkq5
RifZgvOUDPuLx5sJl88K9ThnOq2sTMwlx7SLbmvOsSi5avyky2PbVQbpSDctZv55
iyZp4qcf2B+8BsZb+PDq1L4pIs29JqsqPTJ+qmWDzF0jgMi2Mtl2AuXfgcyaaSk0
gSn1L9ranROBZMorVZE6sbuf2evaRtG+L2GnkOrLZKjaHFmBu6qPq7ZMf29IpEda
TzEOeOHjLnK0J7jvu4KlfiKjyjjbWTEJthWAQrJhQU0825CSqfNI1gyeUsAswlFp
qVEFLEJ9vtXfEFMlErjR9QfS1JxTUS8emL+pRE34Pj7sDMHF5d3M8v2nPEA4wR85
1Awi3KLBbpFNcaPVXrZh6c07SrL81U2WrJHYMGc1EgymnScBIjGT7sjTyMoesarQ
yqdZLk4xGdkQyX2amplUT4iJrkhEtpgZLJliMkiD4iJNIOIvCtHPOCwotXt7quyo
stfsooJJBbIvWUpCdZskEDnsMRp0aylinVvmd5fdsvdCeyMkJoNnOtp4n4cxHD9j
gSo1mMdVTv3R7Ev3cMDBd0ig4DsuH56xmCwY6VJwKbuf4X3aX6aaAEMNMj0KesTZ
wMhKLFO7Iq33KQK+Nz9gX03avajR4RTagDqgSUC8vi492Lc/sK+UMF32EA6ledx3
cE7BDUuOq+uH4PsH7x3Um5fjeavUM//RBNcJCqnzUT4hdyacp5hQ8fGyZmlWpJQB
LBRIf9Bgs4cZ9CDPMzaVzOOjX1saU+9Wj278c40Iu36XN3mJn6KlzkYbT3OIWT68
+C9IigMoatG+C2pH90yZSrZYdOyWH53eL52HJdDIFUHzPRBNRsTLGmT1vDVGK551
Uy8INQtboz8JQEnUFFFP3EmRqOsujb9nto0DQ0crpBoDrWTSjBdtxjpgiDKaUOO3
+Qmd6GxUSiSxlTqLTVyQZCqy0LFAqGkqpo1gtZ+cnvhG65h+6mIKr6ODr+ifxN5n
knVvEb4XLHqU0SQ2lhq7s5PIv7X2pgMCBSiDK/7Tw5u4d3IKhX95B9TqzRlFKxUI
aPSGTYkm4VuCQ1FcmI+QHld1kjZao1BvI4pc4cJvUSgLHN4Q8o07dN8bYgdcQiZP
qM7nAmXLHxP50UyMONdIQUedXiIJb6svbAr/0NPiflYUmfo678AnXJbxbZmb5aTo
s6STFZE6Tbrc+u/w5da30af2Dt9a5+QddvHmvhu6mU88zlJm84c9uoV6IRHy8quA
J8ILuxc0qfHpoTH2AP0hDIXisxzRcEKvxAB0hLHCTTnN83Fb0h3xfVGvh9hVl3Vl
KTydGw1CTKnkMppcj0uJ7V2TzTqhFhVbt4zXdHQe2JbevFUMH5UKDMfsgzgVlCvI
EPbLuyGVtS6KqK5WmTIiCugahxwb0VjI9NKY6M0COeN+s+jsw6yKhVoCTFd9fe5/
BoYKa8+QYBTLU5uOE4BZhMy3op+C0R6yzsLc9wm1vMXEkTfUpk4H10kfur6HyOzW
mkzCnv1EGLtkG+YUL385fbkFLJKx5QlKaaHM01S9NxS+nw723cEfRGTQKGN+K2xY
M2B0maMXXS4Y5RbwTPNBqjbde/kerHwl0FVLL68hY1BfEMEPun+G1h8ILQG6O5o4
SUFsSd13dq+Zmp3ygngeJpfmuDLAmPSr3hODO002C6zZcGGE5TIQGaZk5rEA9tew
OKc10d7/4mi7hYzO5KqYXv8cnyljsMgo/rV54MLzou5vll0s7knwPnjOvglZcdpp
xX5kKdJnqr101x/TqfGFKM6Tt/syAq+lb0SDIcjgEBE4Tu1ui3MT6uln3L8u47qu
78gCQnAgdndBis2gugAZHAJbGkPKIokD1ZHOEiiLQeJdV5HipX/uYTThVX2boIJo
t2rBFDIdInE1NmvafTEd1UDlFyCTABAc8FYsVv6BJJdSvXOkE2IKVVZ6oVhiyjRz
YL+dpkfWAcaiWa9yxlkfoYGUc2dmjh9y2TH48WavyPKzrqhVdz2HHALM0VWSz5db
Vi/KFgMZ2lmNprbrqNnIiSVLhQcEDsRR2mDdBrq7seH1cLZigK2mch4KfCJOzWsJ
9xRb/Uf4u4TKqL75VT0InngKF1awia9Ug5480j0ffn7XsGfXM9m/zr5njZEmU+AM
8DxlKfipVUa27ZSVx8qHHkHTxeUhe3O/ju8/s9/XMOO7BALLK5ZkkqV3lfoPRtoc
uvA4Z4kx5fyU0PKEpwe/hlpPYrz1R1Tv0sJ8XHkG9a0CepulefRBf4psIrFCQfeO
NZhlyLrGYCxXpwN8Pj4QOlYeXmF5U5N/gDo0ykQSI1tu9f7levVYcROYDWtHyRc9
JB/i9Fr7Ez0/bWPPSGeumV9vC/dZaYeS1bl279r7IBK0RoCunattgEfWKbfg9BNy
xrfLpz6zNtLggI9zpBx4H+iPMTN7qds208x/5Ve3qNgI0+n6ykUiCWTAXcWc4Wdo
bER4/xb0hzKWJyWgVh86qhSd3UF0CMMHUTr1SnzCk0FXzVw0Hl6HkDyF/Q+mSsta
q+tnwGqAR1T8GjVKnB/qouP5FRLujZt612ELyGoPpST2J1W2qopDdIAMGC/1vdOr
D3H4fPo+d3X64pLgCVwCsJk0kzfJJmE6XWhRahvQ7J3fyPn5a0V6+LpJ98U1Temr
JpeADlFtEVYkstgNUbCYo+sTVVPljF49Txlt5+ObIrsvbsSKnqOyWluy5kEOkuKw
vtnLGJBIrVw8ppBXimdil5da8sOSCyYThvL1J2OotnmHE+eD1+IG7nyMQ+cdZ9Qy
P5U7h5wXmHlFJDCe1E6r0Mmv5nG8KCrU98nxTWgEF455SH+vNSp0/XJhv6dA0hJe
zqU6UR1EdVGylxCD9jCmi5FMK2DVg1svUoFICg8xHZWMi8wNqccZiQ2qJJp28q6N
C2xZUlsCesmezy3nuiRMlxXKT2ZX2XUsk+596JE4PCn+yc6z9QIOeC0dBUysFFEE
DjPvJFXQ53tGrxF6znAQto6QR4gau3k6zZI07pC+6Png1bYH7fHa6hoPxXOeqeNA
PlATgvHJFK/P9vMKr2A6QSKrzX8rv93706pE0ul2Cv3DxF3urDTAcGWZ5oYOt6OO
s3wdmmyj7UKnS/PGNASHms9jeq3GkOVf92qxDjLiU+8YpB/AUgLCpFQoHaXr8OUo
Y2e4cZEc9+mnZvnvyo5j5TjX1k4G/+oBXTb1MPOhEDGqhLfECBu94ogJIo6ZRHt/
9cYlNvpooA3N+WbnZ/zTjdfpkjX5Bbov3Oqpr4An60vLDfD/W0UcSfSbHpj54x+F
OtFHMMzVwF7mJKQq4paWeGLBOUAJNw+Y86/podjnzB2LNp2ivUkOvqJaPTfGB095
5H8z//UhH+sHf8d5oSTB8NMKfYIwXgORkKpyqUBXg2XnDw5VybihF25NIMnhggcB
l39ydyIs1iuNPZbLi0O5yrN4n+18S8Mw2B+kMvUJbQiKm2NBsLmE4WC6lz6Z4GJz
QFSLAhPwHel0d3+KBlIAb2GvL8gFYiMi4QL0mV8ZegopJnuy/SNY2lMAdUp+7+kd
eJcjr+ufgKUs1TDEI28nspgx3fSEtrenBU9dZlYcM3lEXpIhqoJhCnUiikL+udcV
WUEkaq0mR10VgVRc80hvcGJBsArTGoCJ21twyHztE2RZuIU/oDkrQlbr3IQv912M
WBEaxCi8BWTQqHDRVC57zV17/qCQPDwkFGUCBFAyH/rzMUqsvgOFtDjzH3zFMje5
BKJtn6pxK/RQG0ro0LyoUtxPXE2iHC4iwg/VrAqA5xHgfymY5WDaMT5fVviH919Q
u86tHJclja5SjZsdiakuIAZ8C1J1TrVbXH5fYDf4ykGRvVT+K9a0ZkuRJ68FsDZC
E4FriStSph9EX32Ckgt7xHvwIklIvDqdjFjEW/q3hVqeqTvMpB6VhG/ySeJs7NvK
mi+K7ZgeMNXWA5Pp1/ANDLtJCdMNjTexSfg8zV5A9LkXwclBwthJrJNI8/Hm7/ix
ywTxFwloJdEOeNog21jP6bF6WaCBtxkU1CuzsbHN9c6MMC4sKdTrdNs3FRszk14M
mCYptQL0vxihLH4LCoObg9c52LlztXRTu9uQg0/cV/OEUsbWuKaRv65MOswNY7bd
k9UV7YxdiaejdD8hJvDI9pWwE18pjBPZD5BN3QHOHHW0N3Ht5RTRPfcrk3fcwKSM
x9y9E7RIjnqww/XML3Zs/NXqpZLY3tH6/2sYsCcrmK6bLDWC/BxvlNJwFWM7KYO1
eGnP5/xYacgSLkTrFyYrpUAUQXn7SG9ku6EFq9sVsn1qLN8DXXAP1CwLqlzO44hn
D3vPhby0Q04jZThnxwUFj7vFxehh8TDSTojHujXs3dab4KRbBSclH6S6i5MwvKNH
4EM2nfWys8epgP9yp9gp0XZBsVa2mRq1udHkAV9p+loK/JNvaPStW48lOgyJYob7
6g6AW++Ll3QC1a2uZgQy2c+XUNYSIHiS2+v44ANAjPBFr/W5FIhx2gNJkUeMSl/t
r9YuKdNDrtDujXgCVi9qqHeY2fkLstqyje8AJvb2OiUG51garmwD1v/ANJ2nSCnN
dpghLy3rotMjP82RxDYVnnoQk3XMHJzA7y5q4ZrAYoSVAJPX8td7z1Xq0Lm3Dm5O
co9LGNdlg3Zae8yTT6fgK6/6X9OlkoWvH4vSV7p3rDZvfUwCEqUj6zA72Koq/tJO
TT7/ZtfYWoDOxNWyRO0FXOsifW0serQ4dyR0i4TNt419WgDf5dz6ifLth51RtPA4
7BF0KFtFPeJCJMzOa2BQUhS9l/PlIMXlgyN2leC51Pm53LLznunykPi7l3YXcdOS
khbdxRU7ZATXCqJrNKD1OhsYAoDymsgKjHR/2YHqmz1R+Hg2SSgR1OSlO764GW9o
ZXinBZ4WUmaQO3mOZ9xPk2Lh5F0Hm/t+fjN4zY2BxsXD1p7mZtGXKYSxSRdFDfns
mMyT+QCIC1R88htMEAc5JNwY7ZjZ7T3G3wx6PxV989U40wf5FksX0jVjjYTvDbMj
V3OSCtsvVpla8yGykM+2+DhDKG2drUq9sI5L86F8P21kaWhe/jfhjKVIOCB1Z0CF
30WVH6GKxYvk+mDhqW//H0S6m+nPR74HMBQDIRbfVD2FwNLM88roocFM30qkPUu8
O54W28VC4uEiihJmCIk5mgVUNrd0h2ujerVNKVxmd96OxyRdLDIRxMHRvnwK5Frq
y+8VyxiaeQMcVEZsMW3OBhEv7/2vemJjXOO7UjkgeNMoTMYbu3NaIngG/JKHkJX9
jd6O/N+vrplk+XamOmHGZTbgQk/Lq21nMKMRzJNxyjn6HkAPuo6GVwJHLPmfZhwG
7rIhB2QjpVRUGo5Jex7F79JE2lZUacJpAqe6aVhUt574fZJDlZsGWn7X27Ssy7RP
vD+c2PlD7VGoeK+1K+GYSJyFN2THD4I7mkOqvyjg3Vg1T0UrV6tICSL9pnT9KLVc
EvS/i62Kq4JakPelkCBT4oCYYp7vzy9PLvltacD8cBtAYhgvQQ7SG0fLZYs1xXcs
qboR+74p1WI+KC6uI4NtGIeOCfKHik8mb1Rq5+wxf5GbbysQ/EZhUW2jd8Im8hLM
4VerGZ3QcQc3U5i5kgghxeg5ml2uwRljmo4oB2oPeYhS8k85Ompy2jcIQnKqTZXu
7lfvyC2QG0mmZvdo3LXI2L7dvu4kINjEVwJZzRMVCNC0ui5mJe5i5pPWSCHZvWx7
OBjILpzR2joEwp5ZPtwBCTpB4ooXyzlnaoYmbTtFDbmy3T0K1a3ATU0G5ag66goo
54e/J+fhl4sTRYUsof605nKYdlUS4EgG/Hjn8t5/gWG8PLOO5PbiLpJRLGgg0CXp
9vBSzaXjZgysfM+edv1ocBFcUIwzehXRnbbi6IAIfLg/vfrLqQgMpouMNweV5YkA
M101mZEweuikcWRxAxxrVxGen+7C6wtm1/s1CbC2OI1shhgx+D4oXGsURHrOoAse
sk0gCrx/lblw3WJzSmC+TW116exniteb5YIkv0AUQkJD+tqnV/WkTF5JS5FvRe40
2n9YePBPasA7xHKTVeB8BICxauHOTJjOSWu0+iBmW5ZE3IikE8HIoWVnc1jhM7x4
GpM+2jEp7yjZPH7iNeue/EfH5OcrjFLrU1wCW6CuHx+KPj2GyVwWp0hw/C1nj5vH
yCSM5ax5wXVmgP5Sl9ySy3NvEqOiTQNKJ27bfz8qsqbAcGzxW+R42X3WjIEzhRc+
WjEKi/lmaBhBzHeRAQcBGW+5CP7n05QpJtlgEB4g8VMHh4SqePYSsFwSH99bM8XL
13qeJeGKhy2QcvNA33u3dnuffQVwYE4/nKPeCnN0iMjdrmNN3OgQJ9mitvlZZcH/
RQ8IHjpex3mg1sxASa3s2gqSLThXZ+KY6bvZiroMyAWqL7rXby8/uZ+Mo/HiffRi
8Dz8ynVjpKJ6jzG6Ew96k7y3YCQk4nmeW7wjYEdn9mW24/lRKTOR0fwFlVJk19H7
Szope6lpBFT+8tZmNDZKLMXY7ohRz9/3TvOXZC6F2jGRIxpZxS0nWnVjncW4iVXj
iaWJ7V9U1s2lv5DLdHwpRreadtFW7+6w7m6AT8Q7aQL/6QbVTyy9xHltybheZpsK
5QQpLXMjsDlTE4uaEKpUoVYAnoW1gx8cKa2KNgXjZse5417Ux+trULATEpydn38N
bNyNcbkkwT710lTCO5ntCdOAY19816dSLgOQMQVtJNJEqsb0tSADFu5+mkXKOwrm
GtzEjxpf0yXWyGK/nsl165nQbflu4oz6NHPcMAdyLAAW44ptt7x6QJBMgU1HdmJm
Sm5Uumto2zXvu1FQ/p6vWl1LUjEtjS6O+AKHL9WFmtA5syZBklQQ18IO9tKJW4D8
S+Ey2eLZU3MrAWKiAYtzeigLIu9uLhwi/pr1Y8Tequ9TxIYXiy48hYCvjAHb5diu
4KktbXP9GBH0qe4ldyIYc59Rs2NZBWqg7LQfB4+YHP309ppxK3nn/OT/Ymu03BeX
Astx8YEZ4H53yZefzhzbOM1G3eQclYGhew/DKVZbUZCYVS4uKZXfJYosYiK8O2Kb
eHNBudlGqFSKc9douKHkxTvOu9dAK6tldjdh6Qc3iVXTk7SC6onJhRrGr0EyBsxH
HaiXGKh0VuwZyr6JuVPcnaZaaaDS074MjOkHfUv6+mylFRpi8nOhX5wb0NaNSOad
hG2SmlYefjcDMKQHzgL9MQC+0+45BwT3cAZlxLbUhcMdyfk8S9vVuFm1GcuENYEs
qGR+Azr28goHlFIp6re3HOlvfcSVyKMC/Rn9+D6/QPzPdVjIL02LEMlJXpXNNMsn
hh9e17291w2pj0ssYnARjAwE03foGDiMhd1d9c8NMqZcqxAu3e7asZE9sg3JibwD
ZtUpLzFmQGaW/Orf+H/LAL4nCuet7UVkP2G6EE+fZo+OtPHbm/RWEL6gPBh9F/Ip
96XQox0tVuU7KGYFqg9OzVPluQRk09XuSjw7Fm7pvPvpKR/3v813JZ1sOT4BCVlF
Jzj9tJtYFzi2RbsmVBTDjfj8GlgSyLN3yeWMz9DvlO2hJSuKZx4L0lMTAe5c1Hw2
JeyZVwHHEi9paBDSj5NEi5wiB7ktF2wykppmcwcFzd0ISddhPBHuV7GZUCxiRhTW
B3XUZNg1Zu902sBjRdHMY6rcCQ1TYYH9TJRNZnarCF3IT/0Qw3VurkNKnvmg3AxD
WIdNpeP1v/sGr7+W78qhiIblpLLEGCrCQrEwvaRjeAQ7pdtsTOSwTni52C7cpHVQ
F4KFAv7o0gJ44+4s388lRKucqmowOFthm3iF3PIW3CFW0kdhxOwV3xMce5NPwyxb
PUqqsfdiW5VsOF7OVMSrSr8HzqzA3zoEZl5hA4qgDYNwoDXqLNQgqWxMxUr1LQcV
rV5iVUBz3qQ8rYayYErdFSu2GID4CfoOfj6YKdN5BWv9JiE+DGmNyzYsGDNI1/38
P/S7rDbL+AG4iSjhMyqSuDLLjpn5n6O+DQrqUk37PEfstw5XulVSt1/STEWUGimB
yIl3bu/mKQxw2Yy33LffUSEw+gfO1jkLtSUJ9fofJ8W7EpW1igfwS4W6PdMOJfpP
n4k2xcBchVjGI1rWgCzYiD83VbKIOY4lefgNJER1IfRUQ02g99VI54u/vhlz+XTH
P/ImaTpYeiZAav9qaZoX2SkW2RZGNb01DaZuAiCXb60Tjm4oaWnI2Da+l+7yLBSh
GPuqQQ5jNt2x+5IpLxSzHMsK7ljGJexX6r9jZeWDd4OH6SDeJrbCTR8uMR14WJhG
fxn1KRspR2ao+7F+gh9GlpWaJDSgF+q45DiiBd+mUtgVJyy3GLr32w/c85JPmPhq
Qdim3hWD68vbG6MgAfCRbnwpl9DIq075conm3XCVfXyJENf1Iiu+brdz7wCgMDgu
rSzFoZ2b/xpgxc+NNkFPQIw164ySBRRn7gXKj5Am1U97PRKrKfeq+v72HsjvXji7
ymza8e4eD+uXFVGRP+1ZlbXawJISP0MUPqAPsJJhfJMGOQLVY3+dh50zZl389F2m
Kfu3xczK7SIa+gxJ0Z/wDamVGb27kIGI1yhkWzF3dUwnCH9MaGyP70aGcSaAooOs
4fTi1cMUF3Z7Y3OCNChzSfASFRq8Kipyb0TkxBrxxEQngJnW0wVDl/Yh3juPt9St
CsN/3u2AbVh3810bfMW3edXCO9ZTvylifzlykgZQudKtQi8yKwS0O360VjI1/jW1
EPSTIxQmcCHtqUHNMLY34rPocxZfPksIHFiLTQK1Gragrt+RNM6YK7IzPHdgWQeH
IIpCZv4yDUPmET4zyv8BzvoF35mOI9bOBf4OE7mXvmPYby/sjH8BVKQKQU/TAAMy
taqlwwglZdVxa5XORZDohURE6Gtst18ub+rLw1/klXNW4+XemoOCSbUbPOk4Jaao
01LA2syWAQlcqurN9BUXBuVlnqPjO8qwGdpWCxvhPvUbi0hv5YJPrCRpMwwLiER/
fQZidarZww65StQjj2qekyikTCGb7L2R6jeMI184/WLevmZoxjCf7MPNfMvRFhaz
r5y4wkB8/ZcDWHMC+PcEtEnH8ocaYOCnICg3Q2cKMvymblnSdM+ZInuvP2j4voUW
uV9Wf31iimlMsiQuGwb0B5FSHcLTWNrbTl2qOUSkK8dvHw7qyLHDQ/oG5lxP2i6Q
8VZwLIv/C0D/8nlFQpBXVHXCmkVv2OScAHzBj6eYMDAM2cq71bpFP4F6zIgAtcvr
qorIRqLtnbZ+4lo9jOtlXdMCuAJuihp5el49cDJXQIV9EfaTrjDpQrtcLTOu7P6c
sELQuNONCoPMCrcsSa+7xXksn43fTnN7pEuqECiX72jZwtvFKXU0VyQg/p3l08O4
PbIzwwaetKvZTKBlqDoKr+StMQ9IASJ9gSAG/yqbZTPaot65ycb9dAVIp45B/pzZ
Buvr2LigiQ0woWCQo8uMpMLncNONl5blodbDbuBzuFGeMOKZaSxS1TVfgIxc8GxB
EUAX2Jggi3GWVIO1zdexoTlQBhe1w6jMFMwV9JHokNI7TtFkEmtwXyfrs+eqqvmg
34+m3+EIybQ2RFK1z/XSRdChXlRfdnkVbTCKohqd1Ar8am8+sbz6VVmPfGx2puzp
msXQHXi8JCsfVtLGl/msFFONneBVeyWN5kqv5+Xh/KuKLydOwRf+hGskDbXjAF4h
ufmQof+ojSLv5EE36Yaaigsmt2VQXMCQB0yfmPzrlzFNaN9A2LdovbODBBGL39cL
VeQCu2cSx9ro4zc8zWj7HpcYpqN0EMSNHD5mlBbUFCdgldI8Ggdt6RXMJ5SDrI2N
6oZeK4ZVBeu9FwUaB/FwKNx6sUO8lr4ZVjr7tB+VN3Lx4Puu4EbDZtQ+of5uB+WS
tLMeOh7yCUUnIARHQ4DOIxM4J/yg576X1bRo6V8Sr+NpZgfHOgq6FI2Ig5BQeAoq
xiL5Xja6AQTM6QC3USS8P31tMsC/DW1EMl7vCjlSk2oLAtrJbsnLGIo+e/99pNJZ
yITcN4wtijj0gkQHBPbKSVSUpRJuZSA2YOVMshwQ9tGyEhO8xfvVlcAgPSrureel
V7/jmawjlHqOsIUMb5HkAnHWuLan1GGqfeuX1n4yrs6S/RdNC2c3WkCqgtV6hQCh
f25HkRB2rYJIkWj5I5eIZlhmQtFUD2TczhWE3OgvrK5MOGKMaXWTPmyyX7odADko
vLEvA1sW8w7ccvZO5LXAdaEwkPvpG1i8Qevo9IaC8val6L+U/0dY1pZx5ULJOI7R
VZMZ2xM4AMMig04a9LWEPYPO+H77hcrQjo0v6/enYkgVq3NoZ41xzSymsO7jCYtR
rxqTRAjNPUzfMFA160PvYyj5htPQi0MSylwA+lgPCGvAvnQVOgnjoqeCGyTD4XIx
8/hS35xP4NTcvUhAQv7kMEuPjzRvCXsbH1fGcTaOdiJgMvlweSD8IfRVBAEuG2SM
MqKvWHeoLzNOijFWupbF8E56j9CHAndWIFju6fIGYMXkMgJ7QWNCPnApV4h8rpAY
x3BmyzE7wfkVvlgknGYHo1LePSx0racylJRYHPGu/1pzIIsVn+fgZUuq4kSXnsNa
JeTpJX+0NM0Rqd6FkaFOQgv8bP4lvIhUn/V/iZG+L53YiR2PM3ET0ejvDOIIm141
3/rq3IJ6UybYn+PMR1VIgmYuf2kgNg7/WaEAmqBZjkB7mkdPtLwNzvoLABCSO/4D
ZguzjNb9wHUiaPWNf6BAuYf1sr52p106/yOzP+NH5wO7LZgBf8o8+IceoTS5Nwjh
6y6T5uBQQvpgWvwGfH9LSenTSGSOKARFCNfTdeeL20O1ler9BhvDGmzK5LiWvIBP
s2F3h3pukeLGsJVKcG07S/m82QeDccDiWO048PwajiklMqD07rntI1ZJ2WD8xiNM
l9E7sn4JfXLmNA18XRHkDqiw2o6xk+kNSsiBtzdUEc1+HcrWv7XC5T3xfETMtfk9
ZF3VVuS1foYhopQJUIGgGytr0bUjSD5gp8o1OvgxzAhEP/bWWzU/PWJMLh0ZCByK
EGGLaEUzKt7vf2Jd/dXKTLWvMhyUb6VSkTr5ZpzS++yHj+DoOS9/NzGH1vY7zoK7
k8jI3OBOhaqiCORIWAvlkj452OK1U81/sqNE/T0jjdGURb97+IB8mhLjOdDlhLmd
q7oAwJVatOkWVJg+06FBZKKY25bSkEHjINgOGJ5D62nBV9LrkDGaMzKmUl7HVZI8
odLZhZu2tUb4wkVAufr2K7h6grWDn3OPblEOfESk098tdGziU84/yQHRjYQdpoxQ
VPyA9d53ronsC4qGOInKeDLihtEfabtf5DmgwKIhegswZ0PjeCeTjpTpZNLHGmKe
qQXCpyKKBQzi96LPVDBoFBbhjC01MRFkcjYUPUMudruqKJJ8wkWe9YvrMlpYdJ7h
sC9m0fOCQLvuj33RjkmD5dB+nFbO2UFk5ND5/551MCw7+WGPpONfSFRlLGDmy+GL
wkV4pT7KgnIv7eno1k2vnRHSOpUVKQs/hn9ZMfQRfAPCkQsgXebmdEUCxvprxJLv
yelBT9gqRBkYwBvaUBxMjV2fbwdx0gQCxK67ty2JiS3MEZsOKVDzWGu2DigloIHF
z44NsORdp+Q7VWprrtXo7kb9u6AL8+lSpJ0VDUfKTPJHdQnRE3lYLNhNDVQCFyGo
c6cwgJ98+HGYBky1z7Huu3t6AbMbFpQvh/m5/F5Klt4BV5oRIAo/ffnGt0Fis/LG
UryWtnF94V0YSLQ/wfU2M5ttqU/ChsZo4I6vUTnmP7TzAa0yA93yyssZ9WCKryMj
Oi9DPqsG74lAvnNUYK8cDVan/nqAmZBiNAIqMEnNM4xqTyWrQFMczGIVDxfvn9O1
oKPnNRU9DKw/LPy0/u9TuwA6N30LS9OREjoogehT7YDqDXdLqMaLwmz06K8RAWsD
l25VI1SGFz5qV1g+9e8ZZqacBxzVM1lgCGlTmmLtZmsFMk9k6tptNFG6qLDEe0jl
4iHN+jQDLQEmp0tC1xg82fFr2Vp1Yq+uPf6kxcxTNg1jVKljxDNpirN31gmzlzXw
vjjEfZ21i/6zGjxAv+cHntnqRPqena610Cp7a511j86Wyj9nGzWTFBK/mrqDUUxs
We2EafpKTpzR0v7ZRmsc85DZ0W0mMtAWv2m5iVXCtJi2l6J1hemAqJ6wZGRJ7IzS
zOnf06V2Ge7IoyoO/2EiLCxsvqJhYC14i8U6pS7XpKGOjlbjSVvFe0MXN82SAM+n
uQyR4bqpFlUwsy8/eyegk6x5z2DNd1aM3k5Ogwp7WfwmKineQVhTa4Xnz1DYzZjO
4K4f1ZWU2tMv2QJ3iiqkWBmqWOgbyOLWRUkMbfkAYXs/xQgrqOtwn48gY4RSNXEK
HbnqB/qT+8eLrBZKV3nwP/3KlGNNuxbKs7o/ORqZb0z9mThIky18kS3Cxhr6KNDJ
IZQXzyDrIBcA9AQ8TC5WMUIfyN0k1O6ptyOg4QvptQ6wfyBvwSxBACzxVMXop03j
WepU4Cdy97JVD3/0UbyIYzB+UBrTzGaKSza6lhDtH/ybsV1N0/okakBoZwKl50fq
QLZworLXDeYDkg2eWNacP2KKtlJH7HyBD3uOJfQJc76/hO5V3VrpyR5UjAl+l0He
dvVatrHpk0CdX49sdfYy1FLY6cifst6/7tn27UNoHw4QDVHzHC5I7tnuQ4LAa333
Qe42fjus0hz/rDs0epzMR4Ku3Mc4qtvzCF+o/9n0/1Rg9nLuRvBup0UJAKBjQtpb
PR42Krm6tZ5GDSAIp6sXQILtc11dgL1WlrWeegWgajQdz2fTFY4P9n66E+alqOqT
3b2Mv6VatogLJWC0mT7z7rFyIGQV4+vUbkUCPGpTc4VvIZJiKiBYkYN3PtBtnzQh
dLPjbQRdVXO4q7CLiZY+RZct6AI9LgQ1X2r/QyueRDEg+FOz720ByE1GolsLpPDq
y+oMMTpNQXEVc0/2cJVInzB70cNmDLaF2obK0rkIkAC8YepMxfKk2xFRrF+/th/X
lqwSaTDMlXggSnBFSO5TnkgPIhXTmFLDbCAi5OVryPlv+OzzJgHKu2NspPg18Nw8
9XfrYkGf9gwhkHAt75l5nVF9gNqq4w8FDBzQY4ukDffhYx/CjBlt4NMXmCcfkUyh
/eqk1qjpYX68cVCsWZUBr7BoJeaimZ0RGxkk3oSvdGjJBXCr7ZBaH3SSSkchTqIy
6U6PnD/HSBU5AgJXrcOF+3+PbVzQbwjPhTyzNUrN9VcZhCidJuHAVRAf1k2SUfTs
AkqWjj5Y7LR5Gha6NJuEEvQDNLabv5sKJm/g7XYRjDwvyePNU7XCL8SeYkRYch3t
9O8t3WV3n68ODFBVQ4UboW7ks8wK49re3sHqWHfmvRIoab1pbTctMFOAJxOe9nhu
T0ZjvlEuSwJQsJ5hyb7qR6QkSrPw1+6ZBUu64WoJbXd/e0rIZz6+k6zgTBpN7bAy
nKePCksOZmAFSNAxh4C/y6/XRKHzcl2oqfF7rBkY+jMVyh/3xFC7ciiXwQ1luyee
eCgp80maNLYhr2UCA/4u19RSdgcdaKHx04Vj2q5dhBYe1rN2sR+tXVXrYCTQtcnF
tJMftqhWm3+hLniGuKeQnxzK1sQslwwI/7IgHnJ4m+q8IFrAbCpkq5g6uF0LStAM
bfpOvj1fslKqNd0HepwOfu3lQS9AHFxAotbmj97YeIfsYoXWQoNMompfG5/MKyP0
I6NOTf+zajW29qqjhSJy6p5WsW3b6FlfJxK8eBClmpkJkLwzoP18oLPbZ/S5Erhj
bnqio3URKjor0Bm2JNN8ZXfzP6wpK5c/iCce7Y3hSr41r8YjNGRnVAL8PE4TcUK5
1gpUPxfiPsOCmmB3W2GV5XBrZ8Go52rGUBZw9mLCZxCHHhPBfU05WcEaAa7H3y9V
xHN1UsX9iyGxLqcOwaNqSWyXzr6LUt4dgBNxkLWzB3+Et+FG7Tu/xp0UBHo7xXK2
0Dmxm65jiSjcnHIbeoec08+GlEVa2rofTu11dDNtxmlv0C7+w69M27b85wF7pc9C
/aiy77PSugLRyRyfuc129M1Md7OEveeKELeyCcNrjoXL7oVtte2IWVRAFnRP3Aoq
rqy51m+Ni1NEl1eUoHh/rHO0hD3wYqvSBYADZmXD9MAYEkm/He2ZsHrRA95R9qd8
0af4lh9TFz8tmgQ2kwyreBT7tQGyggv+cG3kcV7SPj7L4uIcpw8CeUmBRvoSlzxV
6DUYE9Wsh/QjKIN/yY2S3w/RipzV26cDmW3tULf8+ITXFyH0Jxa3mBL6q7DVkd/7
NQ3mcnkY9yqG9mqsUXUjXEv+OngXd0VW5r8qMn6lMG+Nw7mN1L4sUtOzUu1waD2S
nOMFCJF/ybhPEO1XTajUbvyySIyedNwuhPxpEk9XlDq07x9GbjS7Nj0YfUfud7e7
kesoFfvJpCO0q7yZdXvssvONzFYCHVhLd9cYtE448pyxjPNVMaxh9RPRsycw22my
aJdbCvnPbw95JGUz/cHNJZOOoSFiknegt1CuwpofyJTH7VH573JpDb5L03PzPT7a
PMhqQ1YKr5ULOs7roIPrTi/AyMTZFYKiN+pF7QkaJdXEt9nEf7LByEgJ5b2Hv/38
OKFYi9yM1h5YlKW+0A/KeXcjyKfKBwajfFMkrJJ0Vy78Cp7+KTT7D43rbW3NZh4u
Q8kWZRQgczb0o2wtMPtMYPH50FOLSu6xDWhrTy3t5PzQ1IPk8f/doY3CtKyY2ULT
NwXUAy1oRsh7tepg3EaPPKoUDVSgi/a44B+lxjBcUDnCOqVvpJhLr7xGGh5O6wfp
3YyniGEA4amlFtxve6ZgdaG6GyzLU8u6AU8Qd4X3P0xHVgSp9je3B58HX4tA8HSx
g/5YfQQw9xcUblwagyb7BX3b4NwYG58m89bBCDzHnW3gHqmY8lNPwFPV7pJOc6Sc
N29NZohSPinIDymJOX43hDOpf/QiLqQ6zXn/lRDhjjGZ2WvXBSj+zYxh3x8dBENp
FXR18jLYsIkbxAPGHwGm2SXreDD8gbIObR0nBnUn/doRbkcgJNnK+3miCPbzXDI3
3trU6BwLE9kQHbwvDaPNmIJCYk3NC9sY7wAtKUpwzRs6ZghK+wemny7zM6COiH+s
dMEJbB9GPxb6rI3fAsa2DZj/0A7GERgQF/dnhLxNva+/OD7MZ88OVDNYqwMHPGAM
dW+E/jgrTS4sObeC/uvPSADLKjdsNjxmys7MHxnDcbO6WNSacO/saJ/srkk6pNcC
fUpjIR5YhTVlv4ASRQfFKWLs8Afwlesxz/9IOAxPM/Kmrx21DWDcY6b2O6Vo1RaO
nd/Tdpik6sAXrD00Tiz+L8b8ZNt7EVZN2gXTe0YINHgYUek6jQ1DR1DUm0doQ3ph
k/B3KhoeXdMojapGbCYfJ44PtZjhnhEg8ifQG3zmQFTLEKliITHtysYGgPazmX2B
txJ1snBCkZ/VfzuF0PnlXy1t+6tn6aywTNnK7oFuhF3UBv2RdHU8zSctpZEQQpGK
lfkdTs7Xaj1pdH4T4H4O58kS3PcYxPY2J4IiryGQbNq+AFC7ujWmdyZUvQ+F+3pq
BtQsprvqGZxkz71cNmYJqMJcJ/8FaeQxpEbHrwJOkcreyJg+V1HqEgWwIbVj1I78
IUHLrnuLeuRwvVZbHhqxJW3hAWNQ4i4SS95DU6vKXkdnXOfBofjpifFEh1Iyescf
vVl6Qh65TkuEVIUKH+bBCxKYiFDBfuZ0roIChsDsJNJ7WpzG0frE2GdpPcWcN8E/
8bhvCzmnQK4gg+UEevXTizbq/RZNhncdJwmqwuYPfchZGB+gyPnxNWNo82GYWyJp
Mmw2hDg8Zz6SGHbouUWr8IcEGa43rt7qOZb3+eytpE2ZRY+x2kicHUlYjeuknaMs
+LQgJ0SK0zHyL2hBcRbRsLDBpGWom9uMA6fzet/GOzr/IW+rrhvtsx05E6qjdHb2
NYInsCn+T3zbPnlSWQbqurWyce9wubVyDzI+nZWZBOmmdDamhg3dUOg4XXmz7vhX
kIz/tgZ4F/+kMokpeaCvc4hEc6MS/m9LBC3Z3BMjL3dfcZdbzwZSr/Rv7n+MRqli
aGyk+DeCafD8Cae5ioz0UqTRmDUc7/wAiVy4NE+Dco6sbUAGSb7akzjKCPGWy23g
o+L9fRSJr/Yh0pVAg71GPzRqJix/bCE9FpIc+a8UP32zWDutDY+YUXU8Nt8OSNrd
knw1Wl5YjRMmgXReNYGlWmoWQYrcx/hZW2V8KwtQ3cM9/T+8o2eM/dNwwAjtM5fa
LzleSvfmgZa4DLBAcg4+05f5R8UCxVdmjXHem0R3brzXGBLsxy/VKomma7dfkbFR
03AG4KOT8EPPmvZGAlBw+eHCo93eKIFTRaNS5AniWUasdcjYdG1R34uQXmdT3U5+
/sf5yn3Hh0iL6MldZ6zUITXHyIYI0nsGhCokcAQr5+41qOhCAu86qk2zO5k7gBYs
33u8T2zvwW5DI82rz6OiYZB9l9VqbtFWGrTH1nIzzjDVotEBBkS/hDhUMPnlZrBC
1m0NhPtkyNacEWoSbhTp1MVp0n2v6w2EWlNjkw3RS0VBLlt4VOE6Tza2ovEs3ydA
8Ra88aM99xGvBl/MdHuY+1PG2OEnaQtJY28IEmTISVjrMHH35ZpN+o52gu8qVtfI
U2IrmN/Uy4pAqwNDfzCCK37BEBUWbPhF+QYDPBtV8ny2fXwaGRlK74VngOe2qgYO
o/yB24aFvhrOaIZxeXzWTYn3UQBi06FR1YO3a8kQSf2OQWxqN4uWJhvf/ulJymaF
V6bNXcJIArjxaU4t2WiQfc05OcDumwyPfV3sgZYu/6bhZyXe06GA90rQp24T5VtP
xm6izWRYfWBF6aYXd7+4MEMjdZI5/3H/x2Elu4Mm49QJgyvO+i1gwieL/9TQwoCx
yxLAWziBq6Bl+vl8Uk54AoX81DeTxFfhLeS8J6Ka9WQtotfXhrTpER7WtZuxMREg
OjkBjZLyapSrx/GGHrXjA6O2I/GiJF16mWgEPOuWAvL2A/ltm3KIHT5lYO5pmWC2
mcJlOmP2c1twd0s/aLqZIqs63M8pHKNOV6qThVfHWn+UwdxsPdyJN54Pes++Iol5
MLsMtywAAtXJwa9sXUrZCiJjq9WYQ71KmzY+UDjuTxFwNUJNqrcuqY6ac+Nq5toG
kxijYUhPMVB874+Uf49WNQrTGK06D/K5lS0ERhIJDI2SPnzQD/sdteiolnJxI+i1
SvtBjdY9qDFmn4TPhOEBXAZzxUQrkSuHcArsSqXnLjAag61NrC8+GmM6at/fdNeB
4V7ss0t6oenr1VzJCHhfZ/tCCg3bV5vplE7b6X7blfekXA0yNVMQXQcrMrJiTjQ7
fXNuwthiTI4cBUkn1CQ3PxENCRqYD7/sLOo2HGr1WjZunA6R/+lEZsbxsMnXTz2p
laAaGC+QyMwGEwaZqHzQEiOobRr3xJURlDF0pFMfDyYJ/NSmtG3kqodW2o6A0VX7
Wg7IhqHbYUUDcdLFHqO822o2RDlLcnYS38OASkEEJQ3K2wGl03kf7H4ZUk+E9tzu
WrzAZP8tVIT1I7Zc0Fx2bcExZUtXaBkj11iQZRVp0Wxl1SD9cIwLQlEOTj9425Px
kR8+Oz7CQ1n5RWsyXWvf+nKmD+ZTKzPDY9RVxzMjTSaGzIVyAjzgCQzi1iZ464a/
4CckwOhDB86k2wZSwIOgYxSaO8Ly1Z1pOMQzhmt/uJgZx5LKGd4bAXFy5eTe8Dfh
yX4M742VIJPS0+kiX3lRWUW8cwx7UKbRrRCdTMrT9U27UXaBQsCX4Ps6JIhPZqHV
rPkubQByoJx7ruvPA+s5hcN/SZa4A+3TNVGoTR+dyGs2Ahl42EWXZn1BHds5rtu5
KwEtQ2ChI9V1djE0/J1PsJjbQnkVCkQSnisyAHulTWrm8PNKVLxCKBZHZsNjFnCR
vvEnIw02IxgZinksVTMOsgxMU0FHJuGZXWDDIKQpRveBRjiph5H49+1uTm//cIWF
IkEc37k6Bn9tu92IHcwofU9r6HgIvcleA8Xw5dk+xsr58iE8+mNBalSDQmCABiuc
WrjhZZ9UQVjWptGjUyTArPsfg2yGY9pNuh84bF+cGG31XdXJUmpOhlZYwsHnOhWS
l2DFTzcs9fp30g5Cqs1J7hWNzVvTyJ5i7zhyxJWVcPQtSj+P0WmKNxnJBDfCXnud
a9sB6hzLGul/kyhMKO/2P96QHIYy6X6X/S94thAQiIu9Xe/4NcgiuXGS9pWW8dH/
VevY+YyMHgFB1x+16HAMeM+CCzLGW4s5VyTBw636qVjKQnRPrsRPERXCHcmpHnZD
RnkEBMeYggMtip4bMXCmECIaBMyvqNMNgXpCDiw3IUIr2We1xOond0D1AT8BhbTB
w+u4+cp7Cuy6n59iBAdkRDMwI9RJvqRT9/CMKFopV8SfXP4/8T7gaRjNIKKvNOGG
Yvdj3gzeFsTxbcj6RE4T0u6+6V9JECXrUuOsDHXrFiwLpgnNB2r7MC/03MxZ22vu
0bnJVj8lRUk/1rCoQ7qfMLf8itAJrDykq6ZfL7DVgcegR+MxOSFRNu7GOWbsxaxX
n3AvS3ti3agQS4RfikOAKQ+j0+PJYixi/VSy3isGtb6eJxZA/aZkI5Fo9c65/LIX
WVJr8/hgX1QW7+l466kp70wzgOfwrBpS3nnJPELw7YVM3MNj+/YBtBH0CmXUe6L8
UXgpkJfcMmDYPhaokkMdQAUX83931c1k8arMviHWbtzr8+0eCrmgh6hbdgjaV6K0
oA1Vo9WGU00cDJNgcIIpvF3NdAP0sUA+LyQo/WYUiD34Ux2508lmNFb+sgQbEr9o
QrzpD6Z0NzA8JfOuEYLNUMhjsMyo8UVSVy2+5VI7PfN2hltEc5j0mtHCTrXnmBZQ
e0NRY+wWJ8qqjSLyXlQtCqav+q7LpQAMw/sA4m/8I8vLQhRd7aKVP4QECD1PAfpz
/MR6GTOVywdK56r+sb9tyGGJjoP2kpFN6E4vjbUXySiJAihI+Ag1GQ15Of4SZPRm
J2WkRMNMGWbeRzkWs+c79kYBwavqR8urCCdMQUCCNe4uoqbt77/40WztozEQlI7u
MDHYpYYqOejnUxmh0Zg+dhbTddP/nxze4U7Q+3dJAFzrNeFz1k/PmE6ZTBSYz7If
uh5nBIIke5XIQJt24dqHvyUwpyPVfZDZgzwwJCGBqkKIEXkPged3iYzYk44VNjmF
HPc6MBlZ4htrgyXSaT2xUbI2uM6ruHEVvxnOQUPuMqAbyXyHXTe9saqeGD2bxH2Z
EGTIjpl/U8FXfDL0SUlP25rWN+19e8t1zLd6D5UaWmuEyulQD90qfVUNpFnvS6HR
TnZNekEtCyDzhhaDwXYqUy822NoRUAKH648DJ7BrRujNTJC85B2tyJ1GEZDTR4Ia
Eq6HpEc97oePDgP7EcJ+TaRqnWZNMreTTa2taZmPJQn505lz1ceLTcjONZ9c2Qyz
O93pGhqxFWckF6Jf1VFlTnVJryJ9WuyY9itQel3lKnb4QJf+RW4+jAH3ZmiJKAKc
2+wpRKTAGa4TsSB121+OJhMXVy/Ss1KOkvE6bd5FKbqMgrD3H8xFY6lcAsgbcgS8
gcVWb8HbEUrqrZC3HOBlTB/DysuEbpOms9HOX5nH7VbPRQsy53lv+GWMkzlmVe6c
LIaKhBIDxNoo0F/KHWk9jCJkRv/lE2WZ4KOhY8hQ5aufbHahAsk8cVcxRMm+wNw7
wEYh5KBAQwZXleWa2w3wVdTUwEdm94Okq5b9rY642us/y5n9LtodNRWhraeL3DKB
nve6koFAz5FQKoJEfgo1ScBkz0dQKnxqzbwJUDyM796LiUVTyniHB8tWPWOvFSqy
Go7rN4k6tzD/y87p1sMb/738dshSGsCf26kcUO959hlLxScQQsGXjzEcI5nfMX//
avBKaZZnp9jQpjTxP/nksGQNiiSEe9DuyHHpYuRPvdm4tm+TQPIp6AB+2/IUCGV6
AlXqWxBRf5r7VL3a7HTY2HNUvpeNf9JJRtTAPrEtGdtjDT2EviAR6sIWIpyVehwe
fL38aA7GhptK83I4t5tZRQhGRiJ0GL1V57iNqhrsDopBi4OZNHD4AtrZPP3u4vFF
JxrJu72W6/a7utHjDpongnYnjzYoAFfbZYmVT9t9h9LjsoP41QsTGwSUA9YRMQvA
Xuzmt4PbS5SBsKyiky72PSBudYQ/2s03553LOgUui/knxYgyvdQB3tROhTrT6sB4
t2PBNLWaM+UvgY8PC5ianYJUBONb4axShbTI0gzaxR0zy9tLYPp2297vi8GFW9pm
808m5X2cpbFva74KZaWPlzBXszKMtWOuUa7Z8/mQVQVfOoOKVkPfvq2VhrEMjlq2
edMEdRa4msTPwK6Z9///tzBqFSTcl3zoxAWf+2Abwgp0DiWnIC2sWr3r/qCFQYjm
RtT6Xt30RO2+nAXfGF/PZtDLH2H/2FQjftZSBO184GnMvOh4EFrPK/6vY6ffco4E
EUE6bMTsz869XaA9dTlJUngksDa90jNuPJxYbsTk9B7HOtXk73QGYtokG+zDoLK4
i6NZcLuUaJyJbQUqpdDRVGZswl69JNQkReOph2ob/WF6zkkPd+Uy4GzIPfsmHc+O
u3TEmyTqyIKdjH1DBU8SLlmoQt8P6LaQvr7nEc11A8UgzhI0auhDiJpbRLdu8Xbx
QEG5jRNRpG6TjFz3SbVkgzTaNRyqCZUf0EW/JqZ2fmkppXGMJ3HYyuvPC1o/Kteo
vyXIA/n6ucm8wnFmOE1uHRK5IS1+nZ1IOdJUFJJCLsV5bgkG2yeLojSs35cdmkgS
+VQTgPnAq168tRDwNFT+LjgyvsVbysz9E7jNYRLGErv6Od8KiKv64uB/aSc7bSyM
ByQeqraBXrjzxsWcb4XyQ0NypKq/veqnqceI5wuYR/JB9MfyHW7XhoVGuuQjuB7A
8w7rbsFxasxEtICjZBNv7BDOUBjq9TS64digBo9Z1W4aYdM6Htoc7TUqsO0StymM
LC7fYssdBwkfC1zx7hoS8+GR3l1TscGkwvmSWWkLT/TBiYqNNoDcwtAnIZwnhFuZ
hiKk2PKQIsz0HE3Wlwj16C1YFRUEsAJmHT/H/CeL3lciVnuknlJBLe0KDsnJGHSs
0jCnRLXW4sUzNCji+1mn1kmTQFYXiq7wh8LppUJ+BG23YijQF8L/zlhxmN3DEk65
Zbh+catSwggL8XK1qZReiX83GMv3EAGXhvLg8cb4o8ZeMPQq5WZQ6ZvJ/AM0S3MG
oyS9I6O7uOITYsPuj3q9v7wR6hLwgxmiHCfNE8otapH0wghSYWY37Vn1D5McmQ/d
a4RVcXHWTMSkeqhJLTfxSYC4bxln1dIiesqT8l+SJW1AjVLgRvAR/A5A0Se3q5vy
thU1d72Jj8HKHjhK/RhVpxt2BWs3HSnhjD0/zWd7FYmMfmo858lCh+zT/lTBT+Z5
VGUJ6ogFg7tXWnWydlLTPM8LflTOLfvu0hpqV67M++o7HC5r5qD+flacYuW571VJ
8urT/+5Pbzde2pXYU/fBL0mt2koct/jWaLX0ZYT6lbbkRosLxtVdcmEnKWN6Tq2Y
DWPUFO3y9XeRus1ESGDKxgzCxUFpGsGf6Cyj4eJ8M6zHgvz/BsrdKuwKCiYm4nKx
tNP8TWIjf2dO7mfmPTjuVOdkmEbmPGqHSA8da819kYNyLKdDft/yPbm04PNwOo6D
1P6oiBGQwXlFHq59drKYK3hRaJ2A5/u45r2cJKY57gbvkGfuVxZShFTgBUTkYfYo
LaY3y/W40wX3SX5DmqTF+CqMxvVWM8bZ3aCLMddeu5mVm6l2u9gBlGoKgWdBXgIi
sHnUvjBg1HQ9JUZdOoCvn5i0CoL7vr5Bifh+B8xFPXCjMKkibnrJfcZVvW2uxvtG
D7YjOfQGR2P3jhP/6ylYX0dWrCxh6qgNUXHcX0tAFEZ+5c7fFcL/G71f+r7Qmxz2
ykf4Df9BYuOB2kcdcaXnqxl10/RlUgCsXOdl8/ckOnFHp2ls0HVPNeSxLg/2AS/m
DY8EFT+iO6JzrKUEHjoH8MZXV+zvTvdzAHyj/4lvkCuy8HA45zt91PUNrp4xa5nu
eAhTjfBV3gxTSr13fm9B6eo/ANx43Ux86Mx1vzlIMsZmM5MwKu+0hF01QEyCIXR5
WB82yvgUVNQP4PKAtkm2jIpMtBhb8K//ziMfNi3STTg663dARfSSKtoTtihiDjQE
Nb5RX7k7ekV8gB5XCOfkx/5wn64KteIwg14UnCmb3+7cMz+gH7tG9zPpkX0aGNEu
GU+OTWnMqTdx59PUXey1B0XkI0siGVXjX1IlFRYiN78rqC/npiexythzV3k+WZZg
CjWXGRfAAs33vq7ZNUnkQIT9W9KaBYJQzjDkOjjcvuy71p3zAMhYhCHf7F8wHci6
hdQB9ATIX06lLwhOGMYqXYMwXfBDv5wM+BCeD2RcWCV1pZcl0E+mwGLAE5Y3eatE
lGUe4eisF5NE598DK8ecAAJr78FoTP4+Pd/SUmBY3JW0IEyHa+46/A/vBQEzImL4
qfx+ISIfOIg4zKRSNb9/l68lvok6h/hBqddO69BZLzHrbCCOTz55TzAkbCy2KsqJ
OeVZfcj90j0/q8UeC37T8bKa3GJ4IcI0FVuQ4+Hbnx8Inl/8sr3IIgVoef6XCcjC
HPVDfmrvkeu2njjsVIjqZlyy6VmH1had0N7eOX99EqacEwQD0zh9qQO2bRbgp5CZ
r81jPUvCi4zmvMbtoHBs8SYY85Qmj92cSajflvUoT3/6GR0gC7Ytr2Cz2RDGhszl
Hom2rOQhr71Dne5uCv7cehSCivlCgBrIKLUjVjMLi+vsQcwhSfSreUfsln6LU+Js
WGL4NpPpFJ3t0DyBD69mS+GrsN8vBi/j9yUD2bF5VKWbxu+30+ienKzKfTReszUi
P3jH9OyXxzy9M/1L8uMHAEvpwtLtGJwXAfvs+hHYKwYSiqLL1Ok42tuXmSqUe+JP
yODF+FR2S0y2rwdsSnbMwiAMicJHsWFisMltiq9Vs0xyOyIEzUhb78HyHRci/hvk
FSlH2rPhhZ+Q+OWIEICviqHJjiWBi4FLLjaqRa9ZjMWVu0eYeOi1xg+6znCroBKh
H/9QkZmJAb7n5eH7xSwvYe66wzu0NqSkkmFZSfADxjPmp9vuNYzVlf7NEDkj6K8b
Va+mnrunMnejxLArgVCz8SQQm+9j9iF2d8vud1dlrS53+Mqb+JWYiYyLAL7Ttq6i
jc4XNbdBvFSD9L/JHpCN+EYWRpPY2AW9HJXsiD39wDLmUzH67sVUlhQkj0lTMcSk
gts/mq+9Fl0eqIa/acb/vym7C+/TfFYTpCKpYMOwFF37paQvYO0vIN/OI2sE9YG2
2M3hXoBRAAIoLi5swdPe0SuU1DtKwYPIEtWNIODS/wapx2MNpKaDzCE763ZbC88s
0xYToqxpIflcXT/sP/1FA+RDlsm9L8wfMmWKlrlhZiD/p0iXzj5fkqBmNw9zcdZA
ZhSfZ7hGF+XZPFnn7Jjdz6uUf+0D4K1AINaAprIGKkBmCtzMO6S6mZeyvJUZp85F
h/sKP+io482rqeTtKESPSTRYubI1H2+Gq2wqinyh7odkgILXds4gqG9XPqSObVq7
DNDmUvUe/6MPeW9x9HWIjRfJKf4VRoXPvIQPmjaaGYmZQNTjCwz2gfwcWYBG+yCz
/uG1agkYfgL6fGn5EUTf82sBVJ2ZN16qf0aayu9lxCQMi3742aFIKfyyrnE0iZfP
/7tbuLY8LZ6BTlfBx7fnDrkuEiQUpS/JdD3LEa3BZ+l8tBkASN60k9tMaYrJba5I
pZ+eOjv7UsLOHNvACd7fFDca0TMngpAAL5xX+OC3ZZ/6bEnqMPoIcTLWSpaQZzOe
BStNMSNbgJlfBTwWqoFWZi/f8/HKYcFnS82PwduuwWTmGW8wNP88E1QMnYAcxwW8
wi1I6TmYH5vA885QGsFGOrqs3bTCwFZ3NzDwIx1EGfjCEB6rUhg5DnuLWxNsHJLX
Rgqv9ubuu+YDKnA68KQdlDxemg0eCDh23gWQAAGJa9vTU7OQx5nK16v6BEKZwr7D
apXYGs4EhYQyW5PfcaZNezXhxdVVFC/TrBE5qAGGcoVQRc8of/yHkER3mg9nEgCs
c8w3wN/RW7Yctxxwf/8cLLLNzVWrHxqOMZ0PgPmeZMNX6nnp5ZpSivPrUMAlpfW6
7NXhXTD3JD66wEGpGR9TEBcajGyuO6pm4MObxhGEb4y5e3DsKc/5XijCzWWeQJBc
5oQ5nFCoPDC+RDkNE1UuY8tWdmbXytZdRhF9wIH2OxnkJA/0XHwl2rkzQ/VBrNnh
S8pxvh1QKzuv0hg54uR0KXZjPhoy0DxKlwviPt3tIH54FrExs6sNseQY5u+5KIvV
kTQ+/E95yK9KhyqrKc+PB7lsWA7aP3gE80c2J1hdAU9hL2jDZZzHvD0j75RgK1iD
JQlk5KKgvWLSA1RfsCbQgv3tyclQRATM2wg4nhzqH7arO5dIuSpbZ+Ug8JTINQAG
2S+jv0b/TLhMSVoSJ2/X372ngS4UWwQXe6RtjZVjL54jyZKSMUXPVLt2ZxLKk9eX
b53M5KYAMyJklGjUODxEws41ipSruTmzqOPgA4lXETxHOHAsrGnyf6dwCCT4N74Z
xzZPuNpHH9kAR8ldO36DvSkqNdxaAsuIqQugtEVALQG2GM6UuYb5cGfqUgJCG5Ow
Cvd8zwbvq/cuSZreQkqxNWh7YvNjvTiM+5bZKIQdz4h7KUanB5eoBV0CVVl37+DZ
wSVpG0T2D6zx14FlV89zctChrodM8d10tSDLU1nASgznIjNY5Phuwj9rwSazS+BG
pH5AuN5YzTkcBcXCNhUMqBQk9YX1Bm0iR+X4nnhDzX+4pxk01vJGxHzrQAS4MTvq
3Drtl/nNKuXXmLpVQ7rq/YBupJm6vv2R2kX/uH6Dsy6w9iXzrEz/uti+hoeXW1+P
XDuVN+jW2UjgZoLizlZCF5zVzYXW3AvErS5oKpyNF6701sdNMXUYdenq6uQ3EOUG
5yHgdDwpIA6yCoTQBpxnEfmn+3zR9uSttGWG9CzdKZgwdYGqbpxzNKaZscyszqK4
tCJFyW7FUQrrmcKE6OTKOvu8hoSSmPYtT0+bWxpZMWoUf0KjDklESNKgolADUppN
SD0iHoNNg17nXj6bi6LoFWmv5XdFvR0dMnZnWhP9x+YiJc4xQM1HbSqcf/7WnZY1
lZQTyOkykGVPnCZNy0tEXXx3alg4EgH7xqkUtbBpcmJ4D+iK70fxZNQU69st9RXW
Mlp4dDTB7uxqTVTShO6vRaUbNHWdjKLX+mdLvTBYMCXS1PxPCqTsfRzeIx18fNlP
Mcy4SVtTHAVchubZVFWLh0/fdV3UntJv5pniPmC6s49ij6FTn2NZGbORhqA13gTQ
JRNGkll8Zo3R0ClAZzpyWYmSs7NqrHgFmH/Q0E8XfYo6dt2DroiF7xCbGDFOxKDn
U7DG2SFp3lphMLP43bMebguON1efzJBSTQKSvipELHnbCn9+BMMX+uiJabKZbOc9
oXeSbzHALwUx7Ds7IGpWCET9J3ObbNdOA6fg7w7RBUCXb1B9M4QYUPxSFoJZKaER
GLwZFTRIqnDuWBUJc8pNKNx4aDlq2tCPE3kI3xAa+S1fkx0lItufgD2eAAGFYk75
U+Znk6z7cR6DuyGr1Dbt4ZtjRe/C+GHl5jMKlRHBKVtBChXXtTFtdxgRS/Nu2qH1
wVE+9ZHZyr6VvBbaozqhF7/MNphIuyHENP+oMoTbgGk0jOLeW3vwXd+H34WJeT0C
9skUj6++Xc4VHjne8xeE2N2jN/1SEjvggcYrVI+mLx3rOW/DJD8Kj51B+q3xOIXQ
k38XPYCkGPXwNjYUI/h61AIuTprJUmxbWGLYWbdwv7guxG4v2JeLsl5RLhP3+XsU
aIsN3/DQJ7cGorPEoQHStQaC8mdlEL4G4PwARdbntNE7jN+3w6EwVaAbUJ8PZbXS
BnkJfDA5MmV2GbIVD4bm/oYAEjRXlgSGlAo+HCrHyHs7uarr17XLfDJ+Mj0YHSTl
FkO9EKDF3DFMrDExENTrMMShWhhPtH7qEYutFbuBV+nct6xpAB+upNWIfoR29JFq
tzo3xLehWi8uO3hLB6q7pqZYezIPMPWbxPHQQYB/nmGOR+WFffeLnbfh5Mfsu0AI
4kaf8orpNiEvDN14Je1cmJP782ehlmz8wxfnZ9Q9k2HjtaVzcW8EUzcMF/Q9fzaA
mS6CnIml2uRHKkZLdxFdf4AkQaivObtt9M0K6E0dZbeUUntGy5YXFHvHD8jTo95m
87P+GC6OC52Rj7KRV6KZb6AVpRhcNez3o47YGl3CjwZjioc9JVnGmCCIzafIISnM
gyPiaycOvkb5QdfY69ehhc8aJf2N+Dw899isAeeOlAw8uYsvO3Qcdj8FbfoOEEs8
xL48kjS1zu8kSZKnNOhH5ZpLIXqVnC1KlyDQYQ+Rb2XYfpAWlHDRxZtrvLqxqnuo
m+ETA4gIUm864efAxESaszN2gKqAJSNO9PwXRfrd0Hhub/wLtYT9ut+BfTf6rGE2
6a+xNrpGImxvYSrBrICpcu64AYal3f6kl0dAy0gfX8ESujQdZN6e2/+wEi0ZO0SR
8oRK9/hDuoa3RJG/FIdDop01ysryQeMu3tQQ3wCjrIQ0rHu/UdouNq6Xo5g6EJwy
MCrCtk8rTSNsmqT/NIHLd+kJxseN/c4XL4maMH5B+q1/ga1PYwOzF7BKdt5sRAF4
hlWL2jWP2j9tAj3CwplXwcgHHnZ+AJ8znYrO9jjWu48tEZSRFuZ4qeuJqIKm18pE
1DMeQ2kiWKs+Mgs/G24uAw/giepJFwXZ5OqyczPsspCrQFEj+CmcJjR9RDnRgaXJ
7OSLw7sbhk/hoCQ3ZyRXamIzRv5uyO+C11aOkD5z9xemoZjBEmrV4hDKKMWouqKq
XYCA5MOwXr264BKT1JThE0Mx0s20Ak8sNrjL63w6g+4BTpYOYh3z5d2X4e2Ssqss
pfcjWdOd+5KJYD1fiztWNJaByGCJ/d6r7C0TGq+pud/q/dMdQJJRHhUV04ILxYDD
XtlBlwgxtPL2gWPq34DBLP0w5BZnwj1wG92pDO1NQB+HwjFZbz2Zl7b36aL4Yl89
aDU6g/wF7PDQxvNi1W5iaLB0As9OTp0xWvsEeGqdbyrwYhh9GNf+YufG9naB9tgp
Hn+Rtsfe45Rr9moukhOXl9eYDxnMxY2ah1O5Sfi1ZwIqPtIsX3IUT2Rh90Hn2DMg
CnMc+v+cA27Bpghq2XsV9Cj4sZ7suM0Xa2zanjvdf2/ahLtfqIamCBAPxbeST4ud
kvFdzI9uuSBtchFqmu7TqP61RxL0PlHGnLzh3jF4+B0LZNIoo5G/tWnH7Vif+lpm
95SGoWvjqcMf08c99jzFJ66lGVfuR9bt4DtIoXMx7kh2Lore6bg8HbJ3lf1pRuOY
Y2a4RXyUTtRN/I/m9ycw68V9rJmQeF0cLkwNHZSB0nsdw+GUajMiwirawTfovsYk
uStPmtGWKq3Oy1aieNUJr3nXxRvLeF+3WYC4H2iKStmvI7snsKqrEQJbkHCEQQs9
cPmNDiBq04qcZm4Y6bhSrY15orm0kJ41t8bMH5lvDguD5sqFPUmpGyQsjo6hp4Ds
UWATsaGHh0wqE76gbI+VtpNlRoN7oNQqAPuTIRzTMJSDIEp63slKKmAdfJgjpgde
OQKgtdkHUdqVgh9wzbDra4U6JvS5EG6zcBqvZ31zw99ELlQXrpZIoFXLF20KThpB
TWj6iEDPKrEcKRm0QTCRrWRUb5lQI2MgVHk1mTPJJvt34jztAKelKoewMYNRHnIG
lr9T4Nktd+9sLROnqBbSWTqBHBTFjKFLr6s4vLJqdiqzTiyz0aPUcO5ll5zyWvua
/bOR5SV/zsO7jXAPQ2QlQtD0I+Ad6upEqQhygLIjfV7pj4qBzYs4Rcur8GxB5MoN
IVJqi03Uch6vzjuxEKAiOoiuSyCHCEPXTru/32z2SwipZk/5Bm47aoIbufJWlRcx
SvTVudGNMh1Xo7upYnJ5h2DgKTODD9hj/kjlprGDEXDTsNVOXTdlJJ53SZKNL3Sr
0TfrN5Fwkq4UeGLXfi8/48KtkTG8zmu7/xs4XcWF5Tts5mw8x9jz3I77gNMi5E/0
eB+yo/Z+CmS99yyw+MZaKrESiibu6ZSAjoMvqfi6OeSKinsB0KYTmh9KzWYwqfM7
IrwhLiOroB0gMrRWB/wqlIVxSj4mSDqwR5JA8mRVJfBaq3B5QRxbjB3x6p1N7X3/
kT45vMRtou359OPNviLfYDt1/Ee6Elkcg9o8kCipIHuZZfBnFPuWW4GBRgUJsiTw
7ZK+kPnsP19A/kNLHCWD8UEKycoxDPUq01IwwbffibubLU6qD3t+7vznbtLepQgl
FmBBLP8aURAWgEQn0mO7pEu+Xxbmp4/Tx4i68nQRAuZNMv5PEVy5rvAD4QiSH0fA
SNeBm+Q2mtTZQ8pi7poRbappyZ0NaAZIcgngAnNkgvaKYLCgylASboCGCXzua8Vl
XCcUYC6KSErdn+MXzalN8FzT+clpk+25HEp+k9m8CnwPY10dR6LlXxhV20vhWNPQ
uCo4AUhlK3kjWQgMWv2TPRmkk4ZuLAEjh66Cb5jhNQc74bICGn+ni72TAuo88jkJ
J7FQ0KVpphtYx7oV2yWg2hwZRJ4xu3ISHIHm8YO6UY6NCUK3cWWMDk40w0ZjTw6O
PU37/hDIaYDK2IyFkJ4WGbdgVpyWog3eJTwDsp+JuUWFORJQEp+5VMT0WCFYFLTM
PqBCN0F2DAavUcPiIyTEmJg/O1mOaMB/fEjAwNgOrw/tR7ms3Hb0dXCP4r/KMQTc
ZDPr2rXgO+5nFM+zcNYMK8/PQRDff4q+kuMn0q4Ctg/3eRooRSCX9cdnN2H9ceBb
RTo6I9D7Nt/I9M9n9ykJHFix7e4E3YhWZlFmOucl31XAjZ24pmXg1e8pojfznORe
oUURrgL4vLa0uGGZPQrg/moirnlII//ZRCXU7PHG6dulQPz90zBPd5jn59Ofps6w
G4EX0zz5edgq5uQZjeIxS8qaDs/2V1eQ3Ay0C10clzfSeIN/n98nCyOi3Mp3kBJF
ORXt+2FUM7O+WSfofy2Uy7CZUijfCGY0qfDuzy8zbRAoYXcAMuXFR532Yec9NhIB
jRscjgn3EhVaDmci56NsiFbgeX4U1A7Xk8SvpUGFUDe+kqvlKDVd5rpsP4DtAwv7
Ti+HdR4hmjSc2stSZM3xrUvuDl/SfLc4Ov7ELzGpp5HYL5OzQHVVpBwXPIayl4nn
SrCPY/3qun78auTXGcvch71CeTmBgQg8BAWxZBjFhRCJBovMF2RYj6OANBvmvfrZ
0BQHeZOCXvsuanxLHLAf5T3ZQ/tIjd9nYCepg2nYmc1UtpDon289UYcJ0MtXnR4L
R2o5gkRs+i+eybJVA+zlnE8sOCqXfDQLqwkOMOcUMpYutLfp/xS1FOuiSR1V6Vb6
ZioTy9UQ9th312MmfbRVyh8byKLiZjbbv9lMQiPJ1NdhP98Ed7A//rqfXildgN4C
4LakjxVEmnp+9VyyIBOzFKdJFvDfZ4NFW8gMOzLahhbk2wVNT/pLOc9S8ruR61vP
/VfCgONISCDDTGdGJr0mtIps+QI+za+OUb+s4STTl0G1nYh87HPmSpxj1gUBpBJu
4e5MSkkdtLCTjgEnI65p6Rxsb1Y1lAao4jH4cArLlt5ZgDzG3o4/2282nR1O3Pjx
uPBVinXwEFhp4VpPcZYYg9IxdND830B+yKG3v7NS+U0b2YA0eUCH7B5K34eQxrGX
xnFv1331UA9RopD8op2kyf3pGs35u/4/7jwUSI91f4zSHzfCHTPquPcxCto4kmdR
qBh6xvhvpeMJuO565FmgN5WOu2B4JTz/2l22it3kXEPLWfVm+7QnjH10vt6vyz7r
5IXqUjN3KdxAFhcyQbsCIqKNPSI4dFeFdrWfIyN6DvLB2VkfCcCZqZ09Ttm2/fcZ
HHAoolXsg3YOpcRS60u9akgC04RH3RW1PRnZQ1IFRXgvToPcmNAuAXCQiiM29rlF
hXVFYOZHxEOgJQjBDUnoeJDxuj1+KiKy0PUZF1NunX3+oIQqm3Hl7ey9lbMDo+I/
dhubWLABnn5Oxi7YwExymGYfJuhJi4G6pTjaxlS8Jps/JByDPw50szJja/nX09pK
XNJgWYUeC7083C4yRm60CmRdJiti+dt+50f2dET0Q5mr5FqYbH6JjeaTf22ICXN6
HsjUHYrpJVO9NuxCYsEYnV4hJ6MOatmZugmM30HY0o8yV3okNtPuxRMUfJBzWvRV
5tEUVrWsxvGatZjCNqOJLYaa+LRBPnVzSxIBxsp4NZ1VGy3lvWOn8XMI+cnG1jzE
aB9ZggXV1iDrx0muLtFH1RtgClL6jixwunbCZEEK5zx4g92RVdDct3NzMUrJqPzz
RDgY9d9ovvR0yXFUndEqG+byJxYnLhTDY66fsowrU0WWa5OAd9UD7RD77QFacE9o
45Miytb9+kgD2m4CcS7HyTet1hwK+Nk668+rHjinwCeHUrKB8gHc86ER92voJOE6
pWnqM1vSu3xhdywAtTvBDroEdqoMEFmb9hZG9tS/PGX8KqO0dLQyanD927qdBt0x
NtkoqFqjCzWGYl+6jpVPXE+U0/08f3YSvMiN/wOe296g8oJGx4LZp9UjpsJIMb91
QZuOPPzfZmYCszH9MCRaVuGRQJeqaBDBcC/Z6HH41xIoONYEmwtfoae6scaM84ZA
IxgLGtH/Z2zTOCQJiHr+Gkgk1ZBUmUEOwIkbJwWZud4gS94phbf2w8GSQvWF8w+A
9UuKVVYb+YEWC7+9IZMVN4vUFNkUn6qrVsPR1kEp+Rs6KVud5f2d7WWqmc5LoyXA
Fpxvg58KZ3q3QMPa4NE9G6WN3Ja5SJbg0TbrnEQlgtV6/yVcz3bMsn2UlohPbQ1u
sK/U38tXA9Kuf1XaM44bMbP21eLWmcvtBxekaqv/8Q5bsIEFaevU6cDCJIzTmt1X
T2wJIt7HR53kesTw8xzZ+DgYWhNr7iVih84N5KKzRlqn8z+3bgBidkBX97BpQ2hT
Z3aT0DNGVoaXpqPCVDWLmCaSF1QFNGyu8Hnxy2r+2vIIPMtqVKMajFJHfoe3RSPD
7f+7eZZNEnbfGNmtBJBBxzuUbXxoLyEk75ZGMJjvo6JQ4KhXOCgl0YX9aaQJwRX8
p/28D7KKvDc9BOP6xTQHo+LvaPcPt665W3O25VnGUQ0O913MaXzg3IHAgERb2t1W
tHulXax2YpksVAyv74n4LpqMeKHAHDFsptxLptr5i5/nB6txBQ9dzHRTVKgj0rLG
BtjfO/L6O87k6uXQV+5vj/A2kHgdMrpJlff8Jfcf1jl7M/eeSdLzr1oPz+CV6LSh
GfJgYelC0SUuVCgZqW350J6e34rB85wUWwuntVEyKBaTdxznKG9XRbjyYDmbliVS
squzAfz/CllFfW7lfXkbP6tvMlUV12MXWfqsbv5tJTg6bJGXaTo8VlXm1KPTbtrO
dJraplo+LyWUr9sWeamKzItriw2nAQ5MeIpkv5SmSaWdlagFyT36Ym2LyVhnWdRs
LQYZoCPLkWIHQAnicnXKWh4QHF9AIt4Yr8cBYBV+l2VVLqzzMYqULhmlsYswgSQ2
y5XEm6O6FBZxOicGcFaLGnIKOjhz3lAifzn5WfbK3t0W6Tdtst75UmbWCiPvL7/l
gNFkWkuCQGjhF6yzg8WhvcKkCD2rOAIwSahBCqZZKyiiD3q+yeqjCItHkoXH2kO3
OqEg5ViCp5ltc61+P8pyCbdpOYqisuiigvt2XtwpAIZtbu4ajedYcXJzK5urY+Cm
Vxgrs7CY+wa81FdHtatQC/Gj3GTT830Byhd4Euf+KlubWiaeM6Htun92kwXkNnnr
kZxkFCo4bPgsauWK5gvxh/yhcTIcQDr4LFLJtJTkfqCAH0+7tKWApWfAF5/LpbEU
QHDWd4UUGLr33jHPLV+3RdYSOXnxz5rfm5YLqaD2Ze2CMCaOyQPIUZycCkpf2Arg
x6YNq+n3tFgU3FF6AHEvMNJImJW7SVvqW//s8FjtbdYdnHhGWiruoHRD/mP60u21
BkIg72cPSRX24xbJREFnugjQtNnihi7QXM6eTfIimAvxFt6WxUSrCrelZWEE3hzA
JzsLDU5L8jONnSaS0wP/dKFQ0lM0HoGmBm/oRRH4ez1ctarkcZavvk421869g9vc
r2oa/VlD9i8HOZPwv3RvptTD6OQ9IPPqyhbGqNfC8ImkqpskYFg5ah0eyJRKA5lW
uO2BdM3Ptc2Rxd2AayKq6ZgpIrCiYh6Di8FYmw8gMezdANF++iKaVcLR8HroGwty
1ksA6W8EBIZ5BQN9saNp1P8yCKdYBPOrrk2wI+qJAB2Td6iP28wq12Ef+RFdBszw
naIyxcTtcW1umTZCKyVZXHoMVkEL09Ds4SW5jvvsP8C9H6UHP7kZJgZvfthAOeOj
VF83379gXjqmfhXOg0lg8C0TuJ88jduUR9mn62uHVUsDnwaOUyFBcVQ6plEsjfFe
wFKcn6o17hbsU6JDNOkgrruWO80E0gNmeIDmOruy8KqA7i4VrGNuEQ6Ts766f19i
3d+UPBNuUfehxvYR7X+0VMpueZSQr6eEhp2Oo32SAuN2l6JbpJqB6hA7rJmQJKoR
6PuFFS4lyNTcQBbYU828LgsfPWG7oqxD5AXPtz2g6S1BISENlrAXfWfM/xkLvmoh
b/hq+m86mzDUzBpYzwm+Ri6wNGxXayqsu37fycTTaGKHcEOxWME/d4ZDa73C48AD
jTmxE7rYXj9xmUIYLXTJJSW4JQQAXfQslqS9P25KaaBCVWGweC0hNE5jPkgODRWz
oslvQ4N7ije6gSRqb5FfLKhkF0ysvXVf//nv1RwOmOLWx02mdo6sMMJrk7TmGfSq
UzISYbYR8bB80eBgiwDF3KbohLVIKdNCcWbFd7fq8Yfl/GCQUhOy1gpRIqDpGrVv
i59+ar27fgBN0qFZJ+HmTPk080259jXZfvnunmZknIqZSjd2/ODwBuSU+pmAooPE
8rWh4qwrohMp2MtgCpf6bupuFw7E/s+TTAZ4Eqd9/mNkHaBwJ35925x1ABlBGLPZ
Om4uJpiQT2SDsekSncDlKP2hnIOAag9rvPVTXadP6jE3k24ISU2tu4waby0ow9nt
ilpxvn4wYauvJf6FSIhJaZfSD1FKyKrd24ZOWaUDE/0G9ZgfqfDOPw36Na67UWy6
zdyn3h9KZKMfz5pfxwubvb51Aqm0fFzDG7LbC1PiCPHB8rWWe6Z+T22c0QOnOWt9
UR8jocLMlh3EQdooJvQLJXe5UbYp+Yl8EOsdNGrrlM+0Enod/yJUQFQ0r9qGAdxq
OzGuzkya326N2IyDmECEu6VhZeGmQfwyWjt7ZKngXdw4O4UQklRMfN3v1uj3LhaQ
2/URiC2ToC4HcWurhO/hpdo0brKEfIL9oUuJEyq5zZLRpZca/FLiE5X2B5fiSTjt
Lgg+mNrGYNyR9NWYRzrdPLwn2hwy1R+J27iUb5ynSJGw+gT4hl/GTvRUkE0b87GQ
owe5013Fr7veH8Ozl3muf26OC0Mp+rtGeL7Z9aNmE1q8ikLdnJ3NQNmOW8J7lEmu
TIpuBlBjznYvQ7efUm44hS2O32oDg9OXYImk/QRxiniP9u5mUThxzOtv6z3+IWN8
SL3OVMfIz2KmJyxx0g4izcoxwWf5xq3iI915gkGqqqAlM54U0YYoiyp5R86gK06q
rBXO/Gje0HfMiJOV4ThE55/BTTVNIw5UKLq5+sLR1VntKd5TFou0METsQ5b9bZ7O
9glA1jPK8RnZvojqMf3epPpgzwpO4IXKMpzH2+rw1e9u7tgJGSAe+lRz1D7LNoUS
TsFaM/FQE2ck4TijJyuZNyn4JbP02o1y1tP3Jym878QBqohdb2sm+I3ZLuSPOrQv
onqbqL2845juQJwljt+mTIfvLKNoexVSzWvHsq8u5Zjc230gAIYQMO+ZlLpmLpqK
RS6z22qDwdOkrFyrtXZ4b8WicojOcPFei7aMCf9dWFcHZrQkUR7HVVZfumm4nUqA
WPGto6MtaBSgkp5MX2JVTvpqLsq8rv43Y6DlXuzc76plW7gfMJ4lv6Eskcf4I/l1
cUE8qxcnpJoNj9EfvxN4zj7RFdg5jcsSo1ebJ24S8SZm5cf38tvaMfby9bf1uje3
REozNi0WhqocWJW94797qHIhZ4KHi/HaFqeWeMYFqR6dALSOXiSG/RpQC1IAOFdn
hcIxp8QzX27TcWFzpE+1aPq04pM5Io2WKHVt38bMPgMgz1K50NOrdLmoHG2vl4CL
LX0prXM/3/JbCdO4nwXKS2s2GtidiilAWvkpnFcghwm86SqoS/ugIKQQN8aNJZmh
/D/EgzNhcm//XRhw+2zvIeOE6pqaCEYuqoep0Fpah99JNBjolC224TS/wMdDZbY8
qB2tg1QMiREGd5PahlZFncw/DADJugLp6gQPhr7Kqs3bRge5fFZozGufkSPBj8Wp
FPddLGu6HRhS7dsoLYVtgB/2PY+A8es3ovYNEmfOEQDcmkagzbDn9utmZBrFa9Y8
JvM3Cm/6EsjidSnS1b8USQe3okba2nNWZIw6L6NXg7YAoAqc3jEe7MjeIOvaevP9
VWUHIVLq58Ad3V8O4J62mSB5bqEFzE3D19JjYiqm8FZWB+LylR5qS1qxM5eUskBI
KMCK1IbX/q5eEfx2X1Hnhz6Czv6GBIpL7H/McYaMDx38NI1RJ4QFXdcXLWSJUeig
I+w3Mi8a2ZmzsPURjqEwPNtrdTTBG1uqXW3nIcJ5rbOrMfv9jfTTrRjyI538u8Du
yjHeuYhFhKoG/kPsvFV6xq9/llq/CZff6wZU5qDYUO02LEmcPKCADAQgQ1a51ovY
WPj7OcfTmX41Ns4rFjXhFGXZhiFNIjXrFgVhhNkMoxnkOASVC+bBaxeDesijCPZC
ODyaX8sBB2ND+c8mMFkk52j0vUGaukteG1e3/gEz8t3xGIvfcmSG+fWADBFizzUJ
GA66gmLDEFdzHugCkCTqtKSDG1W0N5dSnliXeHRdiB6y7VpPoZ1+DjdUGrIHI6+3
MQaJRTkSV1gJVB0EmbdJaUCMiOG0o5HM9JkyHcezAu3dQW0MnpVu5a9hVHUFEE5h
TrA/9I5EQHTUzbFIyzf1PdFIYc2oUnspwXNNSjsg8TUQhycsW7egAVGO840OJ38S
ks2HYKqXcZBBKshpDivxTirpZy8HJ4Z+uBgjh45z1SWH/UbCGqC7ZYcq/IzGEmr0
dS2IKOKbVwguELRpczrXV5jhag1ChIf0zJWGA8q85tQWCYNrgcMqdcUBFEjS6pbQ
vJR+4vYWShu+lcj3Em4BMY9dirYl+xhGBHZBKMB3QemWV9C7a5xSvDIDk+Bedzj5
aT7CWdhY4KezpXfUbdJysE1Fs42tlTne5tbsRq7VqAtby/ku4Ms75d+aC7slw7b+
QE/lGhDuY4mJDJ65qJT4acNkgPg3ncMNy/kNLV0b1CLTsbnT/IAjVpMvxN8+1zr6
+GihmniVMoz6DO76c3mcFWK77T3j4jBx4fCrtS4nC1FurOoQSLHo6YlczFvLSR00
l+U1i/EuUHPZbHcYtZBG+RiwATLg1zpBDzUaOnLYwU4rOv77djln6J+oWZxsxmn7
FmIUnIjXB1gY4OZeUeXv6AhdUmhILri1ObZmI1K8lghZlexNhx04I7EJvf93QDi6
muCfVZ98qiEALG9OVuYMCnEQTRmJ87TPPvepSY+VxsH8mN0V7bZ6Z7ZkJ2eTslF8
5v18hMFm4NTPuv3R6oud5Iss7widEK3kCNjGN6+sONbZdrXkghLj4TAZnUmE+GmE
l541Ve/3Enxnu9tHf98YbSw76jJpdcPPhDcxIY9txmo2ljAn7wmEvtKtRBe498HS
kOfXERM65IcbdenuyJ659JxPPHxwarYGnLoaOinIdIqJ4a7rcAbGNVUll0iSoCok
x2HZ7XNPT7vlkSdPk3L1lAas77zgPsIGOZ6xnAAww247LWtr9rZigy+HwYzJ65qw
Ozg5tAI6m4GSsgaLUB4CiG76ld6cTOeTsrUVvAOCdLQnov7FInoAipK2N/uCvyFx
wFN+rcZqTrfxFQae/1zXGd8Xk4U8Zzpz++XmlA0l1wx3zvHSeBpfOL+iM0Xfql6n
YZKH/k7chW/C+H3C8emJ9PefwIKymizFAMGKppD/ATbQmNSzREMEmAw92098Aq2B
W/fiATarMp1bGE1igABucxq2z4l4Vw3hXUzdNJFRq04FfH0LadX74thBaQZndwYx
xjkPAFkBWjJpWwitmyl/NVUootALxkJ2bJjCRgYSqC8UI64rE3ZSq6wy7STZ5vO2
KPNj6MDHaD05VgHq7TQd6l1Oxyybp9b8902e9A7t191BB1oQnPSPIHNEPxNfXgfZ
/xN0amc2Cu9gm/jYYY3SYqkO2zSMSZ+kLNQB2+clGtmayExZNO9nBQrGDz7PJxM0
kI3gg10dVrhlb3VP37nKU7PpFu6RQA0N0gaztV3JKfXZABxKzg4XamywUsMMoXYD
ff/homjX9/2GgxmuXkBhd7vdCE71x0G2ZoVk4sKz+Z4eyKG+TMjnXbQ2GfB7+ech
DAxXDQt4Om2FGlvR4hYD4yo3Q8iEq6Q13VDYQaVh9ckzIGXyeJ88A9LW/6qgJFng
8pYRI2ix5Lcd8RuPYPwX2jhLsFKLSQKMgZUVVxcZdiOToraG+x+9nFzhncxqu07p
lnBJMEDEgXJga4y9VoHCSDJIX+eg2m7Ged3TiSCPigPXmeU9FHkqIk9yo2kNlJbf
PlHIOX7sx8wfou2CQEpycTlxT7INLqP71NwykxPeZQ199SCSV+kqs6gAbCr+rJ5p
J8SD1KcJoLNB7MZ6l3iSSF5sWWVDfjGe1QOHedECebMGiAHsSWg/EM9Vgw6HSFSQ
bErCGkO10epA/ieWvJj3LBDEijQrlBmJLIfgghaTNscSufjMqpO3iQhA4kAqTI8e
C1UonqBsws1QEeKWGBiuT+4DfeWd3WY53quW7IfNXHeMj5y3jJen9K2k+qCvywqE
9f5eebSz4y7O+RoybpFtosVzV8tI84P6k6sF5DWf47XLZb0bXpwKUj78hYKbf8jc
qtRlVGp3V/NjW4bpiDYcVK3ooiceI/xbTnDRg5LDhOX3+39ydnsyTWdqvoavDWkR
Vk9xlPSlO8dfZ/JTBcClQx2iIjZ2XNWN5V5869SMsuGhsD+EV6NglbMTfSlBT0UI
/a5iEevFsxd6EYNfWczFaoLKY0qvCI9pm6BVDo+Y9RncuAaxlIkS9uBbYgT8zN6t
VN9+G2BrGv/qmEPdp4rW+W5mRvVLSb4JE5Wxwp2g4lXDsv39tErPitXBMu2USOQs
vQje03tDNzQ720/8NSgBWTc2omcKbUkxYoY8I5ZIoh0mD+zovJW1/lccAZNjtLzg
obTU8U+MfRJSqdPADpjcszF/zGTjmU6tvn/Rb7d8X7PrQ72U9aRbkrAA2KA4epJa
Bm9JqnJ13VYlc6GsFpPk/sGxfdmf22Jn8BEF5218M7aLgK7qEy4zItj8dU0yYCLB
HY+NnonHHPZmU5sY4ako+wQmyvX0RyOlHBABLwO8/llB0J6dmnHWI6n3x6qqDW0/
jOBK4U0qhZaLPXfuI+GQnSJcT1+EK44/5Y6GU0sYrSQzfkwJdmoagU0TeC2SWHSK
pOxkvxTNU5Jwefszk/mxJ39YXBOdnZU8QCVAAlEibjMlgZIh7hhpG/jrxwaTxrcN
JKtNYVkSQA9aV0yUP40x845iwiN7ZDwYbs7GNqgwXWN6kyXxEBKLzyXWdlzjY5s2
pSeBzV/cSEd/BkML0i3dMF3NTG/YsYV963iwc30x2gps0mLMkIaHJ33y+dYhWfxs
CITAM3YDo5h1PsTEkWAmctevnAylT7AJjZ6t6+IiNAi9lYqPuhsczz7og3tjAIjN
GiAL7XkyKr5OM3lz0w8Dje8EjOgrDn/xxhALZTghceXOF9BFTohYDNytkKZdvjlh
URMT8Qp9VLRkmtAqqnNJ1UeRj6nKiF/QgeVYPD9pM7mTssz45M9GU4OdacpjL3Y0
57vU5j1Glr9xnFRHI/14kDOIQmjKcBT/6mcoaWvzy2m5dYQYG1PCC+VXMu/vAjw9
lZ7rynJodh8i2BhrJuZye0mFV9pHrtEJUouj3cUCALQGagUAyIDyXn6Q04U+6Vz4
Uw0quRwx0W+8ZoLk1Ds5opp+xpqGVZaGFROpGdSzPTQ5i8bA9HU93dl7oEEgX2AO
yuFMxSXq/XBdy66uiZSOoZi2CfoQXMjXH5vX8oRFQzq6TlwnLIkqSy3WOoRYj9Hl
Fj33pCembrxwJYpQcwqcxsg4JGWWglOOXwg+KJ9YYR0OLlr/r4VKHW3BZ6EzRW/P
iF2ZBqPkfcenwgt2kG7i8YZvITMFkHV+23A/8d9AAgZ2R3FPX1mhFEtx2WkUY9OI
aTROgINyFdVVxln/5E/9G6RJBEz8dJ/9O6SBfX6O6Lt1DCGdjIh3wwDhMbgknghh
Zio5msOFceReqwUumQdIl4TF2OdE5ubURvt15NWuH9XOLnCJOV5a0dXxi2YEbmeh
/syTzoJNE2td9jPUwpGpBUUXFzD6JIGPbBu4bel4F5RcVSAwnWaO/r3qidsXVb05
Mmb2R+8K6om7gI081Xh4yH5PL8G1nt6EUOwf4kNABOFtuncl0+Uvx+k67LOXObfG
EuMf1L2GoYhs0bJlmYRVJFl3ErS4DWG9OZUVPNtAtnmB+SxktqmHUJ8c94vfTJXt
vEosSyPJPRDfuIH9vAampOZUUIP8zY4cUYWLEk7ZhFotVPRTc54MCMEfO0fPo7Rp
mfC82bBWCnBkptlJ+u/54n8uz5+coXtHzc602Ukbeq14SgZetb4C9HgYNr+pfMQv
pFYllsryiCPxC2YVfQXBwaqXYUOzAX3J0SaHd/RtX4j9Bed+xNORX/G2IGfAvT4L
peGrabiqCGS/0BMXruSGqs5KhkE6W39WNwCGVRK2Zom5FbT49N4lElIeYFsfVDiw
yHJEe0MwT8hYEQX2TEVPMbSDN6YbKt7pkrYobtSpkBzwcIybQdkTMQRZAIwoAzR1
llI9xlj21KPaMtPrczPjeGYydeeUTBbcz/kXx3KmFQ4RrToSIHzYPSJMB8CUaEOM
2p3kFBB8Ta9bfFq3MHoyCadoqBp1ET4Q2gJ7qpX1U3swUyC2Pu3dWc+1FnrrtL0z
5GE/mNJlSTFyYvWIkiM/O1QE46qYRIpdNTyow1vsx9K9OaJAIy8Ymu83OH6EBf7V
WhNzrKJZfwM7OK7ZLm4O/tgkHgm72SSnPQBZ1MvAGHhkImpufkKOkgHy2m1EyWWy
7s4cT+vHUqLx5lTWBH+yGTlBfBmQ4b80BWXsbyCxh39JxU60zcdKqR/gEXO2sC1z
WqkVEFtUenXRbsq8n0a19YyfcLEGHpCsYz0Kvt3VY5+NnDGCLpoOdHlT3J7yiJ2C
RQk3HsqGxEmscPExqfTxN6/B1bh0eH2zIJRXOeXsMR7gJpQdbQx5wMWC2+FlqHwT
hvrLZhqyz8hNGkx3JNuTP+tZDy1eZcdIzr4s9z/8poiFd+0UhHbl0fPGP7Yn2A6r
n1DRakZ2nIUrTrJWlXx6DS6r1fRDgDHu74gqYqvWffx4deMcWXn6INoaPn5+20Cl
ziR3j5sOo3Jn0QL50hKxRcsFzOQA/61mLO9zC9h0UkCVSt1lwn3iTBaUixLfVWvd
mXrieFZUEIgZc9DoHlnRczW4A0WryPaAaWS7to2zUjhOxB9/H00sF4oA8/FzCohd
3+rCiBMlYfZ99okj3BZbWpVFppRSEshg65LF6IafkHaSicTtRS6Ee6EEhTJlTH65
dlEOqHZsNCBhdG/yRG4jUGpeoCy7CaxzuuNqvB3DHrTYzhZ0mAX5Q3mFjypDfoPn
QXFoJ8iv80NzbTAzKVGIZDcWuuQnHQXLQccqi05YsizEKHRNJzDbkcLJ1dzggxmV
jDQxhlG0wWZ++HysVcGtL6Ea/tbBuAE/VLAHFe0QrEO4IbMNbaVi/xpdQvRAvLxa
a0Vx+xmOdWZfWECM+JehbzGmxl6ZoyKeoHgR0+7zYGFPcSsksnHVq6nVhPS0lPf8
vF7Jr5xRGHCS0kaSwmVhsjHPF9JzmwWK/jnHNL+vJ+3XAG1cUqqRcs01Gz8oL+cV
bBcPGyX504ovD5fFR49gVVDvyW+4l8cSNdC5mgbYTFc74fLDuVHpqfTh5qJYe3h6
wM12z/XOpvCPdvzg0kyrvLWHOrLivN/KC/2afSwrzYtPu/kndsmq1iDPD3D9Iy8E
JCUWswFotUqCz2mNHZ0shMiuw2JMF3UpQwIJ5vh+FH5xgTk27w/LDk9Z7Y4xrvRH
GMrXwfaGuQWwPM+F3eaBS0bsSu93+Bx5taEA15yJDog94WytJn8SadYWo6CY9DPg
BxXuE4QTUaijiBYPkCipjlyXq5HkiS5kXgWhxWh+iD7636XHDVBifUXMASeh9K4G
VrnlWa3eAPliDb1mReTu3WYzlLaP4SSEqylrBwALEdu/vUXpfqnBepj94hblOMJA
FzNDwVjlAlhBDvVDxRCu1FjQiV6/E2cK7ABO5Ht6vqIXW/HZdWU6IQMSyOvTbzrT
L2B3+YJlbeFQmF1wPs3Dskno0Kz7Gl3I/GORAMDlwjQBPXT3CCxI3Pyk5aGMSPa4
zqrRuArZ0NHy04DCpkmP/bz8gTz4rYyMtCLqqyB5LuPD7/D03IoBF6culDlgwxjw
iG08jrbxd0FmIqUwkwEAOaOCW50BQowUwfaNCExJzOaLZDa9SHs65l4EcW149zWt
0p3jcz/e0PqCHOUllu35HxArI2+2qhhkJ+YGzf9Fyare9QRXgjgcraPAJ4f5S4bx
KZbxSihZu7c7vILLAZZJP08QEEctsr+wCq8EA27EqCd+0wNYRdyq65nHmW5bHU5v
akjlczUDBrx1iNRzZ7JaWc46+Rk5GvLUN37louKNhfMGRa1QGLhdamYUe6ED4mJ2
jrtKAhY03hzixwzyyHkGMZ+jJDKZq7x/B7WN8qF8X+l3so7g9oyW1NSDHspQ4Z8f
V5xq1c4m7YNHW4SVoryWl0ZlK+hqxUmEiGHCMjFq7qQLV/Q8SluoTMwlCPrOHtoT
8UcR5jxEhFBdvA84NdOek62XEuIshPtafgRRXZSjT7fN0EbzQtxvWrX1QjnF3mc7
uZZLCW/I7QvGi6Muf6L6FR0r8KZ3DpAs8EJa1x8/PTT7RMqAzznWgSL3AWaLU3df
tvUBWBFRx8B1+9O5r/7KJi3FaNNmu8/chTxSOLlc3DqVWmdZwW8rodw01vKOd3X1
fgrEAH8uapusx0bsaQ8Ea5vgQK1Tcb9XbhDrgRu97yVVjCKE2KDYYCB2SBm9PkVc
2y9M+aVbCuMC9pl2ynINRJJ51ShHEPCpRZWRKM8OCY+lYk9fLA9yZHKrZUiii5gD
B2QMciLVX8mwV/eXFGEjvuYv4632uW4iawDEmE4CSFg07Zp+lQXUVcnRosh1ai0p
ATgAzvXh805H3mrZYpK1aOcA9DQT/v1cUWZ5S++ceQLphZz962b+sHkbWKja8DXz
HZ0m5eCYUyrMVdWZGZqkM2YNcoUjNQR1/mKag47H9564V4qWLeV0ydOBAn5RPq6N
FWdykSfrrpHCZ/b2nJI8F5aIL69wz7nQHOHhVVQaDjg/wxqHhGouVUp3ny3ksIL9
nCEFh1ieIROI5bD2cQsi70zCCBqjnbBzcQu9K1BpbrjUGPXR89BdDwqYclvmmuNl
KLSxU0ONp0aJRwNITeFLqot5/rcRxRUCeZH2tyDUjwVXqBh+ae0mDMSqOokd0yt/
Wt8Irhoh2E6DSkgY+xTeX8G0nzxTXLrvZfVtL86pSBvkg9vv5ddzXTrJ4TAWmRh+
uMou15cdKsbhLsYsY8tl6L31ii1NC7NHqsVkdkeio1rwO4JwgB+6YXIeH9wRwPJF
YAdvmUYDymosDbDbL7xPRwTlgWYDAabG+SfYHcCg5+xK3S416W3HFctNpXArz0ta
vAGl5Z22fMQdalPR/EEj99LjJfSnXLFa2GBuOZGG4yCxLy5CgBsQ7dbv/U9az1zP
i/w1F0nr1Hc/O9CtbJkbjdIp7+9ram3i7g8LmO+GB3ojhzskBnqKHMQKJ3suXWc4
fL6cOa4t0c5xGcHo+sGPHILhVs/3hObDG2Q6OXULwjX3GdssLvVXr1oXclUnWgn2
4nwIQfo5jVyukUzJPFLBXYmYZGQZoquM9yALccC2aY06HNoaWNKq2UMo+7OPaVyQ
YjF5AMXvTlU5zMwazyM8mPgjoVuGeGVgdJznHXlqsjC6QWSt41h1XdGt1NMcPBd6
kD2QZGGWWYUIcHWMXtzybzw0vzjMSky6JVebA3Ou7T+XuuWYYaaX0rsnrgLsZhlK
MZOLOt3gkcf1UCbWZgO72hjXJ8QbIi3yt5b1joRRbpkesdI3Dw4m/YgfnNJ6Ac0/
rD5kHyAiubiI0CfmVf/BGHGqjlFb+ycekMmlPo4UgI0yntM4vifcv4KEH34H9j4H
meruyA3KPykBXtQk2N9mFcWikLTyz6S8pQ7Z+GmFzSj/pxQ819JrYFrpdBPqX14D
xytrvBwOZbtDu1oEZOrBS5MRiZRSk9b+8JW3U6wLVCXwyQkxJADV5byzStE+yojE
ESAFjm5C3mAGb63WuYScM8jDEVcl9hnsWyNO5kDI0e1aGFDnKnj8rcq5p1ILbTVv
H7MFUOlob3oSN+2rOCKIjIXpyE7S5gSJY9vcE5TnhJOaaH8r7wFw3Ob9sWDhS/z7
UUaM7eWi2mjWgDno8MWZEyxNnTBQCF3IW6FjOVKBGTCmWHITuUf1n6yC8khSOfLe
PwSkk3kpcT9D4g4BuNuToLfidPhycMPuY3Fsefn6jPcnMQ7+UtnP+XXfCc968N8G
nldhUuyEUm1/dK/5o8hHw+zHCKXc0u/qkdF55fHgXv+HbyqlEltmdDBh3ptZpQLc
UNJYah1L3YGEpVJAgCvRkVL1QwEnQZMYQVkBEcpDahINh2eV0rJpl/++rKquj20Y
8SocNd1tdssOPwQB7DWTFQzWKMXn2rk25Hgqu3wgcu5/pmZ1uNu3ndz/rD6HCRuh
jYvIgUQWNI5AYncR1/IqvA4/ulNBacRNRVyaDW0kuxrcuTFxIsd5ZsNrOhzqjQ7D
apGiNGP4WlxsUyjp3BfsJRh6UQChMCADoolpK7LMjvIiDYOyreXZTEnoeih+/oHA
eT5zgCvtBUI2R6gnLcxOVpjtB0IFsfE4m52QE3GAZvqfPiw90sQLuLncek5d26Yh
kOrB9RUllFJuiXQixxJLD5UEI70J87g10ssZoU3nn00ozvIFTen+4/E5DRrKoAVE
2gmIf8TjARuHu1H6wqDWt73HsXzxbZTMGnTfU/jTTaxOC8atU0CN9X0yG/gpmT+B
f5YVAzus+mzfIc9MjAiG7gn8k3ZnAbWLpS4JZkps3HeD0meWR/qOjqGNuUkSoq3q
07pbHE56oLjsysNrMlGvlK8mmEE5rlCFuCCH39RpIDsnbVt3LL71hcTqW43TS+bA
BhmqNWIUSRosqon3/mJuS+TIwWhkDzz/6f81RyEdEh3rmhb1MP9AfYctSgwdK07l
REQmYcaLYBIkGipDroPWjBj3lK8QRjOmXqqWlIT6twhjE2eFmsQhoXHwKUt+BQD6
zuI8Lg++9McJ8jVvWj0j5MhwmeYoeMexCweNzV98k2VsYTfp4wl0OBL6dCMlzQv1
Q46cr5R4tDN1SxXY8dNzhdwOjSsvKiunvlZIMggvNRP6a+Ci9GcuDM8hIOP+IQY1
RMPnz3SCfPo9LgunHX5V1XN0ddDr/TGvsJmzHj3Tdr5ISzKGR1GpawNB2WEe4Xeu
Oo93F/lN4Osvixna/qEApnUnOfv7Nk+rF8T6d3jtkVTleCQYeS66ZQC8soi/pwvn
7FjY7zMTpf8ZqjsPn6UZlxruOCx9HstR+XzUZum3JwP7hCGZWRFNDlJdnBYPwPLx
8uZB80rzrO8RLN2GLj/s8UZmbi7H6Oa0vYuXBfNYQD2MtPv1ijZgJfXiIUCMhKQ0
zA2r6Byk35Eab09P5sddvHZjkplidFbFmtgn1OT00mm0OmC/2WVcFM5hHf5Zy3O2
saaMhVw43OinrvT5tSugzosTmX6Njmf64JaboTy1150/bb6yWO6Y1JW2FdIT1UoE
upTfd0V68cXJQCCfkkm9RzaEWwP//ZiBu6gPZicc1badiwfXT8Qshflezd6/0cxu
B+0DKir8cCNBu8W0uin1Ag3p92dNFlzUZ8upphJKmgJzP1FNpJxZ1jgdF2g3pu91
4eSkfUb98j4PGZLEC1J2n8sh634QHIpn8GXGUcGYXWT4Msgz+//Rm0ONwYPHRGZu
LUElSTBaSD8Nx8ILUdNQC1aVMd3R8WFFlivKCjy0/ZFnOooqppT0g2oT3dJ+l0eq
nKrAj3wuvwtqYacUjVsW/U7EE6ItoDgju7gYadnF0LL9yJBH2N6ab2zWixP3tXTt
+5J4f3+5F/0nS6QLtzmFbvI5/Ro2wSQlLXWbXHpvuZcHK65QnRgNgIFsBO4Vb0/K
4l6DxZXJNJ+3tpfFnsev4Dp2o69STCRktKnZoBemFc6l6ogLx2X21CXi7EYi6zs2
HUW7AuoDuV1aFuuq4gYgTH/JiLAiffS2b0DL2qUODAwZVhffNW0EIR/LmtInyq/Y
dgxWlsB7p5DQnRuo4SKTTyBdsIo0vRF7L3eFxrvRPRu6uMSKZnalrcOrTQ5h9z3A
pjf8jYMB9/NFuYBJDFsDdRiiIgaMwj3i2TPQhiO5tDfSDNKTVgT2X/H6QG3CnIA1
xhmsZsj83fO4VWpo3yJnXUkb02QDnqtLjKQ/jqaVzpdJ5cWDzLh/pAA5CFy3UsCs
dYJuGz/t/e8Nrb2xvrS7e003p1vXLZqjcVSwpopMnWqGR/3MQdgRaiebbRyzDfwo
9K+CG4fERPaduI4TR9yQ2ciL4x9kOsN4Jq5HZukvlltxwcD0UltaWzm1Z7DE5QxJ
CY1SuaKrfOwPkz1yYU836dJDwF/0Q71g8ix6mstK9HgLtWYMQqRoa3ed4gW5Fi14
j13PogPgLNJLNSnWcloz0Fvmx9ib6ZxNGc3wuNuoa69Qr9xRUACJNKgjK5isFF93
HIJCb325nYR5FOk/hwHJy/7M4mn1RQCvtyvyWrODJKX0k/74nUF90b1hpUqaBOAb
bkLB684ZlHLgWvQ0n5X8xXFGb30Skf7qMb88rfGhnWSqeW6EJEyiOiucrMULBG8x
2nzw7CwgLit5U6E46J3QH9/vMIAIZbjZYJibHmH4C+B3dQaTLLWBJvgc2Aukp07d
KVvjQUyO9SKHwfIQ2+LemcGwYNvp1CCBmW19IFPa5X8NhXfwVZxMiU0ZYltgbbjU
x00YxP0SpFdnQmU0R6xvTeEEmGN8gcjg2GD0on8TBRtu9D8sxQu0AL9NsDoBnlYN
0f/kk9rWr2y0NWKkzt7i/1iaj6/Xqut+aQw75JZhid9Ezi7BiYW12NeVCWR1MaOh
GsvGnMl9Owv/0CXiUCTzFvCW2+FSVQQMOwpu4CIOP/tbmxw6yY7CmTX4arwNtA3O
XIB9i3qfdVpUa/daUWmfiOoshEUzKS2nHLM1aKkcYjuueEU7r9SOfK9TnC2xW/3s
ZRKkCRk2+dUualuwNaYgAhd7peK6FDJwznyzRM5/16Wrhowky7A70jALtU3wZFf1
8hTTOq78aFTJpOkETXogQ+BHbaySacXst1RUarpbhdRQUUctvZJj8ruk7EPByBe8
UwAqKe8lULukpRx1CYQIjv1Q3Dprz7DnJYa9r+ZBkoze4d+gZSvemDe5TPW5dOb+
J8mZgdoDOzZqGWQgacgvXg7o7wD873FIagE1l0Z/ITRiZ7lKrvN2DQ9QtjB3qPe7
e+l2olnaZHDIcppr7lvXcfj2flPFPYSL4Adci8Vuaed9h5rjeG1T4fY7QC3ZJd7m
a/oSZxb9cvVGCSVfaeBe6SVPHD5NCB2DbFZQyKbBEHyd3uM1ejCRK8Q/1mtd9Fcz
P4lspyrNZ1lIa8piOtzj/GRuvduUnToC+10alfJFiqTwmxK0kG/Zwc2jENqI0QIY
w1qtHs6vx73/VMX9wFqdHrx8kweoMzAk6EErIxPQ3Woen6uh7huBq/ZOoNVdrtNv
sLShma+EnU+Xnldlg6XQTU5nTkctAJneW+NaZ87x3pkMtPzwNxHVTo6hBh1J2l/O
UI5JubQJj5msRlNx0Zrhx+hMXX+vzY9nfHXMe7pb0vpDp60gZnNHyqimRxxyau7U
Ywy+94WX3uQpOI1Id6tfXUeUi4IBjh9OWyVH+mzmhIpbNCdOn5a799k+QpsZ2TxJ
7ME7rgMn/gjFn+ZkOBJEdbH16xv06ntyhKrS7kc7g2uzWquIqRZy5LgqNGV14b1Y
khFJvoSbPH4aWi3P6jutooX7alCTYlzEM0n0yw6Do39ETZr4P2MmT+gKKbxzUPIo
e/iewSgFjY6EPa87tDp2jdDkALt+WX5lISioVmWpfu6j9px5XbIr2giGXsALUVfA
yqiuA89E2JBxfNqGG23/l2Sg/kkjoyyKaC1JrbA9XlfSu1/FhrsoHwce0nJvRMdI
FlVNzrnuiyolvdE+IMPFgcV7KmpYCwSsz6u8DLvCtamBw+tYWOdxG4AEkINRNJBA
C4z7WyoWSvgxiTSjFnSviaN+j66iBN+fzNPOhHN1vr82CrGwP6VGPEpANP2TEMri
1GselXph/xLczvDrD/6iTaJBliDlCQvYfSk2LeyUStMT0IFwiek1Ckp5DJT9qt3+
yux2zTk6ZhwQtM8F9/2ko5lc3IW+9W9PWSTZ5guJoDifs3Q1/bl++HJQ0VWZVznU
6I7KmfORfO8cDBG+Ss54RkVF6Hmqa3V/zKbsm3GukGboFy425hVJgtVO3u50ZFto
V48eCWr1BU9g7VEEAQBNIIAok36XbDBDeeycRfpoHqZFawMFSbEVYgtozPbQT6oF
Tz8Ec/5DHq6z+C5RMOjxFPW/5yfdgzEDBiP11IQvE4asvY1UwuwmGwSYmJ8TXZz4
HfsAnCJRT49RjxQ+zLcZtParV6Iiiz7gDk9Gij3OiWLgqwuAV7aM7xKk2f1GXpO9
gKDiA2sP/5HIoltvxgLBfcOA31U38d+kiIyERs8fgFDQdut/xvzHym6d2s09jx8+
PsL4r0HbUUukOQgVSmkIkGlmVILcZyyuLn2FfqudoWIp147/TUoLtD5N6pxiwt5x
3AZuiVpSuMEEjk9QtvgW18QxkUXP9uYQ/NUT1CMeo/VK9ZLm0CxpJfn2stJslEKq
5Hz1U3NApoa2bZ7xTU0OU2wchnFHnyaRDXiHuY6ClvIGdZ2sxp8kWTC+veJQsP9w
BUeTKu4yaR/fxFiLyCRGPRvphwzNe+1x4UxfOyqOQun5nYAGyNv6PQPZl0XZCm+r
Ej1VQfouIXqUVNPO5hqePaPUYru6sxWaZUws/gALWBNCKOfE02R9m9fitMvgRMjq
c8PqnE5a4jKtCHuq/TR5zzlI/QVhfJFSHtJe6szgZEN4zxluQzzS7Rlq7PlffMms
/96upx4UhwxZrFy+EZs2L0g+3YJUisn7k52ESgWa6cDEAiG8Y4xKimHWF6+FgBtt
dTiFcLlx/0MC8byIUHXO7DygWsqeyEO2rpuXqBFLMMR+s5etRdY3dyFeMrk7V2qg
xTsg1q7AnKCILBEL2nnLs5D3pZcUgKOjx83s8CcE5I3GJMs4ZhCuKTmYevygaQy3
ULaekdeQj/PCPGCIuK1kCVFdvtV6ujN4WhA/lye8UoheVWzKrZK95cXfSQ4lXZRg
g/EyCoqqhBrE4a3Z9FLfgdXxb5XebqieUBR/2vMDNMMMzCwsj/lH7s/DAdAyzLfC
jgTI23VovF7fZWO15kbzvK69hkA9xCvr+QvN4gB1jMrG+LNUBOufCIJPUwBEnmDG
3egfEW/jey3PNXYhNnwCIeFcYO3iznnL0mmdNW4WDXT1ikDx6aXpFtaf9ur7ECNn
G6haajvI6XU0qhOQfcbhvv9UoEy21CDDuJ+kxUDK1stja/lWKeJv/df8FTQtCTJE
+S5ckMmoJ6bn7pi05+Vx69/FsLKymTgVCtARK3I046RgsGtJkzv6WuXGszJFWdbH
cikyaUkfK3eJ2B/5sQC9zu2bbXzJs6usLzOZ7txu/OlqYpDTp7Y0Pz9J5QtPWVkJ
wiO6e9jAdD3xFKFffttI4CrhpnJC3tVLvfuBTkelOx39QN4+c3wnI9UPQj3JVbGz
JWwD4ICZmKRxRtTxSwEAGIzbi46UfiYWDWt/k6HQIwC3z/DIlFtUWRwwL/jywukk
kMb4mlvdBCeCUJsFSZDwQW6CLL3KFcClk4NdbeH1pMIiQc5bQO905LNEm2hwPYcZ
SYx5CtACErL4T508x01FKrHdghvf/bBrIes9xs8aVlnYP+YCqOVf1LglbwTZB2J0
m7snLE3sd7wRhpx6d2BQa3wd8hgo1CtUSgYV4OTPk8IRA6y6HeR3KydTZKKdFSGV
A2uvOqpHvkKvhGai2j/VPOweZi4dVo4jWdBmy6aYylWKag0fd/uR841PABAT6wCH
T1aPPU7OoozGJVtMekKfBqlYGdhnumQz+kgsuHyDriqkyqou4aZSKoRciFnwV89q
gfV+NONkc6TyMwtRFgeNUMVbWrVywk5zNLXCCPN3MDBQp3KNiGwl7xmJUBARNLUY
CUG/LomdRY5cNKp7ao+QBIqjsG8I2MOzpN0hPzJ4DcFNZus1+iLvDK+c2R1uMkPq
SdlSs1EjBQWJYfkGsZMmhVyKrsxDi5Y2kPeViUB/JyxUEhZocmGh2FWxU6MBg0ne
Yh/iDSXpwYqsCmQRb9EP6RY/tEPz7Dz3+MCFgAcS5y3NM6aUD/8kyOb6npXnDogu
BgJ/GUuFF1TxrD76F21ZqFN+7xx42l9vLBeSGcXnTDPvsGoVZy663MXKplPwdSiV
D8+OZeWuCC1Rhn9cjUcS2lTL7/gSl0u71808xcyGXuTwbzV4g+/SzG9hHhgEPgWn
eNb85y1qk3KLVJaQCAG6E1HhYS6WWkTBtjzmyitwiU8K44PDorh0Zx67C5taWqKw
BgDMDFidRKoZzTcMAPCe5IsGzBzJnHA7vbEblo1qQWpAkTN7oPhadiORFQU++U2q
Mtek7ghETZlevi+33QoT64QhtUBw/gwYQDKjZI2+dQuSszdOyhGXEOV+f2vCyx2U
rHgq3ewwbjk8z/BBfYBXftY0k0OUX+6mtnJHyo8180LMnxR0CRDcRMQnrvFz5MNZ
SB3s6M+SEPgt57l470OBwpfWLJJqU+MbPD+qvLXixk10oY/7jcdyz4Tolocbg4Ov
fDNiTK3YdcLfYHkGbJyXtLDBj/bJSn5LsLg4D/4V6sGucta5zL9CJ6lTf626cXon
penlSXYUu0L1BVSRYtdGn321so5b6MCbN6+0ZZ0EInKqmMJ6YNdWX6s7b9wbNTw+
ppTOscgKhnhTK32MsKYkYq2SKXeKHFYwUUg0h2ukZVUdeVRyDimDas9VbffGCGLC
Wzo7DLCO42L+C4b5namw0iUwHW7T5VZfZTcSAcsr0VUwN2FuhRo7qV+IqTg00o0K
Zh+oWiepfxuffxBJpaqOHFzCCcm9LQoS6jZkm+5TwpfmYRbLE7cHNVZusC93WnsN
nE5q2wUKv3Fqs4id/8XT0mRPKIRSYbtSlc50FW7St6oCBnrbPnF7ihr/guuPw4WU
gJfs42ynSqEg/nTdgBJNK6/FAkKeqxOvq93K9ON38puztlGGKw/NtHin2OTHHBCN
YGwR0iFDghTxfZGV4HTc65Wr+3tvqye+/1pCLDeigXOgryO0HY08y7p4elxSu9h4
tciX79h4eGMeQJjbV+KkOUr5X5hLY1FDvELZyM4YqhxktD/uvkOSlDCK1R46CAQz
ASP7825ssuLpw57UdZlfUXe92vQQ5Vt0bgsGDbIJWnweiyIkm05qpOWyi371c+v7
ttQGVId39yEwcJ/3fbubSTyRkT4Q2T2PVbqXekuhhOZGaMYTJ2v5iTIAann8zqdw
WTGCwU+LvdQG0DF7rIp6Tdqros3oMXb4tscbo6awUEEvsP0pB20xu0TL8z0T8cfy
BrCCgyDMPXVyrCLvsNCdce9eQxdkz490a0JEu+sZqdMgqQuYusIxjNRHODbmhB7G
zH7l0VfP3aUFNz6QCTjPUX3fHjGzRFXMTxbIWRaKjwz6QozT7ouZdwrFR94xCm7n
DwVLnPtmn1p2mCFVa9kJugZyELb762xeA5i/1H5LkVx/Cjq9kRX6R+PZyq4N+qs+
lVLNj7AWk/G+TneFXUknQBDHdWEEjDpQLi4E5p/efyl48XC3xqjnzG+kWoeLXbgQ
HXHnPskiWnCbZU6K6vduqbYz2/k/JYrDZ7pV+FHr3TTF4foSuZYWBJeWBRvYe4yq
KC9O4LBP2mYQliajWx1mu15Ho8GjU5DruG9nIR5BFD+74G218CadEhdKfkxz+TFM
3uN5riLPeHVuSAxBB6sVOzmL03BAXY72EeGhSTRlRmot9vsuOZjhzcawtYgQit5M
LfCHkOFNxA8EcKhtFaDfuRRC3hsPxvUKXrAhrAf08jo/9UxMi0MB/0n3dihI1fPl
7KAujUM2yZkx71x4GKFLUOk7+bI9TxREUG+pl8gOttxitmQUK0+lbni1VSOqDwqU
CkCaKir+ZutGWBxN+aZiDXGP6CjW6f/gSw7FfR8muLD/LirN0h7SMCFCdYkSwW8p
IOKqDqYlJnkPCa7O3CqOugsgv8JEILLcrHkS1GtQyCo3QA98bpoZF/CAzl7IIs2z
w9fLqCvGafw903ei1bDNNuUJKb2x2zhbSBnP6yo/d4xSjxUdKuQNDTjaFZdxbbtz
YMYppPSArRwN7C25WxnQ2/0Fjk1yM9WdeZ2QLOMiEZE/D79xyvGXVPGc8FB85Bkh
dOyRKIZPI0Fw7fRbBn+I9hcGkT8exMGe7nyje8fP8WKi8rLAKegH1G+Gni5wdmvt
ChwxtRPTd3BtVd7U1+BNAYb9J8qa3IqoszNP1CAQgr+ORY2Mc3hPH1/tmiEUga96
hLvxYcEy1DhSFJ/CdP5w5jZpweCNyGFhUufnx3Gis/l3QaTM/ojeb1riKjHlEk+j
VywAV6/0mE2y3IqyBzcV6NwGbLjAieggFohHIcrQgOVJnISpikN6U9JGtHSyVbPj
yG55jy0Nna/hW/Ycn3ZRt5Ru7NgPpXn5f6RS1nTNvqnkRqMqUlNp3kvwEyvdDsdw
peZ1df7xrcNgY+NVrXYbYq0bdenpC9kC29tiQTuOGclFC9/ZWmq/Rwv4d7kbnvAN
m25hE8bo+FiCF7vdmG46D5PkPVoLCquLY5NWZ0ShkWXgJsJY+MNRKsWDYTPh6SDR
44e1JCMm375iOqsasGG0r7yuHdfMQvoQLSpaHHNv02dAkznba2hOzkS18dHUGzpR
nmO1PqiPNePeQZLoDaTM+QXlITJiaaw1dJUt52G6kOMiQpJ+kT8OuazGgzbg4ZkO
tK4YGQydV5PelhUCyGcQs7CVnHXHFN6LnfI3eCTzJP0YtlighHyNcGlAjJM3DdK9
PNMbdSnJ8o1DDKFCAUs+ASe22ubevucwGAtHzPsBvrbj73JyIDLypa/IpM6wB9FV
zCCBXAWi+rQ8qfv/p02lT/snzT6a91/Vta4vsjL8Aj6dhgGNkyS2mXX6zKsL6HKg
KPLaT5y+5iM4/caSslhc72193e7SMV67ZBN2nm4msAg74dsXAaaswgWCLwsMBLEU
pQJOLzbKIfPg+YKZyspHg9q0HEXinR/7Urg/PVI/42+bG5dY10dnQeXig6/Sr57k
ySHGNRENT9z4hriH/c3OzMR5P3BDKJ8ZQODaZxhl4TT5T2VU+1qP7iUfA/+kMbP6
iDUjjsOOUInOyMAxC0ptsKouMIYyLnvxcCOuA+ASJpgwrfxsn912yeuuPBO6Q6qD
hTyEZ801nqmC+L5eV0sCEsIAotmzhMowfvQZmWHN+pCB9ziayvyt1NyUWxkRQA4P
Od+MpZrhrJpCi2Qkrvu/OqhIAbkZjKrtcesuW2hHQ9NrA/siYwORXXoOdrvD5XQl
MuQRRD/LdsEKtLuxesbhOL1ZbQJQGr0SlXpIpJ2IqRHhXrhLRQuAwjPjKa5TRc3E
TKfyXUdQozv7t87Wd2abSTmJLZRN8qiqlKCflJowkpf2d+/yOsHuSzdKkedZYR7Y
XMVCkPY6IqIp8OvtNKWehVaiSK7QJQv2zj6WR+wgmQhRz3OrLBWDN2624uzPH8rG
OLZia0IVCwQzdLuJ8ZI6feG8FWA8AV0y5G1sjaIZ24Z6IravQRquOepdz+tK86t/
4BUlz88sDG+MIwhTCu/FQvBL7E3XCih7FTE1pLYyr4NI/jLPQ717oPu3wz5XEqTY
NINc3pUTg3OZRTNAxBCrTr7JQDSFqJ/qU27uH0pi8XDb6yI/6dvGup59tYxmNek3
zSwPjAC2kmn+vLEuZYNxi3JO5jAjiZbut/YTiPADrcN7p2y0ts5j8a9RgIrkyyGj
HmVotPhGxioW+a/Dg/1K1W1UTpeYmPVxhKM+r0XNQYoMf9+1YJkBi6z7DY8MLRNx
OUWEmBzfVGYDdAACFlwRsJ2v01nMUaY3XzsCCd0teAcvSKfGYqjhtZ856DdJcX7B
6+6IHMU+CQM0w0LC4EIPgQSz+LF2YU2BUDUFhCADYAR0gyq6QMbnMe05le1JT/Fj
ANtQzBiaiNXTg+0GReQPBWkq6nSPYlWf38F57lYJL54xXH70wVT8Db1R1csLs96p
PydsgN9HF86mqwv3TPISPH0Ddb15GIx9JT4qMN5J9uQEACKQwYC113MnrN6zNuku
j4h57IcgnefUaglMhNna9wEqQCQGlEZdYbHXUEv/HRNdjeBWXo3hGF/sCX0ZXmAo
3ZL+liJpKibb/EiWdW3PRiMfjrpGNq1w1EoqyMKCfnhpsJLsW+8sQzrpYHmeAtvG
NOTM7cItRYe+3R1l5a/zSHgRTN8g1/NtqrUXj0bV6aQj6o3m0aSuTkWkjNdLAOXU
F96WI9zAUvspE9Nt17f240W8auuffW6wq3F/wqfh8Ph7RM0fstqZoxUIN+oQJOdx
7zzI8/JaOpZUmeaocmOZv7xLuGP9JPBnL7A7Wpo3UVaqXx3NdLfBzeDz7dJoLX1x
V9lAyaWVZG1mAOkRQ0S5HXsKbTYlRyikCHSdsXsgnK+S0oneA1MC3319mIGQ8+4v
pAJxyBgwXn+kRq/TJyxkhGy6HR5l+l+ffW9S7lWmOHj905Zqs4rnZUfQ3P3rocSf
fU2HEg0B2P6X/OeJBFrwSIwIu1vOBiQgZo8KlyJ5a0mk+dVI8nsT9gbkdnBMlmqT
XShaWFS+MOrBgA3X+HMJV0BWzX14Aak+e521E/JbQG7YSBG3HPGFFklmNmVSFBXB
4pVC9UqwuqM+lGuLPQLJ77DuZTEZ0WGcP2gN7PKjtxip2SalOkZTqjtNolvslctK
OlWHxzOk9oDERcuAbrqMtMc96Qoj+d3BmEOiTjAvX/+d/SEHENzqQnwgNjMOeFWE
ESmlfZV8Pav0xM55MFtpBEWshpZue9yjS9p5EZBzUosqsGZRPyE7U82PnHZq+e9M
mvfH5lf77MPWNrDpMVOTFVXImKre26BSARdVMvg75Y7IoGLB19shoPqV/leEgQah
Y0MU6AbsZgg5q56YLJkkvsXEgZ6A4CDsyaA9/JEU+atJb0BvS6TtiPR19QkCDgM1
lzWKdLCs8QuVIJ8wKFftg5+qsSO76o636zPDavDobIo54BeIRFHNWJeDXTmeZEmK
OwbCoX8Vz6cOgQVf/wWQFGJVU+aGKhIypae1mppsKrgK/NzPN4qZnkarM71JZcK9
RahZ/T9GX1XbMeupnTkkyGHYekhq3XGCPrLnCWu42lws9pTTfBiiMFCwgXZInTy1
xmqmnB+iC3bIFheZyGeG8/z52kMRV8e3BNIL/2kBXF383fQvUa6lB2ho3snUE+sn
Mp5IkHLuwcliuSA2mficIrSYvBwTYIaGyVSqLQ78pglK/TSyO+u9f2jxnEuU5nPw
n9uYgpNuE1tz1HxkO3B9cmNeHrmRnnTV1f4BC+B2dYxF418VzK3eYJbwRYJCX357
HRPdpDjprmJK1WDbdk7K0ZpTgedoXLTV3zqs79GyUC8Xtu8ZtqhZPOs73jUC7jmk
LUZdgqSsrgO6O2fT2ugcojo/U/KtbinLDIyJbpHpv6iieKjLqKSuzdvTGkvnCjMO
qcC/sxGJ2USU/Gk0A2lM5yalL5UlnbuXYKbB+I04bpdqOdcRFxmCX7NTrxj4ROYy
sJGkMntUOAPrnyAuEUqKOpSd/iR/OcpRrVJmTpuqLWz+UAV1wgg4+2aMOy8dIJPE
Ds8eA7ylqvEcBn2lGlpHYAGOORNbDsPeDmfs7ucrioLN9lQZs5qaVU+yPFfRNT4y
RwspvMRyxGVyo1mSEmuAXVhgKS7wIsb6C2htGF2bkfUJ/caDvoachZlkp78AxcyC
gSOeasYSfAguUP2DKdxnjntg7RwOuG6NtwoZe6ZrQEqlKaisblLFTT+uqKwVayRC
N/fNmj2UV8NDhBNAE/Cnapdr8D0uh8jfW42UJ/Ol7FCV8ElWrnBFJ2crzWlAglgA
UX3Zpea6zhAc8o1Rj64AcWbqBD/I3T127Ep8mIfFr28MitGlLOumRov05j7SmM43
tmykxsnGhNRq/6fkoYrMwf/fkJ4O22LTjbpwZODTRQMG4pVwI/e4l6CTMV0otspX
fk3EXwTxRGKQT722ii6UcMr+oUsi+/NelZJa/q900KedVMh81W7qqPEktdD51+pK
a8recsVSfIHLUFJ+CUR0M5GaDtuq4NDS0MCFoRLt2IU4Zv3Z6jVGf3pXB1YFBp64
qxYTXZ3eDjr3p0UL9xwr9G/zvztVHsAnVU4U6YpKRogzLRDpZdhEUQDJLH1+1XqV
G8SkJuajTZuDoGjwIhMnOVDgOE2pR8Zy9PxlHH4DAnJUR+Dage5vbxbSH+yx3Uff
uaO/DzUE21QGiyM+UWUBWDRdEJhitHnqzNN4JSY/V2yHUrR1WED/ZIP5LOaq3LEO
390IVtToCNTuNMcdQYyPw3IJMFshfjoZTEBsJko65pb8EfOd8iOlGd6v0384CyYi
7OX+ChBuMsAzY6laN22XauZ2Kpo3Si+CA66C3UfJMtEImB0jPHux+hJEgQ4PJo3F
tH/MFhkwWC1TIS7X4zvjp9EaMa29D+gpe6uMF4zGsulMSoeJbWmU64nx0KuDH+8u
pQJxWKumRtYXo4jjr3DGyUUbv4rGANvbkXfXv2vz2vgaWeN9BH2XUsrsmpO8/16D
7DClWGHKok8poNuBWlB/o6XTriLFnv1wE1DqKKeCVh5SreGRYL3nneT9yGl1Z1KG
W4EYvBrsFu2iIWR2oPasBF/+seG2Lu3ayOA4SsAdWbb1AJwarLLgg9hLFo6NcQ/U
c2WF//HvdT3Yb6PfoFzO9RCfwtzp/Dfc0InltKa4Y7ujrmJpaBgFXl9v+KgtHnBZ
3qqp/PS/EVf1Gjg8YyscbmXJL5Pi6fqimUsixhyGGh1CBNxhLOzG0U2oE+dFmbhM
sK4u7cgzpHHnPmqpaZ8wg45RCIZpP9yAjVVSxKIAgFqZe5ITv80mcJAziXIvhQ5l
R93Cq61Mwj46t5khYRMn+mS+7EejJ51vJmrw/ert0XHFqdqKyFuCiN9RdX7BzeqD
wO7VcNyQduMDHHAlWWaDVCcDJ6FGCHXePgjH3OJR91883pXySIAQCbMzNgstpoRk
9HJr45sZ5PyQnqDN1KY0X8YTR+5BznJNVngezBSweLObK3ptF5E6rxp/lG6M7Wuv
WtrKYI4UiLWUbxNXufv2EfDjVA1G/VPAIRfPcDxtPatEDGtGi8l3lBDCI9bsxuCA
mPVF/yQzVOwdRJWSWqC2A6A0W2mTBORcQ9lgXhAvbWo7Az41IFv2DAGAGsCRhp1f
gZlN4f85KT6YeMD6G5e18Tc5eX0omBX4/+bac5+ftnHR6RXUhJh9F0Ro7/nVrK1C
1D5ITjvaxXSGANmZSkTuoVJoDPR3dttxHPRRF6Sk7XIEbtJ/X/6T4Fo0Ib+l412u
gsjEM+GEqCG18VwXcw8nnk88cHCu2a6Ji8X2e5QqY+ncjKbBqnXy/LpGiGkU2ngu
D6d+uUDEEFUk3XGpfWquBjifVimRnSg8Y+BGYPCWZ21E/TVP1VgDfnLJGtyDiXct
GPPdO9WSN7Yqn6J3o+IudoJq+J3BccKcbqpRZOOE4yxTuuFay9jkc58foW6PV9kb
zOaSO23Pl7ROoQb1mucHuE7fduBV6NNsXTeiBNFX8nLWjCPfIVXMjeaxC/dlaeHo
eOT1cLwQWZ7VSfMjUobl1X36Ig/5ks2J4WmcHVaUATLiOnuLo2iX0XAwIHv9AirH
3mPyb/NVaW+u18SzOmB5S99MmwhAEgQFFlKnDMI7IWhCzRRGiQeBHnouNoybERuP
Wc4tgMva9Dt0pnDmkEtDZZKivXSX10gJYHFOyfChq6dzhLi9ZNS4VTkxV635aWQm
c00+eVXJVel+7oytqGCVUcKZxvYs2bpOjMj8qGTUKV/eZ/lOfCGw6bva/92OrMbY
OE7vBAX0HQ+GIoJXglsoEQPzI2xnJlya8wkeObSleR5zCu/o1ewnwB9qlQaT4gAH
GRiieQqIeUaX8DNgKi1MBafeN5cdbAA7VODUxbegA7dWPZklGZp4W3zLrtG7t5cp
Cv1W3lwNEDU5HRbOlkbLxLJXj30R4e5wqX6NvTfqZu4hqF6E3ihRsZRNo0i3zIj3
HRV/dRlaHJx8sEIRXoIiC4YmYE1UclSFyte8vikkjxYQD/4tByQMBIuUhcgfbpBe
JW7sBR/zoupyuEVyvWD2dYxgCDznOAz4iTpuAD8dqgAj+oIGiYtN4kJybp0eeHTM
gCBp9bOyD6oOaVyqCesLMTSdWK2iygXgzPuQZwgqvqmCyluaJKPWQwy2HxpekElH
Eor7kkMA/mU7P8tT9hdD3z96jFeepkkT3WeVelmgzF200zDTHX6EkQMazlQDrlHp
kE0iHfAXM0UC/H0BNFqbKaGOq525Dl5I+Dt/axnMBmX7AZjwVxFby+SINpA8MG2U
Wwks88DdqGYzormlBw0mvEbU6n2fKGn7EiEM9HMHoBZvoZ4ka3pSUs2QwderUnMl
+fbZLXB1F45E0zKACLk+hR+bM6FaeBWhYu3iEELy26dVoz/6JgHvTJXe83pVl/AH
00kxMgnKbQFWgsbLeWJv9cwDxrNrGwOsKey9nJLXhuWmvqvzXVwd5UT0rs9oVIQU
Yt8LV4PRNDViHgW1xEJhIiN9aJ4TJefKtClTdhhnZcm/xgt+UTdzqU68O+NJ1Mmr
zmIIe98lN2Fyssjssc3HrF8GaIMw4HNUjfxbnmc1Bx4YP239HfkyH1pgXtYWbHYz
UeTnJ3jOeZmFgkJ6ie2H9RNgl6m1LKOscPjSL6A7xd0tmitXPlCj+owQqB57+RVt
ew8Aq18qrwHYcinODffqIVON0uBGkravVHKMtRV8wZRKgZELTuKj+j/K6VHjfban
VxGGELPF9wgJVUWvBQ5BdNJMNAsy3xJvpUwymn1mqeR+hWon/p/tsBoGINc2Tpsm
dKAsjEl6VZDVgPu9IRCkfGB3lik0UICxhnRCfJ8un8goUvOrbgwUq5CWIQOiwS0y
BPkKvRg2lSMPhr9VOn+s9MYWXootXLwSp8LwHy3rtPrufzBxMn3tfJgo8ioTaW+e
1WVBCf0E4WilBCYP0p0xdDWbk9YvhziA1kKR1FNpAEANkoUw2YRZk49EYmcXhrC5
KuTa4EowFYKPXs+x97Sr89s9NvrE8zht55M6NHSG5PyObIkJ4nHeMlzJ2xD7LbQH
BwMG/586zFaPlLSka0ubk0sngWfRvW5hoduEtNtfE/RkgMA627ur32WMFyLIpTsC
OjLt0RIp0oTtXJYZj5spbLmxGt7vjYpTYJy51WVb1433/faXEtL1aq+UEg89zUNf
nXS7Y7uFAuG6uTpuUlSzTfVoGEXw/4tmI9QNM1BpA7GFcRcgsV8po1q0Pd8ccLqx
YjrJBLLCN7AZJEOkm7p4CL6p4wtXuBx9qiEm5sh8yE6EHD4MNkyyfLlS2fOYgvCM
jA3Nxmxv71riYI3uFMkBUnsvM2Tk4Qi9KS9n3eRWW4s04jeJTcWxJyGb0yhizNon
2hsnsfIQxnbMb0OPka0/5O2i/il2cSHe3lL562osTfga8ZqLoHuz4sos9SKkEn8C
i1W/hC5JuPjF41xDoyRoF4+EQMzGDtHktUrNAYSqlyYlOp9Z8m/Ikehsuj4qOT9W
+PE8zusjDBK28rOZinjcSQDJx6gOj6KXKJOlubQ/W8JTME+BwsKROmkC3xadbxKI
dO1wtiqg8bvkbYWyyZ90NcsrqYJfg9QpaI+GrnRB8FxgUZ51ywgOkdtVDiXXxSk+
RBRhOhECviQ4mRbO0Op6rai/8ZM49fuAKhmJHtoDc/29emb3WddrAPs8WykKHDPh
op8q5pKqzusBaQL9HDfcWlixZc0r3H1va4sm2nKZlOQbKp1lf7ADkKx3lKfFBPmL
U/aR5nWHtY/myr+EaiBcTddVfohhMnMO3dR0otEyQmKJeGbJlNowEF3XwDFtfHIg
OEshe0vTgtnzQ/5jAHgSJINuEcj6RRMEXWMOx2NP3OvlRXkXNexOZD/XOLdaQLtu
tjArGQ4mWVJYHd/spKcGAfLa/bJxFE9JNm1aThgnU2v8uI8lqRWVQUlwh4NMbskN
uS1KsIr0pAnckemRbT0sYs6rrDBnzcbFkiYBUdCy5bt+NFfS53yEfdtFonbyFU2+
InrLgTPQ1aVoOkc9dGGvk+sT1QXlJnfO3FvCj94NUQMR41nQeI2Nd0z/EPsG/7zC
gfMbOnCWY59BgEitkuiR8YFQJaz0ujq9WOR8+jV0WVpW8LuOAWRv/x9KY01V5pZY
MI1yH1R2x0jxmiFWudXJm/XCSq5Lup3Cc316uBgbcnkG9owrmJXH0jh+wUlU6W1b
D4RZX3ThasWVbBf+h5FRqX2ReKjjrtIsAR2i+PZFV5T/K+6bb2pMY2/ZJe2Iei4F
b4XLlVPRNJEoucN/01QnUNxa28GTG7Nhw6tfU2t4AWUXJraHgvaUeL13z7Wf5Att
2kAOVG39ho6AncTOYfMxWKjSu4Oqlj+qpgr1SxQguLfdM38mU3lkeBWgF1NXLNgQ
Lx3E/loQRB+LuijdsK61Q7t3cwkVNdHsMxPdDz4osHfNm4u2hzYEQdGOhPUhTjYL
w4nYmzsCotJSliLmB2kr9OVI6Q/hnkcSunKNLwBLykEed20hqKIQzNNTIuMvjBWv
8CRLBTzIN8EinuX/gSmeZe6ZWqjRoNUzr3sI5CSESUCbtzVUjKbmh6nvxdwXCCoe
KSyNE1CsXgTPAtvkaQ5Cv0TEYxukCZYHjbyOmKPCPwr7EBwamXJAVUL0Ci8iWqtK
xkQtDDFZGMWj0fYa1IzlBNSG8K2MTm4x50XCCxz1qHHUp6RC4sahyrpqTALavO2f
8BeF7C/WPqeRxpTN69sfrATpmx5eHWo5CGJA6sJylwM3BZ6n6uQ+EW2hJdmGL+n/
sft2IAgyYgEs9FrIQxaLX5VCvmmBf6Zfy8qhMxQv2wqLuVDhcoTXLvQHWMKhAI+k
QMqnvbsE2IFsjNguzPPf8eRyAb8Ch38r+nBMZWGvmWrgjNCJFXvbBoRvROISDUSW
eGKiOhocPsRiWKjiQs6dHmbSA9N2K7ospIn6Z2O+W0TSXvajmVodYlo+qOjnwMpd
DRqKPLKQhHuqMYbIAGkWwGkRXQj6Ih3B2lfLFwJpMo40GGuvgdqQEhQq7Ii5ZpCP
I1vRwoaiCQPrP2JkwFk317ZpwSLOnFouz7Me5GYVwXOIIr0YXt2B1/sJKxzymkuT
QS0gGB2TTyDET8+74HMKxzD+b96KiRDFQ4wW0OC/YE/ke7M7M1jrQeaAaDalaJzS
F4SMdiG1SvU7a7g763aIn7n2HOUVgqvk+ZMNzJU5vOJkXioQmAyhdSPxBW9RAMWL
hWNCt4hlsqixJp+qiuL5NgNCygGvMNGVmCCAbPky44vmUlMWX+ocDYDIu6jPRyof
2de5snVVRfeZTQf9leglJd2k9HpZ+NvUncP00x3DdBx8l3seBopiRGStXq/s23FQ
jL5hbrKIQyVmo8/09mkhjUVzY2x2Fz59/dAdWPeSx8LXmfWBnYSFvpNEFuPk7Hdv
cHs6PYbKaKFeE2AlcxlfiYug4EsxJB+0cagnVWU7+oDsItHXv7tvXb6aYvn547a3
N+ailBwLFI8vEo1TSvx7n3QCKSMAVQ4PXCUMHg9M37PIiP+P0dTK6uUsbBc+44uM
FhNKCWKGyo/aVSc60ZJr/pi3peb0kf43m/GC0ggc5fTHH2YSo5mhP+SurHO9k4EU
l/k1Z8n+Q5j5ijMux1e4toxTg3MKfGo26pin3dC0jcVBY8mlVfrwEjSkTde++kIk
Eap1lhWs2/nLp5owEjG+CDh5FpYR3e7Gij39+WbGAltJgiFTV07152HmUADE2mig
EjNm1HiNJblnPiexcf/zt+gj/yhyTzBNuk52sJouzAhBaRPIdv1uteFMoiC3LNtm
l8v+IvG14W4BHslUhrGSPniEdUZV+S1tPU4b0JDXGQTK4J3PdzYvY6x8OFdbhNf+
CdGKCqzff6MS76Sv/pFN+XabT8X/F36x3OkYhDydTfIuHmxeS5F3znr1lt78hYhG
6/L3p7aWxUO45cfg/YeUXcgd+EMoLgAk2wVCdoZ5p/XwQh+90RfCsyoDoSm+Q929
3vaFUhI/GrKw7vR5p9+x0Gt8PC9j596ehvioPL/9W1EHKFBSq/thGvDs8iuYkQu2
Lir+R+3QbH8jiwtNat0gWsoXdFigLtR7oaKgTIwWCDrJ+89fE0enQcp4CMXtHddX
J0g2rSe5JsWyp/1dpR0NiAwW6I0a0naQt2olwwlaPB4tUfIsb/nD25lgwXZFrALw
dXZI/+k2HYuGZzeaL+a/iDUt0I6swcIlzz/ta7TPqGTGF+k1SU3g6lKgIod4OFWi
3XA3QbzI0ZjYHQHgkrS/aoeG5CIbQ9kxuPx2DkZ5PDz8pJw5T16ycbLeqpmqK7Bs
PiWmde4c+uj7SXkK5RXLjWvH40dFYHt1erDb373xk40kO8RTDEO2wET55ZugM4oJ
0jrqqFtC12BsKQzhi6DETykjl87VIA2KV6GnUrN1gJIOLRed/d/Z8vQh2lsGVeB7
57/93D24xUX8kpk/aYab42zrVTM5Rqpc4NM77U58Tk3iHw+MISo8cMyzeJUhglzt
h026+CUGu+LB2ePsLMo+t3v6hLLwdaumMKYVQtJoLoYQxBPDRas5dbSF83Xt/MOO
5ltSK1vPENMTu48PUdjjDOv0h3+qqibFi/iSYx913LJGjtJEIiQlwJRCrc9eOhlE
YFGVvYhHdbI83jarWDLlcmlxjdBPTH57dap7RRzXJZLF1/7bMjgzSttB2XvVx7+F
IavgblLbE8WPdRKJ7OBs8nyp79c2nKIP7UzE8cuLGNSTIKXFYtsRWO4mqsm7IwS7
vSNSOGUpkYAGTZVeN6zU95HRQGJmEgDwlGtC60tj4UzBSKwRPir75QMuptvSfvwf
wODKpmNQ0lCtMfTVkz7+a40X45poVVxDmF2hpzYTmpQ01UYea/0vrxFeWH2PTIct
GbSIUgh9WZnIPDGCdptNZZE6tRmbQw/jmbWf2bJJ7T91eXcuVQbtqln4g7j2Lj+h
zya8SpL16CO8GLlGm4wnZJC8omhIti5UEwDAoO1EKVMqRuF7JJhw6peewC/If+Pe
V+BYc/SbWmNRs3gH7wuvwBaD2v61P4+05Zn/OsZAyocE3XZvtN2WplcxKtXYLbMX
Mthf3LvsETr9FGGBdwtkL6nvXKf+VYRXvkMqnDVHWBSr1JgzmIO2YuyFYI4scdvf
eRz1Tvhumr4xEdX78EfGXruiztbfffvEVM/L7ful7F/teVMPzI0ZTGLJFnNFwiQY
WPoxwEvwEnZpvhVmtTCTgLAeIKHF2ndSwUXs+pwzAY/L1EulOm+iq9XeV8IZ+tcA
J9Fe+A9CFkEEn+SDZQ9Lxd4g5leN4qqdmHwNL89r1mHYhVULxDoMVWdRykyrmbuy
KZ/ZkqxssigRuKax0PatbRBul7HFc98H2rxMekLc7KG7/1IgDu5o0e8KTlFQ39yz
Rt3e/3IKvTrLqATwCV9UsxWrGUMmON9laQiOSVHiTrRCDhwJJI1NZxTfQ94KpqSN
v5x1tourEWjAm+L62aSr3ITOTSR78RlIhg/T5gsPJOrG3G2eBTVOP4DEHOCat+gG
WCjvvEXf7QvktRufanLRkL87tIttILtgQJjPltqvN/xQxM/9nb9iDI4vm4QqICHv
g1pQStocRtf9l78zeEzKo2dipzbuwTnkBHZkDuy/XgS79AWeiQjCp6P3i3zYfu+9
V4AuVS57N+GxtoquZx5GSwg13UE/j+4NmrkU9VGVieHXC6qrXXL84DSIeBi0WWEW
Ty45o7Ac5hxacw30ck5vcio+Rmfywx+VYtr7Fthii/bpgs+uEPHXNn3xFtgJWsNy
8fDstfrfumQmT8gsgoVUu2pbu70gkQWrxusY9hoB+pvWzE3lykJFK/BN85TZdKz9
D5RfGqThO42/4948bbqzMuZ09eCQO7zQDnzDYVIuD4G1XImEKQQ16SkBWFqQ9eNU
QpMLUl4uN2OolE8H7YO1acNTVai6SU1GjkZF0wLZXgrH/NP7/qC8mXxIVOzTfTrC
wVak/AR68SyghGJRu3LoKM92OwCnkpf2YrtzMkEuM+nTWxUyJlgXWwp2YfVp1qTo
QhGwmbBF1x0rd92JtzU/KKEWLoUEsCmZtesodHYbseMQ3RKR2TzEmkvZlwKLwxag
kO05/XP74PCNwnMTLTcP5fbQdL130HJJHJ/NgVrYYR01wzlU2AbpMEcvMaEU984I
sZlAk2q8tcshHVxvaTfsIG/01fHD+wM/wHMItBofPcwzxj48IS+QChCTT1hzqZ/D
4BbZOoL75AoroOAHQ089HFGpuqnw5BYhGC6zUZuxRrDu4k/gHMSjhjAbgWL3F9PE
MRZzTO3l5tyJHp3NXsEFsUdaGxHy7hIj4R+ftje07UfnVsgamxH1FEPkS58waTwM
eulIRY+vfyPe9eJhJCWD7QuEBqu2cvbvDHLaVonfDpfrXk6t6FbUV8Az4rnoIbD9
e2XiayfS1vYZQEHdLiCiPtaJ562x/FxUloGVojgaz5x9PzZTP6a4ycsPRg784TTT
c2kuAv43+V2edVE1XtESN0KIOQySQwFHJtN31PgMqcjNM4UfS8JYShGdTb5IQcLv
eGcsc3UnYlZFIXQf2er+8zU+rKZsGV7BmJ8mX0gijX96a1SCrEgZhSIQ9ulTjQSe
9l6391gAF0iLh2avrw0g/WywlI0gBa63iVPfGx5ivDzrTrDwRETLHvukfxRHaI2t
dlgQD9fu9+9RWRvh7xzeEaEbS3SaBynwlEg2CRVWXcjl73l4BrzU4nLEWCMzNuSF
d/MH7UGvt+P+ip/Q4Ou6am2UrTTlQ794yre+RrZvnd1w4pGC5HVAw/qLP/xUR9E0
h5E7EIF2aTsxFMnb/Et2xeAHLqYNSBwmC5Xgb0ENmUqiMgrPcRC8oHFllm0Nfqym
BdTJc5QQMWMX6bTRho64v4uNlw5/7MEiBcETmbRb2aQyCzVnOPAIVo27nm8k/FGZ
nyB2BvdNAaUsTnb7rc6018qo2h0nl4Esz5jxJhRKzCU4jRXRPDAK9wGIdT/YrlCT
E2Gr/bTuv5Z5JiVeVPtdVdNAWDP+HEg1Z7wXyCmMLrFlh05YoFOH7fUPjo5b6I0B
eMC2z5b3oOsMpr3hOsU99GSm2nElXjlHoEuoknyjCr2DfzvKFaRMoU5AnaG9H9F3
klSRCMuBAZiLPU47+wr/1MWUhAnYaURE9bGctECt66tYdNNM394jZGKDfDrqfsWh
VXS5NFtiJEcKthfPgj4kVlpPQyGjnn4aHUAxF3m3imCmZXd1nmDh5JvChD74eZoi
Z8tnixkJAautu5Ew+gTtWkqzdnWpmQl7YGbMjVLafuUKEVQFu5kS2QAntwjAZlZb
NbKplsE0tZeeKBwGV3ItLqqLM20lMIDMPsV+pjxh/OMMJVjfa3Hc5zSgU+GPMEv7
VzhM/JaxiEW9LbkESxkimYUVOKqMwGbDIPfk4waL5jd8s9Wm4POMk2ibNnSgqk8E
hXAu8JzpennlyYb4szc/Hi/ZZXlEbJaNSz+tndq/XSSSgvuXmK9rxUYmPmzZATZt
r/i6Z8d8ixn3lJ4qofo9JqwSq7QIKfel8VUIi/0g0AJc0pHTrPMdkK5ku+nQE+kJ
orkrfKKZUG7SLfYrPpnFFtL+YiTOmOuOwT2Sh1UAKkHCYiNSkmFWxqk47CZMkt7W
GMgM2O2KB36gK1r5wiVaNFf48RMJToVvu5tGnTgiMgT/KK6uNTeJeqEGV/CBWAW2
n7pE59AsynUqaFxy57jaSPJVhtwFKHdC9U00ulOjyyA2TqbBhbm2eYV02c+7lCw+
POASVoe9cB8iCnyMa4jR/ptAfe6AYDCMwmGWdV5ZyncPHxG94gs29j8WyUW5/OZr
1CgmcUC0N7D1p7aUVYPpIefiwc9WbXwRNHDb656azW74qfCBMj72jMSbszD2zJsa
0n65RC0Rr2Lu9Ad9GBA5J4rhmOwmcIEXXUUPk93ZPb1+yF1FPzzOjweAJSuG7S5i
4ryAkQV5RpMhEqqj9VC3Xv64ZrJ7s+QOT7SYlMJwOig/Pe2dM5DqtC5NySqZaYgO
oIk+3u6U7j6DHauW6+XG1N0vCOC4uGElI6NvCodaN0OU207Kulxr/OLQruoP4pRO
q1OV+ycPJA0Trlcw2kQQErTgDjrHb38Jw34G4G+UkDQbFaN+PRrB/8qz4j5ZiI9q
kvrWTe4AoF+QupIn6Nqw6U3He8JgYZF59FwW93bcw3cS9Kw1cb4oNWzJQtgdiYl2
5Lx0Y/Jz0I5XSXtLy6YlvR1y5HRhW5Is/IVfhq58DYfVZsagmDUkPoYHGI1Y5jeS
ddA2IFCYLYcYoXxSZrdObrPfVb3SnVFJwdo2tqORS78gwd8N7NNXtS5QOCtV00rU
eZZMhM0NA37xpw1itqR54Kx08xNSOvNkjYWNgMqpBdli6zwQE1VwllizexKTZ0Lo
SYBEoRzvKyyYGv4k/6FsC6eSCY2jpHgkvRgCv0D/hiJM+vEFSdYMBXL2GQQo9BYA
/Cp4I46Njvjxh1MOItR3h9M9hE0bl+PX7lwl7VChLObNUvvSzofEzRjwmdz6M0DQ
Qd4UUnVOa3vxtEmikeQf3HWosLA7JKNGJGZUHbATAYv1lTKX0m+1WVOMadxmZsIp
lPgFDm8zgp89OcfgGHS+6yW0OO20kZn98poX8ICUzqbIwJdaq2IZZCFzZZr3MiUz
zLLo9B9r/KBwvgVyjs3VZKDX2+pTwVGhOTcD2IVQbEFK9PZL6Zv6w/1c9mwl91Bx
7i1e/Os17Lb7U2S73E1PCInOpq1Oc26uEJrZCs+v3U+DbsUWzZdO+1t3WpvuPb7b
xayCCwEN+5kvrXZYbJRGSqGgwhb3gtk8F+8yAkuuz0A6b2d22WZoQ/imkKtl+xlu
ksaRGGJLLy/nZCwsWOmAf4ESAA8/YXrmCfAVr3ZFdvQ+JowEveDQPVK/nQlGJ6t6
MVZCr0NbU6WX7rS8oQDxbdDRFrit/YhfM1HH7DMgbPxExBRNkr8cZr9cXQ1SNFR5
OVkstP8vr5jY87M9egfM5JwA085yighk+OGWFi0GvA3l+R7rq+TA27VJYXY8LEk0
wVdqDWPtaj/bJD7519/zy4Jkq7wezwGDlDqMtmdjxh0UsU5OsX6UINsgzUWihsyc
FNMaaRB9emZ6+UIJJW7dHyWlkFChKAJS2c1Alhn1mPKtFtZ2JzmowhWEJgpHqxSG
f/fLhl36nWce8b1kkh4t285os+q7PC9HEfZgnE/pKGWKtO0XPLLtfZfTaC5XDCmr
8L6dK0C+MzOdIw2hRpwMrMnR2Sg5cK0CpMIFbBVv+EoDI80ob6jr68Mzc8QGmM+M
Zi1UTsDFeGQ1a5O7Y60ry9LY+oRVssTYMpQEnosNPT2y7lU3JmW3brMO2QiSxSwq
pOVRFB3lHUtMY+910F2mOsOtPHeV4mJ3VXfE2Fex8giyUaidzOIdehBskpCIotGo
IPMLcCtnh3zyVdyOf2998xQ4xuevbMvXXi0hWia1D4rU1CvtfY+keBj3Da916rjr
hPTY2DY/WHjlBrP68krDRM8n74BYXMBmx/mlwNGiuAM0wcMCIusKtelpkk6mqPl4
1ERsNrpLmGd5BVuoGoAb062w502zM8ASoeGLUVHzRjNrOAbFpMRYxWKs/B4dfnV6
1ffXjkPjmRmkM/a8LjrM5YstnbnKrOpTqwwppCKVp5ORQ8yr8hIyojBUF3lUfjI7
AXt7Qxxn7MFUt6FvN1D3UZlUtF8CDAJ6o9v1HCwZ3IrTfuPsE+o/ELR8LAl8H+0l
BA4mnMuKHpCYmHJDxJuYpFVHMuDVP+Lpa9fUXT833VeyMV+gz5Yz3+u2B0gqjg+I
qNWrXgQlznUKmRS57JH9xh3giscFjzpO6nGxPqaxjnlqL3MA5RWQoOE6xIfXjf5T
5B5OJZIi6zc8IPXnqgWpv9xP6ach/bqxu4kgyGsl7QFfkaDZXRdYA0QfyU9Od4V0
S7v/de4T7fIJ/5f0wP9mNFkDojgschHhmOQ3p4AldrcwS8aBd4/cgGxuuUdcIVl5
OxxlPMJsoHZoDcYkOZ6m0+scQQyAvpc5/eKWB8UoJUJSCPKDO+rCu7xchXr3gmVW
iSXpEiNFHACGhsdnUBb3RCj/NWP0AdUFLxXj8aYTtN3me90eBnRRJgJ5PI8q0lA7
Mz89tVR1LjmVMeKvyDMg8odhhg0Ig3TUp4KnIcrN3oeayknlvJTRk60/ctGbDcJw
vIb0P4Yz/0KPaBHIl7LsY7dgMs0SOSUNqJUbnEQPf3F/7ZNJkHPW+vV2DQTgvfJE
A4PI43KuIZqTOrmQHaxep/krcyZPyySYkHhTPPPQ9r5W52awzP1V55cOWhNbBqgX
9AS8lKOzwP8SibTxd4mGxlI/XKNmXKfvcckxQR2XbrdCpXpgD3uAdHUYAeNbMMB8
EZ4YHdnNCj5IB6LEsGoLHunnF7oOs2VnVJO79HOJe49+5/Xm7QwnIflwvuaYF76F
PqI8c+1TAiiCXDuui76xxqEaF4KQ/A2QN9APIBgOpFUtV7INVW1eQSFA46KdWDUa
L3ZOnS+n8feF1uDlqpCU3FtU2c3TAxQzHIXEGJPX5sW5CCyP4obipUYyxP11r39M
r2Xj/7kCseBmwcdX8hAFtGZbAFtEgbrg+QZCYsYRy4hFGKPC470Qa1GKR3bOgHv9
MFX/wQ3+q0o9jl7V6BuuPYddo2uTKmyMjmWL8jrOm1X5X9+yFwOB9CofqMznFaw4
nBr8QVbWucHGQfc4CwHEGWvDDSrzHRixDcRWPsrK+/rJGQSwqULLWum531NcL/gp
FX/F8W6PISYGFh7CcXtXg2+ANc1+foCoMNLHj2nu7Ijyc7qj9C4knyrE78rsFv7w
NPsRHaaKO8tEIz4XPhbQ059tyz1+N2AEo96dElRjKhppdh662+whj4DnI08THHI1
0l1XHl2Q6PNb1KVwwo1x1929EjwbieqRY8gC/WYF7VmsWXlbSkgjjOPruI0zzBnq
v8Qysrd4frF2U0wfOcYoQaMswwf6L4yWdbfMbhCTNVJPKt5eb7npPL2aqXW/C4l6
oXPaCVUF/tyRsDqUrNN/9CstArBBi+2nVmfImxCOGgb3ncXj/CbsPqj6DSTzggtF
eMhctayU/BfXQqjQuWOOJwnZsyQjO55XUHl6oxrtVlV67ozdhmbBrApDr453ZpPw
yQVpirzEp3YekviMu7iJV6IJ3gWTB6oG9sB/pBW8FgJHK/jt90FYGtVXI60NaDa3
chOHPHpq/YDw4jCmwL/CinVmpK9i5UAN62xX57AVZlSdCOWSXlAU2Bvd1BvSqYK2
u5waxBU1zLXNRNMPnvVUXW6DHYBeas7+V/hn/YEAhluoSd+qjECmMmqM9A153c41
v5ifmM/ETianHMUCkG9I2q6E0eXA8A7Vu7fXzv7VWcx0DauPh0F0xflRcfqvaOVY
H/sXr9MCvYLn7irhYiRNMWH3bgDlT0SPFDjW73VuzmBe6h/dqCEXVWwCWeSPe+Ua
NWTXELQkrQyLi0CSvvrJWoTBcHJF1Rxv6CHy+WTDu1WLy8nQuBRD10AFyYUOsTtO
S6Hor/N07UYqfItni6TzU5VmnNFIFmEuknYEoK9xhp1aJLGxqi3piuSNLySFQxb3
N4Oi4k/llyU/Ujfla2TBDSmm/bMMRrhdypKgCGD8dXqStov+G6OY7Enc9b2rHf12
ivkKZ3h9ad4sYK4660BP5zc8izBlhMnS/iONVcG7UgPGTq2cE52jqEQz61idLL/L
wWiYcyV+PlCoj3SlGnn+9EFZwqDhBpt7pEr3aS4eFMFIIcqvBWTsm4qcp0wLBJbe
BCTerh5Vk8GkZjr9s1svvMTTMvZbIsPXcsoly6Ue16cOq3WvFihQ0sS/jtSp2ji5
5qSfm8w7iRSN7eROi+Q1rFL18KGR5e85sqxSazIjpQ3ZNbMEXrvzrbK9pcTDIVYf
I4mg2IlA/JU4rkxk4M0YzzifWGOuYE4vTw+bQkVIOQ6iaSiLi+KzCXdLjmQPaxGu
xI7P9165d6Wl4PWKuK2B5HEwkphLSdoZ697KY3/7vNeXpXSJJCIrkWpHEM5qTk0X
FzTj2m+7feBXxjImQsDpcPTTOeENqvAuNsLkxc5ocTFHqPjoBPJEDuA6fG+mg9o0
/XAb542aG8oXN/B8l4PuW7B0ClZ4vicLD96XNhUUKZ3M8falDtZcR4hf2cmrwb3g
qYKmxXyjUIsFK5L3IXPJZJXu8lF3b2MwjlVZp34DInw1R4ZUxbw/J5kBEFxldrDn
oZSXjt7vZmh+nR8A893KNDJUIlxDZrYYc1wDGQ9X5DeY3REr+KJOlNrCUGZL/6k+
GwdG1fYfedoGBYQePsm3BCCHiqxDjawU5tvr/EFq1k+W9rwivAUnyDYxL9jBObSv
VJe6Mo479DVpGaRMPLl6Zt7B3JhBWGqCNKY1i3YOyB3Yxx8Ad3ajCUpCmoiZbg4L
ne2zgNNSni1fFT+5XbJevlBSYcLbokfYMHiiUkp7NlBNPFxF4f1I4BUhkb6zLT0z
33PfULx4r03DKH6ryuUS0X9ICox12no0rX1RBNUc7YqFAGzhtGljxM4nBujCnywU
ixZ2UDpRIPqU+BJ75wz7iM5f9dygGxcHru++9V0NcARHiAuKmhKpL7yLG8BXIdnm
upY7X4YNo1fE09SyGXtpB5QrgVVa8omq48Qo76gDNll2eEb3f2XNAXbw89lZQ21w
z3BLbYe06SsrWs5fqh3WqeX7boI4Db+0qDtkkIblWE68nYZ6rvg1VFKndju88Yh3
JHSVzj1hmzkJEJqmSYmXyZXAYF6QFWQiwx/c05YdJDRUJvB3Otrd0xbGqB2sS7xW
LT2ugvDBy+QcdV0fHKOPyUxi829KeZrM6mfuSzPOxeJxFDJTTHjIBcXcX2lefE3c
rAkA/UW67pu3y29zYprTJhlG/qJWMha8kkVee8dADXoD6ls7fo250G1PrC25cgH5
3zuWABiMzUaLBd/S4qJwF+7h3E98uid4c222RYK/n3aV7C8mvntfARlJ5wwCOEpN
VL/48yRYZ4/xjIZN109Egs7jtp5LbNasy78oMxzxBpmJqWLqqwE1mPMILeZwRaLw
HmZ+3d2YQ0s6e5ivDLxxBSW/nBVo/XnlevETARCgGaiwitiERahIGnSBduqCV7oz
yTNvYcPiCPFBTlD3Td+z2jxi2GO2yIOEe5AfkWIJWOE/ySGp3aXGiOjxkud5oQv3
17MZvVPlZNrdDUpa9313WZmzHs1PGvM9MOHpjE6SJ64VrjWqx7tPbO1RtSTVagt5
1B9EAmh50/aVz2/CoovDZkX5uXm/IHQoIcOH2mRzPAf8oGEACvIwclu69kl+ViNj
0lbV0bsHNBTSmfegxcm/rJJOb/S25SIgAxs9+n594OBURIkZ/+BFmDm/2RyDHFf6
kv8cr0BHobU5g22eVmHtYPITkZqv7Ft5OC/qGVZ8f4SIIjQ/Yl80MQWCKf5IXfOe
EnmEf8CJn67j3WozoMzZLVr1y17/yQELP2mAR4IqoTaR4WzNh7ApubUXT/KzARpG
50LS/cYgmdmqs0K1orjMGb4vfle3SAl1FSsKpOVvg760zv8BePKO/hFcxk9DM1Ti
1AcwF6x91RVcxpDdrwuNcFgBZm5caQDgLSlN7/lRAtVeQP8HrsCwLzFHvkb4OS2Y
ea4OCUt9BtcoSIMc5EDa3SM5FyYjEkwb0FtG15o2ovAMyi17i7JrZHbNZa3qqRzL
Y8Jw4L4LTD51s3oyX94wZ+/moQUVfE316xYyPT6HLAfBMYghKYj8PWKD3JxZSvXJ
ljzdTYGJvG0zsobmruvuVCdI1SeFzz2TW1BwVHgjgYPDHIZBZyPjpMX+etbu8jvf
+29ppjwDOtdYLZqG0oQUYUDcIgfdO/B3mEgRj3Of41LdO+q5IZ2eK2TmW5+eMGBX
VMtVTrjQ3M/Rh4tkyrZtaTaO61KO5NLhRjW2E7wRVjnOfXIe7t+Q21/FKAKBJEfg
N5dQPhBHa3zjWbotDpT+nub+q268p7gefoRRZPYEeHCt3/ccdVFPNYAbjpOZ7LyV
Emvz0Fw3XDUT0eU7jIag3AyJx2w8bCYAqhFxdUqVYU5NaxG/vSxJxaNPuSZA4KUm
YlYfb9OfLZjHxTM3ood3/KeBvEIFLP0oiZn2oHCw2oeOMuP+2Sxg/3X8ueRH1FLR
7q3hOl95ChnptHzB9DhOAmknHdG645pNk6sSXktbVivZjRzIFSZemLm6MP2elAn5
GkJgy8SvNC5ixpsl14V6W3ek7mSujneJ06lPuh3o2xaIvtGtT7lumFsTWmsu/ETJ
yvEZOLi+p84H/ezQKrsQmU55S6vyV082bAJDVt7qp4NKTZJHCFHHgOpS6Fb76F00
FoH3yPXo8Q0r7l2CeEJICC/eEANd780jLrf6R8iESnrWO6IQ6/yBTSZzksNecLmT
KLUk0gjX3pgtG0aL/paA8Mgt0QKPWfXfNcIHUOdkrXYC3EAnSIv8/pV6cok7Kf65
Lhf1WNsC23xE9LbDbnSpCVHdpfsPNNJxQSrUCMSbvzKGq+dJ5jDNNKzFIBRiI0H/
gO1bawugAIIDOXOeNPuXmu9Q3dTSepJrd26F5uIt5D8bpv4M7VBQY7keMxxOPc2h
2nKXhmLV77qQgpaGL3TU1wxpqhFsvrIDtGY78Nli3an9EGC0axRoEKjksfQJXCWI
WWXrsx9aydVxbDVugv4OqtG36OkFuZMOLJTIXgb+rzrAsu/J0qgQoJHCLnE9H+Xc
UNHnc2t/NqRLH0zkQ+Q66GvVKdUUOefwXB4sAbRSlh96h391mxAB/oWp8J0OWtEo
nAfBG0xNvRfqtKSBO3kh3vUNX/PRswADRu2EeUkHXGwvDtmdupFgJE862wgRYcgp
2cSJh/j9OsharQCNS1ZghmHNNm2V8Yia9nFdTBI30U1SKZVbBfP2Ezuvzlr2Ahrs
JS2bvTanXMa4pUWFVZu8f1RfPu/auSo2BTPW+8esvVrSBZ6bVP/2kuxAktlLlStp
4Q0E3H30g0iFO7e4mCanpKU9POutJ5jqDJaucZUg/QziJ3EwK71uYx8mQMc/O87Q
QmZZT75ohlBGRYG8qvb8aBg4922hxYdUqHnAKfuRNJJmrZX5+3yb6LEyj5pZuu8e
Hz6yTtupFlTX2FKGXWbWYWm3enR1/QjRpHzY5wotlQbtOpISTSDrb/wu7n4nNC8z
68/vVsVLYYAgA87E7tOnHYuB4fOtaieJszbiFI9ssmUvnbghxsmTJnU4r0FbUpr0
KQoSwr1CvVhmVCmtXTt4LL9+lxlO/eDKShye19GHcP2rCphZeyjzr9ct+pHZCKXT
P5mvbcDUCnvp8wy/miDSJfPQ42YRtO03VoexxEFlaUalTHfzxUIxbNrZ1bvJam6i
RcROVspcesug7kc6p0LmHvDG5RXiGVSEq2/W1N25dzYtk7eShXmbwwJH/1YHUPw6
PRAqQjJT8CDt7VYgo1krh5ErmlwgGNCaJNgUE4B8sTdhuzdaxsBiArrBnlj0xX/n
fzZbEWeCtObMK/bjGkzGO2941MGIvrYyBKvbR5mRHS1F2lmu8OpHLl9/B0hkt8vk
qm/TWv9GHHJHAkehJcPihnxs0hhZsTy3Gps/BMaZwvWk5ZM4jqfD7HBesKaak6RP
Du/b4bFttHHh1cTfS2MJG/3XnvtHl9A1Kz/n4m4nkz/MV7DWYMlZXhnskzNEs2mK
KyGD9FDoBPU621pU1UTbZi42rXjdL+LUKMFBAyuSgVN6SDRcBol722aZWE6IQLTO
RkZk/n7aSqaGWE70rXFFpcoiqhV7LVBLf84iH2UxDETQa0n9Tp8ux1VH8O3PqbKs
0Hh3ENh5cS2Vonc8g+2TW5QrCR6KglrO7SEt2iTZcpELYxCHiV5WXCdm7oG5zrxt
eMrVXkOF19VInsAOV93qYdYh/eq4vCZdeQAJr+Ji+0SGIWcfFalrFLBCWzliBTSw
IgNUr138zXOBAGkC3W7FgfF4HVoXwnCqda+h4pFnaqBqyJs4809xOJGKKGHSNlBG
uiJ2z/IszmHDqmXYHLu+mPeEhxvJPcO4mM7atR3JZHXMx7cFPaoNds9x9CKgYv22
3IDM8jSek542F2L28VbWzN01o+Xs2g6zILHvCZdMvBcFdObBa88kyARIK7Y6et8I
7VsspyrKAB49axm6fGBT/bs4qJZIIxI4gxWptyP58sqwtfsot4y8tcOPfSLiqjGq
i6qD4g1XgUr2kBndtp/NSN8Is6g+uZx/n4M5Kw9fXgLROkJJiyIVkpNOrw2cnEmd
kT96/BRlh8vHbVIfjrh2Dmoo0+206UFIMWOF7e0eWRFyfqfFgI2dUpM34Rcby2Ud
mbrLho3nRwe+FPtYIyD7E2SlATey2UIi26jhGfzr1UdefKxf+B+PSjpblFzGm+9i
xBWAxTJw823mP9fKxXx+8pCxg2MIdCtlNhxLfs03cth71gaFFBL+u1YxpVOziT/k
ufJ2J5Hd1QjNL6dcXAXnJTstVpNlSK6PNucsbqymQm3gU7wA5WAKqp7fH5WCh3KR
goZUQ7f+K96NqsR0rmM+njmRmhN+UelIwr35reNX0BUlpdVq5Ohvc8LbrRV+FLqL
gpAlOqSrpzDAtNgKKYn6i/q60t6+kXtKbb09+sVfxeclM3muVzJ1yUESFoXWUKW6
iu5G6joknmhFJpCcAvwHsG+v6wHSrknO6g5yDoLUxpA09zHt6kbtePL0wEuTRS/3
2o6cQUjyJU4qqhA5WI3128nCPw0LFJsBr2J+8T7xIj4bg7jr/majhTqrehl+hZLr
DJbozoVBJxhBlnPQvf5fzW7zFmc+94IVoa2weDVJJGINDm0pW2iulVLd/oyRgyEm
B59a5USgb/aLH+kHXABV4ymEaOTbfFZXthO4hxADq24taZOvozvQAdAwvWRsjh6/
frqYODzAXQTZW/8jWnGf3BUa+Vz+kuAamEeZ3/KAudy1im7Y324hrh8aHOFyUf5j
Ou6EG1WRBjYFlDhaqjuiOb3KBO45ZiIOyoqG/f3F3k5O/KCUrjwloWwMtfQxijyi
wR2f0YLBIQ4wVYftcdS2vf98a8tDYU6pGyIsMMC2b6i60BIa9zJ3hKM1GeU5AcYa
jvlCXDkwLlfSK/3nVSUXVyv0GoueNMvqYAdGdNg4sQERUGErbJsf8mwdHdeD62sb
2fxlYz44azb9lFejQBvzClU3f9zr02Cg4yyLCsHhkoV27uzww2zaoix6dNA8+cX0
CzqHBqffutGPHBhftKuLWUHoYwKq1zO8miBpgoUBEb9M4MQslKsp1UcqWSZbV7hn
rIiOxKPzyyOrg5cGZ7w7P3hgJbDIg7Lbn72HHzLPXhNfYYqvzWIV/g1FAhVfHw6T
341Ctri2Ha1oMfNL0az2349ZZBrifNJx8xicIRxrY5oPqCcSCksN081P5YDHtGpH
wvX4QKtFLNGdihsM/e8QX19bopoJt1zEb/URUb/A8Buo71BOgDAty9M3CkYUKSsf
LuwkDrEzY3Ey1E2mCJQ1s2FHupSU4YPGVf5W4td+Ivo5Y9zR6tzFLOZbY9m+NcFC
0Cv8kQ3wbugX1H7gtCWVQY2n3mU0MRGwfdUN+gal8Zcu0c0iGw7Y06qKMrelMuoh
SHP7mpByDy/Wd3CpGHwvNAKrrfWxq8sR2w5vNqQi6SYetkdgf5DJaw4Se+gyFd4l
+lx66iH2oG7jszklQEvigdo9ehqrIe6Zqy2IxRSwkloj34D4G6RIu/iZZfUXSTut
dMQyeJOWZoq34MeHo9gI4J5cdQogxu/nn/UsBMn68qTl8lQ+6/QFlD4+EpVK/afg
jogBcQnEsD1EqmVk5mwFOE95Aw2WUzgB7UwkLtS2EwOhuQMPEXuadZ9x1aRzW48y
azwrGYvYQ9Er6yh5Q+A8Jjkvv5y6aHmKX8tWrFT08yLgj7Zx9EWE/SrRTMQf4Qvj
vUFS6bwqdN/p83bf/6QEZmz7s6mh13W+vSJLbUdL2HAyDLSNld/Mc8WFbdQRn0Nu
p/zdqTPcfT01iNLYXzKDCUlFSu44sEH533jMjiPbDn1gJqpf+Cm3T0F+o/h1kHgc
fRKi6Ia63Ib4gRbViLVXMWFEGDI3eUjXgNH4riuEPLXyDLu2T71k2g0klC1CzGdC
LjrKaYRZnDOouyfUXA2eW+KhJjNFF4J2kBPCoSpNsKZeoxvu79f2uSGgQ3LW0wCx
WtBMhnVywNIhi94nqSf+ci6mi1ot9PigL8l+3XfMIC9+vYQAfHVpCaylHHjFvJiJ
Ok+kxMwiCVvuy9T36YD0VM/FQ376FfIZPEWTyuUpCeM8IBqxX03//zfJNfenQdHw
nXGQ0CC6ImdZrBhNmsKfDKNIikq5rGyIA3s5egYNB1vmUIobp1LN7MD37omf8MsL
0YL9qa8yhDT1orX2Q3jrJIyrhJtlKFkLCmz72jWRgPEncKnnaELa1hlm7z4F3AzJ
z6hatHjHikrXFN7eHgW0+/SSvdvYxlM9z86F1eaagm4qwabbZU81fDnqXvB/ov3/
OE6t3fESX5sf/TMCeZ8iLgLxRYoy4exitjukyj9Ut8hVAEtjMLArf3WnJDpoxACj
b5cVS+bsdALnOGZOHa2W8Rwtzd5d2Hf5NuapJICCVbL/bMrbuEht5vlxEoJUbr2j
X1JrBAhgBhrOWhdUC7bwe3S6SmamdTtdW/NOXM7z3ETwuKmZYqw3cFTJMjBM7UkH
IsfxzvodTkk1B2Pb1Cwman7Z+TrDhD8cwvqoK7dI+v7gMLC6on1kAARm6xiaOTDp
koh/VPsCzCmKNEneVdiYmipbFf5Nezb6P3vv1jwy6YPTnRauWfjN3EYq1VpHyt9w
/jALkDtCzu7c+owcJ0KuKMOwCw756A/nI4rL25lFKA5UwdXjSjodNwFxXZpqr4Jh
8utnC2YNn0SXwUiFQhLFE5sDrRX3JziTQaiZ/asyFVnJ+wLweP8EBgMBOWMGEHY4
AWXlWqFXJYyBy0oax8tU1TvJ0yx+34mHVmNDyB4MBFijPwvRNNEM0IgGVPIlkMfO
s80VcKLN/Cdn/zGJimffn3GxMlPt2ix2gWkWt6/2j58d5gpbuaQlRROb7HOyi2F9
J7xe2aU1+nhC81HEgAG+tLJDTib69bwDNDLgeR2uj8mPk6RUEsOhXq10Mm06dtru
8kw6RYYhY4lPy1fY8L63nnIigO9b3TRbRQl0TX2kMQsN30voNZVT4VLQ6aRzgiq1
IWf4BRTDrnf9xvNvtyvrG010CT+bt96hGdGXkb2Hfh9H+B9MSH4qr3MYZ3vcr7+I
zvvexVkdhu5xfZOlXanjeGzSt7ZK7GWhO1uHbHnMH/la2LMRoypGMxbkBxVP6UHu
fAvVibbSXiryF/6Y338DE9Ocf7em2L5zrIRTQ7pFjArW5iUlHjPoXiaZaKbiEPw8
D8SQAZlrGeyhSrvW33Fo96XfRQAnFc2tFq6gU4w/jpFl2WzPA/8DqXXC/UqBj5Dp
tvEQX4qaCBYNKmM/IiBSZdgi4nvFNUI6qvc5G6wl+sgxA+ykEpWvVTrFHBRM854S
xjNcDAW0700tzOkx1yNW8OPzIYDIqkE7BGjwTub9IBnis43WhPEhWA8NggK5oKC0
xNUNqHYW1NzVdQ5nct1QqChOcV4YSabaZQI6jAh5kKH7ZicZ95FU5nvn1xUaHj+b
1kaXvzSvQl/i9+aaPqbAJOdceEy1V4Iv/K4KIXtirwFQ7ZxIdKa6+X9TM8gm0KQ9
zojA9WgTSahfb3QZvzjg6t69eAkK0wutrmROj+FQ8qQ62WtQn9OpWNUuORE2M5IU
NWPJn2m2oYYm2sVTjHlsl+dWJjRi7EG21TXXHc1T1o/d2qxL4DHS8sq/k0opy9/c
cPFH/iC4htb4Y3dphRkODhJ4pWkyOKUmc6T38SiWnEQIfkQzCsq3PWXag07wSuZp
4u5xUHkad+hgoEOOfxij86AUQ8Jh8TZCs+a1ySjDRZV2/l6eZK5P/loRxF0aOall
G0hHiTpH4B0OWRZrdtmmRQFulBmGAIdUZ8WcKpck/m7OTvpuGG20FH0Q0g669yK2
hvrAFq/rXMMS8hNz/IqjXxhOMshMPV/AapS0mVwOb2hiTH8zEPl0KlUBEkRbA29x
+T1v48Ng/lRDmhtUPoJmAiB3MLraR9t4i+7tk0vjPJeqU+lJh9mp1XiZOMGzBHED
SEvkzO4cDrGRd4BFnLCLOt4EprMKn95yRtRmSINVLNmTwn9x+949Hycyfu2u4jll
MVbgIEbXbb8NO5fegzpRM17DRFtg3x0TQbQRFYQzYgJ5uHH8bK3nM+6kSertxX91
hff/HPRhhSx/rVu/ItgwgRSLTyAdk+RyCF0IdSTY3jYWe6p1l/wpt1E8Q1NMJnjq
mqm6d8g5wixoAPbcdkjFdJ64AejjXic39AMobW/XdvWH5zbAY0EVIzim+CtY2KV2
F9DzJPcH0rg7e7YF6BgOBlmN5BVDk1p3ijKjF+BtrpAyuV3MV1hzXc2oSmI7FT74
mLsQnsWgl9WZTxwNE9Pm2lpCx0wCl9DKi6LsY6uQF/KuoMhpH8l0TRjGZ3xO1QTt
ijnniZ+4ELc4iETEMrRgucLwnzz8HcJgMB15dxcx7MWmHjGIQx3mQQtdXtyacY/o
Y9+kHBSq5wU70yr5ILsw1gCZ/8KLoxOEVVl6azwPN3A+HTXs9lsjgChzqpOwmdaa
7aIns7bUQtFakLcnBu8GCkDnB5OrWx7/jeTiXMLH4s1FFLFK60HzSpMqs9jchGN5
BN3WBMR4fNALrK06taiIMIBMWNHtPJ07lU6zs5PP7mwYq0OcjqTmqDIlMme/lvso
uJcOSG/Ej/0aoFUi4phbM8i77Kpv3jhqwNBtmhbDHAHE2T69w7fT8Th4ZhXO/SKN
qHslLBgtQwrztGqbKlT9cxGJMuAyPDl+mbbT4CZHhrkT22OyOrnYZ+YdFFLdrGn9
QaZloJbBd8Zy4TSSTqXSOvF8ns5wvFqJv9n3zCgVNgHAK1nq0BquugingTh2YRXD
/r9vcgvmwM0u36vrfQW5E7WSODAG8oVip6erJQOXiMoYiWaI7RfDeS87hXe3z560
F+JViPGCAQo+yeJTHHav44cLrsv/PpQb51ZXSW30ty+eOBajr998mB3W2wWEooii
7yEmKUG+gazucjNMDLHH669IGx4irL5xaDxnY6VSizi0ia7JjTPttcf11o/5VMIV
fA95AknO0oOXFvyy2Ppw4st0UsR9h0pgn06z5XR1GXE9I6xcMJLj9YHgybTAoP/e
JCeqD89/KmKnL+WZCUez4exf/wCJqdfKf4pALNw2t0G683RCdzFBAlmgo9F9iBp/
XbH296msESm7WXoxv78Tp9Cl9vKBPOtolVXWTYY5ZiAhgGxjv7sv/1dqrNfetxB8
AjBqpaQzW/uzlmwLhHd37NOzPZAS44vANT+KxZImZE7AxAOtvspJiZuOPhS6J0Ss
jr3fO3Hu+PGK6YNS/btbb7FGWBXMzTyKtwATyD71oULHWksynZgWmXzT4bjptF1z
ErbKH/NyA/ygPKeTR6+VsVoAJo/hCvhudyfE2o2Bs6AQ501m+8EwuUMym3i0t5RC
1acYrrkU2jvC5lgw+T6gMr/Z9aU4FsiM+le2RDjALCwwACHdJn6S+k2GMeIh9YB6
LzBw9+btI8mkCPAozJSo05C9K/BVweaRdMXscvmwHy2OwCIO0XsbNG+4wfo36YYq
mlXF7KRgJV2cD7OtcF4tAgDN8Q62ieAoHVLeRi0+6/jdSMRgpl0zYs7mNjZNXkjt
Te6xSkRiCW5cDPUaTShTEx/OzcAashnRWXPGBPzPK4Y9lzMWxkJ5jdtilYrMmDrf
3Nq2p3docDR+cGmxhXPx7XLjJWi4biR3WnKFQQm4IYaIOBimLsAbmZHITdUFWhLV
cs40C7JUo8fvBX6PoYkrZljpktfp45Nl2wK11w1NYydtRzG+LcuGNF8+NfL0i8cw
Kj5klLRGKoLq5oxZsCFLS6WASg09s/w4d7Bl4kUfMjZt1l/IUF8Aa0mHaT473a/j
wfUJ/uLavaNJB4iaXIn2iwMUdsSjNC2clCaa/KXhsVq11nEOySMCjIq2YB1kgjGc
RcLEsTh4KGChHy3zqCc97GXThB76CPtJ0+IXI0l7LI659LY/uJJ/2ku0U6Qf++Ty
LHL811OX/ygRKepAkxRo6OA7ch7PspWWJFEa3o4CohoNoEvqmxFA5lNCcAdjA5d1
uWyAgTRId/I4poZxndDRJOC4qa1kXOP0NCs8P+jd2oZc4IoZDGHu7Ft56ZaLmtHG
lmNIPY+3Xs8FDSvgBySUljYlwEDHQ4UaxnN/zBxiCYf/4IEexPbWFWrbmjbAR61K
9euXWrhbYwNP6CBmsXPF6vmJ2fNiLA11lXRV4U2B40//Pq0DmlfKJkEXwCMxQ6i/
R3PzLyMm/KL6C3kjSY5tgk0qfO0+EZdyDzOJeAvNr2yqaEth4d+DgcnZXFEe/RAo
Cmg9ZRoh6gpvRedAl2Edfpiuiuod1pSzdyaPFmwpAV+l1gPuVFVAWcU8l8Om8i2A
oveyAOpa6czoh05KG0neQtY5wFIUU7089DyDJAkPzqXvpE9vbo421nGK6AGmqDzp
b5/ymuFdTV5EVLjUc2/QY4LAe5OPnYplZoY0uBctOm8w5oGf6zFBsWGaHOqTaovP
ItjJATs3aKonPAy4rajEz9PL1rh0chgUw/phjhP3SLwwMoS1JPx/Bn8ljQJ9QVK7
aPYsXCOWryWFlNUOSZjQKrvyQdmia82P35hi2R9152Y2fYJB+qQQEQ6ZzQ5fhqwm
nJChs/sGy4EVPr9gPEEGatI2z6RFgvbnjvmFsJueKd/dgCmS9YAGknIW4fHt5pmj
a4j9uK6kQ8pwZ+anjBwk9Wf/cG1FJXSOrz/Lw2hf3a0vKke0R6ESLPXLW0imO+X3
/92N34tHsnSmKojjJXcU++ty/tudeKtVgeBpCbijpELC7azCGNWyk9TszYvZ+4un
XJt9K6NnNJ2BXzFEaRGebEVnu0+geEpsma9gtSrQfRFTjo1x+KfnLEuA0Rps5XXI
tm4QJlQ/rZuyY+lv0iJ+H6D2RExPvoFIlsQf97e8RHIPCEyvIaq2zvHz0UzRTGpO
+nS7wT6IdHb01NT9HGra4qnKrKaz+8eDgmWzB/6esai+iEZuTmtxXLnM+sm+Qr+R
8oxUmd6QiHH1LWRu+y0NRZxO9w+Z44Y2EQG++3QOXfyZ4DTPIo5vWbZZYZIFNrsT
IPsGWV+IOZnmdY6jv1TX13Kf7fDN18fzI/SfFSIR9DM71Wh9VctFUVm6dcGb3qx6
hmafljbEUR97FT7Qygv4tFDaKdxuA3phVZBru8Kicc82nhOMPJEn6FmIHUxq2N7N
2JRIENZfGdbMHNnDBzN7jp6/BOCVCNLuOJKCHfXM33kdTrHfcWl9Kbako4NHlCT4
69UHKbCUU0idBmoZ5h29MgXABg6RIFkAlbrXeKhvtB30UmVxu/mkjlr+OE07LP4z
v6lMeRUqW3G99A4InGujjbMiagiHEKIVGzOw0mQFLqiuMjBRh3gZQaUSYV8nGKw7
rh2afK4l/Cv9YYFBfpM048WpgcnlaO9ngwFJjn9Dah0Swr8XpaUw/6qGTb6RMTSe
0/GCYdHOCNGGaja7QV3rzNB7+vmdLcXz54TyF9wtiV2X0kYbUB5h5JuwuIf9A7Yg
N5KfkRCwEdaC1Dkd5q+xI+mZZa3Pu50/d7I9kKFFceQaHp+uBGH6DLhV8CkaOiZT
8+C4S0EO2Bp1GtNy/5ALc+3tVApNKYgg3T3dZmPGJvPTN4EuqCn+ZvlbGzb6U9jH
8rpuGg3XApplnIpnkLzC4jNqoR9RGJJIhQcNKENdtBh9IZdSf27F+8cZIC1caJTS
TK/RLFJ2svGsSGX09vns9Wm9oMc9cIcue+dcOw+1zEhBRHSah4v6uAfqyd/TBbfX
97WcgfZOe+/a9uj0Ui/ZMUppHgvunbVQI8asZgUNYE/15ltV4XGMxeyVVDEVF9ni
XTCiLzZWhgdTwmMealt5hf/+QBDsuH9XsLtxOcdY0SJQlBw2x2vfFPje0J5YvbZ6
kcQRjxLLm17o3y+216aUaCxeji7qVSF2sTL0LRK1bgEDkNZ8ZWPu3VjKQpkD1UgV
GCWBb4+IB3waauUKYXFtpsg+P57X0RSkkBRQ9F+MZDrLpWnbwp7CvMSpdo+kaLEU
9F1Tf0zqdiyZiVKQUoo2SKBTh4ZhExCgFLnyUeSS+qu/+SjZUVOPTmgr3rQ5hvMl
YyP8Or+9nwAn6Yl/Mv24/juZFQsmWwYLMvksfm2zl0atP0J0PY0beFtJd+LcL08r
siWsx9j0B9PcISEXghJDKPJDlABiydxPopDOvJ7RXNWH478xej1ez26W9GiYQ/Mf
LdZ9orFRHqhnE0RhmDCzkDG1bDKzd7wslPVbcQmIuRWQFKBf8t5oQ4CliZ4scTxv
CMeLlzYNhidQQ65U89iMmK7IeEu96fvDrp1OcNh/OBYhoyiwj6Yj3ayxgftqG8OO
5DBPTRaNAGjZaykZJ+AJs89Vij40zjBpL4R3Kwg8ToZajXVAPLMLzT6jYOfbxLJJ
19AYVfHR9aO/CzXfE9DOuNKwWJDGdo2ERWAtSl051DFGiIQcF9gi7TJNuO4TZ9V+
xCaV44jpUDgAf2nz8+RmSvh+GGt7ETbW2Q3xQ5p1dK+EVBcEEK17Uv4XC/zXG/nd
8XCVZ8pC9aqpshBSTxExKvIySwbeFzOgK2q5NR2isqrN2lpv98CzY0mVQPbc4Off
G7H2XXisw70XhYRSSQtI0f7wQl/WjxwiTs9QHWa+81nzihqpDXpzGy9wILDfUFuH
VegYU66jwOwAWTQqsLJ/+eIvLvj0Z2Kq/82D9rYUTedIt2pkSYpO8N8gMloBgNQM
HdE0X6ahMDCBebesUS53evbhDP7CuVlQv3almcTxYuoecxG5zYxOGh7zPFcGzomj
JuqkpC8fpjg5eB/n5dks9h1C8TxRhKJW+nf9b4Hw/tNN98VrGUrUpL3SEQqDefrG
8BE9pRn9YmQYMHSYfNH5sY7CNhZtGWDk/VjfdU2G+bSZZRPXdFW6ujbZoDjsMryL
mhSbtyCrge7KxB66xVo5C/RHGo31ZY0Uuqg1e1Yv6YX2WsnZH9FQ6d+Ie3KyPizj
T/dzGZojH7qGHJtiSIb+NY9hkl3TFSDWbRydyfphavtKCXx8shY5VKL0ldMHbojE
/flLuBNREjV62+Ol5teRqcDqtUM+EV24MGe9PQo/HUmUC9kJhp6wRb/dm3oF1kZb
Os+Z07yaxFh4kj856w/rkE+Q8u7mTx6F2MPmFPhUZcQndA66raR5jrHvVmqmgKip
nPSAo4V6U0R49Zdqc3Rx8oYFKzL86JXK4BGG42manmXgFB0fnK9f4DnH5moimYDE
UuBIE049+/Buip/+ostan1yEsyU2DMhfVA4mzxK1SUIh38+di+1/k9XPFoxB54gz
DTpYwuth44DbM6orY1DeQ7Yu31xNmaGcT71GBzh/4c3APh9ZKf5/oIhH4LRQsZPU
y9cQr7s27ZRTtqHpSbNSpdNOoRqVKS7N7JJ4WV8hueNYYerM55/IJVYC9gRCjSdP
+6ekaz5H15/BoEd0lMFXRqFN1PYgym1mAvnUNLPjPFGHezwP+vdzrSPGBnxz5P7K
DhuNzMDdx4ttZQna+zPRHpkZ5B6okZcsqw8wXQn32eONwrI7aEV+AMguPd9TMXOM
3j4atHVJwmsDAWOnusnwSKV60HV2FHoDd7rM2+GXFHJ11lH3pO9KTIaWuI77X62o
aDZjdlaKDyY3RYo/IOaQnW5u+Uy0NBzFgFAVdpd1PqTgU04KmRxTf8HwWOFWdDe4
wrr/4Azi2omIkw6UEIE++CwQRdWLlulCLBGfSx6nuKWZiW5y7g8+uRHj3KUw9rmV
4ikm/7njDxQ+zx5a0qWyEa6DHIw6xIi3P6jzecbe3dqVozWfvnT3toX9qJ1mOINg
3CLyW0dwMwVbdqyLQI0NiK5T6wBHNANUJ/T8qb7UtiQlhADTeJRvy3yC2wHWTuKM
DuPO5kcbHjaIylvFhHfc+PDDWJk3xEdU/YFnavF/5mtHJB4wfhwDcgVqVxIWKzC1
1b4bc8rHIMk9jWxrNtMFES7Et+ELzchAUCZAV+60w+mqr8dJWFaEyNkiGg+s0fkn
y+Umb1eLs9gInwX9IAVwTEh5hhVCqNj1Mqk7g6H2jK99RvjJG9wgfjXsnW7+wsOA
k1mLexzAZG2A+/wosJFX8PQhgBpH9AM8e+S/TljroYDduKC0Wmi4c9DiEJipEOEt
C10jfy6iyMOIv9xUjxcoPJ61Q2kGGL07ffXASLWECP6TLF6p1RzZpXPYHngNI7Zv
fypHfgko6zH8xVI+B/l4rGRTs0bLl591i1jXBCGWAVw2NmdLeuzaij0clo0qddil
btaj7jHV1Ja70oYoyncZRY7AiZXjgZzaDA2L93lbsrTz+LKB6KYmURdsbKpjfEzq
Natf4rmouSBD8EYxrPnpJHkn3qmdJwxLpgn1SjBROjbya/7EnWeyOY1+7VhSkVne
9ls/CVaNq2xKxnnRybOvdzqikev+dZN9kwC3bbTc/khRzpaMhrSfYOA3Btf8d0qc
yamxtP21NlxZGa56sMOst1LWvwVt93ZY5Mh1xCyS2NmV4L7wbE2H0Lw09m+1HV8Q
DEhsi+v8QeYU+35Dn+UWDjQVOkKzkSFwNOvQoOMxCPdFTYN8HAD/DDeFcIEIc/q8
5D2kksJQIDBzIiPLlAHF/EhJCAaUS4FeuGWCwCxkE07HbCUkR/Vvom/UdE0oMovb
2D/zeF+x6tMTns+z07Aqa3u3cqHPYutiHMK7/w67TEoLyf2I1PC+oajLduWQ5vOo
5wBUjECCd1ypIoEt3L91wKMlqB7ihl2vFtezDkvRUoptpaIYx3IzDc/AQgYzZRHv
/j+z/v8nuO2/VtRlDnA2c453oNYEMumB+Q/D8Inq2ySu3DInUqSVSBAgIz1yHKTu
/ACtFKSFa/Fv7WrTT/E+ykEuYmWH59QWQ1xgIkJKkfvBW+P1sxFnHpASTkLqlLEe
RVt+NBJjhqRpZd46ODZIWDP/H2eQG5cr1UvSfAoU8VagcIa33QpKF0OsP0ko1h6k
/+EOeibjTeSrFvy71XCnoEAXIcheWnGDomTTZEU8uYpgn3XQUOEU0DPJ2ivgAfGp
J5faLRJGrSFL2BAfYimUe5yxZP7N8a+8FhAqXdj8OwfsvyvQMSaBbLXuoSTD+rsD
d62YGxLOlxFiWjcKBwuQS/MN7x6PfJfdeSAuflvD0AUHAHrj1GxAY4xHXF8Y8JC3
Ty6ci0dtfVO9CoCyDBAgT4bFNgnTcxJiOIIb3Iv6dejuyuYMcCKNgTjtALTwsKAD
4M+XnUzwrBH6zHzWR+o9dEpTjf9bdLNbGwpRKII4iUjRQW5YHRZ/YnDFJL954lUs
rF37kUWdS3u4H8DqPFnDgj5+zIPNSy6sU5/8dTtip6HM/nk4wTBoP+b1l+3uZKj5
JY8MpcA6tEZoaxBD2fZ7/spz+K29wBFPZYGiv65N54J+uhhWpwUHmZT1UQE3TOE+
ws6gtXbHFYXMdd+DEh00FhWdhzh4d7m7rdwi8doXXvGQAgqJL22W2sfi1yp9LLOF
roOQHlVLSSYU1Ju5+SHKIjblznu718/5qJ7n4GAHxXtii9R3OuOzTtUkRghaqUO5
LNvn5ryu7wtg6ZPCm9Qk1CeoWQh40fwuNG8KxrPFWFHFQqBj8SU4qs0ybSOJVucl
C2EGAP3wR0XGjM/t63UKnmEEa1oRiRNqZwLQcQWMQ8KGFPbYUbrf7xOrRz7nqUw+
kA8ayUr7QgW5bEyWEi4bYZLRkW5I+Pmn2GK0PK00ZC4mEj/O7v7ttM5sSjIxYg26
qoT5XOfyUwouL86viV+fQydJDIjCWgYMvd4/wYqbX8hLs1ZLjaO2ZWCImxqbX3T+
T91AxdR33MeGeHIw5aeZJ1XK7nSweUt0BekWSrKI3oN9pg07dNap2SiBtxeGv2eQ
zjoCdTX9D1gzW4LZgbTHSUYDIZT0HVrQQjOT2m/GRG6MYFSyCMOFY6l4N5rbaSof
khXTHkACVacUwvl0s0/6w+KG1lZYVxa4VXm78iEfOMz4dzltW9s/EfQ8XipaTGny
kFeDp9mX0TU3JSRlQxqBQpm3zB4pUWjzqx9y0eVTEq9Cs4Wivkf7+SJ+6vEOz/0q
iwPsstzBKgnNiWVBy9bZuGw/j/b8W/fYvndGzbXguqjLS+cto7122H0zvfI7LyoP
ox6XtO5a1DEp1iN520nEh1n+o74XzNTJNYlZsLrUdP7QiD1M0tt7f5PaDyYHKrFj
5At610p7iAWhiKj9KjnJHEPJGOta1yJlB6k6h+kKeYmclUcyV2EWgfaiTnpZlpOV
0/TvI+7L4X43qGLDcaVxMNy0txCfYThG3PrNWc+jPXCwj+R3LcCVV3N+2asUeUI8
thKLVL3zZB5ZlKwyHENh0q6CW9QiX4499LRymitFziXqB4tFHVpG+FDZZe1skI1k
YtTtlk/RyrUfT497pkvp71JvYOEyTWk2hljm1QwfMalGp6/Xm7EdNPug20Z4ldA3
4armrKjaqREKKd0AkDGnDXMOTEvjLVeFoh5Pso4mxcQj0u7f7Fsnm19XQtb6EnNA
DauH1lGMUPU1UuZ974n2dxKT0dhlEyoy0vAReaBHL4z1To9wzAT3qnBPa7Fqt3WC
UIQSr7VgzRRtFKHZZxb+aTYGZs8iGhZ9hvSvwVB7M3aavnNMxkr2jiI1POnfS7sk
W3erA9Z73YNODJjdNIuEhnfc0hBPy9k8MgxWU6gCNElod9mSquaHmokiWF3QWeJL
vOLYt1Ts440DDq2wf2VaXmn1W29wQ8UEPCnl6dWHJKS+st4kWzBPvT4rK0FbKUK8
cMIXvV9nVWs/cf0T8jDfLiY/FjkYjxGe+KdRhiDjtenTe1Jf/n6PXiJfLZWF7+ry
ZhJlU5c0sxFP3vC+vQFu1QQafYMRZgW+BT/bF7YO9hFR/QIuq7rnrIQBTgp/dVSB
lqHJi3JvYLiCigi7DQuZiqXOgvd5Lb7zqsB1CPoeim3UkqehuMfJ1BHDo2wCuw6C
h9GCtLSXiO6+46zErLgiOlSJWYO8JxYAdWajSf+wfQ7uACMpO8V10j9bRY3fuRtR
u/dja4v/3aVL0TYnAQ0M6JCcqCIKMqxkTbqZbFHNB7sbWWCPL2m06vbc4ef+0OJg
63+igEOqB9CarsNKVPMjJk0A7J138EKbSufJE/QQ8EATaUYPKI6gVWBY8w7ROnFX
d4EQv9QXDzOIjdgTvN6W4Vn+Bhh9TJ7NA3uKOOtUjMhBOl/aDz5cd9pmbmb7nU5b
rKf8hcCmpyXXIqU8Dsqy3LMqXebyqguE0JLGS+iu0otnk1JRVw4v/Ie4CHnAiNxV
2a98eEsMnviqrLOt4LLlP1X9DnlKVjdCFV2tXcO5ko0vEtEzMaYoGYvakmiySHZ9
LmFGInusVYKvY9PcgV9Qrod6Bibr4fI7mCZF4rJCw0aGhzROYadAFvxZO1h55YDY
/1KcA+d4AMd9gbxB1VJU5cMqEWw6OjbXHFY8vhD7D3TvSfMqcN0kMJSF4rL6Ealr
b/b7V8BFkC2nj610Vioba9cISwM8hF7dqMPcxXZSwDchqJgk28E0Zy7HL0gLN2zR
iQgS1B42yLVzGOgtn0ibSVQWQ1GEWux5yHGd+Zu4VOc/d/tt7+HR2xYmd7G8ooN2
ZPEnGTT0rWoXfvHbeNXCsDCj3VtXaONtX72/E/vy4ABodTUknX0sRf2IJgEaaqex
NlT5uAISg2RGXQ7lyNkvXlDuF2cA7cdA1GDlByEDr+LCWMPcG4D5yBBrRyIB5Gbe
JBGRXfVH1X9RacOnEVvqZ09yUZOwFeVLBbTE8Ei4oQpjSgeAhaUyncJUlOgU2B+A
LMZqfy2sEvN+C1YgFy+8sS1SrQSpsI5IaV4NK3JDgCWirEjAvOixx/tahnkCAYKB
3WG0NTFpAbHsS5rNTdwDkQZxEECwCNHNOWRa3G1IGUjQieu2QLn+ld90qjokrz1R
31qCBxJXICTTH/Nr1RHtpC8WeY+4zXxu9b6cTYa7jnkzaWsWpHj49Q5woRR3k3S7
WjdsHQSeIbQcoR/gYsyQiodEYlso53Mcty8ED5yiimgy0Rr/DejLb22cg+70hXsz
DNpTX0RSCWh1H4OV7ephYKgsK9cpNP+K3oOTiU8/bByQ9EYATuGJ/g3wOf6nFLaN
dp0WxTnt1ERLK69XhtFy5GmMPSl73VBvJru2IkJNchNi2LjEXQeoEMziPllTFXcE
mgPRwGN7MVnCB1/hfdpSvztegqnb3JRDz8uxPhAClWrtOAjiETvUcmPrJKYSU+5g
XJndgvCYVmogQTLoaZvrHRAz+golOFTWJhJLa8VRjz+9Fd0+W6d7efw779jeVYbN
79cyFmiwDV1viIGaM2mQwqwOlahgaJPsavmp4bl8TlZmKzOe/O1OiV8f2mM6lCnP
bfcBEZ9/NClqgXu/Gwa15M01+c/UjFwVAOKHnmN12ouU4YB924AYowQgiLsIHaT0
/sw6ixdxcpjN0VOzTuf21NwS6GruaxBB9RqXXvcEsGceawWiWB3dUD7U1iblaKkH
ScZ4huLMgnDF5F0JV0vMly5Jqdb2KOgvwzYasaPnsJGmi7/b9nAPldx8ywrsqmKt
vvdcoXMGj6f5SD0yXQm/kVIZUQoUQiwUlxs3pQlGjURa3JuSgH91tEH19x/R5qW9
HnfKunreRtYJw9WF98PfppeLXXgGAy2d7QZnlgcqtFzT0fiZvj0UmurT3zcwmq24
rYsDaz4ahN7FnGvb/Mlzu+zQ1syoVAKyBhCDQ0B+1XA004XtKhEhb21NNn8zaWUA
KgjlX9KFI5zsGmWx9c1+BrO0vKGB7+dWweSsL6b9Wh3OP+zvQcjTdlJZc3JnE8m6
3ypZB7LKPr9NLkVwCMcTo35PZLGr72/EuPJWrBJNEWUb19JKuULkUlgXd4Tr8bCH
gj0uI3zBWbWKIJTT/Ti4cVNGy0IH6bY5X0qFgxSne+b7BH1I3fYRSNqchMaTu1ZC
DSqB0vgbz2czcU9oAX9zcXxKlramwR6DlgRFc8DJC2yOnSfSOkElsamwYBOsuI3I
3Bne5q70tEyeTaTVf3OHhHYsQKt+EeI8jDD3fote14pcOiuaLtxqRKm1z3WOoZ+B
jdLYZLapgPaq6YmJFyPqpjJDZEo5f+0pyTf8/OPBHNZS8eYIj1AnIWEtOMTEJxeN
7SHFykOP3tN/aVEDsoaNJNTpIG0VocX8lfa4QZ1x8fBuP6OWpqTEu972hts+7/jv
0b5QqWNqq+a2JsNwYhPfTRxqN2Qju66AJ9pxwI3v8so37wAfQK5OifRGkxC9rnHF
l3qKWJ4NqujsWiSMuAJheVVeUYPTEGyKU4f3DwOnmu6O0xvpx/XWS8gvsFkjz1mb
M2CZqKKwdyARcQmr1nSuwyF/1ox/wgWY9Ikh6gHTyAvODELxfxawvh582XlHTS2Z
nzycbB+S/INnh4yjoyfufty7hvuYLxJZ25rNYY+cGO8E7uskWENFxUNaWCp8P82Q
end+1WSCrieg8EgY2r+FBYMI8BoCVNYSNNLpqP9vqYty2wkv20AKLEWFA+M6+g1V
bR+x2v2yxCvTAMyiSTZKyMgWzHxp2LcINTf4TXErZjk7kprekwSV5l44Kr7UUCY9
/u6bP0ud147HmyK3kwSMOit3ppieVEk4xtvIivkz+D4d0F94ZQ6bSg4b+uxMGb5V
AI6apk1Tr+qBhnByWkA3zX3ab13D6QBCu9pL+lCJa+J1DzvjX/sE1Pl2fTyFL0Vp
CD1d4BnEXpHaYDoHi2mjvvBBN3CtedehUWJOdW2LzjecuuTMpe68U2nP4JLpNxc4
1U/NekDGExm+Jj6wmtxYhamB0xK4D6Zp4UaoDoqehcDqRBSgJrAt/BRIC0qwUC2M
wYwFqd92mmK0Kyq9vTSEiX+CgkY9u++CIu8Y4SIM7JPxG/x6f7+Tpfpvtp1hfkXn
v4pmabnY0jLPcAj9NgjDqVxsyaNKKtpRQRHv1rRWRXaF9whsrfqkDEqmjLUmfpXS
mo9NyHJ+bBNWVsT/gh7+wW3Mc5om8KP4507cehkddsyZyUAa/fe2JqzOQ+AkBJ8B
ephapZuj++kU4q0oTgEF9wwI/+4sOiUisvbeUQ2plkfBjEmyJ/kywmk2/0FE4uyG
In5ey+XPATwiLDkH2J563ai8c1doZZZDUjEmIyoUMNArzpxuELx2R9Gn3+5AE6pI
+1Zw8e4BNODiWH2i7zI/2PQqiJYNZ+P7jSerDmCDowiUYfvp0ZBF1VJ4VagOjHFv
ADgv0eDSkdwARPT6jUhMesK/t2CyVlxFOpxnL8YFjjaF64ZDf7PNPaw/PtaAU/DS
voEPW9YdIrRE/rF72o1aYGxiRcKhiiaCXneWqAm8Sn7rszZF3iitWvWiwZDiwr67
xwoblc4u3m1jzB0b6w8OWDbFqoFfMzE/pvs5B/53eh2M3x+sUlQc/GrG4SS44U8c
vMuZQBZTwLAy+gNqINBZSY0kn1gchCv/6BtnAKLWQZqpuShWZmBpDBCYg1Uw89hG
nSssgmrSAF5K+UwnB9nkS6euYCYXjJupc1fB+SwaNSc1mIToAGR6zmgLY7xRbbVD
ywJ/trsRPVhUMnbI1eP4VE35hypNBrAymGEEmWVEZAqbUn4q6gVmhpgMPsggx/NM
IDvLONNj/mPBiNq0+s7G4MDQrTbEYjWwVtB7tqlzJZPdoZHIdkP0vETwNJBS4i/G
3q+nAzuUMM0jkyvqpiG4XWLn/SOaTpP53VTriz2wU9Cva9y5mvV0Y2Lkkoaf/GVL
/gaaY0cGQ7bCeVaB2QRPhOP4vAIoJrYeE/MDYli4Ev5O9GubIfz4mA3S31CdnO3j
qZf/7eDDVNpLkcVg0Ig2YGHaKz9lWtHqWy80j+V7TCCsUY2tL63CPnKceptHI1Lz
INqkW9PD0/eTvO47k8LLlNv9hcyhQBBihXMz3gf46OF7EC6Yn+DCTQ9Dz1UBGJi4
JcZmW3/uqIPgxDG2hnSMPMHRaHu5UlcHcttqXjdsHCrgJhJrFtaK8+fNumlO1kSv
Dtx1lRstXh6hpbWO1v/JPZs1iiFCLcXROhPOzTdvG5LLAJP85KZevAQlXxI0qyfO
dc7Q/8M9XdWQV7FOnGcuYQsXo5hoTb4xfQRIcbjHQAqgXVmv4AkHbHs1N8HNqBG9
T7BeJnHbJhT79FyTY2MXw0XULQVQacLCOWv0f8ckl68C5LjBmKqBQw0OJ0wJxcS0
qx/UBsOzcqE8X/fRf4CkwFKo4l5Z2j0mx12WaszlR0wNC+GMA1CDhZr1WS+aKx6E
EDnR3ZegsVKxZWhVb5WM55SkFx8fDeIwI9Hx9YqI9Sv2EvcMfWFrxAMUSwd5m/Eq
gQdzDFgRAxbFXHSodDnry8TYipkt3M/8oBJFfvYvjmxetqNM+g7XFkpUOnfGwtAU
z6qJgWToXUi0ISZYF8sP3KJtDIHUwwq386OXTTYgFZjoSpHlnMQ8Oue5iqnLl7hO
XSrS1/JGixlrW4w/ASmwSW1uQ8UTPg+C2HN4QI0XjHxMEx7UnVYRXvWLgMEjx0fy
sJkUDrRu8/IjAH79k69qyMFggLhrdjc9QV/WRJFSOb2wFdhXdYLShV6FHkLVVKbp
/QrRlZGxqt4p/JYsTWohlBhFV/wyfkgPhFYF8ZuqgDkNksnp6wE87MKUNnXkE8No
ymAtkYMpIXveM1Sda/s9uA7K78eMJzwV3V3ZnpUEInZ80w6vIV1ekJRY9lU0+LSw
ooKfEhxa32PxVELlPoQrvfIogT3YmUMNBzQfdE7WFEV2d80FB5o2i1WtoebRyymj
NMfwAEVMQ4+dX8dd0Cck46Zic23QuD4I2T2vbxXTzMaYYOoCgUAy/sOcS7o3cLol
urDhaKo5CskMHWJNPvDx1VaUgp8lq5IIe70+1UgRxgfmKBZC9fZj7JkcW7uikGmL
lW9XIQ5bn/8CocsKq5sAlsCL7K2Ce1thnnVAMPNb09sxehzm8sNmdnw1RKl8CKNc
xvpFwBx/dIevK4dPjJuYt2RtephF5roimjCpadAfLQdmyH/weIgacNvKE1ld2H+q
+SV8SnyrcVfzMqUFO7ju7aSGVSuHV9AfHZ+MHjj+iaqhpPBLya3a+Odeh5uEa2jT
B7PON9TATILUFlCVNIwPZpsKCU8hMLVo4DcfN2JDzMlJuEo/ooKG4/wE/HAboq4s
5F1WSLwIW0zKvtnq1Diuh4sXbzrQzraXZFxOvhPx+iebCxNMSAgkfA4RI3+eZnhj
70zRG9ywhJnZTSrNydRrJAHsINSHNmac2D2Og/MPMJW5R86as5+M+xcGhoPYzJJ1
5Z9XJ/SNgJvzh4b9UCmm+6GEAD3YVpgVHXr38fAdZ+09rPaMd8zA1OcAL/iGNBl3
1cFvTfyKElEkvkQMClM/zWzPKykKGuY1eB0ifqU4H6MJliZP67Hd38u7lVBcErG+
hS0avO3S1g0G7aVJ3o6guq2EAmZXUOvB91PC/9ESkfo5r0cUmx+s7sPT1EFbvQh2
1dsuv5yc/RKYXMBQsgZNz+vpGw/B4sLBOWT7Pjkb5QOfztzaVNLd2H98tFTB8Afp
baK45TLt19s6dpupw2Cdzf3iXduWibn17GxaOxXInfeJUKFgbGX/Q3Zi+XGzs+Pp
bxnquxsgTHXrxfjUkP8+VT5Edra56ux2cNNAXA/jVof06sTkK70Epm8W9DoMzp8h
2+bTcc8q3aoLlt0AlbTrfreyPeTFQipqvin2c101TuJ/Z9olYp6HEufbdoQotzcT
UEVA5X+eV7zfjQIDKsTVjIF6/xzVOOJlu4CzAdKJOuoc4hcWfKWz9g7u6aVg9Gss
NIMP0GIsd/y8B2Owna/qIeqQTkqL7w1MZjURqBj/JJ4T9KZbcfizSzPRDQLJFaIj
rpuJTaYpRlDMPfBMgbAx7iXzUOhylUh9VSAmy3SSqgHTfIROybIJfJ5cP6T0kSEI
0L0xqHxab/dzrGRyIZizDJppeigvLEbGWLzyjCxpiIBas0LP9D7G0AXf2J6Dx/VR
vWEWHwrGublfEBQmrYlyg+0wEgQ9TgBoZWg9tGkVdhcs5YRnkq9OzRGC1GzGKukK
g6/oMb3trUh3dK6H5IxIzzDJFfDApJAm6gGQu0xuvSzQEQbjWdXe7QAXJF43MhPs
WR8RY17nKO+9ByT0Cn+/LQr9kd+Ljr4jSv+mVDyGts/t1FIUqRHh+sCpS7YH5hi5
eumAkHXCZCrRSvGQIoOhyxCGPjDHLdiscA0vR6g6OGcMPf1sZDDaoFMuLLZutoUE
wAbIqawjEEiuxXFXxiCbPx8RvSuoJpzIDt7m2Dk32iMmxEFCJNO/+Fouz2ZjpTis
KFqS+wClL8jmxDgKvyMPs22p6Yj3Az1RJ/DXjQtUsDaRE9Bzk2Nvx1krTkMsQU7E
og3wl11tfQ0E5s2ImcWL5h41UkeQOJDIyKQk7VyCYlNhCJLWiGxg6fIbxRTHfnEw
cMdvM0tKiXFozVDrpV58VF58sf2bMqx6r9lKsduO0rY8d5ohQF+Fxn+ag4X/lQU5
FjBIyK0fOFpgsu+UDYCIk4N1a9ggTksT/Ne6QXjPMFvuwhmwK50vHaAcdNjjbeGT
WxA06xsnB99ay0DJM38cQkPyB+7sjhN6GBEiWmaioyabpJd9CVi3WvLt3PTps+ab
0uk0nHaEapI5HeMrgn3kCwsH095K06qwnahA5S1sLK4nBhYKLlbDBlmUjCBcjRBM
auoa+cKSSrmoapDuipjn1WtAIfXOCGqjPRUsFaafZHzfG6hIH2kETAji2DyoN4M0
AEMLLXNWxiACTb5EBAzxsK9eXSFv1NyM/ovVz4BE0Uzz6EegBRxHI5JciHQdVzZ6
Z/tTeWFjg6llnlGOyAEDv0z3AQyTV0hZwzD3Qtt5KR8++e2m6b2VMfpBHT2H0zl+
hktXHMnuoaohT/OXblVAa3VD2jAqlKGQj7LUezop3QTs5xlrqaHXBPs6CJWET5+D
MjY62fBwdVIOSgba04zQi2VfGktJQgC089g4VAzQPx4f/L07A9++1qflJAoikPde
g/5+etip7zoNM9VbwWPHEMC1zPn93Wm1fFVih6S4jKnOQQvOA/sJHGguZRzywig9
/dq0Jad+NLTSB1AriQqkFnkTwvkHIbtVjUKSmbekMEwTPgFh7r8LBTFj7K7OlhEf
2nO7V7b9XTBjo0m2ii9fieukoJ80Y+vw8yWpR1eXlESt3liwZ8mqNUXMuxY/NVck
kS18oqoabNByEtWXDitdNbC1J5tCRy4PmPlecM32nWJKIFD3zFegFSY2DpepgjW5
lZONOCkDSr34IM+RgoUimJTEd90L27MeHF01c4pbljPjqdOOIaQ+EEwaj1aWImBu
Zve4YgUj6e9Ev3NlbR2Xi3JaAqTww8AQA7eECJ/nrJ8quYP01Xuf8w/yr/uTo7tS
COsJsHtgpqgRg44hY3cgzw7EJSP+CFQ30IcW9qFpGIxk/GKISX5ahgzZuKXD0Pk6
ensaFIt9oUz2VJO/XGRDnwQfxQ20jYWn/rAisPEWDIkZHNyUN1z/bOgbgcVESyZD
l+kIFM5IRF6n9Gs4zEX5k2V911l3bxarQDcRKnEJtFoqYd/0Z2hsztkFOoIDiwG5
SmF97EnxbKNpI4ZX50UG8DYmOPiFEVHvKM/SwjoQeu4wRelIwAFxNPEZRQyR4vCJ
iseLTH9YAnKxizCkhB8O4BaAfgnpN42XcQMxyZ40zXyS+cIzCqHebJmwkuNDYJRP
W6sNYrH0matv5YOz6sBzCJVc0/lnvP3qnp56fcZQiHygR9OHbRHk6hnoPsZ31NJo
cTeRDMrpr9ZEXuYIum+wpPckW4+g72Ft0O0IghvVIjMh6zOloWK7Lat0yoU+VAON
E14fH2EnHZaqzkiNjIJh0dy8cBJXW/VAWeQkXfz3MrJ0Yi7Lfz6316bw+UZ0KUL8
kWWoB+cQFqsQ2EedDS9d9Satgv8pfSHGQR+L7tmKZSaVfTXbdzdAdnv0dVB3tKqn
QRu761dn1EBwrwtUasomJlepQoEBC9jOrX5U9eaOkXmMiLpFLiJK07x9Ruy8qXII
h/ypSYJ8DUt4Os0wggC2Y3jPBvwzOTeLvNczw18EZOsAKQdGW8a5+Dx+9LnwtDE2
pJ2YdjA7fhFtc7rgWP0uFr1swhnfsCLTVSmchKCRLxVPAEd0LUFiH8Wv2m01YxXY
L8/07r/WxTeBYPFS+XoORR7sG4TLqyTld+OHLEsYbpW6LDkUyFnAa8ekSwNUcz3s
opXQ2+0F4oD/EJoQDMqFOR15FLnhmr4RgECeDAfNoBsSGMRxbN1ChYkbV5rdkyZ4
LupFPmPQrZb1gwCIHa15qVzFxqie6i/9BzpkgCcMFZLG5RdpKvoXI1TZy+gZFzg9
Uv8gYzhSqMZAHVlKnHLFCeiQ1islT4Q6+lShDLnZeSPkmd8iTp9Ga3qQD9sDpouz
kxSkSQGgxiu6GOoeuE2t10lHwuIpFnw5NB/CNz29NnWrPsXznOuce3CZ1hms70eD
E95FaeWfelDE4KWwuLcBaCv5jL1MKIT8lispLYHnYFW96taUFT14CbMqRf/2sKvq
L6OO7oBXzYn/qkPUwoSUg6gM1zWe0FdEGKN8HY7fYIaemMdHQstQR7ASgAljesfF
4EVpYuxbLzT0BAFC4L9vdtt2LEt0mD9k7fbOmYzurB6JE3ppGeQoGEe+cDk3Y7rV
+LoQUJkVAPogQjFRsPX6G9WKu856yFp4DpDs5bQogFmlnA6WsOjgxQihaE7jtnGr
sLynFA3EyK4IEie0jtc92kcxdzu/wTqzzFIWeC3YT5iJ29496BIH3rQVaot7Aa+R
dDzK1FR2PLkcut8PGENqInWvvpYoRKEdcfU7D7E5UfA8Bw7tqc52WUzU0N+l9DQj
NCEKgX/PeMwCka7SVM9OTWa9TZJqJhES1xScg2B3QgCbokHe4qNGD9xgGpMcD70X
einUseNkBQAMNHPqE8xTyNPigr7yJVrp18rmupmb9ql287BQgDg5vWVKz4+z2xs/
BhW9py0kxororGlccMzThLk/T9O2mDTF68CRB/KtBXQKFAnHblUMp1Hoo8IwWb3H
aZ0HNsLRQCvvPXgFXZdAXEFoMoG5ZRSo7AzsNtuS+o+6+Kn92g1YXfxodEOtZnU2
kqNgGN/Mn3GAy2TIEC6h7N5Xdakz/9rk4RjWkaqEODj8uxkoPmDq0gzz0LDZQKxe
XlnjCl4U5Wmc9yjDmWRHPKIdNDXmlHq6KMgZnTOvRehs9wJVLke0IrwnFNMTFYEI
W/GX1fUPyIPgFKdDWTJnkp6hgcMtoynFODdW8jiX95LLPp4tpIFwjW0Jy2QWRF2V
OmyDfcm7IJEX0FndBFh7UHEc9JBJRHqJRHp1Sxgvsn+lY2BLSPBSIzotlPUkkdO0
E2pqhK4CqU8co3KsigiUTtPW9Ew4q+BlYBE3FggKwKNoDTMcCM4QQcT+fdtt3uy4
poIbUt9zTGcB/c4QNbpsx//KP56Ri20QTV6aH5xoq8g85Pk5XLDR6pMCbuoljnOm
q5PXZi1mlda2MbsYiDUbqXRfBb4MlZwA/Iaa5CjGlJ0v5x+5sN7x/w45PCjzok83
ZMzZhvDaMlwWguxMEZqF6kljhKX9+Tu5TvV3L5zYCwcTEN9fVLIsbNN2IH5ak6tN
1pQr2o2HeCM4NyXsUuwdoRvMNqUhDCP3uK4u9Mo9/1wUyPMO+1S+DC3+HJgXZGYr
A4Hz8KA1iRZcHtCmYGo/iY46CyVDBecyX7Y5IA0qIOna9FH/VfcI5l+Svt+RIXnD
orB7llRHipIR8NbxaQ0AdEiWg0fWwZy5Q5EzGOdj4lcjGZ1XHRuPhHFgB1PD4+C1
aPiwBgz/46b8gbHqrAnA9P8cK1lnwz8fVX/MqBjtudmXpe+DfHN94c+Z+5LGiyKc
PWzbGPMtX7225rcG9wmEUjw03bXDSit6ZtdV2h0xGw2PKwGFYWenYxzIABiNxwrK
YZBL6WColdX9MTN0g5W++yD7qgqo6RKDZ/esDeoacSxyMq6rvN9qHDbdxxczsFK1
t/O1K56RYd/nuSYAND5er3B7ciNQtiIU9+gVzFzuIGHidVRbcXi6Rj0OSDj6DXOl
qFlk9WP4IIE9U9XEt67g/JaCnQbqUPuw40yoG86la7LYzlSlg6EBYlPVME7ToxZn
zZbF4b42BNJzda03YLVC4NUcKzaanTEg6Dce9j+e2u1ONTbF5UI+pjb64ARjlllT
YJ692gV/xb65vPw53eEWXTamYfMqw/JSkT2Df/PURd5JM3q1+JoA+Z4UDG1cnWt7
8s2XWkojsir0GYlzxa+ynOsMkfB8+4YoL3XekXwsFrVRR01yySyWyUsApY7GfuXu
lQ8+xQh1RNsr0OK9ZkFxtTIgEV9LQ7rviIKYrDX87AT4jA/Nbdfd5+I8QAYEucAe
5JgZoSnLyRs8JxbYw+5o5wGqNqXn2wjO/G1fmQHFabwuhf6Y1ZOQ+4fNtKqI3w6p
Bn6E16h0Wxg9UGzqASPo9v0iaT9E2I0fzZohNokxN+dWI4wMEmstj9S2nDI5ur2Z
YEmzBvVbwWSjfJzk8J8wdF97+ji934QybcMu9WcdumNgyLRSmdYrLxWn6SS5RKh9
PpGT/YdQ9Besyt/06PkUC+5r9n/sjdaOMwoEuSy/WK/ivvZ7ngy9yWb9ivEzik1y
9mspcs+Q8LIs9oyoASRbN0Rsjc2naBf0WRti6Dk0qenRajtQl/vFiaxrWCBU62bz
FwM9YHlB2Is8UNnlh/Ty+JKW4QA2sjMQhtJEdKmbhEf1cD7IPYJ//ylFB8+B8uOA
8Fi6Y+ngeViu6egGptAVbEKTH6r6gx/+0pCPTQOozetn/Mf4zUQHv93psFWCrP6v
oDt94eZAK95mwOIpDs+UeSj5zW9gznsLbyCOe++ky5DhhktWpGbyobRtWvPkgwgX
qRSxhX+1ikBW9Q7HfqzoNAgnTNCWLJwTCXXqf5mMTgjjKcbPpoFr7/kmfseSAy5A
Ngq/BRksBvB4bpG6jV+kUMPh73b8TwvhrldEJykGuLmVBrNEmA8QZIhBRPj4vEcZ
i25gOoVoKEps49jmjMFOwCgz7Nj1PmMteZi3V2Jtr8FlKTb5DZGsp9F1+D4cSaCz
URYz+mcpN1SGM43nxkLKwRKWDlgOFEYJyRE3GftEPVvPOt9tkTIWLVUXCpJsqZT9
B8u4iJg7aCWiIuHKOVDOfXEewg6JG1KiD8EJ7Xphv0FRlpz1LDkx2eUbSpvHIc3d
4anC6DEl2LbwQoA+0gca7UbKYvbLxCw/1Uuhrel7sEQLRl0BWxfotO08oGvAalla
vOGtX8LAPI/PN6pIiw5NIzk2ZyK1HIlLhFzWfe3NiughvVkKj/lYSM+IQNyUoFZu
/KNQOUITcHGy0fVFV4mUtck/e5/t6jSJU3f7YpKbmreWXtUmX3ss+Nf2ouP1C7gQ
3rQvLhTbQ0PjaR4+W+KFHtx6khDsR38CjbjQ1ZPj78RiMuUGOKCwTQjB/chJjSN+
pM7EassVjwdEo/FztnrhoAYMsvs4fh0gfVCpY+PCJCNLQEx4i2nJan5f7PGJkgLF
in29B75AEfKn2D9JTQcxbto1SSgy9Oe2WfGpNBEqhLeqj/HBXOMhvNDR5En29Djc
+gkNE0vFOQgCh+r2pQYLn+BY+EHJ4hr1c4uWnMUhOH+SB1rwDZzEj4ioYBSb8dm9
PL9TvGKURBI3ybAq3tM+GqbDRnqbbDXoiu3DcDce2OeTh+RY+oAoX3H2zH7VFQcy
DtG55GnqJ2WCKcwZZNgUYfTFUENFA3D5Jec3f4yIrYqDmutulv3gf1Dadqd5QEJN
rLVTx06Lnu/OBir7Sc91XxOGj8pKinN7yjvgWV08tfpTITLoeZH3LCpJwCuAsSzk
7wZ4VdlnreF3kQx3OqWOOHtbKZFytaMCajGcdDVxVDnPHY3DiqaxY3uEKmOa+ajd
S+iEwwtWT3Re5M15RBb2LljZRj3freM8sAQkFyh03xLoxHf1Q0QqrtjSuuixWUa5
lob6oCdvDbx2cJcO95tekouE/YX2EfRk5Hv48Qn4LUl6G+op/mZcFQVhhV/qNNRa
1KUMOrft5y+MTgYAUpS7u2fyZg/6ziMZzytYzQEpMSVswR1RJRMAAmbBQyYVx0tP
+zxW35zmr0o0Ikf+41dflaXwDluPkPEKyMca3ronTlbl+Zbmy+lwrimi2S/BbBTG
9NG2+vQPhcU129uUixyy8orz6mIttpLTPRR35JceQqCdsfgqOatRZosLuGyWpotd
r9/jjBq46wG3qrBakhjAknVYKMPll0hOXrsGM+Aa2BiW611yvtzdkXt2Su7s6vCe
5Xr6NYh9dmNsxAynZtC8yxPKT/vo630CbVjCEUh5pRv0iEef1Fn4Nxwr9OVjlwtH
jwBJju/bgJ5q/91sjTzB4/JBNLsWGmnlmJeTKd1ez7QunMtUmVPhJSXNVN7kGt2W
yXuuneMXsSIG+NmbYgFFxp5uVb/B2ObuxarJ8W3DmQdJa4WtA9NK2j+PjDZsMWSn
7GHpUULDQPywGS65IA48AmXNLIYh3CACSMjf7e2xwvTmQadiOfPvzT9C80x6x3UV
6GbYMWmfmIDtiY8DOAwrynIeIFoDPd+jqyqMhI8JD0yV5REYylW8EYcfTuHRcKG0
uZ2hxE/bgk3Aq8CVXyf9xXhBUONYy04YI87KSjf0SXIA+C5nPP13jw1FWvFYbJE4
oTRbj+qFhA3U3maBQtWZlHlErZVPh5AyGqNO9VyQH75zKH6fr9RelkDKvyV9+BPn
SxUMhMuX0RSP9oslv2JEgvHroVKGU01L9EJO+WKd8FVAa95aB90riw2n7LnWmB3Z
+ADY22Blc7yWgPKmmoLub7w3OrNvzKGLLvqJTotoHNo0qaLjVdyNiyhrkI9daovB
3EZDIUF2tZNlVtfYChERDsScz0f0coUWFrADqY/kkC13lxpEuPa4UlBz4OlEP11H
B48ouuZv/bpt1mI0L7UFRMhpqDkzy6j0WYbMneUN6PeX06leOWahgDbHj5psh6qz
bXUHixUf/hsiNtQzkCiY8j/Z46Sxf//tx7wX0K/0pGEaQkRyPIQgyjfWaarh/pDg
TbpkjrIcqvM0xjSaTCwDP1utt/T4CFwf450JQvIvyBQrNMVXUOux7H4f8alHjN7D
j7k022pPXAGzJlwTkSbBGS1DnNLcRefdFeEm4hCH8XnGzovQowmabpcLX+T9uMIL
992zpLHWrZAvbI4Q8zeBTeHorbXFqFzBxxgPjfRi+2BW8Eu6ayjulRAJ7FZe2oHz
ErQGsq+ODQkFeI5awsT1XSEq4HH/Q/zM2XDQQxJyLQZ4cPmdVvyvEBsnDI38N/J3
Pus+u0iVoHOA0hSesvL+rAUOf5fNPpHh2TNcJ8KqLqyuJ/QVqfbaIwKSVTTaH9tk
zWOZ3SWtFLWOE0BWwWPZyjglRY93gTCS83q1aTUVdP5HtruClbB5Dp7Lt3XTj/h3
vLXd9ph06ySNGHzHpeaXDnCuQRPHM+ba1UYNkU0R49F2b+nkqVvv0mT0YtLJ9S//
McBXEVPFpA4A/oInAJmL6Y3QxJtK8uhlYZD6ZTWxL4x31GUoehj0lCHJoTdiLlly
EFzpCbpuMqSakwV+KrjxF9fte4kDqn4io0bYAfkHiwDZ2BXZnQ1yMnObdLV3w7rB
jFYZc5hl2FfcHiMy+MFw8wlkXkb/4xRyVJ3rQK9lHYSmteEbw90NqpHePOs3utsv
MsHnD1CjPJZzZ9FAzXSHaA3CHxl2J5TST8oM0vnzv7r9E0zAtUfgM2nOXTgg0CPx
7ijnaIXdxMEN68zRL5dBFmhi9/3zRXFySVtrTAx0pqzU5uaxn0ETagZUz41TabAB
0vO2cGqv5wdLxWxK1DBzC/hxElxmHrLZVy+i33aX0i96tJtn8puOgQmaRY9rRA/4
fhWy91KZmRWj1BDYhm043w/SUcDGGqLZDo9aDutMWSU32ktRllCehkfew8nPmTCO
a/WxFVPH7XxVbWyf5NMTmPf5ahUhfrgaU8ilRRf2ByFfywkUA77ckqk5yUCZH93Z
2ksbu/ZfiQr4rSLyjo0/k753HkDW8q0gUkJabGhY6lkmorquK/RS2yA/koEXhOvz
GxY5CmfdwmMTIXfOFzT2zgoKH0NRcWQ2JD0fdZkYNTedoRdWbPJA380Rn8QxMHcf
3DK7lHtOGQBP6qiEy8N0BHBubveJGmArraPbbqHHdz1k5XHZsJL63tpHvM8qGMGu
pgQthIOXfJbMi1XfZY2gCmC1RzXzH3xpW4d8EdCxSpYzxw43SYQxgYjIQlG01iT1
C1I7DTa7ZvoHfM9QnJbnAeQb3vhTC41s8fpXdcY6wodAVLNG0luxN+5fPDv6RkDu
5OqgCxA7FAktzkD5AGENPlFpXN/sNCgxjDh8H3vcbc1jyUndzJYbGhPriqPo5aKb
h3FE2niO5U6Snf78NIyTYYFRs7PTg8ospiteahmhs22vd4JGt2pbrs2rR+XIhhTl
y3zGVrfiLMea/Jfjtbdjn5OuVLvl5dqt0gkBEpw41Tt8zNeQkZxN90W3GyKvq1ff
KBw1Ylhl+d8UgOW4ClfAAfV1+qluOmONlcPXciHYM4hqdiReh3fBMJVN0T+PDCQs
TfhlitMelJPuQgXDPDzKjbyBTF+8kaCMMCMZilwtm44HtQgvxT2ZOflUXK4Sj2xv
1LPFPF82n0qejpi8WQDteWzZa+PtmhiOA63z5rTKUpU99hLatSBI9rtgl3JBuoWE
akRH2HPmUUNE97pT5ZH9gmvtp/kEl3IEow8LCLgjb6fRe+5vNcH23BfKrNAFXxf3
hRQfEAMzhediRAo74DXtWA7dYeh4I1pJ0ecVBo0ECFXRTDL00XMdLonEeoBOfdjU
rLaMsn7HAIXY4p+3NIdpvi6i4Au0Q8Is0xnPHN3EzAe8drMQwvSieEtODKyyOQwB
nstX19Fi+kSyCxuPrP7hJHABRs65fhtfghngfEARRVEZq/ly80VFae58g4arfXEA
PMnSQDWCtystL9BBJi/0S1JRsNrMf+011AhPsEDv7XWgREdcgQmo4piJeVpQLOPx
HC5NvPu5Iaugtm/LAaO8+94c9a0XmGGCOc41/m52EM8ei8/oXcsRgVAMZZIns4+l
4uxexGeEedMGkkBXBo0Bbrg/Sez55Nnhg6QhtKERfEPwBtAV7oex4I80K/rBhmYM
hQz+jChzLrs2zwMa2oKJBhzwCV2DgRN2X39BKXTlP5PC1kQ1Ve/P7ypSIz9BXSfW
WietIBGVkPCcF/DnH9Y+SSd8x9y0JisntB6OyCFzcNxlkfSbsXk3xHc3vkS3mBhf
rYySwfsMRuTWrNgT5on9aSqAo4lF4O+x4VeBZ30wyDR0AFRwprA9UJ/IR7YqBsSA
uRVNV8Mwe6q4nxDy3QreUGkThGuUOFmuWwts9aB7QNr0MTULcAsPuO2oraOu2ci9
CRc3rpwJCRoAa1VzPw6XMULQhTFtJA7dDUA8jNo8/4LADz15x/jIrLcmIpWvoCT4
WKJHz4rCeQy4UpYayENuyS0z7UadB7QQ1J5p95K/vzIznZectMVLCj2mxmEB0U5W
UNlXQOa7O3K7sRAl+1P/YJko0WMZqhlxEbrorwz/W29bBfP60N5vEb4V7znUfL8I
yIiG4OqrC/QTf77YH6zFOrtPVRKaJ16dyb3IhX75gwemvbHqm/inh97AL8HZp6OC
56HrP8CbqMXOUc+A+3gq858/jzVoTXUDD/FrePe+iOkUSlgx01NWbVrsswRZypXt
Ynf6V9mwKowzG76PXhPD6Hq0qmaOwDp/Tr4prvW3L6FvPAGAQfzzJ4gweu9NirEV
L7NOnD2ts3GJ4Y5PXUwhdOcBGt0xX3Jqs5dmXBYti79TOMi463GI05YTbxZs1XiG
kEVd7gv1PtIDbkEVvituAZ+/iC7dnAntfHcP5+S88YsDKviINCP4tmkHD7z5/b61
XfpLVXebl/jfdkynK/Qo2R4aFxLbQJ7f52ANOdlj16ME0N5yrAwD2ZqZ0QmB8VgY
JGwPaM+bqsyBUxpLaqd7sgG0uLSsQAxCWoXdHrGYUioiFMPw2O8C2QQjIRDRo1BE
42KZqYLvKFad4wCUJ3y5+S9CaqsZVIzeWaGwkQ3xTEzC5x68F6QrJF2UonA9EZJ5
JsJ6orKlf6Qy6s/Ine7PrX7UxCckTVEDuRztoQoxzTnTIPxvGz8uIK1mcbDdGlDN
NXuH6hkUjvj+lrdWd9L2+5VNoHehYZbkd7PmaxGeuNF732Orflp+oIfZq1yw4IFZ
IJYetMGBOeHkzR9DrP2OmtwYJiMTsYxODdrHi/8CGQYllwPUdW1iPXWGYnzvdqmm
fzYFxDwooUxbNI/4c8J7/FAJegFJ65NeYampG9PmHdjDUIXCYZ81eiBn4FGUsUAa
xwYCnuceuKUnosSfx5Mez2i+ZxVuYHEoeMIH08dJD4H7h698hKO5VBbzM91Rbc96
NlL4F47M0tWU7GHEEktCGBGgzF7pu/EIoMK7Lb0ALfWQZwguvmyf2y1Uw5HZQP5w
+KW36QaKcBGiewex6JCMXnr6xCMXGmeqaFkGAV4iEo9khCNoxx7HFPUceCNfX8lB
9/YeRVRZihZxn9XBn7oKTbw8d87NKk3poj3yNCoAOgFWJgn9L4V96NanbJ4GlVC/
jfspvew1nXROLcW5vLWJt8O7vTzlrdhUQZYzG+wNqKD4jEM93Ba3jAkXl8wHV9ch
jmLsd3Farcp7xxXrAljS4bMOGnL5yuMl6Mvdb/4VG061P9wWSQ1vuVqiJYGFo5SE
PAyewYxBrZiwlLuaFbOkoMEYggG1S9x4AxiAPAmNRABPaViPo05UHFpqSSuanX+o
BRPcbh3Je2Tzc8Xt+kBduNcHbrmWegbN7yRxYqlA3W0hjpIc/a7K2KoxP5snSg2+
cAxxik/kgDa/sY6IZtiJqM5rjRZ6Ezt2GkVao1Lnlc2rRvAzlUiMJi7lwv48agGg
+XpWF3fvigdFxp+OX2Z66hWVCXErciaC1bTK92DnV4sZ/hDcFt2cjrgUwM7DCgvE
mWyMdFuHQx2EG36U/wx3ii6heFP3x9aIX0FmNfmcdrdQr0WtWsC4tyNDZOYIm5x3
SuzbCldw2P2NYq5pMiEj4fRjei5kyxbcudLEQbtewgI6d/fIdz7igUVvWfPXaCjO
YKtczZYWtDkXgA8UJrqhe/w6VEy/cdz5MUVZkZLTlNEWwli0DS7+YnyvvdYqQY4B
Gk30FcYvRACJRdszciJjBmLJK2IUpA5q0KRitLVMxvd4zkIEXunt88c3X29v1p0c
RYNa+4DocJr/IFWIjC/DYWVqRasSGh5xn6sRMHsgocH0BcgYqIAl1hScV3nNzBHM
VAoL67Xd2f65vW1Ak5IyVPKk/RXhhmlm8KYWbUygCIK6cd0ZwZKMnT+Be2fqI6bn
exlNPV5oL1M2XHjCVVFmRVnISeRm7p+yynR2avAwWOh1D2aItauFHTr67CxigUje
i2Vwh6He3cMXgVNVEGm814G5nulE5W2GHUYcApbtCcMoXyOOj2Hr4P4Ngc1M/6ko
hq9ggYQ0d2U9QM5MklZNxZ957W3EZhEs34Phs3GxrYi0GBb1hvBHS+ys5GdMy8Dv
vH1eECwktJEtLL+GEuVgvrtCNbqUQj9o5m3OTa7wHAPkRx5PtpQ7avBTC4YwQcQd
pQJTwH0wCUFdrBMfKYEpNWVyDpOeWL7Ss9RUvuS1Ck6YaRGsZtAGQy5pLVnhVP/z
b5ZrYQiIIieGWTZoqJzR6KZ0fc5IOH3+7RQSS0SvwQyGdTX6YwQ+3C8pL/FgSGAG
lcnyiGSlQ0OPDjWiocY5W91XP8clM5kkiiHCALBzgFgJlsinsQTiG0evr61OirSn
/X1TlER1A6H2woPG0PEXr2Kex0dXRgtIHHZdBAwLnP7slS17fAylhcJtLpqdzdrf
c068KHNwtWQWS6pLVP4Ho++1BsdDSCuTXRWuXzu2Vim7Zjt4nWh9TUwFQ9i6yU5V
xSwVLQjft1QZJpc/PHNk1gMvNiZsTgLhBBAVRTWS5SadeBlhfIxSnf3Ey6JLzcCY
ZZzk7wI6/DOwmFUFTTDeHlPpeZcjEhRjEY2Ipl+35jakliU+dVmRnDeV7wInW+D2
zNwgSOXyBxYJzi57MPUincbAKP98SORdC/kCHK+sFq2K7HDpz6tcSY6MUwFO/SpS
zm67uBANpaNtislDaNWLekCA3BCBHO+3wooUFU87+O/CVmXtBO2p1UORStZGKJGo
C5aHATV1nvnWDYZ8s3vNNBtRH/XCHRk6ZWafVNIvTyWtRwHt/AnyFJBptJFOWSuD
l0vd0VYYmKg0tNja8lFeF5fw/g7nUSribjdPRwZg/enmxRjrc4Pno8nIg/zbdsnW
WSGHrsD49qvB4/zAFN42PIwfLE7K2Bl944yOenLykTHnUB0r1Mgidzxa3f5BlhQa
pWB5keFlw5eA0DdcjLZ8pY3TU2uc6YN2pFsPWMGgLFGkQC3+mlp2iS7CiNClUiw6
/l4x7XQboHJCScjXg8tyWi0S1TM7xDFIiu/bjZeIpoO94JZoCotOO0WQOUvw2xXq
ZtE18QSGsBnsysh2tyZlN6nUofrWOYB+ZlXa6enFzkyjztJ0icSHZDNwY60J/bmZ
tqeUbstipsY5Mo3HC2setrvz5ZagvlPzLebi5/tHin4/2vgMcU+/UOJAayUFJU1T
hcsoyvtV1ZIl41PlD76XTtWoXLPv6P+6zB0DUpK3nzwYICxcO25mXQzBVyjy5OE9
d4drVIoCAmY/OqALVAD+wVlwEazbVa88YIHtKAEiANIruVLF6XEeiUMzpTvE0Jen
aKO+OhIkIsHBTHqkMb6VL3rPk7s2o66kO2H9WarZNK0bxgiMMQoFmuu7PZMcuQY/
8eWor+DmZOs8W9cyS2VvSfyxTea4NNSyYb74OtsyLDZk7UYUOPUGtiZgOEJCuvff
tw3w1EjTJeLJUrBiwPOMlwipH4ZphFWTBfMuH5Ldb6HmUbJBaGWP2fI5kNw7Vp45
Bff2MTtpGeCe+MSLZcuN5LuzJtQ9MX5x3tM0lH9zbmWB5xkT0BJpDlFizrlCjPUn
OACtjvTmNbuL8yfgzf+pxP3OXKeWkVcxVRtO8AEsj+PH1JdUFiC1VECsVOQGaD5a
gJkCLWiWsi8z1tISXyYGgouBalqbKABx5Dh+IXM0fkudhfBnx9/IXO6wYKHSH2v1
nEaBUYLvGRJxRC/CqB4S/ypJRm1x7JwRFniIyn5XJFU970D3a2ZE9KzJNpYu9rZv
+O22amtw4QFe4dsLLyrEhQKiZLpGUDy2bY3SE6fnwKV8xSdUx7g+aH64ZsdGJ2CO
iQrXD8YW7vv0szcGZT92F1NGpmHPyeziNHa+ccmWshFb7Hf4yhNafFEJZCGnoE/k
7aNVg8bBA9LDOxI/YfrHZW9r4zHDRfbcGcJjoIrfPMh5aJxxDjHha6fyMdGnQYJR
bCZRQi3bLc22qnBwCkFmyRUcFiwbreXRSJfbcualUO4caC6dP2IbtNwGENxgSRv2
iofGCI3QLiops1AkKraukJgBS2HmIyeJw5Ekm2f3oEe0On+tBnGTmIxXPGeu/7P+
XDbFJtE1lJST0pE4VazJ2zG32zHIOzo8u8pDFEklSeC0CG14xxRq+MxWJQqfvzN3
nE8NHfQ9idzFdyanh758EQf8LFGrNj1Ygq4s68XFNMLM0JfHkpuOq44e82Ojsjs6
byaT4sekVD4WPsZE0XkXqB+IIo5brGDS8jNnT211pJpoucK2p87xwuW3EAEkEku4
bLdZAj/CTj0RdPjG/gvakx3crj2HV4Hg+72z2zKqiRYwW9qGlx2ST33EO+TlcDvM
+kuDxreew66+pVfJHv4cqZbdtnZhHn61Z04cAdW7CUOxYRgO/AGcRXE5mHs+PSCv
XB7W13AKtlPrIWmAelTtpPi5/RIeqf/x1AOuvsGN5mbX2PC8Thud6bPBMHWfNtlL
aN/4Mn5ruzdGeRG37tDCzjSx12huV/SKtCKy/xxHdFKvBotX0co0/QKR638EDD48
2KyUw58OQqZJVg5twALpBaXeckJ65cEv0Am52DLEUYpNerjw9KbY6O0tvWaMc4c8
3FiG7CrcNSYZh8PQkvH1iNSkGc5ySj4AdvKWfAtFBpz7lNd2uT+gsQoOJKF8GhNH
49a0I/MW/Du4YPiqWZ2baeIczk7AkReAVtGfnPhOB/Y3ev7ADNc4IEXoB01jd8ns
n8IJhsxV6zhe0o4PRLdkOYeGaC/UEY6J+4RrqpJ6eqKAHOEVU1ni5TLsZ2OOyZae
c6QOBrd+RFp3n5K8MXGj+e1UvtmWYGnFyCX1OmOa71ym1qpyNYhB9V2/DlDYyY3B
tAwFjoQvi7b10Jrja+/AiK9ZsNtSVHP2r4WfsU9FOMP4aVyhKdARPGF7UvWLKpNQ
tjqJWdZqrDqlXjvWpddfIiIz8YWapDivqeFFGjxINJOqr/xcvwS1k8xIody3uU3j
S0MBoLyl1F6Zt0TvPcQMb7Zor+IhGzBGMkxLMl36Ew/E7QSNZ+OMaIiGsc5zxhMf
ey6TfMdSEOHX+XJZ34jd9sWQX+uI1JFAs5GiVEHl2Xk3erc2cbzwXAtCjSVn4e9Q
siodT1u00jZuis8tKhMBMfdfxqu+P9EN7kdCyi0TxyLnTwPwPoK7NzQ47PNefWyb
HxPKZ1UO9rBthXmiOkP+cPulwEdRi9JzgvqW3DqKmDFipL3wEIePFSMdV0L2uc0K
/BREcZ5W+aZt6UcfNlsBHAR78D97fES7xS1tcPwGUpqdmlE4r3hgsJwKnhAXh1tR
yCheRGQtV9ZWQIZEtf4gsmpwVwjZ5u2JdUGigvsKL5jruJrR8C52NDcUbbOHiRPo
haFF0yPHxy7IkKPqz+FnXqM755u7X1R4UgfXLOdc4KHgFllWdQWbjHcQxw8GopTI
vocTnaqc899PwEBTD8UdhoWETVDYcMugaLcceG+Z06039YNKdM12j9fQuinhS0/N
Mm1nADt3jB5GryniPU+VCMsX+wNBX4MdKnfsWcphlnMTf9Q3gGZel21aFclOpJuG
2Wj0ythBRjH7XMMZZwzjoH6pXypzfZfE8f1VitLziL4IyM9oif2mc2LXW8fNvyoj
/bqaZOKZ6E9S9wjXJoTvOqqu1oJNGVLJrsDgCwCCDlEEpTxVrbUiHF2NxcVxofAD
yJ/ldFVwqiCi+nvehbbEXCT/ZuLCBqXj+vLzStE0X+IfGK/wu+0+gIC8BkWzJgAR
khsHnXxwY0x9L51ENsUNsIWr/5JFYObYTuYAucomtj9s8cR/6+r00s7y1aBm/d0r
2jwJ85pxNJUL2I0BXM4TXMRPzBgL9LKDd1f2E+pLCmcfUGr+J8EYNgFIYGqlwmON
Yh0ULWmb6kFWjJWUX+BOx3aPNYbcNNgNqQTEYiJLsMKW/hpU0SRX1A9XDdUR1vor
3QZmJXxtpJzuBnXELE1G/xOzCtQ09x2odtjhdcgldbhfBhCMfOlGab0i7WupU8xI
4tOAXE2ohSgBykrV3WqmckaoFjK1AKeNePR/nExxYdZlXzv4DWBA/LmJRWjb9Jnu
E5agPYmXsMetRhDRffP6G++ZlfM2I5+WnzTyV1AV/zycSFQhFwxkVPkY2tguQ5d4
G/zFvhLDc4GUmbEbyvkzotEiMZWb3aC2KW2swl+iTn7qfUCyqVkjyJcrpwmI2rI5
cK2/5XYmRi4DFpeqX04OLh66k9ilSfrYVCqYgyvGmSBepJB5GVcJcQRzexldr2U5
Leq6r2SKB+wUDF2aUuazElQdbaEaXFSMg27wyBL6ItsSJFZtMwe9XE9cqe8iSeeq
/O19IkhiDyPmjX+ed+/cYBjYkkwThmnXzGL9CBNI+qynEEbjNdQN7T4cwk9o5I3E
ZVWiY6WG5eKqgMmgDPWa28jbCp4X47cEU+oVn+Z3uawRz9FbQe1evwPemKsZTbsd
MzhQ49Q20s2WWnYHN+E4jGaEPe41XOj/jlJcqe7a4YPFjVbG2ktTzc266lEE7nCJ
9Gh2m3xuMIGUN8uohFGpYkX0murGLNxdheXGq5K1QRXoSTfKSFcctwGEOMqksq3Z
Q9r5zmpkGUNoyj/RS8AjnmIUeYsVdhz6qxZot+6nFvAajENMrxD64ck96FAgw3Eu
lsSutEFuW17AB8LXwnNp6H2VDCfTjgVTniZ5aHubw/WevQVj+T+zJC0y/89axfyR
Q/ReXp4TFowj6uX1zxg8rLgGBTnM0xLSUIYLVNbFdMWSioMqtibWfE7k0Ur5B+J8
r5cM5Tsfh00a9yWVS0WQSR7rLLJ8VgGeKapwI2nkPGKcytn+Q79TIUaE6HWjgWsG
IJDzaLVLYQ+McwZmeRfcKZeKpFJrNl0g0JHa7VoYuyh1cuUCY28yHOXJbZh8WNem
xZmqK3bTk8HhTK3Tnl0l7D50RDqQhgjEEW0SR3BeQyv0N+5ymXvvRUmsdqp8oAXU
MtaHD0LHY25/ZsnbqKkGdwSJWCXipsz/ITnik2FjZKb175dbvAxdohQd7OscLD3E
AT9A36yXZ+rwLYMK53tAZKiq9GG9/8laZfWLGRJfKsWn3LpR5nOOTeFIGnVlcGQX
ftMP19n7v37kyXTAQ6fC6qYQzydxzg+22C9IwPZHV+ZTKWUZdeKss7CRTZk4+5oZ
xJ/AHWwm67L8GDlMB8+fyHZLtrihypv9X0aC63Iu7RdObkwkdOjNrkgljRlWENxg
vIUskMKG0hhp236QqL9lkt9YIgXxHIDf1ri2t0iv3FrJ+Ue+LCp5RBaho6UCDGnS
tU3SuSzzcFwGzyiVo0QUjEyKdjAy+OsDhpVsoNFmFtMLuYGUuQCp/EFF65vjpkXN
AvcgDmFqR407aNqVWriMkbbkHpgWQlCkKAsBtdp2UQozsXvkQj44Fk6utFzyei0r
HlkW83d04S2sSSErAGDVfxA+CJukZcWYK4d8mR67qTu/cXXtT+M2VWOMX3Icd5uJ
ezqaXRJSSzpfD2ApnDrpPirMd6wPGalI3jHUFTAVixvAPvrktau1OkyPgzZcS0MM
wYbsD6zWdtLjglXErJV/wrA0TbEBaglj6UWSTjj7W0jwaauqCxjdew7SIpUdTL1C
Aa6nRvgIzR5av0XyT7mF9IqYfAyVHsLBAECx1e9bYKZ3JzOBhEQ1O1K0947GBJ7E
84RXEDPjJKyYAPEN5z/y/zuXnmJEBtLHDVdwZFIlSQDaBPLjNozipC4G1OUMpTZ0
TsCCovmknIYOoqjv5KYKipHuc/r2j1PobPDg56KCWy1G+OPP8WfqBWQWMc0Cc6Wg
UkrWo9melqFcgEo4fcPWHYCDrtR7yygc21jJpEbSNA3+gwuFVQYDllRud2BiqvRk
YzH7TmUO3w0eTtagby834DZeunGUtvxnXhcV4IqbkNcWeI+Mx8vrsmzMf8DKmbRC
otHkBJ1z3tGphk9+xd2p8P0zNOF7vTU8tyxB8yWWiIYjvj052IOjwqC/zC7PUMf3
AbwKP+ftV6ZnuIq+2ltqA4xXVSVWeReJ+FSGpyyT09CMK2pMJ8WNSNA/MZ8E7nCH
H5eT1BNgpLYT3U+Bkkx2fcvwik/yByXsqCOtJAWdbI3pg9kOGPd+F6XqwhpZzU73
HM53gNNpiD+QiwJ6ah8cBJYwvhWrizLeqPlRAF4U7RvknL0PaHX7mP0cFV982Y1/
DlHbPUkx26q2xxqDs05RvYcB61wVQVH/hmUh13fKMPZXEqphCoK39yp6y1CSzx++
QzM48cTZbz5/Dn7Ixxy1QMwq+udMaVc+dkH3e2TK7OSiyH3aNSNmrvTDtKjUdkCS
StYe7C7SQFEw4dLnk6C1gTKJKKUV2acYQ3gMequs4RAK2x/yHMqbg3XQAjJxMkI6
KqWB2iYuseK/e2gnG20v6DgNHAvBf7kNl+yF0gWoU8/eEILMSCiDjuJDB3N6/19b
ouTjTe+TyBbAgdGUbo+Dnha4w/x2t+xwkRUz8imExB9aOpMzxuObkwxsBMW99IxB
uinKHjxh9FR8DFVPJ47wpyYf3XBAdNTG3sVJyB+Hz7XBhN/ilIJby21+ekGXue5j
4YcasD7+P3XXsMiwlc4ewN92JLuzWE8RLcRP1oHd3HLF1J5gX4JkoQGC6oVVuYeo
cJ/1SboJOwFU3eeiPTx8mssbIS9/B3KY9mx4MAaZvQqfwG1hz3M1FCnypnaG6SKD
qRjDsTiHK2YLz7F6H4lX38GyvaGq9cGHUTmEiIw5ZIyIjZWm37Qe+NnNeEQq7L7e
+++ne5TL4DjxR5up8Xcg7ShJnaTNRkcVvbjHW9lEvdTB32Ym/I5610slv731MfsG
wRp8sNSnLqro0wK2tHod61kurLcfnndTDmzt7VDh/7n1AgOiP5qJ/AtnS5FJDgyD
mXo+J69/5kVnrBvKh0sYpTuo+00hQvB3i/9vq9Y5hPHz8DMsP7Ys4I9rYWg+BCUX
Aet3X3IULnbtakDoi3zaop0dVNngcQOVIExenlredIKpIiXjjAXgtW0FnpIH8ed7
D+uObcjv/kTLgHdaaKU6V+pHZZ8R73lnVqOosas4opDs38MDIYOW03oxpRH5kuA6
6iXY+G5ibECPAtVtV5PP+Mamk3NJKOVdqPv5Lo++QQU0RO61xdgOIp9+hXV7cMX2
R/5LZAQkvpqTT58ubVGUmolmg2xnFZe6ABGkj1S8dVX6Yz0iw1pwWBh6jV14uWeZ
X6ouLxArAwcWTk/SK6m/Zw7UygsfafYIb1edRr2NobjDr88izADTdRsur4vwISGC
E/ZBilbXWGHctoeUUZP8UqBKRg7qBTILSCiU7n5njChPi+P5EtJxMxni4y6xa52E
qCQrolsQAj4iOpi3//qMrZ56D6SKMfrP5YelAFdla10oYcvDoISZulzw2pNi5c1c
58AxIGq6NJco7Nn3W4OtDfg7i8McFUwX5bZXj5NS8yIObboco1phfeG978ECq23u
+nGHDSlF37UhcxCejla394KOqtt+KjT43MlJG+PxiA7695qyZ4gWLAWrlvqQJwKn
/TOJMZCu4NgX9J6SZnE5mzWggkb+2Jw0uhFC0goGInB1Uz6kI0KFq9HIWfUzbBfV
8fTpqucEThNkeiw7DX2OpgCZxV6hD950gNdBA9TPN8aH/j0HwjXoy7Z51hITWpzZ
KWCXGSGTwDmT53tZxV/IM/xe3Q8WEq0Ju4ggQdA6mIpsUOC+z7BjIi88kIbSarUz
ab1y5XH3GX+WY1iipqoYv15jnNWzBM8+CsUIYQ3ljkEUZSkWFx0oTlDsTuGqEWWj
K29WQjHID7522tKz7wSySD/49f1Fknt30SS29X7o1HCsS8Z1JNFWFsvNFw/2LlJz
SjJJRbMvR42m9rSZ3u0G56Gi5yPyZh6Dg2bqiMK4t5pEy7dovSLmruCxo49Vr6SM
CqggowKsiE94Ron/akWGa1Sj1EaW5KgykOeRHIfpxXT9fEtPTYOAwFNruZvHWBdv
iotMszOIik80xYy8CMFmv5PPRZxv3zBYsB5vQyyI5GdA+xzVHfthpSiSwKloZVjH
tML0WuvS87JM9aW6K5dFwuM+3bSgVDgzlq4GKN0PMGeFIf4LOd4saI6SX/ynWTyY
PrYUcdXfWSyNBdbmBHDlAF/WONtgBOh/Ylzabf+E+sjjXSRVlpsPxukFIAQQqzkR
JIHiklj7kUGd27Dk2GNdsv5F8bfD1kUszHRre2OklwFD8tImtTaZMCXDBXbuhZMx
HbRjzjiiGtVjfqsRCf7VvL2ixopFeyhVhX1Gro7nZIS7DqLBb4Xh9ZWkSthfbMkG
zlXwn/aMZHQdxW9pwA6GKPwYKdDT1Mn/tqab1bGmW1jSHVCVeSFwa9Kn+ZgWKIaD
JRHjapj4gj81bufBsogI+HsDEmErKyUup9+0CIkF2OMGbsXblo42dyYYXmTDP9MR
VCEZ7vqt7cc/uEvB9IAdo+/l9jAisBkVouTF+/K+DFKcazGX+psImJxJ+CYO138M
l8YaVFpJU6ob3ZlMB5xn5x8AfybVSnEprsGpD1PtVNsWJXj6UWqNrL8NlrQErBMw
te4ow1fNo6QbwDdhH4sQxgtqPoU4jGueEG74uUwGHlabILFHvZt9ZDqutg+4PEGp
9Pcv9M+c0QxL69yhg8DKreeW+JCx5pqu1o+YAhHfKUhkJJiU5AbQpnqCvE0YFQXD
+K6BmrwsQ/aliFTlOp6ZC4V+N03eRDn+1M/hww83OnizOnEoQlAEeKKUch5JBPn9
RPzYl7Xf87qtVitL3hRYW9IJDook9XMx8XfOex3bHf0kiEQq5YU90EBfItQRlusS
ExeouhggtsXCtxgfAD9ZSgrH5AojHN7W+E8iuNdAGLEnnhHd9TdAXzUSnIW8HiAQ
F8+fdDG/sPtCDvBGJDsxFitqBOVWG7F5v1CHv29361MWTK5hT/EDMyeIWxKOH0nn
1hzS738JhOf1dcCN42B0OkNmrwpGPtbVJ/QBRk31VCiPv7mzGfFCpc+ct9p/nRwZ
+Bxd399u9YA22qimhCSR5sjaSc+juX+02kyOGZXr8Qtv4rXaqSiq48pKcvyboElF
rt5ERaIF85bdHTYzIDopGZAEu4uQh5TkM9yPGvSAY6Vf58j2tVonxSUDg/PMQO3Y
Pm3ehQB2Zyc6zPqA9LAnoV2rlvvqKa52j4/cHAKjk7n20+3JO80aAZXmKcV+KKhe
Gnxv+O/jZR4ih//Ue79dqdW0xGXhCQKcO6LkPuhRzr+HYUW6rqIrOUhIlJOfZ8nh
c3VivrRK1YusV99jvF/4w8H6BwCKnnTytqFU62D8CBwiWTw0uAdW4JuG9TrnY0Jn
baWs8cC4CztMaxmj3uMVDxGFFNckIQWp9hXT3GrKLQY6nhVVnaV37KHWTDR4l8za
0nqXSLis9RMp61iC8xSqfdy+uTI7KJWEkwaDwRSFpFgK3NhkVHdsVYb+mU4oBeWQ
dKv+cmQ3qXRt5MYqLA/0kemWZP+Dp5lWNl+t1JdSWHD9n8nbQEhUOD7siCdzgg7l
oCx20hKnZsQO+LokhC/9aPeJQ5Ihp7HYNzXo0eYA41Jh3+HOD1GwG7yVVvcndzze
XbwYb9dxWWyVLLWVfd5Sx4W0i6WY2TAa0svSTSmsurBcKinKqAJ7vejSQr/XkXj1
6EPwibdKIz1bdrhhN+3yD2XxbvK+JbWLyq/aa77x6/VRLpbjRxkH+BUIm5RctPgR
P3YP4BNYPDcncolsLxuCQKqXeHskFUTChiI53Wq1Om7zWA2EA7m7aEv0z2/maH5C
GQ6lI/KL8n5YuWH6SuqLHRFuK5Yv+MW1uNAdh+HUswObtoTui7MWTSOd/jLc3oz6
JJUmnZs40nMiw6afQJ5LLf/K670XKAYG3pfAfOMF/WitMDN2ZCxUiw8SAXTG6IT2
KrR2xD8Ah/Ss/qeTjbW0VAYy/UKiXXgpYqN9mUdzdI4WeQlp60fWQ2Y4R9cBKofx
f6olRjcdc7MzOYBciQvLPP/KZvacUX7fzb83JycAZHazXDsOBCsANYaAahY3x7PN
vNcv8ZwzT7+EnSpxwDV1V2PSQ4zts5m80rdBf3Nczw41Z6ycYxZDxLS+fmKkmueJ
khPtumse0R2vSS3MXtjuajExJMRn89he32fQrQBdQBcvjR7k/ZvT4In8wgeCrir2
iCjQpxxRo+GX+yRtsaT4qVOlefi706OfzMxoIrcoP0sBAm5TN+O34SxIV46TA5qK
Y2YotqtTgiZPZzIZUBGIXVHnVXa+GT754UNS5wQMgicg6H2RCOUH1LvBb9VrmY5+
oBdFffPiX1ar8k3BC4sHa8Apk8GPGjEub1j2GhN5HqGO6Tv82T/s2kyFp/Ay/keA
Izt9pRmCzt5dpPe5W7+71lAZgUWNOGbxxdeEtMyL70VrsdH3L/SEwasH0xDF+1yf
u2UgaJgl07rf8fdXDkq9/dIaBwyS3a9ct/jmCJ9wAhElVjSEGc1n8BK530Yr++Qz
+YbFjZWPyt24z/wJ1c2DRJTq9hTU9w3VfOdvJ/L0HvmTIBg82vCL+kqhGkPVtcuw
oUx/AmwiP9TrVQdtFnqy+7660lefLhmWjHZrjGa8Q5SfWPgVFUYjXAydQ06WCRVu
tV3pkDiVVBONmBc4T7CUUKLv91I/Gye1QZ8IbrVsPGtdF59snh+pNFN5QRuoot5t
YcbqqGqQ/p5hfsY7svs+TDjhYRjuD6HiVT+n8ZfmddmFH5dWXqghF4jnSqKpX7uk
di/QtA47xd59TY8TDEuAG/aYejgyvNDJEzgo2h01sOdX0EUBdLsUGbHanbaRbnZc
+JPP7o3RfmGe0NbzMCDROVF/x9w8gPSUhJk5rPbeoBJmEmy9lohEIKPgWCHAzJoD
4bDoMG6VF8q7tKjRJAhB9mHqTZmAyUmAPUqE7Y6tx0gVVE3qRBh2+f3krfce4JhH
D9dRTstqsOOODbNzbcppXf7HcjgUBcZltiJbpDbGqot2Jef1sJuq4N3gRIO5H47e
aXJSKJiMj/BC5hEfK0RSH24toLnurB0qg8Q3lUhnEHYMCqj9oe4paO3BBvb3927T
EEfPhUdlFE13QGsfjhaSKeIPvq0x1Lx5rM/IrV3o1pPi7JAp3eLSTAImJAzkHnKR
n8RBxDfTveWZyckf5/Z8y3vuTVSDSFLcYV+LcmpNHObjrTb5hZ+nZ02ITLQKvwjP
BZlcZ8T7C9Lc1JfWWj0g1AI1AKpx/Gn+z23WdYRNLOe8K7ZnbERPnK090MzUngOn
Z8NJyy+rVHIXfAPh1ZisoSiboA3TF0wCN54bZ/K5A/3gqC6ADRbcAJ0O4maI0hhL
8SQ3wrCGUNiwgT140pvxRlsBidUxXZyt7fzr6wv6u03qQ1e8XcjsAawQZD8I7Yak
sFc7bRSJcFwMzN2ldgxIrDL59rv2AD3GhAsers/aViaitEUPQZlVmpb4IJDOxfg9
mufWqz69RNSTsIq6hYj786/JK+tFgGMSL6xrAhKf5P6UtZrPL/Bw33wyNPUPSx4C
j6NPcgLgFj7GC4s/fvO3pqElPLgNgL4nsz7zDoQcHjdnXpZ2WdtvuBZz64rK63d9
v7QFRjcolrhezupw0xO83KirqDQWjcAXsxJ3TMNpmXL04+U4cGd9j/6r3L9azOhE
pflyYSI8lbztCtYmUooMxlGKoVmadedjChvOKaMMfvhEQlKI7vmhtzjHLHuLGxHy
1x4Bb+937AObyUy0SB1FrPJWciGFrArsR4qnHIVqy0EMtve018JF5KZfvsP+1W8T
ozFKb+Z9HfFlO/FlLZ8qnCYBYExGGpEaMbHAoCjWQIDsp2Npicdd58nW9k6nciRB
qo0+ZCuj8wRtRrWpBVBXcjhSoj24GKGCglEOPL8QLUZbf+wxf4J8T7b2wf4HbyKp
8iGOEE53YdLwFJRQLPygpQDxRplvEhPV+q0xvnZWuhnYwCgpYM5mSUZ/Vyk/46Q/
ydlPiePhY0OH4O9KPCE61SDxvfJg8Ds0tGLI09leiGe22EL3zc0YMdOmIREBe5Oy
rOy5LNiB+LiwYk8eveWcYRFalrqFBXV8TzVtlEWoBF5zEJQYV6+dlk+nFeCgl4By
iYPS8AgPZfE5v5LBQySEVyxM/0noHuRdxhdnBoIzXfag4MrEh7z66+apYxGI4Zgt
coqz9qpetTKO00WHOt5deOOp77YVyl1zI0Pv28j+iUUePtNKSyxVOWEQwLre0qpE
yCOqOjcPay6F7nkY4eu7PBe64cjvgolP62BJ/I8Vrs/vRaUkHFl6OtOPzJINy3/L
Y86e0wlY7DQCfcXcyoGtvhgRVYyfByOj0yxKz7dlvT+t7/A2BH5ylPG+IR+FVP5u
72fzG8wJRYIt+VeIN7v878zjaGbd/9xUyy5UPjJllZXtjjS2QKg1lTY2SZoMUnam
Vr/Iu9ERjGZXxPPiWmNT5mNN6fqmR6SfbnxXrAXvnvgXZd/1YqRyGUgAm8VZY7Fc
zLvQtjp5B723w78F5QuFMmprjFGUJZedOpFByAIFXNT06JNbNschWaR5ttDldpcf
TCUzxYjDuVY2eboRsLHEwtS2pO/dtZXI5P7vC7MEAWm2MEg0rzK+eCWWTft6b6lK
NuQsGZKWxcyYtDUyuhhB3HQA0f9sPtm8RQlZWspgaJaNuTmaEwYqpNfz7kj2XyTt
53ILs7LvhLnMpSBDkeEOUj8F5MAuduUoe+UNA1OFcuhxqixIVWcZWFwRIzAWj0Zf
jIBqnfBEU0EyS9Yy+Ya94xEHmG/fOgmhoKqxkKLxdowEHiRt5Kun5aISJtXJP7BV
c1RpiSjNRvoz7ECvioG5MRRcy2HBso1YMzVPTTeEJBxfJT60hxW4W/Bitt29rXWG
Wf10mhgOk0IBSpEcsg3IdvS02C5Xx/kafIk/bykchQYJNDjLMbUtTjhFRmpsJdHi
VNQ0JuDOWnNMxM6DtNk/i3kiGjhg6VoDzZPOTOhZglZuJ6ZYaCuzrfQMbIKwkeM3
tgrxCNN3+8jzwXhIfls3dTn7BYf9nyHx/+Ltcedupl/WHkoz3kk0pUD/oIvEQrvD
Tc2oZYpGYgMQgbbZSasLCLHmUYl1W/gpm2ompRXhcRsFQiSazrdVuYQNH9wFQqQf
7ZhDaBY7/hFv0+punSIwKJ84QI3nFaR0iBUmyG5kflq1uOfhunvBBQIxjBounCcK
Elx36IIA1C5OkHzh8IgaUqc53MQ5qZGvy3qACeqYP2crCjr/F/CuH4Zfev6JnzuG
cCMuJNhfALa0Aod4HH+UHUHywdc3cuYl+SxpxGtIQr6cNPm/TnWCjrMyDjKrrZpb
GELAaRgj/OONpPQID4uwta6Q6QoVJ4C7imEjAGw8WNSsad/fv+1rxeceaiub/nr3
v+GWRoDcSmFgaoCUdS/IxJVT9YUSaxaTpw/KL09Dlwo+GnPcKflTph1d4b1kf/zc
U+QVmUxjylH+ogmRHcrChWRqP08oLb3dmY9FuJeem3EYQUqQdtW8XXV/eQPMjzxM
ynK3duWO88JH88PHXJKqILGY6rjHJm4DxZL+UNP9V3MyGy/0ZjZZgY6hRTJR0fcU
kE3/Kul+O5usZ9Y0LL5AN1cvYH7MQL3LuykDDhaY98/Xrp0Yby9VrcPDJQlx5lcV
KO2jPEol7fetGCsXzENmpprE93CJOr8FBznalHdQKKn3bFj7kNRKJ5U4IOzXBVzf
ohVdgwKUK28JV9/90ejl3AAaHjtCQiwkIJ6sJHCdWi5vJFHVgFP/fNveWNV9m4KU
uHmEeJy5FtGEBiaR0u5j2QdcR0IY8CR/nLD2ztnEPb3y+NyQrvVituts5Pqe9jlN
XA3PZ2JUKxW5AS5J92V0AGzef6qtsE34+3sUZ5JKN5aAH8uHCRc47NSWl1dsJ4CL
L6ZlglKaoXHV4JWh/Qh68XRM1OqDLoX+DEo7I7Q4fhFH8C7iHl/EY9q3XkibWVMZ
41RBLP8UhhbEH/PwoFzecLJc/8kRjORz8LBmsBpPh9s9wFXvtG0cavf9a0vRhlQb
d2b8kMSeHk1doF512hpFX9qAyzDxkf4TE/LfKVnkny7n6mvzqbsr7GhLlOQp5yi8
0otEglVkmgo+gkhHZ9HpvUijY+/0wgAeMtMSglsjwx8VujIykQDnBDGc8KFsh4Zl
CrXTZ/zoRcrx5Z3v+gGGPZr/a/qy2Xmyc551JirAUSjETc2PbCGFW8A3/QKocz5s
mLwE/IwAUY+2lXFL/BS1DilLz9y9jV2dbLWlzfkUKBxmsE1Lvjr4XhvvK/hHwUoV
vI6UBRX1Mm0zNtrk8oW7KD7HZEPARc5citCQeWGTh7j29MjdCN7TnFQyOmlIjsdm
H58n2qPUol3DqRpLmivKmM5Xoyru5RhLM/3bbGLOrd/xxaE59iCDTybI9QgAh+B7
mLH56gNEiE/a8+i+YsikpLewEXQHknGdHqCs0XZH5WMGwz74cQrA2ke9+c6GoJlC
nEilSlzLw1yGoXDbEz48GBkdjXmeSE91Uym04+RSzDMiYj39jbkG6FVaribWgzCC
YhbdmkdDoW+6VRLDxafKdKWXQHFbX2gkb3s3AkKFETdq1FD1Cj34VzozPqmxR3qy
u0zOgZ1GO4hyfRiPL8eIGLnUfuhidl7L91LcuhmzrKkU+FpvAaKSM146rRtm96/j
FiY6v1GYtBJTfz6d3jHGGApX11umXdQCOf7aK7HnDZXKGVoCjb68X4i+ex5iSQ0a
UmnOndjOdaOmCTfnUuflyF+FprHv4mrKDPgHhZo1StQWyXp1AljLUtQWCozbPD4Z
1Tjd8cCZD5UVdcvlBa4lHJHS2yG8c7haKxvqrm3rSavB5K63ik0NaC65+A3iNyu3
pcsvXN+6ie6XVHtMk7cEgeiRRIhBLB6uSc36ulAcdiegzAJ9rqJQ3wdJeHukHFLy
fTI9jcAcmWGXyDNDAh7t9TcGrF1Wx1Jz8TLwvkwMG9VpeMm4xDhi90OdwoqVuRAw
4vVe8xq5/IV+B74IxkI6vCiXMysEDSyZfd2s0EeMoqgaWIDJB4dJHhTEUoHLMvlB
zcnEXCvs22Gz/ruhEsJHpkyQv4pI0uxkoRMSHYEi7Hs9M/OLmvVVtAE1JWZ2id3m
uMowlqu5VlWbj4i68uYE1tGfcszD0PQM37B+qW0Od5U7XNyBNDN6gWlKEQOnbgF3
MwZ7j36sknRFpGyu0Hp41/iUHNJk5b6VYE7BR+i57cXHrZ++QmHOncjFWsaPbAwA
DogCW2TopMoXNBIekNf+CXquAl4I/mespSNGfK2UihhJRukNxIG0J9AEFQwxyxQu
yiylNl5fY+SCegkL6P01cxL5XTNEC6Nn63djdFgjWyLk+U6+cotsw2mZFzF1ve3p
/rMjWm8DQciErNbXvQJmPc87ZhgtGRgKfSbZtJj0MB16K+el4849L6npkuCc7XBj
bJ3QtLDjWKDTwZZaG80KKvSnHM6Qii8S7d0Ku+JT2TQvLfBTpegAL6XMoTgtoXJc
6TfzV6WwLPe/G6JCi0xDFyqe8vt20KrJagu9NTphyVrVWygurVlw6pHlQswhoE97
7PZ8BsVnIg6CbvEntN1PU6DHwYNRr8obtIyrXBQHo7hfCkKD/C5V+EUgG4r/tzQk
MaDrT5ov2A8ak7n85rBMcOUDVN10kBhig7fZgRzlYHIg//SYIotL5x3HRgyHijNk
IG0xZ4aCXaIZFxc/KgV8zZoQVroocek8M190wklY9MIexYJocKV9IQPRGpzQXukd
9LcWqE0Kt2NKOMqWwp+tMf7popXu510n0UmVTNVdSPR5nMHN0wI5fVkZQtUETfmA
VOxW8fPWCm3bgbj2afDRKx7VwGF7b7m99meloGAWddZRi8KYmPKK9gp8Y05nazZq
8mkyLFCVW/UG5nGvYJMVNXSsGY9C5zIgU2/1g5Awght1+UFWxmnRrnJFdBx57kDi
YUHRM4qclR6w8uMT80phwcNr4KZjCHc8MkckqUqBES4fdP2pfcL/AGF4JtcE2bxy
ogFsyjH2hBo9ATie7zb22WsKPBtxBShQbaUUi5+7u7XlOftjmMkq9N+hyrP2FGOR
cNNePWriDFOxs5k8kK1UgOtuJ9npsLyfirOi1gQXpj1sHYiU0AshMDcopYakyEJm
LYRWytyRuwZb+IzYMAa3Ry3PeE9qAeNZ7xoLV+zrI2YKyqDtpTzcTf0giolHc/W7
EnIfZ/0tjrGEvqM4R2CZIYi+dvzychCrj5oyxEsbPbzWeev/VNKQ88zAbcRxJ9au
wxv7QHEILaakNxn0+SB5risO8rObQzl5+Vmj4BlV05zNgT/cGPqhArGOQizSEzWz
04f6v87ZxpTo0RJFPyz//GdrZLiJYpKVn/ys/cWtvyOmu6cKJMwN90ORgnTAjE32
3mRAYH4fIyiPVHIAXmFiKpMdZmx7aKpQrqzHopoNJQkS4IDqiONpzs0hYPtAaoop
MVvz4emlDtQc0b1HwDuhCOF2NAEHn6Ib29INj4C5n/lT6n3aCI2tZXZIPJXdDgX+
sF1Tvcf+3mTTwSpeXT1VAGJuckrcgU/nG1bs/BN0DHOX6/LfNyHVMdwlvX9byjn2
4DXrgoP5K8gXct/pZeBMiJVhgKafF44VM+gshOdBLk7HQ1nMg/sJ1ZhZX+GFsTGa
UvvKhjlnLdTb1o/WsahZZM8aeSPQLAlUowQKWwUrT8Cl9kWcF/nSmtx4ZBeU2nNf
N+8sAr+tr3zB77fxuES1YLLD06IOXy8gyTFHqbWBF2NCztJ/kyARaeV0Ke5ftOhK
XQIsFUX+rnu3tNoT0OqROJRgnSzhUKytYirNZJd+grEo4bEltAqZyxZzVI6HRWPy
ROC5koFHG05oPspiV3BncEANd+9Uinkuh57ThjWRwjJsRWIt3nO3Zn4Tf4mv6a5/
nVcxLW347JaduouIDl7P7QAQvc6vRhfKemBjgusc0wP54Me9gZYauInFesbGc0wn
/VeTRgvMQDTgnyhd8s0Fo2AzjRxc/tflnN+IsNyBwPjQxFb4ZQdWHe2FHlgTIxQO
lxZ/tI7QNzEPa+h1tGJVRzHEehMmreT7EBv+fc+bNkiZa5UqTNo2MIOZljhFVigN
kEzHLv8ZIQk3fAYMyq/jWh+CeFXyNenQP2Ux3rUFcdaHw7UBZWpXInOzJj0DayE9
SL+/jp8KqG7iqiTHzV+DC/3PXm0RZSqa7YB+xW1TRd/c5584NyWYw/u7hrhSMcMN
zk3kmigX2bXk7h8eDteb//mkQhJgXvI/XNahjHreZSzfOcteIEFam/roN5rySSEW
4/xTpYim5H4FAvgWGwhnQeKG4+ChaRpQt/rRddxbI53EYanO8QbDEgoPHAWQd1ZP
2u5GpV0HxeIflTRuLGT7f+xwgg5TS4u7GmHrapEJpHODur9SFYOcVKWx12UoOCR/
NtQ4qnySX0EvOskZFzCZSg7c8Cz2EIfE44ZYwKLUhdx5V3Z6B2pMOaEv1EPNmn+s
YwsonE5X/DJfdRRTed9D86Ao3QQCbQS/isvDxa3OIDWiTNL5930U4rJPTGEekJo0
97rNeQvdyFpUrfMXQPbBN3e8kiHoeF9V8RufqB5XyRsQ0vTzvauq+3Jdcg80rzgH
mb0+vEYFe1OaUbOyEiJMc+4UVRuk0wfLYnuvVbbStLrhvHEZWjyokmOt0xweW6eL
cjmejPlr30AzllDEXJqeWqj1u2IhWKvxnurYpz9JOa+z59gdDoyJGKaMIXFTMY/b
Hcq77FRe6dR/4wf4NAWrmNdi8KNDD8oPcGRH+coTj0XgSuZOiJb17XtRrxPVVUsn
r25iBIjMu66cx73VPkYpL7k5yQVU4MJuxYVzTzH1RHjO7B2t00Z9wbzFfG7qEvW1
fYvwOFfC5GK4bfx9uCwC8BIsy9/yd3eRD72ZgwEKsvJpHZnEFv/VO3cug66r+yIR
/+2VPOmCOEqSyg9c7kzwchN6obw5phORkC4TzCFy1tCtTB2OA8KPXeBE/gCCz6Di
NZHlvAuN+DR0BeX0Q2emUrknXoG8Ph0kjHp1fcDxnE/iswbWBS09ItY+/os8zwXN
hrwTWxFXoMzplGAH8jALGT8j4LIgp+pJL6p0uvIBQDD+s3zE0tWebYF3I+C6vQ3w
nE/91UyU8MnFoDyuTzRDOeTqqL4D/s0JnLUWJRXVnlaRwJpspN7i5897y405gyNN
fu9dzdK+s21l4T40RIAvN3rNJtCTVWnD4inTrgi12NJj70z+BaamWTJAUnzjDVGy
fGBqd95LF67Uha5bThKGLHXGXQncGOmFncSQwGeyIVKsIv0B8V4Irl2R6SQgbWVj
CsCAPbnjBELS4WP49oecSIS0kTKH0i/SC5UBhU1Eww3AROjM1uvxmeqKtGhNlW7c
4kWBFgdAnbBqZeTmjDIIWBrId+8sdTVB+hfoqZMffJK3xUDgDj1lITHHo03PvegB
auG3bZB2uWMo7c3TH8SWBC1WWfsOAqLdYcYOcIlT1JMw1LAazBKA4vLrYDVGb4aJ
Lgoz/VRHveOu0fFf10SMo1j/VJDP+U4N8vlDEB4uKw+A2QjnKHHLhojO1QrROFOO
gxFpmJBYZwGqx1WC5B/+zr6UKlXO8k/lzTZFZE+0GmNesjsaAELBDiFoCOovEgpL
IzIO0sIGIcpkNOvEb0yPAPF2emMQZRKJiWGjXxztwNDScS7vRmfucZjQmBUWN4eY
B3Ii2Hg/tJb6qPfWM7qBxbEF96l9CfBqSr+8HnwmwtxxKm2HVcB5YYLRy5vN6i6W
etHuGw0kn/fM/ZkwsTNl+/SSuhujHOxcHXpDNzzReIlg6M4d4kFD8J59mPiB5tGo
icgy1OlOnWEvJKfrWHDe17DBlpe4b+BowTuT7LOiiTTEYO+z3zbplcuC5eqfIEJb
PRCFyZRaVKraGxfeFYloY5CaFImyQEs21ryHBdzF3Taqqz1Z1GMLAQjeQoCJRaYY
9w/pbrcfIA8YwbRv5eaeWTI+VEu2Y3ara9zKLyOBWttf4sechEQx3RppCrR1jFzY
qQxaQjkQ6FZKqbpcciMC4Z5WO3zrSQr9YfQ2/JA0Gu/lQdU2WABsOJrqC0mN0R6P
+75Nn5+EJPk6dWY6ifqlgOcYuZ7gY+tGpKWcThBtPMmPkbuPtqGqSbMdccTb0mYK
k8IUFmL1uQYpq9L5ggJaxoIcTvF0fHc1ZHRUHoKon5IMVQL3QxMrt9Fyea3HH/kc
LPWmeT8+Jfjbl0zgsqQm4fYe3HK6AZOEu9aBibO6tJ76XRudNuj1qUGISovsSZEl
l4wOHQwJDRIAcPXMimiTgYMXqqWvV3VUcTctnYGs2vO6fG/ccDyzR7aB/N6sQuD8
1pZOcpBBkbaKrlMPJYc2snZk7q6/9pwU5HouLeSHFC2Qgody3NprGW9f3srlkdon
INn0PHWqia0Xe9m8rzUqzOtUdb6673JdxPmZM9getQac+ETbDRxP3GaOjVH8zXfp
NS1eryEa1nKK99CYFUx4XaNcRC+F98HiSzwNwtqC48vJ81zaoDbl0eLhZzg9REDW
G/V1UjXz20lPVYsPJC3b6t2tmKe1u9AVoyo5pDB13nrr25HmjaSzlSAAAttl9paO
insNGNOAezPugYBUFbnq3rUl3u31uvD6NTgSZhKAwZ405yi42YbqLWcorrlPcRSX
flwUCCL9o/BdpiD//o29lC36HB1hWX/wqk9dauaC40YYwGs5Z0c8SfNYmnI2/p/K
cXtziARwZn9qJHqZR54N84S+O7vLqxZ7uGCyrHDmb13LPwrFWvNa92LBJcVYak+l
NKjTTvxadSxRFrWrCtQ+str7pBHugx69nziTD2haBbdeGbJrT1aM3ovOVOh7O53c
JdGZQh8ORx/ebie6zTOjbZeuL/KImYFtKYJiGp0rGJgO/slaVzpNcSXWeD9Tq7FA
zCZm3PnEMabhzvziBrqokbjeW8EhnfbWtsBVPCrlu41R5a3onIglh35npNL+CvTB
0sOInEcm2j8BDnzW5Oa9jjLmH8a1RBFfaDTs+x0tHl9V/+5jbs1TyQRr7oKwYFK7
5/RsP7bG07b6j4zav6BqQ3pYjuoKurlgN92TmUgk/KHG9WW3GW63EQa0SgN07j5S
xiS/SfAc+3C+szUGF4TTzP+KZN9Mlfee+ywgi2w7h77ERxFVKdedxKegBkyDHez9
OfvNMLVqctf+QqIXx9GBU1X2RCZWVQPMzeIdfltoVrpeR5OMhtIC6qL/DCYpUsLv
CielKo2nbrXVkFcnPMs6v8q3r2tsFcMPni8NoIHPjos5sNcfUqjARg049PW338Rg
66DmM7WEGOIrNX4BCjzQT+aqx3FvKliCk/4CSkJMC4PXG4kQ7xh30AjC5GkK1jHy
UmdfqYh9RHzv3w9UCP06OLxGqqKfbQ8Ak6dpJEbw1oCvuN3kqVg4wK3YZsswzZeX
BuFRNA5HEiUUXZquTh3ZDBhTBEWpRbOTJ7xDOKfpCKdzfHZqtbrZqd5wxKydv2Cg
hmeKJhVhtAN5Gh2UYemPovdFJ0L3ZSj+34VPHBU4oz99JU1IaGeqvzUboDz2AFGD
ft5JGR7PQpLvrKYCGo6FO5Ql5RuOL79esuiHndNxQRD2ugaP1QJ2rxsKDjL/kv6G
eSMRBAUNs9y0VWeb8vLk/+PSSpzgFycPZYd2L1QelZNF3X4Hfw12hq935SDeosVr
NmqzT4ABWrzOcwJ9hM6PQFYNNLCyd1zvyks4NAlTZQDi8/ZI3PgYCYjG0+2mUOxY
HHjqomUX7W493+NfKt009AWL+B87ifPy1vgUle1nytsshvceK8myqU1Fk4gq4xDw
79RJ0/ScKO4uIuJiqoKcwsYcs/jjaScVSHBack6kRcNshBDzI2hPVEC6owxCNReN
go3cyzgflbPLG/263C+Gu6ZtpLT1eLu+Qo3+DXcYA4ur7wqLlv0UQ+n8ne+M0hGh
vIgRiB352XepzkR0wNUDlA90STcJ7WEYCk7A5C2hl1lYj8B4IyxJmR2ViMHdKQFU
2j612TRMwxqGA8KxWEXsCznHU0Q8Vf7Mlt+RbHVS8H0IvJqnV+mmW7qScwYy9BLQ
lkmXmLB8py4zdvg4aJ1G5KmF+F55dR/it2nlhQizuMovP3MFiEDVZ9zvbP85QBPj
DhS65goJTR9to/Hqv82xSkeMjC+/Aoj/AgiWACXNgepoSCQ6iFpS/RxgPVTPHRD2
ywS6NYvNmZoGFEm9HDeV1J4VwUlnD8QBv+E8buhYURT509ccleyccZL8D1qdA5iE
n9YW13cHg1Cp0LZlwyTNvVtw+GK+QEau4xA4dwu3WdhyEvZ24GEYoS3j6DnokA4c
XCktmNdkg3LmyQbhltq0bpkVNJPZ9l5jUSwmLehH+UMnobaPhCnX7CTqcnn8rvMm
jSjg9hKtTU9YAZAGsUvWMpfJ6KXpszsrh37I5882zsgdC+RbLGaHRYKyGjEauvIm
CaQNVODet0L3ZYCnGM7q+IIAGQZ2JPg2ID4GZ3/uUbnFIDU8qIhUGU+ropfeHys5
eDUbxrJNgjqLROLSN7iiiIF80/GmUmGtZvnu8VAYtuZPm0uFls9hwznXjbPQfJ5C
hZnM1HTWNshUrJoPL4jH05p8eiJXK/yqi7gDuiSuvjN0tolTtcec8896A6D8fS8F
MHeKUADGJQrA7Hs8TfXwTZDyGpTSPI2sl13npPyqZ2q5tmoorcSH0VoPSE79h0D5
PX6QnqQvxFqs3VaPqoo8YjBCN3tcR/5x8P8/3//um4O5f0ovE2H28y0JdQqpK1Ii
66tlbQJtBGcMXArt1BiZT/sxCcsKXDvvdPiMTuLg/tw9dZdf+hxPvUyrU5u4FFFf
nNRntL4N+2RbhI3caShh/AXi6RogB73trJiaWWltg31zi8Kj2Wj1LY7Kt9iq43sf
NAlI3nebTtmAr1jVd8D5YJg0WVOmhBIJw8SZttSK+qWOdFjoDPzQ7QC3lhwlzaF5
qGc2ehiOpwa82zVlCA+EzKh5WvAQtJMnA4trPAd9ygD5yyAJNqQDZAq198xt/O+x
ryQ6VU1uUpdygzyyZSqlJcXRealLWYJgqDd5YsSbCFH3ylZLAe5mI5F/FzhNErTd
aGZV65+g9v7dmn3QNoVf1AKlpSIPsHD1M7G9VTJtBPoM1KdpeFCxmE+IgZCqCIth
Zpzj/g3r0Rxo+THyaOkKKYvMTDrW44gzG/6eBA57u6Bi+TpAExCCuYlHJQyp/tgK
o0b1hShcS7e3Cyy1xQ0/im7kzeIWxTlbGCTTkev82E7T7avlBhMs/1ESjRj+Th95
dYzYr6CbpaGHkwB7WbNeRI9s2kp98xO1TDNw+Hso5yge5/GKiHgHhD2ECtt7jWaZ
4R6tq3V3+bs/a7hQGCIhLJAjAVHgSMXAW8u6DLIIS81uW175mQIM/dmKAqBDCLYP
G+YiJQ3Ihei7nkDQqWSXuIT+DD8+2RHxzY+9fepuTYQcRLTxG78mRtn/2zMYdAtZ
2fbYWK+CoedC1sdIJPk+PCjswYkihLAbfd735EfZhM2O2XuMQwlXReNXwgJUR2kC
xkz/qiWdQ3APQv9z7oW01opVrKebJf+eS+GKbmDlohAcR0XzgW5pQK1HHBxDnWRb
Iq8x54FAk8gkn4tdJckSLI/F3gvrMoFfkQBU6zt4hHy+qMFO4l1JMXr2FA8iy8zi
D2cpjMcvD2MaAk8ZIcQyY/ZcgWQE6pOil2qJkKUBHuGlxAi0Nz05nDMkrwmy4ixH
OT1Y4NPNZdlQb2naVhsRVV7w3Pi3P8GeCigchYMSkAZYy/I95yoMonIfHbm0QWyX
Wz9j4aTZwi1HqFO/M9BOSKpBD38WLoznLgEXV6VmkWMFFCsKXk/J43+JHC53oW6/
BycaY3rEAcrqxsXZLjmjw9ixqblsbppiRzGeA5TW5vf1oBd27mTCE8aMttPh31Hc
ggiOaKn396EkqgPGsR9TpzbM8XvmUHo41I1xAj9pEiPM0QiAX97e5gIsc3z8noH7
91sy8aDOOlWbQ55ARg2+PKvAzNa1G4yOqCMYAqNY8HluXHPbBaJeWubaunNtqS9T
oqbauccZ7lsjf32MhzjdDSfAiri/92liz+XAX+Z2GvDdSUawcHynkFXUyTy4/EPT
ASxrOsM2PlyoO8M+EUaegQTx+tirA5hUJ+u328lgGiL5vV2yV4PaO0pBIqfGU/75
vSiLz7wVID0fKtg61JGTakDUoXbEOYYt6wQ1Eak8WQ9ao+SLSEnAFG9xGbhWnl23
W8qIdKhJy5Iynyb59oPhBvafDIx4okoClCvnn3gE2RI6XcXmgwKMsqcSdrjZZqNo
sEpvdRNVUcnoEFZ1A8+Xk2BHdzrfUXdni54V3QCX97fvEhNsZ7rU3cUYwzd70TK9
ZOiwhXpbTu1fE3/PXMUqoFSqwqPH2hrchUZiJbjnZNyD1EFa/a4OtGyeKgx4kGfc
bFxH4Wd1gQsL4jAQXBey3x8SPVgC4xz7JCn1ec5hJhOiOyfoNVRP36LqbPhqLGz7
yRS3AEwzZDi81f/cFegDcdODB/JAbNgyRxnEiN+SLKwKtb+vGDfz/zS3EIReuAHz
IBkCq6OUxybyFu6Nxd9Wo+zX8K3GufgLOPOTCWoaqMPotT0JRXicMJyvLxhkVfzR
WAQtK0phVbu0rIVgvDumrwCHZFZyDuEfsIy9ZSt+2BCBZgusimGV7XxeA4lfOtfq
kr8q61vRmU38OSdAo14vbJbk7GSFEp2KEfdL2pZ74kN4SYDj+RXg0nwkJqHjj6B2
mjouMbQ/FGTqXza60Cp2gjx8HDut+xyoB6oFZtsiqcSPdbKBTwJdjVljpQ0wEAXJ
4n7cfMUMmN70W052+YqRuptLSHJi/uB4JvKMsO9LnB0eQ2regr0S29LRiqxA0KZw
8bjrFRrhnlNGg5+DMvFDshyfRuT/r34w2C307a3VWsJ7fZJxdX6dsg1ZI3IXG4Ah
Ejx1V+55A2H4arnzbXr/cZDMfTp/G+iG269CUTKiO+5KIktG6uWx7qO0DkolP8Zn
vQy4xw+QKdWo92W3N1CrMpxrZXPeV+RX0Wlq9KTwgIi+02NKoPNcPh9tHmV9z0RK
/VqG/tiESV0weCNpFshcaWduWOJ1UlJznUE3QXGWnuSdeLkZjMoPIw3xV0/S0wSu
fJSFqQ/aoUBV5XatYduETdRyzNBVKjDq+NZ01+uewtx3X0wsbd+kYPU3lghTWDl+
+eJYfzll3/JV32xoMlROSLIB/heSwAuIXMnZP2jqkF1TyxNo6xZWJrEE8qumoN5L
Mk7se0ICBOCzIE+c8oP2MA9/VZfCGhdFEQGLIqI5AV9x6+M01d8FvwYXW/IuCgx+
X3YWK+iMPBl9F1/awNYjZH3aY0kFGQtbvwf8FLxvCO+CqWqkEYDPwmf2SZpjckGe
XIXmtMgm/Kz70t1VwrzQ/7eFmCSsodGCRGKML6C+OrfekbM8mJhJE7LTBhsS9ZyB
qT8DZOahASuK8sENV1W8AsxH56Zr4zDqpSyU1MzVu5EUhKY5eGRR6G5MTqUjcK9L
vJv4Vs6DRvvJXjjdDfw/cIZ0uR4yARuA99H7aYsmXaH9cxrHs3lCfp525gFRvnER
I3WVskNb9P2pYoE+TKfELO6U1P9V1ktn8WjNLtMepX5KGkl7yjkD5leBCfoN/xrA
zw4pmw3+8rGfPkxZFSsZ+2gW0TETGwZaExNiaDD50Qc13MfRru9+QRyaBGU1a1Nq
XJYmyfs2wXTbfkOxCTI1RDUUcVG0iEt3xdXbJVapjkiOxh/HPqTTDZe16wJyzIwQ
5SEp8B45sG6X7pUdJzxrrTiu8SLdJPJ6GY+DQQuZBn2hJDGnAYm6tN5RY4yrwkbx
I4sg3/mfiVC6I9Aer3ThZ6fWqZFIhHQHbn98GHcYZ0RqOuYQsCPZ0mE1ILIsRDhx
JR3c7GbNeLg2ahdojBuZVLCBgnt0647MtoLuSh6T65ChD20/jEpbF5l4tG2Owc3p
ACeNjft6U0nGGKbmDquqvs5xQUYwFhEIkqydtJYB+DVJwm5EmjhKJgqp8eevGTjl
7rHHgG8NQo/5HZk/3vrNsr91IXhCPbYq89GcNxV2Nzv0C8FKui61sNkZUAwiBGlq
fYIoVqM8p04UPObWyOh+foPSECbE5w5+teGg8XVoP3SmzF6esjFh85g9da9l7Z0p
O6CcSs+g+DuL3c6HVCOF8e5aa+NVukGLIXwETH9s3RordcDUscpSa71yzxf7nmpy
sSK9ckzbt/VvfBbL4vDjcfkVIk6/E9/E14cRdGHN08pAhhebXJLtBprlslQhL56A
rpRqT50M0PnXrd8vwDaBOJwEGEIG6V4BikSKpBuxcJShX7vC7f0TnfunEBFqG50V
bgnogr5zTOwGIvzNkJR8t8X8eVDeFL3CEebndNFfptMNsdtsWZ5xeitWk8HYjJSu
kNhtZEgMtjIYadoq+fiOB7Sc6YrAVoCdFArNba3Gz66wlxJKFhn+vsEhMkMPbxEa
Osys9DrWNbOu0zXBd3Coj187n9WpEv73/LR95IESsSkIeK8yEB/cDEq81xYTRDUd
Nk9GrvPh3WaW7uzyP6mkKnxNUTJt2Np4FPpcRRoWy1PXTAIQdPzxS1SNv7gf+3TR
ve5DhGSxe7Ct6fFpmJoFzMz8rlkdjEyRvfikgBFjjqTeyNTKwrnPIj4OrpnGXh+O
l/ULgrkz6F50XBQaauoxzGSJxbUr0ZKETt7gvKeLYqRroF8VrffNJGSy/nTL9BtV
ncKSYRraKkf5tJ5FIrA6UR27uNyqLVaLcL2dPa9shWvktfi6IIoYc7WJkdwUsVxO
PyvmVBbWgZ+TE/CkjtSFlbAQmxIb+IiKHQM7H6T7AnvTEZIqh0eG1BNSjYr9JfVq
W8DFC+cpmczDhER+jCBHZcGpxXB+HFugWGOHtyCjBUPf+rx2lXq4oN11U/MJewCr
FQv/KkjTTTGYSbmS5hpi7hfChGVFGzoWpytMvOM4q8U0EQTpu6uiBERYHDCJEwXB
4zk/rfSXyzfEpga3emH238snYUJ1Tu5P+Fm675lgz19Zk9xQ0DGxTu6mBTiW8wo4
fhWwjDM0L4g+YB5p/ht4114BEJedodb7ftTGpKqLSfoox6+B6H0IkTR58YSd2hzr
PTXrxO6se5Q7hqF9Ci1TnpVRmcnmeVfRguDmaCLFr+PFN3XoKFzcXysBNqbmYXyH
6MmeLtFW1++T88eH3sdbUuN0DEg9Aierl97/26G+VzgmzaxAnvQcMQrrIIdOwgKT
JFlsVkxXXoSnSV/wdKyEYP0D7Lwi2rKmRy5pSDxPlbOr7gg96XTfybvJSvBVGNDh
K3W2vPpMh7UpMF1xRM9elzJ3PuvU8L8VT+3DRA8jStxE0RE8EsMQ8lU8sb3IMYL+
1NZyRO5MhJBSYdU+ybOP913rZyv5zEIDC666iJWFrUPYfgKiNmKNbrTPKEnzHm+V
r1TaxjXyk2h4MpLYGKXeUB/Zl5Wj/VecXlVaMrGXkul+exF9zlxZQsD0+1p91zFd
iLl/Fv/wXkvm6DYaaoZwHNPyQ424FjN9a0ZEI7q3goDlEkJgUdXtF1OKdgHEFHDU
hhxiYIi+TE0xTcjfpf8alHcluPDJQ1B1OUmZHZXuQkTYyp/brvg5OYiPJqiQ1Ui+
JHK05B4VYImpjIflE3N1k3o/BBqX6z87WN3126ZncKBTJISAkPjo8UeZP+eleAP4
JjDFX2gwvZI95m6j97HbyN+QfyUuvytl9HONnaChjN5FZ9yjArfeWDOGNQZUjy9G
cVzYUP9+1R6fLsl2PGrA1vlsC980m4XzKpQbnnDq9S0y1rc3PNiY3ZdPLGzrPE15
H6zXpVWhRqaf4MmCrrvuXomTtCwLXd2fwoB1vr30HlFh8Wn4uRsgW93YYu4/Lyld
HZ8WeuB/q94j66xqFvUYyhPcX+iAOe2J1yEtQ4O9FH1Lts86O9DRarmVNqCUIeWi
LZNHx08dU0JVcb8ochhEA3QIQcAiVrJb1EbviuU3b/CDTabE8SESMHlF4tezQisf
0EtK12II32CxZstGC9LvvggNsjgUm5Jak8IvnnsUcS+k022SGsskuzqQ7BtZ9vA/
I84TTAFcaivzwNJeWWi1x859Y6/TdP6EjrrvLiRN5fTVoYEgEuwLCrJZtoE3ehmQ
GQGsVxdPZRGklpcI7UA5ZPOXDEsJcrTp0LwMlx1llUTnz6DOL2rFMQGDSDtgtoVy
MEFlE8wsolqOqeDWyctt5IY2eTgEke2UaLlC3sAA3+SJdin3ITAuY3hcVj4DBkL0
nedwVPnjBWQuKvFx/JmlLoiibReXCQEuvbDA0+zAEy+8PQXOOoo2xPmNvJz+p3Zx
sGki0o4RncDyzPmssXB3erMp/x6GcJoSUV0vnwruaVZQmEfBDB2+t/vEB8dji4Od
/E1GkjY/N5Rh4JorJdg08s+6S66BSCZFEx6ZBfoYFy+ntkD4Rz4Iz4QBOzlt+JbS
BFUSEcNG85syehI+uKEsA0IiEpSqlqJWduNqxh/CY+voOj/gBP8c3JDo3znAhaQW
DTNE0pQH/kky5IXomRgnePoHN6CzUCZw7qTyBzF8dZ0o9sZhXsbfV8EvzzPpXgZp
TbH5xgrvGWJt8VSYqpa8KvuSv90J+CfVP9FDZ3tG/ce4Io944USahhE45PYtDlEF
8SrpLFkZKyZT9fZbUutVRn7NKbbA/zr/MZG9GMXjhI5hIf4eK4NIon6DHlheH0CA
ZoKuRdInzN2PWC984KXOqGcgXnyy2mUXTI00Uo8Yze79sI6740VAUz1OQSWNCOuI
i3XNVq1f+wb2Sia7qLrIiygX8ndva5kYTMi22st+thpVVjLC0KDJ9XuVvI+ZGKM0
QykDP4zoEoNORyhJsXo4BT65yQdB5Q1Wn63TKtWER1OkYs1ss2JCYQzVXkevcmzl
V7fwlAeIrdD/YTsgyu7fFYMACO3o/0iJWRBTacZefE3zqW3rW0cm8GzNTj75JMVd
CI32a7KoWNeTS9cmtnBVHr8XlhAOuc+4MRzmNQJufXHWeyKVbkrpd4ZzZgh/wrJe
AzvizP23egPXzZz86ZpCJO/tNSR1cscn3nbfTtjl3PPQZY/HhOXMYBDW1EU4f3E4
jIQ9hRHz+UDh1CbmP6cKYvhipLlebS4zJpnWT/qNK8QkYwT7caS0fnegdBnKBPrT
NZ0mGT+V69ppNazzr9bnyQCy3vmTWl4aBr1mflWtU9bQallYplZkzBUuKee7W34w
ceIl1Xhhet8/CiwAjK0LE0MNiTCmdJEWPfv8SaMbtdledtrNwoHO+o5kSz44IRaW
EDXXDTj0tZ/5RH2ns3MAKRgbkp4nNquh/K4ZRsd/8W9OylCZP3rpfBw+xLbkLsBO
YlJcXU2SpMmeSESKLR3KBZFyNTq84a+7K4X3ALPlHOOA+KppRpLbEvx9wsvvtaH2
rrVby7qNIK5AH8+PtYz4umg+5hhL5KCoaEflJ7WsgyH1PtbKJVVLVmELVEU7PE91
GUQoWB4xqj8RO0X0CGfELOxuQr5ABFvvv5mal14fyQs/qUcX8UxzIUA459NPx3q1
nFjGM290NdiObImjcJaBORyNLFXulknJevodc8lQ0gYECmMT+bTsTmJ3tEdiDA5B
EBU/KepXiWsSLJR61YZXjeviUfXXvyLv9xjQX0Y2KPb6uNKPD4F8p6DgEGWdmBR8
v0gv0M3qdyq4rDo9xksJ3M1G7t6ysd1Y7MVAz0s0oRY1wDqnNWdIbcUP6xk3qp1a
bnNwff548Kt5g30TgLzSXJRniMx/uXVQJ1OHQQ9QQ/jgE6q3qNO5pWJBJwe6+Nfv
Q39gE+KaXDNS8045ct04kHfPJZAg/HTqBzyShuc3E7aM3XcT37F47o1hvKLoeSRn
qvvNy44AHHbUyP6ntcMHkY/nkcrK3kLucVP908j/PgxD4lxOianB8a8uIaGUm0Jp
3kPt04snzzh/uBj9mOcBsMbKB8/8+dYbm4scQFUaRSKph96snk/h6tLbb0jVC+8r
P5qKzIgWYTqhHov96nqWk5Fh4tPhosmqcwx7/YPTZrPQv0NVQGxnZ+WpOA0jf2XT
j1iQxp4XVkuP5e09PzKyoSpbeYptqRWnLMEU7xDmZrxXgQjyOE2lp2BuzxvoEZ3o
DSvgAUlONRoeFbfRVdBKib4m4AQJl2vSs4M0jgm9hCjxAOHFB3ZvQxWSMoWQ8Wkh
3iFHL2URFA2kOCUp6CK08XwkIuwxCnCm1Sge54VjFtpZtQYMqCrkcDQ1a/PJhrUf
JVApEUtFOSbTj16xFUazWrzD4ozZOnr90QhpEh5xKxkhJ2QgQ8RAm9n21BB7O5/O
DfgWERl/T5Z34JFLMHsq8u5rl8g7LnjBi01urFT+GNNaQ8kPp/CisLsCOzUlCHlS
msm6REw/cGOzSASmxqgFIb3A99ZLl0APwS4wd9tDIalQ0m3Z/lJPbeZntFZz7DPA
wLes0gB1wzdi+DW3C+jgJumvPw0SZALZ3yYhHREePQM7v5MnF7YqlUwd9cRNin9p
bB/7Wsk8hDu3Df0GpySEDt69vUmFWV+QYKB9T77avcnQEmr5FXFnIoIOsxmFyjjN
X9CTpwWX+uEC+vtj74OlOIe1hw4Y3s6C20duSe7T52EYteY32VthiKl0upqy58IS
JAWq0NFUUAQrWrkT+GS3Atim3JclqCgM0Vb7bJb5hVyEaonBU9aJ+d4QQ7Bjc1Hv
KCtHa4UfqbkQMRzZmsX4j1WbePX891+8xapWX7yVQAKDekSZblqYQgnyca1o2Hhx
UbRzIhgIkeYt2/S3ZZZCh6L9mzm81fETAJd5vOAeRk7zsLWLzzVG34LjmroAu7Aw
Ig3wGZGOxzFRDBW1LqRhMrzrdRb5dEOAE79ohKc445n7nFQcL3YyotDpSagrMspt
cBWhhP8FAT+yKAQ0x+z0Yih26dC875r9Ma/QuZUKY5JoZpjUPedeeRqR2gVG2v/D
dym4cluPr5wyXgROMsCh/cgxqxsRZksGHjb8ZQdFArWi+dbZ9qE5IJ0q+nd4kkQA
ZPdRJrF31G6+flIUX017a3D+hjCFcFFoo5I2WGH5lHTXzWqdzPtqZNQ6tjjkVSXZ
8wjSFrBsD6AIHAhRyA/CGVXG67L/HdYVaBvX2qpUkhvZ4XS5CBg+/eYdssFtqBXG
eY4lc74j3Wuh5xE5eqrnfgMWMYbTSaR1RP/FEPka7cuUSVJUBLYdv3QUzMce+1oQ
0xUvdLqBJ/ulZZWvL+mOiND92qAGZP0n+kYVt0c+/xyF8t7oC/tZup6e4YnztdFP
1eB+Qdf1Y66CjMq0/jbicaf0bjqJA2pqCt29sPUD8bVumfjW1ufDMv8m3UZr3yWc
5JtB0aM2Zdc3hxm84AINueB0A93uH9ixVkkZg8yHwI/Aav+myRyJd/f93xPuAW3O
gzYLKdKuhzwOSdZ7go3m2Iz+jjcgDtY7TEYDQFO3jGnKBg7qYbBUrxxx61NVlUas
L1/LsfVmeLVwvntX1+iEw4em7SU1BF/aJrucOIgc5Df/ocBFpiQz9UGoRbk3ECgh
nVlUGW9jDVUN+o7hqNAQnZFu2Y+Bz0aZlhdoBq+j4bo8encHnwOB6x2NqicaYIf+
gGdc7vaChY/bBH2Tp/0bu5HGTZyWlGyZe5AFJzmmA9s+Q29BY3pH5NX7Axq7S82A
Rzqeby8e4nt/Uqk5h0nIdc/8oe2sePrHPtGv9prJMMCRpt9987QlvODoCuhKZfHj
wbYHrYpI8XwImrtezXKeBEapKeBeLV7WLdCxPg4KrgX6gy5qBtoSjRpOCntbb/ET
62Ks9z106+lww0QlJtEqaTL4Df7t/w4KAlxKDwlMQ8bBWgkY0vnmGFsU8Asd0o1S
LdYEhQCjBES/ucPhzhrQ9Og/Cn58vlx7EwaDFsW8vGjVGmLs1g+sVAf0VFyizlKT
bBDR7AKYfq/VfulPZHiqkQxxea7jHO27jvWgVuVwteVIq9L18SewVTj5ZqB5tzw5
UVWlv73lfFN3j66xvRAENQW2HAZJHCigdUwWq3FEFWx9nIkqru151y8XEdylVvlk
ZggonN3jvt3hcENXEjVjk5d5UHs6SHYYmShvzFnbiDJFv84rGMaCSUZ2uim+YS3O
h3txsrB0mSJ5j+XoC/tRHF5DbnhDmor/GDejL6zknNK44bTcZllxk6ad124AOA2t
3t+66f0MiU4LNGEOXhT3A3ZRl1Q8seYflp+aDRhTrmOnip0q798+vFGej82vc2Pt
1dqxbicDnM4dCBs3KYoQfJ1Iy2m3OaUhiPreMs47yLUpiXVHxf4lGYncGyIpae2k
XIY3mSa/OVhhx7XGeZufycBV29+5Kaqzp4jvsifVe4ugT5g3OE6KTPwUU3pounbA
sJnY5BO3zUvonMMuAwrCv1K/JOjd1DL8CrTb3ZKWvTc+fyNW/DYJwU3facx5a/1/
hn8yJNrgStcsG/qRKkSktkcyyU1dBvxL8HYM6OwmaHRz6dNy9fEZEbOoevpvUKy9
U/Wqp2027d1fngmZLzNrBc2/Y+gff9ZCoN8WtqsVetvzQ+zovrGPfjsooXkxfnZD
fh+P/xrujYSTe1+LV/+vE1axv8mYt2sRDhK/oQrMpPBk/tpB7FkdUdtcn8Nz44hF
qQ4Siub8B5et/NTzyAacXLhEaPvD4rVj9Hcduq6k+tVCeX+7R9SU96W1jaOko0UE
5Rbr90qlYrN6a2kjM0MRIdqTUMIW/kqEW4VjsLyqkS3KLDl9Azzlty0kk9ISVv9+
mSENzw98wU4dc1a68YmRTCaMnDZTulu9kSrcd0t8BgbLOG04TPNwgExkCwd9DlC2
jb454jY+SYT+DbhA8yluaunnvO4tp15hjAZqhIDgB8O5be/Ccnsi8oHcFoF10UUx
EuxsHFmMcieDjT/w2ziqtz3x2303RKahSBUnxwUaiTOlgXdWy0DKd/7xFrcM74Lh
O2/cdR5DierEsqbZEKT03FTsTKfG+VN00sC/3Pfp2UcE0oPwrBFvVCNwEvGHNyV/
XiZ9xDzO48K/1WIUOfjClNgSa9g1jOZWU2wec79o/6/Nsi0JWWRJYUsjb7hbMyaT
CGUbIdspj+m35/yTngHSZxXL8lYP6S4vdL/Ba2o3rsjHR4lYGpiNU+IjxeFDtD33
BrhRXQtXTm9Aei0l6Qq7Dbra9dp7xQXa7yPsCvbFW7W6an72kkX1/iLECdfWI9cl
jhOaZdf6MwkYor6NCm7aLXbzdwyBoaBeQ8z3FuDMJyRhZTV2KWJkAENogyW+ZthJ
MMZtsHBiQqKQkYf4gWaWyRy7VPjCKplfTtPQBcEfbVNdbGEh+kNjwIttuN7vmdZt
U74vYJ7JhbcQYaz4W80jANekRvcloARVlr4w9GQKj8oDbrtLEwPuqPOPjPSeKyhc
pSHcCU/uqtSG0c1LWtqnrwFr9lGqNd85dM9wBh11ufGUZ3E8iiiLvXyVmK0KS8IS
SISeaIdv1dz2Es1Vd0T804/TAC1y3p7Ny1fbMIhWs6aDP2izQX4EYSLa2Jedix2I
Wh4MyfmYr/mxRIu5Nr3CxgbKhEZxkLG0sx2WuF5yHala9DdlHvvZUeATgjeIRhA1
ozjLvkO4sooJBN6OwdUMz2FE2kiiIr6Q29kUjODR9+mNqXw1WtQaNAeOTDzjNI+Z
7JHN2wdeJb2Sv5oAt91OoL9X7gsjxy4vKVdsNWiITrqZqNeTAJjbs4JiDITDkwC+
d+yz2dwYnnXYgxjzAge3ZBdyqfP9FdfNUveLpnG5E2zhVSYRwQW/npgBITfYK3R0
gCcmr26OJrfHAK7hWgiMnqR4/O+9OeuOPwC7Dw5DX3OiZM8bI7UhAq8e4BEL41QY
ERWRz+fle1scL72IiDdvN6vIyzxolUlheM7P6on5/TSiV44sQKmDCIOkkuF5QOd1
XghTsNMJfh6OmBy0iC5Cz+X7N46KWoVyGrEpj6eOlR6jV5fWF/Bm81RZsNicv59G
Ah9bJ7DrZJU0VXyO4HYqzOiptFsvAmRGAG6qYqZTr/z9bnMyapw57FtxXR4408nM
O67xHFMoINiz9Q9enizjeybjdiT/K8zNhwNmLm8+/6N2hicJqAvgxLrGza8I16hy
7atjCFXSiA9nWp/JOYDfZoimsf1CEluDPMjL+X33pYmWFZzsYZ+DOPFTXb2PBEcy
06bAAHzeVMKgHC7mxRYJVvPtXv9tOE+RCk5tj2ixfbKKWS5/OVeo5aaUSgXJd5dX
SoF3scQci09Uf/THP3nUdUcLekfpyvDIGx04ihSidLjK7NXkARbPXPxosd/HK2Wc
bvhjm5TbGsTI6Zi6ih+tebctiPIYOmQdPhbIoiXt/hC12Hp7Pov6B+58/Ej5c8nb
ZuVc4N30c99faRSmV6bobwMfqf6Q/8fDXdQoPRmyNc6SEa9rs+lx6tGpd4R8v/09
YAjkn1jZ9z0qNY7w3ztTTU7U/6VKpKbM/Vfhb2J/N5XIg+byzvBhMuyNHXnIUPHF
oLpJmoXzyn/gphdV21FZMOkrLvsmGROxlFIa+DZHqs95ZXRy0Mhwusn6YJ5ZozA7
+NnX0f9UblEGP3r3ztaeVwi9JU9Cy5Ovlobbne45Cu3Rdq0IbBg7NP90ePT6lVJD
kCLZ+BZhnXWIDuHv98vNzdOHTlSLW2MvIoqz6g/PKB1tjayNkQ1TIpLwf6+sjEnf
cV3qilvSjRmlfu91Xd84Rkh6+4jl+lOE4yuFgYvUzK2EwWApGAEr8JxNDndy3etZ
VINhHdSMWj9R7hYY+0BHDwVL4KyuVkU2HQ4TR/2kFipO43Lp1sY1OExMKG/ahtkr
JG+IEuhPBsb5Rc5EEYrxDK5NYFBBBbiugZKNQO0CBRJestmHvKG/jLnKfRsFGV3s
scr5W9owVJXOQxVeVOkbqe3Q7MRPT7Oq9RX7wP2Ng/m2o0EFzSfV9QR9ZviwU4Wp
gwdI0mnVX6ay924tE3MHO7thrP6G21d7B3L0IGwYVlRVokQmr1g4uxpC0cE6xcR+
XZjTXm24tTGBsReOraRC+sSb+QUwdgg5AIsUIw/Qp7SoWtBs2HVw1LF4e9/gL0g0
7tp2g4VFCVZBJtBgRcmaUbxgcj4Rky8rYvDZ40rVQbj7ryAMhjAa908Lmg6+CO/U
zdhJxBhk8XA/ls6oR0CKIerCywGn1lBlW7JwevUUvQOMlUlIKUzbRuX7npOVoy2u
5uUm6m+KThMaQWTq4YKk3aTwCb75L26wS2qfMsm+mrmOUYZ25IxCyvUQSmvV8ptU
5UggYaKR1qZX81Y4kV0tdRRqYfLcJSODpZvw5YBnuPZn5zIkE8ziF82+m1Ba3cUq
92yy354KkHMbHKmWkbvVOstLtQRu2nXTkotZ2OvuqZyV6xxSPwtDWm9V720xo2l3
E+sZa6xQ3mwDfOJVtyY11oF+jNbmoTZse/WAa/702dpoIPoMu2XltDHwnHq+gPR6
MNNtgbHHazl8ooO6btec2yjOEJY3bLHYvo0UNsoMXkjg2thB4sI5xnSVkqGZKW9M
wPR3i6SaOKdLnDXxmG/sDrOsoC2uDxLFALv8oxxRNV21bDtIPVdO+ceAPqlteGpW
Wqbk35URLH+UVoNvtxFTrdUIxnY3rLnxxu+aWmQAqqMDNMRwnsjTjoKQ0rOYv/37
6nirOzCyBujRveapBrhona+esVDCZJHmVg2ZfdVjzSNd/cxSqEKbKOonNPN+D2pp
+rjyHmI79hzHycL1skrP71CYORey+baqfSgudrm+oStHDyonGDRSQ6DWzPbHYfsn
PWMHms8EBxqRbSYDI1FXW8cxK+E4M38hVVSgE6FfcpMBa6339QATLoAOmZidqUCy
e2DKxA/MX1PJ/PHfMdX9M1WdGJuGU7Rse6wTa+y+K3D7zRTk+g+3v6M8EBXlO+jA
h2k2aaTANQJ4yU+rOF87136NzfwuTL8fXNM3KTo5Wgc3psBkbkBFZre8vg7k8t+l
wny4erbiVUGOSySzrJAodAodtpipVigIFJjqw1xexajZoqhgo2X5ce9mXHlSzpgN
tavAdcJ9/Q4/mxsZZJEsi5ZF4a+7RmlEtN6akvT2iKepF09fk9rxTQojUXu1Lp9o
1HgNqqeiFM2ZorJkVX1WYRVuS5fVjpWM24RvVQf/CKC9fhCS+I+/alDmiRtIHBU5
QiungVQBfSyKbLP7zuG9zF3jcthjIWDAV/8Fg5emCFjXENcDNz7W/BzcvlG51qab
wuReDenDZDl6rcBKX/haySA6nOieE9ODYUX23g8XLfO90ounHNYwIPhXMmi2bTmR
R6fNcUOtOdLgozgMl3Vn21uLKMa9Z0k1dqPWzT1Tr05XYc2Yn7VPQvA5YfkbBogn
VQvXQfBOJm8dNrTfB73Z0yKtQpcrICPI+l9haCzux/PdoHpPhvJ5tkzbzkXRQVBn
6LY3Ddk2gm0YbzFk7aXUfa+s/N5+LPcajA+F7y9HA9yPw++7Hqq3UHK3WqXpqVqb
DKyZTakY+v7wj5PDBTLTnYtgHvHp1rCRhLD4lTtIovakAuPcdHIYb5ZJrm0cBUFV
+npGmBdQMyb3wiyPMpxKkl+VGf+WVgMwh7Bo5ygnPPP24fBrvGXSVtbRlp82STrL
gIqN5PH8uh2JnF3GF4P3GHGR8CD65wuHYeAnPLFPWoeemEBMtrpdH+KBrm1Fxlgo
QUaxr9S41aAw1VtUZl7Q0W+HOnRjMa39gH7NPI356L3Yri+Lj5NeUVj9LpzEmyoT
23rDYb393wsltAvqYKxnikZq3E/twr2ewZBrMk5Y7NwAlPGgD48fDAdP1WW1o15Y
+clov8uSKAmhRhRo89K1oNzXn+7SCZqVan9lbYdD25/wKqgQNcRsJ4pUAf/NcD/n
WEGUv1K3Fq6Qfcx4E/fWEaLzU9ugaN7iflMueC7j4U5TDKsYGvS9zqIQDIpKbTr2
+rTPAJKNxtxeFx3vZoPLHweWGgxlK2Vmdbe095kKv12wz1iQKeoCBlhTPLdFIaKh
9PrVkVpSWblJJkfGyKdIR1knz4idMQTRqCoITidEmbQmLyXtOFSaVZNniI7zjkat
uHCvQVUp980hMaWFVWcJ/uNt8uGF9v74OgVsTs9xgQnghJ+8ThhGgpRf7R2KxI/w
+VBoQhzkYSvYKb1FcRD2bSqAFay83LyXsGa2LjERa55PjqMYUCpGsM11caNtkJBU
Axt4doK8Pi46io13NkYnPjVD4AvmVnyHvB9QPsAolyAXa8tz8XlVycIJ6w4cVRxm
YrktZn6aQjHSWYzdqISt86H1q2WkmYgwdjYLWneJ8FbioLwxEkkNsi3/h97GM3Gf
LS88Yimj/wO67uwZEVVsg4+yE8Nf5KxLH6WYhqcUbKk7ve59BVLv9/yDI2dbfvHW
1D/n2RwYK28X9iwfKXX+7RiK96Fpu+PUuUEe6gd2dMg1XUE2gim2qHW7yxkfYfI+
IZL6KfWFcfUzXwYP5obTJFA9+fK6K0Tmovnf8VV6QL7yGYKxcqKzhcvOZep6uTAy
soXWFqXXbJ5vx3X3Maekh/tuUNWsPSE780iDUaxHP7Xr/WLrnxEH/YudnJUBJBeZ
pIa9HimaEL4gkvzoCmGtoLhPKuIm3SMyAN8hCn9ZnguQ3t3aywoNndOMpsCvR1Kl
IPuB5oqBHLM4YSKNKD6boLTVsCmyFVVWgDxrqxF4o5LAMSHQ3fLVrx54N6atWQew
lmJFkiUPR+K7KB8pCNPomRRqha3rx+Xh/WyvGNGEuovDAE3n9CPBRpfA5stYCgpC
P3tP1lIIPNaLN+rdjnoBZQDpTyP8sG/CSGrxym2MzP8TA8c8983HLwXq0AxGSyK9
Fb/+mMl+Th2V0a/4jz6AUxwbB+jx2pIfxklJ76yqPXa7FDWk53E/0ZS6UfsP+H9w
D3fHtmOcEGBg+wINYJyF+Xz2yOT+eNyfQ/pACfb+rcoL/WKK2bZZV18maTrPT+TZ
z7Fd3LW575gyAF2kjYOsfLgxZtZxeYMbiiJ9ELM3LkXj2kwjlR0PCnKWM6Qc+7AI
QrpcVRQLwPFFrx4xbDw0WliP860wX9VOz3mQ54/Ak0TtM7m1AUGDJjMqQYxV9RuE
F7Roa5pw7p8EhgzidBIyqLzJG7VKQIWtVQhB+IOt6bfWV5QsERNwo5b0cOo3xSt8
CARq2HYQ7En4pu7G8bBPFh1c0sxYBt66zpe8O5nxPV60VCN0d0TVNubzOIh4gscS
/6hkqIClUHDID5N71jXXnWB1TDdS60zAJK7KAWJ/lroF/xQYuBX+M09SijiiXhpG
N+27MnFrLm120BYgBFNnYME/vAxAVYyS0HBUGUncsVbITZyMzmkj3U0fKc2RbGa5
+gyO12ScgD5cWbV6A4L7kgCx6x1jp6nxTTAwzFygMS2a+ZG+o14DGFyqSDbpzLgj
I37klhQKwbdgkwPcsXvpXMoo1OSGzuv0nSjP8dZJfJAPNatNxtdCmMKN2Ekn2pdQ
IfJlYmFUQQR3rhVzEaiA8jj7pgvL9D4iL+z2Q2UkHD7Ix7/GaTekxxzkCs251nE8
+AJcDxyo474wLSk6ib2MUNiOKSQ6AzdbQayN8cm66awzCHYJ7DhL46pffBODdUR+
sQ/uYeSx9H/2TsTEAin9KypEWGLqjO5sOrHH5atnqyGN1Sd0014opO7lJ99WGJtM
sxaMQyRRCuU2b4PFhtBNUYwPiGbpMig8bN/aGGnze0MhPxA+x41yDlP8oWB5x+S3
h6H3nf7bxypUo8GCN8ncWVIn/mstIarVQQTL7Gule6j0/erZqyzSenIy1nz3hRn2
aWrR3iJQkdCEXJP1oI0g0vpYLuSYM9fS4Ft4qFHSxk7fTLtCK3EL8JOp2ZB93PCu
VUKEQIJs2quvtgL6l3IxTLVsohlFw1ZUR9NdIErdRfbqSGI8T0zHVU8s619fk+aK
08F5HuX2ITPufVgkz+YmyO+Nt1M1R9TxFNEzVEtLYSwHjHc8O8ubqjvh+EtKjs01
K2OHkxiGExtu9xkQtuQRXjPVKHNPAyue8MsWJqVfHhT/LQ8EGQ4+9HtD6C9mGhvh
BCVPgD4ZtZppo1+X7qG+vut6KQhmXcsBzXrNOlFj7fNvfrIadeBS2nWVCWrDdpLN
5UaKw6NktNtj9HtIhrKexqYGqWYrwKQSG5MUgpT4EamLz5xC5DD4sTK4f0f7pTbV
+ZpzGtZ3vpB0TJ1QPvH3BNqCf/aj0hfNVhl4yhIq72WhjLqO6zGoGB7yu9kw44hF
ixfd8nwSLwpQDzm6oeccOHiuSxysT3ol2x9ryehF8R1E9m4MzTMULkWl/Rq/WOKr
t1rZdMAC37E0tCIgp5bE5Djmjkk1Z4D/uhPOrROVxxkt3zw1K4FDrXpDWYPeh0l+
kCqqLH7jNkAF/tM3S1AZ6LxluW5Xp/oDq7cafMggXoPrrSsyh1eEC/R72yUjex+Q
BBVriqQteUPAsuf1fN7XkSLq+aY0jfHsfX9FWyHcbHqn9tEFDNvEPhHdVA8oR5gZ
alFZgh3yiqlkVlO4715BjsZKbaYAxhK0Pet3SMrXxzNW/wCebaKEIZ4bKT5ttOAO
/fxsk0FEY4kyU7RCle0YgNqZ61xCEjRiFNwTwO/PigvfkvhmHaMDsRp4Ji1JJzy6
50BqX7A7nLXf4uCulj7/Zb/9WER5iqtUrxZonNWCv6uCBdkA32O1LjJB4HXJZprw
LZlnY0U+GwyRW9K+Dx60XgoOPLoWgGnyD/JHvRcCu0z73yfYlIk/IoMM+X2NaiSW
5z4z+7Jfve7UXhayCEiwyZk0ZnZCRBiD476njgfsGabh9JCccrlF34N3eLO6UFiL
Se+nRFcaC/283HBIaOUCeniM7zEnHDHhyhmnyZn9wMzSp40eDVzXVaC0U1Dxqyba
1QQ0qoGqZ3j73DscC9d1f7vZW466QxPSVNcLBKNAWoBrZA5AIKnNeywssd+gtHHX
YM4XYaqzmFk+2DlVI/m/m3qg88PWA4clCxL5HvL8udf7xsR7/5dBwqGEcjipurwq
rl6ojy3y9t5GP8tRt4zB23gNoTkY0/bUHgou3eR1OH1YlbGbOY+dVncV8u/PUd1u
GTSfjDobnKw6bqgriqvFad2h78U8Bm1gmGOYoxZM3z3ip4irOdGjsWDodT38cg8y
evLKIwzg++jysHJV64DHs7hkg4t7mp2pL4nVvIZaLZodIP2UF29hjAhyv1UBBSs8
exQgi3GwdvlvoX8EoWOBMRPzQarbc5k4XKwbh5w6u/pvwr0Q+PlISWaJC/jbLWl5
jW+mfZGYAxvbGv1Pt2cYFqK/QF3WL8+ijjJu4MJftX/JVSg8DgdTAuI9znQdFt9O
fGLy6kbY7G3DMvAAhoaFjQuNrYtOLsYFYrS5Hnzrw1+bY+v1Fl95gIXXN+hoxCVY
8C72Q7Tq4Jh4BUScaHpGgAcy7DoqqyJ3/a8gv0aVHf6xsvniQKMvO+CldtgrLjZE
Nthc+8b1eRFmz0DzuHgPu5gGlUCa3v6gQDJvDf2vXJnf65+lFMVc69maelA9R9zS
kfd2KAIBQCXYOFMn+v9oefojNdzNwdRSunJ18zSbcPYsg9uJc2J8a3NrtWad/yMB
GE5T+6XDku98Yg7hej+mLG57S+NrsB4zp+TqrXSt4MzTiZrH9G+QqzxvwalZPloW
+0LyNt0zMXeNEfCQdgWt/BoyPC79mxtx3dH7rCf7UNtCKruKACrAVO5tQOhmujtB
FHqU1lPSGzmeT6ptOEZsl/PyDRC0zxIr+xhtyNkP1et9xGyFIhzaNbPAUmVm1/dR
mzKsGfbrNCUaFTFjXmpW8Q2r8IS8kzKRijHb8jrSWhzq8V/dJiuzBTSqHLJbva3w
NhJVg9aM03yvBuf1fE35rgMnBORimZsVDc27B/SHwkpi2Ab7+EBoBp9IpkOAmdn4
2c5zyA7ygvpUW7OqlY7OK0SEIfqIWugvUdjxlNSX1ccpmi7IqTtiYgNPiaZ9hSsA
ZXjRZfG4/FL9EAKslCSeLbdhMBCPL2na3BE2SwoMcZImtazks2vbK2qvEV2nKm32
jTCFt1F2fixS9/bORbdvc66bXY+SxByC1OYZ1aaCzKn/SyPlgQSutk0OBMd2c6Dz
nUyt3S22zFEeWhmsy269wELFA9yS8FDdrhDh9zGlM0chEgAioTYacptXkKJ6C+Pm
rpk5fLfvvLNBo6oMQ+DC6Gl56X5pe94Pe7AiUYM4WHToFIygeizRU0KzVf+o9IB7
Nkdja7J0xROj8qaiLzJs2OBkc6eLHYyKld0GLXYCG0ZXrDN4Z43hM3YazDGYkP8f
AVMF4QrBmZHd/oURQjPWd9c/cAMFBHEI8MEG8lLkYp2ESZEAm3ZQfE1x9i+2aeAk
kuqbQ8RF7oFi1u39lOur0I4Bw8RdoYnt7lsgO2y7PJQTcIMD79xxNWCWSlOxJ5VP
cRASjLO5fMviS4GOzYta4Bcf1Ty2jTi4bhcCX1zg7/j3LEPMCBpeu0b/TblBcGFT
iaBfUZvEg7mZu+zTZwLkz4CM1kHYXQJTHgSGk8AgKccD7Fx0nuzGUqVSL4sZTujV
/mP9CzTsSxRvMoZF8VyxKI3UjiaPDIiDNpiaceKQr6oj4gB/V/dCKStD9Ou6jQB+
Vp9grGT1Li7JyKZPCyLBej8t+Kd+J35k2omC7gf3MAkiKTMGn4NkgbHEqwkLdLqr
SifMW/rBM5YaxiVs00m/P67jfHR9XoAvRbYenJ6qjLFW7fqOk2Db70279miyTznf
516R6kVhzEKAnXyNBuvOC0i+FF6LxsxLEqGvsL1Qqp278fN6G6Lu6hndWCZLk3Qr
RJEVi1EwhN7J9cQbiMOgXKxIxHqEQE4blVFrOuOESpG13ixlkj+uJQuxv/eO8EFo
45MomceUS1WDwOCjv5swneHDF6/nPYbhwNgVvBZNC0EvM3Tv/l9pxrQ6hFqeOxr8
k7HQS8InUvtwfXWg5a1KrEViH4NtENlExlDZ0VBRPjGV4Jo8YbORVDOYQKBra6KS
vByvDCzlsSEF8i6htYD7ZIezI+6u8w+6ySfsDSESwPIQe+dmpX5hMdfBvhZ6Jbg3
VUs9p7dnpTVS7Vat2xW1LJZwf/XQR/6bW62lQ78t5ngPYOBSX4ATrHujXwlxcxVE
WB6lawZkzFlrqUbkOZPFcIgEQBzWtDN+tWPCcj+EAGVbtcCuj1iXPm1v1is0F/w7
c/iba2S1uxvKFXT0kKrA7CJmyvcrtYLAwh4UZCSxwOFZFThNK1NK/vQFtqNLmqCy
F6q72ibDKoX9ZFVu2iKEkvaB5lrNmnO+iKt206V97xGe91l0NmmnuigRAjKeishW
8ul5GYO/uBTRjhEclfrc5GLxGVm0GawJZpUlgJ+LprZaJiN3OOBV6CcsEfqZN2Xa
LOhaap5EjiFnVugNDOL0Fdx9G79IE36sLa8X+/RPwLsFPAcphHDG4Ks+jt1/JL8s
ktV2aeLAWAso/VT+EluM+0Uq9mu3ynNs7nKbyslIdj12py8GGTgehFiQOXb5JnWT
PG/77tlmkoeNJlo57Xq5NlR/dHm9H1lzcgxmWRVKbmr3STWkoHN/WEYzHdNEF3+P
MOfCzGo80wn8DUQUiM6IgHyGrx75+0iXw1se+58s2vl9b8QlZ2RbJDPtEnKRH3Er
7cBR0TFt+SL2WqItvCOd3cPl/76nRchvr3U3rE+9RksYnXueAmGxCWeRg+Qq1pbC
4IEO+Oh3ufcJUl7LrfQ0P8IN/ARvWWKSRzaUu68s/e2w3pv+VmzBUhoUn/2I5vvy
vIlbOxPQF/wDJC52lkaPNnlecsuxD4hsyRngBKx68cQrzo4dKHE6myIbpZ2v+Zbj
bdznslAUfp+X3DYRxgbcb3wyxf7U4+03TPHhVU9tmnTUxUJUuLuwYeeJSJTBM3LR
hAcXjmRBSEtFwWJO3ATDSubMu/4t9cGVSScdndHJUA+8YA3mObbd1uFQNPArC1nt
ubNPW8Ija96z5cUTCfoffxD02NxiP2K+84XyMN0D0sWD4xYfCiA/c+jhRWjGLTZk
CX78KB9qRHZ+mgoDXwRliasyQJyyOk6zDo0NL5VLnZr+7IvwfHGw6Oz1FJ5o11MY
3xzEhhwCIb9L48JEZdzfAakP+1b90MoOop2RkFIe8+HgXFUBZ9t7righlJVWG0Vv
Xo21VSWzLRQ3FmVDXlZkPwRvdB3aNM4uGIRvtdZ8BoxiysogdqKd+BhsPsdgTYs7
wgdCC43kaQDoksW4VAa35bY2lZnZaQuP2Os1fTyXjKKtYFPBzka1mZfSUiuuFij6
gQdfRFSY1a6YmcdAMfV/0Z/D4uZnmLWORWumCYLBoxhHYhv2HhWq8tmmBoTnPKAi
V06SXB214CR0emIkaJVvcjIptVbSY0WM45ngY+ccHKELbmOZ9X4If+HwOoxfiy5b
Z+Blbb7BJhOsvDKd1OxG/iQJWU6XhBmn27U99Vx2wxDs0EpvBhDmWaXn1YI65z7x
dfeacwzm5tm3xuREC1srzsehiYsRJ8dDoCFlSUClXo5DnqAboF/wqe7Y9zwso04j
TiSatWeFwEsXmH+FpvrdVRxPyMgziW/3oCj87RN07zuPgZD07NU9Jvzu+VlBd5Qf
1aFm+JlbEkjO9d16rdRagKo0bXSv+dFrTdJ3YlZFq9nkgBKPeRRqU8OJTEme8NDh
aXpiYM48Y0SvFh2LiwAwOF2DqIa1qD67LAyC3CO08oMOsd0w15iMGL85QC1Qd8wI
wO8VdQT6pMC2oTRCvU/0I+LeSoJZwbsfEzRCWhXOZw/QXtS/jfPwScaJisDSMpiy
Js8mRrCl6MkExQYuOdSh68lnmahw7HKekqTZNIufvHvrhDxAYXS4BA8/hNpaYbfe
yDS8GJUquFZ3KwGglOBNRDxAJd38w6w2RGNVzu4A7hlyOE6NIc3BlVV5cz36ApLh
rNRySCccUXsSwPNBoQ0SumA9wdbuPVX0hB4EpIkzoIk1nZ5tcJp1icqtnr+ovWs3
LNx8tesQOWz+Sy9LHGYcuBHYHR05YPUTOzRMKkpiXWF4jMlJovqDzm0jtssj0MY1
9g8oAwpH0hJR+nZAx5ROpjte1TFgUW3dGjgfsmltikLmIbY2WNlvp7fbE3RATOi2
AeNifWbS3ZCoWAddwMDiQQ9UjkJEk4jVjvt6NAyd61YNXMpqOwcBkb/9k17hFVnG
20QqldR8NVIsHhpOyS2ZStQ/8/M/CwHWDXNNi3LFUdw235CYTnMZ14Xp+QWJTIhu
7ekTn6fJ/jJ9hOAI5t94iCOXLoPxj1ebloAS/BYoszQziLvg0JtUvI3lV1NVgBR2
fmvNhAcWhax7gHQX6R/IpKBbzmx6ZiwJH21k/YC5rHAWaR4MtF0Rd1zLb1W5uRAZ
zmqmgc1awoZ50QYdneQ58eaBj4i+n41usO1MXAcvKkK9OACtaYayTt4xCfrp5q7l

`pragma protect end_protected
