// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
zLugsZFmUQ376DHN24FvH6rieDyoUDWEVnxl2zrTRcXzpe9SKi5q0M1L0KIy
FAgiBrZPiAf5YIXl1l3+zrqmc6zza8u4zl18LfY+ZU01FwdtB2eVITVOVJKS
6+tgE6tsaPkHvyTRFSKBX3+QI39tC7nG/3j71YSg0qey/QVGp1ijTPKXfAh9
p0pXdCSjpJSgBWpJU2gPw8me6FJvOz+NqOHkSOUfp9CnbCrcxNFCRvyjZVtZ
jO06YnLsRtQxWxJpXTbgrAxVyZyooZN3wZuOyN8KsVrcYjQDHYXmkv8lRbmT
2/2Vhf5WfJ/tvFl92BWYe7S4EuXAbIYz91UJ71JYRg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
gzChw5yyRfgEXTxAeb4epkHEI7n2jFr6FQA9ZG9QPqD7GqDWCByGvWQ9sxfr
AUg9BeIKU4kfUnutMmRWzLGNFcA+xdGO4xSTWFTvhV5ZiyO/iyxVmozzcNUv
7X5vZ4mw3ccJiq44x2SLwC1tzOr8Y+x9FZGhzI2pAXj+FOrslTBrt7u5KQyo
18Q0e1XhcVTWzAxqDQL7kQH6xr+a/z+gAHXiPJPpRAiJd86txZJpefI2/+v7
POs2VowapcvVspUbj4170IvrZna4klpUEKTHnpflEqDF05NIunTLsZlvUFIb
h0n0bHSNEuO1TRczXMme6BsANN3xMj6jJJ5A2KdVmg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
RcK8uDxc7KdFQIT7sjJ3zGeNY+FUnL8ZFm+pHQPoeSyj668JY/+gvwhQ/Ffe
PG1xAhwYUVFKQW3RkucnngSq04EsHkeMvDy18BVXAnwTj+TB1doZviQ7p4PF
RGw/OnA3M3QQRafwvgtWmpfc90BuAMUwB13eGdQQ69Q4KrA4thWOYVd5l1Vn
MvR/Azcaa2/dfzlbw2zzaFQupzXujqKv4+fih8wpr//vGEEpbzvQfD+mvAo1
W/ox/UHQmjH4fTRo99uJDg6Koy+o8CJmpdQAyjDvab/80VI88WR+kg1EHehu
2OkJAw5XGvaeuFrO22CE6V3r3JH06fpUCfDm91VvVA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
OvkwHWCxe6ZWCJ0AgkY5t3mO2DXDeL1c9SE9vqgB3w7NthtGt97kKKDjoRF1
zTleCNpsUGoJtWOM2A1QoFRYCbSP0CIjX1ySDLGM+Azx78Q776K0EtKnm4Pg
wukoNj90LEH7ZKHtNn7r6e7TIA0zI2pVFEshRafe6h1x37rAyJw=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
ZUsBt0gciFZLbmaUeuJhqyWBTAr+5aXnKaENZYz67Gp3MNTdJ7HhApYFLI6P
7Lwo+uJG0ZlFXc4yhddboM0pLzASUa6AgdJVvYSHR7pCy2G+Iu8zmTaD2qPr
1YXl/stfZ5c7TMn25brIMn018Z5HFjWSvtr4dHbgQctQ17ifa70yHgU+FaNm
mXa0bDT9Rq/P2DijipGX7AMhR/d53XpnF+O9r1n/xtIcQDZJLPoV4LylTQH/
sGN0n0+tICMzI0cGi3UXi8b0AnGQSVQcOPGdtiXAgjZCUElJuRjUecskdFIN
jYQD6Jqu+gjvhTNt5NvhhxKkSK4DwOwAyT4dhxaVjZHYcWHbUEwGhUpKMDBD
q4D9/UZnXAJmJZvgaRiVPVX9gC4z+XKghYEHvMohwyl+qrcgTv8WSOGcPt2E
LdBZFw5ABvBxZQPbmBs+uLG3FmaNWI4Sl0dZyrMQVRG8yq/2P+DKwq7g2oDF
OM3TxQrEcvBqiaEUxALQklslT8WC7Su9


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
rIyj/3GuO+Znj2zoFUHVc3D9ANF/5iuju8zgagH7MTn4gLzMUNgj6hKDsxiB
XZvKzEmSEmBDMQY5y7aN2QXigzBcucCZWhdEg0DezV501hBjE9VoTg5lwj55
hEmSDuPcLSCCdlqzCNhPOxdj0vb6Zx8+Yhwn9mUm9S5uc9MYVQ4=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
eUmBkHBWVlCBnVKZwETbDC5fKtNjzTnds5157jt3AH9WqphNzv7P5jEGkkNv
2zihttAdQ5CiCU30MWsjIURXBW8HIqcABJMnXsowfATvgwkbyu6uwziRPU1D
EVd1bqHXpS9L/FZeHkTVWu5OiPARHd4M7+/BdvlXxkMMPMACHmA=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 76368)
`pragma protect data_block
Eadi/ubP+j1uc2z7CUQSfZWt5WiFHCjZ3u182PlaVguVjXMBDxGBHTbhFj93
s6ZItvoCHqUWoPUN2vC9IbKVvNW6jV6FEC7J+k0Ek400TXWhItQktGwiZLKa
/JFRb2cqcKJODzZN94ozR7yS/6bb/YX5X+wB7LpJ7lNTj+aU6fjBGvw4PDFL
U8Wc34yPoGtxL3HJvK+u2orNE2gazOSvnBUjQ+4J2WjgaL1/eK2Zr/zCrsBQ
zsX2CJHlLT8si1PKERwenwZUfZti+gdoHSFGFLPtXtSMouPWHn1D2XUaQ15K
5SKMADlJJcl4TObbVsFTuutPJKMPj4cZ9bf8SSIwGDnaC2gyVkq6GJyRIIwW
w5X/th+HFG0zgfSw7Ce1D3HU/1XofE3ugqm6Fy1bn+c49zRrY1F5BG70Efel
M1ALaEXdeDYaUGFmb64OlCIF2DFUFArCSVwab1Er1erj2n4bn5IEI+oYKWiD
+cttCI9xHvFZqOAaZEo9jUul43rtdHokhNGjbAS/VkaK9QgzAgJG4I5At0Kn
E5SNsZltnjoD8/MEmHShzt1bOdmVK7pJYBtw1zjNBGwlxs1kWDVWoU/P9FbJ
bY5LXXo1UUsC2F/BmniOByowP/TUmgkvnW+dX+1j/60/LJ6/wOPrZmh9cdaz
P3svDKg1PQgq230oB2/7gL8DGSrvX8JT6+VlsScqDs3Yr97BDrebmlgE9Npf
lD9lBaBFyCVwUVBE9sJW6X11WsCCQ1XmbeSjonNZ3opvbBGI4x8JaUTSPkM9
qf9z6wG0K1yVNTmW9XEFxhVeT5JhXPL4yir+nZSCWq0tK0bQCMcEEUK/jZ10
A7Rh33NTksstuvlWOk12QXh25J5o8bbcOQonMwlIdTXcGYaJeUv3LF6PrwJa
30NtczFM7XF2H7YvlXEbTg9VzqUaurd8YkTXK/5UMrQolJg7Fkd8ranzJAjP
LoeXVv3+w6ukk75QfCM5YwkfgJxTOTn2d7EETq6/VrjnZYulHBQav/0tZrrL
V0ov61Xb8mnDi4R8R/0AB0ueXiwcjL+G6rg7KlZ39deyYeOP8j5U/swh3Au/
nMP+RTgVDS9TUdKdM8VkvOIS3ilbjZiKPfQe2roruiyy3eoM3oLR4eKfQ+Gn
uIshhyThS0YeWtR1Ew1IpkfVp0mqqsuZ3G0Tog59/clE4m4EKhHKes/QcVKL
dbaAIMlIEL+3D3yuxrYlvOVMwlIVmarIgfZtXD21rtK1XKo+muVULqSvD1qH
sP+9rqCvn1CVmq8a+XLElPEgM6Nwj8enP/NeU86je4tKDW2HC3pcNEIHKg54
mFdNFfMqa8GnMqSEkSUm4cQ6vYMpSJRHGGassvzxUAVSRdXQyskV2sk6ZXSs
a4Trr0CzYxilenseIVv+krTrVDaCX1Qw7YSXiJiyKu44QyjZVVqMOj9C1aUr
gCiVeNzuwzwzWBZKueuWAXJ0A3tTA9p1jlThh98XziBEQL4AlRO0AImt0tpj
Qdbc5BqWpdA6mn44btK5q718DIrk0i2rWqluaRyFhTCDwCHpi8unA7Pb1Cbv
WuytIzan+/Jr02NG5lfatfGxCcNLx8ZkhcbJ4KrFEb1JuopZ4rUoCTacfzOd
lj/OVTPnWCPLD3HwPX6VSKihYgk92xT76wFbOU+f4YUSmDas7fqwk95gTq9p
ghDxU0igcytWNklfl7ZcsOJ/pVbkmzYaCeBM1zIgHTJcrzLGkhEcvrKYJRbU
6ZaRH9A7flSzSK0spX28x+QWdWA95LH5iie+97B0GFtHiF9W4/bnmakiJjOf
CKVMu7p2pF2MrUEfIO4JvVgoV64HRaH+eysmP3FVs92kJEwn+BbUgjhmJ3oY
YfDqskQw8iqiaYELN27ZI/1jW/tZ28Sd5+i6GoB4Yu1N5gdZMNgi80ac/Dts
Hnz3s8rlLWzD/dII18RbFDTSMIH6CQcEvIublW8OVHuEH1QGd+BFgTUF8mwl
DVrzoSIJnaej5GXVSPcsW2FGlt8UJ7hZCultcbnblK961lspMWNC/u6jxxl3
2rKpnA+BUIkewxRU5SSHueYcGkd0nX7/XFRxZB0+hmJ360V5D9pO58uZ8Izv
DxoaQUf5Y8Dn4Y883so9XLet7zEVWrYyPEN2xpOj1w5KyaM4Gvarw+peDttK
ysLnrmM8WdndoyFD+OowDXvdoV7jQWqLsdMCbXyxgtKoqEEF0RS2iXJYunjg
ZgW0UJ7Zm31s0fCwn2ok/SRCZnRkMxffSUpZJwN9C7sMavFQBra/dcZfJcUp
Y5oCY7CMPgl5oowZnhVZXPNQP7PkyYdutYClSaAMeF5jvwNVfT3kHV6sS2+n
LtOXTucJAONeXVmsxZH/Z7WUoCLFE0yYE4KOkxV1KHQw13WDfmfVtnaFC++D
AAEt/eqwHjhF4gCiKoM1XhR72x1x+OekZsxSg12jg+TTYRcTo3o3s8VTvRF3
sfgAc3n9X5ATzrnOGmexLqNW5cqffvNIF+Gjb77PJWCPBth+7c26ioDjAL3M
Yz+/YevVw6/7JF3knChVDmqv5kKcR/Q6IqOmrpM+qEGJYdY1M5y3najbznho
1dV9Gghqv7GV9N8+164005IKSj/AIB9Mn2jleq3qqoo3A1GCPpcNQHl7YRUj
DnA/xouAiehS8o6kgkWRcAvLqZ1cjrYew6t2MqFEcuW9m7POdlDSWOJ3hr/H
Dvf2fiP07ikGmjN4D6ImWH6aYT1WFg35+eJt5Gg+JFR2RVjC5PgehCFSWtVG
CymX3sIEvoKmcMSgIr5vOHSbctiRY1fNjoXhtxqmSCn3RcRe80sxyNLRN2F9
pXQS0vQxCMaToE9P+rTn8mYeoU2zB+CEpl1enZxtyU6PcBFZg1mxgqlzGLqQ
yJTK9H1xSAKYdwLUcIMj17lPmiq20qt3w1+/+PRw4rOPN66c1OOfnRphV7e3
05hy86JU940+4MCByqyPkw/Vo+Idky8T4rvILzlsbXNN2kGORMBDet8iNCjr
+l/FQLC7kjpXIN37mAI2Q19w/nDHUHAV3Ld3H98zgKr3rgkC5yDCUMCoho2R
hJrE7sWCjln+c6UnsdAWfoKmHYdfLBbUPj8paoSkdOMjPr2p3eLgSOAoq42f
SFhr5oohgl2+lEbp5D1USx6wmWHTzvND1iD7wxgWbvdFdm1p78mCFDfP8/Aa
tnUg6H0N36dDWSLb25h97lUQ7xKRqkslqpXOyD/MMnJyVuyeC87qqfXWb+Ci
VVM7KJNRunnShuRY2o9eqsSDCsxspW1DjtmQG8KxM4F5GYc7olwlAYomEjhW
CSkew2IVnQQeyA9jAMEIsLpQqGF7rHHNVwv5O0MzhOYK9bEqIBm1jRFICxlL
H7sk9EucoGAd8YVbH2noiwP9ln83fqJ7gUZMdH7v0KH/ne2f3SbJqaw3oFnT
ZOyv3Vn5vfeUGw2zqOIVLJEvOa9sVYiDVfg3BnFzRM7LMu4niM4QBdQOOnjS
ZuwLYpXgdL3lvKBlmNdp/9sVveK0AU1pMxHCokkPvd9yzmQi4rfFdrXUduh0
CL9ABUKrb4Gv2CaTWT6sdNtreyJlUQ3TayQbVx6Esy2/mQiRq/Gyia1kYvAq
+D/kkpBUYJ7ulY1fD9FUozd38FnnrzjsmYghqScs5i9IrzgMHPLQkknN5RpK
TGv6TPaZSudqGkOLVfZIglrf6DNyJZ3F80sHDVIkR7Tia5uX13mptC5ppZCo
50vQsXYQXTV2um4a+5zTEOktcerwWEzShtaizhUssL+9ArVR88RTVY8hg31M
zMtyQxIG4E+x8net2D8bZe2R7rV8+06nVqVZgkIXEWFC0nK3eP++3XUWsTZr
0U8ybAlChHHFAdzdcqA6AKB0Cncv1h+06V97tbkRcr8dAAx5cxscXFZdvGIm
9hYd6M9RJbTFFE8hsRxybgivUZYH9bWfJuFD1Tpdqgpe6eGjyb421gsm8qQ4
Ux6xSRGYHKbqiVWovLDuNlji7gbEgxYvli6aT+GtmCuMzPum560VDVCJszDt
6O92k4bwKGlh1FLpr42oJuAONJBd7zM4Rx3rV1wHwNHE/Yeu996yp8S6Zg69
yKzvJVeHu0Vwe2gGKYUuboT6lQ6lIBR65HEObVomhWR9yMCS5HJX8VfbkiP+
FZlNAHPosb8Uuz6+0EHu7npm5f6ltlC7gfAcPeC0SmzMk3ECIwUE8K1o8d/M
QpKV4SPd1dLGYhaZU6eA5cYBgvs6m6KzgmPU8qV5/b2nEtfK4wlW+KjKmIBv
j3XyvhFZ46DrDGD6DhkAzxQWc4y4kAjF1uH5F9kUHHzF+NwbkSDBvuL0YgQ1
4t9mhqQcz0QOqSICjagIp7k/Bk+y5R+sd+lkKpBqUOuwxPChAXhcTvhexasm
o1sx7J0AUsLY1PGkfrXDO81rrgoH7/nJiq8PvNT7yGG9X8yTAeShwv9j4SkR
dKh90upm0VBU7z965mdFfSEpr5wxEJLH0kySoUx3iGas8gFDro3gzCRLZJmU
IGsm3wK4OkcwxrAnqotW4KsT9mpZvPrUVTvV75q/7nV8l8aLcDexa+9bJkHG
zgF0uOZ2zZVquh4QPJY11PW+9+WGnWDTTu1IGDiylEz7ru2Cab1WDjTMXogo
FowPCUvCC3M5RQO+MTcXtD0iBUuxLOR9DZ0rVLhP6XkgiVPjW4FZNGslgtnP
jOHyyw5lOKN35FDLANTRU2mTN9nIzMkPR6gJ38Dt4uL5veRv6xYJDC91HkpQ
KmHXdYKB7VkrbX4VBYnBt4KlWWybhdtGwXeTi0hX3gizzHxzsawHNny1sDsI
qJKhDFpjy/wEeSPKiFU6VqlY6GDsR+AGBpdmD8tch5oM4vEgEXSIbgcoQZMs
RdNVQB1ch54gWhDj4NYam/Mq5oMTAix1lINMhxoOTDCm1fEdTWzLMWZfeAsk
CEEpKm6vIwjpfug/OCXf0kBtIjAc+8bKr02hoLeRhYddSxR0PtMboUMEIIbz
r0eK0UdNBtWimmKVRzy7fKSIxdfT2i8cTDP07kdwnpKG+soW2OaMXwbBuoQ7
7WZ/KsdTWtB3tOe/6oYqYTwX/z+vASvqg/dmhTZUgoWfrxkvF2rEOU9DQVA1
TOFJfCoFoxFmoPPpfB77KYq96vum88P2XrRv4FmnufDoAwre6IzUWUi8t03x
sPaW0m7kcsGOlETXTc14RwDIT/Mtn17BSqtpx1UB1ZoMr+yb5Id5sx7VQcsU
qTmdWrnpJQ027PZtXNip8gXXxQB1ZQuqyvgfdZVdQhlPq10Mde23OppvL++p
N6ZbyBCfdMM8CHDCpySkITCQuP518JbqVKv5AZkuSh/JWW5JrZd4Cre9J+hr
zD6HZd07cHg6e9exygEID33B26PNQl+2PyZgUZEWxkliGyHeAPnU1ahKMdA+
ZzrA4iEAfRCAh80KbTvLU9Chfn2mS0zRbZrP628oP5JIRue7NS8hAUAyKh6v
pRZRDT0QLEgzX+Cd2cNdpUnJSgGplNZ+8/KEkymQ3vhYy1/f/RFHDdZysYyk
399Ojr3YdDKoTYYsRTLx8kafH09+yZiXhDrz1+/pPJ0FzNfutaJE/lwHf4kj
q7A/hs3Fnut5KhDMDPCX7ZMy3iIPEUhO8Qa3aURxg3NjoM2VEbP2wV3UGapr
arAP81tZ2NcrY/JY8TxiUiPOR/u9xH+j4NyEpf8+zE5db3CAIpd3+ciaLE2z
5L0OO2/Al32eZ7AZvjiVM9rEq4SueH2UKrtpez2sJmya8w1FsQ4w6leOst5K
+Nvz2PRX6v8I3g4sWm8aEaEoWBusK4bf298+lbKa/U2HlomuyB3oMjKLmw2+
l7JXmTYSx3cHjzcOz5TY7xRKwvoa1r1sEGHbHXatCUCjc0sqNQWqxxujqcS8
BDvfdqzT9ksEg9hox4wxvycaN+fyVFRn2gAnYGdNXccDxK94XTMqmVgLfCJf
lQ4Cejm16yTa4GcGqPoyWzA1hXYAK2gVWqtQIoVWJ+xw/whCs0o4cAQw46gD
NBgOuZEau67D4si6lWRrPvJPhVEVrL0T6M4vMLR/XnIXXVqezC1CheLpaluE
N6xI7O4NFcDZpw2I13XEri0py2ZVmiZjoygHsbtJw1xfsRA2nThdPGKZ4AJe
2Wr6OmFA4+cVLlwJlno6DujV//3HpnzjOJgDVe18UcvAD+c1CllZaUUelBvO
psZAGIC+eYKnIfy07p+cV1p2Z3vZ9D9kG+r0q7bCakxNk8eQIJHZHM9qAED/
v2ShG5KQ6K7I7TzdbVN9BrA8QodiI5jBgOZAwYeP6KY7/zs7yfWMd9XDKOcv
UG/1rAUiQoam1PyhfmOroHtLOPN29iieQPHpiM8vUIC79XTvUWYTAVEftsZh
qZUAKiBjrvTLLX6kkN5C8Law2DoPT1YoQxNOEn5U8jmPxfV26Fy/HqhmAfjm
/m5anabwAjQnssuqZdDOrbjwOalCPDDwxTq8X8zQfFwLLtS6b5V+r/Sny+uJ
RbYuwO1JXwBIJ5g/E2znCshl5zXxZLyROM9z1H2WiEtbPxjLkF6Cofn/K6mA
QzuVvdupTyW59VIWtejbFVVpwmZ0t7Uj3CVbpkzSg5o+jZ29enbv5yF6pj1k
h9TZlmELcxlNqQBHWyvDbX6x4HwPCT26G/4SwejWqJLHORr5YwJMXriOEvhE
ROsfzRZNzLdx/aR0oYQF9A4gV8OQa8nAhSr5Myb9ycbN3uzPTQyOrN2D8dg8
WjqD+ea6EE3gYuUfBQdda9weuPw3QEBJumgxRNW8deseovMwfoNvLqysJCAJ
E2yk6isq8ubcb6EdHRni9SvM2fxwH9h9XtzxtNq5urCTelHuQ6a6qVV2JoRb
9AdFyoT6ap1pPTR/PYHgwf3xSpzsGxclwoxlKe0TqbMScHRgBHM0omaGnqER
v4ghntmKj9Y6JWBJKfQdf1yVpcilVkeFl16Tn1aqTrpS8YGAqLE/2jgYxBDW
FR5ie4aph3ye2HIAxhky7DMp/oIaCY8IxCVnxBzjy7/CxB974sCrrNyo1Zmd
+PRH9PyGTz7VgmnnLhfU0nwe/oz2Lw2SpVWNqYifKR7ARdG1bTDHYLSxz/wT
N6ROguyjCqkXxK5cZCinnVKxwyivAt0yC0IX5UC7zj4EUDfnpcFQy5ekOVcp
vJCvC+X1OLBunOu8axhj86k4kHuvnEZMsgJGznqtsfQzxVYqVakvkjDZAXr9
/WWgHsXZhX1ZAttoV67y5QdY9LQwmZesAQ+KS4JKoIOECFWJ01TUZ57dx6Di
HTmPdsc/klV+ln8aSlcfDLyy43MKaklJeZNilhEoxMvSC4CxB5/BD6ywVQbV
YzSA0Ncd8OvdhYvcmeXsy3fwo+vlepkDBDXAKfT4aG1Val8Xr77bJ37o87P3
mlRmN5IAPedRwb/7fXv3hhvKDIYn++NnKOmRq5HXBJ1U2llUi76/yaUIL3+J
rVB8l15Gms6c62BbYl/FylHEw5QcRBUwcv4OZOij0foQvTXsUye7oeOeI4KU
Za7aXbkjUgtMVuqf6Kk07Tv0Wd1bxil5rt2BobVHyJ3hahTbxFhYsnghXhuV
sEVzz/noTs83a3NB3S5tGdah7JS1nvvR+G1MhO9mAkk3ID1TbqBxOCyMA2MH
+zfsSbqtVOw2RfbGUlnU1jmRwEWPdJSX4fvnvAeatz4rjvSHUDiEGOPDUtSj
jepaNkMNJQ3TBIStAH2Vht43jWgufQK1EsbQiK/2axI60dG0Z6Je5962VT8n
87Tp8hrHUt07aXx0ZZHsdFeVMr0cLNqzpdKrC03dCoY6dlJch57+tD3e1vrn
tAoD3efDY7cBO0WFDafVc1XgLzZgygRJt2Xkv3TzT1H1f+1HK+DzU7DISyiH
+fa3o+uZaV5bsLiVnP8wOE4CPfRHDvAsABtRKlMVqBR2ngwJ/Aq8K67d7RVu
Rr1iFT9DV6GtGLOIInCa3DDNN5JaIPDN2W0gHg6PAv4CKO47S5DCm140HITW
lodJEDPrCHqkU1IrfjhyHbRUjgRVoSbrEZWj8NtpgF6byZJHRQ6EFzKBWzNt
f3hGAK12jxi7vfhgsQNS0bX2QA9I9YcgsR6TA7N2gqgCim/PS2FoijhJqjYI
lespRR8aXIBPbhZTw7PKytTNnDdiArHKKS+6Tx8/kPgHgXFHxoVNxD3oiOuz
aUZ1DOh592ODEtAIqbDeH3Tkq6ND112LFkVE0hTgr8459AL/ObFV6LisbAD/
sCH6vLiVUf8PcNAF6ZZHMiz7WqT8HsxR6uHITNZTrkym3nZFr28kBAvg4LUU
QWF62KwHAwOP0am9DpMrxgdCSgZYfMxGb5jVipPMcYLVVce0OY0FwSqrkdt4
919RCxVm2LaUUzmd3O8kfR6mKv3P49fGeyhEySoAWtuthmAIX1SqZe6seSL7
n/EXetix+Qt7wMC7omrnuwzgOw2xqaFVIZZBwWk+CNUSmuGUqeOrvT9vYdd6
SMF2aJpVC2I9HeA5Ou9uetyzK88Wsi4ANZwceXEMlmEu0qM/PlBYuxPlXBqS
UKOuRwwvdkRHnElaTiHxtlWPmpiNQWkME11RVRTbSUe7TgIvyLzYY0Z7h/Jg
1ylMLWa5lk5C+/HxADkFqHmrN+cScLECtlMlxbFV/rVSXH6Z97nL3ioLvyoW
jw/PP85XJGPWbMOwoUBgIa1+CYVBt/bvPlF9WO6Ayy7a30hEXSr2JyvSNv1q
I0gEnRBbLKwl90pdacy3aFXpRm92lA364cPoCNZXNPV2XcJ09uGj3HsA6YZe
bZq69g7QvatoUpFqj84jhgpVnvqTCq0uKzs6T0ROBfN8WtBgMTbP9Jssq5I6
Y7luPhOWNcJR1OASg1fKNWrggTKDbbU6klls+IuWP1l/weRbhijVINe/KRbL
9VwHyzJZ6UzcwmrKMTmkMStzfPLePVy9Tqmda+bOjZsMHMsuya0pMgeASFQR
CAGKfS3CWcF17t2edMPx9tjpGj9klChXskyWVVUWLl/Nrq682WFYO/1abn2j
N1M7YSa5B+TWdiK5u6YEND5FBpj3WdWo8qgBvqhOEioYgqJIptgVsKDVpAGo
4+LyyjjHSPveWWlo0yafkUPYrFmo1mZrFkvpnPJ9JYoXaxFue7ftw+MDJzig
W69+jzWgLeCwY3JcL9m3F9eJ603eq+nPKrjs5vgKUsYmN1jvXfzqweiC2v3I
FaYyK6aXD2wPD+vZD7vQLU47ib9JlFCCqtzEzkdhWwHh7bo+n0v0X3NEb1Al
ijhgb8yrj2Yn8H/41GoEzcxfCBxZycTeOqDYCQlNO0Tir0102U1LCG0/bb6T
9mQLyhgZFzemp8ixcfSvIQwA60YavDoGATchCO/A0/CQPMePQ06eNAIJPmtN
QHBNgt4h6xk8zCa4vDKYXQbg6RaA2g0Y225aCqB9GsSsDn5bHbU/SBu37pL1
BlqrVuh6ItYmUY3Ys5m6QJ83l2IkpuEftQWxxbkg1lqbd7V5jBXcn40JR8Ka
yjEZFHiAx2k716PosBa9zSvQWl9tw5ssvwZ+sxuufcutMu4lLwRuuMJSb+Ol
hKtdibcrVChNRLJv6NBlHYRxbh553ft67yJY7CLRyqNh8IQjYO23ALkjys74
b35ynlS1uLevNf5B8U6ZuhM8IYdbG5/Vqv/zdbxZiBFZ3lpcZsXNmzJX9yb8
yuFVhdtgBXTkgO0Rh7mFzZzZjZAzdQyhsXKkfj9rWfRZAF3jPXokqybfZW7G
BkWOA1OqZkypeG6Mhe7pvXf1R/RphWzMdzDIf8rqEHCGixFpnUv+X6iL7okT
+xJlI8+usZmdfAMUX5ev5+ZKkdVK5aezhOzMEjlR6ZGyzVpOUxvKh/u2iex8
1AEmUJC5mmpibKlb+tTC2igUx3H3HQ50jOAzBDHYIBN+Jbc6w/QI7+BINh9g
M/jZxWmvZi5OU5VqIqRop75nsIW0Dyb5H/KSwuZbrwCHPlTyDMA0DQZ10Xhb
FAo5/JfhHKfmJJ9N23GJPeP6HmGViNBENObpJgLBjuqHQLsOCvNoBUMMgSAH
1w5kIOMccxI2DPQVfcJRZqb0om3ZRBcoj7ietLethFB1hc8xzV6s2+ygN2sc
/rtt3c55Qu8KiClxG8Dul1lC7htXDqFvB69XOhEPiGV+JAKJRv9RgE5uxVzX
Mdjsz/9j+anwEEtooPx+/bVgjg1qFTZ/qL7yqdGGS9eGem0QfRqTzHyNbTJK
FcKCVKGVEHWmqp4YL/MU916lfZjw7lZpBfNt3pi8NrYTUzaGafQVMFTgcgi2
1h6fJr6j2UVjFOaZIdMDOh4ExHB9yfKT06u1PMSv69enEcennOcOhsYSf1HL
1kSpnfKIgHPxXeeiU1WNQB6AtWAXNsjFr+lOFfnwnfyzg9oMAhKLJiMegttT
vOskPIuDo+dk8/bA65Ro/MXEYUn7lTCKvmghKwiH8chNSbnA5I23sd7e18XP
so9jvIpfJLtNY+JkYzIlC8+N1DFEGNOGPE2eoXmr0Xw89+Ps2moFVjhI4seJ
sbYNBghFqgjZbplwWHw4psZL+5QfB2kZECBFTagwALk7Es4qYYHIelLBUzyG
dKs/umYaE4amDwaL4Pg2vRREJYA79zed8bJCAtOuE99lX1KcXZM9u3n8flgm
pNTCK7p8PljSVHcJPtSALALFuu0qW9wvm9wchzUWbuN0d10Prl7oaMZ0QyyG
kcIePouAAERMde4l2GkkcDTEr9/4rXW312A8eg9Uk/fjd/GTAv5CbHGUvs5x
5td32p2uNiEgPHGGOdKkuobF/1quBReVndfS/frTjAZ2VoV5C1R47i66pOw3
X3NfdcWGWD2ax1Dwkgm5eTYhq9wSNPQtyukejQCq1gS0Up5oX7gnMM1hssRd
xTwht3jPnPTU9ePdUTXYaH3DNPa9UER0mZf0siivcrtZQ63gOuq4Ejv19bwh
b1+bUiLZylGpWEf7sVyn49cljC7FWvsdzdkeFvCZBfS4+sKPd7MQQwXr75Sw
c/edaJdvjCvwA8hEy0ROQFl3dlzFzrwYcWhrlse2zd1UXa/LXvH/RFnbCrYg
MEv0qEl+xfr/OAj0bmV240Dj9+az2ZaMnEA7kW9YvxGqpPpRkJbaR9vdfRyg
x9ZeTnGdAe1UunMRdo0cHixpA57cFWL7ARYqHGxNKhADXacx7QSd0Ra/j5su
4e60nT0BEm64QGtKLCsm6ec+c95Lfq6I0d9NJLl9k9MQo5R/QXg6K+tS3yv9
xWrHaGq1ZZM6nmJio+Vk6a6nIxfqwqctDPao4JmxtgNatCa7n9vj6nsP/IGL
lbZDSxXnCYp6YrW9VnnAwTzGRfY7ZqN5Dp/AJSFyOaH2H93CvbiRbx26xdWO
/IeovTxSba8tK+FgsSdGmdf2TBzhyb91TYK7jcCrUuNJpP175xEWUSn+vcN4
YMOZJ/JCQAvHjyMJFH5tgQHnLAs1MtwYaLe8vR0D1GAFy5P93KzTHG4GfCTC
JnNLHfCO3RepUbyDzntaMrX5bVHxlBhVbWprTqg9yI+GLN7rHPZQyrhVRn3H
NEfcXQnpCCd02OjKPzLjhou7tVY50jPCFlRKlvf2YoNWfsa4xNn0QxIaCpqQ
MuK+eex642T432CHZXbtCpnCSzFNJpb2JCxy1yZa+tMZ6c1oPD5NR1RtRdfB
BQiQ6tuG9hfA62rCSUJxAmI+7zfUNTyYIAhqKdvQsC1rnSBysa8nyLDEUFTS
3hpM7VF0aDkAkUbgm9VeP/+pcbwXRFyRGxkUa9DgzP+MMH+ZnGmtfDxaf0+y
Eia3lvtYKpX6noEPTTgUI4oC6H4kaNrMRoBrO8OnDdvBzeMSSdzh+h/zHkOS
/SoPXRBf2BGKE1tx9YBl+R+qyYpggs2rtRFRDzRZ1it4zFlrd27YCRZ9twJb
dqv7NW+IWybENz9Kop5D2t5mxoty20z3T/T4ZYAlNoTOqiwl7YHC0/vb/zop
pLUQrJsGSkT4DsUAaOOheO9mUvHClIfETa76WErowWKEnmYHd1ASogEZbTsE
ZQ7ISaDkMiw+/miT60Z1P0bweaXv3wU3LAJWpAcPb1iPR35PJsneLRDfiIX+
nTP3z6M1gFPNhm/zuv9VFYFlPdq0/5BWXCCA9+3+BUl0vul+mwzISgEb/Feu
fMEAAQRKGR7Q57gYcyiAt+/9K6qkqlVQ3l0IMVFKuPguXbh0iM08VxAwlAxq
FW3l2zHqcZC7Enj+J6t5UdGeZEn+G2YOHfw2iXkaQ4DGT5MdfCZVARC/9rkG
PfsCw5LALfCExtIpoUDfcuevd5BcsePA4A4WFHSDLNkR9j6VL1gLZ/S6txtx
p02NGG/tyu8vDP1WDFB1geQtAksJvlXwCuqyWt1/oy7+493LuvbeUuaCA6dG
RPhVIKRdADE5mD7/A62PbvEFe/XK+Nwq3/FXbyJ47Qj5uPYC9ZU3ymoqJwUh
oZlaxNOVyiyDWez70gsrVn1LTkpuKV5FZQ61l4MuPIHBi6M8a3q8GgqamfL9
e72l9op4oxxO4W5fm0mkC3LcHsALUy4Gs8knJ5pXJEmSwjMHL2IEtQHPqMcY
/eyfHvvMthBcwl05kyHt21dA2ocoCcIxOLz63oXOP3dAeR7IR3IAHKWHYJiR
b1ezGtomYmiLQTWWD+pNFJcyO92tm3eBMuW6UDe+95FhjLfaPt1dLUiHmquv
TULPkVD9qB9VrBFXd+oQFiCANJz9fHsYDY8X3WLKIWptR5mhGedF0g/0aRNJ
k/Fr0oMjAOS1TCYYq9tq35t+fK9zmQveLLJslIVSMQgvt8xqaXcKRBsP8Og+
S2Na51AsLWb1mwzIuHqwH0ONswRjvQeJ46ArMaTTWkdb/SLPn+slS+WNX6bu
MRDIBnLO8ws4Po6E6/tITTKhvJjVfktmLBPYE1MwzAj+jbikSLQuAVfpeyt4
iqXG6NLX4zyDkzIMNAZlQ0K8AjEdygjDeFct+r/SGIRAvA1BtFFKpsIWGIuM
0QfDdEx2Q+hkJMQOHL/PxtuSBQAWdsqc3sn3Jdqk4l5gKHhCbVqWdMQRXyZs
+Wqr0Oe67tVUDSI2q3AUMGwS4NoZ4dTI1TztvwnhOaVEM+5vh4znTrISPnQA
aRgbgAhDp8axcRx/eZumQYCqgRDXP7GMWRUlnJXy8Zi9F5luNraygfoE+6oy
Egjkt0MMfZSwK9s/0vgXAFbCtEwD07Qmra9NjEj8Uv8Z3IUwTZl+/Y1MHu4F
MsPiORhnn8wRriVTNryuQlQ1fWJbL5pcJQLsughDqUXFn/Zfvc6VwnBam2uu
tkj7QIKyc0zyGX81S5oRNtfx3eOUVF22er7ssrqE67ijp51cvx+fedTluMlS
QAiHON/PmeqyWggqUoxP+mXhYKIVrGWEOL5ZH4c2pC4/U/KJQRG2dpV5iQcQ
QkBhAvBio06X8CQeKwq9kznjuR/zNBwkdYBRSd1NpzK9fl4roxCeeTc5fXfV
AFhpqq5Jjb+zcvyQC2508z6e0tBpDvHzNtySe/CmoJwtgxc6s6945Wfq3f3N
5akc7M2GCEsBIOiKw8PAJ9x/lXi/3BVeMhU8C2TB2hWWIu/G4OCuSg1ObePY
bpLM3930neg0KkeAk6at+oB7igV/8Mb47uEX2ZUGfQ1bNJJ+/7uGvUqKKhdc
LXMFSBEEKF/mWRszRjTrj7bBLKohb9RkeHAI0yahUMiXxBceMIF1zw8e8viI
bt6K4uulbb4JIeXK4ndrT665JWhJOTxZphUW2PCqzqSqWd/eLSqFcBbmewXv
5rhWrVGlcPEwcowQ3sIqVz3vHSo1XbRoBSANBADJ+WWEjTZqK2fb8wv/wZ+u
Dy+yd36rupxdJq8oHBVBvlV0j5QOnp6vobMoZoTk7r127WN62cxNFshi1K3A
+jhv886kwESfYM54e9cTbVkYbhXJvLmjY+/gm9xC/DNgL1vwMzruVOdfrzI3
wnu2vAGIf5VooC/gniitwJ8KEO4cuQbV3BPNUwCxmpwJgoO/4iIwx9/mxWxG
xmJsF+l+nOFoaHotqTOC02HBEAsiEAAhw7ToKyAWTtDmfsTN4oJG2TX61kCC
0TX86Ob8JpmJaxWTBfmBta8oOGq7wGo9t3/d0IV7xKGuozHoDRJLKLFv9OIt
T1l+XxZqr90NBzBdtgFbAZ2IthY2CJSYPIFXxKpi3Y6Mk0p3V8svLzcmqPM/
ddp7d7sGCOiqwywAuWOJjIZecYHDMNfAxaXgAztE3hBpS13Pai6LK0ZbzH5C
TnvG6k5RdKOzKcTWZhepMZerm8rYxPlCJwZRIKVI2Bc57L8/DmIizyj/CyQk
+XZPt+OQV2g9EKVOdjXAF3m9uPtI5eD03OXHeSPirBStw4P5j/zfTerx5l72
qAPGshHZyEoifibrRt70PYUEczW+4e8+nrzapwYQ9wwoZUfTMLejWpLBYG60
PNzABHopzjNDsmG9PrLgTavps15lLE49CmXOfWxG4OnR12JYpyDDfyJxg2Gc
PlNduoWpwKGADWpESV8S29bBlVmVF9guG1lANBJha+zG3V5k5FYCvqROjblL
yytKWYxZyo2ok6GSnWzSVLn/PSHmvqkghtyqB4nFektHn1xRtmx5faHuNAj5
2eBMFxPVKZn9QMrPjKWPZvM+8oH1p9drUlOH4Cca1OCJGiCXPRkxo2XDTWIu
XV+BkhEdWkjY6MhIU9kn3kJ6Va+YINDm4KnAZLTq0CD2ePnHUap3YjZSuaGW
CfmrPWe62HVSC85RQTQZRqcNUnoDkBPd2OPTw0s2EHvTrSv9XhXfN3+6gV8O
QZ+WpGM3/2AGYE9WKw0MWFgTMGIDksdnBx/R19Q3KXTkLDIRe4ZWShkwXtBk
pp0kjML45aphPKMxkHJGeDDGw+USzdIztKyqALoEpVkD0Rpm+07i/tZ9+qxb
5NcrOtZ+7bZMys2UnFn8m5cfGAmN2m6q+bqpYEsvnqRx6qQCvY+3iSxdf6kc
J359zmNQIOZ41Ar6iRSOmpbaXR1Sluvsas69zqT6jeb9p6q5x355eGN5yJGS
oF6CJ4rMEPb0Bv7xq3vSrmZGMRQonW1EsyzngYg1RKwIS1QFTRExzKuId3wT
xY51LVmGYAscLnkr+DPquss4+aQhRZJLccwZGwgoo4kDO+YAXtYo5+E2mzQN
FlYX2rc5pU0jQZ9it2YiD89fH38qMPy0emglfUAnvXCu24lLfNooVMv1GiVy
Jx5FYz5jAsJ6HdIpo5oeJMujHpH27z08lnmuUjLBZ8DFAsjbSGqLeYdeUvnL
qGK26mSxjf05eybpFrmVx6dyAbu879cYo9GpY+4Z5GgSjybAIi7wExbvsKi/
YkrjNIX7n3z5I7mHdjW3+e/63TQAHB6Y2nLzQeTmEv5XDUTSlM35a3hY3pB1
nB5vXR2Hwl/xP4gr85yFs/7qkAigFnU8Ei9P8YwUep6OCebau2pC9c9f8ooe
dLUs5Loys8Sblvi5JjwXDHhheErd/QqwiC5H2fpHtEUPOAuisQ4otBbReQMY
EoyG3DN9mtlFio+mNlL/SqNV1jTPU50GhnIoTitBf2VJMZf9x0tfk5v9lUq6
eQMRkTOBzIlZKwWpBosT0lDQSKCsLf2aEHr2j+EU5txTrS7JnNdPBF6tB1ZC
ufTsina1cPIgNcX8d+KFdiHIfiqz8D1jRPfWpnqIauYcmknZw+qKXwad6CoV
TInY6hDVmyF07NBi8bB9VVWDXI/gIwA23tCOH5GN/AAjvPnYwHMAETW318xy
OPMsDOoi94ggeSa4WwJd9YU4JRgNRI9CsTkFw3vPzc9VIh3125Hm+B3sG8Vf
eAeBlQwRiFk30o3qTo4fQldpc0bIqlnWaFeUMn/Ken+Ajb0vQUkUz7QeLnO6
yiarczxA1OW823zx8UphisVD9wFJZkH6tQ26X/IwvdAZOXA+k4rcYocLeI8O
4jFV+LErOfKtdm3ygj+5V+omYef0yYNUHq/y+3/Rcj4CuwveiC4QRjNAQ2oc
iY9BhT/FzCXNWpbkcTx24dvxSp7yj+b1Ndpf5SrQKH3sLxZ96d/CDsBwADzu
STOQcdxgS1+2uGumQGQjJ188fxU/gbSgONFFV42fGQ4H6Giy/6bmv1crWlvo
U4A70EBCQi9euicyGpoRNOnnO3WWoJTuETTwd/JpO1sEPk2bJtYrq1lnq32E
jth+TDn7r1lCngojSytl7IUgIlvM5/XBOYjgnizU6x6EarN3bDERZUQen/8M
s/m8dTozE8XDHoKUQZwj9rvGCV+hCnxJLLoTv8biiSJRFrr9jiUP/96sdU4v
0Ebl3cUDqv3+q/tBnQaI8etyIi8a5UlK3fTR7Fh8e61PPwORl+XMnFXK4DNt
9WpeY+nNY/b6noIzxYzW6ZV1rPRhhPTwWByXgbbFhXye1uNDMl1GqKXtsvc2
LCya0Fk3RGlQz4/r/9pGs3/kzYK5hgBA3EPpnu1PslskFQUhnXNJnnl0UFQt
VYgl77Ez8QRpAEOygHEcHGbdo+zFApXjhM0CYP2jd4l+s7fGp7nBbItQ7NtA
s9djk2JiB+AvZ2ejcELZcxaLC/dluXyStVABfxRZOyhamUAaoZlP/ry23Om7
cH+K6iL/CzyvWodzGjQ+o7nQFpxYTbOETOsT2vKu6zvtQ3ejCMn3GGSWB7Vr
O3HprkR6nzqdcLbvkDT4xsmkWEpa8FDgUM/3StDy56iUpe+fAfDkyaaA9M7R
dfeu/lUql9IkIjhUkm4PtkiiarndDclNeH2ujlnNIc8vtTXvxc9ivW4RnNWG
6vx/46nhi2SgCHUvt40hmMW8ApRpbPHwId8SQ1AtFMEDiVNAXOjcxZu55yXA
CBokRaWmrdrdl8qbApki7D6iroDEPg0LbxGDOF46VD0RaeBzppBTkDgj4fEI
htfPW9Zf4K/64LUVyJmoXfebuAMeYQoYxzXy1Yk0HphtfJrfeW+EQr7X6wUF
fW/Xxwga3U25V/OdI7BlYrgdRVMMF8jHGhkD1XRiNf4KJc4JuxJdW8hP7kwk
/y0PRt2IksNFTThkKnPaoUFU+grpIIIwiqOnADF+VXhgd0qmHEqgP8c9qD0z
LucT8QFC3ML31x8ojCJaR0uNIcIXmnzhvegu/3agfvHL836o6tl29WnywaVk
DTNnpWKEJgL9jFwJN8fzLDRCLGCv3+6RLL8DhudAgfo854n+YGhoWYLhoi+m
Fi4QbYyjyrCGkL3mY5k283yYGD5gmqlhEQJ44uf1HTi0mU160a4mrj58nYbf
P9VDRjSDgJ6XNO48k9NPjIv9ZYnJ16AifxdD+yxh/JR6zIUqMcSyG46wa9wy
nZKXwS71/sPPGQ6XHFBVc9DMH7Mv03B2+TZ8PzoriX39lmqlOucXpgSfdGBg
49EFvMosunTwm1571mHDEKeyb++MnyrhLo4DobSyY1sigx7uJJKNrWJoiP/w
//Ocs0vvKD4alI0USS9FATguZYw/kqFvxIAcXLqqMO/TgrHnLzWKMVsfEuY1
haTH7n7C37zr7NabsJy06RKE8x23kmVVsQAWyhniwOe3JF7j+iUhMNATTHpM
qSdkOXE0L0Fg6NOXxYpYWFvq8YeuUtiFpUTkjUoso7ac2cK9kpQJd9/EQSSC
JMe5jQ0cG+tgpTkl1zfYG3g7jDR0BugtnrTsk+XPCuCFsW0+X+s39U53Rh/K
SqBgbpVnS1lxC27h29Tz5Dfa+mxjWS0DbRLLqqeK7KXzB2ckfGgjhCd0tEdK
3z2YKlfP9ml/GoF4j4f6OG64nEl4MxGwuEG8aQdleatmRUS2b0VL0hOVKUNd
5JPSpEQGl1RJ49teW4KujfSwKUbCVMDTm4G/Q20TUcPM6d5nXaq7c4LODZl6
AUbJPZ8mkB5WR+7VCWPV2sL3qAbE7rGzKb4mFRymuF2+6OULDQnZ+ERSJWD8
VNEmj+2/WGGb72AycnvB/bdpWvQjBWbe1KQ37AZT7LwimFqUk+IxEw5ZI+gh
wK3lCPfy/PawZK6r+U34nSO3PWB2Mp6OIk8FDVQWSLlo8eW1LxiMMjovE9vL
pQe8xV2qt9Dwxk8XXYDCAL78IFltjzl/xfB3GnJPOpKUygEz4ObOCXm1waBy
vPrtu9gFTkuMkDm8cTBiUkkSpW6SvTg7Xs5gy+dgO0ool0rl655anYQU/2Ru
82vrlKmouaofaFMlIYn0oZgdRL02/8JzoSA/Fi+l6RJMWMjlYgYN7/YxIPDq
sTr1YLEh1jXOc8ECPuabOmE47e0Ft1b2W6OKu1YWokmXRRGWMCHETyIK8C4a
BadKPtGx0S+r/maUgCciMuV9JpFZd/PTnEDY1Hxx7xE0ajFx9h86StD/cpCG
2kt1o0M4vqtjb6/Hl7DnUdfJxHAgIoYKsLHP1DVo0koTXBFXBuk3DgYhX3Rg
m15MfJH0nxHcKoNWmTM2qkJqcVs8Hppryspc0QoIyeCGzxWuLXQ7ytDVswL3
WdVsoC9K26VKGqJ8+dgQa5C4JLulb4Zj5zId/r5jUS0nqkDbbFcMVXv6xSZQ
J0eQVQ1awjYi3gHBfiYx1zYY0LbRZQzYpkn1cvjMnTCHBD9OMngTVU50f8Lr
TjJC14LOJvGlZbFq77YqEkLsLDuC8glZmqmXsI0KUKpBXgX0kkKaGOBRARxc
v8USKmiVNPVUiAq7uomv+foxEXfUPlgmQeInOJOmPP3SiDJ2HRQIIoAjYxAX
WfhSJ+Tzn+p50+E31uDGjuiYR8TDfdnvAgffZoieEkw6f3bSgNUlVPaye8ZE
FLjNj6tBoHNbNoHap6vOlUITP7N+R+eUAICDIY83RLN2aMDmYs62jVGTfS2o
nJyy8Sq2/v0wH+M4/zo+Q093T4YpLXBcFKehMocBxuk8mpve8p3NYDYisnv7
cmlYultlPyqOq3eFFs2VuRf5fmUCLTEqe8ehWAyvKgvzjogSgy67ZFUzcEkp
lApys7oT/qU2jNMulJc7ftR9WyRwtFmkyEZHS1yeToqrtLdDv5F9hbR9d7oW
ebsYrVE71C2T74XLPpAEWynrz5HyGl4wgeMj5/slWcm6pmG2JrsP1shjLkf7
zTNHm1212STOT7U3Z9id3YqbAOZvdclnro82rwCwP+aza5s1wcof4Y4EBwGb
CCl2MB+bhiajF3bsmOfBmkLNiBh+D4iNBunVi3faAXm1ofNvq5rN5a5ZUsoX
/yA7d5TS0+YDa9i3k093YAltJ1uZRq0qyytHP1hZDY1jauCX1zDzjFjmFW4e
SCCs6S4apCKsRPx5TWndNBIrWDM4m3ZqOUWGl4uux/fKMElCYYGksBzhqWmn
3KmhMT1KU4ZV3wYNuFL61JbSSIFLeRhDo/kRol+bWaVvlJBe/aKLIRkAYKvR
mW2LPdpo6lYE1b+HkUxs5XLeC9fZqoPqqgDENDJX9VCMrinZJ70e5GrcbLM8
Vp0udeghMQvgTIRQVtpzBAMNamfpBHsF0T53ima6Hht6bfIXnWAtoxfoZrwX
w0v+0X7leKoRGrfbdm0rcknmSmOZ4n93PrAEN6Q1g0krDYGUe8K059hTISJn
AgQY20rIij028+e+LIATdYCreAKpoelfA6vMdzktFtlWPpxtGNpJUhKbYzJh
vcLTlLv7oz1OhN4oNIY6M1LldahrPxbU/ikJKNTrG7INhpucN6eykfNMN7Su
peSH74jd4juj4DGIhV71hHuEWCiq67iErjEkdD41w9ekHWJLoxNA2M2L5c3O
Ghj2jY6BwG4bE4CG1nEx8xLt5fQgAyBMUxDdDIXtBVlRzskFEpFnoREGyRkV
GdDVs/aLTZkPE79dYScbbx/dJuri1XYlyxvjRAF9s144KnbdOWqARce6fi7s
smmj99THmAjby25v5iJxQPm778q9c5hMySwIbdItIto4luvJa3WeBzEg/BGp
D3S6cYTFDOuE+L5U/hvfx6YYQY10Mqomld8TdE0KmgaxM++jtODtpjK5f92r
bkSKvR2N/vk0Sx7utwYJrjXD4MUMDeugb/w3teDbzKAjPG9GXzT4PW6P/dPh
XxX9pONk5yVVY9ADAfDOen0M2B3w7jFBmewdU8q8EaophBlCjyOXkVJs60Ly
GShqyuQuwP//oSg0LjEBPv4UelHOAlogzOQfoFcdOh6/ne1cgWtqC2FRdfxY
FKpKzx4PxN4FVsELRQ1FlivE6AEd42v1nfEPhRcqh8Hbx/pw6fC0G3fB6idG
g3OuCmjmOEHxB9ETi9Zpvwo/Gc/D+04MpS2atuqEd96KwttnWPvo2NbuzZwx
nR756b5n6wMlY6GCl2AIsvNRINX99OhpegeVURTImAbRa0E7QkhzdBvhGvgh
Ny19YwraFfd1uJHxdhRTFDJwmGF9uDNue0yidjPPXvu8YzaKLb/+F1CV2260
gZbabwaogHFYQ1ymd3MOMppItFH89JvPsn+t+LlJclaiin3525qRXC38LBaw
Q02+yP0J7QIOp5ZlA+DFvMuRIHli1S4WdoXnxdRM9qHiSp8FY4MTLKso74vG
tCJaRSoY+HMAynAQYud+xhLL+xCP72ZdhYqirlBApCuPrMSNe05umwhflwIi
pf1vJA165aWt8Ukv5sVnVHiTl/D2RP9PhnhhMv2y15oToDoPcbwUheGqCpgc
E1B3lOm5nfdLoD/2RfnMxLmboW9Jaml10NIG2F4+9oZ5HofRXJKH7AhnLogR
UDI8J9I2BCrH+SEPp0mj9KyJ6ousEk2APxVMdffIS4OXWUfwiOtTO89NYmCG
2N283zw0MakGrtXCjdJ6SpjInKgHaGLDIv8C70C2GH38jFd9R3RT/WJ6KltW
EuUisYfDQ3ihtHR66m6Ner6ER4wUxDXVzgmTDOpQZReNUN8av+RR06li9y1g
a66g+lXH32nJUm0u18UnjWyd5bjrYo7o6NLKnc0eurYOItcKg1XZIo0ijUVE
9qRpYRNa45HKowhEO3QQ1yUiIEcxhfiYyM2ipqsdXcZnELqL8mlOQddJFr/V
sOnCwl/cM+ezMo90X5J39qUDPo6zQVDt8/FHnqFNFuv06g2/Ea1s1SZfutXi
4nKr+YVpb9wQ5dTkLDnIihvXVN1js8Vng5TqqplnwX/UDLQFGFEuafrl3TWd
Dyzp7PI3fy0aicazjubmi3iaDD2bSq1skOigFrvhcJHvXXpmKu1B5XtpmodI
hcYXwcoNokv5FlIS3X0YZNhyIREhz0bn/OdgOMEcl3H05MBbVOBUkI6Qj0DM
mnEiJsZlFYcj69qIZZj5m86Mt/35vGxMgh09d8IccvH5Rvz42mkq2ceK0rin
S8IMCJ+4SflQFU+D9ed6WDaQDzjLfEouY2EUk13ofuXEn8MvyDCPYVHYFfj3
XOjcEDVng6055hii6BgLmI2Rn+cn0J6oeqz6Nvw0zOP96vrdna/Yq6dGjyrn
MiBYjSKcRqH4snAU0lk3QsWVlQcQzIrkECFnAg8TCrzwFxgAMen1MhWTvPBO
KaqYuQkG93Zb0Udwma2UuYrTapkMt8VsnGC6q2t+r+Pbm0yUpxy2krAp4n3g
OJzkgWH0A2ZIgo3FFiWrT6Bu5nSLXtJjlp20NVO1SS8KWAftexEUrX6UjHYl
Do1BylM1ipyof/DQU9D366eeOScEzDivABh+b7M6dMIiJgfGBr5wdrTRMNnG
H3nE9JqWoAdRp0NUxoA5DlIrGj8mxtKmZ2htQPGFfx3560xVNk0kov9EGSuT
b6puThApIA3VcTUhiYFuHEVEt064uRrqw2GMxkNzUMOR/b/HZ8QxP3a/NvVp
aydocmJzHRZBsE+FKLnAy1cwLjr92i3sk/Z5meHUQ83Zswbgfluwcyg3mnIA
UfsvDg/sbRsmWC//egdABMbPPRq2OiuOOHeui8sRNoAGKx84DjFp4NifAD8K
hAqNh4ATbsrOQTUGTJz0+InByd0fZ3dGwX0A0/+z4VCQM4OSt4KJP717com5
/Ap2mD1k4CrrqUgzqsbmhzC+y3oY+iQYDgyqcsGINtnKfh2Vg5LUizdxnsju
zMiVD8L8m242cP+QbTEWTBUT25xk3uaDCCKcIQuCigW3AXeFSFoXm820QuSz
4G+cS0kc7jVovg+sqzDAPL9Eq8vb9qng/IuxXKZKx5uu0dxMYvGFZlieFKie
9sow8dDig0yqIgAP53JWQZBAjTYOt1s5hGvvsuBPSZ/kQ8uSp+a2lDEombpt
n/pNUTLPJqzKPNFj3w4R/y3FV9LlmMrkhrtg18i0fs8TvMJBA+KvL31PBdM+
PdqK+SLZ+gTvY5SNfDILLJTxOv5cPUFwYZFqQAawN2/ptycBKJcsP9ekDWiW
rsztqo7WqfKrTTb0a+X2M/TV4+ljsWE8K2AjU4KqxpE4mdWS4PPq28K+Brc9
oGelmlXJqweYNGRsWd04BN5ZkKXvQ77pWptVGaJQI2NDZic4b7HwP2f9Lzje
RTcV4Hknc2DXSYyjw1WSbP2osq1ww3wO+J6+0oVZvgMLQ6f7NivlSRz9FPCs
4RQyYThzvCeRDX9TGK36Oj5/LvH27Tj8BOknj1Mx0wctFfJIrX7A5Nmln71e
B4N899M/wu8zUUC5+C67xabBoAx2VSSBNgxsyMTThf5VnNc3HGKsilDYZvk1
O5sFn/B0ATCkzHZcshRD81/K1X1BKZY3YIekRqjCbUd/clxv7rFui5XQzV9C
j0lx3qZo/PWoO8JkrRgji7uT4JgoecVut0amzthYEJbe3YcWfnPrVCKmtDRw
VD/yz4MRSR5xTg0nhW8NGvB2OZBNHiEVwuR6CWzopv7ml66vOrd7atXzYbB4
30Jl9B4QkEj1C+pO4E8nUlUsdS2ebUaNthG5bugqaaU7r5SmkZo25yWzLQhg
kXUZmWd28pUq3pEexVK/XsXbomaJVezXlGzskL26yzwo9tTJhls2hAcrmHrI
vYPA7zXpOND2WnzVLvlGtsS/jk202IABS69K7cfXRYLL1wZuhvUxcgVv2/qH
ucLlTqW87tyz6kDZRh+wS5r4K9Lucnr9Z1LFlyc+RH1dCwanJwubVMUmTdL8
GvVY2MWX24ymZZ3Y+mCjDXjJRFu7Wgb5GVOOZfoCmFMdW7lYcnOS+o4j3A3T
cQqyKxm71Ks6X87rJXsmU3YFt1mC/1D6PzCu8IdLGHmwWA3kTS87ip9e7k+S
ry+npOLz0m8cfcolsbO82gz7FzgnC0TUraUVnkEfIm4LHqXavikqKI/2etaz
Rcxn832M2bIZ5Iucnrspx+rR3HpTdUHOv6KH3ZChGgUy5BDK8IaKlsXK04Xz
1ZNDI1eK1YMuCOD4aey9BXmq5FVUSqpMbGUWlKI26CgL4Wb5KgbuHHv+Kdq8
YFAzkVvMVtkdyq0g+Op1zTvKmNgUfHX67K9pb7RFjojiLMrQJ4tbIzx51vam
V36tTxQQHKpeodD0w+ErulLwmQ2BvWi96sueADM9NRCG5hvw+7K6RoqyhEsl
q6Vt4UogQhPpbCzVesfZm915z4YUJrujwEU+oyrFVJYfq0BrxI1J6F0YpNja
wAOPvk1MBf7e54ytHhZ5fJrRgEO8NBbWn854BULWWdIvxza4Y5AC1WiQWohl
8b8049pPfXDkIYz4GcAi0bpv0lQ/5nJSAXYjBwr89GkfW3MBL5PNQQy78lMX
WRhCExFbJ0khH6FLBGDn61SK6Upd8ARZSgBOrKSwyAzJYKmRGghn9XLv0ojG
M0x70IAsEHHbTdBCjJ4oFGeQa8gtVLbEU9cCrbKgvvDWS9IDwJkosKeowDuq
oUmhCprYDzqYhErSc5f0nxeIgaA+JSCGBvJmr6GTNa5MDFVYooORST0fKKVg
U4q18b0NzXzv+kyp52lVEYgZ8AYaigN3MGnun2lc1IsECt6njXf/7SKh5uza
uKJoM8ivE0y2hpkuRhyGU443wCp5w3pCAWEzqgHsW+A6AC9RmNGVjf2PDQCV
NVazHb/oZLljXYbacWON7qJ51TIVWErXhPj0RSdw79UyE94Bxaj5OBHICaBy
fVC5HMFWvDh81kxZx8M5o5gnVf6ibpA5Omaq6K+AqF4iu35dZQ5AK/dwag1N
tHpopa1j186gFkaX4vhlQwHFJNtD8eQj19CMHwpaGcNQcGirV5bFreJw5OnN
xmgljQXSby3pQNnNxpjdnPFHcokXNemsXshJQwe0JWo9KbQsy3GT23M/ptG9
RRVecDsv8Dgzd53NXPKOvYBEc+/2IidnzkkGJCPwvhhIUmL1rE9xZNAikKGK
F+jXoAcNW03IqrbCnZrfxo9uThtDGHmp1m/R0OSyB8igeR8X39wLyrtcSSWs
9tAXMfIAFH6c+0zAB+MxipyzX/0buNkGBAT6ibB8s+irZBaidzS8m/YEV+17
yl3+jgt1X282ykvNTNqwTs+eQdJjaA0wKNaVuA8l+Xy5VyU5LL5QN0kEKSab
2nFI2o/zfxWlDN7dBK7CohFMDAt/v1KY9Nq4pDD3VtovoZwxBqTAFIdQBv1s
HSBIQCSOWnh2eId2BbTzuqShbefH5UB6TOPku0LHC4v5WHJ+yUugtgOyNTOE
Zw/X5XYkZFXmwabgBI3FajV6vLpGqePhFFxAOrY3pW2XuW4jc9R8ICzysdtN
7ijN6GlVrZ/I8ghaSKsWiljq3mPUCrCOQicfNWIu0oNsNFd3XU69i+G4EBXY
AqpJ6rr1LWgdLEH/PNwPI/yrHKf7/vnYZvSDtNvxeDWaWzGb/UbwApQJLfD2
ZryjViLCBSPkWzzwTu2jFhGJbgOFfoOzKczY68llOcLxLRBXqe4FzoAhq86O
RalzxWesgUckKZeG4euMsdvvfprhm3k+0DLa/rywO37v1iPGanz8XI1tmLbX
BWjMUecsrDQN72llDznm6cKKYp2iYFfkflLajcvOLpRu6fviQkXuD4bvZ/Bq
W0RGeKqi2UJblt52h8Gkhtm1hyYVLxOagF3rdvMlYMgC+jO/e2DKYeY3tUd4
lHdXGixtUu4ZgpRK78iFGJoJt9h+MoD8ph2rYWXXk1vIofF0Rb8Z+XBWI1By
jhDSPaO9+TwdMjghsNTLeocRPeXVR4O7yT60xeLY/+W82S73K3Yoilyh0URE
hM5myr3M7uZU6xWglauu6tvrlA1d1heqdIpVI7L2Utg6ujIVGZGTbQq6qb93
lSKYtu22ERDJhFzpTsz7cQpdX+x7v2lWwDHYTjykEmvzThp8lpldzoyHV0Pr
4BwEYBrT3mkg5XjdMGwEog1qWABWwo0U3ekVWO95l7v+pVioGZbpLnQu3nq3
hfVXuu5fmJ2tD6IGYjVIBiebg0GlkThu8EXStmWldgnYuLgndyGkxuknXWgt
uzD4D+pkTzJEX7lNX4KKDg5nIQ5P+Er5MltW0TeHJ/jN+L/eX4SiFQDHjIJy
VP46VYJ8bcMK7t/03qWQqBB7uc/p4AHxwLWueK/enYlMoOXdtF6GbSV9k6eq
TL2qbzfZHa5/LRqfhu++BxrGfSVcXU+4JBJZeaJ7hmXq8tFbDVmmaaCSxI7d
da0axCHfRx3+hU3Px/lECBPd9ZcI0+RPNZqk//5Rp2I0J+GmHMvHyE/uAUf8
6KpoLbgFjU2ujY9eB1JRJwojNZ0UzCwAZ5H1mvQ6sC6vKUPGb/GBoXI9JP7i
kPZYbmRSl8hmhw7f3d1NEyMUliu/dosazbzvIUI98088f1J6Y1WTsEtET1xV
BxbITBrykIS2/tWpowb+O9LZ7lfH95VPKveQH52bt+GMUQyhlIws3mJ+Tr+w
BJOy/Ej6gxq7J6HKFFsIp5u1PqZfz3eEikxInS0dqDZ/2Uw6XbY3IWyp7v7z
/B+CBLcpTQWTSMTeAUkEtCR4D73QXFXguFHM94l1JbXYowEtzUf3OPHO3mAe
tpES6UZ002N0shz94Dj2MGEGU2Q8iQ0nK0G3NPr4oYna+n1ZNmBEAlEAL0FG
yYNMxQHgdEFdd06DUL1d1PsUqHu3qFDqYdPS27MMmhbIMSibNqSnAmdnLvhc
t9yMMnrY0gMJ3fIOxE1wMwrOFokLJDVWuh57OsNR/15tZ9aBjbajVd5fAbqM
GANBcxvXBoV5lVaOKmTLIHlN6RzjSG71pne/Fy4cNkkNMnFWIeWm5O4i98Ns
yRC22WY6ssUBp3975VMi+dOJDTuO7EA5806n+ZDTHKqhyiJmEMZyaxEQw2n8
Ud+0NlwQtl8VPLUvCQ5gsT5B0SMr+cqO85pKmI1LH87YrJiunqX/50jRwW1Y
TwlzbERd1vMNGVYMhzeiAQ8UpryV264YlcGeom4DKhsiUqVuqSYnf/pmAtF8
I2FmllbX5JdyHRopHsHL7wntkthd3YXIckiyb9DBkAUX90NhvPRaC8+FAcv7
v5cX5Ob1lclHhuF/GIU1TXSrWSoCg6fCmPRgS1fhWenAdFBR1Qum2XmXTcUf
VLQsHhUB5UctWqr37Wpo6B7a42eFj1yzKI6aIK4MAIzOVLxMo5hMQ/TUhGiC
ruOOrETX1knXYEwE5dYgIDUI7TLHmehG4HRa6F3zBRJjGRG3N4aOFkWy2M++
C/QoBw+Uct6VRybOp3DCNrVnfKe2vdvtcECS6Ys2eP2pR7bfYt7axwPP5vMp
eAjJWKv1Xt5VdRnPBKw5uuCavmor+1cNQmpVODIW4ocFBIYHWZXXJgQBjWYD
AxY7fjsaSwfCQ3cECn3rLiqNGie8ecE+r/BZenQJEJxWh14BKman+izclqGr
j3sTgTRcAQ74sq+PbLv5jOzhhyVPImwIzraA7HAIiyQEwz+q7wc15q7J4v28
pfb5OBbZxY/RICJDP8Kt+iaQMhJXv5Y5xVjUgs9xlcCI99FwM1kLbvec9dmy
Mb+1JjKyxiHiUBP2p3qdLzuAx0SiR5+e9y+FJmmIUzoKYTVHBAuMeD3Y4fHj
xocvs05cw/U2lsGNhGSRGjvtsz+yo0QLft2k+mB4s81F8KlMuDs3wVDBBl8k
yRL8Zfdphxhxn51t9Idv1ihBaMLkEpkP8aaNTIInw5yOaDlSHwsEi+uOUbz8
TIYUf6ifgyUOq6AvTVXLpZeo5TN6Hz7QrzNr7wxD+oRlCrAD51eimK5mRMtD
VNDBp5tlLmNk8XrjMYs/InhM85yfdZknD8y7mZjyVNxbLFWGtywA+hRPKyho
L/IEG2CUxJW5A7+Mv8Cl/TI7MkP37FNhm/g9NAaq5BCRLJAiDQ7H+6D0fwfo
lShSldBAZ6kdNMSLHvG3d+QWlmo5MCm4ikW5cbZymfWUgkaymaZN+yfieOhG
UpK4x5a48XiDN9mrwNQy2PjbWRoOYWV4bUjyNjJ/JLjdbAbEd5MZaJLh0r6j
fcWgxEEMdQMW8e+2h5D8fDy4LKhGyQNtwKvXAZMDbwqk3TJFlcBC23KR/c7q
FHj66NxoQgNlmbHRgxh3MJ/B5hpEc4Ew1gkrRbD4xEWbfUSfB1X5BiLJbrZa
+XoVIFpEpNvbBRO2S5OwousyEZK8r5KgCzcOKGvRmF/BsWNau6v83dE0n207
Hy0/PlqZlFpA272QOjSliUZK/+PEegY+XWu6tCAcR3BubU2DiMcHsvHVzkAY
DyhJKwnla1HO2gL0mTtVAbGqPgxEHAqu0gSukvbxEjae1dO0fb5LtWMF4bTZ
ENGqlLZISyVBA5X8vktTaOpQhuVycA+LARapU9BcE3XJ9tiN66glz/uGbPYn
Vx6mmuDBF29KkutLekoLxaXMEmpBpWqP8SsjeTv0OA0pXqEoxz47CuZwPdWv
j88LW6XHauO/Sq1zk+QsMwoR6f9/wwRGeKImN27ova5Wwn9YYqxLX5av2PAo
TdcFI/KpYyhg4e1dzx56U6JoNq+Yeo1x1xRgP9eZjYEmr6y7TN1xfDFX+9ZF
30DeiGC/xV3rpawB+s0FlW84/S2Xl5Hc9B+I85c/WLM14g3z6W74k2ktfacz
34y2gtSXqfHW+BTeiaB/PaKtTtVSFtvi7K5yTWqy7TknXuRjIVR4aZr+JtAI
KaSbqk7UqNnD1zhqHw1wxZiKwRREf2zFsztZl/aR8bhhL3cPO2fsBtIbQ3F9
EfpqtNAkfQly+HTpgl75fCamfb+zp7bIqgz+z6O7TrFCoqAu06Qo2xdG3ZWZ
4AvdE5iF7JVP4hnQzeFvMQy8YX9jA1Ymf59dHS6qXCvZqJU2LkUjnBUxSWjy
iznNc0oKTilJfYubasapf4mhTG4SE/sakQ9CjIxfzcSOH8H1X/k4GncHWt3I
NO8zLl5mZJCbinM8w8a8oa/cIdgXbj+IPFigu4frIpCpIws68WFxQLl5Qnwn
44q33qsfb34StJcrLavszFngll/SzO3ajoiXFn9Ou/6FiPrvNa7X6LvfdeIu
brNe0EIBZtjZLkc0JesIe+xiixGhkPgGaJlvvaCnsw+y/RaYXFp3BYohEWZY
HUhgv2Hi1WDbzcIoj7Dy+CEX5mynCJy3wRzR+AeHctyL3oX2l5z+ZH1WFTOo
ZK0GFr/q2PmdYn+HjX1d+ZR9Izv/L0KwotoWnraxB6vunk5y/UOLWQ8LyXiL
UF1wb7gwUtwu1hEuLTHWr0WLxnN2ojhtsauPY9cJOlShjiIn/7kG0dYSvSN6
S+3fAv5rHo9SLYe8qAgXD5poiZ84qHXJmxOkDGnSbyB/1binpfnDPIbhlZiy
qR0iyxXg4Vj84Ru61ktSKOMAimyyq0369CHpt1PqzEhQ4mk20qpuT4fcbN/G
HJ9nkDZfFkQS+Jlj1rHCoWuJC9/ezR/kZNaRSQB6zbAeqUDPpUtsEQXkg4Ys
/K5B/SeULC+YLyNuqyH4whKdnpn1F0YccGIpJYXs/i6EI3ZHXnWfRynPLwz8
rVz1FdS3yrbs/ogI5pZahvjUGDnJKal0UAOtOy5BBqbAqTpmM+7/+AP8Y8HM
P9DKaZOXYg02qZOc/a08ZzA5B4EMhnjSmjc7Z88BuuWuiXfVxQS5svUdhSXA
mlj/H5q/5sb4pKPcHMla2ZD12hoVfqYiLszUB73/Bl9AP0h5Q6g6EEc12tgh
hS2Elf2Xo3mMvjpJKfrdBv94CfXPpIwbXq3QcD9fYVa2S6Xd8IofGDm1D8wM
hZCr0f5JIXw26bF0kH/hW48f2bQg8EO2ymQWr0UkS/j82KnDcWmHxSQYez8I
SWWopLM49RI8Afn0o/OQ42lR6KQct5DtkjLLL2WbtcMCUyniKxNqtqYlSR/P
HKdg29I/OcFrx+kR7v+DjTLgx10NeDhlaalW98pDsteVI0kYt3IQ281YCMIV
QxTwMx9nOBfXzgC+nJBk7W/GMIg1A4mwYQy7faMFbICiNqXz3TfgJyyhmCrn
Rf9M7x2z3ssTBQPdCNntsHl5/wgivdPLzAlvETXnHa8b2AlFpiJ7R+ZD5qNE
MuCZzA966uPCLQvYff2L0sInfpgsCL//WLxw9wWyt02Tm/Cn2+P3wTLGirEr
1tP5YvzzrOTgHgvwuDv+jXUsA0NVmc2O9vj2X3S7n/HxSi2Iau3bjJztCWNE
8218i3XUzayQgsVURvtn+UTLq4p49qtW9/UnpOdo6fVUv/F1CY8wf0uREyFE
tVdEXnRAk2c3Socvb3n3II6UNRJRqYcce/kMLbvtoCQHV+QlLNmdvdNO8qAH
76EwkIIXM6V9a/TkwpSMf7pZgK+l8/P5ybLD4xdpK6peScRmmOteqzp50qYp
3xHDUP9CFPIRaX6h35FhF5faPNqc8pU1OM+Tb7PoHDSjrILCCybvbb3xgjz/
RhPaKETAhbu8+sB41DI15YLSaS0qdG24s47mMoXHOGCJ0PaphaTV2mgd+z+J
Pw1JkLsdh/kiHi6adBAuwA2aOzudpGxJdrcsTSoPL4ezkZKB73ugp35QbjwQ
xdMlxWyAoRMMxZqyD0Bmg2elCpbA0N5maErLhvhoDyncD6/UdOLElcotXIZM
fI4sVJD5yeF5xbt+tPFlg54BVcAGbvZEGyqBRr6oqS8X3IxcSYbUDdg89+BZ
chCWB1HPaqoiI4Q8Xwa2MfzOL7lUTxUviiSP5lsP9iH0sz43IzmzMIG/0nCY
/IgCmKHoDvKZnpxDCursBiq1M3OocE0nOqN6aIshXF4EXIGUYA6XbkP/E6Ya
PRoc/d7wNpYWHsDFYClZn+dwL446J0EKrglHg7pGBF+S3X+5DwsUlmL/5DI1
CvZfv3BI40g18hCTbFrcqdTFggEOjO1RKuYOVV4uIuoTZHPH+2jL4L3RENxx
WWxvpXPM2NKvajs6dS71DOqlm/lm47gYlu7i2pdF3T3KE58D4D/LtNXo3ylP
lfLhsFuD1L3Ppo3TMR/PgkB6nm9ATvMSaNm5pACUA/Wxx50TB7Tr6AZlCx5w
47DuK/K+rATNUPaeMJ2meJdDvWDUrWXA5d3qebBJvKQLNi9L3gPmiLjI+Wf4
Yq1QzYlvhlciWh8QbnTlMGawE/S1TBKZH53EBtOM17U7ysbZEPzMylfQUa8x
9VpcTPM4h82wLWnu1Oz8XsHynljcwh2TJFgJyZjkDfl8l16E6Q3+see47ygb
24lV1CAI5fN8b67qyom+1bBXmptH8VRN6QPFmH8EflZk2VieETLG1ZjlBX7g
uztOlaeiu4rw7wkfs4tjTqyhIi7AhDkWYmwtjYgTR09IqsAjsM3p7shMEtvh
WDASyJfhJuMEYfdkBZXQqCz5B6xrUpHjiNSy7nCCoUJ5wHICYdzxm9I8BKJi
IF/snLWc8KvHRujvrq4GeSZ6Qcv48gPqVzlVMXAQao88wpOCPHLnfrcGoI6I
jfcdADTXP3dXu9WWajL+mc0EBV0bKSWyIdlIQnWTlE3LlVJZfzRpHMXVY6N5
tR+dIeBzItZZBgQXARAtc55/hZ8LweDbJA3GGXWvvp+EqFdUELSpXc2/bUyO
1eeShO+C2rKR/GhgCoZ40WwjlS+A+4b8SsTBaPfXgcj18vLvIQLU+XzmTGRn
N0VphM1/W0bMdbtBWNTF2p5wVVNB3sv9nzXkkcph31gRhhqmLjAwTq9pFePa
+irR2+/9A1o+fcotfOrXZ/VttFUcupzLoGG1OxjfX4K5UBWIttjDfQ1mihGE
7DCJS9+q8w+1TsDE0wwIKOZIS8TnZ+Fz5ce/Ga2FfHTiKGgwEnxgw+BV0qqj
Z/hvqsngO79ZUARhGFfSQvBQI7euR5njCmBNzEeh9URKvWMhpBoVWfAUGo4j
MrgHBncNn/N71N39EKmmkHvwgHBcmSlM7kUowj9sdvi7RayE7hR+a2mg3MWW
gvKZCI+dYx7vn02k/iE/sTQx70t7+iJwZ8gDgFn9Lr+H9akOdf4vvvkp49h/
4aySMlA3pCy/tTU1JQ/4/uF8fVlBumgk6IS/cu87LcBmwmXsjrJ/1bYvAx40
gVjzaPxCgz9xPMYG2K8KBY+6W463SnS0R02sWOnXWBfymhcFImPyLnXXGrJp
ykqHRZ/6ij9EG4D/YChNN5U99//gDxsvmrA9rXPOxlJIo3ygjT2diE7e0AH2
XPEYjYCb3KXXZu3D9HWiG/r4q2At4xo7DdHkR6/GvPqotpaZGkITxHbpvnOg
0lLDCSMllkdF00dXYLzZxPG/rv+RS1bysEvzKG4WPU43fObYc5IVUFkXU/z2
UOdN51vNmRzVyjNQqIpSUSQzS1ZpkzV1A3htgNgafXvJst25fXQU5s+ZShKQ
QZMXb3Oe1FWKPQ3m7oPINZvNSghI9BAZDA9vFw3uEEV0scbMpVZTpaJNM2o0
n5B+ATewlWO1I10ENzDNrgm6BhzrhQafpbmjsbkZ9tBgFkALxf+/AOOpu1z8
KOe6/GocsFuVu2e0C2sIu61uAeienYrGNPsWBnBYFZtuDDMMult/5NAiymYq
7w9uxpt7mReZRatigMy4+2K5LQv4MDMsjs1qvgye1owhSbLIrkzZtHN9gSat
D3JcDLafGR14zUNvrZ4sC7cbzfWkfhJE9WVHFzu30hN9qIbogWUrsE7fC/KH
K5bPV2/hE18DiYgXDLCr5GyDrCnw3v7THpzSrVNgxua+1YW+pil4lAKYfaep
drwFfPDpWRwzsMflui2YWwUYlWFDT5l03SSehOoC4JcRjVglTAYX2N5wjsqy
HQmsY5Y0ntfcr88BRNxp9KXbDA+JkuvBey+eNePODSo6rbmX3jkpK3oxEMpC
AK+tXr6272/9++oFy7zfl3308j6dimY9WfJTMXYn1kaU/MXlzq147wY16tWe
Z8y21Yx37XeE0CvhmtjyBfa010uxRge0HYPKt/aDOFIAXjqbWjtYVqTUNHz4
XHlixdali54FvwUu9yl+4uc5RmaQu5uWt0O6TXFsrSL3YiNH7llbSkxDu4Hs
5Qcsn+kwliebAt8MTZI5QybzHQv7ylNiBS5sxlcWBxWew4RYFhF5DO3n2Zu4
yuz/VrgpFU5JFcgXEn8+e5f48mBhZv2vXWeCXVg2abeZtXfTKxlUcHaXUrth
OSU+M+N0HVXtUw4pjyDE0KyYxsOlAV2POWLSyBn5litBGZIL6Hb3Gq7wPkkO
9kvcmW0/nKfvik8nRHkQzkMW8Jb03Ds28Lz3c3XMkf2IeOU3lKQGuBBXKE6j
6Bk2wvLefxcjYESvllBaYRurjR6jdTFOTL42t331IxT3u0OA5A+PMww5MvF9
Z2Rd9QQmGSk2jiBgXsfmNzjXSGfPOftO6uTR2q/kFlXMgxAPVu8uonnpWblT
s9jGYCrQY3WePTcC5rIRLEjc28i5rTvc9Az1wRMKD86W7YmOVDB8qdBLQDU1
1A+M2GsSjEnk7sVT9icN+JSf1gqIonYNWqDuSfxod718euoR3PJ7jr7sh+XT
2jlXLCP2dtuJu0M+QwxvUOcmxF1QVXCTeViV/H5ydqpu/QFak6P5RZi0q9fH
dLZW71mZTAnWUGWY7xUmEoi6BpD/AkZ3n13yPGvupZJB1yX+xYWER3xxcxoU
kP2BdhNq8uHsbgHG8hdAQ9LYxfLL11DrAUW/A+Sad4yOmh1Uijr7dh6f942I
V43EfU5Zri+uBiqhg7DxBmO5YHD8UAzUzprZRMhg8PJZIquznDlSv/wDmXA0
lnhaBnSotZVQ6Jjoz5QpNfgAnXFFi/SR0zN3O7thiU7ixWVMf8xzLKz3Pgen
ykhJrDEbV44Sw4PIUZ2j6CitmznIr3P7Ke1c9tVBvP7moBli8v1PBOVAZHpE
GHNPmffriSYU1McKmjmzy+UPlA7Z9fSKYps5ms0nvF6NNjp+OeN7ch9laMtS
DBY221izbNVkCH8xxF6KGmPA5ifHmoy+1SpFMPvFg4UNZHOY+IRFhdLgqm1j
RZT2BIS0giySKWg6DaKZ6nS0DMJw0bOJ+F+HZv24oktBdacWBqjBq7ymmUHo
Y7d/g9nUp++YR34Yjwag+6sIrOaPfURatMR7lTfq7c7PY5do4ZMeEUqzTbWc
/+BEyni+Jg0IPbE1wnZXFSQKkObhGtT1D9GyPoLH/TxoGVoi0SfkxaS7abCy
MnzX62nd545o2OjHry9nRUgZzxnQaRTE8MRL4ibvT0pW+rqTumdruac03lhZ
m9+KdnK4iyi6EEsQ/fKyww+06dSRuiIAfD6Z+tD3292+AbzETasGn8LPI1tu
6PqY6ww0bGDe/HdmkCh6NEsFN6abcOxV1RipqpelNdcJWJ5VtGm9AOLBPAzl
d29nh6I6pt0TLy2Z7+YK/bk/BFmwrK4te2aLtnl1BDUg2GLEsLUw4zINHOev
5anqvVEMNDogcB2fsdv1pXf/9f0BwFDXaO3KrN7GJIPk5oH3wcFCfxUoowcj
NtbWs4rXIbSaZadgs+QAQtXpOjvd/u4ueOIDSgFZOmyH/Ebd7Km1fvyxl5SL
Bvfyn8RY5jr4vDGAd/nDLQQz+BTBQYiPOaXS+KTLyTpoTcknrYgULbo56/1V
RyfdZD74GCwhN22UxJQuW0WcrnXStw5OULNSnqQsco72sAFSim+HJ5wnjdwi
z40lqZmVPjpjq4FrbeBxDdSKRvvpMtLUZzfS4AEf5s52vbR5GVsuO+3DZN+I
j07YHyvQacCEmWFfndNSFzLeWrxejtpEvbY5PS/dpcjW+be1YTy2hFJp/2xx
gNimc2cZyL39iOg0XMaGPfURlnD3VqdX9YcrPMtZs3N504Kfd1d3GvWoQzNV
/h/udFewVgSDW13blUqp3yEgTv/cK7TezbvP+VBv4tWcq0p+kfBSynGdgiXc
ggRF3QDLZeCSwv9eQk/3n+1DajL2TPqajmZsBRZuJ9/FjxsMHH3oQy9GO8+n
paJZVvvkQuRSA5ZlWKc6MeQ0ecjSizQpDKC+ljx4S4Yb0n8k+2f5gSYYlMNQ
JB5AvxSaWTBiWTR61GeEcYsVyL/FT8njNATzEwZbYTI8JtMG1m9CXSks1Z0q
Da1vb+pA5H7wlP8qicss5p66krzvn+I4vzm1ttytU6P2DUPElN2uejR62X2t
WhJ2AoooEm/SXDS1x5hb9i3/ZwCIYEGU9fNYudGCiGcrz8tmgzT24u/Xgaq5
fTunlGtKr40fSQKf/CDcBHRE3agGovsVBI3jarX2SF23yGkGsgRK9J7JV7sR
io31AqBGD5e5Up8cLq3hYvIHmT4EaN5Y5RIYy1BF+yrN/6Ww9WGR94sEdP8G
BXDnzbW47Oo1S3xicTT1oEhE0PjN61BQcHViCqPB1+/mOg/AbhpGbHUbv41d
1VpF/u3zyHpxo0QttcfltFVv6V1rTFUIHfVmzw8gRge/NJI9pyAWaA0B4yus
amqaJaHWjylIvH4Q4qESz1Jp1Rq1uGWXZOdIsOd7zonVByU87HdZOtlVWZ+Z
zfF078v5TcMcwegScbaC2XI9TK6Rn3rdIaF2FpvlM2gB0v8ny82+cRVm/s9t
PBpj0dPMcux5mW1thPMuDJ6MhjgJVFMctBYwJeaenWCvV4ABlG9+TqGKCQXd
a+3u4dAtsR6jQq5xvQxID6FerwR0riYYYiT0gm1nGLKwJOa/gV2hV4od1VB1
R/vv/vz5iAAbvBzpgFF4mTfHYYLlBpo8eVvImMqPaTNrOKbOwxG1uoghwyYh
t8MTaZtbLkwgXCGNDFolfDg56jhpw4PJSvPkl1E84lXifE3tFCD6OusD62BH
YiYXXdNO+ekPHsBdkGjSTMiMlxDJ36oKAsBKPM2HZlnY+USDec4EcyPfDGyN
3Rhq0Z6r1ccPEg9AKG0+t7EkyzvwVcpfMsAshpB7aA0gbRe212fQdQuT93WF
pgZ7UMlyrgnieEHq0EdEkL9bPUlAG0EqTPrJxlsqcoTbxPMXFJtZNCLPaP9A
jubR88avardMpdST7iACeEVJdGEbl4jE7G2E6Gb9TGCsuyYT4S8f6ESXqcDW
5Rpo8NdEiXT84PjoCc6UhGiEwrhw6qAlsUn4E6pCzjQbu74V0kDsMOtsugP0
F6Wh/5NCGDFyew/ekVB96BrhJ6dM76XuDkqndnZ7zRjR319SjrQMJBFVn1sx
qoxJMoEKAOn1+Gn7vSYP8lq4uSVGTpBHw8+xE6sX1+Wzb9WqPFnF3B02A+yM
BKGy8y6ndNqz0T6enIOjqkKVlj7f7Mx5sy7dUHBQoLvFWDdCKH5pK6xi2iFy
vUaYMfoU/sM9chbiGcZ/T5LRCU+bxMKD3zs19StJANLHhGfaHAax5ML4maDa
kr+DKcUspOmnfjOpUZyi41SgPAVydFAe4fOG6jYTkBYsfxeH4e5d6zUA5vAo
zptmyg/nv1i2565eWF0/lBDsCXzFLncvHatdUNEdIDK7LXV60GcidkR2aL9m
JM3WX9dlhRn9kpOiASsOdboe+moqoYqQAGvCcdpfboMaTB2FZTJ7YNLUq0gl
zyLB/0LUpP7HeNi9FBQzDTKubvOKuOWoJ35q9sKNB+Ae0diWSVBSBs691+4K
M9BCQipgHYPWRQuenTZ5MbCaPIOKvt8KPVqs2tMm3FmYafSSaeJYyHbptDLT
PuMSC2U7SR/DVmbshxBhX64UxFgcmLWt6qyyISpwzXWDRiFQlhwCCee5F3Qz
mlFMBcLaHWIASLT5dE7elGVG50xzTuRqb08O03ISBzj62sjdmLQla76FKhNX
CpWZcvJ5Ga16JcukdMqLekBTsZkHFqgEus/f9PzmDl1jie5Qon93pUzj1Icc
ZHqSNZzScvlh9r+2JUggHBbgo9GKU1mxRKJ+a0hQB40dDzyJy7dCzycLW1Yl
F15yGANolsjg6UtnBtVp3MEKJwTZECSRaJTsCIzDQc8m0E3RiGKoqQIEmxHT
N0Ic9cLxHwPubt66sS5ubtLtYO6MvgsFhwsaqo63dhU8DfHTU/iFXzx5Twwc
qlu8WSo6ycn9KM2X/MOyZF1YPZGQ/6FH9rMEIbuU7YjjEwG4fpTDU260NEzu
DRUEENUjdeWB8o/Pt0mGKFuYwZCoR8LZUSzdd/PHTk6GhQxsXy7KUUHh9i80
jyNs8g89LGQHt1NU5IoDUv5ygoYoif8rAlERWtCJB0twoyuo7Y1kYzGfyAkU
qQyT02d76HS6AeAM+FxO8AxiGErRly6QJgWKA3SxnnWud+UO3ZdHZjGHqx/G
KjG9TrOs9+cKBaOEXVgDh7W0LCVVmKSrNntdASpMvdpx2QbO5T0B57EWRSoR
EsQH6BOQEYZRFkTzR4emiCOgbgHv6EpuuxwidNmWcGi4BMjTQLWvxoRs/jyW
MsJlxuD1PoxxsufCH4Z1dpqygnzHvFG5fuc/eXHLzZinKHEn+iPQvgcJwNGd
GYxy+ytzkAaIzVArHLIYZArfjqKElHyzh8EbryvI7568TslkNGqwpvdP8jNP
pEmboN6qdI+LtbtN8+0hZoyH01i7SnQFTxIgAxcNp1zGUOngV6tfbUeokywC
KIShApvkRSf1BX/4AGO8B+uwUszWkeGKbcAvJXFCjuMqcVXqleJAdlf0pHLB
K0/qXoGvtnvZ+0nIrEyejN/P37UkufLx3rmKCcPhRa4zqXExDr+H41e7s57N
uPqN/GXkPNyMRHFJl0934XqwXWuYzeTVjzg4g/5VmnLdc8kruzEet9gOyQap
LYQGzJ1FvwT13Ch9yj+AtXpHpsiIRn7JdHZ+bX5qlmoFdadoPAlkEJ9tPdCt
ATTU1D6qhQZjqdOwONS5KWEWw5VpHRSCeH8o9y8t/2njpx6ZYWiIpYe2K9Iq
qmeeEEAP5CkoFYu9X5TlI3DWbOiisJrU62+y1O50+4nza5m6niggWHEynMdL
mZDomF9sqI0SegJmPxHX3anyeE3HaOoHby3JK3e1Zv6jquLNlrgM0Z2ROuh1
Q9fcy28NN8xD06RdDZfaCGzy71aHuP0nX27GhL2P2Rqi2coqUuN4858Bc1uQ
KsD8HmGNqiHv/RM2AaovZc3zQAg5kueWtXRAiOf4EOTrDh8IQ91Iq55ppM/K
6dWvddr+LaVIf5x0ZJkIg0AldoPXbjbv1J2dcH8dd4diUh4JTqe/c14tdWk8
2+MczJg2I3C6XqDYX1PoSfY+UOaU5ihAcfQ8zFVbei+7h9uzhSraGA975Gce
GDGdzX6K9T+Vrdrgz1MZUrlARe5+jmuP4vLzT4WOdx0MIMWnKD+T4ZA18YCT
8dIpuMEv4xtuvm1mDf96eC4R4ujR8xfBBeXIuYSJhtf3El2RatG81V7SbHcd
TXoRPkiTQAmsjyZVG58t2PpuY/rK1qescYsa44rH0R3pH2Nu+nzEZESwzoid
KTpzf4QJ+F5ru1QWXb70Hc3viOKy3PL7XKy9dJ9U7K7iV1PbXb7ekIqHyc0y
pwR4D709NixelhyeeXdMkevALHbwILLDbTcXFOTgVCSZtZdfCfE60gjGXWtU
QvvSTeEcDpRPfitUlCCV8J83/NegC1kKh9Z/HfT6Dywh404/jX+0oj+Z9dtG
EQqWNOVIUrEPtIBV49D5VdqQMDyjc6rlBtefEhHT8ClV0Jr8h9k6U9F7i2fl
zARIidTpTJ3axhISaqLa8ooD9KCIyeM4cG1xEk491qMS0DrHdY3w5kby4dg/
P2vxPGHnVz6UMFkJn78YTI400gT+GY7WR7ycFH9LoZzLAdNfp0pbBynkOVKC
UbO1hAqg0s8wNMvlqCJEnu5c3+KZ+2obDxVyz8Bp/dGSwQ4Fx8AMbDmFuyZv
A9JZyubwwusyHuNT4QPxEUdlFn117bTd7rrO6JYRyEYpDFFOe0DpcwKZmtuU
z1sDEn2mTRnCuidCMTB2pvoul5vPuW7TLKYkMOMrTr5raPhsF682IX8OsMUW
e90FLGWpG8JPRM3C5Q5NgKiitB4v8cMmsp12fJYAj64HPPjbRCzQq8okEyke
Y1gz07P8l1EZOZtIRZ3dFauZbyagl+m8v7AxR+W6ZDaF0CJBflOLt9lTlK2V
HJJo0iahPYdJKFGhNDwuz9pgCQ0cjyMUwH/uN6rGiKbCozfu1j9JhF+kWp2T
lPx8dZN6UExDAz+ZIMf79T4Nnp3Kx6UFYFChHiGK+aab889xeY9dfnen/cBm
S5kq7b4qH117QuzDPTjV6vQ2CU9t9ZRiSuItF8Q94u1Y0iLCNiTkVXeCMssL
kkGsxf8Y+CptH87uuXia7gSmTCq2ivVVMVGaCGHVdjehSEHkwNJqolvXZmYX
LSMnhfyw7eIwOcd4RJpYFV8TisqPJlSYfbjMz7K3IudP64uChPGAm7NfOm+H
uEb87N3P/Yegu+Fk7hQKiUJWBPt+1kaXGbIbdhwz2/f40Ae4f0wvZIVwurd1
dYclcUnC64uTTM0g+ofPZz5e9IRFxfMwBLAy2O3x1DNzRjVpehPkx7KLX7KS
BQEd+XfCiN4yAB8whmVGntnaMXFuBKUCMGhABxwYSylLfkcPvY6Lda1WZyeT
wqYCFJFimZoIRLLJpHi7tAhd3ynL6FWaIajWbJm0CGKKq135jCgX4Ao3plOh
IFy1CAB80MgLbOS/MN2kC/QEcvnn4LMWqkqvmtd50eVQXUPXQMgeFr5596dd
JZvJMDWEOR6K1VX/H2XJ4WKQebghkHgj6JXMa8NZvjWgQkwIYiekoLGgQez+
mJoNEWgjdHWeiV1LngZ41AeEdvwgOxlC8DzN7ObUTIS6WFcPGV08ndnmv7Wg
QseEMlviio6bYLRvI4A29H5K0C7DuiOBAbORWeGq9p5G3qUZCB9ykm92+EGh
8E5oMl8s1/tFXNOr/xAn3TkkvbC248jaIec0ayZ7rnSIIrVCufCxD1JP/r/o
Ac4UF6uOAhCvAAs1IRF490lt/sBXlNwopghJdnapzcXOxu9chkUkhjC2WkNC
MUBZo+oMewBf5O3YMWXbW7QA2g4XsMzhZLzFpVzThYK+lOzWdZFp2U1vGHm4
jFAWpAv0bDpatUTLYdNASYTOmcI2YYHXXAVcpHBfuNqRP4NERdGPozXREfwC
vbvxnL4XXavrVaIOKneOWdyiLsQZAyTJmDwRW5AomeHUe4WTIJPJq/cibL8a
jwVVs95C7U4mmX5UtUZT3vAkc0N6eIsXAYxafmKp6fXZTzu0Nb0ePpzwyaXk
aqyfNKSDiUxKoMmQ9UKhpKOuDPNeUCTYSW1q0Q8dJleukon3xMl7/ahqhhIH
qqJqsRKVZld09Bq4dp+wcbuvN25hePmmKHMy+QUn9jEjRWO46m9C3MBjX/t/
TdiDYkw2Hfe4naM9dcEE1fz5yW1tya9ld8y2579vxb08k+oVX57oHaW+uJGd
7qaCNnSU2Z3oZew1E87Al7ZyR7pZhadJy/q1QTW6TnH8MQv+pIexyH+2N1iK
E/rhbxamAjmrG7xhrVHvTAvQNY/rz2UnHTkg1WLLgtIU0v09Vfawo88VlgRK
KwKUobISLH8Ucp7FOar+pefalhBHN5RTAwn05p0B8focd0bYQ2irXBVwh8dK
7RN03/c9fRWBue++6QvsfKyxC5P2/SQmQAiAaj9zBkaM7NbOw1dFeSxsiSn3
LUY3hgIVAGwArt6ewYWf8RVPv/VZgJY6JEE+AibHByxBxCPWQa06XgGg8NxZ
lyfvaJj3Hm6F4XwO0BVBRrknDTdJyZhI1BQrt7euZDHiBlcg0GeAOLXCQwGC
tcHAZAREILriQ5lhPRBcF6srZhk77DjiU692rsEXbm1A8Kvm47y1Y0XbkcJG
s8bKoqPPzkmXUi5p6jAt32CsD+IGiymYm/o9bAxFulq9up6XPpv/A41fkDT1
9QXfQbO+cPvK6N3wp+QtMOtOotqX4F+icqsjC99FKq3rnhBITrpmw7pN3/EK
+OB+cH/eeL471MQSpUoWJzUm6of44q07XcCnauyeiJP0zmXCgX2Y0B0i8oRp
CnjCtEgLCSGyuRttkTjNSwIreaq/6k/AdDFS48s3adsHK9ZD0/q52TXYE0ds
XLX5bxAvmkwjPjitnTcb1zwCMM81/PNY+d1y442Jbu+rKD8dXyWVAoMx+265
JNDECZeAebClG+ayb6Xa16z2nfpv90/IivAt9xb0pfU9NcUmXhzwrxyjvUZr
Tu9wcLFhAp+HnWaK0LlBXXgjAB6rD7wIPUBC2+acLmnFyi2LXdol9aWtvTwz
RTA39pAqB+0YRaA3v+J796PbrAYakFyumWKQCN7AvVTA0bJTMycSDzKaDhOD
hH35UKzmRosVBgLsLCOth2RWXnj6PLccyxi4Em3/yLwDDRUTBdfBurewdAsH
0hWl8L0ICzSS6y0vVJj/Mm167a+Pg0CBFeL1R2kIrJz/6AJKwYCjo3I3IYFW
SfxNYzJgauJ1u5yKNvt62XCthiHydX+tDantpHOoSjNjwOmuNySYt/iCj6sh
w6Kq2stK5VwLrWnrlQSCJ7eFaBarwbK2LMX+PdJP1j9i4HU2g+Jp7gERZptb
17YOZAAlEsyANb5VZnt8lPVz+8uKrs8INzEqcnk47aTC4lORPw70guqJPozf
c00V54pp/8KP39ZSgYr6t851cyarvXNIiBA/ZkBx9Tg4Ws8yfvZ1+63cSkpe
2Ptn82go1oaIIawCFqYiBiXSa7CeZqSYxYzkdKOdJBdokpx6Tn4CYijI+inR
1+p1qsb6l7XsTP0afL01jAV92Cg84hJDfCUnX6CIEnsERR/IbFwcLRnlii5s
XRxbfAc5+NxAsTaJ1Mf6PW4Rwz5iKKn4+2mH+r6NpN9RtSV7LkI4l8vM55L8
HM6dX/wV+yF9l1AJ9MM0kNE5wkwW+nleqhId9KrOcFANt1qT86Lc6DLooTrJ
nxkeyn5gnZuUAeVpO/hkxDE/CYTHJYHQQM+2nSmSUPs2A5XgN4KihWdV3pJz
+sXwrp9psG7QU1Xm4bARx+i5oQax0U8ws66PNnk1bCPwLMZ5kC14EYcWrYRV
N9FwZkjT8qj/+CI671k1Yu7vnVOBBY8Kf5EqPQ4y6WCrPPp/ovCRRCYY6JP2
RUXvR/8IKRWVrOFZlCcvSloiYKdLSVCbpRPhdFxIF12gz3embsR+0BMTsizg
n1yDYKKDDN8f19beHgiT5JkfWhV6y2+oc7tsQCT55FqA3A56OViH3sWBMyVW
JvjiNP2+/GS6nRs0/ZJ5uOzqRY1ZN33jEi5gd+ZzIPlFPTtNWI3fEPO9kvGo
Fa5JD5Y9vMuZy25xPXUc4koicDUD8DAKxmnj3LKXblwDEGothJmEbXUtI2f7
OI/70i/J5HN1OWsInEJ4mX00kfvXJkldXniuoTlzxyYKSKTbZ97U8rnWaGBJ
dY3tcVhv8VCOFLQoqhDP2KXtJhtOjhySaNsAdoN2/isKElHUGq3HOmrGrLJ7
S1mAuyPVnurOYO+doqXPSVB/0ZzMztWcHTPnjEuKzqDOuW36onDYd2gQuDuF
DpIJ/n56OwbhJQdn1FTJ6DToTTxTHYZZyziLT5XU+FYBvRqpj9M+CRpRiO06
sHViFaw6gPB3dxhAmqih5VIpvgeancG3dK/sxvNIv2sJZ+CNDD6vDm1mafbT
QmLC/958iRtPPA2SK9ppKl3beSjqpdihBXF+aL/58ehPtX/zVIFYmYHqF1ww
/+ohKH3a5PgbRj22sALSVHse6r9zJhYmf5loAMrBtalJ9kyQ1NP+wylSLLI7
9sA1bJdYbs00MGf9oOHrN2fv2+z52dO+Zfan0YxHuqq7rQXUSHTmcu07ZlCz
STi/tOeToGyMnF975Ryh4wm6S70a9JQRYFnud74DHjvjzuVkcnroJnUJphYH
W6FOBJ7d/MFSEN5dQUTkejd/s/Yx4Lr3hhZpHbYl48dpKQQPTsVF5x92DC2c
/MEaA9dtar4J+ydmar5MV7da6TXGq1Tbz3t93kn1F9ya9JQZdHTvkoydK2SM
YIGwScRT+rZXElus4HRhIZmznIYSDIyrFA8nWetDc1L8WRUBB+CfZdCx/r6h
2l6XB4vOJoNPu278gyX6tf4TnFhw94T/rA028sHk4E3h6Ob03sM3+NlzYPxF
mr79pY5tqAjSN/fnwUoXjWpxIdf6BPWHI3C2s2CbjuOnjF2ytkNgXJtOTm0/
ohXm1uRFLYRdeWzj/Rh4nTYTLTub1Nnpo80VoSS/d5xcn9q4uEwzoQ7FZPBn
HflwsIvwpFpFoK0gxyvzfOebfLQ9WDdVTNtfx380prb3TqjObR1XmeVIxFpH
KQwR6FGNbaObpKjWVUp0qn2zZ3sQ5fqHY/mFCXYm0FMWwyv1c/AYVWnzaNaS
VwaCI124rDCAxH6yw6mUQe48kSiJJcuVA5UWFZEMQoGAn9GfFmIZlotEGsWU
2Us4k1ybs/dT5ADbw1u28G5RcLF8WfOaXva203z5ppHDAbPVEhxgJvYDuOT9
iylWuuxP6XpEEM63o941MQlfJD8HBqXjMkng11PrvVaGFWlEddTW62oR8kqU
3BAXev9VbxCgJAOnisRrZ4tfPMihImJUjCPjzBZ7qopA/YRAMzkrrbahGCNl
XZ4alkgyOiNbhVPusetQJWiACA7OztwwrvJF0gBJ6bP0Tpivot1inh6OpJ9o
eLUklr1TwUoP3AZSoNLp1eXbuDHRHwWyV8mI94ZGbeb89wYv/UA7HldRgdJb
zIgiwE7hbEDiFH6rrAFC/WtcrbpJIGEZKDSi4e0zcPePRPF/zFmCa8MGqZ1E
vZ51MEC1AoaZbFkE7wbBwbkDx/JeAsm51UzGFO4rezRWQUP6yuDqZp0zcBcr
Y/90yFZc26zpz7j6cCxEpybj8kb05TmxGou5qrZ822XHnXfyNc00vhMNVUo2
Q5kLM/VZaKpMYylV+oOHdSwnMoXaXRAyDxgj83viwGfnWc2/Z0GkKjqDTje6
Pc9cTUWPcinM4et+j1KJla67OYCHyA0P+pieX5NpKbrF2HO01/9HhOj07S/2
75JJmGHsp+fQkVSyyxCBjntO44KvlGYqI9xLq55KLKoZZVMD0b0wtZw3vi+Y
mGt1HW81MwxXyKLx+y6BSik5K/Nx2miBs931VcMjv+upfs5S7ezOQoEJdmU3
XDm7/YyndTx5nUlVoWsAQ3mh/NhYGlUHvKJCcaGaC7ad4SBK2zhfrgIvxetj
dNbS0Qbd+FDFzPFttwI7w6LuiBiI0b2A+LBCuXYU9h46IlHiSZ/p3p5Q70M3
WM3AN8OyKcL//T9E6ZW0HOUXidWTCtUlgI2PTRdNrYDKiywmufGvhalGb66m
9DjVMdMNo1Djh/oDrpuZo72nZeDVRuOxg6xYadXMv3dBoZ5W0k444qmsU77M
ymGAr+Z0vXdOaujW+KACD0UQ0Zys5ucMHwQfGkxFdseRNK/SeDFUhNWN7K1Z
BcoYv7/UlhynrSe+kVYbqDXW51VaKiP9kI8CwZ0yceYC5nI03Z9BTo5TQTxl
XcQ8YuGZvODNps6rdtOujpc7lwYj9azYi/jAhrvzmbZjBNpTE4uBNQKckoOS
TyztRpYv8STLijPhFVak5291dfmAqMzG8q3ofgBViyWHAh7LKbFBT5KCNpHP
eqlFovwRq6IlzVlK5Hs5Frh54KsA310qDEkTT7s96WuAKsJg5F2EcBaOVdWT
QCUm0DfQ5TQA8rSSvv5zGyMMQJNQKKCKfZ+5yat0s7ZFx2S5Fbni3mX8KiUE
iBp+ESn9PdWavQkENVjSN1e6Bo5TRnUDfvjaV5ZthAJcP4RdElVbz7is7Jup
5RRAv7IMQFkxD9h5v96W0SfusB7C3456LCm7nmd4zweyTKZci3ru9XJgOAtH
D55ko73MX4jTAZ0RDRwAkKxVIQrXuSdS+ZInxb1qvK3zdwIMvvrEcrUpZTjn
ymrzepw+L21B9IKIW2VCEcg3sLfEjpto2M4i8g22ThY8yEofvFvV47bHEDwX
J0wVfac2MjBpX7tRNgqbUz46sci0+dKpVBT54FZJIzt28KDWKd0pcQzo6ADN
1RY05wDXys9ePwUT4wu0JqIJGwegxtwbV8ieEwdDFVQn2tFByqxRyP5g5oxr
salrgMRtSWgAp0GYYHxoE+9BOE/Q8O1nUGldelKKtVjBGfKhv2aErXLZHLnW
yqZR4PcbpX4EQF+ZqDBAE+Q1Kdac1pTDwLwAH9+m2Icnjv4FRc8VDiKlQf51
0h4zLnd3BKvPR3O9Fec0k6inTt+Pz51rmAffEudeJsHlvNE0D5oURGOxQDBc
PVQVjlWxDstUAWEgTpFohQFMkL4F/eD6rDdNKHgR2nrgECGa41P//vzW9F/z
rSzgjjJ4xQ+zl75QtZx0g3yg3zgl9WDK5+4TtGjjkqtkGpWUKLvEBVSar1K3
7doKbxlk0465fD0rfb4MflwA2dP5KnnzxrmxG8Fq851znHFQwh6yAY/5Uykl
IS+ItYUenfsmatTs92Juwn5N040nUCdBxrFFizMae6eBdqlZDx7C2aIs9lOZ
RpPXsUS5EU6u49Udn81MnYD6RUKDDu6FhaGSBacNewgbMHxQI4T5S9zZF9L1
06Sb8NFpnvnND4v2F37F6Nvn+WkK4KaA0kkO3YrHV0t4OByaLN+XqUFc1in0
Rl1FV+7RVEeK4BpfKJ4NLYsQybbJhDTo14BB70yjreC2dDJVrgdV2pK85mhW
a2ZprBSV7iCbzVPe6Lai9CD7ShyYCNaHauCsgzAKgpopftRnAGCVpGeQlgtU
MRbssxi21tdqxNgKt/HNOFlA6HIdivNej00sHv83xZwsRs35khE75DuuMR+2
mY1kAypClclgKXBvsSGS2oM3CJrIz7HrwjTAG+VpQBfXKIy/GesZ59UudTTP
ic5DfZ9//fxmjJy63+wgFWuPFpy3vnV093DqEmdppO7Fe2mrlNwzrgSFgGMJ
tZo091AbeNbpmel6RZax8sQ25cq7IK5Ued8OcnSw9quO50yG8jUGnGzR/GZ7
o6YXVxmRtQoDpaE1fydoqOEMRY32+52qhRG9eVlNs7pKIKEpX0EkNlr1C02V
+FL/tzk+st6KqX7L2FLQIGpDcI+1fLDIX4Q5cBZaz2DS5IYjvbfuq7Z6ZDmi
NWd74cGu9YHFpRiJF5qLIkSMXS6XgmIECoLGPT2/ETlM5Fd7vaPVzEReShZM
DjqblS9+Hx0pOyuO1SAcOKaO907s+pEn+q2e71fMOkZvNgESW695dyWW69aY
armj6EN1xdPRWZxlUfow3WrdqDSKZ0UePwRW7mjmnrQ3vVZgntrX53x4TJJ1
2KMdbgfgMn29a7rTWk2g+5Ij0GpmcADyZo9/DgZSYg5+iXB1Vcv1ccs9X+ZV
w8UGMpyW8iftc1gIi6/8jyAem6c8YHUjZRaY96u/Eis7OI6dlOKzN+qEhH2H
+kIO/AC/w+48hCG7XuEw0d1wKnjCB96tqaUNOaRIsohDGuiNQVVkfOzuHLCH
FB2A7ITvM84PsooOvsY0d5he88qRBASCZJD2hs1BFTUSu9noI/n8ZIq/9yFA
a9trXTy75i8TxBg7vxvKzrRNjTUwiHFrSKkBG5i13UimurOD5Hq3iHPMvjSH
TrO0INX/Dt5wlnEHCDfXHIKBEbVQGEpxujRY5GZ2ijsgx8MbnJWdqvHp0AFX
nRwpPHXnSEGheqsSjkiTn9UbUMCzUvsHhBnKB4JGWjyhftEhnBBfJWEpZbv4
TtnHK+v9p85wgEVn0QfwSIC+c+sszazb52S5gfqcwbo+2U0T7cTOJ8glvO1Q
TJ+asa1pg0APwZHnMN5o6Vr+m8oLcKuXwCMyGFy1yNH1N0CNClvjCAkzNBAc
eMts727CYqnCZEy6EBj4Z/wOkhceRvm6jeigQD18V3xPmd27ay0r/zNeNuId
W50+rBms+yMxDnEAUzNU/t8R9YINj7fCGwUpQxz96z15Wb/wUkwdFPxzgCKj
jsxbp9VlzqUL38hc5KcWjLcPHVIwMi6oZPrEdKZSYDG2S0jpHg3ciGs1SJTS
g2DFTtGNdhW7DmO2yIYcQdjSZmWDlMW9PxWfHaBKqSSofMl9dqCxfg81RVIb
ykWjW3jHFP6/YIvj9S6kz5iPheLZaLlfmskSal3BUgEwwWruy+ivzsdZVdxG
fy9Wgl0QKnN9lAR6ufeNy1ZOkiIGrQZ2kS+ejB8T8hpRDzxro3XqxOXTK7w7
AOCZenrgvqnmYmCpPQQ6JEsK2IS8L3zy4weZTFn52RqkoTtVnumTTjpctlYE
SvNotGNcQswLV5Hv2W/9mEv/hx6sOCEPP/YOoBtN8nElonwX6knm73K2kqSU
B7Hc6Qw7IqfWS94qsip+gw2dYJtD7EygYGYfJZllSAZPLQNodhS0nxnX9Rwv
xxbF1o3KlKB0Li/yOVmyzavxacYw/r2UWdBQwBEE+PWoeXZxFF3M0zkHNmrl
IQBiuE53dPBKQn+eaT+H8W0cMnuNgxeru37kyDyCF7TaBLEyv9TTdH7cPsrR
bOYYY5XNYpEFUTsVSwEMk4NvFeaTGj0VJrMr9wEvEtu/njFbXvrzAUcb+S9A
DoGkwauxWwNtDD2xulnmab70LLgBl9DuSLrG399L5QWGABh9JzWFC4hT+4fD
3gQYv/mwBD6dIFph/BBaVmaIAiyil0BFbA3EZUoprEHDlWyoYOnTS2P7AA2C
ltDO2AbnF2CpH6PvdjEfN1IK3Fzpv9OhQuQFalu0RFvBHHeCpPfVTK8bDVAY
asw9P7npZMO4WxqVyL60GfW9IPZNiaag7qzKWwo0nT8LahCSOlifGvdLGOw4
i9twkJcq/fdXaLFYmr+TIItUhRqqx4vTqA6KQAL8yxzE0Fu/I1lg53JMl0Kf
F3gsGCWYIgroKKTCrcaxHFMzYewUTm4tZO/BJlMgNbvG2qG7+4s0zB+xsrWF
jCe484chaMCrQakgr1tSj4Rf00KSEZe1J6fpdoTZqU0ocAMgWBQmmuBKmhZj
1SZpIpqVwq89slT1HE02LAoUs0I2681OKHq+A2eVzx4BolLtNuVpODCjMBgx
oABO8LbLoe60pStAax1/++9kWAU74DB7QA87vMbzQwW0Vh/04X0QeDZ/UASU
hVsUBNTtZ8DjhTTDJUkd9UOzlEyIC8lIF4UYP+N+7WStmX1otny7iaGZNAmN
3kQ1bslj45hcWiawC99o/ZP71KT6BQBP1Qrz0mW16Sn7BvczEcdzVSDdtist
Q1r6WRvuGYHlGy+wzPOS+1uWlGkFVxcMCVJYi24Bf/W5QXabRfBsyXnHNWiE
zdN6HJ4YjRZnK4Mi9LSc8dmwNHd3H7o7ESfBBx8db2kJaWLIhK6eghEmpsmd
LEpPuhIHMKt/SgvPJ/yRvnkWgS08tZhVTNosgetOtMV39kJnZrz3wT7nrYL7
tBWyh3fPqdtlVIPmRvJ58nIuXoAXfmBNyf5kWOnepZ0c+9ICLsGvULGES3Sy
ycCM4sOGNpMJU6BmO1Tek7cLJt90HWWssN1GTqgWGrpBCvZmYAkfupJJTltC
a5sh90EUQDC5LWBUrbkcxmiZWs/wwl0/kpGOIX4mfr6pcAt6pcBdTREzwCxg
IDBTcUj3fBGFWkbWaRf1i0qLKDknVkoeMH25zOUZJTAUky6rnwfGrIExDY5d
iRl5XuitOps6Hwg1FIKAKfsD3TAChOF0USR44Ef+dldXB5HAhS6ARJUJvFKe
alOHFRQUlS6WxNMlln/BVBVyTay1qa4EGcMy84rZLA5eoX3iQMaBuRs6dusu
9ruH7DIM2PN/pB9HZ1cK2bFt4Olcc77qJrHnzK68QtyHwndzySugB4C7PXgp
bbc8dp+3D2wOEKH31jpfCYy1EyDCcWitrXbC3A78J+xPC51Sx15+hiChuRY6
V3GR3g40EIk1tPIMn1Dtj+kPhBq97XzV2K/5siQN2l+A4w3wLKey+k1ljZgk
G92MwLADjO3rk08NZfos5oLHY4rI6BK7Ay2zIjeix1tH1Vt9Ds21ZAM4ubEt
inqu0DcetJlPqdFQwJaG2ddKt4SvoRSZMuuhejU3OF/PgVLuOw+9/+v8aVZA
61hIg54O6diEkLDvwXcuFxutqVQk3QHCAcn7p44sGh9PthYbg4O5qxa3zfb0
75mhWnL1+O313+E5dPohnwJNCZOkrX1yGD5rM9+lNmY3NtaEr5eHIz1p9JS/
UXYJPxScBCj6c3NiPfwymJOYhwwxOdYuDo3jKx9CSTUG0cZXgmxRfaL/vcdC
PfKvsi6skP1jt8ed6hgEBSsIUKauCBnvvLa12kgofu3jSQoXzL1SCgvUYLH6
V0IoyQRq6trDjLHjEVa0vnk7zjecvnAlH8QwX6t0uzflvzSAemKStVlwdKA0
S7/D804OJ+yBYmMzRvSzvOZpMUy8XB8hH6AihUuJElALD0s1TVUyY70auMtC
EfsXMYA0H9RB0aGaYNLqHDd+ADMXdbRQY7MPVVmig+elN+ZfnlfHBTx+ixnh
6YOxK4NLy1KTQwse+8pRSeFcuHuJqmccrdR1JbRqDXCWjQOsQCxES4XUIFjm
XUOYww+ZNETe4WHzidj/zjLKsc0+FI9FBUaB3yZKcEFCf+xCavaXWSw+RYts
E/cSxHMNSSqnkApguWQQJ30mJ5rVMhr+M1McpBGa4Ni8ktswieCm5oda8dz3
oQw3x9ApmtGrJwKEhdpuvhSCxKf5+AqzQk2oYR5K0JmZKjxxMHLaflV2qU4c
jQ/isLBL1By258kBbhv03mDSZdyiKPPP8EsuEfx2/6L5CrpzBpFWb29FlXf8
S3UGA1RY1GAGB9/PkMTEwWb/gvgpxIFpiA9c+102Rm/2COcrD0vBFQygk083
qi69hoOoGoWh14GsiStsGWTZo1yWxynb2+dLxe7b7IMDKSwUxbfSKtS/XK1N
EyKamn1FdqtNHdWEiEcC58+O8/SshViHplzgF6PskTeJwnyuX4kyKo4J65vk
58vaAzoBTxDhv697+U+nOpd+i6cLF1+WJ6cu8I+CKi0ByqnkWUCP0upcMZyP
wYC7HlLg7dkRtJLLsV5x6fu/fAs1ebXrcIiOJq1xnKUCMCESZM/lORf1ctIY
2Y1bUeheZ/6fri4XtKAEexccOgLYIj0l5p1V/W4t9rIPh8VKw4Pf8AO4nkPs
SKnt7nO2yOR1SPW8T68wOFU9RsBxB2O/8l8SzAMGXpxiKPYgOtZBsB3Kw9Lm
JwMldgpUUuJIH1qOsxN5/QaUOlWYZ97wMPG/EMnSJxe+9XwhYfzPbdkAWrPy
sNlLCka2b64Sh+g+3VNvPVc4sgl58G89KfrzIc1VG3DPd1vzlfnNdJ55Rxbw
pPhXlHuueF4oqC3WMjLhoboyIr5JlSffNYcm+o5YR3zgIUUvsJZPhdrAGU7Q
fTwE0RZhti3MYOzjZXcCAvp790Ymkx7/3FHrVr08v1Yq2Gxfy18WqArMySGw
xJVWNuN+gGoLt4lHbzZ89It0L0CPrjbOUIMrUMafYjHiaI1sPTGlEmlM83fI
i3CfXTRwyr6YEQOoRiNWcCNQ615uNvfIXjBi4Hfj8OHmXb9Ut+nuxhmBRWXi
xK0Oi16i4MDZHIeD58EOHTLq6J6wBt0M2+ToVYvo7Etc+c2ZN5xO94qtcG8C
7fFroHp8/0wF2cUcQzWH7UniyRVOf+szP969jcwyZQbWhg957+wHOIc3MbwP
B0JgvasN7xXR2808jFoBQB5pyGQ3+4oOpzk08gOt38T6uFwjH/STwfRQf+h7
1o6IzfUlKKEqe2VK6eCyACkbnuf/F7sLjkZaHURfXcNtXRXq99pIPQkZPSJF
M403cYSZmjiSdXhNs6FY/piv83F268Y3561MjlnivrAEUZe0l6yLh/wINlRp
p1OxF1BlB6Pa4X+3AZ9plIhJgjcjCrVRrRZqFP2ziFtSkY+BHaTD0cuYOY6z
1Rf6yTsZikBCM8O32Q7Nm5uxUI0bYsyNbmw6CvXAwmJ1br/ph1TNbxIUwSmF
PiC5a+vxOf+nHB6WZLPUBxtTT1KWTpst1I7gBWKyzdYec3bHZd15ztNUmSll
7BQ5dCnRfvKqhrdRr5mxSfQwSccqov03CmufmCyJUk6TbmYhoMBy3LHp21gK
+48tQjnsjJCnY3htDpHZiLJlyEFpyyPRMpwyOftZ4N1PsC8ZsEUSimYt6n80
pJsIcL1xc8HkKZ0DbjF0oOboyXpnvu0kNTf2+/V94zaD4qL4sVYJ3vvvuokS
rOds/MhThIb1A7mINvG4AUEsfqIYw2xabGjr7tJGQpogv+IE2DzTYjWZltIu
y2I6ghJKQTnzxDE1H48Hnscz7aEdZOjlboAfjeaHiRfAEwTRW/px3VMm4nmR
BxMWgcvG0ibbWZHAj0QZx9vJzblRkuxz1gEqNlSrKrm6GVaDWAeyQkrZGFZ1
kkhykzjT+mQ3YNGbU6kazMHoLrhdDrHlFUjcm6rf5r/Twa7bdz8aupki1y/c
1Vcq+qCFTzjXm4QBazglvLKk1AcmAyQbUG2judP/PQgGtfRVXcg/0PG/8W5/
cJL/orLwsoLLYeOT6dhUj4F7xKyOVCVVQbnqSynFpVlgVGD48nkq/XHotdto
2w1C5BTb0s1Ox0HPfw4WuJOxAxmAxk4eKLvSwPjn2X9/AMA+giJvmu3xoRta
ztL1jO8iz6r/uKeN7wHLMlEMd6du2LW3PgPp1JITuZzJ3nOJXeWlQUmpKEru
98C+kG8FL1Z40fGhal0Y2A6tnHrABVcNOkW9o5WPS6HODhhiQ3RkjSkAE9Gs
B0BHVaQvq/LXQxix3LaO9YTgNMzFwPEHpABXs5Mry5wZ8K5x72vxl8Wm0JnB
LkdFmdH7ggQ4ngAceiktyQB1tvQb4vppeNcmRkT6vmRJAV6VkJctiwr8Yh1Z
4LKCKen4VPaohlFXea265TWJeQOFaE3Cw2uQ/3xwJkkuVYxQC+wl5YNjglM2
8LsT1vDh9gW5GcXqgcw9MuCd3iBDCdhy8ebEHcuJGv6UYetq7WMSzFKgNAfz
7Vo0JGlocaR0HPKG8NokFWtKGKYBR5TlsaSiIGlx8LOaAvT2CFF9D4V6TZOk
EI4+1SMUv2FFnyykIi+N0hL19iQjZgBc0TCx/eKyJccMktCmX+7efYMiQJv5
Ua+8kHFJhCHEinmJDmrDDCcQOIHDR5hD4xxDr6MSlTKVGz4HB6HMLG2sEIJE
haSwosMBvPT+/EMJwhtXox8OhQnyQpO9tYF09j+ehD82o0nXrJ2hWNOIEDw0
h1grVujQzkpZRqd6P5IDeMXG3QT71S9Wvt1wbJNDV0YCFa9599HzZ0I2NbRj
GBw28azluMjok9J0r5DUqvmjnNfLkU+pIyoNj8oHFJ+5MgqxpqovsWl4XZI3
+kK395SG4limNQFlNaySumZ2bqbBwkMn0kCJ1hbROCUEgoT5Xf3xkudiY94V
nc8wYgc7xeshRlTEkAR4qjOE9erizF6lgrwF+r8QUAWgh8il4hHD4nZsmYQI
yrn38ilYUwM2kX2gL8tuYB975AHZ6ToUaUovVd8GJGUIo8WxwG+7u9NYGjyE
bum9+dkTqdvstqRSJJbt/waPZfn0igqXzTGCbZPHCR5cWhARrPaBVWhCPxYV
UIo0KsrUAtdLFn6cCnXclhiqucBkBftmjGTfnptFV7tbgijdAzchZK+9ZOm6
lDlrm0CSkuwHJIl3x04pwC3vCS7RIm0ZjhjdS2yWC+WRf+ALZJeYJaMpqr4u
S4cULYTFEj89LT1wA5q0/Zn8xrhNYnypisiflXVjjy45rrlS5btohRnrUQVa
3Q3s1rm9pd0cYVBCJCjWVLdokiO9IP29P9ZQU8LDK6lSAErDRjBNU/qK2pPO
1sVU05ZSGfDrw6ZTHz2V999rIYfgoAwgYAt9Ixgs4kuh56H6VC64aEIzUqbh
3bGJ2HX59kEa2eET3f+D+euJhoabRaNn9Ge/n805XuUNpWZt7TU6LGsG6DGk
pC8Kp/K7vOxOMo1Lim4vL5lXeHwIswcM3aqkfx39qz0S2AIpZKroufw43/4W
nWGRTm5Zlun+O+mbqtwtRhID8+g5wj64VGkl2cxnEtBfoJ2eUaX++KLU67LI
x1hrdgFxF4VxwzaWSdKTVDbHzoBWz0TcWsCsxVWKEQXqKj0NpRSGxaky99pU
OygcqhkMZauBPUy+PZvLrj3bImHhQlrVqidN3cl9/TqftejWrIuLk82h9wY1
sTu0E/6cyLuNzrhftaQsE5EL0/xvwowF2TFux/5w6EXHbFuVy0ewUluz45RS
g434mowx1++qO8lQP6PsjYYI3CJz2Zj/UklbCQKWockYR/TVEriYbWCLrB34
Sm89W8+6H2kSVPQnQUi0LdhfRhN48fwgmkfHqpLnGyEOeMxZtA5nuj56dVlc
0L1sVq+vNK/in7LY4C96Dy6/7y4/n3fi+Am/eNozjeawkoFEArEW2oacQQ7y
nBYGaxW6wpKp/JLqunfakUp9w/k70EBOvEv2F8p+gRiVrtaPf/mayjy8aKgg
9ufR20MroIXuYkXivD30MGHMh/i4YYOcUT83ECGSrj7dM090TIVRQRoqCxCU
+WT5qqGNl7I/Ie0otA0YfDFiyPw+b23IWL7REfpaYLX2zCoOBxi7x31ZK751
lleCUSTsqkRap9Ln/XW+JkCChfg8YRRhLwgXLWQgCzIje7G7CZ1Zj2T5Z1sI
kCFPGwG2LdJ2PqKn8VAfynNsb7HnI1GfxxFecg955BuX7Suln+/x24ncKGTF
qSumHsKRcZv1htPAirXs+vx6rfbq+VeDxVDn+TYM3dxRWZbJwHBSTaW9EiP+
diP617U3aOxoKXuPmvMRpyT/sAgl9V78sIvb34BWj7gb+ICDokdyLVtN0J9p
+M1l7b+De/LqCq1PjbNbGQDEBaSnGGDqdP+DqnDN9n8/8S6bLJaez8ddKPTT
WM0jWyx0KmgzYirmjVFq+CqtD7Wzi+dn4/eYN/5Y/IZHCOwXW7EbNk/S06l+
r+EXfCAIeZ2s4r4YtD2t7uA4xy+2JTCAyq9wTWWXZrXdNSEvQPzD/fqqhR0n
asVgMZWfhZtAc9EtIuxLMwI7vm2tOtHz0a3Ds0ov0XJLH2vN+8BzbtxlNrTC
7cfPE/XHDE6yX6vf5zM3OoMRByB6lpEN3uThtt5Skx8p5LDM4qfJYV3Jx6xb
dx+wW25whYtGA5S/9S6zupDIFL0uMudKtBgb8M7X0YS5rdEZXzPx9BxaxRSb
HCjfeok1Q0OlzE97N63OsL8w58yymJLK+VAtAhEgfayxLyzAgoHyRHaUs3d0
JqjZNTk6p91OmqwkXCgXdJP8MnLgdf4M2LUqUtZolxKLTdgMMwXG4J7oxuy4
e4sYWEqNOo/gA1uyexRNm1cQYGhagsAxgMcROuqjmb5ZmwmNJRrS9O/o49Cr
FDteh1OnPxlhu0SO9OXoABrLF2CuFaQgbXMqH9B2y7qEGVBIPTPuUsW7c3yS
heGLu8/JpaV6U9i+RVCSpxjMNlbUIR637rMk/aGLNs+9hVRGZFMUVDGsYWq7
TNs20VYieJHU1XH4ItQysEBKVVih+7fm7qq9b6NInloUMaghchvgrQOJ5iT/
iPnG8Ne5X/q9vWsOU+d394Hj7rRWwXoEpwEN02Y+L+S+LCi4nSn0pSXjfc4w
BS1KRrVx+ufueZaiTdv7Ab56Ls111D8G1BMQXL8mpFeq1lRnV+8d2kmoGK34
Om4e30uxGKwYJxZ2iRkSfdq2lGIO9glafrFx2fZ4rm6quUb/Vn60ofmyzYj7
r5jGaAQTIHdT2LrqyiksWZbAGghKyHQeWrePPyBIZEgyQgBwhSqokQM26pia
juCZrZmbb2MhiODP6TuffHX9JZ4pg7Tl0lEIQ4NM9/Km8vU3vVZ/ONSj82OX
8new1tWFHKVckouM0xb0MuGdeopPrna9U3kINNX9OHq1/UOxpsiVBzKJrnFq
hnSUvVUEuqUmpO/gzk+PN/Zk7j6pNems/1YljQUbuJKAfEpSb3lqsg/Ujcpz
BUI/78Nzqvb+PQO4dgGgK9UJPDiZD7ghwVumbxvnxQdLCImhxykaAnBDG1px
b+y4ijs9cnh2DNW4IQMLp+Ug9Zp1GEIWXR2TOvPYZ6tWtt0Nfyz5Zgj16n40
nfz/DzjR2WPYI+B0UlVslYEXJ1Z82U1+It30wBcVKg7bYaErcrFxIVYKC27I
pkdTWzJT3aEDB1sGjNgvDJ+zBw6ro3qB5r7b/vQB5aVGumXbD40zAyBhNalx
CUEHdRvTfPCBMuGPru2oRRxBj1f4QvToGM82OUjhL7wtmQcCHjnjoDyZ+PCo
2rCGNigQbpvAG7iAQyGSFdn7KK/lC+EuXIvBin9x6ojHrGtc3ZJVoChdBr0A
P+4Ks1kkrxppoNUlEF5/uc32QycbllNIrk69dvTJNTkqJ+NLXonFV22MqMOs
MhW60t1MwUZMb8z54wJEAk46Zm3iPLSKPsO0fAeQHQJ4Eu4kHNkUGvzTAJ1R
lyPm7+wWiOmC5ZMnHUS+kz1jMm/bvua2EDKsd4rlR/PLsoKc2YERUQXogyG5
y7IeNd0JKQZzew0IHUmCYf2q9JJ34xcVIZqRituuU3RRDX/GratYnENpXk69
Qex1iiKZbGsUGOfWdH7I0PyOaqMh/KH+VCf5G57NS+Mu4A2fM1f4ysEb2J+5
tSL3lkl3A8bnEC3c2+bix4HfB917JzUGjX67KXhuOMPm9o5ZW2mL2F5Qtv+t
96lXHYSz73eDfFVTCqxhOgkGtD3+D3BRVwEyK0sSeEkOCXgE0Y6ZVvz+odtY
BE4N7CuoGzPV2v/YUuA9rRS7FmIexdvF6buNI+wAKG/rZfy6IwtfpbQDeqpI
2sxnCLauknP0AgZt2m938c7ueCM7/spzbGqUAqXsSLa0v9viVHvGGvVJtEp/
7tRb4tSwaS2KTpJQI0ltAty2xFXvlJK5z6aTRYy+IrLIyz78b3sXNR2f/cBd
z1w6dJTP/bCRfFjW04W23sDYJw/1VV6avCuLhGpKsvSAZ771s7bTMUddf3KS
rAmksSjI1+Kl0fm3xttfDz08Tovb1UN/CvS/THr6FkdomKQuVqul1vZ7mCjJ
l0a1JbjI8ekK58vd0Jwh6s1cWOsXeZfDysRUa/pJ2iDiWW9WKyHA8q/2Ner6
xOfVFrkJurfxGnSDyRDfM/Z2bjJ6c5ad4A+wvONQEtD2RdrfbU+rIfheWWus
6qWMVtbOortmOwv+CT4p0b84ZYSGJY701vfHdw/5SzQDPtCSjonyjvrYBEVq
zpfXv+InKKN7U54jNFNAgASaBhRyRj4n6hXZJPmse/o06EGRCVcq6NMXshup
6bhg36QcQVeAYo48p4p29M3S0pasihkEjNdY14tuSji3iIr8y4k9GbEkelZn
8KpbaOu6jwB0uJy9uBKBNDnrXGhsnUZVONkylTxDkin/bfLSkPavD1wH7DZl
jp/bCt0aCONIC4goQ9X4O6zDY4IbYv+dYEoSY5uJobQQCbTw1VXGwUKYV8Dm
rWHVAzP6x6X3eg59pQknRJTLZc27dSqv1IU9h95aN9B8YPkMF7YzKT+/YKto
7D2XqFWptPHLgRkDhIDGNEcOwdhmah5k5twILSkmmRgBk6cl3Psw3Bz+mY3A
xsUDSfHriTjg50K21sijKh7nIHOjCUwwMwVwFODHy2r+0JkF+Ern/x1d1PR1
ljSmrqJ6HDLjU6HNMMH1xRDnYcrSqQ2uWVFTRCPHoMkVO5U90JiVuTj1SYRn
cEAFl6pFiXG3tY7w3TSE7tz7u1Kc8YUCOM/SQGKmjewdPdPtZ7C+4q3QQGN/
QNF5hry0rPtNmHcM/Ip3glz6+i4OnPIIgTgjUcE7qxs392xl/DD3apYtYFFw
GD8Rp6oW0aP4T+1ItPteWcYwRZqr5UXDW+83Z4KSSoBpUoFaczw5OlU2SGt8
SueoSSdJaCwF2jDp8c39N75uzlwNH0E2AlIw//n1HuHDUPmQ7FphMS192Awy
SpQpP49ZYKoEfMcToOJQYxxthAyGtIhSXfBV+ZyJVqhC48xccb3+1ZkAJQsQ
SWcWLOhYiifd28QvOC6BS717PbbeILgue1/IPHa7UXrNYlJfqvC3DzpURNl8
GGuyvtU4O0W+C8OTMhY6yZbX3XVpbWYfzegGcH5UvwST3CnnbYKq9MxiAolY
7r3BYwxXCA8HWpwE9p59BaNACmYiQ5pYAwcjJa5n0O429kdgJJJnYpdQ/qs7
UnyHXMH9xfQk+NOCPQqhB0Yb3nan/IP7M0H18GUDJsdaCRD7oCc4Pyn2BAM5
hVWD6rfu9B0H8V9HXZFGIt0LvfP8fZE/HU8P2KCj3eP7nlOj7uEVnhNocZF1
AnU1MSEXcxCACFzSAzyoIZJfuiuA4vD4B3kLhfLSKzBOuX1wjH1UYJrhAelI
Sih5Kr1H2TnPc0aLogObB5EFLBQWQYIjd4WQTcHHEXiJ13infgZRh9PWM2yq
BSXskt1ZqhZHfEbbrSeW8gjD29eGIhihKLvfkmM1XE3m8Gv6qMZAIDYezbk+
Oih+OII+TL9HvyLDrNIWnqVvvKEbp6PEKi9ooNtVRf3FYh+jZB3+g8ZkWHmZ
rq8YC2oo4knKl8lBRL0LQGriEwZ2ouupFA1q8eFHXD+1wKvzb6Ibv/D70MZO
lNAJRoZ3RARRGtJZ6Rnj4L+xXlZMvrjKIQhLZh4XJD8rrYrF0JeCCfuXVk+H
4BX0rqH7Fp83GJkxv6WGOZPf/7Xf3U4fOPIX9KQM98jVKu3mxjEKjlOCe5vd
HIFm7GkrFDkL58CAPcK9lmCBN29V5LkAu+z52cz8xMODBnRl7ayy0EdI0rt2
ItKlbF3iKgTDP2Xh6TgG0L1Bu10/iJ2j/YZNTXzbMN/IvBVM1Zt1EZc3L0jP
feevIFUaQSkA0yUeB3a07lZhopi2o26pWpPfvXZkFllJqUV8jVVIxtqQ+jSJ
5+65NrrrIGXiNgeOnfL5Z0uAjzyPO5h5azaVPcW5kRkbe8heXeV62AtHt91t
4O+HNYxPrdiKEZrNlzLVL30PucSukQSdVjFs5U4BP4+xwM/8Z2qHshj6kuiJ
ZF1gwUwCEuDwf+Z0EUaW8/6BRjaXZuANTuPUNkzys+X+2fkB+UCe2tpgisXb
KPUAoM6PCFeFOAXxredbLiUHqNBadELP/721vUxO6hfV7aBdxDba4+VpXNr6
khkbBlE/g0N7AAjOmFctpIjfhPNjxdvGbk8L2wMGgBzl9qmc/28gWZUhqCzd
MdSaVAbDkE2cJtm92CbgDLJLr5GsLm8IOj2j0TQvR8RDJDEuICZ21nn3m8Vh
NV+6coi2wRl+CghBC7NukIdp8lYIOQaF92KBhuaDCDU5JKR2Qmu3rYMomDTQ
+arM8PeaRWRryXXkdaPlXAN3ZFUErnIcavvNbFOUDoPRcw/cFGI+5IivvQIk
LCLsJ6oRusSHja2NYY+YE47FdyuEvReaDQO9C5frG+F7Oxnhhl4CL0flttmM
kQCWTHJnU0AuxS01YL9uTFOk2rZ5HqufdOI/bFSIKHoeIX9ImmF6tRPmxuAv
Riy55hEENerQ00aHUlvfsNJ3fxJTvmD+SnZOdVn9yTF7VGLf2dWb/hEouABB
Wqcjtc1GOIdA2WfjfEH0t7Vt83tOkkDwaSN8GJ9X/4sQSkWveL77tjHwfOo+
HofBkM21mveHxbp0ibFNg8eVjC/oTYxvDBCQhXkEJ6Xq79w3wfbTbXFjgzfi
UAu9yLZsmNN1HR162302z8Ycf64H3jyzzfwuEMLKdh0I8TogsvWQBm7N5clY
E4eB6gDv2gcVJZjaQjKIG69Ly3GpTMSHae7SasBBsoON0V7CjHHmDWmpESAk
+1gVYD2qlyU+Mm85lB4NaWlAgDz2Ff40qV/8YGWHfng0B+AvF1W4dJQlIi3l
x7q2plFL3d0+r879A7QZgYjrXjRHz8sv0nIbXZbksp+qk99l6WJNuxDHCDK2
w0z7RQAN9SMsdxe38n/jWm82NrLin7K3GuqBKZPBqhHFhr6NA0aB1XiKQDy6
dP4AMmUREVrPVR2+imzF7zSTATvgye+nHeHH67kPvgafiOB7fmey/uloJ8AA
a/n2FF2h/Ef+uZmPEFZtfAVdDZfEA5sM2nPAhooI3iwejt0TNMxtsJx6g4lx
KsWaEve30+QB22hYLl90wz1No9OXTeibH7ps+F2mcUmL1HdepUYfgDsuRIIY
k04pAKF0OZ0/p4lC1Styg/IZEQro7cms0rEQpzH09B6iwlCUPB7sACZugSc3
XZMCDmI2oDLdkpK2dJ0bQO7mRUXNxfNLa6Q85usA7U92vfmKthPDwjyLmLn2
bjU3eqwXfjBJVYeGdsxxm2GD0aDqkJZzC6/khfxNg7rXK+reey10S6yk5crR
o2JFjSbV1KMJQ8VRkcstwlPwsgQkqOGYAfu5NESrQd9h1CPBPUq7C1eZx9nf
rdHT+VraYH/3pNVeeqVMmCYvZt8sZMxTei45YCXUcl0HBlQrMRlPuVKycxfS
m2HBfHPc/J0jvax5/lG+RopwD9bXpS9MejYPZXyHWs7NC5L+sFRmXEnM2fXu
Bs7yDiS2moWZSFXmw5xIMzqUbkEs0EnBo7vKQTw+5UqW21lG9CN0quQU+Nxa
Ua5AN8DZ9u1K22xe1CY6oy3AVWtrP+HnYnRYpN+WdMpDA+z8H5YoKowPwWcY
y8Ma4WsKGolvnlOpN+0qHBqETJgFkaYIE0ZNPgozfIjO4UYZqyKEasvB5nMO
CUt9KvKxPqLqMGRmRr8MedkhcuUJoXvB6iW8yirQAkcI9I12/oIEFd6ODVkC
r/FFLg42B5+6c+HlxHgZRC60rzPSQdz+K5X88ABh5CHvAFyI/LGXx5/Iiu4y
QN1NAXNXrrZ398EnXPWIUUF7SFWDsHLYwLqsbJIsMbOHxaZ5ctH+97urcoBt
T77UE8ZIlp4iW/HCC1VOj9Z/zvKND//RmLMEKuhJaPkE685tGnp8Co4RwB01
I0bgHqZzbBCZrzJKGlgRrLBBNWYCm8Wqcu0I1yMjxguIYEsH4DU5VN9mHEsz
uzLRafV9/JQsSxv7mwUeJAfAAMgNqMHmBnQ0bJ68lDdCqOCZhKgzB6Oxh5p5
K3cgFMV+MuMsgnpa3XuePcheuTuc5FOyFUu+BwT+cdAwEhWvRyMPgExkmAaL
vRf28+NrVsTVT0pk78SHDAYPU4QHQPtQtmMjNjoCw0nFoQNl5tGsZBwDmIwi
U52qn9J5HS6H6/IeJ+MkcHNtAeMhOzmIzXwDBr/65ODCPhqprac5ttwBP9DS
D+uJdeDVde6HvD9dl8rDMSHzpr8JCk1GAHiUC1D+ylbZWec8V8pymNMopCB2
eTh5x3jdeP/FxGEsYZqHR0VKUXFZLvXxoWUd7p//ZyNU45QuQEt6bTTsyWGk
oNYy2MSid5+DHtjH9CKGd1UgaMu0t/eWoLcW2U+xkN788PDVSF1rByXC05rS
PTf2HqqGUW1CQwqw2x7FngPCQo2ci1G4w0WYJYqvZ6jAJtZW3bGGCY91DRLs
k/Xtph5f+CMI2/Ic5dsasrB1nOotqBv2MaIFgcCFUvoMk6yuXFsc2nhIYf8H
wo4VWGCVnw4eqndZH7DH8uextznIuR+D+Ib0/jYTEWLSxAPbVNfHqHX9aGeo
DV6hS1f4iTRP3H1hxnjowSYhJ1joldq0VvtkICCWdxkGwMCCC2mMSgHJyoKO
k1Bi8wDUo7YUlYVxHhCxeMc7OcxQhk0eCnhdvzCCnVNWzaMGhHgvQ4w1a2Nf
qTTMSB1tayqgfIykFbMoqjlSAElB7jjsXSGsRH4l8s3vv6SGd4PKLPHGCs+s
W6mJr6a3OHDDOEQ+PaWm5fudcQVKUJRMRI85Eqt1kD4Z93IdhYXcLpBGP2dI
9YiV1qkNDbaqCubqoEW8BxO9Lnhb/mrBh1HRR7P8dKldP27EVcq5INipAqal
ha6HI91JHVY2x23P6nacq7Fb9na/9CNJpJl2D/Ib6rEVspKrR7OM3DTW6426
qFpJbM5MWZiUfOMjkbqUz0E3yAikR54fOceK1dpTNSuBvxYYtXowulSQ6JNF
Q5AZ+R6PvPxqFsu+lCxJcsDWLz5M1UybJZquJ5nrW+VcTzpEgu94nHiBHjNN
myk8M43khtJjPGiXDDXatS1nVvMspSMFg+qAP7oWiOVDJHciU7JHzTSzyTMI
9RIg0MFKiE8DFAVWRl5+mt27aPoxM73TwHSEG14qPt85cAlOzRYfp94CSbW6
blT5PsOrhz9d2QgkBg5AukRCWqolK+Vtuq7bF2DxOqlibDrgOvAix0i8knRV
wKvMT3b0dZYEU9qeKCEv338ogTmR+7lMvSIvpLuRNOJCxcW4iaefHR1i5xTg
vY+zEr7Yo5LbBUPJ8q9Wx56yL4qXYoDqvHHnjxvFZvnEHXd/7Cuo6gXCTm3r
1CcVzyWjTa6iBA8FATDB9RqGjW9mW8rxo4z5EtqC7RXTo3nGjEy0cQMXAIVE
Lfu4a3wigJNjAcm3iZLAzEo6vm+LmYkcSrihrc2mQsgPOL//8mJQF1mL/DVp
BAGFeDwe/6H/lCsmOOelDcvG+eK2JCcqhCr9wzuwGHbrXA9MzFOX8EdmBco6
mLJ2s2czunVjGTdwYveSp4VYkk5qXArxR2mspB/jMJOjwOBUBYdzSPKyySle
ON8A/qICIkKoWIl3BqGu+Wtm3R5Crd6XlMTu+weFQKrlolxJtGFAHD5MqZx6
lgjRkP2C2nbkwi5WXJCmHbKfPhD8v94ttQKYQX1jFO6rM8+qU0Mu2nLaTImZ
JDocgpEC6X98Ub+Iu1MoWgUsDaTImiLqKVv6cOpzNW4kaKtLPIxV47iZTlCS
H8ouHgf88Z065ernFLJviUg32cmyXPajCd2t+XIwRHfIkG+iaiogtzRZGbxO
65DJ+bUVQyee8VmYgOYML2eQw/nF/eAhYYHV0ATWYd1DgZw6+yGFmWoCONV5
Z+vReBXLy2ovYhawCPVTXsNB1BEOLwSJncA/fHeIILxFDbAzgkD5Dh8DCdeq
E5ZTmXBpDd9b7tvY+Hf0wF/kcnhy5yUT1yKQphUqY+Tv3qtirkeFQEKUNv4B
6+lI30yfS+5dQ4evbr3HQgqpOmKgMsrx+n8vPp8xKfyy2EM2V0v5MUqAPPqz
WUrdGsunKiBnnKF3UfXq8SODMzYuMx/kFmx92KLXiDXuDKtsnC469lCrUUEs
C/3dMQv5wLmRAkJz5dA9pn2fk2fa0CD0L5vmB+62xg4y/f6v+ib68+Q5tP/O
sEiZHhodYzw3gKBOyazH/6/wzPMVM7iWNggMYTSyLdbFt2PvE/e+RY5gKS1i
JchxX9xD4nOCjJ5MubDf1n2qZ8JaNMk60rIhiiteW0A9hJtRKV9cB2xsoj0V
T8yfurQhw42M7RQSFj7u5XazlmUxBd7SmESO8keWV1Q2CEBxJJerHZ91pxi1
JckxSSfGCcCEFvJks7gWuXjoJsOqMF+mW4xmyhQWFq8LxTukKDl6qXXRRLKp
qm3xqFmdenqMybj8wbSXqMCJ3Hc1slT1Ct5M/VhkN/umiHp9EjmsW4Ls+Xed
7OwlcGuJm9NpXC2YRMQz9bRIaGKhMwq6StbB2UrmOko7ffYL8bFWhgHRoZY7
QwjuwKfVl6g0pCHFVAzdX5PfCjZQDQ02/+lBxUXabCkehqj/aOVM9GtBRyCn
Gs4fbhuy83dOzqv6JJZ7ArKOndmr/l53a7ItULLxomhjfzp0b3oMa54O5gsP
SVhuoarJrr06YMlfw5KixWS/NkRhzRywfulfpAEwRzZE9QR6T9dQ8oHGCX5K
Lx0ogIV2z1MomVb1mjMrSuwQs1Ap21S6RROCjPBs3Cz/XEEOwO2HaPlBp6aK
kCv51RpT6yB8R0RvuUnmkuqBo32WNlhEivIsW1+3Nb2BRmqSerTDewHB2CcI
KspdlHgBLlCkYIfY+5KkFIz7Rtv14Y/HAT+FqkheqEYz7TjKnj/m+bdIt8cG
S2dK82To0ygd6pJQWmaHBk5OgVyClwYW5EkPm7f9LIiwaRe4RDemF3mNzg4j
t0/kYz5Apnl/36cqi7yy2gCNm/IjtFihkuW7N7iSP5dnHGzjRUlvV8+8kPz0
lPJTxA07C2nu3uceFUMNFfcpExTumj0p9Yu55SXqvyHuTzeRTNb2EjI795ao
9RgAHyZLSXBcidZW3KW/vHWe8r2JiQeI7IcKbREtZ9LINQhvoB99dltF/E/w
9bHk0Udg2W/zaSQG+jZ6JnGXYtN5GG6xuiwjAaJ5Nh3Ye1rISo8IBK1xJery
Y7Q056019lp+mdVbC5tYXb6YH95V/haw8NSnPbgDLfd6gh7witYjkUgNmZYK
6YcNXLejeW41Q7ql/Jdiuot3vUXCTxaPIJu1v5mwBojoB9LQ32EiXYBZbTis
6j4wooLYvP8LhNUm82fese/RgHdP3ZCoENw3dfvddv6kxUMdCBgmDTZ3XPxh
4WTm2A1xCzr0P/sf8GEIYfaf2raJgDGQK4Rrv+vLtRzUdha4c10VfbNWQ7ef
mJZ+k6jEh5xhJXej8vhccYh6dmfMpx6lxxMT6s2MVETJ6pa5GedjT1c3YBy9
vhXjKxdxXsc5vLwZrenGp/OfyYoyfU2//yX/ks33PASs+CNKRLiA09Xymk2F
BZU5t1fBO30Mpvr6+E42qfgYefdgIfWNAFmuq7Hiqq23Bf5Sssht1N1L1iUN
09z0CiMwhL+woLaPlyDHFujqNUn//p0hkEuQLQoTFtQx3JCtlOnCQ9dGzP65
7UnRz57EvBFTv1UpAOkt7IFKM4Py03jU5XTIv2j5KQt4EXmfJNx4xP8P0cek
Kzk58Fnyt7tMjv1Qkckv70mjtMsKMmCPbdIFipf7LFp1UHGBUGfIMU7aPeQn
so+2yy8iK4R/8inh/zVdMxWqRE5cz73KZAOIyxGrDiGQdpvE/sCetslLTDQ0
OIj5PMYv9UE3Z3Opbfxy8ZQKVlYBVHoK10fCHT9r1QzeTb9XU/xa5XIBNSsJ
iTSUc0sBEfx6frqv2xJMfzBf0IPIHzxz2Dr139FN7J8No7USsdqwgXmNwTz8
xNns855DKOl5LctvP/Uo06q2PJoYm4vj0aJ5GwmCjt1yxoQuojnt/aVHq0H0
R4EYkKQSjAInM+bghT9ZBwngJ8j0yWPw7anpvt7ZRbCaHGEulsaiPQrCFJZZ
E2y9Mo760QvqoOpPxG7JomJ7cayHuu6ZuJfVlFQD+RCHFXrX80FRJSWEzuDl
ttaN+4741t3FCPtHyty9HYwYURSr9LrCf6psT/NXzBXoVttY7JB3BDz4Kk1q
bjX/aQOu7+VYjX4tcDtpXfvdMcZAEQ8cq7szidqtMTgH+hgVLDbWoXO1fEtK
z5L85tL1cX/wMu0RNdJq/APnhKeIOmqUnqWQU1eao8c1i0acx1T97p4I8aHD
EqonZ3kP3zu/SB8c1weWrs1Wycv+n35ya0du6sCdf9GZIK31Uw1xbjVn6Ufc
3474uMhJL9u9R3ZCL13aXTs+eJb2jxT6lO6y++EeZWyy4vC6S1z4jwfiNusG
hSMgkpaRD32whlqOghuhuZsNfLMkqJrVeOSZpge47qh5yOqru2IsrOByeno9
kYFl1KJ/nQ9NzkaQBmwXg2fjDGt0lcFKUgMSFEmbISGiz4wW2ePXB6t5edAO
vt4Y3Us+rv7QdwhRHjrMmAPODIlZrulhJ0oEJd+CMIecaTJG5GVJ5pmXnC2h
ANoTUjuT+TI7dviuZ6xkCACC5qqxjgzH89pkSY6kuyI98ZWJejA4rn6cFTpa
LAKK1O7HbAGSg8ZE+MNW+mtMULf/C5kyVRNdiIVO9m1RSjuCUzrHBlQfhe5x
LGg2aGQSt8djfckrtrxFoRcbL2S8hezNCQjqtxC15osAC4woG/QS3gZjXkXQ
5Py4eN5RR0lSy2a86CZzwdHAMW9cFgmVSQwM5Khss9FBYeDJSfgBBFXpvAj8
Ojj3GNpwKIuC240U5dLRtKcsh3znm6Z5yqIYWeXtlklviKBY1kxzur21xDZR
TlzMcO53uIM0zjJaeWTwBkOMfvTqVUvRy0eiyqchG3YcxRmUS3r1xiaaG1JI
zov8uvPzhgPDgdlOEL4E0EMCEpsZXUiMzfNbaNNswrxnu2xZEWvQzOEGdc6o
RpWNINS+BxTuLAGWbtRNnNsobRint+Mng6wTe6tp/Mm4Jp6jlcK8SNThMmXq
BqDavXkLVgThNzEIYlfbV9iFwL/IVnLZEFrzIZJjVsHYKF1KShVdOYyYre+E
8X3fivc5PqiT0tHHgcpVUcqoPqG1DT7AusBSUAWMiEWpv+ZFmy73ENrvfJhJ
ELLeaUbiuuWj0pFMMJ1PxFsQPRMz8c4+6JD4zsmRZSsBVGeXlVUUTtTVxqUW
i1NUaTO68MGGHYT1nIMcI8/rbZwR+WCR4RABDvRJ4A4e0MdxahK9BtEDGcA5
jamwLdXSPkcUcRgYK9lMIRQkCZkQejA5MRdnvw036NdCHmCAcPs4iKCTzViR
xldpkhy8rwcwd8GQKQ8Ies1oeT2QRbI1QtiOTqws2W+wclds8jZNPTZW1Dkc
srAW9qoBg5rTjm/NQvfrArv2Ab3wsHo9wuvvNEh2jEK8Ti+8PH18fvU2XRWP
16101aGYNMwxLWGDrASpg9gkIUQjPbiAHiWOMdxzit/WCOC5jNpFZuOO4mGp
mtgf6V9KogqoN41kZ4mnfDZ/soYaPA16EM5IfRRywPNyYn2ujdYWxylBAT2P
iGeexS2kl6m/9NyvBADkinecPQgXNJbg/NGgopi3P+rhGWF6RgC2cvPM1TJz
0WKpdYse81yuithY4uTmrfkxBwRtEOU7PhgFHt2RRjp9uzrGylQwUFVouGev
/m6vCRU7VGyc2jMk7Um/GAMAQ7t8vfUqMPB8G6VUbsiuHaYeuFIM1OnRubgh
JQ8o0Y3fTCmhUcm9M99x29Iik0uf1DyGgJPdEC8NhmnlHc173O7uKf/KuR5n
Ts88AcwqF++2S1IqF4diuWrnW3CvEDsCU2utGv2wM/iVOKXet8YVxyD4PkEF
ZconKHJlmjmSM6ElumFR5J0Fpwen6Y/ZGMMBS64cJJ4GGXVgbu9kihwbQEDo
sDQ0MEnn8oH4jlsYRUWAZPM3XyVu+FG0AXnX5ogTUjl+C7EOgy9+aDHh2LLc
TFYZJB6WQEFz3yvXHXvReg/wUjphnP5bemy4gZpVfwJlgICxMbGMwPcfh39+
+IoQO5M5uxpLRgfrc0OWd6cWsmqfpANSflIQ8c0eh7WGkFWxQwtRDJqb1wlZ
SNP4Xh90nnB6+p/eyAZtb3y4auG8pgjlbymhDkI1OIoekoogVnEirsetJiui
3mCPLFefFZQvxKQJOP8wvmtmxM1OoDl42RiUeQkyBDyoIXyF3JV5zq0SlIOx
5LvcghwuOmbqxbpEUUpE1dc4gmZ14d8FfeB6iKUgMidPzZLLpG0QCs8iBdux
Py52Y51DM5+AzAXkiEs6UvZ9AF/J256X7MBqctE3SjPY0Zsk7EoHYlJV1sqw
m5xnuuc/egNE1aSgUs4J+nLd2OuQecxOhdL0rbcQtrfxyHsrC7/ByXO/QtWc
360V1ZMoynhAkfFNSZ5aZc7eLEka8a8LUGBkn8wwZY9JGKJ+fPH3UICQKA3x
6bFPPnFX23Q5DmP3/SbFiDkYDF77a547YB0FoFTiu+zfSDZlQmW7cE2OULTH
jQVk1C6U2pCAKAUiLqrIQ6n40qvjUY+EWtdfS/VNxDZlwbwvYXlJbSQg1sUg
RF83U3c1yYM0M+dt5+YBBhbhpIKFWMW4OUyGZO4KcZHaM5hrLlH3uChc1BjW
ooWFfiHejPeoDp9U0rSFvRs8uO6yD162Rn4anbijtivh6uPi4su8iy8En2ux
XM9E1JSWvXD+mBVbMfCERSKOl3kAE9HudBbW6qPVE9JxMrZPZq86IwVJcWLi
6H8uzJsv9AhNrNmV9DNJmdjV7oYzNQfZEiLPXkSNka4hfMoNcDcZ1YulnnZF
Q/KSrnppYzP1ZEG3k17WkIRuzyA3GRGT/ZQsDR/M4FoUacoQ+pKhCgf4YRmU
2qf/ukpvcGLSOEtIw0Yb9iBDjO4OAbvr8o3Q9i9K8M4Tjb1vRWvm/qKiI4OV
PhKWzrwq8XdUINoYviOUC1F5LEr/sLOlnI/hbGNcuB/ENSQ2oxMgUau5kijy
xzLK+qMsCvgNmxH9/fGWDTiIOoj1ztlMfZQJJnye0VA6P2Pj5LCkjw7+5Cu7
Zr7QIYMdSGJuhNmztUV2upnxi1ornGfkg221wU1IgOkSFcJGkAS9tQcMcFAc
WNRTOUCWZNO0rSu+gBCDglForB4nKqHgyKiv0iotrkmqlPUfiTMhZJt2YduZ
mH0dZXOKIPeB+MrrSuqT9y7QHOWGj2QiN4VqxGYS1AdPf2IxHMCKDuWGLd0u
7UV/oG6l2iwexWDHSTusyJRkPfWI+q2rhx4h2DDnaS0dG0CCgyLvWN1NQkNV
crQs5bqL7BvDU0X2EbPKQLhZUuDxC+abektK7ywOE+hDSAmBxRPX3TNZVwoF
Da7Tmt5gqq6vINJPzhHSGI7E1xKMqj75wz32qmvZ9Glc/5bnBcGBtyQ/xm0O
XqUKZD7DGoBCqSFpKBK1bu2ee2nlwRj0pZ3j9bmFvX8C6xjotT9vyHMbZwtU
KNr/LjY1NdQ+xyDxb3pVviMSR3QnSTFWobD+EER55GTBhC4I2C6tkRQaxVd6
NftX/ZmGulHV1jbPT/13W9WjlB5miLxp42vfAAPyUtOZOFOB73D5nx3eBQcI
+nUxfuCktFSqR1z3ayQpDquGAr5O+vgf9fx5GnmwMc/JeIlW/4DIlQ1obTs0
BEqqq2UapzBH39qMbOE9zoDGHUHl1UbLzgZaeNNOKxDnJJwHdY3y8uCsO3BQ
MBhpzcd2AJb8QTMqkOH/ZfTbs9A8YFMz+rSZW+uIRIaYGeBt3nO+33DUYm7s
cw7Bu6IeDftMYQQskWksaSoI6wiY0id5ZWAgJk8I0wqzudh9ox1NmPc+jqUU
dJ3lbnWUyA2BVa7MCIBybPylGGi73QEjA5iDrQ51qnz3Er5t8wSXnbOAhQfN
2rq2QDe1IrimiIlAgnFNQZwrm/g2SAUENQYqohvBl5PhG6NgTi9CbZHRd6oU
JgzU819XkUqEzDUlsbCLnmpeTpKl9VfEi48l1JOD4DWgnTpTsw0M+XMY6Hq1
p5j7YI7ThatHSeBo6xqXkNLjukJLzuohkb41dsESru+DWsfjYH6fbcDYN+86
gOk0yumuk3e16E68Q9EB4MxpztFgzA77j512cFDCJlI8RpIqEZbpGSf1gX/E
93e8wLqaMMWGX98FxRexUTPEmr0u3dzVpUDvY+CIgL1RRSouly8Lq6jedBAm
1Pg+14NC8AObkQv8vz/7attk/ezkGDi928dA7hc/a2NchuYxtnkQIWg9kEL1
NpT3Exzmzx4FkkwVHCXPgIuNDrZBI20TwqlwxJYKIfAX8XSPyrx5/Z0w2oMg
Rf/WxO1VkJuBszzzywsb0i3LzMCJDWawS/tN2PJIWwZpe5Ur1Ycsnpcshsvk
qr2ewjygYP1uOBYD/u1ZqtGNW7Ofa3D0zViJTyLuNDk8o4qt0Knr38aLNY27
c2PydPE0NqLe5aZMnYrLZlBoDMuGLnEQbRvizSePP8+pwBA7a+NCYvgAXjx1
Xa9spxweARrR96kkpvwm1mGt7KlO8OTuo8REZjE4+Tk6jKPLtxUbViuZik8h
WKzZGFNR0gv6cgMr4BbLQerogRAB2Dz/NLLFq6f5oPw7gwdVLFwlPH4LNY4C
tbTb0SQ6Jvlc82pbBKHvVclAH7uDa0LI72Oe3HOEF6XcPHCnG/lU4WHriksz
6302grUQGS2FWI2L51R6djPaviTVN+zIvffpjBa2MZue5jg1uAvd1N9T8GIu
0LCUn7DqUgTGtdxKbQolnl2aUwZPVkXl1Wqw+rCCcLoFVdC+7m/k7vGavqNK
c8CiPpk/TGLuU4mQg7N6J3iuMnIbd8IEi3rogXSaJjLngfn6JZr1dzSqu6oE
ewNff9DajxXBuGAVDwQgP969bkuwQoeC08cVEm6sr6u0fi55BGvKOvGoOunm
nrAaqG0ybnBQylGbERVGaPCFa2wxqYCQAHomhLCUbXJJ85X6528R+RY7rzqV
Bvz0kEPpcDCNkj77KDtJqa/1v70UCHSRkpbRq4U3bvbNNqCP0mjBASv94CL+
Gr4w+++eLSU9jjnRv6m1zpQcC0pG5ODwhWql/vxdDj0s0jQkyyGcTClCBoUY
Bm9/kXYcgqqyuVK8x+avPNS+Shrojhf7a0WCiBGW4t3FA2MvTDBsgTC1EkdB
u4yJHKn4d3IjiPfqO3pSYcETKqRsUSDMf4DbJbfW9aEsdLnkh9c2ULeTFnDe
rbiSMc08WltTLG8b51q0QOa2Sh4T7ldUiTNTbTRsnUYtJ5501ycDNQefSfFt
TYoSC87QgZHNNtgeyh6POz4bsPGLIgNJiCtVlMUbfOdQlIMWKLWmHb0Nmj/N
I2TObv4CFehlrGcdois7V4c1xKPxtpVOzuPLKNFV+QecdFHhs0oVtd9J008n
M/T2yb8icYJQnpfUBKfTdrxq9yHGtTWmzemihGtUx4Faw+Gq0/Gj9xFJ6BYt
MxIZTJbk9F8xA5eGJMbwiz+2Jy6tHWvhVH2sgwAdTQtMBy3BLBLA+dXu/04M
akJJ1xk49Tj1YT6m8f6CuYbpiaBj8ZfkmEe88k7pe0cd1gW6dUmT78CrV6Vy
HuBaRk5Dg5DL4gLNTQJo4VsjBKAhD0+XuAWdwCvuJEmIeELbJtD0uH5qXVrY
HO+zkGCXRNG6EKISaXTWu76puxStm1FTazUHZRSJmMVV37j98AkJ64u9nF/j
0Ikaf1sw7pzAwNS9wk3oYJHK+PXvdiKb5yx6h5DQFPcNh1ewdD/MwxAQwR70
cKiu5pcBw6d4Z4wvOokkinhdi7bj+USimA97jlNQymySpxPg9kzMWD1W3OLh
fMYpBG7NhW4bbBMqF3c/0qnoRgFg6VR+hpnXVAW2Tiky3BnqEl+xlyem9Kgo
bOuwFFpHBW/DnhAKjPIdq8EPfrl0Y7j0c+EflBHVsuqtL6+KEYnEBP7Box+l
8WsXsGrGVqLHguqBZgSdzyHXlymjYwkAjvl6LOdZ9IeB9+nxEUOjva7GpNH3
kovWSOPfgO6fo0e7F9GEQU7VcFIKFaF1nONS6d3+SnXZ5YKU+GYjoi4VfO67
d36gdaZ+aNPdR/GUAnuOvHwfBpN49qpZTiR8yK8HEvONLZO2yb/fHxy+A+/w
YZhE2VBnsjWokGXbqzVjDh3Fk4U5hX0EGPlKwNHdeezYQhyLNSiseDVv9ztD
m1jz/hj+rxR/uFcqrAm6UEEgCbwC1KGnGbG/IS1qcK06Q1fg9AN7CNBXDgJG
g2JQD23B/JsJ43yPk2boD651eMDVttuuj2DesK92G278/BoADzjhNMAl5uvP
HVYHBPSugEFG4yjBW25OmcXuRaJpIwiomzpPey5pzIR135/cIbbU9ZKpoxjR
XzBlIs/pvQMJQfBAsfZ6ehZDF8+xutZ3456VQuWWDt3RBmR0us5OvjNKlWkF
VI0Dc96Hp5knMQF+OQthVLUQ+cvUffSDcACXiwwKJL340wC3vh8I2Zigw5do
pwwOpKTMaB6Cr13ji1QpkgqyJbTYrkug+yRkrydUrk/1iTmMMQNLuw6nXwBI
3gdHQbtoaFItR31hLe4kZS02xj3qDng6M1xJ1WUY2vurIT6Hr/1GpyibrhQk
EAz6ZLehLBkRXbqSJrCjXUn+RrIfOqSKgdyP7L55dYR69v8RUMCbfBw+gVhb
L7iS849mJgIFsswBdnac+LiPSFo2AL94noykNZqHzPQjNaaqOPytg3EmgmHN
p3p7RuOllNfbBsgYMz9INrzP776QQv/6FDaX3Ey3Y9Md/hSXhHz0GhuiLHM4
jBDSLtWLBuDmUOjVGBG8hmz40+fAo/k0LiFovRKdNhAbPmwtPZouvr1lIviw
VV3/ux4tijjnRkgciU5fimRIiwzL78nk/f097ZTFY9UqcOT4EyJh795K1iLt
zsKsICawPK2NQTQ9Kj+SP6GpXBFk1pbmgqYhWltuv+3rBljKbaZDBcGdG2vw
FxHy1lpFnu/BP4HOXzdR15hBmmhHIDb9wo2kxfYQxkWL2tiw04oJ8BLQW+V2
jfE+XaSlAw9wWYU4vmZFlCC6uAQgEPck6myFzVXmZ81N64KSCA/4XrAsowbk
urq66JtaScAF6arjw0C7zMmOce3IM3QzzjaeDi669UtCWiWPvSX9frvtbNvN
W+bSHTFnSy7SLmRHzKrKQDgWCgmGQQEZjr4ADEPzenLkGtewo0vzYF7XBWqJ
417RNz4qbfxZ+WSBf9GS5kPWkJjsVFCHn1dMP11TyTEoamfL1ynlQ41KZOmq
9n2fPJq06S4rQ+TeJhP+BansYnhdOQC50J0QxJaKfo752UIGHZ5T3CVATN/Z
yArUYxnf+b8YTlOdwnboheLwU2akM8G01DCFM5kZ2Kvv7aEmfhmND5cSLQI2
J3nxTSo/cDol/VjqHtVNJLlH8EFpYp0OzjdF9QAuIoKyrejK3mHnknMqLHVx
dz/2X8QzyN3IhkRo5N5SHNfKZSwbu7ycsYiPL8gLoet+sl3jUue60sQjLwLi
AlAKsi4dgWxBge1ziBCSdxEtf6mnUdDe9kjOCW8jrxz2O55zOLiimdG2As9a
nHErWsv+G57OdBFGef5tlo3DxAHQpCInI5vCiU3Fbtdh06HYNCFM3FAAIZF8
xUZ50FhqeYfoLWUqfOq/fipF9SrX/xZGlqHJvWbBSgxN21CQ3Cu0yGC1+XV5
Qw+IJB0fzSv6v3LknrZn2Pt26r10xZiCxJgF9BLyAaofN+dqNpYEjPwP4Qqd
Dm7PM4FhASa4ha6tDnfihE5lkCroXqc4EEKI0DShjwCGetfP/W4Lat62UbVB
KrqxTj7smTre6LcCrwo27w02qUi67/3sK+6HiBUs0F9TRccEYjaQ3ey7scbN
mRP4UDPpScX3gnL8N9QaO4RkKNeHcF82pns+OB24BTGwBMH7S0kU4lpQ0GwH
Iwb4athkT68JIxE5fnuNQBCsGjHnwT2kvfWFGM6PL35DNhImOW3wXxZnxt4u
mIOc+w4/3W7UEXaTL9nPHFMxekak0m+KrQOueFEpZYJ5bGBValk8/kN5KQcQ
PBXh6eIBugiEiUEmORcL0WYwq3GEFw6p75xatlMjqAVg3Xi+yyRQCgzTGL+v
20G2FWAtNR3OoAwkUUSRWBGDh0YiNLivFdhqqNBqKThrOWtzRJE6P0zSdl5C
cqRSdJhVe/YEb0rq+nZxo2vvlkdRq9M/vDZpxPNzZKfzULC2P8+GRINIf5k5
bAy3k+ACtS9CbRHcKQZhqhQlkocz8rf6sfCS8e3gDAC193kFHjaYHEWn4PTo
r2f4dOt+ArR3HS75GWxrYZ0pW5p+qw5HX69SYkCBFdiLLHYulM3d69tVtlCa
XmEFgWejJ2LSX/kAmQkyEsQ6r38cVFpj1W7RbM/effzTZFNV4qzxaZ3x1FZ1
CHxGci6zsNkpy9Vy6g0EfF/p8W46VAEuFHhpCks8gtpTGizb7jte2fKbipo1
CIbJfAP1ODa54KwvETfX40Ms5VtZKqb1RaDxRnZBOIQLSFm2VzKvGvMK+IFv
a2D9OZZnfF9VTlxJrwLAU9vPju8VqXZYGgGXhQK4pskQsiHWfQMioAfH3U9w
9qgxbZ9V6mKS6/og2dQaTiHm+C//SD9lUeknjSJFi3DspbHuthB2AWirYG9l
ZBNlTwr4i9Hwz8a6MG+I1gNZiNLeNARdIYju/OQNTpct8pAdOjIdD/Lx9MRa
cak1W8pcvOLsnKJmi0c/9NcaeCEjPK6lTHioQ3otw1sEYWG8pQ0T1wDB6drN
azFikg6E44mmpuygGPw90fwah5SlADNczF6LsHWRc2GxcYZ4kM36MPAvuUGg
FMb+i8yMlcsetI3BMmvnkkUX9q72/KOW3OHYgxtk1/CF7BaenWCSoYBdDgEr
+4bxGUvi/OfMA8qZ2CnJcsvp1j+rDJsDcfn06fgvd2PzbeM7dohsOKXDH7Yr
A7XfcMvARNBS3Tft6z5lx2bm2xHOFrQGEFJ9735DdYcd0J9BI9l3/m40q39I
F2uMa89dpjVFxBsL9025qtAROBTf3Gph6xrscbghTBCHnUvmjxXyqmpnqRMl
2tSAWvxUJ7dm163SGa9UXaySgL3owf6T4S/ZDQqjWPQg6qusAVydxxBsQlpd
Kwa+yh9t3X4t+8wHIIaTYy70/mg861yQL85RXbnYDYY+WGIslk8jFGcZl+Dz
SVVGKyOICQt+qcELLMh2rkZgRGA1D6We0wXQz4tenCI8m5u2kpXgDzDE89UY
UtjZZDxek3F1LHu4nCow0PRSGxHp0g4gJjupI4Dsor8mPivvbxS5jcgXvRrK
6WWbs68F3UCgzvuEc0ryeY92lNGW6gWdeBK4E76p6md+8Ck5AVapwJ1xHzpF
3mBO0T9gn12Z/4Pfe3Cq37LTHC2ULXeD12K+hW0PPc+ETBJkvsavhD/ejaaN
o9nIrOCkUSQfZJJJz55Nze2b3ThJ3+vVM2ztqiAhtsWJfcFHG19/AHNiu7yM
oHccjWlkjNCq4BB1/pSgTk96r/35gkiZvLC1Ul6HSyaJtWOOxquze1194gzF
XTzMWy3NU3xQWvmCx6EXXOWdVvMdHtpRph1876rFXLIeIloPF2l5llbm9K1b
zhspV9IotXAVVT2jGkydwtvYmbjhV00EN4glDrCfosrBYlB8ls4su7kBvJXV
UPgE6PnUnDc7lH9dICiE/k+507xom0pEh78DUBNiblE1dmT7jOd+Xq+jUHYk
EojqJUErEEiRXO/mINO/FzYM2NlPTuMX5mf1RGZ9zgstNm39IP4vq3r6iTxH
L8SPJIFLzMQAeJdSXClcsAEFuICdkraVMHmq3p4T9C1dgRK+BZ7kordYaSha
oSJFDCnJ6Ed4iaNY0JQrfuPYhSum3RFTtRKp/JMyAuRuduY9HUgy+MGMrQ+F
SkvAJdK6qxJvH/TJFofhQIFQ3MJMjBPKsb9suEKW4fj05ILAv1bxY8fMHu10
UhfvCuqkJjT/Mhmz5iGrC2wj2nzxd9DBWEIg8P3E0kcLgu+sQwFTaUSaHoyi
HUCyha2JLrBPmnJviIicPamui6bN0D/5qifM3s1Ni4GYML/vay9mDXq2TI+7
G+PFWH4VFHID+ERU4W6S6m8kC7EFnuE1iP/uN3ydsaDXvlkzt+15XB8qdz3B
rxziICGUinnJMz8RuwPy7DVGlqYZ+EFeb6ml0h3azv3wkskmWgoTUovhrfou
4yFsnoUK1U1kNFjEK58Le4QBbWfPSlmRMNseow6/Iz6QgAKdWygOyD7pVFVd
3AELpWaztWDAaZugc4LjcgmF+Rs8yatY+jEp/+b48p5daKNlaQbcdW/aAChP
S+Omhq/qWFCtXKds0eU9HQSefq9vYqkuCNeCYeb56MGXBVTZm1e408G/aYFw
slcfaiyZhnA1XjV4UUSCwNQO2hvgSOxzQ4i0I6r70fd/39SySbpP9DfVFCRf
kSLbqAoaGhjJmrsiHkZ1MfzM4ScwIDOIFjIS61Ezdb43qrV25XATbPk7wwMi
bq6UJV3nzc07tEVOf/SKMd9N2OyVsRCOAavr7RjpgMi9rncDO1sj9kRbrx86
jYj1nBILPTSau1xX7G7tvH2DGeFv5DrUG6mZBFJSyQwLYLyRhUy29JPE8cwv
Tznj0gELotAPn0Ltw2S2bE5EpKywQpuf8tL02T37PV3D24+HJw2r6/+qq/il
yyAKhfIymffNKOn2Jl9ZENqmywdZsfChfzBBHMq5XU5MeUiZfrNWo/qjxGZY
L6HPuCfwrjFwHr8EfDGDpJWDO6e2BEikxTAEk8poLpfkk2kbq1invgnF4NVm
cmwhTS4ALfxbSVBB/gwMm3KN3haqsBqBLC0y9OU1c5upmJY64mjvmRUgeCRC
XnjTUmkWtOSLQcAjilaG6TH0RHN3LDfx6vMWLYyxbvPqvwbtbZJa8lXJN/+8
jkn8Dc4L1A+YyKZiu3LOqZ0d0ra9vGa/KCYzuiibBhVX2mHOQHK5QP12TCkw
VkP5SDgwVcrSrrIsCXGvcixa7Cr+bAYC+bhu1a8ASK8ybL4Urr2ZXwKh4Vjt
sCK71qBQNsqM3wo51zF27/q3gjvDlmWz3cgoINjeQeDd5CVqkvJNiOJXSvx2
ZeG5ilz+Fui85EBwiTqhKk2OoIK9Y4pIFrwjShKGMLNXSZTybf2KIHUcZplH
LXhmoOFgf+/Y8cLO9Qw39eHy/IzhsbR4IoDq/RBtDxYo53UKezalk82Y6jsq
kEXIFkqKi9TLcpSgPLx5BexLma/hNjLg5BshM5cxr63FmRcnZXUI7HJfzL8r
oC4OqRo2TEbOfbCDAgUe4iIS2Twon5DhvUhyqAN5bYkN+n3dCmWw9aNjSdnc
jErOnw+GJHRVT4AcK+vpEPuakhVlk2dlVMYiB9PHPx3BvRu6hDYJ+DywiCmi
WDWb5+vFqM9kr0u1HMHqCOeaRm7gOonO5GUo1/S2xmI+lk1JdlnohcVjK4lN
a9jIjghsYN2p1G/1qIodNHMMBc/SU/YEbDJDVP6clDg4T4a3r1lHdsDfbI2g
Bg02m+HO9zJ+YmmGq0UTL03mRKCga5LmLwqBzjc56Y3AZx4gXKzM4MB4iHL/
ZHDgdTPFeQkc58XUThYVmQZB19TRSqLEFG2H4TpN8eJx8OqBbqe07cnnQdxM
gAeAwztszqxV6IuLAenqMR/XLNBDo7zjTf8kOHs8fen6Q3AhFp1+cFjQ1/r/
YFsavUsw78cfkq1rglzHaFG99dilIltHHv+Q9ex7/w8HMI3d3sDBrafN2mx3
zC5yvvhNpZ51DG3BBkV0fmK5+DCqEe2i9GjKtBPJsQpEoToYKH0h2LZ+xRRw
oajSGx8FwN5bQ1uvEXbLB/3ihNRdLgmnaZSKnhkiwZHb+v7/++wSiDpyRUYP
Mv7bxTNY1/HIGHTYCv7Vp9zVH5n1SgKkTeMDeDvLH8F2CJfwnLa33abGdSK/
oC2kBbi0uRCvXgYC9WpITBp+C2bM+JJZvuyHGRL7ReF776XypUQiXkU6BFg7
1DdIQGrykRBTsTMXKWUWRJ1qwaZ9iS0K47KBeR9jBLvfYoJPf/FRpc0UAzGv
EGw/pxiPP26qzVTbJybnCq/mqO15DyTpOApAGnnLYsfyIId5LQtkc6smJXbT
u8osLtZJx4TuoU4849ggS9jNn1rQdqzY+00bVaVi/rFoacBq49qzDjj0n5h+
8RRkmZ6pdF0OgkH37K0a/4ym6H8llH9uUyftLMrUlZPI4jY5nbxLkX+h1hSF
NzT6j5Z6/716ZhweWtQ4WbdgNyFKRynVhVEiVEoUXuMdyTdTkBxJV4RenHNK
NPShURAb8dTlUGFx+oy1XPuybxD+WIijCZs6Fic6bDiUEYu+iGLfULz2coAB
W/NvPiV8sIyAoCjTIKKXWg0kEHtMXLF0Kypw6RnCUvVWEiWVPAn8w5f1xI5N
TMR07F9IXA/vcTw9+Ix/05y75hGlGn5rSC1TdKkKEGz1hH8NmCvkfjxYXbDz
J5oGVRQORcGNI+vjnGUph5ycPvuhI7WUuxr8ZloV/CcMQK0Ed2W02f3+7ZhM
eXFLLwWAGYJdCt679sALSwOHUs+TYkKqjVLiDElVTOQh+Kca4FTpy9hjDh3d
90CeHRq/h9oe9jDlTkpPgaiZCGRIBcoTpeILmRAKZ79ZXZ3t9gmUKIVkzbd+
D4kWj6FHre/9ORMeStAhD8UFqTo+iaSpDzl413b/kI6JsWOdJYxMAQkWlpF5
SUCnJnBFBTU4V3QQ6TqX9jHxHWtT0h6TyF4Klbk9AvFyjjoq8E7k+X7MEySX
PE/BGxUw/GgFMN6lCYKSaVBUe9N3YuGiuV9EHGNRjngA3YBqR5v0wrqJGeRb
k/v8mpXFtNnZfcWcC/F82ZfoaiqmZiOFVWiuTsu7PYgOuLUYtZTxbRzAZIlB
bvkSwp9fOXCUxLkijYMmvs3JOSf+Pb/CAQOiNsz8QrlpQUAPREYyiOabepNE
2CD445eRAESIO5horVTzmLU3lXs+V+nakYKc9ltRVT7+P1q7Vs4AyPrcoYEU
A+mmEQfCQ1QNOdb67UHCIpFyVStwHuECYOS54s4tWYyXyKjaaPGjBugMPJcs
B1LDiwsWT3zlTbv+NfbPfKrjNxJnkBacp5z1/rcVDtCQtTbpnx4GyTpLmOHe
lul0XgiE1vP3MxX4KDV8p+0RcPPUy1ZwNVOT5842otHvFFDzEx7c7XZVR2Sk
AjJXi4qSfAXKrIVwMqV319nndQ5p8xPrrc3V/jv/wKs4kEnyst3XMn5C0iyk
1Cg9rKsR85bCuZ4ZeenRXU97SrqLuf76/graeiAvrADmObGXeLMPGAXNgCFg
ME4xRvQ5nvrxIDKoOiJn/2Zv7lXNazPQjaYWsI8wn3i6eeg0lOJj6Fh1kKzm
BD1B79LRkWU9K3VJdksiZnkByP9jsuPMSlPVG8uZhGXXy1QqRcq+Vq/IQBBe
VM87hMOsB59ICVqYeBtPDo3JVYZGRKXmFNFx5wQ4Mc62TbAf6Tt5TSSTgRq8
P60uAtEPmiOeK7GVlUqplZqJN3xrn93UhpkS6htfCditFG/iuKan1xJ57jau
PNbbSZld8W/QyGjsRlrlXpqiqDIj/B0tWeIMFMD6A0nhxveh73IuYDGon4Tp
vb6bz3X/C+MD3RbxOk05dWdami5vuVkPB4qQBIxEJBX9/mfX2boFwyxVnvSQ
YkyLlIIGmlSyk4RzkldfX38hI1nnPRUpIHNH84NIr2hWN38YgXIz2sTFz0XL
aRa+levTK8TkHYRCpZHcl9kJHHUoIXcIJ2qDVK45AvxDZi9dZNPiBCEgKNu0
T/bCMXCpltCdFLB42IGQlJbQK9LyLOMo3mNwtXVNiQAh/orsoauBVrEhHEpz
yS03u/Up8PH7YTaJECC2RbcGE2ZBdvvZnsbhllbuIBSy1zaaUrL1LXh9e1fc
18bJBVRb3aaddMCRLMoEISD+FSoRINXHAGJWvTX8l4qPmhNlwRwLGLRrCyZ9
8pR49QN3Q1t+PV+XldlJSIPq4HjuKb9uizhc5w4m9vyeyBW0qwTfiYywCVam
Nopfr3AQrg+g6+683eiuaxRgCFz6YbR4QfSyk6o1pOVZUDoNNkf6RsHoFYQK
SCb4tMb6o/Y//VEjrsMucy6GfaRgzk8+GULDtytX4WXGk+fI9cuUibv8QVEP
e2KpRkZPqRBHOeEkXoq4/KNvD4EUGL5ErHRUsLJEf62lqzXaTtBMhTRUb/cq
No4/EhNBNjxHaXH+bQpDL4ldT7ogqENlfyAcpZe1ntUViS9ouPI1nqbz8PDX
sN3aLfM0ZE2tOENa+drthqEk9PVh8sRL5oaRTwJtJZUFCIpgbi0DG4Ur0jN+
W3VM0MceIQMaBDRbMT5h6vDXQIlknWLqmvAR1ahXwEhzMrQfwFUblVqqrx5W
M94ox4+8Vh7cQS4XmSvzHilfd5SakuQZgh9iwrjN485iEnCw3HG67yRwiAUq
M9FWZW3Sz1nh7BAXsawwAxn4E/x8A1k2PAc8CTdVDGBy7kX/BHcvKJxeNQU+
RTiDfyVON21AmYlsUuo/EWDIqyZmjz9Ch9OBM+mXBc/dcFcMDacPz09qYios
kFLGaPVAHtpS5J/n5kIvP6nu6JAlk+pzRX6aPQ4ncSsuM/3MkE9c6aaR19/U
AuHN2YAXDdgHVm9EeKw1ePXI6NbLQ9a16Chz/N0aLOwGH2K8wqSpSn2RAixE
Lzast+9WrgwzqIhWRrDN5ID1JtlORil2Zk1w/VqUW6nx3BVLNepmfjGKSt2a
yAyEWP+tYfv7F7E17gMJ80YckLOW9E7JMisKSm5NapIcasr/dx+ljpRFzVJc
LxSyipdz88vIDNHR8uBw35jEdYz1Wt2OSGCtofRChCOVBYZ6JVxsIa1sshqc
8+e0UzjffA6NPbrhWGgYSJuP42j3D2yVGTM4EYzO03znbGpgdU+BlOdg/dH2
jEfLtQFGAr5xjUkJNPLCIeDsR2O96BGKRE7/bZLse36kkria6DcOAuYAc5XM
hVoF3hAgf0oPFpxlg0g9psY+RSpm+eaeUk4auBiH60duWNqxSpBrpBHwuZx6
Ln430usqW4zWNGWQMi4wNp+NhDKQ+fWrKfAHNI5NBTg8HyIR9g6GaYnLbtqL
DcHs3/ohD+Mb/Ftj6vADVP6bpLG384vqaHeLGuBTqcOzXqWF1uWdH/zKm8rn
9ifTABHggxSkegmMg1v1eqT2AURYfU6S3cgHG/2EgPO1NyO4/aL+zeBpUDOR
25WZIdTfTdohalT3CfavBubjL13l+xh8t39hreAi5Unugh7SvvTpbbl17Egh
4X7pT4GJJborct9p0ShBed/iCcjoC1xjFUUYgO2z+WpmVV6tXYoHbrzAf/eV
p7kRc90jr5ekGlRBcleLnOUbWIiB1Cd1tV8/TYztsVFq/PIWatHOFRZwRixZ
D749Ot6TJiHLLPxl5fJyXe9ckwFECTm8BMISD3HMAjdO5b6SAPp84ugG2s70
16OpZewiUzgWm3h+l+cp64umPUS40Gnc6Gj5Ifx3EZDlYzuKnt6z2+WxBTcQ
VO1R9Np+A2fb5EFzH0itweaa2Z0vTKifdRefGx3F0CxkvPEWi4QTR/TWlkKH
9EZrTEXrWvV2KyYNq5Pvi6wiTLYxruAPzZENyDWhBt1c5U+jmBVlJVCRtdRm
Ph2BG70tAIAk3ADrzR8SrzLKmPaEfe3URo/VL6Mbe1pjToocny4rFh2Fk2za
URhFoS2UgzZcs0b1scqC0sCyK1F90KiiJR+PiNRaHK7mV6HNELXDlLnmhhsq
5RHg0XPUvBLo1cRxcITSjhrlRxhd9L9n/a4jeVYuz9GvKGwk8qZNP+dX4+A5
+zKI9lRr96jX1+kSdXAP6BAuKcc+L4U/OI/VzixB53F30oChhKHBtxrmGEFu
QBgMmU9VLIF82qad0T+MUa0oSZKJvW40WSiTz5NvsoE7zfE0EFx3cz0hY+z7
422iE64UFR3AlyYXmj+hAfgY+69jRic90mflZp9+1s1JooHqJ4MGKmW22MrY
MKOSW/0epp8bydrMpQITewa164SysAO3zOPel5Zip6qT2mZUeITBaEbS6yoY
bbZrxDqV2l48ds2LNz1EAIHAEmXWs93Kqv+TrjRwbVtEh+X624TCmAW0G2tn
7wsK2XtWcrp+OnPV/9i/jY5vN/5umDKDVTBmLhnoaBh6t92RnRCPo3NpheVc
Toy8hVm4hFMYWy6anSYu8qIBjhEXdTt2fH6FroqzdxsglPbvfMh2Q2e1+IqG
teuiwWh9d6gN/vUP7S8iFmOfUn5vPq6xfjf3yRFeY4ZOm+8KGvVpLRWr/hMV
SYfR6Chyxl9mQjyJO2nnS9F9Nz7/QQBZkoacxm73NHQP/JZb84klEmLMNRVJ
XuucvCoeOpLBhEAkpxeJXCNq/DWx9E6fCl4ncbUUmPTY49JmXlwNY1IceHuP
z2zjiY0aDZgqzDWzO2fXT+dWRSODTqP0x3qRpPRGzWowtSVOfAUQ/6ay/udF
eIfnKyDN5tCv97TV1ZnMwYd+zoSYc05kjLV1mLb91pc9Fydo7VV14eI1HUpl
dqZjJ4I0TTHrUZ2PT0caLug6n3piiW+F9Qj8ZMoDHh+KyLHjokR9empnOaIM
hnAYb99XPKNY1Chcu3ZwLrjbAZpJBFwQJspzSYckuZ7BRQs3Z7oFhmzT0KAd
JBF+n7sP0Rgcj5GlDWJ/ZPX+49A5h3pbbDcV96wLEjhsctckhC7FavsqbVks
XynTxdsFFm8xOLekjZKH8aydDAkI4r05DQfUhFjbVGogLGaCP9R8IdM72a00
aoPwA8tuic2Pk6cLIh1fUBeh8s3Eh8i/dQ5hRTYytGTA8Kvs8dH+JXnnEOBM
5mEvbQicrTBtglag8L00RoumF9uORuhapPJb9G4nsdAbDa4jAzgULyocMYY1
UvoGCVgeKL+dw/8b2duqwg+Eeu558Cmy/SIh2QrE+H9vLBo+dQV9H2x2+rdp
+Y75zl3C46XgLJ5W7Gbg6XbXYFfppSYy0UJsNeiwLF/mtReDUKujnsIBdUh4
Z+PcpP7SSl7LdXFEz/eH+T0/84E8lF6xY+UQBRRX/7J+aZw+0/nfEX2Y+m9v
WLl7inbkKLFKlvi3S9+Laj4KGg2qPfo3BEJ/jr2RF3nZDqfYH8CY4RP12PmU
00wm4lNQeIySCX2m+/H8n2J6sEL4BWWqXC07GStLAwODljWZObt5UXRgOIon
AGOHbWXYufFpdF48La8EsdWWf9B1x+mSN1+w74gIKiySnkFrDczZkPaW9UOH
q3Kj3PKhwrR0LwGeRCCt1KfJQKM448UJOAMFZD9/U67+B5a259eptVxb257w
md4dRv+o9QSK76ljM4nY9IslUV1EtfQcKU79WQQ4LOIqJs6WDD7TQfZO4RTR
L5HSh91Q/An8rzfkqVfX1wR8cw7baTv3XCQJJ3TzZFo7LgfGqFKDKU9MS/fT
Kee/QMlq8w8b1sZRBixqrsDY4dblmQBeGnYSi889TD3Ar4j5gex6/+DC1Wtl
3h/2PAJuv8Inva2HnkcaApGWVIx7EYU1zKSmGnWrhM87MfRoYKBRMR87SCTR
XVNa+sF2f19cdMw31bTnk1RMoyHQ8+0ds0oXOA1DeyOhiIHlTZ4TESJo3Hxk
urEHjVy08AcDvus8bDZUv613Gcuu3KBnzMOBiQGyPugRyuluj92UZ4LcAn7f
H8spwOjI2UDz/pBxW4Jx4nQg5dATbzcUyhkS1/K48wiMhzg9Yyy6jbcbOAoQ
Qmyb3GUwmr3O0Gi21bApYn+4L48POnkw7pBqTS0VGmzZTb2uovwiG99b/fZ4
e3olo1Qq+ruzeFT7Xt+8YB4548FFVz6uNd+PPL1PnTccvEweOfDhF/QT/Ghc
xit2k0h0qdw0USxiYh2fSnF1SZbufV9YXk/m6vq2vBHqvUelFjB/+hhOmm3O
lI8mMgVmaqKVf2TP1/Ytg+GwuEoky10xvbxgJJLqjCa95f62nIj5k7HIq+zI
ml2JZuNuhsEVGU64g+gd4e3pHu2tCP/vOxaQ+VO3CKpDHMfN+eWG/rAF7X1Q
SQzL4Yz5ZAiZi6KQfHVLhQpYE1cxpFeln1Y0WprEqxGwyaHmtVv525zkd5EI
jUbqXJcJvPBt0mvOw+p1NXdzRMPfbLY1teB3bB9hmHE/qKw9vqX4G94pIVWj
80k3Sk3WCeuEx4Kza3bsbpL6alwifS0KURe5SSArlaW+LVzg/PUkEvsnUqz4
xOA85LxnURtVzHJEcbB+mtcBshZa8HrPvZSNZMa002hIfPKW1xQ7I72XxF4k
wdbAKq+20WuiSSTjATE+st1P6DkooGC0P9rkiYN59j3pgP7RAhIgZpHtQUTH
EkSg7Xc/SMOhysaurEa2F2Q7r3mCT/UAO99f90naUyc4TbHhggg1l78WO0en
vdh1frPeJ6Fe1vmCuUkctUqNF7ii+j7hqZsr6HquLt2cBB5m2NrzczeodYGF
DQTG4zuGAgSCNnGYVkAORxNCyYzCIEF0pXjHJdHioHj53QT+1kzJJSk+h26X
pLwH8oxx3aC3ML7SJmkvXviT1uWAPIuTE2hgzPLtWJGAlZXA/gps4d+11qz1
U4psIlFOpyZSIPWRdfcH8cjYQVUgSVG4yG2Bs/eslmPddyLHIc0QWPtQ0se9
XyU67aBOZPxjtvJArrxmTwujJFuNJOZ/+UhrbU3bQLbCG6BNj5El0HDQsDja
l8Kf3Gwm0eNwIMyRsNLzhMfvdpYeZOGI2zI5WDAQSAqImqbKd4nVmMU5n655
JummWb30fznFOCgMDo8sr7sTma+HJ1oWOXWuuOTv802BXwCd+F/scoWbdRji
KuwQifRLHHtoSuvw75Q68tygCd6ii6O+woCbJ+KUZuMZmQKJ6pAHM20IfLF3
UgF80+yBOLW0j2r0F/hNf9t1MYnkB2MSVqT7Bg7JgWi0OPFV9LFFdNjLJFH+
Z0NEjWA81Mam721GHNYpCDq58G1J41t3A4qr/T1Zkq9P377xPXeORVqpQr+k
RdJ3kKzZaZuWAMKeKdcWGx7qU8OsIAueW5y5CYjCKUQ8N2LB5dZTQTwSAJsc
Vd1f/zHm3a6ABEM1PyQdjzTz+oAJRPOg/cy4Wdrq5f1cDu27sLrQqso21Jky
TxCjLgIC6wZJ06I4Ht9jwUvxjiCCFCjbrWx0nYPtsC4/Orpa8FdC86jttlyf
URYoGcb1npsV/bw4ieWWLgK/61h0jRGxexrM4yfibUrIJKNtUb8TnGeuB6F/
zUQu8bHs9eZU8DR5WkHZswo6tvvp7pIUKcIYh+kDdv/nL/lXE8lSsTP4BMls
YgXxtDWZFLEd2iSijznysT8OxRa4tcFmQbgr+kYDpva2/lK/l5EiGN03wrf9
w2fDwgKVXnZoq/E4HN7b2zrlJZd9l0Yil+fZOIUc5H+M90C57jrHvwbBRlQq
vy/IScd42PBHsPhJMQ/N/1yU/dv2XJ3A5r41WT4IXLExW6zP/03qFmUgPsrG
zlgNWq+uUmS+ETBJnd5qZKdquAxo5OZrG212IROCAu/XewxaVffyiA6pXlsl
NC6zyc1D1Y5l40swpNA5DzH5EAZHSGLhmQYa35bhx8IXi1Kwxsb+lJlbOgbE
tM8kv/Ev0RlfhJKbu8IaZSd15gaEQ77klsZJctibca4YS6pYn7QM+kq9Dthf
PdpGO1s+4gI1vN96TzPp9QpBXMf39yE64greN6BZHvJKG51lg/O5D7hhgsIG
xwA1PdmKGraupMrtL/wOhvgotQqTutW9EULVZNNmb5B7lKt1VyQsjh83V65A
T5ZHDQOh8sdWeEh+lbzq2fhLaK2MkOng1XmxCsp+zATChcXNUkMKfv6zmNv3
uCGaWldgIjXgSQC4qabOpmxov5OFAkjfj2KFHeleykvENZitQbCfuD3TE5xr
thB1EVAZPOZhMpUTy8KqhR0YyecLPqlld1IkYT081lTaehC5Ub332GvWbJ8S
feKH6wOF2ntDWtaKBf7W4qqTCFObY4xLEQgIqGqqsrw7yfICYyYOGD6/xnJ0
zmmhVvlpkRca2fTiAIXn2+gMWjwf6Otf/DZWmKmjLjjuHyUJ0cdUxdvZ5Fem
jkaFqutCL8DM+DNFLOo9satu9phFFDHpMVNT0T4K6aF5MHxMJOmO+CcIv2lC
X1sQYDzok48DCqoD+KNY3/eekxoT69rPhZJWc/ZYLdFaDY5CLPG2Fqqb6QPj
//RBuupCGexvwMCr4meW4vRhP0sqOZK4Nw5I+Kebnmgh3iW/8bdxSvmw37+h
Jmlrqxs3S/kABm02fPPoCXc9549SJmq3hEKP4nrx20tOVv91XOHjXQ4EGf9Z
4FilY5SIa6ifhPpHtcdUvKDXnH+eHkblGwvzGkbmXFb9QsvmAxHVjGrOOUxA
EhoRBJKOtA69YHPc7s7pmb46OTatGDEiuahIEuLHKVhZVJ/4H4iGIjIIEUIK
guLG71dgT9OS3tv6/rvBJhL7C9Tq4PSfsQeuUkGt/ZHJYWAdJNxwl4ozPZHj
H3crdWT7dwBcn5Il67HqruE1187T/Z0h1aRpwWgkd7LRyLyXasTTADDdLK9v
ir93fcZ3qq6dt2LGA2CiZJYV4/oS+pHvZh5AmyhD1DLE02LrhZgkUBxh/Ijp
IeuOCnfvVPxJiABjTKiLcBmP8Yk4H/CWSxBKjRQ0dOZQx28jFoZMcaPcs3OG
lzPNc19widefuOgmiXofqtAI+nTrNT5JnGKJ6dL9y52aKl8O8DRIKZuOfrZK
V12btdXptwFc52fDE/2cchpapNybv3VrZ29uq49dICNJITQvXqZRmWHPXi9R
UXpn+3sdXo+RHkxOyg3Lapzna2hymoPfPl5PQ1M2IMV+jf1hH578v5/b29KZ
yWCbL6zoNFoFKoo81rlZScUsABrbYU7kHBJMFDgSuJrNQTiyZlfb/5voeUMz
MQvquNxiq8CrbAB3aT91zTPAu3xNtanvio64raCqntXJ6oWbO30aBiVzgwq0
y5BwnoG2jUM2kdfJLotT5Psg58ySylnlDytaylhkbQnmIoX8EzuhIVueseHe
NpZLiBJcdV7YSwHx9Rwz+lrs7886IqJ2EVqb+9AKcPdrbTMWkaow8B7cBcKi
YBxvSnKNtYw/EyWv5gjNJQ5joDzMwvg7XE6icjaEgdqyt3PAkQBnTQ/jyUaU
ZSDAbBfdENldusC+6XZPtMoMqdarfnq4Lfxlp9kZPmS+PBZsao9Kg6FWpRj9
nmXrEkFRZh4P9QZQflEnfHoqGrqAHaKlAdQpVjnt+//vgYxtzqICn5Gky9QH
bVKdixFsRrh0hAB+g7j0v9xK3ju2yywANIfKsIV75SZ+kbi+IwYtc3psisWK
LSYV4/XmAsNlb0lfd+EMWD5mNQjiSJLNqvnUCxdCrElkucyxrlvB6syjoqs9
LCp0j26biuMedaEp9rPBnol7DzUAj3DVz1R0ZuXye7YPfrwYgx2d7B4ysbIh
PIinuxFh2mkFYoSvqUSIuODStXfx31CoQh4drm5kyYMRjgFvKjD9Hj6erHE/
Ezd8Wy3BOinaVKnqaSx83Sppo6c2LWQqMgXfqA8jbs9HMroHdCEo7GGxV8i8
E/dh6Gf8V8w/ABg+7CkMit7Fh1vct9spaPQXib3sHQpIhc7b0MBa5wk25R77
3LFpQRo4KgLU+ZbsV4H5/TiUVbbXHH2v9IbeCkmZOh7a6qHZThHjYAMbb0eh
AbUWwqrbLxQ5dP/W6CD4SnrMMKwlrhvULIykUS+6SnOIfE3rOkuYH0b9Vw1K
Im+/PMMsb7BWLt4QhstYpQrWDtOfNDFuwCWLJMm1LkP6a+gMeU/FwvrJ3xUC
am4cleZccDuxdsrV36d8l/40BnKCsWDm+PnOuqZtPYIBCbRyMICM2FIsbgSe
Ww/1JOJxjRwcZs8kfhd3Sp+2VzSOFdAEX/g15xqSRYklztu904Js3Snc7Arc
3YdK9KPRIQFMR4EUeTgZ9ygTqi3TqS9ZtFx8UR5f9ZTIv7bB4FJ27TPFMV1U
1N4W6Z7L86Jj0pH4uVX8baeLu2j0pPCgjk3ORMpkD6lcxae187jwVmzUdmTK
9MDoCke0rJmb7JlXj7CC8yIcSajgAENytEC2aK4UblOo/E5F7gW3PgwQz+Ld
fX6PSy9UlMbPSc5ysLrDwPvhqXK5ZniPrzkrq26igaXg1/ilo3l9GwkLvIgk
Ja/Mby9sy2LZ1pegn5QpCS0Ee1zg5zlPc+1T6Rizvyxr3hTB3ZbqqZVDwXoz
0u2atlhIJCmO9FzWE09lF3Q9rhaFEjVhjISHY/Wemt6HuAOgnG2ek+hTpIk5
LrFsGnlb3Y6oikTXq0lFJj4NjHb7stoYK3PgLX2G0/edvpwrz2njSa06zUvL
cqdindOsLFA/T9ALtxohv//5+qD2QtOVMKtn5yR3/zGVwpNx0mYE2Qnk7Gdf
1gvo/0Cjr0IpXp5VzbNBOjEExTPPMtXF5jIdEs23zrmN+/A1Fd1QiZ2Bs3Yh
JST6Qc+SWkbYZI3U2xcpt2dV0nbABntgTHVhNdVJhvExRfReKgMwbVoZHGwt
XFDMzmqa+JJtBSmXAV12E4nfFXJtAMIF9G6MljdGfhGt2YmeVUsx2RxU8v5O
q1u7lzh+YTr7AJSdzyMVA07nbSTex6tbRTA8tBTUhMa5EDipyLhgeZJ2hhP4
1FZeEnurzjXVQ+EJlwJgjpgxuIVjFCqu97qbHJJvfc7W7qi6e5E6jb7bhG+p
9uSuA0c9Z15+PTmYa38Y7Z2LM93XoBoj0MqVjYB7WKg3rIoSctchLTWORASL
bVA0XYTdJoGn/ZWhHZHHO6i4EqhbFawRWsE4vH5ifQLYrLJqq36mi37ImKEQ
u6fOlpASybpyKq0UshxfWAdyyvuoc9qJxjM7erde8HUD2x5OovaXKfg0Si/2
MdfC4jvbNWhNBhT5sDqGoo3yImB1rt2rC7ws2L+9T352jS8T752RH3riDqO/
3JQ6muC9c8Mr/iKqFH0+k1H4MzbbGmEr+QOgOVGvW2uTYCMPftaCt7YSMjq4
SyPRoENgh+x0mNkIOnMhncdbFM53+QQ8cQ8VIFwpfyvRdY3RzBj7qLAslEbw
mTayolyUWjJnyr10LeFp9hYdZsnkEZ7h+s2F2r9EOG8iBiUjKDJ1l+dieEiP
Jql64FysBQT/WQKOY+sDRsfdY6lvWovKeewhs6DZu+3T8I9T93MmyeQbm6YY
e0kKJknusFg47U6ryr8vxhp4Qu4oLEtOshqWp8+S7ke6A3ayz9amGuq0r8lJ
pPGE7Cpefe9S4dpuJbmwi1WCmnTKzd+xGi7I42gqKjNyTtnPy/Cn3X6GxXf7
rgRvopzpTYCctgT5Y3YIPKl0dC1719JPR3UnRTm2FHbycDXRepca+hV4iY1O
J25ntsAfC5Tdw21RmoB4RkZDXKLwpjawLxNVLDC8JRHBmPDxFykXocRkJS/Y
FFt4qWjfsILdLcEmc8w4VkeIS9OIE0+uxyZKeQejZkR1W7+PXPF2NG/bAKGs
akklBW/qYCtAA+nVWJ8nCczk7zGdKFSUXwAi7Uw5K9MI8rObx5AXlYkS2GR5
eaf6YAntf+pCmOGAVXIoxfmvLH+nIJMaID9URhC/QdjD/38ZEPoBUFEG7Phm
yt+8abaOE32j257HWo869fpCeQQY7uElhBhGhS2h1maEzDulVBqL4ux+6015
TGCjipvMwakU0Nzh1JJMoKHHYpBlZaXsjkqQBAZTxj6mkDGDj58Or/omg6AE
SiCHow+APWF/kLbCpnZGA8DNEuzM0t9vir/W7ZaHUVNtzGnfNSUxTo+2uRgK
Fl4gIqAnvzODGa3HjO6bxvdKlwKBh4+PdLHLXK1J1cO0u4DB0nKQ40CF8WSa
91EaOzH8K3jqtshWubsfXRaucgYoUTts8tgVNN+EFCaQxPsPS3rY0kOf6wuG
zSE7pU8hAdTZdHEjN8di6nXeK8c9aI8QuLHTNp4/wu6IngVU7goFiMZvNikh
4IerCsN/ftIdPFT/szk4VX/LnQ2uUDvXdu5Dce4DTUzLpfnwYRukfQGRAfAM
rtAaxnu0cwdMNnH8fXAyDzWOalXG60azT2o1ZgBM9aBcabUTgjU+PcZF3LTR
BcpdxVIkS27ZKmDJIy+iPAMMhSggoJ1+LxKC9rVQUllzUyBuPmQ/7qj2YEdj
CpWgj7MpU4WKwooApWXo6GNC6/hMviD9Yi5Jz/hwpewVr43TWrI5TIbL0MrY
8J7ZT5EU5Y1JAFnDq3Fzu9P3Ogtax0/kii6NrtQv3Y7OUlLVUX79nPtOYa4Z
U1f67ajJg4Qy8oV4P/5vRQvIolhmUktTMJ9LuDUvuiVduj2sB2HKZzN/RXsc
1H3H56XZSSfzGyOdV1sxM/4Qh0txQmsDhP0F67LC4SDALAtTY7wQw2om1USl
PJm6KbuuDA2ggGNASEhg+rlRwibAxmOK9fV6T+BDbdTCyCFmmLNrHIHXgeoG
Ksgyc93a6ZoDHd9hxrsZCNXj9pT1Kq9PsxnjELl1Np89Cf1c2ewhrtn5ZUhp
NEF6WgRScKuENb3pqG/RLik+PWl/DE3hJTAjrSYKU8c/zfAJc/b89bPQWy7p
qLeoVGwd5MUijDnGFyNsBrpGyZ4uKe0TVV8/WSb2a8wqCVYnb4SasXz0t9Q8
6xkwFgNnknR650fFz91TCl0MyE9a+yHtC54m8KkEhzzO4OmqVsgTpY29UgPl
q+WezEfPj57LTXGIhUi0DEUCSbK+gf5lJWcKIF3V45Og83Y5YfAa5dq2HOSm
6VNGunNOYcRQGH7sKeJUOLg0gfGhty5yIhtmsUGSNmzwbmV3T1nMJ3aiIuRO
fdLj4NSfRpVQSvan6JftjcYvcI2p0baS6n86TBgnDTAJoo85VhlCwdln9GVL
XxybMgnE4RT748oh9NnmvdcMii8DEroALIKOh22I19IC4lpVW4XunsZLeJo2
OLBdvTkJbtIOQmrmavfwchD8jGZmHP3v4yv8NXMhDydwwuFYvWulmGxrF8tR
So+3zPRK2CxhqGQbfsy46lq8cHVeQF/3I4caje1lQHlu5GVghcGNezsOcCOA
/6bWgS8K1aip1jiRFisqr7zwPDLlrcoJ+iVr8NFxD7ukMZnau+LafuB2PNO6
e8+xO0X7cbyKGZCdzhNIgn6bPIdyvVOE/mzA9+r07Y4hJsmXK234i3OL3IFP
L1zx+i8RmLv8Q5fETE+D4rTO3RFjkT47XTDLyqIAfJEWlrQLXWLCbwbe8M/r
1jsz4Qq7wKEs/3SqSWGA3btv/72kCFcoefuT8jCzwnLAZg+EOKqcAsg3DYVL
6ACE1pj3uapAXRByv1LJ9O2d7ltJY9gYGpCc+fYo0KDNf3BtvyY9qjKPgweH
g9BSoVgKxnqvSIQq+Uhbi/JUa/txB0ydRVUvdNgYAiKHqPyj/VSkY7OIQJIf
A/WKZtKHT+8v7u7UbtgwMm3OeZlzkxyJW93oLx4laZCj6yrL4UN7bUi8YZsJ
Nv2npa41clvXyIYNxiR4ULh+x747Bt3dd9PvIYjPxxlaABXM7qLCGk+0TTOR
LtXiytPGtuKx4vewhzNYu54t26fqpeWNH5FyaWcJO+bDS/x5XVIy1eiarPSw
UEbHHpFSwcmKLo0vz7QQHYm06pTW71XquWyGvXrw8at0ovaX13+xkVrzrIHM
qoyTXLG8hJl6eZKMpJHOqeJqsU/h3lCmaxgZj6sldhh94ztETzqbI90A6+7s
xpR53VHBsBv8EdBhvOWKeeICgtCu6mTBr8dBVdLs+Q0eB7CX60R2uGBMpjtX
5jyc0PxvVoS8Q0IImrrDMNhxCn2UEQuXld98Pw1ghDrQGbSoANsFLdAT1Imt
6Zjc5iPzljPeiUaROiFvZuIkdiJTeajfovBwUBPgHlp3U8yrFJMI/286f5Jx
W0RcrS0ElU0lBH9Rs4qLI8dNygbklzF39guM752DVV/yB/CFA77ZQ3JvWFLO
R1wq9MVUe4h5OQCaAmxqt+rX6yHV9QrOpx/wmXfNXkpGM+tm/Y+Oq7PdmPff
hZzZ/7MWzS0o3FRBjAq6pc00Y5hF6aXglWJ97XmWPYEnDuBLkP87jafk62zd
DJdERrMwMeGAMExyh6apAOEwvKoNG/VzuL51+0HGXL1GjCcoV1duwj/O8PFo
fvTQpLn8mD4LFch9GYMFVVRz1CsC1HMrAUtx+/cueGfw/pZ8O09wDBghbs7B
8qcNArV7DsMfpG/nKbS4tS4Ia6pYjt272CQ5Fgh+Uc3jL7QImKaAoYlWQqtc
tq6ys0wJcKCXWBZ3Jkjgungk7TEO6R+g2vv5waoc3Xr0sFX1EMqLOxj5QgkI
tvrtW8+40ksaCTU4uLJNrCyqZ5kdwNgrO3rbWXcGNR8xe5+jlRdU2yqXqIE0
U1zWaH8rtgTg+EwsLUEQZuf1qDZWVHP8KfGNcgdgYykOU6+t0pjRVaxssjuQ
KdJFjUyKt7W/Ehd8auzZa35nJ/Fw8PHxbQyfNLU5hi9ExYUORbaHo+LjgGvG
tpYRcf0e1Zw8+UGdzwJTDf49SSRyabokwVCU/ZlRqIGtBuWQdxDxiWKDspDq
ASmDoX0elaBNKIfWiUuinFT3+NtL4obbuMBz7HMrHLYyi3S/w3v+P+fBN+nF
CuXIM3UJum73+tuXwSNdo9I8zKNUiJ7gs34jmOfEij7cMLqnMn78tpjMPLYh
v+Eqyc7L4dCmG12mpPMW4qJB9syLKmVkN9w/1KaUCEo7D5IHOuetDKhYavjD
j58dTNXuPhMp9Ddy32gPNudKArFEdw9+b5kuLj48ZThbbcqprM2mXi0SzJY0
Unxs3XA0j9Bp+YqJUJYh3Yk+9Sk/9NWjQ5u++4iVnn4owgG/isn1dIjkG1Yg
CpaIaBwTJnR7dgsgblU533h0nlI0TtFu1X+zCc6EESVBVRSVKDr4d1IeiXFR
7dU/WTzbdW+4LUSKjGiDayFnoCOsW+MLvpGuMB4uxXrDv7egHu2t8PsZACSx
dY4qZ9lwEquAuwKL+dU+paRuUyibRPwEXFrVgJlbJnzEqtqZliqhxg1kAKNa
DUI0u5AT/d+pODbXJbWeXRiiUjzMjdcMQibW2qnfpl+cNdDRpH1vWwFgq4AR
IQ7Lfc9nmiu8WAkzqfRTmhId+Z+khOGGQZ3lN7TpQW3ef0EQ7nKtH2jcZF++
8X/S/pEgZV9yNEtXnTqTTQvWknMTOhbf/DmBXk2ix9ckl+Kmy3Gxlg5ovM3w
21mkkoEqvFX52QI0r3H95UIduEsBmjD5u4BLbDhZafUrOpzXIIPaLaqNeu3W
asod6n1fpVLa5mMZIhx8Eqp21hNQvOoN8AIZhiovp/a3L6mOl52v1Z69HaJi
wjwllXGuituVGwYnB0WawlKo8R00Z/goxO8jtW2b5SuKZvPM/42GPkBpXhjs
0df98MFqyrUTUxOkwhA4lG5G15JOpaGAs4CgYpnBfipRTTDr+nhSupNHGn9v
obBQKn3mu9C0A2hE88j7ykAhAswlZG3CStv+ZsNkIUzMrM93HsLZMcPiDsFq
7uSwLXLl+cpwAm7zVh+Y25l+wp4RYpr0h8pJ2HUAMeA/07KEFMuT97+MTeRx
RYQ07itictIKJbr9e9DcvSzr/hNCa9CJSGuWVTCZB7Y3xXs+TslFOHbxXRbV
ZMb+N4hjKw3y1bS2BictcOKiBOnWEu6I6j+U1SbT4dbdmYBpnABX1XAhQ/OB
+OPoTj87+3g797uadgDud68VGWrQI1TrKZwX9eAdeD0spJ/hnYLmP0LQvW7U
t/ONWQAt4nYxRZe/iMGrIQjCM3AtCpXB8eVkx2trgaMi2bkXuTXItWXjkxHN
AYsog7esEG2uyZVv1Zk0dG7PBEebLWs5z0nhqiWygyxpc6sh3tCqjeKQc/Fj
xsbzWmGkHUhl2ACOzl7WgyQFCcnra2Kcy1+S8EVDbpN6VeNxmyQV2OYurc+k
jdnI6P+F03MGFQhnv8dYL/i4PWKQL64QYaoXRy8h91b7uAcfTfyTvH3Z0jgs
M5Ca5fpZBUTL5OSrViPDemUqzkMbP0ZGL4RwDB8tXKJ8tVA2Ti66wTP9LHMg
Y0XRY0hw1clhxwaMADDE3Z9C9cy97S11veQQ+Etund+XTtO25fLrgYk/UeVu
pm8w+3HD2Qe4bS0CjyXiHkLw9aeaHaBvWRJQPtFs4fzVnyWOYLAPhWLeRjYt
1vVJlqCghIoTu3AL1wNezqMHE9/TQay7+5z2aD2KbGik6jc8lLHx5S3JVtfr
KdyXn4rrnhZTbv0DkXDbnlE91QhxBxUoIWJGnytdwfYgmDPdOJJitJ+K1ehj
xrTS+gjzK/2jMsV7lehPXol4Dy+i3ClE4sWdduDsZI22FaVh9KjHKKx0cU6I
KyujqwtSVLSgwEftukmrUYmuB7sRLHFg5a2rCtKWShmihvtlG17NRCh9LMZF
ywhuFzdWkUM+KzcwS4VlVKufQDVgjVBWqy4AE/fWx3CYPl/OsbOcddUWhiVm
4HeQQkLn+F7tAqGW65KjgYjzyfzElNFdN0Gvyc2RyrO6ODgNewOyZ09gWsUd
9AmrnppgG8faBC4un6YC5QycEOk4aMoeBIxPpM+Y6Uw7seD4GFP526au80gN
0m9oAt3HPU0pSmd9AeoMDtKDccEjPCxaVqRIVxvdicJczNITUleAHiUG6goK
uKrBn0h90/lhsLF6wQJiURvzLU2XFgSBdZFiTPeNIP+Jym8csJPQ0RJlWo6R
QYCnMzJYv9vE+Ypteph34wmcNWhdWykCW+hHAss6IwERjkZXmH1A4xe9mODN
CmQL7T8ar8ih5AdS1z0JsP8uUFlhmHUvkFqdGwiyhFN/hZmtiZJqBKkkxFBY
QvAQObWeLAN6VqtkTog1XFN2tT/YoaUvzLR6APE1mOmtgU9jXlJtCP06P4wp
Pmjg4kDFWjsZasIlHV5WpDmvedHYcWPQgt0mcLjcqRb/sxtsqamSlX+RTyP8
4nAf9Jqlc/NGQ6K29tsDEsWkCetRK7uksLnksB+5TxO0ZA/+vJBikJ3bTlS1
72qlKfNsteYCYmVvsoY1jNlICMJxqmmxhkX1bPVBL1/bI/m0Fi/TRdkUTFP7
ciuEadf12QKWWoGhwu36p7BeTZWSUABvs4ShSeftPa92Ks7X5pgBXjitTTaA
G45D0hvd+BBcgXXAqYTIPOa3CCy66Hv4fSBJlFPPnY0aJKDNgpqgH8jiAV4i
LcRiTHbIvqD56PFbz6zOAzRDpNgjwXoR2qCShxa+RUTjHFjDVcFHhp2ONJ7m
AR9B/VgpxlsCJeV8xp2vZdEFHuapTxrKmyGzR+rNEuwIrrbNmwrzx0DD3Y8q
vhoF7rr5douyYPYGimRHV20jaku4QnNMJr1PBorR6ID7I2ksCPdv55RnhpbT
4aiAHIYdWr8YTYW/KU5Ic+QaRyAn/NLdlA9K9XzVXIU3Sy0HBvH0hPXsnMGm
iYlfhRU/9vnsa72ln+1/fuIZt2OPif9o8VxI7m7o36XBnIZUsPlITtTpmPAV
UIoRq9QX2qpEVKnekiCOa2bGduJ86CFve9QRFEWkTToZsWzbInnE01gff+0n
7TCwd1xz5CPI0khviGQXMiMHnDzANbudVSXJ/J2F+r47QQLbDF4jnuDhriDx
79uDE1xF23VXyWhzP+EE4K+7cd9Tx0a3YzsFIjz08Wor3xsrxaZjf5r/GreO
c94lfByShaBPzwJakNKeYetyANwg+atQSL70aJMw7sItRPr2lt5ZMNqumDG+
F3dWbJ3tPAF2k+Yo2nEZvPw5Aa0ju27zPQEg+y0bRVkcCyY2UaUg9ryrkfpZ
isOEWLyCQ0E1ABFUQw59tWv362kX+cDTk7KuZo8KwhxxEicq7+KN6UD0YToZ
KbJh/UUZtFgzxy3PYZYtZJK1PAbFBbiPA5IpCYSNsVWv92xT9X9PbkUKiDM2
xlnJG46S6Ho6i3LWyC0UzdzjI/OyUuooytu0H8m6IRTqJ07Ahj0ygoBsyowC
6l4S5ENmU3yXKhVNvvXLZmTDlYfhsAB39t3f8FTHQUebOfVpDoOq6TxSuQvt
0A+gBHAa76AjRvhZRgjAvMZT6v/mCwxrxdd9p2F9fos+atiwAMFFn5eh70hK
bLxNoCJeCKptag6RIZiLi3eNcwRNdlcvS0mR13vfSupX9X/4290mLPdOVE1Q
MXmYlSEEJaeYMrMRz2kEVJGAyK6yd+tg7pz25zGswO4ZWkZ8u/c/zvCAZ+AR
aGsvQ+VE4vcCGbdGsOZNDd2slD4WzSduYKto1eCKEb2DsjZtmHRtsgErpFCx
z0T4Nb9GkeGNKWd04cCaarXLB7YM7isEzuO4kiYrKP+U++UwGgYW41wKOs0+
8DARtsBVKURk7b0g06xUgkaouJq+za0KqhYdeKdTMXOaIGgnRM8ZetNK/cOC
tr2PafRZTeMDZ6c6XOeXSGCSFcajJbc5PnKQubC11kXs1c9RSHz69vN6JUe2
ob9lPNqliaAcQJS8FgJfb8XVEqVwsgaVpup2Fm/zeH6M3GhS0V7rOQsHT1B2
QL9CLJxzPzCcx6V1g2bLzqi5F9SEVgdfp/nvou/sCbplJ4vNB5JAfD2NfvR4
sFZvbvFMy9xdt5s+/9BGBGxfjcQXcuFOsSFI28UZFp/7q5ERdZcqNFldIr2v
rfyvLBeT4Mb/84M+eZ9U2o7Mzo5YSnAAM/s0k/WQg4sIgRu/ZtctisFEY2An
NSOu/+SJX7BwHtvyBSSwDnG+FlY+Vtf2uriDMxSRkClfSAhwsKmU4NHSE04w
E+7vzYqJpdRmUmWr7TNPQnvYt6ERTFxL/x8hTrSIMpd9Qi3del8Df9irYW0Q
9NBi2oJu89PVHj7/H2+0kXg5sJUluf3HdS6y8yKDElSUXIlBgGS9K0floriE
XWmMMziMQzTWtDwtVXoo/41K8OjfMATiAa+kt7MuvTIeOT451nhU5Xx8sy+p
cFACCKTB1D8IAUeOw5HGNDfb9p2Af13cWduBZrctoNBcpG/drrOMLXInHD8g
mVIqf+OfllXcZWOl7E5MRNiQyKmnlHZ9O6fMS4NRDqju4bj0jUIqnvnqaeHG
ZdpnUf7TdY26YtKWRg8h1jf13niMd+vPOP16aB+UFsgJge41kjQyrpT7TiV9
mpUOdviFaOHrQo+9zG5TFh0xXEGScR6y5jLxMI6gzKDxFSk6nshjFJqYpYju
tv2nABwWhcIpMBLyYbD6Ovd3ngWspMWgS5tXCtq9EzgeAZcnPiTQNGj9qr9d
fnV5nzpNMkbepg4/FMIeKlCPIbNZcCgj1a29TasDhaBOnUQyjTs5DAInvVRq
0pJs05vNziMgUBiHzDUPBuP5z5el4sIa3Aw7yfqOwOTRsAW8jhv8GzZq8HvV
8DNnl98P7ZdQr3V/fVOqpahlBq5+QFwFKkfceWIA2vQszb0jA3zJDBsPmTEG
AoGFs3LGe1eBSSL8RKjgXlUEtn4LKZ9prONPaJpC0lnLVU8VIYUGW+13X4wx
G5iFHMMQGZFh51EqpDCLiLK/1ZpU3SPnz0FKa+1fpSNkYN30YPKZc/foSyCV
wNmNzwV/RrM5l7wI0NvysRL6VOwtetxPDz4dZgqSnN5+G16ofCYP8m6/kUpA
uI3uoTjf5SS6Qml1lzO/DcKqveNn0Ub63zcYhp5nkrvuJ+TmdB1e6BJ/qjQt
i10drxwcOj81GUNuHnGzOj6eULOFyP7IRttViRKiWm1gssU+jHY8yiwpe213
EC//prS0qno0uqrUGnVovOviiSPyzDTOhJc0xvyzcV+MVwQXYlyC7H284Cbv
0PP1MvXxD7Risf+dBlQGcZ4Tjve6lgyavs0ZSWsRljaa1w0CedJm13an1dm9
/JMY3GWlzl6EmCOLvYR61u4oQquTtC3OdQm8H+dJqPi2UMWWTgpq3yJGqIqL
UDq8oRTt3HRxXXJXdW3SyGalsoxwsFdUifqP9uH2h8YnDSvRv3Jd/PCRX/KJ
6l81SM8PXgOC4N1ASPz2Nc1Z5o6Q7WG4C0f0knYCLBC61Dy3KNuV8tYnbjCH
DOuXNeizEd1jb9dzQdBLbwRFXDN0g6aC1YGqDsSIYqnhpuUQz1vwaAf6Zd+i
ULVGAOSlZo2y0Fkt4bMB5IcEZnAV4/UP/kd14KeNGigFe2yC4oHiA0wTbENm
Zap821jEp7gqDgvp4puxykczHhifnv0M6B1agbqAF26iAeqV7vV6uD4c4Q5q
9ij4lRfcOD4SA0aRl+KngvTtOPywIVDMi2a1CeBQD3sq2mQM0ZFGopficKpD
Ms9IDDAEQb3qCTD28StWEosdHkyM8IQZaHfxw1bD+hMDpmEbHwqcwouj51Mq
TtvPtkWQdJjCgGfr/MlWOHWlX9MfZZ+w3ye1ZFRQOCTfOhl9fCKuaHKHAjQn
qR8AHOASM/CP7UV1t/GhVDznoS3j/cFXePjqsrXEN//qoLI4NJN3TmhEZkq9
tVHdkHsBwtOeaZhJ8FV5qoKhcEJYyZeecrAOTJmuR49JfW6BkcV+KfHLvdmr
mFsQVN2g3hiVZSUiiqsRgmi03NRoFMu/as3l9Sg9JRCZwv53T0dkCgPvdEDk
ua7y6PGJ82oDG3vfUK+nOkb/qBveW550HvNYy+k0/xJjhVBGH4X9rk1TaReL
bIKdvzo7xCAypSbowG5JDrl99kkICuGYfTGfXdCShL8pbuDiw3+pqLnJ1307
Tu1M3Qczzo7iNoIXKDtCZbiJvKp9NXesBb7O0qLtZR7kaFES0+ejOu2kU/UJ
/0WqGQXd+EvAry3TTVSSmoAlv6wxnBb6Wyf7tXdRvCylii1Nrjp5+zZbuHGE
Zesx9akmrANf5r6rVA87V8WyfMQgSrKamoNl4sc4kNuhdyiDLkd+crGpy1L0
Q5Hkb/9axLvoOiIv5Q6WEFtyXZsxjzISpPkj2WdH9g/NeHQXgkHBosF2cmu3
nvpKQFxlJN0ok5db5MnNI0bQzY+kIgChNJ1GyLQHeYjnkKd6hxmJGrlOws/l
9HcC46nFSKEdSfuJcgTL/ILQl3n4E8JxZ/fy2nOIQmixoapqAgNaU3Dpn1aR
OjGKZG2R+1bjDygwM5aU1yEu8uI/wu5NWsh0c4KA0T3aSuNZzwCqyNX8byPS
jkrkxJwYUsiXgsRTirzDEPTFksu+DfCGqQfAJbuLXbHlQCGBR1ia08YsCaN+
wGWlue6rKyVXQz6X5lzL4vBzlWbNHh+2cKd5W0OYN1KJj7HCTl/tNJe3YZt7
2gMnQlddiqSDk5eWseuXkJ4ON1/j1dGqqkLNRguuzRmmCYy5lHLqWWn4b6rN
D0HMjn9MnP+C42DQ420QkgAiazM/fsRoPScn3vUnYIWQMhB9rA7wj3D8HJKL
OpHUuDTmU3Mm+x3dopU+aVaGq9BtdzeaS90qn++6ZkOU2EH0fgL/WEDPbuli
771fPZhc2UbzmF3Kcl0m2KLy/VK6eUfZKOaaDDSig/ZXGAJ1Y/ZMRMxRlJd/
cIgDI40CgnHW+qDpKaRjrBmJwZv5RDpc6/yNljTdX0TNPXzY6wu9JeB3QThu
IIHcY6/x7uwTu6PUE9XW6JO7064KsW+tvZM365tYqeAfl9PqaoWIosWuwotR
XVjt5agKiyk/nIrVu+vWAukddPb8AwwXrp7tNxCFpLTsMqV1yRLdQ4lBkd7w
BDlSK5CGLvWOwbbigo0Y/hVM4XwDsQDakkzfwvxuLk+MiyVeTZFB1galc18J
skW9lke/ux0IalhUtfgILX7dZ2gRl0cXSx35huJbXT9sxqw26yFXLdek9oG/
v8l1Fc7fUGmeO5Qs07iRwQeiRMBqGGT1jui3CktFTfUzxPXdS9htlyzrLSQU
Q7cPIXbgvo4gPR7SIrzAKM+k6VFbe4A+nWYf/XIkm0rteYKU7OX91Sgj8j/i
qZ/yVTcgGNYHLn6TnyvBPo0nVhuo/Yki5pZpZiCU7xvCfu5z5diusiIBnukH
sftuML00yBwR6tdAe8zu+OsOlV/ISXS7L7QaF5PjD3Pa32LGQU/neb7K6bC+
QITFgd+8b0lUuyLV4XmlGIBMAwfQf6ctajv4p48VnEtp+aKaKHHrK96dG5od
nK5S0Kfkny92UDKHdfnpOMbS8ytBIfm8+3bLNZP7lfuJAE3HzgH/V5HRs4IH
wAWl5tlUzHAL15DNWbX9AiE+nR3SecSHUJM/TLK30Q2r5E2rj20Y/s2HZwGC
s1P1EiE8GBSCjPYM0NC8LS7ZmQZPKpCXpZdrPt6BdSEe+B5ifhKkcicBB2ib
7fz44UIXaJuWEZSRgLIc3D0U3wSXyu8xU1HaidmdsPPMYx2jbuKQRx4dWTs1
R4rNRNLehcoENRx/SVRcNgrW6I/1GL0/qz97ggBB2HUBmnxg/24+8W7Ps1Gq
E8CI2Tur8qayIv8d88qSMj5zLcrTTink7NhqzAnnRCrHbEllmcO3EHUjIK+o
oCioPE7QghK1H4Uy7CZd3iqdqqT5MazOGqC2gde1ktq+NOxdOwbnfTRDkuUi
huiR0k5V2lXrauP+XRUvT3Zu8u2SP8s8gUFIt6bPMkyeyw5k8dH5YZwGhQmQ
MjmE71EY/nEFzwgEKNmH/JXGv3QH1/1/2T30+D5y4oKqCINtQq66gb4g9INO
DPFL7TJGVeS9G0KGqpCdOIX+49s+e7RLVTtXyA41XRRGb3pKmrn0c2ip8/2s
iY62Jov38Ia1mW1A7fMddGkTYfwCwsKbNZ2u8E1qI4yvMC8V0KYsRXbwBoDq
vsgsL2uAaUnl0K/iUOj6DMF0B97G/Sbktlgrn21BW0tp4QPU93N7OsInmS9r
JP8BKX7xxya7BM3pE9teZCfHj5ZP1gt2jNFpmgKPGBwiAxzYQF64SuYKEbIb
WkVtJWVzoFOmKQTACkA8raFtzyXaA644btzRTeaME4+2FJyz0q/xL5+3YCy/
8JhLlwNhiQDwHtRQaIsbbZBfQUoH/WxRNVmVT8qYRU/1uLNDM7rE6KrrCF5G
Qac/fAcffvMfSDVlUpaSQvS9lXwl6ditXi43jyJBkyXuJJ5oXlaAgBjDVdxz
0zuo+lD72Y7Be7WBKe5Rpv8kbn5kzv8lrElHdRVfZ5Y+qZinHtlF31tK+fB1
LoXu2RKZmQXBtV8lAvJrVC1ynxXL1UzzYdo+aQ1MB+jTZrvqVKp09kOrgbR6
9nRvlcaPFEuH+o8x6poLC6bJpcSBaspIDGqRzi2RPWo06ErugzVdKWsvyOcs
+i7ch208AZlZxyut8FbvxYUDN31OogYxXw4tE3rA/jA5yLrdLgkVk+dJhmnC
atZQVKvJwOg5xcjq2cQiFmAWhe9MnM2cF0zeD5Tm2pTguq7DX1+jWHsVwcGo
qCzKIYEamntMq0wJvbuRZqQt3KS26AHgrXDRHIDPdO9LUJrqsrgQvXSgaF/K
s2QVS639fCSkL8D6EZ1OmGn3KhBSrT/iMjpAIS+ogVHCCXD2BizQ4bn6U2My
xJaqCf1gf+HjGwqmmhERTtbTBKX4WIJX7mjJP0wKiU0gyiw0f0tC4IPE7Xfz
Eq0gA+3TsILt/cPo3ubjm9eorxpTBlhnJCPwjMcy6dgGtsiO5qiCFv35OqDJ
zBoTfi5KL9UPT9AjJ+/gwjnPe35App+rdiEAV7jGwIzR5CMQOd4D/5IOuBUO
RgszSix5gfex49DN2pltiGXt3iO6mLRb8kHOR35LYkVOcWvBctP/kYg9KM6h
WFc1jTEt8zutJcXYFyfDKP+mfG+Ce/FXM7YtSpi/nCTGVqYc9ylo9G9UhHdA
1Qr6/priYhOhCb6Kbx26/iuELjGHRU9oVw/UNOz63qzBggsKo1ggVFPu05KP
ndNobjqww9MNjWFweHU4lZFbQZXaUjRQYD7nRk8/t9Y2smM69qxgPiTNt0QQ
CW2YSenn09jy9FTCF9FZvUC6SRZaqKwnY8KXJkswTw6Jqpr12dMSeXstg5XF
dG5coB54VKx58z29doJSy0x0ZCdrqLipLfP6ztrkM887CqRiGOkJw+rwVDqo
TBubwx+4Qa8iSwuvuyRIyJxMBIYmF3oPOiCXBGIRJI3k/+jXZPCJx7v5egD8
Sz3F1+JA7prSfevBtWihOkF5Mxchz95CzBPANpeXAFeoUe+p/3F3apPg5Zmp
PI5FG9BV/ww5opW0oyNMr8tsSM0M1bY2R3MN2E04apdhAxDB0Yg4+HkxMStn
XSqV2wRop6+Q4UpowkPdslIAXsYMESghqGw/3IaqYwWLa2Gb+vrAEcea8OCf
NL7ZxbiWia046xuzBr9U84Aoj9Bh4ojsIHM1s4a+5WyaY/RNxBKUjW3T5jMd
cpQc791oEBMSL1DgvViPg9clWRUZMRz8P2bdh8bWi4bUQIXCdbJjBOKgh2nG
83S1bHfOyBmqCrA8bdR/I/b8aPfFykhoQjmBEo/DTQjyq+dy2a0J2ezTqQgq
iJf3u4aGvmb2FqoC8pgW7vgHgNahPr7lzbFDHrh0Cj4eTf4DkfZjXOaoEhPh
kqLsbShakZEisnNPUMnnp1vzB5pTXgRdh7X02jNS9IbRO7WSpcmScei81eIy
XFOnnAV/xoGbQHyh2/CFuCVtsuwEXBv9lIHFJrhorCdetztpiHqIMHT2TfdH
xeOaVEPwUVGxqHgZ44DMvipzLvSoL6880jINiQ1ahnquDjrkOI4fG8HkZWJF
3UJP9MZdnnPCymmEOzKNENK0OBO+CmSq0FBHOjpkyRrz/n3mPEqYJun9wbtm
VIrVVWlCGb322cLlkdlSCB6zMIGfyXJyWciyrMVwMb/W0GRXHmWin7XW5tqO
YfIPIeQ0wPk/wUNRYsG5Sw8zUXTUBPbR/NZWVaoAAVRKSo7o7vsCAN3xgSsX
QjAFCrKXkSWZR+TwlhrXvie81/qMI49hBilLa44UUqt3PWjGRtewqMVWPdPN
rsbCggfW79VCURxcehYQBw2VqJlWMB+oC9/xKQn2RajDUBv+kUfIOQLf1qFJ
T2CU5bApbwyX/jWVCuKDlDztbLxL9egeUmRoIetGJ7QbMw9QDgq24vYM7Vuj
9HmkhjBADBu18f1qdZLp9vdyluide96C7ULTppcvCKua0o1ErWp73qMZnRcB
NMwm6T2wME0n9van/JHGHzLvTe+tLY4FLdzSsP9g680fHi5HIfh+rMP6GAuO
spni+378lSHU/e11NTt6o5eCI5iag96IA5amPaKonnc/BZXC5WMBkFXMEOuv
x+XpX9jhWXApj/7o02oszuc36haCTtLBbMabsp2+NU2jakxgjHu6FPexE2es
TjeMcU42b3Tp22AAm6k9ZgZgEpFX0G9IeF38r6ORibY+2UFYeTBro5thX6dG
Av77K3WuGnBgdJr5QnkVf+Y6WAKA1J9IZs/uGkpYqsHpWHlHnIZiSmQhoRUB
MmWLk9tkBTf+sSG40L8WtC6TSSQuDwfdCJh000YgACgO5c/Sot/4t/SEji04
ute7YNvfh700VK3U60xGWRxZHnScSpR+OH/qNyrn0HwX/ZZ/TQdewxzVt6gH
QgUG5crZQzOajE5TI0tymc4y0BLLftrgG5+gSdVIVcPhGQpw3sowTkBGgP0e
Q13ysIXEdaXO0rUmJuNlg8Lxt1BOa7MV4poicr6TdW0o9VlmlKcqiWS1m7PL
pMVoyR2XBwo7lctROLVvUq+jcoIaeJa66Eal13p5UWE/BbPtZWFBx3ZN3HLK
kwnpvGx4/5DTY2jlpSZowU93EUuruKbWxJI1ClDWDcL7CflphzHtIRyCyP4k
WsSi86TViaepKoODhvFdnI3KJFMcOB/iBnNY5FxxGlOw0YILIcEwDc8/GR6B
QHpfI5Jg1pQYc7YHXYYeoGgq/cwClT6lWqdhEzZ7T2Lb+J2HC+niWUEccxPV
UyBhlAkos004ptIns5Tea+KTE31/lP8GX5+kGnZglsOjasWOV5Vrgd8b6k41
y7K/WybRFVXye0xM2afEA49lQyp8WtZpI2gycAshRaUcYKpfkZfO63HyLKvL
Lej3lYkvF1yxBxL1wyg5w6pnaVkW9cjRjQcPX2wuCYRtaQEFdhb2HCGgQ4wC
TfE0JeFVVqubFS4ArmbVBZb2U+ZgigJfxHJcGV/pBSbEEo6fL0yPTtXK1ZLl
K7GuGGq2uvD2wIhlVcLccqp0w/bbCRykEO4h8lt9bI9tuDLFWQjvf0t2fRA8
9FwCWEdPtnHE8wpBZua60geqXxj5yGE+vsxAqIF0YFeEdlCWPAvFLOeXavej
gDcMEYkUEeAia80FetqJUKbABygoWlpUqLcU/VqvgT4LeERGSyMjBPn13hh1
xNwcSyD5xzvHRRM9E78GBagPs3v0S6bAMWNcvIzktkUvwWi4XL/5iZp91TdS
6Y2jieKtYGYEzfHgXpXkOBpXhtxdUs90FMQ1Tq+WvljyMK2KB8VLddyAo3LX
Aq+PMoMw0RC4Vp+IuDjGPS5AnHUge//ts12aMU0XedRQbrV2RneV/3/amxX+
ILpH6R3oZlbMEl+U2fzC8RtlYb5odI7N82GIJLy4qiWJ1/CUpmlRKA/Eveke
RgLn

`pragma protect end_protected
