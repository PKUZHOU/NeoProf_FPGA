// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
jHqbINCnA/RaJI7hiNr8DbgANchRD3Cg0jGIAc51yVjU2dVIWgjp/Acck4qqJiI3
hrJCkqeearEvvkLSZdI1RNmhyksEqM7tmlQsDUQYZJEf1A07Z3RwRhGJUdgYpSOw
10DumxSgGn5qfKuy22KIs9d3fWKBceJCRPvKrXjP3zc=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 1408 )
`pragma protect data_block
Xe1KJOIceF3IJFnKOSHz0Kzw7Va44Mouel1dT66+qfQT9c+hjn3G/bug4B7L6N9/
dSwe2uURQeSOWEEgX+JjY4r80HD9JYsrkruNQfPNLeQW7yyX/xF4MmNoeaMQ1cP6
/uUmYIejkYh2Jbh5KQz4ZQdaA1uLgQvLKLoIJkayHShM3Mp1Y9nV5o100zjj2Rg+
+tMHxn5N0ONcucp1rx6sYhqHIBbonIh2Hy9wgciG2M6MHUCwUqEwWo83XlgbEAvE
AMVsILGP7pCUf8WwtqGaTs9MWRSUTjzkvh3vlhMGwQv/NnUGPZmTc5HF01KLNalI
bZo914RNrrhnFLmGRHq0jrqWpMB+CfOnEVKL101RHPAUSxRu/4/SRITqn00/y3SU
qEyVYzSxoe+V/Qh7JdOSGFp+K/UHNtwftIfrO/i5oBULUUr+Hf2DnAiyocNUIu1K
Z11HjuoNCiLvydc9hoM8txRZ4a/h3gUMRrdvf1oss/BeJKrghDCcZn/8UYJZm/4V
AdigAs8jgWXRPFvU3IXkTTaZdltzK68jD/5gKqIMbgh59ZW7rTEKZQAvF5CRUkuF
A3kxvK9sQ5w0/9YFF77eI32Ek36IU1YQFVJkLYP5675yMS7t7usi6BRE54v8UJI6
+ajBHYx8e18NMIP0MNqcDQSIYjPhwmY1RtrhQQ2x5hZI3aP9H5CSa0mVaQ1lx1V/
YR78PjS6+Sq5h3ffBPw5WWubJnh6BWw2oOYi+11KjhEYStqsL7v5uKT6LK0csnLd
hqV8asAzQ2S1OQF1LxOIEA3jdZ7WZX+OHXxnJsBkDovSmLRFdYoij8Ok7htR5VHw
2tzM8Nq5bI8X+PM4BK+VFGDhSetAX0RPUkVO3KDsLqh/IoKpyeqrVPbNw4Eo4daQ
u4w5LeJst1LxoDetcTDUUiLKGt5oU57NRwtpnb/PR1Zr8OyvRwL4vQSqjrFow2ob
z1r41HVQz1sRD/6OsuuwpJNmiz3s1BL6Bda9FtPbBY3CCge9lSi8HUwfDftW/t/J
6WuEWArc8W7EL/k00M0PxU0RPtQ1T037Tw5X2d8zFqb+jJ7X57ILOCXtLyW99TAF
a6w6MNVMdh665GJMtTOeksqQ0Z6zI3xRRS0Y6jQGaG0J1s4Ju3HB6qTFLZR/kD3/
lOo5FCd/LFif6KsaFsrXM9x4evVqzGKRZzlPrTUrTjgBnFJwPcURIVAHlPbqSChi
m0o8lQ25xKRNOyBWp9wR4hHcvBJ0UgNnPyRzJxLcMnCVgHAoNUZIGwaatdMgwp73
avcxJHqYFfnUgx969aH8Ht3Yg3qwDo7Kk9KYsS0u7+Jzn7DJMoXsq+jPUuCXlYEv
7TZF3v/z5zTQYuC4ZWvrvYyc0WCs4tP6KQTURVaDxFAQUw+hLK4QRflubIPgeZ9F
jRqdkxeY7xvczMUp9b6JoLJzbzj8LKSUjjqd2h2c7uDJHNcN0AvbAk3351TXp2lv
LraPBflvJBjY2TakXGdBZPcsILhuXYRjO3D2tiPnEpJhn6RpGaPj4YshDOGE6gAy
C162Zll1kND43ooiu1xaFNqzin8VT9CFuZsYUAkc5AdQwmMVGbkTvKzPqZzIijHk
A4FiaEAuZKM1uYqYZ2wUmD8xq12JYgT1gwtnY8XlydBGswwK6bcSDDoTsZ41F0/M
LN8ztyIUQu8hqgWeB22eYgw0h1WkYTiktxs2eIq8Ma/1RcWnZdb3w8HG0nvUM9cU
BYBTh/d+SLL97u3MHoepR4Qjusr8o8JkTi27wSeOlpdgwlsZre6DMcC6KFRAH+ro
qa14xz6b6t/xS8doEv9Acridksxnzz33SqgRWWfNbhcRCkQnlWv6dg22z62wFCNC
C0Rs6TU038+FvPpImsJt8w==

`pragma protect end_protected
