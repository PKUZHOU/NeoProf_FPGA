// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
I9Ussi8KxcAZbfVCjIiB3d7Ywcq17Fa5XXdGde+V5Y63PTJY/bT75I9hlwDA
QcDN8lLZVaJuPAhF2rpaCiVMmAZAMxQUhL/3HNT0uCyZHcRZ1759hzMSIbUN
721vwtGlXy3EjJ9SNIyaZNEVHp08fbUZegulAPkuDLcKZPbAiQDzFmKeNnQ9
3ZvXrcd9zy22wHjU6UxMcq9KdReqZ1qTPVvE/dYrQ5Feoa06PdWoyV9tnlKt
tlgicqeCahVA1ihVrQ/fTv705l7aMK2ciU0YZZ9ddzGEoXqQe1+9M/WJK7Ik
kHdo1AADlRZSgtImXiCv2HIH63sb3iYHXsQ791b3ZA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
g9DPoT4y57EZ4/woaJsgB/xSMTZv96fsay079W89K9GPonb2Qd4F/dAF4VWt
BF37+9FRYkefy1ijM4QA/9v7eqHXhkfQx8a6ssz4EiBGf4GlW20wjw3iYMM3
LBRCY7Bt6zGrxmaOIdr06BmsShQ7MykZdsSF7FKjdP9KpIrblHwx0E+RtCe+
vh0rY68yOzF9HDOVQT1UsAVrozGQYcs0JkeHslZ5TsqYYHMo3d0T3B+lUHUV
rx6WQqdP21sT4WDd4z1y8S+05zUhsw2ruxtGnhzUmGDsp2sV4UpVpONwSGxy
2ReIos0K1/pWRdGyGSrOpYXmjIZSNuyqjscw+iwyvQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
rey06nHxFEKoV4E+JxWmYKdRUjL2jYFd5qyUqq5mK9Bbq5+dG4Xrk5Ag6fa8
a+sl1g5jgeH/bt9sKPyVY++XXDTj/iqpnsY9IE4dezzvC5UHsz9T1YyEm/Pk
bR8tsswBU+qos2Q7Z77Eu9TlpVCjfwC9zO64mjvo6VVR6K/fEmVfmMVG5IHX
+13HP73mBuawn0aLWXhEBMkwigvGkFhpgMTuZUrkByOfBSV2eEdRrzNC+CrZ
4wuK3KBBz7r1z9PYDLqshLa11WHldPYnu+ZF1TrFsbdCtBSuJ9JcrikeD91M
NwoTAOpN15eAGyYTx2M6iyGgA44w4ZH+HYF7pE1wMg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Y6X1op5l0vcozkKSyUzHrXilKEwzoMcgjZSaDTxo/f4u8GxHzpCsTur/16F+
9J+xseyGyTNFEUdaJOgHNwRP1aJjz4D3BMPDrp43cFQ0ofGXPLtVCCBGLOzy
t4AtU41aB49qPJX959ariM6wyShIDYltH8p5pkrQMj+WGRdofAY=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
oSlyzmI9c6SKkwkuuXvPDVyOQuIs6mpnNguEvUoEGfM8pTNhlOyF6wmBs5ia
E88DaiNzCQIMyqgsnG4Xw4x9HT6iydf+UgsfRc5jOvHojCcuWTG7No+A/Sd4
SnLuoWhv88jPOekS803qVbcRvCR+pTH/qty9e0nJ2rgko40J1oQkRIPjWzHT
Aw7NaXTenedEg9FWwAiTMevurWfFWqdx8vEWD8ifzf78WHQ1zayzb5dB1+Sh
gtMiVkP3ACYfLCxZnTfltKZoM3k51PZmTaPtS9iWVoddLVxPWXL3H/d4DHdF
LX2RTJMxoJxSiH1qK2TLJWAb3Dga5aQGYnykijZFzDuZGLaaZU6DnrD0Zzaj
1yXaTx4xO8imYAIjXxsqPipUyIhvgq0t9IPbCCBb2Or69p0ax3qIYOWcec0L
D0Jq41pxOr3cE7ako5pMnbBgfG/r9yLbDuZpirr9ebttRku+E/rkAg+2DdH/
pyeEP4Auta+rKS0t39EUJAN/RSD2XL3z


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
JPle+EKoM+iuks3t6gpRXqahgEbTe6tnIorwyVeF8AreVFQGPn5WCKG/XvFz
NxYbQSZqUadATl42DUK/uM6J35sQVOSruLRplUFd3fQySfhI7qLPk667eUws
bO3vI0FfHzl2Rx+kWKgAuvVRXCEDx+6WyYTAkBrqExp/uyCZgtQ=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
qN1LkMtrop82ud3RsP2RMyi21AyyohCL/9PqrU5Vq7O3MZMVFVrsfQPbzvj+
sVZM4/4E3DgroPcsDY7+XTG+z3dxnVr4ObWzpKd1KoaNdNyLtva51RKa3Ql5
hhxvxuiFodRxO2IcTwgNW/nHrk28kkbDUz7y5epuwqeqDtDFfo4=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 56928)
`pragma protect data_block
Y8q7RA7iEZQe+eM/C0CwERsjs1Kxe+AEjUc+6uClYgacyIJuQ6W0yTaqPCdO
hFxv2B/1aVKD3JeJfY64pGg53xbQ9rl87DnVJzKYL8C6MIzDdDlzEc0o2OsA
1Tfk2mQ9u/SzXMYk6vyyUJw61MuHU2AGuu2KcG8O9gpqdy4G+k4reNtoQJYS
ux7kMF4KTi6wEBRjFaXwSXCFtBi0xPfF6yvagN+OPkPJrxb+2UrYDLUDOAI6
M7aCDmFkZPaKvMyx88AWEQnMXQz83ResZrVtLtAH+3ziV4TqZ6RJezi541iG
Eik8C40roH2WRMrl38WO/S9qY+9F/0vRRHZhmZvOTN17ocpccbeeWYJ8m9pz
oce+zV/hAD0PxjgvjTXkiPTVbWrUu78VHBSZDGOvsPPz+ppD4+MyhoqhJUeT
SP+KhZBh4yf+3rhIxPnRb2vo6Eh++SmZxPX4XjDiQva70GtaV8rM4bBgDrdr
GL7dUTZMb4RsE6HUVku34TEi7AXalvvZAvBFtnwp5gzbTQ7SCXFt/yvtTwMt
nrHfz2wJ4Onh1lb+N4F5AmgDP2aFC5NlFTUD5HH2hCPg67516C2DTX1+LIzp
hr8U3wPC6FZcrN63WlHL8zxH2Ztwd/Dp2gwHw60peS63wqx/n7BMStMYA4Yj
YU6/9FWfoZ0uJmrnjnybfaDznkILvnpVy/Aqf8jF5/njmDE2WlQ4+XyxMs81
Ct+1G9/7O05YUAG6ZwiyCAgQa4z8oIAXzJ5EGp92LuUnZi/7vSz8zy6gEGeM
anLWw9N33KEELVdEiPggiUb+JsFWMYe6eBWOHjEROl1F5HYjkPBLeQTD3e3n
LSmOgf2YwTBoS7DkgGX5B82SLjqdchVStdBh47MLMGBmmxR7k2J+kr/nwAhx
jy/38odLke0rxjO/F4kxu9oHORbw8MEsQ4Z2J/JGz0FSjp0Y8YmYF/ZHjtpM
7dzw61JjUyuwGDZ+C9v8ebfezMaL6ZYJOI9dacMvA952NRp9oGTX6RdOp2WZ
JZ40UHmyaTDWEQQMhjsSB4/0QC6xtjDSbY1U3oqzrFPBwm35Quoadnbf3UOL
XWSvFZ9+kMEMX1r9ygYApjWO1hPkRE5cEDcezoFFR86Uy+N74uiDg2KSd+Ef
tSYrjBo8QGXMjWaTvUMEbnqbjOBWDTTwcg7lJV+DKt8qbyVhotgisVZP+X3d
6VRQCPLu5AKtVG6/TegoeNEGnLwt1dExhZ1SwWD/kT7NpFLXvCBqSx3zgm5w
WPhwSPmQeZstgONrJ3cPEkgwTNV4rh8u098q2ZHkzx6i3rGTnZPTFBKz7WuR
lkvWosHhs0+4I5JZgG+aIk2qi8QTPfeE3owS78bcRbfTN/HGoaWfoxYYp/W2
bp1ha3edCwyd5n5Vt/BvTBKjl9PNSFZYhipy2AlUrfr6cceoR4W6mvh2GI02
hs+45//ApK98/yofQP3MgDC9XzeJoAEd8kFjkEjuHkLXRh7GWQvYayGxQOAy
WtDNKHQCJiZHUjNX4pW/D7xjR6XOJszG2PlZbZ8wHK7KO/Z7MnEMXAH9rJrr
4mMkcLwejjquBBorxftloEBuOq619MKsmxNuPkX9vGDeZG9D3zJeZpuuWG52
K5XFAwFneJD5xpsu0Be3fAc23tGH1wXBnznqx1Yabu7xn0IWNyOTfqDsLG+J
a17J2Fb5W9UuAG4OVo8lC3JVPPID46ZQeOtV5E0NSxWbukD4/kACpteWP6JR
FdEvEEWSTgFiscgc+S+ZU7B2+8dW22XYZbDqvYN6tGzHnuXhnQkJON5u56JA
BUBW6r9JH3rbnRWq8PAggm2s+5nFRYd2srWs6Ioa0sAH5Hae1UuUtOfomhT7
isgBKhTLH3cAnLTMJ7NzuegRQZ7HOPw/xJ7FZpkvKOOqKaJwXojWr1/xLWEN
715LJu5bQWs7mXYoiY71w1JevltBSq3wFv3UDlJWKlJP/6cTqnSE43cNlx1P
DXNNpFhMj/lk0wpILPX6WIy68j95yvoJzBkSm7j/BuHjaIne2lG4cPTuwvYF
+HeKwo+gd46XIDd5gDkzGtL5PxfGsEHHOKtsBHq1cwj90svpmMivpou/X1X6
huwyR4JfZO+GHtOipxfBWEAGgELDVPXxTBWPuEX6WKyoNgXlE1A2IX/ZB6mY
rpRPNAIDlkYNy3rexGUcLBEPjFo2vFk1vlVGvzy/nweb/kwsAFALN/ii9hQS
isYWKduGOsNYk7Q8cvSORUisV4coWSOuP2NsFJABKSszSxAJ2ZFmnXciWZBk
gpZqD0GRdSK6afmY/Mt9rIqqEo5Dp4WqndSs37ORGXrTtCBfl9xYEJCeZxlb
kRENAEP1WU+CclPcSw8Z0o4r/y2fx72X6B2zFg8Ncqd7ga5E/RFjTK996N5k
j9i+25Y0aaE/brX9ui1FGJNOtKM4RfVZ5zZDNIbxXgkEKDPXhx43KfFHAUz+
mPLB4Re4dD/fuNV8ilQkLJSQ2ZJi1YJr/TiSC3TFYXImZtRe8au6Gbzc92BP
VpkUsD66Uc2ZsQscTIW08+ovW6dmvI8jA8nTEkNQeCrZW7kEKMCD1jxu2IeT
grlWWqnlYYd3GgxllpiAozgOQUMcsrKIpKvPdaBN+aMQ9XaYfV7neXcmm8nk
UyrB8xvV9PT2QVVhBOYQ1N9KY3L4zO8wFIWcn0xLcEaZ10CXnaFWu8Xk3yEy
xrlWKQAJccRw7g4qNXhaIoPyhMATIA1s9XqDHTkKVRKPfsP7ux74MTvHwXzP
2fegoMGFUroQ97iVJ9K5ijsrLH11dygEzqfMjbd9OLZmeAeZUPtMdqS0uZsu
ONRJMPUkHgjdgdozT4RdlunwmLz6x/F3z3/wvByPX+eNX8aWV1kuoUB5Xga7
IN9cIe6fTFM0ju0Cd9tXT9mZdkSf8kSYHgTGIOpTkzocH7xDLyf/wYQPZZ6H
2BvzbD4ZnuPtstbEBOC1MscBHKbYofUWfWWLi3k87iuhv62joovgw57Fli6F
AEmFYVkphZUBimrZeVdJmPJDjJzfIjorkW4zHmEWyeRXzL4sXtzwDcp/r1J0
MImeOJe/nJ/B7d+NPhg7H0RwyESTVaUqdnKMB/1l0Rq9UZUNvb+p1vRIqWCL
g09sc8V8A1kznf6nCd1J4jQDqy4vTu0liOni179gt7faNSySGapKtQdIUDIw
dQ1O0qkYiFMGtfFrkF0COxgpHIQTlfm53aB/YU8IC60NIOnjPG8fyEivw3wP
qSYhKVvZ7AkVY8u8D1dGw4Oaw+A/GUb3la6FWVdOWzmD3NAeBuWHacLzQKkX
WBjWN0CU/TX9zYltQTmLXoFsEnMh2sv8R9nsypMMBt1PGEjTBego/v/GG9C2
j7dkpqkgg33H94A+QicSNZxa04wvQyDgSTRbBNTUFBHMraBLJAGQth8metbF
6xfRnBj7KuxwsfZWsUQtFO5MH8azoQoqJBSZzqk6f0YXeDQU90NVEuf6tMir
Jtnz/a+vReyWFD1Tlt5Bj060q0iPH2oVVRRsaWp2camLBbSRh39YbZmHuyEs
gNSGGR8l93CqIyTJWuq27HwgWiSeobyifmyftlH8tKFA0tINuLSQRUlBKTTl
h+Z2IufA0qLPkqMMwYF0TcLaAz3QRhuMrdq0GO/6QgiH/AKlBDS5jrcC4Da9
A5HPiHUCZzEXj0CrPm1mAtEM/Xtei5m/+pbx11H4HRRWRdRHNaxkByspmv/M
YfCyU2QbuoP2t1i1eaIIOs1SlH10VgqeSBrnCYjQuCU63fNoRsOeyGwzMWXv
Z/7jm1WQr1ZVxiK4sQg0XMvNnyZY582p5jlTLw+DFyIyawMU+Y0v1osCvETW
75lq/65FYV7xDtmuCtKg2Syr4i3pM4xgdDmaXeU4PyR+8BC1aszKoyFjuKwO
RyQr3ovJordWyn8UBwaFIDKeDvLxkfMzE/Imn1qDgjc+lQbD0yYP57sJRk0+
tj2WhVAdIWw3Urv1fkGORnGcseqoSsBSnIysNg0FjteZY5LK9kyqMg5yikRN
pzJbMcXCJNh3361EEgGmdppltIlBdBithhbIvBoYsQAaQGCDCUeDXLBFNC8p
vchgJpffmVkVBYNDaoUlM5aCs5WwY5nG12mhVzEJW1LFJJRMNWcurAzeXPBa
jLLKHcQuSqksacPub2Yt0t8b5tSSZE3cHYa+FdaFOrRVAO29kMDxjSPDDjdc
kM76B1RJKRzRehBzm9NVe33WTsXG24pOFGKf9JLz2hoJql0/lhHk+KNJI4MA
T0+sagY5GCjgv+7WEJU0UbK3jQ4DJPqydP4GMXSAsYR9gmmh0XxPZprvhKw8
W8/Dy5dWpZ56UfD7TqNKni6254HuM5GL8fmdxwMz2BsYClL+QD50oKMK8fx5
uHBGuxc47sqHrSvhfBzIKF6JoZnKxaGBQ2R13Fyxx8XHRGuns/N0SaYBWAa1
NyM/FP7SXKTDsOlT23iTe1vfjGM/Fqy+SNynU90MXifs47P5s7UV5ZbJ2R9Z
0u4KnQiUTBZ4/P3gRXSMa+8czBh7OFFDwefKq5lx5U9B9h8dVHuYTwbxAOM6
rTgTU8hyI6tCGpLit5WcVzgR0k01jKpvcOYAwXO6o5p56iWpGMAdhxkY2qol
v9bmURHkz0k4aE4BpIcLEDbCQoiJu+E4vQEVC6wdxz8Be5/jB++/5GGkGBxQ
+ENcQZaMjEo+49N2VeGRhdXsZJA/mm0YGDFYCV3tPThfFk0ooqNE5LBH7Erh
v+S4zn5HaJ4PVqlK01eKVFZcEDspeyRTPrEoHFOpTQKpfAvnDg5+LJ8/ebyK
fLkdJa1Ia5qQaJscYRFR7ryNe8C9CIfPuK+YrQymcNaQVuRrnufegS/pCWKy
RgybpKAkkf+KqgHN5HRp56mi/2F0karmNwD8CLygBlTI9zraC0UmixRVRszz
2Bi5jQVHRhB6LMC1Vh5hzLLlMC+00SDr3o8niCj1x4qFdyqJo1jSsXypwAK6
zrkMPURi7QS0PPJ1S0dJKEpjuLQuueW1aufRdVQEhxUVTD0R26+EM52eWwnS
g1USGRHLogatyFEKNXR4/QIBHOTcllM2ENNKeEau2kn//8qkOqGri2ui/nDt
lMuKR7c/6OrPslFzIwQWoEOIU/fc7gjWQPMXhpommw+IVBMc9v4F4oyEvpsS
JTdty0KgnqwmESXHPaDVCPmAxMJeAleNc9j5Y1GtaQMnw3PVZOQU4Hcl9FhY
Xe0OmuqtqK6Vi3/5PB3sDOsRyoQUwzmy6Mvck7K7wPpxQ2jGIcmJ3mCb4S8i
I7EC3os1pqbdD2rlX83pj147CNOPdD4xNraorxTs/OD+iflfeegCH+0OU8nk
M8HlcX+b0BJ23vG9SNHDVWFnQGgypoCSzOApknXFTMnaWfYa5V0XNvh1kk2X
XNoGYfO3keDindOI3gBX9o/pyISDN9+zrSBgriY7k37irqf7JZjYuSDXqx4a
8uLE3linIQMYFuT1cjTMXaNdQQxeaj2+kOJ5/dmIhsuZbah+I7uBQdNH8/yr
Bat8jQzXLKc7PYa2D7h0rWNqnu71dwQpcf66auFLhsqdIAqiqxQUD9J7LzUH
p9xho6iqUin8BXqJBO4dbeJB3RMQKgoADvCfSfkgyx/p2zzhKCvH/z6z5z3z
LIHlhiDUBeo4wz+KvmJq4xiUlZMlFuAalN3KLKBtWpDjn1vBolHdgZU6m2oa
59kRmcclRN4UDjsiFb/VZZkBM8MfhG6auTfT2Hq5uB2LYVlYoWpqoPAaWmBb
Djb6qk+032e/8WzyuMxMs5uPBTy4dRocciQyMzFg0CCMKD8h2jtCP28qD5XG
0ywzYY0miBFcFi6+rT+OE9MgIjzZuh8WFIydxMSFUHLWQrY1JibSwIRdV4bv
f/3CFJPvQmITWRrnNxIjNZASXGxubLwY38bXF+Ohu9yv0ELEO/pJshBd33rO
YZM0/C2TOQ8I1wcXc78Mh9Rr8Qffpt2nzBn179EfuNKe911E7A3wHXA08S0z
b6rycLU9a+wwYzXf9/Qa3dDv/wOOqQz9gwDUNqaEg9FZCH3z2R57h6rYYo+h
prtjkrdWh7lKIQr2G5mZVPJrg9jnNc/TH6QxI1n/oDEOqrB4haxjMHhNHiBV
7Hk1vVFxSUzpWJ+siAKoKexN3Y5v9HKesJltyJe2ev51ymSJjh7rH4usxt0s
vAw7uRVveiN7iIiPikfkDdwJFXf+aBMwydFNBut2K9OEe/1MHS6XF9aHubzM
MjekXzhsafOTrbmryeiUP1xjHDIwEjgT9/0kr5xB+SjxxEhEPqPFdypPO5Rv
jgn6WjB9sguTnDdZ4avXwSrZ1UgElJtYYi4WIq7pzR39mTpEULfMlkKiggOy
f+KeNZ8pGzweQF2uaSNaOfleMzKuJTx6cDEW/nEUSjguj2HSyFxdS3AFo1FF
h+XKGwSmQEvqQvAEPXyoojpMSFKxX8Qd18j3A4WjNIQIgHcNIVeepqyQurhb
xN2gpuKGzJhv9Ja4H9RilAn0mNuzOztBuRog6JLWdIaBwyxg3vTrMQWlw9GJ
1yiWyJ+EHDfx1Gz+25ytr3/wl7np7EpPmBwL8mmS/oK/NwfAcptxtHknW5mb
Ww0oUz8WKhMh7yGFJr6WD5F6qwaXZ1+ra/D9Rdg4lEWn9WMhi04lxokVRVvT
T9q6xtQFwvrETKZCKCD5rZBQA/1SPr3KJw+73cpX/T/SNyHRWUrwXM3ok9tl
N9gw4xpiQ/E0VtPTDyBRdJXCC5C0eBhdKdRSp7C5zhmVhjuVvhU0OAOX8K5V
4KUo2KKjsEi8yY66b8R5Irngqco95JC6TNrltQWnXZMBjfd45PYsQZJMqAqU
tm5a84m+Jh4f/ClSqDp/f1OeBiUWDhOcM5E+4mRQJwCM/DkyQbe0+vbjXiQa
KmXqdQ3BAVvWe1d/TjdS3Oz7n/UbnMfXHb9d6OthXmnUar4cVVSxgXrUA8EY
7HLqdO3x12dcf2IdiSdJy9lFhpZpgEco9PKoBNGlvJ22hj6kJ4J/BLz16E9c
CMD5omeXMWOuwSppTECNs/bzhS4d/f86gmQCMo7gPjWrTFCttzmRsYrSocQY
3FXq06d+YsyECmxTM5K1njzN5BXrW8wUlMF81C6u1QwxVA1qp4gbuXGUIfTF
AeZYQbzYRNSlJb0xt4U8SAJp/jP0YfJRVXHZ9ucBgFOKG6zBTfMrI06nplZT
t8+/jwFTFRA8JnKIdNo+lRrFmYrBIbXIdvfgb57hrfmAKsKOVpSuXXoxj+kX
Y2yoVpP4nNkRpuik8k7SB2oildOXpeDBq4JY0yCrcybokx8hwvHjeGX8zidv
J7aACpmWf3lOl+OjIF1gv2mbLchlujCbPlPll6EMmXxjFarCwi2NfdBme/tk
oHCVQrUL120ulU0a3A35cZ5Wz0ixoKiK94TL0qSs+OMoNpTb+OBdG2rPzNER
BMr2eCqOl0VSgKDAV3DVhKS91ica0bsroThE3eNHq/say4Bb91ANigaEChnv
e5TNru1/NR/1AdL1iNkP/ff09VvXCGkBq+HVYj+Yda9BD6+1/ciI1MDIB3sb
I7SgA+I6NzABXqCNOdRONd3PcTuOw4jK8QrKGjx2ACh+L6UD5p3Ep9MgDFYY
9TJB5BMZ/yrTV0M3u+O8ms+LFKYYA6x8VQG64nPyUKkni8uB+Zof/zUF3I+Y
v44WvcuvxvheOCZIuLrNM1lfb5370RMllr7PzFG8WOleXe/06KSpLoq3vm/W
wiQn5t6mTXJneluNhZL21Op6lQ8q7c90+9bp6bDec0oqpRGVpYUn0mSBHd+X
cfhhV6iH3Y6Af2h/aB6yt4nz/Mf0H54pf6QuCEa7rHR9USVDkZTLz1FQUFGl
pBPiUHyEK3zgIrb46do4C59EdyHAcft4qVf48is+sWP4h5ZRfE9pjjv4hRLq
2kIcvRqXPhgvuvlP+XS1AO3leujVvd8i8diLcoOlcGP4sk1AfbY6KHv15+9E
AqXD5Kx7uC6IcL9+gVG4luEleeZ8PfkcWifG0t33dCq08/qs9zHtqoR4f03A
CtLWvNIcOpkmAY9Iqq3r9Vp4adILYv/WXZ8f5/K8RLvITnhFXzeLHnmAnTIR
guHBKvxO7eqN2uhbYNUdCoGdaMiBzedUUijyr16c5EY+yvSbvQxUCImYZClM
3SbDIZujA/dUPNkHYkcLHY7OdDmkDm5qCslQL7TxewgBVIcO/gDs3N2ow3Hy
zowB4m2wgmWP5ErQpBmVQsvEgMirZhV/BwN+psUBsnZjIQ4Bp+eKbDJ2f3a0
O0rxpS/1iFZUwpHDGCSDNSizJS2fhxW1/+cwCrQhLO3svuzI9/kgDhQkbboy
j0haR0umzafN/TP1YBtgL1D1z5w0f7qT1sMyhu/QZkhzN8/BC6t0vfxRNIXy
VWBKPG+C2lnOGalXooiugnrUDSZkxa4NJp8oL1K6iRz/yfKzb9PnY0B6KuoR
dbOS6OnUG8OznnBnX0coYZfObNci1F4Ompo6bPc1r8eAQ71Yv9mH88710qJ/
6421OzRGXVCJ06nbcqqB/TTeqekbsnEy1ZgMmQqSmaM6sBF3BmlkyAY2i0sm
vaz5OU3zbcWNnCaJm2s+VXznE1/Oyu5Ki8xVTDnqT3vuyPOJgKMr7jycYG0b
+IDy9Qzgza2CaqbG/9beRDbKEYa++KwAzwZxufdgXJhtjGBZ/f8zdDK6/wZH
MA81ECzZHORjeGUFKLMCqN751UKa0XQIiZ+0ZgdSxdm6ir5Me3mOCojCwOy0
BTsbsZkIxoPSjNxvulm2w55Pd0M6GkTQ38Xo8weTRVOtCPVltJaKnLQLB5jr
4xUwERV0d1sdPqiqs/n0iVoUXmv+JDNM5SEgGfDTUzZcitiuQ0nO/snyzAcE
Lj6KiWARH/1eGwHyLLjC87VGjMhqq4wjES1O6ZFqYnIFqfpoVUgdEt5BK890
Q7Ei7qkwhEwBtckAte9IbIBepLlGmupPSx9cmkoMxfT3nFsdGrGWD21O7lti
HL0h2La/dRCAB2QxS5/yb6hnVg8CifHUfJQwOKBs+4FD+AlyymIry0T7Sf0i
06sP8XMDr8XmxCkIwossAJDqKd/DijcT9acnE/yP2wzHaJ5ZVI1QDybLJzmc
V6XLdWjgIl2ibr5mP9wXIRz2l5dYkFdVi9sOgiWQP78TSPWJcjc1ipa4WXuq
BpshSAwwtD/Q9qb+dFwAa4XoELficVxrkv3wBJIurekXZyiU8DTCmglNtj3e
oo8Prx206fLP5i7sv3rC40VccfDgpOn6EpS9m+PBOslC+XRDpb2CqpWFQEgL
LzwZkaXzm4+D72c4vOPd74KjSJG/aqwjtCV1eKmWii9qRHLtfB5/e3+gdGFX
xC3SAODVdlEx/j/RSkTrOL5rP+Eqiwj1YDJJmBlt0J3+RVVXU0JUXq542yfy
+p4/chd6PQba5HtcCBH442/4PhaSWAyLVJpJLe2mXI8rRE8pjFdFIWgEVoa0
hkURYJ4EFtwjmm5BzZbUhVsXRNvOWFRrL5l5Hn9/Yi7B0dyceitQiy2rJay6
JromcOt4OsFBOGeBvPjs0thFLEatnoiK74RKVrOxzMu9I5sLOhMxD9oHWwp1
CkyUmDvNZavG3VUMI2eAQFieo1LVTFTdKpC1EUmX6Z+YpjkqihbhNTxD4aRy
SDjA0bjddzdeiumBV40DCGRmPoMNqjQTUVKnZ39UxRNszzi+LmDt8BOXFD8l
bA6UnwKDv+BcuQsWUtcIN0UYg3IMojescIpWlCIRx+Etf4rtEl3FkPZ7ivTC
XLst6MqE0Py8HAKIm0AH4vdx6M2+KRyaIL5MLY+irIJPyrxXFMNS9RR0PlKU
OU2IM9LNfzvSNyahdQIWiutND04CSqfYHUVU8GloLZfZPuKTt6yMdq9eneso
cXtuI3SdLvITndetO520U2Q+xDqFAT/YRIdDoHi6VhvdVYbtytHR8s9k1XbD
2eB8wTnKLLnlNgzVkvtEUZF8fPv5DTFTL7KmpMXAaq6b6xTW35VlHq9yic6c
2OhIay1sbSayx6ymI/hMmzAYDyenWwCkKrZ2j1xtz68Vo/HXm1YHlxvXqqOm
gvJPt4A42xAFcNkgdM1ApQpkBhaRJb3JIXfJcQfVZH4j0o4V2F+qFvNDNchR
kBzQyPRgDMaKoNm9b3995UM3lqFjSGm6YaQd7YdDE0PPDM96lPdXogvg2rxG
sDQShBvXJXAeC3cdig4tzT+PrkW1pHiMD8CJYuZYDGnICH4weDKkH+QcZuTs
pyM0AYTi+s/UoqOgrcjSKjIthinlf7O4TXpySC4B5IVFvqTQ7xsFTY+RSsgV
Emkv1/I8TE1DviOer/SInqX7CTlO2hli8Tlr6jI2/7xAv0AfT+1tZwL4j5/u
tHAD/tmtefHUKvlyP2WyNgzFr7yanuLbTpmBACPsTU0OonriyHdgvqIioxBP
gj84ohydY80JTuRs7ooLSPHCMTBCTiF3+Cvs00lmNVqd5BzgZ2QcxX5SoF/d
BezN6/2c5twoyJipNE7pxUOWr2vs3kjOeown4+MgFDiPKk/pkEgott5ILvyu
XlalgTz/MTokqrNGl1nblVchC+IoF28zKzTOEC+7mx+LeXq209ZBYR4Fe+Ps
pfJHK9JMNfk5PfSFFac2fCsZhy51EUu+VAO0lI4hlrO1k8ZpdoLDFAmXiDI6
qsUd0Ir9VuZUUxBjg1+oCNvvVz9uxD/5AXZv2k0Nks0eNsD1R/x6eL6bqDZn
0ut1fxESlT5ic79tBa1/WHmOgD0xwHHVod0NJOESFV7b+YoZbiaQsHMVK8em
eQ2QHqSMIe4YVuxczn16lDoTgy95VCvPBuCd6ANRZ2XaKL1QhowDSnvF2h5G
CREi0Rzc0BxtCi7jXj+Ucevvfv7a8V7+VjWGvpm9/ObzOeQ4GXItTrDTVi01
4+BvzqjWcunLV4OUIkzUdj6M0Tsqvr6QQb7kt3jubcT9cmxCy38HtjAAhMUW
Hzc/QmjmZp7XQq9sxlrbzDlaObRMGUfG3aRlkFtvO+Ysb0Uvt/UfN0HAMp/L
4fnB4OJi2skAf+MxSsJYTiyJBH1H2ZF7NNke923bJ+b2LXXudr9Yu1lhrGwe
AoTmbuRauFI8X/KF7U0dDTfli7r41DKu5AytZPDhTEt8TK1SuWb5+64kH3ra
YwP38gna7Q+gX/bB3czOzjAp6xO/F4GMUswRVrEyclzat2+KJffqyB1X4Ix7
GEUgPvuwLHveyAI3k49FGRpkbF2GyOGYY5tgQV7Wr/TCTmt3EaC0x7Kmq20i
ZQiE22ybIsrBE3EwLBugtai9cr6pRXynGaNbjRXn8rKhS2KqXS9rMuCK3rEs
I8XKHyxMT5jQDH6Tj3nn/bQG8zKtPkYw81+BUBfn179qx1QsiNjKIZaN0tky
Uy+tGjoTPBg9G9t+wX68c/Z/v7k7vZeo/sMfIPKPQtFV8TS/sijNJmzWPLFQ
FLKDQ57eI1FtT04R41+F9Mvq0sp9+stvWOxRWhtMHKEQc3AJMDPdkJMd3PUs
cDv4vZeU2yZ4NfMjgj1oaixYnkX4K6jHdo+X1NxBpvcRiZe3HRDDKaW3XJjH
jJD2j9m5F4+zU9CKuBL0BF8zMC/ZY60ekt+nYBjUTTLDAxJmZ0yiYlOe/xGL
/lcS9CVIECIjwAiG7wPU7whNKYTjeuSycC6T1xgcOYJUbj+HHhH0V1ai1Iv5
jlk1cN6LaoJOSHrOmqQvRoJ9SXuJBP+BdwyEQCNjTXEZSw4eg0OVPU9u4XYS
eZT0zwY8Lyvsasq4QK0/zd/beSgGhkSTySsmUZxVuiolrOWHImUeCXWUpyrT
XaiipvwoKJY9AQlG7yxH5e+ZKAzncG2o2nHr/rXXFG4sAnvRRZn8Hf74dXu7
zrYx5N3Y/iyvd0hZRRQ97LVIsLN6O1X0R2BSTAnYQr/buvRPwBsuTZsf8eLt
bJlR+ijW9OdFQEWBEvJwqKXOSXSb5gXBw5sAXM553DXqYQNLgzxtnWQUuj6X
r5HnxhOxld63YZkt0LslfP9eUnJT0NdL0vLxHjPn1mS9ApVLtqLaMNfBxn93
R8pbTkJK47jEt8fDKLQvJQ/MlDxhbkUNY/oB5uZHCffuGDJJMuvdVoAsta5n
44r2gBqn6x8lnD9RbNPISqWaXhCefYbTSnw463Y+JslU6gqUjBQb/iTvXIQZ
yNEB0t8QN6sTGdt9J/3p0ZV1YGipDJ6ybZlZ7dPWaVgxaF6KcpnOUphNO2YG
hrW4F3IOSx9k8bIIcyZ6ip94y6UbSn1DQvV3mUGRNFZ0wAiuFaKnqJU+QJ1u
uK/jFYXja3dmkkgeQz01ESwL6EMmzjEyyvJZmPIrP60OllGdC59dVPg8aQ8t
RXdBoDzI8FyQB9VpqRHeSPvHxPd/xR3VUE+Z2y43ou1P1MKp27efXtIvTlFx
54qGTxtuoRaqEbHiQws7tzfcNMSHFnpSDek92qRStxlvDbNZ1DQU+e/ZlUon
sraRKSUHatztH2+JnBS/2iuH/OnTayTy0wcsP6VduWqyDxzxbf/4YmAdet22
jz8/GaPGgoWwe0r6UvgrZZXzzBM+LFD/jFl9xZqM3txb0ujfqX9SZhaeuqj3
KOR+Rrg4w1C8XstKHHPFQIVm5SlUTF50w98+GduspiUrRfvsX4BejK6Wl6c+
9PSNOyKvDOv3QRvpU7R3dtwuj9Sjf1MOHi16cjdQ9rB+wFo+QFjcDCuVXiG2
39CK3lMRrKdEGR+AXqB+/2T/Pb7BRi+2ZwFbkQ046zHJZVmbL+9N2tGIkU5J
4VnntDqmviGnnMsvN+dxvARdA00iWOh/qvvMi1KrFNrDUmJ/W+dC42sBUJ7E
5mkpU3wvjDKRJ9eDZMT9MiDFmg7ui3vYR+HpovsGCEFFLnJtDfnXZN9DzNdo
C3uB1G8qgY3SaZDad2kBRjRcHiWO7zwNenV7oVybyIVujzP1WmTQO7MMTy0f
ECop6yhQNaYJCFxyt1vqbjGMLH5vRq4grDo/eHK6Fd/XUVWp6z0FihXGdg0J
GWos268gfDrrjzLHnRohiRsINxIs3howxoVSB7Iret/EMNXnRUe0QKy163KT
g9A31P19EdGPyNsWaF6aJ8fkC1K0Ye85iXxCj+yrVzwXfKe0/6F68V2ZUf31
bizxeFfEluN5b3o1/kxsIJtrCibstmnVtEvR6d5lL4bQXvad2MlfmVX9KvGk
douK2yfd8bNLZmgHJg/Fw/fo8FYkisPYTS0+aTew+wQIzJ07iZiFlwE7xIwH
r0HJV+vxenZ5nknep82XfMcEZWzuS3ZAp4/3Or7qkEBTAMy47oCv3O+40sYP
EK9J7wGtMPOxh3r/ST3buQcsJ8gFe6jwT4lEiOyjZ00KuTVOO/ruExFkc1qj
lCgk9BwzFbH2cLBJ8ffLoN3gwcQbG+QQCmQvi2pT5+Z8F4y9bQd+Bnf/DtO5
2Dq3Zz4T2Njd7gf5e1+KLitJPWFMIVWv0sz8T06BwkKe8LUeXwz1u5BbpIX9
fyYcFRa9G6czXJ4AvFogqGRGKcTbpKKzI+S2CYn6e1rTqhoOb2oiR91rwcjy
JR+h2yVKN3oRt9mf33vi7kq94h/eW4KpFcL60m5NSIDXyraTBltL0viAIYR7
QudTBiQul7R6K06HHgfVGE18Yk4OdL8u5hJlS5lLRGFjRb7ab39WV5cw2jly
X803ftXWMTW0P1Xsl5vqwU2JBuX1Q9ssNmIkJt2rlPrSuSw/dBqF7c2KX+t1
Jep+jPELGG0xFzkpGrYsxVv4xOk4OTw+TZZWr1hrR8ZN6jTTBauD4O4IKlVC
Z1qzXxCWMrUGeDNot2lFpu227z9J0t/eRljTt9sk28TJo9+zkrGeEaJYOQbc
fjoqjyXePgFLvBBKn3851Sxutv+koYWLhfU554LsrJGJ5oBnLlUVJN2A2mG8
YbTGBy8kqYm+UzYK351u7BMTd6RZ+Y0M9+tj3gStuCLYGU6TT8paTDiVQi8y
Lx4y40cCB2LMBCznBB2R9ShJ2kUxiGSC4448CueHZVmDqq3i+jrqhL//ta/y
adAx5dWh1L5pUMO0z+GW3N5rf2tk1LT5f4+DkBlF+XXcyBalFaWiXbNaPgpm
9ocW96e+UdKl3t6TQggsbvNctEOS6Dv2gxea7Yw/z/Df411n8kVeVjuvPU94
GjE97H+f82qAdnZTmxkwrnMBTXZesJ9waqeqy4Silg9r6hbY6NkGj8mw8wW9
vKAN0Qc61LD4Tri+hFKmcHQaWirmGnm4Fori/JAlFQxYGHb71oHoNR8h5pC+
mN7ruXontyxROx+TeC6YbOkHiCv41etv2vC5EfOlcDU5aXrpLGxdk4BYiSlB
8oTP6J9fT7DJRIlBj0MFw+K/KdmoE/L3qQcm1nXDGRkmh2Yv7/PNx+ehIJZv
Ula6QWG0kMhVtZZx1a7fn1++PSqWfvVpio7MMNDh9/kQe9HZjhXSsf/ALubj
uH1ioH546wkG6CnfT8Ii3Dlx9//wTDC/3zSSOedAr0Aa7F47sjl4KsturtuN
YYJjVy/0MTSIVJyvblUnEG/ezrSCXbdE9QeLRltUxnKFabZmRRwLG/A6BqGr
lLzgFxgVJZov0wKuqcvr4MR2CcBtyMmvCUnoRfhpWzQ1kKyfOere00XaxuqR
KtTsgVIBcKBbdeKFqi/xZFCuODW7TnFshp/uNaoTCubd9sbBkS9C5kxwCH9Y
Yi6gY+XCIbvtb44u5wTus8rxQh4d03UqegVwWjNmvBKmJ8rk8zzZRTY7VCZk
smF5EenawnV8ATkwb2G8g4Iyos6uscUiE4sYHu1q+zYEu7OQl8bNdBPh7bKO
A/7VOjKiWzX53DiU45ZdGy9Zvh38qQgLu9L/Olc1P6v1tw2NK9axcrtH4XkI
Sy5svBED8tTMFlawKIwfjMKXGXfRKpRFCW08USZF+cL9EpWmpcs9iFBtnFAb
XPBAq4+1egqEum5w/LehZPQPVD97wCZJxFBe000vNGLRcTWK3DrByh3MobsK
1p4B1zzP3KQ+F7y1oJaRPZ0Nfm1W/65rryuych1ueRhR2TFRR1EawjlLPtqN
I1PBESgJyH+SNc9HUYkBZuQLjG+P68WjNM2Oe2OoVwln/z+HTroW+zV1khTI
ZMeh5UxoPPJ94jixPdUcdQU9QPPWGvSk6v3uvjtp8E549H+RNLnQPLdww4c8
kos6Aga0SqwBv5FYOrv2ofIrTagx66Az5DtUMEhVnhtj9x+w7ZWmT2T834Qu
7dHfp777mrY3tWUN3t1I3oOEXRaJ0tmiBUS7H5t+PIxNQLj+rUBaOXvP2e12
/gVR1u4QWZ0umlmRGK6rziZYRU5ZZW8go42+E11TCGiha9VH+p1+SVej3nhc
TR5S8NMqA/DIusV1+1PYiEs8RBarCrt7US4AcAx3Gq2/J6SKGvkC+fhP5Oq+
tiQDgdShn7Gun3hleG+J1xsaZsB1FCVl27LGN/1naxrALrETp79aMlLMXnB8
G+EZAn4bbQZjfII6w1x1p0Ki0XDEGExeeLrx2WjJIGRg6JTxaypB5pb+keIc
FH4mzTtC6K1BuJAEokD6Ktl2Qqv24NRTRaO5FjFB06SnNCaXxVjGaNo6ejLL
xxGcFaAqh+LR/RnzXqzXaLPaIAlMNJy6k8eGQ+IAv2fvjO15Lthw8f1X85Ep
fju6ltz9wvhikiy3Nh7eBOo/gOOMhf/ji7sgZhuxhVg94v7I0Xi609WH/9ND
fxV9jTze1b3eGLIXrsWT4LJ/ayzIuKWiYudvJhanwI1+TIkx4Fjww4kC7Uj7
pJ85hhmPjLHSPueDpdRGrspp3T2UO+irfAlaL8xlUJ2BUe8E+1kecoUCLmDs
SnoJ5I7nDjVIOMOqBr150LIYLwqSkYhA74e2jDIodRhdNodnGVIIV6atjXnz
s99tBE5jzfDMKk024aBlqPPKzOCz5lUN9AsKNSxLeeARM+AntrtwhzS2wMIF
gVU1aBdBOMmX9LHNvBjz7FYGJQjYJEfmtX2ghE94hr2o5oGahjW87wp78gsV
Mjo0Aj/LK+6P3rN30zNm9zgwG89HxfqlBeVo7pY/hVR1EPgFw28vVYrXELJS
Oo5cJXiWX+46AZMu7+Bl1eA39NZUmt9lBvC4lvQRQI68wMP2sOGjIEw/9vu+
wT7C/QLQRIGm6+uihv7RiVma8i9joX+9VVlpZb0S4z+gjggLQ3QibvfoZ5st
FJX8pulN7kU2MPI5it9U+vVmv5trOCR8sPchxNhSPPCs6Rtx0EhMkua4RpQ+
+qk+7/0XVyAX6TN3vwt8Gjx763OlnT9fHGMwYHe+yUlLX/O/MTQNTOZwE3nU
liCoWG7KzW/xDd3VV3GA0xhUkWO8UURsSIHHHFsZWN3XcAnqMjTpkB56+26/
UwtDXqsnkhbzlPwxRS12twtnTxiVUiwGrBmK3P+shXKmHqn6XK48OyTPzx75
Ry2I3eXq/3nwB6QJxqSfhxm6sUzCXynlRLAWrLjeLHqEA9GkKox9e8MzL9WJ
XYxRzROZ/cfe7ADD//Q/HrD6tUB4MV6d+SBG1I2cw+f1TEVdBi69gn+lNpXd
SEixLJxa2XPCY9ccMHgiNZ/B+htH+M83ox8RoWtdB9VoYE/tdtwqmQBY8j1H
HNYYBcgvePxljiXleQ2fZPLbYRftYd7iTKpFx45kAgjhxCsdZ/9zul557Pvt
bZTc9Yv9sCI+hK5va/lbXCQfzfhNzNIzmJb+JtWmLXOKO/Rfb1sqXbSVqagR
Xn6/j76e1vsenHNiN0U82VgSLK/SLa6KbuF2iEoJOD8K/LXT0dqN76mNTHZC
U/wvEYCQ7T9hEB8FdpScGTgaC2eW6LSZwrKfc5gX+1P9u67pWU3whTxfqzx/
9QpSdq2tpEQiPAVFlJsgkvOC7awy8JH2pEdiMkmdfZO/pza04gdDzDwegNQz
tOF6momZramVN8KNsdr3+1MugfIH5zWx29+EFcbG6bfZUHd2SqaL2fRcwHWC
3pz+I1ns4BCuJq8v/PLMwqlq9t6nGpB1ykLAIcLh8wDS+H5Nu4PCGAVgSvH4
mS6rTdXdYDzGuEAoHSCzBB4dePIqdYtbL4l14SzJ3+WX48Jbk9VnDYgfezJd
+ht6IRn3j9i6teEh0B1JS1Rp7yxPbjnWID6zainEkkwwiURYed8oH3JjxA9r
+Rcwdjy5DHyPcahA0bTdPg5TdDg+pLxrKEGbjX6vkNqptFtv92Z3Wf8O+scl
GwDQiQdDkARCY7NOgPzlCD6F2/4utZz8Xd4BqxX7n779r0AZ6GXtQ3k1MgwR
E9/G5aw+dH1WoLQFWng53xinQ5a/CB7uPpEkb1I7QGmeBec/f3JplWH5nfR2
nQxZdsnx8d7uOE2MUGoxAP+1dt8Ch2IpZdk3txgqdG/5703wrytWtPpXMn0w
j3T0SpKx+wk5M2DO3LEDDhp05RiJbZWm54FSnmzMBpN9XL32v7LRT1WrSdg7
g5MXvDjCjvEZ/O1AskIJlyRTZflrMZTmewEeZMW78PY53sBgsIRr9vINU2rt
F2sUY2X0Vj3sZwNU+KGkHKNR+kFg/twVsNp1ZMqshE7A1b1YfufZ4xs/kbgE
E/sGVGMda3jmJk8N3bzJmH/ST1CVv/dzfhw/sBy/aP4YGDBr3c0BGhLuruo3
abjDfcdh5KDPx7Dz06qYU9cxtJDJfs6znyRK3aTQlmsgaouIkXsEeiAPSRxh
4fACxbvvJEBdsbuvPvC4Da7LEZSvOR3oVnHh7to9Xpn1Va+tRRSZUdPw9vXy
sGJY6IhNgS7l1HpW8/wojOKrZ/Da+QIdyf4Q2me8QDz6iPDOAk8fO7Rxq/Gx
dh0YQs0IQPcL8h/9r60WEJamF6VAdu52d4fyCiUE5x3eO9F9Pru/WvVSrGjE
+pA0Sg9lMSeEythcgFxDC3n1AzNH+FzuSlOKlhsMvgdsUqfxBM8xkLk6YFZH
3w5dRQ5Fdqdozl04mJEN49znAphlNLuHpuOlDzqQymuKSnQlC5g+lSuEAwlW
oHYxbgX1AL429v0kK4WH0pSRFO7YhUTP6GLny9EkPz3ap1BhpGjzGBB5Qf8z
D9XRuGrBw123n+zYBt3yvW9zCISBekQeA7SQEA8ZZyMugkSo6aCfV+detTAT
ENVSjGLMX5qE21n/PyD8DuXiDTaJzvQSmk2jHTKO9nDRB1YqcjvixIjQOZLT
iak9IJrE2Xod74SO6SOJglPyvb/IvURwu8bL9wChsU/SuG1sMkHlOd8odlem
zr9z/kaiBBowe0sKT9S0paK9ZxmjiuHF42bIfCP4LGi89CfaoON0yfNQxVkn
9h1nTouoGOhilINx+HIWUfMmmAfZw10U0K1OwDXbBLz6i06FOEKE6qTXMnuI
bQSl7hanOorlJsRA4WJ8sgnmUJCcfMNYvwGp/AKyBVODW49A/lw4gdo2VVgn
DvryHcriOGxBLYNwvJTnCxj3dojMlxUtey68srCtHcaSYiO110lRQbCwohD1
MJz6JUmn4j+mjt3zFESiq5HnwE4atJEN0VG65FQCti8+tTEFnZjYFfi9fVpM
tE2JH4OvxxeTs90X1BFoInN68hIhFBwn22sc+qnhI170ecSzYbIQ2lepafAP
xLkxLpSZFteE60PF6p6XtS/m/ElfuHyO9hKaSi4FWD/fgtPgWDjijAAEqLDg
y8lRqkn+azxlOoErOzIbUMwKmELiiMEX3/zYAx7Gwcnys5y/WXoz+AZ7TZFm
ZaTOAHq/CZkN9HWcsCH1imuRUo7O2LkIocLl1nYtkT8lhhQQ/CmMGPhMO02B
kiu9v/JT+n4Iyo7H08dKubItuxxeyPehch3MXflBYJ5MW6R2eCP++YnrgzDb
+q4nAAaAK7JRMb5Vvya5Y6sviI/o1SbK5yndP54yLMjol//Z+ZRXbKCHVGe1
NwH6QXf1jo2Yaqjjo2gRYDHJQkAzcmm3s/issRZMI8wIex8VbcVHsFKS8z1a
skY85Wypx2qUdqZDwJpuWrnMbp/qEtVU+x9cjgVPqR7duQTnDjbH4cOm49IH
8UjfLdIikvlRC3skqAankufA4J1vmkMLNh62Oib89slr2tzY4L4kAL6RirQK
WdXMiGi37cT+z/6eupygA2dfuOiRFYShpM2hW9GZ0VmQynP+b5Iap8o9aYWv
RxqeAKf0GfJ+puWzg4xH9FHh87JFvy+vdLMBJGG9mBomWGVuhV2bqPDtaSuG
7SDDTZsGFmwNEOBF1WnJCtgnfzlvei7y7EPjSPhmuynxeZhSEuvk2NfedTSY
nFdQY0RkuJHG0ssJjXFlFg2EFPQKrRuLJYh/jzHhEWom2mOaqL7Pw+8xhRMM
nSg/QUZzM79dkY9o2NzPHldcv/2QCzwsbw7tfmd331xtNFtaB4XEzLQ8KJn4
pKtVd/3DBryQVtlZ75mgRFgX/jQ0HcBoRqKnSon+5gQcP75PHOmEAqmexu6u
hjsDeF17ZTjhIvwqigTBTyexEe23jpeKEt+/pQ++gTQfOmTstG129/ImvWNI
h4tQrbPnsKaTpGJ7SP+NuS2+Ffqj59t1sWbE2O/G4JzNkgXfmoGXeW5NZPXo
YuZMgvtiN8OMsdIkHblXoYZWl3yL6XlUP0mbsfQJZI5A5ecSe8oGQKoqRl7G
y/VytD5k7Oo2zfpO2hvAqeXwZt4gTlAIIQy6IwX54MWodeuOWMO7+FsxesTw
sL708obegKwcRYbRNsMImQpO5JcbQP8d3vakpbLok5A0uH/bvGqFLQATpxlK
NNi3TWOMsxTVGjmIYUNWrh+nyNH91ynivfcpdpKXj0ecIeaupZr21E/P5iQ/
e9Ikyv7fL3Dto/+OCTd5UnKuu0q+3D5o0oVDK62l5w+izEbkUIGVTZCOL6WH
BGbZkYRffNqVFJK+vvqhmf4GYQep7RgzdZh1EnvnivQbM0SK3DnCXLjfaiC2
7M0lfZLr1mzrd6IrE4ShHqqTVMLrWrE0gTenCjK9Rfu289KCYBGAkrEaamLS
Ytq0B6YcFmYyXu7Sq033eB9ZWyfitTYpotbcuZ0gaz0WbGH+ZllIkKdCnPMD
jgUsYr9jlOMPCdRDsuFftx+VeQmLBA8qEEzpnX5MYxbIXm75xWF9aufawP+a
HALyOU1vTYkLnCSKPSik1hyG2I8rZyg3Fu4CmpVvfSyfDVZj/45E0iFww+W8
yaAaF716WdgpkBC/k4NqDmiLqile7HgSn7Jjeu73gQhydvXDZCtN1dQIEG5g
yRQGenFKZTV4RMoaB77tK4csyz97v4GRf90nv3y1BlwFqUnCEyX3KCssKg71
1+4IM8yPwO5XmvdhRbFRIBmJkrT+RtsTtBRoFIXSGmosXH4iE1jaXGnnunVu
Swvr4nt5sazq4Vwf+Vn6BETmNZ/w/EWMdJNkAhSOOTRq1wh1EQ+DrijPd4C0
aiUp9H4lUg8eAQpPI2JOtoo3pOXzmVFdoc5e8Tirq7l6BnjqECk/EQxV9TaN
UBZR65hrti2gw5z/wyOFpRQLXK7FgUJck/kRmtjdRLabzq6Yyrof6H9R6GBT
nf5YKLOWSNeJOpbf3OFRZ2z3DXwrGX6R3sT9ephDACrTTjrxVGwnX/+SQb8P
6XhhZXTOd0YaK59mDQ8EsIRotyi0i1imkSkGMmfCfumiDjRaOQAR+0pD8nZP
DvgHqek7b0iWdVpRPWl7tvLNG8wknfcdQExbMQHsRo5VUDp8gFI34z2QrePV
rJGegScW6WrRnGQCUbyMecqcOY3airyOn81XyUwUjmbE1QTeZpqj1b4mHPLo
Z/cKGWMjd5HgQyii/O0OxkAvPAGwgI7kJJXoSmqhYXfT0SzIe5mdgwgOIv5e
JPBFq3ojr7rbIPBuiFgaYhbtpKP9uaQvpL0QkOq2KNNRFzSGrk6ee26t3Wi7
unZx78+Z8RqA0AeRqVDg/HowJU3Wj4LKYTkADlRqFdaoEOsQhJ3y8KtlaRpW
whVV8Zzb/cUUEGB8/zgpetvo0bLtpjIPsJocOmv31kHkFxSFgV4vRs0O1trl
SKVdQ8zvJNDuju8g6UsCu4bqGhQdk2LtmZRW9GsbIY8UuqnW5dQ98b6PDwbU
a03Wn01Un6K22yio/cX4uJyrYzFQ9yvxsGyjRsCG+lXFc68dEyBd51+0/1Ks
x9k3NSc3bH8Rg3iTkJ7JZSM8K8SLAGXpPSvmPYJOhAhEwMvlVZrB/Rmykwm6
JXc3IB8m2QoZ5BYMEhbl9PNoLoulhBgRCpnnCg1e9YPPwqpKorLxb/OAnfIk
sNfbUzaYenUvgkgYGjXZ5d2JpdUD5DbYCPEdXy+O20XSwjIeQiNsvpIv41pZ
jrIdOUcbDR59dGgowAlo5Gpgee4shZlJa0d7BNUI2OCAG+N/0rY9d4CAVRro
k3n9U8M1SbolS9nrLL8iS9y1JXftH1sFC0XAqE9LKiRfLdsV9Rbn4pIKHaiZ
t3VBHStvjlmIpvHA2e+6nsP/rCB+d22k80bf23Kn2aI94EcYuq7X3d7BK5VS
719CJT1lu//ZqEksyl/37eS92/P+QmIO2rXSv1go1Kkz55n9zDHiIzSNfYrv
UJqE00RKNO6IjRCEd9NUvaPvjlFJX73EbZcYqwdmeIu0nX5Pd9DfhSsfSwYH
s/lVg2R2HZ1CyS19cOikCmzAmGZBHwa9amkm3Tj6BA5exrVDkGH214uQF2zp
Efho+k2ZQuNRImw7X0vxaIl2C3DVEXraBEQ1drLM/+t/8rM7/xVCw4MHvyyA
Dp5XHFNOkV0IAcUf9mtMUqpcYdBE3DcUVQ2tvC+5ELUOOGrTT0kvmie83cBx
rg0Udknd2M88N6VHGl0yH5QIW6Hnv5BWXmO3SgVRdz8MTvlEvCz2o+GI6PIW
F4QACow7KBaI/ScZ7Mn+nJ4YOzEz9OcmK+4zkVaNDdWmHIwkuzHaYId+boXh
Z2p8IHQfKdup3w+s8qfDLCC4l+7uoFHSiet2QWbyw4V8LQ16mfPORXbeXtXk
4+P8PvEwlJylyyCNZtgkQXUB2rjWnb7CfPSjve3brSEwJ4Ok/yxH+YXWMPkq
OAV7eGgZeLntOIlXhuJbaImbdNcnGoPSKPS69W93V12fT7dk5HVyTrkQcSDl
yPOu15PyZwQLm/R40p7KNE+SHe8Juc+GrU9KTJVD3Mq9ur89dTdmKGcILbpd
26TrFLy1lSir1eQQOsbIllNMZEQbFcXvP0/yATCF/LmQE25A9vDjpCdSyC9Y
9aDKS+N/vktYbezmh6Fk84O4yOp59o6JxzLl2WqkmbC7y6SICz6q7VKM0Rl0
E+RazFpSVFCMo0PQSmUv219wpK4W+TOjOlYlR1b4UzG/nle2TOm2ZigzwK5/
ntirpwhTBSbdW6BVeTGcijhEsYvw8+Ts+x4IJw6VvWclLLnGxJ3VOnqwfeqi
zK1D7kwkp9aE1Fsiy0jEVKSzwZnfsiNXzapGFXq1oZR5bGZTYTuR1OSm3wXS
7fkeCRgWRJ/78YWVabAMytpmA9+ucfKOk07P1kFwIVx5S59u7tBUNAiogDA/
WML2CmD1Gg1emxC3ygo7rHx+AiGLf7yM/wY8BJe18aWb/HzfpgYkm6hYzYPz
gcNF6c1pFEdBJ2ytMllZl+fqS3jyhtkAz0rroaCok4PGJNUC+DxXuwQyeCwa
nsgts+IDPRKPzbmkMEp788jl/5sUxg13mV/86t7+jRetJtg8QZ1AdITrjp56
DpPDCSSfI4eScvODLCjqdV6385eZdJlaYq30/LvvW0rw+ULbgm2/EF4yN+32
XqK5Xb1VR5Qoi7ErfSzigjshixkm92x398Ib2S0p8Mf16p0vzXKxwVh1Co4s
lDKRSPw6YMueFh/8hutnelZtB2b8uHZ/I0MLDDuWQuhu+C7zIHJeNVoefcjG
gwNJIbwhjpe0ClF8cskT7wpDnSybkRKpgX7ahp0BzisxcFcKyg5tWOdf4Uf8
bJT24xIM8X42YesYIgv7U7V6e4KzM2Oo9fBjvj1WN/2PuiAXaj0g3mVtycQc
Q1b8LRUXxUhQ6kt6Rdat+gzVeOyYubnm9AvcwJEaBcfgoURYH7psRQMpYCzE
CpX0PyrfRCX3y8NYW9hS7XRN5xnaoFPgu0vQYT1yTA1974n0oUxMbRhy5teH
OxriNlyzqAjpHgHrhwsa/qjBKO2OdJF9TFfg27IAgro0NY3XQzzBaoQPpsww
fjLigD+uJU0w08t9lHt8OIMka4QcjCxeQUkCPYWWevpyoOcaAdIpIpKfqWcw
8t4p8F4VSiT9Cfq476aVCTkRvblcNSX1NNmWDfhKacO5+36e7bYyFrqjhLI2
0zBk4XI+JWPwBnfemZRw60yzgIyRcEwKCDhrDrDlT2BcAnbEv/e96cugrZKU
30O053x2u83AoHNYbMCHOgbPpElNL0N5omC/9yEMSYhghA2GdsOS1GQkYvmM
XT7JSzZgxPbnhSdmCfG++yl4gtzUSsHhtBOORx8oQHGSaL2aZ0G+XMdPzrY8
LbWLTOQdUKNUJyZWOLotKJDgpKPMLzZ7s/RfqblOH4DJWfu7HarKBAJVzk6Z
1OnbPDm+R2GmMbOJwyuD8n200k8pe+C1pcn3HRlCFits2ueeCcYgVJLsfMdY
LMXb4vlW81619ornOoH1D2PGney115OG4LqWCqqzQNqzCgxnLsF+YSaDestw
KsLdLeuIzczXOd+Z0jxI+r9pnViDzeQQhSlWBr18nlQQcOBL7EegsYhN/0ne
lJaMYh9dHWIuwoPAWRnHD7jNOgr3xFP5WM3CNvh4ycHi2ptqR/RntW33nW4f
cyqQ+dAvYkMw4m+72SoDfStwzFiho62h0aryvgcU8MVy8IawGDrEFX6wee9j
eLoQwQhdvFpDvIz7mgUWkw1R9gaAH1zy0SN5TBRclZFwTBF06HtE3kXgcNoD
AT5BOoCH0uGn8DGUagZnSG6Da4vpAb8rfxvF+RgEgxCvwupNlX5QxApG4Kdb
P44l/JDELAvg1HkNc2d/4acAK4SwPwokEssydTQYw/MfmcUyVqhuSrlatvfQ
6Ycd72WL10i0DcHKH06z1Mm5cLMtj8vKowYQPF05iDvqPPtrmqZmie8M0kzq
DRWeZXnmtDGqIoGU8lbxn9iT/ITSpjvM4tVX3DdMDjE/NlK2AMLaCKNQWdJ+
UmN2AYW3s9LodmE+cRjKfwKGVvWRm514j+K01WbdqT/jogtVFILm/B77z6BD
amHcwTkKiwYAJvNOjHHBAwi4pNTi80n95TpSBj+yOj6u31PcXy8M3zjtwkb0
iGPrYTKWG/zwdqHSukii1O9mnrglISqW5Pai7Qpb1UwdKDjOqbwKFxiniTcW
0H2oRN8PpROzkFa7Yd2d4CxXl621XYgr9R1FbznuXb5Naqiv2u2KdpTgixYo
GsjY1gmea3WNBMd9cGYplGNiOSG5KQLsRRADIZbXCk/OC8sTFZbRPSsHQKCy
9Shx/9P+NqVGzQtiNNPaa1KjKamlFij8mElfBdKqk3+4/7nb7T+fsJTMoxf6
8tf2FgseCBJYXS6ZfGudLg07xABfZnIYrWvo2knOO8xdxUdKUdjcBV8R9mJZ
+J222d/TaGpAmEAmMO9ixeH18Vxrd15U3LBlt0dDcvmU395CY5cPFm/Be9eX
aZpmMpqjlPioCe9MrkvuSKVw1r62pbaMzyVxHNFVEl34lInXjv0qu61/hfvU
1zpa+Sl/3ew+CrVpOgj+Wcd+XyK4+bEO3WiE6Ma6l0+njxMt8uNIVH3Smd/Z
dtDXdP9V4sRLAw4WJAEJbSNAHBdDsrxX3nmdgOQwjkGPmroKGddcStfLImyz
PI3KGdYka/w1J7rGYWDoi2rtwjMfHPJ5dJd0RtYC/CHCESje62EurSq0xYDj
tDrSjdLiiRmqSnr0Cp+STCbpZNbkEQTR4YdI8dIOBChO2kTdrAD8SQ4lPeDE
EwOnXYQ6lVRxbyBGjrYudd7W6RmkJG1wQFLYnLTP5KWofex5F3YFuAHF0LFH
XZCE2/GTtfIX1ym5gLWEBPS3GMe7kHV23Wx4l+v2SDf/V8KGqt/sYCtHa4mi
s7SJvaF52egxmvB83Rsx1aKx2AnmhRqUMKF0nPKRUGVIrst/b1YYggP0xijY
cvHR2G4ikBpY5+QbMcuKI/iwDE2yppn3OLLnmw7pbXkzhYClP2btyLUBOeVI
b3pJxX+UHuWtmRU3fUlzQuNX23CNP6FYV8q2yyL2ko4AZz1M6cg+FjD9A8+3
YcfJ/LYUqk+Lflb2jtEe0+cqHC54N/Z4FgZVaPohMGRk8S+i6Vl8Rxh4lChK
UXuXCrStV7NWRZTJ1PO/enxRxD3V+mGj942uKM20oiirBliqTfEH9INohWX5
vpgQwJewETRCUo2bheTHPCk1giS380qn6v/3KZCsdUFtM4by+a10cCcaM5/5
OZ4Wj3+M8/10wU/+O00G6fkuqLQ87Yek5S6KoCt2RhK4oRSIp0mUyrQdENal
LSQcKLdy06HtkGdx+JGDl3oqiCEnsRtIuX/+K05qDAquMK6i8YJ6lv92ezBq
+9yWf+taUTUPdwPm6Y2U5JXl7hrXpqoKwCkb3u5EEY7bm0l1x7XzsHaj8V8j
mlnwJcLVOW+kqKyMO/nYKl6ciFMxxiDS/mZf/A+Wbo6TdvQ1AEtaKsn8y8Wi
+86UgTtvq94TPGAVyeRLLgTvwk0wiRKrW10hDHoWth4oRQm+va1pBJd84xdW
E25k6a96n0jHmwncSFe56uJ2NLsJrGqpDUdDUHHX06YN+VOSc5vZ1E1u+6HG
LBD2oLuHVgwXkEjlnnh5nbO0JltUefsG8A2PPWKxyIi9B+fRXqhf22kXnY/t
XaHGsWjV/icUn0Baa9mjTnEbg5bUK+8BgxjOepiIIOlACsy9isiuopMFOz13
H6aWWN/AH95JwySNu8mVexcDFvllMJz3eUofExQ35LTbWK75baL23VH/ZIru
NJZXr6GjqNNTRH4V1XLrH99rF5QXTSgnM+1axEhU05OWn01l/M0KFmwT6k6R
gbw4V8LQ81RFBkJySaHTPNTksKciCi/Kd5Nn+Ixbk2SMfHhPeBphRcJnR/5i
XSGlSxVKOIk29Y91GG/43RAJbeF4pWyDJ1SKHJe0xP7+uCYrt9nYA7+vcjZg
HDS1+ysZ1yJ4pvklTwATT4FeTj21kT6x8lAOX+7PW3n41IDuiuOlKGIGfaSV
oU4GCaqL/uoaAU4QkBpAca1fVoECxy3O2bpOPZaLerUBrnkhs4DIHtWIhoIH
rwzbOzLYaSGpmerXLO8LalCmoNvJcwjX592+h6XrtgHSvA0tNR1lHTjaczAt
q6AE4dJRvwSHPi2qCIWwmtIlQusTVlhdNcPUAUyZqnYsSZRfcbJx1+N3W6To
TTa+WvgvX7ULgDg1aecBdtFFYZ42jYhjVXmsE2ex5I8uS0sjUVsxIwrwap7s
vdc/LjOKlHOcMXlTaOePYQ115lvB5LtmIJ88kRIpejo4631Y4ePue2a6kiPU
pZrsidrhrepjDTawynIOGXh4dJoWz1SLE10/moiRzRyMAKbos+3vefZefxTT
x58YGf94wyUEQhLxvJN6eA+AqrQaxX2d3A6BDwxGIgCNTdVsboDOBu7Ckqwa
B7HnqP7LWkazFWWUL6X/RioXAN8cms8YtieZAL5RUhx7k1gxJRg64+e0dOME
pALMmRLoI6aP1QvMf7pnOfKkZJI7D1RJNg3PwCcGqPmoCN219ohd7eFLXO8f
jzjzpQlCj4Y8dKgmpPIsrih66k7WP9wFcRJ+wPHQL7P6npfhxPqxa7ejKJjp
DidYj5+jKigNs2ef39r4dhIjMMO9n6NbMsXaS17YEK/WpnxGWQGH0t/yedIm
qlzAQe0x6D+09t6AR0fvq0D9JlVSKn7MuTg+k3V2rDsuqCHngGpiTVWYGoxX
la01UCtVl81vDa+tstK1aAwcbLhvUvYgu1gR4LPUacQ5gnbYFIFX9RQVDDHK
MaNp0hdRVp2WhT20cSWdbKbfXZY94bZytWQgm4YOWAYt4YZGQMkzEd2hEwaj
TyTKGfsjepFOeevSSh/fsd2wwJH63hRQS03voUPyj7X9udkv4DUB9vkU3aMN
+DUGsLHemH8GZmiZusBszCFcw3cqHFNCUW1A9KRqVtG5y87A2r7mpZ/NoynG
Ti+LRp5JVT3NTVXmcQBRX8APHokY8LKzXqF/0s8aBA1/b04nJ/Ncfp17McJl
Pzb7Nph6lUvRRaAntJOEAD9YiY9Jjg5ZAnf7/21Ik5NW/CZvYDd8pre7M1YU
VeVu2SyRkJb/IiSzPts5NzqbKv8CqQsSEp+zDdeGzGISWR4DLmhg2auAI7ea
hadWcMCtSfLPK9wgr3eaXWJUuvoT7eefTpnbn0KCubmelJUbTt+eTw8W4kP7
sP8aBkzS4Glj258NhSTaaC/TZAKf+U0o7cABgawpBsqQtDX49v79HClnSV0t
AERTipnVr4p4+N62FA7URyYCPEYaud5so6lG3dNCIN5h19xvaLzemqzs4AOp
NDW6kjICG+BM7yaa3UgtaHUSZ82gteefWRZv5H1EdumEQpOeFY+0CcyKteRm
yfUBL28L6gc+QTUHSKf9bfukH1D439aBU3+/f0B4BGPvE1umUJLUa3zZYR3F
MRb2wDmzDYHB2nBhSOXmTg9+JSS/fshtYKOC35jC3MOsHSd2/ZBGnoHHm8og
2G0Ub/cpGmvlalv7SFhFcVZSME6qG9JPNqI2n27s4425G36W7cFMItNR6Vw6
P0q1mBjiMvRCGvmv2eA4zJtFPD68R3dnIHKzVGPkhkzp6i48jmSiypvIJDTh
gwjCRY86eYt1znU1mzV17oJ+lt0PBFOCYmOWJiAlyUFzgIlZfYSQ9kYAJCGF
BY0dlFpm7UBd5xmAqOQ3XfpmyZwPjK4mb6pZMvja2WdHgdiwxfQGjD/E6Uke
ahWpzfmG2EP+BrFSlI+OaIR5Xz0jRParvc/fOmGKIT2NDLSZEOqNCnM2GSLy
E+t/07pc2OBx2CmtTWaIub3H0qAU8n7/ojy/HJXC8Zet5aeeGV3Op512ndxv
XRe+oVCkxiAOyDqKDFJCa/Jbdgx2qVyMZCjS0uQhzH8daGgjzGJjbrgh2NAb
S0geTA2ccPr2rKV8hqhYFn4EjQNimHD8+xRleY3kX1Ai+JtYzQKjTnzmF5An
uHo+C8c3lnVQ5IRymW7TD/KxffQHIRtGtJbiKJ3silU2S2y3qKmW+vfVreYL
BU+wRnEAPVQprC3TDsu3ij59099OxJVSPavnfyrPEAv+gaIJyIzpLdJ7gUOu
jdwOjnJCEsoudHl1qkUm/fxq5NuBuS5t135Giooh4yqj8pVLktCI6zQeU8ds
h2OYVADaQrM9JlCe1oRm9KD/lj+kpg7EfEFwEJnBp4DtPvT3mZfIhjEVfOsl
NMhX+oxriXHK48Q/+C7jXVN2fsQMmbDpRvkEIsZ24OkmiRHehpWS0U814LJ6
sYqirIoimBiNJGi4EXD99efB5GoTYhP42gtthQnREyKxSNVWS9UhQxH+PY5A
rT2XuwB5lLeaIctsNCdLlcS62TLzN5++hUBv83iJ9yMe6MILWYNRjsw9ytGO
x2NBnjmJwk2mz6cTdbSImpE0KDm/A/O42u16ocdFxDTLbLA1eYOx4ESi7Ybj
OD2zJHSp6CebmBY94URycAzVGc++kO//3v5fZlAmKQNvMM9j5BF2SVq56Vy4
Mey55ohZd2MslOXutHT+TgzIM2GE6PJjZvlUOFXPZe2/xEkL9G9pn7C27uX5
LaBzb8Z5mOZvLCUHpRoriUJqIqA+efjPdLHKX77V3bMNERxevtvVaOQuG8Ut
bRYNPrf3TuVjG2jdCorj0yjOrJaZ3UAlb1enL/MD2lg71bJi3iM3Ue5JeDLt
qNQyYeHcfS4qLgMXCeHhUoKK0VuKeoenSzgLaRhK1dy9N7IGiDOgY3B85tm7
eqkQms+GrVcnPMnie2u5QVdU9F4M+TtV9XndMQN5flyqx2ti32DSLnEINGdq
EGl0JQaqe6ldNfOBmelGvb3kEyo2VDqVOm3vxl/0Mn12/0Y/LLBWBPLf/TM4
jo6Dny1gOVDtoOMQlCewGjsU4r2aEeqZeZFQiyLFvTqegVKWHcIlnH4na3zq
S23PImI8oPn020ZwWWGcfpAIIEpx19R1bNKbk+viBVvR7Rdc3/mZxnKIduJX
ZRcFRLNw9bk3uWoTlHyBhnQfEoFcd5mZ/PaCdfBTTQg5qf0tlQV/1eMbPygE
8CLXQGmSbTAYN84GJRPNF4uj1w8Pirz+vKtSY6/zu5REGOU12dzPtHyKzd8P
IWdrheW9fbaMZkAbGmnkvJWJqnHMgR/ZIeS/WflslMely8lAk8uWvSXN5qRQ
hVDFk39UoFD0VHJ7jMfTvhetDhyAlpA8JedIr41wPf9UisBkoP45GVqSsVLX
Iat7M0hfPQCVZ0avKGrfMgA6kG2qy8xThKKtAnM2lifzEn8X7r5F/upcUVVB
3ez9dvuyfl0IE0lIaD6H3CWTgpoqWnnRzC8FPCpYsPd5p+s6hiS6twV/Nb6E
MpCAV/WaCfOEgsXrZiGSfAzAoTR6f4qkWu2SOvcXVHBa/cH027EMB/9keh5B
8RkLoAfoUqciko9kkr4GEdlV5IMSijpaqTH6O8Hk2Vtp/uJY7c1nlLGmeT2D
MTGo0CXUvZBKEGqt0OFZkV35q6uBbCCs5nSL+sqr7KTZjZK3Kne1QdcZ+PdK
nHPicrmRcYj7tTvgebuvUDbesuFQOSaq/qhy88nrYcl2gE8sM2VrlePVDO92
ZzqsJhjqwOXd/1zATdbipyk0OZzFeKwtZ9zGO5Zkzxp24qI5QY+HOB4IbrU4
mt5kkKH2AK+DSL+/jnV0zkRY1b6FyBpzIZlTL+EVS8lrc2XlcN40ffQtmhju
XCd0fkcLI8gAzO/ykenp7L8+BjFy1tX6RIOp8PDz80XPI48Xn5rvTckgCx+6
Ksh7BAiMfW0vxCNlyFqM9G4rw2PRudugABDIHXpQkhnWJp24UE4Xpz1vUqhg
zcvmwFiU7hmwIMaypWdCiMeNEuFhWbotqHf+uY58kvzI44t+jDcfMNkLi+Pj
pVg0KrcqwCqGhty6/s124U+IHMM5ufFlBpFPckHi0SWa+v/CFHJEOrHEQY/D
I9Z/LPqtDeHF5ypyNmvlCZmAs1CUrUde1jpU27Ug4vCaQH84dNOFl23hZ4FP
Eu+nmpZYnl9SAO/D9wLNIn6EC+qhzWRemIzHXMXXa7b2l41fmxGhQq2dQExo
gcAg9RCmzYj0umHlFUz27aiXUKl0VYkVxFP3W7wN1PUbIfmFZLyOPd26GTiK
lz9cYbrNSZxDLWSE8R3FOqaEQYaEwj3k+TI5YpS9Uj8w/eSL710TpecIPglZ
6OkIgZLkCWtJk0tPrm8bv6Szi6ObhGOx2Oec760ka0C4eJ0FZdr19ofluqgE
y1/ZXYQNjbxDGdekOPbY+qIYxEcAsoT+4KRsEm6DZ9nObw4HlWej2jTvrzeb
3kIjgBNIZoKEDZO4KGGV5d/iziyKPuqhauo4jjvHtg5XLUdHgVRq/QzXCEvR
akKeEAWfEikh6Fp/T3IuhK9A9clxqdVLGcxHtFtP/Yrr9hJJjM7j9uWa3/4X
8kux0ooTYgQj9RHeBmGsRPDYt7+4EbbIuBPIxDsO3+uqRV/cWiTI6shc85tN
l7n9Kqmbegwl97wJf1YWUweHMEIIqAitnhdhq99CA3Cu537ft1r/dgalUlWd
G89aauWvEa2xCJqOaD/9dvfQ0XdviJr7swxh1bDvkE+Py3wc3qG1n64jKbkU
J/qJKkAOCLcBNJxZLJ6Vp3QQQAUF1gSem9cfQArnpqWMk1KzeOFHjlOzYudB
Ggi3HYf7WrJo6Ffhst2ZUyLD0xtT7AHFj6Rli9aKQzAQ2YjxKtSRWbOengaC
zoz+DefXwU1It10++oogH3yMm/dpaBU71AyrMhiNY3R2CqnF8PiqaJx/CYmF
rAId6cHyzSBnCOv7dMdMHVOEBG/VJEo9wxgflNuTCzElMAmS3rLnC6XJroCw
5GE25tfNBIYWFE0YjFoVpgRo+db45HY36CKXTfhFoU6PK7GpnEN01yDKu9oJ
wq4Ed84AFYM6iH+S0gUdSv4NDKPLlcoiwH0OJTBzANdFqbP1a1a+0TI/urwC
Bh4PVO7U17Hh1F7Ksf/OWaC42KQxNEGFFhIoxni/tla1gvPslHZRu7x+8ya2
DMOMGeM4++juiEgQ+kkmPJMsKbpSZBph/bSIPcusv2TC+1382DobliJc4/n6
aaIayuBtDaqVQNEbhwYU7dghrHGWMjkUFKBaYE4k+8WgQaGsm5zpimbPSa1w
cPw0wD+xw8ApaxWVWz5lW//QPEPbQBOBIqinzcfgIsW17IZ4sTrKxpQNOJ5U
539Rj//gIkJCWdZqbDSc0ZUY/mnSHmP0Aa0CrWuct5juuDWC7OSsj+7hMYL4
sb3PXuSUTExPMi6ojOMzASgLcAVCNhbGRKlq4dEAdwNLEVW+4x0wvOHQY9so
/8ulaFjuE0WN20Iqmsf2g/s/tnR+btoP0QpAt9XNOd2LiXTT0JWCkWymPToy
jeQ3+DhQwX8Fha6fC1ON1d0UMSqh2hxHJ1S1NOW9ZYaFjmroQ102QH2hoowY
gnej33meAc1vEnXi+jz3v7PJM1zuuCB6or1cLiF6BIII/fimtHs38ZwybRrx
0K8YUe5ARAbz38GZYLGIQLTZ76ehdjpsulc+5V0p5uRFlMLfY4G8dz0cXykV
R1TW4mt4UybbbaQC2GELG5grd2WSjU+bqoTOp6QzAR62iTrM7g6Lokz400/4
U0Z1hlnz2IHYf84nZsAZua/5osONrS6gmDchZ8ce8cVYqdl+CzIa/kmQOom/
ZALB9e9zF6f/i22G9zj1GUtNtS5JIEtaBg2bCDqXmufXC4+6KOh1/vfvC7hv
LLsUL51Pa61W3bxYuEHuT0Ht5afZ+UtonjHKK/F2bSSOSL5SYXFamJFdduZC
PeDalBwSMMBis/XpRo90x77vu0XKA7BYNZtDPiwXPtXHO6Gs5dOL2IrUfuEd
9VSi34EvdZRHT75psw8MfvJstfdQP80HTrbvK3gL4kpB5A14zo9BP6liDE7O
faHgfzVLSz4NWZiaVeCjs/zT13dNhmKV7E5uLJRzMfAnWbtwsiII0ZS650D0
+YQT+K/DrP/zz07E/xQMeD0XkrogVi65D1CaFFHcakwZxYluDDWx99v7KYpY
5t+EuXRcFuzitO3kIerGCtWnwQB3wGAN1Yahe6lE+9nK++SCSI5xTGoR/DgH
OeWzEvVasmmifxhfJ1SoqG9zHWhCzjXf/UVJkpHVyUELvVeE7dibBQoWMgVS
152XqGs3fw+4slFJcJvAt+G4giFywh7wNgNEK6oF3cKTBN+0i24pu0ctjJH1
lo7VhYczrJgd9MYQLnX1B350jP7l5uPmgMO3jwwq8XDFoC0+KbfPoxWZKkUR
hW7w9oEoDq7KTqzza9YGqDcmdC57GlJjU/BuEcNaT9qPv8FsVfIvqrzjlpxJ
KXyNuEUeocak8flQhLkmFvSpiUIW/fJC835SvFTVv2PKUGG5qjvtTihrGvj3
kIf9LNjvHsNXi2b3vmwtLhbYaeh+Wshxbci/P8f/XFeJcw73IVBjp75sWBMN
it0x8RZCLsrFF97J5nhCjYGcpMijFWiFEX1utj+Wn/oYumCM/W0xZXcXjppp
A4+QF9QENo9WiKzMkBcmyrcTbcmYbLFhJfCc37dexuI5pYAWpYkedVQgHV1C
Grza6Di76e+8toFJrB2T4WmSjYSrrCXpHrF7FoOQ/HHzVH3fQKkM5+3rOPk0
XMQuPW2XTkYgNomR0QDjFeUzSlaeIFmtzrNGEPF3W6HEsrUn6r3sQCthhnV2
HtxtpUd9HN/wOgkuc70aSn2fTYqk+BxAxnnClVMpjsLJPEQ5rV5uB85JZX6x
dzsqfIJnwVEXkTQxEMDHHn9pGKZewvt/D4xYAJO+cHdEP8KHUsFiYamkXVRm
oAsgkZQ8oXC5SubAOb6Ea80hO3U19eMQHNYOgPhKnw7Ei0arBG+i/dAXVULT
MeFxeILlfKQwAl6E8pPTszdtLVV/hqSIREvfBdA50MQKfq3+A7iG/a3YQnt+
4Krj9yMM5nJSb1NFUowF2OndiuFA+A9ZzLDOe3y9AoUGc65sgp2sB3b3EeNW
TREBQwYZp8XMVKyyztX53fCsUstQIXnbmGJACHVxJztC51XqjmernlyKTVpB
4t+yqyn27DMNYCL7vjUJCKa55hRYO/I6Cu1fZejtU34CPd4T2f9ZHLMKS6Tc
/ub53MRBHnItnmrkLOjmWQ00HD4hK3cqkCJkNif1QANJ6iCYNzsG4E+FR3lA
k20JUXPdkFdkTwx6N4yzwFIVaXEgOEBfI2nXWo6Px1Vl4+ISPyJBbVRf8DkM
mhZnZ0NydRYMUtwhnihr7osKOFwiKJWUEDWHz+oIBUtG3wroccZyK7YSQ/Yg
RLuHh6R89hUBw/TdwrlxYffUqBCZQQFgL1OxmEtVXpb3qwP+L7erVa6qm2i0
UmC4Jn8Ct45wo/ThCxdsXT9WRPNwQxJUZhjHzLfIUTCKccYvuSI14CcVSAU4
iItQsKfm87ISAbkXU88PMZmN2LkwjUQCRSnIvNBP5vDE+UqzgRlu9GgC7P4s
xDoTJDnr8NUf2chZmu+BxtJQGqs0d7P5rRfHkw1yhb9FsnIgwaLy9kLpTL74
1aYugFkdqlBug64iLlz3yrda0zqHn7qJgOEC3mRzAc4lYplhGnz+3LnASEqG
OfqVZJuklE1K0BVsNkKkurYfpPd76ioLPU1dJ6wiibEJPwv8QFk9W5C4stct
V7Rem46CNMdwMQQW6CKT1jvfZPuhRKuZg6Km7Rqy9j85/KooMHn+QIBz5ec3
hXKTL4oECU6IONknizZDRRoDVjVA1TBrnOilGJ+qBVeMXZDmyIatUEOL+qvG
dXoknt7VNFTJHC3PvGuZ3I0m5TQWceXQAm3KQA1rDIJhpZcY3+Ho1GlQL29G
KxXdGLgtEVFB850byJVUMDvpc9eyPYEi6ayu2Np6TDcmbe7C6OjsGQTKw1+e
tynZQW2sz6SRz2TKGIgkfTFTfy9yRU67GHGFoQiyHCfSktfNxM3hPKPdjtiG
/waedwsh9l2DbKLlKbmUP78s+bQDm1WnFnfHBVDdKb0vUX1K5/eWUCNRyZid
QyFj0hWhsKMmOzKfWEkPPrJTBk6d7U2uDVn26WLNLjG1t89kkiaeplUh7qmy
b5jXrCcw9JpCn+bX/Ykk60+O8dtDzl/w2UgKl+9fBIFu2ifm6PtOTe9RFLhN
4EaGTcxt8n1IlfRAhc9GjgzTsJr0P4dNcv1I/NOhsvK9Ggmg7kbDSqQihPyK
L2B1IVt1YzEVnNaXiGMHgkINEGPRHIPErgKHBYZ2BUsXMZKWsQ9n1ugYdd+S
NEsDPz+IF9bfjM3NLL3Vlb+vxcOrSdfPk5eu0lRg2M6BbR7pFE9q8A65McGN
5PZcFED3pyODR7HMWtHG64f0oxejE2dDDSHABKFlIt+wTdfYM0rawJXDrlQA
MvrDJqIPHJbljkp+/4H8JJwte/2C5BHEQ8+QZ1/HHBPmah9MjK3A2Oi8QCfn
nXX8lfgcG+93eboxAD0QiuFboiZscFBdb0YPku/sNX3uuJICGOwURHC/1Pwf
+ecTx3ONi3nepuJTDbylDqd9rpqdQBqJ3Hm9R03B11chNQ5XtfJvrNc7H42p
pFlFSKPdOWvcGms3v+iry6tw/gjT6/VjnexmAsdvLiF9O0+zyyI0S8X/U6my
MiMnh9NgL9eVoP5t/RVJ/vIookL1E+BJUk+5fR05H7p0QftpFQAI/pg1MV+y
AmZAjCgHrKVLGAyndI08JwFCIo57Jg0fg93sEz1ntr92JSRANwhS5TnGcE4z
rSjsif6vuUuyScQo3ccIaRLKKkjIgD26haoWZS68X8M+HJzpG7762ay3JdO8
cSimJruUT0VVX6SQFFx1ESUTgQiet4YdbawWG1om2OnX+ubHaclCESvw1qk5
kaLdm6aGI1t3tOdYcDHM+rx5sdfVPcreqeuDQwcg3Qnw/qjtdfprzqwY9sab
vYxn1zvRYhxttt1FUDui+U0S73fKPiAljHQ/v4+hfjCgs1ENjChiSt0W/ag3
8fmMW+q1jbYIeanYeSbKj0jiFGEbGc3wgPR0u73xK+6MMLaRDoipkic5Vpng
hFiZuPG5aD7hz97UvA1H/dYl2Tywx6SkWuBtu+AxOxFavjog+HsKgYkmRjvf
aRTbnfSTRAa4cTk5QzmV3SHflFKxkNkjPL2rMguP0eJSGYowx6uuwRBSfLMo
gRRIvghhusXY50BUJfG3SY2/Q/uT/YynfTT+vyFRzUy+4ho924D/Ul5J9Fc9
IXwnIg9FHkMWt7UZ/b5fFP9wFPSwyHtlbIW9TpnXwbxw/35UMBKmsXkrjj5A
6NGC3ZmoN3GAt1sWdzEqKhrMOC4eL/7Zmns6kC6wlQTP4Q/aSV3tt3twxjdU
47qAdv3Aa8qvjzNW3sLndL97f7Ovh22TCaoyf9M3aMmS/NzRdT0BgLxeJVvP
THC4dAdFcn+WHXaorYaXdniyfoDPO9jFWXe8FGwnln9Zi+QCNGpkGWNfRJLy
FHvBhyCqlPnr/CpD6aHE6lqcxv8g5lI+ZDb0JMixap4iu/mzKjX2CgoDKx7x
kSXG+M8Q9JwO9d8ePQDISsM1mvOZTv+6Ca7L8H6M4Mz1ckYFJEVxU/tpG5GQ
Po1p3spHIIyqweDd6dfMIMLPMQdBqSZoLyfXcN88+wOIddm5+1u3c2F6VtlX
rlyrAJ/kkrpoWLnnH9A0dDkRtDi6l9JvhbYE85JWFK7A2r6yLr4+8d/XGpD5
+zxfiKntK7Zs6jI5GEY3moN/akaZvtTQuUWUPzVEtuF1fJ6MpTHxsfJPLyFc
HGi686qr5heXwcRzXP89Nc+XET70JiQsEiruhJfA/YuZ2keNp+jxVboBH4m2
HoTx2csGOi3TBT8RF+CaqOY1tIDS4n/7vLeIBdbTB634+2YEoRzNg48B2Nxn
eADyEwUsO8hRCC/pyHTPUW4KSHttVfjhboWyC/WhKxcb1p8bEEn+DuA41I7H
3rj6apxs7iKs41qRssZMBO2z8+K/KJwO2s1yv8kDid02SXepW4UhTqy9+GTa
UT6ZFf1hk+XCGQ2X3qQJE2X2CXcFv018mFE4NullNwQnmsnkHhg/NMcS/Jjo
sfvq8PB2R4wywrzKNnHIDktwJo+Rykwg07EY8PIf3pY8Z2Qp9FvQAfxUyzp3
OaeyG7Ul72pgm9gVqennZ52147TxZaAjNOSLjv1CVXLhi0HLYazr8aCCulUW
Z5/dvZ189dmgt9h3cet1fyrq/lo8cj34esubZX/8wY2tbdOfJEIyLcOHNYTW
Y2bqUZot85poDf3Rl3JSx5GWywJmLuDI8j+P6x87jItLeR85SBAcmi7aV/gN
A5k0/ijtaE+pbEpctpVIvZCAOqW2Y9omOoeIi1pAGEm/Q4BEfSGSZOthfULb
exm8dvl62PqBESExbL0FaiCgw50owBMujvZLmhIAfJ9Wrp5rN8htfCjEzoSw
K5554H1C2hDD1G/a7Jk8/2DmgoE9K29AclJkjy+syi8BJN8Mjk0OPqVEFKp1
Rk2mCs4MBl6PXl6+uwWQ15xJn44a4zLfNzOXlcK+r+sl9Zunzout1xnYh1p4
zmN+azGPTSgKtjJGix20VfeeBMim1GDOc/0bCIbdtkOljoWkrQ6XQqZT1S9w
KZhDUvWb1AA93pVZOpdHz0z4EhZQHDF9EcSsDUM7nL+d4mPffKdPtwAaP0p9
y00D38pj7CVGZe69VLR7ulheJ7R4bBUlVGHVhO0l1IMga/sSPnjIruQfZg5+
5JQDafIi+EJwqC4sQmX4hqQMa2fldNWhJdLRyCEyKla/kbi3E5ctEU9jREL6
/sWtQ2cDZ21XgaGImSM3asSXUe/EncRVIjDvzKAkrPWyn6ECUL4x/fC5xHOq
5NGiLpnshn502Z8P8JT2qsEUqJJrposJUWX2zGfY4nPwnrbCEDRkPn1mIx37
amCbE2WkIdrAcobafEK1Pd7JU0bOPGZz1VFxmbMR/Aavs5BaconWZwwm4uDT
sJ3eFEq1bbPeuB6vVXuVs474zGVmzg4xxwP/qJ7J3s7MsLVEmf9GqZlHqTkn
w17KOY1HI0D81EImrwcLZt0hteTnoz0n4S0/TPOh9aZOPMvy3CBzuIINdmq3
V/0vX36SDe1tA2gUusSuyOBa8mfA0EFOI7xMsEXM+xeXUniLOl47FpoNt8xs
aoFwLpYRtM0LVCTGg3a+6zeI5d5eOftL9zAqIfg15BCe08eYkoBcI/0AAeyT
K+IkB73b+LXtGFl7ea5KNafZyOWl1J7aKp2oumEfN9JW5/kplaBuqDXviOCN
tc8wJBAuNW90s8Ef/Tk+hEp9wxGfg5r9fdbKdCyEj2Rq3nBfcQ2sC83voxt1
rhmlcqMH56wZJo/QOYupBKNjlTLLQ6T4OBj3y+FoesJfSYjHn9e45cqexzG1
u4Vt0o3mHPWafZmEivRYDdCF1LpWeF1+co4obwAjSnYOz2vovF/gcR6QoH9x
318Sk5Ri8HuiTrSIBS7h7xYgl9G2gnaDQmi2sl3x04gx45u5UdVbXBxbGNxq
+ht/UqUzbWe8pQM5JININAe/F6A2SQNMXvcoL4mkxIz6SleY1gVe5Wt3aW+0
w4+GNbJ8XG0S7Jwp2bbqjafQ3RHa2HTVpphfiOnrJ1BPsjKx7rI34CDDc9UF
+cdLlc2NH0jkGAgduqftx1IMSuIRaQrbEaOEi4i2N9CMfb1kIWikozIi8FA2
WBlYY6guG482Fxq33T9oHMJGxIuW50nRCec7chGYSulidqyiGcFy8Fa2HeQ3
knQ/2X+ABLMiUAjD3l8HqAZUnhJGsVz2SmmRCqjPf/52gKHx5nDcnjoSANva
tIuF1p+qIfKoFAm1tyebejfXRkqpMbKGwKlQ+dKWV8gXHEElaROCRHH1MXhb
6uc/BGSaXQlqOktOMPcB/zD2zeqJLvwDeEung3bpwudT9G3ijMNcWFK542fS
A2lgfCU8t8qtYE76Low/lPiJnk+xTJulvJmUjvzKAjPojCxlYvO9Z1ccl/i7
5GSTuR7jwI7Qa2xNU/6GB2gY1aJlCHj8S+9FiDnSVo0J44Cw4Bf0Vr7jSQIn
MkHBcndWTwgvm2UHlytaFFiy9lMFHhkqR3U5KFNVG0yLFssXawWCz5ZPVLNt
y1HTjPDXp8eOOlqieOUOWZ443c7zF77+GJvFb3xLlAKdfwYhs16emf5EM0hB
XCL9mu9jXFagm2CPTbVMU+KeLtplnYIUKskg0mz8I4UbveCyiAbqoisw+MMV
p7djNVXHnWNn+byqdUkAh7QoHd2GO97DtppBJ6NCuhBLbUIR5ZNg+HNPgZd9
/DnsTkp+0JSyKJEqjLe3wapRzOTNHQlVOs+dgxWKaF7NdHG5fOZsFkwOToKi
ZvwYuLpB7avNa/Jpuc4fTWL0VmJytY8/rEp6l6BZFuy8aSt8vMBbVp+1n3oU
8TchvOCDqpzd8wNcH/Kk4SAle/JKjOoiUvp/snhseSSDLuwJYIWFZxvwy+tQ
Il1vhSHgaB68g0jAkIc6+s6tSEDMLDGVDqf+V0ETncQcH3EKFhAbjXI35LYG
x2MMRbhyFEgDO1nfL4iFRAcyo5vka95FSXFKGrtUkfM4Eee/ojsEwGicMcj9
z230IvSVtQNljcOklmCMqh78bqA2/7/3/6N+DnX9xTU9voLGYJQOiDK5U7v6
nx1KcBWQVT7gPS8XshGWotI7LFv6X7f61aXF7PUth5Qr9q/JnM+dm9rKyM9s
JdkI6VQcsM6s+yYuLVL375RHad1UgaAvjZK2L/pzhK0AHalVgN/4AjYhCCOs
Vt03+aMdati+If4xZ9S7EgI2wlpQkmNSD76H21nT3QGnFNsq5OahtfMXMTsR
5xdUv7eGDacE4+j+maUbjnYwkCc+YfJ1d0LfVlJug42h1yj9/rqhD4j310Sn
5b5KZtnrFjXer0s0D8oIoRwlDuOUDFjVtSLjjZG1V9FIutjZX3EVkqlfdCR9
wXnSU+6/faZyi8R4RqdB2GR0KZu1upXecxIVZdbtFTm8CnRTALV4Qvnl619v
hgLSscLwU4221y9hNjbd5rFXGZf3Q3A+WemvnU8ufixQmv5QCpnYAhA74cD3
pua3k74Uxp0Tv2Q/gODSx4n3O8z6Pz9Dvc6CpFbDEHf3jD5n9rkVKSodPeSH
qKqjZU+QDDk+y+gp7JNrTn3ss25OQQxntgfX0KAdmmRfTt2ultH3Es/iQZmI
fHlX9mwBfP1KVMvcjNpN94630noRNa6m+Liq8Wqe87NfcWSAUdgm7kqtHT8L
rcwZOhXdEr3Fy7PiZRpGknK4YIi9m7HSfUfUzgZkYiH3ENv/nJj7EAiYD5zQ
B+2f5xMjCoWnKl4+g1FZ17LzqctPURfxEkQC7CTFdvEQhm89TMA/hs+nVGTx
OG9cdQ72hBgRR/D8jGp9Q2fpBMac/5Akdi8sRTkZL1xozoKLbDQgPQ2MVpvo
unlLIPD0Jcmqf1gkxNos2F/9F4HhLH0xDPdZYhKcilrm6rgfETdPUu0GrFSy
WDmtHu7UkA/kLP7Yy/7A9S5p65TM07/eq+bJNfQ7X3uodrVkUNoXAxPvKaGO
mgvRyJMZsuPywXd0jYcpwmXz6zxz+2KMzl/hKeZIZwbLWeW3ltvg/2I+Hl49
Eg/8SA48g802lqlPSkNT2k3DMu1N4o8qJMO2iGgKLSrOi6liumNv7xX/WKz3
RRtqr+Ph0wRL3TdbvvnVwo6i8xlF4OVzhJjiTcslNyQ2VEGnDfBJlrrrwRo1
ZVeqVnKznJVfjJYkyDyZPSzt4OzP4wcFRb3HPzWpVVgKRb3lrDHnOnZN/LzS
ctlwZwf6dzfjn12kXOV2UUWk+/0HLTW6zAZKVerbxXPGUcSdxuY5ZmEktgH8
fKqxQ/+HogfZJoPYUpnjJgPxwJQkIc3ixfBkasZB2kJB7GLOumkjLcRLIFa+
pXqcRXhdUQp+NOPSvwsNNwjr2d7bEDrY/oRPAWo+zBmzVlEXBRX/sN+ajcUS
M2jMHbfBASlNh07FU0YroGdwHiODOsxf1Bq1/5nRp894ouwqkAcSealwrkJ+
98FVVlmxOEFkLNPZReezCCsAH8xSor7/iWqc7CXu1BQ7pFnedD4TG2Ks3Y7y
CCDt6sViMRSUfMRTBmo7kgrRfusxDekNt9Lrz9xd9IPt+8sf0+qwYiT/U8XO
Q1dXgXunS1h2lJ+qsBY6CvGXrxXO2xsbm2R/ojOOyanEF5jiG6P0jLNjGCH2
BtuUhxQyHZxYpWMKSzcom7RSM4E0ZUErftyWn1J5sTzI6dRvOQoPHRCruIwP
lpaNIVIPsMUBRGuVVA3NCK+3Ae30YT3DIoipYhbKRkTeL2RRU1MOAchZ/Uhz
UjdBK8c2tCdvp3BL7cQrMuzDlPBporV7NZGWwm/C7x28d1cw4KO/UQaWkfQo
U4uH/JRhaVivsHBHS6Faxvj2AF2/HJZpx1Py2p/bL4KeMdUjEQhNHbJcUqqc
KLu/e52Z+voyx5KWNISFXgJUW8ORv7iy9mP4un2OpcMzTr00efg/rSKX01ln
HYuOGhmQ1CrxHj0FkXNFHqssU88qDo37fsbJLLo58g324gahieZypetDRJR0
zHlzS60zYCj8CRRa/yQCPjDA51OVtVmPYKVinMNwJJ40uyI/QBqf5GBAGmj1
jb1acjsXZF1kan2ZqKXDE9U6q8dpnAldzHgYTp2GmSJZqUhn3R2U/V7iS5em
/E9L/weNtTudwh7IJ0nqYnnJ83X3DeqSObUo8OJ6+pNmA4oMslQKpP8MpDbE
2h6v1kdwjfTzf0rCe+twDJpXW2HXs6pAsKYTFyDi8bXeJDPKZVMFbRYls7ra
mUV/BHGCBFGufgy14VPQXalOQND4yDU+O7ldYNYuujZVv9JJ0CZ/ghK8xFjb
pC2mRAY887UsA588k+yKRoKpHcRFmlspbHhKViIRhK9n89f2fm3uOBXtF4a1
V89+XcaImdXkrV9qvKGEQKfcavwSFOh7wDSbHK8LBlIQ8WE1VQW5RcZZYLR5
lVMKGizxjChuEuM5Rq495yJ3/aEH66zo4tm5k1S8NTTHWaI4ELmCqKRPIpWx
fJugkq3jWIoLyU67AlPV0bE1JlTgv0riZ9E8PsKPA2LsUOZeoktyO6oLl+/v
QBHMIA/wsH+GVIX+CHRNgdkLfLgjGxIaCx147lSFzaPXfW4CdvJaeAfX4PJi
XAs5n3kovLe3T6L9AJMMDTN+qA47vekwFrFBE4TT1lQbnHeyba0OlzoK7MnY
dXhRi6YVUd50Ecc7MJ0Wj8WUdslq5gSvd6mkcSDOJbBIh67nW+G/RbNDdtZ1
9FoOmYveNnqQgcHa+NIZDvIl89l5OONPna9USt+LVX6qX2ln9k5mKpr/Mgsl
NLR5gND2oJhLLYAOIdP2yYAu+zlv5zNQwWwIpITvCe8YC8eLx7IZqppl7lyJ
0J+VJw8ToUEops5oT1QTG2R5V9nezTVioF7J+VxUoNcrWUzoJXndN8/e2AwX
m+EfCn1octWi/pAwNA41mJN8jmvdFEy6AJAynOOjY8qY8uJF9TOu9+HxqGaq
a3ywGQlFYm7DqYp8f8+foRElSHf18Xd0XzJDFHJ3IHDfpsAVq+APf+OjHfxB
o6rzLrys6SDyCO8Kxsaqk7ZVRyPVhFXx8NxZGSrOQj+qW0nLZbsx2uF23qJM
oWL5OC5+OJUydWiwK3SQV917X1y1TYNiykcL4tw1g09JkhXxCssaYp8otcoz
oTV65MzhEqsCKLmW9xMWZ5fCzq2r4EwQqJDSFJO0UD7gzeBIp/rTb7QbX7ip
TAFnx+PSB38vLzItiMWSPMXkND//s8PXjGxHBu7QgUpABbZ3iZMU1TrEUvyR
ohEkv2spG+R8MxjSTUrUS+zDGDipbCH9iYkt7tYyPbbokMgxsBSWRXwp8mpK
EPzVPy1URNHofuTzJGnUeeZdDzgeu1ndihkUSnLu6Sp1HG4HjbGSmXFdaIgv
fOBgZYd9BqLx/IBuSygcsEo9kK3NHGsreHVHWTZnSNj51lLr7wvgY55/YORk
ujVtNF3gXi68AoFgw5o0Sdgnuk2Q2h/Ih9+mTw1uJ1eatFWqlqLo+QngEZTe
8eiKZYShq2k04KEq3HyNESnQNjwJgugRe5qTf7MhaOyySkvq0oJTo8RtQmAP
CM7XWKeTNySh44jHb1vrRUzVQoPdnvSTLwwaSaGYjqdXTMKgYmn30ZiL/Ri8
s+UhL4Qsf8WRncRUG2sbbUP2rNLX8KdjnnXHVz4MHQc3/Hq6vyHdP8P2Ws5p
VofBUAEqU8ky3nkEykKqjBJuPNb+rYkw67dBuGV4QHs/zuEl8jrq3r6FXnPg
UMTyZjfw+U1XguwemK0Cc3bGBr9Mrq6xlV8y/lzoHKJ6QKWbul1QnRUrnUz2
C6z7psIT7Y/D8q58ejqDtntrcyz+U4TTJkdCsmufn7mM22twDMJY3O9JdMxs
NyMeo0PCl602reAZB21K9itN6IY5nvLC0P01H0nx8mgRF9QcvlTv9MVbkyPJ
gQ9JGOXFL5vS0H4AOErEFRSh7CHpuERK6uZOyIFO73iFwXN/D73tT7idxl9M
e6P70HrMFsSj63xEQoCHrr1wcsC030fbMwDl0KPREKD4J+Hbnh5F/qs+TOFZ
1InRNt80e4cx4mi7Del4YVq6Djn8UMY6QMRrCubhRqZAcXOeL0u+qLLIjcuW
mVGgTP5rwj6dUVx9+0LaAipfnpxTNVic7VIFBl8FdtIVW43ajc/h+vVv0eHs
S6LOh9n3cdnASI2r5C+zSki4JBi++YMOVucE3prSAtSnBp+BCkrWv4kbf7ER
G1OgjXxg8acjQqOHmnXSsKELz69HFw6fxFVWeTPqsEoVTbtTkZ9BCxJJfdie
LeBgpNMSbYAI1jQKTMixEP17Z8XBRDYMqQRKd8+F8ZhX4b1ysDZfEuJ8X2fd
xKeeHfdOsIVg9+jB83xnPqbNZqJ4WxO4MI4NvAODT5evWM2Zn/6SZjIBXASu
Jhm3RNbV8sF6IkGW+0wVnBCuLqYPnC0+vDQQIFNmhtFsDJHjk6G3gxzgvq/V
I3OiUa5VFKDEhPE/3BMk97TBnWFt0Mm43f6/hoCz6kaR6YBMwRZja3zCFyiX
zEqpbhmuFnkrC4rZz/7bRLyerAY0o8U5+pi7G3Pu4dBJUZWyGS8TSBDQnISN
DyaFVQciSrHDjOeTdBDHxJg/2PfTta7DkTBU1KUXAioPmFlBME5mOF9vPhOx
LRT4yrAKzN37wc+JIN7RI1MAueNsREvJZuObCjec5+xPxbhwh5JnwowEcpt/
z9RWAXmsT28m1AvpiaE9mIOwXPyAcUDpiUsNII+O2W3I5OYdEA1vlyMCAIKv
EZNuIC70FzfsnYEPz8djcCTjWPigw1EK1rfsI4HeSMc9hjhqOQ3rRGYgTL9n
MNTmELTwapYIqWO/MWT7mRsCtGzR7aMqbgb6dpV+Ro2SNOagHxrxXhYD0/+e
abkiYc8URPA4wKixnamV+ZRxOq/3s9XhZ6vDRvuO1097sBTvi0HlmHw23iMe
5bQi6ztl7nArwGfJu5etIGuLNgPgLIcky9Y9Si0Q6Z9asS7jnU+/Ixz6dYhz
6LAUUA9mCm0wXmuMbTmSbb3amNyy+F3LRrSVSUlHsBwKwgexQXe9u4zFjT2t
qafj8etKVN2Q/hkZaQjxGom+YfmKBFvWbGeEGbpeUa2iWnoYxvNjSjoOxaFm
kjutJ9avXE4G2YxqNhwe/cdDmTRSqG8em1eKwAzNZrbn4NntxHaR3O1loE/r
b0sG2CjpBoj5E3hr7aKzUu5vu1DbC4KFskwqXTGB4QxGK79cfNdyqP78PM4l
2q4438nO82dKccMR0o14BxpTF70zrczufEFELCu3B9CLm42DGTRR0C/XHge9
ggekXQQfFtMBNtIzhQ+rg6Kh38fXXmN9vRdjjAWcaRC2HCQCrLNRXOqitYZT
CxrFHTqQrTXvr+v5onbRxxeGtXWoam7WCjRhfSSJ2gXRpOvJlD5ooQUNS4u9
/YXkPNSO2WSJBx4zPAcV1mIPsOemP2dsog+0L2fWJmLgvwChi/aNCjAeiXPT
87toywc1aq8AFkjzHG/cj4TwvU/86umtWloxcvqu+02jBSGR9NfCn/Hm4FoB
8qFiC5Tfg5Gzk+HxC6O4gPsx7ErXjkHcibGBqW+McWXWqLqCrKr/C4cnqNuH
WcBMwTb8LqfMRt5Qv7E6ri230m3DFUMvJe2C7PHKf6pYh7nvadsZOszZdoYG
I8FL7lJVUPW2CY/AZ56TArPtoGUsSWabb8Ekxl1L1HwVv9GOtOhhXMRpBFOl
6Ir/Chy0qiNWYlOTrWmskwb/mKV42bugYCjrvVwUcqd8cnUAsH+CZcK+JkYM
Ao7Luh53X9AXiE5PrLM8oyV1lIpBSP9T1x2Xloz7wWYJs5c6qo1VA7Lp0f2R
++RY6V629zHBubfUf+j9P6OMED3jBlIqg1ExGcHMB2Y6JLplVw3QeC1d6Krt
xREQL2rJ4LalVCEbQMhzdLFwHJU7a5A2OwBkxEKjM5Hm+I4/3CV1Gp9vPCJJ
fjqSPpLd7HsLINZiSuozopCQ1/8WFhXcpFzIIZa2WTxhegLVu5gs68BzkgOi
Cs8VdxG9NJKr/VplSAW4Od7Yk21Aq1pF1gwoNH4wdyopP3Uglhl2b3LimyaS
+PA4YBwb1xXccbwjTgdxfEefqEFVuHS++03L0LPCbZ88W+7TFs8SYdvLUoqR
vjtQFr0DYQblWOfPD2TL10DbQZE1IiuJwoKhd8DDV1uM+xoeMayYwSwhLvVj
m4z8N0crLIyodYRcemrM2L7rQ34c1rPT/FZ9DRzR9Z+jC46hdo099/y3E1kC
v4hVdvztobSbnALb6CBIVpqFhbn+2eJrxyVu0XFOQ8QcD3eKNIUO42C6hw1R
gW31BSnBLakX7dRQvbN5FGCAOlJiuF9XyFqFeFoeZ9CPivlIjlWXc8mi5oRQ
azQv1OcJwaAdbO+9fpAVwjojNVEnyvtEVj55IXL68X9dRhubCTeUCzNBcjOd
ZpVX8J+aWS3io6ZK1SCY7flE/ov0v6D+oopWebCizDLaq0R0smuycTTfK3bC
dbpUQ/NwJiiGg01bPW59RHfdu5Xb/iUGodolRAv8BP1iBSvgcgqPGY6rQPWn
h+9axyNYCtsyUurRxAPQAhRXm+igs4TToUtnolwH/JD9xVBLm+X9MQ+AGWjb
fphRM/4Wd6vDr2djHEnyvl7WnQ1EziftL/rAou50RgBZbG+uHde8sgXmQx4x
3xSydbeKOxgOo+t6tsUZk6kVsd1RKc7j8NPPx4+/XkO3z+Vh7fE1DHjV0Pjo
Rp6jyHI/Nzs1xqK9iTtuQAvyXxiNy7Va3Ut1v8O8szDBqQRg9j0cHPVdTd32
37HF/zmrbx+f+qUDfxbEPL1oRsxbglBNQHl0RwqnmrI1xzWLcHHcpNuWYLxh
DX0IVWmK8CI4SiHFboPl/sqnqvM6COyvvHDlBbViJ97xKjPglTyqd5UvyeAw
4FpdaT1iq7pVHWNOxTSEWn4Tyetp9fojS+rgiYUMAH3/o4eU2/TYDiN4byRN
Cof6+6y/B+2KHvQthUmfF5PmGDlR3ShUH2t6gKqDBleMrL5plIvAV+jK56h/
fSKA9PxpWRvYVFs8m+TQVdx8L3zeqnNgnmlS8HZJ2+zNZxFlwwHtNP20wzil
Ax9iA18vOnZ29fF7cSWQg8CqqlqKDfRNpute/xRmQBmwX5IZ0jmFBOegOT4O
Zh90A+RIzzIdldBJLM1zxpi0yaMVCU4gA6iVHn1ky3aiXfWR3L1Rj8FnurXY
xsV5RoFkWk9OJokJpGwPJOvyyCF5MXXKMSWuygb1irXcqH8KCdLMs1P+Jnd2
3YV0f5urgU7apNRhZG62HaPDA8CRBPslnovEBED5zLsAWXaUIMjeIwwEv4t3
Ezl/NNChMioVBowBepz5iyefaBg6xBgO4RzWLBMyq0N0jQHiEHLtq96VlGID
dWP/5/+dUnW4GoqYDmTPm6cLrcnVx05zLEiuSH0MCb08Gl8iZgvgqfRfIdtx
987wrJsZMQGGoy3e0yLuMcOlRySNMfYJCJc+qlZoj8JwbHB6u4bi5LgBve/0
s0o6hecaDH5iQS+TSAMY2bXczo+9XP8GiKqebaTyNUfY8OSbuMS1CR8piJEg
y5aHkVbRKGiJr9VFW43hxr5lARY4ANDanu3Gm+3i8VTsAV1K+g5f1oFbeh3i
Im9I6caVp1JmuL3mHzfD2Yy2DafwS/h1ADc1vJr8BvFtmj340hfROSY5hkY6
fskpyKGVHRf93XPJoJ81zIEswQK23ExYf15psp9aE7Zc9KyVOi0ki6uXmySZ
zn5DtwV+Mu6SffyOy5E+tHFDNsynb7kN/VEvhdTnpMnBBdWaRNLigAw3qrvp
eNlyPnUjS/4/MUzWsRUUwHP9lvKTwSIQya17Ipo6nr95eNCiJ+TrTEni6x6i
YP7UzzclxPE8em0NinaNv15Bz4mW/b+rjRmc+cbtccLfmAjQJpV09yzdO4xo
CnqG1FXQCafgwrGnpHXnL7q2/qUpdklHx/bjsqjWL9fDFVOzsj40eTt7IrSw
ljaMPR4J88RxOu4NpnFL9kQayMqSbKrzmCoJJU6jOuuJrgbquetJY4FsyO3k
z+kw1AcHfi55ZIvTgjXBfIfTols1udFG2qp8GqP1wAiXtkUImQswJ/cdnQmh
wicS5PZjlBt+JKNBneRzeonNOLg0tyDhw3YF+s9IpiYP7zhbQAI6SWW5Ap/K
PllKXTjtfZA/UkeCi/cr2m+YBvQQtMDrEBZblEy0bflk8k/jyyhiJdZ9QXTh
MybT1EODvKVVPsO7T1VfowmmyC8qMCs0Nw7lqEyT3LHH5E3BXDAvm2Iu9a9E
DDNp/dc1hgrL2DvIBuU0qOB4CyJgDnlBik9rEnCjBu0aRv4QvVd+Zw6Dqlx/
zPlcFavQvuau6VDiT5okN4Lb9X+QQRPYat9RpGs7XcaKoaHvf0YyXrj11iy9
lXO3VuFx6eMBywiLE7cPE6PTNksZ9aXfmKcgk5tNeU0ZcIAtF0GlR24ymld8
sU4HzrC/y4Zmy6VMw0gfigNEEcnOdqM8LbPSzoTkzGV0DvH8SeNnM5Rlp2mO
7ulfl1nNGxm3j2C1HCAd78cE1SbOOVz13VDmikzMPpGjvGX5GGk++55ETtIO
lrIjl1UaeXPZAH6E7+tgnq1Ubyv/F7wgiquiFmuGN6F5Au7MbdiZdCDAzLzA
/pf5ZwAZtkaa/j8Boe9Q9JJruMB3+cw7xN+Attk8QoNK12ygIyJ9R0HxZyhR
ipbSFnnklje5GvdYPGB/0c4qHZWOdSUPdMnbYgIzFN4akydFWLjUQLK1M/ip
BQHTdePwO0gA+gZTiq0t1f4DBA4/cRDOj3aZw3FhHGAra9cPdEDzKGZk6ihz
2wSmINW6Ewo/BOTBioORWFLn9zr9DQyjlUv8eE5fyJGaKzEpNmeOlrYJRRw5
PZtdItLAhztH9MmdJ2KsYjYS8ffyWYiIcjuyVMpoaAPH3uUGrgOgJawc7KHO
gZoLA427K8uOqyd1gaeWa0yME9xHKb3oYLvPdxhvnk7U+Z95xPRfbe47rvaS
FSh/l3qj19wrfUOeOjcobTV++WqEyQsOtKTFZ5sZDwKeCKvgoqsG5nPK8xBx
+c07w8bp/jpJ6prgD9u8qF+2OQuyIJYiM3/Xl+2b+JDRUmHxVJC08F266Rdg
zyHv5WMcNjTRtEdmmS/AzJtt1WntyFNa8ImjrpBpsN8he9++iDvKC3B4KiMh
X6bt4JA2a/kjULbcyApy5lEjkwxSCY0t3MIfL+swrH8W3Ncf6feCQnBkJu7P
RYdLNGliGe/NX+Q6btPQjzzrH9vME2bWnKCqSQfKZXdHAg/jgt8v6SqhTQar
iK1TJp03NewmzpUWZW5npo+2vs2TfNiT8cqnsUvfmDeq6TxKq01V7rSDR9a+
IpgIxsmCEoTM4b0nAi1ild5OwgdnfyiMhK8h4Ze01UoU4rAAzYeJQ6dxi8jy
Tf4/OmI/aA4abEFBSjdLYn0iwd4VhWCkj/54UVo5BtyubuQxiRAPT/t8Kij+
3n3rtiEhRVyU16XME7KSmcINXAvQLx2qq5Mi6OWMqhuJzxwOAWCk9z8eui2I
wzf7REa8/qf5iFoJ+SrezafmYVioXRPddmHdXJ88Wq/DMO+H47E7621EoFXw
Ph6YK2jr26gGUMVguu3MNRN8o7AfyVXpBXjmGWQ5GGstsNzL+gzJJui5NpAs
KQS6Th06T2aNkA7M/Ii9w1Y/APvxy3Ud/eweQGxeuLfte9IU98i/ZOBWHk55
jtsZFG9CS0XJiQhTzTGvtGT+FydKG6sOcJJnQkRmHK9FWbc4+DQAUWFqaftb
KFp1pNMuiU9h9og/9mRpLknLKm6f+7WPtp5JCnzaHzVAffgKa7WQKb/b996a
/53LCaeeMvQ2jdPm/ezludg+eMVEmGTsgLxgb5PHdFvXYJfPXEr+i+QCvGf7
95mICvcSccuswuFHn0ChIVdiw7uVCsWgYVzlP79bcGCzRZ+zun15hSYe22VA
cwkqwwC4u5fGaGMhgwbdymBVTYmBdSkGFRGEtF9jY5UmjWh+LivpXgr7HWtJ
AcA8jGy3bZG204DcgHvowh+1tyq7QmwfUEnoebkDm1EPqOnYDn3h7gL9V5q3
7OeNGSzz6j6lglD8EyH70EYZNGwcVH69m2uG9iahkZL/cYru2cTbtWtB+XiC
eZV8jeatPqs9FkGM2PzBPJfOlyaZh4EVwuA9t5ZBwi/GPzxve0CDzyDZB9Jh
wmu+xo42Oy2P9ao1RF9tCVF0KKbGHPA1J8m544h5ArdzOGhgy8FLsGKMdFQe
iZf5+RYIQ0SY2D81ZNixa7VrF2FrANBo5XzKdDVTrr5Et+Mteob4MHirbnPX
Ff2s2QuqmCi+t5cOXMbhKPy3BnwR/kzHmEGxj66MmCUr0S6WnKejwy7M9J/O
nM+dwPI7Ot8bTfMXtvZ3PDp2XAPT80CikROdBkx1/PQWtkNOMwK/0ZJ8UteG
UhKuyRmRVlVA4J0Id4LlLO09NkKxt3y6FFXqWoxZ/UnPzf8jyJ1Pzmpkjhmn
yhgCm4OQEiiHBS9IF41HYg4ZCQKIQ6V26MEI4RUDjnXzPCnNNbXBobksthia
jdYzhpAPWyV4wqTFKTGW5Jrmo/1++32q4ZVGvdxvyAwr+TwaZMT3bDIbaSmt
cYiv0eAaCpIXWc9aCT6Do8+OC+N/WQwGAutabce0/lP8uUGuLl5pn/3Kohxy
ngKtfAyfUVRbDjE4NKyvPX+tGZD3O4f0Va2iyCYTNyQ5uowFHdGrnb/TH7AP
kfHoRQuJGmGZtlekwW4VYkgJIdnzXzg4Y6jWYrzVZRa4CsZW/6IK3sjvt2QU
csBVeJQY52BZKFbLMP0sGr0LVl3LNEx0kxgOizJfav4VvmnH1ujBTpxaYcma
IvDUOTlvNXQoQ9A/SeNBRtnE9pV+RAwiGAdbsrFBmLaYr5e/472oO3iDAM51
4T7VbeQ+VrBo8H3D6NLrEds/6gEtVHk+/6p2s+sWi+Ksw56MhFlGGjQVEQbg
XioN1qZjsgdz7Rmr4OL0KsqRYttp5+fDqhRktbCGhR3PvomxV/CvWcR2kVfG
j+CFnbzmm2BEQ1PIwz0q+ME9RbfsDmKVcoPmLxQEbpVX+At8lB+RUQvAVFyo
dJNbLv9h3ZKtzp9cCQwTYXfI2ttD25iOhWv32kQLH4hZwr7GWzM4IQaTtPDD
94O8f5Q6tVcb4qDiSQVj2L/rJfL5epe25/7crWXeK4aodG7Ha8MFbImYlqxj
FmjgdpPTFnjIenuRqVoPRaBYMK/sotwTxPm/rYDUFtNln7hWPu9vlOUgnIHu
k2GafsRvxYzvVTNWn/TbqJOJZNRQ3+7SCLC9sL0Hj5/yDBs6aHssUe+iPsAl
wruBZ4DEnzmKP33eqhl+1aA+mPH822qw7C4YZsJV9oXg0cE1Cc/2xmrog0/L
iorTQfl0EJUFbPyGq0dR3UzVl3B9LuDSjJhLqTM9mslwnLjRzETQwIulv1JN
z4wEzkjX2oV7DRSNMOUwGUB6OWu/k4lmKxH4pPMEq8lkN/x/HIJnJoUwhJAf
BDmz+5NKkjkPCFNqkD6Q3eber/QGieOZWZOBiBvyANHjW228mRjvjAiCXG49
eGSdlDo+xrOORkn+ytVy1zldcTqLJIrojnafEfjYaMrADkny4GLaxQRgC0Hx
VvD3TtqqZ6SyDfbOqlFJyeQW4wXBKvBX8fFY3dTaoPv88Pu4o1k9JVV9SQh0
T2IOIHNBw6laoJkh4xtH1Ur1bWBXSQ61ChcKXwEWs9NnnZtXeHNGICWLx/oR
6ygzSuoD/29bHuYvCRYekQ9VlKWy1nMWj3zdXbNHekpUku9nq85NsGHzphB9
mLx98l0k4rzl1p8y0GIa6ZRIx3mxYNb+UiBHj3FFPPmev2X1X2O/r8NfD8of
wJYf+YrH2Db/Kiro9XzfGfwny8b19le00PByw9hnGTtlIZlBbx5wr4lKfFFK
iOu8nDl8cT8KtX3i03Ks2HaL+2DaVmkXZGCAm8TpJISUykLcFJvB3CJ9bsih
JtRVKkl8gzvUJOCw55oXkPcMAIXio0Zs52L8GW/QB7KPhz5E6EqUEpkj+Yel
4Xgix/dEk5wNEKb7ZAi4l0Nj78/J4NipxSj4n51OVE/y3J9fbokp49maGpER
xndgsYRDzYNF3X5tOqJENsIjbGq34nmoYZTD/6umEYAEDTAnoExW+odUcjm7
15fqDa5mjeQ9mNQor6La2F9YJvIwMoI1/IXvvQE14HQ8EGok4CJYtZQlb3nv
2KTyG4964IBn9i4wPWbr3lzh5EccQS3llBFRH0kq/Y3qsD6sKVRsdl6Uu70A
8R9Lx4ggNxWS/Jdns6y3YpWcMEyd0R7QAr7XZUiCoBc2uw5KqzjJkBdAhTmx
+xw5fOguDrrIZxdwwZkhCb1oy2XYxnY0+K3KK6aFabbkSp4+FGLWy8k00bTg
zI803TdFBXPL96WUQRwMBD6Fm8VEei6VH/zZ4ed9qoOwvZoKZXfFIdnv1Z2m
qDhLCpGfIou/h9GR/OUfrPUoJjNg4K9e2uZcGqpWzi4atWOl+yv7xMude8vZ
7fSZVyxwVRJMFTjfPIaCQlhV2FunHxapEGxgBzX81ziZW2ilaY2LT+fj3Hd5
+KT0tJ47D3R71r09O1p/4BN485w6O4TxsRUWDTk6KV8n86tBLdXLCKjo542R
D7I6z2qc5fstBK/PB5eJd502sTk5xLTvKj3+VUGCDmLBiXbNJAyr1q7nMjoI
fQcz3UeOqEVtCbyNP5wDBa9taDSla/4xuG2Y/YQIDcsaDrURFg0pdOAMJQvD
MT8IoO6V32NYqAOit46P5uiKc1QJtpKFU0tE92wRHUFHW0VSRxRxGCN5XD41
gKpjrHA4pYuUDdBEREqI/r94fDev3pHmXrOoqg8dQZWXGvKpv6gKsC1LjR7v
nDx7OMXmhfss8WHwOSMmOT+AeYCSsJ3bqhJrjJrgZx7vkniQ9va+EfC0qPxi
JVu8RjTIUP4gQdWrTtZUBSmO3bpIgiirJgRDwLhvJOlAhNSvWWTAePpnwDa7
yNN5xkaGj1Sq7aHg5Mqhvkx/y+wDpndlJ1ddBMbu1/VVC9lk87Wc6gq5lf2d
K12Iiglns3WHQlYYN1rXMmfvrwKbTVF+mONEr8JM4cxtPKhJ6kyHnkL/YwuN
+Je8VEcj/CdblX0a5OjJ6rahjvYNhhTxFtfxFlKSOil09jXL1/+H6aJkLLZ+
g4/bIWm3KD77zFOXH75tfl7O1nA2PSCNSzzqu6H2CgNoy5UyOy9G1IsWlV9k
nuvQWjpscgzImKmtyCP87tzIlKWhYyOUEyLzM2cqlIsyx1qr+aOhUG0vLpPO
cNI1sK+zHZh0Cc2bHrJlHBt0S7RRjtM473LbHFfd5RLV0MtVNJr3mIC2xS6g
YUir0f6zBdWMg2zgAwf75qcrLRkYGb9se0b8ABeVl5Dg9aFPiMfP34AzaR7/
Ub3R3m7uZq3IoaTTCQatrgtdMtmTPlcIOwVf0vx/Xms25cgGnLongAlELSFV
bYACEln63LfX9O4autILgL8FaFG5t2nlTgcrJGMkJjoqbcFxroRo44WsC5+6
Gf+8+AS8PyG+4soGSft7yM/aGQub4yax5uVyY7554pmeCC4Qi1/Dr+o5XSFJ
lZNkdSbt1c4Au56FI6Lo0UaJ0hcycgp0X1HPYxeESyLMfD5PihI/z3Qb68AN
vo7DSiREtTyDbu/brWuyHNygz8OekeeHn8ktp08GCVMm6x+7wXng+xEN3wTB
qteAIYRLLBgdDZCry0NaBRwSwHee5ylYAOcIkff4eMji7lc3JSh84vDjTG8e
jaomlI4Ma16frEqdeUe4As9D7v6AIsDiH8FD4LcjQP6vdjvVqxdGiT6bXCBE
uzNGMtfPuTwwyvzH6n1mQvUZInVQZWqCpprF2am8YvE3m43UrPgHqtNIZ22W
3wZe+WH193+4R+xOvN7OgVFG7ij9lT8MT84Ln/CfxClWh6U53RuAsOBpO4PY
K2H1+gykRCQ+Mp05ArhtUjDFUOeyqRxQFw/qKjEgmfLGUZJ73UofERZv7Bnn
XuuW23VMLWAHVmSh2oCyKa+0mr/q9hVrynyuSVE7a7QWsYlCqs3T4k1/Ny8A
aaNV77RkgLsAQBCpfGFFTvN9sVkxOQafLSB9SQR0YwV0unuHfjAgM8GhMFzr
VXvjfV03JA9RhA2vKp242riZvpap85VaCLlceC5eQMIwXz3A1RHG86aOSpao
V7rCJd4EZg9CEUHQhZEExO5kYQpzblH1ATkaAIY/xolYoU4icF03++zZLI7c
s229oj+m0Ohcom/R0iuEh2S3Y/ikeBC1uYX5ncJMLopCzF0v5wFx/Vt16rWs
XFHIoMf2KahMq9BGQmwHfB0j0lhz5UraMJV/5T6jFljFFDL/wuqR/hF8Caaq
TSEq/vJSWDK33NkmG1CwW4fA0sQWXinEiYVpmYG5g72X1f8y6yrgriBDbBw2
aL0Q6eRMUJk2JFNtkgvCEQ5HMfdLXwuz8L9YQupV5pyYCjVNgpDUeY9acmD0
fNSOUvpTtE1xKPqUNSoCVRYjdFmyBe0kUy07D1spDTxaJRG22nbYnrYxtPJu
byB8prZmcG1dzWhFM3m9X+tNixYByzPtoVgqyfb5yYdPxA61xTcHEf49S9c2
CivdBUgMMlceK2vCTGtzUe/36SyuRzNeFuuTd+1bYWeNJelN2JUdg9NWXnUg
2/g5aU1yC5JSr9MReXdzLhpGvP95Jh1JcQaBODSL9GMN9Eht3fofbIETE0Qy
/ylIiLGJLFQudbfTrGAR+ZUIE9qhxPn02dwW4K8vfXJQgSwFgwaZhV3IPrSX
glIzd7+QImv8EfcoiIHLmprUY4YNWGS/qHhw9fdXw+/UCU6snwkxAR5HFpuG
YSBF4H63ZhCEpIx4+mmQa0VpkqzxD/CyqcFi0zEHKewbBqH4E0k9sa0c7YOK
qocTjJFPUsb89UuU+RHFsQG5argnAA55UHn4a5YdYfFlIyq0nTbsoyZwwAvG
51TJzo21dwoTVwENSsRSLhwWh6nmnCKcoJYbwV0h9/HfJm4FSnX2fNENX6E4
deuCi+lZ5g4hJxZ4UfwzYVY598TWiIR3ztQYXmoRocuZuHoF83dh2omROaGQ
hyIzhzba1QmavBk3wuqbHsSfZjHU7XTzBUduwLyMDIjWx5zY0iLoJY13PeyM
ue6h7p8Twmy3qnMbjyoQQDGMpHltFwhogk4vrpePLddDvpZgrqHDwdHLpOeV
SbqXljN89adX74qXCyaxDEYpMyhoM7NScSHFBu0+eqaSHMD8FKY9JpH/t3C5
sqxiG1UHQIbS9/lzRHwoertmnwF3Qu4R0mtvB2zrMUvihT3nPxGuUg1LcyTL
9cyh/YUA7wBLM791dGcib3g/SGYmta9tbzv8fc6kJICpk15iBfVgt+ij7Ckk
qTmMcOPnLsUjMbEkwe1eG7t4DRmtuD24TwSi9vQuNAOH2/Ku3wSY0QVHZZ9C
AEGxpTaEGmiJPLprKWvps1zEsesyDASRcCc/K2vFgB1aVwnI6jEJ+TMYHZc4
/ocnKSEAZACJGUnxgQEdMUVBw2UaD1jmsguPxAmYlZBvRFfFY9XgOFUt4lF7
DzzmvC0vsCdc5yYWE1mPTYjt+iO3aHvCsLI0XszK8d2W+yDjXOYnZ10Ut9EB
NckxeAamkUluv9KoYWQGlXgW8P63+PrLcn64Ch3rEND7s7s9pMwMSuYHHO5c
VARmN2RELDvSYcBqnWktUGRipPPyX0aHQDMkkpaNaErh8NYr6wzoPiFMnB+4
nvmYSYs88GluEVMEIEBfPKd8Q33AeKbUgxFmTr5YCEv32ZBjIo5GVZ9mftUw
nc0lbD/hqH8FPMJtB/itiTljFXariBVn83zzzcIaTAJ9V0GMwCyMqK3jhPA+
tnMpw4qfs3dgEyLS9k+1SLTNwCrolfSQ6bR2GXFhlv9e2P7snsEJHNMRVpKf
cKHEXpFHcR7ma9MNqZoAn/JbGY0qWUuaRjP3Rm7ml+Oca+tAhfdYzgMS0zFE
iy9zxJYlbayK3HS5kZKT2uCEb2MYwMDdUmERT9gIcYbbucYNk8qWis4Kfxpm
tZJhuHLoJIS3/weNvAfGeYYi3qIByrBWrKGwcHBT8Ctk6S5B1qnBuJ4Cfq3u
9hSadGy/FiIS4Lus3iZEGI8r0d7uxjv3O6qEnjrr7pP73F0lFyuQqA4pAh4b
fAGZUMPp8mtoZegRlji7uqgLgjMviGaN8b/1cNQnBs5oUDzv4t3xvBS8O4AZ
MgSlWLexA8mGf3xbhZiFMWYqJtrt9uLIA/GRLnfk/9Q+SUekEw/CeomDBwsA
ORLSKVpcWieHsZeSH6/40puEaI19mdG5n5d360zYhkdoUbpV0xPKWNtcPi3h
jnuYTCqTfXsdenGcmZAMx5E7uzye+lUjKE5OL6JBmVrEgq3Kp3t0FLcZSmbX
h4OD3LjNCJVNyxOtKjCnWsp84p8efQkSVdbduxXkpiCYVBv2p2VdlRH4w7oA
LPMqjv91dJfenSl4TQTUtAnY4OTSq+7mzQc6d7Fgwx3tFUgLtB13zjF/BQ0M
R+3HsNmihDuYdFRgDlCwUMmGfoVP5c9YKTq4Q+fwO8nnsSW1B9d641xbkZAY
Nl5xggzMzIkp3JNrvlpkkxmt41zuXValzT6wDEQEsdzlQGyPG2vhF287zE9S
soHz+UIMIEaqq/nErot9VcBOzN8lExNKN2Fq5kCK5knevGKATOGbrEokPmxf
w1XMrVCKOX3o5TpJvcYVz8ShXfAe5bC57+9QOjjFex0z6RxqHtclweiqV22M
SWZRH3Po1Xpb1DhGtJC4XXXRr6I+Ff9t8nGdeoiMj+vmpWZJoxe4pJdTxtBW
mE1bZt9xHiSORqcBC+jH+t2dJqwueGYwj7hyTvwpNgzYBpjEyayfReghT4bz
ML9yh0opSWaOEmU42vfUmf/4b+OKQ5saZp6ymZQRZIlGf+UfPbUHzq0+3F4j
RLQ9rOctaHHd1Vdf1z1Sht3ssEYsT6YoH5xyXtBIOej19ZtWlnz6CVukJ5fl
9z3EMG9qlyqmCx5a6wx3SXdJ7FmVhsdSa2saekDlg/Dr1/usXG3s8PjdT1Yl
6UZ7v3EFvGYPxwf1WHgp9EMfoQGJjDD9VQ9f3fUQxyYjk3EBQVuYnKzBRI+b
5KrZ10ur7CM20/2dwUdbIyoWAS09/bzssF5ijxDkReojpD7ygc4fzD0MdpNw
J0QPeytyLuWKf98YyNM4Ej/RJ5gx1hiAWIi5zZ0oybKSvkF8rxb+DpXQC/oo
5vR0v5r9Uy4DeUliWDiPO4vuM15Fge0xSWG5ElkCQop4gd1eyB0QlZNgByJ0
AwxC861oSxSGYg7hlic/t00BhzCtO57oSvD53gVVxRCE7aJB4jztUXkTtnEn
hvXXgMfkyaUswFJjKIsCfiv1rObiyeqtTPManRLlqc2Kts0ntb0pF0Yx+h7d
n8jxM7zwgkHzNFl6/wrgxZaRVaoJPjMHT1xIuLy2Hyu+DJSDEhZGWi68a0HD
tFOgPbFtoWWVaBTXEA036+9zezh2z1BNvv54n215Gz+ztYwYTYEAunot+YZu
kLYFh8LpHHyHitUnny/q89+npF2aixYzvVrkGstCKksX/Z/1eas/iSS8VU//
s2Te0dY0VUihX+LFzOGtbQ/u2aPlk/wK0Ji0+JDIlKp8Qp0PluRwsiz8ID7a
VL8alnbsWwDgr1nv/iHQobZJA32C52dQjWe51dRUGgZ45Do+5oOq8Z28swB+
5Cfse1KYOU/uEwwRJXRoYXYJk+ouek/7hWCXf7L56YA/o+uz3G5InJq9fDlr
aHPYajOJanctdZLPQZiAu9BntK2nr/PNY6GXYJWFQYBFouELvBxScwvAUZte
4YBnE9veUETZSEt//cHoQv9RI0711j+CHpHZrK3iogJzktHF+9NeFCL+9aRT
5TWbdquP/YcliHctPlzTTQJEllmxbMu+OQ2UVzs9IwC/xP8dXJneEMN963uN
XkyPjOPZ+H0yWn+mZ1Rm8HL+ghiCkG35tbhpTBFpQ/TPBCxZ3vFQx79iTuZB
MNW01Jn+S/RYuySdl7CItEsqGAqQ57udfQWwt/+a6aL7jkppIdmQoM6kieRR
sZQRW7PgVcFL7IgvIU1OgIY8BPB+hY671GQuLfDiZYbeXM3gjiMW1ZpLBIww
Zm4Qnbz3HTECQgOQ3Bj+okfqi5rzbcZdqAzy9MawEWH3GWvuQUj7L8OyFzWU
kkFQoAExWDtjbVTqsYh/55d9YgZQj9eEaJS3WuZHt4kx5C5erholwPg5AjiF
FgJUsWh01Sc4ktG6OAOOUuImZxoPP8nXAeW9FJ+nbLMaaNipwk0x84KovO7c
8UCN5oH7COlJu20Lm//cEU9FlHml2Y+u136AnADVKlho8b6f/7XZ5Q1/czdI
ewpUkxx7a7G3BysuPECaOX+s1F1nr6S2pW4ZZQr2++cfClwnVSj2Y4U3X+jw
8RV5nTOdlibX+hyTcDeADE6K3rkLPqHH+QGvMaf1rChIoPp/+r8z9RK79phY
oVuPXLCR4WHlAtLVwfEiHpF8z4/CdgfDwDZe5LRNTvoxSdI3Uh6NFXOLIRmh
sfiHFjg1cZuffkKzYJDG35V9uIBMMk56pkRJrC5I4/9r5TL0GMy7XYpmBZPp
9XzwFsB7Zk76ZoZ9rWvnjHmtquaX4mzq/B4gdwgjqx0JFejQRVzoR3tS62/w
4Cl6qLo7SpJb4teHJYLfisTyWp4jb8q9xrgtJy/Vh4297lonvltwS4oVUoj2
W2FAerfFbaWbVAXmvlrs0zEmAmT88y0p5nzAjP4M8kJWRcHPst7bXK2wvhcq
vpJ4lgEueQHyDmRe+1yQuqEi/R7AjIGuPqJ0kzC5Otvn5yiz/6GUYlUDewbi
hpJOdVz+OMRm78fff0NfQ4TDJFZ69up8OOJ6pFdz5G3Fv9eUaYil2K5mfStW
kDOwis70tq+FKHr4z9sf8+GwncaZD78qf5K7KtbDw4+dgcvDP0d1E9mRgTuB
umuBp99q3jtodoe7gZK9HHxlRGpnyPxCkCT2R++DyRMOsh9yu3qgCgBo87WJ
4aSOMP71dxQ1RidIw/CbvYvP4gU4H59mEwu1wfzCUidxQmZQXNM83uT43f0L
C5wfgKMEaiuRxNJBpUPiyv1YLvd5/upfXD3wMGan0E5BmGnyJet1XJVqDebm
mXSHBwx3SyKKgCsIdM+aK4FN/N3jpKOuDP+kE+LDarOQQlEo1//ZVmOZZ7/3
h7enMhSsTIKugos+1mOboTN4JrvzWCswwDU2uGK6xNb5/FmQ5tLYpgU/1vzM
lUQ8evgL+2cKEg9+pNKVc3YnPtwxwSxJJba2HbQQVMiUGPiWmsElCUJUd3wp
JyM0yzePmCvtMk2/HBQxpNPNVpjlftcMxGa0YfN167qxRT1ZHv6FE0jmgEp+
CX8a2C3ddy6VMyfODTnyMfU24ohx8Otau8E4rXCzZzx1Aid/x76Os5jTwh1s
wdQFJKGY6hh6l7GEn1W65BOEufHjTNdsiL3wCxpquUeqtqAad2VsM2D7TBS1
utGpe0UETCOKDB5PB/o9wKsBLACLkj09mgpqBi6CdrWFyfhpfnVDzXZzKxC1
rpamN3SlIg56HW/jN+H1KviX1JBMpQkNpT+fNhFTpZ9IiDz8YXe/gL2Ppm2a
uRAicKwj2wpj2HaqvdvGU6FJPc48c0JmlmT7X29YfH4YS3SSuzlyv+dqeSwR
MbE6qNUjBG768j8sc9maNe1Bru5em6yS3aHm/V0pluWWLiJx3SaAfO7tNvob
97ZzdG+craAvJeBm/QQbqvh2N8DDpkYN0hDQsfsHFRa7+2bCFwqIQ3wWsZkU
K6/Ga8sG3mKtHkbkVkIIYmEUS4v4Dh7Nz47rJphoe3ck9vbQ0ixnc4U9yEsj
+Cvrb73Y6b4hkhEql9OI3K/aiEOjypD4vNIU2ZldaYB3s7vmoO4q8wiVS0qH
lQdrqiaISORbs5wnzA2zw7wCNmLE3GmfGlTVHfIP3nfGdOFEyEh4AupwO8ep
lRyaEW0RLts6dTDSEXUFtGiPgB9LVkY4biITW+xr5BbNpBkiqn2ATwqW9dO1
oM7DXS1CsZgLF2uKLbQRxcORG64Mj/pxbPOnXPDRce3QJ/9uF8jR6RpGLKPI
YSxoxjcHIluC1eeeXTd7ttVGHO+NgmM81YBf2vIYq3TTQ84p6IFVjix+7Qxq
JoXiaYCJrotb856MI/mvk0OeOvXR9up/ckg+7OMw+hI3sz4vE4FezSwuEtIq
2if5iRa0uJQuFrHY+ar/lQeFAiF9FjG++DDocUIM98RCN0Zyk7yQVvmrfv90
TJfQxFDLZLjlzm2FMGfmQz7TJCnky/KoMYsVGxIK3kOzi8jqkAjqetroIT4U
QuilW19hiY/lwHEfpe6jcAR0lGoxeKsMUtFasmXkcW4bdJhz3MxJBQHxhPed
N5tDGWEYa7AsOqU7DSzRXkFotBwUY8qHCOf+gzEVexOpbqrqjV98Uj3/vIEN
tn5OY8THZwtadF7rQ4lJggp1wvCNQ/TNf0YC7cbU2GoRM83sr559dtKCPEmc
jV3k0+K2yw1XA7NIpdGqSydy1VKbD1lFyzFekbxFrG8X+YK3wULhBz0doynW
1vyw7ooHWJEj7vn1WZlBFpD1OrC4PrsJ4FYPTW7nCitvtAspM5INC32FaEIv
MaaPMosJ04iclcE0yDp1BIjKEGxTSIS7wL0FbpFzbSGTDIMnUMRK+0Lq8EkB
tqte5gDem2ZNSx6Oa8kVVg80b28UpWzdtLMq7FoQE1NNA2OyS8nsvGLEZavj
zN4TJQIbEE+kReIdveJXN8E9dMPtJhZFrI/WJ/j8VHNHcML1a2bSl700UDMR
vKUrBqB3RHiKPQ0t2bX6+/p55qDl8UKBWxIJpCUMcesROgjJDQlCv4KtszaT
VLnIvGeFt0UNw49xhFAWVy/lr4SmLNXCSbCX3clIfGPL2q+QELuc17pDUKVd
50+bg3IhjpzlVn3JDAGs+4BBLbV5pGGa97LIFQaRCvbIVR5f5GV8fJF2oYD4
zoYJr0YxNfJc1ZLMuW2+GLXcfrEBlh3eIMd+o2kDrUEv7oUhELxfa08WjHtd
+l+ooUnG0M4rHGlbQb20rBHv3m/P+wSUhD9rBrUMDPOHPQajxOvsQDPDRCQj
+yYMlnGQNVwl66FQO+zhEEn8vLLwA1y1ONgotOpB5al7VAwA7xygU7fNypYS
DcPX2Yg526KP5/ibMPHQvRKiaUs+0ukLisTInasiSotBaKBquqEjSx1bnDUd
80Z9GxqIJC9qrjxHEeh4QErc8/drPWeQu7/803YO8PLei4oUKPfCtFpIQ9Eh
ZSVHBVBU3fxwSAOVi2LqieGJjRT4kl0DccIFIIEU8WSTovAVOIpn0IBfcmKo
tFhKHe17XVl17ak2D3juXEpguuJR7huZuL+EzMvIl9Q9EnO3uncxZjGyODSA
pgkA64VOBcQQrTyL082pzgKXGARkW0zzMJKin1YZ6eLMMCoh+N9zlfbl8tkl
3W8BfW+2ORNrqTesuUCXVUKHnw7+afFFHPOyCqke4EQWwAqtMn/FSpt4NVCg
q5dVLaFdKhZCm75U14y+m4mIIxBS7jeBP07sNtXRm6i5GG+0zXalaAanUM5p
OebHyMSLBWrhA1QTaa04ZL1E5+f0bFHYbjXqRukWM+OVCqzlYHbhoe+Lj2ez
xyAn62FeeqvZRTobbcxzDFnWNR1JAuQg4Lo+ndmN0KCwtEK/zUls3loDFeMg
J/rfXNiU8Ki2ySNDZd5+EsFEwXvtbU7k1J+rXgelQvJBRE/yaHRfArT+pPpD
JXUU8unN39iAHZ8wh5x4A9qGmNFkuT8BLVGamjodlFVwI9z1/KqE5v8hX4De
lAc0DWhGXOsjuQy4To9BbSqW/M4yRQtr+wQPZ6/BpSf6cpFwI0QlYm3+9wJe
TdLil/BVaL9SMLfhJ/pv7HsOMr4UZ+sLBHZXvXGBz1hB8aS8rDMvW6U6JAV3
ige/gk/vvbDYsWajXo4EQrb/zpX6SuzOKQlREUos/IoYQWS2bpGQ4xORCIw9
GQEdLTR/0aUv6HAQ4MArUOwTN4aNq4c5gJMMTkV38lyX4YQORrmvKNhoYdlp
vLD2xLNfa9fAfqIjMzFIOo9JxZAj4qQyiIHH5+JcvAs6pfesloBM28uRIWB+
D6XIQhifksv9I9H805vQXcePzSjN8GHrwkLsdKp0tbEoxlJhl3Loc/aBM/rd
Sjm/DL4JdkeaAT0EVVm7J/P/xsuF6teXeiFwNwcdG90c7jhWQ6S+HcMpNERl
tTUInH7j2oET1AAaFlsJWZQpwPBrUXMhaygyrBRXLHOyeIMBJx/fZZx24sCF
5Ip0jyNYtTMtpClXcfxxnriyHv2/VKrlrU5VCbH541Nj/ZxH3EkLCvK/G/jQ
80Ds/mvXiccYAR9jAD4LXcqKu0tHQubolr3UrJK1rZBTaWJD2s8uTITUOgP9
BCLbNN2yFS1dRXt1SRNg/fLGkA3Ex4aAKKdWQ5NO2uXijF8eowkY0MuoIkHc
tsHkUapViRkP2G7cSbEsKZrwILRavbXz0wzixfO6/TwqVFU6kdxSpgFdfqxm
hMWkl2OJSEb6Aw6Hkia8W/uQ4Z7K5zO1TYtNsiPj8YSfaJDS3xjbB2foQFx8
whqkuFuSfGDPSkcwJdwk2rQYE8z/PZp0nt3HFsH99qD6FZB4PTOXbn+kTmvK
ZFqkNEf0rpi9VVQCZdbZlUbz0FuyBwIS1BsejNe3h7A6eP6PT1o9rIZ/tj4s
2waxLR7LKFB3GRltMDsz1O23AfLUkXMpPsP2rcsHe7t9CjnLHOGZZnufQk8l
vl2pBOuyGC/cehWpsPYyElefr+t5t4++MfaOA/KAyUaTUYXJg+cU/bX8flhZ
4lnF/zcVEYimjm2wu7P1YLkf6affmyQ5VPUfUnSWyD0qHXiGgEATJnBVZdmZ
4UJsik59QVgG8pH5Y4JEsh2I7kmrgJXk56oEP44+yJUQgoVH3DWWq0qvE1kD
cMLhd5hGRw541r+AywTWQpWGPHrFRShG30tmZhlxaAj7gvqd8EkwNaIQMQvG
qdcOzlAbGWXKct9mHHfI1TB5DtFSocoBfGcsCKZaGRPA4qx4pJR+D6vt9TpV
aZOMBLA5gTmz+4hVk1Ju9PnPFqYpn5o5W1E3RLKacVA8QmTdZAa+EfEaKFNt
oIYAQ66Z6jeKDUDzbHpA58EyJoEUOXIhRsaej4Q84bbKGj4JL0slxgJaB8V+
MgMQr0/uTFRvBw9J4F6ew//pSyknZNiCh6dIxdYMtFvN2hPmnUwhrx/d0nPh
Hx9B3UYbI1uU1s0jqC/ZBKFW9od4lFZR1Ipp9VzeQkogtXrn+8xz9/tKuLmU
VPAmGTxv+guGgaAnB0w04BZ4VVp6lKTu6vGXifctYw1wJhcYmbKpADxoeoGZ
jkicGbuz5OZ2y3U/5rBIpxFdVaWb43VkV5/Ae9hfIG8JEPLez9Zwi/kSWKrw
j4tMceg+w04t7E8N2g6wCpGg4rqwm0BUxOmrV/rpRAjAXploA0HL6IHO96yB
XOBumkhK6VhC6A+wt3NcO7iFeTSJqzDNQ6XtaV2mp9BVi+qqNyaN4Rf476El
UuRxLyRlzyZpB7dIeRVZs+wIRQpcVDI9TxpG11z8WWl67vl2HEnfQo6ZnT09
s20HMgCFCnURXQ7g8ftaeOlLctPQGB0ECpzIFWUXaQOLk3QQJ+8maqkVuNXY
dzetanFZT6QfyYbb/ACxvY+F0AeC9w3DGBHWdLC22n72w0bve4H/Sy4yEq3X
g8UWsZyiLqaHmiqzp9+09X/mZ7ssK8wnsD2RqjlORw3laZoJVNI89xOYCeKq
XbNluVOI+tGvwDMB1CXY8n09CNUzhmkwXep+k+b7P4OVZoHU1LC5532iNIiq
y/4vkhPQ1GNfl2DxcbiS1gVF9NtyP0VubbR+J2v9px/DJrH6NDPrHpPuo3Fp
z8OhCXXsMrrWjDXkHKmICJbX7qAqdwG+s6kDWE4T962L0MHVZxJu7ZPHHIBA
M3TN4UM1pFTsswJ5MnaSXGaiRVtf5Chw4vn+6gbkbzKoDe1bF/9WhjQFumvO
snnVTQ+8IX/7IAC8F6BalPjwOleaibYz3769+hXjTwbEIROYYxKPNjumuROo
JGo2IQFry/ROy0G/5b/dh7s7Pmy2YNm4DFzf7Iy4rnvkkaRiTjvV2D1PE5/T
WT+KKOHCbzzx4aUPLkEoVHggQrHaKBbRrpMUwe0NkAqx363ndRZZ8439U2TW
WWYvrTG3es0sfQWFyqbCupXwpX6jH/N8zSyQ03RNZ9GU53bRLqYjNW277RC0
9KdnyzllwaQRJW+C2kh6Tw/607MYAr7TRAT5KAL/LBU498IFB3lSgykqxebI
3rCFIthE73qZOic26FNwKGMx+GtDkx1Pr7FXIX9T+vQsUpcgfVY5ZkfYTPFF
/beCujZZaKvHaOnBcSIfpLc1jBelGpc5ti7Thr9vGMR6wRudc6R+R9G5U6ig
76+zFO3i8gwrbTDXxNJv1UEPzHzAW9gGAT+gvSJMWHrY1EVWF7brWG9MK1d6
fj9uzgTx8I/tqntXmLRPI27IY+/FwB6cOpsR3z/1YFJorzjZxjHPSyGHBhUo
1eigd38ncfTVu1NaI4a3hJHjtXuCohwuwPMvArsvRRY2oC4vIuLedarOBzGv
t7536lZkB0RTdHz+EG9txU4maSUrNnw3SpLH9B2XTabGhc4kNaY7glFdR4V4
i36izlzTTcyvW/1K1TlzcD8/opOvF14MX4b39fbJRU4KP0GOUWXYeNp7l5Fr
kAmcD/75Bw5x60EhFBlcZrFe9FKXG6hc0z2YEQY4ojvpKyymdJJL+SlYMRtT
RhiR4Qvlz9vcYg9EUVw5LwCv+VHBwu/ZgHFwG07N4BSgSC9Ad0iSe0kD7gtc
hpA2bAdVgr75daA+bp0j5R+E7u29PvQB/yLfwSLtPph5zXgL/sE/doaJx5Tv
p24Ejf45rsBQlLNlMctdGWDC4d+uoSVFK7y75Jrdg3l0tP9R6dttHaAR39Eb
hOAwDTT2QCQ36i/2BSC1qqdvxcYDDbzREk3yI4BX95Qn1RP+qFipEXAM/MOX
+Q1YkdMPYRfO3HKLxXt1YjFU8KfZll5frITxjaZLd2XOLslS7kLiKQFgljnW
3Zc3jk2NQC6uQOQ5hgVjskcMPnpD6qOBKA6+4iIXGLwCjQbN8u+sAvHTwCLi
mgG+SJPDcY9IQhc0mkS3fy7ho8SBANINsnCHH5Qxzz8NxrFbKVjFcovF0XcB
qIeA5Xb92Ku69ViyrML/WB5I3469QBkMYR+r3pdO2M7h19ttrk1hyc2d6JOE
i2ALijqmmDa74ORJWYomJjvKx4TyxDUMejOG6GW5JWYqYEWa6Bn8H0mixfrX
dH+0/5hwfZfG48WJK+IwkO6Bd6l0QcefwqldDZpqN5nJ/TIaz+SzT2OBTtN5
oZ0sQunkji37Xr9laB4p2my7n7pphJasZe7DuRaAt3CicuJ1miG9tw6RvJtv
p7tsJxWnG/fowwrAuFDg2NfXVLXXQKtTdqoSSbjL2Nh1gP++lZEylUxqkzKD
FdZk51vWj3Vf9INjqSprjfry+/jkIH53ZCZoajBGTQxEP6OGKWc9DkzKeJX0
GRDtmh6J/ZkKqxYU/cB1lHTkxu3NGJRGi9AG8UaYHRaxQGoBEtHEhd+ctf8s
KuAfiE4gxUfk0p4WW69XI/O70msSg9vEmLD+Z8dYIYhvhk7cFRgFApKhts8O
jN4LLaaZLlJdj76gWdYzF/Ec4bg25hJ+lGa2eE31LD1NtSXy13TpE19GzGzo
URrhIS0bz6LhlTE/D6SQVGefmfv6JU9WnNggk/Gdjpu6s/gt2Ip1ulEW6FwD
+NXRGf7N5lDlOkxk7JiISFEITtxT/bZSEB/4qf3E+ut/ovjbXqyJNXLVHZQN
7PR1KWIwy1GpHcHL1uKI5xe6b/HF5VHD/CF+Au7uh/D0v9Gtz8t4f5NjU/LN
t7uah7WYCtiE2HqeBL6ACuSa9iU+USwHUEbJlSipB+jDqP1gdylg3GTrowTd
Dyzvh5XjmYZ+ltRwCKIvxnYZshVmWzgsxyO+obFMl3zEByLnWBidyGpZV/Bb
0NOpADuRyJzcil4UD8at5SCiMpp7N79CbcA3kwCc1OePXvegalU1rujHiR89
OAjo6khDtGXxp7ghzMPHVDfQzyKncx0r8KNaE0FMafBUXmK+FsWB+GgIlNgW
TemvU7R8Slo9dcqeHp5fCtcvwbX3QA1kZIYz2WosNjne5W+UqB2hnrHWuRrh
W0ov6wd1F+0SWaOy986/n8JXpz+QTPKRiILa9gS+A7cz36rCxAAsVXV7a1M6
ZhdBJSqmgB5gtdY0DNLQP77e1gdfCD4i1rH6NGpc+MeW2XQEsEXia42C7zyy
HAzahRBrfcxTlcBkncMGOoXkWc9BniOFFVKyGEm+d/AP7SNcuG+tj9vJ+AxS
NvdKe+hndJiJWk1jiAHflEzU95iN1hdiI0dKCvKiEI7z+sp3OVprezk52AOI
KWvgeQ55Md8Ed4ko/n++IxsIQPODAsJIfzvcJR5lmF8V28ZOz8CKJ6cfmQHt
ovINw6dhFuGxmmH39V76sAsUktPlkF2X1/G9jdjcCjaUu9q60mB8q8zcFho3
nXyvqIF7kldxvHPbUqjmE33VvqUz0LI3YJw9eTt7phL272ZAz2kEn6IQQaRk
/i1hCapzkOvpAN8axlEO4nKOgrsmIwAdkLB5tfTxSdNQVWa7MxXxe3kOAXAH
R873mbPGrjSZHlzhmqbX/oyaa8DbwHrOz29h+Ld7YIB1qu1ctpMyjcNEGmgi
bzcrtqs4xASX1arM9L3ZPBGV6jpv4ZZ3hJN0MidEYyu3fLQOd5G6qHOLSOSc
QOdbZNtX6Ws5azQGS1kNIM2kwwfb7nJdcbVUvLiokMH04HxkXb8gKNJ+meoo
3OGRk6ulGuvb7k/puQworQ68/xKs32dporc58GByapTq4UTCsj5liplZMc1t
lQ+v7is5bU0YGUup3u4P+vjNPt7iRXKmpQEapqihCjo2KQNe3ZJsr/MobMJC
MHGhYW9ppG9fRXFarGOj9AKT690+dlh6RRo4g2qfpbHr8OyNUuJLFtW/lHIo
9fweY4iqS2jbcIsYA3eIGUy1hEnXEqkgK6m55byVvPbKA/13uUyymVbh2jF7
VIm7s9mgrbcoTpuSqTMKUVhmnBkKfpHiykA6AxZNbRj5bONskZt40Wocu5T+
yblRKau3SGk0dNhQePPT7RMMRbEVodXqwYJUjqh1qU/LgEgbX3M+cK8k4pFH
zOYrR8fsBGPA78D/ffMJa56iRNYaChb2REXTsPEqpTHvF08cIUbT5I8SG6a5
JNRYMSmGkubJAsTOMHkdUUB+U7pBZnS5EYadE0fxShYMdxeR4Xe/qooN/cJO
RMsiiPk+vAfkAB5Lk0ewJJD7NP61xlitAkNWcTGm5U4/xzm1WqKXSYbWhSDB
st8fKTqNTFpVlNIprW5zvX7ZsCo3I6ExQvxMV40sWpbCi80wCfm5HXbe2h0Y
xa2RPXdmMNSsG9gcvyWToeRhgJNVa1nIvZjqyzmwzSfQ2gQDW95Zr0n6Tglg
PYP+sGdJWGbmh+yHkwHlWL5IAmkk2MhSYaBn1sETweF5moKb106ixJCimEQV
Sny4dT4AuwjTZGv/8JBedsAWq8Q1fPTiWiiUfPJVvvnbSdn/Po1U7gHuvCV+
QX/zXFZJnYOVzXUrwzaPLzVKCsHF7B3P9WRBH7na1H0AgMJQpFyi9vScJUJO
onkApI1r1UoZxLRqPGzdFwac+Xe2oTqbmN1VxYS6lZkVU3qO4BI2WF40B8eC
xqoq/0XkWcHsUB7CIMgHvFJi6QZvZfrcaCRyvd8shVC3nWYc+KyyUPJ3f2Tg
o7vNNzC5sW4LIZgtV1MM42YS2ANsdgb6xLwsHj1sTUUz5hkkuphmiti1v0mi
P5ffmqredYontZkAJDqiC49b0aAM6A7MBBYqzY17xUsU/GC9C8XVbvoS4wFf
mm4Z8WAVQEAHHLPwJooL1TUzKf719Wt9xX/2FS9S3TfC+yCIU7wlzkLxKZF0
DqW21HMpzRQ4g/lXLXNYKY1zoUKb6a7pRFA/Aq0sCLwobkZABMJUSs8YTTce
cyW9EAKcul3Xew73EOekzk1YRELl1jiIN35JThTGqbGrsFmRJwWgG+eayMdj
T7gkIh7Wrtzfc8J3YM0g916F5Jjs40fMkj/za8l8y/c0kbhvJu8WpdHo/Kx8
g3FP1qsz+X35NmOReqvYFn/TPFFZSMswXhnLjIMeegyy544v29UEWD+a65OB
vdSypXjnWI2jw/qoe8W00Bm/ClGawI7nc86RD1W+G+Zl/WieB0u9ERp8Kfer
vYcpdzB8KrK5GN6c1i3h3FN9TIFIWjoZgmjjDlkBmZB99gPxp9GcETpfTiqP
pqhtHt5bKbdXykull2LRF5gamS9YaXb+CSYkvftOp3TaD8T4cmDQsw8XzQXY
csXGvGB915ZRdpQgXH1w1Be0JekPlITBQy659x8D4LeZQ8f2/l3YvhxvfY4D
RAeb8VbPy4SNUVAer3nFMuOs0af4wEBKFEaW8Iyih77f2PgHZA3Ek9LNzIMI
p7kUvo0nSo5Wgn6vJ2JUQUZ7a4b2unkbrjkk1QzoxqvhyWXg8YceAdYUY5NO
eTmNblirKcIKu/FLzzzgYKrH0B3BjiXK1JcYvBuzNXOzUkAO9KU55YUk6Gdq
IWAeDL2FlnBPLPV5alzfw/WcXhpzl/H0XnL32Q9chUDn7+b1SeTNwusElJB8
I+bf4BEPwdoB9nzj+C7UmwS5sKEqw/F58kmj9VDclnX1pnSAKfFlnowEWbWj
+Nyc80sOHMMm3mw30EgJcc1I02zv1oiygxNnNO4LQsXJXNZXERyTGEd2p0Fw
Ln+WswBuUgunIiN78Z0kjsVhylayoWLdDVBE1oIfweAaCdQ9ZccPWdSOs8Bi
qtzo/3yy1zoKbpuUgol7MU8E2wx/M8znLCaYF/8jZNpbjAbeVqgzHDIQJ3nu
GTWfYzskItDEvtJMYbdcZXm+6VDA8w8VpB40aFGiS8AWE+hZHOHMTAuvImIh
WW/AfCyFeOrM/TDdyRjnf3zL6UpbsI5k4l64Gu2XXZX4fseCkUt52oejMsIg
t7ghxszmO4f3qeteyBGvhl67r7OMGch94hpHldLZvCh2T3/dX3iqXDQkCcI3
yfnHTPikWJDNArGnC0sVf+UcRjeoYsN8Q5j3TKIZVVaKTrIyYQ5izO9wPzRo
ShwOM7wBhjQ5X400qTtrIjkhE9MltJPZFz8+xyruKT85E6KBpvbSJamduMUS
uTawdjVdNzIpA8Rg03XRkUjF5sZV2o/GO5qOrKS6keeFsjUd5R/xeWib7mEL
Rvp/x5dmzHLzZp/cmvT1YRIW65oAgk/8GqeF0Q/Hu24TY8UtAXK5lByvwLFS
zrZt/i1u2d1ryuOIuq0sXaQM1vvpJhTjWRIHJHcvVOgrSTNfmjI2osdV7enc
dajjEUSmtCUktVqxJoJvn/A94iD5hYE+IxNU3ImPmWwaUOiGRQydT+YPgsZC
hQ6563EVglj53kydh4dfy+reNIOZsyAlQPJQGujs5Afa69gHZLvunGQ8zBP6
p6bEv2m7CXX9Fd4nzM4XeGmpNYOiNClta0foaFlJCM/dfy2vREl8F485vjMW
AIvfq1m5aI8PaBUMvBws8XuXCjrkpQD3anaYX4NpzY2HmPhCdcSqeYmME8k8
6GB3oH47J/9xF560+LeLmRblDntGdLpaV4nApyM7lT1ObHc8IN73rE099qse
9PBzS9d/18SRViF8lU+jYuBbgsKGAVdwhJA3pWoDcigXhfqf9m5nmOnTYbwZ
ci52cHGyLLRpaEvWICRXHoLprwUm9OOaZ3OZu2XFmbq0z1eK64xpnKzcDkYW
syTbyvjCuE94qEW/kbLHHXeR7fwV4u0UsuAQ8F/VKddZv1GkaxCKLHSartmd
YxmdG+qGJ94dpshw3SlHAbNPWS/YiBfCcLZVrdzVA5jfCsiq5egsuM7h7mD7
M2Vl2F714uH6CjWIPF+3tvFHRTC1junrd2hEkztWYhXNcc4sZdmzoZUvHFpA
tHMA1LUwWEI7h3I1S44pm1PfyV37n8fQt5sjAHkaOq+fxyEJ6+CPZnnjI4Dm
GvY3dvHhawqurC+YgotNb6Tw3nGGm23AMvf2gQV8DB8Y7CKGoOj0B1ce8gGA
FRg0zue3GX1z/TlzbfXPLCxFalM6q53TbuLRKfW5VWYLs+0E9V5i78zsWAQa
8QjIP/uTj5CkxFz/+aRvpGS9/NG+2qNAwkDDFjWP0ALDeRNQdsQTCNPN7dup
ySsniqnf+CaZLbQxoXFsyZXA+z5doz/202JltALl7wdO1NqWGnZyUnSnsiu+
ime2Ch0Q/eTJlP/apaVAdLKomZLcNVq9roqvYxNq0Q83zrou9x1nydNk8alK
z/SivjpiJZx1FQP+ohMCBhxaqqafciM56hurvXUkEqYPzhLEdCZCGdAibSP4
cFLeFg4JlsXKkDY2NqSuSspQfgjlYXDmeS/fBQiwTHI5ieApDWpw05HSoJGv
5Zme6uFKoq5PBDahAQ1/+wXEpGhdbdSm8zqlTy1u9+BJ97cd0xiOudzl4Cz/
zqaRxyHAE0NSDntQGh3W1hI9bt9CdD9RPVxRBoMMHr2AqGSypOBzybkI8/KP
0UOX1aCIVymELzmRmbm7QLTdDxZIhtsVsdJrbrCAHfy0lEI3VbuECESXSh5y
QM7w0W0WD6oBlUGvsEd5ylSsELOmqkLABPaNoCWdE4UFG2y0imeKc4pcDRfG
KZ5LesrAWULfJfVzI+nOERGJSHysfUB3DWJyc3LdMGRpddSbFDoZehYygy4F
OxAziL3rGQ8tMd4D4rqlCE6cH80ew8piBw3Fziww/X+2NBfYiPq+s4FC3g6+
J4xXZYhkX6K+dxHXzLGoaXAmeZHmA1tIb4syzrSslK2b7RTloJ7eo/AHpnn8
mepihY7kLQ4i2wlFVY68cw3CdJ+hZjn/nX+Vdfc6bXsxfkLbLDyBU+A/7TWz
UrAfSBDLRHTANhXgBSbAEPp3OkAQrvz3n3LQcggl2oqOO5Xufo8qdczW6iYv
haV8kY24862M/y082dHWPr/C3RreF3S0MEjhs1YoPh9DSTAsaUgsHJylQuji
SduF4L9UOs8PgFe7Bg49VaKE2jmxTcZlwBQrnn9VRiu/nM+ZLCO4aNiSrt6j
J2KhFCEznP8/XmCr8qodn9LWmGeN5kMw2/xu2ymcjNtusEEZU9LjLgwgnXdJ
WikM4hsiGWckjynNm5E3A2Cd4c85fJCnxPy5hKuqbiDrNYfdRkqQhEmyHCvu
W2gs38/QwxoEfY4sCHsynkocRbJqIbS1QXUDwEj9VoBlR5Jcggc89cc42iPy
jkVtPGVJUb7YxLe81AgivHWG4RMhR2yzv6NTwogqQjbTO2qiUdrbSt+S6eoh
xVFqJAypjfyYBvK0GjFxKrJDRvm+hbKsvZ9EPbg+1H8Too0w4GYrEqI4qzJ3
OpORRYt9FGYGb4ZKOe8KLgxavmILQY2XTfJ0lhwfq7Vxjm1d5Z7DXZ3sVFAZ
MtE0QKIubVSdyNWgtJCMFMheoHUja1MzyoZT07VIU1RbEmjilGSYNfBAFa4d
sGXgfHu4MCUw/1eLpP4WkTpx7fJRaBxRbcGR4I3fGxmMCuJpUMiLdL8wBdB2
4tHvwFGNry9mEfKh0bkOhdrt2hbXrVsEo3Mso8k1O0xrHaQ0tFMGiYeRt42T
rR5DGAnjwhN8I/j+kRFsKg9I3WaiMayj9gLvUGPOyd41MOf6mFV3eFKT5dL7
jlMqW/uh1rnXidriJvVYTNMKzt+Aynb41caFCREpvwF5vPiOAFpg0IST1gO+
4loUSM6LwWhodBN8FilTkGPpeaGHgtRgN0HxVk1yF2XXo+2eiFM0MVY8IP+3
akwmGemOJ24tdoe0pHov2oKmwz9e6Euj++8z6AgHQRZI1mLvJooOIg/M7XyW
/0ifJ3+p1w8/Zuhrgj0LoTuUljV6ScncWqV37cVCYjTHcf0zsTCs0dGJA4Vw
8lBhfAFdXE7VTqfHikPnegfzpTlf+hvag+iRMgWYLinLlaiZXB5oNg+KeUig
oIPHCoNB4eYYfCAc4ze2xAMv/znAuImt1yvk1pH9nxOXwom5I2jQyq6Eujci
LId5EXWuBgcjgN4PGq4tb1oNkA4B1sXSjr3DU41/hb9JcQNvxa5SNAWArj8m
mMWphFjuO0uA8SZog9D2pFIfBSJC/d8qCMCYuvLE5wu+S7JMwMhBB2t11Hhd
sl3rY8vPd1sSVwqhkD8HE3g7W1c7PhLEtvNfzRHtUx82FaCl7jzrQkphWZyN
ZT5HwpuM0p6Bh2w3GpDPP0SwMXJqzeQYcnWMY+Ak/zs/osBjRxzNlqnUcYTL
GJbF5BYxiDRtx3bo3Ay1ITKbUMtcfTRAethdvXh8ccq3FzwpHOwHQE7gA1kk
CA6LmGZWg/ULuDYnGYMAtmqZUf2Ia8iabeswTmLkyimGQXjBfdrixxlhGeBn
oEKOMI2U2u6mLxNCebVXyRaaEq2LvBVWzDTR8uWy/gQSjFGWUqKOBOGRaSP8
VTX6RkRYkHru0aBsOWrYjHjLJdgsxTYiMh/1hasRQvl6d9zZGRReabzC70K+
34nOqONTa2TnffnkaugugrxRfn8Nxr6FBWjBpqh6aRsUYctD85M7U1pOrKfa
QPXECssNlGtaKA9GiG6K++qaoTdqfPDF4yQogpb953/jzED46ZlwLdyWCryS
/bd8/ozxnccO9EZkMmnmVA2ClI8iNq6qKUepYO4gF3P8xtxQieCCZTnSeA2d
lVOoP/ctuCq4M/u7DKrtp1AKVy0gvj52jki1hLizFcDNPkIvK3CgxPyTYRr/
JjuGrM4yGDs2f5pYhXt7riWvtBCG3uA6Fbbi4TE/XocUakTzbeEoAvj7rvmU
eNYQsgpdkV4O5Unjg0ZuxRHVwwA4DR2PSbqotsekyDPeN3xbWs8ydDVngws5
x5nqjj7GOQ/n0yZxZbUjreZm+yAiHMGGcRQ2AdgDD0RTGWUBTe7SSQ52bLwb
+tJO0sWZdwNPt4mttWgbvzxN0BaFMjvL7iK8KVIfy3rfz90JKGV2/LMV67pZ
6Ivd98X9oybvNz4eGRP+5h0azBuM1vMOtLjzezuaKcCDBmgxlW4Ws0GARSip
YhVWhNtNwYFMIm+qSdqp7KJlS1gcCprXjzY5e/DVmgVnLhWIjjMChykbryqm
xXqXdbUQfy4yQ5vKGMljXtvIXLnebMrLdboVZLwX0GGcI7YIsbDezdFzibvZ
bDJopptCqCew7L3h644TZNSeIAZ3sYkRP+16hs48OJTHing3sfBdC1HYauWE
RxWjpX9tQFbveGRYd3ZxU6RWaKoCtD3/gtvH8A6xJ8ZOf3QKsJirsxzBIOfT
XUCJDwNIDj2tDwzku5WULYy/zqnDVzqP6od3DRAN949iU1hwFDNtW5Ey/xpI
5PiJsg7LunpaJKVhkj8h06YfbnTfKEQPDIqHnzuesCKIKa2cdHoqT9ozztY9
l4yvD6gKmm4nOqNb1OcbvfTYRRi86FiB+EnUHUiCyVH3aP6nHwq/D02JfCyi
bDin6b85ZqWE34igiTvHLQAiy/ePYNaNyQVIxAGL6NOwq51QLeCKdcBkNcrv
Ui62oGzsNsiSuWoFPNu3yrDBy5A1ULOTpbcpxpX8EyFrLTLCGoxfA73l3uz4
48GrakokQEo2/0H2nzLB3zcFIJQ/ScWE1CJ7l42DRCLa0VRE5hcqTiB1Hrr9
sxTId/ZAsckYRdxDC0LXUiI98HBTARnXUquKLS9yH+YqGodgH+40OG7z3hjW
tLM0Bh/tCJHovZK5SuLaw94JiSZd8A0D5H+/u/5kmQlJ1V64hyKUysiyC016
G2s88Lu6LSuzYbwnTH7uguUNk5OdNhPaxMByG7/bQ8E+pqaob/mJTemauNG0
b0U4DKw4py/WDV2R2Tf9ioVV3oyxUNWnlrmYzqiuoQo2VAOhONUhIRF3m8l7
Z2FsZZmeF01tYdbgtNBMdXK0Gv3wUJIaik/dukeATeeZgSbiQe55X5SaQipg
CHDZY/p1qSm/SzoJLO0e5DnRIJ3HNvpYLh6qKzD88jwfYpWALQW7pFMGfo35
bJPh/Xbl9hIt4hI9bzErZ6OCSdIcGpSfMmaHOgEcpjQbDJoCjN4sdxKiRZZL
HC2ThMgqcEqAk8Xw/l9tuJyx/wr3XxiI/D/foviF3yTUT8mVuePFWiL4GBYU
kC8/jP9G4Nc2VscIqX2LJvE/sWx0yIPGXBfg2HW76d77w33gnVhHEN6yrZFw
HO3ZUIp/afLAzqumePoVMLHcfrYIyjRTOMmRF+EqnRUzm58dMetjwvWmwcGE
cZjGdZ8e82GmiBxEn/jEx0DHDPSCi6OVakAvegh9rCrlJqrS1rg/T+xPApGk
4jhwHj67U+VKfDvJhzqnZrphBNlf9bnzuMht86kS3J6VlmGliAbWfBs6aJUf
ytvlLaY0we+uTy+6YVjdKLdsOk95JBDNi62/1VvaUG8NF/Nfr7qw74eWuMqv
A9ZpB+1CUy0r2HrWzJuIdso7+qz6EgJo+2qZ/nWOU9RG1wxIEP/l2DXKdNOy
SOyA03ns5rTUYVcuREOxLV+TNlaTgnjPuseJFsCt/HrAc3/7L7/zell23+gS
mDPObo/tUCt+5D9FOdg8KBWJE4OR3rsQcQyGz5mO7+1JER8CMUDI+yQW19n8
sIh7shMt9rv6d1GciawrS8fmeBiGS12eAWaTUQ7gYUajBz1ZM29TZMYciBBL
G1rsL8da1BisPFbqiF29RTAwBT5ljCBpwMU/H7T6/+WeVEW9pcPJ7EyEoDXo
J5j7RkeBS04MxyO0DY9NsnhVYkC85+ARjFoCGui5espa8qoRewLOhoBqznAW
qxlWXjRRroL0Yy3i0MdMhNhcYC+kqR7lAUkb3ATN9VAguVp7tMtomPGzAwg7
2UFTMzXcBy6VX3RdDiupvJZOboETNkCUv5P32QihqNgLKlp4ZrWZEqFm1HiI
KjyLaSpK5dZ8Zo9sLACOe+swkvoQ3cLc7JOX2gkQcOvVEtoIagiL+XMpEhyC
W4JBXefKHp9gTUd6sBjKJoE40pIKkxuIFNWBye2BQJ52qNvfcSkuSCRjW1vD
rEXYov3qIAc3SOvdhj7ykhjDkBI8PETJgeb/fFDNPN19Ilw9PUcXBD3N1FX9
4VF21nF1ahyRQDtSAOoLQi26kv1+7h/cJ/EcANzIk92pH72Ga6mF2o4dKzbU
Trx8EzfxBPcESL/Fi8abkpiCliMyEMF7JzWinCLT0ZWYMEKLgcgxzlTT6WaV
y6ahrDjN3xTdg3G39NXzLOHnL3Gqm3AYMapNkoYEf1PIHri0ZSCLQDHH4wzz
l1zyBUN43aMQ5rc5bVGUXLcqK8bZ+yWSeyQjGYVunQihq0Zic1AHWJbZ9rMK
M/dNU8/ltfahNT6PhWjgjaNTpMZSiWDYpGkiNb55M4bSbiMKD/4gDoff0cCU
frZmsDXEOZTvoOdDe7K1SDhA4V3hzBw2wkoROM/IMOBsNiU/k7wyTEeC1yC6
tZeW1X3X8uGwJOmzCKneEv6KNdy93hRhU4KjM/4qrkNy0ey28Xx0KiXnOY7N
v0eEVmE0rpcuaOjQAaB70S4oXb347TJiAzV7erbnKzNK00jiwvp+43TDYl5L
aMvnBbxNgzeHe/GiPjJ2cFrqlpXTKlRNUKXZ6Ec7wahW/G8BpXi7io6V5K0e
JnRnQ0pRtQRDD2MiPa58TXGcSA4W0ufMf777BHakyvyonazdAgT2evJNjBnW
Aw3q2mcUHJsQHznKl+x/m60bflSt/TSYkUqSGtfu9wRS3i7yDQoTEG0mEODA
1+/aqQHSRohqPwuD/81DaOXCAgqlEoaO6Rk2lg7zLBh1Pv/QIEzMgVD5wKR3
sUCo8wEbSqggWYSsHf2v7MiyO2IpwV4zQ8Eal6fOy2ATYAB78AxNczr+qVTE
PTCXaMkFwMniB2k1b+0Lb87/lHM093YzwHE2jM2kBeqWoNWNenPu0MrmLA3F
FFL16y+mXWOCZX5QSULntLKDk41GZZcU5KIOHzFP+3hB8JPmXoapEjNIip83
+eU9Zt+f7q/Y1tqg5+jhuFLIdIkgSfY/iJPevgLE33Wk5caqjh36vBjF6T8p
Pkx20xc+B/szFPW/xtNAXXgDTx43bHxsMAE5ARatB09Cl2jpnOuMGHBNFCmu
sENf3LuwwqbPxFrLDiZPGTJZX03W3yQKk62YiIvV7ZhGJH8UADsSLuP04ZdF
e7+Psyd0SqBV26ZqPMS+fsyeFE1qdxaNm3mLNgEpkboBynBNQNKZ3NpkQnyh
on+lxLNIg5DTnbCbYajUfku4cA80gys/2Narl9/lZgOBEcE05rVOM8wK9X1W
ZQcabZpkXQ3r3j88iSBxdfMFByfT5/rtgWnC1qv3wQQTSXCjYc2CTQmK51he
bzw/u2e4BvOOmqp1Rw6OA7lB0b3y5w9D8ZSmvPMsvEiE6dxmrbGd/0irXLLc
K3qEIrmhRoWc69CFBHo2uyWDqNUFZlfI2q7JFUz6KkgH6Ap0zainApRJskHK
jBkMRF7S0doqpScoKr5sraRo94StUHjkfEDYX7Shod04kAGitcUfKd5rPTWe
yFidKeHXg5KjsIJHRDrAz0ZIqVUlBT8YC8rmJgzwAahpWaO1lorDFZpH73CY
24WX01V68WcIP/hz3MjWABO6GL5DAa1/72pQZE+gJyDVUe2VzQflqjQU+JEp
bcb62kJsxY2BqezYVSpPEKdUJbsF0Vo+gKpjCd6VKPZL+4CCtmigXiH3bOEZ
5BnRsL7scxgVE5jZL3iEXsss8Dl7EH/Dcr6BRR04e5fkgIgO6F7u5xaL9e3W
gh72KGQflPovKeAP16zr6wRtn1LeNz92EHZ0uNn9+kyERQFKSENhTPZ7v0nj
MEmiDy0ilT0fx4SNBIvgGF1KVbGLhHKEMWXbmAAcpeV8BSjGPj8QfBh95weX
v/fC

`pragma protect end_protected
