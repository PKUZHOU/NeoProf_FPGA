`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
PBebM8LxBQ9gd/ZdFB1nO3H+rwtXN1dg+hGNWY/of0nPQzRoPe+BEwlvjnIJMntR
swk96G73UVc5Nm8uGheEyaLsuckF/udgpQiIrnzx6vYu6oDQ+WNEg8khsfPmVHds
LoU9UDKSRKWvloJYqoHnCoKDt5mf4sEZnBGWjq7Kk0o=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 91168), data_block
eaacYlrQKSbXf6DUQsdwHGvGKZNNTKJwMaZtQSGeNSemMKAFI4Y+DBd4F5luDP1l
44i24bPx5pdEwMKxCjm3Us/bc4SJWLauXS0YGrn1LZdkTZgfYII5GPbnJERzknhz
i9umEriTtrzrc0/ECbzBzCRArdaRhNrBmNStfT0/cNjUHdp9BrKnvO5kB1k9phiA
fIiDfAjZUNT7+192ITdc8o/xV7BXzZcUhMruns0lsKzW22kz3C4g5DLXan5j0wdy
K+LyPARxMrXd8ZIMXk/JqPVuJmmC0EzuJ1bLtevP5cSOHjiByAY0s4bCh0W8bjRp
rzRo8KjliSCkAWV5XbFlgGv+1sU1jrBDI6n1vsi5Ntj7Y3gAVagWlnZvMQJSCVer
fFtFQgC19J0SP1mkdBqOm+g0L9PxGQJVLUBZOxQN9VNs+blefNBr57Tg1taYJHI7
TvMDeUWVcoJrzoYtQmS3lLnkYlYl1zB5+L0Bxns9Uq167wNRICO/iFJ1tgtw2Z5K
t+tNNkNz10eUil/9LiIDDGSR3rla+cwbZp61ekJPNLbeOD9KdBAvv4Jg0IBiNft+
XHn/T8Q1lmrTb8Yd8Ygw9kiw1DWHPiSMlWzC7eb7XHKonfi3AiqJ2GNfEQu6sbsi
BDGgpXOV5lwpXpYpO/AEjxhBxWNS6Ux0lxwcA6OH0JpXmRIMljfyroKbJyOCY83P
DqS+bGlSeaQQkFl4DJXWjhECuQJ2ySFPcG7+qNkXL3iWvIWCg6TTg+e2dyJPVB6S
F3zDniMKMgqvKhWJEbpjkN6WiqC9Ygsvnq369Hm5Pdr08Qgt1gGJbctmxn7mWLAl
cKodcTScoMk8uN1B8wxoL6amv2gzVKj+lc5mX7veym57HpYUw1Jnwa1nEQGhb0hv
N6eN7fEBFgVG3IwjQZPKqVfs8iQr8QQG5mskU+ym3V9WcDt/BU3up9wEA5MCKQ0f
TojuRcraUu0k/hZIJV6CiG8o7Tb3XtE/x9H/bF85tTeFLwYCQf8zXbjB523uUkfn
EO887XjPp8Uc39FmRwjLOYaRsoM1GsEXcWaoH/LSh10XKHAnz+1YObw0llqxbp2s
+PG6hygiZhYmL41mBI1lnlrlnh+apIdacp2N97IXP1RzzwIGK4wbSyvL+mAxWyKn
rQ6gkhs4cz+aUf+szrvGDHFbFGhgi4myLcR0tNok1fJOj8mw/6YZhKn7Xok3XROK
JrTNRSf8s19UuTqWKjQHmR0Mrp5idi2aKwgougFLekhiO2sv0j7yBw56CEgexEg4
jQtgj3YmVMjEkz8TfL1eDnYPAbOaH+u8iO+I4CPn2qj2yFSWKtxOVoAd5BEaYefe
BArsSCqxTwSeHvMPgEePcZD46gilwLYXsSi8KauB3I8KmRUWbK6QlU/sY85qN2pa
eOnWs61X5eI4CqWVDWd8pR3xK/ipXJ1QoguRTf/Ri6/XhE9H56RDE2sqcBGv62IG
hLPVZ5YL2eUqoQ/V6MBhE+O4pzJzaEayMjG2/TzRmxEpcLX+7+bGX84ahDkn2Kld
ccOZZmcnMjf47HcdbWsS7ttB7Yo8472nm2iUcea6WH8/h9SsvzhvJcIuOB/sdnoc
vqnOTeZyo2VLV2MsF0h+dY23/Ww0PRxdPYw8Z8HqHfjWjythLNMmYGtJrJm4GKdI
eEhT7Emc0H21gNZGRN904B/4ax4BNGSreHiI7JfN6xHkyQX8BfIFQ0t1gbCdchvg
YOo0iXM7JAYraO1DEvuMU+VGA5cxudPMy4Epf+NglZe/oHPoHDP3lVnUwkcAHOnN
wqixRHJQ2jnaRYOyQHFn/HZl16vcpRsUXdCHPX76mE9Chf4nbQ7aad8x95rUr/n9
60lNxgfRcc+lreA4z87Rmwp6HHwm/kcmbIiONVO3LWWjDyXPONBWD/P5HgW3f6/m
+AmAC/1+hDBs/Cs47LM9pXKJbhvlIcnpZvFZLQMWEK/P0kOvpAwG7E9R0/f6dta9
DiGkZqu9evnW5ppYOzGCmd++lWmNEbTxd2L5cB7n+C+FY9cvfHAT9YWtpfyJQV/j
pVpTgNfcGgYbl8GFy7TM8tGgm2BMgGpscc9xfspBPsaFJG95LG6JEFh4DCMiqXuo
xxGHDfzHFtzjwf/HMC8v79DEl2GWznW4jt1184/NkhfGdjXCEjt0mUmmng03ubeQ
gvT8RItPP6aAmsXls0hAsSm4rFF6AS6YNgaee9L34O1h7zisVIPnohKCR1Mn/7Ke
6vjfApn1rS41JL/+bplTvo+4v+w/2/dxABMA3xQURnMu8RQuTUwRVjGgpU/qU4Pl
Q6DcH4X3GSFJnpKLvhEoJdfmnwjWcVDe3cHGYhmVUoGIeQrXwXzL4sfbv82f66OG
vKauzHun/Ka3uZ/n5F5l+th3U+DVvVF+PHeI4tr0Gn+wAUNWiyavIiPpgapwzxxD
RYqEuerdS1OCCNmb0TObGL4t2q2X1CyIExoebcI6PKIm/mnWOFc3F1ygNald+Hkz
hZU9Grm8mEi/kkcYhnX01bzRGjVP56CaPVQeXEQH03ZfcjhVZYu5QhTk2oOmeLDu
laYk+xkSZxZrnPJ2DrfjI10zOC0rdE7xAKpo/OeFrJE9vNW4IZ9hnf3V2GXowm2k
AMeIAcm2cUz6ppaBm+pxBJ8ejPCvHH5o5RgDre41SkANdXJIhDyNP9/i0seRdwtw
0fV6BqCFjFdgOXK83IT6W8LmUEzild0VaUtvjgnl11KjVuWsSCgKk1oQ756FDR2D
EgLguWwFPwAX0/lvdr5oROQh1bdEP0Pz7o/0z19V6cHWJQD9KVPe8VP60BDxhpK1
ijEO8G1Otf0cHAYy67+eIMwyMs13g2PAF/LY+2sYYtSsE8xLJHtd53zTy9EZoikF
4dHq/iGTuuCd4e4VbwVE6zmwD7Tqo6RE1WO+HU5pWgah0dYEzG6zV8eeoL/AzMUN
V0trDd/nC+oK5wJT3I6cepJUJFnO7oQR3E9f9+thMw3w3Lv2GTEVHHdtmPTfMqfb
/kOaP7nJvu4b55yBHtLUY5CH0AJYtJYaeI6ZKvMijcryUv4lMjeKujz+GVahLNia
2Porh1bnPAK4T00Pb8qGDrKAwMn+vYqhhTxTk3U6wpOM/KRDoWGKgbJy5o/QAGRb
0YHy4NQ20BzosZALNkc4Ik0/HeC61R39V+NkbOmopvNkFcsnJrjfuJTuBdqYjvoy
CDKuJJ3L+u+Aqp2I3bPbA1MVFkINnIKSrvzBFYU/R90MBh8qu2aXTJQjPUSnU9xl
+92dH+EF5WcdHjIJ5UF8Lzs9QLeE0TEooP9efgaaJ2E8noF5go8vKb+dcHYQUQUv
vI/jzZPH44E1bzeldc9trevIS9B/d1pmYcpApYq1mtTqsKriCci4GmGpW7W43hMI
yRP67j/AqA7Yfh7+WvMxQRcJlUD4BYBlY8ekSAKbAXURoh2w+nmsxNjgLYZB0F/9
HR26wfjQHfPvf8eOG6ul3pQXlK3Z0AZtkeFV+eD/A3rQcg6jg31Yw4nq6yJiar6L
7pvpaoFC+NjrBYfo7is9zEs7hnG5uSMnwq/mIe8PArKu1dF5rQukeSXjPa2td9ks
XcD/WsvrJpiL39Xbbagxql02JR6bOT4XFC2dQV40/NROHhw7MZ5jHd3vHDJBl+io
4r/EDWMXz1lPv0ZOtv3sYReC2k+KzDVqlzqswP4yUZFjGViOMiiRY5m2yQstdxKs
+YL9xFid4LIv1A/t+NfkOiUC+RRzaB2YMDASpdC+m0hxidi5kFmzDFUC/GFN8bxk
e9SZCq3hB42I2KbjEidjr3nvB0QtpH82znMnBkYu2gSh4F1hWA+Ffg0ZqmavMlBK
usGpyg1TVmZx7G44/8bdp6hNDt6Y71LggrHothtcLDAAO537jivFdH485dZ/rmR0
BKHBTFb4BQnQJFHsHP0sW//uR3j/A4OysjIEZxbYHbIkZqKdruLF30P9FQqWt0Bz
ufmgs3ihP+VxAE8KsXSdhBfS09gG9vxL4otiwYmRnc8cKrngcIKZFp9pkPqamBTV
4vu7OQ2NVinczoEESR/AjMMZc68MrpLn+D87dBv70JsuD1ElfxoM2QBenCcZ9/hD
86ze2pXcss/wskyu/8b9q5usjZ3hLSFlitkdwqj1yuYSB3rd2DNNunIqhlo3kA1c
yF6QDZDQ7X/oEwC6wfjn0SaDfcYEiaXcnnkFpJmX0vinBBllXAlkGrEbdWN+vuG5
XLjgh4qf6BIadWN0uE3DKvviRbahIolyS7riFR55BV+kQwqz+YvpnrKztGruGjkQ
uY0sz79o918I9Dl1P9lYygMUIJ6Vn0DKWVEOVa5OngJwnEAyyslpCjuJlfWa8Ipo
590hVw0AsKFshoWpvCBRqClLUTh9AMi/cxhb4EPrqRvivIwyL1ZzUiRucY5lY5Vo
8oPLbUCgytp7YRY5broqqwgIlFdIZw6qdKmxUtn1gGE7wSg4IGAryBa7kd7WUmwK
50M7pFl7m11UoFXUHp9AUkzWeqnTUx73/bI2FBpmhrW4BvH0eRHKqRgDh9otdyvT
t/A1HGqFqM2xHWTU1BY9+G7btnOaNnd1mYoby5xxXe2JQoLlbo9dNujF8cGoehCm
H/zLnh3lhKSxYjWqdpX15H2rmcd7QwK+ARPTGXnBdFi+MlHZuLKAndZzOQBnutNK
+/U+qWW8Gc8E64SiJkDc6JmZpqR66QhoYA8qqqU9hz8LBRCz1U2u9hjwCZTU55iB
naj7J6eaMp4ydgPejgR+bviPXVphdeadj1CL361ki6C/Ey7qYMwqaxH705/TTZHE
foaAKxYvVxYfqE2Wa7UGylRZnkPdcpPVtC1AgDbB2qKaduHLqhHYEGEFUhYL4I32
csZK7CAKbg2GrFwnoNinPb6cEj2UvUKM4jBxD1ksHPsIzOwvpJTbWGxx4OYCK1Zc
nqRiuZd7pYSCKA0U3eN0RTdeQE1qjuk0SiZGOyXfCflYtCfNY/2cp/976StNa/YS
fLxrFVDSSraKBBzfKTqisbnVKeKQZOiPGRsILHzeM6Lis+5hk/XyGbfdrmWKTI3v
A+YAtOs2LGmyU6WrfgdhvUcGaKYwpYLRar3o/c22btjbi15HQH54DrxYTsNpSh8a
UKPfCSqrEU8NDfgg0DXW1c7ULvBjNYPx4fJWKhlBwu6vr4YUySVrWDsjHi48eee/
lfqAyRlfWsZgu5X3XY3l3RTd/Bf8ypmB98HI3IOeGabQbsrtO5YcCB6LOy4v8Ojg
8MEN023faFX5ffpi/I8dTEEdn4EqagkOQodjpBBQZFSpzKKu9V8FVMYoXH0tuo8N
4O73+Pn3pZ4UtNB2ymEdecNZF5p/y+bv7WVxUDyiUKVsa4z2ygphsSPths5yDXMJ
t0RcZEn062fX6Qd8+Fq1yCIy1Lhth3ddoB5MM2iHRk3+j4EPqbHMxX6LwwRO+IJO
dMqddeKfU8Z0yy8uMG0GmoKIkHr9zgmWt2Rr30rcUVyGft9rptXJ6XUOwDMH9GZg
ar7Iys+pZ1ckWFWD4qL/HnMIxPU6eZ5NnbLXgAAXVfsblrWbmqVHuqJycEIKrHj6
Jno0icvDDiJKvZa0jKJyZx7trqM1L2A+QoKXMFL6bsRBptS4VJhrERhVM66bAebL
C7fHsa6EcLTcgWyG/sP7rKK+AILz1GApYkZifOPwvSpWBYW/2stDCWlM8NnhsHGK
bG9ghrk+1LCXUMZQ+2zZB1SnTmNNHJ9nZ5B9NP2C302JhPnoRZHEq9M4Lugb+NgP
KAP1roUzOWHP4YV/GFhcm2qArQnRWphQTiZ1exGtawmDNrepsEdL2+YSAGxmC4SH
H2EVcI01FfiOoJEo3UiVZaoHs4xffUa6i0VvpVmtu5QlesRmDHINWUwvs8bRpIQW
40iLUu9QzHaZazipAymCA5EqoUZm365Moa/DvvSITBNTS11AfWkNuUG/WHLpeF8G
3NiWPtvp0Bx2e652RnuMyk3UB8Q5vf7K+vtrk1WWBqSlhP9VD4/74VQ/jyAytvGS
BZz6W0iZCaqpZ/n7kW7PlKv63VxGC45EmQxbAhuR7SXg212EH4A+fWp/iBwuyTxx
zrLJnWXD8+kOMpFEsZG5IdhL0oupFqKS2DtLt70KRDHip1DlkSkdC4SKOv2fAgiW
AzOw9yDVBAordeoWXjsz6hNgzCJTiU2VDvCsa+DoWjiC+mlnO3HKJfJ76r4yGlFF
AP5+40AqctEvZATdbdtuPeQoTzQuNs81RkoJNMMBelmHjT+zz5BQtoXk3Btr2Msq
GuciMOdRHktgAnNAi6ULyJ+aW2o9lxTmIoFHWgo5jqhS1BjJGR3sjYQRuZjRyRZ/
95wC8KvUYHWEwj4pVK7wQ8IrCpyv7+nlQuSKYn1fyAKILu/8nqqMKOb7pkQ4pctd
f5OYtRtHEgsRW+Zq6bieimkezX+1IDU7r3F6p5yH+uoOJlqNr4P9AqRMeR/T7YsX
kG5n23sBIYRiPC2sAALaYyAR+dBCN7AS9qPMjVHHMRydF2bVCfnjVgmsayTI7ZXT
3d2yDtlJn+ZYHYjNJZ+TitMiPM1U0TPMRlcnq5jB9eCcX/mQKcURHKebpYkxC83u
yl83E/GB41xJIBumLTEbts8Pg3JFQSLqFgc3BVDrsiZecFFvDN6qJX5Cui1zMP5s
HCWl+Sv1vPQbAKNxIB92cW/OfUM6g2VhjyuJWyDu8PQoGm6SsWmpoQtIEMKI84am
vqcI10ovOws+DLhh/d2+Gse9EPXSYth3gmcS765o1VrIyNkub+E7Y10mGmqIFzl8
Ts9xGpUCtXRIPIBtnkGo+rUBC8k32C1uhrkGU53w/cH/X7fFHSqrDe+SXlN9Zy6w
XOzsOrPryhBIGVn9/QiOHS9ozhk8A4py/IC46XJQAOqOspq2LLbCRvgxzp2hLA/A
35bsp2qopZKwu65o+Ix5ukn0rLi1zhLBivXV8B+NW67khkpZGiuAyu5DjgBdpLJN
YarCqEecCl/8EMtU0r3x6Dn5oV7w263empfqhfJk5FjbaaN21QhpgU7xD7CtaMZN
OwDGleDdsBaOMvqMmgXLsDvWVCEnu7g1yovtbN3uSIg2BMlG1pYOcORasZRSSFX5
LjANunOY545gY1AMh93HaTf1Bfs+WD/7eHjTp4JWlS8THpkOjuhF30cPZZtuVyOZ
/W8Niuu4ImX23bcFGcq4T15SaEEUpertv1Radr0r0WNRyfbjfAHJJCp4QK7B/96W
0Dd2iG3e0xRxoxDNLCdXvFWIzUJRn/r2QZZpbJ3mcUncaukmyOdcH3GpCSLZuRad
vq7ZLnr7ko6GZJoeNFP0+S96bImEOyEjohXb2w2lnHU7qkKVs9kIsUvHjpLzen7V
xOadfW+6mOAKYMU6gTtfztWmfrf9NNxgCOPSMQg4ZP8FUX7xc8Z0FOqdg3t6bffb
xSVapWSev00FMqTY6GteWQ4OErbYLlzaApYGh8ECz3LQvwUKtX34CpX8XTcLEfln
kl1A6yJD+SGjdZUKlCqgpP/ENQgiVjucZX3bHsAE0gJAyeSr0Ix8X6ZGgwE4QTXR
7ei04itCNh6bJiJMq+Ma7O3k/sssuLuh1I+hm/c03iiOBRVuBQH3KaNV90XqBBjQ
M0V4I6i6DCTyZaII/CC+vUh/NMmcamz4IET3tI5vJdNS8rIf5ivDqXO2SDDdJBBO
9fQX3QGOKAoVC5yUal4JIVzlG0g6pauFcP3fl7pKqo1vya8XFXMEOqzf7TMpEPlt
v2oNEzQZJPEUqp7jaIHhVmjsOD/54fSZlKuwJJKWEpbCXEvQqtxa8toU/Kx2GLXm
Q/jDchM1J36N3lGafbgBAxMjwS5jnWnkXxI1JWLIj6r5fqniSSmSS3wfv3mbF3gg
vyXTA6qCxhRWzc4YENSD3llChryHhSqkN3Zennl5lVRN+m0Z+PU/l7qdWMuNSqKQ
5+3fDudbFL2zFKPjgJ4x3KdYlXr5RIHg0dYeEzXEvB/WuYjuAMFzpvrMKux77hHk
n6I9gT8r9XnkBMF5kcZYgi/p1aqLxrPBZ9D5cyHlLtGre8WFzgU96UVMRQxR9pyZ
2isWY0cnobMSnA7QPuB1euMOAWpnzbutpguZvBVOPgJmF3O6DrpGOEQdWxNBM77s
iyuh7GLHYuJf9QTwibW+Pm5Voiek8R7XGs7QtlCUWzId0GNe32Oqmmjj4X+DdCu2
2hXiZv76dULPU4FtvMv238fvp+thY9pQqkHAZRskCAQcvnw46tqxfrYqKk0ZJL6J
BP3cn4IabSd+EIMJ/ppwBlrJ9sqZ++M3nZRJTXfGIK6ILJHAEDjHV7HqvJvPH7Yu
i/eghxqSdNsDuOz3YnGMOAu1sJs5Rzp1LM5awWXA0HvrmiWxaf8w+EqgrDc7RA5F
djdMEoIeWcbOxWSLJkbKUFttmT1o9BmwG3zEX0G8Dhix1yVUPnkSPqcxwX3B/vfP
mP/ToEuno3i6MAwoGEPK5/Laslz4OwgUN6Jnd1Dm4J+M2QN332wECL18Fmmw2+3I
sq+T9aTVDwtONExUU3sMXcQVj8Tm0+OaQWjvK/UdmZdRzXb71GPz0psTY2EaawXb
8LbwkTYryeJ5SfCZvXpwKXh+A2x2kTy+Z042LLQtYLn3VI9dtGiqf4tFU+jnascD
6evPojJVKN8M0EVfW7xDNfp0P+jPN80DmY0xZw21SlTwewEMyT7udi0/h0nZ4RaT
xwgxrxAA7iBfAq+FDdFFkCorS1v9tQ5pWQRjnqsRIqv5Fpyp4W16xwAMLOCTw4Qy
hcIaKVVqYJjE0m553rr0FxcxYSBwnsaVUq/M5F/BYtruI/ikMQzipY+Fo3wzAxo4
HUrMZ0Y6KtJVNH6ZllsC0MkFr7LLOFnKlLQi7yoc5HYodWv28dFs2lOlzdNd5SPI
T6OT44N9+LoNUID+GGdLoILvZ/dSLwZulHUGjZ+2d+SlSn9Gj5IPsD9d8Q07XRgp
nV4/N49BQntjx4zz4w5f3JabTSUWgWIiEM0Z215BfobvxVeNkleRlXvaWOCLD6Ki
0rArmMWq0pPq/EDgIb4jq/2c6GRumWPHGQfYryyJaHgdU54OTs7BNK3mkkRHS8zw
R2hLKLFNLuMRn0BCvDsGhe3cLazOpKvRaf/Y2DUn4WZFg4DIqg+76+RQgBIjL1v1
0v8Fsj05WsPI6+HM7Y7VtTvr/1Rtj2ERdA+8Cta5MR0QUEiVIks5eogOJZhxa8Jb
gKV5s+kRBYEsCgGgC+cUW63FEmkrev2T7etnk8YFpCx181VgZsfUjxcdjBazaFRw
mLTw7QpAM2OjHXONHJcX/RySv9GEyxmCitg1VsSXlFACck5XwmQYTz3xSI0X/kjg
uuV2FuRde1GyDvkSz+RtNHSCyRmpzavAgTIT+Y9dmrQNcKOA16a+1CmmoNIUHDeT
vu8sAdQvqwwWRRp9Ya2hvFqjv7MJ9AFf7XzQr7kHj61w3JbgGWUUwFXAakNY2gTO
GQvlpyJ6ocKUGrQphqrtG4Xx0QdgvGc9hBz0Lqh0eh8G4carzN9tlOEXw4WSH7EY
uNhGJueawLP8Php2gaxQqK+OoBJFmiZ/C1o1JSfpr/RYK+in3GZcs46Ea3KLFtf6
IOn2EozHSOIWtuJm1iW43oRpX8PpYOTaMRxCux5TRwlOc9pSHxRCVfwOSvNXZa3Z
9LnIv0WR6p7kCYki1HIXQZL/TStUefDU36fmPttrewx2r8jNeS4cjL07SRJGJbq6
M3wc4yzuSdl82BYz/impsOO6jA7bC6CwY8dB1LoRY/ojiTkaqIVfVQ8gKdDUhVHX
INM6zvNMsCcp4iRdpI5K958Phpv/EGZgu4KZfQ98VKtxz0Vew5byN02+sunl+dWm
6pDx2w2rzDIpGsYoJGYJlOfAfwrQ9LlrO2/rGa6bwO/RwWhvhX1z4dTraduMokL+
OVHGHonHTYnvp+oNDH6VacIm/7VaJhgYhiVjejIh1M4kv1+QF3HZXsWUETqdtDV4
h/jC4IuxmNyJXcw8ZsIy4i/GTpJrEZhD7HB7YMHb0NbEip97dVap6tqi+q3cwNtU
dZ5VR6WSdGCz1M4URHdD9EXeMGR7ndfFz0CL1FymTWnpokfyR+5qbVeYO9yBO/oR
Y4+/kMh6FBVahYpJS9tOt3Zabkun4zX4RzD3UnMTf2Tnv43h2egqKE9eP/E/K4Xe
8nhGbM+EfgQhTZk4OrZwNxVcDly+J0SxNZrvX7dDEpO8S9oxK4zpl9xIuF9PkjAs
sDl1zbz507gEFBDffBIF322nzKazt74ZfTYZ8AZzQii0xDANH4W+GO+3Q4bpF4+0
gV2R45KBzSx6bPEgqD0Icyqj7KFUwxSJc2Y1fcMmvWKdE9hSfN+NzaZvyo3up3wE
gUUv4xUyizsY96n2Dgq6Vo+VFY98fr08Z3ySNcg6+gFnZsOxQdyHSG/DGxgirsFs
+BIqawqknxqX6VbKF4Joysnk9OD4t5nRamGTDN0cumhS51SHp6br4xuVextKDACe
GN6+sCr61+I/KyyfNVw7Ym1XfXjqCYYnzRvWe7lGOr56faV2Ur6u5pbpOOS/sZIg
aRHukIW9wG9hpMVySMmvhSiZb4EfGISEX2Qe7s7g4zifYsYOWMoFxsB3fGos19eu
Ds6EVy6RFQoqIcNz+XpK3ShN4R5VjHGvOayN2csYehGD3s1pXYxRoZDaOLDJJxlX
tkZyoJsclKMi6gN5rIHyvkukV8Tif1zEJBLTSGTXulR02xYfR4Apw1Z4CelWMJ9Z
ucIIkG6t8a4Mp6HG/7O6Z+3vMyD7zXppvYAwiiNnPZvRQ4ZQQP6oSjqkChhRv9I+
YvYMelZH/LuZ0rM2Lxz56HS/pedhsmsKZRqRag2yQ94ybU5kJcD9xxjNBCdeYfuf
n8Z9eL8D1kVYkjgPXn27MnT3pozmzow9XaeKZn9zOOz4f0xvcQUPzUi6XUBHxx2Q
M+iCJUuTDgOjVkYuGY4vtYQB+RED9ETCzwsSQUvTQ3Edc8gMk2UgOhSxo2Rh6YZn
y56iq4NcT77qkzc8wQmAlpTvh7bSYqRunqWW2gP7yiDlaKT6NrPIDqDyGxgWEhOv
vFu6UtoyDNR0q9EqTd+8TKa7vVHjuknya4dt+3Q3BQOoE0k7hI2OWcsowLWEDJFK
zRxPAoPszmhF41pe9KBRr+YJhWvEYH4rn9LqAzT12UXygM9hEcei+BTdUA3vg6rO
BF3zuQaDi+QDF92DE1o2tFoWW2V7b6NbzzFCAx97LDeK2HQxolOm3yGBAn61Us9H
LQRbhMIjnmyGp6muA5Cb1ldxAuLnfnkyqkoFB6PhuBzMzVPMtah3Ee7TWjp5T4ZF
RvUZONeMKl4/4c9nHq8PwPm4DAPZSgA+5L4/U1wg5jEfFS3YWqVqkYaaRfceygxq
4Yt3VXdpQ15h22r2dNJQA/XwgdPsYycm6i+RIoFUkPRgccOi8MaA5mafdoCQ1nbt
o5UM/0Tu5tu+rLQhVQ8vrs5q3Rspvrb4OGhxsQfTmWgxHVqA8V04vTZ9FYpDfcL4
qXlQvMrNyhtTNPAVMBmvX5JPWzUOZlvIfi/yr+a5OwvkJDCFH6BZPVBWUETsdukP
SVM7d8aWNU2reg52BsMwkN6aE7iyBcmi5IUtl5nmOJs5Wmme7ZMr/wWi4eMq74HF
NZ7MOs6Q5mDJM36SlffA7VHKZmdcPZYawY2fZjpzJN142eGd+gvXXppy5IORD3jS
xj2AeTho+FKagX2B4ZJT4EWyso/33S4oSIOdUTz/4fLuM2cic5szHnf8MBEOUhui
ElVbwGrkM03qgPRWAeeGO7gSsAxfWuqk48I8aqFdzNm+QE9zvkKdlvLBVPF3mw38
wcOUMPpCvdvhq14cuWnKENKOsfleDFVWy2mvZwVYNdYTz+GXy+Um3IiHxZJsEylJ
XIzHXyDwe+uKAjTm93XEtHebYCLjiF2jfBP4zjdGqMLAbeQ7/qFlVuHp/rfUQjWI
Xrlkd2JSjCLGM4GXhB7b/GCNks3IJIUoIjP0Z8nxKPNTH2+KRo5KXRmtkNN3VW1w
aBZUVq48S6k9LIVYQneZhLPL4CVjEYR+mqJ/AtQNw8NR5nOXxsyLirNvFJXV5liX
HCEd986uKE5XlOyUfey7Bc+fcHuc/GCfBJxog2NpLr8ZKzN6vH+5bQn8MFrZWKoP
QUwP7Xpg/d6Pi038g06wgl522dLeIHYNH9M59+rVIsaq28wAahjEUk06SeGnaduA
gputMblRbjCSnl75rRq9yzf1qY1HwHlrG66QOQfnNaXhyW837KuGfScTKzq71SCc
OYsYaiotKc8xP+TwK88n28rvCh5QPyjFHpPzBJ91fBspR49hAwF7iKzcr1DmHtC8
1GS+WW8P/jCtPuwroCFmFDRcYuwHVHzG8pFl58PLClKOPvArXzsSkL9D8y09XpTM
Wf9f8gHLEu4sukqSXw+BNzJ/3cc2w6Mir/5hJeNPe2X0xzKxURBkwnt6H7bykt43
f4ZWlLycqXyyMsduDHO7WQZfmStlMZzAEAVLVvldHlKPKl0m9WNU2G84JZoVlAsL
axOtJZbLJssckIHcaHMEdQrBzkcjf6Nmli7vgYC4bBdemwc8/opTEdhuF9ToXrjr
AVMSh8z/spA79oQAIVe8uRzFyUjurasoaCvPADKLpWW5tuL4FjjPeoxEIsrHRTuA
Zs1aJqLHnA5rVLX1H3hO9xF3TKzKv145QUvFxtzfp+Zubtbw+cE+o9m6hG+9ICbT
1//M7AdtSPgtA/pyS6SCy/v3/2V6URJYaq4fnPD56DFmXv/YCT4EPI88U3wAD/JZ
Pzh2Ajet+UYunzZfkDb0BRifig8hNDLwN40HLA29IvNpRKFE/geq4td5egPptVxX
aR6RSJS4+BcOvqWp3JpeWIsSeQslP2TLS/hMajaFiiypt6wWkNmlWdScY2oXG5oa
68S2ByBm27u8wq5qHF3DXtcV3ZLu8M8C0FKCwscMywEG5xquojm0uzX0CsQz3pSo
TT1Kcibg3D0OmsrOJUcj51nVUH0C1M5Po6f8e5JsR8eS+8wlKuCzoXYyUJPcEl3N
QeqY82Mxr67fQIxEdVpbuXE0UGk/jEm6zD0bEIgPI03Xm6WF9OAe2xwelxlYJiiP
FHB8WBYWvoaJJD8zqKiCN3sUdHGqGGhKIy/MDxkhyFqC7irl9Cre8uRWWwNx4l9y
4VZ12BPEXIDo5KX2tF0ZMPVtM/hyMttFLl4Gq68qj2CHILUn5Jarh+E9i/XXDx9H
kasQbNHnuilK36pdDu2sgSiJ4seDnX4r9RHQ4ESIkgOogz8rwCErq3NEWII5dSqg
2uxzG2LcoPUCMAJZtf/LkOULqeVvpIb4umXVVF9I4mH2LVc6jnj5Jjr9jSvqkxSO
xFbW/JwmYhbN7d2j3uyAZeX1Kk0rB5YIPizMqhMOA0EXhpKEgf0lmi6z8/gtp0TB
sUJJllunRqgkLyKsZSYcUE3wb80YPDe+k+iz4CHmf96g2LGAKpJXfoWxmuWtC7IZ
ZnXTZnGnYW4axrw0/woF+ow8+M5Sp8VNEbofe7MY/pAzF08ElBNE+YPJdvDOLJII
EWUPlUOjTtXXhPbYtN33dHbmjfZ0p6f/B7o8H82d6KKDA32tP/NE3ORTJUzXZmIu
1g+CCxj0mO9JElpHRHZIPsPAvkJuF5DyzzRaZcp3beWlW/gZ/jY/ADAylLe/Mq07
HQPqseKutNhHxru/qNVH5voFOWv1na0FcEyr9/zhjdPqVREO08RRaj9B21bWl52f
soxsI8B1kUAkBTbE2xzH3UFekek/yPU1z34KQCjsE64lFz4WwNKxpi9DqhHdWloN
QbYrvVWLKiboiQ/lLS7ZT/miIEia+Mg1wvD2YM/Lcdrxiqfk1fIf7xvv6DqL3kyr
uIe3z9aN56o9jsUHxAbh9/GHN7Pc1bJtsmn1zM6kvdWrULwtYXZpZD5jpNikgW11
3bHJBSmap3+3EpDaldjePeKMG0VaMN6uj0qs4TtZi8IorjjkvVruE0XdiRI15CQd
/UdTjh+gxWBRm/X6FEK5hxo1qPxD7LI+IYf4V37p/yPTMI4W+b0FSew0HLn75S5p
3NgXXFYgQROdmMAgs/O9c47k5RaesNCCQL5RBmbPq23s4E7wdvoXJcsvQpA/xVTT
E0riyzm+ihtVWhwBPmdiKako7ryKA+4qQpN5JOEmfwPXeqiyCkjkxJHQdRgTBv9x
8Y180j5sXDw8bi60DCujBqhVeCcU95WRE69rDHe0YmPCKk0voVVNVkTEeLp8hSuL
ZgVIm3rSVmSzaHPVdv45/JjFM7k8CY84oYqe0UJgYXsw2sMgtw9M8rKR8Dg4XfTV
xDukSPo4SvPPEK/uW78n/yp9VlF+DLWSp2azDY3RR5RfZI3noL7KCfDokgpP98HW
VIfbNzXRzcBPrsPDXE5Z5ScydjU5dbRzNg4frrt/P+OvAWEqn1F00lNhJdrczbDu
dRs5tqJJI1HMjv5CmUdNEgDalzYXGwh5c95SlBYmt3bDNYQNg9F21QVpwzmvCJRP
QSB+6NlxJUWTr7DG5aG5rg15r4b0XIZApvQASc+CXaHka/5xz1dMyE5DZpYEnt5R
OdAqroqE35917qflelv0STZAbi1HE07V00mOGjRNXMqm9QfMbl4mpp569W7gPFAN
CmvgC/U90gV0ULRTccjM5cYPz2EdApTr0feQ4hlBvNYDLjKBrY5GLGBSfQVAlbNB
Y/EuG006zKw+wZYr2fBOVutajkDQ9wTtXQlLrfPKkO8ywTbwYQDojQm3j1iW319b
ML+Qz3956FdbyFOEDdUUaYAG8PHAVMOXK0uzKglTRKqs1+KQD95hbj0eA159MHnT
UBJiSisZTyLYcOW6QhWafSXXsoMG5UFqcEAl25VuYocIJ1ZikW70ThDdpLdbmkr+
HiM+5d4b3EXeMesMAcvxcAB1zAViTVPwSzpidpx2YYyrP0t5nYAa+wCHj0Aa2Tzi
8+Hfg0lC10/qvA2VpuXeE288ltP/cLil+GbwSz3/lxdgDG2qyc9qzlP8x2j9b0s6
Xy2DX6RQ+YUNnC/dMiGgtd5/Y+U1aAvyziYcd6kyjQuvOFsnZveh9fSTPOX6cqCj
WPtvkMjeXkHSCj0axh+rd4JLBPZ46Q6HGrGZ7n6j2N5huJsUUjs+d33YKt814Or/
r2XBHZlgSGNbuw5UautyAmhMEf5k56uOxqnqggSUmJA/BAtJx71b2oTTXkneV3Ef
doJSzvY0JQFwguqQkgDfZGqrbHqUWoAJYh/sSX2R4fpHaEGSpfoy34rHDileoX28
ZQI4BXtO+cbPkjAPZszB1prh5HzeY02cJnLe8SKHbwUvrX8LQ6SEFFj2/yCeJ+FY
mOro/a+CbCVxUXPKWpJSdka5poJH7LxrryrQw2KiiQ36RubEajCQzbjfLD0WIlWc
53dGsAIV93H/5GxP2mAkgvQWcQ0arMSU535s3HVz7T0WIaJ+YrDkkl5SvbYtzYHa
8qoFodyAWPYEZGSF/TQu//3tiZDDv/yOccHDFvZdzsDJxLktsaRGW8kre/5TRE3T
roz6fOhxKhsUGqUFJoRX3NiGZMYbK7MHWXi6nnKj1MYOmf7PYyr3KyBujK4kxlhF
6LA3dg/gZGnfvCkzc6xXYULOT3+gmM/GrV3UBUTanf47apGX1mTMjARSd8U0Gm5d
0PvGvR4XPl3PY3HbucQlfGcDFnJlbbtiW0lM+PYAuOaUQQgE+acmbFEhPp0KtuEr
LuD3QkaW2d2p3TSRQMPpByB82nkAP4mqPf0xDTWGiGgfWYudwTG8Y61ys47gCl1F
ANmUhXz+lqHkGpto4Wzi/8E/9Pes8EGHYKY1h3PUeV3ZFbuZVfcRbS8fWpHsxdtz
YJgKIvU07K0qZFkagbDrqgB9n/xnHrvEBF7YroLMOjjC2cpkm8B/eEz1ZSKiyN0h
GT/mOOruTJTE4/Kdo0/R54ofSk6bofoo15eckiW9ZtKfZV/j9+tyKL3E75X1cm4s
371KaDumbH1XlcMQb3A52rx6q1ZofMGeywvP5Xa5bITZqYEfB002XD6ldA4hLkmL
MuV3q+yDdtt7qHHg3K+UFzpAaRNTnz9R8o41BwlyPBfrM4vFBeQDrBCpEy3Lt6JW
bB/YVfV5EP3NDaT5WwMckmMWNQIts/PLOiid/5aNKyKvXXKINqUGjVkLujpzdeWT
ZBS9l9YI1L9wr8+Y2n4RGstZN42bPfSWeAHBUXBkp9ctivK8G85J6+Ly8MogjUYh
AaMZDFK47/KGAdpqidKaDICpoe1t49JwDbX54bSOEDXzqeA/UBLHDWxtY2zc4Ln1
0lVCZzfetQPTkTU/2/Cv0sFfyotgHmN4OupiWM2PFYwLAWXYpZ/v1pECO42SVNbf
BrahyK+Z/e7YgyJWX5qT3SubEd9o5eXljheGEwVs6M0KpOYKNt7BANnh6yeqgKHp
2vIx/cfs4VM1siJ6G9Q6ifUVJniTQ9thKA5/dv1iytn8SFJmvK4BCZIjqS8Ic/Zw
/ypDEFqyzPa6xkSlaNpDLKUKZnl92KunkxeXfWe0iUmX2Rj5BGC/nX2tK+n4m/cL
37SAxu3lZ0Wq7OihfY1WAhxl/BLwVFYP0T+iUJRAhsvF195l0GrVQU/2su9GRwbr
GphSDW3XN7QbWkrXCUciQNdh+HuMPMbD2wzjNi5XoDTRCtlEzUk0SxZvntWvGQFV
8eBKnRja0iPj22Okcg3BJRO1vJbcaqes6cLN/A1uzbp4bMq4LV2LZXxuDzB+Soj8
vzR7ZXKJ5Ee3zVj2DLcbSTKc0Sf4nbDnC11qMNslx44OfFcH3Ew86TlX1kPnMk8R
navHTyXwtx6m04sD/U/fKHN+dFsuMQWY74ayow0UwWlKWTuGIZQ8rOPEhgPan0LH
m8D+yvQhLQ30N2m/GNZWa9BzfreakQGAlIH9tNh1rEgPNkYokQFHEsuAHTmbQCOo
FWYW8A1i8Ew1gV5lRrorFvc4xn+Wa3YXpME0kLE5kA3wySiKzgffS/B50rr65lDh
3nAjjA+L+bY+UzDA69NcHiv3dGt7RfwLp0kd2/IPDofo6kRu/W7rga/xMCGuY5OU
Sc+XMVuu4ecxWcMIMOxg1Bt9dqMtXklNjk647skqeZ47pT9A9hE/xFHv0IN24ty+
//3t3F3wJjNi5gE4+hVDRgSAzvY0w/xfH8i0TL9zHclXjmTwUPbZ5xo8Jyz42WGa
VB42cTqOwAa/TyehN0IK0k/8Exs3VrQCqJ05p6BWFNIDBaUFZWgwkdfdBKu4oNqJ
F5OVhthbESPj68qBGJBRcLAYB5gDFe1MCeC5g3PsHY4eylB1h2AJBL5fg/HD13Hx
rBmKcVRFRyzhtw9jYDvt+MKGzxxqxTvGS2WfhNlcFPeidlpRk7PpuKaqDKSzXWBr
TT9uL+PWbQ55XZEHzJAxTC6bpLCDp7o1lqRTk8I23aNvV2RvmePSltFTKms8IbpO
GOMdMIxbG2Tq+IaiiNYzivxPeZSR/2P/5htJvvqKqSZXjnYFHQu91jmJ8PJm6Lb8
3sElEfSYeW07lEmCTdhFdWPdEjfys6iyYFCpt4d+I6lcagqK3ExNz8497BjGbT3N
r7LA3JFa+OGcDaOsOUP2nF1gSA54S13mU8VzmW52/KERsWzfaEqD0jmHTxb1djgG
/69FZyu+Y6cuqcM+U0nPREigOHiyuj2cAitvnIOS08EO5SJ3glOLYXv6d6qpOlsM
WcQw3D6ZFmHpxoE3U6Pv1pe91FadzL+QO5zxXLb8J5U8ZvMpxz5yUZ6imsLK/MNF
ys0WLpvhRELOlC/mqWYA6y2BXnpUChhwCv898fIxODF048/nx5JuclnQQKe99JMN
oPzjvvwKcbaFYL+gpFrUWfAunjdXKLTQqptFEVdRwKIM7X0zXPo7IGe+NnnScCql
1bK4CxbLE4qjh21N5CwDxck/o3FUfd8e3QALiBqcGCK2siLIRFMyIca2tskQmuZc
FdUhJ3I7hRdlM6mcSvs3l/WIhrYoKe+kCk/c+rvE9KY27I1wBC1CK2enSpIr9GwL
4b23IAiNwsLQv2xbEFQtjlvQgph2CZhlMbt5pXJFFKMoAHh0pwvOZOo9INjRQc4G
PcxGLwO9dllx1wsYt7Zdf/hAQrn0AbyGNUfxN7PsR4y1n680RnvpJ3iGnRPYViZa
+HjRv0vroswwnHLKG9IYokyuuQYHJD8sqGtSFvo+IPPxvQ5UMlUH2eUoO3Z5EG2N
f0qPrE8JBMvpcQnYJC1WFDq0THABYu+1OBSnOXOyRU2YG8+gamEPIU+rmW0AT65e
ZlDmtxOcUckxbirysbmLrC+uSvLq4bKAfF2v4R4nxiPDVM3SOypLTa9M0WfyvQe2
1HwNALDWyQJie55czQq60TYjrR0pa1Zf09pO2gSeV4KJOCVQnPa4VJ60ScaKwB7v
PXr1LRQ0wq/Hco87agKcOKyiDYyOPDcqRudgWQPLqytRyAlQnRTxvRRhIYji5JyE
+zhmdWpG3Xy+dMTbg2QtlCSu9yc5Z4iqvLpIki58l/y1MHf2qAm+7/Fne7ZuEku2
esRXs5jLeX/gkdE3u2pg5Aq8wje1KvAECObLD0yUnLXE1vnwOr62CjT9Ih9ZOeGG
gtXbMkv3JF7PtIEu2g2MdQW83cQNJ56cocW72mmnzaB8cp9R7NiBhyao3b/XKQzO
v79ksW/T2j3a13KdO4I6No5qURtfDofCtr6jMOk6dzcaZqE5MVdboTz4VjY5/34g
AGyPvkezDpkHiPe3nk5TsljyR2BZ0Q9gmkQF97Fj9rJqW8+hhgJe6Vh+swo/z7Zi
pa11D99kYS/5P47dEfuqvwF8sOH0eTQgDgVUzY2xyhSWC3nynwoIVaXM7arD+BJX
tfkamdF72Mc3MDigrzs8qcHlJ8N7eFrovCR20HdGoLOK1f84mmT3I5syCBE1G6PA
7i+73S5QfINxAyiwhndtrohMZwW7gCnuoXcKhZhUgu0YVU+J/zl8jCVMWWaciXGy
iVS0sLaocjdXlPWMg4u2ycDr6uG7CrH9WJk2G8rR1L4+oGyjExYtvY2fZYOZZOBC
o9z7AQ3ABzpek7UrhTohgvFyMnUtZDENCZ+jc64O1x2MYwqvyQuZ3EPOrUy6SGms
pIPA7fv8ilDCGdZnJyseQ6I+JrF0hOqJ6eyXduLAGRe7THLqG1FX66kfDPmkAQW+
eAJ7npK1rLLxkPROZKap2CpHSpMH3JubLz3npKSVlrGK8LrH0750kb52K2LGq4Fe
1d016/fbAxCn5LasDsWCYPhrfddJaCpye2Gq/PaSHi6ZriAjqrou9z2VscsYBYjR
hGY2KDXHPGo8eqI9Ohd/49T3wED1aQ1Wzzgb1J68Kx3zLdnkSfZlTtu8CZv9gjLe
x79v8CZLyPMHKuUHqPyc0+vijJA/YEliipZPOP5j7katnX6Ng3cZ+kP1vqZagagV
3Dg8kvV+IvlYnMTXMRUMBeM2OLDJCyoPnbkurdQEKXzZs08UM+a5uDpPNcTwRa5Z
gV56vdjzHXg5qQCSzc3qGFTVp5uAAjF6qvV3q0ozpfesFvjA6ok+3JcB4PylY7T5
gkMoDj22WaCf9+RN5ynxsLoR0Lf4K1PGIq5mYyHHUYtDzuJ6O4hgYInqM8lW24U5
UfxXkAjtwJZymzI0aCXaJj7HoyCaL8MNQSitSFKYr17gKlSOgifmROyutGVIr7cS
8IqtHXTOQQpBPpxkVqun/BR1nZYkGAuQtUWVFpwdCJASOrM3ySr3xZ/fLqR2BbJU
8gToQCpoU8j+sEy9scv4M59X5eZPdsn839sb8qCyH4x0vYnDod2aU6L7iuP1MDW0
6tlWUrW3nhM+DLY2xPOvabVU7amAhY3kzfJi8YLo+sLwtg/yMBNp8j2YC7VcxsXB
boYgfIMwbGNU96zOARTt2ved80BqXSB4k+4W+6lEiCJJPk04Rn/Kta7t7VIGBl8Z
GJBexygXNQP+49xzucaTbVspGPrGvPzd2U9n8XFeIkgwgJ0Ccn6jr1536h48jkpL
8gkX0HDnTTd8217F5/w2a8LruBvNuGm25pd0fQYL0acEVj+cRDlbE01d+CE9gzPs
ilhc+44SHN2aGyULyZJ1778TRdrdzLhTnb5gmNPz7n8NxfVp6BcLjRnrzaFvFFnC
pXnXuOgp+zi+ZliyK6ooLxTZuE6WWMjpXwN9v59BfNLPUphKmbX4+EiaRWmySXrA
Siuz2+H6wt0MwTOu3y19oSUCY8swSYziZpU0HRswluyr5Xuv6jPysRihwRKBh6jm
yCT9FBWLCUkr8e+xRP1rnztdYEh3izH7b0s3U6D2f3AjqNBw40XsPxn9QS8VGeCQ
NfM7mptcJgxs28uctGqjrdTsXNg1XPKeFU0erVlOiFlTWQlJ7R9B3sGS9gs8GRC/
J5wUGSkbIOcfSzPp+5lHXWf1cr/8/mC+WBKooz8CnIfcxM5MQfSprcQIs+Uby0oj
PkAqvLlDnIj/5VDnDHenHcdUj5nsdse0J6OtZfpFL5g73Xv8s+ixx3aE7U6+k9eA
AWfP9DCIy+CZl1oAqqeB9udd+1um8XoSY8Hgv9EAY0qELXN0/Dt1Fx/5MDTJApQF
0PanOP7qHN72DGmvXW+gYgHj8szigRsb64J6nj2wii5dpBMVADjFXOp7Wq/+0adF
Aa66bMbJoldqQVFKddma+b9NGGVebBOVzN0gI7YtFViQIBFm/wSJunqyhPXLxV6S
HknNl+Ny4AET6W00ji9rxEJ8fDtWz92QFcEGUnMlYD6UicdpwTurmk59uYqsa8gj
gvfUEYBnHUSqMW8iw8akTlbYJ7LrCscACkL5saRaXdxyy/eLPFW0x4MhCaZIwJM7
b7VMiNU6f2qBA4bVGqCAsGOedftbm9JGi9WnPl80HwxBI0SMaE72py2TRF8ZwCr9
w1MldA19f3uJu30Tp0Ackx1XOP9gHxpMe4S4nTb1Rbg/Vssu2dl8DcviVzLeT+XG
nN3y9LunpVP0BmqxtJX/aB4CiYaXxc3SQ2IcjjeOiiZmJPS9ppDKjLw9yTkdc8ml
u9zoibsgFzHgHjOV6TxXPpr6RM1uKvsQacmAmoFpj1e8mxdikSUgKvCwCH94wJzH
O8B4wYaCGGt2651JPWDbBEC5zESpivduddsnMnfnII/AM0IFVtrXn3uFeJmdHfKF
L8zdPT8eaVhikFqhdh97zivahgbN1pdDAUoE3GgGaVFIVUcW1Gih5Et98UhsZ+lj
GsSgScYHPFJ17GGQnJjexbGTD3+lE2X55G+D1OdXGChuha8eNXSICZk/yjcZVxAu
qSFt3cvUDQ/M+HXUMe4RBxjWtcEKNUENlOGNKCctUjFibgb1c0robokbHSOgdiai
zvOI9Jeu9uCOyXtONrhDXFZlGrwhm7RJWZtWceY+yRMPYm4CVhcZul/xLjrv+tN/
uz2s0Hwa1MkRpq8ayXv3Vv1UWowJ78q3Ivbiw39mvII7l3EhOYVST0NoWNh0Ynel
nGkJslN9+U7ra2OiLWZX03KjjAz43N7GVcIBdmrAjzBOQh37pXQJkHamDs/qvQe4
j1GTM906Qye8aW8zB8BXdQreMYiqEZWivA+UPuEVHVXhp/XuIG/0QP0q5xFZAHKG
5VhUieHgUI2vOEV76oNcIW3OrmGZV/SY/aCcV+0BXXABxImAgyeOYvDhDPa2IWJK
PeS4kAKVsC/CtxBcaJvJM2uEdRR4/RmoBnvG0Scxg1lBgUuZvjZGAaZYY2wuSRME
lFixF9lLN8fDmoCX4DFxR73l31aDZq+DGNGHFveNqWdVrJjCe1uJC1xdHuBMDFwa
GtBGiWQPfIYLqtRRPIraE/mTeF89m8rRoRDW5R0GTlwJuQ05I0gvltCHLuIx+j82
g+CWx5D/SdWtF4BPTqe6E4znM/M3bw1/HOp5jIoLe3NKMAoWtHMiUDJA8q1IKjXu
l2FH0bc2ebOUHITKWpfmLTbTUfa78puVhp++P8aWu34FR7BkmH2jc5aH6H2z5UNn
0Th+HGZJz5r5C9OK5l9nnhFncZvjkKBJPcHT26w82EKE7/e32Pa4qS48KD7Qg0fF
/mcoipbYXBYXHSUCFhNYWCOiIZkSeBThNTqGRpTUSlDbkqdjz9jo2kRPkl/loaqD
IIFVTYlmZtzpEmUVkIZ1wxcNLUSEM9e9DdAzzOsPRd0KaQ7nvB181xxxyFXHzK3s
5YY1jzBtmO90bTA1J/M+bU6lhdNqZPp7Cmh3u+7UkxzfnvKjtZTg50c52JWkDN6T
K2ES2GnSAKc3fKI3ghmmGXoeTbxrom1xI/G8RCcssvuk4YvMVpj+XS28wumzfqmO
KaUQsTXO9FLg+aEbeaNgx5Nkxu7XG4KQyGj11jPtriLkDLN00GlzSWmFb5pi3x6m
r/u2CkBD86wiHhDVDD5LRZL7gQQMAwKwE9on1SEuFzxbP53qHxxCdc72AtAoGfdw
ti3GM+86ElaA4enTbtI9UHRZWOo/aa70YVgMOH2yyrk2dCMS89rQ+WRDEAyL5T4u
W6VvTXDJEuHYgsNim5GvlD8RvlZHaib36lmnyIPy4VCkJ0CQie8xUSWZexAxlOWE
hpe6cMDmdTvEI5BtaVdaJdpom4aDG1BlIDeVak11mf3sqfwQhtwkr7PgtxVRt7MC
LOQ4m/+EAHiIQ8XTtt0+E4gmq7pC+0pze3Op5Lkldxz+nvMmFh3oi1mkdHT88+P9
nfeLjWqndndecULmTfHLdbOxNIk5+Izsnc5+YhlnVCKEHBm+JCSddOS9HVLGxDTc
yD1GwhMZi7q5asvPI7rYKxrb+7bIIgvu0w+uAXNEt7sjVhSzRbDDNTVbdiL/kaYN
lqs/XLoFen84xM9HJYjGgwdlcMmMUYTe9xAmbwMeaCDjdMdWv9RVnCd/UEHOASzQ
wJ8jjTEh4hKjGDsX2zLKDILIcpEaIqcKbBCcrbT6y15wtB/UuqySGgnkcD0LU66k
4gcvIVsIhm+bb4D0rj5Oj5BdpkjreDKfhRaY9Ftvm+wChh1OEMgVh4cLGPtsmSA8
QPTKyBr8dNVJGm5kgeetozUZyZpIVOHFkO3N+iBBs2fRA7M0qvr7S4AY/KBAK3O5
1Ycz5dixGf2fpaU6SJo+WQePw+mrn6SchnXp5ncd1on/X1rzb5nNuc7e9HFEnTwm
NcsNWCFT2lGyjdO3slrrkLDF1oh4ZhczdVilWltht/FVFoG9cRU9pW0gS4+hEVU1
pdEZeBRFYMYwo9wCtZJFlwMe2meol8cU23Ba/ZTWZeheDGV3YVAdDIrjmv3aMEAL
01JJ1w6JcJQ0cd/Aw0O5DS9h6Mr8OCbiZaBdTulino3LKA3zoB0zvm7UPYznKCMg
QSsYm3DV8D4okQwMbZoqq4EaBkBh9ixIV8ZQFKRR73aIgnfh64X8yernPMJV20R0
eAcUMp/9pM+JFcz85vaODb7t+BS0WDZo9WZb4HPkbyNKgIxpd6ws93SuREKhsZZC
SIbL2aN6TUi2SiUc/ueX9rkTzhIfBA302Zo3q30NvPqwqrYg+PWMyWOKJFkCzPz0
MFz26431PheOInF9iqpuhp5YeGKmEgXFIQfezDM35UNvzChBoZCQgvhfaluxspZF
dm5Ag6bWFnmRBVT19KfkjKY/BfdvOo/2zgkvWIY1CoznkC4jBtYKFmSPQz65LpED
tNhdWdfqw+iYpCRwigJewpPwRd+r+ozzr4Mu4yLgvL45660UoHQjyL+YTJXgKU6G
RfN9m+YN8M0X88Hpedn5Tu9YWBKvohghJ+6M+ZBHWk36JsmzRj7FXQz3PKFSpTUo
eeiQp6u8SmfVq7COmVbSKusXoVrKN78WyrJBIFYraGg6hzJ6XLckH3sli+Fbq2P9
IonAArhgnPMN8jXihqq10M9SfDzgA+Ygx6JJdpxArpFFtl6ZPHLRwudW83rGAgue
fgDKIZh06jKaL9TECXYkr0h9yOw2HbvHkv7MGzLgLlKij9ok+LIq0S05+r/J7VNd
2I7Rw2yrykSKC0/lkuqCgEkAxrk94tmoRojybcHwUcG4ixeuFBvZdf/KarnYmuBt
saxmsWulSo2CZVpEQO8ELRI8CcWfLEC/1hT6cq74QQIEd1IiqdSUQxDirnTiGrIN
v56J4taS0tMy4nffguMh9GEis+G89jt5P5v3xTL3gMnfatATyfGRmBFVVSJmOPMq
WNTGIGTj24usxDLarlmT2F9IS0/YqIRNsRcgm3ia1WyRLHv5VAwXo8g6TpabVL9T
rY2T7SjrRLwEt0h4BAL7YDVmzH8WrlCo+qfyL10YH2a4MTdp270rAQXwMdAWWqaH
LEonscMVnFxhtqXBv4OLwZJXAR/G48vMRLlCuLLiGSopJWZsX2dghLftZxuWadV7
WRI6kDMBZWPt7xAScwnIoB+Cbp9cVgIuNYFes9RO7xBWRtq5iFwEaAW4JkoyKQ+6
tnh2gyB3lfG2sM5yYose7WIYxZOY1insX1dThAqYznWkZKXqlQ1cjk4Av3ynTOW5
O1dgF+FhU12GV2CH5oAzY6ecuLTDM6lSk03C9p+4bdnQuzVyPDGkZclj8ZqLioAf
A8lOx8ixsYHv2BMFcel+P65gcE1CpgRSFEkJH/7A+zXi++gF953Am1OhdvTQu+CR
wlG2v2qXDaAZ4uMx3Sr2YubWXsZreNWCRPicA5d3n3gNoAib2YfgpEZNi8a6fnqY
4qRqJdLNPpD9lzimEFBBkbD7FzfHTqnkZZ3mfpHJO7AKWZUxuzYZVGB4xdYdpWoS
lCFkeHEyCh8ZyhX/EPrKO1SoWLxdMaaVDGwz9/sWwm5tJ+xl3RkKyv+q3fy1/zjC
/lE/jJaBhQDBPG+HhIBPbBBFWF8SlO2k796KAH+1tiVAlk1GclI5U/6cL6wUpUQS
anZMJovOBs3MJIRcRVnRYa9514m5faoDoOcYtLXCU5kSC5dwoFr05xUzZQlgtZJd
EgQ+e5DYfDuGW2F8+cmjXVzT8/Pty02RardMr0qHLtYE6+YfkRU/QSXZ731xc/NY
snck+zE/EKWus0NWnLMAHx+/p3Ex10c6wrlPTizYp0ixAwiGAUYXsSPqAewTha4i
V0+VOqjFxZzt1dIEDNEZHt78MvYvES67wmG/Gp1J0gXRcn5kGdDo6pVyrMESLZzj
F9QypJqGsPjZ6NoJcJABtYPrbHaWhrnkF5vpQVfTtHKsvIED4Pchb/0ia22V53xt
ouRxgUSlao6SAPEPKjUh4iZPt2LXNJmP4845ZiMEn6ecpdULjKiXGzmjqKLceJci
asQkH76M+d5+YVvAQluvny5NonzBAPqkeEZDEoY5xETDKycna3JcRFvXqQqdtiwg
s6/WsxQNPfDrT4grURUww8G62nsKZTLRsl6/wu6X++P87/8V7INlaj9MMjLbwIq6
jBqc/HVX2UOmhx/pI4j6+GuevPZ1Ghy+H8fp7ai3ojPR0JzI212CGwQx7PjLCIMm
K6hSrnsP5r7a55DtYb52rv77FXcGgd8NKgLs6gMLzgpCHmUsAU6uZFz9mB0w3GMd
nJ6NfU6jrZBStPFBHGHhZKRhsn68iIvTpgKtjlCJrByh3/TKFu/p+IVKNRldUhHm
xWHdM3Z3Su/VLcWNjS3ZTNDzOBeEFpfzbDkovKaTcXUF9DyzbkRIPVM20A6YX0Oz
tYlWtHt5X1rklGH1ce56YckvBG5z70DxAXq9NoXfJzzwOLsoeBP4QV6c1bO17WKi
lTih50mR4Tdk2OrZVz9eSP1djavrza3rLWr56I8ndXRPxHPvj5A9iJz77KAD0OGn
b0bV0yzABrZtNKeCwUjPgLQ+waWu9h4XsdGb/1DrMN8/jEJzcTZ+TcCR00z+3Fct
cdRwi8jaRrvvP0foC6PDhAndrgWF4aVBCEY6DZ6E3sYxmXp130fMwtGi/BiSnEjF
CYLzjsW4GFzyQRrGJEgkaAhzM8PIM/8DJdZkofPr1bLs1+DFlHPDmxxXOz3xZtqB
i34LTTJRA2v0hjMLzEnFSu8dXoYC1qOwCq0qjiiRzRnGSEFuzj70TaMIAmsFc9JG
en23NK26iq/gTZfCgONHrVYo6R3e7ZeH7e4hcKbn+2LMy4zryVRqXknaBFvI5xlr
NwALPODhWEdtk22ToWCJe6B+MsBlhVmO3KFY/LOoUUZpeUOc6sTxOk1f/hTErov6
HUAyFrEVzEi3+RpyvZGoCI97c3pzNMRXrP+8vqhxLYRkhwMeM++Hby8MEo+apcpw
4ppiM4KsuFDkgePJuS0i824CxJbuygxX/voRd0Pfr0s4yKmqGjga81oOUmdp6ic7
+at1u7/5xJtviJtUZaiJfrivtrRFqKnAFcSVoUdXq9lsOQoOf5b6OYcVzxSF9aLx
FXpvY8a7ctTL5uT1v5AdXuzWhXTx3v6ltwCc/UJNOBQaMk2GbV3l3UgEcI/amVH6
0mjw9dHTvXu+QI5cPBjZu9EJ25HMWjK6nHbP+KOjZJ8HkriJ5VRVIo6bNxqR64jJ
hXtkkyJDHvWO6zxG6vaLBz5NnviWGkkAuEn9EbciLwpBv/y6brBx/ud4F2SjFmsH
1U/i+Rup8gouIL7rKDitttDEfiZqUIayZVzQXPAD/PlekYSu54m5sSRxM9qXXUeW
FrripVc9LWPs3dK+xtMV2i9jney/tyOxAbE5OFWjz4pWTtpTL7pr0lrUQGEiiF+3
mC5sYu0PznlDUuIh0I8Z9HxsadSD9QQ6puwNfxXpQpfsxbF8VdjY3+eda8EM7jwh
m+rfmOparFUSvsxIDJuAL8l+8ZqvgQ+Sbne8RPQ07b+9pao7Y9q/L5b0yKO0n8aL
0u8Pk4fRpn66bhlA5Spkgnm4i2P3SQlWt9ZbqUqCXYOmNlnv3Jh/O3CnFqI4MiMC
QRcZ0+QM4qKPWBe3r0pJAjKQk8ONk16ZM/vSYLwltb+gl8bcy9mY+xc2iy4Euviy
7RhQ8W2RFzIwjnxgTISKAFQFLq8edeg+r0+W3/bR10HivsOrJmGtaBtsv2B1hZz4
Mk+EyU2h7AuoRwNYQGwDMtaClTJPNvACKEHw+2E40qAbW/bDLQJSYZfsu2RzJcSl
DHKTDyiQneREfFwtO7teRNEK9syGpUAzbf2i1x1grsQfLsJCw7ztO4+l7sLZKRKt
ATGjo+EMiM03aRIqYwEoK8/SFGvNjepnoWr2iC57pMfhZMQzF8FHoKBbB5PF2RQ7
rxa1JImNSDZkMO0BY99ToVu7vM58mfc4acThWQFCmxaNNoMZ8T157S3sbjeL2YXk
z3GRK+LlYq5U9Pte1sSVzXltqfBOWf3rFtFkWtL+NKWIZia3SQ8A3gehqYMdfU3F
U6OCWUN2ICBE81m7E4mntWibK14Yc78s5qFBLweZQs/qbdM6JfOdaRo6oqYviCsR
W22MPEfQmljQn0wM9/tD8Uz0QrsKnqJcZCig5uPYeLlfbmmsd5iIwrbPa9LUT+E1
sGgZkS+81it/x5aSIPQ+KfWaIUJE7WUOqepAgV1cXV/R/lvhxt45PE7OSBJeJZD/
xQehs/+8vEfXw0Rbqpfij/3DUxF0+GuYmWCW7AS9SCgaksST2XXnaVZkR9KJeSaM
wr3VDqnJE1HGgTj5RRE5XSqNNgGu2I5OgNbBk1vLX8MySSurmrIJWyCIGPJWgX4k
kgNulN3vkxzQ6aRcLtaJu05kS7tTXJpBQJrrmV3EBMF3d0Ru3zDRuZC1J309yk33
EEiGf0Y43joEkt5IZ3U4RZeAEbHlcGLd23aDnsmX91dt0FuAHuoTLozwfdFzLey7
ZF60LxzMP18ZuFEsAJtunwmBGr5vPA7ehAOz0Hmnqi7KGBGvgiPNEiwmwPt7y7sI
jXKHWh9A2un0Ki77fuLAdKoo26RFnPpXirfHMnJnhMeWF7o7PWFbltgqezeNJgBY
qalpZqudr4vqK5IcXlVd9DwpeFPaDc6eHX7n0gq27D8a/jHsoQjdna93BTsywULG
NWaPL2gMBOuUYFBYwTH2iiJtdgWB2J7z8b5AX3+VCc8V0sT2BnaHRzS4qLRwUcvg
qexkLOdj8qC7oTQFHCEwzCR77PeS1CUQY9qf8N1jqs+qLF6uTuT9CsDBSAy+vQQm
OBWyHvVM4jmbS7+ODQsDJHG/RPIf5qjM41H5Pu0opeW+QFOPrS63ehMau6F960zz
aAqZmJHBOtuWzk6SHSNwdVq38QUV9yrVoqkn2BBfe4WYIjucIvZEjwzbWNK8gp4T
/JD6jxJ61gR06NDQa+nrdenl91QFi8AqWLY78iE9PVgQQENkRnV971kRnXgX6Lkx
1WO0+LtKux7ROA7sWAPTRRpJN/AINl4oD49v0UT1Ry/9vxIdtCCc3Flyml3jwzeO
5oWJBHJdXjhSvtLIpEnJGWJBOl5wxUMF4vuiUkLHZ4oBM2hiaEwO1TmTxVJQXG+r
+IcD84l3pH6fRBh4noxWRrCurkJxDqxQ3Ie7WIzlpmkHkZvFL2WH2Hwq3Z6tE2sv
NIhNDFhcMf7qnAC85DjHgOneGdBBLYTywRaL3axO1XaqV7odId6d0F8XGAxA996R
rtwoGzV+7XdfDSoM7KIGGcjDnOSmy8GdbfJOPgAd3kuA2IxqofWLk/FaKNtfYmSK
5TN0F5DtWeUqYsXrcPhyjv8qugrHYWYk0eqzV/hJ9cKQVdp/3BpnL/aoO/BdeQJ5
umEZL8OhjM0yJCImfS6Laut3odTJD3YKtsizvbmw98mA0gfM6fx1C3fXkJYjwDYt
LtT9RonYJs8R5B3WwQkumCT4v3zbG9UXkOTIidrOX8017P+4DmYbx925DvXMY6p9
qK0nxIHo1Vhbz7GdJCBvbd/N0F89zdxaFYRztV8qV/iRk2AwMuGDJbpE7cVUjBPA
L1JbthiTywBqN8uAKa9bt5EH48FsHhFhyBb71eA7UKFraPlokQYADs0VXtL6Cwp/
M3hSr1j87zW4OffApquB/EC4DW+4LxHIkDA8zyIdbkzRSpLl5hBaG+C5lRg1GfOC
vaRCTrnOq+b1hXhCxRySyc7kjxh8QHwkqjakiEouwfXM8EdJDcbQi4ETc9Y+/nZj
CGyoeVG/wwnwIFNQ5/7XQCPKRcyhaj9f+7PWNh1P0EKmq0VzDMpQ/qK7mlga1Eta
Ohlh6sZFW8AQBs7xWwIFzg9rRUWu11qVLXfCPeVTO4vHb+ItywvkDStgBqYd+4p4
mI8qFjuxDNRCzKyNRX6jGAUmmV8EBSlA08RyE2qOusaxDaUEt4nc75LP23BZMNR3
9ue18ob+U24C9wxYAv3aVYjCLubAcbNp4FOdcDaU8Pald9h+od4lZirYTKXMFJuH
K5K+94e2UGbaJ96KcVWHZITmSj3snCeu8eEdP33RPWDygy5v5cjMbini+8/mMgDu
FGFFdqhCGRHxocXvUKKrIygVoWvKbEBVI2dm/R2YZowLmjyOpJ0i4+pkWxzyI44T
LEqyYowW9OOHxHhi3pd994iu0kg+6oI1Xp3r87LvZjx/yIFto6m2bf8NocC8TDyE
W5GoL7AnTX16cVgiLWmOOSimDHh4RgK4eQTpFN090k1D4MDnvzCgQIVTzwHhu7N+
9gAjYueHXplbCBL9ghqZ3Ib3+XTmvGLpQehuv/8oZh1qw7G/mfFPQo88oCIxZLvf
0FA/F+7sC8zaVUZ3jdwMBHrZnodj9KM4EHBYm54/fz5CQ5IVSPgMVNqPj2Elur5j
4BvkZZ3kBp1JbZ7p2QA3r1jJ0EkL2gUCBG8MsMLEjc9F1V+n7xtXYbbDXb37dRRW
B88IOk9PeG0ZHdmDuyPg79dNiGNHz78SE5g8A3QW9YiVdYJSMjvYD06vkvZ5SsjL
UI7L6I7/NGZirt7UIKbdB9AtUy0eutLSFymXOB7OB+GuI5rRYHfC9eq8DMQnjqVN
vKs9S82IR8djuoXSW9jecz0FrQJSUtM9+uPwbMdE3/IONDWG0faEVj1KaVf4Tpv3
r1RyarZyTVFc8YDmkz28ClepkSwunzvRW4jYWuZ/Fvf+fxKEqL8a2nmFXumfVAOw
MCuvW3Fewer1FmAiWFpMHQhXBJVgln0oCmefm5UhywPGXY/gnSK1LDMe0gDuot4W
eF007oaTBh1rP9CnZYZTsVEkLAUkKbjE8J4cgHHZmp8p86W80FATqReke3okI+w0
gufLNCDDvEgU1+5Yi72jhA0/nFpc6r8u+cGmk8c5OUJJanfifPHYpVA7HBYBuGwH
sUG+g9U1K1smKxa4itzQlehvN+audNOcyfE262daORg4niaj9JG3oKnXEjLSeMh8
De5eilR9rTngQlTud+d/C2+0PnVTRAxucye7Q8a5g1asmbmcvvr2q6FANh/Sn9+s
EVZo/CS2mgjewAsMls95NWQEyjXM6WfiKDTGKKxk2qXqbvMlfz+YHTP+ZIptbD7D
Jo/TcX1oPborzoqTgV8NIRCYbmT7nOCf6VXNGJbR6UkU3f1UbVwPAXItyeHKgWYl
al2Qar5rVQLt3D5gvcQPwsLJ10GRpoX2Gw2pTDoLfhFH2uOvXA8s+/muAe4JLhxo
gznXtZZ+k098MlGCMvCf1dRj3Vv66EKHe2vUZLrIz2oSAMPe3hU5G9ylHj6fKjBR
B9idEadvuFxpM7di1dEGbCT5ydKWZIf49TNkPMesU3Uwsx5ARYeir6vXcgymYa6Q
QIHt8q5cVRs1xGyhHRV2ixuJ4vXtpeCDXiwXkjgeBe0x0Dss9/ARpQG8WHQ2Vmn8
sutXrKk7mkq34kKRUkqRbhT1PDYmJ423ZjCmoDIUY27aM0U1+TputUqVWHCTauqN
h3ngKgvbyoO4IPOVyP1DymJp+H7OwDtyy9j5eBPR6jfMZPVwlS8XmEqZiS00HI9g
kSSdFBDzzEp6fKOpYz4EDvK/5RnviGmdz0Mbzvyy+aopGXHxZwymluA/aGNhjlyy
fmB0kap15NsOoyZwVzt7GW0QTP1D0AYk3pTUyju3nsJ1qP+q1LFgbdgmFkp2NKXE
rNDrT46hT75nFwNAI8Pv697myze5eOjNtgVXEK6r+ePtqlTULgRlSm736A1N1Yt0
7WlNjDIrexoXxboqcVQakOHUaO5yYGfD3ENkgqkrUGtsb0OmckUv6UXwhZYbXDtV
tIS4yzAh5p2Ep0BiBVzUaHl1K+u3L901PqGGdk4NGO9F5fjGkimqi4oh8ZnsgWTR
mqsS4EdI8kuYue/JHfdgXyabyhI4iY7gAdxPoVuhDj7yfmyaFx5uV7RE7TQV04W5
DCv4UPfTLRuhNQuXqqe7cbdJv1rbvmDkBBi288jN48L0aw1isXOujxdX0V5P9T+9
32IEAef4D0xLdhU5IOb4RLcjrQSYKgBWivcJluk7IpIoByN45/cQQxpr0YLOpNKR
gAswKee5CgCf2ajVZkeoMIcwtlGT3RMhjtWDpsbw5Vs1EtZ0jJZH1O/Cgc6cwVE8
jzuTO0PrzBBOKxKVpy0GFITiT39Qb0RzqkqqPjoOIDok3HHpMWejyIgjqVptoQG0
1tRflPaANB+JXwRYofSbL3rl/SOuvm6Ey/JhbJgMh4Y4apdlaylQm+RvWZbB3TiD
8uO+ylWq+0qJMlQDbSd/it6Az6PpCBMmWn/k6sxboEOdl1oKId18M4Hy8eoMl1+q
bII/C8yJ6wsDMq1JK7cbNrfJ/Jrj/NF5/+k4gE/iYqsFbPhK+JayKriH+9nodsgD
dQjC81NNNq1ExG3qQPW3ZDxcHzsB5BrtKYPUVhMJ9FLkvVnNECL2h2Dq/rCkSeXH
Xvnt/FNoyj02nXUg84rWb2wSDAf6RL96M4fpFr5YUdbYH+ZAW0f3qZcv0EMbYX/3
La/CYqobGV+iFSCc2Fvcc27qG1TtiU77/eWOFxXgPFl+k2C2PVt6w0SpjPzngTQC
bpwVo9sYCunRKBc6dA88q6/AYjOdFy0cRLyKqoVc6zdoCFxnPuhJ8t3PzcZYSL35
+QnObsQr4VAk7XTMzZj8F6ydBQLyjDByD7NQ7DfiuIR4nklv3oGi1MQD12GFEKA8
/KTcYHW0X9/LdrUnmQeKS+tFndWfu7Ngn7JM11ShV4svIMYJsisO5MDmQLpKoPK9
tj6TSawMMM8gzXZMKZAYMkMdZkFZNBNZjiH01oUKsr9PucqBLcxC+oqCLIlLNFgx
Q6YLg9BA5tUXwMPS2kEA8mywNx6qIDCQzAF7NniXIKzlZSD80RKJU+/v8e9BsiGJ
FGSqe9E1qGYtDMRU9TQjYVM7XwZyR7Zp/OWDSIPIGuWVW8qmNlWUeERlSAXMmwt/
468TCLi4iGiYHHtd8bg99Q7sureByQ4xCZbTHEojwvnSz0f4szB4REAWWt6cOYfF
gdWX3IvjyEFawmEj1REpv1WJHJMB2EF/GgsdWmkMG3hWM3Yh/dBGu43o8SRXMBqV
8mpxGplZRju7uf/ofxC8PM1/qV2W4EdBMXqM2uyMmdA49bxqhN6PGBBQNdFgOTnQ
PBOUwiwVtt9FDUnwBQ+ECJGiegDTBa1Ea2LZ7qNHqiE62qvbeQdkr895Nu07liSz
/9VFMj+XVpoAUdwGbnRjLimLP6Vi6YlVGQmJtoKu/7srQmjyS1wzGXgaj8Nnjwv2
mghbzFZiZZvGbPRrNjiLvfIoR3dZM32I1MUkLqG+eePqec3/8H/Zz+43xI6q+OG7
HKqLgTlkIUZfUbHGNSw/RIzfarqYB+yJ+7Us7HpZL+qHZ4OkVoyP4qTVifJDYHKG
G4umHTInwZylFXfSkwLPmPYGhBJUcMUmYanUesGmQaPffWj4/WaUuUIzCJhL9P45
2z5xurwZQJLL0lNTJ5diaU+VoWYNCXxG+bQD/luOCbWiy52jouato4zEUOwLYHrY
eDhy5+vDyNK4wrRqy87YuXPt84N3+Bt0lg4gU+4JenQuVTr7WguDotKfEhhgzZlY
P+SkewZ/LUnYyd3rfl50HbEo7cj3yLMab+3gIJNkLOXJmpDw+U9NGesdu/LpLtqT
L4BgO7P7yPK4cvRWL3tWtfIxZj9RDH7HGoUW38h5Y5+ek/3ti4feHgC8iDNOn6Zu
y3j6Bj0lHPlPs3eW8CKIJzRJWXkzT3NMoXonUFzPqt5zjAt5gZ8SPwJnRBI9EVcQ
oTIGpPtnv+B8tOR5yF+VyUyB828b/GWr+WBpQzVq6CuF/CXabqaVx44xNXeSczOs
KbEYh8Me26Dh1AelwrBR3c3l2k/ztSo6VRfx9hKa76OjaUHBkKaHa+a5NV2yTEm8
znN2hMJeyre2daOofl9X97Yj30R4zf7s2+dX58R0cqUFhGePRFNGuMbR2roiweZc
IT20QsDmicjRcadgqpRsHUQfintMOKIIi3abarveJubcpnh7ffUd65+ZZ4AhHfQM
cpJMiccfqq/eMc3k6B2UZEZd7O9CSMoX2Ib92TQZV/Xn9J/H82Ee9dF/jDqCDQKE
72hQhZ87w+nsXh58VivYeLVn3uLXnvHkKYoFRie18Os6Q7NIX5kFOQYDYrXVeAIJ
9J0jYERvrz7ycuKTNuAJR1EeGDZ26gij2j1Jt9IF151+7QxUuFBZHf4nt2Ms3q+s
3r/9EDJXE99sBLn/AZ70YuXMmSPHpFRtGm7Oy/nvFLUpjclaa7JrQ8igXsZ2Rcx9
GpxvgvfngixLMF7U1WM0YpFm+xvhK4KM9AKjSBoW2Jsg8KbQ7HLYz0248S4pBBa6
rUGa2SO9WWadMxiTx8w6Oc/jdcY4Vjk7FMEnsjrx9iUtrMIa6c4f4t3iCJK/EOy6
nt7onNtIZhCSTYkoF12wdu7e7VtnEdStlF9PrYcIKrJpzS+9Xzx3iV2nrjp1Reea
jpmIG/SrbkVTZ8itc+oZNNogZk0j+sttOK81buOVUsWSpxd7rH6AFksgG5esFdNf
R26HsBBzP6xI1BOzuY3x13TDTIboelwLS9O4NOpDCVubG2xg5dFC1IjtNS7ZvvRz
6UOwgdGX51zBggaQrr3UArTgSjkilUx37MPNlYM5SjmC2gPo0SW7C5vwuywhNaT0
MZrE/V7nfvILQzS4LZlCugKhJGsxrjP7JYycEIr2Twri5HgpCKhEuboz/olvXyQl
Z7CMFJpdQBDS8BD/l0TYe9kHYLPHf1GOV0z/s46qycFtg6TvgM7rGcFwG0k2YqdP
/Mbx2Eo5woND8g/PHPJE6V3AvRYnEJ6xUAkQ5mj0R1TnXyqNXH8RxpogXgmF6QBZ
wWi4CmXP3aQLUQoT/i5Arj7+kHTDvXOv/D4JDrySlxf0UzdqSzPvfSS5VhtP5bcJ
lnu9xW74AnOaxGEHh+vu5/7S2CNOkV9clH444tvUVrWJrjNHilaO9Mam9rgdStfd
QaOZAdg3JURMR9/RX6y/ifvYDPadq/FGpZJ+gnq5FAjsIcfAy9BoQDRcN5QTMjkJ
n2Nsqaql7G+pzs/zsnQGjG2OrNBGu1aAvFe3DGkzLcKAUkgggbY8e0br7O3R0ybz
AKBkXXD+HiHlkyGU4fodGdQmPWe3rRBuA4/zjlfXEEdrEKdit9AUaRUxXHpxYBBE
kJ9VpbkPPLdEH5Wot7LMbTtz6n6bmMox4vgd5eB8ZbOEG9frzzoPiSljYUd6s3be
Ropu5B0YmDjwwQaC5WbEcB3tFUQtP8Qo4BOVziycdYCeMtMljcAkGfY/Iqou/BZv
mr478EGSGFDwHbL+2nilzgia0B3NK83SI2WLx0nSU+/bPE6CgObPtq9kCpBzgXfu
T3s6PJsF42/LZh2MEd5WLrvXKdyL1snuhEinVnsqYIKVo2Bh5hLzcHn+7Cip9CiD
wWoqUVuBKZ1mY0nkW5YSXX3B/vDO0vq+Okv+VjhWXA/2gQ4t9RLREydH7QBfkE/K
/LctMm6pHNESf8VanvJ4at+LyzN1mkQk5UCeQzTmUqrYMwWx+hYRDll2po4gSttH
HA0dV5BFwBHjeNf5Xr/sHHXwswU17CP/ebJBtaoZL4NkdYitPjbd4wzCpi6xu7JG
vCEeVT6OUvbgxcQwePCmbHRNcgRv+SYxpDv+7H0zAxjIatWUuyzYdCuYZK5/sYDJ
UaagOMLMu56NuOK1tUsYbURGAf9xVykKk54MmbTATWbU8QJUNfX0SozCJxcqMMHI
G5rJVSs39FWxhljJRB92PkfaU/X0myWJrqLEZmYh+klBLs0JmXOqd+ZhuCrxhs6X
ZS7valUoRfXGaQDFJZnVJllQzVvDticLJWxpjC80kntWBkhlIKz+sT9jfQXTG3bd
NE7oLE1uL1uHM/V1y6jB/kVXib2kWSOIwT47+ZSaF6SA+JYFWLl1Z1n1oMFDzZrB
DvPXKkyDOQkFTlVhya1tTACVYRTSVcamivs5/QeMZLlEHGanZZw1chxZzbYQPlw1
wRN/CDmHs9gwVtGysYnXy7/3NtQTEbfvFlhTg5Su5WSwwGg4UTqa/BKrvji6jv8h
NrXTKYGeLckXdKVkk/TNWkWOFcDmdT5MOf0he9wQXv72o9fyKRRBvrpxhfUQu4Ll
1kC92kNAIKRNDubVRqBBZQNG1n4Zc6YBdeWhLsJYxRs1rWYCdMXfVzBzfeRxoDE3
vMzn00sRSP6DB5sQ61baYfD8brukoWONTB056lmVoGKeTjTTlJTG+JUX6YIOzSUF
6vFnLKG/ZpYqg/zyph/2skxOeHlIJvoLoSz8w0Szbaa29E5YXYQFbwBDSLD1jW6C
Iuf4po2XCqLmwqYT7wo/gowfmCt5vRNVkTQaC8NavO2SArMI962P1Yvzwtj+2s8Q
NwkAw5Y7cdcnx9CGARK+MBOkJ5XEj0hE0x6WpY8pUDMW7uduA7AcSl1zezbR1dS2
5pvNmXm9NcShavwnTXJbfVWCKLIsLrzQZjJfjTfVSapJys6i+f17oW/wrtaqtkE/
MrbZMkqSHuU3R2XYG10XyN4z+usryTtSVgHAxz6waCS8OT6Ll5NqgHxHCMeJaUU4
ZBY/0vNeV8rl4FmT5wopLsrBA0rSJrnGZpLzed/DN+0gZCr2tM2iHHJiVN/XTIJC
kXh6NUKxEuWmGtvDus6XVzcFSvciAfREJbtsBB7l+hkodhXcEiWuIfF9a32Ts6d1
AhL9B9ZidVSUeUYBJksIN0Ax3poLwxUald3naOY6KnFpShYeTL7TagvRzdLftXA2
OZWdnvJr4bLKyuscjCdFpJaJ9NDtQFZdwir2YPwdiVVKVirx2aIpjKAeyHAfwAsm
7Axjy4TRSEprC2yuIgpm7Pau7zJHKHimed88UteXkKr0G6S5zIGj43LXkcMEvxmZ
o0UMzKIDze7SJTSFSv4ZdLAJ5rT4EeU6w3b0bFB1M2GxyM6S6faZFbNOyCxH8vZ8
kxxZ/kMM43hKsR46d9Nr9LTT77yN74LBxkd3SMjYkUVx8IujlIZlY0abhKcpzX6L
wXoJjlIqXzWQ2JsWhiIBDXYHE0sOcURRHOVYFeJpyc8Lb6jHl8m3XJqq3opQiE7k
UR777v6kUETJ2mQHthjTlqvj/1s6tISOKdjDLtNIPdP6TmI0X6xigbgKqYT3X0Mj
xllVcMuzSnUFS1vJZ1z9MIx3j7LbPspDcTN/gM4+snDPICQbL6ZmtVy03ibDZsZz
VFFGD/6nzfkBUe5cGNLkZ/gpFa5W6mLvoHTyO9euZFOuppbE7jUZLZz1JGs4aQrr
y4B2SUAb4L6gIJHpk9Lv9fokSbvnfm9q+QbXpAe4R1D/tWmCWmdmEGzrypJ/Eqei
naKMCknAAW/wYY80RBSlh9ocj77JWieyZDQIGcgByWgjSAqVomhtJrvzmAf0ce/U
omXGgh5vQwBbWEMeCavrKcZ7v3pCoHdDvsIVpALY4F7qnNpzbDQ5GEssHOfqO/bv
I09IOYmjm8wbPgUJsb9ZV8MgKxa/WAJA9L3fs/gyW3iJEQArJacQoVYl6BT9iybH
13ZVMMj4gcxYgsVFLzFgmF+ZREO5Vkulu9prEHX45njwmlVSCTcv1vjo0fDh1twS
r+ZR5yrZgxJwDB2dzZdnFYlgyUtbDkXRTUrN5cA/RiYzVflcbIWJDVT8VHau2kfu
vEIN8Fr1GJnS7JifO82cgAhST9jC26uE9gFPSs6v1x+B0CiAtxWyqXU1w7MiTvhT
HUE6fh4sTvDdfgIMeV2waWCmSP/H0VpKKbY4Wt4pAUgN0SG2JYW65D/NXop7Xere
MmgSi/mXADsUwwHZ2AT2jwoH4eJIAMm0yIgjQXVglKi2euZ4wcBELFptuWMvsZ10
EQeuxoCswNa9vgpMigP0zCeWx2FxD+pj5gbG1KSu7N204BeVsVcMcln2W54lrIXQ
bfyDUyQltzsmnXLjf4alWGEo4DFDvQY000lbzU8WzAq9kqDQC9uioazBVoQrQA+3
5+GzsEVGhXk/BnOJh6KDNJZ+m9J0Qnkksb37jgNv5iDlKk8qmWIJpdcqNWA4ISPM
SnBJAra+cG70yPMJGXagW3YgahP8LoyZgvyzRzTEb6mkpjKmO61/1JmRegkIaHWi
pUaSe0YlnWFkbfVD0EN/7xCLmumKDhJQrKuFgP8T9RxrxNbdxub3lcWQ0sGwUx8Z
2Mvu9BHW/aohrmuhGsJPSwHGtwTsNXeINYpZHidi18OnPqtEe2Obzxh/TmMCpdxP
1ON28TULr2WyVj2XChYdjILxkXCZM5BaIZu5u9skUpvPwbvlxNJKCzovdfaMX2Sy
MAmxupqe2P7fz4wPGVC4dr8zDA0JC3hUpd2B3C5sGuXsF9rPrrcCOer87Igz19+P
9cIlt0mR2TRZ7e4m1C2eyhJCO/PhhVM5YOSlfrs+06bFyTOwfZmI+5hSkNyznvku
hUGqMHVCZpTaUIzn01E+yf/vC9W1KtVWVLtJC3J57M1QOnZGW9pjIVJDxjSUnrme
rn9gpWcht8n6zjlIB7jsX4xfQWcv9RrGvFkWXHSiW7pz5xxJnxP7X/DIoQbhHksC
Vy1+6CSOq7Kg7/cayMkPK+dRObo99FLk10WrKlrds3NQ7OzPSph/8U9rz7tVzzBS
wiPMTNgFdLFtcv/rkRLW/kyD/W8sFloz2VcMKwz0z43i/J1axHmKi92u7KdCPbJW
cNpdW3VwXYprmqE3b+Gg6UkNQcDkfrzLG0LkXIsqneqm1dfEZldbXIjXlQWBaVKK
RDEgNcQWRqlxeit3B50BS4oO1+3WJRKwkUV/OuDzfCNUpaN2yyzJoRDUr6ajMNvh
VXTwop5Lx6RGcMD8WkZySuij6YbAVs3lRDX5TNX/irEA1Skj+bqzk0RjN1TUXphr
COOJSXpjtKjFCRZD1V6w6Ve2oLEAVS+y+uq5uQ5mCoJyxxOUZ+ubX0YVcVxwD9wp
DNc9PdzIsz1aKdsGnePGm+yGR1PkQRJ3ngA5ZR5WmP2Dwobb0MMIdkcdnRfUWPBQ
K2yuI4sJFwo9x/d/rS18d6QhJ98BvS3V05hbPNG+LZ0m82SYZWm1ba6T0xB4MhRE
2WRYDBlo8Jc6cPIJkFEaNzBfhk1W8skVc7tdjwTVcPXRlDFyiI6H+Wv5D93gTPzx
IMjxMEARAsiRh5DCH81l9v0RcQjpNAfqU7dl7u/y5v0RnAzrQ6QtltZl/VZrEKwZ
edWcnuIck31A6111Q91+ABMVJdFpencl40JvDS7sIxw1aelo/OwLPRgTLEXHqMdn
GIHBCB2GFtgAeN5uwTz7e+5o2vTW7toBqyyUefDfH1YRz98ZDWhNz7zltWIkZs1T
fc5NGYWdzvQWCSeiM+wDpdy+FicxLxLTgf3M+kPI237TZk5Dx+sZAgtRGrqPOCV5
m3WxY0bi5FtQ8cumnhpV8spEnphR9LBZ1Zt1JUCDpokrFbk5L/nJit8AobWkBFQN
WmBr6hpeqHfshsW7FsQ5eRTmgMxqJ9pzmjKnn8InZHQ7VShk8eAR5y5gihlVeijf
xQpdxZX7Wj0AkZhiGS9Q+kHIv46KetSbZ6qb5rmf9kZnLVIYYStEOTLFxuekpjIN
FDU7GA02pzH7fL3JP0GAzJSpOZJB8qledQH4VR18CFs7STK4aJp+0wJjpcVSnHf9
+Kxw/TwGdz4ptd9a/4yaEjkbKVI8Lnvq6WCzgQz2w1b96PgXdRi1IDGRH1eehC79
bMuB/kHU6hAnhilXzVk9AdWI5yx8KO9wvwHMD4FHEOwefPk/LK18sjKjtPwjra+g
GoGNx8AMvZg8FynGPLkHZJ9/alyOrfyNI4D/sTJmDWKwivm4/4V9LBsx+ipMdMtk
6hndaeqGD0P8xdPxUBlD5pdMX4FfX2/DM9Tdzoh3HBj/UGcJcyeqdEg5ZkjfBvv9
7Zna/NwZk1FWdCR06mc4c1aTLtpGKhZyGxiIZw+4IQV56MOb9eNnYc40M0BI/mDY
+ZQnKAJdApn388ABDkPEHX3VR7zDVfsGKmYZX3qy0pH8Ps2+9R7RICmv3/fjwNtI
JmRIhIF5vf6Un1OvoPFn8YL9GRrD13dWzuq0MMjvvc1iXL2JOxgpb04L96h8pQBj
7DTegzWh0MPC2CM0x51UGJNRhfIS+SYSTg7cXAIV5cFe4Ct9bysk7slmP89MAntB
/v+nmtZYphsYJ/l1O1YvPksyLqVMIJRPhtJGWQFuBhPyrMT9uOj2reGLl9ueZJRm
0HdANuKj9RW0uA69gBMfIEddRZw6ORfMTEiuZwwpgIzLC2AKZW7FT5TS5fguEdjl
rpG0mIuf6kLp3aNkPOONuMHEYYGIK7L4LDO5FmatjdWoZaTJgDGDyrMx8DHrFPqC
4dL4PYZ/P6Egw7rtQc9Iqt1fbubUwc3PN7IqFnTnxldjCmxiG96TKDnZ3keQ7Hcn
slG0ttmUJF7n4r0R8GXYsr8nkzJ482eJ6T3vgG/OooGv5CfSgFTPVcgrYcykZ5RQ
EVMHUtZn4TXTw+/zEDKIgJxt3S2G4a7E6UIKCNrTUweEMF81Y6snO+h7Fz5N/j+e
XuCf3QKuMO27blc1mPrlJ58LPf7Ax/Tlo1MfJcMlbmaq22cbXkMXe2DEc2DjlZ75
iI87zipp7aJB0iHwNxiTU1BVSM0TIqOd6DDOYMuV2EYIRArIyPMkli2JX3A7IhoX
Duc/6Q5WNjFRpLqJFhjugYP64XtPkmHpLrk1FYQcZvyl+TdKZmd1L9GUVp8ayHqw
hUdCWqmgFnZi9cHwxRIeO0BJAOVdxoScsGThGRuYbyCZTGcAHY0Ioi5GFgOhuSru
GJC3UdslD2eHcwn7nD07BWy9p1p5r2VlRhkljRA12OyLVIp8tafN8D7jSbiLQ/6w
PuYXAIMJcAF5SHG7f19FKRYrt3XEJcL2sUwIM3OtXyDxSLWBR4yhf+oqGm2V62aB
4akWERo/1KsZoRIW8ri2xN9oGt+UID5X6lId7nM1f4HVsC0Fnsd6dv73OwnQMU1X
p0mIY3wPrjfS7tY3s9f8CHtjJ34opjnwJGLaHgBVuoprDS6erjvNQrx2eJ4xmZDn
vtUs/nKzM1/Xr1eva4DZwV6485YCiSSCoB3GmLlAw85Ma3o52v43B22hWRXP8SDy
P6IQy6kC4od9bdRBd+YZPG1Ftgcap12O4/u4bMMbUlQixJFp4gufdFC+6thZKqKJ
FT6Jg4kBPTUYHv8nZV4Ze6pTMVXMTs1U/G/vfafIOXZlMIJTkn+VGvVUzJZ7cghB
hx4cjc4rsny9tTgf6R6R2+o3Fdk3Fh8/nwt4M1R1DkaTfi+zGlqy5MWiVMQiYHv7
Z0s+Eg6QwMjzws4kkWIHhf1ggs6lfM66VzpbOgznNAaMBgwAZ6RhdnKHuVA+ftxO
QHjB2Io1MMDqNhsHxacDXWXf1Sf9YecXjs9eZKHCYQT9Xy0sh6R6rVpD5g2ZMHVw
vUoOVKQwR6eHHgK9tdhlOkgos4rDU+MBfxiIL6qnzaU7r4/u4aFtLYw/RHWC769v
f/AkzLN0Kbbc/vG6F4Gx7EkXDTP4bX4+Fu5b1NXA4p63WhC5FSiiqeQB24WdxGDK
YtMtokV6ceNMzQQBWq89xlTYi8bzEFMu7I73eW7aora2MMMb7YOEsCaKDEYAmGOr
M0YwfDIm/4LpbYlPAKF+XK5uixycaLYEKcmh/vPlEHHIb7/9X82w35BJdVncNtrV
SGMwopc4g10o+zvyg5ncHuQKbKV2njZD9Q0s5UiKtJccICchG6u/06P8MOVVjOek
IxHen8APudTU062vWL5HbxUkuKzTQYzeOWD0VcircTHKMamVpPyM6sYz7WZrbQBB
sC9UQbfwvAm3ErYCHnyOI+owsqLMhhELJG2dtGAvEf1JCOYWc3O8PLig87jiRbNW
vx8B3lZJPts6kiJRGlZwGc95wOQ07RbnQhJY6kYxdS06mX1Mqp4eaPdSBJw7AEs2
BOQHSLH+1J35n3g6zl+4JsnweueupK0UAHHoQMHxEc7qLLowFp9qaKVap4lMuzhZ
u3nAIhuq9e//c5IglmV62Rnb6u9jvK+ltSZ7be8skmoMYRFE8lHzj5uP0I4uX2Va
Ou1I2XvSf3BtkscMVsoUk1gvndQCIpmWXRM/4hRYjz+NEaZp3/nW31QFSI/Oasfb
T/Bt1G3x7Qdvx8wfiWDZadHNIM72sVeKxF6aqjOYOBadE5JE80R/TOPEh62uNB0W
NC2o/WvpLp/pJuomGlAfV/4jPVvAIhuk+fwdoNnRU55WxqNFCnevjLVxaiSzttxB
M0QGYcdfOaGvuGIzokt7YhFvBdrpbYQolSdp3aXyakRo1U0b8bPcVIFNgKreDvrX
As1Tce7FcMUJin39iGBO+NtjtjqCwdi3AYrVOIC8eiiBVx41PPFygp5dYN8jtAqr
wO/hzNPo6IH05i66DCmR04NEugQdMxHwHpgQFmvopetRQsdFHqDWYM/01vpLDvOC
4Bo02/BZ6/EKXBgo0poWrEqFPMuYpNaVGuGeHDjzV5Hgr8eJSYbOcdHEsG2kG+QH
4Pn25c3ZTl8MRMGBYR1nru/e/OvKJj405FXDDyyPu9KOzRoFc61rkdPpUPsAWaZf
1owy5WCJhBNyKBkfmvCOtVJm2J7QXE3R/tky6qP/bz/aAbhod/gWU0pvRKQcxhdR
K14rWFn90DswFLwfZuD2EN+tab7ze2BQNQKczM+OFDbf905NseJUMczbHxDJ7z4n
1tU9KIpSyW3UWN1c5HDbRn2VBwBoTpP6LJfkFyJfwjwJ8nI89L41tw1YTDx+clVI
ziy2cwAWWmHTzlPu6C+mkblKv/Rkc4RNqkyXAxXONQbggMmr7FV0cDahTj70GIQE
Wk4xadF4kHbhc0ZUgKNK2eInMd+qNiJuiWpL8s3O9ccROAN9bJNlz9ginQo0383G
UduiH9GXufKW2dHrBcMeg7dUI8saDtt/FnG0chstg6lAOH7QiCK5IWqL8wbB29Tl
/m2npUf4hkXqy6APSenFNH6cJ3vhKHrVqwqC5GVYJQewf9VAJ5YfSfeXFYaNgRKH
ENzYp1v392KuTj3ugj3WO1lFrvT9uvr79EEtZRThi70GdpUWX//KRzSgV+mc5UQm
UImoeEMikZjvqYdEQn5sMcxuFFs4K6J6s7eu91eWm4QeNmNkxU6m7bymef5Gzcpu
XxeWfGkzNN8G2TZyievpngr0bu/JKXzEHXonP2242KSlgXGTroTy9T/lwTThrWsI
dcUU/PQ7i97AiYLYKJnCTLfezrfs68Ms8+dyYK0H8pgsLw2C3BB64ZdgbOj0szCr
yIRvJ5p+FVLaY4IHwocVMtadpmhAiKI1R8kEUD8/hEWi1R49kn/Ngx2teUc2oneW
FeWMVaMpF05cocZlDm5X6kuggOnAWXuGG8T3nxOI4fXQzu/T7LzuIfFMSUKWKs0f
obiXNE1Mp9aUuYMH+OiB1QVaM2RpgOWixcNwKK/OhBlGLcQf9YbAvOG80WA5dlGu
yjsuX4ERNLqY+qCg6h2FLGktvHazBM5dkMDE+FuOpLyFM3uVH2At9BoWDAnFFtNw
FHdNQ90ltQbjQaPph+BwtWVbGU2RbfN9vhlXxZb6fVVfzncQs6rBHipMy31s8fkm
6LAU2BWaAwT/7aV/yQ1O3QO+jEByWnNHfHWR+Oel5YQF/s2DglORLfnHXZFVnDT1
WwZUyQ133RPEM/rI7sHEz7NK8u7BtpU7ezxsC+gHw+RDhLSD4k6AZ64lkqNeDnmg
71RuPtWY3Ed/vwOUqMD7RQwjjlDgHx/jiaKOUd6DfT7irlFx5NNnwYO4A2RChoIx
LiTE60rOFig9AzZMWtsuDXFImbMG8wPYSl3+8k+CnODKknBK2S6Y7myg7T878G7b
Zca33QZPsILupXDDSTRh/NXHeMUc+wJQozv6oUs/85swnni+F9WLaxX6t/MYQ4ks
2jYJxQSGgnRDrKlOVZXsD5m+mIhNdi4yFUMoF6pm3ATc49aBLMuoT+k5Q3Z0CakW
i9Zx1527brpocUikH64m0pz8BjIpzgQanJLuAWX+tslseTveYn8w6WgvI6ng9G0J
BImDzkD4o9BbDlDTaqPwQvYp4LB9QfsF2oiAFzNGViMKG+lgCJzRyOGTHzjs7eN5
jEX5/Y+5vtz0adXrWSqXnvIXIurShDH5w7fQ50wPOkGb+fdggJ5uhzIYAYEjRsep
85RnO9KrbebqT0+pJ9JdQBfDb5V6teockOK85svJe5BAZ+Xc3EQ0LWhhsWgIqqe+
v73KyAniIPzPD8k3XiiZ6CrbcS1jNYvzLrtgWjAYLf7krHg6ZtsZnktikzTiHwfv
GsDf89xx4QcfcXoSZV8JtqxVTPWI81J1YF9PwLPAIvmPseICk3PK+GnsmHk3gnGI
FRKWXDjo1TD2sWk1PUCAQ1VXdOtOmf79pzAs7D2ThNBJaGToAoD1jteDKwldHjHF
CHpbak9qeDg/K1t30gxNWwTT0K/KxsjjLUbFd0gZDI+25iVwh5cTRZ/hqAy01f+8
rLqiDTWUZsJCBc7xQXnv7lvagxxZhQcKZyLFUGJ5swMj+6xU8Ljc2mWpKq/hEY56
StHjRdh3aryNOJDtjJwzz2AiuEmzePhnWBfuZmhVSJY/WSI+fHrjWzXuAMKRKZIA
mOfptcmS5Y9om1Uu8H2aOkQCo84xdmuSDvl4mttwwDHDxi73hcE5aAC3ZVHB73u5
SD66tehEsWnaKROSAJchSSG3cy/ZaWCL/GZ+jBcZoheDrLtS2jnOmU3bKnbBMAIe
KPPrIpzO4eM/5bZGuO1DVN6IJWQJCO8esa3hxPvxAVCvZINVVWiuhK/yDolcBxvb
WW1dcGiEO3Z2laSQj6TvrQp16lOXIq4lOgjw+sakgt4Vp4W3jXCKSdv5UEYx3cYd
HvFsF0dah1X8xfZ1CQxSgkYD+3SEzoKQCaT0Ac686Fjo+Afh/j4lgPWV7+O1GmwB
dslxIZFx5DPxdumOFb9EJWiPvfYvbS3B+mXxrEmdecU4vsjP8UWdyBPAXl8JUV8Y
Zz1EwsXZwAXatZkV/EhaXDoPtiV7+wumclBqrTp+0DegLpuPjsALC1Pjpiw3796V
jd3CCs7TQ/O8ubIG5pL3kbs9kyfmCfKpRUSUFXUZWPMDn+RnOlLCQthdpJudBqDo
ywS4SPKRwaLhywFG0xoUy2aurZUIDA3nL+Km1hHRIbqFqt/0a4zWRW3dWwsNT5in
slgxWaqIQzXYP+sJ1bUfiaj16MWZ8jb5GqjuswglmurrlgLzONdh/h6mi/ffbItC
4qREnZE+M1a4QazV8RP8epzHYi1NClrzvYJE//W7FschMU3IjNoiK0g/+oc+pAuZ
aQxw0V+FAX62+Fs0VPnyM7sWAGPhVM5eKZYp/3RYoO3dQ0oWnl/eX2EK1jRDLSR6
wPLgPNZiShyqm5yOYA7nvkr7ZFGicr8TZSGbebJ08VOjGO9SGUL2AyX66mvSJSjP
T3uyGf76lKrxIVTH3tNQRGmqOzjQtsBwN/OPYohf+RCa4slzziEscYOnrNcoOvDr
jbWgHcrDFdVqGy93EHNcaQWYDTDq2YbmkGi8/nABotjd9LDN/I2YGIqUDjf9wK2a
ZAr0ExIJX4ydglHi2kvL1VUYbmZu6iMR06vfPVPknsJMs2Wl/QrBW+jikt0x+bHz
qrigth/DtyUciaUJEF8rFhNCHdLnrapa6XTuYuq/HYCav1MCpFyQSVMeWAm0bRjT
g803YG+v0bOJ7otRhC7gM1eiHtfxZVCTPrDsShXFsozFV78sxiNBfZhxIGXYGUAU
ezmyXRO9Y579kapUhIk0DPXJ2mXJDpRUNfkoxemsGB5vuTRulxfCA1/M7Wgw3HW0
y4NyyjkUU2il2CY7xDiHOaMQF4/z35g/RAt5BdTT+Y0LAyDIDHbq7iNyJtj4ut88
cU9pZHrPynERbi4BiHmcMTYxq2xp+4LQIYehBW5ttgtuSPCSCVNap+OhkhiTJcwW
WvGg9m+AZXIQSSRkIKwt6ur0CmCgbR9+bJukr7g2coH6hrTDaMoWz0xAVqxFiBbN
QYq+JleCWXN4iLuc0y+qvIiaL5v3Ky7swLM5Ixoc5hw3LyHjhl3qCe+1x6YMRkR2
wJk1XIbb4W2ZNs98rISJ17iveZO4l1E5Ad+uN08EVRHbw+aAtinuyL943kGDnsNK
S8oCoox8IC5WU9YPJVEFzKKdVAPd3hQrEqcmX2qqmuzgcP9I7W5LOzHsfoK0rUV0
C4z0/uYb06EJNsq9xGmOEwtcjoLdOdeWbkc1k/PCoQRlg3C2Vif8uWx1U1E3jxM/
BuaQjx6a0Y8GYX+LQR8tK+vUQUcdQTRhCNDcbIIu8CGZER3RNVic3zzpbClysN9B
v8Zx2omcEG9lPgpIM4jomFY1kV9eFWnxneLBULdL+EMJ2GLWcSaAKBxUV5ZFpbe1
Rn0kILv/NHDbWR6sV4XMm5EMU8qkegVCaBBvPireCcBve7OfimzjS4AgPYjrCmd/
5kmokdtXXFLlAvtU86fFYqIn3GwidsrPXtKfx7pWJpj9OXK05IuKqpk0nPvToB9Q
rgNrLSrWqCeMsrjn5C220SbkzdZlXTBOWZUrW7RUUgrmXMTOZlZyVW2YLU5fvmzu
lIF2/AIjssPoAxlVFYorNpMWa2uGViCGj35toWRnVEmRjRAy6n6Yj5EISCF1n2Gq
BCXGpn2RnFKb+Z8NpuRKdKvCQ9xZVGkbFjrxVYfc2hMuSAUJ2+xJsHJtYxvzN6RT
gJha4CL2UxL8wBE+I/GAEL77b7OoSErAtx/5sPuvAhtOgtyBOyZNUMkJdbQTmN8Y
Sy3G3CEPnNUsmgBob+qAL6oN8ScsnVQrb7o7uu/XSWlw918QGFCdMGIB5Y2QYCdY
5ZH/4gFzN6EYn9d6SuA8ZYXeRd31iUpM1gK0Y7yR2zZOuurhbbTlhAg7PZk0knTl
75P4P9VCVJlrLfkOwrRTNqQdo09ZHMeYzEnuTHr/lSWpg/VIDce5G2VDNzPUusSY
T8epV+QgEP2bvwIwJF5OD4/bnBtr78aUMsW0ubbG+S60/zK66iASJbQ1k65+8kqh
10e6br1U9M5T58zbBWrLXnPTYkAWK47vcx1RzVocSiHmDhsZEfLse1D4yLb8VUdo
qtfWltRd02gTu7OPtj5tXpIPAXt0l4e/qWCya5d4+85uyowo4ydgoBR/D+ehfzXb
PHL+KwubqsN/eeHROaWzxV8LHa+e9P8zWn9QAK78pDs/TBXyKMcKRd8+tAb+eAAT
gyBzyD292O/QuYDIiZkyAp0fwz6e/dvB7Vf/K09mO4Pyb2wDkqFRZGtYz1Ii2WXk
4e7HZSmB2qX4US/aquLRJBjy4vqXagyWXiB+djrwbYczQtWaFBvqX0g+RrG4nY9C
oq2tbWSIqSVYJTii4ynW3/MXzYumoUYUrd5h5DmRJri8SmLV1zYQp4sHk3CCFpCD
I2GDSYNcJCRHAcug4rFdLbLfKr9ZuYYT8vvD3lWxcoChn2WzJdBfOr+9WApUeWIN
mBb9cX7u75zoowj0qH9bOIbA9gxBlwyHSEkeHJ53j2Qt619PUwmJ/XWnG+ThdJwt
yf4xZ5SfdrIUo0raUMDWAgKPlRLob7yrJMZh/cQoypNhUg9l5S2TzK+UHSv9Gdqi
xn5AQl0LKomHKQm38rxHSB13DIrx9+Ami1LW5koGuy1HOKA48hRj7yr1XHV0GvC9
ccb9MEF7hwX0ZhNNYb0JvGQPsXdbYoPvBqa1D0Rl8KwDE5pj7NCEIkUQ6rCh5fq6
2YWBg1US43IyUU7TrLFpaNQ8av3DmhK2yoZk7tKN+ZFASIR+j05eA+AmiUeeo00O
1yBHdE4MxjinsZJ6ZWYomr/1/0J7oGp1SbhN1gjBlyBgbrmyNMpx5r9vRwefd/Lq
sxOJc7sCyvb4TmOSEmLwLYTJUlYFNoX8cmOb1aqhR8MJNd4eROkpkRxMoB/1vUzG
EMKTG4il7eHslsYak9r4V68C6dr++kl5+RbiYqKtBethYAI7NivRqMckLhqL0vzf
VXdXHOQXbEdDsJQEoSpaD21FL+QvlB1NMkY8ZJe80M2rcgiIOESvKBHjhNPoZ1S9
XA4hwbbg7wPGd2tSf8rkJEQbEtF+m3+BJ9liutAhUckaKPmdmYWyt9q6Lr/j4VQv
TdrbJyzF9CvaZVmsl2Z1az2Z/2+R+zmWdUMijYAWsYrU0zjDQ8Jn4BRXSB/gt5pt
tE4JEJyA/BTvabON8TJI3r9GfWJuUCgucSDgt0zVe6X3oaaqqw3PK5ggxcz3dEfF
fD2QiaORD/YjKzmesEGprHdn60cJvFNJw0oeyYsuYc6im1sXlP3XW6h3OS5hSyBb
Xt+ZPywgozfTE+J/YYxlUVtkes0wKqwnWNmRkV+u+0snfbgSQl3kQOvqbVvJIUPC
3I0oh/ABaSLsQS8nh6Xdv8UswW6E0rPwe3owMa2cDhv0QymKX/1Zczwx3w456VDP
TuyUPpyGpsvqsQsvTsjtgUl1SwjdbWVbCi2hoGgR0uz/2KXsero0ic44RUWs3dpr
7bmJlUCZuGKD1mWELxZPVa6CtnY+OoEKKKgd+x+IS4vZH+oDU8TyIscH1aOcHkzu
TPX92b6MlkuytYkkQk+70U03Tq7Lmo4UdS5Pa6JadIvkiwtLsd74lVvGXmrMUBhs
kua4h92k3N/AbF0XMUG5Ro7pW1pFqzMhg12ayg2Q6NddK+EN/HKT6toNrONeAZec
nCd0ctxRaZQKevzOX0bgVBb0ZbJx3p3L1rDUpVoKByyZKJFx323R/gZb2GO0M3Z/
AerzoCB+IULdxVH0uqd9K+m/VWvocf9BWFv6CZYjM9Nz4vXEE+Cb7TUmbUD0lz0G
oDkxJAfy878zic6sS+cEDjyVtFtlC2LMpjxehGzLWStr/13yg37Adii71SU4baNR
M4js+j0/2HAP+iRjvSwDJdRypL8d8vZhAfW19LWz6QL5JMefEy2U91V9VacPxtJd
e34wb8kwDWBQPGXA2ppdkrZ4ygc1CKD1N5d9q4DTtk8X/xtbcKkbDJ2zPz+WiuEJ
8y0rQBOvW0JQdGufX1haO41ub+sM7yFJARMwhEsZQ9U+zfEryKmQRvCPUu7r6TLc
9ZL/iydYYNHMzVQ6llD7P9DUDjd96f9otpCr+a8rugRYQC2qzIQI/6zcbqCCvA/n
KG5tyB3GmZBawcU8SjIgPboEOyC9aiahP1mySlwPXZSuYGLogPDsiZzULOoCBj3Z
tgY5ekLk/9x/jIIgfEfK0FjO4UVzuVDPX897KIDuiorL4paoJHR76YVd5f+wx7od
8azLn/EtG+KTbUO4LujfTfxkjJrl481ACtj/V6Yqa6NZ44iqFQ1o1lEP9wUNT2IJ
YkMOkI12ouKFgM8c6x6lsoWXn1HStJQPEDL0ftd9lO36+HdIQbSAISFXDMVkoaTt
XlXHjjhihGX9mpPuj1ZkxNFRcebfNhYyLNxrJHqCIy6X543X8WpVayaxDn2YmgEF
GkE+6tMy8Ol7oKr26FkAaQnvO76ePJN7191uEOdML4yKaEjym/aSYnU7ZM4+MVu2
IEgVWfAOlbqOYqwQryF7nWtq9+RYyhfQevMxOKx/N+GKZ2srNGSzY1wrJFUGUi6/
Yg+mDn2u2zlWaEdoGahfm/9Q9TkyWbrQuWxlI0YMep/8o1f+U8LVVfj2BSEQ/eQf
YB+h/pmtEknNPEIh9rLskpBUQ5rW9fNOYEAVC7Owfns7jesmf50FFR76d0sbI2b4
waF21EjCvTAv+dC6g9EXtEdxi/JtKkFfVTr1cfsZJP744K+Tv2LZ/iKkNJe9QSfN
uvi7jwL74mFCNEvniLxG+e1ZFhACCpmnDyb0NvKJS0R1wAh9flYrNRWXX33GnoaB
Er6ktMf4GXcLArOcsfc4+QWgAhwGS3vu5M4bTikfT2mTk93lgbMQR0MyawZMMStD
elmqK3e9IEuu51/2CAxQV+U4u1z7FIsVhyExMBTc8bkfyrgFN6YRxo5QnFjeK2k0
UxUPy0bhVqBSAAFCxFwhd5JXEX+PaFeNHNSysZRH6jPhcU31fbvZEzwAihcfaUjZ
4jH+ej7XV23yS7rHK8vNr0X3Kqlyi9M/qeZL/+9PZ8NXfn0nVjGweFqpD9XL28Lo
lyLVwNg+nGyXrAWltQzMhfzqBfoF9+TUpseo0rB/rFq8AVygBfNZsUkO2QASZs83
wp63fcztSNMOkUdA6QhJdWkyEy6ncEtgt4kMQfKIGtwufxQCKxpISzDSCoWX/i/P
wAYk7nAcTqbXZH/YBPBIvp2vLEVepVG+wOy1RCAFKNWKv3yNYK1y+83BxltmlOzl
EF+l1OLpKx0LcJosfMTYgNTrpCKfv2utf56kxL9YWfwPtpUmDMhzvC/sYm8eI+HG
33c/ak37ihYT7ugvUygaQKZjns+zobLzeDcIjCrhGO7ZbcQRnX9k3OQf6lrk7fDY
a8cenj/f28iYhnrN40VojrHSZzwS+1htLK8FY7GA1I0r7ikZ5F5FmVXzmp3Vkkl2
d0/4hA4BG1nJWO7whmujV/CTrjivXNcHoog2rUxcSfPybhBau3HHcOBJHw52fPyi
DZd6tEOfeOLED0Gm4RiVZlEx7H2CN3F07MD1HXI+Nu4P5M+4K3PIi6leE1x6OIHB
yFQsihdQvCnp0euV4u4WLlN6ezQQx5jkrDMWMsHNih711CInnue+0/1/K6srQpo8
kChlkWn7fARt6QZDie4bVTk98HDeCNq9pkyWIbbUossC80KG/M/MeK1yfxRD4VTC
ewkFVu7r+YebNcUYTlRCZ4PIfwa3kYeFYu8ZxmsoM9ZCs8a991Yl5jRO2rszN/X5
f3tijd9YzDQl32PJ6Vpf0zEBJRWKK1ANs9ymNx8Kl9ic3txH3ebdC3PxaV5t+KZK
nAbbAWV90ytoLBxzJL3yhoYzAUfv0tXvlH4iYb0WB8BWnX5Ys0Deaut1M8GZwJhx
en7qLXzlAS26g8wFD8sHdK1LoILUfeDLTTAqXa5+KJCW53sH2018VAALp+UP6Uo9
gswSLydXnfWLkavWOstJXJPHowwId5F8ZZBBh5cd+PMrxKe16UXqNsfCe69EAjBE
c03c0yBBoj+8JE5Jlnnw+36JDtk7bqX8AeqeLOTlL5jA5ezv52Ngvp90r4bXNZu4
cR8xAnpje7W6qYqTZ9hEuNwHZ6liRTzSJiZ0kYYS9nwI0LmJwEcTl+oyXk/eW3Wo
osPqy5V6SvGt/a4iyef8Ty9XZpJmVYCvmwjH8M0a7HVozuDaqQY/v2uzs7gXBwUk
2OvJYFFQGMlKi7m+0HRKyn0q3PZp8TCVBHYO4yxeifAHxeT5wc8smwpUYaDB7R9o
wcRk+HKrheCFEu0HJcarY0jz2VVGJCMCu/VIQd67Ai81JVau+q9CPFtEQa5/sv4d
Mqn9MZnpbtbssqdxR/ysJZLWfdDojm2+Xmr4yHXyp5ciIcLVil+NoxEc+C4DFXUw
pCb7ah0gYvV/gA2lE0/5kVuTPbSm8rqFNryBuEFCzcYEUGMzr6Ug6szEoQVERLyH
juUS94ei4aBKikt4y7opCsiSN4zQbFCbRCqnXFPEJC4WE8rECWEHJMLTO99qEJgr
Bffyk/bkw46otIiLq69v/VOf1iW9mtoHC62HGFhxloOz0S/Clj8Wz/88jFHBg5G2
6DKNvY/BjJtL6tA8r0UMAB3YfJIbNFQ3wMXdDwc4Mr43PnWYvoLI37t6RZJmUQq6
QyNKxbfA30zzqJJud7VXvOrPxS8v+PZ5rA16uVhwxVneK2+F+O4YmQ1LHizxjxMj
NSKeguFjM2Dds6ngwjB+CwaI3HkzRQjjKuOigVjtpqtxlXKvRUNWQleolOlBuEkc
Sn+1qutyF1WY5OoWHvbLxtr/VN2Bzju+7hjXR5NTbeczL+zOAn3RyUxyXO4hrVG/
iitaV1oF6zoxxXBcFQMxUpYPUvybG1RUgOw58REcOHhv0yO2bABXY8OhpJDEJQ+J
hMK3+70qhd/670T5kk5ugWuh1KlTouGHzzJTXYcyVIbnS8UJhOM/51HwV/zfOcTu
BTYAhl9CAMkF1oynMQhX+5HLLsXMb6l6LLmlMYOWvSM9DoptoqHv4RwLWPH3XKid
eXWfzKUgRGzCg1s5HZFdi155w+xLiXR7KH3r0e2/n3AwjVKGpotGdzBJDNghOkin
5/Q8SYDexKalsYshqOunfvXkd5HNAzXUxWOoYqZ8km7L08YzW20O2ZWv7SQHASnM
9oxA2SxJ7vRS8Qs0rYz6nxTl5NOearDq1ciyvag8bdDSPH79SOF7d68fiThFLZqb
AMrFpThVX9J/ZOUbcZnvITher4LNoFXx2ALTnaq5QEcGK1fBz2FpNzUjWD9QGf5c
UZGjHJV4A+gsBnBzO9MogExKC5dFtlALX2MEcMhBSnFn0s1QI/UsFu83YNNYq6mK
SAzxHMd5sgbgxAJ5tMwol9opegkoIVmasQqbLrijYseUWr6rMu94XF5N/jHx62Aq
qxsvXWgeLlWS4AOe+zAR5EzxsU6NK4Ez9mZSK6jnrXqr1MeO8dgE8sAUZyWfGDuh
l7GRb6dIkxaaCY/nBhniiS7BftjAabJ7DYtl4olBuJJxaNBZtQub9vzwVWjrPPCR
rREY16omSBVXuBkUlDh28oP8vDl05MTdK6dRxCv4qqy0GTWMeqoTlFN3FWeCiFZu
TVMzYdBqNDEtpY+C9HSdps4EOHnHkeNO+Kbap3aO78cq3BQVzUhuTHiv/9cz8kCS
ly+ykJ1FppfE8R2bjufmsOTb/SmIRTYGrkQb3TKLNWSs97O7dXtSYkUilyewRhMP
kdSSQZqGB41JsN6hqFIvrZgO6BngEaOo/QbkqnCcpIlqoIaF7xmJsHdQk/fkN1Qw
kfcl6PjY5RWEANKkgtTXQAa0oNleaYgDNG5pfo0o8A7QR1qBk8Pdn6oUNnMLnqeM
130C0Hk/lGzkV4es7yxsO9GlkjVV0MZCy4Qs1p0/958bzG6hWk8R9IjnsfFq+6kO
ZJuI2mS1MZM5a2xU+Id3/WAu9LC6o+PYu0o2mWanc4+ZRIghW12q17GOFezUJYmi
Qy/cUS/ENPY5myAS3EUCyXz+2atKK8rbX+Jo8N7cSKZYeoqQG8kPPx7X5Sovy5Us
Yw7IwmJIP0Y/uLl2qzDlW9GhDxgOYFi4ASZQORE796gD/k+HXhVqjqOpll8bBnFm
gcMKHxFYXr+Lt6n11XPEsYGBZtbr6L1M+kDv+de3zzFKdrTa5W4jmBGUeDBBFc1R
F+vqOzsgz7UCdEeOVNXuQEpwJLtpS3xWdz/v+uRAmVs+E2nAl/ulpCpH30lsnD5w
DfMV58MAcyHO7Lg1CAe3ka+zf3zrvoAUfAWXgGD70/45+Otkv/76JSlxU/sNVh6Y
8bx8OuhU0X66ska7q5yShbxu4Io7fLN/RnkIbfGmB7ZWOCNIa/aGn4yVJxoq9COc
ODbesDOLzYq6BzcrOUF4+YPwSZxMeDI4RcyvE5mchZk0/zANMWT+sLG6Yorym6Nn
TkFrUNjT+yDfITHaGgSVetLbVx6VSACs8AOYSjpBxKSj+o23fPLwKFCgHcP5Xlag
6K879V8TWtyIX1NEhP8W52LaJ55hvOaZfm1XCaxFd+w14B32jQwTvWvygzSRNwdZ
MjUlkr6USYDsTC7JiqYHySLJsO1h7DC5V+Yhx2fMv80WuDTyqEuOO83mRAe4ZSRS
iYvLKWL2p+jU+6uD5g6rov+qvJi1oX65RSlP2JOGtkxBESvcuyaAqb602insuggv
yce7lpSjUwD7B33Xa3p83l38w0pa+aYEC6KsrKbLRssOobGb81rUaqoCLs77fQGs
XKdSnTTR6BtrxwzrnBVbhtKFM7uzLGHk40fv0/sRNAhOblWI77Uf/iVkmBQkHExm
7o8J9AJvRYOLjg0XrYh0QXcNHrqGQbWxvv+tCKadjkT9vBzOmy0f2ku+pFDSApys
2A2Pr4Y5nJ1QV6s6VJGOJffQUYMjldz4/oBrpGWXTLo5p0Kl+pXFSt6NGDEuimqL
4eI5RKlFohbK+pbyVfOCLeygrNz7ath5Wn28zj8Yez5jfbvxLkxB3CAq+kw6BXDh
6n0Ja8C/LhLs0fkfQImd78L1XTw86Bk+aMithJzSJnFlYT+qSHmRRc2clsJcjX+F
ETz/VOI7LU3YnTU2ouNqDV9klzw1V/pbDDajBHrklKU0BdJg7AfKY0FiqawO0W2F
HnI4Ef+EchbGB6IYpysqEb8HhQAS9lAvuWHuPMB+3KBPhU3udXk+k8fN5ZN5N/2L
7FBCwjfOJYhi9laGSGisudxUrbIehed16TQP6FCBgxZ0veE2V3TUEr9kAmylNDvQ
LIX4UyrlX0I1+T3uMW9jp7ggaGzc+m8bwCQX/612/Sol8uxJPVeVCNte9BJVh3tE
dQDrDuaIiqr1xtLTg59x+j8f4x9XUg3nQrYFpbKa2SUWAp4FzGP3m6Dk4bCM4Ble
zhpd2XaY9WwmZNc2Qe/DvJ7UMGzn5BbW8+7Z2+CC9WYsRO/C/fB/Jyv7U4tyYxql
G1jRTAfKp3GocTR6Vb0fQwQei1T+VWHcq6SDwWuXwmX3PJ/LUkKwkeKF6yuiTaUO
6CbeTCjuC85gDje48yagNv99PprgGQnGcYuDEM+yioWcMRE2aVUzzayH+2OF1Pc2
Luoj20PbDKPoxdZbnBzLEZl7eGKus1wyYdd9nzP8nvP7J/liDGiY+3OZi6oJycDE
YoVveNZOSt22i+ZdwWpP9htVNkUj2FJapjzU5AOj1QWREF9joUrw/puZV9gEq3E/
WSAJT6f/6vrK0f1V9zG1RSV0xKhyfi7I23fWqOPzFAWdY8CIXXqgxMj5ZUzrvpbA
8a2XvSw5kR/cjnzo33ObNdXLFRrWM/2AHhFP+S5GjaTtQc2LmDdeiEshW8Y00jEx
oUh4CICdqVjJI8Sw0GThDTbMKPvWfoK7HHgUbIXQMF9okgtKhY8JLGzo429bPpww
VUKRPjxX8DIuddCgkGPrfZfh+bDpXKGQTgqvg9bxOGEIxZACHFZrW/l5sIg4RCx4
aMZUYIxoKQPmbv1zDvTzmM/Nu+EKxFUCxYp9rSMR4UBPK2igyCkE1xG5ReVbiyzL
jWHPqT+kVI1ZpSSfBYGjPFERwEHXwVnk/1EA/EpQ72NHRnqkmo5DijTNSHAO+FXp
N5iX38y+LJgZO8UqUC8MflNf38R7WxtgW2YmgGg7eJO9J00qyDUIvK4Da/uqaTEG
wHwiRb5xTwtV0Gne69y55kTaaQw7KJFNVfsWF8gwY+GyYIEWskKPe59SlWW5elHx
lK27dArMXAHISkM8KDjr+xNjQpoMVNNPByUQR2Fk64zrb53xfy2DlfkfeQIufGvl
erFuxO8fVPpXrkN4B+4Xcm5ZPInUdPjgptff87+K+JQN+Hax7dnpYDk2EgsgnAIe
jMiGHXkh77Cd53DlkBXGo+yG1SxdOPG27iAmPzDhc3uO1vfsrt9MlU5WLgylWsZr
L/Ldk1ixocGGnj9C0hnu2FWd2gSog6CxhDzxR0eckEfxCVMiE6vHpYfwxF6rL/kD
AR4Z/oYWFfTvozyA7Z5GB4x/2fINhV4791/UzMtk7iX97TPOgVMcDldIJfx+VPgo
V5aLOOsdv54Fnixe9+aP9U/eOklySqz4BRGLuLXxu/t1EhXkRIZ2cM+s72G/3/dS
QtKn18RgUH6OObWoPBfdDiChlLJmuRPrDQmzfJ0uBju1mVs3cSE60TSXO6e0TdjS
rNe8KyN4U+v7bOYjyh/ZaCTAEMsEf2IVW+RWlEz6Y6pxjScuIsChaiHCLr/TKRrt
oluuvu7QXCn7vZzJM1O6MI0jbwW2k1fHoUggoli3SkaclfATGjo5hbdSZAkitmBw
guk7VI7IWVnvZpksTkdth4WbQyruMtvyxo63fJgDfosKJehqRc3e4PZfs6wyIvnm
1/MYsG9+eZa+mEUZq6D7Q4nSJLDzJv0Wgsi/+a0d15MfrF60qx9KZRYUeirxOSF8
2OQgIBs4CUWpjB/STgHjtwZM92As5boLxxBjmt1mpvDMq1ayL5/o/DR8IKvZ8Sku
R/SVFn0WPdxVP5yy9gNocNBKlOZ/LHCeEpXwbZ1bwiGYoK8ubGBaJS/BNvn1u7JG
LkU9vztSP1U1CVUTKOt6osV/lfCrILdwl9/OUZwSjLsxcfxEW34M65/rBlivzdEK
1wQrW9J+5B/Nqg7Dptz5Adjrs/yCWXBDOlPMK5o3mDaJtD8Zeb3Ftr759eex3P4A
15NuSYVTjsmvxhOraXt+2S+YcbwKGa5P9aqgnf2BOiaiLeIqmoMqxn5w7q9T+2uY
wBZu21dU2MzaaELSETgOUtTbtWFrti7XTM7oFWG8msWnrczN5LqCDJuNg+zhac2v
R1tOcEkgkYVSxPtNvB3DeJJPO4CYamnQwRGfy3t+8Sma/pOJdP64BbN6M8m1tlix
+aHt8l6OOHRzVjHQofJosadjIMpa/5kyI+DHiJyKM4NU5A/yy/m7mCJNnwHKeZrW
jg0hXwFJEaPpPnG9z3zMIgwWWfW5yMU8GcY6J0KPgO0xq/NdzmsdthfUaC8nJQuB
03VKX9GpbO9UqCJZi6yiMRfyDzaUUX5PwLhccTkZQ+cF7WvTBiu9HS1MWYbvs3GL
AtRNSAueXuSLRnTQLfOmvr0IhkXv04o/R8rCNJMzr9OM9qP4qbnv3bYIAxrIFwO6
ZKuKXFXv3aCx63GwPqXKklpAFwPp7lgvARYXBWUJoIMZ4hTmTlhYMRgE6KMpJGBO
MY1PpWM2hXm5Gii1G3EplK9fsKDLuZqIhzdV/5mURYL6YFaj0N8pwEaEb9UDN6A4
BHpL1y1lJNjBgmRUFpLJjHhS2BeqLpDAU0fY/KruL6xytOlwjpyGOOxtYx5uT/PD
7ZlIspzvZaijZlxO8N3/nTTWDYpe/hKiUrL496lv+KY/fT1AgJmJURfwYAWLF+U0
sOU0jZLhkoTxeNcSdnQCI1maB5GToa3AKfghRiGPW53+MB6yvVeMg9+3ikQhQq1L
NJw09fz4ifB0T6+b+HjlhDkHlAHx01FpkpMPIuXg/YwvXICFIkkLQ82I29hxqEn6
icSFdBUpUh1Ndc6dusRN+lSOi49PXsN1LD15oZuF/8ES0ariEmkbQJ32G8TXVIEH
D6xII+skIrsQSNJF80lkZTMAsHYYP/JAbWweqwTKU0ZOJi31231+pfoL4trasQCn
TcXFq5ofefTvA84JEsc2dKjPjNse/UU3sSSrlwUV6MMZDCblJVLyn2BpCFiSQGLO
SxZeumvE2Jqhki6QHFa9wanamzuQP4X4Hn4Bwngrt1jwL5ylAuO4LqPp04/4/VCM
goC4aHC51GQRBth+HVUcQDafaqsp/+3bgb/+7oeLC6Ds0IUE3H3J5lYPaTLNM8OB
jkAIh8o6yfWb4oiiAWDf6Ow5YRFAyl0WX1smJYI+isHecVe+MGlqXcpt4xp6B3mG
JZjIZEMCbiHeWCZt6DpshlqTtXJaRef3TbGycbE4humWSVvgF3aKZNqvumi7XcYA
/6fm13DFTC7etplijbe2Rf/MMSUxE5d3RGsakQpknqhTGErvuozSu4XDW/EfjntG
f7NepZAJVc8DnkK+wq1+ekK73nZ79HX7OMXZyO3MDFxS7BE83//MDQiQ08ASW3PW
N+Ug5ZR48iA7fmdOUpQEScSkiNoNXdD40MfcO9dxXwBo3w9V/o8acAna632Z8hBF
5IAQ9fN/dRqYCj5dq8xANIbo4cgrUFYOr7GMOIPcJzDW94iClS30vUuLl48ZpQhU
S3ySKE/aA1nv+MLtqq3qiEr5SkrOd83AotGHBIi2kDFzYGfBy5Cbi12t4PUMr1l3
QcyO5whSh2aY+5q5h+FKkwT6qcsGJ41elsBDONrDJp2605DhyswTa+qw85nU59YI
EpEgiyMbuIL7t/i2KjVQbunIYBwwrqgD/9UrU36nLVamcuh4eaHwk2jfREFb344E
/M/B3XnYJZheSBPMgLwBDFeiz/04wj2VCzMYDgx9MbGxpaE//mpqWEHrCrwCVz9A
WNQ3ijo2R96rNPrIYGwg+8i0pNIOedAeEj9crSl0ZVlmog3qSrsuLVCzLI6fbyWj
QZNXGefTlhCHL2YHgqGFbxewWyjGugW7abAYq6dNbiiYRM1HhJVJ3w97SeeSQOSm
sQ/wyTe9y6BY07Vj35xIpIXX3B+gUIhXkKSgvlxvVIp916HSd7+/GPB0NkDL0KcK
aLuCZVd/yNPHJsjA7iH6xb6M9gY3VpqovEgJARYj66AigJpWsyfOutmYWLf6hcLG
18eK5JsZxw9wiPpvzpQarFGvtS5EB1+CwpioQEkxwMXlWbVW2Ln0E5yysSGIM4vq
cZeG2AxyokeL0QyngMPudGNYYAF7c2g7QUCuu4UkOOq6cFewh/Qb6YPnD/jATQKa
tggtmZTw6tqeoP/ZQBP+6rZjhx3lvhlmnbOu27LNp4I+/ymnEYea0fxmuMdqx8Lb
BpxM+wJWnqOb0tgjwCO3JNKyo8x7xi+nCSFtaX7vcGxctCt42tblOjTw4fspxsvi
RdvkvTcHVq2QOYOHz6gcYBDCdE6cpxo7nGtP2XdJEitirYn8aUmcEGhByLFBRxcd
gUZBPDdgtES0aeb2tpeUxrFsOUep/e4lghQDFoZeRwgLdWS/x2KiWLVp5TJbcZlI
rcV3GRCFRZUt72baRlrF5VxhQSn9XnhbEAt3Z7wUlVe46CUFd6U7Uv7MF3gxcnoQ
tLEXdLcRXjtiTgrxeV5FfU9Uws2VuLJGrkD2SRruiRlekNRbhbVWgsJo374dLdAM
z90VRaW6feDAPB8wcNu4eDxpBj8JN3SJ03couZ0jVKQ59NFJhvK1HUdxJUyjavfI
HWSdaFBzDsSABXqKNWhsmCe3PFnVe64Oy2vK5rr34y5X3vuchGT6rEPNBVYJjCpw
RyPvnv1qdO7d/KTICWtGz1w3blO7ETZhpWhQ3bOA0dqoQtkJwQ+6jPcumad1YVxO
Wowk50mbSV405PxTbPiuGr4eMJtvtL6nSa3JGt7blzfwMzbIf9sTzfcUC+xhCOn4
i8WO4iDPFMouffzUW+h/eQlBKsixCUm8TjMQlOIe9aFBpYF88M/6yVvg9aWIjd+S
X/ZG49WRikSalkkFNrBy+SnOrL9lWmK1Gke6p9sdlp0cmO/6/p9LUFKKHhudK7et
zt9A/s+4jK659L5DJ3lexNvm1fR5LfDAjUpi2vy2OL2L0896HHqFczz4eCCDndYS
6U992rO7wNmZLQs9b3R6dBJkE3ikDzD+hPhKmHYhvAKVFJiH6KQr2vFXZUkl63G8
a2Fg0od7oQXygLqcdkk3mF8Ds+dVl2V5Mpv2cV91vroNCUaCifXyWTtNSn7VYzup
9Ktq3c3/wO8ma9hpQGccRJjuL4PlHl0DH0nmgFx+yTQYQi2g2RijwnNU158CFgrR
hF2mt/uKc+GBwaAwGtYzFmg0uP1XM45bEbphZvtc7WHA3QQt3BXYvR7r2On+iM1y
xst4wOcuyaIEIAf3iU13RX8/onGoJ16uZWND7kQkXU/wUlRq56lpw/9pdMaCnTSU
A5aGSRKkHK4d87X16FMa4PBDPeWEjJdWqpzFFU7W4qsUVZiW9nxWaN71CXywsoXN
HXLiVeDRaObkbSHZwuUw3hHvKPtQiTKGaJP59tUbFrF0WRkNOO4O1qXdKc0Jx5cv
mMhC+YUm+Jjp6rdwocDXBwDYXaxUtHn2tIkZGnl7zRfTrXoNub6ENzfwefIL3rLX
FeN3LxyCXZs7JksofS1dOFZHaOCWSdUmvHMkAApszcrE3JRtIK6HgW360ZlJc4uc
vDdCyOavMeeHScY8+NuWqPoIBFcIW66FQbEknzpGL8RLly2lavBjiMrh5bUR5DNI
q/2mmOGXSUeFHyStB+/+HeyN1wylFCo9uXxjRcksL+a/IN6Rm4lgmtaCM/KJv7Rx
Xf/40Rw3A0nGF35pPLgmIKf1NI8vx7Nq2+M3Y2t6c9f3Be8jZNlaU3DtFuneWYlb
ewzTNGuoRkaD1FoawTvx/8HIeRqYC05DuANb80TqWXw4nqxUA/k5YXrGoeQx5F1v
O5J0tJatyUacBBvgFDYswDupc2kQAbtQyZnNwet/9NaStXmq+8cOVN2tchUAj00D
3Kb188Sw5+fJW2s9ieRYlsGZ+AKM1UVOcSD0Wl6ztsjByIz0pzsV3ucylTQy4TpO
H6+i030liRcYRrfn+2oQX4m90do73qS8TpU6UO1+ODf5VEUNa5VarIWi3qdZzSAM
GEvJk5cR49dccl0giBNXE8yCP1Hnnodg/xUMhYRSV2sKnzJXHBG0c2GF63fub9r6
T6/whrdoIojLrjdBe1tN9zpQ3pdos5SvZIjaAiWaXRy392bG+62JO1Gq4Ay/NCpZ
Gajj3jBeekN88IP9n2IDY5AaHZN3x2lIQb4NnC8Ijqi9SK43wofFLe2oQg9DerTx
sFClkxsW/R4RYQLJo7Fd2VWv/stpsNRVNMmcVmLdHc3Ni1a8uj9zeQMjDHKuDye0
SftuHK3sjiFHUgJHuGSCUUYYkrfjFILX53Uy11W0+jWPTUtn1zvUy3AgM0wsFJEv
lmnopLle3PKFkN9Tbf9oltKQaPjP0nrdyWxUxazdYI+DCPWSmHNTKxoGqaeVlqG7
nb39rtxNDxAFajA4PHZU4W60BEKjCE4qfuUfS7gylKgRyZY/iVHvJ+PAr8oQdinI
t1Xfi5AplVf7Jadn1RpvxrCsCO+Nys2Qb7a5OainosppfBupp5dLukruEmDnbMba
4RgtjRHU/TrVdRj0YBLyNx91HFYm+PQIDvvuZ/S6Ru4T/Z14/jwPjl+YnYLkYQ9p
5hVHfWjSvCuS2RG+iq/SgWdAABYbraLHPpCepTn7a1wzhm3axjnNLKs7jPr/c45e
KZaZz6GO8i9ccp5JSDdsxbDhSVhEeX06ryGxbsuNmIGaqxjlQ56/loagNtoH3MF+
EFQmAC5xw9l89zjDmO52M4Y3XKmgTustQEcM8acnvsOqRu1q8eBGcpj81+3e54tm
zkijAtPY06+4sl2qRW6CJxypw5a3MxUHH6HIVRLYF3Kpc2oZ1Mcwpo77xgWHKgJk
mWz1q4W0pq/hLPQ08vC+CkMcrvZgkonIOa1tasAykAFkkT2XCYYkdmzie0DZWOko
EGDfDaT8w+exZLdmv0mvY9Wv1XVXJ5IxvvQ9lyKhgYw4prel8LDLdektiy4KA0gT
TNGnZ/VszDhKDSuxS6QMTuz7BOgsDUT/tRyxyUmGm34kSzWWLvA7wNrKYb4pPDh2
325cL7EnigG3ZWQBjQKtle7elZT3qCWXLh1SgLRJIjfXjXGQaWhchRFfW9M7HyTh
Ty2k/YFJhnknmAnxDoW7V9AJYF6zDqtApwNfnhQUSkJESUCEDZUZrIlWsRVMw2l+
l6CJe52MknnbZyek6oajdPFioDle9/JnvYPOYLVQbGL9e6R2w0hAUjtVMzTZwCIc
raQg4vKLnNxHFvxBtDwmpq8LSZUHa7fG1PKMgV/YW7mWzXPpTrKy/3Xc9eMKXjbI
fluUbCIk53LlCz1eJTPk1i57rVuoBl/X2vTa35Y+OMBosuCkrjc2GTM0hU9nkWFT
ZgUg6/Zq+3dmURJweVb4pONR4Wvof3DjUr/VgjeV9uJXmiIszjfzGbk6QUKroIW/
73EEE9Bo9hiequrByvnufthXini0Q3hpj98QBsabCZNgk8IGQPBQPKip1na8jZni
72Bo5SjR5yk6XaPempme76wg0OaTae3g/MMNLjG3O5TPf0RzpHjhjOtENkrdVB3w
j7dWz/WVznvpKuFuejKyRumPgDtHFJFePWw2ozPMBbu4nlhNMT7ybgI/cGi/VnNu
Ie/aSWoT7m/x1+kyVoMVgOqllWSSzBUcevTxrNH/hDIVu9iS+13zi9hlpFrj2vD5
+/RgmQ9+FpaZB7Z0rZKroDovcpA76aPd8usw7FMjFea8euN19Cbcf98bOojE/lL0
MLEk1a9iCaR2vc2B85ozCsfh3L9mjmWIM7dQMgclkZEmNlDATm9H4AzT7Ovs+iVN
0W/+AkNHLN0paVvhz5OCv9OQuVg7vw2oc7fqwOrHpkyjsE9Xwo/TaoCz+WCqViR5
dyADP5k+7IBbka4YWmbqzDMmvUhI/HbU5eiJHljeAKGvLAE4nT+8bu+9i9jxiuJ3
Ak3mQ9jj8lH0ANDMMcf5I+H1EzUSh0T8NoYMqS49vIsRpBC3h2cqPHX4laXRNyI0
8LcyFh71D4yWkWqGCohLQABSEtywunftavBqWg5t/j1rujJ4LLQpAYryLnE532Wn
qApdhwfX2eH5k3YSM8MKQgOS87UQsHb85tNEHfysGemwnf914a37lr/j/7hbzfPE
GZXxy0/fMrDJOb23XoyndI4h4/nYSFJrCUgjHaS1Otl+F7tRYNoVd/+3va0bzowf
/rQBmrEi+GxI6T5xTxMRwFsRABO38CbrcxTFR/n0Su1Pwi2ljhUeW6q5hsqGwc8V
ePOmSilAaz3yyxgR7LY21BjDyc7dsM3tLs5Y0bdr72M4WVu+69ip8eRWMmJJYFgN
qW3GbDf/3TbRvlMUm5CIFM2WqijVn23jBTSv0pBdHTYgaIbEbUTEqF1f7cdzW9XD
FrWOi4ai/eWViB/WHT78KhnQLcfp4Xgm+IOZScGpZVvlZQH73fA3df+Mt978FWfZ
quwmQXyzJLbg35mi/0/dA+MBDEWss7uLhTdnwZ+9lkqU+t4Lr2BWbpWNSzHDoNz/
oWNyl5Y8WPVnvPlSPhS5uisPvi3PDe+5VETIQ8yAjlWaetpXKPIzCnmk9nZGm2w5
jMIttWGkzHhPkL+tgdAuQuycfIx5MN3o7+vsONCmESz67OIlAEeSdeyqftV2Cbul
dM9XjJ8cUDkDRaCwzyVDUBHBBz5+WKbBm9Kfrmdh1KLA9xOXaylBNwRv2tp0o6Wv
c1rMdh9t9OpcYsdsSex/JKUJwVlsxppld/0CGtmGo0bjkGUOfbkJDn9iZoXb3YYD
PIHYwAWA1IOF1pOa2EnDLQH91BH7XByYmC23aMcyXvhgyAPDtfk/dyF2YPHPZ8bl
5agn08nImAPWgfbjh8H49THiPpKrAfZiZKzA3sEG66xgXMFpR2U+V1Bpj2xbjFNN
AfNdWNZdvcisxOkX3gn5nuI8Ui8mq4Vc6Vk9KPOyRnKY1rWZqRrelwevpjnaMK6m
0RU/MC/KVkmeqz3hO9MGkwPvw9gwwGEMRFo7rzu/yKH4asnW/MQZbCr7aO6ukJgx
/oRWJ3vZAD1udMAfpHrM/gl55kHxV/7X5/3D//74pCfcdmZjA5R20vaJaBhOsWkK
QcuEbgSLrDHstnix08ZWq9sE+6XsLMhAelVsbGjzLcWNx/fEEz9g8eShpaMmjG4d
NQe8Dz0NmWUMYWvwXii6n/9qbfP487+IDwqNTmkqnS1sIZ9aAqOBp1FBWLPyU05i
qdguDicXPIV4/ILM3Q+aImUbGwImo9shXA+LqoXlJGDBr8YKVfLK7VjJOdQ+qnuV
0FLmsJJLej/ERmFQP+Cyx0brQhaUDWRz6Gb6eA5mo9kZPk86NKNtXLK0fq7PbnHP
xCubPdO9+g5jG2FTMBjg4IiDyZYMd0OuNOi6wwcvkP/JFG4lCmfgrYcKieVcRPmW
VUErEIDtE5a0inLyCinhdXs0Is2QMpoz5iw/6bAL+vg7oi5OZP9dd5XA3075nf7b
MJCo1urizEoBGqjcXDmlKiLsbpzfKZpb/H3L5RnKe1BlIF4lwuCcuP1fFWbPXTVc
pN3T75eYXN3bjooNA71vcEVs1IZcprWnZr4jZZyWOTH66R92PPiTefJPyTDeLoc7
rYQp+3YYEP2GHlvZUyxBWQ5kGUG78itTsnXx/e7X3kKjUzS69QgtRUmxDLo4ifLz
U6pSFpksewdMgeqHFsnjC+j6pes5Aw+CRpz7LBVaMHmfdWCsIlEOoTIswDRWTfBh
qu/AGGTvRWakPFghJ35QgJ2lTH/rjBbeQDGxq51/e7nS0/a/2Sa3nzsFQUFv9hv8
q9eZaK8HzyuOXQJLZuNpcSs+l/eAZV+eNJMZlEmuy1tDKPGaKpv2IWl8QzOt9Eqm
CjgUQylWpg6cEBduFP6Ac8E76QyjdkImxI5fdR+UFvz/jqODsDPCGuFKfTYYNN24
lGJ2+ql4isd6pZMad1aU9x0+xl1mixG1pKtJkOXCbxhPOPEYLsDz+nMq4WXHgk0I
j3iL4ziExuMRt1ZrMYk8u3sXHJFJNdjDkeNVsccTLoMWNFcNJHQooDT7B5oPGktM
xGTHDR5x5JjJISFh/7ZsBVbNtaLLQ8BlNzsjeKbsweQXzQyRlgjvLkTFyceniWy4
RUK7Xi4Q6OtsOlWVaPRXlZ0E0fE02MwxGpnesbkFnZD2tBvT+s69jSTImUA2RxVI
HmW03uOdf7Y8bIA8O1pm/FGKhJdUNLcTa7NACDDcTipBrXT4TeKJOpGwQx4O8l48
uMJGguLkmc4z8gc0XKCaDKzCWoecYgWrMNcUbG2oSlDbPDC4PPxs/VxHwQpemHAL
y4BMGvqvKk066DWm6N9qcqfJDzgJdxPS2jlqkDf5ZLuf1DPvw2Lx69UNQBJyys6r
dAtcDHxb7K/W69Ryq3Kd4Af5J1pwlPDwL7tGKF1ty6wlzTL30fZ7w65qrINiw0Cg
H07o8OiNFKo1UT9+T3sBD0kfPQhAJVEKzMyY1gMBwJ+WKr6dLeamn6EZxlUJVzdC
rahyF0h21h78Xd58yFe7ws10O+/6gy/C61+G+1LLKwuJh9d/5bx+jJQplXWDhmZh
cV2eDL7Tn/Z5yDnOkKNenMnJUKdWl3pJmDnmgGdjpveHZqVfbA9g283uLW9aIYIV
bq7+tXUjgIF2IuISVcgJlnXOz0BWqMAFi5gj1gN6sbwB8seYeHYLAjpknWB/0E9F
JYoGIwc0HVQXbTrL+RwEe0Db2TcObbkafi0kZQLbTM7WF01SCAVhOs6y62doPt28
QqHwGgsfNxoI9r712t+hHKW9YZtAXnNX3MFRXVpooDvCUQdfPWOW6ksS8wSdcdlN
zil8VGyrBdTFL3qrLQ++wZ+jkmngajwQE0U5YEXfbBhgMcqu4tAgB0bVv3tUDGu7
81cwIGzVsca3J1pI1dcVjL+13u5TkOKZDeZ6r4Wvh5jgR+yuftcakeQ66S8O7SwN
Brt5uEXJ5Ez8XDreM/IVwj6QYkT/rjGptmIq5pbAjLybsl2lCVRsOiLJIVNd0Ebu
DGANJj0O+kT79qH2Pnvl+kAxW1eaFUjLHB81y9yHiCKvTtrGa7PNXl/MTGWvNoEg
BFstdlnYmWQnYnMEr586kqsfLRzlsn0esaw6uRQB4teAt2rWCCd1Odz0n4Fj5V6P
4XmnUJB2i7193WNfFE5fgW7siDUzRaEoazig4jgWFrv2sZfsHvjkq9rqO3huGle4
naCEmqlg0+DjzcW3FulKZgDuPVMjA1IZTAlaWT5zNqEi9tpDtEa9HaAJ2y8u1TTK
hicYF/F1MQxpYULD3HXf5hSolur1UNk9yxxhrW3Hvt6r+p+HD5PmejopG+LTqH2m
5mJDRYPcNA582C5nsjLpbtGHA95gl3R7OruiEqAWqSbojyRxHHj/FnYlYIlYLoy6
a68Z6pY94Bg8n4bnDd8bvXH0ln+/vMOPkOM7ByTU2Gv5CDnKna1At8khc2WeFL/Y
B776Glcv4ixqAqsHvncEAGgSztDVO4wNVGjFmj5TSgonUDSQb66c5Nwm+9Y0l7Z5
kxBBu200vp0iBGrnqbEhSxoV7ZjnB01LQOI6n/HMzLaQFGz54o5JOEmIjfEKuGqr
otU4NUq0Gr4x4dLlX4ocoietSYCpN/l9bD5g5fyPvpYGh8LB+l39h7235ok62zx8
TW6wC3kMqlcTfKk6XXKEOnqFfOVe+Ud88Vur6XtULOsRCCMJqU5TLVCIyoICIERT
WOTzIxP9Tcgs6M93robUDaXo2hnPhdNktgKJY8HqKeeVGF1MevAFXTv/XB4qVhLZ
+sgWdFrRkRwmNvVYV9UFZWw0n8q0GV0+bMSmZAQiZXLTo6T8Z/8KiZJxvFPOuUpY
HwwSlagr0k+MkDDOQvC+FuclDfp++0DrqM++agueqoiV4eKoaxVwTbPUMvQU7mKT
g2OW0ir8TnZvlxuvUuM+EoQIQYHJRixuJ+B3ukw7sz8zs7Nno6VWc5HB9HFfq2mT
tQ5rRJCVIfEGMtyo3xTL6ITNTaEvqvzGEi2gcFlvIN55BbWA4VgEqZuNlvYN7Olv
Td10br6d3KJ9albRJu4ckjKWOEnPzE5S60y5Q/DetjMWB1n36GQ6KzLEcRl26GPf
9LiaAqoEmN90gduNzH341yu3AL2Wo0og+gMEe7vWbqGLbSkTUfzXisNcjimIcMOa
YB1IFJHx+6+M1cfXncmmTNJ+JSVR2Ir2ocpNKmo6hPoyxTlHy2UHFw4jI2pFJ0RQ
9qOZrtCzlDggJZe/Mr33Jm+Oc+h8ucNdITmbM62ZoVmxONsUcdVdlhkPGL62+KFV
5ifq5+ZLpaAT1bYYUzLDiZrVyusYd8wRhB058bT+L1wjwmQ0S5rA5Apsjjxem0l+
cldM1b9VS4wJkzpz5kUrSqP72rW46dOuUMqiLDys1zEjKTAsoHhIGz+fxThYSMPJ
Pd70kVrtFJfhGAG1PH6l32qAiwawyqCICn7RaLT+4nvWcUnSwqqUlIT8ZkxwS0UP
/jAA/rHBBS7xgYWlox/rExeE22LH9ENaMaJjwvgaAJZbvEJ9r2KP3eDxM5vTR8Nf
xZMtr8/rwS/vPOyAwLVXiub+g8Glt7MWb8rgAA15s4EX1krTUemyicmm0nKi/aZq
FNjZKNyjp4V+M6WKBQNUPANl9b2PkBe0fF1ekRZfKLkcYvbyHazenXTzQfzSoPcn
BpZsPIwSHeSONK2SC3c2UU3UwXn1S0Z4ToqntBfvAwq9oo6nCuOPy7AXuM0+PwDo
wo/CARMaI+B7ABgCsfqQoN+6Dvz4fXr1j3QQojbY9GbQCgks8JhdE+Jr6luK7NeM
6o7mfNpg1ZHL1NQF1h/t5GYQ1aKu/y8hAuMr2ozz2oA0/cHpisNRicoKge9AqrKM
jcaIDeUde9E7fr2KvGo73XQ0e3gbtdeOYPerSENdS9W/RO4YlyUiYyZf0uhYG0KG
be++upe50UoDX2APow69R/Lu+W3YVuwr/tr5zTOS76AZVJTO3i2cToSHVfTNivsz
xAv/XBKXjAKZ9Lj4COyt0M99kX6dbS2n+r6WKkCEyw8uI5qcxirmRMoS0YvX532K
F4gswW6T4/A9RKZUkmzfoYQ2K62ojD/S53sNYMFKoxbY4bSL+wfZ3q6rG1OZ+6/Q
8oppO9UXxMlWwuspiJp6WAcr8A0OOY36uVe3ti9SCsMbV7ESYsJ9U9ARVWnspVfH
K+8N0jnDXg6NdGWP7I6jlrOVcE9EPKdrLMl3kAp5vK7+YPdI/ND8DOPEUae4aqox
nV0JoYAHDkB2ulKtTUepvSuqrE956KdSu9f235BqxMFPpFSoE0KWv6d42zGQ3vS/
HZfesYDP+8XzOB6UFkjLsASvxQphEQ7xVhN6/t9kvShQqcYhjOLO9K9HDxunk3Nt
NBLE/IPRr3qwFFM82hhr6UFYkD8k3pcKKaAxbcC3AHhcHqV3mNHJtJAY1mrC4o35
oOSJvvYduT4o0L2tnpMkVIxJT5+8evO4rLBVyNjKgCM6tEZ6Qnqhz6ATzOCEpGOQ
MsHpLsTJUo/Xs4hxGAw6LrJpa8sr1UCE1xgBqyqmfHdQVoA637SWB4vzMQ/Mu0mR
QtxPpj/RhW8fUtitmENNMOYchhXI5Lz5+F8HhhZAtudWDl1HW+VTUOF/X+S4ohXL
DolC4nBs5coCXwPNVOK+7mJmEPvfoZjr6zczfnArnzhbmwlbxy8bvHYNwCywbzVf
VQoM4B5NVojP1Uti7KXZYWRl05WS5VY3RXVt6xC4JGB6qm6jdHWHFKhCEvNLXIAV
o8oaeAErSIfEuzi+JUW+YPaGywqeBD0GnhlwgjudOXSTN6zb5MgW+sRGt6z/pza7
6zm4qaacoSEBUz5Q/oXVHde4hKwfutSn1NnSbUlkMYzuMOxTZniEBEMHaQ63QZKD
GX1Fip5V5X+I5g+7tuUZYDf58+izdPgheHWD3HZFqAlIy73EicfRoetsytOc3cZY
8XuM/ZqjQ15zNT+tIANuorU7hs9qxaLIVqG+Igz5Z3AyIo5TOnwRJKMlGwmrt5mY
IIUbfZfXZdtuMabwOwH6X0SZYcKUaufPKAQVpujTNm3gXjeFb/96qJTz2KxsQPwl
flSU+j8czjkX0bN8Xq3PENwhgGsbzfFiv+H1QNk/89klFIIRnFyZXlOli362FA/D
bTO/VX/ElU9iR3XjocbOf4FMsMiMQ5QIWT6M9NRzIq7xILMCEarYZbcd7UXIAhMG
cIl3aLAxTyzcBQVR89D4vTIbeJF6lTuSDzsPYif/P/9nDd5HPVeN20B/mwjURY/j
7gzAy43+j27TJ8T1DauHqB9PMROwIPNACVvhOOQ2mCD2pEyvl/gTX7BbGtHqT2a7
utj3iPAxGlq+IGs84hyQLAdJmmzOfHOIlx8pwRo508Te705eUvsJoq4QMkZYXTCI
I8cS4pya6KdDRFbfXXej/vsyDwKp2vtCwOAufif8zti7F9tmIkNTnQ1DK7Z0WjOr
pZAqOt/Du3O6xMRGLszsyEJaaPKd59uLRh+r3d08/4js/y8IqPFVDQVUPNAj7yql
ztB/e2uf8v8Z9jdQbXRFjJu54nJore4/ePuG8ZQsqSp5BTAnXJU7MgfSOstuibm0
i+bBrR+sKcYBDI46gqCMSezZqwF0Zn3jb1PJlO4of0l8TIyg0rgYIX86J7frI+vt
fbinTZVI+oKlkuQjVseW8uIyXba4SCqPVNaHSNRDqne9eYNiLEVvf4aHcaV0mJPh
Mhe0VE6l5V0gquFCzD8LPvHod/MMgNm4eN56zyj4wK6ugrmXTl7zW5D8gm0Ju9de
YsWyAL4PZa+Nf05QQdMqlSf6FWUCoFL9yGL0GJIOmZOlAFPyX/HvC9xBtkULDz5P
zSbOw1JZQoETQJsxYC3PfgMshapaWQL2hsZ0Fbd+sQpEXfti6JZ6wQWQpNqoZYbi
FQrA4nangG6onov8kwoGiDGjZ2KoTHj5pmSXIi1mvg3uvZNTPUjq3jD6nYozPJWA
oG1m48YfmTfR5wqLncBpx3SgC6ZH8tT3yhCefUZWor1F0mbV9J5BrzoQZfLLzlcA
+vvHfJczRoKnUuyGPeUEo5fJUANYifAGGGxQg+6klqvjRNDMoymkzMi2oylhuu0g
VLqPaiwYlv800eviALowBILfbRNaZFJG8dNSOdDe23cX/5vlxYPC883ZhPGbc/2/
iCs7ksswBZEdsG7W8Pun2CgayVfIc8zJBeKVBer4PYxAFexXWMmDmEwiEdUvqkdp
3FgjmkOq6bL9dQmymRpxAepCTzLjJ3y9+WZiJs8T98SuBNMYrzXljdyVRg8nPjwt
GUXMD2U5vaYZveTGBtwYf2QCXhV2TDALDuLh9xUYSuIqUwmBdMMnDs3S+UBBr+JD
ny9AenW5hTkXg6jqanq+riDMK0GsqHjGAq717lT6eKecVm54ihNOrzZpR9iUEz9u
M6gw+J8tN+Cpr244J/S78EGnstKZih8BQGuYWrcvsRPygV2bSy7Se3LLT1oqvDC1
vemacROk9LJgbxlbFej1aZ3fBGAkIdIlxzhS6U8dYWzptw86kHgEgUgOMIJ0sYV3
udTQNQOr++XIxPOjHvoZctt/QPBYss2UB389hhIsd46m/pIhJKJSzcyyutYRt38r
i/Wp5gnJiRFdfmeueFqfxKWCoaY/DVWigKGDJ075Wbl/UP7KZYG5NWAjqqV38AEv
c/yWQy5zRyUjlEwNZImL624xE3/tiOvU8U4UUulCAjWzSLlvcyWM1UAdxyT46mdm
jPWpagkj3KHgYNjROHB8diHXj7T7u0PKLRkSOFZ5vFEzWUc1fM46/juE8G+ErIXK
FB+U4dq63ifRGzzUS1g6jdQL0gCvWeYVHa5EhEc8A/e0bamW0DaMVACnGNGf4rW0
2HyJKVE5hnMuT9KjGs/OR0SrV1s7hZw15lfapyUaikWcaTDIvxNElZexMxHOxbej
3hxGuucpwhWAjpQLTe9BdeEwCKO/eJy90B50E3NdZ3gzkivtxLknwvMheyJvki2O
Dk/WaJyD0cczI0UBNPR0f+OY0OBpyHd2m6QTcsdMaq74v7iQnDKsS1SmuxnFlA0w
t6cj4DSUVVRA212uHpC6j38447wDRTgWp6S8c7Sf3hOx5DiyweFNQ+GIiTTAx3zB
QAXX8nq6RaT294yv2qWqZtu/RukE6VXpC9viIBs0Kwt+QiqHraVzEa5aDmvzy0Y2
QJSSJlXQGWQhZVeHI3pPdyG3/L8uDRvSZq0IY4Ye/JR9hbLjrTiTMeGqNWF6Lyy8
TagyxquJfIdzvffn8iTLl73B+LhF4euhAAs9jn9M4xKfoYc6YPRJq9hXbl7iaxQH
3RJmLkB5erQm/2/IO4jIEX7fMVe6d6aTCbjm1CqQY0ujimnirAeq8mbsat6nNs0W
9C0fL9ffF8XvF8XAHWHZQXxlQ1TScU5j+XGdsFA1IbFaaPXpB+XnkVHNszm4vHRq
0Md9lqZ2zxkQMyLKLuxC1H9r9R1+j+EXtWGXrL+q9vVNPKJUd7BsS3hb3XXmsEYu
fLgUWOAp1PADCyLFtF0wlFewu74xXVu4rzSIG6P9HcxMxWugxGMss+bcytebsbHN
M6+oxThmrpejWGQIjmGNwiNYXwonyrmd8/Cchdo7T4RrTOe8WPqJaN1x+/hibi7C
aK24nP36ERf0HJgI4YLeZ68rc9rBvcBIa4pimWEuuS93mSVggGnxKrowTU1/NJcY
6awxkcbqa3jYChUYeg6KhdZ0Kr4YlAp+wYjKD/Jt0xbVjzTHAcosCTZc9Qdj243H
L8Ew2alV1GjIwUsLlFtiNtsor5KXlp2+4l9gwaTTfyOHwTj0Dd9qs/U5xUKpjNIT
3StSHiYgyacaE9qIffv3SUoOcf9xb5mb/tJu4akga5dKuFXf1rTnV0xrLR7evDg3
q/GPG/Rzfwj0h87w0MpkVz9KMjdc+xKDkfu5nlDf9BYaMekic6nj/LknDox1JLtn
AzICyc1hZyWMwxRuViDcTHIJ1KL/b94XPfLvLO/1fDdwH1yU8RZnbt9u3JJdFtYA
TmO6kmc3Sz4cmcCj7iNuGINznlGKeqT5Qh9H2gwEvDmbLdrYCsXKGGqWEfjpMuic
NUbpzb7RFvILIzhU3NnZ8/heA2fp4704LUCHXqeKPBCN5kZc4eKKRTGjP2RCUMfY
YCTwTHfcTrmUBN6M+VbLGmnyR6ItTxfG3LuDu9axyPo4lCjUSA/AAC0c3meYYjLt
8ew8sP0ySCpeGghiW8GWIofZsMXddYWFsfPlUkGgv21Hi2j1QIQzUTWeBfi4hiFa
VzHO2A+HEbfmyYDjNCcl2A0ZvGThKB7eyLguuwYq2TZYev3gPYcxILuVAfn97hyp
g/o/NF/jJmONZIREJkDAEq2lDCVnA3Q8YMRAFf4VSPJLypA5livO9LKeJ0faotP1
Q1rncwGXh/l8iiz+lDsIIqG1m/7KgKd2s/qpDOPworajiwJ0GabvbhXUiWfSfBs0
YdPwCOTymIyHN4lJEVJPy+LCuNWGX24BmarsgM1jKo8VNNvLgZMT0lk5cWcpkzTc
IKdXIcr6th4NOxGSS4T0/YSUz52+Qf0yzz5Gqvg1DGORhoYWE6GHsyHEeShx/fQF
VDo/z08zC4/Meo3A7moav4/uHRBIwbD6I/WisGV3clOY7NhFZNJwX+j9W/VtM75S
FgmESaTJk0lVN7csxpsT+8LmdKU+P9waPH+sKzLgRT4a1QuIL9BxHW6bnJ4hhLEZ
C7EryeJ8MbU6W/vzmyVMBeajuaHNl+Dkcv9VlI9gV3z0egUPmqNPBEgFbe+AwY/U
46EovpTnAYMM3t34JfvG+b03uPPH5GOPhajvdQV7LEnlhp/zEQRrTR90NuYG1vI2
PWjUMlW16K2UjMAyDWtW/tFx9IexcyLAGNYXf0ZIrXGzuIVVUvAyQWtCwgjC6vvL
/cRWzWm1F30lQzOu+QIlbEwm9W+jsuNp718E6W9Xnte2kBtwNzCwUR9e/gLfbo4H
bZoIDYn6NykXa67oqiXDjttxwyOBlUpiTOLWOb4eN5djruP+zxjSxpEzStJkhoZ0
f6iIfweFoWopbLUzd6i1IGC7IgA+j6oxU5gYJMhaey1sLcCEHGsccwMBYZQow4IX
d4RUTpkbtkC+RlEOOlvrovaWMFxlJtLuwt99fzl+x9dmx/aYjIZFvx0P7hHZUh3V
VB5PhCD+KricnP6+piq9SJ0PQveV9shhGKoK/A51drH39ic21sQngXgT5HX0aLf5
KVZ6Y+NTnmbFT2UKLEq04pdE1ugD6+Gv6xb9kRs6CN33KiKoJgB8ohwAvI9SAgo/
eh1RBRdX3qpnxlqNucXmDpcmZu5Tt61UbxcP+q2t3PtKXqUxXqPE2fTga3jiHRbo
ou1vAjxYWE5DHkN/4dYD9t+un1Dg6oHf4Vom07ULzW7BarueRVuQJoIS1KgzNHFZ
IL/EW/WVNGlnJschnE+vBwDPLQ4cJa4U+Wul6UqOjdtYQMQb89RTM69i0wQUJQHL
xTjcskrn9qC/CNkfNJMbMZBzmaA+uAtO7lBpAx1sbzMoQ63UZaa+3Pgs7tpb6Mks
IkdHPhD02+EVEfMFyMTLDN99plfOBOt+FeHYIQWnM0kGBza4T5fzv2p3X8PXeFdP
VPCAOtFTIqBOOPzeVR12bm/q4mUvz0FXyjeAWn27j8spVO1b2EFnD5TCU6ZiOx+C
tBp62Hip1F6TWFGkNC671RoW9GhrBfQwtqitwWSTzgCrvi2UCtYwRAM9splsRALX
Q16X6qJIZZgL2+hCTe3M13uPNJUNG0LBIrUBvDz0PtlSPhlaEfuv0lTlczUdhGsO
ZaEj76oAZbJexCC9oA/G2S3tv1BW19JrpyltVKZxcLVbkJJmUEcHrlE0RH48LE7j
ye4zjnJk+prHajNfPLTgpHmYUGQTvdS7DuYsZmAxITIPr7hh1lzQNFvxgZ3YfSmp
Xzs9T9waCE9lpskcCMCUNlzEPWi0a8OiR8lJY8fiXdIrJ38lnWz8GDzqACSXeBrp
jHDbiOEMOYy8q00y/lDaqDHWj6M1mzGDN2csXYnyRv9HDnbOHjij+yIp3szK5KRD
92zFzmtxnjL4XTd/BYYZ69C0Ste0VIAxBEPvRQlslkZVeKPwj+Tl75E9LKWr1yP1
PkrVvWedATWx2UidJ1d6SY00jBJ3JjTviEHG8lOgkjKWr6yBTqJP9eD/ZShjqRzF
cM4QadjFLpxcht41vY597MUJa9cLEfWchpA+7gjw9HtAc6TiM+IXtN+oeDPV13E6
szWR5n8znl/ne5QT9VrlhDPBRu7n0DHrVwCjrj8syIRjJGtOVm7c1Huld9lrNfxN
r90YfRYtNyI19QvonAf3DH1sS7nC7D1+uiPrFrsc7uTxNrneSNd84/M1z8d8l7VT
AgXkfLDiI4uEcxKy4OqrMSI+fFfugwVNaSC64H14u/COj1ucpEaUM7PmMXUegT6V
LqPeu7Kpz8BRl1EKl73WFbyG5w9t75tCR9Eht6YcIDVNjlPN7Kh4sXt7hTKIBCwH
P+TBL6nShA/A4C+N+0bmQMigH/x/7bxvbfDBEopUcSUVkm1xBKJmcB6phBECh1Qn
DoDDf3VoWari9WaQsp18zYtSMY67yRYQ8snQJ2I2cpgTIxMWsNoGGwmXEflw8Mac
a5kGFc15tOiSV6FjAr5WSkSL+wa1kJKR/NUP4glLDm/tOqjCKPcufEeTjl0bsHPv
biXD8e/hheFwvq+lP9oZtA5MuNDlZAV3IOrxIgtIdP4hJWdXO2U2pHjCAG2zeChr
H1xlntoX0LfaehGXrzZOIaFuzUskt7Cz4mqosvvg226yJ8JxiH73IRqgQqvOrQwe
T+WPCQfmlO1KhQ/1egwinxbo8+uOUyroTfIuMFQQcJdLKEFkXkGJCC4Ge7dRUPnp
X0RZ/1B+Edp3NMrT1A8otXDEsUyMF0ci8cWllGIshniiFnR0NbO5qX9uIi3tOxhn
HASrkD6Gba5AnSOI2E0zBhjLUBbSetmvWhoXAS9EkVMcwXksQZbT4xe3UlDZiOwV
ygCdhGQkQD08HwaY8v3Gtf5X0v0NW1I6Ol69zckm0g3CLcr9KfsIXLvSgzQHZKs9
RwXK55fAdGfB4hmltcZQJIuRlSmP4f4WtJ3m1yTfoOQgbKR2yftqIkl6ICngeWd0
FJuI6b5MldlEn942/XY1BUjcwaTpIpwv1tj39FFgZ4FUBUo+nMmlHfQBSq6PX3RQ
MqE0BONmVSKOVm0Rs93ipsSMuFWYAEnuWsZFFviWp8Q6kIaF/Cuj6IX/Ui96yVuv
vHNeKTBo+lWWoLuJw5EyC/d6f9NGbOdFDdI9N46066K2dLJosaKdcI9J9zsSoItC
OC7dQ4nAbrwORis9j/UTMDgFb9mMpb3o9ZNfQOAag2TFDsQmOg5h4meldorU9mNr
NbuOwFrHQ2cNjUoMJZ7+LuqTFijWK42dT4hTVhBhCVeu0uGuGOfTvLQ4pH+xPDHS
2z+iRu+D2ll5YJbAS5XWAQmmiced/4YWCXGW0Pl1I/RSXMPK8Be6HTGx3xORjoFm
na141P1Y5I+yLRhFGCUCXXpVz6XnLGTJf6RDF/ZG6ANfyOg0/Dtb2+gBnRmpl94J
JK5dLBWj7BIj/Xmf25tBGy/smW5IjyHcJBDlfa6lcKTJvCoPJ40IdYa9Qw1eTTEU
GgffWisc/gdB8D3EFuuPQwI9IqPA2K5iQKBMQsik4jas63Q2aQ273wqnyg5jEgE1
8QWiNz74OaINwDxbUj1qCe2qWnniKEriw3x3ZhbKACLnonpyaFp1WpvLpB56eZ4m
bFm5MegQNCsEn7X2OmDcccGw5zxQm07ZdTija0gjMDqxHyiuY4SRoghcwZADM2Sd
WdJEM4ge1KjqzBnkOak6qz/KNyE4D0V5Cs5NFC9Kimiqm6ESeWtH3Al58MLUam0P
5CC0SFknHlQpXMDSiv6nKs0DH/OhyvkvqjadaYjngcBWelulWn84j7s84q+hffWv
RobD6qp1qxUNtc7kduSJBLuRWfJn7Mc7RripyUO0llxEyP9n+INGKf5pQ9sJWP3D
o2WqPUq87lFD/6XKka4b4ATt79XTp1Wb4bc/OFIMTFUWey4XjPxCJ54UVoZxsiSX
BhnRX1DRTTBsQG+4r975sfXgLjua4LWmJmnBqa3+ZmX9bfGosMH7SlidjqgK4ku0
Z3dB0RrvCzU+SSYwxD8/EHbWynAbVop/DupCpNmYdo3HGP5HsI/AKLg2MMCdzmjp
F+bQS2Zv938s3kBXYFS/bur9qHcKZmw6Px7/VvV0DFVEkU9Rv4xJb/n71ODNDfE4
mMmBQpw4XXXObCPLlJYcCOpb7RETHuqV6jiICpnhAANkKWv2bkV3RbI8hDzPiGEd
ifDfqhrWgXxC3s5vzrhCtA7XTaPvV0SBRRUHLAmRAHq18frz7gTHdV5RQzprLVF4
C3qWArD3ihvC4AXllgw4Tk83rEyf8yNqfiu01b59T9BkoXpDWUp6UYp9FNdiiCXb
CDR5i5kp/lMugVqo7K9zcAhvAqwyDFTFIbhaX4YveXto/bGq3w/KvvEzz4iE/86Y
01O8s2Cd6htZz1stltJNqEGIZRjm5Qd1lLCLtnykLCtOSwOx93LeAxzK8V7uI/AJ
Kaictmz7t3WuyKVjgWBII/oW5hDJwaI93Undlw1dSBk/RO1ZRj+Etrm5c5ejyBgR
XFB4uDvC1Bv0ce+HCgm8IO1pxV2tujOBSHlL9t7z6Pq45/1HyE5f1zMKv6l5wL6s
RlZHBi3ibeue19StZsMHAJJcjBR4fJsgsZoQUVmlQHG9/gyWYuHGCzDL26ItOd5G
CZl3nLIwaycY+icgOAMpEehh+R7X7MKpTVvMVnB5+5lLahJPMYBbXImVN1IW0wld
oiWh7AEkO6TJQKGelkJKSNOwhSIr2MTBz6GzfTPHZXKqyn1rsby7srMw/4krb//z
t6ymHMrE9uX6ab96drPV7X86kv3KQzKb8mFcFdVpUpvpwMovqpK0r0xXU4ikABI/
LvzzoUjsxilDjb0ZNzkapyS8g69EE1BU3QYpML52KL8LIl4YZhbAOqNgl3gjKUgq
6b53o9mzrI+ofjxm6lmXfZ0Wl2XcSwiKohGzhqhTQtpeK5JpdKHX5UEUfMC1Uzf3
Nbla5EvK42qvjtgBmeBQJ7voKsDhAvpx0oOLAhFaemY7WL7cfH0MWS1oyEwPZVQ5
wk4GDD+Mr9iOC2EVHCij4h+GIliNvRJ0iR0j+MUecduGJI6T/6skfqu/zqd2ZdI7
86crQLkpAIx5aouU226zJhiT7j3/UXt5YF+z64L0VD49DgpUJYfVklKIcuGXwQ9f
dalB36fZA0PnBYQpl7EoAjbZO8nfNyLYwKI63JF1Z2nTv10WnGvcFn1nW+CYolFA
ZgfA6+rFh0nUHsCQSOvg7mFx3JqzqYyUDpz52u60ggGOKLfYP7Q03yEdRhQu6ynX
rAxv8JtVpT8SDr/YIfZZ1kc9ZbGEInrxGapzC/m9w+ZFX6XcYXxI6iBHIb4YTTTa
dut+fR1cDYDu6Cyauc4DcRbjV+FftZ/yQ7sPDQpSueYKCNgrTi4tSdjKguZfujqY
5cqPeJiUBxURw58uBdqzySMJSZGA9Gkm2L0QLe3emnycoONcm7sH9z+iiS6b4xqB
BYUMoPWhNk5ohkvekvos4FT7zEzp0BpIlK47kBTC2Grbs1SYfjXOhY7iSLw4u33n
ERr+ZmgX8ZWcFj+m8O81+150YcVzTTZqjGm8BhsReDsKuCbgiqnB6ucGotSgatSq
3Jl8mkCPgS97xceHggN9LG5Pk0o6ErtgxkJZ9qtW8BH55VG6lunk5YOXrCPUvOgC
raz41HZCTtCAGdzYr9mYm7OkOEeMdk6mIEPE0EU+PktEUIHDl46srVuz6jXwugpA
F9c81aNn7O2lEpSeyysKreHUouZgvjJEG4njAmTr5d7Pdw3TyZhWV1xpxxBU5fkn
uJUP8xHQRcRxNq13x2ELeTpdftuYBzALbR6IUJm0liQzBHA/vf7wK38UgsrmkCD3
XYZPiiAJ/TXXLQohn4ddVXCyi/jgrFXtunUnafuZV/Lxs1GaKf6NvWV93Zq+6kHv
DKAkM1QHEpWuhhFsgqNbWlpk/f9xKCZRiEEW3lUWMarKHRYD2tA0b6tpea4/KqFH
lPxkjV8FJMnDzRFla95NVnKeHhakCuu2ccJeIJZa6lG3iUW8nITkS7HBGWAYo7gr
Ds7/7wzfSDrdKEDI4uq1TgL18g64SMCQbYSWvhPSJoU6WjHEqJc0Sfp03IYWQGKh
wx/J+SBVkGpOyf3c0mWt6MfQkxjtfoJeXC1um4ra42Wt03PJh9Cr6lhuhPjV6sU7
kZRH/y7aSQSn9mvHBG+N3Uwerhun3b7jseeIu7x4fwkBtmCBSZag3SlerMyKJ6/A
KAuJD9i3SYnzFMtra/6VBYeedlDXzIoYgdJAZzV0jPGvPNG7Nj35SCM31dkWYiHK
6dWphHCMBc1PMu4O9F3SUBA7s1xtrYZXB5iTCd57NaxfaAlRLCt+YbqIpDap8+o7
hDNTWYgR97evXdU6VGUfaNtUNUwVhmCF+CODO2Efp/aGWhvH4+biAGPttBv20FOW
/f5581TbDfbkiap58NcUfvXHlN+w+bi5A4zUSBpagaouuwLpbqH8aLQ81TS6Jrp2
i65kFXxJ/2cbntRuSMZE12oAGCNybq8IeueLVf2jhCovJR6/XET8l1wBiSAhBQEu
bDmq8hf7Ee47JwP0AcZNZ1ljiQrkKZ4kOjY5WqAokMHkbRa0yy9PRTrZEyA8SntX
fXgVAPam/qsAfW4Exixw5Xb9xb6QrPogxNdQC2svWeR4bq0xUYHeC5MxHojCob/d
2NWKUs4RN5oXPnLVXCLNpt+pJpOnNMu6Pu5M6QalSw8IeyT7CB5e6GkcSVoOG7a/
Tn0fKo301OPVWtMqHqMzAOjBVE15aEMAVNWQeOoKbtDHI3DM3gVGMNbejVoObEhA
Vj+Q+6yLIU7/Qsg5hBtLCA9xcDaG+XGAJKXwGO0GRfEnzdbkkTlyCCylNKpwUNyv
MJ+FhBfoS7V04bMyQmYEybuT1eMgVUsmE2D9Q0DQ8sdknFJfcVfwKUv8JYwyM0RB
0c/U7st2z96KdFjGe7pQ1CN3LfLgTZvbMyhic/v7DXgHQzPt2xiVDvbpX2EqVkj0
po0dA0TpeCRO9uK0o+0IpYb9AzHePip5j8G5YwWRJo8KhXhuXaYLa4dPF4oSfMAW
fDlMhqDuwCv89yJU9iwkSf9sVJRb05I6dF4mzQ5+abE9zjcYhoK5289BBgxedTLO
rdhyP+8GHgOWq6VT5VFhAh/0LjQsQJ0D7OVLq2ICxzzk/c1lpq4kichYoZS6zEZ2
Rom51b9SNaVLmeY/JKk4V9W7CWEZTOsJ9W7qYneGhXEO+gEZjy+5/sGUIS3fxkS9
yLM0f62U8Q+mVNS4PcqePTgrpRvDT2IkenBcwS2upHcFnkq82EJ015e+Yz783DRf
VdriAWpwmYUcuCpZQJm4TL8HwuCAZaBUWloRFVYF+8spvQI4DUSMLnbBSZFaTk4b
AkSMiSqEqkoklsK6TuO+z4BF/++VrZnTSc9k9/BoGJe8i9aoFW0WSPWMka8TXPEK
2YgfqhMkVxOtM4x5nLyzrSpuniJ5aalDmJdj3ldhfgJKcxBpIXiorabCWFzjIw/j
eAfPiTElw6wl9QDEN1Ug9P29GGVe/jcUSyhafl7+YKW4m6bwR3Qe8Erp2ziIjGZw
QSJgokg88EwtojP/trKK5aXIoX1ySEXPTcEP4bwDsG8PEc7t0S8cI08n0k9s14Ch
mKJV39/DGQlqd9sRuzpbMH4k+r3O2f53bgUtKmqzB1OfOX4SjAgyprOh/bOE5ZgD
v/49i3GNr3Qcx7A4TzXFScgYgYVA40SRmC8k+5NnCV7HqDzY89YHy42j1aRZNHRh
0IEU8Ag3ATwxh0xraIjARhx3C7DbHeGk8rg75RDflqGrtWA2AEvxw6ZXqt1jHNHO
rdOm0nydRibuVIV1VZK8QChlpdHIIcwgmj3K6C0KMRQuQBoHJ3K955LCO4Sf5n7O
6homv4F5HFFd/nu5DLk3JItti3UAO4GxnJTsq1qBMb3ckfubwgXHImkBgIpAzboz
fikKH0NYoXReQW9xu4/gJYOarisJVoixq99n524F+uzNjqeXn7mwCbmOGYFp7Oe9
o4uOWWowUko7BhKK6KP+NWZxvRA9qFUiYm/o+Uk2zwLTVHUC+XWW11S0kt9tNn1B
maQFeDkvmqxJlOM0A/lq8JRM41BwJ/PgD4xjVIeD2IPcTs3iCpkdtZbGiiIy7qNQ
WsWhH5VjFyn0n32r0hr3CichkRNzV1rQ+kmucC4mk7YbGpHDikK7ohWaDs98R/b9
2tyxO9kigvCGxvJIf5dV5SNTFwuPZEO/+MEhxXjsCdGwFy9yjTImu4ctnniTCBC5
owLkPvLJ7AfJiQlpJITZz/gPiFjKqwHE3TJlSB7tUESXk1pGkXsd9aZs2JxX13cO
4jgQJfGlhi//+fiKtaYfC197Tk8fdIV6jUjikBZlvNfKNfGXyYMfe+qg8GEw3piC
pvIFrxyH75pNu55eY0QWi7+PcFhpOHuN1QfhvZHmKOWYthuVr1B9He4vTlYWKZmc
epIDHiEE2RH3VmI9uqe2v4J6KL9x9K88e/B1AqMSxjG0l9ZkV87D9v+Bniy+gqVA
bNrnmJHOTprON+TCxjSSJ28Hs2p0RaP9cJabIwAFnCEWkj7mBSOC2wBtKT2y0i18
JC7YaF6Jz4qTqU24Qp/4pUvCIk9fNwkGExops76MuNvEPIt40N7kmY1uU3kUulbr
Rpw/43ykF7zd1oQxQ/aNMqWKgnpRcwBcB5pjO9x9eazu1s/yd2Mub4Ii0JtTZKRh
PPtRwfEUSl+GqCMzPsdVNhj6NUB4qdJR2tzDHxKT0Gf8zBCJdylwyaQwP1iYJME2
8N3CZAosCbqTlqS8w4MkZyaBslrjp3DWuisRm6U+8A2m62qi8qf8qXC/lwjwbfsh
hKKBEm/34j65ntcPbDCZesoKj1jFPafYFA/QnZ+D1kV9fRurZx9hQh+tIl3rD7qV
or2ATn7lPRDHq+6MyqNOl/F44oUANjxd6FY+DNTpJZR2hUSNV0bRYQn2Lo7KsLAt
IeCC5AChLtKEo12VDCPF7Eueg80+TJejGELQ1QHfAWk1Tl5PvAu+i6yyvNHdimd8
mSBBtn5ILJRdI9cuV/ZuS4yV5D4ZUL2NDoq4yA7667KzywkAm8MLTlPxNqpGQ3F8
I25uMOlnv7itiZzkF9lPPdtq+OAT2fFXiyw2qcNmn7HA5vyrTqxo8qQJ+N5u/55X
Ft7tXARUU5oCZP4R/3ifiK/oxVoRYSfNBH9iefMeN/GElLbKic7OlO6F+W/AWS5g
zXO6rIH0v+90X+1oB030csuONCXpmz3fsK8FcMMXhWszveQH6TnTOFlXSPiigdE0
2fCO4Hp/EXbsgy8sjp58jqrITI2Q+F1HjLTIAMXsbGJPUtHdq27WRbg5KF2hBH9a
WhmhKpi2ayY7jyANM+K+vY0pdCWQGZLg5FgqitvrjQGLeWGIzr35MdD/8s72RTbl
akuoVp6YAK3vhPrWlvPf9IszsSlXtsNyWB+WBL4UlRn0P0EIetC0LLE+aeayKiCh
qGCgucl+XOrz95TfdQD3PTmWYTxdr0E7aKf/YI0JaA6Jlou3FXCWtqvbYOgE+Ng/
aCxBA1dAZDtJiQhyyjEbpL58RW4vYJvV79bO7BkHS9/YKqaPERO9kJKJSMn69ZGO
wguhCsTNY5M5MeOSomKIVZ8FMr98FMWoL5tm5ZremSQOc2faweTdeWGezn2jrRfy
k0ZoL7sLuaixP2VsOWz7KWTEOZR9eR5fqvYwMami68hAvFUjrFxD3m207c0M202q
2PJxYMqGhn1RcABnCOvnTJcmX2DXDLW13jZ+eClFhjNruhknmh2EcTW7MuYI2x/n
qMtKe6SKMbGAeBjrmSxXekrdepq5iBbdwwU8jqPKa3x8g7Is17tn8olQZSq9Bpvf
+lQXcwOSlrTv+mL0v196W7NwbkXVGNM53q36cyJw8ToTksfvy9uLOR4AIQpI7dpg
3Hf6Fm+h6kTpCNdJZkIS0jOZnEHFbUcamb5mMk8ky6PbnK0oPsIUl1qEe5LiifA8
2TxtmeJVvFUqsRr9sYWFtyuAmtDvgYbjPc0b0Hh6ld+ADslnaMPrGFsk4mgnyKyY
BjsuwhvPZRcKYvWyh/IphzMmhF+3ykAW5ZDGg5TEpOMhK7gELopq3RQjt0LW4/zQ
bNxXVTBgzCmigeEmTe7oVms4ZDqICEYrIXPyASIIfMR1i+nMwdnaTqzUKXDZDqlv
rlUmBvUusySQSVcWI1K6cp7Tdi6it/Hdhf8z+8NmgpIx2uRmUgsrl/J9yy5cEgRn
fdCAfI0J35Pzamu1XR6z+GBgqkac3CrGoKiyQ/MSaZNLFVeGzcbR1/fg6/Iya5IB
OQCoMD/OkJfYyLoxYsjrXPRWFHE9JNH9umdhQgSKf24BJvZIQdXhYreaj4nmaLRm
qTjuc22M1xTv6edX4JCsBLmpxVAcZWG1v42xp3LaJWr7wfQXEawyUw7ZqGjMp6GS
zN7kxGTB6NbQTiPTUp38eKJ4LP0FWkh8RJqpRc5MUGjNZsrafpMIlRN9BFL2JNLG
RplkdQ6qP71GihgPkrIWF5G1fdH6obP2FxSxSktc9iFT+gmtV8FRfpT7N63vHH+g
ptP6RoN8eaGawauhK3obcy4IjCJSb4OK5D9aQOz37m33WSnGFre2Jo3X4ikl/hgQ
U2H/znd/ou2Ft/rL3rYmDWk7m0zxsiFSw5+9P0jS5DNjcEy95r5ajDl1QhirZ9Tx
IjVhuTHLrUM4GOt4JKTBcqmjR8wrxjqRqtAgbjYdsh0ejmURPw0oPLC/rJ/zMIHo
PlXtkelRxQIlSQuelv3ckkcG37gZXx9nl/t6kCm28CQmUmhICdAQ+H5FD1qunafV
WCuJzMvV7mUNByXjC1AKq7dDfT38aOnX0t3Na1TZDUJaBmC02D80nyibzFbubsSL
/Ndx6E6XhnZ8yVEN9nERY/Gtd0m3sg6spfDC5h2/MN1n1eXYDka3myUTlrR431ob
V3+LJLx/1CIpsQE3UN2L5GNDAwSiyWNf4HSymTigJOoPVNv+282d+rTx2TSPRzCj
LTLbgEVymLfECjaltQUbj1AhcatdtO5T68ptGnn57SfGA8S5SLOE4kXOca0er/eU
10SS5AWBBgiwGz2vFtzquasZH2n8s2PP6FDjbmepmGcNAYizMPz0pzlx6+/jzJ0W
znrqoATYN+avZ3WSRKVPXo4XslIiLcpoclbGBd6knIRlGjDUUg6Sm0gQn6EOp2co
Ll9jMzcE4a+jUTtEC0+Jqv3SkF8vpVWvOP/RAhFalYlXE6FQ3KRkRdNubEYsi4Uu
YP0ms1xIzlHn3AnJTTf3C+1TtfSJC0p6t2z7qUIueClmLNhAUgO2hocqIJOKUAqw
YiFpoOJjqmS3NeOfnUU8xJ65c9xTSA3XPLGaat8ognFMgVoSsKnez4GbY1XiY2aQ
9eLQXZt4ZcqcmYC7imtK8NOAsNy4vmhcztduUK9NhwpZGnm/bDd0Qr4IKM87UtZu
vGTYMQqXWP/9L4l6i+aN94oI773i28ds0g6Y54b1TsVcsI/AOIvqUym4Q264D2//
4l/VbDIcdT1YEz17oqR/F0lW7v6QeDpGX4/e9RTMmzvOX/BCMLTCILflrv38cz5p
E/HFmXACFeWYsmdfsgD2afZLj9MrMThW7D46l07BCBPWTz7Tz5j3mDlXRGVPPn+R
ACSyS4WgUGIxbYAcEa1UxXr345Zqypr/XsLRfoLwXkQG3w1keXq5FFDfPL73q6DX
TJ5iu4Qlchcfior8s8fsY5qgOvOuCmv+u8BFjFeGrMYSToBGmnHaLg8LgS6BQ4z+
uiVKjXOcNd2xYn3K8vbDN/szsC3u7e0TktV3kHA9OhLO+IoRDiim3RX4zbO/weX2
c+2lPA94vUr3p8sGtMM4SQO9VEcaoddZgu/kjSK+GmA/rbJiXyutZ6aIv+iD3s10
hNXibF4mFP9wSs1yvMc1177liY2iL0vLXp37f9gJuUNgph2JLPPHGXKxVElmnmf0
6zt3b+cQRTWlEW8k3MmY05iEPi/IwMx1vSaB286MREYXMDyWLZAfqaDwEqxBE2n/
vIt+I719l9qEq23OdiJmHiMMUnLbm54m7l9niXlSsTus7NkVOafMr2RjGH/P8M4R
9SnaPNIqYPckHpl3QZb2aFONby2MqxO0WUYDU7Cla50r/tGsRbbzoyKWcNZfQwk5
fSr6l32sjtzVn+BXEAZCZMv9vN8kz4Rj7IOLSBfhaO/1oOXkwYLxv52AWGLswQTP
tyYP06q3UgB29tqMtn03zdHXnZeSiyBFzbl6Jhcb8Di7PebqrC2PKT5GXrykeLfO
hbNdwhTFncIpdlIgJGNsaDTHCDitck1NMaoCFAmEhXFdXJHf6s5MYGypaLB1IUrn
uIILpxkMC8IGSil2WFWbe++u+sGcWVCHHW1dmCb4YPjP2S21EZScnedZ/CfpzWCl
5IdFBStfrJsvlY0O7h18peGSnvtIznZ16W6+TYb0lRxwV2E+ozTghOHBjuuoxaJF
j9871F6jKgrGhThPI405fJhJHNv94ipHlcjQa5wem5nqQElIMVPvrbDmNRIz25kJ
fny9XwR55PI0CXSpX+euhj8zSYSTlW1TWQboK+f1zHKNLsN/aAB57cUsNzIv6RNb
0mdnOK/7i/vcJBPT90krMh1jwl9960VRo6XT2SSE4QoWFffqeFGRm8B0jH4E0OsH
qmw1qtIYo3qPLCzfQ2kAQzZdy0EtyUKfc/Wd7WsVqgPSa/57dxhJLs+DEyrYXK7u
bXADhSm4lJo+HLk/DOZO8QMVaeHoGFVmlhAB1pQ8eA+Vme+M/fzxu30IjEgqFIef
z321pNXG+NYLqJ5cQsSWm5t5xZBVHbQcDrJUM1Ql13XBbZ63nJyuzeiMzLPnJpGC
oGFOtUM0WXB1eVSr2ODA3GrJR7lqtNGzEG9ww8XTeeM2lfVa5jgnHA/wCxiQErRC
IcircN+b2pLl9Enh+oLa1mQCf3/rucC3TvaUEyQ54BJsPZLqPrpE8kdj/rf1lmwt
hTntwsof/WjTOmKq8pt+puDbwsMH/svAWSTMabhS77Jwo/rR4sj1EkwreHlW14JL
VyEglc7vTIpFBzvyhUPoColhFALUHv14vU9kNNVosKDYXZMm4HCA2qaywTVCfK8Y
ML1pLdNz2np+0AWI9ACBgucQm9bSwUDt+mYJ9wfq/JRU9OsUoTDcQHDrxIig/5/T
oifX1pgwhZtjINKpH8VnQ8D9KZiCtHtF+J35x2wDMxvjFXh0l6+NQ/FSQGKvku/b
8vYF8DFnT86M8d5OqAeWAsYjC15wj+c252YuUdnxMgQVZEc2gVNWhCF6cct7irWB
j+puOoJPmC1YDgE9BNLpIVyQoTzh1/c58Nyx9x67ezODsh4HUNjtwVwoSp6M8O9/
Gu5EqrawNFWj+Z5z6EGVpSnU9H8KPFIYVm1whMGgcAD2oo23B5l9o22Vv0IFc0bx
hbhaHhdsyXyabWptK2deeA9MkiL3u2XhktNAm2nVhJy1MEEBYUreBppHdt/BYcY8
pWr1FfU0+XYI4XEUB9e1Mg2ndsz+Bi7zW4xAkJPwB35WpcvYqSnvcd+Zf/EMsI9u
V74m9MgPMlxRrT8+GgvPs6+PdYMxj71UN1gvpVjYBw+8FWq+6WiCzHFKovmpoIuX
lvJvVjjrNfxwIx/UJpDQkclxIlK7aItAe3+48NeetgLosAfsdZOvBKXIFo6SHHfI
wihnKkJjf/QkzAH92pJ6mskHjmWqltyLWOacm6mtCw+pxrFLfmbneoHkUrftw+YW
31Mhcs+mY04dKusGYchAajLxmXsAMhpl4fxBkGqygGfpIT0PqdaAgE46GXfctAlk
YkKPKGF7VVXVd4dAobn0sn1tiXgzi056blPZ/PVcNs928r149nZyq4dRsDLKqTa/
9sTPqqRMi7XUwccF1RPzjhp13nb2bRoKdg9kIWKWCOeeFpeQ7FPOFZe3Jeg4oflt
enywEwLrLQfRMhkIcmzDyBsgJCOp3/olSW6fofTh/QJ3Sptxkid59kMtiWuLSCA/
ttMFdKc133W/OEAdjnbHX92v7/kFdNWUbyx9+yyH945rI6228daB1CUvKW3W26wf
io0gxs7NgxFiQhwjQwPmJLseNwQVjpl2tajFIk614SUHon0PPa89Jec9cCKumOuj
xyax2O7GpDVlVggDQXsR55T6Z5q8+BACgmr9W+60ZkFONnmbpeeElScGmnNnbjIO
RRCMQYeJgnbE7WxZLtWhPWKptkCwZMK3DgY0SbQonU5erbO+yBoMioap+0YLtlJS
kFxMtJTXAURcwbXZcPO/uxLgPzNJfeFZETG4UhwxAXClWFQB/IfTbrKGFpC4tZ2V
2JXA4cKt6FCs76KxkFh6DSAZUmsxMCwAeTEJFYIrAUwhwTLaaS4IdKhcPKOpV/eW
uFPM5XMBkK0vwvJaCJzkacEYazlxid7p4jAiuiWE2CtwlDHsCD79TFS25snKvo7B
KSgNTeoiU7dgjRwNchqK+Xo/CIGkLDhTS5SX65Fqn3tTasmFTz7FKKSgjRvsS2Fk
OjhQNJ8/A/sIhFBYP4ThAd/U4ieLZYT4SDO4AprIcfKBBYDP/FWSKDzl6msTRKKd
Wxq43Y9Pi564oIp4b0M3iO2OQxOcXuMcqKaC4JD5GxmSEV32u2V91hWKPwmT7sCr
Mk+pWQ8AtvMxzpc77hhcmkWpeZ6MphllawRP9a+WpO6KLKXhYEheOYD838icqX0f
6HCziY1hLj+EZdoQ29O410NMKwPluiFRlr6Nu8rcmwFVMhKGojP+WolTYTeUSjky
QPGCN9OcW+ZGNUvV59uvd0Nr6T2XuAsKfreFH5UqFpIFMN4jqSVZdixJSafUWx6x
RB1V/8LOd22XWptHB4mXymdGq9duDPapQs9AL2QH2d98nr8GERGT7YMW3CwU6K/o
8w/Bk/j2HmDQRhp3o4QHhouPIAZo73ciCi1ksy+XM69DFel1z8PEV7acEgu9bboB
twVu3OdUO5sX2EnvmKCR5VHDBVAHrbkLapGVEBZ/WVq1mHG6d9M1E3pCvI83/FPy
UTdgqnjvq8XsbEeBK9hRGq7gPlBCdG/cFm1Bsu9edotIk5AVoAF4Apjy+le/DG8T
N5DzjSIoAUcj8Abi4+lciI+G9JDsp8UbWY1xKBmmpM/mTWcuzN0NrX02ueuf9qwI
+2B/1oQwCOpqeJIXSe3VLA01Z4s3aYfvS51WVM6rokyPKpugy1T28N+AgURJZtun
l+dHZzIW2YAxS8TxUFM48o6eVCYqIVFOP+LxMkNPMilAOIqxhyN8KI22pgSc5mNQ
uwTZH3L1GnGs/HTC3t6Xgdilon34QEfYpMUv1OYptgfwlEdIBnbcbxZruy6toD/y
QoatPQn6Vz4DcbObp4Yom4/YrnImJfBro8X2lHf7Bv4Fj392Ip/0oDLnM85/2O5A
rsVW9XKinheVLo0SuHcxnPGtRuHFowRYIh9ASGoA3qvFAQTq3FWxwhXVgX0MiohA
B/+uhohUdLAveKiSTtsOiZN3Q2ZGdhDnD+29LERaRVsd9HUGWscsaNF566P5Rj8G
cLSsF2f19t/2FaMsmnLrtVTG3CGeGIfgGY3lDKE6s8R++m7w+qyupj3pJ4V3WaVQ
z+TAP/zc1I12FqyklNQsCMIhgh6Of11NseDgz3UG7mP1WLgdR5Q4m1ixle8eeFZa
nj1aFggtDOSxQzBdzNm8B8HycWFKgHPGEZcddEeUOyskSsBTOZL1tK/rUysofjNa
JEjnhx21HkcmPWUW/2fQuuXHdpf6FSSkCVUMvFDj0NgYVDqJIDparhBtJEpRSDac
0E/cg5iqmpcHaJc7fxjCxhLo6NRGgy/aY7ozqJYGlMhzE+Tx0E0M6HVGBysb33t5
mh1pm0x3kxCWlFBDjIlNl7/6Xjfl93TtZJb2znwEtNVStQQcLsgUL6LVGKUrBBH5
sPhAKSrunjnWum8FNHXF0YXuyEGcl5KKxbSZBB17C8E4yeQAffb6/hdiotyMDMlD
RFIvtI1ghfpkTRJ0udPjKZZp1uKBsU3tw9hX+W1MKWuGPPvYHVoZ6uOlifJUNKR0
fktI1tQDOWffDanizkGTupF+JG0i7QkghwtxeEzak67XddczvePmup72tL5CHbmz
q4D5CHYf4istEZ0l85BEnE0+USiWC36YUTiCuV0hfFtxnIE0LKXCq6yJBcTPDdqM
17qAPPTgT2HQ+aMzQPt8geqpw/9YygK/Lx/E4mENxsmVX2K12mPjlAAJzXyvWE0a
GfwcI4K4J2XUJiT2CBAHKaNyeRMn5/H9CUjFpblMHF9iH99E2hXxxDGkzUtv0w8u
1Aaw0J+umvvFCoJCW6H+jRuUZB13j5bX4TjQ79bcTdO/scVS4siQrL1Wy1TwiMXr
ThDYuaQYf+io38K4OwWOBOSOKGx42gpKRCk+eSM9xLEG/8Y6W+BCgVmwzyv7D1PH
ixXqZJrllV9Fm6qDTNhh+lMwpAyTsb3C/z1krbPU7KOtk6G1DL+oUgPStAP6MvZo
WvFda0oPH849i3vrVH2vlqZd5zSg+dCLnt/PROGoOsOsQwGm2o9DeN8T8gIlFYDR
IxT3aJUZ0DC8frYgXPTyVPJRHGmZVvhAmwifUh/oLLYSkMbrsjedMnUbjmuDbawJ
vs0SWOJSBGeJztbueSffNSDNIB7iF/RYPy8hTvHBhAi8wVjl5eevfGCupNWRGMQR
cNuICoAt9K1Zo9d6VxjOE2AQevkbsUdJ0tHb0WIiYknFSCJ0MR6CdErTCJf40P+H
lhA3GMFjmZUwP3ElqrG8h8ANpTG3/yn6V6huXxb82dOtZU0b5AzEDJV5RETD2ViV
oAvwUQJh31uO632cmcgnzka4KyJoesJ4cK9SKsJMKI0kHJJOniquXwxOM+eULKjS
/TnC+ambOusoAdx64q8ajGUPZmq0MW0V4uf4lqyzTQ74rhxPQHTqFsvddoEjhFmW
cNwbZXcHbCxr+uRDGNg32jzeoKQZEc0nJ6iYXCMWuLQ4UqyVpeDxpNgodtx4Tshl
djPi/fd3rHB8p2LhM5PxtirDiW+yA89xaJ7o6LCU1lUhF69s9lKhwxekW5S5FpnT
i7w/qi5/RdiE2EimL+el61Smp+CH7GCu32EwWLhaGO1FDQms9BgTYqchJ3M5GetK
CRkFfAlapze67Ln4BedRvPeFONsSY1bw2JxbfkOQMhcjdMcPE3BnSAKmHXCHD73v
8P/APNjcFgGVeg6Yztz9mXci1jjbuzROi0Awu5Y9q/+C2QjaG+x+tPhPrFOdpvKu
GGxKDTLvPqsaWCKCZFseVUlAnQqs9b8R81T/IErV7CYuJDjFTHQGf+fmpIBWYbeM
yh6UQ9yqBQuMQFahcIxRDZ22WyiTuh8VCp9BkRFRLpOxWP8L6a++x9TUOPPQgOhT
/Y2pZ9Nq04n8W9mei7HX/QE7HUVSFUPj+EADEQJR3/ohAztBBou+6w9JTKDU75lh
RNfXnW+u2vNGPFYOSSPP1nSQBfIfQ9BFChbj9ugD3IjpTfdJmzdJDBbSjBC7j0fQ
3uQ2LKygp5RFo2V1NY7pt8+nJJ8ZWylAfgvJVejgE8xJzdPjzCwf9OycljPSoX6H
QWMy57f/PW0rjdlYqxx0Lvp4w8rao72O0Kzaq4Q+KykzrMIYcXykOU++MZzhrRO1
j7PDvj+k2tT/Vn1to5NlrwzWv6fGKOs203YVJDgQ71anFTj4ZC0iHUtsv8zqiPEk
WgKMUU3m3d2033UvSHsOlInXQzkIEKRscMsOY17G1bswiVHxe2GM8lOo2mSL7yay
0aKX0S8XD8Cv2X+Mxjkvok9I+uj50F9KNgX+EXtRJZ2hV4oQtGbKKFB6QnHECi4L
eXcj180KuesKUlBOlTsC06PNU4hlwMgzPeMVFziY+t2tqxe3ttKWxTVwKh/UCYaS
aiJMSXDCToZWEUhuClqGN8iKajmfaEyyzf5wVo0jAqtGSnH1AY1/uTu0pip4RF/A
4//8hGSdIjFd6JP6yX7iIVkcppN7HrF7OFE0QK8vL/gZ+cuaCbu9CM4Dd9HH+LAb
ElcvAxNjQ6qzk6VjwMimUY7y3HQmHggQOKii2O1kpeXf9kluviZz/hY3b544d2O0
T93Z2McE/ShQq8jQ7nX3tZMfmO4lp0XnCU0rBzUKU+49R2qZakz27AYff55vyuLy
0ltt1ae4TP+uouNMBC0QWmqEIFDImRuiJtdNgbrXkGC5pJUwjW8eGuw8ze1sg2Jp
cC/PxIJ47JBskMTk4CmaCZugFQcKUBkoOA0At7P0lgVsREZfFXIwh8HSN1ZXOmuQ
dy7Y9ziD5/wz5akGlhfrBG3ui0U4k3p3Zzr2J4SnAuxy6cpJeeKp+VY7v1gexAGV
L0+OI8OzwbWdBX4AeGc1abawktanLgeiV76wJpuu9fXC1YfbpXpWeUXiZtgYnmxy
acNZoCKiGvF+9681hLUQSRHtrYZyMKw6xDUh2/7GUp07Ji8VuF8DFqoNwro4uW1U
vd37M+e0CtA6P8BEX0k4DNhrV0jhvQvXOL9f/lTuR9JBPVSuwzVFN2HVhkNC2vyP
ZV/o11n9bsiLNXfl+7jLZLkat2S97EojgRxLbu/2pYgQpVNRA2QEDLugvjAgBgyD
Z+iCy0Xv2wm+z37pIYDOBW7sMalv7Uh7inztbL/bLgdIKocLMjnJv0Hrr0QeSgN7
1CsFSbCdJAOjEk+dxq1cnu2TdZjY3WFBcZCQAw77gaysB1fM0bOda5xsdGoIEh2o
p2tCEwLP/SJV8MAk3xXp5Fk2H7yP9KlSB7v7oOLocpeMsu9sYF5/JUqObFx8G5VU
Q+8oFulLEHCFa1S/SHqWYJMFHhZvunLKtgaaEIvNYZEcA27mLfR/Lcloq50nfArA
ZjpIZ16YvRO9xH7vZJ5ZnzeBOVyixvcza4kmCrHHlIbifmSreqmiFStlGrVrUMtN
ixEWIDo6TvGuaSh0v0DpNSRUrGaNgcK6QechFZxuAGLNHKGpuWRfmIpsTb71YfbK
aFXeOY9l14eitOVWL7KSDle5YsR8zzowpHNIfRYPV/T1rLT7z1xss12vnUFeIh9h
LTJv2p2/+pxbUhGl+mWH2oayKwFFi0L6XKD+DFVhSmtaY9+uuKohE3A23wDqsI7v
Xe/M7rLiOqvVd5Yh1ScJffYqRTI7KsY5YrPQSTn+EJVN5F18LM6+48bhanzstqGs
dw2+u36uWIT+LMPhVjgMbI+5vK8p0FVAMv3usEv4hKjRYBLOFR2o6EvlLdt9Wknj
b/tresOoZEsPlT6+u7zr/E5OPNDSc6cABawBPHJ/GLu4Yr1Uq15gnOYlRMfJKhW2
4+/FKW7O1u84Kllt6Wmi9OJdNmeBifCblKqMSO+WK4iXtxO52d32Bj/JGgBsoaol
K4tjbjc24qnFuqAfA+7lnq/6LmC5WhRPttXUXslGzgvIw5JsjmTIFXH4Et5SVjGN
szQ+gx7UDtAMaoM5Ce6c6CT7I4l2wM4bR4WfTq+rRcArNT0Wcqa0XG+GrNXpi4zk
yQPaKHS36RraWvpGjsOuWCkKIFtuRWZ0gQj85VQ5s/2FvW0DAFXw3hJQA+T8UzZI
j4NyZJFtpKoOd8Gt9M4Oqmr6TbFh9yJZ0qV75AlwCdSV88Uk3gnWocaw2g7SkTFq
kzEUGtQ7PkgZZQCU4kAhKntT4KiezZW3puhPKA+qg8brTNoc5IZmpen1iKCmBIpz
fTJezLtA+Q9aKRp93N3ALWk1oUOlHR7MmL4k8zEiOph6GJb7uQXcJvempEgLYIqr
tRsUiOzB+iFRlNPyyjmvSXpACF1ZrIkBy69I3dOeSuilJZ7gqrDSvaTMzwxHtgyI
Zfh5p1RROE+t4W2JYi64T2ORIBT84JYgkaAMFs3xZnwVx8wlsRgPfCAFFLcHAp3U
hgKVi6iBJoQ44tCphflIhMxekd55us5qDbGU7AIm/MzlkOYwFCFR2f678Brbazlu
h3S/ty63VBx4P2Y/syAolFxB1xsPdZyhVm8snby/VGvgbXu1q+JP4BoDpYtu25lD
lKragm3EVQlhsUetsRXmcG0YLl1zSEIJiK9pnkcCTXDcCXC+wvtI95WQzlruHD8J
haWedd0XcWn+ZwdEkgrfIQPE1kriqWeKPhIWDZ4OEiyZ3efD0ch83pOWljAKFS5S
NdkCbO/Dh0mzkymc8GTaokvs4gAzgKwmBFIH85mMIuQ8yBkYYw19IxAJiT7qndlJ
eKCcj1wEIibjxInsSe1HNjDU+LuNJ+YjcG2VQCG+Jm96EdWoPwkwLX3l6N0z73Lk
cEnVo1r8ikT9+3N4nq9BpEx7KEJ3j+CgiX3Piq1PK1wYYM23leee4CxIyCwIkfkJ
OvZdPWjq+BTMl82STYXx7zj3/QJSEoCmcxIFQxT/6qPcU9D59fPeznkQvqFPAygD
Ks+deANsVVTP+uCfc/M1ueqN0p1NtUb81Mpk9gAJvWlIWdnIyyKcTAjO7SBFg0Hu
xhhugaxVevXwK5qZpSKl4kLqmjM8J2gLBjTu/V51q+IUGCHbk53nxLIvSFuZlI0E
dtcfdOBzCQy+2KPFTT/4Zd1Phv3gMa35r1gpqsRX0GLM3RB+mzRtHGCmU/7Ln3x+
H2HZ4qQUhfdJ5NEbDka4ei5H+z/XbiE4nGSUq5C+Caq6uDgBkfDF55ioKjmZs2tM
0ilBPXetrihmqxK4SUgHeg3JQ9k3I82fvn/G/ZWdrlz/CeYLAv0ATXbi10rWB0L/
qlD7CX8tQobNbI2aEDHwDOfJX4eT1bpHG720K3RVvOImvP/qkzR749Jc94W5y3zy
IKNRMBL0bSURALPsIVfNJhiguWWEQNhdbGB+D22TtLDYVPuMOQRp6wrdr+uSptJj
xcRzWMiDxaVcS9NEC5Au9E6kIYi9ri1fN/fW3NVQ7leunuYu+9s80m7hXrOug8p4
9zNfnAG8GHAQ+wN5GxnjRHZUO0WISMzy0DCCdU+pyeAtqAFootkxykkKvgPpxf5e
Bn1gDhGI4hq5oKsUyLT6vfe+ZEBs17Fu0J71KC1DRCjDwJwbu8RYDlr1Bv0bKlK5
NXgSqx0iZUvDfGUKyGmBkzSELl8n4AA6XlpMpo9QczmTEyjOvvVWbvtcxwxAGrP7
h6gJ3vMAeumvGpeC6E2T/fem1Tx1v2S5N+yqwMBUq8MYx/Ma4gYL8GcdHVNEOxhI
7Iu1ME7jf5YQdYmIGdTiQB1zCDjyXWSNu2SFCkC8Q3wrnmieJDHmrTQGV3VxwHvA
EAQdSsPktruWpAH2wOsp0sOvZ5rHuVxQngziOqgL0ZkDsDv1d62g4FGLArULw7oP
NPurt3w7o53Kp5vF97NmetgdGrdda2GcZbVm9rXBHWdTh/d+SccIfDnOcbsryT27
78R5Zpl0UbXGYVTULjTVzJdTMPQcCbHR+FrQfWONN6DM8GxdqyOQd8IVMiUnOKjA
HqHJ/sSzMs/YCTQVmTmZL4ohQTcABD1TKE3RXzslcNqom9eUugHuUotNZIWQ2Ug+
/N0Edg47MsxOS9UmZ8OovHdicEt+d6nbRVuY1yOASl2mXOPCmDDaS2pe7tIvBIN3
NDLIxOWIR8Kr8zvuw0HbMJ6GxlvgVC/3Ah/Xj9h8l7n64ZKyNad3MUa3nR6q8EWO
78Em10LEZA03S1uAFZVIHp3FlDoLX9TMuKNOs+odbHuODlmYOXdLV/y0hiS/M7oZ
sKVyAOrqs7hsoHPsY4Keq3aUS7QCcpSbgycw0llUZQBs1faK7qIKmRU276kcyEuo
3aOYEqFeuQ+F350e09RPSZgtl0bJzTtyflpVbAzhOEBcwi4nNzjfoY+4N7LUeElP
SOBwU59+dSuk8vtOFwViJXMlcO2t96XZG5zbbQiYipWazNnw0TqfpNt2Hpn1AdqO
/OWRUe2CpYQku5WZK8tQuSBCC56iAqw/qfZYi2PDI2O15phwgtw2ztPr20RXrMkY
SbtJWPz/ueaW5JkLN5g6K6uknRBszx1veif0m5ZSDu8vHXZZV0k6s1m/hUczhi8r
M9C1BryIOqmqPLi5Kgl3a43EZwk96osdXdC7qHVlr0h6ZW1AehZLYa+v6myX7VD+
lHxZllQIVvImwSiNW//5e8IPVX2AdSQBArqKpRkexIK/IHWdmyYHbOfTDvWDlFoa
V4FMXGQ87nkDpDn2FTvwUBzUO2mHNtfqd2WTCNpeEfFdYhET2MWYznTNXJpxR9fI
Yy92T9c85LaGmeNRx6vm+rkc0olfPrsLqnskTfkvqSJ7yMxd3Y3dyv4L3yrzBzCo
eNIF2mv0GYnjdejvxkViHy6jzgiqrId7FDFlek5kr0HRvqvOvPHlBUW5bLSA0Ldt
DYFO6oLYNCVsHmvG+7JVqWYDtLObAjgw5d1vbtlITZpF0m7vl7iPzqerl0nvc8TN
eP+ytMiSc2dxR4/RbkY+xLHFWNO+RI++KzFxXl5LN/hYbNLxPtUXTfrD8p5LvCGE
XDYXODiOcYUaDduKNUUd2n72VPkOAXkhbIFLTeb5zR9PDxzdX9k+K+ldyaHwDh94
n607VhcEfB4TLe5U24UfRsiIIAOwGpSM97B2T5+lCAjDnOxlvwBM5c8ig3QE7GEs
f3Sc6CX3dszgZZMBUMtdJ+eA+AJlOnMagAXbyKdylgQouAR9Z07S5iztVQ5kw4YL
287NSlHIb0wZGKNUF3H8pY0XzvcUyt6CSBiZc47VnIGHpCcHGKdPq8nUTxIWcg5X
eYSPqs6Nzu5E5Q6SgOrKZzzAAIQN1o0uLHRu8vhD6wQ2CB/+exQ+LsgS/p21BUom
PuTwYupjCCM1Wj6S15L54H7s85evw1QXBFAG+ttK7PaJE2hSUmI0JpnL42sj+n3L
6Tdk3c6JrxYOEVAasZjt0L5AlxXEVM2is187ZiJikY+X0sr9Xi2lCp3lx+PiI/I6
vTu2EDc+kdKtGSdSTLmg4X6I69DGLX7KHC+Da2rTXo4H8TzTMy9B0bDZ7iskdiMD
ePOHX0oSzO8/Pv6Lfj20nAxWZWdXYzdPPm1G4noRrXlvyE1gPe67s6Us6VLnJwUj
SO/bVDj0uEmQloQHbpXowLecw4RCW2E1aq1k8fKnU9WujqJdTHjlEjT6VXE6uMVy
G3ofrwjyyFFm0ddHBhsL3d4o28g8/qZgvgexqv2n6QMcQegAPLL/ViUFOemDf+2R
HYW1ULuL7CLT37KQvcLvMrHs6D1hkjcjIfzkpKJ7oLa6rYYjvZazuXOJDWVOJoCJ
6qDxNKwBtu+Ve5aVR8E9gvZzKXD2GjF/oAcs2aGk9gZ1H/yqqHJycHbKfYZLx757
smfFp3oXfPr0HhVUAlfrX/dwklB4UvUxb5V0l4chPD8wuz9pcakTySYYB2tT7yq2
ctV/JDD0G/V7vrULZpuIBZ9rfUtibZMrLZ4705MWnSZ7fGERPDvU+dRVpwP6Hqt7
JXNt9l6IcPdNuXer9qsuWmFGsH+lkTz2OJOOtqTcVEm8cdlNNmesMWjGu4vySuxz
8KrMhXF0FIw9RImKjLUlWnNBWSDowErcEd8UBCut8xoBziz3b4Mjmn7fCehJU2do
jXj5qTi1OYRWVH2WYGNH8E8SeI6T7FLCZ8m07sWkhhajn+28rHJKUVb8dBPkwVJo
jb3pEaL8aFiYg7pjUonfBmGU3aXbnT2IsLMCFogybPd1ibEDkjlWTZvQgf0blZ6M
wc+TjJH4NXB3J4bBtqBTPrgCyOoEStncECAnfR3QTdAGbPmm6dNN47QmrJJlAtVM
RQIDd/9tLVQk4LKzcxi1ZqjJGmqbBUmaPab7U0Li5a+QR2bxLt66uNboLhy8J5Dl
72K82UmAORx3C1YAm7Cfl/EW8WYd263Qto2dfnNoa7Cj3n/7sQbd9f33e1tqiWh0
JWVL+2lnPBUEzFjXFkiNBAHiEupvBXU7bU60sC8Bw1jmP8g2beMhgpN6Xb/7lemk
9yka2TGfjQDdLlVZuEmwGAH8rQ+YN5i7wPtCvu6aKn8qT1tccSb/hBPrn8m7UQdK
nA61i43+4vHmyjSRHJlmJ11tXj7VeYic56gTB2m4PyUe8gZCBxm0xSzOlSRoQVf2
cfKnoMEjeRCdEh1N5HilwqGzrHukn8bAkwBLwb0LeNHTOpLHOgCBNFZGAZogf8yN
VxlNVsy+2ZFTbQPDCiNfKPXreWEpNU6eEz2XyMwdFWIDIVGMzsWFFbXHy1iZTwcz
wy66FffkeZjwW3gthfQ9nOiAXVV5hT28xYmo9pSRPmXXUf/YlJL6/BI6AnonkO3Y
ZFenBo+h4YRzPKaEN3+789KzsfpTlxHY1mcu4cthXRy0O8QZKbYQlCFK5xRXjSS+
Xu07CCepYETKEJuTqTgDOhDyur/Jze6BVvj+g7SwRhH4finLf0IEKrKsgYytYvc8
QdL9ePpReF1D1THnjQdS9YTks6YrDXCJ1Cp3Oj1S/pCuga2GtbLHipDNtceHn1vm
ewlSm7unI4EziLxDPfFd2EwnN9usUL3gceVUv7MDTbnePeM/x4EXV5r693k6wxnx
z7560orB7nO7WZ4ASn8D5QTbJokhdbEUFSqDd3o4xYdCPd1JOfh7fGdPEW4iB1s1
n9sIkmDZLEx1q3UjvFL2Sr6WRrxa6vjcREboEMAibViC4/qsYnmEsqyZXxjRuMid
cLEqAsL0WACb9HlSgSZCadi39xLer9r15Ae0HLQkHuL0eTd76m12ovJdom4MYmYp
1vhKJhUWT7nnCyGX5isRGpEw5YWxUgZd5g1iZUHpa7iWKeV/Du4x2XCESDPiGSqz
tmmjadRTL6H/Ir/qRqgzNQ+Hunxw922GyO/vJ7iDLJRGZ++efmZ/IV3AqwWju8iF
HKj4k0sjVch+hk5+xVo4EOdKOo4XDGaJLnkxsjVIk+Wwl98c0Lla2vNLYFr1tBLX
gBu7bT1/WP/uv/g64rjneu9ClvFUBvS/12Wjo+1GXEe/3r22Kq3LnNQ6SV3PlMVV
GxXEmMkDk1ybpxg8kiHKsIOm43RaH4wrQzLXfJN43kdlv5NZA0Oa4UzSOroaJoth
ifjf1/w7Tk/poLxWC4IAjqZw6el/AtocBB+2IoVQtEuITvbS2GzXLMbhGXqy9wx6
7Ryi9USonqhXVTkRfnjKv2Dp1HqQLehX0hN5hqVJ5IECRMnfhAw7sx1ou/82oB8s
8/SSqoAigAB+e9Z17WVedyk9nGZNC+2cwM6AtoaALr9ZvmyLwX7N0rT/aSNIhutY
hlaGqhwHBB4EU4yX7y3mKFTrZdfGdhKBUAj20GrcCZFMdgEDkWKBvAvP/DYpwxyC
AwP3vnV5JKZSuOzgj0fhyxgKHxOtbC115m2rinK5V8lrriby8UimgioZloBLhbay
HyIKlabTXFO51OD6sE7xX7YLeLVXE+CMvbCwpLAieLAJwWYDzrRefOJfUa0HY0ff
6X/570YKt6bhS3jplmXZf0qAggemaQ6/MhNu7aQgkZWKCur+nj+wqMkXQnH3dK7o
uoiX9WifQzkL1JU7pdj6nWZmTdQSns9b5IWyo7Dunte/eZE6rqh63UItry4vp3Z/
c8gb0nKQrabpz83gt371hDviT2gXLy3OD3lgtgexb8Pka6eBVesqBKHJVAHJ0yKj
TtVR2aqpKm6O6TwOqHyKvl53AUarzjgDnqvO+CB2vx28hDgC2HJKj5zzW6E0Us57
cwKp77A45d83iMHBtkfApCxvgwPtS6yfERROeD0w14bLs9HL83i/dmK5OSVi2uVU
fnKKaMzjYJ+UmCrPD9a6KDTzjZbKVoqiNpg/9celHBiJ30x/S/FgDYofnEssqFgh
KInolRPDylNH6Ecn/FC6uw6oAKZYq2HFivi91oq7+zlet3uw4qloC0jTLDaAd28Z
XW2Z2eIjaSaqoQr5awLbkJmR/B3gMQqG1mSnzTvxyKJ+tHFsluofykcZ1/8p0VrG
tqGNWQ5JmP6UWmsW+M2XSzULGY3YR53kLxxgs22b036qDfYJd/M3PRmvB37Kt7DS
Hz0nhRyU23Fcx/DCB3ZZr52Q6mWlO2Mv5fPwMenLNeg36Ln/JiMp8AV5tNdI5dBX
E1usMSwOIEYD3Qwv0JO8fFCtE9af3C4sT4RuM5kwMjR6XON0tfsUvyEOa2asnCBv
eTOWcBevScbKbcLCeMZCpc/aDr5m9C8eduJ0XHbznYwZoszUDRigtAd6uXY+JrTY
ow+ZdR3AjPOENwmk/QuT1tJ4H12W/xDrP1tL6W9LingmVS4r5nZGN03W/v5c9RYg
dsLYe1iff717Aoz/u415x7hcHOS0/X9mRoZKkEdPEiDd7h6lX5lPH8MKgRFmaWeT
9UdTMLaQzozDSfftHgnVyeaYgNQmbF/e/CcMDLGQuEt1ldwlpjjQYeScdsMxvGrx
faYLqii8592Squg4tQu0Lw9ql4jpt+UNMvtq1+SVig+sRnxRuE/OFMyyBj0H+EdJ
7M9YySVTvRVOwnfvvSUUHK5jr8enJaEUepcAXPHZ+nQFrprbazwh5fqkfp1zLFk0
9LjN+muMBwj9Fftn1pBuIdkB6WDC5lSOU/BHHpWq18ja+oDz0eriRX0/LpQkDL6O
lGMz0OFdqW/TbB1E4ArtOZtKx7PVGYh/TpqlOrl48bkrfY3VQrQ/D0GSOCKkI9Ty
o//dUJcaYeixS40iGzT6us9Ogg9+0f+gZ3EwlWN6w8zabqNb1IRNnKT00ElVrKyI
hOt279Nn5WR8WYcvCI1vSQUlrzzF51Z+qiPt3PX1ibmNs71Ha0AZekTsHbHnTV7M
A+ZgqANvpZFXN0mS7UzRKhEJBAYe8ysAIDL8mVgGnC6jJuwkALoxuDW0Qs9rdTj4
kEH4zNqNOwKhPlz3cnmzA2+6xROhK2Ra+rgDHk+xCF8JYdhQ2t/L1g0dBgcVRGdH
XO3rA+DoJU/ghhzOcadzUgg2Ee3jBGZPPhHwFS97MxsNJtxK2AMrof7S8TMlMr2B
sXcb9ksQpoCGTXYTtq0vjFSsniYmZXno27cMq4XQPiGSmdkzE8iagJAcZeX7JJcw
RzLLl+9od8xd7ulF0oUDq/p1hrRxLdsPiwX2b/UP86PbS8NiugfS28PMJvmqtwwS
ykf5btUlSUXkx8LlUTtRUpUmNVRUekCBH1bsWoOtVp9XvqDvWVTmfJF4jz8hTomf
HMXNS7VloYSqTsyGViH9AMOTdGQAaxJ4bwwzG9RC+f6XMo9hYZo+UaFkMCq/sqzO
VMlMuf/2rvelcgp7+Annq7pXJeygaLryxtmVbB0abPrUOfPRLt9NPzIneqfkRxhl
FtRvRdB5P7mc6vycmPShm+HZ2p1Xy4o81IpLwaCDXUe5vaD0VZVwqJFExjYyIt5e
4eSfe+ikQFrtQXuvRzAH19txXOIfsp+uKE6yj9BVIADxX7hSzvTcCLl78viEWHDz
CdAZA7ebIAU8YJ/aUoOd8FSag13/9xXp8dF6x0JQfrbwo4EhGAW5CsGDQAMDcm56
6xpjsNkFEROw0AN2zluQaWVBIyA89aHFmyozFx2yICxQ0E6TiGoRBe18nzEb4dUv
Y1VlrrZhqTGlmeR6TFdffM43LiuGe9iUTZv5pilXxYzOzETsh9ueIEB9SrsZFBYP
x9+AGSFmkMwJPIy0CMgB46Wt0s8TKMe73QXUdQscQl9DH9TQqqkFpIeNcyZG3Ee1
850XC6+lgQQopQ2YolFSo+flBuWptyokrLfRAZzJDcUpJLlju6YlOvQ+FiGL8lHW
Fkqy34ho+jl5CXk7iPV+V5O7OT2hGHmTcSoG+P1lkrjslKg8rCy/Kfxv2B8V0w8v
2JzEqSNQPss6T68FuA2CdSlJhZIc4JJZrPePx2mi2nAoMxpVG2uRjh237HmM2uV9
CFBvdrncgitf0hsH3HQcRHa0ouh3bqG0fJegmbCEEdUMSR5/64rKAYx7yTt3aV6A
LjLD7hNR0n+WAuU7Y4K0+LCRxpwnPvkOVhMTOB7prtzudxp4jxKvyvlemhA1Avbt
TjT5+IHjXhof8ymxCpJ3znsZP5QvNAjAypOdQBFQf94IF1GY2DxaJESV70oC+3J3
Q3yivdfyfFO6kvNfKDDshWlSkpr05lz7quKd0Cg5KSMs2rDyKmyMgGPy7dVv5yfR
0WxCSdiAoNE8W5WQbfNNM/87Ye7OE2/kqAj7MFKRH8fDqueskewX6G3oEF38I/pf
8QlConLcz4yEoEoeSHJFhiZ6Vi8ss/ijQwJpJMXUc2jXw1hi5t7/n132z3nXI5Je
EjTZNoD62yQtw1fQ8a9F0m2Xjar9//jaYl7brNi56QMwJHdUdgbEgCsqnJBq984w
iBu1+Sm3W7K+x062H/fOVfZOPkFmRwal+Lse3aPQGDR7ZV1j/MKDAxrUd32tj1+6
cDJrrTaaZCC0K4NVQsEuaN/S+POWxppDBOVZm3iscsDFA7/7nvGEL5ugtBeGNAvN
Is96TPvCFut8Oj8oRW8+wPASvHKL4ss2TDbPI4MEc15K4YooWHiB+HSoFTRBl316
4wQRsAc5bnYuzxyrc4y8tDmzABM+lzkIvkkFlyBJOBs8smMh1BNRHrMrJzqsReJ2
5P2d85VmEZtw5vKQ1WXzx9WvBtx0MB2VTc5JczDKfk3667YLoZ/jPjOr/faCpkQQ
0D/ZoI5RszoZKNPJoXxpOPQbFeTmbpIwUsRErZRApDmnEt1qQ2eC2hw+YEjQdcBf
Bdq7y1Sw783kozv9lVye6ar173IjphSonI09zFKsOMnFHLibuGmK4lSvnqdU0IDQ
5JjiKlupuJS5MckQWh0XMaEZ0IwSqtRSjlF4UuYaw9wMYUjkUhBHnEEWgqbxpYU2
zmqk0UKy9d734QaXizPozj5r8kT50YRL0WDeDZdsOoLLnXeUKu8roExMve7USa5e
K6SIKHiksrH0zJoOvRvGStHO93wwH1NOBZzkBHIHfsz4hqntAkqmKnDo4q7hLnHV
UaSOOiM8sFUwVI4HbLV4aqW2fXQ4mLRS9b7c9hOsnRZWtDhFNCeNAYHDeY+4D86H
/m/+HPPvbcD8/1jW1xL2yNv4WtAsUSghiQaya9eq4deRgnxZuRnomS103PUDdAUg
GXjc2u9TfoueI79203DiDQpNPyDl69pvuYgpoSl7VCdfuu4QvKoZScbhjcIzsGmu
kDmOyyA/p1SXKmDVgaZlnp+ofULUa0L9xxGzgpJBIX93o5/XSSlEk+BolNd1iAN7
eLVx5eb1B8cvKGOBb0nXrECjeyKdtJ1iNkgNDNJ/EQyS+Ty7ksYVya4mera69ny2
p2PD0+cbo7tcH9sa4caBuyGH2g1zDRu08ubLlFcj0h/abVOjy1K7sDbNjm2LGg9e
+RxTQk9bscsYPH3leMnc4LFyX/ueWUpB8kYiwFt2a+NTd9eqGUdGCEHTkt1GiM61
9GvCBQHqCmHaf5Jv+fcs/Sqbv5J4hPAC8ws3yZmKb8u+JOsqoqfyXaJRFff06dVQ
nARmwx8XILbx6fSDCrNpX6H+LGQI4lcWI0pbwKmOkhQfYpsG26cdMb0vm/NmoV5P
zDPNj8Tmr16fY9vkrhxU85wsdR2TdZenLmLDWiEOn/hdE0yzdTtuO5Gp4Nr6zusv
H/8AIG8Ie4Fm75OAqIOrg7R7L34jIuVBrOviY6ZwbFWc9QTmbkMXnbAhFOgxnEC5
vpRSGDuwZ5TARl1iXqUX6n9rSJBAHYQ9WhJv29fA9GD0jBfbbWEWIMAhhe5pNihv
z3cbvC7qRyaURXZ5kzD8LollstPygxkGdeL9Qf9GOSGkgfz2TV7W5mCzrfHEELyL
J86iIrHOal/pS9UHOQM1Xcg1K1NRsUGznwIMVZvGnNj/y690/mFwhPxRZ00nhAIN
BROF6hMb3YBrPNYZ6VaqBuUSkNuGqCQfRqejACwn9NgTVD+xMSy2rs/gwga2rLP/
9jtSFz8yzmPy9n+Gmh453D/T+fM91I1Rz2xs49e9UMiLPNQaQ/j76CDJPwGcYWPX
vfIIDlyhw3FlKf7VwGsbNstr39us+cftLXCpgLRB8G0nodJk59CCQBqjx7qg6Bqd
xS4YoVNKXqdf7ZTP97qJHSoy0LV8y9K7p3LiebkOUsj5Rp9MWlG+I4B9pLlvN4cj
SSVtosnjFrhWIFge5c35gCdI89Jwp9IHs5W2xzBtZ1lV1rVAsg7Zw7+evw/ZAq2a
Fh/ayW5jskrmZVHHNeNfXeYjHEL3wC4O8BS2/jg9GXV8+i1cggUmwh7ifeOiWkZ7
J6Coq2PI+1qRu/j9tdnvOxHui01UYFiLq6MyMeOClBiWnKdKsDL1DbNuqN/cxtQ/
Kv+V+LvzeoqZ78YtXrTH904mFB1vHT0Xthp1ATiE3M5jjI3nQ6Cy0MaXCf850qtH
G4KIchDDfxKGamztyrbDUyiUGmwoSQCcZcTENBlKv2gZ5qYa6vXztHa1pVWqjd7V
28G/GHo68MyfqsSaZvxq92ojGncF84RGfvELI12jUV/1pvDIQabk7l1+gjoMoJbp
a/zcFOYz60hmmvnfbzu80j7gZz8u0H2NvrlH+RSxNYGG1XXUppddt0hxJsy6YGua
ziwQCtHqPFr8inj6n9msX1DzZCEz2PCt70yrrs9WV9K4t77qjC5TLJqnd/tB6GBa
h9WsP/RK+5oGsDCmSYOgTU/MOuGeaIIdcW2qhzMc2fLoqaun/EcYuGB9pg+kGm6Z
zuw8yAKuYgf2JFWWb7gJwIbFv13VrDOzZvmbAABxBtLJnidJGyCi9n83jUUnZzu9
dSvmpCNf/5l+uDDpeqP9+EvGcysNbX29N/iKRflkucUxJ5O6ANKdb/dP0tGlOkuW
9jomkHwU13Vg1FAXVXtUIUz87+YuLUgFwbYnoEyOt5xhA0kY3vYQ0+VSQj0hdwy3
HmboeyD98JYEVlFqlZTs9al++jPgPzDLiXc0LAt3wxnWULr9eMR5GbNdL+IGarqO
aKjXqxeN2DLsSxLYACWlHnGDtlrRi7igQiIsYT0B3ywsnpkq1W6a0iGQlKWRmSBn
0zo2kyLib2SGbbjsS9Ae5doBBO0mYkNkhzSZPc4VCYsy1WVPzB8WkhojDRaw3y8Q
sMMHfnF4a7T4byKaGdP/YDP2wAHQV0e3ZUsTngvUiOermzmQp+aiRGx5Ex0e/7ol
WizTm2NwL7QXxuPqTwvzxjMvr2H/gelV8l0iIXvFvH8U2JtsMiUoODy9h500JTj5
5OP9ilfUVpJFy+QlnVopfq1xb5sZ8PSK6+BPR/Hax68J0UyGZLz9gho1PDQWBXjY
9bY19dxrIiwXlUu9biPaBk352GDzK8Sov2jbhMl1IY2C6bnLedd/BwuDcYxZE2Ot
T48cJIFEzjnANqqYM2pnqS4mnO7Beksh/XE9tMjjdb0Q92grGTdsPg56HmpyT6dm
w53OgHzfIKvCKzz195v9ggHn9xPRrH4RQ702Wr97fE8iFfA8q/xoRMF3TH8hPj4g
jgn25UK1SbkJN0WtvlOpLJp9h42/4ecpxCpCCv/YvBSy5/JuKxg6kCf3lZwhiXYV
YSZ6pqfEzLCzlG2Iz6Ebfy2JobJoCG6nEH4TyblWn9ZeLmntpD+MJF4JDfNGf0+U
80Vb16XBiRCnG10u2uQtU9CgJATFssF6FE8f6jS6kKFBbtrM2qJ6WhagbHVkjayP
ESpFW40VogEsnwHzGsFydKniEeMDYh2FfANQsmeYY1lL/RyL+hiU5q8UUPzQ2wLO
uLMz4gO4GRdzU3mxv8Qi4lVmTrx6ffyzPUghJvHMS5Hh/y3jhn+hengWbFVI8F3L
P54tWj8xfUPvrUPS883UWNAPe3JS2Byh5zz9/lsdXMvtOtlFW57JvJ2VvFkE8IkC
WW9Mel61dE+kYwm6+MkK1ddTgATCNvytaCpiHawYpf4cHvKshMtcYrri67qxKyz7
PlABp385X6QcS8Yl2MxdP7oXbHIn2XAaFIlLYnHUsp7lIKABvMwzFbyfzpgHRFGr
Cqd41LSmGFMh9YYW1xQ1DGMB9ZTi86/H5/pcDmrD8zJJ4PwbS4NAZknBisPbF5Xt
awlpn6iXsWR9Bd+Sq0y3qgjYLmz9QMSSdSYn0r7RoOUOtWTchtKHEe+Rv/ElU4OC
IsTH8tW2YNJ2/RfSzLbk9ocTTfeHUtwtRYk60PKncu/Cuh0f/UlK7E93EJ5KBqTK
6zWnfOOcMlN/l8KVYo4XVLLCcrEgSDrP/9qTjuVM8hxQm9X4kal0YT0MjVgFflI0
hgbrtwg6FpnzWFBkZOKCoJoi2gzIaeiNLB5q2SQf7Iffbz1ibzzzxJGQRADf6nRq
H6o/RfXSbXx/Ah8G85yTjeQJqZmnTtrJ3GwhBDoLSPx0279aGke2L+ASzSR8nrCm
U4vu07Mc7QV4RixXpJ63diZvLw9prOEzNFhdXWBYnmba4Nn+ubrfPQDxygIdOUux
xNpw9ygIjc7k2zgOuq+rUcCmd9ESFP9piFpagzo7ZoL7VzZR9WhpHCIDuV/LEW8Q
6x4PX5bz5cXNmsnsUI80BV+/fLPoDytfdJegiXxHuPGKeem/rkGKyOCnAvofiL/q
NVbCQ0E4lcVlofVr+hu1yO6rHX9GCQqNbx8j44LoIg6eGUtbJJmyTep/tLn2lseC
3GnGqS02XqB0zqrefwwxGzrcf9XliBDzkABvVgSHOzCgBx4NrS9s5odJhjb+qhkF
EIb2dFMF19qeIIckbNoG0SM5FGb9GB7CIqzkp+BAxi6xiXon7bgiVfcyXAa5vXa7
tzakf9c9v94mNOHLgFo6FKDQoeLtOCpZs4FW8gHxb9cgC5p4Dn8j27r+WS9hayRd
P9Hfvd9AcS8zPgG07K5Ulq6sc/m04oksFu8XSQgxIW6ixiG30/GQqSr3B4VvI8SV
jXJMvqTZ9k1IsXvq7NAFUZ4qvw+4+u9aI93EORoxRxXC7hNDotUSbxHbuiTv6K6C
ElJyixztn7RPxcKPd3ZXkitDtDFFZ1SpSy4AYzXbj/x63U2gchmHdKEyEVR1WKjt
2icmUWc9MTtT/rL8f/cVmqdar3WNh9tMz6R6TLaIWQKuJzo1r0jyBr56SZ9jV42S
o2PsFZWxie25tnPgZbJ8n1Byerzfeil6wUL07Vkjln8gDwVp9/Oo3k3+xSOQi6qn
mEVD3pliPR6FQoWRziY0QO6+zqJa5CnJL9x9Pxzo4xHK5t59cHd0TZ8fvfqY6LI+
EcQVArCVkp/VBWcnN61m0B0VPvEYnaDILPchusp5v6QcDZ77KNv9gfGwPX5bK/V8
dVMzL5y3nJMa05bBYkBTsweJiCqhlbG2M3Mj1u7Jd5daZGcAhYwtfL7gXHRRkTd/
yh+0hYZXFtSHe9T6NPZpIJ13aYC++wk/XQND6uv/NURyG2wjQQRdQ2RCcdiUHRNS
vTLNKD/hglHN8xYHVb2ZXFjZiaaEzhEUEgA1w5mg0S/tQE+fQvG6cOILmAf8vQ00
TCZM86nPfPmerNI6mbLgxptIYlup7H5ZT40k93RenEOUWxzYqHu7knfLMjAo02nE
EBBctSJ/Fk0RhmVwxaZIU5bbhlZsrvzUYO4zNqU95CbPmUrWvxniY40zoz9/Kr6e
Lr37bHT3GNltH8+1z3Ht2w8ZZJv0XWaV+OOexNf0DnP4XfpK4gv9Tuw4njMC8G5B
ZYUzg8GG18bH8ZXfmyR+Q2Xpm9yKHBCAxJ2JixkUUHo3+cEUdEEr7cV6PmKP6ut/
T355ryRVukt8/3HWqHtbJ573qmBR9LZ+aCP8YejvnIYH0cFnEK6iLezRxSlqhtD/
1UfmUnf75uW9YGFb5QQHIuCmvkJe27dHcjl41KkrQxhcsT+dB7KarMBRArC70xrX
HIPDPCTbv8HPFJhaH+rEo+OSKlUZcyTURqeV3sV/PwYw06nKFbrANjcKrmDfRTBc
qE1NX7DwPFWixw/7K3/DskgWQambKJg4piwwmGvtj1qPoXmudk7F4YecRXAwg916
oDNIk55M6R+8YwOyIUeeJGV9m+x5207rTQuek5OgYYpZn+qaAsDT/GRP2LBAsTP5
roDhdxFV/fwOS+2TsP57HADz6oyXn/mi8ovA4BNjYqsH1D3eHCo5po5u9St31rz7
hcbFWbeBAyvKfgxTRRrZT1sBgdSC8ckzKb3jpo3tNfhibrc+YcZ8aHOeN90SG0iZ
xYtsKcGzUCY4VWD5JsIe8VI8NW/6ltybgWWvFQq5T0Qe2oqehWPnR4fC2Y4NQNWI
JphQBx8Yt3YvKTtsOwNZCCp8As/H3A49829SanUcwASqu0NSHPIfGaeu8qgexhqD
ZumP+0FOAbc5IGe+8Dq+g8eusbsDfDCU7mx9wUk49OOwABT9RLwI7Y5F9V8tNpG6
GUWcWY/wgj8C5ObIATiv0lMm7OgcwAbiWSAP1yegPacQeJAJKiSMGg8Tt3uTrq8h
tdrJUDUCUcgrhH4E4kWNjT0kbpWzcXECQycavdGu7b5k4keZcGZP4AOf4Em5hfQS
a8M6BPyAiMMHWt9wc4LBtaUUpwxkwlymzeFWwh9J2LKRfAkLXJ7nwxMVzzt8njfv
w6ooZ6Lc4bMWPnWMy+RBzpdy//keX/lJELZEKZle8ZfJVdXusz6EM9AozvIrSOYt
ll+PqYu/S4cgFKGDzeCCEy9O2JUTdkEAsnzBcYyGT1A4KAj4r9a21NpUdiGv0jCf
3ovLU6GdkdZmfcvsS2asxOxz05kfNk5aOenFUySxMVa49e8gJq5mbLx8xKvczSCy
+GU51A/hCUelUwovjYQ+XWqtZGjzOKQ5jQrn/fbYROsZ4XDiVwpeW83oH8JaZkBU
37KHCl2aj9jWP7WLUgQ3aOYgsbssuN2BSytQWrdmloY7d/4UxL5mkLHFuibc6TEB
nlcPs5KwuYpvHZGdtDg6y5+QaI7ydIGBYJQ2Sv53ppKja5FHpIWM70KGhPwTi0dZ
IHfjP90zVlb8kV6hrvzofsgMF4Q7tr3AL8d2ol0WwOrMWfkqWeEnxsZ/Olj/drLx
3zHXdt6TDTQPaw8jGHsuWSWCpQC2UKyUh9rD/fpaX9UQwASmz8ZH7Vm1tHPrbTR9
RhG6Isl7D+rDlnSeQjdCYJ/zc8UG8Y1ikpUOoLdhrUD+ndcpb1R61bbVP63FSvnx
VKndJGMgLJRxSiOG5BZ9bzqOYY7f50t5Xw/vl5NtYE9E2/HujDf38FCAOBzOui3B
36OpgLD2VX3zyDHsJFnjT2N/Co6r1C35OJss7BE9L5ICfiX/K+bw7nL6CqGjEvBG
u02AggQuDvtm0X3tTaVS+JqeNI+jFhLz8l9jFX2uaPG8lHALXNY65og9+qDxMvV9
NtpU76Nvn4wzlZgMJezKeL0o+jlRa/h0xNNKKIm/3b5DF+4qVyeU7egeh/2eBI+p
aJ8plQGQtz4sxhlg3HQpAB5yMw4C7Os1DWpTPEtPb/s7oA6kHfWH/oER/XilV/Ig
fHZSrdz07JhRTpF8AYUbAZfz4u/pQjxKBakqTM1BX6k4HKc+Yc75sXpp0lvr16qI
QV32nK1zOcxwSadzIFZGdJKROno17kAggWTsF4G4uu7PWLZNtwje7asUtL3xZbYm
1anBHUsI6PGMEd7f9MzAnbJobL12KOGhmCS8/TBEecCfjPww9WRJPW4Nh3BJ9Mib
Y2CCiRP1ZLoUEDQcRDNf/YWfdbMVRbJ1F22agojYIIDGAYlTPDvEzoOQ+0NMvTAF
ifcHdtUTlL1rClW7AmLpglLUQa1iXNI3g1fw5wUsshhSCAeN7G1uETk3EvHOcIAJ
vCuzUCmHC97/0FSPrnE3ptYo6bJ3dYKF30eZkzhpByJjpcUebUrIDXelsooyt/qd
+4YO0gCgQoATCbj9Fhh1xxquxTUPfnZWoPq5EeeyJbxcv14FiY9CwKxc+F5asu4N
0kq/Lau9NSF6XWgDflA6Hzd0mwpjrK12TEu1t5bLdbL730N4v28ZrlE635rdnUKV
rLfMtRN6y4zTD8gdXfNYScnerOs+gr4bDdUnd8efq944dWRUDI3Y3UCNTbPjwXPU
dfvi/Qok7anAwzp3hBiMryhVrrLw6RCRouX4Cq1qZUTmX+Ulb8lWI/qshG/1b5BQ
8XAHe9D/ZFyTR92ykSXFYoB0+KjdVs4DkWLCrid+NuFvP3aPRicRed84/HVXcWnu
/cNVVif0edO6fVb+QkgzJOoLcJqlgE8bsRXA/FkbpAhgi6QGRgAqwXxkdvjhQV7r
qZ7G4UnnCMBJ3gAhSjqMgtHecXrN+DjxalwmDeAdSJyIAeC5U2FW9UU2JEkGtFz0
mqjdNJ8LlWqvlp/BUCgVXpkfLqVUmxLiyY6b/NRz0+zPenj8x3P10Kh5UJywRCRJ
5thhGYDzXmzaQ9k5e3nNTU9ErlndlYg9Z8ItLuLedMR/JmAsAJv0TFFsAgdWISK4
pgMhbyahq7cvGyCRyxWiFfgsOi9gauXkwu47SiRQHu3hkiEAgZtC42AQIGPBghtb
YZUfMvAuvBf9LfyDQVP0e+KvcktEXeG1d2/7DvD7i+xhKS/AgmrLskle8n+TfFlo
ObE+yt0NWFz2zz95pd3kr7Hxg9RiFcP7CNSrx7Xrngkv3/CbWtJU6+oC3UdxBX6P
dpsh8b6mP3ASpjyRE8esqsHJPIkrlqATmdpA5peDrNhTQnpTOvwMSQ4j/pyefNrZ
OWL7se8cuJkH9ljW06mNo9X42PBmtA8d79MG+Sy1qQnODHg95JlLlgde5GiYaOEp
yfWZazZVkHxz+fZ9fclpgN+MOVs/I+W+EmzEILjEEfXz2MN9be3WWKgyEyQOYcAg
cuBipjYCPA4xpKMX8J41UBCRWeDzZm1BY+CfYoV5KiGx47GMEsccz6XEKv7n3FVq
C2gn4fsPQryX0ho/V/BsPY7YG06L3raAj8+bj7BLYx6rqcErL2UzZArnYTqtjc1Y
nA+bdM7LoEKrXVM+fCplL7dQK9et1DWdoVO1imRWfHMfDTlT/U4ChSo35Ch4R3pO
JJeNUKwVkh+kmfpPWas03p4BgGRD5/mZY5n9kLXCGPIZ47+FENkrEfdeRRtNW41t
AmRZ1QhNqJGzYh6LppmtpQslgNQ7kTESCg32ZRb+vtsWBd+MqawH+anSBGo0bDFE
8NOpLP1mpQQCsBPCTZrrjSUPJvKISfr/kyaJFTUVHwTKEX0aBNfVoDrs1QexhxBg
t71LWLss45EvtAYJnpz5Dyx6lMXdWan/Eb8c3IN58dY8BdJvKSgF5mpGeWuCnrAy
+joz7OOJ0JZk1XFTPW1P2C5OGRfqQbOXSUpZJ8XO9t1yTRQRHiYBUe7ijYEAVsaD
/CYdRH3au4zd6gcykHJu0je5Fg7SfgN8pfEAIf5WP2QUaifRDHVSwUlD1QGmuk9l
gGfq/x1P7EwDPuGx31RX1xEI5tAephJRr0I/Xazl7jD7mUutg60oGbOfhYAWSPn4
zYHYNVWeyoQUx299OGPCQfhJmGExiahUFGQHyMQOWChT7HHaRLEbSTdx23wBzE4D
nuQuGZaEBPKVASTbbGxByoHDv+pihER+eDzxJyKdGhBihFGKsKuUwKwCZr1GDcpp
MnPZOR1iErucx9XQncjX/+6n/na3ilfnvQNc5qL34fGMgo0egA7Mdi30bXSi6aEy
/sVydjstuvvfIpOvvgLKL2NDFLEwcBqq9P+ZVYfK1/Ovf64hpfuM8RMEj5s19u9t
KNF0IAEM73Mrhw69jbwb1J0NywIiERJ68ha6Pb+qWs2Hoxt0oWbMJisFpKn45fXy
t6UBJ5XAqi+xwq2tpLPURqSHTeCWghOqGRCS2YkOlomam04rosvyf1vdwzSG9qOe
Mm/lhoCii6CcmTVD2urGGzRIi8QN7m8aBKQXOKVr3++WBTWHTR5UcMeTbw6N2Kng
rMols9XKk1uqOzcsXEwYymO91bVOlR+mUW/P4wPS5Rbj/ws7JN72gp0oKpbtz2+k
Vgi3BZMfZJJxRhcRsool+vV6vDMof9DrD82ZzKrDjkeZvz5Wpp2lVjdzFvZQkHzl
I7w/7DS9gebeUU1sV/ONZ4gasm+nyHsfWFhY0q8oW7xS1p2UHRB9bPTBlj7+aeWz
3qrmnChpWPk6SBLKzIciTmZEumzB/Dt+P519C9fy5l2PTwrlyQkbkSZpsMvrlXiR
lARHHSs2CmzDb0m0oMAvR2yfm37+iK4jjhiqXB7mKdhri2dBlpjGP3P+Z1xgim+D
xPIOeFUHb1j7bIMY87wKHyqTd6/T7mt/J6iBs6pMl5yGpHPSBt+9wCZSURaXXft4
bqZIk/xNPN85FwE2+eosdKagniCDFYzv9Hr7Dt0Qm83lgAlywBVjNeTDpPRDfzuJ
rXfX0bGtePkuf94kmIp3hIxHHFp7Zrybg91Ewxy34t7FRtiOE75olfFsxZNrTeKT
hUvq3Hd+MoXNF2i175INXefHXgNpCc8wMtP5cu2KI2Tghc1fIIAZuSoRnU/GyrvT
6+paS4zK4I/Ln1egCaJT2N1A3nX+/KtO+LXdLv4V38yCz1Y/VdUrXz7IgxI3x/RF
FXT0tslBjiyk7qEx4uSXOUuuuCdSPJwpwT8dF/gBJBNn338yxzgBjrKtQop5TogY
1XIJD71gHf/cQ99ysWT42hOoXBJDNRLE/+bAjZrg5fQ9h61YC0w2eg+Iu+ejWd3A
47aHfgQpreoKVg5k9gw1i/fbUTCvAxkyiLqewaDHBs/i5IloTcHduXpJCIXz++bL
KLF0zUvvhivhvlFB3ATaxkgOu8c3FRCzq7Khb02kxQYtKr384zv92UYAv3ssKo44
Bo99/gQhEGnXT4KpLnfx5NkGqgx49YttUaNAB3KsNq9rw4C6Jsoui+WufXmodDbD
6gcMnvV9EOxFDGINTWemSY6QxeRd1MWTbKKu3ekf4OaDuJLC0AvwySrTp1xD7I1v
xKZbXsuYinKRoUwYN9qSA2F11I9xgZgNkxbcFSmvG6EwWSIB6XGkfFJuX4Ogd9s8
ZJmV1LBOyyBf9o4kvMYJDKOUMVciLEuLx5Xpse0rzmBJqRyAU/QVkxaasMmhrvMk
GcRN5IJDL2x5eeIeYXddVdB2QrEblc+Btrl8QTngpwrjUqxEjJQIHu2vWQRvIfkH
aFS2HmwQQhQQlpOUAKZ5kpyw0T4r75m01UcC5zOpRHqniLuy4TCYeXAkLNVw4uKB
R/7mMDc6RX/J/TWpna243Mbh3rHKky4DD+h8VLbnyFag366SOT/Vh1TKGPITsqKk
6/j6bqir5IXOpQ8/RX4cy6MxRvOfSaoT5d60hHlmcYa/d56JLGWX09eRPDlr9Dd6
JWkHGUiqGqlBk619EQD7g7Qu8qwq6NXFwrqyUnBKR74H7YbzAt+GUytVEzZArSpQ
oZyKxL4SVY2msBl0VrmtDy8F5pU0OOrm4YXSVSquraklgo1IYoE+QKblp+4AT8RR
a75wAzbNRloHnI3AevseovYKXS7iYkzKliGqgsiohbK8Zu0X2VVRvvq2TCn8qvb0
zMyxoggH5MxtZwENuuiz42I04Zp7q/2to7n3F5DtMwt9P1B1ZdqDU4r/WKwC/WaZ
h7pFS6kzhpmOKZGITsJIYpgRr2eUppU3KPKqKuhHTj65tuFIByKL4Ha7tawdwl6J
mSX2tXmfAZXwTk+8T+r1kI1rshRCHZf13ru7zeGYXpp8Ys71LuMn6pmEEO7J5gkZ
fVvrMHNosVMetzOtmBwhxSo4esWUZ/sCFFZKybPZBuysHekvNbZxvSpXTSM1uI/l
goyY/WL1QCt1G8TG767keTi4ziStAGp+L6H8vYD2F+sLj43YClgPtxqtF4QeGW6A
/35vyoCxsOPHcc/RblOxO0qG5XYYAnzxCfiILFVmh9dQ7qrVtq+/ek9CfqCH2yDN
SsvhV7KaLsp2KDfiRbFraaaGh6q/vptFAbhWrRJ7XyEQYq6A02faJ6YckeOGfxK2
Bj3LElSeycJoJO7vtGSThIo9rc7hkBlGBfj1jbntE89z1aCChp3eLPWYV/wSWdLl
VCnd3hgpyCbmUJRa1vFS9SvnxyHqE/40s9kLWCBy7Pl79Qns30P0MBaN7nPntMZs
RvLBN1ty4UGnUyEfBPrBc/t6YGlEBHnms3yd0NygQPTc12Na34k+RtBzpsnSvWbz
FsxiTugq1SgAbq6TJn0otQ4YiF0jv5bq5+nzjq/XD88JSkGAx9ukb9U5EXN9AH89
qV68lMxKLFtBHwlDEdieIeoDHYz+cJM3FFivxwkA9PQHDddSnyt1ngMEe5vCnzak
GaRg3bGHG1E8cR6YV76K5vdSj3+WT86U6DeXxvMYS/FrcryjiyGYtFAxtJZ+nJN4
xXY+vWvRrVbHxYgPUQFYt/lxWG1QgimpYgZXqKk+ZQUHtXH7hi90dey2SM8uGvNq
QcoNsLo01Kx1Vttn41D3hlvUj5cWpO+uyPBHW2IUslDaJuDwRnYbpnx1oI/QqypB
jUfzFXHC6wcjEqHYmmZ/3oIpnCtKNAElQjdOYZhHnZah0Gg84/DiKsNf+AwebMWG
ggxSz6ay6VGVZdUQCUSCN6YuMmq092oHIeAcevo6IHf7nN6TQ1I+mDAACUlzl1c5
kjGz8umD+c1lVVilVdwZ/jAmGmKUGkxEdN+yZaqf45dh992MNBnVBvv2I9iqyjG6
U+r5t+Jt6Mp7nlpKGdD2mSemPMMTrqwnr6FwpfRZoCj1f/W0czK2RKrMwbAjhqpI
iDfYRZaSevxxlIvVDLi/H0+7y4ixAI7pJKZKMMU5H99Bk37gVvGjLkNpsHVcefhs
lay3+ScBCOnJC1US9BDAI13EiBegpImF4A4/fT68xoR25wRer7MfaYsDiYyBgU4a
5U9GxK6SdY8LYc4TWEZbbXTttTKi34YD6+Q7G2T2BLyRoF9BH4Y7fnCLZQGM6aTx
TGfjdB2/26tg8H+J4aCW6JWjo9MJM1eN7vLjSxa1D9jRocyVDea8urgL1ZXQPnCm
vo3qQ53f8d/IcDhaat/r2t6nm2ZJk49E6rl/Nvk+PFvjqR6deL2Bnek2lbBEES6y
7O59PteEHiIRvoMKN6O3P6mThpITeBPBcQsHwQtFoRj5IN8r0r2Y+ch7fzHWf6nG
+lQT/N6HvIisjM/Rvrd2HFaoqi1Y+Z1eX0ZWiZq8DdopQg4Ba+hlOzW3icKdJqMZ
ULRIY7c74Rwy7gpP+IXtqNAHb9iOBOo+olRz3aqaZAlJ166ibnYqUkytPi0o9UYh
+v4gpzQtkRt71nf/CO9v9qtRcH9MpESl2JdVNnZm670wvYu2S9O6T7hNXazTYh5h
JzOFbSLbgCDHg65Mh2hqhqZA3S31j2ld2Z+sIRvMmATd5XA+qanodnGGNDXFPg75
9ku0D694/95xBUGpbXrLAD4LaIp/hgRoHQ8oLlAVeXBnAM9y14eUy87Xo5Bbvr1o
OFStHMPApYbzo32nJwpuw7z50ort1n6DexfMZBjJ39v//Q4YE/euoMHEfeD3poXP
GmM/mIJDLIHLDdTPMjCzUZ2NsT16Ufj8+pHiFZd1OOfsXmLaF/J+rvSBl2TWOBtE
47MRyishY+K/EZkDn+I0u8M0Z7L+5Epdgd/1gIq7cN1y9P5SDCC3cO52jS6g+xs1
TGYNwnzln4kgL463bfBnlBflJhkjqEWDgow4xecWAkZ6WvGW7qWT6Jj7DADcV7cS
D3wbKcCl7WjOMZSJBKTktgxLbM14K1E9+cyv2q39ZmYHu12YvV9QQ4Iraqjz5STL
pxIEv39ui9KyzSHdwVZZnZSZfKvVALBgEKbvr5ykE2GXu5A0RhCW7k+PERUFOctC
pEFQWlmiiLiawLaQO4pvHpxWgVepqBUbhssC2G3JZekYIWCPqax+iODGag2vQlum
RYMlh3XhE/ArHyLl5kpusj178wHN+/uGc0VuvTkaFjMLktGZaMnJ8R8Wm0gBRo70
cQyDYkEbrmYUrfcmfi5mOFheORFev8qQMUtVwOLT06tn5U8BDBttQDyhxiJePPcn
9ckFE51CLr3FsZbEGCBJKqa60YQ8/Rdq51u8ZJfBTR/ifPqXDb+SymB+3/udGsq/
aST8rxMHjw8ZoQajbH/aGM3Yvwbstk8CnVQzmJlgYKiEKJHQQM7yDH6ZlWJl+y1t
p22/MhlYmD0btcHuXW9Ux0EES/d62q6XIfJA/3KQ7VR0RhKex8SbWI9h1Y+IRmm7
zsRDhkVOU72QHHSBk/M7tnIAf823xZm1G6Wx2Nqb8hf5Mf2mTkzPLGtDT1iYUlKL
R8Lk4cvFfE01etq5R1p42TmJXpgVqAxdFcuxBCp/DG9voYi49UMSA5gMXfwa8lei
QpPK8CI8empleY8pkYe90uztuQXzH3L2JYerMf9M4/qLwHrVCRDpUQRBJPgdH3g8
jiPyX8+uOO4+tbGclq1sNyHbA6dQjPRl/7bR8T1eZwlo1oJ73rST81EJ4X+YeuXc
7T/ISK88W0LRc8MPsXH6k9SMh1J/tdUmEFFm7WTydgBGFZQBLIFrRKPZ7DH1Qdya
cuij+ASfV6gFLi+YNw4/F4DI5RLwpVSBo35nOGi+RN2xomJyOrlzIu+gwKXeTBjx
vhOoXNC8KoF8vROKG0ahvy0fLet2wD69+lfxUQ9J49EgjvRpTjkTus5bdNuOdyAG
hl/jGFDDF5IOPgLDTycTSYEcH4qG8Joo8zvW4lP4euogf9oKP0FHhIwTN9D3us7J
sy1QG3mwSZmF5uCLGxgUCweW9/s4PJO+Q3nO6HplCfbvP9LyzwlPfdcsyf0IwNzl
mUYPAZtrGrT0UTBcgB5khUYluxf14LevmUra3qmti+UlvTt5mP5UZENXFMFn2hkE
CdlR4Ntsk3BLNKNZ1SyAilSlnMPA220fYnVWbPBME9fn9HRAQISE1LO3ZN2+o1XD
E41aEYxw4vmBqY/KESbIGmkQhFAgHzhgzdeFM8/V2fIdHp/p3gZTRjB4oCI4FBm7
l6VgjLPrtOG2hUra19VwrOx2DLXXBEGbqqzPYMaTwQuChA1VJkmfk9UhSoQDIVgb
KINHPx6AIjcyxnfUqrEzutrxpUNdmZoU9vym+GxuIPpqYUGldFXPGORwv0g130fn
YNuQYBxN9w1/JTsospONXlysr9fOL1PWIIWRkOKmIA1tOZfSbkLXcc7qxc3JaRAO
kN8m1SXoTkvbTaFtfR7L9GhHiqX1/hbQOtHdQrWfofXdhg2tBAYz8OxsijkxQ/af
h4pDa2JRa4lzqTRCSZpe4NEYpg+WnyKEXS0isQtjO7Cdfycw7PBfWki11eVwzTvc
893tuum5ogMYjdGI0cmkEm3bAngawef+r7BnJvi1Uhziqr/JMoV8ubl9Q37n6UHf
ZBp+m6aimCdfosJsomY+3run+86GA4AvaT+kRDGC7Ur++Aov11dzKzRJ4v7sCh00
bbavcHxYmU5X6MXxKd0iV056NMnSrc4GexHuykIr2tPamVeC5OINgQjgM3tJcNfI
7fLtOQ/6umvwTP5Yl/ajtLUURojSVrIMTVzRtebZIOtSyU3mHflagTADX0bI4M7g
ZOGaC8Ts0JrYHOxfcjpLhU6uqXXDkvE15GTUdGFaNHrx2X1DbTdwneIbvNK0at4j
t9dSyquLH7JBr+WjyZ5moRFzikn+fwa4talsR+JoGg6vElP2OzKPK5WMp6anw1mE
KGRWt0lccAOcPuSAqt3m7SxPFqgeF35v4e86Fu5g2GBhnYdJi/PKGGbzKvTb2pht
OETXvsI+Qc9+3p5lQySdM9lkaPjk4VYRXvuXl24SzrdIRstmcpYmORfeDBC5REnM
cKv7Y4nmIltaxxPbkZqrHJOKliMm3iOIUk9uRP9mJkKfL0rLrVc/6uKSmaQk67/N
rnTDYYW0HUIyyLM7DHXDF7c4BTlxIFKoouPjoaHBLPIiaG/r9nWSyNqpu0qjrleV
pp9pxLuiorYL5M+H3dOOTd3gBmMwBxo2DshBQLPbqEc2sqrZiBxH2rUyf1WC0gpw
dVxkgwf3mHWH7y5nsnSbiJ5kjFxy2hjxqBsfL6VFaFkiscOXBup1A3SsyBt9zd+Y
LHLpiOJWrELaUHhW/oHEetlJ75Qom5R6jZaCMizFjRO0sqMyBaY9wHF1ruUOc7di
//wij/jTBakGWyFAinKr0gVo3RKgQsbpRsngx8ttzaTpn2+UdsHAqTqbIFopAq96
wt/y7wh5G8/kaV5IUfHaLFEnV6nwqFI3g9v62Iw5UOoutqMfhXL/5TzAeneojAuy
/dSLeoWlMEKC9Ie3y0WoqlckYZl7ZXBEf7TFSzyCMHKOzafJLLA62L43dhkQHHDg
mthRDPdw6SCXtHpGoydEnsnDRf+gT6Q5Xo4fM+etbnuYqxrhKT6qAmR42tG5itWB
PQX547YL7Gre2A07vmZdsLrmUAeUoToARXKNOoIdiNbe2z7xaI93Oq5hl32sZXLu
YtYlJ17dhmDMQI+gcWMuw5J3fl1XBM6dI+GjI9f+TRcPUi8S9uvhPVJtBIzOKymG
+HBdUyl/Z66FKwFzFO6VIYnGB6NZRdSOEEW6TICEpqAzxolp8U/yIp9cFjbE1V6C
CYXR5fglnCr9sK1dNfLHWfiqc9bfK/e5+ALFnsrNo3Eqx49VOl7Nreq1GALrFKs+
77WLe4Ex+DQ4d5DGVUfGa4gAceE7fVWGHb7HX2bRzzds2IN5pW2Nu4JJIWMNO9WQ
ovVYB4YmyvOE1dtgSfS7EzW2DFxNdOPGtW5/T7mt1IJJXcygjCP7IttgSZC72j0V
3xkBL5Ik7as6Jg5UFq0tl4i1VnN+c0Q4LjPKrNG52tVWTNKOj/1++iggWgfG6zMz
5KHdwpAXq/tgGwYTHZTAweuLD1nwEf5QyPllXGHY7taS0oBNnJ+mt7uSZalm89Qn
Ns05lJI/ibbtK+xTQ4VVwywNdVV03jQPFTQZhCSklsIVU/Cc6QNh6xOy1ec2JClV
tIZYDvavpmtppmtn2tK034JTvSvSmeeWoJiY3C0b+KOJmUQsr+OoTK6dWIdOYPFL
74hnLoVyFfpFegfpy8Nx/SQZWUJlMqWJIHKgl2Cej8mDo05D2KWjbkU8ZFEWsPI3
3feXuLyFCE1RuxoWeHlxapnhQsjEWzON6tHdjGSR2PM+/8HAViRgyy2dSHXHJhe8
UsTE23ASYNkUSmSs3kuLMILPGieaMEigSVesg6WsVCej2M+LmX6DXWQeE9PafwuM
bF26de0DFMoumpW9vjFCH30Zb2FicG0PWALeRk+RNPVsuzHjudDotLL7IXji2cWP
9EwNDvbtbBZzC0gYalndJP6lrQ8S8KYWLL+waJ4e/mE3htFyYG8/Qut3DEoyc+3G
thy8sibhGhBGl1RUpJV4BUqlR4x7GJvq33LfEhsCMHOxZ3Ttp8CVwyD62aon3rKD
1ntsMWRpz8b7Jd2N5B+y7IzRNlrGm6609DxthTy6/rtsVbjOZu132eGt7z1BGdPU
VTldPp2YCODAQUgTEKZIE0sRrYTTPT9tDdj+bl5tJGFTTOI7QgwwROY2aJ4o0ufz
SKmtHcFtspSUvyYabkI4ZxcEatIbD5d2Lm+n5A9iGP3KohvysMPzNs8sIj/QrnSm
yMWyP1ITN45SAAScUcukUFebPmtl824Is4i9i7x7yfEyVqMByWu1ZcHdtwNBhn+N
scChNtw6vcu1VDJOH4NpMfiCVWot14VKqHLWfWBXGM2OiRPu+qegjr0TMBVwSQK2
WaJEu+CQvjlvTFlG3W+cRYqUbR09SEyM0rEsmjK8/uS4pAhieWfux/DdISvhURF0
+/IEaIh4LM/Ah44z+yfAKaClKTMhETxazv0Rx1IKTVF06T7afZklMVcr29pwXMeO
lU4wvZKDrcO7Ddr16FEpUFHaTIyDxhozw2ZKtmAjj5hrBdKE4EXPk9HZ47PBFJD5
U89qIkfilnUTNGjvnQJHLQlvVhTO4/R0ryAD84H6hucVDL7oxE18+e9qbIu1aXT3
LoUSeMcOnRjCuvZ6oY+jojBq2VG6A4dB8timp0KVVYZNFoa4meS0XAO6IIHQbHu/
9KNOu5SkcANkMBrPc+Odjc3tB2F/+JV90f4DjBG0v3xfzf0ixjjwgHTeZJg+ZlGZ
lP3PvcfRAhZktBXHVveS96MxcAuxpjUrRpcSK/al6zEOV1B7yvaG6KWcPPpwZviT
MyEvVbI3oUih702eSe/WszDgb7/xSoMxplFEaHRpeyppcIfdH5fr0/CIX5/hcqPU
vuWtapU/2UpmKp6DglVzCuAhjuPoYCY2dCAkXLhsfCfmGs6WAUzZcN1iJUK8YSKE
CWDv1LGJws8u0i5Z1317bdopPzD8Rjj7ihmjIVoNlaZw2gdhg9WwfFRNLawB1ve2
k+APh32WULo5FUfK79wKcqapuVILTzrvu+SDvRoID+JzGbTDLD0r0k/abo5CxczO
2lPe/xYOiRR+Cozq+c/6McesN+cnkTAPOVqB2UH2cpN9wnwUlKj5YPVFoJKBD/3z
Gl4omKpZL1Wek+2liw3BfBnRmSkn9D/pej3WrVY7/8RVi97qnQaatCXvJDR4ctSD
yAiMRNSD6/K0wFgpYvoeAReE8wR4rB/j3DcsIVrbd1zFWoO/g43//SJy6WMDE+2T
tV53LfCqFWCtn0o+Z2wAn6FsxuUeabZ42nP86nCE6xGcbAPZC3f1f8GvE2tfCDf/
LabG+dRtC43W2wrKtnm7O6N7Llnnu7F/fI0ZKOCzarGOn3+PNFJHPlC9BZiyFB/K
pwCJWkbZ3rvvcrBX74jZxH+C47C6WZExsyp7D09cTthfdaaOKZSU243IlruNCRjy
gqikg1n0MktbK7ldV4er6G2iAaNTpcSoevSoNSwe7PvXLdLX6RM/xIdbP2uniGvQ
FHDQlGoYeLWFP1xIXkATyE3L0ZGhWoJPjNgNmsVqWr6AcjVHn/hRbz2VjBPjT7Nx
seI3EwCBqAIBGs7lzr9Wk6DsvatgsIR0/UgXaRGLsb5EjIol0KsB1Z3mNFaatOij
dfAJ9Jqxvx67ST1y0f+GFnQ7N8PB/PbeSuoh5YmsBoQWpH84/S9EbMYxmAAZWfOH
2fFETQM0ycD+kB4SJ6UjHetjSwb0WIqudTAQd68qdbBKWIul6IZ3CMttqR6itK77
oz4RmPuaf8HlCu9eD2u4cQanllZefyH7eaiI2GXa8DfG6AvjvjKEzWw06eK8aZoa
CaZhrk0mBqSBI1KFBmBnHzsOluu71fzCco69dY39VILLjtzp732nz4c7xBH1boTl
R8EEolgKu3moYXazCIBck0p7NRH0y41fbIgmWhGlQ3l8/x3odqIrhE4VPBG5fql6
Wr5yUygHxFZflzFCJ7AUJHINfDWZarjzyCo0F7/vyCe8jQNc+DUZZsTr79I2Tyow
soxPQGTmZujiW+cG+rE3feUTmkSqeHZUE/R6BKoCRhsUs8s/NyyucfMwnxjMX7yq
T0f3UXHwSYhxvo1cplL4siyaeUmbhNZ+8bbKMNwCB9Vu6pXHbl6sje2p0dcNBAiw
ycHp4vTyoZ2KUCgCD3Kjhnr/NS2oPOI/X0uR42V+bFhL4iAnsJwEJAPmbSZfVyAa
qNGRbT2v/uN7dHcPpO+TJ3Nb1b5Doipz/eFnjOGXki2hOuDpv/eLNlNVaE0OMHxp
4alenpxIYMCGtu+lGBbjCU3ZHjwXHEbxUQXpxK0JB0tY6DufPQP4ZrNjyg/f1xc9
5dXSwFQyom4g5Qho4wmnOKaUR8LdvKjqRWIz7Y/Egm4cM8r8jm6vplNe/13TLMkb
db421y7T/E6ZIo4LXRjZhxBzz9OJ7vk4RrbJF8591Ygtl4rfgBaiOw0AguKxPZXZ
Z1O+TLhDnJy0z8kDfy7E7DxySl0A0HLg9KOS4DKPYCLI0xVOkaBjNxQTNInlWZCj
SW+dn4oFe/D0J2gVWxacWLi7Q87ZldUxg46dtt2YaJUrRimeIMl+aJW5V8soPNer
6oXu+U00ssnNM6bcqyxrCT3U9sBSFTLmnnONLBzPIKtEuDN5vcrXStEFuGFVVefK
mIp3l0SDtwFiO0sX4nWmRUJuUpAmrV12V2dMi9OwfiBQiJYgr51AO5UvlXRRHYNU
Pdkord6q2JlYft4BrC7Q2wT55yrJY4R2XmTRYz/V+52ER+sOB0gzQSJHj/p8bwUD
mQ/pH8gj2/p3CXdPy2GhXEg4ScqeEKDG2ZDWu2h85azy/0ggAyYhBs7HFGi2bcnD
6RrRSeptcN3ahogp8c/RxaR0cDpMp/yozJIK9oD3eg+3ZA1g1a0CfcgUW1gN87gg
69XmcUx/8yMC/6oY0YJSpyJBs3xw+95TVejUZ6gW0EzC9bY1pHiTSqdPzDbqKQ2L
98lV2+Pg1P3XD1cTpwY+O4V58nvMNMdAB06QCJZeQWERTyKLqhdX82Qjt/7NEjYJ
DMP1Ib8LG/qPFgC5Uo5wbnBwoeAH2m7yMMobNFAigdPeNozFKOReS2Wyr29OLpWx
bymasOgIngr7eaE1En1QydyD0Jovg7xJCcnuaZzbT4YglgSXITVbwmE+s1OIdDtn
7L/8qSCq0ko1LwjdMyEyORdapNHljoOuEn9CJ6aQvuWPWMW30+K0eSWJFMgTfURN
sB7O67Se21Yc3jveFhpwoj+/X2qhWmVwdU1W7dM2s39hcJ1xBX4rLx6kjGOG3UBu
5bxoe6Lvd3PTWZg7UoMIyEVNE5Nlvxfrvxn76vVF1/mjil+cH108Vi3+q7lPpmDQ
nLPCdnYhk91F1YYMykZ2nf3VAbs/Ugl/7MGEGcf+FNLer5+B1jAMEjsdHyq1SntM
ozkKv2sI7ue7N8xGcD4qoxJrUKLvQgtYME7J7V90VRcHzGz4COFlfiBEf4rkBB5F
EHOvMTIjMXmN2VxL427wN33WnSe8Jvtek6X9sBoblxF9KzcyWXzeBR8DmG2sT3MQ
1WfV6ZxC9tzSVBSPIkv45zQn444gk50bl7GCUiTrg+kuQqoIJlJZ47Z6nBtDXTMq
a5LRb/UVuD46yJZCre8g+ifv1Rqan5kuzQ1xBBI0Wrbd77mFcrL8cUPtNda9HBdO
FEvy4rv53AMKawMKBYR61ncgQhR9WmclcZoVtA2/hHjYiaXpfd2mrPwyh6lpE4PI
ujNHVM5fN/980UEdBUHuugGPMnTM9CsJatfCw2yZHEa2dUJhVyBtXdVVP5dEB+2k
AZwNQ+mWVXgI+hmf9LqrAmBTvI4RHtY6Tel/A9etxvpXSJZ3jARCN0n2fErIU0z1
BMEBONDgKN70o0JgPfq6yoTiGGf+/fVueUu4tNPkpCZF9VVivl6GZgwzhJ99Lvr9
aMsLGRufQpYE2GuLreLtgMoAC11LB0foYAfYRuVwQ/1K1I87aM/jxRWklGASc29o
b4+8NG1hVprzEcj7nh/XoBUVxneFAWvdSblUPSv5EmRSRAPia+aH6zzdjqKROcpo
H4jBREUsXmgt1FClrN3U+UmIrh1WYs5INZe9dSB2t7sDxshCUwyrb8+76IMg6GBo
FiFDHFTMejejALapDuhsJwOZI/8WEbtz0jErh8oOKtJVm0oXPEPxM7BQtYILqGiW
ItDvrKjBDsAvCUapSNiygcXwDnWnvWqEFnLjlRWwIqicMSijX00ly8U1uUNgrL/O
y7wuQbZffctM54vcvS8ZbyjOpIxdIUvW1WnoSW2NfvNkMDx7CzgUaSkcYpdH8RlU
lonjTIFn7ISNWjRrPiA/qIZtKU62G5JZgmGrytt3fVy/tzUwzEN6NCHvj3jHXZqG
SsgFrZonzNphCi91Dndmu6sSc2OlLonwpUQwMgKykRIeNdQIE3s8QIgB8dKLU3hi
YmA8b77LIIglLzz2Go+XuqzcktjXLPsA70sZPqmP/Lm1Czv7XEVTJve9NUN3Ydwn
exsYohs9c4pUuieNC/h/+GhAsaU99nLdCyK8gpmMjN6k8aa1SV8U86obcONfVlNZ
Q8FqQptxd9EjGwbopm5Yx81WBKtv2EVh+2DAblCUndvUEt8C893C+78NIlo2yfJi
HKkwrFURY9t6tvveAVXFMopV+v5FC5u/Q+G4P4voFIL6UNLx8Z5J6n/68eavwwEk
BdIJ3SDWxErUYQ1RbBLAo6EyBVljE+bUSuEJ6sa/1TqcyK3OwqYnsiynBMJk057s
TyKrTX9CqW6ObiL73wJiK8wNI8JhAxWcF6V0b0PqBy4SGUnN3WF0Hp/TmRlD13bF
Gyiq6CN/0ON6690mwdnU1ephZyKIy7IGXZeZGfnSOkWdIllEh6zdN+0Z6aZCi0uB
KPxydegBrXA8QlqiBQ19A/+ok2JyCQMbC/HwNj2TYrJusj3NXH4bo7IdZM8idqKC
Hze8fw20uvIK1EB4JYDJt5HnUBI4O905eRoX/Woh5yjPKODQHI1sVIfJT7dFjzH+
cRT/fO0rt44GhgXQabLlXqT/uRCRCh9yS+GXdfM9NIki+PfJvcCOk/XtNnO0Lfoc
ZIF/4pLLjpGc/bY/IDO53l9DUczeLNnS698DuFfH9N12M3HlO5px4eBCHkC82wa8
/8qKXqaPd2t8zUMx44Ys25eIllB9yqEKPN9HT1xyN16ayvrw5Y2bvwUTxJoEbkf4
p0xiLlXyBRqaMy2EOjnJOa3rL/OVvdcMNTuED9qBv1mMKdrbF6WFZzQP67Wbdo1H
oYHA2jvAlIosmOQmaLxl++/LUpO2YY/TaBmzDVZQuIgfbnRG7OQZioCIhzNV65Bi
/OJFBSIGBNvh6Qgs7xyfpLuC/HkhwU4ipFIOD4udhPNTzo23w0QDTNcqPSoOkQTz
fP2Db0KrrrJH7usYVxorIw==
`pragma protect end_protected
