// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
oiyBYnLUbnxAMG22a9KZVTy70eYkMb08WzDOb2BmWDTY/3iJsWz7gbGkF/x2iJ5Z
EvBqY9U5RgVZgLt9M3cR08vQkR3xtLFtFsjxL1CuFTKSSMQGzXbAkdD7m4YynPxI
EO3u64AdJkcl9/hwyJ0jzYApYyI3qiB6Ou4O8Emi1iLZ82jU31+eeg==
//pragma protect end_key_block
//pragma protect digest_block
69qwfOQcIBf+4zwkOYFRdAWjmTo=
//pragma protect end_digest_block
//pragma protect data_block
tojok/WaFddk2aOzNkA7SrKC7us5kPEUSB9JkwG4G2+ZVtPISzE2wp3t/MK0C6a5
qbkXs2EJ2HWNBbWI4Gf04TNcv4Sz0z8yEqczCJipAm8/ddw1mnEiF1pvsAYL2B+S
4f+5G7SqV5jp1UG6q0mNVAIp56T96PRFfuP3dfhdgpEmUY434vfUo9YG8lTi08sJ
Buk6GOTjLSVdYQXLViSsPQEjYbty48hzaCh7u0dCrGQnuE27AlQusx/ds5dN6eVc
nzhqCFVHSEqyH49BLwjJk178RZQKH2lajSmv256MD0750fWIXR1YX4gW94eN3JD0
+4X7QoLi3TdE8QA2aJAkCmL670M17VRIoJlX4UMYYjkg4bfs/5gVLf5WAcAkzZ1l
jE4x1AsZv3YwouGjMN/Mo91GWut3duCpR0CTfAA68zVNNw8QE/ZnYe6+uuFLwz9e
gfetMrntHPYgqCD/WKX1uR4SLXldHEuzAzQlQiBKPqxCkWfUM69duZ4jrqSCSfUF
wErd00vb+rHglkf13tlu3DanG8JYNM6to6Vd/wzDYZ0tZLyz9X0+uTW8OILXRwDf
plwp+WJ921mKMBmPuBDAwNbFr7/KA9+wd/YU7j8sDHWZcy8WoPWMQ1ZYhp4JMeTT
Bsht46Cl9qOLmUIsD/Pq/gcB+1AB/g0atJB1XaF1LeU8yczxm14NaNY8RnoR1gMg
SgqXL2JjOd+fSNlNObcevv9Y7qT7sSrJHf1kttI6rWNOqEYUF/4VQDVZ21K2PzFs
MgDNgOgFK74P3embuci7FQUWbNyi08ITSeydP3v4hRCvRbbWqVF5Ub91c9nZhyi1
MaPPakvQGohw3KgTDfrPIplSpMOxvI7DtzbVxcbIARI7wp8FIVCsHPwyAPwBJLSb
LA3XkGPpkjTeaK7v0lTxSN/Y2aSC55Rt9wv4u0GBpSH2yQT6yMdGYV6rBzhbBWmy
HwWrrynde9GkpSIs2B8pjGxcsmR+qyPTRNMbNZyT3051aLCu+Pma9Ri+apO1/dsN
Rv7lAIDYyTU40nGTr9amfX0pETWhJFHLKcysBHV9+7o6F3rG3iik7PU9lh8SpAQJ
dHHliOaWbC5+UhUJG2TMh+N5rSFkoRdL/lis8cYWBIPkzEFEVTHCgpZphfS46vB4
WtFOZe59MiVYX6C21pumvfwn7YBWmifaECUMpAt62iWSUTE1NouhxLe1gh/631Pj
nOb43S2Yx5EhtzbMmqj4PZad3afCDR6M3NizmOYq0eDuRC3Tzk34MR4SYWSG/eKH
e6g/FdvhNPc4Qclyy1DHq9Fr2ANaI/ZJHcCYImowKDaTZAIvXIJmc5mso+orScuf
X+BEtM2L59R8FMIWlXmVI2E6HhzJsaOY5Ktn2S9zrIRr96AyHKxHWFsrC0EaJ6Is
UFIcLtk4ejYiFBLmMgQOGVx4Wn63Sc9AY1bqiWxySfJxbNhtRZSreFsxPDvsllz1
0I64NUdpAzB1K3nO8nTwK/9KFYWbiWuF0I68LS9qW7OCU1W8IOOkwAwkYE+uC4IA
Rk/oNYSsAs3XgEVWhxSyWqoZ4c8Ydp6yw/Ia553gLZVJkY8U2H65CosP4g0WO0wJ
wfDqhqE3XjFrUSnd/G7WHC/Un05bhak3OPAL5F2mQuoHdjsueY1YLU4CNk+SCSp+
WwMhowLAyT5Hk5UPieUZ7+jhw8vm4TM633ZyP6qyfJdF3/ms5CN7Fflrexu4Q+Y8
F/iz9aZZKEiTVAcT+IRUpw+NcbR+WomUC7knveEsh40x/5GaaX2lO714zjSzoSRX
50zYDHXGs9+OxkRz74WfR59Yp7z04e4xkyHPPETkZMiMV5fJN0pXLlmu08dFCfL7
Dv7olJLtKo0zH27COHV16Bf9l4P1B+zWn/fa/84VdkUFh1rouXJVrqrxTNIZCjTn
VXMMDMULWly//jMBbk74/rys+JKSKnpbQMNqXI4dntQA+2sOSqL6fdyI6DfttYw6
ZxoFbdfZtoxR7sqvRTWt2UigpoPcP2c1ADFk1SdJryBVj9rCghsBGM8G79pVpcgr
oPci55Dp5dEGo7FI5rLLRjMaVWaDJR0HnU4lYnHMDyhdAMf4SpiYUWUHytM8eLDm
N2ev5MK5gCPKXQuc8UrCLYuxpQSHSUurF7jP8yRBc3NfjuiShULPucM4wmHwvDH2
guPHPMx15frVCeXJXazWHovitzRkodHgE65se2hK6Q47kzN0sZJb41R0U52E2ilJ
4KXIcGK5dV8ugoW79UEefHdjv078P6AVWfHPhNf9noZcVUh+mZlWud6SusQYrLsg
EyHusJ7HIrl0nG78qM1qVJs+Fs0T8om/kWir4qY/7fjTsFlmd6WMyRgePkD60yjh
7wc4dM2P5YfhWPan5oQJfcHS+euCoa9viA+pNY3a5RSy+Z3AjsQhZCJzGBwiNLvs
4Mq/gFUFUn1hryVDBUx3QCNEyXZtzXf9KcsCo2dnKXJBT6jlggKtk8h8Vp8oixCa
4tt5mZdtyi9e94QTjaFdTT4EyLgpmSgqHkVv7XJj79stmjWYkqfsGJa0ooG5HYaF
yFuk2g0AdXKgdIBPTVxKjEmufrQ3e+moTaX4nXjjVojG68xgWDxVsGvpEIqejsP+
l5JFmAN1+suM61YyVWdc135hIWgymUnO5FzW3vCeUsY5mUy0EOqHy8TycjUbbvnF
UJEY9fsKf23W0x06u091/k9o0qvSoV60XuUJ94Jr14rB1pwsOPjqvQCfyKurMAi5
Sx9NGhkePTDSFJATRa5MPEQSWsH/wZz2xhdbLRZpabhv8tKlAM+PmGCqJwcoy5MO
9S5PWxZiaQO4qEI4eNUH6hYWRXpdZYoTChvewm6PGP5Q7OLKYtfUIsdZAt0n/hRv
FvkZ0ziJuOZPtNtaBA6kgSxlyIAhDLI4ilMkar5s1Oa7I310EG2pbIxzNWGIMEJb
rXqlCCMqHg2lJZAA6fNut5+479igmtmmyX5HMaa8XNX+vpvfXjj66YuPSwobqPYz
oVwnycxhxw64AEim/akme9BU10yzSHfT+KdVS4C17882dnUUX6cszPk/Nk9tdtrF
t2Oo70QagB9RDSdfdBhSl7mSwxnZM4KjUteDpw1LBVcX+aACXhfezmXzmceqekSq
SVKIqhoI2abreLhsKbJn5AsDB7G2gzRGRAkAN96SWc2/aANnDvOWqV54ZkZHzaSY
yD6eylKCZQjhCx2uyIAMJSNs/zaR/lZhqGSgkhAp7BA7nxvrzmUrC4F+gdVcAdca
LdpFVf7tWrQqDvcOD8Vs7F+/EFJR6H5jNS6NWIwZAQrTTy0TDv9WDrApIMzYftfZ
zlQVTiYWc54Vezh2gNy/3xy6bP1ZyeYgO24fehzaUQcnJ4XcXoSdOi+kaXd+ADvy
TQ2GFYjacyAwhINZuHeEmPN+sGZ7YuSglOLfydkINHINCsxPFEYyDFORuG9bguD4
KPrLwOGEHMwKGiXkQcwFAoAU9UVKemmktX5Pt7t0yN0cr+Z90E6wu4+CdZUoLLCj
adwT40U+HE8yhWsbIRFh8TXjMSpWpiZRmXYLtnMuVHZxspo45hIg/dVPdw7SsB7q
+DvW7wsoCkOnmXuOqvvyMY0nBogRmIBWX4nK0pzhfEdAeBcnWzaOUFpgSTZPWMQf
s2sCEocE0u3FSYKhnoEwF4qa5X3crFky62y89gnPoerSw5sbT8Z7bW84UIRQUDQE
N/o9qjfKPNXeP4CZFK33d1lna3uJeFyrTvfQ8tryJ5XWw5hPAw1ZzFjSLcZeqwjF
FngH8HH2mPPwquMft6PdOlX/TPOXYpEUKxCBeQDngGaOElb3myP4DDzeacbdtY2h
8L22XSWbl3bhUTmX6zR7LdapsuWAfrZcjKTSfVdeE/VcxGWkW+8pYqMlWLw6h4ox
Au4hexYTBwhgWBgwchgOkefUAk2zkttqhUf7gNvj6Q2o5beBYSAGoVTjSLpNtIYE
RhpoctKJAU5yWio+pZDJZ1Y7kEQsxLtktzj8YATZRTB2H4PyPuolPkAeQ/uGPiwe
3L8Q5vAHvXF+h1MKU5lbcNjbp65bUmdlOHE+ej/ACT5Ks+rkFjZzf1mTdFUyH8LS
eT072YFxflcrcjQb6AsqTdVnvFW0JdG3Or/jg1jQtrttAjdRd8ZsQdVIuqDlSQtY
1mNsCd+QCP5rAP1ywKWzafoUVS+WaZSp+qVYxCHxzx5XDIJO+rIzXA8Ud48tdY1o
ieS28bYsoHmqXrBK0Azj2HAKaAh0QH/b16rm3lhutueJc53rILwAPKtbxynIhQiF
bUkcqr//MXK3cY0Vb6KoFjNhgnQEkXNsz4Tc4wxSSHdEv7EaKPpILWpUDnvbGZ2j
iKgndjIgRSBNBCklPl5dC7mPYIaHEfBFejE7cJ35ggTwh1/E3v8fOCficiqGLgsC
sqeZD3DQYQpfnV60aka1j5iu/fSStRRlJxrc7KrJxKlHgt6wPqW2P/S1bzEk0Go0
ne6cTIWQjq6tatKWlmLGYXUn8+pQD/IbTRMLBD465vjrkNmrlUvTiI+6agFsVI+e
mDB/0Wneb2qOxvvwBAgCVBObCzchFASp6Tj/x/9I/QBCuSBrmpP6s6k681QqnE4c
wsISTZhopcK+Xt/7Pkm77S36COkSMMpa2zJJjqh8nxRrce2DvqnF1Y50a1bWLcTr
SmOTPZRM59LB+41AgVm+VZGW3aXpabMJyb6hgisx0VYHHJ38eB/RTDLkuVTssdT4
KdxUhJPL0oWstAZiycU4APi+ZC0dZyoRkwou64EuZo+s1l0L7fQQooTDeU0QvMe/
nVrn0EDsGFBqNY7veFpRuJH8mJHNWAIsRojhTcYhTPqv3QznqeHLnRVbWpPMbZOB
aMQYoTgxeAmfEf+6PFQ1vTULfb//okIs+qyb45Sx/d9R/SqINMloWACzzTt2sRGr
jUPpiffrJTOWsh6G1ZlUZmeKsvphqbOZZF5zQqFH2Yt8eF9ikYdtqiM3ozPYLNXw
oUMYejdF9UjP+Vp/l/NmSWLhsTPtj18H7tKFQtnjQsZxdEpoz42AqpQZghX3QBEE
d2ayVNLoncLO1l2uhRyKywmJNLPeJsKqkFaxef1wBOo0XFCAxdK9JbQsuJVCjdxf
2AhbTC4Chrw/lmTL9zU8KkKd4jlGRPvCRHF6onPGO1P6508TnJxz3l6u+G/jjpX6
hfnq58JW8dn1QFUchuogivG8NOWVw8xCPi6FEv1Ld25kOx0/LbH8S7rumDUjkbhq
PsRfXD3PKUQ5K+wu0g9U75v/eyVGTcAAmqNDMrxkQp3SGj/JRjah8StE6cEc0Uo7
ZpCWgdlclxagH69ZPDT7CZKbvHFg/s0hnFxc4gD9Yil3EWfXPvNQe5rmnXHG4hDk
JRxGBQnF5/F4i/HmI+D7qV0yCS5tmZ/zuFDAD+a7J3jamonDnORwTmyuxXDSdTyW
MzyRMrezfws5NfAuCvzWPQL7srvyEUZYWCHxZnW0mN8GH+htouOBySMfmdD8jurf
ZGD5EGWzmise45FyYN31nM4fhwUJeZAhhUehele1GRPnCtjPmxS2JL1F3F9ObXFi
pk8gcVNBd+TmuFeaoAmRtJrvSjAOwhYbcSlUtNm9T+8iYBHsEKzrDcWEQeXW0kpq
spcUNwJ4BU5S6VoLkG6q2uo3MQbBn5XIP3I1lXff0dAVaE1NGMXlRHjzI4C1HsHw
bALLD9WiDBa1PUfv+vJ0YvlhpT2v5TAWHBHprmqxasOWi+Rvs0RSEYSI+uOPwOEG
aFIQNsBz44VfVsKe+RxVxGOoOLJhljIdnGM6B9HJwf7TdFXPqRN5JUtQ+V7idhUp
xyrGa2+kohrjOnMmIMLRFt/3pzMthXNJKkKAKUZrpvaS+HubkuLH1GRKiy9dS/sV
1SqSAevZRR82NEPkRFiOZpnIVzHXhcu4T9O960tNxrwKXEKYvWyfYsFbweDUt+Br
nD8zaUNgUa698XiphwCbgF6bnAAyJMOt3F8o7w1osNQW9K66h1ygYuUPHrzzWAXP
R86k+UXGbS0QEkt4mn6nbW+qw0B6fc1Ok0hKqo/OXM1X4GvYMlgDby9nU+nqv380
554IRJipoCO3AwgYyQoH2oiMIHRg0tDNq4AOGJdY6CSSbsef+fltoBpdtwicPOtk
Q9grEXzVVXFyxSb9WNcA+6Z5lYbIdpyjNTDqBFmUQ/jSkdV1DPg93QfA0f/Ksd4j
sxCLSKe0ph+EmymAlk46OqAU8/gDhMetSBqCVFAQ/PqmDzku29Kbx/TVbe2kBNoc
iIwJvp4R9844idaPO72+Us1A3upfE89WG8w3S60j1exUAAiYiiC6pd8hdlFLA719
//k9VKVJcAeVCTVz8JvHRbOtg7UjW3kyFd+y8rYv7c5twqmDqDhJ3lC5iCghZ7+0
E6yrEKgqxWiqUVYPPITujgKhWQjcv3yBGzJrmpiBxWOCW0tzJnYihAG7kPG1vZrS
FarXCc1kfJ4sPdRSfLOXgqrSYsr5Tb23HQxDA9Ak450l6mo2llqPY3hGys5yqAnJ
663Fz2ctzA5sY4EXu4EYA6+nN3N5PKpz7VbL0VsovwCuSxopRgpKjacLNa/HkDzC
mYo4doWnBrhU5kJpz+/4n79tfh9ggx5189U2bVHuR078poVrzuTZofj3frCoBNWf
QiA4/Gq/j+jp2eVcLpnblr/YRqvA/WvX10JD5vByxXNIXvFglwE7P7rFX0RoHDRn
072v7Ysnl8HIkrdeocWCzcuxfLleY/XdPFWQQDn2rIhmtlq/TPgelfBxOK/MKR11
B+pPPzhX2z/MWOUEC5yi3OxUQ/N+cRWWFKeai+eGlNUJ8FvEjM8ozYKeL4MoxJcB
MDBVL/bAkyW5ftZZGjXbnt719+CDvMImrMEq3pU4iquL7xYjXbvzOAoYGca8B0Jy
ewVGSCSC+/6EZ+SIBrblXfyo9IEHpQ9xZCz3UQiEgd124QTYNONxG+mcr5BgM3Hk
84ZHYKI7vBaHr2QHAlwOZdwAQShgb5yK+2PPbdnxJ4WdJEAc/dbOAIdKPuXzYllM
6avrmCe3WDj5P6VXXMScBgoxGKELQl3NzcckaUuuAW0Zk5lkL72LiDkP/ICHgyQF
SFUONMeF5BlHQGcOaDEJTSXAzHXHMFnzWmDx0/IRqVddiMiWOADZQ+7CsIq4vvQT
M5x8iJq3Tb3kTWlT05o5ua4srbTVvyApWMnfjFFLAbAuhuALVKAbDeFCpRuJMzNL
tEq0ah1p3Wl25wN48+fCUyB5TdUmmVLnNN9LRezVtqUIgnfxNqZE3FHVNv5B7KDp
Jj/y9SzP4z83gyvlpkOU8+Bw35E0sa0ethOnW3Lo9OA8IrbTpT25D1KPf5bQQO0P
fhMwjrtYCB1AxCQmavPg1483JYiSUiTpS4p3eIead8KAidaINtslFvVLFBpZn1pd
yFjjI/Cx4Kn9QRHEP5bUvPsyq/oMZD5+TGZ6fICdb3UvjKH2qsDVtmq/ZkTGfZfE
jOYUpN4fA2mhTIyK5NAoSxJtNVwGs7jtJxYX0R6+dOtfyFuxKE13WiiFilHBRlXm
cHPnpjvWD3ddHa7uFdqi3bEXktHVmOBF+Ug+9c33ysshquamNDE+hrvoe9LFZ+Mj
nM/PAY/+sm00XNxBKfiSoqWtAvQPXhnrZwZcb8rF7CIG9qmSyuUZ2SKTr0DknsqJ
QqZ/qA3OSQNFFFlOFRXXfxVBoA5eTKwSzQQfVtpOGZOgqkS1BawKDZaEp94CLApJ
9fK3IgUmBgLZvV5Jw8hcS+Wz6PdTHniOGnMUQf+rlWXA89jycwjlHMSuiIz+DvfB
vIyrYPWyDlpOr12GXGeQmCd+yUa3G3HbGd4CidxIpBMUUDr+ebDCLQRGJHmW+dcL
KWrFeDuE/EbY1pRe1r9o+6O+/izg/1V6IToMQZwZRzDW5d4CBaa5boIb9LWnOiHx
cJTbbfCA/SRq9/opPsa/s3o8ID1NzBi5c6O/ywEqD7YBtfEv1hsKYRYd/EGYHMKM
IQLjKyzbGwpBEqSpj+puT/mgBnmaQNXKC3PWWOH4cLXd+4bSnksmY4LynRiCCR0L
ktYEVvV3fd3pBhXQO9s4NJTpJM0hWTx970gjYNy3WMYb6nZ+Wlwc1euen8LTl0JM
U1q0e03+kfgQU5zTF9AT9OESMyUwK0Ct7n/659vNQHhBu5ihhD2gj2OKj/wuNfIz
T5H9QmFfA5Ri7n5Km8yBtCj6bhTQTbdB9xPhkg5f/5+APr1mtJgxk9DdHaMZt71b
oV+dQhFl7rpIXnRh/OSUCkzbwqD/Uy4W5aY0iNBSiiPzscFl+abd07p3GCej8+hi
PkHLp+Kg9CsEE4uZhYW6CDOLFkAZbBYE/w5osU/X0t+YmtsFhhY58xyA+Zcfpwky
YIJ+OiNzykgDPG0Ifi38nhmX/LwEYGBU4ok7qOa9PkSjt4QXQ2ZwdQ2hCufuY/wg
p9KtoVjSsi2avs8Y8DkxqCReSLetoKuYvulUyaEvWRg=
//pragma protect end_data_block
//pragma protect digest_block
H84q2123O3/13ppVtlyfRiM0krw=
//pragma protect end_digest_block
//pragma protect end_protected
