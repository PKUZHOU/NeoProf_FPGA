// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
iLAJ/S+F5+0uSxSUlfRkPW14R1YpK844LnjqvzoL+i4HRan4vkthqrRQdhM0
zBC5TaEDvxiKRs0OpIeURz0DgkT48xdgcYtwb78Rz/INFsgKuGI3UrFBlOil
6BGUiC0D4Lf2zNYlcgSzwz0CVCpW04TORQulBGWlvIokWx6fMQkOLIZqRh6i
QYxcbEmO97zIfdbhfAnH9DcYWAEdnH4iX7/og/sHRpTR6UmQ6kSh/fxappPV
HdR3RR8EwVmC8I0K0pwKOHPF8CrFY29aUYC84HICJ361Sp5j0d7oHUtn9b/Q
sDeN3h7+L6NGU1lkECOsG93pe5gJVD0Gy4hINagWVQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
hofyz6nfhLZ2Y2SvEy2a88PuBySanFD36qYDBmW2nayaeCKkHC+OJXoxRmn0
y2yYHnjhddUy4wgmtXgeclacIdxmgGnPv70PHToGpr98HY4LSbTmTE1tjWUM
SqlsnimvAqU5JdPCNID8XAKEez4t26ApXd41cD6UdNNrcjYpGV0lTjpW9jwh
FaZV4Ef8oTsEFMx2eCi18K5iOIWypcCF1WtuK4Pq6KI1R+HB71k/b/WLlPxK
W9uRhTRoOEG+qVRQThoAqusZV1pq7SrjE5dWgr10s1ZXCQ0Q+/N989Q9hQVA
yRWnA72Rgfw5nTytX5Km7ltYk1VPVZ8CWJI3LbCxIA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
oeFY8Jhod0U7+fTm+ZFDyhfRDF+MVtdQdzIQXSKYqNcH618ofnJ052nKS1Ed
N+Fa0Tg/80RUJ3DnBghC5hsD0l5cueWoBSEaU2JmkVQQeqVClO7vj2vDPU/9
5/z6w8Xnfguc9qeUoZxT4CDZidDeNvc8whKRri4XDG7QfAmHmURUCzZYGsKx
HsjqT0gsIH+NEaOqpvdwfIBSET2h/57GRS9q4l9FUSZf23lHqdfIRbOzBwOo
Cc0DlKaml/Hh4QaWm2eUJkgmuujKYylYoyvAbMmMPNvuN56RpcNYfM1P/o5p
WHfEOSwGoOg4pZQyJyw9U7e8TEbqXfTgJtotHIdTYQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
hhohgV8KGjC0g2c0M8fojXPqz0LwA2JDm7stHkdu8eJtXlBNEdSBEKrKavRG
WOdLkH4BMaPtdHo0A7jXZ6b3hc7fAc9tQjMESv7J9672rB8xn/ZdsXTFhuVN
yRagHUG4DFX1YnBanV6aOrO2TrEcE1M6WlDp17bsEmGo1Mrpm04=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
xc+EBHrzem3iEKoz9EGA/HmljGl6s52/TeRP+gLw8fUHTMnlKTaPJQZFIuBr
+fMPGl7hrNPdIHIQdUGq9roe2wnzsJdLrOhUJ5lPIBXYRmYkY3hxZpY6OYQ4
4o40ojR6b11OWxYOquYASHgsPaL1JtlXZAoEPIATK5su3bfNf0TocjnVwps6
LxNtYmkvZgdoZ+NrxZO4FjRBYNbqhnDP/AT+RgtKIGhP3EK00gEli2xucBeM
gXnJk49Ze1SLSDtm5VYVJnqKOkjdH2oKAizhZRa8b7v28pJo23Waf+cGG1sL
yr1+PdXBZXNA/M4cy9cBa5eBuMYS6Xeb/7xYa3m/xjh6CRO38HZ+3GeRERp4
8dsucXptaPT4ku9t4tCaDpf1W9hK/l33DQ9K8hFOHSXBWIOwQFM7sq4Tj7Y8
Sgo+2vsqS3MwoDZHe8i3hibn7hoLokGjeYfZEmTdfJB96qUasjnUS6tKP1cQ
SB7BDsFSTEgAB5p4aj6hl1vHqtuGqrNV


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
BZuGKWeefGenZ1LlFgq4IfeOgdlinKAXe2EOHPxfUenujR6devRkF+w9psTl
xwffDZ2SstWJPZF74aiznygV+RQEwV8VfwC84F/xpL9gKY5RP8OlSbBVA4UL
QVaswelW0MEygrmlhncmMx1hKQvcv0V26fL9EJBahtZwnHDCKhY=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
i8XS/DcxVkRH3+BLeq0LTLc11QnodUy5yTlIoTd+lKeg9b6Ja5tXvgmhB/YW
0LEyNqCf7D5mU4eOI0hF13RG0wJjM+TE2ef9UgtxNAnYH1oe00f+kI+TLo/i
TvjQkGcA/mHFnntnDG46ezAxxerlsVb76WnXIGpX/rrUeNy62I8=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 6384)
`pragma protect data_block
T6VCv9DQbwzZP7x+2dnsTFLC7aaQcaYr5o8fynM2i1CoOMtvu5jYjn/uN79J
tKlCWn+TAaOZhlB909H2ZiLJe6njmPj6hq6znT8G5U2EAafXG5/AqD6WaROa
wi0hfkizAoRc6r0mNgaKRql/R2A82ZOjY/zSWQg4PkkQvjNwbrDz+R1NvHT1
oK9gmRH2N8rTQH0qn0hzFH2FRqa38L//Dn1iwMMjLMqj7NJfod7UqcLaLjy9
62irh8/LbyTp4dXxw08LsQPu7+6iEEgvwprzaKs3sMXEnuDLEC9aaV4z6U8V
/LAYqQJt481HK/InA+isgBdFlq/nFtkrOdFEDw6wSI2FZCaZKqcOasUW4/rm
1LnRA5ftPShv2UWaW0tWigt/jSvQBMRmS5NgLH+KbTAbb2D16bTuiqktnIOZ
IPqqUmh/c/SNs8p05Ke8TZUycwopeHP7/78cAZ0gxvT8yums6E5ufEhnCreP
e2d+uaRcyVY1TZCuqwQVZeU9hGWVXWuROfLKxgyytPa748TUy5IUoytQ6l+N
CGr3IrUdsChdgEyjOzI0M0pCTWjTn3HrlnjJCBwxIn3XgFl3cfiu3CXBew2+
mJIAxl5uOcI9HmBuVLsAOaI0h/0YcmNIz17eNoNfjbDDu0yogTAbDk34Ezqk
VCCgzcCw46nA7cucc5KydvXcyKvlXTtXjUrAn4zGJ8+JgpxPvprCNEly7Ie7
zhzr+CX9Q4Iio25OE6V28nZ95bT7f+8IWSE0ZyYOeashV40QNmGd6CNBcqRH
2sINYMqD0iESX+OWUgVknIwQzAfJ3hEVL3vWXFqlhZLz8Gux8Vgt/trsshLJ
UdliWh8A/MH5F/Dd1u+d8I+D8AZzW1JexvGcH/zjaH1T2mxIowpMci4ZIzcE
c/NRBp3BdcRrvsjSsNgM3TmIXu5QATBa2CL3jfCXVIoEYxO/cBcjfVMtQuKP
LzVFmZWR928YPgMIZfkiWdUGPNk12wbuUrR22eWgf5FR4SAiFZRqJJA2SavF
ChRVri7y8VzTwTSex2OmatHx/QlF1qagoH1dG35UZ3LgRXGp2G15A1FCABCs
8wmAB+XH7WuRyp78RFx5cU3z4hVXxmf7TV1tB4SRC0SieYdydDohrmN8J7pQ
R3AwCTnqu7YY9AH71qC8Pp041gw9to410XLIrSIOpnMDgD5Y3OsyLH5nQcah
uMpPp2cmdiXOngi9x7BVpdXZaFonEkuFqe+oMtl4lwc2cw6Ocz+Ofxqv6ZLB
7tWZRjSYYZ8z6eojH0/mfuCBEvQ8/Yh4qoDhhkg6CPu1jKVIcGPc0bBFRnkd
Wt6PLPYVP/iXm4fmt+X32sLw4EqXohZenO5FBEgh6mIgYJHxfxEUkXO3ALQ/
amMeiIkd+WuH7FsBeY5e21ogAxvZ3+yazgK65r/ySCSeNIsQkRKvIGZikzyB
AVLJfdXpmnNIDBNkJtQ0GwiqvvkafXxpJN/2h40H1gXfCrqLXMAdquivGT41
EQmuqSexWrXra1a5vp2bV2Qfq7QAHU5CgqqFZKGgx/481hxdsFm5uM3qzODN
oyWcmXFROInRliFJsKdM5UKCDtlbbTnx6Pe/Ps5MK6PdKAXl6PhoX93d3+tk
LR0y6UpDEzXMTXEIFXKkKVyarBaF9DBe/1bdtchaA8yu3QxsX+/y8kDYXFCx
zpmv63eecLPSE8VU+cA8ldSsU1dE6iwPfLjA5iugE9X8tJm6mKRXe0krBTDe
YWNUWCywLL8oA0e5e1pSAqMsklLl/9GklZFBDCxMDOlgyG6UgVMwAvGw8ts3
g0pRK9Q5nlrmQ85gdE1382LR0J/DHPQr37csrP0C6cd1oWPIaodRv5hg4HiB
cUH2ELbKf0GZfeqXkgQAQdV46E3bQB3TGvw5tE2ykE3Z+6WqhqVAYkUd3AUG
E7pQ3LtZQpBDFw53fDm0VoHpLAO3OUnf0dKLn9/4ewhEqm9psPouQvtDGzra
nISUvggScoRCzMerYTBXWBPIenMfzVBEelah5zIP0anKSlaOp1G1YMbHfRKd
H1J70VzTuYwK36YNni99fHs+Pi4HOX0xOzkp5RgZa1UnE2ogqdxuqJX6uhDC
3ZEx4daJ5/Zr5zd5WDnDOZzqAgLyRrgk1oZFskxgDhrpAfXDeTJ71SQcm0Q7
1/qj81X8ZUr39lFIZT2y8qvvVfbJfqUrEvyyG3tHyG9DaW+b5FVD+aVyQuhZ
gxPumz/yYfHl+cCRrP8Novo+bMltAYQxtoJIwKk6Uq5P/F3BDUy2LkELRa3T
IeQnd1aTzGLP53j/Y0jZK2VKFmKTJsaPz6ZDb2Stqp7Wx7JuvrNruV2FQ3CI
O4A5TSlYSE1U4OJ0O2Q0/w2lmuyy/bIF0eMtWOc7iQ9T6CX3JyuA/6svpLVg
iElZGuMq5ro6dJhvDOaidadBJOw/u2eN7TpxfDKj+2fP0tjjDaDqsHkPfDC8
fjsapuo7flIlnsJSL3x5/RHGFdAVoSO04rUOm+2d3vnhQ1k+Md9aKJmcORqk
2HYnyf9rI7419NhR53Gi+KSYvwvYq5JuIGdzrPj00J0EDqYuW3SkjDpGk08b
6vy7ko5TWiLoBnFuztJHMZNGeNb4w0bmtrIPS8QmazXpscjdvaZ63Uk0GY/B
NVgR2LmsMa/5HTB+QIXUd9wX9ztpGHhmBCx0hUVy75Iq5Q4/vIzsCuQMKN+c
NR+BoVwG/Y9dj9vUhDP3CZ36VG2e5Eb1O6743qbnYSog/KEDWb5T0u61+t21
kTubApLcd6j0anC/gcZ+BFpyal+oX0wnLTflrrzehbo2VZLoCkwCrVdDfMOQ
jBvJBxw7NMNsJ/l75f0R/Ur91g4mCRP19m9nCSeLpBFFtdrLBSpWP8JCZ3yt
2VSBrJUc9eFPMlPaFaF/HcxFp2AFPAFzhgcJygkSVfkYGEO34gya1xUqNPhs
gFeHBk5W4Tovn1ehuEcgfTL01zwzEAmieFViTRs/nFuRd9KVZa1cDJcpax9x
z5kyLSjIpbxeHa3GvIxbEoh6PEjxgbJTyQeWa20ARbSqjjsaMCJYoyqtR3nZ
13mKxUT24FehE0isSPZfFJdK5Wt/+o9FbTlgSit9yvfu0mwWQrJ9JN6AKmI/
9mcYuqRnWgD27iWrp/JwJaKE6Uu0yVPSW9wQq3rWGPzpXNNDPjry4u8BL/Fl
tArBf004wkbPM1g/FNYfearrmqL0faP3VMDp4Wlg4iXi953R6Edu5cC4HESZ
ixOjKnHFA1PGYm33AFlhSFvcMjKQe2ibiCJSPGkLJgf6FEYCAyB2mxJyk78F
SlNatDDJqeT/LWF6er0w0lL07BllfukrbNFj8+MRJeq9k51x2Ssuznm6StVd
bMEHKtY9T0e1APCyPTV2D5TDrhp7SwHlJiRaxg7RcicRBfSLDYacVWO4QB8o
cf9fAiLTOOuWSswFmphagWlGvy8RMaSZMOnZCbAV4pq69q14Pp11YH24E2NV
HtxIviL17bVHC8/B3vR/lJsXFsG0jBhytyLAWkD3sJuqKHWVjOIEhOiMX1Vh
VLsRAWEkD2pj/ZXm77CmlomE7Yn+bRg3nGUv3K8LKaAE4Ft+FgGb/4Lr2t+n
z9zZOaxIaEK6Y0QKr9NMzcFJhzPez+oP1WRF47QfPHYSCSb5hGTjgfMbwqCI
VcHTv/WOkeWLouachzdr8FPbrERRCvf9oiyDaLIcgxkt4X+6XFS0SnGmS2j+
sbnOiKDBinIXnwTDy3QGXH74Q9dsM5r+tzObknCe5Jwuw3quB6zrsWbt2p8U
7ruWGF+PEvtaRjUdcp1jxBCz6qbX6bg3rxmphdeFUUE6T0s/V6pMD3kgv1Op
ViXXgtktEfqwbYlOSmD906B6oepHnR3u0te1BuAfUiPCfFitgVg3L2/VAYPg
BPTwPVz26OXF2lvzkT1JJeoer8jcKL32vcMMIIYZdrt4lhtDKz8VwrADnZDe
Cwxta0+TDU9hTfUQXsSw6OmvECtklw8ilk4BFNJ0DbSB0M/8egj7WbUZngCm
pwAf2bt3vOAU1kIxwkkwTeXHgrW4c1TX2aB3aaFpcvYOu6HJqqcKzop/QVjT
LGeg5gNJGAHTy5EB5TBvXr9SOv8PJK24x1YYHnBJer65bLn4KY3Mtrwj7/Uw
Rztn3r+yZlM0VPZz6vlSxdWeqvvKz4EikxZ1j7mP+gRi04GYimeH4zcA/5Xv
YoQ105iMxOpCAr2fpzQQsbu56AJtKNXnKFFrkWiJxzRwhAvzuoyiW7HDRJ98
THroAq9Cq/dn4Z0Hwt6SyEbElhtoCnxigea1lUyIwXdpwxxJqbP9nAi20Wl1
DCNo50MdFij8KAU9TQPUEwvnR59Jr6d9PQb0JkCnWbI7pH3GCBalAoREJ/TL
xEpharr6KW9sjB8Bu5F98unbQPrZNnIAyfTOWSfp5NtLLG4FsQ/s4R8LO+dD
HkBs32EwniuxZ0xnzKYaGTXyjS6+2UAuDcIdqtJWVPGcwgT3/S0UkZLlAyds
CS7OKCsVJZFrgZE9SrjB2ix26BJ5JMhQTtTU2bWRIhgHc/xRzbKI0OorXkzG
Nlm4HYgwUUu0hxWXJUyZFsAK7eenAbLpOeGTjyCpHcOtyWzPX4FiOEuU4qcm
QxM88DK8D9m81Sy59L+syZKw8aaPSzF0cG5dx0xGCR2PjhE//GNO9N49GaRb
4yQcO9GrfjMsf3mgUt9kLLIwT08EUoiwyRmN1SDxH0Hn8qhvFGWuEkmh0TMj
QLW0PNjlHAOzR+30MtGA84GQ1CCMEbB9LRVFBjTce/fVNYGg6isAUjOLGuJv
9rX88ocaD799imJzD2cdTSxDw6m091WVErqxdlLdRcSPqJQi6JbxZPzaFAtd
RiHYC3I+c0pgk5s/MQtQ4Dd1w2iLGcMK+svX/gMZZXzpTwmq72FVV9nx6/bm
bRcMrTKNMwSMnaaBqQlsA85kavbaQQ0kAmUc4O6qMvLZeG8fXWwtE995NUZ/
ZGsABSg+Fib0PXIeYRYlBhAAbW2wMBVDZMBkZlPT7FWRw55D+eynuLi7AbHd
Xxp0ocaVuOHAQFBDFnzk4nn3IfDV0y/J2QG+Yn/BGiwcMmQFbXYK3MvU/LM/
87GXtr2QQwW+wwTZ5PKUXawf1Ko8DvO8ge6J5gaLcDJuw2kc13tOl+RYkDWI
OirSrGUCKpPbl1c4ErcbGe69MIFf4bV+dXt5TPOpvIeGIeQUjrIksYPiAVdg
qWqBqF2KXCqOD7IsNoeu9Q5vVMA4OGUyknW38dYSoGF8Vv4yWFcpsRLrosaW
d/vb92OeSQEa4jOevyaZT/ZJBnVAPjCWFU1BzlMjqfuFdl+oQhYUaGGlU+IJ
zXa9u3ZJ4CfEf5AvakNcXXTTy9c9URXitHhuy6Ri46mcmqcqZN/fSKUaosgh
hU4ofAlwfJz8fqh1LLMcGNY66RUMxqjgMikynM6yOfeUjnT4pjcx/0Dy29/t
oHFiVE4hghDyQ5+nfO9fPfo0eumXJ9Y2kgVA5in2qoaqpfiwcf1uBOsilfG0
Ft4HUqMUHrbNyKWC0ZjiWD0i5UuKw4BGrM0zPP//g/SwYKBfpkRa9CDOsGwH
Z/TFmBKNrUpRCDG/mxoKKynejGr20GKDiX98vfVAcRhkWxSbpAakTk2hbTk1
Lvw1eFPIPVKMqwhrf+cluhYrthUmkfwJQ/7PvattIsKBkQcmlfhZo49vz1uK
Ex8GoMKTGFclhdiRacA1+kWS3i5H+LaPKyJPrywpVeDEfrTPGozOd0Z8jdFk
hNxqd7WxJPTNPup2E2xWbyBhA1KhnWCL5OkgRIwNlytUc4/kwFzDvXiBcTyO
SsTAf+5NnXSIyiZgAnzOizqWPptm4hUfk83TLkJR3tEURxuVBlRAFi39R0/4
Bdn7Tc9JIimUS9JkQOMjpz2gWOi4khJc22w5jMOfA/6d3BEeJNgyXibCWbz3
xtSYdP/btZBn2ukzVl4fvlPQKy5DCVOWXQqH6TQsi0QaSScgAdbNmko2qTro
lNFDdOV51+LAM3Isdgcbgd9A1dh4x+9MoYsRm0/GbA+pi3UfB2sIN+ymA3zh
lY88TfJPD/2HrB8ACKzOmJBd6D1DT6uLp6U8RCPadsp5y2U7T1A65nGxjOaO
hsIbc1+CAwRTZqNBQpdhd7A5uPYYut2WdXhV0+2xfeIa+2Sf/4l8W0RUQ8OS
PFu3jhUG+YfzmJhvXIlnaGNB3zXpUvWGDSE4nU/YflOLURkRQFCjVqL8CkPH
5JU86R8Y18gE8aT1+19RtvG8di9f3N1lIBPMFgMO/6/IGyTbBwO0+rS3NmHY
v7cgBIo3x4KoUGMAW/sjSdQIxh0iT3duk/zVS4T1O/5a2JVcARcmiRdkXR1g
7hgoMecgEh4HD2DbjeRLSzqccSRtkoxnAAKLAT6tcfvikZAE+7XFJEr65Co0
3YndIJcVRhtfJjwYUOcptl5f4vxURAwW2BizhCtzCV7FEe2SBWFXBn94d0VK
FK9eOVZe9gb6G5Y/X4w5zIFiBsFMou0qQ4+6j1EAXcl6cdCtJvnuxmHmra8C
jgZPZmksqsiAF/z8/MsxyV1kcc4GitqG/eGSLcciHfNq+w+yWUoOPUoj9AZA
SJbIpsftawI94NReIKT2t10TmqVnVnu5iNcTjfLqMAhlqHtAjf230p5UOhMv
MhGUvy/NFgT4Dom8JwXE92gG//K7GAOWH33DBfYpySmxJxOoWjdUlUAdavCY
OnuhX37X1xji/Lf3lLXqzGdyAy/9dAgRGV55oEpl3AsLgHiVC3Zbraln1c8A
txwkKe1yapjB3qcgV5c/FP8X3+XTIfBbYBSWdlzZgmzyFty1OkSGFvQTBUEp
D2L3ROfA8SsYm9nrFNcbt6mHpcnW/bEd6nJn95gff0r8IwdOFx5TUjdRWGGK
ULT5JMr/CKsg0muQGNWtSxrbk9Ya+NonIZQxu0gsvj3p5uWb+9UrOE2nzNLN
L4wkGmKzsbg3e1kdUX8Gc0U0G6Dp7c5qQcs+t+2FCsLq3J757Js7wU5Zeg7g
zRlzXFLteb4rssTEKHf/EmEc145UWqpdGelHYldPdHSme8avg9vFkxSSIKLT
NXNU85jqu2554V78MmlgUnM9ra1oeUCfDrEbbB07BIwJK+b7qZWob1IVAk5f
gnWWYEeTUWY3iCTH31lTAw/6PSgirS6F0u5l/afhHwoy1lR0I2IbNNP9ihkC
e2CKz8uIp+NX0JmBp2rsRfa3k9Ie8E0gmasxHhwfItJcT708xrcy577zZ2xd
h1Wx9N7w+gYuY3bnlX1OgHBsBx8X4qBjtZU/cBYz6K/JFs2Bz5fbm3B/T64A
M3kRh39OxMltouwohRjGw+G8tsgmAAFqpo1rz9BblP7q1AiszlulzTjkAFRk
h2JaTvNuEeLlgIgA3VowPTON9bCIHAORxBmWln71ObD4qxRavG0SzP/acm1q
AJpnt0gCbQJCcRSS4K0jS57+OZX0jwNoGcYws3HaiNjTm+lIDZ/8Tf2MAn+u
kN3PJVGqeLe1cCbS1fjctcTnYjZmjp/Tsnq+P/PXa4D5QY7W+d666b568r2u
oiEfDPmMPt+VfNq89K8XzmEYf8lgOlSuWWkU0xfd467iF5Qzq8pwvAi3kQ8q
flGKU10Lrjiin6KCUagRC1ORyAecoci6w2cOM6/8Jpszn8mSLynBo3PpXa2M
rfUCIuz8MGXUZ+9OWFWfACXql3Tdj1aQUX3Kq1Qd0nfqgUobAZNLThmRPGdy
zn8Ml0ZDIDF1NDRjNf46CXpxnc7qLwZGcHDbpECpsNlYIc5SQk2cHN0f3hGs
PAZ1MDzRA6rp1mLnkxpkJ88EtL0qmTB28BhCvX9sykXmkDGeEgJZ0oSEKW7C
dUd7z8Eu9fHpe/z6lP/yFoB+tKlmd2OvtAjf85OC9WYt4fK8zDURHl4Rhj/G
QkVwXOB6VDHn14xUqfRDoJSsH9De307+93fKAfbrH9FCiWBYRvupQ5doK3lS
kfmDG8pV52qshGP5WZhYeLOBqN1UN2q7st34Dquz/SEvtU8CPXTnlMQTwjjb
mC7tCEDPsNBbzm/A/DOP73DHpkXR1Eazkozr5ZXQ8g3igtuBg0qdgjtSZPl7
vMWpM5S+G02VgQkZi16ZaVwjwfv78nBgY2/Wnhw0OdYXDCMzV/RCC9Pheo8w
zF/nlquN7Q6wzvg9q9YJxkVjg1rt4QpoTsnsOjLtMlxXXUtqCYun3X/8c5gY
PY7J+NFz/w3p3NzZt61/vmjXZLf7skoNtB8scvoZgiwjqZoXvndPShMUmosP
3HFTcWjAJfpHtafN3KE6tKtFXJNbXCDFZ+wjOnluogH0oBPCOpHaQbH65AyI
OVW/+UNnB1JLQxa/Q1CNlRBerc7iM0u62u0fWgHaCG9jdw86rhI1jIp1FlRq
b+tZSCIZOfMOWHsuUrf2wF9ZATvnOusqkPUaLbdyCPo86QbNaG6FwyENQ2PU
FdN2y+GTom+bClgunw06mHzZ1vw+OsZJAMWBoKAbc1Y/rUpirhzK

`pragma protect end_protected
