// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
bTZqedHGXY13L/5rAiHbMUMXizuqUAv8fHJTKKImdiUkLLRYOBJ0j08r0M4f
flHA+4tGBqWyBaAKCcF/0kO2QHAWevz42ho7nouyNh8SvqbRlRwKnLNhA+lq
iSn9NdhbDpYU1dnsGJEAZDHwK49mT5u5E5m62s6848EZS391jdq4bEfREENf
TlfqVMN31mbveBJ437aAUISIggZy8FUlwsfVj5XYaDWS1pMKu1orJJ63Gz7U
EUS2QHzMIkMxJwmRvW1nYjPDB9tx4RaS5RztM3/+4LEwrdq8nYSDElTXvRp9
EsXXs9yCDK152zx/c10tJSDNOj5q6pnn3pCP62HsIw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
JrWwPiomzGN7KaW2vFteVYvq9dwCvMOH2saGzEUnY3zVxhmaGvmOBmphJPJ6
2iBeBU7IOxaYtQoT5ZLLLLLzPM1qAR2rOIG+6A5pefmdjIhkv3u3H+c7i6Or
bWNOBZckLROyA9yWCPJxCmSpRT+9fS6JnKB82VlDQYUCVSv3V5fJjuBx1sbn
XcKHohSfF8KTvgMsmC4HHkSEDuyP5X9H3tH2Vg6eVKZN9IJDpcjPsUsr+H+x
ZCixmdQXNtOY/tDzEqTKmWEH0pV6EXkgDwdBxzU1IPBAfUICOufCB4FH5VSv
gb6aQ0G6/BdRBbJkuOlf0Z9CROhRZj2fwNSmVCvjLA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Uar7fzM1JqX7ZWfZzc1SGBu/qjVaEcgI5tnNyRw7MNsC3bxMdrURAzDcWpId
K2ZtrotmbjRWaAxKkY3D+4IAMlNtOdppxR/ZfEf+hUUalAbJ0AVKlIHtBAl9
mQpTA0ivxHYiROgaFmRdDlgA+XyrY8+VZCK5UF6RDIH7eSr/nLxyuUAF/MS9
qGgA6e/jIGhqLgDYp46Ey8X9Cbgwg+1SdlsMPKPRMRBD2uyPRUlUqRpRbqU0
IlRaLjegIAZr2R0HOfa+bEUkXbffiNGnusN9or3E13XiQL3QJKUdODkkBECb
7lSEwnu+q97w4dodtbWSUJ3M42PsnBj8BRBIE1vcfw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
sC2PYRm9Zea5g7zVDnsUGYrhrad1yE+lolRAKVkwG6dhyNmAp7CzpOf/it12
q+rO/rFifAo4SVcvYStGMattKJG7e4HLcnP8njySzn9nR4Nr6a4rt+bh68kv
7QBHCGbl5aq3H3tkApu5+f6XXt5sWlLKu/QPaYF2F5TGUsDXJJM=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
JwbjKlvhrn9mPMk4xAqyUDU1n64wBCOG6Ao+ySeMvvU+SZb2P1P+7cmgA9lr
iXYOh/Yf4jWZgDPhLc4PizsV5N60Wlwpfv+v0Y+2WMiA7xsiIjqEn2yhzAgZ
Pe2nGDXE1CV+e+IPWl5W+OtQLAZelJirN6xZ8V8PkDCtgq/DY0y2ki6YDhyv
xiCMrJxYZMhWAuWdAflN+Hc2Bgofa0NN1Uvxds/UV90uUwYo0j8dj4RbzB4K
jPBUb/9tcjAtmrxAklVLmF/sdfCh2SCXyzIbwQij0yOX5PdG7MWN2v/NZDgQ
NKpIzx0FFzM8tkbjtcrpa2V82kHk8Ou0hElXxtilVq8N3Y7YwFcrZcmeYqa7
hHwIWBzpt9trJ2xo34DRMZj0sxsxlHOdb/OAToMUjdfxVJXl86aTndATAm3K
YM+xDzimkTurGXdq9wNfXXxUxHy/tIVn1/VjvBdWJkiMt2sTDiuibR69faCY
w2dZ2HkGq9MPiCTujRXhyGAygLkigG3k


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Lh1x1iKq25CXNSUiYu16+Et3E0hJXKAkZgT0YoN7Zxoj/+ZqE5sGYl7tqm1M
BY2UMN5RURqzr74V1VCtwffpjGWSj0iI1mABodoHUKa+1jEy6aAoJY1pcVy1
qg3HUTzyFDhRPfvl9DkrfKHbLgg7Mt9PymnXo12EOhLJXsT/ajY=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Ho1HcuKvjTsv2FRxfE4gXCWxT4mlHOT7ZiDppzQ6pnTxzbN8G+CO27TUW20R
zYuW9VngcQxiPM/zgzrmmG2HBgp3PVwRF600EtwL2Ugl8fCIyQOIwiF6aQqE
frcpruYgCHGG7/1VSeg+jfLJAUe2j+r48CKeJuSd35tIB0r7L0Q=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1984)
`pragma protect data_block
juTzBZ3RX54yQZDXria/I9F6nJrkbxSoljGZoS8uRfwr+xKMMAeHINSjcyiS
Hmo1D/ATu/nQuYABMmnrudgD7GkQKwRFK2BzGNL7TviuSrXyRjw+udJCxLbW
f7+jGu5xtCo09EzYsPPpX49qpiTN6KsGfSH9SeEVYvQHuJiWdDxoPY4CkXO4
DjfwKsKqzipwPvvcTIYwJgLVRXHAVKRVRh7AhabIDEJmeov3saE+GVzB0MfN
b/Qu5+Rsgl8BWfjrN3IHGlk6TQben6U9jPT4XAcW++7R9Hj2VBmnXM13YOjk
1+c7O7Li9ltAfYzvLMxSV4rOXjEoWGMAr05xEuxRKIIzHWxLjjHZoc6TajLd
uYnXUdNAywGn5oTptqqPlxJAtVD7vqDcIuujNOW5KhzpKBwoMT6o06pJIiwn
C9EWpkc9M3m2K/1IWWx37O1LKigqBkuI06i5dDSj2n9pnYvnCHtRBqIe6lCI
NnWsi33GIioghBM+h1Jk6/vEyVlkmK3/yXF9IxsjzJlg26Wb+unDbsA1fiSz
l7s4JWjr5MbCZC3s7x3uMQU06QcrcnLvjzYVCmI+8eMo6UWJbfCbKKjQx6oa
X+XD34QDspPFGO98/jWJ6bp/yABuud33YETkjDktKClmxjlDH4kyG0gKNZVU
4rBlaqaJS96kwHHghr+DfDfjfyJ/gh2zpllfw3J54jDsu0VzbULQxV4spERR
VZ5VK+ymKsVryuLPfiEpyHvy+l0Z5J8uWkkzULSoBHksHr4Iy281aTgclZhW
RwiMYSzvw9R2deP0UWBPzsJmbG9Kui0OPrk9KBRhbWm845BIgqH7EmPSzUfG
87N9a/8f3FxULnU9eiR0jeknMRbz+cidvntX6PSk8+cvxOjXIY4o1Ct/mWOk
7eZNTO1VDoWvd7Fx8f2uOqDzg9gU80IYXPRLnYwTO4DqSS6os86VZmQ8Pb07
DtH9EgWwTkslYjiSOuApULSTP1u1b0jK/I8BTIrxd6mRRhNJya+9DfwQtv0Y
fSoszwBrYpONDqDgr8NE1tiBQCUnj9bbiuphrbQQfKuHTtUoveBxnSidSXzo
YO6I1Wpj1JsXGgLqKjDIFawqO0uW3xBgYhwrj6AjR1vUzPIa/z3maA487OXx
FQuWyT2ORP+HMkPaZ7Qo10MowOFPo0iOPgAFySHCxbB/CSGSu18iSm6115cc
TxsEDgEWTlE6ZjCEFbGC67TWWIMrZskgGB8/A/Sj+N9wgrBecmhBiTFASm7g
hdo4d5cQG96Vpa0zWeZcfi9eQ2L8mKiH093Q8YHkn9J9o6vZ3txquqDfDJcW
B8K/nEUWeBKs2vJO4N6UW/o0wrepGJuiiP3W3DDjA/zuOmruwM68HKC0+Pue
FhF5ZMmCiFwiAR67bAg2DuHAV2O35VDPphBsVLo6n4+jgv93misZLUs8k2xs
nRfW4OaWbiczuQ8aQ0whLKvycO0kmI1sA+0d0KYN8lHugsNmwlCT4v18AiBu
kF63ypKZZahh9kHxepaGdUxpvSzqPIM6TybTBJS+0C/pVaOsYKOCPCqwN1Vw
XRcm7PKrmtMLnidBFz9M3tp7PYoB7TVL6gBAHxCEGmvcSKQpJgn/3ojGzGl9
CK18+Upv7jFZjunlUYTHLLERHf7HtbbH1eqAXp+kuQRfioAStAxJPB71aolB
nwzl5w555hMpZK393OhEnnxJQbohZ62j0UF56eyZrcQ0SKzoBCfx/EDASIku
Ub4aKrZ39wFIN3A4BQVemXHXqssRkiT8mRxVIaDwYIz/vaDK64Lc8urEgFGf
qSfzOtuFUv4uCxGN42h3VW5DdpC2en/BTO8PieL1WpA8q8tiPedCQ8xb7ZIs
rICjOxm7wZVkU5qTyopt0YH1/w3whTwMUIqH0/nfQP+FI9bQuEZOqTOb+Hy2
w/Vc7kFdvLqRYR7Vtjq8kJffMbzjX97tPaUCa59DMLdMco180JWf688qV1Uu
uJWvpAat0+slQhHdpkZxPvgafr2wx68LTvJT0Ah9Bt2dAPgi5Z5ibMZP2dtN
pb3HBuOHDy0O/FyTUaITRz2+vkBhodCy9Cn2Sy1kQ54FcZ2EnjRWORsIawe4
X5YvLWEPSAp6BgX0HLB5DIb9b5JtkYfM8YQjVAS8rUcSrsqq0Ec/2rC6UJBw
BrzI362KWx5p1ezdTMZCJiy7WV5weATTq62nW8rzFsk7TOOfGULanU0ShEEr
hrLbXx/pB6yj+eVE5fQAcMTtuHvjvdRTEswrfrk2o/UII3FQ4iGypqdqbsBw
mXUP/xoq28oCpK0Hj/uGRYUDFFxPHwWgUpwnwJgjHrM22B1ytRymJYDXB/G3
fc7J/rimv/bJvMLZZv/O6Y3Go9HSgmJQ/Z4rxfp217eWEXeqgTJ/L1eiPqMz
E0dEDf4jj8Cx5gzt8LwVp0JeKY+seaXmwjn9ZeNyfyKi5LUCXTErEr35oua5
IHVLcsLtHH/1EbYNkGN1mF/pjTXjlubf8OX7KzsSQvSUeKepREOnvTWykxsv
WqDmGaKpgnUsJx5m23JbQPQLmjJmOGNPJ4AZz+JC+LLwMa6ZrzZXu9CDoVjL
3n5QOUO30kLVZ1hRGHkXWu8qNQrQPpbkTJzvB09f5l73wnWLQgmX+9/0KNTy
aTZ03g==

`pragma protect end_protected
