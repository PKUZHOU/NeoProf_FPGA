// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
hs+Om/SQd0djaQXdsaYI3o67TPDUjIioy8z9vtMLWksYJvo4gXyrmbU63+aFU3GBUS1m4iClKNMz
O2rVCyT+rEfo8kTjDlNMK/7gevGT0sjy2CYuHQygVUrimWTyJM7LMiwNSMroMyqp1YmaT8tqRu9f
/hqBeUf8D0tuTD0rYTkRewTRPzbafR4eSCphBUZceqWJqbm5O/ry7aQ+VVsVgP90nr5JGbo6Rr61
Jd0TBEQpmUT0V/NkLPfmrvB8FDGitD7SAFDmbORzqHh8tRVPRjQHpS8E72yuNzTeFea5Lj+zjLta
V0iGtjsqooHHxu8REm4q+oUk8Kqb/Asu/oE3gQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 4608)
01xgJsiGLbhDbO4lHFK9z45E3MbJ1i+zYGbZAYPMQWkUuFK54nPe2LOAuUqAJKzKE9+7evuxIxID
3OOhuK/O8XcWNTvkP5T9KuOwpCLSKW2yDloing8X6XyAQlAo9CcZNMpMI6ivtsszWaBOGbZVthsj
Q1sbZAhXVwyhA7Cwfo03IGrisk9pgwYm2fftfjnufEiW8Iez42Owzbgp2YiAWmH+2LgiXJ9Chu0K
E37NRYLQxEUesdhFsjbzSNceCJmffRprKzJWAkAKz5p4cQtDJlwm13nClrmMaAV8Oi8fky+o59Ge
jCSmPwfiHJ72Ha5WXgzF0c4Xu5NAnPbWw1z+guOD5CxtTW5J821O94cn7bhNlqmfcTptty1OAhjp
Z60KHHNe82XOFixp7HL+8sLPc1zq2kl3HYH6FsAJcI9SAal21gPdnWfHWbt70Wjzgy/fosdQXdCn
hfqnlmtryb/n24ctQS+fZZbibED46GexO7omH9tVEULfleG+JorktOQBmjqabz8LLQoP60ZuDhSd
/dEnvYFbuISzauqSYEgFma0PbkFXI1bpfi5gxHi1Ns5tfFhJ0h4vIjbUcdoziBP0Cx1S31dz1JPM
BXhMVKlRITQnNvyBaHbtla+wviiwKVZIF1SsSDqCxr3FTEpQOFtrp4w7SEleMS//wm9ANVQQv41h
Cd9gR5LPdqmQU9RCYmLKIeGEribdAQfuLLsJ3ACzGL1ZpA2pkQE5U1O9phGp0gE9p1J7CRhZybTn
LJpMuy6gcU8HuNYvWuwYqcGoDJIput/okAlSK7ThEtl7AxfjN9RjiLK8HStQrRjuQcwDeOqq7mDY
oLFN507pKrEJELOrJ2z+Pa+wKh5yQb0PCPjg/N50i9ksLZfUFbQO3ya1IjdFB72GjUiVMsOha9uW
RpiqvVFyAPJnqkUNspCa5GgJpsq45mfPnAZ4+rtJs7OZ7B7Wo8UsNzyYdqhIZz6ah+td/MlOFeag
OYEqL4fItMQYIL1sAm32MoN3gTTa1PwNEgRpu5aevm7HkY6IFg3F5AFIaS1gcRuLuZ0Vp86Koroz
wdmpuIAG67PKpIgRzp7lNUO3unZvWDAWgCp16VPjsGrE6uEOzWqKw8MjkY5bdsVFtyKspC5YlAkg
AiNNM56jq5Fmi0i09fvWSYWB18nJRcBqJuvPJxsFnr98FGJJRLPcOvI40J5UAeR422L+bRmThJk7
o9j0yOoDx72R6KmY2HxvcnsFP14FRxCF+QCSsqZZRVtXd6Lw9z5Cnmnhn02THExAy2B6egtKSq6w
QnqN6yKlKwfJvVjb1aM8gp/3K4xHNye2+rukscjsnnN6fgOAc3NMrUtbDd2So8MvbwZDwmK2aqTZ
VsLsu4M1iKdUGeDjq/M4nX+ye/cN8geHiuG/7k5oI/TdK0kRcfCKkSPt4LrNavYdfw6mtyKeaYH3
286/wr+V/m6dmrKWNWzW2PC4s5QnuKJOUJT9rTtLyvtyuXzlSt/fMG0Mv7NwLiU1AL1kpqmDC2pN
12C4Ldq56AMGuw9yWtX1FbSUq4jggZLPQbY3w7kF7xvh6DpiO5GMqrC0k/FBqYTttYI50e3ZGr9d
mMlXRwddi82ilr81Wx92gGV3pyqondA57OoXK+9nvRheLy/PdU+ZI7KvltpaWlkUx8d01IOoyyx5
ozww7ZtDxZOx0MmbyTh6D8qg9q11EZc4uSTiccgCbESPxCnBYIkB2++N28NQRJREDULo9PqYTa39
67xWCQXqoTHXJ593AgHeB7rzo5Z8WjmqlRjgOzsgXNubx7MNR0qEfDR+6Wm/vj51N5pjnVIy59Ui
nW27sR70jM6G6tX4m+rN9HQzqg0dA3UMGB9Hk3ook2hgdG5os+agQmAqS5VQ8fAXTC6od7FUOLBc
HtajbMBIe1KRqh9ipeZTwJCF0r6BGBjJyjDfWAMu5jLoBXs34h03FrxAsCLWLuds2LBv4pEtR3Z2
NJI/YQkKP1YbHWkrj8cjnZV8YS2gReaY5MKTc9eMkDEV4wDR52sNipEmrp28vVETu5IB4CPixHop
XyN0NsQkeGjuJkol1yzskzhdQkNp7r5v/On1pakDvmOT/6r6THZ7VzjJZd5S/WRMiAifjIQv44TY
MB14xB9WUtPSxyVPKWi+p1uvK/aVzvxxcrcx+xh1ZONJu5RO0S0UTaZPyiWzZBXbdw6bJ4H6RRET
Kbf6CYjjYndjEDlZRPAF3z8la7/WfijKBuSH73V/qrBduQocYhJ1fIok9ZBhFctvUVgOXOjtVE18
9LHVgRKrkFfp/6RY3Il/k9yzB32c3FPS34zkKw7wxu+W2XU7Gjb4nXy808epCdwvtUM5myw/T23I
JiUzldxUxnIapusFQQDniW3pW1X+fbXoZcVmZ9LONHuorulTxFEoZYniQyg55UCXdDeAb8H+HXDi
bsbuYLhQgcOtZyMkp6HeFAsOvDVdhVPzgZy5SG2D2+iu4TqXeOT/cebHfUnBrRWX8fr3a6b0Oief
rWkfyWXGHq5WxQQTJQUxf6WmnUyEgC1YQ4T+3Y6bRjaYKJOIiIah6fwx6Onx8lac8LjBYOb+ChNa
q9C5UtTkawgM9+RTXuFjemKfv5XhLH+nDJXcGviYY+sOtmS0/rhG/Fo+K7W2vQwKBEB9Pp9tvZHn
JMTgiZa5KK0g937+CHkWQl563hR6/Tux/q38aAdHoK/EgQiW8GCooXSdDCzVVlCpwgQlEByjToB/
hzddNqMq/u58URpJ5elGhyBXktK/Y10bUGKWqBnFXrp8gc/9ISTqWEYcbCG/ORj5cvvVs4t43fhl
Y2Ct2RS+qistQrhB3G7NG/8nwDjkJX5eZJ7NZjv9E/R57sDj2qeuDI4G5OIwJ4djuNvc34ZQqvmy
XJK1FPKky1UbQ8sssoBYZJJiK0xgHau1p0gmdLn54eQTRQLNx6ORP1gK1QiGJ76pXmGnN09B+TsK
masJNoqJN3WzGhItCifykOwRqMyOci7vsZTxXBMsp7q59fqk7CuCVpYNLxsvzDkbu9QvXRw2/ZSy
ryhKi5ZELaVeAa7zVA435EYIs9se6jJnMTx9r2J14CED6KBjixaykxKkBeyIxcC4smSlhd003ijm
1Gm7OAnijGqq/FFjGcf5PhUNwUxIm4PISMSrvHjkwOitJozt0m9TJusr6Dx5bMARvMySh1DBZM42
G3O64dGmveQ8M4t3pB9uIlpYTQuueA1nW8qrJQIbqReaU8GvSXqw8J9VZ/vh91FBlEhYasXz2NpJ
eqLJK9WqdfqWn6RUeFk02iQB3islY9AxGzeJhhTnTHGs5loYPGosTshUiVC+QoXFOcOuPlMJy3un
fClSM3RQDBNKyght3fwUy0Fynez9xZqaD2DmWF5a96ywjNnJ+3qlzcbleYyZT9UVyjPy2R/yCDgv
B7TxAzvat2nri1yu0l8R1VlooSMjPCOrSoYuReumCfjA9Fx1Uhd4dKiWKOVwwKlknQt+tacx0xRy
RXnkv7PGAl9yMqLrZzlx6sZzMWwPUckFCBDis6rWiYaiht1nj9CagCXOkrft5XeV9bU2jPwK5PZk
VVmUu6ezzrD2QPU1hwipoHHKGNxIQnG8hIr9zSo3U/9/e9cS6DtvqUM191lp4h3NJPQXw7xvMlpS
MSpbFJxCThzZ2ROTCHrWqTd7Ar4hfe3I1PaQ6VnFEi+HtTiUyV0whoNz4ryVTmK2ZkGo3hlB3waA
OcfUvkrc7YgITBjKb1JZwhxNfsysCwPe7Y3b8xdZIU9LI1UPW1A968RB24EfUoXBQCh1d7JzexQ7
+zCqZa5pZuIlvufgpKOiDp2T3c94t+F3ji86UuD3U+sGblhhiDZPy/xI4DwOIRpuJkdriAFCyoYL
Usx6LCM1uOK+42gVix13UiPUTc2U5MhBpLI0ynvfLN3JenKHYKc6fTDDP2Ptt+noeux5wEiU5se5
pA5wvp8PXPOiq8evsciOxlVQPu7TBz8VNvDSRwJi0CU1/N9AAyOv1MvA6Zj/WpWqmAUYIlL67V/P
cJdkFDxvgMHt8DINU/p/px0qs/oNv3xB3oesuihr629ZU/koPQxcEHYS6JOm7hbpBciriBS7psPT
PoW3J6KADjUoxmztMgBQWXrOwJHC2q4SIth4VCu/KzbDqtqLGUzMSy2qqnoCUhZi771vf+c/Q3QL
k6X7Q324gkhafTdtcxZ7T+CApsuCdMuf1XWsFZlhuNW2S9DbMBUhbEHDOOOh46o1JlQeRnn07TgL
lo2AtTXM7l/s6UyOwLfWfdHk8Yt9Ci1ePtCsDGsfFdGpPIwoDWVzzzc+GdDROZKVr8+gp803p8iY
JSEm75MPs0mGdKUi5FPkWNA2ZDB/Z7al2pRscqSyZDcJB8c53xAHNwDcwNg68I6oS8u42jdYPaxw
hvgii7Sfwjy22f7/2/7vjcSP+35rOFi+UFcii3lK+ow0s1IWK5lxygZpizcmxqcM9B93hu+TWoQa
HlFKOvfBsj39WJhGsyXualRpJqA1WtIZiUQAB7w9Z8IuSsulJOBKPNF9m+TuC3fR7irI2LWa/uIj
Nz7lWr8GuDzSVFDv55Bv793HvWDUm44URbw/1A49m+p56sdbFmJYNY/B2lXNkFtvqo0/6exi6bw1
Uqk7dib7+YeEkofFvic8QOcVXYgM4Xh953gXaTTNrvVmMtXoDkRs0bDU2gXiik7eRSQ4upFKXbGz
LofpX+KNpVLwpJ6jKVfV2VUFKLaC3/8jOcQIqDh7mnCmUnCcLWRd1qTbqgq3yOhbeFDU2TMN1xyx
LfJv8wFyGEDkLFuuP3/ktkxTvcmbi9R2rZofz/GeYvxTKLgNjNf4I4SWtjWryFrIAe6F+67ujMz7
N5pIPK48uUm7e1MUoPI2EJ+5uf6y45BzmOWhRZP9759uo0it9Lk6hXKNpfsPolKIAQdMyf7DQSnS
nLy5KP9BH8CD30d2/mJA5ovkaGTqGyYtaQh+ucjwo8fUs8UncmTztvqbKhyifxIQnNwNdYtD96mG
6K71DiWFmKhbo70ehOFFbXyyqEbLIy1K7GwQOBfh59lJ+skbCGPEoyaW07Eah0f15W6/LD3P337o
HGLLGu8zYrfAiMPTdBdWf1C0BuKZLGP5DvThGEuPcrla7ULZvTpFaS00s9Lvp3GoS6Svi/Y0tRyW
AtCafsafoUyegfbULmVRWCjbFsRhqsmmzvfOjjXb4jFClTviCXQzgc13YoXyPNJCAK5rvZHLlNMy
M19G7Y47rjrd1mnEUBndQlChy3o5qmU9deMgWIOneLEQGCuYEVwZ2l503uF1yCefqoHL+Dhi66a7
TGAG66F4r+WTH3/7RrNUHzwAIQbnAKbNqY0hw0rVZyMlBnMRTrLnAoH/+OWjUCxWPIBB6aFIAS3o
w2Af+FK19AbVdVVOhzGBAG9dqyFypjT02uPTT0Kt5C8N86AQ78vR37jYYlr+Si727a1M9SdLYUP9
m6+dfBUnNnZYwF0/Ve3JIuttFLe+f15VoZBf7GAhutErTY60oacBr6fSnKzwzitxWJ7DYF6/wSDb
QEvFRDqSgQFgw8qmMlxLwMO0S3n2GdSwRN6OaBcC/vhXeisLyin0u4TtWmD23mZt/t7YDpHPu4Hm
++8CStzIJlRJ2IsUFJNYBWKjptKXdxLIv6CbOmXPDZ0uAU/2f4pbgyi/uXgxEoLVdv3g//mf4d29
FVEBlObewyHhJkTpmajYaLdqwGisPGSzq2b9vVzVMrd9ZvyaVHlGZHnB+OdaZ/Jn2ihIZFI51+yM
6pPKO8strvFxkfIZzWGNBXaYHmxsowdbX03BphflsJCpDjNz22aQf8j7l4a65kpArcTDGTVuQj7a
XFL12IjIAFnewXciLbiHyO5jRHFs1U+qCduvJBsAaAzMzJKid7y3LrnKLtZ/HMoRE5ZJYC6aihtt
l4p2Etebr+Oc04WIeBM9MZmfFdGJfUEJ/LsAxbxiBLGJ3+0t9yc+0AoP+f4tusRWcO77uoWNu/Lq
l8mXE5kHxUf+scom3T5ApJ5BRiX87T0FifTfDKLwwHkrp7ompBvwV+sJbVX0B6axy1T3Y+zvucVt
mBZfXeq6NrxXfcbT68CfE5bMSi4h8xiU6vQv/QgV0a1uIJXEARh9TG2ZEKo/EbAp
`pragma protect end_protected
