// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
IA1Hn5YboUutfPe5daV+mDPzI7pzNwwmRR2UVHUTqp9MvWva135ujqmvsOm4
KJczHKFetEE/Xej/e6Tr8QqYB+7wR8HYVQD3EooVNsy6H3LMPXMg2rgtHvL0
P1/zuP0N+05jLu4AZ+kmeOHIwIFDV7Cf/lIubCtxehbc6cf/Jaa80JHWRBfQ
uw7wXk6cOXb/Gqu6hSkS+1OYPF5GJEiWqPubjqyVIRf9Mm9uuG/QeNjoJUVH
H1Mw4y/aLne2+u2r2PLi2md1i3J3nOvLmstwHz3O473WOUuJ1pNIe7GH/RI1
VhCCls1yVS3t7vKHyYUFkN3kdoY/62sEdeHN1rdlZg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
o4GNP14+nsaEwV4GSupj791Htx3mUaujB09dqCIaig1a6KuLHHGw4y8CepYa
gbwMWL7970mhqHq90MKoVXAaRuVdilgpLzaP37Eh1EkBEcEglH3QKJMxiELI
vrFGtYfi4UgltEf9k8QkSjnYlROA6DmX9c5tX0jO+8tMF0zcJ9UAX4m2bzt3
YsL2vKolqnA3/FIC1lpAnyvHAxs1okRpd1G+EdCf3QDrrlZRiwGM7kTsjAyG
/0fJfzJaigzjLk383DJ+fF0hnGVM+3HJmL9DRVSKkQN9A/fLn465XZ6AGuuT
uamy8SCrZZn/dofqTuGdrygpg9HTOgRW5VDhI/OkAA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
THJlvjPjMM4m/pOqihyEtgvkD22BerOVcfCvFchK2jQfAAAGXxsh0l0slFm5
7d63Pzqj3+OAJmFyyyb5SRdpyJgzckp+xwxmz1QE9bqDZFbjgoYib2lz0SUW
F55+KHFq7dgqDthi2DUD4YpS1vQPNqKUp1AnB/tSNNSNpbe53TyU0DEdKV5X
Z1mfj88x+CeXDISxcK4bsVgyb6wb4Vq9i1Rx1QS90brYvMZ+nwXT2oDE2ejd
Y3IaH1ZGejzdK2ynbDbeMvAcYNXj9F0fG/F7xBN9CyP/BQRvt1Wh6u9tvXPg
OSGIPbnwAaalbvBQgKUtCr4QlLRn6F6T2Aiz1ueA5g==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Q06oPM65YIen/ywo4JlvHo3AcRs8vU0a15o8zO+8MXxOkB/xTdlSlzu35zLK
1wkpkKn+ZOU9wToI3yngvr3RiGpiCUjcZZoGMEdazP8FJzlwM4rJuW+iLrtx
qVTIL7rSRd87Rwi5hCxs+DH2cyZP0FMHnSLZsRenv4XCQZdC0S0=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
WjP1XwX+bjQ60tLaaRRX9aIj12Ir7PCPjivsLuN7ZSH9w/Wy/y77GzjSu5N9
f2gDeXOy+oges8MIoeggKkDxjMKpa7FGX+15IQTPEWgiODnZZqP7FIofrPRF
qrwGL0g+o464RS+Jj7VAutzTkzJW/YoCrFHUkQS6+MLw6V+Dvhs716J/xbLZ
EKjjum98kNC2Au61cD2jjOsx4ImrE2kxMxpcg4ZVjabZ1rNRjQHtJOap3OI8
CAM4mlbZH1mOxWs24IWESuqz5tPCffp80i9gOc/bJ8QK3vvtFYO2cNF9kGO3
5ajz2C72YaocI6dx0VnwjusX1pdI102FTlXuMPAytWVwO/o3d8z3uolfWLg6
jWOY7VtRwFDdK/7vmT1hF87KyJn5O1v2g+kz0KiGyAmVkXxXz61Xk7t2+/F0
aIE31Gj2nWwOnvAo1+Ras056NQr2j7XKUpZOsyhtXV8lIQfE5k27d83F1upA
ZTG0QYGrUi9bElhWZnUxfQ76FATo7SbA


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
BSQ2R2yMvVp8RQksSBBTj72HpxeiJJQxqv1kIAfurJN8rQqN5UVWEcpyJgv2
mduNr1VlkUXN37h/5qOknMTOaSrCvuANsmAPDzf+1Dg/EN0yZD90vmNi14nc
XKga4vsYgtYLaEmX1dDoDUmTEfsteNKNoGOtk7KnmSPG8G1HqH4=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
O+uf13OzNK/ezXGRA4bAmqmGmgYOceGFioqGD1yjhVfRYQymi9yfGr8UkHbv
XBUljyG8vQWyaYLpewJMRFmZIvnkzC3+wD4S26S+wZyEqVw0Biy1upX3BH7C
a0MjlmeufEkXwFyUR7oaWjRm8kXDD+jSlOv1kmW5WCFAEE06Rxc=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 15344)
`pragma protect data_block
tktZtucdcBSPAObGHpvq5RPLEdfrdjjuC7VjyOFOWXEWO5hn1xWvwWLu+gWt
fZ175O3ZwzM5vHOR20vdi0tTZGy2d+X1HGB51EqY5TV94zQTuV5BAONAF4iq
edJZu26Mb1+qrI3Hf9c5C48RGHQQfzl2mvey6hgPy+GBL6azpDHvrboj+S2I
5rN3FWuX8lBPt9Ox1dbLweHFpTXMc0IfDHgadr9jcj8A8gkD9Jrw8nLHCPVG
7pRkmIgUltIz55N3PpRPnw2siFvEYfwLHRH91KNqoRgpv12+mtx2x74pGLkt
UOVqTS6VhsWxbyT35WVV31nkzsQQ5Rs3v7XxofUgIWF1Cm3qTCnEcfDCJFEU
mS4Rb8MLIrMA38gqrS0lFcDCRUIrKdih0nVQbYCChJg6th1Cl0ypzLxIxIaz
eFPs8nqCOQ5oUf3uXweCHQHWwobD0/Fsz7neTo3jknnM0x6UGdy3/ziGxNbj
g+K+h9hLIKMZPBdx6FsZ8VqcDDtT1qi5Dr2pwB6j1jYtlqvZyrQ0Eile/Vpr
jr0gt7zIQodo+UMBoTuoZW3QCyD+1UTuqx1/9o4GNaZdVyqDcmMyeJj6HtGV
DyDbVErG+M7LGHxDGz4QsCw5UD/KqoW1DGsWB+70iEqOA56aytIB+skwetc/
Kd70qQuSErWCq9LDo0KyVWQlIcZ6t6N9i0p4XOPXvzYPNdYoariQXJukUsLE
/vVn2AxX7LLL7GRFq9NmIuG+pwJ/xUVOnzFmHRPKnIvXv+glBM9a8Db87184
q5KbEruLO7kiP78667KagNiinbMzdc0FHaY4sF4nV2di/pxiTG62SczvRU7R
en35QG/8GvtpEaiJDrBXbmQN3yghrOEykPgnIr3lFfhmarbKZE3E1tmOgFp9
uXTbjzAjfdCWDiaD3t1BXwQIzr4nH++BIFKYrCU0dnlQogN/IkwRgTO0xe2W
pQVpcGrUAhP8fJwfPgbR1WVFZFy+O293DFs7kWNG9hdYJLS2LJkrVki2QxqS
93u1q0iMMpORVrN82sCtAEpSTFE+olnYDlhwgbOFhN4gngeKIpQ86zpxbVE5
aWq9TxPp5sC9lv+mYL7TUJWWP0QVu+wGRQrUcZZ6jVd0GjYHqcOFnzAlHDga
adIeMDjgWAYyXL6EYSDwgVviWaMDRZy/tuXWG9MvGgASViYI4zR2vL0NlIi+
mDFoIRdaY8t23LpPT3eDeTQWRGGLdaUKjV6QQw0QNl/z6iUCuQLCrKEinLwt
4Oc/jlNRyCmt43vgR+/EEay/bFFKHXdFPRfwxaVwXei+P021laB9160WRPxH
urnHLAxzEi95+y2ePfU81UVZJym89u3dcFu/10Y9+EGjNetgqasnb5BaQymn
2mgoXxjlVaCFCb01vBjy98kfCpLZKPxCBBbMClt6YalbdDpfjVJCdCB4TCjp
ik1n8FmefIR6lv2nED/taOZ/+nQ/BfmOmc+Duzr/W/6w5d05B6LcZHVTXqV6
NbSH+7cksCKu8QsNtWOeS3DCR+eq0BLpIxyDvZ/2RHuLEN+GIkjRwwYEKr8x
54ReBxjyKkN6BHG3KcDo30nqFHD1RfecKskU+rY4ZKnI9wbJQUBOmo1Ay8oO
DeECTNEGVa8gc7Aj7L/vhEK+Ae7bqL6Ul41WRHMf9WTuSBGHibJZw+NpsT++
+eNH+8SPRx8maqdPybhBbiSiKIiJPwezZn5ae/eRIiqFDrImbOMLUzpLxPtx
xV4PEoox++rgI7E4sIcroIagm6KgQLYIC/NVHTh7h4s7E6i2YUcGHGrEH9s/
dch3zvp51bWn3uVarYNqUGkyrbUDQKW4i9o1rsNUurwu3UaNSBR0E3w7lbH0
QE/pDgkc6fIWVP7jw6fSPOqLux+uco5F1ntshi/EhoIPJ5x+8IgBiAwoE1ZA
4Md2DX2F+thvfsfs7Q8CaGU0n6PnMti4TYfHcyWCdaUDBIUV9YEg2QCTgzUe
ozuC+LglzkVJwiEvvXbns7sPnu9bjJJwqohpg7Zh9Z0L1Iw1ClLkFo41RFVH
025324koZ2OaqkwoN1uli3MY0o9uIdFuVuzpdinhxtFrxb1XRy0JHjg8TpVm
ko0QfeHdxwFKtkPY83lsXR7+5bv3Gj9XrhU/d6opyBfavLbh+WnRtWgMB9SC
V2Ralr5kwi8y7RjMFbkSnebWKHui1xt0b8FJHBhbeUcsov6HZbDfFsueh/JX
bCOMkXU7vxI3UGYGJPBokq9vTjN8NENUOMmMm/HBvhYydSy8Mdgb5tfN+8Fc
E9htz6n3FF3H2cUZxUFUu+mQg2dd8QJuXqsKgQGrZNqCvhRDQll/py32XwEO
Y7fKFaxILfUgHgNiwA7utH0KY7gJzp68TNJ5zHbtPr7YcuCKreuRGis3u5lX
3lshAQu6xrv3LjmlsmsiNFRSlb7Svybw2YaFUKs6j9skDevc6/pwz7dL8FlD
f77ahRK9ijDe6WoAG8I5XdwR4x7aOCsY7MREAE1qE7nFIOkstdHjO9JK0asF
TC3yzwdB+8i9xrDm+DEBDQ2258DIeXJe49MswRZuMn04TUCgECTR2nqu50Op
Rbvobt2lA3z0HMkA9Ob69lDWmLez1JvOqGu+uHGeuK644zBfLz29Czy6cH+C
v0L+wDyDUc5byYXhLiqsNbHzX5DkyyQSYI6KwqoTGFuW9W4ixUtt/nMSrggL
sYRN02bsxkw8BGFwhTC4AlK2Ap2tFZxylPizNnMxQplqNKzFUuVyaVXRKtoa
Idjxav5BB9X2dVOGxcLuVCkaxiwJqN/6ZrLklco7Fk6DGIeCcqExiw97ulXN
dsJjGIBu+3rzMcq+HhOsMEeNsT/QlZJZVB8YsCkgrkX5dNdQMOnUYG9SrKvj
+NuzW9/F3C7VAVN8yfFJJHtVSBj90paLDeEePsDHITJuoYB9HDnUW2RDVBuA
HQBUMJDdUmBJs6Qq8wrUG0zp5UW8OF4kfBZV6Ba998sbOFLpSvtXDqBPcpas
NIGX8rKijVfJ81g/e6vgSRmUOj4XaFBcEtXF9q0V57bgng0+Z0eSjmKuMSE3
Za73VzLnd+d/3a6hpHKUnEMFEdnyhgqu38JWfVgrYOrYbxHahvIJEfVdy9Pg
3o/g2EZ334lRNJReuxv/pGrzY40cvm6HLhMeHZBGT0QGjA36LStJ8mxsyWqN
OERV2rUkFHkMx4Cz+ffISF9QGri2KeDV5JfMtxMfAP35WbI/V6c8u3Xd/1XG
wHEANnY+xLvst9WWRaIXysCJfNsUpZL+wvCgy6/UMqYk6NiukRKIpduyAcc9
os5Rn55eLd/8bwBLGmMCyx6XFpPVIZFD5nZwXz9J352ZBZMmmEhVT8q9P3tf
qkH+wWD6wf0rKmzbWO5gQW7oR5s3SaHPPRpcksQYQT4Yxv+W2GtuRmW69c/m
27uv88lgLfyMhsIZRdgebTHvScmhNYxyQkzfIGxPpZ5GktoJZUV32QMCt9uo
+yN27q/qs1dmKujgM4Mvux5KhoW/GiMO5rvnZkML4XYNcVO7SmKp2eWMzQdh
J6dF7O9f/q7tNQ5oe3KkMHywHVFy0wIEWFwmbrAbLBr7EUbmMmheox8SjY4+
6QsDr121d+zCOcYqVkk/t52dc9xf0qTIsSSxmDXB+jSB/U3kXBPGua940+QF
dNa1YMzfrNI5USgstWhEkZh1Gr+x7Pa7oGwqPJimO1fNxT/8Ek0fqJsioWrV
LZk8KmSbXJJ6vzvlfDhv/tRyF7ZSuaY1etAIvaXwVzdfEXmvVticjGtgZxzK
z/zoWb+Bs7lF/8T9AN+pKKKMMKI6sflwKHdX8+dcMwjepO+ZDYDD7EUxoZOi
eB4+al+BU0CXXTG8emDX0XqFarut3XqSGTxBKyRQNLbkPBA4Jk/xHSAyNv++
EQ18W2auGg6yY6iwbO22uy7fCa5KS5dddfKK/SGPhp/fUxp8f6U5cdUAzwkV
OIYEhs4kwJKnGs67Ztj1aLTLuxA45VYld0mXlUeQYGCCBEcK9wWnloWQDYja
oAT5QT9vFPxX4IqziJreOrYLQlvlY6gxENSCGsrwzQE+SsZXBUYVZayPjDPJ
vYgw1uhZDZTx65VHwDU1rudkSD1PaWpc0iatJIpQlR8fJ9MglmmAM2FIatlP
f2OgA5OEqyw6hfjawrjlMxf0/egKzCzgVO5eyOUqWpL2UVs6NY3sdm7OSF7h
TWvwOQdxlMAfJ7koJWytmFSjYOagyOevjUG5kFehMCwZ5wAfgZS1kQo6FKaF
vQKXHE/1p7OPs7KFuROIfikq10j4lUpyC44AADb/MBN0EBkp0ZVvn+/tuQ/l
4r1sTmLgNhN6EU57MlCX9vr+xC4C+v5Gkbqz7KtX/9ZlV9xVtwyLzFGHlndZ
Z23Wd+SgdJcOU0RwzLeKy7Wv1gTg/0C3Q5AYqx1EnzQxQsJOzrn3oUMoQFHM
hSUpZ1QDWTy/g2odwB2t8t90aqbrf6FedQbIqYdRGqYnM2xzXS+kBFzZGT1h
cVJBqYYCe9uys1xWVFttG7d18CwOv/EdUjGztEpZi/Wb+N8CIbHa3kn6JGpx
fTrRGyljgtEyrjLHHuQDHm2X6oOdV3DqRmEdcwBZFOaOq+usM0z9zF5TneIk
pw57oquM9BcC3/inZ5Mh/Vzr5mkAAsM/ceJiy/0W4BO3y5RBTdELzZAWhgx6
4DmquX5Mii1CqUSuEuoFJJ+RSbJB8EeAMkJGfaKL5hg/vUtBdStZQCxOtd95
CspFtOaeaz9LAcsJX4L3yNpI8mUWlif3cBD7+pgrZBXrME5uK9kd5+NVwdsZ
hLK+Z0iX8g8rToqDiRf7VLxwblP/SXN3Nw2mEbJqUFeUmRHeWGqm1h03qA7/
iW2Svdq4KbjX5LWNOhnlExrzM5rpLrzPmuA9ZEcQwzyA9/1DIRyANLpW4VQw
IYfuiAOuULRQoJqeymw3uTAESwQ5wAFW9y58b1YKyspn48wAJRzCOrDDzZ7Q
LPFjAuIISB8LLJpGBLLCN7mbbr2SrvjqexGGrM2qAB3B78dG2r+cmk/zMGnC
E6uZgUDMjqFM5WgLFtV4bWIxz5RKki/do/fWGBUxhI7C845WFNiXRTM8+50N
6ALK7CjgiWlfx4d1lbb/iWd+eNx1wrWyvHLRvNqUUDT7PluBHSXYzCsg3fJ+
1Mx4bdmy2jp0zQFm28NlTt+9QWBfTbu2s0id9WsePl90DlBGUmQDx1DVM0lD
V0aeFNDMgYf886JS7ZQKFNmpEsyKGK9QAC7twNzm1g2OpeM+IKRDUerTXYIW
UyBYrk0JT1hy/ZO7JHNx55G5WYkmsnVOwfBEm/XyY+SixZU59jb9DFqoQhHz
jkcWp7JTtuOA+g7FNB7QVcyM7NtVLgbsXFzBnOOyXGUyBxYfylW2mKRcwYXM
7NRqQJWvf+V0+i+hOuBH3Clc3Q1c6NqTQQgcj1bX6t2WvSETI+yFHPMuWFG4
k+U3NdVGb19FNsnKgxooRTV65nqSaYQ8jnfwqC18w7bLM87pzs/6dWDGobPg
t/cxbTc9zcWjy3acWmuSUKHMhNF8bSaD9nabu3AMEaB3WM4mnQZcxlywFy9R
ZwRbsecJEzDF3D2Q9/5gxdSqv4I8X3hDPwxIK0jG5ul4RbryUOrm+cXQB9dP
myKcTp09JuZaqxeLK6wrP/1AlX6Pdr4LtISAKM2ae5iUNVRxX4Rk+TimMBJ8
DfbjRq0hVIIGf/IFeiXdW3FNJNYs2X3u6cSuDap4WDLNrFBgNAfHNtwkl4Ue
dMGh3k0WrQ2J0T3Gs49L/2KnIxMRqD2gIZKHqZ6tscOTlnabpHcEEIqG8ZU2
qWBIQt6rxzBj92K2eREtT50hRJWtYphfJcpfF8644jKTcxUTSX1h6OjmF5mh
oNaYi50fJOqYufFTv3L92mievljAXbQFJogK9BxOZ9fErLTbNbIFj8DgOnfG
nYKDEClzNUZ+EWyBQ+kBmIksSxXQFHZ84ouvhm8EjW8zHFtrC9TUEabDEnoZ
yNsEJNXIvSMHrYpi42iBTGFVwRR00Knd7LKhskuNueaiT3zBp8PFLU3J7Kfl
Fgk0RZSRbNs7qJdABIk9jLGk4o5KrSs3BmnMId/9csyYPTOPgCYoyF+XFopm
py83JySFI6CfYWAmOQjXTOREI+umzvZ8ZhZykF+3vE5mmphxmGlYyvtTx122
oBQ2CKGMMK54BSx177t2fy5WxyhiF6a4xka+tHyMl6f+G5lBQGTLiCy7cB05
romkINckhGtC4EJeN85Cih9g2afTrwC32AKZ0AHSJgq3hWZbUb5fBqUY1jsC
JOz1NblZrqTT/uo2uRLKYRKqPX49HoP8DX1o/Iipz4aiB/br63u6IMIQW3DZ
rpMfi5xPeqGSWvVFjLAynDkXEQ4uaIHDey2vAFuvvPQHeXEFtERXLvBOZIJ2
g0d7YDKJHvW5H5mbi+cY4YnAwQ5fjyyfWnqSZaCoMREqFpdpg7LnPasRf0HF
28+g5zSnVnP8GqHUsvBYoiWJfUixFhP9HGx7XVYgpk0iZbBszoWdTyqXaDxD
peNqtIl4US/7RhfBx0WS2MHMEALiQd1UKxbdWk9KSv/g6chPyhg5BnbtPb8k
ruGNvYsKIaMqiomJLBcoUIaMmZc88Oei4c8cfLd/zLCHuMFuyXr/ThuOJnPW
ugZLx3TL1t6xJGynoyaxxIXEz+IvF3/z5uLkGveWmze6c3VukqBFTWRv+Wsf
0Szz8fqvj1ozPzYRWRwLDD3GkBqc/jDtB3MGwEbboCtRlV2noau9QOexcakG
NXCmRHod59Lp/Cqz1LJ7zOuk9WkkIgmmDcUuErYlQrBm9qg96CeXhHTBahHR
6hBES5fxXChxGAqQMeZSu+1Sg09T24OzDGyCGe+KZNDRLAdw5yOFwqY9atGW
CteJIAM3BiUmwSVPZpqSxlAKBUSlP02lx3AH9wH7dqzXstYNBWmofxCqRku4
RorAu6fHW88h7zUsEjimKyERNm1pbmVc3x/qa4gUp3VHR0tpXUdwCHM3hi67
WiKc9/UXwrWSC8W8I+IalEjKXLrDGpFm4vOPotxn8WbvHZgWfPu7ZWJLx9Zt
Y1md29nFtB2QiV/KCmXKAZgztOlENwgMrbxXMT9NFWHiziUhPvyKsHb1jgR7
z+62Hp1hDOnQ1tysoPAxarsw/62DVnuZODymiUMchVuoJ12doIAtC6vLXcuh
TKduMSYBfxBspM2MoGhaVivIgDTk+4MDkgAk2Uv1McLZrLtYwHiSrmaHTtLF
XUaw/wM55PcfYz96HgenYRuv+1t6P/0tNXavZtl8lnnp6IJDn4fQBigyzjYF
VVwkLTyTYt/u+iHSPOWOA0nsZmDXssXCeDd12QCnFQX9gN6hTHslcjRMmxiX
QjV9AC7HU/GKcyU5UCLBhn2PTzSpZJIAwTJ5hqImty9AL91h0Ak8+zgupzHo
J0yHZze8nosQxeSqp0NBH9nyvMRVYmMiT/7teMc+UA2kJ684WCsVczJBjYEC
odBT9DYvHTwXa9JyE4OkcaAJg33Y0HrQzoF3A8mTWY/I+bim3ZMhwmEV9JkJ
K4Q0E9zeiJd/u5JF5mlU/8VfkZEOBZ59Y5qw6JIGQu+ar6z8WcGj9O3/HVVV
E9QoGNtbrg/bN2ETvx+sdGs5CIwhB+X0ZkhnYoA34C7z/XxEBzSwOrl4RPzt
UCQLuqlc4cVsMHzfLSA0WFBI2o2uTMdExqAjVlSFO8LR9pu/9/iMywGPB+ye
qpyX9YW/vBXZePU5JmWRTr//YgTl2n3oaYpns8BwnNJCNmjGxqfU8Zz+3H+5
QPFtGQOQEDUd1Qf6HZ2vrERauEM27IIPv/YzJhyOcQ3YePdz+CEwv3h82Fqm
/8yKdXPT1Tzn8oUFflRz0kXb3L7y8tDqemHaX6aZymv5AuRjdaXVR1DquJPk
5IjaqoP87Z+juDyH5phvW4Skmqrxdg5u+A8eamoGYNQJN9LZODTKOV0FfFAE
iGDs6lZmQPaRrBQfvgWleF3YdQKXSMdgaermfBhlh9Us5vJetHgR38fgRhCE
KxzY9+XoMjp5jERiGrvIlrlS0h+3if13OzoAX0cmkcytkH5DYsKMcJZVKDYO
eQFJSv2eCNxGikbNSX+F41TS9xEFzowKO3Zis547v4A3f1FRuIG6BfHmQlGv
HgcpFaHwtIlDOsIv6ZOzGuCBrW04cFdZovtOOQ6Sc/eZ8AzzlJQIDVRlfcKM
7+xol1ZPZxf2posAdmtpPHp6MEZYCEfnTbHaZ0aJNKxbUOq1MOxtJiWg0URm
N4JyEpymrZVpfSrSU095cJVBuPV31w6H3teCf921jrHpaEOYrEXWLxzfsTo5
MK/JRWUz1Q2dxhWEGAtm4zD+tznRXT6cGgTWu5KKZB/N59dlUXM/wWDfz0FW
L0P7+uvXxLw2ipzzoxob3higLvxyQYeMOZs72bUszJp3+FUPf883mE2AAIUq
SCt+SAKOkop8O52iE8WEqtSRP2454j/F3grL494nr9+e0FOENkltbYnBMQA1
FTIChXoxVidhGPCTfnsA37u19enNSxEq4/5MVA6sB75DFEUIg7iqCLHhzH5Q
LEGpcvOPBfUh9jBIYN7Tm97T9Bzh7TQ4o3+2v14OyFAtqMMb4r61vUH83OJv
Z6+eZdoIEtL6N4oxzx345JNsb6TVf1fl1ZZ9E/TL2Z/yM4RCQy3XHiOilMvj
nxKHGU5wyK2N0kFiB4kvR7uTL1oDXziiMatlkMqo+QNRByYQJ56PDXtESF6/
VLQxCbZL+HvsZIwYFAepGS3FxytaGDEptn1Xghb9SvVW2YlLpWsPO3VYlla4
trGfPtbLsp1netdhpwxPrYqjdHJUiDVBWy9oP/OPEnXL1B1xrAw4jnH6T6XN
vBe6xg4ww3T2q3kB8fxkGFYQCOm5zun8BFmKQaEBI+bOI2WFqTSf5ca/q0D/
QutM11UZlEqghlY2i9xkzQS+ygC8FNIK1w8r19GdzYGTXfxO5Pvr3ImMvWPn
AXBls1/xlwA61HYk52bMD5ZBUqXzIDiZ5CzZyYRpycQAAxSF+le04EeINpTB
kri3NCCW1hlAv+7A5INUi4E9TeaQLgtfrtY4n/qkQ82HViY+Sw5iQNTTQji7
mErW7b5yJywQX9Gk0jXyGYYbYGArk1V2gvRbVCbSXjhRCImW80RxN1Nwdrgw
KVCaXV21xg6ZcLBPAgelP2LTrWZAw67A0b3mirsUFa+O/yF3EIBrda9PXsm6
CoCKgDgfapn65JH1q8V3gCKnPjlnmRhJFpJ9aLZFk4+7xFa7MEUi4hke4iAN
3nXNbfWVOd5VnihJ05ldfMydr4zVYxu1jiUyhoQi6WzhOF3CVHMzBapVI2sQ
lvXItK+7rAeGrbl+wHs65JpSlu+NUWcZs+B1NDPWU5FAixRjfKxxy4rBqUu4
KFcaZTJtsgqkOobDhUWSjif4qiayorAjhl3POodcWpV7Ram4GCP/C0637fyC
2EWCRTf3yF7a+eBu/izqbd2VITM/oyyme9NqmbZl4a25mgajUe7GXmPvIJSw
DxiA4s1eOVGngnUK4VYt32zncyVoDZPNhTRUuejxlx1yb0aW1UKH2FVWyYv3
Nj0naDdWNDb/YbTb+x9/ypcHOa6yMx5CuuYF14DB0mJPOhz/ote/tgUb+lFg
DxftTcyeKAhF8zH2Kuz0r0QL+5HqbeM17GQHgh0xPcsB1bSNuD2OJZ2/kNjI
OVzWgDT/wwjwuQAampt2uBcd7zRogfvFyir0fakMhMaHcseM4MkSDGo+jhum
ns42yGCBgZKxANCEp+QGfkOc2HqEyu7HLuylP+lxeu9C59giBdXiA9U6IQRQ
RZ14hLWo/UgNxbkQGiUU6612R6epUo2649ZJVwSBAJlDk7tqlxQjOB5/VegG
ZNd7FsWpgxvYm5dcNhPzy4lGrS5mCNhi3FBo5NN/qsMhtSVgaItAgzL0Kf6b
tkOAC+0wAP8yxuNbBVdk76jxCGzVJb7lQrEQduiDyZ4HIZlGW54fKS8kdD9H
hUXhFITFcwrBkb6HY3hdQjbDqX/czt4sbWEly9ZmpdoqvtSlkcLz9xu/A3tc
yRcH1Fdk7i3zuzqyJQLZvMkgrP4uIhMn1F2P6tu32hBOsgpREk0G4bRZM7R1
1OJFJZijvMTSP/JYY1rKUe9nOyKOOZXYexV3TUuqUpDc+cp7nKXWgellr8Ko
LM6wnFdBKvT3mWgpex47CvjtGYNvNQVZ1Wfaxg8ChM+tJmTJ76eYB01AZxc6
CC3WjNr/WO/FF1YfDH5WPf0lCME+bEoX4fxx8OBSeaT5t/labma9q6/gjA6U
MWdhmRzn3XZP85vAvABJiPXou8GSt+Jxvz3kEu/kTOlgc7c8QrPyrP8j4Ms+
EZoq4CieHD3cnI5miSwJDg5Q19+1x8bWYkPCfxnNnQGhHJoD4Ii321RxYVqZ
p2sFx3fZXdNg4nQsdrNn96LMGWHLeAwpZ/2hTl90BB5ixg2Xim3m2ncx8wPJ
dQhUqTXjlpJk6KFCIrOdxI7IsQPOdCfs5zXP4evPzycL6N+OC64Oe2zYK5Wj
O8lro7YlyrzqoTD4LxwXh0663Fh6k9HB/PYLPPns2PahC0GFMOMJiacCTl3D
9sRX2OCHOvsAoEtDzba7ZLGN5+aNlhTzFz7f3UuVCa0m/zESvDHSfLPUqtbp
gXjZvm+7z/PZrFCvt8voK2Z+PKlahwBeWwjy/EzgptmtzRO3xpbSurMqjksK
sO+qzKHESFcyvA3k/bOV8/Dw7zO+EfAD2njc8hc14w4C3YKOaWEBFZA8laMf
m8o2F0sxyoWht6uRcvEX3FOvyqLb7rIhEMNWAgtZiT0HCu5n4nnoUeMFIXYt
BwwlXl86MO+JAFJhMChTSrmz+ggSkZDFlJnFsJGz2/gPHYuzUhasIAZzF2ls
Q+YTszks3n7hF3+aVsq3FIBYEboVwyUECWB+8u16i6RXW7fUl3ICt7HH9agv
dKXaF03UkjUhuZXFrAvnjmYv74ItxMH/C0FTSGFiU42T3GTqohb7T5HVqQH2
h5UauMd53vDLXPRvcP3hIAgdA8f4qVaaDm3Cpzxta8QLD0G0vhPKerZldUmj
e0NkuvHdRGb1ArV7HoC+8hA5ArewEA3RFI6JsHQtMlUQzvsDmnRn0frhf7vd
06WL23F6Z/bcDvcOh0L30aZKGb3235j4Z7RKCe/I4JMtf6e0eyFjQcBG/zYt
h5cFCeXdGs94JHgZkild8grQ954bd4A0pcfA9IIhRBeAn4daAL+8UmYJovMn
U/rYWnnwmrdD9t5U4KLiQhJRIG53CS1bk3wACd4iePxMen9BKCJnvR87aV/l
/gdnkwy3P6rgzQjHpVhmMVtzozKoQIlcFDKBz8lfDr6PqFXhf5jq/vXxkHBS
bVGRQPnEOQdU+/wFQ5YBUOYBNoyNsyRqQwaHdC9Qx/6V7YPbZQvAsaFHdS8r
BBfzn5EJV8wzs2jdT2E6nfqFj9q7SOVvoqdayCyHPzPrXCwxK2xFrKuof3f6
0GRB/xkea/GVum6Wt5BDN6FsVl4R7nFDrIpScBRj3wx3POd4mZq2wThYw0uS
iEsRb/dH8yFyYBfwOolMdZjeOJIBhaEp0MmO9A4thw8yB1RpskQYUw1l7IUL
2aitSpF1uUbUOF4h5hi5uTTZwarGUFsSPI2BmflOvZwUcYP9HGuCRoDzTM2X
o2nsxIYkDNH8AHHdg9rX6SfAbuPxOEgNgjNVaPEsO9ZXXH2Fr/MJutcr+Bz9
gVK8zR6yR2zW1dXBj1gBiJTUJ7R35rE6gphViW2gzfpBVui36VJuwD/1VU2p
z1SSbHSQzzy3ERy00Hnw8fSbA/0KWBfWSXNBoFOolnDpKJ2oUO8/3O6grpJT
wRdEBE5m2/+TJopRaLfA1FGK0oEG/ZtSQnIl3OOIMRmUTWNYB0lhfm8EvY7d
Lr50k1Yoa9wwLzvtEe36wm8MgjH7JOQ4KEFuQo2lYZW4PyaWeoloz4HdiMqi
sS7C5XyTF/v3/xF7I6b7HM3eoT6fCnnO8aXfQXi3ue324h0sUIeE+kJm38Co
exwVDP5/gymQ5LCGbqlslKnuyHkZrAsVZGW4JIR4eLGY84puO7ikp3kJnsZ4
6iNpA2hffTvxkaoDJg/FtDnj5FfeAaXmTFoBZwR4EDJ9WmrZU4S78TF9m2kM
KIEJSj6NohahF5wwUtHqYxcL2cbs0tl0zUpmqqLsrIwljK7kdCQ5xXIKlqIj
/kj0QAURPSx/v4HFDOb4mMkvg6VC/5J4Cjd3nO2NfWpImNMWSdePDU/hLPc2
mFeUZfghylQv566Bxbca39n+mhxFC1jYP4MaZVBUSCiVumerQT8SuS+gZBf1
JM6ZP64tUQrmU9U6lPk3ywixKZD+9K7PaYiwmyg0ez8ml3P3LunWDS0/bYL5
0BRXOvNZCriM56HKdL0XGz09or4iAJQCLgMsa3puQ73YCfBV/4FvKUNpVDLG
1W1ZlIu332oc0OUM8yAUXpemlpXY9cO+56xNX4zHcvbTiaFrzrnPur/gPBW1
K0W8cNgVXraWlSly2M4qwzxRpucqmrviDrPXO0GkvCafpsKMIRkm+LPV147j
w8fagQiH0uYK5CNFy2u3MilYxuOQUVWoti7Lfias6br5SYrBPibGGI9IDjF+
OxdETrxNecXkqxl+0dMKe7oGLMimyBt1jxETou6wZu+Zyfwhh9V+BXHYDjwY
2r2Mz/TMdNa7F21llmPl3fXwP78AuTrOYVjv4mNJnuN3qc9RmEuVMu6zZVIT
FQzPvnhuOzXwxL7OKri6FIf/0BwFy881eLGCRdO9kTPZSvScF/Q19+Zpdqz0
L0RIDJdORAj+QEAjydnQlEGcwlA1KrhPx62IbOw/UA2k3Q0gYV21yQYXtm2m
bqwdt84aM5NLJQWVb15KgKW1NaQK24mfR1cdgHW9BKGdw4kd0mwySUIe4wJ1
PNVG9a5pkbfSLHlCnyiTh99s4Zpej2tjQISpnZYiOQ75iGbeTkIJ1JRaRDlw
k8Yfe+1TV/doQenea54bu0SH9JPkCBTF+g/qbQbk+QO5C/ngjf2uSgV8pqka
gYR1LO+eHdl/CGedLTJFdg+/tqJPnHGLp63/HFE0ZHc/NaOVsvaXNlSaTQ2g
CkWKhfiCtNrYq4bgQhmGzNwxoerWCyuW/kNYEF7zyWJxhbf5V6MxUPbPkJcd
zggDTEbkZiC1lB9a9RvsO5XxReVgzOIqT5B++UWLKSrfEwHGHMCdzywbgpcr
3rfpS0Ae2YCB8ly1mEPKj9Z1xeYfXvFzswyjG1dhF0S0pETge8rET813fZAa
euJWuQ7rdJarXooGF2ojXw68ThbRa1WLnwNSNoj4CV+P2PNdxO+PEK73Uk6x
fQVRbfd5c3H+4cr2CCYm2Zw6qhcT+t1ojwjK9IzvvnZhrVrjjdkeqqa8flxG
VPOOt+nKGW0wGS18M69p04oCFsCyExTN0REyf45//uRs6qBe4KoSmWiYTm5p
pUdyVc68tyc86OXZ8oHQkGhPQq78bnddYVPUYp9LDFHhbv9xcuhRJF9foyQy
H44gkCJQ0GlnejC6GcNt3VB8/EZ7xCk9Rgh+tjXBdcrZSVr+poW8lYi3lixT
aiLDzbxHMRlok+Tmdh7z6c1G7LOXzPrXuKPDaipunmThH0qDM08v1tenI7Qm
OW0sUZfMUoAGLX1VwTOnXghgltwgIP33+pi92dSYSQ7cmgLSx0f7Jqq8ICpn
kiToIzQlMQTmN7WQQR48vrikPpl+lm0qtegk8N8Uxls2qiqmRwmvb+W+gdID
veRZ/8LIYfP7P3UqOraq21vnVHNip0F+6fT8VvXNQ2Xx6Dp860E1cbJF2yHz
NOFCYemhNqT3nRuFpZINEwEiNpMPmVBV6MaHjqbEorjY6YegbFIn8Iky5K5O
wpLPkDG7QBBt4IQRspo9vCaNtqgjmZ/FI0/5iVyss5tkaE22pS6IHaJNZWoP
661fZ59aALp3qcKEuK2Ojg1Gpn3f7qGFQlhhWZiWrW7Hc1q/a1PLSrYcRMoo
DKhOe8u+90jeXka9IQme3ScX2Xexy45YL7XBA29IaCL2JV3fdoKjGd0wcB5V
yT88UO0nfkvAhLEAMlgAZAXnAwMe2IP+/plKi5T839JiXVjPYVg76k10o38G
nOMsqh1DGyoMMvgcKJpseFeW99KlnJB+UtNyK0eXT5vDry+/B5wWSD/LvT3g
rbrZqi1g31Zb6aQH/Hgmk/3mq5v/kOy6xxYoeMJv+LL7FmduczWUqWfBSlz1
SOPcJRg6KdPOUOBE5PHezuQA5lxFPkdLgY8FG79LvzNLz9qCM1U4rW13vJv4
zyKRxoHZuD/pXSdpE12hW7ikVCqC7UUpjGLyEtrZlWerLnIIc7LUcmwqbOtq
wVZS89YGwBqLedVvgCzMGYQd1vIUPgpTlHTOUjWB5R/FPXaXj5e1YYHAgCEK
p+zLOARikz8q4Lb9CwXterK9S8jhFRAx0EkoSi2je+M8k7QfqjY2AdYx7Nhp
HQ3vfsPBY9+WpiosdMC7FXks8lPA0KXdhBAp+QQqXQv7SHDBh6zMxoH3017L
IMtw4zGEL0imD/2sSEaG0vzDt+iKBL2oIazebjBQJwJJk54YCcgd5Ww3RMA0
te9r/IoMo4V/UlRuM65YPcvM+V+se8FqMxXbCydzmsMs18dNBElHIVd0h+ch
r3PxClAZyyII3Kg5hYOscG9k04BscWrZzHgZNU3rIEWP2maVmQ1VV0jIpZps
UZvm4h1bBAJ/na/CxGQhyDuSoumk69i1IauW2RmbRljYHwB9q67hhT+FR6st
RZpUP0Soj3DucbUqyhma7zBzg/1yO4jeSSRftiOU0A/OUTsuQASIGFNVw0Pe
pxpDQaodk3Sxvf14BeqsOvz19aOvYbmGHm9KHNCCSldjn3OEC67AgVj4+D2m
MGIKnpeOOm6qqiRnWZ0gCWB++uGberLr/cYdRhzdjYNM+ZKPHproQdVOOl1J
TJ9++8P40YSXYtSDhgyJTtE/9sG1IYsbZueHWsff2aViXs+q8GIXoXpuiEMN
WW8asHZ6/JxJpCtE9RgHbpSBwA6oXfJP9zOYdjiB6HVGfZBYy7wmGGuh0UxC
Wi/2Cuq2N3nFZwQOJbJ67EbNUGp8fdCpsO3g/retO5S4qXLp2hEqdS1rYrea
uI133YHZRjG8juW6JA0HNi1qOpMQZakVoqMN+VuA0dTbbNj4cBhBTXjkJTQm
5SdZBIs9v/BW7Bfa6oILopvl9CL8pkDrC/AykfL1no7oT8w2BsJoNULSkwaM
DNgKZXKQ7pdmWyKUn4+7YGQcoPzoPMoJuNR5al0f55uoddEhwRb4kwUyk9UM
bPh3cULKj0c/qsLfZXYN3Kc06vnDJZ2nFKLd0JjG3UnA7oI0XtiY9e1KXhUS
pbTo7R35yF1E1TaNfBnDvuC9XtCD5Bus9cr4Inh8tN3zWdIXP+6HphlFr2sa
K849O+gaHbkothdsM2lw2kv4ww9u3hhBsLem05uWC94OPza3tH1kgyJGb4JK
TkH/skClLC5TaLCGm0ztGbATeUXUhQQp02dVRMWjDfSEVqfBCLSwipTc/eG6
jkDMetQjCkti/6WPhk9KlTy03940nby1Cl8k4mDMeYwLDRpasVO/fX4dPiNo
rHZw36bQ1SivhRxOkdbGjrZIEav0Ox8CR9woO0VatfluTEIK7r4+IxshEcIW
cUzebk7jlegT1xpGUrA+KHzgHvtvuW5uz2MKR0mVjdjwlOX5qU46hhWypwOQ
MawIfrKgIoD2r/T+ABuOdXXctgCvcOT8YKKH1aE8QVZEqqfVyZiyjc/52OtI
ExBb/FMIi2CjAWm+XfKdX3k4XoDXplfBDayyuAJDrCAPcQ5JBmEzl2JdLms6
5HrgA22skZkB+nfd5kQ9ldDIovJKIIj2eJ+pxSEMGkltbDLqeDy7AZ75mz2m
oN/9MZn/p6KwAgNhxpFs6/Lvn1qCjTzAU+uq7NSWG9b+DfAOGgi5ifqHYSBD
c2HI9ZFGnMJ9TNdgRQR4I8TULm3AfFUj8de7Z2ZRQ5TLTZNs7kPuu/7mbpDs
N3bq2ComS3dMandYFdurFLQS1SEPKA2vOVSoYoxxaJmEbvhZq+WhuJJTCxHb
KImW5z1UHfoomMsBS0anmwmgYQcm4gVu1xb1EhHJvNRdoRJPk65gSnveS1Le
wA9E6fB+OIRC2Lbj+W169IS8Dg42rq7njAbGLi8DDhJRZuQd9tLNQ+ULhFBo
zNoGXC1wCmUWyZEWKxZJ8+jNAhDyaftKXTIE5COm+s7EfiX1CniIzHRFp1Q2
kDZOkdXWGBEWpOAb8ed2H+RinigW3EN/g3VquZR3gxs24FiZsh20aBzKqISL
Ts4WVtuJ5sQ3/R9f4nT0O1nfAD2COalD87/3J6UbMpcQMvv5aGeQwjcurBy9
hSCnoAHzCfOK/74NChp9ENvmQRxY5Dpe8Aa/fkTCnKW/hKss1PHuodWsZ8WS
RMmLr5CNNKzxJvzzRrlB4kNdUNsySJWL8bfDZH/GWms2p8iSZRGr6MC1otQc
vzVu9xjhyblTFQtEyQW2CmkSkm9hNgL371zCkFny/6tQgxsnZ9eCbKR/nSZa
ERk+oUsqyHK1eWoGOfshLh5VK6+ty5lU4AgIWrWCkHfjdD0VAswDvyj1kx0U
l5iss0ljjDmkCR+OQc9MD5TWQ31LhQmrNr3HE89NOoj8p0jMSjIQ58+LHrOt
rtN5EPaLWNIdpQfPeOag/BJpvvuKRK8xdXiEfNZpibGeavDNOiwLCw9Zx9BT
V8HPDRyhkDeBZrKAejkc5HbN1GzwwoCD2kILGpyhNk1QVC3R9i0hLm8wYgHC
4VMQCCf0Hy+mKG8+sICAxnXOvLZSXlAA1M8Lkd4VCk2UutrN+O019OMkQB0h
hytuuXRirvYL/Kq29xwHjBO8lm3VBoB+H6J0NvXgAEPfIKEDsaJvQzCVpbTj
Uum6Z8GJYb0YIKzRmIPQFXbupSNGDJ66L6H0PmC2ajsxmuHY70HdQxxycAMb
dGsdgpXoA3yg7nbRQ4KBimXBlCildZS6zYPZT+mgp9zh2H2qYiuA2pWw5Aom
zx79i6P4FLGqFtRzRDipBE12d4dzRv1lxX5YLAqKso9L6tadZq13VXQkpoh+
1klhi+PMveZHKAirLlxipIm9gR3alfsCJRR9R2jFQ+PxSeOaTx7rCCZpayp+
xsBlq271tJJrfgs2N1B4X+fSw3LTTVjM4KYMM+YZtAeyF2bXBfZorocBEby4
xt/kF/avTnUIucUEK7X5SxNW7buQLf512pgxrNZOgrrTzX2MouvOpIw90/Sk
fcO/0Q3oJMOglLO+vW0cG8A4s3cCgExFdimtGZyy1HEpvVPKit0Vj/dBod1t
V4hE7d9NGfzN2t10K2Qt/bMO9ajbXSIQ6MALvqye/qGJN2de2QZvKSfXGC5t
2nA4JwlEb87NOUDN21Q+wpkMuwi9JYDv8WhBesIAvfeNHJBtBre6QT1LdmHZ
8LoebxL+HEOQ6G3cTlmQVpa0oXZXyDSaoP82ixFVOoNu4diqTgwgWBoD31tE
MK455tvkI2aPFma9ucuxBUncfM+iW6ju+aaIA7soDjEbzSuqxu6osdmnUeAL
/q9M5/EM1H3abRDtjLRbB7y2gKynsmdf2FPMijr711ySmemdLCjlizZLlr3B
h5pJFjTd/ka6BkcUkFvyEEUaqwc6bj3wOEQr3oBaNVsedU6haxlrWTzkbGB1
ewhT7HgvwNlBf5jNdNNKr3+jGkRSFaFTunUMuiDxuzBUJTciAHRZR+2ssDSJ
RU1SSyadr/bWmMPHMFznW2fNggNqj1uREkHxUTx6P3rKx8u47PjObgrHS6a8
X3tsjf/eJGZ0WViwpXSWEdzPIbldX5KTTG5VcIWh761/41zJO0ohAihZh79U
w1RIDLqzjwUNqqhfeKeNBJMxXXgvsT6UrGWb6/o+7VAvu2M1IEwPpQ8Wt1xO
uNT9c3+JcoX1Fu7cdiWt7j5377BTC5SPJDEMarXv3cDFbhYGhqNYmiaRuqho
E6ch8ghwdi6Mk7W7DgEqtn+umRr9osFgHXq0MbmSMbNm4+wUcBpbsf3F+M7j
4UYvFBsht4qKKk7cAIKK0s2JJRYrKemWwbXODqrKinBHzMG2miVcZlKkVOci
gc3tEjv1/WTvmEaqOdLy7Y2AYnVLgofwJQxkyIQDyn+RiKt9B6p7M6+MMbPJ
SBLiJ/TeAjr1bn3sQKfKColeHw0Kuxxu+zPexGdl5dizK/NlIxUPvfnwuRB6
fvBWCucrEjtlj23guXrxyUlBznhvWJCMDvDRQRbUZpyWot5njqWM5ZdY8EPr
zNH40FVSLBIpxFbuZrbqC2u/4xvC8r5CW8VmioginM61JWc6Qo86IPQZTvN5
wfXhIqPBCgXrieFZ+yqt4oEm7PL2lWDAIW0Lg0q4trM0Cj0AefwnwSiljj7m
klLz1cG24b2zgK5tNssafIlJS87MHX33fw/L8K6Gc3ScfJfdd5ckUshE9f/j
T5EP4JwS7fXglti/3p9cLXmjg/NXflYrNRQ/W00RM1ISlElS6hRWMgNkuImH
ef1UI0MU4xiqjWtIAR7f+4SBd8zIdhM2cG405qxNccW/sYp0lgcGeVVQ5IsE
G0cBh0zW6wOnI0sTSG1/LiaiElfbngYEL7XVr8hNwy7yqlPkVDdR9A0BTfHt
+MwYNnEBFYmL+QM2dUni5B8VIcMJaL5j4pPmSme1VhY1bKjdwxpuSEy201a7
UGzEeHPJHP1SXYcHdddn9ditpqLmWFWOwme51wjhJwV61kyqyXlIWeR3QuS5
QfgUk9lQvBjPI3mkbbmdJvTrFiWZXCmmKPFA9wt5wSNYT1QShhXRcm2rc6fp
HC9nA/dXpumadNcYqD3FqvvRNa2yiswaAKTWf7koebYIGSvlU/tRltjmxbb4
R2dfYfNKpbtLli0ss/ra7dgf+HW2z1KSWzxFzGtWr9AqcucsBRdHVgWVKdUh
rVEw33iL22cRszfTfUWx1R5aZW/g9ta1GKmezCc7p25GGigLa9xnbYab3Q0V
ZdicJBHBnESfwiUVi/nfvTGVt9JUuZCfbk7S2O6Mu7zYPulRnh15WVeSjyGh
hQUIwpvBXwOOuPjakJSr4D9cOaOqBipHVLA7wwC5S/B4wzf98HKInUTf0C9I
6SbD2hcIJ84WpBjjYCqF/ki369kqw90iZp7xyIfxgazOB7YwlAow/VSqejpS
WqTCk+yE3xDAbIntxXSlBPLzq95LpSoQow9EL/O5Y6ylA+6uNZpZsLAWNAO2
uA36DTW782BCZc3etKGCs8GzFeuFSI4TrofTcRYVg9C5451I3OkS3zWMuYVO
/Tw1ATbM/m0LT3VQ/4wDVFeHWzTFUEMrtUBSq3r9agaSgydNEF7HNce45rHB
UfwjIfvsom8gVU9X3zTTQ4cjeyPdsJpakfH8PDVy+txYfXtWDTeqT9yseYSo
dPj5NaXiWrjMQP4ZC2Xo/jhk2KvhyOTHJJCJHB6Wyy7SJP4Wgu4SFMVJ57n6
ILi49+7Cz9EG5ywyI2Woq96hPXfZHBOZWCrqA6+p6omwPCnXoxA3FC5PDjdf
moi0RnTXsjgFuyjGzMFbkZXV8AZDYnFdbE8l1pI2UabJPirB5P189W16+BMU
AUzpvcuCbrWgi/vOvyBODW82pYbsBaDpR8k1nAGteCAZhUVNRkrMJmNnlpY5
qTHRdgUH/3zEeD8UEprotn5kQcnjNMijW+FFTeYpgfnJUuMkBvnOdsLlMsqZ
8gHVuHb9HpZ4Ts71xjil3ZsC/fWAnSNDn3UdAIZcLNQeNE00wBWffujYmTO+
s0basxwcoDc+x1z4Phz0naK+XctX/Jz/eRf2rwAiP7i78PUII8MRJ19/SUs/
yK7QEHR3EA9ND3TqLZKo0ihJBL3giNGHpOi1E/MO53pK5R5K5T+5+yF6C15E
B/hv1TJuwnZs5XxdAFPC7gxhPHm9uH+P6OppmfqSEpg4De+cHx2afcFaw2XQ
BDfj8NPJ4/lm9832WObqZBnF7ft9TZJIldj7THxc2mDpy29UPxsFkrnsQBaK
/soDKNykcrkVQf/gbcliHPtrUjC6DNT9SRD3DJpmD5A1ZMpusVv0rc4RIbxB
Qr/wYLCKD7blyn6nTVQp70mVnMSSavTysVPSP9LN+af85xVglxDtwOJeRMlZ
IqQzsyHyP50OcDj073cXml/cptyuk+GyNkTujj2k9Hywx355b3TxJanB71cA
UdofkxCUi4rxovRcWEgUfeGCRlAGbwzw09yKTLRAcw3y8QwRuck6c7dPcFNg
tzbjCk5AivTwefmypKyBb2B2yY7JAcqXAYz88aTz7QziW8EQu8NHkg7xQaSQ
468ffcr6Tv6l9X/LvfreUxb0allevEzprduKBUCnxbNHy1yrodwh2NaJSww=

`pragma protect end_protected
