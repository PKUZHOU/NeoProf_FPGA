// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
IEMaqOKEy3aCPd3NCV8UBNoOY4AZAwtBw7t+IElLV7JeDfSo04vnlbCBsfnf
/dLzlXnCPuR2UeW+CNscN6zB+eKk2/HqWW/bPCCKNXORAC4ZY4iZmoqe79WF
QvutyklxfvFiC229oNrCscF1sGZ4/6gHeWXORUgEm98jB542SxrGwFcgVhcL
IipooSY7apjsr65Xrd7GfsGqCPSB22c0eh0LbkvzfreJgGUVYY1jJ5/APp/+
HHDOq+akzbrc6JydMPaK807wm+9okLaUdEJIlJXlZcKCw4Ih+kLSef9pNGn/
hu+KsP/A69Jpi4E5sHKcVbiVMtXUVxZkUzXrippJaQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
TbfHv90QWyjSt0In7y+gYspC8CnGXWfE+GT0FCc/Ii3Q10TroO5mOwOWFWc+
ygp1915heqJ2M5SZgXRv53aAjCsstjaeyYgkEo4wZgBYWOIfmNunGoQfAuwR
xn+/VghrCKTFEJ172pne/7pgj1hWe6EoHwFFYBzXtBWT+w1tV4sxSh36C43U
yvZ0Gi2O05kaMGE0BJqB0s8zUsUCkQnbMWqfqmpabfUlmkLdtffQd3Nq2Br0
fdz/A/hGpJgfDsE3pd4hY1oL4wAOqwekM5vfQcUU4a0Meu22dvtqyInzosYZ
nwI2ECKgMJHO/bduCGLvJLbeWUjhJYtpufKXfw/4QA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
FiGwg64zm4Ge+H2vNUjb/ld6Zhk+G6Lk7GXFcuBidevIM20GJsXE/1NEceY/
sNf7mrIiHDMkT4LOt22kf7zKcIU8bP3sscLi2oNyH/PGR+P/GffzvokqRnaY
IMizgpirKe+NYZfrfQxM44cdk/XCW3H867QNzwpe1SSOmf5t2Q5hH1eMGxCq
dZADHWKwcr4PQKqGKZirJVRZfpSLuuDA4yzB7p3Z3Co9jPIU+cXyCmL9XYVz
/FLyDYDqBkG+XvOt/qwfD/22v4X17cNNIF5jsG+kBY4lVYHl2d6RfPnuK/GA
eLMMCQ0ZkiN/ypSoonheXksTVb6fOnwwmYGK/wyqXQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
NAIj6mR2ZWA7ZW+jWNS5BNbQlwBYDlRpIVd/Xh0ytyUuJVcqh3JEspWEmB3u
ltAbAANO2DtLoDD6SVius93oT97QMT5hyBCVNYF+orN4HSl5l3HxAE8ZLsUY
HueeQsGiGCDYELM0xOEB04WqCl6oWjpMcd3Zst+qHHDSMBGOx4w=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
wj8kCYMTLxs9kYfKzA9ZT7nsdqn+n+1qnlpkPZ+28cBmXrDbl8nP8GGMOZEu
gw8JJxOmxTjds79sMxfV4kY3p/Bzo7s99G0pKJS4DfRn6Eropjn9splw1qLe
ANBkkO8jt7mhvKoYfdHCwUVAvy1PcmyuMq5DYly1MuMcB5AxbacRLSNOhoBi
AIbduK/oGUmh10enOFdCvcPw6+QyRuPZAOK7lOHiKc8+nI+Q8E6gxou0a1Dw
6Y1TZNpjwE2S3AUyo3tcc1IQoQbqlPqjEJpEww6TsVydjMQEkfhmJWos9Sld
90zvg6ypp+b37X6nAc1ylB/ax9uupro8iqrTcnbFGdi8zloLilGo8nNzWiiw
XdyB4fBRRiZcFaRnEs56OX7xor4AOVKzUX7JMlAi56o6lHbBK4V6iPeXXvDS
JhnR2C4IMlAAsc9IQBPWWOOiMU7i6cKMUEEYneg47tFZv+SYcy9yhp8oLFMJ
MsilRzT9xYNLqLc4LIsWX+NNX897fYwQ


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
DvKeN3XqymMCcZR+jPERTdvREcrek0ECqVww5PPIGtktR2mSj+Mf0O0iSalS
aezW1voGGTnY62rlXAVJ+D78qU0iAY4AbJNL9uuI95jhJZOAAj1ArZhFerNv
PcoE6ZUJFRgPR1wHdKS9UAoRcEr5PZnKWECwvNALk3blbR38rnY=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
fhcNVqBR+yungiMJrTx4A1as6nmT1Wzl0bblyekqGG1byYN4hFrJWAir5LN+
mYJrXtXh60dfe/H02rkLNauZ+5utBA/1YSE7UsmHThFMUqKf+jw+4Li083Yd
Jf5qq1iBhyUwRanXt/eQZ/oSraa6PzbU39IBotjQbz+vtoeJLDQ=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 536976)
`pragma protect data_block
P2gdEURvqoc4adg/O5kaHhipgjOZkzaVWiTQRLUHDmFkQiijV5I2QfO+mkhf
hTGN9/LLUXcCS26hni2jigs7zzBezK9zYs1V9qxSgIlogVuBUKmRAJJR94FJ
a0MsAExle58mTsczWaWfWmqcXkDV+dcyhKDmGLdWR83RzBLGCyGm/FtjJigZ
0phJRr+p7oZ8KNzr45A1USQasUrFmxL81m2f3B+IGOasV4hjrnDvA5xDQe5N
M/iJQ2VI3p77B4bnoWxEvOaTQChcGuDp5qp+3aOxYcdZFFFppZXyoN5EtGNw
pZg/cL7QCqkKNPmzZF8Q5Lktz2FGm+BF/ZI0NbkHEos/2JtwetXg4dpRtdBj
y3AYlC7EJtFtki0iVh3hG5u41gHm8tkgVbW8A2Xl/7b0qbs5uKIp3V0ryAo9
7lokgrTusEQco2w8G0iol9JtBsDnDuvB9rdMEElTV0xKUpBLIChUG45eaJL0
ULzoPkfbpGjl2LXm3451X+ipeWMjX/rQQ7DpHCP+QO7be/C6gyjvd90hpX/f
ZvVHFWmqsSGnAfN1gXOVp7SbvtHsM3PGDqvZZvCXEfB6k+tvR4AyzWhiFZrf
nL3o8D/441rEoWWNmcg+/ZJ7N8tKWFmZe1OCdfYTODmkMJcZKfVFlkq5eVML
YX25pxz9TyBFPB7DLAwg/NOx3Lfrdn79TrU8D+lqRascfq2/j5sEMP303HK3
wdVemgFNGk3ha9Fg8p6Tj3OPf43VXJ+lBtqInqlzUBPJ/IjplKyZro3SBnca
3AfRJBxWZ/XUpZ94zLm5/jJN66siWWBJZxNsHnwmPyEan+BV0QtD7bpr5XtR
6MtbJVZvPpIQLTGa55Zlon4X5XjoojIcCYhWqs+C76odRvWl8Upm0mmUCYwj
/l3CRCThS6eW4xlAxobdGqYtFAMDYbq9jDMtM7sRfc2tUPAsA582WsS/icvm
AHFMYBPrO3F63HtBBnYheiynocwmZGuEkOLnTqw08+dG10IJsA5aDKBd911l
Ta/L0NdfQmDnLIHWT64gr0kC56lAWGdl2lYWxSGQoOsGDYF7D2tFIGSu+9De
xzMriYm2xJB2M/GRAJIXQbAgzDx/Su0idbOHXviAeQ+M4Z5Zvxu6pdW6u8Eo
B7W7JvnL/NQLQxTSmsuTJtgiYhWjEsK9IVWDb3GAy9wBfpt8BrcnM8NvLXM/
LJsC569MLmm6de3rfVr+LEGe7q1ec8NPYj3M6kSKj5u7vxePzevYkr0rfIWL
XkmREsxtG6T0k/0wMDiNEDE/xNT56gWPRL9JfovSKrZBY5+JbmU8tuDohBpN
gX/e7pu6jE4pfFwCVeaocl3zjRlxbwacoPzA1gRbCzYyQAByDBhksPcxDVXz
X+x16MttGAQYrAfSQzAirSdI4fXxZOimdG6jYZGKcNcFF7JzOYY4Xr2VZdKM
yDwdYu7W7OqgRH07Ln4LA4F7qD4YTcUxOsFMb3Qvkap1ATn0kMEn4lX1Qs9S
NFNmxq/Tbk62SmbA+MWRp4Gy7Z5fAnT9VNuFARXex0vmbWrxRJjOFB5AGgmi
ZUrVgxF3KQ42s1fHSBw8Qm10V3FR0MtBxjXaNQuJ9o/xPp+tE0rpli05QylR
6myLGcYgTcPaAybPJF7EQ/Qt6bKjt3mIoDUTiF5PacVH1XGQZoj5mkByA1zV
7H9lcU+VVFxQMEUmQ+23me4bILOZ2RAiU6JYk7DcOuGkuxQuChu9nTFi5Ac0
5DxSN65g3ahMSEvGXyGxmQF2unDp8VYP5besg7zRf/lBj+IoBdwgnGrj6FU/
q9fBOVpm+ux5SMRnZ4Rc4lheiAXZMK7gkMLCcOFshwW+55KlaYqIBbnH0WCl
IGXSvZFSwBd/x9dKcDYkBoeLMY4cMpcXu7XYP6Ff8RzkzcpiBBQ7GR6CfrFz
3wJq2ehyixuPivqrOHg9GQnlvHK2UHU28XQP3CgWBy2dxZMn6ef1OcRB1Kds
7waG3uJYsI2G4OUWq1vSePhY16nhgGqhJPB99xk/j3efyk/55fMYwKt0THXp
aY5duJhoreQThdeBoXWggEOEfXCKETkxvZ0yk0Sx5XjmhCO9kbq/kUx8YgQX
n/MflCu93Yn7INCqPBo/MHAxfYz0GGqPkviYx1eAKoexjAKvI1apbPvLJSsS
eQpGkToAq/IKQnLG1YuSUemWIFiB0GiVxKShbrrMhyAAmYioycy8MLZaktWK
EIfKud6W06bme1R1FeTwnuTfQiu7FRk2i1lBd4rNqH3nFJDxNcx6oVAYJXn4
laaYHMLYSEjOUaIu556/4c2AdAVncqS4ab8uZ0jItpa4NQ+4ZMueu4Fwcn00
/YGTIN9qsLG1ErlKsyL083HVIHUuIstIo/5WgVL2Kdk650GmtSf3WZDL+rEH
qoxpoRGdowula07GgIRbavs1bPCN9PFNeKWKKVrzei9RiXyua+vmtzlVYZvU
u8Tr3UlLJc9rq3yk9al2Gwv/QJrY5INbvcyX5DdDP1aobHyGL9EImHIrqI/S
anxEc3dz9v7k5mbA0ZvfqPqWsWSFB/Qi7pR/wfKv6jmdM4VsJXNQ+bgQopXl
PDw3DeWPwF/MaISxZmFGR64k7+Qu50VFaGcWNUHERyL8KpzfTFC/FQs1URkV
dv2r3rQkU662jTYPvfghhTrybfIaICwyk2cukCBu7/Lahilo3ctq6hr+xHRR
+vUjoGk4rolA1wNRdM3rzu/lKlQI7B9YNQWOMmsKSTW/2+kdMU6nBK3RY/t+
mQzoVN4cIvIRYEm/4/0AHLR4c5jaXePMktmM0XZ9EpSBTPBt3FCjE2BVkQmD
ycIlmqBZGYKj+ZnmfDACOh6mCVVPh5Lw24yqCEHdVMepsA1jbUvTNR+plZqx
4ANshmpPfiUHf9HNuDnrrUEoVNMbTJAeBynScRWttokRZSeqGXSLn777dDgw
mdPqNTDVzjPnE3iFR7giPVKYERNpFvfkdKyho71uq19cJhU0b3eGumSy0J92
PDgfW/EJYXL6ecb8L4Kamr7NRb3i6NLyVtH9wvb5f7fXBP2WlDPqW3NEy53a
lQfDryywydHxrONl9z00lSestxfNizvl2YKrs/QYPg5kx2Ygj+kE72EQVox6
S44epm/eJZphr8blyHdUdyfpeDy7EkkuUjXofaTTrpZo8Nyn87KBcE6HoZ6k
wOkL6UyoPfmE5Y9dxwmj8dYU42+2/ciPH+AfIo0rIc2ZR0pKMJZN3xLXr7BT
hWscFfFXSAvZy0oy9eb7k39Jdcn+aUOIWIfhuXWpfJQJwyMVBgwAfxmSH6sB
PoP+o8Wc0LADAsDVtCHXIRiahalTPAL23eZfGWf8L9B4GwrNqn1blSCoj/v0
KPj79Qp5JvzAm5u9JLi5JXoHbninTNXL9PaUoW5+tOdWo2kAJU7VaMnOxPH5
rQWOCr4uugMAO4TxcuzzKIQZSwCUWXOXhmyNaWiBQPSdb8JmLe8Y5J0ZvQ5h
G05v/6D4xaW6mMMthS3UPFJxW5X5UOaqDDozAq8kpZjDYWNpaSWKqVSIOWZL
XYt/93DpF+MV3uJ0d7JedGdbMaq0giW2QD6nk2bIMnMhtUwZfA1du6zqmetN
AvL5J0Lz0VIAa0nEMF64PFrxgeHkg941dnbKjdXGbwZcaKQ7/CGQZm66G9EN
/5lEThS8xz9pgDKBWAMtdy3msDVkZFXxk2xGztLbCdjnXFSgmNdoYRx6XNl3
EYhlJp1ac8FzySQy/EfBOAAAoNeWljedo20TuSwz50VRM89SC1u91RYRE2u6
2rpFpbzKGcoGQM/e4pMySkXKwvausQoKzVRltZJYm3KRotGsJS4hxu2s/8h2
QyfTwPUOkWRcp8CJtcia1jVo/W29h5nEG2cWAN2ROKxR8ijnrXd3aKJxlRYn
HNucxJpCnIRoQYA+g55lIqp/7KYDskyk5JEDfuu/m9koacmbvzKVDvm38Y+h
30xuOWPvLJexnwDONCuXYzSvWIgrUTrfrD/eSFLpGziLrhiE/pA2TMlSWhPM
bBNZIh+2D5ar9rO53for6PH70GudKp6xaXxkkNIWVhpQXMvM5hgJ/jMHLnol
XfX1DC2zuPlv8kIvmhOisTanWO+bJvEUH3b/wWN8dtA132bwT7/21kbQk0oi
6TlQPlvKjH68H/ZAmG6Zkzu5ushShtmApCFrhLCtzW7Lu7Ygn59V6moKH/jA
BfUhbpFLtUX1t94jISJyCSHOdlJeHLF4AXg+TEDjLXu79c/h//eH4k811ziK
5+Enh0MAvNH0Eohax475etMByD4PFgiMJ/dLwaTz9QTh5LIk8veg0ZcTaIaa
H6+GYcK/A0ltGAmc+gYgRFfCDNy0etW1zGfWihr5b3NjUkL+31T2qylnm8cO
sEvLAleGSxf/WTj78CSAb49m4soVu0SYVx7F4pkQCz1Cd4yvvAitiDWDNpdA
KjFzp24sOHJgxGKlr6LvfuChlzW/oKx1veZcbv9SblUCfvCZMXpQTKEdDGx3
utsC2mb9Yk5qX8P46UT/mk6N2sKD9KJcgz1BhbnZlEyTsYkvrbmjKEfqzFE6
ukAbEKMozO8kYPlqhHQt2eyNpw1ViZX8g1ZkR3Fz4PoRQ91RKCNmBcPArx5a
+0sGykwzIciAId1hmS6sEkOlQeOJkXRQjetFVkGgLVReHSenKIY/+h48t57R
dee8d+tRkf8FEopIteX6WYjc9KifvmH8YqluOcJu3gx+wMXXv50+JK8Posur
r9vDwqraMeTBuOONNhcCTMUGeXHSWsoO0jIOcsEebrW9RiW4kFWUPZzwhjKe
fGSfcNed/GCz4Si/bjwy2KNkw4OOs4B4dzEibEQSi+i2MH209KtHVxsNRCFO
KT3VEYGNzcL0OEjIbpH3GGJT+zjd7O9EhgJdMDXKrS64ur0bxpjtsOQgePJ9
6XV7b3a68c5aFOEkszunVn5oWvX/LYjLdhK3YagJMktx4c3gd/WPBGhhMNTk
mVDTNg6AGKirWFEmXr0B47YTESW9ndz841zTsHk8cjiQW5zs19emDdrS7VLu
/q05za0B3dCN98IKVZuK+PQssLfRwdzMYOEC+XSr4bWqFfaCEmZxxf4RUTea
y19n4iSGkRWDRnT19pfMFgFkEhODYsbi7JZq6qFY/huaYoYMUIDaxy+6q/NH
VEISN7wL7TYSYY7n/32ml8V7WH3/mcuRdvPlG+ygGfhFM9p4REalTLJ0MPod
ebG7ydDXw1IEbyVNc8cpK3aCyvf84yeD1pM4wTgYlAucHRR3+cwRHAlMptaW
O76wA7xHjcliMzibxErkP1xhXMTf4lf7JtUc3ZtK9eQOdljF6Xvu3a/RNx+l
9kwinVBnucaqbVedsN7uzasdusVgH6FPWWr4YK1RNmTD5+dPLRimZjAmAYCi
NcxjAcJJep1UjRlIOmjSQ8dcnUJ6g4xK1klww1WtrrBEJ5P3q/6eF3ANfKhx
BhShZV2aeCItcn+7oqQmhSVkcRkYRzzjo7f+AsgZk9nm9gkftLv8vsaMx5M5
0X+FsNNLKKlUuB7NlN/YLmVxu05EfFUeu1IFF+fP7+drcCroQWWACd4G+4Kp
1BsqELpk7l0oBqhYxmklI2wOhaHdr2C/jJ1NS+hNHHcnbeOIspbY8sww+VxV
gyA+um5JZ892dPcZAy6ikQmAZ9cJwWNP/6vmFK2ZxG1p+43XGNafdoOgJhKW
6JqOBpVer9aF9/JIspwSlm1ZHdDjCuQ5984/NBNzKor9rNrmFP1WC+wYeRPk
Nr1Zv0eiDYolCPdrHb13SKyJqlL/6gjRokExwu0UEdl44HLEKzoAAa8adMeW
DYAqi0eNlQH+SiGXMVMhfIy+nK7aRCia9Ishoo05bqIsq73qFBKhygOc/0dQ
lPP95A2xJgJpx/fD/IossZmZhByUQDvhsXCGbZOImAD+1k75Xcd2PN/32xjE
R7oORvLIGkOK5+7gd7bAiwO9aLe/O56dUb+6k4IEnyIsNnQ1yH087Zqhz8sz
LcoGHVyEKFQy+tg6sfqbGB1dtPpVIsvdUpFL7/SR5wwsADzi+P6zCLDviSEF
4wToRz3JakYXPFU6ZnvT7XPJg9rbY60xKm57HAkUYEjDdAN657EgAfid8pTI
E00cmg1xcesDWVYmHnypAGWC8ZlmPBnBKseokw0wCWos0OJ05dQot0CsH+o0
GCSB7on1douj8Qh/t+4ZA8UQKoVeRFvHTrjtXJPFFdEl7WnH6CTjv36IAZTg
9uO7FJJz86HSRvKr5iPUJBT39pPNo0ufuNc440bbREJEtMxjGYBy0O9/hPh0
NnyMe2zMp8PNDK7BvIwzaajGcMpSv5NWWhwBgeFRwS5T2ns6nf/JgH4h6YMX
sxOKcGi/ksoyvOBiRvidGU+uB/xFRpKM8rOeidVaRNDtq7bQ3QxnuK+Kk4dK
Swr54hAFX6PrPyo4nPi1+li+TfkEAEzUevbbdk9o3Z7DCDv6jscIOWHsj3KJ
nj5Lzvxdj5D/J+sXs0khOesO6b71chDLfHGC7TwHpLbVmJH0xEuRc3bIMwaM
xMQKKPdubxBEjUoqTRUFdFHPsQnRPzgU/fDzDGkQV/CTghwdkB4Wqed281ne
exz5AhWb854YaADKMW1De3cxSxCnRkQsvseR58rTYO74CQlE1e/etV21kaf/
JY381WpUUBfvJhN6lOUKAZQtgcgqH65yXSE/Vs5Tq9VAcH2UnZOSU7dQ3OTx
CqjgI1L/Tgv0c5O5HgmOhR9Ae2OiceLKqud4Ntqh+gJsuyb7BWb/fKOK2q+E
cnSP5Nd1Ck5ZzDGVhJrBQrimnAgspVHqAZSq8md/rQc96ozOl8KObu13QRbv
HXjIWe5gAXbDf6cyh5E0pBH8XWTEdemq0jt7LUhBWvL9zwOmfFwi+xG8syEl
u8nW0bttiZmrVwEs9Fuw+eaMihHLOd09wEtnSZkR/lwGJBQQUIm5V0/b0XbH
OwhCDpcazl/6WQLejJL5c2s9tJJ/oGqwD42YlvM/xynBT+OlgYAKXZtWXma2
SI5E5DP3llcS/oMVWFhSEQf3I93TVb8AEYL6HU/fVZFqdEm1gw+zdPrZ9pFk
CPB01/x2t1LeHQ3mlDOfRaZamnEnFNx87sijxUQdfdHmKKdF2O/wH7OAD/v7
QHjODdy3sC8545siCEE6jMHIUBmyh9GEKIUWipR21buCmETWTEUFdiiDdSqj
0kURUCveNreQ8v7j5FDFf1eHrGRyJwT0ufO+LXWl3R2kZvptEemHq28A73lY
mgmueewX5fCieAE9/S5l9LDEp0Hysh0vi5Vvw+VD0k4bQRcY8JCHdXH6MYyI
EymOmL7loSQzie9sPN/bcN8SOvMJYbdK70zQMQIVYsNZE/4tBKjZsfMFTExw
U6uwV4KjNpNHUTjzl+NmJfIbS5s0ShugUHUHp5Oa2d0Aw++jkF6+yzaGHqmO
Ko3kDY41OO1epkc4+O3dRpbqbx2o+ZWKsyR5GFHmt5j1N6MA/Xs87ZVNKjTG
wLzoq1RGB44KrODbyqgw4m0C5nEO8e8zqIe6wbKinLq/6gqbcF+MjGuX8d3Z
ILPkbOxvL895+dUqScFSebpb6f6QQ9C51ez1hRK5S4xZJ0F+aA5lbcFk83F2
rc4611EPK2Wl9/JWlE2vNSIsANIg1pSebN8t2bJa/SCiYX4diaaYS8pSZyGe
RHIxClNWLJNndvXlqHE45N+/qrgv04F69ra3aLegaeFME3pJSau4WOWgScnZ
r/XUpW7SSZX7jjx2py/RQZ9vZoo9Rl/y5Pa0r09+AtH99ohqCu/qv0tyXlWS
0HbIjKrA1gnU1ZjDOxc2k+ujiOCi/U8vkMh5iMy0Fx9Be2I7P7knlEE8aQim
aP3UemTaZOEEWqifblN+f+bmyRbsvEauuOyF1aQI3Xamk4Z09As5DDYWQF44
jT6ZmH6wAimhxRHGfSYFDPaDy3iMoHvs9wIt0E/SiRQVDB6wqhNytQzDEeqw
IG2nMCAn/OPO3W46zW465DoBCSAhBDHllMBegSj4wDMzLkBZ8T50Vo2KCUZz
ifg34knro4pyMaiXgVl911mp2wENwUoOVMLr+2wc8S0NVKzsPn1t1tGN9vWP
ZRYLehh+KSoUXEtP2HV1h3ugKZ/NqUE13jJvGocz7nmyveYI3yGdN25jrZE3
OtgyD+NSkMONxzsm4ZXF136EiwDbtyAIFdVFCd5agkyEGdhn+X1ptIFgEhbv
q1qVD9mXqoI3eGys32slwekS4Tqaqeo1smvxjv0eHlIldrDXFI8zNIchX7Z1
XImid94OQ83zdtZbe6ohlnAJhOgrhgj8WoK6dlpQyFPn7SJ4mkDfJcC86e0n
OjvhoZgcmPDMr1xGLNyfbupwCbaCsgzkuE/F9pbMJqIBu/c/Hr/549uV+P8r
2M/n9vlJbyMsw1Wt3yeNpcJYGuZeLA6UUgo/zAdC3sf/XQjHaZhf39ag2z9E
+NDYybAgdmVXqZx9A4Osvy37XA8lKamckP/saaKX7Pxd661RQmnKz36b1ugf
3FaLmV0Wz3ARDhsd8EdYA84oq8nNZwxdQQYk7ieP4/ORavJ9YznJy0tuVrd6
+Gyo+v7sCCwwlXMcr3YeEavqFkhe1c0XVwdB+2EATGhuxbKl43neiGsH46rj
1/ZG1/XOpVctmR3tvefwoF2h/9p2XSdQT4b/SMMIoj2qVPXVqvexfJ0/xuoC
x0x078IUJ4TFxmahXJr3L4Pw+NbGx6u+B8hhdV+znRADDCpQ8dPPghQtV0R/
hEVRzx4kDYGylo1l9I7uSDaICRs6kxd24a94i32lTWqVs3bxFNlODSxKTd+F
JY5GGoiR+Lv7qgwWfLd//G7MuJLFTNFEDo88N5oi3EyvXUaXe0IBtkBTOyBv
/8ZMwpJ0rvKM9r0OwhcuIP3LnsXJuIFdhtvws68vm4RkcG2syo0/nmaHBSol
nsULBcBJjB08zGEeAVktAgtJDo/Qu3FcsPb0wl5R23VVcDAxQPZo+muD0ESX
NehKUENuOETy/dHSw3ZcIbIMyo4LITXtOcbrmQ/jNdGKF3rboUiC98jf4Yr9
IZ8oaOuqeWftRkL956vfa+lUMxhuWNyzPWkeAS7KxZppTeeZbVZFRZRtIXGE
Y6Dj20RLs7/DMtu6VZmxO3rTmjRjpFhc44cxSKKgBQ613+R66snmYxlBNVjh
HnE0dowj94sjbcZG3DWI7RQ0eq4I0n7tLiyK0A7LZ0gwS2RAtMv8/0+cVi+/
tIaoBTiJRyKc45OMLW7wGt3W+7GzTCVYmGkPOGq4OL1vtukDYv2LBi7O53aO
sjnSbCwzBA8ODaJlos8GpLVnK1xF9MxRmvqNrlypClALDsP1Uz2kEayaufDM
hXfK4QKZYDFpQMBEWGGqyqrejmtOvFjuyOwc9VlK/ydnt+i0mRJY34qpVQWU
pk8iXnJ13FBxfcLnEce6sC9JBEU793RfTvzUA9CNTVodH6QRafYXjp8Cxx2E
r8eN2y88NWn+hJjPQLoNpYWJksew2/QqaU65cx2tf34aRg6kiPZ7/Tco5qSK
M2gfENMeKr/+WgYptfoYXQstXPeUTCn9LVxWHMhqQXrgdOylOtJG4NOqP1uf
fnhLVi+r113HStxHeAju/zPPED7lgCZwFnzilij+nqNb/CuRKR/4nhHIGhHy
FqFE3MRpwW5KctIb5pajlKbIG52zwK8fMVG1LJmsyWfo9AXWdG0BzsU16a04
HuZEjugh4VsZoRTvtEYbdW5gw3gEFIWO8XD3PvALS17GqLnHVybKxwrvgYE7
4mzqx0sVjBYfmgr5q812ltJrEtka643bQBjTGgVlgUhEgpgbfFmkWXD/KR1P
7NvcgzhQ6hqW1nWi0AwkttZbX7RBdiAKp0TXd9E7QAIW0wT6tumaJ4IYh0Xs
6Q2OwNaCMVnnWf6OwRXaJkKHnUeYvRqSiF0RWiFETcKrMc4JkNmQV2DnZCbR
Xm1HOHIbrRD1hb7VZyXFivpDjjVFVOHZJY3YynbTruwtONrV5hrqpp5/j7Eq
T3KBHZruUdkKTJflnwpelcOmfQeKP8nVmHpEw2w5GMzup6JCtQwFwcQvtifR
J+l2brsI/MGj2SwL46LiXc09NeI7LRPv5jyBhP4EnpW1fdf22CFSYzkzSoyo
DDjCS0imfy4o2v8rjQ53BtRp1JZ/BAeYjkdM/vWEQR0VF1ipxhC3bzdIzFE5
wE8V++/6kGP49X9fXcXcBjoH/4ebjvw8f1Qw9Hlj2S4ZPriS/ATckkWlJiFH
8TwiVBkjNGPKWvTuo1G9tOO/hpQ6HhzgLOqrooVwCapqBhlyEbZuQAugm4/i
kUitsxipFjP7itoycvEfgpGbnDBPmQHers+2O4Zopf5n6b8S12kviuXLbIv/
t8oclF9Fu6zmr5kuLPxFFQueQhwDiR7WUP+lyKYnSpxt+RjbbLMRCSZWlSTI
o50Pvb76WFPAvqlDY5cZGO2Gxj74wW5hY+O7Uio+cdpVzXLuChUjoRKScR7h
BeXv2dKGRiSaHeckZaJHjGcUF2UfxskDaCfeBlieT9J4jhY7mJ9IkoqjWGpe
TZAGxaxCunHX7UK18a5juXGNq27yXl614fIn11jE0+Js7U+EHpw1gfLi4FYl
qLR7mJcc/KAylmJ1i38RJ5NWcjHIEuNXg+oXMJIznu19lgSDJp7A+DaJll1F
FdQg42sRi3li5fnbz09gdqTk617TX9844fPG0F2wfkHLamwj8IsdbAToK7Ph
5jonk/jTyJwzFOo5OY/jZWvXcRtlQ8bB+3vb0VZQaV1/7L8LRCWs8iQMOWfq
aKSQ0Hn0yDxE8KqF2vHRB+aj/dzrF2qWVrJUcszXftkra374KSYXKYypLn17
wt81jnEtYGiZnuCFlZxkqvDIHUSLYHDhsybX1KgnKbYIr509nfia/hwPxZsE
B0xtTm8UVNF0HKnFWOxBW88bVDupEyjcWiVbvJo6JKmAlzny9iSWt2IpP9tl
ORRm976oGeJF6w/jUYLXhyEijXYDTPfuWpx/GLKLzrEw4Ss4PoYIqmAUY198
ubgCURhKlcHpbiNfIvTbDV3uVKIsxESQzpfJngptV9ujDedrRFxzvzXCznyO
VdSxsNl5PhaF+CXEVU2QS47JESTAXCgWT26KqHEDdug49wPq2bEaTSFSZ5Yz
s1jrDERvdvbP426+RI5CGPUM/Mh4CY/ZyXjLQ9XYAaQyGeaOFYc1XfPE3Cx2
5jFsiNQyfepJj3LpYXMRbqsYgLlmGcDU24KJTpppuFaBf1AhykBq9IkwtkHh
Ucii+kcDLacwB1AbLazT0MqW5yom01xhbnA1IbvJw4VD6/Y5gYMIijb8NQDz
rZYuuqt2vq70knsm7YcxibJwF6OCq1mUITqBKag5Y2vfprJZIOKn8DyTUN8f
pbMczevWrODVtK68T5WxZKJvC9RauDGKXwCymEaJbMj97B4IlSYy5/j8I9JG
m0m3464P09v/KWI6WJw5QisAJxp5B4awuPDzAa/HFvcdWgNp8/2IZfujq4Z6
ygls+JCsxIZjND3uKe1ugiGmiPved2kVmQhjb5xTYDFKWc8XedfZORpgxODv
JSl7DDZJXFaHjRPi7WoUfBHA+9c44I48Q8zzkrs4Hrj8CI+t9aEs0Om7ELLq
84yUKpgXPvEKoxp/4VJr2qyxVS/uf6V/rLFVGPHZym2TZ2ZTFRH/uGB9fkTy
rb857d8IKAN7wciNkL7KD834A1O3QMw0pOJ1Ncze4Bk37Ollpsyzvdrm9bhq
1z7nS5krtde9IEwek5j8abqDUj82avHDrfPET2bCX3MSkYi1n9mQnr7t3Yyk
c8LHck+fmXjYd8ATpblNRI89pWNnubZYcLz8NTRmUXMkT6M5tpVAKKEPVE1d
dOhk3h2uTuWLqxDGMhxUcG9tN710LZPo6aXJzm7cK0yzB3hc+8cV+KiNURVY
ROvaEpxe92KcLPQ7nOQebgwzgrBXutD9SWiIbzVQ5tdCm1HRpJZX9FPeMHZh
OyspuXahvP26uyTIRDndaZoqk8DXM88RyUWWGl1cxcZqzg0qn+UAntwUayya
quO6AEyjYvWATxGnHj2MSLYx1dlC+KUvHeqvL+Rmn2itbhLnSHDTnmABBQm7
pX4azaUG57ra5L/vlpUB82wru6Iwpp2bSPiqXnikZew+p5q3z1hzYM0CfTs6
n5dCHX94ZEmuT8ZAvmHcedn5vvoOjUxMeI9bvQLccFcmKTp27hsgKrOJwJ5y
8oL5Km5GLsOq4QaNXTfhUOYZBNehOd3a6CkHNiin74JFT4cmYSEf7nnpKQSX
QkzLbuM3COKe6dI7d3mj2i1I5iRJPGfW2LNq68LBJLosIPQkV40E00F4F5uA
HGGJCpRTfPAckUWw+wyj8bwf3kRuELE9iQ7J6WKdyuNJPQ9yzd7LMOIEXJ5n
TAx7tpWye32o69sZYFA2LOQsJJd2QLMwXpMSm/vHGnyJvqiw7KQdoNGrgT3F
iCrKz6J5s61rVjUzojF7Yys7w61AMyVfpp2E+6Wx76Y+B85pYYTs5OgvUJ+i
6msihaVZpkKyc7fIVDusAXGcdLGu3Fc5WYZchDMuPLxJE9nS6rU0j/IL5KSy
bwFbJf7rSkN1QP3TTJco8LIBJt1luUmopLnEGV6+7iUs8PEitEMsJGMdHjci
fB2JDKIZ086aIo0NKVeVI15dv/atkTCYo0XaEKiWx663EWqQRTvv5Y1viKr0
4j0bUmomU+ilOABJ4HBMc2lxdUM+UHZF0yc/pOb4Nc+ykf1LFsFv2Z7gw6DG
bS7WmGMeCaDHDutxW8Rh5h51yY1r6FQ6OQVMDYwfNrSNs4nj2ZjpSQfCTLG3
FUVVlf0HJlJ6u+NKJ3uoZODz++3a5etMGUkAknYdhH8RA7xBqMWwt31BIR1F
UKk+OIcnO/oCDL4CCpdDn4D20GSLcd5dwYJlmxtEZSzvaRqkfNa0eRNStlXz
DSjseSVPanjQYdaNGIrTjzbs7H8R1mtoq2DaCVjtPfwOpK8jnCOrBZ4qqxoO
PploeHj7U5wqpKs0If7h/DpJezZkamD/cqL3QaVLG0xr/nmSGNeMsruBjHB/
VhGQufxAHpUfoLew9HnvwLcB4IkC/yX236A1pkIwdIc19vK/dX+hXDhUg6W9
eTKDpz+MEN79RF9VXLIseEvfIw3EwHCNIyM/0F6UWVQS+yACKdbGgbVrh2hz
357R0DI0Tgxa4mReOJESzHYLby6rI98DDIW5nMeR4E1FXZfAj/+ODIpHRbxa
lh5x5yED3SGmZk7DsgFU23wGD9m8+yHGbjw5YsM8CnvZ5gOi2FRjHjJy5Ti/
Lt7q+TgL2dHL2q5F8yC1FaHzhkQsI/BY5RmCfCs3QYFbZ4kDbQ/aPijSfHz4
zOYvSbCJwcvnJXHrXS985jUEKkVrtO/ZNozTSAsJqP0j80gN9xWzZJDrTtNL
XZWgLruuzkS8f8K5d6WJi7iYXxRreuhduiqkXlsRUp3cHblIb7n1Wcb3vO1C
nPq9zHwir7/FhtxO9uQUzo4eIXK5w4B/r2UdBTxDSp+M7ziVg3gHuh2oFtw9
kqCEU9hv+2kDr42W2WT6yUzbFltBOsk5S7qI0SXQLbqgWTpi/7LlvBiUckD7
beNF+T3QLZe/c1Fznr/7fFA5XGRFm1n4RkZiRnBk8cgtlS1Q26z6MtRjueF9
xonIW2JupTAoscvdlkP37EbUZLkaFNE1qrBg3Eysze8Zq8QjBhr3wGy1ynOT
s9xwGWNtiC2EMW7MxpKkTZyoZMax6H5GH26ooh3qinp/Fw1zFGFz+fIAgoaj
HjKCnmCttXB/FguOwRC3RuwCWexybNoFbqyZAagraQVK/2OwsIJGLKNL0zDt
4/zcVyDu4M69HIAsowbAlhxEPgJs3Bdq6KTtYDt0YriyXsDe7w66SSHDS6im
aGgkpqrouASbtGM7pGqt0IhPqTmMuv24IKkJ2RGKLLNyHO16lErAkYjSSzvC
WW3QvwCymFuJmR3lpF5kW3dOq9N7P0KbMGw84bZD88g53A6V9oYDxOdunK6J
+BN2bth0NsuVkSjrKIrAgqm/FstWbSH0vgNXbre94uaLWMi6OC4KoQzW09EK
0xms1GJZGqShQu7g83Cdfr+gzapP1VH8KYRUFiai1prwQmcH/KgaVGB4V16h
/FVYmGMDUZVZmPJNC3aP1tP8xZ+QfaEt5VHzr5XqBzyoSq2T3AE7X/O4vbCl
l44mtylmXzQkbsOPYN0r0HlLJBRPJBVCYG3Nb4+QlVKrqz9PL617Sxm+pxfd
k0kLs1Ac+jGYfqis56QJlDY7u8ti1P5et2uQALpiVJZuV/baCyesVypMDvh8
b7BhJVr+E7827G8Thhb+GhLVf5O3eQmN1f2Q1D3Bh1zbefUck1EoCzG4DBPn
7o7ZY0FK2I7g4nIQZIICIFBnw6wwuWUz0QPITyVGNP5tPxC/NQPI/8iEoCPP
ziqzUyRxF3JMu1smNOQ8x83UcsbQcaSMOhYlWpdzIUQwDLooD2DQqQZNjaZz
ZXuFZR+5X5ueS3s/4HS/JuZBL2SGIfbXNXTRhbM6UDO79IjJ/Q4n7ptZjkxF
DqdWOmB6nqVzWzusQv4FsKrPho1VfZd+RQH4yjHNcI76XElcPdjgT4sDHFWQ
jaZbhLVFUAeICdC8Ma+FtMfKSzmxZxiKJaIIrrIrzXjGSLELhXhjGTBmv1Sg
hTg2KAgMjtkFSAuJ0pMsyorANiC+RWG72rCXuc64kByyJZTIvUjajCfF4HB5
Mz4YuWKOpVMOhD42yqXDitUMsWCgR4Y+yjZ/MPOkj2bwgEp1dqyQhJ3yEMTo
hzEaF9j6UB5B67je2/ob+LvslrZ6k+z/o43IeGII7k3f09EAjnWY6BjoN5FR
qWZ8hucuy7Kpw4vm1vlL+/DR1jCySt7KCqVrdDSpZC4L8+tkGEHy2ayHujVJ
Fh2F/U/oN9cyXGePIwPW1pWRGu9XB7Rsn7E7Av8Kkmu1SMUjW8W4ytwr0+MF
Mqznz+l/+AlbwqHzGmzJUWEtC5CZ9Ix8wufhFFPhiJpn7yWykNEbPbnFf9gY
KXdwQp9tZtFh/f/JLk687XBxqnNdeWFn8+Pq1uQpC8zuqEnUD9rJT+IWerkA
26y1jpOP4iogMf7Y6mxxufXYBtPF8MkxiRiR0vqXpiht8mnHdHhc4cIvq861
7vdvbgRxkdG5bOyijc76qyeR8OP892L1u3PPT8Z2pTIuE0x292AB7aYZ2NeT
e1WS/Vtjk5H99C/CBX4Fao73Ex04Njl1rJclVhL+Ll7qYWZfj0e/yQ4Eav8h
RC3SvKvfeOZM4XcCPg3VxuEAxiQUchueRq+5BULtSwQHHfOIXCBw0fthmXeX
0yhzbxUCP/eyPkje4iCCWQ5iZpRmnivdHrN7qw/mp0Px3mvowoiw1z1iKQR7
f7Is4hx771P17URs0n0DizaQi1Om1B40BOb5+eamXS8iJGYOdHG9MKdXXYjk
2WDAWbv2d92RQi0aYQEP98JpJmsoRT/NfxXeR8MMpF09ZQ42tThb6+7hoPt7
kD+vSM3Sk17giQFX/mKpHVtx2C+cFS2goL8Ja07mPRpkgUGq9UP4YBlH2u/D
4EWWibyaYoi0d6vuvFiLQIZhL8A6/RpOO66sakYxnEwOi/Ed4j+CebHhgNyU
3L+VvwQc0QRG5oszBS4iInxkNP+B7ubl3/O+35M6xS/fzPWqQdFj9o7TVVXo
zv1+nd5wvNRlfTlal6MfjCXZqf1Vqpr3NGW4Bumv6QM0edmcy/t2wHzmlAEr
V0dO1PpKV7imXv2yv+dvnXPslts77qI4T7/tRO66WbalbczOoVBu7JKtxxdS
w5jhO8dk1ZTjwnfJc+ZkDxw437KawmJtm383C6suu/xFJZ6QNlWKho48WOeg
ATQPqHb4jfE0g7Z8ojy2bOSmVj7c+9TCu3PDea8/m4BCRQwRykHRP2f6BrSf
7P91aO9lJkEUczTRB2XIU0nwapeOomYO9ufGFEI68p1y4bcOKwh4sSc8U72f
liKIdHpZC/gdXGQ6ghVbC1vZ0/EXMHW6JmrdXsedH+laL8OhJtc4MVju+bHg
x9f9PNf9EcSsPJlWKOoUI5BD/lbFb6QEmvk0iKFgI1moYveSC5MXt1IKd8Wq
hJOdbqHBnf5uL4Tmi88Le3oFWFBHwH2rENFPw0lvCRJ1z1e3oettaeEJ2dIM
9g8My0YDuST0Tv7ZsK9CVjj6XwHQwQ5mcEpn03jDMnIqoz3ev/WZ2FHvc7OL
fvVNRhcYaVbzO0eKBi7bnyxJCa0ndGy+69mzbSODnCm/YB0xzUYVxaxaEpYL
6JOWN01693iKcnx1z+pdH2vdKUmp7xCro4jhHRR3csfOUYq0THh4Tgsy2NUF
cfopwziFaaB3OzIjGZiQwLxD6PqRiWcv1jVw06PHC3WCGrmenuItRycZxXGS
ofCwI4MTTi1tlUuXb5HhKN3lkAfUH4lrrAJqVfgvI25sdXxSUa4U8kS+ZrRy
RfywBpkkmN3LebVVZUQLAwr6vpt8P5mSolgHEhNRTSUYSWRijMR01YOzXkHY
WZvpQOU3gi+efCj1UnCxQgkDOqyqI/PMl6yQH1/zGNDdPF7hpA0ZBL/h0kaO
xVJ4GkexW4MvaVRpjWjVhcOT+fK24ZsDc8MzxYZdGRg6lKeWPaeXUsv7ry0e
QOa7dwkUsBlPFB5rAQKR3wsZYqU602zYy3rHx5IkixszWqCY3s4zCVQ2QpRe
zMyqSE0XT0I7/ANEKGhB0DCtmCgobel05rNCpXnPIKaIYm27tTadCBKXIccj
ox8Y+DWG5iqhKFsBdHxhFGs6AGSQ7lnoN349oUisTStVGUNs2SvoNgAhp5PS
pU6xQzJvqNu3qiFqLfuoPU+cv8MaQO2LLpiuWSpwsKwqG3sXeGzi2OLJXhq7
GMj/5ZElVa8ysxAj8+JuSCzzapcgzRcN/nFND3JzNAu0LE1aBo5aHnmTmbsf
rF4Vz0kFVNR6+GTLsXXhZn9bo7HG8zqCdm+6rr6TvspkGeSkntP1tl1eomDB
jrm9c1NDcvoXPuSHL0ORSHYI+ZDcodlLJMD6+e6OaruBSa5X8kZOke3L6M/s
pYGXIgNPepHMcpCuJSObkggezzjNZkapYRDLNVniXGX20EVowL7h6TA6tG6z
jFVrvD/nQOv6sODOVS98cxUdbrkb9TzB0A0YuL86H80xlAYLvQYduc/L2DKf
W2Na6bp0uYFPxUbHdFIgDPBATSIBpkhtJlVf9ZcnHOuk9Q/x+tnZN0fHG7XT
mdWI1hz4wG9UdmOB0DnYqx2hlKfDEnyeGYz9TlHjtknEoGT4Enp7BZ7DXWGK
DV9qsgwdn4Jyb5qKqic7WncqZyWy946eKLXA5RoZ/0BgCIPQS+nXbNmJ2t5s
/mhfu+RFSI+ko2EWr+GJT933H0WJkYGIgdAvEmomkTHzfvV9aVMJnEaHQ7KA
huWOML/2T1A58ZKvJux4579kfF9EwU6/tzVyx+IAZKuhRLgW3iJ8hNKoUYdQ
G6OOKHcXwslqbReFghtTdUe/0b6nlCIzdHaHrknacV9y6z1dbubozcAxdBvZ
0SXQuwnoYJBx2w3joTs8DQNPHWx8hC1zSU+0mrUg5nuVc5vllcpqplWO7H2V
0pwuSD2gUYY/nCIWEH6CkdvWA5Ih0oL/4WAlJxXd2l1hLt2LZORMC29eSpvr
yAE0b/4bwBHJZ2avQAwV0Uvp8bxkPVCzCKgulr3yz/RxTsphhBebuUNs1ycF
x4fCFcSzyycolRWMxFAjx3IZV8MgRyfOHNa/EPaFd6LWl3UVWMW1CuAt8nAF
ghaBU4ls+GK2EBEedL+9/bOcuV2/IpKWtJT4IQKTYL2QzYbdQISlVDj6zeQq
/99C0vp/0Vt6UL4k3tkAmmkgx+I4c2igEOjHI/HDxft5ES85ELeYbXmWHzNA
jfSG6g35sZRznjLUsNjOR4fBk/uquM9ItRGVJgqVIBnHN30MfxhgzaW+gDqS
qc+4oFrEE2Dd0sZfTCu4FINiOG4Q6pNt6haLErHAeJgYYOaNS05+HdUrjUu7
Yb07UbCJe+46pQLk4xTALUUJrAXno8IRhMiGEpUdUBM0xOcl+El4J2te2kal
jHEUYbWvkZmWlCRZ5Z5oAARA95F1s5GXqrIb3YrFdDXYMw48H9WBStsBgT4i
7iBufmu7zdcN90/nm/sZnoaKg6fBgjaB6+umGur6wUiZNsz1PrNHlG8zf8+u
6yZI01lQs58Mv9gmCt31kL1mNQPgUmq4tuv1SUBmoHQruE+2izh4ItpnhlNY
BCP4CuKqGB4T2o6fvz/f8N5ZUVpCgwJbJ/t58Kun8sssCWjuFxWAzs3WBDlI
R8vexbe7dCdLnGL0KQiO7QW4DMVUFwAP2WMEizGV8iyI4nlF0/i8GCxl/RdX
knrBeW87fn2dmi7viBRiXFeRRHYvsPWtFttOVJXkqzS2lqyz+u+v0mJnn5Ui
LT/FSkbMktLtTwM8kyk3UMd3mqOPHEjamNwl/yfsgXAUevT0CmPgPAmBojjt
9oic77al/jFx5Itk3Jg3AQV1nFn8sSAJhlp5a2qURzXE+3scnCSbgGwf3eIn
0tUCMbiML+EorRVibTAZCf5UHq1uwl5ZpstdDXUXYSarAg8pLwFr78jc7R0O
XxH1TI1Y7g/YMIsqTc64cqIHIXAJ3lta/Zw7/Ts+zm83u66vesCF6Dzv7yd1
weiytaSC/tP/ajuDASBldTaeIElgHVu8Z0M/80fplHvHUeCAlR3c+xZhShY3
64BOLMTb3OgzLKLLVYhguHHT65V3WkDKWOajCmWBf+39PY2KLxeCcH4tyd/h
hX6bVCBhVO0Iri5R4IFxCG49l+gLKu9euUaZCplzUvi5NDEEVzDRTBDXypp2
EahjQXHc4GJdz8niZDJknLvscpeC1dBTkOo+cFMMsgUD/nWs+x2dvME1I7tR
NPVZg7Foz0NNNRvaNQNIGvwml5I1RVujOOFv1tdqyVoUCujTn4aAw8hPezWJ
IFhzA285gJUGjGk51r+HYl+V/0lKMUsQ7SqeJQGaMJ4nji5cBgjwnsXwiReC
G16WhEQT32qzj8RREqvZ7UqvKC+Ca9+P01neCbffeKB7HiHGeCeyxnwkXSBL
no8zXZc7g2nMLLyfB82uZcxPnVLSv66l80OOQF2HNFbqLiWU8h+6zkmlRvm5
nu5CmJuJXqtY9ABDVStAT4dNDm6rf579eEs3Vv9VltqgLacpYfeENGDqtnl+
7p7O685/YB21a+bSi8Bag9y5rbpAlhAXwVOVRQ52EQe8iap+4ccGBKH76YwU
mqpUnE0gMxTdtdzvqbGMKv50KiEArJco+SZk0rVnv8fqb307S7pV/Ky5mLT2
mrDhUV+KT5pC5f6TIilapEKp+yBgWHQOBK4ANAjwQiAIOklHJNBOVCdF/gg6
b0D+cV54TWPoHsgYZxEu4s+tui2sA4oqM64c4q5eIx3My5w3dYaCYZ8bbiA0
kPV13eQbjlxQ7Xl9Bdcv9qYTaZACYqsfIXZhbi68uXtcERFyQFyVrnij3dQ6
C43qKGkL6KxynHVj/0lE1o0a+QJ+oIzB9EYIvIiHru/FCFbeSEtXylULr5ae
mIKFXuuHITQ0GbBR2JK6kuhC9VNmlXCJpqZZTmaEPrtlGPxAF4c40LWSKVaK
3fzifoNEwnL7dtW02NLw9PHC4fVQedx6od3JcI8GSV3n9aRZkApln8Ar03M2
fYCoT9V95CLRXL2N1JTMuhjXrJAmy9C2mm53falgWz3yp21AwP7SxmD4Po8L
d3NPd7y8uuQlfkgZq5t9+GnlPtVKbOJWykTRvorEGNnpb5BM4TCT5MIO68O8
B5oYuvuR6S9t+dYvQuUpXlReN6LwEy7eoBtVq9ftuxcwVzcZLOY/MLXvjqWC
NM+t04eKg+a3jegXq60u+qYsLN/bvjFVWDp6+tRxubEirV0Uia54ULpbxokS
aJIb6wPG2eBQr5CMJfidiqeAxPHzZbNLJZvrfS0KMB0YO5rP/9QXDBvObPGC
vhx8foktyVwDq8cdl4rE74YY+093dbzndkFdR7uXYIYzF+2DGNFASoZ5CVkZ
Ll9NWjKP40jCBnK7eToKdLjNitPMYNmXKwnLv2T69YncfThWLq96MLh3RatM
SAqkb4k4oz6W6QNFt4+e1/MCwsUxO1bXBlHXK4s+6Qv+i09JKxpmrZKb7ZTL
+mAmrgTYYpRM91cdW/qwUBi/k6hyjSedVPdldvWFP2k9vZsIi77wxtNT2+lK
Mjr49RBAm6ra8Cqkl3ODlDYG3ITd9IY6YWKtsF/GcFMJmY6v9c3nRcEZ7L8F
7T6OaJC4EYEjedPB6dEBZMvMG2l8nxxS+8Hw1I0/4KEtXga5OQrDoaW2Qz/d
xgGCtb1bVW6+ZUH79lkvMsxYGUHeOttv19vua1fG6Y0/HhBX6tYCkT9u4xoG
zOMxitr/Ia/kbphnFumm8/KVXsuaB/VZy32RSvJlV9nH3PXWbRhA3krZVzdc
Ml9PDczxjDq39aXeXX4fxFyv5xzJEo4JfqdkUC1VPBkujQGz+yJUVKdczNZz
qGBok1GcnlvjJOOeCiYPavMca381tRzr9sxnxg6yR1M4i72kl9dxKaw7hw6l
ISP+5MkZhg74mLNgWNJfvPFTGvy725l5TAOHXh/Fns6dlpzWfjbBlTHmwjmX
If8JnGaZk8n7NW5opIOdq1pa9jmdg9D5BohysPD/e3bdM2a0SF1K9bybl0vY
exHUl4VT/BynYYdOl9yxrStze3JLh0tb9PQcm15UjRf0z4gv7C7pcVQrKorm
rO4b5kHp4dMfYsCcLtfo4wJdF/suySl+kR/1Y47TGFFyV4OYk74QhJUnigUB
f/RQw+DXvkAu6dRAaPx/6Guhl6764z43ruPK5hpyP1gbJlynBKJzVherHbJK
QLomWa7XvYhD5MSVOVLj5furoet3IUEzKCKm3g0+5VzXBgquvxDjF5YtLs2L
hlu8k0nZFjCQ0o1KKTXFr3+MZ30KXjRL0qlQ8vY5br3P5dZ0ZIlvWdvCVnaj
BEpZaT7MWSfRqUzgPb2grQ1LRvVMr63x6FevGmmWdL/UMDKkKu+X1wZjQ1Zt
TpSNCcd5i13FiB7AB2apYnWUpcS7AnOwgBBEr0yK4fvvbBk72wGyTIUOayju
/dAiFpfVhqaUav+K5GH2ilJu68qAhSI9TxVKUTZMVTPqjPaDVUElvjcugldO
6uEVcBA0Nmrm5A/2Da88sm84kcR2qcpQxCIWP8lBBYSxCTGQxHrqhBWnw+Nr
uyLLs5uB+xOOvmsKcL6qHEi6OmmUAKCMio63+tyhKEbr55YnoB6vTLN9B98Z
UC5eVatN52Z4gWFYZVGnk6dUBk1t/N+xiR3URbpiweconfDFblx77LSow4KN
fbs+vfQCHMYz5NIB3nYPhg2caRhbrUYTm1j2DF9HqqT8ij/1/gTm1bVrNbPm
EGgvTrRlVG9dk90tuWZVDsCAV3dNhWpfDab5Yep6nMm+BHt+OV3vjCRNSWEU
q1+g7mXI/6YhX6UnLY16KmzplKdN65Jjusv0vIvU9LNWD/WtgLJQwypBipw3
G55EYjnloG1IIMv+9PYwjW7QokUk7uWNZt4QSkv5qoC3Ciy7psN6lLWCW6T6
a69UHZ8pxB8Mi3HOpBywTALcyksMa5bRANe4Jv2dTAWdyZpvZC6JvJvvo7h+
ABs1dwis83HuFMy4+tT7+Q4aao/SdEpZf0VPW2sShBBZlHv463Fwy8K38bzf
XazoVTaGmhgJFvfUVs9xDPBZh9kPKv6ew3+LBa/+7qZRGsAfVc3oj7/GW5Ah
Sa99omCeIi1aMpzyvkOXu1Tql/OrJXS9z3sGjWkQpj2Z620HUp/Q41mBTqtd
4e+6+ZDD0sdWscgcfszsyeMcyYwlE9C+RxYUYlX3umzklgoO3XbwTNRVbvHG
WSN4U5QPWbFsiYQHFUvFh2guka3WPYpu6wvldNv/ve/j7dslrvmWmj3m4jyc
BgjdShLRBhdNU7ZcKA67B3/VXhwZ2QQbELbLoZcn1gUdjx1qQefv8akHa838
HB+brUO70vrqxc3YSXBWQ5yOyDFcn2vTjO+VlkEPHa1X/zHOdF6edfWgyoQB
XY8dK1kXMJH73JtYxsB9G8YKynZafbgF8aK4tqBy5ydr6enTH5pRE2sK0U7p
j1G1mqkCvkgKiN3SUfCv4rGzTVuP61YaEGS/F0z2NAJzKfTKK95oHRzc1qyh
wNNObL8NiS5dlr6bASpjIFxS+D44XHRx9SHMjV0lv7uuHORi+LPKRAWkWPzg
Qde5cRxXkR+3ZPwEuLvSIHa6LTmlqNl3lOjg8LUswnQqrTdL0BPArmFcnjjc
VQk+Wt50ujSKafw2mVnQfdRQjVK+PVHuZzjKexHqFwNOjKIq2Pj+9uexh7aD
eWvtHtJBy/uHXSI2JAAE8g0Vw+mIWcng4QA25lBzSPWr1FhUsvvWbkf2wMTI
sWcGkSqPPb8PCPVd3k80cYbYRcxDMbJzXjAOTfJ2m4k75tHeWb/dhU5DUdpd
y7RL9WiZLoZpZJiKE7+Ht3zq29LVpDBYtpWUP39k9Wb06ak1YnFcAABwe149
S9xaJ89KYVdZtJlBvKUD7NdTEAAdSN6wDW05nmuBJbO1wJbhMFQshiWyL0X5
lrtNGelLzuNaH0xWV9OhHqoHD5JKWCkb5dBjWOi5T6wQcC7TbdDZX8jh6U/I
olFo2oFcfnz2cmmXLta5mJbqrm7Z1hnhKhGNLsgLdcMdinSu8TrHy2y+DTBG
UTJmooF3UOXynHsmhuGq5VyFuc4Xymr6TgesVmCUYM713x+aioV9NbDGk6x/
kQG4wGXO+57K0NyscNix/dcv0gONUfUiC0Rasx1+WKTX7URwla2i8gbDqkF7
aj24DDw1Phuf+X/21kX6gQfdx1o8gF987sCKXtOHowBO0UHnE6/GR/VwOJH5
L73I0LNrY4FmzxH1g4WCVIdDUd168glOhKLuKy+RPJBZnipUcRg0u/tXsUu4
S7nAkN04koiF4R617BxAAXqOaNdAG13fEu4U/tYtaia+n+ZIhQVWWGZRBG8I
UXm4FjcoAYxVDGdtly+BwdFufyL0KlHQHG1VXSY2So3Hhbt4aiz8+sZf1fuA
ASbAA0LKAOZ6q3rcrtap9fHtYStZIUjiOqdPhQ4V9bWZ9l7lDJRaXdJVe4HW
F/GiEiqavS9EaG+X9ohEIFamxK4IztCrA371o4n4puF1Cga5v1WEia/76Iqc
KsNFZk3LoAYHEdBfk7im/KCb+NJ5wniqN+iAZ/TTbMHuJ/XSL4WgcGlgAYfk
JcHKEhW1+/bDp6fT6A4cuRqsLPXB39T/Fl5awdHN8aDM4c7+9hKsPFumld0P
RfSFNrAUh7wcL3k0EtQcyuotOLGC6p0525tVeOgGIat+oflVB/q6J6WluFNg
Gw9x2YjyIILNpE4YF6BOG7XuPKBPkXJ4Ujn8ud0jx4JfwP/NIOicu/U5fFvs
mzpUAsDhfUqq3E1d55hvAjCm8ssCa8QldkLtaSnidRDqkTZnZ3qR/sJzeVcP
1/uOjdl38nIEUwDWtwi7NuCkaa+c6pFia6VkqTcDp+SampRLPYfXBkVSFizL
oLVgJrcJS8EFPQ21obyUte3Q3V/g+BfpqfJgYXxnr6hE755xuGLAkzQAUbIR
mQJvJvjdpQZIUKQVUyCsmbzXgBQMUOmamB0VkiEBgjwbeHDJ/gZXR3YmTrau
LGcJz522fYsfkIHfoewC9ESz3/95u57XBGxGiko7hlO5PzRYPvPEMalcltv5
aXf7pAVQu1spVDoRZe6FYaJngChmXzv1YrnAH/DonyISmFx9kDB8mLC/scEn
ziGmuCXiYCEwvevjyJqdbGbAyMUluFqV3S0PC7fc+2/+U+suEcxfsCHB4N+K
6FpbQME34hXrRvP5Uck4H5e7dOM4Sw6wJsWH5Cao133nURRFokEQbQcW8fj0
XWQOzNuyEqb3Ix33uZ0+OW0HH5qM6fYNVgGroj/RXdqQyhH9Z08tbxy4qm6U
tQuQHnzogFZCHIxcu1KjyHZNfspXkufR/xDsBlbacIKJDHFVr/mwUEju08D3
5vitStjCmD171zbrwI1TfuFfF+Rr5g+Ik8ObDWFKHML/AEYJ4sFDXMkjcT5r
25vaUDzUIIaK3Vjh8i/UQVTqV79melO7kzZyng7XXDtjrc0MqGY9uf38LWf5
xv85A23hj4g4owazOF5zmX7VgnC/y2S28TcMjBUZKdUCK3KUAs5w72TZLOvY
O2/USAT0/k0oN2nxCq/YHXzqjNgt8eVyBcWR2276i/YqAlXuPOPGqF83Jc1k
ksNpJ1XIqhuenLHe1Au2jyx/FmzRYIM++YKv5i/Wt3m7Y50kAyduxqaUqhGR
tA6yXTDEQf4mE6JTcI+TgKiJmztZvzA6hKrxIk+M0LlnKAbIwHEMh5li6AeN
NPMYaOH5nEvoSa+X0cYXJVIAu5HtjnajZODapHUvUh2rqJ5kBPuvHPubg0Wg
muGBEiuR3vyY4/axvfnD74iXCb8jGw2xGFg1dHqxO2gS26mjE2ZqeKtcByda
dYrr3SWzVGC47XonTiyUGpjlyf1n21cb2QGkL8/LJY8cKYgasVj7w1S2LXG4
P/vsGr9xtNwutA1H44MOcJ13qTiPCBMCV0k58UiawAOcEObxW7fJys714GE6
Sk4QGuZkLZUYgbSKD4Lw8CCRgYpRavxeTOM3eRpJvoyA1Agdtv2nCQBcKFgV
rcpvkXfNApgPxpGBUlkwoFBoqrSvXoQ6VS9U5QWNLu2voCgBY7g8cWMiuz4x
qN06Mn4Ehg7fWKQd3IqdeylglhsjTAXxPwmKeaA/LPS2uKaeUs9L/cfJxnqj
zANQXn91dG1OMjscQC40inY0PZFhCeQtaKmMbasOV6xmfHRh58nzASyEyv1r
4/FGK2R4zaOWsQakMnNvLeZhytWf3JWoqAmbI5E/JC4EhhJ6056ljqo8PMP2
IsTO6exN+B3pr6y0Sxc8qFsKFZqcBigiw8Ffojd32fV8zKIxzwBxX2ZlgsF3
a3KTEgzmUQz/xASt9W/v8Ajvk86U9skIRmKNS21EMofs2wBINQMy82rjmTSL
aG3LiKsm8bzA+EhTliBcYGWLe6hRFpfkyz2L5tVVqgf7g8JtkQXsFlv/jzBV
KwDkr2RQxjNkTM/jXha0D8FjQ5CyKKlHRaMQICFHFq+nn4thXSe6LsJX+86W
UVI45kut1U+oQ3gS+435ADUIrizVhJVKGr6qEDBuh8kpUoU+dS19lqpnLh5n
SAmMPy0N5CmnVvls31+6+akrwyA0s7W3nkMfxSuxRtt0uhFvLunTrrFOH+MC
N0GnYdvLAZH0pEHmLZuLFlivjGGfm3lkQpMI3qNvyxqkC79vViDL+QtYCe8Y
Y+YK113zv2kSfOqQOPbPHC1bYtZa7OIRu7Dr0iDrAI1q9igbx9flosA2eYL9
qfpHtaJSR3Z8lm5dslpDP1adhyJqY/ai1lgsrlkdUhFdh++QSchkg6PhuiHl
faiPYzxT0XROehzveYDWjmbx+dIzt7EkcouTQsxoKMnEnOjyS6B2CXgnvtP4
lV4CKNntNRVuD6vFVvynFXFNBKi6xBmYwDy2WnDDKvoUhjF4bzogHSCd/hwY
M2r10EXe6Lw9KVzsQlX1JVrxBGwOuhrs49Gk6PtgMVOdX7eHpyFJJdIUMZJT
5NR389URBc2HdN0f0L4twaynY4QNQjK/2s0j32Kyf7bwKIPqVI6Tx5B4v1B0
SJEA9+CrXD8NQISGziD/2YCSx/hifE/M78WlgxC2gHW57C698gdc30TzNgA4
LXAhISMXFtsIgU8FaDnh+GwkKZbIcq6gbOnBBDfpa27gPM42iBVgXzmqAzXX
BHwppTDIKEr2+K9a1jL07QC9v0JinolFKMUFFZoyzlxyae3MSPgaQ4U37m4c
/L5S2T93AaK4vXCJVpSUr3z5RjQBXiZ1/Pou+apSFWdgYvPaocyUwNAHSgO3
bjhbnTDc1u0EG+HHZcCBfK7dQwrHR32dVncRCIf8nXFTXHXeVcd1vW9ClNyX
cfPbE0nTgPTCDQKiXFH28m1cIkJYvXMQ3w0TjkewQgEOdiIAisz7R5vMnCIP
n+yM9qx8RCgdp+5TtSyOVVtlD0H4KeK//P0WFomJI3r/qhmRjgBoSAUDCJ/4
GFdbdEMyFt0xmAuf2pGwyD7zwCPe928QnkamGIQTsGDqwC7tQTks/mKde0EM
9PrbNee2h3slTrIHYUmV1tNMfU1T29ef+t7xpP/LVHtfkvwAq601zv0s9RpZ
fYgrXUZSpKnE6zkxMGcy7DDAecERyKdBGhah942Vy2vMh3p9i9q8bvucyxIv
nde190OsmoIorQzlX5F+aBac1S3vCZZBmmAcoW+zvnUf3IGS6gB0xSc/Sk4G
0uyV6JNQ7CnnusNxNF70imBiHWYJiiWRgkkTPmunKqJuKuXgl05KNzRPghzU
IG8W1hFODV1J6Gl006dYKNgkMSDBdR7UQbRJ6Rrb+xY4wBnzOHdGmtiDDd6Q
8/i7JbO2mNijOfXlKpb+oiVKARSx7vPbJij0pFa5EN3tRuSGDdJTsq+Q2ePy
86454cgyYiLv1Nv6IbEpYhxTjjLojAyg0SSBwwdYCHZxjSzI9BvMmC5tmu2S
iVI9JiM1c+cNwxC5W/2yPWGthRgWvdAJAEUQlIxdxR6VBHI9fjymqY1yxi6A
Q0EBgGcN3PI3Wh2cqtLYwGBrbi8edy6SjhKOdhxDDXMuui+B/mI3n1WIXdic
FS4xka9y9uVygV4w8GoYkx8yer9xevhbJTLwrV2NWIvvo2w10vG9tHdAZAs5
5r/lyxEZLnaKnvEoxx5Sfs0NXttMQoQqsNM4eGeknqseRn0tLU5yOubHzw4R
qbx5e6nnN6CsvR1yRNAUsTd1bbTvwMlq8rEUBqEueWWyC8WO9l+TiMLoGwo8
A329OEQf9lmGerwsJHd7coSHlG92X913oEt+b+plzJ9FV5FAjoeN/Zgdmpov
Lpg+yhfcJiHUMhYuyA57YFh7k/xiZJ4a+8cBa+WMdDySKqNoKF0mas4o4jdv
B9v4iX0ESStjvHDmKx0g5qiuxkBuWzgltZOBmEldC4KRXaMb1bj+cg+Qj3lV
BhmiczPUMGF3T67xVprmlyBa45KYM5NLbN/T3j8dNNLxFScL9X3gKv4B8FoF
FKMbAeNf/idmuK4wXG2kxflVOa1k+jFQH1njKNpN8fqXHMspt2zdYoCGQBZS
m9eqfl7I+Ys9wGDbDw9M6dM0pcdtkM1KMgzzWE35zjFijTnbvfEuBftDtRU+
8pCFsy722iaRpRX3UYbe1Po/fY7kQL2IHhAKOoQTzCqdhqE8qSjtPwO15Psf
d3EP0HljP4icwlfLYxnXsrD+XgTFS5mvYIrwFpSut/QrVn6uPcdUw05Fk4Rx
kVAQvDuphHtR/dI76s/ovJwpF1Ec66HCRDdxdppJhMANjS2BbvWpqe/nJGZq
ajMkuXzme/wEIAzCLyXX9Tj9SVM5RoFaaFFA6YxTxKhuekdvIcty2pyVIiq9
aO5yN6xXbqJSbp6/c24Ts5zsmoa4QMamDwbffYEAxOJ5gDw5iMWgpGQvX/ip
XczoWIcnNOJpDUuxzT335YMdidX2noL9TXm97koxZ2E2MApiygakL1wNxTk9
cqkod2e4WMAfPngTQpfWEpCUru9JazRkhLUPS9OtPij3MExXPLOb/3+hVkHA
Iu3zstDmj2qvW4k23AoympqpsLp+sxljE3JNOy88GI1rS5y4Lkm97+pz7CUG
gwigTE5NQAq4j/mtwURXu61DSIDw5ulMr6fbY9xFJDq+5HmXKkm3uuClLhWr
BlLHVaAsVQxrO1ObIOEu1heqhWmgBCJmkOYirz4bZz/1bz0sjXxw5juw7Gwm
2JgFA6wngXnM90+hyUxkkskPRBwwq4wzdFgPIplFihMLIPSYc6NHYUZPHhpc
tdHQkJ7Dn7FNIqbZBbNKJ0/F0MeEJNXDQafJg4f5zQZTtTQU4kIZQjsH9ews
EkV/QUjLFZOsI49pLjCqn608yJvqeDlrcSqRy7RTk5Lzf55J904gEu6vTxK5
EUB3KcIo+v+W/LPRIG977dyUAp4Yjm2pH9QuyoeXSd1c8ps1NsYFZ1VScpXd
vUcXwHNoOnn6K/7ZGgExG0QELxuLw1c2QaGPelSYEdYfT8LPL7O1m6WRHQWO
11MKoK2PnMHTOP5jjhvSiz1MVqIum54yGy40yMEWU04ZKBCKwaTET1AwER2a
U8CoCI1cC3CdMVYUb0O26BlM/GPFe0PuUpgV9i4zxK+Z1CbcaO+00yQK2IYD
UY+1y7z4EEswrUBqhj2hBiLRYsw6cledQhwBma0JLeEInxyP1m7oSclR+uiy
sy7EygPa2NDk3cDPNzwHdv76gw4+3ztmVE3OowOJYVZrApt1TqOa5GWa/dWj
NG8Mb6Wp5Lf/dzXJLaSdPMvW+tddeopjltiZoWpT3gS2wdXMOB1n7aBEaDXe
YD/X1XQb9z4QiTdFvprp0b3Yv7wr3+/JwdwwxJvMMbabl35b5oNlLje1fm3A
r5jZXAjOkBdkDbTNodrtMyVn0EmaWq6nEAYwcsyB+dgfDmoBcjtIYVfJWRhO
3gu8qrzdf/y/u9cfdYctoAejWMGuGRzrBSpcRlF4jyQdLhf2L2xzeqk+ot/c
4Dpegm2AECfs8S5/uoE+yeAunQDMbodb8a8NKsw8iEZVn2cgzFYcL3hkr5+C
bowCnlAWjL23Vzkt2uooII7n1olzcZeqQYq2rSXdHqjO2yq5+PYXB372a3EU
zrMxHAYcV6q+1jufA0hZYMgQYrGNt6NzVfraqn+gHGMzOMxtoVJRHLVXa6pP
Rc9l4pk41L4HpHd/q/OJG7Z/QryspfH06M7QTjarAeLtil6xVPZ5Fv+wjKQO
ItEJBdezeSMiw8prYF7b6VO0fw+bCGCZdAvzIBfSZ51XIQB71WZCkMdWGRSL
RzVDnRoJ0msOh3yHR6VjgDOAbh1WaeT7G2uqDnVVADdA7AoksUWoo0vPN9lk
l2Dyg+q9CakgGh0c31/UM3FaLggehgtoc8WIEp1/KIdq0XiaPjjx1Yj3TFzQ
GhiAqPl2PfecIhQe0sxzDxjf3cqTqxNj7Vu1TVlFAkQd37852OA9HHvea6z/
jEfaSD2WjE97WE0Hy9P2y94l95Sf9ksPEi+enp1QBnjxZUUZRBVVgo9YBA1l
irjaR8aSh9P6TGC3gUuDc9P1gAPhrgn2FBAqv9badvm13+pojTsVxHyc7YfQ
bYIRabOnQkq3wDqI8SLno6q063exn4KmkZFEmdNP1uNzx5rmHcUTLatnJjzf
OH6O0oBf0iAz+DkuPU7MCFZSzpJp8Z3TqMj05IVggbHUL+LEQ/uwXCg+zMSm
YU3WfaVho/qiDxQV1teGnllkoZvpRJBGCEIMLtAicRzWvP15wF4krfGKUyS5
6OZOnMz433vmdbiO7Ghnfb6phkEXXy8/KDJ1rjutDmFtbF7CMwTJSGkb7/5s
BwRaLaZtBqCBX7tlnHeMcbc44CxxHmNkGVmiPPh7+BQoeVmqauC3mwrhM6Ox
i0X6Ir8EeOMe6ePcuAjPcyqRF+R73Q6kDmChz2001WRXEz5/Kn1ExVjYHEhk
Judn5Rn4RJ87VaQZc5WGYqVa6LkHeb8Rx/mpz2t75XHEstv3a2R0JagOtLzr
0SAgtil1DxkWdk12Q+uAGyJZ7T0qHjfYxhinMsZvZw8nyoNh7nflKNxT2ToN
+AqcOo1smCypXI3Pa93DvZf6Ibn41nhGqFDouJqdYkutBFLsNTceixI9YnzL
A5LFBvKUFL9sZKqNAr9AqSQzmx3ZJiUjT37P0bvljtgmoTYVr3z49JuvZLI/
aVHBMp1KyPBapO1M6oQ1nV1uJcJMt9nBH6i1FRvc0uSUzZWUddfzDjakIvRP
UjeAtssl6gM46u80gMlZPHk9wjT1VMsw9UiKVtIt57ZVi0vliJwOhA99NvSd
gUC4ATLUI6wjeGxB2IgAOjam/+izG4+eETpZ6xaOlJ8QJ4sA6qN+d3uy0KHr
siF+ElBB//EpOoIdV9M/OLBWHQlezMb3PeTch2ztQosbZ1YspULcp7msNeHY
gBGifXv0tZHWCHxY0NT3i7v6qiIvrXVGtFMQITl7MEFcn/KUj7iJpw9szIe1
5ozimuSjxOZMzK6ZVShh4ainipprj34RoPn80jzjv9rPprEXRKOcYJb7qcPx
3/LK29za7zcfxIomtJKIS4HXOdXg9NWpktc8p24tsB3qLaKzAqMarP8z13gv
g5C3IVNYZeDL1YmlS2zEwjUo3v0zOVOr5wDeRRCvABYTT7GqYsNTWZtVEUR3
2SJqAbJZfFFtuZd84dLG4uTvy0fD65ArV8zXjEMtmx+px8uy0J3fB0ZC+vLZ
Nciuei7eURCoJ3W0dcTQ7bA01IGCt9L5q8rdNTwHlPbH8kxHykYMw2iG3nVi
qa/naxn7P8u3zy9LownJ6bvMnnmpxrmwbqROXyy6kwV2W76pPBNfLXRBL+35
Si/TIKgWLl9rxuxe2SaHmc2OUNjBuXqrITUjaecuCp1c6EKVpCDaaDF1L8go
/K5OcLCfCFTgRI4L2kcqXdYVVEB1YeRgcItr3EFVnelx5Nm+/QkZj7AF05KK
Qgl1DE9XU7Vj0kg5XiLFRZEZw2UEln3fqmLHyC7l/WtrbKaGqcG+76LwaLX0
A7bRE8t2F0Lzr4HKiIEEf/SNlndtfVvi2L9kRiy99x9lBXLlwc3We6p+v93x
4hZqGWQw3RvetS25k8MkXEIDdZDQqi85MdLbBsP3hoyh3rdZsC1DiWEdrqww
nPugk2apRD/1o7ZCCEESb50EHP//ufAL16DTevwDitMbXSQlTmMqk1mY8mv2
WMprfMFvrOFXQv9Z8ucQBHRBGpHMyUMYtrLfgw0JFtS5I0TQDFY0uah2HS9z
vNqdB5Weo4bTOmxUGcqvb2FiALpniMzcrmncvuL/ErOX/ctd6PqNhitpxdBz
EOvGeExyb8Oj5RNt+yAADIQInXxwhYLa32pmkCykW5cpOOUtN6TOcBS/Qfvg
/p0fpdGQn3Ruz1DUboiUJNU7TVSYpxfY9+fEwRfaKFaAHwj4tnDcewN3kQ0N
Ez53DE2ZU+lSjTJzMNwHAOEibqxURAgONtvfZGIotaxnRaPH9hvlbX2Jdycn
cELXvnSYysdleNrncRqJm8gjFkPKNX9Z4UZWOGtOrIIWTbvNqAxipKPnOiGH
8nVeg+OWPYBGY8dkjQKTGH8fPHwQtfbQC/E2XjI1RqSKwmIZze9YPH7nNyeo
wXyCzG9w8WsanGjoZuPE54MOIo+eCjZlL0KfZ9Eb1tXAWTBvN3+h8cgpcADL
lWTdqK7N48cMhg8dk+c0GT0yAurWn465NbIVMTe7s9x5x7VrIMBurCsXJWtf
DNGP4hloPb1qzCiWvHUdXSqsxrw4waBDLjlauCYo8HtWLEAjc6bVG8s9GWqo
t1vwlqTIoIDEHnztwsL+FWwX7x/YBh75VP3v9XwhX5HH5gNaKFI1aruDE3B2
o3VNVh292T+lxda53k9+HjWLuCC13f+sd/VMfXCN9L05xPPxYkHpdjf+qL6r
N2P9dg9kXIqfLL3YErjKFRJEJKoiTboAmitJZ7AaafiexNeSC3iED8lczera
whLIHED0IZE2SoimDVhl3CtFruZbXRL27RPqVhHfmet2HPVncNjZrApTwiw4
RlMl6WolXFY/WL6wd09UzFKPky50mvWJFCjmaMc25eLbOzC9/8zkOROYcaIc
adWz9rAmkmvvthjGWDnLW3UUEEi/BKgYGUExyLlzINGAeu24EOVmcUO0q/8M
eEMoW7sZL7V+Hk46rnM+2z+713nwweoBelOOrk/iCoeMrEZUaHzgog+0JQFm
IytaVHWYkhuwU2vxDEnOWjvD9UcHvYzsgCIPkdHpUpYL4qDOnGamcIvwqQOL
+R2xCwYKO6etMDu4y9GAs56cFeKDDBitD5ykPq23btgz2gezo89fH3SM5GD3
ct4zaPL87zXUnmLqkMwfr0ocJpCekMfL3/FmqqyAX7EhS2RwyZ92uhWmPvmx
GZ5I60XpGjgpmxEq/L1DxpvoDoMe58oCWdOQPLFbyyj8FSjVqDbvol+Po/nd
VtTBn8VgYbjjRKM4iWbg97xMx4GfHmnUkKaHwCLAmqD98/BpsO0ca+Pu/j5X
HagsCv/QRzAaLa4pHPQfTfs5Om9N85xyN+rdwz9ZGoCzLkGVx6EoHBTVtaE8
QgnhqIkE4woVbyDD7PFEwBsDFCafzp+cW5lV0GWP7DEONC6+P5HeaC9hkmb6
/NCIhkr+xR5cXUYsp7pxlRwV/DJTMNAXnGN1kA74ey65dYIBIoHEoRm7OyRG
dS/uX5bQhLcz6LkuofPbIYoxE8+jBYFE4IScGmKJ0HieyiUOnBQcHhFPkVHE
4Un9kCkluZGqWH2yrqtV3s79vHaEQj6kkhbrVhPQEs2YiTAyA+C5Qkofo8dn
YNdF2NmEvtV7cGtTZYtH++QlSCkEsRLg72bDqRcBOlyVTuIlUyHOMPwPIWnJ
nRAP0UBkxLkHnXnER0WoO1Q5YWYt1CS4ptz/VIMcCGRe7u7DQcMPlPTDtmZt
Wl5HXM/ad/XigNTHgcdi7W+AYb44gcF4Gck/shPtPkV1rM9iggKguDvW0OuX
rBdrZp4fmMvfO0auPslno/gAzW4YaKembZE2IlivKax4gIj26Y5OfwmArPSL
0BLGXptah+MUEfrIGoXYRB08bw2URRIZy7Fkash+5shxgGB/f20p8zvzf2WY
V5J4mvFditlJrqWaTalRjoMkHEvYvAThrzu5tO/pzrujbgf5jrpvAnN51zwL
LB5Bb8XEnV0wQutMVmT0OJUIFQ36K+Mu7DucLZmmsJwGX441dNMZXx8K37Ks
kTvM9y5ya5J2xzV0xAoDKThXTc8eoVrh5p3jrXs8RCJMo9BmS2PYQrYlc3Qb
4uMGuOs/BXx0Mh+MlqMzZTKzFTHKT9MtOOuaWOQFI7C9PULLil119bIewmkd
ax5daMq/buvdEcMZEmjmQbtFcVjMYWT/dZPmEkQ7iipKW+elgatpo+vA+cJE
saTIi0HzQyFtsWwo9/r0HzCFK+ytwxmgSUtuIf7rZ1HwUs+F/lglC6DUJthH
zGQ4BSIWjANjQg032DK1l+CCYkKzMx0hgdd/7uOyfUUDX+NAj3VFHBVVA0Ez
Ib9Ao3dYg+0HUdQLgAh/b+EK54slV/bedxFke9x/6TJgy+YPiI+U2IRORrQM
t2myvdhFgFHOipT3Tb0umS5i+1ttk1xvtGhV3f+gCqhSR6AGLvpNeeD4jkrH
wAam8eAMwtVl144EmKTZYx/yfpsmbjyG4Zk/0rxgwnH/sm8GoJzAPSP9cERO
+Z8WuYacLrEeMbwZ4/jdFhvsusEgcGgfgAUloAoi6MAJkM6rHeCM65H3x3+0
9UJWT47CGpyKrnWSNe/2r4JmCsH4NzCysgNrbPmqjQk9mBOMp3MKiDqzm4wl
m1r5MdxGMH+0UlvIQOjXFwxptyMb2N5dGtaks1uvd8S7qXcwTY2FMiOvuTjJ
m0QSkph1IPkb1/U+cZZNzNlsgVeP04CU1+qvL/Oob5fCthVRUP1uuDwvqa65
8WxUlnoWjFW4a2ML2MeU2bjWJbvCj3p/GcA+yc4nbC8URQki6vp2illDCwju
VJ3tQ+muOoOC/LSFVUDekyKWiJzdBxjFm9ZyC+IpoK3Rb1rJ3K9Rybr2oM+o
GzAjhgsRJXLnXbqyt4OQ01hPrxbze6Ef+eZA/cuSRUYeFlCsd9TPR2/06r4e
2dwap65Cf5EhnFw1Ez9zle0b+Bumpj3JMAnDHJZZGUPpj6sk8uKWKpdbdGP6
YwncNoJiNtRh155WVUYNgdPhvw6nA+42GaHfSKcZCCkHMjSVltXhzn1iuNki
wOt8FWh0pnUNtw4+G0gl755TcUZTfH0sf+1zad5tVAryPYdGt1K51UggDMSU
Ujsrf+DpJ3aR0eywPTfntymZwPCr9YDxvGCE4BfXKgszxRZN0jeuLAIVkthT
yFfE8swGT+WnyqFeEPF4m625TYKpflDXk4rlxBNGZ+BKpPKTXxiec7tBwL7t
ccrEomnG3+TCwynfUO/IQ8UEThhDx4GiAhLh8BCAwjzKtQbHE81o/9X+dpRK
MMMv81YJhA4JJo1AdfxlKNL12akio338Q7o3B1fPEok2hF6T6Hzr+rR1yEhB
JhN+Htz0Vux/3VM88iBZ7zAflvCRoIP2RapoKXAlcqpJOV8BfRewQWqnIzx6
4D2KiebpjgVFGyDL1aSa7xzcJbk0vwiN2l2sO2N9JLpkDhDJmxXOp3RKvWgF
5bQiuHoRXCyOmXsBUjQHXXNXm2K+DMUvoFMV02gH+fuFD0Lx4Sjt9qtsPZW+
RozhYkyUyRqFstrbRrhBXggVJhF7OZSSgdPhK+OM3V0ip1TQB53Dl53Se9ep
1LzcqacB3Vd9JE8EKfLTF/GXgCyaSBlu02/JNsFVnqaj6BNguczRRO9h5+Pb
UJJCdcEE9vCpIaIOKR2TuZG1GnqyNwsCYp6isx423h0TtnxnyqYpOCje6Mgw
vmkxv1ZfO7I1PZS5K83EjbNUvU6Z9cys0usDWoT28lNftlCvo0lZ39o2cyBH
ABiSHws7+K35c094tU79R1s0Y1ow9JUPIoFKOWvtOAYM7u6fa1sPfWaFC4za
BkdTz+iGyDEjrlAEWm2ece1aDOpSjVLsh6jU+1GvIJjWcB8IbKk3QxMKsvMV
Uid8QPOzn3MgPN+E3G4uI3dlIDF2tIMyEUAsn9CKHv2xRUrB2YTJ2VVk0Rj+
qDSdy1NyGBQL5XPtjhSVa3jljAjkRxz32C8j6coNMQT+W27S1eRcLWNHc+3B
i/ptmoKCiCWa61/AdBhZ0ely+Gv5ndyj2uggdkySAymUf5OYefmSxQ+9Gh6Z
M0HVLm1K8oIVUOO8egAYXTTcNqL54Zy5dWl+p3GzCn9lB+izucXLoA3pj8zd
tep4NXT4dXSg+dLRv1qr0aCLMlW02Fkjk3CMkfZJpWBkFgiOnG81xTjNYIXR
7s5NNyuPpAld9J76yrUNiGnaCEoVsKVd/Jnuo4+no1YKO2aXA+VBtPZneJeb
ogs7e5ljSFdvD8Z35XzxlFsYCmn4vMF8im9uQVCB5ta8RGDfy3+9HWnPHEaF
MUNJ0Tu9U2MOwgo02qa44Cf3p5RKysfC3JHaARaBpMMVAhT8NC4tPTKnJ0Pn
ZONLFH87erxQIrMO1HfPI9vmcJnBWvcxBul78jUVCFqhMqcbktoWl+g3DgFh
D1q3CrxEjuZlxQfN34m4crSrbsEwThhZZirnZrPWiHuQd9t9ImMphStS0BDb
4KFU5fiBVUYVoM5YKIoTI2XFn0v4HjWYjhpgkNN2TFNQ15oEnPzYLiK5xbek
NEsgi8j7dny5Cebw2gN/ARj6kUgpDTV/p6popj1Z1CZzSoltyQ66DVTqadoB
rn31HssmGVtkP6PjXsfPr8WrTsn8/jV+t7YFYVi0IyUv96Vpl+dFzzkec9lj
mEjAg3veXB0n7NXBFK2wBrWLAGr5fK9u5MD517RksCcRFJ0/ilL5/uW3Zt8L
1woJKCuub+Sl7g8Z3uXl2EhaI36OU2M2EwuRz7qbHGClnGRMcNBOnZB8E56h
Q3y9y5ox/mYqO5JQs67LrgSe2ldamZ9PgB31z67Dj0L1psfNMMl8sz2QAbGi
S98Mq7vr/24ja/6jtVZI3It5dunwYrZOqqWjdEy+zeiNM1Z7XZa81A2j/1m5
WfeZUksus+ps7ACCIkHJpiUn6QxHKyK1Yamoq14Xmp5ds2VvPLvxXOEo303N
xeA7g/M02GyB6tRo9iY1UNjXoO+jebvXLpWXhvx71nx5cF7LjcOkDWKHxFW0
pOoZJ/zoBGEqLId+mA+iB6Ar4OYmJS8a8JVVUinJ/8NQ4g1chQ/lhVMbjRYc
ZIPGggf7OHk+meeeHKWK2yGuFPN7Xd8qkCaNOvExjv3mrZouf77E2hfLa4tC
xbH+PbhsjvLHpAG4sCECZTVNYmqo799Qa/BYuFbk6aIREcE5vUFnGChnHo/+
5by/TSdno8SSgCtnDdxLg5YCgMMFfYSTGueSaZPgANLrJmm9nHLHavLL2UuP
MYVjaD+LWECoL5eHiTora4+8jmIEUXC5qGdyaM7W6QWrGGwN/bmUG3gqeJd9
LezG2FcTeiYSuQh/tO93a0IzDcILo0Me5e/mKVWn1BFu74tJ4bIh3Owcz/VQ
ViEE7hM4QjHrTF8s6g441GRnR6rgvdAK2Q8AXX88I79En0UQEinYHIXCqmKT
sP/TpV3m8jqajzrQTignwUXh6zarb330T1oBapOHG7PZ08IhaipA5BGHb/Lj
P2Xq3OBGjWsyvuKS734b9V8o7aR8+SfamQ3wOhPfznM9NigzVvn54Yhvb3gO
3AIr6cuUK1mVXyWfudVIU5Zy5f8FjaoJ38Iu3VH8sgDpFNuGGXB7AQaYgTJ6
Q8/0wbM3wzwOn9Cu+195hvQ1f0/e1Ao4m+7lgLi6ViwBc/fP726LPY40B3Od
mpCABabYDqcyWmL14lk52ZwBkIsqYOAj/iPdk57E6PAhW94p1Uh7Ra6ZrBsF
9kRRindFevCRUBichToTGxxVBqbj1pPONCK8KcL4JQxrtQykZ2ZzbkgC4PEo
TLDmG+Gu18rR+1b6UhtvmQ3l+f8EbKRjeq1Yw4pI6xmHiD/M/bsCOF3vrFK2
mQjLZzp5lCxSQWSivNMTG55gMqzBkM1xqisC75cY8kfw/xaQW0GSNc2ehCl7
ohq0QDuLCsN8s9D/oeszqOE9/nMPnu7YrYP2HIsnWQAK44V1ImkGta1RGW7O
tR6CMrAI51Qln1vbUBIlpK3d82w+vWvD5VQaFkbzqdAQVLDaevMSqTDkkNVO
xc/ZdZMyXS4lHMa9/Z8FoIQBbLEK48gAs5qd5G/L5SS0iqb2mzonnm6JuXqM
Pl3Sd+BjQODvd2T5WR344craUhy8/v05yVJ7LN0Re484ViYQvM7KHfl4gDxg
EfDu0hMkTPRKbarWlvP74SrETUBe3yYYnTipaMNKadp+iDqxbsl9BwPem3cC
g/1/psoUCz0fhQYvUNlG8PDDSuwg4QdbDFR6y68UD8kwdRoAZ9oiTjBDfn+y
AxSFgdTY1cE3PkbE2F2QybyWGJg3y4QA7ja1+3Gi/1IcPfoghBBgSVThb3Ar
7xBQcOmukXumtQJEeSCIqEo62XoFxW8/aD6T393+Kl6TNJ2/sN9x3bUj/BA9
rDV/phdqjcgLdRkf/3g57Du82McIiyugfbPqrIIbTTmIsaKLW0OeqxbYBXmZ
WmTLXrjcvhBs7Lm/wskTZplyfdZLuykSMsu2re5qN39kHS7P7rT/6zOzBeOZ
QLCLip0x4jiqElGGyPnroUtewxe1UX3PoCMOkRGvLchwsfLsvpusdr1nYN06
caefET3Gy69BYGNgX2GUTGbr6EaKkBmCy6V3/fWUwri6ZT5REw+do2mOPkU3
cAgWA15FXDL4ExzNtKbkZ/+YwhjW9ZdzCZYKzDoVJqeUth2+c/6NNHgJQvb/
NaFjpaGuzrtaLIiDRZA8go4kLB3vtnObOdeRHSHXJQYGP6cqAEnPQguhOGKd
tSXNBomQiF2dsdfHJcQ5GR0rMay9myTsbsRUiyAKvZhiQs8NZU/TnJeZN8cF
cgazEUDKmCaJZ1g+bxWk7IRbhka1rglpW3cqp8zeJsAabQuF1doeElbtZR1d
Q0RI0c+0RxF/Amr8hfp6b4l6eeOgqvbPCASij07I/bVAmdVkQhMrgvTbSkfg
65sMluMmeIPvSMnrZ+zkRzf/0MkvKR0+0o6MpDM8zpWSPhIqO17tutf3aEqg
jwhlLq7qy4SQgyj6/iJcviDrcYVO+5MjQyhyRSwbia9VxbsSypwlRXAN9/mi
v39IE+W3wtCB/yXqQk6Jv34NwZOoUd154yJCpvjLR1Bo2JdK/qHu5WokoNSO
26JwqquPR1itIp50YuZDVMbPn+DkW6YUzX8/g5E5Xrld49ZVcAiqrveHVDON
R19hJy8m4f9OQJrPYWGBRspG0/dQYk6Baw04vc+gHiSK8X4EdhmC+rjAZhc8
CM8DC9S1GHVoL6Isiok3gi4APq/ZylI8Vi116PWUdRCgS7oGyCRBrCg5MKPx
wmcwHD5kl/Ni42bam3t0sXFFzrTgW60T8KH9o+WtKFtOsrzrU+SzlDOOSRrx
+Wrws0VVCyxYLnWXR/uT+Q3vf8mDP/l122HKETkVj2Magf4ODrkwOnCINCn6
fz2x3F9Aonc+JUbtaOOR38lsSxwrBLsOYPnH8zl/c8B3XpTm35NHDLxn0l0y
MCBrz9XOtziyOu+uJyhjhIfZmi0zPcqV1gdeatqIMkaGjYZkRZ8FHM5K1VLe
ZbHbQn8mh7ToOlHZCMX9rh+FOljFIAM2MwrY6EA46uCS6uTB/rLJzIOw3W0O
2p1267aE5aO7DXGAy5aUIytGhIKxkFQ4x9LDNVdDVi6rKwVR8lr04TIctRb8
LGfKxwdRMV3VpqGzDUSfgifJP2cnfa1SDJNnH6A9+oZ/HS9O6wtP7jrQL7ID
K0FFlQOXJpDEBKPSvv6xZYaHIWWWSDXN7A3tiE5Ps5NDwsfj/w3qZjIjF9jk
vQlKkzCx3PRAuvANNsPdyfWROzOz0Jou78JnjVWnT7IZWrDm5A1CSUtUOfQP
23cJl3v4zGAmNneLe01cBSCHgwS0GrpXL4lPseckZvs0Zz4AtZFiV5elAuMN
3hb6MuIUXhNsgJbkb+KI5X9G9tnXq3ExBmYpKAy/LS6aNxVsHbQcjU+j8/pY
nHTsJX8njo1BHXG6WLomMUaSg3Cm2ldgtXo3PcsIpMVaOU8R47E8EOLuHi5o
ZaIHWdqPnGe8tqfU9EKy3RgD84PA7slit71DUl+FOuLLJZr7NqphDfKEGvmK
p1OClPDkuNDGCOFRIh2L7cAtfdFGj/PT+4CfLJsXGrZjZ43qrRBQNWEaHzaY
8jUSHtm3g3pQQC9mvPZ6YVc/CeSP3yLPjDkgzgf6Gg9ZNh5OXvP098HP5KFk
V1CYFtOOgUR8ajhKHYoKkRWrLbHCzR3RLDeRiyLjmkh2CmskwKR6dCa6HRiB
6lkbu4pPdpcpxbLPTDTh773f3zS8JbQEgazz2whcYn10GzPt0/5mdBhVjSmp
wQ8CrvaZ6FkLlnPVGamqKtLH5/3Of4Wa5M6+QRS6rlZb1/CWwVXeAesITipE
NYNwJwGo6vmGUvzxaapbHyGNrtTIiZBjBvCVhWtSMmirPuJLhixbH/VCmxzQ
cUem7nPq50z65o6bnomNAhMj3FV9niwqpleYDGRl9+tjRKihg83uKJOsxvFc
0a9HHxjrNG2RnPIEe8BUv44ix2UWLfgGCHGwPBGf2FV65eEftMD86qhwMi++
LqICBPejzqPnG2Y3pUfF39OZ5okm1x3t/uRSIcrnXyuaGk0NbCfBp+QqN3Mm
ENPPK88KFxRWt2cow1hdUVdXxvugqZe8WNxp5h5goWB8ezZAsB1VaiPW6i04
zGg/+xuKZoRwVp4QVyvv+SgOL6EkdvlcxzgLaIkTCpBgWFVr2PH2Cmxli94C
3EL9yqVwJ6y73f/BMrDJ64ol9O3hj1Iz91VP3dkC9sFeijO2pqY4S1NNRhn3
I1ofsq891uSq6U3o7w2/OYvlxRdMO5gqx4q1AnRYlF7XD/ApbVHeZbT53E2K
4ox50ZULzKD5hPBrqDsTrflcQBHPNptEUuwzSBWWKYKMXf1aF6OP3VMezzqe
m4DBCHaqzzMWxuV6THOXVkeZyet9DH+i1+fSwWC965W5CGSc2WWiG0spaHVf
UVkBjdo6BAARGtOoZU4522+TLC/duEI6IqfuIEDLYD4q3bpnArYptmGXlnon
xA84gGHC5bxqaDI6dxr9mdTcabe8B3QEHvH9gbcLSOoqqWHB8FpLDY7RvrYx
ee9X7BU+esEm7sjVfdd8GjDotGNLOpyR6o3dssD2PWEaX87pAfmeLhVyPY+a
7/wfot1tNykP20Ci7OYCR0p7m3B/9AMgH29qL+CFo8vK51fwLglAJbYuPkz6
HG9a6Rjjl+Wl80qlZpPmXhQxF33fFFpyMx/OUejZA0wjIHbzDpfsVZw2S4Wi
FLwnPV1qk1EZl4saLrnzycO1wiZRNRcmNnUlw56Rfsj1SiWhOp/Wi/XfVdpv
IKuQ421KgyLHsxDoHCBeugkKNheBHmQ86xWoOqVO8aUYNz3rxrPIvzYunMtW
Ydqx10nOhCx+Y2h6pY3mkGf7poBtk50EMsXxX4vRVsl1G02qYm+RA6u6kgWe
90UtB9OtsBHVOjwYkefe9V2YeAnwalBrH7ywBf+voiNlNv5rGJxuvAwnxY2c
X1qLuI90oSdbYM61h8FMm61sMTpw6fxfgkwBUWQkEB4NlW+IRIIWNRqta+pV
0FEo5tT2FapYyNYKtgasC5Pc8oZPTeNcnXI72o/AxefIy1/6D0vz6shJ64vp
UMcKi+uWZD9+vI8HNviWWKv93oIOXVBKhGAm1yGY3zkH8pw6F4+lZtEeyTRx
mkwmKUsbGHOuzPLydJmlgPJJ6S0ZjhIJC+EOpkw69r9ww+70DOO3/ZP8as1Z
80DoT532ld+bc3gJNLShCr8LNnbKzzjIL9gevI1XvwuZWElaqy799UVyxwT7
lGk+Q6J7bkpdNbgpqxyIeLdjylE7SnDVAvMot5tv8jLGGOniDGQKv6HuVTCf
9fRJ0JBgCZx1AcKjTj88PKYM7GLSC67K70dSbw4OGbpH2E/LnG5H31MUdsAZ
BV+x1rWHVo/Y9Y5MWn1EKuUzDyolhvQpNIOLzUWRLHlb4o8M3RC/BhKfkPMv
9nnl3uLWm9J4YOfTcNLwV2p8SgSPZYnqU1fPnV3RZQlAwd/g6ACa0DG3iukF
Tqda0TddLaR3Pfdu/gvfOUzpgqL85ZewFRz41wPK/x+Oy4oybEpG+j/Pm5D9
u8gZ98sWIrAJ7mjT4hW6x53qPuhLn4VyyjQyXsAyazFb8wqOlrBxnIBuRQf7
60dgarZGiYCHUjxmfPa/z85WrNwx1nyauy7AEOkfpKft9c995EIetiTvxIRH
0YBc+Ijkh9HMPasEe59CbcZGSQbZLxxPlRvj/ZEMC8a1ZgOs9PBb/BnCRbOm
akRVURHrJH0vRfkLDMVR9grri9rz9snHhnqQXJ8Vzeg/X1ercU20devAnLPW
+BFq9HNW4s2E73Khbg6XrEqKtBLbzOEWV/qe8P7tbNBClGZ6iWfXWYSvwLpW
CuWLCEuwrrFozl1h9KdRJc4JtdAoCFUCoEUkXpsnZFKagw7Jmrc401FBaZ4T
EKl0FnzxVTpD5HXH2fMvoQyrdGUPlWtHiUPs/g0D6LgHOD86QBu9QBmmATmZ
Kysg66UjIZj7H7TJVo7UiWFlq3tlqwnwyCM/aUhJCMMQ9P0fgAg67n6nc1hD
0J32pdHAIShjWLS3LCLwtR+WTjKEZfeFgu7XjbrMy1CJeL8OWDyYHCtVowSn
woiF7JHqq6j5dvv/J7GWK+a3dXz/YjiJSstLjOLsTbH30ulS3rlDQv0d/Vev
iZIAuDK6CaKBnqu+WOX5svTxDD7MUZ19ZX8am/1C3FVsnUGZognUF84/7GQ6
XjcRRwD1592QINdtsSqQUTV3hN0/yVpMwIRDoq0wuCQzs1mdzEPK8tfauQCL
fiO25qV9+o0CKG5hMagvC+Noa/Ugwa0ZMW6QNOwYwjlLnYiSnx4vMJUusk+A
8Gpm4gNCUDrZu7pnagJJyg4ENFRGh6RFGf0nWckkMose+SWKqjwYw6tTCq5v
K2Oyabxpr7W+kc3EPyb1WhVLl2t3qXr6LJ0Ir0on12o5TTcFv5xEFkq/VkSJ
4rH3P1qsbV0kbLCvpJ3otwztggD1NGH29inWM8My2l2MVKccGcGdNSxGUIei
AmvXWVdVVAnYt3s5RvfoVidQaV5++zOCa3EfPNlB+qZvkJ/o/DKdiegsvkHt
bznfBJkwkvPRHqXcVqMUeY+xtLW77GOQSmwJnwqeDC8XWFWt7dXl22F/jdi5
B1tb6W2TqLwCSkNis6kn/0XrVt9Gt3hvM/10qY5BSQ1SB+pQVJYyr6tWb7fN
HvFItsQxcMAi87GrIDffPRXPqu93QV9b4aDyJyYSURej2Mty+VbFX0oNV5KS
fqYKD8FTNHmyY2i6Uaxn53l5byvb4TDGdOEslcLQEcjjqHuMS4zBEdfACdps
LMbq5srDADkj+1WK+dQdiMcI81q4k7L71sGnlk1gN0IYw86qDXxQVJgWOwUi
BYSyOvKZSKsOeDeMQHO0mE61Tidu3q/RK40jC77fvx3ygbQt+AHRj1uMvT+Q
+gB2Xpg52iGS0tc5rX8JwOFwZW/dJd1yCLRO66Qqb5YfTiT3zC2C9pumwjsU
aMPLIonPGGf3xVO30uqJZYTnUU2KGo+RFgB2wTmikobuIvzI2qW5rsF243X7
7wgzddfqUoHkQnTIK51P3ef+kz3Mxej6xs80tQ/d0T6dBeJRfTzc/k4stlAd
Ldt14AuzzF2nGe5wndQZHaIYgGzha79vTZg0q27hG8KgxHO3Cwm2XnL1Cpo9
bGGO6jxJhV7DBS5PAiRV4JI0R/JrCdTEBXvwphrwuIflTaQSpc+mIQ+K/nWi
Qnprftk96YbvrIy+wJbFDTdqwU0lAqyTMLnIvT02/5vmvJBje4gCGIa3rRcp
FqSx0zaK6JnHI90kcwiaN1SNCXNieD7wVTuzXSCJcXkSOXDzybsFSvvbZcPf
2XYDy9uPHwsc1t7+ZGix0TvQxMKJGVW6EVvRx0RFeK18p6GQq4Hmt4I3mcD6
1om5rGza4xLdbq6RaBVNxsXWFHdyrhmliD99Gm7980uxiWKpMEeUMrMtFTCT
yl5tTYai7AnVENmnFjrkb2UpsJkdzpZ2mYNv1BiJS+gsY7tTWy/IKq34OmU5
CamzKAKxeszSfqTQmGn79ZxmSpKYdd78/XUytahfhvHJ/7xHuiXU/uBzS0YD
OVqha/pCHD4OOfkHt7KTAVJ3BmMqYkp36I0HOwN5wx/5CbDkodvtqLH1cPg5
hlf50rBwrl+EqnMfw0yqBRhLnbGS+93sjjxD1ElxXCNOECGVt+3Pn9CM0Xrk
kZ+WboPwaAh8M2yGSvcKCyR1pj+7R6kX+jsQchTzIsbsKyIrTBc/T06iEIdT
Pv1X+6836MSohlhfDhnn7VQDqGqb7Se/j7KiQk68ktkmISAlhX13bzRZMvnN
zjF/GEFKu6doaN0BDLVbXlfHEZUJeUx6Gds2ajrwANy9uZEvNn1NFQhY3pvF
ta2F1HEK4F1canRuzCHd9tg/PcVShDsoGlW2bkp+5cvbXTE2f2wjZO9PLruQ
9PNM5VC3KfFIpmxui9Bo7mrJm951QFnPvGrlOZBU32Du+FmeUEWDaty3/MeI
I2kZIOdIejjyb313alaJbcjIFe/b3559lnVwZbUIY3w/GC+BW5CqNQ9dnErG
y3hNPpI3Df9I28Un65iS14+ZQAGUe1BVar2gm6CYKIKw9DYawIG8622jU5VE
CbGoDRRAbbfeBM2Q1BujoT/B//F8Cg1xuY7LYSESzJfjY/yNruP8oZXFzZdk
zhjZ2je8QZGQ54lYlAawauugb6qJ5bnf+huz8eenTAQhGFj2nyinFeQR9jqT
jLA3O4PuKsSCZVdb8liT49qWXq7noSBeKFvQ48ZqpEfOEPubnbRzOpF0EhIc
XaXcTKp8L587sUjSKoDREtSAsyPn+DLk5C4zvm652PTrn8M2bTW8Eq+2BvKM
XM9IoyY9SsOkD6fUPP6pDgKRPhKHP8foo3SPmv47z8NgYm1YEA14/Gp4cvo6
FN6h9ZANnulmA7erQInc/LEFeIPuoZQvGXGhLpLC3dGMLrkuzvm+3dp7kK7d
VJnmyjHRZPjOLc0G6To+26oECzWm9gDHTruX+yoZMLtxGs0+EFlLnA66rrKG
6Hwj+V2T3LN42imvedzL5ax0KPm8xuUj/p4CIzPals8Wm9Hx0SDDp28eAGVV
D5mzmkNaWmXOxbr4krgDLBnUM3tj4jiER0aWWPKK6x7mwyo4fTy8MtYpBmjp
iUUPU133PmtNm6eXm9H4sTbd+JvD/payeZPgUe0AFRVv0SVMsybiJCDjf3tj
1WfUz4BktRdETbJ5nh6xhnuTxOYvnZkwQWgaxjUyHvKDjgxZe07cqTbm/yP7
z+h0SCwhizprWlvcHI/626vVFpFgOx2Abu7PmTj0sr+u3HQrNTANI4l9aLmR
NEt/+3itAI7BhS2596MNJMfD17sUqu0/ecbWEtbsSDamVheRMbWPIPfhNYfM
SGATGnZ8wll9gHC9yhz6XtZHrWy52z/eZ/TCTLW7qoQfLWnDhyxZe4yJweso
TyJHKkwMEymQO4ebJgqsm4tNxPcWOx+Ve+CxzI4fKSl9cIdw91BiatP2Z4jT
AEXjdE3yXMhOgVG7MEna0Q2tFTvUuqwRCOnwl4d4KdHM2Z9VTnh8+RmVsV8G
d6qpbI5SF0Mzwus40VuXM0x3p6g4PhWaCtApbRhGY0DZMLthcdbbQyNYrAjx
u7EI+vmUAVd1UrSs2YxowOxydobqQth4QUEXHHBdIPss4PS+PfCQkfbLHxbq
OtzQsWxFChKcIOuhGWhybmCNn+YtYtgKt72QPsGG0pkln/yVBfFG9+fYIJLB
v5+KzfhE3r+n7GaJzb9dySJFE7JMAYYHHi4msM/94riR7+p57cZaqySYEDz0
z9ZeYYi3RavYBZHH9TnYZ1wJy0aDMg29KB30GWJf8ZocK4Tsdi1/QWB+ID1h
eW/Nc0OiiogEmFfgBVAamJ/OzWn/QfwNUhV9fdEiLpLxa4SBBZYO5IaOcFp+
a9ssyyL/+Din74hN4IMvP+XDQ6/ItUIMbiT69KmX0SWPdZYR8qZz3Ukf5RFl
tJygj6sqHnDVx6evsSKyXiYOkMVSTFOzKdIEvM0UTMAV+4JUhw+b5SQ9Faa6
QwGCexOqFBfat6+D/CG6yb/wgEuQriBzOnp5BvSw5a2gUAA1+7s+RkKyfTGJ
pXzrtpYKqtnhaYxsZo7DKmASqo740dmwGVpjrihgIuxRIDZc16kjeg77US9a
FyplQnykfccy5OXo6ManVhVWlGvSWhjTzdIi0A/DvZVWw22C5F1wqOLgCkkc
UtqhntLlMDtuZwnjFvQa4IkuYPuNkkWWgLsySDOgp0QfZmZrnSFP5z6ZZgqS
aRfi/YeR7S8Cpd9e3aEwg9mdQixSv5VomMSFJno/5b3dZs8/AjQsa5Fi0S66
b+nnl3NH0Cy9rzseRtKWdlIXvJWql0kuku+q01Y8KHOHW9EB2jvYDNUyzBKF
8SkmbJcjZFhba906TnDNy6MEN9SWCMXLFEZEAw81Kwy0nO4pn74pEKLjbcFX
C82L614CohE2jEIo16GV0WVYLWtzYJm3K5QiaYa6Ma+gUCIJH0iZYXeOhUoO
tCc738km3fx5sgibHSU7NFMcXXNTyGE7JcsabMQUeEqP26FQO+ZfMhFZRHIL
QDFf5pu4wUbo0yQh2cW9eAK/wnkm2j0o0oWSusEOBhWI8J+NLwE2Uc/xUtQT
BSB5VY9ttb0UvNc9Ni9i1tS+1QrYrA24EHlI89pRKnW81H8CYjrRZxP9CTAl
LXBDJcPXjhif5QUyVRlypamW4ccncCioxt0DZ2pDtm9hMFoAj/pbLlqHHDlF
2pwIoiZckEts9L2kqqlIdpcIfqRbl2aWkxBaV0xekH5lx0N1DgHNn1Rlpks5
Uw7/sRWKPl15vybtHXgPK177uxylmRoMw5ifkuT91UvBk1/6U0kXQ07hyzdv
HwCNYyFZPpUFzc6fOI+T7E/rmn18zySmbSFIOjiic/0XVrsfAiqtXQxBRn6T
LMQindyHspAKJJn6qfcd+JbqigFSkIQ4Y6ZwEWn++Dse8uGKbCyx7YDan0O9
NpytfimrVkTI+wwiiEYSLS+dFpFQk9QB2eOCVEfTtPNnMTuS6nlpK/8hm0nB
OgCOLZ/WasOV/NSjjoNuSgkJyL3Di+DivrCpAFv/7e/g+YVC0cdi8X1LA2a2
0mbsQPOwLJHi4hYa/AtscHzFxbwz8YZXFe5+qkXNzz6oxIXOUhBpDEbz1N2w
QHMSarUBYPKZPpefBS/fLWGzKcmYslTSB6SxyxspF0zKoNoTIAeQ0LKsfCuB
VaElOKiESCvyBaQo8pfSPdeqO17sG9Yh4Uj9aT7Dbn+vcIzBuJR+IASMgT+r
sACi4QdM1BNnPQNa8AXHKzcTKnFU4HlBcjOfAS+YkGremcbkXsQI+3cYDRKQ
Q6FyGh9NA6lZazMFVPXnRW8gSPVobRSkjSaWHp8sf4Gq3O2fNoi0J/lC8mwc
710cTBHRwp6Xw8GIyNnx1rKykufuHs48MGfE9q6YX/r6cs57lHVVF2DRofLF
AFARUnCxHsNsIJfwWPkHMtI39gcIdGpF7xrZtF6bT2b5yVivG8EFFqNxeM4w
A0pG6qQbI9sluNpqrPHibOwiljnbARVwvad9ZCfs9kmhP3iZpS+odUhP4e2p
nHBlBZMLdz6F8AR64+ZbzUSwM3zCyLPChthOMuH2zZQBeFKq1fFQkHsH2G/T
8h3DR3zMuTLf/xiy59rMZe4cxC1D1m3zixbx/9OsGKsIC7HUrr4d/fSmjqJP
1DECapAoJiBpo9fVtCU7dIq5+lPQq6lrtz5WOd1Ja/iDQvk1vsoEoyPd9kik
4o2d2bc/gk5OAGrRq5rqtrXfwJcGbhN84SNDUKjGtXXc4ESrHjfQzp7XrWV/
9pRc1ydX3nkXYPvUP/z2ggiTJf42UKpJONcYGx17zDM6968nU3A8PmNl39FY
3pNrYMRzfCVPL9JiTzjqqq3nITPo5/Ij8hQfeLYFHC460Mf3zESw4UFTT5Gm
DOvl2hMxppRr9lsJ2DKfL8g6TPU73fpNa//NjDOrJC1H2SyrgJxlQkMyzath
KymkTqKlEKldgTW7FaYW9fOLjFGdEmWxSH5JSD0d71ei7g/Y0cuGWytU8aEg
0zNw1MhX8YGaPoD8itzy3hCzCnyZpxy89OCQ5r1tBNKHH1bAA2hv3dYzO5hh
sBA37EEiNLuLP9fZbZY8eMtz3fbhlriB4efOZVE4RAHUoE6Y8eTzpLWdWYKN
Nu88bl2RwizXoluFWS00a/Sn40lz5LDajZkWkgWWM3SWFRocEfw9stDKej7V
DC0VlgJh6nEbj8C8DQALpwTNOyOeW33Z3QPx+agszGdpnBIQ5lC5fU48wIsw
6ZL5XfMt+1H0n4BOrONIz3reDoxKwfjgcpSlry56owWWrp51zpCVbV/9ig4r
xqODCamxTn3f7OGiynA/N8RDsIYZlfefVLQNZ2+VjoSBQw3mmarFKSaftufg
wnL5k6D5eoDVlTtb3ATMAtTT9EINHQn8Nnly/h8ovARup/C84byfL8iErhCi
haci27EiClA2Swsjr+y63zqaSAX3BTWqiN1SUd3uprH8yDvtNPGXShdwnsoq
ekE1FiSPJxmsQSxWncs2ILY988t/DOmMx7YY3e0+cIqs0iLQa1nLgTtE7MOj
aMirDPaACcONdodvlGFW8ZIb2+aB39AUb4/UCO++OHV2/P+GcWl3ZmD0X06E
+942FFd8a/FRCtKlieK/roAhJDaR5NDTOh3U2OKIlsk75PKfMOr8YU4W/5N+
SeOv0iweCNQqUurUvF2T9dyORUQmz2u9VoxEWTeZVrNsURH8X8rq84+UhlgZ
qQtibcSHrlJAzTbpQZZwlpTqdu6cH3uisv9XVRzSAErFPgfHUNnIj1YoQLTf
yYzTLkWot1Ncg8hbfqIapgDFXjMpAkfrNZztHC5GxKSE53wxlMbexk1vsSRx
qLvF5E5vNhgj/N1NqyUxhO/YQQ86Rr14ibqg12X7w9xB8TXmQJOHW8AWfZ4z
WeG/sQUqfeb919dMpdjdJx/DiPDZ9cw6b2mWA2x/eD0GLHvxgTYLOH3vcMtT
VHarlzgMmtOeKkZE1RXBUMkAfo6jImueLLiDYlD5VDiJbJhu+6jWxshult/F
/VpYrNtoiGI+K9hZTB+t7Gfz/jMWIaYE2OGQnj3O2frThBJdz6dgWDSVNVQj
knjlpOnunOePjPd7SEgvNmp6CLR2uX4iN0km8yjhuG177ev6dCbECNDQLcna
ogr66VmqQp9S4X0vvSE//sE7f5C4cOfmR53dxcuTYQI15wXveGF8iPtZ+zJO
f9QF84QYXDjc68kM+t+IPzOWYT51834u2A8ZEdcQ1t0uej5GacEX6GZnyehq
wmxkDzufpvkPI52zS2vYcIOwRphSva3bz/eLN9WAlkkLvfXch2olB+QNvpeH
9VcfyENirgVZ6QvewikMk0XVACHVMx/cKO0gnGTxs+9ruveAJWrfi2dgrq4G
mrGwe+9rXBGdZm4CjqbQ5kJx3kHVruQHrz4QLpbJU1bWncu4h2kT6sdeT9DN
KKO5eKejO7EeKKbQeXQac7iJVAEw7ZHkAwN+biZbWa2pJ8FRA/rwPY1UoCYn
05JNiDeq/oemVpViFpfz4rZREF/n5VqOBJHB/hRC8XW3aQbwz6YXEll/Quaj
HuKcIe7ABdFtF2wNCT+yXj4YDRh1Lo6of9eMC2ZNsmdxffWe96DeS6potBI2
y9QtIBHW9AQq5Z5RD10xxlAFTtvJSDRConig27tSI3cL8N5Nqy+0vGbXMjw/
rZizfsilhq4//fQwkLpFl8EWJVZ6L+Ht7JB9ehUlaePvCdzSQGmxd8nCKuBq
dnCVr8DNsUhbrx3PdlYoiLjTKIf+9U3EjQAN+tMn6MBfHoRqdIayZlesayPm
Z8fzhQ6wIMMr4K+u2aaRH/rLbCtZIudQng/1zx67lmYzBGSFWcQWYG8Ej9/l
ofXOUguSrS0a2djb3xwc/NteScPUeFVeOmx7wpfpHhf4wndeg1AW4Nb2LhNZ
DqThwI06YNDRtSMnx7M4l1xHjJwUGRpThxrNwToJLXez7QymgFnQ5+Zk2Jps
qC4kMHhfj08zfHlBXYnA9fzV/ZMFLKJ1Y7FAKxHiazH13iWzCqbHWWmEbKTq
4vdsdPHrfuN0VGFWDzQ6CW9A11cuxwkXdtfi4HYQlnPuDI4AP3mnjIIyJhzZ
clz2xJ1U8SqScD+6aQmCpP73emN6zwLR6bnnV+PGusS4jPUmwYGHilukR9bx
E3jrYLHqd6opexHzulfN/TXkGgmLkY22o1v3tGSaPveMvUvITx6k+FDEjJtT
1jJYo8VzcvDA8a3oIlZicWIOIuhmXTQNRaeAK54PvbGdQlFQ//tR4nQTwC0h
mcgXG1ycQoCJon48lqCYY1HW7IFHhUxH4nRLG/uVChxWRr6x+ZAqxXVCReBB
qfiSgi8YCybSq5GMY3l3kFl3WVWul+r8+AuW3vk9iK9x/gOgEzUeGbE3ogP8
vLo0drN1CFDQS9mLZCLP4wCrgxHCyGpd8QgurAViBdH2kXhmavLtU8bzxjZw
5zsIahNoKhUwXljc2gjjzAOPR6SM1inkzb3QISziCA6JLhBoNjk8J4h5BT//
ysyw8+I5N7IGc+FZcHeOkJEdCIdTloJ4Yeg7ymjOS1IO7lgnfrIXT9UQYudB
MZZiY1W/dspH805VSKoBBieMNEZlGPE/Vm+sDw83WA3bvIg5DutfMRv/2umj
tIi/BQHN+GZAUTM0Cv4Zf25MW+0Vv1RQuNzKD84AuPY8rUcP8jd534yLqJ9K
FgF3Kw1X+4eoOS4OaqmmtmkZeCY1qXMZKxFWNqYlFlf0TuJOiWUBNyk/QfCK
8bu4vGbAtTnZt+EuzyozoF9aa5TB/D3u3KPQrB+JTD1MeqOATuOqCooZVRKB
aizwgxHItqpbzUfFHFMLCxy5HBevekGgdhi24xFvmnasD+4B6I7wQbj1hGHm
b8LCS/9KP5lYYh/+gmjJjGLasVW6Uim1JhH4FcVXpKRfD/pq7GX4V59p4OEK
iE+MxBHnx3yIOq8+lZbwqt0gNFj/2FKvJ9rkydyHZYX2/VmR1NwqZjdWzDpq
CFJ6fbntHABvIIrTJ3ay8AaRJkVN2QgtNiFhwqTmpetzKirWmLnTTIfws7RI
VIgvQPDLArUFHP/N7wNoWY8vgpNhv3wXCo6isBsnd4H8d8NpnwoE3tpP4Mof
hwrxPCNhmkSt7CZHFcVqf8VHjpHfbVKhUdBVTo17ZAel3VGsMv6v2FRMFAGy
uhpO/xQ70yA8H5+UpTfE2CHIPmKeDNdltLaaPbP+9ukfBPKOroDnTAWfAdoe
vkmeZiKWIEuyn0z3WiC9YnAbnLn4UeiEa2eifGx/rG4wNXgUM7A/FfhwVYB1
uTBYrSw7hAxyDX27miXxqM2kNEXmdspxASmin/cKJO2rS2lrhgMhvw72UM9z
5iRXKlxfwl6edXlZ+SoIzdy80D1lzpcv1ocgwsU7nqDkgBmARvR9KMoVu1iJ
9CQtzKxUnX02lgV6YhEtcZeZhgpYZtYwtqz1/T5R1plru5jVWabNwdesuG5E
jPZ2E3jIkueV4OU/iuAMKlDdJLo2xcsl0mbLPgFtHLiKNNhBMlH8MU3q5Vmv
5H+6pbsCdAq4ogMukn0BszpLKcosRek8cL6Hn8dBSR1vHn10n23QZ9hMwkHA
GPVsSVm26HRzfL0sdpZ64XmTGP2cfaLmP3rHp7+UFJKW6T9dJ2IbrTRTxLAF
M0D0yuAbY0LWi6oYc5l8YPR67F0B5bJtc2sfdgKK+S0G6PiQBKQEHf5Z9bOb
A1rEyWCMukH4DiZ7fe5vkP/1KycgqdygBOdfRcevrrB9yGT/Yfw7nS3u1wu0
RL1BfhZkbDbcIhzMc3DFgZ4Pfz0rSlklbtbBgtlUUwuTtIv8dzcSPBY5jnOR
Z3oexqnE+CgYi5onG7814FijACAtktg8xITCLcgj7ej5Dz4fjB01qPyveOQn
Dv5/XsZhukN+TvIoCv/YJi+Y0YWTpoGoA6Ita3iNcojMSBy5a8OoYkOzBpLa
fO01Q8/LIQ4NySaGxFluVAkZ7YX+3wpqH3FsnTpkT7z9VpD6E6czFaM1fEL9
nVnyYCuTUKOOviPHqp36FHljVwLpRz2rzp3ZLVnXEaPo8a076OXq3mz2qAt7
I0gcoF9PYXXGfND94ghxcOquwwsmK6wt3Z9A5QHOUPCjSC8zk5mVRQKCZgi9
UfMRgNj+X77NMgOH9VIRXhJLAFuPVPoyThmbcpXDzOFM2hdDLSl0oFQd4/Ok
U73uCr/0RTBs/B4S6TRfq8SHwUFVvmxiKAwGEnBkoK1VxwYUOgrEFhlcfsRZ
dLjiGZvnjBU0spraOHpWxN52YtlDGOiH0Ud2O7QPSC7hQFo3XesxZ8ViN1Y2
n2iVoIn6MmJM1zXtl4lIHn0SFuTU2ori+3Hw+ZWlRRS3Ro93Dq1+AZJh9Nsi
Cjl7crBXQm4IGvXFlLx6FZvA38YeI+Clh60EQ+QUcbb68zJAPHSFoh/u0ZRI
KIi117HrqoztYPohd/v7qbPq+3NPsOhikvYaeFVdQwLm84pCaUwbadl25Inh
OGmMqT8ho4/eqRZBwEFdkwwtW/H4we80AgHraGJDLSDM1XDqMn0xT/yZNex/
3wC/yWSCP/67DI4M4xBPE+g2U8B8PaNcvruGtMynTKsT+APrftsY8TBTET9h
e0pcH0SziEFbTdLaKj7JhVHSnpMUKZnDBjhQw8asxot3j5cFmWeWm12keqSY
M4DqUhspIjxhm+Ra9mPH3Vu/lhTtZZI4FDrOJ0S7bH5ggKdxp8YfL8s312Aw
9+DZto5clfvHFgSmbc0w3nTLiB2hxeCi9yvzowoOS43YePRwFGDEtJr8wuCA
h91plyTfSGHlR7iDp76DTz7nrk04XmuQN8vBkhQn8ABk2ug3fsWmbXmPNjWM
8KRicAPYbSjdnwmRBgf5yyER1n0bRrPrwnZbupfKhXh51lIvSa/GUBkUm8cq
bj87/63Yh6AVSwbXeqq47Lqc1m6ZKzmiZKrEoJvXPkQB9WOF1rFHVKoZJzXB
RKX4Gt6dkzmgY8krcvNOAR6Oha0wpMgWh2eZ2c05lM5KWr26NwSZCtmrCU0U
PLXhP+LZMav7P/9+OhX/z7BAr3CUiQol3cQ227YxyTIxcav7AB14v16RmEY0
TDuI/GnZ/qjIxB+bIUacs5D4SJd/9G/sPMuPdxyRQ3Aews/rreLcTjYhlaKF
d1TUPw79128xp5MRE7QOo1OhLLV+CVR+ilxfPPl2bGyvkhUAw/ldJRM45eJb
lQdfQUblyn9AasHDtz/4pUyplE4sgnE/LnE/yX9Px6yDJemaSGa2+FJxcbzT
vz7tSs3qvrH4L7clxyQoNkD2DHWTzyErnJKCM7h5YBL4XLPVm0SspWH2N7mY
JZjUb1skuLhGzOo16sjvhDfGqdrIo/YjfDQyO8i9CH/LHj8detE1HQafAl5t
sBRn/v4ddNstHznJwYqm/waI+Z/rS8o3MFpSWdstxWr7BkpvxCeluWv5pN+B
BfrklUK4+hQg2s5N59RQ1SEW8IticzYqybEIolRR34jodEy0Y9hgKQ0UhH5A
0pszGR6IWxTvVTfRGYN7jT1KF9189wfFP9tZNc3AvxMhiZgoNkN5dyUA/po2
toxGdyEZNRTQar0bwLq035Z6osG3PAm5c/cUjcp+HjKJmep/z0JvAFaHaA4z
ZwQy/vdl7zRMXD+P/Aj1E4Q98Pwi94XRqdS2dSd8yUpwETMJ20T5U+KTd7RQ
X0uP5Iph6AWY1RxRiuIpO+7aDtFJtYuGHh9yfatOBKTbsDKLE3kKVNsKWsIZ
a2gRubTWKPFRKav+jRbiZpqc0xrNbQdc6cOns2VeExQDOdSmJGQrf3du3Z0w
qPXqbRXIA4IUcakkOGvYW8RreeLjCPDvFJ6ChplM9L1J3AG7MaE3LEgD6Z3r
7hNhFO5EDY8bD6868LNtAHnRPROSMdyvZ2AdTl7kaQcnimjY6WWgN1J+NkpT
upQUsTgCmoPKM3uSk9ZaKCqnUPaG0/6Zz3/SG6MgXd9ZTNkf+hJKadvKKypP
5FuSwhg3KRjRESUM0Z+f0bbjkhD4LriexhXb3hd6oYBQEigD3GNExlWJBrZW
kjlLx2v4fZhPseswwqTBkLdo5obCl/ZNM7NUvR6Hfk1s0fXhRoPuEIqqOWya
6yK8n3Kpg7gVeVacNnf2T85zrOBDxYCOq3tIip/ZvtLNmwLgzv8BvA473GGD
bE0pwkQAtTK6qkjXTgCGz/iDlvjUNKO4T72ludwL8dlYYUqWLQesX76ME+rr
H1r2rt7gbDKH2zF8Ygmf17OIex8CrxHm39rM4kqbV9kY7RFr9snwyVBcVVUX
LmDkeXx85fUd73JKnzNtnAEBoCtl8VTqx2lqo83iLhmR6+SDQLVhqMejnHvc
w1zG202bVNIhqb7qHwjvJ+hgX2NaaMVZY4DhITZHUzDknEhikt3MAqBzKc4m
/P0gsfHXV18let175LUxQ72ZZ0Ci0fdvZ33nkBbrAt4xJcoJx+u7cdHn4uGL
RuApYs+sF2BRNG3U97gAN565MGtwblGCiuIZIM1NzImxCWV1uaBAxE03a/wo
9CBDb/bpJDY95sLLKiPFoP51KrnJk93jYAwN6WsvGZ9Z1Ge9xKXmR8sbu5Wr
eDUpoNSlCEA1wlfqCwFA0NDgid5mCxuEJvyzNxVmUPLh+mgaOeVstsFpTwNf
wTBb9IV5pqzt7v/Kr2zEzcbk7gERJCexOmkxG9Itvddxwr99LpZ+S1D6ZDkl
ILplQ9X2Jc5F950b4qrgYEXkYL28n0fg98Rb3+DryKKzA+p+NFXzGroKYZgE
32tkZEYbkItyBq/IXW1jqer3/JTxfSuDiij55iANbiQ56hCBFKC54H48Yl33
95ddGy2xNXh7IapactXQKsH0av/MDusALdeKdlj4yt72pW3ssu2SxlJ1ChnW
PN+UWdNkb8eIvcGgbGjG7d/K+mrBdTGsu4Ta+U+34jBJW1gigZT+NH4ZdSoZ
eFOajTrh229yD1ZsIRzbOozvokKrK51yjj0VhyatSnunUZNYPa/Rm8zne8I8
Ff2cjIz1omJQSozIFCB1R/dSTnmHgBRNHKTVsSj0zbaecVfxoKxW7eNRguju
giPRqAYJYUF6Fo5x5lIZxAzqlOrUa8uM9SpBmKtVk1G6GgZjbUQZSkzD6vAn
6goVvHujK2JHprRE/Q5IRNqrTuQKc7jfb5+Oj9XpRFw0iOpFPw66BSCYyw76
/gyC1Cg7B/h236KdP60y+BJnALLt5rZN3GFrCc4Wz6XWaIW+wq+dvvYqJ/h9
8IHwlIDvrzw00QwuGS0a+yiS8MWNcsFjnMv2nXdeVI2M4KH8r2JP4koUbR8N
os4lBiak3YLwvhWoZtod6Ydm9H2unE+pJAMp2tES+C4lUd0K3QrCcqX5sPKA
gfkkCCOe7TJbWaQcb8Wd+4URZkgkMaWFGMFGhlW81M/d2cefOcgNa/R6QxUv
Kg6/yg1hA2ZfSSPBti41Mp6F56gSIpChwAv2OHkuIWxpj6Ty3EDtw0g1ZmSQ
UFqqqH4fSyE51LY1aMIj2dGludEhDbi+fZkz1d2WszTt7XHM3QgamvcNnMKA
aWGRRKGbBkJVa8nonHwhOWu8JdPp8PAxJ+DhAHM78R/0zgKUlxZKwG6YCPZB
9aVXXlYD2LBT7CqkjHCmBYTu2nism7CAZeJciIRhOXPJKYyfTx8bcXWY8I73
jUopGdSvQtzNsOz2YkmcQCbYuaaqw0Is+y4Tqnu/e3zl7AfPrJCrUkCKx0Wb
YdsGf784WDyUu+EV6nHe9gv/q+GmMddueEQ99obAclGajprmEdfvSfHZFO5G
aEgEHEScqmtwv1I37lvgcz0Cbm/1r4kePhae6TcKQma7Gfy6Prw8VBuvjyfc
K0GTxgkyW7nsgvsxwNCVJKo1y5nn3Fytz2Xr8wDZY+090CfdEVBZlhsqscE2
59P5PjRIk5syMBYa8HZl2wX1nzJ+h0DnuOiWaI+Imri52PNszWoVjm743DNI
wVmk2BjOhruRqlQswdpvNvOeGyRuKYwOUx5vFZ3nRJPtZ2vyRdisAf2B6Gf1
c0GjdzJEuAaesVQf9a6I9JgMg723Tb7NKUChY1JWcOsnFLNTh5/i3zCuddsp
zUqGR1sOnK597fQ2DP4BP3CoOkC5D48Yif6/LCR51AUDzSOs7AQxDWExqY0M
WgiJYPdHvCinA4y0c636RYRsF9uT1GpZEDsSuM/bqIeA1tzg71OcT5uOeNvy
gvoziDlTVkqwyWmf2HA0q9Prwp+E0JDH3EjcKmLmS/d4ikPs9s9sLW3HubxV
QjNxKS9H0W/dz8bYTDpjSvI/x1SXv+9tE3RjPit0I6KXXnCP2Xf5Om0IDeWg
2N7Sc9pTBlVzIcmby8Ieu0g3aPY2BitESlWCz5lAMJthQCLcMr+B0xoOLjin
3hJn6koRcNl97PVWYxNjv7CFi4irEOSqWDR38nGZCBfy9boygaZQlKMZJTdq
8NIDcCHDJyf+BmUtRKM83/aho53I2eWA2I9+jzlQ/ya4KhNToQlIXZqWr833
8H00k+bNzk5w+LR3EQ6NQgZpVZYm/Bz1bHubaS5VA+FSD1iCA4/Y+rKilhV4
mHgPj+Km/5cfvHvDAsoEQFkqeOslR4GT3j7wQ7Y4icKT1m0fmpa9WrZbh4G1
Y1d8fRZJW8MKd7Z4v3oy5eiP8GSzrkx1c7sSz0qGXeg6t4NxP6e+C6RpYywp
GghhNwxsfVg7qpDczmjyYmh6ckG6YFQUTv8bunjyhZyrcOkgatTMG5z3HimA
f3YXJRkQH5gxFajCsBMwiK9E38jnscCBznx7uLEpFEuf3Nm5m7efcJ4vgGQz
Md02bLOcQz7pfQE7KVjfLxKsobqIPilE/a27/+7Gl8vabvNgq/mMz+D3MrWi
ezlbeRCH9W8y4Xg22oU6f7U65BmTmcofl447Ee+AORLfrH4e6GFtzjyUJQl0
Q4b7KY968IuIKAeAaHWL4Uk/T+uO/EHo/OrEn7KnpAVU3pe1tYOO7/6ZLRxM
q2H5a4gqcT1anoIhKubbvkVzlKGEGjtj/PqZZ7WumefIrU8Vc21ujjiDjviL
ymN7iC3MnKEIKW5jH0SJoWki9OO53lv2MB4sRtn6tNoEglfn0LwOE13pezuh
r91D73JHZnl7AVmPZ+f3Uoal45aBQhCjpXgF2I9btIDkpO3apojarXWdOwFy
fLn5Nk3m3TTOdaSaEcnA7+YuxGjLy/6KK4Pm9StuFhsuTrL4BVoD9fHq2+zO
Mmen7+vjtRUMk0EHLUKj95TpYges+kdtajXdQ0A4PZq95EpzBeq/jZWJJ1PB
/x0GuSetSv4X75FH3jreQ4jiMi4ILlD7t0Z8c+VQorr0sDxnMWj5NuXe6gkM
LAnlx1aZwh9zQ/n1IKPSrfgVlrVbnvkMaOMZBGUCPFpGgrldTlbr9zrzcTyU
NJTmPb/q5xDW0+iOL29BxpJIriEXDjYHcYVIkyrU6NIlWrGko5p6LGguWdtU
aMchDtzIHY945jWFqfNJ7WLgOKNY25zQg5gnvdsaOpirDJ59yDgwove6+TP5
JfTv1I9Y7YSubNUiJAlw0s2uEpNAx+zF4qrkl8+J+iuvXhnPX5rUTQ89f6K9
4O2tffWsyiQGfXblNXqUFF2igM+gQ7B4g7OTmdf9dyhRusWLFrvNuYBuFWXv
aljzVbbKS1qNurKRssISQcSaAiPFkr1SCiqH5TMLvLla+Jb7uzDd9tBU8ph2
ZmCOGLOnk4Ca95b9GWAadNyEXle9dWkBgt170uDuL3P8lqS6EURcDwgiQku3
00JuOBvsg+YDcP8uYqFE8fpFvX3uxOz6oOW9gs/3udZo+5ap1WTHmHoVJJ61
9aKt9vrfGLlc+PQ6TOO1Sxcc0o/mwg1q77w7LNO6rMK0dHia8PlpK+sCTpH4
YG/zXpp/eI7DjUyq35L/1Zs9XMUQ0LjHbPwgjnq2B3bTfCwZoGZ8ekobuDQ6
NbLq5qd4oq34paeHhWvylnUfXONwxTws58FCA1XwP0RUr3HPIfKlmiifsNdW
/woB9G1bYeHOeg+/77xYjOcfz9P3gpdQ1cjDa7L/CMRO5R33cuQ1RQc0LH0n
zxoS0CnaLRV7POOW7c+dRuyK1nhE41EFQ5SwGZaNdx6SEMPESRN0ObWw32Xw
Enz/6rmEWV/8bmmll1lzm/987ZK/vltq+rCWSIlXRWg3T+Lj3D1f9Eqi95r8
z3qIct6XtPVdHDf4fyePOwTgfp56GQ0H2q03+VuVt6LZkWeYgsk6EPcYQ5Hj
495rg3qY2vfoppSh0Mog6OWyOZwcVi/Gz+MftzmNmRoyGbls/rbTt12DUZAW
Oh72t59mDHBPzW71/mFvAIBY8egSvEQUkgupAScuYt+BasEEskXAtS0mkRVj
P4H7d0tT2v71adU3NyTTWWnoLGPpkvA017eSrTK3oA+fcjB5yAYwgtkiNER1
2YM5iKxI0DsG8+t5aZt1nKABD6FE9o0RAIMLe0xrVzIewfXf2MD/+v/CjnqA
mspvMVVGKzlhuupwnSelHaIM4F7+mF+ODng7CjxsL1VEox/BKmsVJTSZN01W
M+9oWXDYT9NiBDGPY+OJ2r07EDBXfYxzvXzPouJHD3eyFVXMochYotntwOst
IadyzSKlxBwcZDilKNEPk28oaZOb8lResbHdZVqcrRKo42ISf6nsdnMlkfaM
m7nJUi2ikrTwLMNNXR23OWHF3Ty8EEv/qe0OA2bi2B579DkyQ65m0wTXv0pQ
uRJ7E4ks0mY2uolhCZg9mQpOAHbjMqjO0qtjb4DEoLLSl0t24G2k8H/Ph75u
dTV4uOrrsQSHEcLGH7A9mU9OpCiXfIaMBZ7yW22LIsDtvHifV3jkeK0S6Ykj
1i1/Rs8GXJU1i+RZYGglI1Tsc0gbgQD4Fccm5kbPI5AI3iaqxIcirW1AeUEW
X7A0JPxiAJCsgd4ElkBvBTj9oBAEOuLnAhnZzqc3DXKoU35GPJQ8D2Tp9HWw
Xa31+yrlsaETBJL/62PoPLb82BUGw9sggxR0kdsHr5P86FTTiu+KGIeB1WVC
/PxD0NPH9EA0tiPXKBFLsTu9OGrd5+uGY9vOXel1I8vv3nlUIzKUWWjW0ujR
f3rLCctooy5IuQuAI2jFDo5vULw6e2Ex2k2S0N7W0kqa0t61njZwT6jjKgIp
0alzFGSUUQEYHM/96MS/Z/EBHvcZeSomkJFFFZHUbA0rT5MRpnIqJj4+SE0q
NAeAM0WH8Cb3jMF+MBUMRuE2HyZxBGU3lYjISzaxEd5uMvbuHpR3bkNDmluW
6P8Pj5/JoAE/5eWQcD1nv/bdh2CBzbPgI109cMNV+aSntQ/dW6OJJLK4i9YQ
L6GkNnD2h9FTkLXnTKvyXF/56ehcBPPZr9Itm0ayrnV81B4a4CJZB/zaPWp3
CVYHy4DhFpS6tdc/RcWR/btx987lzyq2jbwPSAOQ9fsJX47IcagpY1leEtjf
n04V9IpLyzXpuSDZ2B5o4bXavD/ufUYakfCabSNQT7Oa7zDFahqOKaCkKEZK
BaAVULEkltZrHh6sAtVcQNfuAZ2hVE8n/08cnahMkc6t7UpRoN9Bbj+hFhMP
7Xxes7ZmZ+3UDhhDjKH0UKNqy58bD33KtQ2Jafbo6ffzOaCqfWcLdQX1L/Z5
hIQlrsCYycBOJL60OEhVDtYfYMV+3Jjep3aJSwNFbkGdJSB0Tv04D23sCYwA
7WtnCmio0FVtLczkAze3NY95HuPl6Y0SfUmvx+YMsWLbPlec7tIc9Mg7sKoW
KGob8pp6LmG/KUKG9Yhrwci9QbHu9xw2gFICE6IdClDjUnrKoIhRrQXfSQzy
npJZQChrfqIbVHCsLsw4VRj6HkiS9DqsL0FNExwVg3cKzMHWuOKxnv7tPT+7
bDBTKiZlPZ0kiAogizJ+FwfTc21RAyot7NRCbpNJ5ANSwiolmZ7TO+PmQuyf
eAtMydAlGeW2FSUTOEwRMjGLsKtCCmbUbDOeWFmIPMHi+G8I3gknXsyJwcvj
tSkC8sdThuBFNUlsrxy119XngKKh3hBcnfAAxO9MAKy3ukkVLBtBzBJIJuu1
PrQ1j6cFj28fjF8EWxfs6epBMDbi/bD5aNLlOD/ZbuVabHh82DPHREaVcotn
kaM5+Z8tM5rUOCr30KTlNjZ7eHGt/4KOo10f1Gj9KQP8j6eNMXCJZK5K1Nwm
4OlHx9SnaptXfmdDvlLKRb+KoAFufnxgKWFVWm5XCi4liaPaBKRAI7NTp6Hq
vKz+NHmCxxz+b4SkIa3DEs1adnEI2aXGYccWpNIjDQMM2ymZ4Pc51//Tae00
W0eJek/N9v5iOapp3p6g7kqZgdKthkFPgzysfpQea+8n4eLPqPdJ5xqAK8VU
TJ15vYwgQopitahlO1Muf5gpXqm/1hOeR2+7Gl+f5nMvCjKnUUgxiQa/Vq0r
5rlsvlrc/t8hTG1D0XQhUD3sabCto+dx7PHoUFZpOXua/Pb0ZleRKHClOK6J
o9HHoEC5xnjMbX9+sWEABfu29IhoBXFHgN9P1X0v0qn8oyBPPNHRln0i0262
Q2wbibv86iG8PU5zR+Tt3dtvQQH4wnGhTH3BSVLtOpsTwiPALF7SOXypli6k
yVZwesLdTtWC3jvMMO4y35dxtN38jLp/I4N80R2Ze2ydoc4EmA/2xTWPbzmI
UVF1ZXNn1bCmOxeIQeTfBiPFy+Ks4YOR45ci1OFZMIIV+40fKQUgimMZlm47
AH7H5s1ELVqm1DnI7dIQbaFPwwSFu/RTki4PQeUtWrEhWQ0173q912cf5s5m
GMznOEvC9xKWoL3rhFIq8XkUXq4eVhI3lvQ4Z3BYmCUe9PNMxM9CUczRwf65
2VKrGo3lq1+vfY4nb9KUjfJ89TDpNkLVz11E44Ujw6zBNqAVwqebbCkCuzUb
X10am5V0jFRJSxYiKhJ1lSkbXdjmuQNm2zpCDdnc9e0eiJ4AuTvCwqXQXqux
sMm29Rgkf33bajpaYwUW773YC06oUx7McQNLh8+ZdyRDyhwn1Z1N39Iai3Yy
csBu9FS7kh5NnyrMb2C4qYZ49o9MqviJMpMyyyi46owZsjIbqOl6H7UFaw9f
gVc8eilCV1tYe+SlRHVf359RAbw2uqjAJIoTz8KRDNEoW1Sil4yiUEYBJTB0
QYEbYTcJR9GZnYFlZ5MpYuE9GAb7BkBuefwUgxpVv0OByPw1NgAAGKy2I/7a
iLB/zSvBf9cc2bXFA4And1CAMUT9s81yzG4X6NPm8gvEzKDeJi4gG6lZ4mwL
DPMJT6WgXSyF9C2Hw9caK8/QtfkUBEiNDoRZyWmPn0ijKzs1XaXALWC1R+Z7
Eqm9KoIKjFqsPFknES73h8Ns9WIxnWmuOkf3bVFyDMlQWM/B6ZWSpOW4KgrC
3jAvGEwkrX4WMZB6E8CLCNxoMwmorycgozJi3rUMNGpvO85EkCiYFGIhV7EF
KWBHPfd8SGcgrNT3dY09EH8PQy1JBCDRkoneL09rMTc4FVZZqcPiStX/6Muz
wD4VdVCeKsPK4IehmZoNf4UqEv4clF9rSBMoUdRJSFL0iL+rBcNDdygQ20/q
kUQ1yBDRLbU50UAkdjhVh29yEKASkXuoTqbneOp9cwitNu6IYRKXAXu//3y6
79aMnsbLacL5MzCpXbSFYRy+UtYsZkKaSLLeSyjRm1V+l5S0C33d41vFXmFR
40NtJPbNaWvFooRtYLkor6BLMgfQP4+zEGiRe0xKRAfrpNpJZC9k1tVj78ML
zpMWQM6Xq8kb0KtwfPOhJAasjEyMc0YAmeHanAB9A5mPEQtjsrl1p2ElpkwE
PYCVAXiSDEHagE9XiEsaVvwijAnWxCRBu2U0upD8QEZmJLmJPjh0HwnwSkX+
hqx4CdNmPLzbxponIaTbLU2Qw4k+OZ266bhdJa+bSKM2inARF6Ifj3mhJAOJ
sTQ5d5bolvzznn+W+2eV9LXgyDbsZR6rZcb/YapjYaXF+H8F0md/cDTGtzyu
+KWtAbNX4jkITw6kQQu7/hqo8vXSb6RObzfrQ/2sxZ5ymT/ZlLeOkn0l+57D
lR+p2oE7sNde6nAjlVsVkskKG7W8lvn6wQpBB8OcT7wIdb3z+etsvAwnt5lh
gLaHFA6yiKKktF8tMOBerKlt2tTBI755uLaHYguVzUzwBDc/vWRhuSA0IlCZ
0y31Z6ZGDLjCq0mHK+BNxmIb9+iiiQ1Hp5czSRVXyxx4XltXV6Y3t+30TRho
D7dhSWY4ZxTTVNyPznNcknXBxWp8TBMuoXNjqG6RCLeg/Y1LGqEfntnn3JfF
1FKik4iaghLG1Hx/N0WClfiLqpRqi6LP2qoiaGGSGHuno7XNEc/oScNeiykc
ZyEpSdhA89Zyxfn+fzmmEOxqwG42iQ3a1dr4vgsXtJQs6x0vZUGV1bjcSbUZ
ZcWzRkMZ5cQsaVsLJLnFXNk2QHlAo/BIrh21JZAUyqWWU95u5ZE6JulPHB/8
vMpowSsKBb+2Es7o4+6IiXjRSNQIFggP8WuyVD07OWy7eqJx6OAvWxZ0RS2Q
dTZuhhdOJxXMfWICt9gxMhz/C3EcLi8pqhll4njlvSed5fWVFR5t31NCrb04
+qei0+o/EB9nk8IN/J4Fm4zxWckQ5QimLNVjQGBIxHd+R4JQ48ovAiV3XkJp
+FppdbpQu+Y8llq+G/Ab0ulQvpx3DQ39Ag9E1m/nyXnx9DW7o9DHMuYMXPtg
nB1CEdU0Ihw8QjlQf5ehGJikFuRdk5nCsYY5Nk4oIN8OSQzkoZu5zpducZXI
jw4q4JaUCIdohtV9+dtJWu+qTV4ZFrLlaIsyrFrCPZQtwD5KjBlparCKoCxP
/xXNGdzCRwOYxMRLeyPsiS0cSgz9yJxmn/HlCxknIMn1W6Kt5pfGzayQOg9/
i1DZXnRfpj+uM9lEr1w4PAwVGxRgaUT6t9NJB/kVWtgvoW775LAId51cn+Ks
p2FoL6kcuacdPCkW4wyo4PssmDJg8fMaqur1XEkeCESCw1efY0g0RcqnI/XH
kXLmFr2iOBlpdvcIIuez1v/AD1GLl0l130ht7dJvH2eXj527y8SD+yHfpgpw
iJJtP+mj3fUOrZTZCRewprQommGPpHcZ9ksKe4nU6YupDvbTm73woHzgsLBN
IIf69MKLDMr1jJiR3MAbtVeq4YQXBPfU6eG7OsyvoOEWoWxuhjQjIOfq50dj
/7qSpSrNvVs7TIvEBrLxqb3OaCBmTV2A3PJi603v+ieNMniuWweQ0h42/JtW
PKq0vhYZmJARNxv6sLgmRXm6Q5mz3+roghnmbldfO67GbT8lXQYDIZN0o4Wh
2mYKQPsvdzb6Rp+aUU+wPYHxvCAqrLnLQDt4ZEuzAXRepYxC6CI7RdYsAaBS
BhnLA+zprsIo/4Wme6oBnZMhtFThtzmeZIB5MappgzE0mRC/uxZ0TnNwMBO7
J99hxXeDISMlemrBfqzy3ZcxX9xr7IAqIi0UA+BW5yoEaw1eO/702jTLDR6Q
6RnEtEVh6qVmMHlcY5mszYsfj8N8v5mKT25AApRNw6DGBqdurt1ATuxG9rNa
aqmTy7/EBgfsH7rm/MTHWG8cZK8Py98VTeYZ0saYIZ8sH9f6yf2XXz/AFECz
8ckH5OtU0IEoMyC0DpP/6MjK2HohBPyfQi6DiqwD0bDyi2Xk51WlT9qljMBr
xFz6Ghx4cTpFfKza5auEQ5DNajoU0r1ptzmrM1xgKs7xEbVZHNt1r95jonq2
afTaEPRPUHnwrRUbuH4a9BV5UyTNFJu1Q0RrhLy1BUVzmbsgbZUYPiZybAPw
ojMPUYW6Ss01CwOC7A/Muh72/YWG2JyNdx/Q8GDN6lKiFGkmkkMDi6M57cLm
tjUmbPm8TjzNF96ZwPa1+8mX7VZMJioYOXRQ8V/fCslCPgX4kQDgd2564TOc
McqJ9IAP/U6Ud8X86ibcg+Imzfz1yS/5lG2cEGbffY1YNeiKjVWUxOdbgaIT
FNUYEaMxQ6ERpuu6YJGtvIzBEeHnrE9rtQjBCnR1uul+Bcw1Lzu3qUzEcSt5
JfXHm9YgnxUB+61Pp9809i4pOwlPcgd+Ihl8W/NOuLrZfnre/0kNOIU1J7XG
ejJI5BPPctD9c85oZ/ki7TtdigFo3ulJ/cJFJoUflyle1c5Me0i0LOoyxVol
ETt9c9oyFRdWuxu+3Z/9GTUZczm/xBsjYBwxJyeKS1bVJ5MTZmQ8UHMw2F3f
TjpB7c9kGlBYLKFsa2VUkKUfAKwzU5lCBtOaLjFitX70lKy/PGYV4dlcaXVy
K9oag/hOQSDYceA+HAiK5LSOIl5T7BFfwsFZ/sVp2Osn14YF6gT/bOs2MHaV
yZComTcAZ9g18HFJJmkuo0D0TbYXvcnwiMSAJwkxjHPrABZtTXMyWkekyJ/T
yTRmA6HSmGHRwDb0l2/CewlGc1IAEbNS9DxLMWDe5Xk056bnFFzd/Uh1oRcK
SNdjvb6Q+/HCfRE1HMYsDzFqaExVHyKO0qK9QXUCqpEu5RPqtrYa1gxjtoaR
fklOYvKvIDmS8MOl3QZgFsXwNYyLKqQjmt9yLgAMn5DMG+rPp2m/hATA5alg
ATezPniMGBlXYBAZWBd3f69KvyxRZheB19sOa+OaKP2qNxVMkHnidZwwi+V8
TCpDguTAKIOvyJhdYKG/XfWXEy4fTJ7TeT8HVtrgDBgWQ9DOaG2moKOb9YXe
V674YtX3S8TSJQ3kwrfpE9I9j1C+JO/rhNLhOz5SJGQYbtEJ2uGD6f27PFoF
quTstHTR7jKm2FTvstjyPEvqdrRUbEdVbQpI9Y/o9IeCo1FFumdd6VDzeZY7
O777KtMYjb9X7BCTdVr9FwWNNARfyqOx5PMaIXicGx2K1FPug13u8Kbd3qvL
p0tXzwTStCLL5pBeZ6zfPYvjpKhblb29EyT+x0whhlBoTV4J4s7O3nLHW/p9
PNggNlGIPdq/6XjKgxK62C+0lpRGeeNPQOXR2b0uysqT0qr71m+FdKTcRi9S
+n7QcZxcFCNCJbekWAWLsEy2mXaUMzVjv4+vvxNiiO9KlDVuUuDwRUQPa9uB
o8sXKvn+pIGLaH9jpOa8PPH4BcpGG5Dis1PVjjgqXBf74IRP+Lu8+DEpjIVp
sxfJI8xNO6yAlue2iwFY3rh7bdDSskRh7j4s8kuHUc/qt716W1VUHxq5AiQu
rCgVGmlooWVKmvKAZV7LTyRaXSoSGZo3f35s4WUrHFVpLFIvuBy0O/M960rn
qXXkEuLybUBRiO2E48Gg1AMFlgt97NCjpbAGW2uZg+J64g2VlP94oHtI1m1z
cPM2gmNSOc9oTOfq9yW1TtYi5RZaVtvz/v7Rnuov9+TL9pWUSK2p9h/pektG
y8C6Qy8i/hdOFXek8xOlgCf91AtQ80XKlNWIjfJHAUQ67OcK1PPgsTWlKraV
b8KyOtwulCwcFHRPSH+arH0nOgKZ7W8J3pKEeMi2tXV1z6BDS0KGMMhngqet
ED/7C6Fwy3+XLCkIQTk51/LRocoPTkTPvL/0PcIoYhSGWo/RaI5Co00FVdct
n0WbvMi97NztEf76doSFb0pcJ0nng3r2mfQijIv1s9R4dsWWrDq+rjW5koMN
mmUiBrKquBBxH74gmUdGyqK9u8Q/+kHojyCSBoShFiN/K4atOyivPo2Wfkn3
6KTiHXusn6NCsyNpEaP86HeBb5AnzVWgzJT44DoOtPMwbrwbttzKx+CyHTC5
5dzNEX2Yrrkcc3heYGQqr/OgO7+H7SlUdI1UmruGqYg5JpOJFCwcE4aTRB3B
sueh6XRI0BWGvv4nqwkID0GjcQr9nD9j9K/23U5Fz+kdHWdIJyOuzoZJUKlN
obB7FEbh+28rIesU9PXUEL6vQc4EoSmgQtprUK3JvO1lb5RiCgVz7aaTR5OG
Lpiue75SqoojNDPL/KoVaXCgFnIhMUc8bixgi4M0F305flO4cpyKStRF8B+o
L4vbPJK419twop1VnCVXpLC78yUgW9OcY8WlWKbDURAQzAaTyhmhptAXT2xR
1vuNqETLtJDlsIpjyX35XDibQm8Y6hCm6VprkRpAmdePoNAP3aMjQuhhykLD
hu97rb9ELTEqo7dnUmJw/ymWrhvqTf2G9kWWTEBu/hHSqPYUrwA/NVvc03A5
m+waIW3as6W5bbiophHSEM3KD0NCFa9gsggtIDszA+l14ornlhZCXaDcEx2L
KVVM2mFmE6tWGGgUhsW3pk+B+BWkGQVWtoD5+Iwk0daHPqg+rPcHoro/hMnX
4+gJLehJ+bi9ZjnlM7QCkq5eUpMdu2AHLoAS00RpLs0gm+zQaRRiAvSzXCNm
BLLFPm7xPDkTWoNVHEpeMFL4loovbxH4nSnkfw9gv2DPoD6TlH6lMz/C0Oh9
x4qdIS4EStF9e0cCD+PuvrmS8BcAaMgetvOXFiZB1Hox94IixzcgDExGh+2a
bQ2BbXMFAD2gDNB5w9RG6BrP44qhDI/oPq881tqRtD2qIMnbDhCnaoh1WGmW
y2FCEYQtKTSlQLCl/dm34eMUO5qJ/sH7mJGIXx10Rdq1UGLM5R7HtmqWYkeY
yHmZRQpjPY6W4AFDmX49FsS2NuYSzFFHcd1b7bnaW7m/0XYTKjYmM1Fs591j
dXcy9YjR7bKhr9NUWDNFxAQVMcTFg4YmzbA7Yw4S33gJ8woBl+ca60Jo7fDL
dkzkZySdyoVLwglhFIrszPmdjSWPdfUpyDFOjwYzV+dOyqm/wSMopGKJSF/I
t4yQHRNfzFYwXaab/rX2nhuJp8SAOBgTI6hT94aaiaq0AimGtsu5vmYcohQz
sbtcWsBof2+bPC87AFG0hdLpKaJ4itbFA/vsYPk5KOD1KXESqiUC3KgJJwuP
988UCruyEYPoCymU/YtSvhYXNWfe9hwRWC2Hi3jDO8Tqe2gsrc8EKkX+rJ1+
j27Tmn9koSHRgN1oM4wHEdh2vWkTJ4X06N/6qv+bb9vXaVzjaRxyeJVD1VV8
L08sjUYUPu9YcbMYe5abWj13aKPQrNYvnPs1+MNF+ohJEVOls92P1hP9Qltl
yw6+awSBtoxeXZ4tguLV8ElRTQ/NpNc+EmT0EiCkv/RI9MyQGwr56X+vwKyS
fnJlK3Y7XKtaDOFkBHCYflo7pa7VYUFpn41hIeEim9VT6ylSMXU1XfFyuJg9
1WpTqcYUivGZZQzpXXd1ZAm3ITLSPsyjHz/htPVPowXVWH4lpDtqgCs+NLt2
VnrjUbAVhdTynvVOQmAOcwcmin2iwcJnPab+Y8dcBu68yzQzcawF9igy5De9
YJx5JBybGHk7yzJPhdppIBfb7viqWRyBE41kk0QET8/H+gOdY5uzVZPAY0t9
OsKrzUf12+K3ToAryr1xn1afXpC5pT14hNRGOFpWzNuED5jVS3j5jJHPWJl+
g8yX7D2SMzdeHK4+FITgcjEBq0Ym4JJjncXaI2aTmF9N2SXEF87DueeujTgs
8Jex5eti3ZRZSGAlwkoUOjn9truIxUn3iG2kn+WSccOYgwFNUjxJ+itA83S9
i5QX1RM14FFBxICIH36UELgYEtwmLWx8TvkclXQFRi2CnLwRcQG60JBXKYQo
/DWNYS8JvbUi+4h0J42TunZMQDGCzd3jQ9P/qL1MfPDiGkSWyPZBqiGaLsL9
IHvg1/+B7UTMHsXgO4gBoMmbj8l7cKrWVFF+a5fOKVh+OVeE+xZHS77YuuWV
UZkhifJmDVzVu8VxltgJlibs5r72AUFqPEqUV591/HQ+Bzd0xKHe2sfF67TX
dMi+t//nlTxr7vK/F2TkUzHJcax1Zwij4lRQMG/2664vJKijMyogC4nkkQBC
+0hMe7u1IU8KapB7l2BGLINq2qefv6wlisx4mZ9z1jM/fCcYk2YK+MaxK5yO
KTNPg7w2NeSxjsQr9ee7iR719Qd2mrwh/OtnOXYfpC21tsoxI6eAmnxVVbDc
uGBNNAhtPyLfvGl3hHhhawQoVq9/yn/mNFiww2yz+dErKcnjYEGizjjiyyek
H1xXF1AfxiwITD3Io3O3xWumbPojhCHMHqkfi6Ud4HCxdqZzp/sxk/z8ju1/
LoHxybRTFPfhc87dDOccYFQgBUZ049Ln6iASId6hJ3CtOtZR1rqroNsvrzd2
ulH9zEH1nGKLdXdVD5JpVPFzSshjuH1jsNGQccqEy9Uhh8cZAZ5FIsVd2uKh
8VhD6CTfcafix+3fK2wqMgEOrb0aoPrToZnyunug8qa5aM1XSPyVPi9yfRpO
xyBfNVaK8eHfQzSK19CtTdR1bUZVh1ntrtiUgDtX1YetJfRxI4iucp4mgDLh
O83fLEA8QVRqFcYrcj2Qg+5y2xivdWoCXAraZwOdkZFqahHR15vGfudjN+kG
oBogi8JPS6EwyTv/vapo58Zr7XLdHGZV8hCZn98xi4DPqp6RFUssYJCAlkq8
ubDlAwocls/Bsz4SlYAM6U2IvyF5kfLcBuk3bTkdTfUENY10DQK4JQySvyI3
kXtf6XXdoargePvYWgSAS0hPXMy5buILIDkUxfsQnUnrixfo3rMI5XdDlm3k
WMqPfXyOInRwxT404URoXxsuVPIlU+ocwsqbHfahfQ34cXFPKthFK9L3R3t/
emIhCViN5RZjuvrqJKlnUAl1DYCDV3hfLGZRlgGQAUPKqzeK5ncitVaQ7r33
P5heXHMDxig42Ti+s8BaBsPr3xk02R2KT6d5+xwD80UgLX0AbdhyFyxjk7tJ
XtRj4xBJwSPCwFWLbM/DtOYQCvCNke0FvVtloDSyWOlnK6BG8cETA5vIC/vX
RpSyi3arjx6wQKbZJ3aafgSShrzevVFQRaZjFBOK+HH3kXw5WtVZi1FIYWGT
0iN8RNIMXF4AF5cjrZcakhunFgfB32+3LfEbHowEGmSo/CMCwfe7wPh7WCtN
dY+PhD6YSstYImc/6NBaVsrgUfFkx3Wi9ceuSS/faSSv4w52qbEKS2tbKP0N
AWHGChGaGVeZrxW3B1KkFZCw1T5YOzsLu/lR8lVZqx+okZxtEPiXeeVM0sZv
hzGPRFL2pK3Cmh8YguNj8W+2+4lN05+fY5OMbcYOZWeVvwd271IQVQUMAugG
afupdtY8n7wVfS6IP3y7YwB7gX5XS00nHKKv/CvPvz1601W4O6RqMPBXY0WG
WUhMcYDF0AVkXoqGBpWEAcRKmPU4+gke4Z+Un8CuVcSXICmLfJKtvaGm9vdi
7I+9qGKNTUf7IY0QSQGxm/fUIWFf/wFUG0YqqK4Em5/ozIAuc93vW9n2wDml
EDyCImW6Va65hn0XXtXDyE+QrXEnQD7egdUsGDLi+/WvsKw3IAl6MwaCDpE4
1USxwIsR+oIe9k/EX4YhLaDuI/DwLEgNL2LJFCfbTGCthjJBSokpDrz9lDVg
VHLl4ZZblAjPUT4frPbpuiRhJl7ZLgLpN++lfxrx3G2prFmXkB4OGw2B6JNV
AQu3OxwL4jYiNBdtYtxZynoYHdZXZ31yZwSuo8fdjHvCP76Q2yWYE0l/qMQG
CZ3Xtrf2iY9S2BKYEZFgOD3PlYO68A2B0zXOXy4WveiGWpEpq1M38iGz4A3Y
PSuRXcVsqVQopPVv7g+VtBgNZplMTvn39n7sLtSp6GqgStNsXENAJoNlH6gw
3zK0pFFUFOTzRVPRio2n5F2uT7X7My1Y66390cYHahs2Y9SnMsFR7FkX9DLs
p87NoI/y5YecXZvo5m3BFlIIVft0JuulcTln7KPOKdHLlroG76UCl6Pa5C8n
WtZZyZ+0D5RUrrSKXdwYuGX/OuCIoa+aTTn/4crM3EYZr59mdSj8p+5zaZn9
mwTgnq+17Nsw/jR38hgFFexLbbsjzkPOJPZr6v4dv2ZuXyDUXttEI0g38fJe
KieArPTuVIE8mIEiJRCQ1yBLPBe+ahtZFXfHPaplDMmipMXXZi10GTrNvg6y
kU0Ii8MfkV2lBPyuk+ixXhpHslSsmn4vd/aORSNHnpbJYgb3R8YNcdySq5x8
Lm++5w6UGC89nPqCBZZVoUdcL+CwiHhQ3DL0hDr0Toj/mJSHW1uMKISv2vUi
wLak9f+3aTmius0n6bxQYOZHHwk/oQ3Hv25dFvnKZ2UieH94jxxv1HTCmq24
gjxbtN79Vj2cOdcaRJ56P0YVrXTAt+tg9AcxAKtJyBasu5J6y54tT2vNXDVg
BYlBJ/eHuDUhHFk2V+obSzT1tRZW8tkTVJErSWUiZasf5bL0wuIivz/dByaM
50Rvu+3pj1TMVP9g15N9BptmB8qVHrZgT42pbqqWskkCEM6s3y/ZwLYgcCg2
h04G73/MiaDV30idSranJ64RtXiPAv4QMrunn/l+UjWXh5gOlOkwPbgADbUQ
oESpPuo2qTvAuoRYpCQKggabcBOstd2kc7U4S9SG0xtuN8NUk2Nw4e/fPwNj
BdMmeIRyp+n9vVgqyk5mjNsw8CyAEz/96kffaBNngXJOxLM9zwFWi9MXB2v6
xFe11wgvRzCWU54HqdW/HD/8SPklk5PJcqnnDral9VRVn+w+sXaYso4jt6w/
8qk8ohC4sjKYcnpX0+/Hr9FVGf9Al8F49M638DwC43Ml5fhdlMZGtuzWM8Et
0YuMfVkJmr6xCAHHiuh0cCvitycIaOKrRDkvU4hB0vj721KUyPubGEdtiRom
+NFcb6Td/99s+ZahpWWymrDp+rpc+ri4XX07pTpdoHC/n2kGOKxBvasf5dOH
omtEjYI1CIiHzwwoXnHKhwAdwz4TSV8us9dbPf6/Oag5f+vcXbEvzrCjztTY
N5ug+pFSzP1Hw0MXj9BDhvruPVtyZQ/smNsaCgvUwbDLIY+CEcV/Je2CmWgm
6/1IVKer5mpclfkWDofDEe0P+QD2bkLijHzP4ZwHHBBGcSUbcfsU8h+WqQE3
Jkl0F6mmbQmroeqIYXP1whXKj+vrQjvLVG54gWWbTVOIug/KpXAlpVlp1AKF
atmmfbb1ybBTi1RZQUCV9witlJChmUumUUgPRtpCZaY4cSB9ZXD3caTEEujY
kIcpcgKNv+LoI21opCssG9DerDcc5XjbVTn2tDtCh4qwZbmFqYii1SVOAfWa
UfVG2zNP/ihjjp/KtvWVDOw3py65cTG43ecMVg9n8MoCB9fuxn7ZUs4sqpyx
/XpIRyJie/sVmgiYhL3z7ruWE5HKTKbEEwtJi7CaRmoTqrqy5u1Q0SftYjNX
WEQxqM8ulCMhViawS0RkExcK9/MaqFsk0osH9yooLnTPY7BHyz25etnW85yX
LwN/FGOBg3FccYxi1lsc++Nj679VVCOdz2TLlQm4y2ZB+YRDzbbGyWixEb9z
MFeW0CdQiADncC9LPSe5C5q4DJ4uUD/sSsabv23roTnDOIAR1AV0+FrJEEx6
oQck3RT4DpyqrOwlINAD0HyAtNSrNiJzK7UMpM2oZMqYKhuBUKjatoGMJFBl
gb/KPq4eMtINAVRgL8YFj+ERa6yBfgKNkSkXgexktwnG5XFAbhc+9rMThqX7
02VMDMyt94Z0AqJ0RA6i8STNodgBT4G5U7jXOkxjk9H+WI9auvb2uxy35cQD
C/op0HpytlY81O5ZBz05BEkrbV/TBvHzjwhB/FXR8xirqSWdNYcIDNWxrksU
cYSkw1Mx6qV1z+7+hiYqCkmNquHKyY+jt7ffStuh8Fw8rGysPWtkKlKx/j7Y
bySueEHM+mo+3pev8ftSx4iVcGs2uBuUT+NuTEPPcd7VAWdHHkQrn9E4NvcX
uG3AG2rD1lqfh51dlu9PXg5GRBzrSTY225V4sd+phMoEa7pb/eLU6xqilMvI
5PQhPcsDIthAQ5ig7igkPTTgF7DAwdddjDt1Fsh/kXK28X0bW60S8Tc4LgkX
e0hWrTVPSso8/sLFp/gJM4mAeexTGf+D3/zLAfM2tB7cqq1ow0ZE+aSgSlfD
xMtkbiDPvMLOa24/gqtcQpKxdMZwH3Zak8ZfHd1NzrX2BbS9i2v+niR49U/Q
eQJ/0ZPXb8w88RwpMDR+s80fE4aaCIBaIV/reXIrSGxgwm48zwr3GSB+x5ch
c2XYIgQKWf33rHp2pjKdjDOZavop93uZztSLY0eFUSDkYnu4mVwVa5wAHcUK
YkK0lX215RpXG9XULeDlsTAV8kkj8i+jLkxFDwHi6D9H5I2q6IhPaWp9PoP7
aihSZIZuHtd2atEvPUJZxVmmFDDK/vyqgZeWiY3EHBN4ut+cVLkMKTSDVH03
t3hS2fQO94oS9p0M84abau5KAGVcQLzyCpaVOb6B4DjXLYhopr1L9sZCUwpq
WMOcJDQFRPMJ/cuKP5C9dYj7kEihEmRWFQq6d5P+bLC/oXE26ieI0SQ670uw
5d60OmVlaQu6Ldr9/M4QqLUc/On4Hup6t7tY9AYOLnfflZsf6PTOONSzH2+n
BtuG15lA8Eh+LdM862EwLn7F7TZ9G0eN94eOfRBRd0LUWwiZioCTLO85aamb
zdnZOtjMbfkYr2Xv4mLWbPY0EJF92aidf5VauTSmQ9kea4ubBDtyDNr0FOKV
p91qcfriyU3kv1Fo6x4uj2NVQENRC+QxdEOSAQd4JlSKzcIiVDcxWmUxoage
WnWpOneZZlAt9+52CHGP5GoT3MMmH5fx+1oQwFdGMhSgC4jqbjKx4TUahY1K
3vwsc+Rzs/mXCBO+ozpQaMKf7Iw96+31QHff1JvsppuJ61X1BoqKMCciUoAd
UzVsMgbQvPjNaUoMxEwHXby+Y15XKVNdDWLS14WE4MC4hWa8LPJ7npHrQpIC
7/HBr+gvIdtdPLzs41oSFBZivubnvO6Xu1gVIjubR8szAAg8/TJhMeMNI4Sv
vinDrqhP4zphxuqx0aDhZHa7dnnb3MYOYRZTpFxjWdwSPrfKewysmaacec6j
+BoN2RV7SpJD8eA2qP+2Jn1oKUf9akgLBDau2QzLvbL+/SQAF3Sv5Wwa0ASc
v9wq62fK1EL/qGUDgfnBjGg7YzP0Uyg8gzv7oIlzofyHPlZTVGpSdlFMY+bV
YOeI1/vmWEeDw7dOmy0TiB6/UkZuK8qhDKeG8H9xpLszfPqtlFWXpsHFshcb
3s4KfLnmjB26dsMW0Yo8WwmmR38IqcEpP94rmF/7ac9fGjjM3yD3hmOdxo1j
/8NjPGkAMBgf5lQVB2nTa6fCCROomE1UCZQYV8rECNxjFRzq4DFrkAEF6QpN
fSYleVuGJPau7nSFde8PR+6X2BHWieIFjot5SbnKI3ONCQNmVXQL26CgXsMu
3xLM86HStamccYjUwcaAsiBekK5P4PRD2I0NZ/ciMdifwETeBzC1HRIL1jkc
70ka27mTycOceWA5/Cvx4ZC5C6eXO/3vWtHvsE1tSqvwhUPeJhBlRNmX0oIY
YyqFxeWVZ+rCf70gJd7//8I5Cju3D8pzbrqtjiDniomxw8+6gbyx3hHb1RGj
pVcD9x/VHBcC7wtuGt6y7jPfISNYA6AQ3MNbf+3UZ6OzeCXluwBx3BJdFdwx
Tg1YOd9chqzxqMVfOxm7fPT9u4oxaRGk4NzmvaUm3VcGdr2IcdECVgO6jpHr
4TmFuNs2e0xEb+Y25ytl8bFPHQDvttOZ87hZpxu5bNnzYQgNCpBI0Ua7PmQ5
0FlODZ8DXZ6UsAfXh+kKTFQ0IJqARu8+lIiuE5sv4N3nXBD0NKGzrLw7221D
nnYqJa7NHj+1rpSX6CdPm2UJoPnQv3o86PHIGUQgQ4d+CcHRAuxTfLtf16On
YQZ5jU4+Frz8oU6RQemyMSdW8gXmA9Pnu2x0dryCxX8FIj8owdA4rPKDYz9P
AbCmHymz9C/dRq78Vdf0Cl/rTNrVRmRczt8VA+SDwarvM7mLs9W8hqTyuE6l
lrqIGaGpps8HEe1Vc5B/Ky/Fp4KSXJQI0D1WGHpFZSJvPrQPCEO4yaVDjOed
bZ2AHkW0Oa3zoA2878Y0UCuNY0pRQPf0zcjQC1kn+60h04eYBD2jydOhe/ss
+0bgtTI6G7t47mzjSnFqk5UcNZ9grHs/TtdxIX8c51pQVRpOlJdSoKEj359t
q3ss7JNLfEdoqw55AHD8MeanzWgYRp3I03cuZ8EKay6sILdfTqD7HERUjaQS
KV2/RxR17CaRQ4SwLStiQXyqN82fw1iyLxlfMymvy7b4RB9QA8cdOqJxfpoG
HIHs0a1BzcPsVfD7RbSS4h64Vl8qHEWSaOJQmRw+ULrr1JH84UGZ8soJGKM3
AbEMG6YBy819bubAJBQhKsoQpfUM4YQP7/+QDrCdurY9iBv+bPH+ZvRVkfpK
2N3TkuTtYUtsrN0LHRB0NpAYKCKPguL6OvA89UaJsyl8gQQvpKmU/pytOe+j
B9432/V8BnANjqBGBAT2I5J5OZ9cdYaqpWqtUbwug0grbtam/icQ+LIZf/Bu
5cVGoFs7tYqlbTqmpr50mJBy2nwj9+fbYjxahY/noU52sATJkW6/O0E4+U07
oSqfW9ze/Gy7tCm6kt+XGHsZWZJ96gEIT6JJniM+uxDUBfLQ0AhneEodrEYn
P3jl03FCSsb1yML2QVD5XjWuxVyeUzKrAsAhpKD5uZxCQQNLWg/+5LOfWDIe
RJgLykL4bqEK4Sqh7B3ziy6HfjTNsOHgl2aSKcfDa4mf221PocTBhyC/pxUe
xRHjCUd0FR3rMwFD35bX3LChHtxTr+VIPb5VUFh0RI8/rk5AfqlcHNDs055+
OX/tFJ0YBbA/aYBaCGQgZw1hGS9IL+5BE78VvYl7XDQMYNvJ9tgGHOR56CsV
NFjscOVwHyakUktTGf/FmIpY7TKO/btTesrigVXuA+HGO3Zkr53QDmqh5o1S
DnctUXvBcgctH3sjQ8zxWRiZUBlDL9ZpjJYiIGW5cuXpdJPJ6EeJGK2iGRtw
cKbjWVCYSOn/lIADnkoutTJFDZDZUBWsqbLqOz4+cRTazOAk9JmKvDPS6dZH
E975AolkbZAZqVs4RcrzS7nf86N+aYwDo5XrC6OZ6v8ADVTYkBg3CpHSNbhW
nTZ5aq4BNfvT+FCXP5/oWFA6Nr9NlXlah5kknnYuvZ59kN6T3MDMNvxn3D4E
LczmVD56hBsur7ONrxTtQiQf1Ne45ifSo0011Q8mnZKB0r348DHXXZFJBIU7
pmPaTSMFljjArs2zpTV1j2IEjjFoZ1dn37KQAHZkictH7VXK296YKXtZ8CTk
rk84k4fz0yFXRSCPCY0DxZyxCsOMt08vAt2XQ+UjHrGPX9oSVSrOWM9/v/kN
4/0DxEn5YXE0OObk9y5gPsALuIHy+x/+8paZreVam4+drAo1YMQaa1TDDYw0
KyL0kyznFafn2ZhFuzgvuftl01qTWEB37oBvCsImk3XjN1dzsYOQq8wD+vZI
Wdf8tVZLRcegWxkEEkBc+NRfgSpnseo7+DLtVNM9+34EhY9jmGhDKlm9TZDT
DCDnwMU50M7SymbhkggcvuZPiWLiUrndDs9sBzOSft6n8oqhV4xmDM1UNzpn
SInfHeTdevJ3lSkWkXF3AUYJs8N8dWvfqgAuz4jeupqIokil+E3J2ps1wcqv
wj4va32n5p7hy9Ub9Iw+Q0fiUC6KW9uBXNk7Vh2QCez1nO8wFnEEcT//vDUb
dmrHdRo/lpS8eOORY4rbst8GWSIlDvF03GafpaL6x4aZpLjrejw7nhtzyPLN
j88KZbWvEDeI/jaEDh7vcegDMhHB/mBj3Y/LMBxTdTXOPhDXa+ICQEoRiTag
ZLTqifbVdrUbZbCS5BN6kAPcdw3v+uzKcuWuN3gB4u8H3BmrwP5PEtxGKO/c
CCpQRdZbIsz3nuLbZ9iHtNqCd7FfFJdxj38xAsmtvEvED7Y8oU6xgDJcuz+o
kZX6CESrvRQxnkgSjnMjJmXkArbBnjDN1oOl1Zavi83Qp+rMa0erKmB5yHiR
UqJUNixLc2+NIlEBBWk1j5UixPn7P2097Au18Qo3JNZKczzg9wIjQ7BMCQ14
Cxoa6Mlu8QKdd+cGuOOMfJ7kQ11BzidK9roiysxCWwZMUbS0GFLxWGi8dn5G
S+wyTyFMZgjU8g4aRTjH4PiXNoPSywpReV3uB/TqkJYQq63dQNT7Yrf8r+5l
c9TtSwwbpp1w8qTfmk7c5hku9UJTIDgIscnXevG7XNHRpZ/yJJGPt74n/dU8
4C6f3IC1vmEJGGYt9+r9b0dcPDYo0stBiP1v8szrSYkdA+bib5DNMm9qZHo6
PT4ret81bK6Hme8OzIT/+P8Fh0JBkXj1yyPprB8siocCRl+5Vgn5XrmRYmfK
j4FSPUX78BM0SmEo8wp+GEtJTfmjfZMEOcLsg4ZpeRUW4XTWpZtzPOPzs+Q1
aHhbpZMMt6bNzxEjy5llqmpuPBMYDALIsOkrGdzMre2KAZ1eo/Rhn8reAAV4
3UJlrAj69PZp3+62e9NyVNro4oBojJQ5NDYB1VhFS6gYgSzoLQ+5JmCuEM8H
6xzjE4PsjKz9z54gpwDlhFH+4plIK4JpWe7fNGcA1dmKeRArY4xGaQg4ADy0
7lJKWNGE/5wxP5pkXBluX8l8XPJUKFwVdobRh8VmxQqfC44akUtg+hp1pGjh
0H59D6F6gs3f6mxqown5iweSb62rRGlpQjlnmgPQ+pKCPiPmGI6KQ1Hjt3Ny
twmLOyMFiWRybXGqvsOVKiamAY2SXmHkvcdR4DRLfKK3v4SU39jqqb1O8DPn
O6pslZ0rm83RSBbYEfLJIbnUAnYEVG1C4hinr3FecVFBKIev4no2OYn576Ud
7fSNiU5WD0vqPBXQ4/pC5YSvwdbJ71KbQbU/MoKQRqYp4G5+3eX62FssuDoj
CYm+nuQ11ImGtQV5Jv9asWH1OUJtT9eq5NQr/+Jjvazm//kBx3PlLMcb6lgR
TdrSvo6QkGX4AUujOWo4oDKOoqjRxv3nDB3pAL4J1P86/N10KLrRyPYzy4mf
DdW7u+N3UELdi7i42IpUK7hlfw42j73d9RaOA2Dflk8iHYMx+W5kWEUjXglK
4Lzqz5B8ZpV8jaFxnPe3zI+NLa9EdbfeyUI9HZxG5t4t0LfZWz99ryQokVi3
vQdoN0y0VY3q0YRfQ3zfqUpDg1x1Q+Ogib/ilx7TisClNOT7rxwdnJ33APDe
G2xb67+AUHkqAoX3gknWNv6kd//W0L3RrNA5+t81Bp/OU4AJw4bzUpklJAYt
e8ScJh4H9n/XE5GPjHrPqVo2ckPz6nDRunIgVLC5JLpxMcaQVB+iRj0FTX/J
sLUszINkyKfotn9wCSCjiAYqV3Yr1rv+cURwpwj6lOvl9IcBeEdwloN11czn
wYLlExkFsG4GKcfOgmCn5AulrHBA7kE8WkJj4DOirhLkImjWYXj3GUnz8sDX
yP4vlajMBF5Is4DlZQ/mQjnv3JCgA0ZnQ7mwMrabqb64Bwa9ie8mqEfl4Lgh
wxINPlW2Ip75ZyNW5SCmyPbSmo33sSFqalnS1e7eDufbKuQqJEAa/SnnIN1S
+tJmh/BNC7xB6nhJZoFj37bOHhqJKO0BZwePa7l5FQXPPBC5LHX50So/dQxN
H3DHGnqWSrDmnTkpbh6BDdd85b5E1r91V/3usCWInIRh3C7lq3ITsP/+wXpu
rOvrxWqfM3RkG53nPvtynJ56aOc3EUlesYQFl0SjlfUgC1wz8PImVXEo+QJi
9NkhEidfPZAHOSfvNJOPXMqy/4a60T9MHlPDf9iJKeLaB2DhDbdKbNDuH6WJ
7pThKT9RF8EI4NRSDe2QEWG2Ii8dlftp9khGZCI0TF/qahbscAL2siC3dbXo
b1e4toMjNBdivuaZlreLACqWOcAnRNTnBw5/FZSmVQWH6mpSXasx9+CsrEC6
/DnCpRz0eQ0RT9nAwSssfeEv5LEM+FNIHLMuJ2S4a7HQXA86qraDFePjM6Bp
KE0uUpgxw+p3+/Ysw1NH1n6WEl1KrKOqIig5KJ+FY5H2xvTvcBmTcOq9iDBh
mrA0Br7eDJt1jHo1gmjtnqz0SWYx3RpqDvyNTd9R2lk6VKxbgknGzI6WLSGd
u4nAVsYaTCBGYHSniYhQDY5ObctDjj3KH8yEHXuW7akh1U+Wlr7PDX5w5E8r
5rcYZO8hKe0UM8PSJP9BgrrVYtz18HXrnA3V2XUSDQ0jCVzOGFr5BzETT3Aw
xmzxPRXizYcAs+Z+Vb5JNrZ1xYH6SOi/Qe8I4FYwcwRXjSw4nJTU29uZRYeB
cD19qcvAGCW1OJR7QxzkqzGudVYd1L50TpUN3564w7bHflERLvDhXHXgQxa8
p9louiXDfqUjBmHb0Mg/1z1m8/Gbqems1bZCsqcqfKMrmAv9xYzmQzozRYhD
T2Thfwh43sKSTd+mQW96a76gOYn7vG9BSjW6aDK6LFKbwHISBrjrcghRc8QA
CCPCY8bNr7ymbbT54S4LGNbgBTbeC1S7FbR9Gnhf4LELY0zOq8PoscL/IX7o
Wa2hH0TwmCxQGirm47USFZTlFGeRuWbNLSezAmDPtCpD9ia72c4uVwA/iWTc
I8UDMGrTXojAutHN/at/6754P7GCehbC7JMyDuIw+O3RXgaTkdxsrcMWopNo
EtFVpGaLJebF1akIzbLyMZcD+jDJBk+2zwyyqn5IRe8PehapF/LFmnsXnMHC
8WF+JG07fDxne7xxto2182IYP6VMbQoz37DJaFgz6d2tC1Yfdi5UYRWqOHqV
q6vPzVB6+Q14pbXKg874G1PEU/dqNfHJZthVOm6QQqGErEUEMB2zq3jLRIPD
8N3K9336LS2negrjTgWufSs5t3/46Br0MmEpqMwGW1LwbKj6y+6ODzNTSEnk
dQnUGXFxEIr5669cv/ubXPC5j1t4lOgA5TmfrHFPYELJYLrQKLwjDUj2Exz/
aHhIyD9Ig8ZexglQA2JoxHEVpI0KCujC6Pgk96S3TtYlEl1v/y2aaDUs9Lb7
8oxdwfc145JQTBpGj5hwWsP3SyiuMqoOAq9zX7JRZZl8luHceenXRZ3cfFoH
SWxRnOi5wVVC9SrMF1ogMtalQAYL8LnS1IT8dft4YQUSQAe2nH5+sNizlw5J
mhI2EYFr8toOyv2AmfriIVjgl6zmX3d3Xks6Y6xTBWATuGYbQPkWZanTv54s
iL2ghUCOaRXxPY4xqKdKE+Bba5i1Wp6DFe0eI5B1Lj659kdgkgFs6EOSfKlj
HXZ0XmeuIIKoUcoI4qXON61Qtqr8mzC7A5MdrNAsnWZocEYR6wyxvA/Y6CdW
Q8xf7mjdrYJ6O7hjOIicHPzXDX0gqILBim2F3dAKB79wa4RzL0zFRRIEp8ci
EJKjPiytKHJ82w/WdXVHg/LkFndIQvT5uFpMrIAYyhlq23A0ltaGnfjRFqVu
Qbv9qV0pMUQvBbC/ccB2Ja+bhQ93avPAXuJg39hYrK2byyFPnb/cUvs0MQV9
WnzhhlxebfCUd4+OBe5MnsklZBb48wfptmOiqvwrcuH+6F4urTABD7/iYMIu
eybW94OfL3t18N3lmoNdVe4fBCbGS2d0MwpM7rj5Y8LM4TRn0qgqHz29XRfe
XZfVf6IqUKdL8/13Q+z4x6+34c+CI/LxgSuemQBTSDH5zeOprEXvNZgZm7jt
vwwbst5ZBivxqRCbnA/bKmhjBeee2n2z0FiYxPJS6LZESpkx+8jqax46nkz6
SyUAq+uhqBFzIqumN55XEllCvd154on6fN53G5rx9G4+YEF5HZkSnBeJ21kS
DaXMi0s5T2m8wELOnwPnRdBvlA/8Z1Q2eFly30lGyk/LjJpS7uf5t45pq232
mOZZHx+JhxnH1mPWVZzGHT5BqrEJAcZ5Ile3npwMkBuro55X45/1N8s0XN1k
XYd0IM7IvW2NdLqWCD4e4R/xJOGtR7IfVJjsJ6Nds5sooPNH5S0MFmbs8CQg
4EJaNxPmVfnMwlAx0dB8agnzDDLp5wp9kBRtWLBa4oN1eTHPa6674X/TwZUD
mTYP3+FWiMXYp67CvU0TQ5GU4eseMc6IY29657mjSACyxMh2jipKZDAt5Tee
31tZ+8FtWdhG+OsMJEKDrq6XAdBloU71GjrNrmW9XNGm6Pz8HYCULxTMl7gd
utoceiUjHZjnSwlZ1aSToueP4QJ+5PekrvuHt6zapzZ1KuyjIQaI0PqNxBmk
CXL0GqE7g6pNGgnTtC1oVnskUZrtsDOrliQFq/uiTfdn6hTQvnyhV6n7NuTE
4FcBT1Qral1gPgXQEdbRjX34sNez32yOgy9sZM99iVknsp+pLajCveQX135W
waFyc1yu29icbvGR7ohSRBm1iKRhrmdr+C9Qa6zqhWhdpdA9W6FOlItTn7xe
OzK5KSu8gyLBjqJNlX+W1odDvgkfjrCYAc6+Yvx05u3gRuXB9iERovmWTOqV
PC0IwTUTor/+M7xtU8uj3HklLdflrjfTqXpvTo0tNCI31vvspgWMbMq4wbFm
2C5Nfvu/mYvf+a3koDUebN1lLUHd25WMiM//LipCefCua2isAn+Ors1A9A6q
Npg6M3P0IQgcpgp4FsxLDJT5shuz3ZL52UQP3fhk0V9E7H49ZLVm/VMOkDVE
aK1Ms67rUhpZfcVlDrqXxx3r7g3u32sqa7GxwxWdrE0KxBr9cr/k9Yo/g9Bg
w8EmcWAYO66DGKpw7BmBq//3Xrmvx1pok8pUtsDt/cZ0TRxYlFEmoUuUg/f6
0+lnM3VCrMqlvGpm7w0im5giE77AEY85AxpSBottbwZz8tF81+3NfQVnwBGn
MMCbZtUfUEqD4gF71nqz7buzsRvMIHszlwnuzA8+sU6W/Oi8NOGq5APVpQNM
6JMlRhzxu2TThAnpttRNxIO5o8JHzf36C3qbqd+kOK4qI4z9+JrR34TJKCN/
/0xHYf1TN7lc0vyxOcZtQkZk7IY0qRKCjC80IlNIFbdRQflxVLU30evbrf2S
0zdFwnvCRfVDz+Jf4ZoT2WCLoW8H5tkg5JI6J/eBAzfbAOM2nBcjoSIn6Ytb
Chyhbp0SLkDKtPvUckgTSvCEEoBKgO3khQ9ggXoi6KQE/sqff4rFmNqDzSfP
6Hgb44GghoEXKXgA53RZX/TpTGaK6MfPujkQOUJfwf0TKwlphR/F7BULNu3R
emvGkM32Ac6mPt+1ywRVzzDr+EViis6zS/61AoRN+tqMYMcS8GpIQp3slgAw
ZsSoac1jrx9VG5XUw2Ob8L4Gl29TbIH9KcjdEDrzFGvcS/+N4ZXl8l4XL/yp
ZVlHyjfiBsEGdhw2jXxdxWJEBpzqNHbFXQqP/VnwaPGMFFemk5hvPY2M0nuk
6YHNmK66TuhpvgMC9R0Qa1jUj0tnxzyKsuMbo67QI16RpgtoIZq940/ag6W8
m9zu77prKqZLf+XLT37rwmKcYmnZ8tQpHGj71t8cNj/TbM5v+dE8nHOJD7dP
eBqA+T3tiQgwuBl5JY5LaXeI/uQdAexzyu5StWN0pR9n3mIAJ93FtKpNSk05
EY2OisF1WVqN0R/xZwr7ynzpr8EC2VpGLSA157+i6v9z7fZk2sLWrUwZ/rOC
+exKDM9eVaem72SP3okBCeyOV6I/db8LX9FHtafM9DpT8sEJDuzSOhWD3HR/
wE664m3OZ5Db+AxJAGygMEXXK1lqhZIphkTLl+sYi3O09oprlG3GrQ9cvd2f
qpERy0zghA8V6KJAiKw0Qqk/vEQv0NzvoiOjVehwwA61+T1y1EF/TW6fQ7/J
Dt9Kd+96GwKgRyisXTO7gKkuPTs5GE9aSBr0/ekRnoMD1zBjJk1AepQdjTkO
+n16gBKZhZw2PmYKeXoIcEyQlCDIICPEuYNSMxwo3RKKKX4oCTaxUFVlGUCn
9vTOYoF0b01M3inRGRS9iNoFu5heIV1SoXyK1yJJ22aQEORFQdhPMIif5jP6
9g9d5+2iq1nXt3cQC2U8RMc7Y2sk7Rz/WPAG2qFjTCO1EdQCeaRfdj+DwYMH
rn+hZN2F9NjIGN7O7ZXmDHyC/Y0KMTXbHZLZ0wVCHEHojxphveQhzmd/KmLz
tg0UgRdvL+/L6cAwpH3snMmALymtdp71jjbv/THbK/NGGH6VwNtUmq+8LC6b
Y+vE0xvQX5QEiP+BWGrHfI2VQ2aG1QU3VXCuRY2wJ7OPagfRxj9001ZtPzUX
CXsbEv0AgWpL/bTaDaleaCx0z/2VyAywPWJDVvVwu6IRaZbg88HoyJK+UeC5
d0z3VTx6iWrJ9JUHFrxrkVFHhKWiyThEUSXhDkngHPRNdM3ECrIJIrPLcf4V
48Ei3xA+GMSUwDWmrvV9bk/GXdqoAwzVsSKCuCKIPMbeWKlbqsiG3LJmL7vc
Ad165E58/H7gJ3HnFFwvL/F8+83mPuv7edoHUkfuwe4nOTiAnHOMiXcwetIZ
sIA901hiOSYe7eWKr7G7MYw0gNAjdkg80K3veFKzSsk2gga8neLXRiDw2ZRY
oaqbIE1zryJ1Uf9zv5hBQBbRd72DpMthIp7+3qoRU+NH5k62zgkmtbRHkxVL
Grzzf+diumug0Xk4fhpzWzgJE/SYwQwP38Pu/GfzT/B41Dic5earSKtTnex+
wxAJubnygZdIjc4ipV+s1fyScwizg+EheRBG5B8Wqs92LXI/BCKRjgJRO5wZ
hR5CUTxdNodbQOqylW/6K13sON5vvq+MhCIU7SVh5sk9K4I88FTKu60hmGJ8
EkQpZMEPzKGmFkZuknr31Pb9uZ68cyG7jfpQW3+hbvftOyOxtJDyDgt6Y4nY
B0GVTB+nFsNUNM9qvZLJPYtEtKIBwaC0o0fMEWyohvbSHPd+kXoLjVlc4b60
PKIyX2e2dyv60TOh9ffHC0zaSrLvQ3tcXyqZZf5pQffOAiKNGHJ4SSR/lPYS
BCBHCg0N6OqNBGLopv2FSY6OTv+bA6kZyXqXMrKA4vj9sozTWpEDOxSDQTGj
Y+FITtDqNlloW5Lje6bAsghNS5rRSXsn2YbPbx2VSE4LP+9wrgzmkeppZBuG
SfNs9KOxqeuTeUcBWabSjKm+kFexB051rNvoaiN2m+WDbl1ZNapPSREaKV6H
Qw2DeqJEiXXGEDUPJa0syU7WQehxhMeqOtW4x3yQXolh0mGfXA/a+fLvHjVN
xpZntTzCSEMu7ovnb7/GVNv4flosoInzgFWFzNC6KfC5A6g+8gRX7Tb3uFnB
IKmz/GH2480uZoHeBc5XbIJlyqKjOlGnFxz6X0wArxWyD4ccfuHkDTd9Q1FV
jWtPX8C7viPl35fOrVRZhw84g2yR+tMRZHL2aoJ2tNVKI+gotJLHL44x6sEX
e5mDOxFWD8NtI4fBYCPdSGzSyuoCrg+YXf4yGpgTsi14jkJ8C++HgHGMaEta
EbWKowcnmx6Ypntt8PZFtl6rY2sLKxjBm5TtIo3N4BBEk03v7xNhdsV4//fu
GBKItiwhSpduvo+PqUM2aANBDFBs8QOTptKrofzcuARvRFkBEiPrxlFnjC8T
vKhXi+aZoU6ikWXelSwca94YKcLn4ayqGf/QKi0F1fNrVKmy2AcLjfXmuuiJ
Y/jgoCMiTlRrayLlsCNM/VoQ79XVW4aQ6txDghM9jkEeNvx8T5+Y9qqktgA0
ku2vM4zkdZeYtSwcm0BU7/KtvjFYmZSIyByTmSEcAQwelqtwqShNr9Siw26z
aMW7vjNCfLFDFUC9VOCeAYI8ObKw/IREl8MDRzPhFnr+3YGTZznP1JXrlGs9
lruIW99hqrfvNJbXOTSEvoDTEwXW6NGgk+V+KjnzxDFi6dl8TSl81ZmP8mHP
Z1fXl/apMFIXyC1Ubsg07x7LJyw7etoQRXZQD4F45l2CosB3sPWEtBGrwoAa
1GxRC+wwPqwb6a9SZB1UCgGnhzkgkfIOUZLkiKn85JnHWWUKCnVvKuT5r9/d
YNwyGBdmK/JgOaZ0F9+vfILuzFujR79dly1dwmD7aXSN9Qo7YgWvo/7euD5p
lUjEddSOyUVP3qZ03XejwxyCFGFIpN/c4st9ojlHo4jmXlhGVLj4rXlbaaR0
IFszz+FdHf0yXIjwJZQGVkng3KXsrM31a0RRGqk6Xw2OHbYAFIA1S23vfBSA
HZo1ftFUJDV9zByIyWm0twrG73MfOzKoXrytVhM67Ynk7RMO7ujdBrdyuVVp
GKftTx2/UkDmC7tpo8xCcDOP8J9R2YwENEXXE2z8a6HHzr8K3Pr5b0Wk/sLT
3YL9mzWUlDmAcPkvmoDg5TcM//n3nQnie2M5hQFWSrGWjv6E1txaOLShf1xB
FwBB/BQSuNyCtD2wEc6mCwDevEiink8tB9PvmZtEA25mqNeeKLN4IphLkwYU
0BMlzzNT91yJPNsjWWGbMIyWviYPioECuig9iCkRtsJGM6oanvVAiDQsrqi+
93D1byDJ/XqCRb4T6bQVle5SIQh2O8uVOJGzxMQ7tKVN/csPYYtVvi+jaYqe
/bi9RQlqc54Y3oYaw39b6exlFJ7tPay6mvOnZMV+JXgsGaH5OYoyTN8t5vWg
lIc7cjiOjIvUVhv25ql2cCGHFmp5lxbQMhlh+8WqPeKi8VokmQt1S4lYZWqu
GXgMRqnMOwhKdtwPb8hDXqOo27XIE4w/8qp84fpdv6fjgydD8GBevq2z/WOC
JUWnmtH3Gin8+Mk5+QOiwA208o2W0TwpOG4dZf2OWQilwLW1sFtg902KrWrk
uIoUqLA2mewQwFdHeitHpuWL2R3nRNJD4dIsiqMgSggtmbgTp9gTCy9KsshH
LRIXJJMNOa4xFaMCJ6JXCFFCnlNQy09RhhjFKr37ajkPV/EeYqd4emXLkrfz
0kAX2IDIPNMjPqtD1ExyHRlcI5SWD69gyyZpRL+nkesHD2FmDG40ZVBSo6yK
VNcOJG+fR9DrE+ibYnGtl9zm/zXrh0Ml4RY+ks63VN7XZqMf5xkzKeyNoj2A
1IRtc4w3I/ixBlyjvv0ja3NbOr6oI0LcraSLIRCmbQsd2aAM34u8Mmi/Skvw
g51SJSVSHYYcKGEbORPeBIooekys8vc5E+hFC1eUZXbEIaFJX9yFFC42WO/i
VI6tSYkfHPGISeeD77OJHA0lrEy/2D30Qq8mwmWm8k1sszKrbrnBORxw0DKs
VFVsAPohn5lBHcafRdzqz4D+olz4l6IWEl4B53nNd693WuKitOFVl9V6ZG1W
5QhM88Q2f0Cdp5OcGb6FSfcjEL2o/CswDb9DrWf3kX5NUsnD2bvouaitT5AZ
Rn4FQQzztpqMECcXSL0xEv+T57GqE+thesuI38hU8fcynnlz0xmkeHIhPDVb
M57uZICnW+PTnhmkCfQ/zKXaVhpcCsZNlmrTCOaDzE12Q9Cg6EVKAkSZdYEI
obHSeMUdgR3t6rgeHaiT3aQr7QJLSS1HwaMLQE3BWKbOSocmcll+oZBHLAgO
vJE9P2EmyoHL84K5qDcwdc1NMoOdOLtUBBorUafVU8w8807ncERbO1o4ubK2
LZ9imAEkphvv8LQejAtJEvY6vvw2vHFSEAzYT7ma7q9W4jsM8gGKrHM3JUeU
DZsNnpXvP16UNcFQG47lJaTgbHKUlRv6XUBDfgfJnmnC/CIapoo8EQBXNglw
miHTAxqLa/o1ByP0OOuJv96z8AmY+Je90z5PUI9rJqGOy9McW6aSOaZf7n6r
xBlzKFnr035+k/8ckEqDgSWU09lxE8HvniNJDF2wn1ghOpnWbZj1p/c5GFW5
lFK/YaQhX8zyd/IP6wIqlYIdghvBpa1lIo+DaUyZ2gUwPP/uq4b1+i0uUiDR
OcQNmIS2hs1b9XR+4qlCGlLXkbKNIPrO6rb3wNUW1iQ1tDGvg4Nv4NBzwrba
ZdPnt5YQMyogiuPnQCFVspPeComA3SFSWelR/mbHRwg8Qadr+puwHNycZiHX
tiXf7RztRxPIFglp31EeUoGqsw8zz1MtOj7I7ahuG05AdosdxqygiLOud9R1
uJv1Z+TkRSfDkt/sOyEEhBpUlLGsBPySDehyImBCYJmYT+agqbzRe1si6132
LFMWAOYq4dgR30C1JI+ILp5XS0QIbuBtM3jlCzOLdlvmgaog6gu1LR0OqXu1
lORYT4oe0pvoNsyoRAlpDSND4vtrtoStt7xBA4H0njH1A6lkjOhEkSd38Qkm
xvH7LsdV0bGdQTZtt208VyjAV5cDmHWJ/AT+Qow159FLUXmgukflsGDWjC4F
3ctUy1pUvxtkJ8SplD9RQ3Dr8BwoVUyc148cKGiz4kT2LB/BLnYwrJ2BgzIM
mOvtRBNWVUEgQ3trOVow4vkgMIkDgRuZ9wAA6qdFgSBFaf9UWvD5T0YtHrJr
CDnYy+YDas1Vs0N6vSaUl4sCglq2NqKTzlNMdY+25O/LtcSDFmMi6vUW65Xv
7caJ2xWyKx4VmMzviu8C+17o1bEu15fa9MMBABCLwkF1XbKAHqfq0B7KF57X
uOxnRQTvZXoZ3nBeIiZDRqGi5HmCX+V+4uFi+pMf9p/P73WDrKnijLbQV3e4
cB3JO22fFbG2DM1A5EMCrwhQyzt5hMEtDmLr0mbBKMmLYr/6NqRtx9vduBDH
cmxUuy1+Rd5Z1zErPl7QgE+j++CznNxw0MSU4lw6jAM18Et4ay8mOYGbaOVR
0EG0MqUIvuwkvffcyZHrl1fI9DL3FuIbYr6FfgspWJTzXnP2gvYhC3tI59KM
deG5CX2jE+5A4/MiSRQp4UY7JR7uaTrYN3/IXQI3eGqunjhbxNi5NB0fYlji
lOf+qwtEPcGATMnM4I64+0rO3QJekiYEVFVki3xEMEZqlpbr8SYPV6x59I17
RoBc3G7fOcmO3sLRX7uC50Fs6jMYWcC+jipkz1xraN/FkjzfGe3qJJ7q19ee
Kh1MrD5Zx8A3Mv9jnTFdmpeJrxZSIujLEu0YMWSFY2ptbAflAaUYdMwirUoI
PauU0dMQUEKj61jIbWoa4sNgkHzo1Pog5qnqFNc3cWmjPudPHrAI6fyb7dPi
razZ5AbRZO+8RN/D8LXhV6tA8KqYefzMsvwMNKCDcg+MJsehFANFSrLhIDHK
6bBr6esxNM13D+VHQSUvg5FxwVa5UxxTdFgBDlyZslcaurJDcAoNGsIbVZoN
+lE0GQBRzgJ/Vy5TJ5DG72qApqiM/ZrR/QxGaEKLIXyhe4JU6dp5H55x6XBs
zFcQW58XbRMDBJ+tOTKJQfMytHvM9OKe8aCHJlSDo2eEbpJ5VuA3tXF3aYQq
r+JafJG76or/FKV3MSKjHZy4op6LCyuymgfc0Wwfa49+Xu6MBDqqcu4Bp0Cr
FkBS3miISLVasHVHd3lmL6mwHi0nDyCQIXtf6vgdfdTuPxl5P1t0KptAuWnz
ZhwOedEJL6kMf9+oBEAt4KSKQrNx/ehZAQjUIsXBrebFp0BRb9hCclWF9kOT
nGDYFweTNWeQedk0JpWLFkQfCVbFX9fi0LpyBMqjUUbxCWfms9TN3+sOUFWZ
1JIKPWheFGw9zavOpo0LZjlYy5v6c4gvYjwpgUtf4tuZgXoi1nN6ykLiH40+
n8AMd+OYudw3SnEOUJPjGqTL7VxtCdNzpPZIkE74Hh49ans9eNzp9eOB2Sfn
jINpIQV+rdiYIlNfQI9tHCS0pE5METB3768e8xUd8BNkiV+IHmyephfpsdcf
bCVyqItPhFY4aB+0iSvwI+RID3yN9JJuguBj5Rsecew+1o83whdOG5w4iInC
s62m8boTlwIBdjS1/xnMjWcuHakRyarMmuBGiw5h7f6I3X2MPN13a7IUhowU
Hg+a9EqV843mjJgcbi4pLX9Xj2Ldo5coeL1q1t9pbByKqnpIZpVS/nsfG1sU
R3HFzV1lgFpUAvQW9szRP+llKqeNY2ea85jSpFwW10UsTQapYyRc3Av8EHhQ
UrC20QH4Rixw8WmjLFJ+ujBcTDNn2BGlg3LnwJENpRt/ADBWGScI9xAtGmAB
EI9nArgDubj3d1oGNZxCEOJCESjzBfrhKBNgpEnLjgYMXCEauAEoFk18CeBE
YKATzNuz58YqM0Z9RnUKzDZ579epPnBSn/08KfP3GfZonhy17dkDpfxrdnll
0KzME3Zdn+A6MTRmOmONd/Cdc35FiW0H5TTVrioUD0K1rrZ1Wb4jJTfR21s+
w4hwyKLo8H+7pOI/2tR8cONg7P5ieF837vOPXdDlvRDMZK/VrBhlaTpVkK68
Ce18OMzK23cRukeTA2ziPhM5jwuW3QN7No7HcSQCPkPndDDBjvxReKXthSAG
+9tbVKYicGekFNT9jQ3p0Ky/w8vU9u9dkcuzOd3xlRd4a3mAUdhFkeCSwwJs
PT/nXo7hhbuKuLqiPglsMDWf4TnlWhYmQADjuAxGp7EJ5Vt3cRfiQTZirKuY
efNrJuGAPAfltA4Y/MjSS/9IOtNG3H0/3tPP2UmnfRZGSmekHf8XVGyGPN59
ZjfRBtJoT/xby1VSX+b8416CnUbS9Z2V7KP0+396Ac6BeW1b6qQeKdK0HJyz
7rqazL79Q8nXy9sbV4ODNAh8b2NNFHw6LCvk2XbwVCjOLEBxtNohhizLDFOA
TIKIB4qxcjce3ukSluqOhxrBS7NOgzWP0UNFDT1MVIl81mGhmt4KmYSozcMu
Ren7/UH6ZYyzgbLY549psfKO0Y08So6vY3h2saWeCW03mYv73dtIbuVcwTk2
Pctc4bx8fEcpcKgyUdaHfonm7tFhZ5H6hHxucSErsBSQ3S4dDu6beAkNG7+8
tMS3C9mOHRxklPemz7oNTvbjy82+kSgVMtPBfNZtqqvJjxmDkE3Vr6y8aZ4K
4aBAago8ctobyr7SizpQLQRWxUDPQqER04FCuJ8tvxNXTA2Iv9tBlbHOjl+q
ezNyFaHO/AI3/LWQ6/S8E7pN0MGdKuM5aK0fSkMP6Smm2CVXUGFhfUAxebmb
ugyQTE/PPBfzTNYxqDFf7TlgcfGX3+6kfynrtb9In0YtPJP54Snu4Se9s8uJ
xMe2KkwVO2lj4E4FQUuhWM+++eYw7py5fud8+0hMdGtJgv/VkpNQFoWhNmA6
DPE5dP9r21DzVxtFMrSa3hujXw+3nSHL6qCmbBXwwKQnKeyjlVjqR0r0IDpk
v9uvUrDO+ddWxNtXt44EJ9XoxmkNP3iya/dAbZ6nYLm7JID0QzjkI2ZCTs+d
mQj1KxX9/Fzltm3lZfIMUaUb23t4yr9xMeWmrqc50qsASq5rUSUMMGY8apOk
35CYNKy+v1ZNvuo9PUsCI9i60HWJWZlfQjSIJxzAEaOoAIPqz6WibB27WMqo
Y1LTrJhj0AaPLVGkw8ji9mVQbsi8Xe7GfRfIEBpc3BJkE/rJtzT7ZCVMRQCX
TlFzJsc8JcDGwOIFYa3cWsR3jtzlghicwLL7Xvr8yf9ZZ3fBRSIb22KXUJ6o
wNHED6N+8pQWULtQxK0vS2NXJ7ndTfQrR2dbxqQxMt3viORjIiQPHrRs3+Hy
ScjenL3Su0YYeEef8YOYKzO/rJSVVW7p5CQHmRVgh56xYDl+fIikyoyyqKH4
7H2lIbwtRiZNSZ63YEiyMZ4dFITxjlum/GYaiU+HFNCGNO7WByJ7TYUFGnHt
n/rqAiogFV714A41JpJErrzlSNmxV0PDkdYBiihA56I0EmhcnYFQ2XO9DGDv
G8fTR7KgdaWe9Xlm0mOQ9L+se4Ehcj8RlEkg1yKtuQ1L+3xXDWQ+NEwjml09
XaX45fWYRDi+DrXknI3K6m4WTcm3L9MPSOaGdGq8Zpf+LKEDhwCXm3LF9Bdw
57Zn8OFz/K/YU/erKfub4UEaqusyKZrMSDFOodT0aCvNYWnKRBkdKwMV2LNg
MrrVZ7ygsxItz1HxkACt/CWXAzdMraLg/2NI+qPwHxAdScCOLx0P3bBbNRxD
sqj1z14hFxtugSWRPV79kQXUubWg82d9fpNenm7TV2FbdN+9Fn0obGefYq4M
P5pIuArNyKK0CJlcAisPFjbWXFeILuorglS5o6U/aUrFaWZ5leMUDAXQfw5s
9YtPBt7rjPGzLKFvi3ucwVg5plmpS+hJc4X2kzOclCp6rKeeVC/+JklaJHax
xmZT/+3tiWOFkd2O+QLcox1v+jXVgo5gkouJkz84PQVDs+FWbD7KaEJ1Fh6W
NRvtmfyCbD9ow1PiqaCaTblT0/raHnlt2B+KaxpLR/BqvKL+AnH9Zfux1zSd
g1utkm53YoqVIWNKBKySNav9oLGnlt1UaeQyjUL72lWdot7WXd78gc5JNSj2
q8ruY8W+S3VdP3Wolnbg4wRgwrPiRC1LI6He4L6ANYzgjeP+VAdOHcITuYMp
WNbFv8IlnBK6zWy7IA0ujgKr5DCt3+mvXkMkb+t2jcPKWo12BTfhMlTcweEe
ePk51/ymgV2ZSb/R3vvZwplOIZM4c5KBKaGjEuzcvUDoBmdnoFRWLkuWuHxU
60B9p0gHtE9yoY81LCuudtYIgMtu3zVwFTNtZ7tGNhgo93e2HRqO3YOtoiZ5
c0eNdvw0kP47wmb1dqAbrIv02vdLPqM9PqHP9kLC194jb8XIgWk4EQF9INrs
0wQif/PSuiACoU0LLPJmunLNt9DPYdzcUxiooNuT8Nowo3Gusa4Z2vVLEupn
LweY+mix7qJ2K997+0dD2YTd0U/DvnlPrTLxPI2pqTljwPbCSBQNIsS2jqNb
ChWUoIPq0YVAygFDMGa4N3JqixEXaj7Fn2/mrLjSpmbdk/iPHGpwrECxLZ1j
A65a+8rcF2ehP0Q+o9bTBHtJn/N6NiKgv56lBYZy+SOmltBWzR3dijEhYD1x
cTy/gHcvnMDLJuLZCczqCUiKVy7O9t1F0kEGcopKRnG5aFX1ceOcSCJmQ2J4
4pK44xfhro0UYmcusiV0NyEwmyR414QoYrEaGXi+W3Jrh8mYhaSUzQPYGtRu
a6fvQVVedlYjPwdqRhB1Lss48p8efF4R8CQitXdOzSlMyb2gt1eE9ZXwCEqj
S8GiWcquqn4XhepAzkpcpr/StGWb0FrOvHi/hYVFMkFLl1zuDZSkvKSq6dIJ
4i91/tMmHCQn+GXCOTzZ8H+CfNRhkgaS8nfx1AajB0+gNjmNfeGuNZa11KyU
8afBf+8fHUAzt5PcLFZKNUpQu/VVSc1NMkymUHq0KSThOU+22ffiJeF6xPb5
cBdDojq/iJKoT2leTqpyyg3Xo/nJXVmp3rGC819Mw7g8/qXAmPcGZ2xOOMMK
pnquNAxFe8HzaDIu+h6o7Z7ihM8rfrAdvWKElgWf8Yj36k23eretIaJY9yEM
5paYy5GpAdpdqMikPOjHQz9MA40ncyYJ3OaMUDpelYBPfndd65zOihOeoZQw
Pkv1Jy5aMnEqvpGLVfo78Qr20TauK0yb9aUdU3/chX7yzIhYhQldm6e8qgVA
pAlDoDo4WE/biGL1ElcnUxpnIRYH2F+qAaE3f6OID6LtpSrW5A/Ghgl7HeJp
KCF0ZlLj6cvp/Ty63VjcHo1M7ECbuQ2y/Ezy8HMPnGdImTFakhR7SqAzC+/Y
9aYnTisMSvC6S6fUkSs4Sar8/cUMyS9dzeSVZDuman7AVPRRaEq7riOlTiRb
Jy/n01kGjLJOaXl2tbCmCYwR3GFsLzFOdareV9PCATkGkh6x1cI8JmrG1B5L
enMsNkOiDjhGYbN6XnHdyl8was7atqIXPtJHSJKQmDjmSl0msWS0kONoLQqS
eW1i1WIw+m47MWCMEIvId9yQJNuhX5bLzbXiebKUIyvQyq8P59/+XLwWryW5
ZVQDxQidUvjaCCj7zoMjhD9IEqtws/phwZwWooyxLO5Twf+/drxEh+iaTj8c
s0S7oepQGs/6s9HGKFibgn73o9Pz5gdSsWcgIL6nXih3ohgaAzfJe4/7V0Pu
377p5swupQ5zcuuiUS3z+RVlrhKxKwMnjpYVGaoTFrMZaMYbB+PZAVuP6E9p
Gk/6i4Nih1ov5rYGmwwwCbuIWIGyBi0i76LImr7EFLtVfiQLLeTb3UsPtxGx
PnzBm1lmX0ZzMcm5qR7iaxRzBVBcNp0SlqcPWsUe+lf4W7JLdNU3jd7BHbUm
363EaG6QPqA4ih11HxWBBSx7r+UgWnhf/drMjXh44Olg4pLXqjIe3poB3x8v
OhY26nHGGBw11kQMPuOrk0syGfVhrKEX9iySuUYN7bJ7/UqCWSpcuyzdOmlI
xTvrz5NKItq9zlurYw/ln4lOMv0b4QAw7vanILdxLCTgwe49CSk4PuP5D2cx
DBCQ/ZyQ7H3tbJ6nKe+i+1RoyEOM0uXslajSKVCWWBi+nguQsS6+xX/VO7Ux
wWb1FD7KoacCPOEdbC/UFq6eoV6qQEtY7E+deOUCUaaDWYXx7HmkJZ8HVJy0
NKCACR9Emnd2QmwtSm6LFIGM7b5ECRw4NpsJIXYX33i9cw4rdy8c2b6iBlLz
AFS0x4P0ZnDXBKovbFz5avIf17LCeDTWuXJOBkuhQEXPHLr47sBOCL4B1DBs
5Yk5VOCFXAFEbn9doTeRQA0+JXUKyfchAHepJsbPAyk+OqP0D4K2L2oJgwn7
HElrKSSLiW3l6nHMP6Y5q38OksbCkZuFB6vYVY6JrTvLptCrkk/3K7z/8yHz
JpAwoRLzbto7PEZQ2QH/+iG3YFBfKisLBCtSTHdUNwvkCTf+4ECNOoP9Ii3G
aXv9OrGX6yuyYApQqUug1n/VKoqnhQ0S3c6RosCaMp6m6kksxUqXZgqVFoeX
AB7qxpz3ZyrA0Qftz9ETxNT9xuuE9cly0QsWwS5eThSbbkAQvRhcowMC/7Wb
2CkU2BItp4Ps+Ge5Z7IImWSA2pjAqRMEpotX/bzn8yfcFeEv6AW+cRNiluCJ
hMbu7BKgYtRHIRGzxcIIBV4Dp5AhK6Cf+bjX5JLjmtfFalaCdmHxhkW0bBhv
K+ebxy3UsC5zMF4tVUf6soRSCpjm/44E2Sw/ecx8DErS10HLW3TlSdrOWxcN
Ege67Wt1Oz2rb3WBs7zm3L/JwXPUJJcGv+VWuVidWh7Alz7bks2f3pn36ZSv
eY7w1gqfCBVoZL67u3K2DUbj/DbhsliGyFoR1pIOfzibaPCyQzHoDBS4vwxa
eayuQgkijNe+G8C4CW8RHbzfonMU4juj2+KPOjgtzS2ze4cynDC3yl7ui9vu
0TuHEWVNNqY+UIXsl7g0piFHaMry2p3taYy7E2XJB0O1WwWcugv+7WVbN6s6
9cLS0Pnu3jhI0wz8LLDQIj6BGHMUfFaTG7kvNNTT4YbhyXmgZ9Xlp0B96fpT
EwaE1+GgTJde9LPQrkvtxS57cwYzwLrFzuKd/TAv1MJghIRWGG23I+t5gNhv
vFx5ubaPHdl18wvz4QCbm+rNr1fL0SXpkolsmu5b8HuIxRGctVj1SCdGmQCg
V4f5f9p45NhUzkQMRzyozj0DeWL/mZLuDHRUTG9wS9uhzoCuwVygWNCFGmtD
X0lw6Sga7RzBL0uddDFUzH5yYm8KLtuZEot0Zsb9rba3NP3iIIRSDNzv80B0
Hqquyaj6lK4UpLYugGm/K6sOz1Gs90vCr8vRqDRTNRmH/Ot8KeZL86zMxMax
yJkkJTiKUhil14J505SzF67wgzDDz0AT2iIGegot0Bq730ZBY1gXE+E/jTjp
wI4VyumHIRhYJ1Xo8Eky42tPjaPkK/w8E4dulZ74V50N+44Nj75NrTqGvcIH
LGdDob75SvqeX0TR3AJePC3xVSOpg7GCu50wm8dNADPK11SdUTpfhALO4/X4
n8T8Jt0OxTNrBkGPno3G78oND2heM6YbiY82qEXFb3cBq4Y7VabnwoOrS6AA
1lVU1HuMyM519aiTLTijWSZdyCp0nXo1PXYgka0On76Adgy1a1a/2tMbMRSM
F6jJ7C3pHDG9gSM+7gzsZcFJoGPdjTaa7bgoZms+AYMdlGm2liM62HfmBNCU
fyp8dW+ND+3IahswPLkqjFddUcDFOLsXvNLy9iw1KXri6m///odM88obSnXq
Jjyc8Sr9Wk0UbHIoGgjNDH6piGOzXJjjSqTHu4KB8NCvZBVrWuTfoEQ0WfiQ
CpngrI2y7atlzegapup3VRXQC5yxO3G8DFd/EC/fd909CJhmmOps/tD2MWwy
kQDEisjh+27ETlr5TCflLp3xA12KHGlp7ZBmp9GyRyQieGzCKZ4KrRDW3lh8
BuQhgtYOyVdxiB3ntQCNMn/AGFgFP80zo7VKtqhqR+TxwhSn9sz66lOT/UTf
a46HttbCIrZIZn6HfwPSUtjR0sN/Xid6SPJ019PoMsOATyIgQgJ5Xs1O9t8a
KrTBY6VYljKU3oynJKO56prwkfquZJy6BXVzhX8DYo6gplA4xSnPGZ5ws+oO
eFRsi6rDgWAhl3lLEtGFHc7A2robwYv7BBg9xw/UkpBlv8l+JhiMahrzcYA7
whwmR2p50ZZZzwEVTRMMz99Dfza8GZ+PhcXJWygSujA1fbz1Y3b6yMwA9VKs
z2qUvU5h0bWBrXkGUODU6lzzp12lgIaXjOR+/4T8fnoiuOlP98YPQR9dNv5v
QfxLckBEsrzls7j+muOBCV82dWj5KSfST9rdwiyGjuybW3MMsdzjf1zLuxIJ
CF6gGNQ/gOfpLN2EzTwCoV8pz2qaDw+W9jmq5rh/oBP/E3JpZ3Q5UKD7mXId
2IAAds29pqJJ8IKCHtKOipckVzRPHH7stAr+ASEl/WcDwM3yI5yQXSEX41tz
gudFNZcOb6hSTNeV88Q3H+U3qNMkMj7BGp/e5xDcuMfQj9hMkbZwMJ4yfrl+
B6K73eXCgSO0vny10l97cdHPb8INYLyPZ0UvX8iK2hiwXvdgozWvSeEeOVcW
yNoBoMvudj+PhODmFqpjXS1dyz/ZTQ0kKqVywsK/AxHFDnPYJCS6hoKtPAXD
QmZn+Vl03laF+8pZ53OhE97jpX0vVi6hO8bQn36rap/86IrgTF7lX2ZZlBMn
f4pkbaQO189qvzn/CmOU1jlqtjudand9zx5AAuw0RHszjN3nrnh5aXlstK4t
wgUYAMwuu/YMha8RBdm535h5x/NyW3sqISCKnmrmJZsx04Ri2pPUqtD9eOTg
Gs24ca9yBGgTOSGPfhSTmzZYVqvUPzSazHZSY9xg6V6/jDgh8p8QFlQViM5I
e+J5zHLJYLjIeAlfwd9vMqXi/HuE+z9mp7+5yDg77rzQYMNiO+4M5fv/gJUn
57eV3iPGJs8t5egROupASUUJAqzPssdPraoICJWx4aqQLDl3glF5iMZldTC8
dvliefnq1Dj0KL4RUfZ7C9QUbSO/45q5GwirKNN3emFszmPLsn7x9vdUu2sF
d5MK8xue1tR9rj828mvkWpoWDaPiGiuHThnh8yADtKr3MM/sIZxhiy7rHU21
EsY6uEPj/0yCZ8fqby8rmUjljlYxe+VLqxvcF0OSxm4xNSjEIaEi7bUGCZ9i
oFxs0+VQPNfpvKBDlvBPHaZAyy85+SuTDZmxBRXlsS7Krt7I6W9VxzjUESc+
at7OJzEI1kyXQnnAhHPKyZnEyWcPf7d6YMyblvktFExAFJ8S7OeYMZ45ZOIH
HlIls7j8lUjC85hHANk+QwClF8/Dp7WK+X80kOM5NjZ4QchTknuOSA1j9pc0
fWQE7KZ27Qhtm2UOW59D1MgbLTRajhnPbr61WA16IYoEgwUVemwa60zbJil2
IgqKLQFlwM1sxMnDdZAZXFWlLvFZgqaHOU+NCBZmOa3xbp+9oGO58ICxtA6e
rRsKlh3+TAA8PUTS8+io+hfDdR1Oc0zfvzK2z+uUaJDkoNDxMKMjmtapxNcs
50l+QWgvCMs4lJMv9gQHDROVqXWeFXLAOwlp0c8k9r34YIEUlYtLqJVtReWq
SCGe4fpLx/dw9Es9lAyhtTYq4ZfaPt19S98fwvLkvt86BJaeXEIz5bTqwwpW
Op3f/EbqwDvJLZ+X5heeckHLrQ+LGd5kSIl/FrrRFnIqd9DEpQHknHNdNifS
GXL3k0t19V3snXT2Q7qnG8zp9Nt1k9dJ7909yjyP+0J8P/1gLlCwebHGRLpm
O3eWFlz4ZyBqVvqcOfLN9IWY39DenD6WpPEWJqtwcEFw/6GRHThHBkGxiBAb
fmgCi8JmKUuEKkmIiJHjE7o2kUskX433EbxFlTObg/TOaH2rrS9unIJBH7pl
nBy+EwOfrC5jl+zlGXgR+P+i2GPXF5GWqUs6wenfsLvu1RdqFEMpQ+zgP/12
gyY3oKEaGrmt/Bwbfpd4xWkEEzz7iU0K7NUpeJqJqNLtPRSx6rRxX73z+jrB
+3IKOq7+AXt6kMFbjbnUL3Am6k/5A4dlBaeaXjbP+z4X931w02P4LK/+7+/K
Un/H6f2oKhZ4p+fgP4lW8NjpqhG+0eW9IKstLRv22jnQX0qzbvLx4iSgGqN9
cNorDvYgj8ihMwVvgn3jHIliElC13kVnKTI/ozqE0qhVhOAq1Bzs7D5q08zo
pnyPjCnwzzbuR/kggZiHfs26d7DnoI4gJ3DvC3pfhOzcf5HzYT4UkLeAZfI7
NmmI4pko9iZ5GXcOvejrFsFUg11Hos/fMzlrbRWXZge4PWzZnFeaTapx92Qk
EZgwYmVzg+8eznXm65+QXxkyJfA4ImDSTR6a/QsPm0kJ4Pk4B75Wo7YFzc85
dQXpEqrp61TP/aN9wzSy9v5MYBQ1XKCz+NldwoeJy1ZiVzy9gFT3OBoIb7M0
5iElew8/3ff9Hc5PmUnSm0BKAh20YmOSxz9XYhU5Ngu8GEECYx0c4J3Jw9Vz
IVi+izXd9ZzZ1NIcTjZQOJ1TDVx5s4P8H5FRf8pVHzWIu4XmXGkXA6QTA6+V
GhW80E/CzYAPPXSkPagssPKvChrmLOd2L1ugbZ1q1/PmQu9/ItNOi4MZynEP
ZlxYCXxdS/UaJOKnvTwpFTap8ixa7sGqlrPHIogK6E5+AWh2ATnFbDHE6Zrw
N3A+F3X5sEF6SYPK5n/RKLpHcSfEjVqUmKo2JwLu7IpgMo4zIAlFvn5lVzQ8
6nUp/7L5527Hf5wpFMBDtBXkhAbnrbx6YcGdd8OM+0Dc1WTMlQSth47W4O6c
O91WdDt0iDK4p0Qi5eEbybJ1m1tcWflLBe/qXyXjI/I+oQRSUKfy8iGdX9Ql
LKBmL4BXzKxW6XtzSW+79OO1tO9/54eAXgPTiqnmZsuW+CGkW60WVwIJl2GR
MO3CCPuJOxria7YdfWHv8NHzd8MFCINPQ0QT/gu4/Qy1wRlxmc8Mt/s2xMtx
U/m6lg8BXzkf+NqfFS+9OBt+WaR4qzGH53pRTInDZA4xSFI7hPwQFXEeAd5C
lWciMV7FEmiNl542EA87xrnZZzYlyEqtwKbayFBm7kZU7peKmTFnpJYXyNdn
avbj04UI7UYDc6+dPfX5ftDtmg2U7ZqKiSZnbtHEXlNIpz8yhvcmqoxQoxdk
WVoLph58jng7OONOJyDigFuNJl/2mChhYx4ugjlmqcsAQq+b54IEl0pHtMFi
3tifYOF0g4bIHY9XrCvscpj5tHacBWSbeLRjXO+s8nsPBE0K/zqDt7cy7nNQ
4lNbwAi1LLLCFFBwb3Zjg8DsCWcS/TChmgzmrdUeTC+JhFyXV8ScSTbwu53/
6Ti86Z6gh33ww8JlwHazWhWa7HWLFduRCqMkI616PGaxyFQT2ix0xov50Kcf
A73Gx3p9D/dcvj//HIrrvN4lbONB7CAsSLQWY9+pENCoXldfzWs4uojLMFeG
thUHw5+IWr+B5bEG6yvMMVNTk6/1n/gZfkHdb4fWmzoZFPSsGWnksmf2M2/l
otnkHhg31CMbaHsMJ0oNIP+ImE34UIxYxvGjbhVCgPhY1AWOQgfxHfEqougx
/idP+SaBG4ANvLY8V4ym0FNAWCvoZG+CJQCGt/xwnm37bQgyJH6+koP7TUHo
cn9V847LKWOrWnWoDrF8GZdinPc7RXKpCJBVjVM3K81x1oG4rP1EuBeLP3aZ
LLtJdaYqp2gRwSWOsE5R3EfPJMAAPLaz1d4DAOGRRU+2TyfUhy18blzSbSMo
r1rxEVWCe/eR4zaos1SHgw4L5UWEBOJ7jORL/HewZ3ziYbpIzUIgKR3vTUrc
D3eYPQZDsicZFWsPGqZdmDpTbS1aKVOID2wJtPkZCCtC1023xO58LYpD1VAs
BGsg1xR2pHkdu5mOXTLWSIPkV+R2HnrGPMKG3GsepXYXmw7G6Sd+RK4btk7b
JeQkxzKAIxH4TQI68G4GQAqOucQHHT2CDwWGgmbSnXt33Hb/CvR5Iqm+IulS
vcqVikIO8dRb4O4QvNPFSCE+cNYvGIoIEQ/wnfLxMyDtwpt9Ba+VgjlWWAKS
ySY+JBALV1cYh1Oo8u0j1zLf7Kj7OwBCUm7TXBQNqeliqEjTHG2L4XQYp0pb
XxkbyRbopZFLwrhjwAF88JGCTNwaFHFUSlefYoUclM8n56qKJC3GBNRpv8wm
2/6phjQRFudduli3afWFiBZx/HErUgrUc3V1t6agPkISqaNlUTWaIk7ot5l8
PL4R2Kc0hL4u6De06zkFlbL2QAYOGIcuPoWq8sqIajcHdg2XkqDxRyazkUX5
kfBv2GCo+OELZzf+AlQHGln/lSo1W7oOYwCHDX1GUR/NmT4kUobq5Z4rDhFP
fVsybCyyZhmV/Sb7l1jZxdPn1BytCI8un5IcoCbF8YmsJGr9vBlNzzigF7jg
BMTxD2CnQQrMEaF0Lwqrp0U5PrtyoXHaYzp67FwjzJF8BLj7h6QsCjjyG3FB
HPWyXdQhuwwPblTCF7OLCKg80kUD7nA2qACNDJ1FHA6ZHpANu1Z+VLUrUR2H
Z86s0tb5iRBuQOnlvVXSyv+QAEL1AaU6UKG58lxxzx5ZRs/1PRVA/5+jw+Ls
e8sM307CnoiqwwhRMbsEilJUMFMBSuX0rNe8PnCo9Ivl6Hlf/tQJtdoFcNqj
44u2iOLxNVo+HAbcavHRzzmcazob4L9PkCBzM8QBq1c29EikAnnv2AudNwe9
JcXYrmidQ0AfhwywrdPGAPtq6HjikWb2j7i9BGFnbkaDGd4VA/CA+sB2EuIP
3frgi2zzRXU3MkFwRUc50sj7Pi0AOxyV7huigJ0bwIIgSg4XyFJ+2MgQr5/8
IzHD64D3Edz5wJYFaQ+XXsBHZa5EaDzafuL1ZomLBWcuq2I1cVyi3o/uFzU+
XznEWy2SGIujr6gd8/b3TbUKB5R6alrlVCbJFHvWptH+C7+8hrIP2y7TmEWM
Xg444bVzby72ZPN5Qje9dRY+ae5uOBNZ5140Dps3fYCN/LcbImoE/n9V916r
WCMXy9IfNCQFWXm56bBK5JdzMfssvqQwyKrg6cR/W7OR1W9QnWzTox5ky9tT
Oo6kZzX+jyotUC4ps7APr2gnpFO2I2XXZJvQcP8V+rbiu2POJshkv0urumyV
2LxtaoqcmfYElH7XSZr2RoND6Kf1zVX8u8Pdj5eEk1bED8mX0UvrCFU47Lou
0CRd4D55K54nAEsQBoyHbO8dM9+7f6EnRDw6PORPMqgc+TOAkVMJl+4zVR2k
WeK5dYs5jEOhXcFglOMWZ+pxYODGgOhZDsxkbBsP84ulxLx6H6dSIic7KVZm
qflswb3WVFUSSo3P/lg+o5Jpr5BtSjIK62EuHCYVQPQc3M0UPA4QlIHziUst
OLNCey1h9Mf+7ybi6sPoxX5UiOyGNPhSi30qKOLd2DsnO48EVUVfts9Hws2M
955f59siuZ6m1ogpIqb9fpp+896d1UqHPim+uzOaM03ucR92nwhzoB1nefwe
W5GvOsc7R+KmoKZavLYNrV5qDHCT116uPnm1lLUDf80Juye5u8qnvRGYR1Os
oN+6SqZSn4spw0HCXgj4gmHyiMoBfEQeifYR/Y9RWA9bubIDEM1/OQDg21bG
jjaF08t7cptnpJRbR8S8C7bECGdXz7yJpj8fqx80cZg7XY0SrHzf7QhRskrG
q1LzWsYlluuUG5Mlop5vrI/pG/uwDel/Cn/RYs1pe1nySdcsKRoUfr84j4Qe
XAA2RAvVt2hsbSKOdW9XneXwhLM00ihdbFCZQGi0h2oVTvdAu6JhL/cYVE4t
v3v3sMUbaf6gIwTznQYBVhh1vyJhw+w765lYfglHgl2PpG4WwW1BboaBKngi
ew9dnMXwSXb7qNt48WLosq99F1VqOV3LWoHMltgFL++zTiG1SNDta25JiEZ/
SETEpPyX/Tnhwg/Z2AiT/+rr5Y/N6YiLv4Vb0RjBKA+GaGQ6KnMQYdqudhGK
mIB/M6NiTgHofQnSkNWuAPh3c9vYwpa09wliyCf8E+FbtaI0s2MhnT9AVHJH
OMV16AuQF7pM8H36AivvB9rGkl17if7y23bQaU7BDAjxni11Vb529j6YbOJl
UGQRI3GbYnXn6QfJVYk5/nJoMzBgHs0n5+CcyJm8rO0qMI9qoAS2qbENWSmH
1ayjr8i7PnVfzLNfS1XeLqLwStG9g/uSnU1/6hXUoE+hUKP87sUkuSjR1XQW
rC9+uG65Nepp+KZR/+nEbHFqt8DXRA4AUw7SmfNLSwasrs6J3z/1TMYaWeg2
Tufqsp1xoAwSev2PYoPrdz/H4GHTQ6VAnaJ6mgja+mKG1jz4rxDVKtOF/zfd
IWxyh8Jcyp6dGJActAY8TcGoNrHnOSyuco8DdyIGo1V9uJ3xh5OiIwfDftOC
Y8N3pvwNQt0xu2aE3bKXAoPVcOWeBu1qtBrYFxbw/2croKcNQTawODlkQ185
eyVR7O0HzJlUV2vMU/bhuuV/Dsd9/gcMSCX32WbyWdeyZwSmzWoKBBAsxgeZ
i4pGeaxY80gz4xEquwq8Qwn+eKBmZtQm4OvHueDEw4KoWYEGkkbcvCj6HjoX
BUcr4pLwqQrZZQafQxtMKn/q+J4bKMdxmp1rhRuiDI36MD15jiUsEGtWbQt4
rQDL5JC93aDPTqtpA3OA1ojXYxtL3jECM5/YGrRMfKPY35n7eKBcu7xoa5j6
U3NxPaDcvKeVLMYz1abLhYdFCZNNrPMMGJkouYKbAzt/ExpOCfyxsuBb9rQy
oIk9lbr70wLXoNMP3Gc4DpBZIFyPbgEwS78tNlLfyh3WAhkMlYMq1xzBS5My
kGx9sd/G4PRD8LOzCn7lh+lJujDv7pbMbjUTQSDOQEGMr9SyWYa8AsC2y1Bf
Q/V/95Ze9DYXHTlg6QmCbnSL+M8dn6DHlxwT/wkwUAdO/8jHphRGG/Mf77Dg
RgMtEp1ugpvY01cR7Uui09SZ4aryjlAdmTGdz8bQOKUcRO/U1STETKbVG8Vf
boej+DSgNBdcgSZil5J4tyLpkdanYf8c9SqmXqTJM6JqZ9PTIsBirJZTYmmB
v5HgZWFFNrfdYmhJ9NhdioLo02gT3n1CkW9wnloroisXU3jQE4q8VWCKbFbI
v02jyZh8qMJaGbAweJ6z2y9ay+Si/lBBK3Tmz70UV4FsAlh6QuhXVctE2Gxb
WteRBChd9ULfRe5Xj1EXREgx/oifQ5PqfX00Ty/guwiDunei/VqZD2vGYQIE
yCtpibr8HKLdHNu/rWcrxcXCeSH+kX6Vd6FdAr7IFIM/piLYjlJZXTEdxxp8
vTqZRr/SEzHSPMbwvUZrO4PpHrGAzB5o1RzLI0eSQy1gX52VGFZrOxe6gg0K
00T63HVrMovptEFK9ijMHxzFA5MYDqnbRQjFQ2DMbTCkn1GKvWXZpwG5nS8L
cYo2R/9Yg7C1Yf2x3mKLwHtRkE+6Rpm7x1Yfp9wid2t3NfpDYCPJlDsASbt2
/grAB3IqRWZ3nZ+aofrTgZWfCEoibHocQ2PgWK0q3E9iSqfZzVSav31RJoo/
NBdE5bj3wIqCvKEjU7FiUX2F91Ii+dBb4oLYDBICb5CEuIc5UsWukosyoZia
ihK0FKJUdLzRyeGOHcCx5jAxXHrnoNrnjuSqCj4UZ7tTdP5GjAWNMOarJhat
0UKP6N0ZHKzM+A0ymFhg+PqxH4XYt9jyYhkVJTSDd8oI8FWTVsCnX09xvX8o
gOwtbtzEXRqe82OgY6pPdaLg/B7zZr9KAScpxLCGaR5MHX05wtqmEWwGLNfi
wfVVttN5NhSs9JhuXtbSfzrSGpLljS++P+9OvYMNh5HNg2BWQFLzuKOjTl/t
toNb3FN+aeR7GannOQsj37JE6gdsS0fEN6h0UIsTK0uq83cP3qVPuUWPlAsC
hlv6se7R0/5FMQH+zljsIZJd+iS9jMy4JuNXS88bnHE0w9/xztFDXLmKFf87
mazSFwJU3KxLkL4uyL0MMXGr56lghqmPgvh8Hp2gs0oyS2PZCvke0JfeWFGx
rQljYX/ulwNdcP9Z4H3PrXFYngfgyBhITMI37hJnVYuXc6OSXFj5RiikRqqa
nXy8yW3RnG3lBazqdbfCUrtXtk/dQOeVMQ71BEo3b+mIM3SNms99lKM+x/Pr
Kp750EQllyWiKCrscL3kjzQRq32+a3vDTHsOQsQEdYVyr0ZfZwOfj3bfCl9u
8gJhgV1/G0z++g8wMQ4hv2dlp/6SmP51HCdu+XmJQC3qLBDUSZbhewakPwhf
YSgqng7DIdqv771Yl+mL62+miOsE7Qy879IHASvC7RFecG3zcbngmtI4x+zo
1dzPzY2z7x04e64zVMn7GgDFPFCfZLou1cLWh4n4ytSuGnLAownxE6zOxBvd
RZG5jKxmcuVyikqtHCmDx9dce2HBnhjzSzK/CijREAXnYmbBKTckp5aA36zq
fjKW6dfkOT2INnQWAvQWGHNSaqVW+yV3ZVCuoNEMBP1Jrti1hHxYvbJap2RF
tsG+DkZcMVu6W96bh2vvk8vuL7K1q0DckGoxXOOdTCMxduI19tTXWVfTDOW9
pNhZngJLwAnEU16PMQQ7Ix0Ii72b2meETA2lRtGQ1ksDYb+Wbjp2vUQBqfO5
Nsiyo7Oq78uN+6Q8t/BFHjZrLsHVgr3Z2cZPfylZiDNrl1RvA3kzH9ByWxlJ
i1Dm53S4+Xl5EtN9qoqzjUPwdqRBJbi09cLowcERpPGzm7RSTz6luZDhy0iZ
kzNt8oJ7DNmO0VWvRE5StnzCfhKCKyWjtNoEHn4Hc/fIyEIT8zoQW/l7VKGF
WmkSuX9/zQyD+gjEJg/9I/vbwbEJVM5SYbJCpFfPgAvL14ANyJmrUhE1N1Oc
kdIIAGsAWmA4eLt3qKDuSyToc5HQWzDoHurzi6oTNfOLOhxdT98hOAgX33gQ
5ixIRHshI3gTozGN+u2UEVYRDl3d7IAEQKLNP0MuQcgkLArqY+wWNMITz0az
ebY5ujPCZ2/t8Y2s+5WQapqTdmW4SWHVhrTbVkQ1IXobpwswkvfZRarC27t0
AqO7lSf/3mwGydh4jY/s8hR2LrqS5PSpwyhFVcxg0rLkbq3H4TiyorrTxIQc
maRiaH1Ty2CdvBdSYQ8SfehUO3khnasL+zsQA6xqgcOLnHPthNv++P4RTCxD
hc98T1puzruZlMn43c47rHbsGYiYS/UuerQipL4uGC7W6IgFvp4mgyPLbnkP
zYkXeeKS3W5L61ACWGbvDqtSswvjOXp71W2+1Gu65LYMaTiM+ZFztYBks63l
rUlShJ70Qm4oRX454SpzsNlztAGkt36vAKeH6khL2Oq+gGGxlIgzf+J2/GSc
96D5mSHDqqTYSei6B8W+ehTf6OhhNrqQZx2HjOo0b+P3wUoiPQDdB2ss2+6K
YJ4dmvkirUnPcCGkCwxBo7JJGe16/QlpZFZPRbNgxyKvWypwtSqf7VKungUG
amzJGypOXup4zJstb08oeJX3Z94eHQPDP18qk3afCBEqOf6q6hR5G6xC4UFL
UfO0YnwYfK3Mg3hPh9CO35DV1Jf9oIwSioUTdBD/tVO6x2Brp9+tctUERH8j
0j4zcUi/L5ijYF2VMAmPb56qZqYWdCMrPXkE3/TSan8Bf6dSw7YWa8usg2sq
bez8e9QOfcbV/Ohr2bzo4LGVCR5HqRcS8/+u7+wUHCJk7c9lhA44IseGJLdv
65cbJlde/Gi7M+sY9uDK+TQNNSGeYyUMSlM39dlT2ssB4qqy6ndmoGHgH2t3
QY26GEV8yQy5UjlTal7Sdq8OQ0VGh+2xnOCJ+3rk/qXYuOj3ljmVRXO96fDJ
PCRUbZA6TFFMCsHJUIruz/A+WUv+OdKzzagRAkspM5Ww+ukp8NYA5o+lS/eb
+MI+5JZ0v3kPGQgOfLbr77iPm/DUI98oF1CaPxT5AobJbnU5LTupqmn1PsSF
JyHO2nXd4Ur3Zh3wnl5NH9Sj4GIR9ltK0RJIl3u0Yswct/i5cnSopF7kUovJ
XkmbNF41wHSxRjiLGpdnn+ljz+NFGYz3WtEIhaXNjSa27Nst5vBRgk2oPoWn
9xLJDp09iuNDQuzRBw+V7H0yuMS5Hgi110OHdulszb/q/67iv6I4qtDRgjJ5
aqf10iPejieJQieDaNfkwZm6tydBdFoHo+udFeXCaNVmUJxOc3J9jTtqeNxq
V4ZRHAA0etFSnOPf3Ip0zqhQo1JOPLZXgX3DzIaVsJbCsandjMecHU1N2g+R
w3je2DZIGDveYjxsL4Bu4UQNrEOYb+heHD2U2zBk349QWb2jcOcKXE1IMQiN
MYBQ5t+g6GXYo0aGHZDIiqcGCM2tj1u0MKjaOpLiO17TAVxw2vAxFKt2Zpqz
jR7BCUrarkW/IGSEdWA9cAUJntByigUuPIhptxNsUghi+3VMBWmhS9vuDPGU
HYjtdCbqHcaa2B4FRSuW90QvynB6cAeNChH2tzKDm2iT1ZgZkc2cs0OLVX0h
VpYnepe0Tv4TnIMZqSjJtwMS6ZH2O3ePzEHSoE6obohfLuAIOg44otvDJDe8
kfnLCekvyrrkt2hPt6yAEgMfmtd2IxMwQ7xQf3thr7E5dlv6Of26UOZ0tegS
gqxjv4JasNwow4gOH99Y+k0w2X4jFzkNt+C9F72yxsJQmOeBK3JtVDUNFP8x
oVtQxw2PgWQRbXdDd7MOIXNBGUQHw4HrAdsPcSjvK+yG/LFSwko1qx8v4DaR
vMmaoPQZyt6lYDDUC4pH360+Nm9BfLyVsLxb+kFogCJK0PMSq7xnsMhV1M51
dOEaeBo2G5+RrUmY3W6nkX2StLMUNBXzG+ns69LWoC7ck6Gb+4CU0SQAoKYn
rezvqut+ZIrtUidKdAGj2q5rWXni7Ss6TwkGq9+bJzqqOUtg6y/mdHqjUwfy
r+pVTSm/r5+8phnkWr03gV3rvEFKQkjMkh5hjJa1EHDbtoxG8lMzYsKMti7V
UTB3b4n4e8GyUjdbJId+AkOHgMum4oFqoPyvyXU/YAXhjiBNDV78GTuIVjva
TF6kutjAhvApwEOEjwvEz7/SYa1M9UIZpUOWZUybt19gUZySIhqPriYgDEY3
lE644qW3Br4RtonJufM2HSRaeV8EvR/3jw6FqsIu1tSbA8wRkW4n0GUp8mjq
S6mZ/Gf9JOsxzojXxnpZEE3umNdTFcygs07QGMYybgwNNEpqqAhJmpduyqO2
RAU9OtQRBthuJBaBHjYHrkYrLpu3UUBsJUpQsAB/FfJwnM/aaARlv/pZeVAN
XZdTvrSvPwBI076xBI3O+lm+5ak7KqbEtPKI+9ik9ymjzBWghLTlI/rQO8gM
9bjePKF4VP5S/NweyehDumBB7Q+YkUuILJTzFgdHa2ZEFKlYTrkyDsUurcAz
GqQUP2JoR1yANMVmtTZCoXVL6IIRKJkMULah0SIOt4MgiA3GAwOMteyhAP8y
pCeiumzSStvWvAuL/Dt70eG6rG+UPQkK2kzI8vKyW3wsua8ovkC0CvLHAs9M
jCH3Kj++l+h/Z5BzLfOQM6Ew0GICIphDaBaNp1eVwkRNaNFp059GwjpDCwIh
PAPmkY4u/5WtfEhJ1NJFiL6XpgMGEQ7UTlY7mCd1XYZqFI0xnZ5BWyKnzHNk
P/a1UuDf4vK57ff4V8GTq83DxxMVhmEF0Xj1y/ZsQOGxOGXI/f26iNw/Y0gH
ys4kiWpZ01Rozzm/QaOuIoAVlrnh3+9U9K11GS5pdfDr3xhNf+doHUTdZHqR
q4AzGo2nVgjFiWDSieSRcwhyKliFzlEmrMngsTk7gBzQ7FSbmMaabHPGrNqs
/D41fspU9KTJ3ouBexdIuyJA2SYtvzwTYXgjOcx4jTSdNNcMs/ly2FYKbwXI
/9iQdLQp3iGzk9Wr6J9yehHNw8SBynB8h+7YPhhwLiS/oExVT3JYP7AVBKoh
EyPbQeC2qKgl9pOEPArjpwBUpp+Lege/3fiJePtnGzu4Yq+eHmtYIkmrnAfO
mQCosprSHEEj8DjVcts1prnmnPacRxIjNnKUTvYbvBSn6GRoua4VvTE2J7C/
omwrwM9p69uh4yd9J40T5VXkY/H3el1sLYJtHF4xSBSZ9h/cKtLSmRwHWPHr
aE9p9PLjdAnHmLD937RNo9SdvdibCQSVaqmj5IXLfBMfod/e2oPTx1wtGYab
/zoKrHt663N1fDrYUVH2RHsE7C2/Li5MVZWb8xAti6gvfsp821a5S23ymyHi
WuydUAsJrISwMBB18eWiyEHrnl/b4V8+SMmirlV3/lLyPCCCG0RshgUfTYeh
V1FGxKARQ46pGRGdPFT0+gL/Da5u3AIUTjfFIM1IJONw2yatpgOpo7bWKHkz
1C4kHyB9Kq49ty5MX4FDq0OWMcv1O42nMsAdx1uhImKaI4bCvFYT2FyGK02m
oGMi/mmbfx6ryqSuwDGUUD7QDB1rPqSbaket9q0pMINhR4rG/I/51VE8QyZK
xuhb0XyYYNf5KPYzc8mzB8D5YmqPcqfIYKBePhL3p55Q0kpBNpa8JLcB0xZy
7+cEXELraCd2ytNU1FwpjKb254rk6ubBA3enLkNY4w4VhSBUHM1HZ699t4L2
tm6GHwgpXSCtH3FGqOyIDrc9U5BqoeHz29YJDxKxoneHChgEiGbKNDcwDkP2
fr1YlHIWMHkZ3yrHJKTrLs4hkqj9GJ1Pzn1SmsKDPZXoRrZxbfgr9qOVR3q1
xYMBBK/xWVTO5XOXUQap1wkT8+s4KPuQcAiG8wqUfZLN9PggLbU7S9gmkE1r
KNTFncJFhs7JhpDeVcYTKkAbpvRo6FMoBbzCiGhbrlWPlIee6NeBcT+IRG2O
st/Pmgd14mDAsz5Hj7dExGrk6f6aGmh/MFUbg4iR/nIghtznJH3UjWP9dwyi
KxswSpCjwe285cnAENcnH9DdO1CxcxrWnUjxtu/eUVFSjre+kITYiQ+E9YdT
tgzfqiiRTXzfuwv+7YfMlhnLJaDXd0Qcu1pNrpbILhgltgxNioEbdZIHD3/f
xcVqIgcmlQpY1AIpS0MBfOCQO0ZlcLmuQk74CyRbSnsdUXf9k7XIf6l3CFmR
1XDcsrDkzBM3xuhJWbIClYK/mrfnmHjhBTAKnoUQLGhEcZTIkGw3JOsQ+L1V
HMcpxpbo9X7zT+kiPJYAMzzqV4fnxvMmBbRyl9JwBVN6xTiQboIbrNuvuOx7
5RBDvWiUPnoBPDQxmyQT5SgH+IqlOSID5JA4ERlAhYbrk2dhLKsXGR56/lHA
5MSh8DnSM2day1tmA57eGXk3MMwvSzRLAlS84wstO6F9UxAoJt/BSlq+qZOP
8LL2qwtYx1D7A740KXKO28orABRRqVO/UnazFCe4+aJQ1TY1d3K9eEbpyr3l
dH2yYFei6rdFAlhMPbbmKklsqCBRL3lfluahGgB/6/e1rOrgyeUMSRK7TN6U
oQNEexN/ti3vZD1aYA+uZOMjHfIdPfLO/RdNWkpHzZ6VlMaeyxeBY+vkXgOE
6Xuuq22IOJj1jB+qXFwOZ5FDf4qSgvj9qp5Vpuk380TtiKONKS62laoW9ocj
bK66e2VfRGHcaS01BGgMqd3IMwG6mlkdQyNyfTinrfUztjRvHx6e9Thnwv7s
f3aTNRIUG1Yzqh4KDBpUKjvvQx+Re/ais3oU8OYTufcSpE1B4yq5F5Igz+U7
P7epvpv+2Cx6VrDhOG+YdFTE2eo8XrKErbVwQAn6qCDW1I/76arvdG2vhvq+
YRVqPjcmgCmmTGrREzcgXpH+mzvsoJe5Z0Z6FHLHHW/aaDaS9irGPup5y5ry
GhcsjUisFDBmMuTZmCUM3TW0irZ6dGqDhrNHuNbujmrpMrAl5ykq/xFzMxFd
IYcmmVskqWE41WpSSQx+JSIi6W3Ix6MnFFf6861BQkJ8Cok/AxrbT2Kenfvg
Y/y0VEl1KCBShIHL9Xk/5ApRBUci+xKcjyAEKR8MyOIDYVr/6weYsUju8O5+
PAUHCKEXdeBZfotBCHkKI1YKQbi0dFf+Y7vKUBtOfJnG300EXPM+xeyFfY7a
SHFUCWKRcKHC2CCJSkXQO3zY46CeICYhIzRnlvnsUwQDuumR8QFF4WjqcvSR
4jeOjQBA60Eq7T11CyGQekbIZmIEgtINzEJMhj+brlnCgl3cPnVxJiAGXucZ
IPWQVmlrUMO4DMXS8nWq2wyPDHr67wYheI+nrlsDv62QptwFzT3o7VL9BWiJ
DyuVpYI8YrwgBFpiqjE8L6hQcKJJjAFKcwYZKizeR7r3VPIRcj+W23B5kbDY
oDZ5wOe6VeYWpfi/+UGeueqxJbV/xNFUmv+llEmyxTg9tFdIrzbL2nZ0gAIY
qPYFXjecF7YcLY9r9vvtaeAV/PMqYVyyWNbDsxr7IxOvg8hxQX/rWmeQHKO8
ydofaTxq/rGO298EGM85DDTXWi+RSB/mzILwD+APNFAJ3qEQWW0DJZqy4K1t
MZXlIDPbhinjhfrD/cl0Rj8RsdAfDYQALDabsr4crxLmxhbCEUzjVNf5ii5k
2iQEbpi7rbV7mVGXwPj0jNsSfOry2vjudYKvYugBNxoOLE+d0InbAdFeWIKY
4/zQ7WIR3iv9fzemDSwsoz0Zc+O9S1E601dydEcBpV1xWZ+XBukYm9yzIaDp
aEJu0ylMUgolqyQgpiGwQqfJLkwKmp6TKFYhky2Oz5jOwxAoYCngfdzo4smS
zQ4AhZmi1HL2GrfQUMnpAGGbI7U9ELZDUSLOOWzjlO+WWUnaup1fJTkI1sGj
uuperI8BvsBS5MllhAT6J6OveXGhaPNJ6H6qoaQr2keb3Q6b8jY3z5k43L+C
Sk/q6Vc/B9j7V8VWZzSH6uW/QuuCfsF0GXc+4U8XBCqpdHaPuiu9rEreOVbN
c3ytZYm1S3TaFzH4LcnYOI9sK7kSL0dM6tHs/pZzbNCRo9R1dYNj4RleQPW3
wrGJHXDN3gfF/lqLCtKRnP7xl1p7lGTSSrjCe2u9T1W2dH8VuZOeEp1vpo1K
glMPpoXItZ5H3tNhnUsaI979c5dQ/7gjQkQ7a0/rjHx6UDi/M1EJqAdASou0
dmd5LxQ0VEX0H1DhURVL0vGG0qxdTEmAkLr4NGEppsEFVM9VHR0avq7L2G8P
x//SyxaoEx1Ys8cyHH5c+AydISiC9LlAVU5VJZ1aJwoh2b5Dl2NVTG37cN/0
jAvGqIyLtG1jQlxd1uDAOPX5QrkDH6GBrqg1RFKO7tb7IJsj0pnuiRW07kbo
uD6SCEN7tn45TC3Skfr40flKDvVSvwDQk8OTtMouw4WUd7W0R56xjxi26Vsr
cSiPUwVatVRkLeXzim/GhYf/PqRO5/Re0MOfWA8qhJaZY0Y0QxDxT3q+wSwi
Y3Cda+OezsYjaBl4gGM3PSf00MMc+R+y8ZvLfuT3QCBllCvUBgp+n/3FgF2V
qjefx7wHuAq9jTvtz9/MBgu0RxrZC7ICbj9GP3qvyzqzmktt5ZBYSBtBuu9L
QdtsGdLaCMNIQHvUKJINd0ie9yIOuBUBtszu+DIb4R0Uven+4qx3omjg74VS
Qn+oyI8lm9otYJAhbETEhNBBhmxROHhl4pludAd51QE86uECdX/VBSX5DjsQ
mk/e03LMcrPO6pCdD8DmZ7Ih2OcC4qAyl1LCq908ZfTqkWMLNJQHnu0lePx/
xGCiuxuvnutdwodPrU4Bj+Vi9hjxwyXb7sq5IFMdb14oLZHxTFLAg1MpAy/q
U6/2suXtlYzZ4cgW1T0chGery/9u6eSl6zipGgfX2R1nQVHuS2M64OEBCQ2+
kTF24r/gJbCZrjOvbGfDUO07vqxFYGgs8QulQcQ5iZcAp3xr3/a2vxTuc3t3
+TNDMqlmrvu4Qx3GPbvkcxH/DgV34GcT8XrVP/6tbaJXF2goo0HSIc/57Pg4
tj1uPT2X0KVv5mluJU4C7aHwVxH8XE8Z9Gv/q6msA5NJzejljejlWsnyHuz+
5aNoTVCApSvDqMgjz/XXLkeSbQaZOdpsP2Y/SVIF9RaT9hGP0z41I3RJzFGm
K5ZVKHfD9zEsbmsLPAS/ectyK79+ZbNv+LfBSDo98oZn80bfhtWGs4AS54DF
6aOebf/ZhXFbV/jOcTdmAC2MLanswjVd+6/lpgXag9vD0VaX/yvGyATKSyNe
TizmitcIYg3MWEebIlfGYsGv3lc1Ty4ez5vuZP8j/uAHA/RO6E1QjxgRbhVB
tChYwFK/RynYxRWY4vxMAjh5fbppKwiEkhhPMFB9YSBPkvXQxnUCIpglSjwY
rTaPV2+BkIDbgL9lWdJepuOPvpuGUcsnyb3EDfOsAyjrWVUqxhp/nYXIRNRX
BYiYwqxDgUBHXEzfQvsKq64xXdk4/Wd3PIidfgp+lXP5nlHjY0SA4f57zrOy
07mUOPXWQZYl4sJ3YokY9CuHBM1i3u7gmW4vAoH5uCeMmoFDYYOK8p+jc+f9
PfOG4DuP5tNOWJRGGxa8N5uf8te3vWrgn0XAJy1QP7CE7UGidI5ntS9FHb3R
T4eIq3qn7QYVq2ynPWGyjo7AARC4yKae+sB/HWFNFBQWw9C5TppccANOA4pQ
CMUvxXFFBg9Ie9876eYa6t46fK7y7FS0hH+u8GiHB22uTyv4G6Q6F0BPQhav
iDfip3fUlnhNrswpQwynv44/kPmOckk4R7LkvauGh1pWJVIOOJD101n6Wfka
xuJBLABSXegC1AnWVn5foD1n2CAbGRuNXBBmCKEpjV22T9GtvYH72JtI+qQo
yFc72nLaaG94ghYtpTuzrIsmZ6ZDa0fZtggOsYIicFj/583Mf2/Ebu4z5E4G
jXgjqkjWyEIm+DYgfaoHgyGv4eXwBEf6GahgYrLsXr7HP30RxGKhD/TP++2/
uiWPEiOYzxGwFZe8eKz6lwETe4SlkfD3uRWnvUzUKB4m3iGW92gJXyrgoj/D
h+W1Up5OAUaPCcm9msCz+WnT/T5vHm2DrMWnnSYIDz7DXaPWlIlqbvtegtu9
24qA0lWLoWNjy8jYTJdLJrr2NSEK3TIcpp9RVaSsU037CP5JJogidPhMyau/
VJNaZhkFf+ebUzZ8kBarXuNXSrYLpGM9vJX/umUwP+E5Nvx0xxyhQOZLIeXd
sTZtIJQ4/TDQIIp8bNryok2hfalOyQtRDQ8AJ/Q94OCKw7hrPAwOJzteIxyI
QKPHWBRpupdwT9TbvjcKTCRSMBjuDS8ElwGV+OYXJmHwt2uZFycGXmbLgngv
NfFaB2O1mpub088ODdLOGaegPDtThoTLC4rZwXGyC85lhHL4Ja3zNPqKCOz8
Hhm3fpl0awNw8RLYFL51Yg/YNDIfEwDfMQyZ9B0pLZWBSFew4QRl014LgS7n
riV2tCJ55+bM+DHkqwwNosGNPeF5Jb1KC/0j+TcF8u2kI/w6eHJ35CnKjnj6
Xti4G0xEawdhBqlufMhWX0DBXOV9bgFhAU7pkTlzv5tlk8KHBLelkByyJyye
bm9muVo62yvkwZdyoEycrueQ52DgKiYxbUgjfSFtwQYCPT4Cj4p0rwy3WRgO
fk/qcYGZuBxwf5+tV3cEiD64v9YIe04OCQwS8BanK/rVhy4zm3Nxmxd5F3XJ
I+u9/GItnwdEsUn8vS505080j0qV+2WVBJjCeDygeqL3DTWnFn2cVtUTs9D6
2lPGJsETcKTLfhc46MTx/cC9hcgNGgNneDJAjMG2CSu6fx3uuUL2mqfsmpsv
7D+FpmHaG7Ma8WacUJPluKFf2DPm3qFvgcnR0/SGM+7ETFbcr45j6C5RyYXT
EVepj8HDenBYwwTi0Q7kE6jZOXOxOPhYeB/m8VwjKpdRz0bSAEhzaBY5wClL
187qoLBB2IMp20Xg/MTTn4WRRu8nrIL9N2rnOk5MpjTlpmvta6yD7Hjy8h9E
K7krb0l7VO/wCP3803zycb3zk5AbFULbtuVpxCmDCl9z6euL/ygUXchGBc5l
r83gTJG7Ne1f0qPl10zX7Q8I+yuKb1csWe7APhZcuzDBQ53vVShswnvPVAC0
bow0CLmOxRTRC6O2hZArbs2koKG7NbEPy01c0ACzVID/QP+KPY9DghfIVrBw
mHjpva88aFpzt2vAI+D+HLh/oq3GQ3Pl4cgnTSbAzuAPrbzNDV5XNdsGCXk3
ua7/N6ClI4y4a3o27UOFomPyo6bKP6T/4stFi52vQi2M7/RDUV8uO7b+guoD
eRDtigxeXRD2klJallbJWPl3oRD82AA5tb4IG+UxKbJ3kC1dLE6ot4xJh4MD
uQEc2BvFUbtEtz5XZjeZeXIAasAE8O6iQ9/byqQInF+dq0peeMSzEPeCG9wW
lKQttrqUC4F4k5eamUKWAUROmODVYrxRPVRewAnQytwdG6Bc7o6V8FEUJAY9
1k4Kdy6aW/E+PDApPn+FUvlHGb0Bqlh3f97jWz53RFngeuk0BnIOlR/9SARF
Aj/5GH6HZu6Iws7Glf2d+yD+LaTm5iGIAiR5dOuCeR2qFuVt2OqdYaI5OgH/
tS3FiDUuQ68OB7FSTgMj5mnzNWa0znZCpXwDWc1pJCxRwQGygZICATPoejtP
4MVbQOgdoB4SASJpixHc+yHW0WzoTimkCOT3IHxqfvM5WFUj2VHxAOXS5BzV
bEFvGJ9maTZR0XosJG1fpd5+wOLVgmKAb+DhpnfL12GU+85yGs1uZkrjBq9H
fWfHxNye0IID9MEOVfEcK9WrU+3EqJNU9UzZwCNi3I6AbLrsX5AfCr/wy9+L
AbT+1bGNMINq8GljUJB/upXQKosNpeMiZJqvFTw+/j3gpJL9q6sV41ofX70J
Pz2cYXdyKaxORqWQhCnz946OZ9zY7IHpkxUk08hXtIl9VobSnrmxfNXGiGuS
KlpSUzt7eAxwg6ef5/arjYg3akS+wyhu1ejPLKSMX05EC/DJUzORHJDsGeKp
dm/8zPGtOaL1nj49Xir9hZXaCVHOMpk/PvSaD2Day4eYcDyV20GptExm02Ln
+RSePwRI3nEoi3bFmSjhYGavk7kwFxvIgTaMSb+A/TROGczTWUqZ26taYBJ+
6J7NF60ZyD3BmB2IRzqVPQdUyp+YzvAq/9WTmNHR72+iEy/IoSZHIGO8C+lj
X9o5tj1Pd2nDp0yKjWTeir7vUYjQCNwj+Q69nJ9DkLxu1FAJU9MR0CHzI4dS
xNcqvRtJl7Pf9EpB2wNUhUDyj50CTVFDP+EDhsXBovJ80LS5oY415xBlmHr8
dImlf6cZwYSU4ps+X1iV5IBsRk5VlVegq34QtTpIPlPNqNvZSXoV+93lb2JX
ImKorseiWNf7VfQgPo/ybP5keYfLfeG5HOqQby/6UowqZ8epxpSEarHfMbt2
kw8mCcRrPTS6J/L7FA51ZwuklMzZn9kyKYilShE8SnTrx6Ryr8A02BbrFhDF
3fWenFexwSfgWhNFGdSBNlaDJ1+qpHI/rR8HZ2tcsWvj9KOd622N8IBQ4HHf
b2XUQrS5xycaTJjrVlm+lrsJLBdjvkCg5YzO/b/6iF04PQJyFhoPUO/LoNUF
7CBn3p80Dmdvq/PNG1uehk8BQC+SiyFUOMZ4TqRfpp2733ZAdbxTlc3tIiRG
8YydcvMwL7gMPRQLwwSQORTd+CLLU+vXCTCNIWwODW6VfYxAqkhCWXlV0JHt
izITDeTjz+RbFuKmugV7lnTIje20pC4x3u2UeOS3tU6hNMoPGNIukxLjWixY
e0gRtZOcQfotc6y9qF3p/0iENa4F2Bh1WhFdfqCVFRSdCpOJO7koLglF1CsW
I9eBR3YbYXUcPZ13350PjI/lCayuQun8lE5qWF/pav5ji8LWFg+ubPwPSfRc
EZphpw2n+p0W9O1KrNWvlxenqN1GSyzEU7Y0wbmjTxxRBvLNxTNIxVx8Gvhn
LqsjrhnIAM+8T5xxrl9/yWi/fNvY1Cj6rB9uKRpUus07BBWRkWcOpxGmXbxb
/rDzMVZGwnuUSNL9S44MvuvXaNywq1ncWaiVmHZTAIL9l24iRHa6vGQHBR0l
XXHlIejuFztk1PPuFcrqrev4NqcUiR4m90+z3O7zS/tJWg/CPa0kFG751Emt
nqr4rppDwWoWyoLj3BEtxTjA+JQMcOC1moyiPgEorwl3yCtBkWFn9aqJrgmn
KQIM590+DMmBFkQO16bwDGaDP8Y5hPl7lchoK0jKdxg5NGLMk7sWH1B4GZMV
Ey3iOK+L3A5ELrA7cRy1oI9yHlLbualaOsXgT4yhgHO3KSKAK/yf6jOiM7c8
et7lmDcyXI63IQD0iTdH7N+bt6WO7OPH8HiPcOlQK+PPu4Zkgrn5y1ChhPMi
9Wf05tY8cYUHI5Q2J2Xf1lad0YzO/hkRzl1zzpctRsxXupBhuml0XQQEoSDB
xp5s0iyRoj9/i7GIJ9PzkgeRf0n3/hbp/svFxN10MLlNlVMd/ZtJLt9u2ao1
nlRkms+0+fntY4EmamgNJN/zTITxZ3pg/cfBekIgjSMoUVYDPVuscoVDPDip
RKodbe57TsClHWu9OYsmUyF6R2Snuthvvq3sq0OnLjhdthXw1L7MjcyPOx/M
XOfaNTTz5mMU3LOXTiP2VrxVVW3VzJUwpsneLtXlojcU+SHRPXgyjEcCjFoX
kLv6y9GcWMz3kYza2qEqc1c+PaEJgNwBpX6icoY+1+XuOcu9E5/V9gFyz68o
JZmjG9gutHIPzIamwTxWWKi1uUvPxynxKzU/PjPpiSVCzHguqwm60nHgJXPB
Wi/5GNMystyb+gig4DCD71vXRqu/T5f07JH8+XOjSOhgyMnrLW46F/DRO7AX
2BAn/cWU+PMi6CEBO/X7JtY0twHQeaheQ7R5q3ctaFH46d7+XG0hgtXoCC9p
UDpoxke8W5oXG9JSLEWYXyhFAx3izLoM8jJ9aXKLZOAthmkYG/XpF8Fz5dBD
rpPmEpd+AWE/CVd11qUc4t/bizxVjIC3foaJO3Gpqv7rhm3oifnjPc3ieIQ8
n0jDlHROWQBiPCJ63xyuLJGSoEN+AVjOcJEKKOHmlwmiUaBaR1QBs6SMSdo4
wyIsNMwSyeMbg1Vwq0VHeeoaIkDSUYKh5binS4mr5+8K2p8uZnj8FByMxhAu
E9IH8cEGb5uxNvY0iNoO/Ui4GJdhukqcWiT75LiI4rtvX5nThyD8u6ytNA4n
NsJcbMeNR3UdY7G9dWhAhJLFr4oQZw6rFf7pF2dLAnTm02w5IK1bVg5Wm0Ro
nHEudQb/fFb8g+c9LLoH6LA385HwVJ3cC1JKR3Livb1Yzibi5L6a7rNS+IwG
WIl0vO3FV+65rWAYPf7Nw8KokdA/nAaF1Y+QwcvNo1QH6rTmvvBkR/fq9Tjp
N3IDxFyvcC+PJdBqVuDvBRnr+0HZJ4JpHv9YSbbmaBdU72boJk2Ya/HCf9jZ
G9LsiJhh/sXbkltv5V5I3Siefbga3UQ7A6NmQ+MFvLYLBRGPW7vsDfxglnES
fXeFLNyx/ErrOvGT2k0S4UZQd080aZLBJO/4PhJIatUMx5xVvtfXP64+uk7i
BEMqE5oRlV7o4+PU2QfAfeh7BGS9JVBGVKVSQxnqL6kNeVjU9nOJiPi1opAE
1UYjoXnDzLdYQv2/6giJdzuYf2tLD/OU8utd0thPvnFz0sqOlWEnoaqaX2M6
Lb9k9avomoBXOIAZ6GVlFK/dvDJbGVyfqfqJ2kruR9mynQlXjBfScaCt3B4H
sYq/Tx5GmWhUrX5dWWEtfpgyDgK0DkNv+bB8VJTfgiiy5fsKUXhKFrJFsYop
LIdJmKJPCDFtLZ74PWEspKfV8//C6ZUx1ymZou0hiIBXr1PyMp+/IBsUKIi9
A2GMOjQ6cWJHqPgPSCAduMR0xfb+RBqjN7rSXHg/9xr7N7cdfcgY2TP20gTX
gv2lxO5tLtpb3Swsw2hx4C3tx2eSa8HLAChZ0usDvpFdNH64Z/zapPSYvcvC
lBjUhJDc1LJTa1dlNG01+QgIp/Aj8J61/xVBAxcWQoA3hHq3H/YTHP8D69vz
ygovlecYTiwBVNNnbkwVIaDSD0cz2RY0h9TAXPxr2gMhs/+GXpk2vQaPs/ua
fbFyn6dN07Heoq1rZZ+KQJyzOKABngXTATOTpS2irYKLfcDqodkTHtiaAHph
akbDkmcWrBwsWTWOlzvlNtsBAUVKniunhWW/rljE6Y3GIjF7ipvgql3lmZ4n
loNKDiTS+V13P/GSP4fjAYDMdSZ+7pO/KJwV+4ndUL8osq2YUqwqHJZsethD
wKatnVnTtE/3s9nLLsqouNbyY0XalZty2SgL8of2InrSRTsaIL7nMgQ036uN
aGbjlLd4hqNUgyTnV+fsgn/STQIl/yMBxbsVn2ciixJO0kHo+AVmlq7GI800
7TA+gQSSnVhLGW9e57AnwMIrqUsfNARLnGAFb05SYkLUmuhvCUDzNKKDB7bZ
6UVD8kTOi6IFi/NPUYxGde8o0fNB4rl5vRvFCsy7mGW4hAWM1Sqe+17e+I4N
SyASndUTKdSljNk6lx+yAWIi9Wg1s4QJz73DP1fdaDaUyZdhmXNcO/zkLEHq
MejYN4kSPYzEd3q/z0j4yRscOMiUs34B4j68IIDrOnjGU6/EhAWr3FhyAntj
pNXa6QldglR5cOyGXCGlkeToDYlqOUAwXCyvlr9hSv7ahj8gg9WFYr9glXgv
SwC01TvYwDoRKv2jBtc/X1R9Cnhfw+a2a3fT81NnpK+KE1h363RdRYVHh6fx
GR/mz4boWn+To4SC4dEJMSo0rNZ6DFeYDFy/8q/Wp1tp1731dEbtVF1dvqGR
HgfaC3P0TEKnYPPF2cMLslU9DVo9zp4LP2DAHes458lxs1kP0h4UneC84xYa
WbMApoLFSsbZA3qFNoC62EoM/Ovh0hb48IX9LOlz9UsV1FhI+rc4rZasmzpS
rF4KYpQMyx5/rEneGz1WgAo570E9SR7d3FX4bUKZSsFJZwpIeioLkWvCb8fR
WCyC6B0FEZszpLFwZEBo1Egr/TKSw3/rh9CV5+8A/C86oD2VDdxXcACXm5QR
D1x3bbf+7TcAz6LpWF8EqDAstaUHowSk0N0+q/Nb3Uze/mBsW7rpMhiXLx0o
7JeDblii9uz6In7P0p47FbqFU0rIvIRz4/APVV1gU6t3dGWOZg38OY4ueRRX
KCFDNh8uQCIo3Ru3nvZphV/E3C1wfrB2Ozx1w5ql7u0tm7wWJsqdhW+WJtR2
SrvzHqY+i6Ay5wkC7idk6CfqPy+ZNyDx5txTjpYrzt15pqc0LNrAjdCbDHzF
jeUN2mAPWppEMjp6Tmj/cmxKub2N6QL+bh4VHrh5BpFyAit8YU7klPei4CoV
/Sy66BtybYy125RYePKwvyLWlobAhGpDjbhnswXVp/RqrLVmHpi9QxUs7EVM
KmL8wLC4kD/dj3xjmYbibb0nMajZ1O6L+CPU/1JccbcUBABRfI1wUxmTXrtT
xcUQo3zNMYyZuo36VQn3VKnq7dg7NVCRQA/R/cc/eK17fdYqbQeY0dKNl+1S
zfaDn64KNI54yJPwJJ6QWGK+DiL2RGaz1kjNT214GmNxMzK/krXXsX12EOY3
1oLo6ZZq8kSU65S5jzvjC8s1jTj7wXXzFn+3Giqx99TIs29HxAOffXUWv/yX
jusSuQAWClZtQIRQTWdNhlBAcvklYAw2s7Dqv3RDikJAtm2IWwP23Vs/1sVz
1YLfeqw5JyEX8WLZESNJJhvxTtnY+hXrvbjQ9p34TX72Sl92lxFwnCwy69PA
/9GVwl1S7EmmuE14PTAbmQV4E8ixVMOAScVJ35Y3X1bhkn9gfli14dtrXKUZ
R4TtqmDJji7FjrW+eylfpVQO14YjVpVuKndiNkbpVrfMdOJUUHXck7jdJLow
vPO0h2uMQgTUb+ZRFZg/xCg7uoJ9bddsk7Btc/MOY+dNG+EiBoKIicOt5gDA
vvVl5NwuXEDoYSriXAUipdCmn8hpYwrnOWdFS4WdIOGpN0zeWK743btvFUZ1
MPbN3e9jxf5OsplfTylX5qfrsu6dhVhsbmHlZTnhIY024P9YhfPT8o05QC7x
9aOoVkFew6LoiTE1cHalkgKYREh5Gb/lMtiIhav9423qHolLsH4YObHBZqOd
EnNhUOWQFreyuFjLTXCTjuVz7QeW24p/106dMG9EJsE8Als0yviEMavU6yy9
sqdrRJPOIId/i3Q8Hk0su4n/ZmZVwRPGSiO9RC7jhyu8icVs6K7pGm9DwCqp
QFCMHhhwQUFlSD/x+0DoGZePJ5fGUuD+ALuuU+tZyBS6RgNWTi6SevRzC8gL
9JW09gN7qTpp7s/0l5FjPUcDLrk81qgml0q5QSosQohBnTYpoLqOoyeVNege
oP5H3s98HUHgf0RmUrT9H1AEQik7bjunIXhevBrk1TYd0qA7OKzNIl78XufE
opRGxlnKIrp9PD32jVIUnZFEDpVTg/lS4/5PI3Ty+XY0zRNlnz7wxhakTarL
Lhc0MIevPAcqIfwinciExjtYH7lErCpLp2GR32n6Z+rV/ndcjIeHOnpicUoe
BMfejV+AL749FV87BxlbyqWyekUkv4sYDZrleI08IgYC+9j9144ELnTaz2US
Hwge432G0XoWMmYp4w3ZIDMKT1DJ0zgsCr74IB0y6F2XlI4lh+VivxG5zcWH
s8rVGP/gZ6NIaw8o5HAGLLRdLqCE8mJLsA+2g5rGXzkWMXv6wJKqGjx8YU4+
mkJJLGQiKMlr2Uzx0Z3VUaQNS2gvrgg+h7bCKtL/XNN8KwmFWTd9vLNfvq+x
YndeL28ysHTqmtXG8cqiNKKU6tPrc7EBrSH4yk6MMIOmdmFaGpKm79oBkRvb
Z83iQhtqbA5NmJWIUkug3EfikBtc18o7Lz2GHIK0Io4Cavt2AcV0+FYR+2D9
85BM3728RKupLCeADWjdszWGk+Nb8w2V08w1xCFG+SMTu7YTJQPGW0MlmWdO
wx3mTmtRz0Tnq9z6L7R6fEIavU/AdH0ReWNk3E5B17bzRQli7BnJQkm3wHQE
cADcye45hDECwcJICm6HeSLlAMZFfEPA373eTh93OycHyQAEIKHq/IhfB4Rt
GvTSNu8DHglQxDJzLq46Vb6X8tjEB66c6iZBaf0YO3P+n0G60wCEmOlxTovF
5WDSe1PFx8hGhZS2s/p+vG9hvHm+xmjh2Hxz4IjZWgwz97xHk6tM1wtCOlo6
gs9ABLdjINDQbIjXba4acImqGv+gNkTSm055qsthdlPp7qIRGkOCWN3khXCw
5C7GJRGSaGSBr3IcZt8MO9feXuHKXcL9XGPsbhombyOJXjETdwxXkJE1TSmd
9ajqxvzST4MPmTwp51ovowZvQhcW4x1jNOBDgeZMoawQ6RAxNOJakTDoYk9T
mhtBB2wpyFpZvMmRmAD37cVRFkkkJ5CQyZvqSvcmY2VZ25jY2i3VIoUzjhVd
G5dPiRwyHuFuRrHyWreN6JuegrVq4eFLrRDwbL2L0DFktGet07qmohvm2Fvi
IBwcMsVqRdQej9L2lcBPuWbjqMwvcveIsaXZ+copraiIJ7zKnuIPuu6e5X83
UFMCQ3PiDSGkE2s8PBYQY6nn2ceJ/wP4dvuGdBU+y++qks2c9BevYzyS/xz4
aksHCnm8MT1VUGA96hcGrsxIIQ1F/Roy6wa3SxOCXFHjz0QFwBGJXCllCVAb
RAXJRrOG+skHVLB/l2S8e9I0XnB99pBb1WFtdIfXgWXvWxZ3BtYul2FzpyG6
hS/zlIYbzXfEBIN4R5xMmFxQjs/Ow9svc+avheTvAI09Hwqlix5rQwu5a+rr
0s2Q1z2FnGy5R/cTO9ts0k7s20wI78piRugvq1A6Quz/nhKciF9BCoxTyXp7
yPtEklXFAmL6Us5wNecbHvMu87Ma7zvmyvS8Ct1LQ8mOah+aUw0zI3I+GLzN
NntLKCepoCVG9kw5ygEqWDfKfPCexiEFMEle6xYkbuVhmmBLnXyqOnbPQg8D
8jW9oSrlwO1M0VrVK8tzSRQJDNJA/OsruUvntgq/Pmq72iFYfoNpnhWfWJ7K
GqgfC15FuLe0685xd0XyrYOqvmYF8LuaFtTaWMDpVGA65xl3QGZUx58KwXT+
bvB78toJABDAbY7/MDVTdvk6qNE/AlbGviRatcAPjiMzg0Q2YVK01ugcbWFa
QGBJ7+Jm/K3YHG9PnD+etNXNY+HtRu6hTcJiytwbvJ7dz8mYKBnR2gXzs9xs
TSkuocnQDs1HxYor9kDU5u3kQLUsgnydw0TFI0QSIMkSRxbZTxumTrzDYRlQ
hg1iSNi6YM5boQWABXgvWprXzKtiTtNxS2ApSbgG4Bi/gvYIyW8aYJutivLg
3TTV46iJARJnOI7HjwHo6i+428iwuTYVu78THyc/uZWt0oT63CWccPieC8Mi
dr1Jmx64zVcpWOHDaUoZufKNMF9iQ68vV/z93xt6+uxmSQvBCVy3kba1Cxok
zYVPeLnCDZCAJiODi5LgrSg8XxQtjX1y4F7K9v21FOJeSKkS74ZGKcMSfL4M
G3fw28nvgR9wrEmE55XwrbSMV8+AzFh6WH5O0bOBIRrelzj0ypOZCPAOhWBw
qIRkO3oM2023RNRKAJ/2ee7bzvKZ+dyh4czeLJRjBZYmgY1jAbY+2PJnRwDu
CWT4hcbl+mWb5JLfqazs6onb76KrD0fC8pMDijNbu5CZIUSe75PMKJJSUMIm
WJmdrZoHC1ZLIX93z9EgM1H6rFb3mOiGJ4wrXMtS/v3ZOVIv9ncdMF/l7zGc
+B6i0cotrb63xSOLDazmoZBMrZKNd3f1SCy8pJuhP435q6RileEnUGZCZxL8
06bo5QkehFJ6Hgw3cNSDad5Sdl91zXKmIu0BrSEjQBv1GBfpz97/uttaY7yF
59OtXBv+JHW6HCmbZVZDFJANgfUD/7/Ot8fixXBgGWrGP7Lqrqb2sgbOSYnB
+jqk6Ug9JRfWUENfpHJXjM4EfaaP8xX2/jDYb4Ci87QyiS2EF8wh7KX6K13P
zkweVq/WHxYJw2mAAFqYYEEDKrjKBIKuE9npR5xbWY4deHu8lEb/TOOemVMR
4tYCiI/h7F1qaJG58YNVzXAunyAFTfEkJdnIIt3grQxRPgbd8Rd3zPqUhKj/
ILg6mHvh86CRvGeRRqHetZ+d/A+qtOSAKnyy/KJv8+ltVjy7fYkTUKVtYcS+
K2xefpTh1SrD7NpHWZ4ygZhSy35Lb6RxdnYSWsJ668Fhb/dTPMr3jKOb/ShH
Fy9K7cVkQO66RfIdc7fDDeU91s5HflboN14Uyfowl2/IYlG8zPfOG5Yv8RsA
nVHEgiugiuPgqEK9zS1UBOP3kjYXlZ6y2WdWW51yQA/9c1xcrkDdhwozIBP9
UIvzIc+AZXe84lXhfhJSZ/qhbifdbAH2S6bYBOyVar1Z6+Ll8eYuSzurVMn1
/jwCTdhszI9PoprkKtIV3eyMnIhYUBKyGD+03dUsT/v8I2uwp3D5EFVhb+pz
P5gaqdzXqqVYzqKdSrgXP1COIBkcP3xKv/Yy0+BGm8QgJQoq3KiHSDOt738/
hvJ5iFbQ2F7yhc82f+KUJ/HARGJyJ7aBVKJ7PIZKixRn5zTKVgoLb0R5FE6m
GFL94+ZUibpRo9aD/LXPxAF/pEftJt1yQ5SkbX61ftwFOZGk28dzPgkhmkmM
oEkdZndb25qg0FYku3WgIkVs9aUdpyIcQox1RfZe6Vei41qQwN1NepdEmorZ
cD1hwlHJVekX7xXHLv+GxehY5lzmiwbUKEKszF9awyu5GhmgwSa9WSrdoZ32
HKhSzuCopi7MZvSak6d96US1EsXOxYHedwohXuLiTNbdlZnzkMz8HLmQ8ZUi
ciL8W1jAhwhkA6tA+gjwoURnVEDmGBtM0HzRuB5eWLhFxvpyUfkBPmIwLNOI
Fz35zYlLVIGdQpWn3kG/YqWjM9anjNmUJUiirqZQ5i1k1HwQx7IDL359J0DR
2tIdzY7yGKJAXBhs6DPbwX5JgQIISBn28M+LGL+nIgzFb+L/YqqEuC3HMhCt
tIoZBryFQcaB7e/Wftvlxl4x/UrsB/YDv8LQzMyUP4puDjOK5c0JbcZXO8OJ
Dez4pQGzvDjX4Td7IfCwRKqiTUhYfONfHZ7kIlCRqBwDv5XrG2uiNBIX1tRF
34klQ873blIJrHsAibqOCfMpvZsB2vGSf1GRmlx0ZlkFJf5myhHwgVo30fjg
27C5t0T0k17dPlT5+rUL5QN3VGLN4d+M64i0OkbokjAXm/1dOKNdlWQ6h3Hb
R01K+QGXbiu8Goms1LzA3diPpyR3trQrmY2sH9N2OSsJlC8b5ClXKW6TuVR9
VMVr+GV6uzialFC9NllHkIRPEF6RkP700zel4K9/5VDbQ+8ME29XXxMBxb/6
uuunSXA8obZJncLGfz4tVCrLSGYc+0tszt6lBlLUKb1Q+XM88kz9Zx39lp7C
Ldxksh/Y8YAAmHHMyKawCMeRWH0MdIbmHjaTkQrBuS+G5CEPMqy8YZS7cwiy
Bb6r3YhyYymLlyhE1DajoNP3DtfpOxS6KzQOfwW2KYI+MWALC7fge3fkl/VI
7RkKbhk+61qo8QpEqeeKSqPP1fAfgLJx7pNBtjsY7IIcwuM6dTbdWzLL2fzF
yUYKwh1aH5Q6iCPsPIQQ/iq2qhQI7hhcVX4QJiWhYSH+YPrkDtTcpCDi9Puh
TM64RS/7oQOgGzrGQY8aRyDtySFLoYfFjQjV5YrmCoyb9B1fmnXsAbsegr4n
LKCkLTSplLWWVDtxle14vsKNVXmTMiRvD3Zr6MN7IZ7QNc9v4WXAkPFm7R8u
x0z+KNm6o7xg2XdIUs9MIsbuuERwj0IH8VfWuPchtsyiVQx3iGC7CAJWfhPg
+Yu89cAE8oyidLT5dDZPdDmBlIj2I3BtEKV5TSy0XfMHndVEWQ2a/4R/VFpR
GpukVpNPaMkqYiWgfg3/jSegcZsa9+CRUckmEMebLVVaY0CMd9Kpf3gCNQ83
cmNm5QRL6x3Ql7V9oIR62O7aqZ/7zJ9FNu8iBGe0zuZAjlpxKh/zRC1YJJZj
mNHB0iD3aytHEEWPBb7h0IDOm6IY8lI7fMu7CdZPmAXtqolGjVseaA9Ig4uo
hLDePXVZbW14ggH6hCPj8dgueSRNV+t3TQKxtnBVZYNBgZ2x8CAz9SUu0gQ5
YhIcuB/uNRg5tDK3pgXJtJbh6zObDZ7o0M3BBERZ1zDH+ME9tPhzEvEyBsC4
MI/o5KzNdB/rxG+M37qMnT7oAuAGbMPngLpAYAgyEvhZMnRATErjLhdm3QbK
u6hmm6SZyUW/34qC0y2Yvrg9i7q3H/cW+KHN3qJCqDzkYRxUYf7QrsvqX95w
mG4K/TD0sv4VcKz+UHZO07Ji9qDrpYh6Fs0IHw7wLkSkxVtbdOnBOCuPxexF
BY7MJ7L2qiSeTiCX+Kdi14pKLzhe9q77lyqxYntAQzp0tebv8XBAYmnykWyN
iBSS2I2hQim5gleAs8xtWhJIx6KdYo+E6sCRvkw34/IO3bMEEjIwBJ5qndCX
OrSlH2udneDR8sV0idH+K4htDA7YJDUJGz1sJ64oUjFZjDB68v1dYG34UdfH
pJ4UmERGJJMP5uBXw6YX2W1yDkpcUPm3ma//rveh+VhRSgDW30RRIPdpZ6tq
i6jP1FlhUP9X7Olw+Du5Kx3O4ATc1c2sjmrZpwSxg1zbIZV+s3t7vV/DflAT
Dux9Zk8QmGnd9/U1JApOeOxTNXbrMtUaDT9OeLBM6if64PGfgQS3EQiyum6o
H4LpW/wBgvajJKQGa2UmgxbugarblbShvzQJXujKnDJtTN6yiVlHIkc3PlxG
WLCqOEkBF3hp9Rhd4bNgiz89narY2h7Llc8NL+OqP8O3JeMEEsa03L8cHbe4
EGuRARVDwlsm018qQoqui430tyv3AHhN86UkLHsUKhqvVzUIadg1SQiO8oNH
0S+xMRjMqDCWGexwSjycOqKNNEpu/8mgY33JFZZKDBtlHTzgkqVRzNEyKiJT
H92afJZIVWCFBdjEMCOxWfupT4d4qGecs5QtOVYFSENszSOJUJIRn7fHixoc
ZbcBMf7RMt6HTod+xJQoqwTGHs2Sim65rMDzf0i21yF5tHgZkI1GBGprd6OC
u5EvyJZhHKtT2g9+6PWEnkROZ6Jti0OsBAs+w6QK2+zMPysCYvfHRYzs/Slg
twLYpVL4Tcoa0YUKkLqs9HpAMwbNRnjg3tFzNZeychlOhZNA2wAZCXDu95Js
KiEe9h6QKeC5a+ycgqLeMtBfyhV0LZJXuHnQrbL/x2I4wByjHrZCvPJyZztl
rc7d+ko4ldVkB5FP+eg6gLfG87RltZtW7IIKfhNbhHMtg1i71gq2tLGHs6wc
deykooJyMNqStCciZgAbp2vgtVBVLCQ5FLkIaiZC52uezgups4EhWEQqsolE
xqF6A4uCUmNTAhMMd/VkZwfJlHobNBnKxW4043krxiI/SPJBSoyZ1pKetVqh
szqjXUDkLGvsNjZE/Jm0gl6gTMfNlOpjpoFPVK+A58c/YF43zh1/G1vIJWTp
YLEwt2Q2nIQ77pPNiORlsRx9uIaX37pkAVrZOnf4woC1kcnTBeUmQiTKG+o+
j/ebRQwwwxT7EIvIoyS/1qyQJcT3qVVZiCLQJFAr5jC6n2vBqPoxXzHLp4U1
cu2J/+vlp1SXNxQhuBGYabsVfx1ojn9Sw2WLCcfNCPjAqwj5qYUAn99FJBk6
e/2x+Y9sPUDp5sfwc3GIta8brduSK7PZp/Tn3y6J+Ve2bbgnimMjjgue/RNm
pNxfv6J8bUKP8NkbBOCPJvGLgI55SRJeHs8E+wag68SXhAk+S0OBzljPxmoC
/72KhoSlfSvUIQCpxrKVSHroY44R+MalhDlcR8UZHijN0mODQkB0txLmikPx
uHDm4ia1azkhlThCydyQC8avJmoB4mDQQRUvMR2NslE7hCBDA4C5UfhAcK5h
3V8hLFYYm0LqiNPbigVNuVTy5GTd+EjP9PUYHGTfoSNJuTFgAZ3mlkcCC8Q1
3KgrGvcoAat3j79X6tY5luopEXf423fhmL1kkm0P03zDJpAR5o7ce9EeITbF
FWLV3epGQ2LZbjpA4MXXnKYB7KPmB3N+mSdo64KYoToxsf5f3+vklaGdGdbh
5imjoqHtYUoNSCwNPNNnKaPA3AHNN80pSx3NXf/Kd0r/WLwj9BYpU3CBIWJH
2o9XZegCsz8GNMg/XYv+p/Z0ZSSkFtE6J2UOVTCEvlpro8NHfHsjrYLyOl5v
VTXAT0njCrJlfnT//PHRUKKkmV6fy7aJPP4p7eI4yf+I0ubJ65i0VbNVHtyB
in6NciPqbaY4LUQbiWHOUenl8kB+u6ZHMbjSaNOMZXog80ew4Y8k77z7bgJe
Jtr/HrmngfVedqOhPrZyFUw1s/8DtamZktz2LloqFeZQX0ogQTnuWx+z3HfI
5UBbvPRqdK6if2QEXo/vjf9U91nvyUgjIuD3secztIgB0ekQ7wXLfGrmuEGz
54lgDQYYKqUjNbj5jEpKUCLjOArPmXCQrtRcAy+sfMz5rAdnLDHb34RZMR0R
hDU5qUUeKMJvAHjWHjyB344AMbDwZDyWOIKo91rF8t+PNBlhPJWdUjDVLIEI
ay/D7GmsjRT1lwgS7gG6isCa4dJpCQj/XWexYDfsGP+lBl44Ihnn7F2l6xoe
82ZgNyQzgJ9Jvhb83GF+6TgiS0NLk1n9hHwrrSGs0/nOjAUatHVp2TsX7w/F
sBBqNnaYdwnOCRnvblqrROxODIJrZqXrAFeEStihV+mRkWKiBWAT6qMAQ2Tw
sZFB4IvP/loghk46X5b/4DdBgfJlJCAIdBDQrkqy+y/b3o8wfE0TxUv0Hmew
efJsqXK5gITMcmiCfX/CrlPh+aiBFXvSQEjHtK1dZtc65LJxbQ5KYrq687V+
zQQ9MYbHAXOAk7SLjMmD10x23AGGiSc5Qz8AlixDie5ao3f+TWPOwjxWXCAx
baFH0yr3Rn93Z0ueRDOJDmTB5VesrTxSV/HFlYg3mcBepb1hxIJzi9+fKLZh
bBg7OzsFlU6tgXVaH4UlHiKiGyfrZIljAREnLgx3PhnL0QGsswx1CDSMDwGe
5jgB+7deZcheW+mwVCYvBDIWApbCGdB3FqVmKcSRRYyb5fyNselb+wi79ePl
KFLGJs4PK9CQK1MIxlxRQ9qK4S2+YQdsR+k8dp01lHXhRM+s5J091wkFdwwG
lPRkrmglYcE3H8eNnTrEqKYeIi7fJGPHi1XX3VUW8dyfWT+EV9Vq6UHme4VF
4Tife0cE6MksPBwKZQbt5xtNnRBHekvvEAQF7ZiW9Q9YH1sgPGJJ5IKJP0yc
NmwCk812eJy6bbxCpTAQsAAuAooonHjPMvSidtD83ckVch4MWIb7h4VlBaum
KIkbpV658kl6T1YvyMFu6073fcOYMeSRIgHO/18tYoKLxppsHqsOpN7h8ISU
AfYwWpqYkxdKVaBplaxijwfKpOFtSj8K+za0zBoUsENIfzoB0cHw1jVezEj/
qT/WTGyp4OrXNmL2gikuVf3xQFVh7LduzLwj4CkunCTKR97uIGFLoDd1Wh+f
4K38dSh67kbzFnF5Dntvgd3h3Tz/Z0JaykiIJUw9sd1T6pJGQdKlYx1wi6BF
6xwAcnp0CLL4gv3bKZkFQBFemwk5HIg8R1HPwoTwcA+J3MB2O9Fu9JN5KrJ+
gw1hbcJSeGeVQhAJ8Or5D4zRwk8tuVtKqg9nHABwlTZy52IuF5q32Vt3rKok
NDgnQjzN8vFzvHLqHXftD1/6+QNpM7KIyPc4bpaIcGPP+7x7MLi9+M/SGHrv
NOFxRiZBA5OclcpaD15ineI9wiLwxPAGoWY6tuy43Bl67j2JeNMUmdH9I/E9
1CuAfPgTddbGna89RJ0J4voNnvTjD++poIVna1fgWnWghOWKCxX/ZPqD8d5l
w2hJnoG/FMhJvnbqIfBAEssP8bz4kXVO5NJDW3wQ0KueQ8SJu7/lgRCe8D34
cXoJjTi2jchKkYG7RiuyFBnrqtPgHeODUMJJnkiBLrZosXEMoKnxQCpVSgLD
AD3X6Th4uhQYo2RfBPDqOxzGMEk66cMKebnkgOA1OPEz6ZaGTGbByAM8Y+9q
FUsHhf1F8WgVnPAfyWwRq+Gk1LwJdgMMZUnTq5r+y4SkDcmicEvy3vurBNVz
u/dUkW7rgoECV0obGNObKQDR6EAHocKft4xiSnUV50opA68N90KaUJgmzURG
syqp/sPm85jTRJi2UU/eG86sesAYrHfTHn5yzIODDfJ8llpo21BhF4DxoIhL
9IDtOrBdd/vVSQpCu0q9vR98z/aeZoXzXUQPT4UlOWA0GHEhX8Dvn4jZZdtm
xR4OO+fNZN3ylTOHYkO4jsaUhwdjQyrw7vtdg7l/KO0muunSO2cxX6iZozpk
yPjxOyRMsSggV/RBGBaydUn6hOaLmXsieb8CD5Woy/DTtJJ4pWr7TSZ57HxS
4inLYwRBW/Q/rHwIjjh/RvaTjOayMLW5K/lnwmBcMZR3l+18DOoiR1v4Uwp7
rOA9Q63qQCMBbeK/623y3+9ZhyjqcT/6a58hRtJdA7tax2WdVZtwJgppAHmW
vWeGkSJcN9rZSGuOqe3TFJLVwNBJm/St7vwu69xNbkZzg91YhQAMYml6zjVT
7rT/CFAMNVjWwoxSCfLwhgxuwhXkCXZrqXmoano+4uH4pPSKpqDt+nVHq/d2
CVwmYh/BlwqffFOHQEWgPXsAok/oP1vunYKr2qkHI2EvlpvGekSmvnk99J/m
12RZXvuv4e3UcgJOYaWLiovVj+qICs8CFX+CsEgKwfGJXR8c5oa3diVCAFBL
E2933PoFX2mtW/RBwswOkN6iHy9SFpUTz4SVwkh8boGKJpqgJhwcYA2kxHbB
3jQBm0A7LAO9Vs+QEqWmiQSpJJnm5c1pMm2UDFdTKJgQ2eHsPHLQK16j6bqL
8Pi/JHEb3lHvUFiBOA1CJtuoTI5Y63weeTS0ebmLiAxf5wvkvIpmXwvGHFny
qLGVofxH63fJvr0iwLCwlAqwFdCpkLcX8JuqqXdoXSqxpFZA2DpK5uhrYGQO
aV/J/595TUJA1NjyA/VlzlK4IBJlvlJe96NR0iFjgWN32gfgaEqQFEzxRNxY
8jZwEqZxllygvi/tcWkLBXVnV2iM6C5ad0Wb1b+UlaYAB8B4YA4KiW1/1q5l
SbZhu9JfR1xrGvCYVF7IrXTAA5f5+V0jBvV1gWzCY0QbmPMj1pttkM8BHog5
O7AEn+Iy6Aai7PznvOFuBZG/ocRMKVK+fXUIaJYrCXW2Ci4MRnXnQIFGgsUv
q3aGcOqwO1HdNqkkslSrZT8d1mE5+OxQORbheHruW/pVQ8/rVumUS9nnSMXW
OeZqBFav7uxd55ZcH8r6QPQW3jTq5KtQvX0zCzX7yllmg2iM7b5MasD8AUzy
AUW0q6AgehhY5Puo9mjKiT9kOsmXr1L1tV7tlVHMzk5rVxKS35O37EWy7lc+
O73c7pOglNVx7frpaNMmzM//VLXPZ3zm2akay4x+w/NGDLRQrsN7+OFC30kj
l6DceI4jGhRQb5AbUnH9acNVycup7B0zGZAQcXhbqk8zwpOM5wQoFolWmd8f
NcCK7284sWsGduLuNeKZ/qGIKUdQRbcIan2QEP4jRHAbBXf/TppYtyARMfcd
P90Yk/EWgayzszzZvDa/hIbOAcRQ9Zke3ewTKpQ7Ar3cFE8mCN5vaH5xrQ1H
RT7E60gnlG5fvmQo5mGt7x/lWRsGseVTUV8RsjW95F4rYdIYgOxBvv2aCBte
mmcKxKUgLlg3RAuXPQxEY7gYAsKeHX7M5BmSdYfOrgWBmHqPghTDVEW+YbIH
Te01sR9CB5quwG82CXSoCIfnAUK0DQA0GxMfU8FO3Q7r1ZLN18fU6apNKFho
zEAbWddoxV9C0gyBQwUxh1Sr+D+YaBniUwscb96tops02n3gre38OLLrv7SD
zlGMOm4JGWzL7jOoKUmBxGZ14f7dBX9LPw8R8b5meOeUqpj6PItl3Kal2+5i
TKC+D4qMDV7d/w54u6vYw5i9EyGDCTKIzm2Ru+LEYaT6MI7f4XiJpGMEe4kz
JjhoMQKvzFw5FF/ftwXalo7MEXrqhoCfqX6qtPL82c3EAnqXPvMIleq8Bax8
rboE0yGdh/HF6W7q1p/dLvN79iffwF5h/w0RY9sT68/wbzG4zd3jLlOywcAP
7J8POL2zfTuqFoCQhQoZhqkM8waqhRP1WaIAMCeBmQRS0pynAAkDgWqXwOg+
UhzWhKzDxeImuHdvqlpkpbXBgNzgQN4/CAzp2uaaF2fc7WM2JrOW0bmYDfSq
upIpxMIYJse7ITSSvI0VfmVUlajcHIsXuWOWPAFcpPtTzoIx0Ghqx3AZUeHO
+7p1wfFXL+3Kxks5VVvZSLhtwIHSqSRd+3HQtuHVRkv+qhBSbwzgU+rOEfwY
9IEeMT8xIYmhLEjwItroG5hyHT11BfNdHtKeeaN3g8yOh76Vcdwl6Jkzp83x
mUJ+uJ37T9Sb4kB0sUkxoz4y3H4jAWVK8zqbQ5BstaSn35Vu3K9wRnCSA5VI
K5ZpR+ubiId0DNm5Hoze7Mm8LwNU/NdSmT4TLhr6LFES+yNh4YuAj1Wmdep3
6tuol2dTnngqmY5Jn9z7PUH+l6Z/u669S4w3XWtdOkguYWyauJEV232qwwZg
Y+HJ1WmlHZJ7NVkNPf0SsFE34YlMgC0CKX9tGVDNZkfNFvkq0QkY6ExnTpVR
bKcFWRurk9csn+XRPTXFCAJ+Vl70YmMu/OsurtE9I2LlPZJ4NMYfQGbtdvpg
GmK3/0YKr1z9sQDo2DI7sAOrdNEK33paLIZ8IxE+xT10x3flDGUoa3BVz2W8
gJj9weLXho5LvAGTS/lQZKc0mo4UdfdIbYuqGAALnIKZS4fiVahSE9n3+zS6
5d3unVDFi8bJitFSEKVXfX2k/Qf41/o/oWC14IINOzB4yEs4Ir81YTJZ5Cwo
qio1lss08J9mzS9gFtRgGaAZTd1ckbXrSxWRC6mZWefHvIPeXwlpndoLNy/c
fomTET+excI8lNC7v3espFXxCYEdJ9FbRimvxl8kT7gdgqpPv/rITHA6NMCU
ZTSOJPeCUne66C3rSueJerzyFDLUEHExLsRTMh+rt6o9jQ6EMRMQyAQ/H/KF
0kGWqyA7zwz5oXxElDTG1xp1ljvOSHsTViAE1J1ZWM/9Vcfbtl4vOaL+55kJ
YvUnYCWJh0a/3pWTP774yQQKRhpHx95ZHH6OThtB16hzdO3OwwoRi5QGacs6
niUX89OpADS1hEKjp14bNWNvb9UEYz7nLj72JWn7BZ9+wLeNVw5Hiu3EMizY
Mtu2p8hyDNrPuzkO2TGzZhgLXxqtKEuEly527zRgNRpJ5b/Y/LB2UmuhfUzZ
xwRjB1+XN5x18GV1QLOA+Cp0zB8FWJ/m4/5pdy9hBEMX0C/U1DH7CcoRpuQU
wp/+AtIHyZp8StqWT5m+Kx9jI7TD7SiyzxZHNjiTj6EJWb3RuG9D/lmHyEvM
/YbJJdQe95JoPymi9au1Q2SPFbERt7canr4+aPA9YMx4WE+g2hGfk1B8cVX3
vPHS+hPG83Ez6Lt4in2MgVaL1eKQnld7GlbdMgZ9HWDORhUBtwme7YsSic5m
U8wMMqQeX9j5Ayjssxat/CF4CZpF10SCryH7PkMiSPbqos7Da+DzoLYiYRvE
R8faK6N/ZAfQd0/ge/nSxziGkdzP0og27bjGho/ICY3P1P2j8kHsin6v1yZZ
JGCf3l/qQU3uzAAEU5YP03TautYje+NFqNnr3ybuvosrviAt+7mPbZyBXoAS
DKJ0/EV5Zs7rq8Fc3kMk5UsgM046Pi+FgOzGH4bHLbknHg4jchqCblcjeprg
6RXksb/aEYBv0GVfv11IjwrFnT3n0MuPvUISdbBPgsMwpq6wwJa15EM2mz5h
2DWGXuWi2IMNpfkEAgpSm0AscJhfMbq2YhIQGfBRIzHXhdGGa5Kjp31kv23F
FBfVmMipBA3v3pamAt8ua+MLSK9i8NCll2Df7f3zLrnNcZNew+o4hvqy37bG
E+gGy+h9PvdFNnOGHLAyFExN+PslxE9jJJGlOpeF13wIx/mezkPv8xCYMFra
nDnHv6DWCCo1uzOsD+0Q+V63MYzbNT3p8P4tHfqTkIPEBs4niaIaMimT/Tx2
/+jHLCx91pad3XPFQiO8xq+sQEyvM6AAe8a0GXXrVmGSsNc7CFVDb1TfcOwt
WJbwKctrmXDZ4vGtMS2pYkPPA0Zn8J9uhEuaEOIn1ZP2gkSBaFpkziySekS/
pZ7hIVUv9NyS+FsuI5jGzlbgPVJ3bmTpEDjoIhlGmmPTxhMhtEl2MZRMl00V
J1/buhpUxWDO325kfDf0WxvpZmxOiv1foGWZVeGHaDMuJBRm/6TsmibsVSQg
ONEFck0KFlIkOWNFAWHJ3CRuYSULjgR/VpXPuaOSZbnGp0+rtIUCbj8RYp/l
xTNQe9vLRungKrlzuquLNa0har+9m8TFo2v/HuPLow8gM4j9ZgTtnBKYsYfl
lutD7emmLBtkX2kC6EA2F53mz5sYNxnwj5SAzM1sDmOV72+lSYQ85y+e1f/Y
yORWx6Jm4oweITQNAdf8JvP0UPjr8rL8/IQ/ZCaYqJPtQmJid2KcqP+ddP1Y
D5v39ITwemeQ3ifF2WlC4iuwFkASp/mOWJ++Z56U3FOYcfgN7mEOVW8OQU0Q
5csogCpt3RSA8ad2iYcJmzoTYwKdVrwvNaKVMzNYfJv7WjzX35RYTOnUPSKd
vyxpA964+ujTgUlAWvpVr/hraSaR1EBof9EVYJJsRaSXwbuvKRlUl2svND0z
5DoYp5Eiz+KGD0/gY+mO+ho1nHVOFptVoATWpYyokf6oaOBUcQO+VQyeA643
toYpbhfCvY/LROU6SfYivzKqMvT1R0XF2YZ0DdO22V/+YCMKdPfM7d4+AJyp
o7Af0erDaEA5Bb5jQJsWSdZHElDoOjcnr6OrX088oY0CIs/s0ATg6KWDipMC
PM+0FJtlv1odYzMyIveW4xQ99EKjQblDKm9eYTCbDouti+vyRoWNm7XgUVi9
fjGNHhi88Mr7wptRcM++CvPjSwY55I6hpLkYExvGs55QOsyWWjgAjZBNORRb
HAlVCyPMX5bwCrxwRT084OlAZESSfEYXNSmptLBNNjOrhLU1VSaMtK5M6XwM
lkldC3pl+bmeSbjJOFRC4DUv7Er4tMe7LZkZskJz1trE6fWDxECAlhkG9zdY
66dp6teTMVlFaumkU/PkyV/a+j3dF97fCK92t62oe3MTInxCoZY/ftQwGw0c
boVvZ5lZJ8lAidJFMFxWXvUq4FW8mIxg3pTDGG0xNFG4nDQJdA77eXh9FI2i
jZelr8q5dV/cEGCkHQ4wfA30BBZQ0gVvX96ilGYtabJQnfo1Ld+YoUWsbGgm
j9IbQrmSYuutXX6NNMLOloX+tGrNLiG7p3qYfLym+Hgj/hjvjBLxQfBq0Yf5
cWpWIDqehSZp2KLb+jthDORF6g7bGVhlCdsdkXkbZYO+l6cbSxXEOKrhyX9T
ptmX3rfiV0secOESZO0ZYgxI6b42L2ZAtl7LPGsY3eK4XHOO2Q0SJLYqCSdL
6FZBMIm0D3TGc+/sHkeGXGTDBzkRqAggkDwUeaRc9MKuLXJ4rxvOIVtV52cM
9KzGWWULWpe23wm+CUXsm2R1mvq7kYt2riNgz0d/OjwXiNzwsqwbH4jgglXC
PfFXWYRJ+HBZpIdsiIp9teNBqBcl3pu1wdoIuaeel7VwpS4Gnl1J9sjaOZOM
XOiveEgGV2KwbDXezETWye/JVJcm3baPlhPWvVsPViT9HU2LfsYYRZ6u7sN/
TUQoCYxFDBguMlC2/kjfSOJfadk04sMomBxsKSn1AhLRbJ51A/jzKarBdNH4
5RZFOmkgfORMfSb/djlI4+DghLeggyzMMbchmgAS7n16hWV6uYWIEzaFzCyu
Ty0UaZQ6781W9J4wkcJnc9eNJ6nZZpmzFGu/3r1HzWXGZSrMD0eqoulP28nJ
ZVTT/z/czKBIMt4tBm4duPONnooLkwW2SmRA0fSSnk/wlRRzV6cK6po7ibHZ
c67PNqnRiPZJYGpIoDOA59Y9A8vE4U9w2eV5xcGLL8vp5H3jHLiZam3FlKYJ
/rif1Q8khe0vzXVTfD/+ofgr8aD81dToS3pk5ZEBy9kkOsZ/pJ+Saycxki15
NgEmbbsKwGIUkj0V/Owe8JaFSchWgsPNVFSiDZGQCw2aGkrfiCJgSmyUhPX4
o4u3odBMnxYPSyKiiJPbwHu0p7acMuhYvc4kcglskyuo2KydR4WrMfxz5xZi
bybq2ARTy+gmt6R5y1C6xdJj6OIK6eYeE/OvJxxRHm9Ed57ijBup7umfHxSl
xQT6LDYtr6RrYxP41b2T104/OWNGCqVVGP9EOTtsg6I6QgdnLbwu9wsWft9u
OOn/g2bUHPBpGUmAadM4sSz3F3hsZwX4as1zIrkY5X+UWxqriy1/GVUZo8Lf
o/CY1G4dMXmPzdb9IHIOc95uMQyvXR78Xrx042zANYQaR0Qss1n8J3ymVWov
FjW46V2oNNyi4uehTSVhoWi1bq/7JVyTAAY4ysvqQwEKAc8Dat92EJ0ZcjRy
Fp2oN7neH0Lq5ikjLIItKOKIlvZqVQ+iNNP08WhhfVduXefq08pvCS11FT4P
PZABt4ZXb5PubWpKUGlDXOQSCrFvBwSrXWAOpiMw7g4F1v9C2MP8aP0ORPBy
uYn3a6v9Fy7z5VF9DH3tCpZktydrH56o0//Yo8A5RIA9VY0y6AIn7olInLWJ
8AvZ2tc3O6xYcmKfpE22/0Z+aKq3CzRuCFMAivPxVmU4hD1PvGpVLr5D8Vy0
PRr2ZrMwHudIoEUogmLIZC0pGqbrz+82gkIw0HpBVn3EsWO10KIncnSjiSqK
v7o+4Wk5Vs1xZSoLdSADQIroHLfncPJ1n8pnOgvU7owMVqzTDtDbZUfUp+w/
WKJXTJ7W7/JvI+E3V/fQGs96VKwMb75GVVmKVc0mOiZmNEtvhplTh4ieClMi
lZdTWHcXZyIWFLHWd0Ju0c5Ccaf9xc2SC1kWSQgEJihHIKBD+0AlX6TG9Qyy
/iSrlXwZ7bSFjqEg79sb6jW0uXPIAR6z7KXr7NZzAos6YgTnHtK1TnnWCKbL
2QyEOSczZqYXK6g/M1WobNSheoCg6PATs4fWOW+RsZBw6jsm50WjxO7E7jrg
O7VOpq3uowTc4GpsLlJ9AKLT3PWq5zxpSagAXiEAx2WOJ7hYpiUygl8O7QBo
yM1pWQzNJAsfzwqBd28unbCn94KOSmwvOU+gtoPGIcJk2EeY9mxibHSVcszW
wOY1lWx2PqW78f/vYDBJ6ahCOOZEHZs2ga5OZ6W87ZP+7Bu3upuUIJye36Vv
yu4Mdui4W6GDtT0r3jqR6NzVHJF81e7U44LFWAjoBfpn8zhq5U0r+C0XJeUQ
7FWe3jQfYe//zBsddtpwcWzpJeZcSi3sSbiieYZPsIZJXOytGmhdeaYrTlSd
0MRZmx9DbGDYYuMmdYHpTj2pB9UW98lKNzOIsK3DxxV6fb8BsaALx3psZgHM
MaIUXvJgJEnln9NiokH7fkD7jpMpMVOMYFcIm5p6SmR5Ok6C2em13ZsCY5u/
vLwR2AnL1oUomBWj5Z9fYqehog00S4TXl+Ivwz9/cJRUJkgPimEcYwusQ9ZQ
VyC4kGjDSXBn0RbhGxi1QA3pSBYxmZdr7HsnjxWHNmD2yS6PdT49WqgeI431
xYa4jR8Q2JVXT65Z2JqDbCki7MZqHRuQ8X9S5xOOJNzce4d+e3ZC+bRHJBv9
IFnSKNW1gGmCWS69X/jRXu/cMh0pNS0EjzxpfaJQNFKSgMFsAXri6SO6ewsZ
gZaLyOuwmxTvwSxrqvoOOuBut8l9B11d02iz9z3IGsSL+QC52yEhp06PxaZr
DvqhQod2jVJW0MC91W3MnJ9AUqRaMU71RFZBFxBl+5agzGcCExkNXykvAnJj
JTW99fqXygZWLrZobe+N9tJIXPOdDrIN/ravOJt/1UiEBVmY+gV0eoLQvRbD
c51mzVZjCrVIce4Y/Wksa++u25wQqrAW94l8kXpoLRJdBsYYR+3ja1awM5cK
KTbtVBh7Z/1OLXNrr7q8f0zMUASKPoRu8re6blvNwhExIErkD58YrAraZvbp
/4ylBz5dQOIa1jrjLr6C6yDCYBE30M1sBPEliqNSaQCe+efSpZ/qSdvwjL7b
1gvusJmBrAQsoSq3fNzP4BOXIFdSIQwCOlgibGI6iGfl01Ln3BQI+aGs3xpg
v/mGF0XXIKyzLa1HaahuK1s0pdiZSp9jDcpUZY0bbl8XyqazUjBKdcYHLpx3
xfsExlNNyt9EYFtN7ibJarcliM7NoicW4cvC4/WO+VPPiwFON09qbpyNZWOo
AgBlTHQ0KP3JHP/fKhXP1l6OGBQ0WOEJR4/aepLGrpPt2EiJ4KvmFH2WCl80
/rFGMhD3dI9b0PsPsuixlcxavEHthA6oO9gLFetlWESKxsFUCk5mC+w1bBjA
nwLufo7AIuJy7JabHx4QDen+HIs07dY8sPVwJInVSkiRtBhYsIsndNDzyWDV
Lm+jbG6icAYLm1LHX6+h8ESMA54o1uHxm/I3JgHwGJOQ3ZAURQVdJVdMOCfI
wOTloC6WSahuesN67WxKUlvpmlz3YA72tul9RmxFAhKAr0kPkTU56glW7IIM
J9zhhfXyW1fXWRepmdfPQAg38ZzkUJ9xxOSSagKRK9P+qboKNKVTBBuCbqWS
jx4sKk+BXjrRJHfdDk3XPJTN9+BpTIT2wlU4Tq+O9OJ84Ar1HQHn4br4fMsu
5CVhrnRSYjOFAlQnDKM6sRm+qpF04cMQNGp1s2wQcGylAg+8+48eoLVXcEOI
sJ/ejQNzdpy9LOVD0irM7jW8Qah/PKQtOnvWFD7O2AgmV4erJy18JVJ4w+gd
GiHpQreg6JVW/1OfSvF+29pGFBp0b7xe6frVxJ7IZ+Z5/Wf1hVd7j+W5HQUY
8MuzZcakLC2ac4VAZlfLHmkUA0rwknBGgyEUACw0p6SgK1TppUjsQpa0nrZ0
Abpht4EiDPIhKgFB+ZFUzo0O7iFLz3yIGbuvYtW+gqwEzqn43sRIVrVfE+kg
YA1P8LMi1S+MHmSaENyYOTa2FxZfCmO19EERbACS/WXWbhWM0CI9oP/Ws7Fv
PNQVvCHnVS5JMHdeQ+/pc2ljPKfFRoLHPADYXD9bytHuQEY66TBoW7SkljfQ
t7+IwYnmdqwj9X1it7tRl0UDnahaMDuk9KHHZG49An5vj5I9TbCaAPweW+Y0
lkiAYJFuftAnqUIRkQljbWpRg5egeBavLuVkhL3OJ00YEQgHDbWNoix70OA2
qfMwypM3unOT5WkbGZ/mmKAl+Sy7O4JXNrtGbxar4LyKX13NFXlMLZhC1VBy
3y2B9G38hGfFcABnOdO3HI/B5xIPqfMbHbFZ3eOHTawsnsq5tngO1nTpjSQl
X7pKxQ5UpRt8WW5vVOz3xFTdFxApJDU9sB0IrshD9e6fpNko3AQb+pCAgjq/
iZ9I2IrLrArIe6hKmDReSqganakvs+OyzFYdLz5Bgh4O75g5aA7ofbn1/UWk
akUXBmuNCDQwCcDPIMOw4MGXsOtSOlcEl/qggogHkM91r/wWAmty5d1k7I2R
kJwnRYPvQzphYDf+GaLGCvLezktkr7OPzuTen3RLKBKitBmxu2S0wl96D+dp
OCAMH3jjG51Bmb+O2qPvbSvSBwf/AJvcqq8XtJAjxjFZvhiAyJax7b9dwbEg
brQrtQpZXglVrfb8AarzY6Z4IKWhiQaKUS0k+/RocHr+nsfTOpfthOFiElYR
BdJXujhxoZLDErMEwc0I7U66WVjHowutZ+ilsAESNej69CnGMTxqMHBux4rN
rotlUygukDh/t+aJjkqEBW8NJFcy3XRXJyaZK8G8/LYE3Up7xWjegY10tvJ8
IOc2HgUJRVFs3fGo0WGqY56L9YrW7sdvJtEB4sYkjUOR2RttC/F38CMV5w4i
oA9z1wljLtO5leyoFYyDIoQq1MaBv/i/DvaoE0bxbVTXT0UsGOz++UkF819q
EONXfv4Di3L1yL8mB2+XXEGMkS2GAXDGm75KhtCxIqLkCGwZJ1TCQgXLCd4F
zLQGlYoVdrrSV0SSzmn+AbUcgH/OvTJJ8aBstvNh7sCcvSSRtNtk8/LC3ubv
31AtygblscbiCV6LUrANQbJ2zC4gKVj9r2Z+XEmhcqhKWz0/8EDVYBZGhdB6
mPhb2ZxIKdS6vdKYvMXfnLLqKzBNCDQyZYEi4ZIpArDY1i4/aLFmTrYE6wFC
jLM4mWmZgq/oh7R7M8rSPk+e4xzB88+HSUD+bCQH8zuMrtYwDQdomoGgHZEk
GzqfousDROPIdKQ3GJ8tXiPRKqazq4Qf6dl1sySQ7rzeJZIriRSHznz9CgfY
IXbVFEKf5SVf+v0TrpLMwJJIcS7QsmXQ42URIyGwmlfiX3ItuYilU49QYxAK
ZNBc3AbDx0acY5jWvfUyngyOM28K8DXCdoZewWqFLCpgzqW172f+ht6BLlOy
zRO7P589VKTXcxStm4rsT12aCleMXxq/T8iYJbzUIFIj9wifz+Rf4ckmYnNg
uANuBrsCqQJJGHmqMrRzBY6z+GvukT/0V+a9EN77plPHut1I69STxVBQ0Ffa
DaY8AecAQbVcXzn/yvYmaYWBuG27rp+F/NcSimFnu9yR1aRNAkdX0Vughnfl
xzEKDIKqHV65+/quvqIqwnhHpin/X6dW3eRBF5jaWVZV6a3trakXKYR2XKMC
R7B3bmdK+j8P5lUnir8//0L0mNNakMDUIMBcg9kjlhvJjO74daqjPTipVXxu
8rdmMG1ukgBd1Z+wlLeL5dfZDN9uSy/LXed6GpxHfiZ1p9Hss+/GzDfNrfSs
+30p969THHuFu4QNWDeT1b2hVzPM1m5rzwBISCyCmx9sBIx30Yb0rZzE7Www
OxEr56Anp216GlONxyIo5SQv/0utjdSVrJ67EYx/hCI4C/RYgkQLLT6hoXRh
PkDB2rNZiA32b0g0HQLWTNBvOzZ3ME6ZvcGtsY4WrDdbYqfWInsG2sVG2+Gr
sr8pvwmeyI+cUXN/4G6fUvZrnzV7H5w9TPpuhSfZO9jdlgoEbUHYyENGJfOP
4igs1/OhEkJhPVtaXUqK09rtMVeBTnj3B1qirhNJtYDXJLMeKI9ZpKgnGEcU
OQ2qqoz8pT6Q9g8Rxxdo14HbJ7SeIYBYprQxp3ZPSi5y7UbLKjXiq44HIQfO
uEBAX5jVx9Qj8UoHdXEtP5zpddFMDZQrtJq71/3h4ItjbSzaxAUBMEnFKvHT
eiIISaRtQsmSQSOPPxa/s8XOWlVheKxXd4AiS+bZoN/sGFQC+Nc43sVM2i2S
8hUKyzaGPKZzaEyH4BjC/bqo0qpn2L+7pvnC0Q/xt3qdpVW6z739HL6B99BU
WSPpmkaTBQrTc7ML6G41DFaR9SFaR0F58XwsSvA7mqvZWZ43flpWtWhQtGUL
CgdCZzYgmHcQHA0qGHMFFAU0pzDfDKICeo93j4fKh6wmR1atocDjD0VtzrkR
7K/H4udU5/vvcIyLh6T8K1/c8noUauzrc45vKYvU4aYDjbjQK5HC/kGOxtSG
E1Wj3dQ0E+9xG6EX5BOywXFoZZuYpQikK7TwnXoA4Pr7zc8xDy6l2lgf0nog
hRSRftrz7GoaQczC3s74/xNznsPTRrphRd7hDhELK1XbIcDQ6SWLdfEZZ4rQ
3GMnGV3Ep6Hx17u5bSLTU5vhZwAfKfDIB6z9j0/t02fy6zlhdl60Fya6QQ1c
zDPw95KTZ3CQU27+OtxO1MAkosCQJ2Y2X/jaCI3KQEKyI1j1iBuBcG7I5AIG
6lmubv/xWIyj/wL+44IX/MVvh0GuNVL2LRacHqpgHbAwJohzybkY6gErWb32
BxKZKAMPiowpsh51d2J11IUeZ8nrZjQVE2mEuwRWXaOl49Zwj+e5Jsqn7OsY
n4/Af0Fw5e2+z0NMfv5h0WGwv/TggTZBzHDBySgyyVaI8/h3iqioTB9Q474K
2vWxLyWihW097zTSloojpLfKiZucqo5QWa78GxQ4l/SLeOmwYDAGQQ+9WYYg
/qWiXJoVimFntlG5cQv6BRMEAVOCVsUwU6/BKtuEEfv94CkIebf9QyprdUJo
iVaokDtxMutKW7K4buODXsyBJRc/gwI1gDs4CJYifDZ6Hv/kfmzaFvE63SUW
w4bjWr5n5Lx2Qnx3qg9RNVfSv/APRk6TGUOQWk6qfSNo4vwiAa6mfXRY0+s2
aF2Ux8Ri9rzRQRMRZwiLjSYxcO+2VCJQi8WElNHhqy5O4Vj0iD+24ixBB3gq
4JnAMH19Bxyw2PZPgUCwKjMDZof/o1VOCfTBmbjsKdX4RV3jNa70EauztPI/
Wk6rT+r/kP2ddN3LpBYcvVgQlr3YT9QzeSzNCK14Kucd1RK646BKfl8m93J3
GE77cxLADvPn8hAfRlzjdRtw0tk08HnV1G4W7KQ2nELgvEidLzgAosl4z3mM
Zc5CLug5GNQ9yW3NsfHxEsVInilE4cxwzOxeOkXy6gpGpGUUEYJctegesWrV
EykM0aF7BQ+36mxwTHZ9ht60twgwWviZvdn/0hPTV1c2AGNRTqVDeO4uTm2A
mYEBpB6+MuOJ/zWeoje1jeo7yCvdSmLK2/Zaw/jncJGHVVXXOZhTG5AXLwA6
goYsrFcDi6YJCrZNvgqyyu86powey/g/5gimdSfyZAifzOWqp/oBwGsw74Ck
DGpdURA7n5cuzw9kU0Yqu2N/MyDK4HWNethlZCbkmtQIb8GYAjlwGneAMK8D
YuI+zO2qcodVWBQed12OdWbZ3yHaf6Lu0S4SBLdLbd9CEKTB69Fpqg6wCJtX
t14SyxnivraSXKRuTn0BX1yK7R96grEqp3vx0GlCxiScYuuQdV3yXWWQd1wJ
R77tXJ/ccfu4TeFDE3XDvPUKifYtD0HBxaqeskaOvQD/SW9AIZFyA7LOqqod
3XnoQe0HWkozLMO27M4YFXOE7RI03NNl3N0RfZPInGZ6F/Mg+cJ61+Lh0xAs
GOOWUEE81H7P5iJLocf2vajCEUIe4kY06uySzPpUciCiD3h5CorZ4+POJWOQ
b49BXFQYDHtTZZgnjo1QpmQ6nVWHYO9nH/KMw0IrGLnwXamtMciV+KMKM0GU
kuAksuk/VboWWC7IWEDs/ayBHqrF9IYiEx80GrXSj6zS8yf55zpnMqIBxnso
vEa5p8iodSnzYevah5tlASaagb/Wq9vn5mT2kc3PtED5J1SH6/RclfjroNjQ
rpG9rW8BLW+ZE6A4pZfSOrxVWXkXkljvhI4PWH4K5vvba3eia8oJ9R7/6Obk
JzwXFvnkuNMyxo/evIxN0Bi9ZoeWvErDuTDtkS8ZoRFJwJeg3IDdJT9Ar7GH
NLwV9evUvOq5jxWn9gFyWBv2BbDctZKPFSItAaNPDeIXt8PUPZBus2Pf9T18
N7HMDyMcbshLXQFB4jRh+U8DNr2TyMd1MnP62oDJsI6eGkLxp6QvBJQxflvS
hER0yhARASwpgG4TCoU3EY62LWcWmGaqdkhxUPSsy49sbaldSDy3Fc3GInJD
IymomjbxKPePifbHxMOvVTKDtjmF6/DDYmVVLVzHnKDrs0QuuApzBQwnACzl
xAgxcplAvqUONCbFo4Dn3mB8A00F1fivdBGe+//amJ2sSz/tVIcWKq2GOjyv
B3gfVb3hVkMNZRxLDObcMyQP37ry0heuzwork2m9tA+u9gZWpyiD7LVze2iw
eQHuZLN7ASGtpxC9a725hmst1QjGLNBYREeqOiRRjCRTwersKbz7qqERCxOS
i/Dl3Vj6spwtoWIoY+lp0OpItMdS10h4AwKVSS6Cun/kXP1V1Wq4xZKP2x/S
P6DWBUhb8TDZ0DCTwgpkZi1c+InEF2hBJ5+NOR2fxvuCbP1FtfKY53dC8+r6
1aR55XDr4sdUA6gDsKqR9k15geURDENEkfWtAVnjCkkJWp7zAAQ65hvWhP79
LWkit+qOApnOfuBXRakCtRIcYgGpl94iyPqIIWo3gXlgJxq5covX6I3g1BKa
OnaqYpiMoWwU3ka67NqK7HKmpgZNcrQ+X+CK6fSviiya08AVWcMYAHCIac4g
Tlicy3pSn77MOZq3UiceqleRjnAswEJzw9GLQvWxVERh8WB1en/aXl27C+2O
dSVms3kI1U6PC0dAZ5di4LKweAx7NIoiGDtRIIL6BhD+R+CUBCtXTNJlsXVW
3ir0qRQPZWvrBYdHaxbSO90jQqEO8SPr60X0aCeKjPIvimTYFNtJeayrApBS
hlCvBp1jUmzEkopaXM5sfOaoxwrzJthItuMEnx0w/UMzjXrwH6Kki1MX3qp0
ZorOOx+OemD2g1i+GtQDgt38uwnkR/xsOcAujkrcuF9k9T9VzSo0EV/wLms9
iqG3WuTloxcCbRBw6z1uhTz2Yjj3cWYdBhFxpQddJOTFVISmSgCo8S+MYahB
0shrcnM1UnC5NfVE31He2DkIBZBYy5Q0+BKeRKK+aAACzLcgi0BZVB+k0azt
XOqePlN0xjZfvp4uJ84FrRrYFiSO58xqtNSFR9tsIjsVjoP15VCFTvueoO75
wXmVg7yVME5G4Bl25NUUnu5BcgaQjn5rWcbJpx1fLi8zPyhP2ohw8Y8eRfE4
GfIVb42RMDEj/dnaIE+iAWv7RWfmuzFBZOQUOBWnSuAyCWPbyxoSYWVGAzf+
a7qK8OVaXyi70f36/Bve6OHqL5aTMZ+OLjvt3+TM0scMduX68GnAEQgjMpEs
GRCAm87trk4pW/z5EJ2k6Z20ICAFfPaMOaXcjLurn8rVr1RPJJUG8nWkfVBC
Pz8Jatjuc1nqIsFuQobSPiURdAzvDef//Up4b9qfD41Lya8b53+uhZEdrTYD
kZMHSiIPxl6kTjwi+KljOVXbh1NHWS9TngPtMy3jzxzkAApvmDAIwBzKs4Qz
UaySBAEQVlCjlrUlwdhtye1UeCLNh71oRV2mgECwDL0fMWms/072nFKkCQ5b
6cIm/Lj63I3wVl2Y37PKRVytnZCw69ilRcykObyTJFGWlK3H4PkM1EavxDFQ
viQ5gwbxR8CCpzNWoFOGmFvrTXcKTn7roe82bhCTqk7N0lISdjE/wWQpJsX/
+xMmL61wSmSDZusniLnZctFnczghFwAs+vohVj2efuXGxfOI4PbxIOQr0gkw
SsHJ8JVhPcQyWBhEPuxZVvaELtn/Eey0RsZAAIIQNpVdPdMfBtJeJAbiREXy
vFDcux7U0UphKwAxI8uFlzl+LGNIAp1NyVqmTSKxIrMQeb00G+d4CX9hTv/N
brgQU5P2pVRP/OjAAahaUdiJ+p2e/pYIfLtv4Un7BKY9cLNxk3kCNfGpOUrN
XbDO5DYxm1E/2c0OIx8iDyYah6DH6jEuJp9UTic1LoIAwDI5LXeXe3xiaRD1
KlkPDuknMKFiN7d2BUquOEQTTjBJBrW2mVZJfZlRkfg8EMHIctmlxwA+O2AN
XvOymR5eYBXynHHWtgMo7HD7qG13+Pe2VzAf69hHng+w5uFJpwu3TZOsWWYI
2w8q3OcqGnAEBka8gzS685gfsSsTg95rGwpZmLAEEfSNuW0sbMtKV4hOn35n
fNi4ZccAZ27aEuOxNaT8IVn0mwSYkARRYkJJNXSdi/O6xIlRYc7UMgghSmCC
I+drz++KCBFGHk11BZa+4/xOSZUhJE+iPRcCRhgzcjiMDuiyWJnrPzB83ygP
7wKw0GAk4a1i6C3mV6H2KIt9CP7YooYtlj+PqKhIRXW7L2bjE/db/dcvvNzK
0+kN1lkxOaPMuW5yYeOscaiJSWIoUFDqZheAR2DWvLY9WH+DFkwEyBua3cmn
aMIVHPVvrFI/cqVcBBZbdcsOttT0yu/afDcsSlevhIrVT2oK6k+9Xs9muIUt
+Msz/iADsu+xJLTVf9KisH50QFwzAXtaywVgcL5Pa2q7LIoyO0+dM/QBdFJm
YcIf6mTB4j3K6oEfp5LAHmtMBNkslVI0d7G/Oxwb5YoZSj6SKJ/6DMY5nVnO
gG8V05e988XgMJRxoX9acVKy62utxpYsmFWUyg/a5fgXrMEC0ZXFHGxm8ARG
ZE//yqfcm6wK1YAu4HnCeSF8oVX6bOHCezYYRuL0jlNPz/SChJSGypMDx/rj
cfBuZuTZ3u2f5An79xmAWotVI+KdbFECa1LFc4b2wHwgBTTR7tPv1BiJ24OX
vvRjLf+7CxRiVbCHsb1fu4hWc+4maxSIgUrE5G8YuEOciXdL9DGVlIMk4cCJ
+4O0Hl3iOj+hz6z4OgVbQ81GdvHlQ7h7hNYhlNBTI9/vBHxdePrBDx5+ujir
Lt8iC6d/ECKlom8rRdzQRvZJK+i+smUVYzVn0TwfoGXIa7cc4YuIjLAPEMmM
8VrrpWqhG10LkmLSvTD7WPPrEDtnRDLONiFaviS6gAdI/5PC3nlqwvHr5elS
DkzcjGSdq4HBYcMZaiqS6Q+S+Za0aYorbEpKiKh5qPe2E3Z6vPvywNZwX3H5
k1ms2XBUHnQKGlgY+d2RJOxpzYSOW8FcKRU9rCUs8opPS1VW+C1WanPVgU5h
VCZPWOMsFAA2G6p/3DSMQ5MPcg3tyJDkDqxdh4NxQn/J1pMqn/tg3U/2sCQq
EQayEqCWEXK/aCnx7BZJIeWr5GpjSGFQr+kVJbxT3tABSFippwTURwKdT8NR
NHFvLwnfOvurjuK5Zwp8wZZzBHpCGVNN2a9N4I1unLuuccvqD772hTjoejMi
vZDyyMcVxtW4YvFe61KOArXlTmQcMaWBF+tQGXmDzYUIgInCcHKRFRuPlerV
5XmlJnRHm7N34rxd26Ys0yxbS7ivrmD4jLw2C3HvwEVgSbdtpgA477vVMYdK
C8U8IDsWFd4y2tCIKg73IAMNsf5imlGAKNFsBObcjrH0aJ81pr3J3Q6Blr58
ixsYBfI8m38/LaiQkSbBmufvbC0lcnGLtgTiMykfCbHVTMsrkwA537LA6TjR
KQYFXqqiQc0UeYcYk8ROvV0Styp8lDlFKSsvjt2wtlXTmtUon8AUO/218jS+
rn++RhBBDJNOjGhgwncZo7z7FnarYO5LEV6mbVgyrwd2HguU7AVmQ1OvN9J8
Qfh7x+8L68WMnE9KoswxMuxS7lszG36xlS8jYGmq4tGS5+NQC66w6s76Bkz+
ZX6SpRyuxpkjxR7nCEzgwVTBoL13yJlPjCrh8X8IXvVw8jy1Qz9fJKYU/3p2
ttXrxi1CEM/WfMx+CwqWulncpiu4zRaxh21SwBUt0VDLvxJzIWcozy3petlm
H9jM80SWllOtU5IlTyRqOqPsLrRmt90y1vvpieJYGSssmtgQh6jFggvqLzl8
42w7f3EyNIZWSleVGUPqQS80I+EX6GjfkudLwUmJ3ey1t9PRb5cbSMWUP+Ul
eBirEEXIWJE7C/Lj5k3osFZRF/jMSU+ucXLjzfuxIpZcY+YqI/PkXCVmHA8C
blafNy5/WVlhdMnrFsOhcbZc9wRn3pzZDHdInRBnxZO2dZJoggYZY+bfU8Bl
WaX2tG1UpXdHyGCaAXfUZqIo1z2xzPiQSrQ9fldhFCSralgNTACDnyCBaCw3
Kx83sL09xFGHRONhUkfo5wu3XGaShcU/1dXfv22Bjeiy/tm/QR9dNYE7MjJ0
gE0CpLcqr7HwDWAtucgrjeykBhCA57rFdc9cvHb9xlylQQWLaXc5lvKdRB+r
BIy2yPTPb5zPpSmLxafut2Ly+F4ovKgX/+GLJit7PhyXbnxMnaxz8KCW+3E0
lmJSStbDQU6kjQzwFa817iurqHbctslBF62m//5dakjKqzVOkBOcYm4f9p59
PFEIGNA95V90bk6idlqcm50Drliq+ME3tLpl6PnLExBer6u3yibP3ftA1/3k
sO/rbMbsRp0bjO3AnOOE3ftgGKsLLBC1UrmRedRzQTG81T6LjgFoCSxjz7fE
rnCyl+Ljz4AGbJIzPT0Cpc9aq3MdHleVIC106T0KIRKAbYuFAJjn+MrdMq8U
sFjAGs+P0FSwSbXnEGnCUd3sbbgrinocHU3lyQSchbsYtFsYVmdfxo6WzNpJ
Vp9NQhiEKqmIsIbyxPNQ93cEQme6H3ukwpIBmVb+uk4Th7tQry3NeWGpR57d
j80ZoexHibfQMuuS+aWlBHr9neW4PCJ+jMC0Zb6+TxsGeV0APJ6xz62h60zf
GTGoPPzOH9Km8M7rocXjqbRmzmJ9HtPe4Mhu/EM0R0kNV2Pr4LJYAv7Rk6Hc
qw+eU72/HGDJwWIMrbnp4KYeFXXcXr+0koSa+L1BZqwSBmEWG32ecphuS5Ip
mCtrndVQiHK9PIGKDND9hLCTUeMU/Q/aN8T880t66D161g0XEAcSSt6xXaWq
9oRIFjTUaPVHRdXFAoq9UrbpXZOUwEbFHJ6nQ9CyKnoSRiAZ5t5P7hYLyUwU
upDpw0DL4bYv9ho6rzNiMZYHHHIiEZ1JaX4/G/vz6BJwKTVbOPvbl4419TeC
C6m7M3FjnlWS44XHjPyxvcOe6fhZ8mgtsuJ+gqFzhbVjSwobbCFTlm1LYTsz
pOJ1z8djTId2sT8Q2Im+9/ZWlCYPpuO+aNNsEpMCYKWmuYAHvBPBmSAyZ4tc
YiHYynRxO+vnPk47fxZ/LICvyKt/ocVzf1hqDdNKjNXWPY6XUa8+C+ezBUsl
/Gu7DWB6/zOSRYU5BScnJdvqPaWcdU/vFlWka+eltqMNJhHnnHZzJeoS+o34
fQtAV+Q0jEHanm/FecK7ADANNAqj7PIOjEOc7w6yDlBGxGcZduRHjdwv8rSt
65uZLzeLpfocuM6h79uyepIstT5CuM2f0MLDa5U87R3C6foluBiQ0Z1y4HeX
EJXQwyKPtFw8ELCbjvTffvKzUYr/YLoL5S6vVTQGREkUfeRakg7Sa1lNCUil
KQrMxLD4a4BDDjrXI3kDz0YA/rP+uGtFB+lIUqZUKIHZU5OzdSDJWLcyP6Vo
j0frLPJeUvfuK0dn3TtLV80DfX8K3a+xWnbB/4yMCmkiS3ge1YCLtz/Tpppi
GiL12Kv6LOos3rQBvrWx1THr2QdQNxzxy0qu8uQdyLBLzV/unwoJMCxfQ9gm
/gzGiU72XqdHj62EhOBf9e3W8L4MK46vcARDUCi1igvbUSXhNkSdFdlRad21
IyRNy02sQZGBw+OA3YETfeh01m7exeHPtxohH2oEGbKxkbyQ9t+nISUBuFKw
yjBqU4rkPA/IW/mGqWyT7k6J4V9CY3szsgCX7zKrp8lssDy24SC+UcpO54rT
8PhorV/L1q9hSp8wMiFzfYWnwETyKngcp4ZWKdzF9HRY30KU+8qDr6PJqQLV
IBNYPsQE763OcfIgWb9Ho1ZRYiaTrO1JqmKVQWuug1GmLJeCoDjwEwJquHHO
vgPC30KG/NFW/1p+CVPmc7yRDzQKzaLXjLAIy6c7b+5Ub3okjeUR47dogJF4
ZyDhg/MDKBmyYGIB4P4xkG+UV+Qtm+/autPI63/KEcLr05geDiktsv33duzz
ZGXV/wpo7OdkjFWrmkrqPidxBIjOoZ8thXHMizFcFuK74tPhOuRaNHIxgKwc
lDU9hEKRA3BlzIhsyrFQPlthWDcBViFAYJDZG7X6Y5VRPLfXNqQOgh1W7TSc
OQ9irmSKB6Qyrc9pObYa8tKGCmqc3Q17sjHsvKjMSGsqSNH9bbKvkUcM60XM
S9a0VpyogbbIbCEcYfDVa3BRuGcGjwkZqvHWUEXYJRYEi5TJm1tT+ItT5Kvl
GEWAHR7QsAK7DVxLzIa9ZZ7scJFm/+hwUz1xwQWGQsoS8FDglYubQ4flxKWP
Oh5N+Z3gpsimGReYhg4aLlRQHQfUkynjX+ztyTfx0mPiNLZ1X/XYlpuVPudO
dYjUH1V60jySdU0qht8H+VySH2n6YBA8/b/b/hmmkFLO3gdGek94GjPjixah
Lc/iuq6MsY4gQJ1Ly1WaC8VtqSWWHDaeb6CfSr6dF1LvGuj3tus3TpXnzIqI
egDWGhQkO0dNfujSl/SU7fUhWJsC76siYdOBZVHZt7uKqiMen/2DbNyxbpDM
ULXj7PpgiWhdun8aFzxoKPm2snns1HCkB8cygtg3hEjDPsgAJDN4hHMMQ+I1
2RsnmFMscCD02PjuG7IVnNp1WrCwoVjT2V/RkinuiqBeFfcbTiqmaMgkFvlK
rEQHZi0mtW1ShEeW+aNhdJnPxNcRZWKZ70TaRQbcSkYqHFdirsA799bJt+Fz
tdlFqKYuITJ25mours/ppcEpcuYZT6OfuJFBCn5yrw38yvr3yeolRQbDXCXZ
mVK5xwRc7XVqHhVe5Bzry/Ui7FPyx0P+I1LZJ0nT+hnsxjRNWvZ+Sjj+hGw2
FWdQiPY2/nsbBiwfyz96pn7cTooILw88VyF8OrVNqU0w85lxcZ99RdxLKKoD
QDg6/mwq5p+PKMPg93c+ucj+xVqunQxpkjAhLvdCEQqOMqlsanuhVpYX7ujE
V9Uv6UEF/1RK+/g27ILj9CnJ1Truqt+f4BxSCEzZD975I4h/0GIs8VrUaVzf
e9zHQF5HNbcTiOIOlKaamrlxWTJMd+Sgp85y9zdCcu8UM77qivCRKqHElT12
Cq7otlSbieHvJTwc6pkxNFZJy1ghf+5ZNtff7I6bR4qFUeIEu/5o6HihDGVK
cX+VQCACS4wqZRbYgO/qgo7kbZ3Aln4usGocjWuXomYEn33wCEooNayQhQ3j
yU5dYOsodARjJjKAFdUFYCI50DMjUvCrTgPUA7skOBdGomrK6ZsKlO1RUrk7
7UHxJGnHJoZ1pgUU00suMMzxKXM+/lNY8a77EhUevPXaPGTtB8GSHf/QA58a
nQ/O5ZZmpJtKmZLD4e2YepOL3EsYwc+pHa+GMpv9dJzycmZRCcSOncTNK+Mh
la1ESEkVXjLhxQPGlUc9BZYZV/HincfVjMuG31WjreHy2eGjukIWtBKgfTYa
sjyx8hcOdaN/ZXSCp84qfbJNNoXfiFDb82ccO4MOzL+vZp5LbgTz3Kgqp25H
F7b4koqblbgESW2XVbwByYXaC9kxCvefgtU9HfjdQCJ5A3eHn7Ifa1r9lmKl
vspf9vXdYbwypfboch+r3fg7WDK+KonSkuK4/0avYpGla55hv9Ud9UaGi2Rd
BfkPnuaiiyGj056Btxy1Iy7lHJ4CK4Ni3hbmlhTN7s/MXjqUTUWMDUudXYQX
uzUKA8CpZvJCoLcvEcqhT1LWsFhjQQ4zFV/tlrk9h0WWJ//0VoEcaUZe1ABG
NJvBZ9cJC5l5Q5/SRyM7G0zsKOEFHq8KKHGBtcAFGwW0flecm/Gty3/WoetP
iYHUGN0b0+5+FkGe6u7/2RB8Dc05xE9g6buVaF85brQK0Lc91fuwUbxwmaXg
BePJlqyPeVprW+7j+xRszyyTz1ffbYaMLHGW21F+ncZfA5Y8J6fvpcG/rL4l
+b8GqTJxPSGXsouWuCCVrWZ/aoSCPIx2agVOhjZ/xeNH3dkBebuj37D7p4ba
OmzfPW1AImPDKOxOkzbswZ7W+K1xGlf+5Lk/gJAjZoQv5ZSkuA7hs4Q4usxm
SbCrgEhEzi3viW6PujEUkPShPx8kjhuoBYwNioq36E+q+jD+ZvbHH8tz+MFb
N12LcWOtPwl+La98jKt/smMrkgQQqEiYKgxKwHE1UnnVOfRGjwnQrO45Ggv0
i0qYr4obuWO7mhylCx8q3zJgwQGn+Cz3MLgGTSIA2hAWLk89QoidHHSCTqyY
AlOvWC6gMyF0X4s8peAz8nuHyh8dTyGg5kDma5M7qF7AI1xfAVN9EDbci8w5
eFQNoUyMiUqtpflcfeIhf0Uegw9fKuzPFKvXqcLbSqtnScfIGC19Q0EQRRZN
pzfKsqvh/w3muBgnCUvzVzoJOatVIXU9xUQcyp3lsxQ/k77l5zYku+2UB+NG
W5yEh4iTmbQv7b/YaDR7GzuiVPvuvBHQNHgZZT2VZOOlMA0YdspCjCSXgVLs
2G0KkcITuS0kpFkzifsG47cYf/BrnU1KMwyetXx/nTCLqIRd5wOURh7yBBcQ
XJWPlmG24S1L4/tJ/fX5jIqnU3dVPNF3GwPWBc9HzgYVGjNPEoWsMtWz/R8p
qEk1gEt9oLIHytKH8QML9a/NaOUgLsN3jkpQ6i2Mx4XBoxhJvBdrvEXqbETV
fONHa9D+GS2WxMTlMx6unQ98gTepv6l34xR3ADQ/FaCUnn/gLloTLzDsUbXj
Bv8U3NxEM2oaiiFkrN33YOBh6k9cA/b7VVPCtFsvv74iycwfcJL4E9SmiIdt
Zagqdg8m4EzMPbYgR6FTN4ioK7PltOM/AWtBR9PSF1ae6lm9QufWcvv2Rthl
8Azv5xm+5mI0ny4oGW664wFM/90P4YzpXQ+LLm65yVLjam18QVWsYtW3gT5z
oyNwZdAXddwdu/ZlmUTin/qjFknuwfComEZ+Nsi/joZdZiuzkfEvJxvkugHF
o0Q1iuMhKR4iLcZenk2CKdQEkSIAYyQfqOdnmjzVvDSsaDH2UuNcC0iEvvdO
0WKsiEvo1n6pPXykDXQvaT74UYDC4nqYJvPDpsWVCycFlNyPLUmtbKl2WCKp
UqL8jw1oKRPHyhZ315XKxW7mmqQUF8MkOvx5Tf7dIthiuRL5a8MBbNES1Y25
pY8QowDMl9GlvirnFc4yXa3Vh3jsaP1ACUMRNJ+zk8+7NfW81HNeR/JfUXHW
J7HY+GYB4gQtQYSuyK/RdsCOWKXq2BykYVY/Q9p6D5GxGRCNb4Sg5Mdsi7mI
CrZMO4JyRZ33YXJmwtJD2jRQaSXN3OY+xJVZH5mbbhP8T8H0xYt6q7+v1KYY
j+5HXjdAnGNbH1QRAE+EZREPDd1f4gJh4253C6BSpRFZbLtqpcc7+V+q53l7
+XsEwnqzTzzrRsUHdgNXV+00SIXe8a7DzaWwhhG1TalwgGDhKa/0kYoM1Od1
LYSah97YNYVvElPr3O81VptUG1VZ4I3MduXKWDj1il05qVx3zZV2YGfb5CAL
aBaKXSBAJmc4QrddPBEWIZlabrs2YxatjZANWQhMPOM83GtlDhVD7bzqSOMP
F91qGu1W37FVsoyyRDbYxFyKOtGGc4cfqZU3GOmA2HGT8+opOb2YzMgo6bjY
E7ji4BJQycsslVmNV2hbH2b8JLpGzsVoU6AhLs/BLGOpxfGQHnEm9Ehd0mQC
wdgMM01KLSf5pdH9h3DCXvcqKAIStHFp7wdmecvPqtUhMXBEmIshhBOfRnod
RtUihrhyC0nRBjc48nooCa/Jxi2HJfF7eF5Xp+8ABKF7ALXEi7caI+4/Bbzt
4o0bM2/CAahumKczqpmu+HmwkX6aukKM5p5J3SwUycO894ADw5Km/0tk1/aE
zNtEzCOkifH+tk2BUZ7PAX26fk7npAdwL5WzDBQNzkPJNdL4VJgBjrQ+HzEn
kBNvEZD71B4GaZfczRpsurVrLKksbOLnH1A3aq4MTAJ23nP1Z/8Rh0vLpJM3
2PT9u9dRdU3wTK+jljPjGo0ysuX0Gv9+TuSLm4LjwYrrta0VxpJI6i1+J4Br
0qQlt3y8gz8OiXz3uwR/AGlomQpqGprtqvk8kB9/X+chq6HWBmVfgzVvgtwi
tb0PVBdNEApX5XrIigoSmyPB/RE63vURE6mFMCtJMHJh11yJTS5w+Ai08SGk
eMib3q4HLeztkGwWovlDkZZq92BGZPmpV8IfAl4Wi0eoialIzEMqyJbvzC/G
zf8F3JXwtp45A74u9SypQ+sCAyOganuJhMsD9gDdWJBUFHJRatw/t/FWEN/W
RtzG4IvLmLFODcYEDkoETnTjomAnNPaNrjU2BFC2FxeZCM6crWAX4WCRRRFG
3EKeGZH5Gt7t2mrBDIi1JggEs2SGxBIxn2ICnqgHJULOd5ThohaC7PzJKghu
OgeDhwG+HLpPDAAVCwrg/DOEjec37V+OaqYzZ4KpPMttLURK+9OMZ9qpiF5s
jQE0licQc9r4xk4u/ESXzo7vyPbnSL8z9Bf9o4Y+eD7U2bXH1G05zB5ikPLL
/Trtya6kaC+43szWdMQboXfknFujTUvokhBokufxMUYW0bIraP9JSiNeQ55k
jehXoY4T1ri4S5KW2mgm741goTJ9H0ZH8AmFmL4UxPsD94hTBpkg/LmZIfXT
5HkcpYzpNmI6arTzvDR1i/GWzMmGgbWhVT2NDIRRzyp09bbTw7TW8AEbbjmO
6YehEVLqka9XrY/no9RyDKQiRxrBCzpjWFHvr1z1SIzz9i8te4//KOaCIJvq
yEDiE0T16VB7B4up4VBZUSmmJZRAey8wtS1evQxohbjHO6AcpkHorVcpLift
Qz6/wPRDZLMEGC9k5DrIUV4IqzOFw9AL3kaXRwV74Nlu4k0zN532+QjNmwti
ZD84kr17pDUPx6AhMrzjKBKyo0otxewm/z/tjFzBCvQd5ntDMoF/gdquMu3K
HcxpzGtoyfUzeRa/5ClCtlDPjQPZmgWFREPauza8Afqe9ZdezFZg4dYJWIQU
8br6hmUQofn9JSUD2PPGY6kjzeq+vo5rqyt9mnOF6gj21NIafJIyaKsKAcOb
Cse38lcOsT157Oxoekm9Te4a8n/ZHthx70kY9ykkolyJMVNKN6qhS9o4a2VB
pj1b11PrJr7kcqkpwArRjBlbOJR4CQhsIiBlo01zbmevEuXyus4jD74YSVA2
FXCQIm7t2ASqGQCtDQ09d1LRdioCgEjr/ZXQfoaLoRslIgdJl2dbGjUaBzTt
PpAWnSnnaSfr7JBWI0cTGjYXmQa29YI9Bto3R+350c2u3O3O+U6ODfuJCyii
2XlwZyLbZROr0Fze7IPOpg6y8ZYxQMWhY5Dg9pHhneF2BVVOws/LLQfNa8Vd
2EQEsbGLffw6Cyegx57EwwT7hfrz06/cg1b5jrwV/s2d0O8dwoeNhhfJyWJr
aCSpbXD6AIaIPmuGwnCxmMgKjpOGkjPcCMHCRyuC7OdjsxycV+XdPC/JVFCd
PWd5vgZNRDk9INfZ5h3XLFIjvxLPll6/1Q9Nhl6JMujxgSlh7asyf8YhE5Z6
WBrZmYAophwwD1DW2P9zWNmV/Dlrl6YBrQykSP7zvPgm0AG5YXCoQwlkv+Mo
9M5rwvAHVqjS98kXWLOuWYg205e+HZFJH8fZqPSlcap7FJe7NLZnG6+Iphsx
HpsViUcync4bGEnaYxB7nFuUCQzsBhx1hWc0QpwBq3ifAZbFQkVBaQ3azJxj
VhWFf85fn1m0bMpurQpF1qEN06uetN2EoNztxCYNVoPBL4a5vivvmAzweTe6
P+lPiwkRw1CGRNYbErvALIr1wjx4HybitCXXvm0iel+Tuo9k+k8iv+Uls2zi
hkhwJlsX0z2meOlQeMFKtgLFSVl5zPr8pRAvn/cU3WIRKTUF6319U1ZJa56X
rQB9akYrNieN1ZulL5pW+Ax96DogELVc6EQfQKSbMyL2sZipaQsnxdrsLPA7
1g+O8MdnCJ0EBFpXRwpeSs1qDxEMRXVo8Qz7mL0teLgWtEMIIa5EC6OzyzA0
ogR5bPgktgUZ35wetKvEl+RDXEhN2NEuKOhzmwN6sOY64sSXUovXJz66/1+r
Mdk/+Hd/xX/3epBkJ68Y+VlUaTSfcdXmsBSB6HJ80YZxbbeg55smUimEM2VO
mPI5UNS+6sXU7DAFSnVIb8E3zhZ5i4s3krDyPz5J2XVAxeeT8AUY9L93kmNA
NdSywsRNh/4bE7MOGcWdbs044Iq1ddbx+QQjOR7ZAhwpjGeWX1AiBAcvEgC4
zIDGAykf4LvmvE2umml/oCI1OepKHxLD1nF+KCB1DzD3MOMiECyEO8fZSS0w
PMau7K2e/DbjHDEQ2H53rN2NEnOfg57XfqilOctKw7PRMtkYnYlE+l9I3icJ
csoQ2q7ef5NeF++Xboh7zZbPO23Vxo0RRcWZd41lwKEu6ucSSxFnQEwQRxyz
9DHhfQuAEMmosLBP2ZorylbToIbu9BOP4ozJy/dS/BSBGLjt8lQTkQVEktqu
2UUKW9mdyTCBR5Ihni7XIMoYMo3Rfb6wTSOXpIVdtfVzPxa709mX48IuAC0B
cJtVjZuG8us0/RbsVwqX3V5n/LKr3s/47TaUd3WQlDrzMLd6V28WqNaJdq7A
FC5pVVrGOu9+kX9tK6pvOmVCUvOn2WdD9zkpDVkHBkUoRNJ9duB+YLl/77jn
YVhNjjsNFM8/xHN9U5BU+JEFQGB5LOs6IIkQL39YzTtK347NYKlstzROQyKH
LoF80/n0xv/5pfBw2UF9eK9CLuReY1K/k4/KUaIzrfSw3WVscktUR/muYSAv
jhJ5X7GAxXJcx6WtOftDnoMEs5SZQy9SNahmietGMmxcF6g572PUEmOl9DR1
R4rJ7MKgB++9QXBGU0IOjOyk+NgnoieqSJW23u7bGN1hs5kNCezAxyHhpOR6
7cXseiAQH1nplq9rWiHSJUymm79kn6HuNcLOH0pYfGF9zbNFy1zKejlPUIq6
SDOpGmJ6Tdn3i4gqtTjkPHEQi9gvTO2UsYeWQ3my3RsgZGT/hEORGIWEipQB
VAx51uKQyvF4gVdCGNqilhztIkI/5wM7koi9rw+5WjktT6BSnmG5vX6Hq5/k
9A5/m7H42x/Nd+hyDYfmCcn9Z9X/ljRBhmQJiuSG/N2si5OFYZ79Tq8lPEQN
SIaQJxSNhWQU0Ci9dyDUFiBOGPkPNS4+kHJyN7MgDq25Kz51yKMXYkQ5tGv7
xF8gVh276cs/NliFHEU3NtnV1x42n59wVsooJutKcgYiy0CFZwRs/llWfk3t
USM/YowCG/HhiukA5Lli8fe7X8B08a3786Ex1a46tOObdy8ziyMWsd47/+xm
bs8iIJed5qUEIKwlNEa5yhF8hrbftZdJ3zWGme4E9BMWPzHFrbF4Yi3dBCpf
lLWUxIgkme3zjrf7iM+us0CHIyrnQE2OX9abzivOzZDLMI33ajHztdeLhLvC
SFItsDW7ZDmzIM3zUlsfLkCeT1N2KeLGv2AQWfXo+4OwVndNarFNi5EoFJKM
JLR2aKHx51aW2qQGcraaHawZa3Wr2v6LS3sIv5HU8NG6GEF8XeOIRN79xH/6
g5I5nl9Lx2lHtVoAEbTsypCeEdK7frAwq7ctfivYuEMg3VTPLEVyGIkGZhyv
cPoA416qGHOFlRH2BwkSBJcUOmutxSQitsRNxzwpRc3TIglGJKjySxU3wW+w
iBn0FIm91G7S2kWSQxAGBx3RA3/+7Jr7McapOMqsq5+IKNR0TyrG6jMISn6i
+hR4gJljFrzflqjvI/v6gVdJWNMeLwlPXfcD9ziaUbOGJeZqLpTsL3tbE7gY
QQJ3MaWcoLtBGJAywSVg7ltm7yAVCBr7QwKSDulUIdbgblUq2Mlg5RiHaKpY
GH0z8HhhV9u52gjEOCwYEFrYndjieqv5yTlYKnJOaxrAJntSnfMEaqzYFijX
lDAS0865uqqkp/l165J3GTG/ikJ8H5OpRGFciI1XLWp6bear8FnWBuKytiHC
3YdLBpe1iA/uG9KAozsVjODzkVl773emg6i1XvSNdkxNMDb6hkaW0HKbEjt9
Q7hUTn29uW6PYKJ3fRpioMOE9AE/NsliDWtIEmtFbGKM7+dbDL4gUrUL3cGE
DvN1tR3zyjM++LoGWtFaGSI4rBojMHGM1yp4JdrlRQm+7iqNcOQILVBQKvT6
h8th68fqizT2ry5M5NHad8KGM/1Jo1AO1WZ4xSQ+KfS+yOQeXppcG/2WHJHo
soHdUpfBz/3j8D4vFaidfJ72FIGWFH3uSR31EMHHMv+rX4NDRSgvEHlKIM4o
gBKGAO4rgcS1Ut++1I67BvmF/gsD5ebgjOccA78ar6yYP72dc41aQdxlvVNZ
83ToFD+QkbZrIz6OU+JfvXvGZsFH2oqsGYEEGcwD7biBIe4I6epRSqglukyI
UJC7gJO3c/zuF7KWBNEgol/bHCTAKntI6chaFHQRYrjN4UHxKRXYbO9qntee
+cEhYhMkDz816BjqzCIX1Q73QPqNOzrNQZfuWuRZzZ1Lea0ms7cV7OIfjlkV
xH317Gb9CuDSAUpP141S3f38jSNbrPZi7AdAnfJ5qOLP2vHbm33W0MPmDvQs
eDFMRwWlh+w3Bjo5mZDYMK8y8OKEAOyzb5pRDLc6atCV1U29Jf9v2wRzdZpo
4Kamh0JPY0/YMjVVZYzYAbnxkik8rxRnAOJRWsQxxvqGAElwrWxqCEeSEVn/
drWWlfT6l/LG40MjZt+KRWSjSmnSubyG/zjxIaMPEJfGvYqbGchX4h8oHNyo
1ZIAQH4+NRisEPgw9J78fw4qcJ4bZ76jVgSwwyIbaUgNkKZD86OjRqPuEHJw
KLRxYh3di+vHNrYKqSQPqXNY75JP6rya5AJ7HlK4L/U0CT78UokeEw7bt40k
xn6bJzgo6WSPdVP+NOwO8RRDUr1Lq8cV6TC/7oo0C4aCKnPYeYpeZ4a2Rp8F
Xcv3nNxFzT8Rmxjxw1lnk+Ya0CQcZx0SKV2t7DrOBjE2EzhaGMu15DfOirRE
ORSrQgsySIKmoWL1yKaVc2/FWvTYdSkWtGQBGlJaQE7MZfJMAU58xgD8JHXd
yQzfkQvFJURtKdjvNDny775FhOiHbFecUFVNcr9Eqxiprb6aHSc5CMqDaxQQ
HnGi14Y4d871vDfkuCBnSeqMqSf7SWAvyq5cKsuyasFkdoGEo1HuC+Y4S+kO
iL7U+8Fn22vDjkee46qI7lGSpRe/+O4cTCSh70IRAHQfmWNhCu9mCBJxe46a
ZI3MoQMGEdiOOHNDCv1lbm9LgNP14zclvr53Tqlfp3Wz+UQPfAvqvMiz06O0
bUuRTFLAAfZAF/1XvNXHkry0nCi4w6mgXmhSWSxFosrUIjoyobiOpP3PlElr
VzVTlm30pWK+vklUX4d7wGOSEzXB+JeOMaEupfFguztVjfHKOWbPoWexMrYd
q1iNWKr05tI9bLMl+8a4cdZfKUnr3wnF6UA6jc1dGrz4xBDb/Z316PloKUoj
4EN7qTZ6arne7kBzSOJKFkgnFREz0qzpte+emFSVPx/hAc9c5ebMbrGp2j0k
kbIU9jNjNszy5tklLsB2WbQ/ueFiiw6C0/UpdxtynWbkViS9PulwM94Pgess
q3jaDOVOZMSUojVZL1H/95yvf8hshm9FGM3aUTWRcb42U3VpoKW0SlxFGN1B
5x5BTYmaFEIZp4jkQBnhXU5/REtoY61T6NZY0ZhMoRoIiCzoxDVgXACgiMNo
ggULCERQ0kyxaMtGXyBAg8+CVTuyIc42nnV8InfXIJDRLIyP6OWWgBAemtrm
PMlO2tgAGyFC5YcNfaC4PBAhyuj2YY4aru+fJLsiPKr8PWy9/JifY14ufUOh
d7ZR965J39wDwNpJLhLQb3qoQzRNAKOMsbZ6JqxvjsqHMU+GCWuw/JkCGN4Q
2r/bexI1ve89vOp6KQmpA6/2rZ9UMXjDN7fo+Um49VlrOu0pwquhqac4Fynr
5D5Njm8Flv8mwP0Keiygk2y3xFz3XgL3QBEsz2JjSe4l14boDis6M1Gepzob
k7N96M2ihWXIN+IfA5UXDJhdyA1EumZ3bni8x1JBH9U6WzIfpJ4G8Fx3V6q1
Ps5dvGAfISslPWeFANDlf7zMZUIX12kqbyaTs2KPcXG0U06+iZc+v9j9TEYl
PuntXlbpSRKH50oM8/bVl7c14qJJLv5/ab8HAitnjhCk8b5nBvsNAzX90V6w
1HVLJ/1GlEWU344bQP5gBfdcZ+3JNLFXQHKuVnkZ7Q15hy0zYhVqjjUf19nz
ovDbo7ET2W/+HZRWMPxiKre4PZfHq6lVBrboIJ2hOBll5dbZpDTuz7+P3GiA
xG+K5lB2FNL0F+ia5xhtxjYmgFM7v9KxjRgUatCuyTRH0cquqcSwjk5F4uWb
zHd9zaKUoDBs5n8+4ywDFFKhIqp0o1ld4DYGZ1p+eS19nQdnyhiT8m+8Ccye
u6j8JLbi07ENBhQbxBjgLe020uxP5c4v0t2ldQwUMSkJ+jH/4FTFbfSNaiHh
oWMi/MPO+tL1lKb8P5ZEkcqQNAxHBpH2m82OPiPlrFgvUJQ8IX/F89fzkwG1
Wumh/tMO7JteuF7may9zn3KJH3viKf0NOAuMg/AGxtKUZBIS55b8Rfbliq7p
LN9vpBM6QbKXCLObVjUNGj4+xqVgdrf5xHj64omSJ2c3nnKTqj8iiQqGE4jt
Ms8i991WppXchAlVQXB0u4LChAS73grwXyc+PFLrwV2lrJC2x4tFu1v0+7VP
75b2f6/xqN3BIbGswCQqRrMHQcISBAjkfad7CEajowNhhbtLAKANFTpetNLN
phjZlHz2HhJ5TFKyrZJRpEOfmlH5XDDQDN4BxCFk1CiYKr0p5BTTvWts5ngX
CGb4b0D5S6KLs4acNOrMHFhRCpjwMPGgLsah527vFchWA7pX3piMmEZqxhd9
Oyvbs83CE1IZfik4CCmghk90GAA4VYA+4khaN7y77nDMJXKzUX1vm0EKgisy
a79XTS00C92QtzeGf/VwKSkL+LZeQceg9J9fy0Q1p6iYQ7gLWyPboqBSbdzW
kjK1eYhuCa5nivFiXSz2ofVwdN5p+JQeH3jjqM2eMft345ueiRjbPPQSRQxi
ObtuMd+7BoggNmW/mVND9g4dnLlcZaULTgM89H3wf+xqNDTlhreMkR2C8gjd
Lly21AZJ+99G6R76CigODkC89l9SLb8p+MS0LUTKUnox9ZBUCehJzmeqIGEE
9WqRCdQXyPAq4i1nDUUdTiCgInI0l/L6roQkOENuyhWQo8e2cvjjinpD+ees
vX2MR53R5yfWq7EMqH1X7pCCGh3x7hURxjWCk86s6eB4K5vhAN+CrwjyS8/a
nuqQEEGPi/G/AwnWFvii7aAkWArO44q7QOQHjslGnznFearm3Ah+aV+CsXNr
k7ME2m0KntDmxBOSXHbvJkIxXRXp4rzfTwyRgfg6x8X/O1ZbaV7TFP+4W4Vp
7ktWn1CVCIIm/9GRpTWb/QhsaYIDrLFWYD8agbUPfGy42dGdZFKlPdDW8Un7
OiADYQSFjvBqzoSEmy+w3vAPqaQLMYyzRjBeMp9Ukp/FLi8Hb/fBNPntq1N3
Q9rsVtcf030lywm3eoHrTrpZ+Wy8Oi8DN9JHvrjH7TvB+0a1dL9WbTJt/gLE
DFSEvAQ4IngUQLAtaAZBXdK9j9MDSUFFA8LSEZuzlRE08tLKHAsKkpgDQ1WL
PNcw1h+kMYY+gIqpGtMpQPngQI6sQNHvVzCDve8B2K3TJKGQ4PfTGsJK9w76
y3EuErzH9AwppbcyONmy28l2ByMPp2soi+6lerwhY6uUNfXAeuDHyjYMfEzr
y6NjCT9JAIS3h951fXKVVldVxX5WsdXd0RN9kjOY/N6CbRK8ETjQ6GHtuNHK
zNOHyxGYAUopKu04x5hPBbpGMT9scIYyrmyRTcXG0JTRUYz9bvPHxB+JKf9h
I6EqNpji2NRTIQERmKGKWPr70SmxNnO6lNMLYAiyPCnj57Ab7peeuv3rpsfB
H5INrOvgpLLqYXsJlSiHiBoM85jgZYiZLfXrJ+lzxk8rSye3Sa4TfXFKoAuM
htZs+3xNHMbLqYLoZ3MNCdGrNBd2kiEua+HJu/nh4z1tWtCdL4z6CHKR8mpw
hw9qNrIMj7NCNCWP7QDuC06s+k+1AqL6Vvykp8ZjRr0Nn8qRvzESVAW666RH
OYHOrYuWpPbFZ290mzxl2BMdpSbS7FhTdrh9uzihI/2kr/vk3IuyMT1DDu2a
H1ItzolALp/VzDoZYlDmLzlGJLZcxI4eB4lBDmgnfjbBE3wcDrsHtGl8s/Sh
3eDVmgfUkYpqOlWq8686ttV/AaSSdrfYl7qkGViO1JC5z9pEhT9fEkmv8vfl
dGjkzoh40A9HUZrh1QJG27kNvmjSEEorIjUdjGdLGe4klEL4AzhSgz8J/unQ
w86KHy3AWyMrBxOa6Q7XP+FozLCTUJoLs1PQlfEx39bcAMgBHepRkOacRHKO
XLWY2RR8I+oqumOGwDy2dddkEdeOQjapt6xu0IWr09moPIk4uP9bu/IYOsT/
d5EiqLHcQqX/3ijnCqh3SNVkMZ2mB5XSevhAa+cwz7S7EMy9hYGSFseoBBjm
yxOwOs3DMGw5CsnIiwBOvY7zQU9hFcK22UspPfKhYckH2hmPs5B0QXOT0fMN
Rln4VPiiyMJKoocnaumLXu/Dr6e6Fj7thJYn4sjy/f0nUnbTnWZX3I3pIV7K
JfZZFoiPeV/Byi/l8Sh5VfW2RcA1Go5Fk7oV1e7Kd0Qt5CyZLtJh5rre054r
fmYtwUhXWQvHg9vCLohP/4D187WsMFPl8zFuMDtXTDktKXTZFOj5z2YgRxMZ
LV7M0pO8IPzvXzf1AyUjkizInQK+bRTS2VwWPyGb8IORSx/itUwOCaXxUPRI
IyTNtRsaOZIjtVvJW1P+DGCed1ZvnTS2Yq10kHgdQ2YC2cmzM+rllyWxDvsl
s/X+sYF97+pSlw0HaEYOwA0hrurYqD80fAo47imY0YuKcRlgWwrAlDgGvLCP
leU4pqTnH5XOGLfpPWE5eAJLYQWsL68NoY4qHU63CrirBy/feXpQ0dSjIyDI
QFzYOP2lw2tpX1yAHH/YGlP56SRXaotEeCfG1TWwOPuGhhRKZGtXB0X2X7FB
5JdDeDXJ16gtG7mM5MKJVvWCN0djF1rj015bCAS2xOkhMgDMkZIN1tHrNi38
GobwiKefOdHPgwx8CffrkLQheK6Ehcb5FwPFTmvNQeHPYJ7fFPHSsFujzfDN
y59lnDeCbiXqhrbAoWsv60cZ2t2e+lfL3VzBRQROjfSQs4N6USe0TJz+rJ2r
beH8qmq/8mVKy3Idzn+CoZWCH4waP13gxdlctvgvE8HCnSG2DCyccoKRzBLe
yA2LYP5mYPDvevIe256JDn8OO3kb1dYdXXNP5EA00urP1T4JEdjylLKuvAxM
4zDCYF4CyWRupJQ4Hwgo7yyxE/0+HT8IKiiBkmkgehD1k59Ixxjjd0jQFbmQ
8FiP+oQUWJ1h57VVJ3HNu0NUR8ArU+Ci0igIdUNpsna3G1pswfTiedPIpW90
sQusNXz5u/fvK4sfVR4Y5zmgjrc2qo7f/oqfM/7z6pQRDaij8XaOca2kC1Ce
sz0Oji6fq8MfwRZ7xSSjcft/nznvjafrwfhKvLqQnq1fTbinlVJj0uRYpbPE
pKLeP009cWqlT1il92w4+MwrlnQj6hhn9eN4c8k7GO2Evvz681AYS8T5Z17N
oWqp9Fi1qNis+uSmt4uyjXB4BTcwZ2W6sBTtHFS4nbLJh+V0g0Ambdlakmys
JflaL3tNJ43D+rTsvj+THAlPmBZktwqrXYJ0uUOGVChXKkMl9gRYmm4uuV6I
0vB/IpnAwrHTm+HU1trXqzOYK6SdgSCUY5K5LAGUKvQEyhMnIfV5+/nZXZBc
n21uTTsbSYu9XffahUixo/CZVhE7taS3phskxtYeVyoxGsuRM3u3FtKNOl8q
Hl0CSUySq4tnerOxCiyw101Kq0UeECluwnPpAkOXHkWRCYMV9Vao81/jvxNz
RnDrhfjTrU37SQ4u7mRJH1KiUa/HLt62ExmA23zLK7SLTKpHmWyovGdqZHqS
84dXHDwBEP0adaqui/xUdrwsDHsEFgFeHxvQcIA1JWS1ool0F3++ULVQe4Ta
Fc6WQF3HaLGJ4yFawZqPz76bQN+Pbe6n8KOWdr4CYkZYjTBVygs4CFrHaj4n
Y+cojo8PE2GGMLWjHyIB6hj97s7uYYJQ8bo0iM98k991Jc87cj2y2YnSGMHf
uKHKfwQevkAANaBXKErtTjQRAkhRLrWvoKpBMTS+RgSFWNL3XQEgSNBjEi99
yVbnF85smq98PxTpXLZxegAxsZXKhHmYoC+Npv/tQah5D6hsB2fBeJOrv4WA
v9iq9q/TNtdVVp4wzmUTz/tL2aLMeINT0TS/pxGfDML0LPUnkXrMTRxpuyMs
FwFCKhwkSlfJwnUYVuNBmUQyofF/GCGLMpn2VsKTczPKQHtJCiMCiwxHBHPV
SxfztHhS8QWJBxWxkcQxnHsHhQG5NPIizcLMVoNuqg+oZAm1qP2rj9XCc2ja
CV5rrBF94ODRFtMEqoeAXv1jsjSacUv0sZBD3hdljPmapzUipuSZRRIF/J10
5HEkULbpdcUa14QvkJ5DLTR+0z3c+Xz27AIa6y+wRxlFwhzFlOdyT+bcjWni
KY29haatexbzVAYY1LHucd9jwD56HY/N+UnppovvoFXPile6xhvjw6nS21Bt
FXj2k8rwhm3i0PiCGzzQtsufRl/Nlt5aDatNKlbSSilFfetSUrVziPBnpq7m
+L/7kLcNYfcSXvjjBS5fV6NVc+8tE1r/9g29XgMdF4uVSU0bTHldZF9WwcEv
aQAk7U2GySZnghCxDxMAWpMhK3+YVl2/JWiy9zbssFiDVBuK1jbgHQWdpwjK
BjP7pfHI+FmmVi0b2xlfSofMDSIsqWiXpsTqRbozVuFg0cZUFxvc85Nmprod
Gr+6EPurtKXxYzsVR2G3Frltu6EJc8PJj+o9Y5PM4r73d51fUWvD8WouBOyI
KD6dug/pTyRh0zRVrlr+K68QOd90b18esyOeCK04YO2JfQUdFqpRSkWyO896
qnNhR9dNizqMw2TzctGSdNwNWNTejq3/ZkjLCNhPPKPC5PZ/w74MNl0GNvxe
UjM6seCEiDIoeGQVu7OX4XUTVokhLmoQC9yJzgowRTDSqU30NXlHnJjQCEKk
JvhI3y8rk19bulXxfOyRJEfnXjcvGfaZupkNHIDixV2Mdvq+fUsNgpbmJXlO
NpeOjLc9NTODYcLXsaDy/0p0QWoi27TWSqy3mGW9SO6wFH/+FTSdbX19F/Eb
aHUlifwzQ24N9FNszPF78YQzTTJ7RBiDda36ZBoguQ8QUXi5mK3ppRZj1rtR
1E8Q5IG32bLnxVPLOx0VJONQh7Rt4iWr4+qrmAhhNQAOflZ0yPd9xm2wdqtc
l7wAHbhCX8lTQlgDZ2qISHzCyEL89gfOo3A7PmfHMcKrtsdAWwCyckGsDe/7
ARCaxRkLfGD21vE1hqX7kqmb9zkfbQzjL4lRzPbCBUkY4/DNFGkl+FQtaZp7
vZTQLtsDOoEXTZIuUTpwV6NIqxTS31Cxub93YTI34JX9GXMG4vQ1WJGxz5Ep
HggHt/8t+rwkShbB0Jjw5Xh4DWaZp9n7wmnM20yZ9CKb3XrHLfSorn9dCjVC
ng1S02y4zL+XRSi7PriE5u2eUnx/Eo8tkiBGaESspCDd+BTvA4Tb4DI7/xaz
XhXERrRmfxgcuZlArrqgv86yhAjMSVGYnwaz/dnOAiHe8OAwJaa6+4ZxXA8a
frXQsso6KAezUtWdBUG2EagoRb4MfbOeIVtjgtvltQNQfQJoNSI0smH7kpES
BTQ5z5mobAiWxFKn3IRUy7autnqcztuyfOjg9kXI/8hGmmf+L5RmKiVP2kxX
Z3b0lUGA8uPsKXn748IVUnD15k6vSYDiylyTv4tX1UIg9sDjaf9e/E6L5wul
E7BLnUOVb58qu07k8bd33ZCl4fEcIPumo72gLy1YQKw/aHXV/UNwdGnWUUXI
/Db2Y2rsluA7EE2XywTz21z1yWCAirLY0u5BcjdC2as+T85OK+GBLOvx0tjg
003uqybCsZgksZjgXpq921B4aX/AexnAutJdUbcSG6OCtyMGdXYyKeFLDCeU
HxFflVtina8yksGT//0voRsjyJkWdKyH98CaiLPCJHrbk/Hbq7m4XD1joU3+
i5TJ+vNX5zfwP0dmO7lBK7OJT1XfZQmfvQ37+X9HvnviFE36IB4gD/fZ+VZc
Ra8u1ubRP4UTo2wTeUFOf7QwYEJXst1SO/saWfhDWJDDK7RNnuaM8UgKIrfW
KOKPgaYW/G6Z8/iCZUz1j3alhhOAlDtO6PJ2PO8Sfy0nBptP71cm8YPBzjqd
MRp0NO5es2+cHZnYDJoqoVsgzVwa4udzo0EASRPC7Hzp7DE+owwfy+h0bRU4
s4uh2v0JmsyXgygXI7JyKl8jYUUG/ZwP1XX1kefn+zvaiadHMXwX5yGWEmve
ii4gF4VP0FDhQF/+uT5wSxhwAt2ZZ5qzaOZCOT4F0VSYmMRQjcM+9xAxLa1c
dlfNTD3rKcnrCsd3ZHTJCSFRHGx71dR8cdrMHphd4uu7xmDIy/riLlt3ra1g
t6l3XjS1QiqmdGGmEGBlu6VBCC9Tc80kcqFoAcQ5Y/aWgrSXtISI74Mkihrt
EbctAnck+NfeYJ/5GOqhkMla2SwfAh+bfjB3I9PpAkZTYdIMWzbE6fk/YGYv
RbKqGerNi90eVrmZB0/sKcL1uET+P2ZzMw6RbLSyXYAwCfR6HRrwHQFkJdU5
knxVTXPcUXylWOvqEf6Vn+i0qepfmmvLQG1s8DgJmzaLfCEvXl+3Ak1bOJxM
S75viIPwsTYj7gdYZtfJ+prVbC8ZHAob9bIAxr03Rs5no5xlcrf1lU5Ta+CZ
BVnYLifEY2Smf+D49OncV9tci8JyUn7us/mREbDvWzljL4QSs7LhLLdldsW3
5dRJDjEn2nelmnoAzT5X8VPWxD6sQHjfedOrzaE8XT37/l4+sE3csuNIJGPE
1psOHk28rblrBYt7vwHCqyCqx2vXhf81oT24G0kUprz2f/f79wM8QX+RtAQx
3gmBbwlGKpvR0iaiIFL7XS85f7cSmhUqKvdrY5j2Be77b5TdL5CUCZy/THIX
Jov0gEVNM9MpZ2kXcoSVyzUJxZDm3sMLkKYjlERpkTx9v1QEAwGlzu8+hhYI
zJFwlQaUjTanVv3R/W1o4aDP+GxOB6HSnk8b66WeHU8nYQN8uiFu8GKGPD0z
9AO1je0XQXetADYKcx61HZ5mjoBAl7XDeEpl/X3GhuD4/vTfn3hdTV1G15Xi
Cgt5JP5flBBC/oOIc8ouIj/eI4TQnkSAHNhMRH5uh0hZO2LnovixuraPw4hO
zga4TUkizQe/4zd6gxkUendU95F6y/0O0Vuh/32dnwFODlm8evEV+k2WQRgb
c9uaIj/2+VieNmtKOBbMhsWR03roJbDCQreXd2KSlaHOjJ16LGz/HjburiVj
BpyVTbQZw03WcXeg5BVhDt85mS3pIgKsilR1LU3EKo5BIw+gpLJ/OyeSjFs1
7fLWkJDVG5sJliksws2A9m9kFhSPZg7jXULaUVaIi4sVvqv5pKPrDOf8B7WR
iBRxKqvESiXIFoC4Q11RTQJiGTC8JruB/PBu/oG/O9NzGMdyppidF07KihOJ
1M9VanYfnRT98xvnoTfBkBV4sZn9dCYS2T0lsk+ob8Syq2pQrCRTociX8bfR
5kSh2ao9zuLfXzbYTDChOFml7NqeZQWL6mydooGoh3BLeh0Mg18jNkBXHdDN
R7tSHWZwWulNQKNncvTJkWONuIXBlCOWSvuLVSFw/4BpgIaUd/aEx9EHqRi2
LPIKoXyBS0jHhalhiqXkw2/4MTT+xMA9+leaCALS4GeNkx3ni4JoTzVD9I7z
lvYG8PSjqvrtH2yhDzHSGpim3jtaukdKoCLHmigU/CW/eKMXdU/sQatqwGfC
GwIO20c9FTaXL3Z8R7Y0q16wW7rwPIPnHZsCoHGBCCfH6GpuuPsdixFwya/w
/90PVWjN+Nqf4zSJBjJ3VNPoxpaBopQHs6iqEgb7FNGeib+jl/lIxfiAlGkb
2mkdGCiSrpRUKa+jfVgId/cm7uP6JnPL9rJPbdJ4iIOqo122sxFu2PyKmuaI
q+gFdnBNvX25o4GGFJN+9Zv6e+a89DASjZNCZLbuHBbYovTX+3ZYjcX9mAuM
gvpqBl2LFh77GndwUZTJTr7Yc9iF9SdhaydMjGuQDWc+QfPmpj6nZzPuA5NW
/vqXoInET7SAnLQXtnFJfqFhkgv7tS4SQQ0bFWD1cRpE94MZg3B3ahmeIiir
hnQTR5pZ1/LwTBQS3uBSvsnVgrcNz4x9ipbM4XLNCJoKsl4lMiqbhL/MM3Zk
YFWo+LM/DgasDEXkVKgX9DUHhwTbKuBRf5XubshyrAsSbqSNLkQowzxU3J3h
P5iFanRvP1cdEMwk4RlGF7bpf6N+KU8OxosB8p+NipCx6pnxTvfExPSSDjCa
BS9YreBgoB0zYB3uHcztjjqXExX6TcXywus/fN8EovryJCs78w4UEhibfBdq
4TyOzcIL0zU5o+YE7vDW8zJrryL+MmtaIrgttYQGndqx5Zbc9rpoPiIZ2ZK1
G1q7cN2SVKqNaYmzfYXUvgacGihxITxmJx/759D/pGvrsfqeb4i8CUJqJgRa
a+nVFmxDKBEG7Yo4qrXyJoQ6x/Hdmi3ThH1QuUcWufnQBvHimd8GPvVj9lZg
oaFQ0TO6pttrRqjRjf7nVdazSeUrqJ2SJ4X/qRbHVk/hJhPk+ByEiJyYBUJW
lH04NrkJJ/wNpYX8zJ3RDuANAlfglpWTrezUHS8nQxVYJvpDTneAlLGMDoU5
YFqz93GYNdHdrbgNXu216Z/rV57xrfARbQfVdmhwSAp7+sfAlU+eISQGDeRG
q4UF/DMXnd3y85Ti/gD92XCU+LewzbA0aTnEpt61dn//n2gsyoDu7zfotvKs
CRzlmUmLzbVyfWG9s2PMrMvApP73FcR4or6cma2dwn4x4phqkbp3j94UxwGP
0TPpjbzaaO1ve4LakQodGxUphnlX0fgmd6N4qnB1FyXx3dv4i9gbihQ0WNhC
Cw0ynk3UcqkxkYPp0MJxi79lZtbwq6xdx4MIxolUIiwpDtsLUSmVNnVmLG2v
aOD4y89NDog96f7KV5Bqk9DdkJQs3W4kt1wTdYGuNoZ0PnSJCt53UOVhGDmb
PjQbAJZ2duxE9Aq/dZpMzGjknROZExDA7tq1l6uNO80o3kPD5JniUYCyuUfJ
GeyjxVi9SuaUVbBae6psJJJcUwjVMz2UEXN4UN7Ov1Z0H54TzUfudfkmfOq3
pgoxEapYqKmveXUKV5F0I3e5U9Jw9+YrYDSowwkW785eYFGkT7epFYqxXYA/
jgaZFkfS9FFjnT/i5qLZX/SJNUM6B06aoItS/Mf+NFFnjOi4VBQ4ErxVHgZm
skB8PI/RfU+32z1XMZll/zSKnKRc/NBAosIi3vbvzHBVJbW4eUeCAToTzIKE
7e+rWWIAfEMIUZkXYzjVxt/DjV90O1yb1zrkeFua92OVNguoIOWOUCjO7a1l
W4Abb9+s+DmUy/HPh4i352D7hY94JbNOJf9K4RqDlgGoesHBkFs1lIbhJthK
iUk496nikweM+sRxYmtvcNbbbql9h7+s2GXmIG/Nq90iG6gZhd8/tPFnX+sr
ooaOPbBW8yfOvSKOD7b+mZltGQXiMsineQ8H8u+S10PCPzUae34R1hQZdHdO
xRngTcerXohiBEHL61NZVmmIQo2OJljjAcGytTHT0VZl4D81RCQbpcCSXw2O
pixzpxgcaOJPVuVV5oQtDbnliQlwmirBK7YaFlHMHNoMDUvD5Ek+/R3YPgqI
QRbkzFMwkTSFoLxMNT5xVw6vP0rui+oIAowq3gyZ+JZ1BzPMy3tOBwYT37jx
BkVLQRCVTD1pXWsyJYpKX2w1Py2Ou8b9diVSWj3T1ADnYExQ8suDs5vGo9Ee
+1TzRY4laszwBE875kG/nVP5a7fkS/WV6RwKoXkaY6sPqYe9JY2nSuk8JbnD
4YmktdKx3fadlg266Jk0Fftm2ofYDYPmamWLlPoWwKxQTYervj1b3HQGLao3
ezLdlwUoSWfX2XqgZ+SO1oPJGweNxl3U4raME6iDAWq+CCohVL3SEY2iLNeG
0gdiOxYPQdZNuTik2c5AXcvoJ+m0Vc/gegm1YPOJh8prz6BoBYkYzISdWF4M
7pR0cuFVJL+zntcGX9WVlemZo6vjEFX6N7FPJQo57y2fa9TyqrCk7lMKjPkU
tY5RcTh+b21Ikf+bWWNXEIxlvp6bMv+oL2bUwV+gfgGCJEmFWO0rXfmgMgit
RK4W3ZBBkGH3sV/X4AGFHMzrJDYvBH4rFcb6cnTRj5LFwsSg5PFo7tnCvhrZ
MeYEcllwGvuh51zks1JulC9f+Uno6B+dos60Ir0D1/2yIrG0d4mt9gyH1GBl
TzfWSW5Rz6xL/tivXq/YADnCZRmxp4wE4VPJzSDenZpXz/VqcLtoGi00Folm
aEW8jJnQntFWnAq8BYseIQAYl31wPLVLW1O4HepjaY47IoOITpZRJ5ChGFJC
09nQJJ4r6f6wb6C1Y2gnWl2XMNcb8WPqwF9sMqkfEe3Y+g3zDqCB/ZQblT9r
Xt23P1xWYLgB/aTsaDhEb7maju0q3Q9DTMUzqAP7PNexXLFZgGwV3t+gy8Lo
5P93qLWK4Lk2CCPbpro2HR+DAFQki8N4Lkt0e/C4KE7dcGb09n9q/EhBVKfJ
yV27F/AB9W8eI1EYY9yUsU5Dc4wCC1QACcE/xMYFMZyXXghudzXzv3yiIrcs
34MCw6avlR5HzRN448cX6l89REzmEVbrrBDgR32BPYm/QKralm5/syNLQUki
vAnDXW3yx3vKj7dCTWSNY+2NCdQ6WHsx2HuYk87hKy4WQwU0YgGif66iVYhd
M79NXFqY5P+8U8xFtCy/RjBEa5mo8DJqbSr6dgwoO1jCaAiC/+kuIa7SXtIn
A0QvqR/460FkL8HQ50wA6jZROJjpmPgMyHfwUcYYlHiZ4+O2vLKaeuJf2iV/
MvE0NTFj85gSH7sHPNfWeqJ9cFPep9/i8kGPLBjxDknF2wwzRWOH3W5n1/Z7
Avc46W0K7iV5LROS2xTqYrG2hPxeaa+l2LKVClvz4bI+4odigu+kME5u6vna
SjteVgfI/1ZaciKtbJEGYk4V19HGWC8mnXA0y77ZQlX1Szb3C764Bqx6OfLz
62bGSZAIhWFAtaaVt0yRraMcac/2f3wYNxYYDtnMR/Cpb1rCId3pGUwuCwvH
SNflouhw9trBSC3NwRBdfNqRILrYwV2bN5JiXRGRomNXkXLBkVRUdrTZ3Jw9
4rzdEBMwI8rYuqZCuqndqzouoY5LPDgSrIRssgiel64/oviKF9NjSjvDTrSc
SuQzb2ybiNmUniH3SxegMaOe5L6X8RIHtgQvwPG9kwekfeQ8T3vw0u1Hh9V/
VVNkiPwE5KtD01X7/TYGu8tyUQU4cES/RqNE05eASkEM9/h/oe7R3b5Pu5L+
Rj4MAIZ7tv9DtZ6RdKp0SaZXM272aEHfhiExM5xpENAoTnGsT7RI5B7ULHQI
YhUnpMgzYxd/UM8Z2gVSM7h/Mns0kgjCBN4sDqRCHnj9E9MYJ7Ih6OB8eJSr
bUaDi978O+W7lAzRKiGElfzbKKxGpvzTMbYQuWMU+M9rZ6FpUp1fh8u9jP6g
CQTyvqGwxmCAPkvoukJof+z9pAV3w2xanUovVNax32fRco1BY6Gizo1vXF5a
qeVHMnCRoHNszfMIZSV7LX9YISFlMSfmGj2u5Q4YQ2rj3Eba1RqhrTWM9r1m
RIVFpG8sp1hwDFZU/pPzYEW6q8bSL5R1i4dP1J9OexXBEnre0yDCCX79FsQE
uZpQ0pNvWz/pNX15tTq0uwY+KE0y2FQ6DEhbvjSia6bXI70txSSaLFo0yIGU
ZSaMvp0IGgtXic+4j9QXkHbpwn1kH8ygj++jg0dadbhYNVdLjmVoO7LdCr0s
lD8DML9ahCUyaao/RvlCrwrymIRxwQjTqleHsHl3xqbYUUcqWk2egpfKIEZo
YBRkwytZHsTAuj6ZibdZfobpx+/3GNwnqQ/EijsL1xso3z7SbV5Y/HE+W/wx
K9PgC1rSpNZRjdfjkL1+XewQiz/x4L7rXyeaoIRR3hQpxD/EH5niB+PyTFdw
6tTkShleyhHXfOBAAuUjR7EecMjz4ZDzABvLEs1PXB0AxmBqGf9M0HNHYefA
ojPiDMttBiw30bOk6DEEHDBmQr4Uhr+0ZpuPHles2WtLSKTXTqQivde76Bll
O41x8zFVSVY5M1+319xUhlPI7XgmAHcAFeNqDgsm9f/hhODIjBXB04uNdJ7Z
EOSeWywGoi71+obm7DBXuBtRS73rV3lf5r+UicYz5I/ZceMySvObpr9qJ9cs
vhe1RfwUq8vWqWnqJVF6Hx8MawWfdvcyvdWqejhLgh5kapRF96ssfxEs4c0l
sE5ovdC9BtZ/eD7QkvSikLEaD9Y2x4O9KebvV9iEvE1nBYT1HXnvnOWzHvcm
xOIdtT1TC3EnIqaFeMX+xUd22v7VtGiku59Y7+bBoG4GGNt8HW1CmyK+/r1Y
AAE2SLYsvcOgB9st4wKjbczIx9rjrxzGcKP0qbaBSyy6wpx8r4iO1nZ2QLQj
ArLVlJsM44xhV8VoQ1X1zG/unOdM49jqBvCAKDagfATcOab7SWtrC/3fP0hs
oGCHtRtSuI73bi4H+Zz735vXC3SRuKfKoHC2lGxdmyiKb7upefpcIont+/Em
exIIIPQMakonwyIbIgE+EDImAKtn3JEK61f39ytj2AUhc9KCTaEFbKzxTcKe
QhqnEurcmCcr3Y71lIrKOxTYWmvhGudLXiNy5W1/919CnjdPfUgXri/2JEWc
LLN3Bh0sj2LnUZXlvOEIgHUbh5BVWWIsMxmikgCt1vEgy5WguCcqZEqEAe1q
ReXaAP4iaJfCKbDJvoge7f2Csp6onTNMmT7a1iFtoTH6UWKddec1ClVfi15M
z2ORQ0oNt7IsUHyG3Wk620HB/39YBCjH8nW8IGvv035MkD5Eu5rrIB01TINw
Ok6y95ADeLJ83ZmPRKe6ursSDrTSHQzqpTDMd3VpoHS6kS1dq5vRbjeh1G/F
QQKC0GsNbheqQm2o6VsIJfIzLNvhLgvV3WnUb9aHRX5AedEC1kBtuJ5WT3eW
hK/OjJk2oK5NWPRQgtrKP6rlwviaoyoicvztTpQZT0uDTCpFO1l8oqtHpcrU
RP8DZX4TnfB5FJLWEW/v6r5fux9XKx7i/u+kn5XZ6BMg0dsiCZO97kVWDV+H
vGdQV7UiublC4hBIzxulK3Qh09VVqVc2Y4EF2EwxccZBVgQbUR/wv6rdfV7G
MUC2YSd21l76V610gj6yxmmreAgpHRBT1G7RCsCzf/6zm/V6ODG2Qv2Pl0lC
aPtfTNDjsXdS4brmkMY2HIVj529CD89cSSUBdaR2OgT52ZjzqyhqVxbzm6bZ
sU3+GMqCdA8a3wKNVfDSAG3ZDC6WN2H9SVwf3LuUKGr6zfUGVJ9s/awx0oB0
+0MahKfHR9T2wu7I/IXlw/pJR6oNsl0qiJdKwBtPh1tEUh/+WbkZ8fGmxTL3
0rzGttcxnHSuZOsE7CGkVPnY7DcCoSgEAFmIb86/Fw1iRUU7hCqxMvMkgYy/
4OGjjtErGoVUENfS0IuXmI/EV8GdbkdscQDJ3KUm5/1k3FkE7lfdb3tGzUIp
zSuqqnoF/IffB52OM7yBFWZjrX95cK7DA7ydTWne3b402Sxz0Rmfb/DhtE+w
nWVK73q/Siz8Vh4sE3K0orcTt6gi2WQoA9LmeOkpUZdMQFBJ/itmNi4hUhaM
vobQHinxf6vtY1ZrR16jVNMAjGEZiJUZEMSQDJWTXYOSUsBO+Tx6bhQWZBxA
aKJ7RyVB18cHI3x/0I154MqpjpBp6G1DQWhaquED3wSdAJKjhjrkpHFwHZU+
9mfT9qKrQBGJjpDgUNmME1AR/H65fzUT3HIEI+/isDjwsB3XpkciEBeA/fUF
mscmOZ6IgpcHtifnirJXIRxOE73Vu7NodLrtfkEKR1DN1aNOIsyEIkqcx1D4
xRMKl4tyxzCPjQG505iUe6I5kk3s5HDEVVNiuwqaA1RRLUneIV8cTERyyWrG
N9Nt+OyV55T/94UoF+fuguhraBk0qHRtzJ6j4nO2ZvwrGmgpSmw+JheGcuUe
HxgGSQaZeAUNxMO3ig8QrP39lEf012L0m/dRQTphjrGOdXO/W8Rky13TpDXb
blvZQJqty3hgzWHkxxaiPxB2iHRURrAeJlG2WpRsIAa62LkH9ppBJY424AGy
IjgCum1aMdciYKNeZJcWjmbqI1cpRizhSrui+eQeqrLWlfCdXzK/oJgFABNg
LUAyhM647ml88LgbED68tA/z8GVtH9yOf7/+A6n4grQk/f/C3vxHBn0EIGkl
p3d+BmSOvJu4B7kIDRzLbK8a+rZWFGL8PU3HYgaAhllymAPluursa0VqrBEe
sOhG9OMOBBU8YsWoIMvnbzlzUXZzQxlR1oXUy8It7u9+ugBCTDQ6qknHr91j
02E/UEo5c3+ibUm3aaDdYjf6oRuQQAPp37zDCFfypdNO+xsohGF95DHqByaW
CCQjYKmVnBPE1DM1+ZGhtXlxA+bmQGJd2v1Tr9P0YemfNEDm5PcKRX1Wo91f
XbSnV9opXZYuwquKBQ7kVLB0Vq/fnDWIeTKuNaTfjPNyNQQgw+ju8gVsPGLz
uHmbKrA1MIGOekQMOgydIgn6pNi52d0mFA60E8WUvW0qVVhaoJKjvphkrdk8
+gymyJamQaJPN0hvk02SN9s0W5xxm1hw0ZKvDIAG2wOti5T7IY5cjHc024+l
iZdqLR66Kz2D5c4FBaSIPB+SHMRmdQE46hzKDlJbMjg3rYdCxgLOZiVTGVv5
BwfqfovCU/t/IKcQXxmJWkSIRkNyLVUHuSsJC6DSrfi3CwT/tWNtzq15dVOS
qKyLAqhz8kj6cNXA7Ksg2MOer/S4+T1MuNPyGBc7FF6vW1mZbHC2ihCBjgD3
4hdaLl0orNd6Fr6betHp3isLc6OAdBqBcKo4U60Kr8vpDdtJtx6S9d/6rMP8
wfTuowJtuCuOc1UFY8IMOqDOQIskL/i0ayBFubAcT0rImlBrwYF0PSPwBfc/
JT7OjPidJsBvBCdVWgRpFLvjT4c1bDmFLn0LY8B3nhfLRaZHCapGxIUCsRYV
ENTf/VhZei/7IYembJ/kNptzyBSSgr3cFmygo95fEslC5w7NebC1BQZJzskp
ZP8cgLE4Jo1Z/vn4U7rRfDq3fy5/ZE4gSX7FiGfl3ebFEKjxZecxeC0beNyC
yPjoG5hMjBgpUioICrQjduCnlCyoI1aF1qHorXYZ4JBpEPq6wkTobH592iEp
lFoQ2kJZTWmTSkRTdgF5vOMRG2NzWLMM7KdRzmFxGtAeonkNdfuoTNuXjNyx
dqFzYWRAyEm6fEkSTajr2KbEWtP0meEXIMOfSOka0vWn1Rszgx0QJfxZi4ov
o+xB/k5g3JqRtghZr2/tO+SyrpoZ+wxgShr7qLhU20njO6bOwvPp6g0UprTU
JVfvsj67g8VmOu6gMNA+F6ndWWI5YBPgttzcOucJ4bUJt2hmkcmyBTm5T27W
1Nf2u37mstdujt+2J3gBJf1fDP6e1Zj4C0fmFm8yPC11pIpM/sbbcddIu780
crO57Jkf039QN5N3l2PucoxzAHY7Kn3z1QgvtRGyZrRUuNo37FyFpmodNL8z
+YpR+43bd7iO17wtex7QEoN6FwgK3rMEBZYkuI/EYMNhNijGyoiYg485JetG
PVjr+8IfjD1mdhGh9jsz6JFskvnHOx5Ywjxxl/T7Dp8iAxKrEJ+RhWlh+Uqt
MPbha2np4xbSHC/6U+0lxKzbmvJXU7iu+ueqCvODSeUDD75LA2VzkSZamea5
nquz8KxkZBPhGY4fe1myH8yULu7LlDrAt+C3/3uRKBFoi1/1tFiPdmHcghgX
MZ/+qtJs4x6slQ0nbR6oZhv/vZYXGeVwqubV/n7QPoLDoIa6WkbB0lmU5OGn
LNf+8gwc2l3ynbbP7Bz+jvvDOtLrXbltjTcPbCr481knIm3Qo6AM6dZ647gF
CijUYMGpz8iVAuVQ18kSrAEZuaGYB34mjvcpm2TrbTOm6PArhruIulMpiIpE
OcOGAsX0l673Xt4HvGiUnHD2eh/0oLtM71rFgXsed7s/qsSJlWKI4aQmOe73
eGhqTnqEkp/MO1ZgwNMuVqUIw3EcRyzxS9ZsmwMyKvdu8P0VbjIIc1J2Nnga
sIY1YYch3ReHv7t82WgVGbl34qrqQKVk+HzQt0B2pra+iGt/vDbfnZ1y3Mty
J10D/qkh6v1emOCa5WSmLcKHdOUOZkNQW6+7Wjy63NufucwghkJstGrUGXdr
qOqwO8LnjuJuB7yszNcS5wLTfJQpdHjbjdWfiZIqQppHbnEMr/fIYOcj5SiT
TXegkLz9XxeZCBs4lB5pd1NcxvQvje8Y6bon3XYd5io7ApKHUVzFGtBm6sdq
jkaNevxqaiiyKwtekDLVIPjbo/S6nEeR8mm5iNPF7EgaQ6V+555jHLfsFqwK
csQyfV6GqgN0WwCDJ1ckNuOMpGsZprL/yef4oNVtcOmaoxwYmIAHK0I+u9yq
g69L8aJublAH/LB218on6hbpnTtcl5zO3mNCCCtc4aw8Knlci7zVp3ZreiOs
nvFNrJCNT6C4TgcNOHcXW9mdCbQ+FnAN/LHkp0/xIgLAHvbky8PUX2dzAv0U
xednOp9rrS1rbkE9YLw6KiE+UwNnw3B/N7gF+IC4g2xO8bsSOPjgrZOOvkjX
u8K0PwHUQGZm+jo+4VMEMx1kai23PwNABCXqh/Ornr9smTPH8SrVR/VtqnCp
hPnFsV/8CFSTCOMWvTQ+DbL8fbDVU1PvRJzFmuHljetCONy4R1bN24ARE85x
2iNpLIY3jypEKwlL+XI0qUgjx6P5SsN0vJ/JWRgvxuSOVRMQYCMezIzOZ8+K
/JJ2X+v3OllHU3pTLm382vYpCFV1GzjS9GHWnwLkFAAatsQLo3NBZsc3wz8+
pTPHWCuLPcZBpBvgbcq42hz9BKI0xhmvMrddtRN/N1SRAR2Iv5Dw4ZAPfCkW
zCbt4ufn+Lpp2QLn8nHCqdmAy/3GDuNoD8GAq4W9x8axHJqoM60e2U3PrpcV
wA1po8mZOBZ20q+5nZLTEPRUagv8E5gx0g11V+2Bakb+i+MaVjN9CME3jQtZ
oSvhjG90Y5yywsIfUS8KPY1YVyo60UXbVG+YRxW4FOzwb0qiy1zDuj0Afdb5
p6hsPMILIq2aXjC0sysJfiJNkmFHAQ3CN9SXs5ofPRhF8aDqwUCugE7D9PFh
pWi0TN5m+YMxQ8HApFysDFyy5TiEEKv0KsmKJEwctl7LUeZUmR0ylWFUe/dl
KTd9iYHxQgflkOCH6Vhx3fpL7IAFrdW6+tr8myWLw/d8XE7GJ4qWUnepbiuA
01qj8qPRPGl5EtxhbDtwPu8OOntRou/fmAwmVeMbprWZogeLJ7/gWVy9jBTl
rqHYteRP2UX36+gxSn3RSdghrfXkgv11ZHPNn1mHmSmvkWOq/b1MrsFWS2J3
4GjyhvN+PzutE2tdjEB4AvuwjLiDtlMyv5/+Miz5fdcu+M4YS6YSYpa0Fw8B
b8MUred9ghjZvQ5axj2wLc44EznDaIQZXCXKv3vjgUgKjaGhgKVJgiS9Zf/7
enJ1VyoZ/T8o/OZchp5hCOrVgr6pPRbal9irgncK/wC0Byz/FgHwBmai6XsK
KG5cjRh3h/oC3bbxARacZtGrK5EuMtiVOpfgD/KDSywrYQUvAL7b4ghw/pZz
vgBLph2854teUlnvTwUkE4rfxm3w37TAoja0bNVK7mzHcCNjB9IdSvQQOPmn
otnp3N1GyrmSvMBfOSI/GpJ+ZHqiAAvZp2lPSGF8RrG5vldUDDNOV90edAfi
Vlrsr8iloYdc5qXF+AuMfKuUDy2RjDdzh5aE8LiYkqfLSlnNMoCU+iFJL2yT
ZCBjW7XvBM5QKV7S/9Uhn7rDJO4Z672jB2Hm8ot3GA3sqapGaIF5lCm+nv/i
SKKTDv7x2gL0VHzTjJzgNITWGn07tnSCkLLXHo5r6cMPwMPD7poYZ24BQMa5
lBUTInKwzNLiPOB+WvDhA7i9WbcF4P8unUIhOnmkkb66NN7sFk185i0SpitH
ExYphE1BzBVnlIvizkXcMxLd0Hse7msTQ2BeIShl/6jCxpnFG/jipQtwjJxn
tjCsi+mHSYkuwWHdlD6Q9mkaHnBtB3TXGmb2yHzyXvVX6qxesjzO523pPMBj
/UTYysv5MpTMe+S7W42k/bK+kYiPwmZFRwtw/E3J0tJsab/mORxwBdaEYcRq
Z9dGkLO1Sz256xn8A3FjbOL94uont+UyJnFllOqAP+0KJMgI5Y9n4MYSuRuC
/wfqXj97+6V97J6evZr1DHZz0TEdSZV2eqFHFAlQa3CRjBOzvqTGr2Cp3MYa
jPNWqCg7KUXjajBP/fype5E19qYA8J7f6/5msj/UkkWjiRc29gdJkgOSXNRd
zzLXp9CmA/ZzRNrXMoa+NuOApu9JKlBwrnIlRSg8eG7t5+aaKiRsIOXA5uHP
rk8+2qexpj1yCp/aKWn8GkYSwxx+b6v+m5n17gFqwf979pVpVB6cj0p7A8+i
LcSFy73cdMS18Q6Bcgz0N4jxLRy/mNnI63e5M75epFBAyGNQyrHID9pRFu0v
fyezmODMcVhm1vc2Joyx+jrQr8ieDoiEFit7eSnu17LrSQtDM0SZ/YFCMUOo
Gq9jmS9gQBI7dUE7ke1F2uuhovI1iSloL3xDwGc0Yxx3iURKjp+2cnfhGubd
8o3Gi7Eo2bGRVuqb5XwVkNbMGn3646ZmGqqpL0Eodt9dG4Ll+k1pJWXhd/Zq
Lr5TXq+WItcVvnQCWf3FBWBKpYkFU9vhNXddNv3uzWQmomdiLlJm7peLax8A
So1mrr6gN77nVz20IHGNIvOwW83VWku99gyhwpL64vIyF8uCiCJ1BPqpdh1F
bR2L7yFNlcqPOfZNi6UdOFDyF56S9I5uziscT6cRhWA6PHno5iy+tDAi8zGF
mv6651HfMR46wpbYNbnQ4eAA4CXICs9UD+GNOqvC/VqLky8Ju2Yde3pxflsp
cNSk26CkaI5MKJJ6WpRIrXsyj8R6d1hkS0G4oKVlEP0SYOAsqyNuX+kftvec
V5gwDNtWMp+yuN+aQjVv6Y0KrzQXy94CZYRXjEDYmksD30npK1FfgeTOA4IP
mgbb6KuRdRHOtwRjNeXSrb6bnGq4gjSiCOH+Si49LoWEuXnZrZa4TS3IQHdy
8H8Ne6RDzvATcg5MhQhWs+lZmxyZz3eLB7t6KJfokXcerna9F8AAAyImMK5j
j5bJJu01Y/B5LK+tgfuSLzWXFcqZvvoBFk0IxLbH880pT9nSlxGbjJ+ptnsv
850gl2pO15OIQk3CPsPeWD4fD7amGNeIlxh+yMgrVWyBQYposIt9Uc7PyeR0
uo+ZCTCC5Zo6kNEhcpG6utnRlt0SjRIcVn5PmoX34j/6AcNIojOQtNpIL6B1
KGDFVqTtbPmyA5kvu+YTiBhzLw8SRrcPzbj2o4Zla3/bLM+fVSjQhqAowNHh
a6lBSkJ8VPYn8AeGh5YzAiPXaL3VmFFnobQ+X0KVKtsoEOmXVyy9ZlqWt/ki
DgZtaZ7MD1CNpd5DBAYUET0InRuKze6vJladzXPdE/fSZs/cDD0xNq6+MbR3
Zh1mTng2Q0dm3S7e1tFUJcVK9FgxXXFVsyNLxo22Q8VtYzI0M4bOUYg6uM+d
PTJiGV03q+nQMPcmNYXtHuZAF4qIs5b7ychxaZS2HjAQlDLz4mPPQqnBz5tr
+qZ0X+UuxLbeCky+BfPkEjXiriTKqiC8cLkS147r99avD2oC4TMr+TNSpvem
VEXcpChEhK6iPip11qiFqemjDkaCG971beDmoK3dyoQ5KzCjs1wz8QxAxwdA
ocSlehEI7uBXO0S9rrXU4dzEYtJNN0OShWkAsU7XoJWN1uszjSsVIgYNav7Q
AWoPuodLdJOvUOkCtbA5HYBDpQEstjKRTTfPZ8bersEZvz73Osy58jRj68x7
KL1rxE7sYLU0qCn8ZnhGoFXT+nXHJHrRWM0TE6XY0V4pHH0Sez7LfPiLOIUB
7bT9QhDSAGry/MoOdwlE6lAZ6X83Mu1a+i6exRuqY0lLDEfzwtldRdFqalNv
CCJDTRSLGSnC1wxHkaNQVXU+b1IFzM5awXExNtwcgSStaQiF2kxThfcxsR4y
+K8cploKoTdaHVL7UwgcOeh6bTYhszfq25Ohc5n+FZQjXlEmgpHMca5pQlpK
IZznax/qMAPQk/Fvc47yHrnoIjkJ/9/y7u+M290jOnHqCXbvt2EPjZvVYgBx
82F0cnxbS4v+yrfqMqA6lRjdWQGDgd8009pbcs0LXiVx/f7UpENmRXsLd/ja
BdNnUNLwSrjEQiz0QnMZjkh34RZAM9FAW80MDuWOJlaX8ndrTorpvDPy46Vf
2EW2JqdVFhPq6zFxsBGZBoZ23RIgKTcseQwYQJeAGfn1vgQVNrdrVD+c00w/
i2EME9mKVWEn27GAQ55oRBKD+o2GnQqIhJMD8EsuxyHWAymKWyJUmR+FlPo/
pNs2LPuHTG57n8YRqeRzaO3d0J22OrrqiEA4HEb07gCft4jQf9JWzLoLruuG
+mAlNp3zrjXt6uRXw0msPYiaBpSVHmB/M7qs2jEJpOZguwSYTp/+70Topw40
XUFIS5VX0ogxbmIMn8EgYdAH2hwrx6luUSu8FWNUJKaxDUJIe6viM9Gk/LRn
JjFnPHIgVa+VKntJd3PPFQV2QSOveZmxP2qhCrZzWPvbklSKuZ+oqahhhf6K
IboucgnAxIcZW2OuOe41Dyc3xwlk+hRFHmwTf/KkiJ7vQ52Y2g2WZrs9bIBF
G7LHKzCOucDfdQaU5jvy0NZS+6nTbClBKeBnl5djQwma0qQCHmo2l01bAwnI
rOBlcL3y2KNE33Y0bOr7z7V+nzRnfIU4fQnPc2NJoUEZJ4vyhD/u+yuhp07u
hgKnYAwH9Um/AExFBAszMaULd1+Apar5CA+j922KnjY8W0FFwFQJHUvF1+xy
C5Bq2jk/e+UxG+HP8qoF04yhCfHbr6jafbaKkwZ/L2XU3Un9W0yagxUJSKK4
21qUGDGl45lzFXbyeUrMBJMGmLCzOwGLMHTHWStJldShKYC73zQhFg5K01JB
zjUX1GrPqtJqvV7J3Nd2f61dVtIPoyHRkcv9kcfuWgLWDB698dsHWOoq3MZw
fDcdUrIGNmp6YL2Xe66+VqjvQrUqrxruzFxbNI4j7m7V2UWxfiM26kXdAF7p
QnQGRLTxdS7295VNW43nnkAnRnZaHJd2UKUgl+LpBGo5uqPNVpfQrfRlyb9y
kmmXWTHKlObkdx3y12Jy33T5isgsYsnwNkOHnNSGDmEXNa7A0wJadmEySDZr
xtEwFkhKQQMn4kpEaM5CFLnQXRZMTHpEzYOAhjFi+iWhz/UDQdVxOSb5KiVN
OW3L15YrJB1402wTtzDbLEs/vn2rbeIMFmWWrpApjYgpSChuGzC/MT3nDIbD
ppX9OByDDsnMvAZjGwDVfmo2T9Lb/TF3uCVvoeqq34/vDbZNR4IoWsME2fnL
nrNRDNlHnXFGWUBfCSA21nr0XXlLF586Pkz/uCUNL5St4l5V7krPWPV09+aG
95bVltWP7U3owgBgfjI1rFcDJukh2gFJN42zkoM2Fh8SSAa4z7WYYnKJl5gz
vuC6KnlqU0WoJs2gwnQl7hEJKnqquIFlhDJ5NSAhktXOW7qIt1hkvPE89KXX
SrWC35x16b+FKd1BR/DwWoIlLJct4NpK0z7oCw/ooyI4i6bZF7d2UL344tRZ
F0hZVgdv3/yHsmxhBeMwa1M+8l2Un16smdPpGjaDZAUwIM9Mh6aXF1hGolt+
Mz2aDGUohIStgIVUIB8x2g+/H3oExe5q7lY4CTNkOv8Unt3Xo/+isCF+yWZC
n8EUhf1ZGkFXXGPQje7e06lETEA+2L9UtxzXgsfpEo2Q+M3aICr0u5a+HsGz
TEW4sgXCeXACDaaFjZZCU/1afEiSLk3swr/P0rPyzv++UfjXWVg1PA3TiBig
BmWFIBZjRldjCrRy4DWj0Di2sIiGxU3x972hQ9nTaAoQoLPpJGIyVgXH2Lif
F3wr6m5Vms0NyExc0h3P34+9hyvUz301y1s6CR63ubdA9W2p1NoF5f4AxOaw
nkAEy31m1zaWTJc+R7VA+rEsNxnwb2XjF6q64BgyQvdwgEo3bmnNirPty39d
g6NEYQljKt1IuYTn5z9VlXn/Mle2ux3PNK8Z6EOLp38MemFNA/ZVpU0dr/UP
wTVZtuAylWSMlrLmPnoIy2s3Tx78eCBdAdgA67YYYRR3Qhp2828qub2USLbo
hhE6zXnL317YbVrzIY18ttEVI1G7NKY3pfh4CliNoOAt3WCVivOJ/d13y64L
Gg8LuVMYm/lKy/LyuD+Xn+BxuiWah/IrGYpyt6+Yy1gEVxMKQRyIEgIiZesq
UdmkG5MGUDkENF0UGT0tc8MjYtqtBCSnIoXyQfoIUs4ZWKUidpkhIVqAY7u4
0s6PZ+LFrUnsEyjAHziZKz9/QhT41XRK6VoDYm/GPX/kbtSswSo2i5WisYS8
OSTiwyjP/b1jKeYSaOOQFQ0qS+w5o2HLQB3S+HoAxgx10z98Jyx9c5V8Qwdj
QLzjidEL9KvvVwQzTjtXUQLgfmBkzeAfH5547qHUBZs2ZOqAfmFzAVft5Wt/
7OOBUpgtKmu/oDidp2c37at4slt7Qv2YdNMmCTgSVSKICFCRgYXyEoiZKOGW
uqH9/fPzgPGG6GkLUGUhy2W5VBA2wpMhQh0moBly/92/eRrfnIKFnUeVLCy0
iSYEmJRZV40Od0V9QwmpNIMBtz67W0ynxwtMG05YtQOrwZpgqbWJGAIuV5Cd
E02+l09+QVEdtJbIAir+cnWhx5OhfoOfBB1qXWKoNLG4+DTryqqKj/GkIDv1
43Q+352lHnUOvojvPOfIgkIazJt7pTigfKZ0w9JmiFXpyTzXUGavIuiNJZ2p
IJ8O6zZT+jHOVg7FztFqwlWJ0kCFAkPOctqnFRaP2TGbREfAHvBB1nLRdVmt
0gPnNhjC0llxdrN8CNw7SfsVe2EmquG3UElzSRLpjw34bo0pJVPdct3RBJ6g
YyvS2dH8dsH63p5rMiRAr2c4eIIYJlUmNAyqGjuw2PfoecDkQwJCZnk7e5IZ
mYPHF1nRGaRH6HyqJZEfSleGV/pUSvY52Nda/SFDRABjloGgBAdSoHz941jo
OiZP784VxbN3swjt52pwI7iq/M6T0BOBbBv9EJFIRruLcy5MzObfIa00OZlI
5eIu8KvLf8Mt9JcTZ3qSrqbYhSKHHqL3WIRbKgvXltpniUISDmdbytfJYh1X
jmUtRCtMMr+1YEZ1ixjlEaTZH5s1Snqi7c1ABkOeWHqY6+QFVMl1BX7RD8Pd
Yz3vcYJOcN37mArzxtlVI8TMJHDihH4FbHTYKH5D9RRhDgNSlqqFKQcSoapZ
bJKhMOqvw8dr/wiBW/A7GYLYjh899xuQqkTInhyCB8qK20bfquVFnvRq71MG
yHIqcM1epT2cwmp2kKElDAYG6hJu/6akNM2A3TTLLHbO+FVFKp2FmV4QXqef
BAHUVYP1IuzgDJFTLe3mhe2mayCYzFrk4zNG0OirrzD6UaADye4YbiMlMToe
ox9ywE7+AVaHAmvROJYsIr87TwM5Mn63JmhZQazjPW9R/DAkYQI0Z7SAb7uU
VeJoGhRHo05OzlNOxGmpKzYd/GTgPdJcBZGYu8HDk287YYGbj5KcxW86riKW
dCOgav13ItjvSeQM+/HzTFvEb9wxm0PUTScYghI8/4G2n9FZTf4tnGNcPzhE
uLffl8Skpv1z+GKG0iZAt2dlraSSehcJ4VzdvD0KVJH3F5uk3YZSHMOT0V3f
f8KNTh03FjBNZnfvUkCVPHPsRm3BT0R66e7GMqPtd8pMGcp2Odb4vJzbhD08
hRejqbzfcyf7ULVGcdBsNNT8Ah0ewHACEDl5h8hVokf2Sd9ZXegXx1rxbV/s
jWHWs1XadpxB+5tyiH87ywpipn3CGSX+2fHt2EToq7LHQnOCJaz8xrtyCF3V
CsNFj5oLsU6kriMSb5z9I+jrWFxepzvMPdpMCdyltCB9zkwQpTlqPU2rJzI0
vzFiwQQLNrKxYe+V6uvzlw5kKTYF9nNXHGQ+fj4EAywmqKh9bKlERM3l/6Zf
aMBGseu7iMIdSZ9Euq+3AVjYhvr3p8rHy+0Kpj5/zlHrVZM7Sp7/3LDF9oKX
1BLVWGkpJty/VPJH50sHosi4jsqqIuq9oyjzJEcaJlpGvxHZylrtV8mWIIaR
mnfs6z5ayBqAjayM/KIAiEhqCRfqyp9KNAeCUGE6qk/AZxF0mVeCEzwJJR+g
mrD1pb/v33JrYhUlm5wbOUDPZbIx8nBBS+nbLUn517MCFbgUWR6OWCTJczXH
176tZMpEUVu5kDFKE2JSlwg3p7/+D+buGrho1PIx6pz+jf14gGibQK/VGaiQ
rlJnV+pFHX2NdwsKPKFR/GJ9J6owJNBEEcN5YbB3geAS6hM1gTNE8tGp25nW
L/Qgd6RUNeMOyNEaV+2pLkjgTDOOp7Hxnv63LNrKA3/wxKvcbOBS/GqVpIXM
+5TXITmPy+H7Tpeh6Opp0Hfp+0GRm/2Meh4ikgc/mauUMWjo9hLiRC8Pr2fM
fKQ14ZHBv+602jL9RmotP6UaSbNXJU+8UwRqLNYa3xYKPAn9eMUht454tRqm
ee36tF1KELeKgO6COEExlrfT3KCfOVeypJGpWsVXlyf3T02KEgqU7Mmfo33M
mXZiSAvK21FDax92y2Rd5kxkWJV+5rteB4e/bsc5Dl/n/BtRJ9kki2Cb4lcW
lGx0rci4aQy8uoYflVNtZ2OzJYMLUtLlqdyzVwm/+lo8W4bp9WI7f2/g+NW7
eMnP5DQKZ94wXkuQBsnpvDv7ALU+7WYkQ827GUxavRmHLO4OSppSyL0PwmMC
xfF0NvmCBwJkPByY23DMTSQj56sjFCJAdXqDp8UHUOAF5pvESeXEZZyA1V8X
m3tpslxKtvoyzhvGTwLAC79EfsgxbLM3n8umxILXLi5392j+4xIJ9HN757Tc
REFOBtZt2Zdnvl+l3OU04rQ62gXXeOhcvT9zE93BGSFAcR907IStzNOEK7b4
SNrnHa5aszSFIwnS349/q5MRkgWo0baap0gQVv2Oe+gdjew/aUyLlokVIW94
MFRPwK0/plFqkXTsGv2a5/E6rjQPPVh7K/E+Og+abG3jTBd3oXoopfULpRKu
fMyA/4dahWDmrnJuZhLQAa53OnRkgzo5fWxqyE49Epcs7Mowyx7rOJ5mGRL5
Wjv75ti5nCvx7HZTeism8Ilh1mVN5Slpgu7He8P1MANgmKTXkorTV66j96w1
r3TQi7FU9mfwq+XNXQiWOR1f1t89V9J+xvs1gz1ups2c9xwjAStb/0GMQ7Il
vNeuUGuR5RUjomIM798CMKugX0yZthoeVNBBqr255wVS6Z7ggSko6VnEVRn1
Vw6qhYC11R1iEvxyf7EOCGMUMU9m7VjlWtz8kZUpKHpqEikqkPTwWQzbj++V
nahOI+0QOb9qePK3THEYa1Q5IOVls3uLSPO6eLPwQ3ALHtvJrBizK6LHQZ98
iC/JGz8Xcr5EAZTfNwnDmr00QpTX+3Ua7SpD+y1peUpasGwUYojIMli8Trz3
orFnGa1pgjowpA4jZZnrPU8TKm0pXoyEmip0WDmhy9A5eMO9nV9j72MosEQ+
TJwTwbl1RLwJ8bWVY1E74kZUukw6ezKYdsvjMx/n4doHoh279HKQ6vkO3wrQ
s6C1NX0OoJezQRur4U4WAhWmLK3ky0M2tIqvLevezwsAU+PMPEJSnpMfbFk/
ID5aCFbBA3PDZaaJfo7LF9yljIdyOcNOzaEB/0DqUfsHSdO+iPvgXfmLx93B
Vf+a3MMk6IcLG3i1g3HA2kbbv+6RxF9iRTPOfXibQHUJYj4+HWSaO61vt4Es
dKwYxYu9WVCys6iKy759VnxxDo9cQhlUaKG4ZIoxItQIS06jNZG4jnQXHbKJ
tXN9phFZG/Pe/Q4KgjOnOeG9OKIsxc42qaSfi0SSH2q++osvMgGkGp2Y3k4G
zBRRvbXqlz3eaHXSTq21f/L0Dgr/xJy5R7sbiP1WZhvxfgdK5+sBTc5NiHBz
rO3iNZ5XScEF6Ul0ezpJo34TPRX7zRumQYc4XFb85ValzKUwOGj49eO2LeIX
+L1sT9CY3IxoOQdKvBK7T6XY+1DIxCiPZl5+Eho6zFygt/BxjUSt6tkt/6s9
2y+a+oXkPUJaaqA1lCJf5LlNDib8XkteKLREdOaOZEEddHo4DW0aGhcgktm6
3Ea/QfnY+BHKHoJ0JecQVMNqD16RTSTtf5qMqK4Rxl13+etuSKoSyAInSuEh
iq+BD7ZfgYHgU1Y6puXyTtR4XtSarRwTjfh0/MVAIILQZ4NC9KO5oyqkfYgY
i9TdGz6iL6t1T+4QoO7nMl6MxTUBgHaV0u0lPYUvdyV9sLNarFUWFo4Xlj1K
eyJaclYQqEhpHyyR6Q/34GJI6t9/0g7dUVenOD5bQSgU7TvzBvnwelfxuBuQ
63H+HwQE8EWEDlIeClxPO0IjK+PpNgy0eVdCGTTjxvVn9fYVGRtHXgRvwvTU
M/slRc3aOssRaazXiP1iYxmXDzzLdmlW+qPQJ0Jtxt3CLpneI4eOV8Myckwp
8uuCab13zyFTFEeVoPAhsZq+JfwMVr1HOFr5H4lkRpIk1UTHzQGRAUWuONHn
6C0ij2IGdZ6N8y5mrLKIjX6jSw5sjoReWsGx7OmY6IZAbg+LYTphluevvSmW
K+E89OPiZd+xlgqvat4LnEL2aKD9W6MRmWFW/Fz5Qm8r7igIaFSAG14CQqb7
Bur6INQmPUSK4HoJfsF+plUV8jKyDSHDw0EQydptrAfl0xQih41BUnIMY+eU
l2DATjaS05S42yPcxm2yVrUzm9IbC+BBECSSSSNR9ZVBzKnIETdAHvC1Cc6Y
FAcJLemEVeeF5NERdcxXpgKrgE2bGFJ7ALlmbenzizBub13SCwhSdeNdZZ52
hswH/V+EeIaddHQ9XbA3le3SaIqFlCHFmH6fgUyi1dKOPRsR99u67cSo42Zf
WJRdhPJdCF6zsWXgiI+nslPOQ4LkNjjrY+vJfaBkhCQGFPnzbrXASbqzVIB6
0undDbjVG3wtnP+d+BgJjB2ayTxAIJms/innQr1CypNMdFoPBY4+dHIP2EFj
k0ZsQETJF3Tt/sciAcW9Wg+AGiv6s8sxvYp+nSYPZGROgaGGwrF35+iwGIPp
UG64EQ08OrZxWhzdsAKZFwBCpuPLx74RUdG39h6QBK456Ez5I4Q7WubxhJV/
Js5ltTDZOJPp/fWdcBfjJfp6KwQ9N7v7sj5/mD/k0pS3Imqj70Oxh5D8okcn
xwkerrqD7DYBlKHfHdm107L38I34Bm0a7lz+rMIWuh2hRvASEwTfZCwpFX0Y
YpiVdDqwfKWAm+kEA2e8vPoG9trejU5yX5U8dyzDZ7lfNZ4Ijp0I45B4m4rL
+DXc2L+ClUmK+24XsLiyw4P5OLNv+/5nijj7/w4504V67ZAGZzoiWMU3lXrs
GCH7C+JcQaUkebxaQYEJsEGIlvwLSeFvh1WEgl6SYtG24aq1Pa80q/FIA9c6
aVWLiEVUFAjUAUONnvchP98ix7I/hMpzaaJUTixA1+LCnxfa09pzDbRXaueC
VBY1A76FpLfa+xGWa8pt9Y4Uig9WxSB9tn8OV2RBe5VqODftiy49l9+xezGe
5enuK5ky9nI8wnjo5QmI88H8IF/xEggry97hIbmu0QfQ2lt51fg2oxNFVyK7
WD3NfsjFdzezHiyIgLdGMGHaASyv3L7jwXUSDZGaADfFTrBj8+tw7e2BO1bs
2rB+5JqrjJ1TV/wcyEB6ZE1rvEHaxodQc6iGk2y3DWS7cWE4gEz8vRQkE03o
Go6R1URH0xwg09GrI83zxkpCO2EWDGjJ+6IebPfJrepQM9pokD2/Od0SFz2k
Pc8bynlikbH05RfBxpxqXp9jAExq/71ZGrRe6zMEp9W4Fi77IvhEKIIUzexO
SZQFleobGaGvdX1tSY6kwZkBdZz8a8TziWbM3uNCvZycpAe/FVaTeRZ6QQUR
kbs8wafgcqPrXKXt8s158A0Jdpalhe/Mb0ntW2fhUG7+vUH3JjRoCSQ52pUR
LJjHnYe2ELM8kevBa9u9Lf4NhL74yyzN6bEwdetctkm887GoBPMTr+maVLki
5+VRbNm7slX1A6xFQGXrYpS7aItjpHCqORJng4140JqrNVgQp2fx6QVVWlO3
t+CEkhpf8lUf94Zqv/Hzfq4DyEf08sFMr5dDp+IQ0IijmqZFnOtqKHuY64ls
sXpLqUCcG00vP4dDjE3MlFu9/Es++fDy/yl6R18kPV/RnCzNSI6xC1zIWGeu
8phO/LXCfJQ4ximnrUTxXkfkrCKhyqbAWaahRLLsSxdg23RZzGg603UJSY7F
G+n684dhmrcSmUgemOzmcJwA9lUQytQZY9oSf77ZGDPu+mtsowzDnQn4+VZH
o+TAt09FgIQ7bhxLQ5uxXgqc8pC1d5jZaxzas/gJXdodGyaCcejlgXVPKqD2
MrwHBX6+r+FRV5wtAqmvzH5fgIL/bA3WJvCOEMJluSy4L6P6Q82QDfG4gDQF
UhGGmAdvwwHlC4OxaZJsgv+E+cHrb+CvhOAROywTctpgSFB2RRADWSChDxmL
6f3XIrjS1wq4sH/gbEcCcKmm56mRD6HDFqMCEMXHguT/sms4zRKCliHfBbJO
ctXpBdU+YxXSwc4f5katU/jYJHOyhjHH0K++3ijFcc53ICAHEFdX2aqdalwE
+rO6hYzGKVv7Db3w74XcwbUpjuxh6z0MTHngSTg2IDxs50VBPW7nSqucTgaC
b2sRyxXjnK1RizJJw0izKGkd2D2NFLe2Ps4jaoTc7WFSh3NKWvYHVE8UW4xd
faxrvyIlo3VZFTMfpGIy5Cbh+4iiuczvrpbGSP1Jf4j+gckT4eTMZbzmsM5Z
ymd0S5R0Fw4ZbnazPzPzTQsVLPgQHH5vpPfVuEiJUn6qazdiEY+aYsHyfTOV
2sxW32/1k2UHuhJpquDqUa8V5+1inxtx4c/DlxQKaoWADGHy+dppsGJdh/vg
3dvO6aWcKq46qmPZhOpL7rIaKeFIm1HkVJ+cVCumdT//nummuXAI9NZuKJgU
+PSEpfuk/PXHzFbFM1dTKMgHymZ1o2LLyhWRvtYA+FRM/mCme1KPW5WQ3T2N
gF/CKeLrRePVUj2IdZbqTK8MsI8d9ZqI4DtClXejhOP07bpdgRl2zeN7HhkE
hHdyIPd8nVIYnBRNxqc2+QEX3W0t1Pu4Xgs4egeOufKSm1fxo4bKRgqAyrOp
RcKFkGWdjzu6VCCrl+kuz5jZvNKfthmnSvaDbmkz9vSKTeQ2d5pGAMmDrPCD
ZVbNwAfUhXH6xkKFmoOnZVX7DB9MKgqLjQdJ/xbg7+g7Y6g0ibqBS14vt0Vf
+gIiDCGZ+gJaXJUSlhGAk6WsuuMMk29j/0g9mY7Wag4EqY4A4hoeY1tI1wPi
lq7M9PI6igo9O7SUHl5iLFL+4uKSdsFA+HHR9Qbp877lMVwac7tF0YmoJRXi
oO8/7v8GcmDsv7t8SDyofYGnKXbBHoUKVdjfpx1Y4hz9ZfgdcX5Ae7wPUM8+
rHXJfVWQpIHHb8Q6zgVjAJwznOLPtiodqnxSZHz6oNRkPnB1AZmYE7HLg7JU
cCOn5rUxNvCZr1OLS6/Oq5Q9M5NY6IjlrsrOVJYbb7HwstAlQF5ytCP+cnff
N1MY47+o7DVqeZCBHBbcu0R6uNmqq8TAZeDMK87DSY/Jw+3858eGhqJaoSme
fv2Z+tBDcfar9t4I/LYMt7HYcVESdmg02hcAZv/A7FQ2Uqu/GzYihmRqXkiH
4N6NI/kRYvwCaDCrnbljAckB+umJmatWTe5drosoe/IJUS96WI3fYJA4SsPp
wMiYopRMGGKwPsHT3lKA0XZHI59P5WGixI3gvTx8z+3MHaKqpZJfHbSUSVZr
178tGZyMAyYOqBQTA7RG9e/FHqGjmX1WGZdCqff1DKyxuNUtsE9hWxiewDKy
5fN3QajLBFzu3VSnPk8VfUM7Ekt1Kq8VJsLQSicJxa3rEj8h/KNvGpVel1Aa
P9p/cp44FCJhQPFaVO/CdHXdcjkRW0hPvprrc4Abp9Uh68c5WWDrgczZJc5B
Q6icRAqyK6oOZyv+f8QuMptl8eGR6EknhYLEFUs1LupS+LkAMUZodZQzxpuJ
ErO6SvLnsyERes1/upLZxg5SFdktCNp5r3RgNMe68kgq0g7mpuS4S59kn1kc
2SkoXALswZnI0ieYjypod9/i3SIoxjyZy4zdEzCX+JQD7Z2kg2cfhHPB32a3
owAb7ydSn/MZvNRmw6LX2SI8XQli0sKjX4nHkJ/RAVvOtB49gMxtU23vNpeY
0hdpcIVD5h/vVBiiLpEzKmLApwzXm50SQayoY59AJe7v7Qgc6+dtxEXy6dhX
WkGbL3EKV1IFOnYFdoIBR2mquG/soN+unr7RJApBGl1+npfc/lOKj45gHJaM
PghkYsGu3WbDKcezrXft1HI3Z1yifcmBBjYaXnYBdInXfDT69owQ//n6wFfJ
p0DOqh1gSNOEBy1Zg2LjDH+sA21PgbRg4OVw3YdDwTzGvNELWzhE3lwS68fe
yr08csjPU9/F+ykJ5LYkNfA+1Eqcu7FZBkYsED3chHLWPEUgYHt09EGFEX85
ki+EyUqh/6DobQaXYXkphdOQvc4VW6LgVsu33X/nChqxrpkjp2cP6ayVBtq5
lrhx0sTpObba7B66l+JuDue2jN65B4x83dUZG5CZ9Gr0KUmH5cHonDN4MiRp
vntgIJ1zTIYc+QdEikkvKLGacluBQBDaO3cFjQf+QfdM89DaXKq8zo8n+8WJ
K2CjuQq/GKZBpYT0Rlc70EW1mCSrJcNsYO5zp9Xp0rH660u9O2LdIT9j1yZW
dSzCCxtnQM9kNkB7fzg0AqR7FoOUxfrx15Q+Xdd79IEs19ncimCpOd1KyW/0
o8CSPwak+8P6DBUkDEH4a2JUlWIeG0UZpvzTydoY8ITL24vdYYcpiOFHvnqQ
OVe6tWPkkmf9RwfDCaPK3Yozzm2Hnw7nDzp3p9geXInY0BpeWfT3cyKtEFl1
NHJOyZkoHDyYMncfCuVNbePRb1e8AKqB0b09r3bUJBEy3AJ9CyXBpAGr3llZ
TZ/YGnL+T+SEOdgiDeECejv7WjR6b3c/3m1k6hF/rjr7yi1cj47JVqqO5AfJ
3dTXitjs2XagtmueYppKf/RZgB+iUVrp1EtRaXQghNX9EiGXuDbByGe0/Q6I
WDVyMfBxe1pofba3FQjl4enfKEp7MRLoqCtORVsr2G6l3fxdm+vuL0Rweopn
k5KN1B6ItnG4I/Ie+6KtVxDO4elDR5dGbAkSapvlRmKzGIyUKaGE+cheAXvU
rhLjDJPGIrr6+ZdVSE25HG58LdVFwhp09FTitTngdllfSHeQqb+E1Zsjleii
0n7tw1z71Q1dyg2mTs9xArbEwyePvtgBrrsgFyHe1EDUTfgTkqs0pmAlgQtc
mt5kI12BupYlUWkyc6lEa9eUvGtavTphHvgelFh1z8G5nwPwxaHYq1wil7dy
sGr0V1Gu7196CFyEcsC5ycYLqjnx53UwtqH/nfxNanm6/qvarxmuSobyz3au
AqSM5ZJAHYd6lWIBVuqmUaZDv7XmTz63gUI81wL4NjSmjN9Xyj6q/jhEQ70B
fwYR+5CayfsW9geLUcO++svA5OtsjVYpFIHTUUTf+KRaoQ5IT5fjd3YfJJKD
1mZB4KrcN5U2dQ+ZWDddwWnY4ZkNy8xmHXBRm0/RMihqNC5R4BKsIOnCACn2
7AEhb7MzMyKFM0OUI26FPTGu307OCTIJn8EDhrwHt9Io7NpuVXDZm+O0WWmT
EeYS28c5D8l07SksHcAYaPNtkAfS80ETPeGMpCBECjNSrHzkxR4g5zV/MNLL
l9xegX8gFGJ1/9oVEn07atqfbYPloE5geB6hYXrq6wfQc9ccIQP16ZW5JOMu
KjY0uuuEJnLqpN/BIg8R6IaLBnctYHQBKoG6uaxSU3bnIqART4J/HrDlryG7
sjHAg6xH0fZaWJcvz2i+OtkI6gw5YbcaCu+f18U8NJJPGAPLVQ5tQkTyWODc
Ei5NW4JUevKEJJGe2EF3HOXKP2rVTJxfMJ7sh1bD83e2agCi/uoY9cBsfYNY
9Rukl9WON37/o5zG++QmxDUZqNGDdugH/ND3riU6iWQl55iuX9CJ1Rn8WWzp
YpPPRCLQ+saBR/nQHBgtK1s2eIHx56IYsdvdaWy37s/uvKkYpQ2yyG+j9W3P
4bB+0oFKwr/DPPf1HPl8V0TG1T060IfHNbITDIP9MduiXghHe9m1EROX9PZV
ivXKcvlKOFGL8nrBskKdlkleux+0Z7CkRZeH83K86wmZ38BxcmriJ9U4cHAc
2c0BhtLi8+LktIYEVZ5QAyVoRJ8NatHbjdgk8fKv3sGcKisxbBx8J6RmB25y
LETTmdPF1myB126xUTjDaOrbj+wY6sshDnuRA0L+qNv/tcCqSOXh72zZgclb
6kbIaFV6dGTtc1qLQzGZrLtITxEY6f4hhz4J5InDbrlWC5FcJr1azsSNawt1
I3BRrDDIttqYSD8NXIg4iNCKfFkjn9GfZAIoBsyhZ9QcviCvnjrGQ6lX59BU
elSuF47QAnhjGyNQvYMJuW2A/fDnkh1+lnUSGIeNGuTtX5mVeo4z1Uv2qW1l
yTQzmLCFxayYXQm+xD/r6BvgRu1HWhaoVQZWBaeGSI3qpqV+fHxQmYPz0PQf
gGGWdeJoP2IW9LHJqsc4ym3Ounb2iuxrWxgJwSC2XdH0mqJyIqXxGgVbjvUc
nqmOaIiTB2LlE3fk1+vMBD+71+67x/qhnjk4pnGvvFWiezjyT8uFPoyJnZtR
OM+uWAhgNPclL7b4yAVFb4U2MLJszZtIh07mSfaMlOuNbmI2rcKmsg11VThn
yNjaBJgkmUfiNfN7sqR1x+L68tWZQdU33pN9pA0NceoCvKZGTnU28cjs7Ij0
1BrKNYGJu6nfmZ25q7BkLvP2rVocdL23J3twuY8SVQnmzx5c8kV42zRN0jMV
eAxXAntUCycthQ3ls4H3CvJkUCH/hsQfxZCgTlW+0sCdepwKyRmnzHZNPHXc
TAVQWKtewndwXMTDpXpg7W9CpCMSKA/c3AaVtKCLSmAKZmed4mnwGaP7vxK1
FYro67DB9xq3ERFLWPjepY0HVy8IYcr9n+y0paLvqpY32U9nfPlngBx82V6i
VKkNfjQFYZFoIhEMeKv5Ysaqr96bY1k9nL/jtBXRV2anQfgwc8ll8RmOCxVE
WaCb1Rj1e/HjCu1RdLgDpPZx+K77bTOXSOksuXzSO7RLNqJxyY1UBZz90YBj
SgJBS19VT/SBtz86ZNnMEits1uPtyeB9pyjT7JFHoWzPjad9RZcyqUkBm8kA
dd6PqgFOLNgdEeBdYx2kOhgsSC8fQ+5qNECAiOffB3POqLthfqg0bHxOzPXj
aY/xV29MUV+ov/Z4XodUD5o/pXBiPkqwFyktZ5HFaW7znhlKIgCRz4TsaYBt
Dael+1YpcupXz683wBTcN1wxcW+5ZN+7Lvh+rxmIg7S9O9NKtD6diPBOlg+z
vUqMyVxf80OPCmq/Tsai3AfS3aXlToEzZL/3naZrrvC3uj2YisH6ZgIUXVD+
sXMKtc/ULqCMotWHDcYMkvABrFRgXbRvKFw7BUOY5Fq/qdqS9P3zP94lhfcV
5NUtj68yVvT0vPjWNktkJsMSv6GW7AZeYVctSytEEP23qfG5yq2E/TVjJL7h
gSe8bp8AOGzyCEVEdNdC/SgHBRmWhPUSNC4bD722gExxwYn9dLfLXuzvK0n0
ruOWM2RoTqWFfBEqCYdLiKWhTLgi4HO1BfEuaufwK1hWtmdiIeoEik6ktyod
7dTgDq0AFhI2+e7LBcs+NDc0cZQhDmUpJp/ukOVlK1B10QgIBe95MPNjxh5s
mFpaVzDYQv6ZB/t1Xryb6d5eUbt05e86wdTxh/yu5SPfA7pq4ur69ZlnRpAZ
QFy8Yn/QGKaKB4tCFL1jwp2Qo5Cxe6TOmYlSJi+s45//j4IN+VkH0H7BCV1N
eifKI9JXQW7PYwMyUVYkHryNRlE4rfha9JzapP63794A2j6ry/EIBor6P5T/
rUiqPjCVbfZq16BwBxnsKPXHD7s9PocoTLI8AzmzbKXb9tmY+AqD/5U3nJN8
PJsBg9ZCxUYN/gxUlQFQCFjoTAQVRQ+X4qu+u11ZkdQ7mC+N+UUeBkwIJ639
skNUlEz8bF3V3UH9hhy9MGAOCPH6AS+N1x++e9dBOu6ixndlCdzBrAziMj+T
v7gLihGRw0THMb0NRgsAz+S+4sKZyVL51Rr9b0nD6TxTrxhlHs+X+kTjhhnr
RJyLr7Q0xeW22yWDPBN1Wx/Z2xIxdApYkQ67W/1XyAb1wV/f+Px4vYi9l6TL
9L5ubTsa0IJUaeC6C87YxEe7AybExuH39uhptWay180+4Vx9dWulv0SfbIKw
b5rv3WtIr0rg/Joxz4ITm7lYZmEetZoeKv+mgD7SGiKfDBU2etC8FcI/rtlv
Nw9b2VS8X/vqALG9NGTTI9eob5h9kuIsJ8+FhXXdECiNv1TISLvnbQBP2sPH
uonBE7cKp5ZkOE6ckyZ7Tz3ONPgHfa+CYwFVqyYb3fzyLfzEqjoVbTa2vgoK
tUilY0bb6a27CoDqJKqeJYwqh/fKSzgKiNAU32wISQGoZyP05TLChOBxTpyq
YPHqyuE1veBr9EAywbtskNA+LgEs/h9alSpbCa3qR5ODvAk5bRVC+fYXedwQ
D1S9hemcYaHY1GUkNF29y/GVNC2xEBZEyVuCMOHXPhrSjTjMuvaXGren3+p8
fBLRMy9otORoYneMrZXLRj/CByg/7ONqC5b4+gS8ljsQ95zNaj1r3arj5V/0
b0huEoeFbM3ymui9Rk++uPZvq03/HvlMXzzqMBPRp72yXQ8Y7WL9l7vK1pl5
vZF4ux7FQLkBx2pDQ4yPxOVxLPgPPss8VGC+EGR+w+amUqFBt91FVEanGgHN
Oa2q+7p2s0FbTPS3+/ruEEN4tsMbrB4xSI/p7cRpSGvLxSKijIKkcWnnhxEb
V5hQWgZ345qf5V9xWRUJG1KBZCE+sSzWzfvWfaUMaGMd+vWhykKLip6CGBSE
f3Mn1VU70cxLy9biEag6OyDFAd0XNd/wGsstDKl6Aqr/1lnkv+cJZbuB2g95
2RFtDyEKij2qgxxPp4ZUMw9+DcZxl+76b3FpW0LEG5HBEq0WvFhudpUNgo6q
SmQCmRYdP65Jr345XiEKjAO/45OglApcq7XAzZ/K1MOOmyuNH7P7Ivo408yG
kEQxss/akjEOOpIX4DtuewX+6Zg2QKSSvlWfUr57TcDo5gqzKo2HKMsGMEKx
gz2ThyD1EmJOG30G/fYpJHHUJbuKiQJ6kGhae6+lZ05eG9XFtRNso52C1gCj
aUuNxrJnIEfuj+VD4bWuyLnTs5hutuPx/7fpREYeRE+9CcEk3wo6u73jJ+4O
DQEdpkWwUPLSsWUOSGFP3TLBbRAzc3KbA6joUV2+PAbt0eznuISE5YpgXaCr
oapdmI/Fu1niOYRLH4Lt6WvlmQpzjZML54SstJ/hHLan7NFL14oRChlM0qq3
QyKCuKA+AyMO3YSj+r0s/RPSmqiHiHRC8KqUnD2yOWok1npz5xbijeTlAULp
fPe1Djl8svCPCSrYwB5DJN+O9f+lQv7hjFeQgN9ZlVu+Fke4ekv0VJBHV9a7
RuzHcfBjFLH3nKcij3glo5wjUXu1Y5+c42bWh/916SeZvdjKs9aBgX4msiTY
l8o4uRRTfBPYQGFVH5rhfFU4EgbRwmhgk0fb22kYeHcuhmne2V7VSw+hyjRJ
fKVR/Huh9XNk9l5U6+y4i4UmDIGVoTsNslcxGXudg7jnzD7uDactwBmQeg0e
wT3+5HTkdmOU+q0w4R5OdpnseuDpl30uTJPqIljEkY7Az7YTgYhJWDTMDSmY
x0gORzXsbakEv0vaqqflhaoXFt4891EuSMrUEH1mECuxtj5u7IlnApclIscI
F8Zfl6pXrBElLcnyxt7O2rcjX4qa1PV6sSP6EqXGiuaoaIFOni4w/btknyKA
LqkLKWy4MUZ9gbie8T75AEXFdsGrPdb440j+CJjMZyild2q4rdx0ZzgiOlap
sQXbRI7MTOPhuc2Sx2esQdhSaSXkx1SRUkbLEBB7J7QfQXNkr7vuajMHEc/s
Es/F6ji3R8JM0VqyJDCvKJTGTT5TDVN6XTXWRDW+RrgMT+YNeg7KEMHusITx
t611gQiaYpBgjQ0c2hJCy9xLhMxMnOy8jj6ku0KHmfDd/qQo9ZmVBNoM1gR3
1L4k6WeHsntAYNSEUYOWcJTzEWRAN1/+l+Z4L9cL2xgbg/P2BSBMLT/TP4Je
m6H4l3hARM5NlMo6dQIHEQ1H3DVyi5iNA5sVXgv3oC+lZZA33MgZxd+p7hXE
y+wRh3fYryOk5NzttTnvrniB4nNazXMOhE+EWQqThBJlKuKwxQAqMQBffeW4
4eZqYHwDCRjAHZ61nN2yMA+TEzyUWoo775L7OjgKHQ8NyfSOowMgtWuhLEcn
GuM0cU3XG5bKR6QOm6la9nHOQ0Js+sElIyq/LH0Qvts/ODVGWKomPKeLa6LH
RxNmiNAA5iyKlw//hk6uTRjTfv0GkFl2URtqhyNO/6dNspfhpL93FXh4YuQW
Yb3CLGdAkznvfZmSA5IGlAuET2Qg2eqhjOyAl0aTSATFA3QPQzv3+MA6/OMU
G94VA8Lxu4kKgIkeh4Nt8vPCAwiGMvYrzEHPs5Qiv6U+2F+ZVsmrKoF7cflt
JSPYVnHClA7Amg7uQsxACm0ZbIborrm2jBkPPPfiR6cqf3YTl2IFO0DCa5eV
h/r4ofFikXA8oMm36oinJ7HTO4gBWMIxy2DXjnKrrIwFO6GnkuY4O0dxQb/q
WFO9G6sh/EjNuwy+OSvTGm+r+j4y/ugi8DPptBx5DrHC7AA1eOhC3eN6qxQR
8m7cM7R9OlAqzTSmSZ/EB4BE4bq14Ze+2IoRWzH0/aSu79NjWMI9FvihrAu3
3V7Q/NaZg6Zyf5YH9tGxeqU1LV+7Ig1j3GSMH66c8wdZ2ujvYnTww3gK+07N
ooXvqEIbk/UUyL1znDA9VrQRhfnc1dacNA4MOIZbftuG1RrJPHDjCrY6uH4r
x796e7ZwZZX7I3dTDMibvyXo0vCSmb8KPyp2UfpMHY8FlTw833LAvXYnmeZQ
xzFvr/RJVsJuqbGBIu1OskUPzdaclA1AaxRy2Wxx80Sw2iHSGMiCZXb4udl1
gC2Y3Bki+quCKZSpkVfIPGdnNjcWdYcbgV79l7A68uHAQTuybwaHWgrnj5uw
K2+7FxywzI+4xUxMvsU8PsEyz2hMnJPADRByuAi+CPkCBn4fNaIrk3cEB8eA
zVSTyb/+D36VYmU2uQ93uyrjSaVUNzbNiO5MaiL8GJYScHjnfAxT6Z3vXzSq
OZCW/tXao7uQ/6usOg6h/XO3VO3ud6O4BYv/kdEXY4lGNpUpz4KBCpc1c0Gh
GzIx5iuxARbLipynwJOVzAq4txxow9gf951DHyx1mTeBxROUXxOXRmLRJMnx
3mbAcrMgIjdyCZ6v4ZaoUE8K09CL8wXFctTylrwpZUAJspwIkkJORjzJqBh1
MK4va9guWwLmNxHhjIjMMkhfpU0wvy/jUmoYuXIUVkpw6VsKULE5MFEXxctO
hE+J/hgqiVdxzBpt/ECqv2ByWt9PnPf7hMvjWy3ilCmEW1JGEX0YROjmKQYo
SvTlUCflQbOtlyj8/dduVV7q/IMOWdJQxkl7UwYOtq3q1SXo9ykVLKqS7PyA
pwM40WGgAD9KaT+0BhrQ6d6xe6INr6cyRzZsAvg8v7qTdtSwqzJG5ZDcQLA0
rbpw3ZNfFtG/Jl617xWskF1xophoZmc6fiOSeCE32erI4x3kXB8Z9ifBc6aF
6SchMT36L3lPzL6nEkl31ftziBq6aMvcQCRVhp5ma59AZLoHc7hv0FedBX33
Y2Iwjh0WhFUX41aLr8PQVghnhb8L5C0el36mDmB3+SUE6Pfg2AYP6h1EFhPZ
HLYGrJqpccsXp8dkVMtD+mhrWU19dTz4rKfUrnZgyI+SknW3FTWJU+UUg+CI
UR+ZJm6AzVUJALeVXXb5nNpkyFp4EzwoPzYnbz4EFsBjoYu/ldNFnq3i7y5K
L+s7A7/i0YZ9SG4vYWzQngjlMYDbLZtsWeZUXpOpkH4HKcATKeolI3kuDPWB
6vq5UndwWbnDp8zkcY+f2SDk1bfjtBSWpC1G4toOb8vyvkJC2FYNBwb81TiU
d3jNbNuukHRim0Elz5z6yke+7H2i7rh/uZ1jrN5JjoCptDNe+y9gZ+eXLb5Y
LXhPj7fI9vBH/YsmHWHQNFZEV4joJvzl2tVJLaCp5czIuzQ6OjgyUS/O+ynr
ll/lhJH/Ef4HdstXHa0eBa8OECbZ9ytKRDBC/aHZ/XNfoRrS57XRi/eK+0v+
+KCLFUcjqArWuVbZWl2Vosw5UFrfbPFWpxWk+93jURkeMZOCmEb8NwkMt/pW
aMiK2OS/qjnH4X56feB8D8cyy1qGqRqXJZxgkC903hK37d25iNIVRG6qus7h
bB66611Ga+C5crm/6b29nmIkeq0YocoOAXJLnFf/SWEtf1M3ouasC9RPZUSU
V6GpzRFWKJvdi40S8Dq+3qPFVlt4xs7IfOuXsQeqKs9D1V/egiZY2062j26i
JYhYFPxa3l8GemSefS0FwDeOCV3+4fcPir33lEe9u7QQqjTbjReR3NpQV+01
D5mTZCEN/Nz+8xP2r2T2K3Ex4S3/NAsSkLB8c124yUOt7jxbHGE4VPFOIN+r
hHjKvurYreV2yZyRjXwqH1aR+O6uWBq1LJDg/Pm64D3D0ANt3d4h1oEld0nW
RxMAxQgkVRkYU61eEVluk858JT3HwbIthiehkKc3GP87xM0SBWWmBkg3JDc+
yfyfYBO5xCM64LWheCNgnhKP3x8zO6O0JBDX2gzfoeh+RaQgS3w7xz7uNFAD
aeKvBOZ+4Rn1TZzATpQRY4ILCBkx0qaWQRXLajXX60gh6bHYpGvGm2i/CNtt
vVjzv9b9zdfElWDTayarYxp0sLMwZFwDg6KOCZgngJbzV2JRsuTGgv4SOphx
ERu8y4kL9m7M4syQnY3Kjrpwm/RC2FAtovIJIj4ilSQ1734WPcrE3h06ZM3N
lNP7iU37fpuRuJPysjFLLyyXZnm6HDxPxEVNo2sLF8Iv4CMwyhI2HcDvOcBF
nRLlofy+hNNNv3v17j9A4jGRkdtWbChCfbxsD9eaA5q6EffbpAZS1I2m6Kx2
tAViHpK0gP6oIHOfprAAA/LNCezgQZpE87uwsN6fXxQ3efw0rNmDy0+Cn9O5
Nc8T1vMm+t/he6l1GuVA2zTi2b1w3sL+eGF6O9i7O8K+QMnZnIRbc+jp3UIH
Egd3P9DPY1jsM8dZyUl2lcdWDIoVpsb+SR2yGjwpf9mD7eJdwqRSNcxKDIYc
wUYdMN0/ZOw4ktdpK8vkB7n96dBkXDV0DAjUwV5Q8Us/l8jkYbaKug9IBYtC
SWs+vkARjTnUBbZJDiCDc17PuozIP8A84SOrV4c5GJycJYuRZdShzIFGim7D
04+hdfA4Hi6W/FvR8I2bQGdqUXlkCscO4kkjZvON9KRzvxoSPNQ749I4vq7R
j9Ii8IQb2kLD0Wj3/DkAFvpafOTTpxmVnuiYsIyuU4SpIl4pttiZFZsf3Ejp
BAORlWfX0tP9tBJ73sLGQalS9OSOG1WHu0rX/pkDa0XExVEbG4EXZ9HhfNiy
aZ0wrK7Ns3lH8iYb+cQgb9DoIo4g76mmov1XQmmKdqssdOuTCS+4BlQa7QVS
SHaDB7CMANMEW8aCm8Io+XbBK0b2jpXiuIpQQlyD/tlFSS3OEWfJdt7QZ7+G
gjLSOEFF1JOvVB16ezzNCVUJaSjXISVRS+ijNmH1yrT2qgX4Lwr8eJiXjvP1
wfZx9qfanO8u/yNCcrsGKdqALIpzwkWQ3aXDhDHIZKuleGqbqJJDK0N6yjMX
l3d4dqSHtqr+lnO6zCcAte43bPjw2sVCZPG291/MXY2C5/tvmgHkOvOoqmiK
gI8dAS/yDS4g1Ju4XPhdy7W+cncxpV5ikZvBsDnOdx8nY0bmS7jnbyyX9got
ckaA7DdsoLZeT8JKFVzkOI/8zmwSdiP1VGjpdqdEJOl3bs8Bg14/AvCMorBS
4cyS1DZJBZtaZChK8apmWCxXfpaVRyit4ZggzlSFo20iD6zfT+MzebIcv/ic
Gef/7i+pLndKwik5rndwrvEsehm84m/j1QkwKKgriIb/JwabudF0CwS1QwnP
8jd9hq3shAuz9HoPhjAWrEqVDiipyKWbsZn4XT0Nho9p6yPLJwzaaZ5iHQo9
21toZu2CX98pBoEGOd7JjlqfZPHpxidYc0Kn7jhIMeRZxZ/xRI2ow4QV34Xl
rsgvumBSIARwPJhKUr1qgA/kNd3SAw+L3rDCzV3LdqmKvTM6hQJrCPqoNTPy
UqebB3YSLqYu4uACkyu+ra/WFbEpKAS0Z7750RjIjXxdpZlaDbax8nW+pbni
nvtqFkP8UhRDRe5kZKZTOG8pWe0CHvZTGGzsfontjZXauvNExa1cu8h5OdJ/
zNg9ykSOu2OtuhqKb/3mYBNnvEvc8o4woxvzBjITQrsQjyY5gW4Iy6oDqYaS
09/OGR/6pU24sJVDqccK5fRRTjM2zAm3GXNHkIy4Sla085lth3qXQ8ZJ7nKg
DiKgT9NHEKY3lhCPX5uIq8ukb540qu6eSHcSA9PZPZsPOeO5kPi+X7IWimse
Udo0DAJP5H/xje8wXzi1GXTZCr9E73TjYEijw18NF/HDxQ7xm1zXMaQ4wIC/
ouil5ChOPn4k9ssZhFi6Pt7/cC9aQ33EtNrPLa+ZmHqz/Ktp/HSq8ekyc+hU
upT6jMUBwwrrAT/VvB1gYD9aF69KSBzsZwxixRK5M9WP/gtxcNJ4Vejcxaer
4DXfMZ3bLXO76ZDf6isBm8J4bxw6F87xeqEr139mMklCqspSohENmn+JcQm1
KursNDSbWBWDqkKdP2U8wWD9ffnsRtDv/cd1y949h29sx1l4PtNCoj7ZjE/A
UKVdOCuhkK/QuoZDpyeMFl5YTaOrFZkMQHABcEKQC2Ke9gR3znQ7YyxbHxUn
c51vMGwL7FJyltVdv/4LOK0PZwqUgJ+qONG7bXLnGubM7GlKRtmI90f0QmAq
KmE9Us3Ok8PLf35PYo4/sta89H/HsdUNVsvMnY2UQBdoURUVzyEhFbvVNWRo
Sh+esWYxPOFVpqsrt0X3sS2rWuDQvLodaMF17Jm5jUEaKzZU/QNqSzdkz24Y
EZCpmdT0DtQz73Esr+0q3/ubcn4jYqXFEWSPcUWKLGABOs1l3fW3vaQPNHvc
pJvL+BAB0JBYMQ7MvpEjGWnPaGf/TGWiCHhN13NxJw6sxeSKka2512/tn28C
zYpos/fjdeWkoMN9Rfubp0aq2QO70kpukHC3Jx3cAiIUumoErzbJjk6htV5E
LmxxnELh5ai4YR0yGa/A/AsdFPxjDDqxAZnvf/ycGr39XAokm0K6EueZxnsJ
QA6JJ2FiSc/i2HmTaTcwQFRAbqWXpfhsFYu3gx04l6r1AdgfnDAwyBz/bqfO
otARWXyWCJ6YyP3uvWzbYastxDQrkCPOGhApZ1YM3k0pfMEmeIW8WUmUNF2e
O2NSb9YnkjhcQqSHBreIW+KG943wtV/V2WfpNsHmL5mPXENpdE+5ohtpflO6
uopkPToranrnaVJe+g4qa5Kvf4xeFeXHJZwUfo2Vgr7Lic6xFjFCFJdg02Bl
lWoBW7jL7hLvks+uHbm/ALa41xmnAlwxUB0S+ZiGcSnO8XpHCQLhJ1au+6pv
XAjBjBOoxha3leFgA8P1Aa9vxjNghnYf3C/NwLAam6DY/1vEfJFgN7Tzo5By
8f/dgmUs0Yfmb4OsjZpykXxTiNLDX8C22Lhf/Bn/FpkIq4RnBmp+6El0Yxr6
FuE0xTEb5+nmTVkRiCYTAcGvYMgglLKtwWNGSLP5cWyTf/H/069ygERmQfyi
OCDr8+nHTp9nYBdEO83GFF+o+poCqiTRGaLs9U/RkxTBwYYoWnqqn25g1MAX
/os4ekCi1a5Dn9YxHuhBIqlRcln3xCRVTGBO1aHs9p5GNldN8sjw0pOefvJ/
TuzqF2RvQsPZmnP1j944oMTSbkQEXfmz58xtBWOh/v9berFT5SK1hY/lznAo
HNn9vitHwzgE02rpmOWNi4jxNxA0kSpMTi2WbncgqsA1Tlin2mBPfGo/2JkG
F9215P2jM2eJsUcjo6wp9inDDaTCs5ONFNQqfa+LCekSOKg+aYmogNHah1+v
Am6HPITeUeZl/eMXCTkCqZTMWxoE9YwD9QO4SPmfyaYcVlvaOxRqIS5Cb9Yd
2jkXMVebp322Pox3VdhXktx5YoyxkAAJwvBCsrmyjAvonC9VrmJFh7kOHqyw
kUe5dCEse99+tgQAU8psjBeT8l+BZlLa+CCAM9LQ9f19IIGK2JxX6knwaT6i
AKrA1lKkurXRCqZIZiFZbPoJwNxEXEk1uz0ynGpBGOcUM6OW6vSBQdC1Pcr4
5cYiJ5PZCyxn9UDre2XWHFwjplqbLlQb04I19ocLO5xU2Ru6MuKwZdXb2uGM
lzX37XmAT2gVszn+X6M7Y26ZHuMlG2T+VO6xvETDoumGLiWt1mbsiOZQjo8K
hANGW6UG+E6j/cVtnKkWGYaD2KczqHbI0bQWEgcuy3dKwNv/5xafcjQTHewi
ie1ci0MqNDF14p8W6qCkArmJvhtemK5RO3gIS37ThHpmQomn+gtpjZkSoN9n
2qbh+/lf296TugTgcNdodezTum88hN0KwAILPoIYXkvwqel8JyKNQA9fF2Ee
s7X0MyCml75m1cR9yYzMJur+C/y36Ef13P9s32M4o6QzYpCicBRUsgKvCm4d
5NzeycASwkI3uPtIiQyz13yyLZJ1Uqin9saMCJWe4d2OFWc4vIaHJfTlNq0x
L/ghWEMaMmbXUABT//viqvCjz+WRz2oF/dYaO6CO1LKz+u7HR9FxhsWjZT7t
DAeih3rdg23/PK/xHtTkA7Ja1KW7oLfk+U58npLpnZwKtF4TstDanhth97iE
uu/0w5V4zngt54Xo20sfnpgJyqwKDw2d3fnzAlIBiUQq35VQn0B0cjc5CQXl
Gatez1DU3zSlgGn6m8TBAz+fLjSMR6UpRwgxtw175eTYB0jeJee9titZ3j3m
WTR0/vG9NO/e2KFlJqH7agPbIMWr5vQLA1OdVFuiD+ZJK7H5vWAz9ZwyNuXw
OeB/S6hJcGJHktOBnUg/k2hc/eqK9lzyD6zR/IbAu1r3Tq91zLqTqyacxnaV
irRtC682tTXLJRmqRi83xZsoCvp622JlhN0pLaOQKf0NfnANVdBwgoLDbqm+
5kwdnk3iNMadV01x+BE0ecoZkowAuqoq3fQhH+7evAYhqsvlUu5NW+kXV4Yc
kGCC6HBNLEFhyvDesy95N2xoZD+0Tf6HhPudK+oOr/29voOTN843+B69g3xi
UZZy56rLy+P3Y/i0s2qcQKJO/mr/4Ng0OvGdlKfWZgLcV/paMQQpgzCx8Yoq
Bv1A78pRx3ix5vwZ0Rji49xaSwT2AhHvV4PK4QnnvXQKdFzGAH7dC4VfM6Az
TWhbBVg5uSpTGE04qg+kr9NNa/1RYNgUuN7O1HjLyazUf4FTnOiMti4Ndk/9
uZZ0JmHjojb1KOeA8ci+jRHAIeY0966JPymBg69CRjd9i3pIsZTSIvlMlI1b
AavN09XO+jIvAocNvfbY1h4zd0fHf9FyipvRMKrYUAxWVBN9pNZc9+dUPXg/
T35nb6lqsLlxKjd5xf+JrmblQCwbcnenNwceAras0oqfrofNsSHgwhyzjMWV
OZUO7yoRwxDntFEfTd3t/G0TH0pXCjebVd4gIwrnnJgNEleMb0QQnTKZMc5r
AsSO+XWkWoYYAwwoXzAlLiSKkcmZ0mV788X2nZBcNOuNPTG9tSQsqKha74+R
RMbt4YSLhwISsIV2sWbPUpyWTFsH4EPBEwE2iblRpwpCd79FaYH5CDvAli/C
kKjzqMOcu8x4NvClpMS6d+mceWU6n31YM9ugyQSqIdhonbFB9ljIporI2neJ
vYtuGGUbEiCBe2vNLxbH5xeIb8PvpVls/bv+5V+pW2GY2ZoYdW5X/uoXqAGV
e0MZFlGtEZbaNTHMMD9QseWvGPF1S3imAOc0ZImLC1mQ4wrB17WdkzbzdvKZ
WjMkm0tRA+EvbQxsqQwI+9IjknbYfgZQVZ33hp8DCzFs+jQaDqMsLZy9A3hP
ATc0himhZ7ajSRGg2EFAWY2shqV1AkPFopmGUTgIGruQ/p7YRFmPH+WnF1FJ
LgSn/9J/okl8xCNN5+dZKvAh3/k6NuJxuKloyREUXKPglj+5mOXUq1XXHj++
JROxckpF0o7jV9O5s9H2pw0NwwqTuoHX0nAollL4oj6hmCv3YRgh/DmUEwcm
e0yz5XyrO8k7mc/HU10g29nW/MsvCR5iYSCLujlkbruLOfreBfUhtMPtMilf
tGJVwzjajQqUWjdchap9yzfXZSlt1/Q79/1tI/WPckwo6mRi4ZU3b4xHl890
NkKukvwAtefocMijbhmq0szTf0zkgZNwLZeT7DjKU/a5CgfGSajuJ1wjUWQa
Hj8GzpTeeVU5Tz0JOz+r/aQdA6RN0e3+qWDkNHGPTYLM/MZtae7rYcrlhZMA
HgdRwB3nEND+C3fA8aEjyrnoiccTdF3i7uo16294kmxEKObFpFSdq62FPVdZ
VEkpJroGOmOhMXW//Y/Dy0ZwXUx4NZ0aTTDzbmZvMq2iyQfPnBIe5DgZTuQK
blRpWsgt/3BhwJF7Q8pRBNsENPXGdvr0Kmt558dmktyNZSFI0FE8OdJvQUyf
z73fOv7wZhiixjuYmJNu9tx+WBqHw4Sbx3PkuyeFynGUoFfm36xotOHaDjRQ
QSft3eOO1j6zJTEmcgucxswDjgyEU3xZkOxS1WOb7TE7DAvJDtvnRkCs4fZe
EVH/zeylAXHpKLjPcANsiGcNW9CR/fgvqkCNBsnkWtih8zzHdZIR4FQWQF1/
xRFs0+SlIrouZhJzJH1dxMEIHXEoOx1wCwC4nDYP5lPFqpSTXd9JK7jRW0DM
tMiXba9YXH7KnnYgVf79tjrfLxSY2fFJuTO7IawG0VZU85/U0Y8tgieOVfIt
CthW1A48tj8XODTR2top9BsXjW0m4y/r109CaU8G846V5Zw0fYQZdSRYsiB7
Id3p5jDTj+y49a+EGl5WVQo/DSPvPYTR+AmeZMpw9RD7u4g4sa6VF0DOjqiQ
DzlZ8OvsrQ3VTcXPOvQTMD+dN+UjC4e4809gIO+R5ZmPqNG1kRHl4xX5RR2K
AJ7QEkfrsj1gXcuIPtYE6RXF0KU5DfVe7M5qcdCP17DB5LRheuDBBccplykq
IpqpVLX+L4RtlcMGhfI7s+nuz5fxLrN7orEf9rUC75JKrmr3xQp5T2iaHVDO
T4kQjqpWN9/Qf6LzQe5wi7kWj6CaF9Y10vuwYNYkCbYyCoEv7VKy19Aduu2X
HKgg/+VseOCchXClczoWpgROrVwJjMhc3L70gcl9osdCUYHU9nFKqh3ZSBcb
T04YMlPm7Qnpwqr5QcAW07GHYqiGDga/SPeQKPuYNOSjs5N42nkZbGiIoMWH
aZY+2nK3BPkgswlMgSsFdITKej4+zl9JQ4lMP1Bg/iN999Bt1ryJrZFJRZa0
clIG3ZeeKGWMNs3vdvOy0ZEnlYu/8pUPvLke+8AnQcequakAwqSZgcFTUIwk
JeCLr0fY1TnuT8Ko50j/qkCjL0A5RRPJfC/tp6riZ7mKXzGSuiufAT3hR7JU
XhVTV+wKKTGEJA1JTH1GlBzlAo2e2t1+tQf0KS/MZo/aE7qlqlkamOPWFbyV
rjk3FNmdTbE0gdJF0y/m2l9mwpTsRa55Q88hrf8p02LyHmM92ja0ixpl77KF
eMLrKbPIi72TtbcaKpaURqCBTstQw1t9NEdOAESlLGY1ayZ2uAiwUR3SXBFt
H8N+FPSND2Ph5FmozEbm6+fV7SEaQMBAhsqCM26NxTqvVKBBWtD5d9kbLRR2
ie5O6Evxdayt0BoL8qUWA1NCxwVJ1+FTA4RSlfK/xrfDcuqsEehSl0ZmuBGj
4UamvZkhY/ZMR03qTF6JenA4Nqc8+A2AgHgoe4LYHwFKgRaM+BF7LJL7OYme
amEPqzBMoQXBa5PviPPpA6sPvbUH0EqWosMOlJ6642V5SYYoN3xJJDswBtjt
i0AB7doe3UuQzjpi09v+wnxtEx9ndhHm9QK/jaJXDQLJQp76kyUpCBNkMtLg
talysYBensIk0sN9GB/h6/SSX+Y6iDjX4C8EuSuG/KSTHMjbunWCJT3SfWF5
cV1ekbBwh37PzaWS1I1jqP1+OiEMowBv6PMWtUlvY5UcQG8WUP6h16+BogL7
XrPRe1PU45mB1clHbNE8mc1baPg1ULUhctqQdsEg9riFS9LzmkpP3E1xBNug
O+UqPaet83nPAd5pJuYOkk+WifJTLdyCev994WuYU1o5nlhATMxRwmwJfSdQ
BROKZI+FesYwMF9vADUI2BCzoe6voiYmYeoA4XGobOuiWWob+qhz7ktgd8Wm
MTeI+LWA5chef7hCcPBX7+OAY/VB1264KiGUTVE7lWDXb3ZToJe0LAXisEtR
+ewfFUV7rl0Vr1gMJs+YPaFa52EWIeo2HCNIHmloUBYz+v/7bNRktd9j7JtC
4mF32ornkKuCh265LVKbjY84vs/Sx81jmbQLa0ef4CaBkW5SdAEZBMriiEin
HDddIpAeBroX6hDP5dw17SW74+u+DMaq/ASRckVREyka2g/2xMDeQToBZzWw
DA0oT8pACJvkhR+hWUEsbxYSzEDPeKoWyO7cJdHX0dHAqUXn1l339tfytduF
0ZqZ4FOJXh0BZQgBXd8qCLH7SewL+pQk9PxTSg85LxgcSbUT1v55p6gVNYBL
cjXvpFl2wW3t7zOsMJy2P40vp2AmOfUYvPuqImah9/tNjSkDePtkhLxgJgJC
xp/Q44tuCQfw6xqdVy6JeJKif8qK3i2xUAxsAU7vDisJ4u6+Oa8sReK/BDGC
NSJpD8SSJP2iCQM+dhghNgPTjE2Qf4sdG1RHnNauyIvsvLb3Iezb189HCBd2
lAsYbXxzZetOfTZNqEXn5zuiViLFGXa1fh6gPC1kBkSgs8ztG3bhn03we4xX
4IDVYNJ/uqxlm7A2/KDUQLR8x7sLE5p10aXNhsPd7m/t4YRKJsJTQur2f5Ds
X3U62EGshl6YqZI5PPmpuBesqIFqpJfU43kJcIMaVH3wIop4juv/IUkzDHce
XQiCWs3Qb8PFbcPfFJEBn7Q0O4IJj/kBC3zAvs9d+nSpWl2i3F1yfzW1Z2oG
bz89BPpJf+uTMg3Xltjkd2q4InOwNlKUKJD7848LPKeROKGELyCkTI4Wf+Sn
t4ypI5r7HRMbJS3AXMoEdFcSWvNdXsgQ4Mp/uBDvqOX3HQYrS7OwDDo+GC9u
xWRw4G2n952RMt+aEpX1N5sR/IdgwZflOLP3HshBlar3KLURDO9VlV24/Qi5
67qJLnoI8LQQnuIVdyh952ZQJ1SY2y96LuRVBHv2IEI3SJW9np+nADROWmJB
77ZdXwjD+9Gwtzvz24NBekr6i+tcwdwcuSXeF+5XRSOuuTiNjVv0yeRWaaAG
c+YFU/qQOsn7baevm4FOAaV8fkOU6atSUjgRRO+UvPMatvobrET9SN0KzTSC
Peou/g17aWdLX/vOSR9VkxHdN8gm+ZyALs4WxoR7BeNagG2EojPuWFMfEsWZ
96ogvfZ5sVtaKeXTiOY4d+20sakRk0FxZ+0PyQpM+vNfd/Ohu4BET47lKDJs
8ia4qtuZps4vw2jaa1jK5XFRkNe8mn3AsVyuBPbjP3+Ttaz5UyTM4+ueN3O2
sOOhJvt+asO2XntzW82nQd43KV01tn0QNTWrPqafizhHB2lGmH1j0o5DTUhw
iBQDVG2hOML8yMELis6p6OsgjMRgQh9iyGhSxWfPFOskWJ7IIgaZ+kvUR3dT
QuA2gpFnZFTTLyov7gL5vhUX/pndZKEI7TJ/lGC0gx3LZ5ps3wxeYzpJ/yjU
AAb3UunPitW08xumhAEIT4vOJDJyRnl9d3cUZSV5Osy3Jq5NpZNf0x1y0z0r
wsLGoToe4TCDAhsvjrXR8w72ssKsd3MtguSbNvhhfm0XuIOptxWGo7gPkSBB
eH9ebmxT2sTRxXR53q8WPAqfFcHoaMHmGZWgs4W0oCjEsJ9Xl6LRswnq8Od5
6Wr20AJSm9a8yQpAXY2KkLmMyzuDuMEvsEQdt/k1CJd+W6njyBSbEQUBR0em
dyyiupDCONJhQrl4MkDtQnnUCNxC8aMQlB0CN4j6h5HM6WZaagTtHOWWVlF1
QoB+5cm7/ZYxI4xndiPeuleChmGs5e8G2bgG3OkMF+JIZcwoysuBJC4s9rA7
pzjvSYiwymFf0/IuLDNi84OXLgWraZGueyaka7Ty2nr5jTeGgFj6k25cQb37
gH1bGSTvrCNE0AGijeZNZ41a4jGsu5RjxVJ9uRy/K96gZBoIR/+mxelN9OiW
vDat0jOht0M1mEI/yt+rykwQuECLOxLcVx2yoaAVevUmTHPzPn46VH/gEShP
jyWX2q8D7UwWg4EqSBXEgka+Cnc4XVZ+M+/zdWwi3XVroIlPpcqxHlJwF5Ij
9p24qE4lIIKIWkYQ7nFWEiwJNYq3bH/WrqQXj56ksLbiCDYhRtLSfI6ZzK2k
ADksQ5kunlVDnZJ0X3LfADxszK4ta1qtO9bCOG/fYNE0rYcQmtmSJJoyeWLr
6ztU/barIbDOJHzBlkvz4bfMoqGwfU9t8mQckLwBkXhqmN/QR6xYMoahzrHb
0MP9+xn1tRqD4wlhx+MiCWdtqU0TJJaZ7jCBC3r8KRVPevQxhFA0cymPD//Y
UMlOMBi8vzncfqhVpRIq4WPFxKok7SEybIPDCsfPH8L2zYu4ASRo2xQFMfuV
vdrH07LOcZCilt8UZtq+daoZeHNA4pi6yccTMDVt9TSJuxZv98G0GFCq+xYF
SWXbTDwOXAi0SODOsR7U0zBIERO8b6IMMPaFcRpPGD4bir/JYkRNRdnALka0
o9S9sD+mV2p5bEtt2eXo1pFU7Q2TIBPyTrBlPgVahY/OB4BindZ728y2AdAN
BveboHp5ZCP7iP3F25+WK10ccbpEKEOLaBV4Ho5USBVNFsJnejNEkcdr/vVd
eCd3BFVAyU3DRQOcR+uugmv3YGymuoPIX77Rt1bHgSUrywmKqAuELm0ZgSbG
QfpNOPudcsHOF9fJjD/XHRBbURF5ixU3hM6kiD0XT0PmLMqxy+KpbNHsAvmO
uqM28AVJM9jyDJlyPtpFrZmxJL9BJ1wRdQQAXuUkfhlwd9JYQiiSNpC659ou
hYqnVRNTaOVs0pdUcCS3i0r5JVo9aw8S+Hm0rRjhAhzqCzGEzYIQweQIB/DA
eiyj4+foq/p955H50qp6UxDH2y9+J65lAbkjn5hDt7pqS1Vg5gaEudwH40cT
7tXWBP1Rke+zvJK+G1Ds8nXYaMU6a4VZ4SGLQaobq6p5qSH7++aX+3N1vmIz
b6VXMM1zNyHBtOQURRpfdDCu9GFzhg+UDhH/vPBRnu7ttU86FeBuST2Nujfg
61Knz0VtnWuiPdHuf3Grky59RscVVnNHDg4QTIogRSq8+9zFVAYblu5xJaOv
lFd829PnNSXFapa2SLepNdRo12ux0bqjrSoMLIMbSUDKBANi8h7h49V44RaT
eITTNXL0hMqnZzkHWwZ03pV9n3Fjhqqm05+Z28haK3L5UQJ5pU0DSob9MW1M
QZxEijQPSoI7kD9HdbKmG5/rBQIScdD64S0D4triwkGEp5agw5A1tGSQRcwd
t4EBbWeWxIkoP9TIdUZL0XTHlaEPCRzXe76hP1K65SghiRAW1W3J6KGgm0RF
D8UEc8jHTc9Bz1by3Djm0/RkEsJS6ovcjnepZNSW3qznaMiBM5NlkINqsU/h
/lwVrsb64IdwnQKp9B7EImwMlznpv10YTDrSjaqU9WCmsmxNYR4XIN3VU2TQ
1cn5ziz8n0Ypmx8UdsRLfnF4X8YKNwNDU4qx56KISdetuRmZKzvwSCT3CYBo
uNkE3JuAWp+fUaQUFf6tXY8VHCjFvCyu12A4e7uCxeRwS+szy6/r05tQ4QcA
4apdHgi+pOHc8PxEskuJosT5ha1ZauAlHPXh3nKdwZ+AKUXnohb/TMfpZowl
IU7wPOb3jj7R6SHQg++G+IwQUDMDVJksWN6N+q1M4gXHRqzQihff+pbSLWfM
duHm6bGub33K1lNE3tr2pMOQbO+h0bpvqdHOPJL1AxFjX1TMrM0M/P9tuxuJ
hBf6sD2lqAkjVg1Yxcv/s6trvdx6sM/Mye14SdMmbjZnTjx3qWX94Z8e5vCE
Ki1VTQ4PmOYx3CS8ZdT1bcNON8/3iTtbWv71q9riQnpxMPz5ue2EHsn8P+5c
zcS0rfDFGX1zZivnFLRC4HrfDkEtvsD7bYVxhYRhWxZGvaJg5lDO5emGgpNi
eMZpl1Z9UYR+GA9w6N1tnyBDFiGk8XxhKW9g7cDZxauAfC7TfcXECALwddNl
EzP4DFfzKKEtJFU+yPGlFtY1ty2sqk14U781S7DZvHD1+Eax5ix5Rj8mL+9q
YvKszNWFntN8aUBNnnZ6i7MTdQn/Vqp3b8dNpNehwkxq7eeEaDt5ORnXAXR/
lyyYOZV+2asSyUwWX1y88bmbRiYidSS0HfEKEOJtMDp0nJvHB69lBJWozK7d
h4Y20elSAbBaPF7PdNlDHlfkdCyRmor5LZrvS72CK4AEJ8NzZjNN7X6vTW4i
8FBjA3vsH2J8ZKZkTx6Bhj+FUkM0IW47h3Py023na2F1M/xoopgqE+HbLGqy
F5+cpGcC+gKAl7FXGDiA1v5EBKhpF2oH+FVZIaE8uFk1xWrLuFqZLmCqm1s5
r5CHic+DR55D5Yak4bwtZUPujo2d708sntdSWW5sHVwu3wVZJSuS3+VtNy5f
/1Syijrr7B9I4ReLbVlj8j9AeSlADsKtft2kohUZ6XpgbEz9TVdXKYKKUFmr
7h4Xr4ObxzFFgif0XNxcomonaOb7qk8fGlAmXc79fJw319zHnV59ZhPcc5j6
6KnVRKqgwvFivZ0Iv2jykSIedgbER4/2vdCzFljuBPbJzEm6f0Jc1vDzp/Vu
i7ZjpVeTqhKbaDZowAEO1S8J31PNfxnjOLPktquyW8BTkiadlALbc2f//3YF
7MxVAEJMP4wTgAbDCb0F+uM9FibgxVk7o0NimwDy1a72IdeKLAzcRY+seVfx
wwq9xbcCF6pPCyUJ4Ak3kwmXyZc50XXQxOUH+9kq4izT3QXcRTraIrxhnWqj
9i/NwB+86v4WiumfotcJTNtBtT0DDnmhUHEh/0Z1MdKJ8tfGWxiRZ81963mn
DVvXKzcZM7skddrH7HGtxKlLrEhnXx+SnLrBLLa/VCQx2aP9996hfYwcxyMY
XsVFgyfWPC4wYTD4+8tIaHHxO/h4XR1umNqGKGwt+7HeL6mcSw/JC0C/LNpa
xb0Phcg/53SRRjCDBVxhyf4yEYwFj2utqlVnHd5kDq0QXjbzyQgXLZB299Bn
6NXzyYUO2SlUpX6FYty4BE5zZxNysUQBskgfDOzpmABG6zEQCsi2bYnK9eWF
pHSEkOnOMx9/tokCEdmK541gS3HzJ6kcedbYovuz9D5G9FZZIGCucOs4XOEe
M5fgIb2YQKTaGoglXmXmiwEiNUCmLhBAiVBZD4dYVAX8tzfllvifqlnnk3WY
jQh9M1M0fF2ErbjNLGUbs9Mg5EAfkdfWDhEXUPjh+eQ7wzOUEKSI459P2u9R
OOEUc/fmMJAKJxxZF6/zRWDJ9dxbHMkMy4uJjzcnihTpdw8IiIe8deSgQRQl
eb9Pld4IQIfNhciKLrpOLnhc/ijchujeykjwk3HFl7+1pbeRnKMf7UOGHkYf
NWA7o06dsRHpzjTut8zmb3oYe2gPtIlmCqp0TnHZrFQ50bi09KhbWBAm8dMn
7AkH4OiNIKMSm9IHKAMc/+Uw91BwglN5ssoZaIDsnBRlga4aJswbyt3SA8Y3
lpKXCtiYDbfYbnqVNE7jDMhxF6XfUy8/h7nKyArgY6RTSHPld5NhOHIkwK39
LjafXV9OrC/Hk3oGxvjOR0HZIUks6RbARpva+ujpaJR+smZuKlAva2nAR8qf
+uDDRvhyqRUWoZhMZijfkRO5kRWSOKHYCiAFt/2ypC1jhd+3ZgUqjNWBu2vG
+/1czzq40kr4eDUE3YH4q/byNW87jzQNhkT8ISDYzhxOLOH+tvaKabGwgaGD
mUrEX0WOCDJuyayUim8tso/3O0sQDvkhEFHPlFTIgckwC2+ufcn6/kUHtcYL
sIkasaA5zDj/updwPQAgLWJ6ZR/kFYawbpdPLycaua+xy7A0cxJ2U2IwNQ1q
e02e8zD5era1sIX9JjW56Xy0Xf5QI+fAome9B2ciDh4gI+DKmDe6ecti1n4k
BQ/ilZaJ6K1sf4VzPUjdjNE+RAYQ948uDXu+kjcqJLjnBCwJHtYujRXiL1La
e5ffUQw8s5CXDeMg/baibRbeIuailGBXUf+vQ/BECqS5DXAQC4CB7DPuwvio
WU/IwBu0Wv2iztEkYnAF+fqkvyel3PuRqj2WbTFTpyOlRB8GUVVZijatSuVn
jiqJKEeNpuqHFU0pL0RxbaZFEaldtU6khadugAGNaF2JbBSruduovISRLua4
8n6qAFp51+Hh/7rtFH36rvtpstk55NgstauHhT6kW1mXHXMWAUBgctllyfws
9Rll+IsPiiYSWZ1Cw0Je7NYW+ZsLCA91DkS+EJZLz+7Fosx1LN/e1ot1A69B
wMn3oPs/ZrxCSUG+/hKy4shvOz7nXOAMx8RWOMqjnkNPriNx0XuTbNUI3LBu
UWgnqNQR3UyLpPuiCK9bHIaVU8iAcayO5sGk0CtCjb3t6Wh0mbA6iu0HWz2I
QJG3zX3HiOaCvUiB/SlYMJVNpxWBEkQOsX6J80TRgjpTDen/IFzYT0jXkyL/
6ivyc+ELWW2Q/95RxRhsXm+mYSlSIWyO4yGEPpbVlaxsIpDUTI5sqfEawbIi
4Y8nHHgs6BcA9flwDrTNE9oN/Xi+PoPzMFRJb5emkDmNemKNXcwLHKzVZCXW
00bzkjfAYsMCJf1/bLAAP30NdOw5ePNl5TuNymTNyqKiZjU/Q2F5uRWfQ+4i
kJOupoMbiTrKhqu4gog9qnGD8z/mOhLt5aQ05+rhtbUm/nvIlFOHBsrvpKsk
eZ1jV/HK55xK0avow0JDS6jmh7heQrj+aGVHxJzl8WRrg/4SjJFumaNIqQwI
DZbMv5H0sM8Wd1A4dYPsILHbsvxmP9t7EsJCHKsch7EuRjDWiCAUJTuLqDTg
zmiCrBzgt3zDnO8vfcMwUcxqdzos4JQDdBe5bREZC/1ZKvKd+Xx6bbf4CL7+
c9VensS3Op28z5NsjZdOX+FpIrm6xYsm5LJdIhAKUTMEoKeqjfqOOZWStp0o
k4vRWzkb9eptn+TPiZj7SCQuQKGEo0kqI9IUJcREJ6LPqXXq0/hOle9km+zW
WulUwtEy6bd+etwjTn1sh3h1zKt3cF2oNWdxsokaYnVSKipGEa2scjr++3BK
K3KGQpOHb6ESM8oNwJ6XrcvSW6fm51EXH74QZT9cxmZyZExUdz7xtWzaCitp
AhJjJ2P6+rihGxsh5KgFl7QqiU4upjcKb6b8N/6oYZ5juKGHgkf7Y4aSDbOV
ea7BbvE2WKfDV0g2FbgdgLsPuedoRfZrAy919D6VP5DyskYezMjdlFqTUYk1
m4R7GEAUrkM56JOhZfF3Gx7exBxm17V+sfYkQw9Deq9QPVR4fMZVylTtOjl4
jU7cD4Lul34Y9zbKZAiyb+0CVWITFAMgoBnvuiz4as94Pazr1vF2UlftK0jj
Vd8PxYwudxiLdmIzEneGWDnutIvkoxkc7UrjNkq+ILJNNuV9l49RqXDuFDLX
RySjXqjkYWJ8r2Qvmy51jlVVNYwCVlq+WDFvcop/n+kZ3kQcQrmqD9cAx2is
UrvjCXI9xbv2AQxx6dKzD+JYpvn1DaduoUZ2YT45omervpBDsVKLcqkLV2vn
d8m+XzgAbRxFrpz7HKbEAX6W9+cPUDwEGtHtkMDZ+ai6CBkoYwlD+KPJAPn2
9kmK/wAT1qJ0MXQE0Hl1EezgHWkYQS6XgS+WFNaN7+oqqmvJdRo6Ex+ALIjg
NYK/CjWl4P85U3ro/GANvMqlp4/xwk89TYRq2n+UzVJzMwIry+ENCsNFxDRj
Oj+R9UmPopn8b1Ev3UnX9SZELzdMzj2mpfH9TNedulo0gxux2VipDsKRWw+T
WpDUlQKGvI8e3bk4T3rGupdRBihVXzKFKXNellulgODpGohXsbJ0YmGgKK4b
FV31s83o4UQtZGYUuQfff+VuvCzcHg/SWRC/xtB0qyO7viBBLLc9PCwxQYi2
NDfXPk2pFEP+1y552VjaN2LdypWfJCV12rZKThTdisEDO+MKnCqdDk1Hh2lL
erXoQw82n+AfgapYLISLBpudKveC6XBZQ2XIytwJzs7EP27JzRqsffrwQ0/g
6G9lDG7vfRb6qe4rMnIScqOD1LVg2Y/08UTNqmDjFIAdsi3sqdyKvX4Ugu9V
9E8SCEJhH2JyDCNZbEwAN50ob1NqChBdDj4oEKqcZLngA5OT6IJ8kLOlND/+
kHXq9A4HlUf3OdVtGYwp2aOPu2EyuYiXjFpaPzD+9diwX8MBqc7JsyxhMJFq
c6sLYrFg20cm2hPQ1qVkxggeTFfw5qQ1oNcONe6+aEcu7o4VehXzzy3qG5et
/9Fr9BPka0Dxv2HPe2w1h5MKfiTcrahAOxd+ygM0K94+jj8bFTYHxEzNEi8T
1a3X+UxehxVIt9J6av6VmVQNY5f+hOybgEMgGf2VnjofxhZajx35xQO2K7hY
MgVACTqCIPUmCQ8Vl1HydnzWpn9COa60xQaTCPEzzdp0+TBnmKp77vuPuafh
+B1QG4NSZuiGljFx1iSif2Ol0obwJGLw/Qw6A68QB7Ul5GbwK5hRxtaUgkix
Siccs6NIS6R76t5zmh0fZLctrR5OWa33nHIG5F5VDOfhif13h7POpPLrET7H
+slDpJ3Rcm30OGT+39XG49wKGkjlTy2Dn3ss7JO5r56QeAof8GrXMaOHX/Of
dZSRmLD1ftCOdZ7ixchuuMAeWjo9/a+55/SdMg2fxQnnF4J4llc+vgRSle8M
2ZIE662u59JDq6wiLDZ5JVxzu+3if3BuEnMGF+Nn6bSp4Kv1isg8dlpJ1gjw
s+dHIdKEGZvKBO64c3/ge1bY28BtAdacj5pgS59LuEgpOWzJWwVhZS/FxWTZ
SZA6PIGwUv+5LXaD8fizrCdlaxzqFPrjdiBPdpRKTqqLbqdfESMr0V/Oe+76
wCw0NL7087h8uASAWpW1e6xHVwlAhjIW2TOTVBAfhImC/MGTsGiMu+eEsOC2
03n2ktlJJjneljRLCcm5kFeoGGdIFY2DaH0ESrn2JdEhLKaWcfj2TdMMKuqH
XfC5Jnzw+7WaHBaDXHQIYRKCtyDdXKjy6I3Zjz6AsHXm4mSljXkx2UFxbLhO
/7SaVqMWjNqHsDCV00bOdu1wFs4pmDBAuppvORo/S4Gv8uugNicjBRt7j0CS
HXLVNE5SXZHxgiHvo01RgSMcpbshJnS+6ko4ws4vJgr5SE2ppkiuWnhIYsKF
Y5XGsrAIKmGJWW9Hh7I4IcR0TLQzey5wizKSF/lKTmawKSZSYtlQGx2ie4/I
5TBzEDXqS7Ct+EOCm0Y8USimIdpidBsgux5oFXecdMMhA+PoFIM+i2jIZ2Bl
2DzATrbxAyYKbEp3U+y5ycivrM5Pu6fsPW8xfpB7mAxs2MrOPIiY9WehtZj3
K9cEEBkdNtyaOxF+r451tbffrg/AoDI2zpf9ewOqBP/hxkxJye90Lxl9b1Sx
al1Tty3whW5CKSfq0unvGZ+eQxUaUZnwLD1DJ+Nyg0vFys9yDyDw9XYBFrmz
Nkaj6MqWe2YHSL6fXBH+z0fzF5/Ip2VOdIyQZM/kY+Kb16TbjjaRx/kvyAiA
NE8NrT5VlS5vbZ0cCKLyZMnI9a0QepoHvhKJ/VxV3bjdE3V0wGiCXrSTfXqU
SHEMOBZZy6WuiHKX6U5VoI1VPMiXXWYMB5+dOmaRXMUsirZc5z5f9JEImZo3
WexSHKXJPtHjGPJI/ie0H/d6sirJmstsyeHtSm+MSsh+WJlJIogyhoL1admI
74AUR/yYwT81fCiO83QEcnXuWepHHVrt+3aio4/Q33Ayvu1K65E+lis9xYup
DTv2hEOOnGxdndn0NJGPZCzSVwAcY7AJXjzCGoSbBNTLSns2FNI5IgWo0Nav
8ifoGSug4HS6CovqtAjB6lYVPBwf6QylWTV/xkEtxZv+vejPC0NaQ6qUkcuN
KK7ULrNi+ZuQIv61NprjX8KECRyTSqDJiWj53/QlBGRsV1RPSPJJfSaVcEJj
DbenOfP7L9F9TMoQxID9sQ/3L2kMXMM3/JQKKIwBN1BzZcVoh0xDhRqQLZ4D
S/xlkmuE0fttko9rZVgA40zNcgLdKBxhCcq8jF7ABTDBNu891DFwHFM8S4gi
ekODGizhHtQC+wgiGxrnS+nJEp+R0pu0s1w5m2mkneOsSlcyWyJqI7poXSxW
lzDLpM9jlXEVpfi7Q8QUCmHXXLwl1wXjk9YhU929tukTxdyObUYjO/zib5OB
c0At3bFpSEfoNmr8RAG5EzOd9pUttREjjBXIh8JampKUKsBnQqCE9/QDlAgZ
Jlhb5HVl2Ai2uygHQGSsFJ6JoE+ACzF8xmnMRS/4lGfh/DSkZIznbZJ+hy6O
87DNYwBo3u4EDNaZDh7g/369VVLm6Ej5LK82u34/scKrwl/XIZCXZVVtff7j
nanGg4albrfZFx+sK+QDHu5z4d9qI39bVxqHaMsddJq1NFN+kWdt7iUbxHAL
fuFpZwI3l4pNo3wmXYwCiY1i+vdiurLR/X6kSfgK37Ci9P8mCC6t0QCGcNGt
xvqoTUPWbaGXRd0I7E7QQHcBysltU8aHfG8ZOhZmgUShkLKOWLKnHvMG6BE4
V2/15y4HzlU1LOfk9WFNKYDlOWgVSaX/D6/L2exrNnms6NOotNkStSDoKNKM
bBFuqvPrvoJ05KCQ2+aj1v2uIuBB+6u2TQljapBYuMWda2S6HG+pc5cuGY8b
YRLIbDuTuPlQh+MzmtVZpRwCNl0KXyFvhwG0o+586aewavLHCobHfzmvYgaU
qhs0fluiME0Eh7QzHJycoPtQd9CruopaW8k+W/X7mhfJN7Z8+jquZH7ii5L4
0xiIMGI9vKImKs75jWEYPIb6dmJTuo6muaUkvP+iwg2/ohpuag2pUr6NTCtu
6BdPzmdJR5gJ/NystAuvj0Z17qZU88Gr5ZGT6H1Y6mj4tOufvkGXluW1H0B5
HZRvPIoMSOv72mLXz6B4YMlxD/5ytXzKZfxZHCQWzM/ygcckkc4ivMZYmG1i
3zOFo7xC3h3BbHWj/zWgG1LUMDPJVpcG8otQK2aKmMnVtWOVHOCSA2U/39qi
gRok0e619wOxE3FjKyziE8+naLcNTn67AxihsJkGfXc0gT+3fO97COOcjtnF
bfI81OxZ9Zq7YErcf937rY+ta/XYyWFTZ5BgfWVDj0UWBYZHcfIb8ELeqHrG
5EyntZmb0ZB7QwhDlQ/lZfSgXmXccNJTetIj+AAUxKJSTMSryxMICeLVG79Q
2QIOAmtcF9f2shveJUBo6wBYO5lOJI2Af0EvEKoXp/W9DTBa+hugTwJ+jLKZ
pqIZ8xKYcK42L3216NZboepyf695/AebonB6qdSG52u8a/TkEAb9rTITGN6d
91GeIZgB7FDZg/Ns3ceEn50kgHxh2eYIsvUk20gNf5WjpEOKEYGECcTsEvW8
q7XkpxJT+8u70TKg7IsoKrKAGvKqzXLl2Vp3DaaxUjnJ3hhX3JoN1aP1TUrf
ojKhqyJYkK5dvpvuY6p/PSUJG6aCbw0WoX04fIE7PBNiTmvqUZ/YHMImgICm
b8YYWFUWf3DdvbiG596wgFwynPbPC9pgLaIVGMNQoY3IHyX7ouMe1mfsCeAc
lHQPK/Q2gEkZaaBWd4ne4eJir0gYHiLek9YFGPKz3Q3rEQhAYyTUHJc6qnJ7
VuZyjss8F1jCJSW1eYlERBXb2xug53MP0NldqE1D7d1oCp3q0wnOkpSjhTWE
OpTpwU73EKbTNFc8eYjAxhLIfN9/pZGZip3o1UTNrbshnBopFicnWgZnvE2u
qp5u1v8OGJaHIa+jK+ynG09YPpuY0eva2ylYY5Pc4BGkEqU0zx11Y0ikyNky
yma3AxhaYy9jltjFscudTmrPICNrOvLHDDWbm0PvYglAuasZxDFvJxxco8Fh
iJZBuRwN7uqqeapP7G6PPb/+x/SNZzE4Uiu4YoMOdLsGe3AiAVEUu2rPr9Q4
kCJ1T7fTlwmVZNR782aiOWz1TXmxogzLnIPo1jjD2STl2N3UlCqMDS13g/v+
0ri8r+jIboWmzpw8cUX1TAa9f3lK1HpmjejSI3ViAOZbA4eTToQvJoAJ6B1F
0uMzVIqKtrMRje7j4z2wyprUL+G2kelcWW8H3ep6YCHkfm6jNsAKhD9FYFoE
+oVEW3x9pfi25ccjBE3jUdyyAEvzuTaaZFvyFgjmVPH8oIeFu52PuY8dv1uZ
dEib9Krf9qrOlXSape62Sm6NsdQrwcTPIC2b88kcMBQahBYF7I5AAUuaSg38
sBhEfAhqhwnDn1RFIn/eoVYa7fNrCyyQBmtyS/TpCQR3J5GmWz22H8DrSDiB
lhStMEJiQz5/HunhZfkOtKn+hbUqJIXmffDaKySgTMP49tk6fTtce8Tkkx7h
G0lwC6NSvkTvXGXHVS2mmq6uixd7eA2iJCkwJzVxJj7DJYkX8YjDejtIlQoq
ssWDyOnUZui9Eiz6+aw+nHn8i5X9+lufx4MRaV45VxgBuCvzJKyS2NMvER1G
JlIHqbLhlzmhroAna38SwrjbZIArgORgttHKb4Jv5MurtF9RZSkJaJjU0zJ+
XkJ9+zlcx8VQY8z28oNlYYvcsoCcAIecqpTiRa+40mmZzo6SqVrgWydIeGBb
7CH+gLfiMDnLrDrArBEhLoVuvq6qNzj1eWwVXcSO2OBqh/sUGT6uaPg3rrtD
AV6qsNhXfmwocznjfP7b0wORcWqTtuqxnKpM1GeT/kMfLkhFhCd+DoVPkmm2
gRwA5pKw84RuCfB/NX0eKVkcJ3TB4dOm5Bo5MCPV1P54AdTR0FsgAdjXNlcE
EndsUu+XKE4al06GZTF8V7z96aziaCYVMAcvHwa9fw3tsVCx9bGXtwT5w8dH
B4mB9oReJdnzkHrFVgK2wkwMl0hOj8gS8nEVNYWlWEWCKohWAX6S+4H3F+yT
AdpvCfoDfxtp7WRcuAA2+GlqNYLdWPw4miYd95yr0lUq6IHAxbz7XG9YVdp3
a7H8DptO4Nwed6nLcfIIZnjb3I/fevrXqqlo3mcnLotBGaP57cxsOVB912sT
P1FdjVnwut1LQYQURu1L9V2zX+IfrRLpHIKOWM8OxJToJAx+QsP4EeEeZbHZ
IB/Dy7/zKUKf3+ILOe7aBHnAxU8Jex10HKjkOrnT2mAIZuP/jK8TGj1MEBGQ
XqPpKrvfG1+qiO4GXO2biMxn0gMZ3RzpRnWNZJcTJCdUI7GIQDPV3ghusOYi
4O8mZkgz4e/bCN06h7s/Rg+OQgoYVYtV/LzU6Wv9eldDBVIcDAhzvWgsmcJZ
uzFjwLrskCoT/pjnlMKsshdjX86nIopFCS1U0/pKkrr7xfT1CzlixitV9Za5
4GtTF1x81ZW0OPzwmFiVymfsqHjJi21lc5ErHQmrlKtdWvUErLRAq2uc71gT
lXfPOxAhuH3M2OP09RE57M/qrhrt3FgM2biYNap5hM09PjjwTSz9gkxgrZd5
aSQAqjANLl+m9xdJDtObGFV9WR1FNFKd99Y691pcInVU1KDYwf1GKSA3BYcW
kGa5/EitAhS+80RLH2+ORF7QLYzR3q6TM5B1EYZFBdxscGPUI/59DiirBABF
B1WqyJAz6IQzXgiuOm4uRUtajbrFlLSUO+mGGQoDd0ojFJNdcz6mRR5Zni+/
aWlWgUHVyf1h0WMxVEQC0Q47Q8qwG6Yj9zi38SA/NAA7HQ4EvKeLxAetRHJw
f2Z1tXbEZkU8VLo5CBzOCv9uDLhQHU1mpmPPfdQdd7fAvFT3U1ndtxmAoYea
Qv400ScF/nCXFDFk+tOtSRb/BhV61f2+L9pxuEAQQYsUkNl9j01itqfP89/a
5hd88mMCm8BlDj0+sn/ie9k2bjSXE1lU3+r06Eu0ZUFVB5eSq0L+1wUSLkBI
SHhnAFtd2iLOF3VH6K+2gW03fXXU9KfiHtaNFsoTUXyUmBK9wbf5rL9klxLR
mi1CySCEPywoN1+GJ6qFRhn3yr6JLcUuwI+L5uVlJX6fR8CdYqvt2M4n5EKK
NSGbSWX++s93yM681vP1yQ52u/7P13ZD71KlBsGjriw8jE6FDUgR6XaLFYul
Ju2W6VxMob3HoKjyzN9qqZ3qr5KQ7K09CdrfWB1a3diH+HHfnFUjZA3yh8uR
PnSp3nZNQACq0ru2/IlF0vGRRxDM9s7xP3lppuQ5pufLx6KTBkrdPZoeImT2
yX2l15/4NytrFRZiI08NCouOHWKVFXswrkswAdf+udZs1TS43vn/nwVjL2oF
HSJz/OTD0NhaIyN70yb8AxLd2nmVUsuR2J/6lnKPt34eLISAFG3Ygxm7uBSJ
Uidx+OAKEy3KZD4JqWJYRMyACKf+DK/n2EFDwuSoN7q+k/vWilApLYAMd54o
V5EVzqWxhQlOZT+tuQRL9BFCLpFZpfwHq4aeux04/v3BhxB68Ky0HJLSaIyE
Jbtc35UFCpw1+NWXvXG/8YOm4JdZESyaKuMBieD/hGTviQmp/5ZaVG7EnKOr
5n2qzwvjrWIvqdwiC2KTkdEJb3sOiNLx7eWZAvsJ6Gm6i5mirU4TeUSR5nwS
THGFdKLwrwxZssXx/RgUQsb6vSoa9zf/zUSd+dQbY5YtJOj1eC43u79OnYuZ
3hDeCt+wmKXxG/6Fk5ghYm15gS5PCP2vU4fxB5K8LmBtBiOX6cOUysWPVSW3
a2WmLPvooCb/yDxH7PJmXMjfvdrwpM20NW+dC7RcOpGFphUBT+GJ2ogsGI1t
FlpD6BTLkAYoPPu1vh03cssl4/4ye1MQ9/MMf0T7X7PjFWEqUXoDwExt73Vk
wkeZqSl2yWqDWTH5YztYbreTLYRMUO0Ol/RoJ8lloOifVRZkNmo8DbGrcrTD
pxR9BMGn9KlQzh8MTEWxcrx+8YF6YQTfspZVPhKgQdCaTXatlzNCl6wVkEPN
xBBVFjboUl8bOT/QzJ5CrDzzLJkX6QsIuFxkYp4/HLSFvcngnjTnrG82Dgz9
H/KCAQN2qYkpqs/YNzFS22wABEh8nk6tZp+Ie8qwPwrRy6qkErNY1f73mwBt
DMhg+bomfcAhYBKRk8bGqBWZruuGQONsSjIEEXXwDBT4A9G/cxCjkoahLo83
vuRDUzJUGZuMy+PeM2lrRyhXC5WzS8JpqaBEGVir7gj6dqPsODwNiw/T5Mp+
wHZr21o3WODWHtL0WAWxrfZWYJ531DxU5CpObPVXklH4qZi2S9AulyZ14jPV
KDSp/ojwYaQctzWIgDO6FgylC1ZybcpGLfEc3PXT3PolpcxHqrw046RcAh1c
//y7DtJ4OIpEgJYGYJfxeKA8XZ1Ha8O+Xh95dpSeFEcKI5IjamuRu+1dHntr
i/2k/juNruPE+N2snnBA4SUhSYz0ajHkYoSlindGu4qmaAPn9aYh0Mv4yUUG
I4OMqYHiOk5HzJP5RvWkKfmGaPcPrd3I83uqirYb1P97rbx3kg/nuZ3DRfAh
5G6ND+ih4GIlJWNGjNRofS2Gam6cPUZ0IO8vuZudBUzIsFDxRqUvaEU/TUKY
xsMRS26+ZOcYbXjJdzmFdEkUUqPjS77cLhE3O+A4TDEzGj4l4ZYJ33dEO514
ikQ5U6VwveqK9UUyvm/nLg5Ngkjg9BJu1g/V1JpqVb+55In3mKozqSyA7dPI
efr9hzn9/IURem2mWRoCBjy9l9CGjuJ5sCIP95ktFISWGthtB1v5cBaQZbCu
nOxasNfPfjYkvzd2ZqXRFEt3tdWuz5Y1z4Sy05cU5VOwF7+5C4jF1qph0BVf
ail4K7f2YTUT8GJC2/Yj7ZXk/Xo/CG5JeGnr6Za2qe1lmMPAmbmAHnzfbp6H
chjWv3RvLp+OKAPw2M+DBeX45lHSGyM8YhxT5GA7MNRokUM8y0YRYD5GRhpM
vMx87n235ihb/VZj9b/kgg90WBc79QozbQKEHbSCCT3KtEDDzWQPyRMBH6+G
3QvLBeby8n0/dkE2PvRG9HUCsMMVMsGphfHtELEo/mgaVg7AMAqVlaSwJn1N
Mbw3GvLmRp3y9TsLEj6WDqOiA3MVB6okI4mjA6Doln+b5rnWqlJx3S1Q4E97
kJiNtwUJPz5pxNkCV2HX209xlCywkOryImfB0Sd0RoKeJlCB1Z4ayA3DbPUF
g1hFqx45LjpdrBr+YG1dkZrtA3YA0DZBtbwV9lw2wOhbNChaim5tjmGQCr6e
cb4WvdtzcRoQHjU71BgQzvpqMkxeIs0vKjp9JtTVHDgKpj2zMxnkhTct4GxN
Id9KRPVxTYzGWub08K18Avx/qtI98OyTZoGzjfbE9MB74hPrXJxRCtkcuy0R
2T5oP093u4d+V1d6ewB6IcLDqVnjIdzMsP0SwUjsErddhSRx2roG/ZrDEA82
lrBODhBgVjP9TNYah4rKSQ5oiCXwp9FBg3Rvjh/8rBOj+pdUCCi0f5kETkrD
gzmDTx00Cnn66pFct5Kdqs1PEwh1jGMFGMZqt3Pn2QX5X0QSLhUA/L/k5XPx
SPPAOehk7IpPxfvGcaMBCxXP7/hTbv2F9xZoqSlXrmKw3dRfhnDQgbAJp0o3
aay7AOoGRupb1PecPbJ7dYpC+cBwR97Iuz1h9YCL5a5heygvLBgOhlO/QXZ3
qz8threZv5bBUB88GojdsyOlfPJhlwo3Bg+QLrlAw/0WeX9t1z/qp/FifoKL
gdijbpoaMP9csGeHpjyWXsT2woboM/IZoThGK8tKD4rH+i4Esr7UUl2IOh/R
gG2lIu+cCzUL1GRPTbgYfVyA+XZ1QSqLMrXloeWAhjbdD/iCB8dWOdkYSZj1
E6AcfaR/VvJl0RLj6GZPvUSqZqvhdZdq0r/IPEZmA/uO7lhxWnxAk+zbLVN+
UvtngrQLlWaOyTSRvzbCyJKo37kotgoCjciwzEjx8lsbI/LkPO6D9UnlnQEt
XC4rheMxlmeUh2jtqYoe7VpymrchwxRC+8tlu4K+p5BumLA/qQzISHuCkd1t
rpWjf/d+alU1IPsF2iI2lNimihTUppI+cLMP+dtM53ihZYVD9mtrjVCfs25D
WI0R0YjuF9EmmnNHXyHeqMlc7iPXHSmyvfuJxzL4Uo0RZl/+C+Zyb6ncduqb
bOn4mvg/pwZ3vKMgFlyGguc4IpVEIwsN9gQyAjqTYKJXSCX+pe+JNjHdXYj/
PcLmAbhhdld2K2oiiFtK5gPKn3UEY9L4big3cYwm9iDn6THJkWC9DrOHirBb
O96MquBpjLr9bKwR60pdW8ruzwe4EwmWihmI46KC/lk9gewIhTWwjIMMzBJb
887jwSC6lHQ4Ejk6DGyqub57+iQulu/QZgmyQdS/tqPDyPmDOHSP3SztcPQ5
v3qhZgOK96yGv2+xjw0TzYjdsS/Qa9TIYDWdRgNt1P7PZkgtgZELbTwKO8Tl
/m+T3gspplF5T3k/B16kmusapm0g3fYESBN25vEHodbwzdJ3lHTHct1DYg22
TgjQyUGAWlk1RM4W6tt6oYQUe8PmPis0CVQgAHYrli276ENQn/Pu9diK48hw
xHB1bD5Z4Fqjy/lK4mx38oTbZapl0TM4UaULUPKsQraxQ8KX3z4gs/8hGSeM
6m/tUEYECn9swmzuYlEb4gVzY89+9WGHSS+GzboSw7Gzw5oeREHaM5pK8WUS
70RRlfSqS/ESue2r/DWWjotaKfjSOy1W2+/OZPbd3nzPD4CkQtgmfF1+sKtk
+iKXIo9Fsga25d46yC+8lBlUmK3pC6lJvUXvJwdvJgzxV0Y3FC5vEVBzxW+K
B9gnu/5sysYp8A3AuW3E83v/E+iI9i7/UoUaUwG+BXtFIK4bW2i2jhr8BKmD
9AyDourfNUN2bcV2ppvqySzJvUl6dXdSAE+yf7P1UGk/Qcp25NDm2WI/ZqIu
TNJ+0cegAsUlGJjuTOxxT/3Dkh4jWlr0Ilf/cKS4Ab8hty+UhslIl0r7kzQT
6Vbpv+KpBmXS2Spki6P3LkOuOw5TU7vefPw7EKjJylCdi6uPgxHtBrnbSn7H
2nHwyTL9fsHA3yGvhR9PbGq5XiYzuso1eaa3jsQHvTaAEBlliR+Glf4O5BlU
KXhT+hTI5yp2jEeZQpZqmlcF3p6R/wUb3P3Hn6L1Xyxy6ixFNfEUxEDKOSGQ
UWcLxh+fdgKaDiBi8GjobrCBrGFc61X+n0fgxwfz7AjREOYHjvv1t03h4ar2
lexPmQ78jX8KpPk5FdFtrKtB678xM3jlQqklNx5AfTwE1GsH3IY0SY4CgnbN
lmF4R+x7zijFAwCe3WQK/otKzti6hYJnTGyGMANx5puMQUc2QXuV+x4pxISy
W1o4ov7ASyT4xe5fecSSHlHHuFyd83CnvgrnaZpzgjaknCwGCFlgiqjIRPUF
VoI4NHSwH2/LtTTMiw/uQPuZnPte3RADtpAPT1sPEuGm6mBxo8SEOVjXKUSM
gC7juAnACaUcz0sj5da2ebzo6iOyhtyi48cy8mhPB+72CWelQke1QQmHnErO
+rIn5di2343IJlQgx8Y4gK3qDMLVlkKAy6hk3UMUp28uwUT7sNPYKCBkofbx
GSyjBA1EVzjbzcychbtRu4/Au0kOzgbdzm5cwWZc/lfp7Jc6JNDYL9liJjIY
645FvyiuvndRpqd/HnQEDFVCPn6LiBXA+ebSyyc8a5287WX5peObEe+S5ZjI
WofTM3voDRcHCwc+L/ioFpmpH7gG+IPp7gd+d3tyvAxmezE9IF22EEupADu3
cC8L1ENsu9dGDhslfZhbB3/ObgJsnnM98StCRS9nWbYqMr7cObprf1Wcjsvf
v59KvWKB3bBOMaCFmp09cJB0GDa3re26zOtQaTkybPQ2iltB/2yL4CX0Fo/v
36TpGq4VVOM9Ne/9nLBJJM+22bgEbHqaOieDz3OwCq7yrz2Qy0CzZ6AA97al
+PGyUkfCDd1V4txXAK5ohPi9EJl67UcjCwmzxo+twsC3IrTFFfXip+dqMtlG
Lo9op47RgUPeTMzHmFJ42bGGYQ2mHNxGnGWhAvy6dlMMfR1I8ersY3XvK27W
Bals5n7eactWuCe/pl2g9kuuj5/kkxt4YzOg2V97pmW0y3/KnAuW5rkXdHy8
KQs3ZOIC7LyuSdxdM0T9Hue/Jwh8d3fLIPHmGJRLeiFQeU5IC1k4dhJTkdEx
S9T71gGjDy60MOeIylWJrNXS0l56TU92L8t1AV7iC2MxbdY+UrNoA5uMwhKy
QRGdcSxa/DE9NP+eafK/mLuhLRfWeyGHp5V9RkHwgVC5dtxt/FBnslPNMOSa
F7pRDn7LN1mmDz6KFtrerCMtQJFHuYCOPkwtXt+72L9w/8PEp8f9SRKtttTI
TQgi5OfCZJlBf2lEr5zij4H5L1V3HaE/SmDX5Ao29Byycl2NyJb3LLZpEhC9
hMPDYQjQ7CTebC8SB+icvWfN1XSreSpEuzbN3Wcvv2XbqbkrNb6+lJnxw+Z7
3TfrolqekFxty1YGpsroc4brl2ZMWYTqWNVbkNxKh0AKp1qCGktZCe6EfMd2
rvW0Us9EZ01+DV5+nAyNojHKButsGcN95E4hew/d/tq6PLmLXFJ+qZOK4M4H
tgxEjtoEIk9avg1mYq20XLOKxH+zX7pYfjpL42Q9DMCiNFLPYDNgeY4VSxOx
BK2heTY6gp9Lop1RONPT0NgGlYj/l0ZiZdF4W5w555kgDDnXkuZrBNpUEarn
mV7wEXWhVrHo9t9xDAPDmETMIayHCETkDi849OIfCKFqZk5A/j1uTUveq3Y4
jVYrE8fgauB2BLECgYOgYB1Rv7sT3NlhTkbLv80W10bNN5LBt4GHokZquS99
eHTm+Dui7IujJ/p1RuKiTPv5hlCUjDfQt+ht/6jsrrPveiLyiyNeqm2TJXj3
F+xD1ndRtvE6Qu39xJfhoxVgJ+6aWXZzuns2EGuJDqnBjSac9NtLORtPOkD6
HihgpVSoLAYdZeGTYO3rmihC5UFbM/03Eo+v/ZOk6BUaxec0s2AUSB7/bEb5
a9OfYQMye6yWr7kDDf3XbU6UNFm4ZYC0ry/sJ68fQorFHR1krrWyGiKdNPEH
RNqeuIBwKB1EktBcxQ+4KX7apD47AmNicdk59zBSaMLYCDKLusfOMLbhSIUU
j1RUlaTzJbhz3j0NMKowMiZ8M5NkAxTM3iuw7FKV9k/j0scll1JJAco9p894
CEI3BGt+KDJlLy7cQ30rMs1ZLn4mUjpz5QNs8nMyr4tiLKYs4W8mLaCKhU9v
aDvzXuGXKLkXCTOWMRjYA82fSJ87AdtcxDyFN+NHVgIouAR2gdX1P6h/TdN+
WjEtekRedX8YplLMfTVjxTsJ6GiS7tgqhU/EIPaPsPKEvoY6b0LHsTGe2It5
4U99DjgMTPyjsmT0tOmojFAJJSHmoCxMMb9TEOLiRUQEP8B5mAJsJWcckXS3
VfOdY0j7drVLDkUCU3zeeMb5VrWA/yehhfOE9mcSNo2v432is4kP4xdf/HL4
vLNoHyCw+VWYAUZTJkZcSdOOWITAE/5oG4cjDUDif7XO6boeQ44zPEVlMcsD
yEO3N4N0duhI7xHfX8lCFGsgQCZCMa3oC9q2wRfZ3K7rSTK815cbk7Lhl44X
wXVQD45BbbTbDI12iJXRTDxfLPe5HVwv3oD5OQZUT5D/z+/qc8bzfRapHJrZ
MBW391qdklH5AjqizfFRHYZ6qdPo+Sd5hfRmo7IBWCJo/ZDS4ImHWdxebY6L
QkYqE9w55M70oPMlJPD5WkE1WBOLPFaaURzaAdj+UWrBN8THoKhVfFak3M/+
XcRu3EV3yPsLLF+Kb/VzgaCFVG1n/UXfJM8s9MMkJJWp+Uj2VRSbu/eLSBvf
VkbvWZ6iPhKZRsbY6/9t5iNybS5Xqm7LTxg4s2OzsQKh3mJfOzs1xwyXR2+W
V908lplLzvWwbeVcz7wOl9rgokX+i2o7RfIm3FF2yCYljYfcNilVkecQkcC8
QR+bKgprbErif9GC0YT+SYTV9QLjYkX6VyeFo+d0MsPy0Zj02LJkfH9IYvBo
9c/Iz1CgX2UpI5GDujYHdgeoZ6Z2w9eO2PnbA02cZhP+Ed7lckq50BUGYkjg
EKd+wZw0qMqhbdwwpNd+wIbFG35X8KsQN0sIaJwZSF318zkAgAd/LjbUufvy
Ds4RIwOrBrTL6iKtiTCI5ClXNbOqY81dGYI7XBddkHmbLbRFhSzjCzP/s8qH
JoYYlUc223sH3USk6ZpocYe/fa4mgbvb/rhAe1H35UiCsmDlwteqwWYuAXSn
pNdZftmmYtnVxwHPIMCzppAGxZzWENw37yGdV1o4GltubOi3HpPldq2uVEIj
IStUbYuqQlptEDfdv5PromtATWrt/y6hd6STnFtWg51yeKI0xYkmsnPuFni1
W0QixC2cwJXWu8JPgukXCDzKhQRZpHxLPPTelSCjLrVgjzMawc4z8fswdUPl
OwZo3tmxjdrqf/ArydKgswmD+GMaIV68JWjKoU2V4yucWf8X2S3T+2Ih2Htt
lUpicC3DSoNAVfVwtpUwjY+vL5Z8F9ZGCNK5VZ6UFu874xXLaBO+aPMAthV8
jOVAesNhojo2enAZxEd23T/v0tFHNGIsxrxPPTw2Vwqn0SSzIYTQEnMk92hu
j4upmW/H8su5/cJd7/alAQjKm5KnKC3R25US1ofZCFQ03wMwwl/PukIeo3hV
Ff6iw9neuHUvZ0BFusLMBRPz8SerW9hOXu63d5Y/S/7CZBkQs8bZ+wtdjKCH
mBxjoIe5qaIdm83ezbRXzGsvqSx3FC0/6DOC9qgLoTk5E8UKwSXx3I0gTFTV
6ghtorvg/OCAUp3yDiZZt+eHUk5AU42GK/6+JgtFdFDQ+t04oIjALCNzNM+3
hicGog+ir7saqSQMems+bSQBHru3JZLB/0DaJPhHu/q0kJU79BpfoweS6oyG
nEpsTOSKdakyHr3dbRsn4hxAfEyL1ROB4HvNcr345Rtm1NCuJBTCrpCW+zG7
jMPm39V7eBWGzP4ysXPIBahES8BcS/XHLbBdNyVVZdiGO25nrjmjdvfWzX9o
AKkx2U8vP7fE4jxMCAhHYgE3KI+cp0+8P2PC3In+w4KFeB1+QK0MJ0TxRjrr
SgcBSGUBzSNlxdc7a2/wKb9uUpSALXxl7BssbDyWB1K1Q9O3N7cv7O+SGvtR
qJQSsbTkIWdGn4DO/CUQtCBTHxZ7bJf2xjL6l2OUeaX2uOZzxYVW5wF19jdb
VyNZVf35rxboDlExBgByjUrskdp/58iVh22bWyPGX82z6JNBEq+31t4gXdVd
sgjU2gmoBqCMiWsVffRAXttcRslgNUBZF75/RFIfhLxGprH8Xl8we+fpqtIm
as+/tUTmD3q6UapyCRQugN6ehN1N2A9N74n/sPlPxAeywDNOfzyX37tY6cbx
ACGOGMvWpEH4Uok/sZS4Gtx5nSj86L86kbpTi+qbP5yVSUdO7ivGMpaazkWJ
zZW61OYw2KwaIlrvarVYjFjPtUJ15eiCOctAcvHmSbH1ZF1e4LLDZgsMkLhf
YwmzSrwISbxDPp7i5VXwKFV9He+uE4SUuNBauGYgkdsziruAk6x8blScejor
3MRuQPsgPV30sr/bHE3bKbqqPXtC7NYPcxsa0sdGTTItihRypsjg2JBieRcz
sYz1Fhl6h7C15uS5PpGJ2wxrOXKib0XGT12/nrQDbT9XEZJkcYonAeDRjolg
IUIkYc/HRgDzzrBfSeocCiO/XWYM53agh/OqzQV8CEl6V4bLJp1IR/6eYNUe
tlJNMIHdbr44f9FCpzbFKhUrN+xJoCGmHhHRbraGRLrx6BKVZlulxz0kizlB
4HfIln25/sboIA8gKfu76PO6NiKMUr1Aw3WyTzRqPygcNvq/TDoeNMLxOp2v
BM8iLEs4IjPNEGahvwxcD8zWfXrHq0AP3KQB5g22Lw1pjEObWjGWwn9eGBk7
fLwCeYY2jN5sgxCgLSiVclKGZkOxbpl17x/kVmA9INX/+OhDDeQWzxahKj9p
uIP8GrjdZ8LMIB60ayOVNGVMIyRlteyvHzHHA3nWS2CUnLCsRp25BvgkNLGh
HtLFBnRlvVKolI9NGU4PUEVUq8UgbD2/VLTfxybe5kI4ai7QyR4yaslUd+Ln
htVRs3Ca+rcIHsDR6n7ftlr8q+DKqhGnei3vMuY4K2C12L//pA+xdjYYIx1v
I1J1QLCg2ROotm009W5SpN3Ic3YmT4jOIKfCVlQ8H0V+LCEU7V7o/5PqR1R6
hVH7kKw1WRF5FEYRbzmQTXiIycz6LjMJhkbrL0TD6dFUfoI6pIpHwObS7f9Q
jlgmDGCkyd8fsN4bwByFTWY+ULuw/sGExThiLzW7bRZ4HGx9UzylIw311uEg
L76ry62B7Gs33BHdTTT0hcGVbQEeCGcQQ0BHKq9/ncoKToX507f3MCty/Frp
YWhcohycjJFI8s6zZOKStvkJ99Sx65IhluXcJcOh3fQww+PoOB7mIsJZju4V
WK5fToNanuLrzd5k1BmgA4Dns6fM4IcO+GokSmVsnef3c+E0fqhwiYhlt87N
lLHIWGlhitwzy9ldSkFTpmdWNH9Br1swzWQVFmh282PnWZRxAnHfrxlL/f6z
fS5ZhvuiDOVhXX1/NJuUki0PSv2drZt2HO2W0d9W5OzKGZ2h/v99Ykrhh0sB
EBtEA64UQdr8cd4UdwNjMz0CvwWcBPbiN9EKqsrqU6eMbg6vAP5he/5aB7Ie
tR9QkdqC9JVn+VFTNM4k8py7QsZGuDYGNnsJKIj4wTt+UvRiR9RqewRvDOwM
3IVxdL8onhRBeRvCXZlTc5D47+736ZPIvYYDdey8ZKcJ1I4qf0p7ZiCyENBS
GKtUNb0a0yPSR/LOIMUIf6V7jX/qNfqBapfXsrU/fwzE2JMLy+uck0+JLhR0
T8rosVPdBl/8230rsuywRWnJCeJKwbKm4wObDwXikm3xWpaSCC3/+bMy0AQ3
3jlCZo1Pu8sFM1od6j19NtiVA67pmIzxvt4qptS1qJZZsdrNVpRQZTPWLBQc
nWJ1spQR8kk2YfCybhtVt/TIEkgt/RRQoweo6ebaymnXdV0/LCdkuBdP48es
/NhPoxtwWGGxNZ5t00cB3HgRCBV0sPK6ogFVqOL8vp3u1Ut2yrg8kxysOzlm
DIbkTQfytFV8Ez40n/wZ6bKvsCvmDB1UEEFxhvdm10xMMIDS4Q7S3msoFL21
Kne0PDjffB4b+2nTSoG5bW93SDVYxycxpUAps5wYBAbw5nj6UTe7wjMEPBUV
cMIY05IUsr4dUV89wMxoLy8+2kdYkhnxtcw/YTgBKpKu+BvpMRJi9nBuf89j
Jqq50/L2Z0PQMk9qwh/Ei7e7gN7XIYI1798d3qlLjLpr9ouHnPlEYZm1iQcJ
pxcT1ZqguwYeOIncimERDYhGZZZsaYoClr2G8A1BBmldXHZ/gaORm13KDxtY
zbN+cLcHkW8Ovx4VX6CLZkgsTOU+StziM02mz8LC3jGa9afVCtBgx98eUEos
8baD75ZnFsbegSZuxffhFxziq4itIW5G1mOfGOSQ14WVYDAs+4HfWL/Hzm/K
sVhs5LbSns4XqxKV808nVU3oynvqzzEjKMnyM0O11TiNRrajMMRiVeONgKu9
b+XwmUqpKiuyRMCChRv7aXXZF6zhvxCDoq1UrNHDuKzZNTc77cp6IR9ET0I/
fZIBAm2J4IVlbJxk1QSeRq6Kxdsfq6vBfNSqWzm8uYbdRzr1mVgpN09KlTMW
ERKFiR/Kc6uyFJ7+xvkudZPj5NJVQM6Awyr0w0utQCl+n7uao6lww1vhOQvw
pkPOAyZu1tDH2f2YNKZzd2dNQPSJOoFqcs7s42SLLBxN1XecEc7MtZHbHlnn
IgaAqEpX1c+iGsTkXo9RIDpvnmSRRJTqWHTYeVtT8EgWrt1zIcPCkgVKUTQ1
bWdA79eWdnIV2u4OsOks8tOneHSH04LWH2k3y3+2Qrr5lzhF+GzyMdovRNmr
vfuIJicFpXu4bnplyz5bXk0CCSxy9ap3IL2hmsAfmoOEjXdxQrSLUCcYJuzb
Acv4UHD7cRymcs0YlRa0hxPxssKvNUZDrUoy0oWhJ3KNNYn5hpx6mvMYs4F6
4yCtbssLWNADgC0FsGXOm7se7iWZk6Nt5XVcICtm/QfDvLsFBpL0vV0crS/n
NShJB9HRJ9cU0DfjjwTTeMrioqHigOot/ywUdAiClBBCWxxNMJXZAv8zJpJ7
4AS8v33TYo0fysnLpJz3CfOZ17ThflwFfXQufiCv+6b6XWovi5Yk22AvKwVD
PW8EYJm5lap0at0UDcFh3a8gLGXsLjSBzernUesojhcUxNtzICmkFhdiQNnF
gueGQjBxgSMRT6jiX17ZJiz0mMqF0gW65Go+qhkMoV0rPUxZ32iJVRq0E+LR
pP9/fUCKVziM8E4zM+vAo1hUOYs43ugyzg142IQ5//dhvTVA96j3JtpySqLp
YUg126Mgk1fMaHWs/d3lOP9aJxQziUkG3zeg8edZQvvSnMZDTxNwW2ycn9MD
+TzXWV98VHKVWjkd+x/Ht27UYQ4SesSHh8btxwrqn082sTd5dtylw6N4L5Eb
IIoA67lennUca4ZS7Gy8CAYErRHQdsTdRleQTZR4+jDOcIjUisx4dWbNo4wR
CYcfYtDFfBFyRNXLpQld/oNxujtEwyW2ZJS13qed4VwmOxkkPNy5305c6jKo
bBnxsURkHPVtR4HVjfmDYOjS3LfgqcsRn0n/+M1Tf6eb/1mcB3dP4VdG2xgU
qL7xR3S3yAE6C2lJDaXxdpCyikFGSnTbxDAYbhwZVQ93KQvoKHQktvQPC0vQ
Huny62f43y+j6QP/m6lmrn/t8Sl0FIeeRdog2Qohss6xgLVuhevOKh9y+e10
xyYNBDKM+WmjMx8bmNSC2ORtk7f7S3BJFHXqFcfi72sWpTM0ewanX1ihsgWH
XKsprdho2ai/zFPjaGmpfPTk9SNHKXeWGIC6GmCHlOz1YTIY3fiE0u+jmrfc
1hmZzOTlcl2ITt7rDBlaA40lHKLpqRZ80fhqUroRh1X5kKiB+ZMLn0q236w5
8c4Ad132cnEViDAL0Lgg7kDD2u9X7erEHbkvobeTyCNyrhfxZfUPFsDy8OIg
E4xPETLuY+20dNoy/q12zSQAcyoz/N7nPV6QYvXVN6h/V3IZNIbjLUh4tbkF
L54+BDGHomk8wWjqAdGwe8T5zWDWjZPYUjgqBWr/FffBU39zTxYXodLgGVHR
57sO8MzQy/Yz5nfioz2Y9+bvUAyYmEID9ks2QxeDjyfdGbvLaK6m0TKAkecV
lAOQqERUP8/Ee3dfDi3A7UTiKVhjBoAcL6ybMGUb/NCvEHunMgqeQK3lEBRY
XeYaTj9K2wdyFpu3s2tXe4ZR7MJu8cQj5MlURUZ/nKjCBtosKx7vT4MLl9It
NwDEVMwzVEtTybIolWONthTTkNaBe5mPgTgXd0D2f2VQfOVirQE8YP8piGlp
ppR4IwL601486pX6guiQ99YZ+naL+3oKfhk9NlZtKhl5xO4EL1ip242ootvw
PfI6vdZYX5lu3TVAxt3u1Voxm90deAWPZm5KhDxxVFlFAClL0an6aUGNmdPI
F/+OtZ71wwU4ZEPolF7hI7uQgqHIelbvpnGTxrKa1/xCb1kAaKTXgEqRP61h
AXBu/5WzrGiHdqybN1LIiLMC/tnLHG1tlVJmdat6/OHG3nvZzdavSstz2vEm
Wz8PBBwrzbClq/3FmGmVji6U89vsEbZkCI6DqreJCc2kJrFz82E5irZhRA8E
OhwLHoZtdu7Hu0lgbX+uJ7EYoixiHi0AEjKzpEKXYtBH6C8ybgmXT8kUC8ne
Xv8rq+Jks/cfXTo+GSfyX47LlcSzDpol8tpna6ih6i8KoXqrfIaMYFT9rH6G
TqtntvdZslp66/KnjugGMxI65/yjuZsWtC0N2NeTl6Dwd6pRYDgWBxtkAKhx
exGuqLQbj9exuO/6Yinogp7iPXYwGKIUqGyAUBudNldFHVia1Yx5cnSz/DJA
AghNsC/5GqGmET6NCEx1mu33FsrmDmGrUdPvJcIMaI9H7JnM+mr6mJB/u6HX
bAdVHoa70+p/xaI0BKVPg64XyrHMDFBKApdsla1KPPodgjbVhruXTM8ahAg7
t9h7aUb2JnHBrsxBcsnmR+1emQVPBYQGv5U+os9rpFln3EoUq+fRfZBCaydx
NlrCn+jGe+wegeNCRu+cRITaj6O9MPjpgZgsSBjwH4QCjI7v2S9QmlVLsPH8
yvr9XnB3ZuNJxTc3p3WxqgRwUR7MgtLRXCb0O7I/yxRpdezoLke5QpJoxPZU
q9H4cpX4Ga7Dovjuzp1geeQAMwXMOF7Kb98gGv+z4zaGB806tgE5Dr0yuEqs
MedUTz88d/S0QZxW+VePBWqvp3NxJAHAClY1MMCgZWSIpLsKI9cC4IkDJqS4
QahTbgeIYLAwuA4pDWlV3AX2Nsgdej2ANYLV+HE/rUn5vp7Ho1H4hmudjZIo
K+dS51K4B/fXDkYQz9YN6ABCwkzTgJQkseYOlHXyj1KudQvNpi9g9w0AZlui
8QhNzxgxiZvSMAFUzban8U83231NzH+PY+ayfAoT2998TsQFnQyoxVpKhP58
RJoI+0Y6T6AFRPhCNucbNfucKA7BOtgxG441APJs2Y8LdS/Q1qZSnAY+KxNf
4nM8/qW6Kw+XoxB0myeV0BVYX/IwYF8i1NIb+q6utVrUXy10P92gbuLMg1X7
NlRRNVJgGLC+7yGCHRvOcCLfsF+kP55PPmgxn5pLAyNcmp9SilityzI/JHmJ
bhU7W+7Lf1rilZ+ch5PNOek7YcINkMrxlhjkBEbifN09DG9f7tVV0h65EvTt
wU2SQkWkt7dq9sOXesDTaEqxVYyKGBGPSn0jcHETrZcsufKsJqiVlxrn/unx
4y9ZbzIeYkvEKrpSm50Yj+7292mDEbEjzia1DmUOFkxT8ngMSJp5MRWe7lhR
+XPIKJWBQd4vSdxsGC46WY+egRuyYkKAhPZriaLUDKxmmCiUymG6sZQbH+P/
XnHk621PW5Gi6rP1DpTZ0rXCPaMe9oYhQ39m1dHDVf3WdU1iJ52gO8vBbESa
8UqsugqpWlCGZhrd2AiwwySNFkTq/IoUCUea7TT9gk0CT0yXtBWhh8yci6Hi
wuGvp9liLWWuMdcouQUqbjbXMu2PkSSe4cbvMWj2gr28J0foW2ed9dZ7GpxP
ZI2/k9OarzbJmUMdG7XFwcFR8CguQHspOg4Sd7EnbegpnaUNaFY9rpGm66mX
T6ZvWY8pr35JIqKMrl+w6ktwFfnWX8NAuxHfi0tdNRk5lvwAyqLwzVIo0tc9
0doJR3rfYFuzu225EY+OSNqJ0Wbf21mgLEDa28OIBJaUlecGZMk3zZMGUhoi
Kd9qDxwbsVFtAzn/P4zNZdfZHY3kMkvrNWIpLpb+rVtvByVZ7e0NTx8piELF
jsbDT0hm9IA8vzpF/JX8mgPP+TUa+wsmwHghQ5DurSoKmFKC37xq5lPfJvya
0Lqv1flAk6yNNzbOC+WKip5hCoQkHc4VOMrSEKhGWmFRtSpJpg2rvbJ1p+uT
ssO0hgai9/W246p5uALHbvIdTf5I71bN72rI28wRnuMLUJvUMX/brxcWnnkx
jW10sV+hq+C25Rgs7C6B0/TG+W9DL0dh4WhgOviCz1HUvTkolmG0NQfetvZY
MW0yWn0xeKdx+IUZhf0qxs9Y7ZlpxSP8yRVqISTTU92qstkP12R8w7DnAol/
AsNLrad6hj7cXSTuNjW2LPrm5JKShr2Ijk2s1YjLLIfVUcXXFQZVD02jjuSA
kmM6HCqDQmB4g4+fATURmqDm2AwX1WdozIUhgBSo1alyF1heofMhil5nyEve
VMiM5LobJvxQDWwdVHVcbVrkL3ILB7NWl6a6Dab/ugSmEZ4xk4ow401i1LAa
pOMhu38mTwhtHHPozgw38Q24j7bIxbMKQpz8KSxV4ifVPztWGdDwdfM/SV6v
nd7P3/4MgKQfaUTISjtv7V6HMydFd5gxq+iYIY7xKRELlMC7NOsVGOZfdrE0
yN+QaeC280p2XDRbIOs66BE3FaHH7op8ads/dWMh57tyNjKB+Bk7sdyDZnPx
e3D7gOhq3AxPClHJmx8flmAHOaQlVfGHB06QLoCz6sn4yeYzadxjE4fPd+J/
2DwKviX8x2CdbhW5aOk68B/574HB6yRlECHaHeUXh2CkYqWBMkMkG5I2MB74
2BtuG7h2/Z2hT/UM3YFxVLb4zaS1tl5jWe/RiEYx/OaofmGSjOKMOZeKAZcq
dz3H12Y5FECzkwacCGjY4DN+5zDEXVuSsGgUwc/npW9XC4zVavW+7Z4/0YyE
RlrI1KdQ4NS82oVeY/9xONVFAYF+tLkNrNRpTTs4FOCExzZT4et6Bs32S91U
LPCYLpiTfO5Vx/7gehhH5vLQgfVOj4EhE6Tzugv1pAEPlY5+GX5A/lUH9BjZ
bYzHDwWDXAo8YdVB+n55amhs3r97NrJcFJWeok4YdPlIo11aqRat8GlqtOkJ
uTrgapwZaFCm4ZlRshchTpoaz5O4THamBTh66N1OKB1Nr6Rbcf8Kfy0CNJZL
e3pkwMe23hatlflmDCmiee8Qp++22gap015kyL25k9MM0Z8lMzbMoTPUEQQj
WI8754EU3UuiUEJrHV5jzNUJFj1S32Uj/6YtrPgRR2Ybuje/m4Y9sChCG+8M
LVuDdj2x5euum0RwWYdoh5UL8xL/DxYGa1i0KcSs0zrHZ2P+SGtq/FhbgzVf
ojokYstmCuNe9HsN+NnnhzFTf1NvoFp/eTg1Q8zoaEWhhXooZLgDYMbqXiX6
qMB6GFEcoQZRMOjXHLI4hnBleFWIK0YolFsEHOlrKWauiytUfK6OMpbGg1BP
nQ5TU42yyNp42FFHiBCmvdJJxHhAfig7tX199Vzx9Fk6jpIspqTDiOqyen0l
VFYyTDtSH99I9z91pAuO4cvq1u+0R+X5Wm6BHEJag4/ptFYDvY7nJacUdarg
fne81oKwcn0Ze2BagWhllh5wWnxeijGc/0Rn+3akw4R7fljvz5JfT6GmtEM9
eRQ6RmnjBSUEchgdjp8et2yE8fMEouLTmNxCg02IODgLrfkhZnP0kno8a3ZA
Taou6nQyP8rb5gIqiuBIIzr6Sq5XKVn44uawDWWve6bWsfrWj1wD00f75vys
gpjm0mUG7HZEQ1XbnKueFdtByTMWhYk1g9CZPqUsO0MBvuKELNr/svpsMicm
B3ElVYJJHTPcIvJwwYhO+sGz1v1FTRlyH9gbUhp4d7YQF2tCPsbdzVN6R+7Y
gYT+9LTUyPbKfzbY9SfvugCt+ChT7bYvNJBdomK90tYNCfmAeCa8o5al0LzL
qufdBUylonx/hsN9QX9LCkVu4vkkeli2TgRuDcvFNerfxwLXjTU1wT+TM+y+
sAxnRPfAXYvFTGBeHii8oKVVVYgRbih7Se9lmvqRzs7N2llnF8/L8xoFmZii
AU8pzo2lgORbyFU7kJhtIJZIy4JNYKTCN9sNLHNrTm5PSseLve1WYrhUv4I2
DZbnn4toV49nSGeulhuTjd/4MdquNlQ/jn0G/d2bXkWr/sYHn/XLnj8a8JES
HoIwtKj4eGS1FOOiRCuHr+yp02KcDEEPS2QYRFgrnNziqHsJIaHuesWyTAqh
pN5wlztsM7uz8/gMPTgnRxin3h2QGG00fNi0v0hxv5UDmgOSns/+AphojxBu
Ooni+K3GS07rAst85PEt6rA5r0tByWtlXjuhcZAEk7WBq5xdMOnFHTlzCNMO
QYkqo9aKRhB87Oe4yoFDKDpQI2gbIzRsjr0SoaaDz4z2CBOim5uXZDnujOWa
GMsQgspR5QeIXXvkAH6Ry/EUynbF9496X//fgJj7O0oBwhbUxTpQ08l8avIu
IWCQaLUEMWiK5iRYRqAgut7qSWUaHrD2mWj4diBbS6tlqlnnrhSLqgTdE9jC
OsPNhbpS4PGzSKup8T2VQR5pUdkD11xLJcNXr3rCLd+KC/VMvb1/dm8iyqXs
Bc3ynBSamNmt1b5ODVeMhjG/eaTUm0kHou2t+RdxOnDd6SzGeYGA/agqFk7n
lUfkHCUFfM2efmtPa8I1Api0oKh/ODSjcRlN0NnQOvRE8Izq/OdRKrhjN0g9
6BlkiqBeHvlzdrdS4D1uu3h/ArCWfjiimvAQmbltsP2YiuwbZtexGzkZ+Ro3
if9n35/lszFdkeoTIZJQYu7UxCS6vEfQ5jBgtjsOQ/24N3jxvi416Q+bw0fj
EyRnXaAJFD1XLT4z1F8urlcWDv7y0auiJef1oqwaB/5j5X4b0teUGMnEnsrm
xhzzyIus3D50Q4KOTzFdZg90zK3/qVGQFDN2arOa4ZapYpz7QY9UR/1Huzll
OKhi0rwcL2UP4vYJWJkLMW1e337Pep4SdovTULffcCm3CE8INiSAVlu5CQo/
/yPa8izDWfj0iVsDC6005EohImUbfpaRaCmVtbDDQMy9qA0rWzoW8tQKfS8R
J8tO3/tF+mTAKEgKzfJSNEjHdRhKTKHbX/03WzSHgkT1SVDrvSKmHnWWvwB4
fNOz3nzjPbP6qMEs7ysZFZ5Cq7HXu7yQrDlSLFOoz09C0J6DU2U2UVca5ju2
5cHHdtY1s0BWP7T6JeX7M5+nY5cOmYmNTs045UGag7xtc988LKVdTqo2UjGy
CekoEcibYge2YgMac+hiDd2qQdM+ERBGQVh5YQn3f2MN1yWiV1lJvz1fHs/m
0he9OUxWQimftyVn6S3gTqsIjEi7gEQ16HTqT48JYEhr2zYy4aixiQKkWM8F
0W4JLVVYo4bSnFSAhHtpkVSWHl0cqjWL6y9AGNeuAxo4Oiro+2xQy2Aiq9Po
UHbNYSybEh09VfpStmJRlPT9gRVGyeIVdkbOoZVKnU9snAr74W482fX6yCKg
kRXG08PSbRKj4S5hPbHx2b9rIEUCDz7RvdRcO4ViKxA54Vk5O0dJNut2Fh/V
Z5TfH5fb82awKOga24SNoFrpLJyPNF+BUv/SfTk9ix/FIRTGORh9bdPJ6yGT
FkaRVMgHOpGVR1XN9xLGyuHariKEZSdYVFB+mxCdo520IdjfzrKOQ59hCR+S
w+C8c2oMLiQBadG75R5AT/4Q2kP/8jl9NYLcFRrH8J20dmHoj1Vs8Kf1flyu
cFWhh9bi7KQpuhhrgmkoR93OGjIVa0SEr2Z7OJhnaY0odX2dMHEet5jcJOdK
F1JL0ZjEqqguegSaxzrS0T6f0Gmvk0wBAXQAtiYaCPZkG5RLsVbIj/hO8t10
7m9W+z85l/1aDBllrwuYkhmamslQTgSGV7JrMxARDAYsUAh8omw8LWfs3YCg
aGTUGzdM+C0OAVaXaGDpd3rk5pdk0DG4t7oejttJp78BesgonZwmoJo4TL6C
NtdJiHecdDKsZGjZYWLsXWKCgLL2RmK4LokXKN4S3RHLTIjb3sdxnK4gfncO
1YzD7TtbSuTcBdCvoT7iklAZLqYgEmY278t1bdAYrsJ5LYlK0tPq/5EB2p4S
ABe4rVyoz7ZWYm2XU5F8qyJQC5b/oLDIiiiF9ov9L5uVtGMwOJS7P4bCxKr6
5PpchaVaDzjDKU3VQWHc01tC8MI91GpZOeh0vMM0UWYgcf8WfESAcBHH1uFK
uHO3V0/2ecpJ+z2ouPIJeT0jqgzWUnaV1A21AYikIuNNXW9zD9QQBqTbaDKG
wX1W2xUYsJZIJHua/595ubhzSLuqocRd93X6X+aB/FUxFBtcmA9od4TqaGy0
o0yLHnhprvmWwwM9v/IFSsgkVDYMEeGmncpz9nFuC6VmQGQqUdqORg7SnxM5
Ie+fst9WjIqEgEjvjpi7sVQ2wW+Sa+iPiD/h2ShmlySeffQlhBGZ70xHQNeF
ucqnNUwK+pJ8nmFA4bTvkR0nzkf1vXVyCxRwSHaF8/6i3ijoIDQpi7GYCDcX
AruX0CYSkofhdKu3jCubU2QMyY5ZRJuoDpeBnAgIkH7yRo9Ym75FmEbaLf7N
l5ED/TjJdEiMbOdnx+GgGXEzrTMiH4tP2U3j1LddU9yq2lsS/fpVHyUZPtfY
hFLD28jWlG5pRLhR+JQZrGqUh4MVUk3aCHZY2LYJ/JF8ak5QSVcSt/fZkomb
ZQcbPFB0LWJMDPV6JCAEQPGjgrEzPfAfUBsirTfsw8FbNdQaWgSBNDCrRfvQ
GcPBVONK/iavkWRXdNXPcKqdaJRfYlOCAwkBoMCFdvQSAz3y1pJK1SX+kQCM
W3IISbyA7iUuBtymGbz2bkrqsaf/VAkh/AFq0f+D0hQpwM8tCCVyEwWm1URt
Xv8IpL5MhvRc9bHXoQJR3lNiTTbrMNSt0PVvHGB9O2d7D6j0T6oUvaqP54kb
V9kRApG+8QWlf82doAG+8D/Kpn6X7CndAGwG4fgEat8nGGTiNcImH7w9k0Cr
dji21rOwSoNSxTrlVVApJY1cvJJ//p+QQww9gzobDAT2MR4lqGOrpoXl29V8
mXPTrbDRtSYAxQEK094wnB6WR3fksPTM5ATKE4PBOtK65piVa0VGuQG1dg1x
c40ifOIep686C6Fde6YPlk01qYVjUQGGGT9Y4Fw1qWsB6Z3ZhWIf3OcwoLGC
g+JVOGLd4/m9WnQ2NEq7oaGznuUQbvAIGdSa4+5izySyTSTQiKOnpCheWYl1
InjiXH1dkOkPSbFDEXSS04bWIg01c7A0+yHVwbJpv+pgWNu+IcCIXoTEoFKg
alf/ZEQGSW0Rem5E4fj8O82u+8d1ShqaDwRI+osJMXMZGArSIlcsy9XzrbBo
kQashRI17D4PDXTaqqgIRpQDNXgW/ygkimwrv6WDnc4y/IRdjbH5vm4bI8hs
ko0KPeH3kS62/msWHXHwPibv4JxGAfhNBZDbv4sLWyrr+XlWdmPUhprC0qaY
IBiMR145Jwc6SJAa2DByHZ7Zwi/M7eckAETl0fJWhAf+B9OZwevCMx0dU+jh
IZn1o6/HkrCvytSaHkimV1+Idc1gXZcWOnZz8tywiE6Yer84eKpi0GrM7Wjx
NeRDz0Jon3Mh3hn40Pd6fFwTTisOHzeuaGixWifmiJjY5JIbet92w60+3/Zw
u84Y91Vc/QkqWc2QSko6O5cbZ2wv6Q8OZbbXIp4roJFA8TvYjD3ZuBlG3mmO
X9au71fTFy7Lfmvyz3jfZ/VsGeGfqWTjT9AKrBZTmeFA4JFoXaJS8hhmf024
1ZXSF8Wcig5WFC8owbmhSteUDjiW0y1U6EUFCKLIr79sr4JNaZquaDYCgbzn
cV6vUjiBTTHsnWdSxOIZs0ewrPsgNpAb6TszhchFT/ot1+RbFhihFzZ5GWU6
YHV1Y6Q5bdlpjeCFMO3urANJ1chMpU8IZRcmw7zCHBVpz6sfIYYWfQT+Q5Em
rZCf7acVPBLGKykJq+GuX8+RYwxbuQJ9FmEwPes5rMxj4GbsTJuXcXeNKyAR
n+cb0RTasY42LnEOu17kMus83eTT8P3DVD5U6XdIeNkc+Xoa7+HXF2Vtw27j
ZghurJoQMCko7/oFhL8ywvL3xZO9zUUeJ3xXfNggl5/Hl1AVuRRf0fj5PEr5
CeCzmta44/I4t3z8qnRmylgMfumw4HEB283c+PBe/a0X534Lgndfv5Y3nomg
3Z4u5rDubjkmaY6eQIA0LFcZtpjFAbXPvMKXvmiwaYcHBrUZ8ToDUWlCBiOm
/B3g2y9LNsHciKikR4MS+TvJYLOtwN5WEZicwaXvhByPlcXr+eV7i9b2pr38
gtxeCVhUHj92OEPuTn3YThjWUHzwgUkOMvQl+aIoi1Jx/4lfjfnuyXLrTkWq
slZMK1uhKvqv+hE/fJ2c4fkQzpQTUHCAq9DtfXKO05NDjseWSsfy6hIFHhxC
sLr+v6G93tT2smue7cPYWHfI+jHuW87pMZIHu7b2FqD1OLnIIJyFyZC9XlpV
Wvk7VRdcSPDTSqmPY1LklWicHg2GuZm2KIqVBhHLbkjxKlx1iXWRsmPsNKGA
C4cSd4+TkjUlOpombmFvUjrDmdzC/8kv2uNfvTIbZoK8LnaqKLUc6oQEicIA
cs5ay/3nKxz+qeAG8akhsXAOHHZx5jLHi3o+f1Ln43p/TPMKwKA6I+NVnQ6A
5K0INOPi1+QakQhJnv0KRy2Nl3ceQCvUZ6ix31ZZkLLHcglbGVoxcTf5EO4D
0skwXKVxKjFkDTr/dNJTy/b4QI25pUdsrIykHk/YWvw/iM3EbvpXWx9yJcNV
gis2JnBMFLLPuVlGjGo+A/Q6dQQs7Yqrxztdx8IDpjWGMWfpoIUcRd1ReLCb
8yHIembWdFVb8Z66DL3gWOop+SNmqnJv1FHQkyO5VC6jUSGrdsd9W27z5HQl
8ibwtlQEA8ByqdrUbxpCe/mun2KEMbWHpeuO8c3ms90i9yyUSCeIAssv/N6Z
3DqxbXF7RPF0kK5EA5IDkapSa9jUKfS4XLj+fbSxd2TPo5SPdV8OplOz5I7r
RDHQ9nnDzrKi82jS2JFDlhJ47M/U9632Ktn8QEawn04sNaDE5BD9oSvsbma0
3JzyRFxZTChCbayTepZ+cJVcYTM4J791HzjaMB19iOKuKs/Q81A9l0E632t6
/6CutbZ+3LvnP9hj1v8CP4vssFVPTJ/VnOK+thy3EU+pHCLtgWOzVVfrgsj3
AohUX85Nrw94AURGbCCISarg2bTTv+8WA/YidD+YZq+bIzXRQgKz7VJeF8jf
YBR6iPgiL4kPl/xL81/ak6nnK6jquVih2axAOf8PlpBORYF4KxA/SddCIaTi
274rgRN4ZUadtYvG3P5Y0uXbcX0hKno4TBr35W3YfAaQQV8UvKwD9e+P8h2d
uS4pClbp7VBA/Jd4Dvr9sg4r5EaKTn9vsnWl3cdSgY+jtSvPkKOEYfw7q6Tx
LrgC9YMVChbcUKOSrK/CIscq6zmMDwVei7dGlEatNx7/qulytXS2Z0hQh3j1
Fm66RV51wsET+8hwI3kDUOMKNylFX14AFroOfDDKPyHICTqiX4CMEnOCPW8B
9CKITaz+RWDn6VW2c2Z+kdey/Pme0EIz6G+0BSEV5Q638dPow03tosQcRso0
xKDsr0rUOVTLx6GtKuNlP3BuZWZ2AP87KizFCCmtTPeYUk/o11Ic3LcbWXvU
iQ8tJ3qCCpqS/DSot8HUHBwvqx0mYomTdQUuuIl+EsyyFAZV6Q4Av14ULMR0
RS7xriGAdR4QaVV3e3bxzhHdPzA3ProYn5YuoN9uoEZX9zrIGPhW9z8lFA6H
yZeY8Gl/ISH5pgnuqCuPDXreM1mujmd7StxghSJ9DoT3SnFogsD/oc/scfy3
bo6mqOqzDEO6hl6Lo2wEKbpqMH5iz4hQoXTnM3tsckxqM05wXfhhF+hJx+Qe
ACdU/0mSKkcn2M4PSmlfupUK7AgX5pIpwesDftgRzViQIjvwv374bxDNklr5
M5nke26EqsO9wN+Qv/8kjttOL+QYdXyP4/qqqQXx0n45B8/mvaTw1Vb7n72q
Er1xm0FgvA/fiKK4AGYQyZIS5jghuGMCYh/EXBD0VW6NWooj5L+wlhFJ1GZq
OcX6gcCI89HhEPaWKqdckTA6eb15f0IA4w1jidzfomq/7VesM4I/14y8TLFn
K9RKKB97dCtBt0IVdd+9QH2Xen0hWD7qIMM64xiVp9ilwJA0PyRTEnPHmVg+
rBgCwlWUE1jqAHnfSS1EtenXdgeT5PlNkcW4dt7i0p4dlM/j+DOQYkrFvY/9
IBHlc5pjoSdUpmMRAvshZTkVzUFVm6OEzkv+Zi+cRXMXNW401RKWgkqR+ZcK
YF1ZUoJlX8Ssjce57uUIwZse1Q8gScMwusenrAsymFAQA5UpG+VE94d5RTmF
nPZBhaqaIbOJN1W1UaMugXHxrPIMn3ohKG/2kGNoN8P21lPmLZK5B4aYjkKE
0Ygz/RoosjDNRA03cpbYsWMI0UoSHZ8V08jG7ZlbM6AgGwQpbI32QWyi8Jl1
iXcYmIjFvuKpt8JYQsRBzIJt7uI4oz2kN4SyIKfWwLzCyTT8L4kBE4NrIU3/
RvgG3Te1+UAfP33qi84vFfejRAD9An4rnU+Lv8bHk/GCIEtvAxEVClrzpJY1
JmzvITCx8jC7S67wenoWJ2/vkgAOzqBOoBMd6aP84pGv+hXxqksj59bQuMVY
dMnBqcBuBHvWKsjqh8AxqtoI4xb9Pa429Jzn9tRAIAIEj+iXlfIch/6eK/20
o91PuPnf+VXhBAUbiL5dosgybVEV9Uk4EzfVpbWtT+j8hUl6ZLgreUsAqr+U
kAfkhGQ+OdpXYVKSSFXjv98UglN4Lhgdldr+aIboonwe/H/Thj2+W2j5kpV7
LnWuyy10eydZ4hMuJIdWvPFgj0NP/JhXhZjgFvrKEy19Cgwdb4cGieO+8Oq9
O2C02d/nXZhsD/kKB25G1UVBU9JBckfUv5EzCqG9zben7/5a4QPCyJsmLbWn
oPI6LWkKdjSlsO9gzllft8Qt7q5Si9jaRa8hs92TOmPn6Ppo0k9c+LrsFXSm
10CDUZ1Bw0ePyUD6798j7bf/KNLgA1+q5Mp1huhCNS1jpTfHKuVmcrIRVeik
eeMGiqpdBIAVcGtugqbfL4o5ERglPkz/i/i/r1a7ifIKep9OY/95YQ1S7q2X
sER6y6JM8wZs9gIFVKfD5IetXS+r/PM6Rw9lHb/TZjaX/CLNe/w7Jl6QXrAy
axIH+45h24SLN+LfXB6XIXEPsX5Xxui5yBSB0USpniycIEqLx56DILvGmK/1
XmsnogXHVU1o5h5ETyThr6xMwrA9PJy6InpbBotrd4W3wpdEgso8Y97yDpKA
fS+sNlNzkMusDDhBHydHXjkND2YlMq1tK3K6pgkvNIbIcJWkMCQIMt95kEF+
zfazoKI5eBEPJIt1YE/Y1u5BKoWUkn5+uVwnv8iivrXzR6BxN0Dau85uQEMm
PH+YaR6NxYksfGVn4cGZphEL/h8BGsp4lOq9HcUadkJOZ6VUvVCrMgn4C4lM
9vKo4hwF6L2AwdeJ/3ZGV5mvQL31IsFxkcgpBTvbSLMRaXj0lF5n1wE6QkLD
TT5d8S1JuqSfylY1SyWitNjtMebtraAG3JSAn/C7ncsyGEl65QyuJSbPs+pF
IJMK45TFwKtqyX1w+w1irtGRG+sAVQ28miuv4QyUQ0jqi8RXpIWE7A43R/mb
HZatkgUzuKtn7vpeiIo8Ys/flEQB//3nBuvTaI9oSVS16Xui/AqAilkq08xM
Doo+cl3sp9pil6NQcomTld4aciecj+ZlnQg0rAM/9V5g10yNJUntdt7XbuRn
5H9pTNcvlXH6g5UhKi8pUYjz/YHxzdfhef1McW1C1qeFsmJxE06/Z7KrWCnl
nKuiF+IdBGdMPkUX8Qhn1lTxX3Ks5tvjrwSSe/3ZhJi69KWOKkb08jtTbtk6
3U7MZtsm2fxA1nmHdrRbHUhuL+6o3udDpY7g/3i+93Twx6NJ3+Tmyxs4/rb0
dc2G55fVbJ6pwWUcYYo4KNkczY3ts9KrNgnqVfnokO7FdR0lzotohOa2j3CI
csobLI8JA260JvLHk/g/WwYBH3uPolCgWQ2vtO780MLBKMBDpqVsDh8me0i+
0zi5IkKD5EkxXo/3TOHgOyuh/jMMSRSEp4DU7lg74nwq3xx/HFfL36bnIr2H
rvE6RhRzzUOp5yRVeLGSCM+biIvlLL5cOn37H/BQCIfFA27QXFbwibkGWJef
MBBuuIX0KQrS2k6E4hvrttcGbZN3QexigtIhhMtRbv0LW/Ul1TQ8IbOKC+tm
0f3cw53aqgDRGTXNlWzSTM7Br7RduBmBJO5aR6EAIWPMpNG4DNjw9+8cxBZO
vJahgl+9deOnh03OSkLmr3bOX3Pkm9ehJRQtLVx8MkB/yE0HMpyU6qLXXDy8
MRZWBM8A8tFRroA4GNMvrm0YApNDdvf1DGV4Jnvn/qNdwhcDsQmlQjbauLcw
04SHY9bMQN/T3TPPGezQvYBlyMBae1+dGRuG2WtTUhgIchUFu75nHm3qd1LB
hIft+3ienK4mF118qhRdSLRllLym3t6DmVdcBKy2KqB/6KcZmGoLdw8B6QCT
MjwOmba0Ucr1S09PV4qudWBiSO7TRjF0TjFMhT77TKmrxbXY74mqA6jKQldE
cQ8k07LissNihoDLpVUVm0KLid2aZv6n2aHCBRw0r8FHA7t4tKCmoqFtuvDQ
tBJLXzzXZsFzYyHdK7mP/22GKjVz12KKsNGGItl4yCRiLUJhXdsaEf62tsny
3F3sWIM/BTjXkrayuQiP6go1Hxc4Ux2PIFJeGzsEKWo6dVk/IBLop+OI+Uw6
CVJFBkkv/432Ee4tPSLVyHfDSQfBB6gg9zgZu+ZZIEmHJHkSIZVnWfpPoZnh
BDKuiQrzafdIXDWeQDZlTRCmhXuYOgMaM//omZerQHxmsX3xhOq7OtnYi9ym
pXeUFbvUlUYlxkvdlFHMggmfVVuE0MVsBiWj3PNc0768+4d9wCDGSWHKXx5i
ETvrcfxt2Q2JlQdp8tkdQzxIip+JANnUNVRI8BEvpHfcr2VuDVa+Z6ktoJ+V
iirUdxQGF48oaidK5NS3k7nGyYIZ2vXmw3qlUnOv37LWtJ/ahcz4o1fA3kaH
fp5ylwSsQzr2e5OupG9QBkrcWpKE2Lmrc86H3V4QlnYXVgLK9xeYMu4JJ86i
EM6Bq5LZZoqNQlEgtt/y6ZujthwVUXCY+WVnWfgsZH534djJs6W3/jJAdiXQ
oMIzHocsJ4laGFIbKIkt3jDz6wvbRPcPOoGkxNNu2Rl0OdcOD2u635fb0AUe
gU4uEN8goy37xt9OZMwUTBNIW5yPKf76q8PHTSiV9SVTzPMm7g+aS+hJDIT6
4WkyVqf4h5Rl7ydzQanwTyfTR4gyZLX6AdwFRk900lCkShlmdvmndyJ0c6p4
j4wdkgllL6zKoav6Xd1dpFtwPXGL6hNuBNRZLM1iTswbdeXV9b74SYyiu4ND
IYc1N2twgZKwS6HzKZor/a6Vb96LPpDgNQDQUj8KpUpjuG7P/QtPVrWwHeo1
iI5YbL1nsGXABF16JsRppYwgpuEb4RHSv/5BcX1hsJOvDGuqwKr4zyprtGqK
fhrw9QT01edhuOA3foWnGzMWOPL/7vOp52R9fs3RXlGaoFKJKORZpKEYdFYU
8sgsM3seJhfQ/eRrT0v7/qLcBAxKWirRw/AMFWJ9fi/Z+CvtCCgHLR0t8DXV
X1CSCYKxhkPKZ80nIP+uu2mNaQn8iIfmaQXNVepf9JcD8kiBsop30lQoaUeK
sBWn3rUSHw4o42yoYT+aGLIBOfWPBzT3UstohTJHypUhuSRZeHM3+ZmGnS8z
xmzVELxFQJvfxUy6YhF1FhsKhWUSXTnCxUfwrEqgwabGBjqIs4a4PI3lkF3N
qa+2syxZPwmjHMTqYI0bqwy8VK2lBjZoh+uLpX6uNI0MNLwyXcz0n+pLCDbF
T9jFGPqN3IidiKAYFr/WZmlaIn2Y5b+geSyM/1PyyuQAZmspcoduETCNFIY9
wFYshAtyhXSaiaEV268q1SyHmWvA/YkwddspJ/KHsUPAM71DWctDO7Dtqupi
bC53xcr/ESX7L7j4gVGsnF102SFHQL8FigM3G1FkKI951PROpE6RYXHlhKaj
nnxGyvfnX1H/qmCqP9C4VDCLWzS68jKBd4ZjJwwIfKH9Q7OALz5UD43bQJe5
OmHbzxwYBXkfS4+TtukTpoM1gA/cAMlZqeUg4hRWbsMOKwGD8pLQl4xdBUr8
J3TQb2PDaW1tNTQqSgHZKS5zkQQkKUBAI/PX/kx5aks7taKUckZlH2tbbaE2
yxqje8pat2ROCCjApjreMAqOH3pl/M7lEvlZBm+HwlZf8pjcbw9CS9HkrdnX
GOJ68cvwTYz1MRaNZV6ge7m9RztsCsAxNdp0QHHSiBVM4tBdKvMI6vBPfbRD
boXEGUCbn0pDoZRmyVcuBL0BstMLg8spuGKrgmE9aQw+xCvnAl/cboiaupNy
jGt8kS+cIQr73PivGbTGxc2sN5dJgXIYFEFRYAV4wJlhhAY3TIF2Y/CG2kOn
FZrsdiOGSPHXCRSPqAzgBrDnLynmKce+HODXMwsIC8ro894+YB4L3UQnhHu7
MXhmVcJxQb98PuWESPRBgsN7A+WZL8AledEfti63VGrom7NQx8wQg3wAAVqe
nrfxQzgiNQOODvQiWLmLCF4J0IGxHCgJDWE+UN8ABLAgno7yfo7KW6v3Nt9n
Vu9nhctqR5iPGH8IyjXcqt+kY0pMWBD0kD0OB1GuLBiUHA9o44xGZQB/LYw2
+mLpgp5Lv0tp7FBebbHuTOnXSXkHMT9KfzVImS4At0wk9P7GZh8V6XejLzrR
nserLNRasD94DQCygUu2z89P/gi+1CBqW9dKfmtQvACtbJJV6wZTNChb01yS
+FGQYZYIdAS1zrxY8VuGPbWlxzKfYNXtX7AufFJNpFzRnOybiyL2WneRO0MI
8t32LED5LvRTJCkFx9F1oiBFbCNSrg6rg7ggwZDsO2xpaGuybmaiJfwX1o7+
t2J6JrfTrxzH5RbL31SvbsC/1cC0IL0PweamVvHzg2X2/kWQNcdA1ersEK3u
1p/L0qEjdAY/TCCTFOX6b2s3B4MT+lkXvUk3zkRTo1QkC+hcnq9+V/By5LZA
z97PZpWwNWRjJ0QwjCJ7anB69mKVis/n0uRtSlLDBEGFPpNYKFaR3mOgomUf
FsnOCYg+GchOTfiIEjafjQj8hXtiPXqVPL7U6rN6h2lQYkUw5dxxnyxi1svq
t2HERgCXGMJZFcDMF7hxyhPVOJ8y2fWmjBIuaVYQFH7wPyu0Psa2lTGIro+a
SzzkpawpUUwC8g5TTTcVloETAwlLJDK1RIpHM6D26oA/7wjRSAvOMijqk6m/
qRlP8BHraAPJfXw6vhzAPVRpnRniI8uynEk2LdD8zWKAayDefq7XO/y7toRq
0y+krG8MRWacKYavIeWiKlVSQWxhVTDXSLIu5XutsrTOrqROQbwKlkvUKjmm
KpuZdYQGW31zIeaPVDaeVtSycL3MXvbf+ve2kGb25eJhWxlUa0t8/qzzBKvi
FvNTVCgox775UdkyRkktIOCwBLK4QDPqakzlD+0uQ9B4W5d1UvzufNNligNp
PClAZNEUSLor/knjUPzVO+da1OlFuLLyGku9kAJneW3Pjq9YERwCexokDLcU
o8O5GR9kVqeLjPj8mQMVbAiNUg+qOVeM2WkdrfFEiUh5ASgFUHvbql8hKSj+
VY/BdiNKBdh0yDIhkesFt4vHZjjA3YmYFMPs4mqQ/2kTVGOGhtmaBjNgQXTo
3ekF7/eMe92hSXbX9blEboSmiFH4smNYRFCgsSEqlMTjXM4jJmf7rNAZDfcH
0MFe3gu2jPktRqrv35usRRmQH+nV0M/AkWvFk2xfUqW1ioOFsCpjwUV0+1+y
hQFOsNZ1YmIDlrQsS4nrkh4NL0VpD+w4OUzwBe2ytITTE8hjYtEc5uTtiTVa
lC4aSw68SV7pcQnuHMsyBbH2sKjshyY/US12TYmpl+PuCn8k1j98k4TrVnHy
vYY6px8BOzoxmJsGlgskggq8e2mRVgTV33eBxl/RXSyotZzwrki0MoQuUEy7
A7lA4TV4ZGGMYMcrVJVb1+9LKl/IouZQZfUELmXDMCiigHUusjO5/vZylctP
ruVPiSKWzLLbR4F8nZ6oFYBvYYb0WGqnTq3UWiaF0uo30i4VeGu/ABupefaN
DfseIt6B1JavkYOZOL02fhSo7MahvbG+AKDIcaCl+Q3Q4O9jVeC+KYRuwUV/
VC3Xpi1XadR+pq+gdUP7tS4r+6yr6KFqqiNLFoP7v26TcC6Hb+4xD9DBeeaz
MFTzJVR5LF+lGPKb4sRMUwCEvvjPk/yNjVDBLtGkcE2W5QdOlFnJByKnSaKF
EnR+aWfWSw2+1Vhp4+TA8xAyz6aPuaZbMMIv+HINZPf4xaIGZs0jcHKJGAc0
xLt3Zt711IYgJZpT8U10m8EwJ19Z4y/YaJ4ij+D7f2ygDGla9+L4KTYreSYN
3rdWEmta6I6gsf/qVnQPFPmzHVaN/8cptIbOMHTqJiO2kekgaczomqdziycZ
A7Ezh7caqkds7E6XFN0oS37EdVt0NLe1NbxbOIiyHjb1JK+che2E5Hk6q0gw
PGxJpb9Zf8yAR/OxRNrUa1bm6v5JPojlA/2l/JbuxmbwIZpNB3O+JkW2hYXF
qQelKF0+y+pA9dzQQXOnO9TuudE8wqZ4zLMYYgSIOXYdLIdqylJHK/V+DXwe
8R3skBgLfhP33enxVGfJQ1+0pvirNhJsuAlQ01rPLpxbKW5CuOIP7hnezkAo
FVWNRC2B3vfZpSEBrmBHcZwcE32MEsOkHjS4Ic+WaIX1VsMG+UJssZJyACz8
wQFlxi1zju6ULsgVWG8dzgTPPZSZ28MoFPcpQ0RiLmL/8LsUM7YUDcQ252kF
wcq1aYSB//3a/wkuA3LDNTAD0As0SqNyw6Ouj/5wTERM3hyvQUP5znwZ902J
aUe5T0+k5mb85w2JliE3O9xnOYXVbtOVumF+y7wlS60tzI81QiylGxrApI1U
n/JdxGkz91fO1fSHNpL9lHX9uBSDOWbt54Hd9N2QLPTCGo7WDMrUeLXmmn6g
SWPbNgyS/atUQwGZ00qiilcdfEooRuKV/Fr6zZ5S/RKuVUSJNref+nwLRmsJ
UVB8BKLDa+eyVJnVtft7UX8z5kFkj4+CKpOUy6eCcZChLsFO1xK2y90WwzZb
+Y+y/XREtGgr3YdQupEsEcO869ScZsaz74L8vyT6AqDy/q/xoo0BK9Cvy8aj
12/6CSDHt7LeLBGNg5/xHFkH1jejWhKLSyYJtFmTK/J9w8UlCicRWZtK5//J
8rOoT5b7v9WoObcveEWNBXdb4JnaiBpWNdMLIQdPLf6nt1SFgyb4pXTkoC7I
ss9mviR1GFtBSANsiAg+mXOEMbSGCgtH0oNg8Tf83Yh62HK0zeUMCEPxNJCi
iUhy2BioU9GQi0bxgMX0c8xe4TmQv54NsxBDaY1ZfzHBhxPPL7tL4zg+lpXc
BWJ4V2MHrJU4mN51IZR/Hr92Tgu/c7HsWeIJI6qD+UvLdBu3VIxFCpchvnCX
xtowtYvrg3CuV5IAE73+kWrxhYfcMv0oHpWWV0OIZZ0S9S6mGpEDKoUMR8FU
czU7sgzzuSRAGvk1VTcaGmZJyqeUvXDWUlLUXZ7tLIaSLwS683cIIOEKfJmR
Qfo8zNMdrSXuvra1V6SGo2/xOMcCwGulnkQzJnlMNOJcHIqekpkGxM1exQ2g
2hDH4Cqjg9eX+/JBZp/JP1Qh8Panm87C3T/PcFh8jxHFuIkBuy9gTHRUSBzL
tqk7gcy5O8+Tepkdj4xfWkmRijWve9OWzc+Rd9/k58GZXtXD79oawoXjqg7D
0aib+viCiZ0exnBDM4xxYrJUlDW8gY1B+b5jkB2C4h2rBcRH1th1Tj8MGS8T
OvTunKI2V4JcdXhelUg4FP8dBz/hhFVwxFJeD1YDtW8Dv6Z1OruheSpqInzE
SNdDeWcduAk9YzTCFmI+gBivEVsS0K5tEWTll8VVWTq3Yuypz0e9RO7zsTCp
F32SVixSU/X9pMhpazoY2FcEPtt9OSCyDpNUqGO0UQMCqJlLtluCRfbXN8fw
MRkLCJ8O4KdiKe60NoO3rWfXa5OJtFtyvcnevVHAkNdB24EZjYWfQIjHgFjt
sXSH5qMer4ij2I0pB3aXnwD0OZHpn7lMzyattTm6Lwh2znzqFRzySfc6atDG
a39/V0v597QmEteSGLs+N3vR3YB/+UMZHQl0/d8dgfIr39LhdoHMCmT6r90/
jV5XlKVUAh4iPulXSW7tKlNzca5ysphQIsgxxkMoJPhNdm4kr8seiZ/DJ5WR
Kq7KnHNrAMbbPbvYw8ECZCkUtr6zUXXpeZHf9mNv61RbJZHQZ9EY/s6pzrGN
XPnEc0NkEpEEA49WCHhFtQzxIpsmqNi/3H9wtgrRYCuwZ46UcYgus8t5roya
g6T7nWEzgoQxLT4FU/rARYBCk4+95J0V0mxX/Xkrreb5n3sy9MGVq4Hfgm0x
MKjpRC7SJdKcPjMj5pvtykQMRQyrhx4DFr/bNxZS51mbejZjvfSYNS1vXyfj
K0YpTxLwhukLfrUfzmQNh+SGHO0PdCYF1ay56hsp/Vqb0sBJAOdF3qQehwpP
yNlyaZ0zoo5SYLYjp/5UquwO/nx5K7J1qjYlRLsVTy7YzkW5A4E2mvKhLpJz
wR9aLOAko/3lUpjsSccaSsu7P11tQ3kGYPbARGsPG7RXzDvu8CL9NfzWtfhC
fSIcwmuK4BCe9THroH6puFULGI/pUGrpQfJBw9/Rcp9YoJbjh6pY4O/AJPd/
KMCIeXblgQ+nhuf8qdKM5HnHv9gdWJ2UhjuVVWKiwWhdEtTjMZ9oxOGjujCK
2+nnlYHK8Teca+dGk68/SxIUIad53yas7ccYuxdbG8TFaQI6dy273FrEwkgW
ZKdWQbN41d0anBLslI35rMeqQcmymQsnzTBt7/2zISCuLgKVJHgomUBYid3/
HhCmH/gjYdGUfEz3TdbB1FZML5CxrG86Bsm8niidA4e9EbvszvH8rnFZLcTC
eB7u0KAw/8HT4AHXJXTNO09VTxC1JYYlacDdc4qL2cZfsUj7hky3czku7bi8
fn+6cxqZmIJOrG+qsZ8GXuR4NnFt3Uk4dN2SAYPl+nPjjQwLFc9EFWsBZoq3
qUjEnOdUjtPUkrvorNuaib80e//IAo+sEcYLwfSjXqwTS62/acztQeTLhT3B
KGA8aBmfjQh+iEvzmYRPVl3fbIPd9mH2WGjWN7cGiu9gcTvgCGzJhyiLasS5
ZxcGwpg/xxPFVIDukw+fssCBDnwYo3S8aD1JKuwn+b/AbFmfJfuX+GNiiF9Q
krPE3aP/Fz/UrHCMObi2689EPaXeUXAQk4YXBsCjnNvedM6bEiRAJIpTd//e
3V2gMuLhtugvtWttOufV6HiQWmfZPkmHyXOQSamVVIHgzkDDqtAx+IQX92XM
Zu78P437ALdtN2R/Wkcr1AM7KXKNZ6Rie1SBXzJ2a0aEYuXf3FFt5Y+pSmsl
RiNq0sjj1S+KJOwHOBqNsevaC0y5iOj5JP+oq/GTEaHsXD7yKsDjT8scKzr2
VoElPDe873iWHDz9nN4lbuCan/nuaBpYBZM/B2uYKV5imcevt9X1uB3vsG0R
FBMTGE2oAPKkC20lruocdu/f79rztZykEYBme9PqlbGzcD99M4XtCPXLZPEg
xiALvImiGwvke7GvQWPPIo0UPC2351odpgmqhgVq7bKTOylMeqLYUwTvVU3q
uA2b1ZUwkzSZNCSQ+DBwYDvDoJKLCBx2YlzKsAByJ8/5aci8941ygWJQzTbo
c+rjs1+a2yU7X8ZjLQgSoezsQDgRFTB7udcCOt2NTT2myKxcN22kLPjnJk4K
xfITxBEMuy9wJ6QFO8yq8fK063XHxsNX7+oDf2MxUkDeFQvHnIlhzFKooLXK
GfYSK6n+vtuvC9iKZsnVG607KOy/6CE17tT9MDPvT6bs79D/eW0/oSeh2JU5
GLuiwKdNbfAuBPQMEhzFihc7T2CLatuRspe6ETuRJwZ0PJF8/U1rcyfJK0wR
Kkn1FJrGHd6TXMQkU6u6dW38HfCkFlhmO6Htj1kkVXZqPLpUqJvJkeGwwZoV
VFdU9db/M/06g9U3CGgKBpH06WUryVDwZBwg/wKBVAROoXIvNoniFW0OtfLh
V3WRMc/70SF4Gmx+LyWX+NyUEoxeCmHv+p45d9j4vjlbzjZ51odgLtEF2irW
0y3Nvw+u70l7jfNoeRfcGHF27ch95B+XXjQ1BJbbDQZmZjIVkeoSo8R46u7t
aRlVl0K3Myt78C09KSA71AeNgRNj2Cj7TH9s031Tm4cqH/8+DRO5eWne6Fw6
atdzlMscmNQmeUs431XBUKNAa7U1x6PB4tKpDAyWSWVyCs/NvQ2fCT0tt7X4
lZb+pMRLdvx3XHSGj0iu0DdH4YR2DcuenHNPgN2wWMV9IfnQSBOm5zOOO7wy
6WNO8cHe2X05GuodWzFH/vMdofsIvF2GVdD42pMXNJiJpimZL2k01ywfNTi+
bbO4zZ4qm4WAjv9JSwPUEM4c546JF4w46pL2SWtg4zp65ESYRzv7QuoWgVZk
19qbwgesswmCqYVUalVPIg5JVfiETyLqa5GRDUldHDYVPCVqzyAf0qD5fTeQ
VUGV4IUU2peV+YG2Y1hYqu8wm9PVASlKowsZRkKLub7Il6oRcf4PI+TWJABH
9toOJHZF7NoWPXNscM9MjiKm5nvAfQDeacjAgSSZJYgmEIn5zOdzBsnv0k9a
QtgcjMzHZkk/fQ3pMksQeAi9MduKUOZoAkDiQlMPPMwba6jom4/BXzMlDpZ+
Zp3gSXvczMt+ke8YjV2KJK/AcVH23Z9j8RFKbZUT56KyXHizQrswr3Z6xWSZ
4XzpofTxKCALtqCPKPAdGdg9++mNkrneSsm9itpmH1ZWm1sZvLNUKUcofUUL
83sw25UWpBWrTqMkUHp0bbREycucmn8ZrAO9g1XjtPjgh+g+PKqJV8JtIK2m
w47twx0ZCZLbz1/GyLTg4VWZ5eZoLCID+BFynpI/7p2TRp5KDjyzT+CPC4DM
1aYYnLxt1Q2K8zszyTUvBodFYSd+g+87syKhpQ8M9Rg3gVF0Wns7xd+PeBfA
H/hmHTok3PfLzn8ll9skzUwwncp4JHrFE6CUBrdHO5Z63WkOSbsKJe9tqus5
gyQsFMDYD9MOIIZJcUYlM9uWu7iYn9sSePeLPWCG1NzHnGdDoF6CACTlIA65
a6DP1d7FaLBsvpcTjxlp8z7lVYZkKa7ANqR6VWg0WPLS6MnLMucWa3yXmXBf
m4dW+7AKqihOFDAZ7y9FKmZ7JPMTeedF4FETOcHExFQD+lCfyle8M8B8ns0w
KcqDfqSs68/XCcP8YOVljkKEzujsMqtb3UpKBZUC7cP2ENjKOPbQhKbVFuP9
g3G43j0W33WuodVheGW0DjW4GecivCJCEphIsYwK8oV+uZhWMVngo1G5DdRd
6/Oe1i8ZJ9jpyp2rbZOLT0BlpED0TedGsK10QrdSBV/XoJaBR9sCAFtWGWVB
If/PI0tvF4vj0v8HsNWswLEtEw0hum/4mPyr7SgAiq3aKbqNJ3n5TfiiyLMg
ykMuBnWmpVqnAzAhm/0J69GK3TEgbli40NJPXLq5jZjN1eJlyhfLaHrzVlq5
kW3tpzDaL2LEL/Vb82r1rAhwCZGWmg2w0M34scmUHjI8f9lGx8JHrl5qmIon
LOK9oJsWs5npVMGB+dlUQQByVzanjL2YX2crH8rMkdenrJ3di5Q/HgW2bf38
apIzvNMPZTZWXb+Y8+VhVmUvz0rfrimKDEKJLgL6R+WsJTAgr6sp/5wUZB92
rnsCsJELBJ25d/TUXmkpx//yU12VofCZdN6yH7mdhjT1LP0BPxYoDd06T/Zm
Vbnm2TwrDJVc20UyDH2NcyQ4tJ5J20ATJcPwWqM2jYFc3bkaQH73WoWjBPOE
19vPUdZyIIa0jrKI422LId2GmisCVM34xbtgwRNifhm4WHi/Y+Vp/A0BtGmT
gvcu7EfATzqXTug9lg154FRftHRsPKmcGcgXCD7m+Ltkze2k5w2Rtx9U+RIB
zYmSpxSkmvWgfhFKRpKOhv7IVQV1KNwZZNwwV/xDAC4cPuryFB236oSToISe
QNPTHrdH0T8qwb77m9iYCnf4LlPuBOYccgwSwduEzNGDIZnyvnkNvzPQ4wtw
jYt/6XRMQfUwRvbaSh1TGVNgbelkyDJ4P5lqFgyAOvyNiMJXveKHUON2ngMO
xvyaUReLfby92ZImxaCUhxFS0Im+LEu1Ds88ytZqGbPiVgKSUOGBYgSfLMHC
5Hb/5UtJVUgeASwQGArgQTNZgbIDzOfjTesksYNlmueDDtPBlZ49Mgyvt61Z
IpiP97p46DW2FSQR6Uh5k0cKbqLSlK4ETSOY4UVwXP0d+4eFoQESNFOL+Wtd
dSDefSV+qHwC8pAIEwt27r8+9Cx8uVoyZgBr1Don9br7D4HG65jznRBB70Hg
NfoKLwo0++lFR7grgCauiKLZ5uX4eaXbm+oVhsq0QDV5unHog+9kzrWj8Kmz
vshB1JXVyGKe20SEohBMSvkAfj43nUxJEHClT/s5U7THHB+JdcAVs6puYoGT
8CTeIRucOKlDEx9YZQjSj4fZmNf4xU1TVunmEbkKuKBd/NFTHtNwu7OGbWI3
lcRzg63oJ7DzO0dbpGQ9v5dSb85eAqhabmH653xSCEQkCkxrt0odIBoDmexA
6kgCiu2jtz18ERDj6B8S9+fe9ZeIdU5GBVA4XeWNyocyqwUz3UXVGg4kIrC5
mPn32Ricuh7fVclG5MmAYhZ0Gz7TQGQA+nW6dQBzGBtXGCA3qrwt+l6Jxqnh
pENJq467jPWndVcZyEtgbI39mRVd5aR88y12BXg4ztVSasl37wIxipP66f/J
713Kmlcwo6PFoWwIemtgDCqSSmkOXSCVb/yO3mlAMSpDxr+Ab4ewgMbXHvAL
TyoVBvmlJCNBqQc/v1zm7qo9qf6/BWzKbRwea7c4o1j26JhnCJpWDUM4njpx
fyy8fF2750NLgmXnaCB4S7NeISzmVdce/P8WpzbivdeW+geNE3bYw33+toHz
mrWIP8vAF6wyFEYQgY+eGm1a/pHN1CXTsB3oTdg2W81AkBK6mmiix8SZ5K5s
RMxTePHDlGnrRHpWgMl2vHwZKRINRD7e6f5Wn9PiH1RHitX8D38lZ7hOPkDA
YRG4AepL3IdGaG68Hm3KPrRJXa7Q3yjmVYfsxTEvGHKrCdnrmrx/mMiWshsx
QPi+7XUM55jO5v0IjjPcouoRmTXbZbJADTkdS6A1y9wT1Qzgftu+CXJODpl2
m7jDzfkJ7wKJbnTybcjAoJyw6qwOEq+hY90QShLMS44V1W8uAMubVFQhJOHN
VoMu2VXJQdSVa/2PGDggKf6umTKYF1LGJvIxuhqwF42Xti4f/R0504vNc3vv
AZgAqOFGczcArYifm6EG8/1chgxVkBpDiQ+BwY+ldc1aIlfcylLMiips0xE9
UTFC0wzDu7x95yV4QKXAkje/OwnSmcwgaZKGBR6toOkTHSclIY1FpsTm06C5
Dbp7SuEGAIsDChXrJuvVIJlM/mrVhc52P2rP4rFzDyTDXHhOzLfJCYOWA985
NJ1hekx08enAToko17IizSVbHa2o51Y8dQ++9cMHZ3hsfIzCtYl+OkMTTB98
SwQZkAdGZKIeKOGc3DZSgdaBnpuBYlxpURR/pVMEr5miZOmWKiledm7ZhM9L
bEV9hDhmELtXJXcx594soYptTZybrcGJSgrbEu0orM+e0fWtqWn/jPmj3SP4
Hv2UUf3K9VAIxRNKJHW3q14sXWW5IRglV0K1KmTcu5svZ/3mm/+MZM75o/kv
L4icwcrckFMGJJZ24Lpip8HaNH4NjWn/M9xBjFtGUfYgs4U0ynG+wSk8S/wi
2iuu7fj115wGC8XfWpztzZkYFbOjyYpf1Pc9lrI3kOB1tFq4YBo11zDrkKnW
x4ufsQMxnvN/XXh7vrCtq5U2z2nYzdyRzpVrbKKBSVkXVH0vpExd/a4CYcRN
1FpV8t7fVoy0YmbSNcVg8sxuWIWWSHjPVdPyGJLsbP2UNJCqGhM3X2fqIX6H
d7J87yY/MinHqy53ZvVLcpOb9Tz7Zvoxf0WdoByGV38L8QnylDvgRQeg71Lj
MlJjJUlCFyL2cKtyYSTe7nL8YI+qLY301loN6YhvDD3CS24P7Sgnm/oRGKtq
nUQNqbstIZDqAv6IyTo6jhuH+KeRppRumJtvb7+oOmxS4fnQ+gQvYHICi3qY
VVvGpJb7mDvagsZ9C0VUeiia8XJdxUrZVK0CTAaNBuGmuPdlbtntz80QtoNZ
V7YFXtRx1aD9g+B5pBCZUkdr/UkNBn67pAFu+xET30JKua9jA0OJAgdsHSvM
8lRZ19de10e5ERxGbPaUZaAA04Wvwuanwj21Q6eMDakhO7gfCoL2Pe5stPZd
RWcgqamV3ItzZCGjhPrWUtrvI04JIJ6oQztkEQGrMQ5Huly9toTm3fZIV0iB
ZLJ1FT5MDNHLCqX2CzwF+Qt51NVdPWUhLpCdV3YvKMMhhlttvz3K9ktI7o/y
n4pf8n+Fkvo4Zi+rnPxM/5EtyMAGQzdgsPbAA2NC76+xHRVlu97X+C3Qc37A
7/he7OMFcW3Qh+ouQjoGYjs+WCKhXw6RtyRv3axTlIvmsTBPs+NJ9/Rz5XXw
fjLWXooIfSu5uex856ZsCM/Kw9+HREa8quQcq8Fn1STRHm1cUYTbKphnm5qo
mZS1XPT+ZIVD9bfffJRS4LnwREUv/IBd5KlsT34Wyl4mXbv+Stn15RxUB+2/
VjCIVZaa3T0H8wWZlImbU23C6zzFenDJfSV/RaOWnZN4KvASfrU4CoY3vgMn
Igzen1cgmiIvGFyzkCzi6C+W7MKb2m/HIJGsfU3EgFd3XliWc8OlMFac2AK6
ijjt5D72M5iesQf/kkcp8EqmPeHVAezn7d8Oq41cs+dkYsDKJJMTGDkAgyoA
R4gO4MNjRKroLzByV+Bg3K1DT/IO2extLdGOIoik7z8leiwt24Syi9pbusu9
tA/CdkcWboF5/5ChhGVB5fzbSk408dgJcoEK8xUc2vsgQLMLzcziBI+y2ik1
Il0IBtHrLD2KvLpudWdpkkR7tIH7F0y4uHkWOFJ4wwDtM35/izaY4p1gjIm6
mWW8U4ic2bLuzj6AEWMd4laXmvl0PKa9DyDZva4IUazvSKOK8saOhxmC3h4w
pyLCNUnFLwnQwyn/3bsYxwxWqk2fhIyqXRAoKAbChaOHb9RGE2SNuFWMz4pv
EUHPYVEMbPfQ7IU1j994tmfUp5X2wBYg6CjQFkW91pqWRkv0ANnmt0zdKOgp
VtvBEAz1nqF/fbfNYQoPLDYNm4DfaM9r7TIrkd3Cw9ZV0ioqYdLDeD/PHRVr
iuZQ5GrSxfeujBHM2daIj2FDNTU6PoFc8MJFkqRiPo2JY9fmPKAlu8vPTlSY
q7ewzFkrkuhsPzWMWiWN+LUwZWdg20XlO5oGnAFavcoN99tGc38EVzQwkT3n
KcJTi0se0YXehz+XXMX2gKkWIOSQcnK9izCWSuOAO7hpM9xgGBBItLWeXfBq
tkDKMoxtD8p/sC802EUbsdaRl7aMG1PXPfcAcQWrGYLLjpdzMO53iL8OASF3
tnsZfpw/xSDmls/vjmnEbHQ7fZo7oNnnvqoGoqmOtduUusYq9kZ0Mk5G8esQ
T+3XyMTDctV81+/Z6HziAyetnT2iWyHKsNQLVKi/fJeHlALjTiqEhAYUyEFC
X+thVquxpsMfDNL0I+g187Uf4vK59j4UlM+II87oOKq5CmIhry/5jCKZvGeZ
O89Bq+L5whesnyMAQDjjpwrQ0NhBdbBSXvpFoKilfHUZtydiSGi4qsZpsSgE
TqpgvRKcPv10nIG2BzOMcy6KEYDhTe9MPj6WlRNcszEeuWr+INiV0Pkv8Dwr
kb2cw4YjHOs7Umf1m7I/COVh9QrLfKW7S8mL1E6zsNXMy5ZyZtSEVYBb1ciE
y4nEgxbS9bslI90iJO+fVo8BWGkSrTr3TQHOSPrhORhiufgVQUCvKcqHoMuH
536CPtxd/0lIH7Ol1zfnWA3/E7WdoJxbWEUjlI2J6nah4V637/RMU0k1zL+L
si/FOVZ56l4vGOCUiVD4oZt7p5pOg5fH1crnNLGpc+js/RAPehUnm8FErAHG
gp0C1VBt1MJC9DKxwMAdxL0R0MRFWGLTt43keJlE5/FgTmzeqlSpeLkAeG7q
3T7MfeDOtH6kKpugQTBl8H3qczOBEacnUMELodh705LVkMH6ojyDBKXBKn+L
G85LZ+L6iQ6No2BJILsD+lknAUsvFPQXDYjDxyjnl/VQMSI/z4zZgCuy2DKF
yjWochdoO8zK7NaYyDyBedkyLVddwyCzzp1lTpreD1mROqgRXmaPVSHDxbLY
YIU2nFC8AyMq6E7AkdNQJSamMzauQSlfHp1URWHrg7thza0dUqbiTZCZ8yOd
O9EUgCl4RhBLQdjblLbIN/UdUOQ/lUYDrkNzbauAwB0eek3e8Yohdz6CUq4R
b+/eorqyqOn4fxWFPJBrJ7KP2sCMnqKTFIudWL4+j4KCMf/JnAFNIZjs0xuD
grEnvYFmwmsJ/4nDfdeTsKCkp20Ds3ePRh4wso/FovTXpsYzWUiXe954P7Uu
0G32i3FU3YonlshwWTWLet3NvZwiA4pSYiKPIbNGZTv/ATrKsXjU2t79CFed
RkSi9Yuc/nYuXHqvPz0/g+b90motuWMkeLqkGuH2AvYOJuswkmR5OwrbCdzL
HQ/z3gTafW98nF7oveKoaN8aTC3gY/UBj0ijei24eU7L2w0p7EGa9b9d1jy6
nN6F9ty8xO8VSd0E6GVhyA3qOQIjP5N37U9qe9yMa+qa54BBHFa2/lVhSZM5
dMtSImXQwFhUv71jCfywvSPm3IdU5sT743e5UsB8jjgek5drraOXXJFQw/wB
QdCUMJZ9Em2Y/a+v1OIz3KUhqJkG/P8YkjaZvTY17/A9AS0KTAzo8LNv4NWt
quadoffzva50CynAj5xYfpD4xWSlT6ZqmD5N1X2eDQgywV21IPwLS+hGej9A
uXIhVQBtcDslh+Jkqv9BN3SOoDIzJ/mUT0WIzlvNg9cmhXX6cgVxKdTYdR10
ixwIaI8DhXFDaRDgdrTO9kCTN/wJNe8HkozZmlBV4sd9Eb4dTdDGC8dyWyWk
hOAqKhtk7cztg/cUfsXjmzZa5qLNe1V6wkCGwGGrWNQ8xTHM21RZ7hKbRnV6
Twy6kHKhsQC0rqG1hH5+GNZRYg8qECc39VfFbaRb2alen0IjwdgcaA4S7XcJ
1e405+Bp5y9aRwgjpyFeh6D0wmG0387zPU/K6m4A1mvvCbbaraSbZ33tCTuz
UzRaYHz8yjkwMJ5zNLFwhmH4UoQj3w9JS3yhT7z0H+p8TYTDa6aNpU7pi2jk
fipnSDAiFZ+1HwDsDV6US8S1mjNbzQBY0tG4YMrF0w0bD7m9rqTpM47oKg0R
Kz0MMXPhvmLyIml5/nby9MziOwAUPXlh3tBSAO5QlEMzy7UBO1uDx49H8V2o
xyiSODBh/25sDADoZs6VaaWVjEMTEYHMNam8Jeutn7ejTnuoRRIqu1XrVyL3
u35bzvP0BVREEL9ld16InMivv/e1aVzWHKjXPYg2Z554u5bBSuNTz2t0a23Q
q54w2AoQieVA5Y8/WFs4y1unFGawD47o3Wkg1nQVzBlQbAWNELhJXnKqMRrf
/0KCzpmj2j+Qyuna9hbt8CSJIjTgTYSNHjvg2gWnfD0/LcZ9NGi6qxxq1hqX
ukPYrB6QNtJaHOZMrnIwQqLQ66U4pn0OVS9pzex/lSANZcAqEQsOPQ6Fi1Ma
zDDyYGWKr52PIMJPH+1M+kx22NqdyMdsE13eZCMO2OOdGDTgnY0I2NJtKijZ
X+12RhKhwyYd9i7WzWis6FjB9uXHMomI2VwsFesd4BJJmxCbqdIj3xSZkOjy
2GAU3IMnj4XF5n/jVJ+OUb92V0GW4vjg/8zzGX0SVn67rfCClbLNxjVEy6h6
sr94gCATx97JZFXjG2+n1ouf2iemeUk+fVwmMLkd/WAqVf6KdaTG3LBPQTcf
Zk3WJ7WRbjDyvaQLzXbqNItF9x4spaBUvsL97C57XJwf9w89/edHxB2ny7bS
IM4kWD+4g20mKC4OL7AFH74AvIStpOPGGUjRoYNV4m0//DHMKCV7+bF//GFI
ELNwBGbXjMrWwuQNRaEiZL77rMapVaM3FdgZgOos0+KORH0jQejVIb+9hsaB
VDM/k1gYFbAREBwBGjwRt88P1jfv9OPO+1+55B9EbT8CDZr96UGT3OmY50TP
pBcxQ3z6h6/MYhD5zjtq8p/ji6y+lGraLItP9+raJ/HvLn6++Pp1LvFx/fjO
GHq+4UXDtRgX08OSmR63LkYyI/3mAxR3DbT8KvRrqqBdlvQnlQSHf/y0Kyfd
weQs7/xnxFsIL+MOQ0rZ17xMCsx2mmF66sPwSucEjEo57Ajf7ArZ/NfniS7M
Q3HYxE31FXdWmGty7gYp41urSBOZI3SC/KIo8N10tx5cFpGkMqVwvKVvZpPo
nOcXfRtU2W3TQlmS1SFCLCOilykMJxyaqm5/9pEPo0wpgHoqv8jPfNnNXXE9
NNuz3+29tcR6mBVfj3tiamH42dRnvQEpf2q6AkAZk4bbADhprc2au1V/lhYj
V7oaIkLEy1+m7l2Llplas6ihwMR3ndViSuljhdxBc8G4+As+7WgMsjwhQpbc
edsuHyIoURgB9VNUnuZhM2mJiMJnGdLOF1bSASlEigXyV5ddn3+qSJK8LTm4
j4v7hNyzds365jNwqCzKEoE0Y1fBtf2ibYtzI7mFwyjAPC+6hrpLgxFFSdXj
VQ719yXK/7xrUyXlwRq0ek+YL1ItxtEYYZQ7IOB0W5sJ/7DY6IzKD4GSXtXe
pmCJWPYsLxwg1Z6roXU7xLOjmPNJ9o7+U2Viq5J/YqrTANWgrR+u+Lpc2mLC
sHRTydLJocpS5oqtwA/WgagYgDkARIUhyjZAHgCHA2HzpomRMwHRfYNewmnh
BFtRgTfOes8kC8NNHm6ze7wm3axVzJA8PpBmdLypHsSsehEXZ4DJKaHtZxNX
vh/FYPuoyo2TsP0sVVwcPu0KoIU6Ts5k48H87JhZPjhNX4L9Xqt/9tM/aZdr
b9ebi0LJwje0IC59oTGE0VSpiwMFNVOMKYwNNU92DDChGguNSEQVy3NShJRx
Uf7WT4ukB5hz+EhV9zU81bMU4Iy6xvZvA8v3o4mGuxKGJnqUCDTCmhBCzI+9
RW+BwAUBIPMrNgR5cvXCVDMCQfUDVjj9qKszSpEAySlWrwx3WlaXOellCP6S
BYNrj57zvhZYNwRZkQuXxFZfICspKiC4GefnvrgBIJB75HFTR3I0s04OEKLF
ZnKIIJQ1ClbMfyJv0aCT+uEKBxQQBjvNgAN+26r0DT2arLzAZKqcc7ZzsI2x
dPGZMwsE4rGdnViOTNq6F+16XrzV6jBSdHpeOZLf9JZ+7AXVtEWJzzE2wVPU
tQIsgnezmrs7YiE5I/kfYCrNtEnmLh3EjwUz53MT28VHYzoGz64CCUTVjHpk
0q+E4MdNMJe8prW4i878sRrHzfNNr1pkyDtps4WQG5qi+EuAu21dlETqDU/l
Y6gzPPKN1UcguPs1KLLhAICJ50zjccql3AjvZdDz8PsjM3YYyZZl0FBooSa+
+qEdC64KAn1veUw5qUrBSSALccmD4TWb7aYPQOvTlMBC3uUlfgQUEk/t6kSH
vR+R9Es3fVJtE/e/vhAgCLZGBur/j0SQtCzCC5VdpsFlsUCKHFJ+FwhjoiMx
bnYkxkxXXudDdmuiiFdiClDkHSC2yAPggcItEJB/FCBumGm69Ye1AxCqCFuG
GC4t8g7m9JmCn6hmgDN6NKVRRgk8Az12MOI+2E9tMvk7QY59wzOqR9RgzrGB
TPYW1fC5v66LfBy3TUwvjbYe4HSBc7asaZEEFMH1cRLVWzbS6XwekR3XHxsc
nn61lYOPgBhtREvPkYWIDT4PCvk0l+hM6EI7ouBIVHh5J8IeWUyVWMw+2oIu
85ZLZxONuL+9MVcZWkvZnKuvAMsbHG0s4XEwOPAywrdGIdfUeszvWBWgCd4N
0sxkN61dLs0jR3oxnJGkX/Uu/KcofuNFE+vayb1Hy524uHLdQhb9aO1VzKqb
Z/21g+jUPh0ce0bLCndlskLeNdwAQIcjxtjHRIkCmldbwd1tK0Rp4+9hHkHW
YbOl2UHa6TZhzT9a1ehwLpewOHnRy/ytoc7YbEma1HF0kZ9Ot5jJvrfAWXsP
u4D5skolmBQUYCWgIrae1bFDCWBg+8NhWMjg4K5BQPNrY6moE1zwreIKQp8v
YaxKQx7Hqy/j0wOmQGIAhiYl2kZoToqHegrvZi2zZq9Z08F93rGGMDTs4Qra
UlLnQNDr91M1HW35J+TCoVZU+FqrrC5+n0nEtMyQy5HUubzRXBQEaCZaEGtq
xg3P8MKTP064KBnHZ2BDWch0NYsPiJpimrqPadxnXUywvbjhAlW7LDmcm+NB
qgboCIpg6UZY81D07iJiephshTUK9AqAhkTkONyjlVWFoddJXREOCQxVe1eI
1B4zaDKHvmi1YERMOz6Pjd3aelUuEtFwUwv7R2LMgwj5vTs71EHx+cZ+Goeq
RRTB+uJHwJgerbhVUttmJTRMKC9KVZT7n6vJ4xKHmkttE3NDMg8pLtLgqQLM
0e3GXC6Jtq6TYLBovQiaB+ngGCsedHTjPvbEAfgmS94QhEEwhW2ODQyqetg4
jnDRvhwYJv/X6/hAS239LPkVNJ9Roizac8syRnzTrJtUwxu3RaZdme1AFwWC
fTuiMNhY3n9sP9nmNi/1gM3UQMsY2X/cmX4r5Fru8jYuUAtcyAOBwMZJHmHN
q1umPDiATr3Pa9CAHzQtW/z65aHCfB8qDIptUMIgNSAiyXbGZocTFl1ZWHku
WN9uEKnJuZN6WTaexJGmOGDjnGCU2AeR4oE8h2Ugx2EtAbXvqDNIzryWABQB
K5U/Ttf7ZIs/SwHX19uguEN3wS8WWv2sSLrBYqUeXqHmCmXlcQ7hStWjQWOn
eOMxlBQw9MKqjYwo2Jxb9OYH6OvQ8T84/w+ahk2GfBIFNjNPjhgRAJr0pckA
Dbps+yyl0FKw0SQDbVeFxowwntqJXKICgmHmzWIDQWNPpNNuqPC6qOV66JR9
yXMKdey0kJ7n/3ClY02/7xbuxVXJ9OQtFakKHXWyD9CrYTuYLFJ+bWclhUNX
4ZrIWyTiXqsp01MMFsQti79lYXrirbdAPAEAY8z/xZsO0hw/Pdi8DclbAPZ4
AwWgzsQj2SRNbhabdDpy9KE5ohoQpj9SBA5wY0WWxjV72EEsTrVfect5g2TP
EwicfpOelfXfw2Cm3CYiUCr6O5pFyItGNF4Or6oeAZtF1KZmR7FHCpAiQkpN
tdq8f3Q/G18waAMx59gitNxsGDSkzYIxFqi+IIM9f3uGC/kL9qbUbHC076g3
0N6vSX1TN8h2jpte9KjAk8XPHSaxdDgFuxvjCLX5t6pZ6hiJBgy2txRh8T2c
xwUQ0QmF9IUyT1CDWD3BXCj0HJCmZ6ug2sFPaKAOdoJFffeXrl2H8QSYjFYH
042y6eLYidtkbI2b0z99sjZV68pDiSVdqnVa0yHJJHRatVqJYd4h0kjzwRZ0
o/urjalOhtqvmnIvAq0IzVdxo7Mh76otUpmXqXYF9QBuqtMTgPSBCHU0C4cj
jwTistHtMM0yhMs4/lKTpZUAUEwygQT1lUv1PyC3qUTkufRFb2zPtdqfYbb5
nq0nugTJZTeF03ojkY8FGNEjueXD04yJhLdhjvayFzZ+AoccJ7ji0WrAXMqa
dMXZXRJZauyS6eUBDFVdF9DpL3J8S+WmIJY20a9hnWlSc/GLxUEPBU8gVBSp
Mr79YdDLcbApBMrTrec/6RodvTwiJY9EKXwrG4ShoNp51pHUBQw5RDJDJevQ
HCcWybXyNvbGATeUzSf8ZFAxCCetOPqM5QByrP9wzhbTk66OdD4Ri3pmhXim
+tUurHrfuNYH1a6xa1uDKjzpiUiSzYw476d9gZzWTMgjZjGSfMiaSAWjXYDL
XK5CqkUhM22bn6sWr488CoIdoNP6fumaoq4iKDXKoq0I8WDetXLwRvcEbFpf
Sx4CMLu3FP1G8OypeTZ2tu+TzVO0Ddq8I5nMt5qK5HRI3mN4mZBUABe/GyY3
OzLys8U+L/dTYEgDaAsM+SP6HQka/b4tARjc1cKtLJEuZPDUqjtfqvcPlcNb
YaOYFuhb7k1AKeya1rgFKUU1Wt39MPUb72exNzz2ZgJjEPYOFqLxIyhqv3j7
/I10kQNUSAyfoKInGs+95IEHtl1fwuzzJHv4KsomiSeLITMBHyxRo7m2M+pN
Z4r8DiJF59fKO9MboDQDAIquwPII0yLv46OW59SxQeDLEvhkBvrzL9WQoiUN
pHZdCRYgAWvGWHevvZeTpdQitSpd6g5GVNsyFXgRY+mvSYqVN/4QABukOlfv
KBfdm12lhU7woueH1JM9qew6pV8vUxYzA+6C3qtydC/OMKiJIjvVwniAdIHV
7ZPbWYeK6qFFRWUVtYo7V3cWb9RcSaK12Pjgst3w5yuB8IcdBjdFfzQaTBJl
5zAFbarg0p8yrAD8OpnqrH/ZSCOapb7+BLz5vI4VPfodkCuS24ZJtDM3cgjs
OImr5x2CoZrtZwSnz4ywx7rkZuqDAE+24kEBg203Vho2WQU1uQhdoBbOyfzK
Wjr7I4xHxZUfPmxkq3446aQ5DvIRs1Ky7S06D9vTOD4Fhzk8qCNg9bau7c0K
LMqLSoJZwtc7Rsd/M8U5zGT3Q8E2JiSJgwh6SFrxcZJOD+5nq8KSs+wOxsvJ
BpJJLoSzVw6IisSX4sNGJPtoRMiLXUKbDepr+4kb2vfv/1YqSK4xmdc0v1oh
L9gOMy0gxhm+kUNhM7cLVxBiBoJ4PKu2Ip95M+MSYQGio3hYAVksm1n+xfNT
VuRzc07RAC3/yjouL8tkVvuZp4jyGzbGbzI3KctQ3ZaYC9afUjFO/mOcKYzX
/5Je45hzmqHSOeoxe+xpsFvjANAhr039D2ywLCMGimWP22/DuzONKBpLVBll
lnK9bGE7KSLOi6RDUqSgNubA5esGqbohAOwRxWFuxDc8kli2tcyD2gmTrOzM
3PiqsznjuhEcX/X5mYhwLsZSGHZAzRBoZfW4BZEEU0cc7+2LU1UIEtCbBmUR
qK4GbIm2DuU5Hs77JzsN1rA9lNIJwC8iwJkGQdHcnHCLqnLpANKneV66Geim
XN8RCYjTh+4n2r94Fj+8/jhVjErCrg1uKB/I0BryqRS0cozVf1gcnyj10fi0
TH7BGbweviInqhi8miA5No27jj9WZdj4skFbKX7S7UT8+1mvnx1bBH3FwnyF
WBBDT/Xo9MNTiHSjc18cqhl/mwiKTD4x5Aiupve50/UFXxn31bvBnIk4gxhZ
ZkLMeRMuDci8A0IvtVHRXNLoZGAenBClEg3pdSVULVRZZcxEfLLU6I8Xz6PA
HgNmyMmpJ7TjroM6h4aXmqwy5cejbo91W5eXf7JULBfSMi0M1Oe0ggs7Pw+B
kEpBiFWAyUVv79swu+vjfIIwDpvQBntqca/v+Yuu3g1agjR7fh7fTqBr9JRy
DPYtIcPIcuT0q0X5VMy+0bA/PWqyTy4Bg8iAOANfiYzS0XOEyndPJ4Sif9Nk
A8uwkC3tburaBJaVpPlUflEX+cOyWNf4OOizb4TgjGz2awTrPu+t7rGeO8Ax
x8AGAv7/qWfDun+lx9zLJ8rv1Ch+07SVuLEbKQn3zOzXaj/aNfSOetL9sdw9
UrQuASpKW83gJ4+qkHG2jxTZdHYHuF6ClbJo5BZ8wWtLKueQUs1canqtRTsO
AcKZ7ML0N6sH7CpIJ6lOItZfke7sQkFwc7sX/AXikNmiTRdTYOX02rqahCEC
4pG0g+IcEgw32OADxdcrKTdmqutr5fCyQOt43KelLlQAAR3hc/mTOaqEl5iE
7XD/mAanXox6BAiA1lkvLxfzOr6HsYq4r7cbzmc6AJ/U0Dv08uwVLF9iOHme
tPQaUxiAyAez7x5IhsmbrODONM47B8kox+1LpPULmQUMZQGh7Fl2yKAPvFMT
MgXq3uCoM+WXbvNw9vSpwrEfAJU7UEF/oZyoBji+MYjTGrkHkpT1pX/tJRmp
3NjzjGu+3czDzLvkZMY30v/UCBjF0p4a+yEsv/okN20j6ZpGpsAK151sCK8D
LgZHAG4en1DkvmwJ798DBGWCHmKg1t9P9x52rAFxoRc7VGuFo3KjvnQ0MQaS
ns4IhOwsp6hhLl+miCifHwMYCi/FE6mKwcGigTle0CVoNLI235M/7MvaAVL9
iBgjPeVhOyKPp/pkLpmNBEyWS9c9GsSZGH5VHVmvdfds5rQRmW6uwN+z7RCn
BHkXVOsUcE2u31CwUUa/h9y7jqSMk0h6Qt4g/liz3xF1nHAZZboBKz1+vTu3
hdQaKjehz6yRJqWq19EKILfs/C6sTiiQ+sBzZyD4W4Q6QCud/aT2tRwdrTvI
SwH2J0DvbIRZeZaHr0Fl53qXK4aSD8ZoYR6lNcXrqRFcB6uaqKl6t4igw6H3
cBU7P4ZIf+KoM7IalnXdRROdtmYRG80JCpq3oyUih+280o1U1Ek+XEdIPzPC
Y4URI7t7Stcr/erMAiTZROEhiHl3Y7uMibVrpKygb6vK79eiV2SEk4dQYzIg
Ya9sb+K84IZHuOJ5Xahb6UrozX6CDgjdOvZUQemPvq1NZ0pkLPwQOuFo4HsY
qUJhqzCPaUYikGpI0w+wGqHsrQhWITqNyL88m/F/nrVaV9uAykiPMZwtsY1d
VsjgZEgmr3cy8YCqEXYv+WyUB/DqaIsLacEZnPRwvxIjbVsZGydOLwV28ekg
kZCsCtHYmwooct6Mb+owtyoBWJuhUMI1fJmdAvPqr4gcprkgIWNmDF9wBwlk
xz7oq0U1gVn5GdG/p/qQbVdVr76WoyNiRPd2okLfEOdfZlFgzmhUARrAf94i
3Af9xIRtt/6MzuXIHjiIP2goGgSA20pffgYiAU+P21ZMzU+m5W6bXVHb+bbd
Ph0zwTKb7tz9UCy9aOhfymb1JWWDROoT8RA/HLM6BM0h4k6zQl4jtUFFasoX
cQZiICj5U69cmo5VBsmGpnEnsczL383TwULqtRTLnA9hwAPJX4wzuhifKbCk
CyBnRu6PFT4oJz1zNTfLHbaVQA/rvVTDblOhViwlnZAWbH83nUnO4c6bRpFN
QvX6uL6wkrnNxI86fB04C3upAQqRVooxqBFOMoI0tEKJjihHasudvwpm0RIv
8r00FfsORjPI3m+0urs+tBEIQHf0SzMg1LOpQw5tGGcWGVvWWHPNJkBH+nfo
QRdt1CQ/fprAyK6af66dWFT925H/zsWJLjOb3mqs9Mi385xZwh+jMkMJoDu5
ZGccvouTpVb6dhlV0JRM3ijroUPg78Xj/9atH4lbwljBeiJLT+d4e9IhVPaH
KR9hUHfUXYlE7aXCwcIea0YTa7MqhRS3sCatKt6tj+EctwXF+Cv1BfDrgHDF
6c5cI8qDFS7vfM+U2MDKP7tza/LRDfWMQA+nlGGhwzdKApZP3OyQ24TLUhb9
oR2KBwiSARARNOr4DkMKXOfsZ/qq+VMB222PjbWyZ/bHRCDXwhVnpeEMwFJi
OjUo6XXRmjHCF+M38Nv3oSAEw5Yy0Mw1tUIO2aY2IhY+knaL/PXfazbqCOXn
BetfLjOL4dK4pae2YQn3wjRAm+HlRm4cGXP9xkfWBdDkFc5WflKcnpItjcrK
ShOCA2uptfH/uSKnPB49NauOQBSIOrx9cDIARILOVWDmErrwRdJK0Xhb6ukH
mqfAHJdRlXkth4WnCmefTt10qqzpRcWZKPNnPzK12uviEKB46R2lnl9WV5XQ
1VjetKYJf8wBCnohR0PY6Wnp9At2TEkiCwl/DfzpJqaS1JqgAFtzoKSp0F04
v6AS+yu1SFcF9nB/qn24wwo/vFSg33bzeor5NafUxm/9KvxKhyC8IsOICsW5
JhWinISeoRQc4cARilAqretwsOWp2mTBwOryUzCxD+EVhFvkMZ+BAUkvxQEy
Zjo5fgmWGs+T4TIhziDoUKvVBOBeSloqArCluTgRTZerY1k6tUB9OfjpsUKe
DDPgNG42qlWVq6rH/N3T6dTYVWumN2eFBUNQ45DNnZkGCb+qqLLeSltVu8BC
1JWodXdtg/yYoBrjDS4gkzYtKdC7cYEcyBDFC/XJvyCh3zok51GL9hTyo3kl
PyRSWoML9xlJ279+1csfT3T5QEZ2oGMk0kYLOItNXhixNF/TUqZmzjdoqae3
0yxzFXsesIN0E4T+fQtOi3RkwSB9Q9F1speOcgdvwKiuNYOQszTGXcUhmkOM
pIeKWHTX9InhSSXkb6clSJ26lnc5cA5ghpdh5ayxlxbu0g1oILWLWAUoOl7S
G4MFVQfh/19ZV1XlyhzZfV339V7a28EaLBx3gI3Ud84qmUrrsQBsxgTqJJtL
yEFG1tINgooDeJG3QF6By6mOnNEulQVRfOUbGwc2+H5+jXjpA2oFfMjh0MOB
Zgc4DkT1tF/KUexvKxUICM6A/42DFgXzVmFCvxocltJYcHqI4zaFbNMvKiQH
ptQkTcPy7LTir+PIoYxaev/A5+GNeU1X+RDeEX3x3Y+dTN86hdxM+0nApKnD
5hQCodXmEMFC8OR9E0pN8gVZ4R8AinDC4+kxEck6AyVGwEF23DgdJMb+H41k
23r/koKMS2nTNF0qfv4ygVAvhNpGXbKihfuvXetM88xz5/fo/oh02akhvEnx
Ixgpx6xgmesF35t9WKRZhO9FdQs9bbOefXY8EvAUeY9QdwCsdu/oVqIJYlir
zoJBpKgw9INDpC8WRHbVEtKp3haV0UJr3mvp7CqjUT40Hl0d/fSOmZtSKp2O
BEbB4PhHmi9DiFqzltaFf/QdYtsytfjLVPI2TQKo7asIr06QSx0/sk4/3DnQ
IhkI0DLYMr6Y3/BJrdKPLEPqTljQeUd7DN1Fmjwm6AHDxvp1GJHAIFn5z2ar
BV536sq4AI3BCEgFhYzjEfd3+4ZT6FSVSQ/gJ2p6QiZn4dB0TbDzItT68WtI
fyIGbl9638cskhTpK7YweV2rxo3ktzRV/Y2Dc8ud3sioI4X0v0tT+UP2Lmn0
iWjAiMI43fzMoJ0mLXR8SaW2u51n8pvsz68vLj0hUrtpWrZnCe8n21loqZ82
gUBLwXxGmUU89E2MayKzfFYUcGb3XfpHdySDK8tRaBebtlvIkdjlhgU+UsbN
084lILy2qclLNhUX8hF2/1EibSKz4XMb4OHG2gXMQYWLGwsishTEFyVsuGV8
GCK1zouGQ6br+G0BnhQcoekCAPHbxP9Ve/yqpoEeVt1JazBFjpGGr9e3WRGs
E/MrE1RIBzpTa7f9VyvyWf4+FAmRAHqwqZ9IYEv+2V2rFHpBKqanCTreLXKk
uyco11FRbVaqCWBBaLsGp2YaHaWKwdNtTr5MqS5WjdE6IvJV1aiQ8brlAlFr
G2iNQG0COgwbHn2Xp4zUsBENOAnhHD00k1bRLpLyxEpJWm8Yjr9fLrE4bZcb
f8oZYsGHILT1kbwUo7lFu5Lvi2LMDM+XE/fbBKXt1YfOT++pmc1GV9SZZvVz
6Fblf8fZuSyhauvELZ2iDwohasFI68HgLDRjl4+NPzHGBAA8BIc8jMWAredF
ZKbmUhGXGXavGxHkRoMFRKT2JWUzpQxpFT172h1dN+fUmU6N9ThJayNxtwzi
hzx502wVbC2/wur3e3/Mji8pBsmWu1SmuXNt4Sgfc5hRj373mOuNKmYEJgNj
8HAgHx12w22whzRXeVjDr/sVoZl+9MLIk7AVOdVfcw9Bghh/Bn1gtnZU55jc
pIawfRa8xHEpUSq8rjeRKiCHzf39F6dntvVcSXJmlVbJm9HJaru1wA1qdRsD
nn/iRq5oSsOLpfB2Gi1TgR+oFLEJr9Bi/JVxNbSeox6KVTYm7NvLaQ+C30Uy
BX/0sFQON4JkpdZZQ36NsE4uU7jsuusApuc7ViptPqgBJE9O5JonLF3eNqwZ
AU+sGv/GpYwwRW9dCTNwy29zpEapjPviYu7VCGXsbvy21MQl032zIi6o1+19
+qgEUHdUbV74T6bVQMxxP5zUu5TEgRbcCLAbG93JJff5MJTS9Cb1x2czl8v/
R0x4oYmqRm9OwFH9Sg1KnExxLr3QBsDqC+ZZJTq6rHgfDiimwDW4e38Tr62w
eTzOZhVt6cqjj1zVzDMrMxXZyPdO10ht4Rqk8UnFBJ+oaRdm5IjKJsi6eI3y
2la4SxolMLyw4MqtquHMl9GaLa0PxGBo4gQyZLGQDYHYOeSiiZ8mt2rxNwFQ
ZKcJ8aeGT/N7qAZVIwSVCaSAtSXeb5Jce/MEilnaT7sqZE6L+hsPAuAJuVRA
VMab1/x5qCFR67PXtlAvLtevfMGfpqJH7p+HVD79DyY8N8aleTvxFodZMPpm
+ZXFpVSPrjqVXuTa+72wPBtwS7UxklT4VCWomcKcrFB+xnUphci5IijSL5KZ
LYztfAEqPv6SemzP/mggH036gZRdm0x26Sd1IOxpW4cmvWAjCbBwpw+7n7F6
wdnlHmkDsm/JqZ6IW00+24Cj7f9BlFRqtd20gu4QW14iEQ2XeUbcZuXxMrlq
5B3P7XxD2usHfetaHgl+58TWXSLrt/gIkfH/CbTlnUX+oZvsuq35I4dsZh+3
AAluoAfM2p98AHR0k6GdvDrpgrFduYmvqdGwaMuSsjKd4gE1Ubn6c2OT1kFL
URctChFIkVcawNUA9vlPJTnoiNkzSTrTo4SOcHoizH4uTikwjBD6VW3tSY8F
ICd9KdigHeR8yXdivbNo9X599z01riwDVw5FtS3da0di9jiu7+ntpV2wnsBe
Og07Rc29d16KSiC2A6xumB2Aq7efblB8evXlbXl0rVF9MumIZkEubm1SmP6h
UDrg3vM7ptw9hOIdl5K4kxhcES1JevkTBG8s9Y7SRW5qjkv6lrREt1MpVkI4
0HAgqwWGIPaZ61YBw6is2YnjmBEM8MX21D3puFrdID43nznBAXA4/+ZwTF3f
kU2n1DACfJHB3lmSMGXZQBNpkVfQ5uXcOqRzxHSvoIV9WOWaNCQhBuOtH7V9
cR4k/MKNa4OcTlgPt72TMXhozIXMRQOTWBAHP6vGIXZzPTQbOITKVpCg0DBX
XcshDRzzHdCKvo5TZBuCItCgLlqLc/NQKd+AU/I9/hp7rvHvjMlIF73efk+k
TSrrOoE39wUi9A3u8QIXL/SoV4mlr4f/TXrDfRIKIg7DoziTNwHLW/N2cEht
ja4wKvFrVJxkNk8K9XDLilzHD5pm0eLOF4WZo88ooJGJGC0+RMIgkDqVUcG6
RYr8nBEHGQQVyrlxPrEMEYwsujRjqgS0MzqyGdY9ewZbXUcz1KmvLVYUj9r3
NZbXkKCpAqVfFNReZN1X/DN8BXMXCLLzzU/QhLKjwnHO1C7GQwt5SXBOITJY
qSGf83gLjvlitgyYInCL2iF0K29it6IGnJ7KlhknytL/IXqsqaZotYfKmXnQ
zvtLhHwLDaIOtGHLcMdHFM9TcwIjh4acgC90Bsq585y91XPLOmgzjHrLheYe
CXvaCsdUc3LMtyYF6OvW37lrim6GDAFMYtcT4Bafx2Bt+1QqlY/VMd13ZgVz
blVa+Lo+iMo5ec2ggwEGtZaD/iiw5nQ3W2uHUzQ06Pgwpx9gGj92Sa11tbEF
7xvoeKpoltVupNtE0+B4RKgc/cZzWtEFbGJEmPmKsSe4V3riD4x9ibXtvrjg
H15b3iDjAGYzlon4sNUbytcgCCv7OdFNxfWkT5fQPRYZ4DjeW51Z5e5q9XEG
CoKERqEvGZcNPlzjfkODePD6825oxznkZdmuxIZhjMl9A0Dz3LasF1CmIR8W
DYCMUpCghaA0wqbSUyJFrsUrOkbfhOdieM86eF5joyuhCY5ZQNs5gIlVuBcx
zGJpZabtq7VKdhdc8QwCjzPkiAXIGhtIpQdOfo9jEJdGWUwsGxQ1raOs/Prv
fTmO4G1xrTriHKiApb8Hrj9mSdZRaYfHF2aklORqj1jiNGh05yyxTklDiDRM
aoEj/+uhRyTK0J0atSz1hA/yh6pzIA1YiiAEB7y2eUG7FG00/IqV4id4qdoJ
4RohlHcAN8EkmSq06Do0h4QC0cNcjcZtNvZ3n6YCkfx35h54vMlkGt31rAmT
4oTrDUYlkRPbbVk2B8R9Ol50Tdn03Ov9sYwQnfv236F/rtR+odHlLBRM2qr8
hpeQvgywBXLN6CBRva1UL1P3dGpaUjf4fzyu4cAWfqi/MR9/W+kMsDLgxgqZ
l/czjHe042GUzLV37cisDLJhTqKlg6QuZWNu9LGdN45FGj+JnaXLvVSgG+NN
BDfGqfJH6q3/2urY+JtUeXbx8aMcJKJOwDaSmGFewTbqH/PofhbkKEntYuHK
r7eVdy1+gKaHaRERFSnv7w1lqTaDIBn0GeKcTT4cItVYjCJI1WKh3TwSvSXv
smnQs3ypmBCFPjESN5JQBqoNwWhwPIN9a3/sVBEG2mxo4fCsig2JIe9ScHIE
amano5gwRTZ+AzPMjMjlLjHjdP3QIF83ZAINzLRs8Hb5bIyHolzmWZTzuoFC
ORDpIkTsnHwP6ZkEDl4ey0lwL7dwi4z52P3xIxMaS2dd45+gdV8uClBiS6s6
55X0HNe63rRU9xP/VxqVYIFYxwoS5EDK3q244gjc6S/m7MadBu+o0ES/g2td
ywCWYcmeHg2rrAFc8CAhKqjOrfsl52wBbiL6NKqAV7se2XIABOcfjuhHNqba
E9Y5c9MABfabHwym3FtS4kDvTUAZMraIcVRuF0BYKiOPioQ56w7tYTMNJGEp
Gbt4vAo6jWkXcwVIZ7pf8r/lhv0jW5+rczF5oRMa3esStLsONirBUzu1DU/P
lsy2kGUv6kJA3Ts8zEe6s1Wre7K5xL9mLR6DQtpo8SE43AYi7HAkDTnMW1Gi
m5QDHTDHjBxZyUa1PZKpd18/HSHSXSRS6cFhNZEX3I/H+RYqY5geZnFRAYuA
24YSiQTYCcK/tZbBgkylZeFTXK+gjx9P0mvqPdGL/1xkg58a9CWZ4pfDzQa4
o8TFtTdIOoLeqHQzvitjajJB1eMdSnm0DTJVOQcCQ+6hac0Rb545WgZT5qhV
Aatcx0JoXls6brLtCzFGpR8NOx/JhpBHjtbU/yi44cDSfJnEfpUnS2rr2LCg
pjtlFh37XPUzgZX9bnYIIXEQvjZAbCqAUgjM7/HthqONrbSGvyJctdoSQEqt
2AKFxOr0VsxNGQijxJnYmp553YljMBGo3kC1geUe6Y+xbJChmm7bG4BP25bH
RC71SXwjPN3bu/4sYD8qi+XE3mSWaLUC97zrlxKVmmHSEAa/NDpCc9YRQOHC
R9JmK36qLnNWw39wi4yfTyRZejo/xui++2XHqvuhIDy1KAKO6dWQ15At2oyV
UBg3uX10gWdEiKMSHdpXtG63YTfUpoSFnkya1rGAaQrv9g5qqQD4NZmOhAFS
Sv4RE7GRuBb8DNfQR+vJZ1D4e+trXQOGs3HBwtgphuNgze3MFZy50qA7cIcN
5NcnPu+uUdhOi8R0Tr7OA+Cs6t0cLIu1HvQwviyuVGQqhGFmh8tU3GhNzuvj
WrSjPAzJrJ68IGzdwP+vOjEELO04uOPO7hDGGNpr46BPfOEiZaZ4AF+Ykj2M
Nc8OUvbFzddLHK/x4qJKTDAY3rIlSRgutXsqjj0A1DX1ASc5wBSzle9sjQiM
LT9ElcXYm6EPXQCWj2o1Xpuxk416DpK8SJi+b7wikrjCMh+y39UO3OvP/+OC
MuRwAhsazzzPxWWVawOoAYQC+vmNu/UtJ4aOHd7nl/6zBjeP81474lh6ZGjN
n3PoUpSee46ryBF/HPu+HG1VXu87XsEd3lw8EFKazLhkD55VdBmozfdJ6fwu
UZ65BkJ5xfGSGI6kv4KtvHLKov8PS2Pwk7gnwdG2HmDQ7kKDm3KdzN44x2lU
zkAxerZzfdoFbrxy/Fa6OPqHScMG+mt66amyPfwgOfQdrGeq9udFePqMkVMa
nwWtIgST6RJGc3OPF/MhXX79uxtiV/prDzbIwTXdENsL71H7EOr8hJDR5OfH
M9d1KBqfM+dlbaQEPwMejOLflv6A400fUnRLamST2aP1XcYmcovug8JWN1Xo
+SWXiUExSVfT1TNGMEyEoF3MOChMqGP6SC7sDOs1Apb02y7WVuuwhzTnk1rF
hY5OM3rWVbO8qLLSlNzpvOWQAOrylfIbaCn+t48cUs8lA0L2HUVnO/NbFKKg
zPYwQsztZS6fC8T/DY15rv8rnHGgggApSsJL8L1amHwKuFvfMwERAqbreZGy
Hnwx0gwiqJgs9TwOnJJ0ndpAEP70N+9ZpygHMb/FaDoCcJpttwhLsRvsLkUW
sdCPb3v12pfsNKz1TxZNSIjx7XiBwRr2OQ60vUnZ3BEdf9/dTsVgW/uRuMgV
Iupo/XSzojTjRHcD3OWeU2qtbh2N2oqO04rnPpxfQLEqjSb5RY70XWzEE2e1
4oe23lf2HQAeYYtEzY3eSqF82eO7djyPVVe0IuMYOqt85iSUmc6qEowy/N/c
cfH1L8E6TZjwxFJHjs7K51Dhpd+KMWyEVmgKBKNHxcPQ0vB4DdlzXj75ZhPa
5a2jIrZHvnyb3BscDEdYk5Ll+fwMuZLfkZYVRiY7M1GoDiG9TQigVwpA4xLw
NJwdt3OOOAgclYiCDE5Pk5S7Ui/z9pdnaFa38sEfFSfIEaNLEx4BIWnBaqf+
KEehx/Yb0MQBqHy936tebbYW+GO48AxTvB1DXlWluYTLCmDFFG/hsCXy2t40
MVYZSu8QlETn0uqNwRe+Z53awjeGIE9sHceg6Var1c7YNYrC4wC+oyI5E01p
c5Cp7lzGAD/E5R2PShJz2ymASf2K5b87U4A35USHYDDKlPa9rnU96u38EAVy
SW75EXhbSjAB/Vb0tsA+be5sx9DCMWezxStB9ncl6ac0zEqqzNKuAMeWTdQj
gDdmmZ0eKMV0Y2DOFBad+2Rnu0HU1nnZMQNVBHt6TSFFhtRkjeC9c1/RGtyl
aK4UMTB8rBJs01agip9LH5CzI6moC2stRTE6V06Dbxc6Ny6S4TiYtBYY3iNl
A4YvnvKKeKWDjfDdexkPTZe0BZF8esYL3p82HY8zcDeWfGYexEWIjUK6vWQ2
dje64+0mI6Blp2LjlryHWKT8HOGDojOfv+jzqWtHTsxZtxCGk6kATrBh6oJC
hhGS7IZTF5c4YGHumHAdUSbDNjax8qPfG+M9jPDclnrnpyiCdVDbgAvxJNK2
02MUo3gkC93RjihPuC8f0C29o0lHSG3Doh3dlEVkAbI1TBMyyC9Bwswc59C8
BRmMz5xfu360lJisH/tt5f8FHMu4DPR9DmuZptlrE7AuRrRzoaD4ZUTw/ee4
o0J9LBjg1Yd03dQjAefG2cUTxLK327BygZo3sNsUtp5Oh2EWL0c3Prf35Hxl
lifDGDVzd4FumCON6h8M1jxROLviCe7LYh6JgwpsqVU0CCaGwymfNpvguGzf
FezcUz5orjwscXvOP2izmoYF/c34CsDLTWq75pYFcHpOWqJ7dKUnS7f9nuag
qlWrQNmAUQqVns1JSelFFJ84YKZFES22+BnWm2stOlJRZ0JZTaoYH1rm6YZ1
lJ+vEnd2qMiqkGGN2+d8izYP9cvk4riFv3+x5CNI/vdr26DjnW6noZz8Kqow
efZ6nu9+8DyEZTBM3zZSf5GZ8oir25UmLw4ttmsMGVZ81Sd4dI0siDvNEslq
4XNz0wC3YzJRw9qCiSBXq4Q/vf62poBL+ao0q95h91IBUQRm633ysDCtdcuu
iQFmUO5mesjFVxJXWq+OJBAJMf9uXBp4WtKkEc20POYCF91IEUOk98Z2L2h/
2xl12z9mOMWVrwbpoOx8np3jm5NwHd4JoiUAlJ4BplhoP9FCxgfbHUrLrnmK
XQwyNmQoif8VSoKQKKJ6d+MsBmZ2gacY9KgzsIgwGrqsfAeqmDaG4Yytc8Vz
rskShZD+l3qO+qxgZpKbNtUYobxgpq4eMLfxJg/NRA4fWXIKN7Bia3knarLc
p6pD+rYZA+tDFSVa/uryxUq4VmDnQNym6PvMRGhJXy/8sZYCveA8CVWuCYs7
7rhDbGKkybTDD4iyyWEaAEDuRHobnS9ApsjekB1n84KZuDNahETc0h1V69LQ
7Qe4bPbsSoLwJd5sjvCuiGHQdtyoiekHIJ9CnQ9lSY48zwvPxk8s2sryYwi6
l8ceQFmN/Kt8cttM8VssB3rXoskTuXEn8xwIibzfY98CxaoNSgSfaYEdB18M
A1c36yuTIJC6kXH3KQ17CJCO8549PjKIA6My61G7X5Ta2UK8FWCvdJsrD5fD
ovlJGh0PRJGRB1JUZmj0rhATv7VfCVW6eP7nVaqziQd37PrkTEbESr8Oyn+R
5qF9TQJqkPbgcByu8oDdE2vyE9wokDCBiwThBqq5DlgAhXGwFaARBlM5S3y7
eISjgvqeYc8mClQiZ+KYva7ir5TF9yVAe83Tx81lq3SVnEiFP1hS/VY8Y3/7
Pjr0qY8nS3y9Y2E/qEdxz63zvvoH9suodNeRK6+seTEDIjW4eK5pWSRZNv9q
9aatZEywGv/gDICJzExnYrv6l1tMpuzQyvAqR9G44Z0iOjJtAc02p0mqYhpZ
h6KWKFalq0AhS7y3ZGxKzEP8TB9ZAqyzntsf3tYAXKS7Nvq1EXmE8Kx5zJGG
iAyQYsLE87eRMLUbHof6QCVHJSWMXxmKKxb2vw+KZGcMYUKpNXG1iXhSDU0Y
NT2od9YBcY3iqukSh9GPLEItlMM2SJUXy3QKKD8vo5Nuhcdr1CcvDeKqE2Dw
+zJh7nv1xRKMC+dzktegzfb1m2g1rBaKwzzkM8gFd/e8eat04w5+rSqeZSgL
jSQqe6SFEpa1f1iygDc3ncjbw9g82qK3NmepVl334jQkYVzVc34SEdD88xF+
NCkmZ+Qwu3xRrBC5/OqLjClobk1PjQk5ZN2l96euzuc52aduPGHTl9OHbzmM
KKyqPXHlfXA5VSBnAzrn5qNfkPXaUDrCK15AyKRjltoTZ6UsbaH17ODEn3bT
djI451RENCj1zEA1v6VlyKlKF4if7gMiRZzEBhqJXwrwlxJcqsgEPOnMLlfJ
KOeDNfNyVpRDbOW6JtyR/NuXLotesHbeHJIDz4G+x2lDO1ffLq0pvUIH00v9
7UqPuHz/kKUIuF5X+tt+2SUf7ZMN2e6XeluIwT8s+/c7Bui5w5KOoDG1xNeJ
icUFqFL01cEyWJH/137upUUdnKjzJJlf9lP2NMBmRc0BF4kMGOMiW73v+0Pv
fnjE3kp7nAGQ39uvszRdV1QhAmbKGS2uhMkQFzZPv9xqRHzT0/XETqVXV4Vi
+4NyWsjWc2Wxe92aLnIROLZ5c+e7vneylNnUT+uwtFfZCMPO4DP+RRhWsr//
xNEYbpaGsgszRP/sZG1O4at7U/w9c/FI5adLdURpU0iYs+okheqgh1u8uc6B
/HShsWSYu113Ie7qGUJ/Mu4rib0Zv2OPVHu6Zsgi3OG6+8P4+Mn6usVEoEr3
NAZxZkgltC7KRBiuraLlFR4pZpTiwuxfVW61OhSXDEnncSvFIeZYHlL5jLMJ
XAHj5dstOCG9ghC6FpUouSO6vPNIo2IxBYJXiJ++/5Yqx1PiUQeWT8anr+Dy
7iDmBA9YI4zsYqKNJ07PtnsV564tPLHdk2IeBzvNGJQ0i44prsnupgFAPB4t
m+J5t3qe4QgVkOQmbDaLjTEiK4vjR915Vm5GBQNl4SzABb2pkdi6cCNUZYZ4
3F4o/utRlfvwUV43BWThbdDFmJNmXxJ9tup84kBD19QzjOhcXWhKwYwbiiyb
pzHgBxmtsbj0VrGp3fBfUOMr258/GIGuq7+BoDviQQsZHZ/MULu1+zf04IQr
NEO0Vq44w7XSDK/NAm6XjADC8bZ30vaxmXyVJ1HvaNDzlkI6KG1vFqk1fwXJ
zKaUsdahg4C4KpkjyvfhXrAThcBKsqfV5Ie80CNNhBvCjwgsjTursHgGQuU+
VBJSxX6vuS9S+nlEwl9BH8eNb7qNfVhSicZNuK49iS9X9dNkQxnsSxYO61kG
Cpl1V6o7nv9dF523xSUcr58mjU/ByKDGBiG7ywdiLpIPiGItF6l729ReCYKo
2l0IuncdExHxVPRYQCeVwpaqtETjIjByzaVCorycDpYPtqipySKQ44rHNYwU
x/CepDHqyKy3x4fBA0KJnN5QMwEP3wR6Js11gcLzgaVIS/0IyyWF7X++FXMx
ScnxVEMu8HjBj5QmqFOL4A2sZWeS39+wjXc27nw2LhEPP/PAQP36BCqDY1iV
UphnAabvVut5oxlD46EWq4XPvuGAntODSdIuKH2D8/DERQVC/R5imyrhk5Ty
uINKOBgPCw/7WJ45CVp/qcpkw+7HU0v9EApQT6rZA6hDjWIUuCLUhV5D7ewG
Z+sbMdWT5fSbo9xgPeYiQgRhiK7DEm9yAd4r9fuWnpLLl4gE7hKe7qJAlKhe
GNZ7qwu+6OZbrV0EUwhHDiySU7RwC8ouogfrzwZ8sth9o3Lsp0xHqtVabx8K
xvkr0heIEeJhRWNYVLUzG7EXz9ZtCPW1tuKZIOkEEQoqi85z6zOu4EHvYY/L
ByNmGZL5kuwemsvSYRnUl2nM+DF1LGvHgoAu4pYMH1Tuc80OTGogmbHL9/f6
xuxOxYzWOiityDyYsk95JB5SJkdVdRlln8y1echE3UHF7NI11hBBmr+tIxzt
9jZqFyOMmANmESNXekkk8p5VmWb3FTuBUmvP7maPhW6JJmWb+Ojc24HmNmZD
WJqL4mZjEKX9ujaWLT2OuUyDb+bjMamRspVte9JKrnLeAKt5wYOsE2stFI2m
7WPGJx21TM+b57HII2/+dar2m9TVugeQhtv4u3ynD+B7sCPGDlv1b6lu+tc8
BAWDyWAx+XzF8I8czhPcr+AkqtCXVPULv15ckzXzPyqkzSNZ4b4E+Jf7QIQ+
cc/pJ6YYP1wRPvFdSAjkYy4DWigjBjhebNkUZ2DFFNRngK106xhsE2Wjutkr
APM3uI3mH3UIzUAt7E8S8FVShbWArJGUZa+R7+BK8Oof5lCgyIj+bpg1tJwl
kGQORxknQb1N0QmilEt+eEKkfp8Ma9gtGa7EOzNKcKwEK1dRC27el/mJbHq3
7O320VEK8d+glra1DENgGt8dLjGynxy8y6T1l7r1ykVAvWkTLRUE4LxA6tuq
yFpugkX0wekHMJ0H7we6Qtur1tVptqwLxN374PctNJtB2Mk/iqGzPsIS0zdu
PptGmkaSP9jF8dX2azQhNHeKJrYhyTJf7bFb4i/9GhQHtcrA5zyOYwj8VzQt
NrbBiQ0T7He7kjQXppRkDErFIP5K9lSIVafQ0xER5sVShHfQ+XIgcqXezoj/
Mnp/eY4VZJh/uVWo3Q7w/u+mZqCYDhJHDVs0T/FEOFHVWwbUwxC/cF7b6XBf
6plxXj9giSV82W7rwICKA8rJ/hpii08vY1M9e/PCOI1hu/9+wQ3CRnpvHra/
tPv5oXExRRrYSaB32QI2gBWzWe7qF/YSB/H6yxdxLFI4qA4TzDKxSSfDHwHh
rYOd5sBzjzNEtaNRs0HsH/ngiaVw7UqjYPcE/qnb3EICY/NUEGfstxyGfN3w
5qPVVuJOypTxkZJWrg4IoT2r+u9BHGqtHJ9afLE335Wb/Mb5ugVD+huG8KqB
80vF5WWSFuA6vaFEehRU9NwBKRdm4kDCSjwjQ6kTNBgw6mPf2NM8I4g8KQ2D
yzy5eNQ4Kd8I49OHypmaHzyX1xOoWNoJuKB2SAkMKFYpW0sN6jE8TsEbJ2Rj
1GDHI1vLwp24hkzDLtPTOwCK8KeLqeYasPMQkPJUYOedqUcRk6qYGMDhhGjb
vGm5hZLk5LTsVg1v9B+pYLLbXejVyk5JJhbg4Wc0PtreXUwAzxry9/s62Hyl
e1jEJVraR9Cpy2rEeKJHCQybzxrgJhamf+7zYZZvII+Vmo1uQQicdoMa3ysQ
OijhYNdrwmBdBSkyarm1SEimot5NMbPZyS+XujiuQVGCP/lXTGoc1fv7XSG7
RyRdP5fLBVgth9E8x81xJGMHvNKcR7aW79m01auDxE1yuRDsn7CiC7rAHNhG
3fUnNNUzw00Hqe633EwEBduMk81d78fUR/hnUL01rHPzXagbKUGKs8SmDk0v
UJ/ZjgJMIi6WQnx2Rmei7M3gLp9pHye9SeCWX8ehyZrQq0veKEsr3yvex+2V
m10jPCGZPVjlGDJaGs/DPnPJ9bP+g6ri15Y/IGKFnmvCsTXAvovOjc315sFn
5E7b3x+jgWr9lwqOyrAK2Mt0bGQkWyQFegg21VsPZpbt11uTTDnZewnx3AZQ
MC3P9D9BLO5PaaGoz4VCFA63q5a2qN+6zR5smAAHv2VGAyBdLvhEEyzfnRSm
MQjyZV5aXFnL+/CRe5M2AV3d/8LYnKTc09sGQ8Iw8LCc+HD/bHcQ7nwRxWrd
ST0I26Y/l+yYUz5FGBoakLUaOtRW6uh64qkPPSQj41nU7EU98KKPNmF/pNAL
JXqaOWrDuQFuk42HLlOfgXLvWtiMUjcjd7ukfv0MKLUF0gAheDzPVD1FNkwT
KQ9OWaq35SUaB6WnG3qmEoUhSlrs2g4d1a+DNJrReYXMEGz6+NC/6lpyTDeB
iIoO54i9pgY9yzOJkAwVYYjh6VT/h6OHDUDeo3mjPW4i3XgxE7UD64wjtxcJ
cjEGgOQgToHFVZ+ON9rVGsCy0/LHP1iqrkm/atZrPRzzOkj5JXqLr7piVHe/
FG7lpDoS78VzO4+xXu2+ae/DUNZGWnbJi/IbTkLGrQy3teV3l0HktBD0Znyf
QUJuHRFJcBW5QXHC+rTE53YomNeHWvmPb6g20f+ZpWpNROK3hiBtILt7QqN5
DmMLOWyXM1Q+oOZiuPkUtWR0Yv2MaGdwrW1sf5CVuTwNOstb5Cxs/OGC3sPC
hLXPAQzd0vC6vgBI3TQgQOySMZS4HiF/8ZMZEbeJZEcVp6U6nNS+Kc4iEwYD
mmIe5WkMNjLbjlAuWDr427ZD+Rqn0fgxQ49T4jj7qnZLkjzOK6GA57KRiS1b
6wxAmKoZZSJg09SqVkP+WIppyi7dYUZ1yUo2vY7Wy/YPvI2EEErvU9oMbUN3
XaEC2ysX2yIHItn83guPJnMKnS0PvV8bmBv1ExJTUZhO6aJQQFw6ZL6OnEgn
alpmSiNMIBTmlb1LX4Uzheb06U1RnLv3KxDFPKxT8XdLhSFZUa9iujs1ZCka
1mjY46v/V+4cQmuDgOhL2cjE5SFVebFGTInEtRrpoJ1i+ZX+iPSX8RVkUSbo
8vR9UwPGzsksf8wBGYekVxAslhsNtEP3RXB2Nb935O2kdjoKJicBomqpqLPn
kG7niC2iyijwmMLgeo68T+YP/fkOeuB86+sRI3OIe3tp3jccahkonmSypqCj
n0NFPDYzaeJ+UUavpC8HI2tY9sJ+RVP5h4CBNpWGFwJkyo0jTyTB0JBOlZFF
0zwp00m0NSa50dxa/6JsYd7qG6ux4GiZ3xR75EAJ3uFcmJjcpVRVTVJiKYzb
xNZ3bMRZuoaon0wkgJ95MGRxkkJKgEwGPIoww+5VH+eGeTa+Cykn4TDVHj2g
BeD76C7Ta5QooC8uJomJMBuwAKdQ+YuE+qxa0Ql6lDblgIANJDwVfJRbm2Kb
TrAIx1CagOQBXLCooXJl2b4tO6aYTrEz0g/I7owLqY+d4UVRAP4rVi56zS6G
qC8MlRQJ05D6DEydmE0NVQBAeKXRegEqecdVLDBDf3sM2z8ubbmLrZwHqqiO
tLtX1rUpDPHMvjxNtWsA0If2BA5wmMXc0ONLftvgiu/4iPIf913xeWUeP3Ve
2kN2pHfjqNaBk85PPU2scmtgbymTfM3dPXr1WbwRtaSYUQLq21Y8X6pIhAxz
Z/uzcbTU0pukyuulMpim4QwHZb8Ylx/PpZZ6sUKkTUXjHPU4A0lA3LO9b9f2
Zm6/GF3wOaqTwhYL/SpYiJjJNjtKFIx/cNE83feFU9KQp8O/yEy9ZlGdgBfC
fEZDje6Tc2MZCHALuwg9GyWBYDHkt2BGK+UGeGlFtqPCokJLnZhhG9SuBfA2
l+OaedJ1EvHmURyv8tNsbJJxAWAlCfCZCP7RA+MjE5gChHwFhw+1QkjF5TJW
DOcZkdEZrhijO2O3a4uXzqd4YLcHVkQQfdnvYDDAIYp2Z5s4FTeH1aW/VOg6
3hxG1GUoPuFtev9dlYIheTDFl8pnyVnqxgKnTbVKZRRHpmgAdP7WDzo79rN6
EEnoSx2hdsIgJhIf+iT8wZ15tNH1BgHaWFZnAOGmYNuTTl3a4SFPrcFQEkXF
IvIWGaHjGjq0l6AvbXp5fC2IG92fnevmFYDfUkxFLbYUzFbQ1k3gwVts1mFk
lDNXYtrSi/Lgqj1FZzzMScdcHszmM+eYn2hZOIUCu2r1txP7esZ5yKAb3nBS
YFxoTIOFJVR1f1f/6x/lYe9nDMqZJtMt8KmjilEmh04VV6t8vP24/owG+A+U
FJASQPMhu7PdSbgaIOLPyjrViY/Kbs4h2v7dt5c5bg46qIvB2QcIsjBTdeW5
/ML4WLg2QgDjaj43lyvbjerTEezYl/Be6ScGSV4+g/2rIALla4TZaABXkkKw
3pZ0AjtGbGEvA0hgUF+HxTXd6mgGyzAslQdkeUoiiz7c10xdiGHuu1m1H1Jh
MZlkNlIf1t9eVC2hgbBp4N+weEiprBgGMpgdWITeJqHT1XYAMn82eyA40Lcb
K2rGSM86hisn/uad4ps/7Q7vwfF1sdQMKwAdJkbSPg+olTgelq0EUmQLFksm
Cv8Cbpl7B7YHUUoarBRaBTNdAAlPVI9WNmN/yhHJFgROCJF9p4jG2n+VFvbf
+1zxHP/v8xB4h2Kv0B/HgaQSMgBiCsV6ZSlzFK8ntlYSyy3eTooisTcUHKUY
1p/MPHDrOfV0I3BUkXsgmlN3EE+v3pHljgC+z+fyR83PVGlzQ4bRHVxbQY2/
sUe+s+dMPfQNPrLIFj3Hbt/xKWaZ5hl70SBcGIliZwqwC0tLqNfcUXs1LZOe
oBXDNoc9szAXoHtqHnyPHn2/5Ch9lZf3lN2ghHFAgGXWwcwS27UpHIYtEPW3
G3KbjbftBDVnHa98G/C5KQeyLNrLoMsqRoUboS45oUE0BGsGXyUGbFxN5BX3
ushTcKHrxsIxicLR5ZcvmFIR3ZekPlxqbrSb4+zJnM/KI3/gzZEnLmSNhDkC
UyZsK4nx5uvObrbhJtM40s5yGIiTJ35Uvi830pKnFcvK5Q+MaeRgh8QOWNag
cW0gY6JXwd5rlNLlB5pY8EmpRu6e9IyN7o+SUsodh7nu5wGFfYr0oKkizTak
9x9prQBmjFiwuuTCG3Izbn/re1vCL1qCTe2NzrYtSKgUtcEtieMsCfhNCadR
009HvnN4f1RBI64N0ArvsTWDXlJ/yV3MBzvHlzIxUUVHl0mx7mxKld49wZmU
HU6B4HkqkcMnkbnIRTtccPu7KFt3Jco3To6NZE7rA2JZ4YW9po/U9ON/YFov
5hL70NsC1o9VEfaJRfrw+A6TRoUwzLWjhFvsb+SbK7smsKRvWtzhKdYtTuS0
P5CTFdD2+dWPzd5pPaYGbNDG4PGHtmKVTyTHYB+yQfosWsvqRFvMXET0VXgf
UsW4jr3grE85BDi5PYxlzG7XbVA0C+EWPymc2haAhsjAfrwXLDQ1Mhc/ppak
iodgY5y0FqM2BWG00rkvMtKrNjOnXqzj8nO9k474GjYZRxIyo9CXAVxpPHX9
5m1u5xFBmGCbTSR6KSwMTxRb+4k9IQI7JYajOlR5R+cGBt3hRCAvjBu3GMqI
cPi7EmKgPYEkJ29nlXUicbEksq5Vh3wBEVTfF1D2eQobP44W77CujKn3vN5L
5zx5JpCwaCbs1ZuZm1RwzJGXMTNODpYgssfEfR1J0sYXGlNN0gpkHGAp2nZa
u4QITvrx8+GgOhWqULjsaBFkTvgj4QlRyZY+nHdCBjspE8m3mk+Be6o+rywS
2JZwMmRlEiCYs4xqRXyoPStaQKamZb3sOoPKuPatd498oXEN3JLqpOwUxBdX
hRt7+C8SslgKfLPzTUaqNmQ+hSwZP+XhnM0xTVvioVtiCTY7Hf4SjvzDXJba
4SVUDWF1YKmWk29qBUPl0E85yUR9O/ailGHM5JYRYzVvyLubHV2fFWnGXpnd
/TB2YpjOkHtoHmFyiF+LH4wcICODpO5CKbzCtA2tvUVlAdqj8KYxnZBn/wCd
uQY5zdbA4jg/I+qz4szd3k3kTrkZ9l3qlnbIGgOObVcuZ5x7DIMchMvr5gSo
NghCiq0Ezc/Y8X+YlRzsvMb+q21jsP4OS4EN7R6Qf3v3pF3PMF+RNTkojxlL
zZakdOXPp5zzzK0XSIqwcHuOVwr3Ys7pot2Acn//tPFJpRvRpccw1HgWYRvv
nAhahMXFFMY5hhXSvwHysWkCmTO03DBzAPhkj36ZX4ZfMpwQGTICie4g4fh3
eK5AKCxTJExM+Ci+5SY2tWr4CoiJenssGK0BFAwGIjD8LA2ZEBQQDbJ7ADJT
w0hwcF9doqQrHU/LQ28oROX/9l7nuGqUOVMa+RV1ak0C5Ntw7y44SPnMEqLq
1DuN/whTBGrnNCkQvGQi5vIFaCt+5ZzfDtnqXHViscOX1BYHH+JsRW8XrfKv
R1giVeV5NMho7tQMkWNIEETjC8ndEURjwEYZXyhj3E4y3q9egXjczPi5tZcZ
+6Be6IEfpHn+r6G/q7Xsnvn6gRG10+ohDcuBXU7DR3y+2WFJ/NUz5MK67BzO
zsyt5x/MMMKrip1I9iLVNOaI3zM4rYxdBHDYL2V+JYjtBV1Intt2nwYxBVNx
BWyFMFaEqGQf6sr2+G/D1GzG5+zxCJ94bzM0g2DDpPxhv4pOO00Y+vahXuEb
gNm67f1E4pIuAnLfJLihhO7GnSAdVvzyNqDB7zWdfP7KArMZMyhekUoz6CyZ
vcNbf/baagQqhd39+bgkBq90Mpl6CSRN5VBfCUNdUpzBlGW5LXLS+fuDWuJQ
RPT/Q3vjX7PHwJla3Ztu9ZNI2DfD/KLjx8STmjckJlThZeeT5xRKa2D280Uk
yDKKSpv/4X6Q3wn/+Jix8mwqwiICTmyINUEjrT5CWo/8TIINGm+xkM1wOLVi
aPhD2M8acIKxWJ6VAaFJQQvQX5OCVgjpeZxW3keOSSgvOQoVZgBIQk8QrGCZ
uzQYGzHbwbgQJN84S+uKUgG8NCd0LOMoR7WpqE1vf8zzqHae3JkkkblHm27W
19q3GJMVSWxuyQADs5eFcAWsc2OYoNNeuZPteSBPannGj+26DkKBIVQgbq82
FnNhUybMZ27RVVV1Lep6mOoJs5BJpSUs+wcbI1HNBSlHXZ9AX37BDbez1YAK
j759YIt9duXyvLZj4orpDZpA8213SvVAzUatNx6YNkulWdebuVuth9IOX9C6
YhqMddggkj0o025OWqSI1d1VXyGiaCxzFMontezTiUvojB7Ss0aL1Srl/sUM
bh0SvzjyIMzH0uxyZ/mrg/gJ9L4Ji+YJ5YqpjCVHQ0C0oW4RYnoACHXT5jLy
WMqYbr/OlHFqAgSgtIoTU/mcr1u6L52yH5qS6PRo5R4VMyqHGxys1DQwxTuE
MEYssXavZNYiesO7lVbUIUke3aDNrEYEaxvz29ZSxohLmMqZGhHziY78S7SI
xeUrKdofXISfBoaKR7pR4nkbl/tmaS89ca4OajmqVIv/TjMJgqVfhgmgDSpa
cUeJKXgFyEZ8YE+MyKoDrNCuN4GNm5xzRHrJH6Oc+WRah0F+K0l0gLY9imqX
UJH1EYDbygs8MfmtgSqj74BGv6QrIbg8mQMmqFlKyvW8slwRdTOkwouTErKr
atRN8yYSXV05vOBxlqMsUMBhLIupiT0jVPU3l+hDb26cYLrvSnEFVW4jg0Kp
WaY4fuBPUlc1+JTFEOUMv+th1/XFs7issezu0ipwiPUYKFOjs/cojDiNLCKv
hO/L6ChOgtfBiA5heiU7wXUsXxbeAkuVHolWA8OptlOBnZZaefl1tmXgljQb
2+c8QBNRxh5jwf0jeUDb8ktZ0Ug6eqFGEDUuYGO0loY7oLh0eexyyvfL7iVT
JMaKhY+iiGz2uL+76wFeYYDM9LYMGuoyXnoBFwJWVNXxTEw56YCv5Rgi2JhB
NfN2A7BEcRrNBiYxPZujTJ0tlpPlS+yZC3DTuKMpaSXaYluiAoQ4K467JyVI
12vR8X92mLoIVQFDq8mIafnywk/JHSlX9dpYwoU6fxfGgxndfo6JbDmqMHTe
LitNaINz/CasvDoHJ3WplXXgjuxITMR2WBzyUnx1m7agigz8EQqCPRHQdbRy
j51JumICfthE5A43il93Y3iBaHQP4+pXSZz902TtDjnqAzXJG77jQL5JWLOD
4uHOKwG2yBvcaDO0UTMtfSg8AYKkBMaVzHPer6Q/Sdus3NTCMIo+7kFOzy8f
OdVo+JdUlDHDMQG8TwwWoxy1aic1H6RF+sN/mrM/EkvHGRvu2ns6nSda/kEU
stwtWXTEss933hGDfqTrXK8rq60kYGL9eEdUmrzTKLpZJ3otfnkDver/+LLw
AV+0+wDNQatv6n4aD83uXvAK9/4ceknotU0LXJDu9YAhWUItNMZyNoLzrCCv
y7uTzKrGZRrlJkRyLVNpXo9KQlErza5AGI6KvrV7ayEdOQsUzomxim4d+PF3
KBksJPz+LHIei4yyRjkfMN+9cPBpJvRjJOLIWoXeKuGxQpMSlrUk7giPuZp1
aqNcEjIK/h24rhE79YmXXdGh7/fHLxBWETB2XjTYktks7hpMAJT+0FCydjsk
8BWLEzpxYSRLWh67CGmo23KxRI0ofpec5FJPcKHryuia12gJSQydKRwS5I1j
RPfpnuNGIM9ccrR2PNEOcO5MWmFGFwlLinr30U3Do0H8yuvHAlqvQGe/swsi
xeWcVE8U5oZom/RB+3y/kCVhLLD8mw/vyNQ0uytUOSGLT2MyQSTvrt819m8B
FwqzsYc7KtDeBpLyzQ89FDI2oPjv2OcthfEzoE/oWQmff+TM2ainC0hX0cA3
QnYEDRP1pbrKCXFu3I/6ICCzIX2UFfRqjXNqE3FTBBtkzKrP54QG/cBSE7Mv
A/3Dh4FTJe7Qn1XXaxURDKih/1BTNlz8THMQCPLPl+S/58FJTl2FFvDub9nA
ovEdU3aQLDZ41NlYbmTbr8qHu477W88Ap3yN0nioLqu/8n1wlIG6uOe364a9
NG2j6fEDM50EgK8gxCf7P5Z8hG41o+WA1MsFxyHRh25RcLbYQvN/tmOqXSpw
IpWdNBT4DVx4jhNAgE4/4GCKOVdoIu3ynd9NPVj8sEbvSGcofZv5q9KQrxQH
6wqV0oVMGFdc6BOY1mQTSSkOz+eiLHfzwLIMxyHRHi6QDJwTlhKLhZvZHVcn
btNeX7J/nr15lfrnDQ37L0ogDLk65V+XeKvxYLyU9EOS4ORArQ/QMuo1equn
w3vBKqtWppDTJt/HpMfSoO4odNaer0G/9Ll1Er3hu7KnPNp/mGamDr6N2y3W
w4b4INLyo78pgVG930cYPG02qrPjkO4ZN7Gkng21/5wjAZzzbZUve7dCGXZ9
XMrPb4bm9XZBzCVoo+vZGvM3pWK0fZtCFwkTdBcrYGOuCX3LBafqDxkYs91M
j08Z5ZKikowiwXcgVDIUxg+DnFhbUX94yerTCxoDM1r4q2fUzqWJO1qWB9J4
w79dXUTCcIS3oN6ia6gTECu26KE4WdS7wp2Wv2TLCfVxHKvDpwt0Fx2RxppL
3//+iE8NX3+LX1K67WMFCQhT2oGWlPuDX38eUCCMukhbVl0rFfjVBnALxo5o
H6nP9kfUdFERfmsdwXusSQu6QIu//GJAdpbXFpzXhGpKcqguV+zHjF+Dag4X
gAUcX2LglZ3Uq9Kb/QwCki/A8RkzdEZ2soMx9F0sJMJdVLMRr/xIqr2kbxAv
ti94s9j9pPw5uIkapUb6RtNRTEgEd+cAwKmJkGXdW8StStKcgGmqHJH6rcvU
RxESuM94+tsElW/wIKw7AjPYar0iQAv2B1G3TKK4n0eEOEyZUZGWXAWcIaAF
4/vrNJOZ598rjZJM8S+Qa8H/1I/GWHAgmjHSGG5JuHbb4ECxNYr3qQ5GHjn5
5+2DP6rTp1BAVQOqqjAU60r7dIV65M8T4jjb9iGC7p+ks3eN3LFGLea6xxfQ
/tDC8m4TC8KRmoQ35ZoavxKkuZxWNZGKSmVEYIJ41l+3qmoJOecFLc4lUy63
XZBXJ0992X4/QnFgsZ5iRUlbe2B7IO0yC0M5kcfg9rJ3S2tbDvr+N6xrl0xc
W/1kDmms2u9fyS+u2KZoDUyCNTVSixzmZMVaQPvY1wYoGoRR4weIq4O3u5Wp
+NCG6U6v+t8CdQx0wFATsGY6sHFhy41Yw68Wr6c0/s+34BY2HAE6Uh4Lrl9f
xkaiKBdj9/welo7mY0SZp19NB41ZmwatZ/nFfJnWDIIVfileqURvFNB0g4Be
HKeOQEL5SkYuQh/zmG9mhlMNMliV9C2JtMLnr37wksSzckiPg10rKzLWRBDd
5tx7eu+FHpVonKRmf9BytPTUSiVwBYU/QPbrErDWBSc/dkJjx0bdEmCTRY0K
QbhyD8p1Q3V8c6VeUSd3qsTZaRrP8AU82jNT74+XZLFKSsyW9/mwTwDsZuMb
CFQuqBmpE7/tErRVtzbiM5WTYv1TMEsvTSf700No5WIpEFtNXcHLz+AIzI8u
oJ61gT7QDdVaBxsSY40muuMwOcv9zmFypDLPZUrUkWTpa/gwpu9rvuP5/6Xj
MIifABsI8XBVsldlnKmVIAnhOFcypMuOj/5ZUBZ4wDNrsY7jPrJtU3wuVtM7
3jGnPs5Iq25LLmI/qIPhNTywFUgQd+JgM0EwB5/sq8zKMxhv0NRv6j1lch9S
XYrrhoBpVjRs2Lsf2THnkSlojb9CLRTCC22CkJV3QAMXKSWaW0KST8PYNWxE
GUsc8ljVQFMrKpxhXlStO6HYgxUNiWrAXH0WUqyOifVSi55xKw1ZIXYPzkSD
9ecVYvpqSmVVorIFicBlTijEGPaYfYC1kXJldppFyrhRC5I7Np/UmEXlPDzn
fNKzoN/nDbitCi53fzBBTGWUePnpHSb+Spn/geNN04mfGIS3RdaDwb/xxFOs
D3o9oY4WkAJRLvPBneLNVjxm1wH8m9kXCujFduWMxh5xlkiEsVvye1LgLngR
tSaWonydl6KMy4dmkY4ICf+ffpWo4hFEEymwlOVjql3Y6Z0pPMD6PBJozkE+
SdF2qgsSG+BfX7BecPcJSg6MVWK3pJrsKHo47loxentxFvhzL70IOsOhPOuP
yXUaUsTDSOwMPFi0Sc9t2ViNPNcjnKzyK9hk06UMDBPWOvQ4PBBIYUUzEs+k
Ae6uwFAiocQQrdyjccYp+SzjeyRuXfPCn/Yo6264msg79ctm+HSiYZMS/TsH
HFv4WbC2AK9xGLQK9tZy4z2FFZUcz2cG7BdNElaTWArd6phQkrrwmePocZB7
3YnHxhy63uxRQefB1xAPN6NajxExRy4fVlAkxnIjOwejQiXz40LCTO4dkQLs
O77+6Wix2dJIpQGhOqAWOvA8faUtMyhT2g7xfsH0KNMpVe84xh0FXvTYkehD
W661WGL4MSJIRduIBMrTH1s9gOZaj9ZbMtxa2bHFPaQ9Ojvff0+VApkdkCqY
nIWMajLmq8gcs6uXFtVAs7h8RD8RO4Hn+CAcOwMhBy7m9s3NwaN7EpiWreh9
1OlFweJgvGSSNuYREY+JsF5Bj9HAoo8aiUTrU3ZGupoMxTjlPzKO+KAd6gNL
mCT1HIDpEUcaFUxXiNW7xg47ErTcNuyys3QlKkBq/yE4oqNZTOLK2zHjN58h
65nZrSgvVBEsKNAR+o0xWoaqp2r8+K7i98t/nxsyKjs77hoGvjQedMkKYnVw
it/Gd4cn71KmWmmeYtgJ6A70uwl3ay2McOzfmlEBx7Qhodd/SlGrQn2fkfI5
a/3KTNHhS2cn/J8000+iR8KcsG3ArZ0JV0K/7uZfDgpU8sc4S1MnsfjsyNMB
jH3OLC6wT3XubcufBAcMq292QIG7+sISAOieiQwsN884pDTxb2b1vqdLVJSP
rY6m9ZbthpnLNtq9VsDW3yTRNjwyboxoG0EH/pA9FWGjdM374/JrB7lgOBYf
P9zLC46jwAowbYt7h5DRTDFeJvjHX82q9vqusYEM4UPbiYr0Myp/6WHd5VTR
JP4DmPxo++SQtYovnMW2qR2FB+hepy3qEsBIcFeD47h8Ky1vg0PiP6OZM+tO
hsBGB1adtKSgWhhvlb/Sj3wEA/gOw8WhMn07SSTU4/2d55gFNOYvZ0AL11fS
Z4d4J/nTcvVTdUMwfNbtdnLaigfx9GXDVF5mjrNoTiBKLjT1N+Ww1kDHo+5V
4x+mxfAT4xCgtAhqOKQZC5Ab8YP+EEVoSsBHiB48uxUq2gcATe495wQCE+R2
C76x5eMiHcMIF5iFR/1C6wnAAKJQBD+kyS5VDWuz2PKY2uXp5jBqAMM3gnyu
f+IIC5Bg8zvrkhVvRXWftOLXUZhAJB2qNKNisfb0r0AIqPMh5K07EtZfdH94
tg9CUYrptPJjiZ2VE8od7Bo+hPpYPpB+o4N0UF8eLm19K4dFyu5hsOF+6PXJ
83AoyHXrz0kiIFsF/bLj8yf5e2JAE0eMMulWupoCI6UiJHrb/ePO3abLab8e
1bURQJawBc2C/GV48goxnhm24bMbrhrbW/a/dd0y6fuuGLiGoLE3vwRh1C61
OI1QpntXSzLKXD8SZ8cAtGHLO+VhnkSH5mr3xKv8/aNgGhqunFYzkmInh9KY
kBKr4Rx3IJob+mGv759qmM1AE9c/e0d3N8DOsMkOjoa1b8dPm1PNV1s/1wuN
cuaqqxWFOnXVBuWzmdlqWO935wNcqeVRwzpB/AS9NZnWMeKY6erY2Q6+3pqs
yjaP2VtvGzzB0dZxB9x+W3JNKgy4SxiLLzArjgtZH5nqPFx+1WWj6UcRaPCc
wkaT63KDhIvorNwy9qYWCxSJixP1YceNH0qIyfTFzNyQ5Ez6kDs3ozUOlcmr
pBRK7XnDFrzFktAfsX77Y9IXAKaimDyBVPemYMiyL/QPVk4G3UN9JVGsPNG7
LwlpK2HmDheDQ0DmCvPh4QdcGHQ3aOQ+jYUapyH3bU8EDfBolWg1p7dKbp2g
P78SO2ktQzNQ20CQAoxqDOuyVVzs//UUX8jh89ey6sPQumCs7ZVdSNTtkc+D
5ampT2e2h1/wrWjWcB5cpwqFXdqoRxpkScZR6Y4yYqFDHYQkLugx8OGABGAR
+5ZmQJRUMA7pJGRjaDCkNNG+HbSDUtJUltGqVzHxPtvwt3AZp1HrqpHBgEZM
H7CjBFu70JhgDLMrMhNtqQJrTXdNeDmnZPBPxyBoNWbu6zeYVcZsPvMlTYh6
lpWVYN8gPwKdW/PHVGr+/FuY3XUEijF/tBpkfYINuLbCo8h+cI4EmdmLmiNf
yMH4pKxnH6LjE19lYS7RsYrgjvigxRSy/dL2fPHzNMC2UoHtlEgaPCEPWJB5
2OLc0MO3ITw7sanOtNR5gOvwDuBQrroeg5hhDZNEYBQCPK/4pkFCXvx0vPYu
dw12dlRj0WObSJCIZhTwu/sL4D2CVdj4c9u35DXoGK3xXY5FzowcO53j7Rka
yKYOS4OJwwPh12LGUStt+C86dvxCVzlZ6gRcfXw/9evoDeYXMZp2fe4vIKVN
vRDvpMQuXoV4fQqTrcs/kHWTFUsJp98OSg9E0cQhqCorM5uUDhLwnBGgK5mG
G1NneMsrtd8WF5KdLtPv5smbDAMSmp3F+xybQzDyGFI7ZoRSMYzmko/eVsXT
WXzmuDQvSB2OMjNJHDRppkS/B+5lA6EMkOplPn5X/bt5L1KHJSo8zN36ZBHm
ugW4+TCt/19WM0ClhuBZh9dP9IFCX6N7dmWfJ20OvpW/KSe7S/gWqWHhryox
nFUYraklDkd3rrXd1hYdT4Nrj+DtQrYd+O6zMDQ2vU4LwtqezWz9O+HQc5OX
imjFF1PBLz31g0qfzN3xkwiFRO5AkQQvjYfRQFfUp79jPShFqHq2hCeVnNKM
cF88duyyqW6cFtowBzuY20H2wEg7Lv+riB7TK9kHpjtVQ/dhFzX2IFnkLJyT
HiHqRVJU+RuP8CRaDqQq4CtadkZZ0n7iVGu2px1imf6nQ/olHK+MChyuUjZq
RaxJkZGdFhZxH/c+8cJhqganQNv9cSRwisFXN9BRQzqfY672AKgjAxdzNUnu
V4C6sp9fCcAXSzN5bBxC4M+m9Pjd++ftncSadk1GJjZ6/TZs5H2o5D7xgat9
SIL4mV9fOphD2BIxRHcaJ74gDmdPj4AqtNojyUjeZFjDn7opGkNui3xoxhh1
qYd0h2IxH7Cf0LwwRGCL1NtfQMo2hEGqefcOa4GoOQbHFQaxe0bTGvckY+Rg
06gI2jBtNIFCmOFChSjASk1kGLlNMn+iENwrqGx2o3FzbSiM9GkDKVNLBnNd
m0mqxeVIlwA4KkdLBXh6YUpJJI16T92XeyD155wfhRnpPZioVrD8C4V7F/AP
tjZDtjf55z3tBBwWmtMTb0U8D6D2zAz61+2lf0kGKcjVQ0HB1/UEYSXCH/cW
N5sqGAdUWkzW1lQIzEOnvVYr9ZtfjWi/Yjwgn2nv0wkRh0GkCTH9mTRprETY
PReR/B3y6FdDQ367Ho0fSTIjVUakzs3C3iKL3RNuBDdmikO7qgdTnMO7GiTg
xHrSb3obSxIXM6VUQqSlQL6JrXOSGb5J7E/YFMmX2QGA7N5rOoUebdSPGNay
c3zSnglVsusliL3VY5zNJAjR4Jb37OS9SJgfstZYVruZRJFiIasZ/SwnkFro
U06abJjdLo4GvVevXUq4+lf2VqhLal5t92LjnMbtkGNnwlIk1ZRFSSjnXJYy
fxceTpsPBcL4x0PTu8I4DSCRW95miAbq140fFAFLAtagrK+nQldpZqzpOjQw
BpQbLtVrGBhtgHU6mf29xDZjM2DudLSVDVsyDejnY5BrGPFwK+jjCYLaKkci
U+4tvA2NzyDu/5rvpufsAHiEDeJUj5zoysvZJeeBnrLzLOVad9YhXgoQQggl
sunJN5Dk/eRbyy0vjWNUnXShbedYk6p6oV0wIj/SxybP5kPsk16aeyjzgRuL
VlPzT35Pq8xz3xnJn3rWGN5cTOJ++phN13aTiB3ULeV/ccDvXu4DRpsKC1lh
mrZSBO5qpDLBmB/9ELI+AiqJBEIj+8p5/hlg8b4d6l4wTYX3Lcv0wFAIGhdn
ny9wfcmiuCTK/NAK65bTV+/6swKjMXN1MF3Z4JL8dYkO0s1OqngFHF5vsy6/
3A1vnW+/Up8BNVLfpNuahmBtlBiBZkkcaXPeW5Sdch+FpwkwdQtZgjAVisWo
tGKZfLsCGF15GGDv4vb0slVNcQpLilypE6uMZdFCldV5vhTqYQnw1aDbqkON
pA374WK5hbcSW0G1FoN/03iryLwOyv2RNjmuviggpXDAS4ATVn5bcV6A542C
TyPtEDEyVdg42dk1Z47io09EJTO+Dwy0QXNVp7hjRIddJwY6myiynU6Qqed/
fkpglzFnq04aK+CXB5K0A6iZ7vPu9CDIygy9wDEgbeYSjGWi+watz40oCbpg
JRDgRr5kyy4YSvYJuev1zAGYDBGkbihQ7DaLIH0yXvBJ9k+xcsfjUNeOuPt6
fg+58dyo/IQCFjYpD5zg6rX5YXelhz3c276oMkM2riRxehz+izmzxAwQDSLR
Walm+GaYVTs1DkYOl6PvlBEl0GKK6FQtRYyyMaj3MN6JD68L6q4ne8xi/cJ0
UOMIYfi8WcPGHH+3rw8Bs7snD2sWMA5ZcHzFn/FvrJH8pdU8Ti6zHzXqS58O
lLQn07OOT/MAjg4I+joLqO+IoLV5OMqR4FgY/zPGvy+5pfGtkT13/tjar/VM
jYcrv7aB1KkjbiuSccQU14ayLxci/o7WjT4JIaiBBnf4PRUkwEMraBoV5RiT
+MhR13+n4a5b0nVnm4NgBbll6nwm73kWxlECjwxoZC3KDHsZNbE+z/Nixpfj
6D+pU62unU21ROeueDywaDxQVl70cr+xZu1JpaZRTmktzckdKqCle8GmUmUv
RQ9fRXRqYxyEfpVwmEHJxk/GANiEXYZc05ZihmiUPFFSuvsMBGpaMVJDXwsJ
g07rVfkKCeNo3eD047DCCK8s6ta+sONjI5THan/xGp0CTvA2Tm/2hx7Gt4Cj
82fcqOWS4RDvzeWFqHmRW2Q6HfgTdCrcbAW3F5QMOoAG/GG4cD9yot6Ctt/x
8A0z69G+lDfZM7PZRUjMWfIbrixsDWKcnsUsObUfiAyTMxN++2GVCSmBRWPH
yhfakk1/pS9Z3YH58cRlKBb8CJRU+bDpGC38sd0+sOzWKJ7t/KRZQ3Hdf7pV
JfdhQ/w+axepOQO4TDbpAGzamaOpZxjvn9NfIeMT/q+X2PmeAAUNtFs33f7a
srOxBN3Zgq4kg65M0Q90/W8L94/vZw+plRXgwi5x2uScCGXsm7RsO3nFfSwz
qoqJUHqv3QQcSmGBdB78amKoUsgufZHlxB3REDMSisUwNHhz8HJoI3eRj7ja
yPsBtLXA+ALmlCi9f9X0zuXF4Jkspeatoijp+jfTQiCZRhxImbGZN6eZsl1W
Tg/qz53oVd+H+V2oY2P9pX65hXs46KqWCZWqwYv/8isBb9ubm8WpivM8M03c
xw1CKlhGpIfG+z0hWDPpio96Zn7k9EqUkCvJk1M3wjs38AshD20Bj1ijqz81
dmbfydqLIzrioJVefMjb+GPOFZ7NgBpDSwPf8/3um+JSZlQcv2qQTSdq1mH4
njAf7z0mTUdy9aTYGRQmlptnPJW7p70IxifFNK4Tw60cQU1v2EuE7H1+S3zk
qd3WHSUBVr/t1UJuXUrNWl4E3RtW1NAeDPoU1PP/2A7DuFtmPS+kTqP4Frzw
Bt6rF3lTxCnPxUqbD3sWFlYYNB1BPvGlwvevy37Px6QH5LQAHyHqDSCbp/xq
mLqhTqKR9GX50NKRQGDubMCdVfIasEIk6MFmq5g/w1mhniGWpNu9DBmXTyjP
0ZV6JslVPQyZ24J/MBxydfBFN7VIKNRho+tlj2nANxrVlm+3oMDR0TZfRZAL
zjPi/sMUW1by1Pbf65GFOYEiHxE5/t4ybEfVdoSdAbAW66zo7/RUqWY6OHBa
v55hz00+1mjT+j9if/rPqAQi6iBbERXVbznIZSUTWc+1zMaautvV+Ec668Db
zVvGE7OlPdvvbCcfbxuFwugOqi7JOZdGfFFFaqcsTNPIXvvSRF6i184oIyPj
tywHOxnw8XvKVM5d5rI/YzHS5WkEdvkLLHXc9x3Ze6QlefTRiz5zWW0I5e3a
p5EeCRacRxeyf6D1+e1O8IFKo2BepR6QkF0d720Oapq9U0ciPAdOx9HA0FoT
dU3PgNeKBSf8slKpAwcaDrryRz4uPiPP7+Zr0lWm3EuLjsMeiZf/SMB3+1IZ
wrT/OEYtx0gJQ6DwgZmYqqvzS30mQv8ur6q9T2Dq9kTL4tYooRhfXUgNT3w3
DHR9a3IX+19kfVrL2fqkz8oJYi4c7PnTDb9ZljgV0Z5VHXXJfrKB6B4RQ+Q4
nGrm1qxI6Os5YKdsi2g6gUKtiirxgoaberKolLW/f8uPUMegzTDoi+SiKFzi
jgd1La0TNlYHufzeuVAj6E9sixA4uPAOvORF1XOGRioh0b4pzxYOMP4LRrRR
48A+0DvCQVnf84tOXlBFvQs5iBtJlqAvNsFstWi857K52QbohWdaLiajpOOM
5IUnFtGKgg4fAI6vP9TBew3G1iEZIxEY1zQ6bYJkDgLSlipMGSPRsyEcaKVB
leEwXhxCCy6fd0Rnrnbi2WNVK8DkAqLEqim6OKk3gAUymddA44vtfOz0g2Ke
MECD0s97eV+cAf8y1c2+lhT6SxmhcmenkqMkhdkwuUQJM8a4Xr9nVyORWeWu
wA8LaYixJ0kq3prOCtUMOmvidUXRglRz+Azf3IbgaM2my7IYkz2gP5lcByFu
jlhPCceni7diCK5pVGe4IKLROEMi7Js29C0Sjhi9KnIxuG/ipXP7zCiBKhoL
wihs3+97Tz3+timkLZfVGJGIVeudrgkWDORL87Ksi6327Q4Ksq/VZNNJuyaS
QUUIAUhsb+rVt+gRHLODX4fzJ1P9k2KxUDy4/KEsQQriqgnaH+wni2pWIJV/
4g4Dyzdz95gX1Vll1MLz7tX7wKMO1BFCDPPGnGw3GrBqjtL3HQPh1CRU2x27
RiaYp9bpafmvjJrKUxUwrSYsp91YFxiw8jQRwM0OFDy1TXuRJDuMYPLqDRo2
WnmvM/rqDVwouBR7WG3EgGhLukOtMITbwiUksrUpQ5OzoJ02ivAI8T8KeBi6
LADDHkyPHebGCGgL9MtxN8wLGLulm7tglDY8NhBl3/4GzDdm0XkFRbUY3bMu
BVoJtAWyHDZj40pCDG6sElhPneAYVMifam83XwcaJmdL6INZeLPeUY7Q75ln
H49UwSvmaqgc3zF824A9/e2N0djTRXeb+hLC7RlxKV5f9THhjPEEDZu1pJZz
X6R8vPjmAoIPYKSAd3SiX47uviWh0I6Qe1Yqapjb1pAFd0sm/b8CS+yvLBPp
CqB6wIdXQerJ4Gqzq6IZ82wencgy/83De2MsAibt2DANwdLTrtzJLqI0BVkP
BzouuoupB0lNThtaUT1ikpnXA5F1COsrOWbpU0lLnMkGrj13sYNugS71M6uR
VSfemRMZK7OLZ45+nTCw2DqbfoKXpp74QfChjHzDnQYq7xG3ELAn4A2TU7AE
WJ9dpJFfxe71Vx9yYdz/7Z3E5Hpy4E63GkZQr99aZM9hDv9u+dV8uuwHILTh
2V1WX7xBDHvAZo9dVCddlyp6bqYMLeioeCn/4IKR6UF3sypKmC1Lh8ouj7Hk
UjbW3OigAEfECsDjW/FUCswbEZpygvEpxjGrJ9wfqvObhdlNYql//grlttOX
RZ0wKGDsSu+MRICt5oyV1W1h5DIcZesfrfpEgFX3ym5MS3AHBaC4/xsz0LZC
PGOjn77DUAiN5M/gW7X0S99Hu9czpcsggm41Li1gEJrY/dU8fRiqfh8wo8RS
Gdi8fli3/jUcYT7G2CETMQqZqnfApP2LAc1ZdPJEw2ADdz95liPn3I4JQo3a
WknUJAp6JZ07irxjpsI2cDuYu5cSyMKPhL9vCGjmnZ+RCcZCxqyODMmCvYPz
ZGhmbjrPF+LYB9qN8LSUSL8V5SLhStYR0KfEzRStr9eR+aQI6Z3xkARxJEVD
s0t5QotIuVUu6r5dRkiHce0v7/1px9j2kwwObyCDfH5K4kRaDv0pPmAEZiI/
t54Cm2xXiJKsi+0ZBXMMZfpGeoLbbkg1Y3J3q2O1YK9BL1BZNNhGxi6YSMrU
4h2WRAbtnoZ/hXJjFnQMB3Xff+OUo25cx1KAivuRPHnBTGHUtlvQ65JgNmG7
0A3aVhHLT0uOgJ4KKMwBBGCkpFapwIrvCT50tE637FMfCNEHrVzrXZVHm4tv
Bg+qCe6roredleUEdoFM0De6rAs6LvnzSMbZ9jyW6nZh+u5p15uX7NQZeokl
7lr8QrxcDVjzcxg7cpiaoHu3OnCM8DvzSmiA58uAVCVaz2Zg3Kr+phk8+JCQ
LWDh9/X00H8Vp7POgpZRXqpiAeh07kbl9r/w1UNKii6VEtYJ/1K48fvmmKeR
AmWZWusowvJ5MXuul9jCV/iiWGRGb95j5pNfjQUFE3UcHAf2Ecq3cfVNNyS7
9OgfTZYjLMDmjbOiPGdkcacviqk6QWxllkUAWF9mo8U+/L2UCPemXqwbSxfN
7Ua0kezFBwireA7z84NlP5C0URH6IkGS/hk3B1kNVoz8pcigabmleEsIW9sZ
8IrQzkyLO61WAOwUpibZGcFhXsAaO079TpyL+euKUXvafO2mSk5+zkcf4Ejh
IBmbVh32xj+9s7y2Xat7KdFOQoOwTjse54YugcpYtah1w67iNiJI+ObReBCr
7LIMBi9sau58EV4jvIgap3fCUFeAKwCwo0d/psf6tdurAdkw+czCddyJZc2D
ngUvdzMtbld7iEhNUz1VHfhQAH/I4u4Tcmm2BSECwBXwUx4lT4XmGw7xGai+
RLsDEBHFGNsJkyJOrcZwGekEyDsLDKtMBJr41LcaH3wM1FOhQnCPmutaK6h5
D2ywHX2KNQma9IqEicnlOxMoJ5Lxqze9c6uGGHNxPevUejovu3OOmE2fJ2c1
21Z136ZWOIx6YVdjJx8s4SNjq6CmfKdZqencvBQedtJdYsaYI2GXNfviNFhd
yBmfiP8UAWV0yAc0tsXhkDn/r5p/6sjBmPPzMc2YiRauH6C+j5EPvh6ktBN6
2HzOHLFU/wipIIndhhJlTJ7YWOlgRGTpNovC4mpj+ZN+RpTnE4hft3eL2Fpv
QrcTnflazplc/hdOvOUK1xDpJY3Q5nGNMW125HdBk6CFi9RuTQ4RxgoVxHwz
06CIO6EmJKH5A1TRkMWMhCqPvWStp178jZ+p4fZsWvIKKlF7fZGPAup5xjTg
2b4q2cOW+alU5nD9Lk7L7uvQj1sjCv6mWLEUZtbyIh73RkTRz3Ftok20uQg2
qGZUSr9nvA4XZBtpi4J1wLlLIblpeszTNwh2vYchzDzrcmcK9y0/RIV9SPFz
R0rjfTDTsvtNCyWK/QNyJ+O/asCSDHEfhOJzftvAHhws3WtjJ/ROEMNOQM9l
MunuuQZwVV8nDt7VginmDi14INS8Gs89RLGQo5OLcfL4TUSBDZ28hB63x8sE
PSoEqdzO/E2lLLkHhcwO0zmO8aSlK5aJ2AbGQ1oRXxQTSdXr6otbMCfS/y4g
dSTjikmbjO+q3qY6TAum5CtstySSZs6dLd5+jPQPImxS2qrUXCofeGyotd+K
o2F4T2Vbxo7I2F7XifloBJWBnuDDG/gaUv9SSCOmIlbLhcJdGNCSHSTtmryF
scaOFFY0X9DfgMbbcRzeCIfvin85HqbpJc3MY/EEuffeohClnF6F+R5TGhhj
OWGxX754SiN4eMdyNu/53DDV4YP07TegLOV/2FDKm3QvOaDqZKEMxmsaRRbY
aKU4E3P7/VQuY43VJILJ9s+HO+QB1bQRAt0DoJ49PSDll9tlbjJUG280ScaQ
NkiFByucc7LzJmIxJjfD94d5OzLeCvib9C6VkLx8a1NR62qlL3bFHD5bePKx
vwdylBxKPntGVuhZu4qGtLRm1pvDAMp648wP+MCADGyLHmZVaSuNrrDOdeib
n0OAToWYjOUwoumc8QEsb0Rbas+qyx7CqZaSMO88C8FH6r+uhUIqji9Dsh+8
xHVtb4lEj4wTQSbOnkte6gUcTkhcM3+JUwb0OvjPJ+Q95xKaiR+BCR/4jcCy
HdLFHCDUxZ03r062YU+JM4IhkVAetQeehPE3sp+2IGqfyOo/LuXttPq0VeFE
chfENRiAWZDXd7o+Fg8J8IKjldjg1OPTqTjk1VHSXvaWH99QEmdYmGxLRvCk
zB1MKNhF63RKcBjLU9l9Rq7W+wsz2MP2x6JwPd544pSjpOmdU1lo0jx9aYS6
LCHSUehZT6+Vr1NTKZDfXoM2Jc4V2mG3Sbpfx73RjACkOKuoZM4WI5TjyHhF
vSA4YQGrcnUuWMnppif8m4IH8sZsJMAZp0Metg8CyY8eBaTh7vHaubFLTtzD
StgMStXmtPhCyuBlbseCHAT3GUo4DZ6skm3XAumyhOZ8YMJ7pIboPWCtz5wY
C1O6yi6KbHn9texyVEV2GrHkqPmdgLjz4UmrVAh0eafT9/fjA1sKgMUvsoed
atwp+ji44g4ypwe478riLo1aFzCJ+NEBjj/egbbktO2TpTEoXyDQ21znZc9W
2o/Rwvk4vAEVaVzke206drQNTJtkqE13QQQYqmbXZn6Ew6hCfmgNdCfhlOQ5
VZE9BiofKNtrarP+G+x0zMPtHB7S+nkqP7e9AnfD7fhSIMzOZn/PVBApeyea
mqgmgCkCOtgcPTQrRjmjf/Fen6zGFaEaDeBlqU2Bi8qFAUi1+wTYDhF44At0
CTLOJMLGbJn4qdZcHFkB3OW/vc/D5FZoRlKRxUE2bBSHnIeIL/nzF43+tUUr
FTttoUGfts6olHg4eud77zDcjHuGhpJGxo4pISyyI7GmHGszHn45VoU4bAWP
eWUZrz8ACBq169D++uWB1sVedjnBrPeWwKm3zobY23BwR9fhmM5DkpezLoci
4YXrDm50iXNlpGdVzkeB0N4ljcE8iBA7u4Aj3QBMgXKGUzoZF4aNlDWVkJA8
zvOAgLrRnit0dSeZ5+FIQDkA495JF/e45aku9XciObz5BcqAqjDB4bwF1dBx
pvVsm0XzHNEvWL3+eAAYXdlU9L42Fwc28x7NbOBtdp5fdgkRtP0hCjAYRmDr
RtneZZNI4U4OXLEK+e9qnsNwdshrufa2lnUbRI8giXoijn1aDLsKKsgDZbOK
mdviyK9Zz0jAp8vnVyYvbOmTh34sJB3r+sFKtFtcuI66b6HwiYSNbi0LVCez
9thObPMCJsYefhig9FRNCz8yN4KR5Da7jQW5RN4RCB8gnHdiYSzKcoe9y3Yq
BEIQG4hr1VYoA7nzrTsni+OhOSmDT8HssN1UoO0zxvKXCAdGBfDIrohuv4T6
MLGcTf6i1A4uYndTmeSBINQgNC23lLG/K80bL68nwM3IWhlveMLn85cY11F6
GZJHT2qJaxkMoF890Y/xUsYl9R7TEm34uD28yVrugUekkKFU6jcKLS61qOsn
r7JHPcAB5++Y06lgxxgwNlxy7sSiTwVfj30DI40dJw0GWBU6a10dBroOdtAX
9nUEXztJ18Jz5SNr43f5R6Jp+4IjngGm9XmIuCwK1N2HzXQ0PC6kNespOM15
0KNGdZNqD4XYaPLzgGzSIp3DSWy0lR5PFs+bD+6b52a+qkN2uxUjt7SSegv+
4hpZhvEwhdWP1ecDhaoxsY/55XILgcgDY6iKyXtD8107LeqxVeFgkbAUeJt0
jwz3uQ6+HhHJEL+gjxIVYmIIKgFD+l1Df9kXIqfibF4C/4OIxLpncXqBM7f7
0S9vEbNV3XjVvX+TdNW0ceoNUb+mxWtr1EV/91ZWeR9u7CrkB+uuX03BH5Bi
VgaYd9JBtAwX7p5qWLk6HAu8qdati2fi2V9Bn0hcHB2N1HUC0PpicfwZuNrj
B5i8gpp3M//F30cBj1XSB0IBysrF+eRS7MzgTu49hKjnYs1bVtDVtpDzE3u6
YnK0MNKkVcU/tx1OHaXXFAwX4inCA6pnX2qBn1z42cX+7hWYwoZ7coo3ZvGw
9F0uv8HBAkmU3N/ftmNczASpOg+ZDEcqFgezKk5tuzA8UBiNIm+XANn55pxM
vThNFb/1v5qRXS5Sc7RJD+tkk+VfjXv9lTh/l7u3pFRGNqWSyBWwLRYaHj8S
+7xIP0HuA6Jqf9ZU8BGUurxywMO5H21J2dtxAJ/6faclt3tTm0aZQPbj/P10
L/EJRc7ZQniS2BcQNx3A9HUoM+0E5+jGlKOKJ16hA8MCxa4lzdXP36qw0+9Q
9J2C2lhrmQxKlaK8FQPdiPIiUgLbJX7SAXM3/oRv/ToA06vOP1vLicWMB75O
mSUblLAkhzIQTYlBE28RGWuksX1jrsD6053IU83cG5A7G9rynEvkFjwwS7E8
ffjyZ0vh60DmFE0aik+xBwVtUIa9RaxJETR6Lh8qHAu/JXXs+fxRpBC0Urpe
Mu0aAVR2CavGSlJSwoPtQvIsG8i1+obsdqZ7mHxNX8e8rdmZcX4c9OMPdZep
Kox+jPEDHpa7XEH+92LYZk1v6vs2u3M0H700HaB8e7FW9ty2NlnMQJnCth3L
i+TPHm8lRRorCIU5FPK9r+gkk8CSvSuKHQxAqpGHguNCrR5RZ8B3OeuFcfzs
09l6b5uGCQ1NvXcd3NbNW+Kzmml4v0KMmmiMTjI+Vz9h0tYSi3haprW9DKiz
wIfHI0yk8XVhrUeBvDfK6H/C9insSKk7FT6fKrsFIVyJ1ZIm9BMpyjB+1Sk5
dZB5bO9tjfCKkviNnyfws8E121tkqnIZ5XTmcc+7NcoribEZ2J3yOR46apMR
giS873PXmkGIqz0nKEdICSBtsOwOzsayEMnx/ZzafaAUADOj2ogE26JpEGNP
76uw6cJJr4wZLZ5zXg4oFLPseIBw4Ga/0YX9g3idQM8rLF362GmjBfEPeRUd
nw4S/1lUCvHT1rbu0UM51WxCi9yOEe3ec5vt2RrXrFop50bqGozpZ7Lve8BV
r2KB9SzdCEjXf/GkmLXRrbMY+ZZhDkwS/dDMym6uQXCBaoNvH+8N1XpsmABJ
tfkbLdNkQs/irSaFbjoJ59+Ttn7MKr116cEWGsDAtTgtqnBvn/RC/O6vMFsB
h9gNlPryIgEUayxrtJzkYcjHRFNpX6LwbZFmtK5c/Pe3Kkt0tdj6tBTOievi
WSJM6gvhAE8ZWYUjM10NHg/LfW5CcVRznPYmkBf6f0NBJWzp9ibCXqyb2H5P
SapGKpNAsTWH9DSqUJA1InSuZVUprQvy8qa0hKR4kN9DklPP7LpYht3gfV6T
/vSAmMKjatCdKD7Qrl/Xl2CYIZi0AbfJ/yE3y92fHlj42gsLtsyf69ZDz24f
Ijv7cYbSvCOb6ypMt23SXimZ2UI3cI7PfZHm5PWyyIGbIHOwYH3nZqpTTAK6
k0PP+3SMEVFp8q90KKmmiCbnXXyUSRyXdE8m+f2xPAcGxGSN0Wo4xBn2Mcgv
ZG3+o2CBQxGmLXfAylg3RkKbhAsqceQxYIZwLMzp6Y/n1U2R1bJRnrWRsg4Q
WMnC00GNks+y6MUyQnMYLgy2vf8+q3f4os6YXabNQvOSCOzd3BEGYPjVYLnO
7ZSIGy7TRxdb4G4NURxJc6ZXdcBqYyRLvJXOOu1RL0zA0plGCxfKjUk2qPjM
1DmyEL7wHOJT3Jn9CGb6dl2yHsq1RJ/0K1MhIeD8dVg+1jrJAS6Z2EZYYgrj
NZ2hUz58bEhW6RCQRbr/Ligg6ky85Ibg9M+IB80MBbrfZhvVSDbxwG5h/7Vm
/quMZLlBQ+Ukum0JqQ2kk310ChyPbjEdE0dyIyotQqeSaWoz+S4cAysSbiGK
fhy3FSExQ5N0Q6Mybln6vb9wAnpImgoe6WK/0dYyWocmI9ImQGsQdm5cRhmM
LoAFuqPp/0UjH7pX8CCyySyfof2+T9Sde8Em6M5cmt35b6uC9jspso+Bw/qM
qrwxZ/PtVr9VAV79xCXxFeYVUblYpvFDZKYRVGgg6Jaqq4w6SjNWnxZFG3zx
h11gSPCqFqmOdLtOGM9xzKfpaDR/Bbn2xS64OR2mzlPF3pYfYZSc1F0jcbg5
vczB/SfgyqHax9GZ/f1r5U3+qMttBvqOvF46F5oEC2SwGZKPGFsb3+cO1HKC
+KFavk2TNp9SuHjwh8iqFhs+/ZDCBDezi85eOXJoPAU9bvFEYEA3atAgOwPw
crejBhkA5ln5HxBaBScyO8XqBZf1/5hkB0x26erW45/UqN61Rd0ZbXe0MgJo
aAWS6HEuhvLlkUqXX08VDm/E+G9t0gHkrzT3v3yJFiSG4kteh4an3Cscdpzq
nClgFTQ2jF3YJV+cWAft3BwmBzsEm0YKF3i5utzn61MrJeBeyxpw0LO5wGtO
sQO6O5IMh80rkkwJTxKwchB95VdlmvnhUwl81AQGtXfNtfY7Ammcpq5Fd3ov
6S16FR6XYfMFEdCmoNZp2swr382+J5V7PcsW+deudjcEH06bj+fjSGh12vjg
Zu/aQQkCYodPtBxY9d1dQMUxcQDxf14GSoS5LEp3ijhFnniEW2gLizDDnPWK
I8YxlOWsTWXxOtvCotkNeD/ivC6gbsgE4Wmc8AG86+O/bv8tUpbQSyH59wX6
qD6EZSlHPBM43+MYiWtiM6HMXmbKlX4kHSnkSsQ4sfiNasuTeMuy26xF0axt
UCexx5pUdmSTpgjCD3B81ka2yTo4/lDmHPpO+s42UZN6Jc80RWUlT3EAWloQ
6BtjZkZr2kC5S/+taC82oYkJv0uclJe7UayExdbl1kqs/QU4Las4Wo7/F8Xn
iKtYRhgs02dCRL6uB6d+Sv6MNONKAxgVZAWJ508DmBFtR+sTcpVYb5pdEUJj
ncs6II27LFLgyBe103pfp4++F1nZpwVObb0SJRTMj1hh4iiXy8sTK5xIg+N0
wogdDd4BNJuLIa1yqhPMavVEwaFTwT6Y3Y4P7xkP24pg4HDAbsXmSRMAj0SN
YqFeaGAfKe3w17kmCNe/Ysp7UDv5tY72bWN9NJs2AH6xyJ7j83ck26hFdhJp
AeBzmbrv6UVlEI2T9KNPlhtka4ficDMoFHmLGJZlYb4cDe6O+b5mMNMoxuNm
mjzXeVIkMnL2Gz4/MZLRbH7Hb4FCwhjaUpt3OwBwwLoo+3feoXzev3Daw586
SZJNQH6+Fw3OJfywPTQlh43HOm3ylx5KtlZmj1RZSd8Nw+RJn86M16/N/pCz
BJOH8hJCvJRVBdVXHehGRFsky1DGoajF6rcjXuEbLA/6TNvYexXv4Z2339L7
bimrsKEJ+oqn910ICQXVj59xk/7lh4xzc+igRKpJN8bZZYei87Rb3migW7+8
yu5VVjSHHBDkA0VR0+qKkN5actBML5ocsGT8hdYNtenTRekH/f3gipdmXg49
r/ddYXfJvccdNNKd8jJ2T/f+naQtRQERZ1qNcVopaY2mg60KtvB7NlwnStWf
Too00o6M+VWW0e3VXXCmKp8Xnem5K5sQdgrF0MwoyHOYag409uxJwUbhQ0k8
T3+QB++cxEZGVTyuuI4pDeTM8XWowW8cnLq9o9/qe9u6AY7OF8gKTDEZT6VE
FrRHZ5+GrY+dnaDpN4kEf8mEqZ0L/ZsKHPUK4lngLmyZ1KOigrar67HYmor9
rkreq5aR3lADFZTUt59SNQjI4ob8ng+YhWTxb/fth4cZd3ggEOOVuMC2RhaE
a7q0wPDNF4xvDbiGXOkFFlkP9As8FCFqCpPTCV4XdML23LDdmxyVB0iAxMiz
F1RLx+Ol93DlD2MiWWHQQ5SGu9T4Q7y9cV/IqJFt6qrSjTV3MZh0r93XLK/L
aUlsEgpomJX3s1RzOSsZ0zFvla1CCF8ZCIShldzenHj9gt/prdFyet3w3IMr
Y5t6MmncEFsCltWqfAT/gv2I3NNlmDFliBLQSBWj3Fm0P1SSFK2jc4IN9L42
GxuLeMRm5sB+BR1+gRba8MwcFNEwq/6OcSdZgLFYpP51y6AnW2031UsFaLKk
vhPqv0VEMyFy8L0jwzKq5XP/MK1i6NWHw2H2sAV79Et5R6Af+d0rjG9IO0vO
VFduWi2lC2EFkPGhQVbc+q1CbsQp8BlOw1PSdt5g5N710sox9kt2d0Sy+hij
N6zAa5pwrRoyVEaQ6n9LeNaubCfkpm0GmwdT9r0QzML6T3wA9OIVb0b9s64q
xwXtO/zoOJOdj5w08hY7gDTHZrdJlk0etMjwK1lpzK4R1bLSc5FS7HdLK0fC
Bjz0fvBzlcMLa6/aaLGQ/3WA2J94E+aj1wqZS4Bc6OeaXS5I/bjOimHy9lbS
SQw9uHLBpQQ3wcU/dUYfeOlzmyabyrIKF6chLQNTE57n0ChOz/hXyC/SSP+n
O279Kh/twy352SIl9cXJWrdLIHTvqBQWF6pxy8lLEEjV7J8dP1q0SU95f2vE
We6+L+anjwmort0O960IgCz1t7Hou5XR1pA1mCQ63AvgKfWBAbaWMWiORm8u
IaD1pS3oA51aiv+mzN4rhW4WtkAPWq0iQ/TiDhabYufbcgVzpgu0i6tUh23H
kgXFfQB6o22KaVAp7pe51CuZEEOJuj83B9QavP/XRm6bxPYyNGUaVtluED2i
pczyFde0G9/fPv4hJgWjVRBnvYD6quBAWY5VpgisGngmkYo3GwVWZ9ITlUYk
JenitanZA0AQQBGq3rnaHK7eJ+kI7E8/+vTh5bsq6JVX6TLA+EQpNTKnV+Qm
9qPN36AhtCo8kjVXD9rIhMKBNWyPDXrK7rpclS6Xw3xOuQa7YYs5uAA+VIXB
OHbQkCHbXiD81TfbLkbWWzQP+z4cEFJm5utGbm2vSXmUuD1xf1IlU8X73V1A
V8M0B2SD5P72Rm8BJBQ4eiq1Z8LFQaLJi4IdNJJ5opRoeuTFqXsDOQuxo3UF
LSigFcmfW61edfJinJQFcHjY2wQ7paAQuefY+mIdY8R/+LEYCieLmFRHtHro
Yc9aQoXDa+fBOEilZLJMr3brexYjQh0xUz/tQG0BQJkMDQnPKceSvNLAdvyi
rgBbUYHlxElPfWtqORkzos36KxySPk2TmCkxx+kvU0bdz3c/K0NcD1HHDBM7
GNDY9OwtHNj14odok95VTtik4sq0ty0fGrqmo5i2bhZy1nkqaNZkVkr09nHj
i46wPitQQ6b0tfd8GUo8rftzSSNn3+SozemFhr0oUz2Jqi40IUyF/KSBwxYT
45EaW2ch2b9CL2N59YGMwRAuWtoomkast3o69BpRzQzj2wBlARaJysZy4tT6
+el0pKRdkpOMCzhcsv6ijCTlkyZ9h0t5WR8XJexzyi2xFu6syEVU59nmifUm
0XGxLKw1g1iaGhrfri/IpFizyj3lROYrM1iwoQ1Ft1uH3h4reTPqMDgQ2Gw8
5cu6PH9sAjFwU7tfK7V2oilt3d8uuUb7ehqktJOdU+gaTBmpXr4/g3yU9hkT
msXo3yi2qI0NIf4qaG7DGDF0kYbXy462fSpUR3UeidZkoqbce9sT+oOmgBgr
cmH8wpH4bVkR/2haR35w/KweBaqbVbkezhnoEC7dy7ty2JJESbCVkxP8pga1
8PAfniXcg/aKbkyKCcWQF6fbergFLduBCOr3zA+1LPODkzx+W8T6/hn0ao37
HQOS2XjC5y8sJ3wMw4ivKtO+LjeIRdYyecm+9u0JDQtuMMnhxK0DAI2vKIfd
kX0CbvFqC1WnORJkrHcWX7zHiE6qr6msh4QTO4keh74RoQi1rF5FmCMmMRBH
QJuzeGt1XhfxYUUmsJ9cTCPrv7YiFY1ae0NsyR4jU+QezLKUUdiFyJPPmoe8
+eoxLBeJI7JW72G68iH9P3VSfprAKzAM7QYVpftA4iz9y3A8HzeDboGWDUvd
5nCoBkAupQLBxB7HUlD8l30E3dwR+2VWC+9WWpa2WVw2Ddjua7g8XXERe/0i
yb7J5fkqOx69vHAxBn2IJ/TOgzJG4ViTAqJbmzT6ZKQOWtMFAQhVVnZ2i5mC
aIlbCoM8gR3qOFs6xPcI++2j9MfUKwdXu60t3WLrqAkJhbuI7y7YsEN0SLNY
fytWNup+t97izf6EkhoJWfpoRPECGD+9CJGICbNsu8Os+rxfFkpwUpAePYu2
T8FqgnlPvv3RKwIsuj1hUonxPeRYH3SxPRvZy4aBin/5tARSoC98vqjFy3qU
g0mS2eCFO/jJwdUO7gpkKbbeSvF83Z9hUPUOq72Fut4eIGmPScoC+GuPDC73
j5no4b+7fkuxM3S940Ifn66qBMaF12qEMwBx077OXZ5+wwiI0YCRsbno0FAE
yQ8LkBlownocqHEoUFyszfZdySjU/RyFwXsEwEMkdu8/Nz083LebbYyTUXk+
nMh9ik2uUfpaww7kqSYFp9ag6RkZFj6s/nMbq0HwjRLszXfWm5NViuw/2UBG
n5y4j1KsPBm1f0g+FALbqllXeZUKJ+Iw737cd4/qLBYOHqpeLoFz5bG/8kxU
9q8oI5ojQQ/P1625qCD/Zn0OrWNqWeUqX/ZZkUrvbNk+mp/1JttyVP1Hrbnf
SSN3IzyE0W9vbmWGmguKjKf6hcvDhC5PyV3VYMu5EGpkREPIIJV/oHDSbSAD
z8Mv+G3eNZXZqimx+W9EtcSUu+ZtTQVbsRYiw7yaeDlm5rF7fJoT18LbUdTc
4AO3tMWmWmB6hXFlxje3cFuHWilNKoOa9CjyibVbDz3KjiA6hIjaJ5kBaniH
/zZIoe88IzMGUQ09+x/uu1xcAfGlzImGliMxYja9bRRGFRrBsJVvLXa0aQr2
TjhQURULWbl2Vnoq1C3oY0uSNm+ce3bc2yEojx23gTCif9V/QisRil4OoIsi
oUGOV5bVJT8MGOaVYzcQa67+6ZwWBW/q1H4SIsUzDUZTaFBZACgI6B3h6as6
X8slx6POAc8CK/ZwUMp4AHB3t4H+IPCpw8APYizS08GSoRODdsaG1JHmRXFm
rx7JF9Tvj2nZqmMVuVSp63PFLZNZVqLz4kJcfhEkR7fQT/7H6ZgBA5zlCPGZ
gzbirNl7YDg1kYvnSWoQw4jT1hkrxfAv1ghJVSsDfHggr/r+YaRUOMUtGC0Q
5s4yt/PLuYpIwshgX+EOsfiYMNW9Ii+4wxPtBr6NSeMsyc+c0D5F+mJrLKje
Jb0viX/om65qYDBTxuGnJvc6az3OM5S2zoJQvfn9iStKC7fFx1j5UEodVpUZ
nnARYlhbGgNG9zn9ExHd9EzwTadZGkp4alx9JmSRywo/iAeCZkQ/o+Al6POj
JzuJ3De13CQ8w2JrlJ+HNKZsNgr8Pn3Txd7+foBecG8tnsbBRYO5JXVamUvL
Pzff791byTpqBHuot7VqjoEeOSPNJNhfaGEP55mMUDBRHvd0TJk5XEeY58fW
JN8Bt1Brh8THAMZXb+MzDrMXTMkIvbevEQcKTPuEEBgFp7w2cpXy4NI2GceV
NZScxwjcoQ0Ed269I8+ITwL2Rm5YWKwWWT0yKdIVLyIBPC/9QfCRxcOnH5iH
NxyZZvsLKzDNSfMS8ZBaMR7jvge31RBLgjajvw+97T1DBEKToyzPt2lzpQez
lvw8ZMDy+551dWTzyY2HEt7I5Rr1o7IDScLBEzhzOO9h1B1dqJlosISZKoba
0ct6l9pE9XtYmYXSqYpptXqHOCR4wIWpxtVBvRx4YTFgFLNAKbIBt4fIVQM/
UBqlDYBlK4rNjzXcob+EoGnu/o51gQzIrdYjuCq2ofNo/pcuT7Q8cgyXIU7c
yLj+yEnLJGBtAg9u4xyhhEiiZwKcS7Rwtjs3vSsf+t2d2P093bPirUnGdU49
8m6+aolNR93Fq+UZC3eI1MY5vtBXG4UKAn0i5bEVKXA7M5U93zcQ7jWq7UdU
Pw/PfFdSPQAQjxR+4uZOXWC1qTRaIc4F7wsxEe5YKZGNm3810U8hHkXzugzq
pJxSym9hBLqqI1PZO0KhSCp01XNEsqORj+coM07wi+Ha5e/7skLCZaiZeFAQ
vFXrJJvkGeBdt6sOjmttZYo0Dn4tivHwq9Gn593S/9iajLVtnD7SALUjFqpN
br8HcitZwdOUdQ+VSajJrW0qhxihU7lWJQie2IabdINuKM0WhZp4xmijIOe3
cCkOLjKyi+RnPYvdLRixSTzNsTvqJ6FFgQKX0qdGS6KN2JMCo/QYntmpmL7o
WsT9Axrhk37eM9DFSqKxE0dGRcDeh8Z+8R+SuzwfLHVjCnPJ00hwJ6kJjaTo
csYsjZmSdmSnJMCnRVOMid9KXlkPlkiwwPKEOn0fdsq+R23+BoGgYuubOpXv
CbHgRN81ccYaMfxF94zZIR+71NiUAkdnVQn/rCDdpaNJB5azSF6s/IDraa7Y
eP0qbSZvTPwNxmielob8uyfbE9XEf1Njj/tyxm//IaVApJJjK46Un48n1RLy
LMzBh5b0ebi+3WYeKQHJuHtL1hg6b7l/6O8myobBEnPyPRDEMPS4ntO3oJ7G
tiKDuJWO8x+or1LvjaTesK1M1W2Pg+vLa5khvoHwKfHesNJFvh7nV1fcT44V
Ctskjx/ZmFaFYfpUxd6YKNXwQaSpQj7HxhTSZA0elrq+C7ZlEI2WzuIWEq9p
+DZzhN7LspW92oP/CQ3vLHk95afNaIkp9UMGaI/JOzqUgMsUcJdnBh+dCt7i
8sAMLnFycsuq8j4ZQaiGwYC8nK0PncEVl+/bwJ5DthnMVOSJbRxf/OClzxIC
MFL3/lXWSc0Qsj2zLaEFvPPiwZifSdKY+XA6qKxDOjfigdqvYqzXmi1WLufY
sXSLwdK3MEIbtoLSf7zSCi+kDpvMQ5QDzbeugEV+bsv8r7Cew83GE7+oT56t
SD1I+ZuioGQFqXBuecD1eWxHmP+U0OjkmjM+py1T5UBUbTwFIKHZnRaDT2/r
y8GDyaUMm42RiMIBsI/KNhLHI4DH8YK1pebh16qzMCCvPRP8B1F4GrbgA550
uAW8g1xKtBfxY9vhd8y6ziD407RSIUBQ8VJ8kQ0fXZNfH2HSzkHULqr/VwMB
iYO0th3EIwhTuPfl+AmlGj5IxFU5OO1ss84QVrXznHlwQU20FnK4+ivnqFd5
OgHH0eqZ8pZx6uTWmoUE+Xpf2yGv8evvf0V3QGQwGlz8ik5Nrg+lrCR38NwU
9kUPDTssSPvyfw8/QQfMOksAtUvaWxOv13732Fry+gbeTtww8I0XsnkT7P11
9G1+n0bD26OlOfoXpuj6SAGG0P9XBqNynq6+ynvnF4NpeXXcyhjaNSO7DMsQ
zIJwr5demDWZirBoM0ZVmSo3HmiKsdbl6R5VtF9RruHH4C2ATsPayZVlHdw9
wPPbEQ4DJwkPzzbNmOjE4ANEDEHQ8+6kNuHQwASiXvLo5rJVstfs63Zq0EwH
oSn6Czy+8ndUDNzLyLA6wC8kO0Cf4jxhE50uE65m9nD0n9VoqEpKZw8bb4Kz
ndNpPO310c898kyqeH3fwDKkziLrHany7vQYrjhdNLZ6+Ao94lqos+Bwz9Rz
XUE6c2zJ8++3YizWjDdOrCtuhe2bhBSHZQuQLUULVIrdzOHKofkPlGaJ2Ewr
nkO5kWzZfck56Jbee8aTaNBm28ZQ1KEOQwQv8J11cEPxv/ZwHs+z7vDi6wE8
JdujRsqfxYCNuH0uBCHvjfnBblgRYf6mt+VAGN66NjoMr2PlPxtKjDwybsoc
67Y6Bbz4yGbx3uLcWGWBK58fg0UJ2s++kLxz/7KGieqh1WPvWayywx9Pqobk
jAa8vZ3ytaTsEYF3ZF83EyfKKUTTG3nDzdmZrXEVqunaeAurawhR5PrLf9L5
zQauQrh6dlE/D7IjFUTn9GSLnjlpuCBIDmU2nz5MGtZrnqAHPQy0aAahTW4A
Iik/1stMpFk+I0NrhFmaDlNXsk9X8pRv+4fi2i9/pPWh/crv93SpM6nmhwJI
MjKqXuLWoU8/dx5GVOAnrYbA5zqjAIeEWfEtX5rLBSQmDVM4jmkA1/Rrnf87
5zJNFEFskxAtEtUx5dLe3H3aAGZ2R4XCFQCGb2DIAYn2Ldi1RwnX0W+kyMla
4d0qt12IJ9H6xzudyS1owdaqjVymLaZTZMn8NOrJLmket/ZxLgx4nkthOsLf
pq8ARoHILmgjHEKaBtArce2WIm0UgbChKYEZkNNMDV4wl7FcRAaLVRJdwk3a
d34hA3IkPbHNQHb3DQVJ73c9EAYRiJ62R+X9+HhO30epYwQseaGfCjgwh8w3
UIw/ElVFvpB7kVH4Cr3769jlP/1vXBFVSShI1pfO31NJtpBTJTkOptE7Ymk+
TyQuY3Tcn5Q7DD+1lv7GGX8pROX3d2Fz6zr58TlGYunVHpLxCOQs96q91WcF
te+RciCD1zPCBrb+t867gRFkoOoj7V14pzooN1TqBGnk3Lvms7RYeT25xzKL
RAcqHnxJagMpG4F7dJP7g7IU1HeyiVkdLiv8Vll0OHnXh1v70aRMtGb0jqw+
xL2NUwXUzzNuefF+mFwBNT0qt8EqvEP0w4bL6BOe7YxVH+MdX1oXsf3Hx2bR
Vfj9sD4pYntPUAX3b+d/7h/gjlFeKXhMkYQ+xgojYeiOCZC5qg+zzSu6o1Z3
satqrdiyAZVIHGdHYx1MC0q9WT2fIrVtSsTDHrxkEFA6MxCy3XvW2nCb53IX
JwZM7xo5PnJapmMMl3wAyjHLzaRZ0fZ+gGhLyorqpmZ57GFNuyLOoQASFmum
jtn2KWWQPGdD33AdzrkXB4xRXhHdkzYVDcjhtUDPn1YBFcsyvxunSm4CGYCY
vO7BQsxZfiPg3rVVQi3jgYlRYTnCc101bV4Ao3elhJ0Q7K8MYrQ4+A0tQlJ9
8lHUWQUzRPijJ2TK5YDNpzlZNZ4EuoMm+qGFoqSSWxajZfzzTYBrjsuvzrSz
lxQrNr3Y+5eF4U5g3xAa/AknwRbhDm/WZv4LY+vNfFZm1EQJuitP7j/Y+XTq
d7T2165hlJaf9Q1M52pdNBYduqi/Fyh+BMBuMolZAyqu0Ckoj5gbNpJNxuk7
/7BblDyTN6fgaL3N78i3294GuwbPa+kx1Jxcx3bLJoKh8EMEHVheDJBvM4dl
GIR1LspWputFwgkMa1DP1bip3XXf3AU/c1Ga26gV0sd0QzlJy46JlsjS31OW
TLx/kYL/tNJ99cc6jii/eWkRXqNr8Upy+up1Sw862vxXrIITRDFP2N2QMTMK
WKA5dTpiw9e0eagpCI0yAIVNI+CnfQaJaYPCeJfjhREw5vSzZMg5XenNAAxY
9QkUWDwkFznCVhUrK+oGJnwjUzTxR0Q34EKCQD8y3/kZ5EhP59iU2UrDZhcs
pofJXteidz6rbuaWSGr5xh8+wd6mKVeO8qsLrPQ66O+vsxWo/T+7t3bVmdkw
khbuJiu9fHjxNiEIMtVE6dJML7UL9lC0avstNwIgrY70L2E4yvLNbUuMb9TQ
oO3A37e2pJB9SJE0GsZ23IecTrBFt9NPR3WCkvD1jklJaWirS7lmSJsIrKXq
FF9cG6ERA1eqFylwMJVLqykAtovdO2E/sZdTFho+jYjaguluSp8ZG248ibbi
4rD1l81jZp6rrstsedmHobEbB/DTFJwPdu1lruIKcw+BxmbcpQdNR9G1z/kD
DoWtn2w4ww4aRsHVFkP36z2P+csl5FIcjyRiJjKGIXZ435pxh1gFpkOPWDgQ
13aifQFZkC0cwMVF/M0TCoQF2gHGTB2HKwkZUyileR8ZHOe3a6gZGKg4+H9f
tWfytB8dR6yhhC4pL5DDuzngiadP90jOF+Vc8mBQexu9ffS6BpycuVfDn9IB
rr7X0j0hFkBa2DAmkcHWyrSmgHAhYh/3wUVGKhR9gtupRy6FlbO/BXf6Bb80
IKA7jhQOwqccABeX/SVEZ7LI94HJjvPGgZyl0Scpqbcs93vfTgzuCgfA2Hv2
SaIS1SCNHPb1iTu1LCElgdeaZNyjGfmub8zy29tbfypsxSKVYSk+IMsHR7zE
4gbLFezZr2oAIpBkSTBe+04zkTGkmamt/qnNyFkMO+cA7WNJPJ54J6RWnG6K
oGyfEAAefpkqy6V13vYqXcsX5f7IMu+0E/CGyJGzEo9erMJlDX9V1jIfm+DS
7GTSLx83XYzwfxV0c7yQtGhX4TfV5P/CSBeUkNypuUn8x4Y2G57T5Lr+80lZ
pOk5bDoMMIRqwXaE4psuPQKS2gWbR64ZyVv1bnUaE5caQlyxv8CGGdaoa1Ne
57m3RrLrf+NDVZd99MOGNJw2LU9+7AngVaQMmiXjOQ/GAnDsK9nbYG+iRR0v
gsSUV8dNaZq0b+dFWlSHAvmRJUeiDG/p+hKXymxZQyAqoGrGtH6n94rn05CQ
/SHDyjuyJHX4jSFfKNpHlnZZr9/YSHieqF/IDHoifTfnowAcwqI7oEfNc6qP
X8/QFGw85/8vsCW0zMKsbm5QT4Qbm+aKFghxbsV+EDvB2Pl1FOXLLax2aQKB
8V7RRYFr7YIgEmyBDJUJkHdl57SKIyXaSC5Zba0dYjuYY2rmREYl7pI7DN3R
bobAeLYzxek3VRMOLU9YTjLdpZhCfLqEN1TCr862HYw9OrVX/Di5KNKsdVXE
cM5djCmDzXLUDAoEk1hYXDa2r0xkqyucDnyT5ZZREjhGr3j23JJZIYl3kuVF
NRVIj0JnL646uWQ161OH7OzySQJa68YczpVu6Qn/2ki1LGHKj068IoFeRYNe
GzkxfKzF+ftuSdE9u2q2NO6W0H0GVolcDTsUL6GyrS0EGdRNnImolApQvggz
txZzK+2scApYDJI5FJ9hHTzRz/5u6kfJq1HZ/3iA3RdMnrvEz2U0cxyHDHOS
CL+1dWPgscn/OnIozsKkWbXGHKu1K6IACrobHTPQYHjVuItdN1DF4t4NI3Hu
krzpGICrmFOEf6HA7ONhmaX8xP7zOzryB/A7Bhvo56dyNCq7t3wL5RBeAoCZ
Kx9j5tiXHadYITXJrrVBAuEcWICOzxOCR+NAeFSdIVHNSi8FDKc+kEBHvlKN
x7jWfR1rSQS7Jz3RiyaG/+KxtLckQkexk3WIqxU2tH78M4PlhGg7zHgtW7Ju
jskHgBcA0Se69UDPThhB+26P2z9jAUk3paIxqEOGXu7kHIGIyN1ap5Us0eW4
RFSPFmDFFLMjnTe+p/b2uJrebsZyUm0ZtU7tzQVp1y8PBFbfzPMe5R2mZX+Z
NAJmrXKDKvDA2drBckFzhaxFvOYL6dcXpA+WrZI04H7W3uKodoMdWP4WviOL
5r1dDcKJebLoYdgGXFQ0tE4cgKkPeYE50r3YaDYyvDJdG+jeOoOEH7HJZlaJ
2WRzFrJ89ZWMaD0ARXpz0kSPtp+tbSXH710sr/6OFsSx50eWFotk5m2vJTA3
+WW69uJgoZKjZCItqyhCdqeCAefAlPkBPzvhai1gNYa0POCiRatMe8fwa/LI
CcJ2pB5m4M/aByi2AUaiY3qPCs7aXJ21z8lrzhG1p00nXNgMjTEcdJn6J2LQ
UwXvHuxFCTepEhvUpjd+gfAHawe5cSMKHQ8yPg1bW1si/oUAROt7QAbV//+X
opd9Nte+/tghlcY6Pu+gdIW9aOHygBpyzwbX2xq9UhiahVmcZsG31q+4yVDR
4XMOudkYNyhu+HBN2DyZfnZlWb0lq83RyYTNPLHwIL5sccJYRVzsFgXw8SiD
1CtErtx6GS2NgtrE5105hWPwjiYwrrgMHtKEOK3Qp1lVqSBIdiSN7OAE2GFc
T+7tPDUBgT4GWy1D9dWRZDWx33xdBSBu4tvlZepWpcM8JWrV16bGP9hE6Q27
1VVIMVayeDMu1mrc/IjUUgJMbT4+/lMTIOJkDwp9iv9qdFkXc26j+APfF+TF
lh4LNDUSK0Gq13Sbf5taJ9y6L5ORbc3wLqXntiJMtRBNtYyiIncq+i2kbNX4
riW7526OKYZ+HoGGvSl41p15oQ+/MmZgTHHgGBWRYswr0slq5eWkXzBiZRMc
j+qfrtbKUSlyxWPwe6nGpRUB/hO4sGzyGEew7ELzzjQeSxZ7UTlPVR/cdDA+
8sppygrUb0rQYs/rogpX4l8bN87TrH1SVYEOwxhZ8fYVUwGxnBrFU8iHkdlI
qDD6tL1FLTdLtRLXhUHBzZlGAJGrQbjBPnMADL+F/yUDX8+Mhw0j2mTbHmPs
KWTvBaB3BWIy5YYBHN4OPl5A4QC0DZVkEk8FeQaUDAcv1XfObM3ZDlB1W9fO
PLup15tsVTkbcEGkqAUXgWAOioWbrxPco6DYZG1DOJSmRzBtgGOlk/qqUXa4
XcIJJevrwJMtllrOOfJdo6gWkVhqmUykCWXVA7FLpMBwomhWByRhwNj9Kqdp
cSFHol6lRN++ZDsS9U6UnywNuR/QB8QHxxs4oNk2ldYWOYOWHHAKLDygSNFX
iZiYhjsUs3QT7iQMdimI5A/fhVQGWBBT05sE6jomH+w8W1/M6BrvbIYRNFci
Bdu9GmBVieTv8iEjDOVsoteqFGXGi4EynOWGnTLaTuHkO5Fq53pVa0UderzE
pxfRK25KahH+xET5QgSfeX3uGrrNzvJ9UrmjCaZIYEBO+LvnJIgGIARjFrPh
Edegj2i2rkqnbkellbchrbZ0VPY56pWPkTkcbop1IfqbjdoUvdpiT1vggQby
5d8rUu7Dw1i1rIt3mxCQwrDd+/nuWzMxQWlKDTA/0TPJ4qSD3SHS+4unCFcf
Wq7F0nSgmuwmWEIxSb//cSBMhfRklsbbL3JDA/OUdyrMeT94+aDxKZP+Lyoa
r/XgnLlmStHfxGQBfJoAoX9a6x+gHqdvttYpJDWF8KeQ7UgZLiN8cF4eNi/1
OtnwJ0M+DME8dOUCY+PY5c2uMw393KmtB22hcVTaAc2ZAJeunxXImxxfbCCk
WROToD/rmnX7KZr4kRVh+f1pTdnap4hPJowoTZHpIKvtoOup4eG3sOOlW6a6
/qwAw8aZbaonG35lYBiPSFNVsXIqrdxGZ+sAdNMDMBnBG48fDVyuYhMLY+0b
l4LHJnquE0uH4GXJ+3jV1cSDXMd0UREGra7qWAX+MIqQEkbywdB1ciinlnGS
byk63lp8vx6FAohZLag36iQ26tMjkubwc5ZqdCQdBABr5KsgcBtK+aaTgOEi
NRdtI8ZU1pnkgyGlOgv3gk6fmqvy1goRPfOH1UkOaWsaS56VBRbPZ+Q5ifcy
2rpB9sjqctZrgBDn0C6DDwv4KIDVxl7c5K/y1f5EpIXGio1ZSroV+Loiqx7Q
9QJ25dEnckKSDv9WlGbpqQXitm19Cta9mIGLcphvQjmF2QRxqJpDohfdOJAa
45C6O+/2d8f2pUpftU7g8bPj0OLb5/0ENBKchwBCEO5YQtqBYycUKSr/SxVX
nxSSuNnGukoP2gk41DYHv/QxevLN30dnzfV6Dj0fVIXJl8pnbwNYTOFcgJmb
Q2tFD8YuW2OpKfl2Ty3oKRmBFnpK9pmwRp57Qnqs73eIFSEuao5YF1tRqW28
vKgjpi23gXMOfKmQpN00IXpG+M7Xa3FNAB9Ql2OdIDFuiWiwnDCsVvA9uCea
sY0NO8yr/SuUrIzLyOBD69XY/bvymaWc9TpNkPy0j3f0hOaIt54xAac18YjD
XR5BzVXP6sBxD8GJ6aaruWC5u85yUwM5o5g4peV4yFrZP2iQfsE/3kEbZ6gZ
0T7nf0qQOFczw7F0pKhd2s/CNjgePIljCLSS3BaIKwyehoXy0IkX54gMniZo
sBWt9OBBMHIBMJjJS7ZwmPzUCUVlew7GwLLOlBaB53jCF0cDYrG/Cx5Uywfd
XBpCGvIuFlerI1Qv4eh0/o3U7/FbBDqxHROixI6sm180qTGOaXDJeux8Lr8R
8zk/JdwM6h7Bw/+JcXKQythd9xJIVRDeUgh1LpRo7LNvU8gzl1F78T5epn45
Q+bjAA2kFfpoOOf43UiuSGmqodBa7p/+IGPUm6J1fNE0WbZKiHhxRaK42Nw0
Pcuk9j47Dy4wau/yV90LsT7VR8Rxpz2tpVXEOtG6+ADODRotOeEVhULQaNYZ
zPEfUdUh1gogwVgSOlIPgu57KRiH7K6fjX3Il+8f5Wel/LRZ/ZQZ8CwLp6x7
FWsIDTImwX8kKwhHsnoqktDJP6ubEzVyzIiYzQdDwYDgNku+Rpjc9StmmJgX
nEUymXuSOUZx7Esw+fqG5Qo4PF1zTxr5tmgam3WorwIU5JDLkO39xIzhEIop
vCdy4ne6WdYRgbh3tDz8ObVIqsZg7JJSgzrcVYlvjUFDsGFRShlorbIMIyya
ZOD9d3OtSNhjDXzuw2deZmVKDdTpOPISsSjv31+/XFxkWPhiZx1kj1cl8Qr4
dbhMjgfwZ22fBVVZjrNl7q++boRU+KiVZreY3GzNCqJb2ncOYy9Ogu0aS+CR
vgLGTmsTErzZUU19o+htw7Doj6Bi0gUcLuJyTH52U6okxNJkU+ut3j3TyPLr
gL15ytPBrQhgA5yJS/sPQ1EERVlLSIgvfegZme6cKqi/r7JxG13HVBJhFtbL
6tGo//BnOvx8iH1rQJxuPEEL+yBCMZv0tjZT3DVyg3xt3Y2SvxwcCUzC/CFp
hkqXDopIiK3gGRY7OC0GplzxR2Efe3WLxZOXWwiYK8gXBmf6P2wp2BNtmx9u
IXosI5A6eu/zOlsPUQvfU/cNyeXpzACvoH4AbhihKFD8iXUGYx6m9BsYzeU4
V6Azyu/NPCcliB0GnqiU74VFtRh6aT1z42wxEQ7k/KJJwY6pSGu6QjeXsXYm
0da31mqsvXcE4ueTMa773kXV9FTXBtQvDpJnONl3ea0ZOXjiy0GxRC7ZyiVW
eBO9UlqZMsraLiq65FkNlz6kj7rdqSU9dqJZ8W5lkPS16YAVNsEo6smrkUuD
4tgWqr2j865P5AnVGcJ+bafM6QLT0+lerIlaM55O516QKuyQsYvyp9qafQG7
6Rih8bOJvcBF4Ewg6ek7Rvky/b15vwAfUPxCX9sXph8wJXLCSjx+81L9ftQV
tWp+WhaIjsyUUQ0GzYx9MbvR2z9/ZpyJevjOL40sRZOC44+EHPQQhHrLH9Ig
fF5tS3dxk4Tp32gRXicrxwPT5dmb0tC/m2Uh2T0jG2qA5nKZ4e2jqKfhQrNP
bzbCKnNgPewSwMs6Eg6faMZgWRVFq27grQmLzrnh3eL/VX2YLMlGlYNivdef
+WCLeB6i7llq1tYrw+t32PMaOPU3xH3u9/dd099OCxCuacxsEjo6IK+6ZBIW
tmrDETVLI7gpGGIN3gon9XdSfdoPU8UcNinYZhSEugIkxoQw/QHxOP8dJhM+
goCZH563WUhl16vyRgrD19OlSDN+5KEA6/4WwbDM0Tpq+7QwkJxJqJ2zH2mt
7s/8yM7L+1ghzj3uyEWVlKf7xl0RQ40jvdCs5E+nPXNpxxs/FDns9NP2Mm1T
+5pmTXvmzo6n9vk5kj0RMu524vrub78xlBja30Vx0vE0RzZG5x2B4dCHkgcr
aKD9DwB55CVEtoURly0HQqDzkGfaDG1VJDayB5NDUZMisySrKK/mtmjh5rPq
a1d7D/GwfCnnwtIyd97VosXSsmam3tnmyuP2fSmCqOfE16FMpIeoSxdpM/Tg
hIT1a4zvhgGopGV095xfF5EcUrWkgEuedsI/gArBIt6Mo9+Sb+lds/4q0leV
cgp7FFNaFuJ8SDx0wp+oHXbnEY0VtEU2FlnRQvNNC4dC6wplsxFydR9N4L6O
+LBhiF4xWJg6oykrT5J3Kw6sJCf3DQw8A7PZQbM2Cal/2zRgPTv3QdadhMVA
yasCFingPzJW22gwp8M0ZKsU061qiesWwD//aJTsgCdLkEl/F7qUs4FpUwA3
lGowyRN6PRrGePscBQBFfAfc3OAzqKnNbXx2kiM8cm1mdNviNJ0QAjRaParr
du80lsGKgtsylFjjW2TFljvAg16KJ/9H/gVwnAL2CZBeVx83Ud2QlP+gyKRo
syZl/4LA9RbpMkhM9LUCuMzzJGUibDezE9CkJIfMVMQBTsmrVbv8DNPNiEkU
jThjK2dbL2xjhshQ3gdmDwnYMZ+N02eNI7IuZQCUed9F0K4qPTVjn7m1clzs
0cJICpiVRJiATpr/3cIJa0ApXKJRFpVYpmb0OoGN1QYKGEJDBBmu/o3WoIl6
8AVb8WR7R5CuxMAxA+c/iebcYCK6034n/Ajpd2tfxkee4SOLwwYT6IArS4zW
Xf2UN1dF7YBQROm2Zgra0ui6yvfdmxkJf4436fvpGBnNkDWMTxyiVoqHIr3/
9iPztwJS+PWA0DHpulJuHB/koDtWELR9pl7ftKjaYhjF3bnfD6fhsrei45Pp
zCNqPWuvbbOYD8CkD8aJfe3ghW+5sETqvYIxYsP4M2Nv14FK74JXxD7DXzET
5v0A5eq3iIAiLs0v1CWah+kfnLRFVyVQD6GBE4laxUAd/K3ULgEFNjWXWXBp
38elZ2kHClSnce46HgQ1T7hxqW3D89eZlX1e2ThQfWGcX6cE+zXoWCevLluD
Hr8cZlzXHrgB/YJwqy4bvOwGLFnZ+EhS/VT55ZRuCUz25moiZhaECXTnukW6
AsYLqY2DyqRIvmxmx33wCnukVi3s/e7KggNyU6SSPGP9hfH8xperaDEl8Xf9
+sqhElsQWelLUW0S7/NXFjAwZQPFjIkBSUbfcvYX/LT2l3ZjTLzxL1b9pItP
adVbQM+xddQuFjSnL50MpNhdIOHNGaASOcYB+L4h9trOIGS2RPcNojZGdp9H
GIZse8SR3rciE2346bPCVxTHhuLtvmjqi0vLIfwISPMA0IavWrFwRwnuahMU
uvwADMZ9AYBFJtBfD5RcsxfvtALqzvLlJxCUpeZwBaX9x2syOX9/JUjyuR2Q
CWCOpQkhl6eFIE0q4ZjoMhH7aqlhX2mbP6DjX+9BbT8O4u3vDbnJ7ifQY/yx
vkkGYJDXhzvIeb/+KzvPkOz9YPPile/Cy9e/kMvF+rz+rA58G/p5YtKKMnUO
Rha3Y1/zVkZafp5n+MzkodAVq7kWGSA/xYwxAu3s3zrWqYpiQF+lmndwIMGC
WoLwfUQwcF17j7eJ2F05mpCyGGU4GFH8pJ6oM8eZt+wiHa0+T5iImJVDIqgf
cZzRR5OtIrI17eXNuTsiCp4Wg81VkN0Gwloc3aqGcdJFEFXHoMFMbwUacM+p
XzOnBdVdfk1G2detPSe1N6ll2CnplSZ07Cl6iSOK6Dm9T1gHR9R28LTUlHYB
o42UtqW9s38t7orvTvnu+bsznfYp7yW44rrNzVYp/vPiuhO1A0neOuiXqB1o
G+l8RtDY4/wqPwisJRAb46QX3wBOkPDe8b3YuBQFdEwcVqJugaMA9Hn9G+q1
s0nQSqwSL72sH5uI+SCz8qRM8XxdYyWrcnEALGZUGfcZQ0f9JYud/uhqIsc5
IR+Jvie1UnNCHGOkyKcvSAI6P5/pL8Te3OBH1MUnNdgC/zK+bdoiMlMBQz4Z
og4KRH8JK9YRKUXizJH4xPRvCzpOodjqJO6obDJuwatXY8xsvt5O//AkfqzW
BkB7F8oxg6wJo19Zr2x4T/1VavMx9AOi71nrqesHF+r8uJPVlRdqDRKUfda7
+uNsutJyED3lj/KpfYmGSuTbz2Y2byRazqvY9PZ9Pj+lYVSgeiZ1RWyNUTTs
PUmo3ZPpOLc087Uu3MtrXoEY0JIns7FAFTwPjw/cF2oB6AoHToR5l8QmNoFO
9Odk7khwemf+1fOV/u/j6R3ehraP9h90QN0G8fPChGQtxGcS35a6SL1iAA+H
LVPah+tGR9DJGvKD3R/kLFX1FsKCcdUrd8E5mNAjdIl+a1xZEyrcPdYmkaIA
z9azWL8WduPqzEu+Si8Xlhfk2hvWmFA539eNXcA5x9KgZb2VyKaRqmuefa6V
BLg8Si38Sm+Z4lSUfpaX7pstyEZe9PXz+etwmpunm0fh89gF4BfCdGxaPLfX
DvUqOhoqTkRHoFq6Nui2IQ3p5TjkK+hZ0Ght9Xvw91SAeSgJJHxkZYrvMmwy
aFD6BQxBf/saNcj3DpVe6meSO/YgGtmvAH1qsEdRK5AdM2++/AjQ9bepwLaF
vjSjFQJ53EIw0d7i/STm/qIP2Jav3rTt+amzCtomdDAeXiSHzFPs8KIal/sN
YzvquVzXJDP+cj64kxP17r+QcJxAwnJUpLjiIYecWYeLmqngK2UbOOw3Tyd3
ML+A4DJZZopD4da6OLSP1oA2BMU2THJ27ZLN2vyK4D3wbqFd8XBWyczmNmlc
n/SLIkR4AqOP8J9Ov5IIi87Nfn3cZ3eiiS46fBW01tYBrlsODwR5vq6I6WuV
hhTDBJwSXrB65aBSHAQJE+1RqAUpR1OkmwWVRRE0zqlKc7ZoUPvbVvcUrYfW
1NLm5FYELs7DfSl/2lNORBhJPoQ9aYh2pFnBmAKczGD8YM6qSdyCowMT3g71
w0A8J4v3hwOm7HnWuYP1QtvSR+vlJibgUiVUZ88Mc/lYPZgDRdi3XlVpI2/R
yI1D9KzPaHv0CL4qcPPjEmLUPXXMyAJROu4R4a9vyvz79fq3Yyxa9xDEL7+Q
cDDWCRvN5zBtVR+TxRE1+I20U9t+voyFenNByZ83E0vpTWgCSL5EIYXd4xlw
XZsqT0F2/YQ49RE+9131StYRABqlsScrMrHBxOVDeBkSxAypxo3LEZbBmvkx
T06J16NginrV1mNXcOwnjCBCADu+A5QuyuioK4n6GtprQOaAzUt9BnLHfPON
MLRbts2++xAz98a9pp2NHUJhBT+kJzopBfqRhhyc1CECyo7UBK6vk8dSk1JI
lgeNWHBj3gslDMWsFR1lKq4J+KfL2LbPTj3vCh/+PML48LUI3N36akCSPSAv
rK+kf2ElPJG9Ajkg8+XvcykevcoAa2BAreArrO9UQ8psPI7i6M4U2/YteZjR
RWPr8cSEhhbUKY2NU7HI1tQN4T0FxjeKUum2+0Acw35dU1O+B6wuOec31/Qk
n1QUl2NE0qenpvBghXsCzCRlBewJiH2CkS8la8QzDIfo4iqa7QA6U8+P3f0D
eLU+YS/8BfnhDq4oLWWk/d37OH+m0kHUHxt79MW1yBO8JH0Wlr58om3vaFSE
WstmVw/zt4B5a0G9/CqGzk+3EmnaDv+tmZ+l7KqFvJDdpMNyYPte/ClJEu+R
lHWAqfWJmE8/8ffA0jufew/yEsSKJF0LwvqJA/0Jo9Y2bFU75bZMgnKd7wSm
+UU0sHgbE9tDHICT3nJ3A26h8H/yEFZC3TM54I7cY/DqOKQZ3dJf3ouku5P2
54UL/n16TRBqkIwiJGtQRA6iT7inmTe9E7fXCmHSip0cggyH+HfBRYLxl3aD
lCNpXIMsTELX1qBpWkbR2vAeL0R6+lC3BsbbECTlNQAgYVgH2k9QfmyiZcT2
ygIE5lKcvSzpZ4gsf5fHkkt0r6Gn4CxTiXF4+6V+6jEdJQPPUE6+DPXvCCHw
cYdOm6qfKH6rXBUcoaOkREq167ypIQq1kjzleDgtkAzQtGRfUhXPNum4zkg9
0BKRE9o1StiPgsavAWe9e+1ZaQKKiACYAPCoX4DZRXUv1vragL9OYezMTsqU
NPZbzexFZKK4lbvHj/Ho1QOK0AXU3+1PG6tbNlYHifl1gigiKu71xIp2ztLN
DWtwT/W4dZ5pTDdOlwNV9aFd0tp+8Ax0GGuWHNHW1ln7MqI3leV548GzcYw/
u3m/g4qfGViM4Pmobnju3RkygFCD8vnIutfiziW1GdZntwpHofExm7iakb/H
/DKS7YArQ6eFpXmHdv/gv5qzv+Gu2lG1rfxY2C/ywbUKJRNaNTWIzkqy+pUH
+zK3Q7SF8TiZkt1Nk9D0JuimWKIt9IhSQR1hsSpO7gnkJ1ibTD8JvTdxjFwS
G1uqnoE8Dvq8oeGaYzLef7gTAFETUvNmQuo/11/gNumkuzP1j3s9P0mZLy2L
reKLcyD7s9EfGu3rsiSOzvOZOPCiUNAJHWqwECHSiHKSOV6dy+X1OD7fLhpR
t2e+ikhlo2wrmdNsHWTjWHWp4f7vlYdtp5PAcyP7/o3Cq2xjXeDraKe+Patn
ujPYX4zNR0d7FU1WA1i8SToyDGJbEM/aN/c8wenJ6Og4juWOeH4YzBZA3cUM
M46GOu1tWUttfU3G77n729y19lEFFTiyPkSfC9Th0+cAwq/7TqePQ+w/ercS
xXxkFEsVTyPDAB1lgm1qZXhrDdheV0+7tkHVXE8he739MEtp6XNTUMBd6oa7
ztTXtEmZPydoI0qSTn8quFkWGwfWzeXsEl3eQERBhJosk3eu2iSEa2U867c0
0ghW0lk66WJuj1AW8U/u+EvVXpGCmTR9Hd8tosrAAKwJvngeTcGAD20kI9gv
1iUsgtclOYM9ArAM57w5JPtX/gOnm9XBLne8lSi0nDkV35cKcb9byZOy+QcC
kyDA14IgNX+Px8YRg29QHJHD4AqHRvUWH0BMJ9M0ZUWtfB2FsQ2cegsqUgX4
CeKb/UWoT1xagEWq1H6yY9rOniZqMHilBXmyn9CaM32cdvYzKl1rLwFzHXmk
e2c1wCu76nCjt0tLXzqZFFD2NGCCGNs9niw3HFRDlOmrq2wy6vze3MJjYeWA
Q/IFIZkywimKOLmGCwy4HejrqPx/jtI9HSeK7Y++f0IpDPLXNZ6+GDpngXXE
1TeTf2VjxLKw836arIX9H/l+VWXiE2omv763+6fmJOOQ0YeAoWjJ3WRb7S9b
EvSYf9jwCKta0dqrYr0vcRXLSaCgeTQDZDQvXefB7wJUFdHHg1mxa0WOVsuF
JXkypSqFcuw6BNTtEz0AEU7HjUCFZIIKV45gfdezp/VpjyWDIMgIrhzU/Ga2
vqFd+MQRMjj0X8gSwu9Z/EwzELUUl1P0lcanBGuurvGAD5DT9RHpr78CFlG8
rK4LcnIjCiQJml2xxqlX4hy2C/y405WfMGBi52dU+9IvffZuk5TBCAreYwL7
cJBc2mfkhw5I6KyFeECLai6H9Iz2bEIPA0k5qGqntkOsa+kVvn+tKk1aeVwc
wGITDEi06PDlqKKs/ZL3NFZMlHMG1vEmc3WccaZCFLFir5SA9fU/FAM54B7C
Waafs1d46KfoO5bIpcz1A//sAYt9ZSHwbo6n2cPWNdDWX8NMA/FJkgHGgWYk
ObagcsOxTWziwLpff2BoDO1EBxmKhJzM8gkKRGzwhJfWXxBarVzVme53mZXL
TPs8tKBMLR3JHQGFppHn5gbvy9hqTx8+8rxMbgd30YoAIEZ0HiY45plbD54T
9gpAoBLNUQA60+5V8hxsrkS2aiSLW/sZ4oRH6bAevGqDBpHc7SZCzxVnxQCA
uGA4tAlQHVuA7pmgYCD+H/Z55LiTbnGl/4RnrHsacf5Dz0DXE1twDksCIRR9
bbL10KXmD/DOqUF6aV1akBBYZrJZz4acih/V67s/dzOmM04adeX7hpgZvnSM
/3e+lfJzVQmxAWtK8KyrAaHdyqTRePAvmfGxofAGlJaPf/53cIPycN7ZRdOh
FE3N3oeBHX2HkjIkrH2HvMO/zp+CWqf85Or4+XoHOtUcKR94awayoylexg65
Xy4/ChIYguJcJKFq4U4mgoRPEaWbUc0aI7vz1WG2pcLUHZ0hc6Jcz1t04r2i
LlIFF1J+ELUb+F2JI5aI4qbnnSL/PQwlin3gA96bCo/HUxFPOntZHynBuh34
oTZj0kkkKLQAPKfefnK9biGxNDJ6jsnBtYJ+pJyhGLRBfFH9a2Z/19ZdGOVH
dzjA8r9PR8XFxgx59c7Rv/W2MZ7RA5LdnLFjVwWoedxnCn65zdvjWXhEBOSp
JcJ7FPpu6Kl0pnHk2NkXeJxL+trWqcggUvJyQP2/vcqw6ncQH/Oise8t1THr
VnvjR1SrrKMihHBk17hn3sUOGs+dH5xsQKmOQLToNg3avS6czB1tg6g9ACLr
zKseKx1szJYUlzJI+T+dX24RxY+a8/5uKeUb+tucFSxYE/CPaB+Lu45vWjke
1ivvJ7ObiY6FckbBaINFxdPdnbpT9X5C2FIV9ZTOaaAoHaNLSe07dblmRUF6
glDFnG8umimIc6mIqkhw6tSLsNS+OwpidWfqKCJekQfrKZmR2hajQ8ENz41x
ZERmISiWDh1TcZb9O9WN2fwqmoa59fOBzr/FU5OQ6WqLCcL1yTEyxCjaJVHk
QGmjirmUtsLdj2e/oYpordAECcd4WIktAuDy1Ga7WLQD1bQtK+mFO17fBAcK
wAbXJfZAq41F13GGQBZa1C0qd+qYUq4hHkWFeHfj9f0Ty4GW13XmMVKpM6u1
A/+MsilBnuWfME41nNixK2BJaCOpXRfEVvbB3mN9sRtRnxYYhKgizVWAJ5dn
f4jMCTI+XnviSNyLmyRZyU708YWDkS4volTuGyQ+7Z9Hy/4Y9nQiForDrsu6
gb2lKzVTJxBOnsZenCsAVB8Wgze6Gx4fVqzOmDlyXlZ7ykUkw7Enpm9zJWzk
1H68ri/MfX45ERxgI5WkPnY4g0qnFCAC4ys7iMUnYAz7MaMm57wM2bdHSruE
Od4WNMz/3Ezl/xmXk6mSeS0w292VfB9q+U5Mthw5d1VCxqaUhzNn2NT2qiOi
KgX8CFwP2gA/2Z6Y9sEGGw8pCUo07tuWxeY6XJAZH+bseHeR9ThEEIcuH0QY
6bwd9hzHGxtoHkEJdPq0dabCpNdof8SB5EEJ2V3bKKlw7vKn2IznAgQWmK8D
P8T9wl1sWfNbGQ2kCqNbNshfet1IZwKdutQWBLxtTflZDmTk5skloycIRxwW
cjCmt+vzAoIG2r/CvBRTBYFzclIjqnSflBX3MAFDY1V1zrWl27PY+lXPhrYq
vXRichMtjGCruDYGKHNJgZKXG/36tnFlTQSIt0RlavQaKB5zeHfrwJ6OQ28m
ltJNd0d9fdRy/P41wm9EzmIhwN9gNF8qEMdfED0OcwGUtRr1YGEWmyvsXTmj
1lfJUKAWXbsuRlDEKQ2J1aOQZvhNCkRv+3RkMpD80bFS+azKfoi5BM1eebBN
arc63pdMYyhsQXGJq/ZKzr9V9Lb1bwEcII+CWvuSyf77uf/WfBane7fXdkay
PtOPHykdxGaa7kiLxPCvvGMSgajDYkEg4CdmBrf/4Bdd4w6p4ErGuc2GChJb
5DOODVLHs1/2gwEi+/wMi9nUsLS12N0Xm7dstBHddqqgZeJNlskQ6D7o3K5q
f6K4Q9qffNnt6SHN6yz+M0B/m1tBb63PN0EueStaSHFtROEL1Y6BxjFU/Fdm
GSgPu3rSxS8FCPwy78QS1QzGTzZJ7tSGbhTM/MAR/i3dv8cxL6jNdMdPCAK3
ECy3gIIfkasUzXPd6PTjqEHJsJr2Gy1DpUy20QSa3u3+puvls6OBTOw5zZ+3
yewFYZKQG7RlVV/saOenZLFypqM6Hv6pcEejRiCvuR44unTac0dZJGwVx1VG
nYs8hgMvObbzMytVvwelvzGiyVRz9Q2gJtxKPi69rfNuNJMFgdiqU7w3he1h
i7q3sSAIHtI5GWulKgh6zvVMPKggRdQN1HvsdMCoPzIWh6WZgdghx7KrBIbY
s7KUDlcaD2lRZh7x9AGrC9DP2/g2tsSVNZkeU0/tZERHiEXPq4CiAw9ls1Yd
11vwPdS2y427oALq+wAPIckIetinXyZtyjV0uVQ+XiSVxhDR/ZPlKUDnFJ7/
ecya6wPiAzj5azzbJl6Zk+dlHlf69Pqdn73sEPbYkY0LbrLxOqCRCkT/Znb+
z4+ZIzqVvQN1bXfP0W4DzcWONwiCCjsugrbQeyzD/H+wUOROUoaPtpf2z/mg
49Sl35EMjxLJLHs34ljc22Bi2gwOqZZxnp5K0SLZr9WpxlO01pgmqTfbvvJw
A1QL7rLylcFGRqtI71LGRYsuiAD8XdLy/kO3XILvMBRxkT6bK6RIzgkrsvIF
Ze8ShM1rLcZMTxswDLIa6uPU6d9Dt/hxTrBCtdv0ZhU84ZxuGdfHRXR143nu
VGFUtpC2CiTN5GxVW+C6HQSOgxgf1QTllj7n7I4v97KeiQ5PwE+sqcqUVlrk
TYd8LLT4bR4nmst/pCWeHXBo/XH1nay5SANy4I+zOsRAWNEdTz9+9QLAUOYs
y2S8qu5IjKRO3b03jOgcn5mkqKZaOBnrfjBefNT7QjIAjfuRu+eUMWzYTMQU
m9Rkbfni/MIHfYeOuzTZfqvcX2nzE7HKrpZH/bVodTlN7eU/JToBHzuMPfWW
pyHq/v/RuctTZPyhBvK87t3pOHYt/NDZ8NtBQ6JrZtBvnIvIWlz/T4Z+Hvt5
zyoHJI4ZsyjlQClcP9/dAiWEmYa2T3d2gtPxJwg008wXrq8rLxu8zJP+72rI
1GLoFz7AMaO9oFC+oPj7XuZe+tZdy5OCus5SS/jwy+3To7F84MaQNIVC7t9d
0dYQl8QEK/H7iJOkALNN9SF5thOTn8HkPtRn49ohI0zpAe5f0e2gAyOAtIQ+
zZvhR/KCWgqTJ/zqa689zs4YGHSRyFYGbM26KOQjjlMO1tTF7oVBD3oE7jZr
3zoL1CgWz1J409xDkrFdfRKb1A/Pn3Q2RizOvRbx0b3AfD1PNoIt6byylVYA
TUB7HuVbgcQ2BCDsQe3mChLybEsLTXlhTbD1RD8E7VJ5kcDD0GrrA4WUclBM
p/9Qs7r2g7jzpaSpuAovYu0j2qQ+jfB6LhEtqqY9gGCJ+goDG34/+O/MO4WT
6Ktus0fscx+j7ztbntACwQqRcQJY74/IHHsroqRb2fRhwWfGpZElhD3X11Pm
qu1fw7FwMb8lQ/GmgPfnXXIFgAEOi85efChfxajKzvDG1pF6LRopSA3wk6Ig
3AuX+8/uzqpNsoo3QHeE4p7gKcD1NkhTEXdXjYwscVwm3fQZckIIJ2YoIONu
KCy63krfv2IhUZ3rPWwj5qYpJ2rWaxSw7EiH/2/ZUXCnG4lRm5V69fm2NnO9
nOWWTikVgaok+fEHWBzgwSYvmebzRwqdyd4onCKntgdg508PCjypVHyiWwcE
Ds97dmCp32wawGazzjOYHTowzyuiOzqyQe++xoWQJxueAoNTEEYJI7oBPmt9
u96al/XtQVccZu7oJGMx4LYqXS+oAKs4YWRjbYf3BWMBFi9AqoBToGUQAqHO
xvTvJJWLY/einxa55T5Ff3QPfMxmajt6IDEzLSKwS1BH5dtvfB4ZONqHcJTE
6I8FW4v6S8DJBa3DJAZlmmJVo+th7TSbWjosQ2GOsbLXCN/mJ6iXSflPtXfx
UCXlQFCs7jmYljcxFkeLLAOr2BOKvt6nGvEPpfOhu2D2oozRlWrKN32JvVYe
7SFd8tK8zAgWQ8JCFAyuSybAjwBLyPPpUFv9NIcT6gU03eyDR/FnZWCSSRP1
Hnm/792p6wPaCwUJFF/aU22ulNHUezvJBrijVt0FmvOP9/B493CTkxhRvisb
zMeqirdXWyOWvzHUJpfMPNEwyHFTIsyCw+De+svid7L91XYHqXZP64u+KUU6
oser+866IXpC/aGjUZmD/cRPnSKzsVp0oTv1k8ICsloSn+KLKV8yARu6doKT
uCoGVFeLTG15zftbEuaG3VJ1zRX3ElaKnwMFzwHJ02ZDxlemTbtuF1LfnZX0
qc2RlOWUKKBAlZ01ng4Jnf0dHfSNBULqHG0h1dV9Umf2ETky5dagK/AW/4B4
rz61vPsm9FkCTiugZSSiCN6UFq3A2FpNvkad+3OAbHt2hFalwc/zaCf+OA/E
EeI0884dxSH6BYdnfpCTN9rvOxU1c3rrlyz6yUMqcAdYOQ4miF/wR8UjJyw4
SRvvHOdM8gYFq0dH2ZiMgXzoEGDgE3I0VAnxaHgznK4ebRKdllVlNw2inGM8
xtqiWfqY1+x9LgsxQh5LbptK/q4dUHoH3MFlVu4Qz8YtnYMlNx476iOSYxkK
2Wp/DqISkZG3JtMLw/w1Xv5M15R8z1UWUmLPcs3gXDkXG4LT96XyTRzLTog3
e5Xbqa15HI62y7uyC1sFvclckfjqGUbqLL4pdYBoO5l92Jm5mLIYbt71P5Ot
dyJNvSGos1JDMckpd1IvkAnlNzD8rRq/rA+tTMqLsqbpBkbzdZyh49aPbMb5
k+ZLkkGdN441PoMlGoWhSLBXhhlmMoHgQW6DBIh9JKQ73Zsff10Z/2XiPz7e
J3NNYsvdU3evX2hKSAJlJViUpTc6AbzNu2ZqTI83hhf/ENSRDJfgjV/269mH
1E0jkX2jVgFzihEZI9jeNjwLyvtoDvFSk8Xp32EtUvT3Cc07qy7K8mFItyf8
NwzFk/SDZ5qrPTrceyifdctq5l7aqY0NY8rT18a1f3UWZBTyWXHvyFNZI3y/
KLneAUnBcyeAfAKM8OBxScWKIvNm+XDJeqfkQX3Em0V4VM0bYamLtd/ZJHVr
Gq3IHkx8hY95PF8LSCUEJNtovD/XyLzD4jq55I9l0yJRfs6NTb27mj+qSiNE
ebbeNEmMR1KGY15f+6+9P2KG6DcUfyrUePntgfG5H1SDjhiiwXAW17wgojQz
eF/l+f1GJPTPASoCDhYEq8+BnJffnZtltIAVqOkp7Rzi37Cq+bmuZY6ds9nN
rnHnNyBG2niSNNJAF4TyGY5Y479ircVn5WgKNGXWWpMCBqBEhe/QVAkGulDf
s81vgCeBfSYnoFNeFmj4PfLE7M/3qEntJ64J7/wiEeRl1LQCxLPkiRVbwVDQ
dxbWFqtGKXsnK6em49+SRWcS7oHpZBHy822HxaVCSBhhKZ9iTITmDII00bhy
oxzajwcKy1SziiSfiOp4RCiIWhCKVQ3Z5sMv7EdGlH1m5PCJRGAhZfuSaO0D
pFXIjNynEssV7Ax1zt6Jvj3/gJX0kIUOylG1T38OlohqCWszxF3OwSsDswno
gjxRyFyXDUKw04+FsCKQQuLWaKzgmFK6AMFWdtjAkSl24U4+JaM1IGO7Y6dx
yagYjsAyett4dAeUwAcX/1wmN/wkNABGR/IOsqlYuLcM0DfCPdtEYDdYafxg
TJxomQz0ITAM//7mk6qkLH6tdowIS59Hm0dp7J/QSCh4eQWvHBH5UW7/SMQP
IFS3xlA1EySrj7h/aPBp0aGKYPzuQW1Kl9t3gsqcfkmoIYcFBumk3J/n81CV
n66SvWn9eivi+6o7+7VxL/mwjMmpMF7PWTRrwuXDdVxmv7jb9ZROgh03X3Aa
+JJDcK17sFNWwCuuZvSKxMRrVfNrYF88bYjt73teBDR9I6gBSAjwdncmh1ub
uJkuMxWEz3jRF5z7tjd2AbOC/j5j4vRJLIp1liCFBKN6VtDKvs4yrrj82py4
7PqezryeIheAjOxC5Iz/AzZ/3bMMsd2Kh+nAExNhpkN4N4GjeGOPUYEdJFKT
UxLTKrsJUEeN7bo7Ej1sp12I6IwpSEsTOhOc1xup0vRBZvWinkwMtzhtc9Ya
yDy8nLRpRob/v/6TrIq8hg33wuICE5CPQkV5WohG09oVvwsUZLJ0WRPNdQ6s
Db46sUTEDfEHVH66X+V4uRcOdwfjRoxJHwwqounUGRgEkp0THap7uH9i3/wX
awA/CEDSI6qtzzefUkcesfT6Qg1LGlkw1yco60H8JnxhmSElopZe6Fu2c+nO
7CDY5pkn2kW8FljE8fEEhRzygjuftPSEQYdO+P5oprHDyxCugemuDy7OLHDo
km8Fne2VQ5wChz6+dW2p00MDUa78HpJSO8/9u2vAgBDPg1zfPJkg4LkaXsK0
u/vwLYRj8Sz/trScRlhOrTwb4QiREUXNjL6qKztyMcjSaftQSI1PueaeNnIo
u9vkki45s7jYoTBO+iZJGYaqlYiSxC5UHFIt30ElzHf0I0GMBL6JkqHS1GgS
91ULE7yz7Ciw+LhzW7Uw9neihU7oqr4xO7TBtYqf7TvikqZssQ3xYzB1RXhj
rE99QHs+SpMOZDOINT+sqT4mZVEqTjypMNopAeRMr1g8A96Y6TF5FTi4w0fs
Ff/NVhGCJ5ET3q9UoI1Dhn0orVVRUC3458KGL9theHJdIYMAVRysimpT8kWz
O8KQu2Mm0Mo2Z7ugnVSQRt22QLSpuD9FvXq0oqQW4fO5V3niNjNhqFH9p45F
S9dURKeB5STIUFAif/AfQR0gCGEpuKzCBJmHeswtwjNCs8e1UB3l1WLwzl6w
3a/tZFeNAhns47ALI+/gz+s2em2d1PmXBUPwU7PYigmJ4SceJRDZOZnzuYkP
yVhFqLsOc6qW7hSu4Qn0PAgQP652rLQ2L1GpnQCT3eZDiYD7gi5WkkKQtQWW
inmhr4JfhcPhahH5e9K4SeMIAIZTDTqvOztYQ0izJfHW5xs9SNm9tJ+zUgTF
QYS9GGKiLAU3oKv+2SWX6HuEODHg0a4PqGntvFTdh/qF16IWjJgsLILpgJsF
LXhWNEwWxKhwGKOvvpqZSf+Is6mfM60dbGEALduChEnqoanPzDQfUbFHccvG
ggvOdM3yzh9555H3M7y+N49dGE61BM2HcZ2pCIwPReh8bEukdWfXPCVmrFBj
OQMIKd7NCPrzWV/1Hp30VJm8L0l8mZtfjK0qG8sVKYuOjvtQhb+k7QkO4Tc8
H9W0V/SqRNzPwsUQXultUHLQpqHSVfxfC7D8Y1gjlnKy3AjVPehGZdIZeMFf
01+DpSIbShHI3qSCZFmEi7GWIHIaTZfI7beg0TkrAChhJjSmB3omqInUjz/v
VGgIE0OOcyKiIed2rOMYR6AeRruJzBKiRgdKKKLDsvY4AOPzyLhIdwIynkA4
hbog4imkAnQw6Bo9wK01S/gFEmUYfGMH6SUthvMKV2Miy2HK+gzPQw5/wnct
sLF3BrlcMbUyIy8CK1OxDyeiNm1zkBgVV8Ye2CqUv0h4ULkcpfqkdFmSsehS
MJkawjc431RomIQfGV/Jl5esvO4Jdr7q7h1UFy5+2zsg+0msXrJvk8xMA5ow
zOby++UmV7x7FA6cQPOgX+EeCV8jl1iXgsmJy0zw4H8JDj5XOSiP1/aihxJl
v+D5IiXAPmR+AGGAH/sXI2TwP2qV9o2p9Qf6ufmK9Alu8aBOD6rJVUCy6Djk
ZGJ3F5y/gooWr0XKm6NUK4iSmQ58zxp7OWkWcj2v+WxA3dNzSIIRiIESIMV6
JUhG/0u41vrINUVM51WH8W9c5cR2YT7908XXLJZpVjiv40/7st2wTG/YIf8u
Yd1umO9+jlvzVF2cc8C0sjpUxfB1/DEHTiMXGzJGfcAPaGjuEVVOQzGvtOQU
e3+vSAcWnN4q87+9x6LmjWuT0F6LuKKErH4wq6YnO7cUuszvkCMerAINN6pF
6TD9K6r/krw0WQjEg+tuLGJDPRT91QWtlE/iM/wN7OQWn/QsTULUrpTEMHwg
7StpFHATmH8OEaDPjbYCRBxPW2mDm+YAzexkqpFEOny+OTHW5NBv3x6991gm
HlrESQqC/gdYjRbR+73WVF4xa22c2yxZdcYiiJ/1f3YVpdKRfBlfxHYENrQh
a2AxX4NxScvBibdTt5h3EMP+e5IJklBoO7/zXX95xLySSIyhHhavLOtPnvC2
uW950gLSnLktFE7OYulH44FWxhLCJUCeEQjsKmWVXavZfY3RjvZkAVRQP3Kj
eTLMzb4o1Vw0pesXDX/2k/NpZl6GZIwMf75NiGgvolBPF9R/39DZFr1kToVq
bM1NsVFWgppWmuYG5dOzCrQX63SFIMW/m0dxNL1o3VpBAKVECsxpGhmegk89
XaIGiLDo7e2zCFp7QBKu27aZBn9EVjp3RAOgbiapZ70e/GNayXBTu+t9OwvS
1tYNPGnzEuVcCqPqljHuvyQQLe0gpffFJP/NksNB+GLAFupqjmNVBudsxMDj
Qz/SuADK0QBERCb0nvpzeDE7KFWTGJbjA4BPIkvMDvq9iaZdU6pVhOS+Acuh
b5favWOacy71gly0WObct/itVgLTB6eKiNo3ZISe2RUp0XcdQ7u7Li0U8MnD
QHV0/U30L6IOcTBULGAEMB+mK4KA5GWP1KrymCqfAz5Hhv62eF4IrBQzaOu+
iwm/fgeZJHFb58gB7bNv672+ujPMQfJ1w8SWu7P8IxVObYLwqYy22T/w1TmN
fJ0nbUJh1YqJ+zTOyWozJqv8faU9Ad13hLnO8P1RNJdXfWkV+Gi/p0pg6Bbp
MjdmweramOL1RFmYzQl4pU1sBqnwJMYk0lBlo5AMdagdJ1KwoiT486xzamCS
bUFlZbybMfJDo6M+Bm31JgUaCMP90U9YnEIFbjxgLHw73+hBo8lxQoN+GM/O
s2LDzWXD7+NQj5dlFFX55pwGHH9SfxA0CxfMaA4hK6/YI6UXvfQpN4ztalIN
UX6fwxrkyrwbc5q/YE4iWzh8YIVztnJvvKGliasf56prpEWwVzj3GmB/ek2H
fzXmU6QnH7W7xvNrNyD/z6JRJpow6u/hnexNPZV46Bl2k3Y29u95GTCtoQE8
pT9SywCue+9XwppIZjd+4zunUtaHP5KhI7kiez+YgSVxKhXvHDeV4q8y3RJB
A09Zh0mZuD/MkI6++YQDnvsCNONj0/0UuFG9thGH0jgFWVVLeV0+ovTLDHz5
2zys3EuQwzgXlNBU/kzx46tWTFrATQSNqnIeZCJTYIDBzVYEs1jpSR/Kx4bt
uydFXrZLtI+lZOdsE8LFgg6+fEPnKkeWrHfjNm7ucQRsdcZAsoJRwXaTifTp
zo0ems32l/ZgY0EP5PruozyWNXZwk2XsYoi8rT+cnwiF+MSlBrlZ9jc6PKSQ
H6FF9xQuYcUXVC8RQKataofD8qB6KLY5zUn8feZlTHAljkQFmznGKW5RTdMs
25kdzFgwqCu2ez6iCe0cexjZ8EwC04F9UaWCqy3hXKaBYa6MFHBFtUzsD/it
agS7xjIxfqAJCkQhS9H1wfwDYY9JL9Ac7BmCaOz0xzCVa6yIYMzyf9dN+jLz
+gwYb4dw6VLd/g66qTJ4I12JTRDF2XmEKYgN3umQuh2vlFxDfabf3NCzW/2+
4M8ogpIHHt0VprdgoKPn62qVpCD9teSBhzx96PE1CK8XPeqqSdOiKbqxCjfx
uT/znY1fRjfvvKf0gybO6NPsRhwga9jEKzs2xtOmDuwfRszatM/f5vrWjJUg
tstc0L7mFxSvr/BzoknQyVnUNKEs8YWQvMR0Q8RR6l0AfKy0rtJFbvaHCRkI
LvBuIG/OceIEdXbtVsn1kHjGgZ8WYIwHMkf6vpJjGXqjBNuF3qTwHuUXTZN9
kZXfwxmnAHwER/NCNkYaOrsYdIE2TKnQmEgVmkiZnpYQxaGGmB8RskhBE0ff
UzhcKXb2XBeJRVttIRqanZmH0pQMWc55Xp2fVu9rdePwLsNRZyrSv3mfY7Iu
MUQOIBIt344QVdRcbtF6UvNzcQB/VZhmZIrWMYt7181i8fHozKx/Qdf6uQFt
stdm3X9F8hymyeS8V0xOmBuW5hpOpJmAnrY46IXzDruXeX3zS/+QTZOyYSsy
mv6wdZfqCj+9EL7PTf7d38Sd+wOf0rfKnQYYlghzwFpQHqQMHVkx+8Yzb89d
3P9e5sB/jYBDk/6iS52hmOI+38I2G6gNXI7uYRG7g6spDSNyp0ZxnbuIObAM
FydRvv07k3TjyugumZtcyzGdptY/vqSNKYLd/BVyoM3elJXD8ACoZOTDBQnU
jnUszUk/CmJeBEq3rBbnB9DhbwNUEPMklosQD6OIt09trZBt5fticRE3nZP8
zLywyeFaYT2rd92r2x8ZwUZXRoRXCy9iWxtd+5WcnJjHDg/yKZDGC2LUbqDB
yyAlrH+MthyLOgAZKhBir758Kf9bFNRUjEsAjNbz5J38fmBnD/KqRiFA9cpA
6WaEZrJY4zACZvG9ejbyTvRKUnScdH+wc+1c8vNALccPWe6wwnc28Nfkhned
kMduOjC/B4DtfDgILLbMbCfGSKqLiTAAtAH7JkwMMsjv6uQX3pDz0vP48XD4
nrGAiBxrVpgaOdO8iruWOVJmucxo6mJwqlaOIhFlqnpVegHUh0ilQ9nttxjt
uZQ+bl6+SIi5yatrekGoF1jt5kFi7/yWUmxDEGLjex4hb1IfLYuBMBgvMkCh
bESbgfE8cFWgYLfTRsskVGppb7U0gKikuZHP40mU1D41FVXUafY7ATJpr3qY
P/PImjG0ES9Lzs0fAOnpgi78V/LQBjAPHoz1Xxz/iQzZqE+njkF8U4c3jFv/
eXAAyI19TFZDUGB8dzU2crszH35mwWSQnBKYwT+F7trEU7yFG/Bzxxaynay5
ztfh8Z6H8BGs229POPwFt3geurxy3hj2i8pqudz6bRDtxM9W/MWjf3YvgRSX
BpMpmhjiDXzjqcsO0+2AzICjiYN1huGJgXHq9jj6foW1W9msNQfJcHXqD/QC
d2UE/sx0Y5f51uvGYVkXtA6V9xj1vntLVcGFgRUWZYgQloC+7oqb5Z5OHG3N
naYeYnzL+v+cbacpxugaEso5wz1wfBoxzi21XD+e8FAWiWqTynRBo3o+1c/N
+apZYL8R5WmwhUhNfNrViqT3BwPtmO76iwWukeIDWmGR/xf249lxIFTLms2l
IxftEf9dx7gpSmUR6EEQWkoSWyZB0F/pAEmsTiiafj+ErUt5novrI1qFpWtA
2T/7L6HyxqnYimgB4SOkg6KoO2WXc/WW3d4YyNP/PRJpLSpPMjvl0wTIQ2ff
kZed9dFBPRiW2tEUTa58aZ4lVErhtjgaldu5xA3Uk97L5ZDrwpMnJhwZV19s
4bxf+ZmxLzy4osGW0PGW+fD654yRQbFowk1THxxl6bGciQP/VXXXkT3vKDMF
lt6gvwfV0hJvULJ6jScQ42xSO5qEV+CE8Y/snnTWc8rbyX7QRnTvoytOIxyS
6KYZwTGWB7ZtQB8ILMRy+XTGmfd5oj+PKpsJ279PDW5LPVJ3d+P/E68YGMKH
v0LHyimjlaqWl8AjMVEooJRtGcHo9Xl5BRCO8bOSGbDufmC/mjxS6CLHQcVo
iQjrIS74VhqegJ/yBQT3s5t6eNrN0m+qZ76+lc4bobmfGGU640EtcvuCiuCo
QD+rikMX8VdHctUPW5cC2O7gK/UDHBA5OlzUH16T640XYyJzxy3il7De8dWJ
mZAqudJ9FoMCAQLWbSrGDLE8R37FPT8ExFPtKAINjA6BbbJTGs1fEGwaCTLY
PGugOZE8Ef0jgzgQ0S/P/SmEMqO5QyIg/Xdb46sx0tfcxB4ZDw+zFxXgCisx
7+pXkISnbqT4s2iZcWbB3G5FO0dU9tkM4l8rfxB8sASp7ursV5nUXjS+qu5A
w7gWfWmI9+NiD+fAfxME3RhqZuiiP78NA8X1UhDH84V5Md88TNL9RPVPvOc7
X92I70XgL46iJkY7nN4aE+SrAZtYwBZNglBgDuMBjE+lLzhxwrvELmD3xrjN
hH91ELcKPsULCQcvzudg6daBqTfZLl8bA2WOpJg/nx6U51skCegbs1x3b3SX
b/Rdo2Wg9Iv6sBfzslsKLjpX9hq2Py1q6uNuPIS//8rWVeJKL7letlY3zMe6
2e8pfKzl8txIDE6F0H7uXY+NXaFxXC2UnMFAULrfLIleF3VsMBfOErKvmSHg
5x6tcSNBYl0b+wWRNyBAVrXhHJJ1rfCLyt8YaVv2WONpA+mdnI/4Dr9M0ARg
5wpCqFsmItzyaMl1d33fb6/wYXMkCdxKG1vd5JYAB0R5lv8d4UTaEoRQxlty
R/Hfy/rfnK3Ks4lzPL7B8f+8W4RD7rXmn/kGV0LTM2V+EZgYaDKLn/z5ExMZ
EqqxgbD591qreOrB/BA5fa/ryx9ymjxKX5bRvxXlngEFNgcTT7WGALE062ht
RibgDs+aXbfKQesDeAKmD3iNNvoKbXBkeYVyHmFY3FC39bxTCxPHe8obq73U
WY+c+hBViWKSYpmTLGSdNxdu/9p76eVEZudgw9LPZzDJWWlWlJMkShYO/Tbx
pM44tsxJcG2k0PZgzGjmzrXVrxC0rk8xVoNIZ3dCRCelksOKJszNpwvemSbR
eivXkT7otm2/P67LfquwnY9OucKHPeXirAHj2n19c8qxshoOwbeFtKjPS1bQ
UPwq2+HTV210VBNVN/eOekoKMCQijaVyQVnnL3/8/sZeZpRxaq6gRqy2Z6KB
/AxIbhey1eEzzLODoxdu+Zg9DlhE4sYXH70cKPWKWVj+InnWmFuP2Li3DSQm
nsztoM7y/nyEZz9ZhAxrpP87gNRVn21sK27OyRzBwUXnZ7Tn3x1chlhhl9B+
k99QacloyOaMSnRg6AFkQ1nKwBpIm2IrSK/2eWeUiZPTK/1k4vdDROPByI0L
5JRqn8ppu90rPqa4k2kR1RWaBkiG4KpcQZp4OCQF2wEEO1BHNMYRB8HwehlB
kXds3x59lTH4iC7aBNy6ZYS4MYOkWBumkhY/26STTVlEmA2uPiHkAtskD40z
F7cvFZwU8QbOiSTbA8SZMum6kGejmehPd5R72UhMTGuctlBMS/6POj0QmdZk
pD/jHoEaiS/MdzsgXvWgPqRVOghmLj8YatK4B3fEYgKUFKq64nW1RaGfrMpc
bmXmR6FXuS1cBFXGs9fgeFTckkUqTTnx2153RRvTU/XseYA2JGCX57gmzptA
N81mKKUyrnP+cu8kYXoW1sur14P4YEmnFofwElvVnvr9tbgw7MQgIv6fWw/y
Opyh6sc6245ycUDf+UQKYKmgdCyo4QyCY2/w6aMKgwVeOcaHAA1MsNeScD+m
shQ+QFg2ZnyW/FHqguZKA2jGpPwpwo4J6KtcVUsYjHRQuu2O0lBq+CnvP2cl
5TZ5emhqz2kSLB7CICj0rQRUrrAFHyaEy7n4nVUznSv6/JJpC4+jEWMnUSft
GgME1Yzf3Ol1ZXVz3bpAzag571uZCcUeUGR6os2mur7B+FQE/5Ha/EsHHA9a
Oj5scog0Pfti6mPYrL6wFZ9IpaOOJyPNUjUXhwBCjZx7pGkvbnxQtbQxj6o/
XMbutwcwYfSjGPEF1Evz14S3V2lAgV9Fp8UXpcq5MYFHryvut81Ff6l3Vd/A
7D6FScrYMdCxcu6fZie6SnJouB4fkxXdmS0P+zuB7Kpnc2sSL31JVmXM19kS
jVBmrYS6k7qHI/Ja7dJ3SJMcCdtYl5wy4xsi7xGSpk+zjZtY+Ak73eVj9BSL
twqOFhwPXdLiue5YSBEqW1n57xFx2GNmPtxR8t25xTdO2BZpQ4uhTrsMl9yJ
yU+MypgcLpfWixRPkWaw+59vnXBNTdea7Dfo672UruzNoAGHOUBuxbAOVVI2
CnGBVWt5Wa5Dapv9vngVFLNhp2OPo8fCwiXNafIxBA55BjUr4mx00eeaQIq6
6GubVKHbYGXzxRaewlkFkBmNGy+YgMTE/gHX49XmgSoA7QjrNmNmPJ+adB2j
sqgbq4Aak9ZOuSEhiJFFqVhogeO+M1V3GAy4e0mns/dcJ51+2J5pxsjMf2fa
lYgjWWsyIaaefILaTWSdz6E1cCU712W+EMbTOGQ9GNeoDe9s6H620iZtmhUc
yNZ/HhmNjt+fnoU1TutzG+ROZcuP6U2OLegsbsrqPPI9kg46JODcqTfLDK5b
qAdJln+w0WmaYZSa2XEFrkwKWCCWv/UEwXnaYICRid03M4K+tViV1PfxtT8I
sreIUSZ0GPNFbnGuGAVjtncsIAjjdnGlCeUftj4Iu9YAKv3yIL5Q4hepG1UF
nQMigJVsIXTm8htFyySvyOODiXYqONvx9S8IlmhmMNQrIdYKmtVZdhC/1zf3
NG8DJ/mP6N+1Hkp/+hMP3g/Bc2eCRyGDf3WpcQheCIoa0C3bMbEJFQUbqXX4
tGUjS9DN9WE/PO7Q2y8xOhfXv14zb/jWasQ+LcuAeg8evUje8iCAHPkk3/wb
/ag2hDer4xlf4ea3o1EzbQDhXlyZwplfByuWw0yZZly5qAnp9fYZmn7S7+AI
6VMelt13m6Fli6Kkk2j12m7t26ZnT6+q2KwwcQLgiyCeVsA1Ub6ViXBXb0kM
ybYJIlnevABZE5qDp7bb5C47ifbjROojCl1n++nYGudpGW91k2iXh2hM3t9Q
qJxeQB9v4Po1+J/gO+6JUTmyRik0c4ZCVO+GgXodGZtnePYN2CBGf2E8XEWn
PQBEwyFgKQWUJMGNWJ0T+/2It9P2l3x3Wm6y8N9zImFzzDK1kEZrxyhS20kb
0rNQnCLdxyUQxkcY99SI/EGcm4jMLEfW3p5rDs+6S5Ah1ipMQRnIymTLpEJh
6WYfdkAPa+nkeZxgzOJQsWiMgEjTEmTknaY8zXz8Obb5CWjWHiznxf/5q1SR
EmYfdwCyfnAX951Hy9Rq44/bU9BveZY+WDSlkzVGt9UlWr+wAzYYEIpUa9AM
YOHSvBJJetpskkE/gnk7TETxt7yNx75GJ3tgJ2/oSH/r4UJGz/arbAYKtzYH
ShxD+y/KE1kCQ2R2RD1NvkePcz9h/bi+GhqFtIE9Fl/avqz5x6jYsoQDPi1o
GEiLXDabUNV4pu8Xb7DRyN5Ifs4blXREfFoWLsJKLVU1/4nnr7BPq//C00E9
GkZbdXdRQ1StfEf/q322j55W1wX2GOYFC9teigKsScVSHKcJmpqey+eUgoZl
Ro7tCAv3YZn3Rzo/BoZDOVAY1HnCAtvTInejAQ58bwfItzGf/AnY2jKOdwFl
v6gzBgn8ldNxpVsw/Q6w6KuOURhrY2VPNTDqvBpY/eLboadWtilBU5oGrtmV
EAvUUkY8sLNHfxh0e2rKTQJSJV4auIHFoLn7GwBZXGxAhthcbw3nyOOAKNCs
tRpiGioOSBwKCE8wSmlqmm6UUZHkVFll04XZdPMTFSi1lkxJpNBIBcOpHIIh
yKGrgyafMZ7WMJltgYolDxoWEfsjXFK5kpcdX7ve9ffKH+zeWfdTPkb23CdR
C1YyF47i332pN24SF4Zi9cRzQj4nKN+LPOye5HwOrxpjnQ0Gkj8iFVnhTISB
Fl8Mob0fDJ+XocLSsoWZxblTZ8Ezr/HEYFrr/kRUsIW3YgCcyIoKTBaCLo5K
ApAGaRznqjgD1j6/tteYh7uk+G9a3EDQ+olC6kaojt66wC9nvTmyWCii+VSu
Ub0YJtGt/qCcQsm8OMwAJv1rm1NerdVAI8cV4f/q/hJdoT2YaNJHiTWev/8s
dvJE/1mlsYCZwovB9kErSMCrbBNk+F0OZcVEUmxX0x55JCagd+r09qezI0iR
npe+9sIK4q1m24CEpAAnxjbZfDg39HMYcppkrYO2zsDM0KSXAqvbaocm3/wn
bOfsHe6IKQAQ9PaHDCQEWZclwmq16jOiYypoTriyPxITU0diSqwTofFN6P5K
BZ+umce39wV6lTl+kQhE+0vyqJwxsc8NhG3kAG3BP9JkMVpFzuOqFp+ISJtB
1moItCcJYcu1TcDa/UuksthPYeb3Qj7zCPk+/YpkK1+1VybfUPEyfL1xMAQv
v5FCXYGhNp7tQJdhuxCliunGY3dwwGRrv10XV282+UepTGbkFdqdVW01U3B5
hnL9PIz52XX4Kr8aB0hsrPz4Rnp+TazmmPHAL1aiDHTXGALtZ4QK60MuG+Tv
Zr0Qsvx+/SQBHjMd9dS8VRwPLo3YDxwdbh5DPJmLIx7YnoOIykpORK9esyRJ
PYJ11IEX73cuXIyRQEA2VpXKg3NZMP4i4NAwUGcSPCaEdf/eBlDQLMujVuf/
yAlLjYba/mM/6b6mZ75BiEHbkFqQKagL7tSIR8pb1NATYHbvfwUkyoXdBiMt
s9bF4idLBGdcvMSIJbN0rbUAh025+yDMl2eEAeSEEiZh25GCTyumdV6Dsdgk
AJVAMPmu78izeK4GQi06BTNCUbG2CymK+cvpJtmkukqyJKppM2wdJGOF+9aJ
pn/uDacq23XxgyHJxom3ehpDouGgznYPdVwcEBWtqUgrvOU/zVNw+fkwhqk4
nLz9147/HQkGJI6Z0zT8WqmYJMeTpthD/HgMfUwZzdGOe52pWptK4/FXFfkH
qh1sCOJL1IEinRakYEfN90dwEyGZscXq9VaoChCqfXBnfxkdinjrxt/fxF40
3IaaeQDxTIBDq7Eh3TMun6RKYfcyHqgA1ssyFHHk6bRg4GBy7kCtxEoqdnEb
7DfHHXJWAFD3ZfDKHnzByuD9c+gn5whWW1w/GGFuzopV5wKG0w+DlYAK0e77
xXWykW91B/v8yOrEqehZi/JT4N6pDtMBUzeEKzn2Jzyfai0ugYxzgQeMqlnh
l88ggWnQQgkgJ4eL4Yyer6kj1Pj6TbPWqxIKXPwIRZdGDAImJYhFD6UqoW5p
riPIHbLKE44KbKdPHZLy0+RJ2vB5kpydfJoFUPlr9pY/mQwn1DZLQGTeTH82
3BorkBh5eU2bbFuFsA+2fzaduUXVeaqmyAjEBEumTGUC5XegfGw0IF59gdZv
89rJ2tbVKTqgXsZi2uwgi8GKxi3l6cvP7jLajWBHgVzza9/sjRuSI2PsHb0a
Rba6w1wamEImCGThseLgmV3e6XQ0YeDq6I6Jmix5TVa96Xbum3/bcb0eUo7m
+LEVakafhuIWCxE13JD6e1FIdGNlGK2jfc7tKS/xqmjqlOf8yR8GfH21bM4y
Uorp2HJn5SSMCWLK5DiqGrn9xn9JyFojdXr94ZAZaNTK2hWxUQKqJb737+FS
zpHGIvW00eVOX/0L4NJZqDD3AhK7Foa5gfd0ojuZrcgiSJku7ebB8KkS36pb
XoUJ+LUWSvTGKzJ8zMlGz6XiflCSrP4rZXKsWJ507ErH/2mqkQlge6GpxK9P
Kd1kzJ+Zn1aKDcyDUzdEUsALShoxpuPinWrqyuFYX2fPA7G3gA+8srWghmuT
pwEzyIVUV9tTt3GCrQIV0snuRpbjbD8BmdubSoRkhiD/AYJQsksF3nw3fIrI
lFF598qLGqQtntjIN+rNk+UXXgrP1kzWJlpXfkAaLV0GsGZxrakGSX6IIYHS
4VsAETEhppB9QYcAc/UzM9FElQw4Gk/qgm4RKWy7vIZCHrVRTqTcICLjf06m
5QaNfGho9kgwwbDbGmwuoWByyrwkQ6Ooww6WZ7b7UZY+WDLYRAzNi05rq8ZR
Xy7FY/Qj2R9J8CfTY+HKYIjZtGU8bJMLuClE8DExkyVcFqopR1N+hhDw23NY
/OF+nRjbMJC8lfH648gg2dWp016eiad4nnqgDeKCLitfd9wcAQAYq6CL/K9D
gwGly+5nJGs/gzUrNXeLv9GS1EqLSOLAbxQJMVa1O/crdb45EC98nEhtGVJH
mAuCaTuxGXUAb37lx9DvWYQOyp1hj9xB1bXdjZ2OQ0v6v2pEGHIdowiFhDgQ
EGvHBk5l05oda46fZ2+SEs6nq33C30cq6JcOUkymtL/25XtH+J+rT2eClfT3
/wmdY+kwXn/cN/q8GAErvSjgz48usTJque6EyJ7JDzzJYHbUqBbZRMFJ+OIc
U8DCPd/6IfzSz1Dw1AtoLFaHHkzXCiyLRukHm0G0HseReizq+Uc4d20MlNzR
ZLTjLqbauu7eQBS4Qa4CWxO4RUX0kR8eLB/b9AXSX3Z3bxM40N6nbF/y3EWK
VArlU3C5bzWxSICZTRZYTwcfj8Yyk80wSXQV7Z3pQZkIVmqbiAl0LK7IP8F0
yJ9REqpRgpJlyvMMGL/eH/6QEkD332kHhLHSwByE3XmqNdpCb/VT1FtJtTx0
YQSQXJgFA3tv47O8yRuhfdDjFN0pfKhKRxC3Dg42LiylCB3BPPOm6t8EE3tB
3XgHppLalWrALPgAimbJJQKU0Z9HnkrfSRqG6ZYAj7Acoqw0l7udF3U4n9Xm
z4uzf7/8MP2F51jiBYODpSpPLQ5pPpynLm359zh/aMI7xRtiOK1PAhhaC3lK
tHCxu17tdi80Lf1RJprwwX440xwCYsd1821gpabhzd6ovIzITvdBL6tfmEWE
csGxWbDMoauzd9uwe6odToFMk0SZHo0eutg0zpodbGZhKTWiULMzgkb+r77n
0PkwLUk9BylmgnRD7nrQDUtrlZ+7yUrBFVSya/tIIsgU3SSPKrM5w/hP+ffA
0lyqNYr1m9zFLgPFwPqJKlDd56DQR4UmKIK7IAOnHVyBZ6s8WrOXK7CM6TfN
O+iPgCpga/dd7505v8rcme/k8iRaK6gbRCccsZ9TBEipH87qGoQubmx11ZgC
e3bo13FRsZRpgzqRKXYIUkU+LVze6CHFhBXkdmevsaFdcRiEyk1LAortjyXV
75ZhDofs8iC/+uQU4xqEvZC1xpKbIh+xJJB48hWnZpLYQsF0Q5vT5Bl9i2QY
eLp4Ehl66m8ZtIQ1NckkXwi9lQofU8uWb1Gxxp6VWRE8/L9qXK5IwSkVqovD
rErdxawHSeP8Ip7VKyfxyX0rPSF4KuCmmUtkGKiXhH8Ei6EOU86Oo5gi26nl
lsECg0r0vxbiDa9g3QrKQ99pZjjLj1IX9VHrE04jeY9TmmvPnBdQAkvJlJKr
R5fvQ60CBdGxmyo3xgIarQfuq6J18AMKAQvixhQ8trfihy+DkKo1HnGmlole
EQ+C5JhnY4zzicv1lrWCNKwJRZQBoHwgyP/4wzIm6zsOXnv2V48xWkcZhRz2
N33nZ0fHAk0v6MtCnv/9dU+JIuDy92YQXJw7aOP24O/ushAT5zQdHcvLEl46
+sNebmDQMcUkTSh7cJLAber1t7xHPc0GS6xK39jrCWBliem+ocml8CGGLXGk
jskojoOuk2X17h++WyCWPSuMGkyIJv65hgyiGP4hDjVmIh1c6+fZEB33wKID
37R45Pmqzr0WwHU/gbw/Eh5dHDt66GEVybgyIPYKlk65jThkw7ZUrWW7ynju
Yet6r8A4fvyQcWUGiv19o2d1Jl4suP11Qqv4+NtS701zk/oJRYdVu/2vhWhz
vIGrmpYooXHoT7N2Ypa0dV6ojCEMc3oB4DcAhSc5aAgRWooQXKlT547qVZmq
9qIg1LrTCRg9BtrnpfaR8JTEOjUVdDNtIfx2qpGV7KJ2BvoqdobRXPnUQIk/
6Y2TyKKpEjNZh+f+1Yn+3ce4bWxBkxZaa/f0Wf4uxRqBYrSWARFV1eQCmMop
ieDTp/2kN7InBdRZ+EtaTdRYrHRUDi2qAG0uPchfnPP2LndJgYVIETZJOzr5
iPlI2/zqPMtUaRH/baqtdetKLwoCDezw0ScZc/dZJewOgAF3U8gvNKyRn0rD
oue/rds3eQmAJDEq1a9YyjYUxdJBq8bRJ1Xexeqr+4jTOOcyhmqEPg1glKJI
5JCTRrPGvcDytKuDnc3HBDNmEZLkn8TzK0P0uBW7YPOOQi2v/2yiGf46+n1W
SDQr+Gm3TTSQhK+582LjFEAy0OFvgqfQe9FiDEAYDm95gwoHhy29jktprgH2
tAovTSh2Ae6pefEJVKshNhh846+8pOokoAsyfcWILk3Hi2oeFoahbZ6AFB+m
X3otdmcq+G6HDpnfQnEacDgVT0EFzbt2tdMtliRriC+y50WlQiu2tch7gFGr
63NKGwhhdxIfxgiMZbWkyowXTpibaOCuALMmxPJU+kFX9qGv5sixi05kb/j5
sJwld+4gPCY3tEil8eozEDh0jiq2LJjGK50LDyKJd6uO9Z83qisoqW5jWATj
a8Ufaj3LYJPhBP56G8PH7TvxRBKqqo4kr9H2bsF6ctylPOsuvyL1qQnv39lz
pt6y0gh4aFakZSQg2C6V0sNtCJshVHSRKuxShpSRZC/PvraFMlsKDiT7yN/0
UF2Z5vSmBfexeul54ndAOmw0zN6nwbPv53auTpXccqbnR9kFFslWknBQJvtN
XFyq3pKsHa7mLNHfc1xenbnazC5WqEKmk2+w0twsqONpNx9TJ0Y84gnGBfK+
HluJTn6b6JqiOSCN938fXnQ/6K+ILQlH3G4VH/j9B9WE/3ZqRgP6AhjsqWmY
eY8UfIM2V13SrlKnRlawnvkanA8aEtO12UCSu+YcWH3L4T1qayzk8uqAA8Yg
Gdzmkqhes4g35UBAnc0PMEi/7iqZOaRPFM2t8XAn+yaDp5xt01/TuJ1lRpIP
dH/ggf4g8ZSDvh3g0XoWZyGTrPLQ62NSMokF9+nlwPS+0m5JnjSxasJeU2DY
OixBb/EWgKgJCeRLzj0O5+W8NcigeBUAwf2BtMpTBaXHrW8sG7EAJjfhZEKs
kqlCupkp+ItrJro9kOEBoHKMQ9STA93yIwkfJ/fRJAITkBAXNz7K0DPjl3mH
xS64c18eMS5o3PWBx68o1APbQ6gerArl8s08glEpPgQNKz0YM04sEVMjjf19
rL0FC49Nj2QIqd4ILaD6jPbvc9Ikyddt2O3ZRczKxrYZgivqJuXkRV4YnHl3
iO4v1+AHpxGWC5oIoy/jtK27xwonSyRyn0ZwUNTp72rd2/2mJPra2cRB0d4A
ZE/mHhd05aMVQad8VSdmA50lpfrUCxQpXrgvh8Y/rPsY3NO6IKpeKY+wGPo8
HzRo82/LxkndZmGbg0mnA3Tux2d5lQJgNNn7Y5MHCaenLaV+6Cr+1yTr04PS
lRn4Hnh5qsRyScDw8t4kmN8WUhWvMSLScfD47pMXr3EV8CG4XahsGFclwEow
G083cD6SVQf8MrppKhtcYTJnOsR7JmKROonoHzHZ8Q0K0XmKdYOz5uaz9Xcv
a5KTC8X80OvpF0myhp91eobG2B2QHy19VIBj6UBijjPW22AN3hfk2lSrScw9
HpklJIg4k4Gl0b/iIN17C++SSyoMwgj4Je2B19A5XbyAphGO5DgryiC84SD8
f0OK0eIkD2t/GUcao9g6fuyJ8IwTwugLekcClSQXKOB+fUy23eDXSxwvm1tq
zAjY1Zy7t7ZD/1e0p+ziz2tUkNvy5qNN58M3GgwQ8kMWTeQf0LIDPQSfCgxQ
IyQjrMj1fsQfeg1+Q8YZda47Fs4sOS0SrsRgOuY6/XEz//fLmsF61WvpfAPV
/L5YG70wSP+xfu3vWMPQ4UgkA5x2oi3DDicrm7IK93SnhB2gx093zqrObYVI
j8nh1IhY5E95H1M2p5oylRZpB23FCc9VXJVM9VXcytM7SQhs44LPt19kC+qj
0/NF1tB/Ei+3DEs0OL42i/88VZ5Cn1ENz49EPK6cm3DLdoOf82EZcjQuqes0
/QO9P/W8IQKZxQX8g0lcE4xorg2v/oQ8vP603Vdul8poMhS0h9tmE0J3UIfn
tQHWcJO/nAoPBrBkOqP/V7qWxsyHHvQs5KQCKKdgM1KJyzx0/tA8oMMCoo6J
8u1bSJSzv7v2gCfh8jjSepOE/1U9sNofaWkiDij3EmwHviUr2syB1fvIZZqb
FjXdhuE6OxLspZSyrdlnA+9s/iRLGwHftEBxHVVcXVzDci6pqG2fMcpLhE4h
HI0J+D57hYXZPGus5x4dea/ISsk7jxRjqWWM62NaDZCi0cNFiWVaW3Qu28qW
2Ojww1yBiPCen+hFIU0+jWb223CaFAPHVnuJL9tz9i0odlzgAOmy6rQlI10K
ABOAPjcRk3bwT1GU68ngdWS3ETryads8PovJVofWhKV+/s2b7iHkxD4YEPck
bADV0SEaUaYX5DASBIwKggwZRwN08X2XstwhkfRi5wS9OT/M63P6c/gfpUyt
lk9nOCfYxdI3LtJBKvEnDafy2APzHqPH63ENWoonndQil/dkuyGTmNbfD4vp
CnIyIDwJY1u2LZYwXw50+G7IkcwXi7OxZIejHCmB4s24bIMWFpqoEgsPDvuj
H+odFkhyWu1YvDrLktdiMXdCPTf+YCvniRVvACMr08C1a/89+JQy8Wx6NpHh
UFu5V+dcKdZzjCl2ET9uqB5i4GBk0WmTVdhLzGHIo8rcSPMOvykkUO0kF7nJ
Khwu7rDfJYcPe1xoLIYmQuQ0Z0+GG4h92RtLZGL7CWlYD1mjLfHFO2U1hsYh
4qLYFAjiV6Bj2kqmEsTfHHJ3Oofq0s/Slrrk76tFLnvqvGl/Qc5FhwD+o7K0
JLQ3mTPorcnsXascXqiUmHtCMteDdjm8Xa5CYpLub2gngP+lHx9jqarLIHge
u03zbtOkOF9nbgfEwJWu0rfNsdpSIog7DqI1HwWoQqAaOZLddqS9xNpXKgA7
+OmX0mRXLdR7zvyexpnJefkhs82TZw7xy4XyhTesWMwMmzOFYmcPY2Yaye25
2+npZOhjWRE6lN8hr+nxZpTxM8oBdCgNpZK9APFverOIeNQ5/M0kXWHZgGv2
I68to+n/wCvJIa5rYTc20Dxpy3LczBAduHKOOlbS2TwFl+4cqTWKIqLJ3I3V
7kE8HsYwigmoFHGVfs+USyRdsMy9rVF//94JihWh3PFUiZAYuzOnkUHse4AP
Th2PtofNOOa47Psk1Flpgaxu2ZPOWjgm98vMC9Zm+BuZwqcSwxCG3V44gPcv
7+10rEjd33Q12CpN1SASENzeKN9wIHCk6gsD2iaNSQlyk639pgBPjzy0PtYi
+IcFSUVqShwYcu36nsy2EykWtiVAN87dJYgmzcD2UHtPjZi38yelXPP6CSMP
XKebZCm9l0dyrNjwUn0XGFVGQyumWXbG//EgZsJOvQs5/WrKux1+9YV7lrQN
gv4CB1qIQy2XIn+2nBC9PYDT1xSvlI0rz0y4fHAAVcdYLuhnqUZ5URIcOMEd
UpGSnzwiYykouRlzUPmmbTN6s4AEw9u+q6p4OSEYoT7BtDW8wcvA2MgZELfL
vyKeEBdKhh9jJA830WaO/QGYvisnuzvl+zTnibOikoYYVpKa1Iorr6f6FDPE
Hvz+LaOlkA5JoBcR5HaDQZ7NJvwmrFHEGzSJGUSsjB3iiW9EnvOEcZCTSgUz
Yn0KcuDrMj7Nf4zkUu1z7po9SSemKRb3y9jHeb0AJmAA2z0bWrTM98UoeP8b
XpX3ITdKLWG5LcbqYfy+aaoHmkTOqifCXI2/UYOxyomqqzyWl1TVA0F2BSL5
0oC0zZHR/dYD9m9VGL0GJJMjM6pBdgAbNlrhhHYbpdRpw0aUsjqMRuaUr0Rb
2MZLd4f4Lw7b3cK7H0fl/Lbc+KYuAx1DnEq8Nhzlmqft5eJEOZt3V8aL+HMH
er00H2UQ7V+9nT+I25bv1wc11Kahnx1wOUtUw5BvMUU+OjvILblEwoQkfTnf
HL02KYcM2Irp620gAgA1PIOESUW7nThi5rHLeXZ2himLRinw4A+1V2vzFXeC
TZ8QOBxo6s/pE4ZoiP77XhT21XzNH+S+mlx7PCsfmY3C4w66c8/BMpOp9ndf
WAvx38PbiCy+G8eI7M7nApskZExH3n5Z7CSzIpvloBCLkmqUtdJ/fQr/XBTt
Uje3lKPDlLpUqI8+16dm+hO5BTigWuFpPuCgkKg+gs0/nzGKxFsfTCOZYQ52
8/7jLU1i1YO0zxokvMMtwEjsfmQk8ejOpqMzhsTObRU+5JkauDIWRG80yIxi
HDvwUwhn63kGOgGogrgTzeFCio0bZOGCovPQoAvjGqfDwZqRE8sNT6gEc4os
QrChoY2VgV+ax7r1+Lb8opekq3CJelgK5Vw2XhCoPWPLJoCB0LVH5rmt6kfv
cZdYXKZRfyIKA6oAY1yDC+SLG7XB97u6wSMn/PSMaY1PguMU5s6cXUhXUAMw
QwwAYku0k/p3wBi910PFfQVHidvJYK1kB4W5aOzIFMKymTBeZIUnIOqgjBT3
9jgGTEhRLLD+QvBxGBedSznw55/lGLRZ8aShvfmwU9WY9NKKXQc+02Du4dRY
wPJnjbEaFhHuRU3qZtL4CUaWPqYPmoL4eI5OjAqY8xp+mJnZavNCJSs223L6
Q6VIFbDXbIwtcjC5l7EuZXB5fBXF6ECxPC2I8QKJNZSHIa8THljndpS2MxhR
998RUnViiGFTWSt1sx1NkVoVE5dziP+1yXJNNy6PySN6a/+tAVZwSagWHoKQ
K7QI8pwf9r+Afud8sgQWa4I2ABMT5mzJSEBTfvPrclvqCvrsPfQwmMlhpa4b
giFQ8XE7w+0E649I1hlKYEVeedyCO7CuIPcWZqyUxM5bHAdbcrze5K8ys9c8
LHP3BAeDqGbnY+NRvMr5YZIxeHd0jECMG6pWS1/+6BobFGKmbGDRyRWIc+o3
3ho0FRF0DFTTUsCHYqUue1tc6e6TiAvkvhy2tyny8i78qdB96TeFzQIYz70n
F9oAbqD1Yb+a2+zf6vw6o9yPxljoXIWgD0DcP1X5lP8EyLCfciYmrnKpQ7LO
m33IF9j8/I+oFbLbmHtrJqjgDjaPtrQgpJoT7L4ZpKQZ0IIT5P3qe/meT/F0
eC1+bVy2Q4ul0f/k7Lew+XdvcHN9nN+hviOykj5ZgUMtA2XRSH2+HtBgWQpy
x4xdaCKt8OJGPjUqutfXYvoVyiKmR+/V3k4lNgnJP7SSAvuo5QNgEv3YVHwu
FH7U+KRlOchymvignaTPsu2/zSYVhA2W+3lE42DfoQvlaSxdMrhpduWaYuZh
5LgRmf0LYXNndWfMT/0grKtjJpvPjwx4YwVE82JtwPIxDs0TC0kGrWlLmfAk
bbu1/rhndFAsB8EZB77phfJTc9nZ7sR87m1PhXB4S7UF9MN9267od6UHp9lf
do7IfZV9sqABkU68O/+4TWxdJyuoXnGWHRR4apU2o3BfxXEkvhGd0E4O8j3B
VocTwyoBw7wBUThc0Sxi3WgCTMp6T/fqP23D4Hg1Ew8yjMCpZo622IQDSkzv
SAbw/c7GnOHm2VbRNdvPlQ7tlk332L1Q4AoKmcqLNma5V1IHLrRK57xQHfKf
nUSx8gSdnU1r7zWuw18nUdRSWtvwZJeqCIcqamjwNFu47UMUj2At1Vx0ij44
hjHu+MS2gBVEHDcPHrRw5Sksssz8Mj69wht5P143OcFvUUTPljWQEZaWetsz
pRqi+039u9P6tOpBi9HDJJPgNWeIrkbALQR5f5AHvelRbZHVp9DSfBxxkB+k
fwS4cs65pcqp5gRX8KyPaHk2vcgYHO1c4ImpW4nwMnQ6UlDXcZC1ifaW5ejg
gsA+JxKGbWrgSIy1Fh/d4niW900xpjp4r+wvT1Hvm/u4Omwl7akOMCqEurZH
er2xi7rfRlQjonPRP+Si/SNt3yybcpgRoSBorYYkuibWEFd2PS5zQUUHWGPX
vC1CAVI/a2HbAqAP5Xnlb0wEvWwioTZpDrl9WrW/Cj30AvgXmcLoK8r0kMns
R//s2gI3LVaXjtTWjCvDczu8YMoy9uUbTi38V5zCrln2JBuyqB+ciNbkT/am
DTZEJNZbohvzd6t3yTY+EDVTizdIt9/yQ7bn6040E0uIx9cT3Ry++dTYjY4t
mmPmB9NictB9PsA+8ASy58AoFm/YfIT5OshnAP9cfsfd7MxijV/5XHsCn1Wc
M+OP9+LL6QRXO9Ozu58NCqIhBeRxqzfe3+CAReDejJjaahFyDctS17Et6IVj
75QKXO7H3rVSCZRO0HmcjVgwszKmZy0MdOf78p7DA+oVt7IanlfWeYi9NdxB
CezZXPRSfFAd9Z0wKmrhVotz7J8vrn6nj0VN/adxl17s4UcHjr2IGPgitshL
YS136OHLzlw3aJ9p8vCmq7B3wQoy8+nZB/dFByorIHSaa0kQbvJx901D5Kwl
s4JPuaeDv4lIH/oltBd5Vpb0T2a87GJaNX1G5BKw1WLjRfyBtZXQHWBJwr3Q
39I4pugpPX+mZVCNKs06gDbRqmC9mJAAO1OV419ppVDRLRjQPA6E02tDyce4
vXWsVGTCVzF/MFAG6pXEvalGTdnQWlh1MUBm0Zxc6Ix2l5aQlPqII07gzu6S
wlkmJC4dh5qm9noLO+el3tyVHaaS6EFiAzlk+2EtxfCQ/XbZQO07NUqmQnrw
wwljhfF0FHwClZxuDSjfI4a7byIXxfyC5eS4kC1Z5xNRNXsdpmpQoSZuuiDn
UzIbcY/Q6m0NPHjLD4LzuJMPQfoTQu95LF9DSFU6B5HSDahSb+7yQEhehyvh
D9p7deI3ssnaXBRxZewsfsV7hJrkoqO4zDQb8dxFxw0HxdrymMwVYBQpYntR
ryK6KONdnVTBOLfHAip5KcNJtK1a0qzgeofsfTAs7p84Vh7LrHkVhhE8cEh9
0vIPg9VQqcGI7UuDG+dEEoaD4LENr47pEM+OFio6hyNr3tv+RS4DF/69DFBB
3WrUfB+wEcSvHYwCL/V6JaoZ0GZEL2ByortoJjRDMsME1K3kCSDGxTP0C7+s
lLCKM8+NUTGixff9U7hO02ZyL+LwsT5YjRZUQCrWsV5/hrjbJYAngTiDpWWw
N3f/pLOZOFJwYEFY9PeCG7RdjsNJoRPdLoEh6u+vyuzd0Ym33SCGrk2EWNlD
6shrnLco6b+QOuYlnrLJQtkI2APUngPvO+6uFu8JN6S4TfNEtWFtdXVBEcAK
g/jeOHo2YAwyjCb1SieURAY/VqywJ+wzv7G/u59U3BbeL1F88c9e+RUJBBSj
D074YVr5QToAglxwQmAxMaw8qPg16TuQEQsBvyvUcVTOBHvUikC8eqjKfpEX
/SqtXi1EgRoxq0+k3WUk8oHcgedED8SubbVM/yxgVGp0LTE0FEV2uAgYwry5
6IqaRl2dsgHCdfMBJzudube1RMsEvr7c09WQRebj4wLyAOT38fxptpQxaohJ
sB9vyv7tavp+zXUffOA1X53/8EOt0VBfZHu4DkXcH1gbylkerECii1JWNCn+
QGEzSvguEL3X1VwLK37J9pQEp6znq6ybgyg4Cc4btesWglUCkhNeH1nRUquw
tyqEj+4HTkYuB7OJID0I0LWy8P0ViY+N3FOj/BeEkWP5/g076EAYPUcPNJ0Z
5TTfNJnJKub5EsYnUHt3HsIQbqORkpeHQDTtPvCGEZmgLOlxXm2OLd7DHW73
lMEUf489YWj4Eb8z93QJJf+MVXMMaL8bhqXDd1A8+g6sGUvybdHFkZl4wyC3
fTQBWNQo/Syg/nroONrh0544z+XxQ7xKzKAFs5eAKYXvIhPc7QcPIIZMejIh
zZg2hzNGY+ZTOUqz1S/2aI7pV3osafOtuEAOvBY3Gp2VAkuFf38PF74fGpu6
jG5/aiMK+g3+tOHIEc1OVIyWSZ5tQfNGfCA/9B4DxQVDmqPgeSOF4/i7AmAD
MqkQEPHLSPVWYuJs9ejpB+tr84Nlspe89xkc12KKtgIXtXmRF7JDOngLlih1
b1GSLk+Kzbx+dZqtcDHQ+lbQB//AZWS16HrG8spMpPR0n4aXbeh4QxSGlapr
I9/CT7P6qYFYDSWXLXuXl6oauNuLMZG6DYpsUACF/zaR7vnfUiLEIW6i3elw
JH66DfL1DS4uZmxJdWQlUpjFT71ZezLCn3RmctyCpOP0G08Nau0FBk2YlF4D
Fvd3U/A3DciiU0zdMAXPIOYH/uJxzQBaE9qW3nc3EevH/ma7wEd2ssgHCY2U
Wa00sZLivYAfuzIIYxHgX7s7nuaDn0wAjfMFWpesy0WgcvT0KCRo+flGAnQc
MkdCGq3WpVLmD+h97iE3m1qLpxyffGXi9FgxTrj2tKsO4bTixjz/OzF4fn9H
3M/+H21GkdGc0b6P+tsJDby9u3LEEq80Kn5RGZ9lSpYr0E2FBkiwefD7wo3u
LhidvVFsiINou6q56QQfzOJ9ya8Zug+vZPe9+z7eiDlo/5B9zOQUckGpsfhb
x2DHJfeaLpO6RJcGNcvRuL1QKUUq/yyrIzrgl2czDjHjEKF3iU6KU/257CxE
ICWab05OXIsBinKvNZz9FNDGjNySDol+lZ70JpAAIxpdOMouEu9itHrQ3hRc
QHQhLIfDfTAKgcLGhgIh3YvW1a/xaY9rtnXIQdlkbUWcKoB6O9ucPr5BuvVX
2zLkBBYUSAXOn3G/oxjWfsHefehQuGEjO3C82lwCtRlc7A/Y+PnxmP4Q8Nzp
byufiR9G/mtC/2Xc3mlTheo+fr3Ju9TU9HMMZSRtmAJ1nX4knyml8sOMQ2Yk
UPEulA9YVSQSGx3sNFZ9gY1EgOnyzZqSdsfobiB2fIO/oVgxTubRLlOTv8Lf
cdpEwNJ1YMyPi0heLs2e2YrdnFRd4gZfHdfehluJUkHTNsf8/CVbSJzyFaks
OYjFZLdJr57zWeggSWSTIRwbASkBERK0FDq+BKjh+6TYTYYVfdqQfXB/XV1y
YIyOxQ368dc6bdkhLvOkwRNuEX4ATQ8ss+jhJAvh8DaKY6R9fp8ik7zZfF+4
woR9IK3Zs9D8laXISdVNXu0HVK2+HEtINdYiug8Nfqu0i/87OGgycWNeWE2R
hM89huQzAqId5jnMfUIL/QHRRpRQsOxYENwJuPbfKo/3OwUdQVEPSA0xijoo
KTtnkSn7J2dDVLQRuXMcE61TFvC1looF4GkRinZ9Q5yYXJfGasG2f3TkyqyM
gwPrwm2fuuzn8MjsWHXQZTazcAi02TjGd7gdG3x688M3qk5lRbyRZHTQEoCG
7NPW2wM5YbUZVYqxqlI7+skax8WvWQeHXuXXI1giRUGa1uo3dzFVajC3P6Be
WPphm6m96AYANPLlRt1jbIyJj8IEwPZXdRgPTvxWBSS1Iy/ZuxP1JyAgi3T8
f0OvdExWRBl1MJvf6qHW1zH72UwpVSYzHBlgQHJ+654MinVK/eDf2QYosUzo
SffgEttbpp5V7huLhYuigr3Gx7cONvVqI/rHkDRWmKDWTav1zqOLqCVUuR1M
3Oy1NucTe09beNUdHy852TSR2jt7Vna01ACzfp4T907VtMbFkjlft1ixZT+q
hsSNE64hq0RmnQAYspBV1YlOtwUJI8Npatia2Rk24KDwh+FTRrAoIt2yTUmE
CGC2Q6b7MjKWVaNoE7urjFABKs8gljuSaXUUoHUkRF2e10zV13gUI5yl3iE4
zc2/4wZ4zQ4DcelyZYps+C8WIpwA5HbdOYCkK73JUhs60FuwjWELGAurRvfV
e0zLIhrLz7bCUQ7xt3te/SnroIyMYA6JPAP7wzGDvMreBkysPFJzLV1gmzBg
KgKwS8wIjuB1OfHjVqwWhtenzYNfJZWAOJ5VsyB38cHUsvV0ecH/IKn9StwB
t/Wz065kmt5cN0L2baNeLetz7vRR/+hbGh/YdFkg3f9bVmBUKzfbMCr8H9L6
c0cGDCFArZSNfxOeBDvRifQe5sjSQL3jU54RWNSekp7yck85HHNbekUmD8J/
Pbx8G6eUsAIehBxhNBlitNM9gzrz/sWLduD7VcoSPDf5uznIGetjbeV4W+hN
W+JyRsqT4okTe6VCDnbrDZgR6S2yEKbg3g9l1srdiEcmcX1xo+3TajO17n/T
8hf1hXyvUio9j9m6/HfnW7NUgFR/Peyfn90VYKUIE1vFkGt/h7RmOF7Ctpn7
g0LnrDpw/DycYapMxM/Mz59AcJH0gP+d1OvSH140NoKwGE/9VeNT8ragb0ru
5dGzDSsvq6p6GHjyIh6n34P144s5/IHg9uWc8LD0J+wf9ezKkgLIqcmle2Ia
FA4REstBbrSD5EvRpbij2WYEXHfdy124JrKKa7IWjrkAzZbr6fspiVI/sMJz
chxlS2pUik+/jZTFLuwMAuNIceM/vx6zDem/h6FCLSEZAq5V4OnsGGqMu9C6
L9kK2ujDPm8DJkJwYiGzv+1vnPco6h2ckNCZsNZOQOFjrq2NgN3xd5ngqdGP
NfxUkOQmgraGO316a6BXhBZVhTH4DZcE8NmnEecywbM0GV8Be7xGQreRDJYi
Z9jiPWnbrdpm7aHTCWqfx0dpyDE+327jeNFulSgqzdmKpvBDwrNoAYEScfsY
MmpYAY60Y3tzcPAgFuYbZ4jqQin6gG78erVkf7a8L6KgKcbbDvZOagtYpPJa
fWwUxKFHVsX4mwhCztLVMIYaSEhOgBvZsMtMRFSxOZFfrzZYCB9GlxMt5osh
k1tEyTIdY/Na8KQM18Ohuz49zbd6MED+0IhStg+JNs8VN3/iLbjtUQfEEjip
fd1RT9D1h+ni2wOUqqJUzJVpXIw3t02N+RStBCozwRiG3NrsX3hkUdEhSAhV
UXnQxkn7Xxp5F2nHrHtyRuFTzWHrkuxsDeojs2ndJNt6hbY/Kj9xiUx8TfH8
TfF1j0V/6/fIaqgcnZSK4Ie4TrPbVovf2ailE16X2MIwFqvxcKrLzpjDQ5Gf
88t7JvnqSyu+4nbGDu0VO6B71mo1K3GZnbiahlLVWRf+W9Whsa6fL8e0PNCW
AcFaWVde8pb2umnsfGgHUBLkCTnXbFN2+mOip3DTOGwXxb3iCP3ox3ujPlKc
MrtZdcijzXRooQEf+vrnSxEsVOfFBaSyFfxk4cJA9RBqth9omQlXSxS26mnf
GjE8gWQzlRSmaAjEKYUZg1w86DQ2iUyn9cEjxFinOS4qrqKO1LXorr+h0LY0
5g/DM5RlkaR/c7unUPpdCmV7pWMqoBZoWBZwo8eticJNk7QEHmqNy/CQOxjd
+DHzZcwivnTskgXsiQVB6bBSNs5Ou6Njo8dsz3727jz7uyz11669sTiYhpr6
KEGpSdFt0OSyktr07uFUJlIhIh6hcbh99Le9/5qENbBb4bjbF/HbXJbfCNEh
CM1O+y1Ag8k02eHcsIKeU/LeyO9g+aEXH/l/GAI5pfcYZ3xJOh+g9RUe/bz4
0CJebeHql5tj8Tt2TN5Jb5VbFnKYCKC/e7FIZ0q5mL9nGNty6KPt94+sAsGc
K7F+M338QcCJKD1htNmNlDSR6ncYxbC2q3AjIsZVE6NuMLn73K1UDdDKToG1
WkvxK7IZ2777U7nQzxm72z/2eOF7f8Np3AYiRf7iCEHVtX83N6SqYcffVwOZ
dUCVyyxQlsjzbdCvmQWPCMyEiabwu5E3IbsiZRm20ubSHk8efeFi/fw9LHKP
jViRpHGoNGakUGThkIOcxKyKhMO4WsyNcxRdsZO85SI4FZUyXQbcTrEOzufg
hsdoqB1fA6NotSFGc29ajqN/3I1YLIVFm+Xww0zjgFXKdFLNliBFhX/EBTEx
uX0Vg+fbFmW3fdvRg9ErC416hgoz9jD+Ps+usDxLRjj2bKa9SK98gE5jkpYg
HEM+JCIzeU5onNdNLlA/g/cthQfs5I1OvnTNbVhQnPYHKQKd84wH6ASuXL3N
+u4u2q7K9hkyPQFkbe1pJpEuVCDHw5j8aeAaMupBNRBe4LHvVvSRlDL0/Qtb
x7n8QjCvLXgVdbTucVjQXP1e/4Gh/zzsq/rbdu3ouczG7SaiOuf849GN1yKw
iC+XdaBNY9P9WjWq3gc6Ns8UMFlwJwlBIQJEhKehJLH7pY/3/38scH2x3gC9
7Y3ooHn2pkBRtZSY0GBgrnQKKLeZlqOhoFjXuc8gDxNpM6eUJNPGHOuXuLkg
dEvaoc1oyv5kB6/eg/TqpUUhWWvxo3kVEPoyAsSU8/rApBUrvxrqzLPcHZUZ
5I8rPv1zjkti0pjkxDHgEGOMhvAgx5vqeolv2TTEyGvVsll9n3EVHJeCUs5/
VuMiHLFifIwWc2o/sSZRZ9TbLTxFWFSTr1zKDfLof7GdIZi2wZnAXk4Hy8Mg
ikpHjWlbohhkUeIixbZJ4mnF3uGf8blteix42/Bt8maWp6c7Jew+guuXwCm7
lPsDgbuz34y7qg2s4Ch9MQBPxIl0kvU8l8k240Kd0HfL+GsD/+9LOq1fiUpq
cf044jUcW9LaJ+a7pLJeOiTpxxlIJXmhaO601R9clKh7hK4TgvRJdBvcwqyy
Q2j/2PWHX70uVOy9HDvY0n4Jqr86Ng5OlNS3Qkk8Kr6zoRdkjVbexTdvpN5N
wobBPKbR7/KNwdcypYnSxMYzoaCj08/Q4ioGpB5hgjqkSm486DXK4X2DNzTh
dwav7bMAuZ2wMC5uvG6ArHiwf+OqU0AicA1Oc1qv8j4dcZepQ2Xg65K86Otc
8sKyvBRh/0WepseF6jo3Zf4HqtnnA4w2OY+JOt+LK2qtkUktbIQdKMEKo2Oz
mkXkuAhxIbBtPc3WzGvVOK7/wIUCJ4qPgMagw6vemXDcNJgAKhTAU8JFk+a2
LoKiqBXKA3WBK6EDKWg3yEtqZ3Lh3F7X/OSnTGzOvGzi+3229mcki52x9dLd
4YJlEUaz8lujOdMToTZfG1rheyb4lke0B+hP46fWBVQ4WiBewKSeT38cDtk+
851Xj89QcbgOP3cT9/xIzm+OYQ88QWussRC4XUW7Nh2jnHt8TjkqH8K0Ts0V
LdVHSgdLjIhsrXkWJ79aYxtcCgSx/cIk9wja5tn9E0DN0a083rfLjkE7+rye
RbN7RnodPcopCbCvzR5EtI44IH4jFDNCvFJzpVOw7Bzdcz9Yso3wmRPj435M
yzFhqZ0wViq9KWSfj0kPv3I0hOgveMzu9mhC7ltd5b1CebsNK0HEncomafkE
2QeHQQfj+ysu1fyoFr/x3dqcsH9WFJT+CVUYUj/va/uvk8ImiK4an57Nhf/W
wV3fBGOpgWfRw9i7caU7cZFo16RhvYTF082dPszTSp+0aikphVKobTGSlEac
RLUjnN7s3vrBTWi6caPuS1SpzoSCkdQK0TCYll+woHqRn74SlK2pOLUeDZBY
4EXr0w+HjA37prhHVXD3pEeMuUevycSB/m/DvJ5523xG5IxuxCPAzs9mG2tK
mRCzJ/Z50ihwg7UG99zTPDJKvoBjPOMJiL5qers32i2XrNjYlV3r8FAnxFaM
bXboKoZLTqh6WT17bpFdUdJ99B6yXjfmYGxclndiDkrwBBUCqpbWjRmSoEad
kHYNghwz9zl1geR+SDjy+DSW+vHbrMxUTjgiQdidnk+2Z0EdI45ayHcZD8SE
DSSEjXb0S6exM020LzuuOw3dqELRKuKDasgH4MViVFM616u1G9OObcgpXMLN
/SGzKXRQcfJD0pOxj8vbqk5pvwY+JomzU8aJEQInf9TrwZcHbKSRlqfvc8UV
4aoBtM+qtKyh8vC2luI/35/6NWvMC2kOyhEFbDA8Sp0P7s6P/XX6riIMD1ZC
5s+XW0vk31Ubtjcx5PtNu59W6unKw83QQjvE3kp+NJLd6uXAmRMuk29cSD1B
md2S8gyM4f9amcpkGM+Yf9WZkXnqKKJScqtSYI45Dc9IoAroGFkZmKBPLTVv
XnaDHkVDlbZpi3q/+imNzVsTeQW/7rlFJXxXZgFQ+OOzXtrtzsMI/pmckoRQ
NVkTvycyAKbmGp9LA3OQSsC49skT0x/eILsk9yFFEUD/D7p+YbOyekHNTY7q
RMEvfzgS5wcuO3qK5ucivtiFRGYvq+QTibKourpLa2VTSYZZVLCuTPPNE2/a
WeSR/hZOIt0ucC7XbsEUhNVBL3Ffz9uCOMDKEmTPQsgG1+mPEnNhJihDhPh6
6A8f5NNddPEqJWG6j+hZSemHryASIKIvHD7E8YyasXIyWShS/01lt6vUP1CG
Kt4hlGXll+CXOBpI7r/PPPgG3lDPw1KjgDXShPr7o+XOgs8SymeOOc/joaeC
3h91KWRPkYJpJboqJ6XrPNYGOM9birTx6ariDJPsNxa2f4H6fl7WGRI6PCpj
taoYP5i6n8Xb+h7NBZDZNJjoTuaSa+RVHl6dc2V7qpwf+77celdxzSHCznJD
cC7Y/55dVgCMm75ZdJckfN3JjFeLciwFRX/12hQb438L5Hk5p4PWHOGfRQan
/FpNgcotR4gktSqTMUmQs+7cWLhCSBlnXNUMB3wDS6lck83Ufejt3pHJ1xxs
JTU/8yYEEfDUcXq889T4rODwRtY5mD40fzluAkpRF4n1C7xMy0AMXiynfSfS
L8hUs9le1P5+5x/R7NmLPNOsKr4BCpvlx8pBU3tKa63Bu9SbJhLVDrBNs+ZZ
Ns99jI+daPxEl+4OubpR9bzMkXXqANlfOivkOMBWqHpnDn151M5TpFrOKmw2
4G7Txa0UhEGB/z1BiTvB5EZeAZv+KvMY3nb/f6zWURMrQJDgeRU4tkWc4t4k
atvVaNxFtbwdu+6FK1GTYo8x0xr/nNY5Wptg6gc4piKEC72Ku5MFGg7va3Xt
wZCYqKIi2sLsKVdkn9qM+fAGm9R25Z4WGZkn4wObikerYvThdm12qKUG8UVY
/UMJIucdvuPQARqyXKq2xBovgdyQ9FfKgTEUAUiieVZ5/y5AQYXSypDlWojS
XUk8Em1xwqDJn/IbeUGq6d3jwPNWRvQJxJQg3T9uiMJZqkDDVeO+4aH3J7Pm
0genOFhagM2vCjwefvgnyeKbYriEC3GcUxwfxDNeTjY/qNWywuisMQ+vJ6QW
vf9hYbfBLi8ITc7fAfZ1ctggbLD49EzUCUUIL7PgeQ7ooDg4f17SNhRwVTNJ
8wOHF3d7COVknS17fgqRMtEYaWBtJaeUwrYTYtcY8Wj7JP76py9zjxI3QLtY
VRP9XnOl6ThRtici5d+qOyNIIoJUMMrPkXBI2ykoWktMuWc4KUBUT/ssqg7c
d0Dd/m/n7auuAa7nC9uFo3BgVYFMo6skXviUflULkXHBBjFzLoJ1eFaEm+K1
pmvHJmKXC2Gy3QOeTwwpjDLU+6tfrRyZXmt/kbVpLvA0EmiYjhZrVDPYEBFD
N6NRdjZcT/6tNvOWnzlBFEoVcFVZgSX1CxYRLsPm8UX6isXCdbl/+k9odA0f
Br6iTXdVFjtPY2D07n4SIGeMfvG5DGQ0J4LttM/uhyDsUgV9nQUM7Xbdf0/f
1RYSu6kWjx2VBQnnC3ZpFEyibHjXP9vgR+z2JNfoawHS+yVz/CaKnUehI/t8
kZMHaMN04qCLYSFU3UOEYLZv/u/uKGyUeTAfqPyK/Uj1+ni1AkFuJCoroIYN
O2meNQV2loufwlG2vAJo8dHuKWeSWtzQhGirJtU5fyeulbynKHLIms7wMfRp
YNvJOpQK3Y1h83o2o2+4fGzKcv5K8Ym9AoGGyPFuw6DnDWyEbQRDs6XVmPQr
neIXb3igaiRO7XubjE6lrVx+fK0qCPvEouezS1i1PlLozsVg7J6EEriNl3Fn
+uFq3QRQy8dIfaCBf3P3Deh5dNK+9X2yW+Eq7z7Q5VVnqfIrGnIqSowRubpQ
w3JpMhUTGdxunzQiz4d6bqrqVOg+65b9w9cQ40KS1bMA+ZUks7B5svJwC3/P
gk6sDCFPwmeFcVQMllkZ+nqJso5LunLptwDI0F9GrORgzYrdH/D1DkMH21Ld
B4h4tsjBNFVoPN1gjvJveSXJCRG/YZH1r9Cpj9nSpCtRVaYsD4i8wm+5xYqS
Ptfoax8HK4PJUcx/gijfr26oIHU7VXk3d8zerYV4QNkOcmPCOfPu9IsJ+Vpg
S7TPMu+LTx52bPTUYLdlCIb73Cy2WTqGoTGf3m9xZotjHVyNDp+Q+Dh81UM9
ZzcMepK0bfQNM7fhf1+ro7oEPch0FwZbYdJPfZgVqFEMtSOsN+UbE4m03JKB
2BFD6yw8fiNF6dRCaYlZIYmBYiNZPmm5x1GuHg61WcNde4YTc+SnRqpAIsfd
WutnL6gPt3GRaKyD75l6HBUODNcYrkso9mHPo9WIcad6jLGnhUJo97uVjY26
VvRK/OLmFKtGBmfhGGBsft3IGgaEE2FCJcDwzYxmmEqmkwZtDAP81uOtZ1rG
empkGWTCrzkfXxktX8iVvvD4bJLi4rcepWmsA/cc4CCxVC0KEIEn7fVLwq8h
P27V/cA0Mvjni7BhCiRbm/s70cSAM7/mXJgG3h3FfxZXrhMKeaun8GOIsa/Q
ZCQ75ZY0ES8b/dd2EG9yfqGKfNMw9mRGoNX/cZpVSgRezG79DToUEgznDSKh
zJFVq/ZNnW14daLyeeQ9BG2vwM98ubEbkMp3PaCYGtRUr7UFgHAaZfIwCT+l
6mJbBZPnqI8SVL9uYAJC+EX7wZgioKnujQuuyFuOH4OZzKIjQXGkXtvO2wha
gRMPFJs+qUfqzYCekUG4KDd+HuTJeBtxvYJVR/VP4mZ/fZJKhDkuVh1yE0zc
498uGgHpVThgqL5apDeYQiACjqbiP3a/PdlqVVeZgSG7xQGFQS7I2/RBvBhy
GRfjLa5Hjt5Gvrm4oH8ufvpzgaWrg4+5mnzPEYLHubGgfzLjEC/iYR4wz3+J
8dIQRrAE8OeIJd4iE7WJMakXmUXnzAvzasVIU0dZNd2a7wS9yQWr/9xHFJkD
bT0JeJbTAumSTTpPKk9RQrGuHh84L3cpIuE/7K27HT93bGgM12rtjjipXBnR
sD2ZpvVaHgLsh65rOpxrDpU+asFZF+76oP+3UYr0lqbgfN49GG/O7aKS8wmG
28cOH6MgfqEHVbi9uIH7zgqZD2/aaXzVfcmLxRVS3AG3tdUJ9oqN8AKNv4ZB
fjs7B1fXKpZbwkjNbz6Qvm6XoblwGDrvDiaq9MQ2hgwoqXmS6FrHm1ZQA3di
ZA39C2gkC0o3A/srJ+fhlTt015CqlCxW+Ia6oSMo2vlMtjeZ4n3sEdAHgOa+
7B2d84WXWMt4qxi7mLr605TTeUHbgJ45iFFGodvVsZSOHhLetb/Ujm1vufZ2
sCvTrZ4DIUmfmyCFtMR4Jw59ZKErznoXqwfz2B5JWWq+quHS5gFiWHyq36i2
Bw4lTvs+WE7ovHL7GH8i6HHuJkHMqDP/vrbPZiDJ+BVecPtQWRq4zoMTVIsP
LRS+2nbZMvExtb0WicMj+hb5ZxLwrfCb3W6hRllkPI7IwIedAjpHwmWQl0lL
MKxUWeqsBfh3DzjU0fJrUuyBdugRsQeCsP0jRsOhT2xrm7ZCN5AVuR+Y40Vm
T7Fvl/s6JN6JFSjmo3QqrBX44T7suuZSiZJXmPos3zolUUARxW1W43YYf0ej
Qg69EavAna/+CdBvmwePqrI9b+RjbqbeCwDhqgSwZn8MQJ9uIcxHCR+h14fV
1mijjbhjY35G1onVE/NcxdYRNKWG+fpqUdcdRd8ohRjNcSB85J1AXvftI2zQ
/b9uSK7StNg0PpaHMWc4YT1SIIJYfI90AGH/SvM8ZXhrkEExbVDdl98RPMSu
TIvqSNaakmlgItiS0oWYRfKTxO3wJm1BVOD7y5tQFdZ2szkFu6Ayg2PuTUZk
YxBV0cNsyUVdMmDkXfGxmva1NS2pQz8qhsQl5rqJRf34Wf24DQnKC0E/8PW8
pYy9SdzfzJ7gVeKzSDBT5T4rgvTpFs7bpJuFAUxfCZRoc6T03wnB29414NXy
5F74V0fWpANSB/oKyCSkmhobCtb68yW183iXDu1kxrtw2Zj2xIa5DShHnshW
/DNBXABH4fzV6xDuwT6tCLag0hiZwCRJdIR9J+UkWR2JCK3asmsg5uHejIQX
X5pi67Z2zlERLcbq9n/sASk6RIc9VT/xJGciBWBEipltDoOfLTQYJnxh3reZ
uBo70Ylrx1RVdfdXAC80TERslKXmjruvgFVfroXJvgXemk8tsQXSyQNc7GkZ
If0AOHpYS90lNonB7OdNTeo5TvzE/9KUnb0kSgoT+p9rxs3wOP1/fK+t0UQ8
Lb/9zobM+EZm9ZyJMWH8Vn8LkPaAkH3NSJ1E3ZaYk4L/MlNaBeAIFfd0Oa/W
YqAGZ9EYsM2jjN3M2QPN9gDaVh6tMDHWO4tphBIKLWX9oLXDGLSkIltMsOEg
wl1Vw6QqMhm/gjV4kWCZPGjb+fOEVsKqQHO7Pk3w/1FDlbcrTiACGoEPoD34
RsVwEp1lzynm2KIGM1l+Z6Qu/FXASz9qKDylQdhxXT+veMDG00Rt7RORQJL7
Rhm5JHpEvSuFyPR5XZi9vZeKJ+SDnonu4ayS+x8T+IR9Ll6/lubK9otRPTwJ
jViQARfnSE/tcafyHpWR7XxbmJBeBjk4W9pgtk6vmQL20FBbYmh6/6cOCMdj
uGpT4L6POERuViAWUNNOv+7EQu39UnaY4ExLCGbom5vH/f6q+LCCyYiRX/UO
4ZLec2XJlTx5bDFbk496bXLi6Y+4wgCBLT3wc7KtgU4WRUiPwRolJGnaem0L
Y6AxyL0Am+42FscBJPcCJhSkt+Xj6gXQLX/kKD9byOIHGoFkZTt52VHGOa2X
eDejza2HlWkMMgBIJ4PdQa0aMqejlb/h0tmfvUAbrpzbunQOTonllKhVyTh7
ChT+NQ6z6zS2pNA92S9JtqKvNpyimZIJVmcGn1NlHbI9C+ijNntSIzfSd/3L
RtvtUxDRsqF1cKNSEBFcIWDt09xyX9EhxVtHSwcotmZAR3YOiWqc2PTPhgg0
275FakuWQyFNydKSpBN0ZObwEIXkGbQh4xwCsaQIH/pqzqdAEOgfMCjw3+6Y
gwIeJOx5Si5VhABpy5v9vr0Aa8oEjZSPSKeAh5wAIOBEJaG7XLtOdHH+JYsL
zSfR3wTL3oP1et1aFqM+0seEkuwnbqxuJpc796CNaQ3TqrfCrniHeYtUsd0r
eqYXdCVQcjAvcGw/HqYml+/wK9PbHss8XWSYt1+CP8El/l4pNmegctra7rIs
iO+7Ma4ydUJh5YowXU/PMC2ZxeJIFgYRj+BBjNDs2NrHvi5scaY4zbyAX5Ed
VCbH9RrV5S0LJ/e9Y9zBlkFykAajc9hw+I1iQqUUZtUIfQkwFEXrXqW3Eitr
xpvMrdvG89LuYN4pQmM4yUeSbZdAMHkivo3a6fCIhZBTCueaVCw6xaVyxFPJ
AlIoP4FMZZa79oJY0+TXGMtmkfe7iZ0FFABJFirLL/Qew0MvQlgStnpT0atW
WFDt/M7p6ktL80LhVpcUoh///K7v+UCGTfs3+u8dFo2pUoqeRyunAaa4kU0K
h8Ze1cS2EPpq1EWs8N30YK6Pyt5usMhTc/DDz7MRwQfj0OtNuGtk0RsUjxED
HKzB8k0PsqhwC6+BEJmmADNoW6HxU2aNlE9PY3EuSDOMlfZSfdUFUsaiIh6h
2l17cvD4aSfXpYWNP0ksgB25Zqh6dS2qW35ylz+zMIMVau5GloHcJJZ5CYfB
5UPiDSxLKACtbNSzy1kPuI43hbgQQgpoVQPjp4lNNQaQDci4qF/3NnVga4KO
Wn1SGp95+ue3WBgoMpiB33k+WSY83zE7f0Spjf2Sglth/TFjH7m4uGrSscNM
w+8tRwrJ9wmfGAHl+Hee/U4UO7kBMCJnEZ/4QjsypYThG59WzugK6QLnRXlp
EIVYgG9IcradW24w8kgfp8/6X6Lh84Yzhq7sgb3O82JBUOuId2A3zNe3Lryo
rzRIHd4qqaT5/gtz2tGH+4MA0G66SRk/slQd79OIpWn+WtFXju78p9z9iy1U
ByiOrh+m1f6mXXrulrb3c8OXUYT1UyGKgDoTGYP39bmaJ62JPmfhsHnzhDeC
6y5TwBDN/tBUTDbBq0hxzt3JqQarexwH6nQQYWlMF+HAwbtRC5gFyz2GPUv6
j0liKxhjR6s4ULuky1XebvoNaJ+KWRGMhs24p1EJCVSu6+A6d0+gagsyfLyZ
dhGFVD+7SwH1W8l/tpa9X92oIqz0bBrF8TBFhb5WmOpgzrqXMimjeFTPCzek
bgpKFpcI9leSK8zgjJvHBjbWUvVh+L3sGPt5EYjIb7vI9eZEzAdZJeGiRrvs
ysIxa6O3W7h1hnmPU89NRe8JLqV+ZBzrz/WR6alTzdxwQUkYmZxPvJtO+Pz6
54rpVDYhjBDhm5TShrRDs2eoQrddeFV+7l92PpC6GbQz5dHukhz6ZWBF532A
S5DWNV2aWY2R/+2okwvcpVnP6eDHS8Ic3ILFILYLMGgGBrPRhZKTxdjeMRlE
KFL98Q0d9OqvQURPv7u71fEm95G9S+GrSGDe6stpNWQyXGbV6jQ2y9NeZ1qa
NyxDFEvrBVSY+2abOVtbhHbYDcgh4DPbY9bLSZ/CpzHHZHND7kIVuBlEg/ag
W6ABS515Aw7PfnpX5s9PhyNnnOa3LlsmNwagnNcG20LDKEuEjvMthNMcQqTq
udPkc7wctTVyfA5I1913cMBEZuuTUwZ3H3XjCYGi3ZWPaTRGgiJRMuVAQw/m
i8ekNrN5lQ+Q+KF2Um8ClY81k0HYlVpS38QWcKqmCJLalsqQ0YOHOl55SUJB
nbI56Yj/DaPSg8UfLbi+xHDQIr1EI0802/LkuVKoLF5otHLzL9QME/z62sFZ
+T5CjqqbOq/vudYcLJxpaYnH0zzLPdcyEdA6OPeeBo2UDoMbJvE81w1HGxw4
i28j/4TsQnFO8fmH11B1SRDFjUJj51CIPbvIYkIbce+GIpdEug5kB8DzuUyh
13i87ac2ccusAYD7zQ5hXTEKUag9vXhfwR8p2V25vnbYRhT/UTPgnPfpHokj
UaV3kh6C7vVd802kXIyERr9dN5zj4tgHTK5uBcsdkLrkoi3buR1ldpWY7gP2
9759thAKnhW1ZyWPVQQdKR+zAELf3uV86syGQi1VEq2RLY1QZ60paYL5yEvW
KRxoVL4P798jF06dY7aeStmJerd9l7mBfh39BYzsfN/+aNBaPYnSQpl1ip5O
9I1wo87yrIASYoEu2JCji76yngXhc2tRu6WDXZJfR/GMW7k8QhrVR9BeTswr
b7N8EFKvbxQsDFZ6vrAjQAESfOuS+GuIX8ndJuRYuI1N4uopta6Dyqp9CW6U
ihBJAYSZkWU5ON4Rxz8GV0lfmavnF1AF0FxJgeWbF23mxrQJnuHXgBsfz2XN
6qRfkEPuH7TueTxZGHAww4d98YnOKvbd0Ge39ZF80xNmJyAASfKnuQkPOWop
OcQOqy8xjnGMbvMYCdgjkDyo5WiAFzMihLzEi4EOxdfYNz8shSo3yfC817C7
hGTLya/VNHflesJe7ZK/U5jEzrjqDH/M6h75U3pgxHLL9srQbP2Ip+anjKTw
6Qfwuf9fI1UC6+XpBKk8Ds3wy0kBryh6zb+z/nyAtEUFWLvcnq90qbjagDwJ
U4B+dSMTQdPQPq8xvHyYvWwKWx+U8gUHKoJgoW/dPJY0HbZVyYKMfco6huPf
fUNzJLASs0KJbTZwlwV/qEtMAlokaKLqKXSeN/2tPXTfcyp3hWj/71kiP1K4
wIL8AC3U8o10qLNXeGHzIsOfCsiNTPeD4EIY1YzAljlgE02IO+AgzjgINQFC
4aR6lDEqhGOS0qzYcMkQ0z8r3/I0/v0Emb36jq9Fxk0UPo27qkBUGIItNATb
bBHZWuR2jHtWNPBg/SDOwXVVOHputFSyKcMzL0yimjCNoklelVu2bP406xjj
0kM+S6fI0pWLqm5nJGzgRsoze+sbKnl02yyAZVHOmDW+76C8avfuVwJnfnAG
gcuxYFrNEd9a/I1fdC4U3j1DHFB8reyuJEfLorlswWPGQ+zgXWsbZ6kIDemq
21XL3W41GZgX48htW2DvLji2EiIb3k6+IFKqh0yg2vD4W2nQ+4oqpW7v7eX8
ImrdMKUGsIKaF55C4L5tK5IdkNr/K10x3rNjLBcRdUXNaTfv1vjMxtA/5Y4P
+qlvyjv4jYtsUr/X4Kqj/Ry1OjTgskf1hKBam/CjZFRX/TrFZANlPxzkwTy8
/t6T2dVmrmrmANfR7nJaG8dASMhcj7216+iNCZt5siPBOUEU2aI9vmfEoXrF
YvtWt2g0SDUZqKDC8EuZSeFddSpFOhFEQCs/lmWhPkEGqJ9z0u1T8F4/Pq/c
NOZ5ZzdGWT/U7SoFnemsDFdEUYY/RY4/Eorx+jDBTHKM6hpm5lYcN7RcvRYC
PwzTTgKvNyv4hNcoV3Z3H+YuBNytE0s7iZsuJSonTTY2D5G2TAVqN1EqmTKR
lD6VOUF3hkVlDfPN4i4jsmyZbk/EcSXXiUItaxO/z8c4wjTrjoQcWHKjL4r2
Kn0aCV0XumdqoP/gOZ0dhkIUX8P6EWnXkWVijpndjm6yMTN+/7JY3CsUfrp9
ESRF1iiCKlFssQu0Y45aIDHfCnqE8SMra2O/7ZaYrx0927v8aZ5TK9Tux7Lc
Qg5YIGL3FxfJBsQjmKu1s5cy2qJIDyRlE/u0qhtP7BLo1Dpkn2yvITY+lRtd
gJ2zIqWhfXPm6rogFwB9rGPz/l+uxwGzwEHowZ+fuifinqh47fUkgwdQE77V
Dauk5fq6UvOs+TT2knaT2uMzkuQjHVoZkzqZQ1Wj9gK2PpCebkWYovkAYgzZ
/zIwgQgqh1XxSxvCmQuLCPLfaB7sXlVHB73yNiZ9svJfPst/7ri4f6sfdUtp
moB7+Ww8VrW+jUxl9ns3FrGsYifgo2Y5ag+duhnQNE/Y1pSi4AbwihJSCF9D
EDmExbrJykyI75ta7j7OjxSqUV9zw/W6Y3KNXAsyzpBRvsGMC8BOeOlZzy33
8NcoD0V8k7p+zDJ6PgeWF/rqV2Mf07pD7oW4I9p2MvBLVFxu3ucjvWC0Uhp7
LDdTqGgufMemmXYx92AAsVCrRh1zAgFmUOEsd8qc5QsgeEfNhQg6egvTOEEg
5Va7hijnmw3gkgI40YLqNXfbTXGMvHoVFVCif8ccWPZhjhNAl0hIMAP4nGrz
vrJrL9EJvQIwKnNh4UFxzKe9WmRU0SAcORBtv9TZv3vBBKdb/pq6opbnSj5o
JitqT95vFNoH8Bqs34Yn2ScEJSdKnj2wOaERi/Wh1wKXbqIBStlM20V7s4MG
Xw9cBQgx0hpVtY5bLmCJQENIwg7703B5pdhZAK0z8QMYaQyyKAobyDGgTOUa
iRnutE3wAYEb/tvvXYV2yMB+Ln+JUEmobXdPIdB9c4Pb8/mivL/FB/5GQuT4
K9D0GLHCtGqduYJs1PdZ81TKrAa9F9YLsPX5+Rp4iDP/FYcp5P77kod9RVcj
86xLM/kbPkmE4MbAiW5UvLL5Zs/ArnSom+9IVF9yvQlKZooc4hazhBXxx2S6
qZ3OlemlBR4iTNX3EeD360GISx3QI6Fx7O5slYkI2kOj6F1JtJEgvGwjhTIy
2W71UM9kyC8niKmHoprhjz+EYel/36OoT/Rej7htvYx4TFvjsJivE/Ongd9l
bfyhzjchRGfSuBPHuh77grfoD9xbjtyCispdYRdpOG2vlPtYParo7js9EXVX
155bBpfCbQmSTSegd5SmsYaMfTm3szniopbgHRF4IDChOiKMoAzJ9hqCc6V3
+fvE69jde0sieFXWfkupIeHkVghN02B5NSIad4r3B4fyAPFWBUHz4EpFZua8
h9MPq6y9yNoabSp4o8r50LhPqiswiFDmxo/UoNzWZyT/3lJkJD1U8jl/Asox
ecGVu1X5n/EkjEK7iEVlY5ozXGT7MjJzyaptZujb7MCX4afDHCvpmmBboxM1
MjKO9SG3YXNr/DhhLqpwLddp+6NBQq+vZh+IACqBjKZJF9siR2/Zh6UVOFNz
dYlngfChKOQhbGDkhlopkMCnZ6Kvs07TMOCYnqg9c6/0/QFKvC2VLTxJR3aF
FE10bAy9v1DVVgeDcq2CuNkqr71dR32bKk6TIKFV+amy052VbYxyfr+CuQUd
VApxAsf8SILwdp+KQyyM91nd413h9sGj3QwkU0iBGwEjwaCT4Qp0SqDBWKkw
s90Vv7F0X20yhwWM+vX+4b9Q5WLgVOnnJmUXOLDVOJi3Yw1x9U9SFv9JAMMT
avih+gxgYzgpV07WQzAZxeBacEENYdvc9qLDVwEXhAE/aQ1OUBRytCODZngj
Rpz+MHXGTAocS6ucI6EEsWG+kCXxqYfDjM/nFo8b3Ktcc+IYDufseGDq6H2I
lkIDD3x4mc1pchyOe1tONcN7g8/eg7MCZOwe+p11WmAFcf77V6TyZwrOStSB
MHHgSCEFZ9xGg+hfO5XKR8xMk9s/ZnyILlc7JKg5XouuiOqZi9agHVE0SGbz
4BElMW1ikjkdyRBXDp/TzO4w07+o+AQQ2gnvMCr1hiGlVb9gl6RgErKA9nx6
/22ZakU06ZqD0ajnEkgqWL8hUKUOjtDAcXFhO0Bfr1Q/pHPclo2jH3eGxZXY
LqiqnRaSPFO2j9UWBGKMlysdKnArB9jr2vxs6APGr/a6iUTPS6larSXuXuNZ
smHffODTjMKFqfLvLZsbeVIrcXZ8IE3rjw62/fFQZMDt/n5Xg8yLijUnA6JC
13V6LeRFMfYy0K+lHOHHUacBMx2vkhL1Ssh7iI6N7VcdjefQVVYaMbvGnNy5
TI2Hw/BlE9IhGRLAn//UbFNbO/eB8JBJjcNpn/aiqyzTyqiulHGsQQ+xaasJ
IZO3iY6PqILt4BMtv8nUPMe5grls7ScHWrxjgD6miDHcWkMtugsBG6vq5BpW
JNB6UBi8+ezaLv3yXfsLF9+EnA3FsebzTpPxqRoVBJzoaJCRATiRtopArGdo
4zcJqm+PV1SHMa3QSIgXw3coNT3nsaLj8TZ9jXM928pu3RQ9RpNTHbggCh8e
xSRqkVsAgGLLJC55sjwXvny81cnunJjNYfSsxPvgvaojagUbeguMUisTyJIH
fZBnlLO0dmcofu9W/c2hsU6buMqWCe4Q4BFn8JB0QR1jlHIXrqkt2WYRGOJU
7YCTPPni6XO9cJstu62M8CNV36Hfpw2KVZTlIGpBepbhuqKy8yY6ZG43dDFG
ZRvcoTrimUhKMUASDvJyCglaeDPX3XT6pixyaCTmwEKPDh71qgOQ/M56caex
HgsXITmYgqIic5jQCvqIy7uhgEYlJb/f7QLJUJHg2LZBgX5S+M1A6ZxBwPXb
4XctSMgozHYFpU+p4fJ2JCcOdU70vHhpxVBop+Y/ouoHqPT8l4yeGHy0pEN5
JBJcmx+TqW1RlDeoRhWo3b1VIvkm7IwAnIaF1Az8OLdGsTSoiLNcCrDhJ+Kh
Lgm4hxbky7PB+F4WX1jMFHyh1U2nDp8Qov/1Ii8jI3aY3cX/LrFlqPAWo3FA
uUWOcfuJuQ7WTjlZXO3kuhjgS16vBmJ7HyGNCHucn0ZEFUvBapdUXZgIYST2
diL2xf3yIXK1SR+SLd4rvnRdXm3n9LBJ09o5pTLvHBfkuOCwKBM0X7g7tSru
UFQ2P1QRgg542fipqS9PGWNrfJ7XvcDDJPshbs8CpSvtiwwX/TEanhlTstLk
eJaWNL6Zpi7x77G89rVnbEp9DtLezdtOnVhx8Q2H8ZRTQ6g6O/dKfjaXMr26
RxC6sLtTKRBWBiK7b5Qklc1tt2KdHuYFW3cS6VrtPv10bb4bdh9rbAO8kEO3
fprA4J8GqiEvFtj7Qa9jx8RxJqO0ljJV4zWw2oYBfSXCJZdy8Jpv0H0Y+G65
KfYoSRXzGc/UT8KLYDlv7iq3YHn+xPXxXrl/dHM4NYugSFmXnrJqwUtoOGzt
3QoP9cLYVJi0+45S4tSfo6EaD+QEHjRm3UYJcAA4lIeiL553ziM5qFj5vhHH
rrsgg7iGtUoWUPx0wKKOFI1+yOYU7kvrxWiGB/4+9yjFVtTIjqD7hJ5gJJne
VK42xfNxaKEg1LM24evMIGvEV7xCGgRCauZ0J+IUgyya2q76UPs8rQPpOz2Y
cv61di7ajuzhvPzHsh6Jw+r1hbr2w5fAMhHC/DrV3pNsZAiSaqORDhqAMiIT
5qE+VuSyCEBZUGbDzfgqBSuC9y72RYamj1SNw/4BfE+WGaoVeatVrp77rpV0
NNwXLrSi2DMymmuuci1SYyJQGUJdr43SY1jJO8FYnb+bqLJXiV+zIUt36d/7
BBJ0hfo9CmxWzCEaqNYedGuiNmdMPvxU7E4U9OwtVdYYAyPLTkU03hZK1h4G
5NF5JpAFCgn5cs4YwlKuZM93i13DcewPOxeea4qoReXci1dqik5t7xwaK3DZ
s/lvTzVKSs0VBqb5CmKgz1wNHxPAQI+6k3DdWnWlyxbVftYHgcKOLEHzsePx
nAXK8SZ484aYCx4+1dnR8FNh+/pInrjGQf52BMTvMEi8sab6NFUVdV9G2Don
N+XNgLbkxCOgR5tq/C0XF+clw5gdr/mq917MkRWRsHN3xNaDPNxZQMdySt5p
7JaGHf9DNfZQXBQXjRvQjkNuhUSgwU9VpA2ga40xw+hPHBqxqsHRFSP/NNob
uL/29iBS6pcyE1/BaYT5F0Zi2vSr/MmpkQQPr2f2NzvcRx79Ls/RgeThpZTy
zkXsg0cE9i5EzCDiWV/OmquTNx+2wKsAsXY2ebCxkC0JOZZDfwmIcV12AWnw
MB36woYCzKeEwqZUlbU9ybwHku7Buz8XWPDEafaAb5kLidXqoLD0ju/QcKwR
m4VUqBzUG30SuWWjg4paObXX7bVOTGqPjHK1qoWY8yijff0qSKmlsDC2b/l5
RGOW+9CIy9biTygrPfhb3Q5MJZjUgrcX9sonh/e693X74iq9ZCy1M91NKhqq
Qg6WojZj2/8aFF+s6WphvIwnfU00PUng51ttmZ29BuwS8sGA+jp7+x2KD0ID
WCK0MFWfdO0qo3DVfbOP1l99yibutrZnVC8uI3BcBzPydcvliSzNfvjnMAPP
7+uGiDTtKId9DX0izCdthzNbPiLd0jIXtPvHQzWXTFfSa4Jg0JgHS7ZqmiAY
4WjzAq77yQsFsNdGXlyZSn+AysR3jA71w333BR5CG0EPOqM/8CycttBz9dql
KfnEjArSK5hQJWGIQMZe6YDyLaUbcANNdRKsEXd4XcX6QYNI7xq42s05Cm9+
vFGFoHP6V4w8TxBvHjlxQPlXeAdDp+iz3QhUJHDn6UH+aBUyi8fUhlRngj9T
gkP05msAiEMNPh8fvrk4f/GcadiizAdrAsN6bhqjXDXtPczpLb8uk2OkGyCt
+2e5JDKWuxpq4ADDW2aAYwzTf0eiJNzrZ4BOVCt+aPNzOiydXh91ch6a8Vrp
AoSVY230iP7CL7c9FVlOFoMflJjgx9wtnYjcWRgoKMd/zoMXnE6oobkuAJyU
rGC/5K0RKs2A9ip8/grGzYhZ4xiv9exNg68iSfGAbQPqC89nLgsbt9XDQgWY
90op/NJwOM1Kvb95PYJ184KVyGig1q5oVsUaFKv/mbhWRscqoQz8DwhIAJol
M5nzWKNq5/fBiKWl/5WLtxGadBC/fLEivYyPcYb7Gp5pfdyYwxn4Am51P6K8
uyMzqsYeSkexnHhRWFDBvg4BhxBvmPM0XqrFriw/KMKBY1WRqi5pIs8NK9Da
8+96Uunz5A6hc97IZkT9aXPxmo7+AeGXMvf+2YA+BVvf9lMy2DMWo0QVwQ6E
mVrfylxQD8buN+e68zXqldqeEd4xivC2qpK/9JBbN5AUlHKK/dtdlhuQnNmj
tgD5FsnFmxTVzARmRXzRc9YTsG//vMg53q11p2ZvtJbzzIpGOVXVC02Yug71
eX93ppgKIvcdBi8LDbQlLqZzNm2juCOarRVLbeekmb62NeDCgsN32p2m9MG3
y0Y8193P6DqTqYuY8UdCxybUC6RV2ZAEK/MSkDWNTl10TJ9bxB990ASavUp5
0wFp9mWRElzJIeqr721420s9LTlEpaZyRnhIfI4fNF+ZbHX1IGH2zjUqZnpr
QmPyzx2MXzRMoAYIsUxODXy7tJrKj7imldbGxe5MwZyiOQbEfgrUmKInM/rN
3aH+w/77I09FU/IaY3pePv2oBOTl+qWhPXQUsbK9i53EpB0Pkw8WXfjwxV2K
ufTe4E/wdgoIwm/eUnEESCfsFiCt2yLYffubFi2QC7LEaOFHe6XLzQCAwlyQ
hPu83E6iooQKXJm47y28C+ZcAcgFSjgZnZspXNBydkt9IeKJfXVYKpPqoQVQ
r07mfZbfhTfyVeuUCUOE+OktR/RSSgT/AfHxDiWDydFMgugi+zuVqg0bHqgq
dF318JgR5pXcrVYwqaYSYKKhVrwC4xGmi1oeze+sgQXHCIQeklMoZkjoL9q7
T4t+8VZwX0KELDqg86j6kFihxrngfCVxwcoQh5KqyLwhR4Ofe4+173BahZev
mND1wU1ZH7vUXSheQln9neWapM7MpXkdUqjBBx8FFd0N7CBqAoKUEIt4PIal
c+OJaqHSvcxCYcJWyEykZ8iAWBIAef3RMe8f3nm0SmmGjYQt2uNmofqP30wG
/br2JRS6JX29nGw6MREfD9ERxJz9WGNCYgV4qkq9PD/L8EWqLma5K2EpRy7D
svnC0hvP1RoKBZ4/iSAH4qSj51oN1dQLJASknGqEqggtiDjtZLN/AlNnSQqF
/Ocmnrp4cpBAf7MYA5HG9owRI/tOb8JzNeccX3eS0kQHqxXh+MOmgse7s/hm
jNY0DrZAbDGGjhPXCBbbKPkdGPK4j85KpYBsPamUm0TsKIgbxrVtjC0f6aDv
V2Eh/Wwcx3wWjbCJDukGDivr9H1L/1ZZfY7PK+m6RwJGsO7y6xG87puGvoDA
OI8yujEWeuQlauWwBcR4eZX6kKfDS1cXmCrlLAndqtqiIhadwReyiVYKAvQC
jljEH3A7zyBAey8j9OVhz9EmxxFkxFRi5f/NqgGILU3ToaZ8HRrFe0oFNTuO
2cujjQ58LckCK4xQ4VasXx+hTVqeFYrCxN+U78nwFEthXr0xa0QJcGNqMTO3
69vMkZSMVivB6n+skIDNfLXNrc7EnrotwUk0zPOYZMyBypKTzvy5cpWFtym4
2SXzf0OB4DZCj2WNdaMbUIRDoM/h80djKZYZHe12cOajDDEFRCFdxQ1A4oiY
9ddbSeKgqwk67FdvKQrX+a3dHSAjZWYN5F+wtzB7WSlt9dURtuRv/efr7TJm
CObiCfI7yJgco82Ln6jvF0fD+yAXyjyakl0ih324QOsY6DUamdNAvr+CM1Gz
UwfYbh/8/zKZbYXoCKhdEM88YdHKYx/A2fXRPpFgfdnzOCDDihMW2MP7lK1p
9WpZ3Y8Xf66E/h5QXXjIwEGh8wA2rmvZ3LaFvWsIJUzMOuxB78kp641AuCGT
ue17zRilw11xTUjLtNKIbWUlBoBuJJvtc+9lW3Cvv1zg7k4fq6SzlOO1gDjc
WOU0YfeQPmNzUHF34rOVG9PJRncIFTwSV14yaU5lkvbPB8CFLv0j8FvZtxAN
qlTnlN03zP9Ijq6fY5wddVYpUCvv+dj8rf8Xmm3nXvWKjGR8hPEPn1RQrBUE
h0ebeuxIzKzcidSGByvoiVGtW3IUQD1uPFiM/27XcoNKjYsVeMO+d1jzdAUf
ZUUDFBURgZHhAC1lfYMesrQhX842CFG6klRCxN6tF3OS49CHRrgng5J8j12G
Tk+kGp0jlmTQTik6FLi5lrJDL6ZCf6Oy3NqUJTpUYvVFuGz2zSd0vEWRkFwx
oJsYjnk7N1oipdB/zBtZn2ll76aueKLVXGqb87F7oqj00QyAC9AxYexHSH3d
34IYD9RsK/ZaKClS2FWJZWsC72pDphWP9lt6f5N3mY9IqyhC7aIcruOcEqPO
DXMZ9fOefIV323c2vOuDyAmtMyVnOSVcKxH25M5E+K/OVNQ0b+MfFxvb25uQ
3w6X5fXIP72vg82F9Jb0layz4lEq+uvwuANuCLAmCpdWk81rzJLK0jne4U5N
w13t3PRgkD+GILJUI/PMwl2MEUhfWN4mJss8pOu70ezQOJwhQoyo6NNA+ZIp
6/jaiDdl6Bb/SZLAsppTE9syrmeYQV2YEiVS2+dbWeZhz6/BalkSKOSwhfzR
H1SDFTG3BCGwETJ5Byf4WWIH5WeM1n9I5SyEzKfFKa+Gvgd6AcVvwkaVvff9
92qWzDtx0Gjigf7JQXJmAEmNLoF71UCfTOOCu3BVgTcDVSJUkd5r9TjbvscB
ry1IApfMRXqpJ7jO6T3U0yJxbEzinNIkrTznc6M/qqvDNWrgV/Uxd9f1v/KW
4Bb5VKtUwoaxuNg6S6Yvvfyf2gEbi4ANZPHqJVt32sBRWwxNe8unIykbcz3u
FMYODj6Vfjdaxqc4oNLcG4lWWg25907vX+I6JxdZGDtO35cLLgi6mvC4ZSmy
UNkRLMC4Q0qQQSqcR21fedyEY62Obwh/Y26j+Xr+YDCWS1y9Z9dE1YA21Mb6
94T2a3ffnmx1nghJYiubItwGVikF9/Gid36S39xaBPsesKXAZNovInkbzCRx
4F1owxbmCvS++nVW5IR6lyTgExGz1f1cJiiXQgeIcfuFF87JAX1VqnOJUwxB
UJeWjG36lc4RPQrZeFZCM8pETyom+d1zV2WakjjIFCbW6PhSmF5iXHH9g13k
h0N78yZ0LCJESy9y1DqoNsE9Uy0OIu8PBPmNcWvQbLAa1TCAIIB8CJ1NIqOP
ifEs7ZNX/7YjNPCaik66Mc+ybc8ceE8rPNmJvrP86BnY9vpc2JoC4+0adRDa
6n2P2wqwjPRH5zOQHEvdJC3CalPakRj7ngDcseNrqj7Xz2bl7SyPsOah4U8Q
kspQWxjMrvrKa9qV7PCq1PmpG+5fabB7KI1/yqzi1nipB34xrBkkO44DQZIH
nr4wOTsvDnKR9RwGsx76VhYkMF9qN44AM/d5QmOkU529jotfkN/OKjJG4ZJC
EeHDf6SiGAFvJ6z0GPHeW2XT+HB42Yf3uE4wBEqpQe8VtwlWBnu3a3Q3tibk
RD2IMEQ5qeBn03OPZ/w6AqL7JNonSxUyvHJ9anrceTb7VgBth96FqyZsKAvv
W7TdIKhysoy7FmVA9lpfiFH0/zlVsToWffoEFRTmsX2Vr4RL+9ZDhWUDkii5
i8m7FOLWlKpgo1+fpwM5Qbtkh7jgqCUmhKRlh8SyWaULYTLvfWQe5nbAUEte
aldO9HIf0U7plDMx52G3L5ReCo1bNvNMjCXpPNK+GJNfDONvJO4hcY4n93Dy
wJ9MvNM7j15HeQzTf4nxovaPn304tXlQ4/BAof5Dk4egVY+MvFeTOkW37225
qa22xe1QPUjOrfkvtFIeHZtUVNl1XXQz8x1aT9f7PQsW93A5PGoCrMv8OiEk
u4PIvbodrB7IE4T0LhFIrOB4+Dpe07STyrd39gkndEQKOoCG3ge++pXbPo+5
FjO8rrqNZ/BJLb01qXOHIsSrXCGA4iAu3b+87rcnUgV94LD4xmSwU8EHL3AK
s/JhBqPzHD079rUEaHDHvaJlbPVmlj5tb5uFMx737zPuxCNMyrkXhhGP/fbY
jbFZZiS0o+bcVDtLbR7dD0uATdzF32T+THExRHGvfZwmKKvc++NLfxmh7No3
u5VzX206ty9KAcciWMY6YmfsczPV8AVgXIdmJ2C2kX7vZKMA8AnfurBex8Bf
PbxkXVtGepL5pwagu9ApbYqpfqdCchTNLeifo9q8KD+rYnd4BBWddKhnqi8p
cehkEDy6BZTgntKBvSfugStFE2z0/r5qjdM/Oc6jBBIrvp1qR9mZggDLM+fm
LeWFUApfXVV57n/m6VNsVfE3TFYBbjtLSeW6GRk/T4YH2T45w+K5OGIVzdXI
QPo3SZros1Cr1lvDObgLf1ut759Pgy9FeEatGPlm6SEWDxCBAyeWE+jSXmet
P79HJ6qMMkEEInB70Tm45mhXxfcXfGEgYbNmgdNwlFVwYWvVJMRlvF4kgzYJ
C/wa4LD4spb5e455DyiESqs/N8CxykuSWg6JB2x/3Q762/yYtAfjzqmHDI4g
ZUm1l55+HmO/qff7/GbMIJfCkfVzLHEDl+99CijeiRZWIdmVN+QAwaGvymT3
On+OzkvXx98bm0s0vU+Q4efSEQyqC/zk8DrOo1085BnR78boG+YA3DoQRB7m
rASp9Nq3r1Cw2/4728xKfDW5ZeO5XEh7WmBjmRDw0fawETW9wJOJzOXqRMtG
owasLdSPT3pDhFjyFsaJyI3YeTW0sT1Ng1TjrVqQOMPJZi2/RfjZwkkEPgP8
SZ2cSJO8gX6LfzOfHD/Ck+Y3PNCUpU1BcDXcEjBLAcsP/72KaZ+HTUlCQ9KX
7LiTUPzBdYVSnGNmMr0EQGXTYXoFqzq/sSVV1TU/bdrH+eCusrICpcqT+wf9
Glyw8i/3JwCT5i+FcVmQzNow3Xn36dr2jB1tv1X6CSnflG/xYoAuPXniPpVN
3R6YaTu9wbBdxnl+JBI8U27fnL04KVARMq1GYNG0vomqiOaOf1e7ZE44ggLC
XHIrAPw15Vtz3POHQft3u1E/2Yp/W1xk22Wd+QeZBs76ASsGvUMx6XxHOX7o
tEEF/BABw/k5q01wqORrhpx5+OSOXZH35V/fr6meUvqJAC3MdKu7+m9/xx7X
c9xTJEY2IyfIr0wgsJt63odaCHkpY+lyByjixuzGEn/bEKpNm9Mpmi05/1xO
/HCCSY4X1xNu1GoJtDRwH8TMLYfcHkrr3Dba5xnUNiVXDESYs/vg+/EDnDjb
y3WY/5mNHU/b2trOxXv59k4Yp68ZY42TpGRHXoyaDhca0Ph4FvQNp7RXKxX7
u+Xj6xYZY+NdAILHf/5zKmGjzGOBuL5WTWU/+Rlb74RilBYbfx7PazRkzCJe
S+L9vUgMkgT+FQgYYjVI+T3lAhhw8TNqDbF0cwYQmZuQTaMYX1lnMjd3Fnzt
2fGH7Awuwy6UOYIg6wpPfRwRxtWIXtB9aQTZlN5SnjbZtK8lLIZsCHLhzqZ/
hmUsytQBRcU5gUMOg3zKqqbPt9PQF6g9Outb+8CSBN5dDd3DctatnOneaZtJ
728762cGAQYx0AljM/8YBf1dLeFR7a4HIyBDYCw5o/X0UKKhPXfg/vLeOIY2
til/ISnCQEHu3eQOBEEkV0A8wRHgYJ67DrCDQAmK/wsjrG5eDPE0qL+QhjIE
4sS+NA/1/zGyu+OXqa6/aLXDp5hn11Ip5YrpZb4/UZlrPfk81ytU6hfICXby
1GGKYoNdGLbyMqTCHA4DhAVY00qz7JJe8Yg/Lfy9UCHkAc09oI8W+aCz7mp1
7ttjgY5Fn2FFcTmT17A4KLpWnAjxEljAQQEe4rWrq49i8sJwwerdgPssrcte
YVNbvQxUrxU7NtIk3r5HwcFkb+x9GIMTQzTpkbcPathQqGG8jSt2pTIAIDCQ
ON/cg7dR+fHNRrj0+CsRb8V+W9suI7+f/naCI21LwiQoOiJDGtyjAqn41Qmg
PlZGdzJbrlf6jSHviF2zG/YrhrqqnX0T2HvhX4qIpsy3081Mk0UHq9tmTTrZ
8rLuksoNeM0mUz/FCPf8dvb1dkyfGeFIVtPEY1Hb5jOxXmztdis071VbPwuk
GYz3oh/yLf5Kn/Uggmp9kKS/NXKDnso6tgZgW2Xz46pl50PlgBnnTYW+FZW7
V1Jl/K0eT4vq6SYH7wKA3MCVwVtbtYbgTVmJQekX8y3658fKfa2Uyc9wHzFZ
EsSms3rDdcEfLx6Qk8U7BqRfFR39z5LrGpA1MmeONp13CVtUIdx9ePTfbNbh
B1GPd5RipiXerjz0Kod/tpYvwVXa1BdHpSe+bfZNffO7j+CESWOqm0ghKm/F
dlHkCjqmJS8Ws9DpMm95VgJ6lzgFfpXUCsNQzUcRDhY4oCXe9mMnuuNhBxGn
e7Yxj4BT6Br5EARMsZsDJ3+dt+13Q6d1PkaNr5CZQ7i1BoTTX+zUxYm3ch0u
Cikp+1g8dmwH1+jNxZI2eSl/dF2q0a9KylRyjzrKdnWbh8Cy4T+qMIelMDjR
XHty8FnWO498J7JAF0R1M2Bhpf/SFxmF6ZyiRLMaM/jwL3wA+AWpgl2zee+W
Ai1xN8ttl115DrbM1wj2hqhp5DvWvCUUZ+2VqREmr5nnJuhoPzxCYf5v2Q47
OPAVwTCIs7VWyV21x3CzML3HpyF51RMznHqaEpVslmqUejwRT3xys42tfnxy
tvIuQygaCcyOHRhT7pjwlmoEzV3CvTDudR0SPlXti8eDXanaXjIt8Jxl0LKH
PiCsP7P1mC7qoX40aY5hHY05iJWIZfUXrBaYOikfl31AsHlz34xKlGQ1V+f1
94z+IxYtC85Z3TQjezJQOeSQpOFWYRX76ByEcnEvQ6Kv/KR588b0iL7jDOGm
yb2MiY2nYXFoOeSya8yDdJhfEMs5LuD/CVOMUlXhhfF40BwpfylfD5s4hi5G
U9SbDvmM8/hmHqMcz5WazWiU6D5+JuT+YjYLXVG90d0XJwBrgheKPaWjGdvN
JMPsWaY6FZbR3NhyX3yv/sy2BGU2jauMtwCNZt6H2KQ/q6/Kq81GLLNH9d69
FjSblTvTWVAuJ1ad/RQA68SsdILyAMMba/ZStikKFi5/ti6/WL3dQyEH+UE/
/v6+Oyi6KI7kaRDzaEmTD1L9SN9AzaHByUsY4u5dZd/Zv5fj9on7K/bzsqLH
7yQt2A+yt5nbaE0rFKW1N9/hv6UMDoy5OdjPqkXyRFmq/E2WI3U4DzZ0sWxN
VlS5hZtQPVPmee9YmfMj9frBT55kbnv7S3uIoIHSUz3XZyGPm8IRDRqRIe/b
uqn4nPJrNk83R+gyUP02h1qOfNIjdfdb2KM9oRyVc+wZfDxylNhYT8/i6YbT
PlXKB0GQ73S+AURGSNB8wFkYHsedMADT4tmwWU5lQ9NSQTfhGz4ZrExGb9Uv
FOr1qUDPuoLSoPdZ/eINMXUNNE29MQLOum70ZbEM7XSnR5x47kcqZ9rBDUNp
MFlbFwlxymFEEhpzrs90y+lDbmt4njMG/qtpfGQ4RNPFUHE0MJ/FETtGwhh8
+1Dp82O0yIW9+Yx0qu4Vp6mOjbqLwFI7mnGJY1nMMme4KnqNZ5EC7YNx/e5Y
PvMNOp0+sQvM7KcyPfeGArbBZ+OASgO9gQ21LiFnMeHVNWZlZPz34myC6kaB
zttooREOuyBd3QFdaqW2V7Jv9B9xgu81Ye+ZW48Tp92a4O8899BUJr0MSXn4
gpfWVdIx+o/VDbjJbPCYVi4JiNGI6jLv4nW04itxYa1nZkG87wbc7gK1SZMw
NmKm4pjsvG/tFFiBOGkxqlGFHfLON+PuCBUL+BOFtu8uWaVRli8OvhDp/xt0
AxloBGs9g9u+VEnj1jae8irtaNaiNFHjI/3QxRhvuezb0CzhH1gw9XJ9WCYK
I580FOD+hr2RuuPX5CvR6VNv5UcvrbN1vhwDePkAVaorI95osfzl9yrXEJLX
+7ydWs7om8XALFBWZNJ/L7rZTVmshxGypbvJ2w7Peq8RuZS+mBriP7KKpL9Q
5OuAbEKQZ1FBoA7NN6OlyBBQQOAeX83E68g4rJD3uhe2pb8/X6h+hfMQmyJo
rJuyhBmsoM//nksCKpUVpU2dS2KAvpirMtb/RMZf5vQ8unWT1L4/zrYvavy3
r/3e7QMcBA6qoM4vCN4uAaDoe9aelgf3QJIdvzz33hwF2BF47fvM5HccKaVX
ty77upgRetOVTH8bMpGKN/lx/3Ypw5HzdcjPZNIZsXEMBHDYbqS24aL/shy/
tM7I4dHARCu+/dB0QyA2EBO51ARfkX7LqoM9kj0z9uWwC9oeiCag+rTuG8Xp
MdU5pOWBK5uzOOiu3SNqWQc07pQbYl9oHfITnRvdnImZDdmTIhmF/QpIJr5a
uyxPUOXT+TFMeOyLF1DvsDDP56cHQf0tr3JJnV/oAApgK7+7cwAYjRkl+KiK
8Jivem+qIUmo/eSCEzgaTqX+WFOcnShR6uvxteaBHkLgAgxZX/OpAI3QDu8S
b/8p/mzcJ0bJX8ohobH5mzLn0cjlFx/XcL4wYLFyMJLAn0YTvOX6XH9k//Ab
Ms/zj0+Y2GYsBQeLzhOa7dZBTwtKPj5wTOfax+ielSCegf1A8eg9ASvCuQfz
edpelAssKWqyKDv01X8zZOF5SGr7lIKoJ1xWllLW7MnZsQD4UjGG4gbjLORa
NE6QGttBN0emfmV9B6hgNYOOZLVH/3t/JqZRkbihsak3oH41lTQAAxjFWvko
4lJQwte+B51l1RyI7rM9kdzAgk8PChiZ16eBj5fIhvtnVQ+71cPh+Hehtd0z
iCLiNQyEmwghTeRTyWPrJCvfrcPmzlcMAuruDKXkyzjqDzSr8kIyfPFZEGil
h7tBJstXygsN/ErEzAfI2TIFKgLOL6HQz7B1uIHuQqwGZCw6MUzCeFufQaYj
+OjBnG0l9xMt1bAJl+wVvHvTgVyNoRfbPM1tgCfCesvan2ttmf+ghDReAhEk
6MroKBFwJSgHAfa9I5QMdMvwVBfX2Ed93ESNDZ33B2Nn67U0WbwfuPqomPSN
ObG5StFXWeyuwCipQ/4pK+PLQbU9RZAaemzEtNrwV4wC03TW1S/G2zbJy2wt
iFbNMNcwB5O9GLFotzpIahUutQr2GmelJI4nY4WorZ6usjGTM92dVgVjHAZ6
SOA51heXQSerJr2l6aGxFjK0E3tWzhnfZ/HtGv80qjAQcHBcrFT3ZKDngBa7
y4HF4DeFeDgl8oR6OFfbqSrPAvMKH5A28IpPrPRNLdWi37w2EqVTVSXZTW8U
OlNgvwdpabuqQP9ZjoaMCj8y5llcozW1ivT9VlWaXS5/wvO/aOg2N1Noj5Rf
GkYj2FQWF1srdclRlcJIJstOhg65IVINxjuSd+2siGwzJzB7P3r6LVtp4HIa
nA4kRm+7S/iRL038Cr6NUJNDlAMoZQN0mt6ft8a3H695ySbHHjSzycNRy3iP
A54p95mxvxGDIiGdGMdJXD1pR1jfvJVaKCiQjQvxdJoX9ZSVIMEZrOJXkWyx
6qKT+E8hF9b6RHw5HdSPvYpm+N4BbizewEj3g1ZqvCqPm6gJ8svifidGJnwV
Xi4BKjhx/Geh9Kp6mLP2XLj2aVsd11TA+LnEAjWtXd+02w7TCOGo7TP9C5ko
R/oYeD3ePTXNfx9vaQJtXOsa0o4XogzT6dOnYtJmiGcpW0Hk6f1mnllbRqCI
l7XSycNJ9JL3Tm+HnC0vJYACg2ASsxGIaQh7jGZ/ZahT6UtgGaceydEKB5Nf
HgasVOkTw3/hMy4rqkzKDuG4bYjSAgk8bu7q2cxv3AuRZC4vA7v3yRFvH1ZR
rtJLpUWcALuYzbpyyVVEuCIdLaPUGclpB7lb8y9xS+K1G+5dEKJquvLDIB+O
SU+RQLGiCSP+chLDvoLRB+kKxI/pvPyyqMiLSmq5uFaaUpqw8/nYbosLdNbx
6VsOLO7gQ+yCg9+HIkvw3Ct1OkfIxgEFM/p1Lger+4+wP+XPISb0vE7Oqm5m
fdIFFnyVPgIEYnCfB6n9cPEWNlRl8ig9nWn6O+O1XGeMZMhC2gvWuqT8kibh
v9Ku39gd+XXXJCdEJ3uD0F320h5ki07R6ngPH3y2LB10cWIlYZW+z+p0N1xr
l/MgPgyZ6qjzms6qWRu0CggZ3OfmtwEP1M+/zm5Gc5ychyAhBpJ2bS5387Fi
/R8crUbNDQz2FDxfT7mw/pUH5tN5q2SQZlJHFk5FdzJCJzXiVJEuUhoIARLa
dZVrHjGE2awwwpZR/UUR+VRHAKD5YDONKEAmUuCjkW+2NLfor9UqTdNtRYsC
d6ynoRtZ277P+U0X5bA4RTD4UwYwMwgjileR1B8mTYTuKI0Jwu1OqnjzGgM8
nETxu3PNOakcdBzCSKguhPt827JRs/0f244ncw001Tipe5CJPLBfk6haEKTQ
rIXa/1IsSQRbuM5VFMEId2abuGBn6wC1ooF+03oTJ/d3jyLs0VjzR+Nc8ush
HO34TKaCcHwU/IOnK5wH6qpPE1KvczbPeSmh6YN26SwgoMEHjtjESo0wcCuu
jOiF24bhIU0yNCQ4xDLFs7lHj3BPmxWEsqG5iA6t6qxBhjCbsS1y4KAA5lVW
9Qn0kESbv12LwenvPqR0zbJ8CDf1DAYEU2xeYIh/4urMGe0rhe2EQMHciZLO
5ck+PbkDm1cgdCei20WXG/5F86f09Fr/2WKsxVVBYQ+Kue3ozV0CzprhcLdw
URUZ26gVxhqHlcHFFIvGr0eWjU1VppleE9q65JnSVrRiJhIKSSqTUjoivEd7
aY8ybkj/6SnVQF3kBKwIZSPDZT+oe5+zYPJeEKkAkys0H8maAlGA9ZJ3V+eo
f6YNujbN4oxeMtbYo5nwNIU2LP5AI3JoKP3gc30D9WwEN+xrkgKdC9UuAJyx
0okZFg00h/KnddS8oD1mK88GjU738C8c9iII18cwWG1m9weMcKpXiJwXxl8G
TMu4/inO8i7joTzluGdMbgLGzOS4/L2ega9PXUMP4Lk7+EVqXHNWLm86nnr1
F1UifqW5caF5SIcLeQOO//m5vNDOPiJCgSwcDhz5JlT69tW4wTy3ZOByC1oQ
ke8p1P9nCa4gOCwidSoAB2vpQNeSuAHu8yEhTkxUiLo7XmtU4pAkhxNQv7KE
vy4Knt5vjY9KqXsQFYyqHvOA0nBmVNX/JGuVmO/S89y8Q1CdluaVmCgW23N7
lsRuxjVFJgKkdrTaxqKDz5EvW0KYMUwE5qq1VhGbFaCA7LLReCFDT7Ub5kge
wKic1geIbeTKxs003kbt59wV0Zo7lY5e1T2yqjdIu78ShtqQD9TjxBwRt4rs
Inu4v1+SLHdYi/Fa+1YxoqxTkuKLT34tuzMGyNOI5485onKd67fH9LUxohXm
sWs1FqZnkjed319h2CPdR92D4UfhUqIvD6NgdkW+soy4bu0Dpw4i4jQ8ygNz
da4fW+bltyLRBNMPKMgIuDDfix1QIevacn3jEXNTHyu421VLBpiEKTh5dqzr
LZeE9lf57mb1eapVEjob0X+6Tm+vszGtvErmNtH8F6Pimov/w4X3sYudvynf
Ax75cUlB4V7TS4TPTfB1FUqOPiqJitsKTAUROd7dpcV3aSlMIQzlQk880z75
NuBiobfBTmd1WXhlJ3l7Ez87vDbEdmjRl9z/Ni1vTI9f/fyDDtwx9SP0gn7g
r42Ci52G5lSNMNrWrKGayk6F7PbmY4Og+maXkn4J1+05pgUXaaoe1mKNj/hR
kBCPUHEqeMZ02fCDM4qi04GDvB98/kDurQFCHsqql78IfXsnQg4F2VmLtD7L
Ift4D+Hkahyps5BMmfSnDAefsbL4dF+hA3NI0gQbEm5xgt5BskR6NRR/59ab
NBVHQ3mU31iffHJsk8Xti4XMsk2mgLvdolxYbFbd4cTmwYKAu/R5tYZIWjBp
1B7j0zdwCKExqaIhjICP0kxkhsc10vjclT2tP93txu4XogO5sC93amxE9CZ4
z12sUxFw69vb94A2O9Tj9JZ1VoBJ+LGmmXZqFD/ZfU3AcZ4r/+BieMOoAU7Y
m1A2rs64fRegpfeUWcOO1zv9s8GdwJZLOBY0+70m591T28svlVgb+pPmZP9n
YUdWjyDOF2zytJ/iWn8cHkM6p6zItcdLgHXXmR1L0Gel0uR8rY66v0AUdMil
9YExoo8UChF+/aH0LKib4rdFsTXC/yH5KgNnRQVZBBTc6wIp8ujYs9Z2h211
DPM26/VEmZebNjX5THbXu2lo/K6ApxiH+yptm70Drwuf1Zk22EY1Q2Fqcwap
D3aG2pTLr1qlKI3X7v2abDBj5ofghk8JcxJFGPEusHxH48Tys+qUYjsjtt2A
RXtf3Nndwri3SiF7i5GcChFLIC9fnU7RlGL/tGaK53E/BxYgHvvzJveuzDdm
8hi+Off+FxzKm85pGC0y0EnPqvbH4dcPuoQBaet8QSrxnvyQCmEDize82Aaw
SXbtYGcdDOfh0mP3zvgX1i/GfowdP5CjrvDOk6lr1dyG6x+lfBov5pgU07cs
rlsta48C8aZ2ES6VZHBIrywOw/H5DuIJUSLlq2d9x8+mBSfoAumaLzwZaKD1
m6KoTizQ8BpGoZl4l927RQzqZJR3M1l0RJkorC7781XcGOQ9vX+NSN2Sac8Z
YPjIoIVxYA3SnzCoTC+il1TjIRoh7BquHQN3w4U9isLPKftCgLSjeGYCIdYr
3vpZlpdp5/z0pwFZzdcSWgjc+JG4Vz9xx5KiHh7UGD4uLdMe+Z6T7Fu1wdvX
laRIEWE4GhaV1sCJK/riTw0/kmk0GIYd/OtX4sYexADoJEEfE9azz/lJSgf7
7Y7lVjiFXWD2mIgP1qdpk0t1yPs3OIRj5gUYXUhCA309x0NyjNuxHOR9pfnv
LkoEBGlTDlkhWDMpeRp5STfKE5zQ6Cd0xWcZSj+MSOHuUEZy/nYDsq2LJi0o
DQ1zSA+vN6D5VHoB1xXwp1frn65tyT3YYLksbqwy1LCrTsNZyISMj3RWjOK+
+/Er3GF5HeNyXP9NSctuGcCOjTsABfaOBmSsg2WHMSNZDVGNcO999Nr4c526
qEI1wcvYhFOmvY5kW2prUa6tSGAiQKhO0FECmlbQAKsU4b6H0mS2oglibIkJ
N1KSBMNTWxInx8yr0ZlhvPP7awxKy3pc8Ip3PqkiyDNlKmdJUw3m4par9JBT
nWzooOLYzmC5yujEmfei6DqZJpZoGul8EQ9+9+cgsHwidlo1tYlko0I1bd3H
N1oXgw+HQ6KWEogPX+GRnpPmNLREQ+UGO7mIscFZqiVRK4X5l6J/XeGLAas4
timlQLnT2ilLwDr0QrNEk94b/ZdycYaxmwGR+L/z9PCZl3SRq4RRTWMOENSn
tVdhIlfmruCQT6yOKe7JWHwem1fbH0FrVXDgbEJBpzrW1nzQm5+uhQVtmF7X
xlh2BYmeQcgIpPARhEBjsE3U8ZjFQUA43TBi/Zms7GDB3Ll7zAmTMCS7nvlg
irWrrNvEnQ2eopvMUgTaiFEWyda9e7euu/iAhvAldXg5p8n/WNd8sfwWnS8a
6eASpm32mDOewp2JBKq4TbBknktartdELRay1xmrEi0vnWDUXJgvei00MiPC
vYsWhk+BrTHcKRu25LPNWCMOw8OijdXKED76FzYWlskroi33dXu5NZRcZ50J
XfEuOxywNURXplg6uk5V9OHi7ewgAoYkZNOR9sZFi8s8+4QIWYn8WLC/OnYy
kXSXjCtdaxmm/+xz0kQnQUm5Dz2tpp79RbpcbXJ4fnW0B7XhwCQEDZwFuATq
oIUMeEHelvZ98JShK1RMgMXI8xr2dVLb1k9BiifbZLWdJSCA7dSihe1Mt8bY
QXOkpCBF6XBkPRHJ5D6WF98vTaJrqt84i5T4AJECGYYllXTdU0lkhUyEYmM9
djAXmFsK8f1NuakkNivvfMLSN/WlRqCg0Ui62gHlLQTO0rMSWZ8JNXm9eAu7
1UkOX7pa7ER+lIt9wE1afH2yEYbw2LQsqLPpTwf77IZjhRbuT89Ke0bFbzKj
k4xuXXEizzV5HbTWdW0mXZYFdqVvZ+ghDb8JUflkv+FJjXzhWC6LpsUgbAng
eNHfDZzflHZrrHAjDfPUAbQ5YKuFhez6Om90xwuMQb0+g1iooak1+NJ+fn3p
4rf3lbaoxyUK3UdCXYPLP5bHzMcgIHMe5qok7DM3+BPck7awXLe1jtgnjTud
jSXA2WtyzYsJkZJaT93PylFfIHQLHn4L1npu0dHS6/Si3YMLoMyYdvQoWemQ
h3cRBR6XsuOwV9cEkpcVH1moUQLARAvIHLi0mR8NqdEzlTbHg6zI88IvO873
Yh0E6wjUk574bHEIpMmUkcJObdYIiTARJpusYYiGFljM/X00GVPjIm0Y8ojl
7WimzKzOh3j9NIM3qQJtv4zHynnjOmcLjS4fMNzRpJYYNq0j663Xmczk+f39
HtInp+vcgdCm34r/yZWn5W9f4zQJVCNQfIObCz+PSgUITEWl7GI8dOqVxgfl
xMeUfXOw/LwFhxEBPZPN7AUyXCKU7hLarUgiemDBIBTdYTrC6aCNdjRx53sU
XDTxNEhKkkoG17RmHqWbvjoUSf0CqwtHk9+vAoeWboAPicZhjwIgQATkKLgq
Zd5h3LgYt58D3zv5zFPigINJva4dmwnRomDiYqWk7/eeCTlh4Y9GAkbfs4gL
A2aUPhR9tlH3FuPNZLPrJYFpwc3m+5GXSci5wSpkOJSvu5xEkwIQBtnp/90b
SSiZYkLZhoylNubZhzN8fate5cmQlV120RdMJQmo8lLRJt8frjqmVwIViOOq
8KwG9g58IPxTQfGFywcwO/SsR8ukRy8Uh0y89F7QqK/kGcspPfF30qK/0Veu
ntS07ld7QDXneLeGud+Z9bITwg7kZZSwIxKbZ1/ZwBIEcSRNigiqlRxRw5Dx
M4s+jNe+pD404fgqGkPKJu+hx6PW4CRKlsNCWOPp8gBU4uggCD8uVotBmbmQ
LonurQr2cVnXXiz5tFUs8ySquWXCzh3TV+0ymErIkjVu0hgySmbBRkbJ8yzT
PVJvSauvnYhZNhA9bxS6bi5Zl0YjZ56Uh37dTDVFUwknQ27F6Pgeb4uDUY+L
+xdzBQi9j6h4o/cTeCo0wyo9xQQXkR5mgEg/E3iG042Ip9jKrp/4na+kGiLS
F7LKxZpH/JOyuNZ7I0WqMMW+BUGH326zgaA4CR1BvnXLtBhsNUP8NwtIw6Tr
DB2ZHTvKgoea5G9DF/nAKvJ0SjM+e1OSbKbWziyNHKr8cOTNS0UK4nBCWeDo
LB9sqXuWs69ylKZFptz9ToeVnKKbn791ffkmDAWdZi4KEuHJSEgoumFX4J62
92szJIT3tI+AaBAw1pewnTDDjJzQ6amDzPEok95VdAwuRwnD1SAzJF5xY80s
UEPqydtRscy2dA7N5fz2oiQRwi5AGhlo14fFeGYk9ZJGjtsPiryPqlH6UiFi
osha92YIolHCGQMn4XS8Snfvh9Ce78PKRzRhtufU8YzRtA7RqCR1XB3uvUaR
0Nz1oP6E968yZDSqXoKmRGgREPYDCS0eUgE5wM8Kc7hWnWGULixnmhBOxXW5
ubDg8+4f0h4zZtOXpYIWSImF9nPH8QNJc38xc2S2bpqpL6edXUhmTurdZeDk
6+gwP+Wnk2GIKcXI7aWO0cSKTvSuV/ba/o4Caq1o/HrWK3FMOO7t0CG/UHuC
A9vcc94Nt+McuPv8XcM+8BwF81WwX0jGmZ+ahLXMTEtc74BdXDO2ZB+Savrn
irxaV4z7qJREy9Kb74wP1rlSgCv9uziUIsJw5njWw02jHqNeTZO5/jgSwBb0
d7rm+9NxlYqw4Mezt3kMjbjCHPLzdq2uMFmd8HDNKc0f80m1+Fj2ufhzHsMb
2xHoAyTt2auLZwe6RrCr4JULWPCEh8/ucCNwA5hTnkMER3LTxKl5l+adl1hx
Bj6DUPdeqVQj3fE01ws2kqtcz9YzrqE0RErVhr8k4rA8jnWAnUiQN3nXmbNi
xXRa9VKjVOXuft3aw+lkzGPI/TUARPF3SEk8KL/Y8U7MY6cMCZ0up1jDO75H
aSIU2Wqx2DoLWtsxxTMZ4+x95PVSpCwHpKqShUi4OfH+8kZfmRlGyPXdW20J
PHpWtVX+YzwDVytqF8bJwM2p6hmTVv5p5CfItH0xwfxM9yuSPO5Rlv1FGyIs
3ovkjl3U558QKz9EWkhDwN39NMI38vvETGpyjsVHzkWqyavRSqqHQkGNGwt+
yASDBU3oSdx2iBlWih9VR2Jq0YH87/bBLlgrpdyM/jTJ/vSbhn0Y/vkWCQ+r
RhgmdQ0+WLkogc54+r2TM9LhLbIIXReWX4gkSeLdoDKW7mkW1KHPsVwaR1zS
9LpIWTT0hKVb7aHxnbCwS3DD0SPUFTI8VWLDi2fo5Oz+uD4g8ukdvE5cEH5Z
IbZF0WA026pC+pTqjI87y+h8sAp10kr3nCVwWkfMJgCnhR1eLfJs6dj5/xex
YVPdozOOQvfqePMh7osbQnESg0nlntRqaNB5qlMBYUwvvyOZvXXDXbKmXR8L
Zr+V/HB0o5jedkPe6p8GM37h8HDOvjMPmVIurNo269DZFfSvc0Cp2//UMnRu
V41dgZhAtcARioP1O7cGAhHZns5S5mUJDBCNBEdIjMDKZ9As+DaPocIJ0TLz
tY0e4aRQkmBc4Ht++5EojqTVPmjmrIfVskmBCwXbafm8ruON6YaTwr34QH20
Y1M6E5CUAR0ExAYQDIPlGhyqpgBeSWTutr6xun32SjYi82sW0Nz22rkneRIq
JHmAuJ73XZsWHocPV6BWyi3ZU2UT8pSjDlKo2CaXS/5bwWRaiaKBdPRFZkpy
FT6FhiPfHva/pRcGRq7RmW5ERqdi9v/D8Wpg6/KvbEcC/iCERugPvjiifncq
PIiRCkScg59iSJkVn78P7snHmW4RnbZ4E5ftQvD15BzBU4QEoIiPP7Yjjrde
JKGk5kmdyN9bFH5R8enhMNmITzTp7bsGKu+CMmHdvoH7nUIpnQ0/lW9pLIWl
W0GxOAuYryeUYy1CRfvSU24BrxSCLZj8L4EwdCmp8vAAGYAQd+XFhDpX/AxT
cFAPvbDcFRYhwzKYTEJlZojSKD6LRnnMLjVkBjcKplR3FXxphenYvU+LvRYT
OIDMUMjCBFCR0zknIugdKau3uU6JQLu0+Zege5+jWOBIumJ/lX+pVgV7k5ul
QEl+blU8ER7STi1w7QWKX8BTECWWXx6dsuN/k8I/0EbQjkAhfW5vT6hcWmAY
HFbd8jUe7+NXe2MHPbK6BWG9GvnlYkR2FqhS+v1F8eb/jirCvNtJ6m5gI/YO
z5yIKPijv/JgJiRUzkI9wfxnXz7EUow8c5psQAfJnHPCO5dBMjtuh4nsT3KB
K5FUbo8S7KAuuUmZzMrB7w6h5Apfca2XE+kw1Zcj1vDHKlBTs37/Pnc5FSB5
r5Uae1mv5mcqtBg3EQ0Y+6Bh69Cpu6PGawCL6XJCeGgjW/N38mBa3Rhj6Zev
XCGWs2ODnBtjQfPRzr7cVWRbFIg9qtWoQyqHgyk92qozAhYzNMfoUWHtwRAX
kVRhDcyuXTLf5DMMGNLPXWDFAr1dPHHAV6Xst50bQVoQ0PjqzKVOyF929eSR
C1l62GoKQRZ7BPoEdhI4mfk3slbTlH8QsgMFRlNHP339HlO5cRUAmxAPnydq
TE7QQS4RK8njm58L7v7KAOECFqCJxtdv3DUinBtCHQ8XxWjP75U9OAr3NM3p
9eWPBE5LY1D7tM2Wf2v8TokmtxXzAEgRZwNf5CwX2wWg1nipbFQQADocrmP7
3TemIxdvU8jBIFvM4/k3Eva6XA/TKdx1DOloEv+8QjSGamAil1qnN/ofOVCP
0LPzfx8yuofpeIPjldne5wxCRuHbukdagN9OGgXYRw7aesbJHpnDc8acIqVX
ON50P7A6QCsQFr4zU9gfg+TKqcz/dRh81Pw3GLGieDl/c4pNfXjc7gcT25FI
UsEBtyoVeE0EY0lHmvzdBQ8PgWcJJael8B18Vtu7rqe21O2g1zKKcPFVptDB
BfDGuayfZ/VakcO0leDm6qpI8GQ+QUZH7OaM/eightDBUHC8t977/fgrSTfG
lMVEN35UCiYR6UB47NWHBhF/XP7gHZZBqTbiObKai8LBiTgvGzA+tz1KsjCq
e8U0RjHloVioTRwXk+fACPeMWvwDHEv8ZxyPzd69Jy7Lm88fmn0iXjJqkv5B
bCRmHj9IhjBPdpp38RjfuaIRNPOGhUx2je8o2w5K2F1DvYwl0apcTzTcGQAn
juWa3kfAMNhZ0t9W9w5tN86azycx2GMCClMQUzF7MbBmATmYTv/kaG5E6TSR
j9XLQmm6ozwonN8hj14i5t1+uAu78BbSzoieSzC4TGaNapDghp/TELyjNZTb
ojBV2PFE5g62FLIhQ2u4TCd2TkpkiGv3BOx4wp9LafMk1k/TjOyGLEkvCcjK
aBb5JUHgWXJoGUXjgrGPax7KdGytPLrJVCE5GcYvrqoH622lXceLJAsIyWuj
TMYR9W4NYgWpO9n8rzqpH6uHwZGzgXyhpEKSWdWFdnFETkPDc12Lmg/56aTx
/92ifjFXi/MbUnhaUbV+9imhDXVOhZ/zpDYTXgblKU65hFa4QICHr+wlHnMR
S+qb627Y7bw3kcRuJJlPD43t6JbkZuBQgpeDcfh42XDObmGjOgNRQagwxzRY
KNETTfhcfWTcZi0+5WXm7dSX3mHhe82geLWBIc4olnU9lUi09w9Wa882rq3C
25MjuOgtPEX8dHAcp3Talr1Ts3w2xnExNm6XszfaRzU+JyVG6hwGpoUWkPYI
X+OgNJzpgONKCeSqNO9zE1+YC/7NxpWUDkVThhu4hpiZcHxS0eyVmNpmsMnk
7hLm3kMHuxHajrhv6CPf2RxnCz3mcSZqv38aJOP/UGONrJ0cDMl2QX17cR81
FRpUCvx6R80e9+glCogm15E4HKwmmKVigRXVvW3EuknU49K0s0XH1bS78Wfx
T2ulMFTyvoV6SVv8sHXfGsDDSq7mfVJFz4T2N6Q9JfJGjsPfEBYk74iq8sC1
ez20YENlC3M/XxsQjP/CqTg+DW3gaHs6bX4Ob8nIVmiCpDyuAHM6xbHINSRI
cOP4yBo947NzftgmuSrrYji+uUqmr74dvJ9KTpMG2J1pDq+i5CTu7vpLrAok
LX6zmb5RtS67RoB3oN7Cj6tR0otTWhDDVNF2chvnsuhot5iC/YYtiG3F7Fww
uzKauozwaEl5TCNW9bUGsR2yo+aDTCAKa54zSX5K19gkPbpH4xQxhMhIHu5p
nL1Hul3YAAbqli7oJFxRERJHejQohTxhxmZM7+M7pWEtfrdKuwmfBR25KglN
hbbS94gcZ5wfJY74QCoIptX2fUL0TzvLzlyTrLLLUeLM3l8fnuQ/TZIqdwHO
AwwtiPXeQ1WBZPLzn9fZuSCQe5qxZPx6VwYJIuoJ7I9QeRfcxTA8EdL9f4iG
tlOggl40hnDNbCxjbpZtoXhGa4enhkW5j2cxKd9HxX1JOCxSaMvSbvbfHjaT
3LT3w/fgmUaSU9SrlSDk+1kZSlINWCHISitdVRb5ZZ7EdKf3mW3zQICGGKqt
D92nOW5dwOjw/ENHi83OAGzIfXPIs9UYQcZe2EQ6T5lfbEnrEO3qf/eCs0OE
x8Xa2Ep+b7gP9tKbe+Xk4RxUHu1k8Bm06mOu9m28r9uewTvEtbJVYZ/jQrxb
xl5Q4DT5+w7sTezCfD7ZJjY5sONIolJUKuUb5qZ8kjbMJ4B7xTow/kKLdcmx
z4JTuxOPxl2sVRzQSSfjtpBB2UQZATHbNYZTzIaBnPuuG/A/sMfFazBQ9RkR
Y/vRMTgVs4i36TWjCcQN5mKwohnadKSBH3KEwfE6BxyfruTZLlkcmcfYjs3d
+WPD0zSAp0i9zTUJV03K50qc3EMOQ3/MxUpZ+9pb2mF+i4aHBk9SOliRaDwZ
ioPs+7eTnqCGtBfusxqJ7WvgLPwBksnD980OKA7RaDKEua7NCHzY2qWdt8NX
5+mRuWrn68JXWvmRWiNMCR2VU7q2P+JQO1hp/WayImmCgjknclhEDQYkE6gG
BRaW3h8yD+2rbsICUZ7l2Qdef11HvvjSxjZjbme0GOgBEMbVHwk/pOyHnl8z
y6YL1KMSzLAwrJh0o6Fn/yeHiUtXf0Nd+SrJ24HFakaXfdqPnB5qScvmM1Hm
+pSHlfGISoIHvs7rRFC0kF5QuFD2DhmKm1Z3JAnYVjl1bjUD4xYknOaagPYi
xCcbMS/qEVfmaLjPPfWOCghibf2dhdUXB8471Nq4CRitVdBRxsXZPgkRXAXO
DH4nc8AVlEDgV8mslPtIWsnd6M5ZAmjv6OVexKalq3uhvXEv+4tiJrELd4MY
5XgQRD6CUwPfr/mu4NL9MjusjUqQ39KLmM1G0y7l8lYZZ+mi2pALbaUM0JDo
DyPcUfSKuLOCVcV8xbp/RqLTNdsBoKAea2BZRokKH3pI0EtA+ObtHM6HH/2z
XwiHz6w+Fd2QVbzrp0n+dfSxhcoPy3Itd6W77cBfma95/iCdbPJjVPvm5BIC
IMtUqERYMbz96znXe/pr/XsuLChDPjqf9wCcxaler6oRD+BM8qkPmWHQKWHP
VSTYTxwIt/uRLnO4g257KjfTyAl57kEIcixVSN1z/cWUIScs7r4HGKgtIrN8
uXcOJ0+6ieDvY8jhL2Nghj/HFP5Kly6z5VuXgqazWgPFQRXN6CF09njwaRpI
Jkyg112sS3Oad46eB8qLS/WMepuQCAsZpTUj/SQrLBixPJOkgDkDb1yyESrM
1hTC5X9JmRrdgOVs6cYZa8oVM1/WuDVoq+pJbMC2iBzXLns1skQi4uUJ21Qu
PbCeNlSlP1AeB25h6YSqylQgkw6crh5LT97iBooJ88YvlUraaZk5IZoVHdy8
hAJWUiBpR1oAPRYCJvxTBmsksXf0cTH/jWwtxIHA1cHfv+1huaL7+djE1VEs
4J39UVaYmFOlZaYJanSJMeq29lwhAVW0FFffg0lD1VEmlDVzsILEMEAWxfO1
oekx1+luisNO2V/zxjHTupGHEbj8314EjD88JPAqqDgdQz6Yf5PpLSrJXvXI
d6vewbAKRyYVkREjN8PhxFkAxiLkPdfgPgo5twljYhQLsrQIsV9WPYVOOZfo
5Ks6HRQYVAFJyVMUhipGp7TX0Aj7yJip9eOde3nFDlwqf98j4LeBN7PzzaaX
07+xtRWJO5IBmf6lVk/tO68F2ZvkWfMhw0xykJB/Spfb2nMnmslPcXbdlwZT
LMVQHAZwO5rVfuhCCqH9gfhzXEYrZ89wxaUS688Ep0Vd6+XR+BBRwSVOgXdS
JfqIhyRXen9WICRT531p86EansV1iISf5wGiobPVXJBPrjbz+/5RhstPZOjb
rw75qTfcvKXqxb2HDr9bAyTm7eymB9BX7OyEhog4IE0Zi5tWkwdajuIIIIkw
Rd8sUWfWzt7EZ+r4Klm1Ib2H7dAKzGMHFCwjkVDnXjmHWSIQiumo+AYIk/Px
WRIcyzKKI1xxqrDJxf93OgnKdI8VBnrm6lpfoBf+r9Rdnq1uHpRoFZM1M5fC
iHTb76/0YvuX7Xb+Lpi3KGisFxD8r0unR3BVzd/Izcmb7nOljOEDsi4Ite+s
f5SeyuEkg/qh2zPEizzWTNBbITBUFcyxzc8xnXDWa1SSBokzvCkAmMC1OI1B
wlJooqi0sWM6uKvdTEF8ffyNvwkk5LAKvsbiCK5mJ8CrT/S616nYaivioXLr
3mRWf8htv7Vxlk1IkvM9U1XNL9SE5TiMcIJoEMm7QkT+6SHDe200aKa1xSkD
0Wp15b08LOib+t9ex+iDPGP/xHEpNKfWoFEohPL2xwLrXOBdsmB3MVcSQuPw
+z+6A1qSCTZj1cA2Ug7KgFOlkylWkBw9OQIVstrKvX7KM40F104lUWKu8n2S
PDUDq35eyBZCBqM2OmVO+bn3Fg87majsztu8cBPUzoBr/7YhprZQpb3ux8SV
SnC/zjN6rWvKjZTV5dBvJJ+YEST6VgvtWvUPGiwfh3B+tqhiy4aljqOYd089
Llzyc0LVNqoVWSL2qNENUH6mq+hU4SOBWKzl7VSwul2dQfBAiwhoqkm33Pp6
EmFZ44F+8pZyvVa56W4v4HUCB1LD3Yr9aTEPJLD+6Vn4wRcuCbmCkbEsG00e
iMIPgQr//Sdfn9IAMLiDA/HYCvc8XVdUA3N+doghjmOzCLF75L+d4jml0Gsi
qjAdRYy8AI5fdaYN/b4We/xiKykXVG9OmiVE/rW0Umn3FyflJgKP3IdPU5W1
u7K8CmI+H/553sU5Qb3TX2b42EKjK1vfFkvI5wgyOJsNV34LcKoa91Ag1KRu
3hbdmu8s9aeEFrNJhEdY7SNkvymk+q0iW/uv/s63KFiXuM4CLXKKWWpOdB76
ugzn4kWeobJ+YO8IEm5uGG7KVifEwT42F7RFfomgZhW/hbE/m7B+KjgURuqB
OO92ztOOdqytJt+79+1T8rNaJMR/OmY8JhzVay/HVjDoWuPvliyjXseHVBht
uyuCSBZ+OwQvhtXYsO9XiVd2/1OXaz++zVGlsIkG5hRHD81BShGe/Ji/wtGi
PoietvrYSowN8AMFPBWspaH9bIK6rj5TfUPvmkIn6wqEorJ6iQSYyaIowLH6
OimiAV12Tz9APpCJyZCyggMBOa8v0L9QCzr4Sxwpt1t40/vjBypNhjhcOug5
5rI+khDQJY+9IG1M8PCqe7Uvh9i4KolKm9wS4zLXBw/cbM0qAxLVhzw+cy9+
55Oi/G1cVi6qO+R0ghg9KRGHlWImCNGu5UAqzSmA67jf2Vcd4k55mRvgp/7b
pWCbo4r5RNJp+2z/pcn9rJaYobKqhfbhNkyy+keTIvzT8iwBgSoVaNV/47iR
iyDi0gTzDOZLGl6s3HTxtkPoV4rv7gF5uACtbG3t0FOuNJ749PkgCya56sSy
c1Xn5s69YTz/85J5poLMiCjMl09yQ5sHKlCEmVLlF+pK6aLt+6hmNjnCcGUM
ClVVR8MRHwyh1elW6jHBlzo66yF5Tk7WuQghFtBADneG4t4ml05O8ia2GVc1
RcM2UCZ2ZTLEvkY9trx2IOHT4S9G1O7NPCk0bncCt0IECVA83HGHp1BwuJO7
fCCBlbHV4Kf5f2h0G3rsxXZDIT9txL6zEbEIhchS6aTyMC8QEQuPj41Y2dpU
xpYeFmSbn5Jti1hBYhHPLsTTrwhzEs3nwf+9qFbLGH6FwBHLEr0fB3yhB8Ha
GH3AB9nVVM+8MvmpeE/g88ldt49qHBp5Ev7IcI/4HeMzEThFxX0yEURfKiB0
obAYPwZCP89b7bfSY0C9FpX0mUCR0u2i1pNg503XH1wgxT5f2FYTaOzg+K0r
KKB1nNgwD3gzESEGY/a02UzE3y50Zc5we+J/hki5xwVpRT3NOTR2HwVOdu9F
ZkMgUGMzkhYSOt/FfITALzry7VlmGkrB+OPBK32uotB55JZNHgs6FldQB2RM
Am7k9H1K75xxN69MiMKto1CC0vocaQFw6nqpWHfoVu31N+E9qAf6S46FdRkG
sp5eZ+0tUJlLA8DUFSvjp/q29kFtFzYV4tPtpPxsAIWeuLJJ6zOn2VTvd7Ss
pZblolbGMJskic963l5ZtVrIK6X/4UuErZZVE0kIawk2t0mj+NeEy/fiwOZN
1+bLtad4E5apIGrk7xe4OiTtnatSm+Kz26KAsqDJrfdN1uCSyhGikK7mhXQt
9qoGHAaClQNgbdKQKCxq6t11t85cNwPAF+wtOztWZ3L5U0eN8VMHprcoAti/
vETnRE49JZBFoYgIWbKDESODjQGMlpo5g8RyCUuslKB4lgQ7en+hIEwLyo5z
smG5/48C0cuootVYcYmJrnGpVsLGBOOTOGrCr8u/SZUMIAIZTqiw9iTIBUtc
SMByhux8FJ425YMqn/ITjWotoOFKNZgvqrdWEs2aWcANR7sZd2FKSEGYiGOI
cQLcW1Hzn7tG/pnaey3l7dYDHdDurKzWWIhS1jOyHoOKDw4uRzYg49amK0cH
2l3YjR9xQRn4ZS1gTR1Py6Rqu56dsWCG+RvGzJVv3Pt6NBLyGv9u3Iuf5G8k
Ob/CkcIJ2aRsPt7Y79nLdMmb//Y8q+PS61+r2WgbPw4bYCNRd9wQryUwn6jm
nn6EcztGj7HlwC+sePdUhDKer9SH129/znH5wblDw0lDBA7lXsnXEHT2urIH
pJsE3MChOnfIj450atDB25RfHTgXlyyJw/jBCloyRUrtgj5mSotaT3JDZTqy
HDXPMlQGTmFUYFy1mKZesZTcmf5QJHWtyRokY/cyIlTIxM3n/TCJFPSWJjlF
lZ2kdGcRMaTbu9kzrp8hNShLz3ODEcIWHwm+MoR9Q5Rwk5MJ825g7b56GBk2
R5VlruXHfDZmFBZG7z+WUxMa64Fts+z96prekDaB6Dtq318UciVAFmOn4aVo
KhST7brDz5t9wUyzDpH6UIk5RhM+dWC7bI/hIFIY0g2yvB4Xr3WxNXkv4GxW
WshDWE9SHheGdILnRjLGaN3rtYUST3aGmVsUUTjzjLfmF35dAZbEvJv9zqSP
wdQ/6JZOYMRI5/ciCNteChglglQe5QKgXSMVvYIlDqh+QNya8DV9HxXE36vs
R+MVVO8u5wRcbSC9lWo6GAm9Xc8o6NjjZUwU51V9P31iXd8NFxrS4ogFabUs
Nc4PL6izgqZfY0YT4lR9wAhKLVtuHcmX/oz5m1I+BYv9jrYSqzE51NywFgAC
uYuMq8cZRDZeK+O3BD7+qSiLDjCa5wb1UZNyQa2GmrueLjakfsZSspN9IAwJ
ZyyYROimEDkwAqEtQB7a6GfM0pm2FGSOfy4wU4rn896ZhSsG6uNoQshYB0KZ
WylNzKx4CGJ/zaUsUaeNZLRvcEIiIfd7pPLe6bgB9d9Ka1Nc29RSsIfgPFsG
lvAmmPcQp4jYwk4BSOqfhfjR7GErTOXFrySc3L127b2cEXmTilLwos3081tR
6DzHy0LkBjMD5cXVwZH1L8FEd8ax/rG8fdVxgWu8zxd3Wo8Y5AUQ6wGXe9GP
m/cwM1Q8uwUBGd58R7N1CeSHX87l5X3MORxIvig3tOIsFsi8H6+cEyuOrHvB
P5D8y+ajn8xRbrmPr6yHGsTPWm053KzxGPPjNN37BQXouHtMZWRrVBJp2oqX
SHJvMv52CXZyGMwhlFU5KGb8JBdsufF3hqGDK7Pj9hna1Df9IsibQnHU2yqo
wCyUdUzeoIbMA79YMqgnRFjWaOXpK16GxM2C8xumbS0xF+pbwjVGYB2hL/sQ
vNhpz37LJiIB8OtQFuM+BzJahtAmXBqQLrhE5UmHLD8U8y4ZiGgKQI7KU42B
hv8R87RdIymE5tqLCpGgTeH2vMk9yjxn+GcfiWReI7Pe9SPXX2VVNKAoKJOV
vxrfDr9i11X893NvxMlVEewTjFcfcI0wvv+vjqBYd6UUIdYB+26iElaxhDhX
Cdr5HYkATP9pm6AYFOQXS6MdGsHpI4u5hgMuFbqvckKebt87sbl0DOvE7KXw
swyLqNgNQWsdSYbB+lEiX1hfouVrtSQOcO86FwarDUwJdo34n3IBS2ZcEZtk
PMov1TvSCkydsuh8pp1dQXJbd28aXAt7KFYeL4S44+9reye9x4fHmV2F2N+i
tgNk0QJHe2uYrlX/HOCtjd/D0HgD2l9dA2qmEIISeJvOoOENkL9oS6OH4oyQ
Ps8x0TkPfp0XjI3KT9PQYns9WMnMoowDIb7mGb8nSFoIs/2215BNy0/fRz74
DLW5K/+NHPlviiQrfQDk2km9o2orXr8R7Za1Va1ktTXEXuLtpzeK5q6YmWXJ
PNMwq7UU4tzFroaZixoNEUSgXI1xiT/3pJSssA8nWpnAG1IANumseJLQ9f6r
HGAleNROmXF7mYnDh4gJJXwwruVEETlNe5+pFS0fgL3/A8Y/mrsTJjVvZ4Vc
AWXGKRqtuZcnxMkO5HrkwQgukgJ3GTdLyofoCxk5TakSWzsvwtbO45vYi512
cc2eczKXbnNZbG3jH2DTW10uHVPZe6FvE8R/xADwFbZhsIuU+QUYnP5wsp6Z
T4uPqgxEATfYAXCXdUGkF/8X+Wj7AhS34A9+KfaszJ40SCLxgdzekjlsFO65
8QMQOJzwO1AtGJmUXJad+RsjWi/BSDYw7wluXats7lrhPUrviuiX0AeODwHp
rZOu84QMLXo5aI2HiIfYJBPryMHS4hiriRzh8u6fzZnTJT31MP5ldIvYBR/w
qTlP25KxaISg2z9Y152xJFeZBGByxvjgKfHdBxSslI4R4i7aH8fG8175C7Hw
Q8m2IwrPlRTl3VhXOMFOafBDbxU6bsy5k9yoSslZIA67XYrkTfx53dD6lfnj
2jNIzszlIbGb/ua5QK0jxse8XP5Gdj9whCNoD6Fr1ht65wP7YsbbVG0SFP4R
4+9ZH1JLG/g3Dv+991G5LicTjNinUsJeJVKKBFWJb1H114VQ1itnuCMQz6hY
29Lmnj89Js3Fi8gKs6fbzIsWO+SVNDFaFt99BCTnF3d0JITbriD34MJlu/jD
o+whNOTodQJ86qCYhD4JI3OugND9qrOhconZoiQLr2FKts7kVHYcyud4Sa8S
QFDUpFaiA2fxhvq84XacH17XmpgnBIiqhTF8fxEkfgy34gej/APCP5vui4ZB
0c1fZ+dzM5DmVsWt2OCHhhQs5eXETOpFSErhuUCLuUB2vATR/IQKbMjgUhL9
XGOJ3ZfpOX22/WACDg1HtCUMCexFnesyRm2RQx6FrcF7NqOjddo8C1RDu6Ml
LzcXzS+/702hfTrsR5BEdVjfSsyH9J027lfs+qsM9zkSsmhiehYnzblP6a4+
e8sZtgrfm21DCC4s8Gma2qtwtmLZTIBV9q/QE2VUHX/GuL7kVNQ49KtthMzm
MlLZDex2j5Xd6hHoKfyqXm2Bbzzn3ytKBWFdHnmLshAG6NzC5TDXwHqlcIZN
945qrngZeRrH4uUX6gbVurseA9co1xZCUrkyuYLMsiPN4j8JKZS8PHa9UG/u
JSI4fjY/80UrAy02ScEhVvQGd11pqRDB40rsqm7jgRELhuzJ3vYMClzOMLjw
IQR6EiNWw3cqX5MspHKWl5Cwhqc47hevFu0kWgOzeV8hxSVi/M1hs5sqtHFs
91FssJQWiyPH8gImPlNEsgutJmjBg8LdxyCl7MhUciNoAyw37Y6CjpR5VdCV
8UZG7oAOExg8aaH0cIcR92x29VuB5JvlrS2Ay2wVeYz2MZ9B5u9aeGcNVo0T
HT2yqPGmGJWMjS71qy0eAr++Q5bmjb1GQAjivKovrNbDrB3tF5/8AMqINtmp
KdY2mKdzzetEowTvdzCIWQead4aZSDi52glGEkBSf6BkKVTsp3u3KtzrTSdL
rNQdLqZrNFJKuQHTCUcee9PqJVKs8tTOKOUqsqG/9V5YoL6JPSO8ZPVbl4fR
tGADHR2Ifj7tCzVzgC1LLMXl/QrPwHF2Vnr9fBLPwc2ZL1q2uNfv1UPZe/oy
hs8hdQ9ftGgxNo9vr/y18FhKTZzFPcmVtiWdLOZZxQWblFxk4tEty+Cb7SzD
YsYrnGgSUCBUDdDYqTJcHswdwdLMZcFVlLj/H0if03THy311O5qotesvb969
OYGIdDO8X4hHKHfgKFaWRzFsV9Ccgk4UtOu0Y6eD28eRzrgS0woZEEBaIPI0
dALH9Uaigp+g1MxZg3EaIPyrYPIwS+xPSRz3srpnGxKHtcmqHeqok44a/tdp
MgX3hSiCw0gLJ7hhhfht544Lx8hCQzW+l4HUVrWcDwXVURR07sdKTEC74BNl
p6b+fXeaeG6usSFwsw6YXoQF4wPywH9nZaCNli/H4aL5JhAE25huvbZLjcVN
19dO+lwpNZBnNHTmbhVp+vryAvmsMw26fuzpsAR4GO/a5avyljxTsFY6r1it
kvvEhE2057FJwupVhL3IwUz9xpkBD5bxqXnLKxJ6yTs7JrPdihaVMdUR9l63
0SIIQjT/QEBkn7b1ZSCpeHtvCYIU1mOxLA4E3LySxYTPdvWDKJcttYuG+But
IQSekYRHgSQNwd9dzIDkCTXw+6/AnwQ6aehpACm2viz+AA7JetyqT16vlC6V
vOiRTjgZWcABc00MRs/tTnmvvpPwnzfDRy6BmSkm1gOPhMnhhZLS9ILvo9Sz
tbdziEcsSqU33U8udTzTfjQ+QeKM5fqpzbieyVQKWvgMCnhpT42n4kghOvW3
xXzqXtPiFOtuwLvyFDSv2qV5btCoCdFAK8dGTNX1HOYbR3wywjzOIZ9LMUni
pKe4SaI49BpxXKzceBVpLj9c5yya+vRqtxcq9lM2IGPy1muklwn0uXN6EE1n
9d9QTBvvzkwFsJUmeqZ9b/RGGbYWtuuq6QTQAAu8wg7gsm2mb3xf/2/oTugt
D3GgCBKAuCXSt56Z+2+Deu3niUPoaHrqLo/ffG/YsnnUCmYs4MdtfizLnHGO
eO2QvPmr771DGhmuTjPIJ4P2YGbaDGmg/i53UY3EaVQ3BWhBMsU2itT11RKJ
fI35E+XtLkgjvhvWc92w9Zxx7PD+buADHlq0kn3ax9HJaxYLCYGWnVrloHMU
QUDD38cQRPoqf3M9773mvNp8G/udXizKIqAuk1CX5QqjsG58ZBFtHIp8VfeX
6FsfiTIIDg/jcAnvAnYP+mHw3CBYmPas+wWJ3AXKVSfbSJZ2AMz1atPvg2+G
TbTjNO9JuMbPgqOJwPQQpqYSO9s5p9cg/Jz90xsQZnyQ2/1ViKnzo/q82C3T
lHHYEJBypUs+OVvHRsrJ54vURa5cgxuuhY1QR4ypChqT40bA7h3lPOLdqoDS
ks44LmxUUHukrZun0XQ07yunrneQssBMngtv0ZttZKFBytNq9D7iSNTX7Grc
tDJqH7tkVE11IqGvmy4c093qbhT2qlENCDeIjxxGi68r5rBCrhnv2vzMcuug
IYfnxLEYyMCuOMqot0BqHp7F8v2EEdZ2jhWq05HLytVSxC34WBYE0CYOSSCw
rGoFrYsXsfH8cdePpYc7iOZBb+n5WwTMcfT4C58S34HoqKoYN8PSz1sleeUq
X0a5C9tgB2MmTW/QHmYhrd0lgfyx+iMJi0kfM3/UYvWUYOLo/f0qbmpSzSxv
MjIbSxAQslsfeX/0RuiXvqIRi/N9785gqm2EaJUktrxm5+3dtb1RZuYCKitC
8e5YUOxnmh8ttmO52Y+ND6js0s4hnH9AwrSHdnH3peaO7CujHyeoEZsHfnsC
uCD3zJ4BVFBVVC/27bCzkY2i5y8nRFlndNjSDqQN4GgqvURn8r42lHqQYhiw
wLxRrOlRZlbpKeMyAiI5h8cjoc09kvBwoQlzRkNldJFVPEF658+fRxdspvCh
YIvmMj/DxGsVL1AhMdmq86llpKnPprW+mhDrIQ6AHB7wUBfpAsBHc+GVs23a
8eFeACQDeeJtnwll/JU9KfDhWD1FLTIxeO0JnNIvvzhDHUgSiXDwdd08baJy
TkVJoZ99sHt5OISVlmOauYY22SekEh3WFVUoAo7M3BCxU1zOiswMpDlrkR+e
TGVb51AXwhv6aq106zp5tbHYniSwalA1ofR6wPlyjNwaX3ysM2Ld5wqG4Qwz
NVskPFeIRaaYMTU82kR1ce0tMSZkCOaMPylnn8HsqaI7ME/47zICES/8E0k4
qATHQtCStfZ9vszmCDm/yzUhAfeDvL+eZQP7zPXYbDSBscYih4Tg7JcL6oAR
zYH6fzkEYNMFGglveKkLL7F0VSBmLa2xhNogPxVOGyt63WLTszgLRntbeN5J
XE+OK2kqJ2zvSXo8dGSoPtd8ZfnaJfEbjUh8O7nkKyFTQQPDa0HSE8WlHi9a
XxqDfCsHygzlPD5FYxeoLlNGD0h1NXLw2uGKHjwxWo/Vrm96PuOz1hjd/Km9
WgQ8DgoB6HnkeseeNzZgMOZ7hLLGtmyCS76wbn5qmZrte7ob1tPiz/UcJIQL
yjYYptd4hBnAKrY7p85/oSXy/AqlkJuSESxnzA7tYwYFzb5Yhz1fNrF+n/ly
6JuaKGzhZEVTbyqLZC7y0Vi+qrQCyyhAGjLXow+kGInUcilvZeJmHyPWkBxv
AExtp6sFa1Lra/i4qrsYVgoOGahkc0zJQeoYSkVeAUTzm5w6q89fLm81pMwP
j3PpOcdeKGF3MppUIxzyysDPZa+YfMkp40wNOYBgfNMKh+qg7eQ15l3OnRpE
b6F4Xcq/2aZkQes8algsZ3k0S2KDLkDgIw7t/CVkp9gFG3YiZyDxn4WIeU0C
edmQmzAoDRLQ3vBlRTlzmOo47o5ypRLFnj3hL0c5W+V7QXHgD+3dIX5Cjrgv
rUTfPTB9BvM7zIDrAdCSIfAPjm3vLZhq2P0L95P1HNE5PuR7jZraH7VKdhEN
yb2TL8m4uFwgoBnsYU7MF8IpacPR05ZP2LCrquuUftv6u54bCyK+cNRe7RSM
nknEk+KmxKDuwqAzXXJNkPL9SoOVvbmW4+lBEYyr4t6wcnTNm0lDDor1XoCq
iZAUqR5ffY8HEOjFLoYsVUghLSPfVILyQS9SrEUKLwun7vfVJDcpzkYb5/jX
Pcyuvog5c9vB79sztwgFoMEeT/0o6bGL72jeXceZkpablUMZ9zRpA3S1a5Lh
EdD23/JyFsiXVRMPVNSzlT+TV17DTaPVy3Lu4opKmI/Czsu2rbvg4ejawjLW
WCcZFG/pmuhujAth4OV8DnQUJbw9Dudernh8cL1Z4WMdVo6CZGrwrdvNguRS
0pC//uWYZM+Yy3477LMsh5uFAlPoF5IGq5mjgmpyqeKTXw28aCRjTAUwkmMU
oGt1cyMwQxd3WQVSqOkpyV2XBj+Ig0nkk7Et5mtAqpgQObS3uEKXjihRPp7l
l965MGT2NooaXakcpT/LZ/SCUobuYtQLCcZmQ6potbA853AfbPGMQaDNp/nu
vw93j4SG8JPwxgVEhCLmdD1eZWTUpIfMahf3YBd1zO6NVVOc31U9WBkTljh1
+14mcvK9XmeC4eORUzSS/vBERIu8vvRiWhltBZCfNeJIc0NI1Y+nKCi7qJ1m
dB6QQcChbE9zK2puT114vGfCVBYWsv/moNuyoNPJfh72i7HoswbLFyT3++oQ
dgQH2iFjcrpq/VGqj0cfSjuqXnym7KQL6sB575sipXJx1s1vBlv9zOhm18ra
mH12Bbtn1Qlu1rchh8XmEhwWX12VMOJ5vtKJGspyabrlldNTFsh8AErLy7ii
SCRf0jM4IGREY9lNTSMhOsxdex5WmKZqeoTISAiqmKegi4x0zdbLs0x8Gd0w
/niZ3ksvPuYYlR9BEn+6rUcKrvl9PttPodvOkaxGNMkv214/GjRB4TtdOpBY
58tFIi6UV6R8MtE48TR/GVX3AG3XXEvTwD+0S3fB4dqQemfjtYLSldRQwNDL
OtDlNqV1VlqyMbSZuD3YJRoQkuN+kE8uu0ehU1lw+jmp+XmCSeH7/TcYFkAF
LBvlQAgQNzdk2gWMVIE0DlPVjpuCmr1nOdql95++FAdpkEfX95OAdEj9OWd/
gOBc7nqGWjjRfUBWqlPZqRw3+9ZqjqQxxmnGf28GrjEacAVYYRvl03ZUlyXz
X8AjtQnn7CXkZlZXIDyMU9eRcfkrJITqFStjU1jBMh5t+ecGT5Ih0CJ55cxw
ETKgsTPdQGaPrmEnQB/kgZD7MTXWNvPk9GIjNqYYAf5RiNE2uniHgb8gI0Lv
WEW/oKdM8Tm3djoNTpv6hd2BU0JFSqUOjANnwFXpfa7854Q6/Tk2tDqMt5v8
kY7PNPLiNmdCRPbZZFzSEKxCm1B4mXI7iFVHEdWsX/SSgyFMd8Kf1dJtPssJ
Pg60ZsQ6ZEhxEbEU0io1WVEG9KwXTMMI+I7BNdH9QAiIQLTaSbqO3P0QW0s9
diUNID7zM/yftMJwi47Cqa11Hd+zn8uGrkMc2VfcNwcKbDYx8EKFu10J9bTy
+iIyEWAk7LR5cYmrsAD7SjBFwgddPKZB0iDDjcqYQtm6L/XrypenCqMuCGsG
imjXp23c7mya7X4QRlCMZchgAHmvtdzEePk1sSURwAAAufVIIPDwFErHOmik
7Pm1DQW8PZU0simkPRTVF596tOaQJ5t+suhupJ5SjkbSFII2G13J0VU6K5EH
B59b8ppoQkxMpcUzxbTgS6jZJ65xlxiMi9/TTxfUNgPaubJS584raGUn971f
JMMNDT1eNNJ2CuxbBmEcZ1HHDIFjBHjWMt++rBMILdh/vmUc2+iOByewDAxc
VuPbP6efZfKA93zYfWVpQHdNQ8WPrrYGs8vzP9ZG5Yb+2UOXW9omtcvMcqi+
VsNwVE7MipTybh66Nc49/1LwklvdJvUp2GClthAFJcFBTvOjjKfW+waffYnk
TL7wAg+xdSrVEpaP2H8rgCwDuf5ZXShrVhAq+h4vgGDPkQVgwI/1sF2F97dm
MlZne5R1DDhKIx6WtjtYKauD72vT+nS6AqH6DtPr9Xu5rdxWkoMERUeDRXtA
+72/ZMocLO45pCq4TvtYMz23ekXK4q0MUVcAiYqNNCd1cKsby1b2aCGBULIl
+Zr9Ky3gM86pL/J4vaIg6XOTsck8mU5XyYF3+GcMxOkZ9SYesch2uu6qucm3
Cw20YymW+aEaypdluOrGqXKKUAsJmxteP+JsBUzaHmpcvg990TrKXK/gyidW
XZhyw4EDfR7ABTYZngjnoqkig/wOrG7WdSNMw4xrQOU/D7L8ZP7VlUSjPd0U
Fs0xTG5nG8a9zUiqUK9BI1d+y7uOPBIIXghRjkNoUSV3Oo42ZuivhRaodKAR
O3zAAhkjqvMehSq2bHWSNvo+rIjE8YpWSeYGnMs6FpvdWABD8RY1DM95J6B0
azIhyGAU9OzjfqmJOpPLwStcKNz0hngTY6Qzm2Q9qK8Thtju9hrQnyVYFFT1
pg16popFSTWcjZfu31tWczxGKO2LLgqz+0W/SoVscVUPi5DLIOSBiRppvDTe
8mjDzhMOPSi/kn5Uf3j6LB2d0avF0Y0oXi8gCHTvPSiHB5X2xiwCuT+hnaNT
12eaCsg6DzKhBVoTrqHAUWlW1k2N7WIwfaJdm9uMbqLnZKXLwmH2PNN5S/za
Amgh8hVwsjVjhkBv4kGL0jB/5D8OmGEGKoJFefec+wkVkr0YJWMDUaNcO5mB
C+mAkxjCRd5DixcuG4sHFXzAo8GIWw0B7XdEzcbHVu/cNZJdRWbsQw/B1vda
SG3HOba08s4h+XyRrtea0o0AEldLpdM6FD+EtJNmMFsG+b8tbqeyZtxzmdRd
qxtiJEMH1H5p0hpvhQbl3flqmFbxbw7bdYFcrFih1Xol4EzyXLPGir4QH7r9
PkFbl9kdlLRDiv7gbP36QUtqhtoQO+41Nm1Fan155zeJfYWhayyFkeyXwAix
o5QzvUfrOk8Z5HVmvERQfOMolHY/6Sg+ByPBSIsfz4YxaqE+O2wLt/xFPPpe
TGILdB9o9KyR4Jow8ASKbJPN+INeeXAkQg0NEYLjA11T9GdEOd/iuIW/8oc7
KgZAGi8CKF7KNRmvmuqCsybRX1NS8VvaaA48vHTpt8fVLQzAmgw1pMzhk+PR
yNl7xu+PRZiPk1o60nVbLuGPzQ4z/3Yv2JrhATpvT9Ho5JklUg0fCX6Grt8m
sC78Myv2BrJvYy1o1LKV+VwS9N4KXPEbXXz+iJMcrw3oR8N3keSw5WZuoWFR
JEO7bu3yye0MQfUqkF7xUmyhdFrUNNbXH3m7SiNcWGXvuacdhX4IenxSpdzE
UcVG1RWT//HwxIsBPib1zhhBbFFrM2L/vcXVjHin9O0p0ZNZ9BRjqXi8z0i6
6oLJMQrjvHv2E1timWMUxlVER7R+QAiJHo9dOtHvq2CYRlC1IqOQWfvKh/W4
S1wbl/YVYFb12rkyghmG12jR18SUK9S6isLgNaBDhY3yXQchii/B6W4Lbhko
QDEES6wCmu82QJHQDLtiq68t7d2cB5tKvUAmMy6RNuBV8m0XbP3sMx0PeMAc
lWr/SxxZin1xGjuSvYldwfKcStmG1qARn0fu+xtXNq+pNq2j9U955pxpp8LR
GYGkpu/DQhb24arjTSc5ZD/PWpMqSBK9LSpyFWTufkwVdTKOIwl+O2UuP3BP
qvDiHXCnFNxlLbTIM6wkrsEMAeq5njraeAE2EeQmYTDvIWU+OoCSsyeEm05m
fNPm/PznwoNDkKp6PePwjkYGsEFMUaU5PZ8M+dv9j6/rCjF7K/06tTB8HpMP
ojuzndVdmESzvf/D07L86U1r0ozRBlG876CH436XJuDG6lUhLJAcQWFh0IYf
YEcmOjU8uSB3ohKnyVIHYuy4Q3dIBEI8FD3lLE4b15HdbDQUrgVJQP08IzCO
yJzgs7XGhtxV4XmRlPUhZYlxa4gZrVU5eDme6pNC4qdzqwtJQ1byXHgFFQzA
TReVbqfBbt3T7Q72ypvc3h5U6Iz+SiwQXQzLT9Z+w0Jd36ZpcYqVw5tkthTK
j1c4IIKYOBVA+t8M0D++tVfaXp0tpPAJ9M2pA/o2OD9VtX/T4wwgl/oBlcFa
QbvH3hMj1sMuJd1kuHekOzYaykY+kwzqVgVAV60Fbb8opa6uLZUfiLrf4w/d
WrPAcaMbI9lO4TToOZvxwNGN5HDIuZXjiZMST6sH3kcDwHzF5lcSJvML7SqA
YEzpC9T4zz2K/KBnhh6VLubC9WLv5NNl0bqBMzTrL0JMOmW7+iymYxQLeRU4
cQNnXI8wIDqR6zQSTPwz8yIkFNLqARRyQYBIXJYlsghBHTsWk676HIuyM/PI
r6mszCI/mTHFj6Xclnz6wx0rWe6tIRvksqEngXBv/DsHJNUwDulS1VD/5sTN
W4iJnO/HWfEzN+NBDSZ+Y0dQ9OTwlZh6Q8kB5U1nE6uwWm0ImAV7WJ6QlqWV
BFs5gQsO20ELE19jmD/tcTa+DnZruSFhFu792HvHCrOnaIhNRgaltdbnrnuM
ZVSvLPn0cnIKbxeVX4ftVWlWbGZsez9YB1Nac3pmXEPYaq1HnruF9w1i2fOs
6sj5KejFsg+YdblzlVZBVunvOSgsDq2RYEv5ahzNYVukf4tUyqFCU2BI0C9A
6TS6OGNIPs2E70DEGRsQvGd0zlSWNc4e0y59EHN/P4t6YXFK3SE3xnnz0fxe
Mcg3+OAUNQz3rnvvRxXHgBVBublHQCXtU8Qb3pc8V/J6b1PC5hh4/d459gSw
GIzSsPsAv5VqzEyaRoBsu3Y4O3UgGNeOKGO6stywLZ92SLZbwaO/QCLi9hUz
3kq8UySALq/XAnkgz7cD5JcJ/1Urog9uEONm6YQNgIbPDjzaued2rM+5LYPr
Jl86QytVVx9oGipd4UQoKvlZ+YQ6U+SgRo0ijrEXo0PY8i8bsagVfy9LRSiy
IbB0jb22jYlU7j844uAOyiZk711k6VPu40nB9eoaAwqYXh2e4sWm9oNXAxLq
ragjHIAcS7uYXRd3ISbDNpC0yyu8BDLxvbU9d/eTKwoXkD/6HMfPOeEu2kxC
9zMTEaI2HaeTV1RJ5FRiThePhTTS7nIlawbVbbFw/OUpoPjVGg/2nUjyZO5f
f+4tZANu8zA0tJWPx1Sm5+JZSPHVjG1d+EBKmUWNncOOhuEXP+SC4xqivYsR
RJ+PACjdDnOCw+Xrd1qmT2a/XFBR8rSdXeHqM+ZzLOFQYm37nJSN04a+h+AQ
AucGXChiy56icgOofotuUo+a/zUo7SbxC+Kwc6IenjA4ytI+hCOymw6pMrzI
YL5rWaXb3IxwWmacUTZC6iavltZEwvmFWjMzs03JD+zumAFgoigqGJb5W/w7
vqplEV5HYZkxCpuroxbGqOWxffMlnDfy2/Pq8gIpfnyDWJYuw71Dyt7S7sDF
LNXRn/tty+0svc8ISU7sCM54Pn+ivwq5WE6F4B7Ra0XHAMj/OJ74gNL6Lfji
w7aBiK5FhPdmt5gu2sFCJJgyh1GvMSCQzdue3TjHJ0WlMgA5Qu8+prXLwuTe
3JHyEUbnfsuzKsgSfyebeU2kDFVITni3QTfEWkokLzqg0yR4jV5xXSgb994D
74I+R4yTT11tfBbWWqykDUoQePzeCbduI+DFkFUE19cRXFppiCff15KNwZVp
sTWcR3zeRYJd7FIkji8pDpPMz/N6JYJta4X/DV9OflV8LK6ew9O1wvpOIV+F
TYswEhZpgYEekMZ0aU9PVSt3aJeO8vyIPRmfwY7kvfAKJcPTaYev+fzT7qQw
XwwEmDkBUvcEHCQIwD24cmRIIolykuCb7y0j+83nz25/18X2AEWOAJPhaKwT
xJ6L+6EAKMk6VIF3mnXeJ8xP0P68TB/bPSKvVPvcnadhWlE0ELIygcZIwfLS
tRfPS0tSR2GFSEO+Mu60dj34nbU3ZVrqceabCH8Q3Mef+IAmGcxAfzkrUPh4
xog4G1L1QF/ZH/ssRN95rvbtkSl1TCiVAjeTBoqdf2nKnh5+QnNtDDv4EkTj
DaC/vIndRHInHx2uQhIukIk2z88a5e1XePrvnpGuUsJVdxpwwiLO2bXoQjB2
/IuWpvgs5vzGxILqYO37He11O+mhxT8gnb6ZWweS3r+ko/eqr7MpHEuBosQX
xPQRicPqykYBTAXyI4dZS2iS376zvlcG2W5yzc9ln3Is5flfsMUeQ1+89X8M
MPhpduepNT7ewUIkW0Zjw/ZjqVgrC0BHQaFh5YpvcgT6HQu3PdCn6rbTEuM1
Yljcn4WSfwLIWW2omTs/BNRSAYkLzeB49cNKwey2qYD9kceWvLD5ejr2xLIs
JDDy8anXlO8Y4vpT7yF9q5GvZIsPooXchSzsKFYLZpsexvmHdzIPTl5Vb4Qo
EIjtihbCxxfgGayLcqSTKN4IUfdKUv6tqp4LfmEtYb5vlyQUkDNRPHBU297K
0RTce7MOGenweq0L5z/MEbDbvynQgLEr9HNt8sRFT4uBJSppXty57zbAB2uz
NPHNKJqG451xR8IzO7XYKEoNH0fUtL8B4cqGn8PELiiNe5VQsEdJn41ahGLz
WqBlBpFAvL8g+P/Oxwhyx0+SSLuDjycXmKM420B0oFSSLOj6btdd/CC2Mi4V
FiTlm25G72jt7RHgga0XzAjp1PcKu8FNR+ouFIuyySeg3UDz9v5Rr49xyIJt
x8IlYkyYFtJKDXo8Ve2jDvjhCEK0j4C4cp8wKoDJMO+UMoOXbMe9SIqpvqKT
lPQLVkK3TiLbPaEf8RnYoP1JKyQt1wv+K1htuB8aXdnbG1VhlYfPYmQnbuit
XUY4m8Rw1GuZgt4FJLaoULturkuR9WCz/AA6YeA6AAm7dIEz9HV3LNcwmASK
xoIZKG68I6EN4SgRyxbD9J1LaBMbZsq6HhddoziZw84ZmcL8ymbJFrXwTT25
/bfn21s41p5CZxyJty7d17hps0Do2nKVARVPWClXYGtPo4npXwRdnHgUIvqQ
sYcZeq6o1pdcfdinIY7NpYTNfgNDsotC2DSMtnozf2tMQ8V8q2YA+qH5TyH+
hR8g1RKWyWNTipF+ANW6aJUTzM0eIn55Z/g7si1BDYMjhuQgwF+XbW6IgpN4
VsQzXzwINZHpHWATnPkzdSdGuyg5b28oz8lEcThFtzbSox6GLi0usQ0pLBfa
d4r0W7mKmQ01LZO/ENoM5kRhV6egIFpouum+TPXpqmVOPDKc/0Jvl+B0nj2Q
uQhkipW7XgelRHOHengjyV6SEb5bSDo9dpnGHSFUmJhAazlxKLpgPlYrD34m
ZSCEPXtWoBdJQ5ogW3CxG8nWb6DluzjppgNWAAC6YPvbX8FgG/CgFLqF5inO
R2kSvOwL3o6bt0bofOO5vTkJbxv9fr4++ISkSFdF78TVkjrY1B1MuUwFFIF2
PV2nZlRNNQSkq4+XqMpwB4qCmvBpZ0sGn3swRlJWy1lfFIC+kOTkDb3zsB1N
NHtysXgxlPibmwrdvSWvPv/8E/F1Y7cqPKL2XHy2FggMhuzO6AvmZuiJ0YOy
ES6Zqvh9wxkVd3TqOD9Y1EYh8RCcYr9OoqOzeVereTcZ4vXXKnd0xWYLmnUw
d2+8oYSp+kpORB2nRPxrakEE8S0IR/uZIe6swjFKRIf8a4zALLHJ66MIqCVK
NgMRBaaojmNo1GPkqB4xVYDvP6ERNASR5jIc+AC9H6HaEGNXxPkitMgomBoT
Q/rQsKe/rmwZJuyBaaPvkM+67tlS0fEp1PmNZbwSOOGlBJ7Nvvsx+1I7UZJI
pMyKGi6TZHM5Y7WCMcE0hAUUGDwM+eRoInSMqx87FKzx2evCNSS54z9fSXp3
GC3cW1l1dukeV2V3b2dmrLbaAouleM8pbmmSb7dFKRXhCajvtTJNMl9xYKr0
Tr/ej4VQxjsEzGUvhTRKrQ4ahuWg6+Qw73fQtZsWca8gzPcd0wBOxIJNZSow
X7X3DZeTLhOAJfbWTDKzwmesH/ogY2HCpBoTKWTaGOgXM/t7iM2IUaTk64FR
Oj0X5JgbowNNOuZE43uOvILsCBTo2OPvL8juXRsSDIebgEP/nFj+361n9OKx
vSr3eJjH6b1ZqBnLufUaH0iYxv/eJMmfJPAMfopQxYp7ZwASu74ML9Y5MGiA
u8H/bVvBNW52/MORGlRMz4axAqESWzI6UJ+aKb0InWLP4vcuGWLHG2wzrYF7
8+XAawVxqRCK/gqBICLTBPFZaDKOwPQ4HNun5DrcfhlIWCiCzZCF0F9xVE5n
nUrIOvdseOWKi9UIp6quEXB5PrbchvSLdlS09fPUHSNw67YbiSnj/FgdEYH3
cEbAHTWPMabMjVHs6LLFMe6q1dV8v2eBcStpZEAoXbWKntqZbUt0T2TvQ4Wg
la9a1TDnA5VgZed5ryBULc5fgMpSf6JojJ1nPl3zsVQiR0f1fObvMEO3p4Z/
jhWDmN4U+iS5bNUyRMm7dD5srz5a513uUcr/bxQFMk5CYnLNzOsNw3hXQ9x+
Z9r2NM6+EVrZDYJpQWBTd9GjxSCEze/dUfG99dvM4skynj51FAcCa5yUez7P
7wMv3WNaY99e2aGjI7Ga++EfRd2WKcry3AYO6aYnDLPPW73wwa/JAyTEyVo6
XoWQvMJqPAAUcHC86/6u9Du+gJz231aJNdIt9i3q61OOTcsOnSmBNmCZyWzK
FGbIbJpUQ3bhCF8exU5WBa7CEZa3zAfLVUfPEFdJ4p/GdC2/wlyKaaZHW7Iy
+a5I+7Af9cpRXmtnobggldHVFaOsFv5S7inSuj7KkTL1rxMpbdiRKPHwHTmv
LYYql0DhpOzlrD6dJlNomnXWlDGR4BzTLT9Eu/tvaAuRg3bvLM0tySBQlLel
6FNFOA/XHh1mWjHwsEpP6svWySjOIKent55M2cIy6A840Kn1ey2PU9Q8LDfE
ZIW8Ma9d4SURmxdx3105VWsDwmE1RL3gKNb72SDdN1a9q658a7d0MtW6+X1R
a5aBJCOeMZrToisF72I8ZGi6atOtGupw7XWAP270DeT1egeEjpC5ZnQ4ncdn
JQ/3JzOTs18tOXQbTiWk5ZyeY87TNAVIAZhrQw6C6xIY54A42LyXBx4g1cG8
KMwZBmvsLcv/TwJWtH5IA4KolzPsKioO9MG8VbT20bW8t9tCZQ0A7T3oPqkC
OjvJFDNuiz3tPVJR97jYDPMQsdLf7AZWQIBHmUlF8OpXA2gJWtEyoT4j0iss
xqxZMON/YWW8aAMw0I7ZLpfx+IBFHXSoUL47sZ3eTfHquOMNBEhC3/MiLVpW
tUF3tc9ZpRsPKc5f+Oh1bJtoGezNRk5IBC+9tlM7paXaEZ8VJYOvF9LtvV55
+zArxggFvCjsn/qYP+S3CDoakrwIv6ZH4ZTYDT+JxlrS1doo3vqT4toJJv4k
De0LFvRnKuoVdJPB6MBZ1ARM17ZXy6JjNvempSyIiCOTcV/Frixh3YyuLKj1
TbfE0PDDfF8iHzAbYPoFT1vJFr9jphRqA1NqEyJdXc7fEcJ3qnxFraQeHyJ0
RkCI+GnM0He2uh/8MbR/BpYp29yUaDKyIDeVeyxlk2zi0g4rXNaKb3+Djjfc
BMj+UYlJ5L+NJ05tktcrHm+y1uMVWTfOTxknS1/0PIUiQoxYed3opR2VwnZq
sLysBgRyosQaM/yQXNzxL2RRcfdVIEL2wp3Dn3kvq8MLMG5ihFKt9M3Dp/4z
2oL0x0ZD4htWfJCfIAiq83RhkIM93yGdS6lh8x3QyOF+tOLn41m5ZTr3b13f
f9tMHbJ6EW4CagOHJJGiahw+XB54jnCwsBda2H/HkeAFxRNb2P+wzf44zxah
S2pkDH2mAsKwYNKOdr68y4UYoQkfoFWbhBHCatT21RnyjbB/+k58UfQK5pvZ
RlP0VeG353BMpkP78Nl4vJ4HKaRGwdCR9lBoxw19mT57hrK4fNHHSdIzOzXU
arssag4jIyWJ9Mr5HTKGCEEJz9S7vtpFvF4Nh6YHsJaP6+qBtw85htzaCewb
4UA0xNGdwjAdfu3CYqs9dmWz0N+MYk3DFvBp8LmkbuRFzhn6KMe7+QztCbZU
paOeicIOhJzjMJxZ0EPYV6clk3jAXCAGf5X3iSl2dMid55Sph/AjnLShXwbb
W7BbLWll9kcWGRRhwrapuzE+rRnGOdeTtQDXnJrkiU1xy2j17Shrbwpu+bH5
tg1r2NjV3QR8IR7LVX/qRhSYGWduElg1bBTmOj07idaBfR1ZXdEK85YOUcTP
l7162yXYTytbn9FbQJQ4GCecwKjY2RluSuj9RJyflQGIZy8scEkfesX7vZq0
yncCfqKYzpWoZRwCcpqc9WN+2I+EuqVijgyG+2UJYsKfWLD9/cKbhzXWvB1Y
+OhSWznW2M/7eK2eSBc36Kt8nP4bk9hNScSjG6B/RwmOD0gjZ+XPwkVkt/TJ
Xcjn1sEom5ad0Xe5snEEP+Ujqb791yUdTWIngzs+2TutfY7kaJ3gOimwHrTx
Hiyv1VTizvn12aPpU7b2SlhXg7sl/12s4BtxcbaKg4Ph5fbbf5uS9/zE4wn1
hUrr8Jtv7rDPtW2r87fAs8pP0uVPfOtnt5eXq2uEQHypOAN5m/Mo6935bGN2
30c1RVZUCzNKmF1ZtxpqEFePawIUTIc32kgmB5Zz5v9Jg1J+0RXbYCqLrGmm
O7rOES94JMQSXqzdoK5h5pl/CATSL8G72FUbLj4wNOc7khFLsHufNqitAV7d
+7fB5tkEgUN9ChfyFSB5jHYYXak1cfh0+2EHHFqHC+BbBKeoYF+az+8Uz8YM
uVIHxsBSr7rAaZGTN3NzjKH1khJAfYIN7QTadUzLqnhNgXHzcR/5BjU1CPj1
oRqZIRM1xtYpz5L+n4OJU+au7JcHnbGyAyFg+hSQjB7CEQ+dBUd0hUYbFuHh
cdUHFZBHEkWWMQ3Xg58cecC7TmMN+n6zSDKPPJmSi/rnEEqpDvNuhHz/RZB8
ckeEu0g0/RtaTy8RcJO6vZwpnRjvIxLGN354UMpOgpplIZu+j9VEK9Q9K+HU
zVyR0Botz9lcQTZ8eUA0bnUfywOecmZixZ2jmdPtUPRwX3eZXIuEEulg+aRb
crIr+1KePy4n61hMQqjsdHOjS2b6LbfhpNfLq0lY3LjIx3BW+woMNLwSp2d9
or+eHfb8717qm9SsHA/b6Vu13kXieYXslrkymLwEvGY/JGGp98EuVXKwpEU5
pbSZfm6eg8O9N+MbCLeVMnPhXVFsh2uOaDbB2xD6a8ZMlQ+LdwvMyryGAds2
l4MRH/s/B3FqHDQaEWGPHy0mJPU9IQeU1ySAB5xs3Bh6zLABcHhl7vMwDK7G
ANrIhgd02XEPsaXXBqd4ElxoyihKVBdspoMFRsI+sHIMYi2t/2Yb9oCgtqSq
/3W9feX33rOV7sNa/bF3H2X/RxLt8kV+XaGY6i42/BQqw0BF3aQ/JWfBdxy/
kJDQMeIKTkC+L6nkR5VHGkKAQq646SWWqfTBtWhKK1vWHAP6+lQbefM8u4u2
1+pBJVyFZXNZI9aQG4C991bWr2fozF1zcnxFYwsBPVSQXNNfOAvY58kQIIIu
1S+te/vvdl8T1mpFgJoDjgHXkjUT4bfbxM/M4CvYtGmlsld4G2PeGCR5THOb
yjPVWsvMPIODqgy23iMA3KBCI6WGo1yYR1KPdwO7trrZg5vjD+pnO3fQww5a
5AMLcHiI76aKC7INyN54QtKUr41ZTTAwi/b/DodA8u5qnWBY5frK1JiMpxAR
ouR3lC2THxMX3asvqJpeotgHiB/i24J0iMigrJtVB+lLk4MPo6U4EvcIXGOy
Vwa1CGgnYIohyauYRP2gMM/8vF+bEmwutY0aFHlWX3Gnz4B18fMtJbqSs5a8
dUdEkstgYvBoHlS/kkAavOVRNF/00IBmUzWHnwsHNDjN/WgYYdt6AnIwByKD
Glzp+qLATEXuNuK5Y2ylW/nrEu/4hkGB9kLeE9am38lUvv7Sc3bLKRTD6WjC
spwJhVevqgogvQLpfLf3Mzb+OGs+/xfEsH89yNiQcEO1hcyMpmlkU/ita2iE
SCFfMjC8Eryd4yfO4JI9ylQPjPDsn+QIIEEJLNlhHbcakDl2W+WvupfcFpiN
fcOAoMVmzAN2cZ9uQEUU7vqdB4CC4RFiJz3K/PVVQnjE8gapsg1a/hnrVNAa
okC0TZWr/o/sEAamVenbix/v0tsMPUE9ne6MWD2IxjSh5na89mmicDoeIz3R
LCIHE1ntbNBJgp3MXPM/9badWjJODJYyoVsHJTu1YAr8CU4Oew4OtOFRUcdt
ilQFdXaUkv0kf7IEGWF1vbv/mYwLGFfMPoqLzAKDY+39Qjn21ydh67Bz5pUu
lxo5wRIbzEbYiVsxmWRgzyk5/dfOHXFXNnJFj2+6PauM2XW0yhlS3qsa8KkG
2LV9Gcxe3DVUqxReLd7teG6m4zfEvlbD5M3CTIZVxd7LVlS+2Ijju9ghhmd2
N2JeU2j22zJqueEU0uVU5udQchAehBwbTPg9XesopEkfpiE+2CXYEgNRCn0V
+6RGJcIzsSFoqVEstT1ye/qu3ISj8fxN5N1URkwKcmJOzYki4ztwyjmiKZ9q
VwURuXldhyiFlSnnryA3M/BpdvmbKjtQJjN9iCVLiAbUGqvI2XaTtFoTnsa+
VqpJHaQVmIKvpdyLvfzxF1xhEUvRJxoP0WSI6ZPUXf1izooL4LjD8PIXo01t
3Kh51Xq68WCG0xJ0LRXsBvBxoAejjQXZSQ2W8Em3RgkXUVyyKfXNLTq1QdPg
qp3Yi6dRSSkO2uAZHCxeGzzIOM5kL3xRZOgOWhVLc1HHyNf+ptDBkafmU+6g
Nos8d2j7FQgckGOfeSYrKL/ehBrtNfgS5UDRKJkfu2BWGlNO4OTcpvQmeeVc
cLW/LsCPim27/JNaryucEzxx7e+2hI0tAVaP/6UL6yP3OFLTI1dWaKZjZomG
wXQJkllhga37u47+OWrvFCRMRXIKaBMRjj6eF682+jC9tquodNXmaAx8ZbND
T2CXsVFTXLzPICggek0rtLzH6XHgsxA9jXpi6cLRq13bnyzPdFyDCWRPA1sq
xpnUWcNRWFH25Q3JWiJiz/zNi9UJ1o8XtMcBk0P6sPD0FHRKtqaDeTU3mSY5
avAJ07bnmJclbEvwR7GebE2z5NtqQnhI+7QmWuZzvfbscPtPW/PVuzuRUP76
W1AMWsqxJnHMWclV9tBtmj0mktLf9g9kD9chnniGnE8KSWDMgtECE/DasrHM
pkpcSN0DyfIFPIwINu/3V5GUuckq/RT9Dn5NMdzb+LEuUCEd0uC4ePdI4F7j
ojrpKVHWBZuZU2+uBmh7GDxz+BFe2GQKErMR38qhA6xE6vLfinTrS9KfnO0H
9I4S5e0adA8TkILy3GYzFlRxruEuz88WBrN1GH8H1Dd/tRLZLZ3WQT4E9jUU
0kOncuAEZrWAG4/7HEKoC77pTYFPbq328PgPzusQebsE3zoELwkJlwENijGr
ti0JDUs0WtLeN3z4u3SqNmlJOwE5G3r/yv0lbn3SmKQ9KOvtugYVkse6PalI
RgnTNNX/semNWR9eumUGakQL+pN4uhRAuUvYE0WAo47EyTKD4q3BedQl2x3N
mz+BsIpWofvf+vc+L4TShFYm368wkUyubBoUaPx4mu2/uwOzSAE/dOVN1sTV
D6ZdiAD4B+1go9IksD0228J7xzKGqhnjP/aaTaxIlyMnxu3XJEBq/iY3mpjB
PxSstsKuQZSwUgoSoyEgkMiUIBt6wUKbRto4c0Ge70l1Hi+srV/mTu8R/30E
vIzcVT+TY/HRepXg/Lsqh5G3PkgWa4LM6hGDdWEVe0P93mZhu5P4YyvSZn1F
hIp5XGuCrFtoqCUmwlOFlakEYtb36mjRzrr/ygc8k29ndoMW248YwQZRihe5
nTwFu6+8kCgO1Jr0Q60fZd/VPwCK0u8L1zCVQCcH5I8dt+wImO0OhT+jbM35
2QJrzPHtz0b3RGsUspGWQmIX62qTXxiMSLl9ayeu4rGPyFzWCLauzxCxakhz
PpnAqXzwc+AcXTut+GJbf4JXI8MAhhhV44WfpEvvz5p3mY5WmguwpUvjZI+V
+q4ar8W+myjwpMCnzsMyBjPeHVqb6EdyAL+9xPPI/RJBfzL+KNxTCpgGvB6u
i9K1jS697mRb3mt28+BP3/MzHd5kdIg3cn4NicmhW5dZzrnO4rAeCpU+51qV
W+MZ9igHDrSaJ0qtuUGe6QnCYeV/2JCD8oz5y6+cmIQL1E+6orVFy8ZR7GO9
Ktx6V6aWB0jTBdCV/8xanwIXyPXKhWvdajoVCHq0ErtDhS8m2SffycbU/a12
1kKlTiJWyrSsOzAwLh9L+YN7TFN0dDy74TMkJoQxsS7zj+NKucEnjBCg+Orv
ASzV9eQ9CZFZ3pbcVh2PIhrmQ7SPsmumJeWjXYFrPAQ13JThFiaJmYIUSU4q
62V4fK/thOkJsIqZs5tmARmXUDrJurfY196RmNLcwTX8DYMqp4VhvuazDFe+
FNeuYtXCqDF+5pdMabBjUZx7bZb0lKsvOiK/unudkgf9v2WKfQwXCTX9yA21
y6NIe3SHB/8vciNZiD3vuhy0I09WUmqYcOil+yft5NJrKNVtSZJtDG2QvjaY
PkYIuR6i6ECyVnp8QjMafEGnlZLzKH+GkBLvNNfQ6Q0VPkbXSn6XClW8PUf9
vnr7W/nR/RneuuGgHLdJrpmgVDH5KmH/iQxot3lEUTEAUCrvVrv7uLF8qRxh
dGKR7qitDvmmUMC7eRsqy4aUPGL+4htlbhb8f6s4hGekSR1ypIftWW/Y8v8S
0T49VADI2eF59mxc3giJEuBlEfo0hcTJoD6955tHXSmJKuviTXI32y+EYajI
cM2Zili1uQAFb57T5Yzp3wTd3G1TsveSh6oit2w+OnQMv+RUO5T2HW+HRT3G
fhCx1fcIOND3xtXnCh+We6yLvjvA7RV7rwInicO0Fyo/OOtf/Y+TiDVcGrXx
P1ADHbBbGQvODlP9A0zZOs7DBL/aW9z0rktAzOp6oOTMJHZtWiqkp6FVE7ck
OFemHZvjfZ5oBabJ8Jxs1Jdy3DEWztZ8cQHdzhA+0SagBfKJSnBjZ2TeqC04
8+LtXeMkIDS8iu206Sp15lJ0qKjgKO/ANOvUnbgjScAs192wdu9fB/2hgbdE
2UHPHEDPl++Kgq9pzy4b+fs7DnIv1sXN4uDKj9SulzZWwEjLrFoEmaIqS4Ok
/QbkMQqBFg0KB4xbDjjq6IycL0BCglq6Si5sVn6DlArHTfqQ2i2ZSZVW1FbK
3nVNgjmMyET74iD7NeZco4kLLOPE9Vo6P073S7lZosk37pN7sZJlPNgwIUxC
m5xupA/Q2+XDv32jjwwe7TdKxQbEKRFHH2PkKXaokYsb/8kcDzwwBGaAXAoh
nbqvHKTm12odpd72QiRFOT5ZmdrYAtC2WQPtc36go1ZFTQ0eTC5skflj2vVR
R6xWqDkXq6WsPoOB5YcBxGT5ZUW3Vxg1twDvnJxBfgnSsxSinauwLWC4OonN
Oz5mn792hzAseC43rjdeXtWGPjrFT+GmEwh9kcalAz5Avzmz1AhyXbAlvsZq
1DkBN6o5vvmWEZcGQmXIEVBREglxNARWvechkgz5JCBneTZl7odTws5hIK0I
qa4p8Fda2uy7Ce2mvlZ5xfDaW9cFVBJ3y+IILHm1oxe087XJOtH0lLxeUWk6
JONaaQ7D9lyzORONZUNSLn0IWVX8naEncFvrJ19IqSkOBVJ3b5creS7Gn5d9
v0HiO1tj4k49n53fViB9KT7YeHucEd/p21S7tWBheRec+SkP9VSDGU3tYui1
FTxqCELz/t8eMTi40z+lhsX/rtI6JMTxwe166gVMjVExOEwZKRgFsJ30tBC6
lwsOLXrQfXAnDg4lqe/dBBvh/Hdd3aB0qKAcP6f89zOB4HCf2J3rJiJIMa/9
2OdVd8fwLJ3kiIDmr6rrapvjeSc5t3X7JWVVrow88thBJ9yHgwkNORd+8DE6
CV7F8gO35M0lFXWCDZ+vIl1MBb2BrA+Wles2fkE8wBaYXx7nEYV3S7TOHXu3
OSfLc4gHnkJaAOyI7oItW2paLZa7rnli0k0uuxXB1J7lev8hnkUG21YaVm1j
sQDOTuEVX6XvkYWLjMZCSV2gbmYU9qmkGP8sqZLdE6mMvq+dvL9tDolf14hy
RAwkL/0/uie7nU9fajNUDEAoeH2/2E9XJzEzoMkoDNi8fDedcDzb4/s3pj/a
xsrN0k5105K8kJJmgxxn6/ilqhqR252reytR4AM6h8f4mbPn5xGbk03+L3vN
lJ4xkhM3qmyvFcUrYNoi0JJouaomFpHzV3d/VrilOptm23vTPQi5aLhnHZrC
+2aE9OE5ClVm3ZVA2KKSxjQyKqk9jjkBMHc+75jRquKMtDznKIVYArvSnK1H
xPFwT3KwgL3FXlSPM8t0/gqY2Hi+AOaeYjK7SsHSZbdIsPeZkgTFvA5HJV4k
Ocvbp2DyDEZKgcmIqIsRsM4HqLwuqgmNRTKp44Z2dD76daXPVuwp8xxQJRpH
iW6Z/l+xkEEL17MsQCD2V0mQFOiBWlPp+5fPzNW3iyr5DoCjiX0u/qU4vHwN
oCYD4smdmbOG+j4wZPV0MjNQ9/SCD6Nhupa/Gbgwz/SRxVyIJu/BCPsFAAbn
wKNhrRyV3yhZDrWiqzilRWpnrYp7gW7oVLevF+3xDfinEN1tEwUMTfTnDNxD
ybLAU6VVA97K/zYBhppOkHr/b8kT689X0iwVOXykSTehv5x4oclhKyD+iwLC
kfOtI9Es8qi6fOoaJV1QY/AiH4r+91XibZNBlgCk3ca5Gw0hhvSoHSpwXME/
N445dzsdUs+UX7TKQKlPCseD8+bzC/qyji3t2wjl2zgv5zn3yVOAjekjwCZ/
kD08GRMJdcRyEVvEmqcvym75fW33GffT0QUSullTxW2HqdRwFmQbK+j1+ZBQ
oe3VPP3WjM415Q/3J2MJGiHhQ0uaADCSBxrE7ZwpEDhFGd8ckC3tN1RcbMbU
U5W/VbAz9sAZfqoPs8WjwDVqxhHdwsF/Cga9RoXkZwxbQ+HXEJGNexX7F8/f
YqkQuIlvd1MdiFdKT1kdsPqx4qLH9Q0KYHmCTdlRwPHqaUUhYZRwqG9qIhOu
oeK/vRJ97dwe8l5v7rL35c4zhnsnNa6XLZhGva8484ETqW3SKa+LWXdgLifl
vQjL2MLovg7lNPS1lHTKgM0qewZgVHKd0nxAXPw2I+HriAcI/Ugvz2gKkiD1
PgJsoGr7xvQQ4QJwz5z41/lXbHzPkpVXZi2oa/KQ3PTtbsym/Mr8oN6JhCF5
NgpAQ/OOz9Z02JeqeC2deposKde4qqTq6Z/2aYEnhq4y1jxR/poBHg1es3QF
FlO2hrzkjhUX66hpZ7c75JI27bt6SsxpjuFRvfWqyNyf42Apy3Ft/Dpe4zgB
GpUXcqn4EkzA05yt1/0o9AEYlYqLKt10AcMEu3Zs1y/tFup4PN0aUIEyxD8n
jxYayhKivBcByQfN/yDas3mNsfqTcp0CEZYKmAkAI5OkObQ18bXHECtl4QwW
zztLqXdQ8oM3qqLPZ6fPvJ6nRoLMarEWjgHre/0HgIEOPUSjZHbloSQsgtcd
GIAuUhjKr4tZxB5YzHTpEbRnxK1B+lvx0RtP+v69m8ui3bxXdo1jS+iF3imR
VhdMUNNO/ZSzxXYjBmbNutLj9EDWkUP/RkswAfy/yblt73uVbsu36XaYYedI
yDbFB8jSFIWETlFqKozw6/tzfLoe1KOwc6aw32Rjsz+m3AfvHyJ5gy4/M6zS
+cNuJk51H7icucGAZGy/XXsGKa+5vFEqyRA6tCPDgJEr4OUOGwh+1Y0rrDSy
4sNHME5M5zxTn9mIiMZi7azf4PX76OTnE/Z0zeFVHt42tEu8MqTuIWN1YKi8
P1JqRndhbgUEdVq7KM5MUad3h2M/BB8EQ5d9yHjBqLnQXD//I2s9GPfJ9nrt
cPDzkrd6TWNJjZpfAkhPtdbUgc0iRX9ab6dVoBzA2xPA4ThpW9tBu1Be79yF
kqe7MqbM1IwP5O2knBEYrYGRZqm/0FEKFCNN4pHX3AOvlIckeg42QWSysVKk
8SE7xiNwmicbLp0JX642weTFlpEnFeELGvDYkxaM94RX0k53cprTnP9vvllr
uiohLVH9OOwRkhfi0XSEdmsTpk71CqH+2B3lGIEsJQbqoljQhTY3ETH8K1ZQ
OSJIX0EnxQtF4KC0ZtaL1f913IO05pOySzZUSoVvJKBpdPYrsSuPoc5vNq8v
fvwA+KHA0vFXiW/Z+p2hlWcMuvjT/PpsH/52Zuz98ZS+6/YWkjNwxVkH8Zsa
tkgxYHIY7Ctv/otLNYYTxXooc4qLELE7HE/0t59LVoz429tbP8QDsw7d66JZ
pPmXwcPCvkyjoTkoYVxRUwGB/OwZqrXdJF1Gbqipbwbg3ysQX7Dk9C5aqHkW
KVu9TEjlmXCdNHiROLOMR380Y5lzFAPSaOkT8i+NARpqvIuWVqNushmTY/SS
E0LVK136102ms0APJ835BDkdyDuy+DPJqk3t82ITZSao/SoeI7V1yqJPqh9N
DtnOesRwQpEXfkbU5Dh1JKwvNj0Rd4bRqyKnLuNEf8yml7Fyb54eRv/WeK2M
4EOn8UxmEEppZp/LAx9mFpYunoYRKQK5cwhF/szP4Z76y1RtUFywP14zht6c
f6RpQCFXafJsWm++UufLwnjQwbzLP+tGtZdOGq0g0rU/lvl1VIQb+1k73hFT
E8HSZwlksru4zan9V1M7V3yXS1f3mCczqIIXXh7ar5dU2zTZcxLi3nc7UpZ/
0yxctV0XzPjjy3UueFo40AURWOlqUtUBCGzqHPjvwHE9kuZJu7Eiq7E8qW68
DJKI6NygSR9tCnasWg3/8OLIgQV+w+OynUSHrS82pPUD5jxAf6mWrnhwMywZ
6EoT/Ub6rvi1lN+doo8qJhaaYoY6J3ATU+732GieDAOaQxGCKNiRbpEMkUNk
c44DJH92QBOolp4OuIehwv5AwhEfLGnSfZ03W4l1qOK8LBvKzXSXDgru11RK
xikr2kioKF5Zq/q+jct8a7uz/E0pr6paO94YKZ5Ri1VweUuk0kvr3UsbANLW
KBLQTyn4X81TTdPZ/1ZvzkEMYgUXGNYI6RnXNmODPhqFIddnRAxQZEhNhS7F
Zzh+8xcbTxMVKjfu3k4iK/OYZnTDsNsr2ojQ0CfN3VJfBmz+Y0ohJxx7k2LA
uc7VgWnU0mYDlAz/m4q4nl5ioDXE0RpAF7G43etktfAHWT7K6SHtpasme/fD
J252x/dzSQpPeEdRDd0HCY7bKUiZI+aG13fUL9bgdn9hanzwqqFjjHlv0YQc
hbf+x0++jBR/kcCi81FuX+QDQ2H3vV/FM9f8bZAQ+n93dK03ioF9RXQzAJcz
38qXcSvrvwtcd/ZSrdHTWMVZZBwElrpFcKmCZFYvAMKkZkAvmsdVw31rS95D
dastrdY/o4LOtCTvUrHN3RQrKWx86d94cY5M6TP150uQQQZ6HWwv+n+Wqbbu
fUlk+Mjs+N+ltuvXdcT26L+P9QKmd6krne3zxkr4RKb0cPVIDIpI7gV5J0pE
sOu/AHE6fZWq549Tki4dZ753AGCG2n7FAHeD0gqhQew606zeoKTFN8CTIIGr
rG3bcfK6YyI7m5wO/+w8oSR5dWJTvMrw7IRsiixTcnZz1009h5Yo4x6AHKHm
5HR5NUrWzFCYPTvtrRfyO+SkTwP5gsTwdpqTNA1XxbLPSYeoBckhcejbQY3Y
dlqqxcKpaOpryqpjBG2e7owjD4GJOkY8CGP5THtMnGTOwgZQsolDvIM1dFJP
Xi9M8UxFvnAjX9oL4wW8XHSQshvcLF1ahE8ueKIA6MBeMBfav7lOE5XTV6DC
sWUgWMWIoq7Y6QegDF2yHJbwaMY/d+zw7hGieXisOdbCHm4PXj6ZO/A1HDHz
kmgHD5NNXGjn67EP5MQaXtS8yRMwwCbzA5v3wX5/z8wkVWl79bQAHhzn8+q3
TbpVlOS/oF5F5hNkOM2uTQEN4L71CPPvwLFJCrQSJ1UhAJiFzdySHzDC73+I
5SvpnTb+/ky5WHuc7x48Db0NfBBdx4jBSTYCCfm2e6fkTgRskMcAkNTnn5KY
WUZQS1NJyk38cenX7Ydcnx/iem+ZvKD7I78RtdFqzQJMCFy1w3yXGISFR1pX
OsNXXyPpvOxS5W/y8OVE+xSnSnsxJO/34PxZa0GThhFtk4KMSSg4DI8ku0Ld
1ku5/mL1HlEMAUBmamQzsCJDqansRr8JPO/McpatjAlbCvdWlgoIGRq+Qc5m
uZBURuUYG+uDFXdO2+efP/POU+yiFogJZ2WTRIVnbpI9YetnUNvilLkDjG7b
XAgvahn/xozcVIGLKLQN8hlTakxZwpv5Ql22QI/fsCxClPwf2VmmAKGiu3at
ba7phd0/cYYozAlp/9Q1SqgSMkkOW5Qyy1UEKHf+55YkopiSwDXEOR0L/9Uy
MNYzaPiKb4SOO418klXtKCb5bn6iZgjcr8F6hYHuO6fMosuCTjaHt9Sa2z07
aeq/cAAiZ+RQqPwmTKFX+aqZFbhEbyYiZuwQTIwemHuPXEsDoF0oUx99x6OL
SQ+PijYkjq1DygonBZCKHAlk9iHcZyHNq9cG8b1ngrrGTQJ1Vy0g1li3drQ6
jDp/3N+r2BHXytFUX8i+Z/fKQ2SEsiKhhBm/zLXYSEr2Iod9nmuKJegC/FCI
g9mqwZK2fx2DKFXPF5ljBG3Vc36cAdloSGUx8RneHGBB7jd9pH0urEzvWdaQ
ZFISoknv1v5XLH088OEae08VW7q760062wQKES4SoPdHWYjS8n8wfaaPRgu5
oi7/GjG+2RO6zMgYokRZRuabRtNpEBYkumyDde3YOIIhe5gOLxGA2KhnJGxv
UQqVVYeOt+W3r3seJnNSakVf0Zyug80JjdtAt2+pi6qpj+1SM9WzH5GeY+HZ
a1zZtEfMHe0alzB+F5rsUGZctfFWl4yiFoFd06R+sGGz4oGy3tC52hXakIAe
S4VOYKAJ5GUx/VsjT+YzKW5Yq+fsVkNc13B0CoXzzvO8p+62OW9fvCyNeKH0
dbBvYSsb1Pjfu6u7SxtLfsBjmevZIaH6OJDD9BU1t1hctML//a/U58QxVama
8ss1aoNLbScDJPHYfLjMfPpO0gHpjbjnGYtOx28X6D4xYnLeHecPlBma15YG
CWAH5rDA0/C3tXDFvf1oiClQS3xXpMtfeIwEERJTQs6c0e0S1q3+EL6WSAWq
hajY/4Jq1B4YArgtu12kREDlB4KkpeAO736nQ0ArqL4QsjjKtHCv3HjC2Aa1
kGENLpnFZiNo4xRIgN/6dojdCE42bdokkeZF1a/SIPQzNQR++/wBypv6QJzM
dNm0UfaNAGz/GYNPQOuW7MinI6kGqufQfJh99KjhPwiG9bBtTdzdT77ATC/d
CxuXUdsRU4qX8rbw7zSpsJk2WCEUzpgnK4t55lv26HEmCqtw6w0xtynHZRAB
eOWvVCIDlDE/1Fi+EKPDDxlXZ75pG4u9++kbrDKwSZAlueoCZ9acDM2ZzFia
4K2u1SxfQnzQJtSznsYqbjkNJjj1hSQR/6Q2ZoSffxL9U+HfiD1E0M+pTIBg
Q3WtMJ+uBPGTQgNXAgJI8s9KlbXPsN9SszhDagIQ4hf5WuthEzCbJ9XAGDnP
vBifkGGLNRtr86eY1h9L7Tb/nqLc4WTKKuzmwDuq1MPMGayuma9KYxW1oS2s
1fT0MlajSKvaN5UDyohdCGq1zVGa6iDHPm6Jc0wsD1HmTYQuZgEPNEDEBJxT
n3bT68PG8cAXEMWfZ9B9q1rYv7b1geUxi4Qfjwl6lJ12uyUPKUF0TqJtaGrQ
es8/qHggqopdNDu8ctRdq7J6997fPOcJfep2dShirtJstSc3a7xFz95W8ced
ID4X+d1Cr53Lnzp7uQuJxfJByGdxzkMREycP78ks2hwlTeWJVnMZ4RXfZ7W0
byxmGLFoz5YDg9jUIbAeEtsbKKUtMRjwQH2BKk+6riwJ1pyoZU94IQOsCFSl
hSr8rjftx++iOzMyVuJEpKTu6e9QTJr1G3BbE2qzgIdzgz6+oxri3OebTteS
kMI5/mbu7CqL7scCyVuCHLZ7JO66hhhr2saxiam3+Qv3ysAgb2jo1jGePKbs
kKyIFymhAPfxBwH0PgzG8YaOI0E1tPusRGhI4K1khKlsFKXFYz3zmTedF1Qr
YtqzPb34iv0QkPyAR+VBniJEBoiDAANA6uIAiWSYl3aRpyO+Yy888s6Z3vU5
rVVElAQ313B+sDgN95ZqoyhkdWxfKB+SWMTHWB7ExYzjcU8qUpz05Xdbh4YK
ge5QJ1OEGdIyyrRLK552Ws47uluiZyItzNmPk8o//VJaQaX3xN1ABkfKqHt+
caWxBwIL2m23SlEgJyvaHuYvi6uiav+jhA7Nn+iL7lk8LXm62BQu43hudXLx
NvxJoJdusSSSaeHa1mlMSEJa9vJ5SZpUbonQ4QLpq6tZqmGx29OUsMLTHQQo
r2mLIVn4yIWkXvoN80ysApcDtfQQ2gqf8ZIQRGEscFfqrVddcqiF1aNSJJfs
mQaQc7zQN0JE0YWFxd0ji7f/HHUz0hm9DDccJTK7B0asADOn46pnx/L+CJMG
JsDKCofntxu9cDSbXpdOOoL6xEjmukUsd5c5hyZFx6/iTnycJF2M4oSmdj9N
dRD1gEKuKZjfms0GKpMe+CkO2232N3L4+sbmdzq/WK1Z3BNm0B9paik03S4q
74gN6iMUZrCG2dmlqv+suJWZbEZPKWDVR97RBYOKM0bzHeVJVNN/2IhcczxL
m5WvBrYj3QvY4WRGvhMtDLwXxBUWHH77bY1PsKkTdH2/QJWuRHq1pTYqMmSf
PHxVOYhHG9+UmbMKk2a3fw5BCwfln8pBVm379/ztJOFpyGX34qRF3BHXGqZ1
s3SuBR68rHNj1bgPNXAqXjUpXSf8PV1G55b3OA2TCJdsrZupHfRTUk7flZDL
S5Qbta/zqNj1ucg3l0PnQYI5r7jG9Xp55blXJW47a5IrlmJdnBdJRuGtx2cq
KrCImSr8Muh/bG7Hg43m71Mxg48oDVFO3L3Soa1a70FVshxAQYtkVyrVgNpv
G8i5OOl2FoN8qH+oAN7Q0XvjZ7CSFE+aEEKRMHzXFJELOXikFP/FfjOHZH2s
ghGe9640sCioSfG8IeDvfhO/W53N7jwxCKnKZaFNJlJW7d4D603zYMRObyLS
CVdet0Ynu8MZyPCTvvsIPogruCDjB6fcuXHjTo+KaJZIWqPHK8pPbMHQ8J2L
S/bwSwHKipmhFHVWH4WAQBbTvG+05wbhrCjE+uWGlxtefO/gt/UQVbNPpGKh
JIjoUG7sEUwJQHt/uv79FpehuhmGOMWY+q2Gw+zxzjE9qCbrraCwvWydVKnC
GpVpDiWBFV9+tCScPfGkt/V5/z829UkjKXipZGyCrlD17aqNuOhLuhIt0q7t
XBUZVaiDvUPKnISudHMlZbFABCQ5bpez6C6lTJflh5vlGBqxhzoIvWi9WGqc
BXNPN/kOHe9pfJBJmvUQj2Ema8cdtEirTTqRcT3zFPxH9CYt+mxEqzYwYfZ7
ctfK4MNCGB5BGXVxq7P4u/piJMKl3CMZhG9gfSlw6ehk8iZLFR2/VEGruKhb
zU9F2mvlc+mw0qTNnQAdo6K0B78l5TpBB9I79mcOId74s3fPcytACJMfBOt/
XKr4RzeOYTb7ma4i/9vENTkjDWzWCn7qhLvEnV4MEyc1GNjtYkAxHh96qleb
HcJUlOsgql/IdjPoITZmkVcuKx4JrwTadBSUumqg+FV1HJWbswm13Tqc9BDY
Mgz7coJ4I8+LvB6KsSMFYMGU06amsUmcLOYfFg54sm6UcPFwYB/POU61y3uO
b1kZG2bfGPT/bzdU/GCjUnJA95rwQ91r4aYsmq7GJnED3FO43k0lXZ0g18Vr
LbFirgyV5t6cTwb1iW356L0rBjPfZzBg5uEBGStGl5LTvdau0phV67cEfxVW
ca/gJbwqzrEzK0OEwGXQNmXL7hAtImQA800a9ciAIqGDS1XG1GQWBCPvDPkY
9INobfXYvxwlDN1B/qU3OcA/mc2pzMQldYrIcqmaLCeH2i10cK8fRJzLr3UK
6+qDyNS/7rLrgDJFLhN+6186dnJ3sceKnD2HLwIVh9hzTe7n2QLtv/T+3xig
coGkYstZjwe8+sbXdFa+0aFm348BTuPPLdSDk/5WYvYfVP9MMF3mFoLln9GA
bZ+HYbtyzlSITm8zeFxo8ySmvnGAk/Zs7XM+7c2n99Z/imIpOL8ANXMjVsTH
pHorsfxPGjfEd2KvN3TGsbQPsq1wkmYnSrecMIsaLT9F6LqAlVDyVOlmUhdl
vm6n23G4neNB9JvGWkDdLYX3shcdtHpQG+PE9bsF0jBDQSMYCox2TpvMq6Sw
DbOsPmAWbVZjaIUx8/0s2V0IeIfk22TqSd3Xe0QFqAMP481ZcUicxCRTuaH7
e8p+/+vEvf/+KWzn+AMiWMb23deSkrObVZE+g0uu6yy5QOZZ8HvXrbmvjSIa
OYZGUt0EvaZVNX4ksxzGuBY624rL4F/1LQtSxgjgDDUcyqmgruun5ZpU+A72
wnOmdrYR4U5O46YxDmvAGS0fOepAKPg49vtOacMZxoM95YjxywrTCX3telLg
fe10wmMDZVxmyOr2aS2bu5J8HWPGu1+UwnvcnxRHv7cU7PTnjYnwo07fTdfe
YCaKveH3R2KVAlxkw7TKWwG01jmAYFKMZZzN7r7g8AJObxpT6eVTR6KLDA+E
MDuG4OE+W9bFd/ASaPeHSgnQNNzxrh3IObyV6qVCmOMPogmUpIUwVjZNf1f4
KDaZ9JpVSqEbW3BYM+T9qqhBezxMbqDob7IrAYHFePr1WzV0TTGsP2VG9jEv
9R6r6AH2lIAKfJJeOxnCPtfdVPgHr0CfzjIN9IrvYhPeoq4zRq227h5Lr55+
3XK4RRTJdla6+bAtpi62uqw56zQaza37/dMdNWA3SLxi0W0HMnoHul8G2Hkx
73fjEsWUWYAoX4L9cym82p0Ui8A1jqcHUXhYXek6V8BivD49RZN1jWQaxawh
GOn6HheQVG50hYYac6lgki6JvaFKejoncexvH6yFN7/7Q9e9YxPstmVxoKPu
pKGzEZNr98HKg2ORN1sPWsYq+bf8qZEExk5iOZVpaVmz8gTYO+tXrukEwbd9
aaj6G4qnswul6+ujLC0swpmk5ee1A//J/cDafa66lcvrzRDDjiaddCSq+wjS
UJ+PFmolVVDozjWvmR7g2XmFO6pXYEj22gOFcL3nBUv/9I21MXh1VNbtS0IU
dyGrxrCUHLikeknFm7sCF/XZVk1fNvTEDRRe6GZ39gZuoQ2g/KC78UxlAw6J
VOKPGW/f4qijzXqjt5IFjROqDbaAY58QHswMW0I5yHf71H0ndZPgVnEuIByY
BLyqy7DOCV7WkK9jsqwuxxjr58KNBsqGBqAHZV5p3MlZDtWsUSHw0BQJJTgV
BO5GEpdJVq5AAb7VKl0pkgMCO75wbq+9wDXdUrK3eMBAQVdxSJC4bTxAy11A
eELEIwSTergZOyeuo9+3BUt8N4UbX8fqBrXfTq7KmY1Jb+DL5nXYiHRSsyvk
ZqMB9Lx5CiCcA4IRGSvPRVt6Ilg/NR5bOOizqTZF5b3atbZpsJCE+hJZaaIu
PmlhOOVgYxdinQKgHoupcJsu5uUOVnMOUyZye2C5h/kZS9hSx+CzxHvgyHv0
Q3/STQwpCVXLLvyHH2nrh7ftZfmTZmmEBVPf/OJI+lj/Ob2Vc1EZ//aMbVyE
h19RGlWijoflY0LjKz98S/VjHGrAtjlhI+xnanB1ZQJzvy3L9HwvU/S5x5Rm
bnv1jfYCCEMxplM3iESdir16zi8z4Y2CHVUhGxTGtHr1jdyyDgfMHaVvVOo1
9+wKQkKABCqo8F3zAW7W6zuFv1fIm9yAH9dTDVwTNU9YcOewHHzoPfQuVonx
MUL/uEswCiIw1Mn6dEXUXO7vw5SmagarcH1rJhE3WejtzhWv/ycmH31ATxxb
Y+xBfclNkKk3Wc1Mux1IqRS3nQ67c368cq8sJI0d8NP1alBPFtMobcj311Lq
7GWy4PA7JyPgrzF7ELuQRFmhDD8vzTOlzjEvy2liWfuwxWmqBTOpdJ39BrLo
9Y20555w5mTQWVSgy34RRXpovB5bTNV90NmkYGjmF8I3rkJcfac5tXSmNuTS
UduvcHtgewrauZns7Ytp0tifVh5gn4X43TpzATC6TjjaRxIrDMjBrlS8KBMf
XLJ771QhnI8gtlcUNzXZIIMxx5wqrzif/NVGA2Vct1XGicUeXKLMgRZhHR3u
kbKSuT/TJGTD9RhxexQ9taoYf0AhR8QJ1S8/5v4RDGYubJnYcmlEGyugwBeq
rGfyljaTO/vE8KMbwe+hwRfm3k1KmCVXcvvm/JS4QU/EXvB9JRPqww/w9mNO
8YtVkq67sjrr8rlZIFfW5aYEjrxnWNDYYD3iCE9MvqpGQPwxcql+JC0S0gJY
Vw3P+HYNgG/07FnMnJFnY1lxBBQvf4hSDYtxIvklsh6SiXra1cymFE1dyKCM
B98BCjhFcwPJ3d1nL27rz6M0zpORLHlOGNn3/7h4uQCIoukhxAv7/Jt5xUmS
MhHoODCH6rMQl5Jb2uI+FITqLC6/B8LewW5HH9YkmHc8nPtyIbtp3nOGxPB+
06ylHxd0sCGxwOHU5ddHWmWHyDh+3fZ4m8fp1hNE5J0J+2keP9f/dzEqJFdo
eLFD4fM9HuIf2dnyfvAuaKzNUk5em/+M9wQ2IxVka45IVlZo3hWXEzcYSheB
4egY62nYsVgJBbfiZ0z+bS7pRt3k7jhsET6SycXu/S5Da9fFbvfuLgFt4ilr
1mL/vP077q9+qb5cISHlmGzPEzfXIzfYuXcZLyrsyxvB/SJNipx8DOMAnKmc
APwO09vqOrBqjTIO0bq70+rKRErcXVd8RSr0C6vIlO4cq8/z8lhbxCQtJ2Wa
8SAyFEW4fro4hUScl303Xfykoi88ch07/jLEptgLSJS622553GEfSyNz+yKb
5Sdzo4btmXTeVDmJRA+snUmexLX9xkPJCBJIEAhpZxr/A8sRxPVjkOQ17xQs
7bd7XBS3mUfsRvYABKqvNCEZUTA8/o0eqEUaeYhh0C7VWGpgxqjkt1m1oj3O
MM/J6/m8hLmfgZ/KtjDkSTdBZh5mF82VXSj0lkYV6R5QiLAhLng7EHJsMCjj
WcYq8DukfXxXzfB5BfoGU2pjGtn8Ns3TItjCeHyHoPXWkBH/XRlKTZJW6KiE
Iv+C74Fy2KFRmt894oMUi+Y+r+e3Z4CwXaz32gLN2mh3Y0x3LQ8BVjFl++2T
959HxsRbW6uWoPBlGnk45u6LvQyqC1RGhV2m5SI41BqVsT6oiEIeKDJky5xU
10/UZNtSM3pL+/0KapnaMltqfYuMBPgfN/jpPj1LawAzwmhHe/21Nfds7k+S
Re5SI4nU4H1gq8VvWn62vAiBu4Wj2npFZuGLTtsTB3eQYD8zc5iqK/pFgIMy
nvVTdEX2uqv5TQs3HJYoJ1hvbr3c+qf7JnxkxiT9rj7c6Y06VM9KL4Mbx59Q
qeCZCAlpkzflpBGYSPmcdlb5J5j3rs+d1lcN8DHR3jMNYGPFtspoN/cn/gya
viB+XvEm15UKhhvAJ7AS4J18CxcfD5Ez3hAmP2Mv6tLcFKIvW5XhT35vWA4M
yN9FT7UheUouCmfwaOnkalllsXP9yNp47TOLwijpH/E/Q6MqZCrMoVe+kq00
5jojA65JcmciHkfcfP6LaW/1ziqIl2yQHmEnu5QSuB18WZNbpOY2U/+BF44i
SHORZMEFoJucJrT9VQItW+UX6iKEIIyu+r374/kEcXjg7MoXD29n4PTPtGbs
meeSJZC3U2CIL4m/CQb1B2MwImjP4mmJAHr4Awzl1KqhrKCt8qBdHjfM523O
iTN/Y4fAmJgPWMANqZlBjP7HrA+07dOBabxEB/+B8V4VC8MR7WuNYGo+9Ovm
oanF6b8C8KCn03br9HMKO/ZOPQNRiVAPnvRM0xD0P9M6llCu6mBXJ5eoSw+/
JMz8KxZaBegInhWrmPwkGSioQ4im9WCIo7JfUxz8Yr6Rqps9Pw4+WULaTHOr
v8DFbED9zySoJMNY3A+/fvO91NxFl0GaYNzFgZLyPaAratUKtUvaPdadwge2
mwXG7XZ4NOGXEgcFSH8+6fm4NFhACvTKYwNpQDvj2h5jiAvI5tmsNk+NLA8t
vGL3KpE0hCoY48ic1pLrPQg0LhIaSYvZqBj/O9Vvc45dHiQJPcX+riHHhV7X
c8Yzj0aaWw7XR4+SokYbyPInH+ASx/7MAlgMsloMQVHBXQgp/GojrZ3f3SlP
OTj1fHPVW4aVyX8BBUzADTkWa3lWpuSkMHtasi4rSLtF3mMpS4Um/ZiuQctQ
9mVyYP5lXw8NaOvspJFN+NjP5ybBUwrMpX7Yf0wZ+QgvL+UgurRqzoi3MdvF
AmcF19ABOXf38l/c5BUFpYetq8CqYtSjxSHEV8Q2IE4/R5MSrA5p8ugOB/Ce
GZ9FR4KL0GcXsl6gcQgnZzZFyD6qvOZV6eTCHEva4TMB3UFURq7sLitOe7o8
bftneVJizE7sms6uTZWCDkv4kJGclMm+vp4E8/cRLiwj8AhyejLjMWPLsOkb
/uCmEEQVZvbL5IQpuX8ZWz8G2rbTJenJ9Uum0y/boZ7gmQS84+udezt1jvHW
qTcNHaW6TRIbfKuIx4oJX9qQnN+silThsA1McfydFNdi6wOuhnok6kMr9Xb/
FfZdZHnmUrUxtpc6A0IaJemUZlU0qe7tOsRNbrL/UW5gEazpDQFOFDBsvcLj
NE6DlHLotmFr3ZPYZol+mnJpbGWx2Mr9icSZgAbx1WTaW8vtdnFTIojjGN6q
n5leD0i+TGnMqXFQgorzA7RLL6OVIDjhysydgjIo4wgY/CR3CaE6eYNnAY4u
MnHcAzB27Ls81c+mC4BGGso9ZWyvA5/lSch0ku8Gukhe1gcgK2pK0IsQfdMj
f39BtF/AesvoN+sS5/K1li+TpYBXymLttDi3UR512Rq+RkiG2qD9fCfu7MSe
y2k8vqhuyBtnRvIvEYTk3da5AXXH0O1XtbIRZLVWZlK0UhEXz07hSOx5z5tP
bLqTvwn2AdEmc9glkPLPTnuxylmOJNHL1KfKVZTSSzSCPoXlEESN5EvyFwE8
J/cMyJ7+wbyFhBRo4neQNUGxUl8oGV8+z55EyKFjiwJyl2ekMRUHuz2RLtfA
y/5n4exXBt2HCL3qemvx7KjEcFcUCNIj0lc5X9NuasTsn7/Tw/lGkd7Jreig
rr4yXPzDUtbNoCWjinrW393gLsplkBfcA4M5P/KIdN/ZcV3Zc2LNrbmdPfGD
qLwKpuqKdEVXRH/N7Apwko41V+qMbmd7rHh92rJqVlBQy+GaXMDRbRo3Ky/b
2i0Lahc3zLgh31Io+abD2ZIHYrwROyILT6F3B88KBuxpuIfd0Q1+a9EJWsw7
YfKd61frKGQKdY0pgYgL89694uVJsJGKFBp6IYYyPAjglFuletLezGBbSKGU
4EjgTtZBZx2sqdJ9qZMa2LsrzWI4tlSiCv188gpB8ZTv/5xKfEBwAVdHx0n8
gYRS2f4r5FTQoX67vbqaBUgiDCdZGkeWBhDA6X7J42uqQhVnm7s+iH868KEM
qc0/86K4vJZshqSESOt7pYKMwjFw7epjj+GSLtWxlU2ICGXv0NTi1iPFrdtn
fXk/VZdGQOLMLVQJ5jSO62IRY2ti4OiOiixK16LUxrVtZ6qWK9JS6ULiAGEo
1F0dA7EIwlhH7YSiY3i6Qc6b5YUybJhhxjMT0naGncPISCXYSA/UOxzP35OV
BXQSITN/0+rEWRT6JQg+gNptpYJWBfh2t6yQuKYUKfrHXZ9siLLOj+huI4bo
kChNVN6YxgBA3IOpTFUF9ZjlDJwvYr1vM+jwfQ+QwrcSDgU7TrMCDS2yp5KT
ylf+GMnSpeXTQP5wyzLjXA/JwGTUEKMq8t0yzI8y/7pg2dWQByek7EEPnQzd
6NHWJ6HZ9UHwHPT+dffvfMPiYwe1m/YdFEIQFLi22UBNxgMUYy1Rc4oY35/y
haHg8KSu0WfJd2hhvbCqVMCxXct6Muuk3yXOoteKospco6gsRh3cLeFm8Fey
HVDlT1Mynbp/Is1ZT99y94oqAzkYb91k6SH9jfLFf2wHGeQaHuNucAl6vddp
EYUhwNYIP26TCSBn57U6SbnngJo3gm2cBmNL5xLZw1OuHCx+o7zgZHyo0xPi
mbMUjrWHW3kmgwcqc+2fPsnFdiQE+m+ncmYyq5JCpdl+SEHJGBr+3lgbYqYs
GAPgmIBC6JhUuwtckAXBP+ZroEzm4nJ8AXN87f5nu9QUXuMYlzOEIC1GYiYU
iUMmqF/9g1L4Vvg6CwYIUZ0yPtv/qPotYCBUb8MgfFEF5JC6IuBdZVjVIUCF
D+moxLNSCHyh+CdYmrBSVE3vUgGwF0Yr3RvauR205el269emuRscw3C64mF0
5XNJavD1Z+ngIPl5p2lm03OF0iPOEqjv71dheJMTyAcUjk8R1tdtf69LowMy
EnOK71AJhUdWDf9wx7lAf0pzKWIqEcQGMujK3SM618ADIsQIEDaEGbqUJjAk
rxBUaBEuDoIEXJ260p6KpnibEC5UbpwuK30aoA0BpMSFJefuOXWg9YO1J53s
mJg8GsmkWidOCpter68P1TiAtp8Cp5pq6rBNL6okV0BuxofeVs/tW55AHTZ7
Zl/AEG51GK5BBuE2ezLpGk4igAdtW9vRbnbm1ny16zSC+bdSky0OhY0xe49+
SwNwwjG0BX5gk5HSDqwYRD26rfrDhHGK0d3Ym11jrGtygsVWVrbdfj+uKppe
MBfKtMst9i86vZnzWGiG84xNj0GTlePRn98QpNrJwgSUJBttp8yEVJOfzvUL
EsuFz8PlMXAluiGzsMLIZTkO2PtxES8o+YwZTCETVy4fkaldUj5QCkeq4WHr
Kgnwn9xyNBnRv/zA1AUZ/h8cw5D60pi/dmcXdic3ogH0xTX8N07uWam7AGrH
gTdeMiMZPsiW24LNJ0Stbar82GKPrJzICA56+iLRpoxbYxNJslLVslL9oJoV
mS9U2MIadGe98WgbJXe/W2+eem3deODhnB9sT/b9aZJuw8nM9a3wE3Q5+1/3
MjeqsV1q2/S2uzL59YYgyOLEpoeRiiU8b3RFOIdtRmnRjTIOYMZCqQl12ynE
/pkXX6m54nQYe5L5rCzRoxsP5l1HUGS7nnUwEnFEpR/HIjIWWvkjCDNkKOGb
YKMU5BF+8/ymyPFTfgr/a2XNqo9C2gCL6btpsoZTOVtZk30GkAb76F33BJBG
ch4p0PjXs0v/m/nEL7UHBNtG3+x4DDC8m/AwgsdWrfdLIItQDEDkrZT1MmLv
I/CSkZCex2BoaYPd6LKXF+ph0hRqkYWjl6WfBRm4CZtWZaoPD4DlatDzxB2f
8cDLF+SmuGUnpdb2DrogEMkO/ijGH+1p7vppq9neVfRGbhahfILFY81GRX3+
113PXBaX8YASz2PcnEdDfmlane2hhXTQd47a9WVNMWhyZvd94omAuDd6QKcp
2Mg9f1oeZXzuwFb3Y/c9Ld9J0CUXN12l6SDW4GYLEh6f97GCv9H0NkoQWw+D
4EMq662e+VGS+VKT/82RXotgR6oKZUOwvmDnEjZHOw+hbIwoSR+iAldcMQqS
w62XaeonnD8G3o4Qag+Mrdu1J1I1r2b2BfWPmFkD4c0LWHWDKl3rZB1vyfhP
Xte5YvJ1Ss/hg27f/UE8LvmssrdDvKD3KaqDF+MBskfOOHM6RhsXIn1HuXYV
YZu32uRFWSqV7YQ7SovSjmZmNf27pkWe8GKXv7fA7Q9T0ocTfj5U8LihUW4N
cw3Oo1sgru87OZaOdWjmr5NQfvhPXu7IY4vOifsKxXJ1tdb6UwnyvkrGAcSZ
mqioVumhsCsAGBnmQBjcX/eRKTth4BPY1R+64FaWb/81AGc8euCBllviWpYS
NKQCUchQt4Xcm/hj6PdQVuU3nOLNj+FPLdcGJvk/dNMHlWbEspQC8B1ufaU1
yJrM0Hy7yI6jIMn5h1TMYymPHAND4l3xCpDyVBK7tBrBDCBsj6c/9PX3ni8g
2A8dMFCEIYy/0goD56ClL0mfrri06Ujf6nZ4cHv4EyBOdLZwmacphWVOVO9a
eQCcaJBZxzQTp0AyPB9x0mVSA4B17nxDorDlHShoP6JgkGi2OxkBtY00FCn/
BP7jcOVH3f+lKFgeVlphRdSkmc6PfXWF0ZoGINGHNVlSd2L0J/H8xsws2gZL
8BSqa3HP021WvVFzGAvZz563wcOZYTNPpCZ4lquwr4LQ9cWdkc8pxeagDfOa
7SeaTrgzp4s3MxocOEN38BM2UJvwMsA5kwchuG2rn+v7EHzUa3gG70Kl9uFm
YZgUMNs+/HcdvfQ+trwZvgbnhgWD7V3oZUT44+xD0VGjfhbDY2IudUuNUe1i
J5m9D5gp8CUNU63C8pPA+bNZ90SYzuP7aQfRu8mWKqVzQ32vUjhZtHcguPJC
eN0SmTNhMXGlr4TWF9BKh1zFDqy55lYVY8lGKl9D0LNv6fxdxaA3mrsu1ZPb
jmQEcTizlNu0js59nqFkcGiaXwavHdzEUhZ4nXF/mxUBEe/3pp9kTWA89bMF
E302XwZZKkPWsGVe8aHXU1cyr8bJTZa1I6TmRJmNucA0dnStwnfArpbI8xt1
xLfpc9Joif5FL46KogDHh389j0ORbTb7UVEiNYFq3lhrVEwtQ3G9+h0NxRb2
1z66xi0IMHfwnk1WC4QKnznjwDUFaP/IzPvJTwLLmqSGkAOwbPjMDKCcqLMo
Oupl/xHzdqrPGyi/4v6p4Zx0Qv7c50k5QQaRbjsik3NszVHttOKQZHyqAJ2H
dIhUWKaIDAzbV/1T8a4jQeSKtR8AtC9zlJB2GN6rEBg2IyKJLaOhnwyGYOSJ
2VOHCYmnWORbIiuRAVUOIciEtFIis7vskE1hpMEF1CsOxSwcfyAvm24VKGBf
BjetC3kAwEcy0/J/pAJ5pDjJzK9h6kO8caorCsZi+IitMdtYFrZoo1Drgb+x
Oh1EkWWN/85iVwlLvyGI4k/DLn12Xl4/IvJoRkCDkVpth6PV1QFjdnTceyyE
vbHwjQxoNqPlRaZQj0wDpJ6KPRNQeEt+0BHHskZShnVZdNXPSINWIIuJTI3l
siq1Soh4y/cdRrmTwYPvogqOYCvlLrvsBQGLEjaZ2PHEurtyUExgZeib2Yg2
0s7AM6QgU/KgUuQls329li8zSUDRla9OFqSfsZV73AJpfjxgOTVy1MZxVNo4
ch+47N8FNsuLuAMYwoXsxLQPF+BMZgwPg+yPXU9HOFy1QnRYv7NaqzfyBuo0
a/NEjQWKhVYJQFtimoD7C7yyjVA7colPXrlqcvIMJU9qeX+MFwmlCwXfClPD
XzikgTXZX5RDrM1dTT0tWZK3Z4w94ZOMY8CkPCqoW9TNMEzRkG1AZ/VL+2iT
R+aQaK586hV68fZ4O/3907AKeuwQZcF1UOsUACdbt94XpDBQBwIDOAJLWKaE
6ZOZqSu9GnygXDzAyvNDmbWL/71/PeUzFl8zXfNt0ERJALcQb0FBn2fKr1V8
UuophpfXh2IHcc4AYhm1FmTW3B0kjy7mM8x5O5ug4sWikUymvukg6WZjKhVp
aGg94WnxfZ9MYUzn4wPP/E1xSXrMZtkwCQ17SNM7sLjTNN4CBkJ8H+H2w2uD
lCgjUBA7gs/kMBVtNaCCJu/BgoHa5GAQtF7TgoXv3kFJ1fHCGT18BMTYaepC
M8+RhNtrrInHKUugUbQYBTogit5fcIKgEbT1BukrJUqVdXvtRb84tPnk59h8
Wy+ijZouSkWLuvCTHrjZ4RpbgLmsO8VYLi8ZPPDlNEEuM8ymiO3hlyOyXjVb
jovUk3JHIrOBOR3EesxfjnwAOc1ccy4MT3+qeomsI8dv2g0ddhepBqqn8Ibl
2AwMy/EOt6rWZ8w+lz+tN6t9Mb3eblC3Q+fpL2IsbI4UxISZPrjOeNxK7BKU
/31Cn/yuNDI8wabY0hubDgaEYRePJEq1jh76EIUhP7ExqF222463uaK3+coF
F4KCoMwI7zSoYGEQ85HiEodLyKg1CUdHdUu0jBdcXdVfms1BfagBdIw+1kOp
XlMewwumHIXLnMQjjHlg5Ie955TI67Glr8N0OcuU+L8klzxMjvtSzczckbjA
a5OdUlJcLSSYzBwxcy0GebPaRtP5MpLhK2KpAKyNebHxunpSpDJYZQwHWVe1
dzd0E5+x9IlrZm9RM5sIRP794d/KQPb0Wtm+B5vduwA1mPmF77hx7mKHDT7z
DAGZK6bLOYAi+QUedo3XP3AhZFPGiiEPWCD1qpkHPMwRRk+PMTpaGEt2hg23
qcHMzvjcMWfzbYKikcrHXLVSK8STyKL6nOEk6knzw8N6P9dvHpHMG0wci8nk
Fccwx4TPqF26pwAoUIY4c2v5o9ORe4IVs8xYLT3FabJ6E6S2FUlzt1HT/I63
ejwqBs0iYabjze1AZKUYkGlfyMK3bW35YOl1hcLRwidbcYkmHaiq2rW9oyBA
omWfEPy2zMYkw7pUKO01V/JKD/GMhbeCRCWH93+bJtJ7ZEqfxRfEBpln3HBo
BIwhWA36V3dH93W5AaSzuvJ+r8d72OUdjpUgCjcjUk66AxiFRC8f2TXtXuJk
URrY9Y6cSa9RBCJLi4jbAzBRjn38p796E03eUhODAMS4o8BUs+ERxrwqJ10d
sdkXjdZMNk7+Rm5ldKmkdE4CXrb7c6BVKVUJSiQtA8nmbE7YRiAYWPMo0/wz
xBtmLlLsSh6qMvch3xP1xVd0A4l9Cf+GSqenkYcn229ryVSZ+SVWa6cMbz+m
liWm8xfY9pA3KsMgPC0AR+d1KbaCm2LUxR0jFq3qh2y+wZLPBWsldpVWUK7U
93v9R40LTikOieYHX1nfBqLfweswbVR/FlR/r3HP7Yd+9Bk7AB6xwy5MaTfU
OMatNbM18Ftm4JPjY3UnLyj9WPklf/2zlq+93A1x/0XzOW6dlnfj1560rb3Q
A1dQ2g+SuSNYALdBopGQ8qhe1XAebixbg2XbvK5E7sOOXCTKhfRPIGKWWw0D
Be5YHEEHi2T76F8L1NpGJCe9eJj8aGXTxJBNYTFO+HkBl1u3DQM7sjKp1yQJ
Umc5LSnxA2AdHMW7abqy6aZsLkKSorXae6GxXM02MOVoeRRo82WaQzO2WABe
kmLFti/lFheQL/TLoLmA4XE28YFvkssP5KbBXKV71JNZddqja0stebShSD6o
CBIUzfACtUUOMLBTL0sekzG3B8soN15xJe3qwwhn784xWJmKtPBvBE9Jhasu
ccxkUrJ2tCyxVmHrpjZjNBPcMQ557GRgjsf0ayxofcI9/tjWUljewplc6f/d
Nlxdfvae+eDrf3iKsvSWjyGbxHRQRp3hYQIvSqbe4s6lazENi6yrBL+QkuZT
htd00E05tKt1m++bmZ/NpQxeB6gcbMHrFT7sfxeAEbZoW5aINrAj1Jrb/nld
eNQBnYl4ino98jYm0JKfvf+bxBrrPDCkefj0Pq90ernfQC+TbKBiInF1zjme
k4SVyTJBaVQlyMNiwSlKs5gY5GCea4/Jz3bZH4ui1KZrqI1MVIY64J0gt5T1
0sNRwTmnUpI9V693jZa3MZCdtDI/dmNfmRbgn4N7y7cUpTfPVV6QejYCRIjH
ug1UkkM+1OEt0d7jt88fgO/9U1UVixu3s6QfVsqAlWl0X9oMopQpJyrUFcLU
MtkZOh8UD0FHPvBc5XhDp7uGS5gZxWCGCefndY/aeNTEO19mL7aD7hGi35xo
ULtYslQ9JcGyegbx9QPhbHb6KzTQnGCqPGh2ee7iHkN0LSzvp2hM52DGYWYA
TqHde8ynw+v8P2w4sag6Qx1w/iRiYYC7pjSy/g4N+1/yqMyws4s0SFI+gP5u
XdVGw/BOy8+hFr5GUwryqgxzemI/b9eVGIiy7hQpcgJnAdn++6+qoIC6AVQV
mk7rFBix91CA363HYdSMebESL0tHWSLFNfxCtB0wHzHTyCkfpsJ8BUf9+xGI
U9G98IQ8O6RaXOVsshSChIFAqFodF9tYxJhjeA9fC1OovGq6w2piJGK4e8VR
m9TjFldp74ySvXNbkUAWe3NFMqzWW7IvGJvi+URo9/cYJsNIjGwj7hLNOp+A
ifzGUlVK1QovUxlKgHrkVOY/ZJggyhT5ZCyViOpVHC8iZ2Foj707orQ2rZbh
IGiAFXFpS92D84Ri4J4Udn9JKi+mf90Q1J+WfDPGvMYblgHv6TsHx9OHcSB3
JvYP6fPrG+vVylFM9vmXGdOrJmaqSJeiRBYZ0KhPwJdifcDHmVoIyhLdJRvt
s+AS9QaIravR0elHwjJX0BEMB/Jmm3gkKRaso2QYKNrgu8FLLJ6usf3ckFAL
D4UFBb3PLAAL3/P/nLJc+slNecl6uC2riA+MrAjKTsQgWtyJnzDZi8OtNuhJ
r6kgLUdBWadpNk3SNhqE2pQa5FS0pxY8kzG2DalMZpaYOKdrNN1ehmCS4ODU
UsvdkaKwRDR0fcmwbVuDL4KEI9mndJelUMQKvoNDqKd07/EeCKJxoajVHssc
v7zWQuZHGUsgT6bGXBYdZp8mA60P/CJ36MnSCQuqtuh0BxogPbdI5ILz6Xf3
lD+94/DbTPnV/QCwTCXvdp2dNzmWSKjvJM/ScKvA3ufvR418NqUzasOErzX9
KY4bBCYKhEM2klqDKvANY8yzgyksV8L/w9HxY8NxRDEBQG+fv/mEfr1K1UnX
2xBzc8eRezMp/K51T31QYTmZ4QGaKAdiaFP9awFhmNbqzWgwR0QOA+e8cz5V
Q4VnPSLxOy664x9zK27rClea6bXnTshRRXHyuZS9wS5WNHloTWyKv8ze+a1a
ImhQntH9N8eH3zy8PSj2xq+xfV2EZo7I4+PaMCfG0xZnuc4w5HWEmBcf5Tph
+iLV/cusNqAqdeBerlR0kPZ6FbfuZtUPP7WHY5USfMxHpuJ4TtsrNaR4JCLX
9eJa/ClZ9EjiXQiSx1fYQrFq76Oxc/+BBbbT/eLZQ3hSUBFfzrUoumxF8RdN
tSEFNfXYCHKffl7qd0y5YIC/ZvBRguVhfKRATZUOuTRAB95Lit8U2JFwTg8J
tUZrQhFoid8YKbniPWcEKljQvCs5pSVLjUYAB5tNOHL0jOi0n0FM1UMdzLy3
cTcvsB73zVJVIqBwzRmK2XG5zT5qF+Pf8a1qLA0tpFTEOwP0i80oXqne/MxF
j0k+GrrqeBQXrmV0UNcR7f9w1cqeew6TzFAowAZJn4h1AHuuRMRhHbAXHkgw
lQD7uYaJ1CNj1JnZD7Rkh4c5DxhXgjpFvRcpCkzKWh7clfHABbiaF4CiC9aP
2sh+o56qC6M5DDA1apLPMRTqPIz1hqOCGOX7btVkNImrPfR+mUmW7t/W7qo5
Iv1bQ0U/zbFkTImXfySU1vgXn16RNCquU9ipfKPPCzq4RXzHF82wuOctxJeO
Suo4anAU2JnUVG1pLkKiexh1CaSrN1HDea72qkXV2QCgMPit5Qaoq3jHcBhb
nqvgOkFlVTtAl4n+KE9pPRDN6YOHQgyW8Tj1MZcbjSsZbaZg0kf0kQw6ctOD
b5awIUfHV7/cqtvvxjA6uJycHODaSAH4NvjWIVOBKuqGOdDWIyM9fHS9Qd9a
OOxA54HMPxvDWQNnaEwbRzHUBQIx7DlNGH5PquY/prXKie/HJJZbTkUyBMJl
sDw/tdGC0k/LXdb7RICeTCb7hIwsAE4ePOe2AYZPeyimYgKZT2YMWVYlk5E2
OfAC8OVx+lUQyqahYB3YnlCWNWb2RRRFwiGv7Hi3MKzzBjEgPaffR6DQ+QhM
o5bXUEaYUKrnXcmZE+B4wg8hND6fRp+dXdvJakPcufjxiDCvpC6omkMH5yqR
JJf9l94LIFs/bWGavq9hsEovICFrBYOKHj1870nzMOUDGn+gJlmQhgqr30Fs
7WP4ZD3Plml3UelqfGusqXpwBW8cgWhNEsdUup5uVBkdkt1zstch29pNaIby
82CsFyx01FUtc8BHGI1aG+87v4giYeTAOFEu1aqKjT7wAPu88yY5+pG8iTqB
5sRbulwIxPeOQUqK4eQ/fmpB6eQ5UpkJFaNjvGSj7nxLUGHBoq3pzKeNyxJF
xeV5Ft3fjKX62GybEyuvABCE1YLsagaaEDxkrqwdtKlBZW/h5Msge7TbT5Yv
1Ws1JF4/84V/H7V+9fiS75xpyTapTPevw5U/VfO1qKNOM7R5kKYDIhvTA5/i
+utlYjfE6yeUZlwXxBzw59kL3SB+2ODNcku86JTbUaJUkMGZF46aUUMHECNq
qO8BhtN1dUp+KnCy3+0JFhEcJBOkh5N9G2lku6Jn3hSnugVPBXAMSUI856WJ
gOpZVYbzSGS8gROuLvprvDSAFSLeN/1681jscJ7KBwkNQz7j+00Vg4ywgiJh
nnbeS873JdF2Y3Sbx7fkErziX2J/3lK2tmErxrtCIPHzhjdl9Il8lC/2Lh/o
jG6EJqBGqkAiMjwB9n+gNurdUO5cxgKEySeIVSXQt42x7FVf5ocxgayVBMox
EybOV+PPFCVtqj/uZxzE8Ym6FFwZS/EJhYc1i9kMVgft4u06f/NYyH0fseim
fhITGWeNiisgbSX45gc687IALR0Ip3ZuJTXN/1bShgwajiitA6yLWH+HaJ+3
18XB35LSg86Hn8C6N0FBFvbhSN6Qa5lOSMdDGYjj8hft9GaxXwmRxu9rtdy7
eZcNCNRf5qBSoRpDZYPBoOwn4NEiLvmOOt4bdDQ1hk2HJE9eXkLRww9Lj8Kb
3PE6UoULwvHNbN/tw6+F5z/e+FR3dJIdYGvNbpPce4fdM2fyS66FHzGIzKhM
rcHnCKvuoKrRFkBWbBcQ2Bnb+d32ZFhvR2+AR6FI+oNWFlCmLUidkb7Air0i
o81Ryy1EGNdHhGJDc1Z7IT/xZ8pf8kaJUlo1JkxK8o7jhi2qAPAfHtFdwqAn
BafkWmpFxG8/UvphcO/frBeqonQXoQwCA3EoIjGMU55Z3Xr8CjIEA7XFobMd
wANkvyGU9AFSCZXf0YnWC0fUceMlPXZVeQsEPKRv0HDi9EMD+tiyMjtorf1G
ZklGKEnADk+uIkgHskq76XY7y6JqrgnNe9dWeIW0CxWPW9FzSz8Ba4lO0aVu
sbywXCnXfbxXe1+fQsB4mOn3oBA0YNxoppv4nUqN8QJ2HJunlVbOfxYP7ZHA
8NDecSgy/Y6ZPaPao6tEYRWhbZ0gMBeKO7dYd2Kt9w1Mq1pIzZ/x4sP8l7PA
mQyWCOOrbkDpjV0I4uQB+d5ZzO09n2c5Kq0pdmVGed+SzMz2oRHhRnStO9Wl
ucqU07thxvh2nLu2jijO982J6FdwtUWlh3js2w8RKVfwbiYQ9T4QzyLg/7in
XPUi/9av6mochDLCewVxvLvCW7XtBJgnkCzy1C7OhDnB5vFlZcXX6YATnQ8B
szbZN2mguMAqEby/672Znzju84+lJsE5FE8spE2rwBrm6Zo0WK+fgj6Pxcev
0U+xyeen7bLd844zX5nLsx7F33ya9MRy5I54Kwb1hHrU0cQgdGUF06JJPJSu
hGCgAD4i0dEBzOfyLhB8/RYn4FsyQ1s+4cVbu6SQoktoNo085Bta11wpUrKe
Z9rHHyubXZPEe0hx979iDos1lqAQMWIYTUzrlHFKaaivjUzOFe36V0nGJnIl
C6JqpsHvcOuK1D/dI5tFeQAScCqGvH9G+d7avdrSb7IrRZMLNzwoDEp3Q9vw
JA09yJeasdcAPNu81QUzV7CHx3iIp3UD4xvgUh398GGSINxXF0YMlKkxpNAl
zsSy1xY70Ti6ulK0gZOukyak2zFA7RVHv0cjtG+Scp7/9PsFNGtRfEbroUGR
HHX3A5a/D7fauM0fox+rmHSDzZEvzopKIrRmQ0p7v3yLhsaDELX8a8IjKna6
izVRmhD89qDzpB1oLH+TfrHxGGMDjBV7NP0Fx+YlkPp3s34aCqJM7QyfIdhY
/nSgU00n7miLdvX1aNjpmEtZQuuSEI2l/OziOeR0biHCX7Jd7M+zvIBj2Jmh
xzkbUBNZ/H9HnDVeLWFb2LetMjVlMLR3KOm1mLFiz/FT48LiwOMfXBh+Ic0y
dSHjkEpNwunYt7kbDPuT7D16uwf/+0J+66PsjtZnAcjP0n1S56TfMjBA+ou6
seOvFmGSknROrs2x0ZcnL3VrvY7GmIXgEqRq9bp8TdoIT8JrDhD982AlccaE
NykEncPAnI1mVEjCqVJGdDjkV4IBIg+iZXn6LAbmNhUXJIj/51rw2eDbtG1U
blthuYXne/aIEXTmZwcOwCPoLw0hAbYO7hqxd0nBK5Dhh+R3fw/drNIN4Sgx
BQDIyiUx3iE+K/7k9T1Tcj0hnBtJ7Q8e72sgslOzaJrqDCKmwximnmoMqysr
IHod9ShO1skLxhyniGGpNJjKQPrzllC+4SkSyG/+EIdcHMATJ1RZG3RTe3up
UCU2+RdCH1ihYe7HVz6R8xyBLJDmWRrzGD9IjfO7hdGQJLlOh5XucjDmJZnJ
qgQAhHl9NQH3Wg+Vg9aEAoFa6ixVh3Pp3uZ5Vmzv3+M8zkx/UWHeCG+1ba4L
GtWBCdILkragglHH52Y6FripSL/tyvbzeipUV/nsBxRZtFldhA6ZI+FV4vR2
RPYDttHjgfAY5XeDzTWwa4YM4a7qbIRr7ybCXHSfB46ecQxfQ/JdFsO3TmR9
0xbu6ZMIPhGh7OEZPFkGrVmqXo4bY+bO0ASv7YAa9ZKph+fvFrclXz3fVl4D
gqvbbhkdereyr/EQy5L3tlSjXYkjsSVLEasR/ofPHbq126vmmVfqUSpoFUeK
05R13WDu0IU6uEKiJzrNWDu0waOFdkp1guf+qYtlvROdqVqlpkZTS2bg3Wb0
baNO+2bn1/OIFp+oSOK+3mhX1aXfNBlQVuFc8t+uPE7Ci1ZeLg6raNc4ZyPP
4kB/1IVqx5YtojoIwW4eEQIqe8y6+Y6wUuVL2urLUSxbbwytE0wCUXQn8G0q
ybwYDPrwc666eZyNS3QLMDkqxUAsbgis7ubte3+v/9T8Uwx81c++auBGEq6A
D7cn3HSSAFJvO6evRQ6DrXiGe336Ra3IoXXUNIBXh+R2jcAtSLuT+ejD4zXu
xcMIMD/5Y8NWFegQeQrN/I8erCq9ltya2Qg39CZ+Dsa9xPn1YxT3tmjny2hO
n5pqJOgA9XKGubzTV+Pnft/MAwKCpFtIEO1uVqNKnKDKhlrMm5pyQMQyG2Xo
R5lqkbsm8UM/emHN3wY+GUZLf50qMLIfCyeVQP+kOXWR5REkcdqRdenWOByH
uJvamNpvE2oYTzwsc4AUEWmyZJbGzGA0h8OqH9d3ME8q9ogMWerNcvAUGUae
vobVbcqS0YA7ANqlZVBFZRUnaFCnslAvPtFxRI/al5jM++ZHwtAKmRsMu3bM
wH0xfyA2i9DUgzCVxo1PCaFzon92C4fNI/NV7KnHtz/sxDNGz11MUfhHGkSH
5Iv8o9pVw9jsNGGqwXs2saOH7amy7OgkKpaJKVm0h0sGXwIPIffItYjh31or
aJjn7u9b3a2ISXUoB1f2GV23dfLOrs2A9ri03OWm8yG9H4YSp0SlnwBj9ZfL
7PU1MjE9F4TwqE9iP7/yoso2sX+/AnvjS/iEQkqVQzeuAHKmjmJzyno+SmGx
EFL9VRfwRRy9t2ssksCM5fW+EtyvqrjpnJirt7mYy3KHvdU9TrMIf5Nxgq2j
3Pzny6LXvjOBro4Tsm8wRaXBNEX8ki7JuC5FRbgFChREI5IbskCnVvG9ZEQA
IpocF4lUB9whSCD1JKdqAas51XNhjU3XEsjqRhfG3d0X4Y3ChNwWzfiOK9pw
hpeRkWDu7M5cOI0woWT9tXlIExebhjg0/DO6Lpjjs1pXrVBXYcK0X4QvG5Rh
fgTRoki8hkSbuOwroYpU83mtbTOXnAtlpOXbULuCcCtY8KYHXUIbKwfj8X2T
XNvK4SPzL+GN01D9VXrkNGAZ0Ne9789O6SFYfXzv2982V6uJvBUci9FUy6sx
wj9BlnyHNMp77GHUpRCX80z23Lh8T3GGr0OT+ejGWLLFDEI+0X6HGR42p2TH
TCHr4A6dd4srKMlxYcZyIxxjNoEX0my/6aM1cvljKG+1Y3VGqePg8MeA8Hz0
oCL+NeBqc/d0zs0p8Djbj+vqy1C8TFVHX272ytzRA7Ewfu8IYZWvSod+PyFw
jhsIP3T85aGP27Otfq4wGT8IrUwPBm/hfMbcV45e/AAXjVFpIlAn9cZKp1DU
yLcbw4gfsC0TrCIIOtFHeB6jmO4rcs0pZHOOlxZQuTVBulEega5Sdy6RJCxg
YusxHW1TfP6glMxDIFMsSFEUY4pQuaXBqGaWS4yTqcOw+gL7ckHMwjvKO2Kk
1GhnrtXNB/Cr2AFQIZs1Atq2AHsTAc1HBJ1ebDAzWQFBRs5iJaA0A8QLuBVA
w4of9f7Mzmrg+IMbfUUwXJlr76fNHgwW9dVCCFka/H0HAJQQiICuNSfBOEr9
ZJRP/c5QPePWBXPsgrlaCDKasPzSJNodOX6dhdMaTpDVOwk/q1BukzbSGRdd
y9/zusdMpJhZ9U/NuDTcXtkKTZCLRCs9cVa+OnhGxW0ReqUBsHHqMF4Yb6x9
lMg16pBTP79YyDmMnEK45jB+z3fQYs4wdVzbXdkLwbWM8bZ5hpA4IWeWEd4l
EuvBJazKbNzSGrSuPBPnLwRCeDK86m1qlIHQOSocn+sU0fn+XfTzebg3+tRN
3gUi9Q62AqenMsj8/7bQC4Yr7SsD/7xLqu4qI0IxnQtPepnxhZAC6NnvM2gc
gDS4iF6JA5mkubla48Vc46lbtZrPlOkyiJP3PNXdJ2ySaftSjFd7scTKAZav
IE5dUaYpMn5SyGn1Lh/c+buid6yosCZoIwbIjPWrrYAcm8z5HqIIWGoKHoDv
vdTgUHpBMKg6257LgU6RvNO/ZAp4wNoGZZEUHzaJbKmLn3njOuXChnHsird6
SRvrMgtikt2KdLbZc6gKIhY8ApXF/kmDgKUCHT7fyovhqpEosPlWPE9TtvLH
Ih5bT5osRMjTZdA92GP2IUaabXLfKUEHxF7EDzOpFe5bKwheeE9CcWsPnXIW
uIsKfHu19IrNn7yjaWGNWACMciAcirvOxIvPx2DY4CokBrdWGr8q6vYkZvfc
pAVIt+7yElZm/ZtAxHyRSzEtAxvg7wt2iMAJdf6t55AlSBVhjq2xHQH+Pj2W
oNzKF9VQDOnHfqDUKeBnCbMqz5/MxztUKTs8cscv82NgfemwrUEljrNlUPhN
4uLHomEvU9jCHK4X75dFilf70ixBy5sWbaC3hw7rQun6YXQ+as3D0hXcQm/N
MDnbjcm3ZmO5ov5myf2wSvkZ9ZXYo9PmYMjlqXnMSj/WvZvldI/SmDwoLh7t
50B4C5D+JL2mA4MEUh7MgQoPFHCAh81YnBuHAyGiCb5LLRFVaxoFM2kUZ6F5
fuvqNS0uBRgWpQ+VPep2rymptUEBdCyqPhpOrpKK7yMP/xNDlpUH6wn0Klhz
UlhVTSF2TxyJlLK7l9XpRfnPHIz0iTGKC5Y74y4Ny3jfIXYM5DgQnClKFBOu
IhPAIomlJsd3lnexiA3uFaY/UyrtU70YiXBtGEUmewDxkHNJfdQy55EWcdKV
d4R0j1E/6HrUmC7vY3h2CfB85dHSbdxQuBnCY9YN4VBTF8CLYGmFtRWM7aBN
ml7xRAyElTiOVASNOYwwr02g6J6mVrNLvrpvUYC4aZNYiz8ACEacy/CDHVCH
LauPsJkmCMKe2wDGaYtGednAfCEI16xFcdUoxx8U+JgBXOUkwzt7sMX+0vdI
HRidlySguffLr36gZnPiENvA74fU98Ea5aBQ0Zn5SE9K/j9GrzZoAcYY+d2b
X83nodFAKaK8Nyoq2cQgvFeqvyg9oCpECBs+N9NzRJdWbm55WXXLZGorR1z3
YrUBNhU8vCW8HF6SwhyR04xWk1ZAdWW6k7SIjy839y3hT3hYJkiXC6pbXTX5
5Uf9/P+kS+0ym/GOnz2nQ1EoB2RcW6PbqXjYR57Hr+U8pLiXKFy6GmY3ar0e
Q7CoZnu+XlJKzTnhtYpVNqEE45pWvV5tKWo5Lr4G2HfZU/9OoGXtbtRJGx6D
RbVAZLLIVATI5TNGeMEHXu1rRcOC71VsfPKnw77CH1DSkR40Uslc5snbbslp
82lSuyFdmkHsvM7vywkrUcBCQuSX4SH7KGn1njKr44E45AjmVN8qZenZFrOO
ARgcrq/64xfF9JDMuGln0t76UNvA0DhVTzwLk61HuZaFlyq9abXZcUiN3aAw
wPR4wYh9lZ5y7h09Meeb53gfeaMV1Cv1Cg7YIQg1wjd0bb+YmSQ1Pw0kiUz9
BU/4X7WmuxnhM2n8OdGAQhUcCkMYqIVvGk9Ld5RHyLVMKwDqI0mRnuLhDybh
BosYSWdB7GPAjlLx3HEy7Wz1hGd8TyJg4Rzj3CImKLI/Ht/9BpETZThPut1u
scekgRs/HhpoFDd9JeudxlEP4+/vTzOdk/WNdFexmLykhT56mzUAGoUlp0nA
suGPQcZpKbUb2B11XlAYVu5J5kcMQ5HVsLThIjde6NbY9+MdI5BmIZm0fV83
TTCaGHg8yi2KHk6zHN+B+3Rx+xJ14yEDY3lMeQhKo9UmSkjPkBf5H+pHwpxF
f9Llyt5dUf5nxxvhojgIeKBUoWvXk4IpxkILAdR+gvjnUO/shb0yGH0M7ECm
GAPEqU+wT311kcFE+xnZpj1XbOmizEdbLxJyPBdTzyTXVQGw8+6OjiFXYDR3
KA+D0tlvu8bKUOwX28IRRp7ekHyXAZBLlBufwMOslxuOate3vyQwHq4NQxjZ
QsgXcE+3s8lFgbhVTAEh85ubOlkgxDfv3p1ua6nLDoZEon/Wlhorb+vK4Fh9
cLfSepgMQzvsy8PpzXUO7S0exIyYGHLOzil4d3VMDCHJpxQqjtAnbB/MgL5a
owdtC2DZZUxb4JWR7rqVmpoJyu1JWyYKLR93M1pyYzbtNO4gDJ/om0eiTzmB
VRTypLw49SV2a7Mrdv8ls0Iprx5vYHNpOwSWFDBRkS8fYMKCLHL7qpa5/uS/
z07SCcyuWkE7/95FWJ+JKd/a4yH3pABc7sdoWSuYrMgg0B5NaIl230JDuszM
gUn/W4lP8ehCATi63d36EY8EPtc2eJf+GQPMDAxQ3766qgr203GnQsZriHvE
aFI96jGZROZvrrItEGRxUmzoyz2E6IkwAmEr51BYhdQyhssqVDcZcUtiSHwA
PrUEYe8w4ldPYjMkOCR9mnQbva457kxTb5vTzeHFokA69KqsAgYhv3k/Jphj
n9EHixZiwVTrKW7RvRYhA7NYb6/WOeKeGdjC9LupCM4Oy8Jq/Vg0n83vZjOK
XWxN7FNg7xqY3fOGGimCvvFCg4qlXHFoSupZNcS48ce0B+ZWh/INffh+JVZH
wopUI9n50/duEevrD99vhX77nVJw+5PzNY27Vc/9DpWc5YAl4jgtN8A7zExp
NQ5c8XYaAplT/5L2JrhqeMKFg5BdvSIFy9okMNkGQVkZg7On7sBa+K2mW5mn
KpWa0rGhNFYG0sh+WeDfYmpTPyAACDIYfbA1mU+BUZnr0VfefZcu7G8WcZkp
IDv6fdxxtiyfxTunoojAugcbfaHRodj8MLBeJMjKHnE5bbh1IrVRtZniVgZu
tFOoeWCRqEx5aN/s5jKKcVkVnF3uhmAt4v5gZJlyGCKHtUtzKJFfMgPD16fO
ggBoRfumKk8vBEfQazyzcNiGW2YT0r/NSXPpygwF3xFA1fvKfETFUyMhXFls
xPCsSOGZkuCf9x3E7jq1o7ZjB8ogsGdekFjHtSqKdmBx1RJaW94qmI8gxkOd
94P23iHstQ2A94+bKS/M6bf0iOCvp+AGP7T+mSrLFrR4Sy7kS4+mYPIQ61ur
S4xtaxFSpt1t62oXq2HY9nIL83QDgnMYFmxvti/j810U6jd5E4kZf2KDD4J3
7Wwz1ll4lKEVUeTCr3f/2r2GO6K0iAhQLfDlzLp/4IsoakU3ZnbSRjLMAT7s
YQS0bEbNHX2zYyO88/fE1HOhcEoMr+Q3bajw5EjL3wPuHk7+K1CHn0xTeXvX
4e9S9zli2OcBwTGhOALXuRQuLU+85Om+vT8OhHqumgOhmz6rPTWZlTzHIeCS
DRh+fqDjF3KQwODvf/8nQX2l2ZLB3Dyx+CNSSztmt5VuwqnG6VNvn93P5yNK
qOcNS8QimH3PRyPbhYfBQXjUDCZ0oM8LPJyTGjRSVnxBo1Iks+SwGEFUVt2o
nt78wTRzPUN1Lmao3viXhqLASM58mkOch3XISGY8+5WLJMolYkBLsh0dimPP
gFqCbXyZ7a7sdibr/jKIn6yyc9vP7J9pt6kOw4qsy9n0g8Tmoa52+KJj3kNu
w3k68JmG6XTucySwjkjd4XtwtweovCIYdyKdQ9KP3hZVPyZyH+ib1tDztNWl
plTDLTny8ZGnMXLloHV/j8HEJnZ1SGq/e5zLAhbO8JBsqBUtVUDYQlSMZWd9
yhIcYyPCmHsLegZoVZXTRGJesjcg98UQnX+PfXQapopN7isCmryy1Ug6Exw7
le4n6MbKZlkzVHnqoxcKYWsjH/d/ADMazER7pp5GUPKGIfbWIKbyKLrhNSX0
UiYL+ELfnW7hFvFfA5iT5WxSv83lrqoJ0NMEW6vDKY7SgmqELzGYR0xs1HeI
xW/rj5RsYuJFPTHgXlS6UyT98yWj6Bf/fZefkdq7zL9swcGB4ytfw3CNddFr
KygjhwdA/77LulfbGZXpHwalJo9laB9nFGhjBOcmntckCwzY5uShayajGSBE
fSwX3ktomyTwOt1Il2t7htzBIoSDHzywoeCHZnkNBxxmDqhTnffSj0ySNmIR
b1FNfnSEnwAN/pzM1y7dp6J+ilAErpsCd//IcLjojmQ0tmOJWDZQbmOEInnx
uJUe+OXtNZrtLvRx5aKfh4OtniJTDPTE8G4IgvrIcu3GsT1d6y1ArN577PFi
s/dLLRJ0+x8KmuerLUNrzxGilXjQhUaaBCF+kEx6bHE56bjveq8X9Mm48mZL
J2YRi0ac97bSG+JpkkQgIm5Rud75clCviuQDWh4aS2HN/qOJCB/uhOdU6tmQ
WfDQTlra/gDjSxauHNX5+grtQQ+9kOQEVS0sGB7Nwh3D69L1Nr7LLnBJqZyH
wUpArnz60lIfABvMioON8HkUKf7D4+/Snpq8Orb4HaP6i3T7ZgMcXEbkL45h
pN6BBRuUfHhBVwNb8TD+P4N+XTzaCASLDPtY3KTFEqWEoI2RcnQVwOuATUyw
t5pncrbO1nASCA/D0EWOp3yclLWI7UxZDznn7bcW1OvwD076m7xeixgoh2JT
wZctld3jRAQyVqs12l+Zt+OjZ/T/no11+deTPtGMX41h8yD/x64VOo1XRmPs
6Ir0hWm4/d2p36voklGr1OzhL0Tn+9BZm3okyzCiT/KiBufnG2fr/YrdiGWm
URTgaPFntiTILOnZEfHySTTZ46I59LAEpwm4b9kZsC+omw5Q0lIinWh2GyPl
GV4Wsb1CL6bjAmwupow9WjsOZV0M3++Qv1j6aHfVb0H92ypyOnhqlmfM0mGg
wbF6FQbJvl3YMcWpVMTgAoRNpZeQxcLMW4JP0DL3DRVlUY7K8WuhSe8moVGS
OL+ttZB8ruHcxmaiMD9KI9TqLQ6iXFrB8gXI8VoVtCVDgD5cGTq+ScAVLBFW
6xzMzzBcEYyMdUX65SPaU3tB2OBIGj3mXxKntrL1kLF3x5mlEd7GlAMV5EV6
bcAKefA/y2t8HyG32868pGABi11gCfCUgypzqCsP1P9w61GaA2kLMH3NtWUM
4o4UjpGZalh+IQx4kOv+M7CXIFGM7Y4YDvowgePmkhOkaYsIIecn4vCw2PhK
FIHwCJsXuADPiOkOBNiAJfwxjacEmh9jI+t/n+1TVsVQ3ykvxn6TUmioq+Nt
jv6i0VTplWiewW5WDUWazLCFfCfxs9qAe75JAeOJJ50debe96CktjOflvJct
BH1RU0xFSfsGskdXobzljyFa1TVAK5oNADICdg8jnGJa0W3EBe+wC16dr6a1
YkxHENucczjc4LcL5mOOl/SNiiMTda69rXM8hKx/tqYaxL78e376R31L7CcH
Pnk9Q/Vl3GrsKRkkfaKB+Tvnzug8RMrf5ORKg7XXADbV//GZxQwTOZkW+laX
4TIktyrhwegpbp03wRyKZfFfZYQ1uWo7NCbh3wpLSrr2xAgacPqZ13GFSUdY
WZeBhTl1vIErqkVGRipWbtCyTQHIEGEq+UGQ9Evyk3hFUGWK83prOnCG+d4Y
gdrgr+yzt8y5HQ2f9iI7Rd/My29tnJeZ6hAVwDkVsaVOC/ypUqey17/vo9mE
7oBNWgaNUhdfTBTjSJHSz8e14maNjUUr1ffcPxyduk7STW5dOwZWJSmIakNu
Onx+/6VWAcV7wMxWZtdyBEacFg4gUjj6OowSdG0wQJDQpRNq6zikpBFc7iNc
LdcLj5ZEjw1r/QgtUHYn18oQDrrNaOAdXqRLSyDeX6U1v28FPgaW6XVg1/l8
KLzuwKt2n3+/O88bQMRe/6V2ByX0MRW8u6X6oymnhH7V6eIU5ClCADaPa/5Y
dwhdzJCbvfIlwJ3WVqorxfGnNqCUegrfVVboQOOkk7pYy1ksqLVxX9OCG1TV
sGJg4Dg2barvMLWCsYRRho8/2Oq3YDkZunMgRNLAb+3TkI2sV6eoxEPEhwiF
b/1rjc8nc73S+HiVTRHjVkVMjRcVCO6vFZp8oF/NPyv2zhxItTAe3MQDzsru
SxnlY1VAelX0dC9ZhQq9OfokdiAc0En+96UnednCaSg1eY9DLRDxd/gGTVTu
gljIjqC5B0BzmGW0kiAJs857N9fy4Yu7wkt4mzo6H8fE2CDPT0weArZcivxp
FuSiwx3Gia05faxCqUe7LNlsNOGP0Lh+qJZPFlsCxis/M+3k5mrO8f0CvdwN
ghgHEKSfM1ztzuavmWYCLRmNzHBM7tXiuXpq072Cm4eEe1PV1HZAW4VKYsrp
JhXXAJgL9rI3h71y0QmYwBqsU8ir1OX1QfgSAjH1IMuNnfrd4KQNxw9EIl59
a2w8ZhLlGsft20JcQHMLggufM6VaKS+baGsysy0+Wi+rAORw7wp5+sJVg4Nz
TfUnJhiVQxufItiHctG8JV+SxM5XjuwQ8SBDA6tmuvfbtu/bW17suMZkEN5J
1/MGckjXMSdFncOLUIICQaj+cD4kUQgn+LGXb93gMqY0k/ox1+3eaKm3NUhd
gQz6dsrDj5yxuZNDBsT3Bs5z7XSpaYGdwIqnqKfcdXOSpnuMdetlcodwgbjs
SLnOaEDgnggeRWus7DA6wJ/nNqZ4yQNQ97iUytuSV+fW6+RNAFIVqLGOWnoY
CPPirYIsPyKjatjBQ249v52Jvgxh05NjBxP+/ZJoiRgPVvKXk6LHSevB9Gmb
XZR9D2oDclyfZYBgklYgaywKnyonFboAGdiamfEtIpdVjNSta4Oyp/8hvhZZ
v9vgcD+jocxaNWssgUPPXSEh0yzN4KfUrqlwkxhtZ07NpZa27D5NgzwKQoAm
OxVspIDHI49yEoRKBCqmvbHcR4CpL0gRhdvAaOfQCsozSCPfYvqFxwD3rhHe
8cqAzq/6VZiu9HbuYXWuM7VwQhfsY3qcad42/UYL5hQztGtKbMaHpGyJwAIu
aZrtCAWyriAenPzpy4D3MEC6XxpGMdwzS6X7tXkis0sp7Ry4xFq/pebD6T4W
St8L53aGtrzX7kaFnF/q9VJEmamz4hxmYOqgZHU4jTaNKQckm1ykIY17PRmJ
K+SmyaKObcK6k5SaVm+2DFfMS+r7bF/o2cwSnJir+jJVziTTEwHaaDOtGXty
3GUgJeSMIpB3y3bQxO16MC5orVoxf9EW013LKQELbuV3h4Sr32KX9x7pCr2u
42d0UdSol+47gjv8735oFBwsRbvKUA2j4TlEWsuW9yyDU5+DfGUv/dGp2fEg
Ppi/wgXw3BsfP98JF9gAGkPpwssxhBZHlqSOnOi4VjLffE4DWSn/O+GTXQFh
sWUmsfpodO6ivTKdZxh5unMAOK/ZwlT6ITybzkD+VE/FGlsagjTgxtqP4VjR
V6TSDrfWCBn1aEJ8ac/oDFqgo0YzrIe9yByC8YL1jsm5cStb7bWQ2nQ1e3P/
Gd2MxX+L8qc4f3ZwM/Vk4Arg7cd4s+4Ym0JcvMZe7jVwJSbkeuuRb8tFCB3Z
Fv/1Wv6gfWM+Y1V34mnMs1dNUGI/YPOdD4y3v0BCzDMHS8TDA65xsnBY16Q8
Q92h1c3e7R2n4BpSzWKChElEbjMpqdUOza7qsty0xdiCIngiygrZLb+nN4ly
yVvZU2cr3HKJkvqDjovKxHQgzHXDk1K9QCmCP5T8mIGosCc2lImMjcBNL0D5
LYJ+4v2uuHQ3D5uysnJ/2BTTLRpEH6n6EstCgDSpg7Nl4AI4HR3mzKhQaHJT
XpvB554AAOUD6tHCS806cIFpEk6WNEuqZCfutVr0h42czUluzMEnt3A35GNp
NxMrPBEBFwVkSy4d7KK/aUN9hGUw0TO6sSIRleSnLdNWEzfrrniwFimlNtEZ
gDz09HPUS5nPIq2HX4ruIRIV92K4xMFJAjlkFpWQhMZ/ZBj98j9FZ3LuvWID
Ajg23rEh1t8nEdTRjlEkqISwqF50ivBJWi52aPJe1IsflUyTjvzN3aCn8TQW
nLfnqvcVwmKwLoiF3YDhrSr2zx8hKrYAFgHvfnO5NQZ/L0coiI5MipyMT4CR
vlQD2jsZ7iGgmLyv3Eh0Kes1lTQ5X41svlkX10I5wOla6Qek6A5nLqcgysqJ
lzfOJTzJ1cQNzQuXHQPxPql2VplzoMtgzumzJX9qI/XqfY2AKEMYQC3dbySr
O0OXdInpg9kwhHj5NRvq8EFZwBEhRw1X9lATqxJUudd4hluvDdpUCFIcs8RG
FITFcry/2Js1KkHu4xi983HnzyPiUH1cJ+627iqov/7IWvypFN4uya7wTHg4
n5FvxE6yDtagnMvNV4yzGhrskYduzeSoyGTQ74gJ7LTXf/wUB0c7B3yjcRTc
NbI0I/rvOM5jeovMKTjkk2k1DqigBtAGCh9xHd/KT80NHBXApC+uKJeP0sZ2
sYMpSqMkUi+s0aAilndNanmBnLglN81HXFFrzcfsILz3ss5poeBmIajJU6t9
YwY4UCEh50FvFWwPNlCrh0N/1UWpoaz7SybAy7bNQwxunsqn41cZyDXf9x9X
+qP/P/9+00e4xuOmEv16DrGsaa948hNCLNyVFmYvhHFOIQ0AwFGE6xDGTFPv
RFiSzmw3Bc5gR4fYdelPJA6cOxwJbYQnDrQJQQrxvapFzpIe31TUUz8AmJ7r
PIBEryOpyBG7gqJ9nKcqicInv95jzeMpLj89i2cyFMtWWZ2HLl7p/vRwLAl4
LJ6jMRzGFr/YOG0vvJqSwq0AJ3b1j50Jx2fOReccvn5mBYmXzbP5x718mkX3
X5c7a0wImEJ2cWzzqebqHj3ShOL6MP43kroEth12SnKBwfUvyyEWNxDFOrKN
xUPOdNZ1hwbsuVwM7orfo3WgGqJ0i4qThxULDdXNCwrdLDo7/NKYIVQ3nw1m
bqlkhYNj9UKZ95xqQrw20gvgIANZgZ8a4TdnE1WrOjx8rfA2DfUPIQf+gON/
90X2Tdbagax2p+r0Dg4wC1pI7Ac4WbEOgR7J4lJ3WulcoXK4IzEanjLCzayj
cBHpJV9Ax4+sS0dBac3jPwuj3mWa92F2Hchs/Dmmg/KsVLaLVqlei8Am2hSv
c898NIVeWfaGqPE2ev12l2Ztg36oB8IePWAqeC4n5+nGo3pMMfcWBi1CaYKT
kurHfQpE7/Ps/vY9ZiQpWFNkEmTSSYUqGM/+pc7iSzAjoAr60yMKQVo+NTju
KlaUWjLakBvaV1YKFKRwWdC1GeqFzdk6W0yWh//cYkdWIHKsh88Zcd7BwWTl
5M1CNFhgjACXWSkTdu6DLMPF+ttJTxy3xWgb++qstJcpwcT4jWW6yIIUHnzB
0OF8u03HQa6hMLAB4QdPAlv1ISzgEFbYBx7G1bTJX6pqXt3D6HU+d2+al/Qh
WqKE+PVYauRqz/aP2RvSwhtI/COp+2Bv67bac9JLQdtqCNEcOPdl9FjY2SCW
E2pKt/mHOIBFVVfGRtu7EE1zbI4lNId2eomxQV2vFBMupNhYHRpE4UKeTAm4
ntHHviHBCdmCZWeVgBkUaT+CoF8YTzBbtFczMJfbqucmxUerqaiTcAhrRNxf
w5m0A+pXB8iwm6AWmGmU6p6UhZgAsyTp7iyLztAQyAdfreVks6yyF1NFNk8s
nBdzlDMN1qrzcgBVJ2VQhgliBrqMv4ur0n/ovoBsNHbZVXRj6LlviX6bfGhb
o+aT7PqsS54Q4BHpB5iSGpU0CE0GskdynykT00Ckbrm0B9kWnUCvOR1UOAXS
fZR/YpK76L672J6mw2ylkNOBLjcvh6xbxQbsTb1rs2dkdMKY5v367Jppj+73
fAgSzitbh03UTt61RS4j5LcmtPIVbN/oLQ81kGuW6xui5LilcaFrvFAcUkgl
FLLFIV03i2HDStPG6sARD8cNqp8/JHpehMA7+aK5fj4behHhushHZV5b9V4F
AHRTi3TqeceNQo0kljr0Tr2apC3KhjdzlWmeXaBCuRjX8qslERwsbzA5+2Qe
gUbmwpYQZ1IxsCgWRqKbXIPfiWotWupADm/vMYJC4EZ4mZUX/0FTaieewJZW
/BgsrWOiVdDDBbiN3JNGlx1xzWyUTgqEE1FL4XtX/Xm6wbz6pKNm/AaGsrKy
dT8Z+lGzBy75+0PryeM481ePcZ5lumcOibG6ORdlKNnqcO9bOACWWY957hpf
FofGyl9WSanaien2IG8yg5Q19j8Ki4kNYzsNCekTnP5JKynqRG+d01CIwVbb
ZFr30v9fbqB1RzLaLnJ3pYze7OO0/NZK9mox1yYwNV3FIWvdpfF/GYcx1jb4
gPkcQ4sJKQVDYxmSFygZry4GZnhkonPp8w00Oqjg68egV4keO4wZtg8KLUMR
XCoy3TDiJIbExWDnvWPZHsBKUZSPaQ+jHo31yRKNMHVdEFuHRzkjXDIEiJDN
8EVmjrnycFalhoJGhcZ+PKT59JQ4PM0IzfOQqCSSWVGm2qmzdZaxh/+ukpN2
xn4BdqY4oknOdqeoXWesDU6snAwAo5HI3HZVbqd0oOU+V7L6rbw8DRmSBB2F
hB+FGcZR+s4NlGA5hg/l33+JicvKJvIXVIw2y0umoQC0a9EVDlQzTLZ0A2sG
DlN/LQV/REtM4IdrUPre3oYq1uIgYKHdcgx56unlHBg2vSlAAY9LvaTlQCvv
s3VDldfYXTfnB2QYgneqFlDdWbrlCYTBaoPJes69cCoxGdVbuxwnv58dbv93
r5/J3oN/1JfuLJM5XJdFLgfJ0GXRn9VLY/WPzv9d3ha88/GxSNDg2fv7Caju
VMTS2CBHWyMsRaZXQgDT2t41pX6Ie8rp0o0Vs53wwHoTKYWQpt1yCgKSMRE9
hCIPbwvmgKfj7kR9+EdWYhVTzKeoCH6k/P23muQzqyp2HLqW0h6AFK3mpvuC
wxLdF/WqbjIYN+Zoss5+ybMR7q+QbOY+YmHBKOFIgqXAhIwuMgL6/H0ch/S3
MGowncyD3DC21ngg3Lf3xytvbXUehYS+FH4qQVyzFmuLcuQZ3/yXQqhTi1UV
9lIkWHlLCiEvMocw3nbVrhpdCCuqgqJkSFbJArmIHVn+X/ViRwz8TdIabhyV
Bw3IKq2NmSwuIK7wvua6PcLQvr92INZbLsvbB1YFzFeXntVHX8gngnYPDEZ7
Xg/4lGecUXEUNlwVs2gTfV4e/7BK98K5+iYmO5+rNjp3++CAYQYCgcdxUX2Z
u7l7jtoiWSrulOESYq6q3iUG0VN66qfuqnc9gwSADAT8myPkeYY/J/YWfGC6
WF2f2Wi1wI3uU0qGjh75fCFuY3tU8UuLIB/OSZYAjI2yDtS7ze6n9VXRX6i2
ugyEgZ/hSAKtFiZRxJmwILz2xpJfwLHl99ropaUkIovcYtZfA6gCApXuMjY3
vI1byxlOIXM7AT3Vli55lErwZSs03jAX1Ov/BxVym8ESgnsrdgb8yOTA29qR
J2t41XdCjphKJud8k3byxKd5kTHua7x81rR1mgXWHSoiqe4WSt4iWQCfKv6i
j7rv+EL5qoNTczt1v3MMPThB++DQuDz0K8mCA2ktb8N8AsQl8soL58pgvxew
XBKdiW3t2ru1PwsvTNpy7cQCSqAgS5v0u+uMbM9aeGdI7zl7eC8/3oS9+b4/
mLErLuqWbasfGTqN/KpqohXleFV7H1Be5DwYT+CcBt5Ytzuc+b9g7tSnSEg6
PJCBzXD6uvNl/PJU3Ao68r3sfwxZPUSuGXbWLJAEJqrFeBsRJT9dJm6hfp/5
6ldi9tiynqTd1yl7O2rjGZLNOndXIwNd6KAF7T0srKGEl3vaiY7r+yWZwlmv
9t6j1BUd8NRRK4yQyPBaluUSD46WVDAEnD4jRib//kgbod1G+XO//EpzyBzF
67/P8n2RBE8citXjYTJAyS/01rudgehEwIItW3lItXr6SSUWxORyeHe+WBr5
fswzlsFSnrbwNFjTCZR17/sDP4vS9SyjBai3CtdTEkU7w8WSHDGAd7F0UxaD
ucRAAn4Mj6BmL2IFmXyJbciqjb+Xb4rxyQZ4vXw9enWgVWNFvfFWrygy25M5
KrptUZw5FDCdATP4nImVw8pv5jYyEV7Vl46k1UlSq8o8VahzWbhTArrtD6ga
9W3PCnCRo+bDLDfsktLVoyXmtDUoCm9LI8OqY082vTCK2f/OHXFbNcOCWgof
O73MSRdG/PFhjVWJmzDZ1yew/l+KkJGfSDWXUT6BNVtbSujD2jFGK/O6gOkD
Cyk4aoUe+nu2fSxSUmyfaT0O7OttQW696e63u6Rvd0pbupUEruJVu3BVa2eL
PKlrYhGxkACXgQXkrKsJ4PSrt0CSYanhz9vxBjX0pjXaU+oCt7iJJPyLunmZ
M1NkqkaIyzTHuuAyHUSSmhsTefCklOgZGEW55cCkY3hdQuG0hJn0SYryKt3S
K6tcDMdeDfk48FhOQ7VTxxMhOHi9KjhQiCbk6doAL0CEYikvwx+gHdRgKw4Z
L0fCcKjL045CYaVSJAMDLeCOtpNOhZURRgtf7cUOYS4EbE6W5gTinM5u4DLO
h+obSQcZYcsShFPV+k4Do9AIKnvr+gD6XJunvSBVaT4Q8Lwn57WzV2J/0qiS
1FhZc3Lg74q/1GT55Dl3ailYa7ZPIpM3FPxju03P23cNyP0BRm1xihjboXgg
Ve1GmocB0tYlFboGSY/5aNEB0+PGilgCPiL0Cf0IpsvfGHXKTWTSAoalOKG9
u5t8dbpyx+1Gkb+q32+//G729Fab9lRU/X0t1jL0qY3zG+F4RMlzoiDtprtB
itZDCNRHjn52k/23nkUvW5YG1kY0JqiLwNn74VJKM+H7MtsxR75e4jL2coYs
VSIdnpFjRX+fO7ppx0jjLiaj/zJUwdc5JyeZY/0Q0GZS6h/DUc03op4q6GwH
RWANjOgsDb9BjssLjMfq6Phgy0ObL8FDo6r4OVFJbAS//lkmmAcL5wiXIbhv
XdbySNSAYwgWzukA2u854pktYJXw5WtVTjoK2vZfnRRvJWQLtHESeo3NCR89
PBDKzW0t3hhxB4AIWFDn1IkNomhF6dDeMuckDu8bZ0cVgeCkVLkpMRrpVdrS
8Otl3HG79XUb2Oo40KDEu0KLN1w5u91BjYtfyCoLb7GX0Nl6G2j/iTIhZR95
8ydq+cEF98qFQDKJBqWqe+eCBeoiAILB7s4UaFz/jR9XJ/UKYzQfEpNTiWSN
dp8gu16xCSEMM6VOfmjMgvINb/rROtEs5PZlxTzgkDILR0QPUL13CmCgQ8hA
srTB5QxnCQF+H2dyk9If09dTgUtErtpSh0CCbz5QiWDayEC/8RJ4UK9XlgK/
sJ6eTzTULhGIQlGjEnjOQVxjGl2GW0mWVHUxGMQlsW8tv9bk9AVhxh7vcYqn
cT5ZJiFLUNk55xpWbf2Z17xnrPxk8m3RUgHoYY3inlsH+/Z0+1CtZtxQewM+
rw4AC6f6sjNh73jlaMATP0WghL6X68XItpbBEyFRcrL9ewRItavqafQ4RgbK
GbW16hDlcTxi21xQT8VbUA8O/Ey6uTMQwfw8NrvoNtRA1Cltfqh/3W8p/mnU
xPIwSQpayDOXCxlciMBMpu0BBYL/i9NzlOTqqMMrzXH0YN0C8yyQY4c1MZii
rCneD4UCJUnF7G0hnu/vUbHkIQrKLXWMFRjDrB1FDT+70rTBSmdnUZXhGJz0
txqgYvFtI32D51K1EfgYOakmgoE+lFOVSrrDx7SXyv17dolbURO+zdgt06Dy
VEJSbyFtEmCMgVk/Jd2TzfaZzj2Z1GS90DrqUPm25Uy6V4g+MZnJQR87kpXq
1onGaLR0xip0vPUpb2+kbCoX5yLszXIx8K3O9mwTf7s+rV2RLNa4VCgb5Y2f
ONysTx7bVCcFLtCGbEZOtmgpfwzDkhUotVo4Ybqq9fccplVx/QvwMkM5icS+
HqHm+7psYq8e69VYabW2xwYdCW8qj7lKiW3vB4fhHBw9ZnWYmku5va/dxyYt
bt6KFHHCgbI19VOL2lrUkMAPMv449u5Xbn4+dhcT8ITwwLSHZS8qHLMXQNPK
425c+5vle5ajm+1PoOCgsl+JV1xvh/4VaXE//dDq6M0IKEpttrDK0uQiH6lo
LXXy90k+7wzUwHVuwpol5AnYbVvHENIxxMw13R5A9pheeb/0PtMBknZxp0sy
BgruvdfF13CV+EQiub6kAlOjmx431r4KBhpZyJe8t3lYR48kituRO33ikJtz
uMGxBHH7pFLkpI1R15032zS4P46OgcjZ97pJ6XGTBN8izLBg2dmtRr+8BUMQ
iVhnBu3f/Y3qHg6jWWs4rwSdT9afmmaMRqpPJxmd35yk6ebA4fHLchUHuhy6
njh7RqstlcyxojVJVPya0UR/13IQp6rqJNiVNtq9RgYJ6ChYHhJqFg4ctLaM
ZP8Bz6+Tefg8NlkM1b/mZFZMT8rrwoE1ASUPrHgfyFzApdvW2Cy9kkIksfj8
XZuUZHMKOquOrr3vJli9P3bak2jzGDfE7bf4/7OPbuKoAhmIVMukjQ1zGkNO
/KX/CzBNMtwkZTUeouRZkj0XysNjKEDE0S5inY/tVKoTxsUdG5OsRGlAy2bj
rGxEDsqTeMNiYNrlE25uDxq+rxH+scNMI8dRNV47+73FDqwVCD+Aj+txsr+F
gWAblf2sqvXOfGDfo6Nd/ZqxSMs5ObS5RaGZgO5YkkdvvUJn0tCmgw+veR+T
eTRT3i84EPrB6hqaj7yHj9H6RiHrm4mhw/s5bNB84GQvQ5jNNmOARxflKzyz
Lpj/bmEdoCPvQaJ1ZdEEpxIEING+cwuzjzju5MD/0Uv2q9DfCNQ4eF5UCBXU
zSizNlJ6uKmx1jN715wkoaUG2ObLSlyVoc8McYtZAsJ2K7zkffR8+DCeVbFz
fAHSbRl2lOFdGbnOhwYepsPZUdv5eNYOSQRX73DZlU2LSO1tb+syO64TmLae
T+7hLjm9wAXC1LIXFMKIF+u5lSf3YAQOMJghqN/PExdq9lo4w6lG/Oa1D3Zs
Dx377pEnxRgIpYBZWq9IGHtwLPiHEfAHMCoZhXBHsrnSH5/5Fapr5ooPqrIy
SYbzgZyuFQ4XHsQNBcBkyhVfL1HUN69WZ8cD/s1Qw18VyIBT0KZaSaUddKhs
griVNgYGX3vgFlEdwpwHVmrP6EEom3VFwCEdlm38SHZPO7AvN815unjZtHde
h/GhiNcSl29UvBh/B/x9Z0tr5CfACymF6wI6iSJc9TAVQzwR7yNhvhc90LvN
nGMslNky6U3Rvw97uNvSzpRYKqhwDkKpRmVHlyPjzIeKQhcdwI1glVLbxYs+
1h/I8buIeCy4WDKdEJC/vPKmtKPlP5dFoP7YTn9FBz6OOCViVmmO03XEyKiR
CdK59H84EED6Qzj2AvBvDwYG5VV6paar9lk9bDINcjl3pyeZaQP8hZ2GfK5F
U9m/jqGclpN4UpTE7GusGjyzqyznkQyde2bQjb+8hUR2pLRLq3Y5t85nTVy3
nSM41M2s2WPyNJWhamfUuJTiOhGUjXHF0+h4kPwveFPznaJETNJM6hsi2Gsr
rBh5pjK2b9xYMQczz67/ZXP1Z/MirVAqToa4ByfKWLf+KvOF5YPyWdMpLOKW
FXQ0Q/2/o6XIi7tqW+8Gf9ftXkaUnTvuFEoD6/pcI2VuWiCVG5UVQtCsS+s7
A/ghr6CpbRv7qEuJkB386ZnOnfyM9rEP5+1gHZql+P0OIotJz8gLcQYqLcsb
y6iJJcWQIRDRpazP8lnyh5fqSHjupb47/YMe3r/ZEao0UOcl7UF3idIz8WhA
LKkFRNRmVJegmg23U+FKZx4TDr0OoAjpeWWP5Nxl+YlNvqR7ppbVdiPnzqss
yWCukNWn59xqCBvAAv7PYQchoiylsjHcOLCkDrKR7r3ccw394ADQYr3L8bes
WG4bABV7JNHcCynPmIKO1SYRG+PGfI8MfZAI6K7y3Y6L7wemXj0tRISyHZdP
Xm3UmJ8BgM2ekqMRjbf/1Lzk0iq82v7rL/N4PC/R/urrm32fyWdzNsyIm2r9
BvOFa+adDJbIZl3coYWQn1420ixmr/T/Duu2nh40Q78oknhe593t6xn5KNoN
e1quebkNzva7ohzSKD5UuULP6hPFP3Ac3T/XxAnTONGYTPoPmr0wFJDM9t00
Pf0wPDBYKEymkHVSTIVsWL8TMVAz3g8nyTY5dWtmFX4S6kaXIroF/JiZ/qOE
9R3PJ9RTRjBBLpaJiL7+HT6UujQ9Sw996552HcPi97zObFE2WRvwArk5i2Jz
GqSxpcGp/SIDmsLQ0R4+RxJeC5N57S4TV5uETXcTf2G6m3lcdag8omOuekg2
Fs/y6wtLYybbRD3v+LiME9OkugYz2lG4btFUIc30DrB/bTO7tEwOzIPZolsP
GirH8xmNn53ZJg0/A3J9ySwZ+cwsrLO6Bki/bPttjTmsDN9JL5B7Pd1uo+Ok
hSAc7a3cspMFMeBummy2PAbSp0gPlpy3zrGbnTpnCMiud5HQacpUx+kLnmOk
pFKLsHTDN/NBCJREMaWRwTezVv76XpzFaGzD1Mp/CZLNaC/8YnmUXDknnNlA
2nffkOYcJF0qaOBPjle04EFJYW0muXnuMujO1iC0hziRNqLvveZ5XG0we9MR
m5tQyX5cYc3FZJj2dE53xnYRKQdJCkajTwEOGN4U5f1Cz+BiZ61B67c9Pnto
TQsJpuMSZfywvFFP6T3R+NciKyf60kVI5le4MJRO2ZOHyd6pOWa6oM67AZxk
XA0JDqN5D8tL1g7BzcLCbOleuI1YmcLNG0XTNnHqV074iLLCAptLPS8gK0S/
xQOB96RHULIt7zG7iWrcyARS1JeHXfrj7YI+Ue+U52uHyTJFQBFy+7LVcMU2
2cpMRRvB5v7PMJ58ESLNpquvhRVd0sdTph1mnwfmf26fEMcId+y7FdWqy4/V
NBBA8Hcx52f+ysDJy9uYB7yKb8k5N9lMnhPlLm6xg6kNGwJJ1FYMY0yiEXtv
UCvzkx4eAv4pBrV86pY+vQJjzTuK16ixGRAbQBcXF+7z/0r+SSehax3gDZ94
ptNK3+4SgNZ9BRC4ns5PovsXiy2h1ZWQINTuCmTjBOritQ8YKeC2jDmML9h0
iW79Orw7/dI9yym+oqTsUJQoRpR+fYeZVp92BnN9C80AVY8Dc92yj3s2VDem
fJVBrYZCfX7xGgD+E0ANoo3C2VUXjNwuWs/sYYRhf/7Jlb/cf37U9q5U86Bx
ivEf5DhdSMZvYRqcQrE+xn7fjDyDfXBtA12tNkrgzy3sROGYOvyXC9m+MfBU
1m5JZYH3dIhIBqFaloAnKkNatwALodk/y129ZyMpUjhhsOsphf7IHHi3+uQK
KOyTA23L6yaY4Do05coebkNOOqOwq3ZruM/2003UevcSoVf2dkKlvNQBPF9U
bJ9DVceTlLUTyKpsQGKZ4dt8V9sNgHmohqOh57h+6GyBSW1z5DGepeT7skuM
V81gV7e4qjyqug7ab3eMess3cqVNSnb2DKanVWi65NQHI4eTYP4pRX5rBxTX
7lQHch7cyeIJyTaL+YYKBIcXHHxpm+cGptJbBi4HQJ29DnmgJoELSwZXkFwy
+f3sjUIitiwK0NR9xNzuNkNqLTYb2Cxd7hA5InVYKXXMpUB28oQBG7t3H/Gk
1dK84QdafqLHWRTWUWki4gBrRblg+13QBD8yQiAv5MyK+prk2TjywjswBGaz
rjQQCuSSgeejiL5wp1KuQnIl9uKDkK9+cA+906j3GCSQ2RlvZppT8JkKpA7k
6e9C00AzjybiILBObVATc8FCI3yyN0dd7Hs6H06H3Z8aWfR4JR2+Z7oqVpEA
V2DPc904DYxvzQfRJ2S4IR9ovOPbtrIRWbMQ3HvDO4iqEJ76P8V6dt343zPd
hC7xnaiZN4geNoUdz41uy6R4RnEvIIrTkosdyyra4dh5OiNN4P3UgmTH8nKR
9aOIrVlzTObd8WkvGlhsRnvbyvxY3469oTNu4Q/BNgGDupqaJeqbYNUrT10B
uvajQs5ExupQXUl5vFuTl9ozkHY2HkVIDi+KJ5ARAo2szuPFy00I+2Tw6IrT
nVaeVWB843bPOM4Uy1OXXieIcbStV1Zblk/3C4LA8JUZfC6d/EaU4Mr1fk4o
EFXXCor9EavSyx8/9yOQ+PzFaGi+S5DK5s16gzyJ/dIRp02jl5c0OKoQjOGi
dc+XBCbqFJKKWme6ZxPrkSIdKnL0QM/dtTa6zQh3ukoLFOaX9Xu/UtdGAq2M
u1s8IdBF4U8s8GrRbA5p9n5mjDMJ9U7xB7UFamzEWHVD6cSVOydi4xoktDE8
/W0E04909B37CJqYSB1M1A+FV7qucNdhsGPrW7iWTx/b3uUXkpcMIYv0Brs3
3fmIsOv02Iyyv7wnIxeuF6+15F5BMJYdvDt4xJMzXS/iecd78d2Jr4bQrxgv
H9tbGeO4S9jnbtw6CsWuRIPDkITxx2QcJ8+nY1fUtXpsKdyd6VIgiTiRA9nc
g1TAx6BmUV4MlXGOvW70aW4rdGX2uQL7ixRAU/dwnZwHEKKz/gwC97VrBmbY
RldU6GYwb5HH0FZQO0vkbw2TeY7UHAqvhD7JW2eZ8UxiP+HASFAfh9vvkfmP
4zqYxM6outu9aJKqDtTwUnivXTsbYrJV8vJjhKUXooYMfM2R5FvjGCf23s8I
26tNNKceIPgCiSaQRNi5CwDbEar1UL9qj80ckKQFACpiQd83/GfZ3HGn9Dto
zPYmmVk7I3zReioQKiaRF93lnETvpjOJifdUJ++XSLBV5MOas39mNyNUAX1r
jCdZFFF7+1aWHWHxpRu4oGhEA5vSjBiH1kEETiXacxNfTjo4XicmLinglUto
4iyBo+cKEZia2Ty9a1Y2dFEK2MQD3nxW0B8Na3vUzmMD+T5tjT+pcWEucf2r
hrLaqAsbSlkbHnX6day+8NfmvdSXySMm1gBGNzJoCci+jsGUGWtI1y6Fj+yL
q8akk1ZFFN9xMwusP41cLAssYcGACiEKKOrj6Dnc0VVeRi8MQcBWO6mEtTLU
9RN1XfeshG/tGf3eaMeh8VloRgsieuTBv6OzwPQ2sZ5IFrgTv6ukHBskU9Oo
I9MwNS45lws/SQSW+Gsg/hXDF0eNyIO4AIzZr4S49rHinStU3d2zcW6BJHSg
VbJH0W0ocOKoMQTcg2GPBMBCctAY4ZADyDaWlROU/YXivzM0o6DoGQc/a1cd
a4Tn0aKZ7inVAy2Gv9nJWAYbMGZHF91evsxk1f0ZApg8aAN643MA0cWfsQKH
qafnkPxKDUpJHkMDhGjO1WJwh433oApdbSsvMjgE0TMlHhayq99WBammpecW
hBCJVRJGqH+WS/143FvuHNNrx4dE7J9WtKTY4gy9NYTLaDuslaAj33jNlLnZ
VjENPm24MxnamzCtAmuq30o98mdnt6hG8GCmoUSyJBz8NbNxs9wAC8fwQLWm
zaTPiK/FWma1gNF4gQ2x4iLvZE/TzjvWHZYlPZe0GOc/gkypfdrwA427JU6+
yL3pN57iHYJcmTAFoS62gffmKWeoj3PXKU+abEXj6XIJgFRZYF7TmaOXtkaE
+gVxn8n/DmTMhrOcikCRCwgNMVCrHjDHMkCOL7q+i9ZEdogIB2L6bgl3ed6p
zVhytsapc1YeLRA/uoAlWpzk/pFT6nyeWbkIikmfCgTVS15ycEePs6p/6BZz
I/4Gyh1d0jQkkA8Q/vRRc/MfVGDFvyBZ6fscEt37xTjf65x7UOllYbIFc5Vo
pzexdwPB7uIRpSWuKkadJVDKAKDXkMdKs5YaYRIBk+NXrKdVG3R8ebIx8OxX
XR5alztgoHxgpNhO0NSPF2JbA3/In2Q5JqGCw5Ug83huW+6+sSV4ZTYmi/8F
FGx+ZabtgcN04z4PiYJn6tUhOu9ty/xqxBpKuobigosNUEYsvZtddL+E4uuR
IB50jnkw2yHNVyr2VpjLhsoFDX1nre6adYjQiLchjHjMy+wBIUnQj48sWPV7
pnw0fH/Yrco/CPfUEo7Mtu82B/jxdqAcXsBvCyHhuz/fQbaPKLAHpd/pKaQ0
aoeN9fEIle/jEhQvYJ3gFeco8zLSpvn8/yZfpFq9M28UuupAbx8+vgyvl45h
PO2dJKeZyHr6y9B4ra0qlsE3f7aLMvc8wvKUr5nqcXKNahS1lG0Z0+/a7CZH
nMOikrPj25umSTQuY43AbTshHl2vWJDg4HGie/A9MUUb6dYnqiHH27/9N80x
V7KgoyCMnm9pa0Q+z3dyeUEG/GRMrQbzlpACfRTyTKe3smUdjVWSfyryNZ8F
OCzniwtZu4ihYaS5NMp0YV+DusOpV4TeoVISMXtoQ/YOl8hDHsnAFIInRsKa
o73XoIXuO4fyIA/xvhJFxj70vA+n8848CVCjucUIJM2LEciS7kH+Zi1DLprz
ECwmpBZV0lZ07j0WfcnOH/vmjUqJb+LOCcwapVf9/w8jGDdTc5d/Hb/Tz/Mf
3SLH5otH3BxdG2PlKhx0wxhOgv7Env9/gjHDlBx5DE6FBKCGXVxNNBNqNaB5
idYOu+O3uIotZOaxJcEEyc5xQCn5DEkkJap3/ObypyfjIeQW3au6uJUXUFhY
aPIs4hl2X/rC3BUdGlgIF2wwwkhO3cwtrH9Emo8XYpECJPIqBikLnRCWbKQF
lfSZ1eQUhUg82RO0blY7PHwMNTkyUiMbvYS4SoUlzlTCnIloQ36gNj3Do5GG
mn0jSUPlvXUY0zWt66LOn4MYDLOvAUs/QJWJxsRVTOKaxglOVZGa28uCj5L8
T5y5MdmoUV9jSmli/kFYrfGSAkQ2UbGvh5Xl/TI+DLDoAtngWJn4bwrSHXv4
BU8lWIL3EG9NO3U18sCotP2lp7buw2IKVa0D2RXg2UHMJ+Xi6y5ybmsPE6JF
CckRiPMt3KC3LzNNivkPRLNDVqXtgAe5joJPHoekKnByHHkwm7N+rZIASK+8
LO4DFx18mV3h+zvkQzMb4dEsqHX2rGipofkI8/0MeyXUanFKNiehhTVLBzKs
VkN4rHVG0Ie+33qK7+p3gydLrEXxI4zbrNUpIaq9QrjA3dILjYT8q3XZrhCh
YcyCeQQ7hktwXUy9/vRHob0rwkjv/SiNfsCPpNC+FReyPRSkzm2WdHLeDo7U
QU0I+PE5FbpVmzmf3bUXiFw5XuC3efM7mWFxi2nwOl7UvOIPgQU6K+KjXmXw
JYLaZAkNdmq+U6i50J6hgEzDtzwJEfEA+lLmhdbyHvL39kBK1avXAHLniT7p
B8d7Th/xl1x5K7UnlLiEjsu7k+8Ist4iB4F3Mc5W5xItEVMNXr9D4HvmEXj5
VjwFlL1hyujhEv+ewi/SLS7a2jXyE3l2IU9hlGe/EfSpJQjreVRgrUK0+n5t
VFXzRFJVNGTTJ8lDP7oZacYrNE02yaUhJ4G3LxagfoMA7uwQaAc7S3Ki/3Jm
ge/WiJ3drT1AEfm4V9tm/Nx9JQZPd49S96x8SHt+BKRGvG8ToNK320VcTmIt
JMPin4HC2dENC47BCIhUj5pwJ1NU/6ywdGe098UHSXYtAobNZOBmNUvJvTab
pFo5hmSeWXBzNEcZaHA3rf1o2YpMKUDfKr8K8Uy1XtVd1evYZ1cciiKC/ZNU
iGGIJmlzYOmkk7WawvHj52OZcfqVYVI7vKQv2qUmmwTDW66YP/f5PysqhOVF
KPQc3EYSXKdRblbslwrTSKYPZicCe5ZC7C9mjqn0wDe9vBoQX6Yp8w7lowRq
1LsRzLPbMhnuNc3gymOqDIwWPWr2HEhHL4kF2cSskH/UAf9VmtCr7wZ0urnC
Axndk8FlYtbs+wXaVpADrH0UuGV1CRzWwBuWbHANpnqIh+n6SH1aTVVwTlCp
tinBlCDCMbEkgPBwlCYgrj4ObHoD4spNh06mYoPorZaAfyV4O+usg6kS3Jkj
TGg4+yZnarp+mWEh3KWv5TrnPklEL6lKo2MTHQS7JHQ1ATtZ0m7NYrUQCfT7
TYjQlWI1IPNbsVNOS9OnJ5bBXCNO4PDnBlSo+NxGDqqsgNsqUI8ItPt4Cqb8
yyx7qC9VB+u0vP5MYUqDDuWCu+TqW24JQZWzgp/le3kYBImODsgSggAqOFct
XgNwXbXSOD+T4W81ltETg96c6JyaEDJx0eTaCDyPKggKwGqHUH0FHMeW79Hn
syEPK3zL0/4E+gH8XUoavndNMU3MjuP7IcnJWVSav6bFolAt7uY5vzsEW/5X
oaaYKmKzbHt111VP9NcpOPjybq1P3amsM4thgCTXxVqpATM4/18L+nfq3rdU
hsRRVExBTL/CcN6Yc7mgWP/jgskX4qUr95x2pdDqGHprkMcP/rjCiVt/0AZo
RfX2r+Ogveklq3HwmC2BLHSgEpVO93RvOslVxWb3YO8j5SFJhKBjP1UWQYwM
DBFyCXMTLI+WETL2hLnK2B75F/IrNgYreNKDyHJQmeKbQGjGNFCQKk5xssge
KqvWHfH9FZoMRWH6vq5EM+Xf1IXFXtD5FX8FnERze0q7uLGKFZp1RPAcLZUR
fAPrYGedDCpjIo8+WdrDq9tutCs2bbBOAMadCVBo/kTXoXjNEG3dCmzv3xX7
UbFjF8RsUhM+JLTHhQbwQ7nPsfV2vKopJKe53H783zzDuy0FtwxrNztqEGJn
cCsbUQ1eZPeHMXuym8P7Mo31vcZ0Exo4BZ54kJjTdw9kwmm07/Zz2f6N1VLZ
udtsGvn3xUBNsas/b2JlHotCSFnmc7i/TX+UOSobjGz3y/4Lzc3RJW6aWPu9
0jJsTghFCadReFV7d3Qr8/eQbZ3k3JjGIt2812Bkivc+8Wp0qFESGMgAlDsI
58t995W0TA2RXatlySkjrynIldgfHS5v83ECrjP2uK5qd7oHJpqdHwcYTNmM
lb4eJBPBYC7ipKChxa0+OJ2qgfysKL5NvwWRTy6+30YU3sNKSl0Ol/7YJZrU
taFlpmli1H/Psmu1gt252llZAyOll3e8BqgMqYsP6DIIoy3VYWb5bl8Zkii5
B8RJU+n5cjUrO4NsY9stPLWWV//NA2wSh4gQz3VYPdiaCDISQwKXdzVabk+O
s6fvgs30N6AuHnEVw28+NzRdA0Iq9De7MtpaQKUscthJu/RQWTqvgK+4Y+HY
1Qj3MiLZoL3jz9QrLwJAN88GzKo1tTyHh2UALO9UZKUrVtlaIJkGuK/sjKuM
U4D6ki08zBfKudv468TFld/6tz/2RmRkQnX+cGRZRl5qbtEJXo1Nq392KxRW
h4gJAIVlToqacnqUXAjRnlM631I2X1p9gTypvtRQz9or675EKoy5jknUOr/W
u3wCKCegiX2zKYOfQ3B+OvWw4IER6WEqEg7b3kGoq0oc1JctGRHCtUb8HCJQ
CXhYAJnk7zTjhM4WWG8RGtFYRTYMfHcV+wP5iupfuhQ9UcdJa+2Z94Ca6aSn
W3oDLw4ziuoJjpf5NPbQhEC7vXXwVU1Y/DDLLqAx8l5ioL+e+5Kn8m9m9MHf
l3pXFZvi7Qo7B7+EAC+bcEruNdctGKod6Beq+UYBjOlpO/5nQb/2we1doEjW
AyRyzLB10P+sWUvzlZrgwKDzGOmOqYuIGm7kIzEst6OUlFugckG/0x14H1Gl
3pDYKn8ikmrG6YmxRNw/YEL26YwYKkiti0eAbne8fyHgcXitSJA/ZOzZO03n
A2JSidXiCE1qq6L2AZ0nuUhhRO07FI2rNJdRtBp/5dy3t7JQFmx3UoP9qlh/
AQFvqbJurcWB0edkskxPofxrfSO5M8p6HW9ARfsJzpYmuXOTcybRFBbhn2bV
2+yi+It1h6sabx+dlqhwJ31dSqlb0TbpuMMyEG41pUbX0FXeim/dCFaGPjTd
fPPqJR2SBjBiOOGqUiQo33ZL3zQ+53afhy4Dk6ux4nwZ+oe5ODv/08gy+dkq
uq1ZosflF6DbBwb4bw+EG4RoVnlkkxQ9ND765yv0YCF2X94GWV+UUKByXLPJ
x7l3aaGRTvCGnGnUfmkTK2F4TslaBRoiTS6p2DzG8khsykONHyBp2abkz3p9
Qx038wJGKaM/TiuZMNqXyv9W/hgNX9lnplFEW8yZJZJ2qy2YNWazTaHHbNjS
8ll2FCwdKsSYvDNLF71fWRNo7DbaGLItdhlyofbW1X4OE3B+Y43qzVK5hwyQ
2Df3ZhnFCVFPY7J+9CIZGpdrq0oBk5IT3GKxyWTXmgFZGmHcxCOQKIhrDorR
gZuvJ/ITSyn6QPLZvU5RqYfBfwkKzug9oTeKbktts/B7rGAXWVjxAOGoLmGs
86IYqzNifTsXfOn+7zpXvXRfxAH3zR8JiRHaCSTlDm3o9sTxEfHEEJqMZ9Hx
cxY2ZL+SZVhFCxSdX9ItszGQGc153curAc/1cV9qQg6MHzeHOpn7XmZRyUb1
tJqdw9jwBO3OvZ5Ub1GQjxhq3iQI9D3l5NPlZso8Kak7EorhNnd0++pi9Mvt
G4cPtc3ZX5WxaaE+NEBcKczljyybc33xULACkIfSPTlE7s7jplS6d2a5WqH8
frtS5yl/deIx+iDGN8S4siS/iL+yZBg3DztFNBmljnOH23gXCaTsraWG1JCM
uvaQOHgd9jUMchIXfZRehCKWvSw4pfdM3TIRFSLwePV6H3+PsWtl47HGcGPF
TSHYkU4JmIoWB+1loeWErkVMdNmxRA9HNTFBNf/1Q3zdYBvgK6jZIIRKDlp9
35Js6Vm0BuVH2A5uwShjHXrbFoJqdbqe7jZT8B03DTHUW+yUKOdVBqHP2Jrd
BOM9XFORQX/imwwhRl7DWr9BXHWmIK3BypmpiqZFXSuWb+0+ynGmkoziz58Z
BMQ3ETecoY3zt0tW4bgVT6yMf9/cAtYaaq5IJqzFiYTSAZH1alSg3MZlAH9i
iJo01KhqS5/2N7xi2fk0l05giXmK6HLgY7ur9FKW3NH8tFJ+P6hWpf+WWqmC
+65s4fkcEuahddTjqj9oEm6/iGxBvcz9RR+LF7/W0Ak2x2FBu9WamY3BjcE1
DOSp3Vhu0rhSshNR9aw15dKx1ebMfXB0Jqnt6hUKo2YxUSeuf318hIKtsWKP
r5QrOyqUWZyB7yYTtK3uA3EC4OKlUvyYE7AvmHe1GnsSIb8h3zw9BHYCqVBS
JUVee+LyhwKd+5DmcOw1oNRfTgLRuyJHETDQ9vzSoF32LozNSJHKz1YO6NB7
2phNWZ4PBwQ/he3+Mo4tTIrHpNajXcfGVxFWurpNGAMQTLHyqp5FoI6VnXQn
XLxOcx3h1xOCKEXKyWTSz9A4SjjO5NvLmZJ/3U2wvZbGjPDCOA0+kiULgVZl
nhWEOVmmy815AI+jw1Vx2O0Ey18UHa/ytt/xAQc7o5kNaf7oiC5VoKDTK5hY
GVXHo3I6tKrXM7y9SXfZ9HL8QrAZrbGhk0tekYMFGjaMG4RCHDD8vMfRuCDA
m9vsouR0u1FK1PtHQ5apf2XfafY2CXiQMHQ5tXRIDILBYuuplTuG+ZSUM1Bl
7Kx3OPe/HzCaLKVxeMeGMoJA1XGl05og1JXNv6L6wcB7UQmT+uN0dc8kFqR5
ETs9lgK5QHtJOOGcDNmulSp7k19lFcNXW0u/Lc6fJECWsj1mNolTpt6z6ZI2
k40nP3tfR7urvACsiMb24T/DAsXDV9qeFA9sqpV+XoL61rDSz3YNFPnDObFi
3ezDL2s2HGBRuWoLpTds8eF/gWqI1+AOI3x6dV5ok6VBEDpDsYL4m7uzmBvU
gczEELI9778ltC5/cYQqd8OagL/mSKmH9aMB+FshgxUicRAYRuz9OmoZmqXX
o2ypl9Tc3Qd2hICKYWzPEWPvhfG4xR/zSwV3p5IGpxjg/VbDFSGiXW9mHy2C
WAlHrZ8cfnupLXnkxhaT4OQsLrUcO4GYQdy/cbQ0CvRsiltRW81VUzDsPrMl
i9hzGBKy5qSjP1SsS0CRzDEe4+urwg/COeBvkDypnmU6BGjT/oTGFE30M7hE
xqLnmUDujZa6ckmv5yGNhK52VXNKGavisjB/Bi4tnv6tlHJ+jU0+GtBWIBA7
E5xhaJRPxEmwqEXR+ebJ6Cx3N0PDOHepAT1ZgtkOtpH6rA7F/8Ck23SJgYrM
R5dXT4GlLh9WvOiiHyBca4O8XhMGHXs7qcEnhPm/09rSQpaChxidWJxGAnC1
lp6bZwYiiwdhdVmM3ex/lZUJfCEyUBYKkjSPLkkdtT/7mLBGf5en975K3dFc
RbNNZDX8qk6juLW7TtDg1oO+oWEegGCEuNg5dxOjVPdQ89as34zBP9prCfU4
UAifnKPulRCC3OTXjyelU5dTuF4ed/d5RyIUBYsiyrEjZ1Q/iwCJtVVzC8OJ
3A8wJlYo6/BWy00ipax1UtTva7d6Hu2CkUXnkhPOLGAOcK4/YhF/gQ9wrml8
a0KQc3FswA2Ofdc7C/zsOiLZ+kPRT+3F8FC3EY/eFomXQ7EvZsY061wuqG4P
UU/L4o9jcrOhCIypR2hCYRxuDvxke0O4fLGQFI2aSfk+wf3tzC8wq55bDTzJ
Vm6l1ou+7MI4h/kYRJOvHmBl+c6DUNImMFzHWtBF2xkKCzej6a7MPg0F0/+e
rdqizI0Go2WAW2rzqIh5QYlGLQ++SKdBqZZxlV6DA+7typUavv+69W5n+VES
sSyrWPZnJyy+q2gBjNilFSBShm2QARrxQppW/Imsa3D7D/vMVp04uUyVRnZU
chgAGHExCAW1f1IJCWLI43Yejq9FkvAPjTAwVmXi3iRTitQv19ogf+AZFOQu
HlZ/DMzaJy/4ll9kFWyQNYxt/0i65eVaFO3mk2JJNDH/1r5HC2dipGJFyXgp
bMDtzE3+Lkp+/6ROjl88yU5Gx4Q2xOxjuoyK6WvkOj0cofEoVpDiV+1d7XQL
ldR4yTEAEiIXjuv02Rfm4qq2OUA2k7eZI6wMdw2V8opIPxyY0hnYw2JSRzQm
PraU6dppmdkJF70z/20ZVesSX5Bvxjr6/daeJM6IWO6aN5J+kTaxV6y/vXGJ
38tspW6OVIXTpp0VfHGEmeKq59gmAJEYmm41NK6K/kX2jwDRdaCDyUX/3dlv
AondMo1fapmC508T6vM+dLXW3X5cQzlI09wgac7+nNo9c158e+5aTR7ziPRc
8TqQYGPVaNG5eVbefPRyZbj03B/Xnh1dTrQxP7dQqLr19Go49E7da+tD3Uhw
aXDvOi/TKsntUxa59d8Wi3RrnwDfMX6vSxzXEx2BgE6BHBzqZV4li7v5Cffl
OtQrXG2bLzWK3n/4i2mmj1600+g0ud5mzoudHJsTUS+Rys0U3iLKCKtO/BQN
RaSD6ERbdovwj3h6EQcVqAlCexq/aiPOjF47b5jS7K3XJ44WD2ryPeUSb8IO
PjJY01DHq2NYBQmOb9I4Kq1cz71l2qne9fb3IBYrUsTR8GJcmop0xsfRWUBf
EzCiZOtFOU3STgB78GAX8WI/cTHZVpl+UY46eNks9F5goqz+lV45wLkqE5qr
RTrYj169SQ/i+3BbGRPCH5LyDvXogEUDmebXKNQpNmRtY31QlDUHa7MWpZab
Ea/aZXrzuUrD5uBTaYLk7yDBurEUwejTiiQL8fbSGmItbHMehFxY3Iv63qqG
JGNiRA67evhM9Ugdk4tHhjuVmsCumpkQcW8fZc3kr5i646fX3ugGMwFMKrRk
L6PsffcX6KHB6ofoqXcDztPZCULCffNWnA+vl6xM8YjnQ6u+Khhee19MQc0a
pvIfci1RsDv1aPdFearteAQYnhmlXn6MvDNdA4UjeR3VPhZqnxYUrYRpDqvV
O4eRsbKClCubrsG5ULncXFxGXLQfpDrkefNbvJbKtfSzK7AP6M5YFZsIquOE
7WuhluYI2Boqd5BjFWB1hpRExtpYW1uo8g73jAFdqCCMLpNF642IuK1xwN3F
gDUv/hpHY8GmeEAqap/rXHJ4m35mwo+NyAkgCsqk0viAwJCFili0y3s+3T0p
444AEpQr6ywmEybSrjLCANv1EgK0/YUfasPPT6P+LwlcUrsZX3mQV3BREHmg
TKsia4wzPT4YbMkmS3FEYdpgonOCxMmMDaH5w64ZR969XZaQlj/6H82YsqdU
niH4FxLDVHkSFSBB3vFHUXxgYz3pKCjLsuZk8oUc+MOF6AOFhyDxoA1z/f1e
7BJ7lnvQ2YcuK/UWPLOghxqA/Iuu1E2lmUg8qjkr5QJzWYwm8CfVrJKpLwHW
9bNhfXhoelRyrWBKdRYdPLTabIRNSmSaWPWqT1P4Q35ceqaM2NAiRP3w7D+D
nqMvveFCYDOTdtpiSt6M955JB3/QTglUDiDKUmz31/o4PIPDEhkZLSadH7mH
cOLhaBonfonFgSY+HXjrH1qtU9ac96Tz9aHrLAMHT7Ocx4H+Z4aeafPhe/Cm
/XES2F5MMuTklssihkZHVOQRyZnaQd9DB7LfUCAO3aw7NRECbA+cw2pua68x
dEiJdHJTzFMxh+O5QFFfMPaPiK5wZt4SlrOAmyRXvkLWwKgJgbyRF1WfwwKj
2Oxb+MFVkmmr2IfbDUokhxDfg9l1/P6FNPXw0PqAjtuDInck+MqrUBSlefJJ
xuDAW2clLOMo2hTMmK1dgOibO+EIn0cRyPlZ59ENxsPSNhUv1c1GNQdsc2ut
QU51b/2WqFAEBam5hqk4En1ANslgEA4xN3kM9ZtmtmGm8UDSKn1xXV+y4rlI
vy95lPsCPpRJp/joTvG1VrHSjhJfCZLtjpVwAPWTOBG7Fu33JmNzZCfEZhyE
voWw2DZq2a48igBneiqgWyRhxDCWMA18mOZKsSXUuvBeMnnMZLachLcPgw90
RXfAdcXE1CrjuC1hnApCutgudIdLWnFcRV8hgcuBNCwFe6K0PCjxIamsiCfz
gSVeDj87qspT0KknLBAXr+u5E+JkBNdhHRiqsH6UR8/RM/SpW1C5/7xGKwAi
MDWYIL65XnKQYT93KiOL1DffEMEPuHJC8yp8kreCgLTho3vlGGwXTt10ARBM
FLTNxn4GCXXXFkdiL34CKrgNhX4CeOtLdJ4ZpxwLd6yr1G3T3Pp+IqAhVRpb
scutHDdufewSERLycg5B/HbsnVGt55k84cbHrAlT20gCjLrNGUedpDFsDTJy
AFPQq2H5xBOj9ls6RZRL8uroQdFUhW91XBbTh+8eoBB3OgFO5ju9cDPb9ylt
yan8B37yQ3tICDZEejfiCIBt7gC4lRdVw90N4QU7RZ9fJHWgo59R1lsftDws
29XTGOgFYWMZgD9ftiqzm1xK70l6Ryw+kDa5SFsIFqjS16zKI5Kv1B/hdJcf
0jmkWfAvN9/84yw8Wl11FFZDDXN/3W/9Vo6P5gJUHWYndTEutNooXx0ux2iW
laEKjeE5BvCjslE7rMT9YhR8ARSxZigMZ29BzcYb4Yf+He9OTd++bgVk4OAE
z3vZhFukRhXRqn5wjzBViWyuDIPzY9+o+qXBjkUP+A0JcVJyGcQ1qrAMsBi5
zrzxSvd5HINVJzlTi9nEVdt60wpzmJ8f3AyjrzRR4Qv75s99bz6oSRnIjksF
AN4165kPJnror/Ss+vZ7TUEKZphT2fc9WjvOienBitnxfrwraacK9aUKsx50
Twl2x2Bft/E0LtQQxkivRDIGVboLKC+Gz2UFMGTPlWWJgJeKph5/JLMO3XpU
TXaT3fVz+MHw5K9FVIbIGUslLrLkKX1MmAxEhsbJG5mgmMaTX/YX8XfuEAM7
3QBOEozOOIaSZzLgqubQbfEDyh7nl5SMk50oj6dEgI3EmUzpj7UiLDP6n0dL
nxYwc4o3mSf+uVQOpsTGogUh162s9mu24p3ahV4W/Swc15/oYB/n0+NkR5lH
2c5v5HYO1CbE509m1Wy0JV3yrpSAjdn31pddzLUkXGYKROEthxi5S7MtdDRH
ei4/9oCZX57yagXXVWM/Sopens2GB+enY8eeH3EbT0PXUM1fJXfWvvRwkrLA
bBI8lehF+LGv+AuKsZUkyKEoY6ikhatspiMcFkMoGjdv4OmBrtO6G+CaVu1d
9E69bhIu/mCdRykMvErk25eKF1X9mO8PEZBPWuJeTOAvPfVS0PDsIyzwcN2h
rnouVUmxWkdpO0hgYRXHZ/VzRhRGpNm/dWksenXeYatH+y9sNO7eBoFyLrNs
q9E1bjCPQ+2MCRBpaPvVvqGH2vukDjozG6tq5+ZflxyiXrcItoVBu0wTJIKX
TbjkQMlhQ3w/RbI4gFSgz1NJTdAxhizdPMM8EWvS1bm6S7YGs2mXiCqP/VlK
9jZWn9uOfbSizqBs26ikeR7MrFv3RvJisml2f/koO3fZ7uwBtE9mJ8GKa136
uzI/lw2RPLj3IdTv/SXXuROiUolK65wG5N3LjvQLHzgsUBa4PlmhBz2QNfyW
f7CKLUpd3u6vXy0iKbXCpLbzMbvhPn05O2goc3EyiaoOx2ccgyR2Mk2+4jpS
ljtSdl292ZijMy89uVJkwryUZscaKgw1cI7T3nvgxf1ovHvkLw/8YlzuBQ00
ip58HvWhS8wixF+58vESTJ+mePY4GE0X9taitzCoAodJdOAS8QZJTeQpPQcm
oZ29RVfamFk3ZpoqTI96Ojmo3UyovbI+lYfGI6AijP0jnB8zko/AnSBvQ6xk
RHBHNjmq1ujOQ8lnZxkv2/J0lTzIMNruOUkbzEi2P/swctarDR/8O9gkUamM
u619slEd6rJGB+5r5trOA/TmhKqWrbSEuMfcT6XJHmiob1BAoVQXag5NkTte
bLFKgnuXNRbqPWdq/BI7pQVNHl8kZCOQPSCqdAbyOmgM3eCyixhajRtfu2m3
NYIEs9ernQ+ektbqWFEOYPscaiPLjsu5W/0D/bU8xkS81hP3JyODw6L8unSP
vdr27YIFBC8/zOXoBIRguEssZajsGiLb66d9buzg4SRG1837pYsdV2t2k0ZD
Bma4YiGLv14Olz2SvgbEfCMxasdgx910ygKAqNUf9B4ATeoYg9wgu4Es/1mK
izaEQD8Q7zFMutEL2p/mdgAUB9qqEEtV6v6yEMKX8I79i0PHIyglXXQ0vi19
mK1aKZIO47tASUklAGGFqXLWJzOTjfvwvI1dXM4XbzqNrWfrOPYDOvCoUIyO
70k0imhtfHMoo4uqzY1eEtavsAqaWtV04E3Bn522OH+NB3l25/vZFoI67YIY
rO/U/xZrutfuip2fbb9mM0mPJsLjQ5bHcwQfZOykjpsYdeTfj3LmYsWt96cL
uZco3llBGbd5+BPgBKYNQUNlYmF5ttX5iGOw9JT/n11DYRdcT+DqyVK1HEXB
e60qEzpDBy9mSIItdXinjvOxLeVkBg34VMBAUfgtC5x4oRz+8dQ7fQuI2fQz
Dar8J06EuAayqP7zzVwbkCSR8PEoo0KUikE398wr8bBm5zQ1tKWxQRyPHCFn
WvBcuoNzaA4hFnp4lOG1v05wHpOfjy/KxhhE5r8iuDcuFJJZ/PxzWdq3zrOT
xDKlDNF9OiStI2SxwY8mpOSJ+mv/UHOYv3c7TyD+A2OobMufx9hgSxb7dYgF
3xeZpuls/d5hYpRhd6AhNqdIz2RLkNPaHuI8kHhrjxjItwV+27MU7K2+TWBO
4A9UVUp2qhpQigcNd62qPC8fHXsK1WD5jsjd1MhudZkrTmK0gBjmMgPAMVNn
ZnJih1W5ZpSWXksH30F9Ylh10V5Oj55QapS/ah8dynDwi8L0hm+gALiMvm7X
E08liTu+Q4vEjFqNkHPZWmXUfOXK3RfsXXMqfG0mr0QnZNDkceJ9g4HnwdDp
AAHN0S+imEsnsTyEdQqg3IGPxrLHQV/BUqWrzaYgppeaZVJLXU94mUi0weSx
t+wJPi1kCt1CRYk/LG9b/8utnuHFMS/g4aTfByn0AYGswn/v2DwPYAQSLb4y
85FDnbmrpCwNuTyX5aONB/jQ6SyQJhlTz3HkNSJ0OhbtOIBFDjIMP2f24VxS
Terh9KWcwbw3VMT3WI3NaikCOr4CdYHGaFL+1i/JOeVVuu/hRre/CjdfuQ5i
AGxi0zKxWtlizGpL3I3rMBwTsRf1cjfxMTKsejCcKXy9JvqpdfAXoEYEEX/I
ze9jyZ2IEmH0wMXWgZm0qDrwxzH4xMn3PIW8zItcogonnVJbKDyqxH3AyJt0
Y1PPO0QmMDnOdqnxFkolfSSl3INWjmHOdFkzrJw96ZyrfWIQEeNNmZX+QBYy
V/dycSneNY8YMDZKc82LKhwN5U3+ToKQsxZg3+RIP8uDO7EDGrVn5PD7Jh0/
yc1MdOkW1kUJoox+UfkNTfIH/nU/9sXPMS/nCYrs17bnFif0NqElJMW3jp6Y
7fmRzKTX5jyGD+Rrs6cYUOsUp7vEO9p4HuHDSd4oJjdgPi9kmZ6rf9hkNJJp
HyyBsNTmuRNhXfk6hFgK9D5WYmCMcihRly76tOaM0vfiFNVy0yWJvAyMbgZx
idDaRlIMu03f6zt05DWaeOgBcKy20j5pbVVgQqw6vjqXOwFPPsyK64s84YNP
2kNMRJOD4ODUqcSK403cA562zAiAkCvvJTu31Wahk0VT9WN6p6c4Ve9PLK/Q
1o797RbGvxd9pRQb1+eAM8JD6Kfy1MtLoDBt9RuYwT06cd2GtO/FZmvGQakT
ozX+XW5JpiCrNzPYI8YiSE1FSKSSEdZsEpSlnKoOBfXFljE2Gd++oXqTR7F7
bvvFFFPr9iCKmx1L6EYz++kK/GuhuSA6tgcly/KKIzkUA53So872bvchadoc
NnuA9VKK1j0yJeRqdf9lVZlzxdESLugLjKRaX+SbcB+3WxaBAXUNWw/rBi6r
3QyRR51GJBDDTn0WGqbN5GEqwFcypadlBB+5DnTZk/z/EDV+1n52i67fjPm4
0R66QUt1Oltl1rOkPo9IEtr+/y77SMdoRs7iM/qMN44N7Kk3zAopcR46hbU6
IYUisPXLsacma/s78X8uz9MCn+W3YNfCnq3c3UgNivE/y1+Kr3NCN95Ex+Kj
xqc/xBAQ/ZPRY2+3UUwN1CnAoOG2iiawrPX4IVI0PyLeq83n3nOSKUYU3A/W
p/omqe8PPK7Hdgo4XnkmVQkhKEia+qlKv4nf3HOclyT8xYfTT9yasMpaeKvy
YCVTNUDssDUbRhD0BFN9aluXHSe0apKstZM9HuvyoXD2YTae9EjcaM0k+Pgs
FPJS6qTIwiGdhRoxKAY2X1dsWoj8YsgB5c31MFS1XGVyIbmmkfv3NnZFc2Se
l3o0wiE++SuJw5rLHN51UPyggkePBvSlOkKqpEezKKabJCMxfewsPTwvcG3O
FO1Q/okjMpMPAyZWjpgktlAHS25E9VbI7OqgKRHcAHjM1JVMTt7n8fj9+f3S
xVEQoIvNlelLE95CPTKYPuptB4lm1hNScrNweFaNK2wMkpG+YR71n3jryclO
OiX2I6+zhOAXCAKQGQoqUnyWsc7PmWtdfo9P9L/XCVFbpQRXWmqQPoulozEr
4wWyXzJcOnJ035lzgDDkhKc8G/go9KPMEiixcJCW5gci/joix+VZXxag/ubg
wRL6rvWNs3xUPPt4VOPC2BZtpUbT/O1GwMAIZEGa4Bd3xCxSQJ+3ABciaim+
Z23pU+pouTGbkKy7Ag3ZF/rbQvD2eq2lpFvqC4LEqG8M5j7dnGcsmOgAbDEV
T0fOW/WUjFSaieRLnhd/C61unviNQMyjfXkueXHfr6k/8NCV/F4S19K7l+ue
i9TPjIE4BwlS6+j7KhgKBW/x9DiFJrVVW9nhuCIi1M47182QWAHDFXc0sCtI
kJOWmYjzUBhnjImrZdbwmct8AhiUzd0t/L8sZJqtBceC45ztgQgH03f7XlrH
rbXCjL4dC8lsYpdfg3DDbqJhL1f3DqVAim7lGXMMqKn5hyqbEexJv8kycbyy
rhmAmkIAzomWmPkbLZUN69HKx0g3KTycPhiY/LJslIzajSeiOp4InSvZ52iA
gFy7uAZ8ALhyw++bcukeWtCL6Ev2feoRSE4UldpbfbECOBnDrZfjqXIJiQcr
ma7+JSpeuDdjNui4awZ0Rz8YatyH4sVNsIgr3ZZmodOgGFONEJnxpbX6XYwC
Q7UU3Ey7g4Hs/ANu7Dh5KeUpPu0lPj9XQ1YkCYnhvBrfeSrTL/nkGQKKhbhL
drJcQ5ZMU0l7UtLI32I7HQpVb+6dHciEoQTTMY71C1owqH23vSxtqshWL35c
3SHJRmt7741G33R5+cksIPg2taGdaqJ+MS1l9WK2AT2GmQ+9oQxqUawrSafO
7CcZbVoSMcEcKHM1kX0h+0Gw1MGiJ9HgcE18WagnHOhNYWweI2N1+AawfC4D
koPSnX0PzhJyfFmt6xX9tdSIjZYDRg/xkTk5A2MxdTbVWKefg1JCPK7v4yud
tuEnkXcCu5SRP945qTbrIzAL6EoqmfWT/OgoUX7HRaBe90x8Nea9Z4J2/Kjx
vphCDnUpTqxRKtX5a9SPDC019bvy6aNPedwcdgFvc5BGW+9nhe8pWHOGTzcW
5RhxLa2CQnJ485YtZHA8RWn6L6WfSfFKIpT6pB1GUCeLyMeoYZY+M36ZwVfO
QbtNY63WLHSz9LFMLXzkCUXR6/0v+xEFlxzmVwexnzHef8cMXwBnCLt/J4FX
ZsiLQqaNWU7jtAlW2zd65sBMrj4AjVBi1feNJhYnGONrcmTgQbM1fk2Qpfy4
tYWuNEAyadYfR6k+NsrgrFxdhx/LYB5i/QNqaD+nOH0L35deY6mrxSwMi9hi
zBT6hGqkzna2Dn5bYUuE/ePRw3PLvCzBGVx2L9BYeQWP7hyYdN87X0zkSC3U
1FqJmRdbRCUbvXwqsYgjiXg0UDsXRMHIrVojhvmOLKg+15eP5Zyk7VFOc7PH
U14odR1T8ZJ6oNcBE67epezTkJmTjlYbzi7QFPRBxAtatTUFlkJR8rFNEz7o
MHc3Hwe+O9/Lym4W9wbbUdlkJRQP+iFRqgv3zC3MIHBAwEKujTXlWOL09mcS
Io31nmlIhgX3giZyadd3gvqAJoAzHYNi1FSJNHkyKe73FPAvLHsiFXdhM2ob
EiZO9UVBMzClYrdlpeCGxVvEseNUVhhARCctVwgsFvGBb6Yq3asFNpUNOxbM
scueqzOzyJ9xBDuGMIcCR1GcA3nbMSlX7Y7te8C/rerHwvNhzDTcQwwH/Nav
o4fTGNTeG6RnGyLfM1xE+zyUMJD6PPEtTzUJDbHAlvWtEap+8X7sk+R/n3SC
XarkXphlznseRH/X/1J9fQ2u9ZOZ9Pn1g1TjDHYzWVUordyNiWEqFa3zSsNA
u5B6P3Beie1bZ3oC7U2BdAC3GWco4WsxhuVKfrTsdU500ZHTXsaA2SWUW5+l
xy1x/pQSmymPG3hI7rkJhvczUBrntYaAqefTyVX5xBhgZBCOWSIJLqhr3EM/
Ay4hIZVQFOo+RvyM57KFgLd5A2/N3CtZNLUbRMp2e5wDrhQwowVtGAIb6jTn
xVaJOt+5M4+zlxiio+foQl9+J0dniL9Xj6VGmd8PDZ3Gt0pC2ne3ySXT3IH3
HtC3YDnMXHol98YJmnStVjfoUo3nHMbMtnjzc4TrSWLjm17FGXllKgmK4g3x
Yvfxg3eYR/36EZ7CpRmU7i60uBQoPXeUeWGaJqp6IsukcK0JkeVLD9LxVfQN
uin0oVemQUyiXsk8FQ6h2OYr9KovWsEbS7yspGA664qLkKBcXx2utmdDAWll
FW1iG6rDAMP2RgTDdtnOWrp4YF326BwESfgmxVhwEUtI3r8wmjN3isVhdClh
cHJDT2HEpHtrBvteH5fZ6ppR4Pkx/TS1uBeZjyPPwonvDwEcD4Cbz345digF
/X5Do2IEVd5kWVQChrw6gH2DF9NcDfaREAs+TvM4Ml58DuFem6uG7YHUhihA
vipCX7Zftx1EoWAbVN19SmXjHj5SiJTv0HlGSANzBikUSALevPUSx3eB6he7
GwteroFNQvr6GFMvYaA3AmIPLTH3qmU7i4j0hFPevgykSpeucmn9t3eXJDWb
kaMjqyDLK/xPemCON+2UCgZzifX+3MvpzJnHfxvMEyp75XHXWjVVsQ1BcKV+
66sSgtxF61vuER0vdkVpiCxA72Zu4VUSkLAg1oTA763aA2sc3ogMkujBiXgM
+ik9xE1F7Zg7halxXw/c6gVZfZlGzKB3wx7qO35niYdc7MUClp/mSp9k4qW1
z0yeISemNEHQzYluA3Rcqef8NC7hAtfwSsr03fGYt0VKfs0yR2ugL+CAeNwU
JBze1YcA8NW74G4vxJInVmbzgFUtw910tzX/hTIrNwfrzbPUynv1nHuyoCyi
EMiaRh22/tcFwqzoxneAiM82I3cDFCu+t/LKppspeRZQ0OGflwdtMCMYUB1b
q9Jgk4F8zofQJ4CgumJTg3T67kea6VzkPRwzMXMzYTyGcI3mZwwp/hwCcmz9
sdcP8svlaLm/H61gRMk34JlWLvcZ70qTOhxbhciTkx5MQpQN8HA1J0rvNOVu
zz4zxhvdaAdUBmOD9oIWTZJH+pjrXCRTyd0GsD1CgFOgYlJRwRfDi3YSjgct
59Mip42YV4Om5RZh+ScDFxwM73tBDKS2HEyqSg34Bx03F10l/ZNDpIEP8ODi
yZ3MQTjCUwvmy4vAHnCr1eJ/4maL2t/r7sAhSjjIkAs7a78SSj+4jaGktmMi
e11LAf3U7DFPb/A/JRLdcC4kdmJIUJkhLjZXyuLSRxc5bP9+gtT8yipD4hfG
wbSOD9F7ZPBDITzHgtVp3FdP4/Okwvued3pSJ/IYxcFXr4UrbiSUBBKI4hnQ
zy/8+RT0zSwm4WQGwVIAJgRQbOXjcb57+ZW46tbGBI7/5wHG3puuRNgKcCES
+4RC0XBrCrKr05MwxGuaBI0DmRJk27y5gqF8uNZbc5xqtz1+qfQn7/N78NtM
x/+WzxCRxxJKLgxibPhf8RVkVreiswhtx+ys9XsEDSH3rrmVRw+QFbxGu1L6
lGwZ8JyQF7X682tMHPTu5+7pr6z2h8c6YunkHXpyJx+kUA9Ek7rW+zCNpUDV
+52KgvHFZwUbkzLbgbYWaxfh7dFS6JGrKXnBdh7QpSmUilslqw2QvHLGd99w
nIs8tmDwclR8ukrqrDyQO1jFcERxLwMJQADji8MDrgHCqK3s7oHzWAnLYsT6
UCwYn2yXa+4pmoGZVMSvcaZ3LN6FOvAW4eNVyMA4Z9a3lEpucUt6U8OnyjG4
HP0UymE3rdi9kFSk8goCKP+ry0ERNEnYx1NI5YvZkLD1lMzN42LqgechtQAZ
3Mfi32x1f7bLIG67978wrUeOPIcbiss8ylDydop1FlcKFARD3MpRkm6TKL8v
mmKDDV6ynsry4Eygr+0+r59ObNFhpu+yE0pzDijc+fcWG3yWFukZHDkrZlc7
0vCvZPqNZVpjMhPSG//r5iRGUaFdLxVm24e3x+N6Cu5+SupTYCgxNLJmq+b/
uOT7mEYk52/mjsORiNzxGfFdv+BpJG+5jBqPrg3vP8UqqqjIlfSJ80oB65k+
qLFqbBMkL7ku7I+5uk+SXLKwMptPWqFxAAj/AgwTE1PxZYKn1pz9QVMQel4L
twDvdkFRV/AaNrwFSc1Bd3f8OxtzGJn6fQfaLxJy6utT/IPygiF3IAYfCXuc
3ixPyYDtIdMom+5AsMbh+6j6z36sClZp+qnRfODtp1yu/Izxcr+eD6ILFwBB
OR4qgtQ30IqvLbZBVCm46+eGjz+2Dc5x2u6GZD+wMakLHjtS/PXPlLj5zJab
YbqIe+C04Rpex4d/RC3uoM1RUalpVBIo6vA4l7wS5rj8Lvpqt0hI7+NTHDXn
N3SjT3jxpTs6mPfWi2cypEiZ2QpicJCC4+JUXMDKLfz2kZK35qvQxw+jtD20
MFgNuYWKJO5GOx2fj9ZvQ4Epao5yYdO+qyc8kaiTm7HJe1cl0+Z6hDl0SR6o
UzGLZgGN46ZZ6JfVrFuP6LUBpNyb/H9/3N+F2iB06DE35mUHBFeHUeJp87UT
gn8shdQbQ9lPCt3NAfE1wmanrRrXQgXVbwT1KADngCfCh2vAA8h4fq4fL+PE
I4kQguChHPTJenZTWRp2fGPihkPp2fF+L/REhdRnptrdj2nlbc7hbm8C3u8k
2MDnILXmTIflu2TyF7ZaZhsb3L2XmhJeyMOx5DVJy/uUyjE5knzZPfQcu73N
byo8VDwS/ugJp1qDFef9AaaqXfHemGWnPf2VlCQA54wYRKqlpMJy9+tomwO4
ONhW/p6LFoImpPAHPoC/LXvo7qokG+gS8TAphw73kZ+kj38n3SCBDaLtkRV4
WJD8jozQg5JFiReAxwbYjbjp++MHA4ixTY5pE7hGW3J9Rt0CiQ3lzyOPSArj
3PHvlA9175bvvssqwjvcsgoHF/CrBykxXKssgd0gJXsSRx2UNzd6bVAHItsw
p+aB7ZyGNh61T4djj6j0o+2fIi16KUTheN4TN6CyOFyVyAZ7AgCdhdkG4GYp
vj3Nu0KXZFXeATMV2cj5CpqJ+IeTPVBIastq6dBp1NCliJXBkE7yqoUEaj7C
F+kcz5U2EJzEMXEpCVxh6b87SMurwyKgaEURP2cO3TrcWRMNknxLbgQ36pOW
pJy9Exkok8zbrHz3IQDm6z748MaElRcY8f4Tp9wpuRhjAjvl9Dw9LuNCkHyt
yf4QagTnxx1vKjfbLxBxDG7ONW3xyoPh7VaDXM35Fywvha6kGZ/Cj8m14yW0
vwQzsCXtGBx2omSF6KmgzpijkLmX0eO4RJWWanbKcLG6RmVKZCMRiXeJ3usL
8EgxAqijiGSIOBae0aM4LnQx4tYbv5tMIk3ECBXBwq4v6TdI7qjQSvZZWTMy
TSbztoshkMRo6TUNDUZEsmsr9ITjp78ovkptcaOAAgyJgRCjQ9SUH2e70Z6z
qRiczsU3pjT0jjuMAxClrUb9G4dxT/uXZQbVvOLYIREx8nUaBrtE30LB204Y
Qk79vYT/SvQ8v9CPsHAbyuGz9w9UNU0NIZScdTQiBsu1G8hnNNYxsXNoeI+5
BL2UWQbxjGoBPOmJEdSEA1f/2Fver0QVZQcKCxajsOZ6JnXnbPajLkXzuIl2
lEEiyF/hWIU7uHRHnBCJlkcr4nNqUsafi0kV2swdwd7adktE4k+ZEJbMvZMe
bXa86PXO6cEbQ5dC/ezlouklnYuqLvjLxXOTHjyuAivNAi68EEXKfCgyBwin
DbsTSXTtXttYubcJdMczboS0ok2wzur6LZn9Xsm3yaDZjywmK5YIhNAdaLkP
W33ynvlzuZagaVsvjG0NsggAnfJQ5CIp+RsV4c6/qPNqTfODU9XI++jKCuik
vlY2erl7Dg2QNCq35PH7tuMOcdrQWFbQ3ljfS8dvWRj+Lcula97qnUnOuVuD
tNaHpvUPdUQ5H8vLeKdw/i3OXxFSOr5q7jSiugchnoSerEUD+Gb6ZbC2zEmo
MycMe7Me27/dYUuYRc5s97dJXps17hTk6aKnpZCC6Q2hyM4ocKzdrd6+wiVz
7pIy9so7PlDob+Rl7aD6AHq2VH5h/yrrJwdYpoxs1TUMHEpBZBv238UaRz5p
eX/eRdygZdt1PYnAXEskC074XslwzL7fX+W3Fxmo1xw4KyKjgWRkIEs6QQsp
wdYKhqvsVr+Vd0GLhKAneDZkYqm6PsQcnDzlaCLnQ3iK4jKE4D4GYU1y5Tf+
2j6a+ZAa4F+p9ghFFmTeTSZk30KAMS7LU8MZ0oSK9fIeeHkP62kvZMDBVuCS
O5wGtPOn+woHBf6dBW+lo/sw+m6eYAXrlOsjHOSKQiby0OOVdF3CrqgXBe8f
7FuSHlfxhJcuaRJYcokLejBDwta97z48m3E00VHRY8ctj3WzDZcdYaObE7rm
qcEFV28OBXgsM7rMFL+7OgcpHnDsEc+PyUyqXmoznKQyhNIcwTMvCwFdc1hU
zTDy1Uu04/jtrIJP5lkUJYQguJeTaTbDWWyBUGAN0RpD9mnklsQ3FqSpd7Lp
M2xcbTj6kRjI8QXr8NsXpPahyXwU66hwWgljKE8HljI6JuFag4pTbnW5uStC
rjn/ywRaaTPEZGBb3IQLVY/LzjqD4yJbTE7dMMt6MR1trIZbKfUKIp0kO9Vj
EM1VcdXfHzXllGdfNhC6u3iL88CwzZRGq9aQrP0DhaNDXowS0Is8cC/TTL8i
4hXXhuPG/iEfsWoXlZevu14Oq0NdIOzi3rb/aXnar/UMGqGpVZom6V9om2gj
KtrTxj2qlIaTyvbbXus/ze5fhm62cxihGD+jcazK18uU7WK/qjO3MBZKqpCV
ugQSp0NA1SwDBuJ1cA/b6ds9vGS9IB2bJacnJIBge/uUvj0cH29mr/FbAa4z
XjSP4QcJvUd2lBCVOfK3ZgfSa+1zZIq3Gj+wmp2FQIw6LaIJ3kShko2HLgh5
eFqmDKCSMku7RfLIfoooS47vdmAqKephjAXrycH1laeQjtDEPQV9SDDtfp8N
zQJ3y2yvSNFxwR+SDQ0+aLk/4C6M1pubwXSG2XFEzN/kciw9PyorblMhknJD
9gWwtsUOajXStreBW3MVRva2/mpWLrQst8P4/+1xVg0Gu0Qjri+LVcgm1Tjl
Lwxdr7iUHX4Fw+WHspT6Hsn+lCTLEoiG9CQ9+GPkICAZYHwriJ6A25vhHs2E
sHLGeKIEzxMlC4l+l5FDz2O7judtWYvROu+iqLasW/BE2GJRBlCjjK7fvrw3
NRT4JPfpJe3OyoWPHPjETV+YVqt2MZ3CVCGvPo8luE8uW/u8RpPrHHWXpcbH
1zh+on+DK7YhhwZGv74mGp2Z6fqyhJLXRx8+VmJUWB0nQEYJbxR437paNGtp
mDE7jfduWnuOtEAo++uAhf6/0OYFHtElGbxB60OxOizznz56TTpkm03E61ZK
iCK9p8b+xhq0Szfi7ojO5BSFQFnuRgs8ndigwG2mCGeVIup/JNpRCzeAq/c5
Y9LHkeXX9X29k5WnMjaZSMBEI6vbp8y7LRR6wMYqtUqhNs4ruq53UmtdiJG+
EgkUJKFw3Qb/2rxm4Cmf6T8qLj8iHTB64ORiTwGinJ0u3v6HAq1ZLMgduMyJ
x8uno1/31j5rBHRkU+5JQl6b5rfRV39LqitM2QgTY4Ol2UH4COvuXF2aLYVS
+MPwsVEDz5avM7qHFFGzc8ZKSJhZlLCcuZ7BKLh8BSQ1gC6ktZyGL10b+vVK
tieVpit9jDoVVZLHt2JHta3TMVzV4rQKC9ZRVNlXkIDRzAz4yu8U2pfsjTAR
lxT10RFLDlSLv2lSB/rgHkJpcwB9IAJhMXMyNJTpr3C19sY7ZP0HWtC6Z56s
Po18Ohyw2tR9Sd6bBw1srhFmHHCZf4pWlTz6ty6wd4sfAqlmU9Sq4glRc+zD
bbXkxPYxjaEj5KPJEmK5QGsBACeH+bHfOFyM/66AgzZALMNkMNT8iJl1OUc4
XHElyYyv8MqWrFX/CSB84G8/QBPDAQ5CL75L9xV6shI86xWOv/YYEmOiyJfz
DdVrQcZFCoiTJ3o18GcpUE5izfcWcA+uD+N4w4ZLtIsnrijQWqcDyd4eQLJF
k5yxEol8kBNswiqfYV+v4Z1iLGGuUbDIzES+j2krFGIAGDM8hMIjKqYpHvIG
ScVH216cs8XvDwTD1TJo4zlBlOzI48ZSHqAduX9Uv2TGW5He81q4sGpOvsm3
VSPzgJ/r5nztVxQ6UvKZ8er5PJQk8F+f4dTILWiL+Q4VKOp3b8aYQb62VqIe
ZdhbJOL4JmCZ2uPUM4yCR9ihO6xmgg3Y2ft7riLVLcxhPbOXfU0eS7klaS/z
KUohei0YO29c24kBF0sFnkpYWeEmgoSxdfqZUTT3i6rlkcNcDu89OndjQ2O8
2WQpheuYtSDv+FLbM9nx9bQpWF1dii1iaYaTVslq+82I0HMbWaq4ur//RjT/
I8QwSj83isSs482EmQ5QX5OBYKjpZWnzxztoazeZEdL4WjCco8UNH1JmPxZ9
jcMOqHZv8FcrYbl6RMV3sqzoxKijqlouKRvwJvcN8wgjBjDiNBo/wi1a4Uiw
Xvox40JkX7jjGbuN0MS21S89NW+o/oijQneAKRkPQlE70+nUlnrsaCThGvQ9
TCcjtSXd3yDRkOkheDQdd0DbVcyw7FGIOkgZ5R+J39PCXkR/fDtJbwZPD/ZR
SNDHP36V9419ZxenXPjYG9aeAvIuvQOPvMtmGGU3hmfBJpDCyVZzoGzgFCHp
6hCbfnDmkGkpLeLJuoJLnXBDG4bXjpffZuDUmLqWKZGhzlYdKjYlQXM7XiTY
mW0zIv5lTLEVuFEXRJZxk9TsIt4/2Q/OpF8D0xMifOmE7jI2h2zfWRt7zZeQ
m0Z4B29KiN0T5iLneSJHRcFO9DdwVd+xhk0EIBUoUtUlxvGXHpYMiIcJcESY
3U150UjVd5h8tXgUvaWTlWzKIQco8WCx5OZhS8j62oofSBLPe5O/j2mJuLp6
/YCapuSwq754lilXVprBWFObSdExBunGj3mfAbQh3+irF7qAl7E4+zlVCamT
XJ4ArAxP41kBndoiFrFBLt3pYNu13t2TgDZwNW52J27ArZyy24zs1FanYJAs
LTRjnJpUuFCEs3nlAvEhWLLJhKQbdHqnGYh0KZOdjtSf8A6qBz7saFZSRwWz
L+2VZ6rFZiX3vvCfY4wWLqEk+otSys6GKRSjpnMWQx81LuqH4nK1ge0TpKHV
H5TdnVoPnwUaZYXD+Q7zwqqNga3GbBOx0vPqBjAmFn54Q2I0yuwNEigQ0Cex
B1UDuddbyJIs/oX4VgGv98at0HhVLQ2e1de8cdjO4+5M5PSIRPstKZtnpSKI
yHDZxZnCQt1W9roTCKwKpCBHHsjEoYqAZWHaHoTiUcEEBS/ZmI05FsasjmL2
MYd+oVXjtkuTZ3HaVrc/FNhpoWbDjpXxhObBi/+W8RaAIjaSx+xoU/hG/uWE
xC/vH5C5J+K8bOyXfgMep/eZ1N5fRDyyJx9zBaOMXYxeWVUU6/8vR1aDU39V
DC/1dUVI9GR8QbnlyeouOPj03XLzCsssHj+ZXPzWtynR56wN9nlIa3K7zJXk
P0NvJ4hLqxKfoS/cykrQG9DkmNk69gyAuv4/KVfGSaeDQggrXym6MuqaVptE
hCKuzVmCabTADJSVrdJwLlv94B+w6TqD5cHZyQwa5JhzojrBJV9VEsvL0f8U
bwHvo+/hVEO9l9Qih6358t4WStP6cZmKfWlRO6C93dnUgmdMO22i01atPcSg
YomZ2t3Z0rbJdULaf1pf0mRRR1vq1JQkVun3mfz3fc2puU+ujjUpxsOEFf1N
OVGFYpRyMN2RXNPOK1diK5SIKY835iXNhE5K1MTVk79a29ZV7qa6VKbmGp9t
omz8t2Ho1P6suOAWP0YSIAxmJVVlTdxWPqw0caZWEnWB85TWZXM7Cb6VL8Bc
RQ7z0qtLNGVjmDsVbWeVHfHbrbssO3BX8kcA+VZKPAkFzmCzNZrz6s1dskOZ
AV/WwYnacVE2Qbsa7itgLxCcejy7lvdv/vtEV2olEFizoZV9mxmC3tNKnMc0
5eM5nQtv4bOtsG5+PYlc4pEsNCpVMUxwA7k+UWQTD6K3YNHvASH0ft85DcvT
rbDhGD+G7fh/v5l/KwgJysU8CoJm5FWO9XrsS3np01ocC4jfWZ1VwRzT2qS/
0q8LbL9pl5dpMoo+SpBD3cR/rSZb4E8J4Z2oaQNjVQlqHh3BgubtAm4ujdA1
HjOyF1tDBdYut6IggHC0KRdmcIyPlm/GXtdEBAimorr1XqOzS9vEkZ8Ovl4u
zMnKt6tZHSeFyW44hvLRFVci+mlmtnqdrfoLf7IanVkk8Lx3CPybrp20Alaq
g3MFhML0hhnpVDaef4jiY4ZiXIJXobENOVJYdyZbddyjgLhvgh+WweGER/MR
ZjryXghhvu1Nv/UXby0p33f2XFhjHo57m6co6FPw87gDoRp3NyjyQhF16FkT
nBaVuyoa2LRxaZblHlSfNnyRjg9J9wXUJ9Jzr9UDGO4sR9WVXtf3nq4NBrBD
wsnUO3FRz64HjBTLTGTeJCu38x2aug9xCdl65QANW02t4ipCEDSJqWioRDqo
t60BdN8mmBYle+0ZOGl5YYczcmfrxbthohNJp293YU/aB0Ywa/9YMwABZx5E
n5yrARKsyE8V+UTqceA5VikhULAuXvM8avqquQrS3aWn0hzal/RTTASi+74V
Fgq/gyJ3Aq9hFAMaZYbt8Q63FxdFoGDSeJ0zB88+/8D33k2/ZVaqEUH8RTat
hq70fPpeetJK3GtXcTe7fowWlIolKWJRKFmApxNi42UxeBznWwJP86eRgjD1
Gb0HrkaLjwAtm2GDRg+/FLOfowX3/cLvb0rnhOFj5UZee5FoSBoh2Vq0Kq6u
aW7hbvN3eSk3mfc6OBOgF7t4Gs46hmIth2c2OBS7ZHuPakbTV6XRz+U7y9o9
Da8HDmK+eKC5kM+PzJg0MSd+P1O0Tym2Sh6/f7iozeqOJlffffg6fQDrPuXs
zH1ttJ4Af42CqfDpxNTZBmKo8lGE5EaxbKZtleXMxSnB/NGnDzgMYGQ4ygns
V6rb16VtRW+DqoPVMPTTO6MHv7JkdKDwMUayvja+T7AXLpHJdaVs1agksD2e
3kM5OggMX2TKcSorgl4ixIT3f4Y25WLs1AuRvUhVwIZNlY4/fSCfiMdmjvk6
rS8oINGtTjWguoCk10kQC3Vyy7t+gpHX9ppmhbwXJ9dzQRvPrDxkbh/GtVF3
f/OaSS4Q2iDXNKfd7pnC3AWCm3/iVizcmdHDdaKrjfSIId1ekIfYv2VF5diR
fdot/ug+0u6BLOellVRgvP0TlL5GtYkmMLOepZRguV2CKCJ30/S0Tn4zYuXb
gsm13OaOHZUxKpgnZbRCT6Xh3zvhIZcGBIIGrsUB7EjjuXiNUe5jMlinlVWd
kKQlf1t7DbhysFWuYblxDS0dNC01K5t6cJFlCzZMa6xGinBL2KW+49P4a+vs
K0xOH3vrljiILDsttDtWnlCiuUL0lzgkTVlgjpKFkS+KT6BR6GYxYmBQE9TZ
G4UKIsHIQOQb0lsVaR9w1Qhl+ZpR+i/QFpwqUaRKzHR+LgiSHWaYmdtPqbfR
cknwI+soXwyVyxJGDGzw0AJzz4COfjZlz1uV0uKKGA1/L8XBv6klzVnfZgsn
69cJfB4UEEOkmlwemzFvLLzI+CfzT1IF4Wz5P9V8qJcxRd+mygFKNa+u7gB7
0LePWPpowXCz/3UhkZLCxxnkZvQGd94QslOuJok02FMucb83VfZi/fkSTgNd
lrWrjUnEAvWPt2p18/AAgJtGLcbfPkih1zEo1ckk9w3utAK+aZfWgMX2+db8
gXxjWMi/1KCzLvWRXbRAZh9nwwq4Ozrp1zS5FbKN+bmwu+XcmKrB822oCIL/
OaZEH7m1+N+x+hKSl/YH6ttQsvEvs0yuu5TaxV8sRtRlTkpDFWekHX9tKI6I
dBaVlSgixnUTApiM3+48ayRciEZMN/vx3qok3ky6xRcQpXBTw+QY7FgB5tQj
gJZlR89OqsTQjjYBl/NhlM3WAbBVJWt0EL6xiM4Joq7oiTKuad0ZDb0J3kT7
4rz38NW7Y+IaNh9V1zVNOl4FpNdNE0YwnU2OggKG9DYIvWf3hsli2bnnUqVB
at/JjvmUOJXPNwh3VhOYLTwL1+FdSHj6g165cbYjg7m4PBFnd9UFZFGA8fdS
eFiuMrKhu7Qh9lP1WPbNJy0Due6E2pvaN62b4e+rXPk2fb8IydTtoOcP3tzC
eJgMsbfwzOGNTWk599uodGqGIiNaGP6qZFrKaImrTb20MsTqOduZ4O5lMKwy
ynS6BOS0uC6/28Po+zNWcjRKD/pE+xU4/HMN7tMLS0uxrIMc1V3ek27pJ/CE
nF4bj3y06Hl6XFaSLJD+qn+fbrcQjAKOPtm6hfyGOmSWliB9v8qtcifFa9P2
Q6HAQm7NXWqnhv/wc9f4qYMfQKHR0sxOk1ZZusHdI+Eh0xetoOoT9u2Egvw3
t4edX/awmlczB0yqQJXxXxgTvs3HwtN7aI1w/+M864CMS1HWyF6z6SwZ+/qk
X48PIPWLt5cE5BVmDkkDk7uAnQ+7crw91o0crZz+qWz3cPZ4tm0kvQ2efDte
NA9v7MK0aJZx/Ccw19GfizqvqdZQwBmd7WsYTHa1CLSImSl0vWEiGF+rebtt
M+eBwgwbn2wx4gFdQczmf7IZQwwANXTc95pqk/6wbviY51NPF+ECYML6Blsg
JnmaYQ3XpEhTc6JiY4a5OJhiaOST0iM8vhz/uE9LBQCpkC6EJrM5bdBcE20H
AC9uV5HgFXPWxRM7OvkD9qO4Lcgoy5dM80ID50aa6ux0r7G4IjqsqEtkyqzw
M03m6p73QMbKPDu0dYesDtqHd90Xj1m3aqjpXt0RsDnGTg7UQL2qgPIz6GyT
LV7+Oq+jCgCcH/XKk4+ySTpHri3E6eL2BtyC0yUz40FbE47ZYDGi0d28x92e
16wpbE6HZpXcEWyGqrN3XMl/mVdMIrAoVgoruQAFVI2GKOtvv5Sk6ujce0k1
ervyd8mPCNsrc4KZ8rQ4kPWt+b6RpgU7wkQ6gd6xvsCeeyWowHe/Dpw8C1gR
ouOClT4T3oWpJN3kz+ZWYuRkNsgr1x6Ln8ZcylBf9TDTjdp6ULJ2VkOArAkg
hj5hkxOK+L6+0oDixZkkT4Wbqql2fv4cpuOmB2CKeiCN/THljr5B0NQouJ1i
N5m3gin9dF5nQg5J9I6v3UtP8gwhhJMZldqgzD+QbUrS2Bic1nxnsgOPHni2
UfzLSSLu/l84b7VZnwIrTobYyvZfSpw7nkZ2OPc8rm2446aDFYRl1mrj12z2
NYs3WBgerxEWs9YcVQuySyIBtHXVGhKYRB4ixtOHGIfwHV1of617cjUCvbwr
TIwJQ4ASVJaN0ycrtxb6pX+qQTScf99Z0tMBecxyACANyFcaciKSqJgjqhCU
lNcCbqcygYAnScYshT8zb8Va++e2WDu58osp53cUhOmbprzwovipxqHkqhYY
qD2MScaricfRJHD2VPAjLtyHdmxroyTjjSQuirzMXbOoSqhng9pRpmUibO+9
XF8HO5jXdqjd1TO5ts0LroA95vsKKIIGUMUEmz4xG1Zlve91cxZuUs97PUjd
Q0kQR+s934PhFwSCoInnxcWIDIlYAo7dRtk2d7JkSsfvyGWN4ltv+NVSJzlX
JqjuP+eMoIMmrt9n+P8IlUdEG9hz2wq3nysxx9qzHe7Hxuo6DRkHBsB/o1UC
U/1Bof6kzEjd/LCKBuMJ37i1LHxIqGhNJXBh3Gf3KtljogTSRELCwligW1vr
qLDkimjONadHwKTuLBhMV30xSC/q0wKiX35iS+XxLpfufL9blgjURcJB1Ko6
l+H0prWLpKwDC5qJ405/MQtKNH4o05pHvQMVXh4MgRqbxWXCBKACqJ0EJksk
Iysgon7vu+AayBuTtFWQPzrAhrYQK+vgAGsPu61gIP2aZqrz6eXmSu81zrS9
NE0JxXpCipdzI/GNVnBiLha6KQOCVIQWZoULLMybJlNHVHLbcmsIH63+6Jfe
89VRiPFMRLnoBIFYGN9efoNnxyh7YqVR+5zxociYcsyUZ9nS/LiqTvpcGQVw
Wo49MjsomVzv5RddsEO7rQaajxfWnfHhxvlXdkBVn04XD0Kbqd0yblEOUgGj
xjdMz3x/sL3xH9NWYlkd31smC67lGCIKWCYrnJlZQ0/VPK+5rflSLZLHVOr3
t7dn0pUfthKo5bVNPqNLIKddOBvg00xeT1jAB3iia8oI/xQ9CpRes6HaBR/V
qLII3ux9jfo/dHHgBeTvjYLzoMs8lBfOdZLwUUADwL3jJBFYF+q4Oq2PDWpm
e/n+Zimc7DkPS9GxfVRot1QD9QTmjdlRZhbmuDcdpPi32348oMNZfLhxiNMp
ynAU9Vdjy0C7AO/qwievzG5ZTlq0SF9hN6oLsxeBVekuyuU6x1v39Vwdo0ai
6yetJjnEFFcfvcApUpw5sNaB3SYsY2eaZJdeKb1Ef7lLqHkq1HEmuR7Lm0oH
DppQZu9SXUV8H48AweyUzAFLHDUax7m6wjsUGCnkkGZl0zWKd8h03gLkoAE+
+ev6VO1hrvTBM9/B8UDOG3WGtWWU/VekpQ4Nmt4tGGMF4TskRqntbmRmbVfg
XnvpWBQSoFD6d6BhIn3e6WWN8omnm8A447FapZBpS6ogsb+ttv50eUD2xJiy
3R975DSLdYs0+utJ4kGTA/kmqWtXI/FroWrEo0fJSga7zwcLSNuQbgLxOBzz
ptpLYFnykM8FGhwJiqoEB1pa1PYIXwSSJhjc3Nis6yfzOeXr2Be7U09u06iv
jsniclkOJJ4hcRU6CI7ApF4YyhkxjV8LWtKx0VU6ElYsH1t8k4h+ne5czCmN
ride7QFHRgP2pqtZykHmPfiJ1D/a43uvgdl7+5Mh4bazsNNGSkwUvYpAZCKA
m60kFvboqChD6H5P1lc2CILfOFX4yGdOekijbhM8R0Ye/UuMX5RcfM/cj8zt
8iZDbDzWLuBlFmwHlUmgBHw5psmUxtB941OuWM0mWJ7Qum0dEY1mwnRdVQL3
8pkkTT4R1sr3o+KfHS7gLA7QxmeZEzCDDTM+2HEecmYodtsCMPEYOUjkw3/9
5QIMpY67SROcgotdVKT4dYwEssY4xceM4Ha9ciT6bn0Cm0+MuzGf0PRWvg2u
aHYski+XZobSunMUiaElGCwKjBQsumPzGk73tF5Vxqk1TKxKm32fffGZx6WS
PuSohJtvKKnrjGXen3aYuFpt1nL1K1Sj6Kl33Vs1qAUhy2LAXfWOMV8v5LMX
zf3mlvIOqPQ3aazB4+UiNY588FLLqWFh+FAzDB//yPVOqUyv/A7lHME0xR9e
B0J8bsk+f6bmZ0uYIVA5Y8gDXaVuogi71DfU0aT76np+S9qSpNDQ/Rl9mKIY
JzvU1AJ20wBF3IVINM8f5yM5ufd+073TClQqK74w1vc6YsI5CpeFYU2YGodC
Q5VuhiETdV/V18DyEHyxka582TbVtu1XZqbuoDqbNhdlkfpJ8fFTBFudsbZq
M8QymNJ2TWMRdyVE1FvU/6HDnW5TAq/M/Q4m5QQNQg4kHwowK1dsxBZgO2DL
cExm2fWOjevHpEreEpuTSfi9Gxvrhc95Ipr1U8ePtVWf13FHi9TadwguHKBh
lOvNPRNGZzvXtU5oox8eGWsvYi2OeKg0TsxyTe70F+uEHHn/Kqow+/e9BpK5
xzHvoKWDMsXe+UiE23OWZsbaWS5iZ0buMKE4+H7FETYC5AwaFq6SOGJu7jdV
h0CbEE30EPnqvc4qCAGgpoZG+lE8Rxw/qpSs+E9vl9P7IvZQ3tZTydKbHvg7
I40lh48qxNN4ygOlT5ozaV2SvFHSdtyrDrExHymiw+LSWz+Epu0+8KFXd4Lw
9c5ilF6ShY9hqy1zgLfHJAgy98IxMTKZYSAmPSwWthuGV75qfTjEZ3aLOWfE
9pBvLW1jyJO9jYCrX52n5IOWFCRefs5YrQRPITfp9TWCGryBfrLpRPNCchHx
C6oGNuXjx5hYoeEvjEKIkzCRNDRYcHv60VvkKuLAFz6wpysXnSVTgpaZoxxP
ihLv8XIIOseJhnCRbnsi82QIRQpoKqnzFC70glLmj2chEvEXwpn891xwPsKF
66BNzS76dxJolxTE57Kkk4kdKYIK4PCiV840dwLRPMU7CPF/fDunNCOdWp7y
QphwtTpD8KC+uDQaqm2YO+infApheCcRx0AaWTeYn0wzccb/Oo/6eoxjO7H7
P4XBgX2d3q1GhF3IWUGpntJdD+aw21vv18ESRnn+RHky+6dvMOo3ndETKW7V
KwLvubAWiptUvOIAziATRirqPuLZdtOl2122SmJTz85LEul6O3/je4GHk4aL
wns8UCZfUdvNpaCGzHOJ+B12RuD8Zwf6c+vDTuOQK3EmFZQT6norA2p4j0wS
IlKrgQwJlWjug1IfTJEMcpdJ84hC94W03nAZnQlOnmZqN5yxXSZN17ifR+5B
EDeK1au41sJnIXKpqK8nw3ASNsJWo3gbW5SuQ5GNhALHi/SyGIy2oEYQDg6n
miE2WUTYWgeJLnRxSz1YY/BmZ4EMD8pi9ct/O996hI22nlliOFQrjYl8u+GK
fKNDc9d2axwc0zBzj6TBvQiqDZI/qIA0XcpCNR3WPiWKqoU6ATU8Lr3omYI+
d3TN0pGW/Lcl2kbHLNg+sdBceK6AVolW/nJ3zpVCVuvcahrRRPELs5Nkw9Vi
rNVHfg5oK2z8J0QjnG6Wg+V7kxPBTZCKpv/uiF7xvK1J4id+Yb0zd9qrqJsw
kB50IXBivG0zvJSG09uPr8orLpX8LZAwBufw+V9f9rY6KtDFucbCHt5tQH7U
cis59mhRwdkfTb9ULHJ33N2ENxi+5h82YNU3VWZlqWPgRjQ0mnsixmvWbsgJ
UqSvtzyKvk0TPMuIgXsaQa68NK03pH6Q1GuRHfPMX19QxTbvUaAadGyPkXUy
+hTfR5cx5Hf3EkuIZpof5kLJAARwZvoh1TgtKpDchfJU7ta7QcBN82vCPr2p
nCfQfqmxu4t8gmrCaL3LBKkVylb9psrOMbmjJi16lrPHx57T5dyjd7+ltDIJ
Y6RLQlC4OSICsAq269r5C4lvmLfUBsZTZJLxcViJ+3rRyFztI54wQsZlgKZW
AtrbUhaiRh853l9ZHldGWo/tYRK/QzR9L0T7hPJC7qZRQ7mzFtnkKGZBguzt
CsKQGnsWFjiOWVtyjt0oUxKR35ajP0TQ7S4CcKsLF+HWWUcCYHpOCy7CBB/E
wuS8nI7TaSQpDKesq8Y9Q4NGAcgSPr+38gwGlMVJ35D0puPTb+VScdrd1Kuc
JVpaycOYafD2WvadDgBzsv5wWSA7XTMuIYYr9b95Vm6Ew4MIiE4aip3AOCUz
sC336p6ALpttfbz+2cd4X7p0+y4lOOocufCG3NPmNJlU3wYAkZgN+xXJsGgs
3jmzhza9tWNl+6JUxSCEhL4mZhlVkbMBHHoSg/yv55IB+MyNPgdb2Oq6fOYd
M4unViIV9B0mwlDx1YdXYzEtKMsj1oN/bcTVYYBq9/xDnq80T8jPbbZNZGZz
fT723O4sYqTd2HKpK3/JEH7KpfblEUQ81SYngTdg6Ajh1uPidP8RhHcfi9sr
F1oU8qJHEeupvusNCra06VJWxIczOZGYy5lfM/2VbJ9KUlB25/ti+ejHwPx7
eG1OCJoiNqu+xkRyH9bGQYCn5yvmIA48P2gOI13uS8029HjrWh0tsufYUTKa
gVe404khWS4e+y5Wpp+/JKJ00+ChbBVq1qTrHxH0+s2v3a7Sp365w2Im+kc4
m15+8798ntPchsP8whtt4UNhKjzKi6DJv6FhtLNj44Uw/uHJQhfWCSBVtioP
EZsmo76Amy0IyT6dXACbY/bgElylhFt8RzFj4xn8yKHHMGWEj2TMliC2YmQ5
VNaTMMAt5sONjkIt3f1mdToLmUb6Us1eJ8TNtHTe5H+61r7/k40Y4K8jz4Qi
kgvqmrXh5pT4E8r/oqtJw++wMNoRRZIcL7zCNqOptARkm9tlOA9mPIa2/Jj8
FpwqAG4jBWXpYaYRMhW2MOvNyT02THmAl37xYOvqBCxVFttaK2+lTtbG0GXy
k8xJ6WuzmR7kV6nWzid2WPnUe1dgInUjBwJFb36KCcd/+Hf8Z/jaEcng8hCd
/QpGAY5QKxsRRly6Fo7+i6l7rxWNg0I2u2MN2CdwOY43SQXL4u+lWCfhVE+G
ZjkXLkK1AghXq9S72Lo6rKiXselWc1LE4GVMgoCsYYtbc3l6Evsy10GpqyY5
o1uuY3JzcBNTQorC+9GTd+TfGHCVekAZK+1sjeFvf9m0mSYg+9mnqeHTo9YL
d8EF1G8frXp4EaVbRcBdCqkaRc/YaDMBDsJZV/urxo8z5KQRlvBrGQHLS3NW
6dYD38kAV/dZ3cmKDrUEopjh2mKySULMDzix23ONv4jXX7Mg2GjJGaOkFRrZ
LxTxIw1BcDj38wbgdySq4tWLA3H4LBSPQu0tHR7mLftJ6EVHoakOzyD0lDu9
pQ9tI2ZEFMNh5Znm4S+WQwwYizX+g3/kO4UMK0RoROOrlS6HMLj86Kg3VRS7
mS44IpojO8Lw9arzo4q1fEKI1SR5tJC9Ad3hSawHvJOdazOe1Xgqsvrt8TDu
SIqMzeCsmZEDf9u2r7MaAWa5aPjG+x70ztZbyuaD7qgS5dsFKExcgGARvisW
IGmBE4L/MmH+m3fRjkAEogZqZ2EZ4V5HaGcHLrTwoTplAF7zWJocMSQy3RPN
uaLbGmLjJ+PL84cqo8q6edbhW3GcacT+fT5MhMkMSKLend0f/dSvReR0CXBt
JSB1c6XoW19JOrcg5w2wX3Homc2yq2CifOqyZGWD9qM5GEEeb6z9G569rUas
3dExOwQStv1mH/8Wk2zsasiX0yjR6wOebVudsYjXRmiSBgSw0hIt9q7HR5ql
PLVnC947otjffWPEXjWzc0XkENeJ3WvfmwnkUMBwuhXJYeYs2vRec+qBb4lB
EqsDBFs+DDFjb5aeAg2P0+SYmzqQ8cXRvoXix2pmJNLB9cNweCRl/YOibFMG
szXNJnJHR4SKVb37FK1rvrNv7AKO11G9W9oyxpSZ1aLSKjYK7/KCXlY9CEW2
mO24f+Ij/Qeu0WH6gnidDbeNoYnLzy5u6bv2SulUB+vunwSVJqbWkats8S00
PariCjexE8R8+ZweoYAWjFfc5JpHO28WaTctzdX9K3NuZBL60Dx71qJlmv5b
8SAYXQNUxvSBhCAJjYOYfKZwvC2aDCvUP7F0ezPZMlevYA4ONsMHEsElzBeB
hiWgM1L9PGg0ct/IC9Z7Z1EbJYendk672tByuU9DQdbmSGg0BWxl7ZPEXekp
Hv1+g7prQtN7lyWP/51mf4uzyYdHttIvkwArcp/SjUdzzR4Gwn1SI4RvOlX5
t2rTeErSQ9EA0sX64PTT6Ysvne+K/+woOFaICTz/iAJFrcK1+2P67WLGtTYY
BPYyc3pSAn9VBcuU54542pzUAsDOZ7hkyywRqyO70d3DoI12MPrci2pCngsJ
GpFxLSl+I+xgVz/sZc8Kt3ZDiTZBtzE8/GpJX1tZ7wofKK6pO4qpCVUV+G/1
tM8rRZix+OgGf3oJuBPbgjJ55cTl9haQJapfG/RKQf7A22Ff4G2xFKPA4fM/
P/ZKL9HC6KSW8OYy6UUVXTKL00xr4+UuFqh/SKy9P5MIZY3HAvMTw2vgZDQI
Mx0jiqAT/kE95DhKUFEQ30NNtIoQ+uSaHY3ZhA8DAPOiwj8gAkP8h4HomL5N
pgoupaGssUiQ4tIsqi7wOqVDQayruTIgFVj9XPggfVxiN/khZtk1pLW7uppM
wDV6A/R/oEERc82qh5wMqRyqQ60VmOPS2Im8Ogx7J0fF11dVYMb4BuY+rnPY
5sdMMrnOtSHxGKfi8wDqPQOYklAx0iF7v8/n2yy0ThaitBKsXvxfQyDsixBP
1hmZtIq39CSv+y7JwMMHpVyHVk6O1VgAxILcGDd/vjdq/fJIhXfqANAnAmqQ
RZq3U9b38svdrEpCkxBDj89t8gjvE3qgTxfGUypi4kASAYF15XLgvBerDIJ+
QGKbmrc7X8E3vkTCzPPOJ4sHsa+wGq8S/YPUBhI6ork4cvyPcGCOUdgrDoHN
Qsw+IbiFS/OhHBRqAWMww4J1OX9l7bMfUGNsubP2lDjna5SIsG9gOUlFalDz
+GcgXBpLUhPZ/nse/w+4n1DdfYNya+CvXa53NqEDEoxoyn21Hpsew7nG+9zX
74PRV9viMOZph6pnfCWTQrRglEgpvfR/qKW2SdJRHMrizwtaEJs/MWNG5rBk
BpamL+I2L1lY9idAkuE46G65LdHNTtIeIkh5HWsiEpdoOljivVieH9vQPajT
dz1YB+Q8xfIs+sANjF63GTHei5MgEV9b11M4+69716HgsLh1N4WJ+pVDnCeH
MKS+1VJdx1AYR9dQCCNXBrQOH02o9yCAfryVmiZ4pS2hqDU8BD0wiT8D8F0+
4taWMG9TPcNeJercP+FcP56AU7A6WoYWxg8KOMCYC7G80b8dz7k0DD+IQYjW
oMWXpU+xoGP0dIBflPQwucL4Nd5cq/MCaHZfzzzFHbGskjv8JJzvRf7WhjNz
sM++bWEJ0ttrr23cHWTlkQOzen7QljgJotcfsAoJKz0Zh/IQ02wwZI/6n3Q4
PkfpywZyFSdGwGUc3WEEaTwIcMtYx22Q6CuDkviDD1pI3tk36GnXENMLJFDa
P8Qjif9XiLzMi8Wr/8sueKo1j1XH6usdAJqpNFk1uda2ubWz5JTfKQwQ8xhl
9v4npiWag0pkelp43sttTLlO0XehWsvVJOorODrG+9QX6zFuMKhCD/ktewt+
gKdRSgS+jY4ShxutakujimvaZ9/EZGrDekx267kFwijQKhXRpId/Ymt7zZdP
w3sj+bpHU6Yh4AqhZZAeOKWelnRrcTs0IV49sG2mEJJNHOfbRBPri4izDqIK
HzzH/YTBM5SQ18+Mv3bHsVb6xzj6Mn3U5ZlIXykBLsOL9d+9wtZeSN4yvc+m
HPEej71qra3clDpI1eGVTtP6V6NsqEHSGvOx6dvU9pZoJL4xfObKoJHogliC
ZMQRUD7+53crdvv7s9vL3iYRrFd96CqFSkuZ/L4pJp5keqDZ9TfZFw0+0j2o
myc9FW/NRetWfTt7jZFyNIemBHxTqQxO+/TxN2bJfW/whzB71/A+BQsSPuTl
P1fNK1jqA3vSg95DeaRScM3NTXoY8JBhq0FPq/psBfMm5vwM2N5iRP7pwSUW
A6YJdrtWh9UBERfQKy8SIXFXdv0SWG8TTGdPU0WYgLp8pFXO39XfHyVf9i+g
oa9Q7JFaMJIH5eUOOQao6eiR9Z1fpsnLggwFuBcepSR8aikjhZ3KOEQ+4rYy
V1WbfINbiVlN7/jxCjc1Qr9eZK2xo63kbqJOTlplOJ8cZWS0F7QjO+j6QgZQ
ZlxNWQjK77qsesIQIODJBTGVIvfLaObwFPRvXY1/IFiXETmJhkXQ+H8AIab1
ETDD5ZX8okmLbrMzwOLxDY9GhmiNRIMVyJpplM0DsDTILzRsKSP2ayMte+Gv
q0Zq3Xs6nlc/muOu/yNxlnZBxR++jZteUJJ/XT5WAt/t29SLSk4ybY4ZZ8YJ
BvmxLBBQKjGrB13F14iAFlN9LlnzMtDZvq+tuQC97lPM4DWfZvCvCqUNXU3g
2kuAi5V2dXa8jN32FEasxy02kV9Gq1aVBSCHNR30dfsC+XwAprvmfoFl/Les
stT0wjXcl5g17z1lYEMcmPeX/Fj6N5pkJbiI2yUIB8yWzh9w8rx2lrs+HXjQ
WZy79DhK9/G7ueAYdjwTHgN0jPkTLRTXjTyY/9A6ifjBpBBq/lBaMi6NfZD6
fbuc9gTXa0g7os6Vs14Dql0/TL8JggTh1F7BUJqibVuYqvIbFkRH97e43cQL
fu97dHqkmcPmaHHUPl7MhoZY64llvlpnnTPc2a3nlNvkqt78E17Pae80Y7yl
tnFYa+HIiolnXhbKALo2NCJ7OxQ5Q/ws3l+1zYAM33IkTaJP/08K7u2QmJoE
sg0NaE21WkP1xFMmcKOi9JMV5RYhGmssZN2irtqX6sVjvpaxtd4aVTRVgTqU
M4A0zJattr0csovlXKL4mMAazNN6uCPF/WKul6z1RNFtmtVGtGywoQkpd5Me
jQgyksjUP5drVk8xoZMUqyYCyFLpAb6vvo0XGun8x2m8+v410Rhz4Gp3zEyE
n1/L+FF3o8uKi7Io4oLTTaW59zkq7atUnwtP4JBrGgmZT67+JYSIEorom9yV
j59ec8TU+mUW+QfqFsHnyjICZIMbnGse97XRTHsr84ct49kBC9w1i64AAYIW
LYNFkxddDjGeJ5x8ZXyELnC3zNs1ui3Txd7rvLopWB7rvku/cobf0wbbkFs9
znFAs8MGZ8aXAu9meL/ciS+iByPqySjCeasbVbVsRqaJRoef9GW8HK2UGx7b
wpG967hAVqgg6T7B6MjrmKKS83zARclMmGPrCJYlryEVd7wTfsWDWqTugVJn
2lLggokpsEUw/vw/EXUkSxqmuy+pZMLYNGy+P4BhA+4qnonUHN+aCZTS8DVx
iMZHm8ESzy7sybTKuQeB9gGcFWjtb8+RUZKCLhur5mdEqoGEyl7iyI3ijBnY
p68Imk5nKYAVfUhdFOyr3KM5mmAPo7BLKa7Ob3wmzpXAa1KS0lDL4NoeLft8
RmiSbj6SUoNNa3/6Tz/5J7fJc3HFQgmM42DSlAbvOiuvfO8PoDkhD7XLcs/i
j0dWxMiNfdf2TmhGz28uIn9MZr6z6dxlcM44iQRATqh5aGgjHU2EC8s/VPJ9
Gtze6XGZrEDViHLYrOhewUNd/yljBTrNzld2Sip5aw/6YwPKjvbKwzP7Q4uq
ZWdSoyjMVPMgBEiLqg3QcufNHk4ehLtt1Emz+zCxMp3xOwUa+8UF3Yw2nc7m
0+6GdZTU/6Jy7ed6irgBjTDOycv3Qmuu+qgNnZl0qN+Iaxcn+vKQ3Gww+V0m
6bRQKFn0AX7p8OvTO48KUofCuTff64tGVvvOW1NzyhJhnm/NZaOXGxAIxcN1
EcUHtQqznPdJmC0IUkA5cJs7Forl9xH4/71dZ4PMTpFoJFTgFCQzyUm9MZYF
1EnMXp1FMZwzPmOOfeiDahK1aTqaqohJtKVqYeqkKm5WJb9WM4NIgGMR0dCF
DPb1TBmQIBuvwh4/SQe137F42x4uU7orCoCKL18RElpWAw57B/5hJQv7asQQ
aPm3Vcqk8/aLc3HMFo1Kq76tJBRUIVgx1KDPFBJPkLwPS8ODwnbNv+ZfbIoD
eV8yy/MJPm6vyDMNA8MfGHXzFr/7W+FMTQZ2EXSYAST95fC44KXEAoJR8+4e
UGLZw+ctJb9wNofLnmzwxdrjg3Z0lhBoBABzyVmlp4ULv4JFAP9QKUhbsNS8
EXBKvORgFxF997zytOWuzsc7SqF720n6KgsXcSUAtxgeTCFYgGPekrWfdEi8
M0rwr5pzULznVPFO/e3p1Paq7AYQXG+v2oJBQmieNkWU3UqllLJ+usd//8bH
bm5spW4B02HXEwlEtolXNkWSMopk9/NPLgpftSSsL1xXFqezdMbHbPUTjxGS
0dplTDoyQUXs4K3rKljEDhuwNv6xm77BDmxKQiR/SLEb+p4fnZjtViZkPUal
9dy96clSbviJ0IjIPlTq5GmLAHlPZrKkjeVOeBALEtpFZat78N0kCI6qoIN4
sbOkySZqC/fsDF/2iE2n6XvF3EDWflTmXqHNxdBFwkfLo5/5Arf8Sqc0zFDg
VLjk4S86zqJyYHnDsHsQGu5yDY9M6GdNQW94K1g2NQYRjcyDAvRP7AeJjWN+
Vtm4Wjf+MW6u1tM1qk0AzDFsFLGpKS4HvgzQkhaEgotbi/0srzgpFYWjIVRX
eKAmtRHGFF+6B9IOK4odVUUbMkyoQtCMKRjaN9vXBrQ+uikVp0oopACsEZRg
yIEX3fqGiO0njE3vb6q99ZhOjQqBq/Sxf2UAsF+jQ+Q7gaREKhCSrYZ3kSMf
STHCwamO37MdC+B4cZfx0H/MTU3QEW90GXkOyXY/pFp9sZ4eM6J30abyzpMA
u40aPF/DzWl73pCU68+LHvfyQ5SJxNBu5/i4pOqFyFoWfsy6jjJIv3bMHb0i
J7RnSauGAuvUyNpCE+C/wLU1Sbe5HToyzFbWRQa5guBsecmz7uOd1HP4NvAq
XHStINV+ZmFdeeUAXx77IQDsSbHikfIgLdZ3FXlwYjjz5txmChHDwzsQQjsj
IFGo6HdsoMgLmra5Q3zmCDU2bSztIwMmIG2sHLLqpj1BkT7m55+5fIIWrbzZ
mvZOu0VW730LYLvAUunTIVecRzYf5ybhbhVqqnvuMOnDnG1isGg+fz3qb2bW
506Xzha5bRx6lwcK0wY+Wa2nCPdErsWlh+J26r9DUQOxGPhynLPna6DuG3lG
93K+knmTFZSugTwqrDvLe2DQ1s74qyL2hywGp4qQbaJV//3DKC+vnZSL/U+u
O0eQUyK42/C8GsaYgFVtwXrhmh9TXRJF29aOHp4NW7CL1/0hUmofxblaslxO
NMQGCuCluHWG+ud1H77h07pF89eEWZTRXkffuJ/VjnY+dt+ST+/hPgZsRWsN
KKvgKE9uwpAsidLXML0WysvfvX8CetX9OOFpIDy9VJbZqLW6Qmv7M0BcPtOw
+BKALO17b5fPeT6FdDk1emfqdXcYsQIbKZqGjS3G/94vRx+0y+NPLEGEkk1q
0pIuCE2MChF8LUsJpID+qVmduU3mH2Laui1VPE4Mr0QlDea8UkahcWnfvjYQ
Uy/flXrjTEs/wntw/2m5r9/ByTOZebgUFS6GCoRS2qo1mwXHTNf3Z2U9/Kus
gumUFY27gPO4SpeAFD8kBTJZlnvBKJIOhF5kT1VOKqORlbkTyGm64tf0J/5g
utzBXhXSUvBCUtEYPy5NyxkC5SJ3aQ6rc6bH/i62AhLTETesnODOoR81+Vuw
yeEsL7p3x7I+c7oSBTgiM9dafL+K4rrlbpwMNR7+pSLdJPP0+vjhfE3W2OTs
WVm0qXdlbnw537wMTeGtGK8UbhPwCJ9MQrHBkRxEJ0LWBkhp0sEFQP/4D1LL
wbhTAbnfe6trpLF1ZgbYL6cdcaX2byq42b94o8zRpV6JEp2dvEwBo714faLB
KPuVq58G86tpzybvkChiSpeWdZasXfP8yiqdTgpPvy9OoF5esazvTL3bs9fR
9ss7RcIraL3TsPHefyRxM+fDA52ypVqSgoA4rQeyFQn7bF851K3HuJkDOH3k
BJjZms7/icjCki3aquJzsSgITuteiSzwQNH9pbuL2DMNFyKIQO6UQ62KbGQz
0UiF5jF5jmL6kx7vBPivSOQ1nEnL3Oc2QaUXRyKg9nHZdmNxsJjOvvMpeEFM
cTuvvJsQPQjegJf+caCKiAzFmiXreucEGFIUqggsGdZ4GXnVhPdvPle4qtMh
IvtP7Spml98rqCfJRgoXdFk1qCxly4MNIwcgMzPuFz0pCxrESN6e6B+5eHDp
fbxV3TeOEh28Qpe/XmY1GNdGbslZL+dbnC6rQ4lLBxwcDH3JYXrifAUQLI7k
AjKlXilzI1cTdLjfoR6nxwtl8/sTZFevnKn+XEyYjjBMcR53O9Y9gV/l5WDO
xhSAEXetHTiwHqYQo22EHR81hIi8CFWLbarwJhtiZO6nl5g6TUxWpIeeD6As
kYrsn8EMYdJ34tIZoXTxNqrVLMmxzMEDrL7EpFn+fTlPTCM5B9GWH363tbcR
ooNuaOm6+hzdnMreKoIYFvJmO4WnDsDDHbm8Z6eDPerRG5oF0Zs8uiIm92l5
Eo3rLCqjM0AHDFl+UmtHePN37nOR8AOgJ+IYs5tYfhI/GqppnFyDCxRs4g9z
ko2leZ5K+HNdvbZrueArnedGoXt6cxw7POem7QAjfyl5kas53lCinv+WVxgW
oGyYeJb5iKiqJl1F9c/jB7zcFxgGz+vfleJu6t3AIobeccZEb/Gei0s/uxvz
c95Xem6NvqfZvqyRY0p0Rzg49ufWzdNCXiDxYbyGdSZnypQ4OfHLqeDxuSNd
Vyl9jpQwFjvMxRyCHmJthC077OdL60fOxBGbX2GYK9OLpqpOa63sGUFoSbNa
ksGyhZKVM58SFs+zWfMkBYVayUzz0a9di+YUSAZdOvvb8TmbzBLTQn0FNuem
80tnM8vKFXpw7BAPNsjMjQ3UdGHrHEtkEDCVDtaDyh9kpu6ihOygBkPHvjpf
F2nPALiKmi9tljbqyFcDSnyAxTgExr0bjwcylWMTncDxUXdarK59CHNIKxfy
oXuASmv3xOKYOILWXdyDBvlr2yATFq0tnkc3lsgQUmysmEsNj0w+YZ1/tQux
NogyeiNXFcRBt4Xlx8lS38pVJiy4JWTbzrU0a0ZRh0fu1WY0Ih17SdZwUC86
XP87xjX2RMUPtAUHvFsRXsCBObm7H59dsw8U/IN0TcL1dNp+3syoUm3EVRuD
BRycK3eFU7huQ/NFBmZSLjz7Z5WRpNt4rsYL5Wyqfyn08h6SiEail7gwpiCw
y7vp70gDo878Lux7RvJQPWiU0zgUBStbHfJtQfJP1YsUf/yFRG1oEnlxn6EC
k2dhxoufbdEANafpM7WKf97RrOeidqH20m4CHkhtFmGXNe1CjBmloYdgZnUO
SW8Vec2behW6Stk/q9kf17XgdX2Inh4q3Jd5CmucMq9/aKk/GSqER2esVM+3
RBBnLoGPmsMrI7K2r1xHyYiCgGYd3n92LllHJBj3Pap8fGrieW4cdqoD6p81
8ON8BysAfPAYJhcDfEzzGxoapKhgH3EB7sg6Kg9bKG6LEL2hNVGrQlRpGVtm
/v6CoCQEG8x9C7hHFXt73g9XKWEEJEzxBc841rr3zyZetHof1Gls6pbNo1u3
UiNTurdDroF4VkC8vK6XkqSVMwbMdAyAv2/p4bjUVmEjRQa1ioMBE9ZTVne8
bLRq6Ju8l/U0IwRVkeKi78I3osS0OH7Sj93eS7picy5n2qZGSeGZN/sqT9I/
SLEjjZDZFlNCa62swiewwxOZzMvmLSZi7iMtOTY9DlPajoNTWjnwXKL2a93x
QgA/p/ggmtYm/4OUxvHgwOwjzU6DUX99gvMzWVJLJXaHT/OCwadM2/1JQuDw
RLCi6Qtc2T6tV0uHSPefufDi5BCbhcAGUv1bbDXvagYqKR76+M4/oKkiNDdd
dRQz1L1A+OLdbTalDfk5Xhh2f8Cxp0EjVe577bxOCCbnZpmWmp59GvjW9rjI
7Ncrm3tID6mmxliydz3nFhmNOTNdOvoE6cs0OWJEsKkrs0k4N7ETysWo5ud3
aQu2uuHZ2de9jGcESTysdjOtDCgY0t7mQwwlJnR6vjQuyM8Qb2i0CgmJ6jmy
CpZXRKUocIdXz3GkN7UbwGYgeSbXze1g7ZR2Bwy5gL8MlpF1wqaaQvS1D9Lr
38Szv/VW5nS+qCMu3PxAszrwIc+B4ti/99wBDsxmhVjPlkKiOq74UGXvjvf2
gh4BUyytDs/LFn9eApr8o8EtzICBx4AF5R+acu0g73yXQdWVygA+3MQhJPDd
tum8swLiD9NVEvekUKI9l0V/F9apmfm3qTJrI09K+w5+eqSRtPcRnKv2+M4N
WXgI8NdxGMRhYkwYRnhDhuZWqA7mD70jYo0vos4/Dcgm5VBWL/l4zERU5MYn
rGICD3Q3wzxIOlG7swV/APqEI5fF6XOQk6u38oLa7qGgWVUUS4mQYhoOBGXZ
iXNEHg5ypUxnXW+uaSSZWI0fdyNouX3Nw2oRkpq02DovjZL8RnphjnE6dGZ5
0UASUGMV6dmRFPLeU+Kg59Cl65E/dkGJlKsBXIKy3tVA71BLhHJ6BhSm1bRn
W4lFOqn6XR48K2JiVQxPBVx67XW6jkEnmnd0OGsIaB7ECifrgBn7fqlsdBuZ
49Bdoki1ghjqrnX6wc2iy4eOfknT81LtWdU8B4VR7+kfo2QC/plW0rg0Iukv
rUYCQRT7F7Lm+wFPMVW6PmwNlEmHIR0BGS1m03rUeDvZRo99hWANuVdQ6p85
xtq7YpGsCu6kGHZftj7JcGU9bRdlLhTPyAaxZrYThM4qvX03DOKViCZhfThj
4z6v/9DRmvexIDuMx+xGar4OqmNIyc4Ud4DLEPxNip0GkXsDYlLuwyFUD2xi
/ciuvDO3qB+askTFDVCrUpwIDwZtEX7CwZKz8kHE/jRTKCcwCnToFlN+TLGO
x8f+usp2Jg6PJTuXRF5RWT+aWVQw2Peo8z3LNBf/e14d1tcVjfDkrYC4ICM6
wnzpdgwRVW9xbul2Uzak1b+jrV7Tft196o2g4REfwyf46E+WLT5gKjhpa8hK
OAJHVG/G48kPNzZXdaKznu4iZby7Zem+2M1eRbWh93TGkwGxjoektpm38HO3
3OLtxoRLBB54JVuYnqR0mVaIM+5vX4+81c32jyI7ooQQJ6vHzECynK1R+e4/
MPnjdTG5LvQqKYLtLhb7ugD75chq8/ZX61nCcx25BENrFDc7DwErgqhcvPZL
ZMty0uSj/x1K/D/p7ZOEvl/Ulg8WvBP2CuRi0vxvm0PszG4cNhDvgTWuj5Bh
A5KneZfZv7fMXZhmXBvhnWjWGHZPrzrUiFK3aQEeNH24VC/ecQLEV6uNBs0J
pD4m4hSWSp3mKASsrO3k0cxYKqnYGgmUnJTqmLFBT5qAfz0COo4x/I67QCtt
UeacNiUXl4a0wOB9PMAQZX9y9xw1Nwu0fhMn3duIVFwL1QCi+bGvqKU5jxf/
h5qqDCGahIMEhyVTa/Mh+mhrLgq8BVm5+7uu3YOtUpxA3+qSXnOdxpH1UY3O
B8ZQSMkqW2HVO2kcwiotN917AGJ6VlFPcI2ZaDCAsxsj76iIW73nOdTrJE9+
bDf8wwbYUwf7V3fOSPS82Gj8RrL53asIF526Kqi/NciO6Lq1oSXyKOWr8T+M
NZd7VVU4p96aPlUo5HS/S1ouX4Hsu22X97RYQWLaNn4ubYB85+iWDOnqsUaY
YN6h26K4xb/kXOzVrBINcJ6Sy7GLhycIjoWKzVi4J25Fwr6+xd1GWjL3ljDV
4bW3kLWOouB3lL0kH6kJjHB6k2qY/ltsi5ykdNsp2xeNTgNz1by+Hb6HXNdz
WdvQWKaGjZSHZ/6tI2AsSJb5rJmHaAH6LrmbTfYSw+GEcFVsT1ADrr17ixZZ
UbaUnl9O3N8jd/EeSlMGkj+oYeEuWqrh8aNloSVH8NZBjlvCZ7RQxglEqlNj
alfT2we7L+sFC1jT9zAnE96wxuKjmcSxh2oEat9eQOPZ8rKIGd3HEb+UVaD9
CJDmduE7wuxtgvSpBtIzZ4oCNvjmPX0JuT9uZ78SOQCCrh9gSY1+4wTMbdeR
CteBvmD10WNLgiC9TIhHKoBR71vH7ZpKx+GiU+VGHkrAdeX7ggjDAsrINT2y
jTPv4UdPjLJy3mIZIU36KaFMp1JBmWjhNHUTcir9wcHLlEa4gcC257PBFtTh
Mp++ixqjCXgL7j6A/oT1awJsSUjyMTcX3/JbdcPF5FiUGhAevINbS4EKFUpn
L8PjCoIb6WJDEBwX6Aep9MY+VF58VY9UFibjIhbYCDUKifLom+cZSOddWewt
7OZ1Uz5NKBWuhSCYJdylDR+MwQdCUQbBNz9HV4JqAotX5Pl7g+K8bR45QaXn
hLxvurVchDl/mDBkP7UfLPUTQ4VDj4jUbWHoltmW8pVhBIdYT1w01RAsjZ2o
/xDwQh2tLHIUWZePXVG/quC0fi3ywN50wZmqaSqqPyiWTCWRF/h2I4bBAn24
5KQXw5VVGpooYaO4yKuaqP6mRI7aLL+7YIfgRMkS6qCK5GdKzmQTynEbcibi
uK+YEvUazhJf/h/uyUbxLP83/QlPzU48pWj0dUwu+pr4e9BUjqQEwIbPT5Lb
872PnmBrUE+eYOdJBFt+2yRg/6pkUSollRgghogC0sX4qsKzuwMFae9rL9Iw
94l49UQ3czBJuyBqw4Xv4Vw3C5SEeSmfWBYi0l/3gRNqzI7apcGVMu7X3jfR
RgUMZFXOCtmq3d9Ez65Y+8y8uAh/xgtQ2iw9L/QnCrYNF4Tiwjt+9KaeQeh5
I8o+JHjlxXNOe+zPWUr3eRoyFxne885ENK3P3YBufo252cugQI84MCBWzbiX
R+6hJkx05iZij9xG/SfAn3MzcyaV0FnkdDm/7MuZAehMy7OfO5sj2XK11vrK
RM20koBojHjyP54iEbVnc49DzcIccPj/VKFYE0rhwceFpnuFYZTYqLghLrr7
KMyZ4CFCoWvGcEYBXAlzbHSvPFzMyDWLwJ0KklVpn8k0ERMLbSX5uCBPFv9m
LZ3iKWvafMC8l+OJGwhM8CbEC2CsYS7JoYiDbbtm2W6hpYopeNaag/vEIh0Q
JpMZqfpNF9ywZ/y+jz6Jg9aI8bswLLuK0qHPxZgkfiIqCDnQuOn+EEKJSCuQ
8sIiAjVBvdXwgwxOwJWSVLsLuWNA2k7FOA9eRnW2txb7p+2iB6kDMlBZkeZp
On6WfMW4CCdZ/gYXHT1q42RzcTj5DqX9ykwt/z/7zL9j5NpDiyLKwuuLaryB
dTAOWi0GMbWidtieBxnkEK7MA07QD5XHgbAvgs05JFMH31rCzXsGpOM0zjam
s35OBd1voBQVzbSI3VSxpY87P+qcMJIeeA5hvvLJMoREZ1sRnNHyExaPwmNh
dzT2S77fe3tbZUnD5mZ6h2at9YWVAwKAwXC01Cb4wM+q60C9/nqTSdiqGdAk
2J4BEmDLmihzRpuLatbQNLWwHl4KPXR4eeolGQDn9JvHQCSik9aLX5ZWKYur
91aajwmu0poMLp63Mi7VBtmlXIHVUc6uqeyQxBbFdPtvu8fPqCbjAWwZszn1
r+FGjPZOK5LgKUnDCpbqbGiwEUG9wb8mvS1i72Q1DyOm/w5NEicnxi3FSJ+H
WtYoBFEAOziRkNsb1blLMF7c3prsBKDUv/2cPe11GcSaT60H3UJkFlDDP5Z/
5AXgAwJt2DvXZbzrfpoBFAHTJWI5LwH7s56jJQmo8qcaKh/x7BV+X269z2UZ
wBu8F8Ypp/Kukof/B/N+HzwFrjGf3gKVk8frzoN2kX1C9GDGAIAB+1WR1ywK
xuzLFe5VpLpAlbVgLLyxsQQs+CYHoHccsI1rcf40oWDNA7/iisl4c+fqO8BA
pZ+og3Hv28PCIeNwPYlTGnAuCDZb3xB4eW7qtodKOOnS7jwF+1Le09pTsVA5
2uAMFyf5RSiEs9LF/YTr5X+U8SGrp99CT11bAanLaSnXya1gJfclykGWRdA2
OV8ki24dxdbQCPbD/jkEn4ThLa57VJbme/jUQ/sehOew7yqtnVSFD/lsAVni
k4A4S1TOov0+psVDHFWq/liyMCBTg20K6LEoYVW5pOuQAnN8T8lAQ2yibMc/
2redxPEFAUrEM/oVA5E13L13FidFW9eNtfw5mzNaIhOJPGb8aRLRLV5MDMj0
T6mP6s9cpAzzpOuXRTvFNEVhwp0rq+eF+8p+KmP6HZO89HzMdM4ISZmL1jYQ
hXbfHz9KnZP5CMcT9EgEL7dOmmK8LpSJYbyLxcCxygF7POdDtZzdzuXhwTQ+
/ap82y85txQI1I1hOuvQfpGyhudWyeCqE/3BFnuhsNTZ+AzhoDv6PKWrZrHQ
ej4zUXqB45m+TnHo5VVKUyQ+NXyjGCmZBLADfvyq+kGzDpaUN15LHGruN5CZ
kKoUgiYl9NDiTnq0f1jE19784eHvfKgJu50pKKO13HlLYoKG7hBxPWg9LgsB
AIc+xB5Z9+T8EDbOpgS4vgTxBg39GPMFf9iDX916gciKVF2fezJpsPG25wtA
TYCgl/UlXTTQD9QaxvFUx40Q/R0asHGDefVsxVnHVfTku7Nw1fk3jUqwcd8D
3N1N7fXDf69KQBMS2328GlhSFCyW9GeZ/Sjr7PmshRLlAMczomxMv44fipte
o7YF+lC0yS7kcyD0eOy2o/9PAdgE0lmxc/m+YYwGsXE2UfU/530E8hSv5U3i
IwiRnaEKk3IwJ6NchwGUVNModNgY9yDM61bahoSF2BzmnB1tJi3erW7CyHhd
tLYR9+k51C+43jwW0DL4odYBlD/NDAHDmBnRJ5AvOT9eSfbGbgdXBzIel6nV
Vbg75h8Uo64gNWTDVWh162tKsXmUTMwuZrp971X6xVGT62sOTa3ha+m/S1AQ
IEXBvogxYav6khhIdx+H9wcfZU1NVMaWB0C5SvxVpbYM2bgf3KYJ/bBUry5Y
JySToKtbQr0NBvUJEjXtrQRMrHDdoVXpqKjFf9ZRbWGiPnBRRuSyPw7e84qK
Sux39TqkHF/mDlIukE6hgEl5hDy6pQTlIZto+41gy1d0egFoIjQtnYcx+rQG
gL7hZ8Jg/lFvEEgEjZM1npOEupaEg5Wc3W8wqh1cW+oQ8SsC8QFEvzzWiLhA
m2VaCthnC3DE73acLu1SG4qFyNDmZcGYhf6f1OzkPM20Ibb4wNubBOQU+3MO
XgzdEydl/VCCVoWqD9RNX5mxHCbNa3kr3W+0dU+Sh87B+MPL3vviMJ2rYuTy
PYwA2Dhdi7AYMo9c3IQsdnVoGKPIeSKDv30xbzqYs2QdrMRJyZ1R5Rz+LGSy
agNO8aYWwrPJBnbrldjpfC78MfounyGD6JuekSniL5A2rKp/gHbRGukguVbU
jyk45wOuucNPv881TweWh91xTLINeE5KkhrnsJbWpjnak0hsAN5h8WjdfVxn
c83QEpvaGjSVQkW5NiZadia+z5Vxhe45cUuWlnQ/9yj+ImdWHaGjqAB+SKFV
s7qSXZpE9csw6qtyQdVCWbVl5xPFWQ9jb82Baxp8w+prt30aB3t8SAt7LJa3
BEBA4tMcXNcbOGwe51oqfDG5BS4F2iZFWMTFu1zDubHoaW/tkkxflsYYZFs0
kw3nneXQFwQgZ/X7j/btOhkVTjUEdz926L3tcWcPsFMmhHvTCfw8z3Gaj3DX
YpCG9432RgLdjuEUDgAWOJ1RoC13dGmWNku+YeJ8IV3j6cE7FYcVbE9QBLDQ
FoO64TeQDCIqN888EZitfZZ+FbhdWKK2nyDsLusWagxvbuBt0xtl6/KbBcO3
+4IjMhmpz8aoY8qraXZWkMj8pOKPIFwt11kxe3FER1crLAGp9kPuohhJauGy
2NrXCgh8TXu0q38t/wIx0qUQd8Y9YX0OkFy40nbE5GcvjenTwOzkUCNViQQg
S2SX/2ps+xqlGgZW04SoaCoitgP0bxkVpseB8vsFJ1vwLrHA34ICpzSEPkVq
ta4//1UbMncS/IRD+kx9lOyBEv6xuJsJOcJ0jcJabqzYUtBy30zTArZ/605F
TfoxZT6dAgvu+pDYcN1dUHfvF4bQIHds+H75Tp1gSMGAJjuCZVhtmDMkiV6I
jTuzOTWzVYUHeMkQM6m2H1hrFDJnvupDWHZx3Lcqkg/TlgWcaGNfOAvAaQur
HSHZHESSM8oan76++v66QSgmN6wDRRaRUbBpBFeytYy6pz4oVQgYf7JrxCLd
78rY9RDUdH/dncgfcai28oWAP5Cdj4d2ibBxiWw8HihElVlgpk+TAk9vmDHq
4bHOcmqMZ0r27802nYz3A2fnJ8vdqBM3PqIAnVNFmX8ReyjfgLZHySBzuE+D
vlhaTL8gErXj11qwLswUEwp10XGu3J5Y94TbRhjaSnsijE/ELnspcJTBIg0X
/NxMqT2224m+RGi9gXg/xeyzZauObf3XPwnBavD0CAi9Pb6PsQgLHNQ2F2kG
8UfDlIeL2kN0i4IdJ6KSnRz0CXj2qS/ll+pN7r7u4+N4CWERwS5mMs1cs85Q
MSu8xCKUMCdxRAFzItO4EfShGDrjkKM6ZMyfpfie0IDp1BtF3cupp/qqiE0l
M9FujlRF+u9p8V5KBpbkvXnJRNDFQ6aukgloC4lW60CcWwPgfxJs65cb7j0s
pHIN/Gnkz3h50mGzZxjNNpT+3oukHnL333JpXbS97e7E7RAnpBviJQ4jtQ5j
HVvBFF12jiAKIrHB4kNhXQMEHDC1tR0oCJ9e7CJLp0o6JcijX5wckVwbvVhs
g7jrDDYgn2XCCoIOqzvAoYI6ms6gJ+a41DXtELBXhyhkn1RyJNlRFSAxsrmv
n8Gz5jsYp+o1fRU0RvcmbD8ZQQdRkZXVTVoULbdOyX5SEhnKA8X3tGU/kbnD
HSlILucaALrR3L/cRUigWp9stDhZ2M6fxeH7SuFjT7v7Rw9v1dOnnzNHyjt1
t88Td56TWTFYcld3z86H7c8J/7OrPfc+Gk9MGeJzsi1szbkqD8u0JzcdaaIB
kXeQd93+HVbdU9N7BRd4QUq64mCUQA1DZ4gbvbI66Lkx4lIQIHwW/26gz3dg
krsULPLWnFXKSiTO4AwdFScG9pUeD04RjMDGcAJvZPIdEEzhpLjiUb7MQ9We
7qXxqW43JTrLyA3LZdoroxR7poD2pEI+IH9woYCs20dhMjBrkOMPN8vPBEzU
hyw5D8a8KEfPeyl06Z7ARMpjEA7C+dvihujIYn0HST2QJIyoXuPwhkCyMHZL
32Ib96aGkGzZlOhvAkzdIDfoPj5nc81indThgHQVC/sPrTjHGsvzalvIg37I
exBLAwvU9UdqEXlNhYVrREgwNXqn23OW0aGrukN47IzSAIMkRk67g6+TGJPu
PKIDbcgcmDO0Cg4YOT9ZqFMssVZgY8jB5w55ukcKl6XFozvM2RSh5n7lAXSn
SzL7jWvVEwKDnjEm5BjtS67Qf78yh4M5zRgebqnv+xKdqze5Nxvw+ebKBHRO
J//mCbyp4TYODqdsytVebnKQYRR0cJy9YfVhe57/DRTk8WrWuA1YfmLUERdY
x5FIFOhQtl4F85qeqiDlF4367rIxzLkPs6qIIc8Vm/KS3w6iI4Cyc0OO2qDr
dz4xx0i2u6qS/UvaOEyGjwAd9T95wSf9Mi3r+RKzf72+E1XMHjsEC6hY0JWp
8ngrujDcMihp9NcV0ElhMSVUdWx67LyLAlqlFI/OgtwKoM6Cvwq44X92WpO/
0ozuHyfN1NPEziBNA2PPnIhuOIE9c/K7k19WxWZqMfs8/rkF+YkEqoe8h9QE
XYAqpGyCNku0zJj6Ud/P5RY4yiyunXCtCpMi1QPk3spI3viFleFQGDolY7sV
RE1P18Gb2S3B0fGCDdU7dxg7hmHC658kUK7BydmSQKbgDS+RcCQsRvpS39u5
68aa4eFQNfhgsq6x0+62SzKd7Z49Xgd5lXqbPf/tHRYPfglwz2YltnrQcesp
0jQVgSdLvd+nKgcSW4IpSmE4Zljon53iFdvbC7azvi+Q4jFgFYfQPJGUO+oz
u29A00SCTymODFbp6Tft5s2SpmDx9ACjAvZEoJZL2YIeSDoevmL+L5W51i4F
KUvboOqEO/PlNC7n/yuG/9JkiOTgc2wzxRY8MhtAklzU2A4by2alphRAPDZx
pTvDRTzuYYQFZ9I3YsHeNqLwiP3k2TrgxLicFJI3Ct9eUMOGhmrTF5fJSqQz
wug3TiiQ87QwYge/Wa0nKLMSvw+c7KdtdgNQ0knLBloT5BYkEgD00/3jRL1e
y8w6Wjt99xQ8908wVqZ5qpWo+nU4rfizheqcMGO2lUQn0KKS0Y0q2hb076sN
yNFtzhcn9018YPa/pvKjfrVzxkIl+7lxEhQhBxQ3yRKw/Wqw8lvjahJtJs8H
Np31UULbjtzSGnkT0XKadcjj223lRZ0Sy95Nm6J2dyl12aZO9RgnKrYMzWut
/nCi0Jq5SXDwLIJo+Td3/VGnm77Q9vKhLmvGBW186fizk/xAC04+LOBaGoBA
k00r3ajFRyxLdVl5czW60lbgFtB8mS+dI1rma/DEaY4T61n1WvFNRAxhsY+j
ddyGcRP9Enl7PyctlqcHm+l89tiYOHeDQOShqtKAnadbg2lqmftQ8qNWUYFZ
XdPSi4K+X9ldGGe8ER4hCGT8z6EathQ+segQ4BnRcSnyzDzd+qh/rJJwXH6Q
NdwdLZbkWUTN0z+JIFLGP9mZVJUZXvilGAwrrU5WoyK1THxPWCZTAcLoODU2
ja2PnlR1Bwm3N6v9dXgU//qGNj1zLNEqYYHbg5/t06yV5cNKRP6FFVZP3NiA
2wUK3YdKZUoeS/PKLXfyMm46B6RHf5MPqx/UteCcAudYyo+a2ktHlW0/t1nl
+BplbRg2tDSjUmQV5yNOHeLwKTm85Yl2+9gzeQ5DbgDCpEhE44qrO/PO57Lf
tWEB7xOgdvsv9ZIj68uwqhhxc2xdM5AEhBkKGhliJuCBRTCw3qD/VOSQ8kUN
dgfxmzQqQG6QRP73iidt05vCh+U4HDBMsxcU6MPb6odaL52o14TRXraEO7le
sdVZ7uu8dNt0arznZON4LR2aaq7q8wfDKEu73joFBjtV2LhxZ5v3reCFb5em
o+IewM/IAIhwXnhdGZVGQ8CRQd9tnII2izqakQpiovGkCT32MpmrQBNWr0WJ
PSd4H8NMhWa9HD5vWtVb8yytz5l9tJ/mJsoG2ehJ2fepvV8v0Z3TEztAqOXH
o6HqDtC4cEGojcpQQw3PiumwxUI3Wzoroj+kiExlo8a9YMSV6kbZfAktty8S
VKB6GYGRaZdii3y4zvyI9y+jJ/pB0X3crn3ck1Kqqm1y3P8G7Qhg0Vl8PxPU
Mawc+y3MBlJNu9xes5X8A0EJn/xqaBaNCl+SSZpuBrVBmzvy015UQSrbPwf3
AuBvNboIDs9Dm4udVdcqL0rd4Wmy3SF7wxnYwvoKFkxRNNSzja8sRj6/tRf/
uCo9FChcDzbs1lFzM851TGWbAxlje7CtGQSEl18usMTuVm53rfm5kPk+L6VI
HDGXoIjhLlCNE0aMsmn5rXGcR6BIADrBzRAKAy3mTQ2noiPcKVaGhYf/npvZ
4Q7A9m7/kMJA89kW7i+PfShmeQHjwQqCOjcdQaiFKC2H6IXqRsEt+ERBeHIR
+H8Epe+8zy0ywxthGs26e7wPcNqrGSRB3nkf9jIwfID2Z8rWaY49JzmI3+rX
W4Z0N1V9LlxGxvpsDPDx/xERDCnXmQKqxyjiNdIeQlD5qXaDFT+B57CifLPk
sZjmKwCoxQqitZXdzjmnZxVg2eun4mH4F4sBsIcykIfC/2J+zAqIEx8Jic1H
1+13pI5isNUsxmQiGH7+97dK+MaKW+4BRcX+TZTJ+rFSwEuKlCvk6oSyTL+E
6aflpY6GhJOmmrqzdbqLSaoruElPPQN7bRGI4tWbvk3f/bleljYCRHT3QeQ5
ENHxnCOvOYbG1qwhEDq3J/cGgI7N51pU3XdAN3VRCxPbqSNxvkNDrXsSm+cF
9Sr47c2gFn37J4L02NpX/2MD6nOLscQiyAkY+B5cnekJVTkXj48dN9BKA/tu
b/cBG7kTQHJH4puva/S8Hf+btWL5TbxrikJNO7YssBC2Q1Y3p9Sro0gDGamE
3x+Jz3nXrs1Ivhh/2h0Av9H9278MXkczOaMvc5eG7eozxfAmup50Aedq2NZR
NsGcz1ER01aNZyCjYwHJVfUfNuVSIanTDEXiCoX7uVk00SDJwEpLGQ9u12R5
gShvHwEKaETNR6tyRiY5TEu5LygSJG19RDz8sLSB9H4RVE57W2z9KdsTewAw
/lgVfLKC09NlTOHqX9K/8jYLt/Cze6bLFt6HndVZf6Q3v4+oOLy4lNFQs6+h
xsmDERajZKGSX/E6v4SFJ3fdKKrZt6o/2voifxMNfyfVwz6WEEYTDMHm2NOT
6FUoOsfPwkJgbUCqYaMeWd0OaC8hx0iK2h4O2NuIrPoSS6jCL+OWf7qSSZP4
dHKpg5ckGg4AZQAkSdbI4ujo/LCRPKIJ3LjBovx/GGKYY/dwO8pmqBWT31gY
qBlM+v8eEZNDkdPao1wRkwcfPbljriMhP6DbpEmiJwxgmU1W07xRAXX84vrR
k2BA2IJaXAMjBvKc5r+AhFgh6UudOdxqyDsL3CEh9JIDXKWSI3ey93EKc3Ry
0jZiXa92Z9xt9dg9HDIXOM8flaeOqch2HKEtotqYI7+copTa0u/1+Z8dgyyy
leczv/dSwmckXatgKizPBpJFI+2RL5CU2DBYQunr79M0JtyGKHGvmoaxmkXE
sLdEYZUqbyiFH6+IJiKcmPzemfGPLoUVwAVhcEIuWwhQsGdvM53oK0HyGEGX
PgGYbnEIBxz9/xOAvxcvAeYLGaSfILC//jprQUMYFCvxc3fAaBD7v0IlvhhJ
VvQPaVsQKGkrXEZkynBTpofq97haDQzBTXl4QBRRFaehGr7B8ehLBHXzH/12
mpDBIexNwnnARdqcLjr+xnZsL1N7GnsFdS5NFgH+1zEEpVeCqbojO/wpFah4
3YXiKBLrVN0etRInCsphKxuj1tbKjSm1XCTMMH85VRV4Pae5qx8HlC/bwgCv
XZuC81nvEobauH063U0yJD2gJffGekPx//5h8XDMtTuygpRZ2me7qgMfIt7r
TSL5CgJm7Os2kInDAJCkgL/QC3TSsPh1HaVnDC1rGg7QQUyg8mE7MLc0ViOW
2XlHso1A4MeR1eCyK9pJr5j7qAY9MYq3dmB2ZdW0uUq6ZRSszUGNLOg1DoUq
I8Zgo58FXNulT4TU15YuipaiWD+WuRrlV1NYycBR1dAfQg2t3e3a26oDGjLd
4Kfy/uaEs3C1SUXi08aOBC3QONAR/g3bkYGbr/jmj+Yxs5eowcVpOdrHHe8h
p/X/0wj+QBhSm6t7Jk/nu9En4xk8vrr+Lsg9ebuKqC8yLO/PUvRqUEiBDN3O
VTTj41ehsl83N9cpZF8ymBd3F7n4gB1he38dzcQU6V77WOOlagZNWzCkQWO9
lQa//h0lfOCSIX7jGrkAmhLinsgeMMMwRnvMbEIWwPQn9BnFlWOWZjEB592G
3XKGAZuEhK4gQvgVzJXGBRu0RUl5VKjzNyjQibYaQ2du1QdbpKshE7IjzMMT
k/WdmNRSURws+ffGhG9ikeemFOZF+YhqjNd1CkML47mXIx8JSOHQcsYnas3P
Dx7QYKA2QLgJ3GdOgN1P5e9HrBzBv2O6GtxIq59GrFRo6a2xuyogBtBhvIMJ
L3Bq8WDbB/Oh9arMLkDBS61JoxMsZW8IeM2qY98aQQTm5yjswD5Fhbuez/HM
uzyOAYNGMeQLgzah4I0PRQrZ9CBQ6zk4uTbvSFlmZoGnkDbAMeh3DqOAi+hN
bWt35ittKN0UqI0ZbnDD0ErsUCySUW4v9uiXptm9hRPpGGjE3x0pHXMEekXo
dONRW1xsGXrfHXXwXqakR5GM/aMbxi9NViDnagWKrtFvIB/ZxUw3jcek7msG
Pq6ozvMcUP6sjhztfkpSApwqTvX9uIu9Sq3wfPPj9YlEDgHWQdkWMPZpLy+B
EfwkQE+S88+esPu9GTX+zt70YHHs0BM/geEcaGugPe78Zt1T/09ur7DPF3mb
4eWKH7LnDbzcJ1wF/Do5cA3QwC2JM8CBOvbefMxYcYvxYsmSm17tUIgclaIy
QR+EHHXvzaUhQm4o+xVhbS/dgkjB9YApU7qTaXLAusR2uCYOB0ewS6vsG2XY
4vStkJNJdg1y5xcYaFaMzXkhgQKb9Mq/icD3HdHWxBbxM6Kjmdmx3i3u6gKZ
MQWKuXzxDokbRPGnbmXOIh/2pAXBc3phUFAg9qVKrKlpTn/w+cEGl8oc4HUl
3ieuF4+r5E71ttkopKvhtUxmii6tP+zs2jDhLvfgxTP6KUsyfY8Y0EKsCCV+
f0gW39VqzV6Ca0H3plvfpfcQdBovkm/U9Bm96TnJShPhATirZ8s+GUQ20vxi
VUgL6oY2jdUgcCIwyiDFpzGyUKZuuKI2RUWHiYI6jOBFFsK4gxUVMkciYXU9
pVEbtrdMKP9XoMEaB1Y9svxKzLLQ9LR6QJ0jNBVA1+lguMet7KVsNtzwAbon
KeOOfxWK2st6Hw5uGtHbzC7NuKEGGa7ExBohoqNwrjLnzlH3XyYj3w/zuuSY
mTEXLdg0kZYoAymgOsbIZBvPLpNta8nLiKYj2lH/UQluoC03sGsSWE/DeOTt
Uf7RQxrYrU+j6bE34kpTnMjUHc8BvoutQgWtt09Z5L3/7phleP5YnAsewvk+
a0He8Xqd5obC6larj5/F5ARHru8MtvS05K0EXhrUbm5CrRblSZsdesmiY3uA
O4a5s99/yfyaKECX/Chwu5l722fw5xCggzhFw/5YnGzsNMejZDVAZbhnAZYU
bX2ynzNrrYPj+EIgbw1D0RzCPYY5k8Ybjs1iK0ltLqShdtelLXeiPesiEpzr
N/qqJ9JWXG+QqxntdJTn5YtIgriTeUhk0apFG6G+fmWfL59gdemixb6yhE61
6omgOts8r/iDILJRvzJj2pJ5HGk6lVZ1sAxH7w21XfK5axYaqNt9HS5fPZb6
xHGrEW4Ek0D0F6lNllRAb47miRjrBCDhGm/+Vcio2oRpU9KnugxCilrhrOWG
qJmuHY7q2mRWWT/XV6HQ22NwBA8MPjkiarvioGUEiOKCDU33gNCScQP/wDjL
QZFDM6/C9a5jL/CUl2ac9YaQ4audyT6z/tY2tEwe3oAAT1kOoHepmvluN/zo
fAGIFO1Lk4hLUmWtlIc8WOzuYof/eLm/Ov+XGQVdzdHdpr7n/nQClOq6YM0p
NXssVdRVsc69dX7dDGcLsNRNd3kgneSLMaYE1K1sMAIXc6pOEGX5c+4+SlRU
2kfr9t1rONRb9ckAoHYgH2nlVootYf4lKEeRmn3uVIZroiKvfWMXRQm2TgIr
qoGeGSbEMKQWjTGOmc7wvYzZv+WPnQuajMNDbotd7XK2XtitYCfqxpKYCzDh
SwRfyz62KfJDgD9QRULZ1qkZ1WFtrVvlzyRgAi0/Ek8gV5Mevh+bv8vB1tN1
7CeEojSDOmr8Qi3duwePMwMoxlWLXSFvAyGerrayMsjdwkDjG3S4IBTmNXVM
sOs5iVPbsfcvVALZTdPxhnpQ+5hBvnqNZjj3VDmAqQNsJlUSzSY6aTC7SZiA
084mdqiZyZuvrrXBwfTet13Azn0XCk9Z5JGXsJ/5dTb9Y0HJ+SE2Atp/kG5L
feDU5JOzXhRSqtjLyQ3+An2epxbST1QsOvh9cBVFcowW0k95xaJon/NiKuZj
3Bejm1jTOMZC/vL8yLdbhsubpuCmuOQDDeGCXfos46o1jqv4xT+AGAmHbsge
KKt0F/R7ZmsOPfDUNf/PblGbBtSqH31cYzcZunGBMaNcJQqVPbfniczAzY4K
zSiVO/7tCp2Xt3dQcmzmM7SXTBMwepT7eb0fqG3XDzyJJwBPOqZeleCX6YLU
zXYjayC8L3DhczwxHlBS/QFpXw0yLOITligglFda4X/QBnZhKvu6bAHSsRhj
VPGbitphuNRh7skobMvP12Em7C7JJkwCovVizFiLIi95hALwKF60Q1KbsSM1
2EzjS/fh30HdBwzPlhgSTfOPo5Zw5mDHWqB7hrsmbZt5aB2F6FhHptZIwMMq
jh6PcSidatenP9aP0cPv7FD/4QpLgt2B4JOjhJ02lIk6yMKPim4cI9hxA+Va
PS9j0e0eeg6rsSR1wyLgji5mLvTEC89NqVfCsLh4vhovVR00BQQu/5Jllhgn
km2aG02iyviujf32jb87pGH6bFeqOmnnvNE0Qg88mJHcAnCSV9PPq5RAf6yC
0ZbT/OjcpcMABdyKb7EyQw6n5Ug+kS9JryK/hvFaB1lHKDVzB4rlqbiD4t/Y
bZnLJm19SblCgr1W+Ce4ozDz98kb0GM4UCPwmshkOl7vSZavr4AZtsQhqPHK
6R1LXJ+qA8l7K8SP2HSgWrKMr6Ts3nEoXzDIjjbjx3R52x1KTs/bDzgVUi4m
4oYxdqICU7b+cN0b5p4neQNrRMsE581JUSXbeqdwXCg92snnSseZk/86ESu0
j87thUbe/vLi7UMrLjX3vah46rU12K3/YqVksZsvysTM5JIxhbvsVgrUd9u/
9yFd0OVyuAOkq4I8mPw09Kd+qeLrIamdDG5pGoT2W364DrGiClaTy2KAUVS2
QGNs7YUlYDQ79VzkTHiq4C+8M6nhfCOQNrPiXZdd52OMu/paMkLe3TjkNQyO
hPa934Qi72dfTSbU41hQVvMWWWmdtSNbvB+T6VkuyUyjEzWle3hJ0g3REjPy
zDDf7xj2bycTmNvpWFHqgbNkpKLlmqf+SgNvNibJI1SksNAX72yT2bZwSZ05
xPzWqxHcajJlwbGD7AFWGsevWSR9mStsyzXm/50KRsqpgIGhwyCEMlWqP1S+
wgMeQ0NOKcBmdIqNuKoeOwN0nEQ9W86WnfiU7Q9t8Z8ZrkmO36219Athjj8+
cEKG5SGOeNXDMOsr/BqA66x4adRDOHo5oXZMbiQt+ZCeMfjVopVpn0gJFEgo
12I4OPE8uNnnlVPtY0miYiUR+iM6J6pfS0RnC/GQs9DklMdprnyB6a+OuwNg
o1lUJhM/aNKmmIFVL1aWVJUpzgqt5DghGy5JqdpZSwHSy8UU6RftMfHKMYa/
Ke/MknW/KOuf4gO7NSSzDoPd/xsldt8Gdyo9C+PEVVSnMScEmkmuqvwbmi74
IaDsD5zAfdEcq30CDdwRHk9Yz60uzWmz0L1QlCNkCzvKvdjs1PJlW/NiufMf
8nxKDVKlp75AITCuYkHsFjevsHRI5oWhE7fiyuEonNouRDQRx0ujIua3RpvP
0VkJSqCm3H1O4d+lULm5ElH4phCR1wPM9p2BnSwewphq9/9VLAqvUOr6TsXA
/wV0bfPOe0EpJalrRfQsZmPWm6KNgPUmDToHdsk0bEUYJyCh2dkNCrWytQaY
2ZxTsbmGcECe9EVVDM+nMNvTVJ2cgRFKPXz5+e6q0DYiSGk+PFO0WCuaQFBV
XYrIhVBgNrUyEZT/myCtulYzOYO5BvB9UNi0x9vqM9EK3NerA9tZRHt0kHNt
yMpxvBKnxJfINSoZTO54u8DBBv4L0oa1/woixpnnAsxD9QYJGXus5peSTk8l
UWstGW5VtOVyRuqSz0IIwi4O9VOysUO7556Tkcky0YgNEKJACyrE5uH7ndCC
vfuVfRSkY2pIIAAuMIMO0MqJn522uTqUyCkKYLnqSb2jAO5zE/dUR3Zkk2aS
GsbUJKXebS+azLJTBBEVp7nwZ0MW/B+Ies/a/S7xj+3gvjL0aeqxtU6MGA80
zwWNZbnwJlPlmUgP04MZc/AmSCqAETHRHde7xMS10e4SrFpUsfeqSf3wEG3h
XGkC4d+hRbOh7nCfZNvAjIIv5ZG7ceeZdaT4iyQjE1gN1/HfGxLOa5K/5k5z
2YiNwdqP9u/deDwsr1sY0+E+Y6R1KT884zwCKldUT0oXMvhWng16n/Oh7gNs
3cNfT6zXhdRaptdoYSUWhfGxV4XZV082NjpwwVwqyAkbENk9Jid+TACdq/+q
6OoTt/sbJ9ekULVozrVJ/iT4M5BHF4gEdqvRoYMzH99gJIUPAQUv4+Th4ogu
BXwq1GFMuTxpx0WPS2BWIrVUyD7PIXArpAk72aNF9HRCGU2NI9CXHtrkX90D
PobDw89ga46hOULRA6eT7trqYAHtmXxNSStxezmrfYE1mf66uC2taxr5AO+9
25GBM8cDGSoil4M6mBdTmoxu7OPu2JoT0SUIqqaohT3lgumfzv//iRbm9UYe
G2StKtaBlZigarPpN9gc/XeeXA1BJC3z75LOveqRTPMyKnfM1mpFBvtwgsef
cn0DFczyMsquj6W9NoPR9SYNz6YHC5EMHoG9cyFIAskmAN16q+7Z4uE/TFvu
tA/33s2yzdhw85qMGBEWBlcnBnwxsQ9MT1Mj+EoT7iaOVn2F39ZYZZYBfYrK
DZjcghlGAf/BndQl/gxw0EP/j48UeYpZUwBx6GH8cKfCcaJuGChoy77l5Sud
cVLzLgDa1VHN3dgGEwLpJSydEzx+N4fCrvZkHVN01/7NLxtaTOOXItYBcCDX
ohwwejJngMpTq+SGUZ/4BQ6dk/yW9vxLeEJl4uDImlHY28sT4TIoJAZRQ55V
t7GyohQouKCaYkeLohLhipDbmZXgSKDC9Qr2RnBxwgIIgxX//RPAErY50In5
dzLhr8/F4Ljl8ilHZLsyBge8Jf46qaKT7W7Uks8ikPQx5niLaZi8IqYX2qEy
g/ed98KXJSdawKHsBWcTeFkmPypee70Yl+jLuucLEDVYQGo8zJN+ZR+VPi0Z
gVnZnJWFGb/aI7EnOMHs7Oh+VlIUhk9rmstD9oK9OWmQQgw7hBVvOSTmBCTC
c3N6DlHD3/HlNlB2aNRNOqcjIbtVknbGLZ6TGuOgyBqnQoVsvEGszq5xNnud
ISSChy6kp29EUFIqIO4DZDVdqAxGmLfgc59Lmx4J7r2iqTrAQHpzLkt5dkGB
YG0k/sv3t7TFWy/qgyPatOxpAeTij3RS1vZ8MZu2WQqXVSJGFDaztVmZcG32
C7EE/1VJC8HLt26czSMaw6l4+U9jEp6hXToUUMpRLbig4J3AqgNmU3rVg6cQ
69zDEwUM53gzc+r0Nf+gOfIo5aR1wEWNazb0SIVTetxjJMCGUhGZ6mYzex8B
Ss+7Pjlc2TghB772pfTGTfU5Uz+EOSbUNKvYfmith3Vy04sJG/YaZR+68qMU
B3Da9zJ2cySgix7tRWYjFKXM7ulxAJJso/SFD5WBVVC73KrMc0asMREN2qjV
n/XalsxFvPF2W9yLIRk2Cfd2hPUi4lssrm9VlqVX2yxIxXByWXgyhKeTZ2af
keuh+C0kjZOrzoEFIAiIPBrkYnlxjCL8Iwx/d8uFYCr4yHTWreCb7dPemHDY
PXAdFwPax+Q5rzjlG2ObceLcp72MwaDZ+JqtzUWdpTkEyv8pz4PofBm/XSpu
n+A2w2v2WZb9ydyKwIXJ6TslQ4sCfJ/PVwCuySnxrYVZx93JTxYEocpMqT+q
XA4pREtfMTaqnXNvUj+Xb2/DsHt8W1Zw8qAdNgts4igYMz9XLahp+I7djkg2
ulzTznhzRV++SXCgUtpkotnwCcotdrOIsKDjjkh/TvrPenw9t+PFdANsh5Xq
G73fDnEBAgDFmjhi3uQ2wpf4b0Ewvzl9RYI5ujMTfhkCvNDYeqMJZmddGPUm
+y0bHqUKxU0wMpsqW4MwC1yV1XBqBG7l2veYdgcdqZQ7HvX+nViSt/0+O7A/
FdTrSIf3EAKFAFec0pZBmNGqsGnP3SaxOR7hZJI50Zb8FKfIgKunDstwW37U
7dCe6xEn9JOJpfEtznshspM5OJpTjYN3h3Ndm5wyoj1/1DF0Rm/unZQzLl+N
aBKklxIa56aJ0X5619eqgfJAkVUUdBwq3dIhO0s6V3TeRITYyk577alRQtdW
SFobD8EYQq8BqNdgaE21jCMsS3EvUXxsTyvCEL2iPs9d/qg9rBpvNyQHhfaa
F1u3EAb7NLw8hhiXhBeNTW2K27ZrB0wdmjKv2f8rvKC8P7Zv4DKItzuJ/iy6
Oc8VqGMYalpfx3UE8MNvjfDeEjgFC2JwBn8ekPw/OpxQLejnbuPHsKLqUYKY
7dQta7wUIsXy76jOnR3nEtJ90rmYeE3LtebhDJxMGf6hTZo3tnNKFiNne02r
jEe6hzbbVRcfEvbZxi/ZGp+/rFbmZTtLh1VHfMz9SYSNXTC2sMPRGPxfjqsY
SNZA6xwBLPrc5eWM3oyt5ycwTKvB3bcnNIVl9ar1i25MOVHCKPqWG0uvb0za
YYi2X0EGLwhnuepCoRjxxyWQWAGYCGw/Eya/JOeRiZHoPa7is3cxnIPqzkfi
T4c5CaDdNxwBhklg53kACv5FYQTY5FuMEMwvbopbNcU+khuO1Zkdh3pY4Smm
dtk9xx3qX0Cna3/77whXoGcLaNrbiNYIDz9CGmbyuhYaPku95plqxsxbjHQ7
dNQ5p3e0civfcQhDC63w8Au4hTMgkM4IZiBF0oDvrkg3a/zhvuMKmjcAMcXL
/Rin67nDByokhW6ULky8FuW8MADKYhw5WFokhTsQAVHE19mNvBLg0nTv9jQD
9lAAwF0rw0g+BpRXXErKemMJ5dCcajisv44R2nY3vgciPi0gw+cApifAVZQp
uRf4/GNsQi0JjB1d9iESCEWpoeBCeo7oskMBPp4DD2+zwNyl7tnf+gQhNXVW
WmARw7uY4CIjhnPp7vKSzcf1VvppJcdiOBV3GBXuRZXaTR+23Pvdfd/KbFMU
P0kdPyNX2zrqxB9toZpEZdW9vUyij6NTq4HBsw/OZ1NuHSCX45L+3Iw2n4Jc
tRMP9vDoecy/2nWXS7Eqm7RYj5qxQzLbnxzbOHserekO1CrDqzTkG5ea9s3b
PLMal/qk9HC+H4OOGKJKohYjJ9AJ+0a4FWqMOE4Uk6VYpqhWwujZNclgHLr5
e15XzGWCJniiW1Pf/u/jOjnQ5mEvTxVnZUilKPLYDwNUB4suSzpvLL6ZUFao
IjikqjvRODVW4h3L2/A+r/Q7KALylUtTxIjPTnYFUWkeEg1+l6YQProjbUUg
8/2kJwtwXA/gS21fDjroWDXs/HKTRRlH7LxXD6YBOcZWnXTUGJHGZ3nFiykE
gu23pG4fdUvu0rFh45SahptkaOcalN9V5Dd689Cdd9Pg0/qKrcxC+4B0T+g6
I1A4rE5FZSquKPoxHJCWfJ0A/5ZpOu3wgtUvN3zTXuFTr19KURLu0kzhHv9Y
hrXIz7++T4Dp1yaeS5gFY5I2qKGfgS6afDk++0xlb+qFum6Q5d2hzY1O15e0
TA9XJS3hFew0BFglrCWQEqmRx/z3Bc3jKt7b3wxmeX4tOgUCBfOzhCkTpt1n
6MAJgTqy90jx2RHGWH7gWaNT2FLjozkFnKEEF+X0nZq6ggFde10Iem0gXEKv
7jo09oA6D03hN5tEDkjhVTxHqQORsuL9gjQxmdeYImIf2ezu0Ii9XQsoL/H/
qrJ658qLHxfh7zTuz3FP+DZxcdavDAFZq0e08a73PnaH+VTIh06MAxGSB1FL
80nnUQgfkwBqAEKUFf9WUlubXio58eI7VFtbZVES/P8iVNMuRFDV7OOcG/n9
mt5gwLmihftHIerGgcGtvLWY98l0wfyJzM7gGYRJ48JfkZLETQAwLb3crjyC
x7tjPr97zBhWzjMFF7AEaWi9z3sCeEdULqFOA1bjKggsbVOK6J7fDHAfmT4K
zIIjQR/7yiwP2WOs8DvtjVL81b3+uOddqxrbOmKFFT7U3GymHeSOQUEThHli
NDpW8zDNKJodf5m9X6Znjn8eDgEHePYqs8Mx8wDurVLIBDqz/JtXGfSjmDTR
AF9q+F2Rv9cL/5euBfZjx7Q+LRs19xUdCvvLDcpyatLp1DTZ8THF9H0nCjnb
Xr+Op3rvouZmjRjXMe2NToRglyZ30IKZhMhNmxsIw32BbXVh8LwHufx5s9xU
jjEDRlk6VcxLUvQmNaoxROBs1/ND6QOtBuBI3I7Vb4qKeRBfF0l6mYLasstN
qJv1bprWX7fdv3OrkK4GdktLJ4RALL7aA6WFmSRIcxv0Ldijp4Z/43LetgEP
vxjHvHMfqGMph1MIpQuipjCH9dixKvlJnBxuYHtAvgnntKkRBYZ1vbokG0qH
BGMGnfSmUYDqaNrRtGw/OP9xR1nUJp3iSRq7mMSejA2jkOEMu1mHMxyWks8i
qbnjeXaTRvirNvWalcbXDD5YgXNJbJ94Bo7ttEAeCeELHxGm5Sl6i05Abi/S
23vgCeOvA0IDiKgR8sIVPmiEHQlcKKMvc2TCakHLysNekMMCwFyfb1b577qw
LkGAz9UciPuzj1WaZPDuTkr/f2OFZyBG2P1qsKZC6VujCYaKd/X1F+Oak/78
spX8bLNo7XhENF91C1h4Z1IAgQzx0YVXZQYuGB/VUcz2mbKT3SG+ALRIRCYb
eTvmt4QSw9Uf10bbEsR5GRawnFMLOrqMaphLEHH8BkWNkYeVLXHl0FoKqF6S
Frod4G5NUL7CSTE8LqerK4SXsRR2XjlcgfoGVfyfAWta+sFOkgwWI/AkX+HD
/g2bY7Ge8Rx9Jf+P/2jnV/umxpMuAtOqfI+yfJsl8cVpJCyMnhkvqPI3v58P
e6OFvW9/uLs9rD54MouIfEgIAhzTU3ykNTXzB0RRuJHV8Z3Q6Yl19t7UEzjU
Wkw+UVUMMZj1xmqEJz1eCUQ8TofO3z+kVbxzwsSWU9zdJ8jSUK2lxIzx7ENb
lO/9mYLEPx1euzSfu51sXF97bXCfNLLV1AZVCk39TORe3BsPa+zZkY2nI71C
TKHmdEI9pnxEq21nmxEHnwdZ6xQb2Jx/+Q08vjD7AH6gs4+OKHgiANS0FE7K
qho3PJP6a8P2Fr/SaMEEJLQguIuODiQNznLAYGdmOeWaou3AVeJ5YrgZdyRY
btSqriK5KwW5xnUrYUHSM/YNM1JhjbtKOB3Aqm9S4KTU+ozmaQZfrmnNlNLe
e5nADb6Hei1jSYo7S2JhvkUWqZ+8WXVWyPF/WlsDQ12lgHAKiGZVWXz+DiGU
hxurAnwE67kcHf1YfWKxgOXT4wHyeZT5nHwx6SOS4H9rfQNRQvc9Ov1uXeYK
Xxy79dhKfn30FFxfZ+mqUBIjGSy3wwVk15YAmL/ZYoH/FnZiGCionmmE5gTR
Ysrnhz9f/t/Gku5obZfnIHtiVnoa/u1XgAELs//643JnT1WrQ2X5jwjR6UYi
oljIvVPFLXivAaGZWI82R6GiZc4ZWg3WvNYqSIak6tuHYO0sXs59sEPS0XyA
zIOjOPzkBI4A0cA+tNU/nu8wg1LIhg2kvtu9P0og8jiP4RIqX+ufSH95p7uO
4tFzVXi05mjmGcTGSpO9NyUPff1zGN99U3lr6HO+HwBz4waw5pmWf6E1BokP
zDViPouiKStG4aBRPnhYs2gFyWyam8/LbLQGX0jX1aHcMTt0/cAI6mDQ8mSr
52nOvj9IGuU+VnDTN3HO5N4kIsjhtGXtUuOi0kahO4r5kcbtEvFl5NTMbT8s
Tzuhj0GV3GAqYBjPYyzzBhpl2pKW0b4p5pegv9qWzvvNt9VezuOF0osdnPyI
QQDu0kMEvBJ297MiSEkTK9iCFioINQpDbmmkYX4ggDV0eysGzbX/UagX2tL3
t9H0IuG0feNgHKRw6Ne1NXVUCxtqvxV9MKF2szDQ+1IZsgZiReS5OGTqPwrN
jCFU0o0vyOfc2MRtHUsqI6xZD0wtuqrqMZSlan/ZdDGArLU/x27AyMmBEANQ
drZpcjvLEo78ZIAKRcmpyjKWZ9ftAB2rWPRspl5xCxGB59j0mit5O78FvoqD
40gvOdnSlKbcC6FZWmw1SipJ7V0p1+4bg6YkI2RBnVoxQ716jJJdTtbieVQI
0qe/J7rscFe+NFDzAuvfSZrRnS8uu9Q4jtb+fWpXVsQr10tRpeGN2MMajlmK
RpVu2qCPCUB90kxFYXVv+W3YDHGFmh+E4mNf90ONPl6bzowfwIWAvkexEVom
YiRggjLkd9D9GjLM/ZG6YWdaDjbDqgSyXNwa9hFEt4dg7LjPbQl9z9ETsrv3
oGQFGPQzwNnHmh6iwmWMg7yLDCC7rrCQaOcacl+2DGWk0cy9EvCJbGVmgq+I
o6Gb6jX5BEkxAST+LVuBAeYVeNEnJUdgnSkxG3al3s3SQ61/XEl9BriSbZKr
yR0cWuRuFTzTgefM4BIUWhq7PmxMqkH2iKn9j/9TEuTo1hfs/YqFmZ+y4G2a
93r180KKCG/P5JZbehKiCjqJ+KQRuyzGU//xMMMCA3hD5kTHjpt0f31VTZAf
Ga6aJTpSgTm+CTJD1VC3B/lvRkmTxk20Sd9+oHYs3+a8Ccrg47Hx76hf/waa
IFIfo2UcMfLTHNktm8iy/NGJvXD8fJUTkzT6I23v6WtqZgMVfMytorZzwaWe
Sbu87cLvF0ewiziUv4+0Hvas77GwXX/VQqe7CBTxk7ezIPqVRYTMroPhyFdI
JjxynfsJkzp6r7O2R9td7ZuREOLDEPe3yrVva17+OxmFqr3uSOZTPeu0X8Nl
sdP2L6l8GiYw+eDnkL4mzWcF89VLtXv08IgqWA+PB3uis7KyR5k1S9x8OGyh
0bFhweJ91hfleVl80vr0rpvjnv3P1wlQ7d8RXY7Q3oHjlvTHQMYwhk2ltCau
2LOOkKc81610C5ntAqo+IddyqKuH5oCNuLQgEtkQTl+VGAiJgcihnOmxGZhJ
GV60g7+GB7yiKjXPo1ZzmevGlGjDu54J5NO4diT+4Ppp6eu882tOCWoMIyHS
+Ox4JpNUEhttzyu91KhlkxuAJt1zYNAlmDFNJW88ygQ2TnuOdYIOG4+Tz7hj
O6TgEYWevUG0PLYrHFe+kGJHeGVR2NjMgM27cwgp/JBoBqa5B9VsnfcrAnf/
vN4tfWg0O2CucWCxq2U+Dw32PBQEWe8WMkAHZHw/QbXES9b4tcGWMOEJuHYn
DO6rBDwcbszGnoVNpb83Me57lRm0nY4cnP0D0Yb7V8JcJKVSsA8OdQWllzBk
7i7KTNZfzmdKFlWYbzdoYo7+llrez+BmIRkvKQQA/2FbJ3z9YWVxB8eEqGU4
lnAGhgWZbRc2SECm76Ao5qO4EYWuUJjy77z4ya3Q05IsENsqhQDlx2AOQYVD
pN2JZvoAXS06Uj7MseUuq6Voq0jynldSn7pjox8WKolj+XJPeGvHo87mnXb3
nMpB5/M4lNWuIfDHDGkf3nR5U46u0zOQmAYmhF1DcTWR6uuAYTLm+bdddp4D
Fr9+gdeTjAXSGWCzAObRiu7e5vIC/puapRpjgK8Mg13v3WGF6svXaSbVPSBw
UMGtZFPHXSmH4SmvYkkgYXiRFlQeupXSf1px1dAArYCS0NGOPFynRo3vb70v
4BciwsTgEIdPGDnJexGzwtDl5VAD/hR36b3xu61ssWDgpDpnrZETP0eAZXOI
aQKuwWf7JPh/+UzVgIimDV2u0tF9cUVlmGn/uSabEjSQu+zWayiHh/Qmkzoe
EscCthQwKIDx3wZeYXCkDO9SdqHd9Hox9B/nC6Q415tb/N1KtAkFrAqN4n3b
LIQeIQtlKCg/DlAS02uryQZZxUHOFUqMnpapeTOiPh6atsgVhHB2cAgExf+T
k1QK3KtxijLNHow9kGvViI+1zVrdhp+F6zOSumQWS0UbM13KuHojJDQAauPO
lHNQg+vF5d18hndRufSmL00fb5fO5mEHSKAT1A59mQFvGce0HoVJyB6z81SD
1whtg+wAdho3Hz2bPLAOxJILZY91vUgl9yOtcguKZ7GDjFYqgGBVsA+dbHFu
b9Z1kpMDVKfi2gVM6MebtkJO8ns9Pvn9PNcppBzCYS5XGJ3/CCqzftcuQnwe
EM/5bwxnFLL+CNUN+YBK6Qs4gz4fhXxWiA3zFtl/iuKRTj5oLnVO09BN61vg
ItWfcIsf+/XDqxQkpTyslyFoJNH2aoYi16mdC9yIjl0KNFX+lCLOsCuYyySR
8X42sP89H+7Z9X+Vss8FCfiGFg2Gu58JY9uD/WoMfi/WFe0JL6LAyq+sQkuz
SUbW+6f5oWCyekgPJLrkaOv286P++QeMQ/WVCjS1V5UnFTXVgbqVN2xxF95+
kScQDFKyDiO1rWjxIJRmThFnXGEiyETX932KgdKeirRTDQvXr2Qob5ckyiHY
p0vVkiJv4iHuY1L7Nbsx6e1xUt4hNr/Xzc174PDB5dWF2eQBL+N7Ur5dpC3k
esjMyHojiyJzFRO7HIJFgaZBorwYVinsvd6HHlGh2wnateEFjPnSuRjFFrp0
QR2oGYXOqVUJFDsUYcPrXkaoo4gHYkL5vv1j76qfEZyy8VDe9o+rGD56KkV3
KgqVm3BK/5ipXaQtxQgSh33J1qkdjxbLTYUoqCGEmPoiQ4WR06oFD+JjTyQv
ZOf8fWB/dU/QHrje4pgBYwLgjkZo3du7zk2QUcrDapAVqqMVvHw2ZM/Ryvi7
YwRPbsd3nDoIQl7KNzDIhXjIdImITMjTSbPY7xmFhMS2Zi6AaNvVTpe1w2XY
yLWGwqe+mdMe5zmi63BjqE3/sVnQfRbbuUom56Ne2Q41l7eiRxQPvKDKoaT7
4fdDQTT2P1FQLaJmUPWEFq0CSNGxsZfPEbsnN2p9z9k/27FZvI3rwgkGLHwp
bHzloX3QBfd1ks+Lkq/4RApLMXsAf3tt3CA0OWzYW/oQxi56AtQKCzKEaj7H
2+6nzy4jv+9Y5qJzZu8843RSXrRpQsE4qs33Z02A6OEv4HDyfuPnGQZjIbRz
WJV5IoCP+e5p+oZoFZh3qmwAz5uoH7SRV7Zu8W3654EZDcVzi998WRGaJo1w
Co4UT/OARuuk8glAnVIg6yx6WIMZL0r4houuj721nPeJcM1CCG5uah/fqWqE
av7rKIdCWsY+RWCuOgHcYcLNZeqMkHHvkUKGp9lbZKiI0lHPHb0dVDHF53vT
u9HUv4aGFO0JgQ9syrU1RElFL+3N7CwpBKt0NRZJy/fSLjWI737oAYeZlfeG
LFiQVLjhahfWsGyce7bfpXFZH5l7fF866FPdGsdK9AXCXCtDskJggwquROnQ
EKwh5Wua5qSTyzv+OWNg0AblLPFT+S8W7boz5sW+W1CblSOYsiLVVOeYnXLt
zdt7rhnhUQ21Tki7GmDiGUSHkqjjKg22j0P08TfEN96rhqkwllibDzyaSp15
DIJ85T3G16OcW+2WCyNjLPToRIGDWemWbnyYrNclMz/RGxIEevt7VAJhk4++
voV2+xzUE5Y45URS7KYLP6eMy/U2fK4qInYdJd4zSfbs864oKbPRb5FksyVH
tk/sK29YmhHtokp+dyxOjmWs5+mlyPaulHEoYiIgeGdpqpIb5FTLOsEWtHk/
85POZbOpOhGCye78AuaTAW73dvlZ9h+OUSkCBPrSojAMrdy4v2Q+uf4k7lyQ
lgZQjjsKhH5EJ/QPTq7Qiw1XxHb3mp3vd7BXtFWkZ2TnRvIHwteUdoDEf2VY
iZr7iTG159zurZgek3PjS91eMYHUPZvO3rxBYbKO2FVF+lASmrzFoCzjLgi7
aEkkb9GkRoJIkPLYmYLK37ccsMVmwtDR2BgdAiga19TAURZiaTxt3uXP4gIZ
PZZN0xCbhEh2HhAZxAlhIDcmIiYupG+HmAQyp1FMS48UygehqIdZQdNZJ12C
w3jyMGCMig9TnuKA/L/dAlcAL2TaAMVigNqvtW7KDd4+IpWBlUplNxPTDo2e
my+Dtt/XLYNTr1CON6MJ5rVG6UFCy0gsBGr5yyEvRuKCf76wtvCFU7eo9J6z
xOUDFW3opdo2XKDttAVhPfbzNEfzmmPbK+ZXWH/qGG01v/nFCOlvWVJJi7o5
dc3RaLdZKPbGieN9ZKRL7w/Bj5H3xJ463dJ+k4J8fqSWm7Ay5jxqrsLmBsj8
qok45ltnNQ/RpB8LvPddFGy/mGzppgOh43Jf1KND/Auf8tylSUPHOJMnOd2l
Ly4KufPz5USDvoDKjtkEAmDPbPo48gMu+DaMa7NMOlOLRtJTut5uZA1/2QPn
btSi0EoPUHKP3HZ1a1a+YXT+SgvMmNXVCezOC0fkUyd5+ViAmrEUG0QECknT
rYMdW8Q+N+mWjaIpymbC6Jk0B/15w/aciUolJ2Amxg1RMgYkscLij8WzGZfn
vl0CCcAMbOiyJhWDBv0KqxIWzKWuMFnXDz5Z/zj5ec8v8yb7uZksHxtzxtFr
oppSEwNeFtS2fBpoDJPFvR6KI3xrWbfzKC4cANc1KVJ0MMs07l2Tr3Qv96hH
5mydg+/hNTv2+PzUsPGnEZqOtWE9uG+C+fKpX52pJqWOgeJ0e6GapfuvMWXz
b+xXGd1W/inVvpZXGf1Vi/RqaWeUw/NzSsVrStNmBmDZ+SGf0HO/AinkH2Nt
YFBhLFwkbFu3JV5i+smeJhiN2aM9l7/JBZ+ojXfTsqfyoJHMXGubDdcoROxB
NVdHfnjXYfDsJMOJMsB2l5f1q6svdWd9UX46r4K1s4q/cq4uWoI5uQJTegSd
FHli/FfJ4JWx8SM794SJRxFhZesZrKvL8IG2rMkVlaDUgbdioTPFVLPSpdYv
jr/7jumgiq84UWE4rcipW7SVKVK3py8VxcZyWKdDibhNaS0zKhqS55BTtvNx
CyaBiL/hOelWb7X810UCaOKy0KeoR2YpXF+DuJdRXfZSobbJtBMIoOqEvr51
fdYkQHJeOhJ4PyC0fAjplTyy2a7RW58p4qCALBQXqb6iWl0gsFU/V46kDYbi
hTqafw2TKVpb6+BEDI7CtggFY2H/Nwogzl6kLvBU43Nfb2zq+L27T3mMcRty
W+f6z93XaEjnutvk/jvHbqQJHQ7cHYN6FBdn9joQ5tC1TYgdqEyRtJA0Qv0I
al3EtorFDNPf8tTIk/RjRc4EEtLWBYJMm0EBfWnTGXWAsws2pzygnQ7SDPzn
sdomtGqukxBDuzcqhTXTmSocBv6Y1D8mDI5h7Pyb77/V2IEX1nRD7knTB21L
WSvbmCT2Dx9P9MzBRJuwFyt4j6KDR0qY41s69mMw4dfb+Gtw+8qmkT7LR2nW
ADbkqkELTFIJurYckU+/fYcq6YUsVB1Mgrs5J2crNfoKnsgJ2EVr3rlcsOXj
Zmw1aQUI06zxLabjl/faiO8fUhoXa4jYjYNwWrlBFRE5EskayyJLygf/K0dt
QFsuvYbrTuXzHjb9HsdHmXmIUB7UhDerqcRHmBCOPjGjiSMp5MKB2x4u0+Vz
s1tH62ni83guGfTQzlKY/SCAqrlLBQZj2AuMVeGFhg8IbZKL6Xuqpfby5mU7
2laKmOMxWFZQV1ZLUSgNZDSUrx+hNfNOrhmEXryJtTjr0moz3M44sRIZ3ch6
d06XvORSVhnTP5kzZeH4me8bWk9/kmTTHMbgg8TwQAbVC93O0uZmClVkpaCi
siYmXucJPsxExB8LjGZDxjCt2uPYERAHTft4hifofpEv7rcPrBeeSojTqKkF
AobHNn5NsCDBNBON0xCt4Nygwv3PzUlwoo2mErTYQ+n98X2R7kIbmKWexPJs
6hd5yuSoEQoB8JQFXypHXO/7OpgVyl0S+Ra+ee3rfjlnK1W2Dt3RXyJ226ti
uSAx3XUiED8RtLaZ2TV6fTfUQ1MjnjUoXmOnomM1vonCp4JygpKN8U5HFkrF
V7C3BJQT8Jz7uQfsg6+xkhZVWnxXUjNsIGTD0XqbhUAkDC6AHIcSSo6OaMey
84byloryo6fw3Vt/PQqD76/MYqzkf4f/LXyOcPaianBRNEgi70f5duh9UK7l
yXlgpKuo3zwg1zmBLc9uwHHwDKC+mHLJdbwgdoISXcSj5cQWrEUXnLQLj85H
cygqXQrw8ywSZqqGg2V3PFy5vdiYxTb02Kldhnpudzql3lX1r5Z/46Xd5CyS
12+fKpEsb8Of5M/HUI+hyu8fdeYYzJh3gyQJ9AmmUxVCClXmimkfdrgkG7bO
VM9fzAvtLPvQ5dBblQT2k2Ds2bK9CyLWOCCQEaxAPnMCbzjUcB2K+XLtOJe0
qiI4mLWNW4SpcSy2M7WlshWnjzvL9MQyceYBDJVPr1WL955ayJa6t9aU8wNb
9hB7xfoyBXiMzOZsgWlDsUsSf8Bpv8czjmDOVDx3bM/oXNQjsxbMMeUuZfY6
n7iEEKIUrjpvqRSU/ZAJxMkFRuVJYfRsVDyTegEncdcobsSs/85FmI5uJBZk
lNkBciHqt+ZI2b/TK/8bry3W5nRM1ddhBBUUaHx3nO079zHXoNR9Ih/fw7v6
+pE09rswdM4lpYmNgN6cSlJK0WPH4GNZc5nboDDP5MHOHiuyIhU4lwaRoPGk
kmWzm6rKhLHZUyZcWYlbUYSqH2L5gpb9I2spm1iYaMcv0AovEXpCSHyt/ons
GRGBd2o8RSyh0Irp3ErgZ9a58VoZo0bUIrSQzDdu1BBEZvHliJwTRKbEV02J
cgfmazJuRMlthtx0z6X4n6ndoL1ytVrZWT5uvpOwOYttTRPH/hIpZbEF7+Zb
k8VBa55ys6bMsWBVgWSoHD0E60tgdwF3BLonvPfUzU6sQe3nv34C4eybooTK
WTRSDuDeHtOIv5k/SKAITtYL0DSIn7oT3bNIRfpDKLGut4Tbf37Qa/pOMLwi
ghIyxqw8Vk88t4oydu3bwbjROgNXSRwZnC/QdWwqlipXqVljdYCDwElT6QOv
qn6PaRELdxLsGYTJcoPX5ujj/zkHz36NXRcV6uECMPg7eEPpM32BTXQ0gYdb
g23YsLruzTgjuZtC/k4aKtAi/mbvcHhEpVsHrBjutxorbDpxZKC67LUyrNO8
5zo2eZYkBxrYu92A7ybTPr+FMzJv+MwM3njBq+kwukBl3/nuJtDxJiSfmYfx
suRikI0YkDNoNnzvnDfXabth2+1x5z7zAhXRC71Oaqp9Mz8D2mLuCeih3v/B
JEA/hjNrmS9i7o3+rfqntRWf+HpnOJUqhnUeqXinSTAJpUEpeNgdS+4rmqRw
JQm76LiTdio9uh3K2PkahDSg5SgkFTiZpy+Elj6DsH32KmX4BkMqYFtW/tpJ
GTisfWEJ9Dc91kNcJJfr59XJ5NS6cg14Ry2ZEJdTwORy7CMY+eSPfVnfzFww
KZWqbaX0mZcNdKWQD5vwfmCEoPlxbYtPo7n82GA11lrWWgZrr1AfEmzPbE/r
aeHUNuirQlmYJIrZGHN2EVj06yZ+xgk2RnxBfatuUPMQ2LYAbUHwVje2Zihv
bWLSLXfp87Bv9HKgGzVGU96f29ZCH1yOUoiR76tE8UHYXYwPHqTHpxuQ+8NA
CIXGO6EvZ0D2aT5vZdbkqtOjQEREn9T6oOr4IqD3DSDPtC1m1zXkdh+ejN+r
Od+fACF1AgQeP3BqcaqSDPLXJVruVqpjXxn3NTivxDYqlHzs7SUB/N/nNvl6
/wq4uv2hHXRi5yrTEBJA70Hl26IEk6GUqD8Po5eEG8aJU1MH3Z/WsFyBAxxx
uz9hC3sP4XcxCGllkNm2zw2jof21GZgv5DcXPu+hITHpkiJRl5ScblH4F9VR
CpIcsxQiWZ1ddq+CRxitiK2c/WtWoeKSMEbSWIXbC1m9bHpeFdAEWAHOniRH
sZHEE1oUuBbpg7XTedAnX4lXaip3gI9F33tf9gl94NnRZWKVmQNYUyRiNdu1
d4s6L7B6xNDA6Ela/HbJMDKGScKURmfJlDp6+//sVaOK2d80TFLOb8xWKp5x
yEkHT71Ja5YrBQG78hOHS+vgIhcj9HV4VnHofhApuJOqDYF3DZVREaYJ5lNV
HNmmFutSmT2ORnJk7PN7Dijegf+XBiJ/lOB2pqzAgZ8q7+73xPHvYofMPMEH
4YXT9jkUUmufF90c8XktWpaadt3CR9zyLNYXmRctsvpASgjdcy9tqPkOmGAU
UupgbzMA7ery+1ZV+EzTvJqiaTW9ArKFvhsxgD/C7B3C7Tai/PI9frw6noKc
itVdXPh0KCiCdrsrYe3Ymf85XS/+OJVxR+zbbWz4SnM+GuzdNl7k4YcU3K7G
r4sLsWmBNDXboh53qKesRb21ALN2D5f0/ciFYttjOC25RIEmyPBvWHXlyN3l
zBfxkXUQr+tN/Ysj6OtkXCDy5i8fBLCc6Ej9Xr2K0PQtA1E7OT6EZZF9vT/e
qKFk/x5XHPQraA9ty3O8Fl2fSB6freZjNN+5GNnZpRcuH/5YjbOzfRZ20lKL
HDdTl5NI5UIUWscDwU8yYzTCCr0ELRke3xpvxwzAWKVflOEiTISJQM8Xwa/r
42gW7/8uDX7H90obmIi0XZUU4HGO6wkuBOGjHH3FKaI7MaRMVQL129zyfevj
boJpJsh/MGcwd3Rqw4VNx/9pXnC0hib9O+qbJQH+pz8etpAZZx2f4XFk0LyT
6zSuCWA9KxjcTdnxgG7NuGGO60prpiZQqJJ6h8LSf/7PuS2uVc1tnq/Vwxkf
hXW9OBHA7GhAOSShzBdVcXiOlJlAeueV/ewZhYqlFMJ4CpwURpYo5Uegfkjs
6HwtQFq8CzoBJRZNpe77iAKBos6sTPEt0kd1mB/E1am4R62OrAfDUJ6aksy5
+ADGRpyRt/mmfPfdkxJ15gKjtMUFZRj+BqMvqGlrRdr6VZrREKPJIE6YPPZ7
uqQuLU71fUOIjF7/Y5n+mhvQ+Kts3d0tux/wrKvthj7sNUETHPxEvgWEMmKH
F2d534b9U+kwPSxbPB9Oa5pvnw+77AGQ44ifyMT5XCUQr9Eg4U9Iil+qZ4pw
Y5Z0gNnTz2RGDfQ+5UDgoIlX5q3Cr0/aie6u3VzbGeFsB2lhaETCjxLqtBDr
HwkvsmcVC87DQWgudH31SSyBQCks3IdMygJjsXc+ymGx9Rhqu9MIbOV8JpZ7
walRHUQyGdR9PuKFiTN8v4e5C1v/YUScihtBjTSAHl0kxW2dAPEzXNcOs2q7
tXdRao3qmYwtHbOaIPjzmiw5QFG0uGcfbHwGnBdeQuJGh04ap7tYByzFwc3s
2QK+FKWAVhfpfv5VvTWUmdoacFy65H3X1gcOFNb6kFcnhdXlwR7qCOTCuM4l
TjATQZNrziofJTcMRdcGP6F42o682+L5WCffWpwgVWdp3OkGzOJog+9jdZCr
/oFPbZYEFe4PH2Hfq6RCSMUu4f90RpoNGDKq2GA2TYp/ZVR84q2RlR7m4KRU
2P1uZwH0RbIoqmjIZ9VcYtuP3F+g5IuT38QhcrdiNLpjTMdTE7kEUFGg/R1l
/senb8pxvBc9maviGrhlTQXh16SDLQSkFRM03+n0YvamIBvVtUFUa2/+xMJ7
tqT0IJFw51int4nlYT5svxsLYa2IclXiUqKNB4RiJTldpH+Uk2u2JXQJcwq9
HAeyt/vRG7b7C4FPm1hYIfTcZRoP1Hvijk4lqjN5Ma3bXUoNyW9/gGAmKe1s
U9IicjVpdm7E1pEvA/COpTGktDlOWFQkCt6eAp7raxja1d4p/Fj9ojyT7XsC
3Wj+YJLIA6NIjerP2lXmlCNgXlQCRebUocFkhaAAIftapm9MaeSLUDXphtr0
KecQ+r0bJIMk1Dn1TqDv6y7+oCLJc9ktG0dVV+5l8sq63CXJclK4jIyw6KbB
yzP2bdCpMAv2nc22+6wHcEdANVAeTIGZ1NiolO7ANHA4xeJLvwY2VMS7G6vH
kGALxGtNmiMgQSs7Hhk+MjJR5AocAAzp/f/jKT2rn4JiGTmE5Cc38TCWeLHF
ocMtkZm0bjat8dRnPW98aFNl84Cuq7jOaxhGlGFBrGZ+XsTv87kahSYNRcQA
1eji0FoVDVIrBbLvnRHwaExeX5CsFhLuTUEB5eLy8cJIBWRdjt/mLFWtpdIj
J50ldv8rLbXr0fMpi+otI2USiZBR6tIFsAx7QGDeNWrUxFPYeF4sDoR2r2Pq
+zsHw28XFJppsDdoeSwuG8sBf8ZOuDQpRmmu6GxX3FegrrwPdxlxB+bbmIOj
cBSalZzdwTAO9n1zncv6DLhhWll87Kz5KrZiqSvrggPZnvV5KyzDhdgEKD+n
Xk9Ldt6RyhSI/IxoC/bsqw2LOy6Ej+u3KV/v9D3IUh2NsbkDEDgWJECO5LPP
B3ezmXBdW/TcP8AwruZfLEwslNilLGSrs6KwU+rcSc82Mf0rii9nHgVRDkJJ
wrGLvpd0vfilY88TfHPLPik8p11yLAD7RNE8Vtko1XuySuhTW6EAJfzghuev
9lgBWU9XYznZEvUSScG1G3Rq8h9pspTYmreVUfL04ayjiQRTM+7Fmb3MJhy+
nRrfz4SzG3OsgwToS/0tFmOhLsuPzFNtt97dKmUXRWsIeTwDDZiKK7BAQFVN
onklTFKojuddg1XDnr7/bbCajCq91jbqX+2AWv9Mc9cIp36mQT092K9Tt3jm
yYyNM4ftOjZltuMpUshtxJoZKrwj1XM6gXXoKzXA2W8d+OB5HRRbXrzTbVKF
ZaHNioiWp4uKN7SZPEg6+qqL0wSPctLBk0df9L9iudNrFKzg3LIKsPpAKQLk
Vdo4pBkeIvvVEAcPw7s9gUZ425t1duABa4Aqy5tRyXfAw4Zke4xAW8xHZ9VJ
lo7kaJhRay17Z/XrM7LMTiJ80bfcWqzUr1bqlcpDQK4HgEYA4Sxgd9z7eUkt
ym72JWJ9QoxJE/+wGAM+ihj9kWvaTbE7aCSA33FQgyfS1/0s0iQDPF6EIhJh
Eroo6qD3dj3AugmuL7BsB2AFFyRECqWpa8rFrViIwkYO/JDsb9aY5pLhNOo+
CZiG8gBono8dpk+0jYZmQMgR3qC/4XWVKJF3LfAvmy5J+5+Tw2GuciVfuuzh
ygKzNOWwjX3Tnt86D/sPQaI565988mZPFcgoro81bTs5ULIq2QdoO4Pu/02A
Cr1PKbuCxNx2WThocSKxbyTFEmKcOvMS1R+0VvrsK5zG0HHU9Z1yjlfUv0z2
SDFKAaeeFbcdVF66xODoqzNBEUWQuAUiifk5A30WT71m/HjdpJWA3rZRlrJZ
GS20GoFmukmT48C1GWRSoRRbR1MI1JMcL1NqFK6zQI3gSNE56QP5or2QSdDL
ZLSKVeH4+Q3tex0jqmpX0E0nQP/rzw2dUsDvgZ8UBmttvBz2fC1+9EXhqO9r
3jd66QGeInDvAr6FW5Kj6Hp0vNBP0H38VtoRObYZP8WQWA5m5CNeatjn10zL
Z3s6RCcABLxlWBlGaPvkSMeAXVvS7PaPyj34uh41xVhhofXGvz/kgV3rmrBt
ETRgzUeiUx6+HX13zVpZ9vC7nIZBlJMf0IIN6jXJarVZvxAzstlZV4FwzjsJ
q1vaKYKO34TS/rDaOdgrvFCGjbFej2ycdq+H/RhnXDcLf8RtSWE2MXrIhLvB
u5UbVGAbzL1Gnk7ii3GmDgFAyRZZcHKmPk9rQxrvkNAIYzZvy28krxuqz136
7xPdXwr4YKzBlyYiFrRJVOoQaM9T8XJxvqb3eRvnukLiEzaDY1AsY6GlHD4M
j5DPhbs0JMiMeKsY/LjhkUE6oahAVC7QMdGhtoNOA4AGg8rWOlbb6d4Pk4+j
cKeFyepxVOXBDmSZHTJ4JAgbfY7XVC2ayVUXOjl9AF13TbEMdTNm/fpsQXMW
1moR2gDhrLbwgbkTfvrU6DmhhjQp8jxs63A9LGJTByMXL5y3mLvCbH6mduJr
NyUhfWycioyKPw2aMykC4ow1jSEBAdGWR3MYAaJrSrRVN69ns2/SY/Go1UMQ
TCAwBjFe0172f9xuUgpib1QhLCrQi67wpcTs8xHFKoM4FpkrV4pPsy6aVaTO
b9HlA9N3EOUWMqHyvZzV8snEUvW/ArqCmItCBlkgbOjfJEk+qgnPRN9hqBb9
I362+e/E9jNHf4pCw4HPsCAbfb4lkyB123pkyDWR1h8xn1rErCmkvpMD8vGd
OGZe+UQQ+fYbsus412tY8gOrL5+WJHPMkfF2n3K1SWp0jGVrML1ETsDKhsOa
WX+aSETHoETv7pGnBs75INZQUd+0P4jhBTfgkXV8DZt2yeFu9JD6+wRbo1fI
b/8+TECd3lj/BlUjKGPnq5T2o1oq6C3nCDT1oV2JzDgQoMsiPrY+YmfdIPxz
8w3V0NOrD94YsoDN2zMZbltqbpV5SPcUdVk3wwsA7Uy+6q0t0dU1zwnuY4nr
/YvpOOUgTmsh4NNq8rkzKi7ssr8OkqN7LXA9cwmkVb5eSA1iSddX5zi3G6uX
FqLoSjKpn83mdgnw33wjYTVkFiVpvH6y/zZ53+T6WqQuZPF00nA5IdMB0Gth
4lL8NgaGw7oovQXD6B7SXXqS2lNGcXYSnbFOBeQjPFd4XSSJoA4R71CdVUBd
UcclOqmr3DgkY69sNb0q92rICPxENQXUGV7ms1T3GhRKgXwqMSjYXPfeDZuP
WCgCv//YO/nzp9rt6LyOdiI7z5hPJIh56ygej7BxDXRjIjBFSycLeb0IlRdy
1t2oXh9nEXCplbS4HVfXTeuiWG7n2eThmmz47DCmFUZuz7dd8tt+8E7/3c6q
/E60N/cCT2L66VdJslDLvDE38Cbtb8IJyBdTrSw/naHTe1ajwf4kIKPe5v96
PIrm+tO1jC8UFkUJdyZFlUqwiGDy6hkZqaUqaqppFLRKcqf4a4FxhtZIboG8
9+0ufQce8r5YLvyQzbffNsuxfFqCHZoatExZmcSXsDI3rKX5pMs3KK4xpYXT
MIB/QzB9YdqM1jqMKP8jokDm4v0tD2BSZ9AG6hXbVKuZYXRKM2IbshYj3MsC
q8/d4YggkFOQj7q6maSDpA6LZ1DYOL8XXwJB3i0LzGcB/4dmYAnNfeNVUoC6
seeEnqtZsxxmB9MLO898Tn7KO9o6IMoYavsUpgExS4hRbO5L3xX7Esrta4kX
RrDuPJkXwBuyfO5JqqJfgW8CwTf8jOY3PWndqnDFGSV4Anwrkzz1FgXFrbR1
b7w1n87u6Nv/c2Wm52/rf4l5yhu4Ebf+BqploLtvY2/yDsaBRA/Ur/4f/K0e
hmncrLWCh820I/7d+fF9I6rv70RHuHJHtS3B5urA1M/LUmbPtZNJOQAH+6oL
uPMtUUH3sR34YLD7El3Ap17FfifdHyticpmOiNzHr6zpYcWkBNtjZZCaJcr9
FYV9xgI9yiTop4FV/6yO8gRaVKLKUHUpAyt5H6YDXwtO4kjDQPKYWa4xTyN4
oCfJiI5ycXNKz+nuu+JNxlm3XZIGJfWivIzbGj04R1w3T53U/HOTv5vL/XeE
YE50+VqGrjryw4tQwOG7jgbHJDi9qOAnWcPvp2FFzZfNLpqHaaYFoVgm18f/
S/SnO6U7tnq+0nFcEIzzu9gPd9tBrT686EaVjYw+VoVvPWdFDUvUxcniWOQe
kIZEQGODJ9J1bNR/G9fnoJeyMKMR6/izkiU931NUhRhRdIK+7mE6tlTi/myD
s8bCAOS+OouIidQDitqKFjjmTkk85adX3Azl2/k6f0i1TYTSpn09NJKpTPRN
3lFC38JYquE1Sz3r+LQ+fuMee7YTNJEtOYiDcE+qbHQ24w+xLBqRhVJs9VQu
sDkQHaBrD4eg/jwsvRaOWXctHXjFH22CSKU+U/07Xl4EtZ/fRLJEHFYqczI4
k7k3U8Q52/EYInbF44vzsJS8tO/4whf4dUtiHYuHL2crJzs5T9zXQRwEf4lq
F77J5k9Ru43HJXSZF/AndnEZtWzpR0yIhAYqlqtFtaVTfw1o5AJinpcTccyi
youqI24iioldBYQ7Wrez9ta494mMY+nfv/r0PS0lePSrSs+Tnvmh/zroYmaT
S82BdDHuId6C9tE8D3EUQytIH9M3qmfNSRlqW6iyBttzOZFxxB4h7TrF6l7K
cs129BJ+1y0SQfLeqcHnnI+t9Y/OU1gXmbkqtPgEXpA/1d6KnBJ8shINXWrm
zWL/MH1NPtEeAYuDowWCiwLfIy82ALBTgJgKZcRZmmJcjYcMxriuYRP+czJn
KLUtUzoE6aPgh+dai2G8LzijFnIhA0xCRekG1vxDgGCYwUwnkC3BLgbLp8AK
4Mx5XDtnfcgA3acuQDyM4N9yXH4uiwh0DaVxwatvbIAn0z5gEfoCODUuQpQA
W6Ivn2fPzfurt7pFKks25PV8YR/83IAr6U7o/gOWqvA7dWSW4aJ2u+TXQr8S
180qgtfU3t6DpcJSqI9Pg/pyLdtgsH4HPisb6XGQIX0/ucJdxreccIWd6TY1
D38jElRDSCA9yZ/4hlKiD5YgVCr2Tx4L3P8IYOLz40xtGpgcAjzTaxkDaU8e
L4pKCL7rSSiJj7Yom0HeymfFjiooYJPIartkQ38PhLaVVO+VZqIIWRy3mrxW
87Tz+G/Qe//nf/U96DpAz+ypO/iiUsqIRLpkV407iLHjoG17Lp42cMhP9K3k
WSAvyYQOz89mNSHhojOi/FID1DdXWVG3pwLGILe3YAmpU8pEIZVuueii4EWW
rmHYWFv+GaCR7JSeeW6lcR8SSKRYYskoaUSC/aUHEQCUzJzKbBlzvTfv7CQJ
SPZ96cPlHaPSc3AiFRnSDR598/UPI1VwFB1TJoUVesGNDwPXovckO2HFb6vP
rI2GnlN8gDH2Hf++I55cIsKNTMz6yyrDPk1DesOl6iEvJr3Zcm6rV5qasbzT
xe36aojxBhKAvGMzCltFBsGrbAvJKngvP76PYobysuD7IdHxC82RGGp4AhnX
ZJRtqrVrHw3y/NyBPDeEeU0Z2mh+GNrrH2Ob6an7fX4mQcSRo3e8vA3kl1hI
wh9Il6NZEm60WeFg/BdU8JJZDZdclqLqjbcQ4Q4NwucMrihs7qBOuUZ5FLzW
cfFKGuu5ihAZmwenLSHypbCwgUZlvEGaFIKFtNMkgA20j42rxY4Ny5Eruktr
SvWqjd8taQBgEvBfeoExxy+QUMlGzZrZMkYiVr1jZ+JhhBR2tbg8RNeAD9cj
KG/u+xvmH025ZbYSdFrwPwckGgwjmxEO3sjtnRYLtwbnlyUevVCSdpkIOJnw
4gL88TUfOr2LAn7DYlzkbN9owu67TwYqOl3Vjry7sJSA13s93q2RM9PgWjez
wwpuXMMY/EDAXklshgPHnmTx+uqAsIYR0uBox4TDVyzqzQYYfByKE8sigsbv
0Rt8pvgrlIBMaSMKy+NBQQDSSvPDE34OA5rxCQYqhOTf/+fjVd9ZZkX8V/Gb
NGmm/MajNz19LPvOJIeICr9eTjCtCQ0aHoQvzZec/pv1DzS4kDHGAYprew4G
hB+yCiw+kbyzPS4Z0G8xaKYkgH0RzKCLF4jb7KOeHcbPp7OWR85qOK7jGnVe
vPD8pG37O2bUkZYW/9mS09owtI5WADU+PZdMORft9vEEGR8itOiUV7cxC6qc
YUnSPeEXG3n/vpaOZA7aGSXInXIJY8EUygD1B7+uKwI+BMKzQQbz9Zos8emJ
1kFBuWBBoXsAD6+TjkrdUInkXoTp74GfmxgBQ3KjfrlLjjLadBpdPHqSc/0v
2qZDC3/PgsYSTU5s1t6uzJ5X77DICnb3lntMQPsk16B/PfZ/0stN1nZxrwtu
9bWQkdpjXZLFrZdooVHrCaQVXQ9cEA/mGNvn1Yz5cJv667Jfl3Qm4jpQ9Osy
weR474VvvzStg69cbZlO3uup+pngmDTw0byeOqWOOsaFtQZOKvpjjnnNOHtD
RiSr759iVU+RAy+jM8lIbH/mpuo7EuBRpqu7aDrBoY/EAxpnjYHgEHw9iXLa
8TLePLdIm9Jd2Ro0ePW2P8h3MVBvUBK9m97KeClhI2Oy9qI03z9eCcFZGKTs
KNSoWXAbHHdkXjgajNHKdD9lFFxtcgTMfUhoK0lnUTWOhCuLCNdjocUVjlYS
FE306lR4qGmpj5+zTNMoajFcaYpvSueyS0d1YBUMRTXaVJkVcncMunmLpsWI
rOyTRm0uC7Iao/8SyTAbd8eR20y5j8JRqJqXypkSiDDMgI7m2I2ZB/3EvvDT
q3x+IV0iJos18rOCBrR+1iy+1m2TWn8XD8V21mwrLxyQQ8AEenRLWjEokhir
AGh1Jk+Y54NwATqUd0YCrX0k7OV9RocVG5tLbJI1e/PFyaqp0YLDK54/BiL9
L2lCCzTLkl6hUvflfVVn/JBbf3gfb2kAH3qvUEsTR3i81sA9FAqzQB5uQ3dS
iuNJmYtkLkyOHkrjYP8eo6d7ZT1bJJjuYQ9n0IU3z6R/2DxqggLh5jgkIXjC
6rhWz9NiEAJoKBIVD9/1wadSIUDSiG2tAkRBDfoO+R5zpdDEOl5vZvfvaxWj
u/V7yG9xsGwgizPfKPUEJgfAV97fz8SuxRQKPSj7YkKTv2I+7c5Rh+jBxNLx
8EN0fJtEX21WrUIXe5JmW2F2WZdiEltY8/YczXi6RAvw8HUF2FwQjK8dKngb
Jolbh5wYzUBhI6ap/KIJTS9KTYq09DMMB769OgkGwIeAWvA8M/hx336cCYaK
IL5HDRsA4+1YjFe6siGsv7b48IFWbnSk/eDOVeP4MwrGTpzLmOKhMfp/GlrM
FVVn6pf9LT6OULfhqIFKCde53oV9A91hLrs1CNhZmFftCA2Xxs1LLpmF3uCn
dTp6rJ3wLBOaH1SSafpjk/ptSBGMmBhWiVGBVDHus4nrlSpcyL+EcMNXQm6C
l0LYMSaKUrLeCkmHQVprySPQii0bKlbNrltRjwe6HRRIkIl+MoeguRS30YAJ
qg59nrdS9qr50PthQ8zMB81uwLCEaxgEG5jf2uPeSIgxUYqtS/Uhq3BPEvev
jz8voIIOvL2r3RvAdqoPfUw4S4ldaFrDmdOEabZMVtV4Tz+sqqVELM1mXLlU
sfWR0rmJq7hmfrQYquJ9PYBlk4PJ0rCihbVyRMOsUv0+++1Eh4wd+0cVQWzD
R1HUJRHz77nFyRc4cTpLF/TW/UU44AQrXUXWgfoTFZusPFNAGN9b8Lwi5psC
eUeaxaU/KnnxUgeWJsO88m/qmkDC7QmFFhSPnNjTA5BN/YR9Gu2V7YzgBQMv
5+2/8wWE4Yjuexbltqj6RUMZpRycjWncQn99TUBCXWBkKwhoiz3Ys1F0vg/R
zwqfnsKBnaw0AAVCj3hR7cX19WYDML0gpf7DgTUGFzeRkHPVlktBDhQH+izP
iXZFma34M8cjvqYpmoEs+Gj4fc9uZFy2umJkgLI8xlU+MQ4NmUk1iqVnuxNk
Pp8blUiQupSXYdC0MjY9V2r2nGwwHxEXJ+br+ictVln94EE7P/XRfB/+urRj
/nFOEYs2Ua9aCI4Q1FWG1Ar8R22PifADfxF8L2D/8/kXaNL7SKEr44cDt/Cy
rzLZxaynCKh/xcU7FzsUhyQeDIvWAB6DtxULmvV0H9vx4P6jZLkseqbb9B5l
vN3RAOeDHD2roPHQ620ZfipXK96YAzIEc58tVbZREVt6rYfIjtrYfqjS9Tni
osxbDsqIw1cVSF7CTwIR5Kk0uRPZ7/3CX4RK1JAkC4fvcKhV9svL76xSKV5H
bQ4JKBhAXjE2t0+r3oKbCliGO5vJHsONB2K/rK9YAgM9HSZ2T8DjyKJVqEeu
yo5heg9A4T6ENWgioKp1iDcfxaiy0PfjoGt+GgcPggedWcCT9d/ZHGdqKMlK
w5oM3Sczp0jgINk0gkeAzN7UV94I1dJQjDL65sgq3nPQblSZa6UhMysAnWHz
/aKG9JYxpS0LAmqHP9pShSAHSwBPIV32D4gAy7TU/a0dZNGL7g3ssskZkZiC
fqxEExYvBwVpwZ4DqKumAsbfNKdWiufAPOTJnaznGV9vaXuziopkkN5tYHKg
Bbsr5i4D0KANAFT/RRCyptGRajIFkRWgl2H86oVcxt2+GkD0QQxyOwbt4Ftw
NUL3DTjZKrKtY3hUXS7qqkBedgNt5xGWVygCqvULCVXKfWimlv/LUoS2/jqF
wSV6AI1TdXD0QSBTOkUwFFsDCJyh1aCIVoyecWiiYJl9ZhvVVrEjW0XA8uvm
d1W39uCwgCg96RZMT8A9nPsP1TMT2U/AWXS7JVK+69n8GV7mIb33v+QVoYJ5
sdtFbrb7iP1w+aFSOZQtxeFWnFmQMoxHMI9qSZnjpDfaSc2CD280I3JfeEkK
XcvqknI/0KcFxzZwvjDvJ3zj+rHWyaZKZfacqdZnJDz/+aEwZnFtRatypKFN
FnIFdVxNoBNdErdsia0agaR+1iK7how2QB3KEPEhzjr13OU+86PYYf/0ffQw
LXBd4yF0OwpvuJO7qEn3qQUaN97qjpa0VNP1Ay+/5XX9ViyCgL35daIjETPh
BwmLH7ZCHkyunlsFUw7nt9eCslwUPFHc4GkazIV3SPhJovVJndoVbbwxoTWe
aNffE0IJ/tPFsxDg4YdfKY7I4ahtbl2s4TcQzxk4YYR6LdW7PnlKHaZAFyvR
JQD9SOYaVBF40c1u8vz51N60yZhm7tQ5r3NhmX7P22NvY30h0d148Cp8M21h
1HCAhuwFW9/BBunX0xSYECajRcElcUH0JUQMmoKvwQAIhFzVQE+FOtdz6gVN
wqLN9K79ikZr0cu15LFN654FyRGETmXcva3sQ6JZtEEG8c4Dr7S2ic6buLWG
ncbYwp20eBy1YOMYnaCJ35tWpNNx0+tSLTAj6ckKSFGJY1w8Vj8Sbk+ZRknH
JndE0YnwndXYz1c0fFr3knqd5+TjWN+xZuV7qfFGE3TNcefySjNMAjf5nKqA
JRL5fO61wEV/hp5Ez2O5a8FySfrduKfVurmc4SgRBX+INu9HmOn6sq2EgOss
nVENRGTbs7vU75jOZBRltkPH+5EeYPmU9/ecVscsKY4+L5nnHelVjQn4bb1a
DG4eNupCmoBow58WsoHeezLSdRPkhJVGjPIGH34GitEFboXzSDBFmGNfosCc
mZ6nQiTRkCZXzdTqGsGD1JqpEfTcfLbvAq3mHkG2HwZA78KnS0ZfAsTecpJh
SSmPVcLxSDMAIUat0aYZoMw6a/c1iSc6GH+U+dLJvqmRsXCEluSv1euR+3U0
ZTUVA3qTAlvCJ20X8NU83z+RyNiKzj0QeVUtPl3HioA9ylOqWn2mUIQcO1jB
peh+FrvF0e80BrGbJnauSqTNhVljXWzGi6ziE0eRQALBe/eUfF9gLAXKHaL1
W1fKpLdUh54vfg6tTO058dYrNE7dCj9I08XUsT9aAlBk9tTCTZ6nxtS8szaK
8dH7ohhiiBcUNCAdPnPepwnvTgHRVCjnvIHeDCNs4vLN41PJ5b5DjVZ38xpm
i9rK+uQJBL25GbsMioOUa/yIYrSAxNwuYPrmWKpctbgwWxVDRSxFsdcg0v/4
5lsudIAUZfRAIq5AzKxCiMZS8fCwiXcjM+5yw9ToWqaAi1k66D+esYPiV7gH
F880QR+PEibBYUQWltzeV8Pa1cojpSC4RKdXyMBjAI2PwArf7Dwruvilxz55
rLK+lODvSIvZKr0vswAlmeVs1zg2ZfHQCLjTgsiAfvsBRJsWZtR7DH4a2+xI
TleqmQI1T5cv/SA4OzjJuinXQR8UYYw/XI4XlAzi17quNztQgZ7zGZsIBpka
PGNKDQfGPafTtpjjhSOKlVDxtvSgwgnLtsHM/jV474vBTsbTrwLUDk8zZKYU
5ajGx6WaDc85abfMOUJ7XXN47KGxxvy6pgmVC/tYaAr+38cA3KeToHdDv8Xk
3ZoF+O99P99V5EUMwiP7/dyJ7lmojmMQCMjBk5uJmDgyL1edEwalOzT/Qo0b
/qMSPRXF+h4rMrfUidNTSLuYBKmZhPMk4+Taztp5KWHljMWOxLW/1Is+nRzu
ut3FX4X59o1TD2MtVQ+tKfm08eKB+z/jwdvMxhZNCPNfrIQYnlq3Fsd8mv1c
q6EkSQXK0mbsnTG9sJ8Lk2FMscLbkmpl/zC/nnIZpzcq32sDWPwSDi+Vhgxv
iTDfX31+A19uKgscwyyAPMFsdEBfrsZlW9aIS4l44KwhDPkPh9AGVuyzrZW6
/H7k0RC+mkAl/h5YrvPP+YLWTBTbAAZH4fg8swOEGP7bbhujs/gWbDqml6LF
rKMPxinU5kI0ihZoU57CEsYtBPKs+en4pDEqrNI9uUS5B0VK+bPFmNySz/HT
GCmnmlkK7LuxieIs2Pl67w8D0aZEGkJj6VfKpzo3/6mlFW9tr1w+zpG+6J5y
a9xM6+E6q/6gaFixzT5ooUEeF12W5ElrU+qOQkummD32qKCJVDVQEYKSvN03
fQBTAC8M3FU0+LXDrWzSL/ni0bo54tk2Kb46X0uFCsnwUCIqrry9s91QFcDf
3KiqfsmXUg7yr7DTTaYFn+QDO8UtJwNUqGPxVe1zf50z+hPg8N6L67lq0Qm8
XDQd7S9QDyX0syPbN1XWr8Bcill3QUvVlRdmESJds9PzHA16RA9dnxZsrgxN
65lT5Qrzox4lY5XSoPvyCXVhy77xhuQxipbJJBHZhn6iFF5TJ7+QqXaMyldL
wxMSqr3Ak/FiyDsskHBCMJVq76QSeEuaKXrO9t0Wve5qbbnPsZy6pHywV7m8
XYeporpidTvQrOZ6vD6xIDiGbgWnssr/NVofE8uT9afv5ZCNyOZ2nlaTo5f/
qH3bONJ4W58oGK7nEBSW+zaIo8gwbfz2hrU3+VAVbRhDIeJOz20nplIMrvOx
p8WzqbkMhuk5ULmXj1XRDUUOIquGlF8D2Z/zdO6+QhC2LRZYODlZr9Zng+lC
WVP2SuYQV1u2FxU3JB1Lk7xdSvL7XWoqWaU3aGsCXJqI3H5Y+aiQeoDRRd1r
be1MhSVXa9XpF3TotE58lK3BGM80thKbEcAJyrg8bV+pji6I5soySa0JY+yN
APlUEqpnwRIMJZzlHpaUSyuP7D+aCuwTMbFWUYwRDOmuXOmAiltoWVFupUmr
8N2MYfeSH86Idfzrg+dSaO6oVJqz5qvc6PZdCLUlleJtq9kPf8WDnytAKk9x
KPqQmUXYn4ueGEc79p1RPoQYAI1DercnMVLG5WY46CA1t27asnHekXovRrCN
bgjo/3M6UFMsB1Nmpcm6U41XBi10UWqq2blwR9ay/4pXpZolYJjsUM+2cB5Q
flQOU9DeYlO1YoRQ9k6svgOZ6BIZgJggua6MKYNbJSTVG2QiZz7fG6SSe+Nr
Wy+S3+agLNghWSGeQWerCtkk8Z9sDjrxgMt+eizcY+ozoLI7fdFVhEUYvqCb
brljpbQ9+KMy5bg443qrin8/YypZX5uHL3vG+g2KNxTMl7lPq/IHd/kouFhC
mzYgI6zBWqhCBqyeQRFoW1yfWrRC07UVExRXQKgYqUKjwr5MaYxhQGPKT7C3
NEFWrHIDFTj7QoRugT3Ed5sGZ6CXcjbG+MtFvJFwsPQO9REntTvTOHwQvAqF
irKoYsphtN2GG9jLPv5JJIzACaXva7ceNxYV9GNDAnZICFL5V52m6B3mAb4q
oMoe2H8ka7B1daHmoEuBiPVODVwE59uKtxO+azrTqBUsCKEyPG8O9TwSB3WI
oO3/qdlwjInCtr2vtjnsKQjdz4mbOKKSw37URTfHKYwHZru1lQ7gZvoAlvcE
7LVjrzhVe0tm6mgRmMNJUteuXDtfnO4/5bVOjmWfmd9011oiRtb+9DvpL/Ey
vMYpYr4HPXFM2ykrMXqO09H7oH66h4aicZHZ8qBC3NcXcOLx2+tZHgHCz5Ts
QKfXvBFB+UU0ZHH6rz8hX+h05htVGVW+PmPULZum58XL6tFRv0Vk7q93u9pR
Nvuna6a1+hdPJWDqiisE75xz1/4N0XOw9NIejcph2hyLc/oGsEtyXXvKALZu
Q6l7H/0yuGUr6xz/0YdzKGm24VbW+92sUaFm1VotYoLzIfM5K8SieLBBTOpP
YarICuzCRoYyBlQ971ouj/hVb55ilCJWM8JXgoKVuFIIYjEIIfpnP7NWsukr
G77ZX3YXgk7MqaoWH1PGoiIgoNn+UgNvhZaxam0fCFCKA4dRL8kAEqHDX3AJ
aW340Y3wGLTlUF6wD6WHlBEF0dYwZzG3hLoFxNsnu09hnFjLItPEaAhyvEMp
xgcbp71JnibI9x81dR/a6q8pUEKDB/u7bQEhZa/Tlf7kMoJA5w+NgvxUaWuT
sQdbIlP6ph4UPD/45uwjNKTk+McxGe/PYZcIcArxSI8Cw24257IYW4kTTyRB
uPz4hWBIr5//cTB2EMsYdaTxLXkX42TTrL9QOaJEQTk+ka1EDYci2bouQyGq
Ia6maLNdwbY+Fec6o5nbQFn31GaiEwM4sIrslPh0hU07Cs05V5CtJPa7n8Ad
oxiuOSXpbYbMVAiIEYbIUVDgHOBucNZ+E+SC1RC0CNMnNQtzvz4ZjKl/hojh
XApeVF2yg1eAKruoi527NpUytTi9lfCHMoRieroH6Eja2782SQCxogIDvWBM
eIMD9g9yUMIm1k78IyboSof5Mq/IMjGYpHLTOFiL7W+yu8N8pcA/L7E+JSDe
79KWFLvJdzrdrNGSf+2FMX+iiMzKD2aXOgUEyaJjdP/6KOlHoTAssYRO0q5h
yjmIN013sf6Fo841EfuuKgJ6E0L9NN5bh1bNe9mRkQUlGs9I8e1YzBB5Gc2O
LlGHltI8ZnId4AMYRPSohKJSem85Qf1KOsp8iF96xfBf43DL/CzQkYM2FYNq
MEg/yLiTRCTAThOk1ir0gIZYIqEYtafwG6iuNYFDrEeLYxTTRSVu9p/mgXyf
2tnTOh0inbMgYYxhaymCn4o+2do0J+ldz1Blnrt3tG6uCSg5a5pvRYNTIXw4
CPcEfA8bREkKZV01CAlmn+Gf95q6CbVkgGOp+y0mmo9St9utpzP5fNAvTMGD
wQP9/LsNZiQiKvQt+5LXq05dllGp1tmaoZxDV892Sk0qBc2Ox+KsWmja6BCT
L2b6X2l3w3NrrJ16Q0UoT2g3yJK39fxhmwNh/mr+ztZOrwoKsEUDBuddou0B
PZ/QxfaHuhgF+K/c2CEzIV8PSgihZKQ087BZRTQ3HFKvTLeHb2Y9v4ptCUNb
rXmsc0CDe0rjDKCBRrkZ76kGqFBSG8CHWPvnerR71jviNnp1ydo57M3hD6bz
GVkDdMQ/5TFiLNLMelfunVSH6cZ5hx406DIxkcx6W7859HFMsFQBCll77uZb
CN/xtqD7O464LjQ0d/VfCwsp+2PJig4JOYlDOR0LI5zbKeVGzXqV11ZXZBNu
PqTa8pP16Xld1E/HdAS9i8c2WQv/V4/rWTuKC6oybCnT0Pe6W5RQYNOzB6AX
cRG2Gl2MrhorM6mZLkC6gprp7l15BqniAtooJ4xo9/+DGqimvM8I/OcVQFBD
42Sdd1ltBCzReWcImNLFuHjSqw0VdRjki/tvW8HP+/vprtORAD80b35WXjt7
gG+OhpvN8k22NSrerruFGpcbSj2E8ohOQMgUmD4YEHDFXtEXjBZNcisFkh3b
o7zPxh45SUj9wIKUDS6XE0oCYJcpQbyET0WPSdKZdYrPa7THu0HIgUNqb6+h
nW6dj602Sn2ikSdHyGcdwCKeHRGdTssUV/Wl4qG/K7HDiBS4TAb8DEg3INux
p4A8CdfhtmP21Wldigf676rQSKHWtPaz4JH2AWqCbuArHs+Ayom6xEMQVBpw
SRrbM2zrHnBNfjKKjcbMCebD7gcNh2p5A0MMC+qPhxBFIJzA371HDEproHvU
B1QikQXEvvf66t9EUarHdWPB0K9mLWrr6Er/i8IGKZgVWBuiDbk5EusvQDxu
4ISStlCKDzxpRP0X52k7sKZd4yTldAOW1ruo+EZNvG45j2cJo2ZAh/hlpi6s
kULC4DjPlrsI+TTVgkUmm61vRfFFkVxdr7AiRbn+rJGFiW/aUivMCa090BGi
IJZ9TvUMGDWE6A1Vo0UuKf6vQ3FBTnxL5hJ8eJcNALyFKeYgwn0b0CS73lrt
Ekm54mUXWC6ExUxITNwuL+B411rIsaiIWndppLGHJz6wOrQcH6Cclee12VyZ
xvRC1/JMOn/TwdQAKcyeKymZPXky+2/rFo4hZrFePQGmjyS5bfMph3vRHr6y
c19WDRBck5WLG31MpzURRkmXAz5wWUvncq1OR1CjVrR+uRLKMX1tJBrsC9Ch
CM/jFt+t2dvBpCfQ8hjottAUWBpOvFXI66pX9bKpB+NfzNQzOk/xQ0qwUBO3
3AhrE/H5THdVf9LUp/+muHEnHandp5KYOquPKUGvjIt+1JP4SdBylDB8BSnT
ILAEZcF7XK3VWeoAhrj3kzBLT24viPnWCFT+f1W2OY6fCMv723saTJQpdIlO
h6qNUuCPUX1Gv9IDpMEuFUUDJjcv2piw5C8Pzk440mapFA5fMsolR5EbsyxE
YfJ/uElaSnFgjxBfHRSP9rULWw4dL4DWn2r/QXscaZ3HjtHxdka5Q/o02gPr
bN4HWwL3gi+ssChPnU7hr64rdUKiqM+LaG1Qp/zfDjy/YsGvRR7fMiNU3err
b7IK79kTmUcjNuF2xj0Hm2jyKg6p9ZH9fi9KQ1gatUMo/KQOQ5MK26NEbWbS
MrggtGH28pDIKecREGVDeAmvEl5K8SEuJTt2hDKbgjo6mv8bDSJtIfWxf0iV
jLPj4KfBX4ZPduCUkVnXXg5OEY7DwQLp0u8Y/Ne+eFPblVNXhglkLBqduzJ8
/QW6wXPwx9Ch0GR387bWQSeVTVK2fFzPwtUul4y8e2qWyTv5mVFsbeHBgp0z
4LEdJQuyKqNyRqWN9VYd1DoUg0pYlDp30F7Nex/GHia+76pviOih+VeyFSTD
ehE/2K8m2jhfTqduKEJkko3kW3nqvhBU5gMyvsobrVpZ0dkkwoBuF3nXEayc
YBlJhPD1E8ED3gB1fdvS4qxXQbb6MhlYFy+MqCCjC8jx+l6LtZXdON29j3Rg
swyjmvHIG1J02Nv/16rx/h4XJ16guOO6O7TFkG9Cf/hgsl4HpKfyawbZuYYX
5a8Zf1wciFMIup2+0K5Hi8/23Y3ij7N48t9nDDqg5Bsg2WkHSgNKrFztOz+4
KfAUrtamiJ9EHMB0iYFHeQrMf/0oLngl19CvX/6BCgAwtAPyLyKIHMZqxWFE
ub9Ur5mo1qbMXXOoPCdbodx00/uTsqg09Atl4M3kph1//L5FWmN+HBLm5j7K
9XlLZpsb8hbQW8gEvN71fbr/SuvymNv/Fgg+4R8UIg1gnP/MhJg5FiwdZzFT
A4FOEbNCwlOZKGbCH+D39R2otccOJPXn8oqEMst4ZWKUaz9sc20aabDZaZX7
+JSA0dDTSfjk5a0m8nAr17tnPGOxqDOf3BvqP77BG4suLWTXx66L8CB2y5jv
THoVyHXpraalWIOxMFmPwF052r7F8lHSndl05o9CtqpeOvDp3As2SLMjfU2J
Jmv0e1c1gLvOMg2Cb9pZXTnY7o10dYsfsTLlf3FpN6o5zvUS/zsaMjJk/mv7
hrNdv2i/x3oPQdtCi7oRD2HtDiUM1BkxlTDPxEwpNpCDt8NWUL5aT5JQVYmV
l0BxQM1Mz6y+NoIWji+xiYRLLfKUW3Sre0kJu3ySaN2H25S09uVL14trOYbh
ynNAiiim6PbJQ3x9ig5Ui9vgPwnUX4I9x6ROM34JE2UVOu2JYsI5eQhvU75r
3ppf+X2cjKN1YiBNv5LoGdgGoIYlQh5UsH6JrmzsGB1fb7l341NLCJb5qWh7
cG39WRnOUtBbuLwxgpNUn4UHo8VInaxnxjQ6wh7h1/Ov+dBJ0o3vBjgHINbE
lnimc5qiL4RYFUTeRYG2kXbEWRO7Y5UWCmbzLNdzaO1Ucs/ZQed1ChM1me05
BmAmKXeaCuAzdMQ7i0YrmCIxffuV03tsbfoiJuTZvbGSLutV1kH/gG7Q7QUv
oNF+g1OL0YvhdcxKYynVRem/bSV7SGNiJCW+GS4pR+o1w+EGgEfeTdb4Bjcf
QyQBFM3l2UUl0v5yvxaheLZsnQ9hya1SDyEIjx9tO1sr2hUYmtamWyk9R5hg
UQqn1/4qt8LpiOaOzA2OeSbficOOnbSBpfC7+q3+oAR9K/w6KY7IrIDPr3Jg
rJI3ysc81sCxZy4hk0JEomuQj+RuBaa5c7TFE+lDaY97OJQdG1c6kvGR/jYk
qLi2NPzXy9W3ZLjhOM5mafaaSIo1T1A6NVkPe9CcBzHRITGu+rP9z/BI9syg
B8JiqHIFOXHLwmXTd2GB3TZcaJGaPruXoZocuHIHEDsDdSQVmFRD1RqRMU0o
G7w6jpVth3i1wxDP7gzz9AVYMLSnc3Ebq2WMG27FhILdLPzV/Dor+CT3ev4k
b23d2CoHf5T7RvKCfxbyDbbu+VsGzg3dyLg090ZpoXXSRfZ/UruTniTgfb6j
EwymCNhpnNU7o4KgAr/J4hGbvY6fq4eb/ITwdf5d6wnCRKpclHjbbtz1Z+ZA
V8smJziO8sKB9yBMrmXCPHXqUw9AK6Shkw3fiJYbmT9uKQYJQ8ilUC1k2hR3
hnl90PE4fq8gL3FidZ/W0Xxli1FjpCE+Pc6StHlLPP0uE3Rc0kOu0ku4Wz59
tUzgvZSWNwqEF3bA9ATF5AEa6XUoq5z9vTFzgGlNVoLme6rXTtbzrqu4syDS
2jbGyvz8N5gFZQwIcF7wfnpv1llGzg1XKcPif5OjKm57o13W0SRQp+qaInHG
GDGsIPwWds7K0ellBT+571Au5/+3CjmqPnRcL6WbVc4utSf7xE7/zq8E6cuy
lQam/7tTolbdKNRauSWokFB4HKW5R7RWeOriu3fvV8csSwQr/Dm2wX6AVYE6
VQvtWZbH7PzHkh8DhVSH0Oo5sfFejFR8v/E8cNzpbcjykzQmfEEY9tFMqizu
R8saIX8t53k8HcEUXKD518tsBdaqUqUGqh99bfoPwLg69+MTOcreqjxh1DY4
KUx/7PAIZx0eDjzkWS38sDr8IKrvy4elIhq+Ug8RHx9VvOoqm54LWtA2oeGO
AgknqB0PevnnHLp6NuiS4WFvtfZp+366MPAZpJhN3SaXkWLCkqI4dj5yhGQr
Ex8iHmRVJZSj83Rebis+HqPGOMUevouVagJ8JUnPLsaunTfX/qO8PnHagGUa
KHjSzQjJVnVw4Tq0ZS1MjpH6Re02SSrreB3lo5+7p8ZPiWp5mUCBEJPtKK6C
n/eaRYL4OsH7Cfa4412jeYQqP0h0YI5KzmUOtG2S3oKxeT1Ftg+HZdI5mv0p
JM29EEDy23JEtQMr4c/ROLwiuoc03lZQSWSg0tBOvyYCMpo1yzUvGGLTcvnm
MYG0w/ErrxRJdF923rBPR20xWYIW8Mh7YZNOM4x42i/iJTcMMxF3AyVjxNpC
c3HAzuUQGU42Awn2iWEPvKMEtXZFQw/9dk1RlQ3bUVSYIk4pwkmMLU2nPWSs
NIb8azfaYAYBwC0ExxMc754dGvCJZi5ruzjjhq1O3b1xD2BJlHKSxqNvxqH9
RSitn3n09+0UPOUoOZxU/2vEfbNxmgSu2wpCgTPu/lE/88boavUiI1Lahk3t
f/U1DAUbJl/5uT7SV0jDqxrKSGoutTsUHiIftLPV2eAr/MUsHOlKSKIFi4YG
8wPICe+tifS9Tb4T9bmwZ/KGiPt1a8lgQr9oE/lupI9jWYpJnTg5HeduNfYL
cgSqNdSM/6W2lAMgn71tzDS5L4yp8Fwf30z/dc6FO7pYqNQB0/6QZYBX9ckr
acu5CcWZ8hk8aB+O3PGC6u6jlTf3l6HBtQIGvB2KCZo8+i7Dn0mTLTsBT77q
XUPqQWmMtIO7/sjJp784dXFgLjucN0rbpcybiZmUtU18CdzVIzgtkj4++4Jm
U7t3saEY/PStLUlcXto3sMWm9WiMVZKme4+iEkRZxKxoifPtn5NQNdxM3r8U
3Irc9bcSbHzGjGFmYw+vgyF/zCa3jXRfYvk+1wj8tGFlUGrdDCBk+t3L6T9W
JveKFMim0Rkfr+qZt23uPVXX58ln11xRVFNVcrO852+tOkGlvICi/dSx6OWM
3Q0hBTUgSNvaTCJW7eJOs2ut5ze8POQxLvYu3JynxGGmL0vbM2LGlNqNPCzw
TvPfsE1B9u9HFAhBICc8lABrIAFft8e7lVHf1/PspFRvQQ6Tai5vvUTt31YI
dcU+6hZpfh2wjawv+yTrV2vZIfzOo/9BAeKc3LQPXj28d3lZnVmSclnPHLkI
DIKV1e/nWHXzVp3ZEcIi5zca3dJAo6iIak3VKqVDXiNuExJk5N1qLbDYuZ1B
V3K4JVUuJZIXe6VZsNXSkDo41Txn15tOzk+SbRLsJD93edxb40su6DF0L9P7
7EM8XFYI8dxwD9mqwKpx0ZokFvtnGEGed2gSfoh3jyC1aku39fECCvKx7B5j
o17j4WHjVmWahtkSRpR92v58uRYFwhXKVO3nUADMjJaYq0yZYlppDrjVi7/f
6MdPRfIo585H5aIpO13pV4X+yZqiRcF47u8V7fqDJ/nhMJXP2efzvdK76794
cLPIrX0r7NQyl0fxRtQLpB2Q30iBB+/G1W3jcCmNe6vXY3dpOu3OJJ/b3Xfd
RHNFuu+Rmek4ZyU/LO+EM11ZcOviZ2n/65v4R9L/DwYs+7GgT3Np2Aez9ggh
aQ8XcDjNIqkAmsRuTEKHoX+upCvUUoyVxiXW/UwfR3AfALG40dWKygoKQUVY
OC0qQ4fJM1y0I34/SbRFAneeA1r1J8a0qANsWBgKQH2XCS2gwOid4RspjCQt
PpFS42zIDA4VbWLqYRm0F7P76cAbdd6dSf68dKWd3NpLH2d8RJHBuMZIuaMO
6WOmQAYfglnH7EVMMt9bnijfparL97qkL0OYoR9hG2/ZaEIxFetlGaQE9RYz
5WOnz/yxEChLFgteTX6FjHJrAJ2cTcFqP95NfebCMDlRK9lSjEzzDNL4ZCm3
WT1ZfhnPVFgmJRrxBlpkG3mlbyV3gI9XYY/P0AwtVPBMcuG66ehjsGgga8b5
3jL9+OrUSxw2H77XS39KDA+33IK/88WVz3ruYnJYktm3qwMBbr3k8DIocEY+
PiS/wLJ3tatNlAYen0W1bpN1fBUhC1oMPL2ZvzXtXYFnrJ0Y+iatrhrocAzN
HduzFtHxfX2JkiaQc0lmiXqHOCfCZVAj9F4NRRiWopCtHQrRbbl9S/hYkugQ
2qLosHQoo460vwVYeBbfnlYgAGT0DFXTotv+3bnZAUn9xoqHVBWeikJeRqbs
Nhy9AvlcdkCHM3iMVaNUKhwwMJ3MH9dSyxSnmuNOPulcf29dlf1s+6rnRVV2
mWUGakwXyr0PGXBYx5KaVpAIgM+kbcYQ5ww20un0+RfFnKZDZkV7d5kP5xj7
GzQ5Zvdq+whWQF5N2luQAcA+1jMNIHg9dMPZZSxZ1s3QAC8+6+mKBQyQEf7X
byAAthykDvQ4tFjcbhEfJ1t0GYFSIUkh1zWyT6zTUGvOJg2NcQmYfd5/GucT
LUAFbrIIL+oMT3H5JLAIWwcr3G4YIGSdn+uROP3ha+y9sa4RZxGfaTEuJ55t
NVSiLyK3odfY0bB6e2UZGHBcUbcy6E5AweVelclyt+hNBCsiA7eYJeO1HVQY
ZCPkN6Vo6RFarz/AMq2gpk6K4MP4ByBommhhXb/9iB/2vJtQ2byk9ILYa8NC
DaMh0L9VFo8cl4mRfDYjpqJ+I/6yAit1n7GG1NsSImwS6YjKFNQwCzlbjp8a
rbWb7u3Gy2OjwsaGLA0eZ8C13/7H6PY1o2o8rxpq+8HEjhQcTBe5kjhz5sPs
v7lU1jo8gOtPZ+lVfeiHfblbMnGCHzRU/FrwLJ/4Q64iK+E6VM3HkSjpcSJj
RMB4PWfHi+pdLjCt/lVL890fgQAqyptQw6wUlrbC/f+U8vKyv0PWAB842KpM
yubtd/gmap0u5LLStTNnpDlu39OczlhY7Z1Gm9OHogUDzwpP/bT/nB/zY220
kUP3vU1EBL9pkvT/mFeJbQ4j9nu2YJLf6HYi7wM1F9FGClHbzpW2XKTmKOsy
5csaRrY68n2ZkfQPi7ezZYWV5tVzN2t0eQdog59dOvGtZJp73IEz7T1o9p7K
/8v3laY51YI6m4aRRQtf6FM9D4q49Ti6T+p3IBqp4W7ea/eCXzUkaFIJp/J5
BCc5V7LyEuUh51MhY4cg9NS081LSen+2qXvtzAuYYQ9Peyku8lAmF7weUe9Y
Nx8avRxrhuR4ncemhkoa0Ppm6Kyvb2R8zlH368m8SOklB7SSrvw0EewCRTVc
F9PQYK2YbWiv4daWsTe4t05ndQnXERVM3aHgvfo4qoFl4vOms7Ixa/+Vkv+E
6aQ6t42vIkmRA9w8qGE9xzm1Tbevl3YNp1cGuw4R8uiSIm/WNUOimIKUEvmv
sh804UfJzArVdOvifiOsYqZojO8XjQ6c3nmei40+fegj3NZekMxixtCQ4Wqb
s+753beDEvFJUPtfMW6rDPvLIedyccFFBDP7maRBiBKqBZsHjbk+BqdEQAjr
1vrZyMELf7UMQKN4c4vfeYFgt8RPzAk32aX0JKYQVF0k+z8b2z5rdwV+TFwN
m3HlKoLZVxdZJL3Iu9hGyR9Ptg00oI/yIoMPUViz6k8xABai9E0QN1Y6PiOg
91F78pl0AeS1Ij9K+EFmf4r9d/byMZbNVgU7QX3jAPo28kGMbJZmodBIs6kM
cpxnl0JqKXd2Q1azxpyisVoanAL1cZqX+qqpuSsM6Ssq7uqJ1a/FL5r0S8aM
gKchf1BFowdtFSya8hG5RVnEy3BjuqGgCKr+E9XhTLjahcRQNzF6AduzzdIf
XwN9RziOOXsw+BimTy4vvucNGq0LF+7vjfIBVCyQZ6putLYKLqd3CfbuUnvZ
pQpcMV/JYeh0aV+2wZ6zlr0RmiyZISwDH9JGKf5OzuxkExfgZIz26U06P/s6
xChusmP1i40UMIg1SH5rKGi7yvV1/YvBtLVc03cRtUS3YVQ7H4LdR4LH2aFQ
3ZB3A7H/eGqFh1j72hQix3zFwqjGP5vSveikSno0nTkMEmuwvW+qWSfSr7bi
5BvSMAruHkfoU+mJvIVtmD2eWJaShJtzvjyhKBsTnG7+AK4SQDdIOBxvZWh1
b4LN8efW/9WGpYysQyhxj1tBkTv2l8X/Il0F6xii5S09tjh5PA/MBKU4AE+N
GAwAWgrRtCmsTtkn2dMO/jeo2C5GFuUtbxkFvraK9Gzfq60Joi++iBUYPx5T
D0BoNvsPExalMWKSqyu3xJjQPkHzzhxMwIk/7ethE/n/MDMRshD3GLJa39hR
fnblusebUdTZk2jdESLVTAzK9klkpOzBdZSLnowuPs4x0j6ycGypVqKu2S3d
UDTr1INknSf8Z0rx9vpUqqiV+E1ZOjBpKGe51SuMGwynyzEouK3/iNVe0mfM
VAKz4253xVtha9DBRnnYK2/FUr12dJRWfkEsdKfFRUgBW33/bZLeOXgGf4f4
hKTwp8zgljhi7vJXI4w2jU5DbRdntGv9WkCp6VHYAFwzDCxYhVrjqRTk9jmm
1IzXg8c5M9cAw5ogu9x7JKREr0OZiRKf0t7g2kGTdKL9N1w8FtqYAzHUwsms
h20ExLgFQsjD7yomt78JDvOXSGdIf1qtKHQlW+UIcSm8mvVxnfLHOcfo/Ezf
HCodwhhxoiB3pCx+gKv8pREFxGUwTN5I+xPgXcE1QamSxQ84Q1Y3gaxWnqAx
80WIsi5ZFzD13xTb6MpCK1CgVQ41JZlnoC+u5irzdHcmpvpSZfDTbdpjY6YY
2ciypLzlf0+2yxBCMAEqfZg5+lW362Z000vFVeod61AcUGDg7E4g8N1ODiGZ
xAmxDZtc6vsrSDZeBChTpFUbvvLKTeLki1n/JCYewupdROW4ihJEqBvxsrix
bnwH4SLbtDOW278ihz9I0DfemdET2OJsG/lyOmGDjFbBvmLc4q3ZzkOwr/x2
l8Yqp3WUKDzDOc5L5+rsrGko6jgfUVgRpEErnYol0582nHAeXCbE5hZXRaRd
lqLDVnN613QEmQNsX67P7zApWKY1+O93SAQosCg/+t58a3y9IYvNthUZO7X+
Hmphg8J/zpiuYJ/DAxzxk8pe1VF+PGRvRTXZRHR85TU5KIj25SLK0kwlijqm
hSMvoa6V/icI66CJhyZu2+ytQJlOIoXAwAWwy8DNXeqhZyanhq12emWO0HqV
+IqtAtgwDwhhdEIUpsIKxGaFxs5u56IH4PJ+tN+mWncHYMkd29yGs027EVRJ
6i4leTtb2i8oi71sKK94GrP5CeUWkCtP7Bu0R3rKG7/Pr7Mvoq0uEZf8T8mw
dafvx+U8V4losLhcPQB4bZSUod/ecozV1gfRDEC9k5WXA7N8uGcp9KqmCI+c
XX1MTekakadaffTrrFs40vQRgV7m93KGZuIzyXH+FQIGHJ3eUJi3w8CzhOvc
bfvx0APyE/z9wPmOO3k7CFuEh3kJQOR/joKnVc9iwRWxTq3uIX4pt/G2tN8B
XJuw8SpKpM7ZtAKtHn4ZoCrZeBUvq8DpM7ZpAmJQGLtYFZIlJ9iZutAQIeCp
yplrIkw/YkFsIxtDdDanONwVgdzf+EUD0v8Y4DimQwK/LSi/0/txrFTLUEeQ
8fk47fLPaDGUUv7q8N02aMdBpS6/0Yc2vMAAcBOqmX3AYRQeiveESJoXDEHj
wqMPCymPv3dvI2DSJlow9maeu/N2+/4m48q88SnDEjyzmz2ZLIdYDu3j9M62
6Pha5PMci40fkBlbuc8w2BE0ZP3y5At6E0zJ8+Upo3fwEftidlrRTXwCscvo
yjTWjcn3grlmmUhiqhXgxHVVDQQOomVGPppGHIr0GYxNk0piTbiYCsmkFHei
yAAANkYusBsuoHmG9OC3u9IPnjs2pikW6LPYRXThqrutEufqDSk0cbDqpq5h
NNPVBNtbc/s7yyluhHbWdKwgGuJafs20IvVDYlSFeKLRSHQuzh0deDBfUZjZ
pi8DaYHtahP2ojVvRLT59FnSFTceBV2BBg1ad+ktK/tXPZyCaXfk6xXQKNAN
SfdQJtWcSRSHE8n+y3hcEF0+2MwBuLiNxe+Xlr+BWeF5wMSR37tzUXwIQgl/
oD4QAVh38w8f/grUlD8M3V47P8kOR/ZGaj+Sbg1Jxg+nIFqKKhrJe1YWPZOD
pNqGhmmvF02uzIYK+jw/xpdUCRFU1ZLDaUE8mG0NTBA6pVhJPRbrAl91lMbZ
EfYUFOndBRjaWp7mcv2gBNPDoMz88AXSo06wFpPKvu0n2z0xe+/lU9h8DW1b
c4BjTqYSopARKsH875Qk3eGz8oowk3APHpCsXlFZo/kzQEtKuPAe4m7emRYp
kT3UbRZouK39t2++fZOEQsPCdxSzC/fyeJNJgSlIZNpuSMM25xoqsTJEMU5Z
aSYKQFbdo72Yz3pq+a2IsLy4K9RYsbuRHMw04dNCbiQuTTOC9TxGQKAGgBdx
BLXKeU9qn9rWVw7rOZo6Ix/aRr8MaK98lv+YgfigmQk7+LMQb5CQ6ZF7h3yH
LLjLk84qGa0lxTUvwZM5b4tjq0IE1NtFKx0gSgLhklPqKIklhP3A3g8JkGxS
+U7fJrbXXIkv+kDWAzRM6xSSXqGprfC/kgxEej/v3T+z++WiBZbH/HYoB5K4
4V4Q7OFcbd08JGmPY+Akq6JVCSlb8gZJZt6bDvhR6w6rQCb7HMJMz9Z4htZg
UbjSFTE2gk0sjZk2phFPJVhsmaw8wW0eDCNPHe8Nya7XvQ3YTsfpcuRW5d9m
iMfxK0d8CwLXDRf7fazman/NO51/t1QERRXPCVdOxVverWLFXG2kdmzXxcgQ
KLoZ46lHjfXB6zA1JKtqV7y2vZzjDW0322B8tsN2UrZoBRYmPjX81c+oiFnm
8KihDxU/5hmjV0UAI+IadqpPW6BSWpQExbP9elplZsBRVzuQgkq3xqhx4lPo
gofs3XKKBGhC95/16FAJLACOs4oowHwPeUx9S9SJPW9i828tONaHERaeXH2u
9LY65CrMJi56/xy5tT3KeWWDgc7032BkVDmPM9f3v1WowuS716ZJ8UtKcG3S
dJLqx0tEQ2GlOE3c78jFGYgmAdLedFUSR+mdj2RWnd0taVoxoChb03AZETYu
udREfYJ4HEcEjTYyH+r03RGugtLXeQrKEJCH2FG8Sa4/xRnF99TzuPJMgr3Q
BefHQi3crlEoB9optuS0X+Ny5SYAB2K38wCO9FclekzRPk6Coc3kNdz4/jCf
qqF5bR2i0mqKjGygrLVIvUR67bF8xBO0LBbeCcDaYGZ89Vml5t9mGeL08wCF
zpXlyg3hR29srpTlm6+r9tgB3f8H4YXra7bQOtF7PVbdJZj2RcLiLyUJgx4F
D37cLzpLi1UELWJbfTeapa8BaWTNSpNzlrw8VAfpoehGP9x9RITuHi40Kfvt
SmmnlOJDHPGqH3CYtrjNlmCm/GgCWSG1+vVVqONm8CYhXumrYOAij7mywA2x
axWFVNJmpLOyuoC2FAvSrbaovRTgZrefGb6FU/qqFBeYOVpGPRnY2IKdIPJL
b7SGjxzrmP849l6b9R8RmehtoMFaSmLw7xKVJ7xrXhxQGnliXfGVh3+gOG85
RD8nc6h9KkRGqRtOUeGcVmEpxocw3O1g6FjWB2sucz2ZLYBoOnkht0z8e4eO
+N49IgNpsZGdxtKQvZ6B/rx54uLrY8QW604P83tc6maIGFVyJpqzlbdCLWpl
eUYlWJcal4EuQK1+tBnzJ7Hvu3FLHqd5DsIDNMqjYpQJhJIihbOgzKOKXckl
dYQS7Im1CI2JTXD5FT6gxsSFjss3QwXk0FdbU8TAMUmwNzErtU0R5fBW5j0T
1dlcF35WMB963lEeK+dj8q7m3hYCzxFZk7JdBLsyzY2IME6Z4eFaXWVJHO/w
Idtavf3jQkgZIZtsxscKu4W9A4W6W0aNrmvXKIOOUcGmoJrwN9JNPadnuSsu
imuN9I0G8j5P34HlM1ZQv6+qmeeWuNzvJijYlYeW1lIOn0xveoHbw1YSnBkm
c09tq+N9s99RL26WWTAciKweWP12fNAF0E5ZCpRAZIbanhAhKnWmy2yJ3bnH
TPaeK4vx9zwqOnOC+RZ/PlCSyr4f3wh95psMbzd4MuBdEGF0WMKh2lAL4tyr
iZnjbrdvVkwxYsQsxb1vGMg0eaOP5ax1/hjmoFn7Iqep45z3NTp1yIqgaJDu
AjK/Q4zqyJgSvDxiQa8/76PC7LXAALWfRwaWS0XFLXcmObdpqvwUaHV3lub9
J7X0isHiB9CjYFNRNVqWG5RWfb/KMxrb7cibbdWB76GEKx9+yENVJyf4RKoD
3cy80M5RSWGOEaSizoa15u7V+Udx8YUoXDaDERtCw2k0C+Xnw7hRTcuNZVQY
brdBScxLxH/AoB6ThYZaw+7z48y6Z8qa7PIe/B0fR/2oBDTBos2RgstQ/UHf
fYtBVMOP1LqkAOA+v2RK31F5DtLyJZfUjW9j5+hQ11y/zJPtYDqCSrxL+u1F
1EEoaC39VA9+wHrtoB/gHPPwXEd1xlQ84NnzPTu6jnTIttUDkmfAwYVYxSEM
bfjFtsds9YzstPm9yCMc7dJWYK+DhEk7a2MlveOb0MnFTYChD6YlEqn5k8Hn
6cemxlNlCI5Z3giI7IJHcUzMmmD9kmWsGCay8KUkNQhlp4AZe//+Z3gyTfSh
Pe8PdZwl/mcArj0D7j4PJjNIQtZvi2F0wbAN5yfF1USzuS6wquQgY8NCGtc0
7U8hoALBYD3ZzGFs1N2/I4FQyJ6Z9FNMGOw1FsqYfeDnSWKlmHf6yfmCnrx4
bkSFM7fjufVikxJHkxsO+meDZ4S3QOfJ6dz5j+lXSOl8BWfnO+tjX9s0wjod
XI631s8Fw9c6V7NLHEIQ6yNhqlGuZxjirRyBz/1i3kLfUNkwNwkA/sb2vlfT
/WtSBTUE1c2HA1wLcORDHwvzmXA2edjoR4sls7Aq4HRp3wsaqqvGdouYSOHO
zUC25DEDOwUNpa1BoEB+FeApY+0nez0zwT7YxGzOpn2Ys6delAWKcbsjF+tX
aGgAF3YejDiyYB3m1L78pJIie2BHSB/4Kif2UEjqoQZ9jqXA1u9dcp5HFHzu
e8aSt+xmjb/GHT6Zv2jBheajIRa1NotKD22thRpwPUJuUnOaT0UmUGyol090
8RjbQI39hXD71As8Ar4jB8TdxnZZDxNAfSIO671XrGwS5esgsD5W8fR74h+M
Eko1wI2ZuJZXzdvC/cGHhvt47pzxxtYItj+aftObv/cPGVwHiNs0kHSkZbbI
bkTUvUCTuOMFu4tU0mgmXraVhz8NWPRf6aCWZN+II/18I8NrEZpfVX93/Nbv
6tQDQh41Cx4yYkvkNYT6CCiJ2loAUuc8+5ITVCIjEGi960Hj6hCCyIjkEX+a
7Mxn9bnI4gtfTg1851jyUdQ2UwA/WaeHbkNiIwOrhunVKshptPjyXZYBUvCe
73Rbjf9EOBLtLwkhPQg47+k0sJ7Kx5/p00ZnyQhIhk/ObX5++3Ad4SwMdmNk
uXrlb6DgOSEIGTsPDT2n17Y0XFTVeWbjrKMrkEKPj/cM4SL1F5uxTWh2yOmX
9lLrBQG9frz4arjPmiFRLi5yK1qbMbtvjyD96hsMlc4cm3NWaDHb/YHBbeAG
rN3RI4zAZHeymKzn8SGywyyuP/CnI/voHqQDc2a7wypx2tOXjO2x+nP73L0X
AJ3fuQU/wPhRBIFJoQ8OwulRmhYzfMm6GpfAm9P0scwRc3CDQS1CFkLg7UiG
gy+vVVKn5dX6kb5UwezhhzOmy/Vu/wWQobDahPaub1KWpF2PM03r2wzKF0n0
ZG2WmUazrnxhCzXl4ZdrKiYq/SDJsfDXnXsk1sRCWwDts7Gs/faogW4k1124
dezgLbwHdsuKBIOVYpvdTXYARYnpXOpUEPFKghaFx9eMQd8xvJKaoKI+OTub
WhlBQ5APhBrWRhZE3CUOAiewZR/jCvgU6opw0dYgEE5VrZ1QFtnAyZAzW71K
uewiOCrAzjWA5PbjjA+bzQRG2ZHliygXd6uulmrP1gRGrfoJnO2U3UztJzhp
MzO7TBlZq0jj1X8B2aoJJEDPGT10MFYxFu8TlVi6q3ZFUlb6qyo+DNcjUByN
clwqKQA+06li+o+kjesqCQaebvnv76zvaDWeu0uaLHRlLQeqo4c5agpVopco
m4qycbAgQvut/DY/8z3ZNjQSOnEkIdoaY1xOZagJc7piJHz5uKDZwnlnl78E
TTUhl2QywPorA2UnDRJ/4eaEhDuBKeKbcs3B3QZjDQhkidmoWie/eATPJO9d
32Q4zM+Fc0CogVUTSOBMLEq7h60j3dUvKlaRbchRhJHm9Rd57TmNNG5Gzoop
OycQNs1X0OrM337/i8lRy+rcpiN1YqXXMp/r4SUALRAuObrcKkhXT59mcUZz
a3HDIx0ePFttx51bnwAwJHviI+LVG39T4FNwQc9uPyZtBML876PFsGipJtMD
3B4z2SRyp42sGVMJiarmqbwrieqCax00sofWxnGmIpP77m5MRjVCU1j7psHh
LpZwCeo01IC05Tzm2R8V8XEMrgGl+7uluPli2Xy3Svj4WQaCs5eg9Bmh+L1P
6/WwA1BbDK2QAyd3U1TiZ7XB5mO/KMdo3ZBemT7aj9sWjXVVbsbVIbja8eAI
WmStWsKcmFLOEY8Pozpgq/hGasimNzxQblv+GfMzMEA8aIvmrZo24E2zxHE6
nZlC5T7XTMX3NaENRVhRGOx22m1pEHjNL6EmdJ+OTjykQcZ1nrHe+XNaZc2j
BsCLvUCU038f7+vGzPse8jChPTPYdA2CnDh7at01153ym1EuDp+QXTF/Xytw
Z9MqJcI7l0pSE+l/wYCquz75UKHkvo3jOCUH/RENvnY8dNbFTGNweINcqq5+
cMfBXx1P/5eBtvy2/jO0UpfGFU2C4VV/aOe8TU7BHT8PgC3077wDZObGRb3z
bCqRmFg21E4gXsQ4tczy3az7/7Xj27Cv4plbB2JnlCollxWaUPl1BXQWD6ZB
k1vFpW2LOEBmWx568woNRBWNprUFXeA3CO23KBqLp/aFcA6EsPmzwPvi/+95
EJOaQXTLrdG9nxhA0LGEhjoDBMXeGh+A2V8GlqEbduvcCgk40pPSydVKtqrZ
D7xYCA6ifcrAg475vqxvVGO3Jajxt3JEGYXkPXxBp01B5or5+3RCFWhIthfl
7g5yXE+JRR0mkRBDmOlPBG4FSD/kh86IsO7m5CqssHtiCFIpaHWB24R5xABU
6mW9Euqr1utCyWeGve6NDXxSOCkAQsfDyBjQK7PoUVv/lF9AtT8jI7Z7GEUt
1HhJseY/ssv8Ku+RCVnAW+Ckyh/o0On+Kl9rF5YhL8MxAuqWTTEXFeCkVTUV
nxMattMKXxFDEZegXNYUwE9vdQxMqh2wSDjxnRpw87VZyMcP+9WhKCbmlCqK
eiAalq/+uNFraxP8a/HNPbIXoWioYenU0y0YTRro3Utc45CiATRc9g7k2ovB
/Qu5XLvyfpx2ELl4+nVbY9zd0SAWQVgk3xmAUbjBqKez/ThllVepv2gFiM+T
8RuvgJulOZqCmsVzhSVutIT+QGxXa/On0uYgMtglLmrpzZMJQjIAr2sU7nSO
c8RdaGX8Guoi4QR8E9aVHK33NxbUtnJPsNAQjz68X9JKSSTq1GnWzmFLmkU6
pro/kY83lNpse9OxtUuPadPmcdp8Jce/hRG8LJbuwSMf1/THikwWDVE7lKwc
Sygd4qERTnu86HrHHH7i5M2BruBbkOefF6pcCDuxtTV05Tua6+jw0Aa8XsRI
WihQHsZScrklok19Wd8fSIhsGNzYTniuVyiXL3TSXlY4fKtbkL7TW3Nz/40Q
Ep401+kiKv8Sd0o+VTMBdrFUFeNPHIYVbnwzQXZs6/bH8az/DthO2ccyufJ6
TdzNq09JUvQnM0SAQD8i5kue0cRy4pOmAPu8docie/1wBamcf9bFopqTxhqm
DOJ5x8TINEmzfHsDhplHArGsSf4zS3gGvACNI02Ymtr/OCRFbUmeljD2Y9Ls
Qm2fxLU/Maxw5g40QWFyXEn6ng4nE/935Y+ePUfhfujiKCjpHgKRJdXIi2oo
6Bo58XjN+ZIfdHnUT7htK5jjSElu15Ulp4MtVy0hG6hsE/cqjahJn79HEGZ8
5jRv8UT34tGM6XuD+DVn0EPan/c7v3zWWfHzW4KfwiWykVjJA6Yp072eHtkI
au9CluKHYmHKIZbAhQQz7lQPApV3LjU2+v/SOG7bY8Ymbt+fL+ynarSrj22H
NB6Api8v8+5ZVmV4CFNzK6sC+/swyDajDzIDu/Z6vx/OkAI2hj3zrSrMA0Ow
2qsH4F1tV3uRqmDddhabIXle7+XJGEs7sHboJzhDYsUcTRujDEQKhLrVKRAB
0HBf2DGy48HMSphSlhvAQSWnEdCeSs1VMdm4/5eN6umKkLIfFsYtmR9tNuyc
/sjM4TBNwTW/pNad9w3HJ+JH9lVLOohtuwjoTtT/YmBi8gBIHjV9V2tHStnW
5uaLEonME3PTpoqqzRf7W7Vsb58gsGUnBiWINZPnsMsKBsPaUOxZt6TTSdE/
wfdQY6tiozjeSABR7QAc2U+CB8X3df/StyGf8nKJ2HiOSJCGO9UN7VP6LpLP
o0X3FcoTOicFrsuXyw9152NN1VHvSg4QOBEadBo2eQHW7NoLRT36Xix4New4
hfWXuYny48l5VHRKS1eDJacPaAa/ytgrhPRL8VrI2/EHQHrcfYvPDwuyf3UH
Vwm9J00dpXABOtzpgqH+4/3Aqp5rYVHS36Zj1NicnH/LLuGjhqu2R2jKR7NV
O6B2lwrh8aK36sNcGXBOcoCK+yY0ZZ7NrhasK78dnmRCXdLW/5fsyynGUzuw
9/qrAA06znBbQsaYEbASpdW0VxLCeRJ6kkUkKe/zTnvxAHD4ughtxFV2tY4F
OBdVO3JK6WaGlWvMxhXdUETk1uN9v8GuqJTJddXh1+46tvWXhwbRXIR5veL2
cmzagFhVWmuWds+1XjRXXC1LO0wDmdGN2Ro2TQBtNQg9M+y7I1SBSp/KpkiL
+eoVt552mGx0esdwn9fGmHhzBsiALYmAkgN6tJxsJIz1JwI8gCBYXb5TkbiZ
Mcpg+XpNp/iisrhSZcIjqomznXBRXDiq8Rgb2LRMsAvTSphCl5fF+dC88QOC
JS0x7rR5Kydus/ZKOwZ/Cr3YPxY3wttknJHrIdUP/8e4k5adduLmG3HhF/a2
6ZurNY8yThgCJtO97Jy2HyQlJ8ivLFgJUjGwTJtXNbc3O+xRNKzt7EkiQkiv
gqnOUCEirujC+N0jhCjlieLZXFT8C71+fOOlJk6x7rUokD7N0JE7a/VOgjAG
uEjo7pyQ81wKX4WQOSLW+MsZkVzaaJd2yzvKELHC2+fUPOHUKFiZ04VEOdsd
2jsB4vBQk5wEwzzMlXBQ2wwfRALUObIDfYo3c87vYxiOVtOJt9nyUG/uplKD
Ym3dfxcQ+3MwGBrU24LMUPaUgPKbWZUR/SOfUQDPQwgBcEmgUtrXamlmROk7
T6bMtoiV6RNbDg54ooLwvX3vqo/Eb6QgORJueLdBhADXIELQgGMpNdQ6Z2K6
wAbT0WSwCdY0nd4sEP6reuuzopwPi3mWv+EfNxGLl0jtOV43w59ckcZ1Xbyq
jBjazKF0wAYzx7pyTOur0bA0KkebGEbHzZiHZz1RB5joC2R1waFz9kZvyiYB
TbbwSkkpHcj+foMOJ3W9I8l45dB7qN264Rr7az0KhLatrUmL+eqcsYCXxD85
MlAuK7+KlsLbBOOr+H2S0OjO3Z/1uzxVZFloKakHyrhL282vCvG5franbXXI
Wz7WsZeuDujrAKf4l8/owVIKaSVllImAcI1/KDzWY3xsnTUBS7urRBCyXaQP
PKIOxCZG3ZVf36OQj5vB8LQYxzbdgsT1ON1GvKf2U0fPGqmtKtZtkI1rVByF
rAM1apf7tAC5G37VPNeFKeDGzLJftu1QmBj3c+pcBwJnpFxVqwR5X4QGhuzT
k9qG/C2m7XwTKhcD3mfnuRU+/ubBEdEsPo9OXNw06V5bCVaGaXD39/Ml/xAr
nGzZ1BaEQwvsY2MjCmhoPVbma4UKRxRGLQeBg8tnyMVGupRLdoeFSW36v+91
rBdY1GY/kWpMYAyLlsrI/AXFovWlypp9K/9w5dDGeca6WEl2Xp2fi59KTxmM
9FCg57CnWRWTR6EknX2Rtx/+16OwkBlyi+ogEhY7yMl84ZtRR5RXjCsdKVVF
l2blTKg0Bb3jQ0OqNjmXR9k1qzePRKQLPcj58rzlbixR8cd8+CwCjJIUa5Jf
gOWMD0ChrvhLi/EgsUI7Vfe6c6tsM7Xm37mZQBk04Foguqy5qfFePGehwcY/
vR8+bIpyUZGme3gTvhHhobzGx+RcZmrV3+kv4QaX+x70mbvmxeAW/d+uekf7
Aqxud9h7TGPWQ2KBdJPw9cY2Sc60bPOfuP1jM/WYZfDZ3GbkVP1e2GJ4RzFM
j24yZBBSKQFteTc/lfhTSjgfZzqeNuDWoRQ5HVSC87oUkMKdPogwhpqNSs3u
US3gxdaZy4UHUMlNmwTCLy45uqAPzvN73zP1cIGEk459kkQnmmsQCV8OD7Sj
ttoK1z6uG8I3ZXCfW2CvhBSSc088ItVKVo2tEkq7Inr4y6km1rX1j86bHTvk
v9raShJV3mngl13MM409+TnMaJarfYZGes73IucPRHwbSp8Pqx9o9lJo/mFj
OopP1HPR+iAa30OLeIeaAEJ+wr77NX1APa2iq1j6DTe9wcM4CZ5fx3evmdHt
u1mcOfsPRKBfUc0ZxALKP8idfo8gMhQyYb2za5KwPEq/4778Ig8bxofp1oLF
HsTGYX1IFr3CpgLS1LVTwvZWAHFJCSYmSiMlYN0BAq5Vg5OOCeZ/Y3hCm/fF
jJgA6c5tXHLqnRUohSNQXplImp1L4sv4ocg6oFVyYPgfvOgwHR2aMlaSgPvQ
PUumBJub4e9yk9wESnfa/tDJYN5m3JUtl1HcdJB/bua3ywqoPw56e9q8/klV
oU1JtRvF4IUZvFFQOobStUu713ziGuTxbuQvEYDctnVYEpBs4XbJGDI+uWwg
1UrJa8eTnmB7H21LOLsWEixuGJoE4IlrDYkeLkFRMcPPHWIRWeQODaW3xl8S
Qh2/qZ6f6K02x5rNpnkKAHrcf6+8lc2BcGWSNmVM6zyUyY7ma97FKooE8jTX
59TFcXBelcLLE4lTbSdPsuDL01VicoHHV2u858k3+CA9f1iG1SF7+V1W8h9k
j1cjOQHFC1sh6SHT5CmEZ8wAnDvDXV5bsJqtjbOc8SGdVqgPf7qKxyijVT8K
ZjhmXj9JsDNMGnP9zjTanLgKtJVSglAe/HEZ86x9cODpOFJi9Vlqn6e7QLKh
g6qnUwvMwFOx+GSt7IG8kCL5KpWYxGq0Yvdw/0x0UPhf+1YyMgNnzB5o9Zvo
enbdMaI23HdIK8m2wz7RJbdnshibhpmLJ5/X7/46UrMoBd958EACKGmZ4VZN
OwXG7ntdmA6AbyQ3hSpSwI2aZWIb3Gw51STgQZIj5xv4pXXyQnR2yghFgZHI
NhbkllWyJjb2zBCq3hAzN/YA5Vw7P1wPCpPgt4oUBKS554O4vTBt5n10+ukY
APhNasbhMV8/DN2ZxE7d9q7G99uXFhkzS1Jh1T9gcvY/OkjDImj+iTHvwyZN
uOIoNCqYkANcPIUSp1RZPqQeH7hM+gAWNsV+NNK81BA/oxG1Vq77s4j15p+m
7DjhBbedA5OTLQNKMIDEifqpHnXZqpynMXoB02KZH1gzKUxW1r/a63uIjbEw
POn5XM41VL0MMOKrZZ84mripA1aJV7F+aolgJcLpKPURa3Op3p02zehqBRzd
bDLQEkikfCF96qeaF9Z9kJPH9W5lL2uXpjuMKCV6/7apeg9pHprSITXnmJe0
4qUhfgQdutrexIl/ESxsClkFmKiPn1y0TaYwT0XeaEfy4Z6Ole3f2O1s2+n8
EPiF6FTEFKc+LPKwHWnPt7NTBQu5Gkb+gsZU+fDOI11oUJN0q5F3d7xdeOcU
Ia+BFICJCbetRh1u/67o3Ft64J5/PgKqwWdT/GdOWu0N3u9t5sQwb3DTIQtQ
wv/gVjwPdPrCR9LsybFtcumHNrK6EdXayawuknCg84BWCET+Uz54bhHzPgfE
uBq4QXB0sGb0cn40CE6Zkar0dHvDpeATcccPBQIdUs5zKAj3O9/JIahms8MJ
p25/DMmvqlwIAn7GyL/ZCbxruvC3L0PDXbRrCRsBRuw9JzlEyp8uUTTuv8fB
4n4oIylAukH0MSEg7YRFJAHV6w3FnZKmdh7QkQV2FszdpCu4qgu8BCKX8cCU
mgL/BebqF3KdeiDapC/MoCFOGQEkbDVhKyHXlDDST/f8i4G663I2oFZ/9/66
qXScpi3yhCBkafW59en1TEp0jqWfvue23wtcoZZePhEqnwJgMZXNyG4CoaXQ
sMine5B12/Mz46whPlcn/G8lr/lztXYiJSbBbf/E56WjfFAjFkx1kzX0ndPR
GQLuZzNHXQQtQtY+a185Og5VDfrWsU8hFvLdTS8AryIaHZFkmUlAks523Xfq
Ju6SMtgVji5j0+GWfNkjEbHiYbCuKwJbc7TaWiKbjzw/UyJw69yojaeaVzEK
KjLjVyqySCD1zLSGbPDpsF03BPfKB9mWgSXceGeTr40cRo9xZ4It1z7EA4/5
bSEeisJTL8DBrt7ahgP6iHA7f5kNoo/Zgl+BlkrsMWrtiR0mEVSJhbzGTHCO
Bxd5qyhKjM8K0bv+5sLIm93ALJjByZEKKvc+bJnzDYppW8G/a/xCfw0ZBSZ0
EmXemESBxpL6gcDC6e9EeWmwMPdmyRR70w0D9z7nMW72sAXg768wOiyKitB5
0hsOgadNzZqFoxq8sqNPE5YU10TH89l0nhvunlIcocHg5WCoTkcY1/3xlvSw
jfTCy/jDClJB6xbENyKS332BkV58e4XEfArKSa+OVvd1pFcWDd7Kbt6rA/bh
69lEp5ueKLyNEgUjGZuna2yKz7LyXVTmOiGy6vFpoTDLfRX0z8+uVafVPkDy
ATTj6UWHlMCNJQ6Y36fAmndGdJN0W19fqxxZ1tbtEBg8i44HQTTZjR6zXzXS
ca5ZmvmhRynKAX17/TgaCSQA1dxW+t9uA/mdWCxBsES+kTA6cSMmEfwfsN9W
YGgT6uMmTZmNLSsm1Ju+Fxo3J47PQVKBFEeKl5mnbB/6NTFqMfnC2xnFnhA7
wuxYYlI+5Ex41dX5YeKffvOrfpv/T4mzD6Jmo4dr59kOEjO6J0C5xLoANjNt
l79E516S+CANP4ld0CF2nKm87UE/8qQYZqiC/XSvXvyIPZyPHEDzvHuzdlyl
UH2SqB58ctNVwof2Y7GNpjG+aYHF39SP0CqoMlAksIOsGk6La8bveKzIboNO
UWXf2cTHNaZsBhIwSuFEHR1IxcGBI+9pELzM1YDiFZUPQcL8Zk1Cyf0W1TCD
KtnDCUQ1ScN1utAzyVzJ0s/WtjTsGpQntQpbw0e8SXz/mtnLdCcaPJYZb4EC
sCcY+K2LhA8l/rMipbkOPnXdlyVPPlFJKnz0ShecPya9qDDTasUrzXQELKIs
4nDW9LHZctcHlH6wF1lB+449eNkB0MRo73zHoQ7SXT7nniUzerxAaPShQz3Y
CridKGirYzdAkx4cpu9m5m0zRA9bWKIii58gWeX5bvUEShQWx02ry44Iz1tZ
1JIa+PQMWhSB2qwRsyD8UoG0UPj19bsLRhZStkFuUz/oQhOscZcOMsSRcHwd
/tSl0rzJxfqYw30YqfpvR0NavQ817ePw4YxiRkFq+83nM8hmKg0oEGO8JAvB
iqTSioW+2OS893nyoKTpBFu1J46TQFWbzsj88fs3/t1MbRLojbBj/fONAbVg
4Jto36SPQBCY/o/nZkxW8Vss+3xur+zcWOWh49fHZUPXxNh92WoPRcrqeOz4
zqP6iti+hdXWAwYL4t5ehtI8DtytLcaTm2eA7dSDr9AkCAZSTebBK3+x4LHP
LTfYFN4nOx/uukwxNBmScbjGwm4JHOkXygzEj+Gi4IYvrfksG7B2lr34rIYI
pETczPEUkM97obSCEydBc3N/Bg9GyGc9M8uPgKnqVyXzhiUX0aqETNl+chUX
QWxoj5us35eXO5GkfhcDPgR1GgP1Cpv68VO20In3hqk4vZHHPOSr/Xi53Wg7
A6YboPZDKoMpFJxnNWSEWO4Auy4ziofIrCI0KwAxy6Gg3pInIIJj82CpVR1J
NZeRWC9j2QL0MaFKUQp2NeDY1vi5/rQHnhOofWagq0lbccYUwMgDrgRWAf3M
qOMx89L2h1lnj1gwuD9EKCKdjPMMT2M4Sl6C6H1qJ1LyBPsKzCei3EzchGi4
5HXkch3sdiLRhDNJh18AyU4Ru24MMTiiDiYMhEPZlEQ0RRGOqQZpsbVD7wOf
YDj8RxXjWiw7tT9UARmUcElSEGPQnyppw+mrs9j+KA/bme/+C+anQ72yaFVR
EmD2DA56/nr40DsntzM9VpkxOm/QLE8D7+mUXHbWCHbZ3j7bNI0A2HYnw/My
EwjPFh8rZUq4FOpN61BcKUPMYp63LIb7rDQ1PyuWuE8jojYINXh6OjAMkroZ
g7Zk2zT4lfbL3n/c2eb+yFM2jMN/PL3zR98HjS3IjXlbluaW5NLe9niCw3yq
9mOKHJtKquBZSdWemFtBKAnYNgxKWyLbBh0MP3joa/w3AaM9rG9rYdnVwx5c
Sm0jYCZCUfR59zKXKytL1GnJFuWKDf8lsbC1MLOaO03NGzcZDgxt+qBI6pEP
bVMYgLZw7W/mUDHvHXNYLuAH347pikNBB8cIaebIHoh9ehIIF4kufirC3JZU
1MRyeSi1IWrRHb2pUoHaapdsw32JbRp9joMpOAghUeX7igb8crs8DsZdkRO8
CbP8jBC3CphB9xZ3FpJULnAV2y0U7cT2B7xZvsBv9X+ms2aEJKIiwdzrzNIn
xhgJU+ZJTm7pHPQTfABAnCrk8j8/czAHXOEH27d4TuvjiWGTC7KvbjJ6cHlN
tzJy5TcaWKEUQakCKv0jI/nE7gDBJ/q+l5v9FxLlLjM7HAZCL5eu6SdXqURr
f8bT8Xd+h3geZ5nPIU8/Hwgz3hY2D7Q0DczDXw6qC98rEPSmSc9GkSDfqdRx
b822jg39cQtuNV/NSQdL7fOo1rd89wcQ6lm4O0yby3YfaPvFUiLxEytZk4Uc
luFdFRGP09a78DboGT3al9D0P01xZ2iEnHyYIXROveHPYPCPgEINumKcUAge
Dx8FyTGbohbE0RiwkwkLwTMWLjDulW+JgLAlxFI0JYh7Rwe8I6i9sWgm/M02
hUZxac1Hrwt4NmX3iv8A6QTkxgL9vAY93B60PPe0absS2Aw1R9Y6OEUGL3gp
cqiijh1HI5SLZ9K2/Cr6GBpmWHje86HpkniZk298o/WAl2lO6sUlHtJeWym6
Xbl7uP72nnyVP83h3gsRakXBF3m5oeg4MOcPzpWNS7GIOztZCtMjrRxTRXoN
FylDjF9YhsvWEagHwPozwIouyFGwArWpCQwVvX6VmfzseN/qfCD0tSCzp1XO
Ff48hImTBv3b3alySVqQP3eJE0bo5K8eXd1+045hyPVacv4b4MYxV1Mj5yP+
G50BOXkFZHd4zq9jcB9Lt8mfb4srkGhyN72M9VlOSxXLwd5zXoEuMn5PwUN6
7Gw8hkDEctb4Z7ho9HmbuTgpWE7/6PBBRgq4IegtvtiLMYkdVSaU/V6ALNDT
KTeddMLR8Yj1I0XfWm66W4yKJQfaqAek+Bity+hm3tCn9Jyfam9Kylwk8QLe
ECE19hW0BskwJFA6vDKzCgSP2DV4UYIm0uRtEQopd+tKq/EClzY8OBTVZnZk
Y9oTKGE/g/6FsNurp0x8YJsC9kWcKZxbjOXR7L6VEfCohUcuAVCbRHComPnY
I2VJXMA7/9a1vfgxuyS8GaulotROUY4U3qonD8DttCwShHj4uDnoSF14D8hs
LQ5F1OFyAYXwEdcyAPNRywJF0Wz/IobypLf4LtGDaoBHIr/XLsZdIMXu3G9E
cGKb8wko/Regyelf44oU59gEUa7hhilIuOIch50fTDHgddk+9bfRUeGbLPAS
xPCJtzMZyN/+ZlBnpHTBaPw5VB/vCT2UeUigVc+C//MDL3UmBZm2+A+3q/Tu
2hcpVKSNLLztqcjKPV6CRkPf+5ktZ5LGo72zDxs8PkJ5pIg4IoMv8uOLAfCq
6ph7ZNU3bT3UtmXiZBZTQKq+pDy8cd2RpYyvTmlFAfYcnGahTukGQHRFpLSH
JDjEvIsbR2RGl3Ib7kPGca7alBt+sbCejxfeXHusn4jI98OR6p/GQXKUMAjq
Wns2957S2F+nBfY5hQ8pP0ly/lddIRspQKMzGm/G0OO2QLZ6CwmFNi9mKkdw
BNTnNWZdkwJKOHP/+MIUmgop8t9wKAoJkDDv1+tL9vKxBNuJGdioXkch7N9x
UqNr0nAy3ztsJLLhOinQ4ULOApKDts83EzvSaHxm9mWx17Ht5VC/zNRZhQi3
6Upzlx4XjH7VGauDGtY0tYmPHPRacjssuNQC6VQVHA7PxXKf/iwpUFfI3Qhl
OUYQUqXr9Qy0BScqacRTMPzFPbbsEHKpdHR5PW1UbABCJlyI6rcLCmKgXW4D
ICSnoQpA7zarKigQtun5ntZPMHC+uBwGKUY4lni5ccK6VRRCRt8GCB85r0Z6
fVizgEWW2xs/lKbAXpIqwd6M+HPxjSDCJ4lG3K+VZAbf1tpzkVcP4Hvemiql
cBjBSt9SJ1r3jO+bafIS3UdDc/Tbo0/xedY5upvqKP5lBLw8uF7jKC/CfIMI
dvXOlv7XGhl96gYHvoB9XpI4f7m5vfjonj3XKJCmfBCrNARks3CVQiei7+aK
ORGs7I6FKzi9Ar+m629M2Wgmxx64UFosq/dTvOqoPlB2jmm+rS/eJ+BCeArS
PBGPJbcpeMkXyAAOv3l+iTia41upbwcKWcMz1BUTxKSnO0Fb2VLEUApfQMtf
7FJ36vuMr4+4Urwu2ovDzZZWe7kysVRni97zelNBmCEw/IvZd/xecoFPIFXW
59dkRa86U+CcZO39PsVxlz9y+HAK7OeiNQljJLcZ4gmOW06DdVpOSAsWsins
liH9mtqEF5yrhRag5uSxh7AzeMidNRiCbIgbgC+XKYDhEeCPv6wSB/D0i6no
4QRCFNCYFpaMeEwhpkYdsWyxpN9pMfehcCIxgG+gMfAfwnSoPuLQVXq+8tPf
UpcAuzJi+2Lz3UqwCaPxL20XhehLXN3dIDgR+WctLhv6lCDW3CB9x5sWrLUs
6xDMqjLOCG7m3cccIraj96ZBvecWyV4nAeIjoduHISinRgIbeIDS85hv+cwl
1NERQQMkhjP1wgF0hrgtmhMi5aHft4UA2bXhEzPNqpwF6uGxymZqOPpyfwaF
cZknOEjDBs3pOsbd92itXRec/wk5UMlFzg2J9QnHqQCLkMXBBK0E7h0y4fWe
ToNYjYxoN0g9X36ZFBGh8Gm1Xdx81BUrdfBcMKpWzmYvfWQB4hmD6l+IzbnR
itPtxpV6CIMMXEyT0pehXU29P1EGXnyLX0GZL5Rmo7UShQyK8/NmsGMMzWWG
zRG5bzewh8qnds+H9Y2bQpvwdGOUv64Akw+o7DQEftGz66SIgLjbKGtc/gc4
BCZe1Ykfomu+nlTkXHuI6KPnkJmlNsv2MjGbsW9YAankrY9RzM+m80uq44rx
n+jsM4PjKdlHaEblZz/q1Hapvd5Or26/mUuQcDFXsEKRKY/nJyyZz8ZX6xBq
GTN8cyTag0QQCX1qWSpc26Z1P3qyVczDrMvL5ZmDUUuCwYh1FtS2hTIRXHO6
GOjEEVgvbteIMAW7Z3oWz2f1TfrWNz4xW1yicqfT6pm5FW8gIm5McxPLGp5L
MrGZHjyTxirKSW0MuQsKGWWxxbVnIU2w8ohHctKXhZ8NOJGBT7UYQQ1vCUA+
zJKfkkhZxIXgbSyy7TV5TlCfEAM2yTlKoQ38g3Z47Fy8ioyPq5eLOMY46Gu2
MUNW/PDQAU6IQgxdnWaJdTYLvK3XeU6720842cwG527AVaqkC/PlP/xgaJ4N
n/+tmgjyI5WDjwWdnPfxIumIRrITuIlWcxt+F93Rd1/9cU3LWdBflpnve8Sw
ClDkFmxNxUqsgxQLP/h+S3OIDP+r2B9jRIe7uZQtAJq5pWYNeZqSzwV2UZaJ
DAxI+ov4/h+WanqSxKLFVA3uCwKnDyXlcu8gPfL5ECioO3xfsw7ln+6Y4rXT
oozNYVTC8e6tCF9nRt5eBU9v6h33VjOreoJnAb5Wy+TDxLo/xjcmlRvOICqj
Me1cwRwBQN04up+LjmdxB0dqb+RIJuDKdI3s3VwIySREwXCvHHQVhCHwzRex
orCv6rdyMqCzxki9DaXLHL5ypIN9tTjecDkbypBZ+aia73Uo03uKLcVpZr1+
k5thEkY8HXf6H6KNTimym0KcfA7+eEN6oj/wRn2RBynbMwVMwqcYfeacj8dW
ecLYfR2EB0RGBGZABxHKsLxLDGn3WI8p/h18FhmP3jmCE36bk0xz9noEKtlV
dxLqN7CUTJvBshl7A8WIc4OhZCSMYVxUlMZHWhoI8HGhC5EC6LIJK4DVWFrm
n2L0Oj2x+Zn/jVP8KHrZg2enRnZsfctXuZeFT08Li+Yvfy85Dmpq6vdfDuwX
60Z0XyPTGRXVvwFPTegYDXGjTVY8OaoZRtn61NalH3PJLBlOL3IgEnQTscGW
nyTzZvnNWdSAMtSKEDrcv7yf6LoxHkOnwg4n3dspwyvhWoganXDsq6fcJgVr
VBwcEWZQMDMJ8y/nXHreNcr1i3+6US9Zwg5Ghqxr85zzCaOO5hCz9Fmj2Z95
Id6UxEwJ8c+so1VSrFOdmOw7i6S3SLVxPZQaR5wUHOmkD+4Oqr0X2CB+hDBD
qdv1k7gIT22WrdVBvNR6w9ZsDuHtuIUszizidtnvy+VtaS5d5QUii/3AMvqN
6KdazMuIN1hjav3G37KwkzAf9ozl0o+wWYG8qBeJS+L5bumbjhqgSThirXsG
ZwUt7xIGXyfzyyifM1Nvyy/HJwrgBfE0aeJlnPqvfdamPDGH/4Xe+dpl4Do7
5XwI1xJl4jVWUgrsXM+BwfKuaiEYLA9uNEcM18iGge1netnRxWGVheJXNbdk
3jGP/pOg6lxqKd0qvUjnHSijVkAXyDxYW7JqWvZk3YvtbzSCxxuqE1JTk1hp
oeZD+jr3TM7bjxD+g4vTsbXwLXAU2jMWYiWZLOLlYmg/m9qTB469EwKFVb17
OdjhVlUBVyBx691IHfcFBVu5Vz6rKh4CQBwmLTe/lN1fyCVJw/CzA3mQi2lA
aLdm99y70Cnv5SqSrCBOxegRZq3jlCGoORfarA7xMA9nwjhBNK5K2iyXEVoB
tmaWTip2B1/oS5tUFa7Xcfbg2hQYhtlI2Z55Th2e39m09B9QDjVuvZbjgT5t
wZBpkatA6aE5uRaSgzENhy7VpJNwG+IvMNEilUUIAXX7lcveZrE/2LgmOv49
SfygSELzl+J/o/FAUW4hyqRSFaNJEgXC3w60vBmdZYIfdCnleTCMMVEfwkEF
IoUHJk/y+2rXJJDWn7I2sQY4uIV+W6NjUR6GtLp45iF+N6rbWGz17km0AZ57
+sj2SxwfN34SWrqveAQj0s6X2VVyDMa44Lr+V5Na2/+DASEZVeQjpU/kMSpN
JGekCn5pCJdiblgD7h6e7kJh7N/AUFJ+SHRX52Q2wIaofIeNgqhNhfL9zdu5
KVf4/MRCkF+yRK1aNe1e2X+HYc2LHrONtaH1tmzA6xGM+JS0+pduHHpDvjh+
d0WpFYjqjWsA233aPYfjBJHhMosfQxEpnMwSwO1BVqUbYTqNeQ1jBc6eBD3V
QR6+bQXsEXEKz+OMV4fHrdexolNbTE35DUyYnXsvOTpFieAxnnSGy9ux+HXA
v54ZoHQw96mqriQjTKEl3WpIRbbNrNA+iCK1DYPTZKIN2bwfYBH5wxOsxETY
qIldauRgG9Mi5/1ZJjDYDSAoUCAhLylqm2BQle5TD0abScqWs1oHFHLG4YKN
FnArqxuFg+Wa7huNAuk0MR+Gixqui22l0oXKKe11oL3KJ+XCyQ3+yugFFMBR
PLGAaMPcVh+DsK1hULwm4c4rOC++m61zCEIreaZT+RVJkecbkce+h1O8HmR+
ZRmvnuNiiFZuuPTQJMa5MYuRZpteeRcyIH4IGUu1fSW+7jqv5cUHsKMlKqvY
amBgjy5cZKW1oy1zojO302qngdxwSD73X5pqiLFSFoYmzKNiMBxYVzCMuBUZ
igpvST+Yuv0w+tg2Y3jqSyaqAtb3uT2AGzw2mTjSrp6ivDRYHxWwzWK98+tv
sQS/IEoqTxI1qdStxBj+hgT0RGwWy9u/s38IEtP4SM79mKIyWY6LR+JPG2gD
FYmHlXJR5ymCVI2V8dxYRrUal0JsNZnzPKXT1Kv43vqZqMK8QpMIkqiUjvCc
Up7jtx8nmMlH4QhHaZ37IfPTKydaxSH8z6fQMGtrrlyPJKr4laBlBPYrMIVK
g3OHnmXqiQjznfGUK//MCJ7pyMWp570xaSBoitZvmTJqHFMyM2LvyJcAdLLR
4YiNeq6qjpq416gT9D3nQUuWwpCmSpb4FvxcgPTrcZfDO9yQ2eSX5WUniye2
Bo82POK0cIbMFtDL7oKqK2aqsRByUtdhne+2161rbMuEYZ4gv5lG51KVaXi2
oRWtVJdSk0Zv7oGOnCpVEZFVx/9GID2cEZladGM18p8v2MNO+5EZmCRbtB3H
XXS90JbOfThtrdqrVHybmecByzHOvKouoao/lhp+Y2cCZ420XdgxY7rncJ/n
N+TbfJaulVeLYjul+FZONr63+QC0BD94mtKyNJtayURkR95vrf8KSYVqWrER
/1ei5RiFTLfy7pBFd+DD0ui5ZtdTIwg6FqSF5U3c+8d5LDOKifwYiMghgSYe
oJrU41P7Ha8dXqlFTPQ8LizPuDS4ivk3Yuu+/bgbAjjIcJyXNvlSAhnGaiFp
z5fR1glZ1Zm8J8BSupyd7H/PgFRxEXdDgmhB+a4WvafGKh3cYcF2ZgPrVq6U
NNci80hgOlQI6l2PPWVPE3tPptpEr/imx5fb9+SMiFoMt5FF8c8XN8hle3k7
IIeWgdtLYNCMG65BsbhTS5bPdw++agKRkDkZ86I3+ay268a/8PU+G2i92tfV
DlWqhLOxXJiwMcCJA/ky28ruIjyVBepBOz7weBeTaPrC3JePzUbNuXSk1j2y
+aAS13pq7bsz+hJNPf/+WcUymTke///71m1RFH5G3JpT9SVWJ3jCgG/bH/+f
qIQna4vReWFbmmEbH/svH5tICoLYqPjSQDKVrbXPwgwLKGQs1ypQWDz56v0L
86D7ECcsC/R5gUWwrY0+LloqrsOuP3nfzbbkrCvsFlHNdIRFtpywXYIwZbQt
xkt5kxwK23OPnDkXvcatZdD0tbT+CZFpeV9dId5MRK/RLlWthsI7Ix8PRgmX
etCT/VbmqlfAG5bT1+FhQb3KzY+7cFZLlJ45H2jF4G2Hwar1W2fdvaGfQssr
Kcr3FiceMlFp9Erqzx+8qtCh1HtzLTmLwH22iyxGjYrVZUXsXJ8aBx4qSTSY
D8+rpsHELryn6VLq2Tqi+ZVSuPCZu7F7yQKH+aeB+ojqv/Ig83zQKxAA3Zl4
8wgje4O1oNLgVI8r8TVlnkXhBLh3nEnAmbwZwYIrcatOKDqdEaIm/viQclkl
I8uqbejt/IzAN979GMaVHGK38v6hxGXWjmaIhKRMX/KWbG0QjD1R7dXBCIUx
50ayZMv2uS6HWns68ELkWDshrSg0AQEiwI1/13F7aEGysIS3IfPmMzx9J0gQ
BZXnRead4cq/u/Jbzoixz9fj1STmWoAImTuhNqPWvbqSqv7X6caa/FNTm2xf
vQS9NVQgC6Jrit1/vB/6EnE1ZOW90jve/NcOACdNai6EDJqASF4iMmuICZsx
0e4TrisvCJm0TGBeztSexJ9fRnWbP8m/MAz6qiA5LkHmpWidVAK8zrhjQI44
EpXXwT8l2fGK0yWS2psKm0jQTmAHX1AjsGYzGsdz9qL0ZUEff21CBh9nAK5U
5EwKJ9gkPh8h8lQkDvRPAo7IXZutETbcSXBfS3bbSq5/1a0iRVNmqaykymsV
TjBbzcwxnw/EEDNkIvTg+IkWfbj9ntwobU1ScrZ5MVKJI9AyevEKWlGRjLwW
YZgZlwIGsWMwmNnUaUcd6oJ8QyWQVLMsm3RyivrvDjRSXu6q+j3l4cxAeh9c
BLeRvkDez6RHbzhUuMJZZcD8H6DfUFkvduIQDEn89AVIM+ITDi+0hb0dVjYx
3pZofamDYCR84ljw3uBiaOAQijgmvdYq3tXi0HHwCzFY3HUryAFif+tLeXSj
2AmRrNckxlCursxbY7mqwd3pl0s0syYOljatGklAXh/bShC7zrWklKqayItY
L6liYZeObAHFcYsBr8ocjBhx0c/ejOGYhV5NbazHRG0cfYQuQ6+bSIOA1zx6
9okqHc4TgEvcj4933Cddct8F5Kqeq/uKHX3E4Ch5j5zWneyUH/jtaIzfJhCY
RoB2+ffmaLlumVYikTbKLzMDxbvi4ZK2AdkuJjTr90dZJ9yc2R/W/A1dYozv
YgFIhTLpderp9LP2+/6mOsGxZBa2/YagV7Zn8kzS3hpXkKq6s5BkZIir49DA
dcSYBJsFloyZ8GzkbmiRGqFNgOGXrbUtrrxeyiENuOuU5bjuhj3cFYnIDa+4
TzGBSTt1W9pMemutpr+QWO8ddgr22iDxAXhV8d1D+Yun1LFelBIqh1QhFbU6
4utxNYKIrSisuBe79OtkIz9Vrh+++IWfLCdD2IH6ERBLE9wTfZhruYYFX1lo
CciepjTFten9bcojwoZC22yLJuDJ9DSsEumsKSa4E5eVc0WiSbcxhckNIjCS
/+Cmaq5Je+zTsUNdtI9d4feWQOY/BA6HO5VSl8swfxq1yo8PfZx+TbvjJPkQ
Qwwb3PjdqLy9dMzg2oTvn8iNqOCSWS/pdkHFge3xVsmo7/BBykwUPaVGVbo4
gXSWzBrNINWtP4ibojZRh6KpmwMF5pxIZ0/24vn1DW/5cU/Vt6pGiW+p2aHK
hAabqi914y1QUsWgXnMKSyoY0eYtx79iVO9AHZHvS7gfB448s8UOUj9MNUDd
GuRyC4NgrF5IwQKwk1ljTmuQibNVIABgxnZTuwFBlbZMHmhxgExG1TD0PC6L
tHfqRzM7WFoHG1FvObSHGSNC+T5x72XHBHvUGDL/rTku9ll/A/2Mhp2jNEgy
P3W5ySyJG3wqATUv/Xs4PeAwshT5qkV6+TiizMMyKwripoCh1H6Thck30A0N
I0yyq2AqSr4184jyAJ5UiwNsr0mTkfxm9k0pInOlSQeMRAgOPN/9aHbfCrjm
9Sj8/KT5xpMf2eq4bBPM93bNlzlj2inrONHpBVM87NsP4mq38zDGUW7U8NVd
Sx9eW7N0sDkJDScwBCuc4zoR/Y3MLJ8GPRx/9hoWKHs5t21yqk7hJfrHbcy9
satf4aa/zPH9ZGNWo7cCZnW2Pc8tF6KMLUlCy82chUjWiPAKTPCWnP5Fvqtw
YG3c1SBdIdGfCWvSt3NQYs9/nfi+PhW5x7e6bSehTxN6AqM200jsnZBUAlh1
qRCltAShv12i2XBO8R522CJxN4z7VBh1kUZdR/c1FmGFf6wkHZEG74M/s6Mp
LEc0tay7fwg6xsnicn43vaDVjh4Dkg1npJRR3jdgGvmyoUjcZ82M2YW2T4py
XdGwVLNaWJQew0kCkNFkwJTRgfATXzW0lJp8vN/XnRXxUX1/75OZsUyiAyUC
Vi170ovWn+HiiarTuLNG4AuMlVVsGbMrRZHHWV6DLS5D0PHKi4+tGD9Yr///
pL9DCObVhJpHVBNT/rrhurjV1tsublbPJalsdMaVM0qrWBXj7aOyBIJYpaaM
3IHf7BK8cWH6iOuAqwQcFNu6DiO4VTzZPIX4+yrSgUokmPYF+pTQV6QdBG4w
X6V+UrFhA17yf1CSknjoUCK4XIrtya9JRWvq2MkRpTlsQn67P1lleGpspUPv
A97G4NLodX8hO746EilOue7N0iFV0Dp2EfMmBnkvO1KAQCcItSyFvwJOb3hp
6osu4VV6FTTiK/TsxjeSp02EfrAS+NOCKBoSheTmPR+1NKCVyM9wf7ytYuCb
0e9OMorzuiOfv5CrGgzEh9vlbsIVsC8nqLOArBAMW693PLc+Rs8MuzhosZNI
ShnbhmkxlhZtzjydDYDGgK1INUNaM6ZurhXrCrCb8/d9Rliuk5BGJgT5mjzI
K01sHWYwRCTz+izQSkHB1WMKyiooYrzRYYv8aNTEg7sNM9r5dPQ0PuBYx6eF
qZHT5jsCmKQPZLcw+0zjHx1IQpRH7bG1yu83bloWch04NVa6mzMCJYeuDb2t
9/XZVFE+Vw0iyvcPW9Db71hit8Pubr5ns+7FfxobJ4+0fg8OrsGPnusdVPc8
Abj1dDPHfiC58MfeFIaNtqshHMtm3HcitUUt68eJ9/fBPVEvGw869wkX2wRM
u2j3aG87BDuINkryNgYcsudAcObxxnuX7gaco9qcocN4eHLAQaZQgK1B3eok
d4zLQDUFbvQPm5K++Jbyyaz8c+lkOs4VDyY24FtlqLdlaAxx74Ir/IUhvb9l
1MLZuhGVPjx8DpLxVRD1BINoOPX/tKqnV7tVAW8jvToZjdoqvSfUPKPMoIn2
ovqXRaqz7Z/Lkhe4dazH0jGq0b1G47IVDDFtdLnloaKKkPVDmfoZR2ch796r
Ap3A946KMzMrn8/Q6wvAukpv/7wSkoljOMtN28xAiw81mPwrWcBn2xD3qv/R
jHdDL3jd+z7O+ITGUtFuJyWmlPzSwaEtCysKHdwDnCvEo8kJCE/1GmHVjd6U
XncpX3DjlvhrP7jTUtVLIEpFsHRfv0oGAO/QkLXg7Vyook1saRnwxENP7Xlq
NciY6c/mD6El4U9QhBx6d+mTBdwPsGhWNFZDQkUB4zY47jykmzF/FoBF6Jrw
K3834NR9tWdwVhYhdUWw/oCURhP9ciRwrOv/37DMDa+INFtw3EqL7Phh/dIO
D594F/epDhS9uJO+ymbwwbyWv8bs4TsdvMOiCE6QlSiYDrrLQ6KSmVnPDeK3
TpPO+u1BAgfryBJvMEhsAndzvE/FLz3Fauj61Km7DHrm40Hipc4F6HyqFhx9
mUJSYVD+Mt5ncIMxfyOoEt/EF4CKmoigStHY/8TNCpn8VX3q96tqXX/bVC37
IGnKTTC8iE8evqvGZMUg332Tv6jmpuafJXPEvSwkFDdsYqQI5dqBU/+qAtWp
JivwlehlYsgxT46XgVcuN1kCKA1LS67Y8qhiNerEzSIINg44oGY1UVzXTKWo
m5goTvaqmBaHmF5qVd7T3SIO/O1BNNfpZotXttuU7urOqUQ/CjAydspn3R6M
u4o76Yj7lwU7MyXYktgwQdQuUYHZ7PhUqMxiM7pvFyZYoDr8XewnxA/HwMff
6Ay59ev5f+mvqa4MabiIiVSIspAW5F0mu0QnApfvcY6rmQZ4Jwjdq/PWhboZ
NDlc4oDb8iyKmoI727SAyhGbuXVQCUhcT+qlLCiBq9PNcH5t2IxiE5+j7yTs
jfmn/QIZhcV4OPRrymMVXa9wiFEFHQqfYI1pXp1PXU8qfGlxgINYg/5iLiAT
yNquz/ZZV5v8Dn5wDDodRxw+ggIMvD1As8yVdspbMADRKQ06+jmJvTXjWlxM
S6v7CyO4uZzAwsB5mhf1wrmQbjYJCotsDLEZUa7vD9iLKL/IZCyH1InJD9bV
XqIPSq2G8Jh15qZsA2TD/XZPim3ltATd6ve0NqWGFZSdUBQ2gRkDTe2aAtoP
3c/D75tATxSuns8OOymAwYX9ODG1RnhGUONE/CrH8hU5MIGn3atybJLckCYv
gRKyYf9enfsiiQDNUlzyU5y+cEQBGb3ZfaLgre8iYgr25x0DzUpGOa9DetbI
ufMQx6HSAMbp2zJypgRm1Sm33AUTVYNNBBYH/+wi05JD9kFuJh+Corf4yj+7
dKu6ARjOWMXMyI0VykOYZEacyEjEJa4z9lkj7WmjXduOg4LNq4Yxfs4GJ93z
ra6d0m9AHiOG7yPjMh2BsTmhUofI2hBssT8Yw7Qk/SVSwZ8wVkgn2y4CUFj1
bS/AlG1c6OmaBiLtE5M9D2e09G6mS3wnpdWIrf63SqJYBVhAqW3Z8hI8fV6E
HGTDAm9QK0RLqz84ggBDYZLh1gHY/pE2uylRCwLrEhLcmCr/59qpwvfNrIKv
SmQCm0+vWNOXa1B+cDOInF37PcYX/ouGiWVxZU/nfrLHKY4yxN5eNzl+RuV9
zPMbhj+G3JFU7ieQWnpGvqUOqRlQ8UhlGu/RSwijNSoI1Sphn5MRNLwKOL+A
WLilYk8J848ppGKf57nxRahfNnmp71puHgrzbEIFwvCKur8b1us5AI0uxP4N
IstPjQncIOaA4uZZAS+Pmo5DsUVbnAbNE27IlfRFRB6XKFg6lUDTMWLiNYcZ
omyMGSkVTqk+IAdqC5xqn3aEsEpEuRBGRygcJA6uEHTn33W/E12R4HqG0Amk
fvTfoQZstaLjTWNRcp1XfsJuuKeqmMUKm1X/veLCBT1OCfLqBvj6Kx3kJyPK
xKTa3A+nbXL5WfysJUbH1eTaJlRVcA7Zh7H5cwEzIXIa5Kd87rqsxZKSsEqk
+EjEBM4LF9PzvJRIawneCa896NkSd60deTi0mC/xydEYB9yP6wps+QZ2lnwB
X9an6FbcMsbWCA7umEj9uNN2z1PDeFJ2LWD5OBbXEFOvLZfwMxiQjuTD4x1/
KURuaF5+gLJcDTho1xm18buclUYklktwNjBOLeLX4Jgo8QyIENnvqBWA1gpR
fWnX7lMJHhCH+f1y82KbCvexzUPCKBhWLyC/wmH6ZWI+wt7yo3/BO2ni/rr9
I1md7baU+0rFKVNIe+VmT6eE2oJlEl4xbTSNyML3e7NJ3/RJGIlhh1xqxYXx
z3f8aPggTG7YwHPMXqguGglTOaKilbyvKR5BBp/02mdPko3Sk/6BhbbdPmQ4
EVHaVq1jkS31rDnwLCyIYYZ6LUU0eM3OxVz7EA8rPXDeSx35kAm59VX9SOhi
1Xp7z2C1PdfGmfS7H3O4LFjrBMoW3lloT94iUqK1PlkW6zeyK8XKtdThBdg+
T5BG9bYUIlxvSxvLXNsQhVq3H1gBmiaC4A4sW+758waOc9rikYA2PhB2Tqal
bh5PqW5ggF2gcwwjq9KzkK8FPaxoEr0/xh4fyVmdAf5GqPDV+MENEfy9mexR
0ZSGj3KcZV4xu42As7r33eRXXCZnmt7gro46u+a5OokpgK1MDJCILdvcenRm
1EJSqi9X8/IPX6Vqow+GaPokyQmg3cVs2+E3V03qgxWijnrpM0M0+FT3Yfkh
FTponWJAJVG9eaUx1xcxj++jjiG6Dxfq7MyxJgeUolb2lQ52loQWZ+i84ANC
b300a3kKxJ0Tu2T8B/LV37kFacX0161n+JPfyYWpoH+xflVXwC8BXpqnoWKp
4OjFqxYEOxS/sEoBeCn8Ixe4Mioj9WvizYY/EmdC9ND9NVmtns2wVOkM/20u
Glc6kusyfe5SOgkd5HIgPFQlDG9QAHi7hbvFedk02RoYv1xN7VV8r3ZuAM22
UjH7tib6hpzynjVlyPw2yrSOF3EjIVbwu++YY7TWFAbw1FcGT69SK8VC3EHs
q5Oi2luRHzT/InMdq9h2YvnOpPuJBnNt6IozR0wFOcJN2rxxA7hQpqIZQDsr
VSxAHESZ6GqlXBctB5lkvR0eGBWcGqand+ryDfpDt98BogcH1YluZQbIWcy7
G4J9fpoTtCJ768RvBIkrJC1ndjB0d8JOdjofC5PRigdxt78hXwoG7uDwo94k
m1n7L93Tf17fI+FTBbc12FQQoBHEqUVZ7rLVAx2uP/HT4LpnvZwK/2Gtg7pO
e/JvleFLiNfo9NzYXCJPYegDSw+DLjZzyGhzy1MJQsSfL7JVg0mYxuc7LNTx
YMZHy/Z63OowTxAEYnp9bDjz7t5DRGALp/0cUq3pMe7yHhds+/8TnvLnEpqG
E1e3okUawFLRFLr4s+5/Lunjumc8mWWvGBQp/Xr2YAfn3EQ9fVwkBvnXIDsr
zP+YLqTM5qyCVz96/mqMEOZqEARjUg1p3LkLJym1fAcV6R46SDnlu1JzvLFW
hK9ZjWQF1Fn9bu0fqCKrvrgKcQiHsvzPXXvK4YwOzYjkFgo2D7Yod7q/jkcL
P6MRQBsgoTrdYWrhZhOJdc2N8sK4zUtoLcsEyMMSzhbv646B5kvvmLX6CXth
upO3IXmA+oicyoPtjXOkis6DIBvPTZyNeHA2pUuv7UjhhpAxWKUUJcC6Jqwr
v2zCVh2d86zKaVJFB/9MgV6X0e5NLkg6nomXB8ce6bZdsiNN/H5GPWmUEod1
sU1affp1FHO8xt9Q7j8yeBUi7Ao+fiVu01cCXfQS+FA8X5aVqxzYMwK3nsFx
fb7+6p+ydi5dDQo8Z3U0nj1sJooBciUcIgVCGkDruzNY5VJqML0McsMp+OEj
U6jNyNrLPG7OzxjrFF49e/3x7lG3KzwC7hAcRED1BjTF87ZkJYhn7EqlQ0Ot
7+zX/SsOC29XYmeFk0YFjly3aVrSDmlfZ/M4lUeDKCCyrXibPXp8a2C77kqz
wgFs0OrSvDnYtveUJX01khrY45ZBaJGVpn34xua52f+/9T4V4b5BAWF8hE3W
kdnXv9GwN7Pd7aG94qIQXlYJJvrZuOY3YtlUwHTHJlXtAwd245rbuV5Ey2SI
O9K/cqTGSzAOEOco1fmzv0JwtZbPDyYxHCI4QZ9dNUDnIADsCM11g3uKppGd
wO+K6+NO4x11K061767QFnNYGbnhrGqP73IpyVMO6NR53StG7uksiCZ+38aG
0BcadnPY9xjJyobGsUIUeY2hT9AEZuFo/aMGMXTkMIFYYZGkfhnOfYvL/NQs
k4mbEtys0DSemQ0l/2Ok0OrMfw9qQxky5Au8QtbbzP7VDprkV3Gf0xB/REGX
kRJ1DgpfVD7ggDxRYYqB2GYrScrvm1OwkT+aidGjQ0yLXURL2IsPXOfYp505
t/fJT+Mv7zkz+NdfpdHyUVWBIX6+qY59fc98XKOM5KekRye8IhXuBH+Fvi2f
PV81IizdOch02ofYM1dLNu9zhag58OJefSBAbukCE4jypvJ9Sza2Y5gRB2gH
tsj/TZc6yhIGsiBVAIl/xSn+FSHOWVYTGW6yxi+TjvsAJTycBTz1cV54iujV
rrIuMsiCTHLVGKAq4bvicwzouirC+j9gAziZR0FvwkWQZlVyJH1aeXGFVoFT
wcAeeitaq/v/QV3A1QRYz5vtG43lCiXTzLfOfZlSIvmeeGHPXDXxPOw8MV7A
NZLE2NN1XXhsq0HE42rVHADRTuOPJKkbmgGsCT5nAW8IEIQf4z21tcE8zw0Y
lj6o+SQJxYhPPWko1tkka6AJnXWYRCUz8klHaupNsE1iUwqAIfKDcGNvB8s2
TlB0xIQ5Dy61Y/LAcp4pnfkwTqjUgiQ89wKThU72QkJl3RH75bds+4dZfEyG
7CKNqBZFqO5Z7G0n9ZyZJAGwRnqYkBTu2tf5B6bpVNoEiEDxdnpxDWuWyg1v
v0diEe2s5itA44hG0AWzHssYb1M5Ybg8a1siI5a1OtDIkj8iSeG6oMx+M0/Q
HRy335ityRopmCxKGEXJMVn6BfFrenZa0SZp8jwu7NGnfDx0/KrFuSeTogyt
R1qGRgDUW5Y1LPLe2q2UcLmfzLV+LD10kyEBcTR5u6a7tgwXnj/WZIZHgxCS
EOfTf5gWuWltGBIn0FosvUnDT/Ey6cfQTjpSlLfMtN0G///f6u8SXfyzjrsJ
BqGTcGDvbFjegoMBNZ3Aq0xNQNp1nvjQwyBdAEcxw78thUttRO/mtn8tdZaf
qbj0BE3LLX0KNJ4kvFqjoGj2qPcPx3OxYtUTcie06ZOSgW6xKiKmXvXUXELe
77JGVyInnGTwcTaFb3L2RSbTxmMAlcaYOaDzMpiTsLcUCiu7p95g2pX9H2jm
M6tcAMms4k+YZxOVhhA23B8sFIlKZ5fVNWgb8ehITdmelGUOZekdntllz+e+
sd9coIS6dcIuE8VOn8CGkUkBdoRNOD7LbvD9yNgZ9z2LNyzmLxPD8DNZtck2
oz47i+HZ4FT/TuX/zk/BLBliRR3meO4hemVsclokF0eC5BG1X8/YzucK1Aul
Kz/B7kavMIyA8CRQiLPqZsNjovCrFE8Ii1wWO5dJloWNwu44FXXF3EzNpExl
XMrsmo8NJx58ZDmNFEIiDsXh34mqCGlO+Nv/opURZKKO85Vvk+eaJgwqr4z4
NPjQrMHJdnDGahYsm0SkdMyURr02e0PuVBbIsAy1OCgVs62aogQxvOH+UAvI
jQGgaz89LLt4TPPE4yZZtx2BFQeGmdgbKmgK4GARTi0w2YjD+I2mUp5eXxAx
eby0V4NctNJI6RRqB2oNAQoUYnRWdbVCB8Mj4rmUCXw6Y77Qzabncoh39p93
JMQi7iBGmxpzUBp7jD5PRnQxc8aORvqWJAHZZEX61EfhkpFVCkQi3B1HKgkK
fAVe2i2AaVX0QJgvlAEGssvxlP80E49tgu12AfvGmbtSP9IE8nuZPEUIgitg
QF5gZcF60vB/v+ajlxGzclGN4/riSPKU7d0R9G7rakq6hwscZgru4UHzP/I/
s+FuWdJ2ESoUiz3ta3/dzxNVKYWtcABgIueqylqBQvOu4nvny4QI9payoMx/
QbAdu+PbhiEvMjseIDX6MZWU/tl9raFxOJZMLfGMLguxrVr2ra6rLYJ8rywG
ubDWSkWndeOQpqS1XbFwG3NO6khYqyb32IRE5XMxJuG3N4p9ERGrlalVk9j3
usZiKC74ZbRwMxUHQQhOePk4fR4Jq6zmHaJPU/nxWk/xehd/Xpo+JVPor4l6
poZ6oZlo9fjiPLqDfAHPrDh0MLIqIXifKMDxd1RtUhplJBZ3JcbfswjFxJWe
ksGeLOZeUNXMl0t0RIyFojcpBOX6t2y8KWy4DVNoqPKybwwMfVMyxY8cut74
CbCNRYLOHsDv4HuB+SmjRjQarGkO7RzcBaX1qKJXOGdw24uWWA3QWQwHB5gu
e9G+mkvBCbmOamRte1LLO4lgPN073P7o1pW/P3W5bx73dQENUWZzkEARbjDq
qJZHLRAUEPWyuRkNeB7MhlQqWzcsFOiCFEEsIoMrlgVwCXj/f+jQDZLsvzww
J3esr5duvU/9fUDiYpMZMJ7WJNLQgCbuBQkIuDWY+h0YOLJ/CyTJmFryfGQh
SHtoL7OSuOWRgvc8ZEPLTbCcJX9sQwa4LSw8QB2jtD1QiWAZWr2XsWx0RsZ4
SY/x8bIxf7F+cg3o2nxIxQ6xCkC7z7C7nUqq/GbDmNuZxqD1UPR2NavxSDjl
zbSFqcArs/r6h5nXbAsrvjAFHRS1OVXVga5G6tS1xWDHrgXKHmewVf4dVICG
y/dXvfJ/x3GPeDuq4Xr3BC/S00Ke4PuX6JJKufsVvJBsf7W/UHH/00JNyM0Y
EMji/ubp8MuusdIA+k3QhIqqhZR0RiWQrFMOIv2yfyJswDhfY5fdGl237lkQ
Jh1H2vJgKjXJl4ZTGRbcpEmFJOEedF8R4EsoRXyaOUJIwZHiT2/8aVwRjZSg
34mYUvCncG4+mE+tHNI7PnPnTqwzWJ1ZeGiIbA/KLbS9PT6aW6cU/kn3XZtB
mb8hOfPNjefcfCKlUm/JYTTWpUyDChkrDXRrVMMvwFgagVHG05oJP0IeE3nS
40MdOF/JrxSBoc7S9mUJHwSJEZtOuzg9+yXwccTx4RP0Sc8eTuD4KUXdvoij
2FkFewWg6gz0ofb4IBwXBxkCRIdtc0DbVBETB3imw43Y6aN8QeteY1g1TjJG
8yHhXttzKDRuD/M6LKFI5wfgIPqizYNXY5G8Iff4HS5GHHqC1WhJZHRxadP3
eLsyKQyIV0c2woVsqkBjSe81PoFYsxBlu277C/nWLQyVh7kqInW0b0Ku160J
90MsdPkBSbaahxHYgMwDW4anR9iq1e845ACJR1bvhw3ZD4TacXG+a5KrsqED
TfB68qCzMkY455udHOoXk+118UekY6CQXqo/PL6cCS9pCpVzSnV+tR+dsE6c
zp9wZEqoUmA5MTfADfBx8nrOEECYyFBx4CMC+WCIpUv6fj+t1wZovXvrj/ur
tabKttjJer6gqbiOlWmoOOTfQuqtyXtFgUvnG0XyNx0kFEWQ6IY9g6iBWM9H
ZKIDkLd6tZ1ZIGMESg9OW1GyrGIo5tHa3pINPBBtrmqdYyKSVixbn7AIvq+5
K5x6La4oStRikNFqleohvTD3k4wFJ6b2p3/i3UDXDtlKtbu5KzF/G2gtis5I
bZdobBq/CXgjd+VDAdSH1S8UrSi0HDI/zdJcAhc6hr9diEDUqWdnvh0Blakd
CmrLDu3jZUP0KI55nk6ipqf3ZJJKWHc79R9oc4hmmRRkzkDoGixnaD9e7LMW
DA7WKjNQOPZgx6JspBrhKM1m2NnT1z4Q1rb74ik8CoYQ05gYrT6RgXfOASIn
dt1V5FI2AG/NKim+j26fTjuIFD9RraJTpDAyK1PE+9dQsHvU7TRfPN8bNNn2
Xw9Zg9Og84bHp1bxyT2tws05GN/WowFQlSiG4nAarl5n4r8fFflFvU+0IyKC
OMSjNYkBfAnfAduev+zwtpKAmhJHux8mhp/pFxVWUK+vD8trgfQNsG38bRuY
yMYE88Hj49Gyld6McsBedAaHXsEFr3RRyKpw9kJ8zhW9Ij+vlCGdGzzuBswj
JX3XpaybwaV6MZg2uc68+b0UbDUPvOtSlwc0tonroh366P8nwSXrQiZ0LMKW
sZS3c3AWY3qTXf+whTTELFqOit4HeqBlXCe+KhGTnc13ue8Jt+KOliLFGaXx
OdEnnYpOjegctEGE7Nb9qd4T4gg7smm7tdZrl0Pw+D5y/8kTM3YPW3s0OUH5
zot5huF9zIpCuVxkWnI3ZxKHlhfu9tmB9cHBeBbXGiquQe34iD1oakh8u61+
IyKVdpVCqSgu3ZnPxpQMgP2I1tZWykSsJjIDbtNS/ZZgRyBx5Z25sanEDYjy
3IrT6hxRz0v7LHNpcpNtmzt4BKvphCawICqzjsbux2Q7p7v59aPX4Gu9p5Q3
WSkCQ1bRnMfU2VwVmph/9GJIPDRzztbb8jwBvdYOIPdIUTwCkv+P2YfDUVG9
CIvWrDjc61/gS48BCdfjURcOSBhkzRWnpucut+Vcuti0nM1+C1d9DgOL7ncO
mn0eUTe53/3zWGnci6S+B3jnROS+wOfTcTLJj1PjOJvgoQ1llHvXbxUCf0TH
1gzu+i6HdzWJtXEAC4TTNDeTkILST1vnQUVndXvbHJtHRpF+zlCJSkI0NGnP
mzvTcn6jbfYa6NWQN0CqrphMGg45u5vmRb2GRl8tRqAZcrf0huVeMXmZlwZY
mEcvTer2Gq63DebFJt8ws651KoaSw8QIvypiVRRrPwmnFSMgKXviMy4swD/z
o3g8MfrgBaAvPyLQbwS0DnHrDEFpyQNtrE98lj0XJlojWxxtZl1AFQVLlJRS
Lx3voUcamVLClcHtkeXK6nAoG1zsfQLnMjRlEE9DxSNAI5khG6G/72u0N8kr
IAumnrmVAEO1xDv89wvpE84UqH1bV8VCSfFY490tJfqw0148/0ztdu2+m4J2
oFQBnqz0L0g3+5OgXuuE75pygJIPBXo63jni7j4g0OBzh7blDMfsoT8yvUyY
cDJqBm+bfc3i8VoayOyCO7n7xYsb2uTQPKG28n+OPotvYpROOifMI+Gd2Ky4
yakn13XGOx/anervUxNuz9m1p5hx46RO6zTkE/k28IKpoD9QyDio2aFiNH4C
s3L5pfnYz79OslaCruXYqtjLLbcuOkOz+h5fDHharSuh7MsoCX6V5Mjclqx/
BQyar2jmv5Zr/eFHCoRw2dY8k3SbNhF21iIq+tIqexJNzcSUBFHA4tJRsD9e
UlD14E4wSEu+6Jhe7dAwgzuslrnxMKbAz95SRzUZE55X/+fylVs6RVOxnAq9
ZiKC/cz7Dn5mkRQL2xP0NBYgtnUZ5e4q9DxvOvJENvbH4P1Vp8xE7+DhEaRC
//fJsyLVXDNeo1NO//isKxboy3jbftErQO7DM623YDG/Wg1u0p6AZPCNoNnb
NUlJvoc+od50+fCtax4Au1YoehL4R5mffRhbeIZw1uSOM5q6jExb22aNO1Ep
LGfR/skVkcS7zfGm4WwCP2Yq6LMVpDlueTvGy2MaKNUa6JVXNQaYx07CNc/A
O0YTbe4YyTHLf4iodD/pwvSaoA1i9vJPtaI/+80bXiN7CHv8rQ9SIZg9owMT
JLHpHDY8ewhU61zaigXDRNcD05ICwJ4YvFDRWgsvhGyDWEnPQqKsXWqBQp06
whlCX/jHKGR6zojxCD9C9B07yQPfMTVyKXimPll8bv4KFKlX1KQVCqdbfVGI
7hVVmm02u6eA0DoIo9k1tM48K/mRVdCdblJgwqqD80BDkyp2gs/vQwlQfX8g
NXwcOugAX2ArMnIhQ0vtIwu7hz3jprvPO8v/8+oGVmLMqJVtVh+Ukllsd31G
uWbFnJ0lvLYw9WI60uOiMMdTJoTMUcWXNyB9nRsoFwaxUZufg58GRrILIrDf
BS0RV+/aUg0O3cdb0j1+2MvUdjVlq5dI+56oL8XnhbPQBledKBRHi9DWn5iL
PRX+Bsput5jcJ+0KpLDOea87P9RVp35OEXnA9cbMz65TSLRZ8VAo04dzw99E
D+XixNDcuBEvXSPPTeFPfmSD1qQXXDitcjgM3oWaRbFO1GWrO6ZNOFy/vU5F
4DIcM3EMeLVNkURiwUkA2iL3CBLPz6T+nU+hAobny1JGRll2CVgvTYrd40PX
lCTlSRFtGvu0ydXwSEgtLLagnwe9thfWvFlc3nucD2R7vQ9atNF9NYr1m9Bu
2ZcAeiffCCtKoX3tpH1Dm8PTGGGlIJwXERnfr+yO1eWbr2KjxGJ8Wjm031+h
WD8wmKkKk3Xa7mxA8KH8fHwDGPkmiDrfgGT9aajp8i5yz2BhcbwiJhT+X8lf
VQv77ogAtvoKycPc/VoqFWoOOiD/GoAZ9JSJ/zXt9x+ZWbrg58Vi8Eg4fqdL
gn8Ua2p/1SOweotA/nZHq7C+xM9s2MZPnQmMyjw1zqDfd95Sd7ND0Xm0uJbI
7o1gR+2mJ6tHMDJXXFlElPssQsY616YktJ9vY9AZqY/y/uPHjEme5nZr/DMi
riRp82JkEPGaUPlddg2NLQCGSDKtpamNeK+kpBzcVyYqj0aKKm2yQojKSWP8
ifcON3qgdeNpNSdpQc/TVKJV2qH5vnrQ4K9Qng/MNJSh0cMtmlwfYpabUEZs
5FZ3C3+LdEBQIvyyAlB/TjgVCYHbElQdfoIqjswz9Wc3+XcTJkE/WND7UivH
3QQzGaqEjCHzdcblQnqxMPC3jDdDItYi9Fux1pMzsnfAi+RhgCKIXeZACqLF
TjjCCWyPh8iZTlEWD0f/YJ3ueY5BxQ0JrBNdbc2i7pjYanXNrpjWhuzC9UT9
q/qHVApHEozKRxw+bEqlVPpgqb5gJZ95KGhmworUPvGEvKSg2c90ZuKhzn1Q
E1kX2LbbVaQSDazpJi7iMbiAOwNeL0c3eHnYoR+YbTbTMwAC1aMlAmmH7PKH
A3IsjQS0AhZ9yg+Msgyh235w7BHl6wkBO06/polBxCLnutor9Ux09t2MqADb
YzTCXnbaQOEbQeRqeeqFo7CWM2jBZEymHuQRejQ42Bk2R94ckkv9hU01Gv/8
ppL3cUjch94uit7QL5C6ZqzO4LVb55NhjvVxre9RnkKpdqmLnmDtuRLxQFmz
28YPBwuD6Et/s625wkivvSEocg3vArXZODePPhxqqrAdHenKGnxA2c3csLqp
Wm/JWdJ2Y0HteGipnEB6pZkrkXgiRPPjwbJEGrDFp+ejITnQ69m98bRG2fqf
pOkrc+JQ/WLpbpWvZOswSxMSjHxtl7KOZgVCjB+m4zg6HQ6J5Pf1/tUT0i97
afrF7MxPGTjGIDihymayy16/OrAuAj40dhaJgHbxutqgyOJ6gxx5yPrswH+H
6ujCk61ZDIAqwOAx34cC8u79yb1XCl1QFvramshpzoEMTz8GmEqKhQOEV0Oq
HIcSaQcT/29CVfp7zVtUpz/9k7Y0+589GQaOeKbY3kIOAWTYMYWA9AhOTgp3
uExNHEDWfmFH4n9hXsPzLXagHajsFtD8uoOnU4bJX4HKn7+c8AJmcgVMM16Y
P0BkagO4hKPdKWMEMvSzfJghdZyeZE9t7B2OlJvlAKvkTZipgjSjd+VALuj0
+vmnsaKfgRDIAlIpAWnFsXgs/nsOdXjlcTNpssHN/iFNKnv/vvy3eETTAHAI
h2+bLw0QhLWOW+6ibERvtelyCzRijcWlHpKXi1Buqbpnzrel0NfomEO+9zpU
uu0qSHQTBoyo21gQMQkQhDRCzlK8bPpaa8zMwhve04vycVZaQNlwAVcvYprK
WA+RPDAbPM3ZaSFT6HUilUYnGaw+5OLTcfgNR3ww+XxrGJkplBp2r5ioqVan
GKyE/Ke6oKXUqvBo4aZLpaYKHCKwkm2jj02Vi0gXhiij8FusTcJGZVhE0pcy
tsw0h8cvF4fvEV1ny+HYaVWeQKELIwWuyErOg8+5n4HWWCVXyIC/DxjB1XX1
75YQJe75+sXUvk6hiufFegy7DasMFm+p5XGBHPtMk7kxu+ECPPN5kxBRI6Tq
8loQc6quNV0Sb8GBjqgAvg7aKgIL/3OkqP4Kk7mK+IFCWH46HyO3B8L3de0Z
Xv9QRDxvqgbjgm7iB2fKysUyHnlDRi1rQK5oA3k9R+8JxHIfboVa0HepvWB3
FqButkjEBuXKN+u0PFotOhQA4lrRkU4VEKVmeG5I8+QBmYzm6XcBYpOlzf4b
h6+7/CI0CjYU814Me7GklvCxDGn72vIb7ob3F6ntDxB97A6j8HcjecJjaciz
m0YsnqHnG9dB5oF0Z2TMKXXLsjgcDjJURCJDVwp+x1gJHRrTUHA2FJADMRWf
+hb9cTqcJoD44Q6v/ALb8dSn2IPAYIDcvoZxNTx3muPc4xblaWm2EeAakE5C
CbfBoXKy0jQffR/7koOIf0aqfp/3GShdfGVpvf6Z3lgJrUQVniHV8xm4Htt0
+z4bChiXXPWYzg7EuB6Lta+C5DB9tzNxUjhhMhdnCXVdwuibCtI61PAeZ+0g
ek5nmgfENQCL88xNZXKu90y5b+/fNXNDtBt7Z615Ru4WIJibgbAYZftSV0UC
myQtGQUfHUbqyiuJea3q3uxTXXhQWY+IQsFCE3zrZwC/YomvOEinxobZTCuF
u21izp1DZl9Oq3ZOqOyjl+TYeD19U+1y96W5zoxZ7mZmCF+BkmsFcLv7zC8B
9gPJUM0hwh9SZfHoaQgP82AWLb5oZWgC+OAObG55cQiYaseFcNpgKvG5WfSE
tQpd7XfWRZmkZtJEUBLCjcPC7Ng2DBnw4ezT9SX0EfgiYqXmspNsRqvZjEQa
RZZg1PN4seBxMJtya4yH+jRisrr0LVyA5a4UnTaYN4oc2cUknJ/OVqs5Ah/F
s4ZW4Bfqi9T3AVtq6/vUaG8XGUnMb4ZF6fYh1/lOZr/YNl8u/ayiuV8+nuIS
7s7RU/Sbyr8jZXivhany//80lR0tqV/FSiK4tfCCu89+jm7OZUYob1Xlh2V2
atOpCoA8xXpzF2H/VVBd0XaesCsyNBhVULwdP1DWAtNz/AGJ0yLTN9knXX/Y
R0nBf9yZ5Rq+qu28/dxRFs8RIJoDRoOCr69MKks3vbFzQkRuF/IIP4mvdeFt
p6ZFwMMHDcidRbKhXgjSdRCexYUOjrWQOTE6KV7pxLhWfa5g7AK8tHWg70CO
uqP/qk7BvSh0Soe6+AQIIdGeVqBiTqlMcJRK2zsgwIgGk3UIsoq9ZkAoO6BS
dLt9y+q9PhBMe+bFCZnDu4i1vtQSczK6SUjHWDz1BrFj9pImkc9sWCP6tWvD
ABoGB3/3VgskxF5ARhgkNmCD2tif462eHiaBp7WycpgPiKX8toPgU/jUoZ4F
O14tpqwoj8E0pl0uqsrJSP66nwtYSUYnsV79cSB+TcsIkdpaRU5VFBM5830S
xXjZ/MQuR4l6TeJajWr2gXfUinjxkWjw7ksNK47LuABQGjlww3KMe085Ru0e
A7Vh+73ZBqDj/g+bJVRcP8gt6CVUNSVS1Qj2PLsvwJf51G4V1fBod33DQGj3
tLrV4EMB0+m49idd7vMMySsdUxxwGiCH4ctroRt6epAC1niw5ZVx0kPs1Qc9
xsd98tRVmxfAscL3t74rhlJ3fu/8+HpqPLHmaXcuvBMsR705nT7dfy8H4zVz
7EXZMwhKYBNLtO0sf4/7QguaD0FOmMWny6yXTk1dMPsLdHvFdEhKKqlBlXLx
Zdemy/AmZzn5aLDUiKPj1qWY8bIlERk/T42X7SiBsa4EVITko6HtXM4sLI/S
h8WLfmYA4TjO907Porp/dsTfwRGlnvNq9XbHx/rVUXphhqlbj7gfbaSq8o1V
xc2w4boh5H8CTr41Idjed+LiE7PDo+JGW/qDXCtq/fSFLpYdorvecA71tpxL
SI8I1FiF7FEU4BuDI1m18cnyJVdpM26IJ5Dznk442uXgxIqdP5DqK9BJ5PmP
aOjHA/eaBuft5iE/taG9RvjvJa5OjPWRBfs+cFOUaw27rsl8SBdR/pVudlEc
3uU60mzhKs3Q0+ak7bqhdUOIEB/Fnr00qplT0hsRWPmFGp+fci0AD8jHS42M
Mi/Fjrt3ZgaLVcCk7fui/VKWXDpqenNjer4kRXxc20+GqowxF/awA6iNADJm
yRFf/bhzhXh7NhNOcBk2jZVY797vI1H0b6+uxAhX6ZcCOW4lCuLQwIx2/nTH
jLs0qhAQmeAfT+2oQjf5lOEDFRkxEbovA2uKbIZmMgBk8l4bTqfvXNaZ0MnX
zvm9+wJ0ljl6fg71wrX0jyIo+240XsxexA+gSEcPOOdFuqiGNIQibMtV7vUu
PndT6h8Z5NIcx4GTzj5syskm+cIX/dOCAc/ypgk0BoFtbi+YL/uknpIGVw/d
KrWiT0kMLIjhU5CNxHo2czFkABVm43WVaqBfnDDv12DDQhLs7wsKdg8S8VzP
tnsB5uoskZ1IlfeLZ3FdlePJGjw6WeZBKchGjUxlErBKXN49KfDIZV8fy4Jo
0f5HtVjGPiC6+ENisaQ1aOWC//J8yDVjuyFOYUiHSCg/Cv5gRKh21O4UhUOM
/4cWNMta+kPg/S41Ogdf61QsoaQYBjBXCkgWyFZvVXt5FOakRvWY6up8bLxe
zURF1h9e9NT7YOqyqz1jtTWg++dtdON/v3JNvcPMsspLOQl0qOjEJoStP9S1
JAyIKQ4klbj6z51xj5wDqowmPaEKwYg+C/I4BfLG0hfD3kmUFNgcWBV8+Tgo
el+ZeVJt3YPPY3fgsXZ+UC6ucBlLbMq9iy/ZAIn7KxkfuyVeBEIS00i6LBvh
eseNOORvxFyh3jF26XIDLcXRCtRmrwitEoWXEI0QDau3AsL818KWePGqk+ig
d8YBaV3NiTNTkIGctNA89wOvI5LvlwziQNrjQu+U0mtg9CWNKzdoQNCsIT0e
1i/aQHVewnstV9rlS+rIuzGf4XOwD+3Nuo5v3GU9Rpbcz0BFtYEl7ilBlM3b
BZGj6EPEjyUz2ODyGju9asGmmEeuaneKXtjduvaNCavYXejBxk4jbdBoj7+B
zhii6V/wMvI7OD4H/KbI4Ajput7OQAHzUd/5gR9Se68dXMlj1w1jN7y8fjbY
o0neiHLOQ6rnVi9CwfQarYO8Bg8P1YuadprPrercA6MuWO6ETkVWcKK/qDm5
8PLCkR+3yFEmahqb12wi4ZS/rnjPFemtfLX3nCwHTdDNizThvOHBai2O7tqk
eynnwYH4NKJzNO3t3tWf4P1eMlvviiW0xRJ2lgOIAzkR0Q9U50zcrRhpnUyj
Qh3KYY3luM6bsy94jY/BhcweqJCr+IUbsm0XRhBmBUG1fzj8xcaEXfDL0L/h
WQHNJ5ZIDBODrlYt0zC0kz4xwyY0ooYeUxEaQKLrSr9q2r0laNcrS9m9Ra9+
CTY7s423cfMYuvM+21o0e+C5AiaEffpPstSln9xcd1qnb/dOsth7/K1do1AW
iYxnl6+eBE8/MiJzeptVEdEf+jgzA+mJBFwumoO0KGMIsrHQ7H+nCSKHZ8Dt
OGXYfdBnq9IGycd/GFCkwu0EMGd0SLjUDR1JyhjYae9rJ32m//yDDwuZafFq
GMh5PlMuES/hgrMV2reg3K7Wg+VO7bq3TczID78ZIr+9qW6o/Zbtm39j77li
BrU7CgxxqiUU0HQ2mjHT/TpZDjYafDpl0fNUEEplYeUYIceaz738Pg5ATKs9
2pW1Hh1Cn8vehoj+dNWgU2jj/aUSDExiMNJf64U+p8YcIjWXNSLGhdqgJWhf
+Y7YG1nH9cQVLEFrkDxJk0VW1LO0MYtNOw6ZkaWUeBMMMUX/ev8RIBseMmLF
I4l3YtecDupWB+HA/eT9wJJWBrKQYbOohTSr4Hn1p+bvczKgaqUtI/5w0ldJ
EYl8hi2jaDmesp9Mmi1gr0/jPlk7dit94G8OJUe4tuLJpiywnfb5DPoMbNMY
CPERz6mE4A7n5kMjEqqf5Thcte63JXBvmF9triozn0o5u5jm+JjcT3amV64b
6oi37mycrCD7JL6c911mC1qHawP2w0rTROSx1BE/sjldnbSdcvuEu0CmBRy5
zEXpjFEeJ9mX6PfU6O78FpYYcndQkiSLeu5v+V5blSuA+9jwMVFHiDPlm4S1
Zz1qr/JPqf1xF4P3TBQbzyyNkSQo5wULOeLR0Jmcp+u+CF3iKR70HqoRBuPB
am4arCftcYaunDqoDmHzyyZkRx9xuHK1uTswWzUtPnIlWk4pxutrhv1le/Sw
KZ+MV+sbx+M4Fea8+cN/FNAuqDuA6bycw4VQRRJatn4qFgoVkWJ9B07CbPfX
fJLYe3BLXyCEZ8leWjOIB+WC83TQiDSQQWPXzlEjUhFIrjBgysjcza1j2Wbw
Bg+ncwV93kIdgS5stMAHYQh+HcRLMe7hMYocPxyUTqa2JgSrsIHm3mnd6G28
wr7OplyPdYVKNCVj3IEiB8yKudw7tKVhKR2Mm1tCnTmva0+28UttdfqTk9r5
glp60rSbcmybStdXy26TPlydU+jQwhJc1UWXZW/rYAOg2dEQjXKw0IwmU/6N
jVv2icZR8JWxIqn0ruJ9iYbC3tiEaFjwNr1VNeVDRO/ou8ubRuHg7sXHBzX/
R00g2Kw4lecHOcFANffXW4/xIoDpiWy7bgr6sfRMIgV/lGRqzio2NwxydB8o
6yRfwpLUzrfpoO+zexkLwfJlFqc4RrDifPRT6qiSdlvU0qQavrk7yRxTeT8t
GO4sbRi8EvrI8H6L7P0m2/bT5HY9/VUpqKYqaXsoxQC9kLgcYLvNuMHeIOaj
4KNWc0YHBvTG+YGiT5Kd0N/Bi+Mkmduj6iC6ZUSfQYs8+7iAuHhIW0/18QDe
Dsdqyo+E/72G86vdSvGoTCF5iRAGHbNUFzO3GRloQu4Epb5DWH8oa67khWCd
u3+OJatO4zK7SDlmj2p/Kp8hQ2mCHV22Dye/KJ9yUiATLvWZ2v+JDsWa6yXJ
ezrW0PvUkMHz9BklLH9074HJ6h+qj6h+2Nlij37+wYZUYBVWRCt2PAOAx1ZS
nmy+QaDuIUc7Rxrirm9LRS25qAmnjTaecenm9J8fKUDS5TSTaCVDaJ3v8tQF
TCOg3gz7FYpduYDu7WC5Q5+bgqfxxYcrHXKZmB5mVvb8oA52qCe8cwd3sgfD
qN+9T4g63ebfExo98/8Oj+PWv9uq/9foZQP5Eh076FkEuiGAAWSQfO/IRFbt
U/cjbxXEiRUeLgt9SBJZSqD2HZ10B6j8yA5NdmgqOynyNvx0lio+6Z1YAmzF
C2yMtFru/K/4pFeUqfEQyiYfHJfrg65cO2URlQ4PBrg1YvFZ1F+CpvIFw49F
EXS8Z6pvwmQjn0+rjoDFtleJDrAZQ+5b7Zq3ecVmFpsCV1Abc+mmbVzB/Bjj
jwCJSEzEsA2iFe8PAQ7IBh29qzDtI+0W4nwg7e/tAjNhpy+CsZ081u07gFWM
B0y7dBMRgFnNbk7X00g1A5V37mrtVNHchnRbojPGL9J0jGvmLhUdmz7s3Dzz
jgyPaleN1jaNUsAhk/lFJlzGbg+swEsgyoTRm4c/6TepdgAnZZIbFNkl4fMZ
vKGLqbRmRitnHqo0JFknSxApJrUHL8Wf38MHgR86XUngpo5g7zRgO9yAwln7
/VAUYDJUsKsIGbrt0v2vaYSX88yH0Ihrbmqiy/piFf3S1YEePsIKtus8ik0q
v5CmlFONUfQTwFJDOAuVtG2sdB52TbeuHXiqKwYSb9uO/OX7LB1vufm5IC22
Qd5hc83EuhKy9oCMZgAnlu84g8Den7nDPEIVrUfw4Qkxqq283r8/rvKfwmMd
tdFyyW93N2rA2olWZxr5tnaZc6YQF/LtKRy0wwhLXfvAl8Z6Q67FJUfpLXJH
orjAoEVg/A8wfv2jI0Ee58jjYtQ6tEDGl1/vLWOIt1nybmxIHjPVntbbJ21R
pEvvWF9q0YQbM0z+8WOIyh8Fu97PJqAN82WjzSihekd5QCHK67kiVjNesDJ9
sPdha9p6aMD0sYNJbGTry3LoM3TWR2N6paUBbLIghR+fybQqKL0pzvhtTmiR
G2qtCLrBtSQCXoxsRp8yO0RBuksZO9tGDxvO9TVUXLN3ek9oV+NpjzC6s1ok
OHY5tfCduH1O9qX0jRMs0j8zyvMkQyuqpeD9NWiCPMEV4nD1jQZFdOliuAvb
ZJE2Y+LUuODEG73YVpOLWZ2BuGTPBNjmluHfVJie22JtvvRh9ZZGZsRAY4y4
b/bt2n+excNcxjAaCp0jaU1yllVm1T0XT6VtNxiR5XckO+pkonGYx+0jVulr
KSo/lGEqMBkupclliwJCV9EZXFSLRbFXUbFH6tZCJk8Vt4vTJt45bx4i++B/
2WYHtqGvNldYhECQO498sm789x91shD3pjOd5U8mjEO08GC/AJ2C9pjpKwgt
ETgGxboPrfOgS1Qb5FJgIkT5c4a3FfK+i+tm6qOwu1Hzo5D2GkqVl9+9UQ3E
zzQ7TuG0EcNzUoudpAw9gDNA6FZDpYJa2D0pQRmz46z6nwf2T+jFKPWhAm5v
k/kklUF2aSLyuq68PuFiaLNPZ2My25JdNhQ2xQs/rpphbJRjjNiUOqqeb77t
NOi4krMyIV6UdI9Z2Lnj5kFg6Lz7J1F0IjbWBAYgo1drRgHVdDl47y9up5SW
FOJ4Ufp6LWIFGBw74LbGAiEcvFmoz84HofLseRHDKZmANAvZCgipuEqbAzrr
6ea5iIE9fRCu8tEWm5TWCRM49Ukn6IB//WVMaF5pBdhIXork+LJPNia4rVrY
HHfDCOUtb9MNzb/MJ7BEVnC9a4HY37tS7vdm1RZQL2XCb9bxGPYzp/qUKu/X
QqpdPbLNsPe7Nk0KX3if84UG/rfajn+0CN7dUNvELS1Uyx5uw3YpBnX7graw
jifuJPST1WUtAIiSTy3jgHKu8fa1wXrhT1dHEx17bd/yGkZI/FdZFJ0ebs3I
CY3vPocMEu0QRLNYqJGEFZMiXJ2XaQ6pnPucYjMrvSjYJbpupot/tljl912+
qkDkpN8KS3aSe2oIAuSsHWAdqEjvc7L+P+2I7b2924j7hjyqRuMwvB4UHD1/
BsBIoiVEHOlqO9PoOHvldiGFxeCxTDCnpa12VjX5kHnqpUhE5GoL4s6UUcIM
kDDyozzFwJVLcrE6/+mVcKK6wCaH9ofP0MTq0kd+xcZUfuBwOqX3VbGMB12B
9/n77Pv08pyK/AXuIAPak/837NjUclm/70/5Q5jdRh09Wyr54apaFSJM4i0a
o6N00HXtjkYnLfCdPzpNaqJ73987XbDZLbxPzKtBVZT4qQ2Iz34oyULSuTub
T007QMjvuwBr/cPm6YIAQMJr4JGlh+8i4G2ey83qN9DpbNpk7a+AsAGOr7y3
/IIPP6isianYsrboL/MecoDa35bceYLqB6UQ47oJqObGcUqs9ZWi7NcEKI79
ZY2QebLn4z8KJLlBP1qLJIJI+QrgU5eN6rIRunZbdw7bZ0IEbkZqyJPl9+Zl
rB152EXCif7u90JanKEp3gDqAcRv65ELU410twE26hVkSqsyt075lIQsYywC
oahjiSoTD0PxNcvCKpeoSyd+2Uu6viKzaGFdoyc96ZmxQM3HZlXMzMWxAbmj
k53CrnXwnlpjTKnzWs5Pe/YTEBDGcxg1iS6fGPDYzx5oVORC8Zt9g3VFueJO
iA1WGRZ+Y+uX742q2D816gCIp2hSBj42GzpV+YBF+L8XHPdCvbmp4BnYZqxC
e79YVh/JXERJMjUl4N14IeQJjxYLgwhzE0cto5Z/So92TQHnydljNNV/8yXW
+d1DoTzIRlG7GwJYD0BenBmUWKaJo0FdzSrnDvnkuX6QEOMKTeDpIhrjvkhs
L44hHb8NpnfevlZlSOgoWw/3C6TumAEKIULecVH0oky21Mus6yUsYGkN+dUy
Fqhkafiy7O/KvwuqEnESkhsbJf/DlmzKVmbzUknIWlTYtm2lZZXRTID3qrTp
XFpf3qK07xxX8d8wy4a1zfOKeKXwXaWGiTXIY7sfzvPTuN1RIDDkN8NoDDcm
uLW4JT0ZuhytrqMUDT8zOIUu/Z88/aQM2RRcVaBUVcDth2otGPhhBvUiBvlm
hZmpy7ZUHPhi53tRAq4JjWVmQYI8oeH4UYEVx9pJiD+DBbMsFVmFC5zq8yJC
0vZmE8mvWQ5rg7MFbasSvohcRUYNabfBr9e9pE6FyQWJHVl69JZGuW2H5g+A
KdgsM9Yjjm0+E2f3gWwSYkqMU6lTQ3XEPbo7M+YWfKSRvZ67Kf/usvhOBApb
zaQkJSbit1+LuGX7slWkaEKA8n8zKYqNOSvsKhmGEgA289uKCMiGBW2slH5p
60bfUL0ekRtkC8ybI7BZtmKkNNl98vecebCQo63I9veOQXPnoPe1+hdFDOxb
FPSC6wuSMrC8n6dYJV5lYF0dWz4z9gJaz2xpzkeGUFOTdMGbzHO20mtNty6q
CKUB//qcgXbGflYe24TxrCqyJGIVqBiYvTJ9ZeVBkvmbDgXOsCAzX+ui4BN6
qsrXDDyitUuhHncL2cEwmbgdZTNP12lN7t73CU3z9NH3j1fTQuVVIIQqyKi/
w45qgrrgzgw1+5a+AuSFCCyVTeimbcuJ2xy0I5TY7ackZiTAcNEZnIyDkoG5
Yta6XLeXqEMyHRb6pNUEWkqCJ/XYGuqDybVvAZe19ZC7CwRdZ5fMmKUAnqI0
sWfA3kvGH+YNHkZ9Tyy5xpSCLJbx++MJ9C5J44lzUEnN6x4mEUjobuIAa1j5
PgvmwSNHaL30QUxEz7puU8u8F7dp/mGl6cbvccXLXm/qYj7ncGmtdyzBiZiC
uTOOgPCu6IM6P3xWg1tKffLhXfnlkYytvU4oINutgfvhMFF4zKeUi24ynT7W
zqRU6hdVBjTpJVlmDpWL+hcethLNoIHyllqBnYxD+u+tHtpFxm2jfWaLH7B6
1fESk3Uesqlwlqe9yjikzCZREbkDR95H1yhTwQWSPNKGbJuKKZh+tYdRRHj3
aSXuUUyRH8Rc99ZEL0uITuwVHx5jolYXvGasznq2r9PJ5ggol6JrNBDvAhCU
cDMiwd9zQmI/eAE83RFssWdJSK2YMaQqz6WuGaGMwgmKCnOtSxw7RzU6G5Mq
0u6aqPoAmDtRN3vZsGA2Rudp0b3MgOFx3WjarmflcoXfnN6v3HIciL5+JVxr
60BiL4RVjGoo6wG4enqUSXb7/fY28QR7OzBpDCM+RyPoL3Zxu405hqPwluYY
JZ5M8MlXd7JHXwS/xfqw2AkSqMqdEKwxgTT9XZTU/mp4b+vPzmq45rTImoDa
BmXMqGuH2mA9KdZXKXIYfVEYOVwitGDd1e94HNKlHh/UIMka5X9pG6AC9T+9
ym/4U9ny5pMQ8+rQHmWAzwGN1M9pyD6fZNOE5l1DzYiYFK1m0gfZ2tdjF8d3
wejplIHARHwrEwwZLPDrQAzsbTWhU9De+ffqrEXMr8bKdhiljeqbnXmjtX8o
j4S/xnK9Qg0XCrEmU1FuW4vrDRcUEzSp4pfa7SJhwIB5op4bjeoyRq14oAiW
s+q6CyVpFBMVI3pQXbcTbEHO8zj+5hKqXwxE/IbzgaDKZLb1XjyRUFdak9n9
KBOYhOWangxJusbpgzm1ZdA+Wj8PGVHFESTtcFBlNrSomv7Wmj9ZS77IuU08
Ld906/N1QUOFRUfiMnMvZTowNgxSXuwLFaf3waBJFBY2yZXdGZuGceqRNOdE
13osMiPcEEQp8ZtvWv1elk5c8issYqs5vVRcqMQckYEfDuLTcnMSNSCWWqMF
XIfF9ILLAuqIuEd0UnKbm3e3xyD7SpSj5QjAsRMxQ1drwBYVYSEsiN5+f8bj
JXBvqppzuDW2QC1oCc5LA2FlGq+2WA+GIhMqHrmiXNL6gfiNUrcdLuDH55Kj
K1lTuahjfSyGqDAA7uVKuckMRaNaObbeP2B9OYhsKx5vD9SruO4ozKRYgBz9
Q7Xqp3L0aoiPZDzZvXEz8E3fVN4M3Ccd4xUKCT5io/a/5EAWraY8LHGdX02H
WylGPjGmBwfuWXvLB/yTeEEfWYVtEQBu9ex5+bJ9Nts3oq6KhZlatqI0dQ/U
AtdRyJ/HiD+7P2BqXF2KTrwpDWMN4ZYn/C1LfzIgA1o4ZHwNsofEH3n1Mwd4
glXRh1hs9W50GJZwbfT0IEYnAV/45c+1Lud4ZMQfcyVLaW2jx0bdrsaACqHr
DDjGs8JKzGS5jV28n9NgTv282TC5D8WjYUSgwmUBUFr68UPFVGjyTEBWqGAW
ufyvt9r8pwbHtkrcfTYHAeMOolLluJkMJZ7xgkJLJSjNfcTDvES7xbxIO3TH
/YV8YWL5L5dQ6seDfEu80KgppuxSWXbKw3AGBRHnVGJ1mRBjFGsFun9Q5WsJ
50x5nb3XDYmXW94V5IHrzvBbCwizcPzUzPC2T5ytWGhub3dbHpZwrWjib2j5
4p88M+X1z9X+ft5NPohmvUIe6W0ADQRxfJ49IqqOV3IA7hbkMf/kuTP7MdH1
EzXcV6oIZxzlMad1vfeUGdf1NsSq37X8JLOFUdzpCZSU0Ci2Ha1XBCl1UQH7
O4rw0jJAk6Ps81TDItI6zb7lclkmH1oLBJmdmRgMw4yC5drr1lsz9beuxDTF
cdIvNOpRHj04wuSm1xpa0PlxnC0f96DpR/mQvJwg4OAB9wWtKpqFa0p7EQzm
DDYyxSQ+o6GWqS1TlFfaFj3HTc5kcyusET/znn9+asBQd0h6fwc5bYkUsw6Y
iFBI0zZSaPZyXfFVvoHi5mB3WGkNqN2DfqUjZtiHD8a20vTTcPoRBiZZAUWI
gzRKRlKM5rTxyrnJ0aflFbwpyd0vu8F8KRjQx7bijqGfIp+1cIHbJ+oOUVML
0FTYLWT4oTuowA5DzTYUsgKOJbf73vVVsfj04WlG1slob0w03D4Hr06h4ISZ
s8zW8qstDJLavwwE7JrXmUg+PrDRZirL6Fiw0bJSzgXrZDgqwtx6h5k7o1h8
yNk4Dv6O4qZVi2u9n0VJVxHmSRlkQ2w7e+suWEnGW4op8gcyQOjNrJ0AniT6
Xkr2op5zaHqT2Kqelko/o+pjBkp3/G8NES/PmHV3p8dBVDzBxPRR0m4byOta
QOJehWKg1nif5Wnessx5Oed2ZiiFVezhLMgmwizvGCfENdy8NWm/Rw4jgmSC
CGAPGVHi4xhwDpmkD0foIjWVkXcm/D8roJLZKf11uzM9Sis3PKGAQXIesXOd
ufcLNqtM5IiGfvmMHuSFLGN4Es459vYWdTDDeJhcFqib6hIEyVn7qkR8+S8J
63Drko1unkrD4dbvzRerXjbd1PWSuBP1F/a3jVNnLmVNvSupafLSkJTpfiH2
0Cqpc2qxrx7iFmJnc8MJaer1rCbMDPOsC2rg695sPAEmJ7ZnLy4l4clir2Q6
CkbS7splGHq5RZ3Vk482P8sKbQfr7eDTBcMPenJ+K0E4X5xlntE8gRiy4RUz
ESSJhjmr5uQOeDsBZ+jcpKNf12O0SEv2Vmh80aPjUQWPAU5K7XcsOUe2xD1k
d7eSGIqP2iw/fQ9ZRtHykO1htnhY/K5GPW36hYgW6OK/D9sbZMfyuaL1weG1
6AS+HNyjatbEdS3V/jZBhBEj8gzOdOfFfch58bqAszGxsF92GTRNxB4GgV5w
yPoB2DUaGNWng8I1Ucp1V7KezZZ7yjbiW6Ma6SKN/fBRIg7UPtF2yekuvHdF
QRQRKfBTRdhdf01bmG5xlD3KKjLrlRWi3s8xq/DDQs8dLTIdrRRNpAr6Xg4v
RJ+NqwVvtbYUk/TyWuzYQ7NtVJg65jGEDEw0WuBh9Gyz3vw7dJFkqEk8HMVM
BEQ161oKRQFlAWd4T1b5kKim4e88F5nLPfDW5qqn2q2NfYn+F/qGwQObLgaV
uFlMuuul88VzMGG9rSCVpLM53cd+H3c01at+Hwa/XA+JAd5RPeIvOTIzDBJY
Xaie5iGo31K7F8RNv76da5+cyoLR9e24dJKRsNczf0UK783BUwIH/fpiinWT
3uWRbs2DBrtMiky9aoUKBvgxeUXhuPIgyACoc+t5dY6AUoE4/rR0qkxnBbKb
f4v5ej5wa4M1Lu6R44q4vy9rqbVtN7yb9ni97XdqXFVwG3yHN9nfwUsyEqIK
xw4QfLGX9FsHNxy7S74IkoLzSuzYuwkkoqummFCvGH92KgO1wYTJLK3l4u6n
X/ru81o6z/n5ohYQlJfmXRgd/oyYTRT+Y8Nge5tAVTDKd0QQ5ebfDPeVmidL
/C59eVZKU8QdYgGffapIKdTC/F+R4z1qg7wdTev0AqdounhyXO7O4Ru/gwF6
24BKSP/zwXybUM8Em/NX/MXQIBNYwkHdtr5Lm5wuN7+7aCniTkPAk536HB0n
dAvf1QGX5kH0BQJAwMCAw9LjyvT1hvh/CDq43I+iBENOLgQnYuN0xG/OJ8Bv
Y3O372tACx7n6+QfqvKJfH2zkAsQnhmj714LunFlCJpFi1Vxf0geULLEyzeq
DtSqu+yTBLNYzQy7dCkkYUVxZPyy5SpBu7EaYMano30Dv1Q7MYIjjLCYtBfo
BidE9yfYXgLfwaZB87xBapQmcUhDBpWCfA0amPHK0tvUsufjcV2aUDN0g1hP
0aV6houG1RZQOnK8NoEyPwIGR+Q5UBht2nuyNNbJNmwoU850vv5pyNnll8IN
/fSCnfVIAEq2jfIRJFfm4J4Z6f564wAh9GT3Vnp3szfcsYzmFvc86/tobf20
p+Oi6s9jeu99yoGh3CQqAKk5cmKHqizlqU6qoMa5vAdfeBWalYdFBSxsxCVU
tR/hkqPHmKunAfHZVwgL5QP3q5VPrRu2pJMwCLyLzTFRzA4wjhARK0BpRrsW
xwvlcrt1/GmL2qcHQWhXu3JjEQJgVzkMDI5Oq6PPlHDn4ZhVOI5tKU2XzA9K
UNjM5VfV4Ca2ldYUnilcjRzweF+caTQIzBMY20UqQtCY23hUN9RNyVwRTkeR
ZxFpOnnjvcrZZIGh8mdF+hwNaxopBCfj78WmhGsBkLcjMR7Y1Vsoca5mKvtl
61I9JcDShgUGOBRvjYZgEzu4jAv+Zv1fAL/ZA/e8QHvOM0vCYXR5h6p0b/K8
EuT3FAq5XoCpmEbjjhpgH2t/kvf+rAeyqqBrBtx6pMvtemO2LFvY7H36kaul
jCiZ7TxF7iP4xs4sGrOTtd+C2E3Yiu2COtlL2xaOXph7d73rWmtkDqx987le
4J9JQIMacIruHxfjlqeH2xzb07iga8AI8vUplxr+Dyv3EuTwnFUaLdkI6Sxv
Cq2j6PssKIKS1F3xTOwjPoCA4lwyyyAGLdfAKNsh+X0+Ky4SsUi1feUX4gk2
OsJhbPfBeIgPRq3k8mw6TstY6AgPZC+4X/uP7DrWMeuONebH8nSxlN5QpGQV
bRRrq6FxGCF5CWogD+4mYjJz20Zwt1ydRt3HMWYXyuxRxMOQimbGnxMYnXcZ
LbkPLA+peQns9BaJ4YZVTLKlsnouQWF9K3a3x4TwxT9Js/3Y+4XxbMJCuB1b
tPF8gg/KDaCtq6sYg/bO5hESRtStlVk3uHANNGkloieTymEzyJKDoiAOvZTX
7R9zvIQy+PH/rB/PsoxbbEFpUYLHFHoHIM3dtxGxGIcnXdOIys+qgetZwMHz
NfYDho5BwaBomQT5jIo7/7MWyBrp3moQ7Mqoo9IgcmWDX6GOJ5i9Krjb48qR
E/B0/1LxtuNsZKD+afCatvRXOeieMFy1oge2et/zLZB9sf/TtIJMdzK00slb
tAVh1BOioVEPvovyd/l+P8v8/COC6KjfP138oibVTPy8pxCuFKCQ2hkif8Vk
umMEiEym5EHuc53Na+MV18rdb1JI+2NM7B9L6eA736TzEf7pfHCC5msoauwc
3FpW/oBhfjIVRuEHG8UPqZwKPeEAcPe5HPB/AamiO0FjrXMWTdx6GyGmbvjH
9Oluo6n0fHlXFJPsyj2xWloEjwRQL30UufnuVaz976Gkzsf9Eeo86WibHpi6
udu56OBikeexevCBZLat47GMGJE/MSXrHto8imE2z2tXbs53xXsJsFuLle7g
ebbbHUfCMCXOnP3HlifrXLS1pFFI67iCsOZzMjmlzelJo1ZhmLlwcZUA8PVC
tYSuWl6S4049AgvyCAS2Jp10H8kOAbpkxOq7rXJh/B+L15K9ugFvR34Y2W1+
C+VsBefCOf3lFqTA3VbIIX5GW2J0bRScbvWcXTTnAZFAzoNVRCbA2zGo6CgE
164tYxq8DsFVmqZSd81IzONY+nlpMduSm4VlO7gIBe/zp6G2smWZf0TXn6nJ
V7SwH7RbcVVmSoRJ5CCzOMa/P/VmAi54bdgd3DXD20CgbPzqrN/STKR6M/EZ
6O1nb012/Z27zRgFd5DQYZnWIY+ekoXzkx8nsU0N1DTRT1xwmWOpHzxSfAt3
CO5qWH1ta2JIPZLeZmmWhjAnzvRkuw6JROhoHhfB9rNjLUH19YXUqh6mdzba
x3r8NMx3aApe9IBTNnVf29ZdNe16cnx/2xb7CkzpISfdmeWFE7Stm2KglwAw
h46AwRe22w5VU0ERR5y1flkdK8w+7pecX8rp6K+M0gBqrM+pm5+bNu2T1/4Q
SWductHBYYwGlK7UbElZgYwVgc0EawmTtm0J70KFOlT3GrzVtOaM3tHLSYZJ
d/dkjLp0IkBV5SCjuwLAIPAdriKu0+kWqUg3zVYXiGvbVPvVcDxhUXRlhB1v
BjJiTmKpqYjpU17YJ8OXRaFlzUYWIZXZ4hAnpqeandAAgZ5C3kDaKrRGc1dM
UQn6SpUm/zvY5Fua0g7IMWLc6C3i3dZJnQ5QW1s8cjqEdQkJUtdGlzC7bnhh
1VxKed/Hs/KVHU8pjwDS4ORS7jslivJ2brQj2yQk1namYsx12D25qeW87IpQ
h4WSrPBj6cO7THyJWZYzJMjaGAFwSbe8NOGZw0i5hs6ZaFefKd1eyjsJ6/LX
J1u6CWAiNSnAZFw2fs9d9jWZIjNEBHuxzNiJQ/xLIsw0sJZvPjbyPmNnsbB0
EfxaYN69vAlTK50RdUqW7p3wWi7wnhqXMbGG2qsnvFLPJeI5+KvxVQ78mML9
COAh46OwOwm/YUBqDa1R/uUc4dBDPg1cNp+bSUiwsNTfyUO4rs+ulTvA0FWn
hdOwyNEFRwPUJ1or4irTHU0M5I85Px8r458UJAL9Ni0o5Ev80n74tVgO7ljF
kdPvedHX31Z0ScgkYZC+4eRxnSYo2v7x6OCGekoogXjOp84pi11923uTWqCQ
uaKejYp2Zu/qMs6Fr/S9Gr00XE/K5TNIsr6zVzU0G39lhcFb34zDObVAeZO9
PHFUlnrvo1sr3bKVr50aQhoPYkX+p0LgSGpky1uCaDc4SIUXk2+E2Q7pEN5B
719bQqbZyC2epa7eqEbDhur2sO4nz7+ObpGhrNGvtia8Sysn5tN2qDzxk6Kn
j46PNV2c5ir/t3n7p3Uslpa5u+hN6LXZe+dUhiGX9P8mDMI4OtKEpWddTc2X
53gdmKTPB8lPzM36YTIbCnDzx6c4/Ravii/QRXJUO0gqZ/Uxbj8xFAYfaCuT
jfNglwlSLK09AwSER2xACuGJbofI6/pZDgi6EHba75EEqGwYJNH2oEIa/UAM
Q+GpEuyAtvLiPbG93a6InF4o+Y9nl6Ed3NL+RpF5I5jwt0UHT34YIoJiaHxx
lR8bltlbxwudncsOHMvoF7YNgOfHvKqPxGiQauABS4dE8mBWJbzn9IWMoUlF
+17F5wUM4d85VMaJnECzoPEoAEUpvdewdjoXKqJ58D4hPv4dIqJWoTGrjjwp
PvwyZPedBoqm04UbK8UL39t+K3gRBXdmI9QdzzhqIe7gOQ0eVswWu24mevLR
hAPulG7sD2MB3whY08An5dZp2l4HA+jb3N3KKsbRZ0I/Nuz6U2I39na+lfGT
I0Xpt44WDIfeVqKx9imlXbhRywF5JokGtGB6L09yjBwcokZ2VPkR7jXGV0g3
rOolXFRy1VAFlabM7bi9jlppjmaDz8qENsJAkomZ2pp5E0Yg2CM3IOLA8V+q
sr8I+YE8pGFYOlfyj7gNouoTRsgSJSHFAUJ7fiI9vWbCpbmExK+/cra3IV+/
UV0C5cd/gwQ6CNmbps6VDZ0cXZJb5Qwt6Xf0ipTrLBvU3M1mD/K9V/6/nVq6
bKReEQCSRysKLA9bT8d2P+FbYVqiqETumkfPs13YtmuSplvy9K+VD3ExC69z
ke3+ve130BcqucbI9spTTMx4AjlMqb/mi/yVN5RLCV1+Q/OeYelPdzdZ6JZJ
/Iu6ripQ2o1gI0O4vEzlJ5o8FfVj4byaZMy32V7/tIgPXg2jv1Jfi+B6CuJA
HAXKMoCqMThh1ouCn9+o8Oqvm6j9qJ4PxGzDpN9ISOUV0fxn/413Jd54IcNa
ujXz0Hxnvgi6l5wyAtHBoLWRQo+bdi9qX+BQN2I1gIOn+gd49w39jxE7mbpK
zx2TREqlqmA0saYlNYtQy6yt5v2d949wmDxh3V6du2L8Wf5zTkzN/I2IrUeJ
sKoC6qOPr/++v0z2XRJ5nTExnyCicSuKXcj87iGg1cqV7LwguAySgAp8u6Rl
fcbL9ZIXbYPmkFiBvMEjipIH87uEtYU4hK30N0wf+qIy/yuUHde360p5LR3T
9VTx/2LVAnzg58K3MDNH+4vt+HEPOdMDgHcbBR50NZUDTTF2HT0r2mRRCzBx
a1V/CIYL+gM1RDKTG6uZNZRXfagVPoRLKRFgaHzuqn+mC4S/63n44xS/GhyX
A8WiNQm9AkMtU4azDDjTe+2zvrJiaDMaVxCMfOHqfVBGeY1eDNWQCiv1YR9c
z2y5HtHSPIqAfynov8Cbm90CMKtd7pGiJaFXDpfBIyKXodJjfvJHLP8Mbx8g
tOfSkMWZTZFxT/1rjFDn4XbbKxTuZSyH1cbxXYg9rBJDxhev26PeMY1cYcjx
5mVa6qjm5and0SfBMfZiiEr3O0kLXqMloHYWo0BBALrsSaU6hTdLoyTuN/ZE
I1DpwuM2YDuuiWnwpsEbQR4IPt/JyC4Iu1bP2L7M20qWQopt/js3v9qpuBtt
/mglyXvE1pZ07Wn4mhi1dJNFpVxZEY7UE5y9qX33/w7v8bG8GnKtTwftEA3B
mmU/KGWYuUVJpMAjl/Hfczv8b3T81fyVtltIovo4Cg21YAQgbJyx4SIkggnc
bf3iP/H2Y3f/85iqKA8Bw5Q2FjMFhoUIpY/IXsUHLrAARwN1lpedp2ygbuFC
kGqiQWhfPCmm4deKbImxpgjzdsZeuDowGfi62vENiJ2R3BjFVqnilvJk05mS
n6X//nMiL/39KXCSbmlg9ELGIlDKhxGnP9SjP1DFetRD3KKNNjDch2L2xZy9
gj4UGozZzIHLGdxWBzeTvPwb4HrAI0FeKVr+SRa8jFeh1/Hy8APxZH+4sRWp
ZBq4ow/wVQmH/Xs7hsWwe2EwY+QYwg3lmxtjA7yP5o6douCGoz1v+PN/PGdU
oeZNyAIxVnMSpBnR0iIzeTU6gs8dx69o1BErx9+Fujb4/ol/6GJmTsNBkNcK
5mFRP10Y7Rea1oqb2z/92fFKN+OYfyiO3pkLEIGYdJ9vqvQca5Kr+M5xc6nS
+NeW9rcaExbRdRiWDwwRx6GgXoZqKolWSkg14BoRgmJhyMMPXQOu5seT/Y/n
k2N/IoOrl82k3VOcjZE9gdTemxaiBp+gITtJn9wzhOW0+TVB8SIn3ZW+RlXY
AXqseN5Lx/bSaqsZAhAHCk5RM2E5cX+dDdvygs/RMZrRYsf1efXAIeuxaPau
qGl4skoAJApoQbZTVyFsbB4GDtPdBnmrU8ilhdm3cv5XTU3AVmnRh9WUyiK1
+oNJ1/txUc9Rex8NbYWF1eMnd2Zg7+9MFuEJRrUjiUXlUcsi8V37C65wHhv1
Fi5YUxPwy6VUkuX8bSsfxoqIWnU9IB2Zv6+mWM/q68IVqFSDM2sPMy6QsVoQ
FD9GfbbfqHVpI2ydW4tDHQ7L9kAKh56l3j+ehY+2rRJDSLHOp8qsqTQWb1+B
heO3eYgFfzd8+eZnlac2hCnGlFJbjgIfINwRU0DxxxA4QsjeLHsbL3dELlNb
070UwjHQqC5O1m9E/3kEkagpOTXK9Ba/QPQHUk11qTrWzfd/4yv6PDwtsdu0
EZETNhPlts9ZnycDO0LoVZep0pWJ6c84aMDst8BQcor/ODCMmXEid9ryrEdx
XmJrN1bwdetxWA+L1l2W+T3lr1llXdM+uW3LdUE3+T3q4Hakd51MOpxhkFb+
0RZxlNxmK2a9HWTwDQR/fJAPGvbP/7uZFS7yZne+Pv5oWS3oHiG6wIcaI3bK
Rg1y+T7zlf8w/iDFd7FOSQ6wVektrLO6UtBnQ+0vud8uKaviPX4nadzjPe1p
KU87JuJ8RpKH9SNmWZO5IyDCKQVBq7+tp1AWMBw0fFrZIOSfb0yqBaDRZjVF
5gsBnGDZkELzoR5gTniHdvL3jYclvGkDPYW9ORoI/bkO06DfCg5gxGIyzYK/
Mvle5Evh/OuSzR/O/slD6P6WdbJ31Fw659/5G4tWz3Hj99CkhbVQcQELKm2P
Oo08IoB0icnwO37tnGFr6Yj79AeFRfS4gfeoWbnVVrMaDX4BNDhcLtMs8Mpd
nQggKg/miqcI3qa8J1VcFUHvVsja28330sww8EE7cwCFwUNbXp7jznP8ug17
HusNRb8dSo1YdX5XbNMnST3xHB/YXvxnTtZy/dbJa85Jud4Io6Be56XwSUlV
rhSzNouuKMSPdDkKZbDYAhfHoJvOEffUFkM4YaswAoq7pwS78EqEvVcdoqJJ
JzUPEfunEGTqjZRHIxKAd9EA7jwlwFLP9Pw9i2+Tq/+MGLf1RDbcYJIJ3dOC
kqMwJLErCLHvVFWjhALAL5Adee7jnx3NHuOyHd4L5okBnKd5Rhnd/+xUo5fq
JkkxmqFgw0XAbOXY+vwjHnxK1U2AkkPrr9Oet+mkEzxz35rdYf4loXh1t3i9
pqu0GF3bWLVmZyQzhDgRJJHCd6ern9dcAPTmnJfR8JOqslaltHLsYq0ON3+Y
T0wlm5HTcPEhDL1a95DXS9q6ta+h2f9WxuewKMYpp5KO43M8xq8NK38O4pAa
nFo1Id9h5ZeE1SFo88wjHgNXPi1nFwjAynwT3D4XSpxgQdwqvSr3OKOLFQ/s
tJIzgFG8bv8S4hQj7OBusgiRCZLUMmUGDX3LtNncuedQ2e9cbPCdNwBZrxRC
0AtQ/Mec6LyQ8oa5AYVvrdf6Q5Hez8XTnWUkdDxEKtBU0u3SnxOWzF8wKsiX
hkaVegv/0Yp/+0QF2lw09h4YTuJ+6oQg50Q7zhwLPFumRzoUMOhUBier+CT9
HwZxDP1ojw7O10pbcsLBZuAgldBwvVb70CrjvVoa6KJXZM/9Mho5/57H1nqI
mifDYc2WibdXMpYrpBE9cexeRSueODvp6Pf3Mn6g94JbHjyA1vfDNRxvvgFu
+4qaVy2pOlNvb7XKES2sqAWTA7hZYzxxUAyp3dt5GTcu76tMHGkB/djUr+z3
c7DnREXimQOdRsHGthA1cAJh1DZh1BdVfPMc2NYxVZseVH++mNxsyRHMfLtg
EyZgMWBQ5QiwnpHxPtu/0BE6rEBKmhcIfvdLuWYDRw3XfCdGRWfyV4JLrONM
AW4vCQKPoK7+zWUPDbx3tyHQC5H1wUEg7A8iaKVtiq069H7tr/eOFrQ+JBtw
5eUTqTtIkFOVMHDTOE2Fn46BWbWVxwDQ3s5P3vWOYUksvojuQbi4bkQfgV6W
ysfFFSh2/rQlrcCOvvy5FAyGHrSRWqFDlQBsoDtks/8isCh6dBXifutDJE/0
xZLaU10e9ONQnZFOnS4HZtHjlkXGILqX6yJhQSTAlJuaJMHtiRbZdZiaOxKU
OgpLW5U+5cnXzNisx1ZEZnKgrh2VbYy686yIUS//fFXSevemgf4iC8L2ZdPl
Jw96YCnXjo/5YiHT1djnTYnQyOzwF0kprEhgUv+hBMuDQ5lS6Yu6ROivtXtX
Iu8E4bm9b2TWdgVGgC2Dte4D08Lk43DZEXpRwMFgqn+jJ7I1ofiUZW1fmIvh
UymgNfMR7PBxHrsXhknR7G02bIeGqIhgLlWj6FEdcZZAkAqZtDFyi/uaWEDP
pXtIooPFf3qbv1PA2q6gizxSktN0uJw2a9rWQ3TgaLLEQ1WzLrT1/Di+MeFn
jB1owidoaUnNiNGIz+MNbw9gcnqivItiu4lwI+lkbEy5dGX35Pfq8bjcfZLe
CkoAzpg61NaZljP9zeveItBwFVVEf8Qrq/hPWiE+5bm1IUoFliym5G0xS6Ys
KmaOH9pK92JVSzsHpqOQu8GvA51lNzewae5HliNi3ZeCu5AO7P/ZfJTt96dr
BONbvOGKIwJneBPVYpyky6P9JyYvf3Tb1NEA3SoxqoW/Rvu1ANORf2lwTdVe
DO6kwyxzir89rUjtIILlbF+lFSnQBqtKVzt4hOImkXbq+d30WxdCdiMLee4D
WRBbiVLgqwu1zxsDNnS0MpkrAFTV5vKdGKG//SNAKraJRZGfBdwsiDjXY9cB
TSFg2dNNHThQ/WrmsjIgU2h705YptJx1Nw+A3L+glqtp/4KiV1Fte//a4LZy
GdWVL4Yyvcli79YfgKIpAPtStmC8AQbwym/RYhdgS53P0iiGPx2JdlwJzZUz
X3S2kqFd7D57AfsvfG/wJfptIHko114zuJBuPCCqbBHdvE2Wcw9BY/cVghCT
pkTmQBisVRQ5GmV2TjY54BqbotohDRRaHgw8p6Y4VAEw3IOtAHWToTKSWO+F
o7qEdQK/GYzhZpF9LlEyLUQUrPNlmWAcW+zHB/Bcqb7LFxSywn3SJU3ndQBb
Xz1HUWEIwLvmjq3rFNqIEvKw6vu9JbXnhiTtnJJ1Bh1irftMJfG0vjOBTri8
OO8MoWcfFn/bjYyNxokLlTLiKYP/eM4KT58RgWtFO+apcW9f3T3RfAGAIuLn
3aKl2oGA6PS4fs3okw4iiyBfibEb9lA17/E/M2PxzqmI7JrKx5IJXd5kDOkJ
ZsyVN7rKXcsR960SfSreWC/m71hqH7kxfuTRp1lVjjSqEqIFpd/ciE2MIHgt
UnNrT0Am+gdfVMeBuxn0QAZT/1+3BYC0hEvNmIdq/4doa4wE8q/lueGkKCt7
bzG0cGvsn+pUiUnsOv2j3Eq4LWsigkdEWp+vfSosjeFx8K7MVQeYEQsF3ivT
vg5d77VoED2zf5wWzjPsP+Rgm1eehu1YoC3F6KmFa33z4NWdq4rcmzKzAH67
tXO7wA4YHs/NFmFrGJ+ijxRm1TXrnvc9FtiMMLGMTX56Kn2SDlZmTuapnPyC
eYzHk3fmW2vZ6KTIdeHeHJOIVMh/12+aYivyVn9lcdSITZBP4CWr0R4JhDTx
U9N/H0EsImRl0TIywcePfZPJI4k1Rki5NJ4m26ZMMwRlW+Sue47PGyC/B+7J
D4L6IIsFu+takn7e1VCFkZoVO6TOZaRw+afJTxkre71/QcYdXur7126sm+lZ
kFSDIinVcb8iVrtIooSOh8BHD/mGnlxrnkNLASyHrHsw/bDZg8wLpw+/X0rq
8miY8HsvrdXcQUZjSE2PSUIxEOB4ZCR6xy5k6mbiERmOH+HES6bGwMUevIcb
Lqu9f7W7LWCetu7O/KMrLKhmDTtMWaf2dBu2nI79RvagOcXd9g4/l04WFRJU
6kTFQEXC2CfUuPEUR/q72L0DPwLQcRfRsFSD+ttluKXzTB4c/YC18ukr5Cb5
nxfXSU/IlLGJbERx7JlZFh2qHNnPQWt2x3cmljLvHH8FRaTGuz+YrivE5g/k
5fCO5/IqpgQZrFTs6chBqEEnXVvNa+3cQM6Yg9qbIxGK8md/WrzvJvEj6svL
383gQYhd9K36jMEij+Qtv5x3pdIcOFY+ROEZcBrUnwwQAra21vW9DA3b/iHz
LOPmxejo9/Em+1Gi9cIXV7RlLtwO2u4QTjHbgTSYyXw5gMTDQOWGVRiTOtDN
a7Mf44m9sC6/yQ5sbG9bzr3sGX1Ra5rrlP+Bf23TWGZ/hjS/5BLQVyXqEtCG
h0pR5VyP5MFedNumP5tBwAcu6fB2+jkPgQ5zI+cno5ZqFE2W8lIiZxlCIh05
fx/C9AjJ58GEwLXYUPdI8Qp7RCDyJsCB0eZerCGRzrscTdJRJEnYZsZNDBg/
l4jK/M41Ld68IT0QhZ6MhneeFRVQdNxwCkzaRf5nhOLQ64GS/QE3TSynwWN1
2mU3xAqJKsWykkBhaIyGSTevtoGeggaBrLOu9YwLq2SagXdPceDKWhWEwn5z
Bu/hx7s9BZqqNOgpfKxvY/aWcmUpzaexiNRYm7FKX871VqySVflJAREhzXZp
fzhNSgP9lO+3XkqHEUY7dUs2bfuDf7hJBFYZrLRTfH2snvxKcSDDaYaUQ0yy
Il2jZMGAaNRAgI7SCn3vEljGYYEZtYji1UYKM2dAvPWGCBeZUyWf66b7JY6o
DcFHRO7xahTaLEoJ5a5zDJzXAX9gHOa6lLzboXnHW6PTCaiyOMGDoZbO661N
a/ISprSK5lfs2A7I4eQlV9QNoEYkL4MCoJuvzZuYuRJzEjqpvw4qjwb4Q2ES
q88S5Ntw+GJ9k2VBCWyigDOsC3Kl1Ub5LRHU85E8hRgerGbmjj/ONQWh5UlU
C4bAkfbzBBJ/ssX8mKucvqSfZyFwwVxCVJh9gPsP6w/HfBE4RoCRzNZnTpDk
w8OyiCz6jQ/PiB3LynKlw9ngANES+jEH2NoRitOIOFC8SJnEvyMu5SkLBBc+
ekXOMbLBaNewpqW8AcAS+cgmfdE1DuV4x+hIBtXnQ0vlfdZJjakQTuCRD/qG
nuamxIVuKqM8XDw0Bp72eMfWt6SF7qTlXXjF9Zsv/K9sBUrexF4yfgBM1STi
4c+5QDZwKeoMEkQ8L2bwXrGA9to0HCOQTUQFIqSb8T3RyNytxVI92OmE5cHl
VDlUtE2w1Rs2Y5lWReQFXd9awUAZnm6bh8G1YHVDGenvRouFkdCkZDYIiXZ9
D6z9pwHnUPeE9tMs04TbancnUWWxrLVYENaWzENF66vtFNHtuEoMx4yZvxLD
KySjCO8af0/MvQWeFfKoOK8vEXbvIiRNaUmlww1kcNiBYldTqeLi89nhAzYW
JCaD4Cxu4uuZ+/3YGI2UzXcCkxppmAVtzqyfkJdZtYDPt0Sv7m5y6J8Jx+40
P3+h3rYOFRi/i/ZIuHvd83Ognl6n/VcEnUT8olvuDW18H183HL76F55Gn98G
6ZERM3U5Xsp7fq/rpRPl0Zop0ymNLkG4We9resmUAEaW3kSqo0fTCq4iPCiL
gtPnSwWM7+hZYj9khhH2PsVmcuJYsw3igQOa1OIqjDj47gnP99/0AsR7HEjV
YTxy4iiSOVV0qKZzobvj4LcKOazW8u003ZDiiAldrPuci9pwLlDX6OIs8hZb
2rZoeCFhCs8p52bPrCr0raiTvkpnYHDdubByhWCecbMRRdwQmW+DnuGDmiGN
i1tcjdb46cmLec4NBOgwqNelNrTiVk04DzeYPrm7FnYJHQNSaidAJExu7L9Y
FM5hwd6NhDPMUjQrsLo8ENrNQEHt8Kn1B7HmSPenTY/t2uKO9eFQLVoNJvy8
XatOnSMGXv6yoKqFRIeLpk/CDgpNFCgAVdJvdiVq6YyGf5PPhDT4b71u6DTV
rNVcEpm5Yo58BheTTmK3r9ps7BdctCWB5nUikwVEZFC827VTXQ+vHNCbVb1p
K0wGJKzZ2VrB8WIL50E2pVrt2T9T9+n8xm3XaelPHA+X5RgpHh2PVsisejb0
R8AV17/+P7pw7TczCwQw5/QnCdlCKi3BeHqqjnm65dfu7gfjcuXZRS3x5+Nr
NCTMU61OS+5+bE6eNA5bzRRrG3YZdWCbVvGbkAkBRzXH+2mV2eEcauin4K2I
lLq7g4M0ss80fOTrLVrufv7Xp5/cnyDW/rYbZFqyWzHl1wcmQTz8tvnnhlYk
ifWL5ZiuBKHzLKlvTZZ9j1X8XzJIPBn0unk/ZONxGIoK5izXYVxMVsg7DfRt
7CGzmXGCvK0g9Fa2TjwwdmSMQEZQJb7oPrBeG/1mgI7r0AuvU1vBOd4C+D1B
GRg0XYIKAIaTd7/kLsawOHK/0iXIKynfCa5O+hCuhN62G0Hn2xN0rNbltgdm
6D29C0maa/7wJK2NMpRx73K1uB4Go0sAwFgwuKhBQOyt8xv/rOvTTGxjYEoi
dh+ncLGzGo0KM0lVIIWEDH8IazaUwgu16tHPxij2JEVkCN/04Sysnf2bqIDf
S9pjIoO+TCa/YP/sLFWbPDpy0j9/+lKUEyX2bP53C/PvybpF/VgSH1B1goKM
uvjb6RRGNyuL019KgmVICgnb/TviewGA9t47PIgVC5rJN06V2A6rDr2Ig0uc
XhQBW7nEouxw7L1aMtUudvHSbuiWANSuks1bQR9FU8E7Vtqv1QczR5v6EpLZ
y0pETxaPHFn/TIUPfvH7BX24qsYwMISH2Q5CVctl+Jgdjsd9VMMBMkdXPQEK
k+sJa7YyUlbxAIY/8oDAUY19HuQdYaNx2Hf9fYhPo7r9cqWXQQScG7OSAOd6
zAoHje8MeXMo2UY5+peAS/+Pfd2Ik5keH7yOpPW9qOAXA5ZvqyXpoadiw2C+
YdzF13dsALW80ncy5HQa/QlovhqdRJ3ILrin3pOKxLSC/nxsGzEGAX3DOVda
1UvWPQMnR17rwopszYl9yPbeXoe5e6JjS8zGJfb9acNdgFryl3TE+nX/V0ts
wy0G+mRo5EmvEr8xxVMcWI0YuM25MzniSHvo3FFKXDr4i55A2lQ0vowh0ScR
hlaRUnNi9ExkaFk6GtCakZywfIVuorVjouldbpBuhkGI9Jf2Z3/jjgeturNG
1cbIPZNiJi9R87N6KvzCz0v9W4tz0zj1DB9zvpBtxroOKEktissCX5wjqhDr
vr19SlqWufZwKI4oT7JYlcKh7CIh7FlZgWGzowiA4BTGZEcnjgrP9s7jf0az
mfMq5Mrel7ZuardUBKWHiUzRwuHiEwrLRzKSyTv57YXSlCrMapywF0AZgjzQ
mTs5z2SDRXeh8DtcOE+5u2haJpIJMVQAQ96QfUHNwz1m7Ki2nl47E9MFWbud
g7r8zd5AhygUro1z9AYlC6bEMg2OcyLgO8ULaakaczfnENw8H9bmwI4oL1on
gjEW0Z+WUE7tOGHL5aKAN+qy0+f/2BKOQkt3xjAU5eAtik8pf/KnmPS0Z6tj
UaabttXT0HAzEzg1GVnjQCAXACC+7afUdG3ayeGBCtDtQ5q6PaIHldv6He58
QFkvxOYeOxrhPS/DywUHvoAX/rNvTGN76c+SEEU9YX/26vKs+aMO8uYsAEit
6+3tGBJTBJMdwm3tPh1qoHy73FIV2WFpbibREgK4nrBstBb9XJbd+uWIgMFr
wrFs5ZLFDPrCjBFLtQeKy6yz58zDyjtChIJ1zlgT5Ba8Lj6+jRbqKW+SyvUU
HKODIakKGncxiIQaOipJAJ2X6+enkDnGzx1qKARJBn2cmyQjFsS8yZN5Sgrp
U8baNykN95VBVPbTRHP+Ri+csSBWKDP1tA3TGw3GQtXjd4s0t+JNlPVLiakl
QEJrqsr3UaxZdXuQCvJ7cyyj6mVR4i0GMAMjdbBWnzmzd1eWu/LSG1L1ckSN
muu1BvoQuhayKIrEQeqe9CtCL4/wvbK0/UWZBnQIH/WaN1p46osEjxCXzHNj
NRKWr74QxTKeEKxx8IfpVNJmujw4M6s+r+5SZKnm6DPuiDtSFl4BGlsDrXDc
omWehaGDv5wS8VxTJthM7FATl/0t58TpvECzv1btOLlYAaaxtsNEYpEYPWNv
f1mDt5wOTQFo/YE+T2ZWJQHF053XJOsYtMRaZ/eKSdvrMGhIOu5cGJ8a/OcU
Jux/lDTm0AJ3djPAaHc4iPJ0Vsa8ixFY5Odk74xqoEU0hADgZ+1ozPKXwIkn
jLwD4T5MSiSwYrJSrE9GILfntuD/4P/9PbTmQgpJNejPIdLaESO5JOOF3+y6
kLqjnFwRNEL3FT/rlqA7NMvo2CillC3pRY7qxVWx+CAYTL8DO3Q70Vzo8jH1
lgpyfblTN7JUtV2tH08XsWS4gAoz7XcjBPhyuNdzoAySSXmU2b+n7e9z2Xag
lwLFYSdKW98vQwUlNoFesUI+75UmIXpRSGwLOnxKaUQRJYsxn7csqGpI3Jsy
sM9lXhnBu0jNU6hFMLCGfobRQuGQFElMCCsTdRKYJzevWeS8oWWUTBUN4Klx
ZbTuJ73WIwf9pHCGllPhCAvt913qHPuok8n5nwezSHKZZhSt8hdIHJxfX+XA
ItGanyH8dHfjksZ/ZBw2M1QjA0aTwFW1UPazZeRQdhjRcWVRnuuv2GDY5Qu5
X28e6nFSEtrRyxsd9OOnxy3GhVNpo5P9p5xQIRjLewwZzjENdq3tFwxcGRUy
AgYoL1nY5rWCvQd4fGJ6aYyMFxMx9z1qIk7LLIdGi4NLAJfbCo5UYO9t1dTr
hKDVyW3YmbajqugOqu58TOGtzqNWV/Zj83lYbq6KCyQCIMuHvw8/MdHNSVX6
Cv0vXWSnQSiLoNTr2OZnosUjPvAH1kCBrRpFwqi8oFU9Zg2OcgSZGS6NLGS7
LzaIe+7hp3G4N9tcle6KhNGW40vn5LfepMEKG17qsgJXsf4b0XPpd6o0ydY7
ss2aS/hAuYwPzwLajn9SmZ9qbF9mFg3LEXzOwqQtcLSIM6T59drhidJAjor1
n5N3G9Xl+VSiZd44o+zX5MRUZFtrG+R8E6d/rN6S7GwET03SsL6QOGqr399+
K+PdVa/kKYC8MxWR6Xa4xV0AKPvKDYameQQYzd+cOZ0i8f4Q7DhyOnlEGFFG
CDga9NDYe1Knrhcit/rV/94EHoMQm4yrQaE1/AfJgCWBTL56tsZYj5m6w6Hr
zUj3+MFWy05PTnEJoLmQqRJW/P9e7bg0C0AekuIxbV9PXAjKdhn+k2l449kS
zmlVV+pADtIA4sbadUEw6zj0o9OozcFzgflvGOItOlrp8/yjfSPffbrOvZ2j
DSgcQlb9vW0FvTgD6K77zIKjNU+LoVAlcYycLkgEgrIRURTrwdF4XO9D3lgV
2ZdDTFj5wVy7uWWG4RcjJydRBWXKvfcGaVthC9sfNect13GEd/fH/ezxTeyR
SDMq5qVmskuqOFHWcqw1e2qLXhCM/qcDCAcMu3fqd3SWjiV26ZDyWWEzFM0e
2psrCVRoTAKgG9uQjRlumSfa01nDeJJMrTidjhQZlAy7TuYPn39z5NMEXfpa
7KS8ELjNZPROAICDMGIFZxuYQSFjXBT1gUj7TeLWtGUSxcfv630RTORvMF8d
5y5IGJ5rChTwjdGZWL1gmMj/I+wFtudUbFHwSXybBh1u4GO7gKt2M4smKmOb
reWUlPFP4q3Rrl1vU/msomnjHvi59Y1ZgGGkY/UqOI+/iXlMITjZagN956mL
r8b5kjYP4ratm7mQFXpupTPLPRLQw4hmZxzungwb6oZHR+zZzilJYLu2H6Un
piI0zKi3ltkweniI64kEgdkbTC/RmcoQxCCN6zgrWtE5/wQINq7SD6e2gzD1
imF+J+nwHto3kX11VEIvLKI7NqDI/LBOJ+2mqjsZGVAXfeIUQfOX7WT8MN0L
QayU9PwXe+h+d5jfT6ST51209IfAhzM7/TfwmfaTNAyFxosYwAwTt731CkyL
kC1CJbbaYLqX4dfmyPzwuslRQQf3VRUCuAswy3b7t/qOFTw7zttP+Osk4vmx
2jrMHNKrslG5qEENlgYhZRB5r3O8BwlYF27zLFGzyKb4NncNc8uJ7clQsSKY
/ALUOP2P5abS684OtSbglLc/XJhz1XhZUlm34svrIt0jiQxnaKhutJZ+p/ZS
jkS/RBt34FP7LYzpxWkXSCOkSrfiegAYYbrHBr6RYBhGoMTIbbpr6LoF9/hk
m75hkimhxFlUutpOFTJH9RLvFvrF0TXzaSQNambHk4SEBFLBM+u0VRFQYUvf
Bg3ODFX6nrhYODkWvem9WRcabkHFwjGTiUtnFicc4BSQMsCzt+UPXpJirdgE
boWj6yAunPbJne/YL/409F8iLxxwpJJIFHQMr83dgej1araQtXobC/KAHegD
2L6R//SMu3m10hgmgEXbG8y+NaR21KvNsTeg4xO1Fl/OcbxLnbw4xdhdoHA3
L7AEj1xwpxjAX9D8joKuTN+ItlAVLiG2d2C7fSBRAh5Vpt+YkO2+TzmJnjAN
H1U+fdItCGMlMFti74Kk+q2WbCw8DwwwiVaqeVwhzjCIYy5AnBp8IkyRUYBJ
LLZ8kbPgt7GwlyJz5wyp9CshoLOpiQokjrNYZGqX4CTpj2Q3GHOYbFBG3e7z
zMoWAZj45b5BqCNKyyrX+jQVL0PKoyTR8wz5TdjSf2DWRQRM1ariwawx6vDB
UTx0Z7VLMzGvk9w2A6Ek04ki/xU54tzIDuG+/2xyzlYCf1bs2lkxJ2hS6ko/
ExqFNK/P3R41qQYYLuJ2nEf855GTS4r/cdr7VFy8vr2NGE1u53Nl7Scbxdtk
TIxnm5/ipV1/BU5uRZbzKCfT9CBTb1ou8nro06i6TuivjbG9ZfLGwHiOB3Pp
L8NxGw5cyV0VqEmebGbyD3EttUisWHHVedTadg0Zr7l7Y9qHMhd81PxtEKsT
+IKiOvLmKgBnm3flKH55WPoZIhW05Ify+80H0pwoqbyzgDFwlKo8of9daoo+
EGOT490ANwlEw5//k9JHcjmgM5W9O/ObyBT7zFbtVw4ExXDn5qhM2zL5Tx2O
+zG4dgP+u84GcJYQLIzJnL0Zb2D2Q5dFxWoA0kKT+Q4caCUwZd6zFqhVz2jl
eiRmBvBPtVewf9Bnb+2A9RRTKuVBC1W+ItcmcYVkJBoyo4SJaalE+l2yhXly
3gTX4hm5cSYD4J+RVO9bvVD2FI8FnfPxELSO+SPjWd+igbIdr/pvGk5aboCr
gHV0GmSksdy9UfXRFGdzdYjiAw3fXhAvIwTpr9q8xR+oZNSA5TIP+wK/kh4q
F67wc0kzzFq7a8NKsT/9ChfnW2DMbPoXNPxEFt03y9sVxIyiV9l+T902LzYg
7+fI8WKG75OkzBffCoixJFuC25u3pUldVzC9iQRz/MtTWvxHEACyzuxFGt+S
KDOTVE8kSlj9dE5nOnOLpxc3hLdWwN2PVGYN57tKLLIRthrW/JG7sv0HZujX
ytwAjEkECFcrvXX0l4WBd7UGt10TOr1SRzfOp+2SaOFm/DIgd+W3pWeEZRIP
mZJX3oTe+6Hf//YlMz1ghgoDypE8EmEdKteD0s99l2GfzPhZ4rseP4Pyah6U
p8vVYR+8UUgq2Oc8eGWar0HNHPWnx/MxUxFLc/WVZLLHVD2zmRs1Uc3LTCzP
D1J4HYgNwfglyQ9ESOxiNw1VSZl5p5Vcr1R99xgJAiSm7GZ7nNYfKDh9Jz1X
oUeHiMDghmxloDSUX7hkumIGGJWpKv7SP9Ar5uK4YChJvxbbETKfXAyKa6DP
AAWEAgZKJNngCCZee/JCtrjSndFiUyAjtBXU2dfgHG1JF9OJsQGUE9Hn3VME
IhooefQ/+1DAB2tf/cnIAazgXSZpkWGvOkmZhODboNeMH3Mel2trjD3bbk3J
WYqSxoMtR6+2znkBY3sekJ9jtFb1Ib+yAjX7kbWZ79+5qlIZBlDTmKPj9xWd
Ptf3UgoX1F8zLky2W4jonDarZNMFrJVz0X+VHpdUPFViWTx+/sNvh36BXvEN
AZuMlsQCQOzBxpkkiEUGgAtTGgnG5Sc6OzLn9Q6Bg7ijStauv+EnX74Cbrwe
UuLTIsc4TG2sARcfXn+NcSu8x/KFpzRWm5Yhys2cS8Jdiu6jsafx9eFwi7BW
aQpBKNrurHlhejKUEerr1N6EYzWX2zsaGBlqQiregBBRPHqlhIUuR1raSoyy
xc7Ot8xLRUyTPq6NhSIkJuZ11eYjqJfAKo/9rHFCvJsB8DVfVdVaKZF6WsAj
6NPjBnh0X1o2qaZzAW0tnSKduuFmNzEAqfdUDb1HO4NCQoiF6appyvphhfvj
k5yDEEiAGH1JLvUN242eGdMXk7OiheSptHIdCLT3uPVlqp+QODlh3Uss6geA
4CQ16jRZW8tpXurWI4Fqa8/xe1wuKXeUqtXrQkOfiZz4rWP1Ykp3wQpUdCaY
U/Mf896OxQBk3IYGTn+m53caHBZdEZgqEwHgsUxUQ7fS7KAuohoTTjuwwAIQ
SJ5WYZJkq/C2vvyizkNadYX3+BX+wreGvI4ckfZ0yxnsJjD4e5jZa0E0aqnr
FjjESbJMIjfQbgTv3CTNOv51L+xR7YvQVRxNOHYuqXEdrKcr1BXp2XMnAwEE
uhUaIejCZ6KSj4J8lnidrgMQ+XD6640LUZbeZRewQ/EPgZtXH8PLOqz5HXPT
OO/E8dL9x3Fm46uzHzog5UvPfqLmSLJxn/KwnZc+UuLPhL1wcShcF/8zLBPp
GRBt9Ok6HPecL20fkrZZ4HsG3fTqqYmVkHpUu+ldWueHjdJjRlW+mOEt98mh
CFBeLdC8cD89p6wRBOJM8cKjiuRaWZN4d/m/PETWdKs3xOdoWI57BtovKH0R
8ptsCr5In68VmBoQ2GGQ+r3nN4BrbtwMTjt3UjLbLhilVSPQQHEpe5Hwu81r
aeD3wubV+DflxY2iSzpSrY41EmCE+TuSPWDtqcsq6ntqzo3phIiOBBUekAX5
9l9CAAL9BII0/17u2HWJ46kiH9KKPrGcq4NXsAvU66d0WA1Owqch89RaRTJb
d9kRpOspNcoazW5BroSI25MJlF5g+YIabnl7ykcyspm/UpXqiXS/OytzxH5e
2lcd08yfdnLkLjt5Lj+lgEYUQu+nrPP18q/e4r0Orl83lkCs2VqICJcPfdrD
nrpogDWy1HHDcQsJ9cXCn1TbskDjWA1KCs47HeXJMkogU0LsuGaAJ3mvD70E
HBGxlkqBwD9gX53Wnz1BXNQelbMco4V9gu9T+H0LR02FoB5JpIqM1hvdzufV
abshHNE7AI5K4buDZdPvq4RioORK31RO61/qhM0ekH6VWnWN9AiEizx4lOfD
Iip7U8Egc9TcRfEq7lzHpyPRKH/fbwU0GyliBIAVKYWPIB9LD1NBLW5QsHx9
/RU+wN79tgZo1JnP3DvTp/Xo4z2LKRyozOeHoMbSMZPeR3+CQkI+X8wyNO2w
vp4piSRIK6iwaevk/Z9W0KL2a2aU1tVsX+UxvojujsteiYfEWUM9CyiRv3ID
wcldoxIV8cfJNkYeI6IwPc3HRj8jBYsNufqdEsp4ThMtWaSFPHQHgVisHY9I
QrojMY5q67N7T+MgYw66sVSm0Y5oRxEL60d+jBdlL5S6RtIchQ+424ZfUHGu
Btd+Ux5PECWnb2oNfVrCJO0BnmSR9OR3C/lIOidOClO2/uVKy4+5//V8TQfT
JWrHGMKBQzGjME+tzQjxmaum2aFR9h+nl8hKXvH1rSMZ/Z+7fxeg55gBClZr
z13kFU4mlo0VwOvzbF5JGA+6xTS2mKBs3R1AYETZACSfeq/Ua83Zjyt5i4XX
1ycFYmkz+5S49Q1sUcYl/lWRMIHHzs1ldLz2VW37m2zZ4Sy9wOi5iKIbla6B
BWKMfB0/i7B3tzC5eT+GGoj9qXkPrIFq5B+Ww1bWoJ8XInFsGgZ5esH241qQ
mF1HNdpGmXf+WzAdaMbI35N0vz8m1bTb3wHKxZGXEahDF6VmzKkIZ02jC06b
TW91Hn/sPRHBzGMujLiazpFynHvWQw6WGAzTjSkoAN0QUye02tN6yneJXQ6J
mtz7IMYaZzE5IyeKW+d/pBBLA+F5Ga8RvXVx0wXsAzJfmdj5ETF4DBeKY5Po
DjT6ncYghztAS6agL+TlYcF6dehwmii5hd/eFv1RWJxHQeAc4lzpRt8epHHT
Wvyct603Lza8dD2JCCgLeixg/C2zNdDgVgs9xVg6u2O/1sBhmbx0o69fB0PM
x/ZDUwS+uywbdOxiBFE8Gq8RN6n+rpbBc5vPJ4/YtbW4aJ8fs/sn+HgO7gEM
EazN7gIGo0qDjlyO58vgM6KJdevrMHlRxkR42JceKjmwTwhmytW5YJFt14vM
A/8MZnsaBgvlbJJ4Tmc0Dl5zKH+Thz+VOwxvp1N4pCb5iW0ib3df8WA1iImc
V88gZHy3RdcsGi7A4BNoxHCwaOff5VuIjQhedI0eflJ/lDlqiXvtSlqNBfHg
afq+jl+x2kE1YO+Kh7dIM48CgE0Ua50H1pxi7/zDebRzQcGoHsbZIc+RB1P9
K3bKXTXM4eCunNkzpYIIU3nrVxXSnXVbTwPFgUazZZTumhtgXMtBAHX2Ehmv
lC5Ru32ur8vdkryhlaPYK2ZaC8TRY4wpKO096ErUYXJDxwtYljH1cpwKZD3R
8zp888JHDAxdqJ0ibSttFEdgByMpb9ZU4LIHC6IYk9TMX+hWDb9ER/EDlIrN
JdWQJrGZKB9f9/DMjzceT25nBqX9cKQQFobngbiZazLeKhqeTRUOI5W7asnk
KvKkowlKUmvP0REjXeLcotWaMk/b80xWJW1uYiBO/z/vEutLPNwWrBxhwIbf
9Br2FEAMexI1EHBSyMq/Az6sCw12u52uXchBrqIbaeYlMtE7o0NpMfA6eAZ5
ziDU/TMY/1yqe1iRo0UQPFEuRmcfIR8y3SrCFUVNQoMnq1AK0SqJhbo3Wxz/
+KHD8Grjl1Y91ZfIux5VVvCEfE2o5C3pMDDCYeAEU/7ZjRlr9nqQnMUzTJxq
A5BnUj14xkRuRbYtGAbGbNsqnC966msLqx+U9+Cr8c4Yu8wDjHUlQ55SbGJw
JpWX6wknlDpiYrlbsE321hyMvuBhxEsgzv9kxeJ9qae1DIW9XN7q8Qexn3gM
u3E3NNGK07aZUlq8cA0pHc4BwW3y16KV71Yc43/2YPoRN5UyzeViG+V/7nUB
Yhan4ximccAGw1Tk2VPI+0gRugf6SxVu/RFCMrsdtHbXWpSsWTSE8vqTXye5
tmn/SUwaEc7cPcMus+xqT9qGsqucsEyfNR41SR04fQc+QKLt9DvAVjr7cwCu
E6XT9PFg+PwOkhUyL471QUMxDVKTNcotJXc7txX4AcL/iwrxkMF6AU17ruIY
tIjkqew2+r/rxnruZ0ZJKXiuWhZ2ncZp7KpGsZ1hR1qIVwHbPurQKiPtzBf0
brJU5b7kpt4enncTlzFn7vgce64Pix+2KKFPh5Cy3Sdz7pIimnKlR2NR+K3R
59a53xF6rZlI2bVDeKfOJxECXempMJc0D35GDHhI5tRAnNJrREIE5bMCYnmk
EGICuQSS9MH+mvDVvT6Vi4iCSVnnV3CDTYsFtqguABPtMp1zY3uwb+N4aIzO
ssjefWH9CJaJOnEjXNsMYsE+r1GJQy3aald0dSBKuk6Gk0XetT02WrPIbtVs
otxhN5tBhXAjKC9E6AVQQZM16rdZ7QU7IhPRyyNIHZNAR2cm+SBvRb6gDErv
CdmZQfg0Gz3RfifDsv7oL/w2IIucYtBlh2vjwEnKY3kdPeQSTVxxSAs/NoXR
yXeO1n6RrYi2W4iG4nblPkuZGszhA/2EV9DAS/J3QEo1Ohbv3UdyqpyXNjXo
mT24BVA1hQTE7WYRVLndG49jQ+zaawC/6GIfTiFcpOlwLl3e+AM9eaiP4xcb
g9J+YwVl5yn0f2xfbW4N4y1J/9GIuy9wlqqAzxsotG67Qrzk1/avapkocjnt
SWQrFpmezwa7yc246TerJZ+CNGUbQyCP6555q6gxcERbCrvsGMRA6WX2QMdZ
20JthNcp4qkWNGkLN00aFtdwhqpkjgRsOJ4asi/DnoyrBJMRMr5VdpWyznq5
ok+GPEXe6ngdQEh9yk/ajagRLppQ/Kam6eo2JJ1KAqlS7q839HCXCaAK0Twr
SNGaDvcKv8/0iK+WPh3me8DNeVLT0TwNT0mShNRpKxHK069HTr/gN4f0Qr/7
/QEJDCEIyp94Y15QMK+wMlqhRKHdOMTsZfXkR+E3FD2LbTII2ErXYfh9sR6g
ZBFWUVVCgSUqxMrPJNFyqaBenfYvnOsVUvdfkmphLvsTf0FRePKaxNsnSrd3
ste7Z2nH3WL4+GlIu+fHygu207IVC2Ibrc3F9yo3IB4tar8FIZNlKXRC5BmC
/rtcGNj++91dVh8/TpDPyq+11E2FDRT5skoqUIx6dCVXcBB5baEXJJz5PSto
kzlw/dNKxwVcAZxjEEtcFI1xly/AHVIA3aKlesPmo8KCKvOa/ra/w7vuxszY
GERwry7oMo1W3+35OKdZO3h3iY6pI3bykI3ZsCxsSB932EZz/LTxsYE2EJGq
MysgiyJV4jRDDjng3a/foq00wcxTRano+YvZ8iyqBhpxLiiKQwD/51Yp6wTd
2EDLSqnmeMyjz9EIpyGg7/ZhQaxpNs8kK9aFLMIenvdBc6h5BGERsQSWNTHh
P39NCqiJwcjj8szU0/UCS9oDMlNAhF/L8vgHcUp7Et55TDFdu2CyWf6FjB20
eE55QSaLOOlUgYvT96/sDK5t7ZYfWT+VbvgKrCzM57UugMS4d1p5LHYdX1+B
y1KWQMt6W+nJcXXHY8Eo4ZNdH9zdcm0b6Td2OH0d76XcUbC0UhgLFNS7hWIu
GadsUFJuVabjnSMpztJrmMK6rLkrMYIA2ONaJc2QxRSs4Y4kvkXGMCdxq4aO
aIltl+JCgEG0mLFHJqay5Eq6i7WjZQmxjqllWGVMYzhxeBTNriP0cm7abyD2
rtx+bqnxTgNCoLq/XCL09u/IAyukHWK2u0s5HZkvq5nXqT1rPnTYfdotgOn3
DUqnThPUw23SprEVvbVwNd33an7+Qt3O1y2CpBo4KEiGM5eOCNrVQ7b4N+Ck
J8qoPvyQKogaNcGJtREDOyDkYidck0ZXBoo8Sr0iYk6bryJwTXxmGrKFKf9Y
HI9juAywfBW4oJDQVR0jIkFLOez2BRPPgSy7v81WZaxe7nEv7mNRrhLbE9Jt
2k8+wm3HNj3rXe2xG0e2xZzztXCIDMKxssJ/rr1rISuvb85OC/uc1B7tDqbx
8CsVMqWeGT6v36fvIg5pcSdaIs6wGFG4IqWXqaMM7wLVLsKgGPMgQHZqBUpW
srEesyxRECfBTecDesDRKmieGzrwPhbU16V3WBdBr3JEeGE07LPsgB8vmJW7
jR7O5AoPiuFkcaPlOarPnZpf2V73mObowbateppJBXcIiGP4drQd2OdvHTTu
d5jf/mw/A8AoQTzfLQOCR+BEimr3DOXFAunlYgQLqfX3EKB+g5vEARDpNuYb
RCQoXrVGRKsdZ6X4i86GKCL9VPR7ifLbO5UXLuRxkdsLMJtEx4xLSaRmsfkf
imuRsTVxtuSg8Ziwzg29A92VcMnvdWZu1Eqp+MKTfNqB1XCZRLfDT1l3p3/k
soL+Ed1aJkRenDe+wFLMgearjbmrAUostrEvovLoiOSGzMljjHeXpAn7i6YM
EgrWtArtUa/OKTFrbUZhwCHdJJF3Jf1x4ebY2rChAnBcCN/ASG0Z2xCvtQHv
MlSOQTHbO1DT9OO3xhj9At8TlVCiEarXHwil3si7/tSFMvvvwGDiwrfHRpeP
KlRfuiZfZ8mGhjSctOBSlBjOMw9ZZuZRwQaAkieWXRNvnpFcFfmy0p/zwPgR
vECcMoe3BULX1ZY7rQ9PFj+0fbj25dVDDD0aa7ljyGv2SgiMC61aNI+ERv8n
DxRvMLHKCuuqHQQpAZK0hDaIgATYv5nbZEVJfbBANzWbBFtjuRuwpyz4+l11
P/vePjBKxGNVfQjKjPWh1aZqPcv7gyTVLz8JjnahwbJeMpbmlVOg141VzliG
86irxd3/xoAj8/RwtRGKUeMM9nG/Y27dN4q50EgWKwio2G+oc6IYoyw8Rw2u
RmCCVxFmhSEW+u/1ViUvIWhvSp+XiRE6U9kO7mlVGTQUiod2UGFv0v0hqLS8
Ex8Hf1DNCNxXiV5yU7Ckw8J2YvOZHI4GtQGAPS2qk/SprP08bYRGQtKhZiuw
Lx4NV/WbAMMMw9Wsj4Sf6MFwOWsP3smHj6IE2LhxtgRXULrtg6RrLlQwOYHY
735sejpjeAIuLfxzuFKn6I+eDHeX+SFt5kqXeuFk1xnj0NhkrXORZl9vF8bJ
5z8bZho+phJHA36mRD+sc6rlWOgYua75XuKwB2e4QF51W5ZVA/zndMQFMnNr
YUzgbk0R0P0fyDrMtrD+8+MN25VQo5JK/O+LtMUQLqIsj5Uv0bGo6roz9Sh1
AVCALqGl1esSMIQKauBNrw7WhXKu3T68LoxHjQpTHVA96EWyp3n0smLWIdmg
/S78H2z04dVU0D6BgF0mjw4JYiJWkshrEFj+XJfAjs78Gc153PKUFTUmPeFi
/1mjVyi2n4muXjv5VPDrtC0mOeLjP1o77PBh4bdxocYbk/rs96r5LT9NMw0W
68rKz1BBYxbRQ24nPGVH35t1Vyf1c2UfufcKLCRoFnnkEgtMpT7L74FmBgzJ
4nk7mOk+j/QKNZxtk8Afrm7nI385UNY0lmqSo1VJqRZaTm8SeB+WUToGUCHx
Ojn9ABgYRZaWfGKF0WiyJrVq6f6YIxY4fbXo//oykPKzfyKoCky3LC1+BGPK
DmPs846Go2EVLQ0H6vMIo2T8FaJdEsYZ+yI79Ib6/0aFZGTK6JyIiqx3MQBV
tTTh1fBAbk6upo7UNQXAasY4Uf2t8UcArFdAKTpJUWlmTFW6bwIUL/8n4EFz
2WGsnC0Fu0B4TjF3pBnY250E0cjR1jaO4oGG3t3F4Cymvt2sR0t5xs4LhUP/
s2pIN25jcdGEeDICL8mrV7x9TeMhGEp+wRWbFZR6maKXes7ehQef2fi7vWOd
jvBvI9ojv6WMaUwRr5D4MyXCfbLofIvt1j9l2kJ6gbp82PyZ105IWsWfVlAt
7j1iT+cDohwYoO3At0/+tsoa7K4gecEaSj93Sl6d91I44EvOhuSWR4mOWepz
eZFUD/HLQqArj+OdcLo3f1eOQIbMzY+nNCPN/dPuA2OXynXhSDBf6Yxytis9
tLWff79W9+GK1uTCY9QIPkK707wrk3cK0ZZbG+EpcME/2zQRJ3w88ZBEMAJ7
DPWHdQIelp/FLxGbOGD5G1tORbFGhDaULJ4ZCwDN+3VfbiNdCCK99UOqgFUM
xalMsz4cl6mLaSNc1em02yoF1panRSoVC7ko7Iwk0mCvHHqubYT2GgmKsDZ/
vc6vzB4aDR+yyz5jVphcftYL7ykx0oA0t8XykOER5fEajKQaECbH26SSgD+/
Fw1SR5qWmtnLyGkOxMLQ+9xKPuLghEHRCG2IGU7hi5paebFiQ+3U3XXsqZ0j
Kk6MpMnMZaL0GwXvI3hQTPRQP+edUSnYswmZt0oAt8tnIYHnuusBJRnZjhAT
0WooDasfFXUPWuylFrv6A4Ekz6u6y+S9LNbhTyy2ZiTBGCz3ExDaEOUTp6A3
jE4vAzRCKWU/35gyDDB4G+O++QTF0WmAYzL8wC4iLWQWD3HqJhZ6AR6zPHq4
35ZcxUsFNRl8Tb0CRyrtas6eNn0FvO2iRbhq/UkyD0dM2+896Uuz2wf8QKk2
RLI+lIlw4EtGU9xyloY4WD97dohNodszlISBUp77mflRl8SVBk3j2QhY6VyD
kJIB9lRxxYvoo86Bzht8oI3RDkBM1t8Ft0ir2Rq7XO/BV8duCNz416bQSkML
wbM+8UZxU/ufUm4U4aYrlRZr0XPhTacTrnUfseyx66u1IrSZdFeEdlEemD7s
PMOz5elnQ1Jd6SOky2WJigOOvzR7XTH0TFDCxDEkJUrYOU4lUofTdOcJwurj
P7cPb7J7ALYMBTxpInDPNQV/K262I/iUoR9csDvKoQg5d1phD9ja1yY8fjre
O8ioSnkG/eonUG2ytPuPnAMX5lo4XNCWzX/HQTLJ7gToj8gBr5O6XYAbpMG4
wBHrlhvkae/EpbRgPOdTBljQg+dgTGV1Ubqb2tfE4iL+6BLgXYeNflw2wwqq
1I6nk0hTs0eLcc/S4UnE2tKHbNec21A25fDqMqAIbBd7lvNwhV0CtZAx1V24
QT8Etbs9be+whEzzrbB2YWAobiCvMcWWzyXJ7m1grn7j8wUshOOeO2ISkRJ4
0+aUQCH/lnn+tZoKKHlHIPzo2+BTYhLJcZtPzkCYYoMN8LKq15W8eQiAzb6y
oq8o41u/yFUn7icHgcH2B1pEL1AxWL5ebcY5WLLPdScLBWe8PJIfN/+JMgHR
aB3hsYJu6/eBtEMQpo+jqrehCKUJN333mTSUGbhN3B7JFh5U6zCeJjKIloV5
C5BMtgkIUDifnbAMtNnl3eK4824TFpexrUrxTyS5nYjh0ZogC5b/Lscv+p3+
raDZJ50Jl+wlVLUCKw8sLYZVqLCBEVbsATP0wE+6sL0HDTY9qSBREN2sK7Uo
bYysBuDIBc9m0u9c3d2+sEqXZ7ihdvMrVfIolXnoZWpo/nfqH1cHucqoP5j5
VvFDut17Y3rCu7j8QR2wOvjIQBZAkRmWvpNis2YjgFxUwxbnhpCwrT1wyG1/
XfypaLEPbe8TMDsDyhYvWloHnPhOg3w8CnYysTmyUqdKRAynSB/vhi6VrFTt
Ux/159Ci/5x3TOJ0XHJDDWVuR09sqxh0bLKyvIktHxvicORxP7ZWLBBfnfiO
UjrQvbamBXf0ImLk1IBGd7IHPLnyWUQpjDDOQzR6acyxTHXtwRpdKcQG/8GZ
dIx4O5L800qaumVQpUU2yBZnsQOl888gxUIsFTEeujnFIqcX5rQg1x/dlxh6
JhsWNNESR214VdumVCAcRRKjakZ4/pkOdxY6oTOv4Bqkc3sc0k8NPG0W/WS2
2isYaI52YIqcC/TJHMQwywrTO6wBEJZRA2twXmshpf3AcLTHeUsWcp084+os
oWmW6bdLu4H/DSmzpMIKytl3eQwa+QSvYcANUFpYVE5BZZH0zeiX0zvFyK+D
diy4augucIubtM/rr0DU5SJQ4VF281d/s9WfS6eUg+glHIjXXcBFy1S/44hX
CyMiXqaHrb/iy6VhBK8yib951Pi2QMgIZlHY5N4mJN0L8OBc04TIwT+8HQCr
kyYCyN74bj8uJC5hoVRHo4c2S31frRBn1CbYAn7/wHHFm8SA/9yu8xyi6kDe
O3c6TXfj9IWrXDqAe1vtrltuhenK033juo5Uqw5uLmKcA+io5RyBY0AQOXkD
X6RrWz2OMlAu9EAD/LVShPqiFY1nhURm3+BcICAQ2kA8yZD3xh2pDjrmTSEJ
2F7TVx1rq4iGxO8wLDyWaHbtIXR8zCuDkaEwwtPBsbzukc/fPizWEhhuGXlR
jA78e66nW5SHhQPicCfhyipX5o2EvkMJFPyjB29UaecQkPpDflB3psWi8QxL
TNziaZqRig830L+KtYz4DEDmgIr28Dh02uLK4UAZbzsbVH9bteIG/8WZKNBn
4b95QDZ1BTxzR5MSvnfTmFMLhPETOFWxEOpGQ3AD+srTh0VwCoK+phK/xnKc
ykUbm6ImtObtdyAamWTZT7taaxSOMKp9uozZ+DJext0t2QlDSZfikiqSIznd
d7dJ6ipaITOOXCgrm+oZDGgprzVeSxrIZq7GTQNLU+eDkv/0wjzoDR2OxPMF
Hbu2FU/hEHnyTsh9QjhEhi3nYJSb0DbpUdSTwbc43Qq8hPldcDCNJi2bIQwl
6ks+9AQ8yHmN3Q4nCoRcpj7pJrCzex9AlFaDs59EBC5GeeRlUqinA+C5J/h+
tBZkpH6cZYL+8/MDX8qCOMXbGTQniyw0J5RmYBGwU/7xLYFT5REuXc3yBKoO
e2NFh+JKRl/tifa7i2MgwVa4cvC7wPnZt0dIkGfg6TG/IVj8Rc3RKy4Ft9p5
JU6WosI/dx5uH+ei/goJ4WmpU21ZdxTNGKPWbbgRtJ0p3K+cAQBdMgOBGgYR
1YJO5UbpKlBYe3aOn6Zbg8BZFsSafwjMWgjm3XmleqhSchkeY+aJVvqGZm36
H+UJ234N84IzRNqErx4PmWBfVx06SMi06+uW2jdMPFVNbednx8jsenNQrNjq
b0JznIyKwI2xT5qYWOD5T5xIofDdC8wDUXtubLw1IC74/Mg+SozGArred3pH
4boHEdCvjGjL19ktwPb92anixznNwNN0AUoJPcbgoRl2CUjGK6XbN4mukNqG
NcnExByRfDTqC1TYR+lsYSlrgX6ldJDAi/AH+R+hpK+PhAUPra53ie7Rssu0
u7ldW4DjnR7mcm9E1PyiKIvcitSBTyZUhrH/wYkeooJyzaHBd/2qkcBU7xL1
Y9VKguqaWgzXS9ynxBuFUDA0yCH1uCqS42mwkeVjY5Gxvwh16b21bIbAgOdM
R4M6eQB03ZC7SKHwgJ2ywDZJYVTPekREqTcEwYscV1dtf6TFbeNZJTi3pv7Y
+jeXw/myGKBSrxYricJTpppf3JMhqB+rVqhi7YuPM2QDySXq9T8v0bXDWahm
tG7vzDKIPL8G8dZQRmU0PKZ3DV+PV7+X4WacxcW8F1EcjkYKW2j1e016eMZw
urtU244p121LYJTA9gtJL4gG65OpJnx79Ed5ve4BqNyTdpvFXMuO6EBPzHwS
kTOkwPcbELRLGj82GnFDC5EwR6n1OGfAxACoND9ySZsW2+cqXENVpG85mA3X
GZ0RdP0vcN/9VOC5PcZ9Q9AswWs+MDN8EsDvL/Sh2gM+HbY1A4Y0NW/5kyZo
T/jLKe46LKo/1YQPKrsUBat0zmbZcoenWolseytSykwSb2CyLvT+dQuhiJY+
sbjViPR90LW7Zk21pQJjcKQeMNVGuWERAioxm2/HQVKM36fW5nT8L0HvMWdL
Vv03If0BZZi4gLMNcWnX3ztJuQsiDjcOyFydpLvK3jQRKZ0P+5UfCev0InYC
lX1FHndck4NYBUyGBxC1fHNK0444GkAGjXNYvrC0UT1cHFgLZgFQdBq573rD
7jAXO/t1mlh0t9PaXpIrUNnDjomX8mqbkdU2v+wNc2yGdO8V15l2iUoBgPc6
NKa2kur55sJqGsl9vvU+B0diejZ4iOpSHIAwZxJeZmxosUY/jBJ/vO0sCtLE
CYIg0d1BPbDR84OvVAjsGwGJiWGhnTR0lRw0QJUQiJeT33nhPaHRwks1lZAO
QXWwdY62dw277oCF4BUTxDAVnuynNGKD1kII+DTInukpDHillzloJ9GbOWs0
BEkSffKgizCEAD3mc9v4PRCVCQnTpQzYJDpBMwNK9RSk3p9nY0shgN2x4Dcp
CjcMo0nK2ZXuZAys6UML376SaZs/ZhqZ6p6+6W7DSKOc7OgINqrZT98/sCC6
IcFg7xGPnDxGmar98D00jTqW8j3kw4JVLVlS8eaRU+/L6kMVRbbzyVnWR18R
s/tIwzHtA9NGDFnLRch7JOIk5VajVS6rG+/PPt+BflIgoooqDlgtVIrgGn2n
pX3KN3B4NIzhbdyqQMCtXjiteF3BiJOj8rF4+QvTn7zJZFJy2vX4kmDAAP66
6A+YMk8B66mXh4JhSlSIOZcuPXbA6yAEeyKnxt7HnX/kfym9oPvRinnjvV1m
TFAxrKFv7+hO2ibVBUoffA/oJKY4U0Lcourk5Uu8pSORe4n/9hrhHaejNLof
M8qfrQ/uILhyQF8W3/OhDKGLHisOf+it9sAYTtPrYPas6ssNim/i0BOuMFBa
Jj7MePhLvEweHD048DK44A2U64RiSn4jg+ZRGCPUKCzfd6p5npQN8Y7Z+ptj
nUoEDcRON5F/bXyO8C7Gw8koQD4Mp/NQZSX+kXdKZa7oz8JzFQvcbSmloWws
BQHer781EqJYhAbUtlsfh2iqKU56Sentmxae3z5L4sH1wDyma2x8YY86lU8/
mbxFV9Yb0pFn/QnEMEAT5rvkh46UYoaWcGsrfQdf485g5qIww1GYRF5SXYYz
kanr9XpY1GweOOSyV3vNk0dyQn0NxhK0KSMzYL0aXqHxLgUSR+ziduHQd+i0
NY0sN37RZ/t87nGxlCCWcQobzDDIoKytmiaAajqt1AwPP4xKmCv9cawshUrk
tr/pGftu0RnOFuqmAK+pfvghm3skBT2lxKugVFj7nwhdST/p9VoLTKJ4TURU
0abJCIly11+STNbsaTd+NHfQs9E9ya6Upi/Dnls7ZVEn//cbz2kiyFU4RYDj
mR48oa2yv4FrBzS6rmDmCKMN6o5hrUqcbHdhg4CPM6uq+rGQByWA2uIyoDEG
SypUyyURI2e/69IyuCs/+BDHvgfJX6IR7D7RtIAyF9uiniDIvMZ4h1CxCltH
tDWENWoW1YFYHcLr3ohBYBTg1juabRMjZ6Mb2If2uMErNHBR+clpYU+Cqv+s
rv4InKQPHJqkk+weCZw4NGdt4/AOjtnnoV/BmPgWTc+Mdai3CWbb0f7eLOsJ
8bTcCGaGNCcpSR9YoaNoIX9VQGsXZtudVQNY2mWoSbOfEaGFqsT9yubzjBTi
x42OxxH4eCTpb3T8Ngc3T9Q8ZEdzKiyGMEZnDgMVEdwqzbpFJPFN1K1zL7oe
hmVvhvueM7D5kS/1IIRX4/3+YFROecJ/Q9sDuTyq78rqtYENQmRAY5rF+Iob
ilgmhc7lnipvmiFeUTczJlt/iMtYf6YMM4yLyur8vXCGCnEHq/j6LCJSTvG4
DuMpd0reYS13pzKxA645o+NRfBAKmN5BBXSceK/NtymEL2jdfxiDBhroGoHm
xG5unT+pZdsKIh6wexkcbDFcu9q9JXXMU8kOVmCGSJxgm6DdNDUdXJAfevJg
Hkhw82BLWrWa1VcxKTR4vSjnA4aVVWIIqPYgmwZAfuBOWlVg0a3OxdPqOqGo
+gGn8dYLK8zryKHKIvYceSJg1CETLgB5i5E57hyaaAh+JKrud0sp8xfZBnQh
XXmJr43uvotZ8t8sHSuTXHcv9AzzbnDgtNBtKRI+VmEaCElJloJ7M6bIADOB
qWCVRJ/37UfI75iZv1ASBr6iTQKjKrbogg5+SoFAyWvQNjw0Yf1X3eRwfR5Q
jWpSeMMT6DkL2XZgLQxkxKFTn8xPY7IpnP5hcy4ew++6vn1WDtlOSX+IUW8r
XgYjgXt98pDXdw5AGe0RL4KJ8L9C2xZFXTu1VlYv+neL/KzpFzO5B+dIjn4L
GqSZptZjd2tLW9RSv/KhrwrDn6JFZE1k2VlF7/JEuip/3up43I/k6HqyYmOf
YmR5pd49dDDBIy0dOlbJDeE5i7I9s0dZ+UaSwxGOO6CUO/7Rqw+BTLuOLmeX
zh1bkU79iDBcFNavuqFkmvnHC7ozas7nVa4s3dDbXAlxfRrzeVdYqzk0EGzk
JGEgAREVV7vIG+vBRGkOgDgSPhEmgd23gQ5oAZgKT0HvczLsDRo4KwmX1JbP
bBF5phTzMzCNTS2QYZcwqO/VguB082+G7L2pBNmiD+noad050cfohDmIHmOg
gQHu+uPzvD7tIAolv8YU9kwOB9OjH4AaooXrVAz4N/tXSsU5bBepvU0KBQkb
3a3lyQeprHcUW1hNNRLy0Ke1Vr0ai5NTeGzKruoA5tiLGAAfneBVwekXgK6j
81x0NHsrJjw0WKLcDJ2dN13Aj8XP8Pd9tP2UNEbLj/ZZiTmlEDJ5bMXxYxBP
rxi2Ey+Fg/YTSST5si5LiIAmME3kO9zUw5vIasajo+Rzthf7fXlYIsR272yu
Ge8e+5oOQKw/sML1TcqQj0ReX6xrGgo/Orp4Znjay8TPU3ehskDy6KgOANB4
+P72Sqb0Cs8/DZtqCsXhVF/XCjdwuGEpxBTLqz7HoZf0lNVL0EOFVJAYf1FW
MKB25c9jcWsldhK4Z6ixilCHnOYlQOSC95Geg8r2Lg9N4HJwUcEVDAeuVd/g
Zwo4mU5MiNuEqIE2Ja4pJJQWwwu2LnbmrQ1NcozUfTQe8Y1nUvsgzLEUK0Qa
AnzLGU67yz9RmcnVdT/KOwbildDRgqgjdp8/My5RlC2wL8/u6VPuYVAkvnnC
QkQ8lVM+13zZ6zfC2ViM4L7Pu+F3ENqi97v50RARMsyVMZPVzaKmOZgOFJTe
Rxmbo2113oOyC67Xze7zZOgF0UV2pcmx4Nki5zh3af+74LIBAeMK0nEjL1Cl
KHav48dY09IyvF/mlLKKx3wtozxKchpG9qDM6fnj49cU0811JfGiX/XCmXO8
T0SbAueBYFleP3Picbepb5RJdInsuEj6mb9/U009YA1VhkysAODHkCMrR9fM
SAUOZ5zWgzqWlcWrKpLW02IbsOO3IBVJI4imUAgFQqEw/PfAg1YvA2asabKT
e4rRr33Ivnz0QXZaF80Y5UPPyaynljLXHV4UrNxxHOldXXOKZw1BSz2JRWSn
0ijDTIopAo4nK09/CC3afbhwqrDX7bYF8y/ZCRh+Jb+0p/BHN/baNw4GKHvT
1ISnDJ7T8Ery+pohvg2aXEwGoNqdXnWrNuIqzZnQhRR2d0ajTU6mFBHB52W0
EIiGQ8/m6Jn+adHAGujkwbxJL2eV3Oy7r3L8kWM4fYx0YsoThpS6k52wgD6a
ZAaWdVRbsbdu8EiS2bpp1bMSTcMMd1aTlRDnyh/rrle36xiGWh9+GJnjFsZC
kcUjClc+mJ7nRSpi8hewbipI49MVdyVoj/YrjmAgMY2T+QYIrqBA6jMGxb2P
BNnQIax4DGhwSkXUZV6miLxDRE4O+55qTZ3N4kcHvadlSALL+cZfkZH0WidZ
kTwhIVCKhCaqDZfKRHag/wQmtGAskUVXOanwKw1UqKKagLtaWxSAOVnd9Ehu
6T0SIa5vnY8AfRCPIyZpkRJmsZOiyELO/ltIHX9Xej6MEr0/NCCTo2ugJA3s
PoN1vDUTFpkDlQjbNQa2pVrhUKDe/POg5n3gYvzBXWnSTMgzCYEVVZ5XaDk2
m0r325PkWB+nenkLWbxQ+Oe6QeuE1jBK8JNPvjHF5PvZ0Pfm/cjf4/+qIipG
auClURBPYKWixnBrr/aLneY4Kw2yt0+PxC7WbxBHjKJ3Lou+oDYYF3iWGGMJ
gnLdxo6/kvPD5S9Eu31IFb8/IOAc6thwCydarSzjfvZkHY0fo5BlA1Wan6Kq
0rBIlsSBEbmnw4PGvn72Oskb6RCuTN/MLZIQ7dgOU82Rvjj4R2c8LXD0ZvNf
23uHO/EzfsYJC0fyRPwvpzuMQZKqd+S6FyTuW//5tMuLk3RqWuIm4mo65scY
PnnzAbQQZ1p5JagLlBXJhdzAdBbTQcNr/gzOMEktNUcgn9O6VCWZ+AWgnnoZ
3K3NgUga3KGZdWC70+M+3g/PesyDPQYBzkCU8jUeNrGPwU115mmb6+SzhXkO
G2Nv+HQpSM0Ofz07ik1VdPlLfpnejq2vNvwT82gCEeytaNskSHNzaCPVQL/x
NNJ9C6rm6O9+sI/L520okEQKbUsHYTg0k3vMJlWFsRADXqkLDSSVFPm+jrvb
zmRCSvxIMcdGAYF4Q2eHkD93QKQQ9raCVkEWlMrbFefOYxNc92ShN41itZWs
nZGHDGd5DL0JJSepyIOqy2Wa/PL9q5qv1TezGYlmXG6rGSdke0nKT/BUm2uJ
fpVIRxb129jVMYSfABf98TkxdGviI8kMRUM2/OdOudd8Scl2rRCIkNEBXrG/
AZMhKhx+mqWJx23cV4z4tieWRrSc94JC7bGI9P6Ni2teYklCVbkAi0kExYXS
U/Mq5U/4DGHNtcYTPUYJeWdN0aYsCLiKRKWvzY3AVp+TdRzatb5JyWNm64al
OAn60YhKQKK1K+sB0KPy/NFwRBpmOn2dq6GHnRfL6ACqI/UDX9zb+U2drYfu
EVAoVZpL34uhzN0DNffDT7aLFby/w+ESvKoC83U6mKJzouwohaweEeO8NJZE
qTYeT/fGa284FWomi+nETnvbCQz0KjOpL9zzzn5dT7YE/RrpAvGl7qW+UdF1
YCh8Sajp/UNUPhcuaz6Zy2QWVo7rw5YaCVVsH1iEUvVeFcPE/0kvWNZUmzf3
G8RqlCnCG5EE7ynhFXLeqs0VNZzuW3rzhGYWq2dSjv5pRvtQZ+Lu9oWAfFoe
mn/ZYweQa2aohLtDeZq68bgau5FnaOHGVUMl1NFRnMtI0dqsP/M1D4vkZ0I0
2mFIvAvjlav3FEoSGOvdXpGHzOuq7VMpNH8HDwsMI1bhJFEBXrDCdYJZIk2O
gQ4X+YBM7Mkh89TR8ZuJcBRgRPWD8+6sb+5H7KiuUun0z9ONoFrfR7MVv0uZ
Gxmr6ELobxbc28JIERo4dImue8NGEE4qZPI0gAIuXFYmDK4rq6stGBlenK0q
lnUjw6qoJiu4kZhIHlOlGIJATjRIcNIHlUe37bBJYcCGcEYTyDbzW5xkIk9d
7EbJTOjMuqMt+POoZZWgkoZcYObn8uY6QIFRvwboX0eq/QuoBsUaD0FTj4Au
mxO74S4Y25bPVf61/Gp5fcPvdTZ5EdViW1Pgv8yVQQvtZ/Nkb7xgN8jhMQ8G
3wdd2UHw3d9wq21LmZmJtLKZM7UxSynNqyH76bOELmVBy+LZibOYqVezNWHe
zys22adczpbcU9+8PzpvwFL9Yl1AA00MFBeHdhLWlkOj5EHY/b9AE5qCh9Un
fUxmatVNPvC9PflG15DhizPK5W8NQH4CV3+5e9nRybrjDoxFuGnLcc/cNUCl
XS9YSneClnlDJGCmZq+oIBCJPX1hLuLGbae6jAmDmf9GvvjpZHDusCXx+ltb
kgYp+ppdvBg5+2vBDk1to8gME/NDlGm8k887RtbSbUyLxE8JD73COZqxyCsk
yQoUODz//HLWUOSBJvEXzUr9SKAFD1W3hY1EN84e+MXXkWDtIi7+MnXR/N2E
g4zAsmSr+465/9Ttje9P8po44IZ74Xt4HU+nXdtjSKKJcaRABJPM+FHDjlKE
TTBIdcWynEiw7GihXFJrbIwlr/I3JPoZrrie54Qs7jWfSuV91aw98FAVn5Wy
xyU2KREvuJT14jq9s0REeYBGxcgvAoda1qObYYzUeyOXzkZFxuXvWAd7bUND
7KuPKnUI2Ql3xOSSeBNU9OYIsDIDF4n+IDbnMlQ+tuI5SQxlxs9zv1EtVi/N
7c8mpDIuQnXUaVkLN8A6PAPWPQ0UJBv6D2lZ+3Uzav4g4xIppDQx4ghOwKMW
Eedptx0pnNciCGPF4EY2tnpi4qFRA2oZHfRu91gfVupmr3bqajL+0DBX4fkS
J2BdkY0sW5VvQnjFZJuRnyotXKtXs/WCJISHBlHZXajo1pguPxaL1wNU2rCE
PE5Obf4B1xJWClAH6zy5W0ozty7c8pzFWI1C+n53U3Cp2dOPrsZek1J5UmoL
6cMaETnvm/7uR70HyYTmf2PdcKvbuG+p6VEhDY4DVA0bWLIYkse3s4ZfBaa9
Rg+lVWUJoXD/bpFZPR9edllu66la3SmmnsOzF68u+F/qANzCCZBy0Sb0bscq
wRZsv7yUEx9EltKqUdqAxV2LvJO4mAZO7hpzOQMXsvps8jIAOu2sm/SSItLA
NDhrRTVBfUU3Ks0s2kqBwj67HbDg06SoXmmr8NjuegNB7ILEkF/ijc0I+Tik
G1zY0AC/QDZn93KSp4oVfZBXUarEswwdJGzlubHiiX5e6eKHmwVo2gVCzEsw
G3h+IJ4TNdeh8MPIJle97t+uweUSkBwe+lwdhyIwQMhqqNXxfs2IxelYJvMi
blFvloEVUltr8ZykewqK9LPym0fbk4SXrHqfok27Krj/CG566JUaAaVAnlkU
8elvACL6M69FzvUAig9Uey+AnZgWdQ1nnBXfH6EtplFb5Xyu2x/1JkRkzU51
aIVBuinqWj1Zg//tmNUGVWvddtV10QBttDxI6ymKJy6Lvp2bc2iwQNoO14MV
wPXY0Z/6SN9Ca+5fFFv2RQ18/sP3u+BEePBjPcaw5zlFs60b3LkB0hTE5moz
kXQxz+l2rQMMFLNKCPoDfDtpe8kOFMezSsKeHDNdwSfF/89EDZT8gl2+CciD
txnipI0jedIzWat57Za7FWF4oIOe55JkKs+xX1yt6xLX7U05Fe39AGe9NlPp
gUh5VPKna4Zgz3oThR/9Bos2xSJixDnIPLfKO6wnWEU2bfVaHb0mIeIE92QN
l1ZxsmHw3dzz+JXslBhUgobhLifCr9u4NyD7JFQBTKoue+x9fVDnSp10cSK1
T0dUENXJsbO5PI35ep+6c/mQvS0fEc8xpNLRVVMYLMz+jsaPhDP60J4C2jUw
JPrWB8XbhSowmsmj9fFNHB0TVqEDaXEprszfUJTCsSG4JTcMsQiIB5pfrnjo
XL3dafOFreU7l8ahNc+898hD2eCiLcyKQ26jwDE7Th9aJCfCb0F7GqAOydlS
iKJJBgS0XO+9tBKs/Jk/s/XutVwOPZEgZYXc1729xjmXqHzC635jsWMtgnO8
sRmbVDdqtp/wMHPxt1/Tn5GsjeC62N/ymTP9LP2nw/hdIpQc5xX+eAjG0glD
zk7vA8fJn31mbIVeRtd/A8i2zKFknchAxkhGSgRuMujckd5l0fMOGERH33jm
/OUIom/5NxfS1UjQ9EhcSGh5k84xPvfqAK5pCMAd/qM04Jd+yROlrt6YCnj6
DOupR8ZkdpuYd1CFSukliQwIZJWtEfLbI4mo/Bx8cQKh3rVGmtuF2vhrDIl2
lh2vxrLEh3tgfx0GbzOQMJybPLmxhNYJdsa56WGK30+DFI+xrXDpAmo5HEwV
9H/rJpmwluwLOPtCIUQKH+j8LPwx9Zop1ZUZGA83PVueRw6FjUR0w76aSN0D
ZF2GfwnlVIFTkctMadLbRIpRNw04mN5F4yuliwi5Ynk8DK+6TCRLdlJYsuni
yi92v/1D6c2vOAAyPHJBhzxOmcwC3zu0n3bIO4gcsDBK9SoygmzgbOZ60uDO
Nu+I37fZ1ggO8ce39Qqji2iilV5kJuBpudhFS1TEMzMwoCSq8D36IHR8dmwQ
f23UybKPjMD39qZ15IU4X3YZCSOkJE+92wlKrzzJqvqBoJm9lAKJzsaMPXt3
cAPMxXry2B7dhM3G6ihhhbiyHhsZk/B6v5v8vjA+TZtOxF+LSrMRWx6qQNpd
q4yBu5igdrx7Avn5M6dGa+M/ZzkWmDAAthYDIV7FOy7SBwPP3m6umKPkVB2W
+O/klYCHDZ9F53AalnQiK6trQbZaiG7ErdSU+SmDQ1gceYD8fFoJnZqafXp6
b2ZE4Jast0O8YRLii6BZlHeDWY4zBei/o6DibCVXVhyaavElXSXneNyObuG4
8S3WoT/EwpqijGPkpxXsNKTqJh9si7sClZOyrvqsLPzYrxxM2p8WmghSLX6Q
leGvlrGyVi4RChBTClt0govsBx5MKWSGYlhoHPbnbH5klJNG++SIXrIKle/9
qoBfs55j0dZoFh/JvOwDCxtw4qaxzVLz6ADEnlC3JYqnGTdfXm+WSo9gJizL
W3iwGvIs6QIJPV1sFYQ33NPFkLhNxvSb136C5hngJgV6kz70ErPiDS38KL/B
xZUEa8gkF7K0ySCQ/acVPTgTbAq8y/jdyG3plViBeLyty1HsGiJV2FjJ8lPp
D7v/gNI1bbe7MiqoHdqzdfxiUarQj/B7qguFxWBb+W4E1XbJNWKHWLy7U3ZG
vEKjCCboWHOPOXqpGdrawELP6//TwJrC/+Xc+I9N0hwy440ZXe6T3vi584xL
VuZEhAC1QPPpEmVE7fS3KxXEwMHwD6cboUQWCa9AxA4a73Gk3BICaqmM7/fD
d0RB4Xjt/BSQNJmkLKjQu9yepyDQ4EnmI4O1kWR7Tk6fR17ScsrKdyuAIvju
JeIk0XMQcBVtflfQPgAeN4VQYiWfwvM0bOHSY2/Sf4MPEK1fHOb6Y4fX51M/
iwZl6rBcViaz27ZfntprmgdqEjSN1AmKYGU908UOqjl0mSI25tHUtuwqsjly
qP3Ui8eKPJ6EJmZ9TBB4QXlM2Ljs6UiH+BIQpRXqr8SbLE57v8/kWmMLG1JK
qHR1wAaAflKK+vtLYGfo8VweJVlAwf9+Svr92iUrUjacK34ab5fXRLtZB4c6
6lMNyP3Bol2pviXzxu290ojlUeIv3m4QDi/+8fdnO/IkmheP9s6pnWD6D5k6
qoJ8Cjyb+4c0hrFJ6l8lln+AWqWGRPzzHA6gt1qmtPIHRn8Tuy0yqRmAIXTY
2JTMUhFRo5TUxkm2klvGj28PfCAjcDedEremjilWsONenWB+sg2/rFC+32Lc
9o+MkiZu/xrVBxtTgOD1m0Bn7m01APMf5RyUKxa3Xu1MtzvLj2g79fEG6PBC
agQfw2KLvP/2ziFSdEIeVXxKwyTWad+7yuQukoqB2lM0qy8i6+enflly+tnv
khsalpbc2Gck8srY2xOoZZyYU2bTi6LYIfd755GYLlbLlRIYZldnN4PeTcNK
FJnjVBXtbZHA8LPYWAdulCmhr2/13IHQf3+JTuNH9RToPjBKubdhLcCYk03C
ZzAb/2VxG1sPvIUirL5Jw/czM2A2lqj7zDgepiEVJ9jym+0GaPRs2vjhVTmZ
s0MypmnQ/rG4ZgMe603t2FVEz4R/Ifu3Enjlpf26Jr8TXH1NxGOh2azmWtWH
D3xVeVbhZhtnZBqkNE0gqiT6kks19ZrK3n9zpkbDqKgGQ/34vi+ClEDGafgh
qoakF2sSAe31fMqiSDMXnlVi7xqOKjbrJHqyubfXw6C0zqQUSlBuBj1G3en7
Xpx8bqC59gmsWZCwCpfBwnoBL88fVakFjzWT/G3nrEdk9GOJHtVz2hYn2i+t
GmCc5yDNwazlmfXQBZvPKxvLjJyAgqrORSXmo6sdVXVZfK4BRSi9KfrSHWle
TUTIXEhvN1CdlK87laa+j4+l7oS6qhpcLLXh3qWXaDPLdsy2usSwCxvy1WW5
jtRA7mjrJmCBd0LZpAfMkcs1JKgT5tIbxypqbM+bH/WahoX+hKCkHfjquA8E
VnZQDGTjbpB7xkohRm4DbV/suMhz4S1ElU4Cm47+o16CokAjKTe4Vw2I1fTY
VoG0Cx6GvtDe4xYbMMK9Oo0mhEzBiVTmTuTwt8tm33WyTB2zGywULmfMVsyS
d6yjyaT17fugWsB8VVr0zA4nfmnnRwE8bFzLfqcWCGyHjEhsZTmowc6UQC1E
0uU5O1QOqc1uJ5+R6CwO7HWfU4PDmo2G7dDiq0D+h4MEYZjrXFAUMCrYyVBy
u2Kezwv5jIRB9mZRjqTe/u6Gn3TfHRl1hpsIiOMyYhxSvYoT1WTslj1BBq9W
9StO3/P9Jipx0QpswdksLi7OU/iAZthDS3hv8FFIa7d3AmZChePonkWA4nwW
s5FGh3JSv9T+uSBpsWPYqlItF8DeY6ZHcBaMG573I7HYRiZTfSdbbNNMg9NB
AOf89vh2k7tvlNDhvY2WuG+SEnBqFy/uJpcIeGVb0myp9pbrb/Z6nc2LkO4E
Rt3dyeFTjNvIczyUDRnwjQnzJ+RQH8wnOwvOQYC2Pq5Pr2VWrrgTTPSPFFgD
8uGtTaVtHVX/6IVocVH9KPLcNOabRJZnIk4UodSc/9p5JwvEILwzEuHvSawZ
+PSOLNQTtlx+fasXDaoN8HQbUC6SMJLeGgbVYjHySX9jc4gtEep7Qu7oibtZ
v2Kn+VwnxYyAasXqtSDcDoaq4FIXZkJTCIBfiZxcpCywFGb21ku3mun8qriP
KyoTTGmCXbw/HT594XsEsXaJpRegpmEA2AelQSFfIFXTfaz5Ty+f6+I44EWW
TTSiXWXs2BfoxiaLSxgdY44VZ5EU7W9GOXzF8BytPMawvxWV6+JWIVqEswSI
B0Qq6sRR2IHekbR7W6CmHqjT1krXSYOtGomXwQAeLwpO9eKtteo443auORQD
mi2hbsZTJ9vSrcfcH21rUexIVGHiVwjfhXuA2pSv60/mOXJQ8GJCp3el3hsv
kTJbJ65+3vtyl4IXQMLNxpxDJXBWQfpqdKiJuOnhoBjhJJm9d3vXqjvq+uMR
NS0KBQQQR6ejZ5DpO4HHcxXaqLzMbXFAQvRtM/J87fKtZXyz/YQU+Gh8JuXV
hZTkQXwa/74fCWk2MfsqHyjFaIq+r+9KIwLTXQ2mvjAkgU9bcJIEMaRmkW1A
oDa1Mf3QjVBOWpMMEW58dhXqCLgzxiKP3Nk12/sQmBMKVhg7MjdUBy3R3wZg
HUs1zOG5V3/TTqQxBs4NtkC1bESK+DMlujb3JVTqhLAp+9n6OFSFaPvvmodP
cIrD8BzNa0+1adF8Ip9vDIgkxJn1HOWIygWor6LLC3XjaMjTYKMVuwrC2kto
FaIwZHr3Mg2zG29AYOrIuKxH0EgiCt3sZZw6QTgn5FwBWKCWarqDFzmX7f1+
iJ+ti1hQve2N4iXa4sV6jxY34sNuxE4nHTjOlhme4P6Ob2+QktnmZzgJF3RR
uebAP0q+sZJkqP1BQmTcWWeaH60iBsxmMafA9EHqZIyM+5xntvEmKgCISZL5
SG2rncI/bH9cWMqf/Bs0l+qFjOn9x0v3MuhG/24/9/8Q96/3LK3ANiAK5Yct
SsxI03zc/h6/o5zqSoSu7+SHVJjMGS/yaNIumiBz80MCR7PUFb44wSh72nOo
zv94PwIu+GCSkG6VzibhKMec/kpXvfhPPnAQRMNd7Snd6Dj1n2vkzRjqHceW
WJORDu0gTxvbDVyXWCTJk/94S4nMJZSR28bqyda9QZH8zQyqfrfYu01hJM+I
XIGVvrWPK4wUZgH1xV+bAIU4cMIsrid+P2v25Kgu9oORMJ0TPnbWWWora4fO
eAbMrTDkW4xklh46NymXPWKPIVDXc8pVVS+6kQnxAflKpA07JQNHNkpcYxfQ
GBtDRafkBzusrQgjIumO+cFwbQd2XUSjPf1e5TxH1nKWYoQ4gHmy4mbW52bh
Bf9rvd8CB0majyDq3ipwne5UTZjkCabahl5XT7qHs534s0lbSDv5sKEL5JQl
ea11doJhpDNfsLQAPPN9odbr5r3fPoEDYek+ksGZ+nvHoLxdNcJHtESOGTnO
8kOw8HYraZx+0bCA8PGmas5cGU06aYLoZAmU7HpMVW9b0VInvcAPYIHNiVsC
X/ohmbjlrU9SCFda3PtEGsrtXP33OuhVL//BBzpISQpoAHMQDHeywnEcaTXT
F9/BHW0mQXct0Pdxpn2sILZvApV4zMwZPKleGiCgaecGEg30/veQnFAcBSLO
yk9QWRbtvrvwG0gZmfYY71B6XWVroVLtqXSlW1bMXY2psCBs2gcxzqiCOY2L
9QgkogZMR2GG7foz4F2lSrXEGUg5TmgLNJtO/4qXEduauIJVE252MgIQMnaX
uz8Kl5FJoNAIJbBM0ITh8vZtu2yWO1mfQbh4BcXYkZYrqJK6eu5Gc1pSioFB
LcGUj+kwL7nwHsDdRFeZZ4ZBtuaNgyGx9B/8YSFDEGO/eK0EFHfV4N5mvk2i
/MOrKDORHh0HotDlA5kcrpvwXA/YY4LDHY+svW9AuQxykNqERaBS1OD9C+qY
tnxqU40fA3CSGkuWga6Xgd8ohBmf7ssYNaOE8VjX7FSXXxa5PQYHeB5gAho0
XCIBIjvFNsL1a7Pkv7bHywU6giPDggNxvVdO1cnRMs9e4sqg82lroy21u+bE
SEyB/KRHTCMpfT1tTmA6NptOHFPmOJlyZjerLWefBD36Lmk4XXU0VHakVw7F
YAEEIFKcXW1ulWQlAob3i0mGkp0ancFIfRdN4T85Y3y8ZZrj11qDIlP8gYai
yAyPCIAk26J6NugFs2aPO9qQBEKoDyom3f7NuOkIswAxTlBYizUK4DwSJPKU
NbjDdhB6bFpK9J6Ks2iD2zzqv+6/+TZdQa0E8YLA9W1SJpbkOkDJAo/CPxDU
CF/ZOMv0r2Av8mU6gxID29XP5jZe7iX09AyeMJrA+5HqxMtW9fIxMJ6a+Lqh
oiBLyKLwKhohXaLy2b29EPXSCcbOkKkq0n8ALzUSyns/ixfFmtC/a3xKb+Lo
9u3aM1V3IBepVDeROz6BhqYyD0k7ceP+fRVqova3lW5IU9vaEkdVQKrMNNDI
i0zF4gygpvWQfRgyj5J0GC0UadCP19tOglqjskaBB7lOlSyZij1N0HhI8C60
Rez4GHtf+HoNPCqFRMPGFdfHnyBMtRAzRjlmZ2+WEP43Acfp8HNzcX6wxxet
TkH+cXkZdlbVxQ3p0YtDtwHqnUEEf1nonRFpAglFo8F8ZnFfCYIrAOFwwUy4
tZF9N20Sne2NE4Se7uD8qP+fbpajXb6AVY2FNl4875I8ABgRKaE7bKYyRyMn
wBWf/EUI2x4acoDKQCS5aF4haJf7DX4UVqKDMbOlhHvebiCS2IzHZkjUhXft
U6YwxPJFydfpWFBh/RgRLn9BDzNb8FdTiWNdczXrPup2HURulka+YRaFOo+H
Y7w/88t+Rtu7d75moZ/730VwqQkQh4nuropXmfpn/i8YClDaBUGkjTQN4v1g
M26rZ5nfgYAJ99AG0sUnflzS/ZhpBQuwufO1GvOyBec83ts/6DHyKbuKiu9X
NVX2BDF3FY0HCdsu9cJgqwbCNKGCn9vISqhku87YUVj80PFh7pzOlco3T7vN
lOaZqyJLUi86qss4gGygPphBVcDWwNn9AmutyTUEDH9jKbLG1VYidDSxNLz2
n8nbBICiDBPQPDVl5E5X9kxpnbh+DevFXL3yXNfCcTNjMfvelIMmylP4FWcB
+txecrEIRAbbEwyt3aptIpiZi6L9HCYGuuPkVGflSz2gbvX4sL8k9njp1PB3
RUvIXqzPVuYgiBlnI/6HmTRm1BWmIhSGfKdYYsdVr9s/QzDEqgJYUpEksJ5n
H2RYcAe6TZwbVACXFK+33nk1MHHhf7RWgqxRNcR4mYCuVtG4I/p+y0LxkmNC
xA3NpPBnfkawNXvbb4DXpVdoCzX+VqiHYMqiNNteQQhPfOl/4kiEvcUFrBBt
XIc/2zG1/Ynj9L72f2c1kcMBwNnSATbLdFO+CU2bKtkZbl5I32i13emmb581
KWmUEgH12eR5pOx7TDRGWan0z3PsuWStF/3HuDfJrjLMTONiWpE+JYcr4h/G
666tGHV+3gaKK5BnksLY1xlURiZdEWjLAynWnBbJ5U23Pzi/wHnrWYQB9sZd
G3QV9/16NcNqvNBNeE6u/8XZ97LDjiO3tNM9qvfwLFB2BHL0RU+COZ9l5ewl
tA57nS9UjoI1i3B86D8ABpRntZkNrZ8wHQuAl1mOvjnsIsmNv9NU8j1Scg6s
6lSm1uj5SN0ZR7DyiodiMj1n0htyTsJ8LBGEfo4KCoCV/+nMylaU8bpfHlNX
Ukx+0k2FqPb2EOcly6ZlkZf5CjkAw+o3DOTGAY2vKl5gErr086wn/a0JUdBQ
JiHsPKsUb2vrpZk8bNQAkLwprCc6t6WHdBj1M60cBd1FNvIigiR3SNS2rdE+
b+cdeWCPDSa3f/syRMOWIFBLG0frNwn840nmcWMnxwicKNGz1v2yB0EkQJmO
+pDpzHZhl6rwOcUs+D3DQSkw4DkNY7ktDaourf9ztJVLn1UQYSRMcC/mhQw1
qbYRYMnmg0EBX7BAlVnn1ww1SpsnaVYe04Wr0W71Y1E2h+xcrSL62OtP20E2
HMlt2xIkJ3vQYIQds9OsM70F1gj/5fykV28oM95KDRDSJKoGV2/eyboCZIIi
MIcfOEVdvLRZ+ufpPJakG3vhbW7RKIHSJCeLIkYAO1pSTNrZsVCUxc1F0hQb
ddjHCRR5VMmUDb8ZSqnQVxVyYoTygppe/p2aIsjZToKYxsdWk//ULJZnvPIF
t5y/YUJy86+oAykMRYGTJ0+IK1wYhxWMbj0eg/w3TLJsBqe1j0lhNnh7trwa
2pnXDMmVWiqZ7AbkY87aW9RatMySdT+XesZCdiBy0zCvy2xyxTMQuRqCaVNR
+FtcDUUspS7KdGgHjvLtG3EJZqh855xqKzAwIhsRr296MeSsHoB6zq+hmu/E
ZEa4W/kmSWJ4wj93+NYv7j3UFE2rhcMq6t2PeaeAbpbCn+YM3pFDby0kRwpb
F9o4QESSboNDkGYMBGd7cvGKLrDy0GeGNdluGlN6Sn7M4V54cbQXlzYwU/t7
+q8gcRrA3bLGoMi4LW4EW4lxqt+8Qecb/s05l3judTGcCzhO20GWtw+3OppX
j+g+gr+ROI6tLwrVDpv0dnEZyqCiv42h/83Py3YTkVEiIdB+YPVW00H/7XkP
aAsSU83GspSWOKhxffsgKT6U+SpWj8Qgde0Y2uB/krsFdC7+LK4pPBuaR1BD
iSB7gws5kc84NlKQzw4k78U1gIYSsAFhgHrqNsTmSlBdwZ79xnHztuaYcUOM
6zdY6pFrXiZIZq++JKgo00XwtIsjaukpPrEDKy/TgWXAmbNkk1vowdru7Ety
JjXgY4o8+JEWb8WTqBx9iMR5IjrbYjElujQ1nw54RupnK2eRMxl6pukpsGoe
xkuIu7yGu4wyIfQ0HWtHe0BUr9Cj7fEPgq8nLgwKZJds1isfjC4Fd2ntAOGZ
2cvyekzgRLO6LRAYAK2cE8Mwbw/PFriK+o/NDVOKKrkhDPSeKrtVwMHjdG9e
jOW8t8UKvYqFo6iZfLvp7/in2X412mXbu5CcZh7MHCDIfJT8bxL+tESW3Le9
S15txnjoakCTCtgQaeuFp5pIWBdNQI6g2wpwMnzl5EFaD/wbyr3gzfhEyB+S
2LbHncN+mPa21rTW1vW5i229M9xEjLkNAWrXthEQkYJc1QFDLml5dFJu3Uyt
gv5k0BMLVB94pTs0MpkPmbuB5B0BL3aa4wmVEL1o9++pQPVKxYOlg05CCb2P
Bntjzri2w9A/wsiyy8e7amA08VMIhkcD/80gf1pLwqF/cfmoryr2tYuAFmVm
r513tHmnB/GouwlEqANzBeHNjwW2oKi5KnUBvhHmZAQIoEhKTtCBsbXoGNKv
bG/83gIOGqCQ051iLg/IvlGWvGFU9Q1an0O1bZjRspvzpYIVZEAYDfjd4VCa
OKln5MXYkBiHRcpl4z0G8gHHhvb4mwJumKPwgokrsqg4etqDQejD0CHm9rF3
TB4uRYQQP8nr3VSNrFypORKuUMt4HAj91IDrmlGL+m3LP8Uo6hzYHUGLsWdO
Nt+FFTvqcaUPV4R2j4dsW1Ni3BgyqfthdwTPTW5C6cdQrMqZHaVwnu2H89rg
t8WqTpPBETbUY+MxpmtPs87W1xeGNtRUVQCT6BbvRlQBo1Vt/nx1fhCr6s8M
46k6qiY323/+Lfg/wijda+Nw2RK3ubpBpIw5KjeBE6Zm7oesKP8l4bVAYyOy
YZeofaVGpg3h0QhVAM+IepxFDRu/AwacB0iqWZlI/XTJA72RxzJJYCfhGz5o
zMQtbUupZXHxxiPe67s33KdVk5d4iHflymq1tv276Ztp72T70ir/jF98vxF6
uwjLwz9aisciTT8CSNQkUDZDd3nL6azAX8mN5UZVtAr/0ANG1cPMQ6MfO60i
ymoZ3bQzJLzIkqOe7ZrRCnpbrObBeuNcsobwHMRfiUfscqt4jJM76wpzRqBL
OCtcqp1G+pD5qV8lsw3iwNtx6XWoCOYPHhCH/RkB5OESHR4WFjD0V8XWp8BB
p8PMh15fufTCv4EKf+PMk42tPHShh6Z/LeQK8m1LWUolJ9guMJVlO3FssVBY
EZ2UTZxTcrB4n4YtnaMI50YV9tlbBgrLbJRxanznmvKNt9hghPrgZRVCs8R/
3oFSQSUCxQkRJ15TuALFI+5b2GnXdNM18lnF6NKIzh6qnnradvIQ45Z09lm5
w0BF6W7F1e/Tnyss9dZpR+geMqwemZCAlDszs6o4Ba90f2p0b/2B63szrkkZ
N60Y98LRqPh+sQAkINaEd2ppacVx+9LpFJA+HjXIu/l0UoJQvWaNY+UhMtVy
lVhyw1DdHabD9CvRLC4Rr3rb2sHN92wUGDRgadnVFcNE4egOM0vQtE3PFFOC
XmFW7net0+pLXaLi3SSwP+KXAAM0bDp0JY7UViXQ9Qz1gOWBpJ5yuhE2g098
tH7nBGilPiNwfhDT4El7a5WZRdgYiaYZzSzWtgJUNIznOGV6QVwPRlQskwyV
dULqKPX7NFANaC9UP8PtwD0SJaWUjrCipOuRtvwwsxyNrofzFSuZh/7CzToG
hgklpZPGnXBm6s0CaTMQ6pvKY0G5ECe+kvrFci6gpUd6N8gQtQjKKwC95Maj
0e/gp4sKR+OollZmnIoJ3dZfrvdV82MsGMh44YbnGdHZOpB93xYbgxy+bLIz
bEgjgsnYg5CB4g/IE+vd0BcrABNvu2XqAxLyKuz9HS4V6D1lFZly9Yghy8R9
tiJZDJWwyVnyPx/t0tymKfmO55PEAPgwVIwdc/30D2n/nq2g76ZPRzkuRAmH
Ljcbx0/leXxqvoQkgI776yeWwRUMsnJ0hkTkJnuTLUCpekZjOjgV0Lpj+DCZ
ygcX1QIySWA33HcBnGxP67HGWyMIVLUCETkOP4qQbLSK9whLpXfFbhr1S30b
BxmX4VVR9kVpimm0JXY05yF4TyIojE9etOAvOxzMzlMqSGvldpcMGlyHPqQD
ZRLrjcVDxRKHUuSbw7/dSz2bB44U0491SdzRhSqklKSIOxoZkvWU9642snEx
aaQpnZHhaXtCVJvis+CQQrEJ4NmB2MOcc6aAZ5c/Z2YRzsmOkwXk6iwAnXmd
VQAvATABValy498QT8O2zxSAvoFiavGHaP5MS9N0dab6kC87ZjN4GQxGURgO
PTQVXoTqB9TXoqYmvo3U/mPDjbIUmokxMW0UKhZ2qd7+e/VdJBe7yuQrmOGy
34jWv1n5PkWX8ASw8kZtshzFRYyki0/Tupvvl1eP91bLrQ7ZYdQwXxXoxofj
qaDNqUQHuRUOEhUXpwlI86zSAIihRoG7ciEmJjjZm8qc/ZGfbS3FrywtJZxI
zpdCahrfQ0p+/MN8GLJqn3Rv4AJfmQlfCLSLPkIcMzVJqINpXwxVvGR/I1BN
E8T+0NlmYiHGU09aq34+I16j4VGgQz4oqJ6iwv4c3XQ7h3MfboJT4Nr9XZIq
xzH8FRPS4gEx/r8pX4RKr7auhnQAjcpJygFk1hBC+fm0YaoUbVXy5B+i1MWy
0ykw+d75owl4dj3TKvkjqQHbFfTwkW13E5AHUi4WMj/v05QwgbvZGLBwBiLK
l4+oAs4XFPU/Wc86K3dzRroYoVin85BO1LFY44qTG3FlD0bBt8egKm6Q3xwa
wY1wQrYElSCiGrhA4r2GAN63/588p56M+AmlMz5Fvm6fKFCGikRCP09QpdbM
/sinlndSpuZQAMvphtA+yzQ105qdQ+HVXg8itF86d9k5M8jiW8Lj0bE6Adyd
byRFc5El8foLy/fpQ6JsAQGWbVgFAnc70I4ZthIm3PXtt2jsw+uqqs1kfpzM
MYh+pPhkq0phcyELrkXfj6ORgOl0l1/mTXlsMxegGL52WQ/JL/1eLCqm3d1e
hpPfnA0h4sA/gSUImRD8zo2lHLvJ7JVes2q5XQjhW3lDKMSO5m5BaypFs+ya
8/JukxBAs0d2HM0mbwEMSza4cZXp7juZnFtGubU/7OU/4EQi4hOEvSg/6mJm
HSb+TwLWXGYVUnnM8xKrBj12JkJMxuKL7TXBIEkIrC26DZ2UufHUEq6WT3/C
8pgKPDZ++/U6IrK4tMWqSOhbYGcKSIMuv5ijSZVsgqfmCaGfT35nliT+rcCK
HTL4qfFi0OSw50H4c1uoDirdxSBtrX97V5qkLzFRDm0Pn6nkQk3eGK9stQCd
Z0BRWeMs8i38kU50oX7P/7vdqO3cV9togi0IIGw5x2udFtmuvojy1O4SLbBW
OcjHm6zMcsV7y2d9nvbYKPMujBRjqoOBy6sW2cBNI8ilGgcXdCfwSpO4MVMI
Wpeh5/SkAnQCz1ROGG/QNboPpXv3ULWzYgKFuJ8OKRwphQfyyX1FJU4YcaIg
KuJZ8JsLZv3E/Ka9hDOMCz/yISA85t/pONgzOQfVk+v0KxxOrUIZhxzkof9y
ZbR3PBhSgYl36WPiBE64BTZUWeLx0N0Nn/YhMxNB5h1koChNVqtANGvj56uZ
la8K3VixFaBefwzYwlw1X6JUZIrxHpft6b8mUtNq4CT01pAAQNts8+CsePm1
BUxWOq/WZNJ66TdTNGA9eQbHAl5OR0HSLjQ1JGLfeWdNzynrx3oIkfHwlTDk
4rnPAmTW1A0PxZgOeazandgi294eJhKowQrMHoOn7MSUMKZVUtOKCZJG61f3
gjzsMgXprO5IJ5DG8EkEEmGgJHJWBH3/KTO0l16pQOmw6cXB1vdLk8AShnfs
BPQ+ozZAavTOYI/rGAfG8yNAP5SpJvAVLhQt6L0zKkppA4ctivhm2t9lNuui
f+S/01j+9Zhs9iXY9WINjVyAsbzCDWxSIPoCHyu3Z07klH8Rvh0VxVF4ezt/
4WhP3PWnf9JoN+ODn0xH75fI8g9HaMUu6AJS2JF3eoCsMSqj5hRVTcxuObMR
T1qO1YJarbOTZqWzbGKeBrSkWyzcNhw8ogA9xqXQWwWZsf1ssqZ4es6zhp6f
JNYFLoXn7X74MsY9j/5v7DME60olcG1sWiYImgyodyfqhx5I1WvyNc/bxJqO
uOh+knx0ppMq9N1iNpqicaqZpOVjRmfYTrcFAgTouP8u0HYGY/TAaEldCSBm
6fBCisX43VoHoPTyLuZOzK0DzRG/+XZTGGKtz9xfFi9KDVpjvKEBLNQCiBf0
7hfhZnU0FdqkGM34JOExWTr678f9uIBt1dDgk+d8RdmPMFIfoZw4WtKHN4yO
Jm9Pc1YTZxmRWn02KQpXnD7ix5J43Sv8YfwliEQdomfTBA7osAkducgtIyvB
i76qmDquggF4dXMbbP9arrgRLYQVgdn/k+IY7WZJImZU9QLJuJO4KU3OcNTe
n99yBdC1AxJXS1Bpw8CVQTyoCoHNd8GJnAtQGHfEF/gGCE9pKR0plE1mF19y
Yhqqa8BxO0A6GvllrCuWSW2KRS3li7ntyz1Ne9li5UZsmTttWE/oHbYIXI0C
joCpNAU+Jz1hcmwTPDkjknrv1SWEiGj1ZNOifGi8ieGalZnZIc6NSUltBTe2
BqzFC0gx+4NGKBzMo/Th8wOx/2Xxu2mR8/aKgXlUKvvmzJ9PoZClikh36/Ln
Z9FmCe48vqO0wzoeODOXlPBY3XWRozsFFuPrmDEMpo/iTF7HAmpA8KVEMBk2
bCSBENLndUEYCekntpra09MwGA4wp+OkRhZSNqgBCrIRbuf8H9puznMd6OZp
apBFTPGJZwtBx0jC+0DRxZWMIlbpjq3v+tyhfkYyljWHWpZsaZRgGWvacFK9
5x0HlYzRvTmsZcio28kgEUWhLV5xLyCWInb4zoAd54AU82LKzrFsf04c7YBM
XI//NBMaeyURWeeXt9cG9vKukjoxVHuXyVkqYJPhOgZbDFOfCJ4p8MnbMjFj
u2kly5F8K5QbrvtwfdcAQVXmlux3WGlkVlLkUDk8r7cZ57j34St9jqe+GE8V
3lpeOr2ah/vuFImBngG0vX8bBvsl+DQ035F98VcwaBZNh2t3GL74YHs9RVGz
BiKOX2lTlFvvls1PdhcXNnvwZT66NFtS7GzK/RNjkYVSDOHvqdujCz03Qd2/
/4zRQhtfCKNgljrFH85OuhvmSXyrVz/GfrPX3n7KlOe6Phi2rm/eoEetsWwh
RdRPpK9IlUFeFHykGJFNPO1obuIw1YsPFb8HbT3GB1jbyDoCxzbC5Ga/xX29
2OPdO+f5w0J5PcUQ80y0RTdvVk9Jt9tOdyt+iUoyMwW1JDiy+VL+J96Y/dhS
e9k8YSHZHRTMUwGkQa50Wur8Fd1iu/qwPa5Mp+PZ8mmVih+VsUoG2ICml2FV
kwC702SaSo/qXPfsffq1f5nYvVt0CUM5lKmvuAJTSAyjQvIMAsfM/Z5SMqWn
eEOQLAci0pbpCeWozXyCdJMaqnE0Hu8EEcCRzoXBlW4+N0xak4PAhBUNAvel
25DoAYLyvIROVeM9/7ylN+igoORLGg0snVDPoHxj41lFDThKPtHF0zDRYMZf
crzzEqmB7mhrG5SQLMqBmo2MjdQZLhmJ+MOYmfpYuv4hx+JowPtlsmIMzdCN
NcXSiG4eeehrOYzGRj+Ofu0mH9HV+ImOasvWruX9e79sOGpXEVjw+xW+W/2u
lcpQGyalzbNO9cZIW012nszB6RGRpIy6ySzmmsyLz93dimEygGLXIAB6IbQO
6WloCvyJBaNP4Sk5GCMCBReAOZuWseQEegFBKj8+cT+yKCW6t3hGYjt7384U
YcvesYV75aUu5uSTucN9aEAo78xFv+golWySjJlCtfs88qB7OC7jLr+Dofgg
DqRWqTgO1aRskWU1/vhkQa2x6DrRcIo9Nyx4L985RDizAmJtpjmFD/ygOy7l
b+XSqltcDrIpPfO1/gLeh9kCiCOw2VwwCRiX0XPDsDeiz0aW2YArU8xlTKvt
3vyTH5v0pcIKiv7eqowlowgOGcrjEgiRJQcDdfSEO38/zmkGgRY6g9/kTZkL
jE+VHSCfTZd17WcmJyrobSfwL2QLY89V97Pj61F+Z6FvwP1DvQla5IO13HVA
0gt0dOjDW/2nBXhTYQuyqJzRR4uvTj+ZHh5QYpuMCUo3n9gTOFjNeB6lOrzS
GI7ZHcg3MYujRQmtFb7OSXjb5lhKwKxb4x8CcWnOJr38bllQvqk8i1b5RV2n
eYfQb4mUvgXAPYY8s3fhZk4CFkAKBnknoJ+m3TlspInUeFWNAomgDLEPt92i
K/EriZkUAKc3NZvztuWHXuQe9f1f7u7lMxC9PpGipkdNy9wK8zfYXZpFZVxM
V2yDEHhTgqfJL2a/5zECwwHXd+UvHydPR+1Cm7LL4yIp1IvlDjfzpJcuQrJi
rY20YJB+umwyMgFXiO0aa0Q2Y1HEa5GLCyLiT8fvlNEWJwaL57D82CxWM/WU
e9xJgPYW5YO/xQvSEa3FGyZbR9pezufZkI9WWV9KytUNLWCHtLzX2trmbCbk
Af8ZNVeiLtkstjbm/RASQJ06c71R10wQC/mpf+DS4fkXttHNZrSR6IUMNM/y
k4Oyz5edVJyZbwT0oIqXGxFwqU79+SlSa56tQIPcfUZwZy+XBDEh715QezYl
bEDVuvAGvF3WLm5FdBz7vpSA6xRzIJQcYNOUgUEsd+joCBa96TfsxBLiAb3E
s4jfzQZ7s1oTU0GazXs1VIunrGqYw7VkEQb785d/Tukruq9MFeKxmJlC6xO/
cAkQMt/SjJwSzFGLTQiDLbJKWAv/J1LyUGSrUAZ3VnMYLMz19asYIOpnTf/I
CKLVkML1ijVETzMuQM8vRWp5PTSd4Bn3TTOR6Z5e9ky9WbFdfOgkz0crnu3K
nTbYimHiV3EvJDh+wKCRlF3fZlJSB0eBuAsXhgBAcUIYq4FLJcQfnwm+XirW
xmc6IJ96J1ZU275dO07YwmOUsLuCdLHCK9+0EcPdd8/TBzqdj0iDH6PcbO2G
V9NDCZieP1oRr7yryI0KFYoVdZlnxPSc0c7qVfmrROtShVOWvoA2ZHtPrOhI
LQDWbjqDMhSSTQvB4V/vX7maDCIEYpbeu+V+HQTclLQeLHy5a2/ZDFv6uwlW
78/xzLSiyq852SfMTSK6iZ6mLoFEXMxh33dLcmtTuui4bJ8RRa0OUCFJZ1sC
thRpQwTxlPPvB8eu1IGr0O6IIoxtazM25Qv/dElPN3jVbRH0ecuQoSPxdQay
VBw093xSGZ3sydeaUe8b96cZ0OFU0Ethgb125HIONafMnWJHBap/W8ws9zCV
87z9ZtBnBLaFOg3C3ugampd7QWBx8+x4D/5/flPxPoR6ETxW6ehwQD1DLyuh
Y+YrY+dZUQTzcGqe3raRkyqZVnj8+WRivtY5T6aKqsRavLek3jpx2I40/hwb
64d2J7mE4FmBJZ6E1Y8yonlSY8Ly0etukJ5xvVVTrYhZtiKRxDo5V/1mdjIs
EnnF6QgS+HvTPE6gipaYysgWfzDsGFRXtDFlt7ulSpCo7sxNBOAGR95h0I3B
TozwL7Aptb8rOWcUDzZqvSPwl8IxlhSHjSZucLZsKKLuSzVDy4XJOhE3F8ka
aq54LsT144e6imsmor/PfNMYXip1HDtmKfVVHNTq3mZ6/DnyjqGj5KvLmEMY
Ir3enHdNU1sClGUqj6bBO3+ff48PPr0yQJX9rGPC/5zbCVkLW1zwxti+wWhg
zuqX3unz9rxc4rFRSt7P7oGAz3K/5Sax+fS9Y1TPl8F7VBzQZhym25lJAS0T
/rtDZsM/taZX5ZsmsrH1bYko2QOD7uUAAwM0bzu7PPuPZ4LeBRHW1ZC7Phi4
4YZsZvr8RKbduqw72kZ0eo/B374n7887LyhhgcDo30yfdIf3+VkS8pn5ercf
+5Yb5KhTH8uDf7PPPsBXUFj6/i0twMk48Xp+FqdRRUDyrVP7wxX8drfX/rgx
bqbmesw1bK/WbZ6DzWFTm2Va79g6sgrcZ9/ciOVw/bKGVfjA+4Tpju/Aps8D
u8hbteHo5/XAcr3LV2Zd++CRPruE42xfYdm7KFgD6WSnm8cxogYHRSFQCdqc
sstH117N95hg7mrBVdDFmSl843jcVl5LFM1uSXcTcX7GbAi4zcwg1FXoVV4G
Ry5MyxNu2+vawR4xqqolecibJ5xTNm1g6fw+Xi9s4lbDOsgX8K0o0YiGPdF6
HEbjyqIGzYsbP5MZRwyMrL/j89fFcJXo0t6g11jg24Br419j9nLgv2gOXVoJ
XunbGF1/t7UVYWlRs3nPit8eHY47GuA/ysIckvIrNtcFFmv3qcIK+j7CuixJ
cr7K/vA0OalP/ERKK3p3+NgoUwz/UjE36xtryaLoGRmZ9kofL5oOu1YHleDn
Op7Wtl4CkOS4CNXrIzPD6SBiL57KUBqXPXf2zV1YBjLSRdH2aIeDeiNfVQ2O
XHOfrA1QpG9CJ/9tK42BM2wmO2RycbuceCSFWnoGph+rIN4kvvr9BtTkI1FE
yIeQo+VHZWT070wRHg0psnRAwQLHVrQ2JN4OV1xocWzOLpnmYO5FNGrC1zw6
ONYziUaAuPuK2oNbHBOvSBXCYB8rTIGBFCtzD+8nFXe42m/gzYJSpbid4Vqg
39Htwu2arqLecS4AE0Woq8ZQHdVS6BQXkKbiupu98vGkFuTpdve0R5KEFA3D
p6CP1tyFRO/1hojxI3Xs4ras7dvm7U1l43O8e7hOfE+h2OqUWkKiSfvgtcY6
RYvI66gkQjH4lwmYSqn7oWtXf4+CWuDr6wonlOGuVw+1r33ErRSMqXgbyS3X
xvPc+k1sltp9BheViLRg6n3tlq28t9fBmfgnYv3+00lbPEPWg4aWM3Iz6mHf
DM/g4pWJpC8h9RIw/jh8XFe7smSg+5SQIc5hjErkKmfC2lVMpfOQXyXpyidm
xaE/5lpD/PhzT+mAiiYhR9rTaH7bAvR7yVGFC/VU4ouf6yIsyLaI+GI7FC/7
UCW2EHPvxhBZMt5PF2gv/ex2tDNz9b9t5tZ00IF5zuOmQDYZAh5oopuHvAz6
0lS5mwLIahfxgrFNiKuIxCFcskH1Ef2as/CfPj3Zn4njE/BGvS062/9aCQlx
IG7Xk0Z0hwzbHBQTvRIhVVozyaCWyam0MaM4n4KdJcBirIsUGT8Xu4YwAeDQ
PXGFq/4f1n54S0JCb7QviNZgLC49SwtTe5GCrtJFoFVwIupAexogW2e5efIy
GoKlZrioZrGJkjq/EqUukfvtLkRo+fII4hc9BHgvo5y7WnYuLL1XUSkhyPqO
YVbAAr11XCkvyPqNLrQXUv/n37IT/JKLoTHS31BXVBDIwvWlf+0eTF3YLk14
kasS30zbHykEt4EnwxstxWo3VvZ+6nTxejv7eI8AIHHuNgEe8URc3iu70R5D
3le+QeADrRF1afNinLE9vtSOKEoWPLXXavGW3buIXw/wIAkMoAC8TWW4G7dV
ekOs8IxFgu3JeG3YFIWj+4twVSHL/a9CDr5zd7tqD35TFUF7HdGG0+iwAQdO
d7gBvy0ejvQhlV0VHGlKMe32ucCPDnCvSBvbRnpoL2SWwQRvOEYoNeQOmVZC
HxKwv9+ZmWr1umRnz5FIe/L6jW/cEWJ/msVJ6tEdKoRzxwsdgcyilQzP2xVi
sRRcFc6CFQNApMTTdAc+/VVNwtaSj2X4P95tBZlmSlFz/xy9Gdwi4pHJ+P3B
UvqasT0p4FSPV71td1qLUISxGpWURsvXewQY8HoLeiNpiezUWME7YyMAWNN1
RtBZJc0znIJySsZd3VZVpXricQPjAI5Htiyrg65PcqRvEYiBTiWpmNeYAKh6
E1b8Nxr6PeY0193KT6aRReWYapUOfIwQme98nFpaOupTxCDpKTdzdVKwoe54
mRGvDoYQOLHHjboDwFcbWbT7KzCGkaxJFPRnQRqgpCX/yWDjKCJhc9oBgL/3
8ue1oR2zEl+Y469FdwY7jO4561sCtxkD0gW4NEUaMHF7wF7NpVq1mjuWzqwE
/Sogi3tLOGsTaJHPzAGtnsEORnOIV+HJz1ISWfE6mAOSGWZJ5XD+icozX2aV
GdXGnRt7eggToYyObndaaD/GU0ntlUGKqjMpTqFyZRQqLY/yU51fIXmb7SU+
DzuKfekspd7QYOC129ze9O7IkBRLupAY24Ry5Svxa7QhTMXoBzzGwZbTqHm/
Uxehj6MU1aUFmSa31jQ9uSxYD6AcDY4PGwpbiDD6JQlnfVvwNBo/z0XVDQ6D
vdxiJQfejb7spfaSFKv17wSI+iXhHzGiKfqryl5+si6X3QVFtNGmLYn1uJFP
INeDlUzpOvUXm24WjNJyo8riIOm0FdMlLaJFSma7ezK2aQlaujDJOS3o0RbX
qwMCNkwDaEFQZ9BQ4x2biWF6hDhCoW+5sBDR4F7kV1zGsTI7OXqkKdz+dLlZ
q1+HRF4aJW9uOxkVpFuICOYU7zgQcKLsBJ1lpgXkmsEiImgkXNCW4H9Vopvr
9WMHZNIGKxAvYHT7Hb1MoBWR2IIMKliQ76JTeEnUARRRejSJ4+WxdQS3LG1s
jvsZo67fR57n6ZRAS/RkZADhT+861QWmgg7DWccvWZZBU+bioepzNeHo4j7T
9UtgupIt8tB+l9lwjC7YfktDT+m5IgWYv3/QehF8tFiqmAgH9X0aC2tkWGMk
UDgdT292X7Cfg1jles9iTNM1N6ZSDIa9pabQxGK9N2y16I2IJyRU6S5Q8X14
mI9FY+UJC69P4z1xz2eAxDYs8cIPGD9umfffSxSuMAT9JUjKkamP8JYcqA0r
f6nSV+ZkLL2oBU5MzVSoT9in2T0GPQIdGuIVplzieQW6PRriGYXHNRswpXT4
PhCifIWkom4Hu8lZGfNPW9ZCka/cET1Dj9Pk8DyUQ2tLwLknwY6YaoXdVqa/
jsWIB1LPmk5MfodHrM2SZyIyE+3L3gfr83i8vQgPiYczLccRe2EGrXdzH4k0
M5CrVdKAcmJ0+V2vtrSq17XeMMS8sLXuuMtyAtMsY5EXUyshT1j+UMihbNFs
0dLgVJCWOXIeIEu3Afp3lZSqT6K2XaWecV33IrEr0tserPkfFUBY4eg1hD23
ViJC6sH7GKvJqm84emvBIPh/Z+UPGqLw1CFhZgrHJ1YgjCj1ulM6Ewe7xhNi
EA51Ea3Mv9t7Du04i0xyHlAVaTXXfWJ6nv/lijAr3VlnbbpN6KY9A4j1ZEmt
5Xf0TiZNaySrZF32L7x3b/s7FtOL5KvgLYZpWIRLpJfNVxHJnWT9qL4l0POX
GF1BWS8zc9D29waeJR8ZdYgyw0h209iNFTRUf6d4pUR681BHyqAvHoSYtO23
M4ZcWtlG9GQOEQsn0g9VX0tvpyDzGUQwzs/0V+vm1EG3iFLVxj1mdSQgzRjG
KN0yibdFFFIeTHV0tkxlRdWjRorLISYM91/7XyiztlFd+pYRmEfVefWd7hCp
l5Es2QLK3odifw8As10Bfel87N4kgqC7WwGlywbPmdD99/xKklSgJ7BwjiNt
9zWvZMPGcdBPu6wz5JwuGs0cOubRGsyYWCXUPA2PIVEEJY9FxZFB/BCX75hQ
vJ+SEPdItjwcbbLcdnh7M4lbCJmFGIrQ8hXtM2J4RqxiojhGKw7FK14axXZl
zcan8vTNKVfX0Xh3CFmJN/zk/4LUZ/Q9IIWWDBbTPD0Ea+eRWay99fOfKagg
DcT8uzBYpqKRnJTUZyDAM5P3Tn9l2NwtvkXsjjN6VakcB7pBm3B9o1AuOFqH
JmxOrmQgVz1y4ilpaQwMT7nO6Oy29JuOCmGxW+V6di0HyFfJIe0rlLG4UcUX
LfwIMqvh9aDMqpW+LpMXOW/U/ZauzgpYP/s76AO/vjZewSP3DPAj5qa2JaJ4
7NpqFOJHT+Z9R01WApo5lQ3PWOP4zKWGdjHJNFX/X25r5DOXzLumOl//e4tP
hoPh+FlGplylXJbhe4aLy/e06RWScbsOJa2tMU7dYlHg27hlbzFitXp9FIqd
bWKQ9HgR6Ka+xa6FR1IxBzkorZw+29MHHCeYv/R2yc5STc6jIfgY9cStwG+0
Wjvg2OLD0gktRwJ28Sp+DbjF3fS+YLLzD9GCa9IjW8KT10k/C2v4OjpvNehF
07y0tzr8opjGyMe7+qXW1ts6AGfXLmh5zW1p/AMzLKTpuiVy1eq+vGpqETRI
Wt1bVVleM41kvPydXQWf7li5VQaNrZFZSmQkRcPYX4NYORUTb1EYiVvDpNlW
ASaWnLmJHu23EBT1enAQU0kxzk1nYeZ0MIbLybobmQYPCJI4WWNRB7czdzxT
5IonYk9tsQ3gP+kIsgQMtKqn0J5DErNMkI3klnIwgg13xgP1WcvJqEk45HLz
dD473MEL+cNdNj5pfWDaPaZ5+d9hAXK/q+h/pAqUDTqzFperEV843iAkOJ+E
Qnklg4YT33JyrkBtzp5FR/eiKbiAPH67IR9KPh4xTobq86UavY5RxvRP5ohQ
vfO4jvDeY8ga7dsYzlZxQS9fD0uia/Z6BPsgqF3NQh0/9u3w0seZsUyEC+9Z
0wUrDaU8Hp9psxqeI5Ql0lGxTl85w988327sFRr6oIn0JPTKFGmn1qmI4Zvx
jUbbFDV0sXqetIw7yweEx7moiMf8SYepP/QcTQX21YUz4JTxs4Qs9ZKgk+n8
Feki7gKcYdP/4JMMSWVlKrCpyHBEGAiezXuTb5YjIsWRdyIS+kqW8sC1X6uX
ubI9OMxoIEDeGU8XurU/fYOS9yv+vaSfWwOtarEB9ndXGITopihaIfRwtusX
F56R6lP+osjMbnashLTMDAO25Z6PBom9Q4kooI6lvPtLO6BwYfSP0kvWOk2y
UHuzXK26yRraAptB3GMFkxAmS9SnSSqJhgCrR09rbiAfMGkiNR9z1eQ+2AmT
Hnn1RfJZubrPbQCzXH7ZAWcKqFbQhXgAnCYPKEUigdOHoXY0wNGFJ7g3iedF
XrXkn/4q13Tvgkg+I6yJdouMOIY8+LYFyVGI8X/y5FgxQZ7EfGSzgRZEkLNh
VLShbTN/xb0jf4K3406eCjePmzKOdhYwTdSxvQJVCgzJj2VamnNu5bJB6pKL
EK66ggvbnseVVFWQyRJjW3QgA1Nvk6kzCzKlNJ9tDEnuR3poiZYU8dbGCB0k
pIKG9O3D6OliAmO2HC5ifZjINZhVODe/3uXWp8P5yuGcz5Ltr0JC3+vHSVIP
ribgqA7LtyLvKQqWOIUGsRdVx0BqhT/Wk7l1xBzVcgC6TDpcTdJ4mhWd5+/C
TjwzQEQs5ZKoL5CrR+7YNOJc3AyFbJBfcmaYudadiahu2SZ185wy857UL9IN
sODe3PgNDuQ7fhfYUg2Sx4bsvtarFWxSD/ksU79REnfALpoNMfvMOZqmIBZD
h4NRdYuHc+wKXMe70qHTLNHKNGs9SYrnHKsRiwJk0A+cyQoqbUQROG5zIMNg
+MDFqCPDPFoF7onWyxHEIdsUt8bIDpWTExN/32Cf1hYjRqqlMnz7snDHuojT
CBGSS2J/EQj6xdjBhJsA74cn8x0uN1wuD3D2ZAIHctmXUze+GfUaCg0I4iOw
88kEBXP1YHGui92tlakXDky0flaEm4AbJ9X7GeUC9pMhzADI1fRym5S5/uCl
1SuhHeuuOeCZzezJ0Z0c2Xlgm/fV+LWheYr51RPq+JGlHwxx09k3gGQoLjDD
6i0nB5Wz+4YgzzeTlzS2EQJein6KfUkSjAZG0qhLNTzCGQB2B6RU/Y8hAHgp
I6wcp8F6E6Le3VznsQbyzDZayfA1sGCEnFlk9oRn0UlS6EJv4cLFSOaygqqI
EeXBSib8K6jewhglF0y1cgsJvzSyn6PzhfdB0BnbI/Tw1X3hlgHMohpI90eM
x7gejrcKS+DvND7xfcgbKe26wmcgX3bJAFwArvWqkZcgx2TiUoLBt3wLTUha
YkDBXBAD/qxMoWK+W0ZDDa2anN5I+YVT7kAa6wf7gxmxEa5TrQ07pb6cIakV
CWiWtHVPdHCRy1K09JBvFkKE0f3zAqKwrcxVxsggUglDIJfPXDPn7n9A5b9I
miOSVw9VwF+gFESq9Tj/cLbs1ajNCxyp8DAXeZhRhOV6iO7fEQpm26d8ifc3
CJBiXh3uIAZP63BI5EwwugYyIKX+5iojWuObsOeoDho+aJc8R81gnPrRTLfC
OYrD9VSBNh/dS3QBO0Nu6dPIrrW8w3gzTLOtxIw3Dss71ga3lyz8a7149uzx
KjHAAq3yCRRSLoV+7KgPqetLn2SRAojFsuSQsoetoCIwVQNEYzkLHh0A8Snq
yIjrsLYYkloxSVv8FjIYSwE04mtDllJ3AF7JD0TDEfTEWPsZUnYf6lBPAQgk
EJgNT0NAL8e1htEEZ/ISHlv39Sewo+h2AqdmIWRwzsAquv9g01OenHEcYsVZ
Q6DGv/RRol6ka8Ybi2ZZ07qHr8vg+9bgzvlAm+9wejYLO0unbi5dDM9w+Xcm
LFedkH20tZm6LCyBHOghR9JPFgvxLN4ZojVyDUU4w+sWuH6JyW6IBQSpwoSv
3NJ60qAzpaVOuxlJrJipWIGAdR7qnZ/hAwc16fj2drIyAqx12KY6FK1ub3yg
+EfEKbB3XTlgcki8CV8T5ABqk2w+LD0aXSUGbVj3uz+ZFb5mdYplfNcLJbIx
RncABZ9BISsFQHJ62Ck8DYtzqTLbJJgJuBhcoEDRgIFUnpOMcTCZtntGVd3k
VmdvVjDODIxamJ13JdHIiC7/L9VwuFxTBxoA+XOGHapmdMZfxlkW7U024mTS
9E6WlL0RA6p2bL1Vwp33UWAmXCWy2/lXaKOBnIXcI70FOeWJKpUOy1zdN16W
Ss7cHGZoLPDqos9AdYbtARvQ9+RwjEnQeAfDO0poATn3acBjJKp90iGLYKd2
mESTP69CZFC22ulchEg5kjiaUTO1oOnDvOZWTNY4I7t78ZGT9SSEqr1VbpJI
JTmoqKyyNhDdkdwL2h/2goTLj9C35lQgqgLdcxzlBGBRnRXqTxKHSe4uu7IX
R5HB4hjxRfNnRva5PBzRVINMoYIqtDFCKIqi8/VFPWONSw4ZW8GVgT9CZaUQ
NmiFDPp6QWtyi9J+OAkkxrQyUsgeI8B4affRKq29LoaFK+WV0eYDGNyOa5n8
VOp1tpv05pTfLnd6QT4lP5t3QO59Id+64/m3WfTg7TH22q4H6bMQvhgRv/mX
xwHNmd4QlRfgvF7MgqQdT2P+/uhrgx8Os4FYiyAsMwbbMmgi9TGijgr0TXEd
WMZtyUKAxyylmgv/AcidhRUsislq9gxUX07Hl+hz3AEC4FrSIhukeVcvW57L
2VIcXECDsJUzy77JOBb0uKifmB/teXQXSBYJU/0yWrb4LM3v65hHyWPpfzkM
Zbwy+bqyj0k7vwKEx0N7uTWbxNvrg4tkqhkp4MJLLd0zKls8k678rN0rOjpD
vduD9o5R55KazEYzSQK92yJeLlkGGjtNIy0QyOR9v6IBiQRKRj25kv/Jkdda
irpFME1nTatb8rEWggt05bEcImA5MokmTBnPUT7azDXahtYsCokxYdlsyixZ
GoLaqHyTIrFTCB6gfM81dXScT0sFM4yVywGXigChOwByGRpVzipiWNdygdHT
P1KCFF5zL2EI2Ha6//KlgY2gHwa7hKWSk7pyKSye2yjuMpdzqJpJeoc4DI/k
lGtJRInRZFgwjWz/eZEBpaDuR8E1WYBM03YkLaxnO6/iiaph3WxBRjFGpRZF
OsKihJrzcR79Ki13ZK5kcVYYe83H58MLIF6Vzgs7lF09kJKigdd02OMV9NBy
AhdE1Rwzs3MdSktWoRNYQcl488P1frs9SKHUmTaTVFCAdNd84QFRiJ7hg+2I
qlwPP2Zmls+wRR3SHo9k4zoaQknBPZMxK8CjCj/t9h1MUNe+F7chJECDDfB4
G3R11qZvp+ij+ci9TdT9kASxZmJh+rStlc746Cc/TpU3SC4BY0u5ANMDrRxB
2X6QJj7LyNVCGskN/FPHYxn8GN9wCaJuT9jfV8zvWTDG/YLfdBMfA95lTwqf
pBh27a3T55jgx/I2JmuhvF0yScmWdJQExYEduQtNOpQSeflFJf10hcP4yoWB
ztV4JqGxvMeSLTfD8UnjsvlUgjE5jQviRU2D2ClzhvuQ/cfXPPqL2K2OJCSZ
f3Hy6woIajQPF8C7o1k6w6F7LU42Vz02xdDbROpWHv1x6R43fSBAUZIY4AIt
zCkcZ6d45Uwtyd/ivYkYDfw6Uay9QMz4FxmH1WkD8pVmfbVLt9VJfO+A24hh
MMlDN6cq+ovX2sb/RAIIl6xj9drdMT3U6XntHW+cHhigJ5WYXUGAQBghsdZn
WFT7wIV0z7hNpTTwtiMm/9Cj7AOO9rP8hQnRIEZHOzZE54i5leyc3pjJln02
5tnqebVUJ+Ye9/9NiqXf1a7SIfL8F9IG27DfLioawHKNmFpP5ByBykGhPrc5
XiFFOkG1oi2czn9kvF/NDSPX6EmfLG5v96kk/vWaqsdUe2hQTjjJDv23hfaz
lMYhgNsefzPCCzF+bOU7MSmBiEQcGeZoxk5Zj2wbxCuhlofkgqL3oPdgg6T/
+dp6eTsJm8gJCcU1PXg7Ai1LangaaxyQpXbEtXpEy5g/uF/v8sgzmUPcZHkO
ZeYLdkXTjvPN/+JFZY1V4DLshA2swAoHedj+SSkGu/JYpgPspq07x0LAELIo
ptrBmfGGGu5C4vcdtCZ9FK96hLwIJMN8sm1ErB0eDj+i/gKQ1b/aZE3KMW69
Hyckauka2xWoGtFmdHlPVXm7pAYhhVvtGB+lzkwXfnIr/cNmLSR9fTTfC5rx
LLWXiUIO+zXDMrDWgcRFV48e/KAp1YG3OpCF8yw6O3xYqEUy5M3MG10w8dDL
6yAWsAk+BhoS8J+Xc2czV9T6HtOo9pyOfdshhQ4Owd4q+GgJ4xHDFyf+eIOS
G0y59IWO+YHtxbjFb0WJjLILI84QjmSGFszPUJdY+qGfhNRliVZ0VvrhR6tn
CvI1FhArH/Sm+NNXSjeKio5ykb8HQxqcoTEkkqZK6D1oCuwU7pXmOhen/PEd
Wtk7/mmZPrz02cGmjBrtyn/qwCe9D8/QoetJQEuv+SNpJwIqGiMkDGZ9W/Ns
iO/t2OA8t2iFz19YIvSty6x3OB0jWhHRad2vN2OY8dfjvimcoFvoOgR4lys2
z29AfFJKXcdOrmNV//strYyUjK20KggddQQQBaPSeEemX5KfWoVtQHOML8fX
9g4RP/X+h3R5nWoKkV5pbMuf+GfXNmrv/QS0sF7b4abCwjYXwKPKVqSWhuIj
vBr54TeJQSgcWOh62yjRWKZjbPD9OC30RI0oEN7mOU4PudRXcvizSvlxy2U4
N/ALo6bXxSlAArnsYte8SQB+bkLH1wwEQfDq1ITuklqbRzwTQCc7E/Gg0Pek
Iq7h3ny1TrTF0iqbzV8CpyXE32Pz3eDId6KdFB9mwbnDbpG+1dtetvN3utbZ
pUefxaBNCMo2M0x+QOtAZFpeMDneDbhIWkpju9tRqU++CQNqNki2kFnaDTGf
lYT28mYU1rMo1TAhAeb43mWHdPGKKJ0DQh9rT0vzJnz7IkPG1QfXohtShT5i
NhSFYs90NM+lH2FfMEZrRQcFD1XBJItSAiU6Hlcxch45tHjo9SHaXIZtzN2p
cmrZtWDMvh0SXl1pPDsutp5NvmNOxYumTaGNrI2tMw6W8lZT/mdOwZMAuGIk
x69syOl9TCxCWSvaasU/DqjSPDu0tT+44hPVXcbX9WZ06E8LVX2biH6mxU86
+FEUliDNzGh9i4pgtO4WY5m4vEWRbQu+WpWLNywy6PfkA/us6732gpKot1AI
oGfq3ahGorADWF2csvH551141hsP3VO1ufuz5XV44FVaGHMIwO+weHTBFTOE
6icdzQLN96cGAW4hmBZ4bxknasjVnM5iNESAcDfnzRwyxAVCztzGMmC6+OSo
PYEE/MgTywIQYed67zoalFgRwxC7yDZeYB2PGGnC+2kuSPMLUDwDPz/9CH+o
zGpoG01lu1E9jeyM67HdH6gtjKhJuM4pRs0KOq9ds/8Y0Hm1jpn2q3BCcQQ0
+C/BVoFKFtoXbw6GXZYcv+/DY7wKsgzjv8o/0ZQ0iuoIzLboN0nruAx8Ii50
bUDXxoP/XRiRCQYooI0ZXKkEEJQOeTR4CFiisARLqiwdJeWR9DOKHRqtH2A1
FLFe1xHKyAH388kSVCwQR7fDR4cipQIkrIHjUGdERbevBOGOKZT883hKkdug
FnaSc+SgAb50gHFb3d6FCVAFqgltlUDyp5OikvumVrAltP4KW5enJHfH7GCm
CMbm8evYJn8l3GFPWYPNRnIKNVGaNIwuJh2V3Skwdb0rTH1c9KMOPXKaiVLZ
c6eQfjPG222n9Dn34141kPH7sVSyDqHGCTco8yUfZ5O7luoiF5he1M4EnHb0
VsmfIEa867Su/L+/WeRte8eGIa6I1f0iFKPcGqKBHlqlQnOhZXcOAQZGW1L0
kqdg//F8mq4IXJhOFScdOPQsNPvvxD0dXUVNkcy2NF4iWS8xVElMReebtq+5
RbCgOQ/wAW9OFnvWQg2qi9T34LGO4fOoPp8eQBcX7g7JoR5zgf9q5XhvvnQ+
Rxle4CFdL06TbEDZ7THrQVngeO3U2PY79pokp5cB0koDfY+nTiCfNVWBIoqG
Hdrpx8G97UpE5Y4W7MYUGiqjns6SdWVGjKX6SOwaUVYLimA/iDa3SUGAxw/2
QaWndPMGRgSipuqBl9+7SjO7h8zGSyz9xMep3d7W3GLfzFnBsAneNrHVrLsO
espG7C4CeRH6wX0B2+g/pkf9MEyXOLP805N0DaAyAMW8x1GFu7A/HiHz3OKo
5rN3l5p8FPy2/0ZfqTdgDVJqxzeNOj9XtFTMTd35Hx7stmVJQKotrAwW3QvL
TnjRYEldvAD7u4K1XzqP/T/OkWZ46A+a57d6vjz1Fdx4Kfe4CHIaju3HqJrW
c/F2aqRRDVK66VNFKzHiBhsFvOv+6/0emDQVjkn1Z3h6Qs61EJOArFEFL4pO
69MZhryUF8dreEh8No53Lsb3Wj83u8hzAgU8Z5y+TCC2yDtbSpihZOwTSCBb
I2sv1NiT3OHyTgbhoudL9ZZjHfGNFPn37rDkdXwZ4oF4biOjY50/IqKX5uIg
zvLNKy08iiARY935SK6FmsJ4XIF74DO/MX6M+YTT1r7bgcUw9Ch5OB/VbfiU
WmusR/9WHH4dIddea+YDJlVZYu5CuF7nmIDbG9OzIZnpOb7ZC66Lo+uuzvrg
ZZQmG5+O4Xk5eMn08i61vAnGiN9yUtqOB3M/4UpBUN+Kq+JR2mCJZEIfR5/C
Oui1s5OqIley0LEEzTxPICwAAGXkxtuJYZgEbo7Qi+htkBZBMPeameLv9ba3
dgl7lzXU5N0EYjgvv7HA9mJua6hhzCrQEV1+RRNZA0D4LNzFK5AbPzCbxQcW
y9mGXSKEWTQn44wJ8i9hxqvvhWUOTOJJEgiyI5RfISKCkeuyUizu1XkVSrkd
Yb2uPm0+rG6IRsi1/OyFORJYOczlL0hZnacbAtxh+0xnBkQWBCpEw+hi2g+O
YP8int3oyHsI1rl8lXRrUyTYYXaqOMGff74KcFd3vul9wmH8fxGoDe8FgmaO
qjHkR4oX+sQpwLXFKJjpKHgnId41sevu7ssWqC341L1hVP4bbGmBwI1JX4SN
GDarjnetsZQM0TzU2e2J4/ToALJ/55BWYbPKJguf6qnHc0pEyRiGqoWEOSzt
L0ANbvE7Tn4berIke/z44s81sCiaOwiuGqqgrkP0knhiVvnTz3H7vusJM1Ur
doLSlMt39d9e4nS5Nb+omsyX76YFY/X3g/GOgWPR8vckqj/WDlsiVJc3nIoO
+llqSowbioFXY7HL3b897sB2g7EYAtlaxNdUvDZyhk4wiqagPVr/bv/EoWaX
2pkcVVNbqwYP6S3ZKqjVm6/w8H/OdUu0aRlUT4xd1ZnhW/pIlrMueqO36uX3
3esrcjq/XWxlS30aFm721nazWqHCUqyEr/WcHMYPT14jAV8SJFfNiLsXrnam
S+9wEZ1MNAUMzetLot36Wn4D+dOlWpXdOHhZCjh6RJzImK1h5ICH13AHnH5e
sQ9W58zpJ3J8HzAQzEwiTqSVCfySP+Z9OdGmMioUk/BAyVoT/kAM78UYjrTl
lFc2Gx007S+f4yh9WdzDjRSbMm2DzqqCJVPuEfmL+c5T5QsLOuckRrXCEio8
5qbwHN2tvwAA+lD47rlzktuUnyHzhT2aqu0ZFWrbrJnBlzD7kheuhmy2vbwl
pg2+Lu7tl2WIexHFnJvHhwLY/k5pGKQY2ZGtuMzil8hb+mDm/trmFfLi1ft4
ZHnYvwFrKshTRNw0RUkTnS+gcbgw8RMJX/aD3Z6iWV/SeYGN4IhS4xq60cJ7
7z9/MMV5hebjCuSyuneAnzMT2NzgHpwsW9WRD0Qm0/py/gA0Kco7XSdoYM+P
CfnZefRc8+RCjjWvz9X4GxLt8ElB4AHd2AMNHYgi0GWoseOK5hJrRvOPqb+L
Ke/gsFwU4aXxEfMtj+T6vkKhOwjJr5DsOWhEDebpsTDK59Z8Kv3ZhD2d+9vL
B6ywISmNGUehdwCOJlAHnaZ+aWJ7/pvEr+oZWvvYTh0TMff1uJwC/oseMuJD
wYrhEVezkl0DWCFo2Hsv5vRqHSaQVBVKr/kJeCeNjUL8qfyfo32u/hzF17qh
nAlnxk40HsHWd52CwEfYts9I2JCU7zHprd3Mrmhn7l0depp4xMSHg1JADJea
qW8iO/2M5bMtR+/neT7QoQu611lRKHTmFV844X61PsFRSCDVsEP7UHTRg7FR
HGE+6+nlM13qAzFev7HetmlBMUA1vJjRTxBBuU5nrFs8gsecfpUOTGSC+gmK
bSVDw1Wut7pd4+grBsWDv6QIbZ7ESx0g1dYsVQMU+aqoikcGeET1IXusNxtO
ZMG7YYUEWAXYVVV3cWd8d2I1cAVJwfQVDAdhGBmf6LIh89boNb95goJPWGz5
elZfWOxLguUM+1px1W1cyuNXaraHItcN4sTIeWAxTTVDkL9ThLRQ2L2ZRsuj
Kb6sQQHTWGZm8wcJue+Ns5gOfvNf05MQ+tWZ7nTsEA3UCNJtIKdTHXy3lUrd
1hDzlpt/Vgbl3KhKdV1boqwqHJteq4w9rpERYG2dYz4M7oXnBgB5FYK3xC/D
J30IsHksMBZAN7cuPq5ZYUFBbp6MmiChdCf9T09LyjbZfEKplxojz8q6lDoo
rbjdaFrDW0zEZpwQFWjN4j/IS80VeQAApXUJRw9XktQ1mGV1GHm9NEuoRDvq
ADPYdK6X9E14CmIm0gPFeZpkOdy7Yk0jUiNEzSOnFsYZJTFUjTDztNvITiNE
x++Vg+U2lFB0fOigmP2Y6PtkrIjkP1o72WmV8n7ddj5CMOnnSDtOleMkw8F8
dWfy+9i/h7NAzRTzieLn18P0Q20jz4220iydsWRL/tYp7g/EhtOfQeocSb0D
DSoR1mNjR/JeV7IU5bOl2urXQ6GkapKDPR3IQwkAEch5Q+S/lYrBGWZSiVjH
KP/GxnBICgJkUV8w72SowHISBiKr+MKUA4WkuAZ81djUgH9+1fph7rRrfiTE
T+3dz4OMyPAwXEl9jnavLh5Qb8OdC5muZ9KcePthdVtJR+dyWLGXt0Q/q8Kt
j1CZ5/Oj9ePqfBXGtQKxRtvESeQyhHO6VKMoM9aTkpAsTgZtnXJ1n2G8ddAf
k9QP+uwUqv0rdkJmAan/X84SuFaYe13I4P5NMGcNJaGe+02cVhDJei9/FbUW
Jee+KxXo0KXcr0jgdTd8qeFwAMBVVIyNnRBKSBbWrAsL/xk12Gqqo+nTiqu+
kUNsetGrXa6Xt+JOY58X8t50366c4YFO9xWMKIJVddlxB18UkDJdTDvuDT/K
ZSxui0ziKv+NFRUA2IHDAemAzruHK9cuvB5CUGSOnzfQh31/xANYLEYx/h4o
aTP8bdjiuve0k/xMaIm04ovGDbYZm7kslhDxx6FDSt3aNXK72bdpRocP0PP5
4DVAyAXYav6NEF25lfvhuJGVYCy05mw27Sxzp8FxW5ttVAJaSm6D5NboOLlA
kdoW8p6oX4p+5tFP5WHFxkvGnvs7yHIygvR4Vmn2TXRzTYv9rLfh7iIXSBt7
xXGPQayK3dwbeYUjo7x+h47EyTvyKeF4nneaRUmo6mH/K9KC0ZuOpGEm+jYx
1yat+R3Y5ujROgya6LzaPjse65lPssA8OLfTnU4O7vbjaGY5dZQaoMp2yvWl
3P992tNNK+Jj17j+2phJph/GB0tNT7BLXskXOCsSpvccVHj7Bu60vAwn0lVC
K9vckSPcbjGdqqpYOXJ2r1nR3ezwAhyGnBJk0SZh9kcaD74JWMxRi4CVt8cj
04Ne2wIb38HiEVWxbs2NsttB6X01WA8hxTkKn5aKMJZoFztkfWaAcr8z39Fw
EcUDJxG0vev2bQ0kuh2JVrYSJb6DRjUVMv/aNSkhHSAmcwCBw6DB1LImV+gi
cOxGIsE3ywrhQK9LaVUbtzg2vevPsind/71/MxUvsWn9112SG1vvXmuWDOY5
nuiOi43/HvkjnFGJ1ZQM+vvanRJ6b6Ifgjm5Nh87501omitUZ7hchltgyI0O
6wQi0MhiqImt83q9gC0aZvLduHq6LiB3M79ACN34WTdxIVNn3F4xI7RQGdde
OZ6j6nR2fcTC6EbCr+19EOska5lFM8wyI8CmWaKR3iyF4x+li+840U5HK7gl
CXqEufIC4QZfgHBTaZcsZ1Fd+UqgTzUv85yf7xMebJeMkTHlSHkPJ33lckdL
ctsHjnEGcc2OG26F1c+4bEcMFiFbdbme8vIQgAj1hJnbB8anuXIAz9aNTVcx
o8jyjiajYwyVCC3vlDEsEont59ZxoPDPQ7jeanO5bYXm+iSlwcKugxPg2U4s
qAs0LZ5SZ6SsYx1txcAWvbAe6G2+bQq3GFgdP3DBQeoDiLefso0iGwvb08Yx
Bg+GSJJbf12VdEOfQsNR/AeEBoJ+Kp89gMKdz+LPqFjEqxl6PSjy44GpnrHb
B2WzxWcRrSjozYg0DXltWHPJhZzwgOu0Ub452ebvgZIaZ9G/CPrJ+eqE0Kol
XrS7LdnKFnZuBWB4TIbtOaCcO7Y/KbRsu8xSi/meGoegIbQeM/+Al04pRiax
8871N8i2M1jHbb7VSwSUt4uM063YTyOgHSWiLmoqy2EVYsK/reUsVPlfqKNE
kTgIWnHzOUOihGiE6o7bEK+yHYiNYl8nWjSJc8EW+SpD08vOhIxd/FwuST3J
Dk4qSHTI6I6QZ2eSD0wMWH1SxFfL/40be1EdREhGUic5ujKrLtav47Lqvl55
JVbE4U/8/ytVA5vcEHy7UJ6YatAz0+wlFfOhzfKzk1enFE151VYM/gFAdtgf
f4y367L/0jRLuAcalkPGmXEph51WGj1zX1II3BsEKR6ekVmGMxY5n4A7X9W6
v9dDfGQ44SNis0I7hcDRpaAjAw8o0xUu9wAPpGlPrBiZVbaSHmJSY50gpuhU
ateS1SLw/dgeVKKw8Ro3HJgrdwz8Klmjbh6MA8JN1NJIq3Xb3QFO7jHMvgzi
TSNmOc4n834KEMm3UwaTReYLr5C4EtG6PEOyOo0xm5qMEqWC0s6kv/3YUnEj
JAIeJcWRKxqnzDFmAyEnExJ/p+1YbbjMf/x73iUhLLoEXyatfNmJo/XPFxzw
8kkqlUvaYayEzMcWEzUt0578lCvT5FZ/Z0hf+9mNnrRWk97GEWqDZ0k/9zJ7
NfOW8HkWALQPxaPJLUFftNxDaeaa53pzPWmlp3lKfRsGifOO4mfbQ8Mf4qDI
7NIHyHOmrHbrIzocYmq760VcZm7hpmkNsef0plVIs/PR/a0raZ48nlwotITn
5gkQVL1ESFCAqRcLuWkZjmMu/t2itTmX5YDxCGSsTg+vYyMcTfAdwgAUXz0K
N3+5ywyU1YYuuGdh7CR++xtGU6A2QP4887iP7fcUc66e5wK3WK3UQWytJ0BE
+4VVrCOORXytesaS00JIHrJBWu57DJ3JwLFsn6MtkCURShQh0BU5sJx9TyDZ
pNJ3oaVc9UBNVlZBog8+jzsOAoB9/qt/4GzdlxnaA8I0LNPRvo/Fn5YiBuvA
SF6dPJfoU5Yr8td17GH9TM++ccFLwLGurlb+kym074eNu8S91WulZtTIATeG
ZnD8pqzcisSI19/MJrVDkZXI2zjp3amKXW+xyFAsrz6arkakfhjBw4T67l6y
qrvBwh2ei1TT9WtLrSdq1XcbbbzibEJ+uq1dM0BV9ZaaEVKaMwIj8poOl8QX
MzzTca/9dTJ5qabmNPc4pF3wScnR+QDsXOop93+3mFi/K6iteEYGuLu8baOp
c7j099x9nvFs2JmGB6UhkG+rLkDdjy+oEDvYnDZklCb5n0pXM2pcX/CIptsW
Z98/VcU6oLQjyUXPfyVfzWii6wLs+JRl6CXjMAgBhAwsQyscNdYJbv1FUQMU
aAJg89GqTJGOxqji4/YJokMmSXQVywB+KQQ2oyY8+IyWbF9LEWpBdpJBq24f
3evazcqWSWYUlC0kPYFsz3yfJmbBKKOr+KVQiRxuY7L8syqf/PaZn233uc40
IGa36+z4KR67zhrxIg5fVuUZhFZ4lxNmC5cIeODf0V7XzpZT2i1YMtgKO5EZ
o7IU0xlC7hVIFMoLn6orT2/mliN80k45QWCDtY6l0FmIeFbVSh0ey5FqhmmZ
GizJQ/3NL80pxMNBNx0wV2fwXHvuOTh8AmEQrIw/APVu5dClp7lrosISUvjj
HQ1qHK1/pyCqDciSVHQIt4wILcLPd4D0YLuNu4LKFaZHMaboQqsAm1Rmwjr/
65rl9JjS1QzoiLgl0FFajyf+huPxw1SgwrZzcsMJZXxMAGAIAn96VMOu6LXN
81uwrexLxs/w1hcmRhpiPeP3JaMSYYIaZCmepEDvNxjkurNTksioQiPk3HWA
q7siFHRNACwR4J4Lsn6kPPQ2oO3d/YqF8chE7bEAOtLyhicmJ5B0b6X8xavq
BrfU2DxEwf0/+epRLiSUrc0Qcnj2dKx/5FPNKLQxeP1HKWHXrPagE/Cleo9i
NtE+rlaFUmPKAVvPp2jPoqJF4sXEBzk5GUy0Rrk3842UR2HLzJJLIBa2b2xU
1j0b/X7DRq3wLptA2OKiDS+SoN5q0o54t5KkLkIKmwpRORJkYM0f8KgBDetC
38p5KNsXZzgZBFp5c7YEbNrpeYMpurQhQnKyd3/nAECjnqHMR7Ii2UIEci11
iKBhwqfYkDYqmhR1HZiv3kHJbQRYxKb9ybcnqDIrG+iQuZRhoDW09U2kyiSJ
Yko5+NRn54YA4ys5Vn5Y4PBbBQpYtDf/MKvDWBaZbLvpKSTzOlmX1gqiBMsp
Q4GbmCdbcikSiATq4+6mfaOpi80YRauszpg9Sm2U8u3HR3YkHMTJ2uuAv7Kd
JxAfiaJwIns9Ns+7YMsrslwWIGde46QEXmM3dOilZV7uo/ix9SGKPbgz82uD
8m+AiqmVCLDumI5ix/BjmxfU4/7lcG+p+dEl/MJ3MRu4IUOjMgEiBi9povUN
ipjeL9hgU9gl/E+gou694ORJ6LPEevpxlmqE/yPkD1QpPBH01dV+oaeJtCLz
kOolSZwMJp1+4zuT4/fkqw+5SkTdx6hAC7Xo+od/H2I6BFUAIBrdw1UzuXOW
JNJo59B7EmDpoUVvPSinXW0zUfh7EJqlchOmPEY1Nb4DTIk+S0yQBLz2CPhI
FHCIac4pFeyqq1n514D3W3Eb/uz/OWdeGjf4ARNdKJcyxlsTQk16DYnaesBC
u0+msUFG2E8M30VYflaRexRw9Ji0sFw0jxOD+dzxEo/NCjoZd/TJzuM/Gsrc
9nEfhUyXyzZ/nGbXuqWtPGj2ZPjVgJYQ+OIW7YXAyE+9HXguC8Z6JKls+YXl
HgB9mhAk/32rbHZ4X/eaJawaHeB363n0dxuzYUDdr5fIqrnnNYxSoLrPcX7o
Y5lUF9YvF5maCUt9oMX+PTGLD81Bw8T7uiPvOmH/VyYo9LY1c3iSeP0JWXyW
gSU2BT4cRPlQLydnSH9Dics7mD2VLYYNjTONhHr2P/eaHBiNP0nGJckVqPfb
gXBvg2AVVLuI1lvGu6MjA0BXshm3N+AUC/Y7htw/aZsqGBjR4URJysaOyjwQ
jJowZtWclY3EUQz76s5CmuHDB18qGoiD7vPDWFHKK8ksMZVumiU2g5RpT37H
S/0PrV1AkQdop6BZOo++uKxLJmF4Uo/0k7Ue1lJoJAxIrGrjnp8XCc6hywuH
iqV/GXZX5ccSz0FDsmBNN4w70hFmW/CDxvgMgbcIKalbMwXweRVjMPo4q3kZ
Bguk9Me0wa6Il5FZ4H0NaqiVCk02df3h5XmdSe3wI39ETIoR+K0L0VhbbFTY
jaMM9F2gEGni4HJEJEa+aVjnJm6hp5rD8JL5MPl8K+ByiXsWm4/qskAnOxdl
bAs7sBJ9SbQQttIQR65Doo9qvcP2IliaXidhAkKHgiROAHEmIth8EodHL7bt
igRBfKaAdCoDfR354fQiXpnAOCE1n0q1GiJ6nSuLD3i3JuH31QLmIALuWbpd
xL0rF7RSrwoZjUNt3QQkuHwnoaxfDY5j4i6wd0ww6Mv2xk+cACj3W4CASAo3
U4ymzy+yBK6U5PmFwcmYUAfOvRYSAIXIcy8UnQtaYONtL2UN1wtCxA3oKbm2
QImFogJIMh3PVweAt0BvszMNmJcSorzmzt8o+tUCwTSxKRxVXqjRGxkI8cMz
0ww9awI6lmq2AbGGYSnMIKLr+EWXcVLzKheHTcUPdgeFPUq0SOfq86aKWJTc
RoHVUVKg79ayLsajMOWX870mXuZgWZNb+repQBnULHCqdfSXoHtsDoKlGume
Zim7Mqoj0WvJgZCm2hxDjE6z/GGwPZ7h0FMuYl78+GmXgmQu9cGMlkeNIn5e
qRtlxm9/LsPejKa4KGPiPbigW6BWVcQwI5jWXMpeTIEcaRCePk+TqjJ+5Z3l
m5uAKpZHPi1mLZsQ7xg79T4plSuNqTh6pDU9pWm1mUFJ8IKQ6IJT96O5gcrD
fjTvOKA1OIOlL0+x8ogDgOP/3bj2lRybfF5DaoKLjfZdPaP4rA4QviraHCpb
/LL1AOZTZfMDZ6FTFhCalUou+21XWUc7O0rWdR99+bVBEk/rVnMK5zP3aSKR
MJTmA9QhI5vuFC0Y4tRO3hs71woII2Y+aH2R4fhBJ+0YsKoi4CFaKQSl31yj
2gKeFjMjVoDPOg1AdsNCqsHa94EPAe3LO2qvKFarDMVQVWoiv5hfEAy+fR1J
efByPT6KldBzJdsCGKA8uN2dDHp6bkkYmA/jHePuGxHk4XsKdSqDY2qAPkNC
Gi34dQkw6VQPMb7/iB/mvk7BVBWoAKrWbRjzbaXF9GJsH9OtbEGNqvGKsu1J
YSZKk67ANP1F301zVt5suZp/YCDWDxaCmM8absTscwo2f8HlFIhSOdlDrsbU
eu2GYXr39vvdBAkC094w85BsAN/qgLY+55ZyNgI8mtUe02GEqZwj5D/kXEsN
M6Y1BQrH8UOd/wzqyleSeG1OYxPpuviWPwKcW6F7m8onptGm4BcwCF5eAo2A
5BuXRFLN/0/kLXLR4jOuJsJLaF6ycVtrbUNFNwwO9BoGQJxC1yO2SKQrSnrN
tLRaBv7a8xDnASmWEI0y88wsVyOFD7YO1yBeM/MhEjH2Yl6T6WiCI2glCLpu
oPRyWby5+Kpgwzp0VDDmkZJMeWGMadCqR8h6ZPiwaV25uHQRVjkimPzDAqjh
pYqoRlFexJgt7GcT1Tr9LxztOkjYx22K2P7uJuIDCiVviTPft7HK0i/6DrdC
CZjbhxBH/19ze1yCrMkVMQbXllPvIOpGQnJPAveFpYrsG8lkKTI8ruuryObu
A88OnUef7uTPogwxVTChDvq5wxnmPFcQBuAhJ10nbOHrhhZ0f84QCgeP+b8c
Jr4Xs591O8fRRzapBzAzQl6KJr2e/dV4Erg2so7fvYmpuBCoDPhbVbp3ZDe6
PYc3t/H7wipNc4T99IPd4mO6nruvebdTMxqZQeVuJNW+MyDgl7Qjh2SqOLDa
9RtNAcvJDLZciTuhyYUsQSRLBRFtNpC1Apv9GPF5LEP/2S3C6fPdju9i/W5i
Guqv72n0gzF2YGWgEOJNLLjZ0cblzxg6RSOXquWZ90LTPKl1kwwi22a5L6FS
lq9px8QqIXIVC34PB99G8/VZ0//yp5DEjZNS5eHUb6GEQhdnC4kij5vnThBN
jDMkmzRdWhELroeH33/2XTG7lKNsSGgkxqAG8HT2jsBXsCkPsdgGO0eITnQH
vnNt9m2Jym2cLmHusIx9xS2qO1NmhmQ3XbFXlvHhbZeIoz2DM4/9h0YnFsxT
vNMxUVvuyjuTxio4Q8FcAG/YsaFqMZgevu3msGGmbr4cpsxta/Tp35M1PgtQ
dPz6l8S/Ibw/18q56m663EiM/7Gwc2fD4zUEC07tiTEBwUsijeyj4+HsYhe6
EA0VB6STAOEm36YR48p89TGZE8Xgei6+wWxNXsDdSIcUNWIa0ZaiAAg0eyoM
d4tf1QYC1ggtM+AbpZ+psf1V6rBYaUIeKqa+CB+JyJh88GrWrIk6m9egWxyO
n45ix8kp6eAQGSDIDuJsdJrKU8XFri50g/P3iqKZ10WGpUkWoxraFDQnLAgc
4KM3skoGKnpyu4CohJGGy2ITfX7tQkBeDR1pe7kYIDk0Gg8M8JNlhNP1hfit
9xM0Hk8AB8LwndRgUH1+zKem+pkfyr6fks2sA1I3zwP71rFCPX9lliO9Vt+e
cxOa0DRhK+Ft5/1FfxTOSOJRVFqLJD765IHXZySWWAURYrMTM0JVqQdXdxq2
gpd/yPWxg6osQg5H8+uZoqxvPPq9S0LtV3d/N8yr1/EPDts3pJg3J1GBuEJq
tGICm8KYidqN9b89bmRSbs3QNKGiHtpYYIv+0DdO6WwkaKiFtKgU01cKFeLv
3Nx41rW4JEBDtj8p1Ou/14RJ4myLpMQt6UTShZg0b55rFr3AOKtbCR6k3AqM
bvepZWySX79W5s5JNtIaQzM79bEdh/jpJvBpymykovoeuOrhwmrbGPNIKaKV
E7AGTHd6jdInIoCXuThmzZoMsB6anlPhVZX7VCCA2KF6lkGAGcLF6Qw9C21H
FY3WRM9oU00/vEh3y93xrRlFWn5Sb8LpCgulDVOBnRNuXb41cRDIIMZA0ZgV
vp/PXoPrbtMpFPhTznara78PC6t16XBiNagr1YA9uMQYiEFt/NKm6mm09G4D
A2AuxBzoPa7nt8Ye1OTULewgNi5pq1Zm5KsOm8ymOTlyKeczc1/07HZExTue
DcD8dZrtx8pOF1FlXAt9XoazC06PR/NFvsAfN14BuB1y40mHjT+Dontb6nQW
aLFsOrMFdvJb5VpPGFl22rARz7S6t7mPI+2i6TC5xXEdJ704lLwTHGMjl3zI
JOxrqPYni/Bzh0ugW8DBwjY43rzfHxh4+hlCbfneF6DYEet3s786Bqc64rO8
T3uQuA3EY9w0Ee4o0OqpK3LSUkUvlu+RQpAW6bGYlS92L4kBcWifVTOGiQBT
TW6cssgpjBLMm2vOhXTGgT22r8ioMFnaOBimCTMkx9R6upWKOo5NK+y/gq0V
OWoQEfh9dy6pjnEpOCgfvuq+T/j/0LKgw2FZBQGfDDx3ONJby36hHEDRlG3n
slEIVfvujJhTHCfIZw9DhyDM0u5hDILcJxN/THj/kFifptOeI294QbsRbLA0
WbG4QtH7/4ND8KzecpIf9vIrKTWCA9FNc7SXmBzCGU0hy91RO/RXfxyo2Wq6
cPJ/Ja34wc3UgcRZ2SgB1CypjGDgqs8U02fgKJWMQG8WgnF2u77toSjzl80v
+kGVJUO2aWZBJtr1DwpPeka2wNtQDkOdu6lhJh7/PDnZgRXMK6slSsxt2Xnx
AF7Cwr56AflmgS/yadeZJXid0gprOr1LhK8AdPexvz3lrN2CoRTrsa02JQbf
h8HFDYeinPdyyKVAUSuEPPVJa0ajgR5k05wtjto7+q9f/TDGfD+/QocnTEmg
HTAi9nSxJhty92ckmYFLewcK4E1q+vYjgfs9eNngLlTiJ/HtXU2n8B/VT9U0
4XttymelSB8FmiSfAuLhxMoyFyTV5/RwIbGSVWGcaCfKpDGMPSQE4Nu7rX4N
OMSsRqm4Vm1WOAx79DC2OE/TCGIQ8tvLvp35BXPMGouEXP3HKFbLOPNEOV6b
B/xvSNhPbs5kVPrPlPFP/6Psu4BQdy10w9K6C4HQdNLYcX992MqUq+oc6iWN
RZr4nTw+1AA/XJJlNjZH0scqwl5y0wFxAhLjbuXg0PkCJrw947BVhmYmJOWC
51A2wFdB7JS7EQa0aXcB8LhSmIBb/49gbjYnspASqz3grcC4GU8mMWPKbvDK
NxaJeZB9vlImaQ7DSB9ystyMGPnBri+7PBkFDUqm1h2pU+iHN7tc0C3/XvXS
ydkipj4YMJGR+1vuRGLbnei+llcq32Fw1KSAEwL+qmrK763xdXZk73fKN2GK
xBGUpQpw/KMGJDUQR47uQQje4VbiNt1op5lkBlQRcgBMaFyT/Sd0a4c9cHfR
p7EGdjxMNLAQWekbleMCIjM74ZwSosOj7pYbWna1FywvCIbAkrhmgEFk6aqo
ZdPgXiY65/jLWE1sOLnkIt08DOaeM4Zix/fjnLPZUcBB3Dnf8SYYw2RF6FM3
Z+VNeQ2Eqv+SfgWvyPWahn056dLpOCF/jI1/DNCfZb8qh6FN9XREySyoFb66
jRRZWlBH4g+KRLQewAXsFqanEOYWcg2BAHnQizxFLf1kl1lpZgYuBRhY5j89
MaCPy7K1rkiAyT8Zll2Q1r2l+Vda88XNJtX5MtI+foZ55mNV/Bur5zUpjFd7
aa1mn3BJ3ZETs1JEyOGytLBMrEJ1nupsyLuwHrlnNg8v4OrMA2KZGIhK98J3
PdirNjk7U8E1X9BBQe6q8PNKz8VoVmDFmbKrr4i+buinK1f+AFmIRixe1ri6
GpXqg0Ta0D1nMMz9hBfP7mZTxuwoySGrZvZRwpFEXfu90X+4Sto4rfBleb3d
Y//EDzhfR4CMx/iL0bdkfC/bYXR0O3/ZxYAa2ukliZZdhAudp3dB5qRV83cp
sgra4+7iP2eV5Mm0DWMGS17ONSCwg1VTx8/fyky+VXnoJnndDGtyx2eXMYoc
FlKqClUd1jpPVn7N+UDgkz8bf+529Wlbkx2FXC67uCjofmnhIzL4nWFG2sFM
C/nORfpGqOsPN5J0oIpjomBk4NUli0Qnqs3ogTYDp89HlKHdSa4wg1JiVhZm
uSlZVJ+CJsb4Lj6oj+ytmxSOnNe6ZHtg9Q7RdAM6AWX9ldE6UKr/LvbtgWmv
Blo6Y0qV73MP5+anaEnaf3t8SMlK2ltexoOKHLxOU2D4pL8UgiKldtWoARRy
w8dMhFtzTecW5rtiDycDCTP4VPSc34Fv8NlvV2Jp1AZ/C7B1DaemrDlrIV/5
MdJNH6ohPdhDZB+2Wan6OkzAySjDyuFGLfLaZjvG3Getf+vcnlibeuTTLU2Q
nZZmO2aNBAgTOVuVUIpYVHRcnbIIr+nlqYS9HZwz/eY/bwrDcd5+1qlgNRKs
f9lXOEbbvt6Gj6PhAHdRDFvcwYEvTnefGV2bhWXhymBRBBgEOMPJJqoaoO4T
RU4yZr3fb431SZ62eF8cfJQGJPrxSS9jN60nVfhGHb4l25EH5/4ufadUPJtk
REqd59cRo2bzOH02I3ghOYgOtEe2/lt5ksKfFNSrw6HYwhOoeudHnd5OrQTv
otCcHhuYkCQJ7aj3APhuCNaXGsxQJF6/l4OlY8KmVh2tUWqHI3hApCkPwOI2
ui5S1EdDpN0/3VUi7OQcgqO9dyVVb33/vxWgsOGjC0dRrJRqE95cYC6zqDwq
gTtM2MhCTRHNcQnQRu9AhHq+cK3apiDJX0EV3TEDRGuOFP+3/Bdr28mn30zD
HSRx7IGJB9qme3t0j1R3iHMXaT50/D5QS3kViWuBU15Eqk0wWgDnbzLE9VZX
MKKof89/GImsWa7hWqUJz9MnrRCdnTM80LXjgPOJ7IxdczXZW5sSXYvJvg8k
L5RcD4NXkFtDLQ5Xgt3NV9CEHmknG8OPVcoiiDq1zqjrDvRHJSrsPy4raEcd
6kD79dXfVcnTdggVfZUCespfhmbF1JMB2BVK6i6ekEFXnqlE5Q0kj+aNMF1I
/IJ+h0aWgYsl8wAcjPCE45FYAExcRQeG+71cO/9l6rmQqV3shvUgnAS+/NYi
TWWf6QY437o3dep6ljIZYfeE6c0X4AUiw2kQE0IHKrW3rVVlaVXArgpXYT9w
QnFt7yTy12g0AbpNuFpf8lK/dAlU5G8vi8/us4MKVi4b0Ylh7pWdbCPk38sD
6GtAEE53ioMAK3GBbSyC8q0zmCE846TRBRMj3pz/NCJpWq47/3jIyN5j/h2z
7jfFQVBjQc6ibNRYGnaTmHk9XqsujU0LFxwevXQTzkhiGyfUoPScDwLCWmCm
qzJGB3ZXCUsHA5rLAGkXvGAeiaK4+OGhTut4ruEMh2HkvNXVVvqjLl/qrXST
7IAo1bScenpXhpPtDXPXWjw/ZOGG1kC/7mAmYsRp94J1pEkoGtgy3W4pnNa8
1yFbpHtX+wOTk67oa2cfIJUug753DTLP1FJjMvkZUS9UNfQ2iXbzbChOZq07
uzXe1cgULlOnyGT53i1gXE9VE1v1097XyUUeqfvXIKg3GyrGVxo/DcqO5mfg
HIfAOQxudLaE+F2x8nD7CdgAKFoSpVYESALw8YhQLoFJPFd/FtWrybz/osfL
ettFT0v9bKiVW6ZfIyjOR37TsmaXYVZGAvzoD+xHN6c/48sDLgS3MRGR/Y7j
JRmHzoNg8Ur3FWNaezGC/dQ+a6nSoi+/kiZCFmFQUpZpQrQ6jdb8h2vb3gT2
GD9/c9YuD7g1JLMdScBwMbS30SVVzYdRzkkiCJa3+tsJcmjmgLbVnjsU1rAb
VBa7gEOcE/ORI6SMvuyNQZmG9SnR3exbI8sZ5+hJHtKfmqy4tOU/URhPTVsk
Iyzsp9wRCirMvRwrzmPz0TtmaN+cMDd9PRKdEh4kVqFLnuqkWjbYDS0oszpT
vG9dAyAuUKjpXOcSGUbNUgwu12y5skTFbwOGa7vfPSjNyKhSudsUF5YOaWnu
RQaSi/QsVzTHuOxoCL0wHnjmhu1YwmSR5tvKn0GR/lkiGRZ9OB7fqbLrzG8c
QOT2ThFReT1sypo3FfMNc0QnxqDGsO3UBIzeY7oOE7dVOjVmlAEBNk7e2iWJ
DBftEF2N+sulrkNQdh6xv/1BmAC7lTyfzdUfay8eJXJGlq3eoZbjpb3KdDJQ
AYoO+5v/SLm91OMPziVqkjnzyysBukbvKKTEJ67OLP8Ci17NKcAHOaxKX7Qc
hQnKzoiAPwZ+3uAGtFGhxQyYkMxjrv815fUU2CTvTT4vHYzakFJXKQLm0rt/
FRYWltUTp9oKbLnF6XRKetXMOZX6+9epDEn7441MA2WxnBSzJTI3N+amw555
RyjnPSQyDVjZMnT835Z+8lifrf3byY5v9IbcJGelt4V43mOX3wf5TFLa1UGl
/+xUoBC2XtbJG4tj8uLI+cuVliqbX6xhWyVenOnjGrtGKqKo61N9hB0IyvOc
PW3VzhVKl26iAGk4leDj4B+Y5kp0PdP3d3VMzYPZ2VTCpprCbKkSnDBxwkZF
UBRVcBOnMYC1ReMfmabkuNvoUdGWVVQL3N8XZBB/47u3try/zddd3H2lBz3o
feuM/UV3kbocBnmjYVwAgZLMbNiRneuOz1Z4ZUy/IPXy/NI1F/+5CpmC65lI
Oko3mXpdhuWieFCHiNidIjKOARzhiet+yW6d0G2xfcWevQhUMC5/z7IAAGeV
5FBKg3PdZFqRoBfPK/7tIH/rT3Df+YVcBk0pLOFhY1rrOYDKTG/0uxip2ZwJ
foHeGf4JT/Y6PnLjXf/v0H3I4SeMqYEZneXDMd7phUKWEmIRI0fsp8WDTSwC
dOSNNzYhzWElkgkNAqf+IC9FIcBEhwHaiQYL7A666KlgfmUUW5RaGSHednTw
wkepL472u3aAJjhh8nfgGG9nuIQd8NlvqMkiHRChDLXrA07XrxjdibP7+HTU
4JEnIh4GlK6cCgVFb6xp7RoYsD9uZuSukSwTluinI+zdwGPnns+nwqMYqR3S
nlynEVJezpoG8WS6gGu9jA5uFC8MRP25GUmm0D94BKIW26Srn2MmcplaC67e
hgNCkmyqvYEWGmyPuma1kYL5Qw9i02i94q/vCDN6Cum1Mm3Y/MhKc9HxUHHt
P+Sm/TyQzkk2c/2KtsEQhN2t5rObDHijl6jt5yEBUJAxJrcFvp8zhGjeC0+P
750nBFVEm1e3RMgZc5uVIJELoqWOqnhwqvKY9EqSCiaKcN7o+FoE0+ivA43M
JDo8WVvTD4NVKemnzIACRCTMsYHXbkMW+Rr+2OESwWf9izEwIzsPvrTCT2vI
cOAnlEF/dDxchCvFCFSYwiwZ3EsqVSwL91518LGRSgoujxwL1tA5sMmvF/zw
eV+D6ug90APbP4TJozDK1RCSwyhh6rVIDMgt7MurzmfK7D0cn9Zmz85aS0/Y
PhbcS/07ubhAH8UYypNyRVFBhg+Q6l4H1OBOFbR1v//NxTbaCPbZQZ/v8PUD
24IB4kQqRzPzW58yKsv6ow6jcfJl/Nrd6+z1THl2jM0X6oSV1E262aOCDXgh
l+DUHFUg1e54QjgUeBZWYsthJDTzpBEAGqPeto5Dl0dmihtTJTqZyFOgBR+V
TAEq7gZq4bKLrDK+0cWuKOqOd3hHApRGP/DBNXuHjbEK16WjHYGp3SkH/1Id
J2o2x1fotUj3XGIlpSwugV90CbfiMkJLHYSzl3ftaPHPtHisFK6ZduiQrMa6
nXHrdw8pKt1aEdMXIsARkIIvo97M0ju1n+YN4/0wQCFvOVeW5TD8nQ3O2NH+
VASDWcT+a7ULnNPuXSk1YikMvpF6di7imrHTsdT7KwcFflRuan1bzkIRaOKs
3ox+DkNT6QDlBLYTnsHsCn0zJGR97hwy5Sooli5f1zqViPCLShQm8Og4Lklb
pbakWmTBgv8IjovcKepsmjHgjwT4OpGf5VIywuHoHKLtL6HD6t+L30touJeI
xDsce9TY7pGlRHoPxviAwCrtZtV5UczjG2X3R+oSpklpZEKxYKDLh2b+w7+5
4CPEyeCRKd0813GvTNj7unwkiQavo9cOpKDpqiY8RNaQZemgjnxtbZiWOh2O
6GDvbfITzmKyJCZI5vuGllrTD6Dd0a7cdORTzjnaKmi7KGtDzQnSs3ymug8l
Vb6erCPekeoaGGLU84eUloAI2CqcDvzaQi/T0sRdXqqzjUAq5yqeSr8Ky/mM
u9PRoZqK+jfKCYHlR3ZtsQ+rLdK70cRgYgF0dTZKnz5XR34B8PkOVY6ND43L
90egOrIhiIklqnpjx7fOlk0Y2gmmYypYtz4bkP76Q7WIdVHnEjUZzO7Z/Jq7
IRMrT5SSNozA+DnBnKaIev6LBEaeUrPn17cdjq8JF+yKXuyMKmrqBFGABU+i
zKe8CpdLQfT2SDnpo3lQFQFcmSx7C23OMEHWOTfRuoJF5a/UHqmzwT7OXNKE
7JzMc7Hfe7derDpzXR72wKtMeUXHvQ3z7UujqHSnWVjsCEeMeN4+od9l3/+r
krrDFbgXp4XXJrFrwKrRSGDMQZ8fugzafOgu88s9I0Ggb5NdvvToxfVY5ZET
q5UXdrtg/iqmS4qQAGQLdjv0XQFqXAVMDNOZwI+8qQP2Ust0oCOZgPhdoN2v
BrJ0rQHm2zOGK0rh6EZ64L1QXYTDgXUDm5A+2XoqwdeATXwGm+l7oRFuJLvo
g/kp91RmRj+1boB0g0pGtuxtVPwtq2atzlpkCRewPZHQgzfvCZx1ouRTH8Hg
rETmnywBzsBGKYxofZv0rVwcUZ3m9bjjOxzRa8dRJ8TzICSycMtBF9u+D91y
+D/Egbds5IezhwbOtbTI/nSEsH2WKKHApA8n33RTvHYDaxUO0pXm3g/kBYHm
ODOk5nISSFWQuFaYaNA/GAgFDEKKMZzTilbwQ8b75QkMncQkUe5CuXB6xTxj
t1TN8AMrwdS8007GOE0WFbmrAnfmPvYQvkQh6QSxT6a9F57o3wHUoAYX6qSj
aJZtV6KMyRZS9LA7oQdEk9VHdiUNn1BqGCtUKmF0VWiPu+MHxsrzPakbyW0a
Q4q8ycPqh1DyUiDJd2WZgjhAnTLYrPj3EgzHZ2cVWCCqyRjDo+rYk0fwJS+a
Whwc/9pal2gb8WJ7h+83Qheh3nVSYmyEojs9fvQWE9eKcSiqXoLn7J68Z95G
AxrUjEWB9PICoY7iKnRhvGxJsWFkSRNYapuAMAux516weLd7HBeKUXXz70yZ
T7c1f1TKzy0agcKVd8zjKxbc4ToIbFkkMAUvUDF9UEPKghI1ftV84C0io33Q
jJG7qYhw1aqyL/ohaB3Kdm48OnzUeeRON0Ewj2KWWRUp2L8pN4r2UyjcJ7cV
HUo5IxWnkMmbZUAqHORzL9bjlaSn+M1OJO+iE+hMfRwBmtqqIjLmRCipnBNc
oSfUePqqQPmxTdnP3eiCOu1UrGEhX8h2gZpmSd2GLA3He4gQUuLJo0Vu3oIQ
LNxFFH1PrYLpslcJJPTw5cUSKi2ntezdikLP5SIch7H6QcUO7iDswIM+YhZs
uBF7l2R9BzGEYVwYjuBe4VnZfXZGsy63Ad7V6I20O1jlBGqm82mS8wI5TI5N
5nLFLy1bL+izjZB+6/hTukr4ypSX/GGidiitN7bxSFMcafGHJE+sS+mNsDzm
yHiqt6MG5G8X5aJBaG1yT42uyX6L18tp4WOpZ4pMT2o/X4FKr8twaTfWackt
TfCrXvi+yCWFWGJ3IXYaQc+kuLalTgQiMkQuwd7xzbPx54Dxtne8ANY1a5Q2
VtNGCAjXv8DYI1wFip6M1DISlnEqEXxZeodxCof2jwuT/a1fL/1DhqQcm97u
2J2/bX387bmvKZrREee1dpUf+FtB+2kHisQhOxi0JlJB3st6ObVk7KBFE0aH
8HY9hO15O1/sgVjZPD3unYuzwm9fAMRBG11ZOb8Mm+smFHmAvSh17aL9W/c9
cUMOsOQN1KJJ/CQwCpIk6fjKtArgAHvKxoTEGtzrTU1fmGJhHgyv6noetkhb
7yYoi2kJ/vgGS++rpkHpo1jqivL2DXz6mK7B9EhZ79q+WMrLWzz35AeX5l5Q
q9yZmw/jB/C+n849s3IJ59AhSePRjrNYruWadr+M8EaW0SgCXbgceFPmLqQq
g0obVlf6Elns5chTKpGCvX05FKPueHoe8QzR40lRb6hk2bux5YsjNhJ8du5v
Ew0lW+r/86Hkd2caY8YvPv2XtsSz4UkO1CFNHewJg8LSm5srchuO4Mnw1mMM
i3V7nNzzNyL+An+HfvIO0etZUbzADr+214fHJIpiE3T42Kbk1RCr2DAuQ6V5
IWE0/y62CJc02YwIe9ydh/fUGVDcAvEWFBYYWK8mW8saC0cORS4bGOaZDeWA
nnG14H3iGUiQlku1TYQZj04ISvCwcHwyN/Fmr4demmCgOe5QDRyBxs1/sC42
pDaaHzHx2IG9HdIMxBCLdaVABdwHCq71RvXwfvV6UjeJ35Z1+A6dwlF0Ejdt
KVtLyCaWbAFgZKm5IrHQDKuWh+kdmOZPGYHHrrSyYpLX8/uWueG39BZOZMyW
mKsIPoRiEDqVPAVeGZYPjg6iaDYMdjYLKfAMO4OhpeCBgnr1r04O29CA4LVc
/m/E2ja6XJSFltPQKM1Y3Hua4pgPwrBt8oGY09/feUzvMe+BS62Ix8BS5xLG
+a2lzUsg5lsue06QoiB0NRoARPi7u8bZRXx5tL3rZvwvBvulDDiJncyq4mY/
RImCr2Z3TU4Z8jduKK96MtLcUXJG9NZBzf4XLTNM54YCWTxpqXU34YQ9+6Hk
XISj9DlXBmPG628LWgBAT0SDnxkOAM51KwMU4+lNnrS5tQEXoR157s6NPtZ0
NS3So/Nn36SAcYZZ4aFLBJBhilrv3twCzRoUbDZBCddzj2+pNGJDWeUnxsOs
IjvSNKoVJ9LbOm8iZL7j6JzGmkDDH+DSv/+Jmt87NpLer3fu+k1YgOJ9Dv6z
4yIeEzstVUClzZkPoW7QCpb1qNU3hvGe7IeRkSFBPpYCRAiikar4kEHkDMEE
0bxt1n4WZwlxdbJ4l0Fncmo0Y95vl2MOXwX93KvmE/g9Esw1p5dYg+LN31ct
LkjisFMhkID8s3T5QTvrMrWqI8SfYteEt6TJVSnUSs5uG8PWQrXdZs13LRtg
P5WDxnNBCgLYehsvjDav9VfymzK/zskG7iOS9Vq/IG3z8vCH3qEtxnZZG1x5
eIxVRPLZpSX2x0LQUEIvOvwUo84TAPqhzj48Z2PYTQrvtvn8eaj+9cCMfNkY
0mp+Tz1VjOcWKxifooyAaLuw8qa2oP3d52ehHNEXbGft7fnwtpJiec3Dvql7
r4wkEkYxA02B/R/Q40kiyF8sy9ornUSToAkFOfvc6YgMwo+sGc0QmwCH2XUb
PeTZwScBC1/LlIPvbRKJ5iS7enC5bUNUCueJAn9amHInDiAc6llPG6OC6Fzn
69tvD9o8iIEeQ/6Y9nRIQxFpeRzNTnAiBzBSonp5Uusd3aIZU4aDuxbCcrJo
zrNhDRU90prljXrLbpyKND+gcfLpJ1sFcXFD9MRmd/Zkdn8vcnZoPU0MZNCH
VhhVYJcJ4VbhAeH3g32NRUL5aeW1S1h9FvSU5Vp9TOj3gGkM+B46nQj8lk+N
JlUXZQiXxoPY9uEnqY91PwmJQiAQAQe1WIBGyhIg1+ZJeypSm8FxB4NJ1xae
5O4JFVeRin+ZE/OotZHVhGaxPsOxpOILWBv+62gIU10KlqNR3sxH6BfnWZS1
u7okSf+wX3Ud5r7TUENQB/PPVXnTzppPunOV8oAPjHKTN4UAucerIXCgSsUS
J1ZXB2Ejxz30EkHMa2SaUKWgc9gP/BFUJK2KDNwInmvPTOnvSiQkB9pvRiI0
GNHoTMaFPFUlh+k2VVK0tvafaqlGtRmRyE1ghDKIRYQkwFYay+hrEWuYWZZS
6eqdi7OFsIlm0yD2skn7rA+Nsx/znHBFq2o+gLP9tOR/5woHhdkq9ie4sKD3
izRk8Zvu/D08TwEiuaET4M65CSg3rCrxtcCbNIfLOo254lLIYl83HFzi4IhT
lrBai2mV7numV3wpEa664BeqDwpgOXtI1KsKL7FNTfEpdeJnlYbr5nb0bJxV
3Vi9O85cd75TDMpuoOztmQUmBA77m5zyrq9292ZfiXy1EG1UE8VN/abNVYXn
cu7eCkfYXEpZAZmMA2Bwscw6IN0cSBl7iRdIykO2rh8zjLPaEHxkNgqroDDa
zzf6wpZw71w8KJTHrwewmOjDj3IIVWGE9srAQF+EpBfNLwzfHPRN7lzm96CK
kY9LGg7mYCjjLrjYs86kotQTxK+bJnv922609H83jym5is0gKlmuTxHUSkiR
QRtkNjHyNlp5rK1K9+x59HXIJfLaKPnLeuZPPX1/S479IB/yEP3gbWxwvHd0
Ml8jwMAA+rzsKNDN+ZB6xpAtxuZQoJmrDnfGlwD5OCCZJsCX1q1wtkx5c7Nn
R3U/ZBOF9jEICwgVWvess+ByfYFCraUmC5KhkgnSobLReyXYNXVT4MXTgfI4
C7KOMV63fVzAipKVx81+FlOlmcLpc3cXEJKJvNsu/V7+SqQbVkXlFrD/rIJ0
l6N0z8ARQJlZGcZW27PA+5XPf4tsp6i6wRMRPxM8g+wq8podfMneu4a7PaPy
ZqN7guV7beMwRYgv/otoAHUj/tcxAjKBlxH3QX87/NfwHJzcCX1HLPHtB/7k
pun8TRnmwN51jHi+gWyO7TukjsYN1ZKs/ZGWIvS7XGnuspyuqpODZxKM5HyM
bTVc67Ke0VZPelnbLfMdec/duEp3e0MlI0hBZBa5lvGa7nTfxsJvWciSMxO+
egIAjy7Ej+ZUcATFOvsh5lY3BHgQhD0nlYlm5weeHBLQunM5lr/kcKApKk3A
fyD7vcW6VdfnCXsN94yo336dz5F+K8Ztu52igpRIBeE8ktjekWy/vd5f/wqK
s4HN8OXhAn1v1PD+r2LSeu8EdQo3CY+5ZTxnRSHHUqTk4D9yCp8PC8lt+yIW
zb43DHfKMJ2ZpbgxsQLVbda5Besg0/cm/LZvIOSMbpt3Vo1VCH9z3zqI0NaU
INPvUFtAhKGntHuWSMzqVZctHupahs4exHHgk+wEnfcxMV2p2J9dN3g/YeG2
p+Kljwgw+euh9/u4ktXFBV4Ep0zBdmP57DWd+Lr6mf+z6Q8GB+SUxXZtijec
76CjIqUfS1//+zsuON+Jq2U53D8bwiPdO/6h8vkCSowjClNjOfu1jpHwlsdn
Tg0DCUcJqaIXR7MVCr7P5fLZePg2YbHKj18/oP6jX7SrLkArGbbMT+TzM1p3
J7ERyw5TVk8UJXd7wuiB5VBCz8QQU2v0UNYIP1f/1oRMboo/3zbHX46iN4/l
es5fSVU6ETB4LYwowvu4Xi/h6a5xFpJZr9lcibKuk2PNbLLtHQp+0rTZyr6P
unw6BuCBdy8UpbQ9fB9eNfa7rqwX/7MdQ0SZgL/2QRmfQoFGqKi0VMh6Jayg
yUZ56y6m0q7BRC7F8yctWlNczrZ8M5YdC6/jUc0//JZ1Sxupu5Y2ImeWMIQl
4u/w+BshPYiTnstt1RzgCJzHPJej5jciomaKeIpsn+26pf9/OSMWDyvJRG6V
FqGSZY1Mx3GqVKU++LpGTnHLGduQPsUWvTQaydPOgNm4BRCiD79aIH1SJk3x
3xygLu7VQiIJ8w6Ovc/k/kdgXHipIw/18RdZxf97n5KQZFdG+bwUxjG7AuVg
NwHUE5pK4OgKNFffsoSnpJsF1r1EBDY4m10+bLDX/Oc2EL6j3N7aUvvzxa3C
hEo4IPb6xKQCXVas4mf8/nqER6rAIMfQr8ZCMPZpCZHfPPcnt4Cqd9RccyYS
t9mDb9Ryc9ueajFSuSaUZVpMzWa2ovK1KgRFsr6htWBenZ/uav37XcQHNWa8
+Pd6Wf3anZXMf+R1PdxKecAeb16M3QZcoN+hQ8VjCl5uJ0RO8iatjZL5J3mQ
l3KJN8DWZ/7XUxdjan/05z+uNjOuIoodbFF3gK1WlkqIITEHK32XW2CVhVt6
qLFgodM+2f4SfWAcgokCVYLNzFQ/2GIk4FSqggZXZGswcxsVep8Y0pAY+xUp
62CUlk5t3qBtxa8gQTZnrhHl6klkkPRUswScbL0itoj+KG521s5STmrd7zyp
lNZsY4ZmM2cQSOMcSj6NkuXe+vCmzrxznA3LQFiGkS+dDSqb1QFZ4/PlqW5+
X6MCm1FRLV3QLgnqcLtSNNggVj/EV5pqeEqehjBGjgVFpnUeYmGuUwt72iXm
Y6XtjDndDl4iVRlaxzF8N8fxfzAIDrJQGWx/fTcu7DUyKoM6RPDLFjwUYEvc
lF71etccAPhzxSSaur5vJ8N3TrmC7sePNnbM7z494s6dzatDWYSLKvhy3rx8
rhLh0beZIk2dks7hSsxECkNvkURI0ytl6rIeCb5x5QGdwq6wju2KTczaK1ne
+4NRVEm8uQozoO5jfhvjigxifbBr1mZOEKTmK6wN2HCkBJo1wy6PnzNlYcWT
iqqhCww6ufIqf2QDDBVMnnvoK/X8hDtNAzQaA9vHXRd3OdbnyHbT4dj89fIu
P1AUlUbihupEHzguU7KRp4ZMbZpytB3udqDMjgQRg0Ege5ro5JqqiMGxm/Bo
FqdJ+B68fXYRkMYMzE5JoYzQrA7p+Tq/AgwNw9I1iIvyzvwA4YzcHP5ZFWhi
johj2HjmvSxjMlHdoFaRJwoMTyRwoEC90vZR4UBMuKWu5Qh/pjQX3a9t5i1B
RHMGbUXiHuBzKAsSRmKdTaqOqBZ9aFmKKNXyLU5Ed94nS9UTY2UU1fDLUqp1
O2Is//s0ClY/u/nPz70TWZDhdmzroNSq9EmVxNAMnAozVMaePyJgeQvguX3I
EwxKFYgXKCniRN1JJXW3jdLsTE4QuSZpdgygRA1+FLuv5EkjzmWsIFqj6RC/
/Fj6sXtXTcFOnQMpMSMbznN7WfLwBrKW5CyqHRLc83WLSJOl5D/AwPg+Uwm4
PBaQGxmEdO7eMZw/kLPNY1qRH8GwTDY97SrkBk6vOL616aqp+Da/zKdSukNp
biHxVxi+03xi1wNzjG4GSJXLT4UagJGcjb/45lD3dfWRMEuARWdOse0e6DvQ
c/v8X0SjalzqJOEHIVs6cLYV54asAAE4rbs34DIhjO6bWc6jVY6DRyg4Jnf8
u1NI+pBwFsnfVOoBykhew5QVp1lqIHRm4KZ/GFOEhtyZQwNFX6TqB7zWBm+c
1nojoyaI7fjX1LP5iClMuQxF1OVE2vmzXZjas1ZuS+TbIr1BfMxX+0/TskrN
jM23hJ9GqGSJuQSWGrkNoPrZe19MP2AHnbnr8NdMP0eNg4ZFQXb3hJgel5cc
vzAlxfRZgYuOCH4Za3Zm1C7gH17AShgxX+GbVp82HZRmnrgiW8f/vE/o25LM
SKDsQvwBIz3UgQobZ4TJjxnVKMTIAMf/7vuZ7igO/2r93F1AYCkcxNfASw/8
YlRlri8LxxmYNaOtZ6NsaVErpvKxBqNYQB+Ic+6IPHa38WlwPddNglWx0Vyr
P0GMiiFEtf9ysGak2H4hrg+DK0agA4QtFigFUCGi5IZbJIT7zJyx/ILiyteN
oYj03QmY4BeFcMI/oLMjYlhnKN6+YrhJmJ4MM5gk03mJirE4c7FxdWmdW1AJ
rWAIBxMDDtDlFeMtbGFxSEP9bT1kaiXd2685NWBMjsPi0vaF15o5ouXcQ4cY
hEBTP3bJtMByzJO2LMY9VuBbwMLp14SnFCd2177u+Flgdsvv6CU/SmqWN9+Y
2TAWiNK2pinn8YaKxE3RYJ9dJjntRh8APYB7eRykNpi56Ah1qoLtGG8oPld2
OKCTmjsiLwGHYg1xT8M0Jx8qtYYU4+81gZgQiGtZhYxSp3tiKpU/DrmjQGZk
SVhlRnFTftnYLeeQbr0sXr8a67aem2dtUaIlY7zfP7xRRbrW4Vaihaxjs2iX
Ds4lg1u0WHEdz1n6w6L0sFORw3cTBJbldw7Bx2CE5xyTF3uzRdQCq9P211qJ
971SNv7EiFrDM4dRKQcBocSM17E0aR8Fk73/yld2mj9QDKKwIBwu2lAJwz/A
Zk0ACRMjDDt+aTCyfNEol2ObtHjAE+3/kpHy8X4JWpSgxIH/lVKRpBpfWju0
VGh13nCt6SwcsEKiY8IjWKvaMFSTcHEog5b9ipz17wKD3ZowRBTSzfJkqMhk
FsCdhE0A92hJwnX2X+pfGCYRm1dTKESh6WF2kCIUI/51vrxAzF8U7742W5oh
GZadeQVQjuMx0cJhgHjMwzUghWuIJ/IgASHnikxzIV9QQulIlhnzxy/7cRol
gmYBwF8Y2+XxT7i1QGIETwqSFfnPIy+pOaivUmBR5vkAcI6l1wXg/Krk7Kz9
FkyMJZpj53mvygad42NwjLMpOs8LXsf6AZX1Ib4+ZlI7gad8PcuzdLdHRBNZ
WlQ3Z1uz/jI5Zi7cImCBeFBp/fNV5dBeZYalBjWDrcYBHhjDMp+I1bQ+Fwf9
rkf5jBewABenTF1lfzV3IBOd+xLnSI1LiFKvmp41/xR46ljxhzMUc6eGW6i8
dxN+oQ2J6crshFGstsjTFO+ScAsScxn7b/xEqPWo8ZYXhX4CYhIg5Eel49sz
hQjJLX7YPyS2w66UcLwp5b+lNcG3LiLS7FLXAdVnlALdT/gN0P3+lio4Go1W
OSUJZcd8qrb2r9iVODJeRBtMYukCC+EZVrSmDUAc903AiiDV1U0Q+QEXuigg
ZrGHOSiodm9/dKzFTvFhY4ysms9IkHcKzh4zCdcyNlnlicbzK/kxQSTCt6mI
4A1L8er0tHZJb9K9yJ2U7M7hCd7RrVq2CTFKm8GLbjblvPpsaCbAjzzf6bCE
xANucI/6tlngE6V9pQb+SYimwXP9LV/i39rR/RbLqGekQit1Xv0+5hI528Tt
/XWHULbsUPdjiYAS2HDvAMcdcg+dpCM/JLZaD4i1cFIw1eMEO9Bu1ANw25EC
un7iSjwqrxL5FkyOgt381D5HYD7cqDD++wD5HmuBIDZqtMeAPhNEdKhms0dU
mx4nD1tmIYk3TfVNSsv0jsBPstr1avoQDZnndWqbButQynxNnKopj2SuPMgi
1nJY7be+z5CrsFOuCn10SDK+Dt8UfBnIxybcrUBiqbaNUWAOF2oxeOd1fK5l
O9pJ/5+Fgd0Y9qdqKqZFSOinWEZXyEzdypZOR0qEMwkeMcGyXlP0gpGoTBdq
oZFYxmmdF+fB+tIHW8iLkSAt6++g6IRClO2WtMgncJWJHJrPjIfHopetVF5+
Vj12DJ+gDx2tC+3ogT5MkoN4xpxivoe2PaeHKAySIt3h1uvXKoMbP39nUyvr
0TzBVs/m6U4klQv4JzZ2JZaJg6D0M78kxR41GsbtDCYNLA1wYiAQW1MH0nxV
2tF8GHH06/wf7qOK8aXYV31XSewW9Nybkzv7RdIIoWhqg7YsKw8y8AluMu/6
X001C3y8PpMtuzfxNWzv77F4Ji706qNZ/xy2ipqcZQncnYE5Pdldvt1Vk0cE
51vS58RvdoOYZHtoi5CVdwkh0eC3i/YB/f0PUHJzo1VV5C4hZna3ANzlLZ4v
WddQMAVWHoVOFDrOfTlQNAQDVU32zZFSyECB4s5/ftCfdRR27V+k4bphykEL
OUb0odrItLLJwz8YAJuYVALh/zuzucqrBhdwQJyrVDOVTv3bkzdi9rTR9ure
hPLwvQU3/rZCZWxVjSZKozCiPiLMX8VTW/tW7alrSrjUeWJOjxU51zhsW+pT
OQ48kMFLiV24BoAZNkfXJEW1zPWwqL0U9tYKD2FJWV0qNwsTLcPnn9HLU7pL
fJ7HSot7HOqyUW8H8qtYJIF3bo8kajfSF30gfLDxymmmW1wXrTtayiNfVv25
LgXwgxoi9cI2E7S5J8LthF71+SgNGcthKq++cmcK/sz4gklsqiMI3Fm2JwAb
6C9tuHSIQQPtmindonuaISMoSSnR9L3QhLMnH1FSkro6u/EnuE4KCT13jfto
PoR86Mr5T4nVyXtAuMLn+1h62z0RJsVzJL8WK7YrsAQzLXwQQduM4J9qoy0Y
2vuMpBkovAZeqvSuEpp1VQMrXs3EW2zXgooFlKg1pD9Gzn6f13Lc+6tfgjzS
gwslMfiii5Zgl7H5y2l+erLTsEqcOgSXOooMJjrD29xCrPueuzvxOZPwXSMx
9qLA8d48FcedCVX8Ql7P7gSnlN0mEyDg6y0ptbzFT/EGF5hyeK0BPYxi7nfz
sDy33F3xhSvmh6kGFOcseaNsLIvx/Lk5FmRlbl8JWn+zukDMj6Ti8hs1dMnb
KUWN+tjnzZCyTbnGD3Yt3Im5D3B0JgA9Z90JzkP37Fx0PaikJHVEk7shwo9d
a8bPAtsggUXk69ksBoOgj9K7jLLUYmGlvqjpLMIqgCRPrX/Sl3GWy656QNG9
5QsTlwUb1xNbbyzx9rA7CPB9sqGKnm337Q0l+sVStPfZqzKcOtfQtf7rVVrl
BeoZWW1JGfVsTZTp42+zUxmoA5o6vfHPy2hhCooHzpyifWfvjRGC/yt9A/9B
1PjHhsJ2dubXAGuQ6jkwKjxYl8G6/SmUXQgHAuwBbOrjtNv2t4Xy6jiXgKFg
YdBYAz3EFp4WfTvbDC/NN8bin+ekwdCWZpe1Lv/LKE8IRXpIN+pmo6rhL3Wx
fzWo5clLG7moOxNUhY3C/MdBCYExbwfAWG+C2RT1M9/RNV/ZonGxfRTtoHD/
dlnNDJkGelH/6LH+nPk1GmoYrRogVhRGJOk9uy2ucmYlXdslRIhPWb90vLZx
hlluuDPgoY38bKt2f8CLxBIIG794+H8K72SrIMkxC2wbNbiaTBUFLOFXtbzP
WosQimtB3TlUBl/DWsS9RRpAbLyOsUafGA9RWgx96t7eTmQR3isvumI3tpw/
wvVcpd+oFYrNHheaw/w/wjcjVyLsp5j/dnbFokDhsPVWZCAj/BJKoQZKewrR
NpQ4UjXyDD+oLDa22/aEpdqF9FCiwCqiFGNyIMnB5pWjOMS9mbS9BI5AP3Id
Jquv4giG34zG5KmIqZpOMaDHkh+U33Yd3yLW2jc/2i+zIhaBZHZcaWaa+FUm
Cncv+RnWKg1eYeMQ3Jca43fiGJVz2D2Nbb+efFJD2ewVdNlJUzFZzFARd+0w
AOd57B2B4OvQKmDshEdyYS70ITSQBetTc5tZK+blaPRgjnqMQtSZ3gk6VW7e
HiKt/W+Gvc3EvGuqDyt95ZrJ1PeJzS/AtbJ03MAvMb20ezObwJDjoiUODqwY
o01tp5cV7KYCtRbOVP5G+h0KIpoXACNtJYJqcHFk5lb1W/KnXhfrMGOBSvTe
j15ItyR4upqJFTT9l+TehB7tU4sq0Wbpksa0B9WxJRRNWsuByrjuz4IPA5p6
dZvle7z2PYFyl9CREE4kdcGEfSK4C8ML0D6oAx0Ix3cQd7fhAVyILf5HUyIP
A40CEOJXuuozrspAx7Kdg8OacAaCo5gE6/nvDY7N1F239AwepuXGstQ7Bhit
/r7qLuFk4MuPAZStxEtIJuxHGuTf6dSfo/cqd5/2ppP1J166HMb92PaDTAuJ
CAaa0uEDwCM5LnQUuQAa3KDkX3dVvLenNdmAFQ9kpPLofpcslzbjWN6w4x7P
sNzb65I4QoH3nTcTgbtWVEH5MwRMg6s6HABGrVd3xEg6tRhH3XaofR1wlMZw
O89VAA7OOx92lZy2hGpYnXrEuuK6zf3hUELv+f/xHdUtIViMrXbRK7ent6ts
ZX1b8Qya6/52LuR+2+JWKpEky/7qwnLohuEdXrslRxSklXH7MtSunUWl1fT9
tkuQ7dIdVpjzS85w8FcM5hVJXSXsdwDWK6AdN2U2sYSKZp7kUGfkOoy24eJa
Q9lPnBNNbbvAntvvlVCu9fG56e/n8LClHlkkmVKGSZDbPJWnM5a0+3FGGUvT
BDfwTWk7vwBu/wFktTIuZ6FslwEKN2jcIdUnNXdD+t10Pk90ZZu7xDSU+GQU
TAkonZtijwzakDTEh+qMhaisRNxdtj88BAqQjN9s9LkOCQwgHgEBi80aUIar
UWmAnkAKrP06YZbQqlDgs6fiDxjRJfDGJfQwOYFS06NwU7347TjYiS80Ans8
/hHQQPaoLpzWlmM1GqhN/iX7lLk/C1ViT/Hjz4iLVbDjoZe82rI9nLy0OUou
PbwKTX9+y5/5TgE8RCLEni08xQlyvpgb6QEcVg4P4h+wR/05Doz5FaHRJXMW
yVFOQynDKcwLsI07vewUpDomKILzKUY3la8lLyjdBKFVc34ZSKFhxXMLUh3R
fuDtpHeHhdmLmLPVPOQbEoSG2Ao5cOc1+9JM1VePSSs3cmoeiTskSwTuK4Xg
7EHfd7F+PsvjeeEdqBI+gETv1ezr2Bi9AcSnJrABh7KYumYQhDL87S1gUwA5
HTzuhZVAubX2vug73y1OIxNWzbblvie3JTjXXamjIVypook/I2s2hxNko7AM
WKpWX7Z+H+D/YJM+IxQgEXZ0JPJ9/QGphQ7PXVP63M1WjpmNEsycRYas/YLn
aWoP/9Gz+hMFD8NkrC2PlK8BVC+BNlgxo1XOppgKbD90l4I6zQH1leQjj9j4
3S903hINXKZTigh4rmVoFBebEGS1a5zZeIEkQX46VxnSM6p2nzszrvXDAC4a
D1jzLC9QQgQ4HuvVRXMJdTBFNc72AFg7Nqea7PlR3NIdi18Ll/FRoZL4FUSB
Fnwv1BHduSfhf3yBDWmUwArywUFGAcX2ZuFVwQtVA7JU4eT9bAoEhcSCbUlA
Sg4T1/98/oc4wVnpz2oIKbYA6+IITNqn0f9Ha4lCb8E+IS0J+DRuiYywqu+q
/kCJQexHuOVtfi1J0ZK545yJ344ixtQYxAAJW2Mf0yDd6wee3w32iUy+4prc
xP1eTXg7HtaOjN5ZZ5LeWgqrWfRkHAB/s8KXaAuTpmf0n8YkNwzPy5yPV8TR
AX40jP+YZRn77dHW8Uj5tOL0EyTk4lBlG7xBXMcV5QvIZdvpJ1eeBnWSUBvw
Tt1kD6Ypbxiz9x0rMxtq3g3LgBaG3jMZ6nLvmaOmxL4GKqC8r/8cjzIbPvUW
u7GOy65BBG8IckGDAduSRsHFCKekcR1rVgCz+HHAvMumTPG1GDUrSgwykgU/
k+If0TAjnDtNh6bPHLY5S7BqGohOq7gIF6VLcTkKjRM5TXbNZMyg8mny/8ky
D0W+XNYBzVi/9BdEd6iV5J8r/WJTqoHZEBOZybxNb7K9dtWEZ0NJWYEo563p
hxMBdES05ZaK5jYAIdkhabe4mxu7d18kw8rYzKH/SBzduopdA+Kv899f3GQF
GyaIg+agQ+Pjfc6mC6DxIJGvnZyj6xPQkX36TfHCzB0iyg/Ux7dqd3xkdGG/
rKGMH2OF96gEKYiSHXsZL7KBEAWoyh7mZ0gXQb9wq3uPy7qOC6d+oBUBeJ47
qd3DISVWMyxkGTJGbs09C9IWXQXBoMgV6TKCPLXO9mghVxAmLeXoyIVaH/w4
HWwPLSICLysW53wMMG98fxSzRVw05/HGCJVy1P4Cv2tag8BwCYQoIJCIt7VO
kiQnhHwW/bGeQ7/+0WajCtz2xcntXf4l5VdtZSuv8bNYzfcgJrwvAJ8OlMDo
3EfQ8YsBYpaVviDWAIGag2BLv1Ym0uB4mEoiPYWcduK2yCw7pC5OdABlTsNU
fg3Pr7Q1Fr3fTUs8plPXO5Y6/vQ03sNh6vxssCYkhsdvE54CCFkBKGm6Lisq
aPoK3SZvv7pX8t+pd2gWw38TpgQyDh7R2EmPVwrNT3PbiZpexfvH0xJL67n+
Tqw173LfPwQACyM9QWejCNlHfr0DPJxf82iBfcvOvW0kuy43RJyB6w44I1JA
1C5hBbFhOumxDpgeVVpNPKQDp6UOed7puiHN6G8cntVLflOFiayt38vhY7d0
2/nGcSCPbGGMlTqPlqnYxLFPtmQSHod95Tekiq7HWS5Dj0wmMUMw8ChRJyVb
Nabjc7YRaYcBTsG5NGWR185FJ8ygFDcSGYUhJc5q9uv9gMOC2WIPUnOnjmKK
zCjK2vIUUssXVvTu4so5qGO7Ytsjd6m4ntVBZvP3BrgigxKaSH/5taqfP8NH
VYeDvShUduy0jfS70VbYewObLsZwabv1SPE9OfBiOwS+XpfP4tYI4/NiK60S
JsOHVvpZn6CfdhKzF8e0tXFnGoIWhZNRA7FmWzz7RqN54Yipj0nNIP2Fw7DG
pgS0tX6zk3F2euVbEXW8t3nHX3A8oZgud8ZNx6gt62IhyfNvUZOwmczpxE30
zGmyBHlU/kjSyFIVRE2eWtPVVofuaF7bENpGQAqVSevtBfz/maHzFb4LTBzu
1M+gBsXIGIcvxlAXqFWq1KACXBrIMzYX1ht9BhiM+7m4O8uBufGqGLRluDjw
hGdVJhmQryKr9ICenra13UeRg3hf+vVnhCv8HrLvYStPvDPY3Bp3v4jHL3e5
+RVXg6hsHHIUTbAs4Jy7yQ8kak6Fghpi2ZJmctkqA5WOxhjOGfCpsBeHR60x
0KOyEPW3UpSXcvlVd8CQ7KywpD9QcS7xvSFB/EtXmLdJpCfx6mz85PL4a2f+
YxpWYtbGuzJQ33T950C9GX/RZXN5rrDp2UaVvP97n2+KSoDuro3mWuJojDsV
QLmx7K4usaEcd2pPe83GqqExwgDGo9Ue3RmYvglqeFzLgWstxSUoaMv5Mq10
07O3B42qLBEuya19KYNtmvkx9ntJqB2fg+g3QIEKXySstjoruxvernuIOA7C
E2BpcPHiFmQLaLz9+Oza1NvRZEmW9xPHbqBVB+J9VhkBUlEsZDkkejrf2AnE
4D+irUNxOoxYx2cFPY9aJPGNppTuUuYvh90mOYsfPbT8enzqyYFY3en8HFMX
ncB3CplEnvOJSJiyR+aVQUGPjB0w4ShRipYsUPD8lxjkALIlV7NHkB6F0COa
CU5NcTBAE7xOiuOh4sPAxzR3uwM1UHCv705LibZvFRNQ8grukOeN2IHkbBYp
hXM8bUmWTLF2uYfBuBHgDF8Olt/Qs/pkgRr7UgwQ4Kf7lAkWU3l4KET5u5P3
w338Rax0tCyzfmjHia0irmczs/57kQkIkmDdFZrFklBlgCzmE/mykMg3TCYV
sj0pqCN2PQE3C5om0upmW3g6Tz/SEeKmbQ0pszOn9/02aVf51Zx68cgKPPq4
EWt7boz7kibfI3sppsmEL69knD8EkQM4u+lcDO5rvkjXRWhEHhJuojM8ksiQ
TEGJ0qs9z+Gn78p8uDKorUJ+9DLGCt6Ecgm0O2InR52EONNN88SGxUlJWj2A
H5fAwSliujLh6I+vQw2MNwuoRtKQnWMwjJN1wiajl1AjLDqXZpNCqVOviiWn
qZhJHQoNblTEVFJaDnfElGy115JLXU9NDYktei/6qFQFU7PRzOODNXU2+Ic5
EvlyetU2mHwDDrxzmfbuZwhQVVgVLHwIGOuL/pR9hbQ/XjcJoSSEiyxnLbnU
4MwzUqi1ecrnDG9dEweQqGxhPFatFSIyTvMj/dQ8inaGHd8nNYAQ2KOmrs4i
9ApQOgU+w78LXbfldFU7I8MgTck+UeH/kSTR5iIdaLtJzDEBlElviaoF0S/x
Dw54zRNi0h9oZruhIbfvcSu/tOKR3njcp1eHXriz212mb0j6ECX1/NfUwqyb
81QUVZOmtpjNAEO/Ubg80FbPLmOammGpZNcgrtOT8O8nTvL2/f4sgxtGBZVN
9KZOBu0gXWMss5Vr9r+quzdq4JOPKSQcSCeF8C8iPXLOulDIBc6C7L8cOvRG
ERVY0LJ92QeNRHXpXvD3uS/jR9vnYNQiArdc+eyBtdB4YqlqAy11wHyv6vwP
o3J6kQ1AtShbgyiD52kMDzpQ4dfLV49M7po8UwG/rteDjuxF5MnjWsHKdTkg
ys2gfnONTG/lz/ZgGdUa3KJeHDflFNxuFMzNkmfoqI1NKfFBGBIZRkMZMpkk
NcMsjJcW9eWkHZiZjGsEhbGngM2z30oHbOOzSEzikwwZmBArkLSPYy/E0bu9
ZJh+q6/j+Sw2ZdVaaMkfyT1n6iO8dkJZNUQ2vDF0ehu0IAr6Z1qP4XuZSIDJ
KXasZ7pISaP/S6BPGFTaKryiJnHpju5VL7+n6y+C/hJc3whmlBgq4S94nBhP
QDzfPd2E3lYd/fEhzIRvOTYgukBNKXgg/jtU41DNVdzX/vL8nSK4sf1+UDzx
6/OwPqhnlfTdnAZv3Tg5Bp/02Fsrwcs2umRH001Rx9HFy+O0lukkiqgpDs6S
Ub+Ujzhuqe6/ZEUT+tfXLWpSq8IfNh2gcKBegf7GSxPQamQS4REwDW58hi/k
1+JJPdTL/cy9egCDXfbfrG+c4yefp3AH/LcMdk0YD/d2wAvtWio1/SVc71vw
Ks4o+M3Q3QOL28R0hZNYraAfhhTrdDLdtii0kseDHha3U6CPYYuhe2VsJBRD
iwnYbbif4UIjiZ4LOV/ddyiRr//v/TJbVXbvB8EEmqRNwOt16P+Cu/P4aqWl
lUlnMKrFbjZgFdOWs4SFZbBPjc9n5sjK18yvQhA2XRpJn8ZxLkQxC+CV01NP
yCKYkoNrp4aQWebCJrcQWft0JcjYvJTlTaWnbT8H0DmhImqjvy0CR7qB8FQU
a4+EMgcqdVNhB+kGiT7OU/evcm3qLFIXJyw/X+xtSt+rHSJi3xWv2ZpImmAJ
1svk7OrtRz6zxhxRTh+ODw2Yq3sWSRWbnVNCiKdsI2NOM6EVmV6dlmQn02s8
pzZfjZKZ8yJy4VTNycQKc76BfGbC4+q5ZhRc7R2fGqmDew1tchG/vMQPGfPP
g5i2VQI2rpOFT5ZW9CDp7cV0nFED4FfmNtwCvZZc7fBW5v/XbfnRTk5jFaOZ
oOaOWX88HtG8YNwnr12L1z8IqjdZ59QEYiyCqYtngTkCWfF3sZxfDlayoV8v
KIswDYUwgYKu7s4fjnjG7uIjvvCqR6sNvM/tJSmO1yhEgUXi2y1nJNeKqOiA
2af4kqO7ykJAOr5o017QBqZ4WVPt6zt2dyNTFrofVKTGQgPY8IRNUVpGI7qo
HrT7hAbplh+Jayfw4pYBudU25VoZTh/1KfBUr6cuYudj0A0InMRluycXaECI
Tb2SsppN3HryW42I1mBdJN5764Nam6zV8UH3w62u0rS1mrFC9O2fisqZ0LBK
2oQDDeZ84Dghge2uD2RcO82SCdiADHNoXRgST130DBASq9RQ7BixZjHiXfox
RtYAT3dXCVqZWJy5J4fLLir+EjHT2UGcva1YuUCQFp7idpx2S2AN3dDsuik2
WdbZNfSv3Ulff1rXakd0nOzLwgU67qkgsUAUfaCBQWmSLUyVvGnb7YhltV0J
c796ZZt0sg9EFLJuKbkFJBwlDn/IZcf59K8P15nSY50Wm357u0MvMYwRnT9M
xnNND5aIQCyBnJBFE04knAA+ofBKWfAuB8Jjf8HmcozAu0br3/k3rA4YeiY+
bVUd5mnPhB0UU/L49priwaro5HfMnyPCrmDLNI5R9cEckm2mV9WcZBPED2ZZ
gtN40Qpk2eOkWiI42u9KXOYbkCzD6HKKgsfXTXvMqPzQ9eNKTpBw5xyxGevP
AN449x+yiA58o3bRMg/9Ym1kZOcro+NyTaLqohLx4cP5w0o6cgF0XE/lqki8
eUCLfOtxprOu7Bmko46cWY/OyDgRxKdXK1Km+f0+BVWEkgUbrT3AQvZV1Ogu
8mUVuoztrYBIxakFazfPY2n1JLkeaX5NBrQXjM7eIB8YOYhtwKBz+Zpto5FU
V7I40NRqp5ALGASKaYOW8cuPc5TWSaQFa2lqGTQ+OkELfzAlTqb4WBpFeOHv
AcbbxLmQ/tA18xfJF7BIFCarQPq6summy0CBXMliy3aP77Qte4TeYt/y8xu5
UQAzXFejLKSK9tRs4eTP/eef9FgMTiyW17I6MD3OE18gZ9KePdHujhE3CyDc
6SLmHq3KkfFXPoGaFQawYXJupyK70aKkb8JHv61X4RRdP8VKs6HkuSAjmaxQ
ty9iy/Do8IktmDjNDgZX52HvG8BXJnZsezhuw98mypyQFJiC90tk7+fS+2on
8YWOhR3KGGb4UlpxtGsGai0nI2VrLcj6gr0bWJo+PJPAa600gU2chBJ5Tlqw
rVqwhWdQMdhyZN86pX6L4egR2zon1x6Imx/Vq6sLPZY44ZZzdwP2mKurDrYM
qz+VvGvzfHnsukQNgxVDdL0W/r1CBmjRtmxhtEaUqWL9tWHu5T6zsOmQIopy
jT7zLm8LVQEADhz6nsc0qDlrVyaBMPX/xKOlFnzhv4MTaoNoXdf0d0v/Aq2u
sYi5ougrtKM39kfymsMPoTQ/9Xbm0sEmEifFgR3HL1Xi0NfHEd56L+Iky8lc
0LtFfQCDtDhNX1AHtYprQx4lUfECT2yl4gYJjeXvMQtmhFHWv26xOcKVXwE4
ELHrJE+D/QRI38Af9fNypuvVHHnPyOBu8U7RwCUDmCBqzaPR3dEKn05y3scJ
NFw0A9YPJgC9zmJiB4us8HmoLAvVt0PKFspFvTW14MpOON4DZeVE6kHcDcXT
cOvj6kxSAQxyW46y2v0vovB6xWw0uUqgQe1HFISwfFbH3VvZMVRqELgreOth
7ODXJi1UJZQ8DwinP/TJC0fdHYnydnhKsq5b1x1fBr1T5bFmhqA+EW2l0UHm
yl9IhDWt85IRncaG8aM8RJ9PGHF/XuMw8CA1qNB6O3DH6e2tD6nRPVZqMXSK
ZwGtgdeCzq4eNAXvMzpUammxkUTaUE7mARDulrxOb87iicG0/hvqrCOz0zNQ
J1IiEHFUn+WfF4QhCKaez+OWUGQsSMd1R6ThwtgFb5a2V2N+3luPNgOTbUYV
eB0xsZtP7G7p1iTM9OFyL9FpwHGkcYmCgh+a5xKWChVwdji9U4s60HC4Aj+N
nyBaOWxP674sS2GeKzTPV1bjAPInG6Lp+WI7g7W+5z8uoWvitju9RiIede5B
EpLYHb2GbJ7RPtYm/lRuchURYv8HS6L2gH2tkViKRg1Ygsc7agptvYVzWptL
v6C1ny39p+9+xrztmss2L72Ovceae7YqE6cuR4/X2EAsx7fqrZd8z5jLiCVB
ZHB8JiCNDKbnmTJBsn13R5Hgi41ovatyaLXA/wpqOPh0B6P2nqhwz9n53Rdo
Wx3mi47v/vxjTxsIveSVef4xEnE0plKvFbe/aExyFfWe3Rk4th/a8/V6eV5b
7yqjXVjXjWuWQGqB0A47oUqHcje9G8/HVQbfC3Sv0EEV7uxg2oDgyOizpDF4
axn9YqAvtjE4ble8e0QJAfgMhu9GqmQVpYia1x0K1zC2pANMYuZEb6I89Q4l
JHEvOdDw2t9PgMh8tC1lBpjTMcLRUXn8ImZe/A3J86WRBMZyZ+AzM2cHspMp
dPOBJ6kKHYsbFo2+UiCBmt5RP1pEcd5w2F1vB2CWmykrUpjWaolAwAwcg0Fm
U4M1ezxCZUO0KYEsxmVohGxtDeIkbZIEY72IIEvMwrgphfpM31RMdmmxjfTP
9mmMzx6Z9u9fmlIdKhlEsLM+ojbBf61wtvK7GuyKmDl4L/4hF8goxYhEgDYW
a9BuIaxE932UttrlOvZSbkNymbqnp+xbpbnqrqC3UqXecnxRNYPU29rvgnsn
pk04ZVFB4Bc0YcoR7MM20Yj9V0YWjpsV1XH5elqoMPfF/MpFFp4mHX/xb2Dx
MiczPWTuA1xuWZL+PIzQuxTJ0QuoQj0EU24Nl/JSNjQhBzoUV6/Uu7GSc0be
b3iuQ+EBJb/JOOFB8hsRL9QHdu6c0N+hNRMSnxXYzDZVvES7UtK2b6PG5djP
RVCsYmfdVxnTHLyIRSjuuj+MOKRDaiutSVUaZglQ4GLtxwzcewBoES3nzk6d
u2o9PnORshlauveq+IP0Z13XK54qkzZOiEXLp9nzrz0RhjnY/EBjJVxeEME9
56v/py1x2OEACj+TCIliSED6l0ZFmOqSxyZk8E8CwSncZiSfDnBTW4Ytg19b
fHfjaEntNA5+Z8kNrviLEqjzDAC0aDpYmDn4ewe/tNzfdEBRC27Z4A61duaJ
+CZ7eeDBTrDjrOvnfPfDEjiK+/rZJ3eJ63AdIz1COL5or8xAQIxISo5ds66R
e/9vWO6GnZgSSz+Eg2oLKES+pl+zSWleUrLP1cxQ+E/UFJTzudj/ozVJaEcx
2WU+ItFDY9ZHVVhKanWIdK49SL8tWBVfExdsjghsrx26xqcI2xTCgOkzAYxr
adurlbBzRpxaRbAJ13umyMooUDyZlDT1LemD6zjLHxyg7GY1Vrgl8jC7uXUB
vWYfbpoBdmkzd4o0l4lwRDeFflXRJomP6svhHldMXdkNdCeWETSxX2bZXbJn
BTR+ikXotdQYNlAWrvgZGK0iKo7HkoZAkigzA958NVNVYtROoF6ypko0SgE+
A2QFORgG4WmWL4t8E5G55O4ndNt5jHc6J2Z3Y33WScP6U1ichI5M6ib6dhhl
pQkMvfo/rrmb+nKG6Y7Zelzl5RLuUn8EyBYUGxGI7kzO6urJfjYhWFK/+tmM
C7D1pzrSsTu8eDo6D233UJSDxLwn+Xe8Hnv24rQmP4W8b3iS/H4TurfJK/pC
aizCIHdcjfMoj6Pazboxdg/ZdowaK8i0eJocZsY+ESazNaL7nuXATMxUG/j0
8ySSLUH1VtyA1HY99TFrSj18M+RoWpjjpvpDmsJMgwm0tkf0deVw2uSje1vD
mtNiSFfQUOw2s8d+Q463RDDh2KGav7MTiTF6kCWiY6Jed37S0mvAqTyrbnUj
Vj1EilWNg7hWqlHQEGNgdv/zNQxVXqUq3m4KVClznCCCtoICDwHswpFbqgxb
UbCvIE9Gfn9dwUncgjycFfYoszE/4Ltia+5NX++b24+NSqFWf3+c9yR59ZxK
b6mC1nR6OCTS2/X3tSjrDA1dJ0TRGdC4xOpMBIQ0vzU/znE+Ft+s6ZIkiN8v
8N0WV+axFhF9sF6OuyRyHUoPUTw0400XN2zJbbqHKGBE31qgyTtdUbcTs7M8
AeXXYZCG4d1nDMrKR2we1FlRmFY22EgHNJr83fhuV5lPYOEhtSDqT2Yontag
ndcNns5U4gOsSbntk0clCW/OGZNz/18k7VpUlGBvA0R+STtvy498e3gAsENN
HHQNWY6QwqODfztSEiGwOwj/Oaqa99yKigk6hJEn4Cgb1UILIaVN5V841ISO
aNTe80VV8ALAhV+e6CNs2YYwkNKPwvjK0Ea5A2H3vCKwT2L8MhA2ccSo+C45
0Wt9xgwxaxl0pSGrJrjaXbRP9GFaKqUAYbjkZj89anfVt25cRWLsKtyhmTu0
+VlPF096WZASUEu80OeEMk5yB8q59PyD45PDvtu7zcCgNcuzdneAxcF4sywW
53MmZna+zVaZ0/qQ/ZBVz0K0bzGyBLsx/cYZuETb/LrTWGMjQ5VXpbcvwXnf
/Wl9paPBm4pVXGjawSZFRb+9AVS3xAQAxWyp2H3mSKPbG60wQFgUBww9bPR+
TY1zGURXizWo0gUpBKlQDpOXSbR4aO6fgSNwU6GCHL7N9Znc+F3foY4fcsRl
YA5XUwqHlKoovxvohbGQ9usVOURvXrGYQemSkfiv6Launben7Ez6eHsZJuAr
W9VRwC2Eo/sZWM0R/gsdPNm3ucRT61ViZc+2cSyXfLLsyCSScqltc7X+sjNV
oY6kSzcuqjcOMD++yj79GdCHI59Hq8QCZ6CvdH5jW0B2J/Jgxd/HRxaSeh+J
00SQEFkNGUOdtgHSRVJ5bkALh+8ooViiKmkFp7w3WztD2DAEOaDimigQvY8u
1KeJytXavNcus0MIfBneQ7mdkRBrHqVnSrTiRthaN9Z6Kk1RCeajFjiirAM6
KzAjeuM1RVZEgIUHTPo8yGnPrRcCWwTTQieisjnTtUyP+w+IDiIN7K+LfjGW
4+vfVD8Ssg06Bh2E3THVQX7W5aPfbYTc4Myky+r+Y0Y78z1PqTYaJjuid+zP
AkAOFUn+i4OMqsi6hzvyrDkSw2cRM55Lhcslfq5Osy4/rFTgIU4BzYq+atTg
LONaf0eqU4C5jviI+sh+dDFtgDnWoPVuhPeCsBcrDBuyflL8oGe09JqVCOOu
0tFLd7LqrdyEzTlDFIdKbFXcrhWn2HfuNQ6MxdSAmxQ6GtI3M3vV4D1dxAvw
YEdYO0Tv6tkkV1RUdQDlrZzRZRzTdQCtcCMsrQHgM0iFg5hXTrKh1jMQ0gKA
lidg+zxkLtSlEdsHUPqEEdzwwX234sRWaEgDYolTg+Y4DVPLcNLxZS7+kXt1
A1H6n554bRv1lySVp5N7B/6NHfuJwL8tYIbs1QQiKzqREjv+NtcopSJFzBZk
f0mAW8HAqqaeIoiCtB//w+4v8Uohd4fIlmyo8xdBNA7O+77YZlp3B5sOFTjI
crlCudhs21laQUpv09/YoxSp9/r7C72KN0pIjUNUfVENoV2xMc90EMdsMLU7
tjGMpK8C0ImJaXXepzKdnkdJBke5/V3lvVzPGpH1wCsm1kNqgBkZDdP8Weln
6wcjxiNKh+LUs9P3YXDS0xycc5btJbWWxZzeqUFdPhSaRU8I94XraB1XfcaK
8eZAjg7Fa0nLlMV58LnqDapf9zobAJpHlNM4Wl+VkljFZFqsLrvbJFy55RAg
sbQUN85+PJZzVOtY+UfEP3A7BfZCmXcwaZiGNF9RMth3+K+9RY7GP/X2SQnX
aW4fzADQAyboWVzt6gv6I8pl5F4C+h0Q4xLoC4x4t/4+0AJNkuPJHUO1mcgf
PpSDkvIUAYleFrYJA/0Vh1HjSzrlAar0RJmPKUAnKGq2BLhGF0qsRDCtIDP4
5GNBXxNm9aUk57iJt7kUWz8Zs4xSHjU9Ry/R1QtsZPRUd6B7MpoVC3ryTqiy
E6AZemCWzu/ROIb2q9t0L+f+Zunv8H5xGjtmYkm9W1AfJJwx6CKHgb9y00EF
iGAh063Lv5YdDPvxsjOOSctvkGuk8+8hS0Fzg88YLJMtqlswEEQqbjQLfXu3
OmHXSBTrk6oEXviKtOWN6eEeIuMs6C0duNGw0YGzXungauOjozGxsCRw2ioJ
HM/RyVS0kTJJMgt7MLT4eS+D8RzxKL+DdQn7U6zmpLkHYTTRa9J3/zPC9oLf
rHSP8M5MW/eu7PoLMf4ox6SF4glXZdOuO6IDkTCjt/6hmtsWFrXZgu9d0dDL
ELYLU+G/eq+AWv2dyx2L04jw731yyBqXiyn9ZEUcLlu4LBEa4tGQpP2xYOnX
aTj5CyffwqEez2mcfmCUwcJfMMKtsZALG+WuWUowJ7ab9FcQstGNFkvEgU3i
MwwLEffoT8JhR2IqrAw/8uuJ0kKbsYrFZfSJzAJIGQe0CDno0D4rZHT1WZNV
hi1MRdwlqS9YDjI9H/CjQLd2P3Ll/rQ7SmzziDLC+g46u/V7iezASy9qNrP7
C8tXwlCPiiBDFroz9JTWCufx4CG6+PuUUs/OyQVfESL3J5WNvXdVoiF/Ymgj
ltPLs2Lye//wP7dkthofS3Vh32Z42UleiMksyMBln20aN7RGc+tnN05Hhf3C
Ucl+bQ7G9xg9eBuR9wRwWT3PBSGzF4QOALWxkf6Y0yZ9SrsIjboB5THQEWXo
+C2A7P4zpDmVvNDIernUVX9UVoOXsN/iq55u9+M9wtc2t3XPUkX0twIyAtTr
nMk27eUpiwXgjigf4I5eNde0zvjIx/shM86SGT27jxeQtFUvHclt/CMwESy2
qaoOmi9phjeAOmmdYOVQt0Kuo3g15+aujhv4LyekMqhuq+NLzUUehgSmKOtb
pEFHvu38I8up1ALzRBuVdmZFu2WR7pldGRBpFTQ0Hsxh1BhwhJ6c1cZ4gQCa
KXLmrcK2G2Phxelq/W6KoOaXic3/Q4TIhggly16f9GNCr5ezwjUmVs0r1DHo
eD2XXLUIWW39N9sBFw0c8IQyO2binbeuk0IToC5quBDiYlPN7gh4w9rKuyD7
24kAizzX/xwTJMNUiU5wISluvpPWvBfi2FhQdTqPj41uNJj380wV9efZL6bF
qLTsguAE4e2oCsz7B8FSOjBBOKT3+SIr2bjU6P3k9BLSni5hncD+jAtLZ4ME
wb1eW2Cx88hxue0fI4lMp5laJSdJvkyRNN8Mko+jcvNMZrnXpXTTEp7G7dkd
xE4LOKPC1PYPxU30j+TvdQ4izG7zBC1xZ2eXVp3zrckf30vICS5m3yc1dE8G
+DZZoPcGbvswyY4Ln6b6DmYY0VEra/ae/Nwbpth543iocdvedLKiJK2KBAlN
2al1ZXY41RcHT3iuXorst8dnBr7+sALIosh7En48DvHx3877oYPf1zw2VkRJ
e9umG7fyYW3N2NXZE760epwbAmRT9iX3QMrUp99nm33JeXGj9w/RNlwpvCB1
vl3X+mu7juVO/b6ZpC6XcB3V7MKHABqPI1Lr37wXhEamg2+w64WxMp5vYF3b
DXzFij1aBo/1De6Ei7TrxwLKnAmmWcMj23eIA+p5L6A5WzdhZy5u+29ryBoI
Qw+G+AJSUUBHguoLtwBB8GbGaSk3T2EV6UX1ZGx1WrqeSroaVroFHX4DET9m
Qx/3Y2CvWYIhBEz5/efn01DMH8dq5hOYNH8dSKA5zZWPJRvqrPZJ96KSKh/j
L/VFTRTFxGr6LUUvmV0mxxE9NomnWQ5VAkhOi2m3VRCG0CseZvDe1g+TV+XW
dvfxvZFptfiVUAM+pxviOG/dt7JFSpQJ0HxyPGX8mCXXfw+Do2DGM+o3FtCS
JfIxQozHrViHpGEEt4AbOwJUTDc6eqVZPbAzhs1EuDWDby7+3P8j0FZ2PUbY
YzIXJHLse1QdcfFcYxEwmwzUNO3wN9dSqIxk9hJxjDBHSnMeSZaHdNGnZtg4
e2YxOw8EJJ8/Fvwdhv1uQsrZeyr286xPut7sO4/6tU1S2tlZ+JbVI2T9oMhM
SKic7K0p1tzDTTkX68jEG6a7CihXfUdP4Z8y5P9INV0vjhv2KUBLkfYDwUkY
leRg8rPg6+uFwhspAJzR0frV85zn7XZ2zOYscgSZactCYLpmfCwjaGvkOf+Q
6muOJyfW55zyd1pc2MjsFTVUM5QOHw5nyFbdcjP177gTElzdn6sWvTz52TD4
WYG6h8A+c8jrACGU7CzrQtlEZcR1U18umRoDqGo94fdBAupxVURCLRxASZK3
cAX6DqiOgO/Uu7pp5q0SHFFsvcxsglWnCEIX7ytwVhnr3iAYRI3A1jiNGDpB
60bTOoMAfy9xeIs87HvbJnCj1f9PY53D79Uo2kyb0XWTc1kr7dAdcOW7RR7+
eooqesu9sl+VL0wufw3VEc85jHYiAq2AAZl6pWnyI/FF6nUYrdNNWSmCKlhc
NG1h4Du3s0AH8uTyY61eW2Y79NVfMPXj3dxCo2nORaGAAxG0QYAlGUNcnhCb
wg9Q5PL4YMGAz7WcPpXJkwBkVEfqAfch/0Pd8hlTqJqg3VB3rTeKSYTFTFVG
iaL8NiCOpHFyhj1ZztUSAoMsjwFYjynfNoDjaMODUGFR7fKBuxiOm1452S2c
0JVFxFl4t06hLI8lKVvuYMV9vGYZVJEhIzPuxfCrm9OMjW3LEuYtHOc1JYDr
tmlZBIeLAMPJwSF6oJBN1asQ5ucb7jiU08sFqYk7XivUzhvIqdVNubI7ZFma
6Mub5r2yfJbOuGwdZUThAf7weN51qGxF1JPG4961OWXvjxyhbMGSadsoMC11
LDr4+9Lm87/g16VPCApcrfcj8mUz07m+M4hPeGDLXSPCDa7GhJlb3Yg9h/Re
5Y69tEpYYvHDNIbCSwKC8LdTdibUqmG91TjcEYLeJiJCuCmqueXfogU8STbo
stfW8ykYqHleYNGFX4+ooEThHq3hpL2C+YaiFad6Qkc9QxAZ23GXb7uLHm7p
NYFyfTBhGhtREXHPbgAHrIgGOhYGXF28oGJvawvvFUeedl1ftMovS4RPLm7n
Jp5Fhov1wMX6mlQ2YQfoXrSwo+QCqtVSRJhsW2+HJv28jXD37dhzI6eHIgNb
mWD4DE8uqcB3cL+2u1kKx7i1afSbOclgQ6h+KKbLgMlDTnLvg71+Ft0CmjGc
+v5/dBoAGunYoSJnafoW/bemasPvjaqPhLqW93HwjqSNenCo3YsatNqFepyi
aBH/J62fb0eeda27jojg0/00xQNHhStDf5zQWe9o0UG+HlfoO7jwa2FgnDUC
6+ZaVDlACEUG8AbTp2PYfefnrJTM60fA1s+J8kEqT2zm+E5nP3+CmFZjgIPe
j0fszbARhQDZmdsqPnDu+NjcpeyqssBHA6/n/ioiLdDusSjaQ2PvEqoUOCdY
lBcYW5ppgyNnUszkMrBvXuxXPb3F719p8JtfO6i0uhE0lD8DaW+EJdvpiJef
Xf6DFD1tkPIJ7Ui70fsvR/vytMVHls+bkXKiP9n7FvU6fyQx1JL1zMzYAJQn
Kjb0+dzw72ZHZx2md2vF7CjjKH4cvsLMKsaMRO9S4uzFgbtCktgi0W3UH1Sb
XP/V+ws4p4hjUjMzEzm35yXIPBVgWgpa9WTg8uD+s2kcLe2Db0nhexUmW0+f
VRYkvk7CKlrjB/onWPh93PAyxKPLRni3MfeDMUhZo6PEVRSEluIb9WTDo9eB
4dJSuG46p4IMxazsuBmphjC0zG0FSp5sqg0m5nOSnD80bi2msy4M7FqHTuLF
glP56Dbl3xxt2zUMc8k9Oj2uMBYrPje31uwdAgZx+vCFJWsTlWW5zPLWvgtZ
IKBAqgYJSLklb7xuwPmtBGPEnHag4cp0eLij+XOSTdfhbUtwowdJsqGSHRfJ
wwYJDF8TGy2iuZ8Q43kX2QiZp3W9DRcGZmXM2oIx1lP6POvcZr3EZLWu19ZG
rMvCSd43hebIY6GVFceDoexElrBtWKtLg7xeIMbkTIIu+I6tUmPmwYw5JHth
zwLoWA5wE3B20dgKkLJ80Ld+Wufba8i0EBNHCKeWZRBg1s59Cd48spxgKXEf
0Z77TmDtVATONDpR4wkMeAtDNHJ8I5oFKtlUXVvpi7+H7gbPQq80/KxBiyTg
jukuDr+DGup401qkw3JiauxY+EIBmGJpvairV3N6kH+uefCnKtb9m5bpmBkD
iuP2WQpFXoJ69GGbJVy+VwuU+ClTz+izBF8wjEZ/UUA9TdkhqsGPwLtetE0u
/Xj98lM4upMkfDiIWMKrZysGTnc+yhZPjeB1CjNxUL1WT6Td+RjZDnxQoFPm
nSa8Ss/R/t0eRI2w/v7hGd2uE//H6gwAma73j1pCiqNNdRoU8LmgqWKufMl7
voQz4siBykYjiAR/UoV3pfSc2bzoMOdMvIAlRxxkCrbwG1dmthT55xuzTYMv
BxJFVzirD1tQYwWwzf6xDCUrCGoQ8wDr+sCQaVy6SLTV2Ie8eRqG7Au8KcF0
ZyqGJ9vNObVJKzbXCkhbGvJyFYPCSkw6eMrRCuNdo+j7MbfZ2a8PB2sZhpTH
a579WDZhf9sc+HVWbgKnrFj5gTy1Lso/4jIrWS8zQdCtBfuBK2RUSWvVWr09
4L8iEUHyOszyoqDYMBWSSfgDuYguONhqqSG/QDPR4810WY6dap7NAwa6oBTJ
0g4Uo0sD6rvAy6OuwcE3hLqO1ESUguPxJJ1cavTljHJwLiP6Lr8meDFrV1G8
s6g752d2taOb62xdcTYr4LTE//0DgQx3CnXY6MK+wbmcM7YE+zp9CdqFQwBM
b2s06eM9TvqIX8MfKzAbyDxPYMgAgFXzpgz+gAGHs3mmBtX09Q/iaGA2tGcm
ckbcNTHs70ZaZ5dr2MqjT8OeqmS1/1KdfS1YzGMY43c5WPfSIt7HEhQQO8dc
xq4k/484cXQD27pQABPsnfE0eTKJMx0PTduPNDKXAvBupxMheSrBqX3XXHu1
zy2z/s9ZktNxNDCpuxWqKed2ac2ZAH9InTou3cxzwwSE18miJw6mDET9I9Wn
fb8TPQqq91cBR53BOM7zzkS2pwvIkp9qsTgdeF2qVu4u4g4hA1IN/y0ErTUF
sP0odSljmlvhjMxaTk7gKLxDjBV+VsqekaIzqyypUesT5R1LxQsMLoq/OvdC
Ov5ts4Rety9o3P+4ev7clOGPT0CbxUPTTVfjjEkejNoA81wPkMowFBWEcQ8O
py1yuu4GHnir5C25RdZXkLviUpoJXAl7W0kD0z7l0Eviye3RoF0yWWtqqBwH
wRcce1PcMjDn2WptsHyEquhQ1OHDjoknRmaEjFuruSLJPmpfMUq7lNaZeQyM
rCW+Z/E6LdBFmKMnd3GizmuF01TUJEAHAHvGKshx9c8I3pmfboP5XKxhTRUu
2KM3p+En1FThX5v5Jwzo11qcBHpivKG97zjyqoN/NawPxa5DVScSIt5ISo3I
mYiCux3/OAGlgnBl+AosxV8NVS+yvvd6zUVgXTYdqhsUuouubyey0ybvqV+1
2kF6DMKxbCUEhmuKspOu177IjUMnYPMuht97dD44yfs6mnzPGgAKXarJiylB
MzP67QpH/MSR9tVWN8G/s/J2XGkig/VNGQRxW9jTD5xI8wxVZ+R8ANUhzQIn
c/efqMQwsfEbVaTk65kiJ83CPLvKl27H+ls14BrAkJtCv8p24++LuDwMkMJ2
5GYdHm/enqefx+QzVBidvn4lWehVw9PItf64yjz1j1cRXSFmEqwBIc4T4YFS
SVW79pywGGsMgwDyBJN+90dQ4e3eq4moQcPuMRHR2t3c9cUrA0rRhr2D6PE9
pS5hs+f6rf73X49XPTdyWqaxopTxTM3PlBdna4mJR8B7sGz8vUPG7rnMtlN4
1D7LRX3HdSsHAFyX6jPnfbVaKh5KR6+tFbT2YBDLY7XwWLNWBuMcf+Z9Akd6
GEPXwKb41JaixleABdphgNylsBypgu586mo77oqGoOqqdK4y8znJKDucAxUP
h1cuzCpKixw/zOaDDbXy4GZHErqiX4tuK3JTrW14pQjFo1pEOvcDk1VPif/g
LuoCigNiFRF9H4VrX4WoNDzHsQVFizxGarnlVc6f8WwazmyZMFG4C+RQSnP2
evyDVcbBDAniF8nh0E2WH0lUYIy0vxhAYs3fuB1EMFy+9j1dO2D635oOXcIp
5mKJCgcMXfgVUGqb67mKTO/Lb6iS1d7gKK9HiPGK+ApuPza3KDdI7MWEKpel
0J9cdIw7xM5hNBBg4/Ygwe/MZSKGfeko1O9icadC8q3Q2T/7xU6Iy1txEhft
qL/pgXS4CzbZ/FVSoE/bvoNDozOkVJK4NAc7B6tkfiRpCy1fSlthJoTaQ8w4
qoiHva1z1B/QOtuGZcrSKpGId1jS03+QwQ6CC4AuT2249vfLcj7SQPltzl5E
x9fEP/2Cm2Fur5uIIGVP6YoenbFOHMDELdWsaK94lE0gl/zzeinGxj5uuemR
zEUC0X3O9ovtIsRq3B5Aw4w097xCfDUXSCFmZtQmi0S8it0BUAkML9fkULbA
VFeD9fSb9rlqcb82u2lUcjr0Bt7KuWeVlB2bBR/e/kKqSEhOrDtWEubyvFW9
x0Ma2HMUOtio6puS74iQh9QvJJTT7DDFGya5E2pqPT4gdNiflr08cs/9NUlw
z/TL7zfswxKNl1KamI9geeGHx25iamA4y9UPyIRLa5dRFsgdSn34pMQV/YFo
/oTUBw7kKDX80t9fCjLRQ2jdTuzYZlY5WdGXO1ktOBhb6exoa5cv7lxArPEJ
rC5I9PoWjLWLv8emQnumGdo2QzPoJJBeuXuWmrE6+/8shlXXIW8HspYu9BSL
atSNmAAUhD6yY+efkZkKH6p5cfbV6oD39Th1rsLBJCguE3bB9PGR62dz5w41
bt4ZLtkwaddWfASqyVOAIySL1ZCqAtud6EOc36wv8/OI17sHHvvr9Ig5cZno
XPv3MRX09vGs02hJ5liK9pvCay1Dak4Ge11V3bExyx/MmmwquU2jA+BWifi9
jRIfZYKueXvQfeOAaYJqDh1tgRouJYFdjrQ//s/PQgnUEcqgfEuqvKrv/yDC
a89Y8cV2DjdO/VN+9h+13KDJ0VeveyaZ04dExygKaC4+sDWRLz1LSr5zN7wl
T03jrNg07AJhTFb7abEwxL4XQosn0NMcfz236pTKmPw/uGlvVKwqsHsaRNgh
5Z1obTxIpjGUjZ6Tjo9QJZmRxb77GxUb7iVOeTQKxhVKynopY2A1nbpMXmat
cYhJL4/B7+YsF8Rbg+93BG7QPxUBHmq1h9tth4rKmR2LoxI/Jh8PCPWnexG9
lHaZGtRmO1kGBlbETaoAGI/9Z2lccyswC0c61qzPb4eFnNVqsA4Jj3vC/dvW
wReqcITvJ6B2zcI60oG8rtvE7k2EK+vdP88/EDBrFeE75iu+2mSLohaxZ3XY
vz/r2HKQJhgJoa6NVsngA4Vtad15IcopELcbIFP5XWdooTnliEt3G5eI8wKX
TiRuNynDK1H+5udWNtNZOtW2vucRXNfsMpOYonsYLqSGFrNoGjVadl9CAtKd
sWm9wxFs0El7q3EhKVcxAGSHLVojXrofmXZ8c7TUqmwwjK9LihR7C3uErdeM
chSRtc6KVWU2mEbUlVmkLUmx5MR98LvNAc/zV+7lCAftLlPuZ3F+ytztUKIn
vPIFUO/keapv2k5BiFYMOyiOibazNm94YtPnluaTprvU2dM0ML0I39mOm2nF
sl9Z8IKvvWLTteu3FXVpgE2SBAE0kjDIE1A7GyHMUHa79yEINjHAOcXdKKoG
b5G36ql9woaKaw7QX6efw3ijl31hozjv4PtfbDJdrsFwxgvoWDx6VXGsF0gG
dSfwwbMN5KUGfzUVBlDi623CFfzzmPziVE20siaQ46VWzkGWMjBVzJZeT6d9
HQGgj0UbbSPLCSLEB3TO34k/1gq57D9Sl7ApLKmRThnBTQqa5rWH3hyI1ZeA
RFDx+D1W7AtahK124XRZQNtbwGUXvTFYSQaXg7H+1U9RvpnhRZP5h7rmR43W
kkTo4nqyT8kk6GlJFAr3DCk7sX25cebc1xkRZh1Sg2CeuaCfLALZA928+bui
HG31Odw8k/9rvrCbyDAqnNtP5lqC5NJAr+Btgr1o3hskK4z8iCwF+VJ/0mLS
EDDY8EUzaPuJpPGVEclyr//t88vag3B/CHSfm0Nr7qT1eHwYp7iaiqSd7fxs
Atj5MXZfH2mlkQmJFCtJmciDmc9cBxPfeT+esX2xPWbBt5BjOduEY/4S1lru
bkOoFzQpPiEygJjlSnhc/2dH+/ts0oi/zsXWWbUK1WlRPXcAYkrFF8ZcLLBO
3L546iMrOetwe+SONix9dA80RbIc7iRp52hfUXUfn3/PrL/fPMcb7va57f5P
jekhhFPle8mVmdKWf6G5zMneIa0w+o48OH6DrMcQ2s7ODNvlww2V1kPyzFlz
60Oz1BmTpNJvh28cyhZOrtgpgBS8LunJSlaVv39sCci1L7P96Ho+qWt8CxoW
eQ/0YAsHs2yse5oQ/DcltrR6YPVj6Hb/ziGm+nY84VkElbHThCMWG8EuoQQp
t/FaolVebc7NcfBJ8iv1KPgtIL5X9m15HqpqXzPIDhQMYLzo/0ENlEA28km8
p00DNOTJvxhQXGikBKB+CtZocb+49+s5ftnp8vNO6gRU70gtNQWAeKgw+BGO
MuUdPbETsUIJ4eWaEip7uLPSFGyc8OBMSyL4NP1ULH1QmWEghbqVI5CgapXY
zZI5L/1HuWKg0vFiOLzl1eZ97w3J+Rptf4UJOf7ujeeRfTPLYKO70L24vezJ
x/1SLSqQH2faYsMQQHkr5uBHlRB/FYKhdPr0LT02Px8BFxFlMtQyIAeQ8nyh
5P/P23iXWJz/utrxe8TBBOplDuGEC1UZyj+vwJJ7IYCBb/rQES08iycqnquR
O5NQvpocMdIrhUJvwfwJ6L+oceSPmJpK2qCPYX81oyFdHbwM

`pragma protect end_protected
