// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
DMKfscXtXR2Q9Xvu7t7Y+DjLXITTtMTOUywqzMWa4uwrR/9jTvRlO50BgTz0z2Cs
2onjIe/Iqa7wQBAy5wxCGnRqXzirFYPrGHJMkK2jWkBVKg+DSrqf1Nyf9Vd4RyIY
rRg90QQhaiQNuNXrC1NPxY4ew/ZCpQ0w+oL3g5oYLJM=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 120464 )
`pragma protect data_block
0Qt1yUzrhvIHDIIgmFqiTI/SN7AF7+gzzT9iKxKqRcD4/3ZPNhGkaKcc/MU5/gHG
zUizo2BP4MKTZCFHDuyZMgsj2mBiDAZzcybsoUg6eV33gher+jI1trNe0Wcvushx
DD7JwbFBKxin9Xf6JJMJBMkSWIaI9fUUETOgtjF5mm5r/a1VNZAR8zcTX8chpA8q
PfVaOeFVWFoIol/n3JzCVBBU0mBkhbnOMZkuJYqzsT63wRRRKjgYOzmU0V/xo+Dj
bnQBlj+Wlj9c3mR1q56r+izkwnlo2qBrXHSpI41FuVTzZjPw82aOSaqpC5RcQ1Ft
JQZICzEnWazI3+RjRO3H6YtKZxAF06Yu9OB+qIk8yBup5TjolT3swlXTqLicurzd
dUBmeEBCaQaMRPQrhe5p5w6P7dn1xgs+1OzGbldggqFS5Zl6OzM5xYwWeMPyXMIZ
k24PKM9ktoq1lSSyDcD/hfbYqxwZcgT9SZxuGvYxtvAPb9JWTYSPPY75QHnB9a7A
/seeYgffoFqG5msmevm1QopQMcKsThe3frc8AvHeFwcskVJNrNqWwfVbaPgFiQdd
F5zivTQ9zIDqanKwGP4XI2m6SYiNHRBpFwC8i1FN7pzdk0BnMfaRO9uaqmteArfA
ok1E6aHkpZJKB5AdQzYJEB+QiAK/tuLKc9IGWwdcNzv8vVTSZDgQqmCM/jPzzelQ
qFJ+uL+LrjbQIMjZgFsJAiCUIXdtS5AJkPykGzF3Q+DriSy5R1o+REWQKf6+ydAy
xhWjLH56atbVFJY+HrkqOwyGzzAuOZ3UdpBZYZEZM4jorPhm+vi0EhIIIXNoCz6Z
fvyknSZdvW1kBi8H8ky4YVs35fuIVALbHrUvIG1+hVwrQThlTOVJKygS/kvaxWxl
WspjVz9ee/++LuLeGoJQxsWz2Y74dcJtk2rLKKVRfdxx49Xq4Ni3LEeSJetbTylw
oWO22Dl5fnH3GzbOXYt15Ih174DrHvSbOHxs29GUEdFv3AbO2gMCxF0MpKyujTuk
wF7faVJL9IharW4PB73CIspV0eIW2n6nEa0HK+8ZXr6MjzVL2d2TyUMoVNNVw7aV
G6W/NSeDF54flmaSSinaI7hNyX9YvTeszwixd9FJHX/KQR5/6WIpre/ewXMMJjQN
DpLgBSvldydgda7Cdjvr21ihgZSZxKAkWFU0Cnj3YkhAS6rUMqb/kwwFbg8H7AeZ
m/TfugIfw8WK/o6zMSRqAqiREYQpADhvG7gdvoD3Mejt2m8gKOS9h4SyOC5v3Quv
6bocYE/i/R5Oa7UzRtI17QAPp52z4qvzcYxP1tX2MFT5rLtY/aeK7C2NUaU3FzY9
6rwfxH7e/vcdPGbaPTlO2xQZntzy4AJGuO0YcOY5LVwW5lX5XmeQKKXDt2h8BF4r
ZlYg5fENPW1Cobq1LTZbG1q/fmUVlGgfmuQe1EWNsMFTNDRcQt7O0pmG9Dt40xXn
RmZSt21dqtEQFEuyUeS5s0wSV1bU06QntD5Y2zsCBPCSFKprz1uEJ21qYZMaInkF
zOTk5PJRdwz3l4fSK6rQwdhG/QVHn31+lZnM3V6urmiF/tI0vCqZI7fauh6y2ea5
u1T0hLqXgIb+U82TCYxrWVWglcsqsRUT3baWLez6KVgcTWj9fHCQ7IKh9GD8DwNI
1HkXNA1iMY3SVnEdA9h0UACPMajkkk/+o4EG2DIPkzICHSn0eRZ+CLJywHh2GaIw
QAkWzN+RDCwndwcBQF8ztHhz0dnw5b09Rc8R+UIb/QydnL969oMYlrmqhw7DQdWt
Bx1wbcWlp1QnQ8HIirvHmHglzDNQkGHBIwLyrzmWxnvXUVQ31HR6xokdwS1wZ8f6
SWkqsM9FPFFik+D/JS2BqO9gLmZpSHOCGoRl/m0TGZvUUKhioNoEIF25+w0K95cG
4Y0Yw83j8GfHpw9tgHx4l2ktO+IKzBnNT1LT4YJpECu/l50KoGNJJ8V1dNfAoPJw
d2f38HK7bqT6YBndUB4Iu2IoAS1avhO+Dg1QZMMOBbsbz6T3yTztLjErjyzUy2dy
19z5gQ7nI7f6fARDslRyS6lG0TK2gw+4eBwYOcDEQruXGqwVYKd8+kkl1O0fXvbH
D4GpLKZ7zxjuVepULb9f7LQ/6TEDRSQ8EI0/k903l06E0os5OR1ghNXaXBX6fras
OzuA0Jx6UZ53sypShw50jt+G9FHg3QHwjTyLY4ESujNS4Z/3ErvQbbA6L1QIAmnu
Qoe37fj+hPl3Xn0qN5ppjaqwYmi5LCQ3g+ny2xe0Xg2hYwZeNoeOkHSBTxIgv9NE
6jcxTSWTMakby0ph5/ICH3KZGX8yleLrQDr1Q5PBgPbwNSLutGi5v9mtxsyR7Mdl
kx/pV4BT7WW9eF+pF4rJz/TwGHT0hk2LsGpJD1ypQoprPyJR0tFTjFOgvI7xv8WC
+GinvZSTGUokaqvYOIF+S1ROKBio1nZnGjuMfHPrYXaXI/g+cYjLtwj4x44ZX3Di
luSkMSdqPVt1h1Rj6bBe8Hs7/ARdIeSylFMbUuuSU9gORrs2/muYPcOURKpWurBt
yPH7ghSkL+FoWCYFyv1EaSqYzwO0IyejDLsXEHPJltRfWMunIfWDiuZYZUqVfiRF
+ef2XX7tNqX0WqXjVtjRa3psl5RE2XhGzdWlgQDy+S9w3BoUi0koORHxSlL3s8mG
LAkQ4lvHQah9JmpNPXc0fy2pOJ9/uxepqt1eZ0FXwuTuieERwcpSgzYyu8F+tdK1
sqOlbcoC2mMQgfsVQGnkgE6oIG1STh5ShSZ62Gu2emdIMyN1iJU04mJ0AZxuP0oS
ecicxzfofGD1KvtTevFzs8WIXjWWNanl7n8B6xQKaY2uyAX8ecp9b4fhZ5AYaVRP
s4RWd9qhsJ5CikdovBDuP0uIgrNwu2Fw5Sia91Li0wwZzLraq5cFePsTvWinuZ69
r98YQLf6bxyxyWPXg4z2BbwHutj/fOkm+qm9C9Shn13q0gTlqQYmQBIvTYVCA9wj
jHY92FVeJlA53iqZwSsf+6RxCA5knm0DKNXRcG+P9Muqi3KKrUzALUuK8YlBkEHk
Ru0L/oQjTCKo5ZoFfiCCIcgHvS2m6UbEIs8zqiIJNqTKiLH5ItyQbrUFPwwTc9cn
YFlFaSQkMvUUAakpa/fdzNxqCmUse+Z+NPmffMjyQ6Ax001Awr9H0jld6arzhLTg
uCPSO+ktl1A+4gbLJrZB/91RV5Ex3K5Ptu4BtRwdKCk7ybnjTDaKWaCkHEx2dSSY
1CHGbdVwFNTdkJZ+qtGxalJl9Lh5CF+0NqtnxbWG2gRYHIyOTgRwxVXZpa8aj3Ui
JLPYNkSwMDd/Ei44EFKNRr+81lW5ZJQrrLrmboApsD7No8KWx+bqLe9Bo3ykljfN
rsDw7wEAd06Ta0RHVMRuMIqYZlA9FuzTXSPoYuRllSpHv7xxGFD14n4kw39DPk6a
piNgs//JqoMdJLNfqSjByZL6TLVSAfrsnlvDGiCazeFtSZymBe1uiuoAM5vBDWxg
htwltZ7KHwIzb6g9oN6+C1q0jYanszF/Ph1XHwIAKqWH8DodWYECAMmt1cm8+lmJ
k1yVX6YKhEnT6b9/CXhQsdidHqao8VQEOkDix3ARj5hpbDMmRwLE3f54HBqUNdqE
WIMhcta20TyEbm+dfHwz1e9VDeKZLMIjCGAxMK2MHW2ixQIw1KyhweXu6zulBx4t
+55cJUe4DFLuPnVBOF7W9SSSSIYcr/Nw6uZ9F5oTV8yDMh7LfDErCirT8fesE6wB
/T5z5p7dLRp2TTK/f6EfEcr8XVFn8vBxjs+sRkU+SzUAOFqK6mS2OnU3ZwtAZsw3
36EEywjCZNBtpgQObRMmXYnZhFEPST4BvJCDTGDrLswGDftO9SP85euSyf97QKau
ViKLq4wEEjVhucnaT9ZWIBkuS2Do7icuRv6Y/m090xFzlGX+HqMHZ3fgYb3WryfS
FGg1+hokONI31MLJ6pha45FC7yDqO7srUco6kb1CCZn51aBP43HojxPeUwC5EUbq
5Xqla2mvFTqZ99pj7BKEritM5966BbgjMjiQ/bQAwInCUKEpSJ6RbtmgS3FDMc6Y
RH1cgPBJ/K0VpN2TRbIEpkzDuwlWS/mNelH1GTtJ8+gDaq0BpIK7YO1jTnSZGhyL
tR1/cgDEnF6SEeX/01LIm4E/wEa8Mj3xkn4OOL4+XaO+I/4k5LxPk6VGs1prxIT3
0H1XVUEcHDeEUc8rKseBW8PG/1KH+SYVvvhiK8GVsCW1h9dviYmKopYne3XTvJc2
t4yUHn5Ftg4bVjL6rWh95J46gJANmk7dF6hipR0BhrfW3HOLKUaZP3GHOp/9swly
fRLqAzZjNmmkUdjwVeFo1doBzOlwKhe7Bv/hymEegH8Ug2nXYO154ETg52VSGiMN
2Nbigrh5Ga5m8zdNOKoL4eRVQqQrUVrxUVM03+SMtzZ4HO47rUqOIsaS1l5zH4oZ
coreuB5MaDGfITG1FPS9J+nY1/twnwfqMQPPs4PCfKkTVBclAtD3wm597515wp1+
vPt2uaEA0PnjUNvvQ/rvYDreKvHEkh/0LeOtSn8soWa00CscOajOf+rjxPl3dKuM
c83LwaXGS2F+DbDoMqmXN3o4iaHdDh7wQWtXW92lyE5DABBP8GZAeTQapSUtSOPi
Cf+ZVdrtNamKfDgKYr7eORAWRLv+65QVJCCy2nINshtS4j7orLZ0XUK6P+tseupj
9RN8JDwiw/C7L63nAtjfUAjmg29oP32xpQ+zimH+M+HeRaxvb32Mb3k5Rq9F5rM4
q+RBhxRdjePvqZOd/W5b5yQV9ptDUB+X22nNJW1Y6Hll7eQ0l4rf1SL/JAlfWE96
MpM/Wo7ipDTORXbFPgJ/ZGZPOjAVRKMOxmzpg8ejdhMzuQ+6exG4gOb4WYG2OcuH
us/LYAecmGKudrwoo9q3dhLaRTxthHiUHPZdqbYvbWgIAkzNReJdczZGdEpGQGPE
yuYwxtTLJv2+fCGj4vYqbIpOFymTKtGJ8zo0iH2E2Vt4sNBxGxXCjW1Mr1NFWCyd
U1OZ2NzSBEtSPusD8ZfZ8kIi2oq5phGNkbEPamVueJK056BD4lsFDzYClhxRaeyG
upkz7zBvOWsfVRKp1fBTqjkakeu7cd3PmAhw+tIL06WG9/mOOWq7XjLKOTSa9nUJ
4tsomXH+EnFnhJZGRdsqnl6mdUlV/v8rbRwkXTx1dBtqHkEE40YrV2krc7ZXakhb
eyZlCu75j6c6TiTornA9v+dgUxVXznZ1I/3xSsBdLiSi2/zyeA7m2z9LT06Tpb/a
51KykdWlRfW3UNxcyfFQD7XZn912pWNhedah9VZtAO2WmgoqzEtR2O6fmVMQeBfa
/R0vbFozBzVoWKN6Fklv1p2Tg0TUvZGwjz44mQZnMEM/3X1WYTrHjnJ9rRl1JMQ/
Kp7Tsp8hh9aWTimtA6nGTTt+IMj8RoUuWqkRhsrJA6VaVvjKXQtw4WI2KGSUkAab
eSr2AA9B6JbfJtS1Lmrj1ivpFyYbFfqV6lJIk3A98q5cCa4xpX5rXSha5RwtQ2Ph
K9SWjoU03N6PW2NBht6azNMsMEeqWhuBgrEWqk1QFX4hr3/f712gUzyBfIPpOmEp
/UjVM2J66o0DDZjXOM2im3dKXg7OP41m/KTWQ9lsCUjxCmwWJauUFq2WRrLSbZ1C
2SMJ7aOK8Ohb4DrR9EmEnS8E6BuaMlQs/WsRMXghafpGMQ+jdY/v+gvaH9u20PJ2
hCJZLICoBkXCRfpCdLZJVMjwh33sa3lnPTpubemAgLLZfJOcjzafccdT+r3QBTOF
8nbkP/wMRozTZH6CVDApbq8EfSdT7nfY5UXso40kmxBxkcLS+7IbiXM7V3LVTHme
vZjTHx+5RsD0pPvADOINK9ZNKclknXl4cJbnfLH1wIPpkJ7FsbPcbcNQfERm6rXl
32mWWcBXJQ7SMeCNighu8p7Ydz5prW9X8JtE/Csy4xa4xOIuFTTbEkVgk/ekuWmu
Oxc97P06C0+gFuNcP/G9v+TwiIEYnFV21msb1bvhc7MlG1WBRxuiNTuIB5YaYhcI
v1OU7bRu9iF3dszHM0ROFlmoVOAi2e2LA3t2hjd7QCEM974ChQ21D8sQXH8710Zp
GeM+Adne9pGxXFkUA7FGPZ3Pn7qpH/wst1/p8uT1XvS6+ezE7es0bz+0DH4uG7dv
TEZgnM9wVDOTHBEu4+SLA1lLV1rroSIT3dvlBbJSQHj3joEKWGAujv0Sv2UFoiMz
qxA6IcBQ/y2uiOEvCz+rP/Skuf44sddCTV5tNXnxYz655d/Q/kgLupoqB+OoTSMM
hRV95hJtpng+4HU6Gz0ZV/AOVvsFR867GelwwhAwWxuoN4Dl6KH7zTbDd37iRISK
kZ2SXbBOVCGC5NqSIJZ7UhWVYYOfw36tCGB4dpzpEEECsoBbBAhSH0jIJQuLF0wo
QwFzYipA2xKOScDCOpa9iD0qcrVmnslPvwIinSpeplqrBy9lYAUzWuCK2pJQ2hE9
Bu5lcAQPsNkFPjqfbpSWCCvattRL81FyWMEcT9x9Redju1SlLXEcTei8+tnGUcG1
UO8mD5lGxnYzf+Jc4OZufKj5xXqEHecA4cYM770k71chNCJGvy7IomgTUB5w4G6r
kvofhpcJU4kU5ez/zrulC7SqyRAXZOzHmNNaBlKInZAmxRZqszvSGpkiC+Ee20F4
0YyUGRfngTgWomvVR0vyX7CjQ+tDm1QTWK5/DG67JeXQHY4/XAjKFtOyZURIDQH1
DZkNrvTjzgV1QsNb9aJcOhsWvBj9QCbu+OT9GFL1nF2XoFnj5Ui4q0rlmSHa8l1f
yaVnwuXENiK7k/gKZeJH3CrYew4wtKw0AN0EbsASt3FFuXWPgyf1m9hwTKaZFWFa
iOJstDBOCvqjuNVMko9rPyw0hVOKj5eQa6nKH7zC1KGdeiSHPI9qIowtrTGeeCB+
Z/xA8cqCFAKVOGhr/V6u2oQYmdw+ktcQXVxVhqhQkiD2181IKz+p/4i+X0MwpFLY
oUyZth8WzlNTdw3DewV2iCFRp5qG/4+la+CHzJQx8jd94vhOZgVLDk2u6BxONrBZ
W++l8YQc4QGnFr6bCivXRQcyp+4zYS/7HYVuy9ZcHJWDL3oczGvg33tScg4N7q5T
A/IlgOvW93yFBn2ZOAyEhSwdXc/kWeHvE8XJIYoOz+aEMAcrd9nL5CPDEge7MJN3
M+eQjpT6yBMraCcB+0gp9eF3rJGo7wK4tiphkRVJgxSxkOfZKiTKCDxcHNCP4z5o
PF/oT/Bt/aVMrk0Wnnwum0XWrFloiGK6W7NJNVU+e4tarUNOP5YUdA3F21oFiIVg
7IZ9nguydURQtJtRpdAnIDRqv30kygcDHkV5ELf0juLBYCC+pAADOMzCZa9iYNll
8E8PvWKVqQ9GGnPeFoREibN9xcPfYgSHb8j4OxgEZWF9NtGQYkHzEqu6JGaEgXOB
rAsT0Qg1HeGCvpDeDBXE1opO+3U1SJ9O5wdkzCOi8rQDGjIX2F6AuL0wkHCpn57u
Xmcnfol6wFOGh29v6x8d4kNj7Z4NdQ8DyZhiehssGopcR8tIVQ1jGb2I4xEx931v
t3YRtynx/hlNJW2tx8oLJFkA8StW1pltBHgIFzBvyW/GaugT439ptOHnwmdrIoYD
7SlKOlft5X6SIetPVoWJcpncQYw3IOnGMz0hjaRcme/odk6WF9MIqRLw4zyCqrwV
2cNvlwBr337lPl8gYEVm7Y6QNLjrmKuNy8r6DT4toYziWYodYB/ftpPj3f2npicM
6XYM4McbRa/p5ovdw28QY80ISLv5azgA7n1nKX/F2AnluvdnBQs9Q17O6xeD4vL0
ZXQetiFb1Z+XkYRTFDCrDX0gb3U3Pz7HVf1Mc63EmyF+cQ5Ynt9MVXoD4/ENfvWI
OHitVO4DGmIKDWQy1EOafk5o+F1jYNDoWu7VpFKnvbG8t608LXVEh0sTkT/VIT8L
3NNf+pTUEcy0hcGwezYOKO/vf+qPsI8ezYAOAGVF2OkTegeSBH+c9lWB0ELBG3q6
2rCUBUDZkTzmkxUVXZBJPyJZ94l3ccKzD1iBdwS56Rwff4yeKa/5jCA11eu2z2li
Wk3q9YbivWsTiuvPZwigGq3RZLCE/BO5xCkq+njC0RhCvKtQX0yM8SiiP3GGIEpm
gbpCqNFv7Nz+GgAzVXPNL/pWR3BHzpcCwU6Y82nv2m51PyOjagITTo36T6CNuv+P
zMsAQmMgzHSJ3zoDta/IwvAcxYbuz86+V/0Agan56PKLacje4/n7mdYoz6rP8fCd
34TG6VbX+91jG5XhnfWqcZmcSqtG8nVGwTusTrwX/zjLRIBReqRKLwOfqlm8L17B
oDy9z9b0dR7DeGzFU36xuOpcTb2hUWj/LmDL2ytFN3ydtn798L4v/B4ZXU2gNefW
Cb/ZM1QJTUmpONEWHr4TbMvCC6jTIME8nlTrgP1bpNPyxX59hGqY9Qa7D2kiWzcu
lMrfr5YOEZEj9HtIPTgvZCpQn22saWmouPpIBLLjB8zgxLqh/UtscfYuJwmT9SZ9
8YECpRUYJjUItY1zK1KXAUcap1iT9wnQJJtO1if1COeh5UiZrFdq1tWfCQktAy5n
wF+3gtgzhUwyeAWxL+eIzCd3qvl/YXIPKuTrSukWLOSXtaOiW76gdc/hIsNG0uTX
pCyQSXB4FL2nyYqHbDXcqKptU73X7uXPAWVRtG9tBIbWeBaxDir91eWfspRf+Mt/
IQOFk5aZmHkIngflICyldjODU4os8hgnpZtOTn82e4+5hcvHmCND28DnpxpZ75vB
B6xngVdwiecU183aD7MY9DT2wXKpEZ5AXp35uObuQoynWZI7ygB66FIWfY7jiSLH
tsG5WtnxH801e2+0gpX/8BaMcFjUVtAzw5cnpkTBJkEvZ5Vvj5/jb7g2gFuGDX2u
ekJGWvT5AItok65+lVi6+x5RMjeYc+vfEv8cIsg8SuimuH2pG/MplcOLzXQertop
1E97a8fuNaPW0kRsaV5JnRG7Mj9e3G/o7H5QPrSYt0gZx+gUQy+rFx6f4LbTcf5Z
YdtxMIBhsiffjqsdCUXSfBnv79SaE/QAcZUh1D7FDqxyfa5v5Ozf2P8gGFnUJqSX
0YogNQOMkIs9D8Gfn0ZDwCwQqtgEshetOGzsWZunHtFAlpCCW/aQI4k0o10uc9Vw
ql2LMZOrD9wkeiDxZknmmPhjXOP0WHreMaGHybNc/t93DW3XnLneDR00BJD4KaCP
VjPOeG3RJGbvhgglqKdjJU4bkR31+u18jmZzQICUqg0Wljm4AEDpqsWfFAwjQC1p
IHf/cv7sQ855uCwBOYwPvKQXBMc0bmWYdPknhSDM8n1vAMAWFV8TRTT2ldszgAEv
0q37Ph6ZMuQbB17pxYyu/Tx9Z88nSnbpFNL7Idmbtd6PoW7S5jYmsXwZVU6w3LXN
HfeQO377PfdFM960bvnvFOiyW454RSn1tVCPiqrjTM98LY3RC5qxOGcAanr50CdG
Y8wFCXtmPAqGEoCm+TA6laBEe7tbw7RzbVl/caG1zUCgHy7FTjkf9h1hV5G1UlJz
H8aS1KM1Oha/K8kDs9eY/TIRILJAF4O1T5PRhq7/4KPPkPlkgQsZG1wKfbRSoICs
RJplWE4/pFkFOYZPFc0/cQtWNMXxJJESg0esKL3AwqO/HmQhhSbOPfKJXtfNK1bp
FPm/hKpGY/m8TyN7jUjaZfaXP9OK3b9TZqbHeuzALx55dGGwEpPe3eepuBuT9QYn
kZ3ovQnIAKI8XMvbEHCAom3u3d0W9JQxUmoXZf6huJ6OrqO2f6PZi3T6MLOQnTtN
eCY3zYSFPUKovL3am/L8HwGJcTBc/cjUmyFR6Wix3wbvflldYG2+CHYnSHFvcv2H
BxW51Xe8IzjkjEI2PqAmaOPQPgJ7mY3C0jX1LPLwMTPd+3/Bl7b4xtj7J4kgLYWB
ktUg7DVka8A2NNA7o95cJ0Ww71P0PkHT56WErCn91KNHZ9VmWXJNqg9dMVCMcvwO
jey/bZJgXv7GEz99vmlHYHXlEhUPj2WJwMZDVSGI//tFV3n+OkiygmsGwWhN3LBM
m/Pzk0Nv1lh7npHeMlE4jvAryZuIinxMCgQLfXY5ccgw59s3ZwE94jal+C/WNdoN
Ho0ZqtsXL8aWxbATat2PbqknVtoGT8kXy4OlDgbU+EfxmzKmItFXeUZyqpnJzatw
rLjBMkXKXBxrrUY9CFv4g/+u00sUAlOnEP6oyxg4Ntfvv42sjvEBcQGRISt9BZGA
3HygC4zaeiI9mvPqCR1yEMcaVFod6lEzWtag/N0PAAWIenaftebBxt5vvpPDI7yI
PgS9irhTMEM8qPwryIy4knJ+/IXKTuC2nBAMRkY9vHmVYEVN9UPF2Agu+ESVloKc
IUqPq7RKp9h4Q/PMC31me527ijw/A12IvSsYwD7WUKH2neErhT0VG94oRy1Du9Kj
ZqllRsW00zKoknA2Xt60CgTPGeXJyqOHBGtaY2FvZqgd9IqF+dEKt7sRKcPUkRWb
A1TCAuT9okFXQHeLh3XveWXYuarDUsuYyUi6IjHIo9x9oWaJFnqwHOCqqw4rmwJ4
s5ASV03E920FV0q7syHJ2llqj7LbjOmUZgQzM3WhoPVnO6++wUjloT8TKydzTW5O
iwg+8E3Vkm+JcK59rQvlTSFgxzr1SRXkBJG/Wi8ItnbmwKkdWmXH7q8dZVrYC4qK
Omsq89oGOAcdhw6ST/lqpQpYTf3bkJCr32sfebE4GvxThrLpg7EBM0/imsDIw8n9
Wz/lERpfDTsPwzcIjX07t+jCzXYGXDHMqoTUYhVcm6iJlPL2Da5m4AQjeEV8NvKl
xCPux+R2A3lmKgHygNKAwPbf5tE7P/GKBN+VRG8ETScQCbXAnp+MnG4KAoVQNt6C
BLbYwkW3sJgPKDOKi/X87JKrHZFN0v5v3YFmSqtOm8CeY6mXRNgtNHKr2drFGPlQ
fN3OZQtesk6A7R3TPOcRbvHqUIdhXyjtHtA+IMQU3Ke/HXyZpOlg5D5L6ZhW8Zv3
4Z+ZvZMIqA38olBo9IyErKoMH5ZGK/fO2GtMaFkUxcxlrJF8sTXcpS15EeD64n5g
dLadWYIyg7h6qxBV6Q4GKh2xeqIP99J+nFQWU08IoDsAZRJ5bvkMouySkHZbWENO
Qse5uqOtPdghKFeSOUrA57nACvP03GfvN0RaS53CKc6yBy9a9UlLE97NvHR2J3td
w1e4en3VbZ0i0L0NEAwFFikgHiNawaoelJuSgoLhqL9z4rLYQgko9i3zNZjX5LRg
pg/fgypMj9jODUUNaJZXtc1YzVhbLa0/w8DXbm6BI+H5pMYE9Szsm8z+FEzFEBRB
q0A0V65/BefZgnFpO41UjwYJ5QafY8Tx5zFqtp8LDG4c95doeCFD79d2jtGrvo8z
4FO7uci/GSPByhuTuU8xGTPPzbMWhQXcEcyRVk5mK5HIn9DxG5DQEk1UHvEo2gkM
1QPnnGT9NngOsQRXtr4zj9yMSES9B3SWK6bNMlwUw2faQzn8n8GfxQqpH2/knrUw
kT+HD5bjzomPAGgv5UinebQpe23rS/lmXzroAucyFO5OAMKgFQ1EqZJ65SeSi2H5
xarbt81wNsOxfBJMAgaGcHKKDAWTsJ0+tLVY22cotU95HJsjIaK2lWNnnQmSlSPX
u96hKGOvX2IsK2tKNrrD1jCj/IqctoWvXkacwj+0sPGySUqTWn1pUEX596/Y2QEM
MOSBpc6hyJcQM7TF8K5WrGkbXTkgLlsfDQeFbpfguoEE3X2oo4YJblrqCSkH3tUk
KibOQ/flMMODD67hVvlhoN6tRrPh0Nf4I4A2kIYE7Tc5J8soY07lSgQ7dbGbMzKS
e6qEBH6+aHOeTBAfsbQ556vm+zUTkxCdbjrYxXEcmoBjxiC+XRPVzvd5IxKE/CeG
uyqur4Wu+9eA+rKHKFIux2Yo/ni8jMi5DEc3K7hamET7uxavXJscv5QiD8BMX2Cd
cu5C/ukcg8qqDM4AGML1QTGWZgVoUQ3+A9MQLOT9y5fHlKwWUqcXosyI9KjFjgWD
brzzjT1TzniHOJK/pOLKvgXI7dkH/FG/VAnXj7bI4ahYLyOD0JqPxDH81FM1ziBp
qmLH8dIl7Pf2GF/KS7kKp6+jtFJJ+wYglKsQGqkvSbtIsUEK7fiayKqRe6c3u2MX
Tj/SZp/ND9F/9mz9IVqRYkPWM4HgNm2QhwfH1Hoxhco5alKwME/lDPnXvAIUrfwJ
7gak3IrdRPFPmulHhIVdGNfGRZjGTc+n+oI4KzxFYYRkhQMJmLy75bcj8WvmfRj7
uya2VIEXmNtTmZY78JOQxWGgldfhMlx5tIzxs7+oj3jN381cUY8QgqxRdRjxfCPP
RqaDYVe0Od5BEW1xCTEtnrIu5h3AYG0XGrUoMph3kmSydfIbFqIyPJX92PoP89Zp
kn0ip/JohgZdXj4aksD1Ja4hZLvmSnKF5IPlc9OkKBWMMkApyUKFK00mO0IOdaYD
kt6LF2J7QRq59xZRAFyUtEVRhaasAXt0dpFuncDHpSOBGxjxpIMxWc52DVZL2khA
J/ebNMnnMQr9ns9MmIxa6/eITZnAaFF+3TCc5zw0bqkbDtCC46UPCCkqchffngtA
mj1klRQco93E0P9tmSfd6liR9dJfqNvPEAHK5+UeLMXTPiIFV+SFEAiNi3HT2J18
dnCN7TQyhAO5OejqQVVjbZlPLH1qoBoZ1uwfkghQzT/RkABdDChH8VfhUd15gKr1
X6cQF8v9dPcMzFbLA6e8eDbl+0RPY168NS06Puj4YrmAk1qzeEa55d0zra3/7R7Q
CZHayhJYAV3Zn8C3m4erCUXL+1MlP+SK1qOSj8zdcg8iSw5pbCx6VmXJAosUdoFj
RowPZKTc64f5JdOu/xn5VD2iRX5LBeVdOULX+nPi9g699PzIX5J3/nn8lRdeuDBA
OUUGXP32Bs9NYV+KF1Op2XM0cdAJbHq7GEEr2E8FOHYzSqzEsvby+XIz2AQbd6+C
lv5rQI9yFTVc7fbF78ub2cZ62FF9usw4j9cZXAsWU8BE001jawYJYELy7F/p8L7z
Wt5S4h2Ae7rL+h9AhBeeHfCO3Ol9GESxrgyt9wUBSY+cGI+xbnhWj6/+wPD0kptf
h3Ku38DC13CT7jfaNkukO5O6T6T/z/qG4AvLSYNGIFUND8dxLaX3Db0LPr7iKJs0
0wwa7E+v+pcVYWzsx93fmf4kxDr+OdkFLBHwL//naCVxkT6YTQ8ONq1HHUuxuegX
/I8Kj4nv8SRZPxgvA3XFtvcKVIND+M3JfHJBoBxXpK0havSjpPvU9Nrh1cCu3N9P
Yv9xyrKuqWBM0lIQoTOWUMZZjMZWURSFdlXGXTv566aQ+yudI0A4/3mNk7HqtJ27
bZGPdKPRJBL7mgdG/t0wbDjMb+FB7MI/ddYNRZiqjSGSV4cxU2pBI8FM/3woOggo
qR1qObFkKmM8O8LkAKRtbAPx5wHWWLhbdXsYsTkaxv05nqemF5dkQy6xWEhCeImj
KM+JvrBgcfKvnVOmqbbRcYDU1r4qV+liH2ZGiEENYMARKtq3j02zdWK29FZu4gy5
qeQHeliedql9+H1GrqeL8J2+ryCvmfefNAT27KxKrCUT7lxeTwR+NkQM0pujSjKa
WoqmobOLwX00rk3dgoFQ+YaoU2JpeS55Ms7X5wJ/oZwJwknaRxvyApndE+uYX+lJ
ysAr1uF1wxb/LP11vZYc9Ph+l8xYgL2vUjJ0nIX3Dn+P2V5+hhfdvPby9MJFZb1H
hkkMr+t8N+0F1OVehqTmoRjgyMzD3j/ah7BajrCu72zN9rENOcwbaR4FhmM/kz/J
R2MMbQHVxzqf/3bQiDsU/rjPjsoFirw5GOPIdJvOee7OB6T6yKdiThzmz+2nxikd
Jc0uqV4Jhuov4jrdXq+tvFuv4A90YHQksyiJTzqVuBnv47tYHIllieYlwx28az3x
qdj4CPuaaNXNvV6QHOf/PB7JWOydwziR7umQXJf+Iu/SQBaR6Ly0ITLTXUCXaZVC
V0rVB/N5R9HVkyYlWHEVtZvuGXI7m2Gi0T7QA9HUMBORlOBA2V6bjSZQalm3vvl3
Gv/ooGI1+OHNS1wGkTYv4eBmPYXSEnC/DOzh1+IkIBEdRdPiADLxwRr9Cmkmq/G7
+ZlUkI7/7we7Wi/FeWAjx4uND9R3pPaMWacdbZXmiKa/DPEyB5I9nvx6nVAXtRzR
0qPgu1vvkQskbVm66OSvEsnHOJeVE8/W00wH4/b8t8+o17vFA/4282eACU5faIUb
FjdoTbbqM+NUVRIgL3vHcG39sgrwku53rsV8z+prVEinDb8P90+xflcxe/5elet5
48j+SJ1vekAUgtTlAk8ZfuT41FCcSaNkHgZd0G5nipOnLcLKtMtIKgeV/PKdWCyo
E5P60d2E+orZ4nsDsBASxvWJi5O+/NNIEy/CYHTchSODo4d7xSL9Mb/AB7MQ7QGs
nZLhgLdjb/N7Wg7f9HVrrtom8zzikCnweRGe/NG+Q8QAr/OaxdbZp9c6reRCd2jB
dCbDaGoinz8hhLxg1aPFXh3mPCwAF4kAQ1tICLcj7vwd/5yeEAasRUgqXc3fEJXs
+yTbs9VBu9wWsRrYK2OyZXYUGVia+Mry4KcoiIvZY/AOYWT31xW53bxtf5jq3HkR
GHPQ/O73x6fXJU0ZPG7+liNOvj2Fv55+WFqBpp6I8Ylhu+WjVqk4FGfTznXEwPQs
tgnYJ446C8ebsn4sUYBwu3WjveZl3GWz5HU/UArcuZ5IKYuhBgAnRElvx5UbfxiB
aKJ5g1BIrq8s4JpVncRGAMtvnUTV78y+wkhThKguILJc0dTCN8+1tGHUM2UD30oU
BPe7e1Tpker7yGySHVtQlMVsfUhbsKl2/6lRBbnyq7cmn3fV0N/CdSYcmH4uLBGf
DQ4+ZPAnoyRwa4tgf5d0sk+VkCZw4JlQEObWT3oEzCLqf+mrMdTfS3nNqGa6IsY3
0Io5pRlznE407Ax6ffqlk/MPNPgvauszIR/dQmunAkPjDP+vUyaSDkM42nEazZp/
eEUfefQDED+pmegZErjrFjtnrvAj7lg9G1NrPNyB2SQUo2q6DCk1nUlEfbibRtCJ
hrhwtoRt/rRdjKswTB5Ybh8SkWWXFEWfcqjiXfvBs/nPSSgi6HtWUv64ZcnAOAkm
2g2XV8/QmGzVVuwJQ8Wma8FXS8ZeC0FFUyqCgUyMfzWk/vRK7QABPyQ/HSsAF57+
0jMJ+Ch4XjPSszegwy3EEL48IM2h3RSKn3Bk7O/kF25apXweSZvBesNelRnrCcTm
uQ3Cub3+Y9NMM8eeb77kkmmQTlgFQ+HLPNfUyUOliwwOHWQL01xBeE6ayP53SzEU
kdmovWG3iorqHV5mhtI5aFMeLOtDFhKKWjRN1lCS37pPAV9Scl1gqc3r3EjKrrLw
XHO8eL1Ihl8BNCL0yA19fhIRlJx3EF20q4WIYqEEfFFgswazKv/Lec0KD7fYE4dD
I0kxwAsvjoBM16YJHdcGFZI/D2NY9IFl8C5uKPmmC2RkDLaqSYLqIf9GfC4E+Lbw
GhJa64F0dCOuRPFCsq4oFUuqzfpPj6RwRak4xMMemjoxWYXAS/MRqNqo/CbFEm/1
4zspNQykgqYNZvwQMQcpjntOt3MHHQ/mexG6UGUvSJEyoLCIAxHr7fnNHfiJk7bP
G63hNnkqVzoX9IrXzuTTX4PyGLMgtWYzyBMmAZiUaVttdclOqHC07pWOQ2GBcbYj
yP1zLY3xZ6hVGsNhgjnSk45KJ0qJlDgxuAeocGYNpxwj9XKnJfYHnvX1mw6LmXm9
39VjJaqLLAw+HQhndmm6tlMlqk9JNjdPPMTWp345DQ8Qn/Mk3BE8xf0kuak4j4NO
BemZci9dBURruomBe4CAvCG37GHPaNl500CPJMY5ieACkHkV1TpUzdpKU1sWo6rB
5tgZc7zIWWyU26mBPOHPHxejEevBtzwznRUD6VumHBWDTCHakAdm/8iTMZHPCvs2
7RNpBGFD+RQW6sNl6eeN0YiBD53fMZmuZrlnUV33Pd+yHKOW6YVC5lLHpHTt5GYX
jLCpYDulqq+rsUs89jxku7sMeqLLQKyQoyY21JMYTXuYq3CkhK0WeekxjUkaF+wj
XR2r2D2ng/q7pAjD28IDRuFEoB08AJgdl6TnZfW5S9t3y4B+LzoFYyplWdZ0+8xn
LkAvnsjOY4lOze7N+rW9uVHd1lzkBMVxJ5UX/CD3XHVhTVJ/AAFoSlkq0Pw9vkjK
iNdXtwKrPq802U7xzvkPQ6ogBIFPLj+bIFiXjJz/7p9U5zXi4V9R8IIfkeFeKdNP
oRqkAc3mkRsWvyHBpTrW1lJjqms0FA8YjLOuaXZbrKy3jT2CS2f3606WHoHdl7pW
KRH3YVZs85QDzEvLJRaZV3BlouN7vTECPma/J0bM5XCZmkjfatISeGHI1GlEwHkR
3NuPUBQX8XR5Lw7XBindDQhUGuV9iTPxG5myl69LWurZsRBqszKETwOZ63YoY07I
huOtAAp0ORmg1W5r0ylY5RK+EV+Rz25HIF795XK2BJPGT6wMTpKLuWaeoc4VZ6UM
fbJrOX63Xeb+w2we4OKcekCJufa0Z+a7VI7/bSMEiRVX62aRUawt+ggpcOYHu6HW
JKwPZIG6xPHdOH5OS9SqMB+Qz+K7sXB8xTKo+gGPyHPbwFsvPcq4vRXVmqzXqez1
RaOXyCR4B4gOS1fTDVD3lUf23ub2Yy1lNGL7v7rMeTkLszICncv6yU5bAf9ScB/J
YuACcJkVD2om4geCuTPb7mk0Q+vkS2XHZDQv4jUKvaXAUQ6GuW64I589HFd8II/A
+4QFT4Yz+UqkG6PILgE5cw0QzjaMgRIvyQFnDjfsIRgJ8Pb+iLcrofDrY5jrB4Nr
QNHrAaWmwN1r2Iui6gCZCu9H2ZmL0uFeYdHAlX7iNhPNDayG6rUW550KYw02GAkG
FlBLijRlWdvH2Gb18lfsqXLMJgrnAPupuRZeviiIrNgSS/Vz8+2WInBBejA6fuWD
GCqD4Pye7SbcORe3j7JzyXD2WG4UfMuwECirM9cNi0q2ajpRmmtkETurUejVQswq
EBWIsGzdPdhtH8GZq1GUHezSd6Xmi9IqJDkzaI8M4dzPUi+elb1AClIybyo/s8uA
E3WbMB7Mhf78/cW8Ni/zbmfWqae6TFJKO533Ir0pfqupRh7kSjWCYLaQpnskImn7
w1qMdnAkuQ6fRmcarmj5TjxHsETvCz1GhAHPVU+mOTzTwfHNHi3CrhJ4D2dHOw4R
xkOAd26Npd9bBefxvTymEsy3wBCCQ6x0dICUnVD0DH9i5YuM5Fa0KwKuRq8ZYdC0
Ed50yz70zDmmqr+VXLWAMR8ob7rZft+tcesk/jkDcru8zFjX8VZc+My9SuHO9AUz
G8B1mgGHHop/xeTZkfXAAAqjphLRNRTyOLf3ctQVHYwyAfjQhp2OXf4GDI/HBdtL
3MD/o2F1EmtJCDjqdJZMTsmLdv83M3RGbc/FYo11V22az0yy42nPrc6iDbpb90oX
/graRtV6dmM55Z75GJ5z+DIrgIlh8+XsfzFZ9SDc0tgdr0KZlGO3f5EOem8WnGIK
S0gWzth333JpJCPZ7NMeqv5KpC6LiYetUAvy3PwVMMp7/WsbCtZVFHeXAH/5TsQ5
OCxSuh9pxhVazoBPgN8gaHPJyM9hY1nJ7ftqzo+zJuQZJ+f9+ZID8A6WC/j6ucE/
Imh/5HlW0XnsUp1HNhZKt74Vqt4Nt+WkwjK/J6RBMLCej4CD2rwCHdSinsatUMmF
pg9bkKyHGB9z2jVaq1JKGL+DtjjhYO0V0EiHBrCaxqw/TrH1B6KtcTvhcpe51p2W
hZVCjJvMdo8DuEtCf80NJcPNTJXrQivTrbMTvNhGrwNzcjznrbHAhCUSeOgbxcNU
Lc38Wk1KcifQ2i3pReTTkKSCHjBNyrFBGjN1YVs05AKDBYiGosg0/fUBWBDTAdDK
TAZkVk8RxmNXuJJx49bgk35hgqb2b+5KuV+wo+bUjKz9WKD25cWb9LAIsK4zLhO/
z0W0ygwFka8lEKVxrVYQNh2hUt1Ofehj31r/y8PBZXRSHdGuTYZtLwnxmawl7YjQ
BPmfV9Jb2huZh953uP3EZD8VusJ7/fRFDjOZdgm7bj7ijjUZn7wSL/JEeF9Y3CVK
DigyznpsbcEFByfm9k1U8y+cinpVDEMSWiCA8kiYCblOzIRUE4XYnwLDQ7j0EAFH
7pYszOVSQOVNAOec9YjNbGGb8hIMQk6xvz9wKdqsr6eaWG71em8jUM/BKYKWaeuc
XfO2z6IvISWQo9F/2V6fuHvrz8P1imjnfedy8L0DA/m3gOybdNXIToBlpxWb0QW+
POZCPQ8AYmCjqMaNIuveSKB6O828Vq6VWoazMannjGk9Tumr1xjB3kBXRfZ0kmy8
vZVNBDcbduKmOYzBvcPNQFmMCyOh2LbM9uYCm6psl7MBLOXwfnHScRZasURYQ0bS
nnYL1ruSf+FVV6EDlshB9Mt4lXkJvk6z1dblGlVuOm9uNyYv0EvoiWufTB81x3ay
uUvWzCnK/ATMJEpM+gk8syPS6qoapNmEF5cdfXnTAxkAPNtcDgdZ9rTEsAYFlbf6
aOpUU1wsz+vtEuRRFb9l/jtl7vbhFogsl+NBb7QDEUDLLH1ashhKvq91y3MleXq4
i8nJ/Og5xHkwqbb+WtiyvJ1pJmy2TQZ7HVp/cJIyRvGcukF24D0wIwkLR5j7Wzlz
N+gR29MviHe9wc9QiV/9rUl/S7uBIVGeyWEjIokzdsBkEjz0PA2AM5uZVfRO/lhZ
5SdUj4fJTuzVMPQjqDDZVDR4nmmuifCp+mAh1Wrb8Ihe4kNGc4AZSKSdn6f8aDEM
xiJMLKTQglxt74ots+6CM4XQpIAwZJjV0M4bGkDrMhLb3fyADmHAaKLMso8tyV5H
Sken5LCCmqf2ymoUA6R0h6JGeb+LkCl5qhGqIr8pCpIfROU4hXh4GEYMd68z+j90
VdO+K8hr40z0LTOetvBfAsqKKuRdF4phmI1t8ey4P4DkCnF02XJ872HmpkTp2H5b
0MahBTBcd1xTKV2Yw7zOzTu9BpU+xOm0pdNEtge4oYfOC+3pi109Zdc4vInkb/P7
kJtjOHvUPMLHT+ShnIeR4SKdRFH0KvZq9IiueMBpKFwwJbolPeElahCqUYNrt56z
vexa156A2YC/TVGKcUkCP/FufWYp6pOTGN5KkKJrOkF0DvxWGEbCj+kroLvt57Y/
T7IzYnP3D5eSCoh83vKK4pcfe7VzrtytsRKTx88dAWZ/ccayZxnL/twiqGMVeucq
FQDw/Zn8pkvDCBF6dkLPO7Zz8f11o3/geZG7CJMAlx1KOjKZno+gOoe2Zsi3yj2x
2CBsgVcmpV75iX10rnpVDdLYfcgLx6jbEuF9vwjzvoyOL0dnP0InFl4/eoKxq8Y6
qOMYuqOOxh7xeKpGAyto/NUsOQ3imrO4IGYm1kTDma1CYTvw9M0zcBD5HkqTsO2g
ccS7OR1cuGXBYSfIyxjohiuNXeZIgjDcKg624l2W9zxLCM7RrT0bsFXoXrRRPvcX
IcNpIn73BgRofP/nQZbs1iraOKYRKJ8i6F5TVFpgxBeKpC9vLxixAgg7cudjwneN
4vJ/2ZBzUmJTSBZm/FMnsOjDjzzjArK1zJquuz7BGWdRm3w8T+vuGKwExz/RcwCR
UqwFDRyLjKbKDAYvpfEk6cE9GlzyYda67r3OunTosQYbRT+O/lOya7yErCxaVtU7
YHrywcN3Df/kRSt1uLWMvgTKyuSRsHpdaRHVkhmX1WBk2iJDc85Kfnaj7lv4PS3c
zS9b7CVoO0apUbVVLmsyclALRC+LjtuHj2NwfL0juA+EkO2UFl3edDaGrXW4sMf1
rp/eA09rwyI3Gh0ScRNXBa0dVPdIhF0a1o3XlH8ye9bHR0WkfzCehpIrpCfsiLuX
wRCLuBbZDph5Ou7G9nCPoW6/45lXY5qycJ2kwMRVnrVVU0Vtb3+juecevvQC/AUb
VaHR68QukE8hpFpIOUyAO/ArRHUj2prMaFcVmmeSnPqXnL5LQpe1q8dDvd+yCseC
F4jv4CAGVVGX8JNqc22YVbuGYLDcBxBaTGuoi9kic9mJjkrVzwTAakKHmCIw7gs1
A3O3M/ejaQ77EyK6L1pd3UKNG4OoI4ITR/3UZlc8ZliIGMJVdaypAicoiWUyz8aL
MgWda6VStOvuzIyIYedAysI9l0mE+DmYVKWO6hhMobOzsBPEmBHpuScEmBbCjhJo
b8pthwxsfQcFBQk/+Kgcdtw15ZY3FpNj6XoKnE4+M1iSLMZga4ADPM/ICeUFM0wN
3n/5CHtreSsl1jB5TFrXH4MnDGM1dhRoQO0PjupXN8smiY1DzXHZUjaRmihpUp4U
kjU6jVMzrUQbEruV10Y7ZKjOLmgN2ahH+sBDJdNlhBOwP65aiQZrwKOvbpG88mHZ
5tlYvI1nRvu7pOt6dswvBP4dbsfn+xUVeq1RiAPS5RVbXvuUboL2sH0bo5BW0VkT
YhdD3D19bHwiq2N/8kPTLgFHIW+tTmWimen3IDB2BWdm81NiHiV3OnmPkH9vRr3l
rVIOvnuNCurwRNicSBocK+I0yykVifoCUzAHFDlrK5nNMC2caG7f90VussD9uXsj
rSKdkPoJU+tXqQyWBhNB1ydz0sBtRr4iUaGGBqe7lgaAfWaP8l5dLkqG6ck0bVIk
xo2h2Crz5kg9xpGikmf8RUipYB02Ktv7U3kl6ZZU16dfE/fUE6OaAA2HlR/H2Qlg
eBkPkKQwss5YUupFdD+jftN58D/RQL9zy0wJsPD4mgkZZ0E/X5gNQiPrM4RA70Uv
wc52QShnDQq8f+M9U2O2HsL/1dQKjIrhZdp3xTUQQrgeHb/MpRfS73TNXlmi0uPY
NmCbAuhyCG0u5P9L5uY63Xb7B5KHn2b2Ck88a3s9Ab8MMIft2QEqcCTL+YKTaSCx
k6aPf0wavtICpvCB0icuwYtGIy5aXyA7d3mYPBHjGr3wjc7yHSf8vhiCXeQazWyY
9EU4j56mElK5J92qtCntB0TOPXx5UbkfjFBr4VWdoMe41yonubLFwISTCJPWouvy
eD3mhJ0uzmSouHPMdvtPH3qepXRx5Ef/C5+k6rxUK9ib1Xb9zx7ihB/zW9fD/Wfy
R9kcX5Hv+eQkS7jX+9E8OtozQqr3TcZkhxK/BmAjbwBl6gmwYFONLWdptAZQYAci
OncEDe5lQ33bmq+kymKO5aLigk9K53ooKL9xb3nw7vxyMNhhC18/mj323H2seSWd
8b4woLXZ1P3RR0q1+3Sp3Qh4YqhOaVtJFnDzq5+1JtpStauP4N3UIDuQqQMcBGxP
vGEuMsLtKOi9n39NSgVcdQbDgPFNhL5WtJHwMv0aLBV3IgJFd9c9hZIcwptTHKN/
Manc0ttxhHYra+LV1FnTzHCx3CQGPRlL4HZjQjFwo8EeQazPUEjKztp+jyf46O76
LMyLOwJ0u8OBUaVBbs2FqRsSF3HkxTMm86PkgQdM39QYDAPxauX78eBJwFIYYVn8
Jd3LsHC54sEmk1KY0O/TQBgRZ6OXK1D/Xp5LdXAKsyJ9IG1QMlUx+dtrAOnJLm1Z
h/tNynutasvZlXqyZ17pWIzO8jxYIWU5crwTcg6iI+i3IpgRISWUdV2XcSXnwBrm
LjS9nzXcUREO/5kaNTK0bye1Pdo9cNrfzdpMlzrEELTifMvqIn4ZhehqNmDyq4DO
Qd71/W5acrXr53aAau1fdMRR/IiN92H6Azkc9aH/qwD9cmpQSVPamzXMT8utLxWW
3hU1ImVgCSHe0Lsxbu6mZLbMav/6kZNsx50urrhUM/807aJiIgCKFjHoN9Ftcgbw
XyqMxNBF3tX6IWCbpoT44bQkY9Ehq79tIvX6G6L90vrxXqTcClp+zRsnKZoe/InM
lCZJPqxUBP8THeAOPN7dcKn48vmgOHdlE6LR4UNXs9n81gPr++F/qHkT1FsCazZU
aY9QgwE9Xy5NSoDBGSSLz7r97Q5VrhGXfC1Vf3Squ4f7A5Ufyx1s697gwUtUoieW
IU7l++Hv+y76Cvg8bNMB69f6DLmLlINxaQlm3fv3H3V1iaiYT0yMo2a4TUTiBA38
oainnYQQvDdj4egjnpRfmTFocf8jHcJif0v3iwxQJk/YQt0ePf2uxfkafk+3Eb3P
elhHul+8ZxNUcfDSRei9K44CcZKm+ipnESaJNsqv0mrABHYcHMTmneGHUgrakduP
KFXmkFsrW/Yrsr6p/ZWmscUFJFrvFnnRTmCiONx0qMTU5ybPrlv4VfgNetWF4SAQ
Y+cBpCQIWVxiNI2WsHNI5phreSlkimUVZ7GZn/Zezze5D85rDh0M/pT5nPH+gLMk
N4v2vSjYflVCM7d/BU4SADy/WjV8Eo9RONSq+hEcAgI8BkdqP0k9qtbpwm2urGof
k8vzKbgWtsIKxeD4F6jEQ9AE0ZeueLm4Y79SQf0p+Yq+JsPKjDjaOBD4DFnJvq/B
Qaf8PrXL4+8STkGsrLiobddXu3ilzBwsZVpjoPYbePfN6XX1VudNzQnKU8D2CIey
Khh3dW0CJ864q9RvY15h5vL9edtYhUooFZwgTNPJp34zl4+eLkWYy0dRu6ngR03B
Ak82vaPbg3vWhjZI/k5jKTulfgwRWebrVBQ7nUIp5IMQPZstqRbZ/Cq1sovm3uSI
nA9H1MjOA9bEdTOSAJFf0jmSeqf1vlCJ6se1jx3O/R3lIBdWWOB2XXYF46fqhn0t
0pF7n76HeHbSf+NE5bri+x8uBGBs1gzQZSs2b0vdrAj+ySkTPI9KRuiQl2vSM00F
KYqS+KDwaGqpyd1TAAezCizJe3Uw9Mmh1355+cJO4IgTmnLznyyBUNNGBhVi/oPE
zoHD8gbbSE90psxHe1/12+QnZybPDidSeEkFBPxP89zGULwr9VZP6HkfF7X/qHBP
tw+NfsyGOrRoM9YMNzQZadxDaWv4P+ZNPkRprXUgSdZbYJ9eMu/gc9NVWau2FKvi
tQCkLDydsmk9mkfk2GlZnO2PicbVV++JE5zerjvbmAEJfOcyw9OP3xCaM0Ps8Bbb
LmmqorHBquk6TYeA922Rdt+/LWvAuEsibfUqKn/Mx1B9Z+G/5hXZ3hCoN1oYFAHc
7Cjn/Fh/XzcF/QenLdJOrb9Q8K/1HJ+vor5CLcgBWuGonsGtpgGf3UZK2e0vGO8C
G34YuW5c2zi7w5nqg66hkAtLQUqg9hy7fmhR7rKIadDgIlF9zL54dp5K+ExrVgGj
6RME3yi5WcD7+xGFebXmT/1CECmPS3MBcJyuc5AqSvyMUi1+Xc6mfeAJ0rRZt5MU
Fd7ssB/kJhnxBMc/fZte2K+u9HonIaZ9YbrApPQaU0TJda/BiS0sB+/Y+wALQuHs
YfqZ4loD1y5e3eGU9EBChb62Gj/+KHUy0lNGsucl/gEBlUyTWhKnfPcMUfbplzi4
kXh3ZhsPsU4Z/YS6rGtZ57bFSDY52XgTTrsmYvvD17kRDy1eNzP+tLK4cl9zKb4C
XjJS0PLkkE5ANcKBhcyfiNrKlvVahXAcFfMKpCxN7UKLj4cdlB9LMAGNgYqPZ3r2
kleTokS/WWyeUS9Hq08h/RJdYGYNqSeZHb4miyI7+JMfmHTUoKLvqDmIcJhrY1Lv
9+AgeI3wQELOyp3Xac8A9TYOa8wM0k7n4g98CK7Fn9pVG4EjRSvTMsgyI1sjy6af
VFLIA08nPMs6DNjm7ApSqYzdko/4B85W2USZ1GU8q0rnF+siu2iuwzmAiRmJAKLN
qSwb6oCqmEpF6GjrwqbjHMwWLkr6UJXDGKgdtQj8ksBgAInq7UuK0E2ECd2AfJtM
9OySN/x6Dkl2nVNXnBzkLbdGsn8xWHcVRh0ULbHOjfHQDSNRjZlsRk9nCuPuBkoi
nUM7MmbspCAYbz16oKc5PXNw1ljCtarcOIidGs2ZqvQap6d+x1XxfWZeGTXE4bkf
gh2ZxUso9c1Q62ptJW6xWghC0uK1vGJ1mt5Vndd3NPaa7tBp0B2XNe7cJjRFQRsw
BJ8rSJ21qU3K8Ybf9eG808FU+T9p01WLvONFtaTI8yu6iVVl+LYqtBc51gcZdTS+
EUtmHVyPKc2WRLh3uj2DB/19tlsIsd/FHZZWu1yblHFK3i6lFwviLoKHpd/9ShyX
U3SiWJxCoMwAgFaGmimc5AVm7ERJrxeC/ScHaenDK1uyR4b92moV6JNlVBC2/U8V
UkDADM/50EMZkPX0FWCnbYw84r6KLbOS2PfPviDOx66nTek932haOwQQCdsD205+
AQLjTQhMb/xxex4YqEP1ne1bnxwkva/kc+N6JwDPg48Xy55mFAj6G9fYD7stWKVC
oOhbRSWDzQzcQYL8ysvnKkt4dA5f7m4uMI8c+wsU+46MzgcjxtDGZF+z1fW+OAGv
lMhWDizrHRzAOTDNjvOw2gWkEYF4Z9q7867p8BAVP3pBEeIQ6514PLHBkKQc+9j1
KQ7uNOVVOuW5mzxjozmnYJyWeHlKTEmvYQoVdkbo396AEjvqg41EUNY1Z5cn4BlM
CBBMtCYkQtJUoFEZwjbiwsIvwczjhIE0TEnPMuCd2rDW8AFzSRKVpdsCDwIPRXjm
R74B6HP/Ic5BYt6beOcQpnl7dQBQyj6aA6alXX6YNisFZjyp4xWhmECXhjl7iCxx
Mws0mwHYJToIcqYLlICiq39HPzmDV9HarfPHdm329Lyenppl1VNjT1ldJDI9k26i
MqTYXTHI/kSYiUX3pIVu2BUsjMK2e72fI8lLhaTCSlvQ1IKyOqukLDFQDpdp1/R/
Xwi7OBdUpNDQuAsrCx/fn5ysjLLtAakIv23eT0FKyA7ysD4Eh99Y/9kb7/XikpyG
KqetXfH8mBNYJhn0kkWCp90rq+PqDLhfQ8prdiKT3FxI4sWfGTX096Cz8mhNxFtY
AT8tx1HyF6u6J44aNHBv28rTI9+w2/Z34sRi+KkmtuIkTdRUU3w7Yu11CzT3QQmG
Ab61z8uRcx5D+noG9MkG9U0gfpI/6NNiTEgWnR4Fb98uxxtvHBVpLerxdf1r8K9K
jYjzsfo27kFPcwI9tltCtJ6DdFBGkP4cITxBjNFI6jgR9rgjRMugyG5l+qZCkPLA
CPrR8+IVp8HhoJbmAehVry2NMa0SZF2EhzZqbFJWsIN9PhNOymfzoMIpXZxI7Erl
fa2ZlJXXuKobu9n7GYk+P+1acpsI2aHGSwSY1BffZUnqQymEio96e2Qf9pgOS/5Q
Mr+HU0kSl1APbWZdrMimFjB09vFbqlvo/gB2m7BEku/Sr2Ih6kinC9EqS63el6PM
h4rzj0RNZY0ee0Qv9YMoGYAw6Pva1y1YV6aihUXuk32Thxf/C4KvxtB3DX3qclnY
d/a+OR5Dfe9IK1E2uz90SbjUkhPcMKARnhnibEA2e/bBLKp8WZmbdLMa3iQ0jDGG
kcKeOcRLHKE3oJTWLlf8kDyRJinKUBKDzun7R61R/dHqnnAuqvInYkKZDc4erQ6+
49OmHk0I4JsAkNvFeFFMIy1fipBkPnnM1ACCdTfsa2Xql8D7ezX2kd2N+pHwdILn
G9YOtx4sly6tu+fw+8DUAK+p8k2pv/SVSWwEakTi0/FyVVQwQE8b1AhVNTthBW1p
BCFH2mCqjffyEh5nYcSokKjR6x1p2F2MGpgpPPu88WazqnLwV53n5KFDlnyRYMcN
DRV+sHJMeYmxvKAjVfoxYmHkL6Rfxiufp9tdsTfUdbml5rJQwWBmXwAM7KVVIn6S
xNJDpel9DF7hkHrF7rVAlUvlinTj5rfhhwgig96VXHgsDcaZcNPp8C0DmacjNXcs
VUjvru3Z6L65bJuA7xVhxcX4611BL2lhBLi3FshR0hgOp1c5snU00uykUC0c3rx8
4ISTrOUwtONj8WvxqGqqZJeR/TBtYZJ8n/W6CRuw6yJvFRlxMTl/vSXsr9ZHtjiF
5xI6/OsxADGpnziAnYXBckproDWK3u4n7iQWmKRgYwuIZSXRhUZH8qjNUGt8e5Jo
FZSejkcOdwE6lVROf/u4jRZIANlJg2iqBZj1pQZbyPLNoXpRKjMCbigesF0/bt7Y
dBMRbPgSEIIRJPmKGP1uyUpc4b0Nlu5sw5VOdEnFJJOYjaDh1rxgJKsnG7A6ZZTo
JQoctDwNWh6BYYzPean+izYre6PPWWuHvDyh/wFiCDfGyhZGxjyyQCLvmvyTQkoh
zxPZ5JicNe6Z1IubPv1cQxgkvdMrR152hoZlrNKjK2e2XVSmsUCTo3iv9JzSaSYF
n2Cw0E0gIA+dWatQNvfdjUJQkeKORLc+fCmvrqMEtrx02N6HSAdWG5aLpYARPQbG
WwLFSUQyrUjv81ZdSjoiVn10OZW/bMfvKw+Vj/bxl1crpa2gVPJRQY3BXQhqmYn4
253ZSpP5pXI1qgZuCoDOzqUSTOf97efGt0etGBYEqIrYa8F7aOz0D2EtGXh616uP
UQqnVmQfRRddVS5pDhhYdcvCGLM3Q2CaLRjrFd0It1zX/rTbJql+AGidvozmxS6I
i9wJs1vix38R5/6EsNIvvu0CMvypNf4OZvEtrGpVm0BLJUsY1EWg8SiCSiQZUAFP
WEKt+mObwzK2it+4uXLUGBcMzu37b3FPmMtYEw1K1chPFIPYn+kmvuH9ufTJcRir
Utxm4uZWz6xQJYKrh8ON81G2UB6XLPJjoNrhMp3VnO2gHcJJHBnqUPc2yo7abMBK
mtsDoLfIm3xPRpGFbQ/2/wsek4foPcbaDzdPf2uFuj7B1P3QXPy1qWedI+Mqf3xq
4hS0arnLccIdvww7n+H7tcACH7u1YIQ5qQTf8qNBGzp3iA6OJojOyMFdSafcoKTZ
ObzQy1YgwgBr6O9PuipSFcfbGTYcjyxcQhNcGxWQhvkzKUJzhkpvynavtAHUpKpb
kBJSoxf4PdOSQIbvsCnhGnVS/R2P1lTxtzClW0hcut6bLqiwMLchsmZToTSt0y0l
fUUxAWCRxCwi77MG+Cl29Jik7C3S8Fk/oFjakZAFwiRz12USkLBkxCvC2tUgxBwF
/XrpdDHrtIq7MXxpL2JlCMBoL6B8scg2RmQm4vwHdDmXReVV36mGSC1AVLURQ7dc
6YzRBOoxzdWifuwJ71NoSPdUL8azTVg4S/rI+BM7l+LRKDb5DzW/mv/pNCGYGAVG
/00etxrOucmrOKwr1xWRz9PhIn16nvF36onBGFTXDNxC7YRfcs+OF+f7hNuZIxcF
3U94eVE34kF0+4WGRchL3amS2Zy+2BqVm4L9lJg2Ta5amKH0U0AxExpcu4gk0XsV
2aBfIq7KU/grkXLhGRQSL12ndELfakHOutVL3YVnT9hcmIOZmONvhZPlx45gHV12
1lwVO2VWd7n8FGjZBK3xgAwE9ohCnbaB7077+T2pOPjFJ/gkhlxSyLqnCPeJb6dB
r/DWmeptqUjZcmt9+4o01ZrfE9IOrGbZeLWP3c8txSEu1hwTzJLNBumiPhuXLLE6
uk7ivkMRbK/EV6hyu6Ej4Bme2v+KAGpwCEIU93cW8B+1ojxWSVNkjA5n9Enw0FzX
vv0qY0nm7jEJB26Qz8lnCH068CLk8NMh6Z9S1k2+/47K0hpry/NZma4Sz1zG+Lcv
s0mIgtrDwhpZfXKLoKV9d3gVJ08Mc+jQlg+zb26xE4fni18LhPKp7YucUAEg0mza
E3OBHhTakPBiqLLTi0Vo2a7fBXSd0NDTSsnPCkpiuCh4VT8tooyXm0JqwvhmJvq4
c2YTl4AEiBh9ntdle4RiEcT7dFSkY0wmmAqQDCh4dCDVP//HWWroemZLMphuzfiI
ufWUjzpdCh/1cqTNIlYQUWKj2w/Npc3z89nHWPV3TzZWlf+lj9BSv8eDQgY97uWZ
UrujNMk/UVBQuHZHSN1zxu2VcN4rpQDZXzj/Z+Zix7vIt6xhsj5axBm6P9iRm0vo
bhq+7Qrx3alGGyVgbPqI2PQ7s3K15ximNYULH4Ofs6B7h4TED0lk7UchQR/8UUAo
4aSWGRMPVmmrL09rrFb0y8RzE8p8+Et07pI11AU8BUd0AvYvr55T1xRhpQM8fgwM
9a1h8sbETYXlQN2nHDjYkW3kT7fRkF9PRVcO4T1aM1GvpnhaeJd9gzeA3gQKu8M0
VH3FeucE7z0DZRTKNPOZ9I/lXza8afGkjl9qUm77+9MCf1SJZaK6vFD3rU9l96N+
aZck3svbzxVqJbAdZpHBVAqOa+YS38tOrU3mf0MtBcqEsjOmuD7m5akHdRrIiF64
cbsz4CsgnxbvbHNVyK+vgBphfuztsLoY7AViX8hg2UUgKaxhG8wbaVUhEQROOiRO
B1/JnLhctuYXJ/QwdQR3ePKrUQt2k4wMj5KbkZn/GV0jeDUbtbS1qWe5W+Kizeo0
QOHos2mDk2q+38zujiZAs6usjv0cCOr7F2hi/oFLVsSLuBFGARSDwWzs2H5ZZaQe
WQXlvX87mVoQqK+DBj+ZDY1d35/FHK4jvmVttkng6/qRqk66fbWIgkUpsufOEMrl
nvmnSZVgPLr+dlXRZsK0h+Iv/IWJ35h9IT9yzX9Mm+s5ctyPo6146+jnqW8Ar3Lt
TFcpD4ouHTH15I/mGsBp+BsPSvYSNFz+dcZzja8eknmOQd+0xQKzyShzdWFrQhR/
6QAMeQd/WzEL6bEUIyfqBWkw4SfwvHJNXXRmtEK2tLAG5nttAr2hVPlBaP9GZFxm
6w4CrdEvlZYvnMDsx2Tx6zLEysbtfsZ5QcvsYTs23wYqyAcFWnrZko41QhV6hFQV
p7oAlMLwRPavplmFXZtJwPbfsTUfR26PHB0R9bJD3e5DlRLr8HaZ0bsb5+/8kPpN
oTD5mjuYHMC5g+jM8FTCWbwh/ZJlYIoKA9cawlyFYSwm/XrCDnAHFrOKPUV4lvCP
Jo424DuBx/mIxBnx2LlQp+5yHpACQ2cWGvVJfox3EaedMkndlqA1UcWW1U8aqJKr
Mgd0slL2bCnGQpMDkgE5fvitEN9ATZ61IhjedviRAT8Y+r4IAA5pYc31uurTpxt1
Gnc4HWmuM4jp0UMgS5UjGLZhMXb2jvs7mOtf35pM97dm/ycURsHzNU9Fpd4r3nMW
udjRvBxq5IEDx4qgb5+4CaPJlWL1Nv69Ex01VYRKK4dR9uND4L41Ui3aPLpvzPg9
0kZvdWuQHc8ifKlzJmQ4iG/EtDKjvlURBYe7K6ZQmWRcweMggLvuNZSflcG6dtTh
R1JqG5kxvsRKKlQmBIHCSXe+v/myjORSgIfrW61l+6Yz5R3Cw6c4vdgs6AM/wZQX
WqWBC3D2oC3yQX09GYp06QAGvcesmlZgVJpA8JciYft/WLQ6aEOIFPThZngkyPvI
lkzzQ7vlT1cWciAjjTpXvLahKQth3SiLoUKRHvJuOz5xPsMswgef3i/VTq9NCI8+
CIOxsNz1xjs8Pcxb8pf4Nitf/6Ya+2DQNIMvE2BeTMlm55joOwjYCwvW+CmI8gC3
ftzoh1YsvfOiQ0ar8Pj6uOZurOPZRdHzfc61s86Q+vmaLGD2xEMq5P+1s+nVCWk/
uvB6jeHQxg5nvYY5v+vsmw/lnqTZc4ywrAKW+uewd6qCxQlybj2Nt88O0PytnE+g
6IBQRw5Ssuu3JmdxY3aN92Eeve+HJgwsEkDUQU899xKJ9vw5wsdu9Jvp5B2/12nW
KzW03O62Lgv4eYet/Bplh57+Gzyab4IhPgXjAAlkwSmrLPLVm03ZVMSxHPqquPYP
h2DmIRHtMqjDLRTES/x8XWIg/P/4t8Nk/Ve66zHe53yfuyYTekOq8XwFGqGQ1p2Z
V/GvMOQ1fTL+fE8d/6uqHOf9J97NiYeDctUmpqbXuPdowgPhZwzIoGr2oWGBQzVg
ZgJEBvSfU8heIH9VerwvYhwp5VocrKrh5efkeskjGKFUXDFaxcaOmADBHf7jBR9n
vMg9BYGVTF9hhxSi5j/UiOIjjYtO0/y+IBlKcwOuCQ+/f710wGLAaSOKNXkbgqaT
jqZLlZKJfHC/BtyGD8ZXqP96Cb4hB0S9AD4PWyAep2UeA4+63HhWdn5J9/VTq2rS
tz3TjCF/vwJdrPE3D8+I3HHWc8xzwDdy26JyPO4xniUz3JGNOLPstI2Z5R2iz7BB
bKLI+EB9aSdhwRHhyEeM+l+FzlV3VfuIsk1Qvg+6h4L6NM19+zO4T7FBAuqGqEXb
ZdxNoylc+5P/PFKIB5OSeyDxiHbNO1Af0Uu+ARzaz7dTZ4cUeie6e2r5XyhMPz8H
6GzdCU2i4a5c7CIZyS9c6Q2C/ujGSRwyVKi2PCwC3xZsXeNTJdlrF9+BDnqfXL+/
XYjqB21UK4v7VYh2Umgc2WJYmHPPOo8nA2TS16Ty4loGydz31ztcPdALvim7zug7
UXLc80l7n1q2zP18Z9rCf8x5+jlmRcvaEll7ewF8gHwg0UtmyGoTAZsXqSqOQltb
MBzcGKLARB71sKuvGu5arzfTR2wuyakBUqP8ap6GvZZyEbFQYjZTYEk+VoSLqRdn
sUjz+OcLrWdJG+g7vyQUfgohTe1h1o0aJLnGw1tC/A85C/vrBY9MiFUnNGycGb0i
erMlBm2tOBeriPzoSfKeP/FXU2YV3XGX8lCGm4g6IQtQudw3yKE3B5rwYA790tFo
BD4r/2k1qeaxCTJ5W2U6r+BtfOYnp3U23BINM59ZfTJ9Z/sDi+bkpzU3UbJiEd9I
IQVVj8f77MDyXtGRkJ86UUzOdQXYaBsX6Le5imQG5sbvI9rQVy4SWRNuF10W58Aw
hBDGn3N/iB3g50xr4mYHLPifBabk/0yssV33Trr4kvcteGi63kGK8xKrxgTcFmhf
Mn+5xtGr1LSVv56kyGA27Jg35uexMCZLc3y9OKWYt9YvLiF9FqprQ8XNl7jr8Y/d
zv8R6R4c/VLb3O1OqmKyvLdojxzL9mXfXINJLwOBTOtDLArzvoRrGGqJtK5oOk2/
t+oXJH7VE6GfuFwY9hiU6lY1beXyn33SIPysLX8c190vft6r+i9nh6W2V5Blj3vU
lHZzz2bDbw3eBXgTwJpHgCHChFz1KdVz4iFBt8yUVfBMsgGmkinyPmdLdQwUB0s7
6qTf1Rqy2KC1BNhq3DIPAyu+idn5EVpJ9aPn3/YarS7JZdgEYCZfg5gUucrRjVZ+
MIZb77ndLAVrU7KNNKi9j4NT/bj7RYDQ9zOdFqQrdN8ohBdiWbeSi6zdUkwsqSzR
sBkBdFY7cD+itliDEfD5XNEdnbC4hwxnGDjTRHdwGaJbmnMwP0QMsKK9aD2ppR/I
982N59QLeWn9Ih63BkFtSgoyVa5DwaSQUVE+/JsJQiAlZAX9nLR55r9IKQLkdiLF
7UxYMdfkPYv8mScJHnmU3On3PTjgQyk41fXlbv1tUp0wwnafyNIW5eZsOuy1ctik
HDxF/YjKQdf5Eq6gXcmxl8201n4w1UzVla1oq2QNcNq6OC5Js+nA+1hisTqORAgk
GqBzA6y3dN9YiU/ZJndHrs/KbxKaaH/qA+icRKnVOMtKPcjJdeVjUFh1Dl8144YC
+rAKKHVghhBQjVjbvI869jZD0ZABO4lj1TI7gzZSxwwNxQ+s/o3FLcCWSRKWF9mr
N0LHk2ndaTVFoLpJdkpnaOyNITtd4rMQ8yqO2p2DBaqQKk8+IV/1JukX832rnXCY
uA9k5BioWsgWxytXSQ8CTI2q2JK+HwDhgvIQzy4CjMVlPynPm7PtQsgNrdP78AxT
1QW8LDhRrbNseDM8lU+cgTbKPaR8KLWKnV4lBgE9TFv6DVZprpRGJit1219fiAhH
vL71TziDLMYLXMdOLiyzmGKCp2lldtLA26MqriocUZrqRW4VmNKqHlF5UqmzVigh
CL7EGIljs0nqqINSTL/xEVFhe3MlVbzqh6G7zAUIB4OXVxNu5IqWOcCvfr4QACss
PQQaz2FgQ0xJXRF3mLckRE4GJx6BV+prZn5QVRL1ajRsggmsxluat0pBW5BzqSxm
spKmL09anxTv4WtU9P52Bbu1sHWNSQzNVMvZROmnkS8kwKockLP1HucRxAYj+Oyh
9GFjEaXSBjHIyt8gRzMYyJz9OGISTy7TXMoqkv2hmDiZZVp/iX0wstlNgmsMhT1k
SFYGQtCLmTYJ1fL1ddZrB19NzImp1M+aI6LvpBqP6xrH7xzOEpHRxfHnV25avamF
0i442wEf+OP3Xrr1uUF9r7g7KkI2oV6FP/lATo+2mzMEzPiHFt2bNr7LrWYIA8m3
up1JvAr5lxXu9Lq4PqD0rXb/fRKt70KGxq5NuFL4/hboXpJvRjddn7ybu2dmDpHx
FcPMLOuS+6wxC+yWCxy4gbLPFkmPeed4TwIHI5WRejQuLdIpUs3F0HY20M6C7Ndq
pPgIvYtzpCkiMtoi5ERxBkh079Zr5Xek4cVMoXgShXiM8Gl3Yd23pxbwD/BQkkzc
BodhsPKDIbMvMGgTiOkJmpOlECIZC5Dhc+l1pQgoLjJLRPAYj1vSJSYFbCBvWdjb
iVXsOtr0u1hBGufHfgC06thmY4xX9XUQck4BHooBe0FfBeGxiNkwdgBilB2F67j4
UFECVYdT6zGM6rbuePdWR4WH0kdS/4O0hoRNAE15u1LtU7ztHI8+wsMNF/h0vnr3
tHSMLlsBLAIUjAVGr2L02K2Mto0yxWffKevpYYhv711VhTnL7oB3fk914mR4cSKW
P1MwXHD3wtpAfuiWhhaH+bAZiQ4EV+abCT+xUm3HCsjfuwSWU5zOnVAyQeHB+SWI
apSbc49MNVz+85OXqdCUhgRybibJYlXZPnJ+1GBxrLAw3eV8u0RGJW+Vf8kjivf8
1SK7N0bY+Z8H+3vMSbOpdxLqObL/h1RnvTaCxwroEsP+x6RKTuqILs2o7DoHR32r
pMTK4RDKZQLtQdZW6d6gxskHFRODqjkzq6tq2/7jEg8Tj4v+dAV1v+POiWg8FDPo
LOEh3LFcakv7M6e13RrwiXsoqiIVGrWNMZMbMI5RS3ibp+gBe52gWiIG6OhFAae9
9TFGZTHFiUMjsgfsLrSQFenF/gS0AGdVvybxunf4/rP5j4xfjDmJKP/r7djInchB
ROmOtUfaT2B+M0Wk4jGdz2VGrSIhdA/a6oiWx3a8qBRWby9Q5Pv2ktQdvnpHytbm
L7uoshrA0LXGJB8kvmQKNH7EIQWkDYl7AZVEDbFyE659DYsEAr0/sYLlZGdDYfMj
ydiJ3CHzo7AAd/v+Oo4NJ1fzqmcA18eI8aIJ3iQWBPb6KrMMBt9ibaa6D9K/Kpsj
+NZQmiWohFEBCPKylU423Je6hU4mEv/vm/dIqZFzzPtjBmeWburPu7bBpIp+q+pB
YfbzddxuA6Yh2Qg+x2BoGlrTq5sD/0PSOEXh/yKLr+h0THPv0MaR9fMbTVaVODoq
ObZimFpV8UcfZydHW255rUmMmE3PakT8ckxQ1e8qldCutRxZH5BLD1VqjqRteNI3
J3S/a4uvYuy+IC/gCoSJvxsIAKBlyJ8tTyJnJYwqkfCqvE8bV+gpvYis7W0t6G9H
meOEQ8aJ0phtOA9nslDAe4uJBh/PKgglp+a6TgHnvkhVvg44BLEpynd/CZ0FRuuj
aeLNUj6uhzvnvC1SB4SVEIPmXsX1OvBhOWu/W0Yt+LTCBlL2o8c/pv6z4EFo6Sr3
7bM2pRPcsCuLAOefSQ3p1uuBBs60DsaEJrsiLCAif4VaLapVUAktBsyedqtIISwk
Qie53FfeLByKZIGZmQOfAG58Krhss2dqJPhzmVxTZOjv73E1V9XN+LG8hSh6+1fo
xZN6gkhWVLqcDAv3K+pXAdPGJ3Yiryqd8ivLLQQNV4MgAkR7k85633AAjDpm+rYW
kM1hj73FAbOueAyJpHhvv4cyuDfBZmeIaMh4VkBp7Xz+g8wgeWv0EOQ4bvvho9jq
gfgYq+LPa4QsHgyLfClIQsi142zGQzNUzypXjgKX5cqMYmTQWVKgTc7krlwD5DG1
Qu9UdDNqudRblNSD9juKHCl1iokbC0l66xpstnUwiyvJS4BU2Yo2u1sP+vWjehOf
8LDkyl26BrKCaSAbf7FW0UlvYKg+ivzPi3fhbDb4nFj1ZaR4C5P70l8w5KVmGPgW
l6WfqAq8RFBS0/DbQI4L/xYs70zBpnv9qQPoqy8BaAiF/tx7gEFdz7CK0+hw391t
ysrvpAJ2Svweyzzz3zI6auT5iDqPzxrq0Uh7NBd85MnIAvV5O/GQvpPHspRmmGUr
ohEys1OqiBaQwZsjjIT98ZzmtNLttpWXzqQkmKI7BqKV3x/ZIDb4pZi9fC6Vf+yN
Fl02Yt8Ivog8VwpxPWljQXAgbWaSm7MLkTg/uV//JyTmrcH/ufekXgsENOM4jXtf
dFlWVwgTQBwc/EfqpsQjBkDxNu2sw0gGEgTMQ+tv8PKx6jolpDkAbehpGkmCDzM+
2TDtNvOSzjPIttGfXutRopY0zSHxM8Mx71gjYrb4Gn3cTfaNbXPTIxRqs9ixFtZK
ukCIvShnlz265CfbvWHkwsxm2t+bJiy4f7aXAQzUywCm7uH2TTElNt/K4kAS5Yr4
pXmnT1ZtNuTsneYKX9QjOPjvLe5h2DBlJSLQtcF/VPD9SFmjWGjDJPwWDmFu+4G/
+RUyoB25/C2S1+xjL8HqHr3YTH02RJqdn+WPXz/tukoipMnTBungpfL8CZCZ0snS
KXyiMZxksyeUH0iBUMNnrcRLMempBDS5nLLVM1FFF66L+5/gtbGaeVO7Z6s6I2HQ
DWzbzyLLRbV/R+vQoxr2UfbHKpDDzuNNYWoV4zsVAruYGyGhS4LqCnc9V/urw5Oy
IsYeZKNVw3FeZ5VaBN+Xg8jo641wL3IVtIv0TMNgB1JLtvr8KKLC9i4FDJvmnZqH
5/VZYQRt+Ha7i4e5FcHJ3chGGOVXIvBjnev6xHAsML8o/6F2XdxjiYxRTKDQwoj5
UrfOlsofWwdcJG6XQrB0NT/awYIDohZm2Xxj5jrsj1pMXG8+j47YmboFy2Lh+J3Y
8mTbkRA7pr8uO1v1QqY0EpUkiMRmYAFwYgL/YEEu92xd5yXD/31QPl86f8LuHYuB
myIQ7K+E58oW7u419eoNw8OKA27/8Go8MNM0boc3BfSJ8o9vWpqej1FZTeCWuvtk
zXuCxXzE6iDXlnZhOyQYdRz5DympTuzO0+CjaFCCDQJPw2cjzdiBIsL55a96Ef++
VH/E+u6tDvQmxwcGfPpefPVwEr+w17yFlPmoUVofSk5Vxhpb9MJ/IHSoSnWhUKJa
q6J6N61xpy1XlQieoU7eGJ9Qs+5OfrVXkVyX+x9LdQ7QRyPB+P3H+IqpfH2hkFRS
UjcAX+HU/JrYZRKMHJGuT5EDyyFer/JEbQ0EKyZIOaoYnrny40rK7g9HsrjZgvhv
0eDbMRLmMssd5dRGSuHqCRGEEH/O86E48sHahSajK/C/3nQ2pDIm1akfpKnFDrZ+
YOBmDBr0kE589X8AhArRq/1GzlTPpCxOnuPXf1/0tegYChHtW/cCsja14RjpveT5
tqi+6TJSM9MUJSbjSkwT0EwslSz7C2OH6Kl+A0rcDEqbHvQxFFcz1vYtRLrakqnB
NQ2rrxRI5+ym5qOkBD26hd3Xm8xZMtVe/PDB25/RwAMyWICHXXAuCB18vlF4oELW
62fgsQlmfn1ms8MGmsc0ARBdLEWwE+iHaU8bRJKenNRgknbb8AurBy1Sf6GRk88W
qv+BUFBxTrPk7qLiZSkuJ6wqnixnAbrLmJqcQWAL5j6CN9qB/mXNSE7Cd3kwvC/G
kPChEOTk/UABkpJt9nkJb6kK7gBmpbEprgf8hjZfT7G1p+l6ZV4sep9QiafEj0mI
HGGTV6eevei87cBhbedewa0u0+35aA8wP60sR5mqYuhq+/t5TpWYozsEzd5LktTL
42IBkNhP7/Birdq1wgRM8Mv5dFcg3iagAPsz5YrSDsGlRsD9alUHiAHO0m7pX0SN
+wVVAHSYaCwsVksiypezoizs0ajDp3zkInIVOxfsh6OKCUIS9iFFyWTGZXFGIG8o
nKjlqbvflmFU9RGJejwz8LrnAyR04OT3zBvz2lG0jD8FZDGBLQNsbA49pQHvveWi
+TKBJpxnHNCkVIw6aZ8HIKF5YDsVVwe80ZqIA2KpYS401cNdqQK+SbKRUJUhkKvG
09gqCjtithHIdv/yxmtQ8lPDIkBxZ7OQ8brLlV0vznf1FgY1UCh0dRNRatO2GTyr
9PmJWOAK1JBuKjAbyMxBjLhuUZ6BETnkLqixIxwZMeqeeigF9C6KYmcd/jl4PU3U
wF6TrvjWH3+RrY4q4j7NbTy+GDAl2i5jjx1qRZzIxrSLUzfVgHrgGHRm3YYVwfUK
8/LclTliMiLO2rEsrQhWm+EIl+xgbS3sn0/GLg5oKtv2YfWrRgCAjVG+KXIRSAis
YXJmm7utPtJOtOthb2d6nUu3ZL37xCiPRfdbeeqlm5oafCPilnXpPt4BoAnb5H5+
wOjQ/xh5/tZBmfWdadoMG1BafzXo/m0r5t/oDHYVGgPil+4gYNhcuoyXq7lZox89
Y0RhRLRNvix8xcFoYpCqgLrJS7s2scnjioZnJwlfPeVBmv2lUKnkNszH2dK61am+
Rum7Aat4PN9q8sYPUweiwaTtWrrnw6Xo7cSj2ojkgxM4Qe6Dg6JoRVrNRIIVp0ej
fzGlZPLk/vnK6xG7AS68WaCDZomywDFOfZB3Ny/eKVQi/Mx7E48AYhGQmDpP4LRG
IARQRHAl0kpw7sGo2RZyxhE27ojhCd1exH2ePZQcD53cMvzrcGNEAWMWAOSgK9gs
FE0pvolHXcP/jy9rwzzzqBQ85emUY5ynSRHMU99ZpgD/M774XZadIIRtLkDYSnFG
E1rZ4gSuI2x9Gauv2PVgaYssdSZlw6aoLem9PD2CfAKF4FYKMWBCrA3nkGtpmNBd
3lNOgKkI7S0nlZ/t0VMwR6YZzNA6gneHvhTpeee5Rjx0+Z2f0ugDHu3rFppPHfQP
NpWH/MeFocW0Ro8wJ3ZgJmjXSbHc8D3FTwJyFfYtU4nBCc5oT+Fc6mcxq/JJisiL
rQS9AQMSz60mb/hAqDPOnnJsoszgo2ugfLsYAwHdjDYmrbJZIbVTmN9GuKvVs3eT
9HoJRke1j/0v+VxoczqaozJbscx4AHh/gqOnwnjeN6XUJrJijVMBxdw4Nzhb6+2n
CkiFpm+3oBMuV9HvJCcgUEDipM98gnGDJE5nQJ3zQVdcU9lhM12m5ubQ6ljYR3lc
BrFs4Va9h9edss7iwHQj9hTI7feQXsN7TOmb6pURsiNInnkLQPGLR7Ozka2Laitj
YLltquAcVET+50b1ovOH3KEB6GqDcJIYdUeWcTPoepLPQfSP+/Nr8vCdUGykbWtI
OHM1saUoAXzJdUt/67MD7vyR3YsgAkXv3eW+P96ZBF+Aq/LBE4EP8cx6LVifvw84
rE6hFc7dTC1VkRd9Rr6PZh0R9mZ6gc9vgS+tgEyCCR4h//UDGOG0tcaTTvJYNioD
8VLkMWdDuaPVRl7USJtIBcgYIiHgA5ET7iBvnI25a9mIqk3wcm9wOHAHF456hx8G
uFqyHlHa3xrogDXRRnjOVdA4s6LrbsKTv7cZqnhXr2U9Hz35hL2S271W9BgjHUKd
Jax8FYU0Mx33CSYK4AtUiTI1XgJFxB2JEAVic1FX4daexaCYsNAp/Qo+l8r2o3pk
Y7AhXg2jrclyX0jmmQyREKME+3HAvf+qlXO488jMoiRv7FSdUBIu7UJXgNTEM/2/
ipIHOrhE98ujm32YS7Zrha7vniuWs2yTTb8QluwBFQjtgYkL3jmuMdo1ma0gneq6
JrUWt7zzP9ogOv8r+Dcw6hhKePIZkvPPChfUWGF5eh1jKDSbMYhvEPKR7sSmc8vz
ySPW2eH4IOupLTKEhjyDlELW0cRy/b39ruu+BGtZQ0SAgxqi4IwttfxFNpdPOA6K
rxUZx/r1MytAlvhorOUzqdYoZ9oh5059gvyz9JMOgZRjqrtGi4u4c/BBfYkOnyus
xil4LOvhCUzDtf6nyQrFk219I1QIKoXb+oiKE6TsmT+ZeRfieqLXPwZqUKIiHKyw
6cmmyM5XR2wR7Sd9NKbAZJ9arjodak55H2WIHgMpzZUov+qQPVyQ/sOWiM3gLV/V
IV+U9YSGQTkb4wEe1/TFM/3zdUwqG0jo8cdtkT+Py1o/hAFN5jCZlB8slwNlHRBm
jJHtXebUFznTG9P9UUvnD6dS/TyW3HYEe8VYuFHBNA4k8/jf6k3a/NRCkFvvSsgw
vGsla8f6PcBxpOY1ARV7GrDh584ctH4ki8VJsbiqkPAYMnicQM4QuH3QtXFoQJCV
7cPJ7147LgYTmXKhUZ+JFUykk5bgzN/odlfzuekKrkWjwy5F0SgraMtOtn0OOlV5
N+i3PNHARm4Ev1VTe8FkcbnC6q3VVeFgRrRu+rmW6rYTW/jETllck0jPOXoxz/jC
Da27jIGYShOj4t3xSHJj9neSAi4zPu6dI+qWfGb8IcajKwQVmR5AT1RX4HO5jqrC
wiGFaEQzJapo/jAVpERAbeHflx0HSzHzJX0mmnOXaCaCTvTK1IuZPmuScmaN6b2B
BLHF6Gz3NxsC5ZdN1ycbkrh3nYzv7+SqIPK4KE8nifc50Z6jFk8/YVg9wnNlQpjn
dR4Jeu0+X53kVicqDmkJYpFHkac5S/rZfALxh9O8BCdK42ztTI8cOp1oSEh+LIk7
otCsAGAFxXhaKZ5OoMlwaOhDUqQEF7Utmyps3LqYicjHDEe2dLVqh0Op7J8T06i4
3InAwyABKocRh4kO6HXCqKuuJeGjEmJUqplBy6bSHCyURTS1y8CilSoSIFOzVcql
4glY9qTfybd8dLlNFWzISh5CBuy3ayNbJggzxSVsbx9bZPj5eu/uSNvC/XZBGT32
g/8YHAdW9MemBigOoY4eBW09iJVJDtoC372o8vXwYtoli6mLz8m2lSz+7adzI4l2
B69sA2mQc6KOO7xswnt10Snjk7agtbiHRhBW4pth8bdYQ3w2IP84dGY8NZ/rP/Zc
Vo6qkLEiM/H3mg7xNTohJIEUTD0pbzAEc2cQ+BAP3ObBQWcvrLhpBVCNgDHAFyPJ
Yo4VX92+Va3SizviZXF+huO+7/Pb3krUdlxRJyJYubpIX+tND/Mx2D2wR7rQqV0N
wdf6I8gupjEWY04grxl476epa7S90h3fSGvQE2GAbjA2GQkCNmcOjB0Ich8XwtS8
/Rm5+QXRzrznIE5ZvY3H0WX8RoQoEoO3TPSX9PYbJd67cZawjFisS12xKtYKDboA
EAu7ZvTYg8ddWAkHnJTmvi4wvqHI+yLCpI3h6C6kpgfzc1cCWn2ryXPAEms04TfX
UY4/9ahSeQ/rxW3nZeqtPw6wtoiQ/GpuvhFSSj+TJy7XJ1BiWDE7x843mUW9VAsF
7Z72y2vpjvfmTZyzs6kX+YlmxcxUfpdDOZdrUKyRSNVnXvB8G0H1FxW/rprHeyV8
IV9M47Ye+5ZB0QWBgd34pw/7+MPIv8RpIDyucE3a1Z5Mv9Yc1gyZ8EyRDho5ULL8
F5jqjXTZaK3Jk7RHqFrSCjOI4WBQZHKc8Q29dS4dqKVUiBNPuyK0b7frYsK22M1e
Cb2zCjDIRX8L2OK2DkN0fhsU0/7sNAaANCNMl8c9gE8AHujsQXxESQdTr4Df1sbF
3a3BwxmD6lA127iw0Jzlq7NqMrUVk4goJfuA7ZtsZsgE/u4BZzS611rKiauG99SJ
mmKrcrtuiahm7a7c9gZ722Drve2+an6BGZvxJQN5qCrmpVOWUeWqhAVKAQmvAC04
ZLCu3urXsWLdZNFJV99v7iLMGK+qrTpa3RdvJ+sC1fdVu66nGtB9Pr0diUD5Ciae
WE/lwsUCQGcQxZ8ehhcE3iiG5shvSg/OlZwcwV9C4NbS3j5U3exUFBiBd23U3RwT
agJv32Dx/z3+8Cs0y6tz+Joiozj58pz+9ZgdSU7AyrYovl/5Y6vb8TRJy6Jcj3qq
ZTcksPf7TPx6PeNWA3pNPAgzx8gwLOPaszZhc/tHoCp1Bcv4OXAAcbxUVq4aj1Vz
pdy1XMJOntFB8fK9WipWCKLKLgpqEnT2oR7Zykv9vWxWX0ZbX/H8XrgiyApq6p7K
Xmo1vn6BvlF4/xWpCfe3A/ZnSpk9pY/Flf4MX1S/mOUtAAZSouIxYsU13xTJL9LY
UQc13Ecu0Or4uXpr9HyYC3Xwghqqi758guq6rN+Yys/geDeBEHBtmcODT1NWMqAI
Prg0+aoK4nnmQvuggcXwktYdj/dP8ayFqR4/ffXmdegctEctUN6Ih3f3dWtHUR31
hokdtlZalCQTl7WzzQoYNtj1xEQzgJCzRZg8FyP+s3boulhFLUF1y31lMg4g4rTi
ab3+vU2wgpzRV9PpC7XN/0Xv1YxNBns4JeNuVqO6wPQl/a+01bxUiqGk8ziNq5PD
p4NuSyH6xbGWhsFKM35lCL5NPAif0KNYzdM7oqNiBWlxT0r8HZ7zhE4eE+JZpJuC
2Vk+2lYOXAjLO3GcIFUd9gowQwS1421rVggS9SXuix/5qUo1T8rTvEMDE+585hNH
lByLv6/i7GKdg8X1x2aoB6wgtOJZozOUUPSCCICWNyP0o/21XkUxZ+CLgWLZr0n5
vkFwiZEFuc+M7dkdfk7g68R7X04GIQpQZfTrRsK+6EZp7BURiLumOZFagmuBPnP6
I2Mqx//S9OvJNuTXV1tQUcdPWpjbj3jtkEbLKdQ4MPdiA/fRy73XSx/OLeHOtSkY
3Wi/wRDIyibTuqrC1Yxm1u46Ga4Pwj4+vOqd36hpO8lF6GAKyrLtPLR68A+x4ycW
lofAMZ5m/peA75JIY4tweBIauoqM+PNuq/s/HmekXEm0QoI+qiF/3TSvy221ceRZ
giw9P0MWOL490V9gULOezkog5hZmKY+QQeSJlW49cLZ0h1UYJ/nk6wO/OLPIHT74
r516YDCyzSnsZ3AQ9SelA/D3gPXDQRNtgguVjHEwJVjUmr2aXwX0Slq0sM++wYT2
1uPpRJtB/Gbxtz9imjNGQG2OxHH+9ez/pjeajFQBGCJgxDW7VtaS6zKZQb50umtu
J6o0EL/Q0whgsL5VxoHWCVnWfI0tPL0I4wWCt3cbzVNajWX8DJ7+R0bFRswDG1td
q6tm/1eGjy6jD4y5L3d/oVGeaK665Xw0T5sZVkLTaTiJQO8depVmC4KqpnOCVhZV
bCwJOIEOsMIeFgHU2KfFHobkoFbbfHZVY+S10bolWgJeQsBdh8RiKaez4/56oMYR
l8A5D0NMkfw8B4pC0dOqo49MvQG9tM1JUWlNtTqU3Eb0kD5gk7qpG0/rUfWnCZYF
gtMmjMaHjkH4WBqsrN/9pcBxOdmLCmKJbts7001M3lgKhVrPRVv8trmlBdyPl6v0
HF7YTbFeA/Mfv7bqckLD8cUMn4PIr9lkEuMQP/EscmsF7pRaUpXX7lK5KQuZp/Ew
HDUuCUnHZIn0Tqw+oCkrw5qGdLAXgFVi4GSepLawQtWwd3uiYWTLFxFg3OeFcIQr
477qobKW2ajIAr7klit7vkP7+clti/8JeT4QtU2jFjZm7ctkl/KiFT1mxWGiIrSZ
LRSutguJZ9QS9yMYJSsOunTmf826KFQzr/Q31/rzaplDhHfyRH5827yKBd5w5IHa
ONQG6UAoOSNvKdmDcdXQd1D6i+7Dye9ER6OZCEBxhVWHc8StY1MfdAnBkLNPZ5j+
GjxBfXxkthA8g6k7SrAZQlT7e5g7qe1s4GZuaFCyKhadBsgE4MNYLHNuGNkrqYoX
m4WV9QPUPCbjjlk5EgWnk7OjxCVvx7CTY/ShfynJY0W/Xjhop230FYx9DS6g+cZN
wCe/UE6eetu7bRcw1QpDKZpFBPtClgErfeyWGLzcmc5JWG3Za+JhtUMh8NoVu7pU
OheNdGdEj5Hoajc2ELuUDIdY2i40tl2xNOvwUg3d24iw7XPM6wAxxFnQpJA/u0NS
IwVvgcVTsNga0BgUG/+LqchMkjQzq9dQNOCHRnDi4Pdal/ZKGHrDK49awm3GgOhm
hthQ25vjp9n6vXySsDEqLMVaKHMs/H451A9YV1ZgWpIblQYdPAtQX3nILD3KnrR0
SpCjdQqfc35bFKqfyZzUvcvGIzFkuypFYoqO31yUKdAOlQoL0r9TRpAgWincE0c4
C7RmsjUqOY+oHr699xwZAd5q6JMMsFOvbxeBvzBLRke773dbYKciF66S5tDkrrwH
cX4ktXhC54BC600FJdcuLgM+iGzi7iEcNW5b8wOeHX83mhrLWjF29eNhri1+CLmp
JOd/HE/W7SGTfLxHpD6g/GBn66dUyv4sueuCVZp0fJOvMa8bEIqZFS+HCS7OCsLT
dcc9gfIGMiHDG/HRjFxE0My8DlpHieKzCYlws1miy2Q9fFwgvsVYPPTbiSH1yo0L
kA5eBZRkjHPd2TgxYiu2IHkIjBvoboij7JSdQYGa99PHDVOrLRJgYEpoLeFUOQ4i
cJo8aeJX+GRe1ZVoC+pLryi3wOIAt0/M/cElxRvr4iiMXdz39KywP4QInk64wSfV
rusKujwMC7mHXBRT7Tw7466+4v7EBbXR8V/ngIk26m+lKpFpNDkkVVDZeG83rzKO
xUs9od8txNlrmEJMA0JNPM1rqnIQrF3/w57b/zT1kg0IlnTlUlRCFyXglmpHOPxZ
/UHyy+YbjAvTyI9vq4bixAVpu2qIS00KEGByYIaGA2P28T724gR39Oyg7ascbQQ0
c7+a9ppM0+447WWWWv+5zFPXhz9n04xSPOzuUZEj2alxuapl8xQh5OzU/84vCxCt
3p58cEscrJFiPIiUHBfDNTXTBbomcubGeh7S0uC0whlnm3CCOf93gITapATlaIJv
EcFBu12i5kRgGd+UvxMlK3XD8BlGiJ4x+cKbMEZ1rIHw9p8zi1Qe8kJ90tFiTB0J
WCkHKOVKwaxa3Y9XzZc+Ix21Na43mo1GoajaVHqCsPPd1EERx+7OwdzglwBQALxW
jv+yvxoQkJyeJmrGc66STuGD110P9QyUEBazNS8gVkbzGjU8Yw871sI9hxHueAAl
qYiLYVn2y5QsVFsnT7P0X27IuGb4GfQjKwTsXceKSgzBi000q4CyflDIbwUZMgBe
G1zaFiXQ+z6CkQrzkJKUw8SmqhWmsVReg2GqPnD91B9phHbEwc2541YjRoJkLaB1
LL6WdcTGpylrS1Dih39mxjHQrZ4NdJBAGbZ7Ie/C6MVAz8yyrdoEfiIEQsE3ujoI
0cosvwrFYS1z/XV67BJWwXvcAjrT4ui8yfZo9GTUGT+WhbxZZC9dAnTR4ent/gRq
7g425BakKGQUIMb5IczR+A7gDXzyt+vrQD4ZB8y+xfXsbfJblJAqlVbFRaxipKSs
gTaknSJQcPLhFfVs+aVIpqGBBUxrBPBGRNOcCGkw6Uc1WZJbpk7KIKoHVJcGew1x
YlG6gALaqOu7jXcXLxg7PJ4Zf0F1Lrz2W3CmVs227UpRoLA8fsHP6Q5D2jK2WCOW
YdlSSiYWf0YdBWJnFjJuTScmflxvx0SAvXiUcgLf5nnggE0uro2LgJrFHkjb67qz
4LCutxhqD/8qGD94orGLxyE+YoMthr7DzOoikQlUW+Pyqo3r7OQFoEvzZw8tv/lM
dSxT/JCQh0bdZCx3SsYNNUHU59S7CeIzc1gSWo4lga4SJ7teVupSL32FP3mZCKLd
ai5VJfuWqzo1u0B2N4kOpc76Q/Z60HPbjA7nOGfal3B0+ChWAZOOndWa9aZxRNBu
wxlOnKo7Ruubal57SuhsnGYiaX5SzQQBXqbP/nj8sryN3fsabcGThW23K598odt9
wYX3meh8boD56hW9x8GSQY/ka92m6fc6yVu0q88YxBXKCS6f5Uhb7LwdRLqMaaPt
+oq1Cg07GZCebwflukHry0B1WNbzJpehivliaWMWfAbPS4apiVV8UzoZGRuw7y2v
naSJlHbT6k+RI5fNco22R9I6WwP0B/U2cbHnLhzQBs4KttFIjX1A3Icrmo4+HHsG
UW6SpNvzWQNeMjQCRIyp8OzvrK9C5NfzVoMjX0BLHTxy2E6dCZsWB4GUao9tSFXR
wwWYWMv5LqxYIVo/ApehkRFEurQLpg0J7dnebVNQWxUG//ExikR18CYCAFXdlCjx
cLDEJ9XSMfnd6vteYCMKruak3vC5aLUznaunX5b1BIdFgyJBOL1Ddf0hRp5Zb7AD
MeY972Y/ZekqJC1+BN0msy35ffuLB8H/Ymi8LQs4bwe7kRo7skB04ZQyCRwUCvJj
+elSpGOgA0JlU4N3cr827xh4KzV4twQx8uVwlcv5d7GA+P87TPDuYUBGtpLWwqEu
aqFUr+bwA88YA4RehxfsuUuLWQR5Is3BcLR6IX320SrYr1TnrN8RDu4eXLVogNef
aIPAa8tj9WzaVOkwVincjGRls4AG/k9rRmzE5XSdzkQuVlHzTty9fU/ysKSt9aQU
AOgh0kUK20F77I8BmsBbQFNwOkeet0qNTIltdpbaZhhW0r2v4F1cwgxO7iNWBsyY
npjCOm0XTXkdCboMCD77pOkRgkNAyGH+o1Ocqgm/ViKahG5PsIsuFmzcNixzI39/
hE3IyVlw/PQ5bsLfy5Wplwnek+jSTM8QyytW4HwITHotJhi1Y9MICeb1t3SmBLeI
7+kmnJtUvKdwbOXQkBGfdS1gCyQ6y4n8L8xdrhzCQW4PiUqUVu8if+S0WDrlF5Rb
sSnT4uMHMGolLjw7lv4mi9KEz1edea5qG9rJhMywXpv4s9ZFzBHDxjWqxgLvMqiW
VVjzWdUe8+PMFctPUydrKEuK0KY2UticFKx5fz4d/SBYQ4LGNd5nXznXLHZXrAGz
jNrhv9mVumrDtpNlkbHC9j1KBenisro4eH6Pb18yGWH6Mg61vSozQIi79sqY8tDg
92rMegLR4YT/qTtz6xWH4ABfEdPHxdDhnW8Xr/SlQF9pWJ+5wkruQuwGVEdN6ZfH
hLsaXYoa0aPknOoBnMInIGXDFcfcRU8rO3vtVY7zG0CGtvXvZhbjeLYwqoAjHWPS
p8KqIDlU2ZNDZWVDRBldbxR0Xjua4qC3/17yzN6Q7cHdKFOwTCKPOsMuha214PP+
ByUUDd+D1Hw398q253cdzGWqE0IvnAD8FTHwA2xfGb8K4AfHMnLi8iBNSamQ4Sg5
vtvZPGTalol3c0LbpzHyv0zgotjXFI9SBP0UFBNSaNlOldz21di51g40qqrOYwfr
buPlAgwSANkiqovyDO5Nw2B9WMdVlCmhBJMQxwhGcVWSzSaCvfP0MFLlFAzwAv9T
Nh7A5Z344yZqC9aegrwmaRP4stzx/iWUwseLG8uwHNbJ2ZqM3qSG2Xbffy352Xz9
bqzz9C/GTwoh3Z9ZDUXnNcsjj9SDZNzN/7EXsa102KiMMCBh5mityrEQfjYmRTJN
oKsafJmrt0Vrfzhx6zlBZg0G3xBiqlFhpILorEdXo+ys270PlU8nDv2ts7QirCHq
sEK+sRQ1QEUMYUQ0xMLq8g0PO/H0OiNvZIaLlUR4z9aNgdTQDmQGTWftZ0j9oNI2
mrBgm72pl75/0qqDeI8JjT3gztiReLyKSR4ll6Xw8ABk3E/wVlGBQCwSWhbQOA4t
G3NKbHpg7B5qr4AQuzk0vRIu3UMubx96fp8k/wMZ4Q55maQ536RPlUwXRTEOqjC6
lIOWgpi1nuPUiyb2WRqKicPqFCVJ7nhoTmc2xzyhwoTwQoOUiZ9Lg33iE6vbbAgy
NEl3B4uXqdRIcVGTHnImEHpryyhlGfZ8o6YbNILSvJaTQ9zKTGOGxQxQxzqRqjRI
TNJD/gL8JRLnvLEykrLtlvV8ieORoswmzL6AkikXj0YaeCcvt2+iTPc6/dcYQieD
yBsZnwC2yXJkynNvfqkWAZg9TBmpxI53BCTx8XDYRG3Z56B7DeT0F70Q81Ofliix
jQcYxBijK+VkCvu9DJLUwpld/l3dBSLllrpFqE6PqRS+271PmqK9DBOzYLoE5F5o
JcShc2ls6QIwOya7weUB36IkCBe8psqBhxE0zP/2xfK9pnpHoiQJJ4QYIGR+6rCF
tOGqOgR3O5bUaTI6TaOkGH1LgSm5xCF1ZRx6NnSLDVDR85Q3S9hAe07CkE7lUGVZ
B2UX1R70vyj4LbuSSawf7O5ZMjUjn0drtwbdnuURHG1y/hlutZkF2RmGJ2U4NJNt
2gi+2pse0Koqh8QN5nsp2acJbWvaLjNP2KtVF6QURzNY7xczIv0oylwddboeuaFJ
KM74nmLypqZHA4y55APFvMttU72O0o5WT7uJgNWPglX5Z2SgZYJOj2XMpIKS3wyh
rdf5iMf+8I6rMobPPsEdGR24iIMkJ17tE/76IJFTw7k/W46+YCubKF6Xm/ZBa4oO
25LyU7UBc0UdyXbuh9fHsS/P5H3Ivc2wFVUGyY6pGetTAtgO/R1A628yZtm+EIsi
cp0Z27zjfe6sv0FnP9IPKfBaZO8l2UW6VaNq5iUjeRFoFRF+wzgNXZT0dNkq9sin
4NcSnJwBKmaehFGqBalhtbvR0jmK7e7gar/HeVuhglsgm8mUtu0jF0bIQOCTQCqh
Cn2xsbI/5nHRYKM/ldimJYdlk6kFwTu/R5lToDUDwtR0B23pOgqOKR3Hf2bfgNbJ
tjM13gm7MYtCBIXoeYZNMftTt3wY6mIYtQ9P/Fs1nG1YfZ1YpHXnE8SaK+UaPLOH
nNqmUgiFrAt2PGU8NZZft9Hetcn/ZzsvaI+gFirm8M+j5FGzkbOyjW59Ekf8hsmi
xnBUCy0lEjiTximGoE+qizKdbr02O/TAYuM/PLq9mEL/ub94FWkyDrcG0qW9DKeT
oHF/wWPdqKvkbn5CFY0T/miw/RqIbF5FZjE3kr/iiHEUA3UNrn2sZkS9Tt6rF6DW
KA+diK6RLf4ZoXZ3mwjame9osLvbjxy4/QqKAJwJjVDeCCxurOs5bNDVvtpa8Qz/
qfODykvAfM+h6KJr26qP9vUKIJqjExvkYl/VlbgmXc+FV2sHRXd2H2dAbg/vsCGz
KD3GrD/Ostf2LuLR3xDLEwpzf2yIngQuc4CjtIzYsDUNcHr/N9hYWfj7kx0EoBGm
xNzaCJ/OlrNAd6xXch1vaZd2swyUN7XJ2gqd/aRVne+LNxI7CEJjVJv93fouCcLq
QEvsax+M4qQ1yy4GvdvwI8tm5m+t/poTepvK0MKtZvspQbCcNqSUWyHZzml3thUP
n8hrG1S9kJpGjalgPygbY9axrs9NQq6T0voMSvwnPdkmeTicX8g8B9Q+yeBX/hBV
bu4J+fXFciCsNOwGJFqt9icI3TOXKbRwJ8EO/XGaSBiFWQOv8d0QIVzTe2uBR2R4
zdJFtguZ+skIQqF4+fnHhlkoJ/26Jmx82P8qnC6HCwyFnSh9dzGIcyiAZEiPWWFv
KgH+FljvZsharCkPt2Ml+yuKl984HHrwMuqdOC7cP6iHF0NKK0Jq4S5k3YolafWZ
fivmRQ64ELt0KzqJe1ajQOfsxOjDvmPcWEz1JpGgwtqI3lCHNslVe09hDXyybQUk
1Ik1St5mMfUi1fH+Rd5a90eM/oNwPJDCQrBlMJ71+8bl4Ew+FYJcXQqyqQu2NAd2
84ds8rJmyfFB+doEuNNhjoaSY+RJ+o79prIl/RV82JpUAbn/YOn9qcsv45WKfMOC
fgwSGiLiUbf/frjV/a1QDmq725bC8W16s9yhz3uQqX7IBjzPtyIZ5K4hTDkibtN9
50cr7DzlBNw2PMtFxAZ/0GewH8OixHUADTZzUhfAtfsuO8t9frXcIdbPsz4dvr4E
6A/oMK7/lc5aETEAMKVYtYcqUrui/ODSQCCVjlfKogHB7OdQFBTrpp1dk8R4qUcg
hFp0no0wFBj6XaZvLnwHcVaNtEHJLZYgD1JXt1OyyQ+L/s3xE8tUECsLcUO2qMdp
sjk1BhnGOA9VIyjD81Xy2awizHaAkho13s0mj7tMTUZ5QXnUrvY9GQQhAlkIl30/
OnXlc9D7+/kwXbfFt656MYGSztPAce4RcoV2TCmasMTi62f9wnjwN2NlcTciM2K0
ji4AvbZEFJn0i51E1T+IGl1mjUbX0PR+4J9tFTSlpl7xEOYKXZz7cZy3f0uZMdHG
RzDGYdgtzsuFO2BOs7xlxOHlJRD9l2I3wUPzxS0/3svba/YoDxPo0rHb6mAgYC22
f6+N4aZr/YcHZeFBjtBK073KIkpGIh2u+1HF2UopQQFkTRWoWZxCN8VPb1fR9IWg
ihcIxmkuvmDPA0cVk5DPPQEOiGkey3nMVIxE7SBGwnj2gJvsR583w09YYfvLueVQ
zHFq7xehp/uKXvOQgAJJpyczKANSdjR6gF2+9Iu/jKW1olbw7d3DVZZ5EAzj4el5
AO1ptlaQ1JIYzAMYUfmWHnkyRLj+zmyoGOFsrg5f7vzhjLkYLUq5KVhHq1aUTjPc
GPcMwNyn1yYhdAl18iNnHJOEkzFODJTzKuDIsjg2qi2R/vTA2hvM8bzwD5lnN7qP
wehrqZ8wNtwAS+nK9aHghG6BIRzybqacp64kA/WH164EM3htWArgfxiAsPRIWsiP
QJqg0HxfVljsQ3TG6VzVQl5XC8rRlXvfrWsto+fv5dt9k+ApxnsqXMT7GkGK1Itp
6whrXVRh59hM05MeFdzKWJPVHlfBQaVPPAbQeewvOhcMS5qRqsx/ayylB7c3q/tS
MnhHL5Vo2Hd2ggUR4k3/AlGba2qc0ZRibx8vfihlFZ2yTzGLa1xgvmQJ0rlOnYM0
ArMEZCqw6vmeGeKins8Pxaw/S4L+rwIwmX1Ebw/yBmhGNiBIYWrRR3sB4lA0Asp5
YUSTvm5qezQxkASi7gfIvijEuEhnwfC1KtTjNQYHlqFdm11K1xY47Zu2CLTVbwcQ
n385e0j3IEcDe4d8ivi8Bh0Teowb5MKCx1YTk9Rt5cwW6+tEFxXG5BWzuUkfNhJq
AmysmCzFfEcWVFfX2X5W54DyKbWNbn9CK1m4+dv/D2TgJwVp2M4zxsiaoHWPQPu3
EkPM9GjmioMPY+ZnNmvSb+bWWXlwoPfuuhPq/ij/h08D8+4jEl4qTwIZQI3VHPtH
1s6b5+VWYjqBrSD/lsyE/kVdU5mfl3ceG0jc/035P/bZ90j4rTL1Or6TlrIjccHR
P90pkD2dLQx/YMWdbUh4fe01JD1SHYHQje7WDOTdJMuFfZUv7YY/sJwjuMczabi/
o9FcuxLuYI+sxv3bOg5xj0RIK7PffMnq2Cw7kRa2Jm6iz18lCWJm8riog37KXFsh
OUp4A30TJ9AeWBlOUABjtGPfAvvXTpxqjlk0SMd5adtsHTVguA2Iv7dd6ZpGYmoT
i8iJNSSGC5FuDCZWXSesVoX4SCA69QYjctcFqgZ9Nvmahh6+wptIKBsAHCBxPKK8
iU5yjEQs7IJYI8I9JL9Sv9vS7x4ZG7IpadoT3rWcxjtmKTJ9UWkHcdLp1ZJMl51W
eA61XCrd+CM7SOz4Rc2NUlKKOtdRCBrvHmXs+kjdyvHwGIvfJrNJrV3hrFbyznNP
dyMdNDSMqwy+iKgHquJ6SvZgunqsMgq39q6FslNIE46NYTtyaqK7KpvtRFRHqkJR
yJnsVfX20cV9g/rcTy39qrss0T8sM1aWBaktvGVAXyEE1V1UnXiEadKect6uxovb
WnTbioV2qIFEFFzj+KoOLS+nhTbd4lt1Knmqg0fAAl/abyHLUSry94eZiEaFZVDe
wBrCH+8z936fYzYPbXwa8mrkJBjhZm22AvMtmtp2Vz+olv8JzgmSZW1k/5C8cHfd
wUvdBWFW7yRb1PJPpukKMocc94uhdP0MwEgVq9O1rVKyvuFZ8Zf0r95uSj8LSMPP
sIif4rCZwjR+vMJnqJ4keVxmi//hhYIpCOw3atw99Zu0EZt9DT7LpDmmuL3hNESx
ShHQfIYdFxu8CQrGRk6Myl8pmtDVoiToG1iTEx2f0GH+s6WSp5Dcd7fZKoqPL5m+
gRJoWuc8RZCHC0+roeMX1sPsoqpzLIbQx/knU3Ih/JVlHoRrBDhEe9QHfs0u2QXK
cv4coPGdp8hZ9RdI0bTCEDO+m2wsN7PJHB4WIy0Hchz5w0/ULmVZrxB/ls8O/TWB
Jx99ggsGpxWgOYoNY8Gzu4VNceEA7M9xLlb0jtSByeJ6u8B0UlBcbr9Y2CprSdhX
6ulqMH7rmyQRyFECL/mza7zOUArgrcYsrM7y6mfZ/SupMLIRxPnAJiW7OjBSYHaG
1B/Za3Iiho6SOdpb3Xpfrte3SOiwF9Yp3WsStmb1+ps5WL4Ws9zwz/oS412aclAE
/ybGfjge1nlHR/Oyi+7IziVIy3gOvzdYiRmFXYneAXSUM2+RhqhGQaOyn4MSlp5x
kJAUunQ4WZeKrWAG389OOG6aRlk4QBkRN1Ll3isZi3N4V7Q4Sld1E2OX++8yY3Gc
baqm6baY2xjKyi/rijJCNiH/GFkbS+7WQBPTtWoyux1uwU/KqlwrHSWtCsQAm/U6
HsqsQjto+NBmTs6RHk7DKFeH4xZR+Dz/T+MwyFQbqsdEMKNhTJJLlBCe3t6WRYva
Xzeyx6soPhzB/44UwkiFYQI4FP6DqIS4sxRVc3vIY9rnfGGtvVNoBpmuNPm2bHEc
ys8UsXR+smVpQnWHbUeNHwAddSUhkvQfyIM78waKq4bweMj7D21beQMEZKlJwEbg
MpHQZ5N8N6hAWK0qucHKQXGaCQtIw4O/WflnSyqvTtEdFlNt9irB7gZemK/2dLKs
69Pw5v11fUOzfcx8UPDlI2Mi6I/RtIbz5NgS0YfklGv+LILv8MDwKlAXdrJffS9j
2wjRbMlYxB4E0eo7SX3bZ3g6e96Yu1HEphTuMjR6TfnNGEIfzdJ3CEd1QzbzB+5K
DsxtsEKUmzD+DCWMPPKx+ywYrNPXj9vbUe8gUyte2pjEOABSVbfriR789OJu24jg
aE/i0x9u9pxH9T1z+HMq8KnMCztWBSGdgDSjHmbJvK7iAmEEoetLTeWKSVEStjgV
/9qNeCxeLBo/zFXAk8l3Q6c6CBhXRs+JnZY6e5XETzNJ1A7HMUBvXr7zZfq6Ku6r
pEcR0nxPJAWAlvgIQHldvq4ulNVBIYUbavLe4Ddn+PpZxar7k6xE7TODtniqSlDg
aPbQuGlkx8bCPYSBrV3EX8uMGOOcuTy4h477CnqCkDatAt70DrWA9uN6+RoGB+F6
q7nOShdX5pGJI/LrkLtspwX/elAdLbTzIs7PFmS/HAENl6OR016sFOgaQ151k2+V
MElY/5tKeiXVGZweR0x06GuH3C6IIr2uGbaEoyFbgcajP/gtkY1/I1+RvpnK3fhm
d1iHwIeavTan5lmi+dIrC0Jjz+r8CpSrVG5Yk2B6+p0m3MUeE5ByzOTDccm1bYMC
7p0ipjq+zX5j5k7B+RCivdamuyUgbIv75whCoMoz3uYvQvRRbTL7T5x7VWHFU2Yx
+oFIEf4V3klA5GVdXk4XQg03odaEwEtwmup9WdMmrrMzGs/T7ZTKhn5AXyUfgQIO
EYcqqSg0D5XuCDH+G/YPCGerzdHT5IYWD1cgCEn2J1b4OLzw44mK2DZmC+qeZC3s
Gkf7Qqj/cekxLwaCGvOTW/q0Qg9I743GuwTFPFtRRf9iezUlw/RFdW5k4w3aqjTH
QmMSLdrcXj7CN/iglVX6HESlpSSbk/64YF8h2oTzjoGiJRzLaG1W6MkCGa+5zNgg
69r2sJ6CrgcdZ3hIxw6AW2xr93JJ2bCOKVJ+s0oO76ueYJSZHoGAdMeqXXPEPPnJ
2X6iIgABbzH9QMr8EkYAjSNx6JHmVIVVgYAt5Mo3BNfl21/2Oso85MlyszJukTJW
9RlM8NBHTaPaT5/n/1vEs29ZfozMkMtM2I2yESQSrbmDD/N2VDZ2tg6GEtbNr2sA
6sr56ODXmQXibcAYSjuu+cLrYMf5ns9RkDfV5naL67A9X38h0fdkCrtHtv8WUWlj
Rj9Xra/w8tT3BENIOD8J+CxOTwQTXuCG0cYGrPOi2GmQoJn7oWrpmQRyjGYGAIMO
I/hXRhb2AwCQaOAO7Fwm0jZ1ctKHctQsE8PlrxEFzuwNhsTulnbAmZPGefOPJWHZ
kybTTJMtu0o6OKMp0MbtxJ7D7enhDugkN0t/qMpMg5C0xKmCWYxG1GKJuj3HGFCL
1WVncBQTxEzfZQRJZ2v5H/zrtZ7+Hr1fQacQbCrirWUL3cH4JV5uYEhkWHe2jjri
6vJ9qg7e3bcENo+uxaynLfGHI4DJjO3d5GMh2lDRFVVupXCzaopnBZK9eVuKJg+c
Usm9I/fCQg7bBHNj8cJvwLOVdMeQy3G0Uh7q3Ts/WB+JWOqWbKnv82uvZwDG+XXR
q8orUcS3BWGUzhm0IHOVlpsrTTsB+msY4/2hJlFVyKVzTjyPYEne4qzoFf44nICq
cXs20qVjItooBKx0oRx8LY7EAajoNWaUL98+PSxD4F9UBhNTCzeW1b8UmwUd56SE
XE0ICuyQHauMed/DUljGKi6yzMzNnWh6J49Y3qZrg0uzbLsJzrYbZDWJ/+mOj+hE
TOUz/G502bBrs5lCRx/jGyZKVvobBYlUKctXkz7u9TakEAnwZHxCpWckRrueatWf
bM9laJoXQVZkAa05ag1v6B49DUHkVyDudfZ+T7bw6sP7vo/S/c0LOA1eqXi9gb1+
vWuamz7sdq63+rJrWLc5PzETwfgxT5sZgtIWnge9mSpKjZkJ+bjrnhRp0raG4txN
cAT0850hrGyU/ytDFSgPm5syEa1GnRwt7u2y1o9aP/rd8CULRSkxOZjC7Av8opNh
G3I2yWNYk7k+wMeipw1lbKxPwRhOiBVa/ycO7BVQLsmAi3cO+/8kT7T25GJYL+ng
B9hV5vAUMdIcLDjci80GB3VHgJO6QoDkm582AeTr2DfIsVas8spSN/Tr8LjbXFLt
KuI1itnjPdCXbj/MF4TN9mYwC20H2D/tCNDnahyCjicaPzMWNFDSOAZF3b1U4eVV
qCukKmzM+c0k3Wlk7z/e/sQA7XUb/dVoPQm5pwKMyOKSkux7NSorr4WeM/5Ax/UH
Jye1iKFOhMeNLalCMNaqhpCFP4b1ucqMpGrzEmwYSFG4bB1+cgHggNuphy7mTUG8
xjz6HzbYvkVxUv7uNVHw7xOlWMhXfwDBgX8ReVFHQcZDTAK1uNuvd7pxiRgdLvlN
fuqvNWkhKetOxirk1cjOutu3QxOHZ+5GVShggWWW9egmWFzgqjWgKsy9D9VJtWL1
sIQ+4vv8KhPTM5YfDp6GiPwx29/QMtt2sP0hB0yji8ozKM3INBJsUxuF1budImvM
F2RQl+Jph3VZUNf/hQ3uLivFRCZRUZypMX8oS9gHoMLnTF0uggsTC96SjYruOLWa
uQ1q1OpaCe2fFqgkd/lg32LJ6BiS0xsdArP/tNC/g/NeiBGUqaEtVY8P3t263dfi
VSP8ysdCDGhCVQLvqmG0GYJj5fTFov+Uy7iTmz9kd31STTlnCu3eEFIjutqHtD0w
wTZZOvuwvTbIVHC7M5zZLxZ9Bh9RpqoO0g9r9e2E+sngqK8dqj8HH2YuowkuTatW
1HrZaDTQd3v1yuSZG28jiUE054vPL57Xz/sRwpd/95sYxAvrPhrc3jcjDFI9y5TE
MgXy/l3zI5KljswJcQ4iq1eXWgL8x0sBghUJL2/0uXfYDYshUItq1TvsP/6R0NrT
uxNOhbN72KGFIMvTF6O5f3PJgRbXeCOg0TWO+izIonj9ENn9Y3eVLg+GX2/ZsiPQ
0AA5ZniGf6vqKaiBFqhBaWO7Z7ea45dFnRua9PxGZuprGAm6Yirt7FsEtq1rCUpi
shV7/zWQk/VbXI8XP9+t210BMTV2pzOID/ytEnQcnz0Hd0jyKnFVatG8NhunXDFe
jjoZXKnN5Q5qqlfppSkLIJxP8KNeT9TXeMo2TTT1Kuc7G7IKnmavno8n9+sz4ker
UQQnnkgwK88gWKolpGSuzJq//k0oakmPQgr/wb+lvgUvwwmUokUq3wG2pQqey3xz
Xmee9t/Wv+74fsJwjj7TPMoBMI7b/Vd2tdHjzNPO/XjuxkrV+gMib7Vun5+BWxKY
O7t2olvr2oCsHVfh2ezrg4v7xD5jQNXWDq/eDd5FScdcEosuB08pZzHeVq+7+aWA
2Qtz+jmqErrbWj3AWl0f83F08Yv5AqKqNo0RvfXSMEeBy/ZntSdOHlnn3BYSeRUE
6uVZvMZN9sCaXe01K+FZGSrklFgSTEnCK0YUo79/qhgFTLWq1b0l2QHtXh2ThR10
6+hrWbMZsfdrHsj1jZz83TwcJ4m443c0n5aFOdi5uqRjYq18YifvxXNFwxRqNJZi
doA+8cffTatsaJRHYE12QQJBMkaLnGf7g5Qhf1LyNiSnbMrgpvqDlxbHdYbTzJvF
nSevPD8ZnjIweZwv9hw2d3PpofEGd5qUNyDjQXSHXowT6k59Nt+/SFsYuJkmAGY2
gqKLOjZxHtV0kAvR/ikEKbP3ofCyysC/aFEEExPiVZMS5MfjKcnKMiihpMtjC1KS
HRPhkjeNe3eRS8hDwDpZ9IKVgpe0Jg5DYEAptF8XTmrxoGvJ8v3KhnX7t2UZo2JX
XVHp8bks/QNYHBjhpv6aTLP9fMFgEOHiKTh5SEf3J8AvW2PzGp2O/VCxWac52slc
zFJsDOfQR9JWnUUwSgsgqXvvhTi9p4/w+yvitgP0nO1clurJ3UCFVg9yrp8TRViw
23ooE4nMgYW3IMI2pR25XjjR2XUJcXniEmOGu19D2Qo/poCoMET69RTqCJF6yRCS
0JDWC5mCHBK84972jsFL4w7KHuXnoLZT2KzL9Heh63ux/81lOcbMC4DIWRQ9ELSI
O1sszz/0Uf93QTp79j0dhTEFYNSTEAHYdy9TWC/awM9oUCgj47WAqj0wfwjSujL1
dU+Rp0FaB5JJm4EPYdC72Ti3B8bKFVWV+iY5bz+YeZYOfOf2IpeEX17VqKIJXoV8
Xoe4StSbuHTewi/Z5THUCv7wZu+3HuBd0C+56e3WNed/idPhu0k0Z7pr3UULnFAP
/ThJRdN/b3OwYE5Ua+ZQrXA3pWT/1FLh4PZaDMFtlLl1h4Inp+JV4ZvXYOpb+ToT
wiX5jKtSpIOyF5P8Btwv0nry2qS8vwUYBk2C2NpHp+LodGlY5TCsVkJUEASbPQql
XqIbaMMsTJCBD5ZwGYw8CdNpcbc/PHFRL37wzpXuKFilSmJnP4QE+4ZA2c0Slhbt
Js0jMMldkcpuu00NyPpRZcg8zXYWxPVidmu6AGE/8SdxYIc9Gr8R0uWpe4BlEjof
o3GnWzUj2IaQVoGYsIDSL8AcMChfIzffDyWgEzWN2VbRhpC8ko9Idq+rSDNhfBkn
B91ynx4Gu3YfdS0zCe4xf+6oPx7+Stpp+O8itZru0M2fMtPChniBv8FvRoje4CQo
+xDIX1w/3JnW9JSIUYB5VFGsKRUc0+mkb707xUvjYzmQaap+U6Zb1tyNcOGYFUip
EyEBmpSR4SdDCg0V6VY+g6vHObR6KUiP3k5sxxOajS0zu+1rHL1JWJL4litfYGdm
7zjWkYsIzgCo0lmVryfyDsrDOhooB17fNCvgswXLcIlul8/dyjbeAxLsCbegb6l/
ViwYxrCYiGZuBHu9IA3rdZtHWJAhbaCtdgn1iKss9EQi/qCQjmym165ehzgSDj+b
y0KyFMg9EC8kGA6R55BCA1B5oO6dEC/d2txRUQOkAKy0LEuntJurJWG7afEX/6O5
k+cJuZq71AbzBfVp1X6DCesMeETv4oSCH1rdxarSRYmuHNRaIQNZghzJIbRamuks
1Z5yCDfBsbMG8X6Z7qEJ4h7T2tbSBOxUilyqrKx7FKU+QRj8ZShutfevZH2i6/4Y
myfkJJDtAXYm4xDFkGKPhJADReIWac4JGQu5jbdhmZYjlKxmgvXyLniqqWh+IJF2
WXRcsnd6Fl+U5C1HJ40xourla29x4sCQGnt3lulH+/+tmpdoz8MhEFr9CW8raWo3
10E4iiV1vWC3l26zJKfV2uH2FFgWBbfnRphBolYy0U+40mSuAn0ES/fhssLbRlAm
0ChS4WOiPiTDm6ymP7K7GeSFM0Gf4i2kUvneWbrFQ96OGqDLp9c4E1KSzaSGLB19
vk+kPFIVP7lNHqbH51trk6Fp7fOPj7xDcDAm728WX0BZ2dYq0+cp0q3y1JANkN+C
WEtEbTK/V8MI4tEZmkxBOQhoY8VqXVUZnjgPPgKfkUfv9TZS2DZTKyOyu5ovml4k
36g12TQbN7rTxQzJzGERlLF9koK4f5J05cQUpqMS40JFzFQhwIax+cYjAb09ptoM
40Sy/ILsoGcuVnFGanOGp5DhDTKKXg22esjJUnrqhps3OSfbO+2XtZF6HgOGOt2e
DDA/1lekLL2d8L+F5w/PUir2umeUGbhe11+BWFT+/fC5+jZ6226VKF/HZKQQR1kk
Hf/KxQcD1puhhkwi8svLen+YxAlnM16INQOJeHdepQT7DwHrkVk4m2WfEBV5kWUf
9H17lwky8PfTpNeGSBGRWmNvp0Zu310McUBOtE7m+7HTBpBT+k8V+vkUOM0FGNWd
330yN1emh3vW2FTWQByfAFTvLm2trIUC+x4pcvDBRfqHg1oolqxkFpG++39kh7Sz
GxeY9xviTDrinXeTaOpQdY0iST9oyipdU4KI6KnitzJ8TyNGBiJpMnTTsq5jsetO
q9iLdiPNSxMf9yBERsm7AIDlhhzezeAd+ib0sxRPR2wXaZWiphIdVtgdCilvxI70
/uuFFBXrF5yfzi4ClzLDJnp691UOiAM8ls7tl91c3Gi32wjSfojetot0Bd+//h5v
ZSvLEekS4Dk1oOpG7tGDpzG09pUEhiEsBgCDohwIU1rpUAQTXZw3MIoOa726H843
bFennKlXn6tG4HwCGGmG/sR8aW+mrCJnb9W7aUgxtku4Qt1z+bJLR990amNUnAQG
3baF06/c4m/rw8k05h9b1EEHoEW2hAqmzvuQkNFP+OoT/UIU1+gVS3NY/Y6YvKfq
4opnvxdb1mr94bJwVgJhbG6t00xf2EMYg9DYaNgxFSSrqQclGKjznPzHn+/hp9qP
0dQ0ppiK2EqrxLhorkLB6VG5jlCh4rQ6HiBNeg6wQKVRtsYQ1ihpgVlc26cdjP0x
ooj//qRiThGwadzFp/F3OrDeIwsa7hAKYSVD560cDyiqfWscYzUcwiM2l+w3kW4P
d93o8Vtg13IvXg77/V61sYYrlUc1Gz+nS6LJw7YCbCEOra16VN4LyRqy45Hz7xGQ
+Cbt220+RwBlhOubzVMNry0Ekuw2v4RZSdvBz4I3ZyM0FKzvFI4SpYC0jZL2XfD4
1fF875TwW5RYjb48x3+CvpBdlGDoCZV+6QMzRZctPdtqYJ72eDzooeSW972c4fpf
1ndsOtdK2EiBZuSTD/L3gKuOXdivxMmOdCHkfaK09p1u9oBlsQAQU0uFep0SOa6I
qStd6Wl+tXbNfvJ0N5oQSc1BY++mDcQ080iSMe8gRfsA145F/C7jLd74MuKP/cBN
ivEZ7wUiZrGYC/wqBjPT1UZkek2hdquGK+xFXr22THF38VCr2MWJqaBS+hY+m54E
0lfX8EECJTobq7ULbp/2P9GJ4+B5d3nf+bnGnor63jazW+p76ytu+s6VW9+ftdo1
nZHFOjoX/spWGUp0Cyw5MUPWYt4qoNXmS379LjJCRPY1FmoeSwpGnd7mnvAstvpB
0ONyKCBK5u61TiRREWqFI1vu+gKQqNfqDelb1MgnZeSKL6xjmIFq2mzIvw1RLq60
CRa7CDFnLpFJWPBYu2mp/Qo0PawAExG7NLiqHQseEUmoA6OL5gbVix0QKaJaE5Z0
SMjf/+sxadqOWSvzWS4QsxK9/3sGGiPOjGKEDDI0G4acNeIEDlWU4buH07GZgPnC
VMDYjsiZ0hvTSSreiJDNSWVxkwoeuJ80r7BM5TCU/KJKNmHUIM497xJXs9tuijBD
JQODBDAIqqESOPOOhmbQWw+8lNUrHeZqFIlhhdNJEuR5ZZmnzyLth/IDcHNrT7US
ELFgsRrwVXvKx9yfioub2fXI2RdJVYSUPrjT3MplSzrcv/Ix/7Ni0KqL3P7oUhZX
oqPGwQAs1+PpPAlH916XWtn/ar1DKfh1aUUypou8oRopHCKDiCiO7Yvi+3EhdH4v
aABxTJf7Qkbq+nSS4hB96/bX8ZwDEJR0lbBLEhwEqqPfbRHB90pUjpodLV+Mr79w
H4lk+mN+ZPclGoMQHCBxgQlz4PceNERv+L9KBqQ2Da8WnPNlQzYw7IRSkWp+XJaO
yqzsTaYw7wewk/amyloUYpDCGsmATAWGzvVWRMezOXrjxMrJDDL7CBiCKduGYbXg
jBdhjvlAZhmnJdpxES0sgIqWZ758k+YDMB1ZxoyGBhoeYUa7F1bj8qz+RXJhPbex
tE0LAW3gmXncLfQW9yPagbTV/GiLst5lbaIctsXITKCaWM1PxTvXJF3oTeKqTnKR
/4XVH8fVwhbTRHoSxM2/Uil5wHm3bEomClAL8Meyh6LfHkopdGm9YFzfKotQc068
Oc/7/0uio854qGXA9GORccwq7Xd/Ao3Ytw4pkzf6RmeAVwA4iQ4rokW9J5HmXdVP
pu8SI0DzRN73oztjtd1wWP+C9cJFljJomlO5WKbxa2v0oYe5SHv+BdZxmYROVFGX
hUQ/RlJnEqCYgzxcRSWpqv0zDRx5p7I9Y4z0aR68jBY2OUapEA0EZn5QUGMDBZK3
ze5dj1M+sKTag43NHF869fYAMTNwts6/9qCTCeRA+2Onbk+mS63DmglZuvUAD447
Kb3Y5q2qbDu+ZQSTOGNad8qDaHebEXCuxKV2oKe5//8IyakW9RqNwOHMppaMpFVo
JD5O8Z8PMbBtQaG2b7z8Ne0q92QN/RQ70ofiwwEpD+Em6xoZA/kANKl3wmI0KEi8
9bTx3l64R8N60MSG6bIVduRJQL+DZCwSBnazilp3pCzBiBDhgjFYOUq4IVHs7UM2
MaVwLx2oVFLrs8hShY8Bc/Fl4PVQApY2jJtXptZLEB67N3G7aJSjPoHvSRs1jWKg
avgrtuS7tTHyBGq1pWsH+piqJ/InAeSXUcaiw480JjUZNe8LhXUkSVE0bqazf7JS
gWT/ZwYGTO02NG25WiqYa3wDzintYbfmXkT9y3pJbBrntClD936li2i+jrVAzkT7
ldUv4A+DQ5u9FNWEYSR/0hQaQZGszQLfHe5xHkzbR39/fv7tFlJroAXpmgEF5Fyc
WbEUeC5AbWNOyThbK5ILc+MTNM8c5MOQw+M4Id4huG6jwGo8fyuzuOf7IU593/6J
42QwIYEldcqUeI4xyfqnS5H6N9il5hJFXLypfiQ/ljiDuyGYnkFi/bZjgOyqpzqo
bIfacLMuFxReNIpnt1BelcifKpujYicr1Krv0h/aWvuV7sjNz9sQ4JHm2Hf4eT7q
5tr7E+1NYl1+kKR1kkktCs8xMiq5vWqU6Hfmd2cp4S3wEMhAIMO8v9/QP1S5N7Zq
ssfj3j24wwNuSVKRaw6WeX8XFxvEk21UHVe6GUzfvbM0VkeIJwgWsOxCGDYQt4Ms
DFv2bNHnHliskqq0m9upinPojJ0TXH32kskOziaCsbhZtBjbqMdg1NZclrbG68Yw
2Y29CYZ1deLZ68xjRF7fyHRi6v4j09HOnPmdKlIUw7L5gUyFCadD2W69PyyybQB/
ECe/g+3pwJ5qeJFzS0CujoOSxmgRorHEYsUGxq3LRfX2wo/9TNgX45m8N9aVL/RM
SpoTRYrB9wNSb0VPfJ7CJ+zj+/+W1fZJaXJlSQhhUpZPRRn2FPB5xKKNYsx0WTVC
owNXHBzk4bRnlROOSP/1EHxKQWL1D+zOsp3VafqtaDumKuVz4zAaPqqkSRToda+4
DP5nF1fwawSebiqtGT78SlxAPhmRhAVrQZdhD/Ewj57HOY58OEOLq749M0e270WL
wwmFxMSC6OvWx9Qtoty3PQPCeyVIZNpetSsaFoomOJ7nNYUKgEvx2whJjJVMASbu
HafsIt9ppr23LzLBdHSQ93Q9W4fgmQzgn+VU7ejyqfS1QI+5dhLLShSYZsfrTrW3
OMDRXNLr7YkSIRpXVSeRbhI5dHINF+VsgEbVmvRYsAUZ6CFIiCgjWyi3++BUzpOQ
W5V1qtHYWjo22uGbQx9KRI4+DiPpXuhBWvcNfE3vUa4ZjgCUvbGwpy2Pm9LG6kJc
wdluJrfRC2aVfuY1A/fJiZ89ypfcugjFlhk5+RMl27hhvR6FwFWy0QnBO3uRzu/A
wY9zvjpbCc9gpS/kzWbzzTEX0E36Q3qdzLv/V41X+bzJmwVdPC6ZrRWQetf6dVfQ
u+w5g+3TkUS8Arhp1ZxMag06Lb7ymuLt5AqdQJGdbjVwT6uyuG9AsQEZOWVKqAza
q+2uu7Ou8Aoq6fr8iJ1L7LnCwe/9R+mUE+v4BczGRb0sku/3w/N2s93kaIrpDFSf
7hc3GuGZ2SGn/FUPHMLuecNN/Q0e0wJlxWCC5+HM4j9FApeed2XTdapIYE9fM/Gx
ZfcBGFAA+vi7hXpREZVfSJWVMtFwB6K3QtmZNtQTOo2Qqv0HHbT3aaoFLLBWOdhM
7/cjLgzatLZM3gzWUZpEzLDIXJEOo/OiGs2UE+XCzdi4iWPVeCbibqq8H00SktGR
EK4H0DFL4a+PSwbjXr4CQHi7RRCOnf6TcC4IvK23/G5iNNg5wuoVBi1c7InAuBRI
PDtokoHgYbMzfEs9oHRiLziLdZxLFXDvOKCXi7U4alkrMDKJ3RRrqYWiYdGWmxuJ
glOYKqW/LVVM1wYLx3tMgyM8B4kJ5J2BAVltLFMQK3KApEK7e1SfGjZ3HBJT2Tug
ZzD/E3Ii8koG05MIget8Zgltp1W/rLPYEM+HFDh1X5zvioj1IW594xevDuWxzzQ9
NxJvf9sKuDkVx/n1T5/rnDum7FxaX/D4qR/IUChyqZtXTvQwVt6bfBiMn7wvADQI
ZFk/c7SwGA6zNeCZqUifbIUzPIt3WM2bQNh96mMi0Vl29BrARvDuqXCRiagJr2PR
TT1xd41l3gyJawg+uR1QUVDDeJPkz5TcJdNSUiY07+kSOAfxlteXHhl1LURIQvRp
rEzV+iz4khm9ylXN2FTdStw4h19+063jqQ3bQXDlS0PwqI5MYzeU81U8o68yRcbE
iWg2hhOKjf0cb4AT3Z9Srb+MtU7MaxYOn1KUXRsPHB6c+EXIi2awDexlaGTasyid
PfKS0tVB5kPmPbxybLp3Pdouo6ZEilfv4wBceMyZPhlsPdr1C2pWNOHuGY32O8mg
fTCJt9UYYW+m9jJs3H9ITGQZRviz/JQvpMniVZ8VCCPNn9KsU3TYYfh7CIaed2ev
hTZDlVd5gqkToeUfbIt1nmXKapkWNvLpYiy5oDAWjo4yWqo1wuDjHsjVFA7CrN2S
qbuTghwbO2pzwrVwqkmdDInFDATVL8binhrCHoXlAQycZuSpNrDzYOi4UJd16V5S
S8RmkgtR5bSyWyrWGroY4woYT5ROO9Y0QA91mXqE1520DgzQk2JUGqerjVe8gJIo
9zW+uuiXZFTxA+m0bUepjI4R3d00PI/25aATBNu/0XzXaMUoaC9bmCNImtI+StWN
xZ+Qfbn7gP4yWrW33hi+6bPCMcNXQeiyPk8zq8FCUcGyY2+YmIeWFjH8uiQFBAQg
Q257J5iv7ICtIuh/ov11OE2J2pK5Xq6RyJBNuy3RugOeXY3/7qrFivVveq7Bl0CS
T33dMwDdtWuHNADpAjUBAVT1Zr4CiBQBaenL8927zoPVUo2J8cePTkJJisUoNe8F
A4yeZpcwAd2KT8AdvtEgOC/4IEt85fg4fZ4hrMKXmVMgJZIWg7Cn7yzoXiM6mt6i
WTDU9ZePWrMpDYI/O4BpTujazAOJIz/j4DjgmU+Wz3CqkZvkQ3lShbhL54HNb1Ny
phXP9XPjtHUbiS3/t2DqdWWBzoGytsTA1ytY729hwB95bklOMbj0bjhjvBpi1eOV
bd0VFZeThL3bo7SE/gdZ7peZZISEddUg4qZeUklKIDcXt8g0DQLcTES/fW9Cgdmg
UCcxT5rwqYLl5zqT5MOuJTUlt6WTFiQBIvzcVJhSS6jEb21VWx8jTHxR+682nfYw
sqc5wjfkjO7R3FY4xvrfxosAy2x82LyzHdORl+ktNnqfIXpN0o2Id2kMzygXSl0l
EVB5g/nQA198KD1fkci3NPKGn06K4oU9slBMvLYU0LA9Tb43DF50EiJSc3JC+P1m
WdL10e7Ey0zhOn7L+4kHnhbiQyw/VRQMKbCiqH+i+K6VMTXD+QTARaT8UDZLOc09
LeoULnuNo/NwYrmNf+pmFYyKYGbx6RkwUF+7ugFx8wIujT9pq7JdYy6EXYn2ReY/
ljCG49NqHApKA93vwdMs4cEukB2/35L5cdMYHkvCmRMUYRJydu6NV476YBLFP9au
hdKRLA3YDq6WfoTUei1IF2V/96ihcmrj//pU/FTRD/6JD+T0K5rHkFWt94uIWgyo
iFNFDB/Fi+5Atl5pDG/rnZ17WorRDEA9i6Auh8vzkNDhQqek503kmX9kS9xTf3A6
vGgXRefCtly6HiDdz6OroKCDu8efNWtMr7sso6KJxqMoxG1NrW3pOItS4i9TUTQm
72zMRN5+nBEhMN4eH+EXYJbmDjYuaDwmoGKVVgOpo0FQ2SFF8Eo7yTi7e4L/bSt4
olHGyIs1SBjzSblS9LiLMNoq4NSdknSX6SN426R0ec+P6xLj3FFCBUNj9h2GhoBB
GIgnCf+ovs2tq5A771bzQWVZrxYH9gWNMYdgAdF5+S7rDkgLpsk9sfwp7WzkrYqO
ABS9wL716XIgOYWNe/iyvyybLo+xjg5TvSlKyvD6J/0XOIW+GJcJLboev7UJN+bg
r33oSMrfilqXlsdgW8HPm6ZGK4C5/7XaH5WS+rKwOQvUeKexKFeAvaThR3NJSO2F
t5AtshfdXvVn7C6de0P4FrHmW5k7d3wIQKl4wp3zWlkaXvSTy34Ugd8WMbq4ibpm
aW0o3mffAyas8XvfMkEsV2aHrHMWWFxzMac/GOjnraXwgwqF044w4FkNmtcx3FM8
TVlkZ2bF9jF5xumG2SiyVE4E3GvtHgxd4Y1qGJvayomp98Z/9a4pmec1+LWHR6hf
QVvWiRoTFuDX1ajPm8Fh9BGXDqxCGylItMvH6YpQ+X5VBK5hEGH2M+9/LMH9x1/b
d6nQQgDL06vE+lxRSR7vUZSgrykMfWVpOoLJWCQ2Xenfvy0/esoVcVqIl+SsTs2Q
o5fb3JCsCvOQywa4eC2BG8m90J/p09UyAsrmH770BjGzaJlbFOcusqk3hpr17uDV
YQiGPaAmp1eNNrFxbS21XCoWZgD9m8EiYu7Dj7nEecvgVv0lYd8nNa1Gth1OO2Hd
aHT87iAhOb5/pblLVeoCp5eyml2NmyKus+aqkRjfhd6WCQHf4xAdU2bvUOcTPVxS
w+JMxImAym6Oq6gUoCY1IWaEQBixO5AFAgd+ST/+7c4BR6tASMhgj4CTX7OrHImG
ypmejKXdldH1o2jqexeJdYXCPtpAkhHkgkfPl1GIT8tHmZkyH12s+fEUridXWj+w
nkI3IpHK8bQPxsENBYSHZuTE2EvlUKf/rztpQVYO76ggMskwrc/MzLchIla+mSTG
kScjrJcaX6P5UxfD9/VpBcI8QLn99zE5yQMOvdtf6f3ujzveIPkjUvSj6L09hvqf
Y2ByZ3ByRh6+0/zcttchbw4r8uypF/D2IQMB332l9YaOfMB9Y3y67fdzgUIGZgEf
d6pKginQMhK6SlQdSjl1P7OfvzAncJoao2jaGSZqlqYBKacgL8njEtebfvEE1cOS
+PLTJwgLSsYX0vZcQkwMilNfxH+XiKrdURcXAtE++ROboo0IvJLnq6LdvGq+6WCP
npVvpJf4ioubIPWWofmrR1q1BunD7ycaeQEtJGGV2N7EzvT6C7vo99SxF0PctCoR
T+qreA19i7bEBTyb00XWlLD4/QIu/E8qhU13BciL53+e8PCFTIyLySOAkvUAodKY
LogJ4Zo27+Y+tvkdI6kqU/JBp6kRMXBzvnC9WqCN72h2i5cXuuPvfQmLFGF2GlZw
rtdT6uePJLnu5pOq6NcBJx0/fw6HWw/SVSMzvbqpkUmNWIt3aPKQuUs6gOFCX2RV
GgEfcFWjgqFvDa5RsR4nNzkf1vG77CukC3xPqwetBqr5Dvrt1pr+SxWp6P4lpkQt
jaaEo9r7iCY74EOWMvFytphgc1VHVn1gKnJeUCfVNwSkTGcQoC1HZ95OhFfB/qeL
nUxHiS/6gGft+Ll67quaWSeilkEzeKLclfWUPSfZSq1lrMdNb2Qvwjip5z/JjLHR
jeJKWRJjW1B2uDdIw9+sPXkBanVp2Fk/QlJDawrT9Zs2FrPEGqMzOLWz0wn5bZTH
sLoyKbj3jf45V0nhoXwiBxIZkB4cCW4V9Yk0W2hY61c2P8cdzD7LeYQ8js/FEsD4
yfycQqU/BrwlXl1KlIrodSdGC4nQ/hT6pS1VcLeuG9G/2tvqEc+ZMaCmufQy8Id+
CEek7Hl+whhuH1L61xkc4SgnX7YHaaF9iAW2g0KfCOnmV9e2UayJ0uIbIhOch+P6
ozz1+y5fdWEOj2xAo2DXFoH0tm7HCihX+JgIlYnObigQ7g8RNL/T2y0pKpKsmUJC
0CX7AXESJZO47f54qqnnkbzAvZoVkN3jve+7eCJR2092Dy27YojuwllbJwwOAGn2
UGLnpdJ3eT0PdNL5UyB1ZdewlIEv1FFqnGrOQiD9CZdYxls2WtNMsPwDuqJxN8K0
QDwpvaNB4DvfOBmErYJE4aV1/Ewqw6pptTAbe0Xhid+Sd2NSKEN7YVk3XqQEgjRP
s/jeYfv+1Q8t7yPAeHovhiLOjFSOH3Vx7ETHdwsCT8wUSL6REMJkNFEzGw7SlqIf
kI+U8GTYOBJ/sNKXkHrspy18Uz5fPl/hMAQZx9OAXduunhGt6aL2CF0mCfaKYk/D
oeKleCDkDYiIch7olDC4aljYUuvx7sly57onPbhT/Sb1AEdgzP6L+Fq33l9uxDpn
ZG2qt3g9/WmkJ81LvoYBgH4Le8bkWu9gG+Q7usFsYIdwDVz3zM++TIcRZgSCcaGl
dl+nUZvBSOOnILgVV2HWsGgXcx4ct0ane5wOH+O31rDP9iaCwOSi//o2K8nXrq7l
LKjxPExEmCVUZ0FzLQo7BAXysReK7VhDcV07LLlm7mOunXIP5rUv98+BXK4G6T7E
CgGp+ul9fWg2dh01/MRmS62Os2QGLF5CN2VemNthocw5wSlhx+aExQEq4GtyrO+N
ccVhJgjecYjHixmonRnyZiRkW3dO2nyTwq09FGJFf0PmABTAyGNpI3qopE8Xl1Me
fsbUHkvQPDT8vErV0GUwMgWmJo36MM6cYJs+oJz4oYYo/+jw3ZsAY5p9+fM3Gf8s
o9MApA2Yn/RDhCC+S0m7Iru7kPDTBLAViQ/yrseenqPjCj4HpPKuj272toJ+sCLC
dXjI9mAZCSV/VfD6XvZIOHTg0FY9ZXVOCJTeR45EJwuyMlknpjcPZ1c4dhMWBbl3
QJ+WD0IekmSq3pxEL1ZoN+pYBcXtWQN6SSFRD4XMTuFzWKGoQpHtTEd3ET/Yrram
O7EFHDhIiamOkXo5ujKZEuPhtbLBN8Y40X2CN4XGqPW4YEgL9mRbu3lr2OvyGhyA
t/p2QpQ1kpptZOdAEkFeYMfRxXfOs/s9o6mzliqOvszDwPApYGbbCxMBffhWwLGv
Oqq5NFsm/uQrDhpriH1IZogi4zopDJZNKLRjL9PkVBV0L9QYonRk+9MtbWHeOtXf
4TNsMKt1g4jCCKoH0bvVY/7dK2THrAG5wh8ya7SKWC7tfuQ4x/3W4HxtE2QeRDok
2izhyrI5Ev/r3cJFJKsTDg5i7pD+dSN2BIfntVGN8mX9JrUAL4gRWUre53aMU1z5
oVeaEy9sEDzgjlKs/Iu7ZwOaK4bnT6MZQE3Hjo7xUqCCwZbPN5lBwZ5XD9Aq/o9x
LvEuuiwHTkUjy8ZzL0y1Yz00OCD8pRxT+KfUPxAr/zC+VngSqQxPl83/zrfeUKG5
Lw8L/r6mCdbuTLR+akYBrMR+I4T/fPTscOk9RKXZmP3wNRCpvNOrE4dt4nNbtQPI
+kVLl7LLthS24CKmyk3/dIKNjPXdfGF7Tqz39OQ4G/CcyU1qqxe4b9CSAPcmVW+6
u7RCDr4LxIIZTmmbGpB2YsVApHSbQgv7Mt3QQmfqsufUrkiRwW2bbmP+D88imxXJ
J0vKvvbPh+sFiUI4NSo5iMaN5M1jUEQOeIG16YuzfgRtMYa5DEXAJnk5m+IxbMw0
6yEY25oBgwJE6wWUX8DA/PJAgTtGCUoohs9jR8LrOdc3mdLVeWMPAwL9EoD3H5qD
6Z05IFhwte/cJ01HlSnXgZLJ0OaGuxFyaWkD29GxCSclBAgG3gnsjaJ4JfAzuwV7
b9u/1tiEdjAzaR2C0Jg9AuTukkor5d8HDGtQWOydwPzj/YhycF3VJxqByhTJLLZi
Olx72Zv4+URE1qPm3sGfaHFAK5Ug83uLKVHwsVfLyaRLn0waIedpEUiO+lMIvouc
z6lOmJTuut0liD80lD75e0/243nT5xFzvO/w7/4PddSuRuxxuRFnxYzs7QGP2poq
BvF8x9/DVnIRZqt/KBNHjE8+8vNpKOfuui4N6q7rKuFkJq6JAYs5bpfN8504T2mU
2qFaMz3HpF3HWDFCr5aNRFFBrQutWZcW1gYX035uaBFL7dkU9nz5YK5L8kAKN3iK
+eq7V2NMSWSOAXzRnee5r0Lsf7pjIayljwizVL4atzRWAe2h4gF/TLFAXDprti5G
yTAsz8gcwq49XABdSR1qnZAb1s52q/t19fiytePTJVWBJAa9fUzh1yXsMQFVBeD8
dB9Kmjiiehs3qHGuW1TSoEzrhdAtKE12CvKJA0YjawW2uyva9FuA0UdBn3cAzR8c
/uQRvrv6zmvSoAHtnMf/3x9uf+yZqPaocQyVJU2RWMfI1sEQJOeQhi0HTdG1lmNu
+ek2FaJ3NHI3PfbOYmER/GXbubiFYR0835EgbbKi0tJV8ab/CWCDx8woAGkeDlt9
ydJdHYNzTt1c3Sa4YU6MOLh1pLXsA0wYXvIBPD2fpnbu60WWY3pOGgHuLBx69/QF
F+XPOjrazOwE/NSkO9SJsrQqETxt+YULaXjQU5mRCbirwtCISTTk2uNpdhVkXsk8
d/KBddD7EcGoDbpxohCG7Yyd8XQdZU/+8YcvVVDp0YpOwe3Zbmo7c9WpTtoWs2xp
ZDDZ483kwRQvjcs/2lfqzVNHnp+HKfCmFU8xEt8sLoGDFojCvSoCRE4avEWEjxhB
RV8BsQuaETCThFWYFZO9cP9AGbQSUbwTkBJNFecCs12LWDGGxuUm0NFuP4/LwmJs
QFjfhPLfsfcg1rVy7fxdAYSFQAqdGFUN6BUyFNkgcyy5peKO4fqVjjmzaevG0caz
v+gVYEu7u4KSVJj6fbh4DoscfnVSqqN3wTJix2NY0kwfzGbDDHfhehYPThLKTeU6
x0zFzHDYFpFW7tPpalH64wdE/W2bd8sWFDJuD+1cRILcO9Go9ZNZPwum+MrCoWtt
L7oEsOFFhSOQADpm3xbykpxDUsl/hMdvsOvs0bwiZS+ASLca14DgrJvOqh3d5KwB
wZU0FeBeplMH66ZDBHgJjjfX6G/aMd97O0xxX9Yu5rR0Jh8wewG+m4G3+0DkLdCR
Nq3yhKct4XAuc9bzA4RR1eBc3/F7ykNONC+zITdW1Ymm3kcgWxRZOyxzj0KEikq0
Z+UoFQahy3FFGReL/mjPqROuv6VEXX+wCAL9SUoP6W1OE13h+gvq1ky7OeYLWkX0
i//jI+XGKE4mmba8h+xBpGFbKq+ZF72yUFq3IsNUhA0eq+eDbF54UpkzdQ4Fm41Z
2vrzxfO5uZDN6IYs65MC5PqaTvN0iP+IuAsPOgc0GNbhTK/W6sfIZEQkb9sH7Pq+
yrB/czyWivsuFEewyAo2JL3GZ6pSuABy79VbRhl/YxLS2LQgKUjNLQ2mjNnVlP3q
qTgkV+C6T/SLljqEzEFwQwS0JPFs1y9rZUazOzebjrevUY0DkLsS3oLn5/2Yv48T
BC310oNzWdKC4m3olBxIzz59G7Wl89+tlXsFw598EOMT/I+3ZY8xYBCuSwIaBJUU
rCAg34Y5IpDJ8tNOTTy2JefnTnwLIjyCgdL9jk5yGgA4593jU3RE7/riUyr46ztD
0mEL3fbucBZ2nxWpAR1bFHVbRB5vGlAqqe5VKuBeDy4CM6yhMm2nnFaBgRoFt3bD
QTGF1cKB7VCLaPyORxo2zjN28oC38ijdoe7C/yGu8WdXKH6nTOnutQEqQNa0+emr
FGHtJG7g4IBsynL4YRroBgjoGxu8GuKl/q/aZ1Ho2MH2ymdB7JxN3xs51uC/Dg3w
K2JumHpgb0Md069+Txb1gqGfSFLXSkzFx8o3d/HUSUY+Dax5/841Rm0XUMheS2oG
ud0UnTWiQpMeE40Lty0km/MU2xYpYt1kqauSPTPEgCylQVgOo/9q/YX3sc/dEpqy
4UPWuv+2DVuTVoxuEYAhSYvIH4Kv70yir9PxFAR9rEotPQHzHpqCMLpBocNGqWWI
QORrCCKZuVRfjy/75N50Q2qRRSKfRCzwzndn6MEbWYDxz7XQepKKnH1g2j7MaKdG
fajH45vKrA6wQKz9gmKhvPcaOcdZxSQq9/wJ/nPvOvl3tYWxTT4vvQBDGOU40fFz
OePLaJw+0J9pThw/F7QoJcMIazqQsAJkYiam5yXb3o3/C1jcwSpBrCMWpTqcXwSK
3lwib33+n5u2ZyIxL7PSjKXLk7uiKATIoo83kZO06jp7Orn9kjHSbnkpaFKQBaes
NQ9/ubBWBisWnQP9mI3ctBJBSVDErGY8X0ww5CAxt8U1VYYwoeMqhTNuYrF6gknn
InWbLJJgnjSf1/L40qq2C9ql6vP7A5JLphKQIvvOnYyhfsbiLIfly81IBPH08pl3
mjNsOIzyHAq3ikQpfQWDZKF+nQgBQeQcx/+eyXHRKYSizadAwAeqAuHjSJ1ucb02
y7CfWAvdwRUAkGGbZhLN8juJ7QkA5SSnxyMtRfm3WlJwwTUqt1fj8BIJcg5zMIN+
TD7hlkRiLUlicXvSmFTzM5D9WgTpivgwbta7nniX7mRIK8sWCb41egYmmACQld9W
DhdFMGflo6mCd1pmod3lFZN0vw1kvqqn/LVuqZdiTdgbeiwncUrlQF3A5PFpkdHj
WYKPzIo947i1GwAl5PyagUDJijJJd+Tm0EgiE/FSlCgf4yd73hBWh7YFjdO7vHod
rwKAtK+DWQlIZB0KOSauC1thirnzMdyWzEvLwaOZWPDnnI34jte5kJyXL0Hu+N/o
cFo1o/IxMs+mTK7/Qa8U4AwFPJgab+MJn+J1ZtUVDEH2btOnTQblz7FAY1BQXSBV
CJTpsH6ZGltIzgzBacBOXhyp3gAOJc7ekqdIhMLdgYLFNSQ8oQaeALb9Z2ejqvQ9
qm1+D9bWyjPB2UQVQ0dH2aQeZgciW56dOpT+SfxdisvE2hrNioLYjtMdQYeqZaDe
PIklat5qdjzMg0fjGHRAJ5xC8/HgkQQ1w6CXywY2+44M8T7K1k5ULSb6WtkEpCRq
c8I4zGc/LvY4Y9qrgiqewQwMYweBgY0a2XPHTD4XqRz+gnJKbVkqKWXCBsZmg4K5
z1UKOIgZXICnWzjUw8d5CCOiB7t36qvw2ktqWEFLhwHWTmY0+PWj7kgsEgeikZZh
iT6pGeo9BcKhqK9matFiOfpP30qqL9dNREo4kw4V0HwaFakxS7ifreaNxTndRB43
FQFO9QMVvSJ9ezyq8AesZiTYPkrCscKW6JnSPweHCRP6RtU29XuEA4wXfsp5VslQ
qwEaleMmKHs8+m0Dj7qkL/1XdoQrLjCBu5+rqPCAknKuo3FQEQvPeMJ/hzH67V8K
I/VUPhL5uiOGnuVkP1Ht/WNbO1cDsJtnAXilcAHLWr6LARPWG4hord4NqJ990UAp
OJLDeslANnzUHyC4WPmVDy9o7Sq9QENhDcGhmS4QxHQKewbGJcmLNmsOx+H73yxE
0+7qUK2Zu35zPGOUjC/maL0xabT5NnVLaJOqk0uf2XXtWC/V7f8/38kmYnLnxnF2
3jQEL5npGp2lApaKAQ7Lt4Zb4YUj0mdZOAo24BbmsdnXARbs5g60tbHlLkfqaHj0
nJjr8f623UJelT/4Z+XuJioqDDJd0c1u/0H3bcKl+F0l18JGhNWQyPSwPQ5zKPYY
3RNLMQ1elmcF43UDj25dmeN48rH1JfwugrRq3JV1gb6E9kzjZgl/c8RY7c6x1Jj2
uVfcoi1mxVY7Xh1iV/mi46ZN9SDW8HJ5rgw32CO+CqT9gO69bE9Um6Jl4thJ+f4Y
y/ulJuCoyyZBTJFkzBNRjgOCP/U6rnGUxt/IRwb5Hb689BWBcf6gcaSB4CBpU5rk
V1NLH7Rhg9RqJAiUqgLMei+6bLhYFSenkeegRqLVmPavCG9xW/5wUkATribDPcjd
XnGiZYfEGzGnzOGJSU6c0YY7wjnV3i56pore9soTUxOli+FmkU76tAEGrBSKR/9+
+xFUMpO6IKQczvHkRjM8WrShQ7weoIvRE/xnbImcl6NGRjkCM8xeSHG/LQ2QQs7Q
KaPQNVEKylOVZNGsTI8xwMNwM0bZVSs9ELmrxCops6QbbxYNCuvBmpfPz4xAhSi2
0/p0Iy8YDSyv1e9UoWDhqYSoukj1VnPSdcKE3e6kJusN2i0aPDfjenZedNEZabdf
8V4aoii8+/woKROw5Ul93OhKLGhl5XIV/XF0V6QtagxcD4BgaHU2H+Pc+fwhr/Hy
SMDmLhJFZ6F72CoVZ9TQfGRkwyZT/N2gcP4SAon9MLdzhLsTXsmHjCWo2f0V4H7S
9IiOn/2uBKq4J6Sf2nrKIpJa7qic6G7nZ0wVI1/DBM6VrDZnDRD07pHNGrfDBDeL
LViYfFP3baarcqA+IBys5X+kBknn9zphhjVPxVC+z7AiClOFn+3uGaLZ6OikG2Bp
ihdqS9Ig5AXY2YzykciVZIYzjilMW6d9gIRhXbXy7j3Z6tItCdSLpFFPTZk0uvsT
3J32iFfNOU5FsKG7riohGI+iTY1PHC4j+widb5fxisL15V38yt5XQS/ZDMOsNspZ
NqF7f1HuUSxPGBdgU/oRKxCFAkI9PXwCR9V/MogzxMOCQmO+nTr3UDgLdJKSX18a
O4WPdOWZulGIbq1dg34srh4UEcARSwm5llJlM0RUD56tT/zqUtcwuYYtl6SmhGpM
mKHfseEWa6xLxqGfQBak2u94vy8xrH/aJVD3Oe8RhOWKll+Tjg2joSruNiBCNeAC
hf6Lz9PhhI/hFyxA/XmQtwaR4ql87m4gSgmF542PoqQ6eDjUO72ZzrBe3aFJxWj6
0+ahvp2ZIQZg19JbSrk9e24pcRgLbIMQ6t8bnxiM6IXuqVh/QreJ6f93M7SsM1zT
PLYwCyrvaYKwtES657Wk+Zn2fOvC1VfKqWxnIdRgXZRzyo1qLV7jMWlBlP53Z6Q2
AAoin5tSsI1G40y58hQRqs2qHV92scX0+LAA8zOlO+/K+2zB8E4dz4JfXeWIFIpB
hMKbCSg0B5Y2dRQunQM/4GOhGVWX4FsJaPyTQgIunmj4ay7K6nkwiVU+pymBozbl
0geExn7HsvFIdsETl0Orxr/ZzlLgy4rnrpH/mkIV2rZ6KD5jUos0xp5C+Tm11nzr
UPbA4r4BrA+lnbA18krBkBInQ3DP5JvcJrw7aAFEHyo1rkSddalNLElpP5eaB74X
xvjKKZsiKa8uTDWBxgtBMmNCkjY9USl0O2QzleYp6BBaxjVErWpy3hCvnfPuByoR
ABlbJxpuBg+uhy4kzqpZ6LGouIszq0/Oze/62ovcwBWh6xFZgUNEhf8IBZoPtQiK
sYU+h92q/AAk6Mh4PTPBZdNfCtRqB0fHmrbruViwZtu1/vnQGN5rX43HmDXDwwS7
d+ZEpE/Bf1wJ5JNPKmG0TYEVKbzMfJqBqvIOuBegPWYnFWID4pSasyF3Tq4rbbir
HPR8wkCnfxyzOrOg4wQwjByKn/74TFKJjm2/6PgMuR2XQmLOj0RgJuoNWgiH3OIT
iOTi95w2w+M+fKSy6aTOyPvkxC1Jh/WEAPxN1vGlachNkDTZDbLvWQiBh1D/h9Qk
G2nBJAsXPFdP7xOTk+jG5STYEZQeMKeXPghw4SSdsaDNn7SefKAkUV8PRM6JDpPQ
YXUyGZ+Aks1qz/dmYgqyGCoIOM5Fv5MakbkYyd8oleJQDlqqtwqWGHSj3TyASvmH
kB7yQUuwR81lNt+rwYYtvILJTMGNCaRoRPcsj0Z3zsJoacVyyHjgmsmcowQY7q/P
pJ/uwe9sUtwCNJYbwM3NqsNdDkkxeQndFOkLo6nVfMM61LT2o3lZ1uQxI1kzuezZ
NRu6UXIFR25heq6MXA9SO3XRrWHk0roVjfb/uKOenTy5lqnAwy4+7bKy9mC8V5VZ
iU3MwIxCZFaEPA78Zl+rLgTPKRYXKf0HrZ2L13IIjNjd/1GB9UsSpBW1McwQX1i8
MlqDM246s1vjixky4gyXe2GsKnxFXE+LXkvu3/72k1ghmIdh4MAalODo5y7YDql/
4ODJp2ndtREIRDEVdO/ZUJ7e7p44M972rxVCpVdbOAP3p5FyNyv6kEZ/iIZgbwoH
DB+mmgaLPGvsCdXVCLWAm/PG88QW6ElZzYMlfVmJBA5k39srGA2aDggRP4CqDnu4
42MlO2omOPNzEExhyD81uS+IxQL0jBUP3jQk51xK88PwvuzswTxnhhviPRczLv5F
1zg90d3fsKlsN501/B4NzoygGIdGjvAQphJ12p4SJ/tkpwmZeoK/BYW5tUIHHgod
Nu4MPySyBmsE4LUlGAC/YxO3v94d/fT5e5WFSj97fVfH4964aNqec97lmJXPTfZn
3AXFo8PgIuS2Ya3CK0AEEnHkwWZ2WCdmoxLjynjFWyjOotTO9xoEZU9NXfRunt3M
hCPvzFktMef0E5o03DOycRyJoGPcgiQvjrR9RHgpapuMrxpjIbNv5ARheq0uvWMM
UGwWPGY1VE+U+TNw+rNg5hegUh4JPSmO6ZuYXqHNpTSCH2KbLJoOIw9tUR8UFZXR
c+lk+dJGJBeCrEwh+041uNWsfMUHsIg+G15wC2stEV5Xzcu/+gmsQs4+KW+zdCcw
4FzhoqA2bPGWKlnr2eNwnct7n05tz7dViFMwuY8+voDtD7go/CfPdiKgc4+q1fgN
Ua0yLFaTzWmc5e/crWVp3giRVA8cwih3rzNm6wRZ5ovNxopYfhu5s+2kwGPdscoI
am5QavVBNuQLDkJtLqWhSTNiMjUNS+In09zEzYeA/N1oXVoYeCkvAgrv+m16lZBs
G2YS7m+VsWggkFXtleGFtIpa2P96fOPNBvUBKeV1INa9ptzq+VYjTZG6YAXXXhJR
6OYaCkZ82LK6IdICGy2yH7yBwb65lNQ8/xP5bugUCCLGCCQEIeTAMxknO4DWbTI3
6k5Yct1zbAtmr5rXKoAI9+vOHPyHGCXvBbsu6UitGxxYkP8VyL8tuEhQyMt807Dp
OBkoOv4u7ts8zuuE0GykP8Twcu8hqTaeIeyuV+8g96b/Si66LtTdANLSQlYWmfuk
2nAYptyq7c8yPJDSUHAQARudKHf6pbd6AW2GNDV3Wzhjho+TS1uNUIGrNQ2iD272
CA3wuhVo34J8DgUg9kHIE0nIFag5GBMU+1MULnT3OnzH9PMCEMHNoVQFHkiZTd6K
A5Z7CeQWePf5FdZknp0QvGe/c4jZGdUU7U/aqFTvePSpj8WlMPmTrrMak51xLhgf
+4O/zYWtkJjgbYZEqcw+KRW4Tc5VQ3+XCZ+bpvJiCAhCSbl8tORYA7S5ZxP0JZR/
6xx8X/OZY6/QsM3TvM0WuylB8Urq6wb/aXkOGvwDKUZ/sY/rHxO6ClUdYUzea1tZ
tS1e2q6nFuojt6vXkBD9/tmcw/6+pNSCkwp+bsJiVvBI7UQr6XjJVwtc7kN3NHM0
uvLpHboDF3NWGfFwTo44oyBxhfiwzne+klFB0bZzUaKTiT67F8ZAIz7NC57Kq8z3
Q6817fOKYzH+irLmIGufH7+don6zcDCacDPs5leTAszRgKsiRXLFS8M005b8Uzlu
0tOBMQHan2gcCniBbrEa1+6jzaorBOIeBH9IWLCfHjqSFgrPEM0iChgxi2z+0l+y
j++a3Odz5VPXC8W1YmriWrDUNy17Z0vTMWk/sQPSYLVSV/7TO297vgwv089ANCwP
vR9Puiu4B+OQyrBWNY9IiL4uihYaDAKjqyeXH0jslfbHOuELpXlsnzDljJAy5zfz
V8Y6To+eL5jC/ioe0OOhYXvI6yHAldMP2EuYTFlHiz0Flx+NXHoEHhDtKaxdQEFH
bsVaxbwENgaQ9k2hd9Fo2dKNhATXd882zVdX92YCGua8OWkv5jbxG73qg+lH6/p8
vPggwg3oGKO0E4gloIOmOIf9wuTPiYg3kvkf4eo4nHhlWDpxjq7Gbn6qqECodnLZ
dVOXkQ+zJ8ROgiuLjA6y5H7dW6sASf4JZN/ezcn+My63alFSFf3bYJvVrIElEEsN
s/5Zku+wKchPyKLld9xdCBhOL/NOiqko8LfRHDqn7z8rMSuY0eOBgqaPqVWONzW8
woEybz12IAJ0GzQRQ3Z/WGk5ITLn3fFKDFok80iPlXBx+4wjwAK4zg755IMhrOFL
3Ywb+2Fu7wRnPVxnVQJOGCwncCT+xSWN0kDanBnvcCcQcZYJJyNdy8wSCJg80cfM
CDOEJJLc1sbtRKcpXv+ZbpDReEnEocUGqYSbi9fqGrhFdlS+clVb5FY2o99eeCIO
0UyzjloIHwbm8yQI53TNhy9er4+EJo3LMflvbjf4qwpXHjfOJLcaYfVNwiysvyZ6
UUMaQl1BC8qdo9MOA4ug2VQA23mTmtj3+Nm1PKRo9y29e7vkBp7O0Pzkt5GLX6x0
nBT5BB2Iml+qyMdzuAAeLvEk6fcrdKmVXQ1MhVEenV7nDq2aMb+lk4ed1H9aNoYP
GjUX8IRPAEm4HeEU7zP+lgnALewVS4u01gUe/9qGSolBEHU2n2rTpiabEpvuBGXM
SSHErLE5o0D78niMJC/MyUmu88o+dQ5p2YCb+UrLp4aN4vmG4lSrnHF+5+9ZrOrX
TzcrJnafvSR+2ghvBf0935XWRaKZlP8WUxLzb/dbXo+a+EYMrYs7gS9PHnEwCHiE
UPYCmERS25yJ9dDIfPZuyhDxZ+HDDVBXB498v5/fEoCo5qAjPY7xcKV4bf/apiqv
kOKubWF06dE+aJQ0KmzVOTWk6ienuI2e52988fyj7TYlcf9AmrY2TFhJKTX2knGI
Y3LSGJBw6D5TSNnSIBLWuLtN7I58ZLuZVnemXz3gLftfb0JCSZOESbcvdHGlbmwL
cpRmmwgS85OSZH+SZ7Tn/UykqX2WlS9ey2goydcNiQIyk/VdmpBnrQXucKeuj6WK
auKVFpjz/QBhaUjh350Bpxpx3JgSnWpvyfYEdYECeFxUMgjKiooHyM7x/A5XcvTI
z7fZRaE0EJzTkSchwEr6+a10QnBTGuHnXvaFXRRes6NhN0kGn/bfXL2bRyE+h46f
Ny50nSKe27t43eYVHDPeRB1C8O+aTilTiIuCGEFXNjUyqLeQlB5oGBjfYAr7zIzE
53Zxe0zms6jGzmlo2Yes8JjTK7SLwyCnNn35WBu+4o3RLXMblKCtQemOz7dPu0VV
dYAvE/fJGL6sdOxSNwzBeI4smyrqKOt9vTfYw//OfIa3d06ZoPPUvH2q4h8npjQ6
qTkCIPbw3OO0Dh6IVhq8JNYl9KUiuTHmlHMOPh3//OFfSzBPuULNi4lRKVwBNihx
EnXz5belJh7uPRkoUt1XF0m8P3PYmXGtLpRJ/bpWX4rSe5fqSHAKvpvwnoRTtJZR
OAlz65aXIiXEmdYAx9tAmbc/eIlg2Tfwy3RDvdhlnaebhQefgCiYufqQpK479ki3
QXz3OKoE9/G6U4vPtC1e2khfv5YVGqj0+6ySU8smuwrY1MuX0mCc2Q+P6TZrS86A
Xi25cIvcgpjdQ3utKilFbHzdTMz46C6SRl9+A62gWWUtS+zxVlUAVAwUFMIpGGdY
iIYN8kAqX7fhChO65t0aG/BCVFnPWrLCJW4KQwzZH3UZaQsuIHYy12S3uHZXPxlM
4X3Onhi4r77ENSuXCdD8eeN0H0Gmh4JGIbS2KM/j+BsWJbQvY/xgCY+rTElqXeNG
x+fwvDOkRWE4hASdr+oSAuw5EryfRz1CE8jjyS1EQsk42wvud46W+LTeLvaLj3HC
O1mwlB1vr5Ad0JbXyxTX5gkPsbty20RXdxllLEr5fG0nsu/1I8rrOfhGaD8rE/+N
KETWdgEyhOZNkyxCK/GJG1Fa2oK3aMfaoxmqxeh9DHiX+btN2eUb1gb/8estpxGq
yRoquIUuRQ7P/DoNhaBC1gwZcDqhwm9XrMW5D8B3pScYSexbQRKGgGeOeqx+PVav
akWVy2uBkMKDTkGcAQXpuUHeNjl1qdxttUoxyCh/euaaI3bZlc/YZDiVy6DHSkdr
H5X8GwScjX2Fv+BgBe5dB7myqSQA2UDAY0iX6ExowAEjUzotq6PvcC2XvXRbY3a/
yPEi27sTx0OOcpME/HcVOQhCQMOtQm8gxLmDOc/Jvxxyi+birqO6Ac3n9P8NiHnE
kazoBm/l8CGV44kkpQVwH8+piPyvrXGDJciXPctk7gfwNU4DMZYonJ7vE78nIGJr
RxRb3l5m9vNtzL7ygM6sZfrQ0dLPZqXVKew/XlXGCVtS33IbJio6TLLUfugZFO7a
DyzKbIFHWtK8EAlXI/cTEiqJK8n6oBQ+VdBFsa5JpGtxAjqQTKEtsgXnDpJ2LNTM
YyVgHhegYDf97OT3Ry35mOyrbwQw1YhqDYWNTMdjsoNGRmi4knRMN/swEAuF1Zop
D6ucwhyQ4TDBBFMLWH+T2HblulbnI47Op/GuXCQVFwuHJ9rlE+ZhRCNJ6wGyZXaI
GZ30Re3o+LXbyksL/nzgUIkBeXlABUTlTMhoXrJG48sztdWiYasEf1qEMhz1XD3D
T6HMzqzoyYuqx+6uADMlDYQf0gKqnEY29xofgmX7Z6S0RPb4Dn/ZG0AlPEzucmKL
rERccZgbC6BscLpv8Mx5WfndWjUw9JH5mZc/g3/ru8XhFF3wsAcX69APx0MS4XjZ
coZtqjpFM+XrYcPXolPrBwFtAzxEzx1zvime6ar+6Zc6bHjMqZ4Fet7voyTeHtg1
Tleyk3TWsTupQUYzzI7ovj3D+T0OA9hRFvxw9UbLvncmaqfET7OIWlPuZDOZV+O0
F92db+bAVYTXrxsTZRZu92I8nf4O9ZS6/RLbNEexomqCmYoK43TOPMxX1ZH27t1U
ocWDrOtCH8JQoE7v1ckEEcPVXJEQ8KFC58OUIkwI1x9kQpeHc0/SRHfbRBj8zp1H
6DQ8iecGP23STqVV1SgSQ/khA3Vk4HBziR4OzdE30KQidCJQ6S8XIwhen64w+3d1
7JsYnXQs75gO/4vVRFOcszXiKluDwkNMTjuBBsmzsuY/WcB58PDqMR+ppDsfCxIt
jP2wCMiY1F4EzPf87c4hYS/SFZumAPfE8+Btn5WX7PlHetS9gOm85TB/qlGm/EyQ
hstRBxaXS3f+h9XRB/sxA+WUgspzrGYlHKjUXUs3hGmSLQOEbsXJgMTjkgSaDDKl
70WpYetYRb5g9RrfEuaBIjRyUAzD81vAHeV2igXYC0yM+qRsz/loftrn/JPROZRR
aD7sFgoZ8av83+OVo0aUKHVK+909viPZzcj7z5XvRHEkIMOqTh/PsG0fTchsiDFt
+68Qg97KFROev8jHjcjfV+/aimH6vv/FHDEmTY8XfrfpIbk+LVplN9kkdUyVVEf8
myHtvDtJWSP+QbloVNyu+mMRdS7sJh6rKw43CVakahl0cZx8QMlHvxufgtI2+mgd
OZ5f4jLa0LRu9JKas7yQNWG1Uj6fSMww6JrmdJ4oM7zXjltywQfmgaJGeMFfrasr
Qpk0e9csWhUZ5Hu+IuHLwME5fOF2Kj4+q/++6b6lWHGvR5xlTQm5hs3rNcCGCZjc
lswfIzmaUaaaoDySFZ+BX/uvFLLqDm3T7vLdzzaICKstmBjYL5MBOojtpUoz0nZ+
GmN7O2CfT/HG17pBmBNnuJ+jwZXJRYzhfTbOP+NTB3kN4Okl6w06tsK927Qw5pns
2eaEGIjmjjky/OKcwy+T2zLW89rM3R7O7ef5pbxyb5rmQ7IXdM/Qx6EI6PLPAadX
PZZN6ndJ24SxbDULcbCWDoGOZUggcuRQVfFdwnqMCVcRXRIxjq8lbxDAYIh39b98
5Lmm4UoyRYlBJDaFbY+x/HVpyj94HZeIFg0MzK4mfcDiEeDGWYkolF89xscFivIs
HFYm3WVu50cnBSGuyPyir2LPWQSrcaZWmoGbsJDaDeDH8yy8BFmPg34aMmXBtczO
Xr9OMfGbHD4Q4Qn7C61JHp0S29mG61bgwx1XjhTQ9TTKbaMn0fL0THjuyC2MCif8
zd5KQbnEz1+aRqYBbAtL3YqoohKiCH6imjJlYzgoydLZRKyT3D0wq5bDX+pFJHU3
KVCoJ37cqMI7G24J9MElfS97aQQ+RZH9SSWOJHXZdZ1iBpusnz64vzWaxJIZLFBz
L0SAbaLIaDxiF1zo/JcdDZx+ZFabcpl47IyrnRyupoMCCCJ5nVB1RPv+mxJmchqn
d4d5MD+OO+v3zrLAdNTOv16Uhmbq6ckHGxxBAm6OyFX3lzFTtya/Nmjb+/0QsDYu
7BDkcl1PHK4UPZnEF7/yRALczVrlnboR91S19hsX5MFzQp//gzsPNabjv9IV85T/
T4Mc7PVFi7D4NM9jymQU1jpHCJnWJleu8WOfgMzkDbflTpbV0B0HJrEJoSRTRtvq
TkqyjEOzfGUyE3eXqgdoOiixq5hZJ48SXcmKEXufjfIDE5YQfjYZar8xetg63bF+
lyIFKPRauZEhn3zaumAAEmf8lHXfmXb8HTwu3dHkQ5M+fbjZnJN7i93xCixEbY67
6QdkUtcfxxezebahnoOtwe+2+2KN0VPZVzB+J9nZdfOvlG9Z35uuDZrHFCf7AB4Q
WtYFfEvvrcY+8vzM57JISMtlOWfn/g2/2k1fTDze8K77MHdRMLrYLiYdH3ijqoUG
lDTL8hvFIN5m+TLYnt7JqrdtIlL4uRCf1Pi7WGl73SQcjaNytULwFQftttA0p3l4
Nwl0h+nyP9VVlSdbXi2U1PNxx1wqUcVn5OZ79ITFbwfBWG95QRfSb/Mqm53pJv4y
EJqNutMjtNvHK98ReQ+WGaNT0RT64ZaljGzeud/dwomTzrk1NgWoCCcfDoza3uYV
wF1krY6AetOfkp6xYlbdu7XPA+Ak9NYuITBHAPiNVffy/TNj5cEnpVDu8b5jaY/+
N4Dh4MPfBu0SClwy5HbEN3cqXSABV098nQ5mNgJPwSW/F9OtKzgkj7jN0KrW9h4u
Yw1AZRAeCEXY0UIN4uWYp9fVbnAu0bwOh9lT7tR73yxJo7mlFSaEGc8LQbu4FgGP
LfYzu9o0f2EaM2QRAklZfAaM0rYIjsdMQdr8UlQ8f1VNFozUf03+JfSOlpc9/k/Z
wSUjNOTvyykbro+RWXmuaPoWOZlrUp0JKSPp+TQJ2e/MX3cG0k8w1OkjIqe728oS
QuiaCFWs473FVj3XyrP1gDMhgyrz6/+AUzdtxBSfd2Nh67kfXJqiSWm2jG823ITW
7gS6VnYucYu9bHeYqNqd4tyG9XWKKUd7jUNNS0EUsPrctUZCH/G2PJbuK9He7qT7
0HNGllb7BPkY6DshA8NM4I187nnYK1cZGtBGJn39MiGlgvokibqfBDqnUQalRana
VX8Mw8dzPdEFea/jzRB9AlO12pH0JkfCh8LAACTaaPZynh6kZvjemIl24gHzdrB9
SAq3Bucb13X3Lrix2CWTXzoNPhQWUIC45bFlpiEIIQmx4EK+F5oVAMN/mkxLOJzl
jKASe9SDADtryY2J+urG8l30c028K53Af1adHYfcdMCOs+xGfe70leXsfiy+8aw6
K4aYKpJlEnzBthyLweSXKrn0xmpiQIqVBrIAnjCULVaNepIqllFnSQicSIsbciXO
txi7cUK3PSCDaEHzvg71yOwB55PLsAcNVVYAQeFeIP6z+1uB0AZ3O4PGC3Y8jqMK
uJspHqWcX7ZbS5VQD8JY7vdQJV7jGsMg8Zoqo5VJQ7DYcN1gSsZb2S85CztZ2V1T
xkQL9czpxhCKZQrELD4oeluOdC8xY2/jEi5qXV9q3nns2+EGCOvz0ejhi4b30ZFk
k74823teVrhnPMzHdszx05gDFqIrOMieYqX8OlBfDb5CgLYv7wgKXF10C76oT3jS
WCvcWrkCFSpGt1QhESbnJprXo4YaMV+uAEmL2a4xcMNE0qEc0HVTTpvNovvY0rH7
7fK9q+9ai56xw67trdW5t1SLvE3ppv6JIIokZAW7KN/+VkmkQPjf+hwcjQbo5lv1
ArgJ9xMKwaYYwtOnHzkWlTfWdDChyD3aHUxbssiCjxbjZlX8OUlY1V+FMsO9+pDW
xg5f6TH/LjFM6s/PoHVutBz5R983cPTpBN5vxpWGygwdSOQu/eRnLf2kRrn71h0I
6Gn7XpCaGira8H7kzssF+QuE2uYb5QWIkaaPgdUIGLuTJKrBa0NtcfBYD+yv7n7g
s7BL02R0PopK/eURiFqVu/Wj16Bdw2bYZXaFhOE9W9slfQh9EfcuyUo1UQQl4KmD
YlQS+sL9xKcwfQfWOxpHSs/ZZTMHcjZpX0ZTuxkG8ZykNYgN+H1fkAzZoyb86lT9
AgCicVFi/72yYLaBLbK+Xmi7OYmNGekpKsNkTxDmMSv0S3cNSBuqI4yNkIk4KQ49
kRhs4IwBuzuRXYDvRE875HWZNnUzDeoUQRpewLJ6YT+0zMxMVhZNwqZg3HcZAaPk
dmZzaPt/rBro6l3wLl/7HL5Al630EDn7r/k52p2ZiNqxyI9ldYWN2peV3E076Iy5
5uafjNhtyG/A7R9q+lrx1fklEusTI8k/UDMEb2Ue4f5rIKDb3hQViUTdzy75rn/3
UKJEXmq1weh6dz+aHEn7cPd/ws88yIfYtqfeE5SPlQxEfAFmvhheGouMiICMxRba
caty+tWLd13uHKbNQg+N/o8Jvm5PaE1/KUmVmJ/jy7NjhgLXDBopyjYup43q5RBb
SXp9XdCa87tcUDfWZD5X/RBmonjihF6t5VrhsRNX3YbsmHTdvey2YmiuMsxr1jN1
9nG9U6JDcp8EHKqAXYTn2EiAhBG17sr2gvZFyMB8j7CNOzo8jMHTN5JhIUxQkHO8
9uXD9tBogyG9OfsEJ2vwzQ8awqsAP9thxS4kvljOByhKCjLdOuAlpps4B7XIEfzy
txgeQIAdO3+c0kZQ2rBffIcDjzKPPjsIIAezd524/N4ZtpIbKZHtcuyb0JOfnPrK
Y2G8qfp7xlMvmgrsBxFJmfl8Nm1qtx65P6U6V5TM8jGlr+6F3f8h4AjuJrKCLCgX
T4+hI1Isf8/1gZrvZvC/WKmxjnlvxDB4BJqy00GoZCbXCZuAPdIk+v4hv25jX6FA
zzSqWHfjUrGJJghU+HExa6aZ9wft4cYucOhiMkj19m+HbPOxTUdAEPDewlUrV2ED
i+VrN6Jc9xPv8kBV7BJRCkfzF/vAKbGqiNoVYRBQT60+seLlh6t+RLgGqCptkJBy
SUv74iFXLjw7CcGOM0rIYpdNELk74dP73z/AU8o9O8DYN5FvNvqTahJEykUckZy7
MXUOsybh9tBGuiQvnu+mpOt9f27SxQPg0jEHHNcL1cNQw+fKGCqiYS132Q3mZXz4
zKYIfBxmsXVWp/mlrrALYNNVtLO6uFXOvXAFAGQtOGWT3bWl4Lz8nrsgV/OV59Xc
faWwUzh2SaKqbUUJDi5N3w6E67nwz9p/+6NBH2MfWIkq5CXz4Vm6iiCSK7gGJ9a9
nVbIExs/Aca3x8+jZqjCRAD/Xb8EWMlIbbo6hXeD0foQ+FB4DxSeE2PcqdPo7qfH
o8ro9eM+MoB0CEq32mvSV3fuoKj4M5yTpVZ4GHw4lPzqDr0q/YzaU7I5I+KltAK0
b2W27GSRlm7jij3JYTaGYhfrOzJIsVsO0mSVuSf0TI9/BPr2uqrHAqFLc6AeNHiF
isTAQ4gsubodfYA0xtg0gvET3hFfDB+3vOvsYvqCBic9gu8B5YwRKtHxfqxl2nnO
GLRiuO8TUsy1TP2EurUyfb1q0jEvLr4UYHvfPjAvsvPUScrKu7q3MnC8ToEvMpuR
aY3FFgzSFcO6d96gNHC0KG8bTXmO4JccL0ugOOOSsVjCQV3QfN2mM9GUFT90UTLM
PS5qhE984ofCUXbTwyKoktEfVoLkhW3XE2ScBSW3ZyEx6shkluZzepF5jsWz7BP4
3H0h9HAvVX2qqB5Ennq89fGm5bPkjaYdJuTg+WWFZGYLSHS6YEI6pIBVxk4dMDlP
7V/4/5CAKfVsbQw3OVzjyfAsKt2I0AVymbl2+SDsoTzRqa5L9g/jUQgmkASzikyU
0x7/zCFW1IZi81g3LyDR6twc2LgBigNKkSBwjs/AtYyN1I/bwp/I4FeWSFLw7GwI
b8hnQbmpNK92wl3WTioKqZIIWy1LGV6YPGtiSN3A2xS7liChM5mQAQywKO/pK5bv
YJsEU6hHuW1moEWpkBr8zbE+bsRebXV7c3w73StnfaKsGXDd5pfzhb5YhnQX0/hg
dalw4mPMvHuM11QZyikFl1Gi8FMd6whuLWq8GuwaJ2onumATR625s1nRk2gGN/lz
ib8ORj1AENkwD3IM/L8IZ3UYzpqf1lBru4y5mexFhts7tUNDygLgCyRGTOMR3nys
PZLx4t6QvrKLD/xPqsGC0cXCJe3MSkwKXUZ4vGO95eTXunSlPqniusL0j8GRKa1a
XLJxCTRwUqFjqrXrAh7VpS6VWcHAq81yMrUGBWUlfz0gEjwTjpX0U/MROao7PQye
coPnHTK2+X50330lqIkKzW4hkQi+sMIF2i7GPjA8VTu+W7EEVHxUIzTl01M2/Tt4
3PfKpBfATyY/xTEuljvRiqO6/SEDJteQBwfkGx/J6ZkTVwwqb+Bt1e4y9YVqhYkj
ZTNzfEQ96cJMzgyb/SXS/LZzKGyeHuES7INouvCQEOIDtlDGljCss26KrE4WQgCa
+FtNs19FRfTcs5ShIV48qoYVfAtDHCtSMhiBsneYJYp89ndyU7/rSNbzKu5VIdWk
t8inJm5gUC/fA9Nivy76AbACwMYbHBFdzF+o5XQgRCKCWTxWZNK9yd4KRibyNxTN
s6XTZ2GwBJ2YIlVnwkxoAePX9NqXkmeJkGmX4BpYOSOjW3G/uzwrbFZaEv1a0PTu
KXikbsCrD/pjhMi50Rtcw0Je72x7bl4KlYVe+JuGqOyqPv+5DKO6nlAjJQqI7yas
C5zmSAKbFHeoIWFkq3+9g62BsuHEfhow1zKqTOoagHNmbogQJm7EFMdoQC9RR6pu
GTz/nZ7H1Br63BhzLw6pLslIRY7X3oPGbegMw+7unTA9fojRU78EqvWeb6V3SKuP
4e5bEi4C25j+onLQtvXJMNl8W2IjHtPxNUe8T04U5lKS/ippx2xxs//qVjQ/ktxu
ed4a5hVQaK99t+Hzzy7um/rUojkK+ACWDkHA+wJ1hBra3Kx1fDEmdMIMp7OlU/Kl
74iKZsfVB0dOI4oSRH0jMEEJ6nmcpaZjAHH/MqocnG7KatJhA2/JRenF05LSrmxD
BiM3hhzhf1B8/fudnJEfKHapqWc3uzAXA3jH2GaCLNdZIb6b/Wn/frQunmYPMiE0
fMfTmPePM8bfZ0L+o+VTASnSd+xXO0A148nzcUOPrvfhaMkBSibj4+noTfSJelK0
FAbn0lUae7XTKtLuMr5Zzl04hYmywrYOOgXh92Ue+uoIwodUaph3PI4rFD6iygSD
UT4zlH5gdkg2eCPAss5BBEoF6y0F3olqlOfnT2WmS0wmjRkALlpDK8p0ftfsj4EA
PEqSWh90EHrc5Ow80ErXSkeChzBqusVlmBV9ji8GWHfiKYl1UgVWJ6V1bWRU7g3O
r9CY4s8VGRM5+7ipCQmkfeNCEyus6Hg7+AFxNboi1VjZuoduM1cx3i2ndzwkaTHu
WPCq3sSbQCaRIZtv/xDZh2Zvk2HY+2G44GSgaxsfjR6cphTfBJzXUAOBO6+IeCcG
0PwPm/Lcyd1YFUw95PolzxW/CoXFGvaY5e77eL3nZZI05fN8dh5Gj+IWXmqu8dAU
gENaYlAVKtxp0eYKZ3qDjXVknCTrmtl2J/NdIZbH0+1wRhCRWmwxnrK2hH68SWEy
L3QcGAaEQtXTcutZqOtMCLD5BpY4JEjhcIs1kes0D4rjvbzOoy8Ci0M5z8+uoZcR
fe5XpoyQxpKJXVV0atKWPcMWiTK9dWhwQG6mN6A+1IWoTEO1sA3pY6Q+B8+rkaNx
X62HSlyIysB/LXsBX6mhysUEGC7TZynxW63xVXhwOlgQiZXGTZsCapvY7FZgqAij
Qd76we5jdu2+WSeO1h/IjT4n95Bl7dvbvRy+DkhEklr7MmaWbUeYqmtmMf1q66Gd
n782QN6wm3AG78+anIIFHTy4tmdWyYehC+R8d5pVQFI2Iw5taLFzRI7Oyfl13Qgb
QPoeXVWUHDw7b7x5Cmx95wvd6x/KMRKjMbyEi6DBCjmuEiaHD8TeC26w4l5xOlFE
AVqXr6ywIQbL3PXuZ5epodAfBN6mvQz2BqxMx81asSoLX7d/MMo+N69jurST565d
l74NFSZRYVF9Ll+OXeKyoWrUa9pSi7x3rmNHkSnZG0fzJzg9QKzZQypepfXksK2o
/bf7im+2UP5zbN3WP83+tYFWaoaSZVX3Khv1zLtUz+H+0GChf1iclZ8kIvh8qMou
uQHNw4CvfUom5LFupGdRiVNYhL/f3emGhiv3yonrc17MheV+GQDfdwTzxu3sFQm/
PhWr1owaoXCqS1+IBmq6r0/f86aoMYlSswo7fMbSPAb4O4ser7/nzmcZ/M/2UFCC
pcbVifIpbQij4uFVj0LIsF0K6mwsooZNahY+bo/bWXWsnGrMTbZSy+t7EnX0P7M7
6873EMiuI3Zq7Lk96nDf7zKYlsKy4W9vPSQkGAHhMsWddB1A+LNeo1eIgjhKoDq0
i2w4TqiRqZjiKUpIocXLs6BOz6+WAIWhohb6j21loBfb7qXhaGZnu85CupiAjeei
AxHV4SIvClAbT00l9KkW6vtA+bjcUYCnfCFufb7k8HM1hRmH1LKPiX5Kvp0oI+b/
WMWta1Kg33HPOuVGtndjOsk8lDbT2L3GwboHxG5aqegrASbyZrqWlEJS14Xxoy63
8jvotalEX26gE+LIaAWVFv+NF3W5l5jDghpwRYv0F4APrjLp9wBx0O2lmj5YPCDj
SE+A1L+O7XlCYiQMhHHZ08sJFxMlvkSUjSEcxfLCljfPlQqAqXxxW29cKAZAVM1D
iz5aP0taeFu2kOtvCp2J6goUz62dsEnKGMnkfloFT37KXkg5YFITFAyxQvkAKvlF
ZxhT2rVSsZNmNQ9ZrxTAaIzxypt2+uUxqOsvd3fK1q8yRFfaeGIkbT6ZVqanLYme
tYp5CwZnN32/k71sdsDt8IWGuxpbNkVYHPz3jiAT8ZsXljSMj1FGpu+p6X5Jzr5l
lykvJUX8uhFBJBeDBLasIFaWM1uUGzHNhuS1kIHQBhVQ+HtQ++xoz5/Fe9MXWkj4
U599p+slZpHqwV9G+iIRNo81fR0EEfYidbO9s9eN3fv16CgPotPMbWcysXLy9sF3
jIN8llU9O4A68ju9bHJaE9R7CcXtNh1Xrgz6JDcnq/brDJL2hPTF3XUO2H2UEKFR
TfWzVJ3iSuB5qZrqjZ42sjq6dDlt9aH+rSVde+Nyk1kuLSOj3b8Hzl6CYdEw0hxh
60IVS0Lxausr5A6aUleXlt3jsP+3jKno7NQMpP/upw/qnN48IBk4nMZuwEO9+d0y
U+aJvJ9mfC8+E/tOVoyQal3qKeb7NfP8FBW47GTWfu0PH/UPVBdiAChSfKKyCNCi
2OO2DKjCZ7JIbmJjvbAg/gzP3nI5qU/E8UIF9TAuxNGGWNTJd3PLmGZleWOGCxci
L3SaaEMmRcdI7R/I1cImfi9aTJM5KLLMMTkdUFxCvAch2vOSOpvGUvm4qzx/CWxo
Z/v9LwBe9X7nUef+62HhfRbIMVt/ENK/Wmu8BeLKZyEHGj3VPjGpW8gUlSLiLcda
E9heya7E2oLjB0g6S0PNg0U3wf1R8FBy65rYd05iPiOM1p0zDG9xFhFsGXRkA1GD
tcU1rcqE6tjRv6kNddmyQKPm6fMwpVb2HvBWZXqXqCVr3HpKff/iE5xRYohH/rI5
gYJp6bBFhqwut9LPpl8BE4qj4Eui90x+UdBAGloiJbfBog9GTizP490OpGuhn6JH
NZ+Y2GPuvwau9jPgO/Ep7+cJhOZqI6p9ggyuOx8npVTkoIlzlzdFnIg99N5HxNea
d1Npe9Yp0KAvUdyU1WRj+dOlEPYDGSIt5SNu2qd5/5YewxGS+vSLXdUBidsDY/9i
xpkpoTJCMMjrbLhtU/r56mzy9LKRj4I7J7jqd9/dV/v8tmcPc3b81wHRBsF13DSR
w60ampkAP92lG78+C+NkhYr/19GG52s5lUnKXGzf0UC16GIp72Qh4M5kH1frifxA
PaDxVlZSyh4LpIiW49VDS7Z2v4DO9CeNyNaFMpnEnOyq23HYPGldi0xGpsd09AEn
KwZoXTSUAD5kCBu7lTKiyBndE7ploA86qUNSXo4JFqULUcomWTlJ2jzTbDl61HzP
gipM0PW/KAPhqcSigSbotB6iiMZ/+lQc/k6Qq3zTrA96oez/i7Jc8M5d0mQuMMwW
ymtr15GfPiUKVCZDjbVA9taeBbSGxyx9CZAXV7ZUNSSTVBn+1xmi/5CXN3IL/5vl
hPseRYEoz4xdDoS5XApraGHpizqfFl79IKm4UsnZw0KQ4JztP5TWwJbw1fzJjK50
CQeqGjff+7b8W+/qJUdf0/1G8vqZLkEFg1E5BtRHxky7GgLc/p/N/ev6YEL6I/jx
kHz6BSHIWjNP9Oxj7EEVoQQ17J719KCbfs5qKnpRaNrsGJ7lUklN35tb8EVC8ViB
2l1v0WupYZBnvPUoZ5NUkH4RQnoef2f/3h/IXjlsBgAma27TvBx61R+aDLo0VPAk
R2MKcNljCNJxU4D3jlhDR1CM2CJO/xCvSqSMI0LMezl+wHTzjAl/f90ZJIkPBrME
F9DaOT5c5OJ+dIgU1L2c4s/lMIkZoH2xOty273cuDszpo8mkXOlzWQAuB0fz6kLv
Fo1YjMK1xUAnxCpLSuZHtrR1ly9fL6gSD6qtPCGpJLW1jZP1f3dTW9f3yNdMNSmZ
oL2hSXcmeqfSddHYw6HNujPexQR3eXsjkbLEZaTRTu3CZkTzFJPznJgeaqwU+cAF
9nup4BkLT+6zS2g65f1dJP+ufzUDrAqFpncr2TcYUJ1t2J0AdEa4oWZX4ZLr4moz
9itVvTBfo26IjAuH5WDWcGgXP2VOhJUFy8ZYL2M7kEfg6uk7krrOiNLXQaFddc2r
57t+ZvmBmXLWjuk9DVH8mXeNEg7J9DdY3T6HpOOLCtNn8zS2WPBCMfSlbozqWYey
5SnZmtZU8UQWPvEZNZGQPz6BfO4ystMeWL9bsuGiZaeGPojoC+LEenSrtWike1Az
5Sw6nGZ9JCVaE2t8JXeFAl3pKAR47YW27V9klYCNYQg+wBuTRiRBFVbZh6njiu65
U8iUQqOWze1diamW1G5tyh4YtdPfOSnWEOHDO0/TtB+WVbGfMsNhObdhlRYyNe+e
yBNipYAcuBFigNGMHM+OKZ9uWt2rZfk3ekbh34LYLxjJaLfyM8JlMu3FWnfLn97F
OSQtTyJ3fv8DXsVgqh0z+SR11Jy0fuf1RpChoXOycBWGfzacfC44/Aok3BjEDI2W
CYZ1yR8OaQ/TGFyT3l6/oo4Tr6zZVLF51QLHBaWp2mtZivaYYRRQWlDZqpZ45dZ1
k830d8z2k/+9scaOGEaU7aXl90ctFshfqwHZx2rJevUIPZaes0OXpwajzU17isIr
MsMO2UhgJNiDD0OD8Z0mIvvPfcPY1mUZ1Nt/4OoW0yeysuOVmDPzwitP15zT6GyX
fDEZwWu5m5bLczz448cuJwmAXDRb6q9FRl4sB3zC3rNf0vauM00pesZNYlvHg/Kp
byoVOcNbPRMbnAaFm4DvSnKf1rRiCMsyQjIza67tCLipBsn90sMK7Xh/BqNw2ke2
6lxc0QwhOgjiNvL5QScs/t/kDXfnc1vvnsi7dGNSDHPGnnEWKgqMoNIyxlhcCmBL
SVXjmnHgYgtEKIQmXV+xtKuyH73kabOGMi2s6HuOLj0eRCAPyZjjPoecn6YSgKYF
AaH+7gtnvQMSj+n5i2hQn/UrjFDFg7hAmJ0oOcyRX1Cu4KTa639ZvToZDwThEsz6
uR87aQzs0UoaXS+/BrOWRIYHguR2nnQFWTPywrFzyMe0TW4eZ2Nc62jbGF8kwcMK
TQMHL+hL3KOhd3DaWXVF6qbMQLb/UAJUfSljT2GDFxU8spQLyJFsFoRQI3TkQbik
cs/pcfxMef1HZWo1XlD1jHWgFl+vUG3bamDHUMvKbkoYOCkBAESpIr/lams4i9ae
/IS8KPPYcL0aeG68LZRJegwbshqBZdzfFS8Bj0K3qBQukFYLTW3AsdcrdGAzsaWH
Mu+QUjGK3UxmmTrXramd0JMTESq88b4tcV7COIUZlkC745AZv72RehnrhaevhbMh
/GY/ZFvO6OgAvnf9/6JSN/HUGiC6KuC+whGi7vYoQLWv8ddKq91cPYyegEBie11j
Gpq36KwXRWPsoH80/t4FvLitbXEgrpr3eKn66m43tmrTqTcSsddfhPjPDVAk6uDc
FWM3wwIsWgFdtwjAgqqlnhUa9bmb1OPv1CIjjfgmwFEwtC3IeT/p5LKowoNkcPPv
yWeLT8r7Ijtw4rrdc1PzmfGP8bY72LWP0eytu141tUMzVUVTLP+6tRaU1cuaOI2U
/Vzx6C8z0nyNBAChfe64JuhnOPAsVjdxANTfULrGbKdhXaMqew1pDl5q18cSMdUz
kzsr3loULefTCX24vJBhX8ype2kmkCDkaAR/WSolu1K2iWTb4xWfg4u+XfsEwgnI
IeMba37dTIrA3eVmLAmkFa/UMX8UYEx62duCF19ZSknom4Uo1iEuKeQSIXkYtOMz
pscOTJgv09e1+9YgUUkWsh6z1w2cD0rzAki8bk6GWy18VMA1kbdCBVFrnheEdwPk
Z4D+GMY6L3FWEU32+zvnldQc0sd42aDOR/CW1/LV09mjyQlmEtJ7KE6vN9bu6dk5
HuO2QK4gHGOahbFSc5/Rsxl6npr+g8lEqWM2+b5jkGGzYDAcRLFFAEPivC28vEny
Hd4XG5ZmFEguz6VGKYOrXcxyu5jwtQ1mspa8ey+SsSi9CG/StbjduAOtYnCn0G03
FR81rOwR7p4ZngmV83+SjGcXhAd06zKBADOkE9evFa5LjWfX4mklVT4PnvFkykJb
HauiNyKHwX2wGVlSeC10lWOokaFw6Ol4L56BhEQzytRiyw1bYfOqZ6QVIrF7iAV+
g5xsXOL1QuwwIbq2i4BiVSBReYgTSoeB0T+w6EnZ+qJVS3KSIU0e8DIbl+Y8ykCk
bhMN//6n1FE+6zYzcqTXvFjxG6QgXF3iDzr5/YU2EazBal9TY3tR0DjvunZ/kpsn
b/sIYvot0PQHYwd1dg8R+fwvpvfztGmM9fgN6MTr9BBbnwwHWJH6QSSMTz1g6TzW
BoioWrpBwoSIUaU+szfONivoGcsX4NULNKjfa31+0qPMGwNgsy/CVf5AoR2Zc05h
EADjlzOzzZeWGdlUi++TVZp1+Rxx99G3oE83IJhxM9EpBxnbpZ1EpYKy5UIfi5Qp
pY7vZkLKDc7LaC1ZAjB4u4gzBMsMLd4Hcfxw+TSvWoKe+2HoLDQ6ziAy4cLFD10f
6gQAwAJYOBczM2mNeZzjrEtdMeMB4DjNQM2g2P5YiJVko0/LiL0TGMQV3pdRLGh+
Tas+1cBaiX9O7q1bA5jii7rZ0P1fSrcDCSW8+y9EhtmSXS/IEJsAJs+2dEAP3pU6
CeYDFjMo7Ftr8YGftNJeoFaLvdlSMlu9cIy/OonqnaKMEk9uXV9VQXOWQBEILyT8
mMUJEOdyB71B/4VMfvHHJu5tLuSCWH9uqfLRYblJR5kmae2bjdTQRqx/8J/p2Yj5
drPgVMb6lgy5IAa7z+zJML3ct5mUJoqYZTtJeSjwUPbUa9gviLLZYlNWGh4r01+M
SAg+Dq0CSRRiD8lyEqtNnwzIgYGvWDvZk/wOyLtQga2knleHrGiwmp1Ob2vJPjEd
IbYdYflVTi9KMVj0PBuJeCKYFijqh8+BpKLZTdEDWWkDuVIRcVnry1SxAl9N4Z8m
gynGLSpbdqS5rULkKCDQ0ZPZKXT6EfAVqgjR3GvUScAoo+UUgzRFz6HPL9iTh0wA
2Xj0mYQ4Mi744kWE6tRHia953XYdBT90uZ09/6zyRcV2z5C5AVkDS6NJyfnzkJP2
ubMxZu0yJt+ImXhMPhvyckgPpvTh083f8pOe7h1m1VXHpki4X5m3qIUE2nD9AqH4
6wTQ6my8t2HlfaTsWdWEDbLbFuvPagRdNsLroVg1eJRewc2EAaJBIKNmz/1WhPEf
TaHct3YcIEAwnr0jIH51jdFjGy2MWZSXLysKeOwtYYcjEAQ55yhan4YWLuvMcF6S
kcYREEah0io2wLZH/FPKbXCRFU9q9Bcc3DlvYly+IAdGk5azkQgiNPYU2aybtPUQ
5tvHiBMdcz7X+98Ctd/nPFsOsh9SQ23yCMX5IU6Bc+92txXpAj1qV3RkDyUwwhV8
F6Qkny5iO4KiLdVCSapJo+n+ZKYz1m2NLA72K1kF25FzINiXqw5P7YyEzBzXhptP
8f2ZR6w4ZjYImH1Q9Fd7hUYsP+p4JiztRkHPWRQAFjJjM2NWjdnG5qBbghxeOk5V
lmeeTPIWgWOx+gGoROGjn1DjL18X2sCf87L28gk3dIsL+1846iFLvCPiNhaqEYn3
Eu/pKTIdERHz+rETZilR1lk8wGVyhENzNXaYlF59d4561a3fQK6SYleMC5+6/V/c
DJT7Bs2byUbH9M+w4Nv3VmZoP9kHaGqa1XnSANmWT4pXeEvP5FT4ggoVOVYzci2I
15oKZ3yxK1eOcst2cG6dUZmXihxZNuVYsvojDSqtKOF2fIOu8ev7iAXQH9eeql8s
yyDfVhlvT7jL+FEaH0ZxqH9EeKvZf0A9pivGjHek3o7YlN+CFBNqRwZVlxS7Em+s
bP6z8p5RXUcz/OnjWI4s16B3WyHtCSA/zZtO9oeEqVovBVAjx30O4CXVDNEFrvVj
mpxLSG3hAkSwaANytl73KQ45AD9G9Y4/u8tc8zxACEl4wQkkiRHCEwVkAERi73lg
Iu096egWTwg8vhuVFojztvqxeShtLC15TNO0O30u66SGsWjc+1Wev9FN0MKICSHo
FnIN3fVS2OqiS2tp1fZwnBqNzpi7DfBBvmP8AeejPmJNnKjygHt2T0J1rpZiKJZQ
569CqB7jVIiQjIKfAoZm2kY8zb+GYFeMqB/I51dPo7Q9q6FueXD9Xx7d7Qo8IVXA
HRyOUjjQQyZRPoLqbygRxru2IJKuBA37fuDZxLC9G+8qvaCLLH5EyGEmN2jlFmyy
jHRVyFg6uzHPL9pE+kJQukVnf8ZcqAR78SbcYJQ8Xie2sV79UqQx9TRKEGATl+DL
OI5C894NN2pAfAK5XBdaIdKvima/72qJefDy4rdzDMpyOIfo+dc0etbgDGxjbDzh
8RTvACKJHg6e1bt83AD4w5Oez748SgHPrL75Z25OUJcKwSG8fv0LIBmMRI7eCapM
5skXM8snqZffZCB6vDmL5VrEkGV7bbCICv/P6Wf3ioePTq0MEies3VbOksZSKLSa
4p0ne7cGiX7JiArLNxZeckdPvlnxVquFJ1BO+yqRBokn4fPtqgalh1UqTVgoVcc7
V37ZR3Q8xi5NGs+iMa1m5S+BnuDsqFeXSX7rXjHVc+gEGTWCn2yHzi2T5myDMykw
Zh4bFncdIVJyNIxWDybl92x+ge1f7U36MOiJBRHXkMm7Oig5Tc+5sdVXDVPWbPIW
dt7pHMSGSeWftSzyCLcLQavJ8PKjPszkuOo/fqNCUpaNdfLrzkxBUEFUJWtAulcx
DohTs/O0f5tllEVyygTRnVkEgsmes9wfIswVvXM0djYEYAOeA+EoNTwcmdSC0wzM
+HqO8Dh48Rnpc9ssYb2kUKjCNgBvjZwiZJsfjdpSHNO3Xc030q28StmTCNQqy6Ca
mTAAmRGANZV9m/UbTnIDoEfqSXLPnov0/SQQfAShc3auC9595sO2GxIyzlWsY1Nx
8SqyzNHMqSA5gQLL9DzW7zG5s1p6ymwe3mrCRqbG2CJF55UvFnnn+Smn92OXH+VU
k01u05VAbhxm0NAT6BOEUG7PDt9sStOAHLpZyPCUlDcpp6hkQ+LBYE/lGv4yWAyE
7iEwm7BuCQwPdzwJiNlgoQBaLFGFT2NcB2tL06zqNDWDwW9vfw5C1UqWpIF/4QJY
cRhTorLTeeMEoyIjshvUiAICL7PP8taANl10nKBw5Bc2cznZGmETReP81Gh7O6bu
EEeVZ5XL7oIYTXO+kz0ySqo/eXZn+X9V4xleO2H6jX+W7wnXoVuDx7SOjyXBmg7e
j55cAe5phxjFFNwGI4Xnfj167zMaqS5HwibQcl6klPM5hYH5s78l7sUQlh2V0ZfP
zuXsBfUwRUtAOKqZnwG/RGpMTB3Y6etoYjMwO6pWNuACFak6jo0hLxRD2nPfNIeG
dS66Ap1sOd06EPCZ+XcSvhOVmPa8FTikr78QGUUK3HJTuBn6j8wwB6VaoyNEYL/U
PAQOXzjizrfMRyLTG47xBbn0Qh2evDFKMXYJYI+D2kPYWj5+xz0s6Hm4qFmuyHAK
fD+xSoIppT9yFOVxM/zLoKgicYm2IeKEOrpwWsShkJSjguKh6IoKhiskSBg2PVs/
qULJ+oXwRsjkx1owc4vPfpIvOiarY/iap32I6KrQlWlmuWNBAqzylc8I9QZuXJqM
ROf4YyDxVQgKBQO/qm9uGTcRrbpyEHYbG5IjdKh6JIeEK2RncVIo9UalZs2R7c8q
a+SbB89PYdfIzrzixE7Hx7ltP9+vfVovse0ZBU0YmWnjSuJN40nlPaZCNLgx2K7/
MwFaOgVuxiKlRdTzHhqsIy+b1pzqQrjZr01ATnGvtr/r18lgS05jLZeOn8l+Ens2
8OSWOem1tv4zZbBxI3YUIPZzXeWAudKpv1/uVpSUuFq/JIVMveny25IqxdhAExm+
bp2LowCpc7bFbdUCYvSgBaXU6FkhLdyNVnc6uu9pFTLraQPN+qrmrrSFEsZmnbix
7SBY6vpWRezuY6GWUmWguKFggB6PjH6Zk+iwFXmJnF25NaY/Q/nhV2ec2Ds44bxq
MazMgW8c9AW8ujmHwxs0Msvezlb1BceMVIuO7dMg7Hv/ll5/11ZmZbEBa2YPX2SY
w+H3g+Xs3C2lEzyo4SpcnOTJAqww63O0sG5QO/bJ80NBKjuIakg2eG+Np7QD3gUC
urU5wpVhmDf8sZCTP5lvAMK+mD0BRKdsftpNjtuc2k0dFzkeP4VF3+UfuS6GNuQk
K/GXe6ajHYd77nmij8IZjriXAQuQ9OuqLkLbaKEW/VwPYhu5EY5+m2ammQtACcHy
aAxxjHJd08tcUnKBHaH9JtGtGSaV1I6nGa3rb7iIJFxgV80HsvgVBuI2rMSaTTTV
NIjcOIX5McyK3gYyIwLn5yocBtDJ3eQHdGEBM3KgQEYqzJLFGwuDqjpWoz3srPuN
X6rsePL5O90nNXM6fuBEhMvmLCjwPk3Kw75HiEsg7dIs5j6HaWHE4aL++iCWjZZZ
RFOoKbVz+fGBI1r3nsdaiUeSho4NJDInsuwi+3nYysQ3PInaGmaoSS7rnz9fvQyG
VoICtdGK5OFvnb8WAdqxUJ/nSDvwRXeVGvZaF90Z3i/rHD2D4hIQOucTp/3TntOe
SGF0+Wuc1YCCtLONXbWbfkgIMou+y6LPBpWf/MWmF664YKtmk2EyxlFer4E3HgZb
aGeQvkgqVwENXrqUZI2qKCAAAFsgGI8OEbTmX4ko+rDB7G9HA4+qqLrpT2ari9Ha
SI1GsaG1L2+RJmfv+jxvrXYUg+4P3G1htAHARjYeXaGsE7v3tEvA8jaoEoFclbw6
OWq+0omDAFSN9PMNCuoR1qve13xJTwNJJPM7BRkFf3jd70aFILb5NlsfYOTLg3K5
KP7IcESdbfwWDcrxNwiXrqpMhnX8O0mka9mOLp8iZKG8BCI/q/Ai296ABaP6Jo1O
ck2SBYSE0fw+zzWamsEEoHRqvI/HL7LCsrgw45HIJd2sqPZwQxpZBhAziihVKoSb
0AHvjP232vm1EQ+pQUp5UM6tQ2aeVW5mi+2mrp6eKe63oLd0gWNLU+U76U0zeuBg
P6rMUyu7zuron4tzdkOzsJWuiHbn4rPZ9PTTKBDCMBOzagp6jXKC8b45EuyV036W
BFmSshN8/p3ogtAkLGIOHXxyktEL6vOiduu/M4Yu8roV3vT3VOrK98tlQTQxC3oM
yTQ+89ILUXO7EtxXYOStuIG5a7puvBU418+fu5okdrQKBaIjJykIFQhfjc/m/Eg9
faqL79esgvEkzvV0AszyiPAiGCsfBzPvVuh6M1W+wIjHkC59EkqQ0eJmL53YvViM
nGlwcUh2K6a+684khxhH5QBYOs+qL+3ooNva5Sqdi7WeEqkTOlRcVZgp5hIGR2h/
p5g7d6/4mlSoCpTuZHmFjHEN9cIjejQ7lrnmj4VdsO3Tr4cna3Ehn7fGs+XgmSdS
GCgRKcMQ3uK38CDMB279u47U0yVRs9GWJ3KjNVw3l3vmnQsaGmxHAiE9cONJ0G4c
Hlg9uSF4g/OYDIthNzRL71BLm7zAoIBCYho0NGob8wdOAgf+O3ZclZW/er5JGrWJ
M/cnuOkmG1r+fO/Qw2vmm1p0x0MgQELP97HEDAewG7zDMxFF47ZNiupsukukjVzc
aMHFnqKrm9i3E0AYpucn9eKVbYL0yCbM6MP2aLQohbMA+AL+Bxp7uAa7cM9RkHMb
pqTPxe1vAXrGP2unj2CXbabqkkdNrnesd/WOroEmDAmhZ7IbG5LzkEIpVonM4TgX
sdTTD44Ileh3XsoMVUUisL9goVnBu2nrsEzkNsa8pEJZtubUc30UQQvS69mX8LpU
5/qVeEDaIQLPOGHEtkmNWKRNFHjyKxOR11CV0ltxohLS2i5yA6VBl76uEYh18Q5J
vrUbN4f0/p++eJjzbgvTHSVoEYcKQY9Q7wZcUebiedhLey0M2t0gs5UD0AkD7zZO
xfSmylch4M4+DBxXxtCOH4uxoBMny1fFGMKrxs15cTA0b3IwO25dINvjW6ORoVNA
IdCcHuC99eQPzTJMwI+rAWeXQLlWKJ/IkU5VmIMK00iwnhcQ6E9MyUITFcHtweWI
URUAWS4MK5hc2rKmjVFJN4PvLx/kuySgWA4JYso9RP/XvcB+STXB30uNAS83kX20
dg5PxWFkMO+L5UY9Hk18UzX7t4sYL9NM8CfUNv+kcelxg4RHos61JdPKm/29XB7E
GifWUcm/OxweGmJNin/lsBnD9ayltS4rRAKcPKUZMnQjCD1Mk8yM3kmt0Urn8Rpy
tWQNdj0xXvAcntu18h3HkMN52LRwek7obTVFHUrpWL915+bAOUjJT31P+LC9Th6p
QdrQ4hkz7x9+b95vzSuLBLjfSxRYRwxRQ4QnvOgM4lfGlSfZ9XTS4PQx4o/vuKOq
IBKMAYuX0oiHZU2+fVZ+/8Ew6T9gKLW8+6BRJzZWbDSc/QlP4ar8ffU4uteLqaGo
qzz3eu4oUwVwMpg6SPH0761knIrI0SfPHja8fMAE/+Oqa2yyrMBB95FrzerS+sXt
P5eu2d/6nVTRDNDFKzz1lAxY6LPHOhhTIk1qPOBmQMJ0hgmYPZXaOwSpOj7t1wYe
vcFc3aAwkxUi76yAKqWgXSvvuqdYkyD8x3TBFN6NxaojkmiJmb4Tr00oJuMOJ0wk
+XZUcl24ycKDYqzNPD+hWAVBD5RljfGXUivTvQ/+bBnLCSYLrserKEoSX0Wx8waV
CXYl80yvK9Fxp1dKWTLsMnbB15LBEloR/qoCvAd1lR/rkimgmNkvy6n5LvHMmg7V
/2quFvt2LDn+fWmvgQJG+/Zg8t5WGQVZOVZWwNZqMK5RXfKCXGd5R85vLwL7/8ak
1NVPZQI19uUSD7LObJKYK9UVy11mW22wfLukGG1Ihju9Fy8RoZPhzyc1msAoXuxg
3vSswCDsJRtReGmBZIWecpdLE3w+gRC9xHsWmBL8z1Dq4Z/rjYnp0JquLwS4+kiS
8T/YDTQBKxGJTKsbGi9Vp+mQLdy1iyOblsdc9sNY2QVVZxVeIg4cS1INljAn6oNo
oxsk3q0WS8f9sjWWtEQMfXAytETtt/otri1d+/2DbjZ1DuTxJ2C1TyJyyBm4JeVH
ELAh6g1NoM80vFkJt2QrTnUa2gWI8x6Q5zEACywkgJ7ytAZC1zO1hPQ2/5thH+Ql
cZpbzAr0rLlHYb1NZFMqDDv3RMp4JdBM3xegd27M2uArdymkjvc+e7r+EC2j1uM7
3bh8OcUwv153h7EYffrw7LHnqUuy3xsVdW5EtBsMxoRpHTik3raSHNDw3c9jhOUC
bSa15iisUNFfZWEmQqhAZUyPMdeWenlndVFjsRpAwlht2woKOR0IwoOQBNaITOTR
cMdg2vpJUhFTzEk6f6/sNv+gRyFXTio2M5Zq6qCS93MUU31taydAH0AUrp3njrVt
B9bjJmRqcyJV5UkhSRJHrwggLjxFkxPb105vGw37EVIiueKLeAwM/Ep1oYbFi0O1
MXVH40HPcIMw6PdUuIOhSDtSFZ/U1TGaQ8M1bGdcoTtvcXSEwyxB2RQkPW7aT+TL
ZyIzeQMUrRLeorchoUG/edqUn0ceb0j8vW+mGkxzBxcSJIbRMLSX5v3OqHr4d8Z0
kCrjCkm1uvVKnAVKkdDa7f2HeaOSIh0V1kBRpkYgstfwzE0Ch9/mHjpycsMJO+e1
fP4ItKBdvzhRt7LSyuJwFsjSNAOMf7LfTmdlKJWCSuiJJDN33w+Fx383qJXGVNG6
ck/lpUeSYhTedx58xu2Vk41QoPmPccKQjAxZjNEPVXiydBKGukYnCdlemCHefogr
4UVmYIGc6n3bTtNvGqAvy3zweQsr5wAn0t1Ac+jeI+E7RchKHuvgMJZcFZGqUQh2
JYJ8vVhYKner34HmOJ0y4lahWUKyZDMfsQ12yHdTWrYAllK6U/AJ9T1eNDVVcHIL
cNmPDuFRalgb+AsPmS2jEBPjH6/58rTI3uAMYjYR/CLnoFCKYYQ8wwVkJZTKwESu
FWxjOftBB/cTV4y1Pu2qPBLveI3L+05XBpfmHq73NwueY9ymcrLZdPYq3cemksfU
136nf48FEOJKqVzDFIfpyh9l5eFCUvc5X4Gqmv5rNW4KE25XqLIpVoTMWhtIp51I
lCdIQQs2YEY+boCpKFmuUKSyT8dqy+en454beD6BzWtJ62dr7jN+jSffTxgSbW6L
+oSKZDQV9ul842KHjEV+J0j5gk0iwlTVuwvK8y+hDnz3b9oUv7xKZ3tTr9UaY9Wa
9E6h7YJo93nu4Oi16W9HNqHEcjvrzlJXZrsZjpRCCoi4p2mOAd0VcO7H+dGyH1+G
966//gf4crhxKKrFBuvLLD7C+6yddSjzfkbVCgm2itiCbF4wpm9RjkxnpbscSDxc
jmp3zl058bXeQNmlSvb1c+D0raJprcBTgTTjnoyLt9mWq+D6rpZxbSrOK4jLYtkH
5cFRFBvelIQwGgPNOlRofB+GGGAaZieJX7udkyQn0r3Pm133tie31THKXcr7vJkQ
bE5KZdkhXJWOv9zcUMxt5LMudZZ0o2tPKBVm8ZD31ufMtGHtRTt81qnQp55XzWpx
h91RMhfhUHExRPhvmkm6/NksYAJm5mumvKH7GrCGdoYgk34K2wB9MSJJ6wcUQNtP
wxeuWxER49pOm33rndMbdMal4RZ8CZ2DrNGjgNlBrzstBR78MwxFU9raPOQBU2UP
TnUmLEMwvh2LNrFwoi8yc76awfhPAJP4nHrPx2LX/h4Ga/riwvtv+8Ifd9d/IRJq
zGl1Xga6Nyd++w/rxOONYpk6X5xEcLJBnpEtRZtlexiHq8p0Egg4D19gTvtFJQ21
T2MFk85amEeQMZ/YuLe5wj9g/Z7PTi70fnYtGUGxrs24k7akEx6b79IiwM9MMzqt
D5ma3a5GbGbZb9VUlwxrCH5hIHqO/jP8zDA2mpKMzV+YDSibu4RqQ/SXIqeDVnIo
hnsvnhXjySv5Ab9/v11GUzxjguXBqW1cK1IfGY3raZ8UqDzmE3G92tPc07FtMrA/
/KE5PXcG6JRxCWZIwSHZ2ufcgvQThV2WR1w/kZpgvVsKviadYOfXN9oxK2ZbR3DV
Ah/1/qU6iiIV2EgjheWG+qEeaNvG+cZnaNC2QMUGvp5VZpJYQvXrDtEKSttm0oGy
YCSVrfo4hQKCTz1FaYs89NyPxtCIuAr5cf9EthnWVZBAmvmuuylDic3f8hFUeeSE
UXzovRDO5IQ8dhgSxW7bZWVDEGwcYdOmYjSc8P6IlcRP7onKtFeoCGcIIa+hhZ//
/0HLcUaUOa58djtOgDdlSAzXrby41y+bsFci62XLKFFcIKFEDWWduXU3iOJvcm/r
V9ezm5Th0LCT8bK+I4InnJItrpAUlUNXn0Kgi2FvCPy396bIigmhTD9SgEyd9+u6
2jXh/fyPhWFeDztAHPk8gKcrOy3GyKlwOSz1t2ajiXOl1si1TXm37w9LDPeh7lOy
JE4famemHRuYbDpb/2JHvTmvcgoyIvv/H24PaR7TxTQdVkkRrfY4sfFn3e797j4i
ZhofLCQmiaZkjuxWtEEeuC8OIgofdFjUCfTp62CVKIsNU6Z3WnUEQviPJYC1WyqZ
YBu4yxi3eAWBUxnP8XP55ZbUmCX+74PVdzyNl4B3rWY1YPKTaD8nD7Wl+Pdvyibv
PqKV39SnZj5xPVqzaCuqs//SwpWS7kXZfkd3VvyFvfk5K4M0/JWQH/YM3L+LS3JW
K4OireP/5CrqDiZwxf8TVSIL6R7XvSPHP5u/VxptP/vKOXL2Lobc+z2AS+BdQ9WV
a1bckPWqUeO+qA8FecCRw5LjM8+OuKCp1Cm0rASIoSJhkYprWlEcdTyAHvgBkoGz
EY0V1fhZubWhMwoo/ypLroH60CBcOw0E86ZTybOT/N/ZRkE0IOgWjBgkAbSpBcgE
LZRphwUlgteVpCssiZEvOmkgelbZIxpjN+mp7BaOe8RRfhDE/gvh4BERAAQbOyAA
h1JYo+Y0LERusQCZAGc80GWkijHNtKjo6P54EPSTFaFTO3TigSbc5A/umDX4vcx6
JZq5KbgKl0q/Q7kLqOuXovGHY0Q29q6zOMmIIbsGni1oV6oDrdoqvkAqHxQlQW9P
PwAlF8qrYHtAXEgw8QP8JS/y0DsJtijOZ+hGdZFNxDyvjed5JBsbaGivgGOClCuC
LgpFBIoTMYSiZ2q0kRp+HdXUFdureLhXwFTdjO2frUAzVuUHe+FvjOuBSvK4xs4+
Yz8rDuh/3AKhVg+KoQvFRngJ09Vh8736jaZs7yqokRDMNX/A68T7AshVcoqPyn+f
eafhBuqSsCdyoCOV93pWLIAKIFDK6eUvooU4tSALaMAhNUeR9VzIILlBct5yudyt
vCbdooYDdYfexPnT0+4LCMaNw44Cpq2pMMSheEfcUisbtynjdfYkvpbF9+cF2bmH
6Z4VQa6ZYp4/leNi8mwL8DzDDo0ROyogyzSdH5d3CcThK8kwceMZLgmdzsxnSyM4
mW44Q50Xe1Dqu1eHE7qiSdFgx/kGjaHPfbF7jDnRBh8xS68y8I80Hp19618r5IL3
KHmVm17LSCVNNIscfrI4NbhoktHKli73qv/iciDOAxsz1P16w53Q6vd/SpAc5eOc
b+r/cqrCSph2PaJ6n+a4Cp6YMxreN1dO/WB350/xBslmSbyqIuLxXetTmOZP5hha
OTocGOVNs79LHS4oLlO2LB7TS9DSlbCJKpXVmZ7L7BwozNpCyi5Jl1z0uWOIjMfu
6QEe1LgjLAX/M91r/xprVNSDySqnKUkIfE41F5FDiWfbXReNDQmWdh5ljOv8rw1y
0Hzqk5BJo+hr4t7H8ENbW5K6LLLtvZ/9u+GSwvRuZ0QmaEuMWr7IWD2ZzsNK3Srk
w1grYu3HyXXitpTAI8IanR9LTixCAsAiplIAEIZNBFAvniFB4mCIOP0J9/m+SZah
+eJkb3A3aUwtEpNxnFsCUaDE/GXHhSl8rxA8GTlevxiIzVfnpO0+aBLDxN+/XR9A
mC2/NpDzpmqUXC8jm8/wEZXJiIjY4EG3eEtpSpvpifp9kRLiIGRdmNhmZSDAZpXM
8NfBdhHG6EYk3rrAnllqjgmQDDvvx2eOCJ8owAdkk0nXlUey8RnlTqI7pGH7Azy+
5UU3X9gmJ3EC7zNClQeITPiMFOahG50fLd+E1KlsqAsF3JEpB/+vg9C5uplUcEkW
vlMDi4LjmxFW2TUFgxhoQGEG9bKDmREz0VfkQoreHl5K00ZuQDOOs2n1+8bvl+eZ
9oT/lMDxi8DLSH7w8pHT9/RMz+xT0mvhpNsMBNj5w0HpLbZnOaIS5UJ2vzo71bm1
TLNfgaftaVKioE52t8Yue5D6ttqcr+vhAzJUHJMHI3BhUf4GqG/t2kv4xZalhfmB
njENL2MfywHofzc+ruX0jBzz4BklhoHiM2E6qV+JBekuZG8d6ri0bukv+otn128E
6teY0ZZh0DZZWGRsbmeJ4p34f9XRr0fKLCE1Ihw2deehWBobOFOT/kgoJ1wMmgWp
6Fc5MFBcIOTpdkMYOkGToAuw3lIPeJr5KLlEMlNVfsL/pkzKEptJqUp9pRvrLfvD
vKRVBgn+ahPLALLCJKC7Dj/fdUDHIjGKf4E5gM07oOWq9kUXgsh4CaWgYo/k9trZ
UYdF6gj0/e2GDEyFjnQ2zcJoIhQe2AQdlL4PzKCBl9pB441TKQKX7uhzSo75XX2t
4MXfYZ17hlGMxlUwS54YYJeGLh3ZcUq2Kgj/fOLvc+UvK6YK7e8gYAI02fothSlb
7Db7U2d6CtfNtQpHTIL11SkOWutvmRC7I3TRZ5K9n4AFUZtN+d5Uv+0RH00xK/0J
t2LR09lcZRvEnnjE7ZqwUeg0lRcQ8ukHAFp7fFrDWwtz1JnwMZzMPAVbzInQGe6w
pMqG8EsDi5J/4OY0giUTGJPFOboc83CxxR3z5oNZPHiEAGAyTBkFEuX9CBFqciX0
wi5YM71C0RcSPIHJpoGj64ebAI30DgTSeYKhGOFxHbB0vMysPRLNV2mxgtqNVSz5
3wwDIMJZtolw785TgclJLQaY5opB2e84GyrXkW4ec+/LrhdAg7y+WJw70KG9v/zq
Fk7Ko6vPtq0Zp7wj63kWXFgZbW+8vFbJYPZmRlX5iUZZLyL8TaBArZfOXHHocNNK
SVW1mjnaDrU7xpQ3GuafGT5tbSHlH9vm2abcTPg2AY8ceEjmFR714S9yEyMidf8j
uHyW0QJHPPy84FO+tvtYCivOCB1SPaBpI0oIgLkGbYcx81al/KF5RlgRo0qr6abg
onj8VGmPxRU+mkvplQEjvB+2yyP7l3saHRmbpl4E6KgySRGMbPB47rtOAufgGJGf
c30XetTt8cqmLKaOkhtq1wP110em64kUYAEleyLjc4WS3lPKdS8r2nqQtgQ/gckT
cHy8yy5gDT4zobjBGE5ulfyvKvV7VJHJu2NEmYRwrdWyimsgn6bEmg2CiUEU7GHS
f3AWGXkkodI1Pkz6BQMnLw4b81d4VJd+x8hX2W0k8tRKRFgWpuDJexU2EVGUfG8C
genGfYEuJy5gMEk71lkEXMATUXzw5Ls9vQIqroa9f79C922ExJq2bBb2MWK5QqW0
W8tqIEtUdtmHwZw6eCzdBpLOFPeds+QR/2agHLZ/3f2V8Hvoof8jxqk+paqIxg8S
/SDD2V/YMnmsXiVBPScbSQEcfR6zPENM+7Hem0r0dMUs7C7wk3nMWZTYdfR7NrSv
3UHojj44zMfb6NCWdPFkAPnALGhOkkVeJCGafuLuJu1Ivs90XbzB+M81QrFaWWeB
2R+24IWDIjgISj150VdVMIIMffwqUXfB3dABc/igSaxqOOUgyovtIVNrR6ps7HDE
b6UcHJN5KqQkfEwY1PEeueiDo/8VzJiQxmGkcyQT91eSUHEGb2XF7C8xHGeZMQ9+
3an+mdCohLnljBnl2aj6xi/KrpQgSdhURaIQ9KA8i9Y9u3OJ209XG3lUJOz9mEd0
YX0fxh/1cqQcasDshvBm2i1E/YQuwGngCXK56toXnwzCUvhdncl7igr0WT98aqVY
4t23dPMKwlHK0CPly8wSOKhU49XEjCeoWAi2MoSJ79eUBbjrj4B6Ua59Irt9exnS
F98vBJTWgJDqA4jn+e7QUkWSIXXw8tKh0OlXror1yGH34wjS/DuTXb0ifDtB6RPl
JyVh2XyaUfUYGZMefluPH83sSQTb6MfeFJcVYx0Mtko4cqnxlHdbwiAGt/Gt+jIQ
zK+Ib1XsPzfYcV07xp+tpVXO45dC1ynttqVD5guQB2nxxpwLhSVXL+1NmVTExYNl
4wGLzUpzxU9pBeO49rD/g5w3XRCwiNYAzeQ1HvsOYpsquNWIuIcnSBs7wvaASJbB
60uuTe+rsKNyL95Oq61vnuSFqUb0ZL2lWLTUxB6NaPZ1Y7XYhQ0t606FrSfqFPqD
0Uz7OIaYYHd1TRt0le85x91cz4nPidQg/U8dR9Q/16osne6gkRuUBeNJ/VQ374G4
qXCduUI7BAJjPMX8WkOSoMlZ/hy0PPuO9w7/dYDptaQgdZxz0NHn5Akzt6ObGZHI
7UeIziexO2pTo0h4axzD/TP7+1K+BFID9Lxget1kE3aSGZ4VmMbmfMjujbsHK2On
l7dRBx28KivQJC9yTXK/HFo7XJvPb/pr2qcmDCP7fUH9t2orOHsxt7fB4YRcYGyX
W6IaUiVNrxHs9tHovfkJ3N3nHpQVa/rX33/lnWIoDUTOjy2hj62kZvMFBrvGFEru
Zq63lDfTJ+OZN3Gb8BIjwuHeiso+ZEvEP5ZMgHeCnHBkuDJWp94O5EVTHeCQiA9Z
bh6v7KkE19NYGcd4601ZLgzaczhQFhEami5er+gQlLq36SHTLah4Q15ghJcMEPk/
eV0R2VfXNAdWp9DKr8AnWSKDG+twOQQR60+fcBtnM49uvgVa8wf6ZdwhdabgYito
+c0N2mRazOXTV5KeXPxbpl3MOhSEUR8PmmbVl3/0PXDwDYHPuiq9bhYdOBygmRAn
4IN/qi8OvibUpExt0Zu47aR9BRfNV1iLIbO/pSObSJtWNzawBZA9LX/Oa1lneAMI
YnNApOpHMUecR0+m9OyB1g/rLo7bGvAMIKGYm0ZShtHt6FrZfmzcgckAbNxGS4cp
d9UPw4wAsn190WO74ZungfoAhZIf8GE+nG6xNx3mjAnLwPLcOFkWn47MpVoHSFAk
J0pu9uwlDlrtCuFYSdS7mwkflnGTQZvkYQcl5o3dOwfWZWnOke+LREBYWoeTFfKQ
pF3Pgq8WTJmEVws298Ta5V9MGj+VIYW3D5DSJJ0k+SeQS6RYxUF/vibVkBG6cIM/
stjkjckLW4VPCOFMKE5QqK8u1KHEy1vwtLlXdxDkBgpCXusdURWuzDtMtZcNgsXK
af/V+p7vEJMBTBEG8qVQgKaKC/+bRJvPW0fDdeSB7rJXMnpffG11gy9nXmfsON2R
2Fj32uxjXy0ZzRaFDUoxOS0lKAUYe3EL/R6dUFw3DDWxXBS5XJurB8/l8Qg3bAV4
USajGSLdsc5wYRBK8VQ2Vb5NmLtuwneA7YKd6xYzgQRi9+uYr7qf5tMeuK35gtQM
gM7LKM6kiwvaeHBQ7UnepF0GoDFCSj9mTJ/h2NL2O42aYNccmmn85AYEppqRKSNH
PtLPhICbAeMblEITHBlalDsRyQdMJqEWRwI7lRwWi8TDsXs+jo/7hvuuJ9/xIJBf
DuJb+ioC8hbwHseiaHEbDG0HR22U3eqTikCxGAHlCwT0NeYSmLl7J4/kUpGm3ImY
FTBLANN+WQNtQUd42H6qHE7SbeHSIgNAbd8AFLE19fIGXXr0CfEDOuChkEXP1+2/
aTbaqIeWbb1JEamwN7bjq3rTisnhOQxekc/UIIuojdqke/FMz757WhLXy796TFBR
mHGwAivr0A93CZi8HVjY35okykYDpAyMUEun0Dgvuf8YsCDd+k8Rqwhg3H20M6B/
lOV2BHaPqtf/yZs+/iwJUqzlYe+/iGnpSgTCc6cE6xj8T5qaX7LRXm2+/UR3m2Cq
SM6AOLywf6NFY3NhhX77VybVcJaKhTE1zTxHW3u2zQ93dZ41O+Jh9O5BSCmWdxOc
sA4jhOgVHVrzzLzFhNb39TPwruoATu7kZCmN13xB+OGkaCFnhC3DiyeGVsYx9i2t
VeHdXN9mgU5L20GqUHQYta76w9e8IPlkz7l4i2ckfNCxejpHzQl/lG/HQe4eSiIj
jUd1fGDGgfGNXqoYt7CQt2kCrPuR7aYXqD2LaXe4VywAdPgRX0a6AfpYjUt3gQkI
wS9/1KwYwPKlOTQDLGnqJrCXIaayHC9FLMwpkggVPSYHC0+gPffx80BkSzLra/kk
gJqk+hDPmbE7evY0kUEHRSs6lOEkAP6GOH7DcaFCxo+0kaT+gQPxZAXbvSlQvTyX
T2BlIWaZLSKGJuLGmz39qG8MZsRozvLQ05SOIKQb785Ema+5Sy/1yN3tOC2Gvv6H
hLBXybXQrFd4IptI6ydjoMEql53p9HpFfXarz/BqggqFt51uZSHojE7ZVuyxBW+I
dz4Hkoq/aZQU0n30QnHKm54AjhwQkLr1hAmDCa5Lt9B6xoXI5CqW9HX5ZFIlhAlP
c9bUDXdWyJ+Ei+ekFo+EMcmUdx4mw6sqKbsd1gGl0J9jMBXL1JUVsp0PwLJZiSiM
ftQEHCEFKQBhKVnCqvjf9TUEKqpzJHkZ6WN4xRIzFFLWewf6GVVTpWT/LdqC9LXQ
lvX0GQHG57ug1PsrUULS4FawQVVKbdUs/u6cJsS/xXLR1N0ZXJXnyw/aT/y3B/kQ
2S/ZIyq7OwXSmXBxpz2w4TzlEybMRc2r0u/GHPqvRqU/zMRn1tF7UVO5Mgri1vdL
4pGOWwpOMvJndxsLfPFV6EP/p9dyJN328Asz1VtFwHi4NrbdRGGI9gTCfLHZOjRt
0M+aNmIRcmAl/tfhJetuqKdEuFT1GyzduyG6sVmrKZ1QgmJ09iApON1bAzlsZuml
IeOx7H6pXo8KfJg5fjixI1V2peIBcFaoMg9GQGEnvNcQfunZz+4SnTP7wXjeJDDr
tuNMBOL/vwSpUHveagtbMHw02N8au+gIUlR4YiF0wSeEZUH3NLbCzON2Lvf0FjPK
qvXsrY38vOd5SpewrTAMPT6pl0Jft1vQvT2HsKnIOOknQppVOpUkRxIdUKA/LRM/
KEpQNLdLex9brXQg25mLs7r6vKR1DCpxCbYIvYj2KyDQMmLGEfOwIcLzGnKcRrs4
ZkK6wfp7UpinA1eCwTJjMAUJApsfPjFX1WVgoxWQTKZs9PEMhpfdYA0AWm9B3xyZ
zyiPKkpak7ZBB/vhQq9leKcYA7Jwge33e5IsGpwzAvuhxc6daobQlVJoR83jj3I6
BsljmYjtJjXlFmEQJy4B6UgZQF8vYo2GhH+RyMHMpCM1pbZY0Ql02CfhzTGPY6mW
uK70WtRKsfVciuQDleHWnN//+V55GgA5+2883/GvS1B0YBh8LjbH2GaNNYfZ/5Hc
WnGytnTGDVL7svSRTogcrpmx2m1gTlveGKyUesm+7iLNhr7+u8YL+bEpYcqFRYcZ
7J+JO4DQVMZKR+/H4YnTz2617TNKnihmWSz48iml3EzvdhXGkroIXISunhawamno
uGek8s6ECE7/dHiaagcYn2lUtADVgLZTf5i5HEf/a8DDx6ke/ax2KvJ6Xm1bKiuK
E7KB+iVEhh4tTIchC9Neni0w25QOq0lZCmoYDQHNAL6zpL8THQ39gYvs+XCCbXTh
Il10PnT+VluYbZiL4YXNHIOHQFrsmMvqvjxxy1u6tbzqXhDlgMunR9Lz9ueADKp5
DpExURMgcXNEqH/oJIxeV0FiSlvt/rXvUMTAFlqIVPcHHyn0Wl3ojuZ6hJujha5k
T5/qIBWr5StpkS099CS7AqGtjh6m/r8tAxVsiE+Vi/CYi6/c18M6pYa7vkKQ6gpc
vutWSnBpiOqvZ+GspI2dqNFsWvHyrRSNv703enkkBxmP8q+pVcTUTOFVKqzyRuSv
U+/uaVWfHVRJz7bk/3Xz1T7wE/Rt3SF7sUbCj5T+O5BAH8mVciRs9gT1qF8nGz6Y
18H8JNvW/kTXK3ycsJZPXmQRhO3fM9iTYX2lbiJvmLnZzfVi1t0yrZmYPB+D9fD2
fEuQdnJWzM6/pepFH9n5IEeyYMcUU+u0Cz90vU5lkVGFms4EmlTZplQvDlsXeY6T
Nd4sW1wNGCuJTdfCvzDKjR+UUymkgxfkGuqyu4KMqNMjMRMPoqOshmFlx6P0dMfg
AJsP2fWk5uUXfs4M/jyyy/a6Z6dHaHeRgL977Nu2G7gE3912Qs+st2iWU83cQ4RD
JE/zope3mvdt0TpTr8UjZCPz1UsB8K0a0yIvdXI3PosDhnu+9fQbTpGnhiLfHPol
zsSUIAaDZrqCHb6VlTUB64jX/gdY2eufpN6tXSrudcBHB7aMj67qF+po31QgmcYA
PN8ptTUuhZA5yG0OgVODad2Sj/cMs8PsYI45qb8TT2twO6tQekKbLC6JZLTKWXwo
Nobm+hnwA9zvvG5cfgohfKJcjifLmrXpew4Ou7Cbg44WRpWniTHQdCm8C8rtOe+x
LZNi4e/9WnJl1phorB4L9AUj+4iwHbE3FQWADXt3Mye/0WtvKAFkX/zHdBl7jAwh
E10NWA/zNl1hfM6fHVAL7I7C1Dh7mSX1ZxuxMFuDigIYMfCa//9zuN/RIY0YvEqY
u2ebQReYwJDpLVqPfOPX5A+Xzr2Qdl/vmM+HRPaLZ3GnRvzeYUXW9guSP/XK8MHy
S1Ri2PECCJD10oTCtvvPAV5GFz64wwNPXAcOsDm++4C6OAERIAwMsu1QIPilRUy+
TlUiYDuV7iHixKgXbo+cNTCnsvBQOuc7/n0tJ8jfqdmoNDU8y2rTkzTr4ExnngwW
G6FFlD13qf22w66XQc4azN/TuobBb/pO/+GvCxUfkoWkmX7P4RRqULQ/JGUOVvhd
cq6+nhvc9FwgG8F6XnN3yBeC+MWbzZL6ECIsR96ddTPRigmg0izIbQMZexdm00FP
f7j5CilB9d0kUbjQKHeNpDMCMpol0P1Jj/1NguI7/SThbdCsAtKa2pnoMQHko6nD
+o+hpLyn3/Gv1qHcZ2Bo+Gzr1InL1f+58rLReC70/+xSBYK5q+SfbDxmY/K9KFBs
808bP83fA0cWBhp5o+G18AEi+iXsiE2dEb7KxBGrl/HzmTeIyNrR5/5BZTeedCB+
Vy6yCjvy2AfTe41eIyVt9l2Z4kXliQmq8vRYU8a7f72YhCwx4hb8PNNb7oeoaaW1
KkHiulzslfie+GxYwHCMxEpei4BwS6j9B4kuBQpvkvjE/WVKamcC/jnD1ztsVa9N
EXF3EYbFvtpkXRMRjezGix0GJv+GN9BlsU0dSknj6NSsbn/MfcQfKEwkXGeeO9Zl
q9ovIxQdiIUAl0w7p1Zmq/rUiUovzML5obRjYyWaxW4N+X3XMrVypu1YsF1p29L2
KqMg/FaLaFcpLiJkDsRyxSJPanLyMJQpjESkoJ9iBwf1IyXIdx4J6WWFZUCRnXIY
yW6K2/rLTKmOVwdncnR75dIVBcNzBXd14yXBn6B3wV1Sbq4YcCe+tZmNbVaQ/zhF
cQVESJ2yeLvjRVc09i0MKmbJixN/5tG9qUjx/9O6SAxQi7u8vporu9U5vk7e1GQA
lNhmafwUZMMAnvEXrtqwMhr2icEI5+nqkXFWNxdlXWcSiG+MTfW67uZAeQitT3Li
DtlB0s5pQ2p72RqHZVYl+TvqE1Ib2StEWeWoP+CSIdYHu6CQ5mVnKxCRg+7hhuqQ
NsGpU+jK9jDW2A/zJaFZPogzy1sP39LrOWsw0F+aiND6kFWxHTqzNKcNdegHY7JB
d//KlGgvXgl5L53pnIKerQPv/4zUz0cRHGL2g4Wo87eFdsqOivJ16eRRAW7J1EjX
r8U2tFDpRjJFwmDwOJRWuqmMjOTI1QSLC7sR1Si6Tu0YVlkEBnsjjmBVm6BCgAzD
ex4n2tm5qIrbXV1Mb7Y9czLKTv0jq+ZW9aods6zNvxKqJaaop6GRbHRTEoQjusJ6
AEREiUQNqwXJ5Dqvol8iqhthYLPn+mSREw4dL3NNQ4J5p+w0w14EadHDrNqc7Dfh
Ptzmsty8VdwESNvrNrFgho6pRRVrYEAFtbNNQoHIIWrAd7ONyYDPlOqlOx6RP7fO
EiRSXaA/rj6FBI9rldukuQssNrW9fyr7KtvPi2GMNEPXdJ5jJLEzvBVsIx16n864
rBSk6iyW9AyNlTPdMUFYdEsgxXaqhOQzMM+ypL+gk3DZJydVxUDIEKjBCbtKtvJs
FBE6omKcP3gs4aKqhyHZeWkgamBemmwWZLtBPbg9EdpiniTfEanJfe/JKYMnmGmQ
5Lhi46qyPP3rJ/nHOerFtb/4Wft3pDBW3jtJDn2wx0490SFNTaa5loWHykmudZzQ
KlcqyQ4BRXjOCW1BNBPOttiQ4PpESSL2V/UMT9VqsYzfe358gN43tXVgstW9sMYm
IYmuKj/vcCqz9gTWjp4OpX4bH7ERdYL3DPl+Fgj8f8d7nFwzyI8qUiajQHv4N9FH
+11/TTkV2noZqScoVLUzKTJvAShW51y/Vd/emWj5DbzuMxOlEb2AHOOrvgLA3u99
/5R8fG/WdI/cUws7QwzRdv+XhJF4vA92qYF+smG1ZG0/Kjds6DZqp/MVU+HSBIgo
x0j57LnjSg2LlbkxGv1WsJObiX8LgpyU1tJ1rnPY4un64W5ENK0Oh7IeH8znOzEo
OvAeGWCBzEkqiupfIGula3m1VxIgPlgCS/q7H4AC1ZY7fGMGOeHLUjRjKue1XP2a
WTknhu0ZaR5W4ZrKuO4zaRduoUSGqwZyFWJ7LL26fyoClSkDQ9jcO2SxLcHLsCM7
FTiwLdUfpmC9ixf/m1/Phgw3/6PNcTfk8vV/KTnoFlvYxQl0hbzvglFCQ6d1TdVh
DQpLSE+Z/O40kkgIWYopJzI3byzXxwwwUv4iPRxKtALhIVBqu0RQ595cDGgCYTr5
ISsYnk361t1LF6kHV5SwpPpOK3rBWxrv4h40TRi/zZqqvSrJAPCRJPSWUCaRdZ97
cbpGYh9gpc1s22GTaDwHYBZEQfuoe7b2umX/K5d6nmLLWOFBusHDwcxyxAPQUq71
9khame1d+S+UKAF5H4J3+HDjxSGloYJQiZghxafWMDaVOTnACHdoMUipRiOPnNSW
ZdjfifrEPbr0VM3I9kELnxYfxuJtTQ0gkH5VzSU2jQ3xeCdsTXJTkDpiJKkTeYH0
Ss/2oeVSGFYLnD3qtVYU9fM/MNRmGE/gXwLRsyEi1XrFENJNU+bc61sg7dsU3yGz
hdSVrhiXNLYynJqkMGBn8BXYQbO5euzFE6Dls9Xu6T6p7m7fuMb30BzNjc8SgOak
hK+CRvWgB6zMYQdoWs6grFZmNoaZmajHN9eDoEvtBRBym/0IUOyZoLMygVz18O0d
4aeiJjOA4awsytxHGOPrYSDGXAq08URRAhyuxih83Jym/uH0HLQS8cqXSctjwQ7X
JWRwLMqujtauZBIVD/PD7GTX6AaInyMsaxcLdXOP6VrpStMHqkZYHfGMy31Sl/u8
84KOQezxt4M1MUumVS0AhQtfq3mtRTf7QZMNf8X+TIClJKE3cGJNiiNuyymZqGDA
oGXS4i3b7gkp6UGASgCxdv4LimAu/O2xTJTYDWjb2hBzmVp/PdzvxihrH86bGt3v
FKXNpOZlD04ieLDrcDw5yb+YLhYUeoarTe1JbW/0vrbj7IbDUKZ9x2kfzIpdKHXQ
UrxrImsrN2EVXgHw7zDl8t7UZSWOXm3eJ4GCWu4qxgQz8GLfxfnTZrJj8NMXiF/F
SL5o6wyMeE4D4AZGKPGodHoSEs/Eii5Fps5pTqhbMM5kdwVsdE3oIB1OqzjNDLoO
rcZg4QeBLfvVcH7LvCoVcP/2bOMKg2gRzQglzoAJQomdjnm8gs1uaY9nQHJvS4l8
VwIP1MDSk5AUwAnXrqlEEGCS5B4a03lO7mEv5ljtvWNswJPXb1GzsGlqU951a+7a
xa9Gzt1JOyYUWymplwOq4XY/7Qx27QJawsde4vSTMxwGp+DwwCnDalpnhZUYJGS3
Pw/t33bf+r/DxBMxA+lbE3rDUhuWE1+7w4x4aBzw15EaM+SXeb6sBgdLNs7+SC8F
ff17HMFskqvoPHM2IKG3ef4knPKnjSTslQCc4Z6oxkfpZYhG2Zq3M1DfYN6hUFFH
D1CSthK5KDJugsYVV07PAdYw2wu2eKQjizI4hLkm76Zr6m8M/XBZahQNwAez7GnC
G1SBJsN40l4Z9rHzHWlv4/4B9/T1pWzg5JpwcheCxLq6lHdclRWdYC25jYRXK+3r
jPne3z16dPO8JDtErO/98S0FnytqLTD9GKYYqsnTt6y9pFCvikplQWoe3SH4KoIv
wcqV9YtZz0jjruZTx5CwuZ4F1/SDNSBZiySiKARvzOXlQlk5X9ALxDq9KGxtHBx+
WIrmyFfTGZqFEW1eZCTCPuRSVcLj9FzePLgSknh+MDeDO+FgQH8YthX+QLipuX0c
OVnbgDICtemEJwqMukcVfoqkG2og4fZmOdbW1nW6E7PdDbH86KKngGtemg44rNq4
56EAoTdcqnRhUJCRvnwi6TKydF4BoofbzmVDAPAvabJOwOfNfoz7IzTBZI5rfv0V
70+R0qQCNt7WBaeRDBVdHvCFFTLyNt99lkwWmc3D56YCdfgrUOFsMIOKSda3P18n
VCTqpBVIUanyAFu0fVXKLcpvCLis9dTNYU7i9RLeyhemm6Gq7SJGXN5C+ug2YVKn
JCS5iuTGpgrQK6ZCGSCJAS5Y5+Rro3U4f2s5RnmmwzxS9jHXeUGJ904V2pNk0wIz
kh/XhhkPEfGR8RX70qAvGfqCbG/Rr/+53ag0EeHAqJo6j8ZTO/pMxLJKDbkBYApq
ZhBwmLeYvJxtfLBuAb90NN3SVgnXo+zH+WnuSpWxwgD97L20M1H3Sbd1ETCfq/r0
8ZyFeHPbJqykKelA2KjcYoJ79/M75XJMVSDOyqNnPnObX2kEVtl2zeemIgnxkqag
WceU3RgThfLevhq1BvAUvn5L+DRPdFcsGdumC7poARiuyF9lLowJs9A+WK3AOMIO
FZsB16XQtKYAxQXfYotSqm/phqI1mERQ+tUh/UvYD0I1hPUm9gftI8zOUIt96viK
Wx9Z5xR2zp8MiDfYKgwlHPsneHCrJ2YD0GF7cwhgpKcrP78ovLANWapRzWySYnbA
aLWf2RLAXsvzM2DSvlJnCOey4Y9h1DWAuD9NmW5x+XYjqis/Dx5J5YrW32S/WpU2
ZsKpTroirzSMSIhhsGUGWSdIOvJB6b0c3XfFWCe1uQfOR5bFxSxQ+T2vc9rc1eIJ
Imm761Nyv6y7tSzWPkYx+9ePo5Y9XGN6Pgl+4MzeX7D70QVtwuYGxgcuX3Z7VLa5
twe6tswwYvsPICcU/Zjzhb/DxLnNKIptz7emiuFpP5NlUDG93MODBKuai8LlijNL
OpfvdpPzYvF+b/whF6CkfC/0eUF2rbw6gchmgUm5RXRvu4QYcjnrU2K8iSsEFp8G
7tT5snURZ+ljg/6BJG/sc3BPt5juW2Dl49EogYZTsUedvwL9Uki9tD/Nzh9bCgsi
UvWOAd0N6V1yb2N74uOYslVDgteHlgUj3+3+TktrU4uQJPrbbxv1D7Xul6nvid1R
xnQUeOd3Xve2XMg7PPs5zeRPhRUvp10PaJLKqpKJ+kb9solKHXlr7qhBI6Mgn9UQ
zGJxz6piYfchTncC+AXgQqh17S4d0AJzBIqHY5DjTKTinY3VwOMyp2qWRYJvI4Tv
y5iKAo3F1DrwoKgSLpH3nbyColmXS90foH1OYeE9GsrXAOQDoJCPB+emyQWcuPn3
NrHOiQgEuC/mS4GGruRZHavFgiGEr+31WaIhHukGP8cJbcnRb+nUtZD6mfAdmaze
CulmhZJU9rPuOyvfsvrdTQ/jhBqVsUDIt3Sbco9eBEYDy/lrTx5cUBjxv16W8op1
PCFs9R8cP7Npi/3x6nfIVqK05ALR5kL1/Xqm2zZ50QoVOgd3jLVcJJEDg7UH6NZH
VLQevSQfbn0MXsq3k5RK3ebjPDtTf58T+/UnrT8AffSGbMA0Tt/07gK+gH+i8qbf
GgJ40yYcGgllIpo2g/EdERk6V8J+FAojuzWFdecj+69Y9JpxNEUi6gOnYmSZykXz
if4Pjc18hSP6Mlc0wKBOm/4L4BC4zzIjC5sXP+CGFySvQmKAQcpu4XWYksd7Y9yZ
rTi8LHE0N/qz3BwKLEwoonqiaeA1i91YRJXkgArhorDroAfuEx6g08kPcK0eWw9Y
7c5Q/HQdi24LZxyoqAbW84bIQ1yNiETzijXdlTJCmGuRdIRRzeP+6jyCm7vyx9hv
Ub31cOWsJqewijr7rnr9wkqQ6p8iyaFP2w5zZdKbPsPd7mm9qYxqciAXu3ciOVIv
z5PhmYC8Wic+xDxyRHHLrykPvpTjd0pk41BwA7G2Lt1ZQhX83mVUsfbZPCCWiIUu
2TqDS4eJypvqTPtbLlPcZzUuXrWNM4qyKUll8gNuG062OL4vbQj797RXZak5pVZl
AVAJbSBCkpg4/eOjcHTIXTXb/ejorshIVqUZa1Vii2xOWrM1HPBYY1mReRHn6dKD
bg1xWGUPIb05XBhMRzFlefF1vM+Ijn20y8DkZ5xd5aJAB2FFP96YEbXugVN4PRNk
QqHlz6Q+AvUMgCxYjr8dRFLdLVi63sTbM6WXSs6iLb0UaEqOFhPnx69DyMi1IlAt
2D2sURqhGu3hwdLeMtjA43HB1d9zFRr4KFBR+sK8uBMCCmINB1mCF+6k2zgtrz8i
vEwL3p3SNYMnkEDRxawvrQHdsRYBynWTEj3cIm6yVk+sB5dkGf3+wAPonUpcKHRm
Wgs9yCu9G3H4WZRupio0dkmthkDuize01gVgta2Y3iobHLY7TSNmfve6NL1usjzH
KOeEtaz0tnkED8mVUftivrcWevAmdB9T12YZhdxyfpJy3WaIva9wp2pSkrbv+cd8
zX9OfrWriT9ktj2gkYUHCqEEk666I90NeSnGkXEd4qoKmcK1FxkC41u6DThGPEWq
C+71+d3D03FjOngJCx91WhonObpQV2lhGv5seRR+jBm3s16ZIdjexpyEMICozd1O
kWPsB4qdQG7Cjkz/J5502PtKa+8S2M/KcSayzG1cDTxfILlGnZY6bMsLTgrNAzNJ
wu+m9cyj+1TD8ztp378H5vlfV1Mr9plkzYJ2tRFDLrHeHY/JE/eJRhBKLfTxlCd1
oGUtGM5LjFko3RmoMPragvKx7u3gC8MKP6y7fuOJmIzCpu9oyBqDjbzmKPadZiBY
89X+56YUZlxjv76ThJXO2vsNro6ZUmDkADUUVoLn0HPmj1mmlSLSB2Q70y1PyPJq
i88yCbsN1YLVriqia3kFuPNdmq7+9hMLJvuoL0uHUtKvVbSZaelVsqTiPMxI+eBV
WCp6/5MCh23CZJtK2THKNKF6OY28bs1wX9yJ8oDdQ0xQDuTfm8lA9AI2qOnJy/G0
fTmlNHLYnf0nBwM885e8oIgEvLJhTPXL+ZgzXbyf4OlQgv0htIHKTIrBDYLekZ60
iXGSjoYlJk8IMWm/4uqcSkowVmLSClxiaV0PRnXK2gUeItWpkYkNkyipZ7/4gVPy
b7IGzvcVNa5yiPAzg1UPFH/BsAkRxlgejC0qqtavAkmlE6xk4JAysWFAyBmXyeyI
rHrcNdwpfmoNYvtBkI9h7GcKZgF+5KzzZbkKK/H5ARJWgsfSpGGq3ffBmUeVcct7
42huRRhtktl2GNbT7cTvC4KS2xSQpHOWCdmk6A80SNnrk04OYO+lLh2K6/89MkFr
TUnTWVWMBj7jnDmesJ/d1nMmIykEuXIljd0Tc7i7bZwc+rBscbE0bsU9aSVT5X1t
UUwdLRYYd3k+HIw6VujdEoHOQEXp2sv9kPVy5nAMDoyFGC0iz9awn2+2NbhdwGZK
yfOmoGXod5cKnKSPTRPsJiwwP7gRcuHOZj2pItFGDYnXRGObJk2TXvATaJ8GyUTT
GY6uTnqcLfhGrftEX4KLUr77FIQnxBe1DSAbt4DjyrMBX9HzLr+ahDlmRqBk7yhe
WIAD/duKWWC9r28y7ZdcSjgI2LTwoqhXjZrLt9NDH8jpQ8h4XBgqweQywwNYiSsi
sv0X82EDo7k/PEJlCDQ8aRJDsBeUZTHwwQH0HZNBD1zCYO0+datmJXViEv+e1pTP
km+2aKdZVC3BVOQwwIRWfxSQlnj2FLyw7+IExFDUJ823OyW2XfYcFjPvdzBTXLBh
MrPBkbrfGuhyvRG5BW0rqbXoP1tkHrOrnNfOaMZHARzqPy2+4WVrCgZ6Fkb4M3p1
RApm/L3umw3+OLlm+/uFUhHQ742K4O+3IgedBvEAYY0TTGbt0fSrqplUCHVrHCvS
c7PgrgXTOH4UFtLsycTysiWjq18eNeSxQIo7dYeHY7rUyzbUc/FfddKtX7EdZcKS
O51vac0hw2Syh3lGNCBzMhUcEJfPrWigF+44s77mRJP1r4EgfYOFlA++Jvl/QdlM
SqkPsko3DPdMMncZwaMW7es7GZTrSnhyoc0Mvc0Z+su+uOIGkBUxkIH1ijLhNqx3
8Dh6zvy2jTB5SMDzfSEYEGssVorz8wH8CbKJXKqzXVUjJFhDyGCjRwQ5q+SeU0AQ
aIwSVjiIv5gvD3BReuFFCrFJOo3atJIjn+PLgFdts4mV1q6q5EbVMcOw/0U0Ryxa
g547eDdmFcxcrNlvJg3o5lRo2wm2LeEBoqAtvrvC4xHXj7z6paZJI/hwcfJ+XiRA
FaN3W6SsI56+4dIx68RHZPSOiYINUBG4BRZyoqj2ZhCGsrH5VftqCGgSKQ4xTJlw
LHe0p6R/wCqN7tTZgKdfYtIu0JSQCbbCIMjNK4IH3VeiNiQAj29H3iCveaEkQhBL
ZJcKm+eIvsjFLAZ+m5J+Ak7bqD++u3DVBW4RQEYcAnpkcfIUJHPag5Yicu8G4RHa
SVw/YJrU6aUieAo7iYy3vQoNlSAvuJd1Ccu0YsUhWNdsyipPzojQZvxGJvDtWLUW
iNakqkaA07smWiEUHdN+G1J+C8V+gmo6csQuB48mczNDJ+hlS/6YHcSTsra8hser
r+N4CTQPzRajNFxhM47+Nu0xqis9vKZ125pfcIvUE+dAUhBuBF9reWeXLaOLoT2k
R1lMbFGE4FZYHRYMH2qMsWtVlamKefZfsDOVigyWOZ2B3OvnOIwWG5wwbbmVTNt/
6pbqNfsVD8P+diLpTsT62zYLdvldIUKa0sGO1/yUYI1g7/Sab6IQeCV4peaboFV0
w6W34J8vDUvyzHQcE9xm/bJ1L2CQGt0i4PHDF7XjmLhmld7TY8CkCzmbozqZjLWB
E8xjcWZlGgy5RMICCMtm4iRj3cPq+HqPAyUwyZscUxfPXqiVCgm1+la+/Wi3Bsml
DIPX6Kiwcof69DX4Vj3tzIYwoYkjjcAAG05RdsSJsF9RXMSb+VVbNsu9tdQjZThY
wTJkY980S/zHdNvRI+UKr4L+/RiebVFsmZsVK0FoL3atR4nP81rb03u1fLzX5eTX
oxlABiUmDPaETaxcGX4G6OWwfBdh02cwBfPl9OiCn3W89rX6l3ZZDGTfKtx+z7Cj
4wGk69pnipKxCiGGabxNhUpz5MQt2X+ApkUeTeKxnZV6VF1hSiZ24cWByaLvoNmB
CLMzJuruy2SK1bG4PY/iefFm0uSh/ldomgszN1MkZEJxDhCTnTNbRsEFIvWglX8/
Fys0wvJ7vYUdZx+SLXtVxyLPBu3EjMxneFfViH1ltheF6FaIx10jmb9P1i3uhudj
BB8qJeWe1Hc7tzXzeRKBGFGlsZS4BYM/57CYIvYLFuZblgYajOi9JlLsqLu1S7Xm
s5l1/DMkCFClTc/DyvUpzYY228pc8xX6uoAk6p8pBBmqWyjmMrPtSxibARHC8I2x
xDqIr9uvLJdvNjbHRuCkXvh9mozd0rBDd346y0LDcREJk1qY51z+Sof34g7mAMQ4
WYlRjH1cO7olxQOT6sRD4iBCJ7ckeJBCI1YkIx0q0DKPWS+O0w8BBZwsx2WNCa5K
ieT2ThxN13dCsOmJfUrzgiDI+SWuVVT0Qy0YXJKsPj86NUPo81xF2vY/VbrG8qjT
07mIARuqgPl9RcKhwchq6CwkezMXurt7d3vRqqmJHotl+Mycfs/+o03GLsnyLfyG
oIy8w6QcBGisdw/g+0heSi9Hr75BnCKZGAmV/KuSPUyTp38JkD7V46M8Q2gTySDr
9/9hm/hEo5qERZtlk/37ArggyHRhumayVm5oLfKY49Y4FKpNKExHDwBYqKi0nShk
d1SV+XMe7uWuJCBVYx3x08Rwgce+aax0/OLXeBg/lvEuVIvPLeh05rCL/WAjdZTi
6OUtWZkM14oRLK9UVOKIDIbVGSTNeq8ixR9vNSydk3Dkzt8QpjMLFFh6x7CM+Hjt
6zs3uVl0+rzrQixqi1SPY2SzyZudUFP4omz4pOntf7WgYs14JHJx2SL0DA9ySAkf
2xqcjqQHvvhR5OqLVAUTi3EiYLlFYMMaE50SaSsyx/Wa3YbbclfIRp48lqikK8ts
pK+q0EhzspYXNYDI2FgPg8vxMdZk8bUMMAGlJKC8sVusFAx21Bn51oivdRFwl8Nj
dg4vfkBE804VvpNP/8br9Mcda9BGa0gXhG2+1xBWsUYYtR1BOny9XhKta90haeOR
nEv0tLVpqawLG4aUTo5qT3MDSSxIpRn1yzZJgFHhg7HER4ZzcnvZLAqmZvjkE342
7UX9faOHsg5iiI6OrAXC8QHHeevCDXsNNZONpY2phi41l3h32k+XcJRIOY91Z1/p
T21cZMYDWYPw94wpYarckesw8M6+jtMDdhSmpiz545g6lcKhIA0elZTpZU1E6PLx
jJJAGeBjLReTF7AqSxFuEUAwCZCW9EuBIbtGVW1iWi68wpeo2MrTRV/fmnxzKm06
4vSLAmyBp6ibVaosTrizMD3UsluTQYbSKdCHcsX4bZi5xUkl7HAUzxAjYOgTx0YA
wbMkxPMRdNSsBPlNE8Vtv0zlR3Kyyt8gUXCVgOy74k8Ff5rEkLelqHxmL/fJmiJm
tKT6cdtbLA9gf6rjg7fQvKyeO1MWc4v9yuH/L/xHxUa+SiAYVruu5/wP0vXkuETM
gCRo8Zs8II4MWr826xI7Z5cgtucqC0KVKOqzjfw4xoUbikErYMVQknPK6CU/21o7
5R0XCxe5yI4ersg7kkeE2tp6AmS3bYUGymEL2LndcbMMulWEoIUEQcHKY6p5VFz1
4A9aWy/IYu7ScRpjQaIXGxUVShoyrGzejqp2pllF6fpyTfChwxnlkFABWjWcOfI0
IaQc9f8qkyifZJe3DX6VoOlBJGTKRGatEVhIh6NnggC5BKscOOBFUGn9YHLZObEg
zlu7rUB4EFT+Hmx7tMpRIsLG7S7nPltgQQRlPSYx5JOd27pfENIlv37R2VLphLeK
wamKD6bQjy11hwRlYukFdisFHouhHbUbAJrUzN+3TWykm5DHL/fvAXnVsOFMTHOM
cHQEhCdDZTAhVCZB69l41DhkZjP8P/by2p8Ib/Ud+kA12e/FP1tX5zr3f7k9qKl7
UuBFn/KODZGXcSDMwVJcAri+iBdqyhljCbWnzDcYmS0gXFBONfYQz0lj/vX9BKfv
dZ4CkxgRl6KrndANFwymUWKu4G6Di46MLWOzGpSNuYXtry6yGTFTSOtV1TIXEGH9
1BFusOpfhqgtpkvzOXvuPOLKDHalRVqqHQQyA087bpEXLj9hicatM2Whl4uMSAwW
IJ8mt6QRQyc9t73nVLqCLrByZX5Sq6jH3+U8LYHGf7UiiVh11h0EC3ii+oPB6JG0
pQxAbJyDo+Gnc+sjE3CiAKFj3VpuEhrTw0ULQdwN91xfMcUckXLPj9nlhVjk5IgJ
DvnkLnRTc0oaykBxXbZ6RIL0NsOst8GCJ2S2pZXd/cENGb5KCYYl0h7nQrg2npPV
gf7ooZ+UjbPJokltAJUjYnU/CCH/rlSKR/nwOGtsAASetfnGPEm5JuMPs6n0GRfE
eBe/TUlkj+Ezz/e92Zq8m2PGhzCVhu9fErOer0s1pMUVzz0OjmzYWa1R9PusCulc
xJztCMoyIbbYkcfmAL8H+qVPi/3Nmu0U4HpB3DV2tZqKqMLlzc4nzSF4CNAVOjRU
++6MMgHOK7v8F2mCzZU7btZ82g6EZA0OU/K0FZCk2btFFXlatQPMNO4J8AwQvKbr
LWyoaFWUynF7aXmtTVHx3128Csm2w8yAbg1hVUL48t7CbbClX988I70UBhmchbhJ
wiUq4RrC+r/IYdIQUwCFWfU3OMkE9qTr04rgGeZM5yyLN8twvVVSJx2ks2ijYlGF
FZvEUVDR8kT3RQcYGb9TYi5DavqHkms5v/2JuOYsl1MjILbLVXAncxve79BClMO/
x49qj24LTk1WwJzdj8TdrRT6ZplCVtWUnYeahWhjE/ieeapZgL9BM/ZdELu+q3b6
RTFe4WHfzKhOWznGOz0S/aLJBz+ubLZ2PUc6+2/X+h20x4r7SL2UfLOaTTKt2etS
45WdhYu3ZsKGZadL3ugrj4l6KDA4jJoQh9kYrRgqn87mWgTmXkB9/dIiNVV6gj7A
cjMdSneITmW/aB4PrjFpISmNDfDkRkOrHCKRaLTqIr62kLiWiumIRyKhaKTR93fP
3udIpiyasXTea5RdegnHgylbAYUSSmEux+tKIPrIlFpLFnrAdr/ZF9iB5j6w0HiP
aRk8Mo/PxW1PHd/UhVbTUd+jLS0Uonq9lyLtTINtRD0PqyCiLCW2VXhzt6awRaaY
rhQbsjAfHFFNj8pUUTD74mDDpB0P1ZHfE3EIn6Kg3DolS9swqicLL6QKHYtywIY/
tHG7U66sVWn634NvUcuFLtn4veW05bKMibAFc3xzdEIuqM9gZnsH0fa4Qu/AaRtx
O1pEn0MCNHuhBa9vVY2/cTR4D0dN7yIm5OofdqNe7TO0JmlNaMv2l/k4ZSuWU+SA
byTAepUSdcA6dkpQsoqdayrvXbmX6yHBRwkuRgpTkROjUwneQAg4ebBuoFqW1iU3
3Q4v+pp4ALtNwIE9yJgW8cJrYKqqgkE9YJrZn5cLZTL+G7tMxlt++aoBYcmhFOdZ
OXj/gXSa3KPBIpAthICMkdRrA7g0SQCzJsoQYMD0uWCcfIVNUC5dOqOZGistRRJS
2t55lStWVlXfQJrYaLXFmlANBsuLnFJiAMtrlytaDMCEntcP1MfxHNFlqVsBjtJZ
qnn0oww+mLBdEdVdFAP2ISWOkb7Ur93rcTS5Ldj2ETp70Zg6TAocZY7yuQYHt2/g
kjBlhR5Drg9GzUfMSBqy0f/U4uoerxrhBgUsq3i2ynG+f0YNV93bjgnHfPXlQA7v
AtUMj+z5lyf95O5BxfkK1RIPNvVU/wXY+LkmKkNFw9GG/agYeI7bPrvBFyHc9YAH
431n9GUI8v/IYN9CRCGDFm4/HIGT6X4oWR/+uiwqS1KSVl5jA+t2sY1mHj0HpX9o
+g0JX4Dq21FG9P526SgvKGALS71hMANUcN7OtgsRuGrm/smzOnPDttE3Z5ai6IUl
hMJcnoIJ1OQrzErUAqb4lCX48aAvNyEixvBPMhGx62hxxBL2bTixBNKtEyQj2Ile
JaRSpp4oHTH6OWmSUAtGTS3FL8F4B8Q923gaaAfYP0wlBpFoOcWJUzYhexMmUwPL
fTRpeAzFZPQ39MS7xzMasjngq/iPYJ+n4rT/J+DYqOKlM/gKyR2h4iXIVdw8Z1rm
I1gAqs+Tiq4/dimN9z7cODWYvdsG+4PRo+Jpzzm3Md+fiBXsl1HliasONQO/9h6n
e17NMYJ6xDAfMrzpREiZ2MA/4SMS8aT6oVyf4VREC1xZsuyOBmiOthimcC3lstZ5
l3ZexFulh6GrXITCCPFSyTlEyoBsT6iJsZDJND+tv1E4iHV9gMGO/xeKtQw0kQE4
uGhi2jDuGCIHHJ+i1DQF8TOQyG64hRbZ3kMyGfxiQHO4xHjLlfxopObxUvCbbM5w
L4DqHgn1Fuclcn9GYkyuj2nBpTwbv05eHC2ATiL6J9rKxHcIEgb7KljpzHy7hSpx
3DzB78wHC0VCVsK1SOkKSbDtz1+3ZsIgIdPzi0AtDIP7VcL6qB+plQ/zrv6x3Ggo
dgemspGVSUGUebhzO/WPtFfXjwfiXma9AuEnBSi/pQ3TXeuXmhskBTW22Wv9d8L/
QsG1m918aXbqJtvPgMOeTm9bRDYD91V4SJgoNmUC9NykQb6JGYbuLWDCicIp2uP3
BXltChNmIZBPQpGRfJhwel5RZ69WdEZCIyan0jWZ3pjOAPTZ0wy3DzHvPP0wUsXm
QVcVNhZXbAV6sknMEx3K/vSu6do6MqBfQKs+OZF+lkgtofiVgtgwF5J5/8eFWPZv
Uszxf/G7aU/ofbNkzYWI6iUKE4Sz1ayCGxKf7KjhpuW7pffleRTNmyAvJ8jWggp8
Tmb5zna2r0RLgdev7O/pF3Y3coibpREA7ZbYsdHatFh+/0MW2qrl5zuciYm5JlKt
etM7EKYNGY4zk0HFuhPI+lll7/4wwSNl2E1PdR6cNv5kyD+eMCdmGcq9jA04GxLO
n1f2lpZ8FRdIYvInlRz49Coup/AqCycPFruri+7jEXkz50HxYufcH1Zt4d9N4JmI
hzn2jGbaMiduokwyupCMsDlIwbFGM6pawrQTHIKyJ/1yX5mKdzI1kJ1I904eMtKI
VI8tWg4LyGmV4dyhWFQsXDamizuDStvaBgloDOYPi91W7+I69BcJsZntdrRvUo2w
eORAGjRK0hPgcE2jv2FnUY/U+Bf2i9ZKyaGa63n75+arxzIJZx84IanZqAdMlqbT
S6hY0RmyjM7khCNPGTMGkvZHHIgtiRtCCjYCMn5qeHlFJ1aZQYz0WTwluNGcXCk6
IvJf2YdKnkw7PMelX590sSVrJ4eHyocVnZTmB1izT/qALIuR4IEcCV1n8xWVw5n7
dooBdHP1uBJv69Kf3ys8ZJTm/LACPoU4CRdQkScGwazrtWZF2AaWn0RkG/WSRUz7
/3HmrjKhaUqgcpFDP2ctYRTLKtRgx9h1mTbXI11vCDm4BpclqLe0BXg8THcdAbz3
7p7l7/BEnFE46nKSxKpcelG3Y0BRES4z87Oat82ukjoKr247TbvjtTgLWr7jIbdY
gO5UXEKCwN9vfjmHBrlYOySZe0aJlSyaxOTfkSRBJXLG+R2GVTx1CVZJfahcu4bS
GVUeWwzt3kZ6Adjyu3kijiDbAxfPCeyRa5a1Kn6ri4v1V/Js3qUIcQTWYEMPiMf6
Km3c46U4yQbcCnq4pCrN/06YhskalIfQretRSF3p1ExsL6AWRlxYv+w3YW08PA62
O1gFOvGwjQtcsQ+Tc2fyzorEOS4tHnqt0elfJjIEZ6GLvqcmzAhyQ0Yu3D2HIc7J
++PdLk6mmNsT9IyNqsMW1/j/UonB12jksVNW8YJmW99Ld2HP2+IEuhT1L6BxfoGK
3hdp448pTnW+up1jZ5wgUeKgvXAB3HMgX8GGJX5spMluG/wBGs9uU49fA5IEz/66
o1CwLyixUf58tuJGbaprcBeb4Ozs1buCRxy/N2ZAclO1tZLieOdm0mQuRBmi35Yp
qzwmFiJAWcPL3/7cGNaWe53LQW6Lg5TuCLGdueoB6fxiqDvP7MdscU6oxyJFqlQD
+cKkq7EEReO54EtrD/5UDD8A/YOxFVLoHER2FPB1LprONE+J3tYKbvt5GWSgqB1d
A5PLsSgeZHYpjH1cSqAbPyYQbbVb8ENflQVRLJb3Y4nScdWmaxrMYwbJTQXoChfb
eBAaoB24xDICoSbVnq7I1qFjbThClG4FOel6qkJDkeMSuU3YXIcu9e2Zaq2NxLLs
kNaRiOrQ0xm0g7zCHIUfeBnW6jDmg/dIK1tJKj2nZhb7N4l0/H7k+OJxmJAIIr9X
JnFRPlb8WNiR9n/Pzl1VviPPpWYG5hHV4VqudoZmQBAeM/e3+dvUE3gwYWlm9MXX
3Q8YwR7UySf/vdWMRM92HjSfDfRYsMFyfx4ZA1YCX3M2z/GVywvGQIlsX9cS/UkR
d9HUAZqWGqP/HrmpWstJY/JndYuy9nt66wo5UWRz8TQRvbzVkwyeBDXD76l1xOUp
LmpU+LKQPp8w9Xlnbm1WzS5ZP5jNn7bUfyfGVtL49/L2vNHCzuit/yj9K5tRNWNK
rue4QHYmsqDanOCYje0ryVTeqW5YzOl4f4LhSxm7TIelmsrPEn3RHVwoxz+6AYXO
EGzO2QcXkPaPS5IQ13U/rc+1/cjt0o5Cxday77yvhTAzno/I6dfZbbEkxCSlFs72
WLQy0TW9MhXO73oT6TBrr2AyX9kmYf0n1yKnM3qOzY9KwLKlKqczCk1HdyEu6bZ7
y9gF2NybHrpy5NRXA1Ew3mBFCgbQKTSffBxfictQpI8ra+NQlGZ5XDDuWAzWQtP5
st5fkp/ZI0QIk9vNMlhBrU1Gsko3SwWVB+EONMYJYKw0DJQ2p9LJgu/XiafWOftm
QlK11u2g/sxOg2FfwmZ6cNErsT29kZ9DMiprTcS2YDyJTEZT6oliWO1OV8kfhnOZ
5Xq8X056lEO2tP3YPBdXUNj2VOJu8fKPBOizJnEIK3AfAbZbhVNC07oyEihB9j0D
my3WvJAXExR1AG3Nav90d87e2LNMDDb2ebjtMyjAPQOIN9tZoKkO04+tDhVOqlFL
ZyDudFv0Cz5ZILHj77onJW0K+A5hW1I2/sslW7zwWd7AH/PdoJIakZW4r2CPkpKm
yFNGm75gMHTGi+SbT66VZHc+I82D7/bf+U1QqXDnMtJhtneOMiJvo89oiTx8DAW9
shjHkM6zV6kf90xq+miLFFZ+jvaYpA/qHF8vxzrtutUaQOC3N9BCJXPdXxRonpBK
Ti3Md9JPjxujfOGuiUz3GA4ZRMvgRI/WNWD0G3Nu3dhZj26dURBYGKRDgq0XWPM+
i7gPr5wju/lB37ibcLb3Ez5hUQLAv6bYcJfE6FwcMoQpXylzdX76qSu/+BZWcpea
kqXuErQAEgtVzTt2cDunC9fuM+j8CnpvM+C3tupP/xcDMjILHPXjGmVsB7MbAz2M
jZ8JzADiDd/+M/V5ZjPplJDs1kVFk3TJaK3kXwfqwJ7ljh40daOkK1p+uiuGVFZr
NSoBwX3Qy005ChbkXRtdHWDdWAQZ9qQItA1Nk/vZTYHRYHBWYhlMHNmGU2av7wwi
hF2Qm/1EEaUnbXL3EcqxXdhBZnaqAK99zfYIrKhuRj6JTrfJgjN7lzJeRk80MKXX
Hf4NnmkPud2QolVYtM3b1q8mubJjyEg9KGPi85i+H7m4DZ0ZKvo8wkzx9s0/IT90
AsukvEQuAD/liIKRbCkQuoazmUPZYZfC0lWN23bvG0vbZwguuXUmfp0zYlHZPq/G
f0z6t9UL6pdiG9GRH3Ef1feZTTRxJZ28E40YEcboVjGMRHLCf1M2uYV6A+GFrAoe
CX2vzRSJyWvzU4sCp3baMSjy6EE9FEp3nEfbP78+qR4cRWPGpLKKEqP6WP8G/dzF
cNhZguhydNi2B01XL5fbAsoZ7mQgF+AALE6HVFD8p7YQgRnOFp0+j7e54fOaGpZx
hMODKNFnoXnbaFqk1+wMg67HKjKiUBjqAKn7+F2Rbt1r/YBxkyMvQNb2pnXnO2Gr
Ai8iVYmo2OBsrtcRVPP+a58caYRwv8euE0iYkXBPVW9Gw3VGQiI/dLEBFyFoEh7Z
RCYpx29Nj0REbShPDi5S3Zkc6f2WqIgx4vEPCzd2vzrT8hxuUIXk0OavkZw9oQXf
BXN72bNToi8n53pjP9vvUOqy6hRGVQcu/e9R3wzPfGpqCeTMyLSkevmjKAKZkKEp
GNtRWmtQx2n9/lpqvRlTgzMsmZkgXJIHwDr09fzNU0E7O/906a7eP6CDY9d4xx5K
wG192wP57T7ImIywAheGC92vBgZtC4ZWimDRCpczNXm51DitK4EhGwDjQHN0iiJ7
26CuZRZyikVEOrVB1J1rVaZauFJQ2pMpV974boAA3o2QAnZ44YCEkPp9W7UxVy7L
bQ7fa6CU40K9o+0UGk9PfM4RL7crPAV69/GPUOJhIH8FTjyZtPCMquIdTi1AgAPf
STXZ5D5ypxSPm5VrcsgAFSa7g6CJbLtqoTdNabwaqV/QUXauoKb5aoQzKCVCgnY8
VbHRHNi+rj2ZCrHHGHK53LZ5wUnzazRdTvdz6ozGXmpsqWeQ5KlD/AiywS58JeNT
A1QYWQW9kczBOdY5IK2PKTwhJbWS8aZ8aFE2OkPRP5Jrk2FaqYqFOSUkTrs0HXU9
hAkINLX4CfysO5MQ9xn0P8Nnaakdo60AUk2TW2aqYf8umslvtGSRt4+9h0nIfhbf
rBRqoBTZ+XatYlV8QL/ZE+8POR+bRc6+ZsCuIz0QwJ9fKURoroJNFl90MwFuHqVI
A8AvFLpmCqqxdl1E9WMlxOAGuEhYYE5LhOT5E3EB4hPq7JCXMuptTeKLagWJNKez
qgIdmrGCBgEtLOY/jZi2sTHCLpPH9Ai3QWHFIRDX2OTT6QgrpNX0UCTyuCjICfT0
JeM0uCprW3drC4kkETCC/hdRjLG4jnq9InyMuKXuG1fxTz3jCN+MblaFcYg3866q
D/JNXABjh/cHCX40BcPMrk41DL++/L7eWEjuECTq1PsZpKMZn+aDcVsjFhGnME4J
v/XalPBm16/SVII14Gx9Ojou4grH1QhcvkeXjOfc4j1OjPCCBZcRkErSJ+F9Pq77
9tvj5IdzJnYvli634D8nirLE97dq7UzwE2xqRRLvgAANlWOCGTzyyvP3ncuaW/nO
Jo6Tx9GwzRs05yPYpcLiTAUGyJ+1ucP3oMv/k/6g/v7nEARcQkH93Y049QznvWY0
2GpZonID7haRRCmDHNqUCpZ/WtnCcZ+2NyuwlwCDiq5YSZrK2ixvOLZDhno6IQPv
qTVYrzrKfcbgqQB6LmJUkhV2wd2cXyAWDtXxCid8mu//nBSsy18vUZnrslR9SeqM
QZ9kchpgo2RzZeGHogVNcZiWsjENxbwe4yxe4hXLv9fLxxpVCBNCGsJObk69qH64
Rn56glEy1p9M9jOUYtin7QsH4AwnRwTaQ6f9DFW+QLy/csEALLJOOT+pR9LwFcPH
kEWo+yeq0/40CD5ZmWGGiRGUKo7mJoTJ61bE6fTMiaXGLdRnrajABI+O2qcwsxdF
SqwVfLFRSnF4ZWb3ayb9RL+TTJ3kjD/6cQi4jtNjCy306GWMwhiivB2rDW8OeKTc
7MpLnQ3EkeR8PcD6N2d42BUdNLKCdcjcgL5VUPc+Z3XLeqT/vRLnT41KVu+wz9eD
9/69BJb/1Q8OssBaSOF0aJBSxE8Zqjpcp87qkc9rlAEMXNQqqCfI7Czb66LClWWF
aYYB5coeZgL3uzaP9EgQAqlYdcv35T4XOQ6g7eXKkPgfu07+TWxf3FN5EAVBKZuQ
tVVh+ky7LdIIFHU06CtaiTzgDFPPQgbzJnRsiZU4h1TAZ2WHzfBd0VH8YJ5Pt0DQ
JIypffpoT/6w9LTJNBBdekwcU2kLNIJhNyg7TqBdRPHQHS1eBJiLOG8r5kCN6kuU
hV1zg7rE7xDhDGpR/MZGAZn7K9J583QBW128xvk4ytbwf2GPPswv69KfBvRO/84j
n4oTasoveuIfX09HQHGnQyr+MPP3YH4WqgtV/ocpbp8cKt1PF4eYaoLILNltM4gy
0kWsDC1aZOGYl8rSUpZeDuSf+IdT48hWVlLbeL6a6JI9cRrUJe9XsbODdErFVJ/f
yXNxDUI2FXaJnlzv38LADgdQkdkEdSvPGxRh6YJPnwEOt2kMP5jGz8Qr6hCyUcsw
kOOtfuZmRh7h+E1YB85+Wc/VBXqpFXHvUsRLSqJyD/NDrcCotNl7Puexqj0RG8Gu
kk6zHzWcxzQkcEjDqCraYwE3wQPoQjfNnOlyECA/65CZRqhil//gGRKM+3J8khaq
IWdqgyKgMGXOmgbPE6eF395yxzPDZqUQ+QxVGD0l+M1LcAz8csntGgVjp4szIev6
5JdtVEbtKohwxwi+qdF23UntINS1ZnOw37pnsU29/jO4yuIG7kIS8kCQvhlvbUux
xMSgRbqZFDqksVGlui7yV38EShemYh8pP2OGlFGSdKCPhUNEPdEnezklBMQwcv32
5eAycnZ9Me4u6Tc1zrtf8Ufhniyi4cvCZtrPiWnvfr8DarzTqGNH8yD3HuWvTUz5
qQfGP2DqVIq9OrnK5eepSTLLeJOnY/rGR8a+g0ApEEJm5XEfCSabOfETeFx3daQu
vUV6P2lsG+G6FAvYRGLiVFQDRQBlvW62JReHd7zVOLmmQd1nj0VIpHnfzGHXhJcl
4jcaD4KdKPZQP/8mwDDOGlNPWBh5bGHS6O3HVnYAUBKBQCg/Khv3TS4xQxS+tEdB
SSyW7AqZ0ATaEcwY7QqgrZOr6IK3tBHjtKnYG1tKK4vSsXLCauedDBAOO5cL/exH
CDxMQUaW0eqIwZedL7+0s99OjddrfgUvMtxRN5qEds68s6IiEt2f3gz99Uwz+H2h
92pp7KexLl8VgOMH+8VlkMcBJcpzuTseXqULd23zQXCBKFUbEVyKLApC0lx/T9YR
S+yyTgth2FqipGBksVzt9io9bCd72JSdOmbUoN2vgcTNXEm/28vvskM3s07OFZHV
lbiJS/c0kStNMrJ6vOY/qdoEA2fvgk16+zwECN/oXzZzIHOArBjfUGCn/ucFEAYK
S8LoxSJPnTg9OLZ7VT51usmJ0QdbVNPRLEYc8Eze1SOnboG7oi7YJjoga33RmVPN
ZZfYx5gylkJ92F8kSUcu/3OQ2xj72ZW3NYsC1BCIHf+X/Ib2npMOYcyWcIB0ZTzM
OLhWcUSTMZk6+NMZl4gSvvbNSvcT+Pe+gg3Y3/I9xOFAbziVeXjaUw3hI2ACgNnz
T1KfCg9dKC8CqJcBduRXbEk/+f2XG3hqD/wkdNrknvJW5ESX0tylkmeHmieVqbf8
pgHhJBcHgYnEPnJisAGMR32nuXFEkQfvVig/Ongomk9tT50GXiJyXwEPQNQlJLHk
m5SaLVuk56MVkqBS8QVkgVrWq2YnlGR12JKrhCmXNF3r9D5JD2+C7L9Yfjbpvtuu
q/RDtwtRqBZph/Cjyny/JnFxLDvCuKD4E+bKXMntWasH09iHyrRScXolCY9BxizO
3n4Lctdd+cgqiEHpCQvtdZaJMnV2/IJpxb6RQpKV0iJ5O9qiO3KcfhG4cHwAqTxX
XHlSVPGTC4i9L+AvkXgrnBiqhKzYbVvmgAKrZqX00D8DqA3zDpn0kXoQPH66wALF
7TTWYpStx6ifsmUpOqFO39J12GvpeGa7ANHVIKykL8M+/ZcqlE+GtGKfiAcUuPgf
c19xLx1OX4voD8ZZROQE83ZmC8duq8WOuoOkaN81syMnOd7QOH77UPM8qNP7SwEs
Nnkid6d7fBbr1PXEXmGQ2x9gBel/fXooJi2de1BJa8XqctVEzzQbpCGCY34EpvyM
uI+miKQ05WKGTBE791ujvepvnqhZ0NU+EpZAAIS5Gqq3HKeGSmXAyGfkMjfhUAHQ
pnEdhHn+EpFeQeLdFFbzL++4C3QdoFTBiXul0K7Ud74frKGQt7ei5xaFnclYrzN1
7msSVOtAtxw3Avk6T2aWEaQeCSG7AIQQhcpUCS5G1he08LeG2xnixyYoiFXIzQjg
kkHZNhDUGsyRoWBWHNzyIUc0x1kOznrleEMDENG2CIoyNOm0wTubA1snbqjtXarf
Fduo/59oBBmHcLtXQW+MCu0uBvM8NOSaG3UXh1fR0YZ8zIsph190Xz/MyE/oe672
NVofrNNRS8IlY4AYSr2xQV19P8fbOn23ZsflBMObrFQ0qkcU9ON1+k67rZhPSCDf
YNPr1tKW0o7xRwZrlAizyh0g7bj3pB2MJDzbEy9MOLawGT/I1yqrWB7croFxUijG
OA44XLDIkq6G4lfhrPBIL1RDt4FGx5dYQnIXkvI+YNpNr9hsfIpKz2DrKNAtIS3Q
X6oNFBLYyoyrGWIzdxEN1dmwJF7XFVce8ptFa6q4LFo6OXaXqGixGgq2JVdrDtkj
bT0ZSfTFK9bQmzCh49z0M4PgnpkcEFvobG5Y5WpZpAXOqPLFKj19obRXasCa2oA2
KGu5BIfSDQY3tYbf5u8af/QHYGj3KCm6Fv1+tTBLJT0RHG5VX1K5C/mwqN3pmCzB
Gw4cUBzUh9Z15mNCw3xHi1y8JthCGNSGd/pkqPJiMIfV8wU8qc3VqbVpfHkBUijU
lNWbHx7citUudfz5W+Cpr/dgerQ/R3o1Jlh3REEcw7X1umTGn993ixHT/7UPSQwR
ONrUnxXaeBQX28EpTBuVVBYsJOmFBvijg541O0SyDiSXAZOWGZSx8QJDOydUzz5r
DOjZWh/1aARHkhaQEBb0BZC1bCh0x+Cuh+c/hcSXkcXtzm8FYMtZLr9kBQD0uGQz
huKsmdMpk72HlQVS1EPKMDxTqk9MIbHdOgtiHQGSe7f6MAUUjJKbXUoXds4M9Dxt
GzGKjICA5vJ3Y+drvKjoVgz/k0iMzWxINPVJuW2F6ISIloYHBGjkTZBn6HRnsn72
qoHRULAwXcoVXvN4iETFkLamDDbZ3P6CjPQyub2tAcKaI6dNSp7zuINyDXUcWhwk
tsrKq+m8wlwrqw+F087p/6am5XFavX+qqNvBHCzLdC5xdB0YBztQsHz+Rx+kutj9
NnpoR4Yau7skHZKKF+JOrhtjjUcaJbOBGoEFtak/vPnPoiB8xvy7TjQ5UU0mXf9k
ALMza8eSSQhBEI7XqjDVMTro3ZF95TM+K/eYBQQ1MAKxUlIARNn9wSz+BbtVF2Qn
GYj8N+O5iBOiEgfGBK2qo7Wjzq8AY97tjrmK4h1vAM7atQz5oweCcafbDG2x40FR
/TFxVSTM8HD34QjjRhLZYDN3cmvLdY6yiGaxdItB9ZuBabPGqQ5CccLzP9XFrG0p
sZBSpQKCtL5M+j9No0Xs/7ArQdefpLFG6SBGVAHLzT7MDDESs8VuLujbAUpeYVs/
aHMdFawbNl53VTSVgPS2Qfpwq5MUBlbRhDYChBeNc+me/XFT7h4mp2pihDT2/5sR
kSt5Lnb8RfX2RwwLMvCWrzzqnXCSlTPgFK5SaoHyot9mRR7H1WDA2WO4Ops+CYZ3
Sv337N+6xXEJzMOek22ypxRIUbNXl7uQWcLfMgXRywyKk45i6shFafQclWXge60Y
f8fg1aRWxJ7BdHQxZkWXsVIS5cTLWKsC1eFR9//7Pxd3irHWmDyxXgUgEsDoDoEz
FJ/boGCV1c9Oo29KLD3GEno4tY9buDXovK1RMMJgqwP1TZ83EXFkUIwPENcVS94k
3QMg9lub1Ypsks/oFjghK++v0ayTE8Truhzb251oHUlHErFCA53leMjbwq/iuNEx
xr4El3cKai5gKfp1Xy8/UzRyB1XjzPMnTVT7NPsghjnpW0lJJyRjkg6UFW6a/LNl
KboUMh1CpfHkU+JDtp0CB3LoI4ck+zKTUsTJ7OhMwwKlEyexz1F8YIkB9h8sDpxT
xI93mhgbtfqsCL0iD9v3PmP2LkGlEIyR8enZ7gyk8b060yEC4PYkN0lJeyQzxKkL
Fns4YnZ+DnTnUUCpC5GXdSofa8AJofGYYtdJvb2h4YqJGMn+U+gcx2JTgWuqHG6j
BIZZ8zev4KDAzehZRzopN/b8yQrdx8OlKBrBrbddRWXOJACAmZkP26nTcrgEu2E/
a2NkEmECqZd0RZVxk/R8yIOBoeOdTtRkXvz0yd9AgjggdOTD8dDU+iNz2mbn/qwJ
x3EFA1HxHCeWoQnNQus/RlnEF2hIlZvqLcqymY79FsCF49LshTv8LOd9lvsN7PYT
dUMdw4s6ev1wiUobueQMSFWQxku2hbEl4SmrqlgeRu0+cnf9UdNTelVoLwA8J2sT
8Qi9PxUGbxlGCZEWo2hoc+ERqBSuMCQ3V5+NsYjk6cLTv8pWdjYnSF/F8PeaA3Wj
M7iwbJqF9MIlFu2/CnJjeRuKEH2mikJPmSoaraxz+w7LrFUJlVyYK9C9+zABI1Xd
ODLOSYMr/BAdz7viOM7L+zyy9ekPQLEwC+XKc+dPKI1v7jeff+0oqPmStbF+kqHR
84AphO0sixBvh7o+igPrgvcDQ7u9RYhhluoq9a5bm0GAjkOMLnf6nOOomgcF6B1y
rOR7FaWJBwsbJjnNnzAoFUKFjnDiEBL43Fyq8vXbM3soJeV2fWbIWHE1PT1QkLZj
SO0mmS0UqXvxj3ZS/pHrKu9D/Gkv+05GQK0TOTd0TSf/a5yALKtfB1cbn3cAY7N8
W4zvJIRhbdHdoCyB5QVK5WYg6QjpAJaM97fmTqPFpdrdeKv+XnhMxuEj7cNWrHr6
G2F/5PQgyc/OrgVIN5KIGHOhDKeuYETDBUinA3CMxu/jWP2nV7GpCbbMYwTMv07K
vmDKbnM/xHGwgzOzZ9oVVxuYGWjKF932yYMWC6F9CZbJVyp6JiPN3FM9OR1+F8B4
W+2E+TPbbg1Oy1ch3TZPIttiUF/3UwMCsuCjtGxI7yD/Q4cg8XBZtPPcEUmHQKVR
3ANTWD/1zRo+ozAcCsgIjvpFklpJ3pbwaHmR/dQA+SXaYkoiCPvmMzqLIC8mgvTt
C2MzaXOa2dqaG0HdNYE0CGrHYwcosaBg4ZuieP7p3H1840ULp34EM9l3SreigmZU
Fx1SPnRCrqlNlX/P7lbpgIB6DBBkhIfXdslj4IsYWN1bSK8pYEObVD9rxqS4qR6j
dgNz9/pdVLRSZH3zVyJgtaijdG9w4S+kP7SHrxc/8yr9XbKAmae2BNAUj+yHIjFt
udn2wFV4PMjRkFofAlDNb9zxJyPwdNCkuQEWM7IhGpeWRcOt2WREM4mN6emigqn0
BUKYUFdv86oTcEA2jLOp0h5kI7trkaDJoJMh+J/TuLD5Jq/Wm1iraXDuY9wZbaln
NAs/rxZZOqnifz7O4IOHCrq291sFcUfPtiltbH8tFroFwX9z/1GMBIm701wSIXaD
aTkRGLp3Sw1jByzYmvQtag7tKR8xCS0kPKot5zAV4VEQ/FOfctoHNoz8oOKvCVDQ
ZRJLgeZ4XlWSg6DZ0Cojcm6Pll6kqtQIuEYSYJgw0WDW4jpVamwqVZx7kuSW3XZx
TqBQXLlihQUt+0jF1uYa2WRMPhWl1o0s2XpKnvfFzCfzNthblH/jEbUfZn23b31B
m055Gym/jGFMSmNErhkXHcPWrKbvW1W9wck4PNBQehhFvVSYdiPd6BkbfKygC+JG
RL8AH9duReaTNI2y6IowewxobF8eye7p4EES+SQEj+34XCsAXnjf17EkPz3wkRkq
RuyiUy2t8eKFNdTBDV1dHAqDD+rZdU/laK6DKQpcpHmMi7OjvDi2polOaUNi0B0l
ZQTgHRFWSjDFl0OpZlL6hgfI9rNRGmk8NrWpNwInc4tOGVYz+eWeKqfFCB0mDd/n
mT/QrDWR+s7XeusevHcuXqWmreHx4GDnLfHeAwv5a8oy4kesTJJGLCfDZ6cp+5/T
EMDwj3HDGkePaM8hCo9HBfDdVNdwIY+YJ8vl/soP00ad1DdxqU4vaeXJ5HyqjZMV
Dlo2YIbXFyhv8cWc7430wFwK1TqF+8C5MY9+wA0kFKVFxzL8o80YG319Eei01b2z
KnjLiLqmuYXo/q56NTbgi2tTPa6OAgy9r63Dr1Y+5wehjTLVCbJba1azAKz6NfF9
hqLcSxDyaQrVaqLhNXsEsRifhB331M1lulVuVilK1PvoxPHSGIAKmeHSMPiNiq/c
SjntkxjTTfSGPq4IFfqxHWmaMOSAXClz1bXoZ2VmNP00z63jsbUggYtp+oaqd6Ja
tip87DgAp9F/lcgeMzMjiuHVJDIAzcWi5ogJktsr6WlNemxb6y4a552dOPYmQqxI
EHNwJzjjauzjqIPxtumgreNPZWVBZhxUEXilRZrtV4/rsl53TJY1YLGpRXAV2pCx
keFZrq1mT9/Ax/gLEoWqHY9vdvwGBy55CWToEomhH9et4I+N8ABYebH6+sRkhGqQ
t8+4uzSC4Ye/zNefXjVSFGWGTDeCBYg0EgQGUPCFx/nPUZc2xuv2cvbaFUZYPyZ4
VipTvGK2zN/uQuWFq6uZgkZjIQDR9I9Zc2S1/al7U6AJzOVYuyt8Mk+fiZUI542n
LNNHRhtSQOtseJis/96IsfbH5T+fD0n0F+AKuojuqNyDpTeqiSuOqaGl2qhg4zrL
ieKEzUDWeNM5Xqeq2s4ECxeizQ2kvIhj9vLeujOusHTPs1wD8IKWgrNqsg9vCJsz
UD4UwUrkVt0SNEMekbxQmZ2JdVXEeI5apHlXsYMJaB5hnKyOzgvJWlQEqp6jsiwi
gOABVOgMpYTYs6HrR31pD2yBIDQmOBKUcW9llUxkjTV+93t/I2hntwAzorqg/hVE
qUeRfefsdaAX3fjWEw5tKiuZtSgVS2pknMRksoYlUt7D3v1h3BSaWq9e0ipDjG3Z
kPonRAGZEPw14cffW3lRkmhWOU40Wc3cpOsTuIpJyZj3ZVl6l3hnfZvQUJp2feNl
sGvbOfHYjoo3rED+w6wmlFjcjwRHMUHphO65D5hTwFWUHCq/zYlI5dOeX2Pw2s56
p9zxjzmKEg6ieI39zyTGgvdyoG4eCF0JJkydbShWWu3G+4129bCzDXTCyfWiNB0h
UiRgZfHZAreSUnv+s3XaIzoKPQHgAwJBxYWhMn4qc2Kg0BtXDVAuW06lzgWaoLqS
fweEoDsrLg6KBHh1AX1A98Gq+3FlhK6R3uKpteK07u2qGs5hG+v0kj7RaMqVYhGn
8OVDUya/cwMo4X1sO+kESjiTqDCWc4H2kMcJbJuCbEflafs8zY92il3CwK1wgO4m
v6CD06jO2kUxvH7z83+x7C212hklB1Ybetgqq7u4z1Nkmq5Kw1LLK/0XQi+h9U2X
DNxHF/IXUE2Eo/ncDPIZrSC77PnmAaEjpLm2+MmG43IitWYqHvmYUdaINqTb0RgW
mU4nF8Vkh+DtiI4lTaN8qka1cMpCVFlivEqaUYJyuPTmh+JX3MUrRbneD8afBnro
pe7HGoVcznZIkjlnEnAmcewE5GQpic6DkyyBEifNyyNjZJDXlDTQIydIXfslTqvp
40KjUzgTpvMobqlb/17wPD64NNzGwcaFHaZc8Z9i7KQR0lCskTFlfEDKQkxXOvG0
vsqPtld6PoYrJhOYGBKu63QNqGsF1TlUhhXgPtyfYJIHE30xqSBZRKDbXlstvze+
29QptnkjHenY52t+rbwS4V650i3WcamL4SqZvMnHqCtInbROJ43pp8tA9Pccvt5I
IGZ9e2pFpu3p6vbiGSuZpY/HnRgb8qStN5kAROVqnQvJcchUfzCUKfCh3ay/W3ne
2PwgWzglShNClByPuSPgIEA2YxrDHEbEQ4JNBPtHuMKijfaKXBf/XJxoVvs7bs7J
GOVe8nDGmONiJMxvNh+LZFIaa1gpl0jgwNr+vHcsCjUQHkiyLcEiGTzegsum7zwo
8aOQaSV0G3uxHwQbJH47HWXjz4Y+rxlJ/ChxGynXXPTy93S3yQRW3mNetKoUUCrs
paHq+E5ZCrdzijcER6P1hTE5psTqg++HiPeLmRa/IEg2WZjgqj7LTTzVjkJVVRKN
IOu7VpLKaDKCO92FrgiITWL0Hg+k07HlGHG8LAw0d8oMWUVpedPm0ctk5Am5NAro
4mOKG2ecoK5GwVjXVlhL6UAznpc0tPWx37MrDmBz0fXONdP+srwrt5Ss38x2P3w+
HF2KBvkQvSDL5ws5ckeTJWcZYqcZqM2rC1M3WZqwjfDGBGvIRhuDl0jIW1ONfwh1
av4p31pqIEFzVwYJ32xrCK+fU6y2UnozvUfmOFlvp5wERr5hLS7bgMmsini1MWsp
4WkkxTrINQhg0MipSZwWBGiC44BIOOwCpEjpYJifnUgHv+cAHp9RuAPWDU/LEnNH
xHuPLO6n1RDb/wECHoWFRSLYHThpGWEikstdgLrx5CXsHJMsCedvsqDv/uqTJVnz
+vOzix7H0ggstQkNJ4jFmUbCwLdBiyrenIXBVeJHzD+4oGHdyRrXiGA15lwFA8ZA
5gje/K4k0CZg9fBODNVmjjCSzvA2WnLD0J6SGgfCXrWiEr3KF3MOFvsW897nwI78
2mJiIDnAKUGVk/2I8BFawPq9LAMlZUDY17KcHMSLlwGW+8s2zEtsxTgZYLbYVPLV
N7/cRWzfAfn68G9kV3VffkjsWXSSEqJt0g02DFKmSA4HMX2WuxArfpTOz8+60XA+
RTv0G6YuIWMffvdW38HOnco1dacm8YAfsPIez73jTDti3U+GIk6CxHbMtZe09oYP
yNlakgLRVYT6GSyn6VBgLMEcjpFotkQpsqDX5LMxBOUaQQfGYKZFLg5quHP6V/uZ
OvdheBVxHy3uA+q2kfxeV+/j/9VXmPWzzs0wIFcZTpuOEZIkzXBPJCCA0LhPYfg5
dbFp/AagxXB1Y0RZnD12ROf/SUMC65YnLvGHsb1zTiYG8cbU0Ao0zpabsRA3hOBr
D5skKjDdAvZqszBJqFTuldgyv1ZCsX09tbJuPtnQFZg2IyEAk0rTUMi59/rw29xo
hT9QQwQH/dGMNpysXKSfNCvsJymeT9K2p/097qDN5JFvtheTXLskBECj3f0SuegC
bGogbPDsZDZm/97x8+CRXkTlqJksBx0O3n2/Y7Smc7omd/2Py2j/2meVVz8gHcnT
Ui1qJVfUhA5Rhfkbk9rh9y3VH/AAzE2FH9N/jkW9Oi/aR606SwdJay9v8hFSasEp
fz3+eJUiShHVijNPIGMYHPjT1yqMFiSlpVxW7VeMFZa7+iZtnIz4bGZReg6VBE0Q
WWKC6qEomXSDGkEK4QIfJRV4f41LQwhbB3bM8AHxRykjulUzvyTuYbkGxGdG/vsI
Lp5PYPFaoN/HjtPpDl7MOEbYNnbyjEkxHRSPE5yCQ8dvfj+SR7Zv6kMBWnyNwFZy
Vj1GAK9NWsbpDXLWId4A6BjN2wVirVuNdJzbH4Vj7ryTcsKOY0+tOt3KThrl9DxP
Ny/Rl4FLAjV/1hqibNlu7keM6HCxumxQ4XTqecWIHl2jOQz4t1+X/ESHGYna+6s3
7DUVUEfkW4G+LZ6oPEaH2dubz0+hNaTW6QKSGpDDncvaU8AFQihkG8AHm3CmDQsi
ZgDfjJiP5sAKnR3JUXBZV4ak/Tjl8ahe/OBUitKhVzrphZ0gkh21icQEcUq3lH+G
fV2Ij9cbb0YrzLhZhy8+vgp0PzkPXa1Vd/T3RU+KlovZbtCLX2sFplDSemou/sLy
Zjpcq+eEyXt2/0tt++bowYq3MjpAEnNyhxwDELozjTeSOBULeBC0i0sRoji9UTsS
0cz2ECnYyK1nybKWHltykhvy8TTZspNkI/YlVxdjB342wvQCfWnTsevnFTPsm74g
OnxD/t/NgCOHi2x6RdiB1r7lBJSFW79e5207z59/uii8IePPfo0sSGsM2qL1QfE0
PsboYGhUT+E4njWEzUuJ+a9qqFAybUC9F2VWhpx+BGpnbwixPyEdxgbbNs51K3e+
ucU4LpG+/CGqSnVGUrn6Rgq+SuOltjMoeH38rOqp8vlURCh2gdlBqfMzKLKmh+CC
5aRsGHrP+/Quy5w1o+Zp0utx27qLTfkzwuc4MvGTBwZt1IcaqYamg690lZaZuGvF
t9JdAnJDkyK+fmbMzArNyQFNu1UPLxj7h+dWxWb2EiUKHHkzBe2ITkVPV3zuH7Eq
r1XAgpKtrQhk5ArQPu32YJ0UDFdIgKLeTwmc5msuqlU+lXaoSdnviD5QRmG5+g+q
0Bp+yOE73WKp6dBAaQ8+coTIX9FPwJUBxf2wxdxgTEQDiAgcLwriJes4HOpfYmnL
pedbGI9FClwY/BZbJzF5LdwWWpD+wdsqJ77UzJj1iEJBwEmPUxSR8QGmHZissVdX
f5YHWVA5eg6QrunQUY5h74zEQuDrThTw9lA6rBJlCLFA6tObqJvcCKqV013faf8P
sJPYoeztmLniY7rmBuOTidofAFDVCPhj56q50ukIWPRVT2ylM5WvvDVUn8Ee8dKP
TV97L8ypsRqznfFCjGQ4ySRSG9oABBHc1jKahU74VFaQwWB/M1kMyD7mqoAg5b02
cwIiOdGwxePup5Jj3eCkouxMp06NEePWlhtrOdaFAbOYspmcmU4AHF6nXR1GZAm2
O2fg0jmrYHIcmIOmhbav1WGKcLHi6NFPQeZoOY7M2YyflUBVzKtnfOeUPw13YuVk
cAfA/FJgByZp/s2Wi6qbiMFGGC4cu0aQKdHJrZK3LuG6DyU9pg5R7hQzSlUb7lci
LH17UGnMbmsJ3rNP1YQ3672oD+/JpZE5x1BIu0icEYUmX3RBZnSgChAzK24UJVZ9
orGO8RpzEkOmxS9df5IizFlNxVRLjAh8FnI7/M99Q0r7hRl45RH30f09XEct5+Uv
B/7ipQ+GOJKcGkUsfJL5Qv/6/SkTFUCmND7O8aPF1YtI+Mbr59d3vupJqyeKJm3h
tWMXBSHkAD+hf3IOwFyzL6q7FKuENGpbs4k5gxxMlgTph0CZloSg4mFcsIN9KZPG
lNs1s8f5rhAapeKO83IQYBETBTayccaN7msK1pOyIMwtxtte8sMbM52Ag7gL4HT3
cSWX8d16aTjGqUS27+rT6SmGS0ik+ztm/9jW0xXIJPSM94cQ8sDPOJNtY7HrERTS
NYysubEZmqujbqNhYOGEtZY0lOFVraS0GMXUg7sBNre+aVv5CY7HusCfC8akrEjT
jde75OCJh9pwBrNZv+XUpduQ1RyEktmz+OjmBIZFivi+/L+wB6TNyezdBUm3O9SO
bvYhn3OR4kTAe+mm10wFC4dZnXkiBamcmihsEpztk/DSsiu/Hzb1S8I+cbBf1cgy
VgySd840hvHCKkvYWfVqNIX9YVYdCUwgKUixPWsFrtErLyjc2C0Qdl8kIgJG3Rqm
vvFdn3d6n8yBrS0RT4iiHLk9g1MRdcOuOXfIsYZdtRrl2ixCexa/aqLWJeLi5/1F
t4p0Hmo2VjtVHZiXXMILQpWfvw41+zfePFLxuzpQGvi+pQRg9PgadTlrpMREkHS1
YZrBGLUP7ve228f9KpKzx62k7pb3j/kSOmYV+grYV0K6kB+45Z+DsjosQTpEA/A1
UQxVM18aZe6VFZqFn1TZZ4SDAR7mbsGOhfTo4AvTBM4iSmNlweN6C6KzM4lyR1+3
+VYneOIukar/6NB3p3VgR152ToMKkADueRWZ9uKIp3cjM/bbzZgmRV+py2e0mZsr
VlftbRJNk3aCh4O52CkYUjYegq0xwpzlwXqlLBgOKeaFmU04o9ehd/sIRMo+BPB8
vhOtPuQpEHK0jsJ2SeyF+U8AIkVtz/V8WtT5lolypELL1Sg0G2zOaxvkbccWrM8n
nKBwc9j6R7qxyPp+kLask3tAsROB9vIuSEJPolpoYyIPCQMZ2YMXxfxsj0PFmqjg
SKZLvXr6TqUs7M22bLabneO0J0HSfJoQNNURe+Td6WmBbtQu85mkuKY6tgZN4qMt
tBkeelUDOx16GBVsrdmUk4MyKL113+NWks3IyTlLfRWNLpqEZFUBS2HbZFN397V4
YhKfDOhkXkJov2+avs0Qr7tAttBwC32D2QricsfFt4KIQIOWLzzwBQtu0CpWgbeQ
RxPNIxh6YAYxMMQ5yP1pGduEKy6vZNvZtdFVHY0TnaKyijwyh+BbxH+Ugg3HJ1Mg
OB7z6s02KonLo5pjqqYDzWef+qJ/PjXxk0jSMDzSGwAYySG/V2EbkUU8p4DgNLGE
k70hUuV3ljfSQF985b/InMQuhej9GIuC3NaD7MdgSvVgYpzSDMbM0A53V9ohuY6u
iCAQzadjDo/ZcKnMbNohWPB7Hi/19vs/2Y0Gq8It3yoZLPSYopADLrx6xee1+6eu
tGQsMZ0hVcLi0FB71fwO3fp+hoCmZrmT4vMYSFS91fBgVXHqy7X5REaSmWAmojNz
bRMEoU8nSgcE7zD5Xstz3nZyFVt79Zao9LsZCUgmUCj4MiPLIzHR3beEQuvUL3tI
x1sKiAiR8/tpLAtzwb/NAd45FgsbmikqbHZ0CQuBg4OW5/S3NKHumBECqPpeDVS5
T4//POKwsbCXB/7g5PrQA5mEBg8j3M7gyP57rs+nFGXvkZVyAsKykM1WTbiUlAYg
c90KeugOBzKiaN/sMPvv2Qcf8uQmp5/q1WYEkQpX0tXn2jCUiwqHrGImY/W6+qTG
/Hx0/tc6VgVb34H4AEihfyPzBNPxi9fOqcMan8FEw936qetDs7bDmN65fc82dERn
RSi8/1F818Y1z15OCscGCiECzhSqRV8IonfIlUkEYwY1oY3D9olzpykf0V90oAWG
gkCfxL6CFfzrpHBJ9dylmcHrylDA+VsN4Jpc0AtyprtNJqwMPo2oBG1eihVr6p/b
iftPGzThMlYwtaQlU7Ra467JPSK0gUDV1Zp6iaBJrLA0VUGzvZiWgiA6htxJ7nRz
2TDtUKJn41VKReCJ17/MwPkv04Co140WqlrEOEqq4eZxOCeBHrrbbbqQZ3uDhffl
TzfLIOBokGkdfnVqLJg5zZaa+/35NIrh5HV1++YYPDjgyaSsYeI4jw/7s0iGiJR+
8a75uMyQbqYuDF1vvZNVj8z7bliyJ5FeLu9ONmKM4si+YPR/JQGph/SG6zEV0BDm
mvfHo7VToEbmKOnRon2XcTR/1WtPq2mqxSjA3ucsZka7/BTaQQOeB4fnc0lGjcc0
hT6SwSIbFOi3JjGjdoSfRkTC3abmOQaYgmLypZKXv0NE9WOEfidLjNfmdj0OP/3m
efsegh+kxXFn90reEp3uM1XLfEmdxz8uMgcwTw+GCF76eo1YFg6mU+d6gkf4huCK
CVO09CiTbc4w3enEsCebUeJykc0FhSQ5ENvM7OgZMasST95gFZgEM1HokLT2lucu
AVKgkkVkNdV3LDGL/Rsnn5AQqU5bducr2eGjHnI/BcXnTy09XAEz/2ZjF7TinOg0
qVj/eZI/Y2ULSX2KClWTcW15ZC1ptrDuQ68tT3q07srJPm0NHQ8Cw6d+lE1uxNfV
wSTYyRcdNSG0JFTuYKdQi8NxSSI8cUF724nuv150L1t23oXGN8LiJWHV2Id/WtbZ
VFW9T5YTif9pmwOZPn3C1scyfl70//Eu6SP2gbZnyL/dc0MI71cRiA/kX49BbRnd
3dx42X9vm4CqL2Wudd6+B1nqKOy26FROuhRtHr+CWDqFTivHSDCJK8Adoa3jzh5k
g5cI1Xv4K08vXAoHeC8yD06tpqp70Byj+TebnUzA/ZuIhm5LyUILqcq9KxpPs8DG
rMyRf/dBdUDYJ8xQv4nCFJNtdDO6GsXCTbI01lS0iRZ3sr9jhqjQIKJWkehqRVze
tUmwwS82n4ArGI30IaOaQGhWzT1nzzz5LjNsyYLKbzkMgr/RRbw2r1pb74Nv4kBp
8sfhNhahDmzsPSI/AztKHX4GNJqkP7XCAIDBTcrD02Tq1SLItwEB+D/OVeGdUs6x
gR9fNNxFdfeMnjj5QqI0bOX4AlnBeJmD1n4mnaXXFd/IWkUnYVX4MOC5FekByJtb
Eb4wbhvUbkBd4jDs2qRHJM+ACWNIJIh+NXUUtHZaXh7S3b9Ou+F+V+mZcUO4+VW+
+5/4Rxje/NMc4ZZYpKCBcFHAE5r9Fasad//EmtRTKlKoPDs2uYJaiYGXecW28vlH
gfaVKA3kT6PvqSPTI52nzJwynn1ygssgAfuhIADlOmOKHvRsbVxkCKvLk+K1BH7z
GEVmb2K1+uPCfi6Y69O0dCk50MmF0jeRdbzkkBoXPN1p/QUmQAUvYq8uYhrGzVOi
c//yazbZHypYY+rzrVHO3arqhwX5auksdGNXH5oNnF0MBOe6T47KlXksRPV6wbkx
uZF7O4p59OZPA4dnVKm+SuhalLHt5rdq6xcjcWWU1+r5OCASBphzMGT4CCOEIs15
MHMk6umi5UunT2leEnvGd9jXo9VKABEdhzForTaUNYMoHeuLXSoZ/ExLiwCgUJAZ
9HUqr5ENFuriDByQVD3MVvG3FKGdo1wKvYBP+qk8JDFXICGhqRc8HYyAloiaSWSs
+ILskLiNLMDHrRejpTT+0Hs89MdLsjL6pbLK8VLr445L7LKw+uQrtE65Y8LoOhNa
je4WWS1C9uiv3MHH07XuXc4hy4RMsePx7C8Jde6bJt7nLQav56lsnNpMHlUe+OBd
Z+n1mJAdyAFNR9/6r7LnSDw2dz3rRM/X8To7Petdvu/TIdOlj5lIjT+T2G1/Zm2y
yfgPQwASo4YlKNxpFebEZkpBtY9+TH4pytd9+po/3gznup1ou82MG+OcRhMQVcKM
Jtj0JfxGyUZi0n8PMLcGi/n3jvkyAfMFElzXyM2DIVkzL1bStPNzREMPieZ/tEFS
UqXuUGakFjPonTSf91KmWOBaoJPKZw1bkCgtChn1TdRvjmSvdAPYVa178Y+FOpWt
RaZvjvI7EbTkHnaEOUUXtxUt3rHoKfb6byKCzysEYccFH9INFNJrD7HgK1f70lzQ
jYOAHCmoo0c2E9c77uWz3myEX1R2kWKPd9/mrlxbJsAAoz8tQaOpO9zDry0hkXve
S7aXEimU5lbNp5SdsbeOpaYYuozbzDMLCq2ihrBVSH/LPRvGtXjJ7EbSy1SNgtkA
cB4qOxePVCQ55255zb3o9TMtAdt3snIBWbuNhS5YwRcE++wiZsA0o6SwkydKcwzv
ze2ou98+BD7SZ/54Yo8G3HQSv0ET3veb4kVEnqr9k0gsqUoq8h5L3s3Fg1P1Jkhy
KAIzIpZJl3+DEXhWLz+COjS8nefW8KOxU102sYYof2evBXNTVYrtHo0vxuRR+Sdz
JX4hGfSbxL+h/u0qBCe0DyZv6/AzQ1e3LupfXjGIUxxJUGdgBZ407iD5xeXr4p5C
yJOyaNra4ynll0we4syxeA7PiyufS7NRpf94jxH7KTSY2uWd3NtgeupQsI56d3CF
slyPycqHXpMs0sfBczrFDNmsE2vFLKsMGHMHueCS2LWBv+hHGEYEMuWP6jDFTuun
KUt2NjF1jwx98IyCrROLqkmG0bl8fyrfsN/ploYN9W2OlMjeWY7nli3yJeCNlfZH
3c+/ZXIbyjZt0MhvbkczQ9FKFoeijlQlEI+g+tO7SMuS8JxJnex++CPHnFZxyza3
iIF2zf94CzkQ284WQiAy2QWw9ZfMkAB57JL2KcjquRnLstn7QW4Nf6GxdPJ0OSdz
+4HIeBOb/Xh9WOg+bvNnIKWVJKpzQOiucYus/vDEL4N+nE1zB6XvdoK9s/BOJJZN
ys6PehLPZIKzrK5qWHcCr5NwqqnpT74s4if7CuneKam63XIj8/EjaPRyT7WnRpNv
cgP0w2uErqB73WEsA5IfBvcksZLh+lZi7p06IY8fqKz+v5OQ3kPmj3CMbC9OUZeh
00EPkM5gBcaOPNQsClyqrH5eroAHtaBIUWoj/EEh5srbAKZ6Yzl+pgl41WcugvUn
9ul6/OavOqbHJyIPCtkd858YxTVrmoH1DmMV465aFJDOpm/PRfBRI7RLhmQA0uIV
IEu+yNuF6uZ3h/kb5IFPhbSjHiHg1d+MzpbBFvfw6zQ9tk3ik+IohzrcMRZQ8HYp
SsUFW//eTMTTtJwKpSvTl6uAslIdr+QvtnElYWhEcKPXaUQlibwqWbxOnLE6I68V
nkhLyZpW8qsTWUFPSb907GCRYPqMnJaP7gtDhus40b7c9MqKO66cdh0mQjRhuRDJ
Aru2a996Hk79vVAL0eSJwJ36jsHTGVjvkwW/DWCBddfSMaoa8CVFCCFct6GY55Jh
qvtbgUBD2/63LTykH61NgjevEaxQY+vDhCfyh359kweVIyKTkxkGrgHR9sdjyvZ8
xEGpBexgXK/t3rHo5VeTE32oQsuIjvApd//N/9Gzj6dcy8+K+HThU75l75vYbXCw
O8hYbvUfxmvtaQWtKxxrwsPm117MDTkHgK2sDKUOfw+Enr7qi/6CCOsBqcyCaX0M
TGqweUfJ8QPccTI6raPQjTqymUJxXhVrkMeromT9mdPbyMnQvBNwQ0F5qEieOvmV
M6MY29OvIbdJkAGznGLAB7enPcKSvMn6bdbr5WH9Q4Fvndf74CMeqvvXb/r2O2gU
zfVqT0Vl7HxRt4xaAyvtAd5i75hv0dXigDnJ52oHEMCxyVYRPq0nR5m91qj7PAB6
7ov6oiQv0U3q67npfgt7ekV+iN6kSmR8X30tgws1jK2txGFvAhGufvsq+fzaIvcr
VSySGwtQZ9V40nlA1dnkAEpC3r0F/XkhSC8uYWdnxMyntvLFWJ0ZLSTIfNrC9PlW
50pnyD5jtAEbEO6LIJWMqurFdTIbqbH+4+F7GQFEjGxpgG2VTJeTSqvA/u1F8I/C
x/5dr/+27hnEOX/3A1O+qeWNxN7BhRsDUt6Xni1ci1jiaSblEFi1+MmVkAOeGDew
TSVOe7HeIwqiTN1InOniWHmc8TV8NTj/zG+q5ugulamQ0P0rWDJpzy5WFCbtTWY7
4WfxXRS3Pa01RKj/DVE68tdxIUB1OxiIluZz/IPik9+GaPM33VkuQE83YviT96Cg
TXyflPRRREho9gFUQ5xsXfu/SAFPS799I7ydOpafYxNQUnnTHCFxd/CizX/to2It
OLxNSLSUqpMr048gUgaP1oiWhquWMGhrNFnAtorPF8umhxbTYF1997vSHy6PBrED
AL5pIve1N0OfKfkjNRblIJ/U1wNYLPMv5pRj5RzHEBZXLQh57zh8wZOuQPcOx2df
iNIgQdbX2DKTuDCsDbld1JXlrpht971o9Wx3ZATIvu3Q6aNcag9OBjb7rM6sTDfQ
jXeuHNZqnXZYg42qEfoobBVQFb2k9TROTP6IT7q6Uhjl6qSgUfm9tlaPcBvzR3l1
+1MR4qy3By6T2KqFHZmGzsWJWEYPpC1D0st7xcGlAuzew4zzgmQA8t1ip2PXgAke
rZrEz36QUBLTHbT5FseJxHd2pv08/q7Af9sDJ2+pMU3XED6GC+FG4CnpYKvQSvM+
6a+BIJlBfDcYUTfI7MzBI4EBzsf5wZJL3qOCBhhaOFlT8YDl+8xTusUMlkM9Tpdg
kmLDe/vEL3Y1zaVjs779SGJvDYrKl+CduAuCmCDp2t1U6sUDAommjNT06jqqLkq7
HOW0bdWVnq4Elk2klt1c5g9ykhd0MOZn1OgnlFN0cEWEM3MgTzYolHx9PF8sBWT0
u9xMoT6cBYJqR52Iv5UezVAovt25c+JnEiUgGlrLUbSzVNvaP7GIKQwZ1CtP0zxY
6qjMaktMZxIbSxm7Cq7GH9GiOflI9gJlaFwJzu1RTosp3GdFNakLkFqtMhc+3e4+
7PK2LF0EtXxCzRkJ70DDXkI/6gnUfu3n3HWyhrhl2AVdvZRStj27d4AduS3Y1SJN
RNPjmmOmLrpmt6UbxDt5UuXNNTluULDliv7D1h9emRl4wOxqCHeLPnLNIh9Tsgm1
uMeO0LAEtdR3qTA0sPuMdzosablhFiNimuTpApLBZXbVtlMxAl9jU61Hx0PDHtQo
BnpsK7T7cYkgb13CtM5M/SlA9lihRTGpef0E92wXGzbcpVadVNPj2D+R9BtIKLPn
ZmdxrR5mRlJ1Md+bvO5FUOd00OnSNpcGdouv8Rg4dMcbe9s8IA44WdB4/Red4TtI
Ut5PgqrpxvQAPljYu2lE+hsBwg07FmaOMGHMTnMIhpeGDxIrKffq2nLKAWgrnVIC
VIZAWkgVOs459hGdB4Hhn9g10vKc1WFIgYugdK7JVWXOmP6edcTmRuGTD8fw3qOO
Y8xnOW6TbhWdlcKBi8rZ24El4MFOETwCuxxQ1MxygtrgUg4+80P5BISePYR0cNSq
W/AJfrKRoQLWZW74yrfxmRbVz+roh/t/YHXQZLEhkcET7zuqfL3BOoDDVLCSic0/
mCivWatdOh/wRO0rwLoIujN8KxO+NQ7MzgiGUZAGqVWxjKw2pa2Yc3QqBTQefIwn
rtWQbiVelYvW1Xt16WFzJrDYlJpKBK+E5wG1d+VjrPlDJWUyxSSaKjLdssLKTgfo
7PoO/J3UsrrfQi501EfjYkPZGbGc6UoYdNyLvmkVd5DIxVyX5gTZFz66BBtY9PD+
8GhugvS1bS3IgTsEafQgi+s46ww9ppPjPSZfudMdFlJYNaucVnMgsy8FG8wEAPRp
YWc9EOhkRNmnGwAyMFtzLYUMuwiP361b+L2YzcD4GKrE8Wvf80o6IY4E80iQ8YXV
54AChCb3sw9kWnLGLoEN9Ot1sQUx/5qHDdNjrhkrR3a0MnDpyZTDbdT8l1+0qHbC
kn+S79NR8UaOdPKtlOO/P+VfaCAmEXZ6DtZolP20FcvabcL2l2eqxOSZ3pDv98Uk
ffHOqGSxTlFQd62doQHTI9rzUwy3Vwww/jowPsljBCr9DGsGWpoUuFgbytTuDQm1
w/GIH/u0dqRUKgv82gvcB9Ha8rJqe9TkDBIM0ppel5fHKSBKb5xNlck88qGwQJKT
//TSsfD2roY3oNHAva/mJcs2kG0U8srpZxTmRU3Xf7pPABnr3Fe/66DIJy+nQKBD
alsefFO3U0l5MMEUKu1pVcAtG680wgqXjqf8q0FX9wVIwX3qzubLenfutVYy+2QK
lVEKyN3dwsl/qeagfgUFyj+7cc97wIxwCCbl3tXnqMwsmxggmkaXivvOd25GmetK
VAyAiPo541jUPFsacTaJNQwueR50p3/3GU+m3FiLQTdXN54FqYSx90o3p0KtjoT+
5eo7IJihqBP7dUNeHAqJ50ICuSBVZyFFLW3azQCxFFA5ezjJKv5WQ5zEpAxtU1yR
E8KKQHbtTZJjaiR4OzXthPmV95XjZXuCTMyGQuYDjxFnqbVRt4P1yRkbM/wKAjw/
LC2OXNssR3fGwY0xWRPG66WR8XNZP6ziOJNkwKjsfdUw9Tm/TsSif/QIWQ/qRqy0
VdOZLoUGkDCYc0YBeQWY64twmn+ZY5HWHNOgg2Fdb92AVeBYto6M8faW+TThd4pW
rU5lN3omYye6QP6o7lwmEyizBmZ+tdvuzjubxG+NkI1T7UTFiJWV+34WPZjI6Ate
atN+oJwZw1H3jPPu4E9hSS55gb2mUGzZfNOh/pj4YzieAxhuNecolL0QwJIS53Us
FkP3GhXUXOgCGQrJevIUg7INiWLG05qXszj1NjacO0LoQzHwUczGGXHk3SgV6bWi
GGBX4ImsKrIEcNHMPFaZlHpkaZh/S1ytWEiQv1ZFwt+qMyhAUWcDw09uxyi0TEvS
tQGb9wusaFfGdhS4MKubKRqjd9TpGK+Fns/9606862d8O19oX4kXVpY6exYYLZVa
/k0fwo56OY9iZ7+PFFPBtYAsO0pazFqbFxQF5z7Fe3RRDk9xnwALV9+RD0itk6+K
5ThUb/TRywRipvFPZKGu7YvW8zm2t1Od7d+0OLKjt16pEnbL6z+xB64czZbk5U5h
7x0xiWrYTHIHt0ln8m3nZX87T8bn19gCP29K2A3MqUyM3ZSJX6pIxpLo05vM9r4P
w4KeosWpaA7csbj106FnPKx6qPo1seUxNXLlqwKA+ts62uEmButrWj50slOnh6tD
HUJc2t3EiJTPbiArFokZAVvqCIXGhnqPu2lq5qSIdwKVMTwZY0JBGho2Q8xrGIWl
ZovoTP5M/w88Z/567v0SIvuidyX8u4vfc5Iz8CUYpCeu1xzEFZaaDeVZfS226T3w
zOdLYohZieuZE32lvMWqbEYIeHIGpgYeaQuofatrKdgjQ500+DpbQqeWar05/fTe
dpSlaJK78kKhWz5yWKm+bBk3qVXIP9ZibCO+YbgslvliWyDm+sEcuiyT1kOQ0QT/
x+gFg//mI6tzicpKvez/oHUjwGZ+KMeQCovYUqWAeW92F0IYo7MIvx7oqzy0R+NF
MpWFwy72j7tdK04h4W3fOjqdW6sRh2VARL9GBkshT7jfsR53BX8OjaOpTBnVqDdg
4moIh9Sv/uwXWwi52L+gtl3CckR9j8IFk0AyC45Jl7llrR/3WWIc56/h78PfVSFz
Am2GgIpHfLcuuJDUR9k8qNa9j6mYgCvBDWJxv6x/xhVw4C6DAqc+k5gxHsFbzDgP
3RQBcVKgstTApj4cqXW5GFxQs2s3IUwvI9Ac+ohgKfZsf5FyGAbiiar0YtPqwGAJ
TGUloKjSFBn20dHhptn3gXAxLSJM/4hFihnlvaYYb9Fo+dblj6qJgMB4FEJgcEsx
RAryxJIIyXuK2o4Xe07yXd/NWFS/GfzxwxqE8PtJoe2Lf+9GXmYM6UNBu6tkWFFr
20IVZc9ijMC0ZRq3becKr80OwJ5duN9IiBJsL/zX4q7P73vnycBnniOjaMJJz7a0
CsX+jsi7tIe3XCyE8GBwR92ieo/gGZrqZYTegKxZEiQzyOBQt2sGvpWwPkbQXWQ9
7JmmiweG86cwq0Rq8VpBsA1Z4HvrNIKYMBpJq/AIzq4yS/stDflAdBvsSoiDaunJ
woxLankd167tQPOsPoMbgjyQDjOasLvWUIc43qAtY8ShPsMn8XpDrSIwFSSGJa3D
fscDM4gXmZlLuT1xoLqtu0rPTPJzR1f0IAkCz+79FFBJgx46xLzzD0/rdQN2ZCQ6
t2eng8bVF1bR3TugJekgMbPYSEMRyKt5h4As046d6Jvgp+I6HHObBaodXA6/O7Zx
sojAeBiLGxWz9zie5RUyHi97GSXGzLh1WRjPK2qUAoDHPVlbBfVRDX3dsVJlVf+Y
MLW3U3hVoiUY/ApCJqftSNrjnnc6ys+21yvjNSFtWuoL6tGMzHcnAD1Jja00QpGE
XQcZTcfPTA7Bzi5GkSHSr3b9SUo57AezA2tE4VVSrHQU/aMMiD8IrF9s3y48sBkS
jVXDU57Ho/tQHfkJbZsbvJBaU6kslex6Cm2ljunqeythk2RV0V1N9HMaPzsWb+Vy
6wuxXn6o7A5sBXxY8zWRCEN6+G97s2SJ8jKwJBiOjQ4tnYDKevuGWphthBrAhrkS
hEbrprq3KAGKbUWgHRUZ7NyUw6bNq8LJLoC8FhG/BVnvx4GZp42yd07CfnHYrNEK
rvYznub3yAFh2Nb1fYkI/tVBa/pYR+OGRB5rCZWDJ/iWb+MsTfNLYo0/iaIoQj8F
UQz3vfU6avFuJjFmmJ6hODv2SMHvajVQGUPgho+pjR/GGfhv0E32cPFCLo8W9BNC
bS57oiYPRaMtVcWAsVslZVyg/3G45QEaLsFou2O80AkvLPYiofo6v+Ym71+cpdFJ
yPy7PhsUEN/PRxjYdhEQF6G+jo5CjYSE2vrYy2SuMWlNXO5kdXNzlw3cyEOLA+Sf
kR/Wkp6Vpdpeh8PmIDFR1xHDM1snmFPZH8DFfqSf0+ruqdbCGmvA1Oi0uuPQjh2Y
Kc8s0jGhXzbIWC0Khbj13M8WfXzkwpSxjdhT+jyL8Tm8R4YZhAOZCO21W7JRELH7
aQWRD23PPEyAl1xw776rPp4gAzUOgZGil9/chLLBqWLTn6r3Krn23c7ndKwcbzGQ
PXEiGlRJKcT83WsIYjqFqLZTdM++oV0smTUwbLsh/FmsZXe58ULYIioyzaj79kwq
SLsaegtt/YEDXARYuYPbaaRb0orERsdf++3NjIxsbwgJkC7/MZPGZ/duuF0iOefX
hIeXeF6Pz4ur7dewWdS9633l9ugPmNxesw7lTX2Ztg+/WL7CLA1syAcxZMl7/U4b
mMWoLEvz8ObaItUBr5HLu+jNos66CEMdgeeII3FHydX89BNJ6lAmMII8Cvcmf/Sj
pKQwPkeOCk523PSe3P1/2ATLzp8apOdXLYGm+XgePIePLvOMktKfkyzztzDvkwAb
uKoxtePV1RU783hFyBCHp/XJApSQUi4Hp2iNw8UEN+DYySPQq7Ae4/n/0bW4ovjO
EuZtHkxBdQksi0meuH5kJA1djDRoVppBO7S/57pb92Q/QskKOujIg2i5b9j/rSEw
R6kyP/dmAWok8HhZD1jNu/P/GlS8JoWxRJ3bIAy6BGrqNX/yIoAStxfQjYnyid7s
ZcKROqQe84v93azkIkULUv2GOlKKqFJJezT5bxQSRQmFOppf1jqBuuOjrlxZXDqB
BEIiHCJQ7qd0hlmmX3dI3k90Uu9AEU2hXrh2xfhoShtYEEMl3xpc7uWkHfDYaRM0
vRY+6SSjjiYXYYYqO8UFMxXUmXahg7WTKgKYk88qnvZYNRL4AWFz+BFggBGXrxmN
iWVjVK4uIexyOB5YTviHSvz+WUrJ6n0bK+a8OvGI6HRbempG3PdKK3CxhDiFXIxH
p7y1mxy/1T47QQqqjIe82IamtPNibmp6qXs7h8T/Mm/nJjSCnc1XncS0776pe99F
33GD4nA8asnjCBdaevXyDfawQINuJDSBxyvbASJR1j3+Nta0Hg167/ScTbFm7vLH
i27XPGW/eLJEwYKzFXJ1Yli3YW6Lt9IvCoAGBX6pEliGcddxBPukmm8hBQZkg+LA
TghHJydA8EO/1SOs3yMR0REJWXTLN7Ld76JXfCNI8uLfkYPovNwW7ouIklO6wA6B
Fp+DiUQHC6CD7U79/gRvr/sMcUHlWewL5l8yOfdvovelGBK7DemqxATdmZXtuBjN
iq1nWOdD9QQ4Hphhw3Avlv3QbzIdO+Vh8RhZKVvYyZrzD0LX8RorTkgNWs09pDie
gmkDz24ZMRDnUoiTrgCLxRyIJjV5Zp/IyJxHjbKoSDCT/Os5KCZRz4l3m/SNif6Z
ztZxEoeqCV3N8PTDbn5eS482gkbixoGRQFtIKBWiLze9swQIAZR+h2iNAcnVM1v/
5rlOkIKqTSXZ4PEnuYLo28WZowX5NgaoL+Sznz9Ey24zFYZRc7/PRulAIvxKZkqn
lWdYGNTEwFVFzBXyQmYY23B0rU0bIJzm1TDXinmePaC70TSw3xgEtCiAvXU3pFAR
gT9lYvURK58j8nWFiaJqTD1x5TIUkXv/Mv0VWv8qpOt3QN/AdYKMFzfd8qXxkKV4
iNcYNda5kNfo9Pcj7R4TcZPJ8sMhPhckPC6ysYOxbDdktmUdNIOXzfVOqNbaSDfe
8YmdgDIg/kVy4DIPaYhln5CFOyP9W8JxX66Dbd++PZhk7yjuDh/x4kfy1dNQsIYj
ErkOdtFEA+XVcmGSQlSyHZu/jbHyjTwtnImrhkTT8aG/vLTdf0/F88Y14a8/iv/9
sdbFTpc53vqfaOiocLCXt78/QNG6L1j6M7qrGwtTSM/+Dh1tUrxy477qzNDvdOYF
byRpsLSz4Qy38ElEaLeRQFCMA1x4vZP6yBHA+T4FDA5MqxpnqJ5a7S+Fm+8UGR6y
J8BEWFUtnuowlJ6pYn2TXGZnetyIIXJnKMDHHqUXhvGONY9gH0XacreVpQiEoYua
0NZmTaRwoWis/W9dEOwc4C2lTiZtWNYIYnKwVi5nREoa7OXeG/ylpLMeCl1fdX2n
iOaJdROCtWUW/0vdqkT8vf5SmuLB3Qu3qkLsKwuwYT+gajSsV7hlE4SRH8IHtwnR
lb+Fl0LP80dcQaZHWPgksFZtNZAhbIJx4MKSuNrpT4nDSYjLZzMR2hXS3s5BUyWP
AyWTbdlEzRtCxyWEzwE95ny6QNgU8atqmXd1O0KbS+nCdOU3NYybcokyC3HUfEyp
4iDxu8Wxp4CnOpUceuV4kIm+w1oOyKzcPhx/t4CDQrgPIoH+857ic0FzGE/LRY6v
zBsJxHC49BuSR8B8wFvFOIw47G39o2nFQVx/zvQreUue6LuXODYOE7Kf1As6uzJ6
49fBN5YGjUh108h//SbHAQSk+2WGeUo2iXiWMwHSB3wkYUqikxhZx+D6e+xhwGhn
YPR+dB3df78yRO5EAHy1My6WaJnf60yRlMlV+8EfNWmGhAceOi4NHE/7ez8Vt4F4
kATu482juRVf8rsA8LoM7HoZNFYl+Q+t5OZ2BgTNsgTmJvxFJPvvRGiGBkyg5+xu
GxRY6YkOVtoDmiBgwvAlc49bH+HueKoEz23qcVSt32i0OBGJ5jA4dn/pPqTFGeYS
MTTaa/qnDAvknoBtvyTgcwMnzM6+i541VKMMxyANaHAxfjAH7279m/YMQtj+YPfq
e41ARDOyjkua+ieabHNLEBSurFGZTLlOHPmkaGlchWmq9c8MkNJGYQRharFc7+Fg
Rg5rMO5ZHIgCehzSVRa2bPPOSHJCU3KxJrbEgY1PM9dc/vtoXjni5VfsG3Eq+KC1
llW39HqVUCxeMO5vDT72cmhX1Lpzq3x5rc4qE/WMtDJ5e8FZq/2PAULoYPLa/ble
f1xGY7jlBzZaTs5TM3qDXF9gEU8hhcdMgv4XtLj+nYUV3q8OyOqYHVEDKsVmnB8p
h9jueqPpnSIDWA0kkLcsg0sFGOEXc3eHdTYYRc4wcfJiMqlUD0twOkWWbVtLpAS0
AsQr3DyGwMF2EtoSb5fdenuB7tv0+QrxsMD+OuBFcToDvYCytjEsCtQEGhvRiQIm
FIhkAAPSfmBRowfN4cmBpcEK71qqOYUIx85k0XAQuSgPMt/kWpwfgGOsLluWRJVU
f5+xsoJOK2+zhu/y3OBZdkUjX0310BRyQQao94tWhb72nVwStXnTjUQ+vkGBfwfw
eO9o2TIT6ANxjLViwOPmHhhy+mVeIrx91ilOd/EEf1j/EoYZ7PYPv3dKLnBiF0Zk
yDDIvlqYWnyAoijtABBkJIC1kEDZK39fy74WghIEPmtPDv8dx5hfJw+ZiXF+apuv
y+9COAnuIngBPkUvbx+oi+2JwhzdgmakFdiPc1SD5n9guxYhu+6jVcmx3y2X1rj+
dOGdlAVwWqRzAXSNwPzz7ibSXx8Ge0lJL/T2xdE0QCnKBLitWFUNp0oGYIkXQ2bt
31CCxyrDeBhQYazYInE3k9W1CAtdI5N/Vht/aHR3aS62VXHhJBbQ7aGNfChw6iBj
+peQ/F2aVkKRSuJAq4OmTAMLYt7GedTN7JQZGiIkmmAfkEorOul2TC/l2V9Bg9uv
DpbPGbJXOMlrKZiy97W+QzDv+hgmqWaKBAIkIKd6e5lTAl+wsDIxQ4pscLz6xCf+
QeXlnwCGFnIT/1s4kzkYJxjgN7S/es/hXxhASaKip9WcCHPdV7GlOto6CSkSlv3y
h1U0nMC6yC/3k5DoGi5rUpE6U4lvi2+XFdItYsC7iF9pSGrbOaZMigTHrYbQtBCA
7wGV+xF6e8Zv3BCQXwHIpNfA83EtlEM8iVErmNJ8gVm0FFFD8LNsYV4oxVM7ZJ5z
mc2yOPslJJnLBSPKrz8GiSza5MlqvUSgEfu6CJ3qiQC0WYXe9vJNeHsHcBc2o6c0
rViINyh8kyGc9ymXk8AR8p/fARRwEtQFpBal9x9nK/RmtqPyHF2clsLFhnfwUy45
xcV/yX8ZUnaaY+QwpNNUCeZBOQPqEiV3pA61l1N8T7K7VxtaeTA3PAVBqpdJcphW
uRojEqJ2YsVMNikodI73DL9qW7eO4CSarTmeP7sB23KtGV0kPD3Z37O1hSPUCPUM
y6V7JnfJHzmm7GZ+TmKeLdLrK27N68kIXm8doIfxaT7u3/PCHFn1H5X6GEQ0RPZX
bcTEC7KkdGw2J3fZKfzP1MHvabSgaGAWDI+TMucl+kT/fa5uPCYNpzPJeY8/HYYp
vAeZSVx8bbMW4owLiEbmBvQ0CMNLOCSqQ171MpFpHdXUTKr6wVhJouwcQBlAi7xl
dSdQ2Vxnvl1blnzHRdO3rCaCCXLF+sp09hT46v9K+oGNdoXJq89/IsYqenAzOKMP
o7Cin8YwJQBsd/lqkzVkW/Zuey2EECb68yMoLGt4Qsgz1sZwcAjDw6w2ouiO1Fg6
B07NFQYmZXFFIxSlcg1rWx057uEQhnFeLs5weMYq75+BBeKA0IKwnEL7F07Jn45m
AnIT9jDawwnxch97gNNATKVLjHWIWKEleuky0dnn77ro3JNP7b8l33pqjKk3IeE9
xFJx5UlknnHefjAIt2PtUrCdy4Lx9rL+oIdFxW1oPDeTsIXxjpqMQHILLlo5FByt
ylY1xUdB3mYGgdREblA/aWK3luQylFrr2YLmEvxE+hp8aOZFZu31FIohJn6VMckL
CYVNjvTwtIQYjT5jHuNDAv4Z/+cCmAmQVq2r7QaWfv3wE/W5rOcN0OyHdklZjmwg
vDd4FDOT+l36NR4S02vP1EuocGXv+M0L2r5lxHC1BMx+ehemxEiz2SsxGBxdqnJv
iVUv6FLqpVunBZkR2TKc0bQxwz4za+dTzPkhABFqS7iYbDouIYB1CB7hZ/hd42Zt
kmlZOPypvxR4nsrbVAMo8vYALOMEqay0Mv1M35SaUIKQcCRHNwgN1ffUXm350E3k
zC1nltjYEYBZRzep6rInaEAekDaC6Wjg19rr+XTFpePZMvmcFrgnvgBJdf/rCyYh
wPuHZYlwK/UZZHKS+Ejz5AgUYS0AmFqL6iU0KYyjhOzwGcIi88bKGcMZI+5tGSiP
oFauwJBpYLqDY9kATUs8yUS6/nIVdXVm5S1UP+OxVUriaVscviYG0XmgO/xbC3c6
+bwRsuVdIEn24mBJjqMJgXP/O9lij5I2OPJxp0Xk3wmFtQIYraAxsgN2PahstaO7
RKwuvMalRCHznPB4jXYrS+6ACcZlCA4qSb0w/Du+ChyA261bTXkoKxqx5RSx8Hvz
RJ/W9SX23DbGTqg+ICoVaFjFxX2LHrFF6e06MBEQJfn/9qdVLAmIuVsY94CN5Ea6
5RTGl3nJ4nWjivge0E7Mz0eZIGG7F9EiZPbBlNxhrmED0lgCRnWjwIFtkKiyuiWg
TfHWOGfDxYmZw8A/a+pUEPgOgzgwiXEbbNHjRFOTb6bW1XsbfpLwP0Gktc4Rv1BG
E2h8HUGpsQmgfATDi8XnuwVEtLR12vV0kJXoT/xgpszI1iGDAYUf1/qhl9JwKbwv
rS6p/D7zFPoWHu77uWUbw+f7cATwnEuiNNcvAfM8U05nf9ZKKSESIjGmkfnCFI2Q
kx3Cfypa1jGaG3V/yUzXaplC6FFSyQ8i3dxhHG7K9CfPkU8JAbV6c+8sGlDctMgc
fZKT7C30Zaqxcv6TWaB0yBI5zyO1qvKH405uBwaCZkBQVIPnQWzKqB0cvC38xzmJ
8lYd0aF/8S8F1kRHoCzuu8lKUb1ch3PSLkbigUxYR5LISpp1SKvEMYJGNr/vd9uX
9iha5kTpaJAxs1dcCM32GkYIdecyW3lyA480Wh4Gc5ueEBhyPOvpGeFaLTm+6g+h
57TXW0V+WrbZl2Do2oUNbOXCyhiWNPl/Xqml+OjaM+BI6Qtmhz3Ydio5yy/1cHnk
Y5d0FhE/S8j0tS+XFQoy3owl+dPHhvFUg3Fmodf8bKcR3dkMJKIaDtXnW98ViZM3
2nIN1/QClHy3XNsjxgOg4ykV0zftRLZpzmz3Ye+e+jCJnC3ItMhDUy2E61QMeNsa
Lph3dWrh2cXt/vqE/PVJLRN7gbxwcIfvsBLjw0vXzueZ4PE/07UfJuw2Wf+MhsoD
W246XutIm2fiCwI+G+LB/knMm6sZOcKLBSJqvMC8sJ7L97nDNjyL4UXKBxQanF58
3xPk1VcKg0TOOW4yRizJmSlis5bXAkWstOMdSKGrVXuHQ2Mtmes8BZFElZXl5ugf
TevEglg3Z+wujdM9bVdpJVuVcQ4kVSlPRaEkDBtQ9mj9ih3GCVHrF4cupSc4jDjK
44MsH6FoH1XyHJq79RdLHixfFw/7uXJKuOk08EWZDfifVRTeAMx/oazDdCRzKHfi
xWDcHRRnpbXajOwqB9qmxQC8FJvLL7YzY14uNhJudY8Dp/jqeEXiRs2MZUam5Iwi
aHB7usf8yvhFEWy0ro+8N0/qnjNpAs4GpWqMGkJANe82fwDeZtxXt4UhgpaS7W1I
CIJOzRgSD1/+lUwpje7m3PRlkF2Bu12UfsjsCQxv3nANxWAygNgQIi96JRbEEH8P
+WEM2zROnynS56eQDvUW2Ppnl0iI6tFyx0L7u+EGXnS6NYXqJXGDS1PMW1lf4wGj
+kdIW9xyxICF7DmppM7eSwWN6lbCbaY6GfOIiBx5CxTnwkdu7uU3YP5qfm3sk7W9
wnmYjjcJHXIKFoK2wrhxINSA3Ww5NAiEvA7yeMiqAVPwj48YNjfTBkjAwbyibNDK
Oy7GO7cQ2XEFTIua/UJ2jV3kcdLS29YMFvwy+c/vlaNeLTiFsOXfs/0ytHgqCd2G
JIlmFjce6nIsWePfZx74wx3BAoq/KYWqbEG8xHMhXVmYxkh5G8A2p/Tw8yPz8KDe
rlMjsUitlulw2R7A9d0sEAAw2c3bpdy5+JJApUrlMeubcAzIxbFR5/V7U/CHFPrV
w7ducT1tg9u19ACjEPJ66c4UljK7mM9gJvMvLfXQFtp/bKt1hYHhdRw3B1YE/xtF
wf5W1xyjc2Z5gxTGimnsdq/EtOnhKUQmYLLUQ1qmj2Ksil0DKtzQALzl8GWZM8Nc
X53a5b1acW1tBX3SjE7uy46uLP1ID6yUaa5cyQ5xSzz4WQ8C0gZmZZk16OOIAbk0
vWGtTwsHFCfMqFUIGy2TVgBbS6pUovZf8u3arw3b4tzPKJbIpepq8nW6JUwacJmP
XTs5J0soHMA+W3hG7w57vBU/rDhUo//AtbjljBykEYbTtkLoLPu7rv5SUdJDzCl2
+o68wTL0j+JlWlNNAN2ciBqqM/GRqizKIHpJsJMDAMR7Iig1H6+o7wv1Tc8Pp44+
MEtR7aVWO8Mzc9jwnICX/8pNdCklk99JFsYKzbRkxAHbmvKCSaMHE1ToTB9Yq5SG
U07WwNSxLSgUa6sc51ZQtKuoo5eCsXsNbc55V09JfZjc5CxJ17qVhieRWkrPsPDc
fjVADENWqxWjcQqkbEC77Lf5nYBhEA5FCA4z5y4DBcNQE5Yi5FDPPO2K2ddHPVGm
U5ymJCjMGMOvpUuH+Smov3AZY63TEzJH6Q1OlrXNZFpTnFcsj2PVMlLXfq81k0RE
8nIixOkekTVueCfn79GfpJGq90E/ZBvtE6en7Vqz0F/DYOoBRyZldr4EzMlFosqY
H9429ElPwmQ2lPPEZpSdZdpk3jS2l3XhQqZU+iOK3v7caVyk4/h9a07BvOkmS8wO
S+NJsEUs/GFrbTqNh6Z4d+qUvK2A7Ufzxyl2JUrZzJEzCv28tnYP0Z9vJ+IR3Zu0
yUYISJAZeJ9FFkx6GlsP04vPk099UsJol1B8ht9bFtrhwevGmhK9Ba6PPeUZ3VHQ
0UvAVNt4cHV62kY4qBw+VLzGhJ1LeoSFlpvWFKNcPcMb0r9l5+ku4Bl9F+dj3DLD
/0Gnh1nhtyKocCJlNdGTEekzdix/VForIOKqI0FCQjJqYapkkzPbGGitt4ZZpGjH
CwrsuGdMGg4OSEHRgEHmCnCSejdFesOb2QRcu0cwaBoxtSOqhDwAFy/5phx7hXPP
pJjNWJ/pnwm/8APMyol6wWdr+polPn/Sj8FQ/+Vg8iMYFyNrh2hAZYZ4JTgIRuDB
BjGa6fl8VnBlAKVWlCoRS/apanf8Ykezcn46Zt46IZIrDFTQFe+W0gD3f1AANrJY
Dz12g5rOVzsMpBVuPZajhNoL+nXTvDUN1GuEgab8psdmTK7f9i79LQ7RmibPRWe0
0LGCIzztwqTCXNZEdzNE8W8aVxh78b0BLvasV/cJkzJR17VqFIDc3YGhf9fhIWRw
lemba1qNCBb2PeH0cHZEJvb9fvPo3fh0Ig35qgWZi0ad+l74GXQfIG13Myc/NQRP
04NyjDJnpOXu/TdM2JC+lRmdqVy35XLyuyZqByRPmm0YHkp/f4X2RDbLKYMH/mku
1kZR6WAPym7wKrgbgM0JkxwsoKiNe2wX2f7/NFSFr+KjeS9rMD1uix5ZNRIVKUdS
pfIv8YP51OeTrqYD5y6z6/KxGbZeiiqB0DwbkVBDvbb7KbtRlpcCekftmjvH6Oa1
/trschxNlR/7u4XWn417xw8abi7RIVVkdj075voOYv/Pp8+HeZQSaV0v/YXHSjnj
H9fCsnZAyEaOw0g4yKaYa8wvu3tRCU8WjtTKgLcCATb4c2OZ4ub1RIyCzrmcwgBm
1bEaNEB+AIWzVrs6ChUbnFIQizYx/8LPLYsMhJbtaL1J3USC3f6tO9xZK6akbVyN
l1BVJ0zAorWQYBC/w/qT8ntcVIx27U3Gyb+jR6x7no0Huvs65xhduXxvzbqTXdTN
ckRgtOKedlh+p67cudomRXsZOYj0bIGULdpgfPqg8UBoJgfjwQWTtGwafnh/Jpu+
PdHe9a+Fzyct+1VYdLxnP+l2exIytNyMO4kXnmtjdp/WuX+YgjC+jbHFtHao/PD8
Mbn+nT0XMPbGvUNppjZ2oOu4fGGun4FTm+HOJr3Mc/ylmFJbO2F+AwSsVW31qHPC
2rBoBy/TAGXSOfOFuuMR50OVEaOG9+czw/tt4cqJGwN0SX5r7DnL2EYwm9pA96TH
IfhXfKKh3/ixZUC65ed1zgIaLgDSnfVwC7Ud7/lq8oZVvwjW4SyhaAgbkqwDejfr
ATEd+SxvW+LTDo+U5UCfMRUroJ2l4ilZrGkrnmi3rhlyHYq80nMEjd5oGgWcX9Uw
sPnS8c/Zy1dk8xYHqr1eShvY4yddSJVPSgU10ygPHDe/cFLL1FHR+sDa+Wr0Yivn
2B/+6GMK1oGJyQTJlaahKxEbkUEDRKWNJ+HdtYLVIA3tDdtJ3sKm3FAGaFGB8jv8
/3fcpg+9IFHrzty+GLYv6Yhqg/CuIbYDeN6xaNfN+jl/1oZ7Gacxzg6LXdZ6Mtm+
xpPHzfb3hlkkzwfEmY2rkmcqROOfAYUOjrDOgf98CTS6kSXG4t4mSFO0ZM1wAqje
6vgcQB15Kn9JZzTdcLwlbavuD+RhIttzq+sIutLnjbJWrEiRYvJwjj1PT1H+drWx
G3GAylX2cR+bnD0FI3AnxgXk1fuZNZqFJhBbFOe1I+AyTTC8KQZ0tAcU6nGULZcu
6AyMjrokGw08VuNdF6V8jrVPZ3gb19zMiAfrI570l/TJL4dV46tF+T6EPiLvvq/D
cS/PVqZOSnot5ozoucIn347rwGTxCCcOHC52ih6WgbIq03IajKbe6QVKfnEHzSTj
OcR2EQS7ObSCJTd2NE6rPKr/cJxnJ2nBG7dp/ZQ1B4S4URL4tSdWvu18X+/jbW4i
eZYhCda+u1rgeB054ODqPXvDBkHUL7WiP4c+BoiYQG+57vZmBf0PCgK1hocaTNBE
GztLUnzDSOudhT3wTLqsHCyaq0Isa8siMzFpf4u3OXQmaoUMoGDdppiCZW5Qbnho
Eec3D5YZSh8uFy3yXjFCRJPV8c7sfcAZ/PKSlURszRQGgejBy7wqrTiRdDGmAQD2
5uhCKucuXJGSpzpZYgtuKmfTtRNuMxQl6CNtE4ABzMx4Y/Jl1U/PHPpX+KWJpYT7
IhEj2yCQmCYFc+IAJisE3GnXlTVj+KgGbf5TuAFtxOVFd9rXK9GDyGSSbYuW78v4
jvZ7w5gzCCD5PJ/4FG7Ks/wtWak0aiGKozZzbsViqp6RNeJCFQX8qrl9BgBeeiGa
QN1als7vPwgLU55f32BaC5u9YlBnFLHHbcWuG6mdwRFw+x037rTR+nuXCNcoGsSM
jVdPCetM7BSZVZYTcezhXwU8wumYFIaoVolMnUWPAVyqJKezw2UGNfs5tIz0OdeU
tggVjtDTN3MwfPuqPrTG9ZtJwem7hZWwEl7Wq6CLiFOqGhWMz2RRsSroyR+q9bRn
iQ1SVFOTEnDZ+JKR1yA3KPpTESseZqvEhIsbVHD7j+waEas6EL/y8Lp29Itc6Vvn
vL4W9ZVg7/98M+TJeh+zXsxY6ZPkXW+De3Dv9mpiCrk2LJm2LCUpZM7fUTnmKcbV
dAbZUHGc/+nVoEP6Tzpb3DCgHy07ABKgylRJ3iSA+EeGlmMRmnOHtn41aZPFZU7v
gaiXnmA0r6mwNScHDUO4whQawot17BfIkxfq9YhdiNZaVTqqqZhiW7uukGpV9l5L
Ep6qcVM+V2pmqnoJtbNlriXscwtKvd9GnzjqaUAjik3dOLYf3o6KEYx4v/otyVCr
5eJ5oGMVrETaQwJ00wjct39asxOKhaTz67cDuJolqtWIBhyCe8VhBI+qJptwO5yC
hToIlEpT8TzsxcH7PPaB0XLEmy7DvoyFLj3PdzcZ6j3Gi8FY3v4aQXMCUeskf7eS
kQvMuOIIKpcWisDpt4ok0fnzyhNG19DcwHVoB/TDB4Vcl8vk6ujDqpc3s8Rps+xq
3cQb5yPvTzJDy7LRgoiSMayIfLt/1o9RZ42G5fb2JoAypAh9f+0h00dkQd0zcZGi
ma0zqLEHPJzBKt5DHIFrhQPvutdUoYqlTRM9hX0BnMOhfN8Wm6j2USuIam50WqTj
sWIVOZmyNQAvvRdZWhvs3FDwswenInre5Hgv27e7icD+as0xyh//Pkogsqd4/KMd
c31oAx6oeSUttZ/MHG/PRUucs4B4anDhe2crDHTBNT4nn0+w9yBKTGmiZxAcLu6K
BHLeKoTfWcy0J0+0rDtAQGPogI6h60AUGkQMhgki9ua/p+yxxULPix9e53AC+YcD
lpRbV6NRq/MNY/vy75CNjrYqWMBwMoyO56CsAirSKgWeISqyyRIW6ZGTKxyYrtzH
M9S759d9EekVIwk2kvzHK7owO4qj7tIovC3kc5mwNUfKNaFEKbEMf/WgV2CpoxW9
vsOyfSu62mBBRNgaBvkN2pSssoWIdLOfCPs/ekIN9A13vSkDGHIrCsDpQBaoN3b0
sfE1nk2dn79s/Y4xTPSb5LuBdMy85NtM6g47bjRX4fgDHr6AzN9sx2dlVCL3EE7l
tycDdCTI6uUJPl25zASn2OAbSTyMEUV8XVZz5r1FOex3q6ALsOAuojamE/8+LZtR
TY3GnG+26k2Vm6sPyTqWHxd3ZQXPd23dJ3jfs+wnKhRyyqE547rnfuw8D0686AhY
PTVsM6M0eryKotISJJpURBKtoN70Xs09T8MkKA1QRpOOuc1IclzA5nVkwn5rVLsK
wqnQCgBdwu+5zS4vCn3CbhR1L3iXZrQEn9+RrS1I8RxGe2jvRE6+RqUMSCqHYsDm
Ifa3oFcCY7XrsPdRd39erCF+HAMnpDxvp7nJKqHO8eg+y/WjCSiKPjiaKaEH98+3
DvSLt8jg4g/JeZmttaoQtYxWbltzsDSEzVouVwMKB0laCscxCxkCYwpRgXcCxCRV
DO0/zYsQ/OCyp++XWFgLTCGOrxXqZiESoDzgm8Z48Y21iFErDaTb+lBJZGUBtYSY
QB0VM3It0uj+QNt2adk+AlDur8tL5fGKALQvRT5vLqqWRNxJ9uOCgyCqAP0pdg9F
VOc+WTcZBaaiADEMuZdSnoK3+QQ9sZtINuJxFa3Xd0CRSneSWiKrgUe95fNZjcLB
RWlltVXe1K/Ei5u/EPHRswKGSycMD7fY10h2zyk1XsieRXHgmPdgodncBGdIk1RS
oMHwGr1bHH1RDxpzRUgotlxNd4OVuvEifBTaEmXnuUb6sr6PYDodb+wDHUn/Iwo2
QisT4T12nt2X2W76NCcOzXyeaNJbNxD+wKstIne9X/+V2gTdHPnOtuK1+qAbYqPj
HiCDVe+JWJs50WQ/tb15NNDUx9MbLksKiAzydAGxnt1PrA1vO6aDN8otMcQGW1qu
DZUPrN9JL/UDxZhBO6JZ7W/xhGwawt4uNMn805ZcQOtkNRjbqe6YkW/4FXisuONd
RuZRVP9YeoOwTrU69FVnFCLO+7+Iae2iVj00OgxHXxD99LxzxXstEhQDe2KBxhNh
GXMoKtSW3fJcbglyzorfKZF59fNWFkTsURgXWDXU8Og=

`pragma protect end_protected
