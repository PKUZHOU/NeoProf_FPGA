// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
et5ofVK9BvZQ8QseJVOLtYfOWj0Y2cJaEv2WPXmeb71WIJRLlvSom1jmhFnU
pyKl+1RLcBzNB+RlhRLNkL1OlVlAoExlccgqHxFD8hLE1DibBYevw0NxaYMP
qQHm5HFD39CUhwekRa52Nr2Ci+lyscU9keFZmn2miSIvly1RLluM9TSUDQ87
gmvSZi+V6hXqPBLnRNk7Dn1dNLCNRXcT/l0az7kk3aai9xLOu1VxaYLEz3Qu
gGQgP7cZsawNV21Lfef+Wb18/8hb6UiArNKfNe9xY46gerUIMXISl0tKmgDY
ZPwod8svBqCqtyjhaKJPXPXcBqLoj3vs9PLnnt5tZg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
jhdpgBWTE1huf17NtZFldIEQRdabjzQH7FFvKWx8uGY3xc4ot/sX8ne6PAsB
/jb14tGM4A7iHmt+R6HpEoeCTNESXERxjRJ1KMmA8jSeafAOGlD7V7lwDZlC
Qt8OLzf8kz74Vu7lJsW4g44UgUrFXnpB8WAfSuDmSmAhGCzB3JQU4yAUP/Jj
NDgXNOYhvAgAtg4XvNyV5Yjq1oDqEiySDJKq1uHZi1v4DLOacZgV5lGLBKtd
CnAQldsLSfeb5oZCzbMFM0x/XPPzX2WOzrBB76GYqHtjyyuv8UGWJEUjpEbC
oJwIeuLWUp850ULqWla2yhBelAQzt2qZ3X0gLBD8Pw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
OHXrHBTM7vsFbnao70vcqe1G3NAcimyW/R70TH9gzdUmnghsEA7jDeYLH1H8
HBJ3a4vGHbQ2slyRtkxpML+ca+4VP/caQuz/slvP1VHkcXdx8oi8EuqS5WyM
kX6zE1OnMcxnvS+ug5QwiNmfIDP9CXGEh1KCidiX/Nd5hDspvEyw1qbcHQAH
PFHUeam42rNqfx9iQ3HZiPFdL5wxWGjuxLpnD/hl5e4GRzrKiSlP612MQSrp
CWLiKXoX3rehxWRIxZlhr2pe/BQGd5dqri8TzCuFbYioRSHesIdIJt284T8+
1dg5fCemsOLWkxMgW+YXIpMHQBGd68Ce60us8MBOow==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
jTATTuj47eGDuqAeneIqgJXhrOYc3pIYxAqpRxp/Ij+BaamfmzeaP4Fpwnal
DHPruFu/0siHA/6X40m1y9IX6I8voU2Vhoz1kwOn6FnrvGpP7+/u9I13AX4c
zT6anILbAdFlvT0g4xYQHekXOd4zNV+ADFEiFerNweZ2cYLHRf0=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
VZD2twd5P9VLk2vstS0j5absktTmwIqHoyAHGLxRlHhjsBoeudBiMAlGENsn
LuDD6RTHKUn/tTkdR5fR8uHgBdEN3cdtgXh/PdqscqOstp8/WipPG5FAE7Yv
L2yQ1BU/Hes/kr/VYfBudbwCpykwwX3Yo4Xy/rDIg4wiVS8mADsHLrIvLn4L
EF+5IRGvGGeCF+aw++pxRidcTnAl/lwitz9DV8rd6bB6cHdBaOBvnc1a7c0S
JnXPGWrvMyiYj2jP1cNPA9gKFF1Y8wfmOsvCXc/gOr0kIXbS/ep7s8ZWXuXm
/8mnf7StERlazDkcJ0cRUYf3EZeY8nUkoLh85JfKB4IZvGHot/M9krgmYqND
P0RuKCUureLY/ZSByqoK5LRiV4HeiiPVkKHcX2fGKJWnTc536Ra7oKOoFNmj
O412HRkwnP5xoDSrEGYX03s0t5j2PYVds2Pg5Gjg8Oo2hFY7YPKoVhukNqFJ
7q53Vpcwi6xAztJVBddZsPbnPSY9QgGq


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
s+QLc0EJaQyWql9VWlmGsor5VmpsUALSo8CjkJUB2Xmlg+5SYecr8EqHAYzG
e53acRpE0YyzRWiaDgC/E5i8npjjAY1j0ra29qMQGO7VbjP21QUrEUGPAkRI
ux8UQemzcewTNTmvVCJcDZX0s8xpYTib08yvJ9l9K09XSNotKXM=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
LP7ROUwgQiBFifOERL3YLGy6inhZxN6HZ5Pn1P7SLxq4qOZhuU0kRjnMtlO3
d44uA4gOdbiR+ZeOJJ1DJqaD9Yy+o9O/shOUbdpoYAze30X6JqowY1scZpDA
jSKmxDidJt1zEZofBf8In2Nq4ma5mU6Md7euHKfdxvSv7JjS2ag=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 329728)
`pragma protect data_block
RJKID3pLkBZoea6ORVoGpfCMM0C6Zr1mD4RcfAm9dPJTQ+C37t7DATY99gLY
ZxfnT09PDRp/63vGlvufWdSa5VhMMz04/32DnozjsRc6GGF3BARef3x/aQft
8v+jOCcP5bHr9w8DbZM9eR9+o/zfvSgAtgAAhXN1vxnyyH/h5OtGwbbvgAy6
uKhHHsNCnAbm11T/wj0dw1RkA2LJYh2sOEnOfsy8hnd0OqqmZhXBfyyjDWFP
mVP8QJLuxkPIkRJX0g9vyfBfLouY/K10W5jZUy0fFckQCLdmix+WHLelv0Xb
eRO23MqmW2jdf7f8k6Kq/6Rd+WytZv1CWBMTOD3B5kCL2HAitH1OTaOYNovM
VUn2bRhDFYal4f+buRA5fpUbd0g3BQbHd2yUYwqzHsWMyTgsM9wZXHX+MlY9
ZekGS0fZIZtwpbzxUpIwO9oG3hVI/xvT1YUPV+M+a5p60UrxtG7O0cOHu/G6
VZbdV5OpzFL5AEmxS6gAJ5ZoRy0IreeIzTYtTEm6BDITf9DEqMjAaOhKYcjm
xD0kLBTj6MoLRG+VijecBbtq42GhnaYg4l3FGqLxYTnV2dxx8mAyqpA0UWQw
drL+udstmcYBxspkeDjxF3g2ETsORgTmeDi5N6xlxF5dCm8k8WoEa0/REL9W
78pswv4NDSph7mZPxmve94BadK8iC1SwUuhA5kG6bpL0VxoFHG5YTUUf/qlx
WUg77C6XqoT7zQi8tM1bTvgU6r+YnuimYeOawiesHkuCcwKkGrpggTOlZT75
fwxf9ticExntnhqY7mWvfWN4NZN2Vbj7Jxc8AWVHjmUi0OovDsNO1Eo/rDHk
EiAZP8d/BRbrzbWwfLuh8SGZZUoNGH6dE4f0pz95lX3uen9CvBg/b8WUilhA
vhJqU3b2ViJypTFniPOOy6gv8bKAqIb0M61Id1vdGCDorWkEhC7OrxW3JRHB
XhHAGuDYOqt0ZU6JF/vrMdQmTxfGuCso+TJazGjd3hzVkn3ccIXhXKrZbLvA
Ma/qc1PXHUGDBmy33aZ3MswEdr1qPRnwH83r3IB30zmpRH3WB52Hh+9Nd5pB
PvqC3Pw3OGm0HmG1mViyUt/MrP6xl/izd3O5yLIs3nCB8/KL2zWLbZvCQSov
vsW8eicYNRwmlAnVC/0kjPYcPZgTAdSlh8qkBRaVHxr9kQUfElMgu3fW+NYS
C7bLB7TleVUMl6SdnzmH17t3Y0y4WHdj168ChAPD4VrM/ZEu7Nx4LBbTFKuO
C35l6UHohhWJK8mFhDvDEpWk/D5Q6W94sEoz8X8sFPVhtMuKFWl+CHDSi9VQ
FNsKhCVg/RIvfjwQ4/ApVdtsOK0wvSZ7UPbYi9UgAbPCozsxkM2KE1WQOBds
dlj83DMDbfTizE83QkxjEh1YUgVVN11kEhgof7OU+AChHJvOqQs8e6zISRG0
e8++7VcokO0QwamvG/nF5OnWm72lNCryCoJfME415SkX33yn3+OBoGpptexl
FXOoLfQhP6yGn0bqCxHJWNeK7ohaJOF3St6B40oape1NlJHTGcjur7Ztetan
sUkSSe09NSMFkhfKNAWah4gmFIN77FDLl9Fd3j1btAsWg4m+Z/7gE3JyFadI
yBlnUp+RqOOsiMGyDTXz9JIHRIwph4KavjxnRS0GhnRdcnQmHNj2KOULtsGq
R1KbcEVZ1qLr6yEHPaYD+H+CUftPNaNL9avImt/vOfg5xJGl0FSSOQKIBzbB
KoGYQwNI1L/8to1C0wdiim+Q7RtdoSqW4tz5NdSq6fwpxpvJA3ojmMRF/zDy
7vsWjjzP4mU5TzSh9DIqr6Km6AAs/wPini6azXgigSjGYNqctqa2cUuQzLd/
4FpdsDLwa1iTcHfseYvmIYHVVdz/sJUkSYTASIUtBL9OIob1oH5t/e/94XaV
wg6Li8L8QRYbw1ystBvy4bQgbehv8NJ83QTdIQrEvUpECfWvLOmudFC/fFEr
cevWQHbAx10gL4INvhLj9WYzemuY25UJ/ckX7q0KY0TCz1mI5buOtlnJSh9M
sguSitYGBnelAHbn6OwxwR9ZvqF7E4Q/zLGAfpWEL1U+Zp26PfDL4Ae44wRC
2RmI+SX5P5WnIZdHEJRgU0x+0fr/3BvfYh8Gab9zkR7Ut5LXt75SDgGPG445
Ex/8ddTFitEkudwJzSrmninngKYdxobL6JXOsiPb7JoKPothkGuHew/tGaBw
0D8w97eenVLAl/6IHEKzJ5Tts/fY/PHaseHwL0Pnph/w20kvjy7tfbCl7A8T
LXSVtoU3NsYUPbV7l2O+dDcraMqIb4CrIQBpE6slpkXsv1ndmpUc6+0wK0jc
i3L76o60tpjB6jmrB6QTEawkYLQdH0VOw4NK2tQ4mbb++6hmROBatzuJq8Ge
1LxpknqWHCjFcvkXIjY6ZwrgP4bTOMyrA3X9Vq6h81NVNEgRBsru78KLMJHg
C3je8056Q+4YVdOURyOOrSALcxP0h73mwubVBNzJ353zuQdBICNRuSeM8vzp
/WEzGFgfG1kzRRoVFlvj3RScxn5YLUIFdPZ8Ne9Cfj0lu9I5W25Pt4tujAXn
yMulbItjIjjQGpol5UA9Suvl9lgdMdlk0lcHg093LRIjn0bK5c9uSzSI8jjF
k2AmSRTmh3KtUCKCa7i71B2Ave75m2Da5Bq1eO6YG64k+zVjQHylaGyE7bhg
2kquGuWMzyH6eCRakhdGiCi6xsxPXREQyvDrhPtXnIyUff1wq90aKTMtmXEA
ZyJQ8Wx9q/vkfZf0CDM20+w7JdGI/CPUQRTN3ysg4J6GaDcEYTiKIXSGlaY9
4Ev7nxv5+wOPMkAZWtHoTofziKIyMcFXe5xF8JJA4CgooYjzyW/BJ9jalWBO
3u5xKLKsLL71KgOPpqAXD3mXSrf76ePpJxeCYtSyXa2A9uAIVLjz9csvcd4M
KVkMINK7bVV5f0vV2mTHZPUEkqlaFphX8AOr1hloQS/W+FukNIqDgJbKtBXQ
pmgjsARyi2vyPltupXgHtje7O/sFATpHonXKhl7+zjthtNMcQKxVgv8eU/Dk
tNZ0VFTB7EDN8qxrfMPsQl45wM9rfKlUPbf03ct3UdbGokKayU09UoHIruxQ
RPIOR54x/9N8B8JZ7WnwNJ5JBLWQ5TtMfyzXZ0WcW/aYbw/2sqZYA367mucH
Y8fDtGeUcq3wxX8omjV8JyTYtEhjyvlpi9yrPHWooqwSwWUklbmTNorKQMB1
S98B6C9nsv47TO2xbtOBIlDNnJkHMKoCwgS8EYp+H88X4/viaellbzLXW9oY
l/vtWL9DBjCeJ75uHk7we/aVQZd5e3ha7aFK4OOWaZ5eNDmjm2ro2AxEo76r
XZoLiarf3qK/Hk2BXB+LGi712M8ovxeYonOzncPKUDz8WsbqAjcwl55JCzE9
OuluD4oAXYovTcFwfKqQw5gEo+ZnNn5ZEYQuRnf5gWqFrZ0TwOWZLlpnbD8v
fQvWq4I5kJCFxjN8XSnu3oyzl/dhzy+Jg2wqVSXohPo6fuMgp7g8/43LUsrh
ZgdBSjZniV8DojnYXTaUc4wyGXrCQ2bfH/Yfi4cR7Bcetl8/KQQLuGGxkdBT
KUVwbE7AeQOZy/Z9JUSCFKCyMWarG3gEsniI1HmGCZJ18yTxnFeVJkwWn3NI
7slIsZzJu0Q/nYBucHLoiFD7Y7Aa7MLBOZhm/Fj2jaMmMwqsTDNsaunzzxkz
YX/3QkoNbuhNDxu/XBGonkxBargns0Xfahpwz0XhYHLgrPFeCyJHWZpiHG8b
uAGafJoKQFHH/GUzm4sW/KxZFILjE9MQ8XppjdB8ciHChJz9YAJO2zIMfa5I
HVo+TGIkyKKFAbKCVC2AIUREashRVImuUr39F7Kx02CjoeOr3VDjpSpp2pv5
4mqJ4h087uxR1coIGCGAHDVZemud9fiOwLFa3otCwlnvASOmPwrr0T5acV8R
8Y8J/ekHLC3hb/11jLitBnCbGiaOCEo+0aqsHI8zB1otjHVw3DqXg3qjiJ+0
z3s5xKf+/hXP0n2qhlkXGhgNxIscGen5MJmrhgmvvYROjiz87UytRADxVTBd
x1OPgjejc7SpQs/vteMkISpCRnW5tABtRiHnZPanSPH7/NfQPXOpyTfX0C16
hKeHJMNRO6EGPDFwxJlAZRy5lGesEu3QyH4UUOwu9rgziM0pekGqR0rNSItj
aSyu/BvALpjZlCwp0aUdUM1GvoeBbCBbjX/LYzuFeVjS6fex1dFtTQS6wKhK
QEzPjXQqIv3GKYw+jOjSUvrXyG+5plzoANwYFR+HZI498G+ECk2tUjua0L0F
8IB1VvGESHdyhrWi9htHusC2vCT2vNO+Ow/v0Gxe9umzrU1h5/JtHbzWJfvh
YoGxtft2Y+z5FTDC6fKSrJjGnlCW5IcC+Jh4SmSAfL9+72i9PBbva8hoW1tb
7SeZJzDZxGNDtwBmAi1pcSuczJ5Y/dqwFb1x5s5m0hie2JdSwLD+CiCslgPy
13RKwnm990S7KqX7XKdUgkZsoijeB3twsq2wsn1vV4t4Yy4P3AIJ3Di+PDv0
cwb1sDr7fWm0jN3H2LDz9h3TEo74kzfxqWhj0+AQGy+G/zKoMU3/UZLX5WKP
Wpd6m+Yko8yUMJhQGSvUejxsoug+UXoAd5RgGuBFbIrcFxBv8gg4+i9lhMnG
wkLXDNG3lyChs6THhIBWJvl8rwf+x34RkdY+/k6qXJ3tBK7oqW872u/w8N16
XAqf2X1BMkw5EaKyy8yNs1h+kykS9qb1lgI9unTTIynaYQtX69aPraWR9U4B
JfwYCBUonk2MFLvBs10XJ3P8F5aucYO/DFj6+EjS2aKZofB/shZBJB+6Z8sV
z9r4P3Y+dF5sivu0Ua1pnE8B2faDF9AElgGTE9RpposMezWKs4VjmoVnr/Oj
NWXRsYwYtioZpKybK1Xol/EJ4S1KFKE5gubtL8bUDduOfrxDbfVwOlLrFbzy
mb38lkgJ87LorxOCNDhFEoSD35ZwcvOVvkAvpUOPW0oxVny7pa4ReQDXjpIu
kC6oyP2pRNyafbVFrv2q5Bl8nPEbMRAkPdKITwb3TUkuoG8UEonMMvOFnnU0
GCqfsDg2sJvmrK2mGUf1QSPWiFTQiparPsggrrlSq+6a7WNPHp5IWJ3fVLOJ
ISkHV1dD6BWlwu7G4HdGxGiA0/q/VgQWf7YGWGqYaorvipwS7T8ZXdrVmgnT
yJHHKFooE+xvw6b9KqWuF1uprc1Gf4g+VRhVD+4b/8OWnNK1guEsziXl38f/
K2ds1oKZT9uyMJa6LFgnbctvU4BRvUbYV0GKNNLtzytLKbI7kS4Qa1SlEHc2
8vncpcXr5HoIHmy6SlDVsJET9gvbb5xLTAxiiYgwAxLHo+jq6BNZ+JkKZrbC
Ngzp173bLbUFSJO32ThJVpaAVvOmRaEqhLM34JJjq7p/dyXQTJUjMnaY6HRJ
7JonMWDk+0jClehEQVqJY2uPirBPhS+ulLjtvniSrjjw2bU4zLTyTQpMHZ+Y
VvVDVoeY6LWVyprT0FSqmV3jU1GeR9oHiIeZcv1j9ChxEw+YQ9JIcPLAsrhT
7pIrXai/MOHqUNk/aHEW/tmU+tnLGg7q8P8AWC/fZbRp0Iy6b0Du4ylzDOLv
Q7eqFcnGC51RUZvHIxJUace2mpoRyilO+vk5DjlpLuNjIBu7bJy8cBurmxxv
GQXbcgOPmKYY46aaOGj9YeKaGpgig7WPJEMIhgn5nFJIbUcDCiIubhUHdwWF
0lGvmSCSyT9Kac3KIyrX+2mwVjtVDBfGq+UGHyqhreF0oVOfNgPU2sWNVS0E
b6ha59nxpUiEoYah388oC/XOwCcy3TAKAxjbIYhgCE2p0eQCjmhQzbdS7Cel
msIFfOjwYCfC/3th47ZPs6lkiHULUdh23xQwWRmZ36VXQEwUWzjmiIyfwV62
YNacpbJ/THiniCnyWiKp1rCREjCcwYcKjl8kmd2hUKiaepI0vFs0tCXNha6l
719Sfi4pcS3zeoSE0OBPU2UElnvuFZGCkglIU+BjoFheT1O8NRaUKZQXwXdr
oXIY7ewnbffd5Z5THQex+/2cbtjEi9DPwwgdCC8IXzNUSpmCSA5+r1nmjNVZ
b9NWOavewHz3P7ss4XRXzuyFHSptG+jAvea/xZH2VzgXY+9nBoalEUcAMB4q
HIM1p5KINY+lbgd41nUkjahvpM/byRsXNXaf9PORfugKjwu6vN6ytjq40IV+
cU9sjwtEA5yVyiF9NbNz20ZsW4ad38Cr0UbYoPrtu/+rI4aZV3jry5mjYnhv
HjCfK4Mv3cDKJh3RNAceAOj+COzubCLKY6xyNePU+R0d/mrQCNrP++C8SC3Q
3Cl6l4FVlQ1zxX7Qb2rJ5l0pWQWkVD+vNQdXZG6VMtswhbFpXRYoHq9Z5CTN
jxrKaIez/mcd8/qkqVwov1Dh/lztdqmyBhRiROdMoUxT5IbFhRjz3he5pS1J
uPwycq9RAyf/YIphzcITq6GM+KFnQJAxweI1VAwkr/3U3TlYwG89ajhQqA0I
T/vZDeBHsii/Q8NLEJd0Ka+eFmUukYv41f9NOrM3dNf8Do+572ynbcWG6Isa
YVHlwIr29XEvQggYhzwV+YYK1sTA249WOPI/C6F5eTZ7bSejCOTXxEZTg1N6
RTPfFsL7jo5OLfQZZj4g++ojBZUzEkGsqGeXWXcSAK4lW3BmNOBQlz9UDgxS
rFovhrL7Z/+OhuNA+82Fvm6qquqacvVUK9RyNMy7D4jghz1wrgYt3WmdFxqD
fwjdrE4B251tuFaB6O7L+cIdf9OKVK5zayP5I+caQsV7IIULHR1edvekSTKO
OfdcifOUY4d/IFgZhYYt+QK3VV7gMcea+atVPilHkP8FSpQzsxqr00UkRxwE
0Nv71bcTFlOKMf2EaWd89Pj+WVj3lw3PNDNwgHvLUCt6H5sDIHaMe5i/EFX5
VYXQWaba/jiMlWdRV30o9mjTjVC7Hka2zo0dkSGM5KZ5jekH3aLdVLlcNtPq
Arc+w4NvNdauSYa6dUsRBeNbmSKtaJx79F3gROgUO7vWrn8OcC4NKeehtEBe
Cxx6/rIvaoOVKxprXQa4KmdtVuL84nSya0djWFUKY8b1Hnm7U5BfwtB8BjcL
vLzkbQhuDXvI0X/CWlMs//rOGtsTPz+FVpje1Ep6S6UX0FjOswkefGdyChfZ
YUY6SwGMeNR7hc0kbK31LVerGCpSUbjOpCtW1H3vifj5xqIpNIKNpSkSa4ZK
MNm/6WKuxSvVsS1x9lUfh0YZ/3FNk6jBEiA3ZDbCalPFqjEPqHWqhugucN/E
SO14gDstpmovpsq2swr0vErrO1V+E4IAdj9But+6qXKcCDVqZVO2GHublfCC
5/psGPZAo56oThPpuxcZgC/9O1pW152N+EJCS/I7UasaydL6K+8WPcJs0Uhx
3vxVu9LoTnzPB1N86g+gid5a9jhxW1RRa68FU8CXSU7OjRP2+sfszx5mzpeh
jIeVdRmn61sZsbqGLHJek9m6+eRtynOPBcXh8Qbc9+wguHQ2xaj+/16Np4PB
f6T35jYqbayZY394qgbGi8/5yDNey+XVRsRehUPGXiQzN+d3D39vhZJ4HdkK
odPu0bpGwXfyY+BE2zjRcsoDav1/v3+T7frXTvMd+QMJtZ+/uQnLkgt2aQdQ
kVi6mSLNOuRcvqM3otf4fxkDbYPrLk7aC8PWhA9A3A/Cm/IG3N8OBAImLkF2
+jSO6eMBs9ak0ei1gkhKOCwJv08n/tR2kg93dkdEDDVITsIk8QC+ZZiqfKtD
iYeOlH4GbPXNl4qaWGco8edzUrZm/gd2tVLAqcVnYJ9fooEu9x+rQmAEBD0K
6BavAAhTq1cW487eEkjFC2EMBCl95R7FyjCQEMQV3ev9/rAmsbRbWr8R0/SD
W0wBl9EsjJP31uI+F2bfcqV2T9XpMIES11GzryabJ7AuL+qPbNYCxSAwTfgI
FL5z1aDzmSQawaogU0R1s+bnYJY4eiMQyCB3cN9Fvxw5Gb/+UIh93pKaDF9y
NMWe/2q3vVdYu92vpxKC+HDmyXcJTjpEPDMIznGyk03NJLz7yNnMzjcrJ0PZ
E/NtO34RPvkCIh3HRPPyyTYnI6HPSOZJeqWMAqtxUivWK/IMyptkxLGFD0AV
r9cJLo2x2pb2/wxJP56siBXIcylN0WuoK5txQYBv6Xll/mNe8gLS4dXpcPVV
h46A54Ykw0KNszxViqkDloZgmmpfky2O1LLIhWNRPmFybC2sg3AiPEj/1NP6
axoqnlJb1sC+MRY9juyT7RGIFhEyac5TyRymUjSKHhZXjVkoTyzb255UWOFs
GJOzIYwI6N2YafNQDuqdGVwLBq4rWZqYgqcuLhN58UQWrbrnJz4y5Vn0j+9i
ukqUeaaMsttgZ6MkTfAJdv6GM5QLp1pb6MluRoWNEoGzghEJZL1MeBZ5XNgM
7bUPPpRgL4y1gW8Nphnv8/RYJinoT6aCeB3zmEYDsyOP+/RRVlMvYEYxgFea
Gk+Cbf8WoU2QsYy/Wcqg17kjP5FNgO+JimHkdUMHZGvFkBTrl/Kc5noUtXxB
XKShVmGMrinfR2eb2gV/ylkm/DuxfOIDe/j+APonXfvcxUaGlr8MA4M3MKS0
g6yf38Saf+5rQzJ3eDyROnkoSFtM5Gj0SSUFDFXK3dIvoMTZjGR6kbAzl1cc
dTbClLojv1PH1QgokPcFv+r3QBfuYpoC1FriJ9idpsD+tV0HS+NGXLqEad1T
36dCAPJSgDOnNZBfraQ0auF+AIfHSUCQKA3fia7U24cZxGOru3kUBI8SV435
GshNKGdmypHkW0cTWo8BiqJcCA9xDHVSjs2SGNllFR59vXsrxS6lKI43nn2Y
ksVcf34dwc6t45QuxJIcv55IF5vNMHPmvhXx6crY39NlYEW1qSajCgWynZEx
UUlAipN/337D2jJ9DpwmxotJr3fPUBWRNkRHpAc3Zi9NisSBhlLIYxrFGp4T
QDJXvUc5DnQXNAniIp5xdR18yWlkA8i8DE88f0pBK1reYFBmG5lMc8426TbT
Q9P1SaA+u9HqJMNCp87eU3NEyQnEPMa1RBv9PKITR6IDmq76KS62TmAM3hFP
9fu3iAgQO9EaZuK6Mg4QApN9+ot20pIEEGdvpZjVvtcfVL9jJ9Tj0CKjp6yO
gj4F3JL6R98lYE/3rW5vqQqZSnu2Dtotmn2R112/l22iM244kbpdcDt2YMHc
EeK3qDNeoRQVP+zgCmmtIMtPjNChbvycJ78gwMJ2JwUg4XHkOdqPwVnD38s7
zDWJJABjzz7z5cP+iXoiIop0+TCSFbC7zxfD532bgAmX5GvabIEsXuQ8w3Uw
w/uzFuZ3z+SLk9ZhCM4Lv5xY6Qg8K2VQd+rcweuuG/45hIAbVCjILg4oqOG/
AITt6YejpDHWqF9G/hhzg8G+Y1gxesKUgsFtNSaWSjYKu1SdRB8i4IIzEtTW
BVV+PBC2bDbQKd/m65Os0nqMHOwxzGAC/XFnWKp6P+I9RaA9tiJNJQlQHGAR
DjWichhBzTMAs8Rj/VtkvdB2LrUQO/p853nXJWFBOpL+u58SZxQtmHKQ5cIK
n6ArVy6Dxc/1xoXOUNlneMT2sOyfnKzcb0KgCqrYHRlxWblklnueYgM0llWq
kccgOL0a06t2lcAUPjOyaeFaRiK6RUodAC7MHXwR85T+OIuGC+6omEIxWbDE
7BD/7v5ImTSOWPCfSY8NQVDTRs/4q8Kokt+tq25MndfNlQOfLChWyJFeviP/
yLf+jiO/fIEvU2p5GH/CQKEqc1ynY1w/KQxsdPpdVdotmSk+8Smdb1cIlbQv
vZLuPWb+zrsTodd0CPpWpZFciWppjWL0I6nznhslS4vY5dI59+m98YmPcC9r
w6JlqPGl3thOjnzyKxScgtKDalDw74DZpP8Aso77HAX0OuTyC33fm4h6wQ4L
j9cu8sLivHuAuyDf3qYdXzfZWfScomgg36jk/NKJ5DmzgohC3w5BVP6D3I7C
Q2AycTagSLi0EHsIAJ3IDiJ6cCOAOTDrCMOPFDu+o3LPyyPzPt0pAXJxHDsr
9SOIYqIYAa3P61oMy/j5aY9wC1Mt9kq7BP5behg/m3uNJpuUcdGjiDVldbdy
XarxWrXOZMgOqYO4dLo6JjJ6B6t4MWL8TLVATd2xeXZJ7j99wR+V7AHDZwXz
xpW4P6d6LXiSHQzm379F9ANn4zGr20rWbwxcKQjH9BaSMYWXo8YJL26f/CfW
Ya4A0cWp7kpZWrkOc7yHiekkN9RltrGPypxhUiYAzWHDxtUD5OQGYsq57HZ3
uGFmrv9wLud++aNqZmYU9nYu3zkb6TqSjYaGK/6lR0LXHl0xwkS3zdGh9JVP
y9I5kXeP6SIDu5BOl7OUsGjrcnP4BFlXBowfQ1JlShcvLMMxkV5yS/gsJo4M
dZWnN0I8v5SoxRacC/8G2PgJD7Zuh0sSD9XC8swB0QdCSJuMl/3woQ+SixgR
656jKUQgBhKessXEnZnnnjPN5de+u0yQqwVC5LkPWECjLbkrf00N/CaLDn7T
7Q84Xutqwqiz6FVUL5tK202If3ogB76twMZCyTfTLVCTWIKr1uBq/rwgvXuo
3Ukrhp1O9xfqQ3hIdl7UVzrq9bkiz5IfE7vI53LgJinENXhaDfsi32cxMpbA
YuW93AjQU+AheGovH/HIX0Nta+DLNVnRtrwgV6+kLAQJGVYs1QEEBhssyzkD
kLnXToasRtezTyjrJq9/SsHaM+Du2gbj8lONv6hkimWEMfjj3wBldo2/owvh
TDXJ0gSnql3GyW4DeJr3QLFu7IrkWtj+jKJEOhQ623DxqOqL7gee8bFJ75bX
FSWmK9opKPeRxYTm5abognRfGG6kXtVCtJpGzqrWMAZiwanDgve1XTeMPEFm
B7rciGq7QJLRvakQtxCyWltlnvTbNq4ZBIWjHieoPXaIG+hkRE94daFALQFH
s2ki5Ar55Da/d/5OCfEiHFkm659p8NJkK0khT+GQ8UdmfgQV29OWBPaBYqVq
yfr69AWdtU8FlME3ikyqYOxJDH/7XAyr61+jpxfMYOoQSUMqXqGjzvmM/f6S
KzU7xcBkSIg59lCHdn6tbgj/1jv4A4vAQMKKvRqO4x3MFjNbcUjFwAmJBNbp
ehasYA5YHekdzG6I/6W8FhN1r4zT5GIyI0N4lOnRpCGpgx+G91bpr+pCzSvy
rSeXNlrpdOEH9Ousy8U6RUntwjyP4vmTg+Tem/7VsqdkkMvI+ye8DhtwmGnx
BdvD91OVGfKND2GCG60RzkIFhE1vdXGOecLTKqdrCR2IpnvYmN9bwqjNVqAI
3UDo3oKCmSx/NQw9YPos8vyA4jJPqYf2TrFovz1xtlCiZLgQe1QEV9DNXSsz
5R7sOEwg9xXKRwg1DfVi3D94J8NPDE0/uXNNy4R3uzmU+ERCA8lUMZB8mIS5
kVOZ7CWLQcZWE72oLI0am5U8SAU/y/q4cCsZM9HSsmkzp1AJfSFM1mBoRCuK
H/idMbAX37BblLMrJlBoDHx8m75MDg7SgO07Vf3kCNVyTeaBV19K9rcukbmF
Uf2k2iZH+NJ05Ql6CeM2cn8AQSBkG4eLlOwHY0KFlf/STGYEdtaynMqrvFav
/QV63WbWr1u7Da63b2mHH6TIRIzImmU6vCVdM8gAkVfl85Kzz1e9OumEYgrl
S74tYNf+UDlomtNgMCCUQqXTIbPJLTkL9R1pbfXnPxTZMlvHSsmg3IE00ihl
2ah0A57q5s923oWVxU7QfB2Eq2cLiGFHeXd99cOBNxHzgwFTpN8Wsy+phdUr
SUm1aGYZXugMCo8KylwgXhzFO+N866b8FyhZlnUhZyqqtZ0PXrWB3k9yTVMt
48Dj4VqhpHlDCPmMs4CUOvfZFu2xXOx8jlip5EVvykRIn4M+yZAA5DfKg5e3
bitN0yyGaz+MC0q3Q1FguLkFmsuc3gS++KSEt9ZuK9L+Kn1xx1Rn6+s6TuiI
ACsiVc+XPPS+x7bmjxYEsksENECNoF4zAqNZQs34CmxYtikTrEVfvepCg48U
1PBk6x2DjQ+BLY5SNofNC3K8RDNu/Zc1hmA7nYMFNH87wIgMAK8W0xR+kLR0
aLQlhvpsbaE6pzakS+KzZ/jWJT7pIX3RQ9QOZtwPmLH1aqCybWotFPWyLtOJ
qa9x1i9TKeveX5JpLaODch5moOnM5u59fA7dC0FD0wuOq0wY0j28uK9lu3QH
p2dvdWMJJc8rjD4RCuV87cAbHcWsSC2WA94w0GkMUKFXGgPNREmMBmEzNjIi
gAFK0NSjVpC+/k1l++qOjLlK3DoH0qWTUw5HlVOe+CZko2iXGY1BDOLjH9A8
0FkjKSQbz2P9EcEws/zmlfnASyV36x4b8AkzjR+nM35VygZs68YiJlGh25bz
7iUO2eE1mImsXSjbakE1NcaKTb2VJLeuoYOHlqy6BEY0HOlSM2XY1zj2+BZG
5bmpviBbKtY6AIDIVprRpuvfA63nC7faCBcu/loc405bl4+RdPCJSNdWW4Cs
4jDIEycICMO9zKCI5VV0mNB/UYRnUC0s8qMiE9OmQ7kfv7RhmPCi7whWcKKe
T1tK/BfcqFHG+DP5oanPBvrpx4hn08CffZBTmJDLFoqlOlVhZ9KMGde/KsR2
NZKVMNtJ6cJCtdkqS+8cMHr11gaxEboSLZWfD5OmBrg2iux13491/JkEfapQ
CTSPO8M/lw5TTc4uLETOhoMngCZSycYvtp9Bi/2TwsldU51SA9KLju0/emf1
kj0S1T69kX9JgVElgING+a0sjfbn+D/S021yPWrIubiL+DV7hqlhX60fOxH5
14CrRMf364twdwnR31NbELS7B4xQQclfnlTxVEGEXNxqezIbIQNeIX10pSBP
KXtKh6LkRxFty5/lbTkaW98XgwxBiiC7Bi4gwOGfWWgsj7k9XSSe6Ndj2/zA
tVI3OOH69wcxVSF6k7bmkr4/dG8wG3Y7lY11WUL0LVo4rbyaV7QGs2CnS8BN
OhRqs0aGTzZqRSDvNyJVRzJ0F9lsz1JQMsLXm1eDXAhkof5OJ6C/pkaNKEA1
KTz3rqyZ/ord5MDzFDqpWnRNVZEvo7XZ+Y0qTEI6UKU3tDJ+5ByiaoEstuMi
vVpVXdlOoMVVtz9x8UOnJrelNHBoVhFI/b7KWaojM44KoG/15/JOGUDXPefv
Hawljo3GkgdswJuVSBWbrQEEUIBbu4uZi7GHLKnwyj7z16eGOao82SotRGwE
LNDE6ACYvbyVjrWBURBV6LD3OydDYf6cXykcLeycfPp+QWbwGNd/KCnY6LLG
5HSTUKxBx4i8/tFBLe3nYacVH479hWTztwdatKrwfsnnkzIiM5uyufYCLErQ
MMKVVKchvPvLcGFp4oXelr7d3CszDxcEcyMk30scIq7nb5Ok8ISc1rK/T2gg
F9ZS9z8C96OZL8HuwUB2E8XwuzB+dKznkwkjvlocxf/RURgONa9hGDz8NTun
tPzRWy0U18ByHvNLqEfM45TvTpI0Vs+fvwPO0Hn+RyOh7I2BERNhXal2W0V8
MGjyRAvbk0AOlKOxJZlld8cspNVfniFPHqqfD+7xoYyUlNcpqVtoT8zavmkr
v81AmhHRHS4JkwkYkBB7qx5aFQk/qRIQYg9KAVikMpAdF8JortHbQir8BqI4
9UtW38f0/Wy+5FUTDJcn0KoJjTodOGQJvJqD70g/aBlUQGEJWA6lG7kKbqzv
FKzvQPgdCZDzbKmDPRQ+MeF9tIZuA1fPK8ug1dDYmIGiaHdZHCpd4ugFJo4a
xja6618XP93uy6rq7SYD+xd02+Ltt4mjyEmFPummAxc6I9XFn6LDWI6HhkZW
di5M7OAUc1rptB/WJYhbAekbQKdQqkQcS1xUk7pTJg41y/iLknRQ6E97izbr
r1JFeQEza2TmSU272dA3MYC92wOAzxM2bd3Ho0B5yQsc6hy1R+G+KPbDgKZo
WSV3wwXQsKu0wkHkCcBMwi71febjTFso6cPuU9afRvopGsGUBuKZVJQoiGTg
onbP4UgtVOhd6NRl7r8LKZe/IWRIVUpZmRTGcyxSZNKbnadxOgNW+KWk6y2w
dVYUNyV1cnYcxImpmgd4Gd6N5Vn8VC1CMYKCYpPn9gsnyj91fGP2ClTX4scU
g2fhe/D+LTRno/0RYN1Li1oAMUtTwjiwwKZ0u3W4CoRi9S0wSCfVXe360Lu4
/9IQYGlZC2LrkU//q4S53/yMw/xjWCP15+EYszrg8ZQjt0yl0Eoi53TMdxjM
/u/9doVUmU/m453l0L3HGAEDRHUf50tXxUscwWFM18ZsCOUOm5BQ57zjAFXT
R6cN5cHj1R6tF1IWKb9dyXA0fYg0c4nZs6RFHyNTf1fOl1IFaY+95tt4cZ4z
VySXPupMPCdp8+uIj0uY2DstzRibPnuCHtDcYRnTktYtXdJv3o/vl8Snin5Z
cWRZvSGHw8LxkZphHu675ziLR80aAc5vpvCckkj9EGJr91ksvE/XoJfjlsfK
DoRiG4VfPITwmt/grulR6BA8S+2B5fi8+lQYrkL9glr7lTjurxP5xHU3UOVJ
Y28o7kck6idxl2QJLHQAalSWysULFegW8btleIEcyLaCIjoYElfl+IfDwg5c
wpCu9sHZzYMPAnHIwj6XogUzGKkcNZ6N5Ecc5REAVvVjKlUKa7+DIMJW3hFF
tdsM4V7wCr8EakCPWgjbhPPO0zFFPmfmbABwvpOy6T2z0KNDNIl/BvVIFPKt
GQwR/yYL9pw7a8+u1Hp+p5PpphnRH0m5UhRqiGkEpAGU+L8MEuDI5c/pi6X+
wGOvLOA0pEUq/Rb/Gz5p2bDfSseMijl/Z3BqIAutDIM1rZbcJ080na6cLchs
aJeW6T1D+wBsSjMj1uzwvGVHlkUt/Q6xX9ovmmv/1C7oFW2DnLezVSm3KEud
fNmmT5NCYviZWf12tEoltvNu6aVinxPkhAOHR69fQFoMMQ5nZSkUrWy/nWSj
C6xTI75Ltl2TEq7xy6uwNntBeKIAnJxXLJnH6aXTWpQ4Ro3e87fm2PWBNXZT
CmOLjWTdA+sSFbM/X8cah8+HFkjwodaeYjpKm5Pg7z5L5ldfV/nNKuTZv3fx
9I6iyTVQoS7C/wcRyquE2E59GO+j6mf5Hv1TkxFLlsqZyqBYU+cc6wAQMQrI
qyyMqsQV2/isYeS5PvHRI1yRFtdfKvziS9dyDrKlys55TH4xKl7O4nP4dhqd
InfG0ENi9BAG2l7CG6fwv1H989WyIwl7j3fDbU75Lj0vlYp5YOQo5/M9mmOu
C2LprR3xVafuC5Snmv3Z5tFOhY7J3ZZBlIbNpuqygEtOKWVDFb8q9CAQ3jp0
2FBH9Y5su8WmIG0XumPwaEyVCs3g4eQNy4/WftrtQnGAlvUABL/XzhlZ5ogb
7J1hXUO6afQdeudTONPMXBvKe86bAmY87li+lPl9k/DayU1Cg/Dfoxg1a/m6
3+/bPh74yuL1MTvU4iqcMo4tIKSsnUfUcKlhZw8V1PfmpiZpTmGT6zjQsvBA
jS4ISPTnOJnzl4Q26ePIJOCawbR4SUKT5yucmu+2oXFtL4mIuaztJCVEn4EG
IQEg/vRdgxNgJreOR37LSbiDgQdlFQ37CfdSptl7eodkEMrj8Xp3DjQ9skJL
4Q9uMha05PUjfCQYFz+MK2+C/IgfdVJS1gvetVIXChfHfc6oiSEHm6PcDqTO
wYhWbYblBhAuA//ulnlHJtoeV73e1gYGcVJJOq8PzOq22F2V5Lf19pV2vFiX
5DcvjsZC0uG3GK/q4/MzrKFqMcu9vlLTPz3uNv7k3SIoYJT3N5LdgVfhlkB4
9kYeopv4sNqnvRcJ8IwY8Vb0YFE/Q7TnXHyUvsumGuuM4DYUhJnoR7gRmwnt
NnA59EwJk5zDaPeZ3cJCGEM+sKXC3kcHGEDmNNs6kb0nvd7NOW+c8uO8SFHm
tS0r/lHVhZYp3mXcfPb6h+c/FEdBHSsV/ugzBYES1+mT4aToCc1N9iMtDRif
BTGEWvNgQRPQYJj/v0BpFPgSe/xRFu39wPE8N/e6Ct/aFtmsVJ1QhCKTfFpS
akkDuC4/r3nW1e3oCka2nzE2lDnhkYaSEqSAR4xkzE0ppxDe16gGU7zBaKGq
Ij9U9KV+bWFxcpNGbPPis7uS4foD1XicyPWk+0nzXA7WjFpDknNSrWxUv69p
wPWcCaXcRQfqObYW1s9a1Zhz4cUpaENPSidRah/9CSPeepFktotzZxCWDJ+e
7zZKJrgSz0f4ULRSVW2lgVvcBbdqhWxQfAnH8ZAjra6ZOrGMvcuwJTVS+mGu
vkVI0OGwxo1oxowe3M7NJhrlaWoFvITlLczVjCU08qiHdxm87SqOAaWyzNEi
6XA5gU59be6d1c2liEq+gQuK7q5Y1+Tesw27B9MupHAmybXMTXkaTmrH6oei
TVxuAiDTFa0CFqeg4Brz93iooVx+vSxNaN2ZkilNduE3Q8pOtQ2GsZzrARIu
ayY1s6T7itJ1z4Dl6k1MNEEsWFxQd9Hm2JwmSxQbB9N6to2g/wZ2TRBk/AQR
M2CyID6+tAJm66kvEwku+xt6jmF9o1IXN2gd04/FKVSv7QKbB6e/KniuMONG
KpqDovficueSYXTSa13WtfcLZhKujhgGNagEmjhnccm4BIBART8Vygp23D3h
NosOAPZGr/+Z/XUd0BuKLRlTTaJT/KXavE9SHdwf5V8WENHPVRjeX86HSAFr
vGHRB8W5uyaLOVXIWYMwygR8P8dHxni6ggliYD3VskVqFFiiaBDh4AjJRneC
U3vbrAXfEaoYdjM6ZYwDaqv09kcXClfYoVdaibToi5CcJm0geIL9jBfqK8cp
Vz2n/lxRqmUBUdVmUeqZiAoLt9Nn5zdTiIluz05DpGwMAbUyCY23Op4C0ZIH
P1LfAKPkYACNWHthSb6LHFdCcQ7TxYzp+XYp6WOVj0kuUe3e1mQ8+FH+2r7W
ljNyuZ5A76v0Oo7wjSm89PBeQ/aC0M5FD6ENG1ODAtimJmWc0v/uuHiUnpJu
itaNY8lhbP0YyvudIpNT8XcJZ8OVHwkQXH2Aeqfb5tY16PvzRuSocfpuheEg
vHck7h+agsOIpqbG6UhKtz/oNid8r30dNyt10c9nzz+Cw96jB5XrHCq97KvQ
lB4ru90mYqUVcowAgFqAu5+gb6oijJYmZLn383dHf9sm7jLr4gdj+w0wc4kJ
6SuFJYPjp3TXFrrxT2/peyLG7UY1opHQ+JfqsatLRbY0GJ5Lxy9PZlMH7ZFx
RnhfPhyZbd4RRwhil9ySluYyYEpgE0AcCc3oSjsJdqk0TB0Ia+gLBT+2LNvL
eKaOOek0GDemSLI2uURTGf1t0xYLzAN3EVqBKdLZwTZN8AD6oR6rHkOhToHZ
kEQ/5vTb862LislE/tFjOOss/p/EBwU7JjZftNSpxy4N7EpxERh8YgFqZ/u5
r2PXaPwUBbKKcAyt2fzj0l//35roY10EY8p2hFIj8yLU8W6/UB8/NpJsW9KE
wfmdrTwV2mei5LTfMZhLiYD7o1dlMxPntGxWMnxZnkm3rT94vjS5tXX8jTz9
UG5+LkwsKB/xPyqneAPkuEyleDnn0wlcl/oDY3zIpnDpYUOHsOKhJ5Hlb/OO
PTzCWHnzKFKDlhVNEadDLDvKqd7xs+O1XXDsRKZzTMvjM/AixpXNTmlZpqk5
4puATBcACsCHWf1H/GoFp1N8ZMBL0uiZsO/xcelf57ebMTyLmyLvPtjDJLSY
eCCY6y1+bcayUXjGh8v0GHVnhWnOcw+zVd/kRAOV6eJMh/ASy5INLROBVO3m
jNwwFuCAtaM23Jn892FsmXgeXawZar/HzbKKkY5TRyAYUvwXGnj2T/NVZ09d
HwwHRe4ZOBbOkbJ/2AP6ZK+YYkzFmbGDW0laO5AEcE6do09rWuXxq+iOuVgE
KIexCI4hzS5D/CvsjyUN8IUrtx1zr8MF2zMw/N4O/Nl4fBPjnL9tQYaHtpRP
voE+8UDmboFDLswOdnqHtDyUIQKj/5UM2fumd+fu06baywfFIspHrtv4jhFP
3UmEKX74FwdfKPp14aBJizWyW7Slj0lrseITyHEyyjfcrEtctw7TYVIszj8K
uQbwR2IutDvGDnVEL3RvTVjbscXE6fPZ+8ilv/+MjcklR4RUQ8ogl6sp7nzx
B7AGtdWHZPWs5iDEb7cnUGRdpgWPydXu6o8LcIRZyadQFPkGLWHlyNqDQuu8
zTIgNQQc7BcqB2a8mrsVoUxeKo6jfExaW8NX+ANl6SUR/JNyVeAbAOVo+ezs
9XXcxM4+17vJvLZmsAv/CyuPn7IOoAHBvnpW4OQ2+psDjdp5PdTixHIFm3ZZ
u4IlIg+Lkl9a7L9eSiRqounIPHlIGVISspHJZ5At+BwoQvtYH2hK/+qWzpSS
0kxAS3VoK1EVQBO032jaK7Fahbztead11sVSpsIzZd8M5CqlmnpaBHyp1mID
8UJ/iJT8vNM5Q71jv74lMuxEpvZFWkCs87vkEyM7xstS4p7VnOZnnEOrMLNP
M2OPnaqRZMsR0GTMUe3/nUumNlmsvj3hUuvKk8nj8CYlZmK5/HjNYR0bUJR4
N1K5WGqQ/1HEkXXNxtxh8w31LOzvSe7g33ovz2OrlvCqxMi04xOuOBV+8JQd
mWoc0ZC4qI+o8IhMEp7df4Q38XqAg4KyFaSh0jhQaMAJVUIlq3Rw8+Ie2Zcr
l48N8kCXi0noXN0KtVNeQjJymcJ29AXmiFftdipnN3xlfdK8PmwOpWhUtagm
Ev4Q7FCvgc64/1BipwgzhSYsHGyD6ErLEY0XPbsgr6i2VQcng9zThNHdh0QT
KB1jLKvhwyuun92lQrWtDS+M3/87jBlj/I60CQ+FXAScXRpY7iSDZyaoLThq
enml8WTrZG2dY/YSL22X5Wja/3NisFm3jUdDBOPQXO9gLZjRTKZNA69xLFR2
FAkcaqL0ZU0SLGA6T+IdSrVEKxqRll7ikxIF/B85sMg9Ejxo54Kp7jEBwDhf
fW8/ZcX3vbkRCMnklXiS2C98GiiOuDoVGUGcJdQ/IdeFcj2d1VmjAlonIObL
HD6vExJjp2iCDBG+CYYphO45jqL2D+p1DUauMbzvmA9TpG6bkz6T3Bva+hBK
2RxrAhi5nbQjoU42gm6SdJ7B8JyWXCOcE8EkFHxXtfVGO2+9WCfO5LMIrPeQ
FIzFqQLlpvYWteskR5XhO9YVd/m3idPDPlP4wO2+RWAZmd+r95uRa3it9G8G
zDDR6FvXKNjYXOyXXVaiQS55/UjaO8SdpRJdy2eKbFf5pVXzleTZ11o8fwOe
36wWkDmRP8ds8yLPtR56RdAHB5gnvtYsKEfE6nNv4Cscc1DPyPEe0DqXrBP7
L8oa77fkIH+ySkyMaalTczOzhY/xwWpzh8nb+mePMiMD9h4iLDq5Fr19Mp/V
tsSvGIHCGwoPUCXXWu8jb7xtcVk8ayNZEkD12zvR+TuKXkY6RWSKXE4GP6S9
CvhKtrNFKgoJ2H6nh2JV1JjwDzBaaiqK7Id3TPWX+ZyLWlmjaf4L2BlkQtFu
c7lWvJTS4fSYMmLyEiict3jTe7AtjMuRwYLlxBmICUgLV7+qTvAUNhzCtR3Z
d8uLeUZ5AgnQbPEJ7Aj5u1zt2PIlUbpq1PQyEsNQsfZpGodACmA0w0k6P7Yu
LFD0CMtdgbkMuchkFhA6vdGg6lsWirpY6L7PpGbVbMX68rZJhaThZRafKdhm
XRpe9bgqczUsXHZNP66bB80mw996a0u3FstLg1pJklAaqE7I8qa0qGF5dvyX
E4C4hJInzpwLMFtagk/4v/ZXoqxbWmJwpq1xQIj4ym83Z73+D3CymLaAQV2B
yixiNLwggj7giBNp2LQ93CmehTSYrFN2ToCt9ctd1x4ekvlYQzA+YbSQKp/v
oYlBX6ta3KwWICAiSp7Ta1Gem0E8dLL+f7/GFFAz7Dg8AmRYdHTUJPloupdW
Vc6hyo4nvd9qc9k5txvrTLnyMiYPJK+UILAh/cp7QScf0trFCo8rjCNU+ljL
yz42mCEYY6OmM+9/QKVcw152+qbosgHanH9i/f2/7m96a/Cz9g2LaHzYccja
e7JgRxNGYcdOFfEcjQ98ybav1UIhmXFmSX97p4ork8aeRiAieR4zgJfEBo+n
awZXGJddKuWqWoySJnldd9c06KickewyDEfae+0zSQpWdSN84IZwVmqaxtOY
kbKRT4Jmyy43acO2B7GJDa1jBiuiUh3UUaqAYfA3TQgZ3OSLN8ZIJPPE2JGo
C/xazt1ou2WT9gdUfqfJOT7N3tphpcjiwIN+ISf87mGcOUk4OUGSCm2L+0Bu
fJKjceB9ff/Bnlx2Epqrd74YXso+jouZ365lagpgkKjHa1uTP8Tbw08scKWB
pkCz6I/EJ+RA5u+qsL9AMQVYfSEUzXaUXun3n0aaYaiZZZrgDhkcUY+TZoRu
cJqoqa7C56fvjWG52je1paZ8QonGjNWp3kP2G4wP7kOthgKIANmsWAYoJcy5
vEMEqSaFaH9QwksdeP4BAt6vveFTkYTVldEya9yK+/jHCk1JSHkxyQpxWzhh
DpK1P5TYY+RQ1nrmma7HleN182AVioO76pJJZGmU7QqtOOAmcBt7g/vz09yF
SxjPZpU9eFc1ua0+yhOvz0Kwghn8GRJkr2icrC9GO8A0dPO1G6KUzhCUzJoz
hsOUghq+f+QpiaGgZOn/tvBI8oW9/hi67Rbh6rGLdZx26KrBf1yVUvCHHSme
2drW02tSS1tBSsUv2By1z2rCgpxnIOuGEEDHYeP55RxwrixLyli9nVlfMfHn
T6bCHESA5+EI/RfoAczI/xY8SszI7pJiKgwfK0MY9CZP1LIB8SiTLBgKYBn3
gq9m3Y5BYpGtWXY334iW0gXOjo3fDt/CZpcH4cwGtrA6gQ9QPTAPMgRvehD5
FOPLCy8djvhV0pSdGjqOUHY3xCkO9ho4LIunw61g/tHPh2RWKV7owxdysrn+
SbqoJP400Bw1N0PEKfRGT/Ldx6ylUkbkLcNh8WpyAKKuKLAJeSs5+sx7CPdo
b31Gcdb65mwth4FjmvMOFZooSGY3EzzFsX763kt/zJqawbYcFsj7uFczahvv
1DlipN4qPdW1rKq7nHTl2bZ5gfXowkUvLEjnLTPHq3k38bwAgALqS8B5Zfge
KbDQmYwfhUWT/pugKo//VCbAZ2EkSSqyaJKw70sZ0eaHgpkbKlG1GvuIcpwY
TN87/Z7FXmlz4v3Cf7hmbHpgRRLjl47cPjkQlzQp4B4ljUZI6GfCotxrJVPi
4l+bZp9U88n6nco5BJ5XctXCYT06gLpk25X+0nAdbdKkNcHj39z4bjXFWRQ4
paZ6kNVHAR1aXoR0ESoYqAXOy1nOZ60g7tkP7TjmJNl03H9H3cWXVpCIG3Gz
fWH2v7F6B5Nthc81EYqxpkpCtolXh2jLSUzim49tURzL3fVLiAYlxT7fU/Tp
+5l8A9JAKa/MvPcwoOuqH0vwj+cJ0rvl5/R7yY7DY75fIFTJeIEqHAALQl8w
DkUDfukoSWwgN5u7Hx664QhO9OiPiu/vyYROkNGbj7qphuNZe9PaiqLnM/yz
N5hkeS+gQkeGNIS/LYkezKEWhTi0IixG67Ke84e+3JHDSv+ithQuRrNKr4uA
DT0HwbwxudKYZZpniW+LKEE5W7bt8GAa31U4u4JbWhzfHEwm7qaErz7Uoflt
FwEQ6QZxfrYKWKMYXaFyPx5Yrn1Ru92/qpkXLyWHyawbcqdjr21viYIEyIvg
7Qh5W9aP4Nbbd8Qkgj6ccqPKmubWcUP358iDIgr0rOVfCMn0OMq3ajoRB7od
Ho5CDSLztSswgU9HEs2rZYJNgW2cz2eyJvsjJCZSYlY6aup01Hu5P3UIHo0v
PSUX/iX8dqXpooLPSc9MB1PyqJe/piZUGvxlKQyCgBlcOFot9ycWhwpY3Oj1
mwHUt+rh5ltA+fK9heGDmDgVQF00hr/szHJIIJkwbELtyPutcV0rzhZoJAsi
tPuqr8yQrqbQppqHozqFBGgwjK24xFGJFRYJhZXhZNPZHiwHXDlqi/sYbeKv
yfNTgs0/BvUJ7DQX0SNS7Cu7HA5pxi8cxGtP3O1KCfou01pgod66pZQCMz4T
ErhdVtna+dYtvT794xay40t9sWaE897X4m2VQ6gfpKu0goiQoMKS5OxZngnW
6wmP8hpQTxP8Sw3cUGD8vts/PEW0oBC1xYOf5Y9nQClEyOjC+ptLr2B9vQjZ
yWyXtG/TdaCuaxzwqSc3ZjfTtUXtok9UF0wuCkGbVUW5HemNzy3FXi1IRdMq
12ZIvApI+ir8YGJm+KZPhT1yLh4jl3syVOcgCcH3IA3eiL7T0ZBulLspa8q6
o/TrJqA4amZr56dEcab9Z35o0uYG8XzcSVmyND7uic3dBlEzNEdsVFP83oLi
gmkkd6IPsru6vFtPD+rGzi+6YYRapqTMyo95cx2pYvegMe3MYASPDdBeIA/6
jmedYsOFsjvPMMKF5T7MbPDwwyjbYR19/m0knWxhRpVE6ytY/ukfzNWreP+U
FophWELca3hl/2dkZi4DSPM+sBJjUeBKhzz2zSexJuS6ChQ/F/PO6iRX2RNK
mJbfIZUj7Si8X+q8T3FdK6ASz+/qBLsoydKtnOw79C2+2YKWkv4YCA9VLgUR
ULsJA+lPxV0VovqWuPHIvCREY/8JLkb38rg/rWzJPz/FQhOFFYpiBdVXL/lY
adxpQ3chGpeNkRnwRjiJROFlu0pcSzq2HzithxLOx8eztzgZ2kJQLvic26z/
dJzdywmxwUbTj7tAogc5Tfoahn81VS1y+ggrVzqnvKSbPSMqwr+eRqg0Sowz
UnZWadi+Iye9un7D1Q2XG7wW0GDSVsvvSesiKTs4pK2aHXg7fPEdCXTMdSJw
U+jejVI+P7OWm1fr3gFYm/RmhjN5gfVwV3FUoKslatV2bRfc5Xx6dsPLAfHo
wxjAZoaUhgWxP/9KSTJPsVLq4+kgamdxw8+nJwAly5mALYl3Tx96jSOct8kb
BZ2v6oWjLM53gnKJzBZQcfwyf3Knfs6tg7XJuyKBhEZnvrNZ9qG3ciOdQCSt
iNjkSXIYs/vnw7X86w3efsyE7pp52o+TFMDsU4Cd5vbEq2KYDaLfEx4a/ASr
A+FGIrPF87L2ocWp8dy7bCylipfLLGUcCHXPAM14+NUuIlVUDusUezbzM2IP
n66f/LUmYjFDHzoKdX0r3heYnwHTcKj4c3gszQkNNlivKGp2/J+z5d9Ww/Z5
Ta4r4RtHmT6nFLYRMeAJSbm96IAN3RSjGmye70H+YecuRAJq3AFzbbm94L59
iUJZkcd0WKOpFqbeCfftWi6Ur/1Yv7zc/GIqvLvDQf8OkJ4vvbA4OiP5jgj1
z9za3lVV7PLGn6eAvuZ0caq4EC2FVAzrxljpK40ly4Ydj1xvPVKpUJ3TJxQS
L+Int/pZPT4TmxmDOo8ZKRYT64aaC5CYtrCseXBdvY6zb7+CrJdtJWvvURys
F5HxW65tR4UhqfPRIPNhZJENPMzDWWlvB25rt3gKbXD7urXNcRlgZ+eLaXbA
lvMPvMVKr2Wsa4Md8rL+Xy7kJ7Nz/mfJDa2+doM4E2+NAIxLNLZip+A2NW93
o7RgFsQfjsHO1GCka3axaclbzZJrMOWUKeUn2EtIW4Gnoc4mmNNHiIGJWk58
uqyskppPHbZSc+VqJSctNb+jPfoD0RJtTinGaZn20+925w2O8Xb/Fg37MEPm
czJinsgv/bBWXea/56bfn6xwZAoOf3zzZ8Mx5ge9deQONzax3V/ZjbFTGy/3
iaFj/dC0Blv0zHcxjMN6qqleql/zSKee3inkzWe39AtoVgnOfptgsfMgnMc3
aO43qVKnUyyzK9rvoH/VWL03wCh15BJNGDKwDJpAveZpfWrjBKTsqGwIw0o+
cibwf7aOdSMxYY9q27/JY3RpY5N3N9ezqVN+MtUuKRfy03LxuPvy+SzCfKAo
oEDa2NsUq9NDsCabVXLSXpSKcuLlIqlWVKrZ+BSXVejIPC644KyH0XVJqISS
esQvJIuyuLkjriDlnimcZMLE2CQF+7JiZvisJusSEtNNXZVZueUPlkR79VIG
9Mm0yUetpbek95aP8Q915c2rO01Idc9MKkvSqaUc43VhgEiYrEOOH2OGUe4O
dUNsFxOvlBd6ol5fFPwXBwz58YSNV2xI1ERpbgnEeIiGH7rDs3GCfbLjJCoH
Z6NMgkJ3FOVc0v8s9E6SwNrJ9L38ZyBwJWrWiKut97orBG8B7OA4HwyJhzTA
WOceQhwioQ/GDMW/9KpYo9/JFEX9nFjT5F6wBIX0MXBjsH0xRSxlO13rQ5EX
ac1MD4M5Hs6KcI1BKVfQfm2voHvDFVsdo81szlrZA0QilahcAQcOQTz47kFO
bdmAx1nqRK5UvjB45YAkXkn07qolRqrgye4456atJUaK05X5SxqbOP8ps7mh
jSAGWB1BoizZQR9o2pTnuhjxknt5c1Fgg22BJnMhdKc5c/i/EQG1wWQmhDem
1PbvsCyHHF0tiXJq18ZOac/IUZtMXLcKHV1OlWDP8WF4aw4Qw66juVCp0UbN
VcUUleCu3IPeyQ5Y0MDrMPSk1+4oqnls9ZCDdHhWbC+SKk7wrVbNofLpxCHQ
i0W95xnQDo+M8QWcAPadzDWnOmW521BkkjyXjU7c+CIVF6nAxhuRUeydlXd5
go0kXifOIOVvUPMjiyfmoUCgAUc+Ji2ZjLneG+b5Je6cCLoYmE5ubEF2nAsw
BktutuW1tCihnxrTA/ApfUU0Dbdn5RdBiSbcCp3H36FKIHCqXCtfWnepUaza
9HBasaSYENelLzRtzogG6IuhYZaD7qH4BR8ULYdXdBN70gqGvz6X05qX9Qao
jHzgjhvreLAkaaYQzCIZ8a/phnD6sQO+hTFaASst2NR8EUy4553JAdyTTo5x
TDmLXil6+5RyIyKk0+Njgim0c4aVa04LwJsvBD7pyCQinVVBUoGI4LzWUzlW
C5vBOhJaNLjCappbWDkd8NBTFiX9hUQKxwARhsfr7hYmoO3Ez0oc3OhDswBi
BJ2LUeyALsGMbuEwggnUTmhYFlqvj579/49liBVJDqhF6aS3qXGwGnUn7geb
XO0vO7ErpeSGCSuabySD5REC/EU/kJiJhyKOZl3KhLYuJ1hvv/346oTl62e3
gwNyxrz0u7n668WGUiXVSoLib4KPAtKCRxFcPtdHrzgEvumJzLYH989/+Ss9
qOH46xcl3Us20Th2NAK4laWlCu2a9R1ZbeSkyMDVxNDSSLONuRahc+Vfkin6
HCzR03+iNncN0nycV6ej2eFjrmBIEH0UNPxygXMFgSnW+l6CNFvKKa4MVEw0
oIHzMApQSD3qDDkkYrDniLyArStRZjkUoetL7juxH48g0QXvtJIFsFt5mv/3
43N+A4i2aNZOqitSTCBxuW76es8oZqafhVvauibRqLnkkrGBntDUamSaa+Ui
CSUNH10b7bVuwKgeqZ5i5gdKd0bBauuKQB5MN0eThUDln14TJlOUCALza7YV
nzNYWnVT6Rpyr45J+Ke28rhJ3klSJmJjWq/O6KjuJkN/WVUMrLwlJVfAB2tF
Xa9Thn9aVsvXa5c6mytPcajFyBdxBNPoIDkkSyuaeJN4+FjBhtEOZm85luet
Uu/aYhKBsNQFgqPRbPFwh/0IxDqe2VQXcrAdsoFtY8J7L+NN+R1Jav7Tpqan
lLXfauq0/rttdroyXx7zfIW0BX6HkFqp8dYqhAfxadioDpmw/fWWgzYNhu8E
0PzCCOGgiXar+qXFEBMoiNRpTnGUdMpb5A8rd5hAqzBwu0aCzvslmyqHWHov
h5sTJdg2Ha7gaYk935DByu0xtSEXYUtNBANABi93IlH49PnadymrmCqwOf41
s8uUu7pi1e+5uVQcfTYzeA8DrHIZ9g3l0JAMJhwflm7sn/z7to0mKT+YB83i
QhIwy0OFR/ENHlEplgEsKeD477HjkD2lQqjukWVdS+nyd9OM68VFjRejjyWE
FdH94kf26dQKuFURmNXliBPvTg2MJZzz/OUHUDT/KeKc5jAOhqtEJn2Tt9bl
hAqt02AF0GJfo3BmrXSMolOOMsmregG/o+Y7oVG8ptNGv7iEdn83IBvXdfyG
dK2vkHQ2tNB6LcYr3LPNFvh0w87uWN1eKaOSgpoXHCaukbqMP1N8NvjlTSNz
cVoSMQiKrWPzHP6HAWkvGNwaQmy0gxqGZSMOtreKNWKUBYHv46H8BAVEq8H0
GOpwSZYN4D5jwAKuyPaJaK2kUGBFjXTGz6YDfYRUnOanOLF1wdUwF4o/TFoQ
1ewyHDP/d8aNyU1s5qsaYBfdF8V27SF6HG53roUSW4ixoiUm29wu2B6MlyXE
+rdxxHz6hSX1Voy+o6nMFGBMzoPNkqmVmwy3RT5p/Z0Vk497pFQMEmuB8A6e
2IdM6gxPj6h9c8uEC/2g+PUmMhXA+ItzC/t1ktdYsWcEiysOizKmZT+MxYHy
+lVgbKToZSBzJfXy85WMKFhvRNWk9gZBNPWU4+haO4G8shrAwyQ991XWH1XV
A8BcJwfajN3kQJ92xBa5nCKtL8mPKzDRPxkpzI1p0aAjniwqIr7WiwzGAzlK
Z2mq4XmzR18PGoVE2Q4TcpqRZc8/6kWGGGYEay8MyJ71iqLJuZgUPFMCfN0x
KxF29ZPgJWLfLIpGUIr1Ws/dxASotbuRPqQ1wPUm57kQjbEonIdHa7ueWWH0
9ivPUsvYdwxpg0w8xFswIXUB7VX+XO46JE0uKreVmlb/ltXZN4odqz7zdxiB
1QEa5bAJtuy4ZYCRgnO7E1u4faiUkaH/0DbYi0vSVz8MCw1zFunPrFFlGUm6
m2/CSMN1s48a/5Y3ZzN7LHkJIFQzbDC/3ASxoyvMczDURvTN+NnahaIJDz1r
xBOFYd1xDrbQy4OQfxuDNZ8SfdhknWqA8Vbj6YJRf8JOO8CYsjG5QWq7vT5I
oIzlfDbkjR8hzImGgoYd1b7RKZaAlPH7muQ/WHr9tayLQzFbeN8GAGkkBvRQ
TFrdzXxlXOmLboNZW9Nl1ZoccSxxJI77CZptLt57NmYjxUgspfAxvn1gI4UT
tBuQy8Mm1KRdqYqmt4taNmTVtnVPK4ulBKEI9YqmEvN733BbvoMipSexQiv6
0+Yxffv4szBFE2NTd76Onuw8g5I0Jqz3hUTv1L0FzlSLwNAQsjJiOmzGt3KB
wB6YMgVcUjkpkIqBM94fG8eTtPM1WbvFBKnZ+ID6GgC2sUY4Xf8gZXpDX6KD
UBRzq7IorCFZVF1xAxjr49yAGgBlQLvynKwhdUrQndCaUUwz4MBRxUsxmk9Y
KRU4vfJaPgRoiqir3uqKc48nNqW+6CX8ZGcJdZX2IaAr45iH2a4V7JEFJCI8
qayDqyM6vy39xbsQ5lrcGcFUj7fLS5smnXus36bkJs0qF7JfkwEE9F0uqePk
k5diCdAAc0Dd/JmkdL5pzYGxgLR2yv0HpidW6t0cZ0izP5P8Pye21gzTSpTr
99QoBHJg7qGLH23c9OD5sa0257hk2yoIMHLjV29DqS46MFBqG0hALuDoe3ic
UqauQSiCWdepHgpKtBPQcfu7NzF53DgXqzfZ9UY//1ELHJsmHtSW1C8stlac
2Sin3DaKLZRHFLbk0iCDCVgqIIfKxqieGQ36y6of6KfpiBmmDyUuoGE0SpgP
QDsTzbt3JVSMLT1bByZm4cVOKpnDRpyt20WUepJ8JbobaDxM3/5v+Gcf5GR2
gFxe7B7Vs62SiMIYj8zVrYUM34xoQQyc1shmX3sbjFdmDUvOSSnOWf0chYNj
VCkSEhuhRGL66OElrDPVWFLq/4bKQX3aZg2JDjnKcscauLv6DNh2/ff++262
wXd11WNqqLfgkV7ODS+SlrFs7ILRXCFJG9mOf+RDluIg2QaENDan0auE4DQ6
2tzv5sJqbmvflmPrBs6orNO7DYVLYvcw9etzgfjldIkAWfXDPDNg6/urtBOq
9gLDyVpusMWz4G9S1P06O0PEPZrNnQbMge1EmRe32E9w+Vdc2WzBc+ieVbxg
ZDXkKh4ZaZE6ppQAYCcvkrNDlBR5XcszPMYx3ifn5eqXwf/oTR5MH2U/IZCw
CW2RfRXZuzgLNSljZKJficcm+syidlSoVvIUL2AVyL+OJAlubtqn9a706ZQw
1cBID6VATkq/rWDMg5LSD0/XIYkDqunAKrthKIC2PGQb4e40LNAO9Ob6aXYN
M6YSblSMYtXsBbJMI4VU1Sq0KyhCv6449WgCz0uARcAzbI5RDySaSqJBCORZ
bUe7eu3eiVaqMf5No7iiioPbIZ8eaG18oAjUHP6ge9BmEL+Vtmlb7rA2DwYL
cLoJzLGkTkcBTaBHHfOpAY/YFVk/isuwX5WSAe4dIjg1RbxWDULF0SYcBzou
/VaAAn0jAzLWdSiPVAoHCNzxWMFIdB8wG0La2pFcy1AsMnAbmhX3N/zj3jZ2
ydpZv4OnUDitMKQe0L80I8sCu5oWP2M2cnxi/TQ/xXt8oXZ+a3z+ss4T18bg
NQ0DyYiyBdM+ahUpj08e984wdta5QbbOGNTa7bYC7LJXRSfq330MHB2eoANa
v/0RZmYQMqMOA6UHdQjhra1A8Q2UvHI9Uz8WrRQpwfUBKZqRsHhyK7m7FUWu
7axRiK9zaLnrJV3LHAdBNYmPW+ZBTatJwrL+dfOhkih2lDUmt3LWCJVs+uFH
Hj2LN16bikpotNYOeYelPitPbzzw7ZhmOzAZncHHnkD3txknKSmoGHrwTYzP
8WOROrRrWRKZ2RvsXB1tRuJ//xJZbjDfHEHaXtKzqzWHK3SeHPHYO9OEHrMB
vSTtSgyuwW2NaUdtU94tLhJma9GV4SW+eU3PXkSAYs0y9T7bTixBl+7T6tj0
yMaia25xVJsUeuDk1Pm8EcpgOdEpiGqNG9MekfWcLfKP2QRhlbatVDr21Z1V
i07IFuaGsRupLJzl01E1viinRDa0Pi9w+/2kV+L9174yrbWjJc/5ApxTVsAk
arxYWyuwA+r2VDDClpYvJqUsq7Z25ZoHnjIeSM0dAz8AJmA2YFW87he4p+U5
lfCZOUy2vH1iQokFK/CWe6i+VNvdCI660E0Sybgx0zBs9DVsDCNjubKxIBvZ
w5hks3lJ6vYgEcO43GRV9tATXAHSNaMFx5wrGALKeQ2DPl91otwAsytHpJC8
orzEOJA6mrrT7JTFhYdrW5K8CCTRKfBsSAMYFhzSUywhiLhZYi/2Z6GruvSf
BrouQhWdmBtiApOr5WrABdTv+aDu3HUM0NjfqLo1t5gOMx4ARWM6mOplXCnM
GyT05qFaU9OGPkjOWCiMCu0YJz3qbba0sgb6bjTIx63bLsK6Bgw9jwNEI5QG
0UzDt9bDz2AdLrX/a2lJ39yd5LdCviGL3k4OtbWAMdyxnbI0zlNA+4mt2gZN
hCtxlnxqe0pcyqQtvcXFEQ+5PxCo8m4swLWcpdZIx7zjuPDZ1XDbdhMA1i2g
22tlZ5u8uV6AUrLgouZ5E9y0t2fJZmTHKph5B+5uCzw3sPjaxEyK3pOjQ01a
9JDVPHPg7tauUP4QmlakVERSJuRWChFPgkzHUUdXSoW+b9W8/Qcaq+I/mY+N
gJCfgdI2gAROmPWCq2vc9q0xIoO86oZMsodcsmumhPOx58vp7EmkiRXcucME
teguvMXDCCI96CwYyEz6fLahB+nn5089Ihd5mfAwkssOzZ+bCANg+c4Hm/dW
FQbZ2LVSUMUdGmKSgHdLYNQar101Q/EY3+6OpqK+gqB1Uu+dc1YmVtr2svks
rAm5y5+7Ix+2VzN6To+ZCgSLRxQNakdBmyFf2elPlSV+5FZcYpNJNHMw/G0v
LnwZIFKUpa9Km//0ULnlhQYb7NwXsZABYPOOv9Y2PDJJwofh0hL/Dy0yH1XF
g+3yHYnMH9ss87tNwLEqNYkK8WdJHLQYFW8vnK8nMUy3UitrPHXgOAfiKULq
ykZZTg7uN9hNJWvasR1sTfMsWQUUrsYzq7rLAjXaOTiyETlInkrgt0uJlPDg
lLWHDvaeTKJN1cHDupc1weQ8cu0as7SYalwtcGwMWVu0/8otOirWulxgM49Z
UwAILf/LFUrdOlJBnDrxaw5d6LFgFNpZtkojcMMWKNbLbXsuqdxvQ+OHs5pG
+tmt3ebuxTYnM30rcrfUyrTPAgsZPKO+aZHlcKEkOXX3Z5AiajxiFrb/tLtP
JVH3PrKjFItKKGHHedzsAUjxYPMIMIrMRyOXFR0FDpeyNmG6nuxo80BU4a7g
1o7u/+0qaEk4Kl7rqYddy+UlaqhY2E+JybZQ+UowX1eg1ovzRAT69guB1b2e
NT6YUV3m6fihbLQF2arhcNRcNOt2skZH2iLsSvZB7bOpDav79y4sIKi+4Hgk
8dWgUcrtpFpF2GbyvIKiASlhJcqaFJxLqEBaxyf883bAkmXAr93Grbh96U2q
0IrrWnBLfW2IDj8aKpwuNEl+PBcAtpg2V+TTMSCqdeBOKsPYbKTgjSCkF4cG
xnHuiUpEY+ObXzxnylGtCZojWvaSUn1hoeMVM08zdZhHhzC7Hl6+OFq5I3yG
6cwCYYQmlVlJ4juKqvBjSsuaHuN2kLbEazR01uazXVSfTra+TZqCHOEEHy3L
csnti7DTm2KF0RHP4zkNyzy72sOIG6F0xQysd6ck6FaeIO0WhEmUVU1ihvH0
bLnaVDQeNtBg6pZipdI80ianMMhHszkjg8gK2FhIy4oGZyckzHiugs7nYM4o
EdXDlGqZbdC2JFrd1GqDnEYCbS5qYy+4XGcdgAaAPYjiBMO/MTkpwCv7JH5S
/eJyQJR0r7tQDfVzc4LHEuT2U2ILCdzKBnOfw8FS65IRUV/lNstoNgAu/AJU
ASQksroDS+QVnYbKVGu+GABT9NtGaSrjSGlw07ghY3lfn5924i6NKoSozOra
TxHyIcuwvqZivzYbDKx8nPL6y7Z+MJUPpgpTEctAJvnrSbtYIe/5iDIVbu/q
B2IiaXpDCwaZs6M4yRvZJuCNq/bBRLXvkGEqU3VdgiVhv3BWqMGDPeIvKQWR
N6mOcXTMfbqfNhc9aNvVjBXQf31pR1V2meVGdBa3LemE8THmRuMYaybMqj7S
ErJMV9CKIn7eDVTU4uNjNofSMvG5+Lda5O0utDkUMM/cm7F1KwwO54V/EMQU
Z8LpTtfQMggbERQRa62ZWo0/+ZQzr7M6eIdFUk3IWSnVTmPC/1/7WaxXO+Ng
iurTTVkKAAiCiNMyI0Q48XxXo/AKN5K0tTmNv8CKuMYah9ZS4//YV6WU5Ycz
LkqZDxXAFHROdIErP9Zj//ES/tncv1SZI1WFGMcdhu4uRCjVempn9XGLsJaY
4xC4qeby9wX8hDvVu+RhqJRiNW5JX8RNlo4oRm1LFvupuIfvgh2+JOjzdbDV
SnCgmwXoqiGA9jGd3Nde73DOYNtb0iuWN7ekMz1APgCksUVLXMvrAT6A67Zt
ljiTk/rxAbhjZU/oo51GUoJh4lDaTckFMUZadOzM/L0t2Weh+DN7BmPBq1Qs
8jZFsmfrkTFVG6n9YcXLjXeV1ffbe7SRIkAQbde9pLEjTat+qem17OdWkH6k
VajWml03AalXFeGbDTi3rwqvEmLiCHxw0GwBZhzjcaArwWu7x1tx2seIpKAE
NVPGVJxTaU63GfLUEMIyo3jQliBM7PVL+FbFXyD2/dm2zY45cyvmJ6qbctJA
eP3C+npLPrTQS208ghMXLILq6s5nUVRLW6eHdFn/Or4sf3TTF6OOom2b9nP5
dNNInfHjxDVy87kUqemnrWYujgDPlD8/sP/ANd6/K/XGSV+fUnKwMW56QSzK
FbWPGbsv9MFZbj3vF8ctEf1Ng1ikH95Veloaxd18WwqIgBJCMRGM3bcXmEE0
KXuKDMVAdMKuYeSDdwUBG+nKclsjiQKinfrPq6mBV2//a95JGTzjOnaFwgR3
I11eC8lWjRr74nTV+a1ZijHqNoU5D5BvPAkmkGIncxL9Q/U+Csss77VOZrbN
xvI3AYuC30bYj6QzLHlofJGGiIBvZYDYce4wEawREKFHvi4JVYcS2eqZmHE8
Lmi+E2w4Z3gZPD5ZxiHn0EzXels5BxTaVuxg2kzJnifqp/vJuFDJNmBsNiiB
q5IqaHiZEI19MXIsZPwYyTtUPYQzV2ZEN+3Ze+K6WteRhuordJdCM56LGyMl
0yZk3Qb74J+5Nk7ym+G96YvkoDHh9J4wc8wPJDRAOfPLRtghFtBA3UDFNEEG
TPVXwAHLAjJE5/OjLFl26s1bp6+2UkQf/bMZM29SaxZcoHKRvtu0pxEUMauR
EeptdZDr/HRyqL0sfgtOhAq/Jm7WYASDywUi7jt3gpMjS8xTro+gY/XQTTNK
3rbbbd72vuuunTRyKasY95ERVoH5HMV1g/AafmK04DqAnk1U+lI3hqgUvXCu
6OdWJq4wEYC38oF7ioRbx/C+LBPQQi8ncOmgFO7mtuc/Wy/44R47nV5ThMaP
o/2LJ/xeyZyQ1ziKdXpjrDONAh0pqJiX30L8rDE7W7Hfhlo9nxUhEFZapLKW
NBWK0rZKrrfpSYPf5rWtNaoaIUGoiH4KUhFX3WOOPRGVYGLHFr6K3KAFmJAK
sraYOY/EVa6JGUj7gtLsaDj17REJURVn9W+BL3pdLUuUcg1CwVg6zsxqJ04u
9JjuW/lKaNzoWmFZlHsz2J3w6pwwFPTeVFugak701iMnDn7xkZTF0jgnjs4v
Av6njogz5GBgE3jps6Ahjv7G8tBkeey080sFW8YVajxKoUGtBd73CDhYccNf
M2L3QE1QDdningu7d4KzVt5DiYk0qv0t4KbrSkskIcxbtsgNVcN6SSvTanHW
WnTIiFNnN3xcJeSccEkp9F/MS5VkHoRV0IyH/8Lz3UabKSFCBRSzElJjpUe+
6qLFI/KtTW2K1qn56JdqzkuObkw04fMq4Krsu4UgOwnwPP5RAivXUlPxMizG
1G3Jl8687ckL5xF97XM9q5m06fbn7PlcgWEiaVZ82YGXu3VpOH+mSkjqEeFQ
t8ejThSJFp9DwTyWG804ubbq9FF9hVzLfggJ4qVVDulZH8w3bgrInilG6FUp
603EUhftVFe2+qws8TQTlzqAX2rv2rnUUC3zsosaG1tOTkXlA7I5bzrM9dI0
Hw+X/X9yNkQChngb/1YVZ7ox9pgiIwU7mkteXO/sHteuuNw9UiQuXLWe/CgQ
S4+YUf/rdvCxW4O8wA0QDPBAoCHrohq1mRWCSZe0NKdU4nHLAdmmLteAOpp2
aJApYWKjSqjhhQkDSDx1KGHJGvUF1ifhC9KS5pmJJ4RAso0rkKbMSblELak3
U+6kO+1gW0B2xgI4twpAvbepYayCEfzRMHXxViSFco8QF9mpcfqbhLetlCcY
k+/Y8yyg4vWFgZIwc/vPag09oBEClINeqXdXmTeUZ0RcazoDLvf1BZcL6rK4
1MhMFNWHuvZSsiCu0EnZKEhqx2J/QgczpP1L8g4ouxvpqegb5LofWwMbbela
uj0jZP6LPExTvjScSmG9vmOZaoZTMwS/gppS+16N+UYt5KdFviLzBVlPC4MH
X4go28lAsGIaHThM1X8PefkeXN4UU7MYRBU2FXAdlvd5vlgaxPzSEwuOB39o
bSPHIDuMM6X822BHUT2SAYGSYSbxyECeipgQCQN2sDLDSa6Q0QoledBmx04J
27cmKz6ZrHPMZSKaJWkcEBfDfYN+1Legd4Agr7rfJy/2OOp4mJJzjCkmxTRy
ImNOiF9FZjipH+A4VeFf5I3eKuQ/UH40OBLcFmP9JrEo7VCAajHjbEDD/2Ra
DzsGdIt0H06y0dqVuFZ1T7eWmcKuMrRL+/nOQjRUHryin/PCFfTzWFNqcwwB
/GpJNGaEarlZY2iRiyWHeZ+0zQUdV8shoKLwbr1ZGj9cqgVD+csNaIhfNiZR
8Y9rIX9hiAdjp3a1LC0x7fIo+nkbz8H+gmDbR0CQoILKLUgdnZ386rPG9e5t
96hemBfRTzUA2Dc/jZic1ChToJbAzH00ML+xshvtnfpuIfbAOx+0y2/B7IGS
RdkwTXB4cC7/w82pPz6zDELYnbsPVDdilkhzXKm6iO5ytA2Tat/z0WXqcmg2
SPhDx5uOM9pqpv5p8Zd9dFjXekWArKcIjcbt/5cAVECfsZBvgxL14MrhlQWB
wPcX437sIWH4slBZJ2mGcC34kggtsCyPK9Vm3DOKTRctOn/ozusmU29cq+ym
LMn8cwXOCktqToqhMF0kpt6XBT0qQZLlgpbRTBeV7FSnuNLT5QnE+Oo/2I48
Jb8zG2VaUzWJABqVYEgookUDOspYCNLQRIELeRLZ8+zsb6VF0f6PfhAQP5Xl
hzGDC2kVK8s1H8b7j+rMb/JbLLjnRQLj+dUk04Njv6R0YjFpC15w841zBUiE
zjNheJyvwnuI3WS7HxONu7L5no1kbH4F5RuKKFesBtY5MdmA6M+FMxV/yIoX
dZbpwSAJiEbnlAcBJKCnNvg26Ws9LBB587MMhV0QypUAcFSLmX9JjcQkZIsc
lZjPQtL65ye82MNfPsNnIIl45Uh+eJIF5B5SZJEGUBionisvUKbx0a8iJa5l
zO3KdrephTKXrsTn+6e7ChhTz5H1iblsY5HpMCcoS2SNCmj4aiUHFWgcYa3E
KgAZf60EGtlxI9TkzNGQK1yOgYGAqzLSWn9StZpTgJFE6JQcnJMtQ3UMW1fv
pkgYQeHBzXoMJP5mJ+Bmb/25TuYFNTksWbFjhUlvVgMqDAX7z41RM2k/XcBU
b9gsK7O0Eu6wBzEmsk7UUbD2jwddOH+gZrNtlzRb0AyMO2q+mRohx1aN1YqX
PIL3v+yov265C4J5gvX79v2s34BqzE229GwnatYRWOkQUKCyCeBFnZAhKiQ3
ibXnG4KDDAVDPQhw2J5JLU126y4khFVsv6EkoPyc5Ktf4xXHYI1SoV1wZowg
m6YlYMIRX1Z3rkqmYxOD/cn8Vw5NBZiM1E8fyZ/FIECxMW9J+SgV4hkBYR/v
a8WvHHdN9A67I+wUOWhCa1ti4kuMnmBNfn74U6wQCaTQ/dSjtdAy1Ujo7YI3
+x665KmuBZvtqfvguvVJElHzbJjVcq10XuV3LnT6fp1TtkG07CLo2HFUplNL
b/kxw38lwEPcMddBibHh59XMeiCr9xzTMBmXFgoLwXPt5nM3ij4vazlUw3Er
vERpGCu9Iummm+Gz05CCfk2Ag77XED+hDFvEqgiCMjx9DakahyfY7asK/ZKq
PW/07ClHyZNYWjOdFjKoXSow6iPtK4iQ1ITNqWsn1AuQ32OoQjggyUe7NYI+
3Ce49enAf2KRroQs3rr66roptEK2BAByacj5sAm1R5d14AUikQFSWsrgCtl/
/50NkdNSra4AnwRC26frN26nYKqH+Xcl4zerC0atnlfHij06wm8LDu3jswWG
0hLH39jI6lI+Kd5NNb0+RC7NU7DkPIKtKU1SBxRRLHmL1cGhbDMZ70+l4Ghr
tEoUA3Di42WiQ1Logq668q2m5Af/7b8D1exj4nAK3/5xaDOSfJp0eUCw6SnX
lU5CcK0uZ9TbYmaPsIUR/u+HUpbA/T7cHn2C2dt4iFb3DOpT6BeZb8WXtSGt
Vu175u2GTRFNNJEC2mJdDlksDQ/mDuX024cRMaA+pYi1EJdlGGICZEb9V20v
zd0anCLzDvYCen1yr41txuaU6+xvsGQWNIE46ndaPQrV/nzsG0qomp0Qiskj
QvSnMQvVHnH31sVmEQG5HZtzXLqhoM/M3gNj4RosrJ5rLdELM13UWzBD9YqW
v0HfpDUgcsK+NdU9iaKSxkkQmiAO1VYfHLYtbKAo6gWvkRDC8p45GiETkOJu
QVgRlyVxuIygdsALJYtLddLQf8c5y6pnJ+6i6BwtBpKO4FkdaYAG8wuE+fEF
QSezsthpbMDo0Q71H6bf3mkf5J/5jGzrrwzGefVpj/cWsx/WOHZuiq/cOaOU
BaWdKae3QgJ8HqIykPT3Pt3UdjT5HnVyX4zpvTPyspY7jpOPnO+tHM1bFzGD
msrTwQvD5Y0WXC/EYMBmrzLyj9NQjL0QuAaJPXw7DFBBpwaRoOKjsJhdI0ix
NNeHZIXWitE2WPL6np9Wfykeu54x8mD/+AhxsvWlIZ/T48qpdUEfOYPKtv7x
4JdfVQmj+2l97oRWIsYgblG7EcBsUgcnjs4zAlhDqXFxe8EGCft+GLRoKUPT
I0PRGgbWPnAllLRuLK8R6HbDpr/9nKSGdH4Jj3EeA5h7jert/DBYH/fA5MXB
mqzw9WKdpBi8I7+RAeLkkNLmf4uXUlycsqpC1Q2tI70KOcjPTiIryGkLm1uP
auvNQC2gIqM7m+eb/08KPXoOX69UHxIVr8zycVy+tcmpvWZrquYoOfmd1Y/r
vtXZg9OomH61uw2qQ+sBye0dD+ZyLRA1dUL0Pd4q7vdkhNYzZogi9yLzcoSf
y0absz8odxwd+vbr9VY48N6YTxAXTUSKhcFuogIyUKbf0tL9xZHGgh442T8X
qesrnJfpoTECnwCpZPZ2lfk/aQmTdquNy47heIWf8V1WSApThksyibMRAT8s
l/IsswQqB9Zv8NNNj5YZAmUxkSTsOQ4PzgAxbjIgdmuVPB3TfU1jb/VS5gES
n5zFCjzX/7AHNWqt5vnlsltOc/E8IwigoQ9+S6ySS8hxcN9OD8F6Eol6KH6R
/smQTp0FRQZ2mqlvcXY9LAw07+5VBq+JwzIhYqrHRJ1BX/WRrGxuJSN/PXUK
55sK/kmLWkW0mzxZ/XsFHfgmnt80mueBEr1PdABNS1cy6uY3Rm2e9gHnc5Mj
XK1w05HyOqvYxvAF0EyWQ3NZYpZUyewhvDPWXhrCcD5P/KHeXftw7IviTtn4
jgdH0Ciru6CMH/g/k/+8+5wAlPSBTzWqat2fo9B77rQUZIcd+9iywcXJMihv
AdHCoeOS/9UOm8P1oUNtIxAA1PZj4QHXrWxm04tM7WVpTOSyqJStrAoTrdzi
8IBLOMIpw4LuBzyqljhFL+HCfK74LhETQAVIC+by1LGwH9qKE7fe8m1ejAQs
e3LGUxrnIOsK7RYTKKkju+C+nV/H5xyPUdOQoSWZir3elp1J/e6ZSGCeH0t0
xNU4FzFSzWi9tbFFXdTZJed+a3BFgLnm8Ddvny8Kb0wlrpA9SHxrZgldnBFG
RyaVFQHCvxw3X2skZ18cEH6pXbvPIpCTttqNoJRXVVl9T/Ae2qHdPF5oEgGd
XGDF6fS2GZUJjJ3ODA/YJrhGchxWnk4jbs3uvU0Y6t2k8nv/QlTe2DsAhN1T
4izFcKLT+Mlf1RrEXIg1l5cpahr4XocUs+3qdYg3a1Nn8hWXn9MLOdnDW/b3
iwqQVb4X81FGPgbBlVJm86DwFP3M70WhkH9CWrrdx4Y2sXZAMMNE3VawAgEU
jrv4Ko1+wuHTyuRb2YOBgw1jmbZABCIiiW11O28dFD+Dvy2yYZG4QQnVyJLu
JpwaHcpxU6tJn4xgVX6Tygnj44xGapGfwaduOOjBambO4tsUTC6ofgfswv1N
Cj6iLEEPZO65I/+UQAG1ud4KbJVC3SDoUKPpuS8UgH+wnOuahPfAvkzdOnzA
kEVmuke2esdQpIelvaWEqr6flaq9iGRXXFEs1tMsg7ppGd/Iz474mWjh8F+T
bnxLlWozeobopBMSSoQUzXvB3i8Ev9epYu6gHYP3i563eCiawD8klr+BWe9t
JyVvt9q3KzdUeKX3vKC7ecxiH/qKE/ew8fiIg0IzeCiv/Ahzshhuw8zRd3Sv
7OCwa9p/Bar/uuFsrHeEFTDW5ufjJFvH6PJvd+rrT5mN1ewKYtvWVLj2cmo8
NLh/dBHN4Z2xZjoaBEj/6f2L2CdqPV70lxZmlBOZiL8FEXiKU5jaN5svJgCX
YvDsnT5KblVce3kcNiSyxoePDQod7p2myiNiwOi7xLZqFolaLEoe6s2DplTM
431ogdU5H+fOjnXVdHixDHWcQB9iWXiVyL1W+h+OyiT4p3mcRd7D3Du8/CzM
k80fcDrGccLetu4NsdgVMi3N51IJ9QpfQniy5QqbjAX9sY6aAD3YCHiuAbva
VI52JuxHkgoPYYzR000lR19Dtj7C6EdXio9zd5GMrelFpRv5TUJ1w5JZCJz4
Wxg+ZskCEvulUqGbrtovEE30tjOBxL3FtcmDKej0uuMHE5SZrp7UJ4h94bk2
e+G+3/Q2iLG6z8wcgWzkGHJQm62Ti+lcup53q1RAPhZSKiM+Nzjjs82DnPyh
LJRtfXEj4BWd4RaaQCJGLu6MnciD4NY2APjsoPAqFa/Ipz63cfjb6i4K7iZo
lW8vwDbglCYLzgicRGjhBrXPEMefHnEi7JPwBLB5JsMMP1mbyCXehGMOSqTv
ee4U0nLJQq1iKgy3LXTCEE3eandn2RqzIrnLwwxeY1XHahlARlZkVObAIIwJ
6tqe5WsGI18oqnCZDfljWDseDRZdBhS6gR0FnSAzjQDPh5eV65OoD56l4j22
Y4LuUzbn730wTGvucEuAUX+Maq7K+1r+WLSpEOtzAYebmuU2dqSHFidFE3M+
gWZLxwG0dKXcS42Tayew1FmT2atBD4er87w2xWxD2s8yQQ7fKV7yBue9/aCo
LwSiFGz37WHMYEO8kCHbUmBAZQn7L0LlbwDLiofX8Wdc+tvv4bERyvClQL64
7g9b1d7d6f3tXoi7/dWiQz/jbq4wQF0AY6GfVG5cEcb7JqVBGvAj//c1q8Pw
8gm/7FEMT/hzqA3Dgn23Y70f8rmCAvaJRz2VmdS+veAucrHdNdiao6wpOGvm
X7lMyCQuFWMnyukDEbwTxDQ1Uf2nYiDU7D/+i+xrHT/LplbUpzEE7muLUHjE
kzK3dLXWcABL5i4l1xlv5OK62KNuPy8Og7Ecm5MWWoowbsW7P4IuAA8vgF6a
ToBTMtw1kRWohGggkTD1fe01LnH0XlCdHUhfMm2AqKP6tlDnmMelhj9zJDI4
YY+95Gn68ToGr8JMS8ewEAO+7eSrxMR/DWx7ufTLUSBTF6Dca8UtN8KQx/43
Z43r25NrkmkFVdhu2hyC3t4NuF1ToukCAbXUsP3RUWFnr2k7waFTx51X4WEU
K3N39f26d1x2jrUIFkSeDMOqx7HM4S1KiRTE0Vq08n3MRKHH/AhPgl8/DQhY
txTD2Ium1jBwp9RhiIN299OSzaoj7trA1vg0TWVoUD+/eEYFw4+bg+jxV9mK
C2EeCOaBYYheatmH5Ie7ywvDoqxQYQNKG1NTpztJQWOtoVJ3KZB97qJWOAFB
aqJKDCw2iBbMYLQzzNeQHSqlo8pkTF4LzhVmbSUvi2lpuAGkbJVEywkqaRfW
Bv66MPgdds+3+NuE+ootoQnPGDXXHJf0SSjsHnyPoD0XLUoak7cpFkzP/8Lu
KzD1Q4bTsafWPH23uSsdFdRcVQDeN1DC8iHUfE1iu0GUOKJ5cFJMrSNn91kj
lnEJqvinNDRchgyDZX7ukWT6AxAzdeLxPpUaDBfcnSmdQXR1koyOPpBbLep0
Ove6X7vt64gkWz5KTdBHWpkRyYl65L/qSZuhBaZPq4XfV7BVKdmjpCKX8+/+
zbZZgLgzyzRN9WzTn41/Rq9XAgSibd+nIq35TH++rmXsSsTcanc8/uml26wQ
Lhac9mOWKf4nR23Q4uffO8nSa1zg8EEInUOjYP8u9SNCsBZxeUWtAVVKkeBC
gQ5uqsYSDHGq905ijXlDpT8x6NcE/Y8CsU0HNKgtTbRnsUeVQ8+b/Z/TUjJb
9dUITPijWZI//DSCE+OYNsLcp3kHHJ5jGBay4vADPrUrBhbxBIo39aJWtsvv
NBfAefrFhQxDodsiJrTsKnYg3wPintNdenBu7rm0VYsQob/AYVP7RK0k27e3
Fn4MLLBtI5q/wDHqwgABxc3xSjjkehEB97Md2A+I2SbYCdUA9gQSMGcZuvtc
hLKSAHq7hGTbyd49Ogq7V8bmmdwuTIy0RPF7MmnAkSc4gBrBigWoeDK3/hKt
f3xqEdnhs2D35R6MBTx782gfbkklFkhIp7FgmfpQJZ1b/AITk+WZMWeq2/cD
DC6tlj//PfFd7mgxgwrMVgZ1kl03fWDCBE+tCW3FM5Z0teKlQtkfIH4OI8tt
hkpQa8N/HXWf7rLrnZffy7Y43SQS5iTY4n7EQxTu7+nZI5JCgQVGELnE7LXM
aAw4aVzBWyYag43S98Sy90fLBJynNgeTwCHS+N0iul468f+p2H+MQzATVSkg
qDgs1k7rDGgLbUCDz23w4oITOSRRYGeULiBDMspg1yOe6iBSRKqQtmCHEhgk
pfDPabyO4RaUqi5wJ3wQCMibxiPDHJvQSaKI/LhA/iG7h3lIP5g0A1BtffH0
T9KgUwB/2SsOWQmKaeM6EgQOcL6qZG3JmToZ/WwOQ7I9NSBoyQ6MGK+zsyCi
pfr9gUNZdo3X3XDOkr5IfQvk9kwRc691V1KX6DbZuLdj76XTAciEuozYEqBX
twyVzZ1Nv07u2KJyMw1F6zkGWtkq1uLEayk3qNEA8PRqMVrolUjOftIwjUuG
22q3i/vKXDzkkBc8BWrd5e/1E8fp+qkyGarAKbMiZq0vi95wTtC9enJmmfru
1lfgGKmYO/0wodtJMvysapaTx25kwD5QEuIBIdidoLJgML/Wvu/DRDR2WowG
OJAichcRcyuuCXp9ZWEwQOqoI0xyfm4JmATJAqGWlEXJ5LLXe1Nh09RF4SYO
MTKwSKDQdSHPEMhl9zofhGOz2iukzSjSMCMpg0GmYcR+g5J5tNwkbqUiUemM
Gkv0ARGX61Cs/920YzXXcwakHCiTyJFuI0LRVWKL/SEbU1848RiXz+39xbl4
JfAnBY5J9zIdL4mreQwf8VcZRIwAtHpOxuM3CZzIGf73tXGA6KmFW7vAZiq2
Ou5Nu1Njn1Ab6wXHtLaTYo079xFw2oOwXJBEjjy0GR93pAvezWSQrNRAWR26
caiJ7VXj6y5KTSe5qHAk2G0n3WUhQs3qD1RHzMhOtGyOmMrqiOWKD3wKvm4x
mdCSkFgN5zSVZzBEEH7GOUsJMzPiNdPgESJlTIbcv58PxnuxKPvLh3VeJ1Fb
EsWYN+4krYlN5mklvCZgTRGlm3EGZHnEhKoVlYVyo8NI1HkqpHE/rJUSppVu
MhMJAASg1i3ost47urGErNgAgHiOYEu4ImXbr+qKDCdH/N5kLGS86f0XsO3Y
7nrc7bYEh7r7AVVwONvPwLqzk42uDbnJKq57Yr7qluxQTzDsoPHetVxJU9X7
xOUNd20LSgKjhy7QgHpaIFOx9rmorl5BpH5EUlO7MGtxjvGajs/GMrtpzazY
F8Fa+sH9G5DkUkbfdzkOrew2/lo67AmGOEAg7SBvS1tWNQHSn/dOBjGaSkNf
n+Ovgf2YY/3PyTeYB4ciuwoGS4iQi7y8shNJZNp7gT3BP+5HZ3YLBwXBOuCU
PcOIZgnBgcERqbnyEJXp5mn7cieeARv3zqvC+8g3nnigTQG8AdwCqQDg4P0B
WF5vOwupPDALhGTqBGIqNqH2ru1SMip14vAlx82AuOblQ5SlaJLC3J0ZSUsr
KdkD3phXMq+qkc4mP3bCbiPHxqv7AAaImonYxTwmAC0DjZv0lZOcAbTN2eMt
Tm/axfKTtWPTKmHDG21DUQzcMWXWeLBu0DGVMrfIInGXdIyTnrKpnrgSObA+
Vuq+rNobsO0FxH6PDLqURgkKd0kJYYUwwhpw6hu6DUopbpAZhsHuu5sTH1c7
NHL9ITudbdhwuJ7yg/i5zqU6DjdL0iyWDUnDRyUt1fXNs7CeXo3Ai9I/8ByQ
X7NkBTsUZqziFRwbZ2Q86bqMi7FsPtgWHMXJlcLAfVv8j1QhqOC/im2qKYYZ
YLsCZM0w9Xar7S+zZBnY/1ool7eSJGS/gXpntpSrwl/pgY+GJHyaaNTx6B3D
pXUtuWdTi/ef4RwE/U0JxSFt+XD8UK865NZ8gWJL0664aUlEkc1U73h/xXBm
3139YXz+tkafelxkxy70bVmmd2RiGLFSPbpJ91zRVjtKg3BxKkLQkh+IBF1Q
7r6fPYO0qJeYSBIR3tBw1k2pvNBaUU9jI1dOcw4wLbIzx1r4+K5jATSpQqft
dqzd2q0OFIcGOSTMk6BENCbzbjZrU80hlgaT/awO/yy4ANYdyYYUXPkvA6+j
QJKzFVd4y2smhPCSusptaSA6owK51prZPHhZH9ZWwZGfrbTb6Dn1WFP8Qooo
z27RPbPtQ0b/ZZx9RDLAS73WIRgpSwNtT4Ka04+COAL3PxNIO6lP3jLMOFT3
YXTm/4+z/eJiA/AwyjrhyXYklfSvCprQ2WILDdUmcRTqvUE0+Hb1dHfq5eE4
pdRFeFkHVeP9zzly1MkHUMENDAi/UM6iyECS+FkCJnJS7gHzoAMLKv4vhcbI
MffP8kBYKgIAL159O2DTJJIKEgOK6j8cY8srJzrlYtVo1NMvQMSMnVxEEVc8
1nWrml9X53J6ZfFV9jHnVd2z/mw+WpOIroKBaR75flHzzRXVDROtEeU8Vwq/
2s5PUL47v64VHelt00j3domZ8/jDy0echR/g0CA+EsLHru/ODb0LbwEM7Ahm
11JwkFkwPZK7CbyR1MrjyUPGyPdIJvEUzJP+sh8DYry4NyVAF+QYnMrytVvU
Rirp1xAjvM3fBCl0d94dBwJ8AXkp49wBZs04S/ewTc6/b/KBA9L3zBQ2TFdL
Q+CmIqc/xLqpAXp7X/Keow3ActFBAtHMYB5zkRg9gkaPsNAvkbS1WuwWq0Ve
csVUE0/08qenaI6bs5DT52ozIu22xtS7dXKsNxlbQkx79N27puoJPzwYdN5a
HqkUDmtk07zXmxzgXS010xaQ6pNcBRAjb1zVhdSgl4ln4aFYcYj9S5XqH8jZ
FpTtzpADx1Do7ZR3hirneVcFDDSr5um3GbZuehsb+/ps9WqPqOb/4VYa0m58
XcVXrwlMZd/46/dVokqO/mgRynqgoSMSnS8K3WMZ/gwKrI6FsgzyWU55xbXl
SmoHdt/IhVtzU4Z7KrYV6U7FKqcLTt0unXlyY0+BWVGSluMMW1rE3dlVWLPF
gLm89seMeFXcU3eGOd4jB82OD8A4Q8UbhwWMkb/u3OHXfDZxpIf9asxzjclK
37Kwu8xMtF6vRYkHwzBkUx+PbjSHM4zNsZC6qXchQUSdIPg9kh3UJxygTO4P
T2L69nTDcTY9dKmsOjvJkyzTag0kdwTleU5fRcydPRzjqCQhnvh9ybIbrzXs
Y896SbRSoZ5H+rJIe56DIvBUXvS19+/Up3E5zAU6flh+vDgwSEy96geaCb2b
CDXjYnKJj6c3Ryk+Oo/0AtcCHzIvtngYtXjyEPxfzRcnRterfY54/FU3y4Q2
BQoK12SkcH99TNgdTh5TkiaowX94B9waRy9Q3FtE3n1BomzmXeuj9YaoZLUL
/Q36Dsg+DzttxQoM2hTV8GY6t+iHNlFiBgWNTBO6YMvhbTt1LoFzC57LhMxm
+DbOyTqZvDOLrW+CkSwtINGbjf+XzhLJ2/aSK7GRlRd5wP5M+8QEjjSjvAWf
jsokvanIGZbHHgtQqfAZy8MeKuRufZal5pmBYp4WWROMgQ5UWHhFv57SBT9V
MIyAI1U+i8xipCKETGUA/RqLhg52BsZOk4FzjpSySpdrEYOGR6FZ0SfDlP1j
6pp46VJVH586QPujlzZKAnHTzGdi3+OaKZC3JWm7CZERad8rFBWaz6AJe0CE
ef23bMqpI3EmuiDC6hO8zQkl28reiLMQt3Lt2X3EHnUSMFFyLQWIS1FyDe5o
hQwpnkUvKkIYkoxfnLCDZaYVfmRRQS522BDUaWcvKB4cA3ho4scYfAWkSauK
yEzYez3RZWakLjK/aCWtFqKNRBOdpea+Rbv/wcym/X8YT/u40hd/KnemU68y
RfazAilnX4L9w+gEWnMPPQq2iEamg0jD7sQ3SvvSs5pRR9651uu6eTV44tgG
tSajyvZWbgJn/Us2WgDSuj1Zl+rwPY9N3Ru5LEq+Jrqym66e39UjHkv6Atjh
wC0jNiwoDUdErznBo41T+ZQFqOdWzuPS3yUE/ww1nfGDr663pvBN7YeNQMBG
zJkVsQ1PWMK4Dfywcfqa87uQ0ajUOENPW3ppS0u+2WzifBb1kAnOIjI7DJXL
722mzj0FnKwCjIUcVqEEVGKiPflGBBcA6iBEDfaUOD6BzQ9r0boWZ3UGdY3n
+4wZy5lJ9rucOqa+RAkSjCG8sRsVsimKrghawnVq+xH+1+wTLBjh6IcRi0vr
omb1iOViTia/jCCsiA7kFAeRaBzE/XaGn9xjwECzs6VeCeae1zyUtg1N+qjM
cn71RH2QIysisl3b3QWQrUC3Z5YgvcbWVp8jb8XgA4HNmsdi0QpIhQf2f0lD
w66nPi++uK8wf5ITbJYLKYEMHOXQgTt9+2qnMDXJ/TfowjKmk23UCgyMNU2T
9oSn8k2NG3dbq2UJLDCKD491OHkdsJqRaTJcDanENWZNyE5B6lVenV5c/79s
Jk5+QpAJh/Je+HIfxD6NYQPOdYqmuYVyF3T3GC5xgqsNMZj0Ms9KJrskxpRU
EkqECF2kFlMz7T5/P4Dt8jfRQm5U03JmaBEvFZujY3GCmnSOG5tVS951dyUW
YE+KgY+/+b7A6pSVX9659xoNHadv36SiTjVTQksz4pOY+fwIwWikOUfdiCxF
uuvbpTvMAzi7AaGTnKoFkK80c48DfFG9oHaEP+lom+1XdWdNUvoEvAIj1Imx
X0QppX9iqIO25tMk11SRkFHpzVwp8etf1Pk1Y8tua9WwExyWglPjhCAwbnmD
aeJyMselauMNCc+lmR8x2PP9IC3HZ9GeIkwp/HtkviumXztoHKo1ECr+JSb6
iFQ97HYU0kggLvlv0Ai+klKqblWDIdhxO3620kw4SM1MjqmpVGCcAdoAy0um
3Athcr4zaetRL3GckvTeEYvy7R1/JYvYbCvL7JfD3ZR02ku85c1vNDRsyzTa
Pgj/WGOLrCrFOi5jLVSxUYkBdQBugQi6iQmWRFezuDpmKXtUbbvH7e8tw3j8
LftvkKksgkARobTObOgX4RaJSNg1TPFTFV9ThXdzoT/b8vq6UoWphlmjc5Se
uIQDiiFG7yukltfkADGtzQziSQQaiuFF1/GgYm3hY0K0GhED5N9P1FqnG4ks
6iirevrMyJJqrJoO9JCLgmijrTJwrCItWQQDYPZ6nAiffnAhBlp5f0TEB8LE
bkLXeaBSDsyrw/BqmDunX/z9Dbqdg8Rw/EuNYQdC0DQzMnt3/gmjnNUtc7fV
VFlRlDk3/Xcwtr+T76ARfIoU1o5jciyb6Wut5wx2B0LuygkQgEopFvTXOb3I
53hgs62hIq1IRXIlCi6TaWGEWY2nyt9slu8IeiswMksALJQIjvCuOxJ3ml+w
hxwDhXLZ29F1LwPPy/iOnYQQcqz348NMQ6KVlMvufm+9F3IwNtBrSJQxKzbK
LedldlbVg/bshfeVu5IlXkYPnA08tK6IHz0AbthUSdoMCZ7i7j19w/rswyaL
qJuTMnupj28eEMDumLaWzYPxLrbLkpnQ+NbNWNOicaag9O2JXKfwouJPm7st
/zvAWBRbuFwiLjduf1/2hVphlQWsmb2B6A7dVQg0XmkV9iiYetvocnsA9azd
L/2sHooHrdYyy/ntygltp3QwqMehY3Y+azp5yGorC/EWYVOELD3Rmq7Iwjm9
qzy18DYIHFTTEJeOHKtcBAKOcb2ToFMeYLmJXC8x9BqgTVgUqvwfU1bRhw3h
frbZGBvhk9fI0YvwHq7BfaJ/4uCe5/NkfAUCEr7bupj6BnX8g2UMzn2ZjXWD
PcDzbBQAWoDCx9vIQT/lFzY0gTFcCVUTvHkLzbpcZpSe9KZs6RY+zrcxO0wg
dx8pi3jAd/V3YJBau0hr2ikZz6M3LEluOrjzWKjDTVZYy3+Lj2ucwif2awsd
6A01WwBai/jx9u42sT19fu+jQYhfD3WjzxdwOLDyNdOI0UM542BmTOUwNPFW
kRN6Y9fHXtiacjt1pqyJYN+d+ZCNpJsR6JABpYt1rbW2jUVcfKbWTIB9tU+9
zlnZ/b5aOsEeCl25XBUIb3ulf+9cMjjBFiUpad7j7MF+0pV9IPUljJ4tWTH+
Ep9hZZORZMegjN8xuhq5DXI2Pv5CqSnmDti4TZw8U3ez7mAKLBusRh1Y1bga
2gGJ57MS3ErJ8irsgYr/4kkHbR8Xs8MKyklJZ4to1tZ8oLHe0ko/4K5vsSdG
94MqNzz27x+Buo8Jb95gJr2y0i9Wka0Ql7mQYeKFjfm5kdEfHJIzqHyqEB83
OKt8sMIbu0s8xYsR+V6LV2e20Vn+3W1wBdC7qdqHGW73ewu3p0Yx8PkwzUJE
uhF2SrDDkelEpqxuYTH4ktCFwbo3nicP1B5OxoYJ7TwRqhurDkephhbmX7aa
W4VGMblBcc3xKNZjx34wiH8023wS0YnRtFjrEzLA+RN1IBY9UzUBH8GlsemY
a3TZNsD4r4fiZAa8H9bk8BTyYBlqrwjlRLh9ngMPuxuSlPQT1GOaqnM3P73o
xgawY9a/cUUQNfJRM27HVFgGvh0UDy+pifxLiHx1U5SlcsDFtGM8w0+sej1d
er9xDXO7PTMUN5sKxThRbzcfxHCDuffnMvA0uwqlqNuw5jAvKcz1Fm8pOtme
ipr9z2k69D5mjXuWB+8YRYfGLd81RwyNtLVHEQrRNp6QpmMPwj1qPJPIrAEA
4nUKTIFgyIJ5fyW/+SS/h1Z9UUP/KRQvDS+GyI96FHH5K+0iVqYywWkiXuku
j9wMy48D15ZoRJMryGSFwftZQkYxVbjh89+YydplGlbJFLKS8qm7TpMYFCTS
pBy24d0hlLgfak9QtZZgJymIgc2WXjhxbZUM7zeNCUxID6IHUdseSYHcnmmo
7tOQWaqNoMF7pplgpVEy6sWEMy8cKcJwjwRcW4lE9//V748YMdDfuhB4aIQb
ISE4ZOgtQxd1HSyWvREBtFkolZvSq7dsCMcJlhGVFvjtjaY+tywnWJfR9T/W
k0ml1yhbIPL+48DaOg7MFPIAUzKARgAxpWr9SVqhw78zpKHFFep/sTeBI/ik
WE3B+aFwSeDDu/T2oIv84VQ9LMdHdDROzM/9MfcC6Z8rkZLigA0al74HHIVz
4ptjHmh5aZNfFwdbNBq3P0LZCSklj45tYZ+0CM6+CHfZOI9Mp7+2c2m8RxzS
1RWz6zoThUuAoVSL6I0IF1fimAYgor55D61QQoZRxb0ls0kgpx+K2vueraF3
iyUGgI4gxvs2e+gJS61jhisdKc2AO7lqNVI6fPiJb+KmvQGAeN9DUhTv0tZj
hJCbA3YKQL7ttjH5h7VPcT/1b/4heHzDxK6e4hJK6YyYaCN2iDD/AgoAE27b
0mTd4qGp+yxXriNkk846kkfdZh8CbGoTmEL+U9WrdoQ5DmXvCh/TyZGVHl1p
BGRONSeCABVrF+P6oXttkFH2QVTEppc9gXf12IECbbJuRFCx0IZqN7S50GnD
L9P89OUryuxn2gssrccK0zTfPAc0sZ5bwRjjXv+jEtD2Uhpte5Wf90pT1fLq
hm/clZFhJdNh3I5yqK5rDLxKH84MSa9ehV/pRcRnb/xh6mU1h1FCREwihrXm
pGQWFMPjmSX9RNXnxHb6rFZgv74bT9QhO6Zs4n4xD//2ITixCjwFRWrblohM
jhgCDS7XstqDB1aGqeuGiRvU0oCAtZDkCe1Dff40ByADZgj9MHk/S95JZpkr
4fTCFqWahjsTv6QzcoXrAELWMq40cHHBY50SqzKz9776zdiJLPpkcUTONN5n
J4fa/eSG3PWJM1oA95Yie/caQEuxtiOCWRVXN0aZDfST7C+7R95LmcTh6zTW
AAudp6sa3gX2/RSBiq1j+Qr7lzOuIOovzo6vtLjw8Dwg0TqMLTWp/UIuABwO
hNgiv5wHsMYweiyrCo5XbVTy84VVCHCTSRYA2jAmNh0uGn5XzN73Rg9wdNek
TK1O+ekNGf2lpN5bgXPQKhlVMeFCWP6Bs0tsgsy6mnYHDDIycwtrjnk5u4Wp
1lChK3AHvhiJLwSOLnPrTU9yzKCDsfBsk+E0fvuX9B1WhDmYyi7tpjterC2I
fDFBkCgr6D9JVDGYNv2DpMybMZOq0U/5YVk0Mi0Y1uxQR34jdrcwOC09u05V
uQuR0Cik2UZmuHdbFsjzBeegJFjy64IBRhbaus+tiNiMj99/x8PzOy+H8/+d
v4JyFKXyt5CSgYmfJEpWbPyYrhJ1u67YyYVYHa+Rfhe3kf64oenDPqFSWb60
7f0st+3gHPhto0ORO4ctnzt0KxBhY4WGJOF6laekGTSTwJpo3AGJ1DGKWg+o
1cobcn1c7WQmg+yEywBlozVy1qfu38hBfXfFUOjDCUtiN0KU6S2TsjK/xLn6
ReQq+sYl1KmzRhJkDl/ZnNFYVt8EWeMF8XHR5oxx2MehiIY+KhMnPPhLXpNP
LCAJNH5WAmC4LpE7FSLwafd+UtV4ZyXMuCaPIKYicfjkOFEfBFEPJc1ScXpV
I0o8DWDPTCNYK/0f3tpJCS84+505d/1NDxrUVjK6icUxrsAq9QttibO9PT3U
mHaoBhcuwB1SINY6SRiL4s0khpQV+2izeV3RhJ/i2Ky4zoQsdimTkHf2g2IO
q+YSexnWp6foXv3ldTSmp9XwuMDNLmDR8fDlxpjGB3ruEBl54XKyBD8IYHZs
O9gWBUAk+7ssVEdTuhaUFAjZgO6Ew+99Pkq+nmWXOgPb9vA5+e++ACSMj5Iq
3kvfmMyP6FXvG3TkbQQEf6E4lLHbDbNIkGzXN8Vwu34ErECIF2/TGZWDzeZS
41ZuXXFyvGvNOVsPohyPhdBdIV0LmCrN5x40LKG2GKwbYpxxxc3V1VhRfZIQ
MwQWMh5Az82AxXeNKRFc/rF3T5T3aUmb0xr3WxFa7vGw6sf9R+Vfrtn5nUI+
OBWFM1sQ1pe87W7bC1wTJRM6c77HsWefBFShivxHq7Tyb2YFJFZb0VjwtRxM
eIEvzlBUtQJ/Bg6TRlTIPzf21VBAzGALI71LEHHo3qrp8uxIpUl/yL10je6V
pOBWdpte53c4y4g/D8xysnMKMPtv0akzLQfmG1LugfYtYZqm86ZrXb/VnOFh
Q2xVuo2Za9mjSg/LdSEQv2+DRswc9DQVzxGdf6rsLfqti9W2OZoyGjvH+SOS
QTqoe8jGVFXPYo5/E0qRDCz51zP/6kS4aAMKGyhoh9+I2A515RhpiR3hCqEg
3R05RAKVfKGoRpJ4SypYEVHpLnJBRQNirBvcOxvNIeYOYh3USLegNtBT0cIK
e2H7LaG2DcKMhOTlprknHI9ePjmtFtviZpsJ4Y/Ri0LJtDjewG2RzGyOM7i/
kqiJUgaYrvWBeeoSywZIu/L7xcNLKiZpVUqnYSyVUrjB6xI02+rJ2s3wnrGz
RwAh5kBUNdkdmaUYBJwR1h1kZjeMZ5m3ie/M4W0CsSYGa/a0hixxP8f56z4b
tasBbTNXKKjH63kfNpqxEOsgmdqz7OQd8aZRBCHY+5xlnp27iQDLIim6oLwu
HAIDPf2hVnOCbCffzUOIZG9F4TX2wiRasW1Zm6wG1TosETrrEjLSeLd/CKNI
W8OlL/ZU3L+fA61foRc79pyWLr4w00iGLHnSfsVVFmnF6bf8PzdYGatqq7Rx
vjjtORTBG3U0Bo39px0bUzz468DngU628SvFzYlXHXc5xXb+RhSp7WNWqqwV
okeCB9SzfCFcuBcgjJSnkbmaUVpd4NB0QNOXkMv3Qp5ILiLCU15XJ3ihzkH3
74OgRMpyV399AuYid2pxg5GEVEUIVScNcPYA2Mq6ETZiCuaNp+nd1eKd1K7Q
etzq0oPiq6Bm2Qevb0QFK/wlzM8P6GUod9gXZHpGdCQBCibC4N4LvftUnizA
G3YU/3nEjbSDWGteveOF0BpOwWlw04xyX7An0HbFL59aWcO6IefoGmJq6f78
ToLl69HHjrX7h7SkxLIXjNLq2/PyXCmQTus9hajE8vpU9oonYL21yhhjKodd
tU+/MCxuoPVSAJ1Z3cm2cJPY3DjqUCssodViFg/nZvm4gGNL7TlxOF58sZ6l
Rhup5jnR2kWg2DEB9Aox68ieehqTc+XM2ikkTc1P/FPAjbKT7V+vRh+9K7xB
XVDkBerAgzTTwuWfTcvCVLX15Upjtb35pU/UBMQ2Lkqa9MB+qPKz+76tNgDJ
ZgEC2E4lHjoWwv9JJk+/+uWlEax+JbEr6+V8+wpjYTves9ZDQXJPUuV4IISU
nAuJ3rqvqQNcODE+GRzVblu13QONjNoJfPNVvODKQKnzYTp9BO3cLQ6egOsl
i9r3WFG4vYVdKwOEr/BSASR9/zrwt1BbFsgERopOWlLDKN1LLxpfdpIJQ1WK
8IIslRu6F7Ge4oy2/rsn+fpqJuWgF0niSsyKcbuQv5pcquLLFaQspbv0cxG/
jyWBXaa4ThwafzMrIf+pCfVmBjx7o+ZJmH11G+AsVKpPLyW3OLAfk3+h8MrT
69CWvDLt/4F4p7ZBAVJd129Cb6yTgUUNgQ/kBJV/0prkHEl2H4agirTyqJhh
wpUqpmHs+A1122Tw28hPniXWpq+0/Z4Fz2+I3JENSNnGkud6i7ICMttYX60H
W2AQOLCASVK5XR/F+ERUAH02g/MJFiVSoQ2YnmizdIRSrZANPY+IgmKea7Hg
nB/emwYjDxBBR8CC2SaLN+jRPYG+wFL2f/naBCCNcA4Nt7AaBCK8ylb94+KX
6QwtgGe8H8Hqxz9pxZC7sIzCtct6TuG4TnZ7OJL/o7qsBjb9vnw6ZViu1Wgn
rLe5Oul0IsjoqX5PTfUg9u7GiD1JWAvz/ScqwvHyyTUf04V+urdrKXmdX+1B
BtF7UPAhp29EXUSc4eD0Idbg67LSG2MSvAT3r9k2nB45BssGVW+WNOKj0Q1U
DBc1ocAUOt3LII8VUJz8OL+AHSxsCmgIH+cPp1Mfye29HXW36eNxKOhIbMN2
5gv1k+dLM2OzGkNrpOHjDYA7m9iSjU42TWzJ84YyVcowj1DcBpOZDWjbsIFv
ll4kbd2LP5O/gjlIhBbVQebCHETsEhyPrbMx3sTwb99Ca9VaW1/akY4y8zgv
6a0vXbxUCSLy4hUDHcXGZd4i5MKQYK+hYeOtBLKUY6gVxi9LAIWf7/mSLret
UsfMs2gIjxl3CFX7nKq+YTU1JHkuGIB+kdekiQf7J8vycTEI4t2RsITqtLjY
oa2B3Dtoa4KvPLhxgLXEwZm7kjfny5qettaUso6vhUKjFyt2ud8Wd6GnaGP2
D3IaQEOarNXg/bDYRRWl/dDqHeAXq1BizMFZ/y4UrCfPbZPZXnM6I5FVNtJW
iQC/l9JaaUF7+VZQ/ZHj5JoeU79lWIZ5xrBgKdadRCMoFAsRzxYGwrgvHujh
dpRJ1jFnTkMGzf8EvtefZaj2wb5usX7dL/5cg/5Zj+xHC2WssK3c7OVd2pQK
CSeL0ljKVnhQH/PPQmwcbt5cdilbEZThGwl0u7SjEZpMRBlKZtt1bRw/GTLR
8ZychozkNWu+VDj8JlI+AGUOGc94Sj0uOPyV6YMOGU+eXSgUAabeYIpRyUh/
IVRlYTkFXKfLPSr+NpiBCs9P4BSty6FgSQ11w3PKsX4d50VlcAqzFh1Kc6Ml
VnXtSoRF2Tjg/JOYkTkmCQdhzrmXApoys4/LS+kpgbctvmi8yLCldpIB4b83
ywFVFaWiWJgbWDyIfAY1HbZkbY2x+6M0LuuHWbfZWNv9+Fk73o2mbo6k3idq
wy+UiJ+WOn5aFZc8Q2y+sXwxGbxXkZGedD1nSXQH0ziiCXJwVa1sMz+0l4oe
B6fksPbAFaF3EJGJkcjrAm0WpnIywS8QpP+6R+DnVmTLpYdEiAOPwTWDoslB
l3gTovuGE4QSuD67iJ0aNfN5qYKbIqi3Us1W5IFXmZNrM9r/JhVpt96ordZ8
rHwxxS36Sv0uhYox0462bWt+r34CeC6DgaxTGIAPTSEek1KqBS8vNY5wBqdS
g4Lv8DJNiYo+pgJKXRwUD3iPory7Fg/bJg0R1YdW/2m4a9VLeywm4hwxiUvK
UzovFs2wrksddrbLHTqejL7a34TlZphFUVQpxt+0QLQQHnDc3q+jz6yTqskl
OsPWRuFL9IJS1KJ/gsbZ/gaf/AwHDR2yUMWl+/WeZmkOIeFAL/k6gF3g4i0p
hze4uwIhm+CBmCfgCHNVz+DVJ1LGpu+pj/gJ+2xXJDaEfkcKRoym2nW1YQ5T
AP9kn/4igVMTNRdEyLGhwnBjKr77rjSY2A2qwfotk8CjRfPmddE/zzoUgcTj
+FtfFRK0tu/rDJhHu9lUdIAjCgtUDutxCHLYLMLhjMBRiH6HdenUWNqADTDG
SIQLuynC15L1ASsfOBNxgeBO3MCmwq67WhH2S1f0bYYbKeD+m2bKz6DpEN9R
5IKK2CuxGsNV8l/ZhXrux6YCkwhSEvz5Og7szVXLAkDPZ6sQ1Uu4wsOSFPML
5LXcy6robjifEBU67U9HwFIqVURxQUZwtmPfcRjCjOKQ8uEoCHIAlh25EnFk
CqCW6B/N2l30E2l4UELbwYCH2TxogLSGBRwIAmHChY1aZhFLin6I5uVavPcm
jZH0unan5U/fFF3DXJzEJf31uKK0wU5HWqIohmNXd7XavzdxMp6eT0MNMYSW
gVvipdonXKL+UIfX2k66KTQM3blFORLdufCcYAYdrC+f3pjY9MYgIAwU9wy1
W5Ax8CAxKuo8uPf+dBAQL7dwqu3gt8B61xo9i7iYgaRlWllu2tvAw6pyVGR7
lf6ZV1rU1mKBGWQ9o7oBiFLDoJvucOhNxQWubTD4/QS6ejaeNe2sp2B6CM7I
OJ2wXTScepazhPY273d+XcXBki6YqhGAgVpBvLijKVAZUM2bagmX+Jonsb3O
ZOnJY4k3X+F+rzTjCNnaWh1mj7qq5WtxwXb6hjWmKocoxCiAddF1onw8Z1VT
8GVR7J7ZFqlLSsWfZ4kzhbCeUhNVryNOQZ9pLqQCMKc1k5AWvmT4d+zH3bIr
WxoGqG/enkHZe4o4D+FpM4RyC9deZjM0j02wssVO0LXnUNeuZJ0l3M8iEgDV
/0tWdbgayATL1bBHx5lZ6B6XSNzEL5OvISIsrtOXuh3WJBDz4LwpEepoFn6+
n5WG4hQeZU0j/KmXwlbQ5fxTrhKqM3nJHgxPLiFpFbsgVhqmmjfQn7XwhGk5
/xbr0mQgWVQhx+jWejIakvJzuCiFAYav9vLaqwEENWCmaK5mPP+zyO1ftWLG
itmoowmJ0VYGGV5uLJSP8FZ+4eyGCXL6Tt9PKTqQhY6qJfN1x1nHonn0lk2K
CW1EdfQpUEHaWayP02jxiPSaL6H9dV3HAX1DOX4dqlIUGvFHYSsyL+zzly36
/mjTXRoqdBGAWEjkyOOme16LolTMBzIAcSqNrdcnujHpgDxhqVcl+5S6EHed
+v0Yj09tgqkTrhiFaUkxLHpO80gMNxTttOmcdZ5pn50EObPC0EUXNFedSHlS
+cbQmqRffAsipGrQQEBSpx6h2ckzRYfY3h49qZsCnPDCjz0IY6YUvkrI73IN
yAx0mveS36ssZJ3IAmIUTAAgqL2Fz83MuitZW8Q+BrrFhfpW01//jmLf1g7C
kVJrb+SLP8BMVYP+LiazkRqSycWhSGyTb9UkQK5UHl+PdLfWUDicTuo+FAoB
oRYe1rnSxGEIkFLWXwP0CoTqZT0+8SMHDnXks9EBeDF8QOFdqtKHAVUzRBK2
FROcbzlSjQLlaARTediZizdf9OdvN7C4Swo29FuAiGj1JP0W+3lsI6MnPNaz
OJ2C3Ro0KGjHPWOd/i7d88qUC022hvZ8m7y4QZQLmQL+epeBotyQ2ADh0WQa
/kaqc0zNDQ0tGKUCFtD1xwhycNxVg0K+4I5y5+ZbiDIoSzJDvyPhEo5jbAAS
jYX2ZfmH9ANehKQaWI5qqOciPO1t856lrSIkx+yIFIygNcyCconpV3c++P5n
1uFIR2WChsZMj/5pWkRQ/svcrKxfwNhkUTDKuzxlBeL6f/qLqAPpQ2DktGSp
14sCgc8FSaWOG/U2PMsaWQWDfloAlal4+PzMDg3EQ/VsASzfWB0oql/TrTSR
mC1WK8xWQ7K/k8K/nbbKT6tRgEgkHsnp6RKMEAfBq3f3FWoD8KsPZEboFL2z
NWjYh4h9g2e9EJ9J+Trji1vvz1PfrxL69W5+kxbxh5hJkh4wH9Eb7+x+JuLA
JXYnxnBWp17itLMRtTW1JO1FJ+UEYHLs4La1w5RC0cYWum2sY0qTq/B9RK0y
N6gWzkg20RrntZb8XOqqDuoG2U6eQ1kUT1iIToaoDHmLyfRm7RhYRiy6TO+l
4Uf89IBqMosZvgOfylQ0bnU1SxXetp7SIiNlND4m/phDpRAw/qOAyfyTbRDv
C6BN+K9IZrKl+Ecq4/F5DjO7RDiJf9DB206jlsUd6DK2J0kLoIKVgym2SBDv
eeOUnd/hs3Ot9a1zQsf5fJD54oywqRzfromlQugeTW+mXbj5aSjuGTFi0+xh
3iUWc6P0qd5dEbYEhQSFnIxoVGEpOMvsFlitgS1Wl+UfVv/AMUyoFcYuJfzL
5uA7x5VLJjyhUhSV/UpaYVYwq0e97/SgZNberucGwTgl6tcKP2WZeo8y7M8C
4D2MSLwV+ABoaUWD3DwrkY8yAU5dBjai7zknodao1mUIbQTob5W0lqpAA0jj
TDLkezL5RPMx7uarLiHSV4TeCewOZT8eE+tPYpA3IzWid/nUdounNayXJTQc
JOemVPaNOG5SqiDe2gJOPAtkPRtSBSiUxuYduhLbKivfQ4fI+LuhG8R+anic
B3TnAi1uhHovd4Po5XkYeGK+paI3aHLL8txCTz3It5cOvRffDVZtB9JvatcL
Icgn1CF+lvd31wram65ftVuFBDI+JfaKhUKTGmoyy/Qj5XqqwFukEOlks/qK
d3ML7rHp6a3bk1gESWv1Aj5PkaxlljwABL7FhveaYXz1Rl8EnAG9ELF5cTJc
G8OP12cp8w0mrCcB/n5cNFHbZLR9EkBDIt+H002yY6Fs25vg8wHODz1GQ/X4
DIBWgQ5Z7ho+8y+O363XYGNqEHJMz1bjtDqge/OSA0vN8aO6ZNRfXolVZRX4
PsWzpz9dGLwF6+1q4H7pL3hL0deIpBD+nHNBeTI6IgWNL3iEcQ5PDsq7M8pP
DkYIlapsYwlSMjd2WtpkCJqGrLraQpwfcddYDcHB/W0kufmcZnEt7hVEUjml
EjZyYNtsTIzPel8Ij+GPBYpFVKjowk3Q4jc1F/5WD8UHx4zFE0hgec5r3cmk
5kwUDIlN7uw9nZ2oqANRV2eglIdma5+rJLieOVH02xFf31qFthpOf6e+ZgP9
J3sIct8kah8lvW8VVYV/FcTKV1FwQL31fSAuNwd6Z1CiQbkm52xSPbOCUnYX
A+LTJwwBa6xdQ19+8QfOLvTIOnkWE3I6rcApAR7LW6cP857liGkAkzhHKdc6
ketMBjaLVCuXUKFJIhZU647dZt17oMLc8r65f38SkDkLImTqruioy43d5aC8
ktxGEuLqyWnzbjFpSqpEpM2jo7ZQvjWJDKyH5NJ8KGR3dGelKPcaAB497VMI
xXr2PjmHcbOlFeUUXRGW6Ml8aBIlk+AbblfzdXWlsmfhAF1HbxUfw4nZz3DE
Lt9NQEqTZ99IloFokro5NCbEzTMipNmYpwE/Qf+bZyl7ifmN1vpyW60/BzF4
jNxGFP9/a/V8kgBW9Z/bNlt3NLU1dqrMDWmLbiS37u/G+mFqE5Zr0qo+TG3z
E5oBoBU1cTbXTOK7FnUV55A1ZAr4qK/pYNUiSiliUqYU+L/HxhL2gPtRCDZC
fntqOx4G2decCTBu/9bxSiTQ5nblqVew4GM9vg4x2rGt7vDta8L2msnIWeOH
ZrCKP9+qvRpqyg2N3bURgozqiAaLmCZJDd8+WBvxq0BD0aAPIsTqn8mBsNj3
77x438ZSGFpnTgG6rj1KszuywTkmXLUU84C/eymq5mUIWxiArdA3W7gfd+T/
BKTxY062p2frLUGUuYlpSgEyOuPG++7xVZE+ungiLCtGjs26l8elCJiDlrsg
qJJU3q2o8S0ERNoLUcmqSfEPsKvYqN6kKNViDMiqrgaj49bvLH44jpOwrIY/
LPck279G0qy2Bv1fMleCfKpWRPvaAPSOJyyIPJ9f8XUeR49EjjSdBdYObaCm
C4+39ewrPvVhg0eefTF9WQv+ed/h+fStpFjDmMRS+e59+Ka4gP6M4ZNhi6JT
SN8S40eY4Ch1iV7OWVdi24jfI6qU6/M9Rc5YZ7I/q8oCyUhlWwBX0kJhSsEf
rDoWFFVObu2LzUfF1PbLSWHrSYtSqIpkpzwi4eto3Lqj90yxH+Xl4GHoIL6M
n17jse4XFLNjoFr7MtyH40JnW6uVn9TOqO1Oo5MNtq8P8/7o5ZuDV6XFojBh
9YTlczWSNh1tfsLdlGrLvzffnxBtJvrfpiCyGSzWsqA+LrmfN7yxB/DmaYx/
toQ4wx0RupfJvyQ87jsk4eyEwdsqcYQPJtA9NUjMqbXgJud8MRqL21/RCJxk
QZRkJ9mVsYlbmR8L+XK/qBQUgcpZ3x626oULt7ogaWVYz3k8vh5fwIPO1DgD
1TvcJSzEfJ2QMG1fg9Z02O423ii24sAGcDwNpGgvUmT2iEy4BYOAR02HSgbu
xSjkkgdEgy124CkKJ6oqzh2dQVNdTPoDN+vpIw4jfJkJrQZ9A2qsPjrIxb5J
WWe86N9oDs76ha3p5S9DNpBV3Ra3O2Ujh0koHiFnb0weOePLuJy3ASmNR4k/
3yBuWL/tSh81U7zvpA70kfnXJERG2nGTTLsM0DxaKn/5Gb5t2LwOFuRpceBH
2Vj9nPXyEpHFGlN3HC3/IkOYxcdgjmDOcwE7nrywOudVJdlxDY2o+7Ra5NIY
Whh7clGnmfT75oMBsy3j7ECXSck/FbsnA5CdTc/r8jGawBTSnH/2O6ETldGr
7ggfT/p6W5FOq3n5jo7Pqf5B0PFJ7AXioJDd302yTNbOs375bzFzObrfE5S4
nibogNJzc0xfx5J8KJX1FDCkld4TSpBkwrnXUVR/97oDMXE9Vss3W1w9iwH3
G8ADqJVNL2NMPJLtacTMf2CbLY8aZl0BHcHtWKHS++r0/FIYfe1jj8CgwLLE
k5iwKTidGenDLXLr0WI6rV6LMdE4WTYNh4OP61RBra9Ue0DwIBpyMilQ9LvR
JU4k5jv+sZhOy4lz0QGV8Lsexudv2ZwXqHBcxaw3dLCimxnnLHOdWy6yvsjY
Y3pvcucTdr50hyXW9zPhzWoAuTlfV19aS++hL/oQKQrPYOuxFRHmDCSo6FVG
2LUsTveHiICeEqInfgEYiO6nkDMKw+0W04cPh9M4y/v0TFpORsbV4l9nlFml
O9TbDUl5/P35Xygrhi4Q+GR15pMW4zNipSDA2pN+n64shwx2XeITPclhAS/e
7v/SL9bDOwXTdcfLH6FEm4s/oZrQ/BBPbasfSHWUvnK/BnF+ff9UIhd7KJNW
XzAyr2FlZEwiuOYBignh053GNvX2RXbu2PD6MTvBup0k1qSelUAaNKFSBPNk
tQ7N7Yzc3PrJ+A/JIbQ+BXB+oL0sd2MEJ0RzoicPJLMDx9TxqlMChqvcUmTl
TtTgRcsgqol36pWaX3BNi36CpfqxWUhOT3wASGTUDySMvvXo0j3dln1fBg4i
JFbxozXOqmpGHAejkr1H2HjHi5JyZtzm768xsL1CnwMDxCFqoTBXZ/wuwsv+
MWamBYQYECZrPkcrxno7wWwhcpHh7WHZeOiJ2oV/VoAK/gyM5jS14s2xpmtE
iRlPmamA1JHSOx7+EdlYHR5cWaRWZgZoHoPH9Lbf7N+9G15CBAgQAQ1dt33P
x4Q6jXKUEBc3xOguj5v98TfowP/CUSE+91R4Cxt5deZgePJUbETqU0jfUL6c
Gni6yeR7WYoqiUvGxpnZ/FSy/zFs6p0Gn5ADDcu6Rk2NIwLoYbOFNu+bZAg0
/fXoMFqSdKjOb0epX4F/2GwUh08X0/3tUB6cpp8VRlOSroaau3TLmZGK7ZMj
WX7R7OvSA1x4v8Inm1HZdrJIKAUafn4p9XEJmKxFLY6ZhroOmd2bwJUOpMCE
98DlztyC3v5u05UhrlLONlbK/mSGDvfJozxvRdDTwTP+pSwLuCJEv3lbd2t1
G0B0Q0WgEUyMJH22tWNu3tKaUsCHBezafxAZ9dfsUgDaYjdju6cvaQVHbXVe
4OG5GjW3r78P8fPnhYk6OKJQnlrk7Wj7LHk1fh6hcpu+5KXVFMoo8mdB+LJn
AmvEWjHt1p8vqd6pHMuq1R4yGiWacnasm0UU6rlhsdRK7Nn+aLIgtEmFQ/ZF
vAgr7AtEURu4yGCoaky3S97mT51gYihE1hkvozjDi2ebE5dm+p0gNLU9TgrW
cy9gmBi9Km/m/aHtKTu9773UXfmjfx1l1rekIkUMlku1k0iUpXWk2hW19fWv
/ipu/pMyjC/BVPe5ILbs2iEtFzGTOT4EzZdrlvw2XI+76xLiMwmS0TRKKOkm
aRqEQZY7Q35jTFgFM6XGKi98PAb5cy7dy2TZEnjTkUgMCusK+kuFACUv6BW8
D43GDUscFn1iH+CUwK0QCcbCgSL24Q1aLiEvdNvTG6L1vlfOMFSA5tmRM7Hy
VD1SFjy59qBWcI8Wc7LqHkA2c8Xi18dM+u3uHTm+iNMRBSSZ5QCOTo4ewS7z
OeYtetrVV4TVLC4wqLjFZZpz47ppyy4fGJt9U29u3JzJk69l3SSNSVeEpIyy
NtBvHV0g1POA3g9wmbesGPJtmogNVhutWXS++WacaKzB9xAmX5UD6+SyEQ4R
i7l9Eiom56MVTXhBtigSwuoO/+vVs9WEN5WZMWJUdyS6B51u+tQG3uVNilT4
rwn5FHZG9jYC4ZUkgtpJgjjrMqU7L2LUoA6I94kmn3P0y3zjbJIQpvshXbuw
egx1218Qeo4rriCYLIywxKPL7OdlTLITWakmhhkC7DiK7uGEs9PoGUpNJSNv
HHiQPE/aa/vaQB+iaLgKqySDAggr3fhpnv2NXe3+3SvzGtvjpSzDI3CA4bfN
8JNLa1BOiRJtVc320Djhi2CqeGFTpBT8z0ztdWK8a9tYEUdmkpId/8H1bKCn
oUoz4/yRltW+2zCdyQEiyTn3Z2M4C0XzxQJ4QnJ3kbaezXR8tDmoVcm7QwaN
Y/I3zL5SOsttlmqIZnvwDY7eWEmHjESbVr6KyS8/b/OpZckYO7HlI66mEUCu
Qy1Zo4OjbmqQzrtZJr2KziEkILTNocNKwhvK2yEOiNwMmsroAu9q2y0jsYpz
UHvhwx5c8JmTBfuf5Uw1NIGfbz0LHW0XYp1soQGBWFKAZqtjiBKrqidNXmk+
H9D/Sm/0ffJSm5Tn6oV2JZuQamcdsOb8cRFAv3iME9dEbrOq+N773m66BNVd
vWldHhV0Je3CgaLuWnyXejDOZSKptzbUu17WfMowYvAu88LkXi6SVM4Wmrr9
7eh2FSIhc00GCguGwdYgxnnBqCuD4v6vM3EBUrAL5DUx4luJeIMw2PhFzRRS
eW6f150lIcgdlmmDTIIHIT6wH0MSSFX7DTk2pPbS0QshmiGvV//m9akzL+iN
CZAK8vbl0avoYPH6f3XhHQwXmTR7pRyVm7v9y+KJhdulV2EYaeezRR0hNkK/
BOlaihPC7L/MKD+5OT2VkggvhHH/de3TlI7FFKQHMLREp9mKfGaxAXZ26ErZ
AQwAw+1dEcjzeKf0zYlD99qmGAPwgDH5fxpkZsiK9MwuQj/dHGHmVRnMXIvQ
LM9ZHTKCXWe0kQQa6omq5/G+D30Dy9NVPRZowYNzKQoaEy0xtXLTszrzV5Rx
a73H6HaBnPW1krI/hTj9npDj6Zldk/T55+uFjY4v90iAZBSluoiZ6lbHVHXc
08FwbLdQQzy61UJlV6hSXlhOXq1eXm9Cxobj2VLw8rRp/mowID4qQmwuCy7K
gQ01dqZQbvKoqFagJhswxthGhSOfWO0moFYKa2czIcxMMi4u3ON1GkUnTrQc
ao/XenEc8C68VKxpFiCLyLfbbQtpO8xKbtWKS7sBXT/4K7YOSI5Lw47q0qa1
b9iyu+/5itebK1nq91rDaXWc5p56WIZE2YaRg0TupOvG53udQw25QVM5T89D
hyhjTC3rVP/Z5IgNH7tW2114Deymu5Uq4xk7NhzDqgGdyTrjVl8DBSwhmqFj
VfmsTgO7aAE3KFKTNQqhw+uj61rR74M7h06yclgwpMKcSlT8VhoT4dcT40o+
Oyoa4Y/dGvv2ArXWc3P46qHA3WPoULK/S+0RN/GvbmmqMM2002UKkPa4+Rwa
QF/9aVFRdaGx+6nLzk8Wu3w8UOzR3zd3Zb3WSR/d5s+YxNcNt3GiDI5brSAZ
ARZKN/mxMXPHxT7SVNYcuOYzm8tRaZgMcZd60Kz27brosv20ZI5Wt+9UnobG
pYSZSQlPCwJhV1sEKmlylCd3jyi0//8ONY+Gfxs+8I5Q9kDy0ksojQJKHqjJ
Qx+J+ehVJ4s4SA3cpzA/2Fv5UWqCczXr6jcpMAnFvDHoZC7IEiCJ0Aagw5EC
LEItS4pxCEwruVYIbEOfeANowljIIqTDZyhjviYDSTZ8EmijS+3XoESQ0O/o
yLMEiJLzTeMnCvE2yYAFsfi81KhSI0UdLn0wxvCVl1bHA+RWGNAtYPMXMnoE
yU9+YYQohcwYDx34I/AB2eDl86fVe1pQnjdHeBVrxF4jHNiavrSin4KK03vt
pnTBH+VLPzmNT0Aqs4QNAB3BxZ5EQpZfP24vj6c1nH92knyb8RYTCwozXquu
eC+YaEb8DFFmNWFLniLKWtlQYr8hWuphLKJG8EyVdhvVp0xLR4oGm3cXnQAw
NI/el710RI4vJXTcrn6H+tM4Z3LBYajr4djUctJtEKGLd2n5p2eEpjAG3bJZ
ODRC3qEPce4pjWURMMW/ZSYUtIKyE/X0GzqioPq/wyRhhg9mmU5tRRNOVLjR
9ivdjtrk2DHHhPdoNV2lyBQddVpV8mVQuuA8FgEc/G8yJsEkzNbb4Fm4eItk
HnurqjaY1AancMuSWAqxPlhHU2lBT1dWhC3fEpAABcy9tNIhMOqgZdXyxeDk
+JyNcy6nNLubuXQVDRMknbCSR60qi4k1u+Y8k45L3basz7AElqaRufQnnfTo
NhHegmL9cFtfeFRe8iNPkZ4O4E4Ut5/mxyxT2n6jlERWqsuhHCSGm50G2KAu
35ELBezxr8431Aw2X0nnDTQPamGI3HI4TnGlbS3m5IgFVIUsxRqTakCViVo9
F9+jxH4VXLAyfaTrr9zR98B1xLbeF1V/zD63IWbv+EWnDoUZCR14KbZ/PCkD
uqeV47rOYk0GPvqZB7wb9EZDr+ujGQ+3Pw2Ocv6JQAs4fdHvRBLkTmxYUqG7
b7ueirET37SLe59annWIhJSrAkUGjNU9kYqAOHFSsLbtlLMAJjmYBoHiMB6w
+DWROtkWPCMLW34DSZxT/3f3JZNXlZ0Mm8BlXfAdY4GyJH1lLjeIO8wjAjSb
JOfD/GUeH/66M3h70p74DCyWmB2C7ny0Zcq3YQQ7we2GWcgcVnGQTjtFATbA
HZJyyTeanAiYl0e+S4qPHOSyMDj2bHI6K2s7WvxkI43MjXN0HLPd8c0l/5Eq
Odm4AG3uJzuayngOhjbXSOC1OsWoPDvWslxUTZ0bmHSls5IeFV1TQdHZvyrN
7pWy8TIkhEl82ZyNI25Gx+ofLd/9isxmYr5CUUhv6tmWxm0GmbA+zQ5CRIXb
z7ccl50e9ZKjjA2W6J4x4sJe3Imr49PcDK9JSZh8wpaJBhcsijhIC5RvMa02
YApJA9ACRWe2a5zR/63a8cotyHv+x5o+BNipyBCYKCaZi1IUlJQVLSBvTJ0f
6m8NShel41Cr2M9ShG6TzXxngwco2IoLPJ9a+Hphh43hRtgS7q8Dx7re4wg2
65JgaBu7X+WIh2sx+nsgWn26qsg/q2APeWabvElMPgjazEPlb3+BXdXnEa7o
mX8P/78Int2aofimgrTO23rT4I8kODYwP1c6PmEEgY+BM+jj+QoAicO4es7h
oDbSxZd7qUe/nFnd/8jJmZjl0Zbd/mVjho7hr/GXeA8Oz46ivv3OILLO8gUz
rcPIk+M5wDPyAGqY6QHJ6LK/YJEkt42H1QIW0C+W4jpvQhenk7DgiVGJo6lF
z5mvKQtHScPXOtJ5Uk2E1lxAKl2LkZKkeYc5dGFeyHm4LMryEsprvdDtg+iu
GhxOsSF9F2xU/BUjZk60VL5+rGqfNqZo9AB0dq/5k+dw3O9QRy7RILEvF6PO
Iq74nR5//5ISBDsM0MCs2O+vY3yLFqRq8M6na6377NqQHfEqRhFbQgyMH5ap
zFOPwlK/TGZCaruESGTLfnJto4uVO+UNMy8yAPTOKWVH3GCG6oc0CgPsRZ9f
DVk4CxbwAJIQBjdiLsErBJSgNDuGIGFG3R0pB+bctDw5bcJeWk/FttK9f6p2
kRgWD80lwcnsXKtozGexH9PqLemxqXISdr/wgMCMyVdrhDS+tvBjfVpmPf3K
4EpJVC0mNnsydTqOVF/kvwuP3wa1zD1OqUOqo4RKRnZ3QtX0Br1XfJFMFQ+P
GINK4zgaP42JBbG1LyPvH+I/LpXbBiUCLVpfWPo47HYN0tKe/JvefhTwWsk/
rauygp2FuNrGk2S7P6doDk8x7zy6EsY0rzHJkTPXF+27XYJO+CunV2Lbhkgx
vrUNSXgJJCwxFLP4D4DeDfG8RUrk4hTsSagkpltLs+YL1SJMyrzrO/4Ludzx
3klvashJdLtuzHzXt+dSLAQ6QBC5DPeqYIMNDdVJuOHuT4ITjS3lRVt3Z5p0
B2rLo8yB56rm4I2myPrcgPzDjIbhVLsNaDZLi++WBdcCgM9jRk2GANn77bR6
zXM0xSTCRtT1plV1A1qnAVJbfMwbXNdypwFJ8rUvZ56Fl69E06uedAG4Mfp9
Zk4Q4J58LbSzKvXZQT3Y7CrEizDLlS6GLrLHXt7kM/ov2X5V7hhsbI7VRxd3
nRjL+XpvP9xLjDcoWDO7UVyc2SkaCLDV6YJwc4e3W2l5PPgD2uFV8aGccjRE
mlJN8EmymwhXDLb2JOBrYdn3Me56sdnKU1FlntNujDRG87v37kcs/B4KcQFI
riu4WPlsvxN47ds3c59NVEIJXdgy7FITcvqDVmox5L4cfZiVZec39EfWdWzT
+YIC/pwESDFbB7rv0WplTPIl/LoKyjGzO7XZlCODiGT78b6A3yDr4n1AQKVA
70kTA4qxS0+UIbDhJ0wm9owiNpTSH2hbV/rJHgxVNxnGarg2MS8GZxWRb+4V
JP3kLsbBFDrQL/eznuLxxNlgYmvvVpaH75Gn2linYrTrGQrssfzYmNqSQPkj
EF41YXxpqK3bW+pahIgrHpRq1He738AV2axnYGmRabOvGr3Yjr9c6r/QjVVB
NeBFfg4qq2KIVzRFifBXa9K1AaTvY8tLIptcwiUn0MU3kbV600KkDTLJV+li
XJSPZMwQNa2xHqTExI+kJ8nJAIOmo6D1OTagBYcTGh7yY8F1d1jA9T0N0fzj
x5Mm8Rkz5MqSyasGBihZOGMSdUKmXtPA/KSQ9XDbDzZGSEfrErjDUwGPe7gb
1GlX+oNV7l+UuVDRZHbRNhwGAm4yHptNeuPYn3mqFUSupMJ6ishtG8GuAXeh
lTkOactxBT0x3a7wRbcfcGaDFZNaeS6/MIofLiB5dzPxEbr9qq/DiIk80Zac
YrRfdYgdYviXA9JZ6U41RmAF7JUR8WFAJ3ye1RdNsRDo6cwsQpMa+iQFA0oD
BK2uxfQeoqiYPqq5rgP4UG9OLtwpoLpfurdpHm//khxuWpsO/LbHYg9oHaG+
fasA0ZNqY08CqNh4qNc96Ep8xMMTxv2e/JaQ6/8dk1UGc9a6HFwTO2m9n8v2
WQGLJqs6t2O0U6Z6uyndaqCA/Ca1JQtCELQ0A9BWL5gi2WKPpZW+jh5XAJc8
IctrdDOXU4Ny0DWov8qa8JZjW0YEGYJFCyYfOBP2h8IHWmwNEjVtyH5fxvZ+
MPo7aTdtvQQgyvfQc5ebDSqcqJIAGMweJRfhj3zZzUjabcjaDvckH1FJDQ6o
Um1YaoXo3GegRIHzh+JfU15hCLDA1V9NB1Ph9pksLiEAeoBg33vax+oI9/GJ
2V/NuIx8YiJolhQ6k9YL5hxB3E5cAjhljkIQpimxQYiqkkwbGn+2XtnOxD1S
sBF+BoYnKMDREP3Jqf/sORX53kDXe5uEBaDKbEkro074n++ELmhgZwL6JqeA
cr6FY+p+cHq+kyjfW9Vt+bzBSephMcNi7RkX5e9CJ0jsn0Phzev3I3f2+CIq
e7fTJK35VSVPnvqKHcEZqvXrQkSv/Jmw5xDAmL0bchBCskJR0RcR6ao9d9sQ
/VuMMunZ6IHIkUWpGZPPizgpJ+iPUk6osZNqDtMI8NMXeZl0tHI1AWWpD4ju
04IqmQvVBYauFPJR7BtTXQPpIzo8QWqGi7nVqk1L41SdkBSGVus1nfDvS5PL
skmqY3ZSsVO8MX8ylZfPJn1Vw0iuHHDJtYxIO2NK0rzRb6yql4xMI9YlR0Mm
/I1t10VALSMeFyVNw9U7VGijq33+FuLsGtNM2LS8vdKhX5Ui9d7fCgkUFYc9
2xplh1XMqKKmlW0H1RD1I77lMYOlqPpPD2kfPqoDdHkehBNhA7bv2L1TzSY0
ofcaD+X6IdaCKtjfBpAlX/srJN/C1WDNmAU8Ot66xSgVqLgOOoc3xMnNV+a2
UH9iwpN6S0DnyBO/wQu0n/cyCjk0ijV0p3bXLx1urFbo39HzOTbbUUiPJ7DJ
3oQMgJSW/L0s4HmEF0cxO3pDWhk1SggNcEIX1F+iKAl241qr/7JnFm64lqNP
hC9WepdarqtV/brsOol6ayY2lsyqu3tcao3SOHxzbdQzxr3OMXpWVbXmsW3l
ZygNjyhxgmuLX09gdQ4Q2kft6B5ZO6bTzLBL3f/UcVVTUshnL635fuG5tPY9
KLzFhO08/kEK4rfrPRPdQ6676Af6kmYvW1HWTfXg26yO1TgdMFMTo11xvHrm
E+ec0zMNw3avBB0upMhkjAchOmuA8uD7wiuVVtUurbAhoRFn9Og6eq48Gpse
GyhUjAWL8N1EQHz0qri9GxH7ib9NB0G3/oMoag/PpnKp0C2PY6arlT6otdTI
DXrYJIz2F97kJ4LfOLxK+jPg9IakoVUUFu1WqgCySKaplxReUjfYIGuhgeKG
8YXPQWHE4u9fAeUkEyJKJJ94FUxNx1lGVDN2sFKOFGtQkoz6wt2epofp1VYX
EIaBKbJGDjernlsdXyQF1h7lBRZ2AgEyPSAZgIAr/fujH/k652OcpnULnly/
dK2/z1lovGM7/34QUALNbRdRQE9hNPFI3Y4kF01s0CuUoDHATSxjzblXQQyz
4TljD+yCNA0DJ80I1UTz05M0OkdPTxry1jNqfcFB9BkL9RpWLXKtIK1yzUat
ljF2xZuJahXJ5iMdvtjC1Yra3BbfG0tBqEXjT9lKCoIEAGuUdqNuvmvWO5Tn
+ZAI7eyGaRtEXv+tef72LkVe56Rx4dIsC7xTC4JGqVIBe+mOw+eMuUuZdwBh
xVPJfRqK42xvFP3YqycldA6yrgCVcCQ+VrBg+TCa9CSiVfXjaHrWqZ+gYQwY
w9ejQhn0s8vuxHXF9yVi2WOAJN8KDzVIaTyAqtUEaboJE7a3QoRVjiOO6j0e
z7FXSLDGZ19aZ47jygjoLPNOIzKTlGOlHhZ60nCxwrFp2I7oLC4w+6R/B8+Z
nHqQgA0XsQt5FoGkljyWtSAxFZ0N07TYFJbOAkCb1GZHpAZmcc2R67zUnyjo
zP81ytsDMBa8vULyxQOe0mvv9uBpjAcjr9M9rRXJb82PDXCFLdu7rPCCJcC6
QzvdMIiSfs+Nw0ehXTDKtXVfzEJyclevU/AGMGxDj+HUuxBNL4dyYUXJJJj7
WHaD1tpMM8hdUShP0XMaxLzlPX93EkXqqRsrZKM2VkM6O2uDQbc/J07ZeDOB
iS6cKCnBjza6Kb78Tg97O7CgAHKRu835ggVCZFgKLQwf7+gAGBHSHdv3x5T7
Xr3PLtUhtrJqZxHCK2ZrAqxVXkqxuzFKrOdH5JmJFM8zT9PhGfznARAwR1Kb
0+qCS0s/tp+yYvUStYf+pU3AIyO913X04/RaaQRFuouAPQChnnPz5T7FKmce
KYBSKoeie52zk1KQj9QXDFhIZBDZ3/pDQMGuFUlbt8sLoOiIpL7IXtH8Qgx6
Z4PeTrV1CDb7FLtJa6KKJeN0JJE8pl3yF8Xe8QUY9ioVqEF0ohoSm7V/QNow
Hgybv+0JOy87R141mBnZPCYr9EvWb8aJRm78JpdAfdQuyHR4SSI0yAVmiRsb
veQc68Pbx0DMrYQss9s43rLpBJzwB1fksHvo7exdEKArm2T4f5upCfKKzF33
m3H4+pZNHe19HYTAq2ojwwf3NUixJ8ytidFwEUoueXaJnCIucVwA+6KViI/4
oqbq0m1W8fNmlB9BudRz1cWwNRfzYI5hvKMq01oVkIQ4kWiWuR/1WY/knnQ+
bI69KOTGRwXo7J/HbgOgsCpQsoG58yuIOyxdSt3dvA2/FcL9zGzWehClrbrT
+/aNxisAiNg1mzx1ZWdqSff3oNgnjz5GOTv1HdEEG7mfQhwN2AYDdDa7aYZ9
m8MuGHdQxkhM28ionbnT75PKuqNmQJ9ZbXxXpu1PpazUqLRMCVHptOdRfvXm
mEkVx4C3N6Ta+ZowmCrSmcwQ7fqF0U4gNLJTby0X03CYKmyaJZ/UQ6FZo5J4
p1kOQQwajKamtuQyArzFbmhr2ArkC7xYC699B8zhEIh8++52LjQeCm++KQzI
yy30gYBdhAtALiiKhgK27f2dTMVkbIdkbV3Al52Im4l/VCnoYcUINqYTU+uE
q72VOetQLGcMFC25n/NeY4sJsIVGf/cHfq6b43aBM1z/TxULqp9FvtOK52+S
H211z+yqI5ThUbosD7PfBGY4QPg3EHl2DoSHViyJiS3UodRbL1A6ouSgDk0t
OTs3a4AhJLtJmuVMAWL7EUU5RtJqdH1ztANSlsFYYcd3Yg03UYEmRyC0e5E0
sR0MhKEwwM0VTUs4qP1EJWShb0gmwooGifn5kWvZJedAODS37vN0eeaEJPjz
RDXLA5dlrF3Khb6tA8CEEnHYHVZ77Lpl9HRBNQssvZXnOwRI/T6bONYySekf
U5+vQZkw6Otnzlp7EFbYVjVzAaimCWpQfUT2cZe9Izto7a/esnEggNr8oyGG
TlGXjur0zpAFmrDsc2gCnlguEnrvk1TP1LmgWImOwBRNH+Xm27uPJpkBuIZw
YzDdmhexMq9yFrCd5h87zgykB+nKcOwG0BVAyHyaNNZ7N8RJMf0RNcIRM5Yu
UbrSsT+fEzDWS+LODlUyfZwEIT3KCZjxqOqPM2zwejg1suYxDOSaAiWV3rVg
NuNPK/hcQ7hBbcnuUVkqAU9HuZFcSABKAtj+NfBqYWCH/ssEdeO4VWoBfbMR
rjkAQ25/Hrjx6Ae8f3Fdw340K8Ka4hfQCOF1DEvYGNubJy00lbp/lk5VWM+8
kf36kKLlIkbCrSfi+UnokCwDNImGNMVD3LHSjUaIlmHihjGaxkugsoYtqUyi
kU0AIwNGznisoPTCsRvzqySVDQ2cViVoMPlO/Cx0/p4QzszSMIjOVEI1ZfDC
7+rlD9RYrAt+7zjsXcmt64/Aagr78Rmk9EzFOcUK5uDBmUKzTtNMxW2crpM0
bI+HueMc/SCL52z2HMyaA8Zc0OJWkkPUQn1rC07vapsOP03fI0Y0dzXr2yI6
KaTcHMTcamtzaJ2J27i5v6yoZRwsOgtGJPjI54CMdx/PpzSkTC9DGR9/9HYG
N2XHnL71EMGRbjfscLMf/ogCKR/+qqiqGATQmoPV58dZoi+0Zze/Lh/mej4a
WcWGKYrP/taKQA/gKMjZygMm4jaYhl9n36Az6DZAKBJZlIy9JYMTAMhPrIyJ
XgljHleSe44fW2M59hCqKD10vt7NUaQqCxIvJjZMgktO2rm0C68KR82D0RIw
jkyVQZlIZcMS7EVQOa3dn3ipv320ebqPxzpeHMXObwXDSoD33w+nklTlLVpj
eK0jsTpvhs4APv6E1vKs+yV+7zFsybjG247AesODsgA2y8PtjAiO1usAufll
mc0LuAJA+5B5MUNZ8o67r0HxQdSkGb5/hbyt+LElPwrqkP912I2YF9uiunjw
S0b1Nc4Dkih4iNp4pge/w+y1Iw5iBSKZW89OmcnFf7giAJSc7FkIRup1nMg/
9IGjak/NZ6ycx1J9I3SAKLSLSl/SL8QwwY5uTbY73ZemOX5HfUQ74Jk/BvAl
2HZbFapAwg/DzRh+1clYXm43TMRfz9QqucTbyhz/1N8+D+mKp62mw5yP7KzE
K13O4FWlKeEmx/bzdwmwozDWpQsyNLrYlIWgkbBH74Xq40CCjMC9AtLL5i3W
+BY2KQiQxo1iBQWudONdf2+YUhSU2S6jwPAQ1icUjK94d0jKiXysHsqIZWGz
BZcbTmn62TM8l99m9e0TW2j8NhsQs8BcKbwFSsFpwdoYTr8LwzUC15XtJdwk
rzMdL98FzwC92XDN0uJe7WyA8MmhNw3gb/GgWkrSnBsuvuyfNPijOkiv0Yxp
GUmUuZZZCd2v5hr5QdVcv+yfVU++4ooRwocQa3Uwb6gM8TIMiSQYRRKSLSn+
+aZD/VjFr3gH7OjPlrRmhwW1AV2CZyNbzaOtor30FQavyEk8kqTWyjCsIOcz
7hcOjUCB0izvwJktvkj9c2jTQXMCmfXMehwprqm1R7h/iZiT3P0FkjKGsqTM
2bHGmoiDHUWJ08y3ccPF9xhCSQgYquWZLvOD3bRv2HZ8/MafIwHdkPqV58OW
Ed1RK7tQzCLDaCEGr0hGRO/tIOzzvKpmfafa3MY+axUqaFHAqXAtI1xn2mJz
Bf8NRefoxjhgJOIYSmskFJ5jsuJBQ6wMUoovfYAXHV+Ihc9XyFclagByEVtW
J4hufSN//788+zoLBBa1qnPHV5JMdnDEmTQqGQvzds5ovZ+kzRP34QYiOh3q
B+Ws5SyiYIYvF768PhclXKBulbg1rWNeLb8tir42yHQdS9Pqp2D4oUnlc5e9
dfFSMPDj2P4RT2w99JmsQyv+YtZMAJkT7QFz1w8dKKc7A8dnlJeTXWzE52+o
yFKblfodNGFb+MMVMIqbRLxP7mw09SYcCyTJPzqi2YVaNQhwCTi41KxHKf9R
SCn28bTX77Cvo1Jlh/iKlcsK/8qwvixQ6xdAPUQ8c8X6SA/cif0hWCBYbVAO
McV3gNlyzTH/W5cSuOG7V9jKktZWtVrhEIh5hlh8WpM/q5uCsb3Aiior/1+y
/WQxqq19VHhTEm7Y0XpYc+blObgLw8ETSXqqwBIk9CJphFJ36PltfrpLlNZj
5/2BE0/qyoK07KemtfgD1TdHu3iLlOYRdkTASNVH79NVYwjg9tByu6oBV0DI
MqzSNQ1pjZTF/djSxAjMuabYEPLMZrkGlLwgTZX8wNAbwV2Y0vBIDmaLOxmP
rud5SBVdW/atAsWCrfPx0+kBE40sYZ9PrUC8n3Akfbzw6YFe2MYPB0TAH9WL
lmOUtsQ0d8Sc1BWpk40+F/SM4HItYsHemaAjzxH7ZxJgV6Xk1Ky8X5a63I9c
mMGFvCT9swf+N+kIXWdOZW353OpsaJmzxK0TP6CI7ZbJt3hAvPONiMpt5Llg
en/al7JW5ZCQO77Gh5y/c+AKmrc9kFl5ysNr123tNMnA767/BqTu29jEaMfB
ZWBpVKbK9EbYp1b9YyL+7x0SexEArYHUe2OofYgmW0rYw0Dgt968hKTAEoik
oTMwb5FQ3ZLG4Zt0xIRN5xCazz/2Wst8A2dHluCDz3Tpya84ZP1tzVCwDtVW
hFQv1sMoPTbrbMGSCp8iVglUIcLbNyU/FZlc5qBwrOFi9Ooo1ivRMY/h9I8c
eNijlXLgpJnIg2LqeQXEcgiwBwE6BboQb32gMRy67W4NguBvPLJQ+vPJqdnY
1DMOkw/CUCWuXQe1da2RsUO8GSL3zw0fNEbyIpVQZCWOKi+65FeSrOVz5PQn
f4khRcwVRupswJZ1DZcOhkNOfCiSwRB8TdnVAXCmz09D3sk0RgxJVl+CGbU2
PH3ku9p2+IxvZFrBV0hHIFbv4vIsyCDyCWa+X7p3ckA2W71S3/hA/vZnVVds
lhTSO86l1a9+sOZ+7OaN3UKChmTnocVmtAxLqkZ+nmVYS9bMxMN62OWBAW+P
dYwyRxhBX2f066+qY10CCMbV+u6volgVXo7KvE+daXWaKadSq7o2f6zhEKKz
Xc2xJLCoqjyUtjbUhi50FOFoxAxUo8sofCgITFRQ2dSDYl50zSJf8KRxbxzs
s8hWboxM4nIB8poEEiF+pVgr/o35QUi9Z0+VTjTdHtyA91FVWq1pLsDvgnrl
60DRZJwIfk9nWg4n0aAJAMruhOly6ILFuqof49BncxCE2WgKfwIimtlBY9oq
0V5PzkcXGbwB4YhneZ+oFS0eVZPU0DAFmR0+np0PqJz3Acr8hiBYFyV/tfFX
NZpO5LdlU7Rt4VrBl0aOwNSKX+QOZTUcwVonttthyhzZD/6JNGxCmdH51M7c
ldBBqwUgi+FMNjSi42rYGE0BuXXzK3oCTTtsQ7QsJURblGtrh6heXTxoXBVL
fx42iGzmO+pr+Rf8l/pjcFX6ypKoXviH5LrcJS0htphSLS2QJ6gLk6I2e2Yc
JQnc4xAnT6limThXowrkLJ5GQfftGlTcSjOeQFe+x+0VW4jqbqZYgqeoN4/n
GnAWUANpLix3ubve/q+WOk/bBC2jTpdHaU8pSBFGkuDJQbRz5yPt0NejuKw8
Pt0vkfNwn3SKzLTDg0eCY+BD7V1O9GPKvpfyy8gtIoX+3Kie+GM/eNHVQy/r
bmSGny50qO83bIJjwbtc1r/s8Ag6VAX+t/H+uE7qTCl4Jnt8oSN6VMWYGsaw
EFjJRlQSJvPdJVeRSrYAA2KIHfaz0XZQSia1tuHw7vJCW4Wc6m32TzWjClBD
XeBLI4sQ5/J5j385HmYGJ7laqDE5NrKKEOtOThLhdofZmBLdCoS4RswrQR7f
y+Xh0qAyKoFBIfNEFs6yN919cToKHVKBZQAjjSbgUwuRI/dTCtEtCXpU4sxf
zJhR3MSmF7nE/tGIWbW2zsJ/qglbEaPl69uYZN/BRaYaWVNqNx4oBTdHy+z1
fq0+/mMUKO+hkrRYEl87In/A5QAwQeJGbwwNnSQBoJjaCkaRG7jB0YcEus5E
D30N380ZS0XkvRNLqqyrtekbllU7npZA9RdLqNX3Vg63gJMNJpAJ0Dy1Ff42
J+75n5hrx1mit9TauOhtZ0n9U5oCsQh1jSRBo/gQvcqF4yoeOkx84TxkRRw6
9hZvADsojAC0R8xDH5PtKwqXYEu8hLye50rosj9VMGhIV5cmMPYoJOArMKpq
D7smC0Qvh6aOZXD2L9NiAIzvvf+aE2+N07V8qmSco7D25al7fWKk5JNMgY6W
ieObR8kLS3POAhK37O3w8KBZuzR52AzE1FNO7jyul2a9g4v6SeC9efxF3umu
KqInw642FDDz+1MDwLcYCosjr42nhJUZ3VeoKUZaQx+co9efZW0tVd4zx1QA
0lRk2HhHDbKWxva1fpCvGSA8qKm03eqNWxqSEv9tCxu3yD5hbU+P54V1elg0
QNNFIYV5BDr89UXLd24R6o28kOpWspHi5rf1uMOMK+tDxEu1Xft0XzKE6a+I
Oc9IwK9iGvaKF3UJy6DU62tqlFNWNLIwjkN9L61QotemqwVPVRPalOsVWidV
ZNq9ZGQfocZz4FYPwsfatQGmNHhR1ci9ppJfR+Q6IaVMbW4SFcbPEGSBh1CS
2N6Po2tiTTdYQVAOsqoEgQe1CjusmesakGK/EiVcQLGqraofQbkY4I11nUYf
rsCZGdGzJlJWt2AZ2FaZwvos+1m+0419f9y8vnAx89v+Yyfx7ISdgpqYXmtr
nkvwx2H0NyOz7Qa2/1/RPBvj6COgd5BTmNauyM8uQikIwDh18gVhlrcwbmxi
xYJcx7OrfZxSca+xitnF1Q7K/32klpsyYug5aBpzMftjPJOcXfUxEpvvEpvj
HPXPQ5WSHsYDow7Moc0a8jmq3IReE5PiEeW+bLYLphwsq0g7EMD2Vx3Q1I3i
yzHEpCFw/v94D/rJJ0QeTtzrkiBbQ7ko9ZCSCR/YmcdRDKO4Df9z5vTa/002
h7MaPof+xdp65KRrzlFfnPMDO/4ABVhZ6iRcswXc6I7USnwZ87O9Jf5lgOnL
GjVLeygHhB22iwMP7h9P84ASmr1lrVEpNpX3JGM/xVK4CHXeisoyh9MoCeTD
htDC3MvYFKlXBT1LQogmSo5GYrB2RjpHvOcLoM/MA66+s/JQT7ehpBrcV93q
Wqxz5vBHaSIJ4CJ8/iyVknu2OJq+gLax4NIlHQa0TKxDrfDW4TccWlUsN9XU
AjOniPhdL1tiSPzjoKgm9Hnb9Al/kgcwE06k9WFKBUhpwG4ajOZy4iFxRYAm
oaIp8BO73oawbCMe8XBzjElgaDA1Hhk54P5dnAngkHNNDHywNfdK8zDkDA3a
GpAvnAlj8nrnjB3ACcuOaTOTwVAHasPZ8kf2frUbHgPPc6cRcjSH+FSN5NVV
Ig28r0SyJsD0nsUa5qKnZYDe4ZHnSI9ZL/s7TUtKt1ktfKrJhUtxvmkgGp0x
VCbZx3I0CLSmsEWPGkkEuLv2uA7hcFyqFiWaHLyx0/D1Hs3w8kC5KK/1az/p
AywnpihpR2JThvKY1WQnHO1pmVP4fy4/WZmIVJMmE2EYixTPawTzYHrMHCko
8F8e3SFZjFf7PKf1Gib8eHsN+VA9tFk0v9MmexIHXzARCS0NUoRVpLhwG3Vf
tzCniRFRuqk1G5llM6hWgvsYXcbSGNHrgo1yJpSM6QHH2h1wALLo6c0cMIFz
/s+/2DB4U6p+bU/5OB4fnfnWxn9GXjGUAC9llmaxewSjf2odD2EItU+GLgP6
bbz3oA6UNTuvBctKtyRVvoVzhrhcWL4Icus/2wRvsOpUG1/OHk7lRWOf7gj2
s8D9o8tbDeJg1n3dt+ibimsU3AYwa0WrWdqo2oBhhAEFOJDRnPIK/pLe3qfc
B/3hIhGsAALcaZ0q+MX5o8Xna8xTqquCyB20g+RMscy5FYVs26w16rN7JfUR
6rVSzlK30RRYR+sEubQuU9DbezlwDqIbHH2KVgmfzOJBaI73PGqu7MMo8iLx
jXXVrBDVBWXgwVRjw0PUYupOb10ZAV4T2GjOGa5b8jx9WhOhBH5B3kl2J9D1
xt5Er4+VxuozhM+EzFTYOe5sIqpel+zD4iUngHMCb4kDX+m3A6Ly/W4M2LMq
SyP6NaP1gundx/LJuYV/v+gE5fj+qPpzlNA7tX+A4lEeHmBpUt2nE/cah7Sg
VmBlDs7nlJzXsbfbX0VJ3p2T13y4IKmYUUQ5B5j2Pze8oZyo1jetZFOr0zCU
N0IUaSOeYqqxem8B1lCVtIEiZTtb1Kf/OV3vtpxZqsaofFzFIn/dcIV9bmfx
qdJLuXThPsf9ClOirLf7uUJh3fS72E6E9SOjVDS+uffqgIJxFs9US+PqN2L+
RBXfwyYlRNgm5oJ12mklzJ8O71tIrFDcKmikXIjMP3y6o4Hy6ppFBZJJ7dXn
oJfrcWkyndTALnOYXnKFY73ai55s4X4/tzQzxSkZQmE6XjZYYHCeWLRlPdDl
SRhItwAhYFJRt5sywoQTpCxObf338Gw2ZhO4Z2u62jYobMz6PVBucgm8w4en
ONPIjagPzPqzOyTJ0Qg3StCANxGyv+9dXwx02u+c38xUUhV7Gmxh/5y+aYLi
Ux21GmNYmS9+QLpHdTlV9WEdY4V1WAwr5jBI1TqMbfkY5rAxx7N7NXB0Smk7
/VcpXG7dF5mTSo1LN98NlzwVLvqyQoQjesdkBnGQDBDxfEGLVJiA6BZWklXS
8qjQijCA0Rt55IKMwH9mJjY+VFINWiGGxMMgcVWDIPZHFoT3CWnbPqYZXvVS
Mb6PqHECYK+VnnprLUWvLKFgrpMqyC16T3FZ4LOGLLXvK0vTK2N3UDfN26EQ
Td45oQlbS141Z/jlESZyk0iIxdHzHIQPUGj0qzDFuN1q34IDQitK0pLIgFLc
CZOPAvg/DBMz+2cq+X2dK6Y4fvBO82oraqsqLt3onJQp4Nhzc9ViFbYDKBzK
pQ0nqJ13liK8+tEck+QJ5FfBqqd88xYnZ1/8RMToHI+CSkOsTSGQZTyVJk5U
VOZMmOwbPtKuXBQWQ2bcbLNWWRDd5byuFENCmF/QKM//wNv3v0d/mO3JKS1M
MLd6jm0DXLzsC0aSGURi3pY7ZXPTVZkYOVoo+edjpCwm0l+bo7YRdiwiiyWO
t+47Snxp0hSAWhQsTEyX8bWHAzseUyuyseTWXrlAIySLVDayjgVg46+0TK0z
eAauC+4M/c+1uwLd64Oxp5APr7UdfB0sPbREoZbdLxvg0znMJrjWi+6ppw3/
fMBXSbNjfvruq7sMWA9C0WMmiauSwceSfchJsdSbAjIBtB6LEesi0Nz+KgIK
t0LNsNjoZA/R2Igi53DgzRz1wlM1JXz0GVh3M09nooNk31B/Ba+FRB8Sd7Yw
83iEmXzIfDlhAfC247CMRBFs69v+Pw+L/yBXJLuQaNg5kmCGonjyu1MxviMN
rBy/7/q5t6zLzRnaxpXRy0mRFzWyi4csBdLl53Q8Am3/D/J5hcU9ZalebFhz
cdjuEolQu7Jhk+z0HbPgMCRHRqC/iqrHUDIHzUdXut5uA4Yz0xyHonNeu1N6
Q1yf6wHIeGadfiY5o51bkCTciQwnikJdvS8VDmYivLcqXgeJjsGca6bP3Lhq
SA/j7kF6Q8SVn2PU7qLBP59klBHmzyDluCesQQuOHKtL/TbQX706wY2XcUSL
y0tiiqkk4/gD2C8kBGHJPaFQmbzdG5o+Sjmbs+BUeZycP7xyFLGntesjDJXo
jQoIwaZIMRXMQ6WAnNzDPLYd8GmK2lntH5uZyznowSY/UX6hoa9GtYyVOGQd
tmpclAMn6tH6wxQrh6+HA4vW0stuhmNfTsJ9CD6FLwI41oE8o/k83ULpWkSM
a9Sa17vf+C/jN9fKCRwOisXPBBgzMFEQNCrsQ5O36DB5wqgZbb00zOat8+lu
CCdu53oPnecAEhRAGtoFWB6l1MFVx4thcOceEDR/G0c6iU0J/wJNgdJ06LKc
ngu0ltzeZbJcDh3a9EJ244XkiiLxvRmOKHvr3tlUUuEccT+gmqOGlDLSwMx/
nXGkB7l/DB0qK9v5jhny8yBoj4VgityvRyT9YB3GCcIIOY6vuOmnYlpLRrtI
qemzPxqIKoV6p1W4GTv1FF2KtjFUZEUx1QnogQfdZhTAcUvqhJZgq/FGM9W4
fldG91imh8dia1j0owRzb8/3UQcqk6qwh6ukUXlAboZ9SenSONRdTHpkz+HS
UE3CTvF68OXkjiytfQAeSa7Tr1qATXsOEWI6AiA6hv0LICiIK5OVc/Ozkb29
YVM8UNCVOWLP5NVk1t7Ei+nlFf7dJua0Frk59Pi8536GEkxXoAbzwyXMetkw
PiQbhj+X4na2Y03Rtap9xloBnFZEPrUT3rhvj9uAryopJ9PY4xy648ryyXQF
GJTpNl7AIzQnI7SBoPmAcfUsiGHOIJrwdzoaeqphBLSneP+W4AjN6jWiSdPv
UskC5SqdqWCZEAv7YSD5/aEBIhl1GOX75rS71ncO+niAMJNWXp8mKvFuYO3B
31fK3DUl2Oa0sIp6KQlC3tL9yxfP6WCRiH8hye3oEdtbtoNQ3JK8xFswZtoJ
ucQMA00m1PTR3zAEdzxXPr0iTbEnq9h9q9ZeeTufdEuzvywk38A8pXuXpOkz
Lp6GARa0U0G1LR16GPfrDTRl9dg249S5oV4aJAdQfop7pb9ru2N2rzF+v29p
iPJHZoO9G98nQoAKi7KYfxqU7ZLpdkQq3xecJqOsghEnwO8vZ+gGGkOKJIdH
RClpXVDchzgaSTmPB+Rp/DRlyEPh0HE2pPAvjXJncjFtLRpeoE6mZrS7yNnB
ImSOn7vCWxSHp9ISPeaZ3j6V6PeKWpT3oNP2CfgFkAQltuIHbdmxfjdA41pH
D+qsHUKLduTfO9tJo4n7Sl5i4OkJu67Do4lGXRkGxYRVXtBCWrpBpi2rBvWN
XxecdoO6rAccJ6pHXfBlZFrpwDz0gnxauHMUmsCESKPRU8YwH/XVHOSvjPcE
pl1RmBlWI142naJ5c/6z8m8sqJ49cULxiGRfGbcupSbB0ERkTtfoQGCM/FtE
YbQu2bTXQ08KX3tpDpPgaChd3JvGWNDCHkq/u8+fsHBwHPVBoSMYAyrs+Aln
r+5/EOqLN0KsIFQs13mUp83XnEPfpiiLw5Vxesz552uzzX/z8Llxtf60Fsut
0R8Ihwe1dTqezFaLgC2f256X7VQIjkSZjJOvPj2HSHBDcVeIw5GquE8JPs97
PKTeik4YHQumCnbXnQ3qvbCsNlUK5ZyF1/EuKOZyIKlI0Dlj/Yk4/V7Z7Lnm
VfNK4xavw38DqyoTrYORgP881ymVSuiROSefKvf7v5BCttuOZFCnrXTBZD6z
N77vdJbNXzDXAt3ZB08KgqA4d0ehTFql2aScQLeCA5nE/prhBUWKvAB6FN/R
GcjpvRiMHSYCijm/VQEVlh15iQmnGsYRKVVpmlaA/x6QzBUlB1BLedzL4It+
Ja4o6zjhQu4ythiUr+5Ls5NKV9XrhX4ba+CkfWZ3Q/ou+3evFJ1ztT6gKO6g
jeTC+7CyPunf36WsldBM8VmdY2Cq2VF0UXChXa1sZhqIM3AMIE9qZzSxWShF
FPJBF7CEJLk+x1JiQZ1klHdXHS0J0pveK441++4sWUKAUElgKVcfusnENBer
PZYoOOJd12ASH/ZFw0KI5TXX6lBKiEve+gM/r6+XW0MRlklEJCrwHit/jnOv
WuAw0rY38Jflgn+kLXOu6TcC5Gk8t3Z3taBUoamI8HUGmFZrrh+hGTHSaRlO
yY+a3l5702fZy9YG7UN8/mUn5FjmBDi4rT1vdvTp3Rr8iGFiGow3TwhAOcDe
RSuW5OIXp1CdIb7ouWUmL//m5UAN8KUNq2px6EbmPzSTjSHQjUZl1KVctQhp
/iWD9aFKa6huIz+4ZCydq13BJdGW/C2jk36g1SSYhhfG5CRtNpb/91iqyC3V
QcTiLKn/UNXOrR2UD3ptQSkKDVkQYFNpxu0v3gxFxkrrSWLGsU8nFxGYVt+I
AYDtPXevfI+sZYnaZu0UEkwBnpo31se7xIkExdeQeLir+ZSZGKN1fqPhOzEl
WQ6lt91VpQDJpJzKOeqApgV21l4zhEaGse4TgxUfMKM6Qe6VD+2Ii4pQKOq2
5Jndl2yiQ7ptalKUIhOvfAQ9M8F0GKujYf2hoId6zvvvYSqSrLUYq7bh4QqW
ciM23HxadsQF5K0PEKh/QdUEfb3SbStuW8y+uTv/7PrIGTnrNTFGDFtNfXTi
MmAnCkWIXm21+XQcFzwBHSLHfpeHhDoeKYura4KvX8Zr7T+WYeIko7xt/Sqy
i5guuLuRLAL7zzy5NFZy7fB8XOjcVSY8xW8ZEEV6rCvAdBpmry+jCAGtgyWu
deQ/VHXXGwqmsTVpwioHYoIdA91a4aXmfzHy/HF4XybS8mTs9GkDhWzYZqfj
7vDOgWaFOs2lkskro6WWLSP39AumDbZP92MqEkcHK/WqpMGthkmJ7K6q+Fgz
cJbjFxCv3kr94kJSa1eOxjVBzOQf5n1c62OxB1u9Kwj0Y+chVQP1Co2l0JvB
/GUnN1waifV9VmwwMvRHFeIDEWxFs3WzZrQ8fga8lsmamchLJaFBU/se5dvQ
TlotAwr/6X4KZOx04Gv+DGduNws6JaUhTr9/TJV81/xNOkbF+NCcPsKYC5MZ
PFZ418Z2Ey34YUl9vdZHpCFQuRWN71xgIBJDNfcHe8C6eEYswHNz4kq/YBuY
8YlP0m0p8x7FHRBrP1ubDs2SDicoDFeqoMaAD4Iqrr0M0CgWfJwXZMp2Ey+O
7uDAV645BpKeVXvgpTi+/9iVGe3cs+rOYWCT2KxkBRDk9sulJqdyNiPKK/NC
7lNkSWIGGBPDw2MQg3hX4YWrxt/SesPH1410fmArimJ2/9ubJYoD4Nq/apxX
IDDja3l+OPkk2nF8bzEuqdShJfE59tMnKm18EnAWgnkeSrsBnJvHLQkvLiZ1
tATxLCDxgt2CNupYIAUE4lJ9j72VCg22XanqYX/seP+QmRnibKG8VcHkEWd0
NOoeEQXK1wofYfxhGE7YT269q+FX5HKLSXVD4jOUzL3xfwDzTzyq9azkcZhT
M6eztOLINKorF/fosgbyBsGZPWOoG8XDiKl2oShDlcxWHFvGbE9Kpf881wsj
rwMWR3ajCZWZ3pdabjH0Jt+ddXpIw48fe88LoGlLC1J122j45s+AB14vN1+C
CfWZp72Qr1FlFZjagBsNsD08u8FFYIncqWKqAaJgbeNImXx7Sf7NxYMFQTV1
Ig7uamXvhHAVdilIemASY+gvCkVO3iNTUbNDX+ZKuje4xbmv5La2Ce1rW+pw
7eGDANLcNjvomhJoJZ0ibrfyBXbcYrihC4KZIUbp8nsGz2YmjbNZvxje90ND
DHVxrFPr+oCX4tNMgPP1uOOqMCWY8y0rDWffzGZse69hAlJSbd6gaiBwOS2Y
iOImEPvREWnQ144RhFbWuNFWTiMRVqg/YkwZWHjLvSIRbASyDUFK29BIaabG
bX2375vOxNljqQm12NCLF3CqCWebK/EfxbP0q8/5yOp6sHMfncrn8LWkeVmh
WgVvdK9967ajZz3YKp7Xm+qCIrcICB4fK1Mtnz3yfWH/CvoCmAAK9J+DIGDT
1efwbrIoZKh2V1zwmDaA28UoiCaPGC9evm11VQdIoFkynycmAPIB+e13gVva
rkpiT/DbyfteH6tj53icc3GDJNYzoqshxwNKW7649jC16l8Tubq60Qy0usMs
jyL+zNNI75RQlxCpp8bw9OGrV/XAVE0bSNYGWsVZc2/1PtYr4Um/oHE+g0mR
RJyqDTt5DmNVdbLCbhgP0lIxrOKMEkYWXdUtHNIPEzGgXC0x1XpkVQHRo7gn
/Awjbt5KI8EAHrkBeIsFUl2a6W+x6uRBK0TaW5OIfqWcajVCcejeSTVlf84u
4q8GHEj8hRT20KufmZdfMypvfejYoAxZ99Fixv9gj5HGXOoJL/gt8j933m0G
yYAvRJ7x8/kQQdsE3+OsqfKWiG0iG4eukEs8zSa2Lcm916l+5ba0p+CZKek6
BduLr702Fuc9vewN5og/b0m2CUjwSYphvatp2eJX+QfFIGBg0T1KylX7MYAN
JwWjWGoRYujkPveCA7rnRZLKS/4JMGJn2N2q3tPXzl+0DIansCKX4SQ+fdQJ
A1gQckHLTmApRPyk5TsOd4eFDOFd32kOiHTqBWnLbkAxKBO+bcHmDk4Vk356
lAv2t9bJ5zuYBPYmmXS2ABb7O0bJX/L/usKq5sLae0iomO422UZ+roeqq5uM
KcDlP6YwopSLgS/E1JNnZCTG1l7jXDbawm50/rUrX9VLoW8dlmNaO6V4FvDq
yoVBUdMv1HxpyXFdzOJ18Vx1SqC885hr73Y9NOon/VnDUZ9VZyLsX/zAz25P
yRf/AFG50oeiN3j2VlVjrLgZHjLlUUE/Ubvh1XLwmLyq76BjqcRm2KRry+nA
CPwZU7K7p7xltuneTg8omnQzYFsJ1cJRB+wFxV3Fs+P5m+N5yeZzxo3+BeUE
ZgDA7lBlyhL3hAPNKHZKWhy3NlnKtuop0rBrj4lGDzBAzP5uFjx2IC7UwJ6n
5p4PX7CzvBxOtSakNqLy7P6sxmW9DPc51rgzsDlp/9QwGhgOW9orgWh2lTJr
ohmajcV1YpoK7x+/hWESPY9XMgfblO7B1rdyNvTY/bAZKvjioBY7gCwfZFCd
MnCIEx8ERdN9DLnEy8RU1FUAEEgHmuWgQrfeLZqBM7vw6vHfgnlMk6ZM13gr
/Nb6gDpCW8c0094E8KJ7LYcNo8ZpdJhqSCGhtcg5o1HgvyLodyGlQk6xxzcw
talR8pYi1lzjpTEE66fF0NV1ytoy9Lv3KPMlYlFEBtMQZqWhDU7jv8iIUURJ
F0BHy2Pxc2B2FfIungpU5pzKkviWAX2H/UzpUBGPDfEXXT6Wpmjari72xtxd
pwxg7GP8yRVkz+KGWE2Jp+fKGGmrkAKy1v3frOuKTEMZJAESUAjnEnX3Vua4
jxbSI5uYvfXIrZOOctsXDYEbM8Wmb1UTeM1WcpfzR+ViHskw7Ii62NsisbnU
cQD7PDqMqYVvKFqIwi+5/kRP+rbRLnYQhq9b3Fegho8fvDYbK8YToAD0PTNV
+Z2yIbEnQTRi8JWFh1hsO1iAkwMl3xE5UfWGBZOBsZRu276r8oZ+E7dx80Uh
QEcdaNK2tKNT/Xa8BOnikpjfskk0+GbXdCBHiu62+18yeby0H7Qv1OUCnYiU
jI/ureNdtT6dRQDowKbSfBxHcfT65dhO1rRhkCuu5GFs7oOAr5iHClErxeP0
zR11nmFhwOYoKLx6tPT0+M2sHgKKbfAx0nO9gwi5fosxA/O5KUHDIp69IN8E
SWhy5k331K/X95/tGiiQi7PO2/DckBaKomChdxS6Oz9/53JrJJxN08clC5n/
sQDU9TnhpaSpwjsic542Ss2H9wkMgjTPb1HBROybndF68xz2Dev3+Wns0Lgh
irIrg+wkCDXxWM51ueIBraHiuAAPFdH7qjkLRnoADXqGNxvs9qh1aVCOvhOV
vHReO1HTWiN4bd/ewl+/x2PIduPKioWkmBnSboI9THWWUDJ6SodUsM/OIFqn
6fI3n2qlpLcmSaPnTzjVl7SK51ZkyT5pzXYhlAVHvvF1Uje8A5tn2sb3baat
Z/r8C5DC4nIacfuJyoVo+OeOj7rW3TXjqlTft0cTdD7bEICGchp2jJwVDPXy
8SnNk2S3pdQa7gTEOFSL4Np5cDYb2RTv7q3Tixe+zEntOpMHabbT181Xuw/J
s6pJ0jt39K30VYoeVgsKkspV6BFnAeDQ1PVTRbf04TDcJLmHpWNuUa0rXx1o
H11LfQPmdDvI2+JTIGZApXOixU1nkSP4weHnwofceAO0kYSCSYuvWWKjHp+d
sNETU1xYWLpd2Ekg3Kg//UE8slolEWXiyaHGwhrGbxk/wWzPjVxItkVeS9dk
MbjAv0L+XcADJ6fPFdg0vEDdpBUlxvL2asY9/FSBAk8ps5W+FvAYBWb/XkhI
Xtrr8J5z32gUM16hxQSTqby75u+IIZUAllJ8vjPzf1sYEADPhL93XI9ZwiVF
W3cMX0eDDmhAMEol4KcMAkjI6FIuQcQdx6zBLDHS6n1dEiFl+WMXHh4OnIQH
BLia2g4WMqIuhS1pVUZ0fpGSuNsRr5G7ZZbvlkWNrk0BO3qH64LorMUZQLYN
nW/PiXgaIcyqUN6qU23m38w717pj85fpzzEOWFA7x/2BJzyvR0cyiCaFBFux
F71aF9nGveKym4YWNDUoDOqFOzyzTFX7oa3Vj+CxDANbxgRT+j7ksG5vXzwH
bLFO1i3z+iqjDbzC88Vs1DejJQhzZH0b+10H79p3iwrIKn49w95rH60RwM8i
v8gColvoJ2Bzk0zl+M0GG9Zp7I4vmMP6WFnAD33RekyFj3yckNHTazk2Tmjx
gT4LSXxjx6GEfQmpnOrLpzQWxq7rgaspZOCp36DpfQ7b3fJegJ2zvpfkC6MR
YJqHnAxC5dyJ/e3rx0TYjjxRmtp72/H1SKJf/q+5gco+wps7sOCSe1wlkDbc
/TgSgte5EphqCj8XdUqb091a+gWE2CykTVHLsiEfrMLBsAOnb/9KwJpd+3Ax
xwHR3Jm0K3NAJLPtX1yn6kXKKCaTj0iIWL9c6Z1+IaahqCejN1QMUQszmzbT
7i4KB7blUxlBm1135hD1Iw9LPlOA9GAu0YdvCWq42kY5gMcxlXmv+vlg9put
fsVCoesQE+k/sqhu7zmNNoW1r8JlYx+Vak+fX68aARHUIiMJCy+YEA3tV6lT
/bV+66OVRV6CpGzvZyNbfn1b/lD7s1PvjCZD6YMeE0jEkSKR0OFU44lBpwb9
VyPuzTcetEXPUspCcQJDXcHM6xbaQcZKFK91CNc2JIZRPrOwdsBrry5znuRI
0WUzCOcHjibGObPXqZkhHxNXjAJDMZKvFHjmYWbzOeSaW5znbJsc6mkdlXNy
VtG4xalJWDddqns77iu0ktj/Ti9VzHhkWPO8XYhwHU+QbuGp8IsfOA7rG87I
qKimPlBy61Wa6VsbHBgn7D9wJtFEWj/N6g5ANQaOTz3qc+haGru3eWmfYiRo
R99uJEp717cJypxcmpEleVDKLpkVNQqtcHuPPX58kqr3EzGUkUitThsnpn8N
GMcHhJT8Q+W7rShujfJFMh1iEgR2oj486XjtRwJb7ZioobSe2hdXLMYtqwvv
Mqdk42Vqp9mT+hNpq5BljFLEkNoT2t2JYH19kq186yVgPqIxiIc6BE39hw3f
+44F4oENLoWsXC2ocdlwO3lsR5Y+0VqQsZ7zbWGq+vMLKhv9HkGc/5aQNzB4
QOyVHb5biGekfF3KxG+Gzveo+uDNndHpWg2fWVcRHNJE30MuNReNCftfSWEp
Q8GA+a2lQp+wriRwVbo46+H9eWSjFRQGaW/UzPCAFiz+m0USEHAAOdqRDh8d
vE3ttmcp+vmlFiP3xcUpGIYgcYzaTyezWkcRzNv+TJ7daM15No92Klp5FiIA
Z/phu1lesoGhjzwsnxrlWh9JXqTw1g7samo6j2BpRW8Nssnn6g6u4nFpxAmF
rq5DdaIrwKtIZ20p02idYP2h4nwwUWGjXo78Fmbd+pgerXe36J6VuQ3LfjqN
lNbD9QEnJrDGqfJVP4+E4K3g6YlW8SzXaCK8x2feyNGDCSToUOe1bm2obGIB
p76NwnhMC80FCMMHbJTNIOHjaiMXXp/4FoqXPvnvAMDlsDyPKDG1GTgwrcYR
4t1m6R6ewZA2w2sjJD5On6SyUSwJNjr/4uOMN4oivWv2xXLy1KNscC/8iMaa
huRf4v97gh+TVZGC1M6LXoy5Rsr9QmwmJa3eezN0IYqsx2YGE9PSnVk0GM5p
wA44pUT/VctX0EPgGxfx8b1JXkmk4m2VJQOq+pyt88fXn99bmzycmrluWzBo
GLF3+G8c0ac9un0JcHmVZ0EFIYCrB/LQ+OVH7cbgAsaS9fouBQ2ex+WwaV81
5pobeHvFfOYmi+0gfXfyyMyAGkRYHl60JTAxEunWQyjwbxHJWuxDGXxyODB1
PsbRQT0fvnmhCbsIFAP48K7zZDtc6cOJNqY+kSMU9lR9N3RjMnzIa/9s9n6e
AVHWK6jczuS32XjXyK3Lc4Nh9g2UlQFQh8NDjaE8N1v5GiaboGijsTw4xv5T
3rlJN14uCIN9fBeWP8vJ4miEfKFs4fY1LJx45ac8XWl0izACvKMx1mJ0uF3o
FqFkAIsKIDt47GQA8hRThhKBVnGhq0nytUcasupPTALxLuxxrGh2cOsSp82p
Tb9MH6d3cIeaEa5HCTy12ZPAyvZrMrngJNMauWCEFKd0+6BlG6pBqZLrxb9u
LpvaFoQe3whZMKv3563+n2ETOFw+sFXsym33oA+BD3b4ZDT67CDGVf7AWaLL
865QwG/dbskdj1dc+Oq3CFkHfdtd6HzVmwFVkLSlTcKFBEW5lkxlk3SBbrGo
NDDr9B8Lp/oWM+WKxmwTHTEUAiQd9q0DhcDTNaBcAoZ+xaxdr/7H0X25xm+W
nypj/jxBJOZxJ+gbOBfChdI0Mz8X7D0xjjTd+dqlS35rtzQL3ZRnoc0C/ZRv
xiBjLwgg00Kb3bT0ac60WxzNHjFSZKS7tmk4AcvpLNMYwZwpR3yEsGXM4Ki+
Bq3Kl/QHsK2px3GEeTpOJmPZtGUQjl4mlqWuFLkRtjzPvuVdZ1+fES4WusYh
I8ob7Dlk4hMfiNXFxswe/J0EBjeecUbpu+2vtpZZ/PSKLrhv+50RkkxMb3Kb
j6QFTpFaZVznBkv9M7a15RnOJ+g38zQI3isF4R6w8TXISrk23TU4a0gw6Dd4
jQzknmTdxcV3qon71Bd54RFpTkLi3ucrDLrkB4B5dvd0mX04K5ZuV2zInhNu
eNA5B649WHuQQAtlYB2x586vVBdmpLitXVrZSrbivch8fGBad9kVAFJXJbkA
tDbaSNWluPMFa/lPiovPiTWvjkVyej2bZnwPc51xjl0/zth+u+K4zu6cOZQg
yaoETsp1XpSI9OPBcCBRfUiNEqJMVq3nNfs4e+KSzeO4iyivMLnjFlyqRyiG
quTkcDCmcAmG7gaXS6Orkyw1uF/moNiWquOUty6FGDQ/C05gh8Wdeir51YIB
w6/INlVNC2Aqop2sHon8dLGXMUjIw8b+E9Zmmko2pV9vLxQO6QsoFdnHG3QD
KTUg6ZpCHjo8di0pdtiykl1hc3hUS/k5nsOJuukA2ErvAp3aQng9vnBGfDAf
c/q0u8dTCQ7bg+FGzM/GnvdU/EuvLwrViAYDwK4pKp3NzjBb8PPXeG5qTHkx
mISvZJ7Jt+DGUEdGt5etIO6y3fHG0NRmxHUA36PqwbjoWoS4oTb189NE3Jm7
sCSUnBHzjIGm3MtCIGAJ9qljbKNrNYPNuYar83nDbN5zd7O9nHwLDIRD4UXe
MjuflY8imSsMy92V9A8aMvCU8gHRDujUNQXQlME07upGRsvlQ7Mj93GsLr1c
Mci27KhhobhdaOF9akIEjtQHYNrxzYKBUi2imtjPOF+s+Rs8SjBLr2XjMuWE
rXfuzTGyeJLNJhrnL4V1E9ZCHp/pLBayDPxF4ptf/eTzOU/0CLHDBC6Uwbn2
R7xJI8LUKNFY4dDeXwUdhEDlEUgE4rBXimqb0aHWdI7gODS5UNI0tAgx+/y0
XJnxhbY59FM3Ae+Ol0sDSh3jbW+PT204UjkN0QfS6q1KTFVZqj6KMXAS8xMy
FObbIv9ggqEPiDTplQjcAhNGyk4ijnZ1gc2+jMBNhhoiQzNr+QSFbThBKuP/
B8qbD2c7mO9PFLyFzQFHp4VoKOKdbrJvjtU22RmCqjsoLXgNi2TRPXFbjPfX
qh2EGAIfBPIwupmJtnmCK3NwDG2a0w8KLuaM6fNLA1jN/l5LbiI+QGehf6dZ
5NwfCuHDtFqYpvhrT7o69dpt36fKX0ido8N1QrFlmvyLebn73O1XXkXC5C3v
rP9vtEmko5s5wq2ipEzaUKXHJ+nY+qKl7Jh/WQmi8pzsOcvU4h43KgslgqJQ
6DPLQhrgKJFqmhM/lHuizwlmfYYO1A7/6kLS1gU2TDY32T3FXtjkEIRJYxaW
VSTquA22i5AW6AAZV0+Uzff5voDgBifsf3gsN4ajb+5JPrS4cDrVuEShjrjL
2yQkZExHiKJOtqxOJJyZn2l0P1bYbCMPuNrsdL+y8hZNwo8f3hjd6uDJE05k
DCg0p4UeF0falJSTqCowC8j8CDAYe2rzkmTh7AdE5v4M7WHqI89jh/xpfrfL
5xJsEAyfXOXzCa1bLG5g5XGtlbLjP0lknlUCc8RRvNbSkLAASnSChIgjt+JX
zJOEMI9PtQv5UBHKfvex+o7J88aUZKzz5Lv+j5bmHkteybwAbQtWxX2/g+MU
JA9OhZY9tdldMaxi5tVyhrMqKiNxABiVV8PRB46CppDhdp74Nn8g4Y2yUdwe
pn2/LydaJqXm5M60IdkhUsTpre7JBOcoV5ZXKZei9VArizYnm7E+QpgbxP1s
yf/o2/uEmu2meTQ2eK3qoEeY5jV0vU8bsQcLYUCbVvh7PyhwHNqv2NmRF20q
gHpmBikisA+JUGHLVvCr+MaWbr1r5GQNXcnqQci+YHmDclfGDkL5BHxb6v4Z
stgU07QTpuKrflaItNQz9dEQSwD3NDQ6oAxLJF0crK+sqyvl+94Yr+W3uWCa
n+6SCxnW10GM+nQOU89gYYvR7/y3kRZnD4dpvcm2HC/2w1cUDegNqE7XohsO
FjsTzozE1+/ejDZw+nQJn/X9qtWE6cQ92UrR7iuLGcE54vv80+eq1+b30RXp
B2gG9+gAtEHmmZq5wg78JUNWeA/Z4OTzPmk5NJJ2JHp9Q/9mlMrL12qIAIOp
4xq+vnFG8Dwdv9GsDK1SpkebpDrJYjdwVY+QaLkc00ZRXlxe/zI3k9Ji4+oR
8fk1dKwtt5tWOxIxP17boOyvo4I14Pb5klDTTuxNfLKaIoe4U8joJYGhyWZ5
PXFDNuaenjI55n8vDukGvaKFxHIB7nkCIOi6iij8wp1htes9WU/DUT6faqLP
4P2ry1W77QG8DLfd3lzrqTwqj95N3vV11XR48qQihjkI1ID14/jOClN7D1en
/ekg5vh3cZziODFlI7UytBHX4rmxnxN1Ci1FNDlEc68nEn4s9+61DqHDHtlm
s+vb/reEivGRoS29FUU2zJYlXP+tyHR5gkEGiRZbifHekxw5oCwOjZtZ7eMN
ygAP/nYnr7h9reEQhrY0AAJzopUDvLMm/HIk6/P+v7Q0davoLJ8xNDcTgbQ1
UYQhp+lToe1gx7ew0mj+ZHeRvSxwyy60ptswnhiiPcsblyV47OaroKmkKtlc
UdE2I4jBjj5SzcCjooL2tuQ84C7TQZyIQBeD0AqA9JPEh7TVN0zSjyU42YJ8
0OpZlBgs1sY3bwhC1ox2PNvmP2h37OViFbN3+hUFOUCP3v/4euD0oywlVi5K
uSvENNKBXTD3pCfAl2iDdgoR8D+2dklo9z27glTlds0u8/5y5VojCIFy+EXL
0FrSZ3sgRAdJJkahXXL9C0rGraQZHmQLh/XsgedmdwusyaFQIucOtmWi1yT8
CKQnakHxf3gjAEcouk+a3DQBA9D4RwjXrUvtulNbnzVXZxz4w8SWjp7R6KyV
um0jmmNN4zOnyDbNWqSRRg1qoxFux0er2QC3ufCOjofFFKBSgHZihF94gojt
PqLUnbZkpc9b6MpoKYzozhHl+ZNbAkRTFKLOVaDK0p/2Lh/UDz9bKZjdAD9C
1YAR+nyhfgwx4NZ7+sYO2ndoYkTZKJD3YrT3/K2ng/McvwqtCFj3tDs93SwY
N751yTBy8KsPfI1YnJBP9qdlWvLaPHT+uEE/mEVJKmzGul5Ev8lU68PT8i/z
+nj9e06HVTkkNwdRtyOpVKTzT1OnZ4HGZ29pvhWtPDzIkQPS/x2yjELyQLal
k5xJLK8zqZ3HijYKxseVj84hrgNtlzYDJCHRAdmPdIzchgvUOJoyDe7VcNyH
ZiQcIeYB7ojQGxNW4YY1l0yAVpFpB/Vhe4a1ql6NH3BzKEH/CgHRGNXHKbou
VgpdabkzxG0gQ/uxwSdqlV9Mft+jsdxxJdOUDHt2M/QuncZdAxpYc9KESSWP
Za1/b341dNg5MXn5mzWhVLcIYLaroDreROSaMvzEjD8kAzyu/dU+jJNsPxOD
YPLYyShCMnSd3KoQ3dkUYgi+i+cnD92PZ7z2KwVq0cHaCYrTu/gTyPheQUXq
lqcDn5X78RbobXSxwvyGE2Fm9IN/qu4L382mEfECvJfIKb671sk62xfLvFMN
qPaGjrwcXxFAFQUZvYv9pXD91lTFo+Q2JBwXvUofQTmgTleR8O2NHmSx33Pe
RYb2rsBPxg6Uu9gauE1OcxnqQIHHrtBAFPbz9HsDnucOTSA6JjhSRP7v/v69
a6cLHRoOyS5rDBFIkKvmZJ7h3Sv2PxQRvspU7vAQ/YkiXS9kXKUsBks/RgL/
QMOJxes15VpLD1yghkKDlhZvhuWOaU3SPU5oiKbVZ/46se6Rf6NcmOO2kmR7
etUyiY2iNwpmvA8WQ48nFi/JAC5FDFa/Wx96TkfDXb3KIvuzIuFgNjPbyuRI
pW3vC2Ye5azq5Vr+7Idp8TJozbs8s6QkQkSp1Vv4RDjPr4lxSevfvOzXMOu2
J9bRJFSEzcEW+h1ooNeP4wJ7zjtoAIN0N/c69rGJjKn9fSgrxBdcvc1fq3n3
q2e1EuK64WjZ5OsCKBZ9i/AYaGYsf5NeHLEn8NdXnw/wx2lkMRYF/jOC6yc+
lMjtsMxpVDyiitq5Y+eVhYOFGBS2Im2QsvImiZA/nBohJxCCsBbYQkRxYyur
t9ioPeG/s68I4xPPiWxIbMAdCWIDhmtXrqQVwRvsf3PqUZFYBs6JVhqR+eim
dVpHd9gBXemBBf+Fmxzle/kXmOw/AmqtBfkvf+atXBlse8xEox609z2AhAq0
GCfpu58IiW1YtePNYOdcgW9dA6uoxn25bCkobM98pCdbSZ00mvDjCobck++j
TYfIaTIBXL6CALBZViQd/rcEv1ZFeHDdn9PEoRLMeINBqCQZiz3xLXA7k0Uu
1Fr5j+qj2uQgGSa6+4Z5MhIrsTSC/cF49gq/mWQalHxZKQcot9dOXUYOl4DQ
QYidSAdI9qBZPWxFHVqpJ5UAgzsQY3eP8cZOwN60NexxocDKjSRGznsm/LG7
rWK5hb0IF4NLkxWrLJ2TPUEZbIui+XN5IQ/PlxvX8PYBBYttK8q2CqJ3z8Ka
EJNtHkGsfCDDyUdw/TO2ugDZcU3BmfaoE+MqE3iB7B1djA0tOVM6i++vQ4F0
JQxbx+A8CIvzpvxziwyY6oMRCaemBPHNoVJOuVjUx61U62HGEeqih0x8I/r5
6fUUnAnaL0OruYk0CZwbq7U8PATI+XaWMWAQLO0LeHRHSMgLxTtD9ZdBEeQc
RpiTFeAY9oLqJVeXQtrNo8HrmjmHGpbCDfd8+nKZIo2iMxLDL2b9uLnRAZDV
hhTjoO6xfPGpQl3wXhx+M/hJFk65+2JB0jAB6wBUu+rfcSsA7hhTgHQ7rxF2
VGvFfW+oZKDc7C1jzOljZBEOb4uF8A0bdzf/QKF8/IwYd5Q48Q54HA+kV9FC
6gpIeGCE2E7Oq22IpTOkUG+wOXYMckZHvmceBZib0eKyaJI7PzomtGu9CJoR
lKE0+x+cp3pU4fSyLOnxFal9HykOr8JoSfXtcyTeKr9yd7Kg1Pp/jJ5tUosv
nGNfJA1Aw+I4jJP6K1IWe7hu/TAd2mgMI0tqB0BG2P/qz6sqkcFr8QzTm0Wd
O/Ctdmqa1PW2rwQO8ZDJnh37idUEZ4bpVfPzFw6MngjrD2GmeM9vlnPHXTjr
XCl2AwJXxFuNIy+hO2VCcUbMuD0LIrRI3fa1Tu5G4uiCI3DpzdnfxqFX+epT
Prk5Es/cr+PF4kVdpo2fGDgGwKmvGCD349RWowT1UEL3bvzEHOkLOLUiC/CS
lYHk4/+hVxTRzUz7KcJs376qJcGW38RBeFN9T9LIGXUaue7/cuMvSv3XPpMC
QQcbs53hrqFnBDzeMR+Yrt2WaJErBqPPdloNlvZlF0iw2YiJSKD+zuKA/Muw
69BvU9KmFwdnwX/P+4woRRVHl3hLaSf2XVfrwcXACw2R/+pS2TfPtwrdu/C7
ebIqBuwujUMbxRCDkiYG6OX22S1ZmJ6v5h9YAbYQKXnHa9wQD12UbyS4h8WR
85sBThgsQdDQzWV6GwH7EFwyJN4ihnkti35qd4mabYPcnznab6vH3lJLSViN
l8rbc8VszUaxq1PxlXsfwdDn5+8gUhzp8aCLfLu19dHB0B4GGgp9cgi770Od
rF2mqWEJixGx6PFgCKv1kzicZCbj8qLq7iKar0LaqnxW06JVZSMhhLTIARG1
ls/eVflr9OO0SnNvf4NMlZYIho69mWfimRRMOqjpqH4kAKDOU1PtbtoCxZEe
4BHXPpI42xo9OfLmWTVZlpU6NJb5b4zdyBMNMJldvucgjZZecfOlOpfYqM0a
808Gz0OgUn+VTBWEnlKaGWA0EpBBxZI9llSRiZ0BVAfs71QasciZB+D5h0s3
F2tpfcxvM9tYupH90Iko/Iqk4Lkdc9DqEJXxCY3b3+zab2h4kWMVPSAAmhay
bHLsrU7QmO6+8jk98y/Zcj0kNl7zjgKwc5RSZp66fFdSODurmbpICp6/pRbC
Kp6DJdW9mHechcC2GQLhuh8qVXy7ekLBHAgjkwwJmsbJKetRxpQUWZP/q54Y
ld8/j78JN/6cN6KiJxdVxP3VHlKIT4HULZZ6/GXeoXdrbr1+Jm6jhwf5LcVm
Pls/pBPsWKYKkH5RsWi0uXyDvsRj81qUtuE53eqJyhcmEsiG3ECnh64nwLSa
agSTnb6eO2GNtsJMQlXm8fs6CO2vXreDDY+INyKtNyA4dT1f7F/77wGAzXCJ
0uy75M7aAM5Xff2WjwrY3xm3bPTar1s6HHxQIjRpajubALiDQbvWSE/k8WtQ
3JmXlbAqdfSsZXsa/qmcciuR+5MElgYfKKEvSLCZvimRDPh7K1YcNaG/zas6
iFmRa9bEyNHCkC0CLVOAqptJUibAayNQfSkFZ0+RhMJMevguzw7nm8sG16pa
T6PD1wzhL5fHfvJNNFyXzYmo7L/T8myTbskyUdQT2kxcD3aGS7FS4zyFVq9A
HD3tebRrj8d3zD3GMPh+TVTqFCf5FCFKKhtbPsmZiHHl7UqVUH8RhDG6Ot3y
iEEjdPWTlHUN6Dy8bKahxLaOzFCXarkP9apkdqxKl6Ks+l/EP4FiIq5WHg6v
ffrEnmW4F0OlqHqlN42oiAAla9/23CYS+3YnaVu0MEA67bQsyp64jUGUUd2h
NgFo4UWYJ7/PE8D88y3G7z2TPqO/9Xge8zxRxT+ArSgq1nY3udzC2Zn/RiiX
AWl66iLaUa8rmkCvsDLmQglpRZEiDGg2KAId29zqheZyVXMdv+HBj1wcwu1O
6+Fd8/OB6G/wXP6rAHQ1QmWw0efVuTtPgfFb1m9a/GaRolILcDebHNwTit7J
49IAdfpFRvodrSWjKyurMqMtN0iJPIZ1C+X1ApX81d+PFN3vzCDiuuMzbDfI
Hm4Ko2SYBuQYOQ2GVfvXGtlu72I0ZpTPr/Hy2xXjtcJMr7RYAWN6bwqVtiPX
Uud6p9A2fU0nNRZnIGmWPEQpIm1rOU6wNzHK0cg64MRypu55bx6d5dcZzwuG
UuVH8oxiNrXJxUssblrFH1WKJPNm6m/c89qe0nCju5AcShGp0oFaVOwjgmb2
w8GJagObnEwtdUsbBmmntN9lrbL1nnWn/lncOxH6hJcqHJhYJpJDO/rl0kCs
GkMFC7OsKspmRLtb0TMLuc66khvf2zRUK+2BDOWM2lSS3bHY2RYzq7zMPy5r
wlcTlF7/5NlnnW9yWwvv3nlCmUo8nb493g8Yv4DTObX+v5WC9sOMZjyXABBl
nIazg/WffGXNRpxJCelzF3wa4yef6XqlvExJ/KE/rGKniFSacOXTaF/FG++6
bFTQ3TvdIZcrYCFucw/bqc7FqwEAeFFoEep1ledc6zl4cqLMVFOeSZ/ektC0
XdPPT+vcyg95ENq+mQ+uEwq8JCjnCLsT4WGT7tSWekUGfQORfXscJ7GTxesy
1yThB+YAFbbSsupPmPal0Mb4iuaKiX4ZA0Uj5Ql++0yXV5yPbmiWeyC2YprW
U3uhfNSjyQttz3opY9sC7MRKJ9sPTnXh4ovEMt3QTO4uVd7mscUlFlKBhuC/
ZPeS/8xrSbCO0WhA2NdLYXFs9djfhxSzpmwDmHEH46btywJDZco0SbBspiu0
UVbkz1+hUsVbOmtGuj2VbDa71nB3QaGMfdiNQL0ZspzRy+LT/itZHnWTZCQF
VSRUil2d/+I6HKdRUClrwJhn1qc4AGdrZmfz9zvXUq+V4H07p8FvfymNbyMV
DgABDThLzY3AEkZSpKyd02pvKl9iHvESG17JsiAeQPBw/gJXSkIPAoJmDzJ1
DZ+Ba4RvbsY5boH6cgylcFqg1z5cAK2lxEKhhE7fYJ8ZBxhAKsfvXcQus8lS
w29c4riCtFfzZ0sKsdxctrYsALOIS3cFiImH28rDDWyJtytH1QyFz4vU1FtO
dC9j1I6eZfNNdvXm5Pc+d73ECrAx0tnQCDZsVo6vJjQLmbdBNLNUji+C8z7Y
mYCvZwZ1y29BNlXA0pICaxeE38UT3H/mx7EFK8jCI4Hquzz7xZMZxjfxV9pl
HeKB1pFvfEdxwGShLp5aLzlpTNNQUnZeZfZS/SIqlqMBjks6i6r+GDRxo7Fx
ylMni0489DrarBCXBRiR7ad9cx50su0pxFF9z8k4Wgq0jIt5bAzteY2uLFdV
ELAPo4Z0OuDz0ZKAoWlbWvTyI4p6ic7ePXRaqNtFuUAITStRJpLP0VrL0vkc
jMSSFaQLCttMPOYPV1iShsedK/rTSFne0YRf9jy2Ou3N+qP/IFiCbo7T8h6z
TULDeYSF+It5bCpn5NGih6LG6TQsLCdh3DXyAIcF3HrZmWuE3jcWTTCQy6e5
s1ywFJjenC7uaSH8nGXVC5pXJGEI5vEAsxV/9jKxnRuKdyKHWCazLRsCwdHR
knbV/uKgX0Fj+GowWF15zY1U408UXo0KYRZTES2FOt5lIBsND1HL06HymfVA
ojT+2ldc2RYd5iPy4wXGonDJnb0/5/VJIDtSJZiNGc2r1vbylDIfU7GCAV8t
aCKnKOAiolX1xB4XN8uReunA7mItOCyVvjbpfY0NtUG/STKKsWDCRt3n+apH
BWFRV+E/PPxhZ2a56lq0g3MQKBLfqJ2kEtgDZjPwQ4k4F7qGS0p42FeF2935
T1pk7HgGPIZR1tcKpVr7VPolk3neP98YkxgQhCo1B/YTqMlRxy5Rlr9fqsjT
uclM1gz+7e+BRJayczpa5VbDMGEHEyJijx5liw02hYXkxiEyV9ib95wRWow3
th0ko/Wx6SvBeR8m2BjQeV5wbXWa2TJTool74yXk4EHl6p3ejs+n0p26MyDO
SCVaxQqBrxBdjUIU3RMRNzRcWI25rlmlhVN9ddO4CiDVrTi2WarLY1fxrlDj
DFnu659zSpDGcsSL/IyD9/HYZqM2SOzF4TNKWKZA3p5/ckzU7jmg7GjMfTUa
wwfnGFql9sxF7a4Ea+L/0VvU4cKYSvaviYLRyKOybvbzy7nbQyQ+tNHCV2WJ
1HXgoJaL/iX02PJOV37wicoS3wdb4CA4/j+6S7MPURhb/Y8BGoDRAKKpU6hz
BmRC4nck+5PTYAjI1VpqUPuf6gBpfWqWKcxmONVvk0C5jX66VySMsqcNkgAP
62bh7uCpDnPNzl8tXQRmqmAxRS3q7HMe+uFtubnjjlFNMqtyheI1PinxUH8T
CqjPTgXuz/QnXM2daLZWIwHIFCpnOgk2p8zv5wwilGqmqKlTdAxmnUXGDXiA
Ibahe352f2qVeNLk5xHEvJZiPAeMl5+PvPx59iDhRDXospe5ujZL54Gi8EcK
As9EFQFo6h3G5poI5QQ4EVaSBnVEQTL9RnUVwyBG7LzC15LnYhIs+joV4GJr
JkDiHWVe++M37pD//pzO5+PjwAY4xu2n7Dv2ljycWcoz2lVbny3yhfI+27j0
ovG2xo9lgu2VWrr/FH8dbdoWvOBt4T1w0U5usnNvd+lOt3Y8WbhzPPpSGx/3
MSPFvtb/iKPr1s9Vk8MorI/WoId9/HrJtwqa92f8bSdvTsUTK3I3wZFjAmwr
l9WhFjNAAEodSVg+rtnHCRMy2hcrBDnn0fk+FkSUQH9FUoPvlWANQgSGmgXD
Z5k+B24w8LC9bVn/rUqommaH3K1eQlfKH/+zmxdtD6FIu72h5CW3CzH76Gtz
ZXVMY5UQ6wQZVgIqQMIIZgWGTGSNh5l2KnfHQqYiy+at29p94Iy5gwRhzDB2
eG3W7uz/+Bf/W//E/TJwxeTKf//AutTiGf3/j/GV4owvitUOfWsU/otI+Z3g
K8s/pYvb7YmfehiIoCl+THFS1/NzsT/UJhhQb03ArnXmfOpXzATU2ftxAplZ
JCtauhcWTkNNS8UwFAInZAYESucZ48ZBT47psLmpBdwzKNHkR9ve001ALI0U
qUXsFq/7+gJ3z0suVj2bbYWIFcHcGPbk8D3kSDI93YIk+abPA7pmHeP1LbWS
xI5Z6vJ7kihl/+DUyxuXKYg5hBn0fi1ZGD8EKSncNRoVGCBxNgJurDJhfoPY
n6xIZ2bWs/b3J+7m47qHpFUG6jTvZ4pjdG8nAedpuqjdI8zeJ5DiBBv4rMA9
AeFLSph5smeKi09hEX48ntbIOmVb0s7zhEjfek6Y2EAnj4Exyb/NXBn6QW2j
WvP2U/VYx4P/EAuixlwNJtxzGm3dw/NJKq92jmmPz9yUvb/0JAOZIahpkukT
LsAi9a+XtE1fcYqYvUlfrVTw7s9WhFoI92ASH8zRPS8jaJnf5uimRfoLWCiG
Nt62B2v8ySKeJ/Bi4r9kJ0I1QLdfg/gPO1WSln4zKxDa31MtKgHqqcifCsn7
MavcpUIfT1fefNS2NHkx66FTgci81nJrM5SeCD8rZQejc1mYdQKXjMF6+MhW
bFql+4MEF/WRh/LNZ56GqEMJpt0wk1FttudMtUZMK4EgmkquKJkux5uHxywl
86jHl4PcYhck13vesIGyirXVDa8sfIc2YEG1BKVaeU45ci1RUEDhsCzum8ok
DLmXRYk5vEYDNI3bEFM6abjqhjEmEMVmVQkJuTx42eIQkeqtcfMsCsP1hCIu
b9zJ/49A68yITivY7QoqhFAgYjItfA6zVhDo0BBHu0mFS5GtARcwKqB82JPi
OBvf0WzNsRamhimCBOrE4/63vdo3C6D3rKEFZ4zNFvxttyOQb8/1zaM18Qbo
FBq+9L/LxJCB+hazpTaHEOdtvd9DYsOoEXriqil5LJ1DFGX/SLdpu1VOSs61
8bSuUG/fDAEksHXqz8ijdn+hwPJJCw2c9jvGJtojFWFWqaTS5loH5gyKxdwK
fo21fMNuexnlH838eJNjNlqttw0WipAeKihONS6gv+cadzaaBJmMSKF5EgmS
1ManjV3u9o4BIQkEJ1s3DWpvzFgX8fsNVznrxNSd1x8++5mTlQ3QeFLfoO+8
Rdd178Hf0W1CJRI3NnMLMwGLfbIFqSUJamCUUKFtK7ea+ioqJBquCdbyInpG
S4s2Z6cMOlXD1Gra3zPncniJX+thoi9P5yVTVWCay5yQje/gQx62Nr2ceg3i
XsbPUQG4TZ3EFJc0EJ3KPXjaW466irAdX7ijL7an6FWFjAgeb6jRvRxJ6uKS
sOYwKzM2MqH8quNhWjwfBJHqhmVk8jnCAImvoixBGaryn/7VPMioooLUqYLC
uWFzcWnj3i8dStJvanj9dg+i8sfAsTsw/O+Bv0yx0ULmRL7a6dzCbyH31DLC
S8N9eENg8OaNzddwmMl4/E3OhiLyvFKFhR2YSV/gOmfmJD/AK/APgRS5aJDm
zqdW0VfXC616Ov4DsQw1YOisIilBkiyhW6c2LS25SbuGSew5ZRnTVdiw/oHG
msipQMPKh4qyQ6zV5xyHUlLmf4tdMKHn2sRMe6GuPOhIG3ncGAxW2Lmr++gz
X2RPMrgRvekm8PdWogvk6wCIjtaYbo720X83uRSfzJsBnNjjD54+EGAMmfuH
rvJ+6H+BoEhWW/guUwxNvQsUcVhFKIAYuljW3/sHx+U7zFIRRSdj/gvPq1GW
du0neYHngvgH6ZiKUZuz1W0AuwGlan1XNcDh1NF0hyzWYlYmrZLQuQcrfuEw
9F988K+dD9QEZ6gNdWuAQ1fvZ2Q+nbdJxrQ2OcBUbV5md3EdWDEGvnyowr7/
AGI1PBMaF3R23i03RYAF9ofhJkdbGGK8lEBgcO0xoiomKJckqhdf2xYJSKuD
VUfdNWcw/u09VYug0mS7Le4b6ZmAQaPmldu7rJX4MNv3jhdfvcgnS3lUwIOI
pZBsuz3HQ7tznoGfqP95NpvsnuOYnrmHrtUdSJNKlXThko4pbUUlYRz7/Zk0
oopObNwhfOQGnG/TNilGReQhu/RlGjZmBCqSd6g7kzwzVPpJkXOz8BJSHPGY
Bd8oMg2G+Jbu4LM32dbrriF2F62M6mvcTTLNQZioUHuUUT474/G5D9I96WwQ
5S7zfM4L4OgdRrzCqDttbakAfSzKf9G7/nNAYx2+9dBgu2RGCs9Lt2RUAz1P
OKq9gnvRg5F5bBKSczldlSuVD0PxAj335qlOZMfJHYvOCEXpKVZRvsjxwsNL
9takoV731yHEBntQJEZpakk8kuBXpH8B3K4hT+sZWfPxgdGNl29KoFzHPavD
Lu3q70oye+yenpK/hXVzZ44UEAIi/8oG8PGrUH5eRSkjFt+ggcDC6LOO8HA/
w9L+rDUCI9F2mT2Tgb3EhKPjQya8qgz0fhxE2e4ZF4NCxfae46w38OqR0TlY
UZviLqEORbGPPnnDb34InldyfGlkqh7e/DvmI/HgoGFkX1ArteIzjf43G8zU
QFdBjjv1DgR8ODgmW9Yv9NdY9JNdFifmcBgnlU6F+RG/WX4AiXrDPyf554bQ
hLDdFICCc1bmkO/Jr1UElNwARfYsHp+P9EJRpuKbZpSRthbKkZ8lS1FVrJk+
8vFURuVN772VXJAjC6LuxM9FTekuKnqvBo2et0/1rip8QjTVXxiMFfVO/sdq
uTbVcscb2z3I8CdxnQsCB7notJfGA53ykBJAsc4bagMDde3r++wvVJaRzN8b
5FZsxrcvxePMmeOz9dHFo63qHX/RDHOFVbtyseKi+8CzcOISb3mjPomvER4Z
nu6QT35LGEvnCU3HJm3NrW3nQErWQDkrG7TbllhwXP+MqMinisHza3JzEBMZ
SY5lgFVRCTA3OZnUv5z5DvX0jm6GptcGaRbhe3asv6utFZcgf2c4HPNTU0GM
42WYGjpq6hQQyMk8W+GAZnL4HRXBkJ2L6cefFtLuMBG+Be6iOut8hxdKKaSn
+JfllhIyP56gqi1438dSGQ41ULC1KdQ8XKyiLfHU55WRsMJlcgD3J01twDbp
Vf0gAHYwIAj+UtMX4K/2yPCAf5B6I+X2FyGsuPs34lHNkFddRUaxxx7AGddc
s0CIZf7l2Sk8oBOnNlWjNlRqK/114pxrd1Gyml4RH7AGlXPajb0XFyuHfr6X
la2h9fa2EK/aIfBfsqNl8xEBwC6Qz519L57STkzfIUJskACuKHmG+29rBDCh
4ckFlkqptkvUzQvN+3bG97RgO7/WutXPP2DL9Fdb2Lxpd5RPpD07wYjl0QEW
36FlpViGt4NCJDNssvPO4hCLdX/UKZpKbQ+Qg3jIJ+p0Pf3txBDU3TLUMWCX
SWUuHd7sDHghmbTYcjOscd2snPZT/jVsrX4fZ6UJF/h1FxZc45S1TT8wujo3
lMuubn/YKLh8lSxKhnH/ydJommze/D7LusYji5EaCEfIzAyKQDFLjkwUbfkQ
4DKv2DC87ZcoAtUZ5AKxvHboe4db3PbSRugNjFQybdeGsDA6vaXMaN9sLBs8
ev3+9nzGLfN6ZVmTeYPLauDGFrYIPQkWtBGJ9c/xNe2lpsdfUutXrYeXp0RT
dCmucakA1sCaH/TtGHQ/GZksLgLtmfdA+HPZkzAZhrDzjaGQyTfmXy7yIQhz
aSSaYWv3LdtTFcHKXCkDd4C8hfsTITiv1XN5ub0lZdScosRzH+VTPMVsRT+Y
1wRH6tovvpn2qKYyNLdDotb99sUSKz/uOWf8buwgN7M1bUvMu2rZRz/1PMWZ
O1HpdcLRqzaYDnlUrW72XCT7OFmTboKIae/jPjrycY3SsXG6AfOtLrWYVAcm
ttJEwfo0eGfedpE2yH/KBhb0oJd+vZHeVDepy0LjPkl4h+s+QW1KtIPAMbZc
F66vHPiBCvExsRMxs5Oh4nI5D5qaNOKStxzHLSq4LW73fDYvQzlnHLLFd/Z+
aa94YZ6rZU0fcquLPgC/UCOvW03K0726wczvHVZVLYHm93VP6ROmoildy0f5
zZC8/cU0cfDsFvCp/9QJ5K8fe/7F+Vzok6OyXFlXmMauzX/E4Wk17vrJb+8K
Sx6dLIns0CDuEy1k+mDaTS3rNSv2gdnhgeZoAxkm7Vnc5u6eaiTEyxaGw+Ai
7t7fBLdBnwMoVI2F3zhhl+bVw2v4nSGb9TrPZiKUCcU7DEf/zYiE3sUdU23V
ju3pGQ3TMqTvIUU/R0p4nlN9uSIbMqwmkl6vCD0i6AVqTcB+9Pzt61kD/QNa
ciuT80LWg/KRifE1K/S891Qm0vWEZ4CMdOI1X6ZcrAWXVc57mVUR88wdTsc2
M787HrNzHAZYMflv0cviiCLsmWaiVxrE7RGVAGyvhSM+OgAM+evDLZRUFrE9
WJtrYmTyaWkX9OecUeAlAIqOHT+39F6rwQhWmdk4OBieMU2IzsyrENzdOyLQ
YrB4DpIQi4G0JZc/UrjvpPnFXeyWby+DclTH2LLLCuLXKmXCkrJ+zzYUmOKv
DKUHNZvtSlWWW8pusUozu9d8ndabLI4mx92cU0YdTeqDxPNAfqyK7Jg1u6t3
FZ3wSpq6Rh2UZ4he8yxcrVO25Zw01zGilFp1F5UmIYa6E5Xt1pNDn3WGZFJj
m5KW+HbUQcRSahS4GOUUV4Yp59vCbc5j+P2tTrqHdJUK6oXfJF6U9/tVqRnF
kRWQSC9lgP+H85wpPwxopuK127++R4kadnO073v6L3VL5oJPz2bcOrDTFtz+
TKVEIWIzbQttwXmh4QasfnITZ+YOvdDOAnoMsmfC377R/wZ0GwAd3ObD/z1y
5aMp8MFZqnb7QWfg4iqIkMLpfZtncz4+zZ2pR8peA1JobYk4MtKHVILPKiOG
9zfHGNy5tW8eSBYmY2bkefWAQpA1xM33b1j+LP+WWE8KyZOPMWQUk9W7+5un
XP4BTpqphCqAYzaDQLxH5v+kmar/xqQ7E/0FguNW8xdgMQBxJ0i+na6xdCON
y9T2CAC2Cb60ATcxXjOcr1mR6vXOLd+XOirp15XG34Nv6JPQjKGtP/v9ZvPT
OR0pN5XgwOQ8IoCS4bBUi6vEixd32rBeYQLlXI3M0Rnsrqg9cmP0R0IR5LBl
ZK3U2kSnRoP0cB1hoj4hqb9mZSTDsmZADGFGQ7r3SGgzP3NlfftCWwy1Fy60
MEYbTfmvEGecRalmOkuuAcPA+pJoBLCqxE21avB4/QhIJrkzoyjIy5zpWXay
J+0z/bzhzRK9weeiVdS2SDmTFONcLFUFdCE8wltFlP1rLbpwhi17Elqm7ZJi
EY7VIPN+CxxPHVc/i7v8IZkUgRkHwt+FJ5ONQnOGXmANnv7k3X1S6Ab9wdoM
iVo+8fiFsbZUXJ5ZDxy/g7t9Y8H50878ew+yX7/Dq40KoO/Ew94nHsBKmfoa
Q+Uk07tegSo13C7a1/uEOsv0GzPFRrE6XK7ZN1Db2Q7Ce+tyMvbzKyY01HGN
qq+yTW4Zl8/wfPPKXKTziWubmiJtpTjSgtGUT5wVDyd3r48loRtpSwvhHBb4
LwWrLgArEmoEESl4xPwKjbtse2s791Qb1Y2Rf9aSjIMJc3xTVAmWLgqQI9F3
YXj+wqNgFARip+PwHUEOTarcQrEdc6+YIX9CgLlE6NC07JQs+u/T40TqzJYm
WyBQPJLLHbeTnxWBMRGF3Cp6gfndELQtGSXHMxfldnvv4hm65MhQltS3Clj4
0vzs4H8tV4vnSEJkw/WiO7YDq+cWQTyvr5a3iry0pEhP4sTN0035wDnD4ARB
SAV+uHkdNcjoxblf8PbIMTundZy0//4moJHpc6njN0NAWS3zV1nyVGqN0E3K
sM5PNbQGXatv8iHHahiP+XcGQs+UEw73v67zFuwD3xZ9B8TabMcT/qV1Hdvy
0KzizEHdxUFatcTghEECmr96KRmS3Vvy8B0B/lLtnnwXoXg9c2gU2h+FojU0
1v6CFvMv6Z2tic6BTgR7XFaLqcg/i6pCJyfjsFl37zu3sNMUybPp+zvL4FBi
cu3ZrPHVMnpIY7ZPE/nB48PezZJ8kBIonMgpsGECy3BPYDGxl+H0X+S254xr
L+eWkDQtXP+4btFERYKK+YFL8+mq7kki3adW0xKzGCiRbkH6DL+3J3eMwznO
drZruLuQ0BRP33HOMOz1nYifutkUnpx6oCCvo/lRVac8yYDfjebTKTqv4KNz
Ahqnvo76es3n6WrnYbkifc8rRRZByl+4CLsIDBQ3SUXnJ9/2u9VFpo7ytd+p
uRhxMZ6Zy8VXJWwio9Q7Qq80N+QR0MvCISTKgQZwu+V6Wx8/Ekw36G7BX6Bc
DreUpwjWm1qh8/iha9FBcza7p349R1iqkLqi5Es9xpSKl3CX2ZCqKEiQg+LK
1zfznBVahv1tYYUA2zIrAtDYPb16IJac+HCHcG2z46YhT76UuJpMjDDqoDQr
P83Nl+cLjOXrm33ccQ7vz2MdDUjSFBtDdD14skMweACo4D8G+W80WTQO7l0x
OLpsaIveiPM9Tgt20H/0ozRJgKcEnQhOx5bqLrz2MpYUeSGRQW3bbSpZKh7M
qgQBZy6F9qRhpo/8ELfY+P3J4G3ClhJrmU6B1Py1735U4CtHLk7OotsybTH4
aZbXazioyUWuVYzr7MQBnI8WJhgDdXt0L0SQETb74fPMOsJ1i9PrsmXyBgZX
lMnQ2qTRZd6eT0ggmj6yIYJtMBhWvciljXLRY3tF5V1zWC5Kdpx1nlCp/e4n
ocwg5biHaAiErR/8qycFdfC8Z+i1+V62ozexVzQH8zLSaEuDk2AhwAxLGd1u
LlDFfFp7kf2s6eHEy+lwzQguMnYztny2bJC155iDsLnrbQJtrWoqHLfe8qi6
FTGkQIy6PFc6nYR625h8aIJp96M5zSW9MegcsfQIRi9+5bzkoqNCrXB/HEyE
PyM5aPDOAgwuLJ3Q4JgK3ozsKJcgdSGAXeowdyUlogVr40zb02tzseZoKdTS
KOdmsiZoM/45b8fKHHF3ikhMPeDcdh13lvsutT/cMoHAQMs4d2QVOVJNrtSq
JA4qFgO33aJlM9BZ5Ewu2/esRT+uY1SVqEHY5ZyQ3VUte5/3bTwgoPFxMpPd
g1Fm9hGqzMVQTSzPHyHbWCWP+imomDovVI3ynw01iVjDAPU2VKmoVcfu3q9F
0736vfQGSdaZekaaMkX/U4H+uORReejqkWsXBAirJEg7Wwb1d4vBNEonQMyY
g54P05Rsnvtq+AeSDSb6yNhjAoYbIhT//Aab8EG5HK73tzc5JsvrVpfJji0p
ayYUCEf5PHco9giDtF3wV1XC2ig9lIfKEUEl+JtSBk7Et8/sY87FbgaYNQJb
Evg4/cgMpvCN1aowHVz4ezpKsYKSGZM6ofvR3HO+XwqDXGsoYFTVeWqi3wPr
S7p774HdYHkbqe+89mpyeFTRm7YRDBkYfGEKmNIWxbyK5mqLZ0C6xg1Ot/+9
80XZC+ikv5c1gdgkYYzjLiO/gLPm7uH4G5dxTbWENdN/iH3l0pJCarKXNPWz
x30rE/46ccw3NzdMjhcWmBXJ6jdQJrPVJpHZax/LI+sb+avXnkTQa+qFU7eZ
11PUVASu2T9gcV1aC0aZ5LPCQuZc0eMtW8uII/3SFGcb6m4je0Xq923KB4nh
ep45NdD6QrhNMANHNRWyony7lGd5/ZO7lEjSEd/aLabJoQaT0v1fHGXdrD5r
utXjHlI2CMtssnyvyRy8mLZOY55TuUCx4IxR2BmYVhYbS3Dex6JHKhqaTKYW
b18nSHhXFcK0Y1c/DsBLW3/O+525GVnHNvj3yC5B4gdglawtUFQI+brjbzfi
3Nz3BzRcU9ESvucaRdlyPsAl2vVtR3mNFNMbboV9MhBv0UFC1uCosot+UmHG
L0phE9mQj1hujviBY4/c/eCNrbzUsq4yF76mS2jpbxRcbo9AeARJ3V2HqRT6
bOYRMU7sBZABSm+YV+qAs/eZHo02qT8SamRGmT8kcO73VIceiK6O37JcspRt
fggt+4P/7iOtM1Tw7K1VN3EtgeMsKqbZYEzdhLPcd+SOc+LTh6Is1t3ud2FP
nMlFVG/79qpEQgMCAio5G7gJFwL7D3pBfi5GbrNgsDRP0ZojTS6QrE+MUk1u
DqBC1VRQGFzyixLKPEcmt3zkET8vzcwCgJK2IG+IhrSXYNj52Kw+qjKCU9o3
8m2zFrC/J9LOp6x/M1atRwrw98ZZxLT1iI8aa+PiJclBuuI32WRsMLiThvdn
u0eqyqwn9Eq8LvcIc2AgZ/ClUfisez/uHdi/+ofTROvRGdS1xiB7ZP+whMg6
C8BhpSRhTBEMweBy/jrmAVguXBjfm9ZDXspgp2trAJhJftqRRwvIA4pT/HBs
/uQJ1TiOI+DhvkQxZ9ip1+qBX0jHZKcqdm8iVbQ/QaO7tJOjXjf1S0YA1csu
cCwxYbcP9W4kQt5UxI46kRROFcphZiihlt5Q3jiSwmp16ibThniHtRGpq5sW
AymrOUEtW2cPWSAtEAM12Tfn8rY6VLX+hEz0ongxE/LKRUpYYbhI/68dUnQN
6GGSQ3pBXuv9VoSCUVTnYNeD3QPnyVhfhMKkIPVHOdYpvYraOU9lRst2q/IZ
rX3rZtyTv192y2mUkXVJJl2ZjPHPfwzZPGI8HGSxYr1On5StN5dPD1ssosVH
2t+paU6jYdVkPiD9/5/rEiq04fGSkC7sh7tZ8ehMRAN+5cEH+tGdiBIDKsmN
RaSurbkSqCetduKCY38evjjnxx0WY85EuVACo0yEB9RY8ju5SHS8UfixtGcv
BYV/0ZPkfWFF9441/Xo8NuJGJq2WalhghZkKu2MdvDlZvCeIOQN4UwpapNcz
qWSWdGfzZycXdbSG2wdF9FvN4XtrtrgUMWFLx/RiAmUa14Wc2y/ztETT6eqm
LFfVRmny2ODzA7ZPZeStZvCQB87YPLoWn+gHDEsHWdPKsVuzmfUQuj/ONIUC
uTDRzDJ3zmJuKlW29nJUwk7Fs9TM6r9+8bdPBUPit7Tfrr+7V3DvE74ugG93
5rhuQFDKLxSSeWcD94vabN54Fre38MZm6qufwg+pFig207CPKDoDLrDHkji2
hNguSXdC0oJansY86aDoN30DvSf1IvL9PbwJJ/GjvXzaTGFVRVY22+9CfGtl
n9mFqf+IjBeW4+AxuzCZbn28YGgPLK6TRhXYhHPpsaLTlCRtz7v/hJSKz0NB
THZpxSQUmp8VnPQ5eU3oaOus1LVPfO8pMcfjlIZ+/qZ68MZzIlqxQme5Lj5/
acC6ic2ePjlBYL/OXDS+hFXEjE1jD0BxkicLkzCNXuITdEqA/mUOXXe7XR2U
BiehH8+PcByt/dkG3Oc8BfjeSLWCL48ny65bZ9uNfeZqXAdJU+zGRKWH+jKF
p21fo2K8Qz8W0iKFWvkZVx/6+2rnIAMphJVlmrWx9N5ih1DLGXWuedg9J1yt
hgt1yILgmB1wrDqwZs6MKdMDN+IcJzsBx3WD0WWvUt6yXu5zIQsEmcZgc/uM
XCKVHyCIAjHXtyYp+g8Z2wZ66UMPEzM5VGs6Fdj1CHfnreAfkADnWi4tmROg
uiKhSD4AQUt/LjgfiwwCf7SBlCwdRu9nGYrHNpOn2QkuC13Um++IwtcYTieD
UP0hjVyUldoFzMaLlOTAdcBMXap4h/yUUg7VXiJuLB4IGmJPZxlcGr6KQzBu
h5jvPjdIQaYyVhH6IGehI9p3lccqIu2UuasaZw7eKJxRdQbII9Vm3M40a506
sck2cnyTHnMGadqkKisuYnWDUfetfVOWbIL5qUIkJd6Z5Fpu74iLbIFNB9X5
iUUDuOzye9d6DuTIvxS05JIM2ukNmhenoF1PNWwB7X0+7jGbfrtz/t2ISzOm
P8CknlRylACuXLXolu4AJOtC11Q/8WTo3CL+WaittsLNxfCxv4xcHg23tZWu
GLXCi5/ZWcS4zeWL9jSru5fWi4WzbnGMjovHFCgeizIT1nSAJYW/p2MxzsOj
W9E3opkyJS9Zj7E8W/ZJzKquDJfTobd0yWdBxaR1MjX/bhvRJvgFyT5dOD0H
Mi8myeICBDTBQY6D9hRXlg3xshPSWuYiIoGsCYoymKl9dt7XHydiFbtR42pn
vHoet+y9ntvMedCpK3GA8TXeEV6nSov8b4X+NJ3pmfgTF9FwMlh5JVi8uBEm
8NPqbRTqAMwo+aNK+rw/7lXnnNRPqx+hbN0It8VMrL4SqCDeBpWoMXOp+rng
6cbFvcac5UadrfOsnya6oopGq1lWDIGxJSl15tZEoQioziyTWk1s7L91itCI
DQLZSvrAVFwL9RZz7bPWUBQVJ4soKi1lc6TWyJcbf8S/eY47kfnBH/izUTnm
oCMyh1Sd0p/n2JO4nFjidvdGEFUZDyxz21cipwFHdE/GjdQlQy9brevYt54i
3puTZVAL/cr4rZpaCEphRiIPC2olLOx66cJ4adNzNkQp++Xoj72AL7dspJaw
8Agf/pfnPfnkPHcLrRawmy3vbPfWztuYb4r5NZ8Pke1WzOv4a+x01omhbzHN
636cgqjteLIUYQhoN5T6b3R+y/kyqb2qKNTIE2CABsKg4UHUXHlqtqhDWyCj
bqXhN2qk4EbizZW9QG9bwNk/GUsEU3vluJboMdsiRxV1nb2Y3Q8+bYXQEs92
6MCJ8yItmNrShrpRVGAnfR0P6sI7arRcsyDCZ7bVPG7HUwZ2cUNVY8LHf8nR
l4RZasrTIIE881wQHMLRfzL4xH7vhej0ts5vhuQiBzHLb5IMy/t2jD0lPHEj
4padNS3jYdLyGkOf8ewC2HRBZEgncemTUEPcuJK1304A3T/QLDhRCjZMLROZ
Vz6s6BAelehDzioKjWLCZJZ2pokKqDlakUAsKJ3FmDSYvxuqkGizKngk1An4
43XXf3fv00vb1NdjAsrlau/tRvOoCCbKNsirj84BD2yRG+onkP/NCecHN3qT
qpo/7vPQOur2/cZnklwAtfop/CHsoRMHcExtSJG5brCcJJPxkDFSf4txpCuK
D2x0JPVFn2fvj0Qk4MvJP7HhzF85DCPm7Zsf8vtephuaMk3JF1U4a9wbDKiV
uKrldvEsj000pusOyxuDLcdWMTxCJcDTDc5YH2FP0yIH8LS99dgGg46tuz/+
014P0tQoIgznU/Jay8mO1TCCfLgnF/a4WHVh7tRwZsN+aDS61cXECsv86HKp
qmp5TB5I2/N/hc/g0gPU40J4IqH5ws5Od0Kn2Q+fp9gdlQoMSi2nZwZ0RU7T
/A1xKJxpM7uJAv2jUz0l/O7GP+uo0yE1h3ExFkNkmCAFT4Fe/TYQqVDtv4cM
r1xBYVdmbifC8d85oSzmBwTXSkclauxJZPzKMxSLHmlQ+Dx0ybJwlqIdAsIU
4qWB8m3tE4cNJGFKkSYwiBrOFiE03vcRBC/djyNUUVJ/RXnuT/OagROlZrlC
8ZO0GFeHdHQXk8zxRKI+HWr52RIDYHCWDR+EfKq1F1ZpRHcb8t3kneD/JiUi
LXiDN7Y0GmJZtPk8ukbiiz5JUasz0fBReQ3pIMIapApE40MrbzF1YW96PkQX
Hzn1eJBEOagnm9rQ/RMTfoH1RzYPO9I7Mzb5qgCL3d/XsbHxDHA6wBnSp8Mk
CWYjK+GDExzaecz4+8XRb0fYLS00YPsjGeHZl9lBrOSVJxURb/9Khr5w+vMS
vI5k/pFdieevZUTc1yb+UC+32os6XBjGX+z8FFTSXz5vrCoIuN3NCRzJXMa2
NJFE+xn+Le3f1Dl67ms2r5XDIMGmZQgoRzZKUXyePWQB2OA8cVY51c6TODUk
lNNueSn3RtbjvPEf23Y6I8FWsioOfZqVxjDqMuyfzMXLxQBILFTb3fbOxdKB
I5kcjOpw9t5jBXboXHy210ZGX+peiscuUv8ZCW5u6FLR1Aic1uB9jX4YASry
FiX4fh5M4whzqDf77olENDb2LNPkjJ2+DQTrGNPFlxcLoVIzyYEidaRweAl4
21PmQiPVy9BxNISDvE8YCkbyXdvPFCULNRLKgO0p3svdyA9lXSczq+YU0apn
U+bE1+pCkfWhvSaRVuWCBY689N1jb87pl7XMCoyENzYP8kjJnapHELSQdjN4
yiUEAfDk1H0fJ8U3zuAGW4GDGS8G2TdqBUPS7uIPMsjMrhR9Mj5O52no9iGI
xxZ0ZnVi27Ll9zSsjNP9vgdbfyoBR5k+/yno+YEGpkmpMpEG09u0UDfsSG0j
IRLDI1leAcJTbhxdxTUbixSWkp5MKL6xg2Jev4Ql2zh7AceEjG1GFAkYPSQK
UmjbVZX7BlujAE9iAOcoxrNA1FokFWcWpom5BLGplolw4rCqBaq76tSUEYVM
UYGxJ+hJOkauhKzZbq/zOmxBsTBH0gFxGfV0hhAe5bnKVL71/QiyRuNFP4d5
EV/joMycXDFnKrJ2JlAZjMy4YQUkD5pnQxRdcNSg0LCITbFk/k00cZW+F7AI
1mPBhMEdxafqJysMAH+LigjWUNEZZmJ7BAHom37KCSjkb53Y84a4HsWL7xgu
/r9QqlFULoOT8BydCN8y4NmqUo7DVHnaaXOBMq/bNosOouWCQ+NODajOt8Cd
J1pWxI5JmFp32G3lwwfv/DQqrhTXZJbGYWZIeZAP0FfhgWQsXb96vr9L/AjM
lfAodrFqlbguIP3Ej2flWZnnX8Xl+Ne8JZbrIO4ATbmmnjEz+r6qgmuGD8Kd
VHQWNDxZQb6sngm9+QGH/WBxP9qxMMxn7LO/Ld83RJt/KYfWYjh9DIDm+Sge
GppDtuxPp29D8RA9dzJuCHtHXAm8GJ9BGgP/DZTSLpw0P0nZLZ8l3fInROHX
9du7yPn83GnWFE/R/WJY1nmtv7a8iKLQAAxQ389w93TiZwWN+sdamyZ5LT6H
2+kbMQJkJIkYQ88Iqp0izcdCET3vfZ5K5glJZSpd4ARR5bKKQQZXDCXprF1/
s0cHYVG/RgpIYFCRBHtWCstCRSoKWDdYWAlI3vwCBiGXMTlKlOS7udK6t2gz
g9d3Nh1Hqr2u0McNX+Sj7lWs1az1vhnT6s2fXSApF4o/wLjO5EBpfAN0GM9E
LEJ4Qc5x43wOtcW3BmRiVAavZ/edJ/hAWKS5FtzjDtkX6dWybLVQp0C76Ter
zUuGUXRlLlSBS6o5gle2Ru1QRinZrLGce3NsQDcvW5G2sxyQ3WsunW1aciB/
iQSgMjBaszoQACHocnWdMMpgETjT6EPHGu5mAx2+0ut58hKhsixRDnTq5PQQ
BRzUVlVcTb+9sRuiJdDK9JHYVzZU3F++vEVmxMfMiMxm0ypsg9ByafzZfRGY
tSEtewlYB4e4nAATQC31r1dSUoRdwWTutgj6f0iIxOQUt0yqIOnmmFXKrANR
QjB4dXihZRBFQpIhkZoOwfYNiQp/eDC+poau7gYhSU8ETcw1CJYciv6T2GMt
nf3pTuy6/PX3V0XWx+0u9SXgq41qmZj9listLOHTYSjqUUas1BvtqRPMR7+B
zkKLY+9+Us/TZ9cGs+Eti7093u1H53BSyrWAhf0F8DSLAa+j9e9gjokVSxAk
FLKLWyD4ZLuu7hsbaSBeHO0h7UD8eqzm6W+XuUaeszvaekXr1NFSluwWyRXa
fHYJsEeoPjV+BBnaf8LqAr2a7PXg3J8QumwLhcG8B78Edh/1K9CJhSyxGZKY
D3JBjc9xF3kY1n6EochQ9iveOk7Lrg2qo4zLmSdfvU1OUn9BtXaG4k0XkSLV
rLZj8l7/aPhfDHLjs6fmmt22agiYYLo3DINWI7y1LL4PONPh8aa3pvbwozBD
fMB2I26cK1D1THb3HkELGJfggn4krPTotJ32xpJpZqEP622rss3egJKH7ZiU
38BVfT6bCl0NdulYTUzGrltNbC8gf1xPdPnsQul/eA7Htwh5yF27OFc7km96
5iu+hpPEY/eIjbpbG++aPcQy62RHkpvSr0xrgl+5zT9RcLMWkF17YozFov98
dNtQqoT1JGTSIpJeHd5wO3GYfVAzq0CjwRQO3fTT2cp2BOOjSiBhtuzMRoWX
sI2xoe92rrZ7n1TSYX2DsHPvaNSI3HpryD9iCDqP0ux2TP+FEYGkrAa8I8zx
9Rkvbm6N4SaQXE+xHWwQ2frVtZBoPhM0BKHKmApplXlLtyBolw6ipy0kLakq
YFeYPnwkW1OB+Biuxxy5+8/XbxvvRHqAgdIgzzclDU/MMyTswxNRTtsrTuIm
Bz3QSf+JvPgIqRDfjjDmsf+Tm0MX/dVOc9DqVzkVLHAAIDLunF0Jw8Aj/er1
wl71LSD+EE5beBFIr/ahJu1PVfQqngrb+mRuVsSz2k2ui+Vk4WF3BlX7fVJG
au3x/5ac6XFBE19NaDTjBRJj2l459CirRsx58zjSAH5jGHfyTI22CEtId0UN
pY1FJVDRnkvcBSmcSgUdE2MVSHoodLXXUPrDmk6D0ZIFEljtm+i9XAEERE6c
sZ3TV6fRAZWKV0y3lnaidEkQbr0K9aOyn86qF73ZaE1sfOT695ATDm79Xu80
MZL4ABbIVPowiH7RZILozoeguK4XD0n/5jD3ZRT3ARzScvzffm3ZeyQyD37r
hJp5zbaktqfvDbDo5L8YyR28klTu7WQXxMYMw5fw6cXGzGiAeWerv5gUs1IY
ER9RyKiljPp541pGiKV0MywngbyogEq3seelqcX8NeJ42ffVbw1OhN6RgQQF
Mm0uyKDYmAlHMvco/j2Ifu5Tz74nUI84CJ4XDnVmjMImomqloHtTjZr5K1Zu
rLf2qdDsIogS8Li3lIF8ZkOAmtwI3frUXbtTo/cM/fko2xt95yKAFd6rOz2M
QrWbzCDy7sX1OsbF2c+6BMokSwGEVadPkYM160P5i7yG3MJ34HMCN3ab7IEB
grxrrMqlhJNlUviyplQ3DKOkVvKEwX/gXl3NUSjaslfbcQ8kh4r1apYADSGa
SK9Z812bUsJ3t3iUAgDtbBCEGujDvlO7QkQ30602Go+ZySLGDSsRJBgU4ROf
lvbmm+51Zm2V2VZCT6nf4/5ZPPTw4lduF08skNPT9L90Fic8gQYIELHLvZui
4x3N+aRnjQyHrokbyyaiEv+Ik6Ax56FXTaAErHvQQLEGJjICII9TyO1nbPl2
EgHMbxNmgWbKupo1z6/EMiy42kicryok8zw69QBH0BWgrljGgZXUvZZYfGAC
9l9ioTNNaqR0L7Zjk2rTXp8JI4A/DjeCYLZbXsWOLpIjwkeS86KvqJWS/zS1
RVRmPtAFZTkKYhzoq62JGOUqmMprtfBI9J8Wewph1XiMoZhU0jDV3Gk0/tCt
A5G+Mg2fXZ9VXp8j8MW5azVYj/ovlwECEPgdoMvmuRNrAx5g86KPXvlM/HFM
8rYYhX43mJEaFDQM8+sMmG7p1zx+xN9qXHxjnsUXASGrcYpHir/k+tk2r0xj
xs9bZWLti2ac1q3gaeC+McB1CU7Z4USjrOeKHBObUg6U8S3IYurzs9nzM/5Y
plt1sy2++Y3O5Vf4p/BJwlDI7cpG3hIji5AvZsG1vgy2kMibN00M/HsJqYCy
FUzwA8psAC13VkMPOv4DakOc5xAqLsZZf8Wr002HJQw4aDNHgMh88Q5yCYJy
EfAJ0olL9pZWAiQ0YGj9jxoebSezuM8G/MwwshNLTsoJ0vANnDNeA6xUQaIM
hP6MVnHBMZyTYp55Bk6i4Mgi4O+oS9YeTyjMeCKeK373OKofnemCZpicGFpL
UXFbriA23yWXrXrCyPe+Foz1NFaKRZ0Wh56bDInL6sfMGh+eATncJXsp+BFi
H3njYvrAWIhJtORwjjVVqx6N8P5TvubQV7qc7ljdkNW+LbqhaH+2tQU6R+D+
Nk3+GitGEtf+mkuCI61V0RCSReleoNALRVkVVPI4LfgM1V6cNZb1QznPgV6+
aTEkVNL/lm+I3nGWHNy/inMWZT3LFxqp/ld4r+WtpilmC9OBl5AqmwC+irMC
aJfChFl95HkKwvmsqqsdWzf6CBDm3yi5njWdHkuosN6cAvQhKvALizn7kkVo
1MVnc86aPI6bxM2g9llSBAGOoisWUHN2FsZ2YQDA2loNgQZSHB81IT1DkN6i
a9oCV4WraJ6jg7f44dBqsL6I98IqhbOmuwk9mXkj07rzQdD1lKcQplCjAF4G
P47zbBGxMuWNIeY4hT1yvBbvPbd5+rckLRAhDlOY1gL2dtM3yfx5QdcNLrze
Rw4bj+AO/4EVz9smpSyHsBvjeS7Q7+CxhG5lTx7h6J/AnN656uPwtyIfaa3B
cGnV9yW5LjurC0U/85wk3MI6PDVj8fi/SCjSG2Gy6yHayxv4qQKKGRbbWQ+8
aCzRYU7gCZvULh+HJgWD4wuRkfPPFoXs+6ifMpfNZEJczEQOI3cLWqnZY5/b
Xu+ZH8STRssvR71jpRBGaKUJ6EhpsqtuA1GHCSeUYccpPXSLsTXRD+Qmcw1k
z01DSgP/QH8GqhCGAEO6nlq6OriIXYtO02+hl6T9O8YrT0G6ddEshW6YiNre
oP+76P1j92qs3xq6vuDqQ+kfMQ2DmARWwNgsr7zAZdBqHxEb7u4QKFyRx95A
7fj6uGtQLep/5FyZ+t7KCTfvyjGTE5L9YGxfzSkbT5PPdkXrkjegriMZM1K5
XvQL/EJixVmLANSnoWWZxwOvCmhO6UOyAHrmh+dN9JUrOdDBHx5Tu6zrbepD
75A+tDYXSCgdTejmQMDkV5WL5XFTDzrlhTKkaEv6KhCNtaBvI6LeGSoAGwh0
yjORuFGmmCExYponK1Od017mwUIFEw7OQQJ06/xblI3YJ+5M1t4vvRhYp1L2
sSBGZYX7P7v3tEpL54BeZERzR95hZX/4r1yaC1U1e5arlC6SGeWj6TY/4WlH
0ZvIbCUV6k6fff1UaslYbhaQU6z3z9Hf6fWtiaYoirU8EbXM2TtXQXu08xO2
IhYH0WT7zy7dvUtlN8wIin0+XFEj5QbNdjE3BqX0B4ACzAndokOiMHyKOj5Z
hDjL4n/3ZMjeAhD9WUuKdafq5gBMlDklkSEP9GiSv5cVWLnKIiyW/Sya9l57
E35yZHZwrhH1Fh88iknJpeEH8V7cIjVNsLNC8jFdqvWS0FxIyUJxyA9puiPv
ecNKvmy0y8q3Pr6V91zjt5kwvL9f0PQlGaQl2goKsNkm5ov4LGqshR7mQXIs
H/e9BuNbbX1NP0+rs70+jbNBE/lU4DtA16yiW8UgnCulLybuI0fM6kDhrkNh
Fl4kz8vbd8+kti5R1QnQUhBmLIN+YiyLwx3JfqUubi2h4MNLgKzKxUIIKe6q
27kGmsbt63GThdIFKmA1T7ei9O/OE9+QNAKkwOcQK+KNKeMYLw6NEt4ndE7r
h1iUZirNA5tLTl0Xphp56JQAtBnCWAe3fXlKFiknLzsnoOq0DhMY0vgYcviy
PPAeLDyQSC5swJyWDQAvNahUZS4M9fJmkxY7/0fUQpzJIYXBnfkeS/8OJIaQ
YvY6cjcI7o0a5nreEL2mnOW62HKwlPKY1Xu2idv4EWa4oQAj/MMjuNJkQBMV
QPXzHidMjON61NbeMM//WqL2ySEEknV2SbbquklcYgysHoEGsMYtm0dmlYPt
jVKc9AOyQ95cxaPCSzgPr1mGygiO/c5n8iRWXBm52yXmiklSAvAnKI0LCdkx
j9pqriXWTRo7ufkjpDpqdyK/nYxZ+VsbG8Ldiykz4LJnLVlWs8Tmvi+SkxIU
UdZUnyOSiH2rZaovun9jc1sEamCwraU+5Y6Ob84rReTYpb41wLkmA9gGGFX4
zilBtvApHxsFQcPL30sZ+FX0h9k5z4Ci+bjWb5MzNxGSag9DEHmQck6aqq5I
A9f6nzKAfafu3olBr3y7LBMJsIQCIPDv6Hw3kAErEMxAxWPS3hnqtzfozZZc
BNad4QtsBzmsyM3Np0yOM394CUGcqbHZs5lLcdYpXrw9IsEq84I0VWSd5dvL
3hcE3moYFXn0mB7bcXxaSOKJzvk99Wh+hZoWAcG38dNzqctjYh18q0dQve0F
X7MhQAL/3CvPAKfswYRKGk+UKrdbTGcKBfFFfEhVNV2yemGXmFycabOZS6Ko
BP9Ww0KegOiCeznRTBUnRqFIRWXCYxQzHIeUkuGD0ebvMdYP6MSyD2rHMXOD
IUSs4qYYU02JFJEeSFBIkK3UTEmB+7F4FZY5VstKRwTVIkRZrvIjOfM7Vvgj
1ftcDs1WiCoMhBcx2W99EMHlVRU+VRuNCeBVH+y38WV+cTPb2BL/t0XCUYu4
CSEutGex5OGbLg8XMcwMwuoWuACFKWwnc9g/GdqqYgvkQns545DvwACHGoyv
Nm79aWymqxPaGhFLv8mv9/atHzbJYkITFhpU3pGy0iSPe7HsGlvNmvb+Y1i9
1GY5dVKtD4XGPxolOhcBEu7CHMxBV54liA9Z3fEtUgi2XSUO2RTbVEgF4Ev5
oh1hh0LYPw3TLtIYVESjMOOYTkS5ZP5UKpAQVaQAjkgRKWMSc4sPcTmheJVj
yJPiqfZ1XhsZpr0DY5LFW2m0tl8EGCS/UWDiudQrrr+FaYzbltI3ME1Rb9uI
UM/cHqD7c4aWPMs+Jn1SaYL89vAiaGoodvakfL4J+9xpM525cT3ZHkSUvc6k
8QGs7J8KeR0bmEG34A9rtj2fwLQqg39rlvop78IcfOz/yyDRfqZxWLcMmUvK
s6atzsYKj+I5rwspM7qnCbstokCwEO2ioAaiSeT752MWz46vBSy8ZGg0CLXh
AXO+Da/BmPlOR6Ge4/nnJeRLJv7VqYzBYcVyT3Scl3fJJh8LocT1fJ8cLA/k
59ogtdNOoVmmTgDMYUoJWPcvYhZpAEi9sXrJI0J8UuNQxdv/iP6Urrl+pac6
vyIcP/7taJilhRdsAe0rHXWNtL9CFaBJeguGtDWWO48h+PzfL2bzH/ku/Yy7
/ZmFAvkdlZeen6jeeEQqDS/hcowllA2nnMF0GjvoJS7Tk+dws7L0X8BKD2/p
KaPH1N85jAjV/3zeD3qaxhIu1g3u3aWzyhyg2GEE5nrK+30v2Ob5g9sbiSLV
CJ2Zr+L4bem5wPuHgQI8S8toDgJhfYTwsqpjdjMo30svu7d4j0MPhYc3QlMQ
9KJ7pK9FSqQkhglpkzRwdd8bSJbogF0c9+qQoW/mvT8TdWVDU2PNJtkRpFEn
lTespX+XA+gxedZ2AEs60nMd/6OvqlOoiDui8yaAkukuONM2pCQJSsxuJNR9
VcOQNPQjvB25PHp2pmJV4rUYBjaJa1GddORezaaC2z7D2870aCjOKif+Osa+
p3DVfhZkk9k+OeU8/MwbPxmUeGDOL3yWHZNL52MsXdAxJfiJE4OYGJMSdAmr
DdAtG5GsEcNutDJt6w9nFBUBToJMNccvB7VwnTm+lQwappZsdph2/fHRUAH2
a7LBhbwSRzYIEvNFxAMWG68eFGMcWRqzDD+7xoev3LJhubW6/tbS1P3gFfgz
0lzMxZjZ81zizCbu/LYDe5CBvnTO5xXvUCLGfPfi8+IlWhQRzn3bIZaCrw/o
cp84w0u6x+ehK89/iNUWmgEoye0g/r+//FfdkcCowaTJsDSzKXbgmZ0WrbPv
Illf2EIC0SVYqd0vZ5i7JrIB1K7et+qiFRiR229WzeQjaiZ4Ie1bTvLFwAAD
6/SUFQOX7iAZIbbf3nCMWNuIl+wzrpeJy90E1paenRqdsySnySGwzsS22LTf
aFFnBRxA0vDokD+w8TQhRpiwpDuIt59hBx7xIDRD1CaltbU1NtX4eYluDdIy
DfN+Tk5XmoO4rEHpOSKbs6I4QnFmR1BT19/BBdejHVIIXgQApEj7EwpPtKt7
RPnYZrjeD/MzjgMDT2jKdfPk3irShTiT6XDyOol/MWwOqgFBKyh7I/WMynZz
Cs+7Poigpgj+18gjrxApzA4wpGUq/mmD505kPPXM08RU8qdH+UXw4a5TyLA2
UNx6P8nALn11/oODN93b27hW+2aIvClrROF9qvo2iaxzJvBVrhMs7MeRSIYC
c1LIm7slZw1N9KxbzcLf+iE7/E4LS7aZhW3OW7F+Iw3iu7PGjZ47UOOYovdh
eqb26irpBDAOloTwt6u5t8Bvj4qqUfGCycrLswJLSK384QZKwrqd8gBHJfPk
mH+6VF8/bXD+IY6+eXlPr/5DUICMWVj9sjbVykFwx5h7OPDTLN1/pZPbR/Tq
sprb/1xJvOLRnqlwMJRhxo1vVjlURAcpkgkiFwcDO4iDRijl2e0ROz4Tto9x
J3ZkR+9g7ANcMUNG8hpvHc7aMUqwpxi3t+Tg2bkqkSiZBxr9MKY4Br5b/pIg
MgLGgH8hdBSKbf7oDPKu1Y+1OpX3hqDMDAjFGOcg0vrcCEIrKaEIEygRtyPE
SGYSX3DA7JYEhO5Q72Cun9oXKHUFiFRrK7joPr+MkF8ea0PT2Aj2E2I/5Ebl
x4miIzzN2ZWr2cheev5KI41RgxyFyY0cuUs1FwVJaNgcC6rsaD/Am3V/I43R
zSJXnX5uesw8eLyDZNTkyCg7fZsKdNoriAkeWLqzNIsSoFxfVLD1aQTtPuTi
MzRbavNF36YsqQO5k2QgJXd+WI0qzj2L4Ng51n4fzxHWc2Qd7Icp8BAtaFWN
8gmjrF6w1TZ/ii8fyoEdOCnDjsoKub+AjIhDYZE/M2Pis8ua2SYPoUJux32b
hieCv+5rSJB2FVgnjDW9t90suPQ4f/qONR+WDCKZH4mOd+no315Dl9DtCh7/
A6oJOAl70694EQdDocsWV0AjJQsGYiwwOru/Q3ny1n1DYQK7pZ0I/A2p9B6B
jPwLTjZpcPJs6WWQX02Eg2L1Wm+7+lUVGcyKP3GMyWy+vyYyiJPQWQl+UGK5
8her5JU3W6mJVXGO6KrvQiUq9n+5ej46texer+Yp0DJb5tMx5iSgbSmejqZQ
ARituZ6plP8alqkdm43TiBIJOvl38wXbi+WcBaMy4ZfMvSscD3C9i2aROeu1
lvVnUdFiNCEIKhBdO+1+acxRHUv4UgNYD111q6eNVNgx36LfYk+ccZtDYBPZ
Ij/S7DL4vj6eBCzWjJC7rYh2GgIrv/TOxjeVRuqJCC3IfaoWmwMO+jGwzv6J
jPN07qADdw4IcHg0YN+uMCZKjt5RWCWN90CqHQbf97TW4BLNPPUbI92WAygy
WFNzBnvtcBE+QEiJ0/v4eLPxgGi2alTJngoLpNbt8yrT937lwpqOPkSjjQ9Z
GflY6HsMmmczoSMrHklHw3Ms0e9+VdfJE5uxFNs9fyM88wSChI7+62UWeFU9
+CxXYgrEehHyIvb3XZqDDPhW8uq53RQI/EbYjZJ/5I3Ajl6B5JQFtWpaaxDP
Vm3Ul6zTrT5G303aMLSkisPjigr/R0NPnZgop2dcyn157CIQPj30Rd7ZbR4C
nkUvMRMRPj0A2J4owx9YpJSu9TZBgxMN+9ReZOGdDMYauPogmA57yu8Br9/e
FHaldu49o6mVwDxWksqaocqFU1oXBsNVr8BtH6etoZvmlGp8wnXMWmc0CTt4
VoGoWEcpa98414lcaDy1i6yz5spbznIkOyWjO48gkN03iJkYWbLWxYmtB+TP
RYoRAPRgA7r60u2ItkG+1fE0209O0P78C8Ecq05vDFhkg5atK2RABE9n+wHo
JopQodofMLDEpksM0JdDHq+psDW3pldTbSbtPRl4nYbYHJ2+GIFdEZlAyWf4
PlW0QV/L5H18aoRjJAsSH7GBMbUUFvOQrknVpnjHUsOq+4jpsb31Sqt7ZTjd
Xwu5l0J+gaShFA24hbIptBQid1X9TPgyMIk77Nq3NlbY861Qzb9wX7byS5OS
p5wtSTYZuxsnpKSaRCnl5Bjx7wRtq603tV8QqINSzSXMemFVCTdYwmwpZb8w
1J3FEp3aC5Gm+D7LV/DK9D6TynCTcYh4eA5nzccUWcnsquxL+tF/YQ+7tJz+
89mnET7YqSTPhqazxS+v/BQL5LztvYGF4+9faNn8bIJrYLJFlnWeKQmY/tSw
Zxq1rNtzatzMmkAmnShy2uBXYYFSemimaSc4La7hFy+gZ4htQMfK7eCi8k2w
CXN9GjhatdEhYT3NxmEtAGxG9ynGY73V5rNY/re91/TCBUwr8gObCdoH2KA5
npjEkwLz02RCbZF0r6t9aP/5hfkWJkOYcnDCHlpBFN2KioKBWZ1abMwkU8cO
sh09pvOLMjHsXf9liHj7j9rHRJpYhAO/QgFRY1ylUXgs3yBiqB1OZStXhYRu
fsR12h5osm7RDa0XTTRzj+iWOoskJCy16wZhOBHp/pwiYSKyemoCx6zdNvjD
KWiaUZ2zWbJok5AUiBy9CoVRoX4ywP+x/5CcP/ypf3mk4Wggrqr/1GXkZ137
PO1gXrViEmAU5FAyT6OyxvNovgW1Vc7N69T/9gzzLBOP18VdyO2D2zUn4v6U
a0x0Qj34hiIxl5+CgBp+TKX5MbMPge8zsyVwjGnit+YEe5YCio3R1fI62uIw
og/oCXhSsSP4asc2SKeMEn1Xmv8p5pjH3fgJOdRzdHIBHYCsln7LKZ6y2mUJ
f9LwzEmjpYDvfxK7kHX0uvTS1d9+hS2WNAt260N9xcFfamRtFu9Fz5oB3vI6
CwF7mFu2hS/yGW9qSWuzHAbt6xifi4pYPZh3ok2+3LGsw5TeYYHeADggOMZL
iarTUx+CFdosiBea9PSuUQqcmdTewjUegRhMtP+sfVlIzYqMxopM/7J5N+cC
aEq/geH4GmQ5D29OSV189b98xHJXPBn21xPxaL19MQmw3bkEMlccdm/roL1h
aSWeFeEIjw4gC6RaTZFH6c+jPS0sgyq7DGXq/nVOt1I3oGwi6p/vcZOKGTNd
+nkwjvF2pt4PMi3eidddnMCf7EnliJfEPltb63DDuPOjq0KRt1aEJUKOtmls
8nANfRYKBmg/0P0vkBpD4o2S5pgU/DKaeVV+fd4sAnRqcFkuYfxyFePpxMuk
/NsfXLLMgO+iP3r/QRqGNSBs0jnhtVMp36FyRyB4+S1gdyY+F779H+UUR0em
gUl/MyZeh0kYfuJLpmdOUrye32Z88Hngl0AQ1FBIMCY3krNXoyz8u4rgMNFL
88THDr1U0exooeD3X1zjftWxavzXort5pCMKKUJbIh6lOnyljaRhWPTN7fYE
Vs/w6+eFSwzUkiMkrbXv7n8tyMfb0yTneFZmvEjgYhTdzyl61MPGrjWC1hAf
SeT7nitgpZdwmSpB1vlY4QH7RdMNrjOvvLFdq9e97y3807qNKkakDnp7wyKV
A+zdgkEmRaddWGZb6dNrFVSKToYILnRm3VRT2IArRwUgSIkbJJTGkeSvwIwi
WVaRCpk49LUfRXRjL2FM2x3uDWjw6CPrPSQxORTi/2kR4yTvfDUs9y88rSc3
SoExGQjzaC2NbsJtGLKpnObEPGVEITWToNU5Ul1wKzMJPgIUGxqTrvNiS6wS
MffSsTWAF+JZlxeD2Xc2M+hwCFPtDqcw9+Cu72W+xvhWYa3CxHXUm1mJ4wG0
Uf5+rOHBKFTa9XtbBvRnBswG3QqhqTuJWWPsdQCrhadSEYv7vwBeDWrJGJ76
7OXgkPSDSVHbeA9FxnwO4ZU2SdcYvnvW5WqCILFWsb9GmP2X2snyhish+qgZ
jmEycFB7E1rNNF3rYmXH96LKRzlXpYk35B5D0EmEW2JjQnV4dwDQViEi6Eah
crFfcikMwH1xqKQKndgrP/etw/jwwjf/yotl9zeZaH/+3CDG4yw7cbbZ5QZw
jpzG76KTzJTxCe1s6EBYvUcm1AELpZaOiPL6AF2H0Cu4jbCOjhUf9Iw6xXIJ
WqVhJlxzwZmUkIcYQdGHButLAR5HyYpye396PrJ/PsncPE0n7arVf/pFxMRJ
nZrhQjymCCxEtX7Tx1w4TFP06novpS1xyz+0xGKeZEWKqr9+EaIWr5bEIndr
Qczo1jtbNLDr0BXBnGjfvxV5/Btfj38SBs9wQ/4Qwl1T0ww4zJvZuESQ+yba
LMeNu02JjMT5FZ0zf0tTHh0beM7ie3cKz1ru4tcOcSw9XPVHLsJJRDFHh4Dm
+w2Mb19xQRpq5JJUFRBZNu+kRsn9LmObU2poSt5gt3Vlb2f1gwJNdYxPHZAH
5gmOWQ4OjHkEX57WDjAM1I6njHVYWaAtNFe7vwnie3e1Qo+e4r9pIXtaiBzo
y/Qo6wxBRTDUzT9MqBlQllECJY2t11Df7HCCV5wlk9E4D/dj7gULhxCnOXKb
cN3WfalkEcDhi2zzmAIDv6cGvYMPNnUl3iT0V1BOHFZnXYv6GAtW/rDUa4/Z
L3JEn2v1dDrbbkEgK9qEutkmwSRDQkZxVhBVMRVcKhUPFLlTK272swJf9BHF
V+UTFOjxSI9aTgr42y3v05BV7AmlbNg0jj8jusMytyBC/RWzBFq2GpXQiXeC
SPD7A/oROUZBxmo3pWB/tBMbfZSerb3HmFJST1qOlzP0szdvUn9FJvGhZvzX
w5v27TIuNQxU91GS7SWpDsbOHToMTsWiU/7TF8tIr6CID5NpyZcWz4BWq2Hh
eyIplyMvBHEkhRXNuQqCAEbnokbempLE1vlM5MsornmPlT10R6lihc3VFuiD
uswKofNp3zs3ed3pCmzTwnFZoq6kBeRC7grJ7PMeu+cVKKOgwDd95UUmQ+op
WLRkSKbAGRO2wJejbcRyeZE/0fpCq0TQCNGoHP68zS/AdcxlJ9chuRhcRoSj
nhLDS09izib5T001at/fsgH0mbAMWhIsLOn0p1mA+h1yYsWj29xqdckb4Rqx
N/dPqzxSfb+HtFsaWPvBrqHVaG+Z6fxUqzjhm4hxM4SFVeKw/bGS6fSCEBXW
APGTgpzNbwY2Ci5XmU2M5RIui5bHS/9EIspr8WY5VdR5O1R/93f+WMPrVA6F
yU65iBmjBM23dsQBL31LNP+ERr3KUNV6emNgcYzG+sNMJiDD+47RJpO0kVKl
Tj2923EgW8R/SIgLESKEVZ18EnIwFDDxku+Q02CuZ7uuZ2jOfOtIEsC/u7WI
lwpA95PYZe6t30Kaegs8ZSbvOj7wj+pwsI6iGj4WypETf/4EPoSa/T6cGmwi
gPV4SaR1zWmmyP3nmyhYAqmHgUjJA3JV2Sz1/46wkzV00AopIKL7xW/MCdAT
jlnhCI4oRQrg+RUGXpiKT0JgP7+L2nCJ2W/fYG8dAypCJC/1qNDgnZ684H2J
cafIrdsu9kiZyWmWGHCLsHXzk/0CiuxZ6VJMvchvJQzDKehX2xKYwVUrumDb
LNd8LfiZ9PKNLzjDUlgPR5JUNhmRz0//6zbjQua4J/kjnIx60vARwtKbHjid
oy5UVjYpRCjYyLO0mz0EDPvKKCSld7lDnbE7xswSmfSc2NClbZF1ei6pFXwn
o/a8s0szfww/0mfuguOfo9g+yvjM3UYEjJtsxDxk21Bm2ht0NghUpfN1tnwL
zTKJB17c/rLKHejXD1i5tPzaTWJjmbZ7UY6jzoL1bPf7na1ujqdYUY3QWOBS
Twxh9eTGgHHyxV9oqRs7BHx5eHgNBCq1Jt1OM8CCocFxKnx5uHbqYJHSLndo
zXJ7qfEKa9PL+BR19sdsl9a2aAWKKuI/YEc98EzR86mtAZauOu+LSX7bh73Y
MSoS2wAQ+1TDXwxSIcIaSKVS2dTmpHdzWPOnJLmvozCJxnfzVXgl311n077i
LNc4VBZXoShGI2kJ1JIIqAZo8lIc45bsVFAM8KERzxILFNXvK5p03J0JsPl+
8zJ3ibN41I+HUZwJ7dezU8jp+uNGYGfTDLsGomyfigJMMs2a5udcdj74Wrsf
zB7aGvk9U9jirvbMBbJIjYiyxTKBMyQA5t59mFj/BfQuS8/aZAY5MELGwJ2q
ZUiFRvGXwBvaLzpxlL73n9fuH2nB8WDzUDDbqJqjreYVBddzHwNf9I6F1+Gb
1bEUaerjdApoOmNj1PIbtPkrJHk8/bFwj1vv3uX6HInM+eqkOpcnQoAkU8/Z
3ZR8nZWUIsh08BlmuB5KpRR2mKD4sx4YOw7en07Kju7JsyMkjfwsEpKmjsFv
kC5Oh6bdcILnX50XAyJt24ha3m3uIPCgYGDDKnjE79CXfbLC2lRWPooX19UA
SegfJoF1D1LtY2z1u+HvrtMjMla7wJIcqQApC2ZsnTrywW8Ix9uejhd673xa
uvOYAwXIDD8QNM/dCgvkV+eKyfTavWB7Qao70nbSyjjgGy1BneHED9SN/jbi
/G85fxuG+rbvFqEpU6M2LvkRky7fAlCBf1A0JwvVvhrhEBwc8SwfU70UEeWK
G2jLrTlY0UkqqM+4iNne38d+1Lb2UkOrziJ0ifYVqzBChaq84vW1r0KMEtVm
jNevicHEOOBlvDaP3tIh1ALG1jseJnwaZFbnHwXhrjrPA4kC/phT0T3FyAzd
ZJ/btahtsTBdzPhZl9KFgA3HtopkEQqbaKmG5cW79LVG+JruQWBwtaBMgwEE
L3utPt/dyrt9l8rUOCmlgU15h87lVBJTApBsqSAjCzMRKXPnYWLeerUnAD+v
s6OQt0pfxXEQDVewBlcMlCjtV30rJJV6IQ0UBUe3yTpFG+MC2nFzUELKRWK1
uoA1Bzf4XrUGDzqJf2RGd7wnNxKa93Fg1IUkA3abQU09J8FQdRZpLAiLE1dc
WbTAcgsnl1W24ySCc7GLo9msjm2goQKQXcM1nyrZJWIzYvI3Z4MvoQC/mpFr
WeSlWE+/0Q5Cqyvn08l7ViF5zBFULPI1F0HV+nj4GisixpPryWI79GnIMzcG
ztWxGOf03FS8p2e12avHn3XYq4OyjDsQSw1cDM2jcCiAubL41W1uMsDvECpU
FOl61Y7ejnr6pYeevwFrfSWLCFjEJ5wBINs4aCvZK/ZtRX74ekB+5yXS1zUw
nmTSmarFI47ZlnWhb6b6X//jpXvrvqjduIRvDY+Mhz50vK3V8PWD7+RdqbXF
hIaAuJl0zIZlzv5Ep4Nld9kaz4Z/8+6kNZ0EtgmDgpnp9sSy6vTD7i+GIc8f
lYVYfG67eLVKh+Ny1rhBraLCTOzts/0NW93T7+37LVOgWWOEFVAHeGNdtIfF
UE/DxusWMzkMyEHhXkH00EmU74bgL4pgGuugNyVbONMGOpdXafEmmN/CWyFv
T/D5mM7wQlsusUvgzE98qF8LuwYbIs7JGYWjTXiSq2Tb4ZfaTHRtxMY0iX6D
rsPc+XovuQriksg4CFJUQdDFPWmy5TZRRUPVnt7HNbLm383u05htp2RcN/tH
7m8GT5kuGt/OGFiKFYq1VF+S/LmHLABuf2AH/Qn3P09mN0QO6TN+ZK/RY+P7
hNrK4i3OmMRfT8/6RRADWwbyJCBtyM1aNaW0lH11ZtVgvRQ6CqL/W1H+orYK
4SS9W0vFgXQDGt+IWRTUFwOD0jefPU0DFV+h6jXT+USxlo+dLmICsDvoRXMp
ZijiihC5XT4BTOVm8RpAueDy92CsxiE2ip/H69xEU9p4F8Q7rEY95hSJA7Tq
1HS6IrmHCOZE17E2dpjojfMQuxsRIBs9UQoDnUAJJCb/40xMA4jCWdAszePE
MNyqSwk2FjZ1YEviFs69CuKPFDQTvetN/AjFDoUJP+c1stLVh0binudxTVHL
pcEHGH46RilN51Gg5QHOLWb3QYEq2ZDHv97rstIJkh3Wf0qJ+kcRcnOHuh7r
dhNFO497Igl7ZwyhDPm+bWAigkVDeFcL9ji8oGLHMfDqxQ3631bCnYik5l4X
+YTMDygTJHT5def/5yW8shXC6rJitafgBUV5/EIYaCtJ1DpaU55YfN6DbKw7
idJ1ShdS6i9UlQGfZlZISFmo/X0KAFM7MbaN/HFDXtBzmiVepJU5unIIue6w
xPSd+V9Wouu9mQI/D52DGZr1nrk9VPqaLVp2wnKdN8JgE56uBW3xklsHWweb
sXrZx1WQc0JDO4d7XbbT/xnMMziDKjlZMyyzk+0Jyv4tdjVYdx4KdYGvfHTC
cMIhRT+y6IKnlAL3GlV2+jvCKCfmBI6RZ8Em9RI3DgTVOstq/DuPc38QiVpH
5nXSf5Qt0wLRpEMRjyYC883WFY7AF5DkaDKbqjmn07q8T4fLjDaPxbVHLU56
JQmZMnAVRVRFzFIlcaoqkZdXcG927/khbf+LZ4H+vM9munUIVUKDAoPgtz/f
GMxDfz1cgkw2QyvZ0fc0fysyS6DyYlUBTjQU1n9Nxcz3ThhdlbwUQAMAYQzQ
0q89MtbTt4WdVVRe5HpO9QbUfE4El3crrELAyFfWb+htjVhqQoa7ONOsjvxV
OWrdFlPq2VHpD9UoksF1cfViJ3fbEFuD1xqvZcoOsCFmqVaDm+zr34b3WCbk
U/cRRqpaAkljZ3zeLfy6evKghEu8lq9bGqihlxIOCJkncTEOOGPVbOsT/7QE
DpVp0k+Tt55f51UBLiecWjh4tnKIG3oicK6/3rN/wdMEbCRtYelFH9MG9qrt
ngBTOe3YNdY5XEOkJXAjRFp56z9PAn0ZkhPLfheWdZrq5N5PjhEHURyqR5YR
XacISYoaxLVYIyR015pejMX5EXiUGamKUptq43I3XAxquT4w52JnuZ0QrRhk
f+daNd5sCVDSbBnp2LISnznsADKEQNTygaZcIQktWp6wo0tMKBxfTfERgTFz
x2Xd80Wa4C8i5kUkXGOfG7y9+17bPb4fbKV11hvjZ6KfGqdIRlyH4ocrbfs7
yUg66FpFV8HnraP9E2afya+7h82/r6w4HXuP6dChnyM4x7PlbFotuhBvS/5p
SRFmykn/D31iwmhHhGLzQ9x7YdTMJFLowVcL8nP+dWVdL75MBlGEo619zDYM
L2Ti9RL93vqa1PECiD8xhU/UPLKezu07N/XH5We84KLgpo4Qn0WvqNXRxSNX
2yvjuZwqWRO47HItToDfD7IWW1/OrYq1Z9/hz6+j5qZtKTWtmk2KrW5Q9YdT
HvzYkMnE9rrKJNTAn0OQxQsCg0AZrlmGTvc6FWWRRBSEGF47bhBDbyFKKsv1
7ZFWMk0grEPkLHmBu7khHXVyIK7L3hBAaJVUvb489xxsPPtph13DY3heLMJL
i4BW/ej7cXWJTSN5hGT6U708Y2fSL5AXHmTILqw7rPhizWcJDYzIydKYXxla
shdrFeGL4iLWwUp1tuNw+ArXO1Tf9DXEdiAqDGm35JFYbQIrRaa33hIq4tlO
XM/NFULbcRWrn+VA0/XnHi0r5qF6ZgI4gJsYWC1sf09xi0oHrKHMl2ZRPOPK
jrucTcvG3bNP+2p0VXU2mhXo2dzgA6hfwQDzLLW20VxFvkjcEBRVJMspNBsb
Be7mqCPDvm0iPfkZFcabFILUIyLXmP96GzeVXAvl0hV/WBDogYK54OjzdV2m
uKpnwU+y6bTo45QrEVpePfmJS29BXlDZJhY9hp3nEV3rPat2N3nSzezYoVYq
1WS1lnDkD0wMJzm6I4lfV81/HQY6dVUaknTAwbbOx5/0uyQIUeINfQaurC1G
IeqOlkHprJ6y+qebGWh7EGexKnXY2zxNgkQSAUofzs7uLhicQWA48dmw9Zdr
77Mf2L8knDqq+UJzRDLe613XvH2hEGqzDoT3W8ldx32BGW31ofRYY/8Q8mNB
nu2YD9YyColFmYjbH+CX/HcYiFAw/imHCouMsljyIyrXOIzYQmRtFE2GIdul
JiIz5jj3g1E0bu17NMewE9WVPUZT02iMlht+WK6vzV9VlkuNXfdZ5UYlCVMh
qpJVBAXiPI/eJOMtaKU5POcHqKF6feWdALkZ9SqjgX9gHD7rPYYxjs4SXZGa
yaAng7QEYXi28CVDpIIXPDMH8WS015iEA31UvMUNicJVD/4/X1HMl152lLZK
fV/n0G3UMGXCupWHlBwec1d92ZJcIaWPZo2Xc2rE44IBBezQO/jzPQdSnvS8
2lYDWP3wbQ12qxF/H2Bk+BQibYOEbu3UO4v8hZuFOYnzpiO7EkKpZn2UKvrL
0hE4t3kKISEF+2iTV6V9vw8nHoNBxWfCJ2Ub7xvKCqTwpBJbvQ81HqPQKvcv
RxFApwDsypZdP/aGviZzqHkMkTReruoeE/gFWuJ/zyjK/kE1Go0gWxUwE37S
OFFCc3CCwKiF4oiOJLp6+edvu7sbW64j9jnSqx+5VYyEmmMqYmEJRRBRl4Wj
LI8C5pjXAnRwRoypPRa8GVVYhU3shMAp1OQP6orLLdnR98Ac5lVWSWXiwnGq
dwpgnL+uFmci974zr7gehPeO/r0FH5l3RbYnzYZQnlkBZ+Z1rU59ienx6lWB
FumnxjXCLQ+34bPYCZiEMTNKrNd+bV9awuImEsGXSzpIZx+2Yag9GIDJqNvC
GLWuyGB626/4+osmB8Ui8AKXBefkIfZBcSofQHO7DdOI4dC9haO2/DRmUJkn
Nn7p/ampF+0yryHJMUDGD9+tWUqY9Q78Ldx6+CplrdBHrXCFTC9QFQDLWplb
2fsQmDZYp1z4mj1jT9SIw/xAsf4YJKezNvmQ67rS220KdB08U8pttElPARJW
jaiA3dJXK9iPRePK4/WwnIsX5/pIKIb52IkwqQtxdAJYihvYt4aoo1yC+/6M
XahwkRzKpZRLOdXJB52r3Pvoevw8JrqKBHU1FywkHwhI5xHyoRdAu2PSFTZO
TAQChABSQ3/Yxl5a+C+E7q8YBoXHezhmBvV4ABZJqDZd+4eAWbDxsn9z8c65
CX8CFfY3EJFIdr+dyJWzpwLX4cqZzSObmT6ub6R71mcNwYMQc+am6ggcWa3q
wiyXxhNcXd1iOVCFk8+v1MbTFIJ83p2n5XRBRK8F26RuWxSG/ley6rc55oh8
DjXwWFm4qtBFYjd2AQcmC+JPdHgDZpUIe7WnxQhFGrjHWKxzlYPp9ZZWrSMR
TrgyHbjMLU/eSq9kyz4AI7YJ6ifI/L9grUEI2a3LWp2bwCFfCcEmc0oMuDFE
zfYmzK2f1gP6JOJq4vl5WUiwXC0kvReo2900rE9nrq2prfOsH6/LVvZpUnHC
S/go8JSnsGxM81ZvstAYkDOoaBrBGUsRszgrhNxV/R/jeBEFRfm8QGDwOzUa
fsBAQFto/NRKwPVZNUP1rjBPWrtJTqkysuC5kULQ6DCxFWEDlbJ4A+Ls1cZ4
VU9Q0FKe/kKgiRXtc8cdTKgYNbr39NSNYfHSzXYGytiXWA85HL+WO5t44KYF
ljjz9r+BhWGdtO4/psgnAp4ymtKoYbCi/V2KwauLFn48F+VdwcIl24VIXlCW
SSBqolMHAUR4oj4+/eFz8TAX8DHs3Dhcpub7bxnp2xWo991ZXfxxFGfyGhCA
OlwZ//upsO4m7rxrEdj1+8zAlQensrk53Myg46sbOa1NF9mswPunSWEfvNW6
KITACJrYvXDqm3YxXzB6zKmS04u5LF/oM2UnZofvHZYClhta3yWe6bmP1bhg
uojFi0/svOpQw2b+k2W9jkjNuX3fSAa+2UWCaLJD+goiFGCbUB3QneZWF9ba
+glTyWDkvqvS6vJ0eebIEJiBpm1VeMxN5WUCSdLQZGXrTV2RcmzDJGJH+Vzj
wtnhd4FrlYaArMZs5mKg6M/7KWvaGwOX3luKPT+lcB2/Jpap8baqQGlypXRg
oBifmzIj6iuff8oIhdQRafJpgmjAB3CP+rSewbWCB+j5/zki26wVEjXFx30/
i08jGZK0YLszJpBr/Bkgw76g3smDI2Uj9JVpuF1HUhPgCmJnLo3Egg8Myw3b
OLLVPyVeL768KYMp63dKmK6i7W4TD68lZ8D0jEdx8IqnL6b7X+xRj+6Gzx8y
vwAbQAsn3dIHPuh8SKd/s2DOx2XWKFez/NVZ4OvtzUEJ0ccoNnGj2XLuFGya
9kpAhih2cs6ksi+dZ0bB0tCAsKVrIB3By7H93fr20Qq8RzwR70Wh6YpDED0h
f8tWA3qTW4fZ0fD71mYdF+Rvvtt/bAolQos8GDyHOAeP99W9yroIOV9inXCS
FxWHowGT1O1EMrtoojx29hSwR+2H92AeHUEnjlTUTURNBT4kAqJ/h+Z1XF+c
SLMoXkQR22Cx+PpqWtSq9QIwnd6YmJEgahjJFGyd/es2+3JuEhFNo+HF/At4
xZWXiuQzu5BeHrmzcF0906/sYeGnPjW4hABSThnhCAPMxhVnDUT24BNA1Y/D
LDgEAyl85w0paRzAp8kFezFTRylSje1UbC+5tvqzYi8XOWSpFI4rNKK7myiW
V5xZJZy3QZlHQLKQ2nM6hU7p4J+YzrTzVMfgNqc6urOq0QaZTAgE+EbWqLtK
kZkEUXVO6BOWFr5284t1MJckxqNpGFnDIRQLqKk1bp//JAJx3vE5IBxKt14Y
sczdlNKzXE1ZtJPkczUOLZvQmjojfeUyt68bPW5jEWB+A0tN+CZqnNqCVN1D
oxXOrGDBlV2X15m6m9VwyWtWRZQQaSJ6QlnIWVS3xEnWIR/ybJtzuQMRuzoN
uFGq2wSAC/v60oTp05m88hgql9fD7KH9/L3zmLQSgQUYc2Tak0WRQr2bzbjF
wFojg86J0HEDNlscA1nHCk9iRZoP/1ye99Rgu3KwbLmf2wG31S8sRKjfM+so
PHEjM9tQgKULiL5j4iLaJfLzeOj7EFWM2gTUGQLg0fAm04mJnqFsEh+Kgyj3
j0TWUcs5dK7oMFJ0+1eFLxWrw364/YK3KxWk9xw2CRgUFfqIQ8ALRPA+AD6+
Z+pwQn6a/sBU8/uhKtX+BhJ7pZVvi8yyrCm1P4vYgguyNs/mgcoEQHgG3JMe
Z5+1lKyl+yBB6CnxiCsBEZm3jNjNdvU2yFEIXRejiRl+A8MYzeG6AeMYxx0c
roK9xjCIIx9heJ418voqUvog5q1TRRt5NJQosL6P2AqdPkFxQIWR1XTrhtHG
dr/e8wMEGIZ4R3wnY6Ouf0eNIqtiMf0U1oaiVQPOpbIXAPq9hsPTB8OWtibk
VgAzqPnhF5lvUd6jPP4zeZSbu+FwrKGBYOaGGTdCKN2PRGbxGBSdXXM7zkf6
Pse20xpuBzwCM4s6ldomMNr35ZCBpxkkM9oxYHtVB5gmy4UdLxiwBjRqf8gU
FKEOmwTGdS+jb1G/Oms5//bCq3/v0rgIRmXlzMaJozQGkQtPyI5uyVtYcBwq
Nh8I26hf6811aexG4hfMXjdI8QFZRzWpeGqfaSk7YnGYCWGfKCYP2MGQot/C
oVA4iEPDbresOvk8q4FZpMeomSpWqOz5/fkwVoziI+OaS/4LgcJbF1ksbMtN
3HyIYHBM552ojwPy3fIfcJ4fW4HOvmgDklldS8zLrWYg28YCAMdJnSzKyy00
+uKWCiWjy2ruaMNLfN0HmxnYVG/XTYHswE4C07G7JzUeGRezXgpCdvSpe7SM
mJtZ2LcEHWuX2mjzji27IBYFXh1Wj+jxyTmsBJpfSIDSwADGUITBlLplTG+J
4enDsJC9Tld7QelTxjcE+r55+r5AJOLF6h1H1nX43ACpO7E2kwNU/SYNjy+B
i/WmFG/SHAeHCZk0Dz2HRE4ztgIhW3GpHp4UHqhyrs+pJXS/UXqvh9HNk84F
uIwQX4T+LIyD98MXdtaE/40qehcVyEVQexvQeY4gJ90hWBcymQgnh46LziYs
fc3flAv0k+jaXkrWgl/OCOnwaozlRMuT+Mcw9UWrydTtXgAL0wFKuhZ+QMlv
hjGXHXPK12TLJp/T1Ww6n0KMd1Zwyz+oPbEalobf1/ewj/VYPoa+bOl2D8x9
oMcvqoFFN/ygyzuLMc5yQBja8KDoswke8i/XO5y/evCkYqV1Wumeru7nB+B/
fCOO5ATiD9pupEtWob8qg1iJG3sOw4BbA02LahIrQfmz8STxvoVYUggxPCfK
TKm/f63kpjuoRvJ2wYp4RsoEs4ghK74TpOj0orcpf9kyK6d9BGNJMU9g9KyC
S4qu27PVVq/P+VMV/e1ODEEkfORhJ27FD3cKr+dRhlCauHLs8wM/2g1CqGCR
uSTXQ/m4gp73h16/nMFTlXStfE3ZCtmAfXpe5HKPk5+ze1jW9K14zfRB71fo
+6aRjqwHwXvE5CyaTrswGDtwYjnWNg0egMRTEN2bza9s5Ief6DgoRsPgoeKP
c23jrX2CP1Wdhv1zd0KPam+a0GD29qvbKGxQ336FX2286aWjQB2AjHQSthB9
AUZPCPtJ9z0b4LbFcOl5jcoVJZyOUGmZlDVXdq9rqXB8dqqqQRykj86zaeC7
PdGIGgGt1uSjCDxar43vDN/C+r9uP9bmw6rtfW7XyW4Go30ZCHHl1DkYSwwQ
GONJHETA1HTBh1ovVJBrHhNWXW2nY9mvDa4R0DWMyCvj/oVoHLEHkEON6551
GYjbC0vAzBAXNNlxaQUE9D7D91W09GO/1lJoQMxjV6vIMSM0qBQ/i87rzQrU
xbUBBryxgIGzPD5Slt8uKj/z5Suj2SkuiopGCmtusIkjfxesPfNLxEpD3BtD
XjIwIp/qT2+mbg+lmrE+Gpjb9yiBv2nfyFoqEIPtB7chkiTw25IysmRBa00j
NY7BnXxvXjEODNtKC6KUpNfAvUXceayxgBJfNfH0w7H9H7Ut1Z5c1cXQCBFC
KUxVNif9cf0IUsDibXR8a1kJZylTHTbnwn/ozxZoGM7TRscLiQOfuHEibKiq
MJ0h74Lv9Td237NQ6fMPFTjwL3IqXNO2Y69v6qRd6lUcp4jD0br8hW2o8a+q
xPSF9LRuj4Q4hCBUrlJ7tozB9Rdod75qiR7hqROJ6Qe7pfACN2qs/rHeWfI5
JYxlicl/HWo+qz7rmOw5fMY1MACuRjT+KUPQ6UnNd1D4XcC9jGFPLhxazJCq
R+5Khu9rK9PEUzRTTWjKodcHNXKMsAHbYwu1yS0VUYdElGPJjszevbgmihAG
DpJK5IICVEGlhBnkyNj6sT+Q9tSo8914p8bcMXaUiJn7ZQ/gBfHmXDAPSSrq
TvKlOfpG/ysSbw2v+qJmQ5l6GZHMDsTI4ipt+3QUGplHETQI4042dh/O5Txd
qp/Ri2mEp0uoJg6ZELqLvZJ9pgXJ+P+pNlVkZMRKnuNnsPc3wfgYm4Mok7YL
cVF2mHdUe7YZFYycGLT1wHuGWX5jEKIAYgAJMe7KzPyOw5GhI0oVtrQT4s+W
+mBXuNTxWWqULtUTAMXvle+yAopDD8JBdh9QnaR6u/pWss5OFzbBpxRr8pwE
Ba6pLILMd8u/D4G7dlJTpn3K4MGppq2fnJ6EAw7S+oueg6o2pePJYZ7pqSwn
CY2/y3uUyC4TtjGzG9RsO7T2yeHXDMGxgZNRbcLVn9TA9NYY7AROhN9umhdt
+E/AnCDWgDan7tcmvPRusf/c/TOVQ4tkiNT/EgpkgH7UFJ8uBDZDw8ydb2jK
hhn0hwDmE1MJmixtZRJgz+kuPIZVepLaom1g6wxxBqTkVpik+LIEFsK6avPN
PCC7StwS8rmGDJDw4BkrocJ2KL/LUnrCWTDGiFlbr2VZP59eP9MjszQ0ARR/
X0g/3oLTCYkl0mqhgC56MzGU6O2Pd0kSD3aRdeK1Ali5/yDMzJkpteG8gCkM
BvJPHpYntKftuQG1QXxMSIPv5RUOih1ZHsXnTpwAUgb1lUQY/lnK8B50AnQc
CUbSYuUHZw+rRHW/4tm5LCqLqoZMgNuIZ7pY12upGDtyF/Zh1iyngcmtBw6m
6PE8oL618i6cEIeJ6Uj1Swe+59QCmTNQyw1nYirAeDK04x2jNvtWu2esWKP9
EKw6UUio+1uPBEuoFycs72W17w2G/Kkga3lbB1tJFfUp2T04twJlhtkmrSoC
3KMFKQPxtdrKHk5FPdlCc1SS1DlqcsOvjZEYgl6tuzBhV7EuCiiMpbyqWAqa
UqrTuhK0LF5qqIljt91JNb/dxfunh0mjI0Kn3iXAzFnA8jDA1VmUIg9lkF9K
21ps8WX/PZBXZXvJ2J+suV4XbG6L5DOb3+SkO/zEMUheIb0NKqGK2SmXePh6
VxU3MtSpfNqCxSfwFaFb9MtP7MQ2OAG2G8VPa0S0GuCSCGssZ149NmUZKb/Q
E1kF57I+NVh2+jG/Uwx5h243NamdQWeEgpeUrOWUfFK+E7DhkDN3fsSteyFk
28PWGIOoNbtnjxf9rAQ0iyn+W9ybwec1CmvnPfjmpg9tDC7BVXtEbrPRSeRT
ndb/K7I4FQKOMLj5WOei3j4OrPRcrwEjcMR8ehwPdLk43NRqQX57ykXBWpZV
0hiB6/cQgf+/9/8+QfVCmnOz+zGriLfClBVRpBChDRBjgrtbxpbE1sUyOvkm
UNmDQOffDiasDyOLuJwIf631aZZLPeQ+LtMJichTkjKvJ4dDpYqc/15d6FdP
84TKjXosYJ9Jp5z3Y99VX/XWvITADHxPLqPJFwFSFKHMQIfHeaWgUSUKO9n7
CqiQzre49+kHU80L8N5UuBx6FdySlH7LXBph7LwaPIgIKBSDhEBsvlX9k84U
+2TK2wZThKTahiZ0wW27gFYXbBXgBGDdQQNL+2A6BVSsmh9JIhwljOLG+BR1
SCi9hwdYNmplkoNiX7y0Ol/LHpPCAwnaYl0s1wmcsh7aYoLsElRnfTFtYUQN
N4zHdFX+P3XkCTZbICTtFZ6Mm7bGTOczWTyTNKWEiFRzHQewiUKa52wPU1rF
kVfrRr3qAuCp3svE8+9iXHpp8oztR4d6M8cuVnf76dIoxlUGUrpi/iwZ3bB+
QYuYLN9W6LOwn1j4kzMZXS8OpLq/P8cGkIv0WR9/3SeTuAfjTE8U+5AKuD/D
N+2c+dYkEen6jT7x9swO6P+URz+FX0398D3XIE0lMDFvBJ38X6bneTbQAKEU
yLe5md9Bo8+4Pzowbux/RYHirPX8Fh2JbasrX7vorLsJfTIFUI1fP5Sw3D4l
tpU8ssMwpPmEHN07QvCk2n5DXEM9owELtAQnF3/IwFIaS3YnateHjUZy/e7a
K/tP6PAuudzTgDiSKa4HTaFBEnYjNJj2sy8IUuZ52azGlsyRwTeoMRlqxjIO
t99u0UKSSLwLKlXzFVkF77IgJ1KErNxRIfble5qyLP03VeUUMnLt2IR8QAvd
Vdoro+d0neGOu/Xo0NOXBEYY3Zw3a/cxDvE169wQUS2NufDuw4vcAkwW3np3
UdAtkD0N1cdVtjgafVGffuNA1JL1jePq/El+0eX0sFjKDKykFx2K2z+KZvlq
pp+5+QFYValgFhcbl5N9G+oetnuJjlkjPayZdIJI2LFPxyRMBTuC9e3mAiQy
XYNZW8VYI1WbsdienOQHkhaX0raADGSmv8ZRRTfHAPA2fIiO2gOHAmtc5L1d
OlErNdqeNwVig4Zwz8LDSegSf3HmXQ9Psn4U+ZjQTEqQqnVSs/a+1BtDe23M
0IgMIjCq2+jCAPOIvoZEwlaVgGaoIQ2BczVAzz+v4zBVO4l0k1xZNZKTrSDq
IFPsX6Z/N9QNpm9T4eII1o5V0QYN+44u4+WKx2XJDFAeYP71Z/xCnnztvB7t
nvIAOBGh3zkUrsv3OqwQQLeTdqde/RqE8iQHM1oIb6UWSH3CI7UaWbXd/yhs
3PIolgoXrsWHBJyH/2IMo66WgQ1lUViNiyk20TxASQ/lp6LeYv7q6voSwerI
AznzwDaJs84h4zR43sFOoemo+MWfCS2jgukfI7s77FiTC5MFLXy+ijYVM2ZD
fTPyQhHE/E6/DwFD2H8XoIvnW0uyjKEdAPbgQ25K1YOEgyvgVd03lzOr5Yxk
NpqTvBJoFvLFgp71ZDfF5/SAFos4SZ/GN7X4wb7vBGD+Bau77Ln0UTAakdTK
3KE+9fMyeZUNuSaAdz8rAPNt+spA4PeYr0Vn6aMjnXl7NmOiPfhJM9ENIFC7
/waS1jDGEbsohDV4jpsinEO8tgqdvuub4IgYwJEOdegQHGza6WA7GoqUnPYQ
lFSSpMHkNMF52WQ4BLlZzO2GBgc+WFC8YQw91fI+v2H6B1+qBMS/K4NRuQ43
JDqdCY0kfFS3OVcY9Dg+rwHJKauIDcSE0nAOIafOhwocpjln3atvSwJ3Yc4T
0js0URq4YEi2CmgLoDIoQNAWqWs1FnhDvdHhgq/+EKxXlFjcZU3ujLcvnDVI
rxSCgOmwmzXcqM9n5tf9KtkAFgkcDhgElXzA+iJyyLSASKhe9BSLIdUDLUdk
GL66rL5d/yIuDs+N8Hmn/uxD8LKRFBtl3Uc/Yeu1trYHcsLGpYbdfUIvB251
I1rj/kJ6HB8ZNjjpXt8tqpVDIz3YNGSY4ODvHw+Q8WQBGYjfycGY91TJVB9I
enuEuLclhe1Z4GuT8O+GB1bpVWmmjvgB+vWGvqFrYSDOQc1jhiZBPtI3pJDL
ECICrXLy3wbY4BMlRbRlWxqU2Rw/+BuRX1TQ/hNgC1ToN6mFPF0DvJlQt68K
R16F8axzopHoukE57nm/0Y3A70unSTPxk6DQFjomDtMW40ZCEwKXHAza3EpB
XKlOkE3VWSYP6xfK0cUKHx5lhaI/vJMYMaVS93u9coP2ccLIuHLtJa3idpPY
C46HC+5iD3RKpjytdjjOFVZamtAZDBCo/PoNIrbvosPz3Tv858bcI8J41/qD
9+Uyy1a+yXd3XLwZwk/VrieSpmfpKIoTib9oU4KUN8oPTRqETu/nw6daJTdM
DMbdq7B3bDd/VREtIo7tkYATyhAqrz9TsN967d0gRCM03f1W/5XE+9O63pWX
BXRuuYxZKgRPcNtUWoogby3TB2wusYaapcdZC+ChrVQDxK1m1dWygDwZ8x+5
s8A0SJABm2F3P2bLd/N93U5illq1fOgiVN0x3b5mbP/ng5lxhQs/vyc6bVH0
u7c8ArMSGRuAW3Sx/btohf3iAxtszWBKyYGKtMAv9hJPM9AsiQGK5t+C2lWU
xmQv8Fw85BKZmq7BDtEZqkcrchfG1yvzjf8P4DrkXpsvOZrSM5pFXtXHL3jP
4RrkcV72d5hK/S6rfAU8B7/sm1HWku+HXBnshd+7GjyAEgqjgQM44oUaW4NQ
sGw4FLsmdlu7XHRjuEKveDWHxvD/Qrafrh5z381qvv133EqujFYwRxDcdvwj
yple3wGQquYpNCPzjaPHmFQfBSVaHVDIbprmc4hB/Uc9ii8ei07GAhsD3oQo
JZ5R35Oxc8JiWRzn35Pc+S8CsXok+kH2P0q4lw6U53LFtdJySCOzvg/5Oa0c
e9yEVvP1knKEj19C7wq4OO+xFPuIKdQwHbOfj75YSVknSwTme455mj8UOP8Z
dtG8mkN9xlLgcwHpHcwLxXi1JLDmKA53va2/wD/7RB2TG3CFRdJwYdSUbrMx
xl4LyF28knnixz1o8XMEpOYUW0qZxVMfSHzik0PklvVcLzUFdCAuMQVK71Gb
1GkPEyDJg1a6iK8birrZ2teZNdZw+DXrkMoiwqpcBOxCGbjDltQOLbaykjhZ
VqyY96CjVcqn+d2soXEFXfZ8dfXdEhobXcivCJeEi4Qusn9UwzVgTljHAv5m
YTuuQPiiSU8OsD3XuTTSs5Sivp5GRXcRd+Hdy8j7vrgfAUyIeemwnrv2+P1V
7c78U+hy9eByu0Gjpcn7ILD904jasGQ4KNs3n8zVrKUeuv67OsDItsIFGM+/
dOQtN1dCfAKIqSfd+zowFGv94W72n3ZqJluL/dBqOx2/aHdDeWsTWZfi/j0Q
OniH0pGMyL6yFRwXzY1YOGcwgftNuWUSItAshK97XhieqmUkALxsnJyH++tS
l+Dsy7hHiEXho6AZ10g56s/POVcOPeVywDx4maEUIpBzIuLErzQrgWIuVs41
YHsnGzl8UA1W6yA0iBg2G1wOmVkUYiXuxYBTBfNTYEIFhgAVBX5htfePRhMR
APMKogxzUfURbTupdNk9rzyNX9O9OTgVuTaHvVqXCVdxxubEt0pwDFPpq7mE
v3fP/wfNVv4qhASWkrbhug+GFOMj54A9jpWhqYZbiKXvIQ1lLsh8JcBWMChA
edAJiY1EVFqnFFcE/AgKlqZACOr/BxIMzuddXhj2f4XMHnO/8oih9r8YQKMX
sexzm1ySIE+mUnAn7ryx1MGFKrcO6GT5oIDaePQ7cIpyOQhQsxgENe/Mp3sQ
JuEa4FRU4rRV4QkweISZfjCu1QZqUBy5XC7jD0SMEb1CWq7DWGrCDyDLSSLk
Ac/ZavJtPrIubYKdei9znl3cJJIKmjH0vz7UDnARNtNJ0XAMyxGVA+w6FVr7
N/aDLmnh3bl000GYRv5cjReS1Em8r6lBu9MPXijXTFsfI13+DPQdCxtR53zk
EgJXgCYTe0nUMnIM1ODINCVjk/FhHQUpjv+ciShA2PFA9/zQDkzoraaPGp73
vGV+qsaJ3gvLGAOQwE94mqoMwMyc0FahzP1JtfbbtPt+k40e88nnhBRkMu2k
xKqmJE6FImQCroiWKCDi9MxVx3dEU8REzSRm4L3L0y1+FczfpNVNZ+VQK2bg
TnEJdfN7McnnlYaKSyJMk/esiqpBeLdbx8Bz8SfdVAVDbJd9d8ea9LeYu8bg
qMv8KqGLJsboj9RX+Domo+k32NRkG57qa7Db6vs6BSh4/kHCFYUeoABy36Eh
ikBWoMG2uYpQ+2nr/MlqW8NIaqRe7y8BVPWRkaPevBsJ5Px8GovgPJ/ZdXZ2
AeY4AQSd07WJFj202OIsZB6n4LXBXzMmORycMHZaESboV8Ky6SqMBsh41a0v
rO6Cm00HqGCNaO/+38YKIHy1eCP0bcxi6HZrcxXpOvY8xFkwtGU/DhrNZ+rL
Neiy1y5AOY08jTwdA+bD9MZ5t65QhcfSJHdkZx2vXARNlxSMp7LJRnm2/keZ
4TkL0QMNSo//ninQ87jvrAnnogzNtfzZovTfx9rm3F+6CuzoYbsyNRZ7PZKR
r2zUUSTofhlSrWyVP4yu4TLQBEJJ0jp+iW9bpEjXlxKK8pV2ERQf6yFixQR7
KNS1PjMaIAZAQuNkM3muWK+vnCSJD/hIUztHdO837rzF5ubrtO8p3y70l9Mj
L/qiXjNpCsWO6guHH0XHndWCqFqNPTZKin5x7FwV5UaYnog1/DpXLLzF82Sv
BzNPwfwP79CYby5sLbB7EyWGBu92RGZ2tISqP/DaD+P1DJRgERFfe001O8U5
lj2xbSvRM07eFGOPxOjn6IEp51oj+TEJKBBlrxyEDReAlQ+m7u9m1quepxeu
i/sI/zM0BjHC7HVrqiKV/l6uroClBim+qv3e2/j6e8s68fGqk/5MH1I5EaZ4
Rp6MWY9SP63ZLRBf79T5ENtSMPJ9t8SXtUr8SKB3RtmArAOXjaktLeE61Jxk
CmwfjFEm5Kd8JWAn5sNjh/MziDxvdZGN5F1n/qKK2nWSPjECP4Wj9uUi4Woo
uVpVvdSKephu8oIyo1AV2gI/IcuCPu8njWHhCCINyfK0wYjCDH3dtH8vowFm
UqkI6+F++SbGyGKEG4ZqKe3eAA4xXSIDcjEYGenRop/BKv2nxE8av+2wTYsj
RUHLc9kxDghZ5XPCBRiFzaaKEp0Q89V2hEGHWtOrG7uLr4ekH28uQ0T2iHO2
TXFopWV6mRgzQTTnPbHszb8CJTEB+WD7EewGNsOZSBUzhdDBfzfaZEnGhdpt
b682jqKvc03nwZ37VEb2CZmAbe2LaQLmjJbVjrKyQNxR9AnYEUVQDDKwgsFV
ycBE2j5v3e5LFIpbcvEYLVLTWq1WPuAXOYT5z4i1BJVQuuUEqAiEYyzHbn+m
8poSrCZUkZzRXUvKXSo/iA0iXB7AqP/CQawAd8K7r0J0AJFzLP3Cf0c58AYK
mr9TWbIohKJf3TVYoljaz7hX+NlhNINsYOOnQGeOUrbgt89VJqEypd6CB1ps
5DwnQkKbWbl3wQZdkTTeFnNgbM6LBcdjuY3kn3Smfp/IyfbSnaCs9WjtsrrU
iXjd3vZEoxCGGvOce+KZOepQoZ/ANYk1awQ7j6p2lUJnLjGHEN50IcWG0iUl
+jaXu9lEJdwAp3RsaDp5mmgWzVvz3vknUxYechX/fUxxKMN1TtnZTYBN9Mf/
XO9JdHYpujzn8NU3CSppRVnJsEeJxEqmOK5qago+2GiVGJ+qjrGzHOQq1Rjn
1mR3nN2EJeLnZ56A/43DMLDF4rUN2+sIVVLv54D3HDN/zO4G+3DkjtOoI226
GUdokBCifrrZcRdNLwV76n7vTwJn5kY/1QAuHKxUEWcBRishKzcgGrkxNeS+
kHzD5ffgyVWwvaWoc2U5s9rTWzrYZGiO6hKDDSTJt1evLkjT9WmS7hj1bcIJ
lA7zOO/8odtZkv99b82260nojMUnsc9WFrGuUrcMqeVKNyONUeixtwI82RkV
eP+Q0Snf5668m81yLeQLZLWQx0DxALRQZEmqTgfqEuVuntJVbxwTXtYo4Szw
0133QSJeYlYHc7B2U+7Yk7VYJsu15+x64g9zhZppdJqac5R1SVXsC1nay6rb
e8zsM6yU176LIfwRIaWNZfipXPmdXdaG7LI7WHH6UlafXPmD2Kjzz51KVj1b
mT0C/t8NCNpVUUtBuovU/MhtqgRvNdPIi+3HuRryYndpIyQRPQ1QA4vqo5lb
Qv8bmrfMWACAQOSSXtHjtY0nBDwlEklBWym+HJ+6zSGZwrPg3xmNTSoronZS
hAMmYflDsg+RFPi68ZJcWdYIRxf9SSqHWwhua13Dw01bPDkMcofEsgoR9oBm
Wr20CkM/B4wIEGfAB7uXzbTdV2rnsilzMl86u2A4x3zqPZxR+ikLBBa017hR
q/7wm2N2TSQx44vUlTBds0IpC7dS76itKJ+FrmmbljDGlnWlLpKDP1Td5wXU
egLWjhI6l447UTL56gZwFEyy/2AHrT9tQoUM9q1sZ8v9PbwfgSYQdF6fNP12
ag2NPCuNRFPO1GiSUmLd34nUXcXbnGlAVqxAvJ2H5T/ZExzF0B23rb7BHSV+
vTeJElsqT2JiP1Ax1j1vGs4o3O00pUkUDV6gOBZX7Wde7LM4aIoOvpGO0Ied
1oYLwOUztq/t4+v7GHYPOw0MuEEzbeFbhPnQsKPrloSThEPr1+kxLkRd6fac
beW77BqNbH9RybHliULXPn48f3r6Ib3AZB3B/3MO8Hg9Hlt4cafy3gziZ7O7
iFbgIliXGAZKafdYeUCpiYYJ4XwsDBxIgk+UhbOqW8OTeAIIkJkaB42tl8MD
An5SM2xDsR6e5taB/euaq6a1ldPKOjXgiZYOz6cNWkWdzmHL6uCNTp6S2eVE
0qPtt4h2Dy5Jm79VqHkggl2l7rq5BFGdoIalW8nbcBqOJvpDjnaRZ5rPbXpD
SI31NXcOXxCBoU7DMySyuZfj7zVoEyYKuywZom5EEex0jMNl+GOb+QyQ3tsd
g4OZ4Ol2ECEdN2wLZWatvyX/e1YLG35I05XJOnnsChjManIu43oCUOIISHA8
sokivEACA6PbFchPZGS110PneBL/aHvIHZWlsJ8oNbCQrwMnKWKtDg3ph0L0
MBLeoEmRJT6TZvd7I33ytCfM81KYrIH5w8DGn2U+bsBAmttORkZNBgdah2DK
7PhCLbIfByAcqDX4tEK9c1rqaEBJkLJmAry6to05whBBsC8daEXFon5k1HrW
Xk8vbOVCWXa6yTJ439NzcoJcX42cGsK8nb10K8pLBneUw5ymcnLN53kxieuF
a3HIixN9fWx6r+WxfPu9PaD+Gkcj1jprXPCjPjvMydyJ0yZL1zP2o2Ehlp5W
k8XuclC7uCf466GrX1qi/Ed/uR1/zckac6LlIba2bkpaXNqf9J+rLbjmTLmp
ILhmmucYm85S0N0w9dpQ7U8tm/cyisHrpRHR+V5COxHNgumGIx4RczSASsu0
8W1JfkT6Thosdqr3XYGGzC1Ym319n7m0w9J2x7E+BUwd1fa+2Zh9kYc/MpPj
Ge53cwjac0VDh7i3BNUooASmVX72Y0xCP8TpKsrroGwiT9iwl+MZ+z0cCsYC
BV22UVyxCld+yzBIuWjxAymup8S1aS3vruar1jQR6+ON+lTxF8EsU6GvxLRr
00plk3wTEGUg/lSpXR9f9sfxXVrrAz03aNfk2lyIfhGNTlj/s37ja2DeomGV
4JjltabHJ/fLZ4j+CgzwPoQSJjm/qyqQBJLfkkwXFmPJ9hEkg4ZAk8cJua6U
WQ+QTIHAz7RMdfeqnKlS+3+wKoEYJqs4aIlHm3m7Zaug7zWGK1/k8rVwBLSP
zc/R5zEL5HmNZlkORx0V52EbcvuaklRko80r2Os0DbuWXtGc67Ksv3z0vxtt
rpg5ABCmAqWwEgWJTFruqMYZo+ZC6mRqY8+ZPs6yaPmNTM7HQZWTvpjUZ30L
W1ahjUrJmXEA+d7wDpCZbizIj0Nb2E2yX6T5yNDof4Rcx2IbLywzAyK3aXj5
nGufw0HeyoJGWgJKZbgJTnBdV7C91yl0JFkJ4D9oWSYOzFfrG8Cly4fGmMEe
QJ9xsVF8T7E8qN+YKkm/fJL900WdtnGUqjgsd1z+PnjAbVTX+iVA21Kjv0hf
vaZ/6wPQyzfQNbsWfmDkGDFAvFt0YLRiR7ZhqmxLjwGxceAbGpS0Z+39FmB7
aJGgXygNJ4Poew7FixI2mtS+nFkO9JI4OzZzHalaRBgfeAwFB4kjiavZLVO3
Uy7N6LbxltFveB5IkQwpZkU8Ym5JCfzmc0O6sz8U/xMC7ERXRs1aUs4rTO5N
yYnKzRAkvRc1djZv7Faa2GAwmib0bdeLMfUUJn6QnmcEVrZ8JPYRiRKwxHcE
TEHFjQzw4kM8w51cdgBFWpZ32h8233B7ajN2bXnfXU4o9erifiudEjXvF0eD
a2icrdW7KVBzPH42WF4Jngfne8oPSfVQW7f70aOJLpERkArtOS8Z51Arspdq
dEpFBeUU6cABJ0MCzyZFtesQ8CiWYMNJhcyRlylVc3MRQ9XdgmfJgXqMZLrc
8F3IWDnCCsTQSKzpiX2J0y0umk+Fjk5MauS6ta3+nR6fPYS1E8E+dTVS+opm
0bWLrqgwIKR2k7/WKaM+GWu7k/IvPhdecSUkehXhih+RCwXN8GwuzBZSV5Vb
Ssr1LSk/O/geqEhdYi+a7sVuNTzM+DTz/C3lWIibTyYpyzk5UC7lpOU+0Coa
CrHXdgYieOT0JMShmSTR0urE7gDa0s95NdR45iZWE2mMBFs8hqINlCTSrLK7
KGMiXeIzQ8Oy/KaGhFJeT521QuaabF9Y61/DxAseYkUszn5W7nNCvQTkKAzC
p1feX6SPPDKhKoZQKq9GCzSSSu7aoN00djVb1BoJdwJKw45gzcAZrChkn/bg
Dw8F8LTggUT2HNZzA4lDxDOiZGTZrxpfovXSoccVOMso07qlffjfr0UXsB7E
QaYq4irWhcm9pqttB4v6PkhItX5BvdVcB0HomIqzOjuE24IuyxOZ95IbSgAX
utqKt7zX+2Z8Up8WJRqcl48J+EgRuAPdzwyvKm9ibmeCiu53zaVvwyhxSFpb
4U3P9IqsY2jHT8NyS60uDBcnJSe4/0SFN/WYWUBw3IebPHdHUcxRrPLPXKrW
mT0L18s2vNnF6b0DScNJzm+sM4ULS4gBASansCUW4bQ+I42dki89x0J2w69P
/+Wg9i9WIrpmUaWrkmiZ0aRGlPKg0+6MeR8fAof/f+yZJliR6efgjXXJDB2i
k6a2XFokSugYty7Aqb24LbPAALR46tJidppks0if/X3gcPt7JXvN+GWetjrn
N75VKYKR9gjUb0ALtlRmfMmXkrlL0rSpMutwZGX/utq+bbZmMhswJc6qxJS1
lH0c+Ad+W8EvPcrI7GPwoYuXGmoNbmKU7yxz4isqxiiTtPGiS7C1vhYgo/vt
H7O8+3C+MAsu0oleOwIFfYqy0dDWTvCQo6mUWPeUGbzZfUfbIUHYBeq0epVW
G8W+1TKcSWbSq/I/GYsNAFeJmjFDjDPqTIYCpRhLWJPyIuJ+oIYA7DQRLGcO
BxcWqumh7gLJLjWZf1cW5z0qsu9Bg3tb8Ikb4u3NVB4oh/PFR4zUtF4veYQ4
vej635VRN1Sn2quNuLQEu4EYknCrhIXdbq/4sZrX2HS8hvQTJCuKzm79W7vE
pWMSIURl5nez3NflJbANwIT4ul6aUs2nIBrYpOIKQm5F+ekPTfjOLXzV7Y91
bRHdKlNh5nT0hYPR8Zkb7l7VWkukcbx66c3MUSaDaCe+fD7mA0ODQfMaVV/J
cYiHAuQkBH89UFX8wXMoiENGCUvjHa5zIc7qO/Qkq07oErTb9O+sn6ao9idt
/JRCFLSPsGut8ZbF3LoLICf7ImM5wEGTbbLT+gv6ejJ7Q+uX3fZD9mfhaRti
nM2Mcc1KcZVa8e5Se3ks/BssqmzINHEISjyzOUWdaJRFstlYYZ5OZvgD8jYg
B9xiV47TlrJ6ZSLiYeAcLExd1daBSxEcx0V0iCErfPEgEgSKFvSCEfV+GOad
U+E5DJ5BpMZD2LJebLCLuS7JNgGaW/Mv82DXzetjjYr8u3+/cgBRctb02KM9
kkXWTFVuaXdvecm99A2w2gsEHyiyAXKeHsLggI6iTQCLId7rbrCc76CaKxVT
BlunKem87uYDhs/wyhlK1hECiGU2B0ATw3BT2/09AQdrfHY/h4RLkcJbnY77
D7+I9gUOd4FSCSLjFs42VRlzlf5/NrHS6jmR20RZ0OelBn7m6DL6zTv4ToA6
DkKKIbQ0IoV1gLxSQ1SA0KZigdwvgPS3KI2jckSZ5uA8bwvPzc5BH4e6dvDN
fchCCMqU68alIU3AQlOBR0NrqsbOzJccy//Bz104Xbkz7JHei642KZDq+yrZ
ujsfRFRyt1ADxwG2gLzIHkc3xrLFADZ82SMaTngyqLp2la80ytKBqyK+PTSR
/6TtftLhU64h2VvbO8qA3G6XyTAhnucw36KBtLpy1wn48gi88dLtTvFhmykk
0K43zK1xHmDerRTLCdGOeJ1EJxYLlpaSUU2ZVYAiPBAIKkw+fXNXeLdin0lH
TGLYBpwOXVlTRQ6uHooGX1NwR7Uxaj1h/oNG0WjZppSOJeoansMDo3XGYEdo
GNeUzq4tbQADCE5pQwTHIi9UCX9L/CXKaA1OnKzzltRUY691rJoDC2wDK1fM
JVWCdTPV+6AJWyYch9jF4AfZw0BjRweSmM55Ler3zOneBMW7Kwk871CefIZW
ci/02wlnuQhSVPXEG1UyDcriYOBNYDbqLKerUqkNWVh4LaOsTmreTar7tLX+
1fwJxgnwm+dSyNb4f4yKQDdvs6kDE5qcuFmKAvV1x+uYVMgCViOHn0QKHPBj
otwGoszcUniV1BO2RzHZzr0WBL96vvuc03rlV1YbpNyjaTPE4s4pzGEnmEiv
S9KU8Bcf6BhgZy/jRvD9bZHaWhyH+D/Yf/VYvOqF2Qw01a00ovDauEkE+d7G
RUFB//IeGDvK2UVxWOnMzytJkAbe3C7raaG/m195EEA9+ZlGvqJB0JRB9NkL
Pwhz7PEnCkVTt06u3447xIjnBtjQlEhtAxexPgkj/355MQf6QH6PblVZhdFW
PAw0jsCqAGIKcwNni6CzunT3D5GqbwfMwk5inTaoyAYGbu37mpS1O/WkAaXx
oDqVBrq6f59j+TOx6KCtG44vBcHX1KHmnNbi+u1m/g1sHY6mDpL2jZWuOjNM
jZfCaMs9J+8xHMY3ir8wx12ueYd9jHZilpS9HmcLZZ6HFxNFXImlC/WhYQeu
YY6vwR8IenFcDkNokwTevgaM81d+BI3XuobHXpZivLQMYeYkr8u0fY/GPINA
6yrE6tutrGiIRCA38WuzwzGdPDByFWYKX1SJZXONPBioXsAUI1tbF4TiBr3e
pPkkcYXK9QTHrYJAF61oy8/tCbMxf5s2XGmLZ/BIbkdGo7i05adqH+2RNufA
3x8U8EBqB8wcBgP/2IztWcod2c0hos2jcuqu++i+KSmIRMaaYyHO1nW9iriZ
8VbNH8rw7mTSk9LazhGM7m6NMUxxK58WercQIo9exbsFW7HbNK+6ZzhI7I7m
QRp2Ret43VLJiV6TqJmMp/O8Oi86J9l8qEGO24QZnW0rSj5WVry4OiBRr7vs
LPsEff4aAIJj8cjes8NR5iY9AIL25Y4tlcn+ykezPdmMPpuVXKtmhiUAdRtY
tou5E8sdo2grQ7vTSg+zoRcPNOJF8MNrJmVuCsAFWkh5QnjngjDNewD1NSL7
PaYLbw16BAVhaLB45xSEjo5pGt3PyXVn5o+bBSHtFc2juFNdWcUKqRfD3+Zo
KTxhHWpI10bM72NLi9eOgEwLiOHaMXnhJK6lbAoEnczXRQCBpnffrrrAN956
jQeqDjHy6nxqCDXTjvRe3sOEXlG8eqOnyF/07E71163Sgx8AWeer/EYhSGPI
jrPnUn26vxHAHIDXf2LbkU6Kfez9bKFMT74VKfl574ddYUCgMBx6Sip4Kfm9
TDIRQsWz81ypAoqoAmbXXwA71ZcwezD4K17OlA3wE9aNQzv4eQJnUM9rqrQ9
1EaiAoTOaWOXvwZdd9l4s1HGdAc8PZqtkpaJcH+S387kdFYgQrQyNNQ7HTpz
mPAFHBdn4aWIPMAgVsNc/CS+CJ1Tvvtcb6GSvoxez2lyNE3nENSlpN2wiZHq
QL3tFLhNhWZ3KwqQUnLY9w0dpqTkX+7RT4KsYevLbXjTb0ooqOR/yf4FdfgH
MiyBfnj/hCvB9d9NLACHQeomtktxUP8MaIoDK4EUcp0K50yLNrAdIRpcjdb7
16uodLEnIaSPyZggsQDKvqHqzZnmjofsL5if0QoP/cSFe2LV08R/MoOF6aQw
5HJOK6Y8iZ6n1VcneozXNevWzk/Vxue21+Hc3bq4uNNn1b8kCVoAQarc7MEH
PEgefXII/uIZIHW5U/pbghjnt3rjvO0P2JV//Wg9Yb9DEhUziuMoj6ViqJ+A
gP5oGmnKrLFuBAT16rUt14FJPL5qjD2MEP9X7b4sHQqKYg4sy4qy/u3JxJmv
H2pOjZj42KKVMGbOcKOO032OKB6Mvz08J+832QHwFNdZTotsZPvIqmJznT0z
YsgO/bJAJHnNUjAnNHDiXQQMTGDYKNrbgqjde0vcmPiFiVwlO7UZkQE3Lzag
Z2O2xbk7VKmg5ABPwYxUntTESKm7iDmzDb7/4/FO5lUNRa7T/bDlD/e7rr/b
ZjJR3zGyxCJl+/6qR7nmIGZ2CBgusZwMIg8HRlsfHEsK4CphqFPhIQSViocr
ObWxzdgR4fKXrvAoZqldi3FY5iGcSblma+QCW0ZURv4V2TnDWsIgfKId0gyx
xVd162094hiNz8fM7ZeRqMjZkkuhLLNXifzDLs82rHc34z0R8WtkWiLfPvj9
wmPnTsHGIT8EcBSSg2ESIK7/WNwmXBVxqBGETzUWhl0kjoTFXV+wjzV6xQg5
lE+pPba9mNkpufs+UH5UmFfOuB5BEGh41mxaNKOoRu2CYsrfZqrOcm5mgNf8
BcsauAe9MJ8SoND7fM6qP3fQP7z0N0Yw2fmmZaO2Gl1gzPWnzjjlHcFiMdmO
WHzCszMtKLAD7FH9saEaqZfrQMQMKy5yxpaWrMhBmNHDp7e822Vr/OPSVSp/
NwWeFQZdj0gox4m4kbNq+rylNhJyg5COFeAIzkVo4H7XenoJkGZMelYAhTmJ
DHbKxlJb6LAn32NuSP0qi6e+xPxGQBzks2CmAbyG3ilCV6dE1uOBGK+8qTGq
9NEm/G7kn4HrzQOou6ydqPBeRx6sJKuPvShDcR4LauJXxmbeFUWjvXavcNwu
9n6BogQo2IVmwXAYgEohc3dqvvPikh/Hj2uNl6XL1RsPxNbqmiEgnnK/qGa8
m5p4O1QmfhfTmZW8V8IXpS+0kW6FTUzPW6+GaVNSGp3tUGwiDp7JB2hnKgZD
GbcRaas1hXufYkhy6yy3IMTKkHN6pNWaiN2YQk1ldXL+E6TN1E8pK6P3g5mF
mHrmbQ4QEuhHvDrTXTGu/Xfvm77+8CAj0hplqCS65sxkXT9D2wvTgtTRU3jK
9lUh+LRtVOwtLq/ZxqX/KpXmr9wjkk+czcFObVYLdux00Fd/sGPavi0jqFId
iUCwCV/UI4czH3bjDJRtyUDOKU0as89T0fJjGATsyfvwhP4mMdHJLvFvTwBo
DWqOmoEKV15KYxwgChHoFqHrJ+meYTXcfdLRl8Y8vcwDVQxy6EKfE9hl61/g
Jo8DUalCdGG5PC3VI1ovghBspi7nW8ezBh48p/KwMoipuF0CxlSZUR6fx6dr
mfuqJ+5OppnC0g6r53zI6IGMOSxEIo2UiNBpdC3QcRaNEfcgaCmAdSIu/NHS
cJ/EEwpWpUDiY8rnxRfoca4/roPwqU7Hi1Ihxsy784XM5E8KHt90VdY9guNj
JbX9XsySS7E7QKdBOrKq7dblAF4op7/K4qwFlzg4GY2e1k0oV1E4yDQXqMs+
q0bZjBf3HCPzYiu8yyOWZcCCFm84lvHYrhT5DoJxdjgu24DGMfSl/e7J4T5f
zL8/27CMEfS53LaxPK7Yfc6bs/w1fMsEFJZ54k8x+h85OC36BsWDP1O54joR
lEvAC50dP6xS7G5rzlRJoBZfmtUGqMPHpk8B7PmBImh95deP5SteNQf5uB9U
ac0CQytzvlF6XlEesPYnsVvjY3obV6fdUgItHCANVhBUzjeHMj6uYhpMtCo4
uugaXHDJq7ikm98VMlJAXhFMDRuXMDIlceeHfTUWBMRgifltfmN5NGuB0DYo
0iH/gd8AtTwW7kzedi37p4iet1/wiUDbgJz9HB2bzXO/iRreLm+ZuUlZc1Mn
Mziq3guYUYfAZyxjzm2I8AcgdAKVKJM5xt9kBgc+oAf3WP/uWa7LLOgGv20j
Wu+QotFx9Bdpn55YS5iMjGMY430GpclArHGmrb0ZWls+AEaYuCCvQVWnJFwa
DkkJTBQ/d+aesZZY6PZUeKj36d2VNbIbtlWd6MjtuExRqGZGAafkSNXh7k+P
FzAR/owQg2Gr2v/rp+nVJh0jOtZr/ip0gqTTN1kX+/ueirF1FSY9S6jANmQP
8yTVnHE0oScr/hxTPnheeHt6VSfZ9L6ly9X0FvfXE7nUssca2d91jF7Qr+f/
/cEu1rhTKF1tUNZPSkvj5XhsTjR9w3xj/2AMQACpnkezgweLn5ktF8QuZOJZ
BGOjVy3/ZjGN/TmfeBOtVb1n4gLKSPeD6C1VaIe4AT9rsBrj0VHZCeCQ8yx6
9c5vMYlu3FfERPWA/IpOLBqZbe6B6pGtKPGhc4s5Gd1FIO3cxPHUYndPuM/G
x+NAkqEOrEJDxq+8gSpADeve7pOpGJdvQXgtyA8izD1ZCxJRiRl5xJmYoBfE
V3JrL2L8BX/A4pCS5akGVUlXNtosfNsXi8GU26EABJx1NlsLin+pcCIiWcM3
taLnlSPCqyrrCFkaCB2slVPRKKoyW5s8yCToPJmgWajTs2ydzp47Tw8AXQdE
fgITCeXoGWfpRhjfq1MBRRaI3N53uEn00+cvTzg/gXyfYPi8gislfiUyYPCa
c8fXFoQEwwB4i9sAChvjIv6Ukf2UnvwfHpgVwdqLTfZzz94JOVYWwYweglha
+VaQ5Gzoh5JWRERGHqgGTqauXeKyMnN4VABk+FaxFF3HRuNx09ffvZ7dPGbX
D4mKVi3N0m1ctWmYhly8cI30J1Pq1SB1ghb6g1clPGSzdxc+ZBj9JYz5wjv9
Y+hJ6OJCmy0Of9Q3NdlQ40VRPlEMUTluhpeGwJfktNmUxFAzRFnXbuZIhtZe
u6HtnhenxWjVMS/hDHS1H/yiZtJ5i4oeIa+T+wtybK8cwfesEQpVmcwSc3O5
CosIxBJaf5aKcyztAtRnKZzPtmlnvAR2BUjipVxtM1ba7xx1s/Cd5qmqZQ8E
qV7o5fsSVqS8NPRN15vm/rGv806vYXuOMceIGupEoIsmxvVq+HpciH7XIALb
Nn5DPTghX93sFSkaBWHDYB6CQWhxY1qjeu1MLGsbGEA9+Ves7XFt+qKaHWVr
BeSpP3nKUpyIWgMzj6XOjB6I2HvAL0AQfl3is1gk2E2oSjZphvLRF9L/wyu6
zybAXjUbm1cn986WTUEzCFpIMI77OBoX4kioqy7ihbt9mPTWZmMly8u83eDa
soZY+HKXUap5KugQ5E3ma6wxOCa9GRzDEHAlpw0ChfmGsQKnfGFsLBFT/JRv
z7g+UJKW2G3ljQHyjfjpHnF5SeO5p8pgrxyrmSLbBimvGzaPV8aVFaANhu11
+t9GILgmp72HZf0uwtk489jrNRXFbaf6MpGGGafUC6fZFhMxZgkppnyTZMTN
0r9uXINQknNYMV9h82FS7tBGsGxqqEwbKlt2o3D71VVwj4N+0JzIbbaZHRS+
DrxIWN+2BMNekWsdF0x0mp4aiU7rRrWIEVoZAvptgAFuwIyYOi6xtBcSmkuX
zZRqViOlyNLQR37MCJkNCP2mC14pHkLtdbal6LnvffvOmz+p2aJhKfzS21EB
3NM8JQoL303SHhAmhZz8cZH8A2BB9I3v04ieMLLPX9QQLN887p+WVEzxJ8KF
VRvLV9+N2FfkRgQesg0rt0OZQvY271jtqD102NWkAUENFvkgqvEq+7ktCY54
vQpZmvV21wYk39cm/VnCEAWsd67kKED3USD4qBY4dgq7cBJq2ccGdYLe2k4v
QiuZ58EB6yv9uo/dEVHRGqLf8ZLpc5xb5Epwb2mQqJ0VOoH0d7Bz8dGSBA7F
Yfc6SRGLCrbki9n7t5enJh4XwnaX70nTztjF9B3/9Y9G31RUinXMVbxUGPcj
nLNXAHW+n9aq2340ZnwPgfH8B+iLfHC6RXY5Ek76eBq1Kf8N5vJ3y49cTStS
Z3ynXTU9xQnD5Qf37DXAQKaZKcGOXK5odKDmFNXCSTEiFPr8BOng6l271lCL
gNfs1Az+VNWX5TccIx5wJJpQstHeiQWMex3GEGSAxsXku8UahS6wmqcQCxfG
TY2z4Kwf1PmGKUQdb4kk12UKCPV2NJXCC3IbMIjKRRgFVXl8HuSwJL0vhrFY
qUN+a57wxsJ22EjiIr/oH2JYt0JohObaDCTiwqFSSaeN38yMemdxiAfVYNbx
TuB5tbl/nVGQRX40qI1ApdQoJPOH8USEmrPusHl8bpYLzFKZTpuwdbj+sIhy
ZA/ubxLhYgcFX0yxd6WvhB+Rqm7EKJrNZa2IitJjQZwAZEElSa1Z74g9fK0H
F421pnJW+gi/hO5WBBsVWQN4N8J0EtxuLb4RGr1URxWeOSU+6pxBj9ttN88+
oq7a/y8nUS8sv1tQ6Cpnxq+EqsNO4g2IN7TODy41yIouFU79Qw+zPnGqWWif
gNCYvvdSDlQrP9yJT03lllb0TVIffMhT+Er2vPqjuuudogHsxJos/6G2DcpA
ZztGW2YnFbsfFmA5PQHk82CQVwFbhQDx7t5ctPgaYeGfe9zQbmzEO+FaX2+h
jXUKBSPYfnIwZSpLDtzwJF05e1NaDGfFk4JiWEUT8wuu1p1X0C4uZIrEBKY2
TsfFrcBxRzjtmXlx9mbwJgbspWQ4F2wvOC9LdoX4oPcsxnSWmWDtuqPU302P
o92nW4ohNtEvzLbMY3HdD5BttBiwvs9dJ4X/M7W3Ra+UqJgKhHziL/vub3P6
p5alrEHS0OobA4DaE6bcJ29AGj9C7g12jE7WFhJtyPs8mwsVAjnk8n+vNytg
ZDokWhWxSfxy3UoQ6Kel3T0KaJEbz98+LO2j+k7kZJMeZ1JepxOLHgyDVg1g
gRLGpeUpt5k2zlox/i1Wc2mrUJo95iaIXv/ZCLKM0ttPXsv1dG9bS5MJB4UI
vDoWoWNUx9pjZmd715kSgpaDRoD3tzjm8ViQyWwgnNp5kxoYvBkgYzo9o3IG
hvXvqPckJy598Zr+xyCHefEuIgbhsHsydOJOwCI4KCUxtHIo8ZZ3ps91aIAI
GSNm10L4rMTS7ygoG4uoFga4kqjjn+VEFm+PiMQ42OXNWduSTGAHvlcJ0RR6
5fAt1vzaantm7ZJFY3iKIBBgE6Xq+fISeHTtFa9toTTUwj/mTHvbs1IYG+9M
dAT3a/VAOxzx6ljdcCe+B1cOLeLm+XZrfqQh9mCa8INRnx7/g3hFARoTBW+O
r1IRgNQpU9U/4Ja4/nVrvwsw7gg0z0Jd0u4IJzZ3v8g9GMLvDB+uWQWwt82J
nTIMUEeHcgcnVrJPNorI2T1s/7Nga5JBg7S7InQAl+vY5YXeZMNgjT65c0+2
AVRNq/9GaacSwFrJsXOhl5QsQ9678YwhziQJsCvBD5do9nkvlGgAmF4hZ5ta
U5Jhu2PRjlYSiEaeOZ+WSCJ3N1WIHfcp71lYTF7S53Wghs3MbWSFVb8nnaY6
Kxacpfyu46VEs6IUdoBkzpdtnY4xZrFZsYRCI5gevE81ro5IMgGd8NOQQpb2
OXIl+RIbNYVODb0N8+eR0tpZM/ynBoiNDjrSqfRqTOL1tVAxg6XgBYKLlcIu
bYgfYOCXbgjlFHA6pKcFnEIXpEZq8vPN/YtQt4uuyujccz2TZyonhPO0lWt8
xdpSrf3xf/nc6rUW2f+S2uhyq5Wm1pmD/SKURqIZBfYWO0B5C4FrabcbrWwA
v3VqM/Di+3ZVN716p8hhG2NpZyFroyqwKm7Mc4VbyWyQzGxx87H+3oE+fSYT
KebDX7pmI59U/g+/Pt+1zqYCv7/4cW1qK8aNpGqoipqyyGE701CpWyP3cwQx
w8VUiGMxfpea/uAuyIq1wl9VViDkoXJkl0wTNgXteBtrz2U1uSSNykEJ1JJ/
MIWp/DiGIRO4L1xgLHxePqcPWA2DaDWpL9qYGtgZP0Z90g1tKlxUqD8OeV3F
rQOG74hKzbYaodYcK/uu75i6upuDuHsRIWwOemsbl02/iEsVaZ9MiSKOtmaz
jk/cLZcs9PLa6q+imY+s32yjKR0fz8StBedxYjapAl2dMFbjHtfzTV4tUYSH
H7u8XWPxPJwmgTAussdPWWhI84LCaYhPAYsKaRMFPCouBx6fgWS7JjC8geh9
AH6qfSOy90LHisPqy5mM4AdjfLAvcVngWBnUO5GDEgNO785P2HiQC/70QVe2
St7mfHKh6NbIM9IomV/wbUDqpjcGizB57hLAh6AxYqbd6JjBbSKyY4pKldNY
SZYcpX/D54B8SjB/n3a5tR6grG0K3RdSmTju0/jVVNMAqnqBRaQZTzsYvGAP
9kzjoHleDDLX8bpdlQYPkW8iuvcnGvDcJcS+mnJcN7CZB+59phHujp/4CcUZ
Usil7K5obK3ZGEv96WPHxPMtuRZkwzrjsyLmCzjREyBYNKKs+jcrv4zE+FA/
QrRL4GeTwAPwSfH06/WOrWJL4zE8J7vIfuVD88Tsc3Cq7oenyMrBCkIxzVaZ
U6anDHKz1wwcYmhRBWqfZYoXhbzqoJ6GmrBIDyGElaSkHdxzN1hbaqIrgQZu
6TYK8MbLUQY0LgGCQrHnN8KLg4oLNY/dcNDHhaJo9iUzjDw3EB/F/HEgLUht
fOLRpm6uW/c8Moe2EMhPyRZb7zm9grD+k7fqefPKWYTO6Sq+ElIgEfzG43qr
g6dcOcZZgnT+UYGAkdPpTkpsFCa8Ev5EW9GrXn5eJGXeEdKVQsp6P6DcDFZL
pLAZc/MtHwO2gcHWu5g6resdFyorT9f35GcIuD82+DVGFKbB7gpPbdwmcbs4
ANumDj7WMvdwb+I7h3GinYf/V0glyBIckiU+zN+i4r8wtD0yOgCRcretCmz1
cV9hec2kpFIxItfZ51hvJpPGvPFzqWolzUDR9PkSitKuHdxGrAYfv6uO4KHc
9ER/ZXdZgvYE5qAoq+P1OJoJFiCbpzkwjhOkKIjK+qXqvM6sChKhR3B6hbFO
SGb0eD3WhAm06/40bOvciA5xGgbv8SnwGLjmBthPf/pxyID7+Ka0iH5pkEcq
pGJqPPPTUaWKfZOT1FLAT4cxrM9qKOf+xekFlSn0FweOP6MynYo4WC2HwvC8
NLYklNX78tibnbndrI60PozdRyIEgQ/SjkxCYtDQ+h8GmT7DN65YD5ownD3M
46udDXoor1ZQznyHJj/08UxbK+SEgmGBMXCUQMxnvIeKXeb9VdGqTnWv5/wr
7jdvjqJyGx31AI60QddZpmTQuPpga9WP4pGAq5rkMXz5usdqCHZ4vCJTBa1m
d2bxk19OC6t5NwjiTGu1hnmrBmAJO/48WYKFs03TfVJc+Bee59nnmGSA73Jy
eZ+1Z8tvb7Rak53qZEXyHWNggAQIfxoh6NQUj8GlChsTQxRgOHhkalBI4FJ5
lVZqn6dVWocIovKOaO9kPd4XRbdYSCZfahopN5lllvUyeqgISaq6NSDnSBII
CVRS1M4ZW/geIAQYwS6hP42tXnEdJPvneHjGbkkWsEvaNxArmwp/27dcVTUD
65/fQL80JCYn7gH/3n8K/FqYWWStJJo1fP8nbaMSqjThDfHIuARreE3e7Bja
30JgHfkPbz1NhQBib2AQdJCs8nKwlZQnU27jNRIHIzfNMiPsKEYR1T37Zynl
T7cyl0Qx+b/NUqJbD/xsnXOoiriEsa46sZg6iVecakgGsOENZNPL4wXHE92H
7Jtx67+kJIxZHXU/7X6X06R0g7IHFVECS1XU0FT2EH2h/31sMY6qjStmOLdD
7+G4RfFRdt/YkYq4clZoXtoDmtGS00Xzh9xfKk+OHBqBiw21Wu3tsfg+NkFn
iWpE3mr42sLVx1hXsQARPfdYub8Gz8WvWhwyQwPKqykTO2eiUSUV72TAKqkQ
hlZPWpOlRB2PcIvtp4jDdNfckY7mGrKZ5BAKBWdFnYUlVWwP56uHp9XzYrTv
vQ9r33uASE8loQK7K/G9R2NEa2tg6niy9BEOtyFZzswm+DqgjdjN1wDRxUHd
k4i77gCa3eBMWS/KxkHLozKOtSyRN7ODYhnu+p3GAnYFkMY5iGdJZT40iRgZ
vuM/QEMOlVE05lg183EjGh8r0yH4I264gYxJE+zLIKXKXz3/gxnCHXfZ00//
L7GQHOadTADFyweVfQIoyfcZlUumHVa5nxOTUuwYrNRMOrsENDZw0ASfv3d2
U7QmLRFsEcimKe796uuWfYmLCxnaUaREV6i2Nux30RTE/Nlm8EArMbOGoGf8
Ma/ajZONW6Vm8sdgNcrzYMpbH6smjWnuNUVe+oe/jvpFID5cfqh1/V2O9xrD
Pel1svXvlOmBAWG8UVXAmjg9u6N202usB/bUVICb3G6o1o5zczYqrMFQQGqE
LZPqY8VwwUlbqhUra+5Vm1P4UPlahRsf2CpYk2t5YbI8kL7+LOjYKsyXVm+x
Rgt/3N00av54/ZyXzVIxDfsh8YvJDbPL+kg/mckPhmwZdKESO0m8HKaBSPwI
NOjLJKWrEU+HPlHN+dRQWZWPic8NDkZHCGfPfiSTGdEEcLDl2TsnXp4FiOTw
suPSDO4qgvD+yArWp6kV7RcS1mNVzuhztKoMcoOH6fiFQgUe6EyFuAt16RTA
w6rrvu0Bku1HcsSyam8J0zdHEu6krtfTWG0K3tgEy3F0WhqSYafXHy4AsL0Y
DHSjGZtmTP4Br4+OD2kG+KnTST5iBa6hPI4lGdSGC/yp3GATxK0MzgBO8Dxn
2ssaCGIiqZ/YJ9tISwbmw0CiqS3Fsc7EoqzaFDr5lXE2AZLvqlRWFyo0M6Pe
9Uk8UvRkLx6X4GKaIynJZnHu8pFT1blurStuYCyDnGuK+34+tWdy6aCpvVl4
d80f0+e96ZYsgOAG22wk0Wpn5jc63eGI2MHJ25UPAmZobKOGnlFBDoYFV1hA
DSBZd8vVkgJRy83aNwn6rjGNSVYa3DlGAYQdySdTw959C/aVBqFZBU4TOvqV
6Ar4SsE6EfmQBwLNmTLa8p11jEoIQ9VP8x3iYi000CMqX6oU1Uh+uvTUOOyM
XA3Bh05RsYzqjmtQTth9MIjiIODlgXb7ZTx8x4EBn7mro6/53aGF1rWXEBxG
nQSikhaHlJYdb9RnQ8wbAHzzzGU19tqMAff3hdlvQKcc+xYKM1FOooJERzPk
8OE48Bi6+1ReZSZe77P41GkGm/wvhX5IaKk8aa3AcWmUIgDpVRENbyLDCfq1
pTbIsVNnsidvDcG+vO/mkQpBVAnyyShQFhODRK7PmqsFg8rBVdZrl1wPQ/fW
iCd3l0GtjeYEfRTkh32LVEbHcra6PHdu6o4ZHtpjSAELmA6AtSe7m9fHi2Hx
uuUdUkiAAkIn89ii+e64hAStG8nhBnVkGHyEWNXTVE+uZP1J+EO30gvWmf8Z
ocLPvm1s584hD73ZWvhunAxX/XTkno/7KYWb1E2Cwa8D3FgHVBuuK7yrOX2W
VVsf8qXUf6wTt5OddKPIeT1f57KdsfglO35zS+41LJxEGop1TtrgzKyyHSEL
BLwmrqGia3UjeOgDaQU0fMx9+yc5Rq4n0WJjPKjHYz6rNOUd7U2e5AP3QBdo
8DGDYHXvDeGVsA+RUwJk0FbmYJtO/UzuokCk31ZcN6lzm/0wfzXXsIkgKi8G
8r+yjRwrhnadW1iv+Eg37YqxGwkpnh4qeAoJqcxZGwOm1b5xLxAT0fNmPt8R
pgNsUJWzOOzxj3BHBmIN0yN3fCwJVX7WbyS9iU9nzGOANXjp0/aDNym8pfLB
xG20TBPv/pEqAcClQ7Z68WjiSiU9u1p3do9zJljuMEfYlLsFVhlkWWl4Y/WS
wBXxi80rYHvd4TIuWiFUFeICTXpYZ5YiIfjPQG2hexwK9EVZky3KjTtZJEDR
Zqp4VwSE7eVbNdo0voT/t+lvLUTiV8nFqtQ/CMGxGGtChzPeUxIrEex4YK+L
U08HHJ9QSLrR9B8XLSQ4BZfWF+F4VjjGPSq6NqVyj9zUlHoxGpHJUQFKwH9T
PjlMD4VryMwz8lKK2XIZfneMYHZr2xNEwbpnzG7+QwAWLkEf5O/LCOsBl1AN
2KKALr/5U6t5SZigElLncBQjmZHGHJYSf57vbWAAwwW6JaSEfrvRllYj7aXR
r9HsJ61iUiscF1D4z3BKaPld+yNuF5wUX7DeteUiIKxFhgmfQk6WP5fKQK8J
PI4iSasfaAXKIbYFzEtX57zovG1dOEgTN2MEu7l2yTsxbi+EkLwCEjh4D6n+
qBga9CruO+aAQi+7YQQEISmT+91WpaFeAcjj8wvvPEGdGRlzn+Ybgi4ELs6p
lNDWS4skaOnxp9iB/DgTrrRMA9iyQgPAIYT20guWwANrx4W8t+nrEGWXCVBE
Nx0Hq6nT3odVKVuttoRb/VvOCpeWhN1G+cEFelCKI8Mll5Xrh6SHq+Ls7DCH
OBaxq3o7AFc8QTOm/U36h0ShsjpGEQa5Sh5lZmHMxIDGz7VMdwEtCTppxIXK
9Sab1hinh08ie7vBiwAwtaqzzzkYsp5SBrP+TD3bZh7qUNyplll1LZ3z9aX0
WHA+Hit3wBeY3OqngtPSWBhNTowtQtNq+ZL0TMIhNy7OMvlCs7I24IT94yTy
l/rgyneNh05R3SrZEXN+4NAT5JtgO/99g2MBvNfE12WglkkCRy078iu4uX5W
xZ1KyRT82qztJrYIq5qV4upU2JUnuztPL5vjtRzvQ8Oqtg8CQ09HVnDW5RDj
7W3GSkYpbxQmUKoPL4OIZXPrJYmammruUfvS1+zeahX4sSLSwnTbgR0RAKJs
YXbtJ8d+1DGIz+Z17rl9K8GzSy0xTty46Pe4kvOehvZcv759qhNli6AG3ET0
OGlcAWvTojI3lFCC0IAGoHM516/xsQC9f9/v+KHvdGW4YJ27e577YqVO9+OJ
BX8i+HOSqGDhYY6ZGvIOk88fnb7RKf3lmrRkXOEBl7ihGGPl+dhOJoFgKTyU
Gp4BZrKffu5NQzLt5UKfHy4YC0eHsJxytQepeSwxbDM+YL8yd8KpywbvgHMO
J/uz8dCop+mvoH3Ry6hkM+FB3iIKCZlbDat9kNEPQaXPTHgR+DoJ2TUScxLG
HBmducnw62zL60JYrAwbs50vUp8agqTAoPcWWEKhjINF60hK7jWHwJ9BW2hR
5gOXvEDVumIxFZaVUVn/zGGCrKByd6FemW3rjwvxPQ1b3HqFumyh2L3b4MZ2
S2O+UatD0j2hswDLgP4R3QhivgJ4Za+anGgdi6n3efGTd9NpId7LdU9qPgIV
jhHnKO8VhYb6K9Uit/x3iHp0PXYZQzFbzMXbKmz2QtND7WkiZj2xjB+tN9+o
rKk0b93pum9QkdW508sYK6V0xEF5wkhDMVLPyoOlNx44RqqmMzYh0WiEK1aw
TNAIXTzyBvxdBtYTi8/JbiegVtXTDVv3GWR/C95JqPt4s7CYynLgmhlTNrra
mRKTTXL+37G8lbT9cqpgPoN+uEhPJvXp2vOT/08YZ8lzyucyf8eJCqqDDVoh
vi36wBvjPeRonw5/FpYbMUwjneKfp2clAOCzTJdPf676nZ7vtF5RUoS8EK/E
ngDvdTqkJqqcxHXW5sigYJ77g2DjJ6pfQVJS4hpXJzNVFJCBuqeRoFoUN4yq
eGi5ORAU2sTX28GGwm4Dyi9xF8MZNP2Sac+mxdIqJevn65QsJKJT+yQqbvlp
2/xDSEnswOO/zVD86CGkXHZq6xdoPpRnZDSzs8GvS6A9dffw0IgcybDSekDl
nujbMjpKMaf8dMFSEPXLeOr0oRa1P4N/PH4U9bMLyWUa760ANH2rFEFrmr10
lKsmJJPvPpxQeIoK1DrqEP/3TJ3t35U2cLUyLzcHxE6wBoRpNaU8pnV5w914
H3IkcDfDPK3aSx0253VAuOuiTssrAs++Q2g5pLdGL3+TL2izcvj+4kEhDV2F
48ypuOHq/cLxHe3Fm+G1IzCnu47IDXqxcTpfcPD0Nld9o57WJmHmtIRZPmEP
lVsnosVS9bUwhP9F3gel7VPcBW1OaJlFxUDgOUOxffGhJth/gKZgrRGwb+6b
atpOsUctTMl260fM2sbrWuc1dEl/BGGOzkN4Aqj86AMt6ZLJudhe2Wu4Csrj
CJSjgtTbng/QV8dUOBSahF2UqiCkCgdgC6D8aRII/WZA2CGN3XpHQaiDyt6j
HDvBnuf9SebtWDzr64MdGc1/hVg1ET8EZ83UY2JhQFAokrXV0oR5KWAco4vs
1QcBSv/5qTxBaJ8SKZ30fhrZ4T9C3C0Stoiv4Xc4FpIzWeKK9GXxdllQEB6y
Ug1ONlHVfrR8lkvRxjtKQMjftt03Dci1KUKXynGckCTewprsU4dvm/paPkLd
Saauh3pL5f/fR/6mSXPUYSk6Ax4EroJs2H/ygLCfPNRXuluhcz0yzwsgNdrT
AJUvZFDkEtcAvn+2C5/YA6Pm71wB78LwQFU+QlGJIJXJJGylvshGTxkcjCrI
yEyIG+1ZKlgGojxAERo+ANyrsCQFwl3R9g/m185CpLYbbZCPxzbzuaavDLlB
aXM7dtSaycnadnW7LCKQ26jce802utZ7zDBV7HLG2DqcNoDqw0dsE6EUwIue
JL7t+3B1i8I1rz/UVZc+voO33GrL3avRpQrtcc/nSiGGjLZ8T5XA4PE/Zl3/
d6i+r4acxd8yk3izgitLXSAYxLqGxsobJmpSDRSrgFXKoSJ1xqptX0+vfCzJ
ceNKdzET7FxJxw4MREQVOHJqGwF+Ptf2HItUBgNQm6dQE0MF/poV5uClrXcb
bvsm49Wb1Tps4c84Jj6ZPPzDBU+uAqYyFJM+Z+IxawP3RUZ5LdpuTQ0lt6Rg
/za+wFgsnDYaUm98HUjlH/9XKZUFlw1hK/LabQ2ZBjPQhFHyxNybKa3/bVTg
IHoVeb25m3Uh/89YXstpg7SA2+rSzYQP1FXWG8N48FU0gNJMMEYhcYzchO8c
Hxm/d0rJrbtvT71BajT+SD0QlZLHDNbZBmJxkXmHSFj/m6GsYThTOyjKENLP
JbMNOVEBsyUVGUiWu66nJNAIR7CjMrxrCc+pn5O6KRE4sPdzUNuovTXeNDK/
af6Q/zi0pmI6DPU7mi9UBz2VQBEHXUzn3Jo7wUGXPNTSflPleYTKlXQmMWwz
EPfUnHY1Ul9EaRT0OaRhUQ6ReyyCpOKDOLvGC9F/xExklz1QshUyMp/5TG1r
GhmifPetHkNefN7mqHmrou6tf5e0F/4X/kQ0Xa5aRpHk5ODMe8P5S4RtJHHz
ti5sGTMLk6w2c+uKwsAqI3fDuO9MX3SlrxDtjZAXNQcXdRg7yqkwj3wJOsl7
R7nHWKQV8P/26Z1OyXNqj8By4gTZOusup9hz+E3yYdorTNLTG7K5pzhVqj5w
a2nlENurHoBECfwkCeUkoQL8L/Q0bMnUpxmmTZg+L5ffiK76BOhuoZA20hZM
5kSz4ROaL7nyTNmxKFCkPnnT2kefsngrvdI1cmIdooi+avpHfjjg7BNkmur4
yN5semSi864fXNYph53nSogSIzsSHh42UAr/okdzknyLG9Ev9QX+GLiTST2n
RG+qmKZ2KF2syf8nqxrBRjux4p/FDU/mdTpCaieqq1voMSDx9RIO/OGEIAp5
3nVAduVuieo/VfbMV7Ut7MSsh8krEMA9nJESRqLtKPRHb1KQ4ulycWJCN8c9
+/7tbl1rvKUlHWFvoFd9AaFXgTfZ9i+1PwfIlxIlxayzBKCI+vpFGzPnEAPQ
0NLgg3+R8r3hkAKEYDVMsrrhskYKOvKxroclh39ovMvtjaEdDPyxozlFKgLq
v7lqiyAXNB5FHVGpmfL3PBOjglXPDS+MPVzdCgaX1CErIhhUKbmCSbTin3uA
WttjIoecd6XrfZv1aLXzW6shBSP1KxZeM8h/I2/aZsfiOo4Qv4zINOPlhJm6
lmQUuw7qzCE/qLGDvyXyKo6X4pAHWVF/VX49SJXSL3ukMEpttMzInZOnQB0O
4S2CHLhCu8byrEoLdpOEzdw5OplquI56Fe7RttufHhAWHBwPwMeJ8cnfmpAO
okDfGLKBkyu6tV8Uuu7AKSVsL0OwgsFZGAW/HAwNmhre9uxaFZEwnFqMksWL
Dh2Ojoy6oK2veNwX09YOsr8hSfEyYh6HJ1CL/6NsbGOcgSd7FAtcM6MrV4S4
KvTc+dGavFQlBlj1SGwNGXMKkGVvgu2gvJnwObi33aFY8C7+LcpmBZYhJGK0
3ySuWu82mLi7BliqzcNLc3rSnKBAZihSx49IIV6jtH7Kj2vZt26PjZfGy7Z5
Ltn9J1lkAkC46MIWWU+WsAutnylsnF/FE+I4zWmRq55MEhsVsR4+vBYiaD9B
OJgFbqcsLjQGHHJWExlQJQc4vyos4r2/iqiXo48vytURZnfhLtYxjFH+r+a1
eoojc990jrgJp1hmiOKy0hJuEgO21gf05ZRPU9pKIgFU55yQD+Pbo9B5pdWI
NdSLSkhQrAx1DNrwEob3gn3KdO7RsTq17nGUbYIOmnjR7/xS9db/T+ejAPoN
trhqFODeW3kQKJQAQP+3KCnCF5UyKeSoI6YQBjROnXtlCcU9+1N6qlX8v+ul
V0k1SAVnrWEPTjpzakwVm2tJpornfiMCFqbQSqU7pS/iLt5Gc6jS5SAAeJ/+
VZH9JROdd8hvdMKIz9yH2DWRWY3XW7d8uLJvXQal5s/Acm7DWBo5jFGHCn2I
FgmzGd4vzHpI93CmzD0BF3JApYcaYELYy5ox9Bvqv6/XUvLHJMUxKdJNxUFj
LOhlH6qLVo2vKtYiC/I94MUmOxuXV8jRzqmLROy4Uj9lcnpIzrOBWGwtQ84J
9lDXL75AvkzcD95oXE6tdbGBMvVWPPOIHc0Nd6mt5dWuX7bx0oauUZGREBwH
Dcvgu6HvPs5MOxNqtutwSs89UHwzn6mpuRH8jrUnFXpd2WNTkAAJ97HWs+Kv
Ddru/Jw1ZZCEN4diZkxISOqKEdyBkAEILprgaeHY7w4KdFtWmeoz6suh46Kj
MmOw7fX77FnC4wDfW2Khzh7MLNz7x/WpajwHPhmAOiqxZHlq1CCmARyzruRT
9/pYDisXXcXMAy4NtZmok9P8780eIj1YDzu9J7nXZpV28OH+IKfrVJs6jyZH
eWhNmk53pSXzjHxOKyMsYb9oCxE1KujaYSpkkGc+vPBMmFbkI8s5rTQfdVP+
tfBc7RJaZDifPkV6hzoJhpzrOzJSkHbpaCUHb+YJ7pznV2lgSz7TKXGEDwlU
a5S502MReb8dogYIuqo0QaDHaJPKqyfagXxcJCznroyoDC3oa24kUZgh+/MV
gogonapVCPzmCHf5Di5im25cUUqHGuKEC3D76M/fqk1kt9094CghAMkista3
D7NiTyebLhrDScbmotBNnkx/8Homj5BdqdFUGTiGjzQcASn4KyR8VKfVe1Q0
wq5o0VtiuG6zZX914xa5w2w4sUjOL1apuEhbno7WBh1TZh9PIBw1XBLCUiWT
sVD+b9mi4VjaQT+jvs5ugWs45UaXpQxccfEL4MDzzrhQOPXVQDvdPUKaCP+L
C9UOB9oLMIsjL7KH63WAG35mCXl7PhhQMPu0XdQZ+giYUZTCMRHwo0Gp9pVv
8g0SmwK1UbN2wdKbSHzluzhtRJJ8Yu8MooSC7e2s9GLoTL0D29aHOZozLsCd
d9jSGzJm7FHoFmWh8vzNbVrG2G/l+7NzSexv10rWi/muaeGIX7oEK16nF4uA
4EM2yvBIgjkw/wf5JrFuj5VcZIi4T/xKFor4AsVERn1w8rOQK5DJ2hgF2KKY
JzqNe3qknhLhGDxZ2E2sy5s7XfCG5glrr1Z1U3oJtRJy4c83qRL5WemfVuJ0
XLH7p13lb3tacQvOkx6MpdMQf/Qkt6rig7Rj0WY1Oy3tg8KKDS2szZB9oTqE
yvAuMHIO19xkoN2G/l1Gxk2/7OA76hDA0tsDQ5S8Ad2B52txSD0HmKh7p/1I
OxaIPoWTJ8T4Snnw9LRNCkRuRtMNULX/+zxtptlXHftc3knx5SZchIk72nAc
PqL0Oh/FU7yZU8aZa2US0qVTTw9xCvB2GppTWC7+1O6moyvBRbTD5rFEFIN5
umHG4/QLkEEEwIidNw7sj2v7D1MBOJzfip1xJvIeAPbk41w2bbXfR8l0XoPb
HIM6kxk0dFpTuMku8ITFnJuhVByNAZGRRUyuM1WCpsjx9tojO7nI2bHFScwb
xVdeujQVEfU5gw3lgf0nJMI1eRuO5W9RqQfSfyDkc0JtLQRDm/koIWoXOVja
KTLTxQ0HVyv8CkJ3KIgqOnj6TXiwKZ3eRTvLqCggCAh61kfOKJF0f6nZ6BOd
LYNaOFTxZ8EJqCA8MZHrvSTrhit0BFL4xBInkhtO42WZiPx7/STeY26TaSaz
+QIeF7vBMIvjs9Qroa7MYeZPH4u4X/oi/QzKUAWRGnxnYcPm+1+2fqHw6y/n
pW64mTBgjgpXBcTvgedcLMUCxYDqt8OXm8LsE/WQs1w+ecEmMSoVpSCWtSye
uqK912qHJv3OhYGl5tMOTAFgRrBSVGG7jfIfJ0EHzgyxqu5/INdRgIyq9DRm
d1zIe0dEqVMyjqxetcCQwqy4nRVq4iGw8zo9b5vQyPQ07QergqIzX8GlK+T0
E1lArus7COgdiyPDCQsv1ZWHuRmqEIEs4t+OG6Wb3yf/0zzTvP1OLzN6YqpO
ywMDrE+GzZmkYDZNGC8RuAHuSFFlJ10dG+Sysbt6nd/8z9xbD749PqaA5poF
m2ZtCmbnG9o5RuGBqQPgIbufe0VRTF5X5B7DiWOd7xKSeUY12CkyG+aiB5U8
nUIz6UTz4tI5NS2WHIA7oqQgMXURtvwVbvc/V9Y3ub5Ej9z7ELP1LLLEXnm6
BQEnrXAEvOoyvNkXDZXdL/y7XebqAPcJ6E2EO+ijkuMa0iTp3Q1S/NoUJD5V
e1Ta+bFGxWiodvkSWHD9cKsNQ3rihHXjZweft29rQitWBXF+lM8EzaP3bjUl
qpvW/PBvqckpoIIABRWqsVrHyBI5XWG2qU1LrbAanl7TwOnZp4/WOe3Bt62O
Lg+iy83kmGFoq8ifNrqPmqBWQZwGdrppNvie0329BPBhb4hRIWcKR1YWedkx
6OYjrNdmYvZZJlrZMw3HEzYZDooGfLotEGiosYP+HJn/CyRkhU84yRXHN+t5
fz5fPlAwBfK2opNiA8PeYUNyAiPQX2ehHSAhjAI/ezojYEjkRxBxYSA5nJjS
vvq9qD3pZD5iyp2qDCNcgV/3topi6f++m6mJYArjRfdKDz9xhJWzfAivPI+2
JF5tfCuXmORk6jXGm6Smd19Pb3Rznil3nFz8uFOAFUQKn0BG6wJKK1+PUqSo
zvluvlN4/0skQLczXARnZyCpBu6PUMb+eNfNvlaoH+1ccT3iWYQvwuKTJS0i
0jNJIo3bPRPZTFHG2R254Ma1uGFq82rDA2EfLAxWWf++tVHGczzI5o/MASOa
c3OF/VCCNKe9Tb6ejKyNOaXhverNo4qlr8xzElVUm2iDjkjPgzE9ibolbick
anNZf4aeG56hCdJGWrYsFlSZlz2Vww08bvt9+FeCBCPgjLA5T90amUqpxiuD
4veSHrmNIW0yC8dEOEJnp7ztvaynvZmsU37qqO+vmnOifJCl2vHl4AFkoTDn
N6vc0elz9EDjmWUNdix39UXqDZTVW1+1FKVYn7RA2DdJSTSBDjZGNc/J3wT4
3/gxAaxH3NlDaaLbAC1fepaFxRCH5FivdLMUz4Flc1YofxrgJ3MA5dgDOmel
w75i8yO/9huE8AoUC4JuiSgxwtKYi71yt/RArEFCpqq7qYTQUb4URjwmXTuT
k+JKYuTRmSr/6eMLIRx1CgmcSnopcxN9Vb5aXbSafdPeBCb1VkHDgEt9n+wR
y9hesd1tIG4KlxmAHe9xkZSDYX8RnmxHCIZpZZdPzaZgRFtmI3AmYHetiVqc
eYSpg502DFth39OrB4mUa1tHKkzlxdyyivrrVElIbM5B58O3GjySD7v8N/Q/
IxXD5kxgi4H1KYt0H4tFAve082ShpYBTdn0Se2g95Vbsd9PbUf0JHkq54QLX
fwUWVQlWZvC6ztT3guC4tiyPVKnSTrccrIgGSO4b0H9i7YVUgFmHQNXXJ7Y1
ekYHn3I1WkXp1wo0UwqmM/qf8AEZQ5Nj445ckuecKNLrdVZcGlRZxtPCVZR8
de8UpOxILcjB4Jw2jZNGFTIoi9NcPHMTd/NlF93N5lgU080Xe1MlqqMMbFSy
BTMgruOT6Lc+DwKuaCqk4QgWbCOPf8iFqtwPL8lRtOeTtI6NO220WJ3AmrCi
bZawrwDqxz3/saWaB3uPcviv8TUbfZ81Gy4UtXzJD7Qg4ClLNn/s1JVPk8ec
/gENAfFeO6gXx0+mVeWQml6JIUIOkwtdNwXaVGBW8JCi05UrnxsEJ1m4aX/F
0ZLu8wra32VlUD18l8zMR/C+vCNhy/rFDliEE8wiJH61luQSF0hS/zuqref+
++ETAK22FLM/pea4gpsEWxXM/VGiTP6NLrpXbsLaH6Nhi+FKj1sRgiNXXpJy
AcPuXlryJ+PD2R2x0cvyNGDD9PeT/ijaFVlqFF3DamdfOFwul1VMxNFrNVd7
4lOzO5cA/5EOvtxezUKjp7AelTxQMlLqsv35oSvi1IbQD/wDMs/1pxptqXyZ
vgp8JwMxpm5H0jGUaYyiuGSGp/RyhiZoE/mSW6mr2suWmd034vFLrAOmkzQp
1DOJ8lXtf9FrIOmzeZ/eVeyHnXm4YRVKJFWgy/0Zb8TtMoaWcK6d7V1DX0MN
s7AkSe74EjuLyjLPOqb8tLwLDjPgCh8Zt+y/RwId52pG/AAAV53+kGafSAGP
65qG3A1Q1CkyOjQSAFljUFZB6Y96yN+q+WbCHvHtBJNaUsOJaBVH7H0AC7FD
TTLwzCyenJSSCgG+nTsLm1ybNCkhdeoufKWu92MKepsygklbl9a1RXiOrolC
YnPX6rKNpGtL95Q20Z+XHBSEOv4gQXccf/kggBa22ttu7xFtWnJhjrGDs3/p
7eMSYYhPctHjrZfxLb5NpDkaflkx2fUmQRbxAY8c/Ci1WtIYk7MU5l3wCYmc
N8v3jrHjzDTg23Ig5PnfPDQ9ytaBRkHCViu7+AnxZSkHfTofFYzRmpzLlOGk
B9bBR9j0bXAWevvJhGQGDb/aT2XgUkkdIO9J4JAQtF0ANeclUBLoc0Tgn2pR
glmhVz805SRvphVyYg0N5kSkZtNI8v3KCShs2PfJk4BS/8CBBc9H2DfdG64E
6Q9Vcohbv6ndIcz41ouss9B8ZtVvZuCq611O/g+GzS4x/Ag3+g5mUIQD7lhd
vuG8eCIbgMsd+xTQGrRCInPTAXspD3pXXuGZHaZ695GBcY12l5eqT8O6oF1j
ZmKjUtPm/i6sOQANVItO9eELzn7JUltw4soq7GqJl3X9eB1aNRTgE7qc1ROW
RcrE/tM4ZGMI69BSJoSPKBJOw3kv2UNlIA5y7aa0XSH6+hVlYa7l4kMahLeO
pusuOPNp3VrTs3GXt5AV79xJRSzggOl2sDK7Yd6PdsT6fouuVqP+cF3ufvyN
De2S7FsDWXOuQ7jHNIs8mOm3GPL45jfn44pXUcVeNHyffufkTmGOX28Ld0ZX
gmJs6ZOgYhRyO7GcZD1lRzFE7thWsiHFmMcgpNdr//GIxrOtRBBRJsUswE9N
wKSfO/xr7fgf67zycXDpWYOqhhsuyhVarrwawXnVpfaN2ck1k8IqDITmf0/p
mRsnMs1BzV7ZTBHhMTVB3hvzJvkK9wsUlIC7p8Z18ylO4tUuuWvanH9VT5aT
y5anezaOPhImnkHHaFKLAdXR/gbu+1RbVqKl5caPUvdciQlHB+uBoczXZcfR
uCajPdIrJIhH/2H6aA9eRIxnCT3KIp0aK4sjf+eh+whfgOFodZ4n3v3euhre
zmYzODIS0LmJ8fKS6Bi8ehBSu1HJ5ll/bKxYA13HHGhe9TApCefNHyuCoOYx
IHR8ku2gB63g5aHGZ8jV6Ne6zku/eQsnETRBpyev6TO2iN3eIDIFAJJmGc5h
rgBTVyH6Gsj1ZXymRr/Yk6PATLnahoCQj+yKo1gee6QPYvvzXN9gG/XZsyvP
2GzW+W0S5uyw2GVF8MwtGmBI+7Ju0lbhsOYrKpVwnqr9OSulSXU2VdbDX+7U
oWXHf6IO3Heqgqai/mI/WkNWaPLGu0YNVQoMdU+EbCnAVCUNxEVcr6ArbXu2
s0iHpD5bNdT/jDSk1aa5Jps/ZA9coKXMF+jy6+6m6sVQSb+uwUL8Tu0DmBT6
nVy9VRmt/kidOF42n4PJ7a9aA6jUjj/MM173eJuSF8rv7jqjaDe96BgAhBrS
4y4fsDKL+mw3BmB/p/I9WM9D6i3i3Od+ReNsLO9MTjliwU1iAh9mNT04lkI9
2y7wvb071A8SuaJboIRXkDRON5xaed0UyujJg57p43IFDu+A8h4ABf3Qqnzn
nSoVdYbRPx+ATD6X5C7JaG+iMUUmvyA7vSrZRun4vpSNsOvABPRiV2MoqHiC
J8AVmlgo5N8BlRUWVuo6e+9YRe8+LDDI2X6l99ez4KBb4Wv/oeN1rR2k5nEw
B4LLrv2zFBUomufPTIsZJZs8RTEHjzhNq+Gp1cDMVp1mPF+sYK+2m5UI/vV0
td+NadH5Io6pdLvkfSNmZAdn3DZdT4OLTeiSnu5iN1XqZzVcxTijrgN2yKcP
LdEOwUGag96YO8zvKIRvetB85eFJ+QSOhQo/nkwQUq4fefuJV4nO14IL6zCh
JEsU0G1KoNKtJCgha11nvHAN1AYhJW01D/JvKr/wDyIZCvP37wsdWKBCOpqg
ekkobIRSZz/lhttjl7u9hDwQ09RSGjqMmad8bDQBr+Eg3OZ5uN8QmBi0Pk/Z
mZ34WBjU4p6Brnlfkfxt4Ar5bv8re6ujLpcjWFYHy4WsaxCklEr6IurqCGUf
2b/PbKwMJy7MM3prjTK91Qcb8+lhBYVKTd7bKDCnB6g8YIVimuZkydUX4LNX
wx9yGbCJhtnO8/Xk3iPQGleSqhM7pZ7vFfGQFSNWYbfTMGDcp+agPNhuNpUm
kn0oz1wn+SL4bBGHkSUuALLgMRaXVJrYZ2KV5guxJZJ1DFZW17OYqvyRNOvf
FHTkkPQskth27/gwcnjt8yEJpvQCms0foNJYdrqzHuylnspXPgkYe4mr0BB1
qdilJAOa/jWTCEJamAUjdcmxEz5yR5FdDq6lqVNgmNN60cz/S7crIMboJKPH
RX0ldbpBE+i+bK9V3Z7qBUDg1rJQUibrh8C7qIFvgG8fMttq9M94KDtB9Olg
a3mcx9hMcRRyUjfEOcfgVoaaVJmUaC9rU7VtOjQqpQmCjQYZbybDE3UuJZMR
ephXrMcbFdge+IWYocgSjEOP7oQydxSR81HJWEzzZ8PSbzthY7CJvzxAqtIQ
EDH5KCj5ERd2GyL1e0Ersldf4gocNBdsGZvzaR98FSCIJJO2jd83l00gw45Y
2NB9zOAYqp7x+JYLTV9jCRkw9B3jsioLUZ1eMAEQtid7pKQaEoTYdAIAN5F4
hYcHglKR+rMDkJ50MSjxrpmAogmUO1ebMKExD7oLL8O8DQ3DgdBYHVgcX0sN
TZmVkJdzToPTfQNCFgCnS2AMTfDqRBoS6IbcWZ+H7n70PHFc5bPJyZevzJ24
o2BMGsBPiLfEfzG+yLe8L72e3uiHkdhNHJYOHMGtmdOn8VmfE3JM2oDK0dlO
huVYKXZkDocSLqv/wTYvgoQtYJTPkKqbFuzaMvGw1WWzp6ttQ9ElQl6bPPM5
IUb3vePircxM9dJ3OZa3qSIItNwuBUTNoqurTFCI8AN4oSlpZh7eanF7za1+
ZkT8mNPwSa4gNdusNrpZkcABedi+4Go7YnZUrE1LIMuEO4ddnU2eu9u19gqo
bQltXO6IqLPddtLLd6OfghE1D7TyorW4KhUXm41Pq34zSQr7QHmOHGglcE4Y
QZHyfulrVrGKUv26fjInjH7ijglxS1vkf4GICBIis1AXxpR2otNz+ySZGm8/
oht9DHdzp7qSWYYoeEkD2+zWOofJv+GmSvYnmp9AWyS1ytGcne2SveQLgB7A
EOTABNNFcwzLFaiYCwWhr4AF089cXsbzxkF4x70G0qC0znTsznC7SQswP1/f
EeQf2QMtONKmsPkVreEn4sKaL29CnYEe0yA7EKRyMK3tjr2/4cm+bnPmX74E
4nbJFKmyAikYIgXQE8OrVitt+pKQCJL6wf6E9a1M6y/ePFikNSWNXV7FaXDZ
zxP5ewoDkrzmoNcYREWyOobByTxm/2OC7CKkpn6/A1RvS/xPEUE0e0jjhX6J
vyMYuQ33tHdgyBJFUe9JknZfHzKar9Vd3V1xktYg4A/8xteDkPbXT+/qlOGQ
IONSckdK0q3kA4jEVkn78AWAwhbLBPQ1BXTalDvWiASTT/ecAoPTsxmoT5og
Cjn/zz6O3vREPVM9JQUZuUHsxBZ2tlUiLpfRsSpb9SRt8dWSsuRuxxSsCenx
5dh7YAqu8OnQ5Ve0Dtcg4w3Kou9pXGUga3CX2nMMlvfB1JXWjIl5tR07KfdZ
QIsaGchDmRHFIolsTnq0KnIjHXxi2P+bPKoIjxIhokEHbNxs+ccuWIV3eQhE
NrYssnVAtsG/ZGlDYVa2zYQcz6f1Ezad2Ph0slzjp8NAh4khv3W27Cpx18u7
mr/dI/3xhGWWU5gIOy2tpzGtt5QRX1xLlgfQBkmffpedAOwEAUrph/ftXgVR
Mjh0Mz74BXc8At5+wGbxf2EC28WJxa4tM8h6U3scVG1C/VLufQYWWzSsGWsN
hPt1DGHhXmwkGifG2WzPnr+gzVliKqbj3aIBcRZCoIo6adVrVVmcyTqnFLGo
v1eFEypRel1Wy/W3Abiuw3fjzHMV/SmpDHjul9VfTLUqGnLxwcGNz/g0MaIk
ZbVx7LUylL0WjcaJYlwfGVFHAXK5KXSYI+AHIJVBLvbPTR5eZrjfHbsEs2H6
RFnRzSmmfJR0wNgEQWZkSRVjJ0OOuCbmIDQIfChvcVpbYpIePPTwItJOJpym
H2fjSB2ihzFTVzDvoSo/bwGKHDzALHJREhRLSMIbQ2ygqrdxEMfxeO36y6Ax
oQLaIb+/nIiByHFTiD5EjMR+V76vZkG9wfWxyl7F8iXPrhZKwSZ01YvwYE9t
bpfbbPKeBClukUvy/ACWnHhTn26oviMcIGiolNkobrUk7a3aOxkkSisXDZbd
S9q9egRqOJjqP2L0YJe5MDrh8Ps2vocUYerwp63+1189gFAitnPMTdxXMIwk
NBdSR7J5WDXDQCmm1f9tJJND3IHzAeDGHAIwxcOQdTBGONNU2HzQ49EwAWUw
TU1XPQAIIsS0jw6p7XmC1rENePVqRnPCSzfHf0qnOUNyeYJ/7sunuj/yVl+h
Pvo45Mk3LrL8ztIsp5PiEnphnIzfcGxOJSXAJ7ovrESJhmncvD41+bInDJPq
arOOY0uTTNqBAqqR1cp0qVwoivc8ECFWR1iRk8YFx2hK4l64oLteH2L4AYzM
i9Fc5KkwvsSrG0pOvahoS3vw51523lSDn4V60d92aDdbBhvbP51n7UoRxZ39
naI13ZoHurMfFSxkNHVScgE5TyuKtV6ckw6Znv8QIeOErCEHK6FRioS+Q6NY
hWLCnHkK7Rq3pEwn0Fwwmd5j2AAPjWCIj/mPs+1QUOazp0GGh/4cBG2VlgrG
m3SyzPczJ+BPkbGJhF2Ljc0ElQJLPvDBmqsp+od4DhEs7sn4O9ncKjl6sya5
Jvijn+UTtEVtLMyx2BfncPlTN1ILG4RNReu5nepMpj4Du5qxaKuAKR9xrqM2
zvVDAHFQESnUuOqUe4QKelwiscr5/85JbFQ6RlshBGfRvYHEStknru2Lsmon
Vi6ceBtkRjs5XfkvLsdsUY8oDC8kl36wbu8NaxSYYQtA/XeS6x7EUU0WTxLI
TqexIT0MyQH8eA9z/hKqOnu9TQO5hlLrAN6VyHqHW8CFSYaxjwSjU6r2OeLd
SYSqtxS5pOz+ybM9wAEpwkvZtwY5lvxb0CmHjjDvxbZZ++dLJRAA9YG/krhr
RX70ZaD0YexihEliC+Oh1GOirKMtI2QDRNCo+p0Z31bntwWW5dFyEBz0CH/1
avGMoxRZaMviUvpyYhfOP+uk64IcAyoxDjQU0bnyL9tc+g5HvaM1ZqFAKMLm
hquk8mkLThVXlS/rqFxQKuF4RJh8X8ifuc0Do7hu5wLHvbZ6gU3O11PkVrtw
jt9RiNEuqENazVusspy0CRCGvAYsFzyuNgvNsNyg7EfPYdDZXolqc35tVdls
TWhVpEy4r5NyQ7xcdwTIW2b+nKP/wwAZxYcMw/1/tP8vfA9JLXiG7EfHBJZy
mqo78v8hAKfFs9tCwZBc3fJwSbKniTy2PUJTS5YuwE6vJS/VbJvs+4Pwsoxe
8pprPzaIedck7B274mUYBJcp+PsEALnl9ZTuYWltuEuC6jSPIc06IKLT68kY
M6q3z6X1DG644hgAWR1XUTPFp4EyiExcYX3pa6QHsegcAjYsB5TlJiHm6Qh+
oU9DOOo1AApnYrxbxKo+pkIkTMPYRPXvqLLy5hjY34CHhAUBdPEFkluZuj1o
ydyLzU99vsIWOQQ9GXaj7bU5ePVbOWJR2BavaZ0GrhmyEN3sj5NyTaDAU73M
aU8e5gOQuqRrCbo4y+rFKRDRchJjJlQ9km6DUzRVAV0nj5odASsGbNBigrec
dcT5l2KcVBkOZz4NixvNf6Gejk0SiOpJ6x0C1ijHdUwnwwDYArMGtakrzWcC
cC8xyra3HYxMLr7ntGOgoLq58SNImSUyuCMMD85UcsXwLfGU6vDYZWlpiaZQ
khTR6T2QrpzX/D2nVZKCe9rNVZxtkkssBFATP6WWzInoFOStRxM+jEmabp9x
iAcouT6pH/IQC4PVoce8Wr3FByXLnm623KYXXqDOnf+h9gvZEDHwqK1FUcZV
2W++vxS6g1l+9uRUgo7U1cyKYDaYPk3Nf77/zdRPFuDgl30lvM7gjfVd7Iea
RQTmbcEP1PwBZ1UPEfsOCa3nQZF1CURUL5PdBvi+mT5zwgLbQ8oX0XzzrrRU
buVdczAZzhZAr/TZmrfuY0g6XtoFvM5o4VkXACkT3btMuQnet8DzrHSaYYBi
DlgTgRM1CFZfVFpZkjMqpH5buteOJ0HPdGqo11yj7SSkKsxgpyYo5x8ngExa
64HOmfdK/Rc2iSOBuYS1DNipwDXylShPw+NiDHlsmjDzHIKq4jHBDGWvbIar
9jjeLPuofotjSKTaRNZCvmejMV1YgcW8cpCUPfUZMHQ4Fhm3WCa3n0F5RosE
2oQIDal4BCipI07R6GKyhCMO1iRckz4V6Rr01y1R5H6U78LoFXNa3qLYvvWs
/2fGrdm3YbUiDuW0Sul88i9X+kTlgU+GgwAKyRYdD4SOE3UeIwiiXoPU9qY6
5FGo6csPVchMDTuhh8qXi/KpLj3Uchjc/XmSbkULm7mM1M1HmtBO7YU11r+p
C8OYBQbFeqeNlxljAZqzSMTEagcCVtDBrp5zdt1LAA3DJ1dvGvMMcVMEABCR
Wxmjy+R4i4hmoAXhjeY2G1pqmyolGSOdVhejjFj6CP8Z85zjaPSZnNUEgEPp
AG4jnsTWzDR3DtVYqgzhhHIoviFMZSyqtKYgWhYI/NM4GC6nxyFxep6HY38R
7k2xXrSOk8KJIu6Hj7IB8EpakG+0MK1Qa/gx6qRzoWRcxsG1umqw4RbIQLfW
AmUiHFiyvHgknXUYG7VooVWZktwZuOM6Z9EFRNMjGRPSVWu971scNzYe6eQR
1YxribjtCna0k1WyHVOOPibSGD1IEubCO1yVoukJS3Yihh7n3Vqlk9N4vsLK
6W5DStTyWjMnfe2N0NAYh5Ay5KK3n25HR/Q+TrHzOmkr7Ts30N2LoDOSI1zm
W98K1ho6OaAzMdVHTMnqp7Qo3gXw8BFGWEnfFp9w6rDo67jbPASI6AuL1OCu
CB6TEIQaIA2WkEhEijHdu53KIQQ6ndAZWSP8CI3hK1KeoOxfzuq+vgaJRuef
7n0mTh+DpCyEcGAdduSlSMWBXYcuaUCsRjHRL0u+cOeI+jutP9fqL6skF8p0
58laqo89vvufBCRUHIndr/daTH8QVPC4svUkRQuPt0R3hLQ0rwOh/r7r1vyY
6AoOZ5sK0bILGD7AHz/TWiFVEJV0Q1D2gJC+ICqoRHoaDlLlhEbymq6829JD
o4tn6aiXM3BhMor/depl5paqUuQYOzdJW/nxG3MzOhZ6Y3WqkBLK0YVt+pls
nF+BoQ0d04BivcY37cFN9a04469olgx0UUl2QjjJCSQFd5rvZGBAlKCeJ5Ig
a0F45Amn/Us0xKOMgjZoswL6MmnssfyWLZsjcxPEyt/P3l0j/zcbC2GvIgcg
2cUfZ14afW8L//qzAbOAL3XeM48iX9MvCPcm6o3xpqDmNxksnkD0oYhBOjMv
paI/pCtfRMG/z7fWT4jfhJfVGnEsQ5pTdBn5dZ1evJQARH8nouH9Q9HntCnX
Jk2qpfRsOAgABA0x01deKFo6wiH+UXCiKK+90p+hc1bRIX/+gmaHj0Q5QdiL
3lfwFHiM99U/B95JXFkbjVFMVBX4scmpflSWHY0M/LOIHez9RIM35bYCt4Uc
zhLlGbvfDQjRCbe3gte01kMwtlrpDl0kBFD3Y8lgA88kg2eyyuiTDFeJkOv+
NaWPXdMeZQgFmsv9j7Eehnf4YN7zpqx/rLly8aA+03mIGY5ZN5Sk7VckVyib
1oJWtE0VDh7/10cadVUlhMET4Vdb4UXGGOS5iaTK00I8G41JigZkmi0KUpmN
S6JBVyLQFr7pCKynC0Ngxxqe7/vMEBAeKLrdt6Qg0b9r9VoF3Up2tNQTwgzw
DmPuuzoAxtV5WJPakqkYCjdRQDoQkfUq1n42xJSwffIQjzLeDpUqBX9emXjp
WDqn2cBpMdpUsinWcC4Qomn/n/psCtcfhanmzblo/XedoavtxWsUum9yhidt
ym60iEKsJe/9HHkQZADv1h3cNdoZZY2q85Z7WrEspOZxAkiKs4KT7dXfV18K
sEci+XXKje8+rkZItCsVM6VEm+rq6Tsd59hQ5XKHVFAwXExjJc2RHXPROx/e
pVuIzhTOLRHACZ6bd+7y9gRnC9yc5wxDZgcB5EEkazbFs0r+h0aAxfHqsDO/
sPshPNR7v6iuhBalYHk3EynFqRK8Y2DZR2yY0uoFUk8MBdsHjsXhRIh5l3OB
N8NcQf2jKAQtMHrF6VlAIkOZumIqmtjyrnk3rGdfpyjusFEAulznIQAXTpio
XHWq1TW2Xl5Z8y3mzKDcNuilNXgBJ/UFew6AMN23jdcQsFwRa7EBsVuxo/6o
J9DlQHuvkrFXdoWXXMB7A1rdXYkygy2co+v29ipxqMF3BYhm6cuK8qxV8C07
TzQs4DDuezlNY/QF9zsrVqGhq2LdKbGwRo9R4nmdK1q3yBw5qERr37vdCYo4
ZVN2v4Xkz25HdSsfJqcW6SERORqAv4tJlgg6f/1v+x12UrjZxCleF7ae0aMH
5y8nSIQunqgdX98qFISi5xZo3akc/YX/2fy2qLWUTbH9q+Co6Oj3ZhLooduS
QITtbA3cGdKqRcpyWUsimyfnIiQgBvOUKmeI8PRv6HTvisgCPULyVTdGTvHK
65bbZuM3/Hwqiue0Y6/dnsa363baUngtI2u2n4g1Pe0d0ITR27ybtwVvALai
P7K4jyE82S/h27TZqBSRaJ4QSoSHZx4s+01AGfu85a+2fh4nkQM4i/jB8mJE
nSHNIKRXzJW4OkYPJ2JyzdvlQCB623s9AWlpz3DhStvVCu+8XxqfekVqcCfD
CUSXIcI7x8odRDpQLVIMRarMsKdGn5d799TAi7E/XOkkjeVJ9eRy4rB8dBq2
eq5Qt4zFsCXo4qkQ2xvj2wJyJpZBvX3UEJpGwBnO16PKWOASlk0ZUkjqlG2H
xbCR9WZ+udka6Cr32XfhiDGlrLnatlTnHyyYrxWG7LwTBrS/GvoY+XEr4EGk
uhxEILcL+Y+s3Lo7QXQ/Ho5hi8FMsiBRRrTGmzlHdzbzwM/qSY+tOw/puDy2
d8R6fm/KSuT5e4ke8vxU0Nh9/rkg9IeJG92plci6QLkpaa6WTkia7GIOUi8J
AxSIWXPbBke6J2sFJH9ERPpCCB5eG/OMPzXUZA2d8qlJpDQHqBt4h0yMM5Bg
NZ972yzWLEB12jgesCUPAWKSIX/U77rbRzoO4xp+5jeG2+83RDtIFY0LC3Pf
BYqC5ndTQlUg8vdXEzLBUTsFfw46tpH8jlVztg5liu7xnTnI10omJjm7jXDw
TuYrA+w3DBEuA6uiq33Cr2vCReKCR0AkqxI/UxRrU9T2rjsqAwYQByk1ImDJ
b0xiz0hzx4woh8xMUXYUbJarRC7o9SK6A1pTJYaSBEf2FskkyRif/PkB9831
e22VZ+aCgLHCTAd2POe3gizWzJ6r9ZpVbOrsl1jOfaB0GmdJ9v5P0OGfU5FQ
hyVdwBANj6XvXxyYugndhQbEXH0vQnsv53whGxSg6MyK6T1A8AWwse0vUpvr
w8BoiHg1yimQD32QwKQeosr9j9e4jkW2i3YtdTmELI4E21r02B0fHiK6MFhl
mo4+di/9h9LA3XMm13Lem7iBcmRCYWWOH50DeSgnvrgyz+oy76Gq4YBRBSvc
yCNWFwjtUPcrORSE730JzfBqpYuTMxQsDx2fPScTLKhpjOu2tKDJI8XrBalj
DnZoX4YvJFUWs2sLh+iUfp09oj1W1j1pqeVh1fFhxPbpoab1hxjjZ8oJvmW7
CMXYSh3BV3tA4m4F7OIRoAiiSd5sP9fF6huCoX2jqZDYeDRmkY5aPKn912BR
8VNm5FOyk9hPwowdo+2ZrnWcLoamDg71/K0oy/7OXxKL0C9oGxmn+tyExDPt
NpXGhM445d9noIAE8JADQToUD6guhtKl4vZQD02yqYm/ER+N6DZlPG/a9jgB
A/PeZaihs+77FLfZh9s0aj3BdYLQMwzdAmtuBmepUrDEsHQyeJWK0usD+eBT
yW27YZ70owsV2bnPBh/XOG+kUjgFTbTBZ/IT79Gm6FAIS1hKd/qg5/hWC4n4
Oy+AnWJvi7HzldLfzGBAfdvSx9ctheqK0bY6YzaNVDlYKA8x5F5tb6nJxeDJ
dd1O32E4n6HEFDUBaW39p8t3sPTh6KIPSN5QWNWzssE8TlfnGfKePvTbGJK2
AlagRRSldnvVatmYR68uSdov0F53VYJyfn/7gQJkWLyfag8ubrk1gMuag8iJ
Dh4FGjYkNdYEIkYUZBFAuKYgPzYqfA2/NtpStR+lI0r6kWarWR+ACdFQKMjq
NsyTZUYrGomjlWZboFBjlLMrIRKMUoq70A85Eoh2mlSryKfNOJIh+ktUvIN8
vr/9jstEOBmE3gkDyIFCcltUvBxcM3X7Q6txHLNQAcRjrR9F34kFsIK+SD9J
b3Oxwt+nh2M0ZifBykoddxedVIex46rmeA+gpdeNNdqfIyWUCHX8qtNIj/An
krlNkRjx09U/vdPLSFM3XbuhZ5v3kl347ZjCA54VNkqWzDTNKqoskCtlXtu9
BY4L3C7TOEPHfSxpTL6bin3DL5r1ssfgQSKbu/LsFnDPwsi/s5SNIRgVqdRy
cZ82NK5tP0fZG5r3q4hjlXpQFPWxfr/VtxE73+5TOj5LcU3KWHv/vzZx3q6k
L2pm5Hq7up7TjqQM+sg0PhEe2EN4fYtjSB1d21EvjH2xmsWiWV6iOvrnomqc
EY0S13OKXRofN4icSDEOAP2dRRFkTi8hwg82jndlY4nTzLBl98dI/my5ngs8
k31TMcVbExpb+8copf6xuBNVePvERzoax/vqsstIFfxUVLaGJrtvgyH21cU0
yEkjGjgFlCm4PZKbo0oNE2KBcxJA50UZJyxRMxCo9RU5CAE9e/eZhy8J7nlP
z9ZRQ53Tr4V2HBVq1RkoXNrNh4mwKYZh9hmb9bSak+IzeLYSL56m+RB9NuPG
PTAU1BRuEgRQQfNo9CiGxreNp+5n9hb4OYiNsiveG0vC13s7e8ISS86tJ4BB
kDqTih86BACcpgj6MPeDx0lRLdCFgHvBrSDRxPyJbkY9/GJ4Zmt9DCRBDIn+
8uLsWsfaDdRPwlapvKTdddLsvYTAy+Xk8/MrA/2ovBWl7U3WjyReVa8OsEJc
UeqtmuWoTlu/7f1q7XaJzTJ8YUtydU59CiUawvUVbp4FII9Hgcql4jhNlueV
I6i0boQdjPFO7Oo1uP6TyLMlhKX4gJdky2CLGS0phIgYTsZJrERMhKnyr36B
0LlJGU1LqXtvje6uv78xnyzpos0UnChEFcwYHV4QLQEYgoymUgFsmmvY99wU
BJVPzuGFHTreP89wfkRnZBc9kxDaaKfu/ijbt3Zvgpn1hTxhPNCNEj6MqMpE
08o/RnsIDBpgyMrnuNtRGzlDpgCqJl0HAJD8FotGk5CcRyhS6SvJ0JPz4/vM
qM7+3YI2JLodX//Pf5x+9AFQb3fjUSzHlloB+oUWmmPwEXSr/BENl3dzOQY+
yr+lV81bF2odjFTeUWxqYy5GHvVU+1rf8n/tOKiLMeA7MPxvjYGRqceaQ3hl
fqejwIc5fYMFhRG5G9ngOPz5okZx+3EnGk9u3p7Xh0gyylgY+iv0GxVOo71X
sr5SO8kW4wutuHQtO/qI2sgnhcCz6yRdqkzKsXRksRLQOIod5Y6HdNLXCqBP
kPcXQVzwHkBfqFIOpT6+lUtqcgau6bXyN4AlIFDcCKIK51NRE/zuu0AfOZAS
R/R3k8FKHjLxgI/M7gaClJ2VXTR5qlpnXuoLqCX7XogWqEhVElhChyRahIxM
Psu4BEqICV/2Ed76/SGDZEdOzJV2DS79eDdskiubTp8g5bVFVEMZxVC4XdfW
xu3eZ4iJSjdqp9k9PQVfWu99E1u+FOBUTCoeiIQkKWirgnbnXugs2IJNa5dG
Uc9s9mh1Or+Tp/3QlAy/I5FH43TySw4KkPpofgDA7S3OptjX0LMD7sqkzkH+
F8M53Ltwqkz0gNAVywrhUC6hZwT2rwaQPT/hQe9E4pZfUCQYvHH1JN8Yc8tm
NTYfVdZ8KD7Iw76e4q4+ym708eoedhdQtRbrsC1uzROvr8D7hjIe/Zn+GL1Y
oaDtFqL+ytFxFjB81d91oHIgHDOd/dwnYHkj+Gxyez2144oeczfvjhx775gR
4iAyl/Ezro2JYsfEqLih77flp1lBrNt8suV0t6Mveo6b+iw45YOrSpTOLq9A
AYuMqSU4XIYDmlCvthuRsET1W8DD4yc+E6I7f50C3Y53mBng3Ek+ZM/GXH4t
549VwRmy0TUfzhEbKAouPZz233HTwkOwipD1yHQf3KbWZ3dhueDHEccZEtWz
fLIaeLmUDjKnLWHiI7XtssD45+60iObFTmLXIYhssHND15vceLyCm9TlTpkl
33Y1OgnG0V+LUEYGTgZFOeJoz0rp1IoyM3bmN17ll1tJXxix63P0BAvbWPie
9LRYTzaHAOmS8MjCD5x0jPXogP3GSndBWjOMe137VxZ86inuHQW487L7WKWJ
i94365FKR+eMM0F7mVExRin5mWbL5ajxle1O6xd07orv1Jw8ihkHYUUumUJ5
Tad+bcBYK2+p4ERv7YJVU40JArQBZpu5cDT4CmmHFamFAnHyUuTBQvm9NXZW
yKx6MCMUM1+YTZ9RfH3Ih0cAC7BoQoTlP9kfU1LziplqoLc87eO2qdexEsfU
UH02iYzIreRjnJ2VW4pD5wov4aEVXnFfXRVZ3HKwd/Q17OXQX6rQFVx4H77r
NKOXtoqfgA1WTxIqN5eyyIUdhWm4XTJ9aDLaOas/rlvyX5CY2JxqqJU3H0AM
Tb4piRRGuuUhmX7l/lAb/h21ZX8t/HPoi49pbkAwYINmzGVqwX4soIGFX3Y8
/cOXNFQlxv8iRtDe94+mCqfTz762OD+TIvG2UKbdn1kLm8G7oO+lb2pT8BZq
+5PtFb0l5fJtmGEjiiXpBado8aipOmU8zXqsBXJwgV/bKRNxjx/aR+9umRzB
pwhcSZbeJs8OKJtPZjtB6rTt9ByFPpgF8UThinX92S7UjDujsuApiczolxgi
bOYyhFBYlmwo8iezoz7KzT+P/Z6kBYbkrK8bFfSVYlCrL/2ruYVW7ALyE/YI
ZhUC9YCvDhIUsPa9pxwFEi5cwst32F3wscT3j7r5aktWsTvJglmf8kQtzQtw
W0T0MqMOUMBrDdwtZCt1QsoMqJHtLNZbBrudHiJfBXJiaiGDwOz4DtIzOvLe
BmuY5lNnuUZHB/U8qSFF9B2Gz9La+tBNyCwXCG66JhN1sp3bPP7MDpENXXZ1
xX3TjHMN+JMWJtbUicr8x+9tp3awL1SElVDwDxbnQEkGoHAdv3qYG54tce35
+xOrx4CjO4EH1H7YMsYS1IFT896iiJjHMj11BEopxmDe26pnWaPskVfySfpD
kQbpN0jHOtObaTBCen9x0XL7or+XV2qoMxbtRs1yC3aQfZESQkYxFsqRmgwO
INWQy5gJ7kLo8g1lg6CYThjz1ONG8h8sdcHAdY2vGzwz6nfBgUAUgv/Bz+hA
QEo8e92Lw3Xkyu6NNDCR8ID1KKgYQQ8Bg9nCIiyTkVE152hesp/aOUl2qM55
Yxh+rCMUGd+7KBcK9MFD7LVfyMwaWs/67gEmPDQrcKaWfYfiPVZrP/YtHTHe
M/OwyjRnibogImoZCVQ3Py3jxzbicT+bIty9p0SXk8tropflKwo8LLk30QES
7DLpJZMEvFyMirQiR/DGd2rogGAOeRVVMEhL9YSmyhvAv6NOSJ9DzEP/+e0i
ZxTi/sgceijITagCWwTkV7i+j8tlk+vuChZrn0OoX2KdY2nhcTe1hpYKHg8l
ShvQwdA+9VwXhNjgPid+GlXnXTvRJUQ/8qIYwgdq29yv5PovDXkff5CLdO6b
PAY3oIE5OdcRcz/ORV5NMrOnswgMyd9SxO5v4UANZOQTHYCKVHmWmubq6Ryb
SJMhqAW1FSgQk+FM5+9vIa9gJV//ubOuBIfy+OqhDVnSXJclyms+ZesGX9n9
vc9SjwVFUJc1X7Fe5nakVlFtO7geW+0Ksa6AZKNTlI28HmogzBV95NR3sJbr
7QGsyOBwVpkbXeHaX29WsUHgeMmW06khBgbc2EV6SkFLCQ77wcR57ULoIBXT
HY9V4rS7SiQacmN9Enq7lz/UiU78+j8QSqm3nONVUdaAkT/SVBg3jM3RTH/D
tSKqeH+e6Ezt5wLlsjsL/sEfaJimYDxoeeWLiRWmAiU1WQbkkMwCFZ5RoJKz
fLiY8HDyFqcg5Gk4WIIvo8JSSmzTxjZRYoqGO5sumdT+FHp6Yw6JlZjpyoNh
Gehyx3Mlr2D5IPpGUDlOJAL4PkdnwHBrE6d/Hg2tY9nMC7SJejpdvAeDqlGx
m2BYn8J5aqogK/V6eI0B74xBJVgV/EXGP+ajVAXiQCQ2p+lHJHKY1yoqLlcy
pXQ8/R5AwiqelxJtp37QhY4ZCCeSig/zzIxojTIKUyv5w9uzqY3e8KvkO/kv
uIqgISyA9S3bTkUPLN8GONzw0Cb/ObibDM5nNzA35e6xyGI+HZuimBnR5jnP
HMlsS8cOrGlYICzEfoY3JX/5Id2xmOHqypLikEpohBmQ5s8UrKYpSLvPK+oH
znAGKIP8zir8lpDG0SGAyhNkrBKui0rjx3q4Mqxgpip3tKPUnElDCvoO+LTH
JapeRyFTnG4nhbOFYB/L4lvi/OeMvK7bBdud4FC8CqPEKYSZ9qMfBUXBQxJD
zYPk4ywkNgSezN+JDRkwM6ifPFIRnfPWLBxgNeMa2NPTBYvU/aZ+qiw3a2oJ
TyjMAtp3OwbKvP41j+1aw08Eknkp5B5ZgSa8ZopBIMGkFuy7FOy6NxY55CQw
15mUOuUjUBNuWSs9EheVtlc4+PumyDZ7/6XzPHUWy8DJDTtRuH807NEqBELE
zy/M/T6WX8r1QlwBEHhjbuqKDYqEqq1TUyCphiP5HdTxilsNFQsHYOzeLFiz
dyVRdsgDVLkcJWUB3707+XVOFJsuBjeGmmzSVFsVxfI8g+prS6qQ5ddWbg9i
Oz9H3q5PjqDjyTGn7hB+qbbT1p5u+IlCJNNccF6vWyQu5PTDf/PYGLjZWzPc
slYu6JXyTazjlBzMCmRlcz0crI64F9qpB2Owf9PJyDHKWVhdRyw2ptEKaAYi
nQbkGmPp9E28E1ox4EktrKQfJVPeTrjn73C04/BvUnWawUV26cMKAH8E43j3
qFxH8rZ5FblncZJleBKF7XKsKoFT26cwIVA+97KN0rezJZ8uMbuexqk9DCTa
qWOVNV3uTFxLu+pB8K4Jx014vZf6+jf4NIV4Kkw9MroOuH+mSub6xFLfluaB
QBvAL3cipbfFZA5q5xYmuE6rDkByRsHnEsDMgPtYYin4fw21+KTu951NG9HP
oUtQfyY0073ESTWgCTLfSOsJuRn3wrtZ9biCr3q6/xrn+zuiW5nvjbDGoVwT
Cmoiz6rucdzquzLhCTVlRDQdEqNAEU6BT+DCMEBMsH2Lu+xAhEcTA57FDt6n
AdrEtFFERCriUKxChjBMcZD/JuQ/BigGyBvkqpc9P01g1ju/+yhlBZjijN+Z
QaV7PG1uBEz3DQfUg/KjE4WyZH3IfQs+VqEBUs6PNecxBUnNdgnBqzt950Rf
WHffUk33r/5TqGO4ffKSC7K+C5S3qM69/+DE40DiNsxoKtQ+j4eE4lTPFCd4
HiX0ct8pibjf6fFo1cOKX+BN4IE1utVNkMrqFiME7idAANl41TJOltbQAxvx
dX+l6tOvwpfgbbhR0imYJ402rjld7Tmkiq/AjYq02dm5MJonbNG75ufuPNSR
quTxYQVj8vkRhwOL0NLKNEEZGTbGjvX/t7ol/rLg3Ad6UIvfJVMprSgmVlcg
25404g8Cj/GoumdbJGghFHT0xLbkqcADgZr/kWhcsL+b279m5wKhrQaioouN
wIDJ/5GJUNk1ij3jrg0MAJ8ahtpPnF9bymq0kmqQ99w1eH+udag00Q+HKSAF
+rhDWpIt9/5yN/HtpiWzrp8pS/ZgS256vvgsYrw1NJ40uvOFoRKJnCWU5W/p
qzjVPW5O9ZrV8PoN7UHIrSzfrdzfzKj/DPwl3Q5+7QIrdetr9uOYahFOhMzG
6mHqJOtTgeaez0SaI+Gxl8//9pViB4JvMV9UT6mmF4nYQ01UxTy1Z2pmG7aZ
i0xdrlp/TmM0ER+nef5DhOFJGhyX1vrd0hRYuDJHfHZuEpHtzzLkPfkNa4cx
TUeW1e2hmX2vRg9Hf6RY42Rx/w1Ec0Lezqtw6SEtm6hJ+mr/dpLcNsdqFOm8
LTRj+PdGiA5NeFDjqVRCDfjNfYVcKXMwmjQmFNWMVxIjqo6UFGPhax0RpI/a
raMzJA1pQI+PAEqcH/pLOkxaQssCkpBAF3TzgX9eIj2gsS4/I4QJ+EzYXkjd
BitHj0+T+JuM4ZgGn8Vy4l9I2PZtLTg9vmwRnCerem6UNsJmI1C99BemEvWY
thAcivKeKwTTxZ5uD+/QbCXqwvyKcOOe2GEe1iHuyDE+5BskgSplqMH0rIpb
Ik096T6zx1bAr26qzAYBX4RVdVkzEOaQIyG01RIGZ80IjD9LpU+1miLEeC0x
OmFiMN2urkTRWJOi57dUizH5Jgg0f0XtszsrL1XolkBEZJ78APbgcpoVjRHM
vpWH6dkZaDcnSXo6zy7i5wOxDEAvX603uThejfMRq85GBqWa2xd6nVKt4wPG
fyXQpFSyStP4hRzBJoMJg90LBtW1YLn3T+qVqcJrLDozyfbi9MnWf8gOGKeD
+oSuPtNPWLnFrimBvAAR7Ji23sBwQ4hwpVJ2hR9vJGEaI2uzu8v3AF7vpzX/
7oHx850vTT+8WFKXL6+6QhxCsF+UTGRkoZMtAJIDjgYzJEs17anG30lY75su
SdJXkl5smlwhheSdXijvs8E7HmToLWMa4UQRwebvXmf1HV5dCsYOAWpRalSN
4FH2uagxRkJ1hqGAdHoiV4kecOhCSoxMNHwQszn2BG7k7JhDK1/h5dz4WGL8
g5IRPvTebE0JBaZx5FN98A1tFkCYWWuflCrvPIN3h4PJ1hGoIpgGejnLS2mY
9oLdYq9fntDixyoyKzq+iFLy2cRwMZLeO+WaHwLyEbIIEFbzGJ+pfU/tj3E2
66Oa22d7Q6G71203lzs5oULt54/pJBlq5suMnN1cWy7ZvdP5x4DS/4o3DNkg
euPepI5ZqSjJMJWdgtH9NCpKthqbVgaVFuIjsrbqD7eHnl73tdK3hpIZ9eLM
hIcV7T0v0auLAn4smtpMfTZJjZhPCcRR6xFXuWeTj8U1EvEOwb9OC3FyaRn1
T4SRqyLSZLG3SvsoOb5z3Hks4NYOn18bKWHpiLW+VLX5J4VdGb8/rMjPy/sH
xzHfAItBNjeHmvO+G/2ubw61D/3RjcABDdWZjdMAb/nDNa0l/jFQ/nGGizLI
qRdRuGsMtL0tvyCgT0w1NGP4U/b8o2iIK7AhAMtq2uhaLbWXJ6+S2QGXWQxh
RIuarWn8qMk/WV+XOeEaBRY0W5irady5FmaaZdP5RBxfHMT+/HD9VaiTnECz
Tw2QDz/3aNjXledYIhMrPfzIbUHLGzo4IQA+uQU6Cl4nm0c0WLwhFGZWHShe
Jj/UPC7PW/n/+6/rzLJDIT+1B18JsCbzePYe6V7m6xCDf3aXwsJigM+NtJ1Y
b/1EWZs2RqeoWYDCrGwPnhqgWPJ35BrK27uW/ck3vQZTwxZnSL6stJGWEJMg
07ZUeTCjmxgFIAxIPGJkysTE9TkuTKbNUlI2TFCY/jo0mzi5wzHR60ajhIlq
Iv2y1JtP4YNCM3x63S3yK7J0Qq5qE+MUHBZUJLg+qGrrOLRTcvYxAE+zYZmh
ryhQ0zDB+qKjXnwxdpwZnaeg8isVyxWCotZIXGYjOqKecOxtPjl/xwwSZtxB
G5or4hVdVRdXRTf7QcNu2ZL6ab5b7Wb7gw3EKv12TgFkyPu88ZtVVPhQFMLa
nzhQUf6HhF0iVfnARCEKuX2AZ0BwtPFF3h/L7UPZ10h/yAhKFQtzKlAbF9cP
wQykhq9Zo0LRQs/3BjRCmfAJ5xGWQ6vZvOvHBtXoeb58lxehhFT1CKNrCOqw
DnA1QBj2+MTlJHAWl/d4XEo11CE+LgQvMBCINsrZXJF7OJqyleGIuEI0nusX
0J8Mtn3MZNMqlly8gXFf+zKXRnhZqsIVcOPMufBnhwUCDedNhUoQ9AzaYumN
HCixo1hQbnlKKP6dU7Z4a1ybdQhYpkFQS+oW+P1MYIeSalvUVjvvbZtg6Bqn
TJJ/jtMmRZziv4iN0PSNpbFIrRwSoxn9kO81a2NY4CFJt2XWhfQEPhJ6q36Z
c/Fw6NJgJUwVQxL6ZRdb2O6V3jBTgpN/Ay1ShzXSQsmRhBLC6nI9bXH7vb4N
BLdyCbCINXgW5HPTWZjA+Q9spfSPS/kzYu8zkBSfz0a+klv6z+5npUJLdBt/
JKnLvVCZqIr0b7hk46Jjb5PXVSjEqpt9tYUniriW+ubglIxV1qf2a86mu/3V
8FBV8FCOVWW8l3PAP/VDG33xTh4ox91ChUwzRyLfQEZSO8UKMQ1VvyBnqLgV
U4Tsw4cm4H15H2/0RtPPlWXDctbeYsurDAycjRcdjb0Fv4KDq99MuHJ0CriW
sOQmYvtgd+WBLQKEpk+8n7H8hgrpyopsnJH56T980mWL7SbUD1G1v3FtMc5O
RCpberYu2FztxW0ull0mLhbwqoNbEr3z+oYIiAu9nyB5pS2NWCZLQ7NEmDyM
1UGm91qVI9YiqeDbiZ6dtBKNgGLODkyB1AdsYUl44ESQ5VaSfw4ZBOU9JTVB
sF+Mz46uhMIbdQSTrJxXU44oHvFhx84KBJTMwaNFB3rjSJvWad9X0LFX9uGt
3TfofRH9ljweC3//266yrRHYTv5ndYR+Yt5oefn0RB+emg6hc4uQWPWuEkL5
reK6aUj1VIxHM/ne53vI0Pov/msYPKSQS7T8lwmahVHVzmm5J3nAGM8rLT4r
1Ai5vuvRoS8zNlLZEDZHX+y/Q0TXiaTUm/GLjZ1j+ob10RyuJqfBWVFdZsy0
FbY76QA8DFXKDuZHPMUgtfcYWK8d8ejDXV8oSYsoaGpAb3wHXVE/P24XFJqP
tOlqKe/faoGq0DStlkbjWdtDmHU0qoENYixgzy0eSEH8e+RFjxOD2+Qetue7
o5JlPs17za/D6er0b5wPsPCp8iRmRizCc0mYcUhTqkYXywjLVd+jZY0cRrIM
OLXV2ze8f6yz7yoQgPl4B3/r3JTKh8RkuxioQwy41Ya23lzz4alTLGWozCuo
ODaNpy2/R2w4XWwE9ds50KBCBYennPMWzJvcgz3cU2PfvKm637GZRuKePagf
m8WoWxLybSB9tEp9/SeqD1IEtitM3UAJexC/MFXAvqA0WCjFUKocj2ry2YFI
oZqbhu2LQOOPg8aNCf3OAJppBbezFm2LDAj5ZDGjCKuYhGc1UxZCPpMc77Jd
3IBa4gGe8/C/s0PcA3pRpHXc3FkzXe/qCnWSDUPCFGyGzXpIxa4Lkwh6a8mV
+l3IbVPlu18miv88LC3JXspvxOPc9qrpojOdMtrDG3GcUy86DqkGCQrlHdkt
M5ToKzKJfsktAAninUPY7wCZ9VDl17oDWAZMpWzk2OCoLNtRaFooHlK/PtGj
LMp5V30LBCoVpRS0R6kK6WppqKpGsoO8DaHssyPefdynhyx5L6mFHQAbUz8M
dCgMamGUh/qcXLJv4hOiI066cUBljDJtOjbU3MFDcfaGPtXVeGClJrajkXns
OuBHUiW6GiMRMXd8j3si828u5Ds3kQoS/+KtF2slLcAHWIGUPRh11pBtNhiV
IDHNsYfzcGUJQtFzlwDUKhSMfuiSZ4hjgWYh3/gzS8XyFd4sWfLt+2dodKbJ
V/heTs3shKmWhxXzANEvZrU9x/2rOsPQx9ndFCFZmJf3fPGKyEQy7hMMzJmF
dTbe07hmo+lgcZh/RRw4Q53cSGyk+/r8mqEJU2H8Plr3MDudcWQV3RT02HGs
SkNsu5aULp3D69uE9x8icZUvIJ1LqAbyp/NcQTUOp9L6n1yvnaKGEkYUerCl
XQMTDyxxFbibg3lIpjS4TlVAnFXjv1VmipdvlTl1qQQ+O3e6+kWCmZd42eRo
bfcYLVHdkMS6nVeOJ1574k6UtbK8i8PaDiYB9AKY1oryNJvBOX5hCzXHpqBA
WSyk8WfTlBFsZLkuwiCcCfquLEJvKKFli+sZgP4AzRq2OYOTyIUIhYtTJu/0
1ZBVKRtje2K+ZHJhISLl3lYpeylomj2hV8RyRngJwyXM+FH1nRh7nKB13zhR
yHX5HlvSR2s4mciubYR9Wt8oxrkLV6ECEcBRyG7dyA6tgoCkuqJuxOMGGcgb
RRNQAFFfsfxMa4AVLw3vckPgV2wpB0nw2R7rzuSAIkIMxR6hrE/NxzB1awD5
QktQtQsGbqmC8px0PoRYFPNVqw92w+DzxZXyTJ9krqRTdQfcwZK8ALmzRHb8
NY2JjCON68S3IdiLlfgAPPFY3aD44j2BMd9wmYu6jwDmtkxXMnlzM8iLd2HY
q1ZQgm/LQfh8APo0AUPVSBQIl4uS9Og9XUHzTk0A3q9HckAcaAFpTFm0n7rO
s5D3l+XiYjTbxYrgcRQ9AtjcHQtoF+/Bw2rdmho3wbC4IAsLqzjppkzLe/BE
/BT5sBM/anW+4FIUulmDL3SDX7w/JswdJbeKGufv5wDUj2G4AxW0bFfD9Dly
GByQFg9D/W2/LKn2LePOZfnv0WtqISfv4JlRCT8ChivAgLuhEbbhXLFuzcqr
BH/RyhLgFf2CpflSSYxmTMEbc9Cx1YoMLJNyHMp6yZW1n+jcAsTrs2oTP/9N
PhJAup2cGWgK6ZOJD9F91jnuOIp+1z4EB+ct3TiivLav2cUFoKm+6cf/RVdF
/U8uW8PJXHY1Pqv3x1SmOj5k2vTIEnqXZUKYaTNT8rBxP1NXb2KpDbALoA5W
2jm3lYo+6PVv29COZk/Tf3B2TLOjtv3JGFoXWnybzo1QS5tgz+JLpaPMSXbv
IFdY06+2I067IOEs6gBme180rpjVKXnbVPJ1NEciq/TXM7n3JAHt8qK0RR5g
WAHrU07/+myJBkXwW+XBlgbx+PWmVWGJOKjXuGbViEYJGFztnOBgvOnjinOp
FgPDcvDcqya0KJlXGFj6ZSO0xJ/+82sWtCkGsz+Ygu8yUDKH3B1QCFJ1knvG
8DlatysGQxPzqvuozWdZW/ZUB/oLT8eyXVsPA1kwjARO0AEDA7eUQoW7ryO+
nWpcc14iyfg+ehtd8+wsI7eeMI9phAGaQltOYTu8ov2fDTALJCe6wOYe1eTR
uoAe00t3P3yhYJ0HWtpKoXsCSvttE8NLs87I+bIpFWuMeYeTfPYkgI9SU7ni
RARl0oLatPigSZQIeVanJ9NrM4jlT3az2+AaXV9oYxJ8XT80oTBvBkPfQQh9
5iRKu0j+vTDxrwQrQCTCsZa3ZDH4fMvdU3F5MBaUpMsmDedf59r/DUT8n4yk
kQBN/u4CbypGHKWZ4uwKdv4X08KLigk0/nADwutOeaw7NsmblJeipuZCc0uR
7QG3TPKOxKmYg9X7VZLewgQIXYQYXP96/VJkWNdnOJ/DIr3r5lP3SYw/Tamb
Gizd02DosPx4YhL+XlaHdiGC3+EZIr5ME5RsK+B/a11SSCu2JWiP46TEFp9M
3Rs/9jhCRcp5SXMryqZswnx2rynEYL/+6/91ueeJgH6FB8uDBQe0+W66+o9X
Jow9j8+XYW74+96NaQ5kHOQnFKPDOLwWSuQZF1cf0BbOHQuQkgbuPUo8V7bc
O4NJ2gJedkKzlB4kHaR2G2SptWKQcWmMmvw61bnnCPGXTQh/wcIjPmLNq7+N
1XFTqHQmulqInTnjcXZjhY52FdfeDNX7NpKTYPc0mEQJzf4ML/olkIdNjltn
8ly5WyBLgTvLh9zgwnmx8JngUHuvk8FWRC0JDFI2VA2YImu97qVR3Y9Knisg
DEbzyjfIgrd2/i/lon4XU0EHC9YIkwaXyzT9qcq4Rk8ZqZWniD4IgmCmbWRx
iLLLJir5KBHgf+kSg+qLn0wioPIBtmZCZWPssKJLxMKbjcTxES8PVLzFxGZ4
Db/rIXwn0iGO5pDZ9ZGJu9sB0tek/yNpfu7kF12AgQFieul16/tP+jERyf/l
NV+Kam7mugkWe5PDtZO7PaLb9TGv8V+fO++XfSkcgXqAg5Unn6enhb08K5FG
kFc/GHLTLDsb0unYlvTXJpFUGgJuN8ckOx72AIVozcbBQq7xcbzbbjQDk4Wj
uTAx3PIhpu1WDFOfA6tVXllkpc33Gd8qosJJECywko/b6z0OwHKDiieCmLsr
UGx42GhpG4cjFnv434IIlDWX3x7b/ATlSqVx9lK7AOaDS9tGuRc7SOrotJM5
k4Ord1GXxPSrK86ZAhUtb0AmisRTTFMMliNSyfmQ7VnK8/mFBxx1HN2pZOvv
27FQcXIkBllYPStu/kxjfndDof/xdsVzXldbB8l2N485L7Y5vl8ubROpi5wA
BY346OpL5K3x/hrX7e/TZzPopDueFs3nvSqDJs/WZyiRks/OiJO6LE1O6PFM
gWzxHUi/sqZM4uLsHEfF6bMGiXflBoiygzi+fcvf7yeWcwXDRox8IFkydZtN
4gQfEANHQVyeFWHm2rxi9WG7OvfAFTl7VT0q4aAXzNGJT241Zvt/AhRAmSVE
uAqGJWWc3+2vGpy6rNTsHXzTF3xv5JlkBobLg2tkreFANz3yB7BCdb1k/Nqt
oNm8KTz/nFYx/aJCrjJgYf53BTIJKIVeGed2MdMDRs1JHsvYV2a/u9KlnpJc
R1wnhg6KUEcPfEdHvcxJSmtQdpAa7CdEpjvhzZ/qqf7i3qqciYH8jDnWVZjn
2Fajx0tiUoldDDg7yM48dKrhv4naQZWjRPV1kOj1zq/XE6W3rSiW7d5bIZTU
5O8EeKIRgKZKrTz0JqTnSKVc81hmZhIkkf5DVBRJAZCx4tWSmC0bEsKEkjFC
FDNDFXkX1rfmq5obdiGSjeYAwHytW7E8M1phAi5NmN1hujyw5IIXZt7Klv1y
DF+8127MUMFaigNNKYdToFK1eME7V+ZmW1RgxlhJ+aTRxm/kEJo2MOWF63+9
kQo+sY54PFGjoT/b9cFu0jpdiR8r2UVvkuNgIglQkLCgm+7a5h9rgK8Tv1Zh
TnIfB0zR89szZ+cKIWmCOHqBOFeCVjSd2wDCCJEcu6vdUzkHbVEDYiOs05u0
9NnwWNoOjVZRFkYrfmVzHlhfLERizjp/UKJ66Jkls22nv/fxjm0q9fL0WPGX
4L8p9UKZCexnSOB1o9b6LR0bgmMMTSOA7COVnN7ft6YmG0h5XVglG04kqkoQ
+zwSuPCYH/1HdrVmiOUdQS4oi1+DWFkQofrdqHBAeUdEPcXtkcYpVanBXpTw
hQcXGF380kwUJmeqBuvLrpq/zqCaUvjatecCxlSlrb4WJ9y6P4tPJQ6LDTbh
5r9Q7cyyamy0GlpfmhrnpMsxm/yA0iKhp6hNmm4m+3gTPF1vEOjljxY2Cz/E
hD5DH3QlFUdvWfVly//i4mMxpSQpJN9O4ohhQI9lyRSaTGlmyL0Qcu1kXN58
giKjbx+Ku34Nqi0vcRwpkI2W3Mcq5Al/fev3dRFS1U/FW24MzVyO8r7LXFY9
dYvo4N9R+v+gOtbLFreLilv1xgZ477paTtUdQM27SWZuxvrIxfnN4j7VwMT0
Dk4t1hu/kJsh6CF+gXtysD8SvVYdGWrO3wO2XW8r/GazX0s/nFx5eGohxz1X
VYSgsrp4dcMbOdLNI1mkzE186yMr6vrLE4wvv9qYFRgzwotaQC3A7/GbcV3i
mlfY908LtCKevBB2yc69zLB5iQgdcEOJjSyr3hM0Wite8WTeQe6yfCJtSjuv
nYuIY7ZDlfCWjrMZPuZKC04qnovJA4gpRBsSLlHza2CqQxGX2RHXAf6mCTOU
0QzXOpnfYcxWDBPwycwhykXgrmq1i74GKWzzsdMcaVetgTpcn0geMIFeCN+3
cXmTBEwKlNDab3UaxVyoE0mRdNHQ8W0nknLABIrFxB+jhlbFs5heikznpUnJ
RnjtS0RBbp16CzBvX89rItdwwCedtpZzhI8DuO4fR1ntnAB5hjbH3osNwnC1
6P5RkcZs7oZsQywIWi3JLQiI9v51m+OcA99cAnuZuBB7LlC+yXaMWJnDecCC
tj2KXtdMqJyx8Q34S8/6rEO34iHry+z/xz/+lKgZ9CP3MY4qWuMVBnfZx1xF
nZ5F6gSoj+hxEhtAEnVsXm73Sd7Hy1TEFOn3aptxwmfftbT+njTo0msbShl8
BUFJfCSJspnCjgKLJF+C0gWiT35gc0a1Ji2GjVPh83GAn5cQfrH8KtBYdmhI
FEi6J+pAWoVQSeVbvkENg4owuy9A7xWnUW086hbhz/mQ36VydP3e0lpZvPK7
qMH8Z0tQ/2xTEuPw0uj51AAhJz/yy71QqcYUYOTOjS5SQ/hgGjnATZbo2u5E
NUOlX6dtqb0Rf49erJBsVjU7H8Aj+0krxZUhT9Z39efQbjpbi8b+ueGsxUkb
ve7cgDXXarocG+rdLHsAXy6OI7GEwmEO65Y1Rjj0fSdPa6BChhJQrTKovGTp
qzQqZ51WmnHpb36HdVcrNTq+Ndc0tNa9CYp5okmwnv+ZOSD60zmf9LyHMyY6
etR61Jq0f6F6NPReu96pXUfApl03so8HtgucSBmiyPQKgjw9/WWMbbx9WqMt
hj8dm02aDP2ZW8zLcJe2Z6A/OizHmiG13zmfrJDAAgowXobKWhXWGnBqKPUY
mjf/cuqxyUfZQTUM6EhDZjkEigU29KhkCXDdqlYDADx6UkiB1mzN7MfYF1+G
cD3Vre1WWCZeNt8GDvGeZ5OGj20VTUDsPL7B5eth6vQ9xAXSVVHMxEu1maiG
KRSudASsI5+07+kkbBKDU9CJRvyHSnp9t7KuWyxhs87ipWu/njnXUXYzariN
p+xPY6fywbuVMU5WZyxHEz7CRarbtJhAX/ISKrmrCQieiIEG90nzN7QCM+e6
TYI5s57u/2Zt8GXDxagVjsg3to0pFnvfG13zYCHeTs7zIOlqyBm0/HhKHVlI
iRT3f4innsKXJrKBI+b/v+PqC1Nc6RmOs3VIEVuf6JgdsWTf/y9Tyu4jFJNE
pyIjWmFBB4yPp4d4LgVTefBsv9goMPsbITtOIa51SZ0bqTdxhxB/FSHcEv5c
GNSqtSLBLa4ai3W+l4Vc0veaCMIH6cyrwm4InFwCEYG2yRVnbXMjAC7q3Kej
RdP0gNa+MDYnxoN9I6y5aQNWrBxt23n5kBUMtCSm04hBgcyCm32oAx6ErQYv
wCVKyl8QLUGUblz3H5kPpgg+T6qd0zrAjSEAvJ5ODnTs32DAJ6uoiej27OeX
z6CxIQ47Xcj1LUcOU47eWtB6FdeWkBnM9GHo4Of6M/Y5k7zWkKCk047lfeHS
9RvQTK6eMqOQH5PagKocSSVuyXjiSSffl+LpPA5pLxKmjaF03fnbTvt6b4pN
Yv5hfiokLH0NjDNPlaDbZr4dYoKDKaqbLMPl2iiStSoiG0glMGm0YvuFYX8L
zqemEm/GoGaaY/mJwGGY7YLGgIU9O+9MGmchL+TH3GKBZA6RSxn01tjhA+KQ
tkQuh8OUF3mtasSOlBrRbptxMXfTnZjyBcsuNFRMEjRqS97pADjC01pu5lf/
/qomdlb7ogw95fGMh28ZIgORs9TjWFuSdMpIyHaL7xHVM1Zhc1fE8FQf+Sl1
jWiD0PcCWxlC7UVAkv/b9puDCIa1sOZp4WAV9r3mV1Sydj8HQJrCWTHgmjKZ
fjl3Hu7zCDPuS1hOmqCezuYapNMRl5OLHPtrRfqsLTTKPiUiV86hSXA6CSDx
JYFO/oGE4F/O4wg5qPWpkf3tU+IBoXPvuwgYQVxdSbS2au8MifsR70TwJuRS
ezRdXWXmTGPnMtlyhP8drJz+feFFMu4DLMcZHTd+HYNH4u7XKqY9Tws1mxcf
pFnwFj2ulc05bm+aF1yR/G+S0dn14lK/JAPNom1UnCepxWAGKp/X8KzP7Lmp
A5zv7jjitUaDZekaIoDt6NWaHFDhtLySIQqcxrUxdWiym+b8NQARfdMmKWVP
D1EZrz4X9/c534rchHSxrcCEDGu9e4+urTSu7EaxTn29t94dOm3k3WZD4Kkr
7R1ajBBlTl9CMFWKxYMglnix1rCVlh3vjwBrAc+ZKXp+foT3IybpUQFA4dl5
Cvbu4yzqg2GAA9xlLhdKhpsfsQw9HjEfD4lSzddXGdLW9pwPUsmTUh59IcMH
fdPH1JFxwZZVwZyNscw1KoCenb/hX62ojgZOuIJBfU1hmfTR3UWNClveu1ae
zE4L6VyvKlZz8/C0ZT+ow2+lVx5YY3VtxRu1gNub3aCCEKHS7S5bsNcIxHYI
1NEdEBgDW9v0tmM8I+LTPPA//aP4zT6uZRTtULGYBH2NJ9Ej/fknmvucgOnG
YXUNfd4KXhEmO2+Ql1MaFOPt+BAuqb/qwTXWsUzWTD7Id2cUHhomcdlLYg0v
5m9K17KSHfD/8PTxesRHh9hURzBLg5Ihyh4KEaSbyY7ca5Gmug/3/Kx5NfrG
KKYJZnebUldN3Fcje6ZfTmq6nAwh1bPH3GThrsTC/4QFgXgC6IT85SmAsQme
5Xws+rE1RY+sMe8V1f6DsGnER3Zfk9V7FTJ7+u2TojDXF9CX4kGCw4Mq5Lhs
jRuWE0A4GPH/xb21mUqDQVtMeNjFStTwSG+nJaH21xq6H7UMTMSlfagavQUt
Vy0TGhVVNEvFf4xBFjooyhcqYmUcJzWBFqiDTFpRj/S0Ao2CHfTjzYwblF4y
fYsqtZSsMvUTOUpBz+rnQFzBLfb4d/yPBe8F4TW2lMOm77V9poFFFZ26vRTl
2HAhZ0AajZLNh9AzNgm+GIZQbVPStl9qB9yXqBL2ezrurPCqfQtl3I9wxKyw
MMyERl/wDnTABStDGz5UfMImywT6YCJIM4lQl52dirHMIbv0oDW6MtfywhXi
qFYndGLR8LtvUwjSqZR74OSDv4z1+T61DUCQk+XEcL8H+4cp+zUl3cj2lW+M
lYIkYxcnP9YN0NHqSl7LvzSep8p6Yxk/4dfwZQVPbyh12RPa9VJqnSuKxEmX
uiJpyoNnuwGhH2VPOBhSZTqQDuSL+zAzi0DXUhHbVP/xZH7tlX71MIkhMfJ3
dmJKMEjkvQIkbdY7A2+lONCJekMSI2H9AZrH2LgzbaJTvrk1PxlExHBXqRdn
ShgOXzxdXrDnoJuyU17ChmQr6IBe9pbMV2iTVB6YRQgYGBrBrNJIsOU8Jg0/
nnpGU75AJy8L4W0SCG05Sy/f/VaZ09QFJ9vH6O5nsfxMsil/NbD+HsN2OC1G
7PJtopYfxcdnVyOXQeemmW0Um+0B0wuO2A6k5T/oLQrogJH/dx0lVgSmFwe5
H0+FPKSxxzXb7ABGi/pAP8vpZk9zuzGyuI9Oc+p4ggBc2tqMrC5XRQrHCVTs
IFlCmqVuzCOOsXTpA93FoW3M2ixNc/BAWZ+t8vAaITZxM1/U/xajKlEgjcdY
AM3YiDUxDzzeg0w1sogAgCQFft5r72ouEK+0CqfMLjERr7V6zUm16jssNHZr
+SkgNJFhC+yGhgqmohbAm55u3Kr21bar2u5kpneaWVH0NiI8VaGUw/DNs8Oh
alBEf22J8Ou+UbuOWeROzyu2NLe8bSQIiwQaZK0fUrf/eFj40HOvAIKZQsMW
/CQAU5MdHeSsm4l2NXw+bzA/kOIJDuuFqumKF2DEqYsfGDlOqRsJtVEdSEl2
B5mAQJ35xLQ18NR4YYHWIsi3ZkiPK+3FCjEId/liaZe7DpGY5g1+j01WV7fC
xX/Xo4yxdcrUDiFIZePjZ9C7pvwGoCrshx17lg8hLp/49oH5mgNQXPonqTqR
pbJS093XTtMh/x0WcYHaylBvY7jAJBZWmRxcDA81J9j/DJkOmk+vpr9E4lg5
TZdJSbcqXmw7hS97K/Pax2zVFqxJngYg0T8NpWoyU2kNx65sm2zRbcJM6Hqj
ve30JsxOLzuXwH39RLolWhNWN2EH55N9Qs4I2H4WeZKyBucg0lEIYETRuh23
RRC0/2BfAWk4h5qyxs5Prby2+V+j3niwu+7SBdLL7iz3Ay/hNSH63J5Z/8ai
DBym89iSuLEOlZArJKMcToggdLzqx3Ykb5OcD8Q3+6N4ALO1N6xzMcqXXuy1
YW/illT0UQMiXSPWTx1YpvSG5L7K8B6P6y3iuMCNt7rdCHuqzkjtP0Sotstn
9+v+m5FD/sZXQdC43Ivn2npnDCxSqifGu+pZof5nsiizuW/d57PB3aSrYbM+
PM0OlGGpwZ2xlIPoB+TZnM5CzYWgV76+DDR0/bA2r+LQdfaJwDnvYxVfKre1
txAroUT+KWvLPnQKnTyMDX5A7cZbHFN8uXureJPpQmC2uHEfDWlpno4nyI71
ywN2lX5RH29NdV/1mVUYzn+Hhj61LsSIfaMI+3q/ZY856cJJfa/R3UPgOWL8
tuvCVhvHZW4/qpSlR0RjlPOZeDLskDSqM+yJCjR8sz3MgO6TWDzBrKHaPkNO
al669HaKlverTkGdX78Q66Ev8rfOTA9l7kyR6vBVhUcuXIzucscDTotGB37Q
raHEg11f56iC6Iphl1xUKpCkWUaNvNXxSLtn4PN8ilWcT3ZrvDwZMR5lQRZK
I2XrzWURSnDWIeyMRwgKqI5wae3sjpQotwmX0bBIi5EEJCqZuNyZ7K1sxaCd
xBH0AYtVRSTVFXs4vFoUoHpEZsTxJ3Oq2w0zCDHJlGkziFEsfesH8+Jub2wn
gOqugZyZCJ4mWjRAyLjLXMDCzTPHPe/qOt/5HbVqCDcj2k5OfElJ3tnnX3g/
QSCdP04kgYDE5JHPXBWDaf4GY30quSbJQTeXzkV0Z9iAToZUoRDq4ad/DnJN
Sd+BZJCaV+ozNIGM5OQFeFkpqOszKPx0rBQxKt2tDKplfJ7srFGeLHoRGBnK
AhUBGPD2SxKaH+dmIQ68mfbGfET4gwIvuegQjuB2qcXUiwVhxgbY+RBhKo9x
j8jYI9kXzqcU1aG4hyS8dMgASWZ/M5Aj4lDsdyoGMuidmrRjOWge/iwJ8IQY
HMkXQ6qrW+5z11rRqvjNB2qhoCrpZdiP5415vPSEXLmy4t96oKFqjWBxAAu3
RixrLxTfXvlEYX7dx9HR0k9a7XBNsDRVGQ1e3VrE3KmlrMKEWHHq6Hc+QkeL
rHxVDU7utAklqyFwTvwGDHBQsVZXb5t8E3zdX/Yo4nln773ngc4qq9kuIJcv
J43BiuljEZjadiIfiNrQ53jiAomI7JhLntELD+0pDkjTsRzzod+qL/eFKRix
XWBPqOSFVKsnQg4byl76k/L3q82AXUj/u1VkFeYyJobGHy/9ca2JWTBPQQ3X
X2Gn0tla3KknYoNUZkX7WMo3s1HkSEQ3rJFFDM2D9fCQ48uPyhgMHKnZlm6S
I8LBZGpeoPj3aFHSNKOMp7klWahn8HXuImdahSfbzpdAXaN8p8WekTWQolR4
DlQYYx4cnjlXlCgJfD6V3xZDmwHIw2RbAb6AfBbjjtCBG4/NCXTYa1wbrdUa
w8tdN3P0bLeiuJwilh5+jnipztuXpy/AnQI0eCYX9wvwNENMzujxaINwH9FB
8NZQ9/bVTVBM8UyeZ0O3PQ+DHAghxkWAIiJhNIRuudKL54PpSFl2Jdg09l8j
GjUtfYOh3rcOK0HMhgWRxKUxHif+XIQdFPGOe2neSBj4BjcsVLYwyvPYEAuC
3iH0EWIHd8+OQVAPxcdvFOkSRJkRPAfv6EIsVE9C7sE2Tals2Y936BU+lk6t
VTWR9NJpJUXr3gJ5np6NuRI2GzVeIBP0dW86BzllvkoOvfLIyzkRWWB7SbzW
l0g2UYQVZaeyny68+w/KvMxALxFytfAIvpKzi+hF1fsRAXnlqWZGtLaDOoPA
Cw8hu9KFC5YaKkGFb+tTH+3+2CKNLWUHwtvqyxUBZmQJplHNPMEIzzlBov1b
SiOGKeBZ+jZ0KcMYjdPIDLNuAnOXeRflHNf29phoTjbDL07JLOPBSu/4C4Ul
mLvmxuLXb0hNYFJ/f/T+7NKPj1IE8+Pd5ktcB4vDk8G4nqyPOBuy5wQnxst7
a6TaJ+yMalJahFB7Nnw89GZtRvmQhcKpqHyaTn6en75lSX9UtqfBNUXz5QnD
cbXFlJenmjZrHTRLGWWgbLXILFIo1bGY8KJ4xrFssavVW313w1JZWhLOdNHs
HnGvYD+xzltTJIy77pc1E2jxRoET8SAeRETOT/dTGeoBOGAZbBRaPn2e5CM7
SfEcN+pr/vaT4rD3XB6PdCZYV3HatDztXDEgSP/DSAJVJyfBr8t3RBZnmbqq
UzUoh+As3mPWxVxHJ4pwEiVCo2UGzKb7NWpfULIvtu+w5bvZXZC8+bM6tEk3
u8azUUTC+7V+bPWAcAJbfau3UxmTowiQY8JW0lwcNw6z2MbsQB1IdZvDS33+
sLKtej+dyqETlYKSDGIU3ucla+FLLx0T4t7emUwQc9fX0/4vBO6TFKipi16S
JYHCHqD1YzhMl1b1frrGaeXGiOZZa75HpDy53efveD4doHH0Gmcfpx2D1oYk
vQjp3FZImM/dqoaUMSAf29vH4jSy0ffvaVGDS9vwQ0RehDW3F+NMXkPAigcC
jCo/d2N/mtZojgcwwIhAyjLnMPC5EGNRXWwefV5H2ejj+6zIMllBvTsLxNlf
o9vcbsUIrz29I7hTz1gJqpcGkiwbg6fGwTnx1l4rHqKV3eDadIDrruZYWpb/
kis5fFW8qsemwJKX+X1z4tKKaX5FFMo8CkFoxhn+rn1T8/W++vqIQY2LrMZW
PxNN1hiOUVSTsT2H8iNEoGEOjs7qCumrJfGYZWP/D5H64e/00jnuS0Mo01en
rVVWrXm3Q/QqmbcM3XUNJSBSHKKpY4cAw44HPxDEib9vifAFqOacfV9k1mok
MbZf6T96lBJg47ZBB9PdrbeoKhwvkC1PT9/3eB3oSEXF/tIEekQbQ0EfR1ir
5bg4WSwHX0vypMcoEvrKCmxyhVBOHJ0IkLsiYUpjLBw+Wy7LL3/o/6JtiAXb
8eD/2JhL5VkiT/iodt3LAulE7oCRjKlL4sRbA4OuJNqRj/VBtDGWWfW+nL+N
2b+np8cSd+qUQjLzG4lpkKB05+oydF+j4Qic31/h7+isVVMTwIot7c7EKjEF
i0Jzp7EKnD1RHwSiIK2lJdiNrsU0OlaML/V61QqcdGEjAxefR4HzhZX0Qb1F
Y+Ts6br1jlQQL67cvesIbtm8LvYoIuvnmQ7wR6SbEEg5PMxXxkaPjEN47NdK
UlHNFicko+hEi8qgkJcZ6xQbxF0Vb7h7Z0qLGJd2uIST997uiimLhLuMgAcF
5uo0yziklaTTpP0S9c4ouZtHqmz7yac51S9zyAz7DVrtBdgUyFQV4ZY+zjzV
IZyJdXv1nOLXIUqyX8idDt0FEkiVSiena1Ilure0AD3O3/Z1gQnaoGy4fVry
ewm5JtUFoFRnVT34dFIQ6NXi2bROWFIIWljSHDeoJtkYxZg4JexhmyFwjXv4
yGkUSJg7FvgDv+uG3N2ko/nYX6kCXPgFuvCWkZTbw7cGinoeAVz3DZS7Q9LZ
EuTq9ABOw1WsWgO2Ui+1mm6WqkxR99rJUWFgcLXVtzcWsCAav/yB43gdbPvd
D9ELeUMIUJ89ke00YaSR3Ms3cJDarW6n83ynLRUDlEb9YP6Jj+Cq6aBMLX+m
a8yfAnP5cI9peEVAH6Mnj5yss5jY+JdQgZBSJHaQKBR0uo4E125a9fx4AI8c
P7WWGkinTClojgcSqmh4dLtcZfcGiKuzcY9I23u2nRtm/rRekZW55Jsi4k6B
b/tWyd7uCRtzk7/3Si7grn+7lV9IIZPlvXfxOw1h/w7ZEBI0Svb1Pyx97XNr
Y97ZJBr4wL+1KMwuEk/4c1BEG09kTWUmP7et++VQkYB+vMHmgTqEdjY/MKKt
NBfic1riIQcFlhEBhNmepcA8ST6iysfR1oVr2DiN0GJqeAEkna4Fn11i1GnF
Xwv5y4xiwlTgougZFNDT3evv8LhjmmbugISSWGHEwjSmDPBSXfl9dHG/Ib4c
8utFcsLPtGN4kiyAHYJXhWKxLcHfM+cB1JAUBr+JVYx/LsNGMs17wnrwpj/K
217TvOH60pjXqV9WmFXtQid+Q1LI+Zzdk7L5WH99upG0a2FwgWLon9BVH5yH
BFoupPRBGuUTWBfgwl8dkHcmCGHFhN8g1bzQamTO/J+tCN4fVdLLn66qsJ+B
hByFshnNmwQE/IsySYV8XDHjmI4QDx4eEVib8r90fbqeMxw5wqJ6hfTksoFS
0nbkX3RriLWON8V8lif9DstFDH3X/+2IHmoCqjoIw4ZrUfT/OAycG2LDK/KQ
PPW16j6enRUdMphwcVfzrXVPw/ChJyl5UeiDbVqCRyjSTjLCNZkZEGGJGf2l
/gRlT6oJl1o31WB2LJsgmkGBlCIhUGclm7ExtcSK5g8ozzva6mdXtgrsQtca
9GKpIsNJ5OtXHxL1xaQIle2aYuQAU30CnU5B4D7n+AGupznC+SUvH0dDXp2Z
keoCqnfCcJL3KzjsrDN6LUceugzzbkGt9t4Ad7gBcSLWqKfCIRfaf/XkGiO2
HDUy4i0rYZP0LgWjuq8WnR1zbmYjL8rUJiYihcJXVGDGRpdE25kjnp2Kvo9c
ijn9HJqSN0Kmf0KtdthJEZSuHFBXn5+g9QfokZdt147o8v4S3vSHv5kh59eU
avHSDRDHCz8fNVVrWnx+sX6qZR93zrnZzVwc8lroRveAd2bvEX00He6kSdcG
G4VJK9cclKcUwBy6H9sIWj9HM3TlnKZK+K9h5poeynNFcSothXkWozeOr78V
/qhqctqeqQYHmadv3gCFHGzJzX8VYu9Y44RPOcI7dWZkhzwLOxwq39ob2sWa
p8vWD48cT+uxBOCvP3SoNUs0ftb0i891J23HTI/rGwZqaQanPpy9kN2zraDz
X67vSmpZVj1eQbhVnP4Of5QHnkS2fmiWrjNVuVJH9A6bNLxdICEDAsCDk94x
Ihwr8lQ3Mz9QzzA5sgD/81eUGrvd4zgAGqiWYb1Rve7RVNHBJsanm0kfCuRk
AHx/D7vwNtRyuoU47/QvIFZISfthf81g3CYDPjtPzH9Lf66UirhP0inBgz2B
l6ojRcM+GyRYiAOzFDJxMfIWvzau51zjT5XHR/zuB9wqwZ+ohcKLmym8/vvu
BJ0n9C7be6d0c9zTFmx5Qnj65haMky8/CghIAtrXECLmn66l6nV88juMSsxa
rb5ilZyuq8UKQiaEXPX02NDL8v+SilW3j7DFfwUGxFoZZJWcWJLQUQMCQ8Wx
dYTi0n/MYBII59qUqXG9cx7Alu+CAE8QHX5jDFf/L+cY4TCxRYXUBH+etjMX
AM1srQMn8zQ1K9ZhQclG8Az5SMw+8YxV81N/Ddf8K0mlHS8PgVB1cNBDRhhz
fSp8Jsjckb1KrszFmkAMtmrha6K+fumWplhr1Gbr8DaZ2Z91qcorRKcrMRA3
zJB/0WBIMjZsE4Lb+8HhiXZS4ZnmXKAf25DpQ88DkJMPToIhpl5nWXemhIoi
rzJ5x/8u9cecscHGfeOe3JPEl+zh6eWybVHZVHk1efmsfC2nt6gkXewMi9zT
VZc3Oms1QhRLeUf86kZ42KUegqheGvv9xsYgNTMEOoXq4kaNmRdS9WCJc6VT
GB870w+4Q0Iz1519z4PKoDHxDUVsTAhbPc/2MwcUfReLXeHSYpEb2hZaVxuQ
VglQW2jn2R4ICQFGC7OfxgdlUB2ZQE5iYlpSoC/HY3SCeYC48Sc5cbEd5L5R
3zpW+pz9O6HbWBIW2X9UxCxeK4jebsZzMBSDUK4i4p7tUkaZQemQFjaWkzv7
Y5qYuYORfRxJrbij5vb++kXXJbq9pozlznDbEhRjmpEnXNonyn3JmB9BHAEb
9A/h/DtSKPq3u7FKrSdzMniS4d5RdEQ2yt1wyfpuFTozJCZraeGhulXcQLIq
sBKQ0zZlDiCxaTtXmQ0UEQlmIb8UBCVW/mvdVJUYxo/AUgekDqTu8jKfg8G7
rcB/rz8iIEGkQuEJubtfGar02JTe1DZ8KI1KhxoJCTysg3PwxMjX3LNHLgv2
oM4zcXA9SvmmBr5DQAMCdeSJN3oso4vd97Uxrd3Ttjy71Y7X871n6RLIVZ8h
6GGGvCDGV0ThmIJDj+HA/WD54Vvg717XB21aTkvpfgy8JPMkFO8voWOVQ1G5
EXCUdfdeDFOtEHRLrFSOuaEuxzjywIGQiHFGRrjbGEWaXVOQ1k71N+Ahga7j
FybrdFh8ngnfEnkvFrbsPKlFGbLA53lMaM9PI0v2dinVHcmJHW97uUW0Kbu4
SEwT0JH/P92VgYc83faZ5ABvmBFi7AFYHu0l735gVYvs2mwYnzpSh+R+HeYo
JujE1vfvN2pYuosiuwYZvDGuQ2SJVFQfR/L4SYUr2ICc6gAj53bqHf1RCtlR
HRbMGnZeoCKFvintpdWT+gB5xCu38ptBk3ycAG/8+7wMsnhomh1TFSqDcn1a
lHUSfHWCzF1UG06uqSkBRHKhK5ULyb6VfW4wM6PT0nxX7MXB4ILc90wBQ4EN
169QwByd2GZu1vy23bjxUSt6pDpExpkPJhu9w9rcB254k+Cr7eAzjBjpnzuE
KL2MVEWdDH1i9TK7QYQ81zIqz0RkVz0Nkmja9qUH3Qt5Y4gf9LfcrLSu1fs8
/UADO8zPHt4Y5iAxEJxYN5wk57MZy6/dwTQfOnmBL0tOpYLK1JhrYxj4dktz
yRIeMOOW9dL9qnU+mSZGRjX/O7LGJcNnzqCXXe3VgNUI0kOMOiyRup+HN+NY
0KgrVMt8+dNAs3YNW9XXIr2oNQvWHSbMAg3li7Nd2BBeSIpIOPimT2MeyMz0
nESgv3UkKJ0/uIcRM3S1/M0MgGS2toD6iBjh7DSBFhIQIyAOw66wVuyvB2XI
4+VeUvwgHjE7likE+DG1jMH682ntmyfOhcup0FQzGPU1m8i3RJKw7ashkApm
xdswvCiuNI7zXAabKAvTbcK94QJK6aGOXjj/BBjV28NFBv4IfPeUj66Bxk0L
S43gM3p5su1zAO/3kh/g64a/mu2WqdGT5J0cxPC0+FAtkxHtuj18UTkm8fqD
H/sxykXFHc8t3WhTyZah4LFrk5wloLHUp0Lecw1zroCFd9nxkY7aMn4QSXlN
lleL6rNvYv6KPprrWuWQ5sqROYHbfFTASlRJ85khpsVAIqC04FzyhC6NLoM7
1Jo5mXwaGpRjZx1Brpc+MLzJPMC/0Cry8E7uql5YJZUji2zioaIQ+3E70v+4
cmOXHi80qdperrHBbUCNEJzux5fAy+imdMwKPO+IHd4h35VWVevBzJ7RVro8
ePb7BzZs869PXCL2tFyaES1k/PyB0ReeaRrFRsUBegWgDS42RIBja8t0fiVA
R2J0Sfk+VJaRDZrMixr47BRBZSdcJmABN/RaCUUlTDxRqABFp9eKBzZjIi65
cddtDmCdKCYCaYgWGQLIDO3RrDjQ+L4O9oPm9gsxYs2Wo4eC+/cQIqT7RK4f
xH+jyRAOOILial0eMMCc+E7wGae5KuCxZJWYWwuz/OOf8TbjC/iC+5vTrAe3
t1AJIzWkcVUAblRMAkar8WBvXCoaEo0DFC8BGqU/JIa8vZ41pTEvvE2ZVnTF
9qXC1fh/24EMEEHa5U2GnSQg8TWZUun6eWUUh0R70F0kRoRfO2Gs61GX1Vo3
3gBRFTuKUuO9RgH5NJaVdIFdepf5sx7+Rn593AAEF/b2YEBJ0rgLeTXNVLwV
maqcvZXRDSlRgMhcyGz73hpFrvENA3qqZxlMtiMUVUnx2JhR/9g4iHUIPMav
Bh/zof6Q3qTzJw12QYbRi457WeLf9IzuYgb+jO2gM9vUZiXyGLM68+01d5WN
pEuV81rj1+iT6FMm596E2BxOLaNSzINoBE8F2bpIHfhml2K6J8gRyEQj/9Sn
Mbgwj57SRZem1xWewKeEOlz0e4fUd/2EC/sRUopbBmjA4Er8i/Bmo9H+NtSk
03TpQRNQMUJCupftybjh9U644DBA3QafVCWsmOiRAdgp+XiyCNbbaCqFpD6d
UiMX74Ums+BmKaNxwmOpz9ZlQgRWGqLvLFuuZuSkGZTQyiyueuwhGO5ExKjN
poKWChDhBi4EvS3aQr5jDuuJV62XIGOVMRYRy9krjq+bortV/DyXDRKOcnLp
+3/Aak54fTTaDu4R+S7N24efx8LihBKNI/iNPwza+FfW2f7rdP5SSDyzuOxX
njP0E3CkOOp+7E5gu1ltlzr8NtpCtf/DpeTNRHQb8eJ2f3ylDuqeLDSO8D4I
CrPe3UIeT+KZeBOgKtm9E1SxVOxdo+d7GYU0NSeTu9Vu2NWlcLkw51U0OVuu
6UukFNcpeY7i9VooiYwbGVWQCY+s15Aks84oCNcfF9inZk6de3he5nT+qibF
nuYjk4cTn5soFfxty/tdVIxFd/0ZBIZl9fDooW30PfELB+6GUEuvA6xQZzSN
bDqQb/YPlCALqz2O9X11fBGlZYZB6hHqYojJIj8nE5pSW8ey1fK1545XLzel
A6TXkCat4K9b2xq2EN4TVdPzRzLaUDt8WuqWGSwbE77q62XByCyvZEfzbFKy
LP9eofFlrSEgH1C+mJCQFD4PHTkCEE5dCcWnJB5/ohN6O7LZOYERPDcD1avh
j2acyRzfrqRURxrAS+kiw0O8+QLNQ5yebMt6EmQev+uc+nK/xOfaijMq743D
r9uskCmyu8itIlFWjMyvBA5ZZ1aSFKpdVzybjzP68JOyemqECdcs9Y9kzYQn
+qnf2QpOrC5S8EwbIJdnsjzZWjb0jV+xjxXVlLa+5eyEhAclPLHxIjeC9S9Y
dxznH+G8/YO5gap3rVn5Db4opAdgt8ztBSG2DZI8MADlkJu+21gcwSUwXT1b
lLJZ9PGrrYlcuGI494zeNLa/wvEPxf0KbxQtY+KHJmvMR6w+gf0QTke7VAaT
nfWUJEWLp5pmms8lZc7ZheoBQ2+4VC1jVc3CevBz6tuY7IzOWKGj+bbmErjx
OFJsuBg9r+j4T4VXaBsNplx5FSZOvF8JS0aIrflgRTVChu03oHzg211yLbNs
5WOGrdZDHnv4I775Ch+cbyt9/iUvrDNUQ5/JoNBk47Qo5SzbNKWJ0jw65pUq
X31FtEQt+nOyzNX72JjPPm04WHcoHBUvfHjJFU+1JPw68fW0YrdBeK6y2q+K
Vu2cBzXY5u/e4CyxDzAU1uHCRXCdNDC5EtuPjByn1MIO0cGMJWrvzSBFWl3O
rvxITpTucwd4/WpputA532m1PrZUmrZ2rBUkdMWnHdA+o/pnJxXNq2wUoX5F
MVv9sPjHXsDlhUnMWpBwrs/cSGx/VWWKFypYRTkF2Wkatd/RnBS13aZcyppt
GPe0Wkdcyok8aCXWvXBuuj8BgaCQlh4NfkgVk8FRGHwBaWNVMBTX2O/eK/r+
MU58YCPOZahLkmwf/aknvz2VDgdL6HYdmpY0mUqHe1rKAJT/WeYchu9BcYIu
a8H4RPaU3Rz74daSMU235nlFF98Tzf++kRpGL4GxLWJHgWJJLQfHBtLLMMjx
3B8Qh6gX/LeJa6q4m62Yc6BfyTcS3McmJqp3FRwtjkUAvf0luufNu7rL56gm
5aE2ZwE33qUYxMi7Hlks7tLQ6xZ6eYU57dqGuUvOjZPkwufqDXm0L/JnIYvH
DKoaxIXtLcvqCRDCBlf10HmUggCyOnypEofd/MCayu4vooE1TQR2M3FX64mB
ye0UuqK0A8AB7s97jzH2/2ieUERXoKvlF23MpqBbQJLq2kLvd7arXkbtJmwb
STncuCzhEFcxOocktAPTGhSOTtGySYoLrZCBU1B7oIL8TKVWTzvFXHiAOuWx
h4Zl5/eTGR6QGPh4hrgVk0CormPNbNhglxO4nqpJGttyNgoG6sXbX5223Z3G
yDAd7mbDlKzShlZiaxZbchh9Fi26bA1zz+MjmDmGT/b8s7zyGYcpiE4UvUkV
gsaYbR8Ii4Q1yoox5PsECugaDT/S0bmj+6TshHHGB0s9yUXUCs3BoQVzsUV6
t01dN4+S3OSE0BI93PKuaWod9NRiIXy6REQA/E3wpXoQKN/UwaTuAubJejty
RfkFGeuc3uPx1t+hvPDP4B1j6qqwEssiTxwKvgtTj58v1gGKChChSJ98ZDbI
7U09A2157Ta9E+YlGHjh1UlNSUwMTufwbbzv6f3PM3JA84PnYsPa8M+1FWMN
JJGDVBfdRx8DJ4fnLF6hpospUdWW58ByJvKVGF6R+lE52ZbK4+24uj6/+sxF
J5D/LykQ8ShQZG7UPcPEs4UxnN+Z7Gvx1oYbYFmEfKIpgcJGOAGOt+gEWFlV
KlFxy+w/WDhDFmzpFlJvwut47zXussG22NHNnt8dvYN8Xi4riv5bI4rbShOo
z88eroPDEizh9aeefesf2Ri4XjsvZe2JwQFcDNCd7J2IQP/fH1+lpkHDSjLO
GfoR4BEXJnIgM6pqlKmZFTzcwOBuv0heDpJoA7wApLfiy1YDo76KKe2AXWym
6+qgW/j1UPr6VBed8GnyZNYzBuwHjlDBPZ0q05GNUQlyNwNixA9s2yxRLH7q
UtlPqrnkujf/lrPGQ6358uces3meh3sW9N9pBKy9XsRb34x6/tKr8U4ugVEu
24A8+gffHzZ5NzWWfUE2VPl97OldbKL4Cy5WahxCWJZ99exwD8EHD8Y5mNkE
FexGSkb1P2JDsYhjIEk9t9vCxL6zBaSboDgl7hL67uxaZiDx0Y2Uk8tWZMUc
a778Fvmh3AF7f1nl2v9Qmk8V+q5R8DGvOY3y9qCiewSOmK0ObAYixbYef7fm
4auPBoH8sXbc0/zsfAwDQoJLOKlZp5eDDIPlAdPtc7dBBoT4HbC9xFKjx3TQ
7vJWHgLVIJLbK8eeCkWlm1HBYX6r4ypSn1hqxKH/32wQVmrmI3BqRGmokbUJ
mgmzX/pUWz5h08vKQAAUQrsD2sYekiII0WOHvbjbKBJBWcrbcHv0g1lxcwPi
N2lIhz16g0pH+WVgnohzpWpo7HrL+Nr6GmG35EVv5+ln1141ho5S9UTXeLVa
kWZ+Tc3fgh+IT2/cL3SVdaNVCCyezDeYcW1egdj04IyDFdYf4ZzEP/ingxf9
hWwxC/w1tpgBiDMQ37W2xcg/1jMt7XvydgL9ojZoA5ZHHKD6dc2vc+fepOz3
zCgkG2SY+D0ZM19VqFh2GCQ/mCYwYFUaqZHwhfR02HNUhUqDcHmGTMGVqtvo
qgs08WesPGlXH3RODU49J8iOiu/V2B+Ag33XXLKpItiFqS/XgpRJDksGy37m
P+hDOzwqDSNMdafUbxEoF1V2615TDRlGyaSwhrf67/Sw5dLzfdZj9Cr37A6+
5VtYZSz3Tr608be4ZEuo07NOQdwYho1baA+Rwcjr+4FfRXUAk8PEq7HiYF0R
3EuydoebA0zqalXfkLnTanql40p7duLUscKbMRK4D9L9ru3q6a1a2mGaV+SV
ey/fVOJS/sZTRyQnVEF64T0+RWm5jBKVVlY9SPNmhPGafY7Lf8vd8YrAzR2c
6iceFgpSbPREy86RnA6djl8C+RBbNNOTpLT51bhwpsITjx7YUY4bq7g6slcV
eUXGxtW7Ujb7jO9fX0aO22+4X+AvYCrRSTll9rdTkXyJDvY1VaZxyLOUoZ7L
og307+vyjXZxSi1n4k3oTtmfs0NSDyJqNsPdeLBkjP9AmuU7RcPCAFynq2KE
FZFWYXf2hSHxCsIzoVHzwu59JXMD66XLk2U8ZDLXd/dJd6zuoQq0RwEmJDb9
XxdsEcJr2Ux8WtBdbxiI9KyuNqjqII/8tF28YZY++32qUhP4q29v1xhv3Ejz
oB2tOVsvbmKd4Qn4yWazTiKakUxgAg5AUMU4BrR7MQ2Wo3I6H1Nfr6taTaMT
TU8dEiKupe+oIU4eFEPMJAIbjfZ1MmMzqfYGzg3ydonrFL0ssUtvgrkRII0l
hHZ+QSpfPY8hoKBbOVIH8BvMPs/viEKyKLeXKH0VjlRcHpf8Sa0p7P4ZDqMi
cQjWoPu5OYtLJ0cGOYRrKQAva44Dm01J1vVYiRFh+muMMT0sOrOllmuO4w2N
F32YJ2S+sa3tNyX3eIfukvCgGx1YBTH3H1w0ugLtcqqJMG6nUo6bHIeIbVcd
1RI2TB2ZqxLIYKd9MPl6bbwnTJjtWIngXXdHeRBI7AQnCuWoFeb9Y88MHJ4R
wHYvA8ATFYZxYkwrflLadQNPqPi6i61/i8omoln/IiuX3AurVpSazTKIgAse
c0fnHsNBV8gBCCsAEmtj0iPoH85Be8CrALyJ6cxLEQr2NTbDexaQBcUsjebw
pptTmO2bGgKpk57bmBZ2mSrjzlC+iTx6Tm5BtVdqwyZsFF8yZnSx9N5lJCW3
zMAvBmBxqT923l934G0UUMPZlh2rc+KxIkY0A37aGg/U7gUSrg26u+14B/k9
75vPwHsTOly7gT6591lshZxnCK5ERVlwajqLn9yOdlkVuYm6T0ap/2thGybJ
9/L24Vgt4PkYoaafVCJeMCfFAH/QPn7Q/r634Nu7sRQ6A1snW1wiZPJ+lHJR
P4MreXheGnoGPr1LcH/hTvkGwvqT2AtHwg3l417yutIoem3I2cO4xeW94n+h
pMzYiL53KovTzxE/+hR44dmsiWK6MEd+7aMc+QolmpmpngwpuF+7kKt8Rr4s
t/V4JzUO2zMJjPQjguZCOwDvcTizyJO4IYZ+6G0ni2c4TdRR9Z536jcBp+X+
y4/pQJDo2XOjcWk+Q6Qb7j4aYKHhxHJSH33XyV3fLD+nn2GF6IuAIvEKtXkF
pQnOIJqwtgFEwIyoMdKgsduQB7wksTRM5yMK0SublLg6oaObg3VeeqKpVryP
MccnJ66wzJ3+QgMfX2d9RhW0UAJLB7sKHd3/I+Pr1M8mrJ+wjLT0JyVAWDVS
kGUH1uEoDUEwZq40L1VVcyD8YWwKqtY4wL/YyewPxhNigTOw7DlNGFq3CaSw
SXPyUFFTxzzay6kt91OgXAzZJfOlhPF5GhMlE9TIAuLxm6SGLW/mKoZO9I6w
mhNKrEeRwdYGBqJhpDgODSv9FKac5z1R5jNfbmNiApvNBH2a+Rcoe10naH1h
J6kJtUcQOO8RirmlDUeSzf4egWBfdUDtBQKWtDB96YYfnbS4iK9/JIvwwt5U
9GxeUsWvVQpz5uLshVKm8YjsV56shKdYnb4B5xfki15NRwe4AQTeNEYqGek7
RYgXNmyjczX4OrTW6VBSfcuFqw/DTMUbMdCY5oDI7JmHoyaYjvt1+Nne4ys+
w5A/th2CfO23eTrcvLL9ooHuel+83XtQZp/hlfB0oYpL4U+gBGcIpkwSJ98c
uarhmBCBCp4u/F7PJTo7XtxNqmbgMJ6K4NiuihwJRCelzSbC1eNBEL8esbtj
2DgbuUXau/eFLI7/8icmglR2tXtvYPMs5m8wLNWdTayO5ijEX1jZK5fbfyPl
reBNRdnrlv4aIHs1v1D4zfZfjh/LoprWK16RjHzx2Ba6Wzr/kWgcOIzRDEai
tvayZGd72liDMhMeovR081Oihfr/ujGLiR3ZSVM6NF0SLTjRdRRP1MWyDAVy
O6mJfjsBjKH44sbwwZoeWonwbPJIiDgMSz0dU+nmHGRKRqDbk6KpigWkEsjO
dmgisMrZQcx5Zr56JkxfdwqnNFJ0hygmTI+CcDaTzgjXUkFuQJPqlRUQbsj+
6Qm56FqwRfcwigawEev28/HIySBgQ/XywdDS3KO5RaY14hhMHVuOWXjEWldG
oo9L2NsJX8R9SNQV8/KVJ3PUxpVmTdWlTDf+bNzM/NpqrYcXq8QGO4JrnDO0
m/hPBxzport72uG4zNdVIawOz/Iuzc8VaERLpBskiHAasHno+xZ0Du7y31B8
sV8PeuC8SNwVGswZ0S0CVwGdjGTZPdnrIuzFmeaDfMXwius4zMvDypg08kyY
gyHloREfkYgoKrU+5BIgb/bj+trXqsGFl3HlncL5RmOZ8KlqfbpLJyV5TW88
NUVR0MdPA+8NZlNHcRTQRwx9Hi40WifbK4o4gr5mZjLWyqQglyE0a5JYtXvY
OrkdHXxgsBAMlBt38x7dmFMQJvUQpjs1R5cEn+cfMXQ4iCUbhJaVH3pEz26y
YkPRF0uazqUq6cCV9P+CyCzRBcpaxfOoU/bf3upxmz6NEREVHRTzVRUSg8t+
QeIDnGbX8aPlFW46u4KWe+5rJ2uSQu8cjJKaiaOjrE+MwduFkVT/kyUdhWba
HdhQ6bR2swwyz0gUdOxbvRnbQJtcIajga3IfSyqZrJY8YbsXVcTaODMOl7xz
RNRArojL6SXPZVaOBVxqMkR/52+e9Ye76n1EXjSklWs4dpUtWS6SAUOGPwyQ
cZIw+UymuKBxXmqmnikJ/KJiYeZXPjWfrANhB3QFVSJFHj+unn7+cuCKK46X
uYujK/4bNpXAptu1m5nSZK1h2X+GfwWXG2uMvc6ZfWRMZUK4KaK3+p/qliGV
omTZl+xn4l3jMQ0Jwpp2FyoiG3uk7lnwiVo1MizOW3xFZiuXrBjMwDIM/2Rf
5LBh7U5arN2nWy/gg9MyUSykaCbQGkPuy0uLgfrrc+arQYNP/K2Rn8GzHel3
jho308N79brDZEJE0TxsOcoGSkDzBx4dtg/2Lt/tKW73Ny9zZot1LqOKjZac
QtziKmt39DfFej9kxRnTCZ/mdjRQ1SkUJWyD99VbTJi8qy3WYdRKfhp5QUkr
xWqU9/i/fz60VrZcHwL5xieR820H/+jsfhSbVEW342Dx3lzFRPGZfyfrhDO4
H/s85GaeyP3nLa5LFhCRCwFg1Oi4Cy/JAHk+ATqNABQr6cCyVvCJg2piYzW/
Mus5ysiM9DzklSZSiD66bzYz4DImP8LyzIAjJ5LpxU3u1p0WTE/CeTC76lk3
IMNZCLSxk1HWe4u/V6oiLiz8vc36f+wJTeRBJum862LyPwcWgxfhYx8pLzIE
ueijm8vqbZA2l5GbgokD7+5zyZu7BDndBjUcM9IPf4dUeiqKfBk6ULw67Qyd
maqXPo8dpsMmzbxtC/kFJenvp4IiXoM6ZBYtFJtQby/+6nEqGbahwFPS4D9U
oWB2G53w4alcc1Vp43kmw9P087N4NpJXpUQrNUHo8qxR5z4SxRK/0E0Ot8K3
iXzYKs3/RIhtEpQqK/Glk3ULDxh/ZHQ4hp+cn6eAKj5/HH/FRuqhBNY5NUGD
yL4wTA+UQzFu0SkjWkR6Kib08nvbfJOfBR1iIumvdsXAz3WaRQ1gxlcz72lm
iRxjBxMzbCwPF2ywcjwzuLFL87P0GqyaJqfxQpVg8AhlZ3wFe9/sDqVqahnJ
4wl/jHYDZwHoBvM4xFlaj6womKRmHo8kUjsIPdKaM4ekSyCWDQqkFkzO5nYR
rWvXhIdnzEh6z2JCPx/GcBq8KFSBqhZxDSAsFRTKb++Fj0CERexqACsy6ET6
hfKMnHiFq2m53/yswH1AeaFN3+aJuo0mEtgMRQ+NVS1YVwQ2Ee2YaLlyh0ZF
yVwUcW5uMsxB/B9rUpHriLat8/5IVCoqqz4yWE17UWNV+aTiHyGe0fkkO5YS
2xXOZU7DZOpOe+6moQ4DMHGkzMPPj12uRSWiRXCmU5kyUI50ufzIgwL3qJvJ
TkK1C8nHAFr8bbhBEKcr8oYTbdlByHA+zPlEkwfg1Rkc5ldJlhy1jQzpFsnR
z6ywYuz7PLSrJtGRqFOzWTdyANPTuH2JMhByaq351aHohvUoZX2TPddBxD5x
E4CO1mfib0RkvQBstRLhWJhPavRvkTKHzEQGfyfEVU16gGafOWW8r+uoyvBl
Of9vFJVo4dEY7qLHw9EFHRDti11mADkPVrqcL0VBSElr7U7onxHuWkjTq0Kl
XbpDQ85spmqU0mdhvHtANvznhKJxh4MHGQKVO0Z4WyO+nkH3h51iE9EdbGt7
IBW2GU8QlgFmxPY5VN+f6WlYSjgCO200/wt0A+GL+STsmgRa1JO7bUXxgvyn
2EIc31aMgVpkzzJHA4G2s80cnfp1uOzaiD86kTIUIv3NFGKDcT1rM9Sd0vcW
+zlko+79n/dahnYyGEbKWSuEesMBL+0oTzx14jcd/Hw2/v7T6WsNQVvEhG2v
upCaZrPCrToSQLgDha+QYSe7FlAq79idQ/McrpyZzGmHUEt7D6mfj3tQaywu
40oJFb2FFHe02Rat3lG07KvePlmGoED5hue4208n94A2vPycxr9k9mjXJPvr
RswU4f8xaljKLL6Bxkr+TOGL1hkuEpkOoUVSB7FOZQn8NTyVZa7s7T/8mX3k
aQ1BGr62vsCrjHs5KQEHckGjYxdSx1fijyjdoxLWRA63nRm9rM/We4zUknQz
FHnFMBRxRl3rLB3eqCVQkor/JrjGYTDEty3Voe8UtNKUEQ9HyyM27ya1h0VK
k1LE0wj47WfgZVlDEsbsME6lFHBv+pblFNuBxaiOGRIzndeEbJiijiTLoKjj
1RPt0wiN/oZiZJ+hzGiRbGGdfykPCWrKKYDi0f2uLHTzOKy7thSRtzkXRGXd
I7vnnetI/wfg+6nUA4MKa2zhAF7X+k9kVUNa2I2+mVET94mUVooE9g0yezKz
36ggG5qyGhio4DwtilMpCgl9hciSGbWISi8TuXsUwsDQbYlUeIv0QGKD6gpD
9+93KIobdSlUGK00dkfPt0SFx4CJG6fEFS3KdFFuj8kd1lhTFXtWT2nWH+oL
u67OZP3ZH91K35RrmJnoPwnFudFqA7NXM4WXBMVr5PS5XFebQpAE0P2h11HS
O89eIw/ElJvqargcWSCCI/1hPzUiGVWphG88yormz8RbPpfHpKC9vWPO++oK
dkAbD/56djjeu+od+pxgXyVNUN5EkFe2X/vUsM5tCTA9YqgbFlF6F3C/R7uA
hBER4Pc/ruOu2cak4feRHbi/uPy00EM/bkt5jaSDS9c11WbfDkFj1x6cjkyd
bsQng+6619xGiGOunuoBymNo45GRDGO5VYilg0TSpXX0C+VLz4a3vCUTSWvh
nwlGbeqsPKGbjeo4QuTpky1afrFBFyk7MXeDo3WRmv/iD1gqLNJcUD0PY+ft
hmemB7IGGK0Vpio7P8FXERC+EFAURG6y8G+1AEOFHXiHACtfeQkz12+9Dgfa
ESPDEDGC+LR3RA5dZF0kUC9bJ+HYL8t2R9lUgkQzsdWbDa2VZqTc4ogaSjf3
kcdOWg6L89mezR+9dAES5VeE9eR3uSiHm8l2cmrUQR65tI/o2g5Hz0SOIxkU
+qUSQaAzJJApYXevD4kkYLtOk5JZBnkyJ0eBcCziCBIUbB64vtbcSjLwD5fO
GCLXGluLCR9NZHYU9hCrWUb47HX95F1siXzUUjy3cDUPdUiPmY+V0mm25OsK
nFrAeRbx1dsDG/uxyq8JN7LXjrrM7ZFN85Gfs/3QVakyeerYUtL+BrhhL+Ua
b8l0xUlJdnlZdLqV5rYuCMgjSWVDSD/wod90O8/DLlAG4vltX+chqRpVEUzH
kat8mikETA61uhCFZDSzoyIbkXfwsGwH2pcD16TB/m201bubZf59X3TWbImv
+t6o9ez+gBZR9jzeeuc9ntfBBjKMr4fYeHEAtmOzl7iKJYRXnnQa6HFhkEWo
UCM7sHpD9bJDK87xCzP0B5+KIarrX1zL+Tj3ukvfeha4p6B2HJHck5ewoCke
ygj/HYcegF4Hy+U9NS0hj3EfolKiHCy5E0AJMFHfbF6/cenGi/UUyCmRUoMG
pZniiGrfYxI9sD8igIgmMcDSWUyKIntwvIZvcUaSm0tSHnpfVltCh4HTIHTY
AqpQgxXHluwXPvZ2Avgy2954JIEpzCqmQPYVoEpG2avuHNUpJ7IA3Nmn/6uK
MGUSKrVRX0otVSazFAo77pC7bqw+vsOboSSgfyDar9yTJbhU/43l5o+ee+kp
yqQqg7F6msijF78yB22kBresH0pescW+2K8QMk5xxTs65oVufD99hg64fjdo
1P+d3w0blLEiHRpQc0RpQBIvGp2UPvPvem+fF7U+7MjfV3FFa6V6lOEhU3S3
ivn3VzoMjnBIhzTYiTJ6GhPbXdQMyTz0ZWuZchbf9TgIBqjrPOo42lH5lUCS
JBZvsQx5oq0saw5eChUlubJRTvw4IHRN/dgz2FariynPiFUW8p1PoEG61TTr
uX/kQlFK99la7RIlGvxEUbdNNDGczEJ6uOJpS88pDRYd6O7e1tBUHA6FZ3UQ
6CJTTpBHIxzPhbhdfBhvLtAITIxOMf9zQONWYNT46lp9myBYfPIBd4dSIFSe
cckKgR8yk4c12ayLBEqspFghgkOEKMDxbo1leWISFoN4v9BehAE0dszwXz+2
EtrIwJGAznyPrXV6DDpcudYWo6eKDjwfX0kLgpEltLUVYjn37Yw0wFAat+oD
xLd9qs2pwbYD29YBv5DZ6UHoGJYMK9A27B1+DDgm8Mly+8W0A802crmGFg5h
5O7Czz5J4opnBJFAiJjrqo1IANQvueOgOoAr2TVsDvZxJfVgbKgHtN4xNR2j
Igh4ZEoQ273yCvMypN6uCFkuLpwFwnPW0GcyfPSd03bBmgio41sMeU4l4Q9f
mzegU+wff5iq5Zsoez3l6MA61i/dGCmDGoDYz14NECh2L5Cx1Wi+kj4adEqb
VzwSHx36J4Qxh+js683Ud5e7JhkNVi0d9DSst2YGnjtGn+O0Lq34X/nx1Pbx
hV3MVPBXC3PEvD5hSg3cGyHnV9wYHy58Zu8ad5gQMxz8t1cZ706ZrxEaakXD
FzmR/R8en/creanlQo1ZXbYJ9dOppQ6wPEUfaW6zskd25JbV3DFDbEEnBnZV
DW2wQkj/CHFpW/YbveR1aBNrkw3IeS+CwidVvUtdUKDEA2dWutt7Advm0bI2
Y3Pty+V+om9OVykyg+N45a2t0GGPqcljU5h6W06CVVReh+SWzOEuixWoXcOW
pvHzfHoYj0xiGMIY13QIVSYpLxs6Ux86tgjgOlmnzGBTxynrqUnkMkEQpnZD
/23xKQaw375Ld0jeXpodlRPdgDRkfRiefAM8UxovmtwTVSo5dXp3YTUxXeWm
ZQGECDLoCbtpHAgqVKe73HX0GNsq8eBBQdrye+n0D7oz/7tWDrVWjjgw/6yR
fuZrVwh22z9U3bqxXl/1slzKddI638qWKK4FfOzWMTPqwp9PvjQ/Qc9z6d41
/XkNJUxRLjc4aOzY/TzZoXVE5Iso0CopSE5GJwuGFJ+6brPKiCcm5RFOSSdq
uEmKpS3K5jGEcVPi7xm4ds2WQ+mDllMcgCtjLxzUHP7E8AZrq3A+maD/MEbY
kZUQ8Dxc/Ffc9dg2/gSKiUnOWtrS81YQvuANI5xmyCdUGT7CWTicDyJs0aMm
66oiBic3iO2UgklQpcSJazbc9392EfY9uPBHD8uiv3vI0NLTnrYKPUjfrB5n
OXSbrgZFMsTH63yLJkDRXjrwrGf9YY64CK9STyrbxxLo4yCRw96jS09jHUOW
P3ax9PvNQ6gRWRqHr/stctj0d86hmU4Wg1hS102ANG08v11OfuYWm4Rn8FOK
YUUrsiYS6Sn8IYtG6JB7Mmi+EajNRq9EYUeJrGr5cWW5D8JXqA97v8Ar7YZe
wgkSRZ3VGeGsaL7u6e/Vjfatbd8UBLlWPJy4ElnO3Ck4svrBpbEdklJ6zndN
QxOPFnJ0w0srhIkOlb8e7l6HYDamvOCNbul9+YIESM6Bs7rBpCSvTShuKQpt
d+rVgw03x8h1xCD8hPA1ACvD27WUaS+0Cx0J8Mg1/x28hZoYKklmgW/jMeDz
XCUNMkjjK5boLJ/cuZ16xaCqKUnkPeHYOlRUOgeAxmsaQI37HxvjbODSHwRd
9Spnz4UrQX1BqZg1YScB79FCFklhpsvmOBf5XKoNxHiInUtzwe1i8CbJ58GG
JgrJMJCzvb0C71JkHj3lsoKp5Dm3sn7cBoK7QkNBMF7ErrSmcuh+O2Er/ttk
tOhsiOfp+h6vHkZuYqYDuAEOpL7YH+RNy3C1DyAsqMVrhnxyKqZajG2aRoRh
P3Dfr2VCWOqK4DywE1wEOUbq6QI38NElC9AEo0k/U2OSJQ1NyyCgI5ObFdm5
8Hm6hSLwdvPdOJs8HZ2UTHMX1jYQOXHYbgYzB5zD5NGl3NDydUeznDYBTkLj
5swfS0IHjs0n+L3Czeu3c50nQz9VUNypBopkvzCHJJb1g9MGrHAC6d43a/tc
g/Eh3KohomF3bEMMvQyNp6DLcCFFG94rpLiU65pXziDsN3ST1g7aaVxFBPP6
I7DMis36va1HjxYlit075zWiy90IF2/xqvQFhh5D15ZQsxLT/pv5H2ue6Bgy
2CFFXex589qN4NzBsEHFfDxsnZm7DyUGBaQKVU3YL/KGTv9sjekYNwtcyYhp
vS/lS7dlTlfchoJLCB5t969/FCdWrHMlbs2YvJ44OpZhKMVfyP08jkyNaFcY
PIZ5H4zo9d79Wxta2iP70+BXFstcDOHmdcGz1/2ZX/KBefvv6oocwhZ5BYJM
TRIBvgyZIpnlcfIa0dvpCHUf0Pk9lMDlyA/t+RAzNsOOkQ2NOKLJCc/ZEw/z
30cNeFGtZia6LHY8xL7+s9whBEzgWbTv9T2dyE0FdQ2QGIxF2fiTlYkQjmtp
GgiyioQx3DIjrEkANIihZ/pJnJ7jchreAYgJ1tpHDIjPNa3oe18o45AJiJSD
dkz72uPRSI0qvFw/lJH8w+paWSM8Y7xUfJVwcGvLUVBhfQAXLUtbOEXVZfIP
nPnrvpiydKDll9kHHXYXbtrO/UiBtNY8h4Bd6sbZEfzVv/NwVcTWCKEt9jks
dC6pwk4Q9V8xAkooC0PO9QJxw/83cDzQoL+euU1Zvm0x8bOquSllR6wlM6tI
28d1WCjR9LUcmQmylfhk7eyjepdw/4dwOdK/T5dxSTsriY0xeb8OSD4Bm1iC
ghxKlZ9oPgDebHWXlegbtW4Nu/svYxlKbSJcULBSRMlxzDlS/sIKwMaIhLQE
vHvDB+j7aPdU0ru0V/GmtIs+L6f1aX2M88oDxIpDB6uwmxBUZgn+zW7oPOpn
LdWc54Iqbjeclm+4nDj1q+n0FINpDCGcuGm12OTPnWWeali82hVzMGHR1Ydh
YYLa8+HccM/0xByRKmlb7tq3lVj7NbraRYbFNN1EMD66EbkEnuARCyDMmoB+
0TH5HCXVouNZTXaJ/txPD/f+1MHAsWQFGFYb7aeuA06lgdnH7fCyFfWk+yv8
9XBBA6uRcwIQI5Gn3hPFIy2bkuNSSKeb5oCaYDpvCKrN+765DnKPzEfyuFBd
A5yMifftPEnIMwM//SDkvQgXiC0ew/xkLAidatQMIFDj/GDNmMdo9gDRkNAs
sVvZZRDgiWF+2L7UVWigTDs3ntut3CFluiaSYrdv3atxKQKCj4fOS47d8I0w
JgsrIiTRM5JgPY+1l1Ve9PlEgv/fEMM1+cjBylnb0P3k9Z3ea7MgE/CucgyS
eYTDxfPuzdP9sa04ZH1aLX0jhxBAD8B8GFwRY5jMNWXeFeTiQ7K7uVYu3gkw
TgCLSUcliE4jrxMg3vsfuX8kfcUT7Pp0+gXkOl8in6SafWHMRArOHqnAVDkY
SH/vIoohe/KE0Lvwdz27jmypY2E54qbX8W2eEzgViVySeydBag8b9IPETl0p
tQFpKm6aTEHXbLOBir7gp32MuiZn9b2ocspsp9IGfvxmtXwm6xinxdzP2wcI
oWquXW/Hm41+cNcq2qmmsqBgOm7J+h8qd5AsmZp8qlLQjd5W6A3jHlD9aGRh
KRwusUqPhG0fdH2wn6hyCA6ad/YTHHaZ+oLss2HDSLLwFGI7kfI4Cq9SxpaE
cRwnbmj+nhoVyDaa3gWjS6Zdo0YO+9op6y9aC44x5mtiPQ3P++wwz8OZHtsu
/+8kssASZTE3+gc16pUUWGG1zda6UG8vLHk8Pgl/GqqCxABLu2HhjW9IPLyI
eqVpbeQ8nMnGzenGzM/Ei52OwMEe27Db/0yRWJrsZV178P0QT9VJSz5zO4IE
3O7fC+2iM/SIMNcHZJmvcF7BdCPbf/Go0iM5Uj1tkgZMFP0wWQIuFPVLmWQf
yBbj42SSER/9UWOvU07dSiEbcYIOJkMdmCCpmpI9TzxYUz3ohfN2xH5smt1g
lxqBckyf2mIyeTr6mBscy/kTUv0glwVC65Eoxx71YESGV+dKRk3AOINSSu1U
PT8dKw5SX28aVJIapwQA2mz1ih0KokcpPpY6Xu6iFWKyzTgAcOu9t0yPNvFR
SOgQw9YJXekc/xHNiM3boN4ysF4DZjLPvDrE/7oPI1PDDCMIlIQuaMDzpQL/
00pZHnlp+dMVfVc8CLSTUYYUfX388zzcrEDgSHfQssR97WHBmHRvm5begxfF
v+bGttuVhIvCFURVTnv2HqL4qblnpESUgG7ocbC+Ckr5FonpTzLlP/sjCfU6
QeBB4FVaKMxXyFYom02eK027ZINnURZeiGSomwckyuqsOBRE386PGJTsR51O
qrC/sLSPKvB1KpuP62LE2lPTLoeXyPKDjlqSLfCA3otK72+huP6kZdMjk0XV
NKkTP87KqVhaNTNPtuVrtr5OmTvzFhaPbjMo8/T2oTY2ZHHUYcuAMUfVPzFd
odf3wc+2vyZUgOKE6Cw7dymf1r/6V3Q0ks/ABziSclIBQquqSJZt/e94POH9
n89RxXuFidcLVvyE9MjoB3R7kcK1f671q/DoT84NBqjResyJCX8YZzSBdD0a
M6HACVGkCnhOLjuD0Ikyzk4uyoeOGU6hri2U82KTsfsCidlRETzyAZ/mSOpm
jgj51jgjKnTrbMEsro/MDYfp/0R6QOb6LJLHAd3piRy/Qce+E2xsDUu96l0t
u0qLoMeBWxGqShakJg42D0FDbzM/1jVCLvbEQ7e/3feAGzOvGeFpWiYlx5w1
qTQtLUGpYrEHSv2r5ESK8iRNz8l+EXlts9q/SzdG3Ohus7SHnARon2ldNxuN
gJIwLW1Le5J7vz2L222leMww3J3AerQukZI3HvJVOSGlHmff8Nw/fw8c9FnP
xPrGHwCwueDL/Gz2Nnvuwe7jt+L1/Ibe/7R/UEfWUugb8xWM8Xg7sndO0F+P
+u4n9rTX5zIHkDSq3q84Fa4Qgu0eB+jgEAuNmdaDN4StlU/Tyj+NwI9U+H4J
bQK2HUmWzTCdto/MgF0hvrl0ly84azWKVGCNNXV2ov2lNOCOxUK670VkL9DK
6wDhHG9PiVD6sP/7Qvm8a40aAAPdVDgOCCj2AwaOVPu5wFwOJ/FlqYwdoZFi
GsP13c5jmY3sxrFIXjBgyQ8BK+kqRuQF2dE3rIoJJ8D5pj4GSbKpeLEwxXGQ
oRkPbm6cH7KiP1x9eWeFiKE20zV6POSPWkdS6Tu3XPiVV5RuPSDdJzdjil/k
hkzkDl+/FDOlRSqktOGk26NgbxqhXBZnViq7GmpuQVLQV47K2Bs4I7xyyR2U
GkMyRKqrfuiyiqEf4xUVoDmhy8ym/VN/TT39pE1tO1VL6FA2sZHLLNGvvLSR
T7YL+xRFBobLJHFTYr6MFyziTcZpk9NIvOqNvop5+owWqNHcFJcoyDVhOIgW
BFx94dxFjYMQL51WAaHlYHzzurkjYhq82haZLofkuZogm3X3j7GSEnUJrLsX
tNxvb27G6WWquScc7sqgPCEsGCLQvWzaZpBMbxZVuVwDX1YcpSWl+jugHIWP
Tdc1AdQLmyRVslwV+eqhZazVryGNLkXg4blHakEBEcYzm3ILF3jCGZwOqDPu
hsmpHMZS6sC2yU081GOkLumV7QBaxXkxyvkH/o3rzmxvRQwVQxrEuc67uIIx
9VdYeEmNOIegQpJvqtaEZAFJKgdkkuCqckCYbDsrHITHsfICqZhdPGiykFUV
SMdw2UTLmHqCiPd7N4zUldhTlz0NAyJj43aBFA7b6iZ6u8V1SiwdZ3FUA/VS
hT3HycaJb9GMmv6A2zzdKeU7V+R9T9Nu+T0LLCGgVYC9rnzvzW/iLZIOE1KP
jw2xQ/U+y9GgZs+qWb2eh3dqg+XkAqWK4xtSMr6qTwexOT0FofLCORWp/ZnL
5fJSTvMu/VYeVht7BNAmdl7qFEGy/gcGDgNC082wbL4EOiLI1Nxany+TX7d+
0CguJ75JU9s6NbnXCXp2l7tCFzlZlkWorr8lb3kkQ1JQFj8Qm85AwEC9GYKG
JhusrPOc9A2VMLI1dTVZNAlRspDrpvh+IL2qbaEiTUdT/W7wsuRx3c1G0lB3
lDyfRspusYuTCKEw4yfDkTDe7Kv7qRS0vv8bz6D6lS4DsbfZfDtnu19+IDbu
FLcdvdmtmVO2/TPHXjkvaF5Byhmh/Kan1qw3Grb9NVPCuKPbfzNYcimwRtP8
Wno4zxAAFRlwfvXrY27aQ9elzj370JiNL4zKIh1yH+xVa6eXmGSiqZeWsX1m
eFBq/COCgHg9Eco1WpAV+8keeC98w+B6RGGtMewszsdV4loSEWcasHIF8pIb
9EHZjnWfKgfzROkQ9hx9RfTWrlZpVQokc3yE8BwoM3NtFXkxFr0mytEViDI8
/5g12dHskTIEU10zgAu3j40xeYZchaiSmLgUF85YbtAeVNwV/QFwAP9B6Ftn
HJWOB1wgHZrRQQ5t3eybnkJl+Me/vQREIJEoGxhIsBL4bUUpQEdyW8GSYUBZ
cRdky5/mi95Xl28TzWR/WKgz5NT5cj5rJ129ssF3ALwPyEI5SJfnujpWzpNW
5KlB/W0WhUJpCMmqoMvlRGuAtjRAU6QJMIwHf5E9NlGjdOLwkqtbyUq9qkPt
GQ39cnTjYArny6W1zfTZAIw70ViO/gt17JMurCBaI210tuwrvmz9t+6TuIOI
qeQ74fVKucDvjjQ5y2K46vhoI9QCgMsOPwK22NK1bi7au0ZygrWSa9w1Mf7Y
M6TeZfkNssKhY+dFia91Li3/GxTe95OTQsWWVUwNmw1v3iJPvoBw3ERS2yXW
0qcpOcxOoaDCT36mbNJZqT3dw518Cc/58406DYqtLsFL2sss6I69cNYeJc6m
gTM61cP2isEanOKdQa/fmbjeiBDOdlGimzNUYFRIrjC413flTGx9gsF4BW/v
+ZGGutmiABwI0gXR1KDxcIVagLlGliD/PZiWsoYS/F37IGqx6ZCigUeRhVqs
ZKCio8ZpuzZuKBpWK3mKWYF5hvDTpu58mJ/fabZSrbFdNYoWYK1XzlG+GHI2
GHeiJAxGznFWbt0BMwZ9pyHPxoeoTNc0Yn2zU/Q/u2CMhwCRWNUAu/siBQLL
s6w9dEFCqo2DpUoLlpfdJpF+IOKUzUz/17Oe54CwWIwGQ85NlBkDkF38gmT9
BNi9WbxR+YIDIOQZAYL7tTWLchkyLHFRi3h2df7tlIh1b7y9au6hSP68lpJa
IPyaQOMr0g5ToLxKBhLh6yefql99/hOolRvcsblyidNlCaYRIi+HPm0bpuXJ
oApjwMeDlISBbVFQ9cJLK2HX2hgQsifYE8CmZVmB4Ygu/w2Mn65C1zUN7+hd
oq4mPrG6/zcfxiOFBugj5aHp2xkvzXpiqsN7AFjoDDTqr/y4GkSJCLlvhjeu
NYPZDZ/EBxjAWZ0VDBPb8fb9aj+4HBtFA3mgPKnqCKKmb+qxC48EN4W6P9H3
EkBCHyIFV2KluowAkre4wcTbkK9jBH9yoKIJKKfgOYMXMJxcMLRi7zyKq6TU
41BbKTOvVOZje1J+h2eV3dDHKL5fF4VWvbPt+hPcSp2w2J3m3sVxTl7IHg9t
lAXb/vZQmO5njZZHXZEqbD4aW19WuwzHyRUOkqw6b6c5TExQT2Y/VngM/nik
QAkGsHGrYtfBNb6hRO51j1dedB/3phJBvV5EBQHuDx+OgTwFgTNtAyddrxPN
ss4lW/FqIPfD2hvLRgZXWMEZX8s49FWrNJkOTYVM008dssT3FsDsDvz2GoNK
cwt9nkSYmparSADnEij40G72eIhel1UVW9cbp+CIabjzE6J8HYhbhpZYU8kh
cjPTtFCrciAb2UsY8rAf6/vdulUXZNC4qm/suXGwKEUClBe30u1iPwTYqAN9
lnT6OAHOajErArh0FpWLgGgeNrgQXMk88dgzxX4Taz2zXP7DegJ/pvLoR7Qs
/wQa9xJLW7LGacF9n4we53B9fhHyznSQtJeg2ML9QAJ617mKIZVJi7OTXDtj
BHlwu/72H9Ie4pG1b6tLHK+AB+VFYaO92fv4DPjwP5kszFSN8Bx7BFnmkfks
OUUtsNZ8hlb2Foeo7curvGTPlGtwhIcYYqgH0CqjP2my+svuyus4M9+RNU2R
N4Bhs71j1QmYG+dkZHkSzmgam075NvumIHMlOlztUXaJGQTcfnuDfNiZJvvw
NKmJIpruHG4iHM3Xe5u4qK4Rqwp3erTnEfRRqmMJEYPvAepSz5cyDLqaedbI
sSCDi5+xaS6tks7jYwm/Sh2tjxPPQCCimBMZLW5ktNIICYp2HnuYgP7zVCAF
jrw/r5wynIuCBb0Y81s4BbwfEJwAsZkAnHM6VRdTL1I4SExs42wmor5irxJg
DiOTOuVno9tVS3thVgWZYB8eiRzp4AiVFEcxd6pXbVTVLnoKau+YDwNNP5uN
VF6++/g85qmjhoEckOYmVvYpPhJKz+2Pb+C4pI8dkTMA0shZGxxXP69oG0jw
SRnGn3ZoIYjSKDVQvbPUfJMMVNafjtiGeTz+NnYMW8XhktT4gMlc8BM0YUCd
G/89gxnAJCZchUMQpq/ef0Ha5pU777OwlMnSobOZJWczg6iWmaQ/Gkd6zCsG
RqKDLUgfwbzNgYQ8RHiMiaYnEHQYv+lAdQ1Tv+9DuOF1xipptVPspU7VmRya
kSi8TvVC8+sFc+qIKh21NIedDWhDEFSKK8PgUCbTRNwR4cvOr/nqNS3trkOp
wt1oBNptM6mtIPUIFaD/JAbp0MJ9bzFaNdSJpygT5ZhpWLo3eozTcw5tHllt
eJMBYj2CiKxlw9Zo6sCWT4NtAhMd0KnHMyLJUzPfqKHFH0C+Lw5WozWOit9n
/sVjuUE1EomRI7ettmJty4+VAzvfXB7OY8VqjHMpb674ilkBAWbaqNwUJE7S
PpsAfgH2rNYiK6+Xzf96zpFVcWfxR08R6/V2AZ7bit9lY443ipGxEE92wNdw
yQS5NigJC5fCawzRMPGNQvVNdex7jS7Zp0Oem88arMksvV0oYbJ6lDNcmMps
RFt86ehxuvJpzXSZCs8Imqeg8+HqBItjWU3vVZy4xl7ZLxhPATgicw0iKbFy
8zVkerzF1TqKVkDMvCWZG9b3xKBSn10glJ9yOVYBmtBDEy2k0EPTD184s2LR
L/DOpUsfhjlwUlM8YI1PDGK+KGIDHo2tK/Lp8ulZa8MQYOguweQsBPeA3FyH
20Jk4lp725DB2BN5kIrv0LvLMl7dyiEUuj3wZosvdUY48xQzmO0vhGfmxdIu
tNs3B/aJmi7RWfjpKCfcNZHMXjwTt/dB5SKwCM5FDD2foqyn60wsSdOuXRxp
r1vMaZeNTXb6pCXUe811eTBzKs+UAW4+sA9jDLL9klTXTNTNE/kvVlxjLtBc
/Ewdygavlb0FOgaXVdaU72p0mTx3HKLFi0jSrgWxekCJs+qBkul//Kp5Sy4o
n65atUIU+Bkw7bK1R3BPHvbi96kIVV1ozX1Jl8ys0MEzQbBPMWdj4BjdQ1VC
aN/Hsia+S0eFVG3Brcz76ddZSHYYvET8xO6J/krs7MHL5wBeVWPkz6skH2vA
ABppdaD4JxEaD6vKFB9uKAsaa/9f0pzA+09Udf91wlSyUiFuFojHXSRiFKgT
jQOzKLa+CHPzta/C3if2h1Y8akOZoJVWIT6ChFEHVpN1kX4pmcuYlbZtm1TP
1Sv1k2Zjp/jRiYsU9y2BNYB00Do5wLH79orZkMWIQuljNUAO4uxsLh6DrotP
C0nHjYEvPt7mr9lDLk2rRKZUvMS1pXuWS6MbU4ReNuJ5ETshf0+LaF8updeA
PLwHT/yFleM4lF6mB6Dj/mXGMwOxM7WQ3pQEif53LKZSpIOYT0UTO2ry/YCy
BYr8J1GR1l5Za7ksYQmOsJ5GOLqEmhBCLW5Flkn+HlFCZkTM7wEQMht+7FWA
JI14M55jnZGwSefzC5VV3eqzA2MdNpqWaL5nzV033tc2NWg+D7UK9FvBeaaz
dwDPH4YJlZLWLWVJQA3GB2qMayOJUQiLqhMunxISCSmjCOAtphPv1kGZBax4
fzcOwGq75bp2SO+FzrqaxrZU84WKDnrQ8d/dqU/Q02CM+LFnf3hhdMvUknOd
OvQKppgKQZi/ympO6J2/oNHhkCAvaBon/Y816f9iihCDi6Epr49IhfdjHI9Q
c9Ec1/lV7tGG2dxYpdRc9gPCaAdXzWLmkH9uAfje0zXYvxfW+e1FAN8kcJD6
4e4uxt+4WYk4+atn00QpAZFbyF3klXjzcBGrCJBEJ9NYt/zmEzZW26Gw9ar9
7i8rVLLuRyqetmeDEZCIYGBioQH6zkvONPnJHSYDnmMDa9jD7IpBGi8jAYYw
dqEUbQpcWHGX57zViKwLSp98qDQ+z0aUNZqhndvImeQ2Ek13dBYzG/utc+Hr
Ueow0rmaxpPvCD56wPPqD83ye83wEUBZ//BEnsUm7TR7tTKS3qfjaAYHrd2+
sQmI9NdAzMy8ghw9PwsCI/47XXj1l1sjLPUOdUvxgh2+2Kpwabqj9qpDpedd
cy0SeETgk6WoM/qJqDQUpZv9s5lY0dahKLjw6+6mBLDa3VI3IBFp+GIHLGWd
bUKOzzBdTdkx67p/qTUfZSVhE4bteC/tH/cZMadmj6rk3+qTGDjXTsGa5Ry/
ckbbKUrJoJELrGB0uKQzwlw3hzn5g08TZNNHwG52geR4TMJu8RZd7ywiexYH
SYDR+t/eubi1cn5MjrdW8VcUCVjzhh43uEi/pEDcKilqB+fuElicsskmb8V7
qwtdltzVOMa92gknx62HkASj+R8gn1P7rfO9tJp6ur3R0pnO00sBm3wplX2Q
doJFNXzzvQirkYHj6XkhL00kfh/tLf7Yx/ClkCLXb1Eh6u66GafbDTzHLoIg
Gljd4qir8tnfEGOhEbdJuS2DcpvxJlsdnMQ4OO3+Por5fRlrVBgz2GzTOBvm
w5zBiRdK9suC52gfNRGsq2Su1jMM0VvFUq4wbVvdHelbwvN4lMyAtYOpZ732
8QJ/0MpVQGL2nvFv2bQGAx8E6H7J/1Pq5HJQVeveCoYJlZKJxcNz9AcerK2R
NBtnxp5FH3naiXKZlMX4T7xcjD6IEk5RzEayxHVHD3OksveXWhuwygCnTT2X
KsuvzcdS7DizQOBsUmr3BiVT1G0ITR18cP7nfvoXqiQQp2f9nrPTrw9qYf+3
S2wdbI+SO+KvWjwMyvwJJj9FXvwhAFqNZh5FxrEnjuFrVMJnFQmTG9aPCSo/
yddtp02COZbBVM9NUfRwlQ8PtrcpwGOVhCv3io7Uv5D2s0kZUsAWtR5XAQ5o
6T2gPE+rdEHrXTgohJAA7zPK9x19ioWS9ZRhDqJbGoc4RJ9TJdXh+Zl3b9GL
PIrkom8O2DiaHEuFcpg3P7EuAXbstoRya+3DlyxEePHgn37g0yqgk9oV17TP
cBsOADXNwsummTzFAORqB3iiYUfrnBkazq9FQPefTQHE6lB0v4id5sOZFfRh
RgtRRYVLQ7WTAGFA8mDwynLepkVNKQUBdlFhs0FjVFunk90TRkV7Ae+Dkspe
hHta/gmszC1WC9+Cw64u9GMvmXMH0WdXAAs77bh5/gWdg145Oh2fULN/zPa5
vyCbKjXajpzk/N0mD3oFvuZaFHdm/BxiyX6WD+7QN4Pqcf9UUKCUvvnhwvDC
DICVdcoAU/3bTfm6+dZN5QDJXZInbYZP8jwd8A2nvhuEykvG+HStCtrrxbc+
IdF69uySPcwFc62nRmW553X6nDK1lm52+/3FJxd865XBwsNf2oE0fymE+Iyo
qV9xQYPZFyFDslBsn+7JQpUuhLPH7IexGvgV9hhX7okeyqdOmBUaQmseZNTd
bc5Nj8R9ffMVfouMuBQDcBs1FOsl+6mcxb4vB5MiVe5lDregohC6KMnx5Xp1
MltTkUeO1WROXxj2I+AmqMLIR+py1ewGiQHf1OqpfHFsu7G/jLACb7mPOMGb
eIrWLv3+BiJmdmT2k12Lqti8j+Jfaje2y+NIBSfGFvcz2AxPe2iVHpWjPzdU
PnVuU06zVNlscz5d07jgpXMA/E4inGN6ZwQlJmYdiH8OL6x+ZrQjecEbbTfX
+lamEXWB1wuj+FJYvS8xcP2iT7HQL3Bh8Qz6XKfLkayeY3/IoRQH164Sv7YJ
noxl7oFsjlvJGJnlLaXoD308hhRMzWd5PlVDFzOBxHF3BiMyd8Gl8upbbSyY
3mGW5yHpWTqUGwLTyjMSjt+aOzd53/mYL6i5IiV86ortH0XLugdp5uy8TjUm
6mHg94GdPftPgIJD4vWLJyj88AIoxViYnwfZ2jIVAYgqA/J6o9TpROtBClmR
YxN++PC+LLMpSeidkBtT7GFxWrDr7nrKkz2RtwLhZAerBABXoVRj9YhoPZma
nJI2qzodqlwShhFvfw3zuaszO4EZ4Am/nXH3W76L55MnwvxQa77YnjyZ5aaV
kDN4EnI5jQuTorQHa7M3NOrd45F6a13U4kf2mm+P0409h05eeROXborZz1C2
PoXYAiJA/fvE2fT3P1Wy7jsKL09vRAnUyu2BU2KEUvqiCfg4Bw6YOVJAoim+
hz36UM1STZHU1JIHqVjMEOBFaS/h42tR/rX27wf23FiQL7gDY6cIzvdga7xx
PbcOCrL5rI3oRqY4MDlpv7xK+jCk83b0hhKb4JMrsTR5Az3ldQjXTZ02xIad
NjQ5b2RsCvqJQFjWpQXJ67PYoStd0P2HJVKT0DOpzxB5VFsgyAdLmCxtlpfE
OLFl4lkTbVIPr/Y+sGZ7lNTXOoRP0Fj9WGi3vwIMkd5h2apGKJbJ7MeBc/ah
NCTO2OHjIwd27BjufybbywihAE3jhz1q1KIa99z4AksNI56PF3ACOKZk5Jee
/gZmbOftxPn1IobLBrFgwpAvGe/7L4DHh9MbuWiBD783X3sHKXrt2aDEE/Zq
NRmDqvTP2eEhuA0USKbcCZAom1TitC3bYkZFKtwx9AiuFeXXM3/bpv3E3zLm
xbLoDH3KSxE3TikF2rVYueZaiVag6EhiLjPppD+5RcsMY5JRZ1i5GAhyObEV
7YMDjrSNPP+gJdvvmIpeNuVFVfK3TbSa+VH6bzZojuGdDiqhUj5qo6VjPswO
MdcxTUnUYI/Xo0j+J4EsfGpe17nokOdgOOTd1B8W1r3JE9VrsKfdO2cAmEHB
i9u5cGraQZzg5oRadK9F7zcO1KpEJfQbk6MjJ8B92RMZejyKw8KWGb/Da9sJ
5ITJi6hcPPnOknvrQVFg8DuKJHj5ivowd0Xn5tHx6uWUW5jeTs3h4NyioCAf
9Tr9c+VSvh8TyaG7fkXbx/8npku3q0oo0fPkTWYYdIyusN9+3g9PlPTDHwTd
0raY7SmdKEbDQ2/EEiJGfySdnzg8cHau3y4cIzkEpusRIS+4wpLQbaAGQz0E
k7PjdPN0z9YwUEnNVc4Qij0af+NZjVNKSgrVxN3mAWm9nzcm0bPS3hTjnT7S
uazWXlGpPXVXgNhhEDyAsOsI5P2qBQnp1ZUCfl5uyYYD0T7/3ZSq4ib/fUYH
/U+pHVCAGJZQL9CLr5IZ3Ai6/MuFtsYudWxCiJ4oPxsIjy3Ez/D+xFrTAfNY
6QSSUrtyufo9lZA9RcHWShAfTR+QL+UMhJJl3tWZXqaEqC1cpMqCjjrSPxTj
t+THH2idolWag3Q1Ncb9c2nkIR2Ebb1Z8cSnfZNCZMnx9WbrjoIJD28pJneE
USdgEb2pAW/v6lxdasVAfXH3ihDhw0NPypn3ZKlCP/eldw7QLeXCNllpHyRb
qHIG3VJdt+JW43Utl7SL+9jTK8Cd7yCFawn2RjkDplCbuRwzl/pi6kq20SG1
ULxTPkgwOuMJxgQTaiL668HOd0S0CokOQ1a/ShBYxWh/WcAcIWFJu7VK8Xf1
dz/mXWaVphwRYBouUOdEIbeJ8utotoXHwCrd/DaWLfwnr1KuyFhUAc1pS9+q
VBjjIrf2RF3CkZ1r4KIgYDpjQ+MOo2XPQx7CoYC4Mb+nJ0v1ll/vLyZ3mSGT
R+/EoRSrieZCRcoBEAtNF6w+QhEj6tzPaGVj+pSy5zCJHlCmANq/vhokjkg8
F/S6mfjTMqYdwPfi4hLbdGAUq2SKjeyM8BP743OH4W6QXz7a/uT/ZF0MdfM3
OIgf6TYGwH2BiHanVAjA1QojC4chV2cMD8Jdiw0WGSywoulIV2sP5JWMUR89
qA2emmOajJMvh5/hESkw4CC6gjncJRIWOLPDd8SuXiviMCtApK5/+yIpaSbE
6izVHy8UyAMjUg3Jw6Mx/iLXctUntklCvejX8/3aBn5JlXI0NCyXiDfcTu0k
x40LrJHx52qRVWevdSM83c7DxZvjCoD/nZJRMBJfl4ix8LW3WLZI8wUIM+iA
7rJQq6R0DJbm83pCl1MyOkoIre+xtQMKlAVPBPQnMZyzZc66dBk+z1+1I8+x
CsMEi/N6LgqEdYvFxwiAhSqSfBV6MD0MB7RS9ecfiwrnL07AK0WbKbXS2cKF
7byeNNogHcbzEwnZRNO6CvF+8kUfNLhxPO1LbW+QSKlwbwLNkvzCmXalT/g5
ng9NEngpdd1MFD6ym1zHWGQBw4sQHBt1FhnUTmV1HkKjgCIvpGY/TfDwGguS
Y/pNsiMc3k/hmVHXqbk2ZmPHDNOD5G9HJylvNuaNy3z3wuAGqxn5MW+OOz5j
bGstm3cjgINFWTa08KrMqDdkgyGw+vWSzdU1sTkBScgRRLFm/AlRcToqgRcR
Sa2oEBmOGWNpekEvo5PJ/jivv0PZR2Zb1Bf0ug1do9DQ90mGoB1FW9JY68jC
YUE5TdZuQohZYLuqlssvv7oM7d4KNPFxN5UgHkNOSHHH0zi4aSVAX18SYDJF
P6UmS+T7quoNW3lmpeyVIbjqxQHKiJpwBhgi2kO/UnVBEHVVayxhbRN6G2X4
yhST47OlBcopnAJog7XPmrKiavilXreNU564R7OIa6ZLqbCGtHFHtrPiMnP/
j8yBoy0VMurs9xOZTRNv4y0INLC3QmVCcagaorqL+xpdpTpO3wNQf2YBGGCe
EAnJGT14TsA8SvtgnnwyKnq9TJ4uVMEkJ24lBlt1ms+ukRD6mHxz4USv9tUV
TFLD7v8Y32WyNiCw3K9NED9TGAYOdAEw94sE5QBHDVUqGYP7RIK1tw9QDL+x
VrOSG3OQvenvj5redjLBs7ItXhVOt/ALful8LvvZpW83Jzs0AA/1cczn1p5v
izxrXbPLl+WNCVZqzgQJ0uT45P6NdFYyGWOMsaFyvJxf6jQFQvPc3sVKaGG1
LZpP3gh7SySiqQzraDNV7gpPTdnbZihAFkWMlZLr0ed0eQhUBO55hthDsbHU
+Jes0d8N92L5IYUm1O0JPik5KLdCfXNXVTEM4mEbUNDJkatbzZ/YNgRNnH+0
X2DM01rfDWIvLw8pZ0HVJCt/v4haIYHNmYG3PB8bLXl0TSnDpQTnlDj/VJ4w
YBPrddt3gwiC1G6JFJMk5qeyim9EsbGBQiSZIP9n0MSFpt3WjTlMSXu0nlSs
gdpa0qmc8VmoDlEiEHun62luF459O7soCD4fHNnOfhgcTn4tvj413CId2A+G
KJdAL7u/lts/33ypEoRWPnL5vroVWOvYr6WGiGZsiw5g3Y+opN8SQBEOLVVA
LhUSp+pmR7r8irVNuSUhPhWV/H5Y8yvdH3z9qhyUEfYwYx+/0kabAUm78aqq
ujiLkdR4PF4j+H7Sqz60KWofa3RtQpLGyoufqdgQ0BzTLnWlE8/jWB/AzIbO
TL2O9STFcLoFlTeDPtnjccPIZK/xd5VCuxO2rgUn7aH4v5Pps9m31iHy7bQc
Eq7Tb1fa82AWD3AOGRpGqdB0Yismm79pXnhKQmbdSLAzB3z4p8WhY/LuMfRv
g9moL/1toTohxjitGGx9TQfQdsNez+Vwva9WOiFcTbArLz5MuuXp8n89NVLa
uxQbFLtZILr4uMLVgMLW2cCRB4C6UBPnzsW6emhKyGcbGbyX7PVjse8pORHb
gMi2nt89oLCytiOccN0nifjbV9kJS8+YNBzJGM8sGhjjkJDn8W/SAT+b5Xzj
uGRYkVFV6X5s36UGXqhCerENBwq1G2sOtnaOSa7NydjaPJBVXj5rbR5G7wYg
QJ87hEX9Mv4viS5arnTTjeF3905pjbs9Wd9ybc7EnyzdshbJkAVtyxefcwmg
n6jfyyvYWzmCeRJlpRRmxX+NJjCKOrljvdJnQnChbyGSw3S3MwYvgOsYnOsh
XXjZA0piNGt7rX2aHnUp5MEkCkxRXNcWS9zx6pG0s535aemMmyhKDmgrmiT4
OPxvpQYy94WAfNQwKeYfuaY+Mdb0jps5x85g1ZBICJ7cdQVmIrvyKRlUaF2P
AMPcRTBEcxg86VbepQxu1yOyOjVrXvZXt66JoOLCv6sFXiSpoE6zWO8uVUZ0
7ZXNtx4DcOONt/D3TvxABBWeKvhgPINWuf7kuaq4E42otiFV7cy7PwqM7Jzo
dkqokIhm7PzqH1VtPd1RJidbAHxxnR9NLRZOR+wdmWSm95vAKwDx1MfZ30Pt
2LQ2qoP4HlrT8X2Xdldq8WJOEASxbXFm1uDSSTpqaBixL5cMZlS4kb+MZih7
sgq59uGft/oxLWbxw4DkDTevE/2Gv5YOahURM9/8SArwyUQ3TmXXamSbXd27
s8P48oRTSRmepPiRjCztuWs4sRDqLuP+DaqbJtDejQW9cYwaU1gMO58zm+xK
OjTDWXjw6lJbeWIqfxJ6+qC3M0qWYeTgQNZfcAI4Eru0nqclb5wqzhe7cqhI
iPpaM3Wy8kK2q6vKhUKfwa7DrMnwtuxTtHOT4uHInXmWc13++/2a9uXT/+kG
ZVKXZxQBfFcjt+RP7TnZRrFTpkUTKxbwgh/vSLyDE31ervN28QXRuemZPfTx
y5eGqT/4psDFIr9Ux3cfJW1TpjUgJBCP4ZGfEIjDnOoO68zdoz/pGw/Hh2la
MBsxIt8SDH9Xw1pzFRjD3pmfb46bJkVlqxXoOi+TrLcEzipFZY9+hRCU8/kD
DawKGHER4NmuuN6luBWlFA2PXd05ln9C9Yu3L5w7alJX2TyTWrv5eijEGSlV
hSHe5NH0odpqJyC7Q9S/qkcKwUpmmVu9wElFqB4kae0MiNB5m0sDv5wRPhLI
IR3BEX63MvTaLuEVPYargmVTEsA8CSTQQxgZk+y6LdRKu32Qh/+lpyixw79b
fRbLi5shresK4rUFJBwK4wUDScPBB7efkPxVHTf0nkFDIWy6ishgrjwahgyk
+Z7VOaRlHbiijb4CZOTf6xtPiB6M/9dQeMZr63kpcqFVndkd7FTsbbOphQBO
ziN+UawPwoM1Wxw4Ym/OlbCmDmC0Obz1az57tOG2svSeAHqVlUBKcZLOYZM/
UDNJb+RVdXusPAFm5gN+JvE62zn87Dn4X5i6G6YyKHAKbVtoTHP49AixMp05
117LokdijMJeiugkTuLB68IeDZlSh3qRWcnL68viJkSXQSzwENOpvYHIZ7/B
e5BCW5RVXI/uXN3vOdFuYUlsEtlnm8fAXAds9lLySr0x0IR7F0pJVDEb3yEp
I+1SITqbPCbSEccTYte6a9vTtpmTYJq9dE6EQHCrgr9pdSWuAXZo69gPXnax
ucC1ymUyDDqliCUjWF/b85GA69uMRp3DqX148foQsdmuWehcgDcHF5r3t3BK
vGb0H831R5CXoPD5ns6OyahCSFkrHh5bseCbvgjV9eaiuxYFM8BE3l8ioBjp
OBEOz8r/DMopA5CZPA4mB0qVYaRwgtwwakGcJ2Be4sCbBji9FPHQYV4s+TPV
w8E52YOhrCHNMoH7ypx7+B8mTmrfXthO7ckUe/hFWCASApr+Ee4TMbsPYWss
pq37eQCeIzI0YyNCbevdsM9NdvdtXX0+GqjgtzUUbLbDNiKpwtnDdqSXLr0F
D8Wmm7kDcPs4EffQTgTq3i5O9cJJVthBesh6saITQ1okfndXuigkIpJgdyfk
Dfam0IhzXSXykzgSqKcQcB3xtLjXnpkoVAjsnpY6vTJy0nlPycwJ/9meD5A9
194mY51p45zq7y7JJboLfvIkNCi0fnTqdtQJuVEeZE6b+boM5kkrTGQaWliy
BIEW+rll6wUMdQeLABlrQLvbMsuHjq+i7n0mzGMrxmjC/pNoO48lznigd4nk
EQnJY6WkfD6JaIossjFIeKLkhcVJfaURHjfYZTu+fcfm1RcM51ABcbBp6qgJ
WpmDUTYlhthydRwzpXX93qFMG4QPmJklsmh+FNwXoCzIAuBG8KUZ9bgA7Tap
RzcYPD6wHtJiQfId08Ccx778F2VcwZhKwSwsOfo1ztmlSa+grwc2ehfTbgW8
SdiMzWL9hBeEQ8hamMpyl3obDrqwEXTT06+admeZ5pnFHgZriE+S9fEvA+Zg
1tH27zeMSzR3v0wfmsYTrkLInKI6IijpyFDqeWYM+9xhlRWoqQKXDwjkxcGV
AE1npY/Ocba4I1XGUBSdiG17CdvqqXitCb8XX5OZ5xg/8o/9IyY+Z3fAVmCH
IS9H79ghZOBKt6nS29T1mY0nlxiJ4egA5+sRWJgvov9SDtrT0w7NImCAfmTo
IKN73RYpWltk9tqStyb8o4UER4yO9e9bG+17hVEKs8P4r8pFNzB3Cb+4uOfy
NIhUbdKo9e3sNIZEKb/QyvG3rIcILoazST3zTYlCScGwmXfJRuZUu2O6Au2l
z9R4QWjzb0nVKDhN9odnQj9eO0RVGcChjd6layVdjpw7g9W0c7g0LQe0ZaK+
VhIuJ6+zeGfMrmWKIV5yPxfgcma7FbCjQuyGmCvehh2v+8iLR8ObP4lG94VP
SSxbPkN4a8AS3xFkGBVACHlskILdpYP6+DRoRfqbWXwR++fIuO+s2LeGv9D2
0zQprqhe0/dp2BmUH4o2/e4KHZ+hJFvAMuLufiANsPfbcbevWrva6JrwD5kp
z1sbmQrH1njlwpqEha/VrbPKclceLfA1fge+6M1pvhU5Jb2aeHJY5zXLbhXC
7jUYKVh+5OV+IWUHvtbK20ZXsmcv+6QEbBFCvQ4CXc0l1yQQNmafyKZiIdlf
rW4wbiKJa3o9xWS5PdzA0kIT2HMEDeCaHK49s4jNtZYL8ywEHvvlvcYcrPIh
tXvTKC61ffSq7mDMF65/fL4w6yEBNyV5qupg0KEMznBDaDWC+k+qEcesBWJU
FQUoB/RYwQH6pHJQ+3aOUS8rzBjT9CChZOrSMEo6+FllFUtydyet72q1Wnqg
6c25c+CiDycOLqClo73e0mXyfs5crOkdjC45qmDlXUU269/KBOpGcfBZ0P4E
ciwOU7lbpU4GgajDxz5UpT1LjQZB6czkbQ7f+59ymjz9xk1hGkNYyPXFa7qe
Lhlq5tWNzgt8uY6pKGRGO4SHCzVjEjfP394v2EBZCyMMz7DhGnetY7dgAt6S
U2jOuY5UyRR6jutAuV53AqMPybsseDjK0a6f3MyVTU712oX2G8T1bnGe00zC
sMuNXEUKNb0s4CcMYNDgsoZmLCzatirOFEhYOhP9Dstob41BCj4JXvZPfymc
79k8umCm0ri0H3l3XX6i1CwnrV2gvHGPsOC94dnODW2COhhqSJdVdoK/YUOX
H2WkS/GA23wa1X2bgMdO/4JRTEihQh2Ou+RY92bBitWQb68jNNfUsCWoIo3X
K+8RCdyeaFz4tAFzLpsXvkkArYxLt87PmyQQ2UNxAhDQ3NuZrT4v6NucdnJO
R4siaota1nQosNjYPAp4R6UOEw5url00YFEA1B4YPvxz+t9YPP3/jHEWZVp1
Wu7L0G/5tLezM8U003YAeWm7l6WGkOnN/beqYnC3sr0ALY7m927Fm/OxMPk8
mPBD37E8KaA8KpEICc6ltdL/Qs5e0VvRT3BtXTipXHzWQlT24Xy63h687J73
tmEIJpP6X+kqFuJtTXuiTGUnt1GqoSJbqGygkEH+nhk004Mk/7s8mQP3/xGN
0NGwaxHzMk9j4/f7aLyXLY5owxZHkgMENzOijGnrBIsV2Vx/+caHpmdHjbBL
rInyONLD/YQZX+JLHt3OtBvvYI508Y6boLbY+dZ30J9F/3tHIH9GJmCyp49B
k7w5hvi0LjPxgj0i6bTUwMfWogRDKxh26qca2UECCcgdSlqtEDKnVpSCPmvk
3RLQP0U6CTBLLBGLkeyxnErcWDPwCAPkLvZ9X6s8P54W6aBUFCjgT+bdd5y0
D2JU+w5KkgWVayPTdKDqiB3Z5uD2Tv+JmFzWrkvQYmWC/BgkzP9pulOnuR/T
1ifI55N/l5CxAiICN3ZWLI762UQUoB3bdQpsu4Ck2qa1UxL+ix1vuXOU+SzE
BdquES+qYePl4LFdP7PD/EyeWHcn+PAy8++NFhGglZNH20FVko1G8rVJyEVa
yXqm+Vv4CBQH/CQJ7vA75K7REtXxUOEAW/xbvj2OPn06o+4eD59yVXTMc6Ef
sOUIVSKjOsnqVWkOpQ5+QOQLY1bvr2c6vuLG/nOM/26bexZEm3OyRDDvqA7w
btta1HP1XK626wvMHmpq7/h+2Mb0NsGgeZzjcsOq3ARSF3KcrZE/6/66gsEO
gFOxmRqjh+htSxSHLYUwdKDLXi8rdjquCxeobwyFG4O9oNNeX6S9sOefiPJR
huvXIWlAxCbfY85r27A7kmo1JgInB3Cud8rmHNrgpVrdX9SpfzFDBk4W9LAf
Xy7bPgVa4cpen73lz6L2cTQTOYZfrSmevY+9PPc9G8U+f64uXnEnp6tibQOx
Dyt7ogPhPGYgfDV86qsxuf9sTC7vlJeOWDn8yPT/LPdp2WBBhqkMUGwIQPUd
TTWwqWdsEmuKmqkYawQItvq+NzEiJ4xe6sHuEfbjoJlkdwZ9jHgx7xadw5QQ
1MXNy8aXNyetPWQeicUvlccqPGuDwAKLKNyG6U636SGE4hWSnza/sQNsXbdF
+Q8iuGcbY1ZYjdlvUJieOtxkGZYVFwkR38qFAkLWu0VU/yqkUJwXihJTpbH1
ucPyo/MujVvT5D+QXGWGLfItiVyVjKgw4qKRNKPUTwko5MJ2V1qKrpuHIoZz
OlMKpYLA6c7VgCY7O2/jZkxzqPlCgWCBUo3U8rlvz84jd1Fqrnell5RPPhEQ
Ew4w1B8ZDu9rU1eXV+YyU3E4t+Rd+k1tF/FKr7DcjTqRjVOI4e82PyQO5DZS
wsdPqQRTe7gPKSMRPxqHvfL82zV6xdIooClk2D/NVctWpkHWE+YuQX5jEB3N
465eT8b3GjYdr3a9p/0pZNWiN8UzcSe/KCHOfUFw8HHwb7sFZaHwBs2L7FQa
XdnV8fn4dL3kXhOLpDlvKygD6tuReUkg6wuyfONImQRx+NNbwUcOeRIDtuQK
oqalRvo9zHT95zv4JmkYVgRGVhLW5x8u9CADwwrLV4aAMUn+80Qf2nfU27Z1
LzcylGpnDK+SaS9v6u7cGpGvdQxn3MYTZpj2GaE5jaJJaPKF9op57vQP6euC
epcjp2EB3FOsVDzGQt5G6Ny6FuXgOOIUs7wFy6oi6hIzxv5bOz2BXnoFol8d
2/cdqZiAR61OUIl1doisYxSj6AVt9grx+Xlz0hMmzXwHWZFBS6MYLl4FkDk9
4dUS5Q5WTbI2HxjpAiuaLkBoN/nTvIlIrtSrRq7pn9FyKlXW7eUTvA6kPwyb
r7gDpFhLxPVOOzanPCsbXMn7z17xr3OG+51Ead/T6M42uJvkztCVJAB79wmw
anzAiv/TqIPwqjBxNB+UuiC2NWIDK34i8eyZM71Wt4L27cWrZEC4QhZVO8hs
VJ+UCAGIHaCSo5bkvBXU9eq2kMNpDsNZ4d9cFxPRhodL9kyLPK+hCKlEGRVC
or4IgYBzJqxnhrHj3WvStC3ThDPunI8nKv7VvHQ3Jav35g/Y31a9juNksbcu
nY/w2DOa8CSSZ3vetuS2Egm11IT0FAgBr2fxr2Ky6axs5EyFTPdcwZ9slmnJ
iVrtNtw550xqjBlex5mV4Vm090FqpS+Trh+x1LmS5wvenhVpOQveY8ikX/4w
euf1L5L1I2RcbxKpzYv/o0doYrgD/Mory6/NgWRQj6AcIHqmbhfY8VXufFvd
BB3sOAfC2FnimQJQNgGeiRzDBDEAS7976mpwT6LSuCyqIgwvezaSH39HoyLS
qafbK3C5KNFVhajPSENFgtdeaTp2mEI3dHe3hJM3pDry8JioC/xTLticmyRQ
M9p/LVPTBB1tODfPiYNMBPudlTCPJ7xD0ZNMd6eXif6aH8Uf/MhcrZeh03QX
88UBRuofQ8AhKq/uQ6YK2Wpv+U0XwYAUQB1ctp5NqC6MdLTaBKzEu7M1wATT
J4xP63nC4zy+hsVTt/h0XcStbroSEq5+qF5Dkg8JaHW1wRMGBqh5GcwfUADa
oGFU0fxuR/kc7qqjWSfe4dtfWmu4KrmzTZOkpCIIAB5lHPGy6r5RNOM8bkOT
W5RddNr9HHvQqfEuyP9k4wVipke5mXKWfC60TueRftdLSgcltXIxBl/3aeU0
5qWO+UgWWUfFuGhi4AzGk8ypslzd/4HoCCOyJRYT57cHPwTJvowhe6JXFk1X
9Pd59AMQN1BX6A5QQyQvBS5IzfWw3tmFKkQFDCEZsYvQm999+Vs3q/zb5x5w
DxKPPH2p9C/mJRKKGjoO8zoR9dFdPS4G1W9zvbvRelZnSdG5sPN7QJeINnfF
RehCtiwZ4B/7t5i6uN7sIH27EnUOaZX2vBXUwUVnNoaz1z2B97aMeWKQPKeg
8aQwGnLrJ4/oMmvE37Ow3+v/xC98zj6603zEPm84SDG3tYmm3VK6XRe9auNk
DIj3BK7oPclADHEqKzoROgGYcC49miUi8E1qYOXtWXsNPd6LqRdRsUJgSqJf
DwjQTDcpF1xW4enSbgZR1Ol8ooI5BkbNkRF071/MwGDgjVIbG8BOYu63W0Ao
YuFllwMB1cVsssRVWZV1aKvpRtWnpGHwzOmBPhemaQBH4OOTZZzDIIJwGMzn
3072mSwuYibWfJKjgcIsRsHOw6DgehU5VGDRBKltYKWdQA120JWKyPncRTpE
VosTNvROfvGt/NfOMoccnG6nT93kRN2OWxk/N1KHPJyu+M9AaAr5TJsaPSRB
rBvCsVpdx6E7xkMUkyh7noFsXroCBKSDC1rCLzm6FMNTxIyQ2Nf7OTiHPfv2
pgEJO1VB8Mu49LluJZaKR7YBM1ExCJxtRZivI/zvRKKvQ+ueXbsKc3hh8I2w
3vVWk9zdOdKQ5RRqONevhkfR24RreIyi1q6JYlzWjyb0CTsL8JuiDXLThWcY
i7+mB1HSNvdmNJFwhDvdg5GXm3SRcCsohRoo/bi9ARZ66Ezm9eZTMD+8k/g4
EpDeKgQlhEKJqS+e+8bHIicFmExInC+QG9Z6U9XhDAHWAGBrvyzhppQ7R5C7
f3Osptb0hwoyAH+yeGdsUH3XeqWLcL2xeZ3LcagUWW7fmFFI/3H70yINpeII
XlQurFh/kGtwFpJB9kQEW1GI0083QVtugfV79wiWyyQAPM+6OAuFEvEbqUQH
E35th0P2Qm1hsOkKDAx4GXmcK+P/2X+qut4W1LJUA/Y66vNTjZNKPeZfLwD8
4gEVGNSrkLfkoNcqqwfafL6+1R61GBWwWluNJzMW9wTetg1Ft5cSQDfc92bx
NNjDR9Vx9MMJBQzkWQiP9vy/OZRF2HAYySOmZch3/bsf1+pTVrMQ7zBKnEaL
kL89flSp2wMfk7o7Lek/1QqzaDW936SYu2GL7bseql6hc8khouDgDOiZPiPn
nASN7VrFToUj0ElXjAY0Zoy4VysyPrp1mam53EigB7LG21GhW1/ZRo8MaR6M
fcJavRa9XWPfFcCvI4GVfa+tQMlxkBrQuYI/ICuGs/fXqjdDGQVGKzDX5qr9
W5P1jMlcsgs9D94a+igj/Gas/6selXb+bWO/AWPJgOqMu9JLK9AAp8n+t8nm
XgPXNqyQoefucoTqxi6SohD4MjBStxfi3C7iWrxSWbpC0dL2xnBv6WHQq65W
SvTw6ZMqA6zaxu5DhbDaMbjFCS5XEsrtkAx52RD/ZglGr/ZlxNcxXwsEL+OY
QPUU/8Zofb0o0RD86C3OWNUw9N/Abv9xF/Hxc7OWuSeGsRmHHHDLEl4Ioclc
uTwgf2ba2XrNRvZ2YkkvYd3r6IWKdfXgZKaipVwr+JSXXXcXYJwFU70/Fjn6
xGV2643t4BqSzvZvex/9DyFna9oXvpl99fil3GWcn2UPCQmPlBvJrnKC8L30
YZJtCFzsL4gjhGjsm5f284J8IZFndk9CaaMtGvX4Hs+BJr3AQLG2TMpH89Ug
6HuWSaF9dc+VMfBn0er1YGFgWf8riTTe+OAcHmFL6BBFWC/mk9EvyTJtuDVd
ZbMKTXrBITUKpmjcicQMrGrI8p0bj5Ny69mucAb00SRlfSXahg9rC8mnEJw+
LlfN4JDFLEXY727EsxOzTrr8MX4fWxfs4iF3S80WOZO1lq4qVnTBwrEAEkYO
9Sw8I0ZCU0f5zJYWRrPQgKeXXteQ/IWjPfuRyZP59e0No4A2jySnEqZKgcZP
NDpx/ypneU0C6jgJ37TyLhnBhmF6IbnZy1QgkX3r2kQE8j+Yp0/mKO7nRBh3
PMANPui9MJVGLHqg+1uyi5Lm7QLSKS9SfTceS+3glLzyfWXosgEE61kHrMOw
k7sPW3mFP8RfphCpA0OAyaWaxZ32Z3sic6CPal725HZNsY4F5qNcCEc+fYkh
jK5bGA6C4r+M/DOxF5ykQ7NMAhlfcvFPobR1Mn2hfMOj6PyHr+Ll+2pW8fCv
3WZ4dd0AWxGjFdYXtJt+QStCeDb1uIeRH/Ct+RbjNTTkJ5zImGKfmGw+5cY5
fWJ7QmdiBe/27x4+FVrMiRdRyZ0LvC//1ZTGatbm5AyE66wEWUkMbm27yIFY
GZ2HRVTQv77ihz40ugWrxA5aDiwZ1nj+TaxUN1kjgOxl/H9jaavKP2CB64DE
2IDRwz6wOTigAUP50nvweSSED7ajdBqVS0Xci7kAPAlRL1TudUgIfffU/s3D
cmUchTDBI77wP+xZ3ejN6MgrE2EKhkPrauN4P9jIT3M2PhHDf/9Ko+WugbBO
rPQkph1GCrcmAi7Q0nHtKRsDK9wQXFpkpoh/wCBF8gOzG6VhuryPBlSZ/iFa
lU5rPT9NNYFkoHpBBFmHxK3xCLqi95geJedDzeXbADbR9/1Z0TeS34YH1R5c
c829h0YHzzMxW91QFE8yH0WP8Ee8UET+LmRz+tGSN5naZO+Te+0iXOE6wD3c
7/uCsh8uRdu45TW0tB+TCkgEBXeKRFzld3Mnf9SiopvS8sbO06+07i6cmV0R
qfs8pusaqyOAugQqQDcZgGRK5/wTo6mbDDQyFEHqw0NE61aT43SBZGHHLbtY
xqMxFRggS1pzCMSIZ3tMyi2ONudR9wDKF6y3q1gsP6Wy/AS7n99rjjb4Xl+R
ua4clhbD7fkKWn12m6wUoNeA9JeEArHQEF8bvuIsesomUgakkueV3acPUFO5
DPwFePm6LTyeFtnbVsZo8+txjNRF36RiuCS5GunPTwPGcuoPwclRbCEVLx8n
11xvUyCdJfg8gev33OuavkFK3Wt47Y8Lf7/1SnrVLxB2omqXV2JFLrzlXSAe
85k7kh5p2Nipo3AOQshV+qRnb34YhPCFramYAAkY5geFHz8H3zyhDBIxsmCM
2HeVha70umE0lY/e/B8J6xztj6t9+yNz2yuWVB/cjzcTROp+Ahw28DNoICYn
32UZdziTVDxe/PVTYrC0CYPaWmAVbkD/MgdIlgknr1+LklLR6y4K9Bf6Rxe3
LVBUwepVjK9wpn4BcrdN8gIsXNfnemwwrsI82zCS58I+GYdGCDhdaKMU6v6e
ZpyOS2D8sG5sjoKwR46aF1WiOx5XLgEQukATwyy/7TTy5No+MU8WY0y/5wRT
gQPIAeWxk9d3gDeaLMCvQsP9l15QSQ9C1G8fa9gzktRxgmNUFGCzcNDVkafW
6Hbdr3U2lH5Zsu5Z+nUd+rtS9Q8c39vR7s2+aTCsYUyGBd1vO1UYwsJ+1bc8
GD87RiXzV2BK5eQwNRSO4qmcnfVFKni59YX3V/qOoS8jVO3+HaIBjwyJTtIH
clsh8WhydCqPs3WMtfrmjetpzUk17lvBtDbw2sLqbKXNOIewE4Zy8B88vO7R
xNKx42KkctCQgc/gHkVG2CdwKhgf41gmoH4XpSTJy8MmAiC2Nbl+V0onkTQT
aob3IPVhlDxgA2qgBxFo/THTsxOCvSxKJjvZmhGfsUNrnbA+WEKA2l3CxUP3
xxV3GqVXjnBmxTBi1/Ik+F9Ul434gmfQ8NkSwdX7tEcdEXS2Iwsin0kGJjTa
4rQcYVmximDAz5qzGeWD4d6R3cHAva7vnGEqxAluACureavtahb8U5dN/eKw
Z1uK2hggn9phgJh08XB2Mz4AsZK9uSSJkivUnay729khiHLGhzXqXYh2SuwS
9EQaJkh7La+pTKhROwoILZlilXKjpPVVp1m2NAHJiFkvtJvb+Zp67O3CPDW/
n5H808n2aMHDxBaB0QXyBsvm0XV8477m1QpAD5rEetVyIedaLEIvemsP/51y
BOgDj/TTkjEcuQ56JqLfjRRddEtkguB5GDnFjPYkHezCbqjud5Yg0uWcTngl
tamn/VmxUNJolhqIz7F0hxQoAuuW8Xa36rJtBQG51dL7jEGFDxK43Zb5PmHZ
QQjJYIFyt/P0M0MYBA4pfi/VRRJS7lHQ1kW6JwhQSVTis5x7EGJFdF4gfbBW
wYs75z67bjy0XeiMSrQdVfmDrwiwsD73FGwNKLZ26Sw37X8tEo3igmlRJQvT
7PljLBWFbJkSslNGMzIHDytwkdzKNH0n3bW/dDR7ovXy2yXOLdL44F0AVcNg
l746njKsmwo6DzAweO2hSKmCkRilNtq3t9YRCwfLy2sYnc37QehKbuNuc7EY
gUzKcPEXtGljycJqFO0UYD1RHQArmn0K5hSc9wehNC/onZ8zEZE5rgPMZa+R
tw09lRWra3DrB+OZGjJsW/+FGmcBT+aE7CY3mxBi/xkm6yMjJvjm+yibKX9c
hmrsATeS9cjr5VRypYCmRcaYHHE9cld6kxsTbdxpm340qxLxNzTCH/yCnXFS
Qvo+ipDGIJS/6dGHmcQZ7wKOHDthm2hAZ+8Vm06Vjv40rVVYSAqagHHnaqgp
+ZkhGiy4QfeUChlpxZvJSolOaqFKokJhEJfZwoaDY4Q87+pAXAh/KDYY5I1f
Z9S26NHo/r5cT3srP5N3uSQwV/X9LG1s+qjsLBmWWWBFNPk/wzxS0DaYpUnk
MC1LPeFmXYUPob/WVEnDP4VrbehEf/P3pOzPUn+JwOosuobw6zIAYnTVDkwo
Eatpda4qSYtgghSaiDyLMAFsXSEjkCAmJYnyxlPSUhOV3Yms1mpQOR53XJXx
adHvVwBDj53RT+U/OuNViEauu8wcNWmZvnEAdHOrfobGObmW76Ug937E/iqC
28VuUa3tjkUOcgR0+oFx5vvfqib/sLZgEIZFZogCJygnekeaeTql7IVsf+J1
mPjfwZfBXA/GfqwbuSTGlgr5sU4FvDV2oALNYDfbR6b9LqK+Ufv5rGIGNYbE
zEldcn7Cco8QkmG17B4laGmRrhW/FtZN12HZFcGYUPEFQUIwMXnKSL7Acag8
K2tLDMcteah/NM+VPOJco6J/j7FJq+HoBQ3JLfnXWEbVtP6FgzmvxkybNq2f
hr0y+qTRowliI51rv8hYhLgq4DyO39btVwECuBHDnRMtgFrBan0biKSMvWbn
SSBVF1uEgtH647KL47qGSlxxKBVkj9kC05Kqq9CBvs96HZlk/IjVk5dMrlI0
LCvfVWOjfMuyolF57Ti3IAdUtb33jJsGuNQekMKHiRoEDOG+XXwYujsXGnHd
ooSfpe2ew10cCoHKrW1RWy7cd6AztYqVoKfET2+9t7UOycSiYeC31hn2Z3oN
Q7rZKTuNrhCl7SwIC+BdUrACJ2UHJjpv9Y/OOSHq8n983kCTRzSUTDJLxaAM
QKDIHvjp33hKncq5hz4FUMtoeTACVkEdTADuCFgzLf0zs+ylIBiLzQEZvMJG
7k0uOiTpmpEXIbolDVxQJb4ahEXy+K4x+ijQ8v1wvDNUdmHTipq/gEj7rNVc
KSUww+0Qu/MqJArpNYIsTSorl5zu5+kOYsdwf/Yi0soQfYyrCBoijQ3h4IEe
UOEJo77ipgvOEo+zU11RvroGZ2m9xiul0F0vnwC42W/1NGOXacCW/NWJPQhK
mqLtq+/tylRWU8Wmrqczwh98vVRpMxOgEbm/G4Me4FHWuW+jXzcKTl4DIHm+
jQEORTwkRMORWKmFpBlSjn2XXwIq4l513qlNqK8gYN9X9d9N2JCpIIy2kHp4
Zl4olsNRxqhFvthr7LcUQx/3DQ0WcSGzu8ij3Xgu+8993Vhlanar+JQCErcb
9iSabbjRYOzm868UxqvpIhsaMwRbYJlBaF2EbaWWegj629YxM12Asx70bcMw
2Nug2KM0OiiyXnbTm/FjTj2YlZQnY+93SUnNZzdFCPXCLybRPt4664zDSWvm
nBQfDpAjWe+9ufd3D+Un9DZ+PjgDwTmhoqP/hJztbAZgmZM6DiVZ0d1Ly/3Z
PRMs3tpyB0bwzzywN+dUcL/EIblIOCoGkFBUgHp97wTx07Dilm7AV8LBMiFK
siUMC6utRNO7PnFv7kp2TRgF6XD598cPXtC5B/Uc+YuvSfvmKSOT3wFiJr4P
FGQTE3hOHKwlvkEFD5DWlsKvB15/67wr2lwN6oMmcs1J/FwpjJV+LgZRxxTS
7gRwi9aAYYzu7VID+DumnF6ZNL7W+Fih9EwBKiNUaBvhplXZnR9RUsU1IOyj
vS1hulmAwnlsmrYz1R5XG5EWNAETOJ0YZ3L0RxaE8Cvc29Hg6GtJtJQ4DcE+
SW8ocx0lQDMTpF1CAzzDiKd57fozUO/zJVuaGX6+gM6RiCbkQMsCEimyombh
UtZye/+EnICs+VnY65SuFvK03WZz6BofUSHa2JGz57HioRzqon4aJ3QV4p2H
UeTykF7lGNMB25FtxshS7gVWrwlO9pTf5JiTB/I0GX5xEtIykpCE4xTTEc5t
GCxaDqETIKfguWRVNAYLutaUs8ezDNcfBkIAVJpDxmU4MScdZx/Db/Fo/8dc
fvbTgWlEa3gBaFQmg8f40vUjg/0FypsG9Fi9u8Tmu1Xh4lzXN3QKc+Ip5QFq
Xn68vBTDtZgNv28EO8WWxcYSeNSo7VZ1eMo/LW3ofMIwBOlDzzQDSo7oRrVl
/N/14qn0q71ro9Aj82pmyCdRZSPwq4pRWJJQj982tJeKzhrXXjZYNP2nQxj4
W2gz42vulCml2IPLzWUpceA2fbDwELuqa8OTHcRnn6gB9nv3Be243J9KejDC
dzPcA4OpZ0tY12tqhOo/RTXZ00/Hr1LD9i9SIb3tmUEpx8cfBPSz/gKmhUiu
u7Scpc8C7f+C3Fa/DqJc9+11sdrtVITzbyrTW/H8hQIhnDZ1HW1nmQl8pSC1
7qmiMzzNB7W25X4C8/yQW0EkRARw7sI9ncC7AAi/r94FHZdMJzGsBMz0dE0e
o1ZNdqNEp+3VCyI9JxAz6s106aubO87sO1AJpGMqeQT5Kzh/IiqWnfnLPDk8
gDrhTgP5mG+Lzpie9G384ibt1XoQdjmkEHfcRcyKmKV2Cg2XLLO8Kazlnspy
r6vzOhvzqgjgiUh1gW+Homqrl4UqZRkOail0hG2IU8JLcZKk9jqrtlz1WPnk
vyzcLJxHNLQKMk6ZyTO7PlK8GPVOY+UpVHPpkOjeCXjSk5Rid+r4U3cuA5Op
4R8jzJbbSgdTZqtkqsnjIBIjLWIikgEv4SWEMMdRWH0pnUsTW7+Fl1VPPxIy
5fXrc93q6bnTg2YM5VWDjKnr/iKAn93m9ODyPH8H9KY/EGnVqmjqXNF8bJzc
T25mmv5+eFjTs506BsevD9Wi9V24Wv8ZWT9fyA/o2ny580yfLtnHAMyUXD6M
lfeSot/oIQ/RjH51G+592uAyi/RuOBu+2IurRazM+wtO9Z+I7bH4NGgZJ6yY
xhJy3+BYTgy16vLZ71wObqSKhDSfc1BbaXxqAXFwFfGBnUaREU1h6oDBFlz/
2llOYrE2nE61zgz+b0+hh0wBBIWnjS3DyhJz359cG+/eryMNOX9E9JmnZOjD
13g1PSP0DU4EYSF2al4ZNPb2BuSansALZSdGmJr47BVN4fTCArRr5kC7g8o2
IEyNwW+Zd7ZP+i5X4w776q51ap7WmsLsvaWLQNf2U31mi2NhgqVHWRSHBkHb
1tBDOJZ/S1jkSBknJd3P158ngBzSFxnYmEzsYYobIpdt9cdPqPWrPLF68Uxq
0Er4/Gm+D0HLsrkV9IFQqUyPSEgPoefwfLbabn9l0JPFQfUdaua82e9L5UBT
EZbemJCpSoJiqQPHhQLVXzQS2JEu1DbQ/WkQtyaRW0FfeUB8NLby/qOzhof6
YiZjkQpwHInDew+uk8QoRNgqcCSXJGFuu9uUqupQYvlcWtGmIE0bizPX0e/M
obAEPmmhYQwKTMCkmmlySlzqEiR85pYrRV6fQMudAJPvCvmaPOkITthPH9b/
PwsmJivvP0a8oaMSTWgWFgPOmOe1BJIDNS0Y1IDVnWrQhTGd5HvAy5Og1AiV
9yV3iVnyGEWtwFFlMmNLRYBB0WPSX+4KwbmfBl4f+uLL5+1opbQUirRmuCJm
5CD4nsf9w2AVRrNw3N2hzC7wafTU/8aiuy9KJhOqDfzcXKeVZpQrOf4DoPQJ
lrAsjk0cwDG6WhiADrcASNbD/I2AHjq87ZNaRuq4i3F+TfPs87o4QIUG7VZk
GOT7JkiKbKMLh9dA1yO3LmZqzIKmiuZKVxpy4cTsf5Z6wRZOX/aCOh0IbQt0
W4y7AzZ4aCeMHftYc0nwWIs4q2iRfBFGp6vAmJP3FgFMScUSB5bb/3447x+U
m8BTfjvNVx/EVCUaUcvh16PKK/kg4pYgCdcLn0OxMnKmVerFNE2k3+YBBWm3
Lq8bIWwopGMIPI2JvIHml/wdnvwlYyNJ+R/S6FjtkNAQS18bQju6e+OXZurj
UY2kCMenkkr/wfJwo0pEr9crxJYl5SSVUyXhZhEvvQn50+aVIvjmcIfZgjY7
cCyDXLl1/7J7nmMVx/14QbHYkM1ZJK6dc7R6SS3Y+kqVjPODRGNn4pRPxkAK
NpPEH3qvWUNDdcIFGMOaMpIlrDxx/IeSOnkK3NV2BpBCbRro2ZU+za7hLaUF
Rjys982t0KLteHvlm2wUNywAP0x3sO4GdkYQYh0EwAHQPEfyFIRGcFQYdp/G
Zbz0SFdcvHDElFmwXfTemqF9FbM7tzfaE+77xCTYIgcB5VdU4Wsi0B3QVNKu
aExVTCCc6BywQ0bIFybUyp55toTtcNb2RN/E2fv20p+R8LyxvUOwPdnjKUtX
uZdw55HQEiBYUDUYnzHALdxvgx8BOdREVLA4RmbshM4jKtNd5E5fYA7dK84q
d0apCkHLdzqLR6fv59EL3BkXBuagQ4Dqz1/x+3lMkTNZdScheC/SmsbcOsx3
aGuIPBPLZYDNfMCHcLfCPsbrmV+d6avoK+JUlWz0zHL1KxiWExQUIQL5UiGd
Y3LhN7qBm7gKwdOwiEorx36bSYjFKvGMHLB8OU7SB0guHzbpdxir8v2pRjdY
SNiEsIze3fiQOD0lS+OsF3ioaN0dbS2lKuixte1RCzce7y9Y2cOY6ScZiK5C
ALNFTeceoxmKJHc5+BQu7KreFBLioygAXUMNNHsnGP/WDdUm5dLk43EnJ6zi
N9IultjSObAjjW0+6djxYyMvom6Vptre0TUZg9TgHudz15zzflC+qvSikaxG
vDZVK9aDy0IpmN+Oucll0NguaiW+P2aqnwbIzHtVttcZUmCacS2lNwV72hCw
agrp7hWs0v8Pq+2DewoRn76ZhDBw/cGs0MjJQqk/gaw43l0sh1Ox92fF03jA
ac+K1LKEIi0w51bMjxPSBbqJIro9BNpOnhc3FnnBw8DSV9GRMXX3vG9rNDRi
ZaNwjbzyDFFIkW5eESh2AzswXMfYRNbK+6hcylVnrMQ6sg3WNCLAvi+aILB1
DHqKUhUr4dfBV8+w5LnGkNct+j9hblmakcLFqYhHR3tGZtXwFtgdRuFARy/T
+X4uzaYCQBUWAXfX7ly1cJvsCRdYCFjYqG8yIxGvQLLa/uN6hroehAS4qsm4
82xZHtr1jjB03ZbAo/OUOc92k8hdrJ8KTEMrCVIZkupzFVLq14C7gezn5hQI
vBLMxgMHeurYwvwuiLe06jJYZf5DTS3U2i98pKud5cqezE03eLMCiwwAgVYT
wXDdPl6qIdMC4UNpwgePOb/NE2tSHnALu8NBIoBPlAoSq2eSejnqcBpmH5Hl
JF6E62DkKiYbgEWDyg4x9obeQd3BkxXb4CtM7niy6RqP3iJEWVHH/3X/lJuK
osT+H/r5DnjoHOrgwcpuPmhkaQ797IMHzJJ7S+eu5Sg2RF6okKwRKtZcusUn
DA25KB6FUIeTek9BHFsDLU4TtvSKup2zrMt/GFEnBJYE4aOgM8hb8b/CxymQ
J8EMhRE0XfOdwT2c1t7JYG0RpWOJtOAULapbSH0VL3OmWFp9+1w/AXJARWOy
MdpRx/tdvSCcfqqhXwBe0XQQHzRyfBeG+f+cMqjYo9Uxf85SPn4KgWgVkX0r
hFbw3JlM0RZaw7rryaeJzXB4aAXG44O00NLBgRR6JginYmU00l4iKR+pc2gK
0/Z0NlvPMbYGEfDWRUkO9DxTZ4p2L0jNU+VbVhl14FUmFwo1vl8OOxMw+bp/
UxIQdI9VX0jA/8UKuV8eG81pnCsLCuTmtjmA5DAhPKwBiGeNwxYAlpkZpBF9
jn+6IbhGHUXuiCEwLLRB1ufW7zQD8iu6JGzjcQNetFhRCdthoOjgCrZNO4R3
EalTuNREieNTvyx1rIwIO6TO7kkGh22+adr1EMz6ISE1qMyapyt6TsjnjnnY
IG4lylxPLDuygUTanxJQtPWGb3PSLdb5QAhGOlUGP30poxbcbDv/ENNsb/TN
I0nP14wfBWFqpCTsar9x/yVcvfpIIf94tXJqxi3hL88ighJcIm/4aBWW3GxO
uMCfURLrE8twL5qThYna0J0vROf3v/Jd40N2UMVDk+2alTqaHRb2sBQwP14t
0rR71eM5+qEEW5bhFMdwadXtUYmVeU87rYZrm2/Bhpvj3FANck9akSJzbU/5
CLaVesb4H1OWptHmf4AIWuWhi/cknGKfwTmkpOUz5tieoqYnDJMS8Lk1hGTK
LfM39u6h3ESU4+HXRk+hwYg+TeNYyenQzKFTOE9MSPpAAxvi7Y1UWp+ZhIwN
gnwknPedkZs7S6UZOUSBi4H24+8Bk0KegpyfW5om6EgNik7QJmR+fH2mvT0D
ydpUcRvFcuFn9fGK/e+oLUQ7mpjacdi+3HEqljr1APObG73vEBjwhOe4e8tI
CjcOad4t+RmenKm3J383EjyiJyIvAHXFijpNkvIYIewdAib015akSKaAVbMS
Vw5Jvws/srhnySWzsLn4ClI7c4bziMXzGSl6AeMwfczJHRhHTeBsvCqp+SCo
RBAB2DAmNFCBY2W5dsYnZcp061hGYS5siIf6mnY/vMLSuub+qlfciRNbKWSW
c4N1j+t992iWffeJ0Trj2VSKaJyj2UeEdIQ2ZYn9xxet/2Fq/r5WmLacgElP
cAQV7XgkPZ9auHwNaCMjt8t8+mQ8mt9cJm4AIkHaUkOemDdZ1jKhOACdYOmL
EQLKqTZb+33BbdayhBtgUz7zz390A7KHnNx0tQq08ciXd2makoZkMojC/7vW
OkbDK3N82LkzcB8CWA/Fvn2nzcHKyeGoA9yQo3eS3nQt50+fDYT9wQZx52pH
rGU2zKVuQ1yzdkAzk2Awwz6iDnhbrgccPV+JAC42GtJubd7QjUWmM6Unt0Gr
mKhiN34G640HQmZ5mh2W83+St2mxHqevwVXBZyIBayjmizcMnlb5k1YB2lHg
QwZKId8QWJsdkVBSm0AfJltdxAlSY9O+1GV+ViBG6vG/+/9rDuciSFx4xiCh
laX4d+svKayCbYQyPpbbUH/FWmKJ0TRrjGlEOg3C6nCUWbem5GiBTgYBk4lq
ZZ4MYJ4k1vegEkF5x1mpVj0w56mBIciYO/ZhC8v9T/vr23ET9ZkndePAt9ue
AmV1/EKHX3q00ixGbJSYiCu3ag8bPr7sQND8WEbnGstJvendbU6Fe3gfw3cC
fPToJjK4TCqapTHTgq8EwfDSFcLx69WojaEn+OyEmWX9LTA+5TJi4W/NZyAg
CJoLA/6a3UiU2yxwhzsWORR4hD/tsc7R7UIjFSVamiKLmMqQGBq86MwgxwT7
FjlLqI4CK5cOcObSALfZUcuBU2Q8el9owB8lsHT4usg7rKMsGp9f+Wrn+V9U
EWF8ZYeRNcxA0K2keWcC99v4l5qqwXg1aPPwDfTYy2O5zVAWb4JhPttc9NQj
vXLkWO0GbmR/LcgYms4ptMGbX68PksJtO3pWwD2ES1//3bV+465gM+hdYKqY
gGZs6IDezGfvYlfjhkFB8LtgdPZgFv2ngq1+ai3tL2UMPn1PXyzoiITAVScS
YEODyb8Vu4CCHslJ52PkEfTm0GWPnWR6YBKEKl+TrwWD4lJydd6NDfaKjWS/
RveMQQM/oG70LNM6RiqH0RCucCvVu39BkhCxwdbrRvPC549WFcn7QkfVoIT1
cbmHUbZAEND6z/AmR26yI3qdfoeN3mMnWkRwZnokTveMKA7AY5bh+6csTxUE
MuZXXmY5D3sBkd1jsnpXmtf3FzVg9X45cSL34WZdT2rTPmEf79VJb2S9BW/F
Mrtb4lTVHiiAgNKecuYlu2MqOs8nVh5YY/mVd+Nw7IraxezH7+/LOFFNzKOh
CTMYuoImB8Usc2zEoTC8wbjDJV3F5D4AHGiKPOuarUaqCFJ/rLKsNScH5QMQ
c1IbMNYExTZ01HFDXyC0LIRTgC5fFGFII5wHtIS6Z0XS8cE1TrqxTJQM5D91
a74qKaicQU1jEYCgOuGGFq5NE5Ji6ANjMmy2yCFOIXKzjOQ3BduDuzjZa3OE
C33QUDKL+B0pwQG4vQtHRTduo/R6DM7EJY6EhYXB3rN3mQV3Xy+mucCMpWV0
HXH77vQ4oItIxENy1ASge0P1GLzziUI2Fpj86j/b74EzHmbNAd1AJqN20uP3
ra0OyQngb3Q/ozU36tgt9DogwG3HH/ucc5vlqfsQ4vlM9vKWh+0JnNtoUNz3
I6EXsy8kk8In+pNAcqB+itiTzM0xq0SbPJOYWiSFADtuupc1+/kXSXjz5XXd
fJ+ZQ8jGpC7PFloDop0UBkf0kVgoWM4BAIaLT3EUPtAipqAtuIqZkw03w8Un
lZF8QWNIGHuJoE8Nhlut5h4bMcwq+LT1T0CgED+duZ8GpkX/uHXYv1H9Xhgg
MoCUvGkrLtpikbG6wRUsewLc1S0AdGqIYa5+u8FLahEtArOf1ZdsqF5u98JR
rAPw6zcaznSdZTq1JPF7Kwt5tr+SBXGeZVnV9gHRNR3fyrzslWlvVj9f31fH
6WXKkXPg9/gAa/72S8tdvTKt6utPdRT7s0I2MsCjLm2XGgYntE3kiVutbdrp
YVqGkDWkAhoNvd6EtUW0LRszU4ZsU8Cs7BnuAY9CfYWP7cJszE2FWDTE7gqz
+ZACx6Lxuc6FTvh83YGKx09VZTWCtfmKgncc5cXK761ZPDl9ceU7BzpVfAvL
QH7+zIx7nuR5b5b4Uh929gm2WU33gv20jn2qwmJfZ2ej875tkTgmF5h/ctsx
I4n+bJjTzj3/qoUvjM7Ydx8EN6w5C72tP4lH2yCvoJ2R5Q7Rn5YGQB3e/CbG
qRlYr2DEMD1/FVFww88EDvdwiGVlLCcH9bTX+m5bmY2zyqlmslK7hO1ScFsE
+pkFmAIsbAGdycibq/iIInKhveW3zz4ZLf73i8nUISScz4NVt0CSq3+XtMhs
WD6/limjwctzz1nLz6o1SDPhW+ORE7SHLB3FtYQde3ObNl8B1Fp2sEin36gM
W4HhLdoPSgPuWz+vPxLeueJtU5VZWnhhZxpF2hkZNXbqUsvygOfK6Yz8kzz7
dZ9lXoymIj8naYIJIc2vUi8wWSQdJOWbAKxZWsR+muv6kAbiWbNEg0aHemYx
0qUjAE6rChXGDFSuyK3shE/ShHlZj69VdkmWBiAUEjfZrqCoGWFaf9LLslE3
v8XrvLunnQhcoSu1BkYVUECSkvuE9GEsvBq3HE4BRYYK1xtA2JCxcYAPOM8S
5p8Vgf2bezpWg/j6d/o5uDvbi3LmIEjavVIXIlzoCo4S+FKQyL071ZJpP87B
O9wOK/A9w/j8xWvCemR+4CzZNheB96+bXhKn4wTStC8ANifVlaAk+OO4TjxO
2pHqtDsnUOTVQ6Pjirgdm3lqSdE0tqSFJB4/ACfK9zG7tJhmfoKftGSV3MDa
T+sPyVO7/JOael6Sk0t0m5YOwDezNjnYTfSZ5J4zS4I9l3MlfrVUfI14trV8
MteVmR9k5DQSHzpgl4CVhr3Ph7QEwB2qRqGovQ4/fBMqb1+GOvCRxLwTdYwI
z4cgZ1FOQRwX7o+HCNM4Cf3l+LPFtaOCw8LOFI0pCFAd2L2780qfExrvZAo7
wCICwvUM5tc2y//MHalHn2HES8fey4uKX9q3RS5q4LejgDwh5ub8EizaRjUK
IrZrPqrSKNzoa7flpz6XAQ3ro7gxpYQRVFEv3xRnov/uxf2jjSCeSu9g5it7
t0Wp6Szngz7q2X6yv9+6c1fuHDUeCieN0vE5RNKmr+MK+m1r/EQarOTbvpXc
Hdo0/fcUlfpYhQNgqJpGJ72LCHbi3tatt78sgtq9E/pTcz3EN12tndBzVADP
WGvtsTGikl6NMDJKNQwk6gyz/J4YRKXioweFzUKk5vdqry9s8SEqb37J1u6f
1d0IknpYXNjXT/3OdSx9L/Ym5c4tFK5JtgAjPLOwJZnudgLc8d2iGI6LP+Cw
OhLPF9mZ1ShW4fBstByBm44hTLnVZpdQgNcY6qh+AX4Jm7KZ4zh+C/ZcTgpT
jVNZAyTq1sTbPJ/VJH9Ao6zVcGXskr3NNog3ZcGJn5z1CVxN5nwMtIkp6U5/
l6+fheuwyTP6xMqHFyxgsSeXzfXE0Qm44pAswKxwP2GhhBDY9D3uQlo4SOD0
03PlO7/6qRoE4PVx+F/oEQ+CaOHGLHHtNJzVUtv4KXhVf3UD4h/xns1NxneX
C6+sQ6qBGw0q2fz6WRt18HyW3psX1RTyR6aXB7P5ioZz8RZbpbDrldyCmA7I
giWteuDzhx35uob2lrrHNbvo3aaf94nxL1adnSMBxNBr+vqbBIRNlACi3f4X
nU7G77zOM8MAJU47kpiZYbkm/2L+O+XYl3iZEL2krnLLjHO9vkxfqAXvudwd
n+C+3MXTwggh7n4hp4oplc69qO7dG9QVJwTr0zKHf8AEd995stjPtcbEbIcT
NHleilyFwTvpDq5OBRzuAQ4nkLOPjk0LhfdA0nUOet80O+Ooug8CC0uLDR8d
0gN2QSq6oPqZTBack/ifaTcAZsLugWv8Q935YqkdBj1gPOTQWeKg+PLKZoOt
CZfvqe1W16tMgwJsNdw5bvZYrAs5ORZJcLjhCf0amxeHjqHnnL0mGagaGY3l
Maxr5tdXkHJi6wVuvRHIzmv49lVrFpDTzKu6V2SE4Pae2u1dt53loD9xoCOC
6m0rija477K5oum1ZkKNSyK26w9LJrS6mRj+fqV4mttRV2rFwFOVKptd1zbX
bVTPLmTcP3Y+1bXOeEAbmWxKF9oEW/wVYhrlUeNcnefhhbNJLof4Wd7cr013
R3EsaUx9Bjz/0P3XqVdgXhY4phO+mTgMaVnhFSrozFW7vvlF7H7Kd7c42Pr/
p14xSriIIarITZ+HyovVXfoLXYLf4vOAnUwoVx4rwUfLJgtd+RB7xH0tiuOm
b+C5evfnnF+vb8KzyIwXUpo96jvOTe03Hkfsk5knA4VV1er+JXaWTFX1v/7p
RxaLHa9Nw5LJRwZklBI97Ky5/LLVe84n3k7qDYZl054Cmcw7r4+uUd9ez2D3
nI2FzwgrqcJYnYNLWSxCbLj89/9i8X81DlcMeosx8jGBlBSuwf1gzFhr5wOU
4+52h7UKUK4+pqQsRD1UywE5wus5GWvA3YZbem8NO4VzPnjZ+Gg4oMCzdqw2
GyUo9P6yEvYC7Hmc5XnCcVWLg8y+YT9n6BXnDUSjQSLe1z+MpI/uPR8IUCQi
Vm627iwQpQ9wUFeAcji5OrIeSInL+IebnEs3sy5aOuytpNds3zoHI8jNz7V9
HoffFTmd2k4sAug4RUQqlWqTYs98TLMt2xvIAPr989rFVdHT8Nuijc3fe1+Z
jjDm3y92AWv4cecGpciP/2KC8YvHovX+SU8L80IkfHErUkZIJO61QQ3stbPs
JAmoht0eK4JpDratAV9NFWo81zNr51B4zNWt5iDwH/wZC87+cq3Ssui3jN5O
7Tj8KpoJwaoRqhpiOCYqhhTlT+R3gGJD8tM0FFasVrQ8OwKpFtimw+NcfpKX
JTrP43cbpdDIhdFu4SPCKA1TKdxGxqkbPoacFGTLC8l5UIATyeGmx9XyqVuQ
9C8nx08JPTl1ADxxp79LRmnQ21M9kfgv65hOts8gAcAkUQYm6B6jBzOBNiJ2
K/3CLZ9nZZiooKzgrNScdeqEGSFyKDzgzvdNnLz03D3oKqa58C+Yf2cIEvGJ
1+fuCa+5x8I7rhuBFJ+vqtcgWwvRrFbr4b5sABA4FrP8kShdBizTmAKLlokM
p1R0QSLoyuHKwpcUffNo30YnlZkl9cr0uy7ojxrIRFWbturjrKy/5UtoGd9k
RLUePI47pS4LkwvEH1ODAivOMoLVNIWXCRQWvibNnmCYjEdyVGiW2KHNDAdc
GVOwvrOPObs2FSgAeA/WTu+c3MpXzcVUCrTDAOQ1vg/eBrLBriU3cWdWb9Nn
whGX2x9lPICdWpGta7NSK7RYoNElT2YKrI727pmpdERVdB8k54rb/eLE2KXJ
uaW09uorfA7kvzdidtER8ORX1Iec3RbgQKFzwvfEWbWoxlo1QHQrUiOLXBAF
zc5kyHpXpwdaSy+JiXgcM7iDjg1939K14BBl8rrPC7RbkdRmBAyao5dF3XCm
C8GePXQylIQLm/QoLZKqmo3eyroNOKd9ADxT76BSsVTg5irAWHM/7FGw3nAT
YLFww7S3Ttk8vcjQoQfmuJEuCWSiD1Q13JcOc/V5NyxFYy8FBBEYGwXQrmSK
HTj+elp9ArLjEmQNMw9MVZVuRdTTID72uDf/BJpEblSwrM5A7iIBYmgkUPwq
94D/5kNnCNEQpYwYnB4Nk6yZH43TQHDbMDLZrPDEt08OSmkNTRr0Jbr2Prtz
zK7t0g5eid6T/wVYaBJTd8tZTdpDtUWnXTfbelJSzekMuP/3R0EcfPgvmMDQ
AaAMw7GZoDiB1XTLVzJ3SITEWjwE+m0f6PGRgYWwD1M64NMn84zw7Dx0U7KR
EalZjNR2kyQXpk1EbZX0YF0SivujrXlattZ2KAIXBxKfPOnx6lLdSa5UzGwR
+YZqAAgL1bhcqRbluLC5wVbwTe0XgzjK+jtCBkyu9M6nfPfxf2okpXwtyHKy
w4Th+7BDBVXzmZpD/eG9habO8pyWBetm4mr1UWi5suN1PXDsZZSMZWSLiQpC
Dnho5HsrV4XRRv8HH3gg6YbL+ivJq7y+LiWBYYUl0XNIjYN5+Up9PSdM3j0G
zXAZC1LTxeUBH440OfAB6Co4Lx4famLC6uLGVIu8VXVMP2I35zZC6gjV0bM3
/lH+Zat2jeJ2LbTFybiabpAk7slj4j+xCqPPbZH41nwuv0lvZzotLBZkpM6D
hDzJ06a8lgc/47r4tHDmS1plKygDFDwScyA0MXMCZMUQm1DKhe7YzQPjs0rW
8FWZ+JhKcUVM+HfZ/EujFH9jz6MXyHou+OjqxMLZ57r/qEIMGDJUvCScPCbu
Qy0jVhDw5PGyNaEv08ZL6bQVM0Pv+rlolQoolOsHUP2vQ0sNJLSwEzrlBAr5
DpxqAaFLUDYN0WX4Xy4E8hWDe/GndiHcXhX1a3sTaVxvJ8b8uetiLE9eQUYj
7/EgJcpPs2iyUqAVi0Fo98j3a8dQqfyO+/3BSBqoBwzSZGOul513oHeEFCRp
bewUdAs+iuym9gf4ztVey43ETR840/94cSJikzhfs6rhMPlCgOcgRSRPYLyY
g+FJzLCRxYi792gVRUxNbuOXUiUXdG6MIT56WLZ/VfZZkeoZxlDMarifLkzT
vIUJQdKNe8LFKmkga8sUuTv4+P3QEioLc5jTK9XAiCNI/UB/atuV1wxrsBPs
vkvnP3KvwTcdP0C4yn5N1go7lUi0DpGPQ5XBja21PITNwY88YwDdShrIIQUm
uKo6bpE0FxsiPvyiJ6ORzTqO+GXTghSMagO4exbhzf3dNPPc/k1RxzD2kGZ2
I2I5x6FdZF/gM7TtbFBJaPktsch91ItuWvQsvKGXZjneu4mVOg0T6lAONikL
ohKnnYB1XWX+QFEJEusjcnl4hpUAbdpHUFeV4ElmCZrCd/kyXAzDxerJfZjr
OpxJkQ7/8hdOmTfKO/Dk+6yI9oH8ds9dzQaoXAkbIVBX3GWMjLVMXAWuV60b
a9URQhXHznV8JEK9HYJSCNY4k7zp3ZP3R7HuPPVypmkfhfJYHbtITIc9TT4P
VyFGGoj36fT6tULNdlk4qFBHv4xRBU1rXBXSUph9zVNMYjQF0gYV6cmVOk/h
Ttg3e98Q4QwnCojoTiTpEAxJtIt8zR1nnMGeYuPylXTyngfW5TtwQ88lwQXG
cjrc+ADQ9OiTe7QICuPwqYu3AotLCY9w1DbFhHUL/DBkdilVwuLNCdtjPIPp
uyTfJMBWRsGF/wnElZzMzAV3ACH5FnPGy8nMW4gXtR7qCHMH+xI+bKr7S4qZ
X1IngTugUt0q8Ni1TkDOK385UUw2/Vt37G8+mG17vHTXldv9ityg7724itxx
MpmGtRs8KUV4SByM+r6iJq17AFekgWcSDIhp/29JhWMST7HoKl51ID7/+uAy
bgrSvnLOOLtYW35Qzqcakrw/gkqcSnXSmIOPpR2nUeKrMFKZDvjtec2V99t0
t03yRora0H/F2XZxAp49uKn7e+pqEsnloqX4yqEVo8LSO4vy7hz1wxLTm6iD
b8NCtRAtfrwZJWHCm3ENID4zTC/88ErFHCys38DdYwdO0ywmYqA2W1q3bVwv
DU+l8CjEpzPvKe91Ewi/SpHpkbaOCo3UG7PnbzfXoMnEp8k3fSP1Y90dxHtm
xCTHp4WYKVn7EG6nmqvD+1bHjJi77C0y3JObV4p/BRC/VOCeDnxaIIZSW3TA
j6tsj7a4cdGxWdy1dniXLD0i4f0AcrPcLw9wnODuziEXozVNijZTvmLq2Eox
UQKFmtKyLv3KAnvJLhZxUUs1sn0gqJ/LMwP21hn5hyxNG5nD/KMuPjSV4W8I
673ex3IoqL0rpr4n0v+SqDbasbUjilLsxZX/85kSHfIUqv2p0FLjijdmVtnT
82ungLlmTlmMI4GsAinztYiIT1OCLaiCqv/P54cXnMCbLSkL/U2qZa3YbzEC
c+sxjMnepxj0F9BetLKuAkgpZXz2sCO+3PZihqS/nP0FhYPecMJaS7434geV
gFjwv8fOT70eF8O+ag9CkcBBZtAkpSZmLzqX1UF9xyENMUS2A9JWtlV7Grfn
+miD6R4CHp8vdN1oeS25CbEWuhWsdQxxzCqR5aeOFA36F3/AjF7z7ftbHSGz
9FGp1WQPjJkfniZOlu4sylbEOhhdnVjZjdpErvlBdQg9q2Hh7oRLlcCtSlWW
k8g1JkOBZlz++/L2dSk2p87aap6aXP68Ijdq2trFz7RPtDcv9D2m4QxYybRU
jxCaqF1GB8QwJtsAnxKDVgZFqngNbcPWwOvpCn3wFbSwBOZyRJ4wKo9BcsYz
ARX1PIBX+KE8lbTrRgnT4tNhbqRo92vouECHJ3J/Qx4tEltkrx9ItVrMbUCx
wOXO4VeqeWQn+61coa25gV8dUc2cRcQzkXrKLDTHxJFLAIRRLjF+Y5R4JnUT
J8q7k1AEh4elYpkVNoDuDz3/G/wKQw2PA9dAH9prlwAy0R+L1ESURg3ffObc
dA1dnVwjwGuVmMdu3TDDNxiZc6hvTSLFXlMXbBefQdR/2kbVasAYJZMkaxc1
8HpMV/TDlYRNG81Ig263l46bnfc1S1iTYO68ghq0urt1yzoFpf8b2WjNZ+qW
m4q6PWNbVrX08DIBvuL7RFV1yLKskfg7u+lWrk4AXAoCNXHP++kM+DdQ8d4o
7kcUlnMecQ7SMmfuVCf1Bzrz25ltHsjhrEVDxgDaoxTxRNWZzGKq3l+mAgTG
FmPPXzqwJQwXPXxj7JfwQTgaeIFVJ8i/Fz2pbsjF3oHSW2pDT/9D/xyojWfL
9j1Jp/eEvMvwgWj3Ce1yBwEfcxKo8SieaHlyY12qTL8sin0ZdzpLyRpcfC4q
Ntkcqi+xINd3kjm40X46Ty54Pzxl6XZd7cQOLvM6icnYJXsDqKePB9Rsuxsh
UcOK/Dn0YlT0O9VksEi4Qf1m4EbaM1IP8bLbGHCPvvjkjVDIQOx/Y69Fut0L
Sh8mg8xtHgDgk6VDGCcu0z8YuMLvtWgxbv4BsOkbsBCa2FAuBavWE58QKKWe
EMmx5aSp75v9AyGYOBO3lmvYErUEE2Xxs8X95Zm7j7h3qR2sO5PDYAFYCaPn
9kQDP/51oAmsiu2VQGLl2E+tH68o//AjDE9U0q1dOjRXIAR6O76FuHUTSkK6
I0qxUpQ0drlJzO+W0Uy0GaCcVoee0fLEG61Q1eURiecagl8e5tfGfJJyFLQD
8KthX5guKHrTP/trdVeWfxgVg7v1U6Aw14WyGR2ENvf03Wdrzr5yNBfTJ02N
caE5zTdufMnx9PLAWrozB56bmm/jibqFyYE7s5Y7wVRLy2S4W71oNR0R4pnk
AdZTqYnYiTDSSrKKx19++8w/sr8MWZoJr+I0gJGfh5eQdq/v4QBmpxRzb3Ql
R3y9+BC8UdsjQKlajqW168GkvGEbVQqnziA6f1Em8FHxkoIj5kzUPpfQgbZ1
m1eUBNWhfuDtwjzdnemvrxoQdopKcYjJe82F9/1a/yoLE8w7FVvknTi/ZAk1
lt0Y52DE74cilCG4u2iSvWbqDLx0jyTaW3IqVvLTHrO3Eoh9/mZCokF0Y8zW
sj56bAEyTNfczZ7AP73qoSNyEf3bm0btLaucmra0XZkJrc0dKuDZnofchyjb
ufvJQxLL0ug7edlByUwaJv5cn+Hcy68e6FjGZHvyclMeSdDVr5emApVrv6am
r7fCneASNRwa076TWT4gj++Vc3wk74MXH2igO7fGFY9lKHfWuK9crtq3idbn
GVwoxSMoGhAmhaS/n5qP2L9jVkjKSRdxPOVXWTaEs7hurBHszXzrWWbvuycs
x/yafiRBKGhCgfng1nno65etXxhQUMqvukvFrMc5V6xYnH2C1TvONSGQL8nJ
dWNvlBdFb8rXuMTij0r+u9zJ5aNy1fzACPLRnSgEu1yPgmWkPX96Nne/zv5g
gR9mBA0siXT8iFij7S0DG8ACSrFZbwQquO/yuK0QQ95SRJk+y3cwJ+MZHR+V
oojA9WzQVEuaL9KAQuds6n8kUE9yAhAEJjqk4MvvN6bfnEMMfatALzAb1ZEx
HZogU3aKHoa1Yzpq146o/NVeN2Klh5tPVTsm7khbDZ26lOVZRr17BibhDHno
JBLZbNkorMbtJAFks0QsLdk76LPycBVAudRTT56/hrGuZrrsamBmABEJSyIA
c8NHzUZ3+wkYoZBxEFNq4MaTibIG1MDT19XDA3+jsVZ3QDhUBk3u3h9wXPpR
e7NhcOjtQ0iQ63vEmRBbcDX2U/38jk+vqUEHoN7OTSeoOVAtfaoV2vooxKHv
jBbSn6vQz8rQPWxdrdMA4HXPcNIwAr2Cn55rGFe5PPgTDhnD5gcp2o8MOZjW
+QKjVwlLFQKBJKEJvDfsS2w31gsA4P613Y6DIcI/8N7GgvwIV1sHiWzJ0gfh
skFP1JvBhP3tsKiB61z4itCPruvopjj7NCwzYmcLPG3u0iejxcUVgrNQ1WIa
xG01MOVzTHQeeh3dGla7QtqgaHRLjtZAxamlhMLy5OyEQlrfxjU8L/+AQstO
gY59Tmrl2UkHXsTxTgt6e6qO82Sq92HL6/PU7A82UduBE80KV+dhLoLcLyb/
6+hSzIyuUdiFoCZVTKjwNzoG02lIIBdVRsbD5BpCGWSX74uCocqUev2aU+N7
jLGtAFw03IskknNf8EynWRqe8z8vsu5ad32N29Zw0ddG2+h+7M6ASBzOXxtq
m6MGI8w2pNnPzQ/NEUeUagPozisakdAgBO4fRLEs/i4RiWCNtPAQ2Kw0R3VY
6j5FjgTSeBA1CZLYOtm3nzyGOLeIXBVapwJD3N8AI1bowliDGoWqt1vjo1va
Z00djYy2srf9xw+rgg5+RmWiFyHE+/a2wsrSfYRSRJS/erMHTd0eVUPajtAp
l8gj/5yOKkMC0Qj+tkFcaxuH+Pak23v+PhpjtKizv7OhLOXHuOvIgpQt8x4V
bGS9kGFzx0IVpso0G23cbNwYwh1e5Vo09UUsLI/rOb0ss6jjusAOY0DiE5b6
VsTJTEvoc20R/61UE+9eAQKu3v/NiY0+UuweB1K9yl1huVLdlr+1O5UMWUty
jWxMH7Pp0eu6Bimer74LI/0072f/vOD2tlzIt/Uj+gmKkME8CsvT4dxEzTRX
rOIEn0FJmZxfYLbRe/uCCGOhVKAGRkM//Dv2wYcVABVqsTbtPBk1noTrLoDE
AYb20EgjcXXoZBFOqdupacHqIAmF89WAxFYqUp99cGojdU+ArN66zcSDmvEj
ZeQ5qX1JRvB7xAVT7nFERM1Bx0b1MsPmfqnqujcadBDOdx0BDQQZ4u5TZ6nL
x/sTfz3Ud6gHgQ4pD2muWMZVdLweAHXGtytUAZBHBcN4PK9v5D3U8WYM226j
HnzIdydIImK0OXOiYE6tAHeXhe1E5I5fRJJNFwHSDZEsBK9St/CD8yEjAy57
7T4/j/4TUlW9JIdBkBauNoKMME+4CDW6wCqvxbvE3meUTChlvDNM+CJcbbAO
+LBiU3KApyflwYwlGdd1MmiZuuHKrBuaxWfK8EZ3EiqMD8owvW5T/JlxGIaI
ZCc7JbrCFfAJTSBDpwJodAEJuoqG3FEvSJjttRpiqmPIp1rrNT2nwZ8TZNU5
wfylxBQwwPZfVNyD1s6VjLYQGf9YFWcImIYP9CQ28eB66qF7ln5hRb3qwf4/
rAqffgcWFcifsinA8l+zO3q/oRjKyPU9den06MMXkiVHvVoAO9Yrfr1p2W9P
w8rnpfqTDzNdElf9ucHvWaH5/tdP7AGefHa8d27qBFJpLbJ/WEArYWVoK8w1
lbKkFkxxsBMq295uGwEYhhXsHFuir/vu/9DzUTicfVghgRlzbb3NJhMg1qL5
R5+clqeWHV3Rt5lqTAvi1EZJPY9ZrzkDSEvoLuwRD1PiMCQxQSxgUPwQzQOh
Kav2L+2gLK9aROxBVauC+/szTyeMUsiSBo241iVuF+iuKey1QrM/yXoH5inF
wHWOUayqQnc5+6OK3NY6QgwzKZecgcBZoLy8DD9d3m+Rcn67ZYSFcRi/sqj+
ltlIhovriJ/uy8g4o/cq7J0zrfc/Cheg0/CTUZmHIoCjIphcaV+3mo0TZQlX
ACI2TUO2tB/dA48ckQ8lmLCnr21xwmKjwOmq9daperPdZHtycmRTt65ZnEil
5dMnOazKzNOSPpBxXOAaYPV284soiwchRAbJ+Dri2zcFuxS453Vwu5cXa6UH
JUbpJCCfKwzmeyJeCRHyCJ91J3XzpURHAROYrcSEJog9AhHj6zbfHT6veMLD
7r1HgknfAls89+Xr4hadgHAMbcKjo95UWIZYOu+cgfSodfADJYpX6Jd/qXAa
Dt0J1fBOtLnudFGodU3a1XzsZzDwEkYzgLmKA0CgCBt2qrQD492VoMTGlv0i
NQKT9gLD0h/3kYP1MJfDRjoh/8aF8+xUOYaTmkp5pGP2WN69IQfezwv3HOnp
O72aO/EOBIYPs8wP9V9Fglkpr4YF4GpiT4EQkzs9H0Q89p1gzuvqUW0+yUM1
PB85svPew4IPDPcVx5XPbf8DCdX98qRmd2kllA56txNReTxKDPC1RayLg2Nl
UYkHfpr0IqSjjq6R9f4LLcZiXJB8YVE9Cu3JsY5rsywQho1/jq7sjAll+9Jf
nULn4sbNdtVOaPCEWmVF5CkJypOQgxWxrNeBpXnngv6RR0Ys0jwmxUJjNIuG
X2zUNxKXibA6YKiZyzCTY4aar0v0QI4hT5Lr3vAxLrDlJsQs/hcuTgQAabeW
umDF6YdwZlXVzkfh3pqXmO0rsiDxGrTauee27eTGHvO6CYIslS3tFo+jN0Vu
k5W6ANEL4Xw6DkWUm60QrymsshpQcxbyXLoX1gXpLsAnWZ/ZBrMM0EzCc8fT
xF+2Y/E3VYZsZzhpNwxaGtsdqdRxCQVuSLzdRbST1bi6n49L4hOjziZDz3lD
7Xilvbw91h4dqg5tr8BGhm48lRN18Avpabj07ysH6p5kLbg6SsFtaPng/UH3
drlKQLbsIsTrFHFcoGFvssytTIkOQFIrqGGlu4bJYlHBcT15Eyfdkz/ZdAb0
VLxLIbS3np2n1KHy8OiHOLbaJs3GaooKg0feFWjLMlkqj9hWiegmCW0N3nfX
mpq4kRIM6dGpWafwxA9zgeGIMH4pqPDNn2RlIf5nAo2y7rxbp9b20by6hJsj
nDTPGoPKXHmy7GW0hCXcSRA2269PvfiuJHDQ9P/JxPZEaBfRBy7CtyGcH62q
ZD5YQCyD1n9s+XRmAeR/OB4CapSXXyvrn9PloXo5v2afw4PbBl7dryOjP6U8
8/S/A2bIeXdYasCkX/oMDxyHSfru2xAcPtg5IEMd3jSqaawTs9WtlvTGhFIV
SzPw9mY8LQ+e8q7vvMNy64cNhfrfEfEAzPSGvYnehtlg25MR9mYz7vIrbcw3
EUE6uJmhDOxCenYXigfwlS/q8lAkeQZKMQqIhRXZHzkpP9LxcoE+D0rH/SFG
OVr9+jalpddZD0oOrnZszXJbr7VSd2YRWRXNXmGHLpToXvLmbemR/dv/wFtm
6FqrEaMn9OlBVo1Zgvo9Ak3CxXMGW+4tIy8qahXl4ZyBYGpjhlctIRJ/HcBo
w4XYLwnbgdiTnyBW4jBvJFI7uZ9kByxj3KMUZI88LLD5HTVMw5H4RVNcp28F
pRAkPSafBJCTlhBdoAWCrKarQLDiXwfVWj/7aGIHXHNiF3gLZOC9O3oAi2A0
lrCQObbHvDilGUkC/nkWx61T014I3OH7f4E9oZERF8YPb+T7K1bG4GIaSdzd
gluoVwg6XvJFsX9a4ssBT7lTuXCC+RBkQG6M3r+zC/wlHXsChyKXnW1DQgc+
Z/PRe6m37gPQybphDxXbZ9EkbQyL6btPAGi/P+ErQRnE4CEDVIksovaA/tgU
Md+bnhr+TJKj/wGC/wQYAIJ16facYu1IyoUN7tDP2GdBLD4DWyT/WxBbwzXs
Wjvk6wxkKz9FVfoZCWqXczXdUvRa6/Ir8g3VG8Ot7l/ur8dfhrmeYw7VeYXX
KyPW8snZo4dZ5eU3Zm4/ZJsyLWbNg9IE0xLJEMwFpqUtCg/wfNrwNIBZhEJv
vl/9pLvuF+xnrCeg/wNvZj/lffm1GgVviOQzlyEvHwiEPa/iYJEXex9MtJiy
lfqnh3fhYSnUcjJj6yY6VoqaPIio5fu4YMTqnG7Gi5x2LibXkPlVXByI13uu
Q5MK0CtIGIVZKpIc4mj1RVovANL+/uiHq8U2d1L+lsWfSXr82qyf4R6wJrQ0
k0BM7pwzoI+NYnyU8fNN7bqVKOBdEPUGRvjG0gsOgorlp/RGxvyAr7/4Z4kH
ImYrpEnnc0hGqhthkOrJ0bz7kigUo3gx9TbV4YCabmEn+DMmdhbCFwOGRcVJ
2Y7DJMypf4NP1NGQkRWrw1rN1HwhWQlrgMK8hOfPXW+Hmr2SbPvxHKFhxp+N
sbAMApD8FTmPJwixGzNmXJ6J91UhKyBMEk2vmcsq4/KsS6sM+jiDumLz45Na
0ShUe7LWsp1FU5ZzofajYsiyB2mAxvjBBG+0fC5HHN1ra6G8wHf11Em3ix8D
G7HRrTaAGMcqy8GNY+vP9USantvjUjLyx13TjvZ4WAOggdBf1RpzZIlujeKg
nSFQVPZBD/ocI9CL8nJzc90uBUA1Z1+O/xLLIc/srn1n/lgTU4uAFJXwm/bE
UO1/YggrMlGZ2gF0GUfzwf53XJLtmGAppZ26BJ9XAg2Oh+Xw9X1Wf7arD9wR
jeQc/RLT0xBlnqMjdF4JVjj7g0nx7QXWcFCzhF1dh76tWfn+/270gIGPrXN3
egCz27nXJEY3yBcVSK1xXupB0Kw3J4K/YKSRZsUCih4fimrHBkTNMVjm+aKp
W3LYbAnoXzwOlQG3AdvUkGpPXo52P/pGZ3Q+FxZYbxHIVLFX5qOSkKRFMW8l
AJpN1hTaY+gKaNMSor0H6drsi48T0EwZlATbLTn8frbWo6Knf91TsDeI9OEA
c3YTFxobwl4UDpBulY/dMJldMT/Etm4mmyUKeOjOvMVPA3wPymssyqahfwiT
Tb7gsxkRMu2adfyfeY8tiOV5/6vLMYz4DaRbuYTpokxnNTfXx/UOON2eGeSf
5nop2YVunw6+FoNklIckg72ocg6eJMLoPNkVjAl/BZLAkHYGzHC2Dg9CCSBS
x1DhpaqzqhV7AmQy8F/n7UUvVzpwp/ohElACnRVsudUMRLVG1suNreacKdQh
fEKJzgeqZXf64i7EX0mhlN25lwaXvNlSHzb+bXyXqvaEmMe+4vfDUn1lGkHX
0Hzj/DK4hdaCxnr7Ke7mHzM8Nvfqs4AgTdcXUVD4zYVHFi1DA05hLJhqrwqy
hxMB37mNUAD7z/IoUHrGK+LKftuxNIlqjOlmeQbqIPeBvAWQIxV8Z6T37HpX
dB2uEe3QUQIAx+YsJGVIXX881lqm/LNkK3rdn2uBBLU2Ir3C3Knndb+ZekTl
yBlIc8pFQFHnSuE+EeMeqi8xA0EdZkVs5MUB1nBAvF6Nt9xdKGvWtNwhm7yB
igkisjeAX62qoyQ8Knis7vAzIhNYsGWdPGiRw/dQGkhJAXt8Utq3ajDUQMTY
7OgOwMQzh0/Ab2xy+Elri5UVqR79rUeB7q4II+2ig9kkpAZ8W8UoGk75slCB
aE6Lu6r3qznALQ8lXd6gl4DwVAogrx4mBWoY3jk/0AKYRc5wr158TDaN8LsL
2IfA5jZe2zHZbs4VY7zohoAoONjT8J/QUeNADlExJzM1n6SgmzIoAccP5A38
tuGl/iTlNUj2EoQR3R0qBpcz+LE5iwe9wi5maEXdgWIB5RQlnBdxpXmnpAb4
2HGdntrFG9zBQa3ILrnTZpK4ej0j44GBEWGBUy4h7SHzX3FtSmxDEA8Y9A+h
rdw8j00wY2gpP/eqbjv5NuigLbTDG0lKxRUB1HlgzI/M3m8g1YnmU7RE1OCL
0zVku1Ch8xL+j1GZXAWlW91tBj1k9e1T3as0SKOwHqUGOhPRcm6Y5II1+Y3k
hbU9yKyONUa5F3UQsUAKzE+GsGW2AfZ8/XiQN/76w5MIfIdCxOSY7kkwUZLU
IJ/A812Y4404cqTsPs8rsNOitQLWdWmV4w1dCgA71Q37ISLO5vZQBfxh6q1C
+FblvnSm8lV+rvY0bvrN641+rzKQQbSoUdNc9cHUKhgHocYl2Q029s5UnS5B
ckL97hI/FPlDwwAAa4in/dG65pENztcX3Fl6yZ8QzlRIKzp+8HFXEdlSJsvr
5t0MJSik6gA4v6oFIqDMuaqSU/qa48XOJLxC7Bk6rzyaE2jf523pVullQsbH
DxY9MY9+8kQuagdI6ZxLyQ95uRTESBsERb5qb62Sz5LNdwXY7CGynaghIOrE
olNC5szdXHZo0jcveIHPgA3ZA98Mt6P80coicsdEHid8y0xc8CQDM2mevrlJ
pK0adXGyMGJ5Ji5L3d/CoJnUvs3tDivlT5tmd4ErN1tJ0eFetheUuz7GA8UQ
bu3luzgjS3mHGFOSmzw/wHtcmLGtNkk4MceIENc2CoFyx/IWQs88puPkvsV3
MkTPwIDGlZsSBNm/Co8LnPFO15+BLSx20E3AWbW/mOCvlIUN3PLsbsxZS7c1
1a6CqbsRNXg4Hw6BFgMRiHPDUne+OrmLhnBvxpZb4zJPHOa/94kCIE6sZIOV
iWhiKIgo+a/O3rPGvwn93+HYIq/NhPmE3dQ3jBYVyQdDuRg+3/7gfgU1N2WE
rAGYguL15Lb0/fQC4dtXZHwrj8jcHsrPDI+cDdmSXGU3ZNOD6SFNShBaUjS/
AwSoMQvb46RdUcJKvq7H4MJg66xuNd5pij3elCZ/XOM7R4CbtRSaKerkUfLp
mY9IpM+2IK7pj/YUd3fE8l0YYQVNLpMc2vYVyTqNrtSivLlWI9CqoWZxSIxQ
ujnTdsEdUzivMtbDT5BymCSTSHEyEZSHn/TH7LoH8D/uNtonH5d/C5xPZYVZ
01jU20KukvR9C8xcMFv3bXKis7AzW1aluIK4C/h3A/Il7mveqT2YrMFjT6On
RwyQ/CgZEhBKfPVck+O93yvwEBAL4JKV0Y9XqB9ExxaB9IgTll/tooTLmjBm
wf4SdYyzmKbJgXuVIfzyaUzGb+I6DMeYelN3t/9qPV6DObo/THN6jZ8zp/mg
Z+z0xRKTZjkx0nqU0key+eme3V835jDw2cOLpSmIxtcCiM2IaRrPs6Hs4ISH
Z/+Ytc1JThsrI0IQJHg3MoTJcfC/f1ODeSiiOB4OeaLppAL+VRFZKYLw7tWj
jDf+fUm9Io0SYOUVuebP4hRf7IpLjQxWQvxbQ82jH86OJYECR2zkqJqCeWgp
0raBYrrZYBjNF8l4/HssauPb5SNCdmrDlrnbwTK2vR+ioZNwIwYgxB8DAwbQ
rJWQoIoc2hFyDGJ9ZZUt3e8YRELqfeLsWYrsJDFcnbyWMVJmxzPl2FO/0dDN
xcwtFVWsHxBGrLl+/5PXCh5Oe2TTp5wiO3eNChZKF2qm4zHkdjcXPBTWfuWJ
puIAaP53sxVnpWXW7LSjO97mdQ1tgwKmZCKRQtMufVPm3tBLyK++BQl1AimW
2hMjiP7NMzonoE/K9a/jVk8X1niudWL/kYrmOD8O8HoajbP821FClYxeFo5v
mO8ywtb8Xy6TkVAP3g/tWG6zIhORD8NhkhPho8sKZ0ffRMjUjfAxiT+xaVbv
M0hJZcTfQy7hRDzaThK2fQcmikVVNh2RgAN0MvJ9cT69/1kLRcDytI9saQIl
A4J09OlXlrontBST9/hW+hqOwjBa+mAtbmOIQf0ojCs6DFrmAXD++6Mia9+K
Iqt1C/S6rzjSuEcL16se8h0Fj55PEkI0Dr8Zup2DTQS0ZPvKsXvS5dRH6zFt
eoyS4TEqS0+YA571ACFSpzBkKxPn4n5Wnj0OLjT50+DUfiA6lh2l9LqMV5oz
Ac5EZAGJw3uR/OTv8DkLo8IFAhRd7CPvGrCmMbhV9fGlMqm+b4JLEKmonT6P
oU2eDzCm3T3ovoN22x2u/4WBAJQZhHlXG/0Bs273FZUvgHT/LTXSKp52vnJ5
v/9RYjCJxOAriYFkT53ynXj8yr8+h0FPzOnSi8h9qZMLVtoF4K/0RaYATC+e
D0rT4U+NLuZ9rG3m34RoKuoYUOgrBFjepNHNBnOCNWbOFE+NP8JDB/uPy4q+
6Wbxny6XvTZMLTNq5NjKLCY1UnGYtsK4vUGHaToO+27a30dsgu7eF/ojwo19
w5g24V8pDu41kBOqvgz+JZot0aVgJEEi4/6C9KPv6tfRbaPZzD9oYV4udxKY
HoAcG+rRZrdr84S5dWrUYTYTDHHiHmd9eJ48MsgVe1gQwCrHMXr6oR5VoaDi
aKOeBtACxHJMxNUwf9qxBXdlGbR4tGtx3tzOtpjPlxhxWGLMkAayspO2BkvD
XuPUFdBHOlBt7EM/CruWbjKusF8YMQjmsVlB3iSWEwszZow5V3DJS9CK86ya
PDXikhKOLy4ODTqsv0h4iwRri9V99TjTw6q6NtakMhnRlOP5ZQR8CdkA6Dt5
nULzQb1jTvcyltB+l9Bszo7NtAUu3tRZw8ToU131QyGDmyD73/9DJnhpIaBs
LOeBiaI50XRy0Um9Qi0ywoPX16CWJlnqlbeEjmxEuMmlxcNbSi71VxZIL97s
mBk0j4RT9E7aE5yrdUNUep8u0KqPDMeAa+6SaLOfaJKkgmNcdEp1j+u7OJOD
27e/63eFI7H8lH2QDJVTezyvtkbYu5i204sAoD0y2P8+sszXGHV/iFv6Ux/h
VyR36JS4HVqg2mqT1BwFLzx/dIXVclq4cZmUzirVLVWp3Ps+0yVEZ/Q67bph
+tBAToB5ZNJfrDGseD7FTotRgyscDiWAOh4GHeF6VdZNnWbjMVo1uhARHASS
wo9VZa70V14hl8Ff6rsFag+VH9SdSg+9206ercWYKsfOzayPu2rzqZmlm0EE
aKwnyw/YJG/eU1N4AJV1Ar+Pyg+3UDgv1lVrAOJQtO91AW5Yzguc+KG+1sRk
3LWCOC5E0eNi7Rpxs70V80EdYiz6+t5HIxF8+nmn10btc5oCnTr6SNFyNoiV
WqZMF1wlrk57Xop0Bed+S+0raK25XSrbFgw9/y8pt8Uu2GehS6iWezTcvMnZ
xTG4yaiAQSVi8BaHn7/thBeY1kwvdzUDR8gIlpw6J8+5sEffkgv3VeP0q/sG
A7QTGXkQOR1w+Y/3KlCmyv5Mln2dSchLoTNO5+U+lgg6Inv+w8ux4MbhKstV
SOAKVgrkqT0LJlRwP31NeFOEv9TDU9K1mGxZd1SGViTk8+V0DFbXfSzoVpRo
Ud19y7UnkvpMu/T3ugRbzFbHTvR2zvMnbQvpANou/JR1XixSfANpnvLI1BC9
hCUmrXcGTwuUuqfYgJkZJ9pj0z3hL9vEbvw2/3edFu+F3FRFqXoRKBD4vHTH
lkgFfjGWNrvVDNGlylAjKqdMdRdKo/ja1mVCPXjDiEMcYkdUzwpkyk0IgcpL
yR2NkQYu7RIAUsJR1K8HondmxXdDadkNYhc1J3+igIb2ROh+Bc06Haj5SfHC
/egYNqWIUZmzCfZ5kKJ1E4lxjQ9PjAoYJSgLEgAu+ySfnuhynDLKrEwh64Kq
v1X7VvpMjD2u/KRP8lL4gZSidN3I7sA+FM/rdgYf+OB3QlCaXgOIASUvl/Gv
eEDISs1FMk1QeaQXbtEMyeB0KTVR6218hRRCMO9ELLMgGzTsOKvdpeSkDx+k
xM38pT2i/ch7Kzp50kk+k5B/dk5IrueKUbx4XqeDakavUQ52r8KLK2F8Gr7C
+EZzsjniRSW30vMYxqqRtVWfAJwI6gqY6Shd99POy3aIzKnErlcYN4Le36lx
BkjBS5mo46YHH/cwHayWVfSSAxX1BV9UBQlxj2MkPGl6ZGzeany0PnkIZMA7
fF5qw/BpbxoOA1wt5NQGL4h1tcX4yezKMlnz+jpFD/xgDKGXz9dPp4+FIKa8
M/5K1v0Wr/Zc/1/69brnUyLiSwPTwrMmtio/50Y6vc6fQcp2gTug/SgpPV3L
KUSQzKfONCyO/ts4RCRkphmfVeL/QwGPN0nYh3IFyoXFlp7VHrkzLcRX4dpW
GdLDi7ssATPsHsXtzOXxtVOQXEVaMyDqS6zcYxB+6ua8vkcGe3Y5b1tTBBLu
9eikbb4wTDMuZHwprogzAG608tsNBqVNTMQTG24+UFOcxbNDMe/l3uYHI/j8
cqNyk/4bW0Epe6QCoMtyfYHKSNtolgySE3V3bvtxXG/Xum79qRZGYc58K0RT
qDIa62cuhx3f8EQ77NuhWd5OvhgKHeduZ+qTs8im+pFbhP7Rky4IyfMdn1Bm
zEtWMsuRIZMV81bcJpADiwVr4YywKJ8jJHnE9s0F7m0XE51cXar5Ukr7yVuI
Wa2rjjOucW5fgzBFdpyAc+EXrim6Kd22ZuKXZrRTw7TiDvUsB8hxZzHYbK53
T1QWGyF86O4Tf/M3ykmScOh2ZE+sVIMGRGSX3gdjCcHZAEURF1L2b0sbo9Zs
Capfkm9ZY091vSRHO0gBJMIua5SwVDRJ3nOhxJYomWqO1YbpyPS521hqfuDq
IsOOXP6X9xwURWLqzCJi7yutCC3aj/WkYUz722Y6s5FSxL1SLxKbb+VDBSO4
YXyiIPizHPqmvM+bVjYQYVG5MSuicyU+DzDe1TMoKpoJfSlOy1T7TkVjjkPY
fhnc08Z9a7WxEEYFla6PRQamcLg1/E93P38s/5I/pQdtpu+H0Xk8Y6Nbgl2v
KD2QwH3hxcIHs0u4mzyyzQRs2UT+HSVw31hM1UbahHR2fu/1T19xDrylFb0n
jk1MCmP1w5nfAR2QGLxgwLO0MCT2j974LArI67fxdjD8bOAOzjw6CkcCFwu/
I6rMgIu9Q/KMg+rfWyLRx+MqQ8aupdgwD6ZXCot5OPN/bn+MO826hvNwX3NE
n1IJWP+C1UzrSTZEghAJ7hEwK9Ufn59cQRbKwt9EP9Ii3JkSdEdNw+o2WK4E
gRn+0OzduwLzHrzD+fnMk1yVB9xb/xytL+8AIz3vwVU2hUDedvuAJ6xaounN
GEHpK98e/zyFFCbs3wg1LLzBR69fXuXLPNnY0lzmJhTVLbwqANynZye3bWKy
GSUPeNAwKVg7ei64kkCUjeELxW8AGVd2EsgBZ9/GbXjFwvaPLRPh+weyky6x
ggQ7grK8EVsx+vtd1J/CLx3kOQmST/QR6SnpNB/5q9x8khZFRqTJMr/iazPN
jUsKdVoQww4PwR3aExJHg9r+9Kwbrt821FIie2WKkclqVFUtIO70j5WdmWLS
ejQ2bfsDDsbX+lwcKMnxlEU/Igd4LAmFsj7sFEWHtdREIY+dhkVuSp2oEjaV
TeRD082jaqVCxnpmv4Z6ImPObrvaku4mJTeQzvRjNlPP1/1g+K6xIvnbtIBq
2naZhfcgMLjFqQvA26JojSaxAKCgQGXVXacrALLI8RQuteHqhfRjlGT1oAGe
EwuhTjW/fZ8IvGfGz/R8BRZ3rropZo8OAAwNwS5pcMYJT8wQTHOgdj7MI0Qx
7Vhzl9+fOS609ZyNe4gNLRdUj7wyrdSwL7UP3M7hDNLHOzRkgHrn5yZmnWPd
8dvmI1lezIgR/59Ns/nJEy9ASuaPUofr5xuG2sueP5rkEmIrxaj+ZWeR515u
drZgn0+N1lgvyBNk9I6G4+pqEyXkTizPwUCvxLUVzcmej8MgzLUpGcdV0+7z
wLNlr8WsO5AJ96hGeujUUIflRSlFI0LdpFAmwwP69GDJTG0JVYx+6q0KzQNz
z0ryDVABvIH8+2moitx/0Pop4dDmh2NFNQPUUmedsFpdC69k5gEeGxQIitsh
53OF4b5dGRZMKn0+bx09FS1WLOVFYCLyoJz/hnJZAxWf27THhzlOOhBLquwa
hNRIvx4hkf2FYg36MoGxulEnNxfZvVM1XoiGY8JvAph+JKyFbHNqhUS4fwH1
vbyerzCuib3Tfjs8rUGcQv9wf/53mFSqgcqOgyVfNB+vl+rkK2P8xS7grfQ2
qARhyIVZmm8t2NaxT2Ou2+zwPF2CLxrkGV9GturHaQSb9/1wOECLWly8ej/Q
4gf2oY5n+xOh8tN6+M/ij5SLufUZ9RfMoE8ImRZ4rdprrKPGIWoOwrNcuIro
hnyuCmzD5r402+1SaRv4/vao+XDym8Xs6BGrnIKLgTE05LO6zL4xLHx9i8zg
RDubCuqoU45i61OJOGqkgBavYH5mdrzPosRhlF3tnvOM7CH7Qd8ZSZglks7P
kpEp/oE8l4YX/2j3+KwYUmslWH2g7NNyr3tYOlyGf2zILOEFtd4Grq1V0uEO
YlFkIuAPavQRaBLDglra5efY94da69y2NXRXjHFjnX1JHfwQSmc2D1kZLaQZ
UdZQqQL5gqtDZSaX/GFwOjL6dcEOQF7nVSp2qlnpqiFEl6E2r/uDevAp8oE3
8y6Uo5KyBqfNxrqVey1JVbj1pXCN0DLYcUcgTOPXxz2sZuvW44uhPvJNFJ5t
xdteHf8Ij7ZsfLQqeIDaLuu19kJhVwp4Q3yqXnf8Vyh0nhT8EB2LSNfCvrH6
ehKM450tTUinX3tJom6ute+NmKugVwcG6gBFYs5zijD1LXvO1UyPnjPS+Txj
ZmNE54cD3OKYAMAAp8Uk/zX4ehqyhGmBquFaxgmi4TDJoUeeJaGnjRPqh9jo
1J1riLtGow4iyUkcxIJadREwdfbIOt+DprdSoBf7hhcIetIQCCa88H9Q/dCJ
EJv1EWr2tJqUYPWGpBCnLhIncQ9Y9Xp2wdkc2qo3AU8ygqRqsBrTplBv+Gap
xPIkEZS8VbjdhnuPrCyVMdXKhlfZ6H4I2DLeeD5QDxUoMAqCMzM4sugu5Nof
Y0uIOnlzWajN3HXbCYOpiHBy+uEpgEJQUIaoS81L+wIzD4Mu5DxbtjwdacGH
LutspPfLypdstlpeSge/iJ4J/pLa7xtquqwUxWlLxhjWJYK0jrvZVSaqdXV/
Ni/QJUG+K10Pf5Rfdetvf185eLJnSm96wxvXFbC6EUmIYXXR2bpbFXuwUI+o
ieWLx5lXURyyBpXpreTCUX5JLmbfLNZNcgOfkqsBnMLAPlXIcXMqUhpnyI84
m2MKNDULuo5S4gGK/LkDH62/z7T0UXNtnw00fhE615y3opEETBcYEmlDdqkz
r07JsGITlVdJQB0TZ8AK2L0d3DMWdHNs0mGi7plq2zbWc4v35kOBN3QWon7H
kOhH4OBfgBDXwKPhZo31iqktwrRKS4TeH3N4pCU1BoQTK2fwSr4qPkkF0ZzM
Z0T+JZOeoU4w0wyI5aPrJpaRfITCDIFwk74xgM/uX8CZuFGUMXO8ws9E7tOE
sYHPh1MGjrjg+XN/ScUcv8Qaaylm/BfTZ8r863t5DFNMVgA7nvs30+TQ/zTY
AGQQ1eVORWI1WIxcM61gbFxLvMyNMTmMpVZaVuVZsLfNnTOubMVgpO6TgR0c
ILoCOkfNlCCOAlrF5ODuEZ2nusnNfyx7TvgTrpVMf8avPSG1lCn6L7IxG3f3
hUy2zmUrfLUD3i2POsAq/XyCKaGHYPt7s7QuZg14Vkif9/d37Xc08byXoqkx
f4BfJ/c02PJTFGJDj82sbKPfF5AT2QSbM2UFMC/bbrZJh6JDVWhzD8GfDRZS
MlEgi/REmO2bGLZX9I+w32E+wZXSrWNVvtJHr5zgsL+cfn7z07EOzJ3qDvpl
jA90Y/DSr9CiVYPWZM1KmAHnS2nRLzenHlm5zS1JedqmWq0MiQhC/dR4TZDS
K0P9ZZpQbwrzv3VSJoQ6MeUyoo/JZp1NQhHSGU4sFp+fb6injgafNz3TLJlW
TlLwfBq1uDB0EecuSn/NbPJg/LKxW578eOEgpRmonWxHG+Ng8Sy85kTiOD9r
zbIKzPTtRm3aZpRzox5H1UmhFCvC+lgNIYRzYXuG05uKwrB3tesjL5SU8iV7
8rfW5eupoFZH6+RCWDAJnLXcXlOUoDdAeIazK/aLC9LpvswAWPQ4sFE7GrLX
YTeZ1cFzRl9p5vm1pnChyZ7Px9F7AiSpIhgw37812Z0Pam5rKXNE1nU8n+c6
VquJEkChnYSgCGXKiRqLDL+JdiC/ggBJMlkhoAL/8XLEgvri7EPuHvBicW/X
xXhP+nRtLrFZnR9lZIKIrrENZMxv8YNXVtMzPb57lMqKL39jrf+RsTF2CQ7Y
VBs2Ckmt+gagiPHUmWnznExkzpCb+bEYiNENalWKbjA2OW9UnyZuBBfJJHt+
npW+ajjD/Jmxt7ezuvIbkUGw+7UgENS9rQbc6V61/3riEumW43Zil4FzDclb
NDMa/o/EK7UMIrG2CL4IC2NCw6pghZQ+6yW0SOnk780i8nQyrq/tdt3T55Sk
BFWA4e1n3t9Men2VNUrgvEkAiJ8NRQg1FGmxgcNhPBIpWbIl4FeEJSdtkpQn
PbYyrh+BPp4ZZLj4EdMlL+TaPakuY3Yb6McsoDCR7LE/0bBNhv8OrwhRSTTC
TFwhC8mlGHIvDDLucFQkSZX4K5ZyZeQXI3mdETHZQ5jFOzTgyQ2VK6xafsa1
f75JvrhoLNNEY8FBdt2n8/5XbLq8AtPtQkwQwhTOFdSojqhnhKNTStYB305/
aWMn6HXhwEQcxqfjaDHdGgFelqYlUOszOUQImX7jldbIOpIc1oKVCdiWNo02
3uDrDpjdRm56mh1MKkcVwL72Ip8LFIAfjt87MdsQo3wjiuoZw5cFkk6fGuyG
7mzpL8tjKY6MzKzJdW83DbJR+g6tFG/bBK4GTkr/SQxmY6XnXX+/BxQGU0BL
nQU+HkMbUI01FB8IjClZ55a9wqGM8k/Q++DiLY8YubcbVfSIv9LF8dt/PXgL
nbFM7jzwWY3YxhlPk/LYMKL1R+zpXgzDgu3X9b95AXSSEt0YTcB5HJZdHR9z
wL1ZgV+u40BNli5SWSpxerwoRTLheu/Uh24FjAjE5UO0dWvwa2SGwze02PQv
jdqjnDTkSeA+fZxKpEGjRFhOmNnm6cm8G5YNyhe/Xr+2vOPKcfkT8C+VW6UC
CaMcB7sesv5kEwNvRHdeSvJfUp8wHcMU//CY47HTEmE8mVE0989yaa0WtBUM
EUGpaF9Z4xcV1W6c7IrhjN8g+jaLB+GQCjoBgzBTiFhcvEEeKWFyQwnO5Xas
TD3uOm/Oc5Z6U4xREQw3ECiaaH82Iw8EpPUNlt/gbT0YaDXnaUHqs8LGC7om
mbn/A0bHV0X5lRY9ybuKbrydtM+PLp38Q/6ncIdbq38AMR/Ak+WvjXQaCsaK
J5h8zd49FE6UKyskn/Dfo6qw7rtm0oGW4fEHEFCy2UJhIMGBH8i0jQxO5qz1
5NQQ0HiLBTBIeHqSv+GTy5luV/749hytM2fth0FxwZRUXwRbKZUZctaKrqTo
tdH2p0zp8ONJzW/2ksq5G4noSBNCUmULHkc4D4BijQw/iQ7QM9gC8rXyKREO
GEYWeU2W9DjbDZbElTgW/0xTm9dhsEZwQS7VWEEnmmva9Ex5pLTNDHI7UBro
hUQJoF27WROj/PmSCi2rpRbENJ3pgMIonWdWGDHFnCZlov3HqUmP3+zxStdO
E2PgXQYerItpvFBcgDkO1ElBw+i46WUTpJ8e3nEjZRc265OcWGQHKlAGvkns
89s3SSZkcw6GuEa9Rai5zEty7LOmoXNuXD7pXLVu23k0Pll8P3+/Aqy/Dn66
wpLVTaX/jQndN0Jtl/figBgC9m9CGHGcJ5ZOBCTKY9yGknRWXh2MHZ2JhemY
1sq66jE61iQFmz5mrOBvw5pfy4HisxpVpg4nvq83qF8f/yuaiXAr2zKC7mTr
u7CqlTNkMTa6qPGUXqO6U8F06pBsivzyhO8aiPiHWvbUoO8mIYZaO2zokZ1w
3Hy9ErUcxBDE/FaGqAUyD/yr602hc0P6Pe9tdlRXSi1iTZBNo6oZUvejY5gD
T2wk/MegVkWDRXtxEEL1C/nFtaKNxMm4JoSzuckfytywC9/g/CqFbYDjNpW9
w5LK5Y9I+jFmLq9FIm8TgrQrFyR/UDzRDNMiEj5/CBFNPRNLCoWt96ak+Ij7
4S0kTozpMXl/JR0f96zzEBAPI13KFfCRjQZEmwCDRLnIR/PpyTM/0Lz+e3tU
ZzNxjvkNjCzIW5Edz0JaAL3JeGlinP0gPqj2fzw/geqxskgV9gMLkc3m+iAZ
SOO9REOUHZIgsi1C/i+p+poCW50YFJ92YMBPfnhYHufj5fJyy12iIjQrWXiS
QBUAjuqN7JMuAY+Nh528wjSE6cKPEhbyx3CvxohUyWgr8LhUcWew0r0XH9b3
z5jX+5ZAIMRJvJTBXocgX36+gJmKvh3lfm6ylwWbbI0XJTQm7oqz7qDHJaU4
94e0RcSf0lkv/cjxQwoKnouEpbfqCVSHQwVeAL8fwXBuQ2OnAcfnCkhA9yCh
wQIXM4T7O0+WpGQcW/YoVI/m7hFN30MLLi5KqKnVMslCwNW5Yv7G2mfI/NO6
9/3O7bqevlPEepZxDdnNOOlyqYfhPag541cUKkTzohYORZ5ub5Z51MOo+l4X
Gg/1j5/i1nzdl5m9BnlBN8HreY31l8gkBAaoNizO2Myn/m4I2JLzoloc+SHE
zWpY0s6QusQm3GHu2LtkoBJv1Mq3w9ByDCUqyEZPs5VUD3shuBmyaRUB77WP
D9NRZUWRWwPevrV2Mu0VwGKAahJStS/4ozmscUAavJHcNwKLrD+WP/Do++rJ
ZxenRFJ4n2zOvRpTmjWAdT243dzkfGP+D25KG9diDvhMe3ZsMFvZxqUkjLVz
u9nI5+fy52AhYtzcSc707fbZFmlK+erG5dILi0ZrSKrl3le8ejk+IyvLt40U
gZ/4WgehPmt49HZbkkocB1wQeNDGKr4wdir4ZkjUeszOHv07BL66e1K9IrhJ
Ugf0Rri3TgxyS/kSvKVQI1ubZ5kaXU35x3HJ1JOVYRHtSiz+xsg/IbK4ZLY7
/W/6DNY2/HvOWdrn19gvjiclxMFaim3qAc0AuSIMJ5rbM+c/uuEfUjv4Cx1Y
XPDZfye3O3QQBrEZlgsnK8mbPL8ajwOSQTN6CjSO95MkFC6t5iaSr+WePSRX
+Uo1vc9f+f1Ff1M8WKhLf/3NVZ7s6vr7HxCoL7xEyqF+duSA0RxskLOCpM5W
/Gv75oAdUkUkO80VwdUZdT8PaVh4go8MQHgsuIvT09EAluk7nmNWYXEwEZS5
6p1wgDEpp4f8qH/iUXqdy74AZ/DseRI6LLM+pGUa+iLJ5xEMypYjslCwu+Lc
pYi51riMKBnVPUeB4JbK4E7jrfSDIb7SJJ9FkhPLriBk3Ggl0Qd7Lk1+biV2
NFHc8pricgfoK53DqmnoKPMFANd+By6gFZR7XWDgk5EF03PFlquz1d227geZ
r9S1p1muSeLoEJNPI42LXRpD88w7S+UElnUAmF202zjTVV8/FaHlyy3BiiK0
BvZJGCuHsXtOY3Vj2sgxccN3Nom/gSuaIWI/YU3oFyy6fUJfdvh7def+HWOK
/ByGlejLZZoww1N44fXffF/h3tLeUg2INQUzHUbBUcF/qFEJhgpbLU3XFNit
dhOQp2Cgf/VIC/653Xa7fjb0pC0bV7aMjTGU49wwytILKUZkuf4i1sZVudWW
DHzfkgwsTV/W0DKvh5dBUuVtn9OeBlmK2Z9SNQDmcS+nf1FT4FYQmHYfWLaD
Wgg6z0i3MI9Y8wyGh5aU3coy8wGeQS9Y0X0AiZpBFQnUGK0LuhatCH64lVlj
Hw4MZDZfDnXLmDoaVrlYLzrizchwHDVQNdA7ZFZSATVEsxMrvPDuUIpEs7Zq
iFNmyiIaWwMlM4eigOGq9ceRq05tLZueIUI8ihfU8BcAniX80tj7icJIFJiK
SDTMwQNrcEwVr08QJlRGSOFpB5q9XtRyjxegf4SUUkbPZNOyrvokClKdGln5
qBxmDsqpFfisXYfIvEhe0/lPUPitEitiVQCfDuli3Nz5rxrtwI6iz2ksHA7t
xU22V6Dj7WmBZqqbAO4h4Y3tPICawUGEedBYidxTr9apjvqvpKh6iKDZu4gr
OrPgEe24FGkl7ejCIZK1+t0vWR5dnezg40esupj6yr4CmcqKYHuzYcxm+816
C0AYJTUaXl9Ji+/3KRat2PKIWWT8eBH0bZJGocz/b4kJluytlOK0LHgQ3//n
lOOGdqnnE8WdlYUDiMQeDPppg1mzeZ6l7RteKAVcvnr/UyfQHw0HdpPYQ+43
PnygqgSyzLqAc+Cj0FVLZUUiUvunhhkpjPmgztHxvHq+cg6t2/3Sc5B8mTcj
CN1xhKQqvkQwwK9K7S5CQLtZTB9gtMeFGbixF8AXetLZyxW0Vgj+XE+VNx6Q
1DckAZi7Bqv7KaSUOwJ9DOBzREA4T8aBAqXqUMe3ivXsqUYBPdZ9LPWqd++f
BsHlzBSkNXolWuA+I8wUs7Uy3qwYmHD4PISvxiwsjUPXCDEAjKosHEUKwERn
K2Mk9xdhFm1BBqx0ArCHE/vqaMQ8sQr3Vxr42UfRObbBMXgVuynLBxDtbGuI
+vgGMBKeWmTcZTO7OKKT63Erq+5tpum4ipWa+4iX4/ai6ClRTGk18Y3Zyj1Y
jmdU7H1PH/S3u0BpKIGq/iCAWTC4i2Rg2ZP0rtUSCrHlE4ZdLS22Vq0HoDjD
rEsiFG64Ve+DUTwZr+OsAHr9kqSqhqBiQ9pzsMdbOR7Cyb01CxkjUFi6xOAj
GNF95vy1l9VsQhA7TjNfPdbJrXu0cy+s8Aff14kKMxIA57sKkMfZAhhcP2UN
DPNNY6SVy2i8bBS5nI+oV20CSm5BwxeeY939PsIClWAiwNr+JhUygBRtuphV
8QSmbfy8YgAJgHMMLiU/Q4Um3l+VFvpIjxP4zquO62vdTXif/Jjm1553RDUp
BoJ6UlFJcvRNi4nF5zFUXg5HwZEV496KsE874/4ByWRvR8wZ7hOv006rQS9D
0S/mEDUtRb5bBZEZbDf67PmCI+3Yfr15KF0rUA6kMTRdR+cxL4pdfaYb3H/5
oOq3VZGQhTQRGMo5X+B9FfWhzd6tsKWGT9jg/QuGL6/w6NYGBwD+dPgqDLxv
pHw9fJiniZCopq7RybfjnqVIOcYrY9wMhkydHfLRvTmb+REgbZRDkmiN8OuG
yO9Cl+X+ZqiNy9a2c9f60S69W3IbzYCHpRnRXsmNJdBOKDavEhCL1zkcOMp0
zR2fHqy/V4O0MTMB6G1AVEMuhQ0KmCB6Ndppv5vW3FePpFPorsI0aeiRT+bo
jeIo4gz4npkSZkJTI/HvmNP3j8MJ1mqvy4kwRR/1X/vTEbjMn8j5+F6KtqUt
eJr7auJNPI/biCXJF0AKu3149kbjHs+0PM7Kz6m/3jqaOdLLiSUgHlNOyS48
Rr0aKqZfuX7B23hA9d9axKE/Uilx1FF7amVJtbdIbzOq7ud6a7UlAQjbX3mn
ar/WLLtEgRE4ep110fFq73AD8kj24noN/O7SSE/0L3lPUssUM+xOrnhrJR9Y
EgH8mkPC4QZhCrjIV60LvkZToxIpG3i3dlxBauuhYFRtA4hpURCZA1qpDCdp
pAUZfEVCfZc58vWiOc3GsbD0BPkneyoktIdqnG9diGq8oEk75l7HfQTzLMjL
aam+Hd24jRdok3GJIe8qJxoNPxI9S1srQwZeATEIzRJm4nPBvZfmr/MQMx5y
AaDv3X5w2dAz/Mpk7kDtruLlXYFKX3XYot9viOvUx7PmIfy+gOUsE9gONyel
9hD3UGEx7PoyZ68s9sFKRtWx35sQqnfrE5mjfnYdfWr+sO6QHSr+KxzssxrZ
80mn5ZAfT/l4P+W9S4mqhOpzUjpTC3R9/a2JshOdG6dELKlJwl0xMnbpXB5R
DKChrX0BzLx/lBJklPRbcy1ARKTlDyye7VUZbj/UVnxAMTp96pLHIRWiGMKw
HZOhFGBaI3R57hQEBtvZSpWDm12qL/+gETztTjrnTrK9WbEWgYR14nyzOE5Y
TtcYXnwKzsfp3VlqdgkhI4fJy8n7amJjw6i8mgyzsSfvhUpllMQ/ExnaDCiy
Uz7RjxtqYkKJ1qA7zQlD3VusZU6iT+sNgyTvUHeAuVHVo739YK0dbM6examU
JEowoy6L+sYQUkiQMW4Rr52WOpKmqXwtv3YPU3QdAGZBa4R6Tl6I/Ke/fEHS
YukbLGXX3rQ7kMN8AHVXbslPG7BqOgkEbLaWZsBWMyQ5eHMMDabAIuPaadD5
Abf6vs76GJ5eVWTIkzd/zgulxQZ4o6m7dAKY3P4ESSmSjRfxxDoJsLSPw4GA
/bsmPCgkkq9Ez6jjqDyJ/NTKyTgHkZMOOyzIOO+PuydjhgRwLdqK8AJ8rFTs
KkzuMbjjwaQ+c5NYElUhBSwZ/0vCMi4KkoS1ZWp1oS2/ysEWIdUNPE0zzCp9
iIWaQnmctk910yCwh/1p7scxs0xD9iJyk7vSAxsoCRL+6xWQ8YPtGCHx1g7b
wmAUJs8uAJW8Dt5u3tKf3E6QtelT5fwb09Mau+EExTYjiRJ93BXNMez4rWvR
vAEnCVnsKlQuJTJR1kzwnlmUXZ2aDOS/QgV/FOpQlJAFwGfwKtr75oN97QVR
OL646iPq6dekbzjBoCE4pBhD6MgSOFHN+HC/0GW1wzY9GFdH166MyWy4DtxS
AuOprcXQQu74yLZhp0tfV/Eyffl5l2o+udaPWzYgjpkPmi8tZa9Ns/QO0nVd
0WLqRRvK0KTuZMdqFUIVls0a83T7A5VhwHSwo5iOCoADlVNpq8UoVz02MYhv
otchCDYdi71HpeAFhYzShKUnrnnK7xboWqJp4rOHLF0ReBIAcjyQOs7S4b6i
M6JnITaiUa0z0vwnLmNqG60/s3G8kDCtU0rMYZMM4q6Mfx++5aIGbXWzHRXB
/NAcjFE81KTQAlFmNQwff42TaalAGKegJKPkkCa21/FtvcXqJnXQkdXc2iKf
E1Odq4gXNhuY0G8dlUUuM52fjKkFLi10S4CvF6qI6rsvk3Fc3bRmGzb3QH7c
nXHT0GwuJZ6s7zhiWrq5CS11ouRVrO3B58Q+WC+lo6yCi4fAM26JQDerrTov
Ojfx23IWyb3m78NK3YexCo8p5B0VNMCu+j/RT0nS9KUSIEPZCGi5ExH92wro
6Tjl7x7vla7FXPizLtK6m90zOXWmzm7qSOqtfBrbTYXMD1+JKP/bbsO7/6H4
LQbbRedfFauS6qQj3Y6KWuK/gAJAXDckrYpe2J9zuUkHBAxOxuobP4p2/Erg
vxSijLq5f+yXDxGOiJ+t2ECC225rYaUR+Dlf/jdUvYkrhh9Mz8phBkCw5E3W
CmXqHUoqHxpKUTlIzkte8G/2DvF+iZo4dqq8aCg4ZQIILQl5mXT11Mw5qFNB
H+UzHsrxiUN9442urUhxTKGRcd0+W6sezycVJi3L+fjEuLRik5vpMs0AoWCH
8ygETdAlJ+bP7tzGkdD1SZssKFJpkMbpBNy1Emsm6A5LiWNaV3L/HEWcxDo2
pWG8/N3XO2eSQ5KT4Ca5BPPlGmaQJQQZRd8EvleTpTtElhD5AQ9jApKVTopi
ORPSqBjcKzhajVLVJBTEdxBGVDvLfivb+ivuFIs2Zj2kHLtPBlU7MGnpIcNK
qdrIJbzP7wrNfp/9Ji1qOrzBVa8x6eKagC6wiWELFwxFfvjCVsUjwq+qmc6f
YpLUIkZWyvmeDG0C7puayi/yG7fknSgpjaey7f+WuZ+pc3ETlQHbY+C0feGt
p7+LeCFs4KLe46KsuSdN0hMu32StmSAaPMdB/CPttHB98nOU/OB8YhII01OS
36TuybTb2EJkIbu2NiltAVlO5JbWPnk77iSn8XhLNlydKs8SgPzo4RclcQBD
Kg/eaYStSK6LVsHOAqskpkKWtQroowFmGwphQx8n4gCBiGdZ/+nCI5fmCWfM
8A6bk61+zeTH29x9SOvk2xoAiszVm/VnFxYvDropOVXOkjhAMoa8itNYuNhF
YRGtsQO+HqntcJpl7ToXZdvHqmrhhcxLgv45PQDfv4hu5A266Zk2eIh8j02V
U4j4uZEsrkgyjH4xB8xMFFJYaHraqi+igbocVuGW+kHh+ayyaZc2dlTtnfp2
Lrf3nr5PpPyeqPK0yNvkCK7s5gdbfhwEPHMqgvTZjCQkuETCCsEeUkhe7HBd
ojEqIUbr8EgxpOnlW+M9rU3QGgzLdZ96wDPlDKtZvKTyPWNWZU2q+mAY0Esd
wBA3Ha/8Lnu4n07h7yIiy5sJiqSEHNhlNE32b5LncqaMA4jiEFNw4JnzRapR
T4v1xFPfuDld0rVE/B7un4LRI83sB5IEDHmDuioVs3oliXM71q4YeZlEst69
cif6fPxiHWRH+8Q6ZvKM1qKBxREt46kwOIS1Z0W3mkk1oAKLSjFIqQyPslAn
NQbHrrgsVJxWJ2yd8hbcjssVEp6rDQ0Qc0jWilCJ/lu/6KP5JnfHwnAF+VjM
A5x2dllUm78LynqNrdYIGvFIzgCyIyIPRedMOXLfwGYZZDP9MhUasLAn9NTN
wiCXrDRGglkzh0140gGWyBASXr5TVUOyQ/Ek9mCJjFKCyKyUgr/yxEHD5Kk1
EDqPABhZr9XLfjAwYhIN7wQugIakqd/v2ik8ywu5tKBJI3tX3nyb7ZRzmlSx
CbZQtpAWEGOgbUfJRIZgU6yK/pAYJHK92OrcLgqI1cVp/oE44xbF3pi9FOvL
b338gzpHtoPaj65UQUT3/CuV/xhYmcsDclDUZnuztGtcgk406UPbSYD8AV4M
af7t7SxT6bSXpRsR9oblGup/N3kfKcymf/GFW6jGhkYv9zisBuPQ+SRklkEo
+S1HuA5eJWRmW5CQqu1N6MOIdmAqKVWWgP9xNzNJhgZYQEzC0tAVqf656rVW
i8uX/MT1Aap1WaFKTDrWxL2uUlul+3UhIrWYP9DSijH4Bn10QdVSL/XzLjE6
Y8g2dEayuYBEbuW8Zj7ktCEVhHdZOA+N7r+/5pc4UUUcmEZaCwxM8dPNfaZE
BZ2kl96sWAcwP39DtrsPvMhSQLTFfQKRq+RpUwJhesLYFwzeTQikjQQK2uO/
grOcpA2ZkE2k531TzAcX5sNLOt2IHuAPRudwcIDOXfhoDmmbJa9EgBLUIWv4
TUCqqU1PChXUl5fdFKurVI4URRIIgNSbPMEmbuKWJxPvbqxpkbb7sEcpsRCB
0KubXUD5uGH9V9B981hnJ20R7UUQA+Uj3JHJGOErFQb2NOZO7RL/WR1kjJ5F
LB2tz64+UWBxj1mES+gKLChN+AZvdclZbgRpMCSi9Q7gxDFwj2AJbvZ57xsr
mSngAXYPBJrzxR0a2FvC0ggPcloPDtQOzRQOPSPeQy/F+5ECwCEhwaw+i8F0
DyJKturU/6LKC0bXt/9VikTNlXTOpYIUInHkR8gbcw2il/0iitRRiRYjp3hB
Cxpj4iX9QSxFADHNHDaNv11H63TZuh+9cVSQRTvCRXcxzQn356CIbRr5RR/E
W62U5prgn3b5uISGq7RG49t+ZQonPvJ7RQMru8rk+ATalipnI3tbfN9F9Grd
bhwaHzPudaY5BeK5UszFyTbWaQu1658hZQcF5XZmNdhL2wxHq3obqDLgLdZK
QBHZ4q6feFHZzr7ttG8ystw7/vSHuPkUFpCaj4xn6n4R32PxLbP4+FDI2JC+
6B6B9uC9BmkK68eX+4fwJsFNrlTXWAYdPDq/DWFIj4yoBULYqcojX9OfOHdP
12M01o1uq90gC4ZwCw0r1FCkfF9ECFAOKv2JCpxzdcLJThQZYvXPpK4tJ62x
BjtR7HBIh/YY6pQnciH9r6wgwQ5A+QGYQfs0LuOH1wr6TewfOC4MLrqnB3fa
M6eceJVvz8evGzBXOrrqX9zAQ5XdHhAetEuaE7fUJyAgu+qTIwQgul9e2r/Y
fqmxR4QjeTqaBs/DAlI2CDgAsSlIjPArRfSYO+JselJU+9huIlb0oT+ai3by
LCc6FW29IvQKNEQ/SK3OotWGVjnI4g4aCbcNnLwLTVYwDIHpl9CN3AbBmMl3
7+ro7tSVyBQu86CectUcUX+dQ/7sxL0Aiib0n0Fn5VmA4/bsBdWUbv2m1nfN
vL9x5KP1atXbiYSep7GA9ftNnjQwB3fg8+TfTwfvZdLPCGDY2QD7kmByhJhH
HpHgFb8Qo5DCU19vD/z3IMhbDdcBqYQ+XXMkHwDr8CaDbfTZdgDdfKmUdq/p
exJTmyE7yenLpRcSuKkdp6uyMdQ0mgzMXXMwzSI2uO7jKYxL5gShXFfpBoWh
/pdSBt0MkMr9RlUVwvEU9gxVPgfDttv6HWwa55w/1U0b+sdc4+cZj4FnIC+b
yTd/Vj1CFKyiAHRT2/SoOJCfdrOXWeHtn5ZO5Vnb4Ck+tN2jAN1OdsmQrSfc
kV3HQGTuq8Qm13A1cQCqky75Da8IaJCHKgc0AxhoHomOJkYdX5n6xH3FAUAq
n5mW2mdj2UQ3gllIgT6/6YTMIQsHI8nOSnq/ZkH3koBitriFSnuQ9GwOe0gC
QeHVTTtqjQIX7am2TxcHxTaH3o1Cy90P2HB6Xkk5Mzzv48mlglBeQjUXXRpt
z9s4RxncpBrp+j1PvQVOF+l6AeyltDHmuwX2ZZL+aYe/M8an3UIMjycFsF2G
0CA2YPlEUnpT4AykqYx4yJIfxbrvxqAt6RPf3ljZfdx4MGL/VlfOzhXmFzoF
GAEn0OYHS7NRSGyO7787UEW4UoFTBsQLPzbwm/mwVpde71DBNVCfwNddyX2C
v67KeZvTEV0dP6g9O+i8vVFdRFiXgK9S7HeStXUXaBCiDOlNsuH3hzyOM/oA
1646LFvEoblmfPFe011V8WspzyVbx80OF4BOl5dzX60FIRg/rKZn9G/Re1yk
ltav3auSxCnMl+n8n/+CUaQalsnWfzUIYBZ8pj3qE1VoxfLfW1l1xkEmdcj2
3oQ425g/hjiiAt8pznLhAp8BbzSEbYP7RDtb0mzuTrKzqxUKP3SnwlW0K+kF
ZJ7B1LeeDkStzmip7EN2+GRedSbNkyHZfLFAEudRUVr4kUYcADLu38KpozZc
SvLuqp/pOlYT7myCuKX4RJIYLfM5f1dcy0z4gHdakGO1MCqsGsbp63Wv2ndW
1huaopwlmC/L9bt6itbwn0+pEPFhMjgNVb2DuNvNLYDkY4sKZcsm5ktqAtSf
ur/hX+AfTSBzQlR8zWvIpfoklC/eA3eGX/LUGPjiw6w1h7ewlZq2hPAYFV61
CfuPnXc48vBtLVZyHW8/6MQ1JcoFx2UD3c+NtzO1+hnZ++O/vaefsyufQDvl
jiELau5x7/SFdJfwmUFOP7S+MV/djJ3UdzXqX6hN7ZkoutDXbUOscj2cbYwR
FndbcYtq+SPUBoNzxFxYqZp68hejPDLkaJwlaJ4FVjzedDprDJqEAZcRrsui
O9aQ2yHftWNK/4ogQWhwrQTLxOISIngenUeDBCWgqjIE2MXNEy2WMfy9LvQZ
pZmJnGaDj5fXFVtSEzj1Lh7zYiWz0gADazuOuA+7PIy1nkvQ2xmuhJbgOgOY
HdBU32kM6DGos++CzTpxOMLc6VMmwwRVOMfjov3jM1yqWggkFeMOYn1gXCIt
MM5G3Xxxkl+GdjotJhi8q3Jqr9TmKUXnVryhtj46e8Cn2TNSaK5HPc0zLILW
n4lyYA6cSsSw5rSs81hMXI/lFki0IxRixBmr8usfBsyxN2msO0BH/WZN7QEt
/xaYbR+BUcX5JeYeeMBa1VfKdqPl6DwnQhBuGFT2kEwpe+5SW7HdkV0l5ii1
ccItNvJsfSMF9uquyqsT0K9aIlJpPMNjOs85yRX4401ONY5Q4Q+Fys94nU/I
cliMqSfPWol86hMmvsnQpArabaitwcXWJHT+ejZkB+f7My7m2IuK/fEEyipu
1Y+xJvDvrwpwMQI4PKlbxrQQP9u+eIl6Yc7eszVrBHKKdfP3lV4cTUjZeb1X
wbE2nVWlXn1alSG5djvzJMZpBNscqiI1pfSrzrc0KlJKyvSDkVjp9R0otkaD
pWGDy04zCj7rorSOdn8dYIlaPPnZIzJSQwpMdxuZI0jgo1SD0/pxZB17d+gn
k0bmSu6mJGUtudLgUn2up3E3eI4VdhC7TnPlT4Bc8zjP+oVivppqJuplDoWR
jcFhDa9WebLkXDUneH+qyFDyWziTOYXYsr3aCmOM3WV9AMZMIM1VR/hlp0s0
1fmaYNI55GrrGRpEHsyPKG5q9Myw2hSI6i7LGXFKhaR2DhQUHmuHMxseZhA9
kmSJ4wTPecxDn7DvyoejAIrZuDHeA8o6EdJ+vHhAqgKMMnulyBeCKIEjpa+X
1xUR2WEewOzIOUPRaVwYdTTywEV+ElzndDdPC7wm07Iwn2ohzo4yNqCu4LWb
4AkdVrzMEAHzNwRL7a4a3D603uG659WIMHNp6PSce83JGtouCec+OvN51RrW
HtTDq2ECWy/TTYv0/T3o8LGHmRfHXsAGD7pVtf48qSAhr0iAuJGtuLIs4wCB
NmC3mOq8z2uTO48eWycsIQLDvpd5ogizfZygNIvEYqv2pdWeOCg/37gepj0g
II5DdkzfZIZL+wPeVEuICr1tHDnuW99+EU3fm6lAR9TBwI+l32G3HVjfjE6n
tZweoJ2qDb0wpja6b8Iq6/8Y1uvQqGxNQe3RtC+s/wAAs91Wtc18qx3LGp/i
3qqesPaTaUqveiqSPAo0Rfs9mWwrBdBgUKDV9Mx+WMsu3plSHCX0uu27ns+J
T9Ttl6T6Ldzgv/7VMPDLV7Mfi2ZkHRTiY4McOf1gN0HDu8LsjtUNSzzxjtKT
4Rk1ClY24hsdZ2kAaX93YUHdUm6fBE7Js05lZGNX6lnaCWsWNkGuc0/5gBUk
azcNdaJFQFtUYgms0jZwE4mKbp9yKNnF3DiZLpzvC76Um642qxwz1Eo+UplE
e1Ougv3K+oClgO3y/gCyWdf970PHroVEQhwW16BpJHK7LsGIltBm+I3tbGuK
LfGyrxQ+qLWxV7BINTWRW+zPrrHm2gV6khbgp7nw38BXJo7WbgJUfzu7npCT
lHXP3GrYECmtBORGZa8kjcR6vJDsi92YlQqHdajUvkyPEPkf/1cloxl5F2rQ
mf5vJCCIA/clZT9TdSVDQV2AxaDBdbBrifz039hQEu/Fb/bcR06smEx4rrIV
H3T6Uj6FKB28belihWcLm57MMB0VItkWdyb4r0UWc5oSRCNU/rtbq9m320/V
SenzOA0t8m8l2PDQpaWA0Y2Vyq3IYUtZvM20xLVinZNVyjJQke17muRsF8Fy
gVB+TBweriUoGhj00NDQ7skncT+03DuigT2Mk1RigmoQ238JKuCUBNz0jLY+
5Fzvq55Qr0jzFR+6kLgu0AT3suqbelZ9iEIzQ8picP1PABAAlKXy/bva/zFt
O0CdcV+KZ5mZaeYeQ457MpxDubxpPB/8TY9BqS6wMueXz6bwTI1i08Y6ddFC
gIcjfYwIUH4flCxcYc+Q8g2AWIuOqGUlnVI8021o8vdqrBjw+5nyZG3UObHG
OErs3FJMKJJUiWwWyjLsqvR1IqRH4vhzzWn6WO8S2IsmQikLAHU61/h274I+
qlI2ZuYgnIlY+GomzZ1i6KQGQ3bKBLVt78s97otV0rf5wXx1CGDso/V4hJN6
Yb/ugEiu6mJCai8IZx3Xb89QLjf3v3EM8rX0Klk7AQL6yOA1zTu4Qio89KrA
4mFJDX0IOKymCMx9d//qa89JT/wXWW4R4skVVW9zghcSr+vSyTG9Wi8sffLW
m2/6Vq928CsBtkj0Dt7IROJsEay1pTY2ZijhG8Gwqjofy/dU7TcT2TrR7fzo
WDwR36YkGsUyoWbXIvf2KHLxpnuhSOtx0hpOdwgc0JVLRWz3fnu2OSrCJWJc
1B+u+eBdTeRaXQ+hui1Ut6/qOPx1jNx9Xp52kA+uWyqzqy+aLHLbIeJFUNAo
bo/zi9VNRZPqDOxBvvS1u+rF2LsjiPlT7mZuaMQlHyVig4tuPru0T26lE0bx
GG4zjfR6d95/NiuCSxxe0qBFJT/J8a0FYCDGW5S4W9z3i4X6PBng7oy5zTZd
4RztNN9eouxoSHQbti6d/i1ATMTLiY1yMFwbbeVJ6zoxdWo2ArYT8YppW0or
YHZINgEkz5BmYB6HwMEOsbs4pNpl6czEGiV+PFvDEs8Mv5yxdZuNerNND+Vg
pwYgaI+I71WCii6bO4NoM/q2NH9VzZzCOLQT7blPnxl+uUjnxbF0SKQts2vw
u2Pi4tUOxfH5CIEKnSpEqJiq+TTZRz0YsXhKUssT1LpPL/phxZe4Nu2Y693D
wta+s6xwv4zGvl+anQgF/fr9jOwCeIRySS2BEq3T0lVE0iZ47OIiP3QLz2f0
DvY/LIAyRsUmfmQbU/X/buvhc0i9kneY8L7kDHzT3Q/nIAOqVYFsM0IHj53n
viRlFUXE2Ta3vuX9QQdoF10QHKHKnw+sMbNYio96WJ7XmoncXOGqU4/+YbKt
41L7pmh/G2gfUUFZNAEcfQKsm2jgNCF3ZWz96W6GuidKa9qmgthy6eNpFu2d
/qK7wR5XGuht0WFFu1AhtR1d5akzOk1y8aMv8JSFZUE9+aMvwNWXXj5yGgZL
6k/sGNWd7kwJkYvgs+cgCJsP6Cnc5qADcX2SeMxijy/vPPSPqVJaOJ+3/2JR
AzGzUNTHdR/rHskbCESbv5p2GIi0kw3R4ArmUeJGF/H6QkDm3ZbpU4wi/w6R
K6DZAQDQ9WsGF++7KTDlY35UV0Y0Q+xDwXsC7zOzWYIeexaJplu9K2+GzWmw
T4JWSTRkJh/754FqOCN1W75/LLe+ePPysWm5tRylu1nmTART4PDyawEqKsUn
0zt6TNPL0W+hcw1yB4DyhoRIZRXTTL+8mzCAFZGzMRSeXxHtPKbusTj18pjW
jP2UhHSNag0E4A0oT7eyu/NfzVJsZs1uqvCE/696c61zy4OoyVqQls1lRlZz
KgBuo8U0lafke5GPScw5lHufr3GUPQb26WmlACh61fp2k+R3CdHNqNRAo8ah
Dzccm6OPB5XxO/GXb1YLOSnXdulSDdIPNHQl207GiKMVZNwPGq63JoSHYFpH
kuxSE1cz893ceZftJSTfxMt3WoCEZHUQ2IiZnK41Bqm7AlXTgN84bPgwpxfx
c3CkQhwvaGwsrIqV1sKzgVQ4vYkp/4D4tA1Bv5D9cDMYoILeYTPgbmI65gR7
kSVS0GRVqRXK1HJovNP++oUeZDerO9L6KCljch2QcsETK7H3Uly86UhkZv6Y
0w7Yo11vuxYemid47HYPd01iVj8RSRMwNweY+FBiYD7qdej43dboAuAbmaPD
dldCzxZMq1uchagLEBDDGjxV6pw8Ji91/silw3yMdfGGuVmIKqLUXnHU0cUO
x+PrO57CE0ql8+/C1dmp4HvaTqwvaORCmZjtbU4obe626601mzP3Zv7z1vml
jUkMcTphNr0qkEx3+Y9T0yPaWJ7NEKUl/+MxhZ/OsP5aQ8gpkm7LGfeYk6ML
zzCP/YifpCU84qQwC1/LZOVRi//1N/5mNdax2o6zDtIm0ZzK/TLr2dAfFN2R
JNJytvB86t+7M5SzEYOjlBzkgOW+t46tmWJUFRnjMqtSrhTxVAoKsPu+QFoV
Y1qgd/WZKb5r3G3RdMmdOjrsREMjVlXawau++GGdIFvnJe1jQDJIZlfos7gB
Ql2fXAmhRmLnhdurQhvruXaL8Ys5+O3M6QxlJFsUFPuAu5Z8djSD/K1RwkcA
D1igA/VxfvKn03HSOWD2RB6TWjEeXzqDJT4RcfAbShWi7m0e22kVv8J7spU/
Ql3kd+wV0+0CbvImgQeJDwlyrrf6Ad2sdAcPa7Yt6WtySOqXl/sUsDxP1RTd
Ay5vE5EUEOBLYSYqpnYOaJ3Emc+mVVt+REQ76AxmBpO3hJFF92ajmWtqqJFU
kEf+R4lngtGtBWlBWQalSx330qn0QcJ31OLss5Tpj4Kjdn3CSi8eeCdPuxyu
VcqLXNfXa3qQVCogvFVUqfHJoP1AygQrvJPiP99NQ4cRMVOimsqQj5cOFxb+
YOl6RtVTS9PDfNbKH9vB1rH2rwrml2ulwzQ5FNXAvlTMSUR4rSsfF2v9piWw
zFKBHGMxEOqBsvLEKDzaQ7BXDXeBNqXVJ2jTPEMC50ABAJX8V8T1QbuXmpnV
n+acsIz9ecgDffbGp9NdfYFKk6YJTK2VVk5zeDdYyGHi/LJsbuNb4O7ryTvG
lM2wF7iSrnEXP0LYM4nJ5FNPHwHvb0+oFevijk4s3/AS7W0rYWSlY8mmoth9
5EdYeKZyT2VA0yQZjTtAjOL4uszGK7X4l7JfHFJOvS8LRqg3gwdRmZ1PE7QU
P9HD7aAumh7zlyPVSOsWHj+Q7FhUFplRo6iGWvOSrVJ/3ZVY6yukYa8z9kL6
Hlch0xVL8UT2xVCtWbLM3CTpic8dD3u9ahLk4ZZW08mTNnr0+MdaQnAw9Ujq
T993vA29E1A0sUctWu5+LhKpIk9u6AS8oF8AfDLzAro4BouL7CZW9kK+szm8
fbkBYhpPaVNbVulfCPk17Rf7cUudbGDSVd+4YWENqMVgmsdyqG2fU66pqR9M
y8fwLtwukZas47ztN+F4aW7SyjwrEw4YWTJZeG29aTdku3xsM0xtUMPRC5uL
J6wzZp1mOEw79u02h4QFY0iB7ysViHT4x6L9bzWEHPhj1Ef6DPzc0uWynhlI
HpoSG+3Q/5tr5y9pMZjZXMyHQrgBlK8vItwQApAid9ynr2E5xdqCHHsSe34J
Ykgc8lNx+sDzg2pMh4aG2wqjx1XyK8oXrlC4numaC4UYYi0BHgwHm5QOKcO0
TkrGMj+HpdRHwk3NhGLIV0giBf5iU+umsc7QkXz5GXn3KxSruuQ6wZr5961v
IIUcQGerHHvvzxzdIk+Pb1Ccw/mbzym+DsUqdLi2TVOVcXvIh/ZNgjYnXXMr
ZXQlEKZXAl8qfw52dnH8bkCqIkOhBHvaSkD1aChaJf9J/sMAANVEqdNfxywt
rGyrIgNoB9KJkXJEtaBo/wF84UZZoHKKmHUIpeTN9+PAr5m6NYsw7oMgnCH9
9DWB+nUe3B/tHjF7oySWr1DHQ6Bju92zCuEcUggAf90D6ZWwnmqt49ABVW7V
SlW+wN/stIIAvNk7/OHCHhEER4orkWt0e6BVqlcXE2wsolMENZpj3zJHlV+L
FJ3QfgV+7R1FM/rk25Pa6emGBMBVk0ryfTiC9iiG2MsShUbX3+mgDoXZJK/2
s85FNZCGwmE4hU77wsTp/V9GlZMv0B28/aP+bYm70Hp604pu+/bvJL98xcDZ
KRBTm0RBidhST905pcJvhRWVR/7jvgP2+yqkkEhPrvymcOQgcUYk9erab7+g
XhjeoMTM8agc/Cy+2ixD12GQW0FmEyqfruI1ip6edqWeJ8hJROqQgTZB5dvB
dlx97Q0bhRkAOjmckA2wnQI/eksbdBcvN0pd4c9gifqIo8OnTConUopOUM3a
Ds4TMWoDAzD0qdzwrp81c4RvYVK3Gl8yBef6WmKyC5iYZaTuIubiiNb9foeX
1lVojWeE+uPGCMOmu/zUfKHAslXio9gCDFA6sP9L9eoSyPQEpYZUfx1by3Dz
Ph3rwtB0OTQf/ri7FrhwFSkkLLzqfGVnTrv73yTIor0HKh66uPUWEEeMK7jA
t2lHlGD6CgBec16G4LgmUEfVRfHKghXymGCi0Hl7NTHDoA/nLRpJy1xJYDvG
bLQa/InoxZ0CyNR/rqZjxn11B0bL80BKoUWhrzyB43ijW6YV0lmbSLLqbrK5
CfYu81M16jt59i40X2Ds2Y4k6VbDmOs7JvmGtNApOY2V7iiwvvramaJ2zgyy
WbAhWRzRGEHl3D0/a4uweBQJrKcAs8EGpcvOMmOv5AlLdF0bB4i751SsRVND
iNpUcRRZSgQIcRSFXlF1I9ubae+7pjLOhSr7zULsXxMAke0y71ofnzlgYiS4
FYmKafy9SkUsBjQchFWeBJnISGA4gTX5GIO3aw1+OwnxRxYGyAeLu8z5jkNz
9JYp14WLngjMTB4klgrfIAa9Abt993hcVaGDlEqMnZ9MHp6eGpgBKXGb1qUX
lXibJl6ysruhRCgBTbB+9z2pSTPHqQmISKzQLTolZ51iw8jZBlwp3Skvo617
Ahi/Hnz09d2VtSI6hT3xvu8eEC/nX3u8TdbUDek6tn6h5CAI2VLeUNN0o2us
xjB+cz+26IqMevmPWrNv1VhqQKFU80l3IlvfuVuPxElGDxMt0zn2bEPzWGSX
JCg8MVeo/OTI0IViCFVHLNVGP7utxZn4RHgeFf5a5gNpdAArKjxbM8KEij9f
aklZvKeEfC6D6eLFLt4yigzv56glLRHKxvhefnhmAP2cGHFbcpx8622wa4PZ
4Un3lMEkFH7aEELbgI35mL/b3LthIhx8IuNvKPWiJT8u7PFPIJLdh/e6bvUj
IfXD3We88oc1y2mF3zQxDQjrFZa9EeCu/sHWqPcDZtJVZQIEipX00zDpUu5Y
6b9qH+I66faiy2JBF09Ngt5rZHMR+4PGIkGmkp9Zvc7NKJaGrVr7B2TTtNT4
rHxsTiwPRjtyyQ1gEw7IvSn9TWBOgWebU9BdJD2n3xJDn6/Xc+D45xRTW/e/
4CMOWL/QjrS7l9oOcDe5c2h+wQiPplcT1euKtX1WMMxoY3H45aU3SG7tki7p
qN0esT5gnVtlh3Kx86lBFWh/VC3+ryv5Y5OggHELOZcnDkaaI6lFlXOsPR8t
vT6O3TtAepLC+H01i2p4yKABmFUxiBBsp9pYvwz+VRjj8UZnSs1q0bo0D5/8
dpnbUqEPlYYfYIq/TIeGr8RgyUWKNArIsi1TYQM1gOEfBxC6IQMrP7+n1bYY
U7J1xoBNDVK06r8U+9fcyos5JaaSsQqISfjeAbmxzG0jMafQ23k8/2i0hFDL
la1oetfFekziuKi0pjV7Jm+BaDzaEYeawj7Yhej7jWRnGJCF7Y5mTsE0oLVM
d/H/5MveupWUmU1aW/Kl9eOksDfad8uTb7DUIwLDNo5q8HckWEfxjwRKzoUD
7/nDURgVy7vOpyJyKzPG11VDOYt5GvQ/bruV1khfxK7B4oDNznY/UwTCaWA8
pj0iHl1ZqD/yjlgeoOLrblm59OhTq5RkWZVrEYisNhddPLG05pF3Q4KFCxct
CIfg630HWp/AE0ZVtK4I+nMzYjGKP6DTXKlXiL2L7xrf4xrGdWBTWk/ZoiH2
oncm5mU9heWkcSCUx0aSgruriUNNtn4nf2647dM6J+ZbL4TaIcEtF5HmGc3q
HEvVqsF59mlEXmM3Z9v/gJOGWhpWDh05pMmTWNnic2u8G33dAc767FwwSbGo
k+KfYWIU5Ujgib3I/FZd/ezDdT2jTyrag8QxGtIlwErfX5LpiQJ0HM4CAinv
9t2K/TtrkeCx7NuZk5Yu89KQftOZWVOLpQImmdxtl4y6Ei36vnikQjrAHPzi
Ob6JiKbILHu5sl1gBTDDPTODAg0CfpHeyYr21dU0Tcp2SMIOKl9fTuFRrTvN
Qdwq+0sVFLQs83uyOnLO3Jkdz6ZDiNxESQSZPQdKepkTBmf54RaGVdpDRh0o
jQ2miLQB0Cvmc+slIU7GahF4F+SL/cdefspCPX5gt5mEgVaVvPlcaiMsOJxX
g8P6927DPPwS8K9l7pNU6CjO3UEOXA/67hreVOomg7bLrI1KUrRjeqnP10TS
ZKfXwM9R3LlX6wnYHFcGYKUiNAruJ6SRQbkMATBBbaH2ek4hV6f1SFQ2qylX
GvQ/k/nVwYgLWgKbz6cha6qaU136eRbkzgC2yRCfToSnnz6CTjKaPVYDkQ+0
JC9JDQjmUSQjiMWe6osColNduznpZZyPTmLskwb+/1Y7U4qM0DpI3ZrW28W0
phfkAJl0apJKnVmhjr0HEPeIj3gRbFpyy4QaXNXePnAA1u3eY+xVax5y93x1
js9uf9ShbbMK4NQxwtExurYgs+C/stARx1q1XF9oDd4OU2sDq5tK7VpFl8f1
JK0h5GXYq5f6NLChmCr09KbfuYIeiZACBij0K4dyhbc/jyNTMgMB9h7FkSoo
0hZYpep2+NI4/0U8DbTLjjCCyqrfTLRr6qMz4p0U6nwxFypkh3D5MZNc8uOa
MOdZon3Di5gBMM62iAgQrmAmLKPOmefC+/NvFP1odnPsFqrgOkQzi4vPcxpT
FMtQo0K7sFXWl3hwpgUe2folkBhkrprOXan9RYs5lwz5o8XQ82Kv8Vbw3S/N
idOvj3lFuxn7X4HCGJaQcA1VPtGpmt1oxwG4p/KbS0Hazl8Txw8BuaqO9+FZ
LTBv78bN7Qcave6uhvxwlLtVwoPv/LQgjPZFVTf4HtBA5dPIy3nGj9i5Hz6E
B3GduceGYrTrCLQvguKn+dQux2xebm/kB5IjX07i2T+lJ29jpG4T5kP/CEx1
uR3qgNmdAZrropzCruvpFSQLn37CYJ7AATspnIyqbCwsHRDOL6cHFuVK2UoN
spWFGboAZ2tpCc19evPmSOV3z3Vn1KXX4YPnj0XjmoUr9tGF1QudDHALbRRy
8S6+6YTnF8ggDEuX5W2PG3MXTuw8lYmYTHyh50JzCoZLJhS3/JnE4Wf2O3dx
kp9o6L4Q2JaMCOPaNo8M04EnJtyQ2grBh6PznBKsVkhVaccb3KD+GvrSt3Pt
MaKNMc800e523+abbI7HdnxwnVexme25k+0NJqN8ZUQYx9mVpFC2EroGWsfC
tvITHk+st0SJhnzjZC7wGjugw6eaJLfNbs3/zzaZQ5wHjfvSN6VTfqoYscg7
DHTYUnKe3DeMTpHmscFsWSxf2FNSeOM5VQsi4GQTKY8pEE7qxobi5zsDokC/
DbUAA5cqbFgAGuYLuyu998j7Tw6gV9USZFxhKGX/z2CqkGDZWupyfx+Ntr1H
byBQ59cbOCaETygeBF8utXEHPjDmYBLGirfOIuSPkHciVG/yFPY+lkBAgCC9
mmMWIASKb27759vO7VHD5sj/HKHQXgX9U6lUVTaK1tGPGSing1OWc8GZmgM8
Cj7x1nTTCkIdgbX2eRpSve4I0v3/fBL3k0YxNDmktdOltPpAjWjk8uU0f9px
Goba7cezB+jwJcoDsbTiD1bC18JrfWtNNP6jzDsO5yMCY+DGSK7BwaMxdH73
oNF+GOz86uhGmNuNgk6ruw+EVTKmT0DboLQWM3NNVxyZwrbmUF69HF1cCW1g
5nhubqAUP3VtE/4zQ1EhndTM3yyJsHSnduqTaTaRJ/LbkEVlq4ms+Td4Kvg6
hKxUpeWV0Oyg0pcUTefHSshkb18gM9D496r6qALfOvGrekdzUqqm4yDK2CPP
s0LyblzVvi/+lkBbJjZAtIYRgWsKfhndj/3glJC0rraZYCzbPli8zsdfqalr
b4mxfXl1ovu2h4ZI1tblrJrgG+2aD9ePoixdthaAbxoExKcNtDLhyjA+vxft
GiOZM+GJw4gy9o4pW2+SAtAzgntVTUhFovlAaBfJBiNjrIp0OOm5YfFwYm9W
w2grWFBZUNo25bYhz5C0Q/QkDAeBeLjeVoR45r7WZuAJ/zdYQVKRqAO09CC9
oqhoDlpcMRjNxkffeY6Oc68+U6X+O7EYuXXgB15qmDhcCYgF1SIyYs5lU3IF
Q2cJWAyfNgHMpQcswP/pouGEJ2TNO9MFKl4IXNxCwVp3ulmiouOU/jfK6cnG
uvv54Tk5gZyOD3grC7IB/2ieNiqKRwwhllL/bYfc7QiilIYz/Q91G/lul+/z
vJer5W/lab+M4vOWPsRD4emdyt3c0bRvy1AYJz/57E/nn3XymT5i4Ll+St2x
5hUOOPBvpzpHwtojXSt+byCc9HcPFjWVudPiuUIAqWII9UmTqSVTn3LrwZSQ
TvcU+mgAYht1dabTPEiRbTcy/wY+x+wtEELpTAc0+LDevf/CyIvtkaXG/p6G
Ux2mkOBGE4XpXiNB6ASfRR62SyNwIKAS5zajhH1/yDWLvZIqQSE5bpqjB188
OJ7F1iwMqnvxs5ruzL+ozglwZDd1mobNFJfn4gSHr9G2liImZrE7jNRQM216
zCikbw0uIsgzonlQ5ajg6j88XjctSpN2rhI1SZtqBL2u1rT2OQwDhpuzs/cY
1gd2G39pIyoJ2/dXeC9JBd4CJVTdniCuJhjolQImOQxIVJu2TuEBIY2vtvA+
Ywt0hnnAR9ZAudP6TTdaazGfZEUgsvbbYLDS8AEU06HMafTWP8ACRMGpPhe3
0KO4zkrENBFjYv13Y02ffZnXCDvcl1/3wrJPnzuxF7DLRnqRvuL0cb8b46gg
BmbDpF+wYj8r5ZTEA0ttixz0BmhRrZPpdWg38RDOYDXzFty1wn3D/wqGXP/P
GRaddIQjqptJvuZACpKO6oNK4p+FW8Dw2LOujKXYK/ZoPyovBBLHDcLdtgN9
MHdHg45J9DxbhGRCuT4AkvFCe82PcXOcKa7hdUbljlC4z01FdZc+wQQr+IgK
2fdFHx4Iuk55cyREGMDfTsSOES9C7jtSThyz1q5SDVb7L4hTPBq3BfuNLKaZ
Di7rNzej3cHAfR/c/P46QpGQPw1WFZXO7TZKSoD2ULwsubaDFay3gohwADGI
om1qncevGWi7Fw/jP2Sc0jpSuLcCEVxA1unyCXZdiEbeGq9+tzZbPtlX5XdD
iuD85JBcai4Xb3NGrAOcitzqdSCWVAu1p4t7tiNzMxKF8ScOfHaC4E2OzhBG
c8M0LY/wxlStloO/DVJ80RIW2M6WW3UYMm7iRNjWdLR13UEmi38yCKZ1SY0P
z4T9Oat/jWpNIxZomqZ8zDTdy1l0VwohTcI2CZx4aKF1E6HLduTb5NExei7S
qDoYQnVGAYfhScOGK8TMRNiKmg5J7wgXLKl8z6TS0j70+bU36Z0abFG5ndaY
Q1kOzzOgzsLNdnyPVy3JzTdIlSQ57pBSC6+M+jdan3bFZ4p+V9jEgKhWDrFO
sYC6SA3roA/j36mY2XVw3HThtiJlRaj2LS0RUWJ5RctDYV7DzGpvotjnVHc0
tcLy1/BN3rJHWqDyNDAUMBxqiv5zc452lHGW6mjsukxrQXOeUPmlQkRQD4Gy
RqOGOlhmL+rcjAxV32DCme2JgqWxqI83k4/GOMRNexqYu/SMeNKWioyg2mRy
75n9RlwZ7CNmBfricGjkvBCiBh4rm5pXBL8mFRqtdpJdpvRgXc9dqBMvkqWl
UDDQScO7QAvWz2yD4xOGWgYg3DPDiTRzAh0wgcttHHFqhL8i/idIqG8/0dst
89GcfHSG0Vct5hpbXETl7GKA8kfAdsgfJdM7rnix+b1FVVXHLi/+2yXm2V5/
qq17E9BB2NjS80wxvz0UTAq/FG8Cg2vK6tFaNv4IsN4WfoMtMerlOVnjW1lI
1Qzr9lAK2HWw4sLbEZ+lpUZMa/zL3Ar9pFPatoN0L9xtNDYn0CoBA4Ae8gVQ
Y84hOfDMc1zGRKyG9Qp2vPHooHzNk9lPfiaFhkAZDbvwyt5z2+xMMo4egHmM
A0TVXVk1q/FdQFB01yr98+N1/tWRq0OPvNTUUllSP8gCun5a1esIhEukoQUl
GelnB1Z3hhKIon9ukXP8aa9oImce53bGSKipiHyXfnuP5mo0dXbGpqI87qLF
Oneb1KEYxNUreD7BCA4qIi7UvxUvrGA3+zDmEU1Y5Uns0M+b6Kv8TER/FNX3
ta52cW5nV8AHRn8shHXuycx2hnB+G1daH6uOnLtzJ6NVYuezGClJOLbGYfC0
wYcTuWJcOhJ5IiFixr1Cuw/Q+V/tY1Zj8P9Qw80HNbcSWSyLddP4cuMuK16p
Ic9De53mxDeIU7V6Ju7TqovkyP6InQx/WyYd574u6gmdleCOKQ6NtxTlBzwH
6fvRrQgWnIbRL28lKrL1Z9Lar4y9vJ7EUdE20UtLHzT/kgku5hYuUofufRCV
HuH8H8PmGxdsT9GJEe0Web7nW95UP/o0K7T6ZaRLEowJAVKTh63H6rbRpDQ/
qdTW0KRhpXHCCX2267Jzb73AJJkt7xZThAYFWEySMx4CXNJGHqLDTHbMCXVD
VyQlPFAcN7BLY1N193WGEeUcHnEWh9+I6G1tPU5iBPTD8C7fpa01Wuf+DmFz
PQnIkt/xE+xCs1kQPB+4E5olA5E3Nt/d1nawoMvQfo8jqqr629w+IXk1kGUC
if7yoIm91s+zEwT3eQher7QtOAZsBmxw0rcPrhIACv2VDFGqIjTWP1EP715k
wrRTffcsIZS9eL04iKkq01JbBa7EeZ1Pu0ZP0nigmxDlV2fmaPUwb1kFfZrz
RIAXVP0JVCPZNj1Qz3DTvsGpsC7vhL7KPWAuZ4bUhkDAWHOAv+wEkAJ9nAHD
pipheLVvVRsvgZPzsT9VyceHSlBlOTidc/sEEFcTQNp3BI66V903M2/J+zJn
x45fHPx8eb0pTY8JvMSDt7fDER5+VRbPmMxpJDf4BUViHU8terFzGjpkvkTZ
aRLNO7hqe/tJQg2ABktu+/RR+5PxajFMYCn4sgJ376YBErwxlvfjrfI89heq
CJhLkOw9LvUZ/ZbYBteSJ404mn1cdsBkOAxE2Eo3vj3y5NayRlcd1no2JgXY
0f2JzT7aDJ1LGxiFMds3G0s/fFaljiAiJ2lBV2MtZ5p9DptbGwb3gNVfpP5o
emSz3wlvriuL+SMSv+pC4fZY5eLf2/6Hhqd1NWzFDH5ePpzDdPeJJxlaNlu9
34Y0dtgVCUYvQ+GcEqB0oRKcCsfCloBi9bx+BXyMCQ5QXPpeOBGxBInoaKzJ
dcTKSPpcui6VrpnZDHeod1vRhuWhJI5AWk1OFvRVjfar+z4FPpZpKi7z8Yh/
U6LJkWWfDENbAJZWdjWb0hlh7dYISHF325f6YhjPb4dnTXybOtM+ZWA//Wh5
92A782jVcn6A+/WpBd73yQKij+WjpIrMYb+jcwMalfLW4jSSQMCPAj4JNOV/
faG0G/WCSXYdIS1pmHAF2ZWM9sbwV9IvfYhDn0uAikU4mvPQdiKumZ9ckuOR
dzqXdoncTMciCY+wemL0LB/7u91MewsNdimHDDZT5z5KHn7FLCVR4duOc9+C
MBrMq34tVuFsb1y9hvu/Lu8KnRiB9mzUyY1Kb2AhmLevr+ULJcWn9kJ4wxa+
lz+9SGIA2Unnh6szOODwC3+qlIHR8uaJEWWVKoIG3QZ7bEJABDYZBSgWpkDO
cKZ1X/KRdqtBVt1IQOd1q9kQDqlBM3KEDeo0cjj+/ECEAnhs8eSlk6tU+oZ3
Qwl3u/OBt5HdPQBrZZVRy+zlpvaedqZDoXg1Hga0i8HG1UPkEUFuOcc5AEwA
2esqr7uoqeBb+1WAqmL47084AIm6BdLc/rfFua41got2lhc4JACdt5q6mV7i
xXAnyh/JIEVRG+WvCkbiriPLEYCGcWoKIgM+kuN6I4Y4j1GWgP2svM75KU/i
DewaCt2RGhqPrLyGjUQ8Ega0fbUYwKIP7e/ZZ0Bk2i7XnV/gzQH8kDlUOao7
TfjzZ33mUF4BISrUBkd/UppwKnIS+r/AEc2nN1PFzXnq7rwtGvG5LNg0PFzn
HV56GfZE047YM3BlDyCILB4PWlkGZLFHAGyQmcAOAKH/SXTsZ3KlvrlLnIBx
qnbVZ+ZRp5h9KhlH48Kczq4hbZqJscNXxSsAuqG/r9LTC33BqT/GqfKiDzNg
umXiZcj3ShP+rR00ZsnCrxO+COL8hzS+F5rs5uPThb6DUlZ3gikVgneRcHY+
YoFqoFi0l7ruwJhzX4JKL6RF5KFCC3LfH10/NN6mFSsphYM8aTqh+sBy1HlG
9ZEI/8VrruDU4PYw20MMhkDiKEx2fcC8Jo0tfNloklDuCzaRD+pd2k+HrTDe
+Sfnlz1sJRLa7WLbX302RlsHyHZ55wCA6xXgGWNJvVzZfAppIbsHmX33Vbq/
+Hb+k+JCJ+uYzPAqf+3eD05rhMSLibtOSHD1fsy2vQDLM0s4+ZKCM3GyhrDI
imLJRU61wGV5Pf+mMFvAGt3x1tn2CwsHNJOpqBp2PBA5niK4iux6CclP3zhd
NxEXbkUsmf0ONhvIJd2KDNecjUQ8wFLFfWAp5SLeQMKcRT6QZ8BU4iT3+l5E
Dx8rVzgJmFo+hO38f5/d5qmux7xMC5y72RtMyWNDfb9v5sMy68U+EnbJKjS3
s8F6j5MQKOuyvBES1H/ORQc+fp6TlXEM34rZh3rNeTbI2YUJqJAtAfBK/58w
f0/Ov/oYKONjU9xaGZOjpNktGQ/R9XIZ/xQmimSAvTWFBaDfl0aQZ6nsqj3u
f6uB4pDrvFv7a31IQOHjWf756f2qm8jl7l3IzobsaBZatFNx8d4ELZuYYQJy
9/C+lz9aaUL4YDxEch5KAeWmxCZ8/C8fiBOXmRUu7FGz6rkFRrCZAmyoL1Qv
bKtRvdGnIDDh6zUeNg8heaYdTBuAvKA6rvZB00uWE6IcLSI+gBDbRLH4Z4Mf
bXGHZk+kKyyF0nqqb+ufWzlT4EdOTC3lUlVF6Hivjk4SYH2ooDaBonLTnjNi
OPTg3WLobIjEkFVnnw1OVrA+wRBNTyV57XwUfKq6VWFwoU1GG41ZRgvSJhrJ
JZMHhISWTEOQZyDkjxx4PR7XMaqRyNJKkUtHiZpRstTisY1S8+P0BkdcChJj
8HcMP1lSVgLv/IRPUl++rzX2Xd+UtdNqPbk4B1xA9dtBl7U9z04K8TeEq573
dS7OHgXgNO/89rVp4Zo+wBHhlUXsXXqm+tW+a18b7LW0NOd5kXaG92/smP+6
cJjGF+WvFJduimNJ9aARPbbvjonr7ujCT3TB3VKXoEhdQj455YFqnm52TYsi
yJsPPnB78dWTbeMqGTgq4LIvcEUV26K9qq73qZhMEokgW10v0NZOVF2H1mEh
TgdAXbMX+YJzBcmXF5jQ5slvSpLgGLIxI0eLoH8fSrpWjHyEkAA0Ye43GknL
8NMJn20Nt6noM6FfWmfRahuAh9UxjKjJjXZw1BTllxprSEl25UIgbGpni8NV
5mzO3q490IPYpmnl4L2kuyErrUs+0Pw3KvqU7pxY81wK6IUKFZVXXd3HA51N
AnQF7GGUxXTvMJ6g8Xl4a3/BAr73f1MrLxD5Rn7det/llmTePEy/yDRZ8ZdP
M/7XvGXDYuNIZ8tMAaFD39C8KaKyXPF4xTyLomg/3g3ohnA3hjH19NTBdngo
XatHDItkl/kv49PPTUN6b1OlIPYUfM7vp7x6ponsnbXayJ89v2NBuRrbk3RR
BbDr42SkYRL98AtjHn3MlO0KgNIn4UfcFC45A0Ek7fS5NVykwZG0clmnO2kI
V9BflxtB6wb0t5Fd3OKDsBhoqUCv2mRF0ZAVqJStxyzynQ6RAoOupyvuaCqX
lZbDegaf9qk799rHFtkatNuiJBcCriGon3zDwGcbBnGnRQMtVRIlehBEpvRK
xtrlEKSnP68EDeEQg0M+iLYg6vUph5iF5cVxbG2isKELzbHgUJXtziHNnJeb
Q80OvxZ173tfpGkXEyn8krKE0ILJjLU3CoyJJ3mTSBJQE/kiJt08+fO96ufQ
Z2d9bWNg2kMTyz1/658fdP2sDHwj6VYNatn6LBUggBS0/U0VTxcbPJ2Xc9DQ
YN7f1Zowg6PDPLUHmgKXZHoRDiUjy3BSQ1/Hz9wGKclMLABuk1TDf1fzhOxB
5OqXuFp271mk8I+SMzIx9ROY1FSoFMXlY59y9CWJ6zXTJxVDaqzn3RO9wLBf
vEvWWdo53zlBNVRhDIZGGdiKHBgKFdzhp405TtD5H7ajRrPvRI7Qpp5aXvbk
h2thZRlO0RnSsoCyzMto5SpHeZ0Ezt5qIqBjZn+AMVEL5j4+FbSUoh0y1La8
TxskY+6jpuqGgEQ/b9SiR+duRGBZH4WwQRBONqT3YP1fx8YcqSj7riplrMtO
BrJEtB7Pe94ecbW681Ta/7yiLigUfXt+YJwNV/iSlGvPqkc/y3QxL+jJ+KRE
4ZfJSxSDs67B5PAeF5kVLRK+We+LDbkbRaOz1XT/0qnaVGEZyrJ3113cWJWK
nMH2YY1GVUgjiOiGejwjBl0NILIMk1f4j6jn6DZ36YQXgRrDIU8g33J8Qo8C
0luSEFAaZsWMAKawKCgqL+vyN1ulozA3Rl4aZH6pael65aL7dF5eJ7aeC32F
hpLfT5+FQnb/WsKnN3jtJEdGtxJoUNEmZ54Qaj/Yjf7LfxbWBRlNyq0DYh/Z
3aBWPEDZKEwZCAXL7H8M+mqUfC8j3Rr0NTWh9IgVbB49mGoptALQvyIxxbGN
FB/s6bYqSQtCbMZGKE/1VYZEct0IoaBG4/uq1XSKWJIjsGkj/z5OdHId+QY8
L34bektkMvR8ndjj96WcPJGOKhJB64II3TedaXzTr3qCcWmnXw3ptIvgAfQb
qlhu/Ceub270a94z8JmhAifoIlk2iVwejfwx1yaawY0bdydEqmVBcHZzI5zO
bbgSSUbqgPH2GOLhMEJksk1PwD2odGyiD3v0FF/6C4TmWNyMGkmZGp35Ri4A
7v7nL7FEB2alZM7QUllqEU0c61v5xO7FY02jCemuld8Bo4/XrDfBs4i4fVkE
HnZxoVwVMj9cHvcekLYkIvTS6buxniKmqja/w/kBgI5gGlKoGNEmz05bIMrE
e+Da8pIAligvM/FJnl3Uy67bZjyICiV5dnY85M4bJClPL9iWKgeGM4jLtUGi
MOoFUFfIPN2hoCj8cbKJt+6dvyDd/K5xKP2EyeLWDIC+V9XCDz1VOwfI/N32
4X7YVwuGa0CJTIBWlSEAz5+JBfDzUnhinBuEMGpBVg7aWJoaZ6li5kQPlVzF
OwVWRwGA+wRsTLAPTlwIilwxpyDmPM05a1JAkSleh2iTMtJYhFu5SgcsIFK0
29jn/2kpBM57xGAOREdLvHtbf4WqXpnErZG06LxoyMzt3mrGIJuV5E2FOOv0
Fm69A12w0tlHW/cb57PExU1H2jAYOQBxIXX5aWwxoUlXcRgrMsXZVjdAVZqI
d9ZBo5jw/yUYYPhc/h6k4cH5/VLpSCCg6VKlw2gKiycYJgsrbrHqrLqrKwkf
d9yOHBI9P7hJsjQ8VvGHYxSzp62P4o21shytBFBfQ4Nzsnau8N/gpARCZ0O7
xz/OUoO0Nwp1vnzWfr7hZijKprcKWjczy4Bf3OlKzVilQ51Ii3+VCWRaZaX2
BM5VtBcFd4I/zg4SRrs6dSfls3R1JULmeNDzZilWvkivNJT53VoK9g7K4DbV
mDuW0kYuFSYYxqUarSfgU9pvqaCp1phdd3yS9QuoLgRTqF/qQMdRq48G9JQj
eG1odgqh+V4gr/XcPPpf3d3pAwrfCptrVjD8o8tduOBEYztPSox4Rhsn5BFM
4N19mi/ZGi6ih6eFXIexof6bu5NLkrgF9yh0PfnbMfOIuaKXPsASyRfSc4jW
Hbph6hRSs3340FJvbc2LCex1uSB9diNUzc6OA7F0AzPAOD4ElAGJJYHu83N1
JlndhVoSUf2r3QWW/lQo34yDtfVIuF407jBShWHl1iHHsekuAW+sKqdv+KkE
tVhWu+LFa9jvQGDaPqH6qVLclcZefTRKsWWsasffRheaNqyMv2pjQpshXN6R
cGE8JNiKs/1uEqEM7NpEhGlAUugDLaco3wAWZSdH/oiQuGccc+z7cOd8Nhbv
Ej8xfxQxcfufKviNj21ECVs4McFIIcg6Xp6RgskPTaduTuexhJEch/xP28UL
ZBhmBVIjJOhknn3vbjtfAFl7hFU5GJzw5ritYKcemfzb7MTzh7ZgeAFaFbYS
u6IMLyp8Y4nmoDTaXZxCHlE/3Og3bo3AGZGpCWmcKCSrs70RLj+FDAjE9Sdi
4AJZ5CKAUa3uAg7Lxk0jYji78Yb12GgzV9yVKxJ++uyWgDP/zra0KfbKu0EN
M10fqPV6Uoj8ilLS0mBs6X/UU1LpubptWhWb/5C1opgCyDT0TMrJQFwc89Np
YFRoMojYgQyTl5JqDmZ1WzH6cmarDW5s53VcFxNPOFU6wORt+JKWc99GhLc0
ywzKGHdNwnBO0wi/nGYaPgdi2tR56K4avuZMYgCcriHvTpw9MzgYWkm7RcC1
5q5KZYP14yz+YDbO1NqSzIW7D3rDX3FC3Rumc8EpEart+u974dhgYolTIBVU
pmfxsIi5g0zwqLMjrP7CFraOUeDfRUrrZeG97QrP10U0fTRJqSF95TjBZ2Q9
iV3ekPH/EX2/F8BjBJ+otnqgM+fHGQST1KM3SF6kp5K7Gxc3NJF8/IYRNTsy
DYwrPDW9AGD3Wp9+JSv1IO5grcptk71nrU9035ezD9r02tX3aGpK0ha1JFbz
7L9N9NW7NkojMyliEO9E1+D2X52DGUDzDRHpGDXj2kG9FRh/nNs4tBxKhcmC
V2ONmvA3vgWd726KfU7Dw2Uuns/vk4S5ZsE8yBMt1CXKelTcBL4v/vEugVHo
JgPleiFf3clkvcFoyJuIKAqqLEjA+R4xH+cUt9FLAJ6HeFpjNqbsUYI3MjPv
er8p/NrRdfX/IB01QsYqszcrVhz6JS/ilDiTcS8GyzvwLKgwlAqP154ZjKLs
D6EY87/KVP/0gUq2tYh08Ln1PBoDWxF9YF2ycykXc5GEl3Nuwa1pj8LB4sC2
clh6p8Ha2+9EU4LHifKL+faZm3GXNgnOeHyE18Usl3MroGW8G2+DLYORux6S
EGNNo5xDZs4o+GbSUanQ1Y1I4D1ZsRj2EXRSSGB8wyyByAvD1Mcj1RJNjbpS
UdPaFqRDPIOxHNBVeKxQ51SnxCpQSAJkEFMCfwaf6qBiLtQjuzizNLji6Jcq
MyMjp9CiElwn8PcLz7QBoI8UHvNmqGK1r8iQj3MglPGfZvqui+Q6vKvqiNWp
zSUZtNt64gWSTXbi45tPfD+W4RPO2xu/pFaEcNJayjxQYrr8Yl8a9E+1c0Lc
3CUYsfMuKqJikkD4WryylCws3XbeKA7mqPVyFmjgIMAW+TrbVqx2HX0ewyri
z3Acdsgf/pa6yzuJ0A/TVMBsNV2/szwon3Y4Sc9SLTPYz7qlYN6O+gkf4FNK
PcIyv1Ykn14HXzyBLpeeI4eeQD2g8ekc/DZTdBtMSJfR7q0lHRrwmULpcbXj
sKtII96LocolI2N4DyRnKQNYGyICwgOkTeP3lOeM3y/p5Pa2tQ4UxWN8xbfY
lrT7613AnXtUzbUQOomWJmm+tFFm65aRsuKATd99iq9Q8h4IlwcF0QHPdCz2
igZE+wptVRVsF521oV0ZsuVvps/wstTo7zwzz9m8S3PRrzvHY05vzKDUI4x1
uoBXm2DlmVsq24yDQ4/+LsZxAiMpY90D4jgafmzRPb8CY9hZS/mIpp0DrXa6
X2bgVg2WP6/KAuXUs+ibsQm5Q88BckZZKRYwu24Fpgkcf9hZL+NsuVbzYpWn
hBf2pBCVTyjFIVWxf9RoBZMnPPsApCwxGClnAvIZ0R4G5/qY4SNj5fiKNbR/
W6sRd8bpG3QNlTmyhahztYPIapYKTs7XZAlH/4NukkCf8xZMRHiiz/Tvz9V5
YwE13nzYqNZv/OWCSibI9ZQ1mRbGHvU8A+D1tYHlgDntaKW2lbw1XMNSqHAQ
nHnIv3/syGqa/8vt0ZozXwPUGWajixXkv0Lq7uZesZGy50KagiEOIXkT9NUA
U/ifhLGx9zihKFAM1WumMwCUhZqqPwxD5kW0mWysnYrDtBMILjNJngQ1zvA3
oUgdamqHoF+/DKzxzzKqcqcxLAvERVUJ2ijOV7hL3elEEq7iZPLJ5l0af6ED
f3Xo5+Y5f0pM8PYAYZyhVQ/EQgJmNi4gP84UanLHepDEmAyiQIqTMqYOJYZ0
IgZ3452yCAVMQRwx+c1SOKNWryQy9yV8wMhEzlkw7gxwY2nl2Vcnrf9bTe4E
tqwxV5vyQcx1015tuF9c3gSbtQ8CcoLTxWxhoz/YDmgxnkKraNXKyZwLDnPR
n/qZbmBs3ZLpbIB8D631GPTjLccCgXrIUKB1Frq1Geb5nrwm1NC9wOZTa/8S
2V96h4DQIkI7wfYmzXYSdfUsbZlA4B+pgkhmf6O1H8P81Ual8zpS45o+68lw
nxv4osMnJs8Bc7Qk2eNb+uugKUTmfe7pf1W7XB/S7YtziFm/DTq7NtaCeBym
8YcTQA+P0c36HUl5I8ZZSCY2pmHgRSjJm1PY/WMozeRyAvo7fvUQ9thCZsBr
HGrbgavbCJBbvEmElmtYWD8BmSWiFyL8Pbqfb0//FZ7SMDKhOZ9P82HOW255
WNdiRFIvmZQf+Bndp1UNimEEK9ATC/CeS4kvznOpczrPL452WuAi4DN3ffat
pPkNIOYGhxJhzvgBwjQd3LohoVW3UvhXSGw6s6CVKK25A4DY2QpnZdm1LVZP
0mjo1l9VpY6yKmuQ48W3l7H51cMxSEhc+r7BYbzHAiU77V/Fa4BxISt+Mb6S
+fBJwELT1MVgRRpGlXej723jxbdtVzZsFycqE0AxXUQtwtbngBZJk6+UpPB6
/hiyZN7rFbm761FpHr+OuyymdiYmakSvwbcIFRcFBXkhi6FoC8VkJE4EOg5r
2aatZWg+Dl399C7J2XPlTzTL0DoV2JhXOEHzlteZYDrNotkwLvybzaRgXoUH
+SzwuwXGBD/WeumqTIBgEa2R6W6+SPWIcRhOs3lXLU9paFhPhQ1jbRyWdsOa
5jWvFrd2CcqYXxqk8A+ej8lDqbRLqEu/sIOMy2YChfhLHa2jlKtPCu7vnThw
7Y0Go2uFgZG+5CEy8FTSob/3NUe9s5VBZ1hjkL8xPs8JISdES9h73ZGGzD/y
tIXWGpEaFsjZV+8bte1LFKsakahiNgE+9T7DIgr9BBRtn3UwlcqrIipvXw0X
nweSh4yxf1cPwli6ZO/lJzS96ZJjKny6ftDWZqZ58E5xE7jrWys4iIahKDdO
5xUATYuC1mJtKzoINIzLkx/8ZkXYhfABODmw1u76vsXH9RjFshPcMD8bWJ2r
bDciextH/o0Sd3R4Q7/Hfs2mGHUPSo+SiJKF9pmVYWQxndl7kN3A0E1Xpude
GsxMeEnycFG8SvVx8bHxlLpoRSmS4/gnUcFOtcF8ExX1FMlNGTWfb7uVIhNx
V9ftqOtOBQ16A2wcX0wMCXB2yJB/qO/7iG4ngCdguR8hDuWrB8U8ybD/rn2z
Yn/seP3ub6hFrFcARUxgc3iWOoF7Cf5tux5uB1gUh2s40m0ikRgIBVzOvm8l
eZJDp2oNAqDHl6iDNrtn0epw9+aTIQRgUZTjPyOFBwgeTf7J9lCLtn/eU6Sq
Zza3uXgO74i5DQlp+x8hGmp/PGfI0G4rate9XR/+u6HmQK1P132wKgv1XJNk
rkZvIcPNqn79ixsrpvdAazXxA00CGgTHFd2JTbavW6GVhtpY0Yzu7tlJ/ptF
cA6LoheQJcItpV/SwcisgvaNskl3NL8W842XwY4RFkip0Dv5uZF9JU3O/qBa
dHeJudENlSXtDRgRDhUB3SbMq72pWmSW9RRbHDpx6jlv9cLZGgehPhV3W23S
+z1OzTp0GmSAdPBYW8/BuFW61mBqGY2F3InBmKNJvjY5MfXszVhiPMj7ryek
DSCczh7CoNX1qlysA5g8xng9kgN+Dj9plBNyahgzhMHl/u/9BeQ8y0r2WY+y
YyQHAWU0VlNGLVRYBhAR41vfu96J/suIHxhTVkivPwxh6Zs1P0LavEsEyTBU
PbL3/rDvw0DP7yZEobL0cK2E24CdI7sEe9K7Plb/ju3b3l9vvGCxt1SJmQYx
7nX8rHQw/0/x0dWwUpyiuOV7s6o1XjjPuhlkPZE/NT987j9wedPeE4Yg8vNb
DdeVn5b5yVmmpgju5h3nK9ZDT2rdlmJ6o+kUU9fEhWC+W1W+dcZ6S/8GN3lk
oF/ILyrKMUuL9GHPqxEDwzYw1gsaqbFBI5cr8xsIfUaOHihUq+KlXze22r09
U/uyYxlWW7i0y8vRkA3gqG5mswgEmkqnX2pTUnun/DjmqmLJF7bi87FHi8Q6
35yu6JErdhs15obp9ZkMpTrGsgP2/AbSnvbWHh7mHnfJWPxGCMyzdyhb/aCo
bp0nleZxhuuz3JfSx7u4ePwsje8reFU5d3vz656q9S/nEPacJQy/IyZCbrUH
2IvajMpOshUFvVFa2nyuGTDujAWR+JSMiQUQvLOSx6RlA799Ipofmm3x2X5x
vzM7MYdSbtuXHuWKN/2rUY8n7oDjueJpv2TMW1GF0u9ANgZwpZkjlXQUFRHw
nYaC7LwnFvYb/60aKuZlM8uOcKbnhgaFdhPIC7+UOi4DKilIu3XHK/wkjxfN
R+T+Oth7q/6hnIEIrXpQ8TjrexFgYDXcBPNZ01oFChzrQ+VKyxIZRe+ROwmq
AfA0Vj8Vt6G0juX7zC/uinmE2JUQ3R6fZx1Z8Mfc6bw/Omc4czZh6RUTEZA5
uThf6ogCiwcpJaUe8ZbJ5SQtr3tfqXr0yd9qYYK7tqFfUYyjS+PC8hzdZ+55
fH5ftHCFZ/W+1NmtgfMWdLRu8hXxrsdwuQ+LEZannwu8NjazPLPCr31k1wFz
N52ujE5oxm+2PD1okyzN0RHHtZGMPNTVszQ3nx8zGc/pRKucCtle/c3fKq6n
Ye2uANJBgFdBSwKMDLwGtGJnrcw3OOlYuVAvDtJ0/8idnRMhjgJod0ACucj/
qvZZ8Y6rMcBAGz0gYh4OQByLTM2ZCI6kjDu6M2nb7xPTjfjeSd2Q8VGRaakF
0a8wSvMjVclidVJK8w74WmMi20Nw2v8ymzw+gWa5MUtl4j6Tzq6vGPTiEKVk
zm8IN1i4EVNlqdHxqAr4k2K/haF2zGfdjrbiJI8wRAA/BOxppEIqVmsdHokE
vKHbmD2nid8IvW3gGnj86vebBtIEGU55EPSjrWwkmk9wLY40vafN6jGMz1q0
EDnem3LqmnbaSniprIMXltGetm4h6UPbT+55VJVYFVu5DdX8zDaGGMoVqRHx
DclB3lt6g8KIXWYKP3i9fCLni3rY2B0QMbF0NucViyZuOZE3gSo18I2dKB92
ZodhTvlJ1i0dbn+mkUu4gVUBbp3BppJNbwWXjXASK14p/GQ++vlQ9PsYvv25
vJ2c/LA4brF+x2bEDi4m9QIRDGyLrP5AFmZr3fQKJ7HfYDMDbLNGwJUslK4H
ZLhmP5dg28iPeJFoHjZA634K1DAcgYHEZNJT225pTqmvpZ/C7XVLpr69GIKL
UhJ4jByvuzpNL69dhc/3gKDVXSPNnBwnEumPNux8rcCOoAuvye9PkN62W//T
AtuSTTwYhcuo1Hvpc6344jSjtPJrvbp8Ykul8VuzpTsl1TzuQozYWYZ4v71P
122zGn8bMmtgngSfzdxkduWGVRdXbX+utKDOjYgw7ABOyctvE/X7tX1u4KtV
FvxndeM8UyP8hJf0c+as+xMWDbhzlbqHyEVD3Ue9U97YuJTTUUoh1XdiCEmn
2X5bVvCXxudD4JwQTO7w+fpdBY8rxntzMmUWLknft62QgntGZniLs2HsH8Xv
g56/XzzueV4FL5A5IrDlELrptfAnxMpiSHMv33FZL6gkkTh0i+c7UgS9wmKs
/DiOY5O2mzelfSePkZ8YCltqkjOEKrfpT/dRkSbatYkH7tbaHrKKfS+xpTkI
64Jo4fx7207zI9U6XdXFSaBRcHn6xtxlzyzIwkZUMYaAbUYTakrZDSSQb8Qb
IfD2j2FDdXNKlEpir04YhzUlRee/aQGXSQWMsPS3N7LCBBLSbtJcpXA/RVlx
ON7lEAtsVP1wU4V4t1i2oLaOH5uHZ4jSGhYxD0mJ1ftps4okdyPj9ayvEhYm
5QD/iBDqjQ/GFeYxylOKcuSZVtPGO2J1EJlyV8oOaqSrtTRbvB5fHliW4grc
tIS2Yt53gOyA1AKeC5twThtdoCASWCYb5OT2535Aud6ez7oFYgaA3VyqFB3z
EqNRHyid9PehiymtlEIw/6Sis1gCOLmaha4Ij9TbCBuDCMAdf6wy5Aeedm0s
VisO9mzDVm8spsE7S6peKJUrN/4OO/PoV59WxiHgIGCv6rTx5g2cpEQ2fvxU
Se0ljJi/5IIjGkz5xAxvDvhdBPOYigOjm1DYrPR9O/NPkYirG07RQ47OHcdh
GRVAKhr3tZuW0KpcFZMxLXZ+1rxt6JIaXbUI3gvMNPdbIRoMTdq4IWOrF/34
noz3UadWYh/SH6nhIWWdU639NPJpUxdyVgKMQsX8JaE3ISDjFUPeBZL1qq6W
UKJ5zmczLOCAorstcru3UW6KiFFTxU9Ym0BaYdJX9uJRLzHCtVgwmD0CJOjf
0SB/ZAe0T1DJv+KAyRjybdQKirdY1lv5ZR5nPCHygqQffz8UYrrrSiFMHgug
TE/bxCN1tDh1NJjGKeOSRPf2Mtb+cnQo5N55d/0IzRf3BcEEW9MVRioU8pdI
O5dCUE350GalK++vsqKdthS8EsggMhJyZHHBJYb7aglG4aTtzphM0nMr+xHN
O6nWnEGx9J/qd52eb5OTJE5yzAebtqW/4mx3TVBKvfBIWyM1cz/BQBgkFSaw
DyEkg+gC9oxhBeZ3yjhpMxad6WvunpHaL41jzfJnazZwVXgVXsDRvkfjtT/v
oodauIUxSEKsjaMGLJH/FQmQ+ax7xs8zybUrMJ+wRtS93UZ8rzwl/IlH4xK0
4gxxh0IPpb5oJD0oN36AaTgS5Uc8cAMOfNk+1Q/iZM9vPmvQjWriS0UEKmT1
eor6aFDdXxW7USjX55trsVdqq3Z/YQqQMP4OMHQ1XHqHQRU11Zv2IDCT8jqH
6Igtj3V5JdTsiyA4P6bw02vSf5o8GEXoC6Ag+m3jt0fzGC87JouIDjUWAUM9
8O8Iex2TQkesD7shNQEQhpWJk26h8DFQm5h4CtWCfWbfxM2KN+PQKy01gsUL
pKkuxz4aPfemt7IxMujXCnjNLpAcRgXhSATJlk26SwOBmgfZDivCu/gd65vv
CK6RZeoJMw5X3eSwELGrk+o4ER6EY1xLHRHSXtYmrEMu/EU4yIrdpnS5PODk
mnL+vEhSrCMwdIL/QoKqioLcGhrbMBjQyCcZ/CTSgPgDltWkY2AkOTsCCjfS
LS/UBWRifLD5+RyFQLhz5fbzoVXVAghT6PTCN8E5ungz9GH3aZE9n4epLUFF
vOLuBNZa0+6ypMxh7f8NPf+v6+qlrb4mXxbpLAsrQZ4w+fN7QMPAR3Fpa6gu
KDsJToUP9cGGh8wGE0bXBbd0dKR4mdLLins58BoZ639+Bg3FZFSeOX/nQm/Q
dh10q5wrO7HJB7uD00K6jFeaa+ELcAkVlR/Sn28WDFxb0v51Yx0V1UTDRkPu
ZWBwgJOti+/o6Xg+ec0x13B7x6fBAnnqbuZPx7YjbOAorurHs9lm2EH69Gsi
bCIJ+MAh6jaXOERjuqFRcU9qwx+6eSnr4S377Dz+PVMiEALBcl73cMKbgMiB
pN2U21nU6VxZbw8Qhc8lEY1fBycnNLCktnenYwuKALRdtQauTv+xCkbu1v0P
hkfHGde8Nc/WfpNek78RN99lWNFoL463sgwGqWOt29UeXJXeqBjhNSMz+d6x
h5+UkMiStsqL0D1iMdYm26DfJQDf3CiObDK1e0KGY0/pj3EMl75i+meYRrjQ
ZB/JNnuXu3AXyO0FUbvas6+ZvYHXUornA27CNn/GztFDkpHRGU0R5VQszvu0
Ap3uV8nRLrSspXjKcb0jRl4XC4bN2p1FY8pUV7jPzoIjqP58L+m8qKot+EWQ
wbohOQ+d4/Sn+KNSXa62R+OiQgCuq7RutcGxmWquj4Wkxu5odEvQlC4dUk8t
i/vq4NkbuGyBuUOZOIQLI3UeSXJdZZvZTwMQ4m1sjlAkDcUJEvpHDeSL7PFz
BON65Fu9zUmrFUcWNfuNNOKVl8S1jiiwQndn+5Je4P2Bi+P6/KqRYOQZ/oqR
ZUZagttLFgpB4OxERfcfn9ritqDPRaSJG1ZMcnAf8/SeeP7juer3QF9A0YOt
WE3Hz59HecOSc/I03IzITDhmHE8jYvKdg5avHVttvOLgTGcLZD2wDvlvZma5
QRJ1uQWYSH41L0kX5I912vh/ZUUvjGpmGe7TQHkkkUvIuMsWVqkp4DutnlJp
BPFuA2BVHCO1x3EARkIyuCQeccWnnsj4O0gySFKY2K/QtAq54tFKVaaB38LU
kcXvpDNG5Y0coBRxW6cFtm3BT9mYG0ZyIeF3RyaZW6WaaritX0IYl9YlYiCt
gJKJzGZMQddRCUuxp92EkttTtSzlIUNTNTzvT01aX6Yo21POXd4hbmQ0bwZD
NhTRRRZzlzM5GpidnFwOFEKrPykWX1FtJFLd1jLVLGJigI2qj7oXO79K9j3C
JhweH7FnHj9kkQdj6vYvdkBEVTHgffVOhKTnyM2Ukt3lUVnv3/kB+aarftuX
oEFiliFzwVcvTtvr6/nh5CqEjDReXllVTVO6cdLMksiNLh7y+WUcsHrwvdwh
8BUXZBPpdlDYzBgcK0j4rqp53/3ZQNaG8ZuzfQ2oqlw+T9/+5d5h4/7WcpLF
rz+HBnY2eOrqAdfAw1Kkk/ci9jK46fZs0c3VizsGEnXAX7+h8NlmmOJ7p+uT
+My9QZo/R3Iv3lEDismVmU1Y46rwFtg0P2X7Xfw3PX8PNEsGPrFytdN7cq2s
i58gAb2/9N2YC4espuuWUjqqm5qp8i+O+HhVMAK02p5CsQRsXZpI3N4rJdKk
00cJOL8rFvq8uKBiYiw9eY7GYA0j/9FjHIoKvDEVng40gj5joxubfeOvGnsl
/CBPIBhlBv2sbAT9E3gpv6eyTg2WLA2WnEzSbTFGxP6HET0nQZammS4iXDLx
X17JIP6SABBv90edW0yDgnJ5rWns73EC5RGzTzLgiCpZ8zGt9+I0vM03XQr3
z6MM0EszFC5feuzx2BRVJkIHdWakz1XEmEOWFFMjpweBTjoaI7W8Tbv9mGUk
3pJMGkalAQmmXmATZuakGbiQvMecqKdYGwuLbcBjRrNq/iiBOUO6D+a9dEfu
GL3k+P4hKeLWVjYsFSZhd1f+XxQly7GoHG9Qr9rKDMRaBpXyozewGpbUZJiA
+GbMJrgZY4yn1oQ6IpmjbIe/IuojfvoNnd4AAGdzHf47VLkF7x6U5gP1VKgb
79JD1INBS6hJzPLYjwZc2WHPGBillEo2mXHH5ieio309BjlAB+fpwXK0UWEE
jo1u4nA2dvtgTQJ+0YCYAvGUe2SgXRXr/hGZ75yDeW8YvRDqHqGvLyB+Nv41
cc1xrx0b+NJXf3QQQ3tynQ8rGDclDqe983GeXZ2u+r9A5wGWRsqLR/z17lKK
VrlGKvAM+X2Kv+MBDCCZWAbsg0zW2emBkJsAVESZGnygstfUjQCTQVMDqFFH
Ve+fwVxqKUO0ABTdT51XBWBNIztVaymhRBDyM/MOEKL0tx4z79m7yKOxrsj7
sADVgjPB9fQpv9BZpw83boIibSX/xKzihBIMi7BXzOAZVyb5OY+0FUUmdLP9
bPm51/2KKST0ys7J8Qwruk0j4I4RkW34AfNmbXRjSit2yASceQ3AkYz7SpKI
jEzUDA4fseHk481HJhdpkz/ycGEDL0U2GtBvT2JpF/igD/UNEdt4moovgrye
D5u8jN6pNV4xV38iZTQGfNFLPyqcrdFzqEBOjgdpUTQGqDLWbYkiavLtM9PL
Fqz80XTvLSkRFPt+vaUkDtyCObNyN+hhB3GtlynW7sG6Hihb+/D1LrNsuYYw
DBg/6F4esl4WT/2eiGMT2xQe++orMW2rEe3r7xozpCdQFH7JwUCflK5pWWtP
nrwaI7lNtP0HjPjUbJmUtUrR/hd93DtHjYU6eDkQRebAYKCCcNfnRc0fDurX
Ww/WHaem2tuGYyCcaScDO5zUXLzBoMs8dG/UE5q2nOuksZXGkpmKWT/MurCj
BjmPgdRjt89H2bQoGwPfVAJqL6z2p2f5oxlEmwZ0jjMMXXRp3BLtOIzN9kV3
xiNbF3KNcwNE3epC/isxgWtfi9EWMasV4V+cV6O7F/TsWxsjInEBjz7g7M1r
tOjyheZV2/+d805K/sTef06nQzSLzalilizvm25knAr61EqoEPv+D9EI+PwM
On2krFgS2M+OkkSTt5dl7cGrtMPOk+zo4Kd9WQMAaXW1Q7bQMnL8Rh0ZL927
iItXyRmkIDmGEKdWoCWNO+Izeqzz1rkQQc65qWcPfeoIKPYmRGLs6YTupgnt
c9EFfGE9poBORClxN8wKikdx+LNUnYxqcPWGhDs+o6q9ekQaxpV2XwINkj25
+Yad6Q5lrq/rKKvwS0buhTvCLF8loDF5L7jvmrcVPo3+C9fh0x6Az1c/SeCD
Y8wdqAQGJcmKI0ylUgXBjLvrlZjmVP/YLN5ceRIaaMkv6qRJNr782b8O0YqW
mlYorZMZ/XAAf1O6E3kHt4Tmy3X9e0M8a0NZGZ1YMsZ++oUxL9eRAHZbDx0T
ir4qYmnB95ivoN2Q7yu1vBkEMvGYQ5Zm16S+otELKZsJ6IWZ71jGOWn0giTE
lwIAjzd2zqae1DKjKXZYBpFFgnM8gf/x6fapxN9wIr7WX9rvHJBqyBQeHrnu
irZT+th1IcJE5mFCK/epM15QtODVjIQJb3rigmouzkN8vv0XsBgNV5PTesK0
dg5FWkMO1TCphh2K9IYe1Zc5wzZvfu+81XngR1HfC40xZ9WToVm26IzasQI4
DqnafOJVcv12PlGS/ZhXglCtkMUxiHre95npW9KEu9BjVzeHjfCvSas7Bixp
DSb6WpSvElgYYO0qZni450DhvyK8pkjEk+idu2blgYeWTOaQY1xKSGX3L6sj
ZsaPMTWKVi95+V+v9gmmSGuwrcfiTmavXzBYvF61C5906hAwNJo0cbI6ZPMw
Qrm8chdJggDTmSqWgaVVeAGIcJo3IvRlrJ453mvLh7imIjFEkjaBXVCxGE+f
uRPJNDb8FJTxVFG+EExIXwARMec1kDiTj/91O7IgyywYw9yNvKFDWbk53YSS
3KLlJKgy9FxSJO0TXoq927p8gynqrfwezCQQ2tu0xZkG1/A93hShBD/vzpKv
0zOByHLBnX0Qm8wYuPpHQ5XQjCx8whhVoTeUY9vbSL4scIUG4uyrJnCIjlYB
r5z++Nu6Y4VgKNZaGCanJc+bysMJC44YgPmQNDEFpxLKfJlyoUlrM6YBp6ai
ykDYH52k2asUMDQiWs5ugE8FE4RrD29VzmOtAvX96g0eLupMRlNj6CNq4NFF
MvVOU1RRYkIUj4j3J/dTxaBFAjn2zdQL3/z5o2TriknVE6KXLAKZn6EPzLWX
QSjDRPKcFbMN3Q1gJLF0t8/mNvwAsUvRWpQvDf6hMoHVXvrQ2tk0JyirOqQb
BjhLOjgYlkCVp664G4R+p6w41nNuiFjlAy8KsJDufGhR3SN09bOtI3jFwIEh
96mtKVZpBqZELQ54wlT5ZY3McirrFDVw+WjBA6lhK1lx4KsGMzqXHyxtCVND
pzTW+plBHFC5kLAxvOQ6vFTMENiHCUvs9wDOakey+N9gzzpk3vMVTa9aZ8Yo
WE5P7uC5P4MOQrlqAeKT0ABmpC4EP2ejYnLLy8UlA2pvaVn3OW31v91QaGOv
whV1yPSKFuOkqBO9qsKEPGYw7cnMGnHe6Z3BgG1y4XOHHtfI1iUvdnDxaIGc
rfaPSxXerVgVDsca2ZtOBr+1uPI9SJkyYRrbLnNAAv9z9ePqh+mU8uiyEGf2
1RqB/bfnEnrJZHHkzXoYnAB9cd1t3Eic5Tonjqne4A+e6ejvm9nc12my0y79
U3TLP5C4vKjSVQxgFmSu8tGP7BlZqn0SuKtlDoeCehN9ajFyJmF9EKqDKS0w
QNnG7ZfgNHR43OFYxmKPEPVqftrA8RnyjBkFLVgaS5uauZqIzHTUCt31ksyy
ccJkdPztuyYNPNThJfdAkgPr58ceCd1hIY1X3U7lcKfp78K+mWUXDESg8sfl
2eZECb4uNQDClP3RqRJYsMxf/yarMpM7tc+FnUfy7zRld28BbMEt41GUqBvj
e3oy3MWqUco9kgJCUX4nwmOBrQfrX8iZvg6rsJrATqkl99Eg+Ok5HTz9tuG/
ALZluMNi8PnkRqmB50e54ARu0SNGbqqJMTnJ4YzaAorN/ZlRwUj5/Hzh/vaq
j9wEKtBonXK0jUC1mUXcXSz1UamLRp+ucU5qXsQA0cMJIN4mm0JoGtDUDe3q
K7C9LHd8m6CGJKbwhtLEHCHwBGKjwtfbj+HgMegIUAcgLu+1JBqGv5DROm5+
KI6iK3LpQROF9H6st/WeTU1CAG3QZUzHHKRCRlk0SOxpreDSKuY/F+wtSX+Y
eJvmuJlv9yRAMfO35O+S3OCiX5bP/wdKIIbwp/Ou1JWGyE327nrK1jTp09sR
fqx4CDahChWUvqcIq26pzk960Am3fReT6c/uXrUrfmphCgwS0FSsUkcaLvBA
1MYIi72D2LdMPsBBQgzcSJImUgTCDKa4IZY8EQte0QKE10QUZk5jYoUgH6Fz
jWaftp5B04l/GUCzFg7LmCVx+EpllE0fvtKxZQQm4FRuDaZkURN8k+aQex5G
xw7T851Kc7t67XrR7xNczyV8p/T57NZy0A2o+hn3JAQa49BC/qT5YWgRUa4z
b/f8YQ4ysJ8zwMIEezVd6eLf188/y7ztKZYH0X1NAFjzjP3OKujh5ZD+HkXH
PP8xVn43oot6BzT6ygECditgRJ0JfwzTbTckN38DlznBdIS6Tayy2gJ9Vbcc
ujqx9AxRq/5t4ERf3oDWrmeqlCLXMg0GckF9CKt3UY1rXa797wifEvaMMMAb
PZO93Z01QRlhO8JAHIvNvK4WG3cnLxuAi6InUgXSI3IM23OjYh6FNJ3uKZ3O
LyFnbKnTY2pfNmlKeOJwGj9Rt9+f/nS3n4QFCkBcQ0nz5du2oV4PAZmuPQbS
fWrhxq5fKzBXPiXktie9ilXCFGTJz7WiTuS8JRNTonADX6g4y3zlu77vj0GA
V9JUipV2G9izKpPdMJB1+K+i3Yt3k8/7oFcX1RR7+cLJXh3l297WW3kFXv8t
UymALYWIgnv/0jY0++3VXbDPoSM784bCyDSINEtR1+NC5x1RGnTpzn+k2NaT
2SpuN6ClBiO5I9GjtwYslGP4TPBDV4Ts1mMP8rc1t//vxfBZeXpMl+2eFJaJ
vTc76iGYn737phK5x2ipJpzEieSFfbDjB4ngNR5bAmlC79dEgtUsXqOn/YiI
35Ovgy09x5VRk5sDv7GAWkfREJIc1Pj8qLkhkRzzqgMq40k5gqSMTiWpXquZ
ET4murvTewoTC4r0B8BjWWwdiYTXQI4d0PFi2V0wDGD/j9qIoNN1zKhuUGTH
cw3UAYr/i7wysDEtIijrwF4FzDTZCHuVHTVAbpa+nOartqTjL++qarDFuI9I
ZBxPbVgEffLhvW22hyLsPgvM+SgtTYAsZ5IrTyhXB4cavvh39nHvekSJHe6G
r8wxixaiyZr4fUuwZPuOGDMf0ssYEnK+c+mff+f+DgvQiRUWj20IYFH77vAc
mZKNdkEvLYwgHENmEZDYG+RQG35rvqpAawD9dRML8awwoz6KaPXFYOqnGb2j
r5HWajKbIIy8+Bee74Nf+t1X/3BKlyYExIOvq2uTZkTArp5FPBL9gl+RFvHN
FRwCdwpWvpaEuOyWl22kQMtIkNKmtXIX4gtJcHNUlBF8tG1b/U9ZZb9pH/m9
Pqc1/1rMcmDDtZt6HDyTySjQtqOJ+yerJpy8XqXcHPE4dGfuJ1uJVLLATqUQ
pqvIOSXN8JKSn1Js7YEGBwuyVr7YRECw/o5Gb0bDHwqKoW1U08z+HFFFUD5O
e9YwPmwDDuUETJf8/5ZxKKm/UrND0O2C1XIMClh/L7Gh0D6aJCnBjhim25iu
0ZFOSURH0/U5q4iI/6JFjY5XvopI6p6gbB5shpAy/CaCG9A2ei1JgdD3q7zn
AuNXdOjb52XEDKY2Cn667F4jf8kOmzTOUMWqM71eFiKPBGe9mr2bFJ7QjoOw
9kWSYBi1LbLqJxFOald4lQBcZXYanOIjjr0L5GIoX8FopejeQ++EWHNrV8WC
1/DeRBzBiR0mLToOZxP4U1decaU9xqIPzVTLtnwQpUqIjYGL5M6ouJfQhO7m
Dx9RrcvVDMG6NAUqtYrIvgntF4khm/fwxfq2rJvcm6GEFIRQroCHduYMcfYT
IwcIa9mcA1NofngveZslWGwzio6MdYytErzfxLy7a+iAgyx4zrQmUtaCvr14
HrhT0ijDVilDqlbsE+LDkZ8tidFLy/ZGleFT4zm11k9lTme6/5BpIrt+dZsO
MT1jHX+CW+Vx6flwaDjl+cADIxN9eEt9XQysVGQ4EsfRronKxOcJ76sLQdJh
+WeF6c+NuQp0Sv89ZONI9fBFjod5Kf2MhYa0lSEEFLQ2d6HceUc9twmu7U8m
Jqmd+DSJR2P//6VZnn6IIRWNuwFNAgaBIse/gSeV05jAC8ipJAsCV3WPI+X/
ZLzeDBI9jLhwaGzanQPJFDhiZR5T48NY9tHfFsmVchR7n18KpHpRcf8oEWlW
Z+BbTcrqrqdCrZAyWK/FnfwVAIkZuoQiGPH0PPEbQQNyE6/kqKF73LRD13HO
B3JKwlYQf48O5xyzAUrKYCv1UNOvcIdDc5xBpDp17h+VXrSwT+/NuJhEol8u
FSFdGxBV7EXRWzc8IkuHsuE+GttyTBjAWsNEfd7Gq3GYAfNYuuqUqlUTJ+ZP
05hbTwaonfAmi3lZf+FKKB7mp+fGA/87N6H9YxKbyIjScKTvFfCCqJ/dfgyD
xALTXajGGGh/2uLpd1RNbOPeqo66u8ZvdexCvqleWG0y7XbRXWN+bW91xupd
Oqgq/HK3mXVotYwrilYA1YyOPZqjxkDw+cm0lhcucsPqmSyG1uB+FD1q0CDH
q+DYo3Gu8FXIPvAgG65axz91/Z7u77gBdhNcb7j1bvxECf2qlRasN4WGB43x
NFzezkYP/Wz93kP/L3vwu3Ne1SLrgPpkNGR5HCXdrBDz+dvchtGBDjmG/bS7
6dCu/fJd+JdVbuylJTYef7wdgWpY6WJd/tWZjIs+98j16VonqQNjo48rRGCH
PzK7mdEfaM7gRnTsRq8T6nhkTLRzJ+urTfsuf6pHYIGdBf0dAHAat0SkdVgK
z2FJ24Nu0j0DrJjIFx/RRTM/V9m439VGEKlrM3vm60QizSRgAn0L3VdpxSGJ
KQXRMNKXvpJcdEWE70xnPoz3regCj+JYCPr4oMpi7A0Oh+nfT3TfQ0tGX1Sm
yMNdgGmD32tdqZXko2BougMbGS2j/yeaUDQuHAq9K958AYltr89c/b3UGIle
d52KZyRTRSr9wLvg82JNdifzVOGWJHbmnW1ayotEChOXMQyz12RAVjpNLN4M
vZz2ohskSnn1qBXXhakaURwFGiUPPv3ijAlhsiSeD1MjScejFhsoZj/6rqcq
oud51gA+4alm+QQskOTGfZuAuNmWSgs+lqL9bghlV/HwlCL0iNbboTEAsB3T
VnfdSNqzL9DiW1uCXpkqr9X0sqGTH8ULGrQMGMbSAC6lXyqzz5RlTkRM2Cgm
qK8KNnNTvCIJOtj0MYhXvBwj3jGkAmZMs0zzzJqZIFyaFrAURp37Fy+x+Cjp
/2HU/PW+gtAc1Fb7yzd3m7wJl6olmEYkigP7Q9V4plFcF1frzcBjH7pGXQGw
QFbI6uaQumMlShPSZRagmfGADB9cGy36arv42lpws55PJ2i94rqTceoswGtX
1mMpx1BwZUzQtYJk4ygQRhwb1IEgVtrKqdk6BXI5Z3mYQVPViK25auLImN2n
tmoZsJpi1xEYj+ajymup+MyvrdqVt+cjK+dkn9rHmlpHnbtpjPT0rErZLkSB
ecYXKLdsYJF9USBFDcTVtIsPqulToHz1etenE73LOT/wv8ahYBdoCgzVrwqw
0aDfkcBGEYzJasXMvP/6a4QXJWI/17T8GmuepYqOF7XOpTMY7QwHk3bltiRs
KWcb1Rgb5qF6c7Ni59i0kc9SoglVEpTjNTt/VsRyS7pQV6rbHTPPejjAMOF0
52gZkNwS4yMZXhE7LCTUcP7LDdhFfbFuDkgr/7umqhyfAUKBxH0lHWUeDPZc
KJy/LetLeZueo+durIwPmIrr75jZgbuW7pz7EIRImvB4xjIOqajaemxfQ5LF
UNUcor/L6PemeqLAbECT/6asbdSlU8sH7X57cqkl/WN5Brch9Lt/99nNFyFM
7N5iS9Th62OVWFzsSdYJSyM+H6OnGcyRQXyzUdsbUlWVx2Vgf6Aq9+38ZLer
gwA+zfl0fjId1gyGfw6aPwmK3eN8WULinLVpNzNkXtDJmPav+CPUE8cufcus
AT6a024cj3Ch0N6JKOnI5kRFKauYcMOvFjnPhOUQ1vOV2soV9DRNw+sFLUKu
jEwUCARaAIHk+p59XZhUqv1MtqCiF4YG63VrMke1k9ddzssGpw2ydl6kTNms
fVJ/Du1UPLUHE+keMtBnIReQzbqLs9FgKOod5kaLzdLFokUBrl4QXF0CmCae
X1LohB82+k2CIF9rIgbl09rBqdLWDYnhnOXroQuOe5xdIQWNWtpZEldVTjuY
toW6T+7TO9gRH+mXV1PDu9Fz04vZ2YtcxQWJBDyLjUdypg0VaEoeqQNe3OZ1
YPlOr7RKpdUOISJETLP/cJm2AsTYvXAeWgmPWTWBGP3UN8N/+Ky9t2sbzaln
WC4MnRO9Mwtt4j51gGYykc2Q6EWVg8nlBiHFcg1/q7ftAK6/iR203USMpJEE
f8SgnlurunExuYdueH07ymzQpbMftvpSGmReRefS4pB8JjlFMVC7FYXnZSY3
mOmfnhuBFYtYQYhLjCJARY1doUy9AeJL6q3Bkjg0z1UPYcWlKOpsjcmPsb9g
G67wDi7ZLkaLoKNxS3+r007R8fLmktl9HcBHezRA//h+eMfz4mNPoDnZTzc0
fqg68Humd8THVDWVrpKdEDRvbG+PE3Gtpd5LbAxpxVaDmK4s02ihUv7VZRGv
j1e/1nDPPDsGjf1M29WSjZ8Y190fA3cO6bwIsLiqaPR2xGZ9xajtSX1UtiO9
0EEoepw5fnc8PKN91cNyLEI7xOAkzVmsVXyezgOujKmvt3jm6mTw8xqk0Vr4
+WZADYG9wp7LaKGo7N9obo8Ik1MF8mvQ0mPh9yx342I2X1o1a+eH9o/c9M3i
1m5LlnQP7kJO7aOetXJwGxRSKW4xDYIosypKa6h8qd2pdTeexonamUHak5MO
HoBpeKiqZ0eSiKWj7TYhxKr1WJg7grgP39oH2EgQK+bCAmg/P2vwnDRPa73Q
BZN0IHhAzWCJNDeRZ8+Lj5eLdYN69HK1Os4nfJsrcQjTPxkQtRmINGkFIA6C
pGHPi3BF3LuuGBSws0o5vYGsxE6ef7nuQIZSylTTEu7mmJyMqyz4yl41BhZp
3ZyJQzRoGb0DDKbHqVDLkUjtt0yf49LtY7Xby2C0xbiEuh5ptZT42JPWTDqG
sAbd66KJnqCKf00mQ1pQxdyiwgu3Iuw69vQ++sDHJPvPsE1XEGW2REYjAsnR
b186e9xHql7pGEKWttLYTyukJGJdb4ilAM2PVC+jjKD8ukXjmy1aZN+UOFzh
sx60s9c0BXaKOR/6w5cyFU0EyS3Bdd61c5yVUl9VZKKyTUyoaaFr+7PJePyJ
mMrjMvf9xrqweRvMsqIGxkS3sYA/gUmKixvIR025QxI4xSuJcXeZF5bwuZwv
sEyAJ9Coq3xhyDgCmzHDeqV+snbgQx8E3k1ZzO9h3/TLLdrcU7Ief7amM8EC
p8UZEUS/OYiEZkYbnOBmM/QwoS14TiP88uWv7h7R1apBLJ1D1CHfJJSXy6TX
BKjR7+ht41EbF1Uvoy4cwicXGPge8ygx8Op+w4XSJdzv6stJY14c6lkFwoMr
MDybAquAZlIOyF8r969qGAuVkvb+61ZqIWHEsDM95o83VBt6vFhgrLFeKNqz
DL72Q4nofkg3RetYsMvXo7lqCor6wOwmTCsTvvh14sqhkDQStGDF1cmAmpMC
u/hDsOE8rHPdrb+1JRKRZvoGcKWgjLK9tUnnz6pMkbux/npzxdt7EE/pUjCK
mB45IaVTb9yYcB3oFdjGMHf+bTTbY46liK6GEBvu9UQAtKNuxpch9YEEPlX6
OD51pqS0G9mJjHgke1PkiFlSZFxb0qq53Zb+BIZSV+P3R8hoCpzk4zzLZ1nx
ozMp9W2VrvxFWidySUksSY/jnrB8nTUj0g5CA/ycJDWN1HyW51lXu2TnLK/h
DxsEyfS9HtAWJEtsS/dGfLvcNj3kM9AHmdkuPc/yoAakWi+yy5yK3WIlzYcM
4Cribf5vRPEadVLp+SZb27tZdsxP51wbmrR9aGQ1+YN82ar3WG9/C2SE7t6C
Y7S2PbTrpt3JIhHk5WwXRbE3m5a0OLy/IM5MAlRYH7d1ov2sxScZFg1Mvcen
gR2Nva0SIpzTPXu9PfADExLrGEDzZllNYlMvhmyraxxykQ+amPIQnbLCORb9
RyXpKU39D+G6fFgIKCVYzFNg0TZqDXJU/prcDReW9PEfVBJSUQL63zdT+E4z
CjZP2ep11SncmhvuxgNhmMDt7Xp6amf+VkKu+U1WvE7bW+Hp898H/gPB0CJ7
F3r3UiMidOXiF8v+T3mJiDkQvphy/d/eHCJ0cG+Kvcq1exBQU37PwSCTps9r
4fu4AtBDXiP5jeDOJHQ3x2pUD6xth/is6MiUxkLcIbOulew3qaAf6gRBPqQv
xmQdJXLRU/B37h5SRlCiIe6bm7NZUPkn3W2C3BUumvWeFu3mibviIzYmfLyF
/YDOt1n9pane+Ifm6C7UKcDDPZddEun80t3IAtetQznR4ztET7Zu16mgyc3O
Ixqp0t3/TpPxIrbkOME2/aHS6D9cj82DcugpQinMdOMBZIX2BUocZ2b/dXAA
YLg3sGwCoZmZxiYcKnEvZp7K5wePAEZ81gN+JJ1bb5iPq8CJeZ9tFOwhDdXY
XeIfFL4Xsy0ks4dDtJXTq6TgVy1f+qJ1aOMQZHehSBLvHCoHNPm9M/sshZL9
ew5PBP1adtpzV7MOxM7gfcNSGru0nHRHbVqpL9m81ooZBaJbEcm0bKx99SB2
tWGkbi67bXkRMIAzG+La2yWp6ET7Q1ChpVWPuM87z38b+P2QBEOGBcmggj8+
m16F8ry/fi3vJYVEtxsnE4UWIWahE8L+YWx/Ax1QGKE12a7LdJGV7J3KeMwT
IJy2n7eunYVTquctEnC4OFwGEx9guyHvujEk9F63uLuETFpkXtqpKrc/UjTY
+vykoN5TI2+AwqGrtPKUl3dvd6idVaU/8gtkqjQwddFcYfnyJg7SWR4z6CRc
DtZhxrgwbAF3LOnTjDWJW5AWJ1Y05G/aymHy0kPqcUNCzQChb1GXIoOHd0tu
+mssT84/NtL47WDx+WU8LPoC3biN44Yqi+pGZ5wwjSRQpXPcO8npgtNsrq4U
98/CKA2pf2cuS9fP2KWMloKJ3j5P1/ZudcXsfjNpt9tARByjkDa4k2Y40mZh
zYNr4cG9cxneZan0G76K7+lDvX8t1HZ193xFDuseC0BT6Fc4j41//B8hXrJO
0G6AvOKSnHAW99e213MMicmYKI/viCZQtpHiLD9afnAlz9fZwgLurjIK+bUn
slobrm0OkqoqPP1nZPYNT8S7I65wqbyafA99DdRK97lwWyJRNCctieFvrDh8
gpZy5gw+0+Mx47FUVisSiM+fO7skq5rrHMEiRNYCFqZ/tHmDRp1TOQuylES+
Ugeu65dz4f8VbbD092Tx/nONs08sHR7J0M+JL02+LjBOIeDfYk1BIjgXt/vJ
nAVeEyCvI2MsbUgdnoZG0UBK/wJjThqmTmcNd4T+IAR+WKpsfub/ePTe1Jz5
tvZ1Sg4/Jo+oeNlJJPchgHUlrsSN4+UXCNxAk/OwhiNqf72fnxDvLUkmhGVB
Wd0l/VAzxoW9/+W+NTVhIrDGAeLwKxwtkp3VNb6aJWxMuFaHiB1Eyvl5OGuI
SOoEzPCtghsCtzQXvM5Fl9MjKwsHdo4XAhFFD5rcagAX8LtczsQ8/T0FFD24
8XNVbztAwRYXKdqQzdIIIbzylQWpRkWZuP5ZIEdsTm6rfZPFDUPDJYy6gby6
wMZoAml6H7JgmL432TIcMmezuG958P2GIHI32rCBvPEvcXWzLBXyryD+cmbk
kk2XkKQdNX/F3gf8QgaCo/OykwRsant1VM5KA2Uu3ojEO/jK/qrco5xk1oMu
Mp/0B0S6pUnsGzo3ks6uk768stIDB5+VpbXg+lkEl99iLUUdhZj6vWUhhkRi
PPu1SEEgsNGsvdAj9uHin+HnWRv8E1XUJGB6TkS49v31v3RbPRCLgcbgv9xP
Ldg4Vxy7PeS3p/KGF9NBZqtuFSpD3+hh5LrJ57HnPOX/mM8CRlM1p4LbkVd3
CJ8qkZZ99e0nsb8iijxDKb681fevS6QH+8wD6TD4Bm5Cjf/0G0SZc2eWqgQP
wqvuM5HuTb+CJ7pajR3i7eGXSExzVxQm6238tZXGICNe7tMnI1wV9S++/R/Y
VDmFpM9U+XJ/5vpTtpGBBGh+qE5Q2l2iZK2IZRlsfcK0CvSFq3gGBDXK7oOg
5ABt87aYd2PQcl0EhXThTHq5gTUNxULmwgYw79XLKs9p4NlMh8Dss6vg9K56
WRF+Qq9MTva+5pYtu3s1Jwf7AD38Grz9grVxIBrlOktPcHzHa+QiQtl2xe0S
NvrgnbqxDq4XrzvHjx1GtMIG2a97xMY9z9Fwgy8VBg/wscCQsq5aLntP0LFU
a1vuJvhyKZjhh9M0KxR3t4Gl4Y2yb5fTv/lltqpTucBXdZYEeGt8zbpEF06G
LyHFu36P/WA1/n+UIit27IZuSvCAvk37qNeefhmvOVvPZq15Ch1cMAZgJOMx
c6AzID7qSkrT6R43ij6V+CApCtGmfJzu03UGMREd7MPbhJLq9Pa5vm8i0bMO
GZI8/r5jsZHKZPMh1WWxKDmhXHkm0hAxwuf9DL3tG6u2bcGxngQOpCgdXhBw
9srwtiL1xD3Snqi+SK3/QiIvXH0ft6T1Qfmn/naJSOrveI2B9aGLbVG/PxZu
IsmIxvJBcaRzaOXSITbRUINiAe6MDcbaCAR2X2dA8jmH2MHQBH5DGffTFByh
Xr75okl6BUAEYt4MEXASfDpfUHXcnTnFLSXKhrCscimUWvOrWxfgMxrGIwPd
eKlAh9QnpkVJzE1JAzBEMqsGStrNLRpPu1iJQbVXc6FpnzF0APYnQrLTNVs7
o8LE4sshwGezQtroXO2WbvrS7yQeY0ONFxSXuU9feAKkHZlxHlIaURvVwINM
ps2PWTHxj71N2yTvP/GAXaZbkFv+d4VSxaR6o24ZWk5BhfcbxnXPbudHA7gG
e+P0nBizk2bRzoUmIhuBlDcW/tnJd6NW/76JK3l/VECM7BJqDd5YU93zefpU
D74vv3xOpdRUzvrdmaLAdRyt0sZgWVueABi1bwMmomNrUtl7lu8sqbHXWJN5
BmIis3pU0ge8Ok+3T2Xp6v1yPwetsH/8Cg8IB+71MEt0iaU4cyvD8vd2tRsI
WaHeSro3DMEkmfqg8V3G+an4RA5xJFMTjE+g8D2PqPv9gPIridjv+FHZIMoi
XM1hj0+JuuJwCcQXUJYgeZoYjk26Y5DxJYDj7nrRYUwdH5PO22RjYqWOb/8l
uedx7jFn5V7CfanNJlqfr9wtMB8N1WZzp87wx/b2Q3/Wne0W6UV9ed2XBUZ9
0mETL4GEsRgQ8sfoewqEUqNPSq4+2T92G61DV21QeUmRuztOWF4QCU+8znzv
A6CoYQvBoqy9mfVq4GZ5aA8VeRZKTp1VT13hHUwFjasaE2h0AcYcijdJ5cC4
gUq54pwII26CD/FzY8v/JeVSFoJwX+tmY08FIgy3UVe/uEAaQmxweTqZuvmI
f4wJyFBxIjVQgOukJLydBRElPTiZtjZXzTasChAU8slUtVIV3OoMyW7Nr0Nl
ceIFVbjkHSQN8V3yF8HSN67D1O/afPcsUnYqHdBYCF/LoCvEI81sSxTx609A
ej3ONqX0WSQlXY6KS9xNqoJUXTQ0JyF/eu1ZW021QrvCvJaML75xxG1z4XVz
TrEpi6IX+U5Nn0MDhPuMFC3S59EqNM9US1DreUexxOXdrU6UOfI5om8U0z/+
h9Z9kKpqB+VGMjBl6kTWV2eYLdRNN6RU62XJXWA2PhedGzR4+H2EuxSSIY3E
jzvFOVFwVoPnWyMf57eaDtnmVmzLXw5wWJKRvcsGtZwQ3VfDk6wLONApgaxd
Gix+/LV1qDcrKjYvwqM+QHAA0JloXNrZw2+uJmiBRpVc4nKTeS3cGX6+VGUk
yJFlF7k2Hx/p3Lv0hFBj8EyWvV5xzylg0HAppQyk+7V5JltOUCuzkbmK9cW3
wqa4q+Y6XlP4nXNKJmp7nIcIvqcoNfg8B22s0hUxyEciMfSnC75TW/oYbHJG
+zpmfO7gHPdOw25gJ/tkvST3pH9N8fSP/dUbgvrDqpa0zTOxsxe2YoU1Fmc4
4EbleLEXx1RGipH9JYQhO3Y4Exyy/4ZOdIGts1dPbAvPGge3eDd5ARnNMX/e
K4r0f4TXZ67RjrJADuRy8DJK6kOwhiqrMWMZSvuH8E6E1dbQTAciM0Mbh7Ai
eLYNBP4XXmfZ2dlcXnQ3Q2NihJoRtO3PITfAw9wX+EKOFfwYLRHKq7p9GnNS
/e5QvlTYlv41RpNOTXCyDIftNujwRMykyaItxD6b0I+80/ywnGKNITiY6StF
qHZelqCIQriCqd/PU+ZDZj1NFFWuQydTOaEjSx1aLV7k0wTyE2vOtk/OzbD6
JVdJ9hPvloqaObFzM1Hnq8FgNYGaJgfFKCvG15kGsUaHjdnWBkctcr6ylkC4
GqPFG2F+Jx5StywqZHtbJeJ6YzEBDP+ZCMq2tJ/5H0to1Te2rjMJ6ZM3L2Vc
fQMT5xEUWBHQkeF/GPy8iqVdEyyQe2eTamAkMtDIygxSnJzx6CvdrKtFkQRe
eE6rD5fsmFYydHDOYWdEOMCJOW9gRNGBtLOesNYk2VmhG/hkDrwXQsgLdKVi
3C+SM7Ei9Ek8iSh5Zyw1xp0s3adV4z15RoaSvgzNHbdr1hm8wOi6IzgKLmTt
4SxZMzH55Rpl3PYE28RmLfF/TPgYwJopcGcg1J93oJCdsr94hR/aoBg4bVSd
157sCAuXOOS/fsNDLxqyDqC7B7qGrYTrMkVCladGfRcTqewFxUmcbgk6Y0ZG
bG2LoDL5x3FvOiuvxygNFoVkTyGSdCple1LaPqIW4Y4yJJkdWmOP1SRBg90P
aHOJ0JJfby6GPf0R96D2gmRNHplpvewOA9/+Fg6CTQdf2N+60RGVfAigGFq9
VRqqTy40yPBKwnKwtL2eNru7xDSpYHund28jb2Sw3Rf1FXiTVtFxmGtW2Xcz
GRmy4VYuhHrZrLNFais4Ll2PeOJ1juzEhNL3HwO8vy2TYTuZQiKla/r1Is14
T8gXsHCV9c5aaLIwIsaHenKP5YmUtGSBxNV0RVXO8NhODoqjizhX8bfZKTUX
c4uiCitHVBjN+bWtXWS+m/j6M5MsqvJMg7uZyBRIbetRDZn8H/tIww5VFI9Z
E5Mtcj44+dCO4EEcvSG71xvPgu+DXzv0UG72Bi2dmZvTlgHql2p/9Rl+c5DZ
7kRdZiat4ZBGlV23BWg2iXwQ9qoA/mf5Srj9BfvqBTaJgNRAdOFfsYdeMbGf
vIMwPbqyRs1Phm5wuTe6aFkBVueVcZ/7a4SfLkvsPjaKhK0BcXAvmk4cgJmL
tkuslRgdUi1+OAFyUfNklTrRRkI2y3cBxh2tIIda2MUGptk5U+hbIog5xEA7
ud9NRVQjUpBcaBrRfvLutnUcN+xXY8D/K+pMRaaVrQ39ewfbMsdHe6wKy3tg
mhqc/LaCk8RSzGTifWZ18dqYijMVHQswE6pTNWJADtouUlB1vD3EfwZtbSzz
R2hV/eZ+rpCl4/yhalYrvBOYvIJ2mEma53I71LYbSmg3EpVkPNL39rmUXV0s
pcVAQK0wgs5YMg+DWDFuqNQVR1vgJ9nVUAwNe3NPgMDAXSlsderX2cxeb2ns
VqDpo/ybW0j+ETr427AfD+VO7GH2djGns8EiMAkSBudV7KeU16momn/TyB1s
VsSsUIKBPaufUM6dDL+HfPHn56rYmTh2KH2eNAtFme8TvEXb+PCoppe1O7r1
Kp9oPwWuOO9ofgc6c9aplnKp0OMZvcUmJngDqEPpFEoHB/hZAUIbjke6d2Hv
WB0nnk39lqvakKhEh7XgM3EzJWcqDfeYBiHr6WtJX+JIJ9UiQIMuYrQSNgY4
1/Fjn5nQ5xgQatb5iOsaqBJpyZGeNE2DGLpglQnSoscRYEf4+9mGURkTjvZB
LV7smMlFk6VnlGfyiYDyNQwRaibSJ90rJogUnT19oAXOYWHqRZLpSj+Ag92z
xMq+k50J2WaunbCzbZy7psuIzBnz9TeKxVcGiihh+Ohd/C9cTeEFDjXntAUg
CtU5BSnM2L+sLpJZslpshCzw5d57s+E87dgz82KJ9XFFl0zTek/fAEmB2SKe
OkoypYK03oQyR2ShvFLqRSCen5mWAcsy6/1pW5xtrodo9Mxpu3fgD0Ss+CU9
oE2BNs5hurSWod2tm326hQhaP/LnOtXTE5NjOI7Apj15RNzXvvVCEIoWQWzZ
Wu4hwBnEafGdG1xOITNdMoaAI/x0wg1sSbPwc6lgp3A7MQRQgWSRR7m0j5p+
ECySf4bsIsjy04y26hPS+5wycw2j/jGF91oxlX/NPjJlYnRrky2Kbkry/sPX
Mbu/thr5nG5lJ3ds2ugsJkiyYroqh4Mawlk+SNgedyHq0XHXgYINLqQbp6EO
G9I3vsZE9E9bztv6rewlDqfZMgQOfo3KexLWWF+FSq6zA0WYPI7YISMolwO+
OqyEW5zfB2hkd5pob1JoOzIdX1Q1puQ/bs3vPHUubGREdHCbXmFPQgE0FEc/
OKypxNqc0kRcpBbCM/ODOqIvx3zTfQkRuXQUPHQv/3WIs3gOecfnFELyHLoE
aRi4KsrDAyme8IM4SHnOCPVGshZeHTv3O7PWrWhA+PcgFzSyaSPig/g/6rRz
Fz33EkFD+HmBAMS0SABOw3BO/VD0ud58zmAFMQgexhgOVduFS7XD88eBUyPU
v+z9sqkY8XoIIhZBBHl8tmcCSh62LvX0thc4HE+29Z4nrZc8NrjJQQTPIxFM
KVE+eCo78OVt5vyAREdjuLTDZZTF3Sw94Sc5O/FfW4d0B535UynpW1j+gtjE
jB2VXX8xuHiac21dwh23RYr6G+tJc6gYGtYEhNi++RgOdVPN7I4RpcXhnEIF
3rzSnGtUgRL0Ebg6rd0iKx1fASA8UnkGfKMDVaR3gQkbe5y678extRKrkVOr
AmKbozG/AYxk0g6EvyBx1lNEPfZa9ch/gBowXg2Mntcwc6NAGPHuBTQWxMKX
BQDaBj9E9kbWPplZE0d21ThHgYQ/Ef3W/Z4w4wdh26m4aAzU5UMPLtyve2VN
QpBCPxwpIqpdIndt2N6hnEza8jbReV1ZZgL4/P6aP5EmG/ZchRSEDMWyRRdS
jQuLbHLWIuJd0WTTbwV6VuWpHKmizZcCKAFOkq/hbaJdFH31dPS8ENuz2bN3
iU4GDP5egOO7wHy3N//XtG2kvCXf7C0HDjpWnAPZaRPyHrmnR3ArDTwMwlBT
QQlPg2gnv7T/etmzhAKZyHb4b+2KdBlyVzM9rPMruN3CxKIj4cgReVtBr9o0
mEV6g+9VL1WYOoJZbYFLOW+LZxTf5KV6JHgqSsSAbsElZlzEPYLO+xKn1MUo
NTT3uzoTt0NltlTiQqcPbbntmHRCRSCK94d0A5G3uLn2HM4axAduEgJBKY/6
fPFqCloqmbM6x6MHgnya9phv7WDY5cIa8ralKv8N82vk3X9x4PMuoXqmoxSf
nDELFDIj01TOalBDc4U/B0lGgdT5c5y2pvrJFpoVG+45aCyDCV9teAgtP7Xd
7ZeA2qS/qYfyd5MR5UboCrmKKM1mW7rUXPrgc+XhM2dUKPUbbIEbwXiU0MEE
PydONhopwE0NZ0cz1l6z6H6Q8VKd/ZCQpqO20rN4aKNz+b36ucQPCn/2qgJg
v6gNpiLN6VpMO5RUwF08GKnzenUA08oU7jKm3frSs3yz0s/DZD2sojJQd37b
zVq6iTQkHx2uQB18p55Oe4sEWEyHd5eHYR8B1z5CSGWMozmrmGHFJM0CcJ1P
1u7TVT3Y1oggfpO2ZFpOs1KY04Rwsne/a2l2dG4KroSPJ6d1FK6E93bnOzco
e5zMNWBa4Kla26no5N1Z6bm/ATByJ+mZDcKxo3RL+hp0djzn/Uhq10XKmde9
KCflwApiS0yBXblVniVpSRBHNPXv1HUlE7t/OY21XbWRvEktoMV2mQb5WtI0
D3Y/glbHu5+4UWQIUHes2yzLe1gaPljGYN5T3xB2EyoiWh6fp9fu8YDF5EZ4
Dtxh2wW4ijXi7IDliVxuOPUNFQbTI07TVLbKdGr3heYngD+6l8EnYSJWDqTc
W6uldNOCvaFmHGJa98V0OEvPyaXwGzaS/DvhZJwnzsdOXdCpFBwbenkdfTX4
qZBYEqIigXgU9hS3Z12fusT1KqLgV7xegoElnBcKPqsxVJcmQStiwbSRkOlK
X4TLt+202fS8qvdnpu2cknPV5k2wVAzus0Cl8hO+7fhneB8t7nGbFfzHaml1
JFkp71SQLfZSr35WYpVkpUN3JiVhMUTYTfeUpu63f3PLG6hkmwa5SqfHae9S
lvM86BOZVSZG9BsO1UM3DzWME5JDlpvqlCbKFjfvVAwT3T/FPV9dtMMhtSb8
DcZrESLmEvJTOdReSCLByjA7UcCUz/vjY2E4EqpSN3tnEDUInKK8lSPfFZje
uN2qBwfScTM/5xZ5o/fppqbke8MLcp6Oig31VJjEGo4YXnVHhMUcrogQvC+s
my0VEc+Hd6Rju3WnhRgxffxcNRsii7ytqg7omXba4XVV8kJiZqys9J2IfAmx
vGjwOh3vcshb3WVW1nQtyfn47/FeuikejtXwSi9kXUF0Hrk5azGz+Ip/egbp
hRA0EWXTtndvD6QZlRFlUOcCl/riJTx2pOy3m3DrQNAXFG7n43Bplyd2enaY
1GWZVe96Jl8eFlAj9Z6BfgYq5NceXcNz2eXGLtc3M1ghoZxl4i0zNdctkPAr
MeV4Io9A2XmDVVM19q08/nRvnyTHILjgNSwCXM1pRtK+7+w6qY2Nrdz56eq7
a+fB9gpug+LnQThWlyoNpa68Wq8GOHM18lMa3GiXEnGnpE2M4BsQk93CDfw5
7js/tqAGpylcy9jHwroZcci++Khw6va/+p7ruyYA0XlNBKYdCBcEUSIZHQ2h
16MjKFOx2ZirMPVaE9+lGBpPU5Ntb0H5300ByoWGKsJ5eQ0knT19l7d+akTA
nNYo8Sup6BZripbd5D0YF1jWXL7yQ6qdZn2M8t3/gkKfLAgnPVT2FKHsj+4w
CJgmV7VTUuBJuEXCmErPVdp74S6M6KMFPCf8Q2PRWTzx11vO/bM44gFkSXd9
w60DuXvdC4K0tcwvTjNVDbQ2XW8TbYAO57m+msnBMQVkQZDPTdUleXOZ6xkh
cJgibzAC5pBxj2E2GjIXoGFW2uuOKlJAWWtahXARo5GmL4CdtBn5FMZxgnoS
ncCo5UBDM8U3LSoaL9SCcxpSDa7i51fndr71+KGbp/486RnXxazEVKECq4Sl
O4L2yK5yfqLCFFdXRZaL4p4nz0pBLHa06yOGenv8DlZyhrYubvZMYPfxLhrO
NNXpibTbCrivqvC10nIXZcF046fFeDMT+VcS0dsKo4j2+5BTWsZC4jY1a2fl
MYghG2GTpMm17z7h4HxHDvPj/FjqRGnapHqffKzzbXXoUsWna+DLXXkCx2Az
u3MOBSB4uuxFUfNzvlscRBb0zE8yhZygxuOfQHM5OYj6CDjhYDARZqmnCyRI
IXi4XgoEWXGV6rQUvpuoiPqIazAEZqDOilpWnX+j/ksqzcbaETsVDtIvT6Z2
xyWRXozvaRLlDHdl0necknZHnrM2wfku8esBsLU+sd+r6OEvS2xkJ741b6qz
fvPLLoduAmJcW0ttBq4jTPmjCmJkDQtr4RY3APh5KzDAevjiPABe44lSjEof
XNmWdd11uW1oJI8TzvR7EjrdsoH4UzC9AzO0F8640sdox3YG5zTCErej77Gc
SfcFNDWW9L8imuTwoGZ4R0FqWk59P+kGS2zWpoKgU5JZu31eYJwTMuS9/uRc
4ZxvixLDf9j96ZENyxgauR9LnrXWbutqmLznjeujPOHfYQzM7p86V7WYw7OL
+Bwgjsxw+sbRP3OcV/KyIFhRWlXTd/9Dh730n4mKc3XYub1i9QGSJeAN38GZ
pNwH95jYLt2M8UERPGJtkqm+ERbcPmAknGKATFCODsFuCtey6j6r4Dun5msU
b23ZhJJjZ0vO3jk38rFeA81M+AfbC5CY3fWyZXVUdpNkdsXapwZWBF48eLrZ
wi1RvfoFt+Ur8DgUzx4u9lWPUjfWVVsrZFI9zr2BrZlUEfGNbw9JVLugw5PA
KJm8j4fVv63FDWjeHefXPxfSZmYE9jRReSaxPytg2PSMUE8vZaSCKYhitH6y
OujEFc/39mt4xQ3n+5BMMCAKxm1bk60yOaIDDYws92H/ODpVL4dhYY/Oikeu
fUEADnuHRqOSTAN0+9zy26k9uLrsuVq9LM8YNyNT1pVdM1gqNFsxPSLYEeV+
GxFGQk3Pwbt1DlbUlgxwgfMtNKJYnnfVR8OZA51xgOpFwRhVtE4i+ECR2qn0
zt8l++/ipL7+Rss/z7TrIaWBM2U4UUVVq/920z+ceispEh9eA0h7pF8T+1Wa
FnP+B4DPHUYnfGME65sTSozhlxawLdr5Qze3gb2WfKrcqwf4TKdcjNT5uTmW
/Xf0gvJ3kMxZ7p9Mwv4NoXDFt2A3APcBvV5PMpW+Cb8jiEZ/CU6XnGu8DkAV
md2f9trVtyDnpjJKpDPIFt2MjTj6mRGxmvDNQun1vX86c1o4aV7yfO2MmdB/
iA6683eI90lye8NCUlTDlOWlBm6nB6rNIXpt9GyvKSuaHdlKPgAaQArkesXI
ectKPGFxmzLfjpmUPpkPwx79aTB8zxSZN/pPbqlrE6PKwdIdoRQYXdbiYY7J
ClxSCDDvUQ/IsvVs+yG0c9YPPAdtgxbZHcNRk1b/hvoNgqCdjefwTeeHIC8K
MYcZnn/aUE23CEYRwjmzmF/ZikxSqSQP+fbnKvXg5Qx/JcCYVKSuJo+G0ubQ
W8M48IOe9nCAYAhqYK8Lan0fqXsJpOQWlFJ6jmpf13vGU+lvtdo89d/aKJhC
nVY3xGKeEoUFJ/PfzITO3OZ0+tUymgXqTOmbIK+yvEIjvMlTyByVGyZuFEA6
guu/bcvgQzFmEeca7E1gas5/gRcLLBdHDv82CKmnSAlolCPZSiWzyUBGRykp
cy+0GJlVeCdHlnlw2bC8hUgcfnkSS9tvK1Bc1tfME+BeAL5w53dKWEcE1pMU
KCiMhnh32x7Ba+IfKLQwIDlsx5TM9Z4WSaNNjclCPCs6294WF85u5IGYlrSe
SrLJMpSMbkM4EUS5558Jx2teSXjfJul9pvTPooi9mwa+9gy8SJnIv4cfdb2c
nrTUl9Lb0qRiG3vpjlwlmXhppVVEyIUITuJDKEywOdSCAd5Cb4YNu8BBsoRb
iFc1Ew6YQ2f60ssvJm3mTc6wD0gqRq86h6gNwwrFcjYr0yUXzQprnE2zrIzZ
ZHOQboh4m/O4Izkubmc8CIXUTJ8qMKP2O1u68qOzF1wARKjeZoZeCsIN4KC8
rr6/8XQ+L/g8Kdgu9+1QVQBZls52hDnyv+OsdzOLiUbv/g7ncVeaRSu+gMYi
kotHRTuV3IrWQK6ezRa49k5N9mmWoJV34QlW5jeTrNFa2j9SUwzt+5DdACiI
eImoYTo+AKNlo7XIMkr4xExM1JQR/Bam2Av9MR+Fzz0gIYk0PqjkUpbtYiPn
CUva5OFdt4r5KsoG+WN9W2kdu9GYt6Nq2BXq9xYaXbqDQcpwXCLBMplz5qcI
qncxdjJFNaXA2XoZBpugmmIDDJxnnf38lApKXvlbXCuOkbqlLQhHojDU6JU0
VVu3ATIS+G3Lt8JgVeNUCJc7tnzMJY0eIEc1bL5MnRBz5XdQlZ/UfWIUo86O
m23ofS+QwQT3xf04ZlMXvytRtC9seQXruNNz9A8kOEbUj2xQuIrjH0WLcqm9
/Le/3j/93rHVRlTh50bFH5NhYhCI8yVoJyYgDhbVhewe/8JeWF8vtII1BpQZ
2dHJq1SpWq95D6XdBjV4TXe/gaz7BjDK5QwJln19BARuJUM7qVVulXk3W0PA
hClPG1e/nDx6e4rLNRU7waRbeBSTaugO+mcFERriZt7jz/FxP8fYqwbYbNnq
LOSn4RleLnJ0BClVov47badImYCKTBuGfYTdg7+3B9BO8e2ukLkVcH5RHxx7
2T67cWK+1cnUH7ZCQ/xKGW24bDB8Cd9ULBSCJfxY4UQEfjtkvt08AY+nj2qN
qAXI+9XJjqwYd2whvGjFOfIhTFdL3CvejTP21p9lTqFeG+wXRXsqp86aEaZM
tsZ7qCJ9pbw/XFNHVhyapTO6TKfTAs7JKDfpK17Gj7RuEqNybIjFftkfZXW6
bNf1Nm5tZYoP2+7L03ZyafTZpXvgQOf6+jHw/wOnMWWXhWQ1MUC7taZrCDh0
uDW+cBtkD/Q9mc6ChObgc61jbqdqHM9ArrHDegjyuhoTnLqGhzCDWw48PvCR
MgIaQhVsMMXgs2yYkE2kTm/0llux/gqNYgmE8NW1qOnxnhr7FLaRV5jSFs6K
bmdZudk69fSQQCABEnSkyF2MGA7IZtmCu6mv1L9SPtVBh96Au2Q4BE9P9Bz/
0esJoh6Xt6+upkHDrzzHXsPVL2LdJ9Wv6GYl9uETaP3sBkqBM+eQu4BsiXX4
+TnJLA3PJWeR3JNhVPxK9/FYJQQdtCciCiSgfqa6JVC0DEEj+SfbKuKxR0/a
19q4wJRtDLvmBMHvbzZuysuq++Mm7DC9D15Ye6v0v9JiHTpLHkZKSis1uIxc
1UQErul2Y/dpKyiL+zE4HXhTdRirFW5jwVS9qeAwVndU6INH9e2gv+z6fuxL
6h0TgGtgjcGT/bbbS99+lW2yds9Jsdh17AqeGFioEzZlsqHFcKz/ek9kEqK6
29jPr8PyGjSVO32V7EMlq/q3Tht+xQNd6gE2wuEWLgFgDfU0raAHJve5qcm6
/DaDalgV7cfCYxqqMoXF9e8eNNGAYdyGmEP3f/bGUNW0pK1KaKh4zAGogLP4
JFPeBLBq5ujJ1tM3Ay1qAM7dvRL+DcfPSjgVLUZGirXZtsK9Kg5U5JeO1DdB
azJWqddxAVNzeGLW6R6/SfpgGHrE5nPKhsuq5SbkeNw/3eT/i9egb7m8nBuQ
3mpLUAmGu0BAByVbVq4xgT3wflxzTP29yULkN1tnwMnZdIn9IloGCAFkz65W
bVZ0BZbfkjMGVUg9LeGCFeQepoNLxF5ODf6JHkmKgIqDu+GUv+v+dfgqHMyi
C8WivmI7YYid5S9+zhko7RllZGMGILGepuJesUr5enMgHf/7bepg1pVThajO
DQ4tsGfCUbeKUWqeNhLKyKEABpNPPpvHpBMTpMMFLxLOfG7hYRZv5k2CQY7M
HwejCcL5PNpO8ccgbqzcLc789yxfQ8In62NtLpsPyGEsGv5v8JEb5sqbWw3o
Ahzxi+pTdxY8jlo3fqflIQAq1VcaQiCAG1B5+ZUuSrWnAZg3E2mZaMo3YcaR
SWa+WUx3mFDZgeiEmR02+w6PFtfzkNGdBNZGuEbnLuS+qrTdzt363Ri7wpel
fCAIB/CSUBGPhDHuyoJGIjI1D2GDuhejQFdx7d22jw4jPiRSYm2zOoDrSMit
4wxsOJVj1W6FemHbAD00oKqcmAXqZnqb+qhNUZzsWtPcvk9AomY0WYAKOfW8
ly5GAxWA+DygAeNJFctNE4qT542cPNoiXjMfQGliGbbU2uVMabFyzDlnWV7K
I3Ca+R1eLcIsolh1CyI1Ci6hoeRf0xkq9BOiT1vgIrfWuY+DgRvVR8vbd524
sA6mr8HjuYoi4H2U2LLGtu5Q7NpgfAFvko9lnQs2JcH7iNpPLZlTfuPQUHVn
yi1BUI+vCCogpVhTb+x7Dmn3Bsw5/IZAccqnzVzXia2cZHtIpWdjV8Mbnj1+
ZvRMYrwmGIN1ObtcJf9T2c6P1NqKO8JHwMBMtC3jaHYJK2uKmzdZiYLNgaZG
aipX+fxqnrEpXMt/0XwXMZMwmyKIX3Yl6UWzGXC1s0RFCTdQVJx8g0Sj8yCw
VcfTkuRxhn2fFdhT4K7CEk19V8Zw2cGZabKqXtKMb2rzV/RWjNAOGtGeOhfl
vX1L0wFejWbkrQzxsVv2/MfCdygzxtK2NHGNwQ2UxTPUhkcuStPwCoIVvVQQ
AxEN02YdOK43PUbJack242TVv+Q+LS41I5zjSdL6H8X1hI6ZpB6M/VPEOaF5
ClMMr1OtD5ynz3Xob0MAlA6u+vRPsnot5Qs27dKq3A/whUM3BM4UVSp3QewI
9frUJcLsqsdV5fUePhGUzia/e7+oIiOqV6X1ONwW3xW3alIWFsR60TcS5nfG
zmejPD+px9ZpJ5hf05PKkwK6zwU+9nzMfrvF8BP6DTVZhySjjVL7kVdLJXOo
OZv+1clGkrRCzRnc+N2h7nJYJNxed+Hd9YRadYqQqWUSQpGrtp7Ll7fRil3J
p5iTIqbsjUs/lFuGdOD9uDEoP4tn4ReNQv6U+CMXLLWLc5nFuuqnau5r47UM
7LXXEDLpVpUHkJ+Gu1bXQOy+n0SVPT60F7H3DdoBXBKZ5omVyDSs9Ny4ikjw
sOFYwUsKQIcaF+VB2Ss+w6TD25rx9yO9sbzolR2pwQdDmlqap0uYGNDBwXVE
ZS1VtkNE+DiA8EKFoYJLjzIRCecFeV0dKN0Jg9AJwyS3FTBrn2OzoACwd3Ej
BHetb6s0NhE9grosj7qYttz6X/lQ3K+iYCdjwnZCxH6GDxxqbJEFVihn1Caf
cCa+24mBzbXJVZw7kzdaU75+DYLQ264C3MZ/WcCV+0cWa8dXfLHcv53+hxUK
D0wk6XVSNML9Ey432xEJf6r4oFQmOOmm1hs3IuRa8SNoUrsdSNxTcQrMWdE/
Gn/XzIVjK841GNhFq8OXdxTcH+6++m9FKP2zo6soTSpgDFgZQeeQYXWkiE8U
Si1QGV/SshcmkJSxN8eIkAKt6o/SuLL5SaBcHAWT3ptA/RNPQCgAz4uZFcpp
LfTh9c6rBLEdU5BzckwR2u81Ettu64VPf06IBO8PcC+uLhTyCxnzcze86B+D
ersd2wsRV8z+4jkNVBL4JQ9eUp4/V9X+Yhllrtj8T/YeZ3T3+uSFZNj0x0fa
/Mx5ifWfWU4Ra031RR4AOyk38d89G38ewG53Orp+qmppgT+f0bcxUNN5xy8T
xvfX8M2QzHuE90+bBZz1bdIpntBIgBdpJwFEMErDgJ71adkwk8JcelSmrpNL
Usl6ovO35t2BDa3QtfNgVFsOtXjxO1IaQnxp2ziYU8AEnmApI0JiEqBeYiGO
Ob6yybjPXpMxdP7+JbVmOICQsKKU4kWOftc3nSStbNet6WGdonGxD1pGCV/v
duI3xzB6jxXAI9QP9Nq9qJBVxxzo/XEkWBrdpyNM7RNL1rVsRHIHNFLedsb6
RDH5MVUKtEP8JfT+NdzqYEg7Gcj052e3I8VxY1EkhWIeSVKXGBYuC+cdPOZc
f44mzJEnuNIb5WblVUS0rFaxlrWeJFxkJuje/9P+iS87PIMmrl3VYbLQcISV
SeogMjIbdJLNLM391ddq0yeB0Bx+QzIUEjOAOlN7utogpfeM2jrIihl/pncf
Z8Dm9DqW+i62Yam4N+J9dMwxyG8lDS/W/8AP9TEWyCM3tRR9aG6OIQyohqmE
2ebfEKUAzhOU+W5Lwwa8FtiPbui1ytQ36zPRCgzya9XXkzNCuPJZSokyVpVz
oK4MHpuFQe47aMIuKHtDdRPLrmg8X1fLvxMRwu5Sz11ZgCBXyCHxVAkcWWEh
uMWndZDdJL7SUMF/XKjwzj9VPvAqTfN8oq3l4EC30aPjY04wy0Lo/Be+Sxz2
6yVVEVv+zOI/mnd/bK6rHfXhCa/uNrAiPCSsPfW6mou0A7e43GHffb8BgKgr
mM31ORCO5w4Yl0AOAP0Kk+9J4jWSRMOWZx5Ah5GwfygOOrePNnUqbZaORc+l
HnbvS/5UA9p24f707eURuswF6cMt/vqpmH9ONvcr/sOcDKidg7addgUabemX
TRQVSJxGwVBdI2052hik5qSSspZjhoGHY/l97/MO2fRd9Xy+bZ93073/8ZBK
/OTTKJnuDhXijioBi5J27jR0eFPflSG0uwUju+FgORx3ugvZ6Relg+9d2E1O
Q8ihch7aFQXy0kTqfd+z0x8lHw5EX1JQ2CoQ1os13f4A+0EfiovEs8VqzWEq
tS5mv24q7whnfyd52o9kwYgnrims0yJi0X7LKK4TsEYFuaimXT9AAxTxOVOb
btssBXIQ+Ga11KdXNemFZevDIyTQJyyF6FDhPWYd0nJHLjX6ANNN9eLAsqVT
TuMTiROv8rQlZQZXK6tdsjMFHZ9zCZpdVV8CCAdgf/9kLQBPP+SmfGe+Fh/B
ff5S9D0Uli2P7SAFGULPmKhxsKqmGRkEc7dIyvLmccIQkWnnm3bT8QFeAMNK
/TSiM69dWB2No0sro+yBJAEMrc3LU6M40sLPSmoW+AXnM61EdiNsoWn0f5Yy
74qixq3Y6b20SVpY+Jz55marSgMAAgpO4EBu4ahjDZo4TDGCoMJNSBXWDoq1
581LOeIiwMHicQk/JOZI2i45eUJRn26yvYvcb2FFE+3VnHzE47N1wJkJx2H9
VA+NaIC1kxZ6Ycu26y6dPyRiTVN/6O3g4A9xHGvVKI6CvHMJVXeAqvz9Lv6j
UxnJyl1303Icw3KhQZeGhneugoVcHSAHPmEZaibULEZi0JD/pbaKYghZCCcH
4Ay+k4ju/wQYTjcE3i2PSTC9I3ieQ11AoTuW+dfKTh8LeZ4xpK2Iq1Eujgvg
UNrFiuYgxNWdTCI3iqDmjlEYcZ/eduMVP+xz0jGx5HZNbeXSMvMf+lM/1Y/8
PjIoIZJ83zHM9F/pUL46zuHYSxM42S+dM01xdWtiG9VaQl0gZFKQIHtr8HA4
mWooJKBkN8p5RtV4+CcbAm3Jiak4Hs6ljlIumI8E4tYx0OpZzkS7EFaFPAGh
CDb3BXsguic3CharHXYSHr9ALbERccB14LZjKLsnqNRKP9uP7B+yKzL3291b
ummH1J/wWu+kuzFuiibvuvWNJ6ojcHsvH2fNaojna5FkRPx88eFt828kLuPB
/G+GBRV5lEt4NgDkQqs6P39vAlefRFqqroPZAwEt4Cec0T4RA3H34SlbR8HI
caJ4/jzMSBwwQh9rBhEjMHRAxE+QjNdWm49Ie99z20FbX7OZZwrJM8MkAAWC
a2ff/keyHrM4bMpVMlKAkmgVhA2jGfOe0Np2uxYdsnwDaN0lbHfGOZafkS8j
+T2x5/qPswx3Tppuhsbh5z2NsVU++EiBmzu6I8fD/PFRtQu6RfroDnnNJVPn
yenvznBqxltlbQflf56RkXpwT/22tH4xBjfMLTzOGnd3W+wcYyVCgnZpPPTe
qeJ2dx4cjHVwcdLhAaMXWpFnRXcAd3Y5NT5NzeLbsdOUvnk+BFCevZ1a/wWB
2Z4r/WmOZuUhgJBi92Zm//kM+YCWRpst4+4h6SjU1dgwfFj9E3GaAQRZP6gf
/MFow9A/6N6HOGdq5lQn7lseBZiJ5IjUxt8l/f8PPME4UUg0q5whJMTWA2ni
VOHv/6zUuHbcu11FDD8e1fUETYvMP2+UJpuB4AFDawK0vHWRK3LF/5aN77ex
YD8YXzL+RKWvvk3Po4/mS4Demd0r5Nz3SVOw7wsxuC7AYtF5P8pIqxgabAyS
dK4PT68tvFSqeqm1Rok3QQDhzKPtfVbZMH2LxZrv+/Rj7rWBrw7Zo5mjN8Eq
ns9yFcJ9n8SJLwFj7HBYg2peFJXAbhOv3rNlhdr9hCyjM+I1qenFdEH89v++
iNIMx0s4p0l6BfKGOILkV2AEOCjf2Bd1fdzmNQRQFRzVLTG2s1llewt0KWC8
9vViOX3y6aqRKdTa0FrAK7K53T/jBtxNkdbW8D/Rn96Xnv1fEKFKkeAGcwr/
IqAW1znfI6xztL6rqEacd99OrgZji7pnK2iVNwAs+FXltxa2cN6Zv45ro2p0
vHjpqsrnqxNi+Bpq7wQsZPIoVDsrWSo+toSdEEdSL6wbwHoDfOfGDEcETLtP
ABkG9KC8jAAdoF0Fznkv0sxGqZdqjA2YSSzs89MqlT/IaHG3C3b5US9g6IrT
Ui5Qb7Tw1YVYGcaKD4Q8N6VtFKSolUPIbM/w0v4QkwaXt2CNXRiREmOhDHlW
7/TKT9QLjWNwwTxPJ72ZPj7yQCZDyJfySwi1Abmi0axp8SshHMPk/dO9AGm5
bvLoZcFzUVJYFGHb1xNUzU+REBf/UPIJ8v6pU/lbFT3cD+YZnOfJu3g2SJ3l
oFtZzOwwgwpaAzb1eKtGWP0L5yMfz8dkJA686dUbCRsLcU1kLq1r+ArsWrVN
NIaqKT6Iq+YwVZbRBVtDpZ+5jQnt0Utc7yz9s73MsqYA9UIOiU05kqQGCLAy
BgB0P9WWw0B6YcDTdTiIzjWuo124uqbdERKQGzTDqXNYP1rACXGNKKUuowWu
tr42fDWKIpDR0Xh9PDUrxpXOC63oDAln6orgYY89y2+yn1ImW+t/avVYQ0b7
g0vZFmDdqgNbbwlwx3SllPGC4TBv/bOdkFoRGpWzPwv9QASLy0c+yYzlHDYy
j008DwIIf69/q8UKqau202AIMlZMhKKgEoSdyZmI405AdyjyNxrl2JtBYhIO
gHlmIIvjbq3mtr4jciOEdBFmpMx2U2lRfR/kybgolzdtrCjI6UjDZEWycKQY
Fhg6lHcjT0jcQb+MMP8cQTM7A7KorIEmIu2CXVARPXGPTbqXAqj/K/QE3kxG
t0MmBjR8SVlaAClbnKqHN9IOW8vAnilmheR/69EHkF1yUqqBReQdFyvuAvK2
ZuC39hvXSPtmXap/oOPqWF9NGYCcegrT1Ktr3CNKRcloxEDqgZ9f9IomgqLh
/7BgCjRKEfdWCd0W0SywYJKxmeyHlhRNMDNVNW2Vq7OHJBjYHGRAd/y3Pl2a
49yPpMSHxmIhLnYP1FdU3znPUFmzSNVFzGWxr3YXnlnISS8yE9ghDLzfsABv
bihUqyeOgaZxhhz2SPzzwLUqzL083gHg243VLPsA70iW9ck3+rLOjXRn9U51
224u6ccf84+uK2tW8HXeMCGEPMuFgX/WHPWoUlOqdDK/z6EZz6U9RP0x/lLR
uF5ZnnL5nXucNBKiEBbZwZhpW7XksXqZZL9KS5VSCAbkBNhdpvOZrwT6jyKB
mTPE3P0aDUx/E+8mSzb26PwoWomNa8HKqNIRBLLNkwUd7w1bkEIZJcP8JawQ
YBmpJR3xW63xXY90in4jjc9glwVWOFMsEPI1wgqkVm9bm1OS2w/IfgzyugOq
9A8hi6LiX6O3q7/mTE7tHb80RE+sDAFV7+y0v8yRjh2N9uyuvCHFqAOjhwR9
qwlzEIsWoxoYAjUMpOEUzuAH5KiBj4czAxh7aCO3GfmIolo9gybWbT+4LGaR
oqbLuG4uqvg3WvHJAm6Yk55mEvEOUoXbgZZ02UtY0pVUbLuzmZdSG8zZ+lL/
YQ29qUGkBgvq/V4Z/1q4nGlsAQHfLWvdv5tPsAM1UROitE3YU+faf6rX1Ezl
akITECMFL9t6NLdiR+LmZ05zCOxQrqZI62cuZELwNiUHaSMIqMtLkIx2nUQD
QIlyjt8X993wWzL687Ton4yzus4edsCmL/L8OggpFLWf/Eo05W+TiWXsuDP6
AB9gfntIAfTAQiN5dwdvWQfeh4tQrZoWqN/bVFbFcH95id/vz7EJZDOj+4z/
HNd3yhynG68uOTH9LPmU9mRKhrmvak9pwLJxhbpqMps1DNt6LNXvnO+pgHbl
9MJGizex4oQBUROkZQO0i+GTFQIWqxjRpMlA7LT8NPAj4lJVaxPc8Wfi9K1v
l0gp6fXKqADnyNeukQ316sxaSfuniECToRfHal3ErNDNmIh4Na5gHTT5H3+G
OCXyJ6sXPKHTR/yH0IqFjc6zH7CcXt0XsIyCl1SIIZ+sHMoYqNEBVi9+A2rp
G4gdNMk4lMT1lzE5Bsio7jn18sq86FjMUQaacZRbEpz8LAeFuODQ1e5bJn3D
GJuTHdUGNzBvGhif5l+t2iehw3xnWIDUbU0GTPUvDq2V/cZ3+fXWCvS9LT+B
Hk0T78TjsHcI1frf+S4daQp/O+wXOJdSHfuERZ6mKIw1ERqroBkK7LpxzdpH
soT4XyymS8jSWJRcqR7c2QoodFr+ElJDa/bIcybEADXotchJA5sF0pFeGsin
60e492HoPCvNlopF0QEEBMfpxR+tM9j/uDXJGHEPty0I8p3/wKxxWAIqYh/u
ib4xuR2w0kwVh4j+n9WfzWzd+XMiuSb0FdjhQI5f9dfQQng6WZ9UEZbfi5TG
12VkGLxrbHST8h8SNZfLQs5Np0qljG2cADVukurcRgqaxF8qfY8f5n82FgqY
84h5StTjk58d8AiXvRVWDTp3RRG5++r0XYmZgA0ip+jfA2uc7x7yis7CwS0K
zAq2IKK23yDZMj54OSZKmDvrlLaCELByaYvFALppk4XA2+1wkawnGWY3gdf5
qmDCieTh7vMJpZzSw9RxIPhiX1aRayhCQvRsEMiqX3GyLLIUL/y0Pbj2vbHo
YeO6hXScY4GNfhe7DFxlOJEQcp9kdF9B4YoEHOblp6HTru6cwpxLRabe+6if
CVq6gQ/F4FdsJ0098UxpkuJQWepI3+8fWWSY1mz0OCAcZyfrEbgU+SdyBJj/
wdKEX8OxDB6xgYzIBt8APGoXzGJNDm+bPmJnvH2DG69/rBA/4u3xFtz6aId2
DYg1agkVRKgN2Fw6Ln/fR/EwgNOEdqfEDh6quptoxXqFPwxQaxF4QI6diMKg
D4usfKcUniEFjeXVxumZQVT8zFm8tz9g8a1gDrawvSMAR1DdB0kwco6zzA6q
c6CdUPOL5Kk2MIEtyb5pzveVoI6sllH7GDUVSzuRF1PmrDPOPkKqcoXqO7/5
wmUUk4tNqQ/QteAwUQ/3dbVUPN459dWF6GVp6NAb3QsQ4pSsjBMBqHHVnN6E
Hy7P+39WGHgoKtZwt4O15i0YA4cZ32kr+YPtCH8hlSCXYtBuzqqmhl05l1KB
udJgBzQt3v3XJJDDFtS6JCz7hBKuF7zBwdIR71xt5/9iczgy8Zl6qUf0eQ2I
jIOYywNB1zkvro2SBBh0AFxiYtN4/I4RzDQqFXMGZFf2dPw7hGbKYCialVOm
vJ1b4mIqkcEG3hNU75x8+TWLiue5MBUvY0Dd1Q96FLHDZVr5+6x3OiMyWCjr
gPoKQP5XnlBTLzn2J2/Ak2qaYIjcFS9py/ofMpaSBw105Y5D096ncSpSG/Mg
ukUKZ+rsmiKnuDCwCfVZwIVg/Byv1UB3aPXFALjzIxSDgoeIhtgVdngrz6Ng
ufgip7SOmwE7QWmi5arjDaD551JsKRHAAHH2svZHiWE9JZzNZj9UIKeVvL5R
cEDyKf7MhI2t3k6boqp+8SEczv4iQ552PInwMdbYtXwuDdGxVW62rNSoG2sn
HF9EkdSllZ5kXaApjQHeMF3XSWPs4dY36FpRyh/weRSCJgBEdX5Yv2DQxQzq
hWiwJIfLhBV6V8l7K5aXM0xCZv+8hzRuYdo8zENssKN+XP6vcNRyhixQWy8s
/Sdi2RcqdVNSo1/AhQYoZAFRS9vmABXtwCSmcmoAMS/RbxpQ3X8ISwulQaL9
sCwPdw7jk80GLfl8U+6SvtyfXNbQ4iSoxpZCbJFNol3CTf04QlRTy7GB8Cgb
sHBy8rQTdQS1QSQqWt2v9zxI9UCHFyC/DEaHqXUP6/vGl+6gbpGdZNWKiKkz
hqoOhoHO6oxS9DapeAqMOmALBhSymry+AHU870b8JidyrrRCHoUEWJKQ62C2
r+f1aKvXKDQHgUwCjjc6H4T97B/Qgs6x1ZBi306niNQPgGlX4ywm2olpWx3h
PPXteJNoERXIrDfQEVb+ntwJmMIKUIsCkpgRaIzotMbNgjaR1Fnn6sO2UTuF
IOKQyrh/BAIsWmUxSS1wWHbDxezQ0Bm06/KLRDWDuiUlJO6A4AIvS97ZVhJJ
S191U3LSOkXcHz6/YZokalOR6+PcXDHlSppJW8E4DglYj3AUWpbyDRwGWoKD
N9UcCMDDF7l9WTQ3Mv8MgitmPvP+8WhPu9y2nt0ZzMYJR+BwYV6q7qIoyZ5w
3RPOSUOr1fe0mL4MTWsztRe1nVDQ66AhyrAXqZ5ttfTMOebE2hmTN+bgnTQx
PEg1vaaPussWKps9Op9uAsbYvQWcnte3ckAXJ5VLRbC0N+tX0sWnklFINEEc
tXUDRGfdPp8zB3XrGnd+6ITQoBmCqENEVe35+keV6J7aIahAcb1V1UZRPurf
CnI9KTnMxKGxdHi9Zsmm6SgW3sR2+wH/P0G3BDKMQfaFp3YbWvMFs0CkDgS6
iBrzSheZrDeYurZU5m4/WKGzPNTMSc9NfRyIyt8DGTgEykEY+4mLqWSycAR4
a0djX7rL7rJL30oIs5h4E469U2uTz6VhF4awY6jXZbX9qUJXk5D2MX6lCcdY
Fd8UgA55oQKFKyDm3NEDD0sfLBMqO1puvcTvRNWI0awwQiFCjbLgjHjPt1Gs
yCuwMbJ05lkk0jZIdZrti6vGbZuwX5u3ghOEy3EjVuhAlnPgzgtHMlT9W347
rT3s6NcTQRvXVAfccnx5ZuXTUKOQWL5pdwjAeplAUi2KFXcJd+maDD63tJ6R
BAISfnJcFd5bmGJjALRbepTnJ74EJHbtp65lkFGFCOJkUlUIN50K8sDb9M7W
OVBAjWvXvpyVZ2nED7QWw1G54nBBlK8+1Ms1bRS4Y1ZWwxH82ozaAb/1JFl3
sv6XEoMGwC1ax+St8Xm6oIw5oF5pqFzi5pl+xhQCJDNFWe2UuyYCMmxc66es
FmwMZZlNKJXoGI/5x+ApYbatO76FkwWovsNK3Z+eogz2VwT50WB1Kv03xYBV
GoTaudUJ4PsJSL15f3XkRxjiGkwF8U94LveVLTGhM3PQTNgKYmGPoeZpJg7Q
y+9EOj+0Dsg9HodOONnJ4KwTFNbwL6U+q+APMP0KWazVNBkg5ULe/2i4IgBC
mfZpkpkV5XpVsquwub0d4u0mrUiHJZPcw1VdTd8N/oaVLHgjw6gB9SfbzHpB
V+DT0zaVxc81oWGwF0buZNVWS3C+G8b6mXu9rGR5fNyztQ1qtuF57yJg+5Na
r5DLHaNyA0p5m2KJXK+X/94JLmVg2zaB6XWv22MIPxY22Fm/8ULC0DzHmgke
dTGnO2DcwBLCf6NqTNCXKGr8gI1BLuJTtyfqrs84Tk/17Z9b0DNhzToUDwQ6
E2bTAISkSPErN0meCApC5R7EtVajx9xpDPhUXON+RP5cOHvK4mGTRZXoBl6E
TLuFepuwJnRT/enqL9os4ZmYIFnGTiPR1tlntU8/ErIj8F/NCovR9qOfQtqR
D9n2hwVBv62lVB/PxNr9/OBrVKfw4YMFGEE6pHwznkTTmfVYjwnydWDAWGNi
XeojK70sOp3yVLTMZNXDuM+qt/35JX/0Qpyt9TEpiNOnpsP2i7S17M7QZM1e
pE/sd9YGoVYKxJ6hYMxA4IG87xDIn0NC4rPEmlNbRDWty6qmtTzfZ6V+pnDh
nJNb5t0CVQjQrxpb7+VnWySQnVybkOjdfxFhvLhUtVonOyy3CPkqi/47W68r
7vao9Y8Y8xM9aPUp6Ck0Pv1wXlLHa7KYq9Eb7LHvaRssthMXBF+YJAPl1Mp3
4e7NUOSArZAcgoQcwcRY08MfB8nGAhNYy3j3+iyqG8b8I4QOq5qs/ha6ikhJ
Uc66cSQLhqM2cxWSllBl+S1R/0RgEIeOt+xj0BLZ71j7Vi2I0YwrKtSwQ+87
q7TPXQK18N4MTj0M/+4JiKEp2Tra7DKk02YmqEyIk0viTNBsy1is21d84GlI
Xj554ufgiz7fVEPwvzeMf5GAWcLBtKBD5gyg8LOJ6qS+cikusgCB3gMseOy0
YZkc2B0Iq7Vym2XS0oFQPn5/6tPhqnz/0z2PC0K46/pnl4JS5u8vtOD0s7Sn
yeZiOxdro5ts3EgdNR+kc3Ls4PgvvOdtuXRj9LM64cyP8Zbatj/rpr2LD7GM
NyuktvSxVhKbkHxGIVa1Col9thXc+NiSVQT7U/HhF3BtUTCIhiWc3VlqQqqZ
ZOoYGUo/8NFx/etDdiCfeHtEs+Pmn8gol0Dz4GyX72dTIw3ykIFB5LtA9ehU
l2Ux4OFD+YftDbrn+xbMwocqI2VgRuT6OoSsmdDenuHseKT7aBuZgIwvs5AY
qk4iWalleWcZGC51o7XpRQzMM7hrrbmEqWqv8kVSdcnEyv9KNPmpy2mcPypP
Ipe8Q0WX3xkidrj33VWw7dwh5LQJOetox6qcdMMX0g5NUgHUiImcWSgIEY2i
f5WXJxSMYSLe/e7d+T1pffthe3aJXtTw+fv1rdDBgrkS26TRCpNgfoPy+Qw6
7JtvMqFux0rL4hcZNa2RbbqWLJ3/LGNaIAwpUgSE7l25zAwThadLtfKpGUb7
OtdhqgCfIyZ7F/uUtZZx4roog1vecWYB/T9gjICtAcMdrg4rlkiOnODc/0Ez
1OTJH4MIyeMZJq5u1HoAbsBF/5MQXUTq8jqK8gwKMXgVCu33+vX04Dm48lac
QV1rl1lii1BZ9jpduKmU5NslKQUDQDIINfbLw5rvah7EDMrxJ5DkqITuNU0x
bgWkKXzLSyFyxi6ZMYp6EF8kzcE1sqU98ZCFfExR0qx8QYn9ujfKRpVXR7pz
IMD55LNi+QEHV8F61/WPBpt7tg3B+Q5MYVIuplDeUlCtqJJwSVUEU0JEabrO
jdaMdn6IRi9oZsX4QB7myGZKiu1RN48ciZeEJZQZlfgv6S/nsStSzuidsjKr
o87c41eRvIBfcAlYKVn3v0xx88Cqkz2RdjX1xWM5C0GBShaKRVL+WS+qVrGi
IfAjuTo8VVvlyhokdRdDTBeHtfo20a5UzJ6k2+P6ElCCt0RalVzc30yx7jIR
Bnc5gDDQ1UdB+/E2Xpszf7tZPFakUhM7y8GTI1+HXng3X98dttDjFcNUo9vx
JxA1KL6/E3DFhlSUyysh12BFkuS12FwIZSRSXYo9aQZbxyS2wt7b9pM0os+/
Ly6KYpFrunxH7ERvwbx4oFGqOE5c1+xboxHYhBMwKP/TXYIYs4VzmD1WjYBE
QrhR6LVBgfEdn2HGrZLXuw85NWfk6CeFjkqXjWlTgo59XgeQItGmcXlOXiRm
n/FGgBgC1Ip5PP3c4pE6Pgqf9OVlM27mAbl9Maic5UrBMXjeZJL2wlVNh75e
S9SLndlFaBd8MhiCo4gIMOMiB6C+IOgdIcAnN1n2Tl+wJfpHGufNdXSM+Z9P
KZrhU670BeuM4ofoE9k2F/ZHS1TCfSVXJsr+ODDicdBXHPrRbXgQHnsgubcP
XQ1jJLsfIZzgeyJdMSaL+D2j4tTOdw51cb5/cyTfvExk7LOM4W9ZDWL4wO8+
VIh38/wJt2ZCi3/aVLON0a/Cnx26w+/dyeIu8ZEJECTrYaARHRUY8cc2wRu8
PVMHQ2IKqx6JWCKOru8Woo8PdYJT2TFeO9s9cRpNEWzVDhNwCHzNfSTlDgmW
HCeeynqiJdR9LuANrBdi0Qa/V0dsLsltSa/rv7bZxfJb8tKtpq7PID9FDc16
iaeEGW8IHkepGvdrmijG2/Y9Qwtx2kiCJHSuoHErcpvc/MdU59YBsnyVq5ef
w40xAR6SRh9WrOzs0anBwfFVjg1uhqw+zLg5Ffl2kNyR6ZS3pVRm/ATndAwP
bk5vEdBpuC9GIuz/m/2vzJpuoLtbs49MhjPCfoFRtpUjFn1xvFwYVa1ph3Ql
g76jCisx/VKBQNWzkDaEFVfRJzYDit+2Qt+PaRnWL/oXTkARcA+kNFqtMtFV
clgu6KDcHMSNyRmaXcbh1c10fpsKALs0nxmcYuEmWslAJxNOgiURGj8V3Lxu
NVP1Sb3ZogKEu699FR+hAt3SqaN5/+jZxRw/NA1ljgT8hf2gOuBQhie8wTN7
6e/zbpUHkTX2AkUuTQUzlY2rQRBRkdO0J13z6fI4clVNcYjDgsJGaaUPUaOG
HtmmEgTTcWJegDd+//pV4E38Xvz30yOrAkQ4F2qBQTfBFkgfsuxRHpVYQrmp
aIdm3DJh34FB2GeBZXDJEt1SSwWJQPrkkZjsJvBkXc8s7gn4c+iy8q0InJLi
t8hBOnN5TI3Z1u6Hy94YwqWjOw7hrYhr1vL7fMPXBSgQ0zDVD3vqyN6J2y/d
1wnX1FT9lpCLju5U8l5EcvZHPZmNL1oWJ5iz7tCPkLErSSxwnhPLKdW/D69z
VU45Hxh2Le1duAsoFwaKvMEuT6g1Q66MdydXABiq3c5R6iJ84UdMvHmhSbUq
Xo0yEgiXjNH4+6Os6NMD+WlCnxzwPtIfBLw5YtcYWQJ1NUhoJXjPfxzT7BNT
jM/3XUzGDi0vFK3k/SmXKAg+f6Bd45DTGi09P6K/RcaCqNBoUV2kYdPKjWJo
67K/UawFvinclPeqS7P/lFO1i8DvEVjKMFHVwVR/Aq6lQEHug17Fw36gy7Ew
J91mGe/J2giWqRBIvgocuNrnxIUixr5wj1LXHppNarMgIxqjc6/3Qktqosfc
pOVS0lBKi4IB8Mhz+OX9aQqULf5FipnxtecUqdZdcfd1YpuwWRu7qOP9d+Pg
qM94QGcpGhoypR3J7V4eLNpVf/QlvJnzb/C/Io7rRK0xae8Nri9Wa/6vH2tl
9grRxHurZb/BDfLgZileYVHVvS8Lk/1nL6auzTxDLoFIICNejpShafS1wdav
qfER4MAQnYvGfD362ujzndxu5USMubnBa3s/DMGY9CqHUHZB/udoJmHayh2Q
dVl9eHjB3HFpOrdi7HrDM3JpQHec14ssyL4DJb2ibfl8ACll79XG9rULQ1fE
yfJfF6jZfx3vMxlxtM6esAMW+zAeTOvb/yvCxZbmsO4sJl25V9KPGOKb3a5o
vL4lsnwLobnHq+a+tXKbLsjHQ1PT2CqrhhnvtA0z+pccDbONC15CdaLV2HC2
oItNrFbFQ4IVHSgSchF+BX9g+uycdiWCdt/YX8SZUTDOSzEfZQT+4SyCjspN
FI6upyBJRYQmyLsy/VeZ6WHfKksEqpB35Qstgh/l21NvQ7i0DpfrnpfVRafl
SPE6s6y82RVj4qL50JaYIaYzDxz9nfszz2BDeoosFeyJG7Vt+WCC//7Owwx4
LvhlAUpRdN8imFS8S09F92ry+rdFGQ1Np2IGgDhqo5RvB4yIy/jOjKkXA1g0
nLSyJK30XaZO+mzG8IfSY5vWZxTk7NpBCMrG7GrN2BXk+JMTSau6vlNgIxf7
X5jZwPK2JU2VTSrePMK+XUvAtkGGEAIMp3wfg8NSG5WtIrPyKDzQitYdTHIa
UEXDobG0FZfjI9vtDa3ppR11fehit7tuYJCYKkHvs1flZMoqKwVR8D4uj+u2
AV+CjfTks9upKdLVOuWdn7RnTZG4v9scQvrGD9TwRLQKdEbS9QgDAwdDPb1W
Qb1RuO9lpFRbhgzqYtGbW+ZhcEq35jNMU1d/whjnvF9ZhtFTJKL32+FD58ur
x9Paq5Bq5meVJEKHEBvlsknXpJ0RoVwFs3xmntJRQKk1mW0EN2w5qBO6PlQK
BSbn+WZbLe3r1JCqTCYUdLSM7G8Afi1d3HBgTllXA7ayTmde3qMp0oHByDk6
vypU/mc+q7rY3cpCF1ueiZps6OSMjbGWdSRrW8BtHdiYa6A30bH7tPFda6EP
aCtf8RfohOXhbeUQSu901h7uvRTbXty067LbNwzNW78qQKHLHoMscv63U/Mb
ULqSfs1rCMSECMAVY7RwiyBA/PC7PumX1aCP3cXvblqTJ+80LcPE1tHHtn0c
1EDdw4A3s1/7F/nhVerNpVsHmWqqHfB497BCLxcPs1qzHJfTwoXV+lg8qUR+
X6Vt/G2kws/MpGThFbqkMV+8sPk6tL13hjTHEgO6jq++1v8oI8sb/sP6+9fI
ATHIV2Lhxs3E96H366HYSdWOs2WI3gE4lVegr+1blW8lys/VC8ZzUeFfZq4y
LEc0Ia3SYS09mzpzpFV3nGXEuNgT4WE3guX8/VhS97Ys9koS1t3D+PKDVcv7
ZQNpeOupLjar1t5lWIQmJoWVz3Xj15MpwdsmebVcUhlIcBYNnhZ8U4G/b0k/
s0vmv5QBrBKRSKtTjhHu6yEOXGHq1to+HQsKjqo7rVYgV/LblGeX8wN79Ira
hZWspdv0PQk45T85rFuIlbfh/F6SQIu350kxCS5QKHpfTPIYcbh/6P6nsrlY
nch9PnwqdaV7tXdCENZ3iKcMK0Do6OSOESQt9/f6gCX52SoAdL4UWdtucaxz
VSXgN2PoDJ7TcuoA3rWoV5AFSb9CGSrx1c2XOXWOyPM4kDVKV2AGTL15J1Jk
Wqii7zI/6dcfGPLQNIogSexTZHWyN8ebbzh8LbZPEtShwUsEVL/3d3+EjG9Z
YTeGhxxQ7PERQUrgsFcLiwitzLpEiWWkGyoOIUwjB2+Xj30brRHdjjh1UT8V
EO2b8tiJk46BVxpkQKtID2qK72dn25AKjD0hNI3CHjk2e6T9BcHKzrWfAHEW
9lUPGmoHXujavL9Xp+W6QYRX6iQb+QkhLCtHoBbUHnpm2meO9u3EPDoqU/2D
3sPuUTeB2MbyJtUSqWktEd7AkejIG6crzmpE0C6TeEsoAs3g1N46fI8/nO6R
OvPs4UIOG3JIx9yu1FZxfquM6glgaGhQsQ/aX3H4zWKpSQF9MPDR9yTMqGN7
KLLz0lSD00E97jeyXdFO/S8jHKM0ttglAPR6REjOP6hQuhI6l4cmlhzbsGV3
kVsoC1i+tjGFq5/Nc5irZQ0zPLNrtmBx6jBELNKt94me7IVQiO/sxA5mquT1
J6dCPi0NV7uO1jN5xwNLogyJSb2UOB516fsSMw1H2EVUp4LENXSguRJj3MJN
1688++RdSr5/ydufHiIttGbjGHLrQXTfw9NVSJEhjFb1lcBPHCqEMPTkM2CH
zHZt9PPxbby4tFlzpXbWSHdNU0civejLuZ22AvY3KxKc7vHcB1Oaz/bnbS2L
IlfHjRzasXyrTWU12f6P3DIRiQnOfCUFcTQJVCVgGE+Is6eTsPh63moxDSDu
0PpBV9YwbTElNkC3tHAC+8jlDE9xv3PZMA53gknLUyhDtikd/5yFC/kTbbiY
dd1uEvmF3erkfz4Khudgx6iCa4vW0AjW9Eip15I9w/XSmWsjpUm/fuC26q0G
87f0sSBknN6xqbv6Ntbe26jpOCDJrkuyAV2nYsbkHB08zQJfOrbHpmwHr6+J
aASc+dFiJqAGvFqkpbJUYqa+7z+/VUdqypTLEgYYsPIczGevEptLUS4P7cNo
MRDiJ82cHWiflMeSlme9HKzYsKpW/sTn1IA2IwOgRqMeG1HLw9bbXCmQFn4R
n2z+kn8ff2x7Bksa7eRV/Ty2jw0aAN7tgviTcNV5rSXBReeqg7IpsWiTsdET
/b8oT4QWVM4Zu8v4UwKXxAMdhtsZgmLuEMkRyFVnn3wBwbTVMd6VH/VLpwY/
ZiOx1Tg6jVacwfNFkRln7S9L8C9snx1mYsaUsmBbXyjO09la3giiihWeMqMK
OLL5riD4CnDMtyMkkkhWJnu5J+91eGrSuM6piuA8arR3FR3pcXmbcQNhcqnQ
g94YQ0bDATKyI96pgazohG52t98t2mgOpLB4rgu6zh7/vRkFCMRHQxbva3+O
9hHRHP1G2KVR3x7hHU7iqU0wTp087QPUWDd0AhQulPwxuy7rJjcXrb3DLNhW
AXyBoRY9+G1yaHV+qPznCV6/Wz/2EWuIYrc9y6BVloCzz4GRQnDQu+AwMMHx
XkpJ1pS2V6oqa2fE7kspNSAH9vr7zB3z3ZcJZ6Ym0SJS2vR/abS0F8pviKW+
oV+z3dpvn3Q2okH60BtF+3Bd5z6VH5Ni8lgcykWMVDIyAMzTA36QU0a2YfVj
jBpC3xXP3/IxUroUmliNkJ/xAuqFjFEkqCQz6XLRspnIMF2mGcvjvioaA3kS
LHpj1p1bo94829/T9qTsj5FZJNJdDDFXG1H/S7t24KR1pt7feP8nsmp37EfV
gZYs8GW5U07/XINuJLkE3DDNzbGudLcdM4x2By+xmnXQbHXjO14VqmClYXRn
AhNBxbuYuwGEyZ3XUPHgrTUMyuAb3QVB3JWBuTYg7/ib/vNZEmKoyI2iCRbJ
fyuHCAyg6psrVjHGE3kYfIDvMY+WA6G6Ao23Z2i8wiK2+jIIWk1cl1D5xxLY
SJq/INPdI1jyyHKnQJ5R1+UHerVDyBbFfZ8FNf1Cwtzj0PYyoomDNf1nxjcu
kneMkKar6ldwyf1WuTDz6BxoEPEwZWVmplwpS9yUcDRlqU+E30LTrfJ9TVPH
4tNxQCva+ESJPZYLZzhHj0oICHLS0ti+aFMfIWTnMFz3dcsRv1AIvyWO+aff
sHc1BAthfmaV6XQDAZBJk6pZG3/2tfmzxBOlmUlNjHZ7S9cb0RsARttP1BHv
jdD41VGTSIaK04AtOIp9GCHZE2z/2n0UcZExdfyu24wIta53QFpbe3cpwTQZ
6xpuEVH9dPrq+BW2ZYGNu/ktt/l9Milc1/nWOi0OerIDr1ukMmKUCzwXC3OC
j4pMoBDYFOy2IJyheoCTvUiZ6D3ulJnQvP5DrEHPJJ3r6FBnS0EhuN1SZZWx
lk2oWoELPU3Zma3KSnfzvHxDEcJslLqaskV/qI6EnPkdit/dxWl/m1LDkFBJ
TiJ0DHhwwa+EbIC9r1saQCVRKZh+PTCEaenGhVXwTRJigutLzfV4ZdAQNGt9
1MHGLt/70Mr+ExABtBF1PFEL3RPdYiR+2aOebdveogB+jSkU7j2B/P6uj7MU
ZOc7N3CQPYRc+JGbjZyotbVYDh0BvzRIyjlt/PQcnn1Jx4bpySf2qgJe4ZZm
lQA44XfaxF7fIl9Uwy2WuRPdcu1FO9GeKChYTN0E0MLg8LrnWpdwi+qeM8Rk
oBVQMVI41n6mRx7BhQmWAgOBfmwPwqCGURJd8leazUhYPGpFGwRXZe/APAg+
XMAy0s5tLADolQscxtmp8AdvdTesUF3hS0/1B7GNeD5GRW6ODg/le8BbJojo
NKakR/q3pH5HHItwHNTO+OI0YC3YCUVBtL1w36ZO415rGvAM4AcliksMRhF6
pO6NIS4l+iIcztE/gVTe1FoDUXI2q4trSnMOG0JV/4Jm/+onY5Z6O3NP/X92
PmdgxKkoqHm9k5BQjIpPV+uWHISK2mokEIpUz78iK3hSZQ7zUvTa9kya8Xzo
y/bo+/UyJEmogwkXXuuGct2KnXBdHwNO6sBe9zgZTIUm30NKHrtycUc13kg5
0u6Ioj3qNGfXxzpakoqvD04bUjqnA3LeeeIdTTuzGrFZm4pyg7W8tX16lig9
u4GpZmXwsr14C1r6kD1ftd/M97zYqnbRovRA6jzz+pS2xogi/xADBTzztgWJ
zh884hUuSC4bv45tyriBvWFBp6aX9bTbw131MHGASoZCqm67mggS5oDNhm9o
XI2EtsvoPkGslzhj+3jL+m/AVVg9m8axxUAlCyO3oCFKR5yv/N073Vpv5mAu
KFNeSo9f1eUXrIxthj4iNCHtkyCWSEyoff9UgrKwlSLSyJGGBg2ugodwPgc6
+4dYQU5TWJj/hua4CXomHpfTGlo9JI2SPdwQZKbHXHCekSM0UONIruZ8GtMv
Sil+6ckxVtp3X1VCNfX5Rfh8zAB5EaGFekwKaIQEvnWLUvVJtjpCR8UvOd85
9zyGboE06NcNXlFtElgBXiQ2ufpa03dLRDJxv3J+IfICuzsdispdLAvlSdYI
f9s2ruYpEW3fr2kQVHfc9CluAV0fjNT2LAMlN0FDc9ex6zBEudoIYo1xFd/S
j/ZNFshHxStu37+tX7PGVYb41c7py9T8HiucJGRWyf5KrfrsBk6idm/xJa7S
5k9fNGsVqkwbcz7IHDL9ct2NyCvNXHOB13BFa2xn0AThdeKhRutUh1EbZ1dj
Ko8/O0NJA2Gvw4nwNqxvTEWChafUNgoeejgeiI+70REwDL9v5UkGmojreNNV
u5PKsQN84woVzlAjLtR4sRZZgSPN9TGLntvlcKlnK873UPZqH6cdYd2QVKZv
3vL5KDCRARgeq37NTray7ro0EJ27mNeCpmBlchbGS54mwbeUcAJ62Kxa8MNz
dUvg2fOGwJkUyA8ykDOsG6ER36TK9rRiFE87L22N9bx0R3fBAgnloPlJREax
kwOUPpyJZtc3rdTPDZch4fEgPftx99rufBUlRqBKL4ViBLyra4CQcGBv8jop
22QIA1qgyfAPsmvNKR/XF/qhPCCEXwbIs70rBt27BgqX62jPb/75jBPKFRYi
k8btZQr05TR/1buKAN/X9dpWUVkiMDpvOBu5O0glGjNe8HPzZQL6OgZ3KFvw
hKF78PePninvpI7DvP7CeNnelofz3kAn3I5eMbsM2KGqA8dmHK9acLKj50NS
SA4tyRvT1sMtgOxeOSMlc0PVUQtxWWt0Ij27cQUwvLSHW+2MaO2OnN8bMuZ5
01odiRRJg7CPgYsrFr7iXrkq6d9OUUVZXz3o3cxKbfNas5IKeH6wJJoDvnvN
0UzZpS4mpu50hhN6iwo6el1y19YQvofIuWw1MTvnidancCB+LDMg62pJVeA4
fwWUbUHQNcPCRvxM6XDpkLOxaV6/pFuli279+GdcIf9rFksBO1nz58sBwuzO
djS6yg61aQ/24z/p690aOKXptRdJBpDIjDRsv8lY8QLnnqo1wOmW78OYpAMd
uWO0p/Vr/0ciNWHaz3W/gM9bZCIPXSxxjskApV1xb0TcX/Sy6G9CQRvcVZzL
1FPfvr4aDMxYv8hsL9CszWJpFOIcjbVdOtvA33XCR3WxPCdZO4u0zFvV9ByE
rJbt5RRf0GprLXisTSxra4lvhJnUZJC7FP60Qft4X7h+3cVq+lJwZUK/zI0i
IGG57/Chu1ZmUxzBNmRhgjJ59oQMtXkbwwC18Z4lm+DyvXW3yLI8FNZGu1k4
u1UjXkISgmVJ7KbnCE6QIfw7uqjSB/Y+7aXRa6RUTmVnpl1Q54luQ3nzp2W0
GHDds1KVIdRACwx29nTZxRaS7lJTIAsDiIBTKy2qoZx9U64ITeFbigg1gaiP
IxDUaIiuTtGRPdZyQs3jF1VKSPnSYZRpfhV1bWbZudR5i7cm3a3oL/DjYpbf
EUuL5xWylYz7H1vqMbIkoipS7zhefMtn5dYwCGnApIcdpsf6zwkvhg/m4EtU
oIUH4yGxYsjiH2JHAsqK5k6s8uF43IzQbLZ1rfm5xs8JwCrUGNpXkpak0yQI
gXngNmW1Dy0HiDRi3JPyhf0Tlo910UvYjVsXsPbL0aF2qQDiYqghA2BpYtUd
0UteSqAyf9Z8oZcspJ+9cug0WbN5KYdiMgSx3yzOktChO/cCJae8LDnD9Wrv
6cWeJbXjSAmW74faYbFUV5rBCnEDzYnIi7C/wArjXKuojkffd8WQt36WDi4P
L8gdF+QWigy1jiSWXdcch+mgYhO0Dys4FmDXFVyNetx6pJWn8977EZEeSrhl
rRPZFrsS1u2QSmtibMoaQm+FtxNsrJdc+L/j0ymUFExsocGMZ+3GwtXOdHsj
A/exzjlzcRqiEH38IUWNT8nIAMwadDHBzBye8fwQcD56Ptfw364H2NcrIdgy
YiQ1+YIXQf78i3J/I8pFY6+QmqHP7buDT+tBoxx5IJhkFZEgUvRZ2/tZhKXg
1x0FoeLLrz+GFrHSB0vaEYyumDtfXGDRF3uNWevs+c1Fw02IntA9d4ApLr8i
0n/r4wH17CSCE05uJYJ/6PirKwCqFvInS5mUFVDHZSZc0aWp5g1sllCZ03R1
B6QH3hR/ZiA0HOTIPn5fC9EYuPZIDzGy72lTBOP5iUUEpuXdQl39hHw+XSXJ
GtKjs1HH7IppDGzRA6mwVX5z1g8TmRJvCXgPn/Ow5BepA9OwQsxHVOcq8hxX
R775m6zkWaAsFNjFP/GCBHyvThssYZiQVRp+FaOAUaKpjmvYJvwdjDtQKzHq
DEWqFx81VsG6VLIZskvx2FeygExPZ6VNnkFjTjxqdnpHTTdDRzjGIcNCM1oJ
0CTJoEDULgPHgxJaUupznJZ4AI9rvyJ4Qg95CHsDcVLLFRyR/2z27j6/3lcR
COgRGLB+V0wpbSYe5xqS0SBdwFovac6wlCFzcfQ5wEXFd9H1CR0CcVRmN7IQ
3osRM41rYC/+nUkHn1PoevR8/Cn6MwSe1mRyD5Ym0LLvw1tX34871TUTHx7J
an2BDM48EhgTJPzZZouEIc5GCNmlHQRe/QochS4BDoEbTkWG6afBGSolJJte
2Nl49EyeBlp85b/OJiPcd+KfoGDCfkFugAhu6sCKeqS4PfubDnSDDC2SbNKU
BIL0MUW3FwbKTWODdeHiPS1khs5OW1LcZGBnlMRFQfLOIAuUOrtKpCmybGZJ
vTpXopXF/EbzdTKNDrpqQVrxcPJyUKswfBnkxZjsp4YIjB7Bu007bb5tAE93
t7YkavC+BGDXCuhATfcMQVu+JwitG3H9xnRy6GFmrgg0BoPbFBIjMgx1WD6X
FQK7Ld/BWm//UiOh4835rbXZ/HQigizDWZiwrB7O2EJKjpyVseY5XCg6EKmJ
IM7qgzAt4Dcwn7AsgfY5NMN6zz/BbwFWMUhOsHnoWQh9SzDiXPXlHxwL0oP6
8I4QXeDlGf3R1bfM+QUi0ZNh73FUfW0sJVhYRjZVGskZX6tG+RU4dTz72oOz
6slGZUAXqUqupSoaMy2xErhaYkgWn4pAUvwpSW7ZJgEyo1IVL4ve8bbWd3m1
l/LYbBFWq0he7asl7GnEtq5sa/VY5Dilktzs+ALI+oHRNYDWOtMiHUUpzBZ9
22mDq7thHv/OCgUVVhRZi+T7KwhgcV82A82Kf16xSfX9+DHAXJKe6CieFYPT
OvAY/XyOrcQ6pnqRAljLyE/bUeFxVbCxA1+sFhpEVLd/PyJQ/CfkIddWb1bJ
2P3P1DDXa+gWiXb4qvYHzxbR3VlobH8cQbKTswyP1GeGFNmpA+vwHTPeSm/6
018lxdGebezXpJkAdXWkr7xBh+QvRybmR/KTxtZexqd7Iw/8BPn3jw6Hck8Z
WZm46+0Orv2OlfAy2kcK69z/yuUKFUooU/wKUGtYIoVyxqROC26ziEvNIem8
/yJWkcnmUmmya3LeosD+knOk5iXyYYe8MJVyYvpiuBs8uhuFoilHc9LgKWar
aK0nEz4lZHZBUU2eebyin7C2/MzBFsleM51LkViZDFwVgGgkofV4i8TMTIJN
FIYBUzyoDlsrjJFh4y1AH7vEHLCzIvhxVAvSGR0qmNXItBaokDQDDdAlxaRy
DOmyp7kSBH4h9yzHsa2+kHvsVZINZ09RvlWxL4jLJ8EZen7uzqzMm604mIt5
81C1qjs1mIiDfxk2o1QH+xftrd/0/UzakSMe4SEhpTa/sxkvbuYKCvpmTBcT
tpC9VE4NR72y/lJq/xxHvNTJUa7Svh6z5BHmjMtb3+PrIgb4ZcO69v2Uu8Fq
egFrDxNjBoefrVMhvvkJ487EmHvpAA97Dcnrrlz41f7aVn3qVXrrwgR1dmBn
XbxiImSBxAnooAZ8Spg+ikOUSTjFlt8kf/3SrGhxvcQV23hkJJAmuGI5Ik6Q
GEvWnh3+BkkvFvONwkIae6AtHD7Q1SSErdUH6eNwBBZSQkuTylj31vV0E+xr
H3rvCN/ozUYSWKZg/YXykaiLOgcjwsgxt+wtmPbvJAzGt2y0ju/rtEGtK+ds
v5aBlZGXs0XDadutEAoxwdkajh8QC4OMLr50znpOeNwMQgERnaZyt14/HIOG
WpS5fRq/8LXzXsj0ikPW8qql1avpwPAVMON2rcxsKO3NE0W+58qWV4VeLDgE
mSPfwiGGcUmtIIF7Cn/OzVGWlOOYTpJUWd3iOxq9IFJBGl3fqAYwdxv8c/Cw
Pds9D6MfOEI7AX2tIK2gfGKR8Jx96fhC/pVdPtX9GQXv8+wfM7NSz2DPcrT8
8iErKkGKnQmNaeC20YPnfamXBiHNkEJDbRS7H+g9V4JpNqoJP4O/xdPOciR3
wMZOe34+vCFJkTt0BZUJG8O/MoGDaaGMDAFOfqkIxFYCqoLehkqnsn1B6Yri
ML/pRhzgZ2mw3icmEgpUuuaSZFUWl8hr6eTHMOBoYneW46H+vhWqBUTQWqYG
mMx1gyBefX+NLTYaoZKkHqEavHnHHM4VFFFxWuzFy55448QimEhFsgufqXYd
ZQjSjLD9s8wCBJmM6WSQW4fYRzYnyWs2OPMjDhzAKmUYGKqKst9KtBrjJCVf
hw/pPgMkzLEHbnTtJbg5NminuDfasSKCyjKdpLI+idnxY+csPzihr1pkrneh
EcqQeZgLIy3XNQ+hWz5pEDLLLUKc4h4HarrRvKEit8CfT0AOO+BCLKpgg8rZ
p67BnEsBMBPliyG6i+90t6hSpLF/f40gBBr2hMUFTO7uaKSQAKnEAD9NId6+
AJnhpi2xqI1S6NmRLdMaFTGuT+D/E1WlLyHF0BzPAqhYNPcIAZWT1tzN/Tbp
65BhrcLOgrNJmiNs89fLRtOIN6E0geif1zZQzXDiXt3A02TjYIQ4oUNLPz6F
YIPk6h+7wpFUW8jShzq90aJEGvjm9gxU9lgH74hNPYMATSZBi24IJxpMTnwc
x4zUfwYPOhW7Zluw9pBb53aGDkURIlsf5eDsBH8/oHxf+umZXanJli5/Dk6a
rmcl1eRtOZpQosS+4nySqpwTATmlyMrtfLc8zcp9xuQaP5G3C+BInWnIoREe
dXkfbxSdUZNiIufHVwhXN/ssUefRnHDjSrqUckA52ITySwW+GrVV4wPVzg2p
4sDhr13OUU4AC/UxA/XTNcqa08Xp7OduTjYKher6qCtfhcyhBHILE4G5HyPX
ljT+CRvgUjFHK+MdRmyZK2Cj6IInToaXBK+sUo61nFIExIUMRep7a+YDeCHb
WT0KlQjw3yZNmG2gECT7rqydDS01Sbe+8FdK435aOUEgsB/F7wxToVAANWzj
H08k2q3KXA++ygukZ0GGxqNwsZoYwOgH6mkgiKCquGbMdRfimx372DeSuBHN
uzZzbcaxu7ZMbsbVkhALCRJhlBkljnoSomufzaSnKEgjkTiAV8HwIEJgaYFR
jNr5o8SrBx458fQ9dU89C0DjayaoeeT81B1AynVSepNnghpAxhwm99wWkNDq
YWtZ6QgW5cGlMz3tjDR0i5iT7ObRKXtTW2JTFCkMhwgngJju9sqzt2BB6Rny
ZZhlOc6ZaG8zeBq65ALwNa7m9wW5K0pluo2g7/69NKUDUnSYoAkhz3dsRP9Y
l17+FIDHuQKJS6yuQXNSVDNYnT/OP/IMmOVikQpM08I7EqVsYoHAe9nJFaKJ
cMnKmN4wNBFkI+X+Mh5gnrx/tK/n2GPaXiEdftGD3SeFfo1BaAIn3XREANSq
NplNk32Q2dnhfvDTE4E8u/tSWcLBRAdpBjSzg/USr7z+RvPgDepC8FOIrb7C
IKH6Gy8t8bk387bHcs90j3GaH3msEirWc950oK+wyJZeCyUSJ7IJVSF3p51X
8F9f6HQT9WRL3End4jSHm4BHpePo2E8KCWOUCW83FEpRAF1okmuVLVTcGmp7
/V2v4u9Ghx9DM35fXEciDtsIl4QEsz0ZKHXaRHUaZyYtGiLkpwbMAjy4Mc0s
X3+9HQZ+KvPOY/lb/LEEVRSTpzhMAu8aBZtoh9JZQr3T20JIAKGAOwUXOCeo
4Ns01UQHKSSZNG3Ts3Lw7wqgAcozSPeslRQ/L1MYiXDRRLH6Ag25Dd1t036c
ziLx22kTWdjYXfKPgP0PW3yl3Lm1KUkAlKMOAAjbSj8SGZ5/6SEs4pOTX3ZS
Q1VqXICoZ1B3a0j60103sfihwjoehyChvYXsafIm6RndU8BcQ/GmbQKHujDa
LibymcJRnej+jial8eAIt5zPqTCVsvZO7x7gRjdp3Yry/qbSBX6rEkwAJDSY
lP6QbCNHbvUTIEjZQ9fSEI3C0vgKE4CV3+yrOqoc5AZiG/r0tb/YtKRrHFhh
4kCGBu7OhPlTZdMdUlOLtip+zY6Pd6wQc6BcCR/NGI7VWBdDwkuPc2kULIxk
J+Jp5mObi+dWMNEiKuSn+jMe7o5ePkErJVyEVTUHfawaJVnBy+cpPG3nQn2x
SotD5WVUmAd7TZ20UvRx1Cls/Z8pEsVnYuH3UBSAZDXkF4PGnwXrVtXfDFH2
hRBDhciMvIi5QBTIyQbLs4lEXsv7ilPMCS14kc5YgiD/bNhX/JwJLHafG3rW
dJ0+aPRqj6TVQeobFQe3CLIqGbCTOHIJZZwcIq1PlZkSh9ddZkdqoyq+ErHw
5uj9m6F0PzCxFeu01ijch45IxDWm+FU98LvbQ2C0mYaicHTjCmRLIBUGauzn
apZUEm2TAOsb83KbNdZ3lcmkFLJlsT641QV/sV0YRxBiSVKWux48VXcsav1G
e9WP4wANZ6N6E8VuI/nT+NAZjrYYL+fcPAvs+pScsvVRROb9blsAyKNtDtpE
eWwVrXUBkWd0Pkj8g/5tJoL/CbU8UhS+xIuSTxwXovJwpMY2t7oOBTmE8nxP
hjWzRl6K/bzDElgamNxeLp4UZCbvNMFe428vp0Nd05mK64Lvgj26svmPh95v
7/aWyx8ovxT8gjFnNyAtnaF3Bzo+vRTMrbbF1uHU0gJpQxSU8B1LL3R5OfeG
2R7OF8XaU/dm9DL/pocPrDwi3puJjDs/KUt1U7NV7EjzmMwjdNQFG8KYynp0
EDtI6/quZeg5tYfdiEHC+M196YRa975mDTSVR+92pxC7qdBR64cYg6WAe3Fh
nVKuyWoUJa3hzw5bl9Vh+y52n+FsdLzYD5rWSPvPjdSbJidJGJwTtMRoac01
1W0tiVcaiNpBmxffXuVcBSUn5tuk8TR1gVV/SzF7k7OWK2dJ+OQod1J1yQxY
opIxuoJEo1AwOoLtWiDh0cXSHNXAvHaTcdiO3r2wPNGM9C4LtqV8oCCBmOk2
kZMssdjLPBtzWJYLrkasWh5ZD85momiyllYQqLa8QpWWlnz9gVCuwF/7Pc2d
DELg5A6CmQBu4i3JDkCntBXdaRxWuZQSv7t4T+IfbfJjet1cu5XbVwbJLC7p
oVGgTEY6ITho+v4YZjN1+dAciLdPy50s8ksERIlEjNaZDhl89mCpt0YoEwmQ
1vo+Q12DUMEm4d0fG6nHCzt02d7gVPcAyjrbFNKeFQO+2fi92sIrp1Ln5ePc
bnOzKTI/0MOs0GF2CGwyIaDItGCj0SBxToOY0ot0WMuSkp96ZmZEcJPhohSz
CcT2t6X4G30e4GlRY4yPTcSWWreXoDIDXoHc6hBEalQfSUckM8GDc16FPrRD
lI/6IT4AqeXqRC5aFVRI4NCLEqmQ6/wJyg8HuFxruU0plUyVwKxVWE/+B3VE
U7jYhImaDz+yQ0tva4fZgh9ZRAAUnVjpk5CXSE+70IwKST6r8sI+kDuTZ24W
5gRV8lnRDkqLgKuSpurHFOKJlQ4te7aphZNdnK783qVsRyHpbpU2Bh1cBWYF
wPzcpcQnZSj7074ojlvYDcbx/fKwt+07AStkazDAXxDXyyCAnOI3BOZcr+Ra
CdxmEygFJEhKbgAAqW50jHCqF2YtXGr7IEoFaxV/nBBpYU9Hht8ZNqdmGxBL
M8CCCdSWsy4XvSU8Wcmwzgxl+aow8xLtx35HK9MWzXdCFIKYE711O9xQoaeI
qarAZXcuT3llgXaylf3h/TPnWGuqqd3wxM111aHCNFv/KQTsT7VYsGYgDqTC
gm4iSonamZe1vcZVabDZzCB6Snb8Qh0343euvbf56QCio4109AdHO3VRGX05
FW31p3rTq3izh0qge8/nUDN0NPFFW0c8zk5UJqZCvZ2aC7OipnGgGQF9Kfh0
PK4zOJhms8T17P1dRT5JwZ6isMOx4VYbJSPmbuEOY+j0BDDZJOnUejNF69JT
3+4VNlQ95iCRihgb1VMQ6rBTG1dlPWjOlhyXz6z3Gi8pBPZ70GptFbD3IrGd
wsBelSHTk1NQlPNi3hSYDqpTEKxFSEAqAmY/lYvzhUjRnn5DiaYuaN0hB0Lh
vKBRpIpD3c8/KOcv4CqpmcaEuV2rj3Z5XRmDMNeuLqCjb9I1wIoxo6S3ovCB
6gvHQHeSr6Kh4PlCt5hJlTIBsB7EdTZpNOMbDc2Ozaf/+K/U3curmo/G2jjx
P1n6NLlCipIoYqs6uFuDqrNf5qdEvuaTqpSP91djh7iZxP/+Y6qHBfvY58WR
7z9ry5jGbt5hHSz8pumjWr7Vdh9yBF+xAPS5FL/td/P5Ho/OmYNHDc1PMNlR
f9IlDDAOXEP+n++Tj0IDuAApdxvU2hgchopc6XofUKWi85ctVnQe4LbN5p4M
WiH1mYCxURrAtg6BwJ5JrIbFDFkUecPWFhC05H/9FOZYETT8AXNZrWeCWIe+
bLTAGj1vMIerL8ggKwX5Pcmc+EOfjLnjxkQl4TLR0uNy6wtDVHz9ultOt0V3
yGt+RgrCq2bBhtby5P2DwegcVTudgem3ZQXNw2galuWOwvE/6Sx94zUeComH
DOeSvyA6bm2S9jWDN9kP0LErWdzWrhKVFfFjWHyaWouK+VTEt3zGGTkaca2h
A6176PwBZsDWlJjiwxgIQRF1m/+qgnN4TlzPdP3geiuFIVohRZnw25O7oSEi
WoYaMyjoHij+73Oqz8YXLjkVPUT5WUfmEbdlmVlFdA/kgo9L3KmdMRcAd9/Y
dUl1huIc+Ic0P/rnIsBM130jqB70Bt65XwgnJdvld8FgIll6vkOVTXkFINDF
ZRU3N3QnmWqRbb8dIT6cdjexeTNY4j4AySnM0tth42JnX8Da+CUCSjxYPZNY
xzxBOoZ7i2PYP9On3MnOihUe2SjAn7nDX9zWGLz7pvGiAV9uTBAIReqU2BN+
4QEool+BgB/TeWiYsYHNaWqZHXnke2/shpmcMoD1PSY9mdLWwC2Rqa8iKv1k
nxvJBvWtArFPLLZwRRSG6ZlDyyIVUqpOniO5HYRZlwCMNLRBV0fccVYD05Wu
XDxve1I3vQ3fH7W+2e+lyOQpbZS3tHNx7YAGWC2/xsuJGNxksCgPlRpAwvVj
5ZsB/C2GXnCAxgkYsUSoSK/wrkFbKpOa3XxdKOs+mmExbswJfdaNC0KL3fKC
EH9gmSj1lir469jNxH8l4CEeQut/4M1gR6qOwTEDFFC6J+KsUk5QHmSZtvVS
ZU3qaGr6l+DnzqKzT8bQ263s4FoZLwa+MjejeZOHNVfqKRtsqaTLXrRbKNv0
sN3+tlJxWtf2/83smyaHfhI+rr+mxbXFLHpwnVUPpoznZnsshJM4Y9tQwMkb
eZISk9X16oDZHOn8z7ZndyT+kKdbutXO/nE8V/p53aTKsaaxnSk8AwEPMzL1
IMZ+VBoUc5eN+jQS59qRuqLRXyRAmAxr+QlxHmmd2jzOSP5ISuNaAQehJsRe
Oc5qP5G/jNlF1m6t9S1/eFP9+rIoi2tapLG/Pfa0hEac0ZKp0Ao90knlP4mO
5MzBfpEtHnBIRfbEt/zrkhRjKH8RuHuthV9FrpPjK0JI1jG+pz8yrmM5ijSK
Ekn4rPEZ+K9q7KbBsyrs3YXsrcb/tjj1xPWj06RD68uPTyUGu+c76U9E3lUS
dZBfMKDRV6RVgC+uHwx0giFPBrByJ8RzUoCUlUULIYW2ZoYwiA9+/eVNoDlL
k1T7p+uprjiVMkamKmxx3vU3QPjfTKApDPmGZoQFnNZ/czBCjsjKpxkJmmt5
a3CL4VUfFh8/o84lvbU0oWAk2TAfvKg8Sn54+MYIMtCT5LdPc5haHN1vVNib
95gQBoAN3lRbo1RIa2MyBPHOOWYEj81tZwUo0519l44IjZjlXwQuZE5TymkH
SeRj0xViKfm3RAvfpSKYPFp8AQ1qHoaGsBp8rsz8qPdd+U6sTDEXSVWq6hR4
bQMmN6b7NoCadSHWpze3OwH/c9O+U6Zwt7I8wVPMZTXEBQxSklHPBXmUl1pH
0ShEnH89NAl6zvV/eaB1T8lFjvoDDo8LlSc7u/hMHSemPt12I3SEd1ruxPOA
j8SGx5o2pULlX7jwPZhaMEE1sjOgvRepqXMAl4Sdn3Mk3mNMsQSEi9iZNc4S
20y7xz+vpFhGRD0/bwm6rHlGk5r9Le4MqoQkks7zRherT1wrkhpBCUn1pGxU
pF6TawLMpLv9QrZ47SD9M27uXyD3B0cDm6cVlp2isDeybA8TcKa18BTmAPnG
fGOymQYFNybHE4jKEdvmJSX2WtCLtjM/9q5uwDBTjEjCK0rn1GumZbgmnyk9
maEi/fb2DjVFVjoaYzhKxyBS1EYdk30TZ4FQ+3PsyWHTXO9aAffsIRfBgL77
xraAVJPOBxXlqn9MLhT7a2zwkokK8Hp7kPC0cmHrJRjvq7V6HhJ7P7yH4HC2
gXfavXYLp85S33fS+SHvmkoVbQZNtRBuMYLvEJAsMAWrfuRotUt4G4rWC5Td
0eQ+j53ZUonIbP8HWf+Qxf6+t7ni2CdTY21Dsq6b6STeY0fTdwN44jrJjuLk
9K7Y6CqhfIvLfkO7258l2eaU+GhFSsPcuunDlTj0qPixYvwd8Hz0ySODnb0P
qlDS1ygpHT4ykjuq9RA6uQ45cZP/SjbP5HObick8XJnturHzNSm5kvjWKUs/
63nilbKliw+tcnHphAYv2X6+v2908i0ggoxYgao3DPSyJkD/l4rUD1+pR95/
bQs1DF6Qcg+ZRQwlGsABIDgKrbw43nmEYqGhXsG/GfipMGd5xQl8cvq1us4K
U17BQ5CAUC9dYkJOTtvgJQ+p22hvLJF5Hl9MPvWF8vj1+5nDDLdrq1TYRECm
rajpW77fLqgM7ORrz+MbrPPzSU80Gr19vvI7gZ30fHgdYd2s6EYP2sBMvN40
cw5JWapqAV70Nhb3d2rWbrjpMoON8pCmwrBku6qgptF1W/FKKhbZVFFaLwd4
7eeFeNIwvUX+p9Rlu89+vv8hEketU7BwKcqlim0lFNAveiuvrxZQmkAsj0eX
4Pfc3yi0m8nnmR40YpIvKHSus4XU6o2pcp2zHakfIfvYR2FEdav6hwevJILU
FGDC11dralA/BmrpAbDuLfPurhJWayuhRtpJfvyGt59n11v2LKct4IEyke26
C34i5UqPwjGqJRnMjRGURgTcyb93Fv8bC6MmuqKpE+s/rCgeUu4D/TcZihJA
ApRFwjV/SLWqbYQyHiNi+V2Yj6N0JOGYpjQ37zkhCrmoM0LlAsEjVlRwzE8B
w+zDFU484KuquQiuAuqLVgahqqW/DVjZn0UHmYs7/81ESPs7VO/5wOhbiL9/
RpTGD+0p+QFPYurii/AEu1YC2SYSRJbeFIu4/+Z0Wq4xnVBu/VogFkUm0/lL
8Klbt5vAxrshFIvhgabsnDuhDiieHpCaZOJZ3YmntGhAVPlTUpuSAdEaCnP0
ocdv4Ch2GxyLpNWmWeCkYXat9M2cHTfxwvS7n5YvZ7XL7nvUXra7DTl9/seD
piXgIAS5Caa0N7B2nOfEze4VhL/4q4XrcuONJio85rcGfNXOTlHjMwv7iGAM
bVY2Yk5uhdeeGPl/YWeuhrXB3ymfPdHKaxqqmqFLylKdydSktXwpMTYWIUza
KuUYJVduSVHdRJntFRKfFQYSlJm2p0bOyAZZI/sx+Wbc6Dp5ecpBJRD3m3/a
Mr07e0kzD8L9Hp4+AH/rOPYEc7V2FzlcUNkgFQ8qj0B/KHGtuuDOZOcVaRxu
8CenTe3hqpNdYGkQLBjOrt/1H+5rbFbSKod0jmin6AbTJY1OWytDsNyLJcfs
sKnm5CA/TlFYCrYPLdoXvD15bdep9wsnWoLYlPKhx6kjreOFRKvk8OjaTQve
5wL9Egm69RbrZr1b2jZMWttC7cGLbSE9QhNWB2D8YArHJfxCpjO0ueQbAyo2
Ydt58RPfp8rbcgID5elCF0hinnbrVE1TP/D3izA8heKnjF7VxbNFaQBJUtNH
5gOzRDO1TMrBAWV6dgGVKCKO4nM11+7k8joZk2jqdta3sQINXGXgAwQRxLFI
wNZUpyIydHAkBaDwsSAKdosRcruD+67l5LxeX7NHi+Z2GJFgZZ0cZA7f92nx
AbJS120mSKe9tFjkLaz6JSuYfJa3zYLVdNlQI4LTu/A1Ih5aVx9UYiQ0n9v/
X2AtSnVeW7rTXx2LGvqB4ctIa5rtWIM62JUk7BHBtiBhBWQAF7r/AgnOGkMH
fdeCz57rN08eec2SoTp0ArcLJBQg/NM6qe2SBo8jpnkEEK7IzcBX/dsXNg7U
kdcQArMfkiop3ZpoK9Q2cQ2j7KYylLmeuD0IBGqJW76TFEvERqEyLoafqfKp
vaWHMIyVK57TvFlnpNVLF5p7s5G6f/hJlOPhWyfwufuWMEMjUU2op+AvoICf
+EH4Ea4fmHjUxHAq0ySuU6lbZYAcnJsfsGtGsnu9Lg9QAuJG0467eHI6/89/
J938P4FHjfXBgXqmhwcUQYsAXX+oYq7+uDJkHwZXCr4s3U9pzX5C0EkKKZyl
qM00H6CeAacxj3u/1K/nRP2CsUcp5HqdEGJdK9mx4vP1/4mRL1fb6aA0NDk8
YOAreoYdRXaVLoAJusmS4hIFflWLjoMuF79fDdr9Xx+felRj9X2j60WiYHdC
1r0MBgyOu/e7R2jj2ChrvJW8yoWNhQZOTMUxSmvouplHCkjk+klAanNW/Yve
YHhyAdCgn+NYivNwbpaS+MDmmS+wWQ3Gi3nA471dHBuqD79tcoYB4O7fA9jL
/6/KnbvARMdmonlZ/z+OHYBqs3ep/SdOOMOzuNgAjTF8BZVo5VJrSrBGNyVD
MYeiWhUt/9uUuewt0X+HIQSY4fCVwiWq9m9lsnDhCMNTNjCe8gJmyBdUzF6X
2767m5ND/nY1zhlqsvF/d1ZRqkquYZvM2jQEoGanLG+NRvurp3LAzlBLVYcJ
ptA3y9yUfHyGPKmGtmH9UwH9TF06A7aS4eZ/fYZGRC2T5Wj5rwOrGKlbkV1s
LkP6w4YfVk6yFLReRNDyCcrIarej+CBsFF/YW1+JT92tcbKr4EtSzl3jPPn0
UoJHS7t1smR+yNe7ZzMs87R6Bhz5RXFVheL+zVogPbImQ0UUxfxMMVU31RgG
tPr6/fCA/AM+Rq99I+l1+BhFvuaYXmjc1RA0+/fNK3HyWG4vlOiQhoele6Fh
iVoe1yppfne86opYQsVzMJ796VW5AHw2zDsUD/9v4alyRkH4BysAAspXMe5N
vS3sr5SYcTbJUtjEtTScD1erNq1Ui7smrI2uZa4g/m3sSWgFbcnNhh8PMh8g
EPXyOm2lcISd6jq+jpq7n+IKK9eFAC+DBFhhn+RgJYKIs3AHjeA/B8Mw8RNS
v53KdYvlt3Lp7kgl+SPQuTqfzSi6Z/KeCWtkHRPwpbXvIwW63V92ZleyMRGf
cEjThPoEKTqyPaBQlFMmUO23ngf3Iu2/sBDXnN3ifZ1J7MYvni359p1kzxcQ
SJHV/PV9MH9Mvii9fIjw13w8DfolCcwAbOo/3G03yuS84VLQs+S6UoQl88Pu
rY7nrlTvXBlw/MEv2trCSir1yfZOEMF1/mbcRPg39vyclDhkCB8AhebTaJXH
kQmBkxYzM6DHJX6v1rqLQrGMk59efPULxoKphgYa55KQA1ltQQIZwXE6D+IS
SL0v57b0KAc/x6ZJ+sjsHaOzvn8DkrW6q1ifEcmRREWIcfg0UzOkI8zW7YBk
Ex4OPrMSMvinj9J7U+QP43pBfWaG+9T++gSe7gw7XhHVN0U5KptiWp+Xu2OH
bZhqnI2uRidJtq3ERuM8ItnGgTu+mI2OdUc7xAz9q4xxGxYAsWutnsJqd8RS
TaQ+JuIq4l6G2l8bs5WesI9yoXmYnsICivUpjogX+W9jtJRRO9H/3wDu87qn
DHEiwb22FE80y6J9qDOL/9zBkXJJsWy7Xk8zlalvpZzawc1+YpRf5+NOIPVV
pCIlVpw/RgesZEGF7pnxbpThyvfwpSiV/KXyw+u0YYrBZ3fWtu3Sg4h3SMeg
G91WiCmEq24A8O4lroHGAr808UJmzBZotYjngKIbdXrYTE0UCpiMvlH7e+8I
HZ9lrfJXtdEh2VcMtCmtXzkRCDStbVl7bD6HhbKrTDrz/7vs4TwOyB4dl3R5
BpwaTMubE4UBEYIyGU2cPyd0uPgiBZKvWYt+snVzS4Kl+GJeeYQozwyp+DSt
o1ELRaI+pafMDh26QOIyenz5X2M/nMjVkgSBWgvpFsEIhv6B67KUHdCwwW0X
Ov4I/aZdu6VtCkTDcal18hU3ndUzSWwGKFQ31QgI74Dy+VUYYLo4D0zMtNAi
TYFFBJaelrnMm7CV8TQahbSt8Pg96AuJwUEUOHveO0dcq+74ikDHoB8yier7
ViQGwxNzTFUjceE5SbSREcGoVILTYu8wOvK8jv15tONi7/80MTdFh8pasO1v
3XFnfD6KptutjYKBTto+4LLU5NFddHSekbVPi0kiUUOVlhFLD8jbkHgopBR1
qmy9Nlh11Z3WvIq/pAPZIoos905X3trFTOD1Gvsxu9Oo6f53EkirQgEBBc/H
UepYYsF/GoV7Q3zhkGhHoxmfgnZwN3J91QjmpgRshE5nrp1LT2PqH+fXVtVo
rjGr87J6hAkegRtbJzaE0ZpyZUQcOF9KXe64taQOSTGdAPplQM5NrE2ijMQG
91tE9ROMnp2O5UK9aRPdjRanREfB/BDkpODenHiV8yrcOIgdwkcHcJQm1nJ2
DkG5blhmNOx+j4ogyYWNLZh91vsuPf9w88YMKiWCxJVgcEKYFG45UsGuQV2x
FnNrD9NlvKAl93nelX+578YgMejt4q87a/Abj+ylmw9K/4cj8GP27dhFQtYk
4yDKrb8XFiL4gaUIzSjfLRvC1B1Tuc3oqO/PhKw6+A6hxQTE1xBPtaECaJaD
u3p9RAmPCGaRvRh7oU+rO3SvVEtdZA5XihAJqb8YQMy6xDkh06rQfCmT34D2
RZEI1zMNgGDceqJeCqrrI46N3O4cxAXhoXxEuaZiqH8qZgf9kgQNKPQ3qJIu
LhUTCPGvPOIH76vJ4NKtjuQbUhRko2CLU8+EtnSqxihqH5ydlCbIDD6gP4dH
SZLPKhEMxCyP0ecthsMLfjiIVW1zERMWHAHENq51yYNFS4iSTKUkuNciwZk3
AxaYcsP9WBSwzXCyoxFiZzeUo+5tO54GP3gJN4/z4TaUn+9pquwia8C2ytMZ
Y/bmg56caDM7+redtHrNZQrDBh6Wf3H9cqTYGfEhG3MY0Tl4n2BjSKBWRQYX
GLGL0+hWJI0+GvAokt75yQMOcuWIqZwaZop0GSLyRserp4C383SSrn+6ksY6
jci3lREutm7KkY90Y8H/qF8AEBnSdIyfc2h3vCsX3FBn+JioZK2OCGPJRTWT
Jv6Y+RnLqmEwQZu7SV0b249+DZGT4KjQyXQA5W4IXIAJcX1wDOVSl6bXKlsr
HCV/uNWQivPAW8nY6ny1uOL4tjrrtKVWrtTEAHuEAMOHC7WVYWu5qFJ0UAnx
fSNdmIiYqN87QuppLW0/rmqMNA/o4XDfQAb+6/V+dA7cbwJqwOInQ5KB4eO/
KjM7FRz2X0WKdVU/QzBtWVVe32dlv3p6cwIFz1/Fn2KMSQfC7wM13gzY/hLF
RrVuTlf+YJYT9jc/zmHTm5jPr0Zi2XboMetNr+9fU21nkz0zeagNurrfc48u
b39BD1yteibDxFx7T5sshJmzfbmyHSjakSlblRoVlOPl+TbPqyXhhVFLmI6e
1e6hMLnqCxkN98vJln1qB9c/7EdULAjZYbbCGRnyxz3/y3PuqLSoxBMZLgvu
eAykkyvJP57tTakCOFUdr6HsWtNG2lwxoDpl92zBclKNmj8lrslHIELYNDS4
kJqZ3bf6UcKeV50hHXDHBcuDmC53ol5G+vxT8Ms5glnM+HR0qLcV/eo9Bepe
yjIDuqV/ZRHwJGmCoV5xNqqPLKP7ROj5kgM4EDi+vhCgsSX1BVxUVkWhnQWw
f3i5OItU0TwGcflz9H9PrTfE/OlFwMYcmawgrf+FBCUQTTAP/apXJ8WcYChk
de06YPdtYW2knbJHokQBKxwXFzS6vJclTuw3kqSQTicsEVj6DelrQtZ9Lizs
RhMLsNZyuY3uGisqgGJlC6tjOvkkuKWrfbgTP8xOTC+lhrpTtCTLICyjLJga
h+WvF0BRL0CMPDCWiuXXvUWeid2m8nXg4ZHHHwePw6lOuHK2wc8X4z5weAKT
G7A67pu7jtDsa41h5xNYDEwVxljpnHzL1hUHvmryUCHAK20hw97aohTplBCG
VQSrzKwQxKf/IpZzOct+EaFHD8U8+Nx2oYG4DCWIOGnJfzcA9YgT2nCjMKKZ
ehBbAwdggvsoYYmO/dwWgyz6Q5dogw/9KnIxQFQIjlcjImB/rwgQYzjv/CBB
7/7/H3hGZTEq850mnurk58dEc23/HnC7klzAHbNHujSsk1mPhMaWG7oaU8Le
wLrWksGPvV4KSASHegpqgmF3lz3zfwFwFaIOnKI+SoPJ0k2NEUHMbOZSYF3x
kvIPGf8pbcBUDyZ/TMMcjSfuZttPUpIdmfFKgieFBWH8bZsDQw+B65i1Egnn
ZvwB7UaW65JSqQgHpwT3aoNQjcZQ7YalQ7nJPvzyPDpBD64inpTka85PwFoi
a+MOCJXs2USXKWWrBbPBHBMf9hUKdfQ047IJz0H0EHdssDUJUbxr1PdT0LIT
a7l44aIPiW8q3wurHTqd7xzT6pYAs9uhj6lRWyQ3mim+NfYeZe/e+guclgRy
YQtpIMuRVzykuke8YFoY05NR+Y0+4394dw2B+NsIB9wIvxwiX8bKtPMocOsD
wR0f8DClxvlwdoTshwwLSPEMQ7BcNVeS/SUKI1gVUiSVsIhet73ootSTnsV8
5lgSkmjpbn1KeIp0dh7u+WXjgEGipVZJCzX3/LkSK284czd1hYXybBh3b/1V
4Q12PapwzlO17NhVoibpQQ94MKA5ATvkKwe1pudEVYZJ0uzZJclS8KTy1FID
yBXA+/PhzmeKCA+ZhM0MPWFr6LL0cD7tzwB1zKxvLZnZJbNysd7CBsMsmpB1
UCJ1suX8rpA6niq5OuoFKDdwzE3c1IQ6QhDbkfqJ8exL5+v9IIxm36rBlY/t
EeSv1md5JOggKSYaufNApaWgc63tFV8bF5WAIbeAp96fkV0zjdEHZQ+fAOyZ
yEO6Q0NUnio9dh1P/J93+zls0ZVbLq4MHxtTYTVurzoEOjKcD7+POm1Y2W/N
0RxdLvVtYDL2lZaZKjBP9eHBzEqnpAGD4C6ZL6Z/7T3+DzOs3Y553rMmApVW
SJeg7V1LOe0sPg/Kzl4CIRsGlyAv9Pt1op9AQWLkLtSie8/CZhau+t93d8jv
6G24Ix1nl7TWGqBL+HIRJybMZBHMnWf2fucYen9Qr0BdgMmfDdMWTjO+Qm/y
RWAlo/G1FczDTmFIObCNujsU3WEr0muqz9XPaT9AJ8yvJXofR0zhJCaZsvHY
nYZC6L4d8hIkoKBj9MUhpnEcKE16ckk2oCXRjlq6nIAhlBK0AuuZq+/ch59Y
6W6d62+MTbALWu6G+a4a+3NEGOp0jqofiDjpcBMFSuhQA6W6Yv/nuY7eGZUq
CKAazZhtvcrw19L9Qp7UID5uCiYqJCM0TuKyns9ZRkNoF/nr0Dn8eIcrMdJw
IjaNMWY6+ihuj2Cq2zuvi4XD0BNIjMCXFoL1ycOR8mdqKGwvwKG9j9GKJj0o
RhJwmaqDydct6QQ5V3DMrvEGTGZXLs64HjqSfXCv4pBj1NfYz9XT2pMVOSIq
bUzAqr3m+Q+Bxv0wab+LkuodoRlIr01Olop2G1eWyfzgqON18LSCIfZk5FpA
9R4Ko9Z0hUrP2Eig63Zf/cn2vXqsx54IwVrJS2PZptCvIePcoTaMPlH+G48z
Do+T/ljsO8IQM/juxJyZbYvoAC7uEM3pe+jdwz0wcflFnh8GtVZsrQ8OBxHc
pfvkjen354Ycvm559mTpbWwSN1NMzxL9BOa3WNNdp+NU4hgkCDUZi+HyRwOL
qifzdQqg/xwZK12VI5rUKg3hRefRc532ZfgyErHA4oiTo6sum6da0LkDk+nA
pLYwtDosFXl6SZR6TEUJg6YaxgRIKjQ0VLcHVN2m6Nd+TiELF0y0NyS+TsR1
QCAUjzBZVEYY+W9rnPqgtp+NC1G3xyM1n0+UB/AKayl/2VGbFPVaioMgjH9L
vc/1H9xmuIjlI4L5qjVGOfiIxRyqy6ZvEyC2+uKZ7JuqyvJm5ootR6ZKHPy9
YD7nZRMZtcpIvDP9DfUIqT0s5wCVJyhbhYBXyMiF4R+/6Bnp0C8VKWB+iHJD
3mTf1KgKx7awO3TffP2Ovprvp9gnpotsaGAztratwQbhtvYKORny+Wp/0mVS
IT3Jys0MZTeX6gU2NQ4x8HLIcvx/bYxvdpuByO/GSEpHmGOoQ8bvFckPf2bo
kHvyyL0VvMmSDJbezIAGwGvzl+0m+Pu+lRQDBLRn/wuDI/zMdmoGXRaIZmzV
01ga1gA165XNPf/7VnBHTG74xhgaX/zkGkxDLCmGXZongMSRttMzS89q9cUt
nrmajh8WiP1L+Nk65X9VqCD1063t3OYGpS6zHTPbhTu53Y033orWzZKxjiDF
bBd//a+eN5GpgKcRdgNucF7ufRcxrQN1zlXWh9U8qqaGICmAdpHCGL7fOshd
iFjh4ZSbgCZYw0R59R0eRTA6/hcsw+3m/ozV66Z+9V6xDFsFT7Mx87i+WBLe
8uv9V9S5XdU1ng4gXQ8LBhgjxxnGT/7LNk6WXNPT6q9N+W9/pnBFP9CMqgwO
o0cd8JssmXO5YbRlbOM5eXiOnJ3g/TCG2YK6z1HHxz/5jnSzR8i5qV7xyGAg
nyyGyXuE3W99Z8V1FYdOgDQ+tdMUpoPvXESLRsI/N89eoSjWhYvEnDdBRqAH
K9XTXwYkBdNlxiChorWcvaviVtLo0Nu1p+gKMJKPI3P5wmTNyoMmQyDYzkzN
ujlNlpQ0YNoMpKcK5jpwG89GVRZTdpsPSjDsBdLOUbvaTFPONSgwSDBZBVeH
37ei84iqcjlVVLQpjD0gx8Lkv6LM/91SwG9tdyOs/M9ZjZJBMLAV8vxuhfQU
IWuldSRKxPYYsvmMnFI7ZocabmCoxnVzBF0z6zlKPyv/1Q/Lqj7nbMWRTMUW
9yV9Jkq2fe0WU9Dum1QDU0UWlFOyp4PgOB0l2L0F5Cuhg1HALepaf7Chq06W
uJG5owLBo06RDJh9Au5UAW6MUFqHeD/eEhQD9jNqerV7FxBnWfuCxU80w+NW
1tTlrATm/LGx84KG4SoNeH0SPoa1kbSKie3QGlipMmdqpzrdTPgQ1P2rQcAD
iEKG34vFsUJemlPfmz7PoBcHhtcSuJbCMNjNf71rNzeLt/jopJenL+aOGh6u
BqMwlEzx9XHbOGFosEJ57yzTmK7O/CDpcEPjjwgpswq4CI2CC3xrDtvjbns4
TyxA1xFxGBhUv8Afsg/jh0LHa8tlSysxF3P8xYcP+XOJJe3U+jKvsK9t+WQi
sBgHmCGCDwy1RzU3DB5FMSuFIceLDR9tLcDhM5VOrGTM8iXu9IGacS3QLwaQ
LIIuZXy+wk6xlEZMacSbIk7nRbeqmujNTMi29S96i73V3zkxQ2NlqWpBTbkN
OHdOTnpxZqQw6lAgGxk2Uliae3iCo83P9MuEpjETIKWH1mB/Az+AV1EMy4UD
8EWOcwpnAEjQp5GdGNM4AO97LXYaKBX7XSCA/6eUV+aqMlKSjOGMWOy/P1u1
EbdUQ323YHRqVp9m1wU8A+zMqdXDHXdT/n6ByIqeUp3oAe6J5Q+mNAsKuS5j
FmPiMl56620S8gIEKI+LAFRVFBlk6A9JtFdkgYxU2krCSWAxEOKSnOQ7Z5Jc
+hOFKuYLDkgzoDjOva5dFL6wnmeQlbHu8fT3zOLzK6NmAyGUMR1NaGgz1Kfd
ASl9nIrW0wILy7YosMvbL8zUoJ2sSqkYZd31wGftGXM3RUtPe0pJLjwC2cxS
LfRm8vbTRSk0dfKsYMORARqegA16f/fX6MZW1NXsYEWh2wOizh0Wip326HFM
JBkOeNfLHUzbfnmhvImyVTdt46Kl+BBOXow7flTD7ha0ykpBsXgbIn0TMPQ3
y/IVo05fFQsAJu+KFXuZAH7uRY2aoIKsoWav/t3iInOAX0mCL8rcx4ggn+Wr
khCfRDsIXbbbNHHS+k85EbPpkWIFVntQ2Ow6evlF+RCiSNEqdiIrClcBdEPz
oUV0qc2SlH/1xaQNR40TPUBF+w9cnqH0GJgQ/5g2yLjGD3pxLgPYRSFGUmmj
FrhsDlcBaOM2fF9x4T1XCDAsKQHLLoDJ7xzQJChLtCYFwD5ExKr6y5sSVGSe
elmlNcvTXlj8HgRz4UDlUoOZazEFgWtVE7OH+Aa8sJNYfIf2LaaibHfnnwMo
EdFqeWzsLm8fM/MfoZszlrKEz5LIdKc2TQqDmIk2fqkIZnWyfeKwPUxhqrlr
UC4EP0yn7yyeMjKT0u0UstqjmOARylLPXF8XxQGWwnvck7JLHo0l/q4kRumz
W4qSA4921bEqDG+VL6Z5cQnZnGUlFP1zES6phr0yrRV35pDyO4Zhd6jm0BBT
W1BYxoA3z34bVs179wxHstaZzeViOKMt1oFUW00vy/m+6x7qLP2cQb7+4Kqz
sGxakA8Ym1icbS9ZngJ7wrPqHvfTlPRwlErZ7h5/q9S445UDS94BXDVKI4K3
i2gHmtPsyuxqAM5yJOsqp068XizvQSnu13otW1Iwtd2ET1ijbEE37q4e994l
hcIQzslpmPK8Q32ohzLqe9aYq+dPjYS7BHYeSqDQ5n/DrHlN8c/6BDDGYQaa
VMAujlDEzYngzOUJzSXjhnI4uBvz1m3Szuv7fv0F5DR8DQmA7jTNfJ1/ooXS
+eqIoT2QseyPwPBevTdHNkTWb9nLFkLIuZjzfTHblKinGeuBJXBSiO80btM+
romj0J6HV1zyGrExSmAqX2CH3QmZNEeKPaZ1aNf2VSRrhwtWusjE6oNsAJU0
mIp2oPcENCZM9F+I0INXimh/9SyWr9r1NeNxhjSlrdg7bWKKOZWZNSLV6rUt
fvE/41ITzp1CXmpCcZvsQZac2JETggSpiFgARkADcjBCc/e9/C2UQ2KiPSDw
Lmhhg5unHbO3UpNlsYfEBpPAdSWgLzgUXp/dfUS5JpyywTS3saHX4SqyeZlw
IImcJlpm7Nw67jFqmXqsNq8IrEJmJiRUv5A9JYlfORoD1hteRntlE40HsVg4
txt9FInWbW3lyCBpX5/a9pKQAA7QjC0wQM2rb7gxD7E/YMjFFx78fpvZBisn
7Y68NTZnfbpsvCywyQGG/YvLI3GnzNfbi5qBhtL0qtywUzTcmLGQwFQ15mPw
OGHOOCgdf1LAbXX27hVGpL5gtjh6hStAoZC1oa1RFyDdFDJogYz0vNg++7q7
Mi26GgVocLAbgYfcM5b2+BoJPNEwQ5MlvCRRM+GIVrDGzBqRZNfFWbh6Bpkc
AEnTSvQKr2UoZg9Vo5prQl17db0EXSID8b7z0pkGNqDJirbx36Ug3G6Y1pJo
GGt+Xll4cunbyBmyq0rK4P7pCx1Bmm99PfrhkG6O1ndifwTLSrBoWm35Ac6O
cogLVrgF+s4eD/EKBekLUYD49rZQ6hkSM7UIzrO4bXd6XNgwH31yeypUGe4b
KO40VhitwHmLwYHeUdo17FcK9R1asMxHVoChwR4pUTdxfuug6jtCMuFJiUk7
GGZQE1VK0E4m1yWBW0l1WeIFsOBnnntgW/OQy2sedsVrBKUxam4HHrJW3fRn
/rNVIxMkIRLQqeYx0Ft942dK/q+218H93mEUxrb0d/aMVqkYP42MCMOC2sKq
8ic/sLvHuCx3k/1XmlQz9kbcU1o75PFZTk/4ItltI0mRBJ/3sUKKfObVTj2p
zYJZ6qhP3ZqsZCql3HOKd5S670dtUwIzADMjMgGKyV0HsvPdVP4vcojPDsTD
y2QW0pTE0nKlIG/C3s2orlJOiq1nzqgRtJw4xkZfqmWdWIvZKFm6sEBN3PRa
WtzSqXIt1gjrT9rpPkUG1+yXPFO4x/YO3QM5cXyMYzeZmraK6aLOL5vmH9s2
EKeEEnALj0bZ6S19e1Aq95LE4ltmoedQmE80r5tACZw3HCwZ4Q1Nu1XT63Vz
pxjUc1J1reFXlANNZkse+tCulBo+Ntkcd/j0WcSPtlM7my38rdy+FnWPdk3A
tI61T6Hg8uM0JhxPQhoST36WziArcdnoFcBYRTab2hSxKCs/jL/7lUlV5RYH
hkFgv6aMx8QwAam0QACyw0pRnYHY6NG2emeE3btHVTmXpjZU08wsrQnzGLiu
WJ6m7r1kul2+jsDdUsUA1YyG634sHDEpfekOFluq0yGmfa2CW6EWHbmtsJqm
7yWCjly+wwe85apuGbGoQRiDOh6Q9UxjYtX4PoI7w94i6DOj8oe72z5LYfVf
9DhfBEu24FNKsw5VlugysMw7ea7zv9VVGf58ZCCKVErdPxNiVLQ/pJKY+Y+8
UGYz3t6sl3h9M30B4fLr0rnVuihJhx6e2wTPMMl5FB9/45w6rVPGfkEyp0bk
o+UTgFBaPBTloIvNVTIbmGV1ym8cSOz2LUXCcxrjBlvFDK2rAF6RANqlnDJF
mpNs9G9pg12ijXeSL7ZDA+PoeN27OJnqa6jxbumUxUbcnSt2whme5WCZ3L6I
RYw0XYmkFoEnf4c5b5PGDkZif8ZJEAvJCpxlT6kVmiFpXxiNFMXHYfa+DbTs
880jXWpNa4c3NYlSZ5hQUBq9zsHN2Jc82dbrsBUF252fm714Eqh0PEjzN/km
cx7Y1RVgm0ss2C0lPGFIV38qEOmwb8Gwkw5LNiIPZZ17W1XjQ+qzl8Rcms6U
z0x6BHbn/TkdD2YdBeeEjiqW6LYnjqYTUSBKtDVU61gmWPloddCoxC4lFZzA
qpw7YbQs0AAuweiLmuH/hZRJWUqpQggTCQ8ryNc87GEGXuTpZO9J72GvjmEg
Wt9hqNOU6d/21X5H3g1b9YLiI+xADpuuDYauJsEPNoInuaOJY3HfXN3lbf3u
lfJ+mEFhBVPhwznPR3yvdlLTxqt8zGG+hv8asDrLI1+bC8RhipT7dLhAGCxQ
3dvUpnfVm4znYjrNH+UnOLvDAJXSutMLJE+5GbwmQ+IKep+TCXWzqzdUNTtR
96G+Q2C04QO5SMaQJQlmZ/RUkSNWXA8Z6OoV4UqShPG6drc4mrXn5iajBGQn
eLQbV+kxj1NBAt8iqqSJhbmBz6b+GNb8cvaLcAeFhScws0Nq1E4pRmt7CQuv
KR14qO1a+9QaLjvIOsx4k0IFbtjH9TLFOmBjMUXIAO0vc5UtJzNYcFWa9WEW
o/IgWfDYGRm9J14hIrUi2ugOPIfIV5LfrTEtKYyVK8wcLtBmvGNd8GGP++x4
JattW4cL/onMyjRZPLFuEHG1z09rh6o9eSv+7Iq+CJUUSlmlSGHrfOQW3WhI
utUfTAL03tdYEiJYbaCOnJtFlNUwMgGJ01VsIfMNJIkulF+Q6J7h3/dsTDVj
ZHv4A6lPipw7b8XMOCAQoh/lX261NOE74dVn2MLk2BGIHNKqWVxVVSn7cUAI
E3nDCSBNG9sos8PcIF1BGCXsvBN9wxOeoMBMKt1DTv9IltgIVpFzhzmuJi1O
MmTrL60snVch/xhLng5UvnJeSLXSqNwwLXLqr+0GqzNkWdK315aZvmcmQWQd
g/6RUq0yt0dBjGV8McpZppTCZW+CRJjfRVc3q57Q4IgO2g0eigobp3S1DL8A
uXM9JdMnPJXHUJ7d/uN+60y76wWmd/+NFxom8dioS4TIMS5Dveh5WBNY1cvA
uqBxHqeFqWDFi7Mhmg91/cpodbXCTZ3tUVgXVHhKlzjz6GihjordF7RWJWwR
8QJeSeljFSKiUol+f08TMDD9Lt2VLGzSQ4sGbKup3E1CcHreGxH85C4w9oAz
gQ8wvzKSvmYESwSVJwBNBCyBW8OGfrThNJEiBNAMOL0VPPfN7UcbzWgDrS9n
1eqsrQLOilw/x/kW+XuEViGx3HGhSZOAG3EXxuAxFLENtMr+bP3NJZ6XQ4Za
3L+HIZyVVQLmmJbRF/OrJHJ7me4Bv7zh7q3bpa+hFL3RxLAQpKYiiPnVS1ME
c5eMB/XzePvugXC8dUsFiIaPCmEslHj2R9l+EEsNgfNP5K7C/cM9fWUT+XfX
M2LC9M2FZuMd1rAwE18rVFFtXhUzU66AZ8g25UCgEB/MhgQJ1wj+6SSsPXfY
LBN0gpXae2Hlal+5cFiwFgiyjSftFBdJDLX8cpaqm+GXlVacVxUAKlm5/BxY
lLwGc9PZ1wwze0jv7hz3P/+W/KoKs1pNc6yGf11JiueqLNdjogcHpJ3uMEOY
gESdvqxWNTxTuQyEZxVuixq6f7M29uuMqq+zgoHF5Xv/bm9Cp24Irb1jBHAO
3VVYDowyAneNE5DYqjbAdl2mBe61aCRd1Z2qSbGnvFw58IdySR9PR2Br2qRw
f8nrnK4zfd4FuPQTufw3fgK7MtKHFPjWflvdTZ1ZadAgvuZDzGPp/1U4PlyQ
nnx4JHrJNqVzaWEB+WEa8R5PNvqq4dYbVLn859WI4X23Eyh0KVRPIOjaXJgy
+fqeEggQLTPDWkBEsdJoUt15uFmZvtYvSr/my2pEjJWFjDluev8Iw4pUxaDs
rp4MsF0DDLln5fMuR1fagWJhnfTXVdI7u4da0VMk95Ghal0kHN2aCb2uYYXS
oOFIEubIJMJ8ltHJwAT8QRR0e0rgGVghyevuDjrl1FsmyaUHw58CrueD11gs
oFAv1x9W6JxnmbCojV4qSs2tCUGdT6zjFpLaO2JwEtPkKWJzhh5zJ2f66Oua
drwaYngq+lS9NauNVv5KNL1adMVJVVpUzl2sqpYj1TZkkytw86mlnxHmPrgl
/7ig/raC2kGEa6NHBQJyqBZbLCFSJCQEfkzip61QMBAuVTfqBY8ht84V/vNu
JCOyDPJaZympgz6ZdPnRCONgqVxGPkWBXZta2bKnP5uZJYfxxHlviaSimh8L
ACYWV9ScHwcBa/bMODbhDI1pLfpT3PLeZsnqdDtqNCqkOj8I0Kh/gE+SB0cj
YbAtdeLrIYIPmT+qtwXK/OUwFiKhd9S8GB/VoF39djDi0u1Opdg6fq39pD/j
okDQAwrWXQyqUWAJ3ZAmEAwz1lST3yJ+m01V459JFE/DxkIaGUqBZWb3qZKX
DgBzU9q4ms719mjhksF9r5OkOHol5rcdVms6jhFdDPnzlmN1FeeSKxxEQG1V
67VRhviHLlNXZwdgti20CbFh6huji1+ung8s5KSVCNg0y57MiV2mG174M0wP
IULEvYdQJIUbbh6mCabVMLc2NMrvTWDVSzpc1tAgT4O7BEpl151tNGfVBPBM
OoZOm2YmgGU+Mfl0JPfv45z3pdve+t80O5whWvRhRNSP9M3jLKcLBE4Pus33
L647ECNJjSZA2BqJ3ywKxIw75lANQC7lZHbWp3nqLvyjnjKpJBmP27KVS2Hc
Wyn+/IIYB2hsRYBBoauvlsOvjRihsSLgIBx702mKvonhLL13R5toXfUbuDC0
3AzoFHONKK8D+tVama56qp/mIJ0A+aKgZPyvi/I0srJoB9vMfdgoTPthfPPK
3LR1U1jNdqElnQJ/7XhZqMWm9ydJLpDb9LKgm1WnQoZ97SJiswXgBnJXI2uR
1tQaUKn88JXq92D4QToy87IMTIF3MFNIo/j6+oDy9gRWXCyBmCEuldAUid55
TRdVm4jYoPQeYJJ0TOhiIBauFvKlZQCM8Lf8XMhhCcX41XhH9UdkIinhcwdg
PUOzoyuCUqU4xSO07EMzNHc+/JvO4ZVT/sQC57laz1aK+tn++1OPCcjkjRC6
5+NA0alJQwu5Hj3Kf3DjM5nAS+iviHDa55OYijljH3Hw8L2U3YZY3WHK9H0/
hv3w+HxoL/CHj6RJLf2amFyBGe9/dvEP3wPIBcUXOiQXRwek1FPVcyTGCxEn
8G8pdCmmCbcZ0bqBgrGtJlQwYozyOvsTE+hrZIxHCoh8ZHnMjlzH2qySnIwG
w+kzNIkXRvsfCo4OeoHINVnoyOhOf6UoN2s7JvSaySLS0vPaVmU+vpikrR+R
AoMxR+Ri88Ebb1BF29ZlnDorrwAgLLPrb+JJAWjmfkonDsufFI+NpqDBKDgS
skDcMpefU1fC8VMca9ojROSztQR/k65as6XImG6EALt4cYTb6oXDVHhZG5Sc
wTr8Zxd2ZWyACB9zF+4goI2nmty+Mta+Ys6SAfNoECeloE5djE1TUB0E0FKu
TezkdfpmQRjfPBbBPqzuboCZGMWf4uyRhBmT1Jq6NVUseTPGwYXFvLaaJXZW
B5kYZiQXCdo89oTGMzRh9Iw3SAt1LVltaDhFYAZCpRJDdQUK1vbirk0DjRh/
4I2RBvijd/quO/Ehr6oYunUkGUh0pPBk1obRi1LAbbW83NHnxyfYxnc+DLds
++j0QmUPVWfi2LaGrnEPjLg18HHKQDPg1z2na73uTyTfSbBbs8hkRHemhnRu
9rB2KMot9jKINe+z86gM0uCGee9YoM4oHsjjZzscPpsBm9qTyX5o6wx4MQwR
llS1RnPU09T3z2lL4/lKhfU0BEENZ4TeYVtos/U8IDbpUFHXiRgCvSKnX1W2
0SpIGSoMWqkaUaM6GrUTQq8gpKCG6cPi2e47DXIT2Ok9QSU8AHkcYQf05Zmn
I+CJ3PHToG4ym9b+dngCLr/RxdSePCf81mhxm3gEyuXR/Y3TIIJocxP44zcl
+PqwsMkFMqxo3jtxemAmDo43N7yNnJbLBPugcPR25dt3RHoKONrac0nhLNUz
un3Lx2Q3IKQOTPi2o9CRwIflSd38JWU46oJZqgG5YuHj9vmEtAo9q4+vHjoK
rn7vyGlmVYcBoI7EOBZm11cBuE9ltYo8zZVhSMqt2WI4FjvxdHDHGKB+suPl
i7y9NdkwmFW8cv/uuE61Zu/PJMOFY2JLQwcnssUaVWnk+xzKHNyDU04PnfWH
wvM5SrZcoziWitrxjKuN4aCOaNq8N8zLs8jw7TljP9IOnYUb+SeaHeAEwLE5
jVYNnExH0Ro8ON2JfRV5rAhy15rdZosPjjKB1Bl2dAVZc16HrHu6gkcA+Nre
4+Z+9nwM6J1jYu49955ks2ScrJU9JqOuT++j6SbOgycQwvbtDcYUQxy9Vcxd
Nmqf53pFmhrTGAvQDPh7FUTsuwpuCBRy7NObKmzrP2NkAT3qNqWZJ68ubGMl
yGePSXUVpNf0uoJKIzMT3evtf512jSV10g7+MNtZUzJlRwf5AoyO82StPZF6
V1dZvKUKnUyTR1634xTgpj6Ohge5wX4TH1AVvUrpV1+A/aNiL2HLedcCDG6k
NPy3T9W3sO5It+T2YJq5uFKyl4hefWWZAW15qNXsP/DCs1Kn/iJla/TtrmeM
HR1lB7qFDywsFg4VNfs0g23MmNbKa071Sfi6HQeJ0Xi/rm95XBCFm9vk76qT
CqUTYbTiYjbZaYOI6t4x0bdt2k9UQ8NaQrBdZCta6F7ekK1Ut2aDMdBiYU4C
0oqIbh0/pVg+AGpI4zjKsRmkcr9QwBL7GjzpciMNKkORjWjFUK9DgLA0RaKL
GB3wMuN7Ut6gqOPaKs48qyb8OUl5QiTWZnPFaHYsZ/G5Ab+oVDU+6C5yoJOB
nf6X1lXTIzt6G3diM6zW/u/MTeVh4KyrOe702qtgy3/ROHCRXzlAdHRUybW5
BOj1Wg5Qs7EZPt9KuxAamdX/d5BWYAHBAnxHEsXo2NbFeJNw+4flYnN5IgT+
4VGG+oCRe1T4h8Xu8k3/Q+NQzuBorTvlLKolQRf/Rc5mLkHQWj3cFS2hg6cw
0qdflWBOvEwQOSY+GuygkArz03I3hKsK7V0hKQCsX2/zAZn6yURayzdROa1Q
nWmTbsmITcwbQbga9TtdNGMTHLJRQOCCLsTtpVXWWq6WnzpQviCpVE/eHs1I
UnAgFgKygIUpGAlpwGUw7sDf/jxRUyBjQ7/yXIObbOVuLzEM1F/yQhzWiNs0
TLtuGpeIoHNTCqzS9KWuvW65VhRqdXDY38YuuDIn0IEIVDAvwSUIQVyV1JT+
rLkS0R2OBm2dt9CvsiURaI8hxQriM8o4nJqWcj4W8EN6EeoEu8JE6JbY+/Qm
ax3mBzJIWqTRd/UGh696327IONeD37YJExtG2LWL7hUTt6nuEtmN8osACkrv
S026jFsNcvOnT3b6PoHTSp+5wEw4TPUPW239JOTktXhCdcS1P4+2alnqxnkr
18Gf8SufbZwWPGIqO6PAl3FJtuhhh/2WAyaO7rnK7jNX0YH9x4hf3COj+/M0
U03W0fLrX8aYBtiMRFIr8agQnUcXlM+skHx7gp/MEOqJBtNAS3MgzMF5XGlp
Z2Ze3uquMsoI0JO1a9Qw/tqi+6QzOh/HOxGAqLTK+CmEKt2tsnwbwtT6hhj5
x/ss2exfewFUm74Eqrgco/rDVyIOwyd0fRX5wFZtNekefvEddcOKq5yx0Ad8
1qsnBkq/BqJgDq7hnqhcV2xNT7LLFL3563zwOmCdGNSMRse4cNKCsSp/bkDS
9GyztkOBZm8W+vkVU9DIdQJBVElVQTVhMVwjtkNomg9AGLjZkwpaPCMbDfwf
Wdv/FyTQaghkYa8byv+yQnWOo+ttITR4TEu61BKXMFwOigntswEChfiHpFBY
XfTUTp6Tx9PLn3RmehIWwdKcxJKS0hsbO63O5pm9i2H8VPvSlPGFKhXNMhWc
lzFhiboAC2wuBudFVItOHBBw6NrPqy4GtSj9AZVyGx1F+LqpyqW+QY4bSiMd
xnqfb+p+kCLL+ef4Ozaxvt1pNOjOcHC4fa9U0NA71v75DMae4DhE++0YzU2l
0QS6Jf0UUFnra1bm6MXozp91/121jwOBv90uwdUEo+WLKaTyu2BPrURbMSSR
jwHXqdy+rI+aHOxZTXb52ovkOZxzVhXOtA5Iqi1NtfopBbl7liC1cPiw70o2
FwoXTfYe5wzQokgNco0VkTsgtQ+JQrr9oEM48x51vTE8C906lo/cEluuuEsW
+VkBdKxzIAy3SZo1KyltJWuRYZwVkGujEVHFAqg15Gcmc+08qggdSKynGz+Y
XfiEI2zjv7/ypQ6mtniQr3uGfEragR9MXN9mlCTRN3NUwcBsEnnSK8CdOf4L
FNcGS5wFqDOKhw+mx0svjs7vM8PjDDkHt8QoVZHggthVcIAkaw6fR3fAmlRK
wHq07y0AZFVNjom1jc0w4At8aYqNa8d6vdsemhYlma9/bz3l+vDt0roNCAhm
XTQBLrVkYAWPT9jZrZE4cEQZSETgRa0V+A5208bNtOciU3W8Uh45t0f5j3aB
qaAp4Bxt94d0Q0dgO8NyQB8zlSrqFO291a5paEWI4ul7lEsoxhI5thiGHw3O
Aj1ahLWUcdKIKUG4RldFg8mJXBlLyx9qhuIyADD2t/alA8cSGKGE+2r8m4bp
MrF/KV6pGbFfwWeMCZVUHrV/xTNOq8UxxdwEk9VooJKeUgB4e6BFrskiVsfx
8T1UCtvOCY/MFaHrHFXTHt8vp/DhoXL1bVzFkU0CXhUEqyNNG5+kNuetg/DY
nupO8HLAQ/3JDNSAqIqc45C/rir05ryVMjglEFf5eCrYdwcv0hFs+cSFP8QZ
Hb1eKrVjQYVrXRCaKUp0fDnZfZivVG8+fnXF7stUXJxtt2JDq9qzOuwC3J+l
+85l5DXyczlA7K2sVNmn4xiSskLdeaWU8NKHCS4YPc1mumYhk1XotWEvg8fC
YVVHWucSaDcyZZFKaeLGjbmsNK9R7n810NvcQn/sB7uZ78ooEPzdM7zof8jB
cOGNawSICy4KaOr/0lZ4iZLlkkFi63jxqWdkAliDMYi70/xrFQDaXcuV0PUZ
LB+NR/8EJL2m4OhPNCd5ryHXft2Q+KNAEL/h9q3IuQkkWWJMseK0fKYsoFNP
4EgG7LtZhvwyUyzBo4NLGmGxtWOJT6NhkQ7+cAs3J5RzgUtQ96Q3j0eqXfTq
hjfciAYv+DZSwYpsrQa38+l/gNFCks7woZWvWkMPT7VJX2PQ2LBtIDlRCQFM
QuN2cnjNsSjwZEWS37JtKSLYwMckSkxYBl7ea/AwbanVd+QIPTD7jmdOzO8Y
oE7nkTVI6h4ODv6nnYHWwTtv3ZNjXWQW1ZjLbnWB+W2oKDlVtD5EQ2bddjeY
H0Hk+G5yLANbHqdTRduqnIujfwYg4eJEpSW2/KN2mRuOle7ouvgYMSVw3YYu
rh3GeTrY4M19GEBPAjrA2davfHgVY5PPPMfJVoJmsJ8Bsl7jqnGgjAM2LH/9
p1NZcc5ve5Kk/poa48v2xMzefHj5CLO7QBdWNg3HGZjJb8p7xFqckq0dqlWH
7nVA+0I5QMQeFWmH3CyPBdhq0GrEa3vgRVrQkhXjfWVhqYx5s7nL1Qpn5f+3
mnDnmFBb1fHT1+ekQzXZ2OmJtuQUmBtab9I5PhcfJauGQxc8Tj31kH942vHQ
gRI9i6G+rodRv9vmndexpkkVYo8ZxHsaTuZPKTNzwbhNfrSZS9ziHN5e76Hc
b+e6RUu2cHa3VwUat2jH5wIVraEwEyyB30caK/92kTFN5YTbSDTOfYgtOQiU
HTRlirqszn/9Q4C1UZiGOFGJ9b1hz6k7jSvSErGTn/kwSQT8zx4rvu89IEym
oIz3o3uyEfviJzHjmLb7l5j131fyTvjn3TBwElV7mP1oSl6t1qQrT0jmojrv
6dARyZg7NgLt3naEK3KzwKafAMatJfQ++hNpjw8YGiWyX+J+D0b0IQz3h7ai
6Z0SOZBHfdZWfL1cmCn1dxkDzbqQ1Vj0N2uWF3sVi/k7Ko3qqRkcF+9w7rSa
ewqRBdgf4AvRnU6RP4DWsaSAKKjGqwXoIJqgKy1+nYwQjV3jx9M2XJYoVjte
3rEy9rcYMTD59J1tupf1Kc8q99i4sgFdxucxaFQCSxB1C4O2L2h+ofRRlSMm
aDL24sFmpgUNPbEzRgoCdqHvMyURtmh72EtVt95oGEeAOAh14DMNJj4AnHRz
e9dZrSqovj8OmItPeFTJ8Oy3F4WVH6hGTCuSqCTnwaTv/onhxlkjJXybKap4
dpQOqeZ+1lrAOuVf7UX0KlCNBjke0fNXVxEyPYHF27BVSAsvzu+fkaetZyF/
OVruD8a42a+7pj8HDnRy35KvfLoyY2XmrqQlvNJuFkiTjNVM2cG/iT84ZBZ5
6r4xV5QUHZBWjrue1DI9ygTEmhFm3zmv1mjEV3o+wPZ8JFMC4ULYBlzXZI34
mSstBYlSXfCQCGYYXhB6KFFPeLvSBgG4RlLtyiaZrzXDJ5YwZVx1tcFapy9i
ZOjQzNlm3pT1IoaEBe8GCaXgs2G+nHhMATaZ/cn4jV5oW/EWU9ebOHM+jXQL
EnUaBwR7uh3ekBMYjrDT5tT4W/sNbN3Jwe4ZdY98F0cNSpB+g4+qzJ0qwfnC
9BT7TLg3JA0F7EVenZesXx2oAAKVrt9iLTv7yfUrohtKIhcCtYsMxRWl+6qL
zTGd/kltDhCKk6jiMqTQvnGZMbYqEdQKUdJbUZfTf6jPpCEAgp5NwipeYOSJ
LDRF032BGpi7TS/CrZvIz4UuQPTH4ZFmyK8k5JWuVuP6K8rzxMyJsPWzPQeS
4px69vjpckFAs1kE8QHii8YVQ6xqcvl1zfKYM2503iWNJdc9IEQ+rTgfbxJU
DlEFuExf6giskgz+QA3l13QXny4mij/p/hjZxy4Q/TtPuvCQbJ7SbNFWzuDh
NhMdnjhmFQSJl5dJ6YIt1mkLrshe+XW9aE8momsIUvhw6OWeBDo8jKZiqZQi
3c8O/6PRhS6ajP6NMjXv/rprxLmZafhtlEmHVryokzaS+cgHnOBFBV23MuLk
NrEMscQbxugKN0SMKzmf1oyLT7IERYrQ4kdat8jpk3znzKVJNMA1wy4f50MT
isaui/9fo/Vw4VgSZSCh0onUcXG7lqYwVVCmoDYsty8KJnJY22QcDlCrJceL
IJ7AX23EIysEtWHB6xJL2D1BQSZZ7exyX6MH6PTMBJ0SO7eznkcG1vV42/Tk
/zghkZVIrriYLLCMZoi5re9kSFx/dKWgttpN6R4YKp+dXZM1NQnjnnAwdXwe
YvFgMpDVYWye3b3Rtn2NGdVHfMxHEFHQgxGpz50ZFTRZtHkXwBW00zRZyWTz
fjlzEhvlkxb+e8DqCQd/pMSifdxVbKzZh/5OZZS/460cMihDrzHjxk2f6K6E
fQE5XiyTOGoRUyKnpTPmhYrSoBBJuKKWhBXAILRSIvzomx6hhTS9o2wI6Yw7
EwCln3h/vkZ0AZ48/ngX30s7DbkZwLI3piTF1DjDD7ArXw5tqhnvXM9pG/g3
TbU+zBfWBM1hbZmKHfJYJ4+9Qc2Hc9cWxQ3InZ0+gDP5ZZ7Y7BeO8ADrdMoG
dozNUkO4DC3dclQPn1OBducj/AsMPbIVhJ1CLrHRR3/NXz2vrsLSVIxJ499Y
O0QSDHl+yK2oCgilTT09sWBGcKdFh+lShIwzR3dvkDYy3NcLotfmnjIeEcCJ
ES6wAG01j9Hv1zZiDZquI774GlT39vRvkuCAibPf5azESpPKZo3uDud/pHNp
hGrV9dQsOA0nPEgt7qAI8/+wi7AeueAGW6fxzzM+Xu+FrAUdeqT6KHgETPI6
wu8mEuKL+mMxXxdkOOlxoe5lTWTrmOwvfqC7bqMmUSMweIV939aQKeqie454
qDe7G7BYxkv9I+NDGx1fPGui9LOikjUU8he2OZeqDhe1l/VNyi2A2+vCigra
uDEBYfI/FITgZHQpijqn0I+so/PS7Ls88QmILykZC7mQPa/Vn74/eeucYFv6
+lpZur/CbewJeBwyfNgdpzUdKLp/p3vpisbjda77La3RbhNmymUKh/4hO2ig
uXTL7Eg2KTuDQai8EnAen+GQqmeYgoewlcb1Y4i+YPc/eGrvmFd0p6Clz/jJ
IVCa9vkREe0a49bUotSrv+RD1SxgDO7FuBXFePnPqqalhvWhvNFFwE2xiPE/
KssV1oBK+8TqvHPiOisAcsYJd93GQFMsCa0lnzqcwfS/lT17xCNPVrqXTlZ3
YzvQP3k4PytZ16CmBAEjkAsOGVODM7MHipF3fdHru98xLcmIJ8BWYK9jPLK3
unSGIi7+ecw9YCehHlS0ux7Qciy3IF84gahWPpTvRjVhowhYLo1ph48Nwlma
YvCYlnu4e0NryMinVMXvPnre+E9Yxv1k1Wwp9eTAZtjJvolOl03opimkJc65
ALRSNJ5m2OxR3XbkepZAXkmHpzoik/NpOulruB3uRwQqY/XOAJAtXxRb14u5
pyHlFVDJPx7eJ1bIncddJhJpAWmm/9Rk6GnuHiqEJL1qe0XZgHzx2ZWhe62M
7MuPZt+ol2eKGxlYZ3Mlt9kXd6jJpRjsWCSR/sk+wWLKcfyvZrbPqGcHNIEE
mpy/F0kXv+xrGSmChn+5T6EvaDQ/cFunChrzzraKf85f6ILzN6dmfs6QQUa8
/TJ80qxWt5cHWMcDAkYf4g6p55D4bWh6+UjU+ke/Yi0UqTIIiZ7FDPqLCtgq
tyvS3KcJzb4msPJrNLk95VPCWHm0YE2uiDe4s/CTUtjDJyd2WKGsVQWVak7K
/NvTfHeKUh1CXjsy+Hvk3CxbmozKo8Ha1n01a5xc3otkGkey05/bLK+6egpI
uo9oMO3Jpky0S2JLICBH+KyavPn92UlSiem+jvwf30OQSHR2tTijSHNUzNDG
cN81Hw2Gr6JVZAeZHIL5xlgv1CTMSIvBDMjdvMnX+r/LnpfChRhcB0Ea0CL4
YEL/9YtfpxfSLR3lA951QZ5c9E66cs+HWzTDKhVF4HxAZN4r8V5Fq24CNenY
A5klCXrEcoW98c2lcmCcWdZ0W1pD4PrBfvxXQlc38F7AT2dw9BrTx4eJEByG
5EXw4nGijTZ9EmkPwNXWjohM4TCoSMx1KSuFZcFSo2v3VA/LmrS+YW0CvwJs
n1JDWbn4DK5XRxvd3/+WoOuJCHOFxBGA/EYt6cg7S/g3Y8TPYgDE5E2tThCZ
mJ9C2gLucbuGI5uwY1dxWfeRRYqzJ6xip3GXu70BYIvOQ/pVk8wHpeWnj4M0
4FXbSVNREASlTrgXlQ4INEr42PdK+SeWqT2aoiZMzt7JjejuiCRXC3IvRBot
TinuGTrK7lKUCCM9xpoPTRB3e3K0k2nvfhFPxQAXBgnYc10EhAFejGfjxNRa
J++HuAGskqbWdKYOqye2wkJ0kW2/EMofpWsn16g3hnvvryATXf8SfKzZZv7G
FILFINmTaBqQmIPoVYSbyBI3i6SBARLZ4E5CCHZogSiZ6SbzU0klJNoe7Fod
/3/2ZiKJtZNeevn66bmLcwkbIRjBQsQoP5ApEOGTRWg5PqDIjHk19hMd9oMB
Xx1BPBGga7+PcZLO7Bqb88Y08D2oRm1kFINCt+ZmLrtmYzTnZwkb52lLiWfZ
5onUWsPJu2gw/+SYhSsYMmmofom+/Buuz7IYbCdbMBtDEW+XZwr17ispk8QC
yPgWrBglFxum9OQdGk1yRGgXCuFAIe+7YRw/Bj1nzzJqIJJJnLfo6LnXA6Y3
IpA4YL/fkqXLlT7mSnd69q//g8WaAV2i8D1i9uDgCfQVNcOX/Tpg9cAPx+j+
Ah7vVP4+R6QRg5TsQIhinJxn05flyYjLUIvANDuxyrVu0esSIrkElp/Mp1Kx
KgPLLiu844NO7KSl0lH5d94zqpVhIQwe22mO/Pgouf7qLeUIZotOQufHtkSD
HBI37ZQca4FOS384fgcE9N5SEN+bdzkMAjTysDfnaAXx9+WUN32Khr638A0N
aSEE9tqGgoVLkZsRiRDR/kTh7dhnx52uTg/1tTmPqcHDt8zQ4M3A5GkkYn/+
zcLqZuuLvWTuE1F3HVFWxBJ7DRdMttx2yZjYz/cR09GOrKS+5SVvmyNV9cJX
O6nWFnw2JBwqkh5E75WF3F2VVpUkcE5XtxLcP9XcMnzhIf3w4nVLRlWZbWoL
GAWbu1eXuwcc3oQk3DFfY4bxfJNgt0G6APPXun/E4Q+q+EPEERt/52Bavy9T
MQuzONyysycxhWYaf4CbJ8PLz2jjdRyCYlOixTGqrZDX00bY4ZdR/3KH6xB0
1xYB8f6JDgCDUNFamPX5/rKyLaOtPpb3sJ+OxaH69nfFns5245jrCvODM4CT
1X8qW0veT2HFnS8JgMsOvs8vKcZLjMnaZvL9Vi7j4ZcNqC7pJUXJ2mXGsNRK
GibC08UsBdAUSzMb7SV7ddMxATjm8JoOlWQJmgPqb+rgb0npozwZ6vsafvjs
tB5IAe7z60ut+aZbe9TeAmrGRJvFtZbi8/ML/GsUXyBmQmKjyu/zS4URT81M
ef+pPqNwqj/GH4JNw1+M3ohDAqJBl3OObT2SvCWQlkcJgWatotsBNFK+A4tc
5N7R3Tl0PrO5kfj3KmRfPOgPUvv+1orK/rHsCuJkpWFtN8W1LUTZjTBHsBrO
/RxLALJBOx6Y1V9Sn93A5fI4gsXAWV1TXhzkU1spr+CRm2mq6BZcNc901V/B
vkpgjEp2tqhwCexvg+33RNL1SPUzPeLjLn/89tUXdJzG57onHvxviUzfEr4k
qQ4HMbo5lYVuhFrfPQNnho4oVo4mzxzg1N++Dg+A2UyX8SrBXo7dV5OcB5Pk
yQFYfyUJUMy3KnrvpHFO6LByokD902xhS2R8R+FSnEgQDBoI9U9NBkQIHgSv
azGC69MLX8TxqTSWlspEy8U2+DsONyWjZORHDrJLTpkDXfvePny6nAAOxjN8
E3tj+m/OhdLAXIjIKziVu7+D1JSx6o3u34Xadf5zmn/E8Y27fGoQKw/Dk6Bu
vDIzrzgxqhyf2GR5mVZnx61Etjz+PniVWTfuDgiDy5T0fVrp6ZbWKyJMUlYK
FpG1PdvMBvpu3vi4RPdqjOj8E21yYUkX4vHnN3u+Xsl18CZHn2F0k0PfP3TO
R09IqcSUN5SPaOf2XoBK31oTd8OugjRQlmulPI3nPM4THTEEF7dldDhiTaz4
fAqj8dBMIbn/xp8+LTUHpf5tYh5Mm28D2d4adCUP+bNAdD5yTb9lBimak9xw
BJJ4CC/p2b/CpDVlj76vjtpU1fg7NzDpZAEuaz/e0xYGVb0TQ28CASpRtUM+
/kzm8RiI9hNZyifpgSWbVtJf2/hu5M9H80PldpBuNGlpKGsA1HItYiDqTpYg
iinFFJ6ThAqln+/Jaiv57JmL8yCqO+t3XouyZV/lqoQLPXDVOdE2W8ytPhEY
DjqTWj3dWJC4hkb1t/n6WmFC0EPYcgXD+g/OxpJLfsFkavjeNYSznPsbaJDf
0k9g9VEdWM1JvmJ8POmr0CtFUn9MK/lVQG6SCreDLvj12R/vaqmVdVYBnMHg
dPN1HEeZuj+II9brtfw7peVEXmBs+CttmJOX0huf/emb1FCndBzyYr7b4Etj
hzECLCdCMi9m5XL0PkXVgQ8qFsgN7tv+5eTMu/xQUDVkmN6pOQOqirsgdBDi
SxKrlCxru0NOMAqqkNihzJvKT3ZOMWJdoMQX8eEjv+IpmGU3LP6unjzH90wB
SkQauhXNJMlKF4OpGsTGpjlCfNcb95gaGqbhARJoW/UjSDJynfyPYqEKpya3
5NJHVNte5O8sA+KdVwkIMSYpQB2rMHr3tM9V5y5sMnGzmmTHaS8xHnFvXtZq
88L4s82udBsu2RUsBM0LxWTFGcyLJ3ABm1ltAzLzjzr1Y5kaD1212naC2PZD
JCMhSn5X2deWHUdab8IM3MhUwyhYfpTv2Tv3wtuF5yPigSFMWqtGYm8rpc5Z
Rst5DFNopic+3GHKC71uAIH5AyCD1OsM2NUS4zU5zngyHAic/9da2TH+BDqH
2H0mQtrvsuFX4mVT4McpOa1/5pqF6UJZEneZlXPU3qNcUYQpjGrPEHIL7mNr
/HExwbNuz5NSXT3fZLkWKGVz+UD+38UK9faFKaQC+6eagmpeS1FKaQfwYzOB
0Wx9nQxjYmb/mMT4qLm9M2O2Ha7eepREnKrE9LwONvGKt7BSaseklOnU1YEX
EeiCE34YccurHLWNAOgnXsFM+nBJFjPtBeQZCGClSjnUYsfrGQvBwiF8V8Ft
mYTrsyRftDXt+lj1/ypZs0iQSGTnQrBodASVo50YgQjLeOifL0fFAj/vFeyw
op0yiWWmkBj5fgJc+GnVF1sBIg6UIRQ30WM5K6oEoTs0MGUHCjxh1ynfE3x+
piuuKpo5DiIegBCHfCbLM+AOuK9if9l/sZb0GxdGYkxyDjJWvqN9ARl9L/Hx
PcPPVu0wdbfEorSW/tnEXxFB9x5vG5WGhzN6SdatzlTI8bVthXk5181SkFT4
8qz8LpmdSirztHU2qqg0wphRS+VqnE0sq3+Z65P7aCp0Hcxbki1djsRvJxmQ
QjKYaL+M54hjAjFwEoa2JBl6Sic+Y0+nmLGmsQP0UzKswov4r5Vim2cpHWHx
lgPPKfjSqJ/PfRBGMVNpTdWZM5/19UTvTOHuijRh+Fm0JlWI3Sxsrh84j6JC
6glp0o1xzcIfFxEe3Eke6beJet8SpaAbU4jmDLVQh2972sFt0ZFcf2M2CFZ+
J37p48V9gBIlRl2S0xv7v6hjYrfX5oO4j8SwpWY8nqK0F7Fz52ntza8Edfw9
tixMG5raiPqplUPpAUA8kCJX18O6pEqH99rl8EWvPChCdEimO8BEJwHtrxjU
GBPRRasvZp1tcgGLz1SKtSjKAhHDswLS2aBTrnpu9cMTpZ9x+pAqakPvIDWG
MEwiP4KDCnnyWV8rak9cL6SVF5xnWlpU27/ia6CkzL3kGA4ADF26PkGjvwcf
lfkZRn823gAXAwh0/1lXZviKBsaZTnJPHOAgglwKOs3mkvl3w++UqDmTRMBS
2GLkFqLv+wFFWNovSJ9FBPc0bbONn9qFIvMmIv7NE44mxhimDjq8Nz92RgpA
0EmvZYjEJh3lUXV3TLPjEKeM1CwsCuvVuTZn+nhc6irzvAvGlxgeecfpwBgD
ZkHn5YwePbEQ+2cvjbWEwILmp3e3FkPHrTB01A03T5mc4VPD2h2u7zFo5C5s
SAJRjPjl/xFITBJdwWm1TYp24tBtW7zk8o5ALAT9dg4TkfOtsi9witDYFZd3
k55HspQnuiMLYWB5x8AjFjQSNnnmdRfPc7PQjaYGOW1X1BcBQXgTZUk7Fms2
ANfa8n5UtC5ofE7dw6CZVXL4ek3brzT3JLQ2hgqXh6hcerI/fm0biF2g6ycl
w3TbKJT3KiiUXKRvjwnr+dQbpkIVeAPa61Sm2TaNV5vfyxFtlgcYzaBpzPVG
xg0C65BjBuDPQDGJtWpQ4UIR18OLrN016TynZ5wChd3NMxso9i0EsTdrFFGq
m4Q2B+439diZCCLOb4eZNm2SmFbgdgf4PsN2aL51uIapjCjUcskdAJiWqSsD
h18grrV1DI+I2GsOHneFDMr2QpTSTyuPajIfcogM74gj6BN9RTfMMs10jtex
2kSld4xHR5/ktJ1pUyRsCI1QZWjUUJdgX7KmyabuD5Y142Hr0aEpMNuwwz1b
E1JTFN5xS7SpAB7UIWztPmlx69uFFuZfgtAGbMxVa87aC5y+im5lrAXVhiVv
h0q2ERLw6Gd4bVNAUK7/lUfQe3d8tIjgeX0eEI2MoX0QhoDWkT9EIeTdicw/
d+//AqBxwOmOfP9/RiVsK1wKqkE52M4jjljH/GKzkE9Ly8wqkUXW2l2xGvHy
rShGU6r0hUXhf/aysGakrZgnZI396SBwzOFsBw+X2EZ6f7GYV6A5dhk3aLmj
9wO27B12KHqnpAYzTBXhFgRnpu0sZvLiHNPqTwrPA2zqRvq0xIcxRuJcfm9x
SlxnE6kKl7xNt7QSMphoS2Z5v8DdRW6z3qb4ve4oGfGKd1ymghT/PEdPR2Nc
I8Qo2q1mlZTwEy917kJIyPmmnGmielIGRyplTUxl2tnvfKwn1yKFXBYTTkJE
6iG3QgEVdeDzjIpRK+AU2f1QMcrKpziVgP0zUhTys7hYjIPQNrebMAKTqa60
I8TgiCjv1cF59YTzt+OT16+iZF0nLiAAAUh9Xz1ZH+3VvowY0DvGvnf7ejTA
TbV5LiYVX+VxsSK9ipQfUZZf6N8Glmo0wBo++H3IQwmTrE/LXx1zbOKqpu+H
eKTibcG+Fvhe2V6bMnVwAhKQJyTsGF0CopaHrn+H3G4EpElsIyOqHnv9Vj87
Bt9DXpm1sxlyMhmGSC1xHJsgFAC8wrZvMoPZN3W6xcTmalqH96FShPYE/Kp1
v3LkaYd47nXBwjWJdZQ4TBTXSbfGTF1q+P04LLdVdGjLI2lHtCr56Ahv9w8y
72LOfcOn/Bh+zpobVK7BhlQ7aacZ0G/bi67Vg3Vv4kdwAb5edhaZEIbs8Vtz
xdlSUTFfgqgf2igU40qTuj/AcuCscnOH6ggfDZa9Jlonjb9HeuYgzm53lGeJ
APnu7rU/AE4VDDyfxV8pqiGgQ5CaYvOzgyHYRKdlwd/opoKSK9LyXZoqNHcs
aFiccwQ3AskFU9yxE8JQcrOkc8i0JqhjhdfU05dHPi6JPqQlgEhnr8uBQo7e
iqJ/SbAv1c1kjyqWckyC6VqbsZ+S3zMcxXk5hG2mKhLb74cvG1xhcrR+sBE1
qfw9I+OcaBwyDnJN90IYvIUfWZMjaFp9a1xTIuKSaXQjY3SXpJr8C1rE6+0M
EhWqi9Dna0h881bfb5k3uUwXlNZ9wwm1O38tSvKHaGJQoJnek72Lec1pbcS7
UIb/GzF1XmUPrbLvbrzIGUGnUfo5Kdt+gG06XRXiCtK5xikGTZqQ0FvYpGrq
ftKulXA6u4qNrcqBIBLqSHzg6IFpUi9Oy1WeCW5w6CsDv2bBSstoAr6QPVU9
SBsmXZBLGayk8AZQ8o6xPWnQJqUf3RH+AQlwtjCPWfLBZ6kSsNETW7+cK+G7
GpXdFIGAEGysAzs6gMsQyF4f5tUNVi+VxJk01xDrxB+1FPoyGqzJW9JeHUHe
XxHKpBFG5PvBA3lFkHyT0c5aKnQIcvtOyvehiuinE77JfK5quH60z6KJK5oy
whORjIuaVJeBvPb4a4JiYY7VNiAqMWbSHl4RlCCfEmjde3+rK6fmGpCgWErN
q8sTLsidh7eCd3niGD+TiFjRY4CuxA8oARFSiSnNK/df2lACr3DiQPm4BYea
l9dAvQvGPNsWMQ+osq2oNBi6fgjAPi5uIbEMELL0eEF/zaGcuFnnYHYpPrhT
F/Ei99d/x13glOGo/I/0AuDh/8e7jwEwBNoLgrhwuoXpQtQL7/8O8LhpSd9Q
XcUVNw7SBjDpxZDpiI+P4uBWfx+P34QQML3o5le0JIFHXof6VsH9dMfo5l3g
Vyw7rryzuOHQuL5kKDg30gRgcLC98LcFpMa7v/1FfUXkLTyQltXXFGhpEWug
R6PL0nO/v0rMgyQ3S5HGwQFc6XU1Y8S8lwB8tHDcPcRSK4v1uxqkzFICgVWJ
oCe0yoAidXHANt4wfEtR5dDL12BFsZb0ZiHYx+qDLLEULbsszYM+okBX24me
v3sBsdzvmZ6yPedEBI0DIbWI3bX7nN9v7oWByk3GJtTdjA501QxM6QlCWHmw
emnXoGNcIQye16D+yqAQsMVGq3cvoDXD5H6X+jNk7uUciylfVJ/h6TJ/2e4P
enx0n0Tr6JYjn7XdZMAZE2CP4D6CZRebuA1bBzHz5dyKvemxdaJ5VPZK4UOn
d+qsLwQuUGvZ025jkcVdkwCsQrAixzrk+2lSW0bfg79PfFphYoedq5i+9+5w
InXvEa81lBrGgfnSzeuuXyT0lDo2skcl6j3GRSAW4HYEwKQ4ICdDF5JfmEUK
N75OlmouAB8ms4t0pwPUwYSnNGgu/7LWZIfvAiCdRv2CtHTtv78z3KYa5Z2i
LhVJrfvwzlWk0Eo7olwOVaVK1dX7Wfn0Xg8Y6SI1XHryJM/uNuDQf/I281+A
wS+ozzJJJ4ffGfXg9EH4oFAvtc46nAfZH4Ykx//XSHWGK++jw9TLfZmNXqxG
vn0kSMr9Qrngr1Nvbp3vnLOlK05JYTA2aG0D/VMxnNA+/MGeeRVDRlyzZXye
KE1VuG2S4J0v6VRXKvjwGV27qQWEN7RsOpdMO/QkL80YTFftH0wbrTwckqiN
/fsQZ7Vh82YwWm4wpJY9BLwKgitdJ9cfS9nBlslRh2cdnfeYUfK81RpHYPgY
V8tOH+lVw50xWvtwHXx2k/bRzRqMgXuztohNcgXD1+3MJ3ZZhbgCP24GU3+R
bUQOVenfxdqUW/rngYddQwprUcqKiEwttdKQ6WhNzCgRuJebcVI7eSZbMAfD
fe6LCyHgsJm2sDv8loV/Xedk0x5x3BX1/PQl7XsW8+v129MORH9NrakqX8DV
mCiFW+r/WANCodI+LjW4kR8UTjComdjUuVK4z+kCjJ7gz5BoHUfLUlEHlfu2
H8xwP/4HCWjqgh3xfeHqMb++sxO+GiE0+jT/OC6cgmqhuG8tMrX8v7rnbU9G
zj/2hwowrF7aH8jfdy5svYbFLuygALNIgEO8ABXCgFyeXdRNhzZhvXOLHKR8
QQ6ADN/1SpMNyKr8kaUGF45ENkvGk/ZQ2E2NmVUiz4iiXlhTje0+X5FnSLcQ
41hSfOcPdjKL9OFMD///kQE2uRKE/GltCTcqCsaZijrDoJTMBz7iG3p4W/+h
rKQxiauxKl3cm5AKbsBka8RTY5MJjRgqcpcQkHanxZ94ygg9DuDnjEwOV1gQ
SQleRmwcRLcYaUUX2pxCArOQLlB7W5PLarOOVHcwqZg9hzTykaZmYoRXGBPa
17u9ruQdSmMzgz/QwwMT5NJ9s+2moS0YQYFAbn7gqID+8pYMfZPFRC6PD4F4
dd7BHuzaNSJCWaEXrbT7dlS1GdvUZxAjnXa7cZQTd9NTyQ7mI7oWnBR+hrNt
RJSHZD50y/1kLAAkudiDYAj3LdMvZ7VbkqcmwD21E0wk82ccyFdqUlJEJBHd
Jh+KN6gdL+LFvcRlC5I2ZmwN5sB33wG9q33UH9uB2E3H5bWvlmNx/RSbiCIa
VgdcMjUFK3mML1SlRQFJMarp73PC0qLlaVM/lc3nVcpeq5sUlw0heDPKdBzO
cSs9qMbDUn7Xgperyl1hfRcdRDWvsqd+8UfLcrJzNB6G7PAJS3q2oGlMgwR1
SWNicP3Zy+pm9/lU4E78IhxEQajGwpFfJbN4IktoEJqYiVGpsbfPgWplqJfr
gWuzxQuDBw1fvdv9r54SzpE0cqISyOUXozIuQGXNivRRwvyMnfrfsbhik+Zi
jmKzIWF3w0BcRTIXyOgmk4zFaCuOaKU+MuyYmF6OZMKcuN1aQLjdnZ/P0KLb
fdKX2OZP1EozOtuWhB3PSZBIt+3QzZWMMjNh0bFG93rq5vofPshUvvh9QAIW
HB+CvQLs7gHSA16XOMQMK2sLw/sdQW5vqEw018dKxeFqDHql38RDz/OYOVkQ
ZhdcGWqyXDMlNENONQPQqbESKtauJJPhInEfqxqkke9uVGyWVHzFhMu7DabR
8U2Zj3qNr2S+nN44KzsUcdUqJhwnJHvuO7WvLf8uvMjj66hayG8iyD1Qz7hm
kgKYAT3PhT//QliXPzGQUb30RWsNUKxtEUX/bn7++yBw2YvhizemRIpdyt03
KwWeIW7A15uYaaXWRL1PuxdwfEl0u3qcuoMZXvBTlELu0OJq5NfVHa7ebylZ
+cSOgUGC9qdwNm+3eHC7Nobr5MGSTwsBOpSta45uw2URdF5b/m3Xk3qvHeiU
iX+jkvi6ItoDXBKJxwC2MbJgE9vypsTznaQbb8xFnXv+uYm+brZ6JnXpdWr5
30vixFseMMq8DBcxHOFb9/9pKN+oBLh/3Um/FKBq6mhKKP6ixTWV/iw+ln5N
0yytgJc7HkYZSmGm2teqahEuxbJ665buFIh7Uy/knLsCkmTGzOrkkMPGaoF0
v8gTreeebCf/z9wpdgNVNL37fFgvBoxEndOqunxOH5UvGJbVmIBhymr6c8pd
wwWN9KuHzw6CBIKhDpdwrO3Y3goVUBODZtTwlPMUAF+RUVcDPHk8HBbEiEUL
01OVuZLkrZ8GSqXHfK7XHbwqTsxKcZEHmDgKvib+uwGiHVcoQzaSJvHnejiP
6AxGwuSwidLmBLM8sNcfVae8TY03pWdG/pFEB8tNZGLmhuZEb4pAXVF2AI3r
D4RL5tu3ixoRbebLSLAKlzl+v7emuCR0YbHWdR9j7SbhRGlZAAvFnl1+/nAg
CKd+IFHWoblK08Fp5aU2mndg/RtN90yZ0NAmbsZfMZ7/8dAAvEvumpOZQeGO
aynCZkRr+x7FumUsUN08EfGmukiki72hvmdr+R26Du27WEhMyLZ9sr9/KwMB
vV+AHvNt6fNEZ+TGwwSjNuh7S4IBpTmpfPR+k8Gwr/q+Sw/88QcdFKHLqKVc
roFSm7tlrY/aBBwtYMMfyo/9oBbI3RM9FBIE+BJ1PccYRWgRJkkPkQhtbO+K
wuCKFqIOQ/N9jiXvTGojNrLHd9y3fpPAt7yjwY3KJXm5yTvrFCCwtHzM2gde
pZkRC/5wQwbS3PiEJJo5NkXLBKbDjyMYbRtzbbfKPFzLyq+vkbXDNheK/gRu
XAhHbxe95NzfgyWy9s3JtyqUKnf9RG6V9PHv4THjXZGS6L84/NXCbG9OcrT/
muzXUlqo6JB/W4c9bw3S774KThplI2wTLfqJ62TgvlpBiYkbf/LySFO9Gd5U
vKT5K/67zC+9XwdCIpwFXvaBf6BVd97sOa6eKWNvP+/DyDRwPIPI1WY9Yczq
mbXup3IS/tbAzRrghV8aD0EVP5GbTFDhNjV79r7RSrlO2jZe/LmwrE2hk1PC
U653ZofpZWEB3XZVh5WdF5qph9neB0PvWCF3aIyfyFSJvq39npCrlYhDkKfQ
rUXGUEz4s/3zruRCWEB/yu8nqgtNLCLv4OG0jden16FxVUSrSDsk77a2fo6A
D4VwrN2xRv1vimYBCXUb4jMPyWi/FdQUlHdkjyTUhus/zR33zlCsoOTMr+8n
4FfvcU/eJVN1Yq1E4U2guSZ2w9+HmShd1VBVAVLvJ7E7siKNvFlI3pICyM6R
Tl6pL6RfYhl36v3bLMO/hFpy94AgXGVsq0lgWE7j5OgfzeFMIv4c07U5bZAS
QG3nsBqBnoJBYlld6QK6XtBbLQcZ/LmBM1sN0YfkWAFiK5+9hjAa2LpmxTyT
zVKq0iwiXE4UGNTOw8XnVffTLGd44IOrt8is+fPqCqb10gHQl1jIpiKNPCvA
ENYRxZayf8Z4+8VEI43KBw/fdy1guVqrg5/fFoRjWNcPmxmNgvmABM/UzhxY
uu2ad9LOB/P785wEbmgJwd7eTbhFn5X4lnvBY/C+0lUZrEPvFkxD9oiaGLF1
CCyoMEdxHz/WgFbJn+dSIWslvFWu35XxtScJYrHRGNjZfDIUMuGwm+Of6i3G
5bs/RHojxhKdlasg/rUu3L8jxsN0bmUiqj2N3SlTG57URkP8vKFTmT0sCS6E
O9FPEUPnTBRb3UDoJlCRKj5p54xHhHwgHyMi+rGYazzv/kPkHls+gr7ggfLQ
Cocp2Lk2qXeacrnDloewrhJ+NUej45NB4uoMVTN4B2WNRkDKcT5/GfiJD5Qg
9Rbo51m1PpMznGcr6dld5eg9htghd1dSBYPWMNBh6ls2AIs+olN36p4A7T5F
89RrdxeDqcBX1xMUK5MzrDIkrJM6WtqsZ6uVZB2QDY7sJSQa4eAM0+Zi7PiW
PrbnNLPYU4f+Ts3OrUPaQeBnqazbb7cor/N6vKT3X9JnPjZhf2v+mwW5Yz4u
nasifT0s4JGq5P+IoMFv8zQsSeIkZlNvvqjEBi2rohme69Jkb1OWCV9lgXIU
uU0VRoum8ijkBLnIajSFh2Wiq1TXETYZhMqf+7zjXTOqLIwle2xRz8unVlGd
QaJXS+s3UJykDVNMfKbUlNmzBTk77w05UgjWQoscV1/6ewPEk5notpd3fijC
/j6DNo0CrI6q+UFzxN6BP48VWKpaTF0FFXTueHUv84RKTc5AQQ3xXsZWOQXB
7r2EoW+oiCsBtSPo8lbDO/+lJG0NZCdQe3R7akfKue3BbeVrhg5bO9m2Uwn5
OsU4htOkrwmf6/OJ097ImGRY16coUNyDn0jREBVcIVZANtzOCipQYHiZzEVE
GzWWyCLsTDyPmjtB+XGS71vrhLZmy/vXHrhmz6gORmngcMZWpR9y7CCV996m
VnzES2RTNgWHq6oRHPzkm+7ODC5M9sLd/uu/khaXm2cSDebvInw5VvKntajS
MlCPJOZfgP4bCKbCMkqXa8rfCyqku8hy1qLb9dUoqCAQCXPaQPQzXz4Y2SK/
iNOcPS02IuHpNPfJcQhRavVSwMOxGpiaaC4o/um5dXK2hwoQTFzI1m2UmfPK
50wxoc3nKPUi7nvAwSbyopcaRHGeHrRWK9mesTaXRUsW1W4sdUb5m0UrUa/8
gavsiVxH/quuVSBAwjhSnIZo0gr+nTwGEenhnEvlpwB8DIu7vhRluAeqUIeA
R+tNByJ5YfS9g0NJ447GkZDfHRurZ6GUyetJ2sewOYX1pswnF7Ok8RPTO0er
ZJ8pBR8tb5Ha90O7a30vZOPqZhMuMSBW6wIrOsJWTfGxVMCa31eOhFh8/bJP
JNm0FhcuL4E4/bfBqaM21dfjzWoRx5OUu+D02WAHNT1zJvJF0OWtaY4BMsW2
a/+rLYAS6pNqY28o3iyeMVYofcp3lSEYvs0t1/Ozfmp7ib1cpqlvQjh6YIti
61UhUOlFOXJFYigKDTk0NR6uCeek0CtFlexcWt/SbA0EvcKycRXbVpfZY79F
YVg5UL1ndmgvESfRrZ9Jr9LWY/qejV4aXc/F/gUtPoOAyL5TI1jt6NoDiKji
ukH3Yqqh/mBTshOPa0zTvl6zGNU2mRFE9DvH8Ay/+ZrdGU2gvad8upV8+WCD
D4ftgJgcKQrfndF7yRq72td4cpF7GhqJ+qihVzsPvcEI1a9uU5Z63VFiLkZs
UZa7HimZd1aMpkbKfBKDbU70ruN+v9vTgfU+AypJLKe8pY0ni2hMpaLaafi5
CRSmw3wuY/U3nmRWj5dimVwp2D+I8fO+sXKhGzIgaXi+zEW+a+qAL5cenI8g
AtAdGdkLNC9pHJVA487oKqcyuS0u7dNO3CafIlSQXtHRULZmuczLeYB0AyxO
prN7zfI8Ths0DofJJC/BbR66N6O1EW0BcLalKT7tnLJ2hEvPbU8G4BS+KJtp
xQlytBGOHNcArla1ICZwLHcfdeNIMrFc39ykmF/Z3VIQvLMQ3khjHkfkbrAu
v6zg5Ph6KU0PAobH7sEBUhJRhvyp2Vdj+LILOg/HnZ9gbBQ6C7cfDf0rymnr
cmnzg8cSxPyp3w6lBvVHG7A8+TrQpTlBoKRLITjHj451bRwsds1SYflIt+a9
+QSLx5OdlNJ50vsfUxiQ9AgECuZKCkgysdGEMYr/jDt52Y1lLBNoZzYdxK4w
3qitfqyAfCe/nz3efeIlcXirAIpVbISHNiDbC8NPg0tCdHi+oYLz+Ryt3NNO
3+pHNhGejlJ7DQcxy50cPRtonYdg/i1JZ/A7aZwApD17d2paJuIxJV/l8JK5
qI2hPkRNmK5s6M+ZWqcVYGTZ8jKEnd43WWxvCZN0VJSw5GrCkk2bQKp7461n
mADzNrBqUjne1ZBG/SGH244e2U2YbVFfl1S5fhVpuuy0nKgtROcZO04j0uTm
bQ8LldEtTb3mh0/3qx6y1Ub5BqH51+fYd+awEu9QGg9FMLxfatIZZKJPelap
hvJnZjjSMC7dAjJD2QtvjVgPEy1LgWq3jzMWFD7cbijPFzqo2cBCRHy3iKbX
x4ztiPKZuBFn+K9v0JxDzJsz7QRTdjnqp9flV7DKdsNZ8M+3Buq68MzFE6MZ
WIxVkGXXSFrYHsRYO5zayODjJF4WuxIm3skG2a5wv8BrqBxBxCAP1kpezPyL
Pjd5NXRhYxMec87EgvgxOMl8olG1v07hBwCOc7F9CWUD4HVX3+r6FH8JP9i3
z4Gj6hYiXsWzMh5FA9ZzFluBG/kOzOsC7WBPtyDyUNX5o6rbYqDI2d49wNCW
XLU43TKx2w0tNNtd2/ArikNwAGfK0lcgSMY/LyH2drBr0oh4vFo2/60D8Yox
geuNhYWoYOi7farh74D8K0STPix5IZx/KVZaoQC5gBtbl8n+FJimopAynKIP
RIGhFO7dgPysqNvrfCnW3cLvEKd6KbV7+Lu1sb2c6l7J4gllkcNEybp8mg+n
ja19DstuACeDQuBGkyPdpAQFzV6qSNJcMwnyjB8BxPHN5FFSMEHgS7CEfmsO
E3aE3mguMSMu+uhBalvuRmqYjSIK/gOSBt7o+ENyqYgNlcefSXB4ACeOIIfL
8Bgp/SnmjRL6MMtLZ4k3kC/XQBgOmd8+2VwySMQ/sK9Re0/pp6+TUxnbJs25
fmiN8NhKRIgAp06s4/dn5Kcz2Gok4vrhQnaEQ2hdNtuKz6LlGGtiNVMH/P0l
h688D5nRuh4J1aHF5YR6htGqx3VZBtTtfTn7DqsT/V/dtBpM4xsio/sl5P1x
Sn3q+Jg2+O/36Ez/2bzLiwWBbyKDcgtBKFD8+bVcUAvz9g5goPQYp9UyGh09
geW26AcunVLulC/u9l7T0vnKc2vMnTcirlys0KpSC3R9eFEDVb7AzAVg3JzL
z77QL8t1a7XEIpCipJ1LAwx7yPnPK6XZP4dbMYeMurMU11qI+YCEqKIZTyl7
VltaY0bre5wW0i/Ar2+ENNCI6e+lwG4FN26knOOA1cC3v6K2JeYTdhp2MLI3
jbgnhei/itvcyyAUEDNGOfPgHnVhRTl1K3x8aQpRge7e5iKHh2b29ycQFpAZ
vWzlQdSl9lzgvU3Xmy0/yu+qeOSC6GV0y18AbyKR0keGCgQCWueTSXkh/j/1
0fM9ezjJr3nRkgV0nyOxlzjj/vqjh51nRAHeMGKdzHZ2TwxVZvzCFJfYDK9f
iJAHN/qQKdDxlqz+IFoy5T3N1lPjjuRndWc8fp1TURSmf2g4dwRmXV55GoKP
cdqKU26CWntMebhNm81zodED5Nxe/Q5xjFnidASPcH7e9IwECKJB3lGQnKs5
/2une+c0X+KgsRFSXl2gV4/5qDV1oy70dq555wFu/kflGSRQhs+pcwOYnBLl
2np46vRKfDjHvx6XN7qnR64fNpfpBo1RYPW0oR/fjX2fcmeavO8fczUjpyRg
UdeCwmOYdoJgpw2RMpSkB8SfvSR81MvYvndj4W91r9ov08tfEesRR1FzOdGM
CLsmXFYVaDyDizHK89yfvzOYONQxjfnlz0e6qBBzSsyUwk0p727+bNtt6xD0
6ATe1YRbuYwdxj70RYGVtiagd0oCGtgFNaNc1TUcQZTSxjI0atHdViqMWiEv
6XfFSyB9XEZv4+ebkChocLck62jomp8BjaalroltXJJwwJXnD0twgLQyFJ+E
W1JpPW5hACPmT8GIidolXD3toaMmaowsXh07oAiPck0W1aInqw+cEnu6kUQ+
37XJTpmyF5csn7sP01ZIplSRbEi55SoKUGWM3rNlZfAAVJUW5Q1Ba2XPFOaI
BY2W6LgzTmsdebO+Bw2sZWtuNsAdltaiuXLzlZ/bFrLwkMtxMcVTT2mlcE4w
gt7cgS7ORAk54CBRcK+aEbxZsiFwapewG+MZ2Dju/woWyyGnOl/NvpiUp4hy
5HfhbPYWgJp7D/2NoT2prxZkc7QGYAbNFtD2Vl7TCtg7H0VGb8hgOIB4TG6h
yy2Qr5qZV4F+T0H2mGXMN0SYF9VKQTipOdHC+O59Se6+nBsOKdw5Nj/QfZSB
u+ZaUQGichGPX7xXus69WtkcOG15+/UusrH4YE3oDOXEOv30tK8+unHLnoOh
/k7Gb4eQdCaOwr/f1oFeS+nmnepr9ukrpYu2hJc7Ul86KbqO1rfAapp2yaaz
1ZpIcrmq2GMEulyby2JRkVzwG7WpgFA3LRAx/fw9Nhi1RQ3fDw6clyTsS2/6
rCVJex5sueT29Au6+FYkRDBBZzq7q70MXqfry2P8cugMntqrmUmvNtpUguTg
8DEShwm51jVht3fHiFjlDrV5iDL3a0PNKAc6X/okc7tC6TQbpBEfXDgxkpEf
cN0Fisemch8n3ZC8pUb9uT2T6iyVSlwE0PncXttptf9Wq58PdsUO2vfk5zFU
u1N1hmHQgv9yP2xb8xdULIn+yXJJX1oIR7IpA5McNbB6powMCOFGXpU3p+oW
PmP05ccQQ3nLnqLqdpozzfO67cufKH2FOo2/5uQHrtYRcpTed8JXXiv9O7eL
enRbckSNn+TyksJviWzswYbPG+sdwfpmX1WtKzCAznPx56JGuog94MCjrOz4
CbP9XC4feGQ77PmRgRzZ/IPNc7nd5rGVXPb3nEC1V4/Zn7uiV8KApe1xfJ6I
mYMNhED3/K9pxBtOQl4h+JzwyZw/tDWVaL4s73PGU/ewq8rtFVAjyczsiqk8
g2sM3+DOnPtG+WkOl1fr7qUGlFYFVlSJhvEeQhOxtn/05JQ+OPTi1I4GLc/y
bbQYxToYy6jRG89WcVUNWHFUKasFBdQ65Qjk4JDsZwMlszLAHfPjYu77dy+W
+wo2znT4RVsUgbD7siYODPojOqpAgM6aVW0GPc4rOeueSHTVv6s3bFulAMyE
jkLlNzFyvuCh6v2NEtFA0MBGhsLfjkUWe1NA6ug8MYov+bcWQ9nPJPANoMp9
bI3OscXA+6S//QQaBZQktLtTHgc6V7ES73qOttcgGha1LSgICqzQ3wBxucdX
51hG6dYw0Oj56JhuR6aB+GCsbgN+kVwFpUsae04cyydcU02B0SIqfPWAAc6z
yCVG6MnquOqgtPnaUnsuyp6KvUrwq4Jt6kV3aiqHecNgKEFiTq1w4woz6REj
DkSGHQY6fkeuGmSaF+muY74hA3IB5CyQDLOwAi52VxZFz3NwHnu31ijbNugA
5BvLf6ykaRrV6kkJBIHG/jDCk7QMZM/PhTz9nDhTL7QtX26lusLwmFz3rs87
em/iVNWzVWVooMoGa4gYjltlAtc7Gui9yNo+fUl2DkfqUatPzWZxOkAhK5hM
2EA52LUGH+gm22+LmsbhFiZvQB0RX6F/mNC8twcEI8/kRRG6iAyW3LRJrOp4
UcC7r3NwydqdSGEhtCUds1d1k+FmyTzOn5n6kX8DSbUqzfJbrehe5Bitd6rC
MSiJV/q60Gcn5l3F1E/CnrM4Plto5FD+ZDQ2DselciGM1BDLKC2aWincOD91
sO6hM1NSaVjF+lViSdi338k6ldtFtBjXbOLz9hHlnnNAi50nMFfFFZADO17w
X27bGdO8HQH0yI6YSLqsYqfDHD7a0OjegTA1tbuMEhi/OHnqu84QwpDUyn1e
aHCvHgfQlt89PPI4hHMhsPzx3tRT2J8dqbk2hwcXlOmmadHXc1m3o78soGsd
+7NBKCVQkOXfp9qoq8KRuItd+CwVjm15a6eQJBGJJ3E9OiKg2ddZfRF1o+gE
ATXdVG3+RMMR5StiqQMlIMhijQ1R5f2iMVm9RTbqp//kFeGeAbyJCGKZ1+uF
iWMG+I5Mo6R/tnZRYqNEkyJ8M4sfookk8VVVX4ecUfBqEb2QCbp0S0iGe72z
FStY3/mRasXQPERDr9zY6Y+KlzQUEWP8+Np6IHJ0kmPvEkGypD2m6Zoz4xUB
VBqNXdMsqUwZXzZma4znGBvWW42p6P3Xm5YS8x5acFoeMfSysbO1LeWKGHlC
wBxfD3/+IHZ7Zulq//xuwalN2jx04PdXrusHrywxkU6NBW/5HChsO5AHGrJP
1o/GoKUMdtuOuaSq2l1VlpB+5B3UlwwAh7O/VyegO20iIn1gPmpQMfd2h/qg
5apq+KnVYcz7qbgvk+G3VNobKay4oB/t3UtKXBHdns5jwxXiIg2m1a1816ia
8CWymYbGX9GzPXwFbycfg0Z7fW5WhSUs1CMkJRJMMENRMGm5aZL17XyGb/zW
9EDruX0+jUx5UTf8POgEZifoWtPn/YdVGImrCDLTxggTVPxGCIFB5Dq4b9WU
cT42g62b9qQvhSvpxY5ICTYQaNsqVlppTwztGg7ec6WP7PnLZiUdLGJJBD6i
sf21jAzrlhyutq/HgiDZkeJo+ZAfgzOKKyanunJZH5nZFbR6UMFRkH0gtQOQ
WWI1OkjGY75KdwjqppTg7UXOEJOXzP+WVWII7sazONR1qLlG5T2/FqEKc67/
UGFzkiTcePyl5yzZny5/uGxqeP/CVtI4YFrGStzdg4YmTuxdyO1CDxeK5RYa
6F5OSNKmiTUqbWiqPIwTDqsKG4QUumVk8ByATNOfcO/TuTOWOcZ7UI72At2h
zQodm0dbwvBOJ+3tjao5GHWbrGrTo0BtV9F5F5nqnldQyUGR+lFgsUbZIUBm
KhyT4hvgf5sZqZU9Hker28YOduTYb0ckbTZcuCFB8iBy3sTwqmisSvk40GLf
um0SWMsI6iDVycqqDxV8CbDxc1UMhJabDveSWhDZ3tgy462iztm1glKjmpZe
YVBJPrxlij4oucfkysauYXh6wgBkM2UykyoYGDRMu3+w1sgOSHZz7Ak9uz/P
Ann2+KbBMjEP9II60/6JVZLqBOqlBSkmhvhJw6WhLkWKPbbFuXKUN3RPZ9cJ
CpLy7QfRBNFYS36vwdT/njUfdW6dtfHLzrrsUXJeV8iiyP42CehjMD2aOSCN
g+dqdMggsYJCyAQraCxye1yAtovLqqFPfmGWmzvGxYvhbLdlQC7tT59Uk3sX
3DVXA6PuoWhB0FG5fcKKq8mr27hIJ0frs62XLbwgjLanHmLoX/HwgR6f3n+Q
+KUG6PGJrEs15V4tQjkwNS9FUXqvgWQ7F0WLyeV5mVuiv/v19uIUZUENmtmu
FHi3CTHwr1vFB4w92fHXxHLmv9fs9UyURhmvLRixxo6eU0/A91YkUwfWeoga
mKptBCUDi+TNE58pU4aUjOtDeW/S+heyNQ4AV5L+ADtwmeRb1YFIMmCQuE6v
RA46WvVjlv5iAbvQURRp93ZyZ9EXj7lnss4EJnC1nkfTUPhn4UWNC4F+x/kC
sbtfwUsVnpavuW0lbN5HLFCRDyObZyKHlTkET0pIAqcCHV1Eb5Gmv1VCPmjE
MFuzGbXz4UTF+ibisJC2Cx34bcq1DpW+ot8uIvsC3d/lgFR68bCsfXEegRch
BH7/fp0uVr7IL1JThZyluGMQgzFHuz4pBqVd/eg/YMpiT8IRvE4LDopevLF7
JY2xVwV6So0g0Yi7zJcGXG7QAbvP2V1s9NpY53iFEFpXccJ/YL4H/wQd6LU/
pcSwKlI3a2WV+exH8+xV0GN4zynmOzOBmlUaHQ3UdF8437yOF0UgTLFtwChF
slsLbhKeY786dR5chCS3u5k/wJ6Ibjg2XjvCzkddEYnxCAI25ugB7CT62VNR
s5nT9YkZ2SZxd9e+lm7I7yFk56j+mEMf433Qz47C1NEO+jqFyYWu3AuoG3pv
B07Y85Ey/iRabv0hqVtjvEVIEzqfhhhFUDI4UGHdKZGwYJ1bfz09JIlAqL7S
pVSmQMLneNPbJsyAtJmplr6MftDBvhVH1TZnKYI9VywXvoGWBvm53qXiKsXg
+Fh/J8zQAkurzldjiVGIM79xuPuv8E45b0uNE7tiksYv/O3WlPcuuDn3uJEc
d4bCa9B9Tde2WTzb75GjRvmfaKipGdHD0pgB2jxMGM9XOSbMrW0lvpv92CZO
aXlbLf4ADk75Zp4+E56YRUE9KglcFaChTcoJRXpj1cg3Wv1yPSWRFDu4g9UN
if/cRR7/AvZhhYYuOzjdnrKxwTqi2ewF2Vf1nvpzJ5Gn11kKWfy+KmrkCv5K
OpyTpYPP1XDh439RVu93M1TZqtAdIKm2y2SJ+iRxy8mofldB4yQvbLu1d78b
m3U8U1utHOH1CtRg1j8LUvTh6asEok2v06X6qIHAlW+S4mst/k9F+OgzHcch
sAfRB+CI5LOk7XqP2Up/9EHmML5JcGktrkccdboSgZ1CQKQmyCiz3pt/ArQX
uM2yguTAuM5Sheaywjn8xZ0I4idF6FCEKzftsQ9U52f3XA2U5JNc+JPmRK/l
t6CMBKl6/Y6L3++vfb1KWUGh/XlklNN0l2QRjg5hAauOc8AYhrzDxU+juP1D
r+3PDT5tWRHI/fq5mXc3EkpANA8KJu+AxAULC2C1AaQeq8XwqzfOTL326qt6
I7hh64WSdkUzNPH8nbnlQ79H99eA26gJEISEXil9GY7SDfMNMwpygDCmJpDq
xiZZ/MAArUgQ5+uEy5pTizjJQg0S+2ID091xzQcemhrpKZVS4bHmmSSBbCJO
tvr0KYRMPRm97o1+eBasBavEqGJrJHIoWGp7F11qvnxKjLUjNu5NkJsxlQwj
JCj5ZKu1gSI4dR33L2A4EGOsXuFsciFZwjoI1alfi7JCgVeG+pahzyebeBIS
fhUu9Fk06znzLWHBC93Dk4r5ECTZBrMl4/yT5PTrGM4EOzuEzrx7BYm5VqOE
LBnkGVQOK6/q312ZZnq1fWU6WYceYjQvnvGImXVgkTvpUHAEqk7h0nGHwu0c
jDsMbHtF5ULLX4iPd93IDfa6jCBN8kf7gNGWVCH8PlHOcd1TUeY9kaAsIAm7
6S2bEofE0wtie2FW1xIBhU+yq/6eCiukYKwlbDzc80V93/7xydYXxn0VNu9y
983ZRH9d3pu8QpZ27lSU20ZD4aR/WmaOJt5Ui6Dwbmicvv4HRertSyfJhKa0
C2qEDyiFb4pbMDhMYpYF/GtuPtOHyt6JamB2qznKLtej00pt7J8h2aAPLn6T
OxPTldlAOdkMkV35367w5NVpBCRflMaZwV71mgxKPvTPlLRUn/s7H0VWYSXb
05m/CR+QNtr5WKBmuvUjFW4QNAUpxT4r3wKXLlltfzLDO+XMnpG/DkrvCdWC
43yIjTj/3KvR9MoAVEELvPu6h/gh3NBfJleA14OZ4L0SrcLJy1MGe5LOrAFm
88Pstk5XPHTId4oR7wU6Debf8Ot+eG5iFQhH5nqT2HqFMfPCl9VefPVyzAVB
qVm15P5biLpcVNLCjkILc1A3wFtrDUH27oP9umjYidDmt61ZtY5XKSMk1rNS
x/PlH6TCmdM5xG8tVh3q3lmavW3XGbOwdktmHfYevrVHkIhWYDXOBsdT8Zy8
ZMNJPWpVSB2nGD/6mtazAUCjq55bVnW3+BUIvUQKL1GA+sM9VQcqXaupZtkV
NW8eeXpeaRJDr7L7uEy7XNZZhgKAOLbuRyP8nr0LPnpHFk+4UwH7cXoLy9gi
0Xx8LbzvGKJEGXSJa45ZrAEHDzP7W2EPkQaYF4VeVBSJ6GygonLCTUaoy7im
FUe9XmU9atbNyOX7i4cjS6QDHUQBoND577IKUxxQpM3OSyC+VdsK9VMhDy9t
9S2rzusmhs/wU/+b5n+HnyYuajOqjghrBJmVSxUfZGPG9+oQYHjhCDaiCpwl
fi5UnBP+GpNkgtHkO+QoTok7+eommS4Fn1CkO/rtSnjDJmbNSnjhtcNA0dr0
OF5mSACMWR+wIwXvj9XGhLk1gS5MCcI/akx2pKUEGUWXLN9mH0GbuD7MXXzb
zJ2IZEAa9wyC1uIrJu+mTOBbzDQ9L7hqOCt3AvqBWk8e0o95wZ8YD3qjOxpJ
ONV9G1J9ze+5WvUy/M5EfT1bUyciv5ngwSegGfRetJqyYCfhB5jQDEwGs8HG
nGhHfPR4b7JEABwHb9DkFm5Q2mQiu/71jeXciqTfkvgKIoANTH9xRnmFtpOI
Pq/wws2s3dwSmSKcA2fW79f0K9fZIXKleX7WdreOa/lZqIuQ8azlhuLYcoVZ
AXuiQw8jnEbPveu5o4Shk7FU6T5jyxFTXJhPUC/ltT/X7gv5kthHV/Jv4Yrw
LWQ6/YQo1qarlA5m115yNgmurZ92oDTCqVP27AYMxZoyeyrGh+/hJa8LA6Ly
bgcUAY+1eJnJT2JYjnYKjhtvKc4/loliE5zAFu+yjKZu9iolgKLpp2o+AV61
6D2P0MX0VUSs05PcAvN4uLWH9oNHKNbqg17g94cuq+sp21Unt88pCwQKBkKX
uxTw09EdztCfEJyOdyBPFLYSs/Xr17+CBbNeT9evwFAllxIC2/sUievWI7vl
iROeyfWVdrQUu64dcm3St7sXQt/iLETutHz25BG4zUr8+VpGAyGhU9rinJDg
I8wvm3zHya4Yd12E//mZ6zsALRgcDIqzAXspjbvIn/dIgz9/6DUqVNae/N7B
I7ppGIogFFR9ovBIQjOnFe3EGUuNa/LGW5ZozKfy4cLgWVenvhg6soqw+4pg
kdfrwaSV4wOCRY2AWdseHO+fSQMjmrdU+ApmXdOTU/Hp25TB538s6gKqJ1Sp
shyzhNks/NIhV5lRkd2LXzbiY1y4KOw7XfBwybexW30rJEd9Prpjed9TF2fx
BM/BVkvYLSZl2z1Kjdblzst/BgN/GLskxaFieqDegwI4quEQd/rIctzSU31+
tdgsoJSTbdFEfePOqLtfOZjqazm+X3H8Pjtqv3aulduIK4nEXHwVOqt+ri9b
NImHWcBQSVRYyicnLEngUeZ4/fFg2zBJVi3uHBPAsjdiaIlpoiQ1pmKFpSkG
G4aiqiI/AgKJXt+v5X0Xu9adfZ6ywphqnyFv5104+XWHzWVN9tSMG1Fc72zU
/BgSfPI0JLt5BEYhmaLE6G4F9RIg9UL0dSDJhJ2R+IQVQJXjNEB92eNd9zHS
OqX3sRqt33GW+d8TjHSbWQe+zNIqht37nBzQaXlb2GfemjfT/uATne7SkL1s
9n/7Jz6heZ8Dq/E5vH1R8ByqGlC8/n0FfrZmLMdKQ6+DjUB1joLEJH4ouxw/
92F/knUPqt7IisiFwzUJr8JOvd6KGfuXkEkat73ojUbAjIW9umVHLJ1nX2Nf
dAO9qcLDqg7nloUdG5vDfg+oxhe+LuHK8Ji2BfVndxVvbdmUdtV1n2ImBRzJ
aB+EG0l9Q3oysuuFnvW/DB4pH+xRbFLk6hRwrQZRgfOiJfkKqBbJQ02nD7+9
YhJsy2uc3j4ReK3aUG713UgjxtAOfhnXAndKTkvDeM9qzDAckbuRIxk4xw8B
SwsWpuCDHVhAUgNeXc3lNZ+mwjsqrgN3Ya7QjgmeZKfC+oPTTazrzRn5FOLt
GN6Pb+0/dlP+lwxAtlvvReBR1G/GDcQFk+f+p+CijmOaTA9qQnFm30atxAsg
9/Yc/trVsdjcDG9f2BEK0HksJ+x/SJTbAzCRPvd8wgdsVT5FqtkVVwwNqqZT
K32v+J8XFsoRPdp8BgrE1UFvjiKZSRfHwqektN+QFKPSmuKuY9bPPQJ76PaZ
rE+0sx+yQwdLUQT95vW43B7qrpuW1Qn0ljU2tuAAHeZxufEreEy9Uwa+dHNv
KJb9idJQ+3cZrPwcOmE748AGmASoUOjIO07X/p3u5SW0yHcu1OO5Df67Pxbr
KDxnd38z+2S+AMk46C8Z7qv/iyWCeHlUhC7gZ8NW3WgEXTEHAGYpreuNduZJ
BX88BRL8KCp+lwDQGR7ndvBSPgat731ausO4IWzM45SvGS1yJvNxPrZy5bN5
G6KJ3JsG7F/G0FPyLEEQbTDxP1Z1+fEyTYp6eK4XSuCyN6AYMe1LT2NwzyKO
wORdmUY1UFTRq8roeuyuqVb9mb+D499+4aQRlZYA9zv3sR0LXNXIWVqMwZlZ
z+n3+5mn7k7tE8e2YSLtUYTWVIubH3888cBuBkw00pIE99yVUNd6meLmU+HT
pB1gaF8Ia7E0E5uJ+TMayFoAHBDwCfZHSZWI9BOssHVh/Q22o5L5SLiFQ2IY
F2PSD5Y2BsgcTqGDilmY/sXlQuopIOj5raOfUGgYMFbotGu++hGHbgBv+RAp
PPuA4HA9VSqC3DUPIb8RfPC8pm1Cmv6WDhcoA62SARMsFKJNt995snoJwYDa
+OJlFJpjM34kowf55dKBdG68y6jdsGuSI+5nsh7D1fwse/4Zqan9WMQUtNcN
0X52JXo14BQTDMMBrI1Vp1xRoa4JjdARNdzlThv/RaG1DUSUdaggodp6+KXO
ebUndIe9APMqMhsIEOAXLdGCGZPpOnFWbImG0to3EY/AINMa1heL6DZmC2OW
d+PLC6WvUdNamlUuQMf23RIIAypqSNpcRUZY7DgVgQG0lyw5BR63bxNSuslB
FqAoIbSjopxmNE9WcQpe2u00QrXDwABJsiPjvrxyqvrhnWjQCpV6gZ16Ow7V
AFRSGHNwJDQu87CWTSPaFaB14ycZGISNL0EXDptZsp+3NjKnnlJmD2koUQ6O
lwJfsbHAfV0bag3843ZoMyu1LOb7jjwI9Lh9jOgNXYSt1vj1k/S3yHy0O+QC
Qp/vb4MAAb87Wy1laequOFwf9/ACzBO+YiX2/wF5wymlcdiXKq+yGWCsAAbD
w3TG13ldUgh/U67cTORlyw9AxGwUwZxjK8zmSb4M7AR7swiU/WU21FbN1IEl
3FpHBLGgJZMza7mUAADsgMK552DZ1UZn9Zm+ptwT1RSRg4mQC34tHGdfMxXO
Lx25e6XVqcLMECsAMYr6+rlJyTqAM/tg7zOUD6xnsRvjOHKhWN8pTbk8ilT/
a1gIvj8mSGP4FZ8AXwLFZKk4jTmoC2i02QvgTBClX63IrhyUnzcg3Ew4ojY6
1oSHKZOaAIpaPmxa7gyAthI5ucTvLSzoKqhUiiCCQpM8FiwPizYuX9qM7ZH4
Ag8en11nUlPc1URsIU/KihFexoENiwOI+qDaM2uCbtO15SZ6CLxj/BNfLxfM
9jeHU6cL1eQWtc7GqQUWFn5MjazlKgLGbF+CKC4uT0ClofR1ds4cebI03Hyp
ZBFqZ5MK31lnqmujp4hry9e0Fo6yrwkCo08Rh6jLEBqRR7K4YedM8KTql3+P
v3qiqtCTK8xpAYY7HUmJNofJwQNoXnxTk3twjUMtYBgKbB5HAa82kNfJ1794
8Xv9GQ5r1alUJKw2ufqLfGFpdD1LQbCW62ncAxj61PQfw9r3I/uVCRo27hDs
uXiBUebBLSvUJO5pljInEf37zDbY8how/QRTKQZb6qFNwFxGQuPu0jB/NjxN
0Q32CjM8m2EWlEl1v8dx2wuY8O7riPOdnZTyirG8I+wWYjKlYCsUYv5ce5pU
jF5B+QLTVC2rzSOXVTjpGCxApeBXMHJnem/EI8yZzUBJIYfiGkSwhTOoRtbJ
beA8kOpcE6ojlr2zwwpqrlteSH1jskR1bRhJac0mCCVIB//n9NSAUqqL0+0g
yI6k+yZiFY9Ch2HRj/xkyfn/Z7TufYP9xyJWbecikunTwVcVdJ76bZI7nmn5
2/sPG9xtZ0kpQ+ss3k22QvMvcAe6FltkgqwnmuBIgbHFylc1SY3+YdyhXPfP
WLpYwwvLO2VIaR04BZCcL4+wSWEk6JsS6U2jxod/9W+H3IEQkCCqYw2qykKx
UNHGJr+MkXu9EdwDoWc91uFVDMq5j5N+q1jkHBCowFo7/1xOzSHmwok+76FX
I8+cYHShVzB+M+adU5IUI/2ujeC0OdNwoIdSrfVVsLX9pyG4DO9B+ChP5X6i
9ySpKeAoOba+2apw585e6jfuwlnrsFzonSg65ueTQDDFkeu1QuHVHWEUnvXA
EpI2rhikb2wucfwB+tDxDX+oah6pHS1lE6aUihdEjcB9qcFR4v+9SHTYekgp
+18KTqSE+zOGQoTMirWFNqeixDl9HAfpHZqm6zYfLZ1piyYMaC9uFzTg1YnX
91Rp+FwCT1HRzn75vYpR02Cw+L73lfruYT5OPjxAJ72Eh7wqOF5jxaJH1DQG
pleXGvJYuWXwd46hc8ej7syXF7DzzU0i9IQbulhRG2B13wCb+hNiTHJD8m+H
eVBRiOiLAi4rvoigWif7iQ79HX98ocPN4C3L1/jCr3i/emaBdHufcX628vnn
7k3VMJ5wBPnT3B6OnQBZjrgCH4IgJBcsgAZLlrZYK6PNOXYgxHsO9mFvPrUv
PNKh+X1o0n0385r5fr9TRK6zCMpKgp558QAJJMu/z7Hucu60PKKZSrZKFnNw
dwb3p1sZdj6GVY0kZooynKKHm6CLwyjsoyQMFIbP+rSwmSYgoreOqlNm7Heu
16S9P5g8XDfwdH1/xKHEAmnjcqB86gOz8hLeD3fSBYdQEnm5RYiX5hzT96/o
keybuH87UYlTeS/YQi2N/5MoJE2GdmuZxsL05A4rCAD4gbui614cVVle66iw
UFzqCJVgpX5rGmz7/gJliUkyvnNin9igASqQhKV3PAaHzP2h6RCz0GX50pTl
v+KlT4ahcEAI5Wkof8BpYhLYvpUCNPQwp6p59PnBsS6KYBcZ6/Tbu3IH/aNr
YjVSjJsAPiooyfIbncmpOSmkaUfQg74xrpH4SXx1cXWysHzP8MPAJVgWxQkb
YgYxQUJwi005B8VA7A7OUzU9egTacMZ2PLl/HvQ0aNPOsBZLb50ghwaBDy8P
acXWjPfLXRCffV+89C4vm+lKYjlZEgPMHffb2h0MhO3oEzhn6QShMsb5Yfuq
iEz2/AyzGNGkXoqqA/ppylZLxK2HVco0CskVhmDTFyv1Ad2s7XL0eakflYVA
l5h6ygbAEk6+ioanWckem05LgoPf4iR9YjMnJQ5FjwGWsfIjENPQ+doBdHkn
BlvTMt5tEGzi6EV5wkA4MMeFYFU6OabvD2rXD7ljA+4v0r/i+MKAgi6df97Y
fVZrxWxsugXdT/5RQ5XKvVa6Sl5cL22zt/haR9VCeA+z5ZJ29HB1hCVDqcro
zoWhtjYa6lGnENkLOOuk3q4HW70dBPeJQlsP/SmUSzhCJzIQyHYxoGB6LLKu
jxZh9pAJOhR0s5+vnWOCZlDfV2KqpAKz4riolBZBYGcsS+dxmMWi6KWy7vAB
lwVacgCV8UHIvPGDSxsIy+eLJZvxafCfGv3UhZLbggs2m0GJQvNekM4z69tJ
JCSqw54xqKYrzemPh4sPHSzcs6K9coXgMmmxNn95RwgpsnSHG8iJxUnUVRxl
hzID8Ly7bAE2/uo26Mjib6nvLiq4oVEYBI6x/UC3uXlnJ4BarIEN3vTatoV+
DbGo9nD7uUVX8jBmirh0CiBp8HCdqAZDFIr2SFoB7Ka4RGD5OZEkAX5xEfVi
vZLEztUxahlPZGmi09c3nFrIIunslvQhnIU/D0swnLgT2WC7fnzl4zLrA5RP
/+TkHj4J+bMjIAcwc0tyuPYBOmiUpVYlBbqw+1UOb0o+rvcgN6MgoUrXyVDr
tcvOUsK4IYWaGfTKlGNYgq8+AsvBeaiIMqOUgCY30b80McYHS8/ZqtyB+fO0
8LXkAu+k/u0KBfyZPN3eROUD2N8jyS4C+yR5Yzvu+q/TUyWKGCTAjvFKkao3
8vqAlnEEYvYQjcXr1yjPn2vAtos9z6ByMyyFrmqYkuttioRd1fmUoReZ2ffL
oRLJY8ZqCV73+9oB600sGp7off4qnmuzyKOsxGQGu+m7Gl8tzbgAbSeBIPeQ
1hWxm3xixIutsKAiAJxJ+GhWV1k3hC9RpuK3y/rBhp3yUocK0tzDbQhKHfHB
RDft31DaBnflmUfrFLDRCiSYZll9yppA1CBoUNffTYjaEulHu8Zw4qmnU1Em
4xytNPejTaS1Azv2pzd9Bp321a2MqxNuiXQDUbM0mRVFkS8nd1DeI6cZVwh1
CuRvdLyvMuvKVLnb9RoTj75GcRQeEtPFb/YiWP0z4waBKR3TUWYBkIud4dlF
3WYKpwzO+kFruT2ZcUI6nEaicYrRuc6eFBj4jNNs1dOt1GQJDdsv7x/2oFyH
n1XujqChQ7ZTwRzWErktXX5L2Yx02WCdIiiVPUf4edbbYv6XWrJQvCDE04T3
aohwvzwzXYfSriDlmqkQ/r5cboq3BVPLjsF7DipAusy7VSfXeHM2Nc9BsoFD
zeUpPLbAeTlKPVi2Klw89Ndank9P8DMjOBjL0Fs+uJ/i6F73NutyoOlxpBvd
lCtUM4gIOiYVMaNxaEr3SFR9paRzSFZKg13bYLPtj0+f8m/9xreLyVlyrXbO
jrlOX1gMSuP1318reN/5P5z4Hbdd2/50OA7riJiLkYLKNAeZbSzAXoB2q0vm
ZOrJuee2qOgH7XtNDlKVXA2iprmMQnBjccm6o1Kx4ePFNtKftMpZwEd3a5Nc
x1JHfK2SmX8SLU8HZnwX/eIwi2Ppp9ctZ2BSA0XV3uV3U8HsAkoO8YQr4DZP
q/YYRmr0A1vswhoCoaIEkgDZEbv1gJOVF0vnTYEiFSMXmpNUMn4xbHJk5tzA
fDkM9gI0k+JO17dRUiDCcoZMWrbwYdcUbuujGSKWE69uZl5HxzBuB8JsOoeb
ZozZKNBdXZQVBSV/fB+55VomY2RQmBd/kHOsorfLYCPxs5D9c4X8A7L4oWYl
SvHOk05ehm1nANzyEme0YqkOx4wY+YqYMKSwnply7HfUIhRNIn5nGeH1rP4H
7Mgu2CMoi1PGBgSMcSUfEtBdfyYKXCQXFShHp/IVfaG25W1RLZl4iBUV1Z3z
160VICLKocCNHZ2l9nf2mwLs5vG1BmApEO0TO4LBAtqFaHmzkbOM6QAw5S2g
ysApX47cCJ23i/f0NKHkgUcWZymA2JXPVc5Yto4E1YoMy4h/bJIQD/NC2M4u
KMasxBQIQDXEiYnLQQYFDqETc0OrJ8kXvI5jBOkN+sKFr6a0OSMloIXwAOCj
/+llRqaPwD2Msh//fp2vSlPotL6PdTWOfFLOSmHAAtpjogE9RlnCK5EzwANp
ZjKxp3rPmpYOgzAl/6nEGiMou6RQgpNva0qn8XJkXl4hUpHK4iW0huYlI4TV
wqMzf3lUBR6GAR5rN43Q8C+BfMgyAaY4pFfYv9R8KzeAB8RoGIlLmkNItFwf
4nLd2YA2rvEK+3ktU6OJKHZXSlmDRuvWzDhC05cvDEqHf4Zim6zo7aj9HWAg
3uEDZ29CPIOFalFI3HM6wLFqpqpNbEaGYrWvzPrr+t0WxX9FlSfQfRQ/k8EE
rliQ7+BwaLaTYpVGdlXQ1hOgY0ATzwy0FZofAzU67QFkfFfQMVmyWEdNGFtv
O41gSMGJ/+TqVZO03bEYg3SWufgYAM6ycOF/GT6wauZcQxdt+TMd6GWzgosX
B6L/3zEppKVgh97FocT4wa6xbREvJjg9HS6OVJrgMg3cuLyASTSeYWhw/OUV
KZwTxGhMnkUd4IczmN580M2b+dE4/0eF3XfaLc0CsYfzaoIXc3fpJTnSB5cx
/V6gH+IGfvwEHv/F8BPaEs8rXbcvBUJ264Wv0b+tZ3Mnjfsk6M4bH+XvRmYG
suFkuavurULwO8GHpy3rJPDgiHB7y5O0vGwf5bO7wL7EyOIUsSlZYnetz9tP
gugFF2r4a3Yctz8Wi0aqWMpyB/yiSpHOJpZ85m1dJS79nzWIGgI6qX+klPEq
LtGgRIBXePvnbcrWq9AsmmxWiKdbydyWxhA8UlvdrB5hD/r6i7X1cQnOOLYS
BKets14FAicRoU37CXzd4i7zz5vjObq79tMVrV+n+l8U0nL8DYut0KMHks4+
+uxwYb6vNq2cULFiiLAkNC7FhTRPlk5Ot26dshoo8apfbJ7bE8P+rjN9QFZJ
/DztvXsBLg0vrruSnjqgLpMVcHjDatsptgNaDJ6r4lOikPcomsL50JySDbAB
Gi4IE//Yex11urU7Hp6i1+cl6Iikgdmytu/3Yq+ukG0mUxBUQPmwBvrJ8rzH
TsnAUPBaSZJUUFv36JArBjrRyvDXcWHWUrhw51eQvvNnILHeI7sJ7LpJLhWz
aMKCLQlpEVTzF8xsUIVxbfSa2VCWTSzuPcpozLl2U/XC0fFGPqYHiJ7qlAN6
bZVY1yBEcE4fNhbHpXXFT4LP3/sEcuMlKl5BPhQ2IoZSJG0+9jFH1NnzTy/B
jFlRJuhwRuyf3X6NtUTIttM1/esdhP3H9FjLykGL6/NQ47AEiGqYtAAK8xks
+It5MZ0bd2eL8oESeRIk0CVvz5ipUklc9ctPx1kkD08CX1KIi+3DH7MRZfh8
UomM2e5qQl9fmL8ZNQEVSqxzKJTogX1WcJnA4U3sbJiq8pZJTN4Q/o6g7nG7
6Rmh9DrrnP+xv5IpharoY1vSlf6hjtdzXbm6dmBFQJ5VT9uEdvZD7CFGudLD
42Cs35M4huZaT14A/vu9KRQAYqOU9cfJwv0dcMNrBH5ui9F2s9kvmViiGLsq
7Z6rI/2ItF40o36kLZz6qjr5fhDvNv4d29312r2GkCDq/qVtJayZj0597z5Y
a2tQa3B7N5qKhMQklqMda57Dqk9K6jqok0xBaVfx2lQT4gdELw1N+jQtNKUf
kop5X/tBuB4x/T6SmVEgmuKx0z08jxeix8K1+RQdbidHBmwblnTPxVlJ16r7
KJh6JapwsH4kXQDFXR39SecQ0fmIY0glWqNHj+bGRnTKs5bCzIptnEUIAZsq
fdFvuiaijVUnImwzqccgU4Ayaq4eGra1GZe6MnqlqkBfRozCLlAlCk+MTiA6
InRCE+NSlkv++OK+nE9e8RMFwwC3f7q/zL6/hyuynmwaukzeaqdG/E8MRS2j
UJpqL6r/oPLV6BwBJXN/E46dX/KLgAetJrtmoD1WUhv2e1mRxraEBvap0wLA
eyjFBddX/pe96i5vRdt2h2rU03XNA+QXI0hUSLubekx/vpOq6snONAMRjXu8
wmVTsshnUZMtYb4QN+8h1yZMnn+rABYIQdjP6ZTzO7DtpyRi0lV9OdOB+0q+
IFpoTtuQnCgCKH3RAGEP+7Ok+iPVb11wDQwv1KD4G2/YM10JNXTCFtIO+HPa
VmzDPUQV8+8ojq5iAHekq6LLD0KqHIK6TjMqq4NazJZjw8bt4FlhFDyhrWb7
H/bIweIDtXtQFDy2rSMslprxTXXLdq+9lqph1SkT7sAyDBpKg84Z66nuEyr1
PAnpH2KGl7T+IcbgyyOVp3qxDyGISHz02HpZV7g61594e4frKK6TkLcrrxQH
Cjh80C4QPhBetxJZsle9IYYrdB80tpPG1+dgVYfja3czgBj7jhMoxRxw+YmN
ehtjAje5zZvkKDfaYWaPH9Z10kfmeVkzj2ESfXiM9PnYlx/oNXDE4j0Uestq
a5MLQfL22xA4UDFET3xoT8Mt7IpMTxyHXXZwZbL2/esZD75jTaktHt/TPv60
ea2TwKaGoYTvmqFrzmtSSLtgwHPVJqMlTUkUe9jYdj7LYztonlMUW6yCN9j5
rryFqzxuLFRWSiIluZqLLYxq2chcULyQYqMqJHm95LszuHb7PWRfhzb8xlHG
y3qSWqFrvGbKTcTmg6iLaYJ/7c4vS/T8ImkQ8fDaNl+A9eeh5JLhF3jC9dYQ
Dt1YLuyJQAhKMg950Omxe04xEkx+MMqP3vlh0iY1F2BtYAYrrucHU0d9Jjl7
vjfIPjt8xbReR42mEYZAvqy/ceOW7THi7wdsRcY89+IUv36NVGi7aT4YVtZ4
E1+eKMeqU2qT+vfi28D398GQ2X7KzP7xAKyGUuSiKRGHvj5GHnBm/ZSFES8O
H6jhVR0a3k/kVOK7ldTzN/pnqrRZ3wpcAkB8M9T2evDi7vmshuYFUQFTUgUC
aBWs561i2vbd7emY8nIcfYWold9s1PbXgKU218x+jE7m2U5pIxhJMIy2XMM7
DWIay9mNbxZiF+UHaKmgbZW6CVaca10p7GPIgNO9eCmfuOMroP8026R5iq99
DQhZf3WuPg0rtANqhSuzokkFKp/IsWEMG/pFRMidsFVzfV6p8QhtQ5sRk2iF
AuUWyK9q3hCv9B47cI3b+XFIR8ndpf00lFm61gUvD15NqaVD8t3n8z+We2I9
I3kirlqU+Er4lxBsg8Y24aFBKmGinoupeb5+5fjaTGjPH+M5Kr8xVYR7Zw51
sEQJb9u/nsCFYET1wQ2rlcPC41P+73bZCNSmFQGmjYRMUFSXK6MtdnN7DxPY
gEqiYcgy8N83sYXmM3QwF6fO4h+KG/wCT6e7MexyNJtMM0j5MFrSGzFNGzAq
pmdebNQDby2bWmmIT1VeSjc3mRbWiC6smmj9Rk1iNekfiScA2HRH+QqULhnZ
O8NAK2djfooq7/4JiM0PTxxd7vCDNmciCvcl9QHX4mrS+9ns1Z5Qg7Xkx3/P
Pp5wyg+yl04og36crJwc6vGu6p7W8byC6KzDStrvotvlGbZHFGM6dCwtAynA
F1c99jG4gJR8+YFbGZwuJpHO/ADWdGJmmRnbQOtu0WFa6MCpxzr1nTe6Di3/
UfizkaN0GEeWhCfIIrAPhcrSZphmn8qybidO0FCZDLC7WRWdlxowHifXZg0/
NiSZFd+L90uSQRNacBF4oP4xn6X5pcdXmCIpRvGSGtVJKoG/nU0IPEAOAFPX
/TKhpSGX1/BlZsUbIPeXXQJy2k6NkFbm3JPTJlNSTrnqFlh8Q28ioW67ztmh
Olm/B74H/zSdUdBSsa7r3PgGgJ/KAwG/JQKVsUiCcCl5NPbEYBwI3LNo4tV2
vm8eX2l9/lyMgvZx7reZhgh+W8/X94fRIulFFwPyXWYCvI2cwgcm9nE7kwq+
IBlwC8tPOzZtPUTo09jtNY7mDMND0pp7vQXqp42BDBGUOBoAWS4uWo0SmjJX
TS4YL1x8CHdfGy9fxRoibuPOczIQni5faKqRHODh3Q0yetCWojuVLitgZBto
E4L4eIAmHWwvzE3J2oyhmIfR/apgJyKb47+15ELGJiobYKVMXrJO+o+V66Yn
KTk3M/vO/qFSRvdWcopXcjLyBRzWKtpmoCXonhU3udVBsORVY3rLFBQDCICT
6tsz+6jr5l74YAeBqUcp1v3fMlSt61exNfEoQdTZuIcgJ4PvJ4k8ckgmqYDd
udgyzdv/JVW+3D8NERoJhbTI69AQLbkXKEGc1K1GrCDc4lAL0k5isQcYSBEg
ig7TLvcOtsurPNCgzgJsQ0wmv8JPitQSdc0rLahuRpRQDo0dWZcxunt/l0Il
Dt2RNP2HWnPt9ZA6vfy4IvNL686viBpslMkHsR/pArymscxmRXllMhnsqo4C
bqm6qwPsZipGXhZElL1SMOGnCwYLzsaCr+4DMGm0yblIK9iveJ56rZsHa4NQ
cUtgSgMoy8OkmuclWITWGWBBJ9tTAdsnFy/NLVHmgersQaoKv/F3PaFlyyZO
GiXrz9vYzVvc9DbuqX0VKJtsZa+aHbTcPpC5vHD4kfhVBHF9pYEzh0Vtlv6y
1l6MrbIsdBL6U56H87CVcI8i+k6A69e8GN1SrWThlwtn5SYpU5MPU6mSIyvL
dum9E3o5OCgtChrpd+S0eG8Yyf9D4VHBw/G1Xlzd0CwdxOelAxQAuIkMxEEb
yom/dXsf6SUg8vFi+mSLQKO9rKx3txSCsQWb5DyvjKewqo5BnK7NhWInlwt9
BOAW/vQkvaEYGnDsNrxDKsQYSf8N2wapiAdgi/BRSO9TQDemS4gIMUkVJUNi
V/sDaCf3BlwQAkobzlv8WZo/Nt6SjBaJEQS5xx0q0t4f3dq7t3lo951r4QrD
yjBeAFt4H+z1f2tT4zU2eIUisrG5PZrIi5AqSIwhW9T5hWXwwmHch6tTNAA4
Et5XLlUCtIYKeScnJd4aoPdetcjlxamE9pera+QjHHVe21RrgMaCOlDUbkUm
pVllfDri/lJdEKV5LIT+oPccb3gxNs+1LLi3Tk86WUGS6/+t/ZocgWKpHwpe
QA4e/CV6T+wLXDTqWMOD/WjhJyQSpmWDAzh15w5Lomvz7TH609Bf8K/D9F2y
eVy5/hoIilgKNe2FqjAPF5cPSPt73Q13XY3z2FMtSGjiI6vxjfiCYbaxOQZN
xnK6L626MnFv9gen2VZhXmMiF3YFLGX0kmI/FpvRcv7PRBJiPBjfRQzxk5gf
p807mYrgi67v+xCM5utu1VMY2CucbPyifZqlAKkSXNsRQJxUmcbq1wdcBKE5
9DqJoH3BRearIKTYa59jZGhrEeWlMdiH7hkCNqIHkRiYOSv8wH/MCkM6MMaT
Gb+TVNiWn0DoGyLIS3+yJd/NeqgM7pqWREkzh0o03pF+B03fOkcsVfexB+az
AhJsUxtIw6ts3GmcWmfXT4mcwzIvUCj1CQI2nx5fSxOFq7MQN14cy83vod4j
tDaiDyRy2oRqdVflDpKKNpHEwewxfB8uxrUENvICbqXnItCJ0Ckcn09y9Vv/
6wRFOhOztHJywgjjLjlT/oCPGQMu4CmT4sWYg6tcJIxg6d76bSw8aLYv7LUr
swmszTmXfOgU3UgbwAFqLjpBpB4lvBAm1URBoufPO5MXjiRgI0P8fv+5gugz
HkHjA9ypG8QVmB4frWvAcwat4RN8Bmd/QCeWaxGmx+iI81vyQjt26H3ZiXTL
A4wzxRO+EDXB/gTjCoD9jJblyDNCKOkaOLKXOFq10+t4rTNHAIkpXpXmK5Ud
OeFAhnAox7vihTS3AZ/MhVMrRz5oqjZEZUXPpvFbfCnnouxKnupxOKtwe2YH
2A7Swi8nAS2hunKXjvD0M50WWHf5DeP+1be7VPP7wQxchroa3zJwGHS+utws
Neb0VoUKf4i/OL3fxhE9Ccd7AzsxhNE+HmOGxjx0EcoVx5L2MWr7HbfItkai
uPd3QPenFWKq4gbyB+voOhC4SYBdGgW/EThiZF18UxK9yoXIr+jRUPdiLsnt
mnvRs2oJhGhUaAfGZKT4GerUFmpFa+LcniDqQ6QXCxFYMMx/mWvPgi7ZOs5r
APsgWHNvsfFHGJZUzthdKcP0RJoXprxPV+Ju1KfT309aSjV4nUn0jrC8MNJZ
1PQMrHAvy9kWdHOeAQqrefI52DkHu0jY0ozYq6rwMqtivV94iJFwFvO2wkVZ
a4ZSuYc5u818um2pJg2x/TYDeHFIru4tJp7gnDntx2v5Ij0iMNA61f1ahK+E
fSNADsnAgH5D3IxY4iqPsCe+0h3mKLP2tOFbdpCij9nKaAz+FkEmzcmfBzqo
iYaW07SZoOENE4tq/cptwFrdmdZURLZKhH/yCpcY7yCXnqALhF7yCqrPP2/w
fJZY7gfNUNXDK9ld7258cpnJ7/3/26Hhsw5Tez8prvYJ2nt/XsXP6DGloqJD
NcBbbIiDM2WNSGZgquu0nnrwTSSs7x7oTgDjSROQPE9J/h9uPGC0y5D6TCVx
n++m+l1wGva7WHPbacK8FGPhujZWRahHkHwFW8oVPosW4fprxKIRVhL3PhAc
pNor1hG5H88i3Dy/zROm6nDyK394khFcWyAbsLKVe+zhKSK4NJPJo0uuhAgM
B7dbIN1QoJg3/mAxCtyTrC52DOw5GJsSZISAhWO/oFZQbVeDrBuvqK7wUn2h
MNBDQHDZ72HVkohiqYxF8lnQBxyQUNsQobM7RumFCP9rwBtEymyiM4WyyG7k
Fg+6PpHOTP9Dw0ejcJ3AftIRMKYiWPhpGqgjbjgeglo1OJEnMF+3cC9Inzy5
UVTd6WZoNpNdBMLqZJuoIGGc4B3qCEzbmRm18bGrSeMRXT1k/SBlMp44Kwyl
jnsScL9tY0odBnAP3nhwsz1uAn4O8f8WiGk+tEgyRES7WaHhSMcWlK5VTJ9g
ZI5GU2UxwZMr+uEihJYtGEKyRbgqx0kTU0ZchaX9BzQO3weilDWzvesSu+N4
SZTcwNtfAFUwVDbJoa8p9EaHaYIi9q1cCehmNufnS4Yyycol++phh6hCsln4
JLcFO96mAlCm5jnWo07nrEnCOlwAAHDXg+WP6aZA4jdonauNOUiEN+EvIeF+
zlDaN2vptnT9dupP4QvJiyaLXTUWwOfw6s8/ImU7CSz39VFo/gSS9KTO5wAz
QtcWt1uCaupfaqo1+O5+Y5EvbHB5CNoEC9jeIq0pGE8UK71rXD5sR2js0BsU
TroY8qnaQOK+SUfvhirPosCezaTuQ5QToCv9xE23eFtor9lVupMVoudwleTr
a+ezedRn2gUZB8go2OjMNVGXJ+Azmmm+I0YHf9S6tqPunlJtKSRas/q3Ymob
gT6mwOraoccpP40XY8AKqE1PLPT68bDZRby03ti57j4daHUQLPTgY3msW9j4
DzoreaTetfPMzr8cFUAz2ndFnE2njvC9ZJ8W87iYhVzia3w5s4MTQqcTws+6
LHU9DChR8xGbCvj11x+mBa7DGDoQjiAGKrJESYpnUsoQLL2EZpzCaEnsR5vE
ip8UjBMqkeuDbhb8srwUpI5Tf6F2Fg+OFpYvIvWU3m7Zspj7OAI0RpWro+oU
FzM1BAPIIXPTle5LPTj9SmhL0DZ2G+BkKbsDg2sK0Ll4aKd/U9Bih9c/iYwj
CeuXNOd3fLVNFksNo9VoUr/rRuMiik8Gt+y/vSJmGpPEvK7py2E7pOedaiCy
XgIMy92377WoWVhcxnhhNMZee21v880b2ZG5fUrAyYAhdSAS/0msnqqQtXAq
7Rl3RrtKNhhUJvppKWmMkGbwmM2bkTOtCP35o9vqwfI5XOcyB3LDrU0d4U31
waYlRihnQnL5l3nLT0YSBEG46huCSyIhIUy3GeNKoJda6GxT9JvpxijzZ8QP
3EIkJrNrWUhhXX841mGibV9RhQZtWnvyWSxXY+A8ijScWRSTNl0Y4xK53uXw
p3ibz2bQi5pD5fjSCY8c9dmLDeBW9bvq4PGDMeR41IqaFU5++obt1Q7K6hV0
1DZH7oNtjyQBuJGGd6oQM5/oQjmldk8vsPg/FRPoj93jfo/7gkckEtuyW/M7
R7aHL4P9DDWhF/pzibX5zldU5BP2bgca2GsdlBER2EB0f8WOn0sscOun59vt
bp3FecxvC1ttN0Kx0gWAaePYGdppa7S+KClXos3cHk0imjJMzIozkpr6q8nF
Rs6qrLEgR+YRp2iQ37rwbbMCRAepukgqLg2UOzP+KkypoNpM2oOjKKtqx6oL
CAzsTRoA+Wz50QUgGsi366/GquLT4WzCcAwJn/hjFEQJca/RZyIlsf88oGYZ
bkt0Pt6UATr4mnQmHQu1qj38IFgHXdSbTm0CK8r6A30Gy9xbQCjLuE91MAAX
sRvZZpmxzHeYlTUFzy7NFBbqlPbyVI4wPuloPF5JCzmbNkIgVRwM2If6RFDr
etEq6V52TLqC3AmwAQY127V2GqmwlB+IjgYjLdQat3Qpk72CAd/y7hawHg8g
n2NTMYgVaVRKEdl0jGkhSjM7T3Z3CDrWHLRm7zeS639Oej0gfkV6HZ650Zc6
YKWYSpa3HSvpZh/Qw59jd0UyJwdtRDJGYNdTA9nt8u9o+kyp+F+X31rDDtFO
wyPpclPeTV7CqZ8WHDQSkwDzngpIWBUB3cvwS4E4yq0oSiX9axnn7YiPSLgy
xJaEeO6/p7WiFxtT2L+f+iHO//RcX0sIkDiSUn6rFYjYBMbRiDB9TMBL0Suw
p9NXZOEoTU83J0M/7B4EA+ZyKjizKP892MsoCEjn+Vqjaw/TZsa5iWgExZHl
kujZqhzdlpPR8dtZfa3vDn8G5aMc7RP4Tn1k3vEY5cmZxWyc6NPc7JW3MtLS
IzIjSeuEYl/C8ugK2AZp86YsxA0RzCsQkZmdYFl43rvLtILe0mbHSL4lBKQZ
sy7aAQfeQnPRxgG16CyMgZneWVQP2Y0tSIZNxkojgC47nx6SF+nE7cKbX3E6
wGGLyKUe298p9hRsAMpc5QHRiSjj/+oP5Vvjq2yNsUwgVZF4o3/9jhTUXO6C
X5UIoFjCL81t0ieccbwLwjFOLru8XM96uYssbIw7+u16e3ZZlqUSOlpoo0DP
+5BSpWef7f2d9tROt+oUDEoTdy9R3lqie8DhSFs0Q80Y5JpwsI/TIXeVkrNf
cRiJrtxivKlDyfsh+rd72DZRRWUB0BNQkWSr2Pit7xPADfQhoIKmqjwjScIE
2+u5SRpKhTuu76/Yzz0CGCdD6kYA0Iu/J6NhGfR4IdIMlDuNraWpx4OMhhUK
/YBf7Q+KjZ05W1bl2fpxiL+wO+yMovjUGN5TvkvtuXV29ncPJVl2jmaUb/F+
fV+d6i1g6bW7+jb1wZlSRumvVU7knTXJsCIFTsPBDZUV7bBQSow7LsGHyCTT
GhRNpugF1xvVokoXtK0mAaQOXpTDUwjJfi9EvOO/KkQPqash5ZtNhh1ya+kj
f1Zp9+4ZFUbGwWZIdpPoc/o0IoaBvCeEMu89WC5aZUSCYxjkJLj0bZ26clGV
mWVcLRS2VF9fBa5YjbVWYrktTbJZ3hak/QIv9eLS3vu1494ipmrkDfLwUdnV
sil77lFEeMOPbTTXioJrNwEW3+UdWzrtUeEHSr2Q/udatuPB5eHtajX2Ysm0
OuDUboUHzHCBYFLkJfxuv9CgIEI6FegxlUDhIw4amhVmk/iRkpPANbb1VzMX
5S5U1LDhehojxmN7+j5EFkBzQ1FwNiRFCFVKaTBkuZTemIf0n7WWaQBSeBFw
PXZoIUyg7rhOrqcc5oHUlE/SHyVRS8ugsoVr1UktnnjONR+dFQcMbDKputgX
8xP/nwDTsgPAQ7HENbFwDTdJdnTaeJbCRlxBwg/jtFdJ5jbHDyHQ2ubUrQss
ZoQ7KQttnzn+feTecUFzsSYmPEPdzb82k9lI/e30pMbhP/6x2TEtabO2vB4y
+6ufuB3DJKXcFXGfqO3SBHb1vF/PKadjlQBzFlq27SnoAPxLEkvr8ck/ocfk
Sd/hRtHGiOiLkAOyNinn8OGb2T9uevsZNkENpqO9MCCn3BF/7w4+fHx69sSM
iIQay/Q4JePkyEDBEyWZ3KRCn2N6L9j0kkOMCXIS1lUpE8tuQad42A2IkW4v
Hl8H+4N4K1PCC8M/YrwztAP6f7YUiGnzewcndJxRLuo3VkTGiBiixu/Wa07v
ibmDm9UGke7tZqoKo2r4fMHXs7x7vdVCCScOmlX4PVy6NrJWykx0W07cwVsA
Vd89cSgqBk82uNSbiY2b3cnb7l82qQRDUJ1V9sws5uOy8S/cht+uQbhagUQv
HrtRtzuLWC1+aq3TlNj0cSMy3AeXldX4T0AycHWdeAO+moNaHKvM7KgsbGpU
ykAx6J4VLX2yBQsmBxWgMhw8ccoIFuuhLFlbhl7MfKHSGU2jqzBLLtT5uL11
6oWmtYHS7BaUPRaDRS5svRxU/kIbcKiXetf69u2EpKttp/9lS01cGe1btkwi
9HTCSZQdpkisorTG30ImGL2LHq6by921fXCptDossgd+ARMz4aH31q+E6J+S
Z0sLCM2rcLOWnWwOpoyNsLT8KlDtsZVIArMlK9NtcGTQ5LqzbMyBbg6MlzxJ
xYP5GFKI8KdsJqkvddz435kKQLQ2d0QK2IzZ04thESIQoCH6tMFjfuvgWXV7
3fb5jH7f6qfQ/7SH0HYETPxNVvW84WqdBZyEs1CXRvvL5JeUoWqBDTjAGtip
6r5Wx087nQgEmFVlLdz81L86bNYHn8ZAkTbxgpGf4YtrdTNHfYwVjmHrG0D8
/v7a1B+4fRZC+3C6JdeLS1amLLYo420RAoOIW/w3x8jcZJ+iM/aI8czmY/QB
BPg63pspIbXa4nWCINQLOo9OdXuZlsfUSRW/r2Vp5lq2gkGvAMBYDn9y3uDt
oLRnF7kgX5Y56wf8Eq+/UVtdOTKK1ZoPNG7MXspOTEBeIWHHOsrmFWHgNJux
t2upu7Y0eIUKYc9zan87lKrB/hc/oGTUtcWmeD1dJhcdhalzBiUQ6Kmw9Rvn
KU6sdMePvdu5S8EGNON7ztXXLKVwl0vaRPejy8qASiC89VL12mw03HLxuXob
4NTUoc/2TgZhtyLotgFZBATySfpMOCyvapwfGaieliX1L+N9xyt0Zp9qqB5v
T4UGp74GausC+NLstz6Gli1NZE91DIGAvwhiuztTYif6in98Ks4E1NXF9bMe
eubgcBidLEgigkN7KdX56FkGrUIJkfjyudKND8GQE0ioxijU3GEF3PRCXr8g
b3fF7NwPYPYzMksTNk4AG9Pm7M/4trM8rZX8JlOypOJvCyBojXA029Qa3SlH
a6c6McDBhnWcYwRyMDDaGR3KyZtNACPEagD4GF6ZakDELTWesr6F3bISGjOV
8fosQafXpxhg3sgNKQq40lznafEwKGgfRytcYcbeOf2cPZ5SouYzNXqISto0
L8+niMP5EoJRkC/iXuTI1/Kqgr573BoefYeakVpUOBMI7Q93J+zc9/NgWLYn
wAHgwOC/jsV0N+AuwKRg8zQhch1fy5dhypf+RqEsNz7kqmqg4gTjBKlEu7qq
2hn+mdTvPAsOT5nPj8PqoYAuScksjWfj0ouk5NJaej3aWXRTz6kHy3FWM5Ja
ksv/i2rqVB/EPQpvnBlG/a66PKDwQ2NCQYUEhJFoC5uur4Cid+oWwugxcQsL
wEritiTP8tgREoopecsNrfoZbXQ7IzS+2k5RkCuahcD6VYgygDoiJDjStgP+
QXkQMzn0lCqc5cc8Na4yZJwGQQXQoplzHErdb99KMbi5pJlNvYyaFOeGd4n3
2R2hDhOs45behMUghI1A3UmQqo78zw4PF5UUIcWWsU5TD5CRsjMz5RXw0FwA
WfxWai4RTdnoD705T2hd3O58S7zxnu4Pr5gocDk8yymJhzJOMiF6cVMm+KB6
tJiLtwrYPgI98+P9S6O5GcMDW1/HYreI1FIZOXTJw3sWDN9k+9u/lQj25PI/
bTHgq2qe8rHoHRKAIUCt2+I9wBro8jSs7Wfqs+BSDAFXMQABol7n+bUHEPZ/
SJpOTgcMUl9yOc4qgpxoVm9BWrIQc1COuje/ys7M+m0hQyWiC80GqwC5v1JX
BabFOP740b+Sq9SC0nrmjmCiRRoswszW9paBxNv816RL8U6nbiBhrdBfGfNx
AijnoqehykLk0Q92pNAQFVVX+ymlNXao867utAs2D5+ZSnTCXPoLIpEYm/Pr
yA9beMf7u3esmUmUBuqFRX7Zaol6xSkUnKwtELU40BvqKOXYt4j5nx7N8+un
GQyDggvDzcsFrmO3WqVH57bu3MbcdH2DZZeoKh27CevgeqkWi52bw8NYJgMU
E35CsGx9uCxXDlibc5vTlGLLEy6ZcYuW7Ir7biHJ4Qz8k7ZBjZqwafzivNsb
GVuF85gWsBBA1YyLblBi1Y75kmXOUZttD/wdrDBY2BQcieb8s8ZQIVVD52WF
sLKUM3lrbjif8GwU6NKX899+D0BS5Fc9+Z/yP+c1fPsmxeXSG16H5OpgMy1G
hoV4DXiI8oPJPxi6CZKwwAJ/gqXsFcX+NL1bq0RJSs3EAmx+T/GicUPzN/hM
AgirLe+QX+F+gTQUc0+8A0MkObALF8FQtVe1uRhf0O/raoJaEoZbztryjIYw
iGNW/8UzHubDZa4Pzp4OSarHk+hqwFyXXZNPXuIP4RlQ7dTFTCtTqbYPLxDq
wiZy73JbV3rY6IvpmuelY1VkrOR0qbyvNl8DFX4erwCZSrQsVBle+/73RnJC
YpasVyyFnT+pJccpmBSjH2kNdBfnXm6eTCZrqLv7vG//hqtig6hYcc2SEyKy
aD4usI7Sdg0RVEwhZLy0Rrgfcm+ziUlLxVq83mxEl31+4U+l9YTtsgN4bCbL
/IEdb9njvx+5CyCsKD4z72LG8unAaRYM1EN6NMUm05z0/ZVh6d/FdhZnfJ1X
E44eV6BRWPOgxKDGKif5l8pQ91d/q/67gerI7ANs8TBzPRHYSfirJw4Vz+tT
G9YsCp5sVZhdVQsvbcZdwWR6NkNiq/Mz+InocGo0iWw5ilmOoD2Dq5YeQk2O
LByr9W94KI7dMDJxhQi6mS/HthoI1vBwku1S7q++ChWdhB25Rlc0ar9i0U3L
8ssZV9xF7zC8wx6W5EhfsGnCLQ8tTkkc93MY92Bic7BQJsJbuOQcr5pKkQHG
bTdyfY8FHh9d6TMfXk2JK/HXu7ckx5Ij+xx9mbHZ6wQCFmu/3su6XGzGqs3F
J68E81M7bTXN1lHgij906vRW+v9bOnFiohrWncmjXfDfJ/mN7VVq70BCnbDH
r25L7S+eO0oKX9lwg0ZrX+n+VtL9lacZjmnBFKlG1vkUVbTi32B0QFLOFcSO
32MyY2WVsgikDas8DgaRArPKWv4UF9D+a/nPnpaceuI7lqTOvi9KUnOHSBVk
OJNP+LVGTsKeBOHexJEOKA9iowilHZfvF3Td3/U++O+4nNmKEG5vAO6qw/Bn
8/ArZEKRQMT2H1JvAazgKs2/ZFPwhTbBcMRxYn9ODUpabFSnj5MCafprBVeL
w3/cmMqFg+UIstbh/3HyLzYKMbnDUA/3kdza/jJTFmqkJGVec19XrMM9zaCC
EpVSazR/ByUTxyonrVgU6ioHCOSdb5KBDRjOCF7q4GMyuqo5iPJNmHs5R+WB
TFKnhoEfwGH6c5SpLsaKGep4jpeWtH+2Fv3EiO+ZbfQ63Be5Whrv2Ufw0484
da45xVVLVdPX66+fAJUz7wg1q9Ynv3IIlW6YzoSk8s5ww56lLiXkte10Nhjp
PZiPACTz9B6Tsu6NJimEtS47myeDWWn4rXdtQywKukcXAIffZfB9PiY0GvWU
fbteGEQ7FP25lNVA0Ws8/SkSCKJw121Yf457EpXBAXP0HHIe2fK7HyrOetLx
b5VI6iCkOSFuFjo3YyVsfQqoTFGmM3qJ+FqVr0gL6uBAYZeTplv29+WlgNOx
5EduE32Dv27xSkHjYHbUrBz35qPrrlmlR4gpMrxxFTEWQ+byN/Z+DP26ZUFF
On8frs0rErv4yrl8xXH+CoTbk9vYCwzge8t6TlDRKcSM36wiUCiHqefRrUsM
YmXSPcLlDm7hYnNlZ5h9hHLbO/NUotYOVnMtvRAZCcA/wvTygC9sYDDaOXTg
yb7+hLUhOvVFMDjC3CVv0Hjpl62SWXYCHwVAS6ohbV6vDCzPY2peJ3UEpOxw
lXBYnVeBF9Dzbi6d1j04f5CKHbH32m1xNYPrJ1o5Zmv/5NU4VTN6Or73h2CF
IDQMlVpm5DCQbq6ql4wlnsE1rDQP/lJjPUgcN1l0Hd8uGoMYb4spViIbB8I3
J1Mlh3mzpiV8a4WuVYke8SLsT7JbtIbgUH5HNf+P19QIpxTkdmfjffP7Rd3N
856R0ZNU/678ulmOpBtltYo1VLFOvv7o1sOW89ATUzfJoyawXsg4hHc2rfT7
skNqYYhcKyPZ9SQ9YPNDZJu6RCYR5sV6ZeB7vnWb8XK9nnIsqWNPdKKEtmxt
YRoOeEH+cBDpLNxtKTdXGeBrd47zEJLsCX1emzBDrrKMt5JL7ZtVCXbnN1P1
OW0oHoag+UU4El5eMwmhip4iGcjMml8rUk9xhsh4mc823KnHJhsRxawe/Tbh
6q+n3RfH12F4Ou1GfvzRp8+VV5bfKy29jlZwuyT13dU9GpkMUs/NXZrwGYRs
jKeomj/Xq2UdZ6j2tuaF9bBw7py+YRVAfB2aDRVSc+BDZKWF1EanxWmlkRZM
U333UJKZ77wW4u4f025aSGtjRh5hm6qqzW6eXfooQJ9SNyfrT0s05cYYpn9t
q3m7rFSH7N8cpRfkUPqDbk0AX/5XLL9xXwHlMuQr0jdmSa5drcV4snmxiGqf
3dMlG9vKkb9XA1euUqp1X9LEYVQdtYwPeP9GL8vp8V97XzBD/4LesH5x/t6T
1W2MGH0fsfCiccqpVJdZIDRLbvDrn+Tg5+3pMo1Kq1o7xqKDhE2WbL/30UFj
rbzQgZnveoTnrsj332XKlM6odj6w6p8vCX8dsOcUoCIiQ58jnltTCkCMXnRW
75Jyi2nRMhSBL7nC4cv3zg6QFoHi4dfdgFKpDz/jEgG0LpJEL9yFBYLxE5tD
Di1ffdTmlgC9BUV+1wczrMQxhlhscYOV2n6LPgwUQOvVl9sCULJfYVb6wQpI
9V7+40b6ROtz//XBalNPRpeIkBOF/cw9c/aGlD0FIDioHhfKkU5ESZPuc4FL
mDAcblNjJRCEUOfyTHucAJmpGazgq6BvA2H3c8Hr8V47zI8gqZSSx5cZQkIX
69F0C13UerVq5yva2vgjTnz8hnIKHeK6Ka48QOwQ2RhkoMlIN+q2wJM3clOP
j+RCmnWL1ll4K+I9Kypp+IUynrmhmBDe3bFhTDmUuBpJY6kXBaXz+PoAZNbx
hhnPw54UGzR07+EbfDLvDPzWDSMAxL+pUS+Ly88xO+RnhjXVy/DXW1pZGr/k
Q1OKIAz+73+/o4o6+eBBBcmTmRyUHpyBbEVlQWjK7BHZpKKeVGfCUqsCkAvR
HDNw8WgUseY4YL2b2hVTNnrihGNPh2J8k0l3m5eWe21PD9ICMlG4i5dWZbtM
U7f1AcDeGT4CHpLgrB+Fz2kzS6eSDLGNlRJFSK256+CC3K6nNcFk5NgHusTY
GI7E+NlnWLPyZKgrJJWgH9N2sflCLRlUp2SdBBXK+c7EzZNBq7UXAQdTFdYH
jxklmSR4HzuVpjyYUghy0tG5NrmxcEOGZ0Z6ETZyT045nJPngI7mtuuhOmYq
cU9nRVlCm6K6EzUErcfwC30WSb+YLAzwuGghV7yKgg26AdKK9fThAXfMD8wp
dy7Xgaqzf79p5Tqwe8DME9xtnZNv2Bd9Zh1etbzvUlC6t7M5tBa8ccYp+Nix
r5zhipqZvCpwyjmBznLPNrA2G1EIYcgtl7OSM8EMpVv43wplznbFmLmll3AH
f8mAND1/SkaRM8iBQJ4qwIZjBPG0mYe/+nXE57eNGbYuFNLZ+bJ6D4/qBuUh
42AuZaB0aKCJOp/UO1j0GP8eEarIvK+QyjqR+W4LGFW3MCre6BiD5hkanaav
EZqlyikOn/ZwuYkLE+Rf1G1usuZminX8+w/mxVUt3F2scwHbx8upSeZwbJzA
1f3ha+LlD3a0Ug1mvZo7hu3kBa+liHMgOgxq4FcFwh7X7sxT+QU+ZbN/rNvO
oLh1O+aq7kjSnxP/Y/xXPZNjrQf07EvCyDXTMXBS9VqnbNLNEXRYIefLrk52
Mi7h4+LgNmYnGosKgcM67+MEkdE54YB98XC5JQ8ok3ZSif0rRYI85ROK/uiW
MMnYxPXpanpXhtrrpUyr+44gv6fGKqyjy99sAPEgGxD4ilpIANHitkLDpMhe
tT8JBYT+EQtgQxQF75KN/1oYzGQoCR2kbCr9FSxYdY1nZA9jYAnCkMS+CXHc
xCrj+ks69bJZe3UTYiXXvdbt0O4JWQ5zoeWWIIdVGqiFpduVEgRk7j04adqY
t2dhMToHGkkHNu89RsfahEXaAEjSUFgehBaCFjfFaVRIkN3kLuEAS3Mf/XG7
OKitmWw9WOxJe51B66SIU7uBQtAsTaAk6dlvK2NJclUbRpEyByK0SwJMSLNO
OiJ7fXI8pX3UEx/xkZZ6LKZoBhnXHHON6Mbf7fLAIHCZ4gsTu44exYSZAX74
B+PO1Budygs5ju31JFdMhjubgJF/a0qoKVLhGtZBNN55E4KJIdnh5lgT4hDU
fjf0bln3lpvgxRQlVdSRI6vRmNignoaUNbAri5uicjalH76/kOg5DFPTXDeR
FF4bkIRYPc7ma7AyXsgeap/jalhRnroORZCZOZ0y5aFtUYXgKEDIpZyOebfC
J2J43NFtHSovmjWJdtAVhPwe5gOtIozFe1qJ3ykzhR3Bj9gq9f4uvEykHZUq
50oqI6LQ3j872gvxcv4VemkUg1X0RDqO0cX7xnh0fIXMLLAYpbCAI/lv2KLh
JwNZITSK30o27Q2PCwt7QwOoUrNysEmS9Cht8DSxscksE6pgN5BDgbuJ/Ufz
pgxlb/K2SXdcKD9yaThTAP2Fjes9sbmDsXeA+bqqvL74Oh9XfAS6TT0YzTkl
WtuWTWJoLi/R+Z4IW2kF89lYr/FRWqmx63SxpQt1Ht8RZnx6R9DwReqy3jlQ
z1ygToRcH3DaaeKV6EV0HWwJuXiitBpQS6BaZq7QztYe7w0+ML2ujnyzbqV6
7p0Troe1wQS55A0Zd2hSi5uyTVMSfPawtzq1mehbKmfWBrcj2FPm7bOnwMpx
sU9AQwTk39FmFnmtFs88B0FLIVOpEd9EVIONWN4zANZ1K2r/g+LxCinu2vK2
HQjrx/ju8kKNxX0BLQJZw8QMqoT2CvoJzswBYsQ3lqmgjPHxM43+R7MYd5Tn
GtZTEUBUyForOAESbDoagiAMDfIoy9uPId/B6EDcMLSbUiakXK04sJDAQkHZ
6DZiSMsaSfEcquaUt2dxJMqDPwD0vPKWuN0pNrWSKqsBkJVEDuTxwi2QVAHM
+Ci+kQzDjneVGFyLMfGcEqBedj/czn6uQ88ErMJ4eDHerS733JplvLxySxQL
sbXUnSQ54YyWWuNcvNziid6Ykf8RGCEfXJVD9trVJ+QolY6tm1/M4FrF7KQ/
o0828zGNMqzhMc9SKZ6N3D8U6+XA2U+3L0dfFh+1lPFDT0yT/+7B+7A1s6NY
jd+M/slSI8WtsgRSYfkjX6ssZOzI4dtRmZ/b4wvwwyKIcrVgmCCDduEmShel
Ipi9GIEUuUUmiheiw6lQHf6c/p3qlr7OHMIAsWUCsa6eLH+ab/ZFJvADRY/q
OkIsvRdvA2udPiVsrnpueOspXy3PYVVA4R2UbuEvLNxjuuz/53Ku/QbB2Oum
qn+JS4I1mM3MP2CMnIYjcjXijGZ2MMJHeLE8dqZtwFwe+n6MUdP2waNT1LkI
sDBgopLVNAO45JaXGygYISQqgzlIUiOxQMMxTDKELYdi4x0jDtvlmGfTBalR
CubEdMky3AlvSlCpIoYuFiKzdAQA44aEw6PIDFjXvg/cJ7l40Nm56Eb8sZXF
jaEwS/h05fA/Ym9ZJtwjU5ObOHwRxE5yREEnT+Rm8HsIAEHNNYhcTl6wTdJ7
fTecjiiQk3jlv5T2/q57CgC9pPMI3reBG4QZ6wwQB8hJ/qcfwIYS7kMgiXDl
jBJXmPzYmMEyhW1EABdXgjJmLPqvV+dzmBJ/oahznfhRk6w/+qUcm0fpjBPu
zotMCTbZs45xRf0QcE1kepqhr25sxrzaWFpqdbW2Ykg6mbNTVN1nH/zq8Dha
CPwUd3w2WG0+S6C3HWyikO/fRadpzsY4OMihSOb4ee8hmJgQMb0ruPf4/sn+
2r08RvYHoee3Qszy8yOtW7kFIYWxN1TyfO7/J2W6BACnPRhVioH2sWcfEo7v
q8SfzoRKtYIEKRCR7c5a1mohH8GLaRBVB+eRQgOKU09n5A98WQS3880kvBpo
Sq0UyWzC1h4IJcEqDMa0IQLL0K8907Qz3+ddQYuKIIs7GU9uWk75YQ7irF9f
Q89DYyMaNqcnSTK1OPXY0EPf9ekFzoUKXmzpKKhlTBJirWQTg+kvjQ3HRVU9
rRHGema47/rE9550/9LhjOWpCBTi3HXfp22br8uelN2RzlnDWm3eHA46b9K1
jJYl/Dtj+H7eTTYdXXMK3UhizKVHvoOmcvSc0FtMf1LFbZ/8Xbu878eSnogQ
m7ofePCbvFUAWOqE7T7tyacSAWL2ZuhDjWaFqzVOriGG/QChW3izI0FKRVYO
ae0ozKX6bneZrYpZfIbTQISvOWmXe0aGWTaQMEad72RqkWrhF53kQPrcaAD8
O+KMGvj3iYdcYPBSGEj5rkvLbFxbH2cmEhkbb8bAdhWAzH8geE9m65XuChtk
Ba4DvMItHxcIjex2txKYtEo+8dRCd4PjLRbj7Tpt8AbsOYxE0g7+vFvuixRR
B9YgNw2vtAJr4NRx+PQiOEcMcIwDLNavi7N85xUOtydA8rFTF411eOUXp5ju
18OS+8f3EnKkbfZQBqo6dYNEKfE+HA/L7yeBTbO4VBEdBN9xOFqRdJfIyZYt
zznWii/2+J81FUr3YXo7rDmrH7nyH7zYIkU/q286U44BCsolnObW628LMNnn
kOM7g7dpM6BfQdL6glyBzHwlqV7Kkbwg3Jaue+d5ZteqTqV9WXCuKu8H+5r/
ac6a+4uVgT/e39Nz7WZG1OEBiEWz827GjD6FnQ4Jaq0ebWmqC3kKjzeiQm//
Cr/pJRAEzbd8iKtCHKYYm/K8mgKJ6DjwCTl9dPruG8hLZ01pfBAXLhqg1T/Q
E0JOgiFyK1pyJDK4LfRvnLStTL6zhnLF2Um8W/wxmkKYWuG7a/GCMAMqIv7k
fUF48bCj1grkrZQExUUaenGRedyLuanssO4IDNQjWY1i/oJ55rFuk8m5z0+b
gMDf7T/IA9v+O6NjpSCKkIS/yTFJCWhHI79cCB6WIjZ5FMOtwXv+ljmyf7ka
1cMcjDSFJ1x2RzyFVXcPUC4zIdsxdLpYuaNRgXXpPxDAkfbKTsyr0qUc3qYV
b9T6H4QZuH32VeH62+BsJpjA8Sc7EdQRVMfS3iLm5y3PJsWMicsFxo6NlcN/
XheVeOfN1ozwoV2RcUnJpjtfH8Kkq+pfTXuWsAVkuF8qx7DWcCbymgwkOm6F
exBQS4fBXNAM20sedjVIC5xnfVlUKzUets7dBlgUKJYPrFTzpS59I/3MTMw5
zErs9CMjGzEJRQrmxsfEJekmx9jMAVQ6x3F05/2If1Pc7Whlem3P2RhCYGgj
/IfgBWJV+kZIWoNBWugJYkeXcJeE2BpVa+Y8W73kfB89p8YvGYoh/hv1TdLg
++9xm6RtsjAbcrAb93TEnDbD554052rAjHPDYoCoXElukIMzprOyFwnnDTP4
M6gAjZuKjilzY2xnxODYynoj9pkdb6m7kGfT38P522AWyrJYCKKNGtwf2pT0
OJF4IQWWhfNktGPkJK8vcc/R4X+9d+yUvQHklwBctJc/MfUGW+s2h8sibSzi
LU8s2zaKNIOlqCLbfxowGAEqFOaHrt2/krLHbTfjZ9+5kRqgW4NgQstIORQU
+r6XpdCPoRe8FJVVmNjARXabcw01w7lLsBr1gyQ04Vr3ADbIeJMIYp5ScMmt
MYodDwjhwAcBl6lm8+xafW7wRyJDjqG2hkvXIxNiLd6ER7Nbsne3juMe8IL8
qibRlS9WEEeZbH1BH2NatXR3+McGrTYQjYh9IrmMWzrkrx615TNQePeP5xuo
VpaDHBCKIQv5i6Vo6n3KpRWjyLEqC/ZEyDrKk9PkYnnohPDgEG+01N/iXYrQ
un6mLAV/t8QSlP1+G51DyhRZK5O4o/FMmpKK0I9Xysg0/OBeJ52VXJoyyiss
lRjX4WnlbLzMlwmh0tiflH0rtvceNlrrvZkfT2WKacmBVsMYzh6S+lS/L3B/
TQtK+zIuTqzuGXHMTY7R+VfbtnB+ZZtMwdlLiPHfm4hjAOJSuKbUHKecD1iR
voZU2TZZoENdVBkVlFN5hCvMsZqS5HmQ1rbjwGGYgjbJnxfiqcelBkFrji9m
L+cD54Ll+FPsHZ6oUF2P6Iu7WdedRUSH9dEePWFehvajAut2brzShcSRveRf
OVyZ58Q2Rllp+oKleG+VryMWB1fAL7zNAu5TOvLeZrMWwEKhBT/1c2UN2+cS
R4GgIxpxDJuNgxcMvP3kuSura4seKDDhvC6ZH0BXayI5kpniP+PIP+708OuC
BG/Fdy1Sr5Bp9Z/CCUsIVgTamqxee0Sw45RXV653j6DIVrhIx+jEjwEliiR7
GDhuUfOZZ4PTaED9I97LZynRR+/D41VLf8oq33rP7GT0SlVNDxRyId2fL9V4
uBSjuQB+UcPyD7SmoDwg0b2Big7ttn6EVtFVv6IeOk75rMDo4qb4c2IQnv3M
Af4RoVXTGLs8d5wr+YDhxsR3hOodW0ipQ1BVSLWtZpjIJqCEnmUdJTgtMhPL
t8ldONFlxIesxixMkgTe3AfC9KiVNoPnDQroDQAXX6tuF/hQd5DNuRChSdS5
cRGdPMDRwPZxNifxeXc9607AQROOFkp0Vzwqg6o+uCtoOd4tH6uIuReF7nmD
t2DzNdAuxXhwWaT8UsdMiRUTYjdbtw/36NGy6ncgnFqk4ZWMM9s6EFmypMAo
CK3hiUgCXFU8s2jF95IxRoDb3gVtz94VRX/7v33fa6jJ3Roe95xv5FPX+Rfd
II9ESostWMCfNWvj9dX4oa9ko+KRK5Jk1QS92IryxJ2ORq6Oe6X21aD8Ghpw
wc9zrhPE5vA4WLMEGXPT3SKZ3siYdYNjDBGz3fS04F0gE9pdcmXVOPbsrgEs
H0NwdHTnVT9NCQXsdxoCi2YQjL7HZohx/xFq3/X1E0Auvyen2p6JeBcO9Q0B
Izd2gXTPwiKNwXNYxiz8sjTYIBUPTdsn3Wlivgw1Ei2c82IW2A3CLXqMBCCm
+EhL8wvqlzGGy0Tb0lcbcmu+sn1vZ7yogY4VKCYi9fg28xerQQUIB2dgtYb3
RBl0L3ddgGL65WFHzpF1PiPe3GfebMMZsMrN1sA5HvDD+JL1rAVsyTGIgSw2
tna87oBpxYZJGsF1Cqf3WbDc+7/yZfRHwM7P4HM/pr9RgyjZTesOi/ma4tGk
RrttmLx8anUCjU9wbymNRpT7ZuFKsYd0DETRjaaIdGh80UvdkPvzVuAuw7QS
2KrOisFtg8B1Ee76bh6VELttIDJX1stekzrB1yjqROAbhLXDftr9T6ybCSPF
UH1HokWOhWC7A8VOk7oFMOgWt/LFafZZHIh4wQdt/WEtWv3kiLojjNULEqvs
o1al4wx5og+8gZ6qK2uHKMDjB32NfNLicpoHypWhIGv4n5AMsYGSXOed3Kek
+cLGYVS1YPc6Bx/ZdxFJa2Acy5iJzdqC1PbD8YTLdp9DWfXWiQz96Ywltj23
Ak8q72ftPMgjdRAnj46q2hQxHFVz84LPgI0Yt1GPRJBnUaiBUTlD0WX5j52r
nBgItJDg2t4QvBYbPbcMNoBRIW3Ay6IaoriIlYurIb/lfJyYPyVpUC7TtIAB
RMdMSIYMoG7ZuU+MxSyxZ4ehfkPeLZezfXJ0mE7xoncgxjgDOH9SWq0b0ZkS
arrYxV2Pcw8JXwubZDIe6zkZhPV3WWarJe9UsIOr1wPbn0U+OnA0WqSsvXg5
JQFM9Rx7HP31TiFeBqt1pJ0dexQGgYgWqVRQPf0zOgarOid0syzpi6BsSYU4
7wks2nY1Mxe6b6ssTXssKiL+3U13BaF7X6oEBXsctRjKTX1dxHsrgAHy0EGx
fnpCVHSgcy1tkAkpjBivBOa78+/U0RnK7OfdvHKoH63uyFN38l/sK9s4NZTx
6iZCm6zS53i9xNonVcgwwIIcSUTK6mBbQM8ygv8ddZUB0ufhm/g3yZi5Er5F
v5rShBTjQkLRcvse4g6pkJYNXQhpFilVOUQ6Lx3Un3Yx7OpPJ0EMCgIQ6KPu
BdE+/0DYysVWORl6+GpRRpQs79MD5gBAhZ/gxzgfy/dwz5QP6TXorUOPJEmA
C8qvciT/VCr3sPeTMlN8xxnm95KDhUz45hEGg1Aml+WXHsuH9NTS7WiQ85i/
TMfdpRitkSoVXL5ypbpzD2MZ9/hGOJX8lNRgAP6OPQwRfIPxYXBc6IayZGSD
tMCf8Guc8LvmuUOvkbyZhrlgzSeWyzXYoiZVb9Q/sZx/cpUmzHbjveUhX7Hm
YKpezmh3VzbXIb4nd+yIE6URgU3eAI/j+lGmXYjqoRG8RldV4SANrqAEfTrH
apVf7RInnc1ADku5Vx90JXK3cTJHQwpEmZfnKpxLTnDFRrsMfF3VTa/NoMez
71Rg0MjGBS/F4YSkXFCFbxa++oh1BDMwbTgOGBZXKJY80xERmquSybvQU4Jz
jA6hygTgF/4WFFgvXvZGoomBpcmplGNcp6B51czXAj9UAfkL/MUtQnvmFdd5
oEXAIpLa+SaMVDuXyV7gY8pr2QrwUTYwGDYvVmCmFUsh0BJ6CrBLvfVWr4qL
ci5KjGuKbHg/t3lanWCk6xG9qpsvMuCrYPudSEh7Lq3J+sPMSbSUR1EfOeRX
EFp75BDx6J8yek4SnkfnfGPsOMx3U73LD7PvIDFX8NKvLrHDVB3t0rfikt6b
YXNZwigm0KYWnxF1q6KGqJ3Om2MPcK+ELaB3UGRPJ9JwoKgs2EpIqcGMUfPu
yIP+KZabyaEwQVDtNl8+7ojGYyXQV2HXwFsJd6JXqGpIhsd6av1P7MaRPkjI
Y04Bkt+euYZ4kwDXR2JKL4KqWY/d6Z1QCAN2cYd6i1ZwClGeq1qC/Jmqiaf1
UMuJQVVKQGriIxO0qFsKSqsL7MjJalVQ8179SpugfEGGelE4gvog6Yb73PUE
+jFrSDi3QD50Auzd0Yu5K9fQgnRXxLB5u6ERvVKgUes3nkf5LFn2Ekag0Qar
EeLaRRCImaBguoQ1HkF8QK1Ww0kXAoyHoGJ95jv7/hj2PZ6da2lg9A7SKOhE
1j4H6u7mub1Q85Y4TvvFtu6g/w53RNS7FhRJPOhk8mPJzgLhaF2aSyAFpiYI
eK2xO4fer9GK6Bw2YzEeejhOswgJNwt6sqo4bThbO3blHCtztx6+6zQezs1h
dAm6DlPlIv/2MGyl/2wuSyCf3gGBSYPm1IV98l/QIHW0j9iDLw2YtzJYt4sl
IjOhQNL+9Doxsql2EUY05prHcYBnHZLdKTrhLRliLC8amS02BPyvPdmkJJHg
gS69cFTzGh5mVvID04c/ixSy9R90T9Zneri96dhyT61Qh/Q256b8ucrUoyMB
HoVBnwRKUQOuYvqRxt4CiuO4DNLIJB34gbmZlKc9ousAIh69VCHEHT8DElgy
J1v9Y/WDkLsZ/RIGlM61OM5trVho0jtOeQJxSdrbTmW9ew3Wt4t+BhANDYI9
yyslDGBLSixvSqIbq1wAuZ6PkE3KpCde/ReJ0qWwLcilxp3oeb3MVowsng2M
x+GRwaGmz8X582x3OZo/VxN5EqG7PJMrOs4HzMXay/34/G46ZZceUbUjWjmM
wwEh3ctRk4YXWoQY6ZJ/Bs7WoaJVmRrEavXB0Tmz6gFmLGC1fVtrhNeAl+k1
E+2c25VQB3OrgpXY2WDWpqXJrCAOY5whbaLvaAETMTZ52QccGj+miva2fLr8
bjInJZopG2JeME1LrWEKQMOWRVpsb+qgp8wT6CojG5Uu2dS+AIuOuHvjYcuO
Bno+Zvq3+w0N+43H/K1xfyw6YqTmCUvelJNJ97PTLvqT6ASqqaPwEIMvDF87
6WNu+W6sg+Xv13OXh3Ud1kzPH2syDfw0MEoGNBdCLK3JWuQtPmoS4ha+kuik
YnlZ5AWVPmIJtRt0ZbU4uMvGJuX7pTCPNmivCUXVP5gzYZFDa3yazRZe5NV2
M+p3kosz6htNxrhAH52AsReK+Xyc1D1d9Lcd4OHQAYfgdGYf1z59jnO1YhFP
8nlhR6tvMe571wBSFPLa8nP0vkoqLKdInhIfDq0mNA3pT4OGINucNuhteg1p
rmgFG8lrPjSi+OesllGs9MiH+bGi7V+/otLpIA9GGQhfozRfB6FCPcyGrwXO
Md/QtG4JPSncHN7iZTytCBtnMDch7IYD+w/z80OSN17uJxyfI79gwrceDAY1
DZawCj+djt15HVVNN+TlBxuJT68Gb4iIEfa4Yd8UrduhyvVIVEyrjEA121AF
i5Dp6EGOLWOZcGBqhCOwayZyWfeHVSZg4PIW3FXQmZvfdUT5wd/YjvnsJ6gP
a8Y5XUP9KcQlGBPg3wUK2XToOrXcz0MSFnAjSPGpbDc5uovPCw6g6BQX9hIT
eWhbVWRRwARm0zeYCXd5oKZxHQwvFHWbtydsSLPau8JBvhrzPqJyOIX1kt4s
U02TnRjLfm2FuFj3mlSKhluVOfuVtKrkaPPFORh6F1EVmMNPGV7MP0bXqtFh
tPFRhKFkzqtBH+pZJkuaWeJpntPJrL5EskXXjOa1qyVxtIANTzK7YHfGvsHL
PNAbX0HpQxfnbVnUTJyXKEjPX7sfEzlLuisPwrrhfjSu8ezDXit3O5Oj8tLt
7UOCVQFujCDUYDOdipdd+2EgK/cDqkqIHjKROJERxWPI/CwchFElkxX7bMLM
TvIY7OUKg1GcML5BJXMI1Oa3yyK8Fek+Zxm2IYuceKyt0Wb/+o2ZtrMrcr6b
wza2lHVN8/rSVGni2ONAtOuKKprT6iO72fGKGKoSTt1W5soSBtHj6EhoK2hT
tZ5lNFpFVA4W6Lev5DYSFHLd/0L9ECxeMk5LIGX4nJQj/G4Rq2/6KoerMz0F
LUk6m6oNZNiGdAYvLvqTtxCbxMxf/K4VM8KwB12eC+QEbh4EIZ9cSY6ZogBn
ubvJYM8E6pkUCBiNYM/t1hVEIuafZurhBveVSMGuPU/Q81VYJxFp/Bjh6Ke6
6eqPHxYMgwGkhXzBAHSe3tkFsXsKaOeJ9mK5Us05qN3AtHVnrw+O6sFZ8D2Y
NxW365MCJo/DkWDsQdULvbGKXezEY+ea4Zg3JqHd1YeVQyjXvaD7jfI79oWT
QwkqrjSj8a6uesroCo5JCf5IiZe8EXz/PsY6iPLgoQGTWMhXueZghmmhvo0J
nqnbZJkXp481b1jJVBbqEhGxwaBYjjzDXhVrLtzB+d37BLHuBLmaUGqMAjgk
o17x0RF6gJ+FwYzWBM5tpcVAVQ3F1MZR4AaAw4rt33UCi6eGrduyR+dNev69
wg6A+H5YShe7GaLP1wVfbd1arybKXZfjIeL3GIIUccMd56bakF7KMWdaksNo
waTrUT9IJA3FQ+xekV+RNmJM17onr5FtehJ8xVbVyebBQib6xUB+oVfUb1xn
d07my9wHW2/lG2hAwvJe8hS1QGcVbcHwxMDp4iPvnQHfFEvbKVzlCjtw+9Jo
MB42Y5uuBzRFuPn/ThK80QExUUWklurlWHRhzP72RwQczXXtv8KepNPr/IDf
SSpWlgpvP7WEZjpYjel7tbamuQLOJK41UjXWDmjzRYbTgr/4DG6+Io7L+PLr
IZCYRyMT0g+Iw2IA6sXDTQK54Z+Yrd6Lr6pE9my030pSMUhsccHImxVJYzZd
vXOcQ/0A1In5QQoO5/3XxVMHAtmLTt/HhaoAjpr6IfsMBH6/ehzyGvgrsL59
uoU1KcEP9A1lENB3eNk30m9EGyjJ7LtsZ4dOrj8ILctDpNLAhSWKyvoW5hdR
I/KF1MrxR07h+SbpgQFWa6UprBPOmI0BG4yu0ds6SFrZXt6BOVGnk+s7SBZE
SvlxmsYFvnZ00PnfdquY3+M6JVX0qjGzD4XFSH+L/yRdtIgQxdgWJKBnjfqF
m/m9S96qW01uSm0j8DMmNvSSOQ1tty6V0lEqtTY5EMPHvfFfvTvu0FtFMbQv
unXtlTwz/xi9h/rEdcAS19d0+yhvaPu/miTDWCBk69V1PMYYqNwnG/HvWbSu
0Wno2Xn3UIby1d0gYmiNvgXk3j5nqBrRm0hNZBCqWOp3orlkk1+86snqnKeU
VZc/YUXf47XOk+G92KiW94pjkxob7R/01RqRek869wo8XqcIZOuK5JPHYGbb
pfiba/4LfUVXAwhk8jd0XP8gG+Ez7KnGNvcN3pulqP9zuYfKPAn/B77ebO8g
+EpiMKADLxddeh0S3A9xZsfxSJjPSS2xanWmpwSA8+m+mrzcK8FVIW6ytLkK
iaYHk0UM1bL0+EUyzcn/Ni+qmTxS2n2dwsBPhtHHkRXG/y4pON3adpt8mtph
Vc2kBZCtNHsoWJp4OqsjNulNBrj1gWhBvlrFHExx+O91aotYZwWiA0NPIUGt
nb7cDonN51TbNbTG4gCrW6EpTnI6slrPDE8jI4LUwu1dYEjKjHJoR+ONnscx
dTh4CNwW/fdtJ7fjStzj7NK0m9qBa/ht17mulVgDYwXXAb63r413enfJmkM5
J1q7lLFw5/3Nall/v2H8A97MCTSb2EQkJBGyyV6ndfOgDxjmf+tvcyJQvCwy
AaTckCA2kGxHyk2YMYo3W+P/sTRyR+RYpxcXDtMhLiO17pj4xorHYgMo/fnD
MsAdJbArkP8/pWuFm232N7TpNjedV/8b+wcfFFVCwbrljKmHNsN8NZrKh6qw
5z1kDm9lgx3ObCpN+0lqwhlO9zcwKrUcDW7j9wc/pLBumdf20eJ/3dlWmB27
jF6zU/whoovb8buKSjh2kudCMy2FrrlkaPxFF4FiqU0230/FY8FoQqvnK/KY
o+nGVWSRVBKdhK0UtWe3qIaBOOmsB4vpTqf9znvLsNCV2sPeNIm1M4sC1sBm
cxVyLZcwOTIspjZ1ujaY2JRJEx/lD7PbRzGofiWPhJhMC8+GeEMiJPz6CVrb
hnvATABSKdNBVyot1YgHas6rneSPpI43WfQ+Lfnl3kdoIrEQZDfiBIOpogbu
Tdd+2weAYjGlqtN/N2uWWMG0oooaS+N7CYAU0PLL5jYJ2t4Dn1HZuHOTm6Oy
OYz6xPODddgzxz5RjIi48UbqrqvfHpEWw9hj7qq9d6dPX6wCC7a9TG8depPT
R3FEXVsCACfE4Xkdm5n6A8o7Hj2pMRZ+LW3F07tyA7EdThfhiI2YX17dQ0XX
4gppH5l5Kmjynn0cKb5a7Iw5mypVJC+OP3HUJ7UpV3riZYA5Gs6C/L8VnIyV
I6F8dQt5KVjPHgxU3gbpVt/eNSFSdCGiBpJtMO6L+EZsd8dKvymitKmst2Lh
UDDB8X8BdJ9ddS5j1RiNCmMRcYUTwCX8DWhFQhEK3pne1vS8F/5+Q5oTNkDA
j33esxtS9MOP4K7qo4vF5Nhlkmj8F6MHGDLmOVRmtNs3W2EoKeMRN0f6kppd
d5/j+0d+9dhBhA9PLxo/l7urbrQB+rt5vkig5PlTO5wN7zZxSKh3sv+VwMjO
ml3wsaAWbqXxYiBaziiChadHDW77zxaE+bvxPfoV41oaYjCP5ALLY0YYnut8
9IMpc5ooV0QkZhfRM9jj31xfPSsLrINQ+5BbIRKiwYradnUMYRV2jKbNAFNq
yoMR4FTs04khog+m6aSCvtcIBFjqek/x9GV2Q4OKLXd3qoC/8p2x5rAkTQP+
4guvqLCvhOVA9E8ZF4uJEXlUinLQmQdFIqSoKZCqKLrh2Rxtkck27IRjnRoz
pekquRM7TS8ubkY6yUCFzPiDwCtLjJZrPMOz5T3H8ta1QFgWlhr+1gTBVRvO
eMk0TyytyZdgZUiMfrIgfykvzKvgeejvhROeX8o/LBomJsxSGnt8T83JyYo4
+qhjTqURBmbTW02I2uCnXXnQ45WoVDuKf2JMwP1OohT2LPZ8rFwBkLGo2i32
LnwMeuJ3mkYdKBltD/Dg4TI7SfI4HUPe7/Hk5RLVBdIm2SQvMRheNUwCeKz9
xbeDArBGIyPbm9cs6+HGo5+HKepV1w1p3piBkBjwKWPJ91W/jbq0/yocvhA6
1WAuBOau7REXQ+oPhssqWsxKETJVmnnOwUJeZ+Vegp4OnBXuzGVva5aht6NN
LJ802hCyOr+2j/Vi5wrUBK+PwlLEWSsLTOzMj852JmMJBGiLsW2SIj+jP2N5
hoqAkJRxX95rR2l3aF48/qWkxmCDXe+dlqPJ+hPwCtLLxmonb5jP+lnRG3zJ
nvW61XrZWUewYwv9ZWbRmnq//kq1GgXF2+YE25i2u08dseHDO/pZeVJuCUf+
0Qic2b/KUSHGi1Ml+GZKnyrwrNxwZ/IoxpjsvOSdXuPD9KFOhgZqGlNEbIpj
AuDXjZ6F9DlW+Vv8R4YeDkuFqG+KPJnxOjo92YfS38GeAA0u9oecS7JeXRsK
oz5RmjjePpl7Jl+zZh6AoD+uTbyVtiazaUrr0ZrMVc3IPpDLmm9vfw15lVHl
xlL9Kbm+GfeLMO9z/qq2otB5M/YGshD+MSdpfMnczRRBgKjdC17uFdU8cj5r
zFDTtGbL9Lk9LN3kBbCW4rWBEBRrP18IIHl7zlevVnTF6ZaASr0DCXVAk5tF
7bcTy5He7XOiiIKTVOBbeicwjvSIxCwIr6LZKyuKqww6/5d+AWK8y+edEAbI
ZV0i5tTuwP2pBGBa417LA1x6368SnWvkJ8LYl4pADCtir3p/OKuzvZPNt3Da
s5JBzw6LBxxtslvSLanyvNKpL2iGFClIMygdcM23HI6w8gL5/OZPFSOSSdEG
ehSRW3EbajMYVisIu3oi7Lpldb1RjedN2zGlUrkmqcarylpbcRNC1D4ERYof
RQfaEwDdCk8B4whyb5zjRfv9PpNc7lWtOvBUK8whEthqvSwvvQUdJkbjokmN
QLf4FlyKg5VwV0bkn1FvTnMIGddVs9cvtBrUM0/mJAn8KUMijnafZxXXOIYJ
0g1eHKpiEc3DkfL/tfSeE1iJnvUOh5UsrcdDwbwKluV/FnZ+sHqUYgeBHMIp
tQ2U/LXUNmgqPENJzck5dcdqsRh5yBR+DkCehQ5RjVl6JxBEplj7PYqBzQXb
k2YtmmddKJ90OpSmHwMgj2OphfAujRe4fnU4wnmDmRjT6VbMlNqxf4LrXYQi
z5OiuBg+cRKtbdVzhfVnwLaQVPOvSwTs1cPXxop5QPFxkbfr/N71LgMnyHaN
o1JXitt+AX8NDealjRP+8pVQR7KeySBXao93PSP+hTZtIFiscoYqti7Nh5Co
tja4Jky23B101yxKf1B5Uj4Mtw4NPZL22aERpXItcfjURyV5iJYLPJrTL5eS
HvjOEeRwmpro+8eIpRxASG4UFiCgBQP9MnMjf9V105xyxkQL5bXtqfMdrl/8
RUT9hOv8SOa+vhlnjpS4nz4LhT8UHAz/WkEhhLXtGJNEoXecwUQ64E4cePl9
Oyj5LSXX4IPNpSsl8s40XqVJjXkHxlFO+14nA1ZeZgQf21ZpdIKQRjkhf6Tb
WnxDjQEeHE9SeaD6aiN+2HTimrVZVDA8fhG8qoiqqe+2P6FGJ+TkfWG3PF+8
u5WT/aI4ho92sW0dQfUIaMX2Fnm32mM084wu/9yw/HXOO+f3Z0H66Izb9U0X
HCHf+CGAxJ8Amu+T03sgtSt6bes0Pi4ckvqy8to+V7x4bdGc5ko29CvJ6NdE
kPE/C2x9DB90deIsmTP736mXNNlUd7vwJgp4l0rYsoULeZBv8O9fnomTCTG0
KpK3dXX5xa1lSW/tCq7u+ZtSiVVeR1NPP3Ch4DAfWpHmLEKQeWAYPXUlhkJ7
1v6gth/5PVmyLPvMoRFyzNzUnnM7Df4beNbeDXmaO+Yw619nL9zAQzxlvYoq
DYEViFTOsJ7sPCjVWGfz0O+TAx6PaoDiz5jNJ7tkTHOer85Wz6eGy8eXD0X8
Ebaqmw1/XLf+mwO1rFdpilrfP0uBJ140+j5mIzDmMGUvHy3uAcZkDWTXzs1r
p48mfgrZtS/RberONvFkNhz2dQei2WMHRagcnj0boVSoyscTrrr++1Mvf4eK
WDACgDdW9NItl8PYEGC7RoyedbGQQdroRaOyEiY0dDQFnUBiqeCKa4CqxuVp
T9eZ0tY+G4BLC3jc4WXHczkYE8hcB7twBE3T9j2tcL8lmuccSoQniZGkPUUm
CCMaA2PLPdMWXb+csxHUuKtX5Ksa6ciWoqWQ8NhyEKqQ4GjVaO0pqEbtXqCb
zacYm7DQBIFfccMbYq7+ACJPBDy2OHbtz440GKpm17ZwOxNIO9xYURE5Mwcl
oI3HMmIRdmBi4bmYXWXdyI9H+pyHwydCyeLUqFYmbgY5hj7Pc8Vq0jac2lWn
6tuxbWhsXtjKA/kmMzw7EDrW4hS6pvV/898KvJW8Yc3cKCXKf26EQPG8UVsk
swkIB8+jL8O0g8FLNU6JDlnvSGhrRQObdrlTYK0e2N8yi8DU54qQxkvMkrBP
YQVZ4RVcXjuGbXxR5783CzgBG1yFQ80iyC18pgQ9XkOIf0hv3KfnM+GqZaPy
zaJ/1tXDfsVbzgD4dM0J2Vy/teA1UPR4h1QU8RLgSOMqRi1LMO4xpneMVucr
5p60N7hYByqgbHM2L3wjpGI/dV6UeEJLE1EwocruCEnZoaabwIgMkCh2XxO7
kUWrBghgRqx1HwAdutAbpP5gzNjxcSupCEnzfCiAZ7jaKe/QAPEZA9p1FBPz
mmHEhy6dmsgmFd7AFuc6KsyD+ydZq9meBHjXZWFTZgSoSZIs3yHVgOxddAhO
UbvNt9xtxKyib3wtawX1+RjM8viOzocTJ7ldBJf+RcRx26VbmblJDNv7/o1K
rpFqaa6aCFSy1qkUhLNpm99zxTIkgQK52BrCoRC7/q7gltrZs+0RYN5MT2u/
qCRbM0DfbwV+VIlQ2EIwrXgHz0l9BKMNyf7zzHUkb58aUWlCYL4G9dU3ZqM7
R/MZkNVMYSqES0oWszJEbUzFqCHfUxieEvw2nfjxgdLzAX4vyUR5OAPAdngw
NVfh1OskbmJbyrv+xW9STj5Jr3pOLrN6jZhiesxAxybpUang4uL5odCfN0vd
k4VjKXsZkAnDAZHUSxsMf1//swRITTcPbQmbNgiDBpMZMK8CEmKqicz//XrV
EDQb6zfzrxdSChwUqY0QlUeGQJCZ9HAuUGbYrl8LMagQyh/RIo+3RXLWgpw+
Ce//tx69VXkd2dWc350mV/bthJFTz5dMBaBBPKo7rmXOUdDqYyGzMKjUKZTb
RtGrlxavwBhRBfOIfNStqWy7CRxGECax4jhuePfDazejMaEMqegFY+tT/WTc
PCyzCT+eZLQyrRLiRk6qwVjPKam0EC8Ub9YuAwEUHPvPGAI/3WF9cejAT8d0
gKuucGJHNUbl6Sg2SNFz/b6yY8K/Vqz6t9hstRPqij7U7xHVlp74G9sObR+S
Y8d6GHkjfIUiN6bm4adfBP593dBS1sASEH/7Bi/wr7QO6mp9x9oZifDYXyZs
H1QGB+/YZWEgpHZqOmpCO4jq+c+gBFsxZD6DsHTAUfO0+EUe1ONkpLh9v016
UnYF6aEnMS2BIUl+cyWtfYlzU6CEM6So8YwxPu+g8vE0ve7kJm4Bmbv76aer
Bjt3WXzbVfK92kRrHmaac+Uh6TaNff2P199FQTsDnf4G/uOeHgUDQ15PHcfk
O6DZA+u2nLkGGWfN+eC7sr55QpX+XxKdtBtv/Ud6qpEgVc8kqd1qLs6UBle8
xAFCwHoJ/ZcYAicXtBwEdASluLWx7GlBkkGNenIOdVA0rnbUVY+BNbO+UakW
RTHcbNMxctLeEqGeBAmTMVIJmbDI7hPl9APXqOb+XAbAOqd5y3CGc/qY7x9K
gMgjGEsuluWpkbEVxxnnCT7EzRddNsJl8DOE9jTNBoJ9/eXdDNZOk8cdbDcO
+LvNikKBhjN3ZLUUeHTBC1tMyk998wvQCUYYTaI+jTM9idvmBlIXE9wHmEzj
xX5MbyHDJDDvMCQ5ECSF8FyKWi7EcCEmhUL1I5Kz4NGLScKtg4Y4hksGBpbj
yeSaSUlAuYWSPGX6kZFrtKfbGM1FCKDdW0er0KJ+lgkdB0KWbyYaEoJhd8Df
/u06xNPhw9Gq9X+UAn2pFKCLZr0/t+T+E8c5aDx1Q9yTV9V470x1fF8LoqZL
m5Wp5ksN3pNyqTVFTuzHZlfZ6uOzljoa3xVrTApKSO09dSRxq3Ud/8DLSlaF
He5Q+wkTKeH2LcyQ2mG9sruwuXscCu0ZGHECqa/yPk0sE5TH+y5xszGvGDv8
zf5Qt3thzq79sLA/eJZu9DcjAGBeDkNChbLAG8Ov4Hu0z/utIrJikTIJCXvC
P7DTB/JkyWh7rZgPpSFiZQA8dMYblwXqHub7APxgg5JLmtC+FKoJOAXfh/Up
jWEXCly0WnYVG8ZSYQ==

`pragma protect end_protected
