// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
nZTP5OHjLqt0SEURt/xKPWxVetHaQpzhGGW50cHAZcTu0y4X5pCp1l5sfsVhMM9q
811Oid5TTno4fZAkNxkr6UoF2fVsrfXufwD+zCozMIG708yBiHo7wPSEW1EpVoMs
ILxzza258lQh9Ug/L6wkE+0MloDM1A3qaMkvEn0+e+s=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 32288 )
`pragma protect data_block
vqv6NL2bHaj6KQkC74Z0TbUOVj2KC4aadunFVZmskLJOpyQGsfEygoK+yyp38lGh
lp5u2G0KWARg+HUxEonUcX+IiMJ5THf33GseJ0qFBysOLVZOguLA6z3YUoEDz9q2
wGkIncg1PgHyvkoRBZLr56iD36lIkKBVurFiAhDkRcZHzuqjor68C8V3chGznYwJ
Nj3/Js/NBA0HnZPJuB/bYBZF/bds/fxdAPOOlsAOAhId4B+WwezrT1vBH9QRhbO9
p8TLSfleAhk9u84nx7dYU+qhKWiTE0y90dRtT/qwvoZhizKM7VUd/RozB9PVjd6t
IMvJDKvTHpyNLqNZLWSTf7EJieZUMcYkYlD788r+0DuncMme3GUmMeYW9AhR2/Z8
Wau0wJ7jPBRx1mJjrYK16oSG/0Ag5YXL5j2j1nmW8Uwz1KocOloRYGxLKlbruBMk
RxTJ+Engl/SBvmPFt519lgjqAbcRk4LEtLElCuuu36iRNz/1/1J7+awYt/q6SusN
7jXHDw6ywEBlDfUID2LXlG7fiKxSlDzf8NLk6rzmjK9BAvQDlaK8KBgUGsMbkO+l
BZ9oEPwcYH8lRAiAHvyyxZt+kFgptJiswRMct3R7wHPmkTJs1wltjcPMcGO2RBHk
sDS4gFbAhI2/PWclBUqMpcZEMUI8ZkXm1fte/F9g7eOLwJwQIqRK0b7NcAvotX9m
TgNIYFGd6mxehomfb22UGNujxKFgQ8qFXg6uZ9pBEvetqOHxfVC9AqDADTL7RxAS
Tx6klvW+WYn9x4U6Hq+NGvlBCrOyWJpu8A+CnAV3V1caqKjrB0m/Eiux+v1L9zzo
WmQs+VRUdEEaYwzV5eK80osYexm+N9fTM+neGcAbTLz75+XLFN/xFoQTHlrmVIZr
QDoNq/VQ/cq380orpqeMkZ6gqQI4pTslK5KGiIu99gvzsCGE/c6u6fJO9FT4bvNB
qqn27Fcr5gLHHWaHMzvwK+A37pnAXF5V9dwyOlUhlft5BVN3dxpNP1nbwuPux0dT
i9j3h5TIzmYefQ8tJLpdjJeZwNJppEmrtPHc3giJee0bM7DxhS9JPDflEdmqPqdB
ZqYFmFt4EBuBMo2KYUFVsXL3WoFYryi0kZXpgV19yvtJB7wSeGV1ss15iHqvIO2r
sxezUZA2S05WAOJs/rATJ37UYxFUq8dFXtAoQz/+bmxsu+HLmfAtqb05TErd/iem
QW6WCfa1Z9x0cHAfzjUj9O7Ye69Qd6Rrn3+TX5EVT8Qfh1XpmL1Gdpq1wjhBxv7G
NoCgZd+i0tgvkV6yM1nLOFc4ytREE3uGIKHbCcchv0xGnXj5XnxJVT02TjF5dHMX
Q5M1jG40bt3tbNJ+KGupzGtZDkt61894soesc5xd/DoIs78aE18mcq6w+zwqA5uV
IL65fuqmTkRYs/P9F8f52aafKXdpsJzmN3Mt1/fMwQbmVR+qdZpxUkxudkCGL4/j
YrYrfrzdRv9IImro+mZoyM5L/i6oc3EIVQJsodQMltKxqvYaXcNdTUEr8JUr4AdD
JBBqpT8CBq6EY3TS3Y3uXlV152i+/cZzPOWnvVUlT3hLatpUebtVIh4EY5X995Fa
Q2Eqg6uM3NSDkpEY7xfQ1MF7MED6z2dgg/ewG9jNKsa9vrJY8sGrTqIK98NwR4cS
kSxa8GE7IXXOMKKux0YXEdFlugDAaT0Xyjic3aArDobNGSAYC+ZIYD6oH8ZpY178
1MKGB9ofrDXDaQLLhLbvCRG7VbPrdLLA9X+YPAeXqWPfz8y6KYv9H6+wlo6M3ZKz
SRauktmbLNm7mUDcSXKj910LaHFwueS62kLfE7ICEkqhVBoJXqGetEAQHGhVKN1Y
c/Hp7dZvGfC2Gs9ivG1LhrXzC7YBB1H9Jx05mFWcNcQh4xdiobGkKoWPesQEgjFt
a32VOHzSie7ToojXOzaGnccQk09bqVE82M683MhXbGnVsTGoWT1T7QYHodu2ch2V
USlGHlqNVZAwggAyQcv4crqUVM6SUxvrUcvdEEKttbLvUADys+SSImtlDfKl2ghL
MzrQ/T8xeMPl32YkOpX4d71HTX37mi4cPaFF6DOQVlA29fqMTqS/rCgFWK/gfGL9
cpOwulNWQxBBABVzgG2pdWKbuwxPy83WewkkniRc53TiNASCNiUJwNUXtdEYpGas
mbgHDKRMcQA4GsmLGmR+4U0lie/5nOu5QLwAIVJpVf4/PkpknWlTF4nyKgBlsqgD
rOmfDXyO+GG9lXWweMAiVM2+JNgg74W6uwDr+B6fsnW1BbvYI88DDp7Uh0kcvbPr
Bp0Mdq2mYhbaEUMYNmkN+3sa4OT6lXcfuIWO7FiYPBIVKAhaG+Ph1UMac8Rl5VwF
Ul6mh9p9kcgQdX/QFXFU5XAFtC6feyDipjhE44gjCFXeRn5Aw7il7LwuTyrJ07HL
wt3vbWcqUqdglqQzsRe3Fsz8Bte2LPiMxrNkCpQyfxmGfhfdjlz8Bs/0AIULRmDl
XlcetQfsRKNgVh9Yj7hYKQrJ4r/ZfK+pfbnrUqEfnMev2s7wECWVPrP0mf/AHLjO
a4GOmqg9GkixwcwZxA4ysJWF+GcVdiTC94YkCEZuvUOfNvo2odPR0gR5PqvGsJKF
8J/w3mqKZRz9AKOkFOpSXF/5EhQdA+7IBJsOAcnTWoFOpRMWQRF0sAt1uSVHVaKC
pCENJ3znoKJNSf5T5Y5O6v+uOszQ8Z3M7xpmCMaSFIKcnt3XujDxNfbXuTjLm0x3
6yk8s3nBS7ueVKd+MpwPpePB9vz1gdE/yVEdLDw+ZAzHz2Ga/PjPpTiKPMjF5iJT
Wclwru8ZkOs6v450OyQrsXYwcUKDi5IhhUyvHkHxvBghXkahm8ZmYus9wzadH4CA
7G9w1VvDlxYOa6Ym1yOhjxXY4uokgl1JOMT45o2vHZoRtdLzp78Dj1tvE7K8ya8h
1seCrDerDVQsbMt1M1RKmg7vaB3SzHQ3dCP12oo82eJAVflDS8SiT/TlpzJw3Yzm
co/iuxu8dpgadXHBvk/PcKFfpfsAoET7h387iRRABBFAr0gW5KPwHxe3QQ5796hM
h21l8b7DyvOxar84OfmE3RkdPecTTsReOeXeu/4j3oX4BVzS4fcGRSCz8iViIw02
TbDunWvYiXj+kK8xseGR2MROXhTfsmCYGmY6SnxAcSXMxSwc9E2yU27NbZ4mW1ds
4CZy/hrmqf1N78/OgT41n12BaEfKGmIkZtxODK8zpNxQSQiokM4RWaWXck4Bx1C+
YO/iTvCLku//K+MYLtjnyURAMhBDKKyLUvqJ807lLgSiSa/XVcqgiCnSQbLLVwnC
y6HURxax0rflzDk6m1XVxzxq2ay5SMsF1auPOlpq4JUOzLLFjFm2umtHNbxgVLFJ
Wba73UAESWhPq87nYtU3AFUIfACTQolk98DwR1pqokJKRn7zFWUaS9Xu8M/QBGNF
SW7nC9z1TuUxsvWx2AOrwE/6dL2vF//wQcwueNOA7dTJlUdMkwt9pPrFJ2FBYqkv
bB+LnjoEaQxiJSS6mrLOLy6kiPigKjlsqzuXBmAatikdU9a9TfFK6sKGIJpW0XXE
MO9h93vsgbf4AwGRl8mHomNivgkJ/NTqQdwyg66ZrdNrWmekvvoAyGZI9EKCMFeb
BZrjuQbdCusff+ThtR7VpZ3AwqMZByVygW9TWS7lO/30AsExt5wxNTZN6MmpbbUW
A/oYheiGUasTALLS691qX15Dt+8y0lzlng+53t5wa8bZWAGffoNjSlaAbbp9xKxE
rmXzMSmf/gL/4ibl4XRH7c5CcWHFo78SoM30dEG7nXmDll40Rm5WG3YLgwSrjit5
BViSfMpsE5feLR4f5N34H8XFPCObfDNcRXz/qwHgmjl3/9Mw3FM0Ehn8GIawao1b
0JleZL2Uj+BussQ6YknzHZlKBmO8lt32gdNeObXwCQq8hM2ldMIRJdujLyzsKMAo
UDVfe4GlkAA/m0qwRN7jgnc8ctQkd6DFGfX4pYY35BxVFZTZh8Du1klNA5OPdDfy
J8cfd2b0tCpvO7IVKhysj1AJiw9gULckC5RCcv6vVqif5nBYP6KSZ9jXlTujbvFC
1zvndnBzZvUMgHPzlx+YjEm3H24Wt6InX1kJlEMmbZkNT80R5N+/JRVVMwT1c9MD
7ltu+dkDlzrOyC8wJ5yp6eBghPZktc25MQaOgZO0QNQWiy3pGc6Ot5DbZg/65Kvw
XkLAud8JjSrUdkv+8q7EGt7a2es2OkE73MFOjh6om+Jwt3T2lIuSOh5vu4eL4h+0
sGzZ0ZN1cSq1PhRZtZZwW+y3nJJZL1ApNo8b61712u1+QHTMf58yCsJuo0R8YXA3
CnBjzMJt9PtmjdITNQq+LDD3rcs7BDannOYGGRkv8pGGOFEpxbFmw7ke/EJYCeIL
iGsUhwMzJbF79QHtc2tDH1tHs38JQBpgayF9vKXbEzNJPRFYZ3foUOZ02ITyxON2
g5TL8AdASktQEFHyL5kUSA4Y8zlRC8KoPIXUSMdIcejBmrW6U1Ix4UXkHPZ+BUgc
YZcxZAsVoqhCgVlTOFtzio/ZX7zL0jwpLgmQIjSB/3HMJ6+fjQ1qrp4HlUvoZaNY
eTrtrK1e5EEZTZ6jGuR38ibaxBGvo0eu51LqaJp5DpVgE4lIEoOqaIF5api7oPOY
909wfSfrka9NhJbVm0Q8jewNFJGQN/coHpR0uGUoZOhZH9xWomUgGNZ8nh9fTPCV
ypr2iAYbNjuY8+0/Xd8JoEBWuhyU4WqtGA4rKvMu/J0w89mq650XyC7dB45dul+Q
QXYIB8Gnkh+r6J21YFBOA8OXDcZlpiMI2Zdn6fK2BMymGFm4EWJarBZF4Isk0XoH
xbweQTeoCBNR51GUNxpJ0EAPXtUrlT2AeJmfgB3g5PPBf4dTCHc/iWqshAtS/P/R
JQkzgx8pjVjDxe0emz0BLmveAbx1UwHu0t4hKhaB4XzXdtsDeT7cjHA1hbKdL1BG
2uXyFlO3s96TyBC1mB+hEVIMIFMPYQRJ7S93MVh5iMUbUnuq1o6H7fpdc0lfplVU
oWA9U+poLoUQn18HuDIIptLbjkUjFusvDWz2zPoawhEWHKOOfZbMy02WwMDKDZVJ
7VGZX16aieN9nMxlMRpKefKQSJdbu4IpaFeXzCCVjS4/pi2jBefkV6bclzhGSXrJ
q0f/k3nL8IO4+8ikq+0lSE8fmJUffL+Tb9G9e6WjE1w7j6CAaFlRbnL7ZVxgb76n
FnG9VIWeFt7NHd0MFpOTPhvE55eL0Oqd7YTRcltwJ/+d4M11R97sZrNYNZ6I0+zW
E03I4AVOgw8cIH0H/eUoEI8ClTr9KwzOSRXf0MsW/nNoJpFeAIPU241ogfXGRvLJ
BLCSN6KsIDoZLtExIbD1X+Tn1f6EqsfPPjacUmlas4/fVl3Lwqnx/v6I+NCD0vKe
X+4ksu6Hj8AwNdeigJF+mB3TNopP2cRLWkGAACaDMij3ui4cZvCn7MYF8a8+0VRY
uxjxaLmmS2T1DBMRxO1i0s5HQcsAqzOXB3WNnpHPbBHSjeGydAPleejM6nIGxPDM
qYAzx/xg+PYYJZfVcWca8ZwWM5jzSqeu4byVSuxBRTiJUZmTcFzXVipfNR37gOt3
L2fMWT9J6+puO8xWYnOxr34n6q0QTQo2/Y1giKPfF5vqFm3hnvmNfFR3EGztyzFT
vfQTfOUAFtG2oRI1d9U9nYRQxC4YBkyeOZUopeDORRjccHU0RgbGbRt6lRA9pwuF
4t1Ta1lX88rhYYp+Ohe+XVX31XVr5hyuN0Twp1gWuKI1UbtYdNbvpzpddL9Jm5ra
ktfRJgIVoI95F3SANG9poH00jEILcRnZaJ0pY2tdtBpUHwkMvQ1G/fVmX8B7PcGo
mwDX7U+lHIUiwDnDVJjD2A7gqRU+aRxy4vQ2AgiONqbIjJ170SglaQISk7TJMq0C
kHfjUK3iyOaSXrCk8oPZLJC8kCC1/3R/4Az6rHg5bBlL729E4fuKFa5H9BcA92ty
M4n3BwUqcnnQ74Y/1RiQnL//agLTqSyCOkGFs55do4J8mHDoCTZuuj4sdEI+Nxqu
N1FzcSJeQl/c72iz024kOhjF1EPrQhwtrNh1gKBvHllBm82hiUp4pRTUusQZxzuO
yN1XHpofUK1jqwDZNAhYr+9kfouRRH1yJLW2AoLCxxFBioqOrL1sAZ5dHhKaN4OQ
ZbVmxj3YucMjYRiHH29hWYs65GHAhnmMvLIN69XiKQ7iLlX9nYZk9ZEx+yaWHDWg
d8sKv4Symh2+p1Fn0tf2dBU8PPXuKGmtv1RTUY9icFCO6T8jp7a2VWTiexrh4Xsw
gYvN2ksqWEl1H0jZgfHyekLQv0Bxnpb7qpREXMXUym3uiM7t0g5EBXCZh2eUftKF
m7thRZ+4brEA3xTXQ0hG+FnLGtzIRflncyjsTokesoHL6GPHAG31bXAy2j6xsoWV
68sAfzEEDZoAuiv4be0FmYXps3U5jwH5cV4k5Mr/4tYeGMl1m5rrCD1JDJlK674N
7YwoBnL41A5sYj2jZGTY/j3NMgmYyWYsJ49dcjwaR6/f0tPtGju0P6n1xXHQHVND
lE1Q9BFM4h+4jxz0td0k5sY/KEKQloyMRuNnZ5n7yZJGpzUuqQFQ16enKYxInc1H
+jDqLLdoQy9hrePvbj7d4v+T//AB+Ny/j87w2yGjTuTnAKXGy/D8SdWmp3XIXO1A
8esJhkxthZ76bOjIztZ/ofR6eBs1D+8C/8gODEfpmIv+SqBo0gGWyKN7YlDGtVXI
1y40t+BlaTbG12+64LJ4pqmM9Fp2mow54z6mPZmBMYKlDCULszttDhZF6Mr11ix2
/UVtEiVpJVO0x0XwkXhNoAR8w37KehAiT8ozFMbM3siFSM7fR6aSleYlBLfWZ+1g
tqpqb9P4g7p0yK9dUZpxBSaOd7nb3JOcX9U9jT4Bm0i6y8HVKpC5bCEb9MZ7puhd
+Hf0r+dBGGHJUqSENvXnk/kxchVjIv68nAVKhnvBc/Q4GSd6wNDgJOs47/BdTmXC
9dlZW8u51Bp5E509QVnj3mAxhI7EZPrnHgmJEP4hnJiEi2AznKz9DkgZxa1Myrd3
EWgD+E6/1GJjN6mggyCJDralgSMVwsBlohUJhPxjvu+Mbq1aYgZcf0Qn0+Rc7cQ2
fvnqls3rYJVqQvO0cTm19LT4O9NGQ2FpzC6AGBkEyyFJBR/d7RU6hQPNEPNA/7JA
QsLbgGGPaJ0hrsAkmO98DH/+YxYyfYOJAdBUHBjP+KcYSLlYA7qWrWnv0Qz1qEA5
k9XFOmVTbHYMVkCD8AB5X4y56ZHZQmypOKYdZ5qHcdcXbI6gm6C5pM1hikCZ6Nh8
XliiKVoC9LDbe423G+kxUT+2B7qBckNkvtMFZ1weX9XnQPNmpfqU7Rw/w9zWMCk5
g8h9aBuA/Z71jl8RLjxN7ZXKCo/I/HAKgzLDttrbJUCtio/7UGmg8dr60hKDL3SX
gNwjUZI82VPvtuVGczjdfrgl7rtKCmw2g3D5UdyB4/tAfixNpPW22sjkWBlgyPmI
VrUvawRZp5SiNbE4HoYI+tMpjnrGMPGM0p97cS51UG5exCiFkXyqFlCLIZRgjWEY
Z54JSx82bRMjQZuaRtjaVSiNxWv9+/aqg86Y5cm/1RHCwJQoeYiB8EZmwTXoLy55
MJYQW/fb3ggfe+P+14TLGbV+junCCHba5oN89cZ57WRg/SaAks2ez8KO/oiLHLr3
2DkEbr6boRo2BxAp1zjvOotbR20RjLvhOHrzpkJrW6A11zTj7ObxULuV22tfBqso
lFRI2JBtGqQheevH0yGgtK3bgNAVjYMYQIHwVSNNdWsWijgLTke9yAmtYSlKlDzI
BcrJYFoeWSAuaoPU15QYUKOMv/4+r7eTVkKdtbTChfW/+H3+i8cjKV4yoJGSDGts
rAwtTZ3/feTZB+WNGx/J7UnVZCeIqUZTHTUeG6Yzlxi+COVWgUnixJr9v9xqPl6O
1+wSU9OixXwcpra5aqUcG5YsXaEdgPbd9fUSkqhgmcBwswPxwrhrN5wkhAF5T6Pg
tBR76i/07wbbkqJoGO1jwNOZwkS303n2ujSCRfu1HL8w9WTN9zO/i2odA74qe1GO
B5AkX1G/odIu9q4xljMPmS0WUS62YJQJFMA5g+O1jTj2K8H3aVmRSa5c0NACuTGZ
X7ctoC0UhUvKzyAumTyeSH0QMq1iXPu68GX6MYmT8dIll5bvxMrSOaU2uDm9e9HO
zmiB+yQmnZQQyNBI+G40SlLztniU/HXzVeIF1n30FLoKl1Vek+xIsbXIEkYJ+RJa
0pOiOpeVLgobre4Gq4Um5E+9iBOIwZwVe9VDYRgNy79PzEuK3k6AQ8vSWHhQy+Lz
Ve7Nx2ocxNr7TmwQI+uBzVQo0ugr6OUqaczQAg5ub02MVbA2bC302F5CNX7Vhaih
SvKXCSncV+VRZPrdtBe+6iiNp6F6Iur7HPTKvvu+1utU0Y1TmwsuqqsJZjOay/Rz
kNs9VV9hJQp8D70puoKPsjjvwel/w/K3cbYlu/pvxlrl+HrB8hM2z/XFWF7pz/jh
TrzTS2MfLevMvxA1UuIpZkJB599fMZYl1xSwveOTTjSI1zkc713f2aiKY8MJnxf4
PMgUlZFa62YRNaa7d5JQTsF62ziCQXU27vSrniXvG35obknm3LwCX7Qj4QkUhn/X
S1lWRN2RPn1SH/4ouMQ77LpKrefyTT1i4MTJ+gZdpDCTO0UecAIn7eVZKB8mb4wT
AjSVFlvAxmA+Iv9NwdQCznTGQoQvCiUoYYr9QkT3qKqzBGMjM99Zg4ShJ0uTwODn
qXqvsS7nVPmUc1Ww7JeU5JjgkYYeUEwlKnw8uGnfM9Ve8eRcstXQGoV9lqya/bSM
FRIcifqzpB99N2yharVUCaP7EVeaIGigdozYQNEniS9LVeqN5WVb4V6D8KlhHDVf
J4eMtnDoBip/DBSOaLo645ghaW3cvsUn2mPmMRr498f8P1+LqU3rnbpKPDuoN2DX
10hu5qPnWU3v2mPHCD5FCsi5gyqmRjaTFgPDzoCN1Txn4LC+EfWx5freAC+mCAkb
GxBowKDJmypZGmMGWdKVyvz+5A3vXhj+G5kJSQgWtBOfpDtP7+SqvNtTcPEvpdak
lSdn/+2Z1b+F9267fCJ5FED6W1o7vQiVzJn7oOu30EKWJAVeZYCfq3Zyh4USlKZl
Il7NUWo8qcy07LFPz4m2xusODfPFc1e7dAV5VkUN9E7jJzzPeKX/XkA+gXw135mT
tFPfaP7ACXS6GvJE/FxxuPTTofWo6z4HAOGXcojrsz4QrKtZpV+enhbvHE7CzZlJ
xdchhijmVlvkR3urTYKQooyQ758uUh8zUzOv0dfrW7JGMONbUwiV5YOrxD+gIzoT
zCunfVQIxFnVJ3FDuj8GraCPjiw1rQanvs3v5mj0GD7UL7qpMjiO4ZTTv1UiU/8q
Qr4T3tBf1Du8csc/zAq2FIO0CjCHOXzi/8DM6LfeU+iHuTieVjGwM04L27EBmBPn
1k1VRlvnpEDgyIge4AO+q20EZ9dEJROqo9tt2xPNbvtuIBGm70StCPKE0D359icf
FtvHzbUvQjRSwYBO1/Wq0pwiz7i4fEXNMfUj9NIJigtLE2tH+UUqX97QUh8oT8VB
sE89GYHW6WYR8OAYLPW0hcY6cOXnnw/hSeyWdN+VA2ByaDMug5IunUfaHT+hs2sN
K/Onve8xt9E46nBw+zr5HSrq95tkqwQ891N8vV6nMGXtL/OrkjI+evdohF6TiXB+
UGKTQbk9laScb+bgfBX/fDg7MiEfEP3/jpOT81rd8Hbu69AB+DagxHnS2ojJ2FyQ
h7CJyCUEZtpFufGic8mTR3AEIDRlVoQF8QXxWjI9ZhE6dDuSVc3CaG7b3odANI3/
9GNM5thXp/cCCQcuL8JNx5kdZVFVYw7ozowO/kV9KyscFQ1+4v78JVcqgATuUaxW
eA5ZlJVUQahS+qqRaNQWGpDDRErr28OTZvok7U8AnoOoKlGeSRePD6bXe61d/C75
UZv86swCLt7m73m9om+7FKowp8xkATCb+LiLKjnEvjPaq0fVYB2zXkdrqaf134TB
JQwJqOY9yNjlFY3u1Wa06AokVQJpCWWbfGUDdmP8p64j/W6tbxLX6FxkP100q2jh
pNiNndrDXf50Ca024nPOqsra5vP76jn9ufvumftBsJpfYJ1Rhg01IuWm7OVk8CSo
8M2iriB9rZejGTD+O78P27m3pok9JlMpIPphnr1y9UO+y1KAiZTPd8BQ3zPmFegH
yd+/4lenUm1Yqx3UrQ4gWILes+2obPmzGFm7v2zhcaQlbbzKB4I6x36xCC3Hyeiz
nRRr5H6uncbEjmCOrvaH9zi3bqF9KAU1aCJRZFOpLy3lbSMhQcM3U0ppqMxySqrt
GKxrrjDXNZEinHDRfDdm3v/m5D+sdXZRhFZpErDIhEX4mNSs8Gt58u/JW3HxvGXY
iGIlgQO63IG5HGIOrSzPAZlxxcRkUOEDzROI3WRjN9vgstvQZIT/Qns5hmpDVnD7
Nwin9Fdpjci2h4eCgjkcxJyT9xcgF82PPrrfeQuW3QFoT4sv/DpA8P7kQsxkHVtH
i4wMvYObyCTUDovjwo46Lc43WIQEBH1cL+g+vihNyuwLQzntXXtCkDGFL33kFcm+
WkuF+DECbHD0udYh7ZfwtnjFTwpvZ/U/rYIa5Q0RvKFUnfLZvRxF/K93h8/nQfof
NcvhXz6JGe4w5lsQa97CwLUu/hqRfYruGctaw6xCjQPt8sdUqaWoAWc6pY09/Zu9
oW93CHDCtEGt88Rd3V8Bxpyl9hiHvpBxp+akGIgxXr0ABZi8IQpi/gsYpV2TABQi
4l85E2zipL6NXjZgeAcwxoqq+KvjwUDm/BkUtIfggQ059GwfIDirUpW2A5SVBHwo
gb5PXvu9pHPycCCELawShZ8QWENaLOJwGCqvFzZEfNFiFiW1JD/2CN1PFxcGNpOj
dTFokw5x7UVLMevLMLea+i0rCkjkyEY6t+WCAcd+icye9xe5/+1qjxvOMZ/7/ksJ
zlivPGeaOM52Kh5ymDXNyuaMXNItbGjHaLB7t1dxEGB6MILs/bCIwcrZaV3gOYVF
dcT5oQRNgoIdnWpUGpfuktKemkHdGrxwbY9jVecbd0Sn7iAfhaUYGpzekHLCnyJa
gWuO2gpwY1N5/21rZkdNNznIzpearyJHo830OKT1EMLJC0PDC0+ONRxQUDqLz4j3
YlUwyVa/gPQ4jw+htCwVnMcwiGwCDlfxQc7Xz638JeQXSZu4AINWnRuBvt2rVAK3
widxmQsy6NA/oOsTaVaLqwCU39npmBjmAb2v/ml4QAgtagGarQhLWyNqY+U84C85
lJWC7ZiiDp9ISDtadPqrhHtyA1Jq4HhdflcYdTtJW8dtoqhU72d024LA/bRLgLAe
mO6qtBedlJ80JcCRe6PwBgo9OHpGhmpNXdaLYy10mbiSzVBMLZDmyzHXbr5D5GHM
9imcY9VTLvWVPJn2nGy9oXoQAKzbXPS/pYGl40n7evGgVhL9ykBYM4bKPt3Ei9m3
3A4B5MJHSjj77ixpqrcglGJEXy0xtEjEfwh6Fc1rSLdoRLu2UHX0MGVuI7FntDXA
PBbZd7uTrnGqBY+6nZ0iGRvXSts5zJqzOwX8Bg9GeYFxhp5svhJ5M8K6dlT1WRcP
p8ne214xTXRgjUWMglljBc3z5JG2Ckfi8dT8ciyUv6GcDWt93BfMx7izoAK5BSHq
Hpr717SRSKALqWGpdGzKXKdRCrKKKI8Cc/ZfHoyc1EXm0UTRjDeWT8vwqFj+nBSF
LXvA3R0lkIJc9gMFPDBTDgIAIXZ8ZlsV7+TPRWBQU+mwsbZGO8xcmpJeyf82VMvw
dtz6hjUV1AcEgczHMamgqoxNxGPUX+ve77vYgvJhpzNAqo+xntuQbEZ9RjFOqpw1
a58GLZR0fg0dQ8SVWowmUvebx/9GreeiTRlCZu1zRJhjb1TQuP0op4ILQhV8Dqn6
T4RO0GdbjZRDXLak2k9iQk6Lj0DNz7qObyiXPJinaT1Zji5APi5OYBMy/gl2MNnZ
3RRgAQHVOGM+3ojkqPMgIwvhxSz23vI/npbLx1nN5PdzOu1fAPAH6ivF3s/6quJ6
Ouy8JqsQ0Kke2+x0AqWKq7B4ONZcqHbI8/r2KLiki+RX1s/yLlGABI8hGaEXwA7R
0fKQGuKfbFE2aHi1OpW/7YF5wRISNhxjpmenBkFGxL4IhhrH3OMzBQIaBi6X5x81
1IeWfkh+tQJtaKsCTOMsX8YrOUX+vXv3qZXtvmd5LLKLPwtPCECC7Ux+VtI9c60/
eyUWR4WkVR2/G7FKhAbqorA48e6VPOFdcR5r3C+D12NvwaxZfcp5Wi+ZG1eD3AsY
jXeF5ATdiOLBjq7a3veZKdcnzYrqg56xXA1JaBgGCLk//CCvBaeLUhqn6/kzcUAt
G7fEoDLAy84m9pxrVgxWNFITGK8gJ3oRXEQp1YTPGvMzLPQgMjUYoRRqqa5xTm42
GngXBcy7mAdGgStVXkh36uE/x/h2swzvCLn1lcJG4YNxHinRmDBr/S41/gEl5I2J
QUZME9088mONOKA5EyAtNapGMsw9Mn65dwWHGVTyi9TfCgIp2DOD7c3E1PLSBLmr
tF4D0AuU7prx1GvQ5icxlqy3UTcEVcbaBcl09KmL1YerFeh6NLJgWnel08/CVSmF
ACZQhWa5snu7AGJkj+V6jqo+ll8tADib6fBXXnVpHNm3goazOnAD+odqhullyLXE
k9KVQ0RjbRrhA49Il4wOUh3hzr99vyEs0uqJKEMLpT1wyczgu3ZyN/dXTLA+AFzu
eFaCTDzFRPuEcwI57XAakCtW4Vav696CVIqb8TO8NBfu4EsYOGiDfSFyIIZes5OV
J1YExGdOpm1X/6eHpw3MvaA0ni8EsSA3J+VCdReNtY9rfvdOc9w4zBOIWgTxTK+Y
9MxoJYf1twdB4MQhHxyxQ2Hnz7U4XoPW7t2yvwKGDdT5Z6TNL7yM3cAGTPtSUWEm
sS4C35tQo0KvEUcWLG7x7SWvN0xoUFumTu77KFBmdTBYFEvOeTGbgI+hdjPzqZ8E
UIHPHyXMNDKvhk9EjguEKnlt7IABEKMiSraI76wJkZ5B3dMvz5gzSk7T+durwQqd
Fvv75MTvv0XEaRiQGKgudwJPnwh2y9r+KfmcAdAZKWINDTfQc12E9KhCVBKfu/Pr
Esvy7ofliPOn6+OgVk676PUKp1gFdnuEWPkSLthBicRTBbWwL6HAxfMzTp53HWL/
3M+aq9m54Op4buq7ERLVIlsW0LDZ01I6sQoHx+bN7oF+SNlSQT/G1luL2qWJlKjW
zbLy0dKmQnw8c7CbXvvjKG2t1SRu2QAF+Q2Xog3Q+symLjwyU/PcBmEU/2Su5X8X
cDMUGwtP0hdQNdu3G/Cs1UlRUo0PtATy/yyYZN+LFOIM4Yvtc6Xego79fq3Kq2QB
DQ+2C0nzXk5BexY5j/bM6jZTEwIhLom1Jztaa+4/J3MHsOQuW4EZ1OIXmM7vfokk
5YabsxMbdsVSgS7DW9rSim4fp+daUeMHddJZp2tZHvH5DzSS2Jp6QdOL+W61R1yM
OiVNPFNTnOgAJssLWIAYvAmjwFuXpZgmD669dPU2AGyCRvzukIWCNQrE28PX3+c3
xVeygRYA+5fHIA6aHLa8QZfPtK2Y0fN3/G/yUpSlbn/sN3YdIRkHXoV26gKaJdz1
z1a+Fzk7dBaINn5ULtWIJvA4F1Q8rypfX4wY4RQvazDWinZu5G9sL89pnYRQiUHq
2qNvd16RabqBN2pSpZNX5xaMxOlUTrHG4D3Ic/WCeQE1OGqq+B7doDfXko/uJI7S
sWIvW5T3/P6aMO18Zw/ZyMrgBHTp3rS/tl4U1SkTr8rkZcslqv3uM8IcDfpuFP5H
abBPJbBV0qBEZ3Iqf99bF8KMMVyR5uOnh/uj5+ugsNNPbn76EG8+UJQc5P/EK4wN
GUgv/POLzXJItfrVgrQchLxfF4aeR1bRCmPaU7AVNI21ywKqITjzNbRKIfwOtqa1
DmhpOFn4nWxUZ99iXwacj6eqEnTeL7665T5EuLI6hAI5lzyXLoXIM3nQg36pfRRz
iOKFRUgx4F4LrGLBFWG1oTchAyU5QhAN5ZZjHh+BBG/uj1ddNRUTmEuoriS9vw3t
J6ktDB4Rt+y5tSet8CkC82cCup6+PQfzrDPqb27MNvf4S2apL1bI4gQRJObrdn0w
sZYDReYKHNkF1w3Br6KkNcmBzDxAULpBpRhlC6gUU+E4w/xA4jXPNqejop0GuAfG
DstPQ3yTYKR9OjUeeVIq9lMfqBmFVZlKCNmxQTE10wg0qYE0ywAiADbWjajNcGHc
j44WdPAuHlyAiS2wbp/g1h75xyWEpat6dnUwVeC1JdxZEypemWA5SnisC5oXMXlp
EvC7t9pakrf3oo6gG9eXwKtIeO//LgHw3OrrnOzB0cwToz79ZTviKkvqnbdzZxLh
eEJnD3KvBOqLb/CHvJe2/Q67GXN60P9yNcUXjiugzZON9bdmxEJ62CC16OOy/u/G
U+7/WOlEVTblTmA/2CFvjhVgMiElJ7b27g3czRr9zoK2gZjjAKxyj2UmI02ZFtaK
nR7QCU75gWB9U33SxehEoVhYMto2ZJK+4ctRAoEPeq9zskFszXaYq5ewcWAAcgbu
nS4uzmUR4zeXqsmBB6CZUd40Pxf/y/Ibjt3UwFjv5IBSnP2eAAl5MO2aqCN963s/
qcxj8ZmPzru5e8TSBm+fYygNVYWJvTi4R508SwEeY/b/CUaQBxj2Nx09tqNtQsaf
lhhDrQCQhJIGTa/Xg4VIgwn4YGcCd6zXm+fhuA2+yeAa0+EPNhy9gnIpJg54dAPs
iUWpLx6gk9yAam4/P523xp48VAU1+nJQHEysFDeNGkyYZvnOfj4mVSU0BXqt7s5M
zfM4LwIpJ7nXCKDdoo1X4lRkbUjByJjKvNXBkCVl2TToW7ezeB7SZSyRo0Bnusix
uyeCCDzso2HEixJgt0oSDI5LwTVPfqaH0I/UVTjptTEQ1D96geyGHhxMEDOCLQU0
l3fkb/CChK4BmW5Ubwj+eRXPnmwX7bKxABjanToBh1+F5koB6qRySayDBcrIED3N
WgalY8Z4tvEmP9GLpvAie2uGJjemZTOyj7wAexroeM7oGRDHCHap7eRJ/JuSE+2Y
Nn2e1mr2ja8Dh3OQYfn1SU5AaonrBTCNFCT0TNpOE6fSg7LwoUYGSe34RJ2koQlZ
JeEVHFp1OiBM5W0R0PL4GOjClq48DPDU6RNmT5aCQNfge7WZNd/Wxk0pt78IjnCt
/VtiLKJygylJwkeQdLeuxAHsAlC2GjXerkRDpv7LuaADZROk7XbRj9wLyZLmOxFc
4WnJwQmv4z4fGI9NBldf1nzMoSkrAPdK9GU6D+cmSmtTRaYIu4e3IrEJmkZ/ZIWA
7KRsz5ncpoIscDBsMbedev5gNW07iPpACv2gL7uPF5+Qk2u2F2mqIBkZQ4RQE9J9
E8GVv/DmdfNppzq8i7lFqI4rCBHgBtDkoUcgFpRy5VkCfJWw6E86VgEEVrgYZEgU
MEgA+Kcs0iaY+6lX3IADTPjYhmKXh7nWQGjLuXQsjoDJ+maii4kjEwSSndFMwsHa
Gv6/l52W0dGC77cRRSj1WLS58PMXhwP+FV8o2/H+WV3uVM1hcRwpSxMiND++YWvS
6nnzl+drw/a/xSpA/kf1kvsPJMdnQBzG1XZ0ns/BlzPAoIVN0NN1xezMSIANGOzV
+nhk7+Cxf3NlohJlKiTekDj1caIwYoiAUGrM0LpewQkRkyTiEiDa6L5xGSsqQCR+
iw7R+cbFeo4q/lecSHeJt38aZd5hgGWQ58WSbnkNB01PtDbdsMxmwO5O+BOKim3h
HxtpmuWydMnknMcgzzcTSGZCC/W6eDaVq/GbnKWNlD6gH7CuhMf/uZmwm3xF4B6Y
Yz69lvPAkJbpF1oxla+KlRDNu/z8H4v/y2EAt3KGLzjBponszR2BDfDk0nQXeQkl
mJTxDFjb+vWR6TghRKeRhrn0fxrT5HHBqTqFaFS8Q3l+7GYWkyu8glWoUtKNkMR4
bbsOMLlFPY7O/gZajzX9o3vFEPmRKlOhs/Wvo/MIL5Q6Q24PL7XdTmu+5IcrGzgT
QBpCCjwrm/gqTWLc6Sxv/d19x2+hvlqJRvFyzl1QvjBWcSZo1bldaOoNXZAugyKL
6FsW7oewgNAbiG443V4OtN0qE2JBuHKK3LiVnX84rTIcK8IWxt1Zq2I43NQR95eW
WCPIIewV8m2O8nin39LprxOiVaYnG1dVi8X2r1sZc8iqbx79BAczDIj15csJSo70
ltopR81pRI/9mARyBW6B/n57yssE2oEfvkiCm43ZZJpoFXwa4qkcUToQPWj5n5Jp
9kELEeoJPSzUBkuYFuK6kkme+JxJTk2b6UNPC8YsKpTNbIM+McWswRbihFyaitXI
qK5caiBmkfU2553LlznHaBr5pM+y7x7rWsqmlOjlDagf3R55rzKx5UdSztUbEhDD
n0xGZ7IWfZDFXE+tlLAbp5IjiT/Ibkq6yWjxTbP303wX5PZp3/q6Y750wmKKLYLO
LhbQpoVOcavvOTbFVTaln2RPB0aLtAAmjgyWZWqqxCnxihA8K1VWyIMC6r8FUwe+
GVEtUqvLVfeOMgkR0rx9EuOx6cRP6SCNBiE2+iuEWpY2NHaEuC5D2SbRRuplMDFJ
qmmIeKWcduT81mSfPPzNViW+zeNPcIwCCnbZbedA/XuHXJOcjsH2jzVdfxrOh6s2
jNf7VktfCW+3kD+BzV42+C9qPwcvMSE4Jr5qV/kizJFOL4295Ao4KTG52qPb+28z
ZTlqHktd9I8BLJA7T7MdJFEgBPwWHgk3IGcsWxPzCWyTQu4mNb9UkXT6g9VfUqoV
XW9yxcI4J3ZbsXwNNZgmqVwjhae+fLKLF8xhWj0cobf8QWLOqVecVzyEJ+RMRbDk
Br3bAcRyEIfVYDr8BAqlszszZ19goEE2TLoQ6Wr4pSFSuCMoK1yHl0J+jbdY7a7m
Qd9CIPDQdbar4flqbhRaRxgT+LctiZl0NcG6s3iMAj7ppFSib0MkH2Tqq61c79xO
XgriqZpsQ7YUtYE4Mh7FHwQ73iDitm5gnPDGhrZByxPkwG5/+msJy7UaYhf0gvaP
LY2RZeYmgUnk9ccw0dd2N96Br56sBxAoKf/gl86y+FN81YCImkmpBafzsAb8cwir
c+ZLrh1ec67EBkbnO9S4bDtj7PU0RR5Rws4o5PlqePaqucadA4fTFiaQ0Lz1pXLu
vk0VF8YlnW6t3OgSkPPhh6kluoHGpFGqaP15coMlLlUhdKhfDEPy5mi7jvsHkVQA
S7txv6FjU75OUEaUjqPLwbobhi6kNZ06HUsiEoxjr8Lh+xhd7HKGfgFucXjwFCt1
qCgbLOmjp/dvVh6CrxiP00mvdY+8/APrQ09Gjrk00Gqz0OWshajp/363UV23wprT
NUBZGdx4WgMek8azZh/jHo+3Cdm/1H6/gO3Lp6ewu0CiXp7r9sUSvdJ0Ki7EpR9+
r6ucJy0pH4rUFMwhPbFkrqmfzOhoQgFn/GkSA2VfQyhRxoEOWjUPvSLWqlYY6RlZ
iGl5jKQsU9QvrAnvdCaqZUrNUby8uG1ATaMEDv9ouByM6oDLiwFl7wOzftQBUyQX
B6/A7hZwduwgXNoT9SdKPhBnFguI1bHXRidXTr/FVEZdvBUbKGUy7HlzG4uONkTD
kNKHpMUGRlKWIkcwyNwDw0T3RQeT4DjSInJ5meVWomDguGjIUDP5D2oqDxEx+ACQ
kcZ6BgxEsUbZPfaXHa3vmUp0L+646/fWUSdI+BD26A/MRinfLelbKqOn7uTABfxc
0lWQ0vANsFsYYKWWb9d9Q7XydCTDfDMaBPC8zGDTyxW8mt9KVE2ZwxTYmZ4js7GF
ChLuHB7h3k+3Zb+caJ2E9Xo9I+aSSKEEOiTtgKNRGCczv64JC6nlM6r86wrRblsu
NJnydWi4O3dnKIhzaN0SIzejb7qmcRDw9H9spXSTw9nr51msCTIM2Sg65K4bAp5y
2b6T0QKttcOC+JNRvUoeE3qC/hSf4bL9SqCpffj0vdjibCQ2POgm2iJPh4iaPQk3
Mcl92CM3xwPo082v0kEs3afAfFuL1ANXGemWFFMroMOvyxKpI9SLIcvfv299zytP
N7Fue5xLfk1iqEUMbQENo/rgEMe0zQtdpH+P+uGSU3cV1mdgX4m9eU29yyTeZjpx
fD9IEwpJOCkGpTKiUHdIwMEYK1yKEJRsvkL/rFcRIpsdJxm8Gyz2lfiVS3uu80xl
75QGz9DmnSm3lq3utlnQjXL8tUIWlUNfg6kaCQY0NV9fWsa0g3O3fQWKWgAy3oeD
oLlcAOoyp6OVkCedg1N6ukJCAxIXz4yfjoz+hqgPiEbELWqubqgjA2qG5b2HW8/r
5IasDi1a+QUPp9zBico/gju7VSHDinwputRhtO9BybfCPP5lv3ODLHgqL43iXhu3
BhNtaTqhS/wqOjJHgXWi7BGkwhmoiI1Myo97o03lPERSAIeF7jWfBCW6G7TEMEid
PaYVBG694BsQSVCBPp2KuDEzS47vxDevYuR/wqBC1qyqalnmjWrmF5hiEH0PDrgW
HgUlKixk7Vq5uvWZxVNkoC+2CGNt8nrYYgVkS+KEyQz0c1rsWT5RZmK7IPub6xuR
A+OXputP/g/TWjAUD3qE7xewcxxyRFr0yxNuKKtduLkdh1YJozCJngz/G5hCW1Oj
u2LFIsq+Dpc0Q8i0ZIO5RhjdQlo62DiTmNAFZltgn6gfreLtk8Df18mbYRA6AWOE
iGCKbYWA5evAoOq42pkfQq1xCpN+U6AS2gLAp21vVRaG5AG0QG4e94NaV/3vDF0t
YvHV14RVAfrNqZrtgzGo1Gm7phiJjjx+MUjYfMVF6vACajtYEjEadhK+ccxnhsSm
+z1Yqp9VKnlSw6ytP6yl5+1Lg+ZuNyJCeTFNddf0w1h5T1VEmWOT9mWlrkcU3d4i
TRDYn/WrcwOFAZywBNu0fmjrLGeoT3YLma2K/xem9oVZbv1EuVYdrqmfdUoyuV12
UxedEPYUtcXyR0J2W82cnat9UCdX+RXd+K27xyeW2x1h4gZtQIiWbiq5tvinH7Ur
cEhLT+wr2CgbC14FXeJ4/kBaHNQoZxdoWOk26GW9zwUP4sX3ed/TgZ/6VW3Kw5ta
9mU7yRfbOaFyUyyYRwczD2NNJH72LamXpF8zD3nWdZZPNdZxoSYEy4S3MInEN7vt
1DbRbWqXOHwwsc3XvP1VBuh2ng3haN6H6yhcH1sps1V9vQiX8lGpn3mCcetmKHx6
DCXeDhlkq7td8st6bgeXi12Z3CVqqg5jlZ1JgU/N7udh4Mi3JRe87CkjXDsgD2bM
kBqS+ZYlRcoouOyVX+MAZqUpzCWkNsvTU4z+DNIjspG0VIRcjjApcWfrHI7hkZbP
0O9DSsYhRUgjwsdmrjv/gPcojHeta8f22343b+/NGb9WDJ+M4jK7ha79kKEf3244
hsGasqmZiTI6FQP7BJ8gqeQHsHyw8VXuzu3Wtea8lWFgG4+lpt0KdsKZiGeor4OF
9WYKuWxldLJCSUV7hICjfCaBBeNEBK00PrJD3qxSYjESHaL898PjBRpRg2SxE5uR
YEwVZqfREzWl5n9bCI9qFbdGmyeYad2Y+8dwiGDJFjlE0j959b4h8i+3WbEUlU85
4nPWkJw9zbiLOMRxZKtJMEABoQJvaJ98vw9GdFIzZMOYaa0mTsEjhqUwZ03KGbYd
SttAlLCJI+ZPlaFgDiDQHI/isyrrAmvTRFjV/T/DpwywcfCYNHH6AD8y13szQ6XE
e6QhJ82sUk2/ceCnKnCfNI+DNmvITbKmMW9OvNmuaaF+4aBJ3Ehi5nKWqNx2DoN8
4miJFVPsh5sVUZNX/IUVU9fd1vvaBsLB+hOSt29xcxGdPWWs3m9dxIhOrHiFPv1K
E1lN1TjdSFLRlqXe24aLGYcIGZ+SJoZ0g4tovSRpJ7BZfuYrqSTKGIYtfOM6E2OV
4yTI5sDCYPaWiRuIKlwMv9y3RKSNBOmv+ER4YJmFXShIuxNZz/w3ZsJKMtQ2dScz
nkzh0/QN4clWdPNhabBMHO/rZL1I5xkpuGWUAqrsOoeksQXZxrGbxyHmDIT0UHwr
oRaHZ/DsgOHXkfyDh3l2GAQHYtm6eUGZIfCLsYgBlOnN7n/KamnGOXkFtNkpmFCV
CA16At8wVbI5YfrYC6xYVkP26Rrytun/7bru/fGtnK0MJl2Xqs3l7/lxktUazHQa
f8nskNNeZRopSz+W0HtYlNxFNvp8Pl87w+6PrAonMZuc20pyoRwdem7HnWo8t82B
XEmG+Vr1CD2D+NIqML55229VvnBnSAyrLnoK1AchPfSIBIjZzcLFdqvanAkybpmg
AQ7xlDAVXknJ7UwQKGkoX9vHMYW6zN3aTJzIuQNxVEqdbooRf1u1pux1o4O/5pd2
L9kzit9GOMvoU6CcGF+/NqsfW3CgoUvlkanXSn+iUq3frkwstdO2l6EMVBByjwgm
hBWWfzBaTBSQ/qaOduTUdzcmgGABWQRgCJ9oNjOO65lZZWAdbLDEy4kacsbpT6+t
oVSy7VTYpbcXJ/ZTPNxXEuzzn1sopqpJAFg+zr4vQITGdCPoMu9j3LtmCZhqEJh1
cy4KwO9+P9/8A14pHdnWT5s+1ALxxoTbxq5W/cp4HSVPcX0PJZZ6dyOdQ2hMcTMp
XwUzU1Yidb5uTlwhmkvq80jfH3IXel6JhFpSFy5CjZFSqNs5WZ0HSW2TDZox+VQN
A24oADXB9vwzk2oH09QOETa33AtloPnJCHU6bVpjMxjo2bMiGCIIV8e6DZv7Wjk2
JeS6uFF30YqvO0pzVHKQvxuTuIXm2hyJnHKLvdwNlVFq9v8CY49yAbnF6ixorjnv
pgmB8QrlduVj7o1Gtt4vWbNWyml17mRmcSRpXt2cQiBk7Hn+j+5Kx1s2zL6glc5Q
UO/SuzqSfxHa3tgy+yGa0xXndz4UoOvDxePxr7hTlNpAofAYOJ7ZBIZM81AN2Oal
Qd8iB69Nynu/cBf32/atLOJ8MSU6ZP33FAdVFbY/n0cOPv1Ns6TIV5uTikLhfFWx
LH2VC6Ep/Gj/b9zAMKpItn5eX6gVKN8nfQZJtMhALRyME4xCD743A75umahvaXti
ZU22p78UK1QJGOEgIcESLFNVO1+07mGKGdi1kJymO67LoMBjZLKO9WEofdqykD31
YXVpBXMaQ0DEKHkSIxtp+VmAClwYfHoyWzOpO74cfRjo5e+ELcS5K0E+x8m/NeZp
nbneuoDIN1f/5DQOOHIxw23ulPCDeRwh/8afzPb1E0Sd8/YbN8ADg4W/ChxAIIBc
72AjzhRw7VCMBQiz6WTFvKjmuzcF7VfMjuzbayokKasXe0yPXnqUqr5D2nH/oOn8
RQwd/8u53Bz0mzdHISdAapzHoR+INekKdHDvgLUDcq9c8My5tWT4gGJfQ5J+4I0Y
jeXnFpAmfU5zaw8iZ5YdYRDT3vyR+hDxutSAIYlibZNUS4xlD809BWFGx0NfY+RA
nyuiegA+vV4IrXn4BszJ08e4MFwJa4BsAkne4LEzY/d51SUtwtNqUGhdyCW0ZLw7
KwrUsboqFm6gtgSpsRXyVd2byt9AO4D8N+bouTRTN5uFnLCUKmcP9kdvzh7vSymu
cgfxP+UcfXgNxvr+IWWtbEjjiGV/F8alSXn7bD8NQ0aClbjJJ1tyUOrjUY0Hc0kv
HoEdZEyjAZciJaITVyeHj4fmhHJtURgFEXTOgPfY4pZA6QmXs/2MsxX1IRdECYt7
O9aqlaVWRM03Le8vnWBxnHkLA48H6uSeJtjaykYZyzP9IuBuyYg2cKERID23EGbW
RGNR/DBqbbJjysFxaxK8DCeBoIknDJJD7Oq4V42xB+Yngxvo7fWrkVg9Z0lLPwsK
chE7mnLadVoYM0Wdu6J6T4Pu3poUoAcy5LBMPgZkYQ9Vcj/JOlmcp10okzXvnhr+
sVttQgeiG3Q7UBNVLJ+7Lgpi8ZkEC/Ruo2pPPGZvlWJC8x0k4CRRJF8JB1ALEdH3
QI+Mr2pQJ0b+/unao2b/i2RIF2NDL8sMH8PJzMpNKl+NjlNY65+FLH3pBFq36Yry
sK3Ee9Cw1LGgE9sp+YskyqSpDdoKJuBR8ksKvflWQMgA5z6cxpQ1smxFiVyQdVLc
4jKNB3MKHpSvJJzdJsWshHSs/GgnlAZWirUNL45c8wPOx1RZwTOObdOy02/A7WEz
GhmrCNzcWQ+/ujtIcw7nyvHXVL4HeO3weSHm97LzEXW5gAjA4hvPodUkHnyQLwcJ
qIePUHzfGepGT+cbhL/ziVTrUrKmP2sUrisX2qnZuvGgHjoPljxIxOoDz4rj0yMc
eeZ/KzV6JBPL9MbQqiX+KMA/VCk4V/Ct9Maj+qsHrmuPkawKfLNL2c3Jly+WD5gg
I6ibIZ4gGyXpg4XBNQ8sw7xN9V0D2yos7+GG6Y57ldaoenzBNoJeZJ02MDHBARwa
rJzMAtHj3EuAVafSmzJ0G7bBcfNVaJiKb+IF8MpCLnzLmKaC6cpVGtgwCkiOvbcL
pb0Ej454aUSjD89q5siENJjFiQ9sB3e70XoloY05i09s5HSkIB+vX/fCFPZWvCZ2
37aB2d+ddnGsQMxPge24nU6urMwvz7JyUzCgCCBAOG5YSH6HaI5ifWtc3Jpbk/Lt
wrlb5Yl3csFpBilrLBwCmrEm4DNjLYODrtDogD6Q+QPgtaxBiOf3/UT8aIFnNiXx
jyCk8ym3Wer0XpnleY/HGef4U5kaFjgcYF7YyR0jFu5FrcVNm91UlZaKyeI5QrIq
sgecAPX4dZJW8Scc27P6iIOsv6Wnal1Ytj8jMK/BgUJirHSwFQQeWr54GV0su/M8
RXv0+gE+IMTAad9fNLvVnTRXB34C/fWpQtYdOJTiWW3NPp60aV6MzbQZCD9xjvJN
qQq63A5OHIWjuZIx6jBNlyLpWlsHWHe2fGYOpKZlsLiyqQAh6QPylHSHS0mRRHJQ
K2VmdlyB4dpfQjlr10eGSed9949juxo4UxiaMjLJBKJ+T8ZRV4Nn2d684TBubAv5
8KXyzotyUQhC9sTkD4yGRUb8JDRZ+hrgvMiKWAcrw8/j6kZ/2iaCBtwtaHpq3WxK
sQshWn6VwVlSrfL8B+fIxAKRnEud/aPWEAj0QeSMFGutpquYAG/9yQgXDFd1ddQq
jTCI//G0JZyMVR2EwhKdVA+o2R5ynTzCpOqM54jM0PTNcEGvpVioqne6KbHwvm6Y
QN01cE3QJZpUbBA8axdzPH2YiMPCBo2d0AjZu4Xngi3BJ+OWavapJcmK0hvrQZ5Y
YnsoRi8p/wS7JQukvbLmt5NveMUvlon3ajOD5uLF068PVHWzZg/HINX8e6yr90a/
QBFDF6uVxXS49HvVN8Kn9qErDzqFcagulgldYRGBH6/5lGdg8P2rmtuw1SwWpluJ
RtFCg5muNbHPH7pl3YnlZ/Sdls0+8I6RFO8zd+ni/heQ+7KHU7fzZCEwOHnCvvFw
g4zT9aK7nIYRM1yv5TnnAG+K38cKIadwaTfJF3fW3aTKUGOQ6G9MGQCAssNvX23G
WeReKmrjJS3aOF030jhZNXAKamHzovrJYXD8bOyhwLgyWocwO9Ymll5nJ8SrpCpR
ARV2s6qVWj0HScQG53FwgrjQJ8p2gtvmAgCAIlX8Xrk/oa/BK2rBNwlY4iYw/EVw
zoZ7sHlaScST7KdIuXLY3Len+fT0cHrMT4aLiGRWaafowp17oX2zXE2y2FTQDVwG
59n7rEDx/rKKw19PE5JJfH3i/L2vvuY7jXjlNgm51HfuB6tUAYOloODpowOw4SsF
fNTBxF7eTfOaolCWKVb7cP0B65+a3QJEicqUt1zQYl7kK70pwnduZaU9p10ycsO2
OPlWAJrW/beX3NWN9thfhxXRD8RW2jBR/ssC19uhqgxn0KQUoCuE5oHgAcd4DdgN
1uocnB9lddrLcIpGOZhVHkBWllgcn5SufhMJN+gScZWR3GgCan3dPuGFOzfjnBW1
L7UWWvESm9ag6ZxWhUdo3mJB8rBUMfxhkmgFssvIhVXSzoIA9PoL6+OOxo1aG/H7
RO2Ik2Q3lMn0jAlfVJ/UkDoHiI0EtSQuY4xdurdUXTNxJIT/Em6jImKUbc7W10PZ
ZWaEHFkjOamD4rr2KHIyaBIF7Ate1dtkTeGucHFK5pbA95scgRHL26l/w3bDLrdr
HkYeyANIXqvzqAENUdGrmoJ6C8H4z46id0ql1i+FV+YWI2bdN6ARpmBWF6bVtZba
1JHuJ5Jczzh1xql8WMo8KiS8oZJPY1eMPeEGq01RAZRCf1BJ7HB5283K+MmSV6Vh
UuYEPdf89HRhCyM6wl2D0ZvZtwWQyMd8I7WrXjt0MOnGtCJ/fF1pNXqh180imfaM
fs9dt7VYCpbg2ZaCEKSVApTSoZjuifqS/giY6YbyFZAeRgYg3Od0TfjHE53ctsON
htKtdqn0FUIgv/B9R50bMMAGKXaRoYj90eDgP3kWFgEc1WeyJ7qNKhjSCdtcpMQa
GpTfChE8X8my0oJSC5m+/HzpFSZQa6CI/FgldreV1nArNGavu4pXDHYu7wkPRvJc
R+WcalTU94QxYXtz4DhSQz/kEN5pTVrCaMbNLE16AdbRGvdXuyjzM7te0jgTsprf
wllFmbqrL36RWqA5vmF1f4OXgOd9bToDo15L9gzUaYBQvCIU1P9aMmdfBi7WrJ/M
SrMTRFnnE1IZuedCkyjXOcji6IYC6j5WoIbKHoW6+2YvnRaKjqtAyDSz/oYKsNQ4
TsWYZWlqmn9sLJVT0dDrNq83zbi/m7EDKJJmbBjKbxI+8NbaolF+sE7SVb8IoXwF
E2ibQT9Ic3GpxJRbAaPJM5EzTjh6Hn2Pmm/yMJwWNM+LKL2kEU4jbbjtIf1UQ3Mi
f43i6LETstWzkwTS1BF/YFqPIV7T2NT1fGteZQ/16L96GQcf96uVJo26dczdfWOu
h/sr+MJidCOgizOjCKIGxyhR38njjTTwF/xrTmHQ7f19drkdTN85r6Tnu8poBKOt
BueXSHIQMYHRm0IW50Kj9/c5ExBwl2p/e7+oq3bCYJnuD5I+/qWni1uxZbrYXKpv
yIgicjHNFIyW1sQ5PEywktI/og3/6ac4KvUQTUCble6fYhx4mP+uK6Nk4V3+8oIq
Q3dGVKbZZzy8ImA1KLXm5MUVcXTgnvObG0zYcn4aXds6OooPNuDyp/lFlC8s7hI0
fOvuFCt4TdPN9ILmcTsEUYfgil+933qZ+yS9Nt+uKMjJPHyJ0tMAox3gKmUiipwh
0WJGZ01ouxWPZhYw/i1a5YGr7ABRnJBDg5y6rx6/05fedq6Vb6/ZE4/d+lbCQOH3
Yh8gfZ2+TyYdimX541AJWZS0BrwF4fwJ3tRqewbOjyJKEAt/ygTJtYjwyrPjwWQh
c9UpCGVeB6Zr9yHOuwKAV5V/EZguhS51TZOGStRb7j8yLz1MdeYZIviAOenbKx2A
F55Hp8GBi82THxOmE/3tPh4TBjzliwYSzWggjX1ThaD3ukD8kRoXJm1u60RC9HhX
UaJa1sLaT9EYEOVg1Z/q1OsuhK2pR/O5uvrYVHNTUYtXVN2TJHvpEJAjYpWpdsA4
b1pSDFe6/yLhQCBV0lCnyQY8hx3iF9pcynHTzU8f6Cm3lN3KZDlxXkSvzsw9I1k4
jyS5ngL9a8PkoTMMMib8dkybjdlXe2W4iOhpFqee/0PBbORO7tHCtfmTV6WB1BML
r7DElcVORj2giauizkWC3W20VjvPbuVPmDGttWMVup/Dp80wr55ukTqyZFPFXQ/B
P28bfMcJSIB3pVCnCdM2DBYnXxvCmPL8IKvFtOVgucPojUGFaxadRaYFD+Vo2UTZ
Vrb6AHvRZZRG4qrEMeo+aj2ZxokP49rUZ9MfpphRy9RXxTJ8P+stEPxxPlekKAwm
PqUeSyHwUpFs+CczYghJv0Fyhar7J9poH40DNy/2Ju/7z9EPKFfH0W+GS2lhkaLw
CmsUdE2TshOdNow9rcLl2UrDXvK9qPegKffbHCd845iarywWh31Hr9vZkBZtU2TH
7gEYbiSEWJyNl0zXwYyhIt5vOH77SXxKTWi6pkfN8ote9lcPJF8O8bjzQrY1aZsa
OzP8BYgEigET5t+k9uTE8tWJhyHwQK/qmNCkayfleAF6W9mn/croutqIQpKlqPBx
QDK4hknq61V+9GjSgLpJDYj/NFVDB9CNLe5SSxQwLDT+RgvRiIqFj91KCfOzvxGP
WGtqrqA8d5BHmdMor3xh0yZv1IS41IG7Q0VrZi+GFTReAvLo4EjqgyAyfqdgaXvQ
XzcILVO+LLEKSiePcvwgCEhgEOEtx9yMEk7YI8frkRia8KJpsSd/HJ0Tnclyjg0u
z673OsrBo8x/mvYg8oi3dOWrw7agFiOGsZWrAlSPU0+0/TWp2wG8nT8JK+YRo0GG
qQ1z+/AfMTGoQoGlOGUjqtaKfnbpOgsqu7yHtrWekkSKTZirJ2RT8vm0rC6//h+9
b+7ktrm1j0yF2zHbeJ48IjkX/4V4DbD+HwJyhMB6DD8z1+QXaSnjH7le6g07IeBO
w6yHD/SOXO8A1pxZqPtfChRfEq1Hy3jUuUszu4ZTA1Zdmtu05VY/Wbab8oYh9e/T
2wpBp6i2JzHUuf+x6AacfqdsbZxkytuyo6GXTqsG7uCvLFCYY3qGthozHf87PANB
zY/DPr5f1LnrtmlLXHAk5uD6m23R9qaxTfOWO7HeeuWlk/LNE5mBdOnl9g5PQYYq
fp3bmZxDY2mcQ0dHuvD5zVtrR++M2DqElL3xlBay2CEXKI4R4O0jRF/hEsYikr2g
jZ/hdX7m1N0m/h5EBhFSargNLCtXVmNCvKYql03XST1RSg2lvh734YL9Q0eLrdZ4
VHdxNjscO6YKMD9eD9v/GFraI+uXga9Gq3JITRqvgmyxNtm+PEjxtTnzRngqp1Nl
wEgLWyLLOL40tmmPxQ9ff0txO/snOQ8BbUAQGLr4xVlSk4qFk03N9G/nJH+XzJdK
5vKkJSpqexOOgS6uSkhplsDUYsUr/Yld1Ew0SOIWa6/UWzHG+/jqo/u+oSvNxYNZ
DEISLLRpOEA5tvHqYR++pALBir0t9K4omPb0ddtYrGnCpNqgJbXsW6xvakIWS4A0
0kWpDANJdkpjYX/4z8oBnQvz4ZQ6sL0t7gI8P5cT/XcOIpg7LyfSgLlJKgzGyNWn
buNDjkWKQsbED+0SuG36QOj42uCCBkhezY7NB5O2PM1qr8B2LZOZKXDUI0l6jg55
C4wQeDh+jccyQfitAhPrzIX8BnV+V42CSPI8+UA10y/DCmZbN0D29YfK3ynEcuJQ
K6Tv3kPtgZ5Vwca9Oh/qb8URzVSBaY/eYmrasXPXw98XoaVUfNljXFRZHjL6DkBb
Mq4Z37bkll5GYZ05QyBeIkmylZSBtHJ552/2YyVttEtaP4fGSsjNausnYEN4fviZ
H8IEtemrOKQrmWemswFTmJB3vlcLut5XmbIjPYeHXk84ANzd7s2t3tmdYDzE7YUy
UpegnN79KdPJ5ae7UKRe0XBWh2U9UEqjmT0yMw+k06iUpDSGewN5Y2uDI9JZr++u
MFXmTmWAan1smnro+RZcLRoEqWGGTEk/1Nw24PmpbJd0r1+H2JGux58Fe5ou7eFf
2tVmQ6CISnjQujoKGoblgg3q7zy/2vtzrldqSSUAFIDBZ728h8wQ200AB9t7eSo6
jBUmIihYTS/8nrKn/6fSSGiMjXJ8XZ55dGoZvB7JuQWboPP8GKWfQXy1bhN/P6++
c5InKshECqXWkKgHIa6Owjz6MstoZkgN+mo9NSihQ1/wl8FmrKF0p8tRy8BgjaRS
fA8Fh3pkT9K01QASNrcMVHuf9/GRZgNEoIsnd/Y+/quGxj1s5a4M+GukTbdKO6l0
a7hHyLg+hzyl1E8SHYRW3t1CULgET65rfcBHIeQJteWuau/QOCV7e5ZYMDlikbJ5
PuC6e3ntAssdCzi9XNrKok32+d2rn6+blMHsg3I+vhDmPgkjC1NwORY7xYMzExd9
5iehDy8D1mOeTY52S+KDGZt7qDVgYJ8kP3LM9UDsjOocwDs1mKLFnhLuOjvbuFQ+
y6lsrA8PakDmu0TfEwyJ72WB6gUxy42SDVJpigkTcbZOIQePa8R1/wYPmMj/+qhm
ZJVWmXqHNBqs0dxSziX2b3cOE5+ZCu7MYt8DOmTspirOPkRvhJPuOjp1xE6it61B
PLcIT4eWo/6sMjQ5vQj6dsv0/E7+pZLoDg0MuxHQ5cU+wIzpyAseS870yZyAWEsN
IsC8VZclyKe+/95YsR44nP+3B9pMfZDTvEuMXn+91QPk2owVjEt9VeFBqlhGBI/c
N+SmXlPh/bNnMYkS4BoJa5nJo5/ABAqoROXhSq+hk4IWT+VfReJI4fo8Ei8YXhBs
xNtLBWGUWMBTxyN3qc32mouc6+YFu3SkOPYwRRmUbqQWZEHChntOFyt7cKlIKa2J
/MiVd4boVIi2KHnSuy3tne3bTF+v85MZ2g+N6gQlOV7dX1K+R+I8sON2M6XP3XNj
EzT1IxQiGj0Qu2Xe8R69/i3zalZwJAOhT23X35ZgHElVOaU5abm7hcXhJFv0FxoC
guwZjlG80S/TZfyj969Sc03DOLpJ7Im3fT0Tg3Qm+bNybG7JrlxnfYtezEGrKM6x
EXebzLaFLs/9ZZJrYikvHN4pD/U5ZpH2uZaOw5jnIWQ9hUljMM/JbmRX1ETciULU
IswiiIZjLFfor43/uc7QS8qrdQfQP1HCKTie74PkkOAKaSPPIpkBF/1b43yj4eSd
JF9mJl51cJG24Mx+ZUbcZavQa9qh6kZ2/sJZkiK//hQTIgpn8F72oeU2aaAWol8a
0b4pF6yle3cTtdVYVHcyjQ4FTaLLbaiWSXhNX+hV/6eGEmMJwA8Fz0dj88ayCGLx
GNfj5C8L0o8oAcsunWxKQ+R9p49/s0JF9yZsQ6s8mozHMuNH03nHapjKp7xlx7Wd
Z2ruRe7cAgZBr0hzpl99naEBfW2CLCGramnxVEH4BiGaETQ/zrpV5fDUluKlpcFC
wKICt58LZWsi9SJmhZFDVfXR6APXT/dmB7OSpnWeOG8AK5+QuBtOeKGOD4JSLlk7
NyojUPhb1sMgxqX2qg9p8ES491JP+YXYgqV9Eq85Jh/vRzLeJZ9NAanqDpDgiZlk
oay+Mbpb8IL+ehuoYK0EvNAopU/O+gaeb7cJe0bG1kCum0nOzxzARvGCQCwLsLwx
cU9OLqhsQoiICALMid/wiAGWYfueAnnTr0LF2eiakWTJRJwLurLZQ5SKdE4xsqqc
OfnTaYBGts3wKyozbxDq6pmxGzo2puPZ3OveG5s5LOVehhR2Tkc1QkVQ4GqtH6XQ
fjdnsyhEMc6k9ezmqUkUJspwOWJhn9pPGKtOFdyZz87hmsdHOdG8nd/3Y/a9QrNQ
pEev0KQQo9krsOLF3awiBK0h7FTaTv38I4DEsRoQn6h96j4569eN4QaxhZhDsd6V
cdDYWHMeKwBF2kA23MJp8UllAqc02hlXMv6BlVBfmKbdsLlQl/QgeHVv3aYWPSqC
2FZiqAw8E2je4AK4a4upphkMoDnto6D3dPxtKNGVGiBoKz0I0CkcrrcFaCLd4B6j
prUEFLon03YsNG6OB2Z5nGcaubB7PR8xWz8lsmEKVEOEOaorAfMyrdTmdnNQ/NEI
6mY2n5WdUIYOQ2qBDlHitWCzAUun8Ck0Y/PM6p9saf+0CV6V7KVGFXnJGaF0Sm85
bOU/QJ1/1xZg5wNE6swIuYmIBVoPIuBiy2MZe78DkxCTmFvA5rHUkX+GlKH0pVEn
Jd8gi9Ct1Q9hlPv1l/gFlW0AnIeddj8HJYGAPmB/irn7JnBStAglp+7p/3tCk45V
LpKShmZznGncbokNqWFkXBwINNiUBChPGjOxIVtDiqaWuXWq56N6c3/vvAiXjTN7
lGlMwYeB5LCta60TdUJrYf56q6XCbYR5QjwE7vsEIz0gmus6zPSuAHP0Zwsz0Ncu
PJVljg9WYZzEiXmQRA/OKUQu87WJf3AxmAn308t6hBZWpmkxZzMJeqQGqw9F1FrI
Wa2EamCT+80EV5QoY8AyLBfBibGEZmp8z0/k/AeDsI5fLFUmN1SGHMsTGCk2r/qy
2bE4QFUd3kmRcovaftGGAk4mOM2wAXpQwD/KnxyMPxg0Ep8fu1fk5crYiGIKApZ8
f2il042szmfpYB2GXjOuNayDxyc6zOmwPKiGStmW7oJ27bX/lRrzboKfLb+8JRLE
e1C256KlHxBxtKx6LvYodUhKkXampJagka8avuVRyb/tyP+UR9+qzFFdixbtMPNT
CvJJKzHga4wmKKcrCEDGmu9MWF/nNvn1IYlnKPKAqlrcRoIJyTW1np5I6scM+zMX
K4CWiCJvSbi3RzCJDuoD+Jl2OwnJD/CnqAv+YSJJhqxhgnAmBi5w00HP1w+sSqsV
R8SZjgyDjuHDFKcBb+HDr2z2/swDve+O/DLgiCRGpUcjWhNvurIqtEkE16BWRYcG
CQB6jje7kpXnISzGZaSEb03SCoax+o8kOvF57Qj5CfPXrbwQej6nViXqtjaA15yW
TC9cTWYS+/Fy3NNjkjRDZ5fY0lpV3ExhlYxUQlBytKMaevxQF7a5J5OT8HCY4DC3
COgq0AAA2kw7l1oLMlsPEH8/TdxJy9WMtxKDe+ooFgQN7U1z41X0OwQzHcEZL3dp
Gw4i/MglGds/dio53l3v7BRcNZX4Fq/XifHrZQ4b8whKFrlZOUykC7jH75fuIGqf
fS4iGfr2ijPJPUt6brXQYoniNrFOzKvz5ndTkQb5zLTgoMAYou/tolj7RVVHwByx
ini+9J4ph/0fDUfuEPpC7CzGMNM7pzbt9mbWoyABH2dLsHpi59DOms7+dckaNb2a
1+vHdn3e+0oe5ENouizxo+eIJv0Ciyf1ZoN3aiUYHvi8SXZNlj1dBYs9eU5BaQ6w
yVbT8KjEGu+ZIQc7Dq9IXlhf8xc3ct5YV5vOURu49ahOlD6/Oayhx0UaHAcyaWz+
w905n6gY3AeRIQtXKuYYqvYMav+Y3NEmrVmPg92baSqkY3nG5tD2spIwdjXSx6Mv
BkWV1VbfbJlCC5SlMrD+PXlJEBB4r6Mn3LuI6Ajm3OsXFTrOInNu4esQCiit85Pg
yiZ82oofQFF9+LK9/uqEaZUT3kluweKhPBCggvMzws+ip0ahe1uXpYYzcIa24R8H
UEc/0ertgqfmQVldNg3WwfybRQSAWH7AE5ucMxT8eFocoeFq9SAKFrzUyJqM9U3O
VRdouznkR4+cVe3iKA7y3QulC0JbdwOF+rWdOAT4k/RhDEAp+ZCBRvIohMiQTUnp
imotXowLr7tu8opmwSiE0KisK7EL/cChrn6s6NPITgv41ec3HMOIuq7j83m6Gk/6
qdUgG7z0yYSK0/AyNSpHLcMZbVFnafYeeGUYmQuNtSGVKz2m4q/wi7oL9AfLHQjn
4wH0HNI858CIEeRExvatR744MlCRWYqfHpeqmuMovDas3iUoCfZSB8UuSxWIilGG
o2jd900bNCKzy/C24+UQuYRxnZrShCWOJhrUnxWd1Ba2KCvwxybpoL48eJqg7gyE
xDyRWrriOUYDucwhA7EhTPphMlkGjJ65sphyAFsjRgZtzdPNO8Nk+DbfWPV/5Qpl
nE6jnW9mwIoAMOixy2GJgTNMp58fq0wGvzO0qUbgNIiCZChFy8e50syJ1pKDjBNR
XMPFhuCsDCwU0IDnU6w5NmRjEtFKlPQD7kPXLLU9UZG06l5Cd07rZsy6X91AEPUi
UfnRwIoTpJR2B/ZlEXAIbsD1bR86ZNqpInOin6zw7m0b3dUIcmvd41qXGkGb8MJA
iZnA1CPwrDcOVpjAw2FVQoG5PRWJJnFPre8gDGKeneTe49/aZ7NKKlBHx120p4vV
+T1aXJj+vbcZRNpePNMYHJKs4E/+dedunKoyYz0EnBAg3rEoifTpM1JsFQy1rZPg
guBqkhzDb18tjxReJJegJRM97n4ehpSNwVpvHPAJ9P/gLjUto9v64JRx2lit6A2s
C/S8zWdCLyAX4hAJHes7pfWK644Y6Zlhfeg9eRJ5esfuMesrWJY0jyRUophSV46+
dUTi22jPwDPAVj2kNuIqzzHBlCN4RJeLavE/A6ASs2ilGW38Qglb/KZD78ToIStG
vpAalykhVG0C0kxZ7yj98p0gHap3eML5DV3Ek6OcNiTBjuny5XxYFoKODmf73SZQ
Tp9rW75Y3GNltJLu7tS8NJSJ5WAGCXx4XwFo+MDteOnywic0Tiy+IpDZ1A4Pc0hY
OQX5MrB7TwlI8n6J4e6vTV+xU3JBnV1NYrPwqYGVg6jq5DLW5y4PnseFFheHRjCQ
tKFe+//dTcUzm+UXflP/+OXv0a/ii1NrsC7h/RZBshvsKkz/mhUG1EsTgCZOO57Q
fTQxmus0ehQbyYccv9iAy6tnB8KxIS0bagHmuEqmqb6fld+egJbnLOTcz5GapdT/
pduvu2YXF24OWm52679JMY52+JHKBl6L+5i31mq8veJXYg1IYUrQHFlQ/37/AyZs
M7xLsir3tS+AYp9h7vvObT1SrmYwBCTCgb8uYH2JeB0BP7MAmm0WhTCpNR1qpYim
9GhIt/M1ojUevPbJv9P2OKqHqEWh05rwC0Xk94JDfXlv4PzIWb4RTM+IKOjo0DhA
cedwOgvR2reLWPqPLqX+1hG0nS/T/M+G32/69UzzoTr5KiMwcx+n82P1J0RsDByY
KRqNXQcw/4BeVsjlYTK1ud19Tl4LSNDUkBkqxpYDztx24oVxNjaFswIsPU3dgvwr
6Sbo3fendRoLeb+ajd3KzbDT1EBcBcT2Zcge6iNQiejNdpWZOjz3hCfF7oiqpQWq
KRcB3suYFbdcN41/P8EPNS6uWJsNnTu69nZSt5GBpVhuREqhBANLsuxiSI9vXMNP
MZs88yE7RJ6U9RjXHbl6PPq9yWJeKwi6oSCaKY+Y81SrsB3NJfYj2HBEleeaQzdY
G6aunAMiahRY1Jb90/Bp0dTKYp5dA7TmAie1meTebtM/vFF9vi6Mk9es07mOnV4R
wvPn8v87rJacBSbdCpf+pVCwwkDWCcq6PrA1z+diXekN1TPsFSv2xDBVXdkfubVd
FfSVr5M6ekayXmVv+hGzupHlYI7z2K6ZVHEfaX4krF6QPwSPALLRDn+zU+62bT0d
4EuhuccoCJnGh9LbFTgtR98vmEqdn6fGVFPx/29fKM0eCJtC2DLQwx0TBjdLhoCj
O7Zaq+VUj7byze9iExRGowNh6fuUQi559HmVVDPE5OAufPQxVC4Xyfg+sxL9vK5G
4xNrelxO1oKCvb5wN7qT/r42zqOtc5ctYyeRgKPpmFrnj5JnAlKCVA6YoPzD+Hlk
z5vJc4XQLkBEy0C6Ir416W3g+W1IU3m0AyuYUecx3ZldGFKp6ClSUq2DfEQoqNkt
4MrZO1/3UeSvQCoqXT5gYg6DSoz6Ntplxv2yMU/tLHQ6eJC3m9FDf4q9aeNIV/Sg
mZY3Z8OHAko5ILCNdRT+7cNpUnD1PKN7a+KcMbkASqe2pms0XfmadB6+CxB12X27
Ql6mH6LKnlilhbS+FsJQw1aG7l0qc/TUh4Kt7x8VMmRkz0gwpi7I3IShBeZ+7yQM
9M1EnAi/iBcW8DUbLH9xGIR7Dt5O6cRNWwGgrIoCASHsFOUnd2uaVo4mWbxSt+8Y
JnkR1y1uknR2mxp86+L0OitpqWdsQijhqVXs1HMFI3nOKZ0ilrCg+kzfbPZlg/LZ
Dl/yMV3EmD+DSm6jw1nJ5yFpO8peppfWsyxF4PVOXliXd+euhNQyrqUaL4xw3V4m
kBztEjReXV+5GGAuFedmWvzrUZEgjgcfdZRVDt/SFWdML2c0goVv4NavDci/826y
ic5SkDYDpThUkJz6SGv8y5/cKdmXWOWMr+IukTDAYcLe8rI64BR2gb75BtbvZc8S
4ySiZxyOWj1F+QNKzYBzENFW46VGWEJNYnYhyOF4lonOXTBnl8abwmnNxEumcpgb
mnb9Tv8PAWX0in/C/AR64z9nD7UqlmmVuYRJogafw6YJM9JQ3xckxCjrOGijejX/
+yMNfqqTtjTNAFlvK7sy0wURqWCwISRzS1+E/CB7vR676IBYTVieN6ddEkrqVitY
+rjhj4M2Ff3TlIearFUkYIN4nx9Ugq49c15n5DsZqASMxzOhQC4blQ9WstGeYLwz
TofW+uG63orWkgoIDQt0vY+MT+Ov28flW9SLU6XjaWsqHFvP7tiTWb9JLDfdFQyb
LhCtLh3ziAa7OTJP9lGOAsT7D5kPDBbpqK2jgI4KOMXB/P00qKG/I8r4lhn1azuE
A39AW7vPTb3diwrb/YqyCgmru9k4GZ3dW13UiAhwIQu70o65Ur95qKeF7dblB7Cz
rmEc5YWOSw42WCHf8mvSwvB0+mF7piSLAVnjWVbtP2OQQFSPrMWAXroSZec61t6G
Ar9SENZ0oOA8gZhto+NWLqiI60htHpNzGCQ9x9U8DDhGrmfZA4RuPm7z0nmCiXCO
GW0Y/1f6XzTlonbVsuEe77Fk73LgYlpsXpM0ONG/+7lOyecy3jdM3Q/pJqRye/Jy
QjdtOiOlpXEr2cyrpNqcnWbn1Mv1sB5VK4zj/2zkhOyVRoE/xKOAWfR0txkcCG7D
2zE8k1W/LGPBrEp7rQ4y8laRCqINjqhVZK3sfWbhIVsfdhdZjSGE8/KhnNYXEeH0
7htWll+iLhLWfCV2bvgMaKUGZCDQ8deL7fQsWPU3Sm9iL8df9J96fHsccfP/YfdK
KGU4vlnN2s8ArrmMf+5uwVkImsXtyMxPDVC6FN04rx2RP2ej+sq5rXjpkUlizXxg
uD8Eia6DMP2/EOgzDmyOCTLrjBfRIh4zSX6dfmoJpSN7HcfHBc2o6DrhggfnGY75
tKuIr+tdwbu0ckcwkFTV8VqRi1wuZQF/GGY1Vu6VwNL6jTYkNwLMirLWxW2gdu6K
BvyhWVsNz0utSy3O/nZ87Y5VBYpoVGPTQuOkMNZgjATPHpz7snkFRr6YrhqZgEfz
elA3xfMHaA9mNjq1Iw8vl5anIja2qOHja7sqr1wFRaFRya6NwpilYyG8h88yYnZl
xhIO+SEEWJ6JRhlXiBnnz8oU0DuVjGqH0I6latIbptew4egkVR7DYmqU0GYnQsCR
eSE6rXwSByYPPrsF9NTBW9JaGZEdw9LwRFxUVlZCONmqPsZ/0MwFR6QvSAm9iabj
xo89U4j3tks58fFoaR9eE7TAX+OBMBtJkRGUt8D/S2Bkjb9aXGO7RL11iAJWrTiG
mO0tlW1X0UnD+KuTQZzuSnDDcd0lEMpUpMLLA2bNcko0Hohn1ruEaj2spdRzyey5
r90/GMS8VCvaPUsU0XIPk2faok9sy5qjoFUhbNnBn2AI8PDnIuy2448+NV5stzIl
206o2aH1eDrlij9NZjwiaqEyT7nHaJreYSvwoyp+tt3C51X8TXOnahsOeAFiB0BY
+QlDCWzfkY8cgkYJPU3pV6V096viMyA1wa2V1fAdT/iNUhHqzH11aYOBHMtU8tcH
BkCVEbey8ARbX2YOcm0TFSzxh4zyO/KzgQy0xleopArCKoSJFT3TpHIVT76J1yt5
YMLhDx7MY6OlD2UJShHt6vDvGpugWGqua/nrKFwUaUpp/Xk5KlPYnb3PzF73VqqE
m0gV7fOQ70gtvuryFO2wZVqJjfzwixyTh3sbw5tHyjJ9Z02vOCG6gLuG0EkWkO0/
K1Zmid4XfnygD4JEwZPfuDw3HRj/jmFD75o9EujfF2IvqrMPDOviNic1ga9dCQ/4
s8ylsQzJx9MzbFHNk3t/KOXCMhhweSltl6iTLwLKm+0a7ZgVLLS65yeNmX7Pqxt6
9us75mUhzfhsORVTwLeVVD6yK4z6WfMqfBU6f/10Rb4oogQZeHeyP9R4ur2l0t9x
UInp8rnCi3GN4udtVZcJDUEUBux5Vc4oD/I1/o4pDLhCaRZBz3BTNRhrF9excSYM
rIanfhLSbSMZ6oTI4oEIsyQuOz/OrtFK1WOk3f0n7IQtfdKcIW97elsSjFjczFkk
o2QV4cDmfj0TS1HmPhFIJfxMhOa8O7TGcpfTj/nOZTI4Z/rSm78kB30UFgoHL1/2
XUuKjrM0AiuxQq33RNlfpScckdLaYWtQu88DXnMX6ojDh1eR/xZ+UrUa7Xz/nIN/
CDax2l1C1u2ZH0hCASAtBFyFxRw8RWudh55OChZlcHTLYKG3pYJTs2I1m9X+05Jx
38mLSa0epJyX9WqBg97+ZvvvbsofAk+QEZotwqVuhTha7o4E3dk6BOFBEe1bthah
LMbDD8fa41D7vozAbo9j3OajNacTBC+dxauMzj/PXWyJ/K19WH9Q6kRAwugQvq4t
0JCqGs6ifY/0CRJMWa34t9G+ntWx6gAw8FvqBnm8Y0RwTJcQHBc8DQ1mbAw9q49P
7SGl+6QUrvDHlIZfiCXbCSAmob0iSFYfSu7Tm9ejlr9hzlcInuyMtyNvGGUCEAB/
pibqPQXFzRaZUg3MumS4d0XT5hyb/hRYWYl4Oey0VSNBeQ7M70kcK3X8oFGhQ8Vf
y89iiGcN+JuE6lOmdbv1/ceZEX9+//XIHEZmglCKl9AtKC1dUzd1UMcavFur8mO4
wk9NVzOUJl5iCRUWQ7ta5if4KafBYjBXEeyNo2zDwNKUb+uBodx1SRDot9LzcLLv
7oR0QAmcd6T4J875hep6+IKENg9gCQReg5tLzTY0OI2B7YBhOMJ5hibY6dWW8mpL
GEf09mld0BRbrBQtHMOMNQwlFQjeWA1bOVIsW3xPuT7+0urCU4suTEyGb+xIibbK
4tl9z1YkzkGgqZIDIRMSQhmBURLA69cVFcOKmhDEugacSeBqq9PF8ou3IJmpt56c
ngrZ49nHG1qKD267UbMH5zI8Xu5vu10J1fKFfZJVlJd71Lzn3rw0OyW7fhBYkd/6
4kLzklxG6ELmxS8yVEmb8zm6wpKNkBifcHqbfau+/80dakGUEk1paQKBl+1aUm3U
KXwuS1/Is1W7kdgUE4GVLDE9VDJihjKUnTac3zObnxwHZ6oNsan8VdazkAtVHdqb
KssZC/bxAIOk16WUGwLsBSCjV+gr31XDcQ7HxDuDNNyRZAsfWIZyk0vAMlWV6vls
tYCOYAr5TSaXLJg5qy2vT5encjTL6tpXOMbJem1t6qabsN94P1wkTxm9DhZCIusk
umxj3lCBDWjz1eUqtK8S2XbL5Atr6qS+BhMEyUtfpqXQKlP4hPji+p29+2ETX9AE
lx/Vro719BzRzMW3BoqPnXZ/SDnDc69WlmprnUMfpOnOFBwI2JZkejWt6wZlb6cL
e7do12j3s6C+ITxIOLsrzROSDc9gftF3F6X6BvDV+4lQenzBkK5wQPYbuP47IShT
x6q9zhmf+SuLGEvR5nrBgHGTbC0clh5pUIMrbgjBcXUgkxsc5tiiVCZ0yUm0ZBwZ
6p8d8YUJXvzb6wO1f+OypeHvUgF4RVfKrBeocHSAq0ZzlvXDcSZJYVAkoewX2KPf
cM/sPTg2Q/m7IMgnF2XNMhc1kT+rUtTUnVyt+NVfVVMc6gb3+zmCF34NnjTSUUcN
wGJnk4aPKOC5d2AwjTMQVRmt0xyr5Oo4WPsaRKWl4iZ1DHYCvQiMU7yWxsDZFQTN
0SI/UPDX505M97bekTtFSdsBq/tE6ekYHFQqR2r4Aa/ou51QMrarlo0f/pgDG/e/
qYuiWQTFSkYVFH/seKOzto7EieLk0qIAdMLdZ7urj3rPSljHhBtT+g0AazKOsmWg
VclpYGGV0DuZwVKYypaGfwOPhpcF9e61dGXm5WIjuwFJ0VjenmAYqugD0dQ6rvHX
REGNTw380Mdf+Jjlm8IXY9y/63TOi4G0a3EOEx8wBIrAZSvE6HBA02pCGJ3HUQGc
1Mb6XRlO7hBiKmPqTH5eYNq65p7U9UH2YXdLLNQ6ZYQmBTDQ2C3FkKHIPZwUR05I
M5zpfgr7lMfPVQPGkPZDrsVG13/cK0fWF+I4nQlpJZSkbI8ZL/ZGP42bW68pn3Jc
IAzzHRrA6xooK20IPA1lagDmAClsQbLA7vJUNTunxRvxa4wBn6VO2ouRsuI1iYhL
r2rVycKJ++oWF5hZbGpOtUxIKk4zhWTtbvqmp1l9oO1uzo46PIwvr0qcEQi5hAa9
KTzdoG9gakfnukX+Mm6cAaaSEThtgKa6KtMyDCpEr49IafR+LQ3a8jddF5FSoclq
8vTVMVq0C2s+Y3Xlm+YJdQnXVmAM4KLkiaUcLCUNqV7Kso2cqGsw1jvkoKBOq88r
OR2BbaGbIeMqD8zHTNboHNPlLwexyfSP+BpSwW5icqMMxNEe6a7zNVHP+Zlq8RQa
T1lcgwZvjl0vYh9CX3knf9y+FYi35rPfvOnDMSwWrjhU8uynBLUdMaeVXm2C6INY
O/fYrntz6/rHK2pnFRcOzO0Rn91JXIIRY9jnJqpRAT6teW/G5R0ypsMw6ZfWODfc
SUW6ZePp1FSB9/+5BjMs5jGuPV+Y/XQnv0psVIskAfKPkQ6ZttHmKzj9Ti9tcPSe
2c2eQ3gNK0o/fR9DwpuYlntvM9oh/T1XL2cXJSfn6fI10V2tSkE1Pi2rfZNYtz8I
+/5tAtQsLM9M4PZXD1w7oIsUhTta0A4lldRyAUrqgJBTdjXwU0TIWHfIcmoPP/4L
vhmJg4RXc55R62yJZqQu+FdhvpAuaRcDU+rlSQ/lNeflq8OQJmdR0vjG5XweZKfo
M9ZdqYlKgfO1pKB60sR6dZDmQrU0tp9HSK7zixztEyVP4srAvoavWuFPioR5SbNl
wUkwSG2v4yyE2tPlZmKLZ9InMA3AYEyl2Xip0uT0mT1CsXhYDmksFOIEVCbkTz9f
Hw1Z+Xw7iAeHJhyXLstFn2J6dqwuU6V70YEDgsD+7FzzXbtGF5HWYR5taL4IaY5w
91Ie60+oIlI2ztDUlrcGAqwYncsKHTq6IkRpDdpp3ThASK7/x4YIG8ksaeUigblj
wp7J/siBblenZJNo3kQzEPHtPWC0uO1WIMIeWZEpSq/fg0GBOMtda3C24ZCNBZxg
lsUWL3GtM2OWA/J35K1akYaBOuE37fOt/Ex3dh7kL5Emm31ZSXhsk+LMFoiV3SvX
i5fBbHDyTWdQVV7afAMJMIMloGmbt8FJr6iUHuL538Ov0M+mzdzMLWRd6ElS6Ini
uARPKczp4R/rl7mIPHrtKaHHwXBRA5OzNpPTcukczbbvq6edEVaySQz2S/p3s5Ju
q7vrFhtFBHOWiaM5eVRxIyo/tYYTLa/XBDhxSFUtAhOnlky1Av1ecN/1qSsd8XeZ
vrxthVGZJkPdFa1QhKHT69dpTGYYMuDd4lcE2OSjXLqoanPkZfXztPvP6zQ+9NDn
A4uS3mMvO94Je0cpVEx5HARLqULcxl7ltywbJTct56z+gFkbmfZavRPa9rQ/8Dzb
L1YvrrMMetfHNMdqFlhgFDPmBX6KDteqz8AsQFsU1K+o26ON2OQF8CXbhUAFo/PD
X9gaKgguBggBLerTfHBo62BE5B0e6jaQx/DuYv24WGe3cjJBD1I2CDSXxpvvaWUB
aKSADFyu8MRRjAX8NSqNqYx78HJnN9oSyrYCqPkYDJIG/A3Ccnw+1oaG7QpkmpqY
ZCsxWdiKntzCX6Zy7IgxMg141mwx+GyZ9I3qZZoNbh/RLoXwSsTyn3bTl8/9tjL+
6IdHOthFWtjMZKvpjha0AX4531Xrv4BtzXrYXbxGemnqEQGq1X7hjkf1qMIOjSLx
8zPZfYJWBqMkqP7xM1qfB+XyctajYokDh52p1m4L0DS08avjF1JaL5Zdc4xVA7Ic
nyqdBbHoKRj55z2JWDszBzSa56ZfQio8IfFA5CZz5pIxZHm6ZSHpIo8N/nMSiTdQ
zzrKWdgIrkJTWPtHkjQPq+2MaHBV8fWKTnUNuWkhkSaTHAiOYRrYww4hycUqhacw
MuvyoaOhtf9bhXtkUcwmm68o4TjD+WkNlt9dsyJiA1sgQz/ptHLCKY/bJTObdv4o
JW+pirZllYQUS+diKKp39+4LgDVsuKFcMo6ZSdGyFuUrIqQYrx91sbvhhzVwf3k/
qsdGB0Zj6nY1KX3aTiJsbhbBiNkIkU3Evh8/X8sEsrnphLuPLH5oIpLGIFmcpnrM
Z5UlUwKbgh9Jq/V3LpjlOMH1JYtySXDwk/G1dp2YD1DA052gF5n4XqvOj7L+LTPZ
6UE0yb/sZo5ySG4vCrex0luSqzsKDTy0mkCKXOcypYkiAg78fpTw13GbwPpiyFBd
mbBEs2opNiE2nQdWikdsrYPhYGL8ynyIfmK04QWXo3+qBgRgc2xHsWugJIazDjQS
ZPbw3rgBIGajjfAUuoSLWqjc0v23U0Xyv0CG8okVr+N+TqJl8jkmpVUuum/BcKsu
UOhspaFLG4kbMjrv0S4KZoF4PXuTMppOfLFIIdgynGc3mTJkhKI7v8jBne9F0WNK
FQJyCCV1o2c4A1/7TaXwC0QV+C7kTFiw343H3QpEe6caIoi7c9CqDfbkS2yTHDmx
8u5DzH0TEwqnCKisOhoZt1JoSoyEj/+yXKfiHJ7q6e2K2QAuoZZJK3sTyJ/wteaC
XRiy2Ds4iAiVP0GOnArmxEEP8YVlHxdZju7lR5vwZJKmz4hw8o/CbutNsOo1uaew
W3V3NOkmM4PFMdqtuM4W337e8eUNGRyc9YNH3OMKNHjZ+4I2+mr3GNhXjq1KyuN6
e6XUQMBsPGZFYQ+Ko1rQMTYFZfUpqRJ0K7SHk4wgjiRzAscoEbNaMg1CPvBGX/TP
zH5GaMbIoLfRLhb15q3aE+JkecnmOj9aesCicqadhNFbx4JInRJQPFWDkr2FsIWF
WF6MWPlAL83MyR7DrO+OM+q7BfBYJUFSqSlJHeF1lVPeCSwYnQKWH+4eDAC7HPSF
rNFWYwE42a+amhNIijyWtKhpLb4q808KBIpq2e6dssq6L2ELbNP5NgK/mzs+FlTy
+RdRY8wlk9+1g/+dDByWKY8vAnp300v5Uwfo7one/hz2ubuArw+8aYFn+d0oYAmA
3pXUuSs8LXY9eHOR/wK7awBVgN8C6yuxYzoFnu4WH9nJ8VRsruMUml7WhWCvezU0
dN4zoCWlFJoGsMT0taVYwBTUw7rwiK/7DZIXHvgawyi20ECHcEneFwZYnx0bdWvG
IF5fWyshxM1YoT9qZF6Ax2sr9bZlYG6v5tuIDi3jo3czgCEN/OxCWcKJNp+WEiSn
Sw5wtpFLp/JwH44fJKUtMJMCJLouyEVeENAbXOP8sZk89ntWqoMfPia+YDG5dcVV
lJfkyDSefRkgakei2N5hEwRZJozOjlq1oT2w67oNS8MEmWkaVy/TAUjt7rqtLwgT
CFWkz2e5fTDffuR6pCcIH2Y0pBLI/funsibW2NtSVb5R1Wc0CcIHxhDwcPgSW9lN
0O08lgWTg9DtqEARbHQq+R2gEV0Y9nibNqqKN5Qp6jucEKClEIQaej6cgiD2INim
SMwVg3YIVv2HxbuMobioQ/XbQdej2YKhM/lvfbzxN6Yu6MvJ8U7ahWvS7FldW1Pk
vvQ3mDkRpD3vXKu24i0zWaDk4GN8uKjyMft8VCiRbsAclev5vLWhXEzSMzoR0B9c
n8Jes9gZ/ftpRoURjA5emkdw+QGbKF4NzHGVJnhPkdfn7Pp0ELClE5O8655FJK4n
/V0VdFqA1CZTdVFicphw5wFugQEwqRPEJ1SZvqJki+AgaGUQBMy04vFOPHCAMK1m
c5b0alYT/OqXbKAkwKcbVufFct7lGKlWI/LbLcEYdXwV+XvKDFeRQ58TsrGA46xr
9CtchWpv1ZkKkK1hvrzRGHzPDYrgIqBAyNc3VFuyneZHrYD9dZOtauDVA4WByzez
95bCfeLbKlxbYAJnVJQcUbIQ6gsH1VtSxFXnZArh9oPG/LKckKbXMZ05sxkPNzAd
5ejna7Z+VwYZUm0vhiOunqZj3YVg55kSPSd5hutqnb4ZJjzbMzkMTd3ruhzwtTxR
2jrlkiDm6R7uMjIpEvRnugJz2H9eweN+hTXttw0vEWCpF0oODFClzA9BlUKbLL84
JrywBwYwx5bDTqJs3KC3E/UGCnwzoXED0Oqiu8CCnV+4heBBKBMvL6Yt4+yZoQm4
1cqGD2oHBpTVTWcx52yM2R34vcxozDdjubrysBwPh07pTUtZooSVqkBLRvEk5ikG
YFTqU03+S1E3yS4W6pNuAsrJEPeDzF9L+UEEGElPCa0EIFgakl+jWXBHcocDBqvb
Duc1sNSywus6sLziWo2gbQ1g5VXUZ/uHzMKBNm5VQCLfy+8ssprRwr2EmI6eK0CG
H12K4kyTOmnL/qbG5jSEGyqmPpCkFvXs1wr4IStplTpHLEY/KJoVsWwNajzduVUL
98dnmLJjXUUQdQcximmzkhCd4RRjw6nkJ3Af61guJxDrnjjqECc19g1Dco1rZJ5m
W1mZHKD4uqYkgYsyImrCrciyhvzATBtTmYllWuyFYWdCoIH1/zluNCNc4IevsJEC
wKpbahmcPddnm0HZsHG5yvw0XPSYOqpUxk98Gu5iaqVWz7xBrJRP5qhfFwg00u6f
kRnakrVIyPJtm05TPJNGGRmT3Q/XCSnbclC6C0w6bfmGDbPrmR+ICYlkj6d/mjVQ
dne2f+2RwFsPNnH7kHcz61p73pCRVDsnFure4mQW/MeV3TZ3hABQKOBXp5N95Cpl
DJ0wEv7+tvDZ/QHh6iBF9/1jlHQcjpclW3dawEej6bDmForEKrfG0NAeBkNJAnAl
upMiowkuBPMvekSIoiEhCPlwUSIiHWo2h3h/r5BT13RSHTkMIBMSVkGUadxGrnhu
CdKlYCHgNzl2xZOhLwgQOY/tivf/7N/7Vvwj7YOiq/g=

`pragma protect end_protected
