`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
qpbU9KpraIbhLtR6gyGVw47QEMPG0+9Leydv4M2WTX6MGaN9terWGY7iLQ+/VgNF
HR2pVURVZfA0pWImM1xpvA4azajqtsaQjhPYVy5ZJl8lwNncVct1VzbAJ/zP64Wa
ZJwmVxGrE/7+q3Rtil8tIKdaS6oOsnKyiBskk8Bi0FM=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 46432), data_block
D12NSqDjmOkfN39tDGTTToTPcIGDbOIVUGKHTLcHSB+V3x1PSELytYJYHfAbE0Xe
mqLpCAiqanllq4h6Qft9k+d0d2FYNBbQM5sb3fADkJq+mqqlOqs2TgQ/kDmrSnBr
MkrWogNLODnqIwj2vknODf26RHnwpTH/t6lMMN2B1pr2jlHbAtT56GRrGW7GC7GY
bQXKhKY2oPoCQ2ynmFA3fDmfPgs1jypIx11/vL5zRiNeQ70IxK8AWbqXf08QxkAa
1X8ipG0wiqDMj72MUsvVE9j9iTdYJwISdg1blHTmSy6KsVec/brxnZsix1aA7NEU
yapzoecOBUaEX1gqswChBZWmUKNEElt1Sd3oo1IxbvJTMXwHUUGxv8R/56WF0iYc
KIZHvCQGhM5xqSXnpamceJRmHtEptOFiXIgH1f9+5e0BJD57P4Z7uVDpTqh1uT3t
KrFZ+0Zg7/cLzC/xVhBV+z4bmSo1dIEB19LGnXrgT6rME7XK+auBJeUgClm6qxG2
2jVUtYA9kHmwJvqxBRVV+g6YnrWNcXbqGwndfUDLX/4n8lUdyY33yok+pzzmDbK+
wdoXmKbIcexnBdloEO2poCtH6+72euWAWxT3YS6NIjHSjzyeJWvXWbR9BJXxQw2w
NexQTnvcjYUAzytwTI6FdxX4yWUEWMqLQJ93wbmH72qKC8MMzG9QVWAbIrS6MgUi
/4UjLp6ZeniELf2tBkeyOzUcxivxcH4OU4V5OOSaI38ben1Qhyu3DCFnT8ACEsSH
hw0zmSCoDz67Hc95A+V1eZC4hvfyRh8g+H4nwJsR3DSsdDi3pkEzRy7JPfzOnHqO
5sh75ZY54o8MQpI010t9sHAcw90+9X9MgH73h7y77YNqXWpFlhvA7JmSPLmgi6+0
tU38YZD4LkGC0PvSPwlCfL4Rq+TlGfl4WoGc9fwXmYBYjr/pI6H7elb9/+BL+qAW
6I/szS6zz1nEEn2H3hUISlsvOnnXvgzSHixjq6QMtwfq4Hp+QQG10j3/kpgIhxGR
Wg6efo0OC8oXJ7H3wgCZCRP/L4dW2Nef1MK0GcQ9i6HH6xY7JYq/0IwurwRAi+M1
Ymrf4qMi+haUafNlWmykkACFxWdbRex3TN7jYUDbf7KaVHlP6OockytpaSgaX1DD
dPbJcJpFyoAoglXokgKD3emx3SE2MZQl0KhN0eeMkprsMjhDHUtnU9mW42SuLoRw
VVaREW95aU84yNoeS2vPG015o3WhpSL37IXNouw7rbic6DGb9vCLtOC+KfZzysBS
caiMQ0Cdvy9UBTYMU6SUuVOkLeIO0cX6HuutaKV5TG2/XNHNE2GLrMX1aHg3zC98
aAiMu5LIRbbTSNfNEv5Yx1wJbM8MHStvUmcTKsVUCmiF99w08yHc0sCou8cdn/ua
2htEcu5puB23JE8DC0p/eAnicje2skcrd67mVAhvK0k4QY/b6wchMYDsj2XWTXoe
OVF1nT+sYrvsKg4ogkblEi/mW4FFQhhbEsbq6N34ywhKWs4nQiylEzMz8iujjS5R
FYuSPaT9wp9SQCMqfmJL9y3rnhqf5HLqNdNrYObOVi/a8VR4FwM+1imtNbsKRl2B
owIhHF1RkRRCTxzS3JXJ0XE1t9VXaFX5mxBS/eklmb35nEXosm+qoRbbXyOsugA3
r7LVU0Lw0ZalV9gOqjSg5OaVpnIM9rTFPCP7SWyUMdoxyznSSs9TGrb8EDGLaOKl
fGRrDDSJ2o+QD75hQQjiV6RQV0OhhmEx9GKLu+EsKm+gZRzJSkKgGXaYToSttTkJ
US10Bq57jIrJkm5d2+QZq3lM4sSYUkPnyt/U07yBoJ7O1e0N2sHM5zijo/tr088b
ulQ8c27GlHNCaWnt0fTKicRC0UueZlHa9CneaVzBqHyVFIyCzXK6dygXIJ4uA7Os
AXbAlD5BpZ1prgRSWy8cQ5LdFR0krjYsLc3IMylclVHvUDA6bWoUV1gF1LZovsoA
Iu3iLsALmwl8ph/BIJag7YB7sZd71j1+YXjTApjLo4BusLFV8CEi0kkGWDJF80JX
F+CXcrzqnMHbgoriNdURq/zVR1TXKZPAdrOPhF6Z7AgSSjvcA6xTWR9r3dSgx+9o
4eUIDhr3lRZgD1TiJalrjKmfLBtOZymIODf0rqKKHhge2ZNsBeqIbMO2yuiw9r7c
MnyLw5ze6v6ZdRQrDcjlR3zv3fIF05syLqcPqxV9cxNNvHBmw74+c2LdAmPdKiGA
0WAG7Y7W4w9z4FKG53zv7uZx80icoRIWD+kQsn9Y/WFISDaVNnet0Gi9gMHP3Xtz
iQbfbe0PpjrDXNDKqbV7XUtHtZJMRfzXkgFRN2Z9eic90Usr6dafqADfV1VbWOzm
y+lO9oYsnaftEhQBVSSNan7xTq8tmQIur5C4qr4shgxmvrrP9rGtKJTyuChYrdTK
VMQTPPrQ+fOSOZ/R7k8r2KhJbL4+JMbVvtoWtBRgOFyNcMp0kmRryPlTyyMhW4E6
uYL4P8r7br4E7pFMjrv4dSnN7tHk8R5qivQ71kt9TdUaw6lOB+l5pq1o8A/ZOkfn
NIDHckV9O0613JtfiOJDGZACOm8yTdBWbK99SW+3rVKHjWi66ja3bDa1cTVQ+uvq
APUdVyMNXcWSaBSDeiJcjqwe9QDUr/d39yzp16dfCR793vIicdZpI19iiMHzytmp
yn1vJeDKkL3lsv5Ygrr67NZP60z/gSti8EMdvG+OJkWVnhLY+ZjJAf5WiieNnFDQ
B8lZgSgxt1LU4rpWR16CZRsJjwWIAwetqRpC4T9DxIe/XVKrQybdgGzOmIHFJFcz
cqiGjprkwXR4lbJ22wj1TnSM1H6L+Ap/CdVrXNsgPXgfEFhex8Bwaw/ksR42gEAI
6yIzRoaYkjVFSfEi6twNAwoq1UQN6Q0qpg7973nMtW2LooJ1djCkfkGj+l1Btc1P
sCVg/fXEaj9gxDR/89OFexQqSVTxHUyCZYd8JfUTcQVfJpYmsn3F84lqcFjuC5Uv
IMek83Yom9SZieDOFcddyPPDUqbN0XHPXtdVmSUcFBS25YXQFFt5kpv9GwCsg9rd
Ad1ZnFFHo2gEQ/rjKrSBpTAQ6mnCGCRptH7AYkLi6lOD7c1KQXtJwtwAmA3hJt3w
izlRvqfrvAuDkUh/J7k0t/ItujW+jsvHMkF+Npwvt6wPi/1qJLLP25t852ZzS+BM
hVaKWG1wq8Ymfpkx1StP0pmryb0y4Iz3ckbB8ukYtGh5EBWKq97nJf58qOhsU0HK
R49r123iMHxmI8+/G0YlWnuEp0WCyzyy26F/4dgX56EWJZq2UtMunOCdncqH9W/g
S6dtDAi185zH0kH8WJ4cUXoEy51TMfwCMVK8DUAAlsrt7IRn0FuGvNR3OYVN8w8v
BV/23C/UznD+ED98VDi+nQVjF7W5wVCOj/0QR7weyA6LkxDnle40kIIfSr+XvP+h
CdS4ZGu/yl0CjmP68HvQDhQzXKgiZKcGpjklslTBI6mHqTAV9r4Y2gzRuaF2zvE5
jF/2aiTO/r54NgabXu0VsM86OY75p+pKJ0FdQCa7L0QYiW+W0xfteq28oHe9youg
xGcYWRUXBmEFV2VPBgbNKLM5jSHB8KJEUaTa5SW81wBW3VwJiO/+TWq5LXqeraAF
5Ek06i7FGBqw/CwBlF+2fBWGXZ9gwG9T4MiTKqx7BtTs6UlEQm1Jyt4s3WmIv2ID
3nxoLcYBb672uVikHjWv445HafMApoKaIO8zI2mPHyM3L6g6Fsws0P6QCf/7/Rux
sTWH6rEyUkreUN0iNRPP15mAssyqn7CK6BgSITmezThfhwZ2YyXwMjJQuWxqawPF
rABrFMZqHsN7Wb08K/V/98BOY8k+rfYQ5lUNE5ilpRJFQPsFNkdKZ2f4RkLNvw6h
Ab390jILZ7K6m6YHTsehZaeUaGsq+nUQ1WtO7nAqmuwqBVKShLunBkVOMuzLt0XB
l9duujpyDXOlvuSvMKqEKt91jteWKxeJIZ8pyEyQq5uJOHkT/FpvrH+1ybF9z59Y
EPCzBhzhf8AlgD4V6uL2tXz7YnXwDj+9pr0H6UOZez0VRXqmxn0lxwL6ipngM48g
EH3qIVXj7j3EhvHz5mzEHuwEq3yIwxYCkqAeCALInvOzBVcd9tbsDkro9ypoWxka
QZ6G1BxjxvzM9lZaUTSIi4MFwk41aT8Pn2/RCKHdspf1pbY4yURUn+4iW5xN8ol/
/4NT4afKV3F/9tm4JEhWHBePoR3fchXfpUmM32508DnY2tIeTCSgTAntcTcPslGY
wTd/F25tbMCtByJg6uln1kvVkO3uCSmDecDt+nzDAdM+skh1RdgyMH+845D1+LqE
OZSvtTCF1mfyTxirLxuUqs/TFaTtgd9KV2AUvYjtWWPnIup9rOc5lvsdOu+tdeWm
fCTKRXPS5US2Bd8vPNSeHXsb7yJBbMZ/1ZGoZ+3z0WeW6CnvFYNb0VSyBKcoGgVi
RNSgHLyBeVQ99Z0WfCDtesQ8NRwM7e0x6ldXHlKfydhMLjCfWhYljYxKspWLPlLW
FhYT3zRipbIR8ifUObIFfC5+mDm76j0d2EatDG6GELm3cuflymhhJbeWkDyW98v6
MJqdAipQCn1ecbVNSsMa77hv9FeDnwapqcjp1im5EPfsO2AvT0oat6toaRvGgs7i
vAzLoF2D/2Nk44df1MzH9dTEmTmzhJG+urgvin4ozhxnbAQTudcvBpyh4iBnuHKN
3NAbtBZaeBe2ZERwSvgEPmbEbdqNofAeJ71x9lI2ulq/ODmbpYRanuhJOVE6QvEy
WYWpJj/HIo0XlrE7iT4jEwzWrcqHltiGBhaU2yxkH6OTQ7AONZN/+e13ollZX+s/
82IRjOmot6gC3xpBpygBpCpWf7TaQidyNSRlye8GR7u3UWnbMew3lIYakZMoRZnj
mKm/kRr0mA8sK2ZYcUl4guQq5Y0LQ8Yv9aw8Ka11l5y/feNwWRYI7Ufq4/MnhrTa
Dv2TVScgq+eWsn/KS7EmUmS1qRsOAzsA/94Bs6lrK+jp70b30W2TGTTCVJ6hDQEH
SGDvWQCB0r9+yqKA3CIWCttsygrF9oumlVgfy6OpyJt0pUzKoIhVkDZKQGzn4oaW
W0z6ExQmbutOX4PPch04aHy+dXSJTS3QCuTrjVWbRWYXv2M/22rX/1GS38EIi/o+
GBX0jp7DZGzZlC4ZHPLpAdlJexZZ+7gNfZ9WKFXJwWycMnLPUpCKfHjWyZiFTvGT
IrO47TmbY0gIuW7qbMgXm67EX2gY7WyAP58818rgufoM9O+DyZmMN++XzHiQ6ZdV
a3OwBABo6F15JL6QPM9F3Oy+NC0q3Z9ThDnOFl/80d1/Dq4uWFaCiQcg6+SNS3ah
xLsSOQkuQnfVR+cr26TMPgat7AYLFnfClTtZ4eFoMsqjB0lGb5+vlAiNUNJY8DTT
0vNpqU1mgR/EPe62Yg7PgAoc00BKRtJGdpFKaleUxJ1vf2zCoSRbq7mtncPLT7+c
fsGTJetLUM7ul09ary8Amw3+551OWPdttiPOv9oAMVXNsxIyvRk3q8pvTgliKk56
MEBiTgHB3JMKVwtEheknZL6R4bEvGV8/Vy3G50D3qAzcospEGvOQl3/eHUGYFqBK
IYDtMgu9NkxE1UtxynvBitLgqLvrmSiq3b5aNk0LVLup6SNkPeTiVb0v8IGM3UVL
zo4UANTsLc//PiRiQVUQXHB70Vsoc8uftlA+GrrJEuMBRFkBk6D5tluYgtGNZSBb
n8JNg8s6hiyyvNFO+GF+tTgpxueQIyHSxs6oT2SjdzL7zqoBuCckE6BBPqawbnHV
k2hSm1U96IxCNErAVkC5njIWhTQRc46t0gII+vTxuTLi11W9DE8AcEdn/gn7Fqwp
b/dqzG8e6pEXnVjZJh0x8eB6Chk4CXBk6ErJn2SG4HxCBFQQFow2QkZwb9DRPiYf
4SiejyE3b/MQmM/Lt0+aBLQzQY8kurOXxPgzjipKbnrLBVJ5/N3vc/1y2ekXQ952
k/ir79TCXGU1vWtuAryrRtawBf6HDSMqfjXdH5YYKPwHDJ8YVPG7b6GubmYa/JWY
gWJTLkTlFYiV7o38TZNR7GdZ2VoCZ+f/sJjU5VqI2ME5+AqIYXpBEuZkodh9Ym1h
AuuZA1aLyTE5PlHaTAhvX26pawD/r+WBfIkYiylPXHldRPj9jH7y3Nck4HypLVnz
kdqy1k+4kIfSMm7qm+Yosks5q9XQZuoJWNb0ffsGu3tg6IlbOxs11ryk8gNnrdKV
jl2jXv8bSmkyXUAZrnUVXcpfin1WYj73ysHkVpWhajvGGl36khLQIDTGn3ky+CoX
BFP4jyk3wTUMsAY3EstU4DbfgO4D4lsI2eTAKolUbq1JIhED/myasAPK7w2/vEIo
QpSaPtYw/U3mTEGhIUimqHhDzouCeDmhdfjSF1kvI93OJA8PKxe10tL3g1Gn37UH
eA2QzDrmNqoG2hhDnWjuHTkCl3VdPR41w6x23koIMh9zBoPYH5Js8J7SN6vQr8m4
rGQGy1YiltYYsMeT3AFBvaGVMbv+lG3jnuWCS/7oUJzCUwgkZ0CsM9bFuEfBcwBr
Unzkjkd6SrRbF/bcIIlAggKlkZGrJiN+WYN0LHc+pLKa3tpqVXvv7nzzSp9DyTtd
qYNgeE9UzAPkaoIWTlJMImQYwGByHkyGWxgG4qprz9w4XEwQntoAnsCn+euCHEyu
vVDcDeGUm4ULjwJ1n2FFL+UQr+K5coy0/jL5nTvbZgO+QdlfzB/eYWUTExI21Odn
svXiufLREe6pvCrU6j80CA7dGiDoozPJ6q5mfi12iIBy8EkL/4w2bzNUQ0JE2/V4
6ZbznxYjj+WHPPcIrGkSWOriSWO5MT/RCKmricPdGPOteQxuZrYeW7GE2y8rF68K
Dz2KpAf8NsVTdFNNW/Q8MFoAvxmtz7bt4mqORGniQKn5AktG4S0fGFTN5IjZRd0D
N/to3gQLIIUHIysZZZmdyaOBU86xzdByo0GdllPtoOWJVLuL8t/d7e1lfL2pMAVv
eTGhN4YeUXhZh2u9hwle/TLi3moi3qll14vKyKnU02d71tlZdEmaFfiy+DjUNOQG
Cf6kanWIREKYb5vP7i2LCxYa8QElBJUxxvePOdM8JN72vNE8WwwxkRck4Y7taU3d
55nu79ce3Qg00EGEVRHKhYBsZytWuskKwMbKZPNavPd5NtzpZN1Un+2t9bs98w4v
l9LfyAnZfphj7w+K+DeGOIFHDWbk/Am5K7qgJsB287Xxkoge5dJLM1EcdC9GNwsj
BgA5qj6gFVlDi6g1/w7as7tRSMAZxfLVr0sRJWIiwiaFP1nB4tzygmdSSN0xeyAg
aTzuZ6J2xYBhC/lxudC1wj2pe+1WV1oCV8Oi2w22fUOZJ+kjBPMj/iwWgY1nQHDT
awyvbpY4xPu+j4aQfHNu+9PYEf5FlW/iCc1rNP791BNsneRWeVPq+01ZgfRXFCI0
2xYPgCggmvaXfkueC/wxm+YseAG2rEJzMSWVBndS78IutVb0CZp4cqkjQeh7Xb9w
ex5G5PoeBjQDAJXFFwZf56++5eUSOWiqyNrtVDSuiGbd2NNDLCOnxW6JhBkXPvRx
DfwIiw3mQEBSF9CJSQoRCB9i4gKsURynepJOFWrPla1JEh87BzIWVB17F4BIFMj7
apGwwF8jhVldFuB2Aysm1/StDuc9Di/700AZqM66zt+GnFYFc4dbfnHOErIQOVeY
MUA4KsenTVPq4oa7urjEX7LHqMrYH1YTSiSglU1BSXhre72Y9aMZ4CnmTHOCQ73I
RC7pVOvGsb3XxrSjNE6wKgZrcM2480+AZ5hPntD/hooAi8AFWX5DrwB97P/waZZ0
JBHcHmi5xVyRe8oHxjZ7DRglPuTPM3GL3U+BciLQv4fVXcBcT4algMi7R+n4qsOJ
tpbJYWjYl4FJKFVCSlckqviBaPhbDKz3HKJGMX6WGgWKTrk1/kOk/+uR4auPNNuy
fkxDAhBnk2NOkVG2mLIKBjuoZGF05AG45z3qvs/KzYXUWJsUWnogFtpumcmA17L8
z6qoCt5vAiocW+57LSORUL0MX8FcN/vhbj/46ZRKvScsefojrxN3X/bpaPup1qiT
YuocR9SVgV5JZsrsxu/9Tt7FxWEwW7Y1FLtHO/gtNX9RbBzHapL48BuJK2hRIhb5
+KosxeqnqV86p5GcNpAgeAXY4MdwogiCuIa98EzvhzyPGusS8Z8Qk2dB9bRW92/Q
+sKH8WbtQ/hsNWcLAraY7ZGC62ddPIQEcsunpFhuS5JPL7E46uYA4LWzltx2Uwyu
KxV7j6PwHz3nixY64wukciVL33wv4zxYr0S8my0mPWGEKz0s3C6o4w+4G3bOC4P4
+FMwXaYzNxhylvNNWlAQI3VvTcVdvvQ/seRp/PkYSnfQ3Z9qctVkQjyAyfthvGkC
0ZnTfIaRRNtvxjD5jAwhriZLYb0wvSYFzaugTDoYs8+TXE2BLH5mFb8rxJSgjl6S
ppQ9DZKoimmKrBO1k6lsKdsWRJdUbx1xbYUxSicp/CrLiaUlA1EqwPnqqSBYXHKi
+Y0xwYXsn8jJm1CpZHD2pHwUzf54GuUnloMrXbNpIL3Lg6yVjEPOsXMyhJFDoYzX
oUn4N6e5+XDUkgkZkiAF0HSxG5oNphWses/jGDkG+CjThOZXo97ywlmbPEsDmgEU
/1b9DZL0ejk/iWkqXa1bNSqPx6LXoa9l6oASTva83Hscz05uiWLPtN7Z9YrUYrpY
zCb/fnHX52QdwNiycL5ECadsYpZuCBR9tn5gf80rmgnVC1Jj2YgHd/WXuq4OjFy6
ORki7GGwz8PwRj/9UHaW7vR91ndZDzfDIkjlJJRWgEcMYgy7Jziv+fChktJNOTw2
Wcf31WvxOyyVHjqYBzTH1KDPL42yD4fYN3eMRFN6gvMroOPrXfNqye2P9aRXJzq1
uvXUOAbDJ7gCPwS2f9oD0subczt/3xHfsJx+Rcu5MnPK8Hzr067vX+vXQ4lPbkKR
sOBB5HGuGdaLHlpAxeY9sMGPOLVLRRncGMXNkaa/QrDLUAYAB6mIu4oDhJTq7fHQ
kEbnkItok6M3xfFDGg6Qv2akXTVclz96j+EZAO3dQ1hJPVIPdX1pGcmuA4ohzwHc
OEh5ntRc8o0CIJKj693RfmBRPTKphBSwfCbdB7D90EhjtUdsDGR5zGv5qwlLIGl8
fohG5PriuVRB5Ar/yMAylbeXaouT5WvXCH548Vk2o5lzYMZunit6dHf5VvnJNKNM
Y1niqQaXuWD8Z9bceKPQgFO5Fh3NSK6vXyCGsizxGSJl/Gbd9Vs1juw2uU4xDVu6
1YHGNAHTxc+XKJwZ0Kp85MPChmdXyiubP+VKepOUyfk+snBSB0qklf1RMiwBdBX7
XvvsfnT3U3WWDsZdEnu2QwWYER8zMMTl11kuTUTBO9jupNf46xlHb3qX82ARS+Di
ggl7V/fD1cerT79dxSoyilsOnRbMcmwNFe8RrSOXJ6f9JpviyEcTJ6Q0l9L6QXyI
lEnhYKSZv1MTkusPmWN4BqJ/kqMvJBrNDjQnW+VKyLQbRqymfm+MYqgkr6QZDme7
9mHGtHN1h5opwLbooQ85I6Dpz1na99wb/OP02B9dqhDaZfgN7n6MgKwPjStkU/U6
WhIGshqB3nz8pAdGtbwG32oRM1F69VTOh/zkyzB+JfCuzHD5JqoPsNB3d7Vo/i3g
vQmAS5AxEETy0rltJndhdwlCmfQ/kUOMQ2p2M70YMdkDJ0QkIzFteIGYtaQZMIAP
x51EoiNudakhLSC+DlSIih6kNThbe5meOHthyJ5HcxDB2xiq2GEysczGWnt9qLct
KhyOeTLpYJ30DF1iJvlb5XfaIUC559JDqVWfcZY/GseCq+qU9hjJixzDA6sAnRMc
YCGnO62y3nkogScuqAP6iO5ebu5V8BOfYFy9shgUBw0MHa5XDwPFjSnD++scQaj9
h+leBjHF3i+AfoesgX6qk6Bk4UUz2lfLNPlnVW2jeSjcKWdsRfg2o3DdgdmO8hEu
VVkuwv6SWr2RHvIGNMUa5r7piE/JVlDiPaMf2McDyWU4G525PGNULuQgCWUEBhPz
C1+23WpuGVdtoDTyFoTZPJG6rg2gu60PpEKCci0YD1bRsYezvHnbKB0S2O868NxL
XpbLyPJaWhh6Ij3KVnfqp6vg2jzsMsgHqCToLuMR2i+yxxx1NtEBAOxEnNViF/+8
6lqSzM3xpF51VYKSiNmU2J161vfnfIyMBdj9j/23lTrgJkdYr0eW43uDN+aojwh9
zxfF0nGL814PXNHrGNWNWQNBEi7QeW+U2u/Bpo7SWEq/YZP4HofLz2l9ZOHQmcR3
puRRg9kIyIVu1g9jaw/q8nDwfeLTR1MdS8V+H6y2K+iTj0vuW7tvROMu3GdKK+tQ
SmlUen0jC4VefZzxk552fikZfUiIsSaoKokyXKYh0TnAM8UcHFQGon3AWSum4zYQ
iHX8214h5/hKM04nXN1+LRrEyfqie29cqDuPVUmsworzH4q7sQ2tLBppUel/cayF
xN4njbBhbIUs1SMMHOst7CRUTEycNoQh/FHwMQqtaOV4JbAAIPnnSvOVocz1cYhW
hnjRUPJDB7TwVENa17euTYhUe+KfvqNyrCiIvQkVNZIL6Iqv45VfE7795mW2fsnh
GrkWBIP/9sikYrAYq10UBwyL/5rgujdbO2zpW4HyKomg7qxzlAlpbfWfv/TG9sYG
QYBwnjTa5gyEdcWyTjrF6Rt2wgd9gBabN0AODXnj6G4MIHzWLdCSJk3eoZqiByHq
ttxkHO/H3edy3UpuBFerNuruZ3DDhmfAL0w6BsXNQUz0bSgxauVtXatUTtcog9vV
AWmIlZKNx2mvT8Tab4uGv4yldi/i1L4dHHz5yTgH2XhSVa3ux/v8/UJRKHTAWcD4
Lyjvzf9JGT8LAmE1UZnNGNgpjy9Qe0AtcfZuBVtI9CDP00NCtXTEhG25r8e1OHUo
tmgLlX6YaWhfrqSbVO3Ld9W0GfUy47Ylhj+Z3Y0cUqKbDgq3Dmmf7BJxbb/JOHyd
W0LZZucJdC8f/Sr87nCjEOlokqFwMeUOjKnwR/TiGZRi0BwLmjtYrUlUaorlJizL
CbzMt4PVy4GM+w/+k5VU0NZIUWQv0KBbG9ASIODgGd1OJQ/kI85JHY6lXwF3uFBb
31XdmV0zPFi9Kb75+EH1unUIJKX64RjwVlbo2ttsevN0ddSJ7qtCSLbSY2Vx/cc9
izAlEbVxXTLmeY9fvuuFFfoxIc7mfkU6aRBaqnP3QvmPNxXHAkO5l1r0X61NO4dD
1c5MZfl8aC4+1p3TZkGO/JXXaKjEMaLAb9KHgQlVevtBl3c4EN4RbE89+Lj258z7
uI8NerJr+jK8LnaVG65F5wti9adHQY9g/CcBbd9v08t5iUklwn8QYvWZs7+hTfQO
RpW65iTOfH0hldfpUzpj2YgDEdH0WQyxJSgk3I71aPod1ztH+Ro+kdS4nepjLIJr
wTFteQXQrRKZDbk8iU6xD/iDE2yFbBU2r5sZ13/b2xxCVCjAe/cchNZ6NGNzE05h
XgJKnK7OaQVaUQ1YdR8bcxnyTeQGgajNk9jCmkvl2yMAXuZt6auXLEOkEl/8myf2
U8jE3N2m+I5IxjHTsQOgU2DM5Rt2Ph9ZL3bvnHW6ATNw5UGS8GD9JgZXJs5TdcTJ
GEh7EmJdFkjF0VT0onZyx9xcFRUGGpHYUzf7tu1Tac2zl1oiTWFzcYmUggCKz/YB
UgYL9ztRVRaytd1dgypvNpa75COju+Bc6D04rnmBWsKHBFHpjxAu3uqP7Db+7kws
VwfJ0ctb/u2Ne5Z8Afpw6/3KBaBeUZI+Y/klQ2BmESAtpgTL2ZcT57YmrAVLyyWR
qLhG6K0EOzOcJDfrY9AU/4gN4l95S6g/HWxx3UJ+Ql9hU3kCt5KEwyj53j2GahLg
dSB2EpmmoiTi1Fswi2H9rYEiq1ymDkJxSm8pwNVc7eoh/ElurR7koMPGf21PJaL8
/3SUzrKALGrKioZ/uLAieD9ygrdmZ76DR1saYf78mhL4HpRTOp7kFmOHfJk2UI00
LefITZytuy2TPL5ysWD8Mksyl/L2XSehfYAxaHyUziloi5N7M5EaRBqFcpyBmoWy
tkNq/yEXcph0RL81yassDo0m0WG4iFzffa8Iuh9rbr5kH7rPBhJc6P14STiNbwv8
Zk98Qecwhis13rQs1+toO74W0BF8kYZTrve8vOieDC31ZL+pqgan44yEE38owlgZ
gz9dsuy3i3VZghp86QfHJUB8PZeZ1ApkrH4QUcGWc1vcyYiS0+KwkIs2kszjWK9O
//f3EtaVCPQPPTqCFMmiB34xLuV447khrMIednDiNPcj2oXXJw1tWzP7tFwbLt+X
8cFikVpjW/ocjLKCFtQr9La0SeKBYBJADFcCJDXZ7UzIZdT2glvIgKFd7KPZhMis
OTg+RUdy5OKA9hoBP9bqEb6Pfnv2z2ZvWUJTzJWjPSMjPGfKlhOVcwzZhjLbGdpM
4RLQRhZITP1Dl++Zp9ofB9cHF2ESPSkFNf19UZq3bN135ZIqAhuRgw4ldWExoZNE
YKSCScbVhBzWtdLjE0bOP4/30Y0ypbyYcG8ujZYX/hLHwzvcHjA/en82rnAn/G82
c8sOnfsHIvSk4snGFQyTTEhKTvRK0EsIyNYdnget6lzfICMhPmCNS4raFtvDP2DX
TLRu8kMxBfJl98z2y38PAyaV1BK08+Kw9BMNisZtmB0WvGjT33OvuXKZc7xztqHk
FA73X9Aro9GOAtr5e9LtDLdQsLIA96tF1GxIxpdFpRJub1LwBWRxJ+e+UZstNI9H
XiX4vRLUqRSErsyHfO+AxYEKW3IgdFH5U7WDbOzY18QOvjUtDEaGoDg2VsjUh+6e
Kk9Q7OxGndmXWJ9Q3qbLUG+WDMTmeGUJIavXJ9nYgxeffsX52bGJZlo0i8zkvt5q
/H1xqN/GCCAthKEE+bV5LNiqxMIQuKUinNZ1/FgcYRE7k5yH9I8GepASU/fH8uAn
tQottMiM+bFyUC1osJ0XMkKIhMjDVS3QPLSlUlDebm4+Ne92goAlY93Z1k+mACem
tZrf6bfTXRWU8iGBg+OLUHjz7TK//rktCPnPkyaV8HSeSdCjvTN7ozc7gA/HJxaJ
lk/SqiOR5SMm7R/iFnyzKrhRw1Kn/jVZ9zs2LRRdjG5FpqKpX4UT+7E3Fyzx32UF
9Vg0CIY9Hpf+8CH7vagcuPIVyVHnBx9d9EusvNjUJntkR04gEqmzYFviZY3jdTVF
Rx/7JWCPNtX5DqKrSK3vrC73Uk3dFQbw0fEyMU0JBDBsSC35nfW+TyLUFWJ6vdFY
VtcHkjtQZOSIQ12P04Vfou82W2AyNsrIt/FJIaFDY9+FdoOqtmoQi78Et9E9i1/E
v8UvR6ahcYZKtS7MWDbVgdaCMViIeDH+RlqWlzlpyW5cqgmfL4kmAD8EjKkdmoPK
aEKrWNrzhTkx7MQQUClm6xtmw01/NJjRxWddoYT+I2NwMKv97l6FGfQMRGr90L/Q
tkdJ/KC7ZMY/b0Gp7qcAGiyDCMCYX3oWZcLOuPyp3GUuRpclWGKOyBO2W0ljje6k
1GonEHQ9iJjTcIwNwgNmmIBta48OpNiRP5ofz4pQTBsytEvYCN7p+ePNx5RgnCpH
HY54Ch7Yuh4qWtrjshlPoKtBjiTyc1kZuPJdsXcL9mbiSYHAFlszraLiMaZXfcIR
nVkOBouU7Xy0/a9vIpv62lbLaWEn4wkIVrVsp/6iEKWKE0JOKqjCgqGF0b5xE8E1
3nYVilY1MJUMFTS8wzn2lgTcDJEgL2Z5azL7TxdqPYnM4s7vmUhFmtoYDGhx9ddr
+R/azCuPWXjg5ehWoZMwidziR9fmWmemoWUqucyRVRga/Gqx2wCEgXP8xbA4CTWb
0CHbkrdNQCE02Ts0L2EcFfJWT+nd7N98bwCaAzVYG8nuOlsmrEglfvEEC/VeQIeO
QHc9sCjiZ4Xrr3y3URFOHmryKRVuWtiqP4RcVhZ7BCVMYsZ9cXyViUs94e08XHSv
Y8qIzMCC7iYHMmyTQTd2haRHtpp1lmzmt8bicOA2qnMVEIM9YweYKeNB5w2Yv6qt
MfYoh6v5w7j46XWlYJWAEcN+sGuodRzR8slAhe3lU2uKC+G/EZgDYt2rDUQOGH02
ZYgOsb6sLpAGpzB/vQ4T5ZNIKADMzORHRYkBE30l+zdzjRJFIloM4+bJP/ugddKa
nDLcoJBASlum9JNFPsGoS19SlzQfegdenXApS9ok2jibYs1ZwFko/xtx1zrBgOiQ
UvhtP9JWzp3OZX7TIsBTu54taEB9vbRue7C69cU5D9iTbyxPXWWw23eN4yGMMPmj
oNmGYYbWjZ2UJVYdUG+YEedKZsXs7zQmJ3MgVilNRnYkabfWALDa4GDeBso5i0kG
Z23677AscsszfoaXlOuF4PRPM3YDJvFV3JSBKiZE+aZWhrTYxPIRgWO6ZIe7ENtO
7IxhdQXjRL+9NQNREvxT5qSFJKLyixlNlymXFnscBggc8fnPhAkaaUbCyIEuBK4k
Y+fCN/xmRJ7AGtwSg1kA7pfVInSCtzFBpuaY+93J1nqDmvzwRBzhoSCAUbg9Ng5W
ZMVo7z5mV0f/pqPqttsCYxIF/CeLrGA/cpCg889z4ZtdLZaXQKrUJNU2RELckolR
kVOp/RjpXw7VTCAv6cahpXOMVO+lfDTm3M7zdpfj7iYdBT8O1Q/3CuBT108Jw/Yq
Ose9JvEG7//+dqLe3GbYTCdAAxcpYkMnu0S1obRHHlCQeUHQCrnvlhVozmvI1LEy
rbxcY958+3qdc4JH1sovzUOIyBV3+LUgfojKQ4EM8N0E0lZfa7XziivuC1InWbg7
pRasQDJ6M8f9j4MSBIgGhjON+bMqepDpuxPRT+WAncE57T6iXCNuzvcGK+4PcCb3
iP4v+nLFEJU1nEkHlipyWAttbhtYnXkhA4aoBfJ1Z8FZNIeYfoZdtlGSQJlNL/ni
krBOPNWrZEAJABtB7NMAOlwj/ZNZcL+B9ekcnfvm8rcEPRYl7nkFJwLlqfxwyxdq
tQV+74FpHufJy8FA+FNUFRDBgJp60xpjlLFVCsZxmlXAueRPwts84svhpZZ7Pys0
kjX/T9g+tU4keCu47sOI/RKS4ycFM+ZRvRjDO3yG66R3uIZY/nOqHXSLbHxFTjtJ
eIVlAw7r6TUKGCpV8DMPir4U2UNJ4eSPj7ndOTrCqg1Bf3xgMWbHk3prF3RZz33H
PP8RkJE0Rujf7djyQNeZt9yDz9dZ6wiIy+/RlZVI9p8TGCUpXVvM6YjCKgyjNTzG
V5k9nH9fWC/fP0CmszDz6XrK0qNptqxjf43zWaNYfDatV5YZL7Yhk6KX3uHXvenI
4P/XBO0S+wA6co/PSypnZBwKQGjDYRQo+Q7Zc03VwjCsj0qBfhu3LvhAYHpV2oD0
LgH9X7WRHXUHgWeY7eD7f9KivSlPNg7D4WZkvFvMoRr+YRdOfC1e2fC6BGDdqyt3
Msf8isCoTYVJFdDYb7IGXypQDxnanUW+tNtpPYMcRA+DhmhqFyBvkzPkUt6Xl2xJ
xxli7RiTnVz4f7PLayKuxHFg3MMh6FS+IwfhE9gljwrHkeMJhain/FUBRGQXnNYW
EH9vJgw2kKsDrz7Wiqm9NfnNiQhllbCbkhiXSm2CYwUVtVXTZlsY6aqAYkE6hl9l
gmRDWjvdMiagCvRWJvZmLjfpidRwknhY6x8rrHPZ/1+vSDf4N/TqRIB6HXJyhZKX
bL9ErY7lB+BZrDaTPeIVfwM0T0/S6ZRpx+ENXW658pTFS/pq7+8PFABcSEyfq/Hp
+/YLM06bjHj43ZWKtm+UDvDajvapTOgV4yicTPPEZIIVYbyt2OVTdvmMxMOU3BxB
DnWDw0MWLB6w/1dCiAgc6kd1Lx5Ivc/L9s+PdaLWrghzXzqMY0czK1pWJoW9AyU8
HDkjV/5FFXTToLO9OvfeII5JZlyFxZspkmaZ4W+Kg+qNOa5uXFdHPNLD9plAi/U4
EPzP99ElCVQsv87MbvYkbEjcYs3i2Jy3lfUx6GjmEmx1fK27QHNJpvIuXt+Cepci
x6Kd69IGTk+1V7W8hij7a6klB4UADgB6TG0y0ycea/6bNDiCvF8VQphq+24A/7bK
UyqfVFNo/9j+C8O71eEmfVu+cs7T6OHVdlDKv/xk6uNnf6nwksfqKHnr1s0upFG6
88l52D90J33VBtLnVM6CRR8mA/xCr5nyB0LPWUDjkJAcBL7kOl44wxM+PMsdzpVN
lZt8VRglJ9n5hl52gdSFNIm0aKS2GzLWdYmUMsiuaF2dD8EW+0FXiKSjivS63otk
L7N8/pgGpAs+NRJZ1bj0y0Ts8m2FzfCmXIZoFHkfPCbqEfnAs3nM/GqzASZAuOhK
Hvc9ucZlhqKdVmnoWvoLB2Rd1qgp/8V3IesyL1AmI97llvtm3yz7Ch9B+wJzqWjI
K2NQt2rh+QUMjKfIoTIUovcHgR1s3+jnvOfZYLC85Zf33+f1f4GF656NDFGrkTDP
RnEl3Z4Y86yaqlgdLfFyB+ytJzuw3Tjvp4Iz+CO+ep+SAYsJZMyVO6Qdr5EkYyqm
AgvlWrWhEOVRTR2c46FaDPY7HWYJ0NvV2WQUS4vQW8H4ldCP8Ll2lHV0CiyXN/e7
vac5O0+HHS4P84nWaCz6RR5f7WMDnsjXGt44UxTgpm64D9WueImc8PeSHtUoUBDA
3o11ooxTuc+6oDDFXS740RsaMRc+i7NaF9rLqQxKnDNsG9GV73tnEI009t2k4q7s
0ZLGqXeCDGqz3Tw90U+hoCSsEcsP4gPmQd8bL55dS9rYrt4p66N+CfbYPPiQGeav
6gV1Lr+Mrv+QHlWRNPQIbcf3KA5ge5GbaOBXTSVOYyvln0fYy4BlB3u41o3HGXeb
mDCcxX5e44S0mn5gPD0EJ9NFDin/xCYUfCXaSq0nNIKR0n8EuHlgP9nfgG2pd7d+
EC/XQkTXteEFow6z647tTMiRQyn/9OpDKJ6yQHsO4qJY95BcTDFxayYtDV5GDyJ7
HQ8Ga0g8i+dyda6g0pyy3zkuRR9UvYwKNCvp5XcAgrWW7swC+gyDwsO8UVG7t/1F
K4wzilVjq6XIy8V3kjcAilaGVu7AerRM8zi/uYsLmP1Xh25eCsDYhLRs5P8aWBL9
s0Gs1eT1oDOv6I6mllUTwcBeGVIBKdHrFmSLFnVOzxpql4iofDSE71pP8RuO6/QU
kiGUFh7Zil9AFEHAczrGQTUtBfEuj+Pc0PnSjSLs44cN/9YXiq+Y+4RNipXAtl/G
wGRZXEcJAaWQ81HViju+UT7VFtOE7LSfBvGhL5FMY4IhDtX6Qr+szpzrZhiqjmop
jss2ZqpM0nNdwKjdVwrYM614mb8bJvY0AV3NDs00uTh4bS2is2TexC9yW+8rFc0m
Sv8j+3pIpk2TY9YPsjZz/p6PMk+S/MpWemIJmX9eh7jmLUgiPYmhsHXO7SpEpla7
019VgoTp3HM+pQRN1obQYDMfJwfbzyLTophcLEQ/kC9NJWNzgncZDIrmkfXLmjNg
/h9JcXqshDRGUjbj5CMeN3XosUBBNcumGkwjarm+tqaQmPSV40RY4q4OGQ1uqX0Z
7FWV0oqHr9hot6mtdd09DhNfJsWxhrTFlQy7KBE4ozLN54RQ1j4rgXsIT5pGadv0
+r91IEvdHSbBWQ1KIdFGaKhkZgZiKdhA3F51ZUiewkX48OFGNp5YFO0ozZ45xzDL
N5ceyxRfNwtcvsxflIZa9SgKInTX+XIquvlIBDYtJctEf2eW97VWeTL9xAdmEq72
ZAGJoyCHUvKMwvXyOWfstrPmiBnxiBJ7DfDDxLwCh1KuQArNYGKlg5YwfzzZIsWG
jVsRWFr2R3I0K8yV5LAwM/tWWkwOghpVAhaCZVpXJIMC6Gw9VxwFS03rcXytTuoH
kgrEsnwCiVd/ahJLzZO/RkKCOnyY82GksjR1Jz8Xq97xnjsOuHnR5ua7cv+sFbZ4
emi8l0aJDMLkPHyq5feoqPVDcSQwY8tSQ1TgIiA5yobGN115OCeQ+R8sOkWszluP
H+1zKHt3ylzruWW0jCgiowHIO7lJWgnh2TMaM7K3wbPY3b3C6c1vGhRly2wFb8BF
5sqnOgqD90rh9YUlHpfCSZ9S1Salk4eFq9Px8CBTGLej2bXSkcJ3Z5c6covW2hFO
vnM1fl6l7yG1Jb6Rmq8VdYNQC+Iuwe335sp5LSy8cDOwKipvY5kaDN4Eor5O34rE
Y2dWGDehYzbzFDFEVGPncV3yJh57hn8cFQh9pueoPVnSP4OQ1Anya0hrwIvIITQc
/mH5osqBfHFiJzIFSX/2c8f+NrpCs3U+eC1AjxrdG+BGudh8Nb+enyeUnhtpeIn4
acqGsRgVmqbIIsh72wpIAMlgbCJ+UrWRxKXeRRoLL0E1FAvKdSkt5Wh2aWK3XZFD
YXSZBfWf+ZOTmPiShYXX+BMVEK7tyTU9opwAVw84y1AWH2feS2zFPqqaZ+qKvdxo
dhAhTp2mJ4SO+mO33fWyQCjcP2JxV+uei/N7UjaYmhm88RenX2xa4x1d6nDWEnN4
KkbM3FJpEKSfFjrwT+aqU3qzjop+PutVoKRP5c6VfH90lZV+7U3swCO3MQxFkYBY
ajAcBxVgs71NsjW5ke2UjM+B12TDf5qRnCeYuT2HM12Q2tk1GFEo/kl7v335Evy+
aN0ltmvSOLm7dN1zyxjCN1pSx96QY2SabWI0RXEksozrIAS6NjXba+pmtQE4A7Tt
gAUNfDD+CB3tR8KEG733ryknKzDg6C6TYnX/IWOrCqzILM4gjJyh8nHxTXW9EScG
RV+eO0EceFh2wERdrMz6JlMQypUho4yyKBPltoL/FiPq2j3lvgnr2Ub2BYDmt12z
qGUu4Pr3zS6HRZcFTZ5EDxlA3UKnG4HSSsPGU0T8SzYD3L5l/D2EzLhpq+7D+JNF
meAE59SNuIgivZZoOtNs5zy6xLlZT76FWCA7bWxjqt8BhLziF8a5N8LyYcv/4RQE
lI/W2DQe0p5FvTqBkPiMI3c0MQOzgbm6GsyyEmUNfrNaNs23axqf/WktKsm18eSy
EcbqVDduzCY2W78ixy+b1zDYd9Y3sJlU9/C3E/FaG6QeOECkLAab0++ppVUJCcXo
Rohl5jkkxa1v6tf7VeXKbClESmdNt91d8cFmQs8abg5zgAfJhHG+XgJkukuFbl1b
+wB02D6layX6yh8TTh3VCY8EPNVeG73cl9hWBTTp1Ki6YdL7klJD5BF/YF9hKQE6
ZBE8bcuJbosQoVOnR6se3EBO+WM5Om0E6b9o3lE9aMWAaPi1njeByiL9qd/IW2RJ
sbxLHGKWAsoOw/LeE38L7wwgFu4N01Db1xCRvZ1UyySV001UhdWjcAvAbs0y+wto
tY+oveieS+jOv+UhDEnsCY1gUw+ROpF/KwEfLBcLzOloOahreuHtvMIdkuhIRJaR
Jcf+uQYGPBcO1ie/sQs5IbQW7JQDvdlnZbIPHnxbpRuJLub8pVqKvPOdPDdhovcW
fHfz0/f5yQGPPffd205joM2t6u9uPeSjdE+z0YpuF8lfvgOB26WmVm2PlZeYu8Di
I4rCwHYnS6oWA7ZU9/f+6O3U+anLFO6w6rKKCS31k0lfwX4Ay/kJgxUCwvVDxENc
voaLRcfwyDdkSMsFymaUVHtGBchrubQEkBz1g5BQ0TXwZmL8AQIVFzdZXt2ZPPQs
MKZrTBs++7FSqrLRwK/wCjdRkBldeDJwbc8ru9JCTkGRaaAXYjFA7aQj2YMY7aHl
vB/iPyWjO7s1kTzI52CM3DmJamZxwAQPA1EOdz90Oqexv0Pkrg3Fj6nuOdCDYTHv
j51dMO364OKSY/bn1B/sj4f+hy48q5SZ4jsnmxKoXHaZFnrZL1KQCGQr0AsCFMJA
R9l1XAuiqBm05FiW7FjhAWTEaEs2PAPv38PZZzQYPorc7kv0gu1VsPamya5HKF6+
dTh4xTFogtcSm7YZT6/BApzXkt1SU83UG5/B4PfRyHRXqCCq1dE2IHFMZH/1m3cW
7ngtKTbS2IqtDTZawx1Sa2YY1uXaBqqiybM8g4C1bCbQnNkS8MKHvgzWYYG9dOLQ
DyzdS7BodC67MSNu1xHkc6qBt9cUGK+o4f1wir12o7GXkPUX9S3JdNdlliH/X7n1
P2CSQVdflXydxBmeJFPrb1kgIH57S2PkEkh08wkeaPjC4At0eEP2L4cya84+uB4Q
LfMsV7+0P4BaEFSDP1F6lymyQCeP4TPg6Wxz/gW6PqceYz2L0uwEFQiXAh5kOjhp
eiw9UXGNNN1K4+MyBeMJEotJcOaXbi1taEljGHfM497KxLLtW1R8SXeQgV5ehmcb
RUmcaG2iH3ypL0uPbb0hjE0+OKb0xkIZenVcZcp/d81/K/F6e4SLG0CY82eD/9U3
0o3gS35urWr/hAR5t6HJW72+h5drWZiFxHDuCUGmBFN2kVpbNir2gsw45lVyyacG
9MGOekRX1Z6Z7/jDFpDZrjWfamw1IoB/yO0TFu0xm+fIOO+oBePF7ckCtmYNrnSL
YQGs74RTpssym9eEOuZxKmFq3OF/Y8P3ZcVjg7O2hALTP25YIOFZEupYBG4Ai0W7
xfGoSTAbihHjTX/K5JywbfODst040yToxF2Foal9lUun/WCARknjAdhkg1jsOHkr
voNFA21FwJB9AnJL7o2Phc2wzXrfEX4H+HfuoU3rl4Z1SyqzWdyzBb+yb7QnvjNg
Wr1sjEBYBWMwipPpz/BBz+Z6oVi5eYybrLQpF05YoToHteHrkJ5OolGBN8Z4jF5d
ihjVvtnkoEdOpkkeRCWlzMIzLqniaGuNoIWqmBR8Wb4kPUA2ny4yzHvQuHVwqRLn
ISefNx+46jjceN5rz9+il2X5lqW/gmfr1FHK6Rf5E6SwUTnEl5jWjQ51yP1W0/BV
opxL7SW5GVpbpeDM3wLsYr18EjIa0ueNXq58NqtcSYt98PMWfnjuKQvGPqQdli2X
kVthUXvK7tZ48rBRupGhaOpe4v471RdxiUcLlR2UN69LFFPr+cf5UVkZvv3et18p
ziD4e9zDRsPZWM7TF2PX7ryXkLOLB+aVUI9PjQlt/7mbXMSgnVabGqVQU1VKTv6y
EGXWJjF5Jd4NFO9qdp7SZThwgH0jyM7mb1+OuldZZE+RR9HHISsNnt4wW4BZxboI
FHGFtMqKs6ztcpNiq0npyQbxeD/LeE/hoEz8zgYSJ1S928LQyvqNsqjcBHFxzMC1
nCzUq+gKONiayfFZvz9PpUIJqZ7OqsOO7T4Jgn7EJJkdxx/5SIOQsM7wQzkjRCW7
0vufMzhhIlt4Y01FGLRidjARfBozuuy6DBrN3++quF2Sv/yxuty5T4kPavawaIAa
fUCEYf4ZTm07xQWvMivRd6MSKLKIC8o9L6f85gokuroKUlEazq2MLew+6apOLjZh
Z9ogK2kbTX1APha4VUGuUK8k+E+sw3v+6dftGG0cN/roKupfL7brDvnbm4ki/7Xz
kNDtF8bw7NbVIE4tRTs2WETRbr6oZze0sEX/I2AlucEzAqN7KdjrZbcohy5jsy0b
6k/UL4q2uW+gER1mVBDr1eBFjO2dSuzm8Y3voREy84HbR6BAmL6fM9nLabZn9DbZ
PN6jyyQ8kYUyeUjPKpdr+xVJgHewFtJqZfgYhOue2+GnsCrMECCU9be5/w4CsmkM
3H1iPCrz2smvJ4hDEEPLt+prAUDfA9uSw6rSjYNEz7oV0cXII6w2XbJYl+VSaFRx
7fskTLkvuJ+Qp2UbmhCU2VH7b4H0MvXYr0hnvm3jHn2k/AruJRaA88auCf9FDmRM
nysIgjXbTSx/hxWsZ1NECLhVfednbcMxDNSYNMu2MZVslY/iXFFr2kylU8fCv9sD
JNh3RDzC0eu4BiQCYikJXbhQhG7iHU/rEPJN3QbOGgIuBr7EMWawW45la8SoL/VJ
rE5w89uqfeKHlpXvjhoFQOnQp01fblXc3G3dgQ2UPJ8btYwdYGDPIQCK/J97ko1o
npfNeVYbMFEW4XaM7zlK6COPb513SUGx63GK4Drd3/q9BXX+2WgVfIlTGhVl3Zgo
qbL8YDCgfUY1Dx+L6wsuff4hhgAPCJguHSGH5Nz9RcZV550Umg61lPJYWDyQ82ay
jxEBH3KxNj5S7x2zHKPZl7UxK8RsBk+XDvk41wQyW678zaWZzEDsCM/7wUfyTMfn
UEwEQUIEMPkFAGMX4Xv1l4DhZV4E/bRYDmlIBuRkndWV0GkR1TyG2Xd/RmfLi07M
DH/L9rhRvYCbu6sRjpP4kG7mgzi61fOEcrEROLoqoLuWTJKjojVK8fQc+VoX915G
TF/zGYAN1JbIv+KArhBhC5LCm1slGnE0Nw02lXsnTbosmkzdyCFMLiwswyeTIWNd
EHKcQbzJtH/hrG74jEh/nbDmAEnEr6G1H3P3mJqKRgOlEsA0Ey/SyQH6AUz04Acg
VxEdZp2JiYYhVE74UTWuOk4lDc2qLr+z+s8nSnoZajrceSFL8vtnvztZjCyphs9P
GVmnX3QuVTRCdRUij6N6oLelR2YXcyfi5usQDPawy7H1WWB1evVVosgTXdvWIFfe
YZqISWFWsZ7Yb1erqgH6sMwW6BkzvFoIOO6/DmtvApNDgiEUKyKdTdPVIGGDG22x
g2Y9psDTyz8j4DIbH8a+IPZZ6IYHpvJty5AYSyFjca6F6AordrTCq2aei8/NxFcx
dWdpFLHkY2APdQYQXTx/Bwm7vUL119K/hoLpw9y9aJirjnEzglVpBj0h/cGxCeD2
fKY6yhocuccZ/8xK9XTupDNZ/iGT5XzId2nc/d2VvCMMUh5O6lH8fzvg0j/uCHmx
Fke7kK89noZg5dK/HpzlTabV0YGR1eUVDPki7Flnc+6t3M06FNvksLiKiPbioRPu
M/ieXM2cySAPC9z1UcXFceendJGu/j7KdybSm/gImPCVvYaxiopjUWVtlYBcL2KF
RLZp6zrPinYBp3RiB0Lv+P6QI0uOBOAVgXiTXCRcSbFFP3lzBO5diy5cTKx9h0lO
wkqe10v836akaBVbK0x4cSvtRnZ2BXgs2vK79UdoFoW5BDqdEScZOsm2v4wwANyi
6o+9wRgbJre/M/P0OsEdRJb5KJ3608xBYS5oR/GMUjuEAIKJvtF8jXBzqBgJ17Ee
toXl1u13iL4H1T10w8/h2KCSCr/AMIzCXp+WUBLdtGV9SaIhMNJYdHpBzYvyUX3g
RugyZ6EV8ReS7D8fivI0PSSmMYrhIFsQmkukSAnKaiaxF7Lb5WvvYh9u3daH8fRy
/zYQT+sxGmIDas33gK5SBGoou0sz+hb+xQQVsaFT4OYIDgt4cebLqNGtwCQckXVj
6Fu8Bc/mLAvbPYurEyEP88h1aWgOo/WEnkYOmVYh2LEjoVMngyyLiAoEf0hcdzNB
j3rhxP/KGJP51UmYokpcmG//bwPUKQ3nQi7a+eRJjNBdK6QvJNKnyhqDdyRbnfm6
XJ38VrlE225Ovrief5MVO+5bWIBXPn8z6B0GhmT+RHAPKGOYFPRLc9J8Pk01nHS8
wMB1ldvd4nk3gPJ1s/5jakylHVsMk5UoZRrpHZjmObSYYSkDPrWN/S3xDaUkJ23I
UJPc85p+rBWCOtuqgG9BVMDAVvnNJewr+5Tjfntgn6uKGypFBmTzf8VsgUUCk2QL
QJ7MBdWz72VdQMitn67HZZJ7GRx7bYBLpDJ0xJabkvOqb2yDs49+/mv/HcUOUPM4
D0uo2gpn8IFj48R8Xa5xopfNI+bVVw82fuJgmm2iy78lZp143QN7V4/sSyQVpRMy
fhhRCMSnRy+86COX+pni5zLCMCiE2mlmo11EU2Yz2S7RpiQYlLVHUCZuzUwYEbaI
GNblqYS8z8YTepzt0lq1Uiq/aozd8Ido2g1ayMLfz0vToTvMoApOsH5SQWlX9own
/RgZ7rxTxIwp0kkgCIwISFGs0OMpOnjSYOoxZoOW2oRoW2Ak/m5TRh8YmTCmPWLy
m4GjbS7JUk64Wn0V/mWfP4A0y84LDHV9Lf1MCLfwFlrUMW1BVdIqkzne+B61a13A
ZygUZsszKbaVK0rhX3PQnm9ZJfosK7Nm45UQK0Sybj9s4X26XbggY0sV87FEPxwZ
zMTGc3xztCqkKEFBqN/DfiQRiEymISYDGM2kx9QyDqXQANOXrY3yshv0+1zvehCZ
L+NYceVGD284VSbapeOoeRX51X3AzeX/NXEfUgyZlbuI+Otn/L0Vrg+tl+WOruqy
EKqB7v2YI+kZpO5b8DBTxrNbdwlPm2CJSkWqMBJSIVqnqHs3pmTrODWYuzHck6Hq
+fyT5BKlEt13pOSbtdK6psK1fuOsDtIqm/Al24vAc3qsY8EPnqrAQOWFg+FZ1v9J
eMoyPQoD4Dbjeab+jVFUS9VDySzwYZP4EcqVdzDy6lN4lsidumxmKnb3Rm5s102A
7tlS4122iBODik7NB1E3uLf+NRBJoeUIqkJn0aYOC0hMwMl8dNDI4efnwn/N7Bhc
NFjq2P5pQEo8kVFLWmn+X5wPJSLPPmijDmWSUbK7/zT6+VrXk9PoE6OESI8fH6qb
oAku0S60GjOgOypcDz3Xt9LYGvD7uuH/KguGZOOzjsdvygKeTeH8j41Nyu4mkjII
cn3LYY5i89AvRfuNzFB67odNn6vfrZmTXjHQa+7NMcg+RF4XJmUxrvpbicjrsB9M
vG+pCD6+FDXWW00JJG3itZ+UY9n2/sd/jAN9lKwhQWlS3E+rwAVQN8wqK1JlApE3
mnH5TPX7WzXDC591YHPwwDnP7tMD9ADF/riV4qUxDvHKxvoy7T62nAP+RzCpWqUS
HL0b6uHtz7jeqAVTGJ1spDNvejOo0okjZ8rTO1O1wMqVNDFYHElwpWLwosGhUCmy
ZrT2ogRuX8JfeVAbipu/x9UpHPW7pQRnmyJ8I6dduHi9BtME4PiBN1xmAfI2mJrt
YR8WuuhnKYiBTqNacuhWo5x73tH31y9F7fHBgrtBKTgmIMHpdH7edvE6+QNa7fMR
w9N7Lz+3yuFi6SV/OCu/GAFwCoR4AHLejlkkkDxpur8LIrkp+ih3+lX5OZfFavWl
vwSuIOgQTve5DG3TcwRSYbPkyuEoJLpoPaXGj9b8jZ1vMC43HMOoplr6T1fwbXFU
SqLkwvc8SYxylu7UlVdcABThkO1J1zgTxj/6NscJvlrC5UlUFKFFC/W6lelwhpKK
TJzFyZfu3dOQNwIxDJoI+DI5i/ifaxfDQNf5oJG+EWo1i+mT4Fi5D+0ubXJszhT4
99sGHDhj+HEN9k4e9+0NPU2IEbK0/WB97moH3RUM7ze4f7mxp/ndAGYT4W75MRpU
RwLjRRm6boSFR95IkeKzy4Dg4AMSChe2SHYVrumw+r7/vrmYPLJQtVnIVoCLSnVs
5+atnm86FRHrWkLhnIaLAtGxvDFUaRvrG86nla/Juc1aV4E6qCIQCYbmjcma9/Tb
zi+mBk7NsRH5/HieeydA6/tNlM4usJ8+WDjz/aFjjL/3XnpVjeoBYO69kRnPBMmv
Q2qiCgLaICjSAuRwPWEhMJZMilSWIa1NxC7RJPw6dDvU69Yo8byZE8PInfenRWGv
+582HqC3PLWnZUceWHBqNHnXAl1bmLL5i48A0I9lWKin5ZKK3TtKmSkuRSxn/273
Bbj7NyUR/oakTEwPpz9Grnm2XxF7UiX7G8f5sSYRy0CLyxZE5YZAuq4E17/nlJ33
cZbD7c6axzNUGoqSgx/dZQq7MbCK7pTieR3NLxntnX7RsBFOxpQAKQ0q+3iQZN++
9xg/Ipqknj+7U8R+nV2HOc7Y0vLBI75WmHZ0HNJ6xEFobAHKvOkLQdDHjHGsk5Xa
5xethhuyiWphK3yKgr9nYXklXuibXNwC+0WDx1++URZ6nJGTi0jXMatWV8MeIlxG
WbAit/Pt50iUhNHvYEUwxr8nJZ1oUdFW6AbNNshtTgDC/MmufnHDuE14wTrJl1Z5
/EO1lfENdAuHqz+uOfSqg9u3wFAemXHEgU4zbo8SwGRtsqKzhBu/Rp2BgI4invdh
1hcRHAYvT2hRZRPzXuJ8igi/rgk/Ii5fZINWzyfk937GyxjBti1EK08sV0RqDNo3
NPzGzuNqC72qaCqUS7b2gmp8OZXZGcT8qrOc7wZNlhBjt9nUDXRIsYbu9KQiMobZ
jrDq74Puk7Il75OknJqNpW0YoqxV6p0ACySQQPmo7Jx26e8CjOwmPdvGZ3oAZsYU
JqShiUYs8CBRC1/CaUXZnUav0OJjBD5wBcUKBb0oDIZ26DU3B9Ec2y4fH6lfI3NS
LAA2KKVrCZKuvVkUqiK+DnHhbKDJBqcgtlQWedUTcZijLA+fIPIAUsnMzwPIrNzB
prV4gTz/pyXUUNfrFz3jgBfC8KPBT6B842Wk2lTKH2zsPzAtUYImNXaS9NcETu1p
AAL3iusty6YajQNEqRgsc642a3GSkt0lFzBUSOA7BegPiWW4K3izwIH/1MxDmV53
FkTcCqeKovr/Cv/fjZr489LHAO8omogmrnnKuaZrOBZWn1Xn0pUDITmWbuXID5ja
+tddJk9t28N31Bru8AtuHpBjx9fvo+qQCsEXl0XytpNf2U/RPExNNbLaH+78Spe7
EO73QG8qwgB1bu/tLxq69hGRwrH3BXzoM+d9vnAL9wOGN0HsQyoS/Wte/uJEj9q5
6CpFyBjjDgFjkeg5JLDwI0CqwR805iTYE0+P+QwTpkPeBtWZP8U39wa1mGxtqIwB
Vy48feYh22X2lpOg6NehLKZpFI2Euvv2uEnwRq8HNCZO+Zj0ItKm0nbFnTUt2lnc
4f0ocKv5EkpXmEp43l8Vs4t4mCgYN6HJIU4BmM8ejv65kTvjD5IQijA0bVWwN++v
PDHDstfeNr7THO4tppNUihM01uiIOWlj3bzm2NbglBC5TIkgUTZfewP7mDpgWHW8
OH2S67pm5MQ5ggbOaMGUNBEraPlgF0imo3U1ng40teGdFO38hudf54qIvVsololR
78DsNYbqyZtJtYx9hsOAXK1/UpIi3ygckqaJsL9voJAdsJTc+2YbWiYXd1K9RAv9
vl1fMp5fOmziYi5HEj2POfPbnaroB32Bi5uRkFY+l+3DXaIlqevrO1UL4hQFcbku
QdKmQBm9F2egXVmpaE3gstemqRBHS+ZlOCuSVBN4ZTH8XWoi9BKvQcW6A/5C534z
eLcYcajn1aphUXaMAX48iorQskWxVcnj+CIgtJjGvgL3J6QM5mnoZtcv9Y5iF2K+
Q9Cz71NnKZXFzXgxojj5QmCucWhwlLNnqRa88GbKIgm7jAlmV9uX5nY2qGWsqfZp
YjzdgaIKsK9eStc/L59cTBWpav+BmffNq8iQuCfuDFVueMrhsuCjSWS0RLnB83lG
dLdeDny9jrgVX+eQg0c/hgoUPCItkHx+3Y9xMv6W0WNcCnCR1Y/IvaGlz8STiwiB
0aIN9m7RXgjgiLKkjsPc+t1qbWN6l7/yQWxOoW4jjzJOt+1egqgh/8YagJgnBTUB
U754RPZxiUSAAeSaZ+49QZJQWVc24IFVyGeu4OukUntrNJxihYtkXFssXtDrzRxj
lj9ORXGf1rEbjWeGTf5brdKW6pc0U6uG/8WJXkHP1knf31Ya7/yiQlDx3LprQCNw
PyycTEMisVuxMK8F6BwB6C+DOMEjGj06Bg41Ax5WUanMdPnOWoC99HjAMwu5QRZD
c4Ep5+jilZ39FmUD/0egkVLCPlKkyNv3dxV/KYf5WQYNH6Yev3O+BdXzAHHF0qNO
v/FibDLZxmlQmXUMN6hbpI9Op7dZhORB2JSpoJ5lSO7BC6U9URPFfm64GHGwWv5p
LvRmBfCPP8LRKxtE4/umZM7ydz/pLEeeEmHJtkPE3T5prD0RsM2qMeJJtaZs2Lwe
uBDwU+zMhzZCPzRDCaEF4rn2bzNB+Otx7TjaYAFVAfogmYm2e5HQMO4CwsPYYIqI
ksv9fENniliuRAvzn2NyAmihRMjOzWp4sqUYNargO4db/bmNJfJGWmG/R05t4qXt
9BVng2HWDRq/wwCZIzLst3mXodze300wBNhddgqCYqAs1Qedoi41mhD5pIFhiKG5
wjBkEBzaaV/YYKb/OKGLGhYjxsB00qL/hQ1B4nYy3P/wle1O0unKTw5ZGgajLCRR
4Qix35I1ocwoV8lshrGwvvGpNAM3wWmcAEfwjjoTIBshpzsWsT8rUYwjqrfreexW
1P6fp58qqbdMLfNYuDgO8zwXRmIPaGlzrMdywPAgSx34Zs2/mrbT2YeoQxRvi2Bp
zEbteG2O5W4595uIyz66o7ZXjkC9id9KgpFTmcclry29vVzJwFoVxyVHloXqqKOy
tL7K7K6QO461wDthuhBnb5e4eNM9SDRqZcK/73IvZsfKGc7Tp7m77Fyuv6ZtyT7W
GZZ23nrFtI4p7X7YpruDCKopomVWsw1J3G3PJFc5bYCsA2E2s1eb2ymLeo+aUtPK
N/at17qJXF/kASvnM/1wGO/nEWPrZVtiU7LgSZnh3qa4F9Jvgo6KvTCsIuy5lGDQ
J9eisPPkmwCtvNSnkASk7GNpiQNUC03tuw1C3G2sXyvGdF26ioAzclYS8xyRGb9T
u05hFQhQzkZ/D6kOL2gSkJkAUElWQ1eS3jyRGrgMLI47FVZkc8e7zowrnWBrEnAJ
n8YTETVKGJHdQ1QzEPKvGhMowm/VOICCBEwEDs5hMuG+n3hVRMvpqgC3YFk2uqiJ
LwgSZCwwtPT/NfPZ0RF31Tya0jXHGmnI1DPiFi824gkBUcfuXk6yVlxaibcvMh35
Vx+NAiPf1NJNJv4rSPQb918gv7+hUcRpmoNijcaeJy1AERJaQZVno9WBKOZvVDPq
+6Ch7Ea/6yOetxlzyd65ig+TNdBXypXFjQdAH7wCG9U+6AtaVbzxKrNpPPB2hcHr
ZMlbRzMWq2lmbM/2yIUio0i6FCe6rVLPmpc+acPd5XrGAnCh/lPVWYqT3tl/CdYJ
dgxdnzqnd1OObEWxO48xuI7n+/ooRP0411WTCr4sTtJMGLsUDmmJA4HxAYoCit5u
Gy1O9imCZ+thfSCyU11nQprOpr+Tz5mQnxH+dspFmM+KBcBNg0kwVDJWUJtcg3dC
LbfGuSVbPlzkZUDyD9VDwjhR/PSCRlQEv9lfnBfUoS/5StsoQ3WDEq7BBrgwjvTv
0STtXkitpg2sBXeKdIzR59fMRt8k9Kobcbpo7W2lxvfYj36jkjptbdSpTRE8y2vk
yJA8rbX47XDL8BPfH89WNHhiIQaVm2c0FQiwHmyAYrG6GGCbcroNnfueD+Dwp+Mq
HvzD55On3VG5QEMPtjTqlopyzr/qCvRsVF2zuezyJiQr6a7eyWaFvHtDybwJ8EHd
JPkmfkZzyHgmi7jZ8nrY+o9YxXbNW0svxNlSIYkFOVE8GlPucSq7t09LFVWdt4bp
FM/gPaRtc1zjeydu89lkDbAU5sLqVrVd5pPstRgL/h21wd76T3mIjcu59T+nxvsn
NiHUDGtknCtzWfiFvOI+VjRSBMSaHE/N0EYRJsbS7FZUsazkKl38wO34V6j6iRIw
8PSgaKYTvhldehJ8ed1wylNkNF0KhTPV4RCOeCkUiyaEZoDQk5Saamqy0eCFdD9p
M08+I+5HgH5lNqKAFRnRMu8tbMxeY+nIQz7cpXjT9aay8cIlU9FH6OdyDpBogXKM
PCZxM/m3UwI7CO0fI4s1GsrKydwqtpmLyGPUu2CmNBx+vUOdLuBfer/sAvPwz2UN
RdrjVPMiqOxi3r/UiWhqvWTFij5IPEhOwkw9dIjCSBGVAT9cdtwsqUd/gr5W7udg
YUBWUq3mVt1LWq1AyFiLvZLfMxQmyx7B8nPoPJaGVWkWYEBY8RlIpFbx53H9vS67
d7PpmTHV9JeIFfoxtXxf1+a4H3EyuXn54uAqVBC0TeF1Da5Tfm3RqQ/465EO0GYc
mBELJib0YCvn5uI4yBb+t9ctzehkLy/Zi/VuvwigXye1NH1D1vE8QYYk30ySfJwy
XBRxUxjkBDmS2sviu+Msz3MzbIQpOEc15kDVUL52SBXswFFtyaTUFDyX1hYr6u1r
nz4Qct8wejqyFT0woUUkESPZ/fdOFsoHJnkCAGFK0wTgxS+Cwc23MvVvPlxNbpkm
hoezX6xbxvL4ocico8fCyz9k+AEIsKT6q/f8EKIGkrqWem7lDYAnlVQmpVU7dnoB
AcXCWdc/rsKpRGGZuxABoinncNpbpAZ5bOIft6o3zuVkrhIOG86WCcQAbGVIdN8N
9TpydmEAvQGpiU1p26kysqPgOSSBrC2IrrMry02aAgyWiEaO+DfK8ALYO0kJVFoZ
IdOiTwrituiTL9vk9ZmeUQViyMGME3EfMGaLvppU3s48XHEUu4aHCehzGZd5ZEPG
AfsA0iLTQcVFeJl40yObPGvikGM6ymFL78ligVo/mkiuKepHeTroy0npN6vGGpzb
2Pl2GQ0/0FNsBgbqxIXKHL6KwWKpanKFKiVxHiYH5g9FjEUmO3IfjZRftxddNAIY
SFKU5znOOVVC+WHZ/f84fIP3nT6GaHgP9zTkAJ3pvCMp0QpzaANMf0ZyGBMjIZj5
MblxmOJ/8KLOLH2CvyFmdIyD/0ToecU7RFrNjIzB70ulb/Wyc8ougcZjKvysQwEg
zWRV7I5knRz8XvLMPPjNQ6x0F7ROIZLPo7C4qZBqma7Kcn4Qx2NUwJdO3xfupaYq
Ig1o7FDLIqIq5p34Hu6gmQR5ecDkZR8BGCrb0cvpq3itA4eFqT6/wpn+j79Zs7TV
VYupDP6NOQyDDqukwj6fPhTdsjbuBx2oAw1q+WUQ6sAX+jnpQTtFJ88k6hhp8jW1
N8E1GRQcEdt2OT6zArGybYE0Y0CvLitgw6Wl73wTSbt3wNyZu6ZsLtTXL3LEa830
4BfakNTMPHj5wok7edCwksQY8hBHBXoFBXOu8lBjdVbBTAtF5rP2ojdJH6zqz4qN
oRI3X0RL31dTn7hcxq2ha6BQTD+XLJnIuExt1RU3y6kB9wk6O17c8S9+id0o1uCJ
JT0xjl+q7FxSjlx0g7mRGD06vCAhqST0j8nHQieLSoJw37M3CaQ/+vXatfbevIDl
pbxZnNTjUGXIuO8ZWnpHlBjIWGXLEcNnZ3Unr7HOIdtTfVV8WTQqze7IaqfQ8Dv5
RhMhy9wsicC1kCtkL3oG4+/EgyV6Zri2y465oHKqMZy3+JFMESl505xZHlTeP4if
lWBOgv3EiBIVgfCbvrXbE+qyiXDxszq2YoYR+xpYUVlYzy1o8dJvbijjqjwK7tfo
nUvEDxKHy2EaX2qzwXvQF28pzXBeYbRBCy1I3pTehDtUOuPsUMXQscDBXelIZD4a
5s/ekMFHOTYnRYEUk91IjT6aeU1h4ISc+9mTjc5sElfmKfelrnhoxOOS6WGebeaJ
LLbOUTDln/1c+NC+EL9s/5KXYbRDlLXhUCXDf08Y2xhiDXHK9C07OgDBkAh/edqV
tGiC32nZIZ0JhcrUJ6NUNVVMODFwXl1cA+ocgHuIFmbiCc7stTyJlzoor+pI/J7X
vUlaxo8epHH2n1hsr6ftHWSGzHx0pn5QQ1X/Fct4Glr4UM6XEmcZeWcRKOfctrXS
1Kp3gFatE0Sgkor9vnyWFJNpizTRI1d/I4PDRxnyArs4vCJ9BCQbsbIPwEFWzHyO
qJyxm6VD6zFPTtSWhksNFJuxtdTcejZ4QXGUQkl1UqKurk7PTY7YRhEVYz4MoUdF
6lN2y4N3kuQop3lV4lHhAaZs7KVL/9lmG8ip8LMH0k1E7ZGGc1+erPN+SrbP1z8a
fyybWfGO1qcPYUEg7xZ8VHYhoIU3K1snC19rd6Jxhefv1i9FhLqN2iScGNcCcebh
0g+L8Qe64CjfslTvvlLod0x+cuDcuTQaARm2N+wAx8gQNH0SR+2lGIA2L0jWaFYf
TQTgig1b+YNW3pOaGVL2tQcX8RsmtmPYLI5g6nVC1YQJVp7bpsGk6Rxv888q76fv
ZFGXn8aZZSNwFpPZOcIfqS41hl+ZMqy5b4yfW9Pb+Q35xWFc+nWSgWgLuOxKL1xs
Nc7nJ24EXJ6izqDj7HDLYASHzIxXfOh4NIwsEh5y4amZZ7guFYwSiMSHqGaCzs1d
jBQMGs44mtvcXXev+fc4ySfjgT2RWvYYRpxdYaqupkW0KbdEnW0IW/oAPR4DTAXV
upopY6aUG7ZzZ92eQ3CYB7kQbNd2OC/7UZO5SrhGW98fqXZfmbUEzMTYnJOI+c0p
XRj38JQ90HQr8Ck53YqNvYn/lDCkPzBwp0YBLgxAhi7GQKiomSrJaBD1fAXA0KKA
eXtl3ZudJMR/RDAz2Rt05O0AmBV8xJftKn9Uxu1CEc/rj7JMuf98e2AfPeXe05PU
4EfpqnkhR8DzBZV7z1Lyef5+OaXX5c6HTFPQ0cr4gTrxL12fIIpncZWFU10GEcj+
/msAeJOK8y/LbpC6qiGT4jC6ruTxayOYrG1Y+ZVWg7PO9b4pI90wP0E/Ywhr4ap/
wpm0trCZTj8PGNqCPysZZ8uMQicFA/tygpi4yUIiWbbuCxIskOpVb5s2+cXtqbKY
Gw2oCwAamE/h3Ek6GwwMfDfXkZl2Nigctzr9ldVyNYS+tbMvvCmhjl/9O7cSyGzE
Ecph9LBMHFAOQELITVYShBaJptb2ryt5w4/pUPIhqkfa/7Ay/F1DvOxxaogtAaHi
M2KdBnVHs8Ef3HExkDaxjKCoPBDeBxVXyb4+toCu4g12injU3qrijzdcFBBzm47g
0OsMg9o/NzS8p6BpQeXM2v85YogNHqqPTWy+v7e5phRl6PrctlfbOYyx3fq8VV2J
kE9N4Dcq02KVaGsPKYGO3XjAs1NA4hRo5n5+4NyHr9sL208Mh/h1deDGYL2Qsnmg
t3NCEeJeKiPJ31ghHooNnqfdVq5lYTof/m2G+tfR4JDRKyGqwg8nXyq3ZOJHEoz/
eEjIwvIFKC2QN/KljQ6zD173sdP3CfSsKM9vET9VUx7GbnEcchHlvnWn/ZEUjp33
Rk+kMc2pLxInXkd7omv68Z98ksND18BrQV8zyZHllXnPG3hcst53vPczEIjp7Pib
fQqaTG9DZPiwr+tnzS3+8ZJ6C5/N8gxqDKhhc+QaEvXA4CyEtSTl2U0PA4Pmz8T7
PlAQSA9kTMJY7xXhiwmJY0idPixfP0e753I1HkRh2bdNIhO9oZhcLoSOqfqNgl1P
RZlYi46uVWlDz3Z1K+b0keKdUIW8ZrquRuxa9WFSuiVPhCsTgwBrBvasHyyi2cUm
G6H66doloF+xem4wrZkoMK1ORNXTDRsHvAT5QpPFp6WHc9ZRvZ9GmZyUeVzRiKLQ
FLO9t5TGv6cD09FtZf3Glv7A1dgZfUkuq0aSTgAEkgDw5gRyaxjDt8hFxSHP+BgR
vpVcpiYcXEGwl++ciijlZGJOr28GzZtn34p9LWk3OzWVVK1dCuu6QgbYLLTaWogZ
YCUPNs0/oXmmxIyhRSK8yIJoJAhBnJp+QopD/RjYltFFoUZww7RmjjPTAk8toYje
IFpFPWXNzGevXWiKDKKWwcQ8yp+QO6zO++ZdhtWotDBZ3CzJuf8LZ/CIDdCZGpUc
Q9lo+P91V2NyUVM5kjMyuCZDNyF1vO+0hsUT2vmfv9DOM5o5YyoWgrckmoloxw61
FROqHPmIdat60vF0RASDjUCEVYP7NhXt1TgUyZen1DfWZkLf9QLpizOAHwyX5gGc
+huNeP6ua6BdppkGpS8CyigLV3Wk5qubXjv9r5DPhRimPAIQe1zDx5h2uL3pXx+F
Lek4rwP7+QsKkXeil1pGEG9Tx9svGAiP+UJAXrsBtNbWbQ7jYokuc82oWsYEOBn4
vqiAcR5KieCP5MRumitJ9GucELnYziKqEJ5yk3TzM/IH8QanDLwEQfAlYxr3xIhx
VnqfjBcog6Ac8I4h43zcugiQE+0t2oo6Cgc0k8UyPTzkGZY4Nl8/p1+6MW2Cv3P0
XHp6/ysgK6NCBYojC8a6vBYl3K1QDcHJ+kfo24dM6osWR+InHMozd6p1yTBC/9y+
7gwDpIUAwGLRVOcq7thBbzvZlioJ1buHYmB4mMTBOv/JBKSWeKecCsawliiVD1OV
35d2y6WAzqSrmBq2Ywo54IkRbaQex7gg17EMOyftdkIJjzGiI0VWiXEJkOFW2z9u
yI9YF4Y7NUpLlybEV707Yq+dcqAGhkwawJlelD7mPFI+7XvxetUgR8iE2g8tTubJ
HnH9UU3FltmdfTIxxmcQTJ/h2TI9vom/8Me2KDPbre7ZN9Xi39EF7CrrcIzH1Fqw
d65HC2yfS9j6iL/1EzaTX7mnLKTPMCxeaU/La7q8UcUNWwKup0ec76gPJ4B0Ev4V
pcUdLzKDHX7xNjs8TpHSVDuZbxjBa6oo5XxRmWGWlnP1UFA+nxVdjq8c972oukVY
PpfIKkBJkmD0NvMtqzAhW3StziPXLmgcNr4WCAR04LcjXahVWTPUMdYtfMx59iLt
eTq9UiZ/LXJEaA4Hb9/Xcfz4T7Wr8kxPzGWrG7T5jEQepZwHkAH2TLnaXaYrOjVL
VxygFivhnLDzEsS3C3d+k/wtFKQa04gC0fpMJzEUswqP9zObbf0QRCWKQSMt3ymL
Ai/naIpbFDau070tD0Pt7iyJmWPb4Ld+5ZSzVaONRfPKRLy8sPwU3eYJq8XcVPGR
uTKa29sSe1XIo1dOyT3k2dgphVUt30rDvDJSH78TVr5rI8tmTKcY1z2jg2lcnVFF
57j6PZ4GorjxbpV3PnB86dMP7jYnCc2MBjycSy+R0TmVRGdEFbq5w995tVZuN7+h
r9h8Gw8cA0fPP8me04xBgHTRKA1cAdFglTQv7W3pb6tgkmipVZ8Tb+nbSpoLKzCn
rU6GuOsotMNUwMBIJJHkKBXn24StPWjY2K6uvjUZOITOaLuZMapKilOZOJaxDiZL
SiahUBXaiLV1KFdHLm+kVamL1nsLoaSs8iKYl11LFY/1TDZ8opqw6u8LyyYFHOvP
XZ9eudleZf3cMSYIO83Yxx+za0NE/+g7o8RTRJoH7dpiptj6b90MrCT2lFLjslPW
c5asO1NBrb2Gq9pRka96KaJC6zaGTTFuKS7TRqLbehIKQOQliyYEV/jgtmAaEqco
zd+DJAM4dcAZvHCBMAbLshdDAfeo+j63fsMvJPb5mhs3Wf5pOmB62p+OVnf4S4ic
n4ZX3/rTfqtXqAX+xzsJYOUPHL9RG+yAvCgJVpVCI6UoosvCUiA3D8NWyfuS+mtg
wrhuKUGvCJvt64aH+9hCmEBozTkIVoB5Np1lVglcyC7oF8FHGIcR2sIArSPHM8kf
N3cKbYeTLc87ua0OaD0mVl7PJ+yjeHstzjs6JRG07i8AlILwskkHJWgHj9jfwuXL
4aNvo8DLIjpFd6XWSSkR1DtfkRph76XnLCx6e27T+KmOm5L6xfQKqBeQg6EbTlIp
80oLbVt+kJtwSBo2w6LOmc6XFaiTBj2A9EvCA1jhFbVphbTjdZ9EXAy9w0kko0LX
IYgdtD4kt/B1Tvxi1gDoE7+F8GN1wF6BtcbKtZAj2HuRlbOEyid/Feg+dv/Ao85Y
rK8aJP02qtQT29LedKpl/UdXoTa8RIACcpf8/geITa7x6cKWouWzMCyow9laqcww
P4ndyoozNryOs1F8m4diqC9BMR72BGwP9KvdIoyWE3x7iHjnewsdyHav+txYpxf4
yPrrBhj9MvesPgHT71oT2LgfRDUYytj7qBNYT/MJeG5UmaAGaqtXHqLD1oO85UA1
fP81P+M7ni5Oa/zg9/cSxosAaR4hbTghijvGd5QDZasE8nue/OSSAU7E5XkIBgbJ
9rZClscNZ9iaTuDu5xiDUb3q2G1L5SFTAh+geZFiTJejFrq9ESgrByZ9ib1e5NYD
uLilLt+x01BNugtDmvaAFVuoPH6tvFX759/GN1PTXlQIqDCR4MVQVnGRgVEEfxV/
PdeboSB97AAzScaIf5sie4W3oWlrLzZCRT9oXvhnsC93kRAs/42eYyeAnjJUoHzR
cWMzMJfXgI7gaFamJfrP2qY7/jL+Q/MXaBYcf/415T/vMAuCrT8vd9G7C3LZGtLn
oXRo/zNByOyh2WY15thTLmW76Kw7h9RoOytvjizpbhLt3UNiwl6Vwt40swWt4dkO
cOrW9iQ0EFp97ZuqmxcgRHBScL3rnHBbxsln+9shA4krOdnToMwp0VustKH2RuW8
YPMlkcuMdYJllaqjqijDZA1aALJcH/7gbezzNfSHbgGC/fS4ZRTgLLQPnIZAHIxq
gkMIcXU0yEUUdB9uZhofoxVoK5xHwH+wphCRoT5MCygLC7NLrFNrqOJbpl4RbK0G
ROaRiT3KruUX6qXfcynRNaJvSkzi0CKaxGShUu0ybFM6GnxCLGFXYS0oxfmk67Nr
svMOQmY+k5x6UGCdRSMjoUKyjOdhzWNnfBBEGgMhMn2iGFMMwG/0529WLRA/f5sX
vKK8FGWfrpodV2ZGAwoIEOSWQdSzbcJ4ji51d8PgsMhPFdpSRpWlijHigWGwftDi
MzExMMGM8pPg/KWVn2o6Tnbv1xHhrIZf/g+Fjz7hY9IbIF1bFO/MFD0ulA2vqXDA
UKOyf5HAPpxW5V4uXfuLVv81Ymeo1AfaKCcxlNecWnPv2awjTKNZ2x/CI3X0z2z2
/3IExlSfek8ph4Q7DOpB8hhEyiyAsB1aWMSa8q8C4MW6EF4PuVs0bamLZJMSgoO2
tDCVVDqBuYjzRctIKjVVVQTXJ2iTa9LteX31KcOxgMThms6h6nNJHZ5rOcE0ePZ1
gF5K67myEoR/Qg9EiaCGJjTwG/0mYBrsK3n3iFO4pRs7C8BjUS0OWNQTpU4UwCto
jewl4i9Xc2F8JPpVWsx10e5LLal7I8XvgewDx9Jnku5yKXVifUtaV+yLhSkDAgmO
UtE3B7PmH7UVIm01fCpZJF+xdEI3zEa11WAKDmkCPw0JyXgQWT1kavTTSGr8mLR6
IoEk1ShiSFgO5144ABTuDVOv6YMnq7U+3ovLqJLTuHUiyQ8pTjuoD8hKAPhtPOhe
KUnxiuP5+86mE4II2ATtvCHgHZxcOwaBXiM0IKM1zEbwcK9yi/NsU2HVVgQ5n25i
IvSfVrMKxWqfc8J9stbsnA1idBEd6ISMcIJLpy1EuXeJCZLuCKA7ld5rM9saYARi
sz/H4DtA125yq4FS7any/w1ENX39FiwXubZ3EeUvE4Fg8mtNd4kuHclisIu81X7B
4u/k0oiah0v9bW1AAygP/r+1tpvFr1qAWlAkNH7FxAlZ2ueBeorY3UWaTR84Vbtn
4eS067OEtaaxrznW8DLmq1ASzZCidYGUiXVuAeb7aU3VtR5Zg/ADzpTnvgn9Nriz
IMizhykYwQov30qnqYKK8k9Qf0RlblW/57xfcRb3dnw9t/EVPkGGOOae7DSN7qHA
dAQ064OGugckQddEuWpsSjRW/Jz0ovfUmu7RRJyIpuxTRN486ZU3yHfWZ6+OgWSc
E8C5NGTWilG6tU3B1rp1V+PjjjRzabw6ny+ftICYjvmAXxwdCCW8CT6nyKj94WXO
+N/Iqf81X87aoSKc1n97MlCIh0m9MmPf6LRZV7SEo5DPi8QwXnn7UKJPF8OrtqaB
TswxKkgY/zi9yHs1v0DQ+XiN3ZXenaasd7I83LVcS2Hbl9zlN7RiUTQ2JwX6YKWz
qgk4MvVJYicLjCf58PCcG0K6VcImUkR9r45WdUxUeV5ngETeeHTSAu65tuAwjgtN
lb2dy4xqnodpnR4bh8wxPe5Dlf8kIavpy5fRPDmrGL5j+5M+kavhEWBLnYL5noW2
EXIZIC7gvno7X5PxxjqegnWLw4PFIrIN3YCAAjAyFYwa86XhEGwjkPw9o9CzPsoA
8rapmweJGS+dvIcJ2q/2M5a6cHw898yInbXXa8MxaVF28XsdeeIOuo9x/Kj7AJG6
PoY0W8NscyRgMvhh3CHeFRfj/oghIxs1eXeUaRM4DPYPl5GbaNey6XyQ5EAxptn4
MMmgZOp8sGIsAMjQz/gkW//YZVNFIoKxSb3udwgT1asCUC9aVsnfXnwQiy4NU6Np
mR00FOUqAAInJZmQNTuYrc7AL7FSfjS4hW5mST3VEf3GmWUoNsnQQWNPeae7LhaJ
cHDZISMWORpmY0lwMvGo7/o81n3wQyfLpDaOfdsQrgFA3DQSg2SGLOfOeEclUCdL
FFsvg7WpBa3pWJr4Pj8JBQRMuxfeNd6X4q8H6X8eJmogwkJNY5L6ZGcnXt8o+dtP
qTvoBxSv5M/ZEVOhYgfEC9yJHC24wgO35iuWpxAz4wFNunGre6K81XTV/TNiO5i7
ajdIFiAtKvBbvy3AM2i/61hLly2le8+gINwGMnnm0iXAQRhlbszRYOyr4jzUGDE1
KNjHZRNhP9I/gbCmRn24PIem6PZuvtuUiTn7EdqRzicaVfxbx2IyhbM29hdK8Bfe
tG/IRN7xPIsyuaOwJkXXxGBuu7Q3ekk1NBXMsEvCb/lcoLkP+yu7F0Xl9Z25Arn9
NhzwK/xQXp67xsdaLY7aIpRDMogVN+xFILxNRQWh4+GoazL1B/++RK2zqjQQQ7Nv
6KGT8SXT2nIiSOBs++m5XcW9j+JARKDBZ8nilPBIzXRg4U222pfHJDNkr0Pgrbe6
AC+YIofGOjMUb1hJqES3u2hsw5MPE2/X79ozD9chzkdcx0hKqDKRqUiF54w0l4c3
dujpaHaCpSgrfKCN6Oa/GZbAZHo1zC+mujfahya8LeHR/B3+0jb+gI8IFQOxoM35
HczOFNqWwBRwlbyz3kXSEQda1I61k4fODRJASQ7763bLtC1w/bIWfF73ZAKMyryj
GORQqtxG+plXOPlQEk8cPZ7m0lPbWFt3svabnfRPoMvCE6qg1ocmF0NOjKxNnDC9
Pa750VQIGOm9avbx2fjDZ2tvI3cWQUzbm2GIRNJcJn1YnkbRl1Qgka+OTNxmcauB
Ap78ds0BIU8S0kRnxN+11Iz6gCKZ4fHyDPDzmAkO6ZCpqEjjtRUZJWjwu0dmgPKe
FU0RLLKNVCA03eHxMEsSzseVFBIP8h7x9TR8IR+vgTf68lUTJprhAIu/PpIslqLi
eMEIYA1joLuf4b8UGIammvxFIVbNIDVsZQzgPsENyepGckwAmL/kfRHz1PdTeyl7
qoDjXawAZfHVqzHBPiltv3beOmDoVKkvjhjvnDB5lzLPO9Pqv1/Pvy4tzgcTnltE
HWVK4KeLGHcJdT6lK8kL6QcykeGpDc6bsPzjJILewL2ImByI9rMvnr4LSn80s1XG
B+nSyuUElIUZygiPr3Z92+1ohlg5bv/chEM1S/rqn3h1hx9ZQTWlxPrEOJA7Y1nd
2UyQGkbcfYbWFkFhgbO1mURbkaHv2XlJcKU7tSh5T5SlDGVC/XIPqXhDIn1vgrDQ
10kV601j8x5NAX6PRXZKDLcAaaDmSu6XwCfedC12aOh5yhxur2Xm7lCdrPxHmi/2
S5TqP3l3rHPptul63sY+LWOAXlTSGYTYO/DdtBJ9B7DvpIvdOLKDv+T7tnnodlf2
wkIeeqM6jCZ14cjoopjQqpJC2vTZmBNFlp+tzMgUckWF/UKrWz4aT00bcHBYI+RT
zMrcudDYYNGOCF2Ht+5mnlVbjfEXlsILUeBufZnssNGLakrEV/xQxZxHqIHMRZsU
AmhoIoOxl764qtiMi3fHbtaYBztJ5gJlQEPu7QQ7EeNAPSb/IMEFfyh0O6Js7wEG
A/paWr6gnvwkTST/VNYGvnyaFzAI7xsLIca43CozdjU5m9UWNAkh+aa2D4cyAqKo
DmV1dI2P1CUopBTpzBSbL1MkOPw90XYufzs3tTv6UHI6XxTi4Fw5l97akzpm2+bC
6dKNyyll0RB8rtpY1lD7bX7gokxo8qWMhsDI+AAZZv0L2vr9Nj6LsTopmnM8gaHz
QDfJsX0zPMEZ8cRsPIuyri7WKqhX8KccwVFBH7CVsRT0DE+b9HBHRy8vAcAF89c3
h96zg7Ws+AXss1TM17ebvZB/5CD3JK4hpSnuzps3Ld6iAA882vIoM9uR9auVGn6z
VUWBRlg7slMZ6rQLTtRpSW14FfeAsreZSkL6esRM6I10vszD3Wjiq8ieYm8VGeYT
5Oxx+JTnoVC9g0Ks4twn36tIzcot+fe+7C3VHplnwqmZD4KjjNfv7hf0iRT1k4o2
6rn/dJpyfmd3vy74BdiO56wnzlpSBd7CC2aUWkboVVZGiuSPbOdh5J5zklmNvoie
UolWC93o3YUXC27J6NZ4qNg3dVhfBMwIgGmv8siNhLUV+AGdwohC5WDiWuTSFNvI
NIQVWc89EngyETmOpbtNOr1J5XZ0VKS4jEjD0A++Dh07DiVbnrcJl4LixGE3/UWP
c4/suNVFuItGHLtinteBk9xTFsWsUOzBFtLyn+IKVA7Sk78eEYlX1rPCBONAvKzp
JK4hK78wNrZq0Zm7ElslcPAoMzvjIFUx7Ud78HHXeNqLsWpzhKKC7IA1Duxt+o9o
+LwsvvipD1RkcyMQqUHqebRXpPfjZj77TEoERUPiR6nv13Eh8Mycqj/yIizgW5BA
35+ImA2Whvh9Rc1hAtjFudR/uVYRgJx4kAc5D6Z08UjIApdSymmmMvixez2EBdM1
se7awKIi0rJ6BQ/XQ1IxUWCM1C5J4YSAH+05Djmv93IlT7tGmxB3lLZY6U7k3IIM
HsoAssEgRSZA69kV5lfVbmsxJxSkfCkhIFXr8PElS1OGjzmXYXGvjIpio7ByLU8Y
xlqklVc82YRwpbZK9CTRo0SjgiY3iliMVHYb173sAalN9AG8TAKVMzwt9C8PcjuO
3gN1aMGpUYhvxqAcOjyCrxA4fztXkpVCPpLqbIYQaWL8Q5Gl8BAO5GoOjdY0eItA
MOYJWjRgbueJTxcNI37Y9djlD5C/aE7KL9bHWDmVvJoxScc6krYIUohszQG3hI1T
6pJDVKDPezQtql2yKFRwDRD7ArFAWEjELlbFl7KoS+s8lygxY2ta7QxgKRHIoGuW
57YvsFQkYed5IbrI1h3uPKWwebuBNttbxdXoTyxqdgd18iYhBGdBpRvVnQ8NTiCo
RSZFHxmdQWcLpuruXZpCuesIPfmnaZ7xJxl3uXeT54DH9zbcPFDXPdqW2KYiN/1V
aOhhZWRMPXhem/o4nW0wRRTNlqLkBSEo/sLR89SG+1n5fZt9X7bIuAwVo1vDd1oN
n278iRfI+rMbSPkWR1qIX8FqhHMRhtAeoRgYfBJenJQ5nIW25VM6rkXVoZGlGnKf
QREA389LB0RHxIJv0uUci9c+Z8n3489qBgPr5oLhs5x6saX4Lm1vaYWeq964tW6C
A4EHRaVnQBfnIU3UjldbetGWf/1Q5kzZREL/ESJBt71bPQilyFPryd6U049Mcgt7
jTKHv5gSlwuAjoS5nKoYa0C7deAxWL0Ydm6sXP4ZUNMk8I+2Y1xYrp3ns4oir7ds
5ufWb9++RkrdHSTc5/gaD7whSAdDlGjARs7hnfJyPOEDMfgKSBv6cWGZfsUHzEkF
ghnWTOc2EW4abKZ3v5EAv6NjeB+AIbouLo7kt7SWGlY2Dljd9t3LDvBBkYovTkWH
hjgwt7HNIpGIUybPOU9LCO4POZDuMDeIbsRfVyWDbULIgiznFTyL7Jeyv6jbmmmo
nqadq/BPikczj79VYPzSzgo+QXME8xC5mT0OSHV6iUfmZAX6NtZXhXsS6eGP+1+M
a7NDwhJ6u9IjaeCwf/gjhs/joNZYrwrf/6bSeVIRf2OMGUM6dphJcY7rxxzf8spA
RFA6k3MmHqLhi1UWDDtlpF3NJLEIFhJvwDIiJFMxo2RUjjp3LHy9f7VxZ5BSKvo/
cXIRBYmdMpueopcWbGcQUxUzVzFt0yeIuGAjIM7Fgco3OCTEu9moB5GTVDuxyNzh
64fLxVfjiiTZ6hbGVqFvRO9VZLEwk7mE6zPHGiGFGgE3hV1YV3FY1JV8JHeioMUE
AT7coyhN18VZVy0siNJlhzv+p2bPVIIizOuAOI1yezaz5hBG+BR3lGjT08Q9XTZ5
c1Sp+nsepjJMGGQG0vsvhdaE7y3Qvf+MdJ9qS9rkKHzBW5OBxsotcZif5dKvuP7D
RLPox2LNhKJoIGsoj4Eetm5Twdb8yqHkBFkirw1Ze6YYlVBDJyz2IO06anxoVS7R
jYMx4YLPYIGHpNFhgvIcT2UOq8wI+/CQXRaUpoOmScfAiRFl07VCDrch08Tsu2eI
qhG37s1mh5ILTjm/AM1MAmEiqViwiAuaWPITNepNa/w+vSd3btpgoW7XOWOSVLa/
U+5ZA0lFmVg8vPyNA00sZFSwXfffqhbGW1IdmocDiva3UA8+dldfinvKEDTqgEAJ
ypYxWHKnrIqVT92o9eXqGpXu+nQ7JkYBuOc8xoNXLLyOpR7I3Cf0HtlQ1vaq7CDj
W/G60EL6iLD45S6vF0PCnyVPAU5V/7xzjS8T+rojufhIRbCTn1goGEZjwWt6JAbO
fGFqqh7YUdztdRdPo4V0frP5x2uoKwAPA4+3lywlm2CTk+MZj3FEmy1vfP2OzKbl
qcNBvuiGXiEDONs27zTXPQHiGSeaGpRJCyCXpmIgOqx2jBJRohBVFB/M/QW4hK/N
gWHgDKxcho2lYVeywzC5pgF/mOJfGentNVbcx8MLbdi70IiyZUEvyGTyEpAYqq/J
ylKBPpdY1qSRlb18m+WZSVm7ZyHVe1DHl38o16uQqa0Z80XkSNjw5zqubc7he6Aj
o+dKAEJaPmIdM4UrKpIAvPAvPO9jYRVNDUrQ0340Gz9fgyIi0Oc4dEo+nmgW5ls4
QuFzTyxq+PJlK855Wt+WOe+0Xf07qqVZ3U7KqF6U4H6B8kDVuWxdJHRs1rzS6RyH
bupLXFraygVRKELtOb0okuTcC9y/Be9vLAEwVSzGmHY2xtSN3hCzUoamVISvfvW6
ga6eibY4mF9TOJkbQwfjTp2agicWjXvgXpOSoQbRhpBq4JPH7l8UpeSXcBzsNj+0
lnFHJXk8dSKi1ih9Hpw40sM582YMVjvLAvswzXcohsYhUecqjhhRQzrS3aJQAcyp
OizFEiqtSIi8wkflTqAK8peugeRph25E2cQTte70Lk5qAGpczKfho5pIytDNC83K
p5xW0FrEfsJE+r+1Tp5G44GKyTCSWkuQHOEbiBYJru6T5XmDgKTxzDsNdDqdUPDK
fbiMOyQGlliRLfLSUiA6HTKowP+FAN+3ava/O5IWkgZExzs/jHahqe53O9/DOYfi
DpCyS2g6BeOI3K/Z7qUdmjWYdSPehbvsZkFGjhF8l7ol5RpX9a3Gg2xB0UGiEKNW
ZbB4Lq5Pu/tIEed59p/76cWruXaeK2YXqRrn5wCjFD4aKCK+PcIeODQK4mTPnog9
tcVqH0tFLPcXBK0jWu+GW376VYT6LJJbf0LdAQpwW6U9NM6u+SYdVfn707aU2iUn
8/JexYSsrkiy8zko8uETaplu2ruhnuzpNH7FvOjnpcGDHgvADQJcPz9cbdCs0q0T
H0TOZROsc7b5EFYVcMWtNjGvlS2vHYRSmt++6IV3NJ20XwSyFqGE954M0r5oNxhb
L6uggdalGrI2uR5RlYPcxa18Wlzh4uFj4APZwsswaEiF14EQq0yJB6gTfD+4iLjh
EWLIJoPRjWXqlrqKvd9Q+33sIlHCzyQmFHWTkfGfSsUlPcD8RJpr6/m0kN80s9SP
qou/cfo+722Cpd2S2nF/7LueAmhJBc4rC8LvhLeaiAi3mqL+ygHlry7hGcAXOnrj
l7LdF0LbeN4lE5sJ1ouY2C0qYyOhiBmpfgbGM3nD3P3NMdMViZ/I2zaC8Vcu6w3K
0w/QngthpYg1KQGTuw83EUTnV5bRES9bhj+hQ3PUoEL7VVjpoyFXCb0tvxD8SlH7
WMcAUVAVtes5tJf+XAvrhhyJRr95J9BBoUtdhfFwJgJFzNx28FVIxtdIlfnlhIOD
jdxuiDJpZdKuDeUuaqc5+Qg3GxYDYLOWEuwyA1X4iesr+FFzvjSqWw7D5jra7vWk
ch4Vhtly2g5ROP3B39xL9I7ufyT5Py7M7L1SQsoCYbEGUdTCxaqpejOKzewKE8bV
TnFrWesFy7dLV5D/kC9b1HMFTVAAND32s6AkJCVsd2ntcGSoJ4lCetd+ra3azm6M
ikme/r0jatpTH2W+l2ySGeHRjIzEcr778sAxZIlZR/xb2tTO52PBnJv5sKineO13
KyOKGw161gFGTmlobubxkv2Y1S5P/Pct7yi27UiKmW1X9XmpH060lFRVGO5bE3vR
+eVcqaXhz+pCMdV/gbjpcLhDzNpGsFyRTz7Ai7qfjlB2jCmOPqTUkO6q0/EexiVw
TI0SMF990pTTEGZwPQhWPc0fW2NJU4yqPFc5wkYmbPX49ovRABLtV56b5DS7cEWN
zZQ5ZjeYRQ5l3/al5OGKXF9vALynIzklvPrr/05ttQuFOvIw9l9Rc6rWf9osiLKa
25pqoBB+hjM2jcSqVqMu+bzzPJgQ8DaOXdTaN+5bGupPFTeEadUm1+odzEZ1rNU0
c1WFQXibHVi/sz4tmJQqxIBkze1yAKesrT2qgyuzR0zUi8DHeEPA24kKD/qjKcv+
D+3r8/c7mpSJ5t4zJsBhlSvMoH/Hr0gLkN6ad9/GTZ2qsPD6Wi7hZZBvZbLq0IU4
I9m+HDuxVKQWyMjx+/QrPB4CikPL1zCeIiXRXkaQI0J6KmHMjiMm6i3aYk9HZH+q
ZYO092x0ujPa2lgAYmU47K7xcdcFvMCWM4/eL97GKEJ8yOQYP3dRVtXa+nIENWn1
M4JgFbi41FqmqPdRQ5OxGdXX+mVsc3YsYDR7R/OIjUsxzPFTpaRT0qzykROgmytj
IFnZ/S0IkCnK1oJ28EGySCgb11s1WGj1dAZ5a4xVHDKuRcwjn0qUM0NE5YmkbDFF
MGHALwSnxI5aTp+7RnMZO5nOa6H30Ta68MbDYwv/FXeJRkZBz3KE8V2acycvIDjR
wZp56/KDK/qhyNVt/FhUv/XsxBPBgrQFz5ZeiGzECzozEoVcRfqcbLyUiTX9EkkI
cYRpBq8X+Bm+tsudO05F+Rm6p8oND0M41iL/++QxEer4EyKOFa8DmtKn4c/gQgTi
GXvGA3n2PCaJTMXNFjsDXnGGOZYGv8DvJIpGtGTmw2ApWMp8TQ11QaJ0BmeSCnvl
9/rWMqCfhnN7GaN5KuHX37algZdmrNSxVV+nWFoROsX41MfPbV5ccNCTlhWw1D5Y
DvjiR+v7SE4eCK5/3nW5q59O9fSxDU/sgIDz5d9xUDKoPMq6J1sp4h/dZprQcyXR
k1IhEAQ591mZz9Tc4zG0fCe999C55Dsps3wnmWf1jO2v2KIJwTtD2V1sLZE0HFL3
12m2Gs79iFQ0TOawie9H9xymVABl2WlyK2/n27LrRKtTXGT2HbKGj5s20v1zr3XJ
ft7Ztr0nwh28XjaVgQOk9z0EUfFsCsQQud5812dimPZQhFHIGn3XCE5PSaI8CH9z
WQS1gowZjBLjAfYRDLreBfmuGOwf/7OT7V/WkPcF7WCVXFhli8XN7VK/3JvXCbWW
z1YocqV5wSK1VcDKJ90iAx02UebWRH2keFdmccf+IYCr+jJEqTq44zxste+REN8S
oHv1zEj0ZSg2O+e3u/OU75BK3gkJBeEWeUkBQpTmgGhKuONLdXF8NT1mL3Z6hd2h
AGhhIy31K1hUfMecSK1+R5QqfI7QneapEEnZmPxyKrFEtqWgj04j9WUxPM8w8wXJ
GZvanWhaJ+SWgEK4HPMNFhcOkXAvIobNT5ZEC/vUxSkMYikc/zuMKzTMynOvV2pT
V+aeBGwgi4QwpJMi2puwviMnNtnfKMOHpeoYeWKVS/KPQ1E2KXdaAtaC7JONx/XY
pWnBb8qlj0jzCliZRGyuvgQePPsNV+OrGMtXLFylPkck2ERERNVZMsq0bcadXhjA
BG02hQomnOpghbytdWRPfqZK3nPMHKzXzzdZZdExuB0kd2DVGPfevLv7FJnNGF/q
qnSt0PqVyW+vD7xGe3vnbo5UWTkDCpdsf0sJO3+/AvA/wthaB1+vzIgGMS5yMEEF
XxM2yINo95PBs+slb4gNrbbYBEE4nvF0w1v8emP7ksV4pENgPglryXs4wCgHQiY5
vynv2nka4Ncbd+pT5FUx1Y9wUIOIPHBoUVJ6TCCoMSBDZcL1OsAciT95Qq7GG/6p
2PTc+zektoFGHkR6vM+Yml0hiAXI9olWMp/fpBcTp73L+//n6TbsGy09jlPRgrZP
9FaDpR15cfJX5EKddEOp8l2Vp2v1IyDKX5Er/F8K/c1A3pZk13gtEjbqw1dnt1YM
f+uuZUN46S3wtWLUqMSnyQIkmm+8LTTPsgSeRlacIOVSg6xzA5pwJ3fmtt28x0F2
crXbVfhRqqIj8nLSKyOBar4hFZFD6qwq65zWVGMDUA6RZHofkYNsc7W7WLK3gdmA
gJl/Pxipke3cCs4s7w35lWyaVnOd2Ba8FOhzkjHiGwzajD9dAmtiwv9cqVK2os7n
bu7NrWEZqENibirDV3x6Yo2kPszEgFVtXMZOfJ9ap/sTQsd2zCTC3gGwb1GVgeG+
cBBm4nz/LbDgZAAw4mCi9jOdLYD2fIfxEnqYtomZWxxrK5PzEYDotREJyfggDF1P
M+4iqZKMGfIPB+sSmUY3cHi6t/WN3Xm+0n5DuIqcm9/soT8oIZtVEjr1qH7/wW0N
xEWgnNH+NAN1iP2k05ctidp/xVifkTLE/aQjhxaq54zdlsHCnB1mdG26Dfhxtm2d
7RcSbsTrcDPeXqVWnVZaz1FHk+i93Grkoiwr5F9z7ORU/WyMWXgqG0v8pNfdq+Ep
2M6sdhUVaMatz9F7A0vl75+cEVxL0Di6lNmMo8y+/0ozyXRk1uwZJfiRd0ESktmY
MquHEjZAPwjTIf/4WSHIY8/hMElPs7qUQlTpx6gJllonxPoOY8liv5d54/W4YP29
PFnmIHFfA4yTm1PdVbk7Fpda+gLj8gQzhd1+/uWQKJq1JSAe/gptEhXvyiQul3Pg
Pksx2ebB1bMJ/WRaPO8ikgXK2PXaZIdmUrw9bSHMbi9zfLGlJEfqlQ5ZigmModSg
KcbXtgT4yKv4hh2Oy6NXhOe+5fsiuJYdpZ0ZrWI47bPNnHZ1kqRXr30Ae65t1wq0
ayJ2v9H6ZHBRUe85EHzKKZyRpeINBPj4cgd9mjCp0ZpW6A8OMzXIcMi8YUS2M8rw
bFnW5vCG+jW0mC4Ecq8KpeTZ2I8sATB/a4CGs/lXXemlePF4/ric6HfPYxrChIuB
DZa4wjkwIJAnjjhI53P5KZKCjXjy+MaZQt0JSeJPyywbc4snFrUApkHphy3Wkl69
nEbHLnYo2ClG3pwPjNuOXnnLkaCg6IfSYemIvKmMaMAES0gmzo34qoC8SZAQW9lc
JpRnquzDjiby2bvnsA1suib458v/Vb/0rjiZvF9z8ZvEnJF+z6jmASmQhrgf1Kzm
9WdZTc3AUt5+1sv54MiLnvwES4AKKBOpJawNV4Gl+KlTOcOGpJ7MV4+cy3qoQ2v8
DKa3P8sIFecW937QI3bcV+Fn9d7r4iGD6JJAuMZG4CTfHBL0Kv6XAv0bsI1lKD8u
+Yr/YInzIiJ2GTlxrhiY3dxpu2CLjL2rsQjhcOLWMTxRWTdAJSafjhmlwkqeaN84
szwkthTpogU6wBtL5pZaEzqZqigWF11viN8XNx9qhNhnnZ6BQTgzdRQctFq/ORj/
hG8q60GW82HRjsTUdjdKvtPUybg1jqQ7dX/7Y7ORem/Tl1gnHcjG5YezuZT25Ec1
St4rl08Eov0XH3iytKds1VAdcGSn7QUxpqJ1bocrcgcbM5RKok/x2gJVD3XgcjXd
vQo+BHijjTvrj5mx1f9oyUVXEw9I6g2V9YmFiblAlGwmK8HLuft0vk1ByvbVtvJx
dNm990aIUtkhwpvjmuAqZDenK3c4JU5H+AVcvo9wD4BlynAaA8giwnYkqqa/2n08
OlVKdHpNVS/4FLpQTj7jCIJMhXsfuXZv/bWEfuo4DBePZM9CMOZIOjdzc623j/wx
0VUHlCUdRNqnTSdzjvu7JQczXlDvkuZPt7SAndTYV5aVZx+Lqref0noAfzAMvYNB
J72bYnte5R+3JF+wssq4kZqCbOL/WEcWRxEfdHwh4/DoU0XY1Joh5jwOB1PnSNTg
1C6P202CewCUoWKSeVA3FTXS6nffirDnxCstEhOjJ15I8Rv6WsKCJnJ49wdgb9zk
0Ngr0wjiDXvu6ELlzWWunSmP1h3nsNrs0PK5SI1tPhGIWIlNqXaNzHSijy13jP3U
Br+iuxC31oNwEb6MnaoQEVAzR+V8RO3HqfxMt1BFuhMLg328txHQrTzJDRcxGzzy
wlKP5IiA+/JB9pXgi9BjoHfM9QgObME38UxJftbatELXIwbwoTY8d/5ikiV5Grq6
ttIfd1QFvQNBPrUb1WhYgtnU0x5SE/DMhXCqqg8tn57BFWnVddCq4KW9kxIZYkyt
rf8nuWOLo9NipmMDcbolGcpr6NgV2Pc9TIu/xBRqtbVNJJR0euYgXv1JibuRsb6x
UYEZhDGprVLjF84fvhCKrAwoKNT6jmS5Z+MriNYZt33aip5BbKxdyPJIRYWLGURd
ihZz4Xx+u4zGeXvNkZw58yqA5rY4SCvS/MvFbR1MV9DzrCm/xUc279970nZiEMNF
U0c46lmAAijWMWWo3+pyrHZd+4oFTW7RuESvVn6+aSbSRnAiREJF25fR6BiInuUL
sKefXAdR6ou6vgA80NtvGqNuEx6N579RlkSXxCu43+nF5oigBwbbCZVBkDQW7tKR
E8JgCTC81I8hJ20LqysvHcjLYoaMse9Td5x5p7u0Y0L3gHSm3VcW6ZXsdGCDBJAw
Bl9KT2P8HaEt5QfF81CpdtCMMNI6DHhnmPmPUrDZ/DJoonFg4O/nZpR8+jMNGTlw
nsqFMpuG+kKjLucaZh2ZqQZRDAlB17u2svGFgdbnnz8/vh+cHSQfEnzjY5tge6RT
P0bZY5JY3EjFc6Xs4CUU5vjm4t99lNZWsPdQvRxuagq2hv3dXOQRQ8/HouItywm0
EE4GIFwhkiiVcB455EIEMEd8t7EIoH79RiuUTX+obMPYuCZwFsVWRK+xiKe23uBY
0nMF5xqXwnKLeoTSY2/IEP//U9AXyhQZ6JGDCYVs7Z4mrDZ4iJb4kY4GfP4Q0v3U
rH1R6teI243j0+bTZuG7+n73WxaA3LJOHNx1Ww1TaPUjlDoID7kZ+Glcks00Ehrn
Ibsy8G46ig5uFQCPujgX52ZlkpB/Nir20Px1lDcWPl6ivvjYt4ljLxmxA6ixRjm8
nZEG2U8bH+8rL5BNjQv3/nWCRHPAvlNEL+wg7p7SXfCUdSBhZPIfXA5M6EN72FfS
rgTyqqeoCvnDPNA6Wx4+gwUeXO78nTKcqjuEVtqMmev5Tk51K/6rlvc8yYNwdPyG
J8fHqVktCf8kJ3ZMsdYLAf1UsNJXYYoaM1t4LQ/j4eQebkT8IpmnJPn87+AOt4/S
7N0FqooR1eE9I9WCyaTr8yeiIVB6dxp+d+QDhGYLuk0J6NHe1Y76INoa+DX4+Tef
3KbnigpPMpGhJWuamM0xZHwYdx1i5zwtaTNBZ1aYaI6l3iuY5u4j8XPJRlVrZDJF
HQ3WLF9J2DbwIwplvU9P2N3eZldNdVUMPx+3Z+u9owHSQf27KDMUhB8BsGt9LzIc
m0QgMhwZWnXXdBQPolcxf9FRKi8mWzgNryjL4dvtPTY3Y49EYdk6zUqEsSgi7iCr
LjAQfml/e1QQCgBJ7KNlvI1oyl6lAvo0wcy5RGIzxW843i6qaAU1ovSfK87L9bq5
2ssyQmkAeKJ3eXW0PdkyJuVlC96ZQaKeHlsdOkfrH48IbOw8hHNqorCuvLnBqXwe
LwqEwW1zI0FJ8VhUO0h/B3SzG2t8EnEsWhe8lSq6KESzyrW2uFqUJ0kFdFADYPnH
jfMJ3fcBoRQVO8FBtaC4vhHyYF8f8n3AOAGxnA0udL6tcJ7fXg3Vx+0pU08v7kvt
rKNL9owJU99UTUgMGwSdSm9eDfdkq2QBIwKQGMbwsQZlOy1fDxyaROfB2NbwCMke
r7kfMTQc/t7a2dnNUEkoUCdp20KBsK+xM0GPvLdjjNxPDd20/UkhelgwL+DzkyYR
Fsqx9GJQxmfTJf6j2S4BHH8/98Dv6AyAwb9nGjO8HkzqCuBtJqY/Y/oek7yXaWlK
pQBqQoGXfY8umRkpZWHOiZTJFmUahefaFOVXUCKjx5r1AUhkhXCaI4+r1/GpoXMn
Cvm8iRH7HtvDpqLOsJ3hRNaQR8uo75sUb3bHMf0OLJbcS6LF5CI3L/qmepLOMm5/
x/fYMcLSvKtLCZj0FOryVd/qQoeqBCKInViajFebt9VLcYANsd3SW8Nq8BIXhzyI
uiOFxCq9neizSu7CxgOzfwKaDtBpUy8HaH0VxynQvhIrfptK82Qjq8i0Rkijo+ZW
odzOO2K1CIoG3+tsdTEmG110FAMjAQc3XBxef2KoqtnAv6Ph58Pehx9BF/55tu4/
meK6FPy2T8mEIdWvqpRsWR60pg2BmO7O0lAfiqVZJIx2LIMbDDlM7qGO1g/3JFGs
aH7PBHm8NmG5u7AuLvCp1MJZBYtE2K4E331wZBnbfnBRsHlFBdN2Uf66j+QutVxr
u3zB/cOehdKQVrIKiBSjR+5bHOD3ZEhIaX5Ye7NjXZUO7n6MRCOlo7+icPXhazlk
5c7itOreR62rd8RVmhOB4B9CtIj/q0yt1zCMxC+YfzU+DfI098v1z4oWsbiitvkW
vBCBMbOubkkAxqTj80T6WbHxbTS/h0IZviQq9UL6emwdkQcuzPS3w0cBGFq2oOBu
XNrft9hyqbv+HhWYS8fcTRcKJIewL/l1nWg2/75gIL9KgVApen6xUfgUyvbXGMwr
AnLVpSb6XxaQwBXOzSPrxarr37Bdn6In0TtP7NujbpaxJbzU41l5/g/2jIIKa28G
4mf2Se10hdEM0jp+h9fKT/Bh6jpkyef4iwFO392xGoSgY0b5eTXWx8PPEob3sM1E
LPUpHUi/BI0OExes9ZR9okHyzqCpOXVly5WIsUJmXhCazI8Mg/M6xtF4mZ208pGT
jtaJZYrPXGXNL8IxJbODPugJnJMamwI/fDB7Z9VBSFzgIfH6YW1z7O68jWz3Ph5v
fwbDVJuXrsYPtx6bqbyERGzLTZMdVsB9fyMLk7Io6jhtzO4EqlVzX7VBDVC9AO45
LP1bSf1jYAbzmk5ldtZF+uTn2+x/4Oe9Ok1ymVAL347WyzDjoRPWkbo5Nv4mpqWg
vzIqmeZva/GMB6OiJ0fCU34B1VTHKmwSB/Ha8cfKZsUiD1uL9ocuHJOfuEcGrCkP
A7L4IT8NT/E4mELbzYJo3mg3Y0IilNmcPP8NeuzaX3StLMySnNNwXM17m6/HXBhD
5Ic8Dh9+tjHo7NzvVjCk2zww7XgC7DW7Ifn+GKTD+lS7y94EyXDdlfqr/vT6Wycx
0XmGKYjSNtd/H4inihURZPxpc8Ezz/vZEcOb4FaX5aJnJ0pthS7g9JnVlrpIagNg
8xZfOcQVPWHKihEfQsYMW28EAQWnwA08PZjG4YU1KAK2Ov8wsqiKe5tK1eJPTak7
hHQYkkr27/aextb+qCUW964N5EfMDrc2GUDcxkwWLwP4pp+Qp+alv0VGUFSCGq4I
I64KgLdUP9YWVDM6U4MCEDs0n2BF9CCrO77nIwOLEGDh0dsjslheAzIFri7mC5fS
7OsqYwxa7ewqGvdQXNhtwhoBfe3aCmKe5qTxl3WpzYVKtLM1yVw4MlyP0qw2xvjG
ijgLc3K8er2XuupXd7UsJB02NNbNIDX4HzaEdIKEllny8fSZDlhD5xPGDsJrkSbo
BX1/qio0ML2WaWeevKnw7OMDNuZvyXWbBffNriiNd8Ugv/M+dzmb3Q1E4EBlKsZ7
q4oiIX0ogJYjU7wY5XHID8O4fNxHyCxhb725Mo+J6JyacytgtMRIeebBsXEGQU91
HUN+pE0eVajsRrz3p0Y6nx2AbCbRF7dMsNHwr46SXp7Pjf+ADOltMqizZX7wjSBT
EaLijpA4P7ann32YSNsaTmWpyBsaZOMorHoeuLnI0RTpgHv1iztiNakP9BEU0YFN
a4z6oSls0uEIaJLFisYmMLbS76Z5sICGLUdcgEwo2yB882vWDPrI8Rweifvvaq7o
I9uSVyCzIqoRlelad1IIqUQnu1bkMz0nttUsrR28qobhHkg4KA57c/sfQI8QsyGU
523fVkmjStbk/PAv6x9haOKaOFa1F2BbhXvVtz1iUTCA0cWmlBRBLQmtlfk2gZMX
65HDby/fogJss+ZPSZMjmD3cM5ZmPJpZNsxOAE3uQQTuB+TLL/3UfJ8HCyNw2oXx
R33PLqxkw6loNS2594C+xGjXIv7lIFMdQRVSeKj1vAvtZ9ONvsehVldZAURG0/++
KWrQMx71CKH3v8JV88zI7Nw1xpXMVn9LVUBApcJY/Ssq4oMoXnHzfDdDU8wgBfll
G0IqctJXsuNK5s59WnEAqAgxnxd+5bh6qD3wNI/CyscgpfBCR/KgOKhBqmtBSnFm
0rWbuKs6nCWmQYWfNSGofuiM3y7bLouoaqTT/aPxy5to6Bfq9S5ljSCER0m7XTWk
9HwT/LT3gb9pSlzCNuA/c68cposrG8y9vu925UBAtCr0j2Dd9pXDOPGbkcboEhXw
NjsDQC1xLIqTtlVifYypAtIqiXDNcQ3TayKLnfEnMvdOEhSqmmTu841hHfQR8nD+
F1B89Dm/IywL2LwN/4LeIHKlNhr3M1ahGNB+oLol+Emp5JadjxAGZPHCJs4ijIGR
rQfg1l8K4Mh/CsWHoqcb3721wiEMBW89al6ioXJ2LPuDdja7yjtzA6NF6jyTGJ7X
O2dJ7QMnn5dRV1PDzXruXin93g3vkn/XLPOxtmBZMHPGnGtHMHI+wFyycjauPAMJ
XmyAqSCEvb4d1VVfcfwvoMWYbYhHkXXetMVu2p+TI4qBiloX8Oc9Oakwl08YvWW9
kGVZaLFcx06P2Sk4aIXNId1rGVpNYTcKvRfHPX/uv8znvWwtT2YovxovSkg4kPh7
OlV8tKC1Ec6WBcja/SXWYD57GMTQhvFV19s9wcBzWSwKdjHUWfsoDMXrdalUkVtF
QoUclfK36/mgBmcA1SjchzgeDFBSn24hNzcxR6QSMfUl3yumXYoWida0vNPnF9WJ
QiHs7gb1wcAEzLtH9jHHY1RBVuoShrtd8bBwGMf1szBnbcAiaHha33/OjJU7bbN4
xHenKuRu+MV+EMzPmc+30tvmxZ/2p2Eoh1KndL1atVzG5if6CnKeC2KeSpQv92dQ
6/j3CzeB1JFRqLph3wVqyQWl2U+1IZ5b64fLCkaCzU4wD/eZyj6NLLzk5/iK5+DP
kSLyhDC/XtCMyLibV3yRqS8BtYgmzmNvjNPvtZyWwIcpPFMHkfSFyZ4Fl1Xt/klC
AeheE3MsDTOmWRAabSvVRdQ2K+RGqw6++6Mj4BptUqpmSWuEkSIxyJW6ZiiT9aWK
UeWYn7UYYCOTpztFV2YJbXl051qh3JI/E4OqczdbTGJvSE/hfhQCF7+Awo4BFJyF
tiUR+b6YrmxO6r6pdutLbCD3YnZQWQ9atmqd36aQCad9SSMjfMUKFmHBatbBXbeZ
nH58RLAoHRqzqam9WuxwQTvNvp/umPsqFAvcwTQejzgXwBzA7HvBnftbCb4nMIJq
hOflOyWACrBI/j/oCjAGejUMvxsJr9PP+TrCVCeOaboAWEUsy9g1dd9xwHDHtHvT
/WJAWsSXDq4+ybC9GA2nafDRTp1oM2zmlEbp9XoLd1eGkpItJNUqeJhFBosT+9Mk
XF7CC5L7vLIofmpkXN+F0rDsqH/9cR9YT+/yEdX2+geCXf6YPE3WX5JYIuFtvt6u
BLZ01S9gw1zlCJB1258S0cqm57ENqJAC+rICx6AplS07CRw0jlD6L6Gfb0dUuwqq
AXEt20uV34cwcQRD6ti47ZDBAaz6QpF/ATTAklV0Xqx9jiG2Rhh2qdKXhtGOifi/
dpQco4lSSZbBkuImEo5noQwSnurSSTzjNANPG5RSelC75B75uK+w3SeZV3forkAl
IJkckRizO3uGANtcpbcXCXEjLXv96eQcZBWR4iPsnUtHWXT2e/KcOL13pg5JxF3D
96EKTKGa/Tgi7ecYi+OmcmTxFwen6Ucft2roL+ou2Pj/iHDv/+KjwVIIjXIRX+lM
fzdnbbjggKyyGOHn4sTW1J8FrSSTPrHCvhht+NmNFbzH196gVjMZ7yB9KVIWjSb9
0UDNB1JTknQuwMhDqG5e5Beucpto+6uM0F5cNuhj0tCaIjz29YfOTExZzE8A9TcE
B0/HDWU57U/bA9ovXfLz0QQT+xAyxqDKFVwelOpi8hX+9YE818igJsPWavhcWLt6
vRI196uw2jo/F6Sdb0qoYyImeAu0OuLbN+ud/TseieAKy/GK+dy8R+AJIZOexhsd
Nd9kapfctl13OtA2ngDLxGNbtMdCdIw4ioofRMMN/+Bc/cpmhQpPwElBe4FKhzph
7ZtBVsHoEPklmknNF8vTOdgIfN0T9vGPxm48Lfs1y2KVfH0OtYlw+JUjtK4zwJTq
6y45QuMAIjQJf8BK0IwiWkuSWMA+LwCPUeEMkF7FFPN0hcUBgCHMZ1HckEFfCmZM
OOCGzfqx9S6v+xx8ps6HhGyvKhoqfa3sgcwL7NTvTJQRJtIqL5m5oSqyuV10YPb1
rI4RlGhsMa7yAryh9WhivTJ35shKLOQWUiI7Riy0Hn2CdaLz27LGYwGvAMJ5C0eT
hI0ioEAoOn6v/u7Jnm5+UbjQ3zzsUuO9mrjr346UWkcjVQnelkkzmcs9QNJL2E4w
aeUDjj5xhC+BvfYAdVGV05UeeHhZR45P9F+xPej1sRDDTZomws6cnhrJI+oieepx
kr1KGiTw0FFsID+lfTlGgV6DL6ADyJbJHJQCjN5MUA34+znhyoHzyq0IHYKIkpyu
wC6aQTDC83PKiwgT0u5DIOX7v0kGdrzTEPTBdcnIonjDPs2ODdoqxB4u7l1wjryt
cYUQXZBjSh2GWSmU+ut3FHgm12g+JyI/D13gTGXW0RLbHXPnwaYLD7wlR7OUvkAK
kk7h3NuF31SCv0z9tAMuXdwqPFq6nHHQr+39LIB1nNvd/VpFQ9SayMjTBwx4I/Wr
fHCQ2qYl7+ydIuPOoAoy8XY/OHUbH6tc80ijdDVzF71Axf5Pnoqe72kDt0J9I1jC
Q7JU6X7RtWCaXMkDbTavAz4+jW5Oj0fN6zyvJtmRcnxh4TS7ui6i4mYEempy1faz
Vttd2MI46JpAHxCu5UgW0/KEP6m4uNO0unyxlFpQOS5gNeVufg4uGadquW5Y2N5F
2+sqJ4erm5YUoVm21Wp9nbs1u6B7wA0qeGcjFxJdVW3QEE5bTlqlJtwnzVqkv1dp
oLRMF6xvv99qsKSGHs+/7heNpr+ZffNsbbB0jUlSU9gZfULx7p2VN6rAarpeSvFV
GcJj1o2CEIu0Yef//XFNacgiNlUhB/PgopDo/W93mWOB6A7C0fgJrHGvf2BvcdbF
YRMniWxT3ElHFrmhS5LGuex+XvwAtowO8lkRcYNj4W8OQsCNxiAt1XtjhP4Zu3uQ
RLhqR6KY6PmiJ7sRi83CmfpcSiGiPFn2FilymhRFuBEEhrlnCfKBFxAl0zcXmeyA
yj/TXPN39YVQ/ttJvyNJW4qHnSJP1UYQXU+NZACny/OFONhv9T3y3pGXnLEF2qIS
2O6wSnOi4DN0+MKY/rfmwBiRW3XXszCm+xwTvN4V7X/iQvm5T1IVtdyoO+winHN8
t/ijiCO3Wn6Sonc4r+3fqRMggEMz7w22bBQtHBkiPQ1dR8UvWnC+UNmnfoGfL2jO
XlVw6xoot6wM1vQV++zzqij2uuwiqMT7P8HLjL0FNnyu/5YDmrpi68O/AmoZVOGK
XD6O7BeBqI1lUcMpA/f0xvr5zM4fK8WI6BIXHGGmpxZVrOTX8FWWfWOgX5gELzx4
49a3EaIF8EG30lqmokqaWvn7jjyUugNoWZ32Do2JOzLQnIbqMImhxGeMJUbHIwyt
u7ZJWzOn8Fo5iJ6DoPMu/QDR1x7txQ1dZCtHImyHgLNAqJzIUhchGjcQFXImAxFG
/18XWu8ByjVohEC5MMoW0Q0FlJ50Di2biyd/rg0LLcYwDJhdkKjlxfHZA/+wOd9u
/t9RZtsrBi+4rJTHm6ylOXCD4COVtmqg1kzOomoJIL8XgcczpsGyDk1aSXLt9P0B
bV/SM2g3RBg1Nz9xDrwqpq69mZfcygInh6r6nBR/PfKYQ/jGMrf32Nk06jFYKhBn
Ir36WyhyiuOavjn8W01gpdF6fj77b4YM+YCsrv5VPTjEMjz3yKKDOlcSWOCk6a24
+T8VSVJ7lTULiGvTI66W6/CvwZnRs76KcjsAHW/dyWJc3nbni3mfqhtGTkPfwcXM
DIWdAJa3LtueIgn5mEUe5WyriRJanK9ZTmd1E75Izl/fQV4ZN8uDZMhgtWXYbMt5
9qIfBRMgKVHSH6AG3DqlLGbYIJkx5l70CI/piTRVenWHOU6FanNLQ68WiwFh5Kcz
fRBN1GPMCdecVr7xcWQ4dUlB3pxc6FKKywfLBQTmgmTvEP0MLPteuJM4VMkMeCeq
ik9WKjvg1t7vXV2tc6o/Ou0YtUWy5c0QwS4ICryJDU9Ea6jmH3Ugl+KxlmA3bgNv
SX6C89ZNOl88v0UkuUL7MG28LR97UnSSQxQSMbgHF8HPcirSh6g3/FvsVDRzG7Wo
qELNrFV2kSc94vDLXPZYI9wogFpW1Ns6kjbonX0eBuEWPucXwCo+BafRsI4vGFfg
JQywxdZ+9gHwFFgcmIJwb5I7//lKX63AWH20d2yWcm7uQqrDlT9bJayujk9t9pC7
7BGY4koSKvZLJx50ruCQUH7SweH528R0mBu614ulWcui2SLGw40Up5RHfZZDV+F1
LpnyItm0k5R9edGnjayPvabXejotV+167E9FQTC/YuIyAZJwZ/cFqF2Coqakmy6Q
k20DS9YLyoJq1FPFNjscMYJWoq0n3oYyQkecULFpmCxbacDZzbMF95LliEgnEhW+
f68YUql5vs1+3YwppBJLEB/NfODeZohPZf0k359tiBSdCdZYItSVBkWc69drbT+z
7ZotA95KGUbjiZy/OKG8XmtvvwoWB5Rh4qTkIeDKE9k7/DCukymAbyZSaEcpywwm
eyAfBTsvuRERANyRPDqrPnNUarfdLtS7lqQe7QO8wMyPMofpMjH3+LTyjp4ZciHo
Snp9KN6h41XIN94C+weKAvsOIUrJOn2RkIY8qrxryeqRLLAuMfgcAAU2WkNN4XCu
Q/h5f0LocYA38Ic9eyZJFPqjI741qg2JMEhXFhPw8h02mGjbolmAfWaIe1Ldh8zE
YLbPmuv4ScxUhtYB8BhEZPJEYnB6O8ZQ6njtSb4C4jcopnOOlBgmlUW8jtsAAmxf
BJRcNUe4sqvdBKHlA7z7Zvgf7O5lyEN0AhyB0KxufHJBYtQhqSziltHQmOrRBAsX
KDBuPAgS8DkYJDS1fGmz+BcOYigP/5joY0CETA8idis5NSLTNx4ChWIGMVczm/AF
POSFFhn6NVLPOmt9aiph9VwOCAgC44mHAT6WqN5hL7z8OJe0gTgC6Y1XEHQWmEZh
/fBBAqDoI0KO9Kug/Yao+WgzvxwkdOlnqaA5xq7Iv2cTyKtf6o7jWU2zI6w/NBGG
aASHkuX60n6ikM0XTaNozyXkw+fnvdIG20uFdC9YL1uF95o0AVCYM5Iwtmki76so
dSQ7O61vxQ3Uvp0JeL5zy6Ks1AB/FLXkMMYC8/bPsBKRSQfODN8fBw0fbJ4u+A+T
A6E7vY5qproQRHPMwVTbFohzeLkhqRq1axWybrWfjAZwkPZ61gGEk4AO8CYs2PzN
vhe1voQ1/bZwcA9KUlZljlGb5rN740sgtkTCXZVyTvwWJSzJ/W+k5jGJMamCDc0E
YeqxARAmv7SCLYGjiL5ad1LKzRQfi5+HhCIZCgzqmbGRLCgDN6wP764BrXVuCJph
oW0qTC20dV0LmbGE4DyTzjnyBYffXVXpxwfmA0t+Vrz2hVVcpfLH1oI3NZLbP5i4
puv8hIn3UeYHg+DrIBdBxlwPdGgcvn1YPRtHSC4yZsSTLhY1nZsBdWgKASzHT0ng
R4mRiKaTAsvXoXHedBrmc7qA1BodLSuhMe5vaItRk/2d+WWLfi2fSP/pZgTu64Ny
Lx4B+YD7RPrGIqfkWRdhhDtHPINHdjC+vH58iyLLSRP2iZ63JlUZjgJuEaE/vJlU
enGYl9zTVUPfYWKpNyQ2zR7/OYihi8B2sUc4ZsxYKbh4SBdybJizX48IDyh/dn2z
GSR3+XF+dzuK+8Q3XojTm9qRFeUoftryZI0ah0kmIFtAWltaZr4LxO+11JVLlvs5
fOWUOlbrk7V9JeFOKkA9jcKABX4xehpBdnnJXfVw+LOWgT5vkwx0apIB1pQ8OzWy
vnRo+RxBoWmtOGP3DbzOV/m9qco8S4QFhJtkGYLHLxd3eBhD6tniOr0V1MBoqNRs
O20SBFpAycAoQwre5Q3wFHOmVv6i3dhyXFnCqs+8ag8n5hDNwdD3Vm1Xoh7I2psv
4R+4/nt6SEGjNSaXIepxOUjbe12Q9k+W03LADwPF/aafF7HIDJQzzw50ZFUlz8BZ
6A/BEdotwCReIiKMKqQQ9dEtdsfiLL5nCj17YAgqyHuyjNCPN3BBRZn9OrsTQyae
uAAyzNuO2bsPvaelSVfrl15cWeyyIXuN2XA2O95//l5vyKeddF+Dk9ZhDFbu0Pbf
p8t6cSd9JmBb+zqZ6apaveYNEqlil/CgKFTcSqVh8i6fwC9CVxXLqZc1ZWI3wGfn
pQeG6JOhKkLJLgwfuCneEJ7mYzFU+B7BG5y50HgXzkXH8IokK56iTnuGHStWawNt
ydXklg6y9VP26SAqx3cA6ftUEzNEIi9BvlQDt7wScxtBZT6xu8zkdLPHRS8hPyuv
CWUE4g66sqUpcxsQN5MDmFrOCIYMn59/nuYCx87usmfF/mUcqHFBKAdGIYvIO3/C
atTdvQQY9p7+Z/8wpuSH3C/5zWUa0Q+9o3KnurHDOGhYfqCiM37S7ekRk+xEq+LA
uP2SDGvhttC10805DqgSDGj5QzWFOFudNIgVlCje+p6BOkFdSDs2RGgR/C3Dk2kt
PttpCEilvrVw/tpvVXRZANiXRtI4dYKSCm5GLC3lLKwnaJpIUm2cmnJUexajpgwN
cPzsFRcWiOII+AxMs/nLbdVFCfjPL7TkbaV3kJ2ZnCuphH1qgYbi0L8JsPUxKS99
gHLRgnhCRNjhkJmWcZ+tgyHtEoWgXXqqfvRT9L8LAXTs+EGFC/qY5IEHCFA9WlYb
emMeAW4YLAZelwXBIiPcpX2poCg8d7DBRpTsSz+xuSX1JyzVbZJBjFZSoWEuilXL
w10Yhz8UvvI3PsyOPIwxLmCnbsG9NmBjZNeKesy2hG51CXZuBEsV0HxiJy9b8dOy
M1EPNGAJvA5ZCgoFvxpQUNzyKti91wigtfjMtclR6+zf3YVL5/GU7ZkrFci/xbwR
qG46qNAklrsHsj4DRyOYB4T9sXPWJ+eqlql2jix/L4RkFY7dmHxGz30apWmK3sXB
DYM4StsBAV0IuQSm3C807KE2IKCQieRvdSYWGgoBUcXvA1IdyZo6V44OkobmDjlk
DFqvy4JF9nJxD+Af1Jcbexfnws5Jtu0K3rTr7G48jUPfsAaCT2F0hiex5s9Z9Mqm
iS4iGHQ3ymVNxptQUQ4l0LEuE19sR9Q1a2uA5TI/wYFoOOpoRp/5FhjgeDMTuK4c
ME17YLAskPCt5igL5+JorZ+bk0YT9e6vvDNSSzSzREw+9hIsOza60xVPRPLZtr+D
LLuuDH+xbkVeIVDYdjV7y2E59iQTsbikh8PdrUHVfuZ7rQisByVLGJazRB75ny1w
rOz/H/fJjFK7SM0oR1OvzNqAkZ6w8rhCPEZw+w3zg5oUZR2hDwJSAT4UV8+ZtVXC
An9n1Qtj+vtq+UcIpxYZnKaytwEnLJQMh8RTcQ6vhSGVjuTNpmBnaNEgbyU+NURz
wJMr7a5eKJZs7XD7ufjLpOdB34m81Hx1qbFv5TU8BGtJeu9mBOqYHiNLwqig3QmN
GTqJMdEybnEOWONUYyo5fQws2uO2uiFEXW3PJ7XvxJAarSgqwX9hV2x75UMVbGr6
QbESHgfnkwSdbiXSpm8SRD8M/Zg6xreePy/SZcNsYK0uY7r4cTud3uYQSJLbL5bv
XBHbgUgA69JXP4pCVpSJiH3ZigxX5jE0Gt6ml3GYdnkf9pxwlJtfqiq+2bKG0Wxc
+rwvlZwDDcjckHp7CVgwJ2EgEPCnW3L6PHMGeKS2ATe70LID/48g7+uBZOWz6sIO
TDpavbg8F949kmD11l21+EMyrf2PORv9MnsRdrWE1sdGqvcDp1aMJtZEy4+/IBOy
wG37ijgo6vvCMhpoWuITHyeLX1heZn/4CoK88m+HbrUs0kQe1SesOg7cvZCZ+g5V
PAe3EJN2iEPXvIKui6D4RyeO2C83/2gYGVhM/1deullmtQQPsTKeFsZn+8JChLhi
AdEj8aN01rdgZFxNyHUKYnd9iqiVEsQ5q4A9+Fs94fP+TZQCdAFf8IVRk/2mp7QM
YN2wMF4CGTswPGENU/gYTMvOPXG3VlwnbrIUL5ga2AH9/GjMjL5raWvFuefMWsaY
QzzXB7p0KR93jqNsflZH7GOvjIF8RPNhMMNEQP57cMLBQO53HuAtOG2ECI8FWZ3y
tejOPXKewd+WOW1LEcTuF5euTm9q0lrduoAdJ7M4CQRhhIgJpd2SThfQxj3oRotM
UTR/s+rEkiTJflSxZQLP+T3aTbuezBc+wi6Jh2IOFfM2/bQ6Gn8oJjCaIwH181ib
6NnfjB5toHnV1oRx3yznYZxhP8fxto+Rsxe9sczoSaDhbSCwFHzhzUpESQN1ChbF
n/HsIVx7DBS171j4Ch8LpnQO5arajh+lRvW8mIz0OqAi5+aOoB+3lHj3ShJHlNgu
lMpSpM6Gi9lduHTm9eYO/eVMulwaJl6L3djV1FSBjXlA9/aBAjBdy60yY8RT9kN+
UMuGtLgSFpcnnWgUBb76sHsFlaXmvqhWUPdjNjS7kDf460QoaUS46FmVA+hSYSLq
MBMmQ5TeqYLSFt0Vus/fqjfdBpPq1T7KiEVC1rtcqF8j67I/qIpdyk5fH2ejg2X0
dYWA3StOokfbNHIOBcGz/iw7UOcK6ob2NvHLoE2+q47lzU3/+KuqyTwCdwRLnI/y
MMCrh9Zr3RYOaT6SgtFK4fTa95NKdDCbTt/AlKEO+U+QxM25rnsxK4qXQqoF1b9l
nO5ibW10Oml9IoplbNTnT1Zvp2cdJ3beTfVDDUNUKBk+EtH/ro5xxwGzYwWUoXie
D5Ju8DrxedPhT0FA2CW7C/Q3mjkjV8ChSQketANQ5HbA6CRYI3N3155lxbXx9cx0
6rioutKmjQNoejE1rBGgQHuKCHAbyBYxT+LfudK8ImI1g8wJvJ0NnEzfGIxtRMIa
MTB8VS73GE03BXwJ/mHbYLDrqCJuaZMNhEGKISzaiYLcc83ZNTWZaoXomzbk0JkJ
rGSpqMHmfzDmePF1oGnFrvKa+LJ/Gq9NV5qSxZKNCugEouoo9mOwVi4bNSUl5ghn
8dvwkJkFBNBdSkfWzEyQKew2IRVW8qt0TxTkC4tKVrrqKRVniT0Me1FTdRSsj+AO
V1rl5XoVKWuTdHd50JcZnw==
`pragma protect end_protected
