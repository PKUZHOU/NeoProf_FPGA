// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
BBnPTmBvAeWqpdaE/3Yjb4U1ckvM9DH6mnMdErvc6WLYPpY84lhN/UalnpEjrE3UIfFKtCTrb6qj
iKC2sSU+LrLOERPOdERwscTx0OItDUpDKfg9t1/6G4GtPu3VEkr5l5cLZa+NCOzwOplVtjLhx8wM
zNwjMpjTkCnoEdgJP/oC1cU+zkfTinZsi9FA+SqY8aaVUy0x1p0VChQdtlvLu1wolqppnix/pQOZ
mvgkXNL7tJ6BikX5fRU5O3j3k538L1bs0nv5V9tWc5A0o4+ht3rtgqEU5Utqqch/gR2aVC7fzoMV
An8GV01rC0F495qgs+BMLES0wCCJF/bvD9wzvg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 22736)
wesVG8d0HMcA6D4U8MaP+5VhjEeYM2qs6Adys7ZEaf5VZTFXjTQJ9LRRD3lhrNQJH+aQzpw9JK+l
YmhVWApYn+S9QKRfrMmLMKUQthFEHlRSaraaN+2EoUpX2MahhLyvyuC8AxFIZBPkcpO+RaWn2mLb
Kb/1Xj8NB7wlqRy/t909gUNhGM41VirHaZKZIZItrEXGiEduWb2vGZ0xc5JpXx1z66Aw9qSue94x
UWR4MHWPatVT5Hn0jjI6uUaX8I/jvNcuYguF44bbgWhAXltj9erDBS3Wd51Y+GQF9qbLjg53pPdV
ExRfu0L59V5R+RNL43Rr59Y14gGWsc/KOr+nQWLJXjfIlCQgH+WqvnY4VTckCPQhsFsDYVHMz2x1
a1Po5aRmpGpgsYistqxrMD+01Z/HGLj59xwuhZh1tI363wE1JD1ejYn/usESm0o9ZWG8m8GZ75qM
YjZpxzc3S8S5GJt9tC461RjTf9ukayRl1oaYz7baUmioC4t0q3B7O6IebJqHM0Lzp46XKo8OE91h
joqcqOD46c7+GHDlFrkWlpKqF0y8feapNPRtw1gLQzG4bP1KEEZIIW8hw2WdbAmm88NyhwiW6Bsz
fVx92Am1q5yvBxX/0O1dHBojrgrHd2dE+HGkT4IzLZBP3VFFkVGm4mkIL+kYcei3hPVlXiZ3FZr8
9FsgZwH2CRd4c420rqBamtWhGUqU6r7dOzH4nVjIo2ofvn4idxGLQiLCvqDCo+lAipH2eMCoSOlF
tHiriUtAPCvEkG48F6YdXFALaPp9PkcsIwBw0n8LDOHfHaM79dn//jCbB1lTIJzzPob7BUEpgG9/
jUQnHvveBbRxCz9Yo+7UP/xI+F68DI9WlI7VyZld3tk+fDrjYLkw0ZVFqXH1gYo8WGF0ULeWMCb3
KIBACMUy6JHHinHNaUExPsY/rCkcz1AcCAeIjqeDzMiWAQRv1gdgDWOI1mTgEHlXMPMNbr7No8JV
k3xypuvyAhBINs0HXT949+NTSX2R5dCA3D1YeqV+pg/pI+tGXCR23i9mn4vlgGvnwuD/nyzgIiQ9
8ZHuLxanNazVW37L0+sYKIuGQoT8SMGg80j6QeUkNc72kvFhAuZ8SW28fTesTnri+Mh1aK4uC7Zn
s668oR8lVSc2A8DsNGH/zBOVMtEFIGThNeumoWLFTMgdTS374sCFqIh71/egUu/Hv2LzHA2NcmXm
YAg3RH1tqlvzz2Y8mXue8TQpDlYq9whXkC76XoLrV3jp3oTpJcGHyXPfm3AmQ3enyV4rmx7wa9P8
EQcrKBDeuTCReby5Mo5McP7HHbpBYyLSGEjn+CvHK8TtnL/Qa99m9+36xBZzS9QOTdRGJSz3/qT3
LHRcXCyq6JZRTGmZAITBQotQRUh7c6l3jpHH6B/Etgg0gT9P2skm2HhOA3gaL5a/fECQ8Alkq6u3
Udq25uQX83uxME3Y/R810ZMH677hXUlR+V0xQ6xZzubq2PswWFhoAVSAX5PBCskiTlvWlbW/NE0A
DYrYoCpRSEs1QhUt8aHKjulIhjmxMgPudDtOCkkHUGST2hCFgVtwbiMZ2wl+8h6EZmk2faWesP/d
xP5zMc8GW1HrjBMP8Wm/vkMWXoexNKDKQVtkFahTkxW1/tUVF2yAjNTiCvo7rJlQMvbox4UTSXWL
UleKROIUi7SqxG94KhJ5hjLX2ZOSKp+K8eX1DMY4EYGgbEYqcwRW2iwvmkwxHVo1UB7pvP0sL27S
ybPlc3KsL9uCavFnQ/DNSxzF/D/mNjAWTlbc2ctj7/nxbffY/3Rlw/19ifQm0HYfAO1UTlBJzY9c
9L9tQCrXTJgyQ0RGoTC9yIqceigb3Ygrnw3iOH7s+LTroDykiKKT2XuwAa9281MXfdNvFSoqIA0p
BoLfV8KXnCnJm/YruwnqObWDmnthx+/EMr6YCWVNrsQ4qU7ijbjYN3gpZdKgw/hlSFGG5h4ANZlW
jmni4BKqq7P9Ksfu/Wj9ZajviFy9kBx3/BIgFni34AnSki570j9ruxJZeW8VAEJCdwlBNqDDxMVv
Cj9yzfFE1LeanyyzGHmtSf0e/zJfYuA0ZCKZxNVKpf9tT/a2SmECYo3HBaoLIs1zIo7XqVi0D4ur
oYHB6rulRrKrmMioRl907iBO7zE4XkOc1B4Vjx1JVVouokD5Ff7GyEDnkKuAwVIM5Q3YtWkcJ36/
OTqrSlNErB4DgH7itGi0h3HmDnEMhqOT2xpZ3H1MzSZ4pdxFPtXZ7az7qVIzVwd6IN1L7Ta/7ymT
QEdmiTdgBskbaAU5FLe0RMYQIyEf5NeBsrx5aiVrPQvy/wFf6c7a0boQi/G6ZZhTOqBK7SZOwLHQ
UXlSTq5j9mfyhJfxpQgW+CYykgTx/YsJsxBE1JCVZQq25pAxA/upELdJ3UKv1/MJVXxxQDqH6W4m
4zUSW1pfxNcd/EAf0pyyDy53FXB23v9zkHGWmQACnB2iA6K6nAQcJt8IV/qmekDBJymKY0aOwSze
PrG7bUgSMArW6PItFteKgS0csy7u3DdaaRbOCcsDH0QpWkaYKseN4t5uPh7OnRWmWknwWDCgFmf6
b41LxtnNLWHNKzBNNeRK298FPLnqEEA1fixXRnoLJXgR/C53Pra1ktNyVOihJrQnLaE5x92LO/LJ
jbbcFbYgENeyo4HyG0bIQcQifrfBjify3tfTquj08fKf7HDGmWo0pUSkyk7FxLylw62Z6a/yCztG
UakUtKRdjs+izGxjFgHWdWNVGxTGsVDmIDoKWyj7ND5mD3JLlrwH+PXq8OwEER7J9ji80jA6RaDq
ssl5vwai54KNj3TILeyEOUTdnQhecPpWr7adeXWL8N/ZptViZ63lxUC3Q7nIludR3e6So+jBiPjz
doi/LxpQKV6J5t2t5+f9JPjWs4ygZg8AYCm6e2R6JxFcjDvMpwqFk+bFBdsyFA4qUJZ1a51rJ7Ms
uX6jUUH35jrrzSSbT7KvTAEupoHmZ5knIhl1Z7I/Kbe9tKoxWTDZ7g9JZmBv75rWlsWsKLH1UOs+
WyJb5r6/Lx834DNVE8xo+ZY4hr+w5fPN/IyuN0jf+ZOuWOeDEDlTAuqZNY2fX5tNJym8N7RWm67F
MTySHfU8yeip78iFPppZW2Aiqi8+uQSugKfw5feVWTEjM7gnmkPf0V46FPjzevqmryKk9pG331Ai
fTp/Yk1r8ESkpslaYmregVzvS0e/LYgLCiVOB7DgYnpdFtFEvbgDEV1/bwRFj1P1dnnO6kNy5qUx
0Vj2gs1coT/ppMWtJW0wSXlzg/smnYTEcUldbI6BtzD6iS31j/y+R2e7rM3MYdao96K9bjz69H35
s8hKzV7nrXGCvD+ejIq06Du6uAvuJ/msOjVJVyDpVcllkxupJQ5NElhZQ9qDNfXmiE5l9CT3gt12
bZoBBA69R1TdeKJQdMMQEO+2BJIkJ3T32gbdXkoEwSmkKfN9XYI3bLUVvm85OrZx/XIeUTVLiXiG
io/f/NbgFBewteacL1qUiCpRsMPuWfM4AsO5I4NvCI6oUc7d4INMIZBJgkc0PiIUBOVvqMrQE9Mn
+0ii4L+3SZKfKfr9gGmJww5bii7f++/p50DaW4MtpQr++ipJGCHnyEzSo/YqTuP6x8dN3qQmBiDK
PjM/uVkYl/BQ9Zkpzg2+fHxYEF/9HhZ89tCKMlEcmfV6HH6MkD2HycooC07QLNY2uvfl/U5qIPah
ImDSHpmSQFXNdc8yZE6q8cex3Y/a/aIFYShLfb9/V92s4Enxf3Ip2vntqaj0uYS68abQHA/3nbcQ
JANot9Gdc5Ovcs3t3D4wpGzcCIAYVnJk4GVJwkqAvW7lNPYKXB5lkQz5aMXcwUK+ca/4ujNPSqWe
Kd0k5p8245geUJ5nwWNMG6c9nLdJ5zrChczahxT631BjfOpMPalS2bLyGK6LovZVGSnteD0omUuc
v/LiwIcmRFbOzVyO+Ht8EKDi/qIY0k42W0AUnwnePG4xaJYvvA+i30N3vNyGtiVfrIW8zz8ct0UQ
Bz5WA7XVgC13XqtmFMvMrnMrkHMjlkyIbTYTjClCeItlS8Dpp1RdyFRbdtBxeY5EKoqgfc52LkKN
AZV+6oXW1wH4j+bn9FMsIBu0KovuY8nG60BzzVkP4i5JeDsR0WHarq1t5n5Q/a6V61vLfUOYch+Q
aGeUVyrsqzeBuDOE45QgfJvHNZnbRD53HOdQ88PZbbP++m8d5JYYJe4WHDHgczJEB94F8kv3ZVsn
copxYDzYeMP6jxzpbOQSSvP6e6B7xkHcRnmsqu5hCQ5oMX+KBsUYWs+qPfSwpjVU04kFn5SHlAor
KdktqzYSRJZRdiDeJ22bXl4XCuQM3gVCkyt4rt0RN7X3zQbDapdcHQJ/KL4nObAjf/e19v1/y8kt
UxRZofBwZ0gVYN80wtmwmqGqg8Wuqv04hL8r8tEc27Ed17qMjzZ55qfZccJUoLd1h+Eb6AfIfg71
YDvcW0tUEDKh3lv93cPoRHqrFlgo1ccDb9+Xuzp8I5MVwMBlYRwoNsNh6hcwHJioCwtsfyxJQskg
DgytTj8SIt/SGbkmlrdzQHjHY5+z+zf7vf4IPukwXsaF3d2HE/sT8VfpxsqUGWK66YxQpZ+EkVK1
a+ZZmdxeou7y9fd4njxiAyeqzaCRJ9eRII6W5cMk5Z80/k3CE/jv26ad7XgQrGO+35GaSTA8VQ1/
z6KwLe4NbFRvht+aQvPEDXRD3rNI1x47tEnNaXaCACa6DNxOh1BRCMBQCyzgvukyEiZ9qXAGPPLT
a3bRCYe/gdxTsku31Yk0EMBHA/7CWTrBV1vsHSW3hJOR7lwj/lqIfxF9R0byBzShgrpnOhr29qra
T78FgtOcMSkRhOs6F4aj/A5daFORNAMLRbJYR0jcm7hyBQgA6r69JMHqayHFRqd8+/08yMSBTJv5
IdgXXWTalRb4jiXLyfm/nrSAGKrMz3WQZonvl5TBiK97UFKiTvBfkU9+z9b5n7gezBia58r2PSPD
0quaGN7/lQjWHdtKTsc1ZCsU+l6THQ04cRU1pREvQ6HBWLgvC+Qu5iBARc+DiuJHEhyROQworkXc
etjngaAaEabbhRWZnTXYOcKx81gbzHUWD+9n8497stMKxNSIYi4yDExRNP/UN+U1uv1BVhioRzLb
zDEFfdbPK90KgVpXKDs4b0o84PfN7oFwagUKlp3E+1WBf/AcvqIWTN1IW21n3BO+zAf3UNgWg91I
D+OAIp+i1PzphXzw76Jc6YgVd3UgmWHEUaNxVSsho9lGrywnv6jQFOTCwOEiEZij7AFcF2eEKV99
r+raBGLIN0LYTdAkwOibHjOxnfplnFRzEpJ4fF3yCKpk2WbpeYvCAQI1MQWoqctB+uvTISW2Y7TN
jloC+UzdosaFcF9Nfrgb4GfWbXJQAWcq25XEgx0RIqUySzq7yEi50gO/wD1pDMo5jlz+5mZKbDTE
23xtXBOkd6zCLaUh6e6fVmu1bqcCRN5+ruNUzWivsU9tUAJnRboC8/s47MTOoAfP+/4EzbGNitSV
cg1kdAn9+oocIsjXwN+gynstdh/7mWjsBT2/AWDYj+JWmpCX2HL9gSHbWT1Ab69/seX4NUNuEZvt
n81+XMyTFF+mI+FxNlsX8kUoAs5rbErFcj7aGc/cc0NoNhlOmR48sNQ1AvEe8xLwY4EpyKoAnGRA
os20IjZiSGHjfRWgYUAlxr4nPN7uVgHRtcwbk+RkwcxoEFCM53EXaOm1ncwuAFkvIkeM/YP5PmGJ
PZRH3DZXwc098NSIjRnPudhTF8ALVCnU4nyUBOcEKrjfh7Q2J6upngXvHaL/g2+xSG8UI6Rgl/mD
Nmb+XIeWBvEdyC4CgmRq8a9vueJT8eWl94p32O4C84FLyIHFBMXBYAPUXjHbGa4Up/zqWT7v3qWY
wLrzLGhYyjufmHMX8u6MDwzb2GS6Xo3gmqBPPWc3c2slDG5U6F0G9t1e49Y4C7qqbOSZicO6jhLc
66OsfnAdemN6EB7o2mFuMLxaTZsgGlrblL5Q0r6+jy1dCdzRpJdmLtM63g7JmIsgVRhWm8nYgArK
CPMHASRL5sr+F/uhx14rt9iAEVK0rdocGwIrfpwwM36M0twOuSEZDPkE7G2mejY+QqS6QFojNuMr
6Bw4P9ic/UdFZAQPS7oXnKgPzuUDr+v1gw+qMkjgRa0aDYil8sSUPaD86GdoX3SkQ19UOCYBHLDI
v2SxIKyRpbzswVcAKVVZ0eTkkDg/BKHiL2CvNLS1W4LPjIXW1w/Svhgi/hVE4USu6XjyDWbTzt/H
bLqgBxqqcjre2EiGQezZIQhe/xKytov5BUSh0kFPqwatE07fOGKboqhNtQGyZi2ex5rwpoTR84//
FYM2NxsnwZKjvIThZP4fAre7Qogd6KYbNadK63qGqcGHtua6xNPukPFP5pvo3GNf+QO0q2admLsi
U5Keh4g+xbpc7a3ILFvzXWjJ1AMGlARtUJgxTpJhJDEZg3K7p5lLXnFzzIyfqc14cpuvL6NOKYHQ
11hbUw3McJfYx47O0cw/uWG4PN7NmBn4jQyytItAVDzIl89ii0LPcSpIozU8tvaVpNx8ECVisRF5
hdScnxmRggUi4UmWKzjMk0Fa3ZMvkFdEPX7qDScD/VrOHaP8Xen+zr7h73xZqOTp5W7QonuOZfM/
F3Wn9T8GimRuG0G+o3++VxAJSmMZYfWJNCsBev0qsW/xdF9memCYodAnVgHx3f7otSsIXGJhMzg7
0jZTURHRDGqOHTFt3fzd0Eil1L/9WAAyll3CoIeQqdnZYB5ZDMxbq3fN/9BZ8z7WZhYBM4w7ACbo
tm6DRWKU7u/d8jmrpheuTGXlwK3i9HKTZczKuTX1+kUR5o/QBOOrK7AVg1lFfMfJuWwAsNXjTzmI
tFzliyNx0x2tjzzJ9OUDqvXybH8Lw8lo+aHC73h86JsuUQM2fUt6gVnpbRFWt7N4xOzsnWyQHx69
Df+du6pwyY2bQ2lMb7bAHM2vCzeWaVvN1JP6Qi/g5wOmMBxr7eYDdQXcCQJ6oWr55yYnseISRcXa
x3Al/whNXRHNZ5ab+AL4m0c2MQw/2LEkTmNFj51bztLrZVTT2IOX6jsJ3SW7cfahdcRSgpquE/OA
k3rc+gO5cBdep94RIa5O8ZAetoUjO/wnBsSP+5mv4+p1gwDSZBMfVkWdzaQ+Dftj9VMyoYRYEhZk
sDDzKx6towfKjd5N61R1XYvj82ktb8TZe6uHecA0k5xmejhqZofAHkHAHACXNZqb4ZKOzOAzRNqO
RnPHfApL4UBZLJREDm2HP8JMeob/HoFa/xVAeSg1f1Unv2exQ8Jd/Sf0OQnwzmMe3F09bi8CfKfn
ta7liOw+TukyY4rPEHcG0JSpmA5nweq0Wvd4s/XafBgn6qm0vuDSFX+nEP33+AX9ncbrviSm1ofv
1EMMpTDgB/H9j5bqfcrUocesb+w5lWrNFKVOI90FGyqWuPap0pX6rmORax04YZI1N14iVyh+ToJI
RieehNA0VY6QKRq4df//5c3cc8lOjKP2WNZ1wtn/e/otC0i0RNzXQYJM4QSTTNi3jpna6tDf0adw
t9NTfIRLxJHS5H/0kw6KdE2JVaqq3rRpo9d6zPZNai0sNVAE+frXkRev/3bgIdWD4C1m0ibaTQ51
vZCrKjSfbUKrth8KTmR1CXq703JL1yazSIldfnpdUoQb8ZMRcLECUvJDpB22Qglvnnwv3+ejTYKr
yYX7uHuRz9+OxT5Eysg4xZjxb/1eRs6fkkBi0LKMMIFKnzpKQSiqiq/jP+Hw0sGSPKWbXKNrf+37
1WX1xhpzaiCa7X2YTVdFYiox4QtNjSbAJB8/y3GmFPugCVLd0DVD45PKlIm/SByvDVWGYI2A8L2a
l/uEthuG5aSH2vLS1/OfC20kl0QEA5+txSDp4c7NpdVeLTdJfVVffTxSWZy3fO8VKQE200gD7GGY
EskUSQipy+biPS8ruIrh1gEq42CEob7W0/OKrMc4Ez5tIUp8fOSTRR7kgXTRLNPoES1KqMYOmjus
wgMWCNFKbe3qH2pCbajQEwu07XyRGZDbx12JZrPfXYlAuvCVg/j8amYKFjXhEf71Beihh7PKh7j3
4mcf3ADM5A4H1LmSBMHK3IULWY1ACJ+9NNPEDQHAMEhBgYBoS/EszV0OfOgR6sValJ3Xoi3Cq2Z2
kOZ9vSR7912tt6uiAfMIPQXZQEMAUtBhEBOnibS8L2WaTaGI4+4MDvUIapWbeDcaZQ7bDInqLQj/
yhUn9Bu83Tg/nVdKISz+NQ26UjtpxP1CtXKuIcvOmwWGIBSpvusEx4TTNoEPzw5ZLc8YWyGz8xxD
4pMBFPjdZFy6MCUM2FWBdjK+379SEibQUvNZiF+F6mpxShyQfpMByIDjV2GbLN8EDSie8tkYpiW9
xPo80ZURdtnzl5/5sv3dllURg5v9Z4yUljfsZTDUMK3Vru1tTWWyNb+PMcLyQvV7POgMqOWF6bzX
uRuv5Lb56Bl4LaGboiUGJ8JGVtEaIrus+I8vXZmYX9Bh8iyvrK+LfbhFcYXx6IX2gAsZft7lsJ6u
a2sXbwQasCqhdFt+PKVLc43fGMs87fX3ZiNgorUnHnep9LWIrxKUc7Ya9yF68ToFfvXsYW7rlUse
xASSJQgFi2QrdTClw3vLXKBI7W2Ks6QGi0cAo7PuTvL/uTelMR5iSqQiZ9K5eOh24G1XPPb0XaVx
Vi7UeUtBAkjm4gy+f52t8fVujqVK3hHuZZyw76FtzMXHq1WkKxac+eTucVVF0hNCJk8dERazfvmQ
xXqVJ2gjX+66DdNsO4u5e8HI02vjux2mSyfWneO+IpXGlSsOGrQg/ogdHXz5T+l6mMze7JegKhbr
Vh012xIWq6K37omAXnWrEAPQU2Fs3g+NedF0PbRWJIqQ72+FOu7YDlyqr4+fa6HOp66GP1hpxQEy
ShI36PiMMxUJcgtVcnl1hZ3FJnc4lhkWHRooUSmujiOWCSAMgvRDspNb2dtRtS21VqVhEO7d8y9j
Jlth+3Z3MHv9kYz5rPC1lL6teMaO8dB8c8PLTY1zXMCTlvcYpp//exGSAS+ooHuQhCMvWqni9rmN
P6xfQKCpKnd6rM0xlHI5zEv9DojRgfka4veH2uUtkvstSrKk4cAQXqx41kT+1Crxtqf9xkvdPT29
zPMjIa27OdXidz98yi7sLRBCS7+gQdKX5DVM1WXNH9LkXl1cTklczPWdXKy7Vo18oANXww5M8vd4
FomLsHwTUp2yf4PF228xWLEzXz0YguVbxERaO+v76TvuKDJTNsgh+kY/MJT8W5Zf7F8vZ8E3oGh1
W5ra57TLWTCYTsMfPOxwLVmbAMXQC8xqHp71W3w/3LHEflmhrwy1qtUf7DXm1TMNawe0cVEwkio2
YLyv8gfnyUZnLzXpmgOQfA/Mv2tEfteM8t5UqeibkfpV02nXw/jqdV7I+zxy4wrDyZ+9OBPOKI0/
nyt68Bx4EQXUjRKNOHiOhkTt9O1ySjXARC0k8yONc1Fkupv03Y1khg6LFgUjdqyJCVj8xCDnPfuC
GgcLNwaWxoCh2AaX4lUcOMRFzr4od+Va/1t/XF+u/Z7glzclMG1wI/j79++DfSyyjMlf4lHxf1FV
bPmTeDgj0BjJ1EOH3UstjuHMrZkLNE2OOSq871zc8xGMzAT5aHVZzQLFlNcQswNIMULOtip6GFnb
BIhG2ziLs0AN43gzrg5UyY2t51n6WpT6pXsWJpFOb/ptH01r1XbNrsvgZeqQ8iyUMeyc8wtJcopd
kp74Y+zOuVOKaJVsrhIYvUEe0k3Rtz1VJ5K/rE3ePbvW/gkadyvJVqbrNQr7uUBqFeztzCKMacHd
mEvGp7CUwz9FsI+ExcK/89H2GMHG8DdCQNmRrcZIgNIh5hSfvBLznXUQswOHrWEIEpbUCLzJnpho
+zf/MvtCRTJ0Mz8Q+pN0NBicVrrGcxv6EnJrmyC+sqgu9roLj9Fwlw5q+m512cmYC8n+u9jNq4Gq
9XDTLCM7OMjvVQACx6DODBabz211uTiDAb5oTC4YkH/0rS1FOEV7xMGKRO00JslGDNa5KV7GJFsl
ISoiGS+aK/hyLxgjE6YMm3f5gI66CVqryWOUVh6v+IckA9fVGYZGjzSI7rxwSg1pJWWF1TU7Hav0
l8eTfKzFimsB33UNxIkA7ZV6T1BCAQIRSz71m2yJKk+lqniYQxpR0DUDhFgbsVA9E7lTUPTzx/Nu
HTjZMREKQ6HUj9/NPMGXkl6YaZ9A4eWs7nMEMYob4l/cB039bRECLLMb1YJQtKZGHKxKOLpy+VNw
mMCBJCcKcjAxsWfXedekeq1qOE8gM9+z6nIn0y1Pn18PZR1cP23DWzPFVMMwwfMP0VF+zOE4wxVf
vateNFBnfhlhc5ZKto/4HYpE8gawNCxTBvxoYepA9ZRC0GzuKHJOh1ddrtecz7lWu/INXa+wW4wu
bXY9bxiavzBHbsB72nYdD5MUKUEhpccwvzdeka5nXJzPbFckKu4YMu9yZlnH6gLiFLO6YiLS2p0Z
aL0Hf8T8/0CzYcbCicXL5953fdR1koYw/sqNXF8RQ/lu725JTrzMzysAwphsr6qDxWHfyWG4swlV
HnS3F2EHx1k9hsnsvb1YnwWjDg3XmQP5MyqjDYhZMh2ZK+w3qW4QrcTsilKfcAy+XIeY1HmwfQUQ
oayvfTXm2KCdKptY7PdJxhvvfhIrYc8+EcRpK+QqKEbjrepGeMIAos5mOucPsIN3rOKeEzcdyUrV
zwUbPooJW4r1Jo94H+d6PpKI7jD43ZpiCpU4bilnDAIOhG0pMbI6uOHod62s5gu05e+TlJZPSULC
4lxd1PqdV1ospGceuT1kDLKackZI5zlkXGL31UxzCOBzo5EXtWrXww4z8jUz/uoGl0VcsIaSPEtD
GxfOL2EJ38pSywIhewoZnytUcs0phXOSjex2DME8xSW5ZwrMRsWen7b+XCADNurCKxU4bhKYAaK4
Bm4wrnYbcxzMJsWbOzYRqRTYCWPCaEHhLK6GxwY2i2ooEhexRsjJ3zOU1DxmdEQ/yyQC7m7D3Osk
v7qHRbJDZpYP57ZFSjjhpQKSpASUhYZzsMmcfk2WmKR79sAYKYda0aEALwuvpTh0t2aymGggmmuA
e2vbo1Kqp9LosvV2eNGJTvXFY+FZX6xlCyhdHIon1iVkdRTgRav8EY2m0PaX21h0PiWfGVh3959e
KODiHjvSmcqWPS5S0q0hGIaHbUxV6cmTuLpkUZUGSzqc4jKbAlLtyJGA17Kz0w5QVIaH5rZdEZ3B
D/8IvW2C1fmu3GGAWc6V9nVJheiAWl+zG0rvcP50MnO9RZP6/cTe2Vn+fan/F7oLCsqQ2NEOFsZC
QRbWk8T7QEl2uQOMyGOFPyFAKsy/vJhuCc7PziBnV3ktae0n/q6U6zXVLILppQcJHpo3QikIILsB
iv2GBzOf6pfRn1rVd19OKCTV+EAh46Ue5e3zfF1XXEEzgSykxBI4gKtcH0hC8QKZ0Zkp59iMsreO
p0YVMeqlBbqpTIypwMrldGY390zK6boo8ihUC+WAqgsK7w9iCM6+PhGW1dX9XzBREYnRc1Ct6CEc
3b25Wzs94D9mxOJYeso+h8jTwauvzs/gnsqhFG7Qkva9EovF4hpZrbR1VbP5Wl/TWW3683gfWVph
a9fF3MAp/uUhp+LgYSYy6071zFij8JC1bETbYsTjrx4qc59wCXhyL2x73MgtMyVCAfxeS94/apbV
DZLynIlX66eLpBsRkm4A3qfhvCPjYyyNfVXgISzDCtW3Nq6rnIhy8FYKUHyBnYFKBqSAjx+4Bt10
Bfl+w+BTmukM2xQQ0S7Onl3ii4eN7w+dZy0UlMoTZOrcgYngci/x4GihMgKZSptYoFVOfNOEq/Nf
1DRnB9WvJM1eSohST14mGyikLbnapUq/jlQ1RsGpS9Mb9zNCxD4Ni63GzLbscMzcLteZxXJlEM7e
zRtWHJaBzsciOkFRu9Lhk/aUeqbGcHz/hnEynMEKYolZFS9NL5GLjEdDdgHD1kLV+TRGWQIBWtUS
hSIVZ01gFUZRyRtJTEo3QHbWuZJvApzaPUz86BJWp1+KsZk5zIVoC8oNNZWSsO2usSQmGWRR5f/1
Y1suusuKRNZ9pnIFzC4dnZSzp96rahlHwUiTxdEodcxnCriKLAypcKwANrLOjReL2ms4NGpW0pG0
G7cGng9oyrvSDQKFm7drSGt+JALc0Ddh+tAJsyj4l2IrL6KGZlIt7YzByhBI8sw7ddVOMCxOBmc8
nQD16lqS78YRydmrUHiWnaay0cWbCaur/yFIrsoO8lmTH8OeB7QuriBE4moBbLopDAo9loVKvMhr
RHkl+pDBly57jbnjyPm5SIp49LUBIYuQ0R0TlrjC36hCovtklFxU/VuSV7YnqMMJ0wAh8xNODEsw
nDVVVBi9cWqdCWz1x8DyeKg1DlR6gdZconbYPeDK92+2dhb4lypCzkXkBbF8pGiNyiMie9kWz/Gg
IQbWzMXENXEb8BqAB8t3Mz8Wg/Ra6Sh5VOo44kLRw1CjYuRFY0GbzeE0/K7uhagznBB+8zrXky3Z
doEZSZYZyr3Z7GKy+fZottw0R8Y3POV3IFfUacoyWlm1MXJU1TlBHWdjPm0A0TQ1A1ET2shcqiTp
CdxiepkgHae34HaexNo82n45jqfEtBiZZ1kZ5T8Mr5uzkJTW0uRjNblICObH7mZxB9w/QiGe2S9N
OUkR1tAIfRP7faHu2ey6aLas7UERSkV89d5gxpDgGDoQw8QQfyjHiTiYz4Z/HHVN+ZUK8DChkFb2
XqDy+TFER1J20t+Sp/tMMfYl6kjrR/W1m0cA+ejPVvkN3JVYEVbF0XpACLBVlZFGJVmxTVamsc1D
IygR8VZJR0hiVPjHwTeLUL89t6D28u+kKUm8g6jNSUHuXau1uSv+w7ln8G34X3gogE5ndwVlgY3V
InKCRTbOebAMWntmHwsTfUqTLABWQ20fdRuasOWtHCmHWk3ZYeXrq6V6wBikshIAOo4+dhPaFV/1
HNUTt//op7ZrNofd6tS5y1kwmDmyVpplEGQLORMGivFk5t3Hczj1WT9G+oUKCY+DA1l7/rc9j9pF
2EVIjTjhMdnpy+9morQ+Ldzp7RpgvBdBTMUeVnL8qNK1K15rByKc30jIvP50VOjvs2447bKfU2ZK
9TaTQ1a/KLCmZ3HrxRzk4F/SxagapJpllibVUpyQSXNylZIZG6/YpmPu1S7rDDTacOWtrVcRfy/+
Ob75AOaY9sol2TiQSwS4OPx8rIXFSR4bW2nJkxXFRDjjGes1dNQODFvvV7aBCqf/Td4WUHcA5M6H
9k9PHDrl2EgKN7ANvivG6uEoTR8EQt9sYcd1PpzHF4suf2RtvipiFJB/2YMbOxTQQDjJLtdADHSO
jNc+qPtoHsTPrM8dGvMyd2ROGNRqPErzd1t2mOodVojpBTWl08HUxI/IYqOzJ8aYxiNoXMgdpzLX
0PxCETvJevoe4zLtyvEHruGZT6oMLYu9okehBvRQDMwW8Y9qC9NGRFDAVJY9f/ZDcltBg0DifXft
WFDeqwHtmMwhQGsvd9/DOaHUogiCgIiw3mpm2FSGwR01ivLSTymxLd3utbHPVPgmXjuO0vn2vQud
SOt/Xf44nMKZNPf9KtlccDKgioqdwDQYB3Ep8QWVi3jRia95Q3U2baZKtx3aiX0097epo442A/lG
VBg95A29475wLshq+iB6cVg3JHb+xkwC9NyqronHHAkXj7lD7GbsrKldzr/qLHxpZzjctbahCu4Y
QgbsfMcl0y/QZXi8yNfUbOjYf2P8bgBNqHKV0/y3zwReZUDx6orQJC5CpojfipewBrmevxQ1DCP3
WfDjNTc6EySMoUYswKY5qhsv9EHmSve8ucxl5cuCZRGDdXVCSQ6KocD4G7+Qi5LZ8Vs3wPYEIC+x
mexeI01Z8CyOxzYeDYYgdXjcMYmdbnhwa/4PPz5k0VBm+V2ZJyRVNM64i6Athkl2dY5kiYgIuurt
o+b2AGKxplowIr2CtJMdTx65YaMtxcqP+R9CnHZwAGB1HEVRHK6rcpF8TR6yOOHdU49l46YjA4Gq
eCOedgMfKT6vg9WUXO5xGH99L3Ig1hV3AUdtdSfxNiE9CBhCoV+i7IjZkt/Ri2dhn0k/1fc/DxqW
8urtC5ALU4YkfFqkIwKGGNwYyay3yoewUyFLFmSNi21Qv09C60/vWEr2rzepZp7NrGBWxH8K074K
VtiC9kzueiEdl1mtrZWiibnyj248iiFbjuycmFceGla7lLYbGHPdx0Nd+NaVxhoolUSf6XbPTxID
+Ay7DhD4DP6gQZr33XIt4eQIsP/3TVZsiF+HCurSCXt4B8Nv+bJ8XccT8Hf4zaRCpsoMVyA/XDHu
uX3DQgAQMmRTd2ijG/PpfIE7zdQZRifDnKGDPmG0ywYIEDMAvYcu+wFe0j/kH0oe9jcWgCXZQOio
ydJ8dCbv/3GIa87RMVTbcOkMfnzLjfOwui5nTZ52Nx03GjvWoOT0peN+KJLO0Z+kCIgHuQyV2HPg
p+Mp4LH3ICCz998EC6rJEAS61EhM6XEPNLypaLbw4bawPcyTY6iEik0CipZxp/VpPAdfganFY81f
XcVflMonOlprggpvUl6YMgcHkhQQcJAZhUGSCngwg8dOW/SdJalq4BkY2NKwzz9ma0Yr7PLAbQbv
otkOreR62EZCMvLXewmUCXAoMoQ7AaepXiQu5+VD3Cy/e2kWqAI0W1C2Rj//ZcjS6fh3JHMKSZNx
hqSUoemjGHi9t2b4KzbhoBuhvOc4zz/V/r0PYReS/Ru21a48BHOf3+4zhi8nO/3IGPeXRvN0JwEI
moMedZ2AZnGlroLwRiD0zXVcNzJk5Q2YiqW2Oq85irzVmHx4NOLKFep0YxUhRThiL8izMeOVz0Iw
p+R203TLv1zGzDG+u0q3iUOSVkFvIhVDxC9p3j4V0W9GufIqZEVcRHj69lGmZtnNv+Gah5TCFGa9
du5c9IkYP1hOqwGHKrobgXwwliy84JB2/83C80MtK5ad3IL+kTUpA4dT41FF81VFyftvREYI8pEn
ikOETw4DfZTHndRr+g4lQl6TJjM4i0oydtmtR4J8gzyDRIiO9yEx8ifVQ5mh4pubWhmvYCa0q9Uc
9hXVAicP+WUWOq7DB6RWerUFeOCbpNJ/6A58l+U65E7HhojqhFVQTJ1ftz5b7t1VhHEYstY2B7gj
ROa2CC2eWee0DkKD8Uq2BKvLmx1KaVQZMsxPvtJMkCLf1EdsVGUjjbjsL69phSLBgmCluGhVTqaY
xv5Y/iiQn97BjcDp++//9mYwvbUIa2eB/I8gpyJh7IxnHNUnREpIrYFxCV46d3mq4G1LEUZIYI2b
3Hxw0cs3QbnM8OslJs117pOXpEI287CTcwxY4K6o1Q6X6+h7iGi2wolHNUSMaHcE/v1QEDLc9Un2
WJ1qKHxiXUPQlb1Zunl64rF97+y56hn3m1qreCy0SO+nRN7gU8pHMHSvj74dfnldzr2BV0Nwx+0g
Doe084Xfs3++1PQkQBJBVQm+oTn65L/Ybylch5dih04Hgpr2laSG0CFSk+T5n4HJYq0V68al3KIw
O6E8rK+MZVAXb/G5Ip+R2lYH5JwhqOzKji5BeVikZjPHcOaQBjzo5ryuXhvQpMDHcS1f5j518jEq
c28vbeuy1mtgK/qcdX5IoXlM+hjTOyuAyx7jhUeMVrIGZ78qhVUORggIStmWcQJKUWhGlBjsp/jM
RvdCoiI48kRMDws5HfhT/2zXHRHvh2YGsCkvw+NiCxmjWiqxY7j1iiivDL7HVwX5aEQ5USvP4tXQ
zVgs2zRf3AM5Lv8a7CFa8XUZg1nIQbkXxToI0CeiPQTeONLdtV5V4xuR1UyWPCDvivKXKSP61+yd
SZFRc6nhU0tW3ruRat7pos9MImlvClGfj/Xagm8ln57ZDg+0rw8wr90z0AODcQQYLomrVjp0ZGjI
7U//PYCMaV8ibiwUHeKt2MiQjs3f8f/+azPvBbnxIzHm/qNyiIe228XmNTeOtU/EQKXCxmvt5Xd4
/FepulKHvMa1RIyVQqUUze43x/tMGx9HMrpn0IO1gvSP+dcnUpR8Q5loc3mIo80Xp61Mw04c6XOz
1ArvHOAwahxszOUNJp1YdXGsAI/j7oXwyeXdonFnlXLa4bzP0OmorTRfTjKe5SK3TNjaRS1wLE9t
1QctaVDxf6Xzm1CvVb4u51RAjP4v6GcQ//rv2f1kdbGep3aOFPTxdqd7RMIqK+HsIQrd/DJo+rDP
q+HEYr/IHA2x1z1kSOyw4e3EPg4RjHwsvc19O8TqptW7M2wZLt/6gXo40sNHttBu6C/1krWNwLmr
SSVZ4CYvUmu7NlRJYdd3JkQPVh0lRKwLPjL07qqWH1mHkF6JOykCxjspQt+E2yPtVP95vjbIsy70
HLuUQ8/pEbIeDpCCP68QzS0m6IKupZkWNx+v9W9QdeoeSkpNu0znBg2n+1Py3XsbqjgT6Bu0BZEe
thHvMXhlgpInKOMeQwpET/M+xfAySHRP3fFbR+I90Ypu0m7jklPgnrVY/sEp6ClzWR/td51vrZ2o
GYtJ3SIfqtxc4rabDMd3OquAcoYIH2LHR+JGsbW562CRBNnIK0q2rYXu1of9CtcPZNqbNEntcDEn
IzMOMMAA/BurdwUauN2Ttt04WTnyDm++EpRWbcOYPAAww8uv5MycvQm765LX1m/6uowW0BN6sp6k
O9Lyylrc8VeQv5cG5h/pnUvEStKMJRMQGaU7g13LvXRTQ3zb+RTMglfzxsPffqaVKvHI/Tqzuc1O
9iUlBZ/K6xBn5TwomZtgFfdtG3D7sdDFbXWXh5vI/EucPdpSSCK8nGplhErs2mJcRCpD1hsSzYEL
KNuYr4QjoBo6kKkG3vRqDQ9xCGtIjgYIFDxcqG6ZjwupuORmaWQEuAfQkPmw/xXLzsmNPhF/ijqQ
mHkzl1t5HupatqGrwEnbHLGHcBhqWhT2yZE3Cnr15N5INRx32N5+vlcgm2J9isnA8AWm+6b3G/OP
Tn31t2EW1wHiFHL6JAxZPS/byY2P/jhdUelTAWFY0XosGB5NKXbjN9b/CCVaHg2bY+GgOqSpd5j6
8+D9ZO1WsfdNZ2O9pKEatSmBWCRNUdJR8Vt7QLvmXGiaPJfXeN2wkIGFOBdUMkEqPOuE4a/ZC7rw
imuUnSXZRLtkhOOFxcHrt7Wv1jdQxkgjh0deFiJf8D5b6IhBG++/fWghRqEP89R+7fEo/z3JFzSb
xDuKhXkT1pWnjRKeq1Wbzmog7OuEWeVKaAhIMBQCM2cpRKCBnBFjfuSebH10KZB0lYHUsR32qNV/
WLVR/mBCrM1bGIwjyauP5h0Vs40mt0WGDQ1blP0s1Ur2Vqf62zT7aT2Hp6DBK1lntvd1j1dc2jpg
yDSFPHjz7mOLPUi1BUZu4G9gNPZMRPdh+OKAcO3FD1pupjckA/57HKmYnoYaAfLC6JCyhm2ebgKh
iCjjAnT79IeqVproYjRCfpqGcrZHKc32t5E5TSZyDo+fFUsjsDKJet+yRnP1kZ3/IFX7mW/eJHxx
Kn3V6tGd3UUVmoI3CwXIwgVS7ZI73QiZddFGdOQKzchwYYO4BNIl0QJ9E0ILaswcmgAiovyFn5D8
pXlP/ZMTnG6k98DmR7s6XY4IYJtZ+yHk0agzafh0xL5/jLo6K4FGXmp6hc69TwavKp7RRlhFPH5B
bzFg3OHOlAR59VoKmQgPJrnNGj0Z7haHLYBoqtpBSI8J8SX/bSQ19pV2bHeUVAV1be1pax6pPRj2
GeOBYgYCU3fJd7fTfHYI01Hsk79RNQMJ+l2Xb4NaOYPa8rGigPJuaU/f1vAQJUTsu6dTzSsGyPYc
ffsDqc3/6r2sQ5/f0LoswSbkIz8IQNnZ6BZrchZCof+RUHpGKOsse8ZZ2juIUzR2VY46PI38Es2o
hJEtzH0UrUGBE1hgUg9/NcvU8zw8viVRSFX5uv0D0Tw0CKKfj1Hk6+vvZ8HU9Tqis2bmynYgCBxJ
V8dZ0w+6T+7xr4HKo16RPgT0b20iUzygq3FfTIXxU/0O68QHuA+HYf0SLb9w+gPrxHdDybLqwI1+
nrB/eODM7G1rp7pPV7u+VyGGKbP7p9ESuoyWX+Je3EGA0lXbvTJV6Z7f325dlG8EILa0+KuhvGz2
NwFc3rgcL8v8PksBYYKS4cpGeMEOO4Klf7k8ZCo0c8il6LhsI30D9ul1h346DMtyj8z0kXLIhYcq
qutG8Qj/Gvk55/eF6wcqKPl36hnjLZf436cSTtB4YhMHMDQvv4kYyxWQgbXYZwa/fDnfHYtdqhEI
FTYv0HFgVvVPDVem5upvA+CDpL/9B35SR8005uDPpdx2g19e1Q5nk5auLyP1Zi73QJFW1s0VZb7x
DKG0YAdoX6TXBWalJ4PNZMEtk+RpJXl0sIOKXzpsUxhlXHnVmsIrqZhnQ8x0tiE/d3TLuxqmtVt6
mPkRTPDW7d3W7rc5Z8JVDIeH6ZZ9HfBFprEb2PQH3ccvKqL5k2CneK4Ucap4maKl1Nxp1Y4k8V37
fZz2Ee/QbJESuSMsUUZh3GjaZsUQQrP6E933ahEunJyM9iZaSuR7oj1CF6iqkYz2u4PdzDwuaA/x
Yh+/8hxuiGVOxsSCNdqnutGj2iPCWxJ1nGP4VwzDCKjvUfNKSCbiT1wD9MaQvoNeI3HkT0tYhpOK
Ey88zVaUFkQGZkBLCxdZthsK4F/Q+Bx4Lu2WMc7K/upcxZ239Org/D8ZfDDRzIIO9e2aRspna7m1
xDUQ2zhGaV7/oY7nMUiOb5efKMLHaR/hLy/k5QwvrVEJ0WBy1bXElluWVvaM9o0vYUw5WNQlL3D8
S9UMKU2PAdLHAMO7SiVO0uByodiMLNP2mK4s3j9R+fZiWdUT9MqB8Ihvt9x+n3xUX54jUuVSGmYa
k1CnXvc6BjPKBqXgGu46drWDjwI5LaRENbPGAmyhCGgjcZWYFpcaDbpyTrqMh62FzegkCxhTdR+S
/TD1gPqpuy1OOVRph65+hUVmzZu1hUXP4AXJbwsiox0BUuDjit1QoLXLoqqfaRVejDwcMKievHez
k26e9wbS8dplsWCvJJpOlhOfUaefm8+NIw26G3zKqMNCC4OpO5m7U1GI4jQb/f7wTB1qtuctDoXj
VujenZyYFCouRKKxbtIzQCJODI/EM4VfLqgGTX3N7PLVFGl8F7KIcx261kGiGPzJnw/PYqg955gB
ATCaY3MMos8VH4ivClqNslIgMZEkT637TGHMTjAOs9C+vVTG5CJayMnlxSlU6VbhiERgNHmfohmk
7PsVHfsWnRf90+KSKXsC94FyOzE2ZPvewdnI4Httr1KnMTkvP1pNsHF9miTQ2rO/jHdnHi88sitC
TehlTIm3iDnxCNEplhAR1bHn0uTzkEKl5lT/FXqCr2e2qaL6dy8XJZZWOFqL27/RILcw7b/SfrtU
Q8dyueVAyJv3ygvuU9sW/+/RciasopiDUeAVF49R8HPl7U1DF2bgQJmEm3+H/8mUMZTPfnfSoo85
t0GoOM3gq+yFlvPHeqefOnD5GyYskAABGh6Oj/wcmQBTMNEQyEb0unC/S7TExf1OtqjpSd7nRGM9
JlPA7UfHNw4KkwXf8yU3PscZ+P1SjoX/rH4HM/zmNDiw7WJVsQXuM2YG0rq+arQgtaXZwJ9I0z+l
PPzGHesWkejTKb2s0b7Eyu4y83i+pL1NYaZb2TVinB/zapCkdXu1J3yArRDIYvWMtbDZc+MDSvFW
FFucdLvhVBfcPhf4hT0DDQpTY/QSV+PSqdXwYfSkScAQywqZHkcM+st+qGxEg3ZxVPDML7zQe8N0
yXDxRdnlCJNIhGLJQWH7Bbu91Oml1dBs0aHUmQ/LDsl0P80+TpG0KZ5OlXsypg17v+BaJjpESw9X
U9zsy2w5OVFuG2Cj4Vdz2gtvc5m0WqqV1a2QEMcZxSypgqBTDkK+v1Ka8Ye1SVwivDRqY08P4C1F
CHjcBa5EfDEtPpF+6V/j+CPGdmmBIIq967NtHhqhRx8vghVPhn0ErK+g3o3qTiiYp6E/iAXyN38l
HaKDFAV8YJfI7BFjEXFEzAHiEUy++HDYXd9HzsIvC5zTHN7770JTfvAIoauiI7mxkivRW2YxIQ8o
WXQ24lWFL+3/accDU1JO1PvGphB4KYIR0gymtgmDvSC9uJvxXkzSC2Erg3RyMmitn3hbbwIZvgQR
/GbJjXUIWFpGM7bNUSiQlpAMbfOAmFiOua6cvOlhHtBfpnFHuygcmKkaOvk4W5NtTdAbQkIyQs30
BOTOzEE0urhbs0OENuHfNecA3ueIfqNbdHCgUNXiZAYB7/UVjOTXQTU1R1/EahP03kLTOCncUPF6
VKoflfAgJtCMyoDprrLpS74v2bquXWHcnswSd1adpfQdC4NnTc+ei8aHlGE4k6NfHLR5MtZ0LdPG
meO4LO5/be/lQuZuzBhyFhh1j54lamfVQa3LjkTR5zE2H7bU+zLDiRB+zxAqGLojKwtdnlmmPPgu
+2nXIPw8Ex4MssbgwznlWeV6zSIyotFp/l7s28ZUjcvBgxbkn42yKgO3xjMuaRPFXK4kt1E4fmI4
X3ydUyzL9POIZo40i2WSGcJmRw877Z8Y17EFmmJFH32qAXnbyu/9eA5EqaAYHKmg0JytqfNfvokJ
xQAPKQc36zL2wcCfOlRnC4gAholNa5sCfRC2LtfnDFY9do0WphtNZT/ygOoJVwqmRnpZQ6VAOcqf
QIraPXCLVmo1O7sohIm+MJ+6uaLy5jiR6PdrS6z3Bm7U9TT1EPwH7ATc011ZFmJH4nMyrD/cFta1
ALmqT62mAhGhwxOb5pPRKrNQ9VqcRmtScysx8V25wuH0nndXUg192ku9UeMfeOTfdihFt7t5oWDZ
dnByMvTO1eR6PEHaOwXhr/XU85Ls1DCGleIBJfuqGbgfDJd4KSHRZpPC3yVR2H6Hs+AZwa2UOiA2
ltj++izsP/splbFkASJCY8KLQMPInTe02tZ2g91FoneR6N5U2bGrOUVKHpN+wxlWx4ygWtJJbyCe
iCBM/bL0p1ptLIcJLMDWGaHbrBXaT84ohCk/AzeJ62tPsfMn/8Gv+ioN++vX23zlK3bGilr8TYbb
75GC2H/mbfkszDSk5jMBJx068xFqEl6NAmUfa0EiOBIqHrB6HPZo3xLaxSr2Ffp+JlYxcqYO3e8v
soQEllqWFkfkFrQjPiierqiyQzqZHX/ojhfXEZZLC7OAGHYZseZv9JsNdaDOCtR8u56Ned0qPlbB
aLv7OWlkWGKH+JH8yrf+lBt+rM4WQqyIaHCkiVHCP5mKbm2azKn0vs82UN51jtVuwDCrgU2cYc1k
TzGigJ924GofZ0qt6vP4MluBkPI/XP3HeebF0lInfsvX7hGamKsWHIyAjfaG7+3LEPEyEb0O3gHK
ZW+2xC/GsojAGkAqDrM6AJc1M7T1PrWtguIKSpTPorB5jXSlPSx1+UznT6Dj9zrm+oB79ErS1xWb
k3PAsj0QVX+Nsi4r00CR+L1SNoMLKAMFCn4RYnnKnPCArmlExBu6R1KyyahPbVGAfaV6SiKGDtLT
vzWx2K9sewd0hV2TwSUxNR2KDkCsiMfSWJaPQbqXPTHs7pN85DccIxDcQXH1kP1t3iRe5CQQrdZP
ng6juhxgb2qCGrXljgEFiP6K3m73kdJDz2rR31YjMWcdEZ5BtMaMU9sSKP0J0V62YjqAS1mEWcTD
0VwZxFGhYhDH50sLd2j4ca4tXHr9+HpOdLGbJCvjP2Bc6xWpjGKH88/uTH4Eezfp4wwmZ/AElumL
4Ko4fzmhnrXlssT1l26x9oGgQqpISE1MrQdMSxDMtZKqJPDvaNkDC+E2otnXOUZ6W1VVmaFczFXi
3OzZc5sR/Lgc4swAkoI/M8fKGriiimHxd6K4WKu9kTtwJbo9cUdbopyGklSlEu1LrT2wEGN9PrKo
SJGPpd+Clc2xDaFZJG+Xwcs0b1AHNLyXjgCI2zhzUbxYZGqnQ/y28wg7T0AqBbSXWXw9U4xXCi+t
bOujTXsRFPOdLc7OCLjZAZfMK0sxB/paruv81ZUmxFrpj83ebKRdGAp0d4CQFRT1vyAerDR5agCK
w5/vuK+3gsrGAI9QqQzeaAAHoPI4f/oZvXPpZYrMDYBSaibWQM3YEggVOdYwFCE2LlkoW4XuBPO3
bX8zniKQPCjCu8VNg0Xcpu7gykTrtHsjSVrYzFimCl4kheusFf/9s+qBbmQqj8Bj17ykyWSWGw0h
AKjHs7G7tdwn4H75gSu0dBQd6K9AnhfIOpP2GJ0/mIjOh8FK460goUoxP1lbeELk+Sci0eKoIIgh
TWykaK6GlFfZVqVfKG5PEsuYzYTmpZzlTU/Sbdq4c9wTY4Wdr2MvuEr0VK1wJpD0mKWEmLrxIzS0
W7S0Yo0dqSBroTLt0Wot4GTSOXca7TLTRg3Kd/HVd0KCZHDJzIkhk9MUn8/vp2xH6LAZSVxoc++X
wGqOlFQ9nbNLIFGoT5FdDwy4sXvDD+6NWyHrHHmIZITyuXvpRtXVRBZMm0nLSeGvs/aVktlZ3ksV
j07XYE+RXONXhqm1XUxTu2OCubgvOs6UCfcq2XWc2CiyU/Mhz1+X0Jpz+1zz2EWU8cZpDmmdm3Wf
FEUoWx+lOpOQaGCM6O8C8Vwwu4+D/cV7byrhBBQG3KUSpMaFEetH4hmlL/LX6+6TQXLgbYjo0krc
egH+dKf31lW2CjOSdkuUi5yWJrFcxLGO37F1MlElrleCio4JZ2L0amjRj0UeDc5yRa7QW3GF85By
CJhWPn9Al+KrIPJhtGcxgObGGkwOQMbvUSDp/PawhCOa/gXAbAQMmOtTb25w82L84KNx6YmzOCN5
uPBu1j/H+4XpjNTEnIFQ0efCBml2X0hIi4RZtn5Jukpy4RdpNVYtZK1UTHRUsJZJW++mZBFYr+WI
w9cx2FUC3PUzA37FOW2FrVw/Bn/TlVmWTXvlel55AKQqhTgAdmCsgMSn89MgdtBe7A5r4pfutiu4
z3FdhNHiBERKTuUGO7t8c+THadmYS1NHceeOefmVQ6+7EpBS+fZmFtksYj5u0BTDoGkcTRjTnI16
V59DkwMeS+OrnY43CMJKvSSCKtPzHdePpdBG4z0ioaiHcbKZ8r+Yb7HHj8XeMmyvpWZXdQ2PIFKo
DHzU6bjR+EJynzsxJ2mqM+afNq2HKkJxP4l6dR3UsXphO0CM4K6+zY9oi32bzE4hV61I3R6q6etX
AJ/8mg5dxRQaV5joBgoDlYZdacyIakjaP0GX64qX7H5ZA5+MwcrMmTShIZh+FhVr6GHjyXqrNCi+
anwY+S3HO5RlRN7U8+pgoAzRFnOFAXN+7zx4QlQMpH3T9GKR22EM5rMEw1IExkggcL5At7I5IYkP
YxqvqfLzjG0cn7OMMG97XTnRI92V416NqQaR7g75LUXfgMzT4h9QvZX/Pxm0PH3+ScJBex27cTUo
0okr7u2r7lCQiN3Fi9geTEwIZ4Ypi/hYgF7yXVUYISB56xU8Tkd9pb9J5zm4Wu4O2rg8lZQGcVsK
y7lmIx+kEZqfFlf03Ks0RFUlvlbeXBcBIMTcI/2BtDMh0gb868lS9qsHubR1toZCWINCXg468upl
9gZvVShEOxoA9QdwyXHdC4BPLutlI3Y9eZ0x46JH+IdvcJ4QwHzL2xo0WV2QvOOUeeJZh8yaEhrt
j6DXzel0vmvDZfRjivY+eOmhRvBG1s5Uw1/PpsagXsPs8tBB1TSEW1bvDnL6M/7pE1B5Sr4oCthu
0h4GTg1FZMCdBcEfAfPSWPt4puzakC6Guishgiuj5nQcgfKf/WSTkzFEMLmC7L1JwjhvLxcq8co+
r9lZvtyY5ndbVbbHxdlyMlwanswvlVju9t6m8Q5umMmLhzlRyL34mRKS80HRr/wmgk3dmEMUKtYP
KWOUph416F9/Wc7RgcwxyVqMsdnJF/3B0Bw9jwgMlQMkkrzLXq+fJV3MSxxNG9Y1XXcvpgPiDc2d
7MHh/sbm+9aK1vgdvyoGjvZJ4bR/Dbd8UPFjqxB4WiRn6dNLeB9fsnayKc7UqTaANqZB8+PR+F7z
oh6nWOTbWeFXkKAQee0tKHY243mnVoa3X29sHOKYiX/k8FBLuV0yva62NRxjcL+gKg3vlbLe+W/4
uELBH/yaKfltsda+wg2t8VfkFaJeJVlUzY3u8tUj/mfBIfroZE33rvljjSWajNpO7iw4Pjeremh9
Ir+7sZyHNWapK04yxSiMsksAx5hXRZkhGueFlTStlamKx+//ZSiPCeicb8aHBxGK7BTMNHGAg/Co
QUAp2IIVUh6zWVJpHW5JthZ9PVhQOLHgMmhE4N7lQY7vnm8TOVGtUGVv1j1dCutJZRWYPyfoj4CW
+WV6s1OaYOK4hPV3tw0AdeAOR9LPW5InTMLC3i5i8lVkKs4QKx38rIQuiYoNT81WlQyDW5b9bpPN
/y6ov8f9zBvSqZTMhxM1DovtIisyVniqgAL4YAcPzhIlIcjZNHolXW5w7IJZ6j6UV0TVwBCXDMLK
OKM640ZeljyacyKsB0XBioTC2mR4Z9bBy3s9TgT7cH/hxSMJR+QXOnPoRKPt2owSvPE3KWwIW3N2
Yw25t0DEOu0k0SNf51RSZm2UbVFGxnYCYQ3nowyFgb7NQa8+p4hxeHg8bjCQJUeNXj2ivQVeYQ3E
CmDzFefA8+e8mh27zIsJpNy7GEClJCnCQW7p+HKCw4wHNLE2AidjeJO89dP96YmYX4zHKAILmLHw
fTAi9vUkB1CBa0ac6MCxEXj6gNwBLH9t7n2dSl0Q5/nYtpOevYJQDtLfn5xelsilu42oF3JfRBxV
FF5Lg3QMOZ2JsbQQH2Dk+/JPv0yBTH19z8MPGZgEP4Pa8wWXqw+c+IA7Pd8VXajSN0SldOTec0Vs
fIEpsHsdRxC2gV/hopgHffwZagdSD32gNaEoZEHuehajql5PXPTcu0dyodiPxm3SyZHqElmipxeG
sRh1URTeqAvKmm5+4KSxsu2klM84N/vsYfhkaE7/RshpZqcZ1kWCLMh7xSOJ5bFx0Q9YqOLRnjtg
Ob0aiM2eUUYaOiASozbfcMbV+crtQZKAUE2nZgjrcC+pZ0jsorZtbfG8rijmnFk6sZEhXlaPNKoM
TlDv1R7yZXZm3IcVVCLk2u3EnB9D0km7qvP+8rn9nn5dVP7WX6SeUwiFveFHyw215ea54FvNjk8A
vk4hSV7xO5RlouaNgd1m4U+MDbm6aT56vn8rcN5SpEnbvD+9Y2qz3KeuOreunEijV45nN/f8VTXU
QC1uL80DvsJXMZG+7WqXKWYoxpHiu1iR58s154Ay3eim1VMy+KqCblVjB94M2grraOErW+xgmsZ8
CekbjgEQ8A3F8N7ynECxKKLv0CJjUDYuU7DHMHn6lpQs5ynoGpVLBQeI8XVG2PktkDA8Zp+8Yr7p
xL5CTU6oA0Mt0p1xbaRkztd5aOYtIwx0f0bo5/4FukAxuwCRwMQlbuMh61OmBn5KlU3AERCm4Zpj
xwYBs4Bd42T95gzMbTFwsDmz82VZ2HyMG8GW/aj44sMcY2PFJiVxxeC2agczwcss52HGWmJmoc6z
ca2Klymb/ORNYQwWqEYOm4sFlULlQVRhROYCU935YUTSI/MQ3alzZydMyuRatOTiU2hfw53vDs07
xig4C8kdolFW819vagHZcmF226nCYVADlcOs5YfVGFdjksZ4TM5qr5vu91bOMJ8Lq2r0f8xbGKfR
KUZgJkryYN/sml5U/kqE5+u2GEAtiKb/BHAYZkgpIiDuXyPmmxSzMRe7dSZX+faAULZEJ95n+Ev6
C3ii2Lyzf1B44/OkIfyKDX6AiSHtUHcg/VFbIghfLK62iOvgLpq9S61hfMfJgw4IkR9FpvrjIYaG
jbkVc4sTr5yJ1zE3EhiLVs9z6+Iu6Q/4jRr+Cm9dQXVl3Wmb8ZgSXKZessy/Q0HbrxxkQvw8CakT
puJZD3XWbaYtAonss/A7FVHOaOSMFm/eQ4wWnKST5Tw4oN4sL5GlgAgEhehEhZ41zdvG37wlXl74
4lxrHZEViMgV6XcOWKDa9RuoQ1CZLXyj2jo+SZa2v52lWC02WjHz1bnHvcCLH42McS21Tf+/Fli0
QCAjsmR+hlXHPQQK8UypcXfOTg66lIh+YOckfVVyz48PzUefvlYvFmop6EBFJSm4XgPpfuZkS+Jv
eNJUQEMDF0zu4WnwGeIAfefKGI+9lMVprBrBXOmtTzR3iYzGZ1pMenFK+JmjUnYwEqaHy85iF4IB
JfNOGCKDS6Of5oqA5NfA69otElFAMcPSkUyaI0kEQeQLCJDEUU5BTHEbvpuy8FtoBTSJSmqCR4GJ
KyruEaxjSUsY5SF6KCiJCt8Fvo5J3O+rEapPYzxjj7ErPx+9CpBP7PMv8aswCLL7LnUOcX9aS54P
vF2kqIdPqIjSwXS/ao4yQLJxduP0YAZHWdkZSDCUCs/3+nqvf/xTMLhuIKuNhg4dReSby40tUyPc
Q2A7NCgm98UBqf9gH5rbYppyiCnptctItIFL8WIieqpYU9GqUxtFNeWm4Jky8kj08Hc1+aXn34S/
oF8qu1EjNbV/1TqeXtVYmAdS+CjUd4mlkRBEZrN2GDCLhdFZqYV7bYRAvrPv+zfR3Tzd+tXSMm1+
AeOvuDe/odB/Sqws/jB0WOEoSdWYhg0jKajo/1UFuehrcRM7dN73llkDGfMImwJobBgzxV8aJrMb
uTGrx5SoSHT71Ih0yBbrc1IVrNrdZnB+T/8CunMBWv+/5QN8u5SveVMJm+mPoqE/rNn/8h+a8zPC
JP+BzL8BqN4ffEr08vryDchoRT9EDIlfIzNenkh/CGxbOG9mMb3B+h0X6JzrZkfeskoRw2XNnk3j
ZkUT1MSKq0rMLxhaszNokD/tV1hS91x7hLWD2u+r8FmFTubVib6A7DBYSKK31vULoezLXsMi8mz/
U5ipSxGyRzIVo5eAU+2vRsNIzjdrK7DHLJAFhm6DbDt1dWJJJnE+fu/ITIAGOBDVo28kNrwyLkGS
DLG2Y7CzN8Q/brno5usmbN1HsPI15ZbmItfyOF0T+UOZE23dk7Tmkph9szmKqm7TsjcxVaZkOf+u
iVdhTmhOf5YdzhsmI4TK7k4o5L2gicBAcpCzDQQpJa/CTmUPt0J+35rxRdK0WlmsM6M7RnBx0k1u
XAIjVwClJna+BU63agfXuSX3OFkzzK8czuzJxfmK92Wyzqf8Wmbkpm1PZOWvYAFDfzNs31K/QtaM
s5Ksl+2f3BOHm8rYYBCiJmiMuQq6n+Sac9Kkmr76Xtj7JyeMsRIvSRxAukI5aXSdchZeVp3X+IVb
0QhfqYwyx9zYiu+EvX1/uuHX5r5KTIpnVs0j5GofFIdMZbs6oaE2bHgbho72GaGPtMREfdW72oRo
ohCejHR+PAQTb4I5qzxKNB6AXj3yx1MaLfJFj6xFXABnSA62x2f3x2uTaTDlKrixtApGbnj4kchG
uaBEiq7ANYBEpJ3Cpxl+EuCVs22zbjtEnLafMjUzTURa8Xl69rAihT+CkB2k3adl+2jPon3+NgHI
HTkEx0B72NhEorSS8YCUNA1lwwm6C6rRyqBdq5B6WbPjtxt6FBnJiaZSSMgIjbd5z0kiMG+EmCNi
klHQZJao3FEuILcNxJMYI1prP4I5kTOyNdOE9A8D0FGbSdNzp6DP2Dtet6VUJLH19QWh+wo54HUM
ZOWaZj0kN3vY5a0YH1ER+r9XrtsRLy8iR03si3G7gmBTLgddM3oJgBQv55hLlKySO/sCVASJj5wo
oUgle5haOZGqdxl8V30j2RZvybbFuXhPTv/kP5QZtgmJ68GNBWpmZ+sWauADGBHypg7oZKnhDanp
FBYVoFjkr01lfdM6qgSEprBWPcuKnBXFWjV5AKGecBTQ2TCTKk/0i9T9ueCrq4N2Mp8t6hw07/oz
QhQ0dYCjx/EVm17Km2Zdaa06wfMJtdlrs6y0cU1oh/IGlDqBh/tttHFXsheW4a1e0u1iZSuRVyZE
+sARUJzUo+OpHquWjBF/RPQV9d1lUzLiN1zBVv3Xeb6OtTa5PsMG8oUAGQhslj5yQfeRCxWryfqi
xIfSl4kic2C68KBBiUkZO13AUT6RobzaCBRZAhjvdeTCMDkNJYUc/5sIEWSiDa45Clk1zQ+25pzJ
TmhXf0SdKmdTFVbWp12x9pyNTz5fggFLd/sxj/K+QK3sErU5hnIR+CGea4SJjY/Fd/o1HiF9MkyW
u6VaGPzU/TYy/xX/T8eUIJPCpXV+0zUDJDBu8qjj3bXKW8Grhr8X1CSuvrp43El2ND0/EBmto8/b
sVBtVfAUOdax7neTMNJs+om2tnU5JY9T52Qds05zwhpOZoSgZVLfNxwnWEiQNtdRCWC8m5A76hT0
miy5Qy03RP4wcER5+UBYMkMH1nKBeMY9+9NmHiH67+WnVZ4FxUQxqLbczRkTSLTREwiUQ+oRT4Ko
o9r/pgsQ1NebZu6dVjFXJ4qrNeVyV4xz7Qa8zdF+/Rm80+tD6kHYOuxSw2mYA/rb2ZlPWAkrUdR+
sMgZp3p8qaqaXiZQQi31Z40/S2E2Hv8OFSY827ixevqz55kN1vTIvlvxFgZ8fLr8NLwBO5pIt0/c
yk3CeSWrkh91qGzZPUz0Bh7iAKp6Qm2Krz9ZSTSSka9c1zZhHoQkmU/I334ouQ2phQy9sBvkY2LC
2x0An38+ZxEVMXA1RGzmM4PzqMpn7FxnVEXXwEnhjfusV3vbRH38ND5pD+NgdnKCZQ4Nmi7XISP1
zWysZ+0oB3fyzMYZTlPhlenbVolL6QryBFRYGsliSWfiZxprQP4YFycrnGOzJocwcaSGC+w1yWPy
dVAndx2TtnVtXXB/i93I+FJa8Wsom/wkhktRuXGy1jIX2jH1w5wCRYKtxv1Td7ztUOPUSttbBgPv
jHqGldlEMMl8RnFCsYLMmhoaB9jzrPTqGYNGz6tpydB+ux2W9QrGRKHxtEgTyT3Lt//VxrqID42B
1M60bHN24saUrt9ENilC04pGDNb7Fvbuq9YOSSOg4sbGNQsB4DRqYDMsM2fRNt/m7uajqAapKcXw
ydzA/qfYymatgKaoc5j98Zg7z6Sx928kh4YjlQTfd7cnAFd4UrcPjS41CYCZu3cMyQhvNrYctytc
pGP6Ot+vyxUO5nEfIeB7W7W2pBZ17vJ/K3vFh2/xUQyFnyV5VGcvYhN26Wd9AfcaOKykwjze1heX
UuqObNgw4T4o3KKTJ6XLCgJbeaSToC85pT7G6JQQVFLPuyNxW1gyZD7Mv/Dwo59FmmnP2PMkhv/K
yuBHyguLBFmf8TMV34xsewQgLbWyLr9l3N5dvufFw8QzVjk1J9uBs0grqtvWujoiwpt4eGbATETN
GDihC/yzCoc1t+YgM0jRaWMWKWC3wJBOMLWGcBHVjPOMLQArigT3W2x9WPdLWOsFks4fM+VVBUHv
k6yjD1htzj8vGFWAjes3XiyACP2442M5DTraOXZCR8ZRHTyfBhmftQCiJwkn8ExgF0/KMFww5hjT
oCsQE6VNyzNXvwm/NXA/yV5mcwa6e5zB9pY6YoLfVg68YIF9/bH/XPS9vykRUCiEvAjefDn5561Z
tsfO99OOF0PBJOS0mx12fQT042jQd2NWhrpknbBO0ZVIJdHGE1hrE2mNLevWZgHIxo3j0wR+jufb
tVuPlgB3aJhZ73XsD1co0AnO9wlOGN+NpsNoK4ciNC9A+yQIOX1l8VvYFW4kbmtQYmQOt0j0mPcG
4d3SqpfU5gjTD8TWWJyFY4dVZFeRUMgeIJdPP6Rn2zhxFxSHVSFYez/JSN2n21veT4US2SxuaSJ5
LqScHUBix1WZoLueYyeKtteMQwDR0PnSQ+X49WK85y/OSoHrAcOHBVKmi4+FJ/3QysyP3wYu60yX
E8qZ3iopPnWFEwlHPqYnCHGTcP4YUX47HQ0SVNPDHBv9cAG+7e9lUHeahFi4FrkrnjFC0F7CejTY
oGY4i01SXdCuyTmzI+fYmZc4urEUwm6zFu3ziodygCflSqAkJ5V/otK49U/NJ6RJiKQXFL8Bx/33
YHCZwW6umzcERsDgG00H01l9ffvIZq9LQoFqTEvhyxjAV45OCas0QnVymSU5N+t3M734Nb+ZeOpm
RMIGsmjhzFLqZ/1IQ1NfUwAnrSracUAChWPFND8vl7Q1jnaJn0AN8zezneaKqExA7JE=
`pragma protect end_protected
