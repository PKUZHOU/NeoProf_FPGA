`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
ZfsOWD362AoU503jxylvXgzDQtaAQ86zFDwfusSudp5uxAtXWAcDCFkxs6ON+kSd
4O49oEAgNWnKqAonksg0iZiycpC9bkRAqb/Q0m4SFWAIKQvZWD6ngf8inheU2fGJ
89eZ44aPNIvwtVvkSRQhHci40fegrlkKIwO9s4oUGAo=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 50288), data_block
yiwi+RLlwoxYnfSyquRKHIN9BaKEWUrfeV/a+8TN5CCQmLY2HQ+PJ7Lz3a1deyZz
23qaJMlf9uJfnJZONvSojfZT6yd9IcDFYjZKK6P+YtRQLd7Q2m1xPWInSxb5XkWB
DhzOiaAvNi4RrG/cjnSosgv1G+eSsRJrMlmdiv8az5xg6lTkeTsLs1t5eg1X+VS/
QIBsb6+eYI0+GdgQ+ooKmEvqKvtq98VCSzjmF2ycx/cN61GHf5y4EEDOTbZdxcH4
0v9CCyqspuUDeL0c8lcYcA7v3qFKW5GhxodI1D1bHu1Mrt6SRdkOB5KhuAb8Yquh
R99H1xz7NQfzXwtcqQ5MeqZBhrnPlqoD2HWtb/wpCvDJ4l2cKpZQWYNfEpPekgO/
J/fZB52cMTPB9NjPOoeVClXTScutL6KxEuB4G5SwZr0RvbsXQxBAE4R9RXPrd2db
40pUVE9Xk+k0IrNhW64o0UqOdQzjjQ0Z+W8LLZKTs6MhYunmCXgyAVhbhGcVOlAP
Jb8+q0KShZ/M/lR5f9CSvoDaMrX2KZCbvCsR2wuAdiwM0SZYSnv4OxKxKNKSnHh4
IMJW8uGj+YJfqh4yPoHWvGmVh/7aoAPGYNzo8k07b1lHZtmawVKeA9s37AGCm1cv
Ef3tWM9JEX3y8aUasl43Bi97AyeDhtB/LUF5QdKQmaucqMIQmbr1cZi0wSZRsXmW
9krAt9o2sqyFcAAEA5GVqIsN4/CHGvwCFmB4N9wODmIPE5pipk+XR0jAuH6dgKqQ
GWewmuZczb6xfLzYtMcKDNabu1Wn+LoMCxrbNfBRunfc4LJgG7ueAhapxFcBNBQV
sbt9aIBOP5Ummq0vFmCNCftoDaWR8OZwQR/+6DHc8y1pL1eBIlRbSKXcBQSKAnVo
OraMKwqGLHFwi5IGjJoMu0wL2GfxivJ/sXiV1gTnv6TNJlL+ahv/i9TpB144BRNw
F/w94BNJivZemI+kjfxYw6ydVBKs5ek6OJRqy2dXx3xfluAG4PGXNPSQHroZu5/u
BYhsYgwZakZYbHXDqpjHgRF0NUJ8CJ4thQM82apmSDRivQdF9ut8eYfiIcC2Cmhe
krvf0wvCOp1LqLiHCQTJ7GrewAURzlFs1X7FCG+uHFvTNNmwF8HmrL6rKy+z1pW6
fRLCv8f/REbR+3bEHusQ+bJjbcawxMvgWBKISKZWB1riiGuTSGmVc2IitAFfQe2O
yOmlCzqZG9dTdgFnrxw/BmkV2ABdEHTKd6BHUst6PTnYKOFFqBglku1r4hgG0g/d
dIoaxLlEItVUbLWzOT3Stf4yfE++9mMmbNcCjRmmXlvOMANEux3rdAy13+WRSjC4
aQUVBjSKYm0iU6XgteH9eIokIYaAoAEqgWDMmfnZ7ikwO91m0ISiXqSba31FCwwR
U/QSdxRBB5GCW+9jSvrPlgADeMWiIIXZCozGEPzPEZzD4DmNtzaHTWQfHRbSppGn
bSW0AjbFC7Ixwauha806ZgDaE7n013aaxKb9Rv5QDgM5TdzbGgPFPNEKZ4/fa1KN
mv4D0f/b3lpu/WnI4FH1/Qbuw+XDonCOe0s6adeivvJXGXu6w6lEto1JLTdjAosP
lxSAeyzXP/URlL05r5cPIvYE2+VI6hb+pMEVI19TkzNny/aawSozqR2sPYIYDlzV
wirt8+N1RKlMwvd2J0lcyi+Agbrl+GQWWgb2Qt2DR/A1XWtqcmtPgioiO4D1hdny
bjJHOVluIB9zZ4U6OZniieNw5jw4Po5M77R/eqiiqPzYiV8+tOCsE38hVaGWL+iu
YB+/1RI5523v0RltgZOaoE2uW5jnRG5OU36i7E28YfQQGYlZwBZRFSfIXLWqPP15
TmAwd1GBKiQsvvvwFKeZbubRO5/7vq1zONImcXZYRrf+E9Wus+EzmJgNZzVZM46Q
L3nxOdZkYXbZhMiK4+WAJXGcFzC1wT/wKsrIqZ/odAHIpr1kBpzsFGIfzU+viO9V
sMIEFWYr2tb5APA+doK3mP5tlsBeTdxHFHbdkSrgYxcBZ7TbLPzFqcl5T0goPZHQ
eW9O8NQC8RjOBZar/K8XT4CL/qX+40qoig7k0mvZmC2fRlbb7elz5ziLOcRAOE7R
UjvRg0QctLU8HxyCkOUfAa668SqB5BqtDgiEqnOQ56ocHRBB+BP3eVZCt7uVWT9z
MsK2CvQBh3g44LMg9Q4XUJjliMspQreslnQPCTx19iCiUlsqg3gU8dIm+Mve7VuW
8qhGP9EcQE3jpD1ta2ndTgssnfoxrudu/Cve9hGUmJk/VDMloEJPvBZzkGgQNoVA
G945V4oCoubazbABqO8keWWb/uJhlLvLtDjMczW+QZV/mIaetxSjkuE3PVzOOa7x
fxyAKqb87DQlakW43BW1CYzcRuLZTHIILkLl5DXVJCLcmEbJ5mVjlRDG7wtE/c+O
kintCVfkbGIL7FXES9Dv134sQWeGQnc/7DeKCK1/siuR0jZ6pQusT13Zo+lvge42
PcNokkfqoT6ME+9iN/NHjVIWTWm+SJZZWVve2a4fm7q573be9hdfjI83WW0XN4aT
4RVWOG+o5SArkpNZY4hcSBwIwq45uv7bFKiYRu7ljM58pbebtlNO4OVwTpyWaui6
KSTMrm6nDVNaZ4YlZpCRWlvQuB/2PRSp2N4WpyAiV5iZT0KV9v2dUpM12cNDUme+
O3DNM0Sfgive+GebW0gi/qclS9eK6iI55TVQ7Z+iosAu7mIiSTGwT2p+B20GmKvY
sfuj70itewJnMj4jotfyrT9Jq8WeA0NXr5X8DZASMzKCX+L4uqVIcSPayszHp5MX
5TaV65YoON5gpkiuIMN4c4dtAhRK+JP2wr/R3rgrDEZTnGRlSCVmqyTVZ+mG2HkN
yzOZYgFL/8GZFZEbU07JVgYqC44DN/mHHOHYEAiwXt/aAsi5yzG1z5XcwzTo4z2L
Xf2OxJIEDeDPgNPjq+tXct8KLQnVhvjAm4SnnIPt4DMDdsFaoWM5xlqxIu8476Xd
sNzi+7RUyZ5ONlvgvev2beKI5YFIPoVUnj9mwj9KCCqyD7aDZBeEEl8w+HGeCdDp
1oURDfQaZVKl/1SAIinV3QMa2HFiqFTFpMjkVrLzFMEZKtwV7HvgcmCFIXDMHDgH
JiyMV6/UH+eVQPWGujErY0HfKK+Jqbj+EH0kEu3Aql1tZ171iUkVAQQGDmI/+HeO
1y+oLngeMKuj/VIQ8Y5JBAL1t+yUqfs04EVDBT5/gEnacqESP9b+xoehotik60zj
lrtI6aeSnDLXEr/5zT1C1aGOTW8CroULkzp4k2ssMVtKYhTQhsxBLUK+fialz+lU
Q2TnazteASg6fjxBakjOvQXM5U4EiB0iQbgx/6k9cDRNriR1t8vqppQUz3R04/KC
tjmsIi15n5K69ouxisyPwcfbu/GVcHmWRMWiwmE3SAmMMnTAydEaZa1PV6hGosdB
gCBnB+dD0yxBv0biRrauWEKOZb0MJbx2GMGSS0q5Nt6xDZgEK+gf+7ZSKgilmNwo
7M0bj//U0BqvMDmzcosYBCWBdM4RmtXkNsBw/nqkBbB9BqTckqkdnA9GRQ3BqVru
nV6K39ZqmWmoGvAPdxKnjORqrIC6F+GdWEu8j04+pYaKjln2vr7FFoQZiIE3EBKh
zvlxHyMwxctLLmmYQcYTrbiewu9VeNVJZjXL8vtGS+px/0Yt+PQZhl+qa9IolImj
gqLW5subFEWXZj/J6hkmdrl4OeXeQv6M2DhYWzy6lJ/8gCesfVQWm0FqJ7cNr06/
7kKK3+kmGpst1v6J40+CigFv0tojBRDa+VeIKTDu3oOKFimyFO2FXr1TksBkArao
qf0vxB6kRFVZbRVOxoiNgs8QEea3r061pxcxy0jc2lR9VcH7ji1PHOB6yAjxakqJ
QWUoqq+/ZCppTjaOPYarpaAAUVeYFzs76TsNfiPfdS61IL4vpsASBYwO2Gu3xY/g
otUib87R5yoAK+0GRv9gqDkfR0U7hq3lBOF+QDcQ3/LL+7Pgik3fLdWpaCXdhVzR
tSZdmXBqVOLYc0xtFd+5UHiM9WAoJVgltb7uHSXseJMGzT9U4/y8sSWscPtQzj3D
31Mwpg7G/SKaTYhNUIW18Jq9/Co8yTlsY4XPQQYXUJPFX1iYyD4L/WFEZPZ5nGle
/LoVNFOY5NSMCYHXor72LN4DgoWLtzdeT+WJfxJqQY1Pt6B4brKbu2qwj8IerA7n
CVTdROrgAlRNS7rYKZPu7kB2xotIhYo2FU2Gw3ttzm5jgf0XRgrYzGPg3DpLZtjm
e58EnubqCSAlsUe4P0hcBn+IbRaM1oOwbuLwJ5GYlivyug+52O1rDVljN8L5AHR1
Q+1gjWx4e23SHJBGUTkEPkK6iwfwm6KKjreBgJFsIXd3n+VIsCrd8bmG2FDnsljp
3fSIZOH/coocRPFosrnnIealXause5U9m3xtTRoxhlcqcZIa22zhYHX1emreoUQH
NvKQPktHJlVzU2Qicbnz4ajTk7EuAVrA9dYIq+GbPX5p95LBxUKIRYBkBA91mVAz
zVAJskvOFQQaDxXYAKpdgCdAkOIMvp2DAsuMTxdA9OK7lSJBwjdtHUxB2EcUAnOK
Lpl+hjQ+8w367rUTUw81LY8dxgeFws4lBrmRbIrdUL5Cy6MjsKsq++q9SDAj7++H
yqkCgYWA4YaFzGp7sic49WY8Lo+od8XyG1j5DJpFfjorkJWLf5/t96eaBxuH35qg
LxBFfXan4x+FbZoCL1Et3MemawNHXy+LL53MqOkHufNOc6I3iUJRFgAlcfxapt29
w3eZl4sAlO49Wj763c6GxpTmhUz6vchMl3JffqD9jG0OcQ73aKrRyUWNduaN9vXL
YxzAFKi2VUF0WtpBZUGXOtYUxpTtXaQrjoLEcbSIwBI+sWhY1vIYT0lhoWR6sA+5
U1Jm3qep8EPyiF4XgOkNTpq647xYmLv4pFn39A2HQMa6tKclTPymAtjCXCgqlbmr
n2kLpypWmRF3i45ShELhaSXYZQ9BHhnpVWIvYpzzmm2t9pYuiehwQkCBf4XgY4NJ
oD7jTIAMpmXMd1l5QAKTKOV4LvKWY9EpnCaidJfXUxdluDX3c9JJoh8f6DUXhEjU
jsz79w9TNk109m4TXp5OY3cPIIf8eDVrlBDE8e6D5dIy2NOJeh1Hquo2/RhMS7hc
tGRLu4M5DeiFNvl7hG8ksyvLLZJ2DhNtfmZOza6+40vHgpq5FuJ3wzMpt36VTdCh
Tn2yLwv0W/dGtpuFtr9lRFOncYZriMw7hp04jTwzzuUTuy7ahwdkczA4tBm0TDKq
0r70drRas7DoYsdMdjHej7MKs9Nko9/9KO8Qwp9fJHjad9tWQFF9QUHGY7+BgdQ+
HiyzT99dBI44wBzBSGsMGF/UNBzFywVWNwe0eGZWWcZyzpiTXv65wAuVxQXXumE6
3pzKEutYY86ceWo0Ox5+yd1h4mYxLFzngjoymPg7DA8cqK8bRZKoYqqvMaJ1ez1m
c3c3oYIWdJFTP5wMJfQp5Mk1Dam3uMADrhG6Qb+Baqr1r4GOEdV/TdzD8mL7Msf7
xJ47efWvxas5tAMyWwKaf0bEzpgNCfnFe85hp4Nrl5ExZCJ+uCarunaFRH4EJjJm
n7XkH3OBPXa5lGQTR3DltZ3+9CvnFX41ar/DYH3GiwogGiPlXtjIVR0+ZaWZ1uya
03HjQjPIL8gyQYAIdtlf3f0EUoc2fKVA8c1EoPiiEQ1+kMqTPl3u9OHe61V+W3sP
NVRG0QZbTMTOwRQHpTcjazCXyeHC5ovW3UahM4vTxr/KZKXPU0WzTQZsTFBWW7Ru
s9uCVmCcz+7MjQZykRv/nCGk1npx1wXsDxgbZcBG84enpyzLy9xFk9Kh06/g+lG0
YCijDLEiO8EFcN8vLztf8Axa+tv7Wn54ov+PBlmcJIdMfXzkCnDSWKwDv1BId4hM
XBH7/CYChi+/OqlJ9zun9vRIUYWG4lDPWSb3gzOneBHeTEAk9fSKaT9OMX4umwFx
FAr7WojLdFhZbecLoCI+qLNWy7Wb8ldKX97df34A6uekh5CjuvhwDkzSPUK+74cP
n5kgMduCSKfAPwTnKb+nxGRaR4ITaxQUJAx43ShfMPt4qf8f3xVzlALpfHslnI9w
2peDfmai63SrsU00t5RtgIWX8sZIOlkuJCRTwJf/7yxjI6uHbVuhfxG/u5HyHbQY
qmYuPzDOiBvdwENP6m66gPBdbxFQ/RYonKPtm5YZLPAeRsCJjkUZhogknLyHytqu
FBM6aeaB/1SEO7YiMkI7QiXE16QszzV/utO6f0U4JTr5FbttNUeSlhraFXFTf60F
Nw1WClYqGavZIkV3GT1jfq4ejcEk8ELEt4z4jJMrpoo3MvvI1JToeZF3eUJ9rrE2
xyNH4bgoIG0XjtZMOblxyOVsCkWihjvrAAPM2jdgMnfwnVWc0gu+0XKfUfMNFXAI
Q9KMgZd+4CpVLkGGMy4Rgq7LUwkknQpE/URdbih2fj8rrmkOLCdeh2gBQzTX3pbi
zPkPND3ZlB+bHbqbneWYal/RSmCBk8BaTa/24ychQCzhlosfqk0Et8lpLxIUb7Wk
UAgsPT0YMEO26pgZH/mIuFnnACkETi4G2XsbA9+i7P8zsdxv5Ml8uUbLCE4HOvHU
+Us4reF8IMF6HvFMctvPh7xxMuEHwPxiXSI8xkdOWMKWR+ZR7LFHsKvuwGwEKorZ
8IQntGK67o96e6WqioxzWn67tmVgpMhGeiqF5HKLTC7MV9IIZUm5AA/heKWBRTZa
lq1mvIOgIfYcZXaTpojoAXYbXQoRKDt1bQ9gZwOLmmwrNhfHJbWyRyZuNbgdWwZN
POPuLAcvfglsorIWZdZbqEfY8iFBjmIDLviPlLPCKQOMs56Lj6odDyQngiscmwr3
A6jy5lC/lZGI84+wdIk9FCz9pmkSf2PlCAVi/w/6UDPVe53frA0mTi7qSvsQljqm
kW3y6vc6Zvr/YExEQohrMlBYoVScFLrJCNvi2Hmv30SJ1Alytxq2kz3cTb4Wy4Df
gPOu5issdFS+BDI8Q2pvGpqFlRLoyyh3YPRTr6wFIHei2DBqL+B0OjD1eDBcUdhm
F/kvp7udS6X1UeSkGusDmM/nt8t4iNEWR23gmfVE9MYj8aKmilu4O9Pl2D9hSQgv
SOoldBBtlVdbzgLx3CLGByhtFXX+UNrP0Q2ZK2FEzlm4DNcPiPbCssJ7JuKINd2a
DajtZib4ffDCTdiCOgnKkgPdSeKPti8fcU2D9Ie0FOV9Phui9Vh7Op3Ha9N3ygEH
UZ+mDYmfYtnqaSYcdVIkVP3lEdrjNf7ZsUst4rTLqxvrVE9tGeF8FM9YyP3rRB89
q9Isk0TzImS56EPxJWzhGdmqf29aBrR64ofGXWT2PZ13kdOtGPSvwLEeDXanThOx
mXCPnzV1uXjMM2+b3ICKD283VE6zaMoHALDF5pq4YzKkXFGQaZhmBIoZ0EY+KUat
3C4q67OU2OVKecViKNxwEeeo5htumWwMYtXLvErZF0V7j/kzQxKxVgXfvbgzfSVh
Rg+TRLw5j9YEEretxpWzXQf/TLCxNEhX3AeNTJjQlJbZ61VGZVmh/T8meFmnOGWa
yzw3agJKzoCiuR43xXr62HUVcKS/G0YExy0NJxCcTWIBIho7+e/QA/t9dz01pW16
hCj5+JwkZGZrbIsuQYtbd8rVIQXotXP8zOcgUhCIpobCDzleQtokFm8vS1gTDQLj
+gDakjVbC8y1BlOEGrWti0rEguqVhTVRepV/jpeonVd+HruKQW7KsvC6asuQgc+I
x6A5rl7rcKuJEo9a1GaNSmvk3QrFsVO+QqN8JqYnZR8nhHR2wgXWFmdMy6bwkm6R
Hx7XZjQNKaroZBIeO2oidpRHnp2DwckmkUd7B+2YImZ7dpofM1uFyjjmhvqWIhoW
tOSVodQwvQXbzWvFCdBN1fn8AITr2jgLZ8HLiBEkb8zxA0sGjWZ11Se6P93MDYTD
GR/u1mFFZHxWIYrb3a8NTJREFuzzHf14PDQ4Zpz4IoNLMQ4MKu86NZ2ynBJ12RLF
iNE06yOBzh6Buoc1PCfyKXg/GtyV1QZdmLuUbiyBzWl9/qY0Aq8/239Tsga8CBVb
ba8jcfTJkRcFbvpjfW6MZ+lyTfjg7nDM+RSlJPB742PN9jl4YYh5OaZ2jg/9PQ+T
9x1oxzK+HvTfIWFAzfddFqBsLdSgJVTPZIQ+HDKApIWcyGOnxbGMUjtNeAia0y/9
h64+ExDu/zgIg5xVpkfYJUGWwVKIPA9v/Cop6zo0PIZwgmtKE2cItMbIU3MVfZoy
p+f65B14fbi+PjKlOdVDLCruMABfOUuZXyRlzFIt4WoRWjmf0QyrHoj4bPcMQIkL
8qboE+WSu4999D3Anl5pZBtcWgOJ2CzzgdIYcvdPMfOZhShMFVK7z6m+u/3PJnZI
UYHGj5CKDcM0NeIOwKARTi6uk/M67XUPfuVvP+2BTGD08YmkhOx5TkpP7h1i8vAt
W1hBO+Lyf0BMxtaJlVpi0EEheDsS20uiECAvtGWV79zwf7dEmLKt3cAtF3V/0Ws/
ToezQgU+Zmrq4ywRQCs+zMxrAEicXBFqSw/CKl/uZHMClY27aq3KFxssHRmAeyCr
SzbVLTtizLaSXNzVWbKE0W0mHtRAPpZy/8oEiBWNsDPVAV4rqBsg6xSN1d0sxsJC
wH3NKpa/4ioP1tfzTYrv7jgnVtrlFz6qZosCxaKMTgfH7Pw3DUu4hjv2rUUIDnKO
uNhl/FtBtZRRKXtw2TfVYE4WDyeNYeepoLTDConxjisArQXp9MQrHwFsY/By7OKt
dSkeYhPDkr8qpqLJciSnW5rQyySbI9z2Wbp4Q1TIIT+ilrOuYxcoKcMm7Lcb7Kh1
RsqgBceOV9tTjrCxjSBRgabdZ9ngTkS1IkjihINeF7AoAs8yYHmsm/0Pxp911iNt
gFn7lWC08+XuyNFI0mweGb84/rYjkDSQw5++PqC/UyKx9TD5Ua4SKEkHuy96hkiC
ehpKGDY8YZ1GvIOB+DxhOdgtUBeUoO6Unveuax0/FTzz8DAEh2mOOQnQTl+CDP10
Sw2GsagYI+nJI0SueiIMWVQdmnUclYpC/l6bAGCSCUExBU/Dd39IoYkczTedSxbM
iDFKgNeEkel5dKeR818sJIy5JoOuvBMFCRfJWxSv7JJcpyAqPhwaj7Uf8aM8IePo
exx/65O15n4JZ7qFeI1Z4Otz/EqiHR0Ldv2FeGCdmcDnGWOP1xGTQ3Wdx0sxojHL
uWwUCLil0sKFfbCz++pHE9+yLpDUJS9XWzlEYQIfrUzLRoDSl703+JMK3AaPvVmH
l9J5g1xsqscHgHOwdqrJFq/rP5Hpsk+VypkjCP0862C0aR8YdvNKZgvythQmVamf
64K8x7obrO5tGMkAQK/jeQEdAToldddm/3og/8UODWuYbvbBYUyViAYWPkrJS0X0
G0TBB/obSLW0L6ah9w7iziJttX+w4nlsYAYcwQRVoYJpV7rKfDA0RF+7rfEeF0Hm
OeHQEIenIIR4opt83jV644DmmmI3DrB6DLg9A5Gco23UJsRXfsWW2rWXUw/L4X69
S9PwAPuSZs5AG3FjGbn0ofOP4jJx8E/RgUeONSB0tVKP83QyokG0ArNf91/8hlAB
04LqIc27NemN4Edbh1TeGEG/G0/r0pJrXnqgcOtWk5D7/8s2+MPysy1oCKiF5hIT
XucDE4jKeJD59+QLul3edLYD3+pdwSmy7r7W2RG9hFrxLNKJeEzUv5PJE4lxcMug
rm47H2YKvF4stEUimLjbqK7sk6wfekXHfh78mPXGJA0F1TZ/kNn4snrVx00USDa+
zHaga+S1W2EG6P5nnPjjwjeGhvRWO9xmRPvM0yPqwGSWVF3tNVSbHtHAKUgjhJVu
6SFPVvPcPdWbmqmvg0KNjUojZcFjs/i+WUoZSf7Psk78Ena+ptEWmLp9GauhakLI
Ga6MQJySAzR4WZTGiwMKhyVRPzas/o42VvTKx2cQ/UM1Z84Dmm6JkAipuc3LiHM4
j3dN/vQouuwgqvo8xGZRJRzJWlerks0DsxMelqMrcRVguxQK2n+yuqnoxRcBF9lt
9ANDJ0tDKz/aDZk73qvSD7AJgUZFjJ+Cd4LKscOrzngI+SkhlqUMv4K6JzHtNj3t
/noiSkdh/66mXpggvaPKrQWK5Mfk7f1kKQKYOzXpeu3YvuWq0Qaz8fjvWmjFnQO6
R6bIfIe3HzuWiRLNgAIpYAVid/Yef65J9aPFZIxfhg6rLEZML2IQmZmVKA5NF8HZ
ZA9R2AOukqsP3P+C6GeR5vJeVuva1TBW9I4C9FZUNv+LfhAhG3/Li+f28QxUvM3v
h4YmfXGnbcXnZErqms5GT+xrOf+mUUm1rFeeyLpbxdHP1xPdds5Nq9VU1H4lWRK/
EdeOK/gmfKngHoCCXSIsHVjGIH8HjzTYd99pyx/is+wS295R+anibcSPOYEWvHRm
BDxGo+3zztnAx7PMC4XcCDjV2iyIXZGA748iiQk+fncWrLC4QA7EnlZ+zp/6knvc
sS46PgjZ3FM2ewy3qcmU9X/vIHWIJJtTl8w8QRU7oYg8p/C4DvhT7P0tNEEKLqDw
rkhAoTmT26Otg4R0n0KyMXbXTq6s+1UCagXyhqYCj+Wk4c6F8wmAUekKVRP0EdXf
jzxDlhdGrReQ583WbGlsImaJ82uWyYmzNDVi9mmuUv05L5pUNohbgkoQmgr3ex1p
oicyHyHTYn6UsvwjQzohmRySLyrEe/Ic371ofYYHU1zNmxO35l6LWYegtBnkzciL
KSV6kARRqc/LgFHMWuXjnCmOFj07ig8ZXdcQhpWAX2JsklxbyoOk2dFNTtli76EA
hMpjHKCM2GU20X6b4Ajjyul/EuUydPuEAOgmzUaax46jk02cUWJT6U+0sixGA+pd
19hASmaNNlmTns/ZCuzd3QqIlwycxWkkmx51KptAZ4CYYzrgQDgr1dOjo1gbamow
1Ti+oEOUCbkhRcm3FC2clQDdUSJnyIpjiwsoToQGNcKPojtH5vwa5SbRfo+URT6+
HHscZqSU/+cwext2bsIVDnSzxxvtv5tIelTQvyI0x4QPOSD9S7/BhLJHfqfyu35a
NNFQyqljCCSjLtM1h1mUA09RrsvBSLg7R1rjR8VJv/9bLiT1WvJMVU7fGmhFZ6or
M+pAOTZTKgam5bt0pakF9NjQT15SONnxseu1qVBdCWdmt0DnP7LzoyZoBEP8p7A+
Xqe44g0+NuaHqD89MFulDq796VrXBMArBs2F1F2+mdFP2TPdpOZ008HBzBh8LBgH
huDrwG/446Df4YGFKLczULLjiP+O+KyCuTzsHIvQeIarnUbUi/1+SmlLt560ksSP
Itd2gToeboaFTbJZcq+GhHNBq27b8ZBYmHo6HPt19ODCFZ+WkdJoXi8ReXv71hts
B+hvSLXTcwe1VuDXaw4FXCJvFfOsPGIaT/ZwBBOhE/ysmri7KZIs+JWgVCjemPRq
bno//JXQw8hcQ9gWkfmF4Qe+6xYyS9+v4xJEZPdzDIwnqF44WzxuA4gNolyvtqm0
zoiRvPYEfgT6fXvqpiJEYA5fICy3PnKIM4RvxO0O9JMlD6bXy2mzGPtsv35muNIs
V7MBWy0XYGeGJPSrj+PPqNFenJnxvZeCFWn12lnGk2+ImckOJXfZsAnSXRzjO+SF
xrTvLcFGJvGJxpvJ7wCIyvEq7sblaDvbkh7Aw0fAk1Rd/dxfg5V7089d1Ljt6qI4
VL7FTzIUPr+uXuTrAl6zpTPgwe4tzf02NbCRqok41wLL/mbMsuA/8pi7g8ygUhSU
pQi/ZTdv4tRF3Uf3TVNyc1KxoySAmuwTGKLgZ8g/zz1P4fMjhcfQFKxS+yL0mgM5
jXxfljn9jKCfdigrvnnNMBqtqUJVpnWfvdEJZTv5vqo6CFGCV5vPcydpHD3AiiEz
D/PvzW1uZi4nw4G5vp/F0FTSWgrNtM/WYdRBQAF0j0wTz37xQpQu6MHfwN3EEywW
y5Vy2MX239qWYTg4XnHfmDrMVgRjsW51g2cIsk8xZ3r7n/Nk2+KmEGFbXzKamtEE
caUY6GooOAoWT+XgAEClpfB15w7oMOXQK29CH9rWHtxzn3ByE0cdr3qILiEWm0Eh
dpqt04JYHcpwxsmKYGFfZHGb271ftCLSpoEEzRiTcXrwDcWE4elFZ7xkJe9r1yOF
U/ZfS+TkvVyOfGYvavv60bDJBY/sG+pZjnnYPka5jp2to9JEihFDyi8UXQu6651L
WbwgJ8PtDmqfgyGowEKKIik1CLUerJfDlXCvfaKskB3400qw+HFYnfoxCp7tJPix
cNICOXFpVNERWX5EOPvxVNFgmlF7Sx4ePDGU5IrC4JyxiYcmrM0etWBzD+H+VLPf
vuUIT2GANMxhqVeON4PEOvlgmVQ7P6ebp8g6TzgRqczh48jP3D1vZY0Ydh6n4kJG
tXdGn9tuXjcfAidos066HrVMs5KYrL493kKb6Y+Vl6yyUBLMOIQTjwGfvvOP5DkZ
HwoZEYjtngmTd7HJJjQZiOoSqdL+GpGNP9tqoVTLhccmNFqOS5P0Cpvug/zFgVkn
4j2Yi72JLAGtNri9EEapmmI2sXS0TYTGUVxJ+TgrgFzEWrj+2IlbPYdfKBonVOzA
j98vsEmPH5tJkyWrfRutGpj5zGZCOzowA2/26ZFeZYCt7DBCdUewzxj/1TSfyV9V
dj7NgnhhkwjHdBSrdp6Jm0Aj7US/TVHEpGyCK2uUGG2lqKjCQmdWdU2oQXLsrGg6
pq6UNY8JoDvgy+FWofqDMnkbvtK3pe4zT1nm2qtku+taJ744ACCb++u2SReiRGpC
ohvpi4zA/8WUpUj4hsc7FBitkTMfG7RjOETm/AgVMhbYiCrz7nx/uM/oWn0R0xVp
0MmMYH+r+shwAOT5tqCn3NW4M0Ck6BnU/Ic7Dd1sHsR6Ot2RMq46VCJdEQvU5CXT
F4NKO/Tq8psE0pXaj9/ADX5BLJshssdmwKT4nX3wV/t1iyEcu47ADJ0CzUvbg1cA
iIQb+6BititrcVZvmRZVg9VXMgYC58mLlQp2ntMGF2OaXsURsp50FxJqe4YiOSGo
nmvIEnjrlNBn5f737q3x9g+eGLbz2XsXTE9eAV0cnd9nrfZHwcQjyz4CqfxgVjNa
pIxQWVLGXa0sjHDvAAehiUSbBWBWBso1gSZ6Mjj1xThEh/gr5iTDOTyt1u042MO9
utvpoDwhXwaKnp8niJ57oiTlBajkch35Tyy3LcHzG1AjQVMr2/WAprscqDCU1jUy
sXdykdOafWAnODpEqVmZAkWYsLAMBtoGXKa5fm91Z1UEpYMkh6l7JKyvKZ5YDMqy
NrSdFS4fhHv8jsTHvGFmqtilZOFi0KN9cF7AWgsza0JtXHu6PVVt8cdfkRFZodfQ
HcKiNmUvP1cifzaVjeRHOJgHkh6UtnxnMdUZHADFgMupgkFXvuyjsWDSoLOh3wSU
XTngeg9G0ZxUcYqPZ3O5Hdxo4yEgci6E9EFMf0DQ9gFOOqB/Nf1C15Yd0Enmm3TM
p6VJvqwO72aFfb01f8CObIgsUFeq6sBf4S6v2vm/RS3SwwWIpy8t9k96qDhaTk10
s4dNT5GxGhCHFWZ2zk75XqDNMoBqJo5f6Yn5o6S2kcnU2EjGeO6YPccugUF9E6cr
dU5xa+bbbXqEgZWv1pFaT3Kti9yuEbObi1zjCGHMv1xb3gnlYKZLx3B/oRHlEKtI
IqsZQ+FL2uRcuwmfWsWMSbpDIc0lBROxZdESJLby2KdTArbd5R39aJjlLUkiStAs
iitRhpp3nfoQjhQqTM1E9P4XGhLs3N3WSJhYL5wMtD+vjqWfQ1CUie3lJrunHrf6
OWNrRMJpKrpWplz8qEImW5Ykk7XpzkwN6FQ2LOp+CgRu8dQZkZ9mBzEVhf3BmuQc
kZw5bC7I53dbzH9x8+OKEkInaR43n0zFuKgqQtOhn6jxMivS7bAMw7Y+HN+4HRcn
02fVtgBuKio6rVqDkUPsI8/2bOA8sV/HkwEp/AgQjLbb9D/PMP2TADuTSp4Sbr6B
tlgYfNVsSxn7XIwJW1zXDK9vgjvLX+YNjF237iWwVswHRYnorHMQGaRtMkDLR9wp
HQYe93pAJgIL/xLNyKVudvp0Yvl+WIKbLTP1keaYO9zPT7hcmwSy/Nav6QBTgZIc
4o+PWShbUVN/jxFpDQsM/j5QwzTPUh3M+RKnkK+WoSyUXJa+GaUhSuIKDDwGGhHi
0z1mdYG0pj5C4fFWuehZjuCdsFxPiSUG6QNFph/VnWHaAMCKneq5xD3TS5dsIEEh
210oOosKRP7p+rZfK4zLxxXUNeqTBbAXtKxPNh55wVDZ8UnIcyODlWhTWVtMx+H2
WDFbfx7fMJ2RJY2qQcH5MazYEZdrjvDJZN4PU3xx3FK5QGLHOnuQFgxyZEGN9KSQ
mVz/1RfEVbnSJZhIzMAO7w1AeT0mbl5xxQsUaO/Gjmv85X8GT6QrvXPDqBgeXKj+
DOgjtkOJyDHzJZZgLm58yP+799JWG3f+GGpR4JOMwhw5mw+bRpe5+jeLm79w3psG
ROFQE9qb+EjnuU+SpLNr++vpTKIu70tJSSpHEn/vQl9M6yIbvnjvPvp394xOMSkZ
MBo5AOfC9XGGoxW2o0mHvKkBn4/VGi1mMOsoypuoeqh3J/R0vvFzPCPrrxGMVlNi
IC6fpTNO74DylHrCKa03s1ExmCcOnARR3qWN/qx5S42rfRazmR3hTuKV002pSVes
NfQn35ELkr2LQMxXqjepSrTGOVhhu/UciYTNFxUxzGwEofe8K6HpdkhD9ODkny+A
6xelgAqIMdKAQF0n8b3BP8whHsXuBTPgYF2t6+GozCK5trh1hbOn5g/cYVwMXeKJ
9RK4BL3e9DXCDMPwMBHlA4SkymQpvZ7MPb1U0GrYlLKwVQ+YmwBx3Eyy7U8OLLg3
Jt4UQF8Ks8S6mguvaHm/feHAlnVGtAGHz9YLPCuXiW2/5uKJc+6cznrpO/rjTayA
y+QuFfsShxvyWxkKxyy9BN1AwgJgTEWifDfRGta02gYpeMHiPI3/wQoF8JjZxGFj
suKzGA/GK1HBRHZ3UtV4EZDbFCCtTOFBSvNRYTDm1vpN6vuPK6nvVjwXDz69Iuvi
rpgpODBxGkwKHfOHIYE1hEgJujMO6meWsKXl/cqgUdwYVnJn+0NFXcpzy7btDkk5
OprGWFImX4bokSzFyZmcQLMp8flCxFxLBRqqm9ynoodyIYbQfq7ATuJ9tTpZD4mL
2ZJ52QYNwEGvT9/M26tIrf/WhSBBAon4lLvBu2k0aSgXbUokT1r5sOUGZeqh3Tsz
L3bXKAnC9kGTVOfqGmq4eVqJcfwcrnKMyPwmIsT38CUSgRmA/yGhfibeChBKpkQi
haaE8ZIyg2QaidZo2NKXXuxGuvU9rXJe6bPYHZ8LnreP3KvMsgF5c78hZBaD1bpo
DzKtrt1z0ejap14RHf2aKEBlwq4ga48u2Fzw6P0TacCJXBlS0eXdYINF9hkVT626
lOj8BzRHcmo8jc+90EHKxvj+MPpmr1piWJg0KpXxSGTeeH7ZAoVBWQdcFuAb+Wn8
DqXsrZioyHOgTYCVizYCIp9bFEz1TJQKL9KisDqWTKxIwEns1Y3NPuBO1NMgbiOW
0tdACJ5sLCxviYZ52JRveGauIjLguV26Sxp5R/sDRVwKAFUSmQSwgXdII1pgmE8i
m2cqvu7RJT3ZTIMIhL4FvD3ndWab/jdPWoT8uEF+TLWFuzL5cfO/RzAN9emAczie
peACSm0Gl9CIG3xrJNYWHcs/NLcG4J9t3ofXW7TbPDZ9Bx7QR4a1e1aDUm1yUIrq
AzPb/wbWD8oK0dlrZu56cu6LPCjt9YG7YavH8JTZTv7UsfdZjBz8R7Mb2j0o3wgB
fVsVAhhAjMghkjuXl1joGHcNh+lZ3/jB7jCK7gNbtRDrWxCkWrE9wxF6ilueYmZB
OqDEWqG5fJ3MOxBSOG3YoNDEgJItuXASeQ6mcrqVWb+QzGAORYOO8avyYXvUg/vD
nDVed9wOqORC72+veBvTAH5uMiAvknJFaV04fgPdqgCjEbcdKQjH25ug+A+SbtKI
yAgagm0cFjMTzO2OVnhkhEmPodKhMRMBXNW9WUikJFtsH1tT9hDgV6QNlOE85qiV
XXkpg6otucl7oJ9zQ82J5dflBWDPLPnNOXUonzresGbSWpqpFz/0aJ15VVP1n6Wg
tReINih58DtyD19Sodrd4//UPlV5zfP6LVUIlrQnqHlec4YuT+DJxO4lgV/ynD0n
fjkV/yGe/69a6lFFMRQ9UXPignKAfaeoVN1XnzTm6zylcgJB+YVrdEBrp8sqs9p+
x1f4NEHZvUjbZhpkuAkuetC2Z1t0Lvay532QUC0PBQymWludkLqJ/9dON0vyc2JI
W9Jiq5+1ZqyRbWaDDBnb6vJXdrrt+dg7nIIbs26sS3NPQ8+xev+XhqAipQo98SSG
XwO4bWxR8WuPc51bYZUjIEG+1qaDbru6z7rRSYANpMeQ0FzgkK8WbvTZwVEVhRvK
sdXyZ4ZGijOAmrxQVZqktuJEGlZ5QCGRh33zkwfwa+VdLDbtzAQSPzuGcdcg3W3R
hPsY3NH+F7ac21G/ANThzFjdtFVy1+4SCn5hhsU038XVW8jGXDAtwGQnMRYKk2Ka
jTf6C4MU+UfF4YSQyEMj7PXvU9TOq8gQfTBR4Rm2/8+OvSATBQC1+W2YcQ3mcKIR
VQZfhNjPFIKAXJASiNjSKw0fhcgs9ajB971FPCuZlUJZsSfM394n719fe9wM8Cvl
lTPCIpLE/Fr19W/xGRIUsANw5eFHuxaOyAGGV8G9gNZdY9l/Grr3jNXjoHKK1qhI
31LeejD8rH54wKY4TAAnacGRxwKv880loaxiPn5MuG8hnJF/vX9DP0xTsyfWoQVe
RQR/g0nHuQ/vlqPE1s+XVhWRINACc4cCSHedJmDkymUDN5zkl+HQTOfxX0q+wzWq
50SVsDKYInWAOd8hGE2f3MhSZrkoJHWy2ZO+2f6222FSXG1sGhVXsEkO8JZfixSm
pmgXOE9pfPKoOtxQfVvrrCI/XifiLYRbhDRGSbrV0a1upB5TpFgUviIhizTBQsB6
GPDz6oHpmjJzXu2GcFPR7PDTRaaPI7Gxwq/DJyBjquAxTIuPje71b8SPqCa9sA6s
BWlOVdLszHXBEAr22hZ/7QMPUY1AZ+qgj9AyVrbGsuWBJTAWIyMjflsy6uE6Qfna
O1Rlr7O5Spq4Pu7YVudkdYqHQ+0ApIPtRUHUmGt4Ozx7i+NlT8DMtLq2BPX5fhbC
2SP3+qAGIu3qiRHoAvX84RsJJ4o8wDYJA4CW864aKILJiETjFEWGq61+NW80vN1p
0a4J25kG+HdliiuSgZ0/cuTBXFMgRkFq70JGspk5/6Dng+yPqGMfOnrvPNeh5vDX
dWxopxbDx+4GEeTE5ZXdI3baVxBhR3paFZ5qtg0pfYHtPfluDS4a/hzAce4eTvlu
edF0r1EAQQ2bFP5NLcBLKlW2mqcW61FnhX1tsm7Wmqg3sYzDahF2hQII8fzuAlgb
Dr5pQ3Yc/W+lxSevTIUqapfi3qDMG2LA1pzDFU39ohwBoMFASiWCKx1V6Ez/ebfV
B2zpkA8a6/ce2y3sNL2yDVizhwwduesFnKNOoO1u2mh9Z0ZoaLRxCtHhT3Xvr834
7t0hX3WjOeOckvvyuFBXZFV90Bs/lgNpSP1UFsz+3ULzsIaLRXRhp1kw/hukCK38
JON8JbWdT4r8ZZGYnTCOyqUYDwVSR/wwNqxb5/9vPuA+H1/b8KY+VU77yzd4/uCA
dfhzcx33tJ/F1LS0RZPM3vpSWJ7KqJYXNqMJ8+itjM3nYPeiAjr0VBa66BLt5XSI
Rxq+G0vjCI8/iINIulnKvqVSOgIduLmsBlcaVF0KCnxXvWNEtt4WtjC3OVMXLaig
Ifuz30Gxu2sVrnoFTrrEJfQLst1VODD1GGuksQhTLjio0aQ2yQUOnC+jmN8DUL9K
SJ+7/qT8SVPhjsMf6lSQLLXU/RaE6kss7a/uaNH9SiSSd7He0qCCMh4IkY9kJ6Vx
ZAkkOk7OJMmbJnvCoVkedvXEdOhiHDSBbKlDMfYVOvt5T7HF6Y7B3qu4zHVdL1bs
7afPL7Pm/+TMaCzAIkq9wXaP0lsxpjzToe0Iv3SuwVt+wJpFxkUsdz8Y2CdtpKdo
Zi8l9kL2RHIT39sUdJrOHGX6CZXwdsBAIVeAmBpnFn+vG5avI71Pyoheb8mAUpRe
RcW/ENA1wZ++nqL4XCEm+ETob7iW0n4M42xNO+LDaq5EQopjvzeQkGqAGAntHYfu
+01oDsnb1/AFicdikhY+viLmUKfUzqOCGqZJtfeiFbzAqIZxgI5gQhkEEUmUlN0b
XWY3uqvLhc2x/JUCEUwiaTCN2sj67WUHZ1Ypjvk4I5G5idfWmWTZbInzLKBUrgAX
qvDI4HIuYo3A7IDkB9C8GMWwQOAPB9TUnNourSracDnLrrLnYN0KhubTG9d85pOc
QTPyOEAKA6H6t/rqX9nujoXly9Au3mAXIa9ziSDlxWh7nY7OPhfyoncG9xv+PudY
yyLaG4X2oeTbgogPeD0TklSdBWhmj+3m38oCgidGoBwuS1pH3RpSPgbXNgKzYpQF
q4m+tFiltygBlOFH0aJUbJihRqJO13bZP7H++7T9a5vPIJLkI1Xw+4GguXGTabEr
jHTEPjXPPIHM9YWrgOjiusI4BYpReUc9omR4z1SM3jgIPfmQrZgfOt7jNqr3pZRR
LHomq2UqOcmWtiQLFTWF/iBKZcI3TJx7k8pvxmXcAKiHPB6/1TAujtrcpw66oPq9
8pztDW/Bv6wCIEPIBj5IKyYW5FHYbjfUz3fp4YMyfziyFqT6pSqKVQcyBvZ9crfC
IXFI9v00xw9KY4GGyDohdvSIryFxV+Fb79vz35DD6nCvUg/MY4+9Gnvj921aexL4
82SL++xLseaXnT8w1dodKOkftI1wQFODC6GZZDmNp+MRnDV3j0G0e+UL+RdUjLsS
KgEGxS67L7jQodGY50qnEz058GxvPeSdchlWos29omYosYmG+Fmvw1baWQDJGa/q
MpulZnHMRnWrOCfGJ71a+PwRWKyWamNDJfpwB/UZXttRElLgRbuVdltKGSXl3zO0
Ug2+ALZcEU0jQO4OuenlEHCXCZRPzmTmM1JwsSi9y28Rem/RA+JVdf9Hr5C78JGY
oRdo8CDjUcSoGdRptCpFZg5DnHOAjXT5G7uMG7gvQDO8+oLSrP3QhSffKQAX4I6d
H0H/fak+93b5e+bWJaRfjB7VLhaMtuUqEnjjih/VQjYqrfKeNOzGgjJ130xK3dLX
m51TtbR9NNF/khF3Vnl0BJukTQjDTSyhekUIOjDRgF3e1pBurzpaJbVjyEOJcOw3
KwW4I/OVPtZlWdtsWOJRi0yOHXZsFg0c0+/yXeccnkBq1WrDtXF0vF+qHfwDyzyY
X4gR0ymEMGYYhURpLInEk0YGTk3KvWalkHrB5Njv2saL5T+ae4QRujDHtw0Hoe9p
APZPlVGbBNjrY87dGOmEQA/KtzDO99a/wGtwju4twNaLbcvL9v6lNIB/RNuUFKlx
LyJcduT/2xoI8fUIvPVCpWX28iI+jei8m8qDfkUvpAmH/6UFlQ5YzbeWpNqkhD9K
EPDEU8zQosl77cBt6peJB9DHmumD23nP+pjNogEQVvQIpFXVCF6Cu7bodpSE1H0x
TYfI+rpq7vRbPQlCQPM0mJgRMRYeamZXKzxOQlZXqqdkEJ2I9DbjP2LXmKvzDDeE
+vMhOSEFPmO6lIzmyFxDzkebFlWqLawMD3naiHQOKrn5oTzEV16SkF+96RePwK6Y
gNZdEeKlwrdk45yp42qAnZjWbh7wmxpOLjBG3SroSE0f0B3OsXtgdRiZnDiX5Xrl
S9oO0Uo1ZU+IXoeQQOaIK9p6BCJuo2wvyXMCDYh876Cutflm4viGRtlesvLnRBhJ
JF6kQ4mPgPnXjMTVpk2cdS1DMKdnnYQcNkdIpFHE8hJnGs/knBtd0trVfozvXx7I
PbiULZDm186yJJebcFn02LYHt6HHES2RbMpjr06wCDvTqrNU/ioI79V7z3V6bIHT
x2QnLEjpIfKrLyNgg2EoZ+LkF2m6kDhFGdfVQpcgtTkLHHdIALkeY5l4eSnrYqS5
VdaFU6sunSQe8tc1BPHiBRToEupmLwBUT5nba31zLy4zxgu/ag5P/y9giEQ/SgVy
wIncl4wjPp4TnyJ4qeCrkM6KuNA9L2BNL49OrCPYybbxrPxSvdGCeHl9OlO6C3Ob
qrAL6OJNaaEgt6xWJOegVsoFIF/O2C5sfgpIteDp20u43ITHdO0kcrXCWwbUmAPE
0/+t/8CnEaEchA6x0ZH6ML0GYlxY4szaFYQIbIaa2KPEg2H4Gl0J5bvJRFrggzty
7HeWCYqAnblxQXyGTtiy6a40Kq4e+MpfA1QbyNKd15KymTzgG5EQMcL/HMA7+GUj
z9GtkzWvsO1YtAOcZW2UCbcokQe9a3rD4Mf2dGf+XG3JNP3Ndft5SxTetfvJ81iM
UQ2S9OERekCmB90pEZEVo9aet1Yy0YR3x1wsYVfyVd6WQWUriAmOXcKoQ+GAJHEW
aBtfulFuZ086AWY5b+yQnc9w3cLWt+LwEuWLVejYS4Wa6IqB0TfSTrRI2OEe8l/6
7UlbJEcMAMxoUV+8eKGWn//mBlSbxSyFl8GqTrcIIOY1TsIUwwFweJZRwb+objKc
j83vTksVkHcM8WFpmew5N5s7f3TBU6NzrlelgBonpvdv4mYHAYywRvybmu4GYFd+
iIR5MHJaovgDWPkH8AoNAFPxf8DydafkGVgZxtlIf5AqPPnqAJcPI12y6Ph8sb+R
nBIiREorUzycCBliHJDUnCnKeqqPB3sD5YxJ4BUSQ7tN8Sk/6Us13AwWBPdEqrTy
GSryRz5YNZBAvtqOVua9D3zw0c+QG6UqCUxT5fneMmuO5vEoBPDWf9GAMqkTmHFe
ygeC23vPpJdgRxFyNKb2TSENmYpzN4yw2FYvZIiqtR0G9Pn0mOyx5Eaypf045NBc
6KeMKwLhB6IvjATEPWM8mcrDUyZ+Hu64GkOUOdhAhazUk2kcoF42D7Cp9TDT7ZDW
NGHHE/kTsH3uGEeh2QqouLnU8RMrLQwR2nbLaEqHZO7t6r+fCXdYOcIXAOZYb56b
0dpGMSVxlFR2L+QsNJ1Lz0TKXNPbmUiM1S5Bx42hk08sc1OgyoClzlbmkgvXwhmn
NjZgHQtUf1o1nGjVcBnvQEvIhDlu5/U+DVQMpZZOLGBzka3fn9cxTOuE9tjMBJB7
mwsIN/dTr3wZkKmXi2HgRMcB3HZ0FdA/VkZDByC8/ji2XkWmnUzsk6K9J5yoJV0+
LWwHDlpSjGXeh3W4STSElBr4XTxEHfT0LYtlwQPBp9v1ywOKPanSoVdQrGqIqvj4
5FTgWvCiEn++tAUI+qqjR6nawOJ70wz6mYwgz/CJvTJ+nz5AXWtdDDpfP0ugYkCZ
Hi77XAn+I5kuQ/Ci+miJYx5JfDNguNcTwxPVnTKQZY3PG4zKLM1O7Gdulo917xcp
2maNRC3tA2F7Wj9nAepYq6919WAbczbt9QmlqexY8FHFWMDMtlvDyvu00mXXyKOT
7rvrDmh2VHIFp2FiUIIWUOdgAECzjkbeoX7UL4TG/kUErOuEQ3CjJRew2vDdu9e9
VOg6gMtUmnpo3DcFcEPIvIAMxZ4dfxQRVN29VIKNvPukiuv7sH7HeZwxtTdGrlNj
R8FfPf4EFBY9urSPMbCSpm9nnFJ9Y3DROUmCDoQoTyuE+r4cVB2VGKvbW0MJB7Yt
Zr6Q/GWsKg/QEs1wJwu442V3OjLF/xG1bbnwLOEoWRSdYAArk8fThp/iTbf2dpJX
kher+q0iS9H7xvd0ZvUCAv+cYLxnzUMzGIFZViFhEOzhne1CjXfVVTHH8D9Q4xIK
tmqAqmG7k4zM5Wdb/HD7iTg773CIFf0wfbVWT6XGOjngpLLClcg+ctqSvU1lOL6T
qsBK264iyhgKIRePyGt+zImJrx3ecQqrfAX7dkn0LUwwRBeUJ+9GuvebPRqPhHEe
k4BdEMhxS8VJrWl2vmkVm/R4wGeWySTlAvxpounJZN2AsG4+Iw1w1Cmop7Bme+Bv
kE4KDreZlFo0kVrXPRP2DyGIVUHzzuM9hWb7Yfl1r+pwvi4C8cMNTCNOObYvmjBz
SlxurZgSLqMymRAamrfDC3wrYN4JHgO7GGa3+wTHmbnq8MkY/4CGQsKesoLj69hp
Felerv+Maikqlob/3Z+6SO3dw86UaB6/aRwtvGBOE3kgH6xin4tEe3AXjsmoWKQd
oM99avLh5zCLmKT3BmbrIuEi8VF8IT1ptE+wr9duRvRt0ZM0i/bEzg1WbIVp4m5v
1y6K3W48Q07Lrgedq9xTthKywgLAc6iC7aB/ehMI4WdLvhIuL2/fWUELJryUy73o
wvK7LES/pM1cxqiFcquYK+t+uy98era4JP2a5dxE3IgL+qArPpp/XoopBrazPsZv
iNMSklOXWaL4kNbvtCjunWloVe8dAoZcALmbnXpINyGTqgQTVvEymn0YWmsr2V5n
RehzqxMt95zW6IjGk1Ev9eozKCK9wHfkfzew3oDy4PRb1/SYMnNBeirJu1bbWJmW
Du58wSDFwLIGVt+ypA40rC5rUSc7RMKLhtldCLibDuHC1FZeS1/H31mJXXT/PjgV
mAYjF+ULMUs0K5I1Udxb9G5zgUm9AW867nFsuNuVumMO15uzBawcAmumhiAf4KG/
sXyHCJRDjUzJscVWGkUv2UOuxirIMp9I0YMivnn6uYFKH7DTplHOcfDVHQ7NfA0r
ai2YnMEmnIc9zWxmq16dJWEcBLNPXKcB3htY8ckB+1kwBqy2PtlSwFgk8rqLMtEk
HPByr5xEw3qMOHgUdBw5/fj2Ey+ntnPpiygRUYmbbQjPWBVYnxGaviSQiGWFwpaE
8epzghDJJTMD9QGlGyUCyUsPw1BdNGjEGC8I4ExgwauxSddkP/d+LyPlt+D5PnV8
NmeVYFG1R0Dl5Gt0SwDNwwo02NBrwn6cXhjCA3MbxVt5rN24zP8jqPkXuuZCib86
jY87/sM5LFW+Olw6Oa+cQ3/ZSgo4JlkLSMOHIGYSeRdOjRrhbLi4RfhY1iDGUXBE
p5IV0q1Wol/qbUsBKV0UMvkmqy+5ksSVmFEGmbH36T3Kt762KWgU4/eUHg5OK5dj
FBeIjC9yaOEBmRthcB9ZBCYm1na0P2rG91FtUR3Muqj9Dk7+ovGHUVSWxKQPZduC
BG2KTIpxPamAjXzoESfSfaLTo9AUDo6ZTHsJpKKlp34n86TTl6cjLkRoRIyBZtGN
p9JXspcnLF/JeHj7Ze/qNQrv91/RQfOaor+pTd56Q5VJTlS+6/EG//nb0Gep5ufG
7GdwB/hv8Tv0X7JRY6KiIch/NJRO7XB568KvI7bGKJ4rUF1n8P4PTeMHJpvA7oDA
bAVjW4akCGjwqXsfrANSRbktuqJDWeFWTveIGQf8IV4Ml02OB0qWQDPujpuPodSJ
0Hy2VwDBCUfhnfnRjoQSx6FSsCSFaFJbFcwi3wAupm27Lv7/EeKqeeq94c/07sr3
hxe7scCBy2A38MEy65lhf6KL2cx9cIl4xekdsuI1L0L++Dgy+DS8kGkweNaMh7lv
41BXUu+0FmSb4P9MMuTxlg3RIjLdjnJqlzxu00K6OjBJg6Uhqt/S7HH9mxdXFKgI
diJ2kjAdbLjA9yfHJPQZCPk19AiIOPeydTZ2o+xvuuolzv4uQK2sRI8/DozEvo/i
63y3lh7irucM0p7+XkjtvfENdeQ/CEcnK2AySvQTM3IuXkr8afH6eDQ1M2PJMMwf
suaRWWjZeMChQfO4GVFjPxIqVUEWYiIOBfG/s7MhmvouBGaf6E/QUKNzE/NjfGuU
1Wb2TX8+ijVOtLI3JcXidYgiEp0Yqpwf0CQ+xje8PAACoJ9FylQnTqHCdoQnQ5LL
dWLwGMQOMS6sQgoCFw4aSadf9DO+izN++mNt/Qmh2DNSEEGnUoL9KYZ/AqM3yhDP
HOwkAHTT7+6EMJWncbAhKC3sHzuz3ccJnfVJnVVHgBjp0CCtpdBjxAFTDISNC9RF
ATls8Jtnuz8kC84wMP6kKCpQCPKtsQGpuUs1gsmqaNu+vX6fnssEsGDcT/3IVQMh
QYLsrCsGjFyb8gi6VU+Khgdl/nkU5CGFIVU/2Y4zoQczsliUEzCWBHOzxTa/bkU1
ZaVLmxBkvv3zN7/44/bc3poZdLbt9vTdguBZV1aTgp534Qgk7/pGwSgRHmujxjNN
/O+cb/KD3vnORDIt1xpsTdZ8cyeZSL3o9qUmeGZoKNWCSftq9/d80P7ED1vQTm9y
amLbhLeR243i3hg0GUuTwXTmUg5zc5sMHTeKmV+/sSBz3jDy1Ot74riGbz+O8sKW
wAgfiPP1TWenwqp1xt6beYaYI2nfw5A8+A6H8dG8qgllda9Jn+cbQjWo1xw/R1T8
BPU7nH7pZBLO6LLvwLZxerzGV+3K+dSJ1NlE56JK0CRyxoEHFuJAyvSLs4lpTJf9
1O4VphO18kjiSEHla8BHmdY+cNOO8fynUF/X0/SyGIKjEfpH+9Ye1g1V6v1kNpuE
HcKKOhOewFqkXRAyA+d8nZJvK10uyV10Ury0A8CVP8RxFZGDOnUv9dabvNzw/hLb
WTIyqTFXCSPcvD2sVqwrtgOE2NjCKV/v/xtdgnZw/GS15O4WjP4hGZ69hHiuTG+k
0sld6KLz3cxzFpoSoGEYbNasCcWvDPVKQD5xtwHOvOBIDOD4oe+lNGEUrpZbwkGQ
AOZL2EWyJYSrS/YNRrhPamp30ea/fRBm6Rf+BO0AZiSn4QSz8VthJPi2PBNr1/+E
vFqiaHkwXsj9HuRWCjN4H8CvRxHmWfOHNOFFv2ABYxckKaR2KolVz9rqU+HZygeX
Zu6oM8NRL09y05AG1o4RfPO5YaCuHhNLuny9+RL1KsGawtmjpLcNA7dfsGdIch5n
QQgakCK+81ICv+CeZJ/+CxrBfhTCSgnL5EUsGURyms0Ld5gu8dXFJpGkSBzn9qfU
Wfro6a1D0sTTg54h/SU2cOCZQy/SoWS4eDZne/VLmlx2QbxrC5BsRb9lyXCiUWa3
LTqbSynNIPMUmWiGx/esIuo9wA6GOAore2xVqi2BZclUrBZmArI62KJ5UcUOOGWh
m+WRnahzQ+jMQmcXd7XCxUZQedBJlObORF+6yNNSfjs6KfFe9iIHOP3oN3X/hdiv
Ph8/zso7UKk5qI5ZiV/uyfqKk6IXpG2/kK+TF5Y3cGc7wwpVodgz9bCoVc+8PNZv
L1Y8nZqlK8TSO2YtbNM/TCGsg/g/qAgHXWr6b0okGLLfiZar2Rt8Au8IIUhs1FL4
znSs40l/B0qiqMBrP/PMfwceeA+RPTvUGPuu4nzQUxP5ZpC4IhGbNn6JY+eOixiA
XQ729eUtF3Rz1U9On0+B6OcgbogbSzxKDYhnQakEo3omdwxGq9QzMGx7sAzeiJ2/
Qd4E+QoTqTKC3w0LKyFGwQG3F9PQiqii8M3IiMEKV18dfT+S+vfLy2W5wuUVUyVg
C8ll1WCQyA7DZDB/7DXoDyCkxX7S4MeDjne9PFQKEGOYYjQ2EJAfc6znj2JOfHj7
zUk3yOrclk90aX90iRpKwLuZq6hLpCCjlSxt0xG0M7tRrurWPg9ynh7P1+JIDXMV
QzAOnkzyv1mTaxMVDIAiUtIa31sgWmRhjp6L5ISBTn9ftyRPsgIJUz0s+vG6SUXT
OnI33pTMckb/gkSzdynbQbgopJy0RqYAqLg/Q4rxBvKcP76Uhe1ZvQwhwULTASAO
FLwsDzk8hgHRsXYySVcQRJiBHw/Ul+Uz3KOifwuK69z/lo7BstghfXIcXun7T+4s
iue3SdZw3//VZsNc8n1PmZTDzH63JJmgwGq+P0BPIawD5phoI3ffNIgzXZ/5YFJT
1yyOiQ77prLzxrEIcQShfgeSyEyTACWd21Sz0Gv7+GagTPvaBckJYw1+N6bhamTT
C+nqUA2QsQ6SwRlG0DnT/bZ4N4W0ZR0v7XxcL3epKbZ96MPg1gSvdKYVbr8Pdzug
E/I4Xo+LBVF9nZss8Z1I1Zbm2wUTXQ2mDhh5ib7n/r0Vf22i5RWOkBoWK2TIqGd0
ADtgVQ+SBpG8RNLUUiALZvxrskClIQXuyworJmqTvlKKuM6PUykBXu6Qnef9kmsh
Ch0SYmE4oB+uVjQwLr+vh9y0sbTWvuSRo/5bJJT9V/3fVbNmawOE/t2bvFfPjdTv
8MWE0qZF+suyoECdmpS1Sc2Nt1Who6cVQyKgXv5atycLmvDERgPEiAegBbo8s8Mw
mvIxCqFWxh3LXc/92oIjmza+LIxmDTxbsPhHy8f9/jBKH8t2lR6jJEvVXOA1GotO
tb2FSBr84w8v1icM1LtpOpNR1VcuBgvb460pDclXu/N2pIqVley9+5SySXQpo8Cm
EjgqGLvBtppzKDSDfz4FC1w17i/qAtk2Qq76YEoGMo95QiL9/ErAkRlGTX2MrA0q
oFXTkc4j9THauL68BZXsBpZyij+QdjheM8hqK7ALBZiXkE8816g7TWUwzBoCyk/W
q2mAXzP8zxaOwKObO8Mjk/VRq/SbhZFIge0VSUVRIu4R1v1SXEx3Cqo3Rav/ba91
0P9txiCEsnk6v5B/NWcKIEaN5/nYVr/pxHY8hVS97tBVWAHGX7tzzE0wE/GDZPhz
4HxbXsQDdLwGKpB93dXxIIK5pryFathis3ptpzXThz9TrtVz58vMzPYZKfG3hv1x
exESGLYT9dmqvkvj+FXx7hHBdQO6uXZfLY0IonxmKDUcuRqoudpTsyHvR9ChUUwF
NBTX1hSfImLXmo/VMdq4eJfHyT27tc8j3onUzEia/iaJ9FRwA3oDAFLSUxQSkxIO
XE6cGSqD8+85OJUdjF1GckMOZ8OG83lbF5rvhwiRssm0EeKUGzcess8aupIy2OHX
l3mFWNJLQwfirbfvMiHEK5QwcSbii/xYGhJxZllhSc+LBPeRBG0ONcdZuB9Mi5U6
pnxWD53jlBFWZ7PMjO8LBGEnNkBAGSPVKGHg6bYDRp0zf/cmlGsqvYZodWcQxyBR
MH5ntxqfgo+rz9+NdE7zoAalrPqc8NgyBow3UJn81LSeLwxh0Zqv0UsmNijCcT9l
dQjk2R3rTzvpXVDsQg2vW1MkUg9nmtX+wxSpJQM9HqjD5FA5+FFcsirP++1LgOpS
ohu6WFgh8dLm+PR/afN/MHQWP93Aia3qG1mlfeWUd0n7q+fAalUCo0BFSncUqpBC
sCxhnNYvRsNkUR6SFoTfE+ErN0EbuTj+Cy3eqqYgBVplaTAkDl3CMnZLY5qJJKzB
xsAMJaa5I0fJ7rISsPzGGLzdHjHW6hM7w6OFtVbpjAXtWlgswnDU8OWuHT7y/yqg
zx9KYcj8oBLdtHufbwx3VeYkF7r0jqhfmzRSL2bNcMbL3vWg5XeMOrTWazMQJwn0
785aO67h5iH44uykQZcoU74Mpa6VmHC/z5vyrgyQDwVjNjEKiCVQZSW8qEBBQXJi
/hBdVnvQX0Us/n/WAcbQ77+K8Aepzp8Up8eKGyhNrEm/IxZp9EklvO9atdM/YX5C
l+vJp+JcEMkaFye3FDTZTXEbKnFZrgJS1hYz/1wwrC9j1ZUf7sH7UOSpcgi9UnDG
71Oj3X6kwWguT7ABjOptz6/iBXjFa45Xz94k8utygALTj6b8/ZP68oznE3MamBrl
GTWDruYpDbFX/2bF1Ho80UIOqVlgfa7kospn10bn63G9QvW+bMTF6KeaE+wdJW5C
rdyyQ4QcoNPCzeIzMynFjyuXggb3RkD9obby+seF4S3PudZYmxNFsZUp+N6XZG2o
1Igiox2dffkH9RCgVZNH3T1b9woXq5WNU6bjdO8/R7xZbghsLykJV/tvjl9hjlvw
OSdCP9oFvkCE5hXB+1wkM9ctaUFAZ2XyVgdi2lvaJ27kXodo1r/OIFJXEYi/oSfq
GxbWkFcfWuD60oU4CX9tQ62V/36XVBrrVHJswaRVwhTD0tupazGJgsjiX9LHCQ1a
eCjpDo8QdTs1OAQkw7ptzR2N9s8nu5oQI9ybumuvQ5IW0h4O9DlSRrBQM9HPllOI
gZ7TvHqYg/3SbU4/chpaxyAS9cEocPMcM1cNZBc4WgEz9w+YDadhvqIAfxzv3/EN
+3TJqKNiSdYFJ5+tZTK1Sq7N0nf4ea500DgTGBBmC4jvSRAhccWTsFewUInSqk0T
ucvki9Vxb4om3fde4TaUcoTPvu8nUXnREZzg5zhUTwECpNLDH1bZ8T9m8JeS2wWP
ugyQIOjTd5EtC49hiRAJ0KqFYwXfARMbo2rDFRmTRoCQfYYVmVKOsYcGL4ooJ/mi
zJXU4DsjVgrPK+jYV/iE3X8OnhaqbnzQqladyWNAOYgjdm2cH4mcR5BdP6AenUzD
LCGGSAag/734EHhjCA5R0AWYKQ8y7PiC8KkHMghHwX5u3yMT03SLYNK+hO4AUung
37mqMVuQIfSKXsmalRjq/ckmmjSowumjGsaz5SNfGAqaki57ZjTi1xD8ilsoEB/V
HSYLo0/r/95aXEXIGzvKzs+gvxmzcJGzOs3IVJCQD1LQ56oIwE9sdYEgBm3p3ksV
1hLI66JXGHa59FqB/+ZOEvMmeduLR4CscuSiUJtAaLQ7OEVoSKGhzKJBcw4PXV8D
/3bqJAGFoVhq9dwm1y4YOk4LredKw/rJVgIukFFxtIiL72l7bPwt1wYArj14DvBX
LWsqipowOpGWdHwnLPBwChPM0pmLMOyJFhhb64cPGUIkv4Z7Ue5cxlAmvJkBPLxO
urxatYZwhGZq4EgukAPCE4LY47NtEghzWjYV3yscbEICXlKndkCBI0tlbvP5KFT+
77VwwNzA8zG4pyyb7kVG0jZarCbnNKho480ZZv+EZSeqLWmMrDfdjLguxIQ7PrOi
uYIgOPNOY2kZTB0TAYMKX2X0xWq37ysXRYRoMei+UBa0rsP7L+DCQmTmp6YnbzCm
qSXCJSSlbY7H6WTpRXAWJHAzj+rgW8xZwYVBYpP/N7ATFRLs88YJJ4kAZzphWLWv
w6u4P8++ryhIQ2miXgcZCa0Hu1qZt03vCtwaVwVbje6mhit01xzRmhkLPpXOsW/9
cvgoiVKk1wy2SiRXa+bJTZC0xldWbks19DxyOv30cfU29u1sfbHims2lOj1hVl2Y
qDMKYii/yfb9GePb7hF9baKSeV55/WhTH4eHEBSxUCPP2hfGuXEaA4aa3YGB1BTy
BWz6oKUapsaMv8OpD6qgDutRQ/gofsquXDcw2sE1bBs4qH3pKiXp/3HEYf/G4Y0l
yeXjPaO5qWaEqZc6/csA15rOI6/nUEj5Czd26yqzlLivN0LxAZtv3zmMa1i3JJXK
mNSkt8YmR/52GIxymast7k+KO7O6EH+nW5BBL1Li2h57nnJHGzVqMjm88qPmr2jY
/+zKnBtnZmATgNr7hUvWrd4uNDs8ONpVnW/Ql21cDZMeje97CPJXDdwBVhEZ9hLm
5C0MhVG6E1t4KhlIyHAnXqKYQzV5Wrw5aDHTniB3mh7oZldnYly8QL0JPTxhkCbc
G5XG8xMEMMEBKp6YD6zadN0wiTu+5AbQVAXBsyhhix7riKHqAIu9FW+LTR1z7sio
4ghbJQH+7QcVC24XzG4JsBrBugDEYQ2Aq7UnQIu2KIl5NKLT50Aaxffy7qd2znnt
htmRCvTONNJvtzcaKtIraLpnFU0m8Cy4pGDFLIHWwVg1avE2C5U1CHsQIs1RWCtL
EkpJTfAssknwsiVzVgxd4grPgbh0bVEDhA46KXwWBTK1THdy3OjjtlVasql4biLK
CeBJ4jCvQZ4yr5KONGqQSkY1avhw0vKyxQdtcxaxMP62P58tmL3zxccYO75lynWh
by11A36/b3ll2C3oX7sTPnI97TKVNgjuHG05kqOf7yksiNIVnCmsPwxlptuFd43d
GiiwPv4KTlJiTFNw4b4e+ZPi48eV07H+LKscuuaYzbeWXNGXyG2ha1Nt82EDpXHC
/yBb+dh55SB0HcKbTEvp1NbV7rYqrxbc51sdIQ82qr0ZTngX/kQy8+H+afWO+IJx
rl5InXjq9mro2WYwS4qbnWcmB8a68zbax4wVtdWuFigajF72ajtUEpT0Kh9KRqPU
yo94RzLxRemt2MbaFbFOB5L066xkQkka4LOTRZFCN5wHS6e+8kab9JYWCb7npBW/
W3Oin7J3fKVpYyU4DB6qMekKzMvulwkBHlGUs5ngPZVkp9wrbUQXH+WlGbGo1Rxu
IlPtEuv4gmnAeht8TyHC90zPxmjpuYTgLQpnFdwS79024hSEy8At5vxKVaJezgJb
fJM5KXeNT688udlc8q5SJus4l4SSHLfXLQdD4eCXIiBNzgOewyu5O/7pCTDBwC33
OWPZN9eUfcFnTrP5FtC3aw/pW4V0G5+dqB2EHN1xfIen03FmZCwXnNZ5lfpmHrqw
MvNzT1G5fMH0NPQeCJnZnjsx5Wn8pXIGtK3p8yeWt25X6yoCFZg6MHUUgGNBWg1I
FANmxY/kDHG83OGGz/khoISDI6ec5gn3QY4Slsuv/OVZKkM4vVfpO7PvLnk0f1fg
IM+ZB/YWBBdybqT0+EUBy03tLVgI8CVQUStsjRFVGHwwhR524IgZLGtG5lRk7+LS
Fnfa+kqZ8oZ+bFfHDOxsw1iyBMaf+6Ez3ncgVJVWSO5rVGrt02kmh7D/pxdGaPTU
hC4gvMa4WYaExvIps/VvnaPNS99I0M3fJoverL/6fSuyXwmfC2eG9nCyri5zVCyt
AbTI7HNcOWbxyVInJCvD48w2yvjs3g9jLrCP72wyiO7b4SEsE0VJFDUMvT3AUzCr
J1Jq/YHtgfK0ZkttawSEpeYVk2pBb6316NuL9YBxo44VDyNq8XKYkTdfFEhcCZ1O
fRvikcwZFGFM3YwYxuj5N8//rRKOBkVs5q95QEwUPjODmF6bW7vm/3SZkiqT/k27
9AKtKaA63RniT9mLW19C2Q1k0pwZK5qh8H7NXdfUqIulqPrsBVg0AKpqvyCSiobR
lxASyNroq22tuFp2ooeeSS22shmuoL+GU/Xm3/RaT23GLw8Geghs8BNT0FcMYQzq
MdqhVcVzYvAwgT2t9le9NIm+Oscbe+lm7JSrxrKu3cxxlHMwmKE7LfvbkyBurk1d
Qt4bucqFALu7vqPIFYsYCq28EfRgd9SGRzV2cHxUFjfB860Och6aFjj00OiQ4FtT
brlClX9jStI9Hnsm//V39QiP5iuMQYs3Xj04qEOblY+AuMq4L3OhUrmrPJ5ks0A8
zmarVAPJ4b6F2oDbycQRIiOcd9zKbQyUxbc03dWPtlmt8QUtJj9aLSyJocrVQieV
zik6XHndmxx/XbjK334zenmh9VMf5WuCSQc75OjdK9GCq4dnF/ZY/IL6n722jSu+
7VVPEnM/DCakLn5E6PYRDbcDqiAoOi/lt2exr4zctwrUF5Hy20LbWOwfBKJJXiwc
3SxKRiextuy7P8hiMyctxgGCwqCei7QcsZFmy0YE6PBy/sYxgWf12xDBek0UyMoz
9mEJr3yyCPoHGqCVc9/MOqMd6fJntC2BRJAM97n1qrSUfJGDvAArwxHzk7jVjYoa
pftADUOOBFPMERdrd4eRE2VniA7YZU10J1Djyb2kJNrofKi5drdO4amWhBpqQ8ry
WnM79xe3hq2CXuTa2P3lOIyy/4slN7LKfoEgjzAbrJHYEvYe+Jy/YUrRtKHJ7wLE
Bw/it9ZFYeraQd/QTKxq1CGU3srLg42IUMskIfp80NnKDY3txFFwnHadYPo4X1Eb
UrfXBBTQHmuUm0C8z22iJSkl1qqDYRgExTLV+ePM7EchVJmEDhDbxSTGUd+8Vg1f
j3vjKnV5vETISdJItWvOgouJ7ts4d18pbS3upk1YFoE0jaoRmFCambgzr/X0kQPu
xbkrrdzEWmGihygGzy1uKWKn49Yj+125EPtZW+nk4cJJDO2e7JdZpbQNpmOiv2E7
sjhnGNFVobWLhsiA2VhH3ZsLNG2Y0S2FvfVReR0LYWPdIdQVJc07bdOvMsPLiRTx
ew3hWWAJeNeCsIUE8U05Js4PR2MIzrCpNNcuqFtogU2E7TzWLeZww3iRDTcvyQ/9
hjh6gVyxhBMqVvDKJlbmx8Mqgg5E5cW1/E051lxv0JbsrRrikPqHWfGYm4GoWGOQ
V0u6y3V7vW8YRoDSePAoD8JYOZ3j1Vld82RNBrKzx03w8iSOCiOkkCOyLYpi6eha
nULO6dvQV0r5CybLrKhQPKOGLkK1zASWB9ViOfActNURi5JYUC7V6oFBaksPzZ9b
16DCDUHdfJPVn3HYxAJ/sMp/jMsTOwFY35n0eV3CYKFxMMLj6dyK7mxthGsRwnNg
g+C161rj4g8V1O1+9x23k7qf85XkNH3mImxMFQlXcolZVqina8F65pHC3sYDcCLp
dWWD/fZtJd/zvOx0iFz6hYkUey6F8wf73orMQPIyVwHMkJbnB4x/z+kvoKGERfUI
d9gwPH0Ffbu57caJ6hnOkGVeFIEcWyVD22B5w5hgxHqUNUp/9n/r2X3NG6XhH71C
fMUSp1N+ebBW+aTaGTTtaQD81FtT964D/eEpC1McDSdgLw1zTIjPbKbHaqo/M/4U
7wd4v7xuHYDBHnqCJLBaqKVkg+5ipgWv/5JmE1oF2DjoI1VGOM5KZzA/oTSq1a0f
kut1Xo47aiMdIh97ZJJC17eHuBRfIK1h+lGuRfqKcJjwLpnMeYdyba46v0iH1Y4+
NB8co/9iNiXLUpi79+Eyjr6gPxSIFkNCgJPxa0QQ2iN52P7A+Dxkf6q1PrJ0aAb0
pnbiOOEbLnFhJDNkCJ7UrICAgTKsDLadKeFq5E95d/siy592Xao/yARmo8kvWZiW
uVlEXAt8ZKAK+zT2pO3b3uZWRtucv3Ev1H+lbWO64g8/+TKTruSN4C2eK7oFWNqK
mm62iUBdvIbszCso+xH0qbHxEc6Ixq/anSn4sOWCfR+BmchTzpq1xe0EAuChokiz
2xMQ/UsnYZZfPuN+GwhTQRMDxoRutPzgAaQe4jjl1AB07k4EAPwQ14+Q9Pk5lx0Q
S/Yh1cF0O6AuePCnKQu3z4fmJ2KEgJsj7/7RtVIMeY3FYR4745V9e/gby72S6Ax1
9xFlQ3Le5VEfeNRbE3yKFzdlT0QVRvUwiRi44FHgIAqIvAIbP5tUJQfLYKfiAzZp
c45/+tEMKzkMcLFIfcs/EHK610XyjLdlzOQJf8tpsFR0sqsNAZPwuqlMAaQ5qvi2
x9IKfh1460gm0c3HAnR8XxPT7RTXn4VGOtsHBCgSnKxwvHSRVLKG5tzSBF1HF5/p
HcFh48iPHbtYa3C3JQHP004m0y6ALk0TReBRIzOp7QerCyFKWYYt1PLQJmeCUlHU
MuE2ohAC2VzXOvGqL68/C9r32szXm0UPkOzn0qp7ZtxpAHw5BRY4P41rs6JQ0RGr
R21S2reljwfZT/5pEjw9qCouQmY3+OcR5PyNE7y+wLGRntfhb2cbb9k3bvlNweJC
zy1/GXOiAhgnwOsoYRCMXWInpAN7J4U/A6V5lx1OHZseBb/5/KxyLh+wCRWKrMNM
kRcpY72GecUT+uOF0D4PbudULmseuyOYh29lorrwmnUj4ecIyQk1NaceN8E2l7zN
QQLx1aDp2ttwQIN5GaUhOLIa5c+0/BeTJcC5PBWRuChYIWrK9xZDKmj6n+bQJdc+
X3cUVrn1taZXCBy6UJdjPEWFRH3K3tP0cvpJRqcss+qntG3N0GWmQJYMv0wo1xHP
1wdlddYUn5w0GJSrgWQo4beaL3rp3fCQAA4UbySQyiOk8OgQ57qTMB5yMSbcPuvY
yNQN1n2H5N874RrDurMCU3Jl3hWUnxDFo8xPaDNLMflo4JImVQjiEG0RX0I4WXrO
ndfBa1CCzNILViHa4H1Jz3VdUqiQGEv5C39n4ITbyLBnTzUzt88UcmFbQ9HdxFm2
+SedwoOFwIL8AyxPFsCN82Dq0MG2n5W0VW13Bdp2/Y5Vdg+fh3xWbOiPSIRGOQZW
iwY15jV58ra4Kn5RqGvy5f9eMDzF5yl0Gb4wzrrMf7suqzBxX7Z62pGMrJ6+FrOu
sYIi5Ts488p+qkzNa7MZLvktZl/1r88BuTO80JRsmQq8oViJQHl0iKt86z5WIrSm
aViNpY78nfbroWi4BhTq70U1Pn73PkAyJubiVyNKCkVOucVDTEcE+KRlpzzx+NdP
SBa2peG+iLMGD2FF2FtAuqv8P+RJZZxXg2E9CqWXQbWWQe2qdmJfqDqW+ng0Puxw
XNIeCJBQeWBBNk2Xi/X96FAePxkCk9Gv6EGolBwrovCls9pCP6upQQkal4Gy8F1o
xE4D7ZIGs8Lm0z/VKax8zj/WfpRK+opPm0EaLfMiFqVv1nwPRjN/g3DXQV0jXvTd
ztv0v4+PAe+QkzNJneJ98edoRunBvZb8pw11WKs5vI9VWS9GVZoj30sElb2Al//s
+TToXCI4ZZn39uz72eclYAL+pLVDWvmVbJmGdB0WevzCoZiSgDV2MIJNEFXb3jIG
GrMGC1YqcfxkpQIw4cz/rwYtcwEOSlFgUWY59IvfhdcMf3/BG52PkQP7a6uirkZC
c5UlvWEYtEByiSaEof+MWuVphbrj2Sao5YUL76etcfbnCbyMa6FoyesPizS2orJr
m4Bxp7XHwsHvE+TJL2aL/d8UohixYQBnzuGllJSr4uPFRFCESf0tvNc5QwJwANBZ
yKqypogyVwOUvXVl241iAA4ffolsp+SfxgvUEa0x0MsiYYKOFnWP+pYuxWd6eQ5j
iPGTTQptv758qmz8dgLUrTyLMCPoGyZ1oGZmXRY3HHk/qyNbvSRiv3/04tOUecnW
CkYQ5ULax3BoAxaOEnHNzwQNDLOXQHs6uFBEAMROivF+PWngkF6MD250VImageSE
Ujnzy+1U36FAHu83178ep7xLQQMEOtc3mbPQZbj1Fkxc6FaEoNm9+ets9TrNALwU
guKdA+AHYIKzOOVXWZT3ZSOjc1tDuSNk8gmk3/mlTJlordez7YP7ZcpnLk304Lnx
eM3343qO5COOIRGq6ZXXsOt0SCg0FTydE5H/un9mQzNJEicrIcsFNi5xj1uhLe+Q
ENoCKsgx7oIvR0p5ndeUT3MdUDJ/gSkJ/I245VEfilP3J1X+yGj1Y/5dINCfuzcm
++RBFS6N8W+RSBFmLiCDk66Zq0EumvPonZZlwD46BXCZGPVCl1NwIwBaeoZgVDFh
u9jhHf6RvQklsaNB82zppzOH5KtSKJD0yzK7pkq23wKksRhCnEUMaJBS0iGhjE4f
mPKt0z58WcJsS2T2gEYwALw3ASNULJnnLWKD9on8UTl/LCwpX/xBu+Hq74/hutGv
q/oLOr9VlRWsMCbNraTOQDREzEp15KmUvsvOvmtn/Ae0Hc07XJe9v20LGotShboU
O7HJK9W0VtpjKYcHOboQXNPm2+74TTyshi1Tib6F0i7NTIWXEnY51M95yEKc/eoD
cv6z077PeUJ1TAfgrT/CQzU7KpNkC5vhnKajvfxT6uqH7NFyZ9xUaZ/ZTT5hXiVI
Q8Tpphu9h7sc8/NYtxoPGv9wwe8/R4NXDBgknsde13TVYDf0ET6GR06cCkY2EswI
vfzM/tBFiSOAnxzLROvMnzp7ikO9x3OT0gB5Hk95wlJGDEKcQf2vuVw4pIk2U8D7
OueIjU3YE89nkTZNrSdmheKQFmJoM25rS8QXmFlH9TrdE/By4ASPnKPp0JNboT6F
P4xH0Z53pzkhCMX8i+BUuJ5Yf2gBB1RedSQ8SHhxX+Je9o8fR/f9PAlAtEjd+O7s
Iv86zrbDmxHYQY+uj/Vx0sQXGJBCNF71/pfTDvuv56P5CAdIMeX83eYHvAwmqqu6
X0lkrOuSq6o7r0O6DwifLx+KHo5MJjNqJhHdHcCJLC/NDGujVsKwpFJ7Lh9wr14l
iHkJK6ehldD1iWFEKBTOPGsOzj9oUd/Y9FwO1/2ED+joi8YkGz9+DkYvE8aa6x28
87PACmc83WRgfqvAxGjGSF4Fqu8K1Q34/SpbCBHiqfnzaO7XXxQxTRHSUcDpscBq
eBiHmAppTpDF8u2GLZBBWORtgVkuD1v9T+isO/g9hxtdazaJVXptkdKs8Q6tRCzp
p3VxAf3Kf0LtLA6r/MHlQOhdyMpt3UO7WcmFEuzefwMaE5bEEEtzTqrgdrruQC+K
ieSUlONm+JF0saHzW9KPZ3cwcqhcDA/ZBqSV/IuaNb2szSPq57HM/X2VgSJc7rWy
0Fh+ZBrkd9g3DOjAEfswMM1Nh4oUNh7L1STzZtZJDIuIj+06lvBUil07h7+jKilU
/lpAkSSJ6uAm/FRnRXoltE89EIl51uD64NiFCUVRbPp/oD4VmkJAHhuZbt4Mv4fb
CcViIxJGqKR66Jb3dmAAsnVHzQSq3MtrTby0U91HBaoFl3Rwm389+4vm1umR+FzR
QZoFE+dk18mhIeE4rO/FruKF5saJO8j+2Cky9qz+9wcDMBT/vhGdlNcVn1OrFZkM
I1h36lyYXHG1grBK2fZoHYEAAsl9JcaiEqf4psxkVIHFXuW1Koc8G3j1xqkFhAaz
yC5RKErzNvotuUqYlkU/GzAYbFEvWANmsuHx123MbNGWSCEyfWEoynJgNMZEebpA
qEQcbmArYFzxk3m2VJ45PluPXc2pXkhxob4bnPl9mTW+PV8UreZTxNPCO3a2w/Mt
XblchFpaE0lkYp4qRc+etH+ExB0rXKZvSvLO0z8gtbsEcowmjxcDs1k5i4q3J1lf
9jbBJkJoYwTlnZID0CoqDF55C7s9qlvCK2pt3kK2OBuJ/+RAqUu9+kRCvW+0Pv5+
5/5gJDDgD5F8El4d7YKiQKDofoVAqWLaN9SRqcEV9hIUmnLSCJBjbFsSvPkSYoMI
hZuf23MJjexMzOG7bd8JKh9dP9UV63otQ+XTySlSYqJgKUjbP7WyPtu13CN8j7XG
iUSA6BCbaphFaarku4918Cu/HFwDJeCG9KvLv3zytw/jQfBcjFmRdS7oC0UjelEu
Cy+dcCFO55XsO8yvKRCB+bU1keyj02l08IjIUP+6RgGQOoKvI4vgV321qZ2QX4uY
O+ExDRTxMJ5BUJIDa0QZINOv4h1U3PCtnyeE60+8PB7+TiBXUft8n5Yq+1X8uctD
u2Uys+icnV9gz63/2gpv0EbisW0DxCkMqx2xfifrdeU6QGXTp5YWkIWoUON+m2dc
zDtD9iEYnkKpPjAe2oLHFplb88PBUD2W8V+PM0AqniLSDYktcGyUX5kBfxCq94j8
OR0zdrkO+ujdReYe7kPSlsQRQE82CBglKE8+k7/Gdy5U2kD5dSRGso22jtPvMQLL
o3x6rCCpKx6jyTWcB7xcW70RwcQTCVKQyHqOva530B70ZpDvC8c8JyYPpSiSUAsX
pEhs0wElJVYQEHHr5ulK4kFtvvYg0PkmbuXeGHRop1+M/feSHXweC3hrFj63ftyA
q3H1lIuq5MLL+u0CNRUcx2IZaY4btMB5hNsvCGXQM1ed3tMUv3o2O7yYZQjp+Yp0
PNyc20t9xYcp+s56uH/2RewF1dA3hEStZWVCOhYTSp8XoHjPY0mNvlsJ4eVd2rBC
pghEWtgcy1MP4jqOgYaOA8llnHkPQyc+8YNIoRSpGrmQ0CvHFeug4OETtW0kTnmU
sN5ceuBP1o0ieZ7h+DKogtFBuUuu6YRynLRbUfkbJoK7362S4J5REp6MYs2HyLE1
HEWz1+P/pTFiDXsAlDB7XV/hwmaDc54tpdVfmRUBQS9aGmFQFgz7lFAYwNzD6kKB
EJY4E3a7nVLrFcQfNNm1AoE9FCcs0SpaZvkVrWEHm4FWkP+CuKzlbcof+O7P+Pdn
TIHXJJYyLnqN7J4RYeje2Q3fZ0lOZwfJdApCPqLZjiE3H+6kIQPhVWob6/9FcXlC
5WDFx0jkuguWnBb3oAbFjDSO882wMTDg3hOA/1DEn6QN382Ly3rlE6inW+ZrOlkL
VQaxjLg/3R1esKurQLqBMehcs/J+s8znyfwjvTlVUjoNsgQ/L3MXM6loz4b24GlS
aU+88KPq1zrwhqGNlH3JQd9QMm+w9A4Og4KwUe7Ky4BwJDHBb+Bn+37HqtM/kBHZ
WWZ+0uBvFs05zd2fqRvfvtEEmAF71bzH921buXFPks1UCeuFZBQTaQmZJG5dPyl0
5+mkLLTZPddC6zlMP6sx9gjfovhLtcP7JKKv0sgOLv8P5rO++L1zQc7YelJT42DH
auVezUo+2MfeeEpZc5mrIrPasV6CU3E8Xv4oPJmbnXFUSfvpdhv1+Xw9K8fi/R2f
t2AeWyRR8ohs3gjNIR6ZnkNOMV7t8Uvje2yrk/uMg2yG3eBSz7PC0pKXYmUUkoXb
xeA36PxwokMHj17nf697UqJ24Hmx4MmXlwRpnpDoRdf3I6VrnyHoTKl3Soq9B+KH
SfY029nM1++A0Vj2vI43DCA9Gh/nttoeCod9aFfYGYsnlAbygUjClrdqpmeS6F6i
jp9Q910SuZD5blYFxhB71DXgpKRpfBx0s0WpxFc5eNSYCFdLiscj5p9eIWfnY6lJ
NyBqG/8qWPsW3EgRGZgsqW6lEAcZzLetjDTDmauRwFYCjvkK9U1LR2xxg+5mDWYV
pIFrXzj7CCS3SjSn84ynxkZ5j7hjNAjDbmUsUzlqox5oHlNuQHlLQ5yS1DMbU9Xr
4WlLHV5v1mgY28qdyvCmZ8fzPcJRcinPtuvJx6+2PWHRIVdDuioKCBS5CJ1loPw8
DUAWeSrpg6+5oXmMTdvurZA8mtbVUPt0CpvdvyiysGasmOYfpGjX97JTsyP2ZCzR
/7GziyBjhWqqq7GBc0zAJyWudk6izbRnDZZvgUL0kVW+pqfksD6y0mFn/YAipbUp
kFcIK69tCpuUqkw+sGl8cZZa7aW/kZt5yc77PM85VXSZ69XJt9cGFF84bT/emE/v
u3aazmxxwqmm/iC6nZChsF+ZCfw8aeDNA/6M4gwMHu9BJFblXMl7AT6DCsNqC9BU
7fuSPe7uHcCfidfMicQErd4zPFX4gZUF3+9dNKJ2dDOZq0wICFcNbmssUedEc7UO
SxYjDeH9e6yo/90ZaWYOLsd3MwKX8NWVy5Xe+kaxvmIzmHP/57dM0JSb23kzb0qh
vBrwflBS/gL/v8ypBFq4iCAfyt72cK/ASS2l9auYxurwy/nZDicq5kKF58oQMKdD
B19/FCy6rW0OjN4FW5NxURXdMjgmzKr7Yje8PFMD7lXQwDqTPOw5o92rh1Hb+W9t
zvoToZvqEjfDLUO9L/VC9r6NsawxDw/wSMi90zAGj0gjJ3c60qgMzWFT6sAD8UBr
/xtIOcfRvq40F71u+mHlyWDITGmm3KnmEMJVPUx4s+IoNqrnXhOWLK6TcLGvP5Gv
elbQSTV65c3hxaT6HcVU3nHqiac1/jdL1qDNuziQFgRmn48kw7o1QBl+DyfR/4b3
FpEko3pfAETuRyRyATVHmYfW971neRZ6xZ2UE9poEArWjQ645da3Lt+cPHmW5wu6
7H5OYma8Iku7VMWESg9NhY2iGrwFiFlfenoYkiDIg0xXGw+10YNEmcbHYCSET2xQ
aKXGtCkQwenuDwkLMM7KMVKvddA/hZA2WYPwBTVlrBsIRjlVuYMwHV+BAwRUNZfd
DX3SlR61bER7dQM2PgxlVb5ld1cp9vnFP8aUw4Uj1In9i8kkZ0CVuhLr2f6CC/ok
J+L1QX7IuUpGfbttwpBfiOv40KSSmu/ncP6IqHDJiWMYa3GVcuDyV3GMupx5TWVg
QmNnLCqLWtlz/JAEq+ZS5BqKjVr3BCKmCgGTaOrZjoAxqn8cQDbhmWz2rjD9Cod3
sHon0f6TZ/sa3Y9TRw5uzZ7wk33aUX1QMuCWaFpb7COgxua/ZGIgB4D6ZDqO9j0r
AaVWxUEkI5/w2Fg8qpJ4vSWaWlz7ZUjdDxgCLKLLSqKCJ4mbpewlR8nyaZk9zJjA
9ZYmoPjthugCTJt2jSt5d65B7rLaKBMjaNVC9nt4prDPLBHGlvFIS+DmqPqWgcQl
NeDTufSCeY9yz6F6jd8rpHi/BBjL9NunpRRDUaloU7/o3ri4PUQopKpnxNmLxV7v
afNq8YalatBJ9XGi86ApKkzBRaVEzPzG+ywg2C+szUK9yKRRAlsgLBW1QUO2na4d
Wg7SbkmNPmKfDN289zKyKhRvtVN3zhaLAn3Kdp1XF4VCDZR7U7hx5f0jIsXksVPH
dBPZnD8kOA6Gm0xxIifMVDONdJih6M31qASwnD3Xvft/dq5SmR9CO+NBUH3RYcS3
tUnxJX7lBb5D0M+VmlWiKCU80fnbCXyzYk1H/4Tsrbo7KRWYqTXLh2ByEDD/F8Sg
bdjBKsQ3lKh5tZTHEDiacJ7lCCtSXrMOl+XBpKagXRFVRhOy8jY6SKjmK9mLxfvj
RlpzaQgAJwUMg20y7E8fH0dxMejOy7A2ECJIUO+o4/W4I6QU8B91SUweLjx7wIyf
wzyFvoJcUiUvZwXEnzE0QolWvA+r1xx7mTq4h7pBlJnht1cjv5cgFeNfoLRrWTKT
CNs9G2wP6rmyxKNoSfjdAWPIqw5VFE3hlZpzNo8SIPGp2DYnbD4GoYDczRgt9b4d
DRYWjcK8xnBRwbmFKFe6RwG0/91pVAQctCt4ERRsjWzdcUkY7ybCy3xVsyYRHC8n
Y4HAaoESWdDKiA3qEvbsfuDIRaCCJ6g6D2ArGjRY9e4Kwc3Vkb4NS8h58p4wn1ZO
YaeGrABwJBd2n5b5Bpks4oxzE6III0aFBoZE+iR02b/6YEaeOGuJXcI6P9HKUUEb
efYcsHOgQbuzOwIm/ldRR1PKaKPgpRwaNxquhU6PoGteKvUi0X0n+C9QX5ahdZAH
vhDj5ORJQNtsxOWSoQF934VGn4YDGuose6XjvIAadZPg8Nw01DrxSmWBS9AhTLAz
4DLmuxmEbWB1MoQR38WEWT7nebFRKw/vAVRhitlhdUbHk6Grj70w7zY7InftpBQO
OyuMkSLzNbyl9oPLHy5GZUoSzlum/JetaIycJ9Sd96oVWaFv52BmZom9wO6eaCRZ
zQMUNaX9t/SeQAhpUQAUntGTef9z9QI98P01wndhJWGKzHvmJtAkSS3EyeAABcpM
2Y2dhrad+Sb9A9/y6YUJDgs9zOpIHs374XkOeEYgsEg0UQuM4hb/56Xg5MM8J6Ok
guTuRYxYsuyphNYhiE2DvNi493Fa2JOEdQZH5vetfvJ0rcTVWxwTnNgeyGMOSssb
+me5FBy6IGF2gksGI9O3s0Co5R48/nR5nnRVHUyMFvxHV8gP3pTfIEGp/g5QYwYh
01XzKFQ5MEdtaeL60xQhUNJcYKdnEc0FdApB5ZwlBfOC/S32YpIyhTG3iRtzsKtl
M3y558/RScZjfcmd6z5gw51w2AtGfI9l5z+uMJ0h2pUjUXGNIcEqoJ1xT5hkQeTX
Ie4QO1NbZ7AO7AUSAAPlYDceB6JYjmzVKGs0I6iDzjRJAsSmEXwTRo1ovLVPnYLq
OHMTczcJmTJ7gqEEPDaEoxz+6Klkh3PRmbwTZiVj/EeavpRul1SD0ppv0I3w53Zi
WpP2W9dCW9+SDsYdba4EWN4hkNRL0UWb2sWDgTAO84DwW/C/R/gmmOrhcvBn6VBr
BGSGOwYBbs3/5Fvc337vZSg4XkncE16l7qiAyPZ5W2GXOnB4m/QvBHeSApDmGNs6
CuFjXDC4CDg7jhjp4u9jLf3Zmdv7VOo8m8rxJ/pWfpElszORL9tJrJEd3KT9QOld
wxpZe2C9bxt0Xf6anNJESLM4EPgC9/nXc5cJIXbM/SNiix6YXISsZj+mLcEIGfUj
MCujkQMzlLY3BL/43VbT2g/kOLl0ZyzGgfDsnaL4b7pnpq9F8z9Br0ZQ82QqYKp0
fTqzOESonspShdQkgDP/duGqCz5fCw/bfRnBwIQaNaYPAlZOt3smPCKS2WZLr8Ga
+B2OFDNg1p6MVWSWxO0hLyfdjH2yFCHuncdbD0Gxeevj9Xr0mTX+bAOZrbVmqHth
xEyFZ0K3D4o6b+MSoKkEDtq+nStHTCU1FTuq+WTDsXMi02dbNctMjYsJ4ha2y46I
wVVIh4ke09l7IuZ3HQspfQdu6cn3nXsYYmG0B0bY8KuUG6BUSz7hBEeBpRSVdw/P
WU6/c1dwsmDqJEJPsz4HHOUsL5eCFA4n2gSCGDZSPGs5B/epcSAMxzy0vL+YvEQA
TvNHRC7hVqIXAYBhv0v2cVp4giq4rY8K9i16is0fZHMLl3pEFjcKKnfWPqp1g5ry
D9TolM1dV+u1kuZr6ksWlgYD48g0yEikBWo4boq2Y6fjPIkynzjG7SfCsGeYJMPC
4vUj/vvnwkY7P8p3E5kiTwylTvrGrMr5pa0p7g5VVRpTGMcbHUYZOiFjg067Z0NU
mfhijRAxmJY9t3Ddh8JkLH569AzQrzPtOye7FwtkGKoj605710eDAZ0ITCJig1F7
e6T8u+M0aHd+UTV/fDE6mYXp9VTeliBPxyykMPmFz7pcnzdGWzBD9vAmeTr6rP3x
03BwNvIm/zM6iuMkOTRti7MHq44+jgNCVlWc3Ewuq0LKtlCrP6RHHKb0li7lepmy
nCV1xlGfqs2bQ+JHQ1sIEz9FkMiES/vG/7TOEMCpiWWhL/EgFzuRmb8oBJQ9PHkp
8JpRuIbT78TSHnQuP/Edriz31LY+xpEWmiYaXNVd/lfh2UVe+pW8uFOLk3nK5Iqy
ESEqMLAFbrkpLvfwV5sQomeSan0dqW7oo8XX/97Hu2wfiaZaZqqaoq6Hk3bdYsWj
Wdx0VFcVxgiKWmTBRti1gUZ2E8MLN1KBr5hTml+qW+AniOoHvXltlwtIlUtVafJJ
t5ePF+gOjobm7RIxI+y9+lVoGbYBXte15HZJLhCSRflnl9a7slrlESk+RhqtRHK/
mUPirvSb5Tne5MHHUjXMOXoYUWmI/TEo4tq1bOHKwHoF5N4EGPhayKfMPx11Raes
+le7S2veoU9D6SmT0FMVB20MmTsH5cgd1wWoLZxij+752N6qZNZu6Ko10wFmpJLV
D3IsAU107nqatuuxRFoSHtiJoqV5dkNQU62sa1ok6/F3kheTFBIpgJ2pq2OP9YQl
JybVZtTxnHdRgDw9Uv/5uQhy/RZlRwxKUl4HkO+uKIGwb4bJdR4HUE7tkG2nVlgu
KE2GmqQrXenQLfHRWo/ieq09JKSuM9fQCznaLehMZyiCU8WHi5etW7kEW+RbSx4b
OKIBEUjoSrXfjXG0Tw/BSY/8t77yY3KKkj5fi6Q51XPET7NYi5rEU+YBWEM7oigD
CWznnVDxIYMJjQaaccv4qKWTZld+MZy1hijdOeUuIlB2aEv6quKim+bv677wp+3p
deqiXERVeycuWccya9WTsNqh/XbJk44U8cQ0RBHnB+6otj98LIy1QKMvliOy0A+p
7EeNQAFh+MnpqBFwuu5Lcje158+XNh+rPD4GwpJo2r6Hzl9+LS5ppGoklpD0hoP0
UsWjaB5LaCvUGf2GmJqyvpA2EQYwf1ilB2uOFJeWT7fUZ1+emMjcU6Y/7Acw77Iv
cxwTF0iWXCDTml30TowKyJ+9phO3nkXOD2f7s0XHeRuVQ/KUYhJl7aWMRXfpaf9A
hFos8dUcYviXbssrsv1PZ0ZscQZIlhhmxXSwd6k4kIK6+h0SPPq5e9AyMhix4cQB
Hle4JhrOPVID00pUKM/qTFHw2MRIPRDG28zQRpMfb6UW3Do8at18C4Q8AHNbih3q
fx+pPpEsmWHod8d5ASPrYY67nYLb4I9vqOf8psiFu03aIpDXvEygHzpfPbNEigUP
Db9815vWucP3ZmSvyqeraiwebB6uisiUfB5YLaEmBHYWaWjI4rfMsWE3+lvbKeEG
I1amXuaPqpe6uSj4s7uOiNe28u2GRCUSwUdx35OKWxnWYUWUBSXZbaaCrKhX3HKi
Xj+RGqK/ct9+7SURzkuAS6t0yqQh64jssNlXuxTNpy4PlenKtY7d7q95s53JSkgO
6RYLUrXBDoIisyogrgyaJLXfY73X1rJePIPgYE1YLbLfwyGE4kTv4XsZfu61BcrJ
a/kAG0YqUwYpjenBoikgDMCWSnzIJl+chx4dS1gbAxdVFbx/z3Xtc8TPqyO5RBn2
YdS2l3zqgO3uqY2pY2KcYxOV4+ecX8ORQKS+eoiRf4nxQ/tggn6dTOBP3mlhSrUm
9L/GqLMyJ/prfPIBt75pMHW2RPQEZsYyu3hcGw+V39dSo3TpWbEP6V+E1OaD7L+O
1zUoqdjoa0BenTESuLLEwPWo8Fdi2dBYDjBQT0xVlDrFvIv2fYOU/qqQK9juk0rq
s9BMEReM1BHyH66z3LnqUFXw2qxqBEtLRE0lR2rAufH72eRjM29zogRMzhF0Sug1
48zvMGXUBcRvKNyTVB5Ns9H67PP5pgm9aYuRmBSQWwnLUc+LoqHKWFasxGyHuAls
YCM1CjbXCHVyL8srYZznmMUiE58NScxuM89Dx/CQo7+nj6jVIi9R8T+WYC0z9QVp
CmZYtwlTrJJxSzzx/1e6sCCRqKKFdPqcEieXLf7uZuCMsvitniR28HQOdjSQhcca
SU8aQHghv2cZ6ucLTjHhs5dNbytTvNOm47O1k9A+3+8Gm7b+2r/7NVH73QQJ1o1a
6ILK8xRdCm9xMvOLEarueqnb/xqsPwRzTpOXSLObMMR7oRRUEzG29MJtdrKJ9NXX
LUBlvonPLsTJRuYuzLezwB+ktNKZ5dmpn971AYP3RJni9Hjyi5fPJO5drepXjAuZ
JRTjg6i5NELDatUe1jopAt64FetnSoowAoOMvsLtsWZumqN7Urjb6fiHvUeHwcKR
URbUYGjnNBiq7cD/4SgZVX9gLWjVAy+wzbJ24o3tlMrBtAaCuHDkdxh90flKbuGN
nuGGSKLZg4Vaolvq0GbuRViADUMiSEcpYtlonXn9xIQQa9mPJecUvlbL2pk5fbKL
ZyBEPlvH9Q9PmScXQmphqWCWQ04wMN9wyj5izh1VdTBye+3J9jz6f3vYHR2t4YYr
iadXiob2/k0FuCl3CH0UIxqlI9qtZfac9xjJ1cVj6RAzpdZb/oIo4xPb6IhQ8Zyb
5vUpIVOwgtJcTipnY4PONtwEmtzl8aMFkSfsj0lU1CHz8RTTOXB5Z9nE/cC6Colv
wJVdNWuJgR55BCUETUhbUdw1FYPgY3paziFtiF2+BtqCmP+jzoG1N4IFgXTtXfcM
/HseZcUZBKOvCbYeJzxEcGSZ9hgdCxxlOT9VPsspk+Q7DD1aLc9/vZrdEYDPcMvB
kXUusILzCAlSZ9Aetl6PMYZB/UmurI9Uvx7vvnqShpJQTysDNokwZC6G2AwFBivz
PEuQIF1PpY5FmWjiiTkB58lu+HnfkSkSj52QS+40Ywi17HilzYrUA6U6/bCY98hd
K7Qhm02+47CAqmclWHo6g7UyUnnJtlglVWtuslR02HNapRXcL0nssM8jB+ebugdF
dKOCjKhRl6pi8BpQAbbrZ8O515OP+9/ry3tW7N0qTH3Gwp+j1G2nmkLS4Cxd2Lb/
LIu9Rr55KyM7wye1OENbE3iygRNzQpTAPEMP/zmVEqYKfdr7Vorl2QoE1hzcY5at
iAx3ZMlF5lfDz/1Ldr8VnEAy8J47ArYoxEsBLfK8zC7+YilJoGv2KZCFfGgR/bHT
WKLHUD7MIi5JL8KPjUdTVaUP7KCADLZRHumw3qllKM6W/9UXjTVtp5XQdrpW0WJ0
5A3WXfFeLOhVZd0T2C8Me3+mJk53yZuwTqDqjSKzlH8VyTWmN4pSZ6V4+4wk1929
yz0OiNmiMZgJ0RWV7aOvIDXIzzzLIDtVmn1m70yYpkSfDSo/CuGT68P2AnGIQGgO
ns1csd7ZvV5vTZneBFTl2RrWf8/77h1mH+k+y2cnDUj0mYPn++MLWNSFzcLMcdqh
MBebkLxX6dq2ZD4kw+LJx2dMyU/KsFePnKy6gALkdZkjgCQqd6uEGX6qoPuqs/aR
/HfyPc835WAJvhCrhatzL+MEIOOht5E1Cg6Aq92Uvyd+ufguBN9FU4g6XQKII5+g
EylNUPbHfBVRrjUhvPm6TR4Bffr18fiIfV2ZkoxkFbnr8OKK6+tmnJbNPFo/28/k
GZ6aVhIlZTbgUnLnj+AyZHsnC9qPuB7YNnsUTBbiAXiDYjSnWc2t3ZTm+suaa2a3
TwooDemGOfEe8AxBreoraAMsI/d5lP5HwhwOY55awsbVdHL8F+hUGXgLnzU1Z34p
vlU6iaKXhmsIpCexzlG9dtySZUSBv1lsQ1dsWW8bjsaHK3GXSDkS9WahNmkRGpL6
VKLRD3lHIKxTwSZJREm5i91b4Q2acjKYqT9qmWgEgWg5AvwAgoZjxhD6tE5W97PV
2tPcseNHLT6UTqDpcjO8YG2mJd03+K8cubzd/dawcYN1GaUsVqTXmpmENViex0aJ
/W6VTiGKaoyicGidZR4Iqk2UE2fg+rUDNG79eP3huKuKg5k4vz3KF8M77i768Wzz
YfISHblKwUTQF2DRL/sLH90ftR3tkGQv2VCeaZfL/XfVVc4iPHT5ezo9PPfQ5nH/
bJFPpXLZ8SGyPAwvCjdO9p8qGYLAToVoL7e5pnNLhEGMyN7FfXNfmvUkI3fYKJvW
WJ5iXDwmwlw1dZkrf2zsHEbPNIcvoKp2r0V/g/z8/l0xtGiIcUl79kl+e/scRCmn
agSwXUEqCmfmangOOlmcosJ/VlKMa/3HHN3ngPcVND5/Y6Gxz6z+l3i2X1NfqzT2
SLs8bSJk17Lnfb8OKUc+J7uyro4sDj9xDURfDdNyzdK8LYqdLVxn92upSBYOqLd1
s+rGf69iVHDPcDqP19ZUi+iLYM87QwEjd/rLNCn9TDf9UsBGIoPgd2sVUX5LRuj9
Iw1dB9ZdvHT5eV4fyyh0i5/F3tsJ1UQ8O5Sqels/J6+4CXt96U+kXrxtEzA8C+z/
zFZRnTgHIi7D2/pfMQi21iVftnkdGN23MSXzWObLPthDAMkW1Um7iVlAP32IiE8H
JoDsUUxJiY5KzSJVMICvdD2UOYdrftIK1tud0PHpFa8Hwn1dfkuWThy+EadX52Rp
M0jQf8g0H8kqdHIOHB2V+PZ9hC09hPlEFqZy6NACFRDsndjVJJmhBzocN6Q3Mevk
n65XZd+/Ho5pE0ej8bNyWVjnuC0Ow1stsYDHlHUtHVPXP0NcdWkk+HVIatAWk+8X
Wi8lJZxbCm5pB5HzidMmSZ1WPdzcWsjWWU0se3t6zLIxFc0anEXrrR1mikwqt+Su
g5WlUY4vSuc/ad00Xk9XpCUatQPSWTDVmivxPVCibE28pf6NrM0uxyG48MmAYytb
guP8Wg/fm+6U7PyAM751Ct1uesCwFAYYJWP7I+Yf+yFRyc91Z1N3zkN1E0+PaMBh
McwYnc7yStrfO1PNi8LSk1fULLF8S1rTTlHMjNtxG+u2XlEKF+FGrG8HujjLhefK
ekA6LZlk4R5eqHGRViSjarlPYIl+JBjkq+nvAgnGUui9I88TPPp+v+K/ZH3mZTRn
ICSCbmxiNiIDUYov2boY8sRVVTLM6lulFvU+GuaeXvz83jtLN7ENq5e+JqfynRri
vEs6N5ajPo8y/DULR4hsbJz1oNrMXRXfXNu/B7deKifoE7nMZVyWAub9usdKyZdM
7PnBcan7FUKPk6R0t+SK63wpU6SkhO3wEOnAWKP79w0xLvYjAh+dCzbJicNPd/81
3LM5RLhVA9iWU6vbs5A7Wsh29/8nQT2xDQXcRGMhL9t2ILEVu1rmiM6epWph5bDA
k6AE1nSf8eepx0y5MUgmDxU/FgqPcNJYUGjI3dEp91B2AqTLgTNEuVaUx1iz7lzX
iWvLkRd8LxpAM2sse+sVia1Bmck2xefLOmiFZaRwzQb/r3VfCaDAeYM+ITS8D+aH
hOAZ3YBYX4/bssAYNylFt3a+2FI1mQ68w6+N6iEJAz1Bifhf12YTwazxphlPlwRa
ry12GFaMga05i6HkgoAHJMrPQaOuVttgvhB3QoGDbTywLGshYLbTvxH0/uacnPRp
RCvalZyH5UggrwqjJdafjdPJb7VpiZT8c+BNBpt7TeVzYcs4JNkP1IkfczUTm7KD
//H7GrzA7JFMr4K2zmOIAk8xle0EN2V1lmpCaUinIRwtSQlMx3qthqGBNLGwqw2A
WtO3xp8A/Q8tSZ2+Bol3b+hT5C8qO1UF0HAlpiRMJlZHSfg3jgt5yVJ74DmZrVMm
e2OYWX+neUYW8rO1aMzU8LJH6AI7jejAAB3h7akffeh3i1BCGEL20oXsydeubqqK
h5Oqc9hLKn0RFT9/5s1G2sJP6BLahZODqENjKWgf1tWSHVkUZX2MUhvyBzKkrR/s
g0d7CFliqqA/6qfUvTAZDFwchawS9o5Q780slSpAalOVItSkiS/xZuPbP9PZBZxn
27EcqYHO7LKkzmpt5fBwTw1peEbxb1BW2cIR8EtxgUM7Is3EbVCqhZZRX3DGIOC8
AT8N1VNwMOaNcpIWk7h1BSQO5G8VTjyMjg/FQwCbC/x95v4biDLlGosYgNwjxpoB
VT70MZnLWsPdb8aewr2gB1IE10Lsbl8y4El+cd8v5cnbo7fi0RGggbJry7IHNDXI
WMIqbkE7zjLBhFbyu/tWSpdaULy0l0nrUDPkQV47JDrHe8iZJw9XhNuGu7hVi2iG
bx+pZa4pea0GO0UdbWHARthaGkPdx1KBSvJTQ+hVXvdNFYgRJ7UWT14efI41313g
fYLjPrteuYtf0iVhnVtLSAUFCQt/rogxfk6Byoha8bStHIQWbNQ5q79XbrVCQVAY
uj0gmUH5FGC39fuIbgzb/cm2I7jJeFnBVyScG5WepnKPUKak2lG9RLSBQT7VL7wW
ORemvNDx8/f6Wk8i3YUUfuMPs3dHMqRsjHqzLczREBFCj+5OzfWQ736iIghNMyU7
9nGTlNV2trmFjOqcpPcF343Ztaw3D+wsFNRRxTISnw63YwkhQoFMcnnv+DROpej1
0Nw5Ncpb8ltTNF1Iq9QYxQo7JxY0py+hH1xsXdACvz7ELhkj6WBpeidS7UHvR5hz
NBYvic8uxappYMaguVIq8wyehO231oz+ped827k5vZlS625PmkGj+xjJEPJfjTZV
BSHtXlasmB90fC2aVUdfXWl/t/XMcCJQ+OX4Ktc2czeLfeTacIbnxdi7zsq/rIqH
Qymsb3SMwj/O2GCJ3/RhwhJOfUQ5AD6r52SCBugzgj4zsaAXew0D+KUth5qvhuwU
TkGsv4kwv7019FVleZY0Sgd7ANb68d6umiCBKvLaQZM4NYMDPcjTOwBhC56E3EWH
T4S9xMn+LJYX3zeMCL6kgotA/9P0fYyi5Jdm2TUKeWj4YsWNsYLdWd7amgdatrz9
Zt7W4NiI6rmkvl1Dpdx+Ya4cwnp3adUXpaQj0rHw4tZMfwyzn3wTvvu3wwfAGmLs
hPVHXp5aCODMcv/n3g9FA607Mtl47KSrq58YOS1hF/CfVeVpKqUBqc7J9we9BQ7O
6nKl1I62nwyKVvYfp1yffvA/2UFZQX8fGXMTM1pk37HLl034ahOWK6xzFAWK2W4N
jDqqH5yR8eW9rhFxaFXJwQ2FqjAtFQxTHy413nS/zTpyBUOslEKcFzlcjoLvve2/
F+vdMLX/ip+3KTnfXIxgB1SfTawmQYQrTDYV2TN5wqw4C5bpCzSNA0ASsNtUSCna
bzpyPHErUwoEYftW/e5OSvjDcDs+oj6tZQURluCUO+9tYnA3p0+uuIUZC6YbO5rF
R0U2sxcYq0N1p6QPc64qkwN3acsex9ppyEonURbbI0KirlLIYXlh7HX2F0JLZFL8
649PiLE8CQxRPjtGQzr7yDwCVcSq06Wesz+yg+DzTmVYUP5Xxq3BQm+mN0sd30HQ
lqgWHXM55GpSRZDxNsCfZZjTUsAOS3wVpHaahPJldFADb0x0vkEjAdg98RSaSuui
F6dD8agcws+QnI6oxLOEc/lWQr0k6DcElB+ZHg/g5iJ/2TqjN6asvn1AKditpQIL
Fc/fRZBtU5ya3gurt0po2u2ko6gVGmASTMV9vDRtRFMhu09nMXNgA1Hebq3Uqe7g
KN3JOxOzw0nqbYRYs/mzbETclOniV1Id5CyP56kLGzgxrGEG1WSXS8xvxOkVphTH
TE3HWqyLN8m9OHcA+sQgVxvePs9uY8D1xx7IV+czyl4tS5S0JPtrTmGBVVZ/TNFw
+OOuB9KUJnC05/r4zmz7bOEPMGtrB2wufyeHwVKfpZeRqg7D+nZ9RYg7ThA23+qk
Hr8DqdM9gVF+S7M2ODcvqdHRSMDjJnn4GREBJcEUn5WeraCMmnSQ0tV3ZtO6dz3B
jM23dGv4IDQ7QqO5WOzkT0KsneQcg/9obJj2/y4cTR9OqgNdnQsmRRnvPfB5ud7x
7gdG3haaGAsHSZ4fi8q5r35oOKcy9P9am0emF6Mk2h6d4HWvhGzc1yYcWe+ij+x1
29s+iBL3j6vOPcI2jlnkpl1lG6eBOcrnIqFXPyZVjD+rUUR8hhcbRMFe/fm0tnc7
jSkwhBX+dIjWL7CPLeKuX1yZXoRlJqT8MW/7Me+QQ+MTPyZsFEl5lFQV3OvLytDH
xEr/xNPa4ZgegZsAHdAmqJQ6ViHwcl5YmsssdPCMgyVvXRH5nco54Oen6yt00+Lb
nJksKGqErTdRoVy30AQAolM4wnHclNOoYKL+eaTDECHPjpcd4R2MmkrpdHbOxXp6
lzi48obZAuemVd03fnmmdPmVEA5E7CJIAMxh9hKMcOhBwqy2ORXYLPWDZG2Ru+a9
Q03yfz9Y2QN2AG2y8diPeDaYwDFl5kJrSa1J5iSJtVgMawg5fzUZWgh2RtiwezOL
ByQPn8siinu/Ju1BeCkl2RcT8Pm3QH+HI5OsWuMxQlddKknZfFsTM0Ny7FMm0eBf
XMdVaXWffiimtFu8t/HOkTC+J+HKpvlWJss8p1jQaqdcKI93zWvkGZU66VzxIWtp
1ZxfmHvpAIAstx6yWMSb40hm5dr1KVHW6++qNrKZG/L/DYAgjahXxz9fOAAfhUsf
Ag10nWB7kNRoBg1CCUaxJExbDjFrPKB9hzyokAAx45X/ANa1T5PgvrXTBPA90Jri
3/SPiNrJtT9GKM/yMJc/6oRHNmXDMNIWQw5Pf9STvdVV5FvKyrslqyadNBfE68It
+pEsxenR7igJsdT96blqQum4OZ9ScAAEuQIAcTvZZ/nFS1Y6un1Mp4082OA2z1fS
jXME6KBQSVp5+QAMvOxMm580uHB0kYVjCjHDBp0CdNjxRZbjAPqNS3hEafz4+v8n
SbiBlaQ4Jbd+hazGFtJ+Fvruy2sq28Pc/AQMX+N7BzsTfl2UwF7rQaV+P20RtYaO
+3lnNh3/iV+R8fF/W1NO+5BSzh0cyIlMBysdokX5US4TVtd+CXuqJByK4/MEe8Gn
bx54EsR7vy8dYrEAVsQY3Ejc5i8WLYpmS3aHicJQnoO17NfDVeb8m054jmkZqYDc
JcjgaU+JhprZbyYcrtA4vCM973vgcTVKs+daVzbapeF9T/aePbd3XaJMturobj3a
NcnWpoyYWN2kzDSpoNF3TlSxSlJsHHGmf04opCGSHPeKkYdW+UdYs97r89liOJsd
C5BWg6FWsgpw2wN5dXbcmdXJprL/Wz1gmxUHHd4Ju1Jn2PGhBmXtk+DvOSB8di8/
0A9jE7MlXxGm1Apw58Fd5ZzBqsasuMICNaEmMFG+vq7TTgXMgxE4s6oouZsi8PFU
zIZNfSPZ9FoWjkCMI5wYQxwZF6fpPuRMUDUCAyasY6Hp1XN7hT5O7qGKfWgCyUD4
WImz3oZ/Gxz67D6XPiR5IO7m9kMisFwXDLpeN5qVaxa4VZy68j0UYggP42Dbqx7q
V425h6khdmipMFP99ADot0gG4Zz3I3LWwioOWDsuUXB7D+htfj2nR71FtkUgq/nE
3CxvUVnQqXg1PQvrqeauu/7UabAD4Udan4x2p4UObBQ8UlUerXcKmSkGpr/vnBmI
SRr+4w/PICSCOOVS7/Xqj4YVGBOu3udYxlpdgDB/YVsYjnc6AV4s509DJ/bbYJSG
pWDkb1vpsB7UUPrmB7KJaGhjk02qb3KBkTudx98ahfvNDNcIUQHrrYb+gcQjXuPI
vLRwskEOuIURvUMTH2jyotrAcqnRd01f73KffcJo1QFNTPzAIEyqudc3vLpDp9Cl
DHjLepyALYL1mrXOd3GVjgbprggqB9b2/gg6Ik92Vt/R3Www7hQqqdPP+0pajbC5
3k+ZymbLUlZMAY8Jc+zJ4OpJ8/jM5KCwBFSkdgRCcSUVtWRtXEWi7gogCVYUY1L0
JtQYZQFaQ4Kfjo2XaZ0YeO6atR2B9QGU1vHpgfZtFTAUX95K+3Lr3E0bKiccUxUv
I+Z/ujXk5uSb859fRGviq4D0MJQsMEdAkx9cVj9g3Ih22GH5tob82f+PT4CTJnpe
IVrAH7Z42Opf5Z4KH2J7xTFeisY/c/gJ6yR0TDb0RE6k/u1BjgInh2Np3lfWqLzi
oYYEHwhERpkck+8yEqF5mCFU9llQgDTyhpVX48iF01988i+Q4ROkPS2FREIsnpHr
KlXqnSS9YduBmqE8HgJ/ljLYzOp0zFMMelmqwVZMr4waUlIPFYSudn90lnkH0vxV
SCxTp7T8wh5+Fn7fRo8BitPtjx76VBhwHcjbJa+OZkTODItMIBmHYPxMmajYB0mH
R3beBgGlMsvAnSonTtZ/1Qk4a0ide3CjSy54Z6s4fiickzTXwF7hSZHsjrXGoSyX
OX6QY6+guOIrLcrrhyPrIjMk4PFz0nSs0Mg91pPTpLjt6u8/TffF5EifKIN/fw3W
bXxb5vF2B1K+xaOClt0atdfAS/6ILEYk0ABv75Oj0s4WBb1GEfRLk/MUpq7vQcFZ
QKXtJlf9OLHxJ/GypbK2aLQseSflbKq3f7v1WnO9o4DqGH6BnqymDrgt7jxbPGYc
H9ibuwHwyrfP55/6qOv4zsuwBFNEv2fu62ObZ08FBmZbD/elwhVd7O05tGVAhp5l
qhkbohTQM2X+NsE2sjpf3K4fKz1HMr8tqwW2ZrhRBehUxRrBQcbZ1KnPQnJwt5Q2
sBD+Zcc5d1FWlB3tCwIhRjELPDrv26WQNu+IOEuX5j+AyK/q6Uz8TqMCi2G+E2SX
tSkz4pOzwX64lC8RHPydldZZkPnWy17qI6zQH0JVZfK7zD+PvwG5mJFcVYWD6w0F
biYBuvJm87dSnjOACeV5hAkCa/HsnnI4DmLthu9aJDCMWSCn0xlM1BQGSo6vdvCl
Y0N4bgtNkudI1SlnSQyJ15fi7XwW4htD7+e4okL9MBkRtN3Usevim2CPDsZ511WV
xAH4vASl/eWmHW2Xix5IGspMzJmBxuhSRBLOQo+SxJk8Hi0VodtIh2d6X/bzLVdZ
7JZYwJ6DYJFDgjLj4+vm0cfa6PTIIOjEY2G7OPq+IfgAlyr7ejam5BYqbnQPxK75
YM8Dm+7Q+8h888ttpSgBVUjbCGOJQ3J8/d3FCg7BPPh/+SVRiqy0oBaBbmjxs5DE
37ylUzSCYOlrxoOZSnKWMCI8+XXJ7UyNRTT/Ni71S1PWYXPAx1G1czhQDL0+W4iM
2CqJeL7jagM3qgfsCw5VkSqdiiKnatHOFQzVpzWdmckY4iOcQ5EeAbcBDg7bWDVh
ct8VeA2xuc3c5ZV2eGybYjTcpNKQYzGSV8UpYexjwWbS4tzYt+nejrbaG4CsHB0I
Nwdo9Pcf4MgnxYZC/EWmCyw5+iOKxUkQSHN9edG3soxfkwAzsLxN4523lCBqlCC3
2qCD/BHucNrqTdqESYWPbQXrMWaB7chI+tVa8LeC5XfhLXPXsXgDn1V0Z2cNCuFM
h9kdC1issGqhXoXJG5yCtT2voOUUwotZ7lGhfGQOaYmjHSwmOld2scn2EY5lq7WB
n+NjlLK2lMfC0JXg2AoZpwvpDrFS/PKMnVrPyKSRA+/QbBODzws28oDSK2WEyD97
UATCgcFHj5ReTMjTtLn1W+UDrJEzZkcC+ZV9iQHBW+nDMIdBVExM4F6T3YcLboxM
1ff9m17QDQU/LI0GzjLKH6f+IDnQYCThGDP+zFaJlI+cRIVdFX8ExRyJdnArSIVx
IhLa4yu38OQUTq3WKTTDzO2nAe2NOQ17oKB98On/wr7LXhRBiNfzrJzIg6Suu4cr
88QXoK7dc2dPQnUY8u4wgLAUnkliMXvQosKDmyOcW0cksMFXU9Sd0wSVwDBz3Rpf
uKTe3jAS6zYj1SlfUDcNt/OvD+fTxiyyCf6FPUCDKKpDzW6CDrm1Bbs1DGoXBxqR
1WbEXLRQQ+PS+M5tttoQKeXUZiNivPHxFjGSfBqM3DUJgXx2Z3GUqmd0Gc0d71Zz
yE/TEJItBwGuP43ez8TJlPj7v94d/wlYgsF7PXdqIOSbMw38h6qTWvuHtmGN5wvv
jSaWzjmdb9RqZsExjITfjPxlYUh6kP2P+M/vilBpP4CPoNMMK7uDFtZQ9HPBOtk7
p3zmzBXRjx46rZsfHdBLGdv0a9rhKdodEkSuNyOm5cDYXVNq3Ga7qYP5WBAs81ah
3Zpy4Get37zQTKE8Sb3HDE1a4Wv2wPlEOwYA+XiLOQi3PDkoQ/YX5E5GpAmceXkC
NOls9cPMSx8VXNAysZ3awALmq7HX1UnL1i3bgssjI7ZD4J+eeOw7vdPIyYREWV12
YAPgrJfp2lKlgSlc+wvpkDuI05WTc1piJ+kQhZJUf24hRab/ABvlLAiQOSXKw4C6
MTq69KIwp3nltbndSa/ttNtDxEsZvJrH+jXtJgVNKUui00VxpTeyps3b0FkBfR5l
v30avu+ylQ5YSIWYllhn2Xo1Tey1eq9rJiBVpBmgz7TxCfbHsiAUoJZws7cuiqjv
K02FI5qJDTjAO/x13kRJuoEtdGWHr3MEQbDvRHxfqve0UGo2f1W0aKoFijXxhj7L
fSfUcd474EqybeYFG+5q/VqNoEoodNuPhbPCvedqltZrAB8EBIVB91qBiZrON6hE
VDjmDsw78voUovLhcCdB2kKJ5O06u2t1TjgNvtekw9CbZaKjH4FZmiyBpWasVzp5
LyOE7XNcnlJcewPOpZDYCc1SvqmYpFglRgktSSL/3ooSlw5PWg+ragh8775WGimB
sBs2DiF78pT9rsTgfwOJXNdJ4tpN55cQiW2e2Zat+MicZfKN32EZHUdeUc/I4V/1
DKw+diBgPoxfm7pd9pRXAdMINuHhdZt2WUZBa0HviNGBPfOQtzHAhKWb5bYkyOeH
S1SuCeQ3vDbgjM1tmTzixsk9tu0tU90XQpoX19i/MHkTvvv5QsrcyT/KPw4QERB0
4mr33qxK3LzhH6UBawVEcR+NySuDWfuj9xyE4Tgd/F+lt49ZpgRGv/jtSr2IAZ3Q
bX2sBxLEHFoU8mHMtB/xkWJZjF0dHtT0E9X7RX6ruo4iIVjv7M3/P4S4UKweuaVa
DvAU/VgXC/RGRrrZBYVgdJdcv39bL9bCCXa9hUVPxd3v+9HFWWe+ZrYVWlUN0Cy0
txciuZ2bGTvyVb1jtq1rOUuzhovWVEzUXC/XGi1+5EUd1GN1cWBdQderH88FA+Uy
gi0/t1714p7aMQDEAk1Svs62cz24ouI4zJZZUQK7aTC1CiULTFRF7sTfkrAm06tg
A5tmKuHprSsoMnjBad+JYyiJm63Cc+R4N8eUOsp53zmyC3lXIYByKhUjlrHYawtu
CnsMwvAz7Qwe0w1S7ZFG/YNVfRu8iaJhitvd5bY1q8zuJg7vg50tGgM7lD+gYzOf
3xJNjX3/7Nk85HrLRX+YZLZAPkRj6yR8bzyMy8SHcwe6V2rJxh8mhA4pIQ1A7Mcl
b/2gjjxbnDxhlv4tYeI/KGhDOMU9JGqXcqZVs0Uv9tXJ6hrg8XAqjE7MdYHn/2c5
y1DJUQnc2Ti5lPIICQTmIfZ4bqXQSl3vqekdKVS9FXACay8Netsta6lzG1nTSd6U
MWhHjDjo44ZRd7VgsStWw1fVoVpZkv+QbEfKzf5B7rtV+gwbvr8nwzslwiWB5bZd
36YMCUmLZuTMNoG8gAJdltxuL8OPg3rm4bQJRIo3sxALnPuMLVO8tqmkPhX8UCzc
yrEs4eWLa/CnrbkUVevU3rhikY70rOtMfcV+HfqTQbCuF9XR1yPGMjbeX1v6KvHo
IW5vnvC1COoqgcxloUEtl8SO+7mhuZlsDTppoRLm3IXtcsMlI70F8DGSJlURTChP
lb1DJnIx6Lq7oIn+3QL3E5WxKNfXsZNRSow+Tk4mLPpghYpSEIxJbzyDNSsM7CAp
tQT2miNO0liB49UxD/FYllxrt3EOoFhaQOYvUkLghR/iq7UMnimbH/3QPQF+Ni51
QiigaB8BOwXH5EizwDYKvyzcaqFXvubob95836nqGgdNwTaO3eZL8m6SVo2UdL6Q
f8JAw5z9j4WGUgTAImJRq1b+tS7sXIsVDt2A7C/dOox4vTrOfwQpCiGeNF2L9823
uG9rGBVXiXGaJgmj9zOJxB5jqd0DR+UkeJU6XrhE9wuxdoMIo0D0grCsByf9s+JT
BDtifMBOktXKH2Ay4PKxb3w2phL5tEaREms7X1+SJkl9UFOEJoY5NPbR0+JpYFiM
tRg0QAWk6WoC153gxTbUxhJuuc7amZboQmlFDoqXLiw+g5pKJlTP4HpMSkzKZlLD
3Moeg+R1VDE5cEKneHHC4CG9sZn+m8KjBlha2X8MK1kmdHyNp5Q98DGjFeqy4Gh7
zGtuAstZeiaSrRMgSm4Y8NYMTxe0oEyH8XJsMxkQgRNfuBOqQcqfxvj+/2HA5bpN
x3m40u6v0OOs2yfRvpMlH0VqAGZuKbUJdLC8qWGCxAEcyeKSy9lQwF2jSmqNy/GQ
Q3xeOjBq4XD/r9Gb4iVj6hqLouZWQpV3gIg7tG7Y3dZ30x0GqkjywccUJ+bGNzj7
Zbl8Pg65524veEj2t6cuSI3EpBhXv5iFABW+UkofrOWGDXthxw4Sc40BGy8G426x
+jv3FlSlgH/+1neOJsJnGam60+E69EGTqkDKBjjF80xZOLsgyHR09TDrZlgR6uq5
jUtCnWPKkfFmp60o3cw0lC99GMAx9hz+WmeJBKCgZ621EvCM9Aijn4EfPVYU0bOS
jXwL1FpE9DXHqjTykbMD+GpmQbbfu02v9ZYgnSMGs8h4EdxtXHwb30pHl99BhYLm
uEAKZrssNAjdJDqSLUcPEh4tBBK5yzh90Idmh4xHmeaI0Ygyt8rcFMYSEHsCBgHt
r/Zm2Nynl7bGr/biuvEOTNMHG5ERIMUVTgIWh6oy7rm+q0fKobqZOOasJaZH5afk
xqo4W2iVIwefHkJZUPpbMxaD/WCyvYQtdmIIke9RgpHNudyUXPTnTo4qqvXFMTY+
sfKKrBtx9O8166HfsnW2o2dIbkQ1cKIqz20FaKhEkFHRlnKepDa+EFC1j9AZTNi8
K2m0hGEFkv95Y10012H5lkE3sZGxrWeB5Am9UmgF7Tf1XLjCXELi+yThyT11BHrI
TPVqVdlcAk4EUhfCscZFvukScex+O8iip3+HPSVJ43Mnc3DX1OvbnwSQgA57PaHy
7vM3kNUe5FkDQPIy9/K1DtG1DeKOPq9c/aIeoferF8Y8cR5DloxLLsX1EYzieavH
DH2PKPKDC3w/P1aoPivWVCB5m0ggd5FaEw2CtoOVuaFOHtfOUJiKAdC26wSPnKoj
O420DRnJqIZNN/sxjVWwOk0vyg5H2UT+2omD0MMb6mK2ZknrpeoMWUG66qwb4/Cj
1uQBQQIc6yBu+0dSEAAufYcohaklOMoDHTSO9/0HYPs3gpCYlXUjVAahWn3oEz5H
DUJvHeeoLLDASjxLE7bV+MUQ1sIJ8i8Zab3rl0EfToIOshz2JZ/zoH4p+l2NNCms
ymdxx68y28HtrfTXtqC6I7OehuajI+DqCoz5J+yntL9pa5+I8AXu2FnUYdYq45mk
6eaFLbPpum6Ew3pJE9K5puf4cY8I2TO6yqdanBKUOKCA1hCw6pCELJGZjrN4qKzH
2neMG4MuHATXQvvURSct5BwrZg5rMKPj2SA+WiD/r3BYxBE85z+Inu5rQqlAefo5
fPjqRvydPs/0Qxh7HYQr9viLstCivoeyR2yMHPYMfVjBIYFeMbRwCRIvM7e7VyR5
uBFHk5gdxAx6e+yHKsyKHxnsnBRws/5y/tkFKLzADEVJkP/mRObxGadYQFdzDfCq
z2EOYYPiXEj9atqNw3aS+L5YuiCzZBwLqnKq855so/wPqUNEcl0BhbdvbgNqusJm
SGgD+I9gW7QSDEu+04TCnf8w6V7CquT8EM6yJogv22DNJDurXDU4tL327ApCEMa3
smCQMzokBJ33LUhJJTySNmErYjJ06nufJsnhNZcF0kocdjYhdamWEUkYvsUEZQM4
QeqgkS3SCaV/0r/+jQU4yngZ3bCjyofW5mteXCj1XhNLUdFJE54WU1rxEd7C6lKa
N8CSZBC38VIPhv6ncsMO6OY3WFnTfDThyiThrOf0oibOmIV3e8pkvA0FDnQjHMqB
VAxoW/ZYijTQwpG5vLl2AneqVz41EWDlDJiumaPlmM2HJ8peMaeUxN/MPdr3x5Ww
gCdWh0pW4f9Q4FWqfcFej7cHyFbH1d5LBdxnxi7LyGAxbGSaDE9EDkCokQhJkcIf
KwX6KGoeIG4AA81pYgruGVYhFs+PU2ZiMa4dUbrAywZLMiVP1zfQ0frDLncGGVBa
6zpMqiIutMR3sKWsUC2soMp+PSChA0tVanao7HshZ1IRnjkT1aufpLVD1mjEQYJ+
fYvn5VlWpPX+2oK4TPRBKY/bCR5PmMayI/ZZDFHvWXUd5olB6o+inQan25FCnqwn
b4uBqkvIZ9RDISzRdtPUx9T+Gd2QF9z1F2xhSzNzGwAKBjHCzaBO1JwaSko+uoij
5+laJ0Wd5wKB0ljWxR+hxT/1O0gEU08a8ar1RvFKIfD6yl1z3Rs+L+gQtEBwt63p
YslCbxPqv7CLzK+xoXDlGZt0n/TyKAZwaETFDmZ/19kCM4SclXKDgtzmEiAqF+ro
Jy72aS2/JQYZVid26rBjqjp6t/eoKKrBam9lSb3U1+dS11nGFDh+xqnafdogSZTA
jng9m+DyEmN/U4lcWGGwBd8cVeJ/4WnAQtJ6qpI2j0GYYmoO1gyrdAr8+KoKbc9p
1SZg9m/FQmvTV9GGveFbwNfCnQg0xmaMMUPp4KgQOHplbiOwP65BWpfVZfnSk0LY
FJRdlVk7HdvO2HdX9Wz9YPCkBZDOSo4QjwJSCL5pggubB6WNAopl+hJh89pIsVM2
KGbmXy9Rn5+PImQA4t/yeQ79xvfD2AWXOSeKRNke/kcVFc33sAibZYVCRL02JVkP
Ulgf+pe2PO48Z+CVZCZPFYTdwbpoHgwepADu8hHgssP2Yyh3AoVLWH2Bqi7k59jm
zAc6qOD5OKFwC+b0EAZmkcHThLDVukyaNXP3giW0MNXMoVfFjmPJAZh7ShNms17d
clg+Q0p+vXTTNI4KwR1rN35qJVCRx7Vk7LcSqmsRlyGDZbVZiEo0npfgsh0emYwZ
cq+Z9oH4r/qpt34QIfP8IQA3cLtUlHaCyXsNEb7SbtDOlfRh658pU31OSkveZkOl
9MNMKui6JkbFCM7jadji2Q1j0AKWgfjEQn6ZCpMDAXBaIxAFDbmf3bCdoTLoJMic
2DmBomioMZMtShxGNVoB3iJ2atzoxJ9vhUD0y1Z68l1Y7lYDM8wgn/Rwwc4jAMUx
8Li1t3xAP5YL8/u5O9I4mjL6Gn7ViogI6pPUpyEC6kSxFxHWvPZtzykia3TJJkl5
TvrB1JUsq7nma6PziXz3HqlxyxfkLVNhcaPBr9t/BEdp6YRlE4VYQjfV+1/SG/AP
iSRh7e9F7/PixWwmatVmlQc2kI+OkJiGTjkO3m0ovDJZ5HlSgRWmLfLE6EVLBapl
FF+PAW5R8Hlg2bnnblafpthoESLAuVqQ27cPNt7kdkjNkTX3CN1R28y5avQ+4SQu
qWJ8kBaDqqUZ9nVcbLhOnVjn41LkRFN6ZmpDv8xWvJa0fHoXCzHZbasPXWMcQpb9
rwR82lEyz8suwxFnEYgyENPI5pjnXhIu6SO45DNGZpwLWjRCI+AQhY/EdnJR/BWZ
8Op+QIUUqxHNSbQm+YXg6fnOG002OsupBeYurxPzofB1IeepRGDTNfX5VghumblK
4qFIwTkBdBtZFIU2DWIqMQOKkdL6dhiYWihLjBEPE+bP+EfJmaPeB5er1NXHM1wp
1y1CVxIIDJkSDpDZMccUKKBl4RJSNluSTVEEr9t4Vjvh8GljAMqg2JKOVCHNuzVp
NSEiNTobS0SKRwT34tqnCv/GyL+A9ELo0QRA5R2wnS1C5JlqyeSRf6LS4TOtL7Kf
KvjARTTy70v3yqLZ8fKoBAIiX7d/zgW/1qNLs/VP8bofohEiw6S9IWubBSn4J193
jd5fFH7wVtziQLZ8s0JTgNDhYKbz+6mHf8Up9crh9AbYb+GdlfED43SDLXVafELe
FhpkdHfAAVEfT1CZLL5dbFiEcVX1/s2DO4eAlC3NRbAKg6L9NBqevHOYYvp+S3Y7
udgAZYy+6LryIEENy90vjiZW0e95kYxcB5KN0aT2TfVCeHky3tjiFTnaTcfDAgPY
zhoZzuC9FykRfeay94jKow8LypHR4PvJWwbJaGaOjWWLbsOCwNaxKOgnQrbpbL1V
Gj7ctTzmtPnPsLrkRcOW84PTegmUu1CGKLAWKxiC46ctyK4zs+i8jMoyvUcpKXk9
EQh6UIBUCny5CMsQms+28k8Ld/6cxA58Yl01RhHFyFsm8SYERXadLT9ZXQHcb57z
23voCfnEN0hAGxFJgdLzkCoakS+UJ+2PgjN6sRsir0tFUBUZ7DzLtDBIgqv2d+Ya
9bw+CfKWEPZncqvVObZd9NcFRjNFyAdRuW/xrQJoLm47SfdaoS7PUE6olKj+ff7l
zsSfM2HR7Z0CQP05ASbZJggb+36h/fBpaUCieru50fT6N9LU5eIl7aIJ2sX2oYKQ
+1kvCU55nigwzJKu14A4TQU7+ePDHfxNJ8b1rgA6SyIT+yFk2i3gsSZDKb1KYsRf
JewKcYQ8IapjHDQP9jPvSx7HJuKt19tl5PY75fRG1GZ58psHJoHURthvFXJBKHTf
QJCNFY/xOKz4TAOLAWSxR5wA/9eAIp9GQV7kTSSCzh69iQaviyn/Ha8JwyAAPXSh
WMVyVDdYx+ZkitgQRhji/Kj3KkN+X+JgWOKHNLcmqoNJ3Hxlm7K5UGpvgLCgoryM
i6w3025cqedsfnOzwQpi4a5Z/0r5eDhS0/8NkWYTL9zY4HyA6kH4P9IML8hIrtWQ
x1FS7uXYVj7NFz6mYuEhZuPtrPRz39+k6WpR0S4kqqYGVmd/WjzlB+YDTkvKGhI0
vRHF1xr6UDH6Qr4n3zHWq7Pf/DaoXw9v6LWevS2JXedo3p3j6rb0heQ7aVDDTEqo
dlmvdvGD9vMeLdnkbKROqnwWcsuj2cjOIOEl4uhOhheCTaQpAvMLqv0aQb4Uv6MU
W9BONsXZzC8qacnsabbbrW1lK1SJe+D9YTu4yQ2QDxVEr48OCrcofCvToZOFEESr
2L2X72Z3GtSczzDfd/S8KGjE3VxXK7L42FkiwY6YGFkXF7d1t9rEw+/w+03+rPda
1TQs7/1XTkv122zOFyuuXcj3bCtbBSnANNoFFXhQ1lfuofPu/xtZYTJFCzxHoWXT
7BP6uhY7dmlaxg0Kvem5ZOThSD73BdhFRtjcmReke5DIcvCfpFwoGZWhVDHXMOVx
STgirD5gwyrkHW5NR6Uinn+r1/LoFAZH4jLz3WZOD+CmwuYcxWW1OpW1eaMa9l0w
y4gvn71OazRpU8wMtff+gVUUCV4uUgPi3vNc/BblKoykCPUzCWCdg7lF+7GKUtwp
2XTu9dUalS9RJ83jF9qbgTXbz87UqoWxJ8LXzmEF5DW/csceNrPpJkl/y7ZHqlXR
CI3Pzn6kcn3Ce+VlySN36+cFpOAnYXK6CC/Nbgbp9xkHet2lO7MBaBGMb2ch180F
SONDzobtVa1GAvHNAc8n5hi9ZMeP5Zw0K6khm25C6ynglnCJKKNepEeIbWg07tCf
vneJs6Fxe4ud+nYJ+jZJpJ5AEI1Cl4AhOOdJ1kuH5Dqin8iDOcBCEVpUDaFg1/VU
5ESXiDFTWlEHVh5BUkZrTcXd4N9FLPntX3A1fpRtfEddHDQ9I3VlKhWE0bGgWxjK
lNA4K7lYHfAlU/bCox1ab93/iau9FUqKKvGQeMsfa2XgZG9ceWdh8tFfvlcHVmAF
z/mhWl4pqpY0VH3kuAe6Rjf7e2SZs4l50qVzRC4R9UMlcJxXxzE6biDDINC6M/Pd
gPryBUwpVHxurs5G4LCOmIQiw+aM2fOS35GjYKjkruGD7hKvKTfltxHkV7sa/M+6
yTM+tTs62+UQagUvKhtOhoJ2IJxkeEUi4assYC831/TiLx5qT0CX8nKcEiOohLe1
LPDlNhhfspDSbPqFOLGK5wpJw/1TSPbZ/n6VmoD4113vxy8e6jfzJE/eIafjNpF7
E7oNIMro2wk2EbXHBGkyv7qcfVkfg7s+hLcWJ7/6nC3F63VhPBhxstTL75armzrw
pnfzknJnw2luRPzj/Vb+Lpv/oKTLskRutDGvBNQ/U755vK0m5lDrsV9iaIJo3VLU
Mg6imZPR6CfF6cRhEcg8H39Cd0AkRKLDGR4jsl9FasTd6So/rpuo+HNcPX55UhL1
L2rc9u/b2QNUO+0bEC2zmtNjus6y1SMx9pBmJio8WaEt2d6dle/4CYi2vdRc4lJo
xAyFxW9OHgnvqbJtB/HpKVxfjeDKgdeM8vv2yN9KN6otcJ4cKJsflTMtOuCGlN70
UqGwppIjgDqTKK+Ft0k4CLrLnb+V7lc7MXyfVY86EVoI+rOibHJjROmBGWwmn5UE
IjdIBdUkpYPLIzyRNHKCT81LbcMdnlrpYukSCJgTWzuiYegjXh3HGm/Y2QCqZdwY
0MDOX6jQqBQLTLAcYJu9I6X5Zx9PUIgy0AZz80a7vtv6+NMv01aF/gcj6Seftg6d
Cch66zgicKXaIbDXbcojbeXWqN0xUCl44psm3iKBZf64uNnQR5mXGm0DYu4SKSHC
v1f/6jDNQQ4ghlLJl0UqFlR9Z1BiUKkZ5e3puZ5KU4Ik7eJt294A3kGSW+1dsoAU
DygmvrpLMUaBeRi1LdWSjPUzEQTbQEt6+/Euux1OKcCHYonf6tL9ZoAlPXzWGa6V
azjagR/5DlQ/K1JgNpyfdTI4o7peICdEiTK0ISJCmzCpxwSCHz7gbXjlKSH7IgSJ
sB50pAsLEqiCqUJmfS8e08YGdzS/mcFgA/mykYX3BpMMHJje8IBz75xvhOpzfM4W
6HniDx9POi3VBc4FrpijGg6ktNeiuNL4+fCjDzzCm/Wvb2vLGryJpQiXPo+pvo2S
FPjq8GcEKBZs9swrwpfY9ZNMZbKjrtzTsVUUrcqty2ToQIa9IEfXt3oU46yhE9K2
Gmbd9mZjIb05aklCbzm6cE0E9/DuqKIaJ7FKYr29qv3UBtSVbATVNul2H4aW7nhZ
7JB1v3yTtfxxuKaONQQ12/FMLSww4j2Tj1KhrY5J44B3xGO9ffkJsZAQnvGcHPQb
xEiLluka7oJLmynb8lI6HMdqRIdt/lgBbmNOVHSNqX3PjA9h2w2uo7tHNWiO3eQI
7/XleNphQfhUcfNnDCXmsfartkd7V9iqxEU6ycwB51khvvssNgnwpDe8wNcFmEUc
e4V4cK7i0qOa6/m62lOF1S/Dy/jLYx/HGZe0BJGRVS5tHkhP6oHau/Fd968VRT5G
tXhU8K58TM32LCS1kGlreUQX9sWumV4tgXWjs5xxEFySwMoMIuPol/rJ+G1YccuO
k2eow82wzOvrLFqbNPCyAeKJKf+m0bQtDlbeouD/0T4QE3zuRB9XP2Vmcn+woU4M
eg001qhr2y55y9Le1aYGM5rCDMLrBPBdcomQt98Q1nopvmi+WlyFIay5H1EPsmgy
Mdvh7lxM00cf2Qrb1+UvTksWk31ZtVvr4JBc3K1eM+4e2d8S64jEQux0mlpH2V8K
yyPn9EwKJizoTedOUqXOlptDmnKFmZA8vQF1qtTINWgMgD14qxz5TvuMXrWZ8wnW
JbA87DKP4j6aeTjCPp/tDv8p5BasA4ZlL56x17Gfv/nSxxMKofUMstuq30rmNsaf
3R0e/Yjp4B5g/N1dLIL/z73gBiFkJ5j4JNIfsJYcbAD8FLcBa6h/amHUF1sFXjA7
JE/+A6gFaFKeYnehNipS4VToKj1f3tT0gz2nxJPdnC72m17QQ2HagDFUcceXR2th
c/Cr2UwJQ+PB53qLmD69yoGfKwqQSakYRoRjVjax01B7bmP5cS0/pevX9d6biBbg
HhNcRYh+YedmiQ60XtjYC/NKtIVLRb80gIQaaycpF23TkSyvyPmwSV1MLnkHHoMa
ntgVD5XvEPmyEOGR1hPrBRvDzlN2NQhxSE//iV6xWzJ7OOvLfaWld5Sda5LSuHo+
ao/DeNYa/PS1l10cqdoFdEkg7Pa03h0af/heFZn17C8oC+EkF6TdviBNgcbr64Wi
xJe9ZTEKEkgGpXx8d1FMD3d+UIuRxRiq+I6jbQw8CBp7iCnr0OrKifFWMhzrpI+c
k7EWQ7i+mmAj/6yNLFiUKjbzb5Cy2N2IDxhNWLiDpZwzxL8GLYP3TGMGmumS0QrT
KXowIrcraESydM3JJOe6BTSW1pwsbD/pfQNkIoKTztNunFJZ/4TFKkyq6DJ5e6zq
gtq6xHvh/n98R/WACapPbadYZXH3XeSwoSsXAS17kUs8mKlgHkO2DAEeVfm85du2
C26V0kpWFQ4qD0arsd4x3k9c/mjljvWQv/iyrizw3rUhf8hMxImCek0TaYr1vtCM
K8DH4hP4AX5uc3U4rtMBLKE55skPggj6Uh6+jPOxJZlrhbML+j5j22O4eHCdNsJH
cxB/TWvIYy6hdUH9spLDo0u11fShmWRQfWf3JiUKfMXQWvd5YnFXf0e7z7bJCDF1
DGWOR2c5ei2gKi+ughbzyTePsET2Q0lPgywIKie3LfXxYdKXlQ5DPbfok923RDGk
0I9lsWFAybfgqt/QVxa7duKRrAIEVqLz91rmrtbhHMPFK7TNrIWLyM0QjHhDgxqT
az4SsMSODhe0U2kLvzwokKAStRhutSlg4cdb1GQffhl1DNpKWYaNiXfm6LdzZWaF
3pLZ+7lUcEfRtnyvCXlggUONOeJvxTisu4P1dm5HnyiNYSR/i9wJJoie6E5OAFt2
zq90Qsy44WxRqXjKd5AcX4iZHpijtroGyDHRRygFQQ3dT5ycJAfJsulVnuWnVXcP
vis9NBeq8VZYKODwv/5I5jrpLQIwdYMhmuNWqWyFKahFMVXLOwbgfLvRF9C34ciR
g5udf8zSpFvNRtzEE2MMF2b4KtXwlb1V3CM51JU90p++ZbnKVS/iRLOwbzuZrsuE
+nK0aUdZ3vz4ncF7lsKLkD1Gf3GGNYJVm4AW7E0TZuR3QC44LKjbXzKJWOcf43Ky
1UVCC+LtFPTqiv+xNXqaqJXsceIec0Ap65j9kn7meg8OPtDJuW/24VO+ia3IxhcQ
B8Va4yzap42K0OeGD9o6zJ3hKEf7E3/l1Tom7YMigVpw/DdUdl/Wq6+YTdLzJsFu
g193Dfy4riSgtW88sYJ9lbBZF1wkQ8IcROUmNF6hDTNxwZIKMvMKAqrGS3uzHlUJ
ybSwXStf02KCU96o0HWndWOfw3zlDGYL0v0YUPS9iGMWWNvI3N6u/Yobra2xVU9y
pbni/v5SIlbYwXj8778ypa2c0u91X9s75m2n3y9tthfOdgOmsip98Pn8ThDpGnqh
VDBwir4YKd7I6tqU9KKhf0t1qp5t0vvTMvUrUFdB7+PBrDZx9uOfhcAjM/zsUUUJ
1+oGEgz5Bk1S4BPzZtOP/n938niyYP1QRAFVmZuDS2Yzqvgl19GkX5dKaUPARst5
O0WArGAObPm1vp5twTDSOySez6Ae8XdLSbgKR1sK7j+a4DBUZ+RI5hRsy5UstX/f
gEFUWNGHzNxEpTxSlgilPQoTTUP6nQw4flHkIUK9FjvrY0+c8xnInVWWGnaFQRhh
UI4TrQYVhkHUTwp+1M5tkghEDitT63jj5awsqckSWf7DV6/g/jFMfygU67QS+YNR
tMFjAdGJoaKuSbTybS9q1Tw3jh2w17rEebsUKti5cAWbv7bHxFbklUEK2QkCNJ3X
dI63+XmM38D5n0OMD7X4YQPVwsqr2D1eAmRXfwwsEQONH3mzUGdcy5O36+KrnNRS
Ij98MAUvBbjwPb7wQ8EpTtYlcFTkVvggRLGxqFQGwKSBhMZhlS0Gf3GB1CxxPT56
sT9Q2o+461DD5ir0UKtmlgUXTNcatv8Mv911DDSphvItSOXyDx+zxzYk2LXQcYHE
wbChA39LV6koxT77+s8hTDg4gi1GCF98BDodkp+Df9gZxFG0fUub0XBxPi9FcDZ5
ae0XadV5JqV0DpXRajo90FZaHb//gSN8+FOrLtamDR7JuKV4z3Y3gIDUas3CwXl3
BnD5kq18fD8a9VoAJAkWQXWP2b+8zWrqEbfYiVWZc+bbyP4oZx56wiEmG7a6TWrn
pZIBTe6Xq1RHuTOdyD/gaU0t2JyCbGnlkmB6nl9uWhosOQmgMwDgQ8+O8znIoSOz
rrBYDxTq1kiCBfJUNAEtDVOT2fYkPzH25G0AK9Nybiw6I7qrhldUTISX+q9bAzoO
KXWiDyibuqRffUSK7qmQLFxJ16mdRzIF/pxn7IMiVLbEhTmciILJGNypCSNEXbCI
PQpeB+CFTdGToW0PneEXDzQwzmiJq5aSFAFqXTsWudw=
`pragma protect end_protected
