// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
XgvY8X6TqDJWn+Cx78iWgge8LD0bVDMl+aW3r3prd934DWGFo1UreCtDpOXJ
w5U4agZd1nEg1I7k00wmSdWLGHpF24EhVFN96j0c2Zvm3p11fB6gmyoaWnC/
0G4rEzj/iYingFEqrYFW1IrwkfNAn5MU1npLmJWxVH0YZGQ9ip+KqZfPZtZV
L/n7qpKd0oDW5eCjUEPGsHVS3QOL/wAqS6jlmhrGwpY6KArUK0kRit+ReQ2f
FchQzx/bwIicExedgmV+CIR3Qn6ZKtySxsBZyw/wCu3lUCUmmNb1PJcyoWRU
T32Smzolfbw7+TEub9Y/u/09oPZZZdoyLa1SQ1DNMQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
mjo8INP6st2f5c6Sbezm5xPI5Q4zzgpaSIpTPcEYgA9ToUJaZj8BcDDZ9ttF
zsLC39eUM2gQBTc2SqXD67MCOahSwDz3nc5YfWcI7UXUkwKB/y0MDcDpB9qU
O3kLxoNXK23mCEEzLpc3W3x+QjXGQYhlHz1bcHLHFYTW77M0JTlAYKLUQdog
CPTfCGBDGAmvIrscYmnSr+51rRlFMr5uZ0IOd4ZvFSf3uSEf4AzWT9ebMktS
kTLPlXj0lk8mc9KMtsKUgU9Tw6zAtMMs6jbrkeJZmzf6lnhakD4KUCkyU80K
sIdSmUx3pJzlok1vnroNPXPbLYFzfVSaiPz+SvuzjQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
JB+epgiiazcIDKBCnjH2hBDXzB+gRpZmFyuq09m+gqkSaoge6iMyvWZhdozL
r1GtvAiCPvdxOH46hH0/ygLTG8NIvvO03h0OClG5BwUu5jsJmn9bVhl+qQnq
4hmIf7Sphko7mme1KLunl4YQL9sJejnE/1A22ZMgvGj86AEO4wu7sotpS4IF
A9KCf9viUNz7VJvCTimVskWI5MUB+JAdg0OA06xu27eGd0ikXIQquMHF6i2O
kQNb4tNY8XupvB0Wa9rGx9G8W9PC0B1HfJOeYUatGJO3vGREBJOmuRjxTOqZ
W4I1G8mVbpRt0QQOk+WUyUZ3iDGkwhZ9m8kKzbcTdw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
PEibmolh8/B9zB2pBszgGNY90HgVhklbL/erhVZ9Vtu6ALy2xWw95eAutT9X
YvMC329bQS6RLwOe9bR6Hn1nU/XtcUyzBF/3hul8D0ADEzBr1Aw8bjK/OfEp
EtaVTR5ZwIMGOgfWIYQGYGbXl6tdrNC5wEADW1C+3ix+M4knuxc=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
ZU62UsxBZCK+iyEwFmCRzqMYnJ+J7wIcQA7zFfoAxa+AOfaotRu6d2g/Z6DM
xoWYuH3N50+e4eCFWm2JMrChgEQwarb/85c3qPguW7h+D1groOpIUMkB0w1u
7daVmVH/lbeGxBYLUw0K6v4iVptdybb3WIBRiebW5KEtC2SmyrOYv4Jvprog
zlLW1deCGDMkgLGhSu3GCKDqmR8eskwOR3fy0ZmmtzTgE1XW5SoSI05UyG4r
vJv+qKZW1EMXs53GOyYiVexhFMdweEW/rh1jXtUGiGB3RcLd1bXabmI52rsG
easHZhVp8IhGgrFp93Xi6yWoPwT3ezJw6iHEpFUw46QOK88ME0suZGidYC9K
Av4IfTYTQGShHg2ZdF1ijsIkel/Cpb2av4SDKrG96T33wmyHFYnugE6/DWf8
hKl5sh0oHMIVEQVNdx5ecbjDpgCesxjAaD/4qiTe8lv4VH/7+MDDjomC+YP4
7s8zNlJ7/fPDOBE8NkadU/UhJrFpb9jm


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
OD2NiWgHC5uJKn8iI/0WGZ34AcNpafCIpuRxtZRn+8gn+Z0Vu6n4Jr6NnAld
eWSNPgO3rq/k6l6Uz1FMJ2EDYvpRdbp8LWogZvqSbkRh1Vg0+HuU5TOyx6lX
2XRFHriAgacS26VHnuwy68Wzkc5WWV3IDDm0849tur8HwQIAtYs=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
i1UFYr4Am5vm7drF3tBS/BZSlW4BEjlbhJXAWP4SRpdB4xREBUFk+OFQZUE4
zgzMUVtXz2it/qjLqLVsY/mKIo8nSprXyRKKvQMKt7XJfU2Fuda3Hn6ehoW7
OHqzpgwn6DSt9F09m8Vn3fE2aNkrxeOw8plCcfYvI0cMZyj+8go=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 7936)
`pragma protect data_block
T1z4TjhDBsw4m8zVj5l2Mp26W/GZg3Cgchf6gu+39+7lxn/2bbqO5o5WqHqq
wL7BKuxBRBrTnx3EbaBIJrQ6B/jQbAi7Kx968d/CNzQaNnjwcMYwo21yx3S0
nyyHXnqfKEfj41ivLWTU+ZdAvu3deWs34EeQjiV9CUzjTnZZ8CCqRJnAmGKs
9DzytxOaz/dU2H58bunSLy9bJx3wpG/VQBAoj021TxFinfxduXDI7ICleFBw
Iy3tYAT7LbD9gr0czYNBmxAimgeLYWuGvqt+SzVrU59krxRFwYMYnYyBOMDL
05nK90EkHiOnSpo7TKD8HkZgmzChmshAHXBPmgjdXG1+HpQcK0ptlZ790X+J
Va8JUZLzo6Ffmdsf3opcFXmm3Kz1+p10nn129468GU2A80UA1wNgHyPX+oMQ
JZ7DJ1XASo0zJ32i0mzAHNKAwZCcWEdO0DpSOc4oX4eFBhko2wX9mZKJb6pH
I/QiYg27nDGkyv9mS0B9+EDQ+mHpHebho9Rzfd3MfX0idaIIFhpHXmhm3MDK
mq1LEZUK8U2LzpL/lfq3JizkbKBHc58P/qH+Ad4trt62EfGfnjxtwtMYu3b/
V5cAutdZTtMaaz8lJUqodpU9VkEUaaQUlY6TLOh2gll9MHsF/pAHkSgN55jG
3ZltWQJssQjGmvG2ILha0nUuEjyNwrj0bq1avG0Lb1OFAlwKVn/d5oBSQGye
67yNqz+h4+h81crULBbtk0xF45DRXPNT+G/8BGVIIiRmfQEOYvh/GekE1lqg
npOVrOsBtP3l3d9+MnCRNh0FPV1x0ItlM+vaRBaJeW1zP+HzXjWaDe8SXvJk
06UUcSVYsCkQwX485THEK2BPBYUXCzTxponxGpqkSIue9wHiqFqlT2hvkrNN
+nK5Nu+T3cIYeHaCDSSrzMki2LASISF8duHppaaKcNT4QJTWRS+2APfGlwh0
7QFmranHfvKpD8MPFLUns05E8im9QWpHrZNBGb34ZS6eGKlIQnaiPPe0pysY
BGFLIH7sKsfId5tBguAc69SRW98Y9qj6at+WwkrNxdkojIonVnNLxlL241TV
5u+iOPp+olNJuyR5mJPNAbWnd77mz5P/qhLNa/hYwu+lf4+gOKhQhZj0u5S1
daelpoGXcAfllvTKRLx7lAF2eRDeX3nr3SJnJrQ1jPx/J3FvhPKe96hAP2vl
Tp/tYM+tj7BeuntWKCyjEmhHJW6E6NSDSTxPx8nC6fjUFlOvYNccJGf0yx33
mkaWxbhbaPmOJrwDojKBKBha5J6EDx/GP5V4ll7YiCVOyybFET/sGYHprDEJ
pXs1H/t5LskwDP/iLgXTRhgPwCPZTvidfOAHUpxWTSNP6HU3LjiuSM0tWNYO
5jkL/sOwUYYCQyDCb8+SYbaWNGW7f6EcYy+tGuQQrvJcvlUNn/rKGSghfUGQ
6eox9CzqFvHAZ9C6baxDkJlqYnd/fZADqgrWoTxbGvNWl6/XGIXsP7cSbB+8
ZBTzK12t585sKUeghFTMi2Ey3lK7AU9DCKF3PswC/03c/pmhPNB7Zy9Gbibi
eWPTl2EWhEihIcipScnroB/K7SPTk1fyJQpE27PiWfH2XAMNCU3m7zlnb7jR
76vOwzSnB9qTiOUSSkWGdQmvFXbrkX2/l57kFWv2+GKmFXVj/lySa5vmMW7H
R5ophuGMw93c3rqXoXLIXQ6TUYpmSWxfDDFmoDB0QGFR15C0ua5nAJg64MkP
7v1fZiFTX14o+SmnvLhOwRX63jRtRnWk128ngZ5VRhONx8LWxLVEM7rQMWFq
NJun5VV0aats6VIrMrddn11Sm0Njv3rMTj3mZNKNzH26VbGc80A08pe6aqr+
jvY+WJZ5tA6LVMdaLeAbssfP6tXTWaFboSPWSuSdwObeMM08VuY5g8s6L5DW
tg3j5qiEfOsaREynsncLtXI5IEXejpPR8fkzDNUpUvcZDOyQ6uVCyWygJW9F
bFoi0guPqUo6Hxpfjiw0kam4uccibaPskTFNGirpd2d1IiYXfHik2Wz1dCID
B3JHui2nUESU9AmzyX59scP+aRfHOnIsKNOaGL6Bog6Gx0V09sjslvKDfk7H
3H1RQuBNwsWJnHCwFLMX6H9KfFj5hAUuz/B9vUtF6L/KPNoOGWfad0bOQvpU
xbUHadhXBMsqxa+k5PRSdsMY3HbdkoMfifYGyFvHpLa2t8SfYCIDJzDgspcC
4/iPIHaZYH13i0kypLcbPI6bJlC/dtFXTsFcNU8AC1uZdmLYktCHGqsb5DUO
7c5dGB6GoAVlm5em0f4N4Z5Oj7JaeiEaCPPFWw4AsPg6HfFRJcHYPQL7CHIg
ti4ojmxkK0PD9NEfqY5PRiGtgMRtdf1h0ylu80CbfBq/+WDGAUmebr1ciedW
y8OWFj3XXEUyOvA9gVNw76L0hqC5npzNUShGdFSO/1d6w2hnO0IrKykzoNLD
C8JIEYs3Ucb9n2rRgZPdnlzD7RL3EnRiuPGzlhybQGFrxfplB+Q2IiApHADB
2kjvPcEZOAPBt8ri+Fl02icS31tdDCz8k6JjgNgP85FVoAFIpj2VwG+PTJ4Z
UTSOIg73hcW9DLA7lXFwq7NXklqxG7aCvmFPoA5lohOO/syXkv6cIIX9OjP3
ApUciXXbRhJkhv39pxYeqvgJfFTfTxJeWRH7YwFjZsZo0t0j9EDCgXKJLj74
NgVCVFgTyBa184DcvPqUoSMBiGHmO3ci4gY9CmV0M6bkV7c7Yth0BezQKN5D
TVqi4Ftg7xiDzR3Z8PRCO7os8uw9RxodG9ERMa71A3Jw8mpzpKjNVPBZmHCQ
iGtvxksMyQqFtkfBrG+HVbuRXrXweXo3iEKNOBFudStWE0oTqXQ3cfWw3TCd
AhjY5L1s0DgUKNxShS9smKFGII+ilj1uRsVgQzXR+VDnO5eplZXNgmshupXF
Yvocn4ZM54mf2KkdXr5pmR7rGZP78P1Uj8whltKDS9IZTVjYyrOEOtMq3v8K
R0+AmHQRwRvXkD0Lv59q5QpK1mLyu5AZtsk9OX2ktaH5srpFRYfqGYLcH/ar
IaNjFJeiM+1yoMdLdlnZZ5UgvRb2Xpvk7anvm5HMyfJRs7ORLT3ZR/P/XG5U
v7Umz+XmlbuyNTDT7K8aEBOCSYhcw91TmrNEaDEYVgVbJOxcbqzoulWC4iff
mcU6XXKFklgN+nRo7WW3/8NJ7N9iNHboHT2x8ZopK/g3YdpER8mi97RBo+p3
/J4+aE3BHGn04yVKzV1+MuSh11iPDSZxQrMUGFOTkOcysOZzfCPilpUmjlBb
RTXqUJj3YoYzyLU6b7QN6DkVEtTf0N+VOX/eKxvkVu5eXkPbgAhA/lSpvUcH
WVcfWA3HlQUoQ91qjdp0hxS8KRwZED9XfsDqi9Sm1DJEmP3ZEClvxpt3fXwZ
qDhf3CIk7wP5o1mg4Hzhz79esWeKsFHgJCk+pspWy19FVtylZL1OgBtE2tbz
TG7C68FWKX7RD5fNAnqlc6QSIZHfku/6+TiLihI+JyxAoKWow+bzmMGhcBL/
4RmA7rPEUVIq1akJWWeeDkpB0W6a9TDyprhpSlZK6E7SfzYhSODN5zsIY1+M
nG+T0r+xD7Fir8jWbjjhw1XVaY0EI3IjIAOcCgTs8Ljq3xaAExPca66icVBo
vzKUGW+hYeBFvCrkOzfL8eky6RD/itEGm9XrTIwzG7sA7/MqWv8ie54mrmk3
xCI0bfOcnE/wANBFNBBO+FsurxOMeeF47h4l19ofs2iuWAbZZMHp1qSWlSNx
5clJFvTaZSXB0crPo6ugqvrPgdh3pTAZOHBOi0QChxI20+k0gRzVD3PeEQv0
76bIXPKXw5w4JdHSBYQWBWCFHvc10Vc/8rFuC90IgeUA0831T4txN0XA5NZh
t7Ub+agNirnkw6yU/CC3OgBBp2tYDK+aNTxkF/NwwA4NbCaKKaHtf6jlLRLy
xLPkgFu7SInwSPNF/arzfY2s4T1DU3ZsdgnOKmjrBHHAbF5dXOstpMuOKno8
31QQwMqRCQBY3Remvj962fXe96rSV0qrx6yu3S+/SE4s7gRp3TvuP3cq/N2C
7tn8B74f/pGmho0jPVclTb6USAunFp6pBF8tRz5ndM9UgmeJ3YO/SRzpMFlP
kRYTEswLgWYA3mzlLXvXVcGQwVNNZtoi+mr0RwM66gJrXD2r3/IbsE9x3Yo7
9BzZSWVO2gwtdB+tprZ1wjzgKSV75AadLakAWcN9r2Tn6oSz6YVSyYTX4g7h
jfExaUlCC36YBL2j9Ui/GXr86wEDlzHVKk3mcamq26I3kGzD9Tf7fJ4JHIb8
1NcVh4Cs48yV2ElN2MBqmbxplCpzPP7b+GU3syTucy2x6N0i85R9IDvyT+xQ
AOSvbEHtGwMiiiMELtCLDYOCoQMyq644LV84RTEs8gvL1Afm1HqNK+5hqqGZ
RxDUg7bk4p4nkdjCDZtvzynhSixvCFY54Y7kFlDaWpGaVu3ZLbOpw4Wp7YQj
lZCCOSOH8lLlKYEAF7R1/11zvebx8ch3k3B5tWgrP2YTk3DJ1klaJBlbZJZi
3Tx+cTSC9YOc8tRnWAyOw4KPMxclNV3c3lKPOU+rrsF8RacUgpL9pLkSJKUc
ePnowhXEalpExVvmJCVO2TT5YIqfyAeb0+LiFDToleJ4/MzRWWadXJ7Bqj4c
tns5YvZmRSXPVbcCXNZkkl9DAxjLDpv2gOxRBBCyMUtvb3x0AG+lOYWYk8pM
XRFvhafK8d/t6/T/BY3OyWIGcV4ltDaXTG/BXnG+DTAjLQs/eQMCeKoD968x
4PdPNdn41uiWviDXwgmoUV0L1ujPu4Zh+ZjgwodfJO1ljmUY6RVs9BVvYBsX
JNto0keA5t20Lp21EfVNzQU8oXyROVk9sr2CYTTeRpS1pMIiTOmMVpKirxrA
Xlc3IpEk8cG92QwqLZGuKn4NlKjKUU58sYE7fPqHraV4egZ3d+wc+TeO9WcP
zGbAMYEkER2275qU792d3qQPlFF2H2+69pQs8tFvXJk4jQIPhCX2CBTIyNjC
xUsUn99EV6jgPQWWgK7QPKI8IzclKnumxXZKxooOdx60kcVYZ+8afk+fhjHv
PBxED+KjkyR9wCr3+xquoog1QtfJfrJSVy/l5jAIwlhq9shaZdDrnEZZ1J+2
ObI3acHTTeJoQLO9ISJzi/zKDNH6w8H+ACWTrST0rKpUNeO/3De8a8Na4S2J
GqepdEh1V+5gBHx8hh4ZqcICIxJ2iMgY6YDS0msO7H+UF8sPpaVC5SsCJPOq
8DsWQ+FKC2FZv0pCfc0QKuGcTHAHwbgkwaFfqKu6MaF8888YcInRPUqWp+tz
sfUeRFxWM+BnOIJoL0GXUyRHSHnV+EYkiwOVMDkJdaI6dnP/JlXvvmZVF5ct
jScG/U1ft/FdFLEIte3a5eA9g+I1iLjT+W7c06xXvXevn37IIUAaGNopAo0T
T3NKctM8o94PZcnjWdVcS9dQsyLD4M2OICOsifzn9upV0SRcBEjmUnjeYIWl
Beq+JtZ366qngPPEDLnwAaAxy3Fmf2K+Zdd9IuQMqEPEAnRfoALBbZzSW2x0
/I0H3nBaQK70UE4LkLKdWKXYpW0qslHNSiuLvfgX/bTUU+E4C7AmbRpiDMlq
wUDg/wgt2UH65WVFd+CzDxXe3VDP6JbDv+Xaj2B2sNmTZBtyp5aprplNl7/k
6aEFtB5CIJFSsuKamReTEtwPUx1/F5PeGbeHDOHXNFBA0mZ50YE+f+lsbayU
JPyKpzuUnkpQd0Zb381sESjwIsX3H1QnEch4sGRu/9e48GAeiI42WyeujqeQ
KdENVV8ZYMybij4HrJ/VWdHl4SHSziM+HUldH8aM9O+kUTDA5eUP1yvtFFCT
TCSNqfrpdauqqVUWDdkyk0SB5fjqlBT32CuAQfuSmdeyo49Fjldv1gTccL3Y
RbWbu+PuIX84mcSsRXM2EFH4uPwagpWp2guBhJP7WBV33YIYp82n9B0OAVod
vBC/dKkaMI5xVLZGiv3bocngesHHGPn7/lUyrTN7UDlJTbITPgA0b2H0ui4F
iwPoA+J9GzLxx74QNrQSyIykz5ye7vV2iszOReLDhvjoxJELd2IX9L9ZNfo6
FC//SPwhqDNZDsv8isDaW2+SCv4+xsxW/rdS8XnIZcxR8nGHTE5LlkLhLxNF
IzoE8Yo6PMpmX3eibv9JYXyny7NfNZ2hzKJvVMFls70ceAZQGudZdj3i2yuU
JGb/lVoVRe2fjTTr5G7h4RPoJ5p1XgVc8Lr5nCgXMKjgPKGtFpkI60TMuaKI
GyZQlkEq336iBYN9K/h3eq4DJ3/4tVBZD4tcxiZa1RWCgDRu8WgvNXHbWGdR
6fklZ2RjqdNfI+saQmuQQ/vH7npyUHw1bxBYXWBcrKFefdUukOPiUy+894c3
TwHCaHdqnjLELMWmAD4S+B8tAfsWaue7xwRXPE7xlVK58qhrVBq9D9uzo0Zg
nET/M+rHCzwzfaYxX/TYNI5TwToz5gZ2vq3qP1m1dBOAD2hT/ZKJxPU8/laE
5nDzueqOQZ7o0CHA+Snc0iq9oxad8wMQv8kUG0AblK/ehi25pJJVHlyqtFyJ
B37Fbwr9DqvESNIWmbbXFH6LkTaDp8ULRxXO73h+we1b96DvRGgEnewyx1AO
VSUv1P3LsvdiNo9b27z7bzbj+cZNMSKTnHGntCQm4y672Q1Xby6PFPbEWVw9
W1jDo+xKF8E3A+Vr5UQOiwoIHvcxS8KPEeKfr+sNc6XtwK4E9ujw3L+uurOz
D7t5nO//xh/LrGPjcD8MzAViDtJfYXVkQ2YThFN+UmuywhieWR3jDO3hZljI
pXaPBn08ekVXOXzYV5ij/7oL4frlnaIpS4Z2wc8TWA5MaL6QdiqmZSoGWHpd
AUgfvGCSPAFXUHcL6i5u17BAc+zOAd872Qlm6cCcw8t59R2jxLC/5gLdwot6
yiR5uxtWXeaw02MmXaSmRbuNItzE+nY77srKOXIlRfmSFcJy9+FybmnZiATu
7EiiCCmAx2A+6lctsKoMGhV6UCH0lO3QQ8gHH5kgye558VvMZloNiTABAzMV
vCsDcFky4jRa+pTJC9XhAGlo2RWxoOlsuUvEpR9ZAx/ar9o/TZK0Zb8jDvep
IDNM92yCiqwgjS9juCj0flbj0jy5SH4pBTOqiASKvR4Lg2xY/Pg8HEeUpJgT
AFp+RDAnTb48Ew9Od6rPebkCjKqaTgd8nbeRRiNzs4a1wYc3zqbimqnOryJN
cMYy7cgMwcBZ0Ajuw10t8T6BrVj5PWAjOdJ3tmsdmQinc7bOVYanPzVrdkWw
b/xxYZSgX9YwCjiYipU4ewwHzNlkRasWHkPqnRvxB/XBs1+JEebdVYOSQP8y
4F9L7jTA93/uMk+3WTgQI1Tgjph3mDAnwH1rYODo3ZuvJ+zc4Hu3bwCzhS+u
QJ1vibJoEib2zM7ptf6CATzHSsz/mhLWNKqt/O1kDe/Ob1k/KeaSYsY/7AJE
B9hA50UTGRJPw/MC7ZjkgL02e2DuBdnwrFHaLyj16t0HaQrTtlAqUt9qRLop
1laO9/cwvjuawF8GKUHZ6GPeCME8JxbG374DecZiopkY/IRaR1EsY8+cqwzK
v/zJtrE/b+qeI48Q2KRc2c4FYNosOYQevmv1GQT0wuO1WJPrn4U4ZJrnmxtD
SYQY1z1v9bR9u2BdAae+VxqjfhiI2T+yKA+79MrGRROfI70dFUI1ZvjsDPwC
7ycatWHA9+W1RDE65sTc0ZywLaF7BI7SYt+mOeumbtjXsaMIHF1bH78JpEuG
tvdnKjFNPrzpeUzwhso+rl10Acyuo5FzBBuyB19a4V5cF61Eeuxu5L4tb7Lb
yC7A7t1Wn668w4UuqpwmawcQisyBBIfV2MFntspifcsL3Q0QEYwuJZyxBX2b
q7ENVPf9Y4+qBl42ME1m/QgdH0fKPuiV6Zl8hhNm0qWwbJxTfofIn1eT/KqR
LmViy1JGB2IOtkHZMhl84FPk/F8EGImXPEvhb71agI8dnA/SWpT3zBW90+6h
l7l+Irfm5P9DDHvy8bGGoDKa5Ahe2pSmInDA/h2c+d4bieX8pUYnBZ3nXhd/
ueGLETPKXNLAE84UZK56fWEGj3x4/ud2BNKVJkBxOapvOKIGyHBAoqFV/iNw
RezEBl5RxNX0BJdC6j1sz01iIeK7TiuxsM7ZufN4rjKBly41rLsk92QQT/Rh
4GLsyOVdavl+KvREU4crSQQrVzaFXNAMVGv1tiEim6/NnBKcS68C3YQj/sJD
ic9cAHigIDLfciPP7vUwVvSV2CyHYyf/Z+9r3s0pbOuKSSmJetNkotfVtIKt
i7/sqQbVeyeiy3oophmgjc8v/5GCyezc1q0rEljrfU+ii62NGvfxjS+vG1tj
DEX+d86jDxHgTSdh5q5HUbet+o9E7lsZm8wjwJR2q/s+4lZu97m38UAhUvWw
RSnm5tl09bA/4viW4Gf3+58rZu1A8NiS96dR/ruK6dq8S9tjxO1XiQkhXEvX
H30mGjq4G0hnxsAPWy9KIq/roSa9Xxuhfmmwc0rIMzry7OyZGFlakaogwTEg
TnC9MQGgJSiZly6uF5r5lZJHbu5ZuKw+3WdRLVPEGb/sjX7x2HE4yv0AqCyO
26nNuCZLR2ViH1juwxWOw1GMsB8URKHqOlOTzf7MyxlQJ5LTAwDPsTyUIk8P
oVYaMr5IpStZhaVuJlVD821hRDk8WjJ8zqJVq7oZsjH3fuCUNMhUVSVahp52
NvtunSQBVwFkqPvrjUr8AW2xIt7eJnjW0gsY2duc3s3Ac8PLdDW0wnInraEZ
yw/DRn3cDshrxLCkPxK559a+eK7n2u54is8OTf2ZLY7agzUJPi5gwv1qCItR
N+MOcFaAVxlx3yco0OS+jKqjwtQ3Qa3Jt6Q3BGkPZhRK5kC3LLGapS/QHs3+
lx8dNgGLx/rVTnJJaSiSUWtXk5LSLKtwvMjWnME6ss2xe71/ISxB4elMtu3o
2Gi699NuZjZBoV9JknbKMSNq1Fs1uWL88RY4iSe+mqUPvRZjTIbDQtuL3ky6
U9ZTHOlAl+VxnEW2GsX7QTyCM4bolV718Uq/BjrQqoZHSwge+ZFkrGDdiZOF
VE3gf7S81NCSRIuUhdzhN5ylw6VPyYKqz6CsTtXJqOcaJzccGurrNFAMlwfe
t/PojTc6qR3rVV2O6LZzu+773wJ9fn5WsCqtLh7kuZWJ6aHW0urSZk3Y38j2
6yDUMvVsxrehXF0nsfVcoStUK5DG3G1jOHysuYu23pYsgH7SizNxwjEQ2gRx
bmYNz1uhWr0EtUCbudsbU68VXtRq98IcKvY2JW9lS0dx5rwkKFxsQsMCrukL
DXTQmYZG69HTe2jgQRNQZQGgOrvjCLcsRdGUeBBHnDU88MYiovJXIq7uNqQ+
GGYe1NXscjFXFBtgwaCukY12pTkzhh+wzK8CdWmTqRNZ7Ze9m/j/ueS6hnye
+FbCbS/fgBm9s8JyVoPy+KhDqQHcAKMpQIW7QaEviRtyGuoO0ufHQeshsYgW
G8U5SD+5OQNpPeH+hjTao61BWXhohE3gn2yDlFu811FJWQuwpLTz3RIyc0/x
AR1hAfmSKMgppXkrHxZgeaiBWEkvjQmbwsdanXmKGzhEzB4QtOadMtfzwIGZ
3cmHX9eAAMtNkHM1Tajcs9+gFuJ4D3oJ9LAotXg2CrOGuTtuxo6ANwIeE4EE
z3mzyd+znTf7LhU+WdJsl5p5flwUPrd9i3Zqbl+U11xaLpFYuVZ9Dvh+aX6h
2/qohqYYWho8a0vzX0y6MEuPOVoyR5e6cO7Y3tZjQ6mCxzQrTzSn+oKGn+1p
23zcaGyjs04ToL8t4Z2zpn7KXPUFnXAo0LSHGhUkj3kTQqqu0jvL+NGERZqt
RzhTutQoBBXQHkHkRdzwSKuOSrXGLBHlWz1dRYxKU5S5XMHsSzHJAmHhCDKx
W6JBhD65Q06tADtOV+wVjPSp987BGBZ0px3pGpuA0rgATdyRXAabLPdhEVti
jOcHKFgI9JIWbfwuHVjO6P3L1jAE1MxFrHIP7fDzapEPkoSlF4vqRN0sZFw3
ELSgegOzj5V3UEHvoj+2c7I/2lGUgLQW06r2DdPm5BKoou7LxIIISF4bpsfV
2gml9xH9qj/Pd3LKI199lFsFSx6ZBMY42V1blM0pc8CnRrnQ9GKrUmvkiYX3
5vrGtTezahYxfycO6BEJCr48t3hQjCBEnk5RD+Dltt00ZRVh7PLpjyt+GgCT
fSSREp5JE/00gjNvoqW9j+ruq0L6iihWAiXCSaIht4mJFoB6mxlj7GvUEsaM
P/onQRuzIFWDSfdiQKP0R7tALOhwp7mOnr/UP1j1UUTK3YBZWvmjHHJ1+gew
9lyb7xr8L1iChnoLKXM/FvquW9TS+m0cqcuiWqMrrO4bZEdRC/rODk+cnpri
kxKSXPQ/3GcuTRV2xFiiBU+X7Kavt2V+PlyY/q5TX4jbm+HQ+toNP/y7UZce
rnFBv9Je+OgxksEbEq/0HeEoUJ4MTxv/+/Fj49wNPw5nOU4ytxlehYJfZf21
oCHHX7PN4Cxt1um0MY9Mpw==

`pragma protect end_protected
