// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
j7RTdv31WTM58pNui4cpjrh3gllqHzeqMUfyyylZtYKGmu+d1zMq2g+f2nwt
DjAV0PXRwUnxBBf4y245hhcSNFoMjg6q4kaDbQiNMr4nGsv+iE70iJl4Q/+n
nGct0UPtGu0xjsFK+V+N15XobOYAAflcT1qc/ugDN4dgahFDLSRNe/4TCEht
qhKsUsKkTN/ZVMWcEs/thKIUWrVi7rt0EZZiS4Yr8vxxNpCUyQq3Iyr61kh7
gOcwgiv52MyeXD1CFXsSZa9HhUArF4K423B+qTuo5YEufD3VuWr19Yb7gFPx
m3LbSlZEUKiB9l9aJI2KmZrmpJuAhNadKDxaY4pOng==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
II47Fx5ttHE1FQ88v5N+ZVsR6FcVCFRo7oh1qVsX9X75pIdifnUzWZguIVfi
6AIX3uDUn/i0H817rWXQIGkq7ijriwgLkyMcFxx6QeAI0VUkYg9sfGNckcUq
itjBcw94Vm+UPRjvfWFexIHzzfaHHVY+TExWhx2KOo/8OocARX/0wIMBukfN
vDmavxeFBon0zyY93LqfT8ooFYEFmi8zEBoT3NPTA23elp0rRSvnd1iuxhbd
/Tfa0koEKsXtQtvsB3Uxe1SaoLtExC9qo9xPunWX3cNYkcBRIqiTZ90DYYV2
o568rvDNnHE4RtRxf/+ISbC27FOQpugGApo+e+AzXA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
HXJfEkA2RKLaHOpbSVK+OcE9VWDIfeD4E42Vph7V4P2cycDiPxsOXdZisjxW
1jMCaMbz+IJqcTdZA3k3Ezja/Y6cpIUW/zxq5lbOGYgQ/bmOfDgHHtgjTiEW
sQRkVmLe0xwmsQ2snBztcHueLgmDXRRQGnAIyMkZ08gnNU/VwDOIY+KBUunh
iVY8Am1TE8rihKRsDDDbf1LoyPxrr57CBHBdCBz5BXZyXrlSesp3wWPO3iYK
ICKvrhoyVia8EApG04yWBGeXVNSRmgeWyhNuHjpcjfbK5BM+5Co+SRLydinz
LZdYYR1UsDj9WohLXSigWQP0j7z1jndZat70GvVRyA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Q19R6ha2anQKLySM5QH8fprLSGItWHljF64LYoAndIBv524H8XlfMV2jSDrV
OyaBsKa5KvIn4SQEa7DbaOcqaCZYMIn8aAWTXntJ0emfXuAbIYoRQ0jZFDhc
3yGojeIIXBXOWWd+A+3jCdy+GP79HgPt7VVj+I/TPgfA/i4gCO0=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
qjh9Tz5erytPC5ycMgehYttYFcPvE+tJ7nmWaDI//PcPcfIz8gg4czjybeUs
MI08aAOR8D/5hMvDV77Apt/JojGzcbtY/1e5HRiTVn3guqINmSy0eX/MqNi5
y0766d4roIpAEkxPKPxzwPLQBkJP2G6mK2utjl9AKR7uM4vYDL8jfWoOGaxn
oT8nEP/SqzkXLJIV+x1/x3mU/u/NNXO1jWQZHWV1wx2ZdZR7f5CryiIYfMMt
uN9t3RDDntI/SzJ/3QelOPy+1gue04WLvHr7BsCacM+Qnq2hX3FWtKci4lsS
WmTwMH1XBizV1PwtmMeLKlMsMivToKB6FEIjwH2T+Bz4O/zXlSDxIkWOAIJ/
3oBJSoTr1LwEYHrsgI2YDQdERyNP5VuhBRpWuHRctSq9noUV7Re6e41+wvSo
ZyNx2Nb1sDRn33NTRI9vHIrXmTIaXXFeYykoMGVWe0/tLfO4FXV38YhxtaKI
CzVcHzpvEjaVFB/YVrX7PAzSu/vZq3f+


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
dcCtSGABvDJPnAe7YPz+/BFDQGN5Waq2BKHR74zbFcskrtMogyCZJyBIqAnK
D1vO9HahrQzxwCqhMdlRPet0XQO54SlmFMGXpTi8ti2wWiesUHlG4xZjCe84
bC5+mOKmt96UGXKX/ixHu9rXLmMaitO/BlxLgtlQ/CcJYEukRFA=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
eSQqKDedTpCk3Vfvg1Tudx7aQV50dNi7Y4a+OKgkLyC6Cq5NFCsxNVjQHzPU
05TiuWd6lmxMz+d6fnAJRbZIPOW1J8vXPUeiH3kDSOyWxLT5Fz7ckctLkuG6
vOr6NZBmWeThVSp5v8w6Hbaxl8jyCPPKuPnzn+lJoFpd3ep4k5Q=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 27600)
`pragma protect data_block
L0A4/ce/43NpCjr0HGlHB51HgMI4QyUDpQi4hJ/3/hZuyGx4grGRSj9UfpDR
Lb716CSkIhES0q7Rq6XTfJUF3z1Lw3kT7uXQphN21CurnmUOoEF+4XP8k+wT
Jxr2qomxiRMVs+iHVetRqY4WbOVMCs0FJxtGksF5IDP9c2A4w2OK9fTETF0P
Dp791GKcuhcL+Zjk5+Jj78+SkQmVjJugKKPrW+fuQvMzl0mqH193CYGsLESh
mwMplWrVFHTF8KEf0aGwdKdKts9wCN4QlIcoKiIPy2GcS3Kc+j2A+Og7f5QK
nKyvEKqJ1kIVqZmvONPg2QtDTQsPpVA+w6UskGd2gFQeifAc71Xd20HfPV+r
IwH/h0YXifAlgzQWJkHasBm4dcYW7eBAKo313T3mI1DkhcYLPOsPi6LxHHxI
M5PUu0HyL0AFKGp3gv921hDMRZD3MCrRWtwKAuet2SGmS9Q/j/A/0krTXaGp
JiV5zoLjwmJhWeNKKbPBA+uxDG15uGgM6uwW+T6EHf3GCYEJij/BlFxpJ7VT
f3MPJkCIuRcqgCy153O3juPy5Bn++iY9Nz7c6oTLeQaF37k6S7O01j1NvFNW
hdZrYOUbx9UH/yuSZIITFKRNUefTcy3mx6b23xb8XO3NZ2fCODxN7hd4ZZyS
/2t3jVMbbm7Uia0FH45uJP8tz5piczoalLU88nqxc8om0ykA2DVcz+5JgsuG
SGJ0mAiutWfZKps7kvLacuXjnfy3QSuJcpnfnJawrGm7BO1f0SFRRnAeJIFT
ZW9ceieh8tHruxAkCi9kfuVTPOCQsuAlgDlprHuGs9tYPwXnuuwXtKnITHAJ
9322gvbqvkleqksnhA/yqEIQKoDupxo/Ik2JW2VessnTpYTRKgxiFV/t8K27
CJDCUuw6/OmLeYZNoxGGyU0aBlAz1fWyoyP56MyAJ0vkxh1MxH5flqvFBaQn
XbqtGZjkXqtmFWkFbRkfrCMd+auX20QD83rLBpD0zeXu0Wdnijf4shVRRpFJ
YVdg8iKFjrk3mLVwbDO8X+S5mh4p+X/ZAwakdix42U9HoEqnWirpzoMe96KT
8utQbpehesGFYrvhdkNeCgY/FaSklDskDKv32rDs4YDIVE0JCHERg/abpv3y
6kM/6gk5cbj7mNsiovXoRBcEXnpvSsZ5izPaXS+Vw3wRRXnD54yEsLhsT1k2
NHkU+aDLbzpQ+rF6rbwxiHdRfju3z8Yzk4KwM1RAS6Vy9l20XuF2QPct/GN+
ugU6e5/s35R+7DBFAXqwnk+/ktfxj6WL29R+DLasIFQgFF02FdgZ5hF39OBX
8/jG1Pa78NmYLjYutAc2wcXQ7wwUS8ZyA+dFILLMCrcuR/DyejK9YAs3cmYz
30Tp4DfUEK9LAXOiVlXg15vg2V50CLhFU6RosX8zX7SdToZHFS9yrddRHYXQ
I61bBiVPbkER8LxpDS5A0sQYvGnVsqZGJmxdzMrVTxnhyYvpGg1bGvYsvlPy
6p0Z+ANE1u2cvSht6eqZNdi2SIpXXGjq77shWcy4/cbh+Cg2jy8wpujBegvV
u/CHHfrCJWGdw9BP7uzWtPrDgQppefmytCwdFxA6wQ142cxA4jQqoHkbHENl
ugYrk+4ssZRLg802zRxN8KNyr4gZ72ijppAtofHxYSHl6CaO9HI5Wx06h4GC
6Br+fhTJKKb8ZPFqV2vqzOtt3uUMXiDtDLGZd9HhbxysKuH/PIm4Po7jOIjL
ieHW3+qUSugamggtr19TiWIRzVocHB+rAhJs40Gmc8mtw4PQF9BMBD8VXVoC
rFoZcfvMPDEdxY8viQc2eHgM46Rd1TEm+3IeX44imHsSV/JNYuYFzkbAQvY2
eCgBatWO+ZsATx2xjseJMSfGTOPT8qHTXaQqNBxOGu4AIvtkT4IFPAkR56rT
6SqlFkvqS6/hMkqjbSVCsEYDdu4vOXobRiVvSGPMfUeaDtyEpQDYE8pqq+C8
uaa9RMWc2t0fhyyVFAErs2MYYeti3/6IOKb3rQQH8Oq4sOvaU29Ej/zVtLLt
iMDpEDU9i8NJLMn9wO620DOMlVbLBh6GBAO27TdCnGB4vKuBbnTN8j4RwGRC
de1PzwCBMGuH97Z/4k6KLlyTZuTozm8HqlMphL0Yib/mF3SsuOJyvHqlocxc
x7Rl897oW3oN7CrAzCjb03rvUtFVtlxrJVukgsjWgRnvYCL+bsFQ9Tfx3wPu
hFSsYJFsCJNcI5nAQIoUEfXbBdNVk019Cd4+T8u3u4RuVfNrqhI7XNmc0Msp
XfA7WDsNgcDJPN6bd93Qm/qsvIQmRgmqSB+Lwxm3YBW8uhIfO2dU25pLE0vq
PSuYnXCNbo7pPE2TYa8/dLrCAV7MuY9Tr1EtV8Frl0KD76KdsRXy3H8noWDU
3+alFzOR9yvFiZD+uRmfVfLwBQaohOpVAfvNaxUGsSo9iasv5LGo7Q0+ZasQ
+7ETTdmrEhfwqBY4/K+0j6XeSyFDMwIZZ5QDXKvOgYkQPzFSRNufQZcos6hU
ZpFhqUUrC0MIHYY1smnGaLI4tNKIbki1gGOAkBDatERnc1o6P1G3NZs6miLk
OsoYQere8bEW0N805jxw+84mgVHWEtmnp/aF9wxz4ZaoymQLwyyau/OLvxpH
nWMabW8zvLkUGrFcBclWtbhfVeb05toUix6R8MF9BFR198FOubHK9TsgmlCD
z7NVjSG8Ahkuzb8jDlKrjHybacvbvHehG6ehAVdVLgzWzWoDIwPMXjRsxVd6
fUPRknPsVgEbzFtVMBgSv6Ww3A5NZicWshIlToXBvOHiHKDjlXvAEbLEsMvd
Rql+KLmnmfwdp5f/CEXZmv72ljLl9cdUPuw1q10cDvs3TObrvn3FLYL5d6+K
+MB0UEmgJSjjXEGkO1Jjp/DkuaRASyDJKohRG0eBvSXwb4vWjbalzxyR7XVS
6XISQvp4l/b/ImKU34ObDxNMaIE+MTFIzokdWXopgPfchayg/Avxbo3Rr+N9
Cu1CTck+th7+Nm8JqfWtV7LlVVqeVUscIqblniBLMWX4SJEOrdcWm6X8ODgY
Kef1jgjuqdt9uXqTLgUbxjeYATM3R5w93PbvdetE9R71BCGVjcs5GsKLQRC9
g3N3zHpM8n6GRsiW4QY4Ypx7Zk9+1jhKAc6t2SPDA2XieGp1ii66RbtLdnnv
8LWTWfM0aKgDa4S0OUQjIceCDrBa3f/49VUWOzC2/QUQX76Lpl4bapnTR0o/
36CGY9G2uvJmN5acoq3h9C2VSglZ+Kl1zO0GkXM5UC8WHgx7lyScDSPkIdUU
l28YZmoq2TR7U3+rMOwCWw2DcUkxeDAX/phukiKeLuf6x1TU5/ENHgrhX1s0
1VpL1vbRcItJ86083gZ7Y8X7Q9hBiak2ASPeUcPS+1wIe9zM7DnbXs5dBWG9
eDeKQbXCjOx5z5zjgMSWv4yXEmoPFMGdGvhDeCgngXrY3f7Wvq05QbOFfSfI
yIkYdK+LK8+3TbX2TUDeVML8r4TpEmE6RrSgtY8ElQqvqtamU0tfa+dzyo8R
ikkvsHqp8Har7Fw6ExCUXr5Qnu36COIAmGQ6bIYVUZ1s9pgNrDUOuVFR9vzM
F8knFADOqnIBthnFvoMcSUTFLZ/s0Ne+JjmMwSrTV+74O2Onc2lm2C9TvRBd
rwQuvWO02NY/K3R/gBgJjv1GjP2OqzPrr3hRCwdXLWB5T8xqG7K8haXkUwjp
pt8+L0lWI1988JxceAt1mFpDVsztNiJpTgdHos8VsgqoJJQSO+IxC0QcCiEn
97AwoJlIZ0Ty2SQWq4Qm+PDoTiRHkvQSBEwaBBDi00eIFd6K3MdyREsgH4oU
tDWZGctQlULig47HvS8Dv8xVT2rGFn1OegOZeH8UIxdyHMdsQrFSFkxyyjPT
XMLLyjfQ0zyt113TcfMa+3YZQfSgo8EWb48Ui5ZggbtEFfF/DZdY+8Wftwl/
UKDp/pkcmZ4QtUWTWumdmnfblcJpCW3P58lT9n0O0TDy7Hm76GuF/NHW/I1d
iZy/IWSnbkFNjIIeLX0lWRBaZfSk4ErOX2ONMznhYO5NSpVDRVjRvf2CE4r3
4fMYyBYhhSChnHat+xniPX6N3eJ+fx6t+P5KoeB0QQXfgmZwD4qFNqNSdFL7
61OUKDwTDhVyoasaCjorP5ocSmgDCEQgXz+SHVQwvqBvTFFBp3vnfKodLaPM
T7n1jseuHvCjj0NFEweKcCR7KZp+lgqDc9UtIab42VbVy2+zGuBitg8hwqxU
XVs6PoN4bbds10uiDA4OYQT8DD/in3Lj+ULRZtwKtJ/o6ApkBoU0HXrQQUvF
R6qxOUaTLG4kSszwpChI2XEY4JdM63GBvhFnkuXhaOgfC1hkxjSxS25oQb5I
ZG/iZ7XwOfVZwr+NNWVS1Qq03YwMHzBUl7cMH4jCtwgssDZk6xhOt6dm/Bh8
nltZkHBT54ZMjz0S5B+QS2QV8tvqfwC12NxP2eIxS+5faNI7ksLpJ3lBdPcx
iWkr7LNi1uLKtXAJFZ7s3H6mVc0LMPLtZ8QVOe+N2xg2TXvPobsOqPJ1/U6k
CfNjPmUpq2fURnmESs5/YQpkiWzoMoTN5iS6XFSoMZTWt/ybtTJvH5wQXRyX
B+7Lg/2m+zewpbid0dB8IQTbvNTZqeZCBgT9hEJBO1CdOk454e6mmNyHPQ77
ZH3ImyBbucOa5pf9L6lIyQv/4wmWSJj5Xx/fIJKj1cqgFgVrNg6ps/Drfj2F
w11TbKMhcb63EzlJRcLnZzmVzQKJQAIf6dn/y9TlYmOeqPEHgqVZwjhqa5J6
mKE01kRIZxl7oDS1jNKnRDvqFTl46uX56fuxQ0gLTaS5UwAoA0qbzOqCbYU8
b/R6usaxT/YCxHhfMHDU08hZEHQA/V/wSTtHL35FVaAdnkUHubVkIn/EezVM
OxIKuGc3Ro/9rE/FTVw+l7SVQSVziIr7j+48+0uXr3yteFMBR1/nu0hJ+iw8
FvQKa6SyjzlFStWfcSQDA9oCQtAe8leP1rCmZNOEJhJNj6Mze67dnTd4Ez8+
IGg5IgOcXLGshgI5Sk31dK04KZlSithSZSi4qatSpB9Ihs8fxAspkcCY5bSb
9w16l5TNY/4aIRt1PgoRFC26/YyVujlY9sFew2wLkOxqK8+jl8oj+JE1qjhT
ftaSn7HUdqQCqKi8Ih+wT9kzLQjK9J+hIGRhp/yZMHVycGT9CUKcG+TCxgn8
s3krqY+jqQT5thl6cVtHd0Ou+Syek4Tc1qAH4Ycfh3HUkzqW2QzbgxQuoKPY
7YjoNFOxQAdfHP3g65cOZp/FLFs9UZLUfCMmAfAEEya/78sY8TGgv1Vd3yQc
aKGiQAydPntDnnNlaufTgbwm6ScvtfRZI4MhxYTeTu4wM2XJaeSV7zo/hHip
XPtfOLGmkLP6HYkRtuJUeiKW2uGjMsJvQT72oT7Zri8AWZPfwMRSz9Ntiuc8
QqkDP8roYLBqfP9WI1KmlJ5ozxPvxeEkjYvbhDj3mXjhsEBpIOoz04nRlWp0
N2fYlgX25XpJGm/EhYFd4jdXHs9DMKxWi9MUCjj2fArDeeYeg5e2RBDAnzik
MfrSojc/H9H5xt3tB5Wk5GBU7pBpL9ABi70MIAWemhrz8zMIPSejIZxipXZg
y1QS8CxX9y/EZFdUJW7qubZgREZD/vMAPoPMbfFQ8oZH/H7UQYd3bJKBN4y4
zr1U0yeFsSm91cMbXEFvMYEfK2cHGL9W3hR8yVxEJGThWU6RMwF+VqzrfK/D
ym5VICmF+O4E0yfFa73CYXKbLrwXUdINiZwzmpcSruPZoFVruASxnzdwAmb/
O+KtwU9WudsWYVmN54rdDWH6fjTJKPVYvyIjqRVGckyC24e6S2NTG30GZYsl
J4841ThTnvQ217b0FFBz+MEauOKdOmuLwgXtoiN3K8MfPeNWw4QKa3gIEhBU
rKfqG5FmPF48P/Hyzstbi9dhS4ZETiggS4FcG16mafng8eb7A3FamCH4NLRu
61L59+hzTJGmy5UIhFUjC9cVxQSXEdg/LsdA58jAhCqAWZB7/o2qpTxiV+3n
K27KGdMpFL5W4Okx9dIDwfRxSjDZ0JjsHK1NhDEn04ij/O1NpWND18a0R5Fs
xfPfGyNUc7nb2E35B44oRd3olEBVVD6+qxYncbzhRYHl2z2ysYqKHLn28TsL
1+e8CV6Zf7mlGemNodLeuy104w2v5zrPxQDxr8YltTGQaIX96JmgTkRJ65Al
AVU60FafvhY4cB1WyVOTv5eu57NFiH5eFpL4gB2eXXePsquaBLUiXgqYBIlw
+XhM+8KPLfyw0nEz21ELFKeYxqRTYLHsoHWfnZ7x4oFIL622ZP53d/3t3sTe
AoqD99vA1maRg510covaz6IfcjdFi5+1SpCuoo5lwi1XVOV1oT0DP312Ks47
ydLwcxWCPvkhWTZ0PM4ehmDbAwX0QdCDa9c47GmugN9M9QYG/kchi7AKXQLC
YvYyBMecGKnxBktBcURxVN3ifv/14NHmuL7y3bUt5EsHvd6O+IwMdnb7+wg3
s1Z1wmWHXKxJ26CO2Fljfqs8YRySxIkake93up5IcZnKw0VqTBPf98O0XUWO
XyA8q+uqZxJvT9gYlkwff4TJ2CyonNhjfgeWeGNXyQpQjg78BiRreg4bQXAK
DmfvwgIv9ANjab33UFrpJgTLCm4WwC7YlsK6tSjOd1Q/PQgls297P9MDVyDM
piiXbI1DqZVcrlEFltC2BfD00KOstMzUrn70fRKGPmQwcjubTcF15b3bhFgG
XjkGMrlEoI2GU93HV1oL7Kx7Ooiv14XDGwpV+ourkjbD1qSAqkvtT8gNPa6g
PO1ieLG3zGNYNQh2sBXC79+0QsrT0Y5uRWBeBlfTDx1MxM1yOIdPEla7b8T3
YfoqdzKVyNveCtV4VViO+JKsPv7OxnScx2/s7MtCIMhL+vuErNNTVKEGVeSt
+8VSOVw4dLrIKCZiFC21FHdH+gy5GXIrzDIStBbJoCwHkQaJj2YPoYd9nF7v
Q7SAvjwL5kzdhFxaK3gffB6NufmRIOFtv0CR3y1ExtxM44i7UUqcOLN05Cs1
EnmDqr+DMeu0IHFB72u+wwleFh1fU4hvdSYxvROrRFI+FNRWBSR4MOqvjK9g
Hun5aBGtqEb/7Xkuqxevw9YXep9x/gW0ppbC5Fvg9yhRDX372HATj6XhfD/e
8tUtLDZyoy3lK8mgLx6/LRowQ0/32uPT4OawnEm3yorge48okXbI/i7Wi718
tgZvU4hs2lGdT1SuyhByGQ+4uED58OEojt6WoFw+69BA0+/4UyY9enf7+zvn
7BQHtsZY72itXxNVZmpoTvPTaiiJn5BiLGCP1z8/Pvfnz5VhrrxnRB6C1Ykz
Iih44DLJB4UIOysWgW3iKUehz7s25iLfqUBjmosuOJbB89p9DXmRlyMEKifx
HR4PTJpSTe4lR4JbwxkJPSxiqTHpp1mpHuyQrTVbn5w1hOai0nyQpk3a9epd
ZawUXIu5ZQ++dtBUS3B42h6PK9SKvdJF6a/ZtQjrqh0gkAUTnnCHxIt5pBfj
y265MVV0vZWoRhknX0z3AOkmEwjKnkd/bifjbYvFOTvPxZRKTPBOqlGRsUm7
eTYYUMk8BBpRkZMkrqnDNPyEAzDSibmVnAj3bfq8uWMQMbW/4fALKrDgSILG
YnoFqaMY0HtyplXMfaOChrq+pFkNgm2zBtZW+l2XPH6EcFipVzKGWSpmp1sc
D5MWHg17Vnzh4fj1s7lDsNbQvTzgM/CdyfEM9VGV+LZXw1uvR8SqD+DV8vWR
cCa9N3keCxBPmA9lOgMvVCfnyYz/r+hsW7rsgPhUHpo1MV7sy+x+WiqjpK+0
6Run06ZNtpqIPuzo2HZH9+4SbcgxLc8sjpbvQxkSUKR73kt+KJUmWMXzKN/U
k3QWzdyXS9hPkdip5eh8D6mOBm0+X41k2dYQ0m4GzY7D9AIvYFxBIofr/QH3
G5muk9/sr/fl98d4FK3gDhyrTIy0ZVmnJe9kshzOcS7upNhtJ9r7JILDYhzk
u8vOGrfBbQZK4bbDLZgLkyKahIOHaplB5zxnmbgufhXC/eNAqSK5y/WQ+TNU
tANgwmG2HDUDCUlUgS3m/rffMC/1A5hho8yTzF7Ycjq6jBUIgBL617TAKZxt
IStcHCYOdXjZxOA/KEsrDh6CqgPnPk55l0X9K0CO0UlVSBz1m44s/YuIwYzp
PAnHP418KN0P2ky4NGWUySTH7XI/zwQCfpn+mvFUNPS5KauS1Z2xVi4OJIAa
jeiK+eydiOzc82th0pgNdAL/IGIkX73Q18uzSZu9nPvy4xHMrQjNluUjEO+K
TPJVy925zdgikkohhvCV/GH/pfdgNVjgnGFKoyKrubOtGmsXusY3j1fnM82U
D3v1D4TlZc4V/+g77pMKq5QJ+IEEh/+Z7kUMK0fKI65bd6rxeu79w+0J0st4
yz0kl/VfjeorAdY4XiG9Q17zzdg0wPTF7bkS1MRrtMvdcwgvOHtqFgUcm/c0
2LjKWvlw5hTuHD++c4OohVQJncTNfJbI5JZFnLPETujnZShK+ywsZt/ns742
VEB8N/mQ+0id/AavroKnGZBXv5BdHE96SVI9H2UWzzlQ/p7vgcg5Ywhl9pva
H5NlT8+JxdlSoWfbCZPmn7WyQN2t0vU+BXu/0jqZ2fleoxBjE17uoxn/Wznw
moeVisdNBxTrSIBzLFz75cfCfGoJavlti/dE02lLlgJnq1t17ezNY/P5If6v
DHlfvI4+c49mB9mzNn4vu65Caw++m/dFXVWSklC1J/16/MANbUNY5wB+PZP8
+R8V921sddDIYc5/BbBnSSY4FKGrkG0BueLG1KGLSQSLQAbYYzaIt/+k0sd7
koc+6xWl28FMF8u6sjCb0bRDzLliEIgbuUcvNKjwb27wulO32doSHrE1EcYN
pQnv52xssHQwnKFhOY/9bqJpJyxObrq+OdVoWVxgPpmk/Di7ILylAJimSDTQ
3a1viMcCdN/dWr/W0zbh6Kv9VxIV4GOxihbfE5GQC+HQfbHoX4Jr+KYqfiIN
PHkSnjLlb3s1sRJ3cYWj5RWa74YbW6lANomlHyOME/pwjjtemBZ0QytXiD8B
MTZMEwA6AAGUyQyPPodPNLkr5wrm7ezHpLvHbk8Dc2xGKVhL4MKj5k4WmWra
I1GsE90yE+FQkvTIFGlaW4KhxzSw4dx0Hiez/Lpumo1GF8yhLvyZR47dgCRI
DSPzF7kSvEefefwmz66AwEp5k+xzbYVn7p88+4YnaJ50WvoYcE93h6NF5IhV
/EzlqpkVqDW61WafuDV/z7XQA1oD5jnwR7N5MQpSfwz+P3I3hLjN81m8fr2/
zOqoVvD3ID2SJA++sAPXohacpyI2gVx70Op8kM1Ultv6Dxh6U/ezjFSE9jra
gjSKqTwu7lo5464ha2f+jKVv/mzCq0ssrgfpk4bgXhD7E+Qsd6aBDKpw0VR1
oJOCwqrWFK3of6isg5lo38n6Gw/v5JtjwmtfHPksHOwCWSXDgMzzeMwUXnIN
csdBNJ5F0LvqtNW7atpaISmTBzndtrSWK+b/agbTd87QmakY1hcramBdvunh
1NcvkAQQGpJzrdZUZ4IqtbBtF+p5a/vsiMWwDmLKguGcGFjpCEATxb3yVd14
ef8BiVoFkDPb80NOJhlNGt2+RPZgCTeZMJ66hFUaQW9NfbgtcDdUMI35+qRb
weCnIR/hC3+MpnJmoQCo0fMKrT5KhiYKW7liVQfBFj6sig9zqxoxsAnkNOXd
yA636DlMQOFClEf2OJGsaCLa0ZF7vvSJg57LQ3arpE8zEH/6RdVD+Wnc4vgj
jByA5JQnnR6bEThcCDTxLJPwYmlEaEZuHEq2ybEW6H5jNLWSscryTRkQLqi1
PWwTYNbmFk7i4diuY6pkacZn6u85lt0GoYBvas4lyqLfGbrax32RP9A6235J
lIB/QAxU0769my4dCExncqlWWH3J28qd8Ngnm/KZlmJWFNabRKJwPxlVcOWk
nkSYU00s+kbHSNa66R+aYCARWDIM4o/QzPOjLDLcJNmFcZxR5DQq1qSCXhkd
g9Q9ATgfrZcyK9UwFLW3yNChyQmktPzSF7+xcYWV3BJD1o2m9fhp8s9Md9Vu
EKbEONvnmh95cOqbxSmOTdW907D0Vdwi1Mq53L503OKaGbmyh3h/dbvEwlYa
U8xnmXWBHukUOmkdV/MMFumeRSH2vkO+fG1EzOEEepnVojIju7zsxfzJ4Is6
+Jk1FKvOuqiEBZo6IXnKkTEflU0Hv5CtJ25W7jo0Q9qqXKaoeTXF3x94jUxW
aPLVANaLcmt56X5Fsn6ZuMmqybYedbS1YI13okWhsDDbUY0oIEZbXXmrccW/
pQtsf9tyDGvUuXB30n3CjR5Qp0YPyc5Qxki1ub5lxcrok4qttN9yAvMsFLzP
BDpgFvhiCg2r83WlUrcS8b0Wdxur2keBWkdu4PdDnZF/CsD8mrFqlFYIxzmH
pbSOnl3vwVfecBx0Q1hamu/86GmMfrqXgMfIl6mLTeuwN5nGON0IId1rthaZ
cE17FdxfSDk3Dkbf5KX7n6PVw/elui1yY5xqNNnf5juGQc+kaJuGyeMwx8OA
jUdT2OrSlG3NFJjyTHB7FsX2lhuULyw3yTYaz/JnrHYqDJeye0/7P8nGF6vA
1Fap/n3uHjnxYF0blsWQYWCxktvzy1Mul7g368kB8ZU7cewey/ZPDpzoHpDy
2/XF+ky8i3bM+H6yJqr5nzfmWN09ORDmsk1HAc1Zva1VHiorfxr7TmBlP4nw
TEHDpMLM72qO7F8PsYv2xNUkXPhGzPIcCU/bjxcvwxj8S5QHToGPuzQf6MbR
ogVK87BURc74eZAucQ5cRnsN+dKLiD+N3TjzeBYu4mBuTSRiIhNNQ9+cimlN
//CGQnIz02+Vx1VL0l03GVSMeWcHD5eB5hA3ukawkU2vSzqW9GtizclhvXxI
84QcFfO+lz7JglOvETFXkH3Xyh0zwPZsGZKAHojclAVpBHL3eFVqM+8GLAff
/yTVBfZkZCKm1CBiIjcjHoVCKHZvQLYSuTN8zUk0cnEgVD/J5FvX5xd+Gw2y
Q2GlmygCtW8ZqKQ5dKGsYDSPP/+tiUB4Nc63qNxPQoftn7nOOO6yZM3TFSlS
8lqmY6riXPA0vw81KF7qqwfefEk9YpThUaxdfw2yjZOa9CQTBY58aOMOeMD/
HS8IONnAn3BCIV8XJZIQDOK5qpnJkx0l3D08QkAWX6f+GYzELtAcd7dwj/gO
FeTAUGWriJOlH5fX+0Ur76VHNxJTRzxY4LxJDdT79WP9YU0FdMCg25H/RxKq
TjV2LWwMB/dA8UN7j/08Da/qD1Fq0Md2TriP9VirS5fpCVndXq0wEQoBATOL
hXtLLldIvORAqN1zdeKTjYWgS0HJC8qAycULvpFRLjLe1HFLvUOONVvCnpwi
TDNdMJAp2pYv2zyS/Xw9yCkXjj50oE+lgej+LWVtZ+8RrVB9MPxKJw+aJ3lN
H9mrW4iIzZceFPdvc2pdpkCBRS+gtuS3FHOIpP9k/vuVKZ7oqc+Wp3Wjpy4Q
Ppe7B+LQ/VfDI2/HXaLMJfpkKuxvHCqA4QQX+mN5U+LvR33UromdOiQI7x2B
JCdmYsk2DetsbJF/wD2C56WO+QWRrDT1JVNaBPrjzDl12ma2HN5LeHPtCskT
O08qFmdAK0BvsDMBAB+ZtkJguVBe7rS5amYhJDVYN0okH8uP1FlQ7pogZglS
wdDHo4Y25rAYtFvss3c3fpkzsWKqHMonbqkOg1sNzkohWCWxhD2ReHhHFfpf
7W4HIO4xcw1htJVm0LNdOhXIANxYZNko3eNAv/+2euq/4JU60MdY1ZGK/s4d
fgb2GY37/pD2V+/u+L0MRUNVzONQNzzeOtiOAGvzX7xe+J3Kt8ZlVegofMLh
0oII/be95DCDG9+iMxsXYMgIJTyhRLvfag2fY6fubui30CgE3jBkC/WMh8p4
R1/e5JA3wO2fQX7DtWahaVW7o+5GClWqY0jQ9Po7A/N7/w0R4A6EXN3Jvuz5
oKYj3H32EYshyOEqwmWsqj+FmfFHnOb0Dqo4dYGQIWjAuGWb0IQEhPO44kCk
g2jMurT1UG+NEutK2s0RDokE67TBMNymW7lpJOHKyb14OiTn7T7Fg3tH8HSv
9LgBfwCc1yxRGROoTq7AbIea63asNZzS4NydFZBeiAuuSrE5RZ4yEYs8SY3n
KaI6bN1cToMMlK5+O0jqYHFmmZho3Z/TteYpec/YS9Gaph9aTwBPDoZxnLqh
DUJoCfXzqfkoUiydRe7/HWeTVzLytcNf8JdylT/8Q7tV1buLtyEvOVmDAnr7
4iwSz/gN2QOJcpHvRRl74zsn4T5q9f+r0/i6we5ySXrdSZ1zzNZyOZS8z87y
fs2jHXNFmxFMq7XtmxoxRM69cMceLFIo36ZvEZTPzsVcbZdeXBpV4H4ddfsa
hakiLRUyGCvxEtztylM/ZRQb+zXj+v1T1gs4lmFwhhUeAm5slMsEoJ5BtVZm
A+neXi3J5ILIg8uF9DMxwW2zLEpnKWlvjnENHELwE3F+gO23dp9z4v2QukcQ
ntA9+kiMjVeA+5cTE7T5xWAp3WgEM5OaTmCl22dO95K4o6VshTFIEwTNTtbG
K7liR/aILWJOGsEkOaqNDWEKFoQCbZbj3Ad7S1qkxjSO9FIEKp0k5ABFLo9z
f4OL2517xRo2laAQbHa4zNYT7sZyNsF7WJY4IqvkFupP1pvTsau384t+Xuby
300lvRTTGg+pA5uxIW7qwG+VrqQl5dElJQNLyxJGKmffrhMn3BgF8GkRn1LT
c3mc4BSg19krjyM4GLb40rESa3ib0mR/CKL77GWLCHaBNl7Hw50W7hMkx3oa
TUGJl6ALvQcGyxKACctlngqB+/yWWW8aVmFyY5MkCrnJRDKf9bPdYvQ2KJgB
OCbLa3U0cfaWTZF8IryNYVKtPL0BbueeWPiKYbb2AyFosWA4sAGJykZarWyz
oO6uRbre7hPdWeq2pYakno3tekhyj3iNuLHprQKKnU8fucCB1xrx9AHfuH3c
ShHMJctvl4brmcFgkkIJnL8j9IjyOYaSxormV2f+ptNKqPV8jfjqiJ0EY8pF
27Xis9K4/nuJsrSK+eQ27gw/Mh9koGtznpKFQVYtV6uAFxuqN66KN0BRa49g
O3fZ+2/e7Olq8DhlWJICYGrZ/vGKSf0Bws/G5M2Vf0TnKgHwKJs08UTvqqF6
qc5CBbOnfqQMOEmEzPbW/3mKbWMAcVcn1J5tSY5nwgputxoXZaGf5tVWJThi
HXkZ8fNtIEDI+noDyodw9ookvIw0a8zTv4dbvFm7TqtdfqVOO5e022dS45ip
CN6iSSsGb8CbTvLHnTgJi+tOoCNohm39ZGRWXa5G9qUyuGfO6nUicwAZPhhG
qn20D1mk3ER5+n4YcOpnDbs4aMhYDM7tB53spcXRgrbpuLipzPuzxgI+pMPm
PieWKrvAOAlYcHOYLwxDtiH54havaqyt4BtdZchig5DHrbgp2+OJlOVYG3DS
iuGkWvw24fV4KYPTimP7kGWQgzlxake9zJiENLJpd1SpgDdJwLzei622ceN0
JN0480TK/hV5+TkpodDsOhaRk9IzKLJhSdkFc0PLZ4M1hWs9yywICD1p712j
BFSsE8YsA+RLeEc95f2jq6C1IqJqR8y3zr5ri789tM1HhV+PqUKMRw2NQfG3
axC4M22sEJqF291rAvr7GbRIvEjnkwF4q7dj4WpSNXiyuHxaGIa7UD16J/VJ
OZdhNH2iR8jPAdGJzlTilTpt/6aEv0cOrgRI0SHJJEBoFllMOc757MC/zxe8
nW0xNegkXsdAk6bS5j7pZwBi3VMitkHe6l0F2f/FwH/r0yIedWpERAkW5LIc
FKzFFDYXfWPfuxFsLUO3jThiXWhcZNNnsgiCb8qtaRG4wLXGqB7TptEr4f79
Fja0GYCNmgl3XamQsNCj6cW66KkxW44z+d7R1KPBUIOXyneby2vlzz+S9QZj
ljdOLu7Tgq1wPsfCN6VmLGS2Z2soHGzpzmPpbpaCtbKB3aknmkP03KcoV5pH
dKAIIBmT/VJnFBsfjyclksJQFFqNuW8PV26rRIjeTF1xs8goO4wl8BM0H2Cq
wFj8AGOzuZCcSw29iKY3Wk7XgrDUplOxw5vDasKsbeogIGtgsCvDyXCht/vX
gB0bZ5i+ODL1VmFyv+LciKXpSV7hl3uvB5if1KXZXOkJQabsE9eg5ghsmOxu
UE36+VqndUx0NkF0spbwc36lbORKPu29afmvNhYBL2S7HDpGw/Ge1Qlv0p8G
IziTOQMKgq01lcXCX/Kmap9FIiaNJ3V3+E+DeS4G955wPsvLFyGHb8TMyI68
gM+Uvgor/0HunUIc4WoYefFYXTO+U0F3wlM2YGJKPy9pdDLhhdDwiSI4m1Nr
ExYjxCxfFQNG0tN1oFEC9gWgW6M+u/ItY+cT5HctvpDDdPFKV18OGf++unE4
OuUkokswMIlsNsQ3JRl9sxOPOTggZ9C15BKdCAKhDfaFhwC26jydsbCSvPsc
b1elYTkmMMW8ELC6+HvXkEjWWBtgKiUb1jUmr/WouuMVcCGCsKH91Uts7BBF
lTQFo3aoL6/s1Xm54MCa4kjt/OhJIh00ZOm4yRxOfUPffUo8xbhEB8KeEZkD
wDCwAE/eQUBOR+JlpTIeo63vF4pmQ+/ZW3PRZEE81NqW0XcIr/yii4UOQYUK
7URh94lqPcH8X7c1ps2OPB21fFhLNiHrVwnB75pHUVzG3zVsRQUvZJLkwycg
wUBvvhVMrdreYLP1axf9FrAlsgYsYRhYQtBTo5NR/LVG2ZytunsquN/GV5Pn
v/AjZ63J0E3bdIbwc3OO13GWqQ7U4l256W2HqO3qLGRzidXBlTlGIcpQKjUA
Q7+kZPG7lc95LE9mdlzdqwbI3hM7QFbNnc9Gb2VpfMo4jry0gv9+ceDSoTph
cw6N7Hbt+DJ/yI14QS1Gf6oY09iLiX2ee5Tn2GJeZBBTyB7LKT7xirSBgHjH
6hY67VT+D+D592G5ay381w4gIYK5FPI2Uk1CEwKU7COCiEtdsUWrGeH8T6I+
/2rVK+dOAfzE+WG7cEwLhP1s0EIRt6RAkMZ7WXN3BbaepEdRbEulkPufvSfJ
s8lSBjy6k/aT7/elS9nvyW1qgrD1VZTJG+ZI+TNOLI5wDCkxwkiB7wJAvZTj
UZBekCLVvdRltFFEdZXyAw7BP1S8VQhvMxGhCp/q+NrP+d+jKUK1ruPuTfDN
fY8DtHm8uqFbsi4R4JVILOhtikPl12xDfaja+nTgvHvfcHANkyfdNg+YTCNv
oLPWvyVF7V7mrYATP1BlkbawLGib6uwsRWRNQmavcrT1H9PL9OBL78x1D6eK
z7aQcf6iCo2S8YHaegtD0IkrJ6PDoaj6j4Y5hQzD1Zx0yVPUoAVtE4TV5C6T
9YLXDWVBQzpMhxPoVXDWu9v58fVlRnQ1o6OHxoZrEeW0NTbRtHPDk0ocvEWN
dt8ZHmIMtlyHB4zFeigtislwYHB9TCiEwQoHu6Ldx7nuwD+s5lDGy4LI3038
JkHsN9svZSOVlHk8+oexh4QnlxdpF+brdhK/bUaSVwnfBjcUOsamgnmRa2XC
8kMn75gqdGyMTSYoZbq5ly1lMXqO0TBJtce2kaDJD5f7aC0SD8SJDi5v7QcR
uuFUMf2edo7gi5jKvs0BiwB5e9KcaMjS3Qds8ZwjZkbASkZuPpPXzhqEmCcY
xMyG2MPyuE0FqU/ut9Jizqj1lvzAV+0tK1qyn3pJV9Ko/Cgq/ZXiB2mDGkx4
WTDvUGNtdHoJBORHqwbzUc2vCR8Z7wfggIdAeX5XzzXEvCqO0oqmxH+qXPci
Cq0LWRMoM19qLzdjyGN2CRJRhDLRUU6Oe76RGV583L7ZGTh1arV3OPIdVeoU
wLVO3OY9B7Bh0HhCD1PQ3MKY/6GZgEokeFMz1n/u8NfbF4XBHZpeB9+sYLjg
4lS6mtJmCgV1DQ/5vLf3pmTS6bpwn0jMVTpqsSzOvx3tPLx2e7zg7HEvgc6B
18lzSR3S1HcXbsB45milicaY/quGe4uUGk+2PA2UEZHjIkyHGtEazuBrF5av
6l7aNxv6nD4/SXtJjbAjeO5iHl9GNzPNs+RtSLpWzLfcfWVGA7v3GOwJk60g
AJ/iqRVOLajvR67ghAz5I/JgCAP9Ohr7DL1Se/89iPmOrwAzPxyjn4BeO4U6
8Q/3ERPlalJ1TP4Z4mHITUmIZs5IppjeccyRfFqk6rgg2/hb+IKTnheHbc94
96qwe7FLfb8GoZ25K8dLVgJYqzZq8Si1AafXKnQf6TAoMr4+vgytRH4/b91g
sx7/WdovnGVrWe3nQ0+/+wlwvMMNlfADlVsmcsp7lSo79aeF7Cq6xgiC672Y
LRuFVtsP4OhPAJTB7FhSjCegqPAETUlvIkbwHyzHQjytd8j44Zf7Ztjg05iX
s7Ic9ekRc5en0nwxD5swdscujdUzK9HRYG9OnI5XPL7T1gSvUSGxcWZ/QgeV
L2FRAvyZCJAifPr3+G/Cnfp6w7qXRyVSQL+tJEg982PCjMNxO9PgygbULqPs
Xmpoi4D5N8hK04PADGELANAhHUTTPSxG2Z+Wf/vJS3AzQU5Yu1XZBt1qAIhH
+JJnjSDOAWqZfqdJnzHecfifkTV/d+cGBVH3IeKjLSBmt8/pa7djG18nfiqy
0lY03PHrTQAIbkdO+vjSqQt6uVUQ+WYlSBKEskXrpR484Kd4b3YkNqimUIq4
ptZMrylPEYzJqw5hEOXZPFuPcikxZulWtOVcacP7aL8xrCSWb+nIQvPgb8tX
R0nXwfmhjVfEfDGOryDOInsAZOc1o4Jw7S79kR5UgaMNSpOEybGiaQBoDPMl
5tZCaJ6TQPZBxyL6FbCZcdj10frH+IC50j45btqO60OGf/+l/S8b0c9sLzxh
R0hmvaxcH4/Vqi/VER6HUr8Gi+jXTGeUhnJE4qKc+mUn+hhB5QRIgaRd9r54
F2C08Z9TQ74t31PcafjExY8IcABZYnyvkhSuN8BWaeOHXbM0HKx9ccngEfXe
Siri61+yOtz0rC3XxVsS8M9bDTmNQl6AaGDe3Nl/66FRyEG4v+aZz2HTrict
KUYRTfkAAE3tdDAD8fByMeDETq76ACdC4G6AArfcLNyXBwlWfT+HcCByeVOF
UtlcWXRqBSVAinfXKxKZWyvKAgzoILWGDeiS+thleWfVghnnFTd6zWcO3LQd
Ry+rNFGnxbqbTV4Fy+KvkLhUl+RlkjrzZY3Razrn7U9sp5HV4mtVJA1O5xZ9
8clSbXbAy9Zvq0HqgQiuz6iz+ksNFG0aY69MV7i46y+1gfVCcSrbWC2FlRCG
aagQe+m+FLHkjKPQGSPLB5uMPPulBKLHWbr3tMgI0ItHd08Yp6PeBGUejLUf
Rdn2MOh8lfAVdm+W/E5gzfOJe53c8R1kZ6Jpod0XFfO5AHU764wGQyfuzMz9
c2YXmMcRgmQVyGNKJ2TAE7CvCYc2mG11FfU0HWxeflhm2zVoy/l3aiooFG7/
j1r4mUHMhnmOnar+ijEnrVwaWEJrXIrm1nCOi6mB7oXpYpawNj8cAawE8rrr
k0TGxdQQgFxk0bHhSueIR6J9z8eCznGJuFU/ig5xDZvHEN9B6johBX049qPk
bSlh3MTvYhHpPmUcMn65eP6yux7ziN8R+bPv7lgLv+rzw1quXru/QsZN+QnF
KKwRg7IUOTw7GsxF+uYsSPC64zFw9xTM2lWfQo5lSZNS31jvVYaeqdt5Eqxt
uh3JVB3XcysXfT4Eq/0OEciWisR7HhOrKaHrqyg4zjbWT7mXMhvrJzI0OpTl
dK7u+97epxvmNTV6DS5SKp+52xhiAUmvZvoUY7CGI6JCdYqaf+Fz7AP40hzj
t0KFb7q9dZqXb/n94osPU9vRROEk27JYF/V7QYhIFXFlC1NqPZ7lxQXDc9YO
4k5Kc5z79x7TPQUylT+/D80jJTuVGo6fXBThyV2WsvymV9or80UZyyJTmrwy
OcOEa3xCsn0RpjRmJjtE5INxLsIoCwyQbZXerFCS43/MIDrQ6MjP/WRajxTc
FSPjL/5tQjr6K5TVF55kAAuGjVK6Eb9+OyC2UlSpL94PkZHkxFAfCCcEoTIs
fvKox6rFDkqPu5Hy7XAQ7GtBp5Odxr7uzUsLGHZEeglRFSML8X5aEv9f2qKt
9xeZXcZb48gZgLhdCzxfZVAMBfqBnreMWaEDcIgq7ad0wymoIli9DanA5o7g
36BjX3Ck57T+x0txWmJxJloMjCtxwR7V3teIqCNK0mL8WR84cPK78opkWroR
Zs4Be2tu0gsNcuoMlzrWlTVcpWo7TsY7N4UCRUxrDPYFLrmddSt5EHPHf8Kb
i47g/x1lUh5vWt80FbVH+MWibr4q2vrNw3JY2p/vIC14ZIfx0I0fTHpxLqkB
43zk8pKgIOIuHyqu2wNpRUNGn7XQ6r3wbMhpoQbJkUXVcBhhPVPT5m0eYr4X
CRlEiPRyxaKjvot8JaGGywhT8oiaEfclyr7dtCOlmjlLOBKq83LbH712m1vR
+OBW5hOO74m0BGKfa0Q2y8V8QS+XxCWiuyEFezSiaEDhQos5KmJW7iSGQrca
YiT4T10udUtYAikZ2dGUmCEEnE7VHRRoT4FEyAbNRlDnDagyCPExjs8vQ/tP
fargitasaMku4av/nDh1DtdPbyjvz1MDM7iK64BVh2Xczj9zPAOUe/rbYMlh
77bKymhRlNPUJoUMy3xz1zRbcUkyzuqQW3+ukRn1YqD/U4SCVQKEGwn8hwpB
oHnIl17unYlpFflZTYcWggT15ZVKfUuz4xAkb99MZV3FqgfeLtMYBFTIKcEv
Mo7ULs+lHEfrBUu30ah4Mv6XcHmspNMAwi1DEYXKWJyMmYDuRcQU0rEnv1ct
5Nv2zzAy39QnExy4V1AtEjVMan3MeqJ9JhPdKHUuSUx+n6ep3epEdnv+Hle3
mmolFNrV4GcCJruOeN6uK7p0mK1wzsJdsjqYSX+zWeUqzc+iCA4J3yCo5kVi
hGLbqk8bPDdCbx+jPPKCT/xHHqgoZDOtDwSgBn0nASjMxXuWKY6/c/ItfMzz
glGE0m8K99UGZqapvNlvBE299tQ0TJBJWabkfi2QLc0fBAyCMcgHAQHW/LXj
M6Af/wLPA3//JS6rBA1oGcVrIlYr2vWPNWz/JTaKXhpk8pw6kCYHI2iVDqEw
6lmAYrAqfLzpFW0aFr4r8ZHDx5LqUUMNOVPydIE8UA5CccrsMDBBQ9Y+UIPz
IOJcwoXJSUpnQvao9Wzia98/sqbef/ExOlpJmXXXHhycWufOpl4mTBp5QtFT
wtmbR75JzYJIcIcoTntVd6Jeqp2QdpQ1uDe0akKmXUcLxC7Jh0wjkUE4mUht
1PMQMVM15l7egeFRuiogwWAQA+bYZcZ+hdycCnkrf7iKGDC20CMgoXWW3zRP
0xESzTkNcgkczZczPJlofeiKhMITQI8jxee4Btbv66lcgaRF6RD77eMJd4I4
PuPE0e3O9P/OD6eCjmLDv6/JyVYfSnoUQ+7eeiZ7IkCIXMy7cNgQFrL03umc
79sQkxrxdu+B4eoh+NKRjwWjuOmqT2UHNgeybqkOlkH2Hw8grPa0VIoKP4O/
XuI6sa/rk5yXemllloWWEU9m6SwVcxPjVFnllgJhzz6KL4Jt2dF7E1cpOAJB
+X3I0tiPCW9EdTJGW/oykaD1pyEqIVsdounN4Vi7WNn0oJJYH84F6OgbPCb/
kALVMIU1JLGG2Nw3OIjkWoSFxsZC7pYUjTQ/RbQD5G4RE069y0O9LzoUEHUd
6WKy+bWlzB8FuWEdEM7GwwqNV8cyYgRG7mlJy1Lux6XFMoWm3TyGrFA5otYU
Qo67buYyGSWdPf8GD12BGZywZzbNoKoulAFOBswdLtrXcwao3lfJMBUdrab1
1qtMXl2t/lcu15cAPtZO0MgSGe2okZnO56sS2pZ15CYYRTmNazqFQsVJwOUB
ifd67N6TjrPiWUGNqYHTL1eM8WLnkDzN90nBvvIrUHAnsuwoR1TcVmj0tyo4
g6Q/9XXFO9uyxf6cyt3An0cD9VLxdO0j5fBAZ2oENzVQFwYp/Uaa0ERYl3pz
pw6NhYodQAVAbMURKquos2sp8WaauujgbmyLk9r/QpH84ZcuGDz/h64+mENQ
PK8U/GKg5UqRr8GEDLhH2bUZQDXwYXyJGmwz+zI0GTq9XloYU9k3wjZWvHu3
JK3p4+qukcYCXCpcpnPrqo2MYpwjMs97gjfg280pr3y0fiAyzAElKu/V8SsW
DZZHGNcpJFg1AU0Wa5Fe+QJikm2MWi1RPEiwlVcvbCRKQjqokK1mSJwKIUbG
f8koU1cp1rqkHj6CgVKNedrYLykiQ+7oY/rPihj6oWU8VG/gXdEzFbGpuyst
qOB5J64JrQKNGZSaWYHbSWyx5KHMapWl+D94Qn60XX9LugMcrT/aIEF2zXlN
eE3LVd5Z5S4zw1dGqvTU8fl5TosnA+SJ059nDSGV8gLJxO/kBz8OP1ZfsJjA
QYGG0FLIypHiWhCSPMNkSo9Y0IyCwvAWuTqN4ULKE4NRDiUgwcPPudXaJv2o
MbSbY6Rv45hC7TlAvPwpUNOm0VPI20OgtS+X8HI2rLsuvfdhX4tNXCDfr4NJ
Ms1yTXmn7bvQLlnGfKWuGAOgJQq2ifEv24bhgY1xMLKJRAVdrbXlsLd2zctN
F5GX5Ip5LqGo89p7C8XJmkyaQcYqIcQueIzUhzusPjY3REjgFAb8jQ5iX6RS
gcbMom02TZb+ctd95+VULFEntzD48STCdh4zvTv2358VAW5J9y9whMhintrn
ZdgloE+1xKVAN/rovH0gz4nQqcXSlKh/aLOAS9PfaFFJIfMhJ6IHZa/unlLA
nD/dQiPSKBM2Z0Hnr82qVofg/evOglMwjD/TIPKKOceo23k7x6VVMDO2539d
72JZ7jaZtInWH/3m6Eci6j+L0kA2xnqNTeWGx5f3t6cl05jfmvoaCv7/CK1k
QSphdM8X+UXXQ0EIaZ4LlRH/rhwl5MFP8JsbCXwd2jX+xqW0UbRe4z+NJNKi
3y7cJqWiZIROROWjozDnH7rKsItthGrULG4UpSyHu9A0LjdOp6WWYTokiMsl
8LrGoP/xCCJv9LIhVOKheYuVY8agDq0Lm/5g/P62sVvi27ynaEJ+b72Mc/2M
jouNFdLPeQrE9Tu9awG44VvTofUBivBly6psAQ388o/BGXU6V+YBQ44qi6L3
AEA5DDyn8WXEmHxS2JQBc1JcrsYFSCaI0NKMwO5h1/mTXDCq7EQG6CVMWyBJ
MQzZHh1UXLOke9l18y39m5T2lD9tqttkIomT38RxaIEZLjgxzUycm/UijLJD
RmvqyHUSZNVS0guxfpQ5ydXJeJ9ahb+o2Y4TfTzS6lT8FlfGF80DX/Cr+COg
K6+g3jBc4Db+xSS+2peECEzfAiuPhbGQthafiUT2WWxievTDMAjsp7QIce6I
CGKbMS7IUe51F9x+elNpu0PjO8AoE9u7+Ghm2K6CUYoJsYVH89cTJCjxS1+e
D6LNTZPdKjn2ZBAfx6epFp7okiszJu6t3RZpBPoIniF97t2RlqEIs21XN92l
DJieLNyCDAil3O8JUp8jOgMvl28dIioZoQ/mDLcedW8eEa8LKmPxPeIiRL0J
Q0802Ze+j0NisCOPLPCsxztq/Lj4KLrW5cAZYMipZGcABmyBLEH1fjD+Pmur
FbNEMyBkoI7zJQ4A/J4HGtelMcSFcUFWMRp1fHPwhbed1ypFeNZRyonbMU0K
mvuf8Q6fPivucDgtY5PqG7LePMinUOHGAdjAVUPXgxSACIqp5FacBm+HEZ7n
RfcBArfokgKWhhJfh7UVAtA9DbiougxLmmG0lquQWf7FLMXB5XFqSrxjIRpc
3FjwIA3s5YyGy6wyj6DYuagonqxShvXH18woXj9FBHQQeCnMHLHe2c5pTzzs
IANA67e4KZlV62C0r54V23rysxxkvLtaVUOooZY2G7ULukGmdEtW4lwlu1Gu
u9mYBT3BrRSWOYe6IYRtU6wvY4mrjSgNrwzXzL+V1pyHGpbtIM747Gi3F52C
bLi25DDQuw9QQu/yrH+yadq1u1nPMTR4+Tik60L3w06o/XljNue+w/C3fml2
z2AGi1i11qktQeRSraaFJd5I3szIwk9u2OyrqDZJyk7R8NWoduN96HMfr8bQ
tvr1unD5TUWgjZoQ3qrA6bIffG7XBpGPZggI9cA/ew+efIoKCbFvgzfos4y4
fOJNZWgZOpSWFE4+anh5cJYuNF12afjDs0SAxjH5VhtUjafrkIPHv23uxVSu
nROAiXler4IpqWglp5bTBDFPcC1wHTgDar719T0RWsuJHIi2ac+NgYrxBQE9
QuSxHuWqvTXsHG1ajPzeu9gqWUy+JNCZTafOml8Ag3Cu+RKgyHcoJK91FyCK
PrfCkkMChQHiGNTwZ+YTHSWa9/4pMVl3uGO9PFBiWib6/uNIxhb3ewjOnjvV
W2OoagDnILC+rFFTKrEaA0PX5fchwr1d4Hh31JO7/mzIgJaIoXFc+JjZePa0
O5aAJ6+MMkRIbwBgH7D9o599g9nfa9lAiJCoz7OJeBHBYdnvvO3rr6U2G4p3
4LwX+KIZSjGWfkp8WU3JV0cUpiK2/kLXLZSUuUIGzYmhPKJXnmIUsrus6mFM
Xi1QFEIkH0eb0mmXOd+s791TrDEE3sggyXX8UpgMateXYifX7BUT7qYvkhLQ
rf9c1QV3UzcX3geuOyNvsCWruYN5vwoOUw/j7ks5SMVfW9d4iEEtG0mIK4kA
qI4WDVg83krZGTKtqI6T4GGBwg665dlY6IeAz5xdJkvXAh24iYTb1jKDdmF5
NxjZ6SYQZiQOe5ot0Oiy7abWch3LjPiJGhB8uuQXjbpd1o5/RiqQicgtRaRi
mFAmbl5yUCPlgDm2aKoijjGqKSkNLvS3pcQPmKBHeYaQ6rcpVGe0FA62FM4L
gvXiY7n2/1bDRtQWTSYZEmG/oyBUxhGK4MmzXJ45RvRWx+Y9qSgJi3sHhVd2
WkLxRFMD8hIVQi/N9UAXzEhb2NyoAEJ4IZw9sgpD6aWsNKD+RnmhnweNa5Wu
dmmEuoYPyNpLqkKTbdVWDw5RfOgwvtJ8Q1v0I8MLDjVAA2zuxl2kmaIpCbBs
aIfFyU9ckOm84oYurGNQCL1KGx5EDGvMo+d7aFTHJFdGWl9+DScerdyUyTSr
7pyCEjD4BccY09prPSI/aBAWfGaEjw7Umxi6aF2DF9A9E9hzi8nfQ194+/J4
JMyhQ9LBwxM5htZ8adQRZgQ4ckaPtjV3c3owt05A+Q9GrPHTA9mTCIFBaRVi
200GQVGp0osT5FlvXKiSw9311AiYfc4agt6nWPVunspuUNnZxQsDiCOuU310
YDK7v2or7YKYNSRbrETTWipphIVlnjzrP1vPIlEzIUJ6KrRScjp5qOQazf0V
5Fm2cbi4f6zbG77qUPq0g0xTyq29S5r+DNO+yZfsUcv+p7mT/m8mXZ8+1eaw
Fi5Rg+crsqhCf3TL7u/sDOSrWnngHauRJ1zZNBCUI1VVN78AA7rjmyeohTgX
xjnNoqYJyBbjjrUAHmBUe7PghunKerruziEUbWrAMRUVogOG+GW9m8X8mVwd
AgNx159UZ1TQHc9ZXRgm453qI5dwLYnPINwyL7xS0a6V57q9lhwwYc6lLdeZ
dQTdzwj6zn6fkZjFj3NDTGRbfiRXORmJ+fImZP2rtv0rbO01gzOtb9wqatz/
uW4buMKsICZ+XPwKdRGryGQyRB6gYcj/0t+v65j4nRaDaqIlewfr7GFwvRIz
P+ZyOupWeVI3qHp+2NK/RzymPjOZGSmn0ufO7MSB6ZZk/as+bfvFq0+xTg1A
+6ewRQtc/auJVwro67rZxc6QbbxtAXcJwmVLaUYBESjI+YR8Ek0IG/OgDNUf
H8RIKpCJc33NH5UENAP1IeNSPcS0/UoaWLP/XrtGGTz62t31sjmkxbRvnZ/q
/7aKShFbYiCdX8/zqkKw6ExnCcuWAq0kqi/lwv/e1b/gtPTG+tcapJ9cy5Hn
9FwrlRVmXTx5U1W/gCWANahs2kIb+q4NVe6YO2lqCjtIln082i+Njgp1WPi+
AdngA6S4zYpvWbu8/87OzZ79SStVxF3ZYRlqsSQoFzIEENj9S+Nq3mSS9Dw+
3dtsNSw8nVzQtL2gMUHqOCuku/S6w4spDb/o0wJ6jDlj3fczm6ct67wUHYiB
l3frH1BcsIxXkFKQlk2cHURyjo3iy0mpOy9KL5OvcoHoGsrrxy79tyvAE7S5
UOc8zmH2d3NHDcANq45eJy1AjRVVAz6gdXaXag0dDAy9NHqjPHKWSHALMHIe
U2C4txoR+aNjRmYLF5Rag2qzWP34cnJeiXaKASTt0+93yaQCTzta6sGdxm+4
2eFpFkbliRRAdGSpzbdAGCJ7NWT4CEIN7z1jAB5Zf91ixlpFGVOWrA3WDpYu
IzsGQukffrJVsOmqDsBR1rhDs1PTdpM47eUarza1LQFWpOI2FCqgWM8LEddW
+9n1/iRPfEoeiIPm0oaPmb+wlVo5QWrOu3m//G8pntPimSyRMM/AdmDiHmwe
GY3M0NrWp8o1CdgPU8E4xuI3E/sd7sMxZ/0O61YjoImr11WTy4Zz6hwj8prN
yQMzPz463t0xxUMwg2o4LLM3XWnsEqckAavkGCS0jhIZNybwzhFtYvenRvip
7I/4f6mRQaWatL7oms069z+lPq8ALo+TNCZh1dlk13LhSj1MDPDpnHl6nhDK
QdEU9UK/6XU4m7WfuZ2coJTN5Mtuw/JFf3uA6A14uAPXaNKjsC2c2CQebPo3
puxH9XqN6iQrSLlIRlGwdoMO1Z/rqHQxFHO+Ce8ity855pY6AG67tE+9hbKi
K3RNnWOWyoFf/znLwi84OShkJ8vEdUJ2FGKyfXXC1+a8Ajn+aKWzCui8ZOVv
NraRdbIA/F22Q4v/cO8AFT/gP7+9XPGJbr66yJhcJlhfyq91i0rXfHfLti+b
PEgiJZraCpM5ygjMv7Mim8do27hOndr4N0T02Ec3qLsPho0E12xjkbzE1Gwh
h7yogWQljyeoRJ5LhT5Px1mW/P1nqMrFXHU3WCGJYzngRufh3DCRKeRvbqpm
ZMe12I0q9hz0lom/dN4SCuPSG1sitGowYaQ1j7PwJaUO0f2sDCjsNWUXYiii
jvBoI+Rf+Ps6prjxuoqzZDQ85pKG9MDf0/Y+S1W9LpPqwZDgz34IgAj/pAtX
LEnHojy3r5Jx+RzDcCjleHCx8LujWUDAeHhRmWA40hXRYR7OHqv405xiXa6a
JPXy0vf0GpVCm/W8B2VeHESVwJntCfsEsjbwQZdhXxMxbrmDChNRP0BlegQZ
GIw5BkBVt+QFYOVgbPisGIOn7XqJbu4hhJ6x089FK2SIkZCq758hieC35Rfk
ql7zdPJw8LVZr+5GeM+3kITF+O3chd6UoSaLiOWDg6Xnadqwwt0LMhG9aamS
UWa8eX/WBTisHpKGFfgEJTYU2e9X3Em90GxCl9HYyuh4YjZCo1+GUr40UL8D
/E7d+w0W3i4UySm/GVpoRZRS1u3O5ZtZCwFAp5RwbEyxOv7AHRk/IYnFY2vC
7XcxOgQj9h0UQ6i5eaTtxWvVfVxVMJmwE41lOquWbTI9/XCCRrSZvynmy9W4
164Ipe4Ju6L9/Ugrx6M04zogEI1lXCuT956XO8cuHW4kNWEiJskwOH4vyxpi
rw5FHL/EgNKwB5oW53Q8aPu9/0uXLF6elhIsD7VIgAFEb8adHRDylApS1g8q
yU4WL9cPdxo1uX0NUCLgcbNUELgwa9M1MEHrorB9gL7ZZL9IrW6MmrYG6YqU
j+J4HmU/RgtvoMLaK+D5ZQyoFLmDDezJQw7XD1tin+Z91vcrNaC5/fnG5skg
zlX1t0cwkD2clxYvgpMbRh+ZW5wAPJiDQSQUL/ORRFQPG89bdAIoMnu81uIW
Lj/1ySuo7S+ZrgMBb12fnpbSlHrqheKVnsxBloctbnSZy/R83aXLI9wqaqKh
Um9c0mNVfJhIns4gdssBDsu8SXrgHmNJgwGfa/8RvNrf2HTAgvi2igBMDVmB
emPBzEsnjNRVfyG3jnvOHAjlDwShBG70fxO1+su2ygBuu3NXW9aB9IC/c8uI
mUS4xJA9XWWREfaimXBI4+7cuD+PGdcwNXIl8R9+3dcmbCaWBAS4vavM7LoM
L5iM4k1F/YzNuID+y5ONlU6NpDXLK/A+D4ghw3phDyvA5QlwuWZF5KPXUzPS
h9NE84c1pXuNb6c5bXzo9vlokPweTW249+J3IKmbcJC1EuK1MAzmx5kcT1Vn
juWEmRHk1dTEofVq7r3PUFG9Hf286/h+sMCNJecQX+TBVyy/XRUNxKsGUWMP
1sspqHhLSP7PwML8wmG+h3Dzyw2SilhhYWrj3B/GO4Jo0FXvPPF9MLSUwYds
DPpEo5TTo6qS6pP4mukr7aNLQH5di39eFpgrsb04iILTUyvuq+i3vkp3ldwE
ty79uoHrgWV/DLqF5WsozHJKG6wiq3ZwVIquKnol5rhdIF5J3SL6V6nnBY9j
RTi+OTDgizsHxnQFqEw2hfj2zgJ8TLfb9DjZmsgjckJyZpNvb6L+QLvXsJWG
RcSpLQyFCNNxCm0JzJkK1gSQqNn/r+hvRqFklHR8YIb1uH8fgbbMW+RtUVic
J69w9QJZnznGtBq/nVrhRKrkyQt9fBFREm35SVSHRzKjpvUKXz0/fUix8Ghq
AOygpRGeVei/5IXYWe7bvUPJ6Gysj5moFNiU3TyKJx1R4483HD9L4O6GIDs7
2IFUxfezE7O/l0ukXMJLfvha8sOShXLCWEIWj53KIZOMLLYM4G/ARenGrq0L
6tqcitJZzNCIYTTRsk06etHGs9u4w965/Ae3Duodk5ZS8UztuVMbT0VOWoJ3
Tn5NUZ/KgJRpxEZn468oE78+ZwifHzanPltfhWQBU6sgt+3jntVeU+CIIBZ2
v0YXi5ZThLVP6mG1IuRHq2eHvJaB30yZw7NZjHYyXoojb0rlmZ8Q0pjG6eKD
YUpXFyjAKe9s7NgbIYUi3+J5hM5yqtsoJEle68ckHB6uH2rryOaQ/gQpe02v
R6GmiAO8DRkDXnm3PsTVjJXfheEvFESuPQHLU/ZY3jxUi8aG43lS3sYLRX1C
LFXcvbdRliDZDjgVjmVGHQnHHtQB2+MQLcMrB7s7108/qB0UaZrlrIWPLdpN
F6XIAKJFtRmCvA8gKi6op6yxY4gZcmWwMjZW/Ojng+Sy0Ac4iJ8HFtbmTT3l
1An709M90+iQiGVo3K3E3dFvTbWpEoKsAwt/q9OZjz1+Mycsoxti99619oGK
tHQQ65b/iGE6oWSIESwHnMXA2MZ8raBTde/79UsKO4Y+o6LILH04awDPRXaJ
Cd50MANFsALvtQkmPBTmVcY4Gv5nXbHka1Mz/R78tqrodSOYRyXbEtyBJici
qbyBI9GaFJK+6eQGovnqyHDxxU5XufKywDjyAJUpBZDVzabz5mHky3hYeZyd
NBfruDWpd3T+7AmlOCGcMGEeMQoXQNSZ4qRrxS3L7hQt4JJqVOoWiA8ar+N2
OIK2k5bSp4GRWdnFpCE142MmwBDzF6K/+RLxzvnTfWZcNOsS6qPVpK8RCYgt
LEIuXi8SS06PeaBvpap6/hHFE8XhJdhTZgmKYcdlj0JfQVtPAzRDlmxkY0q8
dW4KOSw4t89tKTKt/ojMRruU7wZH5S32UJRoQZfpmIC9B70cHnSQ6WJnDVyW
Pujzt9kfQv9+O38kMCSTMvphQkWqbwn5VLGxO8PGmVJaJd1qWLcW+7vrZ0QZ
RYE0PRQvOV/4t+9oHqm5/niwmSjUncl8eP/M0r3cyeV0ne8Dds6ZNjEHWzCg
HxcewXBnheoli3nlDIO9lWFSpkpHD23e+7oBSSGUT4d0Rbf9EzWF000VeHqF
uAuUBlIsmbF4YBLO4rFOJfSaSCnoEOjlr1WBKwmAdfiNGLb3imOJX9O3vTYA
ID4cdDxI7AE2dZWtQCx2DFM+2+1mf8Iy7XHKmb/7FQQgLrFVVXNoVMEqieNV
fZmHh0Db4Gqnnej42yIiUbv+Kj0l5qzRNvD4V+gGVxBeM6M+0qw73Xpox+9f
/+bNPb6dPrZdfahGxJ+PvVik4VcUYth1gskFScxyQ0fN16DITSIA98k5Pdbu
zTMg3+6YIdWM/z203xhLp3Pg6BfImOYhBAeZXaXx0md6x/fvEkX+wtJ+MjfZ
O9QKVATXQB+CxBDUphzWjYbrvwadF91om7ptpkQrxmRYIlDSUUZIcVsE7cMK
q3smZzf0GmDHGYz08xARSEAj5wqx848pCMVd2J94RrLCq/3SLqFB3WYf/c04
SX1nswbKETPeRFqVL8eyN66QBqCbhuMOx60cKH0Uq8MdPOSe7Si6BDbDWJjt
+RAk8rqg1dKnfqNUDo0X/Z/kbMSjq3barX8+zel0yF5ZeT/vAst4gkSYDYWK
20ItOHDifgbv6a2g6uvcfZJ756vNCg4SX7ZZjO4peufsvS9S2MzNsiYIrOYV
j+VWQST6Db7h2NefUFsv3sK0NCDZsAQJ6mPiPMlIUjtlJZce7m9hye5j9dDl
2c2ZClnY2hbq8aX7wRJQ9P21yniGD9slEAd1R6Zb7zUGotCcB6GBlzGad76x
vV1QDo1AUOT5jKJfxzzjgmDPILytNYkQCzE/HhbFtqRsD3CSiAFiCRK/oa0B
6OoCgv/7NBX5ii8BBkqoaOK9EZ4htUc0OySmMURszNwScgpL+FV3zHrMR8Oe
TselRgJ2rEyMgPH6M3m7Sc2Wo5VJlCMba0AaKdZXg2TgHvylys6HsxewATg9
LZCEwusNnr8fwbdWCbedi5YJ384YmA+elwqLNvT+Vu9XMgx95U1z3VLEFooO
fLq7N6XbfckHw63DjGxAQNkTpQq1sXBuWqJT/ZN3RQNXxYEfkyHbuEyxtdUP
3xXwUVXVdWykQIFUwvnSUe76GSZPDLWke85jqtgOZSG1bZ5wwwdXtqYoMnbV
LQiWV+EtC5NyCs31mD6BOgNs0fUqGeQVSl1v+mHGpph3zyeVPmty/5cUj2DF
8U+F/wmvLfNZS1Q91hLP8ChRcMomt9UZn8+ZQV/Q3og4Bx1nCZvTm3nHlHjU
ClK9+4QZmsnWH7g1zX0Kwfa5yxxUZMu1RZ9C7rLhzwc+ZhvOxNopY4nkb4KO
l3GQvU4WFLg0Tlxq5OJOmEmDi0iVp/4jKrWQoYpk7AbsMlTJ1f3PeVphjKWQ
HcMdCIWl7nizrjywHox/W7k8y09K8S8wqTiY36jFb5mdOAvK+3bdlJYVM9rz
cT63RgxhWW971X8RRYnhaymAvq/fk1TW5lFPg7ME4LLh311ZtfEuvQg5sgY4
pSgspvJ1T7OliDBy0e1rzCjedt/1R9V5Y12mwNKFzl+Hk8j6x5xvIiUt2fe4
TfSHN/9SXxyxq3iS7H1Zb/8hwW/t4JfVbcpib0N3SGmyL06NfYIcq2MUq5OW
FaKo1xsW0ubggvPOR3oHJ5DWRwGCHzr+LMA8QdSSntrxkPssBIcaQyV6d4gg
TbCC+uQPhntVjjB4GxQ+IsL4ZXpy9SVnwVWpRCTaBqg7EEeabLNEp1oqqMZD
XCSxLAso053d1STaCnb6n5K9wpc+xRFyHUK9x9x8h0AEzT8aGKgCJh94wToy
denM9/kxVugkDZKCP6HzzGpxRtfvfp+ckEj0ctQi/h5obb+VhaRF9HE9gzPl
E2TxJBiqUWqo0cFSSHV6/NFTbTBECc9Zll9+reKG54WW6yL/93Q0eFBkHpJB
4jyH2t1rWiCTaYrTwVlKccKHOX7cbQlP8agRMs0r8IRIXubjETVa+HkLPgSQ
uUsz450oBv+wrBoeqGRLrer8zNRSFW8xcJCbFqel/sfl0W/mC/X0/3C5pIfy
SrxzQycJ95vzKunbzAukqQd70JTI1P7fCjGjVu7bjM1Jsf3yHOICqRwxg0+7
oG5l5mXDTNbJ2YWmFtMbatBkuV/IOx3s19xL/24qc4bwGEzD/aHcE7ngSshI
RVLLFurY++KbYIGuD/DgsI4qPu4p9sVAk58ihaUMDdLC09H2SgdagRvpPiyK
d9p4DbRMMmwOkkQSlXINETl4UhDXGbAJWLaLdPx/QFeRxDOiyHFl9AFJMA0J
Cld2sWRRMjcYYSfkWQ4jA1oYQSykZSGuv0RyUPcIuiUHmXcncBDl7wwI/IXD
ofRnA5MvKgRlaTsNH3gnxCeiCP3kNPqP8HR9WD5Q/e1KwFieQUTefH7DJ/Jh
/t5qw4/xbgMtfd0ZmnwK87CIvXeUrMHTC3kjzJyKvnmykxSfHHDyFw8cQCIh
KOqFy7uvfHpbts8yt7DVQZA4mvUNJGayGVcGcZVsujP7iMLmrmRyyASoPgT3
HMyv7vJNxLaaxwrbGr4RamSTmCuuqQI+7z9fTKw1ZWj9YBTmt0jUcqxgO6PJ
EgEmC7msIFBDSlKlx1vqMcFBxkeOdjq05QU5Y5gscO6mLgd30LnMOo2xplng
VbJ1OCicvLY/6Eq5ttMwfH/CJdEX+ar28LMBJ43mqG3RK38FgxoAAw4lSusR
JNFuJDekTcDGXcpaDoj2oy0a9eW6BgDldPPZupnTNkXwJ/w/xFNbQx0gWg02
aj/yLbzz0+W6pmYUlD3hu3hBiQSwz+MbSNNEDADZRYPjFpe7WhRlDVp7EXXt
EgKYpCVBy7K4ylGvnWOls3okRPcvZAeI9nKfMSRvXtf4ue/EmpuvpuuVeQyU
fkXI5BS7vBluVlV4wAk7kcV9LTfDVcNMgbrZPGOBm8nGR2JhAxRa7SX8XdgP
AS0YPjM5DH7ZJYTD2NyU0meK6Mu+wC/ysf/L5sNxWX1PPcSoEeHSRSDlh+JA
vCFwXGg4b+uPEBlE2/kFyGyL3PDMpLygbnNhKCwspcqNpWNP46fqb+kb5Lg3
vXjpAVpxYHFyCguU0AqfO6UfTw2SLL3LB82Ey80JqXGYKO3OBj1HmS+8dGQM
l68ozJIKzRVZE5h9FC5H2dtFobcQ+1gsNMqcTN8K/xyhOdXL0w6o1eRRL1Dd
D796xJiJt7VkRpFbrwa1Euh1mmcgRH0CQh5eTzpEwX4KtEbJ5cCSFA8JQjEv
0gUoWZAXe1YjUNsLjpe8uW1omQYhhxNey7Qlk/+vyIixz3Aw6puiCCy3s+rP
IGk969ydgEywPWWwfWDN5AJk/uazcf5zNEDonV0WqwTbAljrpgmkeN2uRlol
c99jApGr6GpgArjFFmZiP2+MOkC6fs3iE/+IkizI/KpMuTOj7v1nXSgA9lMD
kvqP4NWztr8IUq6+BVPDDsEOZ+Tj+T+mjF4W2iWMItaKfmV4TqnHk7cohRAT
r6XsfaLOpDRYGqM00MKEHJVfcmxlKXVYGEuwyem9LslK3qvRGlMUiIoJ4swS
uw0RksO1PCFn0VWNgEOcGCC5ghiMGEgpyyZ44yfNkXULWS7YHCyGogE9bON0
SyBpwxg84YKuEJcKEGF+8YH7GppnNnL0TId/xG4F4eAr4W7JmtUoDzepiXKf
EqEODS8cIn5rDNTGt7ukK1vuEkUuyIB4tEDAZH+gh4hD/72wxuYRr8eV6J01
RHNWwTM9f/IoCrlCsAsP1qXd4r4YF/2eb1TnO6kQmmMU5J9RMfRju4IqOCvp
y8xsD92JR7serHtIi3m+PbeE29fq+MXZSOK+h9tRrhSksa3hcAkVqtfs5US4
kTroBUklcfyPkuBBBlKk+Swjep5Ha7FmyLTew14yJwakZTbtij+sLC/HVN0P
ijL65YX1lfvoHhQdfPp4a+02n3SAWvWQEBMInQ7k7jA0vcqtx2nxhWLxCczJ
tB67pKkM3nkQe7TGceESQiY8G0f99ZB8ZdjGmxI24WPEggFm37SV/GKud9Gc
c51D9RAivy9klaMYzIqZBOOt3pV7rYGCYAmJSjFuopyxi1LWC3UpfJVVTAc1
XNbzv4nrq5IS+mRSn5wGomwHJpebynJActUv1jkBGATXGLnfsZVRRcu87AyC
VOtqgtKz15ykx2UqNnjuvJ2br84HMT921SzYPg9jWcLBMyjqEsAMIsTKW0bx
2qGUWB/zN5JcURIAmTPgN/gNRVa9dnd9o7WhBCwpJJ14sDS7k3z7lt77QYQA
vkFaxuQ/aPqtYt9LykYmdFEzecMIN+EjadNSbAQcZcFzLy6BNIPR1f7qMKes
83vPqkSz01cDl2Su15B1soJJWDxRpl5apkorAt4bKLFanae2UtfvA6LMyiae
Sm632HKpyv/hlkAh+iNokcM2mAK1docc3ft2FC9XlAtkYK7RRfYCU0UB6lRt
ynvMDm+j98xKObuGI9sGqKxZPIaX3q7q26zMhA7heHEz1IDXphMsfMtdDAN5
HwZzmKgxAlJ1+64kI4DtL6lIQvvT+RcmEHAMuWVPTpuOwi6cBzf/mdP1tRDz
+DTeHzmFtEoO212ofgrbOG1HfygYDJf3fG3C7M8GT3kPYN4WOeMJ+VcH4Rzh
EepRMVJp9qVb5mYOO6NvRrOzFktEc0qV5M4fI4+bh6JpeuP5jguYLWfmTlcC
Z/WX4ompLvIQXyoLnCJSU8dMfHAWYt6TAJKaBMFI8LEkDERLi5AYSSFvPwjG
ZePTWBXI6YXasNeegDlzBW231RxyqhA5xolaw8+DbsDBcxwTl42I046kuQrN
rjGr994Fnf5dGNzuJ3cURsEF8vbPtBizHmXy9IB5+T6yNisNFc8ZtlLSCldq
Ud4aVzrCMsYb7lRjrbv5f1wR0zcLRJ3YMdIpiLAZLpbotns0CtAti68qSvjc
JAiEoYnIRhqvciq6RG/u+stDWzjsR3IrfF+AOhKQSKp/SVgHvgOEaWKwQ3CP
ekMrEfIna4ajx8RbA9mCxlN6flsZbid5qnajd5h5RLKhwsujh9Jk07kDw8SH
/mvh053dkvbU0N3RR3RMbLwFK7124pnib85olJZdwFKbXgKZpKNARiyH6bgy
tiaYCQmWtZVrdULOpWPbZZbm6gz5B0lK5xhaGKJOaxMcgP1joHxq2D0Qg5ip
g9dBrWtNN+i13Telxm54PYeV9VaCLrl3MV16sda9zaT+Y4gWHBZ6jeCLoEDt
de81cLtOuYQFwzmgJ+kp/Mlb3zv6vnoLGILJQjr2teqSL6TpMKnByyd2gPJj
Cb2W+uSvJJenyVkYyjPhLgkzZ8a17d6wu+07OxwxNCswulJELfrmSudYaSha
4mOU2xlOHJkE/WjlTtCjmDU4RxhFKAnSLngWHt25uN1vDf3AlW5PpQPRPNdF
jfmHSi488YHHgia5kSeyoOevFUfe92j3IGHZeL6zLwePut4G8jr4U4nQJDtF
DN5gJDe0AjXg9Q5JjZVpEkaYut4NbLsVUh4ymdwkaQkmATtr527czEghqkqr
+0Aidn0MKZ2uR4sC2E7/24fZcCK6AWLQDw5QrSej6gjY2MwF0q9eivSkZlcd
78+dzrNrqtmg8xMYzAaERRqTg2lM0txmIvkn3rpolMI9fhcqx/CjZhOFcW2b
ecN7AEs4Bl3yxFVvOJIrd1ZDPvCtYSQtHoQxJCTT6dcu+GU3Qg7RjAbA0sqc
6y6Xm3gka6CmNo6LTwplEFHGwxIXNe+OHwNudXjEWxuZPHCaPbcAtTpo7ty5
TvRzFGr1ZE978TdY2jSH9E7KGaq6iF0ZbxKIfUrhCbtkYyaLC7esSkR9ED5W
ZD2YDDNtkmbGHZClga7omAWkiiSblq8MSI58TEzTzA64j47z45UgC6RSM2//
CnNnMP75BBfhby/Gw9wZTeSG5ihks7GkGFvueppROZB5ANB1CMRnzeknBH9f
J4jeTLPABt41eTRe0IpevRNGv8bloF3TrPT79CG5+R62wxa2knYUMlttQZ1W
eU1RftYOEyLQXRvnKh90YqfAoOFreibr4GTwRHaM2UjhXySbC/R188n0rK7p
aCXZKQtSYAD3c3Al3+uzLaQydjvzaaizoSte7fU9LXgUcqw0KNxX8mZ7Hge8
k77bqcS2v1cSPTNjUVOCZOXF986Jwjg6GrezN4kBjEyeQJ2Tcgopxzq173rG
vcog0LHXWXJDlzA9hZu+Jmhso3FK/n1EwDg41UIvBVE/zxJUYHqsNUxKRKy7
g3jY0CXLP01B9nN9U8gz7/ZlL2wFtq47vlMhz8XiYw9le6jG9Q0dh+4BfC8x
VNKnmK1p7dVaunY+3uHGP+3GIsg3VQHuxAagvIqiSpljIFiyxYV/Amr0EHeP
GjzjCnJGZ9dmAvzWeiZUjmx3Q9E5TqejvaYPnzEsx4YY3/rVb+D7fWm1ANCW
a4sd2a8ehuc1eepbiSpOgWBbUP7aypkieTV9FJrSAy9oHl8p31yA/c61w7/x
IwiNAFaG8tP/sJ3vm/Xh11pjXdh9z/36pQv4BkCp7DgqzlIny+B5+IV/P5io
2Y/gCJIe8rJ1KWj+OTmcjm4qmqkc+5P7JdEZCKBys7pQbDlKyuDT+YzJvzpL
XtWMdfbDWQAzf1Ivvu+FkKFhC11ETPCi5SmBdp3dORKp5aQTXuMZM19heB5k
6ifKP1zRZ+REy74QNh3YSlQMLgXujOyzkKMe7+ZltflDvRWNKlBb83+YpJhc
H6/qk8U8EPx/z/CXJe1xwrhw2TWYzIfehzjK/Vo2UMNMiG5jpJqRtZH77xeb
R3Tmk/0RlMdbRN78w5HNagokx8xO0D98hTOxE0zQDwiMvcM66hFhilT6qr34
8wf4JWwzeHvRDQCc3V/sigS5tN8HI8D6tm/z3dC/KCPHP7PsTpSfDuvOJATN
9veWtucMhCCHssVcdwh/k4OmoxdguZfoAYHCpN7cOtr2BOCGLVzWzeTl2c0l
12jzjrxTwkqadNV5E6VEsY34madhTe2PhBAv9WpjG0NKoFZHeTx8IYc1wQ38
6NxzZDfdiqtXuptPz1yEJ9uGlXUfrFvnMYK24KZf5fxUGPb9e+cdy9CnDGY7
ezb5Bhdoyeog/2k0fNLtTycFHek+YtTxgobRau/WSnkJUji2XYK4Fypbus87
GGsXstpPQ/4thfCdWGsGkF6mWzLqvwnr9C2xnsqOoasiTydiPNsLywsdKc3b
e5bCtFBsOIEcON6ft05U8dhvVv7RcvlH/idzhM/TqqQPdSlfBwhN2KdrZjCe
wYWbZznf15H8uq0iq2AU6lVVezyltS/9mcgFnBHbVOFST3HI6YOtVzkjN5bF
b2qOZkzVeXsmw+VC9x/nZDmQtXnLNnXKO3lGH2ieznCaA6m8cW8RQj77dLE5
rxkg4LWBfwQTgweRFqXvbDwP7mkO/xUSzBq6snmGC+2x570QUEnNxslbfBBj
LtMCJ5t9mcZ/7KzjsIYekejIynm3sad5h0+OtxdN6gmH/GQ7e2CPOMJUwbpl
+u8dN0a3DMLP7m1dN3B863mfPHkPAQ+8REGISDfOnr0fbr92qGXT/8xCH2hW
YhIV0OH9mEe75PbnphKiChyMtFhdginmDRtmo9k+/XN6fo08ZzEtpPhooiVN
UxNB2XiVyyKO41dkMCHboO9LmGz963uCuq0NQa4ir+SEsleTsmfPxfQdj2XX
wcu4WhBx0oX7M5pL1ubVsRlCIZ3ie1177UmTU/mgKZj/H4b/DF3l5rPcU4Jo
26aTcrQm2/tHmxB7J/v+zbVGwsEDmr/3jvIdg97lzzVYTTuUkIQaqXVZFntE
t52wROMCmcNz5gTpdhZ0v05suOvQwflQTd3YRbX06mrHBUJvbSa7wB3keXe/
b4ts/+/lEFvNNzXim1U7Dfl11I+Sai08m2l8Nee89o8ZDgmsZ/ey/CvT0sXp
I8fBcrogFbl6gy8LHkT4gFQ/LgDS+qTHTlKW/lQQA/yXkKovUnIJ0HBe6gl4
m7VW6/wQC/NX7sOnZf5ZO5FEeI3H3Buq/3p+bHQLsag1weLDv5PmjJ3v+HR4
JAwoA4nQ5NfY3Vmtj9RFuyJBmrsK0YyTxPf16n9sUipLx8Q3I3PTAYN+QJfx
IA3Vxe4to0wk8iXU1RKV5rmR7nzDbRdK+YXh6kdUisThcmAZGpvLu6INi9Ar
BaiSO4AC/0NWvjGFylfsJpbFnd3JAsCqpRrF8itI3Oryu5ti2A5makzCLKQk
wkbXLakLQhrTUCaVy6+Cvs3BwY87MOX8EOa8S3Gd+KfY1XDy6ASsvzTPzyDw
xtji8rkAuphZugS/PucY2YqqZ60fo7mQtt/gZQhzKcNYd9tfb9Fn6xqP2MLg
danotnU4tGDNHWu1glAvEEZfnNVRdpAmMKFwjvO3cMb+8z2CahRm/FwH7Qzg
CyJtpMeIOdm1FI77M2ER8HNaWUQf/jPQ+A+2IWdk8wIJlCPvCkhlPADgYf7H
WnHH3H4TGZzLAFBAH1cWNokEtHOlxVANA1v4sgGYhNWGPH8ZO72HG6MS4gkr
iVfTz1VmzvHjMT+SKZMf6wNP0zeTtfKavgax4NWQN+3/pz4IX+GfV1UDLmV/
Y9NticZezl0aIKAgMHjONp42TEP24M2ddt4qvEwvcrwESYl+rF4jEIAH/k6S
1zg+kQN19mTdbRqBebT9rst5JwNfKkG5N/3a9SUuZk4UkR9xpSyfnvjONAwj
4A3TlM30R7dGDpxdfg8QHJmItHutaQ7XGejjxzuqQScdRtGSnBVuHZF2H5xT
ugtA/x3hU95GuoRlFO5hD3krGyGf2dBIlHP9EMhc8+pBkkUkpkqxzyXqdGWB
Vw+lBkgaiCKZz11e9Khd

`pragma protect end_protected
