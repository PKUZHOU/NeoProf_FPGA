// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
S7srlgDIqMKQbDI9hiAoRGa2k/rUSWbU703GnDJQyowHmTME3z/ZO+wnUmym9RPu
jftoHaOZN6mEeSuFZBoBd5SwABvyo2xTTBQYhSy7DMWfeycsOmgDvustrTkbRHIX
dLudi+vQhjzJ/QVMiy5cGd+4xO1CRCwCeCN7Vf9z5BA=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 5920 )
`pragma protect data_block
UcyRXx6h5UX56QFWy4oI0KSwh2TDP1vvMKOWRdf1sAbVQ37WWVzuMjkfjb6FUOQo
y3x8miN93EQvIQYuQhRYhcjmbtsitzPiUrHz9d/QiFN0dFkTDIHTPNFXrrHH2xyS
4mRWPmJD+HiAcLtsrrg0U7cdVilbv9nZEUXOaVPnOgeM8cFT0as8A3AkzsTXV26s
qu7MiOOVkO1vTTUJ1LbayOb8rCdpfRljOQsGVvg5nUIUN1dgiD5EfQVuADdejOVH
5qVvZu2+QcgIDCeKBcyBOFJPC2S/5drX4sWtV4bB2QhoS6hAaX4rWpuU0O7CbHuG
iJqWxzkKa7jXlsTdkV71oHxwwi3Egu1+E38ieegOKEw0n89PAG9fPqN7m55bOkI6
oqNqCRqqqGdeomCtWjf4xC6xhu9F+A+mXuKpfJfVn9q36erWxtg4oq2G7LDaS0Zz
Fw1X9EBUP+xx/P7N+wUlPuuLG/i8H1LgHbpMiUtzx9YUFFAU2nVbWXO5lxmqeiwh
/3hS3umytX8ZUQ3TQVNLKRy3Y6EUl7oZiNzHn92iNZiE0bqZCPN4n3UG9TV967y3
8Olbm5Nzj+mOy3FSgCnExLj2X9DswWFut8v42HP41PkmujOPhJunHMgpLYNvHd/4
T/l3Uq/tgVY3psXaFRZ62kZjSCb65EzdwdtIaN9XERLXWBAvT2W6S7D580WgisAE
se5SzHAarMO9TunE60scKMsoxv2Mgq9fttwYGno+LwWyqBVgT+ArpPU2ilCxep5p
zS3NUEk4dnPfVbD7Ig1c+e0XBDv7xua0BvqSuzaqaBsZdkWLLcBtHBzUoikHN0jR
QJxlEc+y59tjRRvwoU5Fzfy/HTHPNAgw7oUsMuSuLxBr9Zh4pRMyPkxoCqhIAPxS
pUT8R8O0fWircFhMDjyC4wSb9E5PUZYYDavhQuFzSgigJvMx5pocEOcY7lqQRCsZ
hS2uE2fNGSwBj6ng11QE120PL1DYAX4ZMVfdLSjfVw2cyw5wajMN6OBcJl3dyD0t
DvxM81cWECQHqWlsd7eKCtxYYd3Aieupw56/sgQTK0t+EmfntYPQzHuwBsWgRLyO
lYHKhP1nSfX4Elc432Lxd3JqI3eK1C5m0BDYZyo0q1RoBjbDUVmkoLNi0dVYVLPv
KcCmeoiozeIaEe16LV4B6x7cGV2jii7sv5SRe1JNwGqc3mhzl+agOVxiWEJTS4W+
PtPhI/3Mpsc79bMuQIn0B6NlhHXGHbv2Xf9+dnKeO8KuCJJ4hjFEkzgfnksZaz9/
gKetTVNv8XbibDZauGh0x1oK2AfyDs4vdVdvx9J1O7by47ggulOxtSIjyxMQUWeG
lEtbDNo23Y+3PyDFlsNPTZyXQtJemMDYZ06RSQeVAFsBM07KLuTicvez+klmmqWw
RqXXx85nux9OwNA+heM2A0FJYpha9SWac5deBBv/aBj7TdFywUD9kcLDwJ207Y1o
QMzygL4tRvNTzHivFP/TS+gOsj353ehutkzKONChtZx9Xo5DyV2UA058d8wfpKdE
ds3KIJA4jGmVJ/Qsn7AJYAqKvUJotdyWBGUUUmPeNitnU83aiwEAIRaen89hAqGE
zZ+LvZ0R16naRYobcsry2JrZ+9WYp/G+EBtjIQ2vNir96e+FQFmcIO0W5tC+SJE0
rQqxYgtO7ZnZeANeQ6VJ0vrrmvWx7VQAAiP4GMLrc76XlO1tu7f6ha7bwH+F8wof
BLAoLRUunRdZJY/KL+SXslsnJhEUI45uIMNNLUHBpUXLKJg8/oo1z8Jm4+zxLtnE
4fvzlsze4EdKqnP1hu8Rh/8suLwHUj9rGIOLqTigDUfP64yrHmkbMCzBwxQSgcMN
ne3iESyIJUIXV3zLl4hIa+tJEsm/2pEQv+3RlON2Lhtee0Qs1SuaCTO4aJuvLlht
FMou2sZ1HGaZGXtgzhDjVOL0l0kW20ISHT8TYBY5kr/0r3OnMYYpiukCGnO5FSy8
LoyOfmdoe2MD8EWEu6ODdBnMl96cc7HWmKma/41gfL1uMIQP9Vw/stSy8rO2q8G7
vjOx1+U3L4w9O3PyLhs9iYbFltuN+ijOG1fOp/3rdiSs/3zpK0qUi6V5Rka1czJD
1iGML34qqDSGVcwvko0uwh9AirDs0g5PgisBscCzg6tvZRnzOFnnWhZMjWSvRLvK
3Dcio+q4gz9g2MVVigtND11NQWe2md5QHQShjjWjXAT5tY4gAwwdMin/ZQDwJ2E5
QVuWLVBNQUOls4lD9g8VM77sG5uWguA3xU4wlpX4Ih9rDGKHJwMqqo866ffaDMkC
ho2vCsOreVTKdNFZ3xiZ0AHQdfuFp7aPUCrEam3XVLT85rDYr+JagYlUhu5rdRqW
EO+pFMVk436QLjCcSen6Y+5HfTH4j136+lnI2X8wHZYCF4novwmOim9W3b2I1R2q
sbz6ul8JSXePej8ErKTyDF5SBBLyvNZWMfajl/Wlm4RAnyWMQ/aKv0RvtCWzZ6xQ
+zHNV3jPrLPB/KUtOJebBWxUfMDQkckt6+iBIfL7QlihKSTXHovYLyO/GtOBYl74
8zq6WwVVm6sCrpLbOQlkZ2CvaDcXfhXhhADppiwuCDbuDO+y2OsiHvG8tj0TZB+P
0tzcw98yxaK7UYa85f1H3o0PBVA3VZ66jmdAS+3Q/weHLwfpXpD45UTTdZDNwuUg
6H5x5QNFc2AH1E7sNQCrScd9QpC/cSbUgnH6VCpHqGFYpADJDGNpA92uIaPDAxQY
n/7JZ7QJfx196w1PA8Ck9bVBjtdPqJJST1lnS6OLY6sWETBqHR79VMhzl8qSf2ER
W4+xpatgldGzOYCrrl+Xw1rvQp8Z0XxB2HEG+IrZqcirrZMmC9xysuiNuyOLxy/l
duMVFKHlwyXeYYchKkLD6A7dCOxsRBI91DnY+MbuIze4urUinpqGtaztaIcrJX4k
LPZhU/3MnMhNlNSewGwiu3VcBuAA/Ry66dVbmLnGg7uGxPrOF5KDiXJ2rn3YPt61
VOQhSz2kXiyvqL+tzyZw4EVZfFCwmY0H2AoLZ49dh5i3lbrlpWEZkkOiOH15hH22
ovmBHr8uxqbw/4OSx5e2tEyLgJ2erAtxfkQYkpQjo//Kt9scszuyWskgNkX88Wya
rwj539RJd+WTDoVgCOQGH5+tA+gn71H9jhZVFvmuXCphYSV0Y8eseg/mHo2lLJDU
ng5fnEwTtYds15wyFlMpPaYD2aCg3bBe4LHtnyju4x8fRn4+l3Z7OMeCAgwFnZK/
afrH6b0wnaP6i3N9pn3SSkVzoiDs8CVF5D+Qc9L5zGl/grtf4m4yW609tarwsgDk
dKRzIQiQhx3j9PtPmvndUd6oKUzzOTRrt+ael+WrzL/WFol7q6zVovvxzHitdGi1
tbQPOpyRD91Z+Q2wuKx7odIfscac0p0VVXZjvqZG6yryBgHQV23sJZGk7+AjcpIX
pQDrJLR+vmSf/20QhZQ0PSACd7egVan19VdWQ4lxXXfcJKSfGP96bw8iIeP45r0o
ArMjG0YyQ+ekYZlBsRsNo6kHBWZJe2yqF8eI/v9tvYNe98HF5vVFF063cvJdThy+
ZuspOByGQqr3qldeMPuitaRMTCny+QGhv0Z1WvqO3wQRWCp41gHK9AdE0kW4yEJY
OpScxorBZSglldiN2pBdsS1MdUC8zR/ASfA+7lUBvGLpYnMNpESq48lO4KZ6apSA
BNB3kItR3Ns+jZAKNizgxk7dcS/3+asomyToASJ90HmKaj7ZcSHwkMr3G0tUBXWG
BRfucaxTIpq/NzXWSpHY86qChqzs+4TgdQGNjbG4h+um7EzRxIdJL847GTSXLzKq
yyulqb4lHRXkbnclZwhLUNHX2XPGqmgm1pC7nPZOnn7JVLEobZrIQ4nieXYunDrI
tevUpG3ZuPguiRLzVQTOyM0SbOHxAkSEf1B2NH+/qdAbKlGx8ekcMjPV7704cRMu
wEOo4U9i1Zk39RvQrL8OgEfKbNre+MBheVwyfRsphF2A03W+XgVy36L6Pm22DmQQ
bb/8+loJyMMVCxEFOaAsrubWvZSJfu+r2XpFd7qtJw9xEkuT2tYuhyLQGu1MXC57
KIC3e+fUWwK5hxC0hLRGyptuX4mEkbQXaZkf6XDYwTvqM4skk2q4xBbjscjo57VR
jB/TK88RmKVb2030NOs0R8pZzpc4FRUkSFY7zlJfzIoZabRTXoMq4b1PkE4B6qHX
GXraL5EhyCBFsj+jn5tgiHx6fsvgp5AdD+SIdajxUlAQOjphV5TZqmymshYYk6IG
WO7zIyJlgIGDFbd6+BKskeaY6vzM5Vlr0RlNtjdYeriSPD9I1TplRER5IJPnQn2/
1N6fyHwnPBb4nQsT+rgLdcVYqE6VpMw8m9TUpfv0ypPpPA3YBZAgvoWYor5FHLYx
BDAnz8ixWk/IWn2pVb6ydWO7pgLKsmvr+39qkQF1wUHNMr1UobCvtcFp0usk4Orv
fSUycGjfRCh6AN73CvDDSMTXfOz7rWotHOa2Bjo10UHEVAlQ5d2lLQfavvlaDip7
FquEKb1Zb6a7zLRhPmDSgKPE3dT+/Vgls2NQWTdMPeH0J/Y0+dswvbVSwMa71sKy
m5mJwSL64LjwQXvcMRFkxq+yD1qJ2qz6zjhOXMKi8A7gLvj1ZHp8z6F9SNVUHZTS
5O1jgft4Y149yR67tohfHIXrcLU6WSQWiIe5N3B+2JHmdTH2n/19SPG1sskSm5TY
dCQEie3tlaNrfBvlkWWQI77k3IZ+zK8QiN+SUjyJhk81Y9UlYEBLTNg+jYHdrG8W
7oxnzIpF/n9dRWY8AVhvuUEXbnJXHnNMoLhRYtMhHG8F2sFPUSHBq2oV6rTKT/hc
POqqmH1080R2jR3oC68K2Kt41GWVqtL69LYVXQV/wfJCf1k6BwZlFX3m5uyiZdk+
H1EPIiDgn4j9os827YS6BdICfB4JXkN/gOoMTNs2OAbgXWkClsF8Hfez5uSWZjHN
Tm+6NBRXKjZv2LoSec9cgxArkqufgebKgnvZmg/VeC19gY6SvoR2ZfJI7HDjnu6v
94zNYySAhlUxPUtXvvUFo7hXo5nvlAYeWxU8NqC21dXlFSe0QhOsZh7WgKMdYq2P
VvRKdId0Dq/Cqf7iIPSi3k8CbOwZaIggQhTaIXN/Ft9wZKkFm/VEnRSzbFFlQj97
9OtjJcKEbeS5BfsVT7jSIdIRnsj8SQxf6E1OWC+XN1iuzGqtn67f5CC7dtW678VF
Axqr3dEJDHku7zndyBl8cXx12JmhbljckpPFELVztHyhC/8UM0/OeI6o2MkJcFNm
CK6V9lqcyTZDkNfsUnNnNHx88/fVErhys61q7sQiTRQp7XvuOZNyOpFwv+gtfCjn
CcXLG/NiAo+WZtcwYqeFUAvdfs+S6KeLUfyQboVxTZyjXg8rZd+Qzc0YmU+15OCp
k1xuC4tipzMPniXYzov2CbQ7OH24HzcjbWg3+MSbbvXx/fRxkGSmP8sL66UlDiue
Mt7tW3R/J098EqyesG/K5K/iGlpPvDMwxiG8l01EyU0c7R+BjCTr5WyaUtc5vS9y
onD7pUnsgY3zlFAhsGLWUTkaUrDz9BePHdjScx/60IUnxkkL/L0kWv5l+sE1InX+
SJ8mZiuvF0mmaJ3Fpr4ieCv8PSnaYR7daSeN0NnytGKyJbGuCQLAp+FE2WoIVbNr
OzYboZikUinG4EhCum4+QxAU7Euuz7QPpM42NGRpjZN5jPyjx4IfHkFIz0pn0UfD
/HZnlIq8qt9MyPHfJmLbgvdvWbfPL4ab+hziCm0zIaRWI/KAbcL75RorCNJlY8o3
u0QeWmIXylx4m/zi+fOCgAyXObfhlvr5B+oWJ+AH+i93xprfrQ5e8rAQ3f0gzg16
8KuhdmlPUd7QI3u/IjIsJWhi4/n9VFCWCVQN5boe5rS7RZkt0nqtbI8+67j84Pzi
9ry1tGqEhKLl46MvCR50L5Inq9f/hkXvIfZ6q40arYaJIMkn4/r66JrWQn1b68hy
tqNbvFi1whq4tMy4bvnt7MBG+fHeBaFUGCGyD9bdXiJU6yscOwPnxL61cp6DpU76
S6fjVeai2OkG49ORLkUNAbkSaSaNpB0CckEWnQfwQ8a0Zx+EAuq042iqvqvbqmSW
hdqjUXbumulHfVsQSzKSA2GI9bZc3zkoMlzBhE/sJwrSvAaE2G40KDMulDrCK7K9
2pxz9PqEZggAM9hYIcpU9UGeRzMf4kT4X9a54n/Tud/PLh1XthCTcSQK9ZNiDp88
mrdy+ii3ImKLHhNPf/PqIxTsL8CgFE4zZCJjPBfE0JJtfC08hQsA8ReKZ8uOH0Lt
UOWmBoucgToaHRZjk3bbm92v8zeYUP4nzlxqZtP8P5a4wcV6SNjaZ1A04TRgcgER
A822WxA3tClVDLfB4KaNjAG0QUBXH3yH4WWw7ZZj40muUjNFwwUh6i6FFyi34WSK
GwuM0i+/s8PpyLQPogcfzeUchezXy8dY8z3SQnWcvG+1IEvZvR0PN87Kz+EUZNsl
rRGRApCPgmEMBl/yGXVr70z4KoNn4NcXt8eipy+SecDbNKzsuaNIzYTice2oJX0K
G9uQwh1ggtfWNSjA/hMMHUmh4a6w4UVDDk2alhc8e5vS6iLAzT6ptaq6yqWVosBK
P2lwV9o2qrkc2xNdHgAmzZ+5bBFFL7vEAgf5zlwXK24seyc2iBkvUGqarW93HseA
WPRXQQDswNFL5hbCzuHQvs24XcMOUx/bn3cBy1tLCczdOU+Dej+EeitL4GrzMHTl
nIjcY8CT1oR6Xn9ApsRoZ3IQt2w2G6pA6KRDXlHZ4U8Vzpb3d7+kQz12agrNvjOm
w7YCFJBbxk5mqOB2s4ndiO3M+Y4gNUitpEg18Mlyy1XMs7k+kgwsDOotUYQ2SjOg
Oz7mCCC/bPfj1V9PqbkK4uBWVKW/4+AmYmYUTbujT7ma0cJkIXVJX+b2+pwUUJUG
vH6nqYzEuPd4HOd3DPcpeWFXIuUUk4i24WSDW0zf3V9CHyGy2CbFwMsoGh0K3DKV
U3ODuAPcyNzkxBiqn9K3Kw3Ymcc3iNPIoq729anf8igsma/UEsTmwU9ISux6Ns8+
pyrKLFkdNghZRlB/84m5dpif44e0YPvyhKzTFs7GXpYRZygvLx5jXTRCTV4FFO9q
Pnh+rPpIjT3Job3q9zltl8+n81fcCslrdayNtbhawy2XaNKyAmgZsvGFsxPAo2Bc
Ts0m3sQkvnFD6ugv4hU6gm4xbPsE68p/jX5iuCno8/m9CsFR6IgjzMYbUIcaPnk0
sciWfQBUxUuz+NFDmi7WeuhZfSuekLD4Z6P2iTx/l3xxc8nVRFytR/PWkquI2DhI
SWO/5I8vlh3YYmaFtVsKarxeTjLC9VXpljhSKw1F6uuHuW3XS1J17uioKwDEarBg
CZ/+sNUyGKOEWxY5nYmYoJ52rbv2phNAVSP8tU+dWp55S42ynuJOJR/vYP2tnUsh
Guq51nIOlY99Edp1uNAssdky6gxHSH8EKF/0N7idWeLqnJzNCgWXEByIaJBavXn1
d9wPH+ZnKE1YFy92e/awtA0lJQ5VV+vjkRjphHWlYiW9jqH/ztxjWRuE37qMKJc1
yHA+zcB9z+Q/TBGfftKQP/FFraoZq0xyztKmvg1lDHxy3lKRUpCBwdOhnyOxLoKf
JCyRvfPwxVLKhISFsOYpTu0taeO/uyk0aAgznzT1QTdXqJwiqR+zWtAgo9ouyF8a
ZzRXcgjKKwuTgAEyIqKe5vSxrNBhstyQJuCc/6U8sovKXFT0Lb36+EUo47L8fQVs
utg6KO4rjtwUVxArgE6eTEKQQYHjeZcGWDkTNQO4cc7fgATeoon48sNUKNcDIw2x
1Wvk2tB5AsrsyjfKNwCRqQ==

`pragma protect end_protected
