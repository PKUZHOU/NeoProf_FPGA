// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
Pac38e3vv/W2vbu0nrhRLS9NQMGyPDIVx6HDuzULtix1Z3tPTTIlWD0Cfe6L2G8v
fwkQXD4nV0/8saP2CNuhbD+Rcqa81h8oea2sfwmixsWsdEKyjubu8QDQfyW232QM
Roi3NJoFSOeem9AKiTMltHdTtqoc6bnI/HrVa3aHdzIL/Q+oFx+3Vg==
//pragma protect end_key_block
//pragma protect digest_block
FarQjuI7X8OOGYPigHtQAmb+zP0=
//pragma protect end_digest_block
//pragma protect data_block
NPssUp04sUoyPtmHGB6ldGWv4ddG+t6jHntc8LHDFAmX3ZGzLPXL8q0gY4ERjCzr
GVnQD9lFqUxenU3sgJa39oxC/cxcr6os27es89iH57rr4iThgHjWj/LlUR4ZC7+m
BoB0J9zhYOWeRLGokyhwaXTdZ9Gfg3z5JHTpOr1qaUsJUMfwxhB/HXJymsj5xuxU
HV16v39dkuYxfoy7uYxlsbc/4eKKCLzzxGJzoIsFMSHvgjrAro8cQkvqZxWVtkl9
6cWISUZh/gq+ecfWyOr8yKhgbjC6C+nnPzHhXXL1oOCRRxOs+zsln0cQR3F0RD4R
eND2TAI3Exr+ubyjV9mrrLh2N92FprOLlwUb39X8tCvsqzzoIdh79jjrvQ54DYrA
ZibUjZQxPlpu+OsKCIh1BW1ofDFtsgOou5HfgcUXvNClJ+IvA6h1zwNi4M48QZYD
lSAnR/aPmYzA0QG6/PEvSKAoUQjG6A0fmageoQy8fF011f+WTB4QKaEagujVmAvA
FZm5OZjl0agYwVxJt1wKLR9xQ9uDmlBTmV5IEjkzzA53m2fH4VlbCMwXWS2KWBZR
KKQnrB9aIwgXUNMiXov2Mu9VhCNbNBQfVr2TovDHcBhkOzr7LPMMQS1gNLUMfxk8
uuWRaPVNKhkfaKLYA1GHKU2sg2LBBIkpX9eDW7SHx1zfU+Y6XRLBqxQ6pfstNqND
wgHAKwUlUbrYLSZ6VOqYjGG35UcxfI6Uy1nKF8D+tZ85ED9DIPZHL8UQfUKuvRNO
4bPEoPjqsCPnFlpMHbx61WJjHgzMokyzsmrJ904m8ubMGRusXLkoUwVt/g2f/KET
w8AYm3D1VqMKMhbPJobutgV5yTAvQVVf0ReolGVhkyYlayxFVwaT/L6qXae+KLXa
eEw3UfbWItx+next6kb0GxqdCpJoiM5w2Q22NHE7+AL5I4Hizcn7/hwHpwyeBkcD
cUzckx/KGdVcjKT/5xJuuGYfXteRSuUX16Mq0PNitjZED9UWlgbfPFb48J0Cj6BR
TnXGBUCDYW1OZ4fqu+Nmm9puzMrh05jsAeNyeJZ+TgBVCnaSxQLFLP8O6t6TE3RY
ex9aVKiOSRKqSjTfpP7y2MVYsLdaN74g4PWnsIVI7iH0G36qaDP6l263qRsxIHMK
3EftJyeWK55O78+9xOsddztQUdH96gbIF3Fi9OSYj9u0s1zLoR3s4EBX1bBBsV/Z
t+22QDj8kCeWGcG8HrRWJBhCoqo8gZy7Zn27LHaS6kUBa68xO62DBUKBFdUIevkl
Q+wgtIx7wUEbuQK5Qhd4WuNQrKOc5kff3GPfbP8IsEasRggQwBjnFGfRtDZQze+O
4Qovz+ylNVMlsU5s/kyzcAZTOfPCS+5jxHXGSsgGMYRUkrhIha9fytfVicJ2pIeO
nFRymwVGo96Xxc999bqwbzs9YPnikEp2ukpfBJM7XFBH2Bum3Xb/QEDQefjBiHsc
+kzHe+W3wKDl2Vy/AzQiyioiSnMDoeaQDJqbx2+PX7X9HgCI8SQXEoXawbBL1Pq0
9BqkYq1DKrnWcAFeYBUQJk9KT+DjJuX+zqi5coFaYUnZVUIfZ5A1S/kg9C/xCBLE
3UdTI/h00gQ8oOdKieotKR4Tyg6uvZpUQE8uGp8fqxJFcEyEU5l4t/v5DVUdmhmI
fc/YDk21WGnsJ9fK3QlaVwraiHcMkkW33JddXD0wnZZ3u/+83Iowjg1Lx/qXBscx
NRkaIjrn4mmcX+Kn1HLaF02n01Nf8ZdYlZxGxAknc/adf8v8UspRHsT628WCM3GO
dCIYt7P/6WjGDciUm2p6ImFrP3itfa+qhizU3WMFLsXmsDHoQ00HgYBfBO32GDiW
HJrKA92iaxOLIA98T/gw4ZEekKyd+kzz2z9FmIcyMyaM2VjoG08Be7alAv9Q+kp6
LXK7sVPROeCUYDHeH8K5qQhKh4ejdLrpMxl7nxRL9HdeD6kxzIwdmC0aS2AZVDXW
eDQZbUPuSI8UHi0b64sGhcWGLoprYN7Hk5huU3jHD4EmVGlmdTMSkH1i0jS+5jxb
k2w4/HfZEXovOGP0eZpDRhz3aWVTPtTgz+lHHwybXQ7x16IOIo6bjcHiq6DOcWxl
Z46C7QTs8toCFcSp64VjLWrHnxwM7xh8a4IYpdTX+7Eh2nDW481NW30ScNP2sbJu
nV1Xo4l21+8RzUX+Q2u6qkhLW88OPVssdYf27EbSPXD50wE665PqI92yaw8eXMcr
H8q7v2nXL2TBswXj9Nv6T+8xNriTPCrbf3iyPR6FCMxiFZ1wWDskHEMVagw8Rnco
IadXzGUlvc+HlB4Qd6Dg+wdNm04oKy586ZR6YjAtLqIllH6RRn36PTBLMQoQZLzF
9LUpnUq9X2CPFoAV4DE2fxWDULB/M5gDZEkNu3JrQPEFC1sUYV0g9YfPtOgceLkd
YFVrFHv663tC7IHiIhquqRUZEirvRu29w64EVYmJxkX5oV7SqZoCxJdb6Zq9zHUq
GRLWod2NNH9NFBMAPO59/Yga2Mmr3KwFvD8MCh5n6YFn6ecsI7OpALTgfUl19RYN
xBVheH1MNVqgLTSSSRyqJ0LlLmR+efZYNO39oinVAmOjKHQ9+vcwQ7J7Q7c0toOg
5VDxogEq3ueeih2ZWJTj7ntnozHJNPLOOEhiUbXZP+p7feTU2Xoct/YvKHI6ocqM
Pp6om9mrBjrTaYONa9cOWT/Tc4IipcDhcws9pZKKr0VFZRSbQUwgoRymjac/B6GF
+gFBP6Ronu5xRSMQF8tK7M78Qv7J4KSNSoFiPxfn3FNgjzsl5MRLXK/dP2AZvNLw
AtQFIXTQPulRQSzh4X1Ruyxtl4BAH4wQwG0ocko6IZrZjY+tWpa4w1rOeJSCZkPC
KBM05L5fOwWZDkD0UKKwv3BwQQ49x9OOqYEBRZPO54y4JBfSu0ji3/pfICuEsd0K
hvi+sQTk+ZWun76b8IU+boc2c3xW0kWY5CkTy7qlVANIwsK66F34ra10kN4GJkFN
ncUb+foQeiyyQso1AjJeEkpEzCCqFj6xubjF6QLVVVbaicNpFZtasq/Lx598MHNd
0hbwfxb9p5Eb3cxWdjN22fblrSY6nYosUhKZohn6BWqqtDZxqciPgvKlSLSHDAkC
R36gacCG2Gz3I/sPG8nktjlL+g2Rob9wQhuY72Ly9/6HOJTDfOaifvg4b25RPZaw
Ll93NELinEz9bgTj10kPlYkwLEJc3j5Wmd6yRWKe9sx1JXLpuB8n4fx6ClaX9g+O
T45cuWKCz3EANVahzgk2VrR0GhajJlMKk2MMKcHL86fV/uMh+lTvZ1LL+1avJZJw
7vIZdGTgozU8sZYKvb+6C2yoWB0zieyVF1y7inYXeEcutevZgubpZoaErgEQwtvB
Frb6anNQ7kkO/zkuG/vU09FWWJwFq/TvZa2RACmgsSY3OBAhXnODBiruv+hiyzTs
KRP0XT/kVLGU1D+HChavjH516cEjozJkkE3hHoWpeANUr2EhJ8A/XEmsoJPOeq18
2/L7CPhFeW104GPmZoBHOwpnRHXwHu2ZWpbF6qkK8BII7bIHJabmBGjnqPdYyW4h
MqV17DTFw4JASkAeL2VwfhB0GosiVhMMMeAm5qbMdiTCEBxjjJ0WEISY1xQaIAVU
gHZByf4PcXtjUlXgkR65ny1/EE9yLL8wPRwuLyf+82ktWjR2UnxbRIhQuRCPTE9p
smWyv85rG89xGVE7l4JdnbuHTRlfYvTqYIPoLiyVGluwnZtDp6XQ+fWR50lKCpcM
vmT2kn+0JJGQNE5qXeDVtTC5PGkRMK4SwI1J97m6f88busTGtN+NQbss92uk7Yvp
F3aGjG46PEMrKVQQtD+/OHeV/3fPAjyEvFb+8koUlut308ftv407kex4tOLsCV/z
7HLcjS69wZFIOVOHAdgkU2pQAOy7tLGxzMMmPvfUIUblxSde5ffd9BpXEqwb7SGX
SLW+9XYk3IjiyMBAZ4pRholRxXwR549eltSFje9kJQUGBT2bIiwS0gBXRw2LEQOD
DVdIVbS7uK09o3EUUn4eGlb18UrwsH+IWY3Q56AI/Fz5zpmTxJHv4YrO0lZpb8t/
3AlORBFoZaOOkxKeg9Ezg0csSbJahgd/4CvAyghM54MnE9Z94NXxwXqyt3eWNdfi
KUedL69pEsG8H2BmeTHrcoCaURRFcvZjufNhLx/ZOO6bCeuBLHCyYE7gBn64HADq
B5W9Sp5w8uJDBZ6ahV6hswDWMmPYp7L8Dg7YuIDbnN6FmDvmVnGycJ70sJNz9GD6
EsmfqLHv53VJnF0evaL737UtONerGSYzmqI1bl4nSn9S6FAuaihu7ttne0IK4DCN
8RynMAa1D7vOMjHGuc4FUhF9X4ZJDu/IouXCaa6CzenFYnSQZ8Kvw4oIHCXImvJO
7ZXG80q+HvnLY0jKuItm4UyjHTDjJ6Hnx+xcw6sWjbNhtbL+H4TR+G5KbSfccTha
B549vxSUsKKha045hleaNuxO1xLciFunjUKW9cp1waolZOcLuoxrtgOceyBRWrRb
GWspa0h6I5KdKlzME6BCXyHn1907C6WDIJ8blT6naRWgncV7Y6sD8QSKRm6Eu5+I
fdl93zrZ27UOTe+1W2Zjj0Cb+gE9XyJKD1pap5pYwUYLrsQItfrvU/U38JjDyV48
NrvwFvDsLDq8zcN7Rci8Ylx4ceqfCtcsZk2XcUok4BfoVftV9bLheeJZbDugskf5
nRTzu8mHXKGEkTk4nw+m/ewCUJR9D/BFbbqxU1bQbo0y0Ko0vsW1F+WsbakzrZ69
UilJAd5oYqJudayViW3VRNFiJv1xOyfVvfxr+dxUyX7G29n9+sH7dWkRSABjGF4A
XoL5lM8OxlirGah5QphniY6rXtaYhjc7BBxfk7VCjjX333YUq/FRAirTNIuThGtT
LsIwvdTCwmMrNeRrFff5qNFO7KDdz2eq5P+lL0Q+OwpPmhnM4J/Ab2X5k0UjXutQ
wIieaZvzOefxmyeXH+XGz4AMckWokErtYY44/TmxwqvVHAsBFTZjcDG+V0XXTyNH
M4N5X2oqep+k2oidoIHirTDZxRrtMtrlCPRseANeSnelK5o6B1uNogzoXswfM6Js
mrSIbdYCmL+g9ktDSB1CtcA0M1AwW30+tkFQZCiXSeK6cWx6vz+R/Wj7j7QWpqYN
dg0gLTuAgCpvzQ54ZbpSC0mamrEmtTLVDYBq09ArSfV19fI/Sw0CMRD/c5Chztxd
g2bZIwWvWQDBihgIz42H8WSU7btDo0hfOsf1Dt+xKAFb8fYQq4NKXl6LT3boxRnn
SOMERkD96/TlO6jt6jTcMCqH5m7p0LUrSSyBONRCHyweoqIkBlU5DmiOnB0kzPJv
y47A9J2p40mbBX/ISg3Cjhw6DPjLlFuJQJ2g9XKERTJ+DyAFKmRFOu1RwXW6Nq+e
MgaTA/r7xoiDpOJ0ox8dLaRTn8q5WUH+vRAQwLk96CKAv77K8TkBcIvd42SYTx6a
Sk8bVLyF4WO0h8DvYAh53pMvixchUQAWaVIKsetMvr3naxr7zuzP8ycecPkBMndf
TdvyAwfbHLv335ad28cvqWhOUuceBjD3SJq0JAaBDnJlvnpa0bDVE0bZkSABgXen
Py/OctflnDFQgaW6JnTh7WISOOV4m7JGzp4YYRwn5HRjg9gkQ/pp1+iwmoQPZBVE
/Vmh9dH6p/KPHv8QTJrMcptgYnRzhzjk8YuFaVDg3pzTEhQMpCaUV+vziA22zTrz
4KnJQ+jmx9q5KuV6jn/qBhVuNy4QaOpXP8Rp+ymogEy/ZgPGoiZYUClIeciqyKr/
r8f/A4Ns5MmUDdTMb6iHsqwhGXTMEZ3nOh3fyUnNJQ596mkXlDHlrJM9fpyks2EB
fWGGQupVrO4iUkrA7Cru72h3dTjMrM4fIrGRNfpzhBNRjvSXVtpqhQfxV+7uRpet
vOD/FFKaReJnQmwT1C213DFQiA7bqlURXhjQFLB/fHnCQHpSaLnC2gVWJWYWGzRx
1zGntldulRkd/WTZFc9n5y/ukeiURse6rfak9PHD/KDHb1FMF7D0XxwnHEzsBBos
ghyes1Ic40v8EiyUIphvhkZN7DNxN6XbI8DiTc2hwwBEy0UJaw5xi6mhEGuI/GpS
hweqPSGRso8o7x1lldJAwLPcbCJQzk5OxrZ8/+F/3xP5/8zXm1NXCr8KKK/0MjgQ
VQiU4BGqzLaW0bdxru18SmairWRoc1f1s2JyB9G1svq0esqSh8/hDt1i+ZdVAfBc
ZTMeISy1VNahLXi+Kcs/EUGYFxk+iP4P3vPpMqC08qfnFwCaXuCBEmNjw+KrRr3n
8ycS0feMoz7ysftJ7tswaI9pb5bXtBHhifW7p9VNX8GSrhaKAeO6h5r89Nnla6Xv
g0uI60oil2DZu+o8msOYNRCsasNPnTcYeGIoDgl0fxAkTRHCT364P2q4fC2bagE7
2B7AvHbsAKEzbdeMNuDn0+yfpM8aq5w84SxfcOgqCm8UF0Xhm9JQ9STmStRhd01k
VpaX+4rmKmlJxJn3ZoArOjIOSl64hvzdeplens7g097fAVBLPQLVraUZtcVlo6Z5
ZF1AnFEm9a/bWyFyQiJYrwS5oA34Rb0O6eHXx4lHVhm/W1+zOkg2/DoiyNSvlYjS
+6qXY2ijaG8NNZqfhTp5Ij3KtVaMcYPqaGwj5/b5BHMZvpedvYnIjnnu1gpgUJnq
PIGKpP9vIHdTYU4iIjA9sx3uRbd4gssss9+zdYTy9C7gDbVe5YNxQIgtMh9a0Lt3
H02nnHX2KsytKzvJdrp8kVH0rtZbWiodFbQXqsZjgmSlwjkiEico0xXHvdjFpJED
0r60H6GjiNr+WAadGfYtNjm+9HshL+KSe7/NpUtcctEvyPiofu0oDF+aBioRWEAm
Nh034Ag2hczsN+fc+hbd+oJ+IMJQ+9n3qz8nfRgYT3IMiB4+Zf3EgDtPhBi87sF/
k22YX+Mmh4dkmHs+SxHSShtR+AiEBU3kOB9hLeZU8/TcAHZ25XiOvgQDaUqJ9DM0
dzOmyobaNIoA3dwM+3Db2rl3gCO3N80tUjEP6Z4zMLgCiSbsZ3F5Pypf4GRqmMqJ
w7Sse+pWxIZtnP1iC50uQs5ADvXsrg3ViWObOEB7ppRXlravvuO8zr6j4Y1e3ksT
v0pKYCxbBjZJoGyxD9aJNtm1fyHb3qiv1ezh58ooVTTcaKClCaG6enL9fQr2Dznk
T8N/JY0tXZZgyA6acZZyxHIm7gd6uo1z7SXBPo8yyyxzAj7Q/PgPBKkW0vLF+g3W
5sA5dm0LMNBJ62paeAbv+3eM9FJBUUp6iURt+7bugmmFAc/bLDmSHONSE3TyCimY
+X8sPCKMZnC/ALchZnbhXH301jQe52j0HkancnfnCZo5oUifihff1c2jzV+fMbzB
r8ED5dO8CHD0ZQHVIBYFRFwF2RmJ+SRJ/z06TbeuomZklIU/qXMJ2DVXFNHsRHyU
qanR1sZ1iGj3Kux0NEcF3JPVVJ2Dm5UOUbCk5k706sDXfZ7aiLAcRiLIwYGTe36w
Drx2WfbIMvb11crY1p5P/c0wZ5miOOY6ASaLJxx+iuRHS1DaIa02ixLY51DT+dxc
GPGbgePEkO831t5ucg5WHjGyG3NcpgZ8HddNrN+xiXkCG8J8nq6M6ED2PyQo7+B5
1u6mxwom70V2f98kwP2tZAtHj3VHWHioMK4lS/32CklmbQ1aRXhLEUCMb5/Igl1I
GHHwW+ynnqcSAnqfYa9Enz0Hii+Cs55tKtpbYecZr5Dw510UUcpAfMfgfZM7MPEM
Jmfx//l7h7Nd/qkKzSc2UW1vJT72oajpebFB5hH4jjf45oNQJpA754wFi2jUL70k
/dJG1oIdEk6f1qA/CrjBw1xt1Q5KU0++ltekaQz7007CuzER6gmeRnkFX3MEQzGV
sa3dhQzg8G/6dBofYt9APG1O32vJsd+ErLPtmTV4aPGdoZL/d4Ue6kzE9Q7zCtoe
FBdMcQ/DugyPmUSGeYG7wz1JDsx1eCa7oI4W8JRuwMuN4EIfT4zpMNNdB3qEMZi6
zyJ4OVX4/YWsC6ZLKhD3ewTosVQeU/i0xakDJnusz/St7H6ra4Iieh+yT0QumImG
e7y+VxLQIXkMfwud3+nLMmabjMPeL7nfbNxwNrO4DvhbI+j+U5pTVye/4c1jptQX
hDUJqLxCR+/5UfrIIywZHNunyXkcV15IQ9LaFQTfVqAN1BbL1vKnLvv1dQjpCLgR
zzh2pmpsOr6MQ8oEAf73MushWIYXaxYMvDXZGgICulUfjEQH47HCRI0ZgdgHI2sb
i8Zl7d0qSBdXa/7lrXPhkiOhAH3w1soPqiTmMLaPVWWjvzx4QOwB3JW7ytCAsLQo
0+RZDVrHPNcWCCtK4KvPfhXPVyOwisWjtdSbt3mvcaNC0W5Maoz+LhMEqWVW6H64
O5odRQeGkrGCWTsoPSd4Bs67+QYrp6qX0l9TIIHORPocZiHSuQTTFC06a7wAghL1
mlg8nvGHd+7bjIRMxRtEMTQK/x+bdnHh/ZAqrUxUoZuHnqcDAhXbntuFKJNF5Ng6
GR+79VUBZGXy0rLdhBeKr+rVcShUK+FGZDcjOoVZmZcATf5ZyBeeh0ShEHUg8Wrb
isMiAfhoZ6Qgx1DSfL8Ivk9LR5U3m1lxC2jBAYzWxXPZ/bYb1ZwuDiLId48dTiXo
CcodhhWJtkdbRVTrtBEipdi9kV2Cey624NFUaOY15Ezh3R80kZe+BxOu2aSveE36
3aiHWvl0KPGuAxzboF5U6+oOE+ZtBa2vrZk9+dKTl2GN5xg4pmXrF+HfOZFh53SM
aTCA7xU5DK7Nij0txutZGUENn6ZniHauB/pwrc+1sjLEwfv6VeCRp/2tqbp/miux
XD3q0+9mnMEWlnvaXPjJzx0FM32GbfWynY0lJ0gYCDrgyoPmd5NhYz4wyHrMFixV
10pwfJdE9XsdptCZxwu7pjYB35FISVYE0xOY7ii+owXsoeR7O6NZ0cBWgEwTmNh8
fDvnD7lcCf/j5B16aWiCLkUtfHPNZp0a9X2nmKOzYmgNDcKZ7xmqarhPX56W+7Nl
1FZWqJhj2owZfNvay7/g2FxmfFtZwkMcyhUAyG2PO6Gyo5AmGfXp+9G6OMdcLtSG
HxHbhohNIbUNZQNCysn2oh4HXu4elY+QFcNKv95noT19nAZXdlSTO+rM7p7mFdOC
+0639LL7rEG19PWl9p1bmDUjJOWUUnPYsqzQ52z7qbBlmwdHBGxxWjRDcJpcmGpt
M/b2NF7Cbt5GD+KFGaLnDy8psX8dXk+bVdZ7cDoBb8x3/C2lE7I/txcqqDAoGUTT
j7Uwj5nuyuKLS3fOjogHFsniwU1m0XPklA/Yceqh+mwn0HbvdjMjh/elLFRvB0zz
oS/70W8aW92cdxm9xU9tHT5xG/gkMHYn+0SF1wcgjA05z22wplT0IPTE5oZZDoMP
8Z+ELgMT2rNLGqGnw8uKIqoeJ0XkhEcujtaeJDwgL+B2/CJEkF9/JwNkk9lJoGRx
S6XepCzcjA4oojxAepOKhPlFSRER1hIBxmselMXqyytO7nAbGcQf6o6HZMVD6FoB
2Ro9monNoadtGcHaWNHPNmjwjPOoq3Cc50mqOuT81J2jmaQyELKP+mPyiHHsejZ/
ysPg1f1gIZSd3FsKLep3nZwZmtBersIkLX65hxbXyfPLohSGg4DMj69uZ7gE4lSm
/karIfsfNvH9uADlhQ/J/KBJya1n8HoexfVgKhowrvtDQzljg1DxFzrjbEXShFAD
EbjxlTKDE3uDPUFfYrM0A/zrgvqtAsCTXPkf2NHGKhC9P9zymhOeRLdHKBSH4QSw
F0bRmEgexbi+Smj2NmqwdghQoiGqR9TRSYu/DNLv2BibmTcA1cYtxD9+xDWPSNFS
6FuzISajRAcg3N93sgzNuBMDGXRGTkGwfZFcGKL6CCBYGSTmaYn2+XoJyO2Vvqtg
x9Y/AAw/lLsdPWmOYd6wPutw/m0LLiN4qCPl+7dx8nybwORkX/vUogUdPowjm6bY
aSglFxi2jhGAEf1XyjeQq90xiFIz6MdC96IoTu1hPPYTJncZZ8HvDHZFVjG/CvAf
FIXU3cmsin5EHnG7RWv9IUrFyYys+/v8EVYGa6fyn6Nlsd6eA7p0+o0rJQ/rrK4m
fUmRbMocvlU7TwTKHI3hWeeSr6RR02JOE7++zeAL9EQXj5/EtKfYY3qurXU0A88m
8yQAGg9qiKsI0EMhuCqsk2PGe+OeWausa8VyWyzRksflSTrDJrKSXrg77eOewWxh
lqWZTw0FIHzajmaDpXKqDgVlYA/NxuafRFsy697G4OxzQrJNLkQQrMipSxYhPspq
GfKCO4zVYZ5+659LIVI3McZAUff1sFUPyFbfQYjCtXFesKBGQHBLibh8uRU2FoTq
jhq8F4xIyqm+5PmGbEp/qwzP0PCzuvD5Ef8w4mOje9A1uvgaO+MPuX7qOioDbSAX
HORNblgdP13ECPoKSdLlRWljfFJil9scr+zfhh62c/zNVH839iEVBfQEb1tC7pQA
w9zQX4D34ATbhrIoDZaWJhnz2Id1x0VZH2PsePyTr6iOiNlQCYg5ul4V9gbfdLAA
xy/c5kAfYA62U/dUGO0Ra8a8/l69lOe6dp8nZTiAUI7rB4gnvqHjElLZ4lHunyCm
rIzPJFX4QsXeHx2S7tXAirNChMQ3YScxuPF6ugOr2pcfCd0hfUnCQ+KiMPsb6k8a
FQM9j/E9w5ook+DFyUbrjkhkFfDtTps3PEm5koftiFwSf0+3Al/KiFusimliPssE
lFnTeZgTWEK+fv/5xq8qW5pD2ec9fJi275PfwAqhDC5hE0JxWnrERS86k7joobmz
C7rBA5cafLqnJnoAQFjFirJbGEbHoncF+X/VHjMIZ++VvnJyKLOuWMOhrd8l0vtn
F60+b1ssTdmNwhCCNL3/SLP2hUGZ7qZ+5mzIAzHAbT8CWJtKG1YkXmDpxyDVdcz7
cc47e42aKXEpvOo0VyRXqr7+0A/LuZKWNraFSqPUYsOTPQ3InjJeTS3Mi+55bdJe
yMpz9Oy3k96l+T1GRpLAIRr3tNiHWFakXmV2sFAJzAeGgfVXT8ZL6TR87KEC07rI
MIWGxTm1jBA8quLiA+etpUquSVlDgugJhZKFRNrskTqAdXsYCvv6dnbDllAPmtzY
GQXPitg2oQFR59nlhh9KV+0Ddjft7lOn3/IaPRJ7HYxvxCuKB1zJSnFSsnARjje5
45m4Fcg9iqP8dfDVjK/kkm46Et/h2ePPfSJLC737r2BOmVnXdXoA/gUFQTzjLxDb
SlwhxN8lRA0nn6/YmE7kgEQ3dgVuNPRjfeCOlEBsG3nF3MRcZJo27pj3OneX4zcJ
SWJDUxtTHvxHTtBECO0cOtZFw+aKYv25/UU4hZBFaVsj0Uq8Db0rwl1atgH1N7kx
+4bpkxSIuTQlmY0+tYgNI7Ju4NmlqEUEN+S32gCF+xcBmw2vhKgfEuE0Ol7BaAPb
7pg34UE/WO8XNXxhBA7wtZEYHWCND6N5mEMiaEDW1v6d62B4Kcutqtg5aLhpEuUv
33+aap8fLRVgawffO79Nbj6JlXlD1M3KmmFk24trx9mLKBVEaHilJCFZr5QpUbd4
7F3GqMq0xzg576h67KSovZqu60yjhUMpGX777IV11sYAdVPYBb/psyTi8/VmgHsh
LHoU6IHikcpusMJdD2ORbmkiC5dIeFSS3dl3ni5mmtaNv3Nkc08+tS17O4f/ThBx
u0lUoxyKOzvxMC1ufii3c1dSXjwfHVOdoxoAPLN7XDAjbW26dwWvJ0XJM+O2gCjJ
z4XrGWJfPdRcr4NnuiXnbVF805+xOWQBFl1nHOa/gZJA2kzs9i/s5pQqOCAzRFh9
gIaGoqkr8D5cYWY9o6qihseI5rt+r97k2qIH2t3Rp80nS6bk5cshlLm30pyvqve3
b6mHHwYJb9+DGEl8NdieAmL6bXBhoFdHNf07/LjYYYn54bMxBsH3Ytdh34f2GQUV
NtVLNWyh8fmjm0a4xc7U3Ohaccsrbap0s2A/KaaddbcuiDGj6wnn+hQiyPI/Dqi9
EsbOShJVT1IBDy468EBc1IxJS3chcBK0DB6J3GIe51UrfXqhNwFi+VYxoLYElLQR
/GTzgVp1hEKzXgBG1q9GtauW24qvF/b9mjUD9DM05Xd/KImgV4a6TE3x60P00Kek
+o5spmlbGppnt5h/yGq57U4G9Of+qJp8/XbhvChGrIpqOU43LNhO+mhbvWB+NFnH
7kty25g5gdJMZRfg82UwRk78lLSm6wa376g2T3n8i1nMalbpnP4AmmyDGJ4luo2V
qABix/uz3lk0Y34uyJMPL26MSjY5lYiLqtlmjRUbWFlFImS7Qvk9aeq+jQWOHimM
TAc22Wk18ecBtmH/3HJPwXSW3rLAPfS+vt7s4aSlQFr++sR2OuNtpzuK8M+ejdh9
SZvgG0UrI2OW/dtr3j4Z17GvF4Q2EpSiOEDiHR6vURiZlOcTh1mO+4LUo1JBCKwY
zVDdgOZZoLQGOocxJcWjGcnrwk0BPN/Z8hpGmKWw7ePmmOIlUEZPbaQxFC6kPQKp
o1w4zz6TIz1FBGcE2MLe4gzguIfoF6RnsZ7+YVr07c5WlWUpiDD0Y3aQdlMAxNa3
s3fMU9uf95OSnTgzK+jrBNBgX6YwOp7tcLx6gOy4YWfI5FdkjPu9PqO2S6zAJ9nC
qCxwIzd00F5JsR2Z/NMlvGuqyNygPSocA34KuldVSippcX686LleIQgmyd9UZ7jQ
eE+WfFz3DB7yvO1nrVGYcAjoqzDTgqmKo5iU7nHJhdeYpXsVMEMWzEp6/5r5JjD3
QbkGKj/w5Xx0egwBPWPFAs+ErcTgZYmsLK56Iw8OmY8PDSNyPxpsgR9DgDzQr39e
LAc8qD4mDyLyUIvu66DHbtjl1unpnfJEJp0hzRrOMwwXpBAB+7B82krxeEjNN5ZE
n+FKVkds21xU+Cttd+mEr1BCJmS9sOXez5ofqzkcfEft6iTRzsv2LHBNuNjv9zj+
B6hQY/FQP8znIrZaT/fLDfShXdTSlKLWog8t+cnZGlGQHDMx6fvDieL96CpM/13s
+ecrTBUc1KSEjJnHI842pDGp3Z2XsWNfFT71XjCau7pJupgS3ECNViPEgS55DUKR
Xpk6fdcA6p25EsgzRI2kgKm15xZfwv1c2m/JcIE/4x2S/IG5uXhkwC461c9sG/Fk
/yHZIg0M2T7MmfT5+QWOywLDBrQz8P2I43uQ0C5ODVCvUqwgyAG4Jm8vFOE8lBGR
N/eZATe17KT3gRmuKZnP0OpBeOMHZIkcZ1uAo1mecfffD4FsYKLDHt4KHa2KQ7bu
VK5MSc6aZ+8qv4+vtqDKhWvYBnEsaWQ2Jbo8tYzH5VMl96ujoIeIzl/l1O1NLRu5
cUW5Ycg4uypnedDgYTnu88G7hHH98A7nJrylNn35iRCqtnv4ZZPw+aVF+0I7K/O0
afDyEWydcsGR9GyiypfxpoABoSS+ltFWiHTILfSSoI3gLAo/XOOzMXnhRqFI+KHx
RbExbuc5gbeKtv7PGb2ypvx/a952hUQCnh41W/nkj2txAjjLmM6lUQRDoXiEq9tO
SIqonagkifeDwEWZXkh9ooge/SZ/WhsMr7CjgRyROUBAIxdG+n1m34hx6tlqLOoe
pnbhCHDyi41nKaftjmMflDuF0kAmiQ7NQcg2R2NUNhGRfMSv163MKrkZpXmczXc/
b+YGiWGZF30L1gBD4vCX8KrCguA/fbBjRc2x9/XhE8HnOr4m1k7olv1U9AutJEDB
Q3Fem+Ox0q+iWpZP0EEHPUp5Ph/ifi/RPpgdHBzUa0rSCnPPOFF8RInAGJrJ41UP
q7/UEOjg2CYIAIlU4+U2jLmnC20EHedcvabLpilPas6WqhOiZGRtduGTFxpSAdjM
E3cvOD0lAOghD1UUkbguy3eHyY/byTrnNneg0HmjTelk+LKKnIPwkuYq2xy5DzYp
PTU4/Y+fEfIkyhqm5cMwELPNawnBm1udsLuMtnkt5ScH4odHm0DgLlbWFDD3rhEr
7lhtc2qrFwHKhbt3BdLP8tpLAjlOd7udDibx7OS/jbG2hyzAxVTYN875xltn6xdQ
zqoclxKOgCNr2pNFYhkCiQJfvgViqSBLRPLmT1WZucKiFqbxw9HAUSCDmsy63JKe
yP03QmSPKikWp3xGnTlEzi+wI6Ry7ThgBvfJHaodHUxi/5TcpHa517FDHxEhHdFD
hJjpCNBSAdNiUzVOEk4xvmI252eGhlHHBBQxvkSXc2OaO0QndxFEcqlXSlrmct6U
XMQPdLzx22pbuRyaxUvFD8pjWrp9oa4j+RMe4/0YpFohixU6+rZzU9Xxhojy/EpZ
+vuE6I3NuZA7EVroQOLFXmhumZnK3LISoDhHto/21z9oxYy6KlC3O0Gqh1JQbier
nS14y522J8KaQ/PPIYcfmniJE5DSzC2OZuRaI2FhzpJxDdMQ5fN9uW2iAdN86mm9
BuM/L68Bt7U4U8oCz+YuAjJV+Rs+IOCpEp+EyGVGKo+mlv4i32Fl/61l4ha7IGoi
cn+RWZ49dnYZvsqTkrJQdg7OpSUYxjEyYZiTCu2AjvW1EOGRX+BJ3zOjFmGRObLz
X9XM1xkQ6wbt3J4YsYnd6Ujd4SaEXZ45aKOpEibseUgATR+bWgyMGtCeUzjaJQ2w
o+YeVsNEkp3bMXlc1KRDo0wvJyb28UQk6M1wSrHzC3Lj6+TFP0knl+vXGKat4+RP
NDN3cRipnyaT/nEubeVJQYXFSdfYUFoNhsz22oVMrUFul1xtNYmR/vemQ5RV+Woc
AGDk2BCQT18yBXRRa0GL/F/BubNDGILaAJBxDBfVtZ+f/UUDr+LJpM+GzH014Yuk
WkjQaGsXTDI7bijV1x4TSCr6xidvcWiSUnaVXf8xdDWsWsOSUgcm30ZR49FnoInx
szhsyeUzL+Mw2NjYz38LRJZT7anDPc3GlOZA+6d07dUh0j1k4LaNLxwgp4mOweej
U+nzzSVO9BuTrO5Op/9HaailGKYP2NQw8W/COIdOzFE7VvlegKdL3rz3W084EEWX
9ykuQdszYx3DYzO3qHd7sNNndv+/ilTd59Iozl5pSyYV/pjxJVFgb6yJd7pO2smL
+pbjVGGTwjKq182VQF2Y8FakT7dyxNVxGivQPwz5o4grUeSs+Bf096ay7fatXuzQ
/CTS6Cq/1l74ytTlPsotGCe7fGx+1zMHccNZLP8FMDq67LVvUM5YuV9wauIrQFJ/
bBFjie4kr0O7H45iUfNcPE2mv7WdbTVZMjd48KYzitZQ+QWPKVXN3Ix85v7GZWug
ygmdv1QquJri2osoa8v/i2UYLLusOHIgKks3O+R/0Vkfua9kXMLYlVve2wyaDBUi
MflusPfkqTH67s0yPOlqNt5D9hg69ukFWscTu85pNQnYVghnP9NfPntGylm4ZpzC
OFZWDZO9hqVosrWPUTl8Ctj6flcDXY0V7rJzFX3B/9/OCoMGlhJzXXeiwysnFMi9
LzEQDEJOwQiHGSxm+kREvrxCBxn0j4rBF1V4Ie9B3iAVK1xUbC04bhl+lHedAHPt
GOlLKaLaL0CMYRjYuDpuYE+LNNpjHSil6rPNsfqFl0Zk2F1EHf3qsCULoOL7ufHr
+H3sCoorNAuun3169SurbLT7MCRjU+5SO/hvuaCJMmvDfpoBDeoKSQeb2VvpS2tI
81WgTYyQUsF8q+dyyAvPuIym5ZMO1wRjFfVv1JLnvCp4XtUNHv8NTRTIhDQGWlOS
MCF0f9ysJa8NzZXyrUMgHxd4LS7j1vENm0WnGoRfGGj1GUpz4IDsJ4vB+hHE7zmg
qGhkPA1UHixKxqBCXL4MlBbgplfCq9qa5C0PQdw4n6sfLVplH7oO+w5CjBi20h4u
+4XpWp07zRRFQDcTfZlO8ihFtjIHXT5c5tIs0qSRkkN/smiO+DPE9FtNr7d8QYmp
yX5VGy1whphJtTKyy2pedLeISjGG3SPq9OpgTtMG2cYN064zAqMoeHfOzHNkaMrM
qP8W7qVZEI6Zs9SF47nfimFEohI53xICJBSVgiUuqDmir6vNnKqFd1qqTlfZi21b
BY3QrQeGfpdEOCPw3Pg0BEgcEbr/6OqveftGNRR6U46kW/QP2Lovrysc6+SlIGFG
nIYp6pT/drHulZMmoQYQbjXVxOd7uenzGe/X5VKDO8U7TpC3dCnFERXev/tRydT7
IDAYbLNUKFWmrUV9JGx4/3pvczWfW0FfQ9wD72X6+hu21K658XgI9b8A0r/UC5Zl
s3CIcC4aZzxeGK0ErXBs75i93XqJh6WMZx5M8leFjOVyLVd2cf9VZe3En+gm3MYd
XFk/SIjSSm6f61GOK3YbOzZUlANFNtN4ZD6YbUMMZpaSm+bI4WGzLFQJ39KjT17A
ghwGMoUfPRIq6Ief9a5fI39lYoCSGAI8upOkmcbyY9OCTC9ICc5MxlC/oxd0ufXR
s92Ul9LBCjC3a+KFJr/xduCcsGY7BeseL9zLPdxA4Lgz6CLRzLiO1rgMHx0NVgme
5UPK26YUW7irKmNx9T34/HCZzF6JNTkmsGt3blFsneRLF4CQQfl0+ekSjdYIoIi8
mY1+GSb9Mj+DJHQ7Q1fulhxbW/QerKfVzo5ghDiSdHfUUXc9hEB4q60VXN1VUy/e
9GiWWJ9X8GFUZQVdkUw7g1QL4Kqfd2uXjNmgYnrNbDFGTwAWKwJFEKK9HlzLTHgN
FSF8Sl0PRrHE1ycBr0MeSukmNLoFiSQ/ZHIqV9VI32Qfvmb25f/z2Zl0DvkNkwEa
dZcaFeuNgIthy5zWGC9Z2k7ugGxRmarxCPSxLZLiyhwz+Go0rwBxIoziYpAVdk01
FNQ/CsHxg6kLXkGJXqHnxzaYQKqdz5lMywfpc3P0DTcU/Om3TbVjIKg7lOEmgjGO
NvWnL4V4PqbcEnhi6MrhFeg9CnjyB3+3Y0y0ItWCx4XkrhEoZDeJopHNPhy+XUnm
SP2W695JPFCKQ9UDjEAEf0nlaI7z47X+oi07fGYCsayUUfd5IeOOxSke6esZtHt7
E2FgA/s5ac9oqzQhlUjF/5bEdwAFQVdTZY8vZcgCwBMAp9e0v4LQkCB48hI+q8hR
UmUlZJa2GQ2XzTvedMnfDcx8ryKob5URkhaMhBIGFJeNqkyenOrq9i8vXzPbiBSn
xXRDUlVLMwMXWO9eEo3EHLdEd0+QDKbi35QG0PeEN/q2gRPxyrTx1NUSbmqaOXMs
U7i66xjpNnSKdGaSsvogcb3VanS9WjC6MfNrv8vQgRH4pkY4y71En2wGQfH9ln3c
dbbfx8KZwzVWmYA1vqjLjqAKRIbi4oUBCCj4Zx0msR+n+If8pmkExtvL5wMGFYFi
05hMYKYrFTIbBxuzeTGEJHQBJW2y8CZCSzuWmIfiXVM1h5jWSX5vLFtT9ENYbf6V
TngpIeKQhMh51omJ9i0bGlQBx9TuUDu1+ESXwAjvsRsEorGQp5rcMKvCgDgrkm+B
s9yXYnJYdUKF6QKtn59h/uM1WzlbOefZCOmpA2qw0/E3d+EsdrgGBU9ySGzz16kR
+vj/TZK6Ok87S2ChxIVgZrXr/9wZ+VjrFhAACO7camWqkQH2QB86cD3jjaHJ/Q42
RCoFYbOWTxhVbwrZTdLTKXSUtgTa4LGtKGYzmD5qfLVZG5LVhAvIXgC/63Z1w/Um
JRfpfn0WfScpkeWcFIZQGDoACS3uVkgmC7kjuAv/vJ0ZOpz0dXNfB3ZZ699W9X76
zRdTgvW76r56Cv2rZfUn7xA1eNW2r05vdgbGhy4WKfpdi0ILPj/+ddRtpKOHssBm
m5zaWmJ0uuf/bhFeD+c6YSvzkHspzCAFiTW6S/49K1Y2CUsp5o4M7l0CpqBEDons
V3Fm3Q9Spg00WnH6nDJXcjWtY4OXcOy6J6pWmG3H8OGLom/LhfGMUzgZSqwTAp/I
A5cI2VxV28xaJRYAa185uWWng/9UbQe1lu8C5E78xH3XSeJOF3EMHiegC2Exe0Lg
kT91jqKurwLqebM2saBuoFYOdZo902MW6Mil7T+zqS67HuaZSjl7UYsYPs0PaVUI
GYKE/grXBXuLx0Vp17Q72jUuhYveGK50kbTuuRLgCzp2z0PHgiRabgiXNc7QdZwZ
hKO4n6IDqla2bQcyY83ZDD1nSSVB+0i4ro8oW1stcy5DHKoyHUUA+1mTpoFDcRZX
ROD+1gyuThVw5SE3mtzzCWcWtKhHDBZLdMZu5eYdU5RGxi5LM0v9Q3qxK0yKzPJn
Z5lYvVgQIxeGkBG6ORLyD/yFR1ySRGDMzESHXGxqTDPQHH5YpT/4dKwqpIOhz1TD
VIuSQNimBD486TOMJdOLaN0IfAFITSaJkAD/5yp8C7ezjC3lCSuqohcc42sBlLAr
6EMYCodT+IEvXe+vWGBGcgzgyRi9w/jSXydZhzT6v9Wwhl9/VIJ7/YPRr6hFqSbk
H+FdcjqGRnyn2oZLKN2ChGjf0lGajhVXDbcypzwq9hZOq2vkzTVUC+n7/sG+vDYy
9STWj6E2GfchUQMXGoOnz4grZJ80GpXsDL11BI2rb5JtD2XqSvkDreRZioxEOt1l
HZTEd1aSgqmaRlsbIUKJKt55cn1JIpeQPxOGJNXkLg7k/1rtqVNmeQt4vFt4JcYX
q/2N8a7gJS+5C0vpDKnIvIl8pnT8tOyHcEmKoO0qjvZNLLQYYwPOVUkF3dOA1SZK
P+XG5rDMowgx0JPZLgTKPcp9PErs2KMZOIXc3bwyaK7YH7HgKj75Vo9RpqwYipML
E1rNDQQ+vsFabMRB/isY4x9L0bqcJlMN7jlEy2l+Qtw31ZVgUJ6qMAfaksHBh2qs
7mB+TSbBZoDNHWO61ztarmdcMno8i9NsSDiZf7xzGxBrPE7HZ8VkwdY5YA2pERLR
zzs5g0LsBoiuomcfzotLrXf39RZgX4jLbVblzpY2/vgjrQTc3Chkmc3xG3RYBKBD
8ClL1TZEA4iPyE/50bxRP0gTBHUxDN/Dx9bkJsF7fLWuUuLD9yVVLJ6HnKowImQk
LgCsMiSd5hYb2YH4fNtRAp5wKJPNoPtHbbN60sth4BymjXPRRm1Md9EKD21fmdpu
oR121Bc+QsagGIkvhqjJ3oOE6+VJPIQUmWe5r1mkyoVthBvRku0yeZvTgscoRn6+
QSX5kyjSAgbmSJvzGE3N69UcUBlxjujrJzE7+EZoCfzKqOMIKkEouQMHW5joSu5q
4w3nRsOkgq4AuDGjm3uG9o2uY05lu/dnc/DXgWn6o6cUpZhz3cQdK9Kjk+PhQwrn
IK2Hc+giNNOAeQnh5kyG+HdUPL3l9CRtrbedKgMLhJZ9E62ViLpw/5Sb5xJGSG6r
Lqp7PPc0UwAuCTH28ey02kLfOgYNyUa68qS0sBGB9BDB9GSWYF/iZI4KV4XxP5Z5
8aTnsDbJL71yZTBUxWL2WMcMQYT8k9D51BJLa//Ab6Z/Tj+0C+57wAmlPq9qYstg
xrpv1AoaE+2SVDtjthOe6IaXlGluu8mZTN/nDGfBi9JyF8694rknmfhXPo0KHqsP
tydxIjc4YyrQu7I3eYNeu3MGTeIJPqfbMweHAI/+BwmF39GLefUj3YOKHp03YwaH
tVFUKvuh4/thhlxpr3VRIuJOgcFtJbcXjdqAOlKfS5DBocjvez6MhwmgGhNQoQmY
mE9lhZzJsniMcDImisHvBaPapGhCfcbtTdMcZGaN62ub34S0asRiaelmVaDvweFs
dQu1QPzgJ72u1Ct+Z8gZ3pDm/Rqb18TH7/auHwHyNtFM2ohmn95VJ50vb53vIUSB
5N36c2gJjc3Txt74UtvxVV7fym1v2w8u+3VOIVirnG0yAnQusHa+sdu2iDsf45My
1dexiNv8k14jhTE3w26PTbhEp3dai0z0dy9g5HaF3yLkUjr58QPoNqhWIV/KpyLu
1N7avrKAG4ouu2kXhly0rdm6p8DoSdz86TIgQor8ugXS5K3dZOHkLUhHwvo7+CC4
MVANGG3u7gWAV3HkzGi+JTHxzA4xaBwbKj5P1hBa8swb/XTUQZolclODn89PsyZi
VjFX46IxgCWcO9oFA0D7t8Sb0YeA8D65jOkx8HZ3Cy6gGVfDs0O/sXswV7t1ttGi
BdkaRosPqTivviFK9WcLZKQMounVo0bwiNjz5WJpkLfbnf/kZ1Rl01DmDrdHbuqk
CSfTgYu8TrLzxQ1kIMpL+5I36lAW6m+QMEUtoqtCYfA1LCwQMaXYsGIJBGca5jGt
CKpt3o3XTnY2nxazN7lUvUj4Ot5of0c/s2dWsN04mqV0dQdT8hQdi4J8FSHqilax
m5BZIrJ1EmSvhYUwOfZ3Imniwf6Xhs9afYWxdWB1eywwKudY4XBxohW+Yf/TrDtT
KC7G5mfICNMkyhOmLDPC2FOeXo+UessSbpKiSJJLo1h3eXFLGVg/rPN6qkv6tD6u
x5mMUsfoXduM68zw643COXzYWck88szYV+Te12sh23oc8ie6oO82GSZaSB4dYPpI
0gMs2FBsdWXznHAiTGUdyVa92xHr4XN8bD7vsBszECp/sTQ9Eq65dO4K9F3TDAv9
KE3k9tvjEmoprC5baZZ8uuc35QbBq83ua8aWXpeNrf8mq4Wbr2pURIHJ0Df4ab0I
yVFJHIIXSDQwKgEVTf38EOxFUZwXnRgOLX/vQGI/Qcf099jA2E6HVqqq5DIhr/6M
ZKcgvKzZD0szsJwlWYYK2Rt4RVG3ImTPsaStblA4isE2whGU4EKGfNDWVvGbBWSf
4wcyjDQboKXOdrghVRzVRKX9pPEKqgJknztqDiHXnDB6I/y+AMY8hISVHWWYklmA
8G/XbPTXMaTG56XNQHl631tKpODI2IhrTeUTQDGmYklbhUplYFYhkKoCQ3DWWLkO
xoZk1CFzEerDkfv950fkbQsN1/OiDo6/OxOZNzMb07RNgtqeLMctk48/ntg+sRE9
wAhz7r0XPYDcPjYj05FAYrGnIP7bOWMCvStXtnuWsbLzwAr6Gv1h+PUb/sNBws/D
lYfqPYqFZz0b0DA1VOTULROgj8VQR9UjDkF7ysri19nt1vjjuRtYyZ++RBiuXrDg
6qdU+2Sai3B9SQuUJFH9r/5YWgPpN1XfpFNquHC617ceKN3fwDt4kJEdsK1DZcNP
a6lmLhxXd6+PLdUKb9JRXYOXK5xwhZismZ3VBg4Xd7tFEmxRVEBAMGdQKNJHpJOH
m/aHlG7F9bwLNvPV3BoWqMTN8vkRDBiD8pzgOPfT4D1lTpoIKO2l37QgIMDP32lD
PSh+KCbBspis+BqsvG19J8wgFGFkcjEC1/XGhX3SkNneF9KVxX/cefXyFEvc4uYK
x4WTnNgpWDbSWIFU6gSW0Z8ZYywrXrXQ11Zj/KUBhP1hlxmg3W4qcjdauAeg0hHk
vJUUY+/xrw3LLMW3ao5HSkh3w/lHqkLpZH+GQRm/I6ymhSdG0aTAauDr6iJ0oODl
xOjwHFAle4qxTVoLfxwlY7cgZGg4Ix6ybBIlmYewT+YtBDZ+UV/tbRr05QDB+jtt
yerVAOZTPg4HG8TvjRz5Wy94gQ1Sjs0MU6R24R1aJXOBB6ynfHPRSfGIitW4suPi
S12+j84gXE9uWVXgkzAWK65ec71Vxo/QDTxJe8lMZ57jqrYg5qnufRYZbYc8imDR
pihIReKlPBjuRFjhVYz5iUN55IY0kzaMg2nmIOSw1KCw3a2A4QjIHdbLBAU0e0ZW
+5a+7TK8dZxbMb41g7kdF9V42hZlSB6hDvDZ93oZnhRUd9/iePrcSvkIMPCRs+3z
RipAqpNn8TVkgbody3xVXZjuXsXCRtAJd4TQfMIrM6NcDx3//Jcg8LYDSIHbLmMs
vmIUqmCs4QMjrtqZhi8ChjA01b0nOPToqf+YkDZ6pjdg0RKf5BmKCTtQy/JHS+dz
+tPk/EOQLxBjJ+sMWKid5mf3D0XGiLNNZMMwVphPVL5D8El96bEWhU11ab6vXQQa
0hLgcns5csr6IlLQaIXqrbgPAye1+f/5vFgIQKyZiULXSqRzhQjKUmNPgK4Gjt07
DeUnXN3rmepOT8OKAPl5mSd6WLdTDSB5GblbAyrrdJzJ6HxGHEjeZ3lvXmYDQ8Ew
1XErN5nkUZX+B6snRkNTcSCFoYwrsVXeRNqMZ7i2nDGkMjv79gWiA2ZtM0g7B5Mr
5vfRJZgy3J26gqrXIdgf2WwOB32WuhCmPfdQOUZvZ0cWSh293l/crw+1hI/xwpqp
JreblaSopuD3qFl8wJRzmEz6QPmWaFpoeVozGwGruzscBqCXM7YCcHX6e/dlkZrm
dB3qhLeQCykBdeA+XIWFaTGqyX7gw3Csx8mkzXAXkZSACOg5xIBsc73Ox4uWENE7
QANZsz/6gdvG/byo2pqGGVvlMqWNsR6mXOo8h8znejZTsIRKqS3zab8PjZVyb+qG
TOBE/ap2Gca1PL0NOJtj5rVZgXeNBBciVruz4gVhN8EIl30pXAu8CBhrBZTO+nLD
WA1HW3ZEuT+r9gCsibiJ86eLP59D08bqzu0gqDl5XR6zpe/Jix8Dt/IozI40vm7g
mlSHfotxT9GFFI+mQmnTiOmwo/NbA+7VJqhwb8qB+nL4CwBbznXvWC4sw/JHQQnJ
FPr4ckfH3pKCG8u99XA052itchJxRSEVvKlr5j+/aK7P0wfyiKUcyphKKFYVP3fL
gWjvmuPLNIDwTjtDuPufLS3inTNCy3Sj6y1pqQwGEn24S/pt6ngsyMG+maI3rTwi
5Qcya6I3y2nFj4ax8J+wMGae64HDyKI4D68kKDP9EWlFG4ZJeD/+5o39vm+XJWF7
eK5VlO41SB9RpK4GIbKvPGUTyuiU6D/8qByejvg9zGPDkTAawAuZqw4pWsS/37mw
5MD+C9Qr1TOSXM2l0RTSzb3Sqv0/S2VUtVEeXyak3CL3sY2XkrN5lcPOjHvGH3b1
FWUaHyVmorFw95MefeQweDtK3Y7w2ROx7Ta9ywvdU66glIv6TNk+TtzIx8JqFnHj
jn2mvCShiXqBxJ/ePoVggdZ9ZpoCHAQt5kBW4sCI/izHIYTb6Bi7X7McxPGTSwwe
BrGle8LjMgTLSC/715YfFCERKIYNmZiJiDIG+2iCnorbBxev+KjOf2SLwDFdBi+v
pXnymPLloyCx0RYTJ1aXcxoARE3nYotcFG8jJExlyUqV+hk0rt8K9o67kclKrK7i
W4HlVvTDOUazQk2CI6+XiuDmxrSGcHedvYhIShULXHKB7h6XNbaLYU5nDSmEe3pO
z1IPtjYxBTvioeYrTNAu9LYJAPjcti1d6tlfAClutdnV8lCXaqZDtHJ5HrwTe4W/
c5Rv/GElnBca7wQmU6cII9Q+sz2XxWistE9FXyxg5p8cy8KMYcf/TyegUrI8YZpl
ApR66xTOEsYqht4nVN3BN9EKeNgV2ej4K5J5rSdeWN00BDWj8D1jqDGv4arab0Vr
vFTHLSNlQ+0hRqfJQMEsUsgrWcs6LNxStCQZAU2ITeCgEUuAC8ZIi2NNRQe4OwkD
BAGoB2a2GUbMAqGK1rXvh+CosrjrdYMDmq8Sg141GiHe4LuQW/wvGNhmbFOAsAdw
ClXVnNa16J3YJy44E15I/W+l8DFaOJ4jI+9PFING5sVxdj/fd+YmEUCdwRyQUpGG
eMPCwT0NDUkY0x6FVKdIymN6L7bS12P5NeN6fOoVH5bBDsKsE/6FtpcaXy4HIqN4
GLVn0uTYkICdWJ8Wa05q4qLJ69m6KXIL+dIb9S9NLeJUKCrEqviN2GMQPKvO6qGA
h76qiVRpIZjpih8GEyhe2Y/z73sTgQzz69nOCQtXYOOlDRkpU70Wnn+ItK/G1APc
rMFyOaeeyh9eK+14AyAmADuAu7t9A1/zx14EyuaWvukwoM/w4MxPcNcIObQb4QE9
MUtPzP9EJYmx8q9iJmBdgSfR2uFls7VfQgm1JydWvsgDflKYdNO9Cy5iZhoEZuZ/
bPqPkkKG8kiqV1b8nNDECnm/q0yBtqHVPJcm8/9XfDgFhRU7rQ6f3N3//7HMiTq7
5wuMfZNHpK03vSgPEAapq6AFOX39zwAYhAlyzdBoroz1cLNC/exQA1Um/l3fP5Mi
sQk5Ed6kk5JFulW3+tIOwXZINf2T1Kd/qxcFhgrr0VE5maP2+K6YPJhZpB2qROeQ
Za1Xg1IDJ+Nr006lS8bemCFR2+M/rdeCohSqm51TCtYn68bmDJt1OncrBt9GrYPF
wWNiVLiStUYjcfYdxt8/F9Qo7FgcuWia/2oqoedWFBzAdpX44iET/InfUi2Sn/fP
XtFJ/XJg9xXmIVwZuYYCpz+9zf0Lanm2vyvSwIaKX5mOvXLATaMBgwIkwuFKhwFy
sOsNzj1sQDug2ipp+2bYleBeyN00jNtFnbCokWIXol//52yQfSQ4jiGlPn0Ut0+Y
fXb4i8z6ALFLWlXajh3gKUKdEl+Hp3C1zyh4IMTczyL3ze2pELbi/Bmds8qReBCH
OArayWY8p6abp6Gx4Dj16u/lnzNTbf0JxKERDNBfBzOvDR1uhn0mUqk/4VEdAZbT
Ez3ZIDqCIvevd9IgZcbU1j2Z4EyiBzLMFfhRSFY9B5VroYN4Hzppn8sRX4PaZufD
f9VLMkVrT8m9eCdov6b4UYbTxoIGFD6u6Rt4Tl3ieq0haddLCW+T5bvTmmiQy2+D
jIlaTwM4zW+KYTs8Vpba1EGrox5P6kwZZA+43uqhHfmMGX06nkQqovgouY0qUVdM
SNHeaHU5ZuC8YyWGPF22arF8v8PMSsZ6vPnTfvGKjCLTvILDXOSQx33J+moO0BFA
snYdV91v8SAJnXG/9ftUa4nXvvWWkItKSNjZi6ui8/4OSQDNpJ3r88Ro4Kd8SK+N
rub1f2AsgWes5Df8D9t4V7cgD7ct7gmGEKNVTo57OPmuDCxEY11a5+lDAs3ZPHmv
Jncy7E6wW77EbmJv3cE4fxnS/u+9gYshv+4WpEAi/7w1Kma2F6W0ORvyLClLuvlG
awSF27rZnDVxMV9BvWek9vtO7Ey6zurQtu30fGJSFqjQ0sXFRx3VP+GErlJmOjdX
0HPVxu3TTNg3Dqwlq+CqdSsrEyj7mKGes25NriyayCI7KdXB5ots84cM5HilFOxi
B8R1bmFJsAEbGTUN+7K94RwpbpSjVNmwz9K3WetsKXT8nZquct5deORLoOIT0awG
u8CTjc3Wkhpwo1hex0a7KpM3/cXQTUpf6hodaUXA/edP/Jjf9CY4axs3xOELZe+F
40MAG7hWa/lHb/WUTevW+mKwIqAA7uh82eJ6Hei6543YcxrQhN+U2d60VgZuhnav
IPqA4wecJLm/48M8Y7RWSuqH6NxM1Pqox1C8P9A3ZKfwJxywqDSC0ThwK0h2bNK5
Ly83AYCnvXqYThosx1Pj50h+csqwePsZxzAtosytDr5TRxEMANBtydzOXqlepjuN
5L8yPZNYwlhKg0voHt/SXQcd5OpZzV/Dz6ozVciIZ0TGpqY22Z5wiO2UEt67zn0G
J04GJNd2yxfIs1hnshUI214r7j7lCHbUgYmtQKkZyRGZRAuzT1hzj4y9AZ3nYe2x
6q1/9zrTpA6m0AlsvPYScEgc6Ag/MHYK8vHjdGZywJXAAFoJzcJI2jtf9Phodi93
ZjjRc8CY40bZyXs5tYUGD4Dg5QW7V7lJXFaloOf4JZxfR4Lm0Z/U9HXI3WGMVQsk
T3FPvapkggGv8gy0OieIl2J/VtLdvMZdf8eZMyYxQimTmVSj++7/PrEOQ2I2SQrV
57mKqWmOfw2hXoE+siGT9dfayxtB2CaKI3ctIlWp+UfSuOabtsq8UYt/IW/lwizR
NkY+QCFFvXdYH74FyabdJjaAuSX6IOUvC1g6nqDk0e6pJzKzO+8nRdADFHqlOwbF
MW6d6mcpJlTvwPeVR19u7X/cNGC/NsMTELDxbRRqYU40hCkcQ0x+wcWslxII0qlR
iq640CdjZTJ+vh9ojtIsjMxEBQRa9X0WkTf4400MU8IucU3s0cLDvjM7ApBU3cvi
ULJX8HzkZukrngNWCXKqNsEIRBw/C0ZVdhuwofcblW27E3FuYyqVNukX0qTOpXTG
DWijX8Qg2Zv+hC35LTpz6u7RoMlW83BfsWHM5BtZgO3xwFD5lqJyH+MxNKYIe8t8
rM7ZdDrmw4/igR04CZx+tFJyKbuVFT9JS31VS5a577nL98jlYmqeV9wws8OVyFAa
G+XwniKWJDrORu4qcS3S3u861s1gIIBMU5xWHfAogOm9/U4t1JPRoX0DOhMbilGz
X2c8+A7u/HBQmdwLgNBLk13t/+8ZT9QKxn68jYWhMmY784R+T80o7fYF6pOpEVhB
F9T3eUGI00xjeRDnf3VxM4y7vPcP3coIrbqGXhWsbkIp5ZWmXVe7X8YyqVnD8XMe
yqoxmAYQj3WoqDBCkDItNUcIvwNEPZ3pvekvZTCdX5vkwHYdsfHSWlu3a7fKpSgY
tbPDJeMLfuc5LDaLDG2NKWfbBmeuo5LjiwLnVYD6UjkcuojrUUinNH+BjjQlS4ES
cg1fgHUfmmXSijNqO6o1YCPaxw+ivnTXuWzMitBcPgWlwzrs0KMseYfTZkcdLasy
G1flKH9LiLjUScVaOKhZMPkY4Zk1K6nn0D9jahutW1cxqK+jvxM/i4j7rxovfjd6
Cd8AIp9YtQTPeHhzkDzqbj+fBr2fSCPcQ0/S9aQHZ0oCagLnmqGfI1+Yycx01/LQ
3utnRmrwS26PYvw9U7RK7OhmCOuh9cD49vGlm5DXiFzwFvomFvM0+6FWqTfdQLiw
lpb94baWiYs5Nd2J5hucbhsK3KnZSMFg/dPyjVW/YbTR8aa0PSRE7bg0/PpCCsoj
YNo/N7r+ciNC1ETUH8DnrWvH8S6no3n9+N+UBij/C2qWw0uSRwAC3UlSAYrltu7O
HOL5V6qWMIGuITjv39BtfiafwxPH0EwfGK8uXJ1k19yTDLvn0rAjH4f05Vwy5LKW
2hsEk7tINp7YvQATLLmrhey1zsk3kmKXbNYC2RoT699kbeESBIjOjAHYH7ZCQzkr
UxrJuOenBooZ9s08c7DuMz/bw7pqhhrXhIb62Cp/8X6gCsOtZIxrHcMSrIyI7e/r
ujegW3hNVtNmlZcse2TS3NarH3Hb9Qe53/xsYIBNqYpcKFOxbcodXsUjPYwOcWIV
VQFHsx4S/UkBlITEJvDy0RcQ7e8vkesrq2oEkQ3SDVsVkE+VoZ7+2bZjS0O9kGeS
QDgVrf12YP6U3IiSgvjIhgbU541ep6Bt8tgGQWya6RrdeKP4fTrINrwu33anvHVz
REq5qBSoqct57YTu+8OUSSO2uZZ5sj8pdT/AvjpCBFUZslu5J6P7nHmBGoThJMa4
/nTVdP2SsEnNk8HcwjHy0fIPHWLAk6YCs8NeXWzE1u6VuS80L/0nB6rin8+iqZhS
hwPvuQjQnolcTlx0qaq7wWzDj85h7TP5xszO/Y9uWgG+E9e9wDJmHrxghd3XREDV
PD75VNu7ORUBFt3tXH9p0TX943EzQa82kXVTe/tEnpWgvajNksxJSOkkiGWmvzxj
w5vWfz4UECt2UsrLC7QazqmkZthLe+tN0UNYpz31rU+ZU9n+qgIsOEPFKsTe7+hA
8PfEivnAePlH2q4IN2RhHMaGBsG1NJ39PW8uCng/5kDIRTj/g0ZqvGIXVo5oP1s/
9WeLrPBeCL5bKc/wdmYxJmjNwZwmK+0avmtxdFpKnWFJOT6de0dj6FHEithmigrr
yhrFaaG9aZaZyGOP/vGtxbiG36h9TnQAU8f2/W2uaFgUduISOIU6Hq9iALcThBjP
FMP1xCg5sgYHtCvVymfNkL5KeHRyM/Jfp3nVPDHRKL7slyQb8ie6YLfBb44vu8x3
dtQWy1Vo0kzFf1Bg3uSp/ga9x7kboyA+WGYdC9QJOZojMv8Algxr9B0fiBucukZp
wevifa0RogZkJDtwa6z/n3NqCvyy11Qn/V+yhCsB7RL0nbt/hROzc01tViEKx6cU
hJa2kwja0wpOSVzD7obTiaDamR6x1PnFrU76n2qDAKbiLGSaB+EhdX5DSV1XjmZ7
tT46LOe6d+q2z44gaV10m5d5aoTfqzJ9s5Z+eOP9AzlSD0Ggv8air7He7rpPdFo5
/tQ9DepZiH78EstVC15qI+4vTDcEeGpho4nQL0q5YOXw+OcTm3p0tfK7DHCZkSuw
rLak6FKXTWVj9z015i0svIbX/Ya+GNTzyOy+BHsCCU7m9VB+XQvqpbI2LEHmoltG
1ePXb2E2sJuh9X8i7mWFS+mGvd0Px50Cbegd4vIYJ8wbOzgzNhyFm5dfaQx2sYlA
ATJPETif7WjY+Ac9v9MF0IaguMpjiuDGrhtJhPmLgU4BUUu3hSz/e76HLHwOTpuq
zGXT7bOIQwLSPpfQcGe0wqlokGMWmXocTYwUx0UKPzu4+yZs0aWIXOIvX9/yAEla
dz+3whxj6o7TAzwzf98IovebSObWSXjLRBMPUNkUvRX8P4YgP7YcPhfzeoT57NsH
KxrAKWqbzp44Rx9OcsHwgQSXD8nan+N9ytP/TR3mxI5WmvRmvZoTJto1Mk95IQv+
s7qCSSXwkPaE/sBcgZkxefk8OaWpBKfjP+Q9PS+wkEaxdNr7+WfuQMXgyxypYiC/
SA8pVdBSiwAbeCLL23uQd2i33lr9Xi1gAQWZ/hbkEoH5jIH5zGIIMP7CB49dsDHt
bUsm5lTPFJcjX8BZprDnSH7xA5eCBCIbcSWKFkDhIjAWjPuHzPuKd4oPZBvCE2SC
GlqLR/bH7Uc2CKopnYZc644zRw8LDZ5RWG3964uDhoCgcb7ojrd6LA8h8ls4VwCs
vDunJT8QOlxClwUT1p+3VD4PxH+L6/APSWFfQNLH2B9iItcqhMiE5oOo3CZydsyO
EeKWdrTViqhSGZFwNQNxfOlLQdyv+l5ic5XSrHrT7Adg7rDQNcix1UsMpKGT2Kl0
rJBDX2mirAvDv9p3yVQ2v1d1NuVB88EpdCdygAZtDVgiwsFptqTjZhXcQakhZyh7
Wi6rOViPNabP9uMEdsbp5m11r6DG02U1gsU/2Wis91jITnPyhsdowlZZNOh8lTDC
Dgo/J6ZmtFcyvpLKMRYuzdF+CEEq7Goko3Pywe4G4aHSFh7B42/QTEjslfTM4wDY
EzyrG2MsewinAiE1e/6ds0ancCaid3byFR8UXHG0ykFeFwX5wXS89Y7jeL5knNnU
O4roqkaez8R2xUeW/PrN/qENrZLjWe1vy8EYTrgbsIpD46pRDNbkS+PgUxj+xk2F
tNXlXxHaTfupakIeRznr+5AiwaK3EH/L0Wox3rynBkkSnlwbmr04PTS536PHTMqO
qwMuGP9zHJL6iAPIKbDRc/Bpu+MXWyJHETd7DRzHkngvDX3oW2F5N4MO57TK1MQb
uHsf8doHz+ZDEEoB2tWnT7H9Xl+IpIBF7ien3TFrej3iyonnn61Oe5JtwzdS6sW1
GdHb3AWo/6RGPKJoJQSIqEBSHD7UOdHdTSMiaV6XbvLiG9WDepSblseClwxw1vU3
O/Zolh1LDejsJjsxKCUqJe4/kP2JLDyzhCgZ5cVSeNcLVN8oUWpuzy8IVXBIM5gp
HrqUBBx5kxHv98h5szfzQQhkulou1q2Osuv4uBFxaJlIuSVtt7fP3w6B0Re15ttH
K0dg6lIkHpAhfrrN8ZqArVCsSJCYzVP1bpywI0QPP1QrrF4/JHAzU9O8/6iIdiN4
IS8vRU9qJjTeSfBRW4coyhde5wgU0LMJZ32d/Vp6B5dADVyIb+hvaABNDtMMaLRL
L4vUYs4viwKDOBi1Ole2kqDac2C1YS3MzMEVbFYHTgUH1QOEEW/KITFTq6Ws4X4S
PE9xLtCWMKHh/oqsTM9194huUXRjZ54ptviJOjA8ADOl2ehq/SzBRNMamT+5F69W
nT8lzhGC6IaO0EMCQIWdLbyWGwzvD8bxHlBqKwhkmPTSzFNm6+z+G2NHhTBwwkUw
FZjuAs3VJvrhBN3Zpfa8Xzb7qELGdP/rZnVZHfRVOGyweg53pr//p0NlqlprLEBz
Mn1OJinESKvDloIb7y3vdZhL5hbL1Dt8w97FOZV0jITRL6LRMg0YfQ2mRswqqLKG
SeGRj3ZJbLhqgJE2W6Pd4IfPfjCvGzO029/TPg/sWv/tvc7+jJ8reLt3Gz3TTKxR
IdAbqOI7Nkr4xVqGDdHrYQ1R5A98KlH2izASsH+Rpm4bdxNeZJB4xTIgryjbcjg4
IN2D1JlwMdTi/Gzhkcy9nCa8S+OmFJqwtTXD/T04qdF+IPWu+LuYHGFC4bORbW09
qO8e2s1IYJ7AGPZR49mKFtKwz9TYkjz6bovVb/sBQRGOblWojpIByMeonsl19fhp
/vd128LgOBANOPR/M9+axhES2PNdT4S5eYLlGKBStb4FlOBuNBLenJSAvj0vBDFM
g9EkT3L0fon58V3rBPBuOOw9Z2Cl4qnnl68CU8V44+i7g5StRYg6rgdDhxlwaDWl
yslFmkp9JvyIHMcBjsAziGHgFmCBkUh5G0/k5Mt5+FjQ/isxmOmHCm6q/nmlRUFW
3sRMA08Dk/s1QUg27oZmWIjVXFgVdSSag63ugotyRqXq2uKz7GqIMf2rsARovXNS
jy1ZOP2m0/Kj4/BCdl3lzt4qe6PlzZtXq5NO5fm7oNcwMr8X+EOJGZ9k5Li9fvbc
CByKq+9+n/JWkMzoje/VDaJr5o2PkbhD2e8pGdSuYdSqebj8j9if487cuVDC8jC3
7RsqjnTkoVqHm+0h7Pql8eWAYLgi2vnDKfV48aESY7JXcKt1Ns9x8Q0w+Kxkh/bh
On4nLC+UxPvUJHOqDQSgWlmhU0O187kYIbA92GIt6DVfxp9DXpU1brFXAFYthLAJ
9B/+Sqte+THJimajGPxGMxu3d1YWH3fCXRmLSLns/mN3EBONoYJOzkOnW2soXCf0
4Qt8L54U93gLEBbIaNfPsTefkY+JFrid+ySYNGORdwqyONVGiHtj00FoKcSxofAw
Yp2hzdv9YjYcHA57IqEambn+72jzXJCeuEEnsPkh4uPc495B8QrWIgjkDr+wANDQ
aoH+uEIAm/hudFTQNOrYrQ/whaCimGWyvqHm+wwP+C5sgdo2HgBA6emLFiaDJc5l
XzSfH/37zRWAIrvKHTgLh+5XVRzJhzqPzTt8vboqluDgHaoxFbcAtvpe+nRd7/Kk
NI22c4GPU6/vA2B3FgBCOrBb63v9pKMZEJEnrlAaq8cm/xGu4XBz6wqdHy/YIbVB
L8K9Pnjid0HbKt4sY5cNAAlQw+r1lEAFgzqhniTpzy/TIaY/LscbliUfPIabYhAV
Zkd1+3QF7TA9cZSLAQQ4+9xonMFtDvE9Ez0r5fNpWWNBWt71INE+L1+A6W02YObf
yFuLsXwiNyODw0v5xAP5VX4bARg5zBE5Vu0q9B8krUlcWDnqQK9XL4SNUQ2YU47i
Bd6SnjvXZuDKhdDcSniJKZS26UJRcbBdgH5Ypn2//p9zdSqihEGKE0m2NSI97eCN
N/yKULBNe4pMmHGzs/75Afw46ww6oEkrMKFD4QwIWjggDyddxGbXQU0Ir/PygRaL
dBtcX3OdqsXiPupjAPJGIXFYNf5aCk/abqtDy/IeqbfBvxZes7776yFoTg9qqjDH
t9OddgyTLH9JJ2Z+fv39g+rlCZLKDbYZl6njahfYMGy0hh8rl3U1vkrALTBg55/p
JOOnHxpxDptVwcjeXM/+Mx3IUKHQ0Am4dQTH4mFv80iFQRRw2KqMxkTjQ848GbBN
bWcDlbeSzZsgKlAzjR9A1gKtNBw9wthMIqlcivc2ky6oyW7gYFVJqspL2RoMP6dU
6fAwLVptLGa7gOqRYFYbfnncRRlb7mLZd/pQfNxQOb6W2Fd0sEZwXuqEzQylG0Fm
YIVssq8spOrMe15PhzyGazfeSRUER3wtWK9nHQUJjIYXOtY/egV1mnldmeyDnLJ7
M6RPfklGW9Xi2xDRC90H/lL8pTacbq5HWrFasHItCCwIUz1r9IzQXm/HHThhgEqo
ieAL0QIghL8ntd2sSH7vHmE5TLwhvd1LWarUjTbCspSAcc+KT0ZBvPwqZfpx+Jbm
kKCpAAG758lb9jOONe/1cz/18RBOVzBNYGeSoCZJbpO1xqpuNCcUPNzyyi3SL91P
NKeirRCpN/2copbfF+dTa9IFpiRJOp6L/K56gdFB5Yry6hHxey9nEympMCGJw7/Z
5/hkZU6zfnI4oiatoZW8F+4eIsexB4fPxOIAoW/4rpAW1BN6Ux38S4UoVw6jfFDq
pwhXf0+kwH0lGyQSijO5v3h+h8r60IgEBaP/9L31zYmrQVmxvfooqls6XYLQpPkK
oKd01Cju2lTTLxW7P/gQVkTdlXh/y5thctafgiRFoUogiBiwdWGbWnqhNP2B31Mz
243yL4Oz/O4XeowGLHWNV/9SxFLfpwZUdSktucmt3aO/zYWsxXM/9se3Xv6/mcAP
wyi0FAdthBR6vWqZuOOWVphhbSxSm01w8XrsooDllWCAecApW4dC2+F1rOho/Hzx
W0m4OjZeMlTwmOy+rTBklF43N05EWfwp6PQWA9wrhbK+HwHDTkB25Ugfss8YZcPr
hVcGhpYfag2dwhHtEdZm5qlfUTBi6SsHXdq3bG0N5UnTVFEMAEZzHB48z1y4s/mY
mlsVoaBmYH3rPJkda5DEh9kUih6R+aummHsWnf11V/leLBs6uhZDSaIPtoUz8FDg
OdfItqdenRdIQLEY79qhuD4K55yVI/vykPFmaaDvA1I7+FIOCX5gpSzsP1PRpbO1
b7nVnP6i0sgAr4Nfi7nvzAuIyy26Jy6bbBjW199Q9GusAGYedBo/4ShFVolIhlgp
d4/7t75BpF2jZEz2SZgOtzQpqmYoUD6NbsBImAHl75fCs6ubiZ0RCG8VCIBMTH4P
32LkFFaOrH7yUR421G5GDTsgHFrr2UvK2Erlaf3oCUBxZMVZPYwntXKRP0PWctbk
aDgWEjhtK7/pA9mTu6zOsERHucJ5QrE07izwLAoSuGWBELa9yYMbzXg1JAlvgiBQ
thu9yZTmsoFHnj+WQg9MItqTexgEm7oHkW2wfpUVsntiIVELQlYdn54DEDepUVsj
/0auSunBtoLkYPuTX3URNh+IgD8iw5b1gEIasR/qfkkos0ScYmFrbfdIFdxlK9rf
Ixuy4MaM4MWsBtl01cCuBEzCjVV/qI6Xpjbxyt1/dR8OXdUBg/A84ZFOQosDXD4S
yILBhUo+oAXs0AfrZCfLTOqwEv9b5yDlrKePB1cD1Ql+rsoW64y29T29yPQWj1sR
zG83icdHlGTRvekNfmZDS690JEO8BGPcymm6a/tzk510cdF+ifeJkdzvrbxsTo9F
lgI5nYaxrDrYAM44UyUv/zsJrQWgOA0b7/atGifCp+7JWtj1urFRCCX8sketAISS
21CDnDFcUAfeJ2uY+0/7Fug5xWiyQEAv80s2gO0OX2Egv6ea4WF6yyusjh2k4rGK
GJC4BDT6LGk7vv84g997CXKI2H/xwFZ+2j0AXhUkS5reOzJrXygtIu6W7gHirwKR
lEXTjTfbclCrwIIdE6/15sJYTfqNAX4W/jB84CryT6Qbzv3aVJsI9S3Ea/RU/hkH
eOBwdGh3fIt9L8SZfd7noBNrJOL6cEOCnJ0CsGaejNOJmKFUVKRF6abIGobJ6IhW
VuAwMJ4TgLjSphAo463soC6rZfrVqAsi6+SWDzNzJJ8lyHLDw6AqIZMKgbo0YZ4Y
32RR5zWQt7v2rIevt1tCLCFVJizoSOQaBi3zWzH1UtbYCz2LqX+MVJlvoWTZ9C0t
QFRIkTIhmrCm9624izrKz7bmVUMAlj5bwZ9b4IncyreuvF3dOO1zt04zNag485iS
FEyQtu0qUgq68EyNYzu9w8CNyPeC+48rmJEZpk4EEaOs66q0UCdtDVl4hifT/zhY
sexzsWbvAVnTx7hwtdpoJKZaDaj99dsjE8owfpwflhisq907xrvW4w6ZnacgNBWc
Ne1R6ZRVMiPjycsHNcJLvKZBEHzXR9Cme6RjzFubcb2fSQB/fNrI9jfGDdjWihj3
8c2CIOlSIHwRHgG08QASmk6P67Q8eP0v9/OE6K3DiP1IdTZ3t94i6ZOZl4oZOTS2
k7HYnGhEWHPojvDJqpDAP3rh5qsxpxK1SED/hE7G1UxVy0Enb5X2Q/TVIaaKmakB
JCZDWa6Nni9r9Q7vw6scp8HEd8/8GAGRRE116cnId45wsk1XC5JP2sQw3SSIosQ4
FA7qoMVdf1tG1iIcWcS11FJgymuUsX7ih24g6jw1MNumYdWTmfIK8E15O4d8/xjg
xFV3Gm2Bkg7UM3P1S50IeR57Wu9M6ACnx3LRVsY8nc3H9F9zmzVtflTGRZFJ/jc7
0I8JwHQ4U4v+jvNwPCnJjfdmanRBo9zOcca8xqoiCeIsbkH/AY54a7uc8tb7bX1V
c2oKqjkEJbXbv+XpVye5osNpWvVPJRWkH9LWeoLIfjDMqQMSrNwEv61M1BciI2ZL
5LzJWVRSn0YgZFm9NpODHK58FVSFXuoNBKO+MtuCJVf3ZliUywTpuOU6K+WyNiiU
JWtJsY+TZwlU8i3DIyftB38o6D2C40eKb87k8KV1isdKcxjyoLjD3FC9WQzAFAA/
m5Goz1G6td2IjrnexWxUogSkE5yjBF3p262U8PEezcExkR5AgIY3HFhHZ7s/rZfz
IPtt/YgzeUmDx0R9e62odyszoDQtZmX9CekmQLETc2JfSlvlV7cJMBU9CXxqF6Xd
ioiYrItx/8MODpy3RyHCIWN0fRub90IyuVIvoYXTL4cqDxEnNBvwCaQ7030MY+a1
XaPZQc6S/MHoJOIipI0se88lC5SrnnKUxAr9CzE0cfzVqVaJgoXtS8NDfsMjpVem
JVUg9PoZqXMzXuUhkoV0/T0WWP+BRdcHqC/0KI9vD2qRb7fDbpFbsUmVbvo0gNQF
WwDHfy0Kmk4GVKYr51N6L3vNGfJD/cg1JyRKve2nV8dzeG9lW3Nj6QYpQ6hQdWcP
Dw5c+BhcKu625ECyZkYWfeAEbXnVZW3KVofQNPPMqq1xz1D3vjPYP1zr2HFDBDjH
0779suDa96bAmIoNp5J8GmWLhIVCiRAtafGR4tBaO1qDG/Uo3+IJCbAtCBCz9A4B
ScSZIgv1LvQzZkhZ431bayM/eWiFupNhQJJ2ccjX8rYi5SllMXPs+5bWKkFzIE4k
CI3Sw/O9xREfDEwh56V4052gUzGBuw0g+6//BAs6n0UZA6UesAEzP4mmO3JrVVI/
nuff5I1Q4U7Ot/4FFQ2IMHjMQDxlSBbpnJyDL7RAvX81ZQvfYYjafSNGME9l+nNH
0gxZThCm5E1Aqlfpmy9T0txq+NtuGlKgnh00P3V/b5KjYroUbV8nmgcNoXcOaD74
Gyxy8lR2iXuRW3sEuEcRlOhO8EeEnSGbdYdTaGdG/KzyfO9J01T/MGVxN068Zl4I
PsdJELK/jOe5Qv4CkI6faFLc/pZe0QWbQNqQACi25wZ6IaIll+eR0HJmv4s+Dm+8
PDWMhD7dxMo0wUUXbMnl2ueLoD/T3RHKIptkMuXAkrlzYkn9zkeEUYv4TzRToq7x
2tARa9o0f9WXBUjo+7OaIuJGXGIVLRLAK6pLBicURLtqA6LFBK3s06mOCGpRcUg1
mQR5t/rG4sUjbdx4UbgM7cMJTRVqnt5I+T4TCk8gq47P2l9aVTKV23y9UIxda8a+
OvbxUtrcPo4dSqEsrBZaFlJxJtFpetzijBuR8DckygkMczX1DkxPCIdwAQqMW+2W
Mi7hCx+WqBgL2aqPor0sCTIZ/82TV1FPxszQNXE5GqAacbNULo02QjZ11P1DLSCv
hrmq3qREosH0OmlpNfTugKM3tSAmqiJOdjIUIvell+jqkaIaaP4/6cdD8AznFdno
5JgYyi/thRyBh80VarsbKvcIOZGQRT1F5vCJfnj3KwNi/T2+gZjFGsQOxcGnVlQm
zv6KGbxLjUEpCBAHTgbsFtu31WpKpKbP/bvkYml+OEviWx+CaI0mRjbPV+hC8Jfd
8luR50NgvWirsDErYObrqAIohY6usliBax1XVNHEacAsCvuDp4vkhZ200a0WuWow
t/oM1Y+enSY2itMrmyXCnfqENHms5qeG7g93+/wBZoDeOqUJz4mxTm/YfO6xbxpY
vXOG7fXwfOLsyTtnprC+bDAsKiZVfB9mmnrT3oldQTsHXsawzjwdeJ15+dhWk+w8
O8Ek1PyDlPVuPhTz9KjC/M/4anB/tJ3zhh72d1EiBtESQMQjTEBtO0sXqa27Sqsx
eUYJ/jDrWFwTrq2vlb/iR7xFpYmgqMtJkpYd7SeksoClEByKJneUuDx0Z91edMjT
9Pf6+eShpfsld1rgSbpI2Sy3FKGBHIqCCSB1jgrxzZ9COcBh3bzPQRV0Q/3rJyQI
ZBE7+NKH7a0QlQBbBx3NkfKZ0h9lpOOZ2byPTeZ3etyU2qdrmjOnHlH0oX1kYrSx
tqM3OFXfL5aLRXL4mnhSZosfB5xbQwfJmAlYUY8JqRky93uWNHkdKx08PWOPq/9p
+oyLyzgMdDRx2jxGKaUzj/PKvqS6pZ3cJEIdUlLTLI5bwKcvt8bnFmpCps71Ps5h
TYLRqfPRQ2E+3K9A6TxDRr1/Cd19mcRWFnu+x5xYo3JmnDUoubzLQ0qH3miaKOIh
GCzxrTfJdmjr0IeIuiph9jLXMGdURyPnrRiUW10bvgRUhmv6Mm4V2XcPtnUm/O4B
x7M6z3DeKDVMY+oPxi1/OLHWLg4HqHKyNEEKStoj92H/dHotJblLg64MoiAVZqCb
IWTwERxOUwUATj0oAmqX5oFHWzWwRDDQ4jNQqSe3jnZmy940FyfF1dcE5kg4OPOO
kYXAxs8FCgE7I28XZMSxt+S2oc563njV2tnF8s1VNLE7OoDpLQkOXImJV+CD9Vl1
dc+W+bzfrJ22iJITHruirBqDXfaNhLnNFX8DVGPnLoEFVkpbVM/fK5RJkC/h4gne
cdd9tg0NP60oR5dNLnrQ4OqWCVJBFlS3FazhlpXp9a4LJG3asMQp0WRlovHrO3Jo
YRIY42bTlHyTldCOBLsb7BkONm8rS5ONwReOyKwflpAfr/1ktvsUKtSJOzw5B6UB
biVT9VDuoDGAs8CcMTy8Yy6DPp/EFizhJpAXjzyElaby2YzWeP+mXfDGchn9GIHJ
w845Nuxkf5xdzo3Tbn9jgndsa+RBoJqRqkPsS/wfGYmTvz09lstBge2dLWLA0OUr
ZuNTV0FZB3lmd7NHk7pacf4G28mHMrNFHUHem32qVVIOvT/mPtPONVdtoxXrbcu5
8rspSYqKYDkJ6ojUJAaZMmZM5ZE+1EB8j3OVz8dzu/UxuTXyLFeLOS5P6ir8pDWU
jFj9h7Swan0tLakrMgSA082lVdtqbkMeJxufH/DSzhEYgTrFTCi0yorP+PJqd1zJ
dN0X+DpFcPSmYTdrFAaVYplFvVi4WPw+2UQpVObbGA2mn7i4y9fdno/zNUOVDuNh
HNACgMM4sdDOgbrqqZMICoSKctoiHTwx9vcTvsKRQJ1qNg8dHm/MVl10aJHxNqfh
7BI07e7YQDGK8gGtvKKodvKBOYVndNXx+vYml2/9gxEAKPNfu2JkpwZoIfWdHRUv
7fn9JG/WhBsG9qqe9JrCg2bdP+ti52tZC3T4AyHu0XLYS4kB8put2dVINoYHv6mZ
RY0a/ttEQiVNs6hE79vSU6sQ8mwXiJjShh9cnF6A71T9TXf+qtsEPXZaUV1PYfBu
SCBszY1Gl/KRCKvQbyul3HUNcL8MrN2SRPdgHJDzqYoh4DSuZttImOPC4cJCFv6Y
j0hWi6/G/9FG4OaFzwBmAJwwc7itUKVxxVaNlguKmYVq40f+q3jdoNt0SgteLqNH
du1AaUMu8BL3UdYMOjU9hgE7LFilnq1dgA0kSk+LiDijalzoMLtbokH+Af/nOCf2
DlVXKi5g/MCwHRvP/kYSHhAxN1lbTT9u6AL/AqD+j6HHvGWb2CXHqGXtvB+OwfD1
BdLcZJizhApGOuAXyQwHoN0RCR9T8rOJAgRvgcZzHW9YWTRxo3fei1DGbZajPD/I
+DeQbDL70wzCvw1bNWBaATf8EnGCF7sLYL6W03js1sMXJglkmnJxbW5bBMa27m1c
dzoaYZ9Rqv76zCYWFEWu48KEo9uRaVjUZ68k5awvaCJAmlP9kNgrwX5uwwSV8KZ6
tPVwPRuVgPqR7CsHV+mvpvlAioUI1SjMHBQWEOZYkQVFYKp6JMDSreA9NcrTskFt
S85cj6R7U5Kk7jkr8L6LzjGDTdyh2lAHCvLSRnfwZG5+Ee2IQIS5Ncni4jxgiTAC
9RER8GVpFLemHABbm0yVhsf46AmP50cxsa1SYtThxnFY1qad762jIpfEwBaLx2/c
q3qHkkIOeEZA+akcal86guAW3/44yhycNum7TtJXHozLf0Lx6MyjNU4sgjyFuCeE
KM+nbVNxzuQKuUeehluBDUiEGtfZ9liSQzTQ0XximtoekE8Tuay++sziAQzVbo+v
aGskcQbDWKgROjJhdB05zf5XwoZnmbTgM3/rJ8E+pTMac3B0/vvx4kIZ15Tn+aqA
nMXDFt7T0ToVPy/hF1VpxK3X64l1f9Bl6f4llJZgeQnQazpkPuncZWOiMbKVOOFn
LHnT9BnTnJlBKaxkT9KFcAAC/JK10TqCXgHfU6iUmSMuNmvzX6oeXyfigGHFTDIk
K2m2sc2ODU2WF92Yz6BguquerRd3W8ezGKaQ9sJLX403xUZfWTVETFGWQ2r6fIDV
voz6w/heH73CYJ+TsHciXx1N7ks9a6PHRyxKbhcm5vG35pMOebi2sfB02QObWkel
CetWaoYTVsDyvbY5DY0YTvkD9kS1CNwG2gzjjbVawNi9QHZ79olVIZN90hmmOVTg
m1AqAEz/PCSLne1eSl8ScZzctmIx9FF9jcvMrMRIbcaYntPYVaa1aniPv8vYXPOE
+XofWh6w7ZICcH3oB5bcNsGd1eWxCThZPD0Q8lgksYEuttltNftiWFFvL0FOZhYN
3wmkpJzvvFiAR5VwYsWGWOqSB0PaasNzX6pk1dNg2r2HmfUupZvJ+C18SIkxIZUq
jwGCGnC4d2LESTVmkaqH6985CPh7s3KZ8z/1J8iWmSlOqIncl0We++W9Smz4V6ra
9A9o5QJf9eVpaYyizMEk8tDcolP+pQjqkCnH8RC/QvC90QtquIt3kgbBO+EvRIS/
qp66OjEdcoVrgBtiDItjQzTWwJqOESCrs8kazbodhJU2oHwhtfrv0NDaRnEP3Imp
tIweKS6+WnDRgxmWvqofeXindyOhaWzxscmfWO9b1PilT2URhbTPqQETtFu5vp/X
tton5KaUIh5ykCJ+AGGYV8KzdXYABxbPHetwi2V38I8WVqekBJ/pTJP5125E+HFv
VQjMJ277x5YZtnm6AX569pFKZDbRLdJb8YJY6AsY3K0gw7pB5OAe6vmIoriVV2Ml
LTPReQQLQbexoob9kpjGOWHK757BwGHcj8DX1SN0tXtTlDJ3umOs6QX0U2yQiRAr
bsdN0TJ+dM6iihxesaoO+aX78NNFvvDC1G9z9v04aRU6krscO8+X4wigisu0XAgv
tYM8nf4jL7rUEcw3HboOtxXN4TdLPuTn4Z40adfY0EcnvJe/S0Zwwk8QOKObe2Jn
gj+cULl+9r+bvsBPFd4w2nnPnOaqw9kJq8PIMPJYNvYmwQXndYEgrP+m7xt1E18e
LkMS2wskU7NcyW6Lvny/LNjhw8F1ioQdJISIHjhjQOjp4MNWB8vbabzViyzLdY7j
OngI9t2avpqqzuBsu60NiHQuijSIVF3wlrdshxa9rPskWJZFrbVP0l5Irswd4wim
ThQ+as5/a5NtNWq/ksX7viB0cojiqFxCGK6JM6ZZ3+yEL63E9rBRlGNBy4ffBbkS
Y7brRB55xuVPOXPgbx1Wr6I4mYjBWg9X85RIyXmw54QnVnessKbGI6o+Sx4Z5p0H
4j90xDSZM2Xl9aJfgOY7r8ost+BTX8gg0JJV736tYYkMqM3KzysUUqawWfap/Yct
bnAyEW7omUs7Iuo/JwwdCB3vZGj1Zolgt4pj2hVadkanpyyGDSZ8+qVwx+r1wwk/
oq4pZdhujA0KT4RADIvOw/X6GGUHc86cycmugsJ07iD3Q6l1fGn6WA5u8ytCUpNM
097i3d23XJJFgvY8Vai3rWYssqMADI/n+CX60RFdEc0cXDfz5T2TKjOuSF7QzIre
AkAejfutBpM2crx1CZHddHo2W+3TCXE6dJNr0UnkrKSYZ7JOp/faUb3Mep77bWwO
+arpT9JPZRu4GlHoGrNUw/0sl+tZrI+KWmuZxiNbcmWwLJ5anyVLLTnbwzGH3kXR
gj6btld/dys+3xgFlecvBwPG8iloitMdCct3uRvDnAEoYAQNgawvjg0SMqqHvRB2
Du7noT3nqwUHBd8b8klXBP0WZSqFmnMZ5lysYFX1RQV++D4CVXgyHoYPvL/GOZ0s
QylZ256iyrodBxS4LEdeiTkgq0SybZv9YExO/T3raoX2CxhcNvSZWFvYNV+VytYa
MsGcMPZ2tZpWuRYG+ZnpicFd5S8HUBhOkK5V2kbJv5t1t/4lvLq5pLCZzTYO9dsb
ZfOA2PPCIZUibHHoDezTINYy9kCApIVGtlMTyfC9mU2eUq7KlT6BdxIHtddnHuf8
maI2JC3jebzimmEWAaGoycgM/6zGheG0zgqxYNGJgdZ3etoak7oAgYXA1FKXx9/9
+jitEpulKMwaA4C5sFKt4TB5NDQ/3sST7z3xPXBbTlLM8RZZ+tTLdk2lCqUpojA1
n5ylueYn4rgfVmJs6PhfUMEmOtjQTV+U2CjT0lJD9TzCX6hMn9BrsJ1HAKvq0m5D
hRfv/1ztJn1qEpyR6rTvLpdrO9zS4HYWxa/Itzhfj+E70LrpczbKy12xAKTQ+0ni
Ps0eEStDifjka40wtGSlKhk6HeIBDlzGuSxT3T6lIfHa/NtnJaE9XnsLHe80Xf4w
FVmZYsD2qf+G7TZ8Dr8BpNjkO+WbX7zbIL/8fbRxKU5aRF6K2PW75FUu/uRpgYLO
8BN2ad++uj/7W670ebPjPUXTg7lZHQhpwtAfzlMO8FBN9be8OaKNo3m0dtl45MId
h+2XDEzXwYVObzXhF9T6fAgE/20D/Hm8nqGQ/wdzic7Adm58nr+vqtS8k4FVRe1A
nv/h8DgiXm8mrEpuMEJcqMfhZIFTOMO9W4euDjs2CKtCXkaN59deLJmeX1mBDdmb
FPislfreV2llfImxR1JzaRUlFayH5lTZ4+iOtOMmBjLA3Dzguk9u4uidwc5wVA11
bdRDmhrmIfq79zqwg6S0o9SBf6VpF0JKoYFXd1gKLospcdWr2KtGxB63axxHhTU/
T9qD5Z2vWR8DPxT6wfhSwI54mFUFiXgU2Zw17q9k1+brxE1qSKbgbaAfzLOT5+s4
SdbLL/LlyUybdJz6JbyBAszuuvUBgjE5vxOnaj3GoICq+RBFX1+HaYWQvTMxsKwg
yU9oMWUg0rDLzpp3hTV2aNV7MzKHa18eGbGg5JSqC0LzjkzHT+uTF63sxSrlpAjz
//TFo2uNR51ZAdsdIbArsMq8Bb0Om7ydUkqvqRFfbd17TsvZIvsyvxVx3aGdjAzF
/N8fGC/o5tvQVkCUwI3iVacxBw0YYJNj9Z69/MRlY1y6i0IXN9hsHjb9QO2X6ING
ueTMQ0ko5hp+qPw3cTjbKTIkpUlyrzXioDqqXNdnxWjhEu1nxqIJIFx6IzTW6MTf
sLH3nwKTRNoybOFsFrcWNmchyJ0weDEea8fV4xzB+j0JC+PZXUOQTxXpIitoDaEj
7u2zmkEwSj8s3NXL87lachIGteJuUrAnlSsdXVa1aDgbGkDBehqvUnOC+QLqn1UD
rfYSNwu6WBWpOqko2mECB085er4OY+6IlVmM4k48JEAuLs+Nv+d6gOKxgFpwNSu3
FSyr5yUIu9Wdmy1cMGjr6OTxzhPdow8Q6k+3X9/qHhUNZ7CDD/H7Q1OFqLoMdQA2
joIZx28KpSI3ItNbpqOqeEL6AKaDE3wPkCPaNVRCBR/ns2P2pHLnz7GZqWxPZcXZ
h1HZDqHaYJ0/Ks0s9GRpqG2Df/vWCyI0Hj37u6xAkOdivdxHcAiMq9xL0iAGMuQJ
E0RcBYqIGBKSC8kZnzW+zKcgxRig0Cp/mjGjkoJCm/9m6V1ppTmoYHdMdi/obaKv
MRJlshPydOUSclzLC50AP7ZQNOkCTwNDfBIp40AaRYsyl/owuHbbNhdsGdoZINhF
QDYsAMcjVH6ePALWs5FJ5o2V66Ni9P4WxOpDEf8tQYsnK6Yg5FON6nk+xbYYPDXZ
kJk9JE5WjtqxdlpoFOoB6eUvn189zotMkwKygueVONY4R68FZHyvNC1h91O29pZ2
adrcuq8M7eITcIlflZ92OXamAYOYcKJgq8XPeh3JG0Bex3IIjx8NElzP5UD6Cu42
Vu1sy0iOG3M0KwzIzs0f/oVxsZ2fRM2ZtuJnLKwCH29KX97knBhjazgMFJ4aAsE9
LEIQwoTpq8zYxhMPKkumKWTf5BG3KNZoESdfpiAgCoV8W/U6UGxh84GAElvRf2gS
lUTRQL4p7TbCxYRKjt9kUGto6hn2aAQmO7HxpL9w/4I8eVVtTuDPZDBvBF6kKPSg
URF8TZSIZLb4FZT0Uy9Etz2f9UFX3xVg2UjsmwlMuyDhboqpX8KzNPUNyLuItiPz
QVPYZszr8yaaZVx5Tyu1i6YWnTeZ24jZ137/c8t9re7YdKlIWgUQgEDryr8bkJNs
R4lIRD+m6L5Td1TOzKLCS6z6yaKZmQPWbOW2bIaWh51LxR5EA1ic1GJGllqU8u/f
sDlEqsvVyh/3W6XdqZ03gfzR0UD9FcsXPBx2girqo/aYc21O/gjbv6xK9EhLZXGK
+H+E8x2+G9Y57VPscnZyRx0cQA29TRuHT7s1AvHQRjUPkA6XM+/QAkUwEuRxqrbk
/AICQh4Eq4n13gJQYHM4gn2Omq/C1FAkVOaq/SWbECf7Qo/lau15hRBLFNmNL029
z2hfB79hPvx3eBQEU4oJta1OLCVu4aX8owab2cornuOceiQgUX4f5IGgiDFADXkt
uJQLqW4suxjLCHfBHMSoFElFICoQIFjCTFpYAglOxODBNDSWbsnJWzLLnZMLK+eh
draGlhH2tlAKpG7dT7XTFkd0t+jr9yf5+7P7uv+pHLoA5C4HUJXlZnC2S35HpvKJ
FQrEPi6oVJNnT3YucDrm/4nY7KV43sSrui33U0NRbbPdB4YocMRMRcrwQ3b+rn2Y
54pW01hVyP6Cb/5LVPPOkaMH12zhzmhyOuRg8C1TQ4oQRcUbvcp6uS5XR42wjm1w
VWMEGNgHKFngAo7JzmIzaISBauEx4J//cf4Zdwwu4r3IPPzcz++1w9FvsvDydlcg
py4Hyx/rAQ1T8w31MXOUrUTV1ZT8uT2QXOg53+425zZLluJZ/AcFV2ONgAFVJyEj
5bjNAyV7eItS2muTuxg3bfR2LrkSeLNKyHayTft2ZkfmRPMO6tdYyqDoVes0UZC1
5mdPAVq2yrN22CWzyB6wWfN/A+Ly4G7jGg9wg/CozNITnOIi83+GbCivVGaolWVu
1zH8Y1vd3RoI+u5LJVPAcZYq8Vg1uIxeJJsWlMKfGYrnywlEUoRCEeu1RNJNNLVV
Shx45m1dwQIp7RB6BX2NagMVvHVRdkUIT64aCKsAZw/X0kql2SI5twh+oQZeyDyZ
vYqCvkISB1a1+hmo/kFIPIE0bfNDN71U088rVnVWfokk66Ni4z9KV/+XNw8vk2tu
U3G67mqs4iXLdbxxQyq/kD76li2TM7k1Y8t/pxykV3hKTTisehdSWKJQWTKaXn33
BQmjQMBE0LsjT8xFq/v6ybr6vq+zLQzrO8sYsNeTt46TRlNX/D1I5/WgKaqVdY2P
KhWgsaa6m3vCIe0ysE7vdE0HsXICayurNitKSlqXFSc98w/RcdkZt0l541AD1MTg
YgsriUmiUktgC4bgPJBngMMsPlwY4uO65mymM8UA+/J0S1+RoeDiSNfOMX5GPLhG
Sz4XB0d0zK8+bVOWxQI3xJUCpeKSEVE0zLxWLDROFJh1WrhCjr+h1OYt+HDlnf5X
+QrOH51lFq78CPQ3Vy9wDMoGsVQSps4/g8b0DJnC7uiJOKdTYsjd7aXUXlD5LFDT
36n3NXLAOVOxJIx2EwA8ryPJVjW7FiQ8H6xXFHqTz9oKLG5SsraYNH1Pr2DDX1NO
RqpSlbQU+rwDTyT8w/BvSahEjcr5AB9Nzw9ixPEx+HzgLWmvB4lwgc7GX053owBC
yeTXZ7ftRn8tUJXfLi50dXrVZmE4ar/ASFbMEekeS07LCHhdx/BQbrYfzhqt3QAz
a7ZgY0tMrC/Dvlydu3DZokNrBwOu4Zor7Q1ONE1QiA0nVu7ja53ftOkq2wsE9/Ww
zqKdm/VXmHrFByoGc7fJX4YikgXBQNbvT+/FGeSO5o21VXaeKjPwozqA/+cFi8QK
JnxKBn4lBIy5p9U2U/hKEootKLPyKwAPeC+NVIHD3JfHeeECFSwvm5ToJJA9EV2/
/ZHa4kq1F4LqkYltbUbMGBRsBUIXnIYXkLl6T7Ju97gqz6tqHL1GZyZc6FX8s1V4
KFsAXkxH93oiuRkhBXQiVxX+PVyXs1Yh56AoMZkKWhwg0HsVbY7xPSIpIn5M9uK8
Y9al/W00pw7L+Gmuy3wor+UDrpi16mdxzwV3sORN//sWlUchDFuzLBgBCCVDKehw
Aot4o2kOa5yHWIa+7+aMUnRk+UAYd5FOKkpkT/yoHuRrFs9pEP2Gistv37GnvHvN
58sYEIL1wo0/kwZiWN6WloyThGg5luJx3u3iHhJjLwnr2dlkHMkbfnQTmluOZewj
VsnVZnzGDHka/36CArrywrJ7i2NUtPRXRzhm5JCPGeUkO5VjSg4bhIWRv0grAtmr
667RuCT/LXgFADd4syoZrLMV8YFL09/w2jL6uzaNaY9Vgpbr5Nf6hLh23knMvEYj
3zSLaBzH1WwtrQXjUC9SPl6xPdKw5gKAaprRltvfXZJY3jPlv87p5omch+H4j1Kz
CSi97xXP8d7TKvtjaq5V5Mh9m5skj1xhi8hRLTEqDK4mFN3e+iDiJaK6mRcVyQ69
3wkP/qoV9I3amhLV/R26RxEvvpO768p00iwqcrG0kpam1ZT0Hjeid5/12a0/Wfcv
Egf06/8ob513emhM3zdaS6AvmQRYtyQKFSsd/H87YZ08fZOe2ac+66gU7o0uWhG+
INobw+S/wI1AhV5Uxy1ehOhhpKK+qR1KEfzzImgfTygYTPP4lS2NCcJoOr/Ml3v0
Oe6MrkuRzNHhp02o0KPsEN4pg1nHdyj2fn3BJJubs1cdSRV5jBFwYzfyPk1X4Y3m
BTLmKBXa+Ok81jb733PQTwJ9+7soJfFn9SWQddGgU5S4ApZghgbMuO1O1Z4jgq+v
r9Wxg2b34UlnEjhaQqO2zdvL3Em0w1wWEBgtbzwgkYZ2M1mzkds9D5kZcx5BPy+G
OprPrbhiBAiRDEdCLa6enctc5UtgTY9Vclvs8mA94DdGQlsBbwUEjCCEKufhYT2i
TD8X5W+mPxiKYdBgzWmBCQX3CmbTCN2aE9kIxjdlAEbO+N3Jkv28zhuCVBb8zBy1
tcnTjfj57WgQ7yh3bjkUl1iL6y5lmZ7VVGpYZx8yO1XMt3RxNDqzn+Z+UuW+IOhw
2P6NJbd7U9gOVgDT3jAjzZjtIWcx3+sfXJdUg/nzCFooxGsow7lqckFR+F+HGwYo
oHlNJ4zPwfmkYKPm+/mGsQo2/F8UlgAlH0xnN/+CGItn9wZywQSRSSCghUm0MrdM
ADrmKkEe8XIrBGtObxBdfmqZhg9BtacdOLmJjSura3tsaQRdNAK2Do0z4Yx8MYNF
k9ra6h7BbCVtO7HYU4K3BBUBj7AWRCXUofDCX5aYaIq5bBYoZBweLSOIhU+nDRQM
1YJl0vu/N+yBl5ibahqYp1tmDhuYrM4vjZb5cjhWZMeqVc5qwevP4j/bRGd9sSmD
84tu3yMM9OSjN4M7QE6/X7ON4mHcdpsGabqqFriLoZghFwx416J5vBdTtT8UoEh8
kj9iU2ZMiiLuIIUWFZVTOmxUHuhqqHqmZOXkerQO9LVsVr7ZNK9r1yvqdiak91+V
O5GolXp3wR+EOxtzArSToos0gz//VnIS//vKAqqaCCFCKVpUIEghEskW8TtlsEK+
LCr+L/VKL4mu+jF+iYzICvwiMR8i0qUBibV/OVDSO1xuPVUsrRac3aMzMU0g2hYw
NT3ClyX8EQIDrgA8MnaACP6wsgl89Q2r+LsNv+fCJyTRK6eSXP3jQgObWW41Qxq2
7nY1extYOkkxvok8AN+9hhNnIe6iOF/dzX3eRFJs2NJWrmGep6poVnQcOl+5hfwe
hwctopRaptB7ZIG+L8h0RNQTDNJRUaT+1/5b5uPrEYMWQUh3VnXz50hhqNb+ajx7
+qTR8gNWRP+79k5bGrCo6FOXDIFvevboUqPgNfXbD49Rf0Y10WtwLJT6uOJenL8I
rUGBOrKCrxxUpuXTj+PGYc3N/kH36Gc4L/XqrDjf2+iZvpCMtWw3oHjWHbTxuBIj
O0IbIZKZ5oWykUL5soOggbseLfaINngRirswVnP1aIqOtd0K4N0YMBBTN55Zn7yo
uBGsR9Rt/tnu70HKXL+JLq5lA2U5BEYin2q+Jht7sk235/w6GS1D/juZwN2FFf5g
ARBSEearzNCbBrxO9wkJTxP2VQQPSU74v9MruYq3WvHgvm914xcdtuwBvIxUVruu
u40HJIn1TddJ7rbDv79OLZz9aTVuvmaf1BHPOyIBuDvLRP+pr5hVYklD5fwJuKpL
+TLVBuVDLjh7ccjVlsQ9jJeA4+j4R0tUhGOkW1dCbp7oNBhT47OxyOGocBcySOwo
b9kspBrIpztuTFXTXdAY9OqZTFhoQQm8zUOQG1CN7/aRjt8JOC+/Jyl9PPSeBMgE
pxAi0m6ByQiloZxaiQhVJre0yA9DHXn2RAkRWfH30hYf46f2FZ8eIOJ7nHCbkX8T
SGw9I66caM1mxfI5Hk3mHb+YBH69J6UvDeATYd4kJEsTLmWwjhzkcG7G6OchzQMa
aKOfMm3jJ/FagDy4VOZf0aABmyl2o2o8kdshXSPgT/ufqsAhGX1Na5IYMfs9bk6/
TjtJxgkAttZlXQevEb79oEzsBgeb26L3OJG8wYl/HWf3bwl4Bdz1LedvxooZgX4d
u4vtKeNhplW6tsT0CYldbGDXAVFYENiWdI5FRfzy4eJ4iNwdQeAM8TvTgb2Rp0my
DYLbCdD1qg1xDOfX9rynFlwcdDzGGjLTZ2V+CMg/exGQMANbtuk3QO8BwMUpX7Ep
hZSVTuzjneUGP6LmArERpsMRlXU3llO3WMG/a/p5v7Z1gzVq43/V7+/ZFeEx8N4J
pYhobCY+ghVGz7lchZncEaPN3JtCGrjt9SRFWNXs6UR+Qbm9rq9+uRk6NK4HE5pJ
opMcsZHOn3oZ/EBJltEGpkBgEOw0jbrK8aQPDflJ47ZJmNS95OYEQNZ98z7HhvYs
nCXrdu0RMyenjjjBxAxwOpeVtNDBktdsnRduPU+mOubTS2GjLZ1qzchE57BQK6sw
jOrhLp17xc2sJ6oEcIM3qK4jAzUVtYqFmHxafZ/AAD043T9aWGUqGCbkvVJ3C0+C
iynRMflIZZERVGLdU49of//br7113bDSeaFD9Ei0C7IUzxifzgCk231mGmBRSaWF
LcKu6bvSBUjAAAffQcFYSTPyoE1HKQ6VUXz0qHdxXXoUcKWaEDIOjhY8nVn5GM3l
0/hUz6oTPQiPre2Tf/oLKqerCY0stLUtV32rQu97YlSsnflKxgOuq55CcGm4jdn+
a76xRSntMApOZ93GYnnoHitL2ejfdZUFQumCZAPG9oYiZR3EYM/O6jcBz81nZDCt
6kG2YmVf6Oc0Tst1y/NtRHk6j9fUCtT5qn8rxMCc35GkOzoNGgT2ROdFuZpQMKEY
zKwRuAi5PIbC7sx74HzaimTQM3wwwQZQMI8+67lBUVimjXzCxFNiFtXT5WmfjJsA
yOgq067MnpTtgBqwGpuVncgtaprgzIlg96gL+6PaTZzR2LZ7IH5fP7aTOg+RpbUP
/1Ef7IUK3pJs2W1kAqKyXuv2PmeW8bh0F3ETkkkMwPjIrg/OF054mOguFz086r1z
4QLuapEcDxjxUBRAgVoM0M0ryPKjwNJLNZoDvj2wvj45x3k8BGszBKHE5Hdww96S
VCCicFFV0xQn3TYpqCnffyp0EP5FO32Sf8chG+GB81l64oJvL1aqL7wMMjZdk3zN
cRs2vw31MdLY4bThBu2vU94l179DwtrPahdM/kW3vnPQ+LZlzvGxbrIwIBd0e0iu
/3m+a5lvswTJvnp480Ksw6aED1FMnbhkzqHZUyTdrRFjEbCvhB+TwEnN7L1ZTFgE
0KBy1uYLcQ2ekjy727Ym0niCZ0hyYCRa/eKggnet23R91DDTwMIGdtjuHb7bkggP
m9o933NjXoIqb4WnlfIRINKirFUAIVYN84fUoQ51ojoir9CnL+BxCZ7HIHqSNepq
UDlVVhsPfxkVstLlJibAdIBnNvxs6WBV8CsAnpuxCMxpbH7vTRAXq8OrV+vaC0Lx
OhFT7hbHdG+3X2s7nE/BoV0rhzehulRJ3wE8rlbGTZ91jV+tAAKjjBIYUOL4bOOI
EwKVu5Y8MQV06z/vCyGDxnsXAp3DPqPCP6ojeRSVqQb28L0WXwSJB19142JLhygO
8apiqNNO8gWw+CqsBm2pekRAulKc0O1IoA5QZ2FgIH0TKyqqOFZEF7Y2U4cvvL/B
q+m7ANlFEONNglYYRMdTeL2dy/3YCkoh/7E3q2G5Si3/6e77ZpiV+MRqAeOa7NDv
7E4gYAmrRuU+K+bunrFdpn92gzMh5lgWLwr6jkpdEnz4rUojp+SyD9k+6UxJJRK3
hftiIbxvGsyXVCVXQogh4juEpqrH/DysAvct8CIHPtF96Z6tJR1bAFcjtGZTqVuF
PRcwdxO76P4xI+t4+xG7Ob9G8Air+hjr90yiNFcKptMGDbjq3MoUxTrMkhe7nPj+
QqaVbZ8h/Rlp6hHbXVSXhvHn/XGvFsr6NE+rIMRt+EOo1Yjw3v6ZBKKeEiMba+yJ
Msj+DB40BABvozkBrA7UMh5jk8bF2If9gFCdV6m2JMMWzkILJf5xh5tvYppZBkPt
Qmlhbl2+y1AYPxawm00er5M2Uo/PlxKafRFlGlkmnUPkele0gu5l/SUaTewT6+C2
WrF8obgIE9Jsu6k6fuMtdecYB8OowWHJE1QOvlK7UV5C1NgjeFVYERNqmAmNn2Up
IBCXlS42LwjW6W3Mi6qVfyo2cLKIN5jJUrRZ3jj2qLic/UqLOOuWa82nBJLns3li
Y0+dr3bMP0RcVUTO4bLdV6zFzxBxabeXQztfe0o2pR8Ws0xw0h+bUDlT/6MhS8uV
KCZpy4jhoXSVzuz8aEmmTGeM2CmhIv2wz1CfMPIm+hHnXYPy0dxK2Md1FUng5L4G
vuTVXSCpodahlLXn4nOh9ozh3xnhAIzY9uPXHpkCUm8luDMyP9EYbdGmDYhLvLZK
qs8CJ62swa3Ey1Zjw4vmvvmKJyn6qW2GFnytfbzTrBoWfNn3UVfbwX9LRMMo2AyU
xIkRrGoIXcRtJ8yJwNErG3bEPO5Qa7Wyk61XRAWOdzcqktxLZzcr5I5ch0wigaMd
7z/hPuvu/phJ3qhWffQrvQBWj1PQBUWYuuRFYx8MS6mCeWzP8EoJx803HKhIDThH
CfvM7YGEycq5gE+/SFNG+LdOQ1BwlTMDazlZ3Zy+laIh6oVYv4Qip/LQomMK8dco
nHz/YPWc1mjWCy73maA+cvszOb8/CA/OpXuzVHj+b+KbknTc+b3zvuJxcihmgdDr
+y0cGcGZEYM3DrX8aA8jlqO3rJL4QJeikCwte1ojr/iPWMdnlWwQSWp4oFyVVJ5r
P2GrS07/mqpZovElcHUDAPt1M0toSMIkaBCvNBelW/Kdlm8KBLtBDMgF7LUfkQnP
1bDNTQnO+68wNePHXi2MJ2tReJO2lyzuOTD4C2sCVhYKi3d32fVj2YXy51UD+MG9
slWpKpzOG2/r9q4a3jGXUEAoCqVDU6sAxetkDerF6yx8KP+45Zx1vMrDHVf12vjP
LqIiinG9U6Xhr+P7xwVq9gg2fAtZXPINzgM1OJP30QvA9DDSmki1IJ6Bib+Sm2Ht
muCAC/VJM3hO0nB2fPqPks7yXxLiMpegKy/OFoKw7R23+k04Pd8T+F+IzZI/l4mC
f6Acpp+5y/R6ws5AuQu6SfIyjva1jfaiYmll36iKjh+FQx0nrW8621tyAG+Uw/MY
o/EFeIRtNzX+cr/n7fcQ5p1PbBzrTQIQJBMmdA5cEHxTB2mbxO8RHC7XpCYEqNsS
EpcIbg8hfY/426JFTR+tm3Ncb2XKphK7AExUydYfPA07xPEgQsXyGRuv0XPDEWq2
TYPq/6J/D+bctPqZOfikUTv0djoTT8mpjs5zT9ICf+dJ1bwNJQ3hyoNw4JxJnMG2
rQWmCkRoW86lYvQlDsC6EjC1sZk7dE4BWOXAB4DPiJP/bkD0vg6VIjxW/MGm39aO
RnecJUabVYFPrVQSDONmcO+UtZDwfZBg++OCFcB9BJZxsm2xDyCcvuzfRVN0+Dxn
qWN7QnmOpHa0IBxQlUqtjy4uDzKk1FJXUcDgoi3GbKNv3L6GWXW8KJ/ecM7ckFuj
J4F7Vxw6lFhsI1SL2596VyCrH+vYn0GHcGDNPhPBKiBij0ORso7D5b+7wY2b0Okj
VZ2Swbm9p0N27teqLOcYUbaO3380KcINBpxnDFAEpIizFX7np7Rel52F2luSJl6e
JLLlzFglekn+Z8qaIJ7u9k1RKmOEk7t1xOPgKgxXgARWH7QpbKUiUSjabmeo85Jj
jxcbKauRqY6oKIZ0knfKmIWKwMQrLViBfxG770Te2z7ZBaM81NH0WMfrX5n/+nDT
IlshNM2IwCk8/qlgzbnrcYR25VG/5UaG8PnVyHtY0f71eadAPk+gO8U0GVt5/yuz
/7XtTgEoGyc5EwQ4B+mMD+9jA8nCYYl7oxPsnt458kr6HIh/dnpgRVnolpU+UFwB
eOjfS5dQKHM4LrnIPf3DdQm+92KPi+DC5ycZ2kdJ5DNJzV8GI8JPQdAvStVsMvcR
KBfe+V5rrsN44QXAC6xeNyJQnXY/5IHm8Fa79ueiNiHP1z0Ac1f3gK8UmPN6JRrh
f7eluJkDCF7tke3z9xmxFzVR9DuSVNHNLIEyr237UADDv93sJp//RG6iD1IJBf0I
/ZZyuhhm+T8YpeJ5LxLk+aEPtvAzeO2V0qzFqOr7DSm/vJwGkBFZzGp/lcm8CEgZ
qTyqt9RDQTHYRNclvB1QPFfDWqDrlW+yu5Eolfdb6TL5rRzyAMpwKr9qqtAr4NtW
JEi0NyIpnUlO5GjC+psbQunLOJ8zrPTv56KBhQhFxbqP78kFjQon8xoycxf71jMQ
HY6GKbIguQ8vm1tLJFTxqo7LaECqMUIjZfaZeh/J4xBcE9IPXjUy7iQpzzRyUvts
Cor0oOhUS1uRCSN9kxr+qhZKHKdKHX1ZMunkBzxQHUCoKXVnMZyzrwxUrLzayg5/
Z+nv8OIOIpWLaoNF3n9U7tmnFHxUn2RzzYmgcRwJ+Fqi9hXNucvDh58vbktwQGvN
ripZELk1P2ILTWWzKZY4b5ShUszOvS8hB/3Yu4CKqZHFx4UW8b+44+wxHRdaHcZi
vsbLM/vu6EDtxEAMCjP10Igj1WVSZbTQAqKrG3LkEDi1mloHZkNkXqW+uI6FwqrO
gCdrByhvpzFE/Or6totm4XEM6jhYDsoxLiaQZ9oR9KDnwg0nnWQ+JCsdFmKZ7jcF
B3+3uQCUaffcR+EQVM/gQ9y8tGLutH2YErd4wmnbd8hBoCMgwyzXqbkPCH/+ZftY
MKE4qOk98b2VcnWx7mKEQXQ5pMS0nto9qY2BgbqgLvSLbYeFa/BhmMWJff2vOX0w
Sm6fqUWVB13T2yNGSIq7S1ojy8a4lF3TUJHEwhHtrxaEpw1/6BaeuyoJR7+e/Zh4
UdSZBwLmUTNq53HfnGhFf5ameaI9ZF/kLTLQHW2rE1aUbWS/By3RfGeOaSsxb0TS
cbtOYaDqQSK2P+0e//Bvy4dW34yehsbyhAMgZgnKYddSrPzMQ8UHz2ZCEC/CzwPP
ZlAglOUi7l6xmdNdDX+p+rCX19wKEQDM8/z3oaDpn/9yRsecjnAqePjnPVzclWp7
G1P+7qY+3emTLzsgBEvE+mA/FVTwC2THTKvncmYMCOonqdLTV4uWRZWxFEZEfozA
XER4JNKJ8k8pa1Td+ckcxW97nkYkMZlL9MoTAvxzq9RlCpe+mrdR0Q2ieJlBa+tN
7jpBH93a+YEDjb1xpy4PUGu8+IFTLZA+sOMR9pQkC+Cc9bsOh+KdETu/+lX/VApC
UFpkFKaQ1sv31TOW8Qh0h2lhneXnkAoFeXCh39b/QSKQ3RKnD2QP5SbiV0NHfzZ6
Mv5ARl/k3jsTbN9qsWKWj+5/XdQNyN/DXnSs7sDmhKgjzFhPCG9V4pHPAqTnUkKd
DwRpp/Fa2+en15+BAL6ufz5c7bq0AWtpf6u/0AT97JDrzFtfUkXb6kLewsYdauqF
EXlddG7urSUVzs9g5sTHcBONaZ6kQDBKbxJXkXqJ9h77bXcKzJzMZ/soxoAXjVtW
UHKpJTs2qZKN2bl4MsymUeAYHYtw6MU20h0DwzI3Xno7zrIvNZZNrtzvDCVs8G73
jPyS0iLfuaHDPw0xKF2tBRUtjgqn9YWLmCyhrDT/WS8Ir5+cTmvKlkuuSrolkU76
2jwcwerHTeZ1DHKBILRigUZM3P4hGLGqJIR7Mfw+HHkjX9oKLHlfjMCN8LMNbT5d
ImcDV8YJifZzYsZnFidqavgnlO0dXaBBrKUMzgsnlqjTJjBB6YnPJoT+7GAp+iEK
eqOI6pzjuzxC1ATBN9VPbSUJHppHfdmYOJwz0CEP4H6p2Ut3g/9J7jo+bSBUUE7p
5MdvD4U4/mxn66bIacyHX0TzEPOMamg/UPOquMRhAEaWton+UoFSGtEhKk7Lm445
ZB9Qb7/ULLc1T1ZNj7s1hjCTnqyogBTznKnVxqZlKQcBHz6x9lYh+yw7UmS4qbpG
ZJbWuPKbCC9j86nYhjHjI0Qrcz3HSik9eBuf9LXFfcIH2z+JMjBnVqAyVhefwfkO
d/FHEB/JoXHJ/Z1PRshFBEGT/l9BjeElHHtwiJ3tTjm2uL8xmlxILq+OzEoqwX96
UKYF/VebsdxgNo1TmEoZpTPUCLksr5ICZX3eAndH808Vffeqd6N81HoExSxTads+
qFifYqBYsMyEQAh+5ozK33zn8qDvWJwAska6Gy6BaPDsv7BVtgww2q83526zGmKz
YvI4R/1e/NqE6wkNJnne5yswXbVqPYJhLzk5ADikt+RtlnCWU9Fj0xia/QQ5cJui
xnbb8s0/LIpg0CRnDMyx8ALQ1Ruq20+DfTo6REiYkDVi4cXA4Cqs6xMmedDl/MSa
xP+6T9iEoR2bAg7Ew0T2p9Vq9wGIlGCfTQOEQ4zZTs6wDE7U8D05nd7dwh/MIzjH
O3JXzzki/PuUxfX6UnWFbk37Q4eYeM8H6rJFOOUNwufth2pv+b+uO0gnm1wyNpcz
6Wm/DKs5vNKYLJ/wLWRyXGyw9J66f08TQOlZBRV240tniloGHD96kF/fSoB5drxy
1qYews+0Puei3PFUgBMBAIk07y+Q6Nch2vQ6J5liKLr8na2Q5MFkJsZrHTAkGXcc
Gztk9/qE6vw4QGvIBUkPBViGya57pEVh1o3xGUVWaltU1BV3/HRfSzWTzmz9TQse
G0ea23NI7Le6uhOKuOKXk+881PGMnDeidNGr5IODt9tGWp7lNqqqPkWnsCEQoaXz
KO5YyMLVN3RR+hwJSX4wErAC+GALCYMR39GkVWKPr8XSDPsGS/9hBdoEpArnNkVK
S3LA03E0PSQ/KCP/hbWthxQ5CR+ratVFUON19TL5huBuPTyRUZKUz6c2t+To1xrK
bwp3oERDmvWGUEPBwJayidS8SGVMK5SnagFIgt3q+a3ukKXErVbAeyHkz53CYfse
+RHJdPQ3S4p+3VgAXjuwSLiFgKzK364gtDnSruSEhVbDnxuk2xOxYWLURk69LVHT
9aJRGOhnOu0PAZ335uASljQLeXyVn943QyrAFXc9w1Cnoy4xVIvuWrPS5yY70BGJ
+WK0DOyrqVmP98J5QrXHaCAHCNDDEhT/FRmY6QNAIocn8JIwleQZdRnENaJlocsm
+TdHL3QgIh90d9Dz3Q0fvAuVXqlq9sI3KH/MqlFAySej4XlCQM8bnHzZ9lt37GeD
JUQmdksPxdjzZPrzc7hcEmmJfaW55uXrBLnDbfl0zuYcwq2/PilcZ58SbSallVlz
YoEBESyWj/sTAQehar4Am1M1P92GUuNFn6WEn/ulY0pnOZFZ1H+aJoxV0IntxV4Q
SO99ldjuKkmruRfjP+4gwe2TYEpP257BiR9OEz6ZdrPCoY4q6b7WgVkXsFUj7hwJ
OTTIdpyna/On1aEi5C8okk6lJ+14qPUgJKrnq0EEgUBZDppSfk7/7Xy0bD4HdCTf
Zd7rMGz7mSJUbf28yctsibmjKU1Zkn2OgGgv1DCUWwlZiNq/30WjIGY79ROsOTOK
VVEesuCxvmzgDCgjeopcnAB9SlflT78oP515Tn+7RsJ8zDkUQDKgiNLfT9p7kOKX
uQVSvJ+mu5vvc6s5DJoktai7JqxO0mNhTmjz3KlWrvokQUNY0aoLVZzhvuc0Bt89
6+APteW/W32Jn2EwOgn9jLydyFKXpKtDhCLplPsmMEFZ4vJptgzqxrYpyaSCMzrz
uBAvw+0muI6YyaqLnEGWdZZ8oqbhkun6eEpozIqMi5v70jxZNk41uXFW/Gfv1PDJ
TPx798w3f8U93i3nvC/LzPlybXpUw/BK/+ATI8wmjvfXpTFWjsCRukCR0TW3ZCXp
X3t/OIX6J5Gb2nOL+DJCHpot/eBARmdQ3WfCY5i8IDf+Wy/+rIoO35tJhm+XxXGK
BmfiMVL79qO0pdD68S85THR+zWey16ueuRhWrELimlXMSK6YLmVRISQaQj66hV/y
+9HSu8ARyjM6XEyJMtiHkyRlAPj/MecogVAGv3EGGAnIGor6legklVWKw7QNxWnQ
a1zOH6nvLcKZ3iUWkiBTaXabioDE3c32OdxrbJ2a3K7MshYfoe/r06LayJcvwygg
A9uyBI87B6EaagUKAq8JG6cJXJZISinzBuOKij05qMzT/R3ioHWVCdhJ3Ts5CiFt
NE0niUY+UXR5+pzIiojwGKZi3aI9MU1Tp9aj9zLZSB4b7N1XuTVyE/c5HsCe+J6d
nSxTdfSKnyCunpBeS+nUkmqZFvz/WIBcEhJFKGTW/zcYJxVwL58oLtLqvppElAN8
sgsrMdlYHG5PIyzHWSTzMvqkxfs1aejdODFtaYyTzgF4lyeKoZQPOfwTijOvVSon
DqRUoM5mxuN8RCicmkeAO8zxowWjMD7+ScpBCuYcBqJWfNICvIc8B1SbNvEaDwxr
sGB4ExNzXHL9Wx2SPRKPhFBPTiNonQ14i5MaKpVnWW4t4AfIhA1099BgeNTTS9EG
il7l1VKfuCcy/TiShVmGrpE6TEXjCL20QdiyO+Wiler4iwGCicJYMPS1IeymrzaY
O6gj/INvTVLjU8ATb9fmYzjI/GV4gSmuRIcQvEpCy9ICCo7Q/izXPCDehbAxAHJ5
qIuSn77sJaqCEWthrO9kz1WIgH7G4pAHxyWi1yXrMianAaB8nTbCFImC1IY7IGA9
Jdles43yTFZ5ZRMChndImx8AIeA3F+lBkYOeeem5hvlSrTSsPPG8ZXgK/5SRxRT8
HuD6UfNOis9oXB3eoJzxJ8TnuZQO43ZkN2K4IIjXD7DKwwDPtBJU8Bh0+Q3BX7pv
mtAhv//Q5SqUbSYfGFNKnFMcRL753fuARRy50zLFrR1pKU0AsFkIIOh4G0TLnDDq
jNNyy+Kg/4JVyFI+W9FFFtfo84GA0Q+nKzTHFphQ8UjQS8kxJ7vKG/qpMqYw8hwV
kp5ig8HqvwDbGhq/6jZy2HhcyTdhVog2++GmcOhRxtmj1rc+hb+7QuLdUjc1QOiH
YzGEy3TFpguU+R5eY0mFzCl6hxDhHEfEFp59edxbBteKa+1sEbaE9B3d7TFJWnii
iKhEgTRCooY0LsYyplN4xhtNgYcVMpl4yMSa3qUzp1vnSDJo4kAv5QI6Dn2FcZZS
lT660ELhISnkbZUWVhDTF44m2Z/6vJ9YMyXOXiH/SlsXDaLl5Xpfe7P3ODGQzhj8
uXC1jIwjhh8Qmiq4zlNmzEn40bCqbHOhOy+H1em4iorDZjUK5ICOP9JctD7IAslZ
RrZ1zDfz2N/gkAAN7ujGEOikHsdjgDwk4ZcSAn7jdpFLrZH2POlmJzC4V5dtRZZT
3q2b29/INBgd+0yKjvb4AjuXhtR4NQ0NjEDnJ2sx3pkMnXEJY6P73vz+bXdeldiu
237BZQTuwTwhxswcZspO7tdjKjZLojoyAlzjwg8WwJKQuhe6qDfwVAs6RsWGDLnh
TEDimzftI50CDYWSiyD8uoAUqDC/kZJHwe0RYn/bg8osd5Lm+FQF9r469U7ZEDqM
+ZfDDGQlpQjIlJZhfclAHUYIOh0ZXHcvtkF4J9uJYNHwhTHwfOB9q5ucWpv35TEW
causUvKZgXgj9Ssm2LVjjr8/0S1XLCEmfYPBnWd+SxeXxJiWdzRgWAWZDAKWPAUq
GzlhlAUrUYCaVpw8q1+93EDq5ZBcistNi/slv8r/2nGiM7rrJ2obLRci33KOvvUU
zUiCq+DGx0S2af9H0TCmoPcsIEoQocc+c/IqHCGyTFTFDNNKrV6nYItXR291r1xP
F6NlL1Bi2mjmr+FKU2+bMqk/L1VmzsCsg1aTjlulzlMZft03p9bnS14HZdwsMdzD
lz1w7Tgs/pqWZlzSmxPkBPRGDxGjP5GpiFWKa/q+YUw8BlOES1qAKGjljvnEz5zn
uKYGICn6MYKEXVjMktdIANrqTSQWAMnJ/1U65EN+Lx3WDblyD8+b3PKOALweQsWJ
Z8ABx7iuF5qAJq53D5QISk0k3h3Ta2NYbP8GQ2Dw6S8PZms4KNtohQoUQ5XuFYTt
VUcrnQkWIe/Cr5f5RCaSHsRvYAGAfITDs1wysk7VptEalclIO8yOC8JER09yF0tW
QBgThWsSorcuGHhnqkS1km0ssMvv5L1Rw29SlOrPp88DmJ/brnoZdx9X+CIusypX
EENARdP3PWaarPFqazNhCSojKZj7jgy3pq0oVzoc9AhfbL7XsW5YSJ2dg7zmJfzE
kpscZOLRM4uYX3qNMEqmb3YnfF/UYWizp3C4Z3HcfHd2kh10jHsJH9v6qZS7Wn3J
sSe7YgXx2w9JwLtmb/Vb8onkeohvbTT1zrGxts90MmNRoDM1QepiU4I5ZYBY5DNz
JZ8xHQHgtj5L5rGi6Ae++ntylzzvxKUyprHtNdRQQd1iavNvWWEg3JSsldIse/yC
fauiRY/ltDA8XEGZ2Nz35cbLLeOQ7rBT47FnoUr8Ib6TK5kKX/oHY1rzqew7qmXA
1CF6Kt4OfotyFAzIuwGmrPoN/IeTSzRIVKgvqUxvJIsZF5xgmcUGknoBXQ/4De4g
KilnQGfJXBr4FCDL1qOvChWSKrh2oHln5mhpVmjSBinR8SDCynGfbFuh+ssN1DWh
gDleglCsf0TgkFDRfwwPMqM85wRJeZCheFmIQJZthbIgstBwZ46z26RrfwFfQhlj
YH18Bso6VJTRy4Td/pVyyBuE/dAZvIMMXOg5b1JDZXocxdTzXvVEybPOp6d3udBh
eGq/mRKovg0vwv5QTaRg9mwnwze8SYHSF4BI6Bj6T00M5pCBpSbtacdKaxpmzcIC
kxGUptZXxcjjPzsGQuDSXSu2Za5scRQDVdxjQn7ikFSGKQd00VqhLWrBtkst07En
fMBWXNhAmESx0ylo7raGR/XS1DfXfjxLcmBEdfTMQFg7hhaZ0GISqGy+dM6GG7yA
4BECc4qJFGds2ujl5ffoNf6iFZKaF9qZId4cME2mdp7w7FIRIOzYaQeIzpfXiwH0
Jyfo3Pvuef3sDdDbxWhOnG0dNTLHP+fry/51IZt8nfdXHlpnu+hPOAWEw8yZrB1T
09D0OJInu0i3fz3uDLHUzZ3epJweHjI6NkP0JzVHOdPgWpJ7hi5WgjbvWOAAr/QR
j7MGnCQZDAbU7SY77qgGSOeC20NUdfYaTXTbPkxBSIR0XN1yKAvb1ZNx5EZkRcgo
LLDERodPaizcUNJcRp8T9vDeYuRwcPC0404DrF5PfgT/DQGmUPJ24lENXJ/H0cJo
lA6dDDzEoh6Djd2xe95w/QGn28ZYuWIUQiy6QPF+cALIZ5hy/xzO9zwMiKSgrm/a
6IO1B8vaDALQ42dDfKDoHyZ04N97lj62E1xOqTrCuAFvZqzey6g6gRCv8j/O+cON
a0NjMi5VuAYO5Ok7HEdJkTK8MNElWLt5XIx8+E9FaDXBOGV7P4xipTpBXbCzSAwR
G/ZYcakXL6evYyjdfru8Z+vIOIZ/oxKWS6GoFzhG+U7utxkknK0U0MeWYyKAhfjA
1TZHlJ+d7M0aHreAkB5++wAGm47IhAMKJRbCkVIiIFTpqIaVoa9Qi2szzsyoeg9s
Ip+6JO7+J84+wSdnMj3oKwRULK98taL9P7a7M0DLOi4Xc1udn8An/hEh0mjGXQyL
BXv1XwwLkpQ5amPUPAYbzs4CxzJ8wzukWRiWHwKVEu/bK9gPAUUS8y2BqnP+KaS0
tfxIjO0t+6kYgL2zVe12pTfAbCR7vku7yj1CU7t5SBtXha1DmrignwhjAW1dnVGM
Fp4ZP2ieSgdy6e3giVMlWeQiEGjfkTPXkVqqcUPFFE8GyC9yDwUz2vmaOVh7FsaZ
PBzA1w+foTQM0HepQvmwwr3f/9rxcvw8Q0XoAwmX0+3cRqVdFvj/NBWpbbaTF7DO
bpVXUxYJVcfcHOoAuRuVNIg7oBW9MBgbiNjc+P9gBc0e+UuWYFFvi2BEhOOcnN8Z
VoS/VSKdhPVOZxgurDkLx76pIXilyjtTB9Pho8Zpq4G6dOHPN0H/ZWjEK36Dln1K
Vnkm5YhJYaI6aM6pNVo6L9JbEKHauzNRYeyQ5xo1sD77jaYyzY25hzugeYUyJTaf
/0iD+H7o5V6rmxkvq3BMAhro1C4IqbZrWv6OrNDjd52W9nasXvk4y4YxDd7neUpI
NifjmmMOx0ublDI3erigkiTfBgA534vqB35gML8gUvgoPrMJgInw7dBarayvDzSG
G/mxwqIESjDW2r6panAX7r/fib8aJFqfT+Du69TC/x+PwvVaYLn5EBdbttVrvaFb
XyJJp/CfKApDeFZHWU24wwuKF+fEjE480DOc6sICrc5JWnI9QDSk+1iJ7wdi4wos
0OEHa38vDhJgQfZRJ7TXcXoemKxxXl42YKftWQWOh/w2oheBp5VKIFlO/ruqXZ7E
M3m/hscsOZaCAum80ecmFuOKkeAZTMR94sPSJnHHNpOkbzdYuDiInWi1IU+bkwds
J6wPIHEC6eoDV7hRNO5+Z8Sa6Nmz+X7gJo1OKPC5FiDfdY/ws3inPmEsdPuQsDWY
ay0Dier6l0nvZqZoFFCVT9YansbFBEiaUuzy/8FZ3OQLfzHgZb+7Op9OVLBRfQqn
sMh6oG+BMAnP2nuokrOHjZ7O37cLd523g665VB8J1mBUyu02JTBxqQmBkrJSZURy
SYCeAKLLtEU/j1kKLjrEj/97PxrB8+KtBOfnVN+qV+dK6QyNjEnlMJeCacgMuE+t
seKNfJOClK1chjKAdxbQXsp2ggSN4fIVbMzY2cBELrmvQcz5JjHoLU9rw2ZzmR5R
bgWOtCNGh8QosszoNaenggCnbDtsZ67b/J2vdqWsbiZNpLsc6w9oG71I4ze2ziHK
TAxEOW4i7LCxB0uxPXmbKLaFNIHYSml+9XGZxquVSBR94TTfMUshCV1hDLE4sp/x
b/Im4vyub4aD1wI3OxMXbY9iOFT6m7jLRiUZtWnooVsJzuVFeCBdLjz9xzL9Ka2p
70s+PSsyogBdS8Yz1zYO2yTPd9WZN53n6sw+WcPpWvPTcXzJfxALjzQaXm6TvL+P
qzy3HSeEVlAUMxZRsuOlf+px3DoRXjNsVif1uR7rSbDDuPz9/+QUV83VLGjisSEu
vJRmsUxeXFy1f3DRsKeDLF+UOe4BLCbzgKL5RiJhJ7Bf7I0FT6TNPwtBmG+/dqmQ
wVUtHW1oaXtTjBg7RsbS0iBtq4jm5shOo5qJfvvo1b9LRPLWsKLibKnoqC9CNiMx
RH6SR9ftn0rTAL1I0Ni6FQkhLvOhhbYsfrusWhCIwig1BLycJkUICY0puwHhdufo
3d84z8ThSwkhXT79YNHRFiasNnqYQNiQmRUuLCeRHyf6OELP4/mUibilZa6hTR5i
xK3M8wN6C++1PLCAR3gAfL5f+Ad8sAvdpPHTkABvIsFND2fXHtTp/0lCZQU75XLK
RMy8XZX9STYWTapeyP+fVDZsiXQSdRx/G2J4J8xWdbhgC3KEA7PrrfSLt0SYYVyG
XeaH1/PeTbgye6r/e6hZJICzHPVE7fkQijI9iUHJiyW/Yvxy2FWNKNZU08/VXV0W
O6EGQF1Z2zTqm0XaAfBKqZ84anNCDuptXmD+RHf6X8i2A0EhhgkyxHKPB5/90cnd
SlkC9HD3g8huJQFH1Bmswezmaz+JZCSaf8mTihVdiVg+qp1iyU9Pki/wUuMk6js5
wXOqrq5ZwyCBRkyaexiLqDATlTxTfcPddmTb4CoFZnxD4Yl2zro7s0vFDVgGYaDR
HI2y0ouugbWRWQhhhx1swGJSN07TlA9lAqo7dWeRdEduJiSddymjphyRYwQ8YevJ
FmOe/VQx9tHndzDLfN1mNraVt//AFceJ0e29EnQymLll0uITX83fx0IxL4cXcI++
bS2PWel5IiJO9wrRS0sYURNomUAYKzdwUbLpFV711bt32AwZTmMYJsVMJQ109SAv
TWWBVWEHi3yMIyV2TcNLCqqdYupL9TLt/axCsaNEtt3tIxXGw+0wc+QyJ/bjmaIl
oQsEgqbZW0Qb/cr6znyuhBOIdD9k84bVUk/YTjvIL8FXVyj0q4IfzMJyRdPwpQg9
c6WDr1G+rcvNaCCI6kFjeQyBdgdWccdoNlYXDWNlCJ8x1jQy4NBtFpfdySXqFs5v
KDOz7872P9zTqwedAiva03iyFUCqs6V1PJui9iJKlkClPIdEvXTWcDvXvoQYm5xC
xtvCAXEv3G1zQ7zwjDZKjvSpj0W07vneMKnwJUUw70xHi3mvZoB7l5LEa3yMlXwl
Nm1G9MdpiB2VQ1N6kBHfLx8WyeKtnC57+1SUXvqemD1vmtkNU19x/jSgfql2iPlA
ndkWEjAazhOxobNl85UlGJaAq0aof2PLrmKYRl70vPQx0/TG6TUrud//ZXun+gvO
4PUmSEIIB4eRObZKsU0e1SSkYON43d8ADV7b5OuIHfHJkLwqfeAQoa8BOEp10tBS
RNg2d5nvW/YgC1oL1/bhylFRxwu1wY1n334FiQglMuExNx4uDS4G6todVkrMGaLm
WiFlpXr2s9/ts7R9uax7jTKG9Eh/ztkvLuumyhesJxYU9VUXS1Sb4SeoRawGramu
UF8zaOsfSxmlwnla/ZN4br65yP9KUbwDBX5sdVtZQ3P+zltmumunFA0CV+rXLgos
cjvTKYQaSWf2W9RNB5O4YljB9OIZNtmM7iMy9drxb1ILzXGECGrRj7LRdSo+Jjki
ofpAf7TYrbaVW/IhsLMZkdPTCUdizaP50/u8fwFYlBv6VW9STH+WqFQgtl5NCgiy
C8osHx/V3ils/O18cC5pMA==
//pragma protect end_data_block
//pragma protect digest_block
Yxt/vHwWc8w6zlb8CCyiu0n6nqU=
//pragma protect end_digest_block
//pragma protect end_protected
