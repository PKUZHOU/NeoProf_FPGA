// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
KTTZXfSIv1Dwjjz3hMbwBJKcxrt2euAUWEa6HJ439D5OgQS4CS1gs7gc7ct6kA/V
710Y7jVqglySxNTfh0E6eSyqsddKbGbQ5FFW5Fs0aBG0ECDMvp96D03cTtBpitTw
7eMQqPfzvKMH6UINjVocVWhVzHNIRdcdjDGAb75txKY=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 34800 )
`pragma protect data_block
GL0fEinr0DCFuFLgpWb72Gykto3A4tDcp91m00BEws5QUaRSpeGBy5u8QYXsK5C+
dwjJQkyrcbxBghhP5G9kizYNA55AECnEWlK1DlDb2bocf1299bIvgnuN9uhmKa4R
n5RKmRoXH6hlrH1c2Lum9MSfM81qiEFWPfkOFtAM6jaeveJwGqksyURAbG+KyOzH
Akg7SvnfCzUneejD9vJ+b9i8N4xXlCeOCNwBFEXNzPOuZC56fNFxBvFvI37eS5ci
MpkXhCud27T9/V22aEISwmYPhxdP2GQPiGrEz2gqVKA5r0p3VugPQ/o8e9bsSW+K
gXLS5EVV0vss+pE7h8myY4XnOC198jZyysiPmlVOaGjjrOHWt+cjloh5bjXYmBvr
muizk+waN2/1BEY+NSb+UIROrKwEB8lq4DqzMDL/Cn230X8kFbw3jGDHAT4tCCH9
u8JnLujjJeRwoWTnWdzMaWykrzPPxOpsxN1jqgqF486vGwGeyli+jylCJmb0nzb8
c7bBgc+kvKMP/wqMQad2n9HPmbe6HOxkucNCgBpBL3f8wwB9eh5uEOwA+ScGc/0q
ftPtDFTqAcUih4G23qBAXwcl7+8FNKYCuVIATThyDRAvyQZgJdyBgWqSdwG8iZUV
xbYz49uusfCiK2sTD9ieK1zFnxFxHNwilampVrzTALq2N9YHnLjQHKFq7jdhysR9
d0XTcuobOfpJm4DIyTUywqwceSr+tNFnreoRZvyTZyfMW8Bd34fo6HYoHfKWFP7M
sq4ddP/pbOa/VrPqHgsyarrDnf4V6CaleHm1vRc8it2jzE3h6knD8OMqt9ANAwxq
gz01cb9CI59zC4+UeDzPKMbUcWErft+b9YvfA/qaSt/m6Cufc0uNwFf41KroTUiY
VFXi1WigYzNfOHfAsDV5vmVxYbX2MlnrmquNgO2gWP1X9nk2TUOxFgvL5+JYLrxX
iip1FSWErdxUNzOvg+/qkyBRMVdGa7B0AQbttxe8HTuDF7HDDPK4dn3XR8J98hLI
5ui2vmhtqCKIiGgZUXVaryCOn9Welt4qjwYYXw2PW71SlK/slfj/OAlLIKsOqiJV
j0Z9/kwGhBOSagKxXpv+s5crAUplqkpb/iMTg3qRhHJHpB4pXg0d6SPvvOwo5osN
wOy9B380Mxq+kiEw5py3K8E8X2T6L64CSAO7fG0AifrO2RrMpDKOT21APLPoKkWQ
n8JN+5EX348a7oltW8G4cG995caAhyvniSQ8nnfX0jJ5v5QWJwWBoauyKPcaDh0w
MQGsxQkI08eGpz7W/3bb1T5egclKDR1R3MkjwM4t15rLVQnwTSYEuSI6Wf8jtOfu
+bytq5wbs5IiqQ9i9kiLq0JsqhRp+n6QkPBkvDYJ0sxAsQdd8+9xpQ2Gghi17LtB
Ww0Hta80mql8ENNim6qpGQJBgE7hW7nRH+tH8JIp1lH5WQkE60COcmZaA1sX+abC
n4YGnH8tnT1dBdzKIkLlmKEQnLIaZN7bCxcgE117bXopZ3bvCBFF/9DBjRa5u1kF
ONnl+ko2Qe+I8kEb+fxN5yuafSIjvRRkk9HttZE4STZilwHfFbaVw8t6o6vk61Ru
eTgV7wQimHXspuUEpobuP5l91+ownkshN3+975GOOmnnFjJjG5AyUYO7DPl55pRK
wqUaDNO8dCSnJUl7bFmm7k9vYk2hTO5IVB1p7PlBzkCZSmlrWAy/mLSjnD1/qb7y
4cVGrpJcgeEWBOobuRhv3M8C0ajQYzAUbZsMGgJo2S22Ji0P+F5jmIH8hxUlMvaf
Pn/YrFsiA35lHXVsJglDDfuArlDfIKuQJkHErZzsHHKa2zn0zd0mOqbyCMJvdUA8
orLjGbsxUIPlqK8eVKw4kKhQZkCl2kopWQXHN3mY7oaOJ9PV4rZK7I7hrhhVhWvZ
/+tC0NV2iGZ7kGyAiw85qCiC2+o+KYOegrbBCKrHHIN/3J3t6PWF49/gYFoCkZ3r
+uLEZnHesGhzRepCxEbXpsGU4RDS/g/ONK4gtwYr053DH0amItgspdWJYJnBhLnn
LA4a0ymvFwyzX1AYzU+L1taz06lVF1pw7Ouuzljja8s8OGqN/3oj+FFPi1UUUkkq
Vsx9TNS4ovo39rZ5ZNp3TwbVO8DhZlFHmEPUDOYr7UW1/E0cdBSPxXmkwO2stuYi
6QFiRUknELSKQKtIyLOaS8kUnyXsiS+h94rMsoTAPwRcdHGVl9an9sUe99Pe/3UU
F6LgxUOEQ8TwHaNkyhqUXAe8L7q/8B51qjLEasqWIPmr9k6XR9hR6KDT8LSYBeND
r5FTzvcH+vpwLiEiMxnpGD+soCpGNLdsDLoz5To/1Rn4XeIPcVKfHM8wcLrA2JFL
3Qz9N+K3CYhtvx2MiXw66OYO3ltv5sTpL3961pWUb/TkJNYTKMTZeNbyAQCD9Bjr
e5xzDkRjyYvug/wAGoraG8tERRKnRJo0beLwc5ZEgbFB/6EsRqRZESOPjFlU1Kod
5jVO7onqxlvRb7FuKJR6vNNqTPPnDeX2CdQp0IzK7z1FbLjw+7w72hHDvlX/WAFe
5IPRVQXdG4gP5bt3rONeulFmoiocMUo8pdMdhZNms/sXmEbrLJKuUD1I8DBVsDDJ
t1z0JrrFkbqAgOrZDo/k4Vy7qT5a1pHT+Oy1/m0JcC4YM6mr92KlxKB3AVQm8MNl
D5+bj7eYjfHlTFU1N9MCVtTW1Ad23xXIjTvUdmkTw2I4x5Xgecu0Nl2sSLofV9ne
ldjjRlWveOMMrgmqliXWBgJz9IsQE0NznL4+NmDTZXIcWzBLHANMLDoDDPKlrTiO
QVvafeFFZPw/W59a94IGFzWd0tCW2V87OTT1aN7QqQdK7AwDdIr3ZEv2Yhlb4OFH
Ar81RPAcj3qtKqumgw5rYkmWbb4qgUjn/r7ZXmi8xlCBcNCwj9bpaIULOWuFQQnD
+70/VYJ7mUUUzw042aMC1v8nJvqGkedIHULHQ+/deQcOYICsGZXnobIQhUSo4Cxb
dONJ1VGp0hedUwRifOC0BAv/XrBdq56JG69Zdy4B5QkKajHKChSv2oKzKxUYkANn
d4rnRiKy+kfR45pXBPYdSYmdUBkfxpbaqhLZ8jVME4rzrfiNu2sHHjU3JjKNgUXa
w4rKAHX4SfATmEWUaN0v4bTLa04atyPaJYD8CD4BrGrV2nC9gf8D2Dbj7PUwVDKv
HrFklsNBWIvTRzZvX7gtUXX7HkmEptml0MtmdjRvUHh4A8JVm9rKfSwTTv5NlPUL
9QEu45vN6SJ2WC1Liim0vkFA4YzyQF0Ed5To7k5Dp/6Usrca9JwcUqL0pfO79jay
1AR0vvHFi+hpgmK3WgsPdLwLvXSEL0pqywVFf5zd6FAdkjqmwiiEypbKrrbHVV9q
CCVbcUYFN++kY/au2MVhcYS9JphPZJiYm3N+/12UFBhj6rWQjdQm3F0pg6UQ78yF
nFB0R0ozplZYCERSx8rdBkLX2l4aEyq0klL/M42la4cu4fHE53BkwABMTSXOWhpx
wV+bStH9hheZ/S/eAUXtBlp0eysSa/1uqSMfFJbgyw0c8cJQJrjqOKBhDSqfL98g
0FxbeLMgRxjLeWaPVfOtRkbWnSGGuw9q7jGLIUCe1aDBgeiIYKomWpJ96RdB8SmS
1igI2O36alSMucBYDxO3GDd57tdz/z1o5Y9PqXh1+7yCxNY9DKkvv1VVGvLSk1yo
pyDrGH6w+/ipSfYlc7prvGN4cGM+YyhCUjKugQpIx0n3RGRqBvvKyRHTnxEQHWDh
3LlL4oSddIGk5+oNj+2x8C7gO3F1uS6z4eKYOZvCtanTG8qPJkFDLZDbAoXNmBLE
3UUMHZ6dkx3vTNF9weJa2joD2o/BcYzLckgbnPOkGftZBe0xrVd9Mg0o3JbkJdi8
SpmY1/2h/9kzleYtq9c5zFtVPU3e8oGo8S0Xkup6Ma55CwJtphKMS2Rf7ffUIJXW
NZOOhyfaw0kihLFeG290Mh3ivr+suBBW4v1K8Oo0SfcnltDgOvgqXoDUNV+AP0Tj
uyCM7IWwelYfaWVGZXVKt71bxgxCtwE5Saam7zL01Cnbwn4VST7khzjLIbbwm3Af
s/5U4OIoy7thS8dxGvSmf70Q3Goj3YV9MXPUEmORo0KGo6Dp2KHf3fpOMBkcXYdD
mm007+8WFcUt9Ffw/Wjt8DSyZJqDfOfh7J/qw7sysupi3wL4ieGOrD9c6BzRDM0Q
kgELSxm/8iXMG+aHqKrO6jti4kQ5gmlh9C00QYiRs+iv/1OlMmrBd5BvzMC9NJ1S
wo3Q6o8gf0gydqaRhe6/v0AwcZFEDqbXk9yxmMSHZI6FheAYRCoHoO3680lv7zVX
RfvisQUa0AtOxB0ze16CneUyNidVKlroUwVXOVn0jdrqgWDfbrYKvW7BaVkjMahN
6WYagHBGb8x42irntm4whrr+Xss1NVfJ+u/w/I518esiiGwIXHUApvKvE2lUKGRU
0hcm0sLE96mkjPdZUs5ir9+nVfcPW1W4lyu9kQ5Ko0Vq5tQh3YLxYgEWvk+jZToS
Taikw4tcnhsHU0khuKyTeNAPLnKkY8PNNmOtFaV5BjLh8E9ut7WxWfklsU02Nt0q
sQHzC3VGZc90PWfkctZVr3+RL45Vd3k7pob4LmIO8kUsrZT5XenSs4xvWqLgOCLo
A3c/7npAktO+AwS7l/cDk+rUyIR6bOS+qzR/s/TV8BVJqHYoXKvaPljmjPptHskx
40QWfxAKyJLnvwagWCwKqr25q2iejKl2MB1KU38S04oT8VaDfvOekZL+FsK4CRm8
vK9+cLX1VeoJgdhkeqXMior/bzFMkfOgH2Z4n63lemA7vAkV/1Xs0ox6AKVbhVFV
YpLsVqC9AYAg/++QpwXvG/0aF1PN5ZLJv/HrgqB4iA6198Vy18xtIr6JVuC/ao7Z
8zS9yfmoI0THHBWfIREAUcG2F0MiPq6HoYAza3mPTSkNmRTc1/B0XY1lPm9WXeUj
LCEExysdMcWAxXSdUQF/Ag7dg6azKkymUtVMCKxDjJWf68yqWuPqqhOkLmMwYSt3
Qraw7Mh9IPEZ1W1tWYoE3y3wTKcRCT7xBzN2yPooP8IizshSrghB5gbFCH2kEC4x
2gqXNg/FHCsBCp4uyuNJLrEOzxYf8E3Q/Xbn3HD/Cri2lrETchxzWIMUMbaRZsRk
7xmNhleJNEIbfhAnki/islBo+cvUYd+Q6G4yy6/9NHOFp90delLd4D//Awi/z8xG
1DK694K8c1HTfIazP7wxV4fyd3PzOdA51kjJCRlqv0+5uVvRoY5JGJN7V4x/uxkM
FbMD1GhP1mKrD82oB8zUkqgGj4IjnHxAFbIDbssUIAmwIZFd0xTIhGbzic0u2WjD
ikZuhm5LAi5wQBMqye/9KahctF4YennKwhc50YIFLevMX3W8MYYJ/IXT+mGBrdWn
gQbPqUMbWPkR5zN9k5ON0dPtuly7QxhKeXqRH41w4WKCAEq7hcEiO+tCR03WrslJ
fPRq2UCX6YXAXTWPlxaoubQTfWh8G4Y1wG+txorVFIvICXaVQwSaOmusjKiuwNU8
lNzK5mlwpDaSqdWtN7n0qDZSoPVEPDnDyJjThryo97jqh/L8lKb56xsz+5R/VoAB
xJz6Xjbkvmv/VSAeXaCDsmi6Fc+2oYHLP8S0zcZwFaQWRtD/m8Ql9NlIzAdC7b1u
jUUTgVolQGbyRgDEeQeWJCyIcA8dtt6mhzdBqUGUAjuCNtGtehgqPKL7o4pIhyHo
ygTnDEHhsbi8Ym5JN1U+5BC6w4WNbYNGyPmVYiMhGCE6tjglTXJqpKY73zsorXV2
675IfylB5QZj60nAQgP1U70rLTtSIEO+5qTrf7eARUUEIY1pyznJFmUA7VtZw/Rs
QRHvyb4/5b+ecgoO2dh0UVKK03RuBP70515P1WsBbhYiuUont3DT663FXvc2UX7W
GEv6lm0zNkLfUgvXaN1JXkFHKd5rYKPIteCCVAdkp7kXAyDTwPBP1zHoCleg6vL1
RFm5Fb/h3iVRcrjFbPCJQAMMOb3tKMkZj8f2RBQThItVBgrRBWGqyHhpS5636OYb
KT3zv4a2pqkXY1fiJNgfrq84GNb9fe7tzVEwV/eNnVwBBeNCFAxlC1mtmYn5aDY9
txn1a/Z3AOqyxlBJULXaB/WZUjMqiPUWBs/KEEJFfwuTJ7FuQCUCuGNrEoJqeCLJ
b4WlCtp383rjlzvwAKM/GsAPdEv1Vzp/pa6C2+Zg9QgeH5/o9PjMA38SO/kMEu9U
84xBsINrAMr6+nPo7sEWXqZ8t2GSsGAjPO5QOIAf41axLKfakhCjRyHAVXiV2Y/6
L0Ye6SHqWXYAY6RxkG9hbUCHrN1CpiHgGm7tuqz7RbGZbhqTaR4XkKH6hDsh0M+H
ah72Qf6bbmjYPu96O/nr7o+1nxcYHyoNI/fWwzXNDFgDhYR15c8801L1FZL3TIjh
GZ4sSkIwFAcHxpD3r4KCvhd8IeWUVhzanWaqECTFssLFAaWCal0/2qq8NbPowdxB
cd+TS8NAS7BRO0DTPR2UflLSdY5e2mfz6/Ug24EaoSisGW9zlrCJuj2NtpMG+avl
1ZvR3tcTDIPXnqeneqw0mO0Th5/gAdetESV8QNN/CTS+LjHYpZD3xV2FFhbnmzcD
6nbNXorMU0TNNdevcegsHZCB3NaiSsOZ5hqq6CE+PrHSZUXS4+ej+dnI4fwyBOiF
cOgnx/2yWlae88GxV6jCeGFqJn70wwtQcSPymeEM6q8FzAaws2m1Ge2RlPJpYib9
Oz4Z//wr1cPfAJMLhTVJzAkd+9TTLWfeZi6+TjT9Lx/hTs222WX95SyvnR4b3KaY
P/dPACKxZEwLJeMnymurWZlfCb93Poiy+hTYuPRT/yYbb7jTdrt+ZtpSdHUkBI+P
dXJDQa2GuwOQEwuUMgNR0j2Af6pbyelTJ+jiqdqJmJMh4eFuDc5IgpQYUMiZifhX
sRCraBLlReHsNTcEAjpUfFDHjaKmhiMcW4hQ6ez/0DRe1AaDUACmieH0lhP9T+AA
QomfJtAJwpZEXNCLxnp68hwrL+ilprckSQs603DqagKHoHeD+SiQIXvcSyMt/SEO
9km9+BHj8Gx7Jlf5ezio51kaG3Yulnt3cck2GiIFWWe+cCR5Zu+ld+HdEhlVFe+a
rFvCI2rcmrZW6r3xzgY2fVMDlBLbkUliGc1vbqt7zvhSC4D0IOq6SJ6o/KuqF1wt
pn1JuUGN07rFAbwDC/3sGuDoNvHddQUjl60t9zbkkmLWW/0Zpnl8wcGZl7tcVZsP
eiOKDlzOU3d3GpNOwDvM3PSH52iNbWowgyOCQ1akzM2Kz5Ion0n685AXLXgq2kvD
lqVHoU+qWmmRQT4va1bMa734GOeXRO/ZuBgvqIWDbZDYpIQM0xztfGYik9on41r1
ep72BCliLIvWmVkOOMbR3afbm7Nng0hE4I/hX/Zrg1eORO10a2uaRonh+Acv/kI4
QilwJncJELnF4vcpq5UdeqqXO/1X2RbRU5Hj2ELe35juG3UaCgfyVl5DFZOYrEm/
XnkE0T5o8UPtSXRdZwBS1tAO/4DFH+735vCj0DvPL6ClZAxo4Swz8dOdLuz9Nixd
Kr1L7RB+KrIwcW/ozfTE+WtJ6O/ksWrrTCSuxLg7WDMi2PZuBhTOrcyJo/78TZy1
Vzx8Z+ftY7RxM9NkFIhuk/IVaRgklUuhlTdA6cM3XeTV23eRFqcDebvTUbydCm/3
nKC//y0HnlLrf3f8SmWBefsSkUPGxHBIVvFcp6OC+BVQWmJbW4HG/sbVkDEs52ji
928UVU4434KFGOXhfsB2kbZXTuzwCb9GPHyN3ugya03d2wz/NHXU1ntY5/WrAKLp
M5b+WiSGtHI1u4AKf5B8dqF3gaTXkmGF3MN5s5i+uDP/vwVaqzCBN0dg0ek/SZwC
7E7jVIa/RhDGkbpN1qUffDVScEF/VujXqBPWHl2FtoMDUQ5GcvEYdDzCA5QfZUK7
qMb4pZgfHXsnPR+m00XlHkWD6/kUfetxI83ZExZRU04UuCL9q+ZQAHXtJYGpCu4F
yts9r0trQO3NAPY9VnKS/MgEgWIzaPzxOE1cwMqJHoc/DTLK2hOJO5lxuwdxcJ5t
jLXa565XHHDlaHHw+guOuAWPZzrxXmg4wFJVmkc5dhEeyf1gZK4NnDx6S4NzdIVM
yEwbFj51c8XBJcRkuBys0pwWBK98Fuz3BnC4dZfUeAJysr62HGMdKsCjogMuRQjD
LXzcFFXnjED8nfSyairefZrOGcTa3pOr6rvwP4CiJDjK4REIdFu/hAQWqTVaKZ9+
Q4CoN9fBDYWbFIWQSLCaPiPRQ2GLu2Hv+ZavMIx7tFmYIR989fpDe2eFKMl6mrs9
Jw/TOxjwuX9a9sRuIPkeW/GfHc323IpWhpcgbhnUnkoDq8l8kmSFeMix1KW1D3Da
K2huIEAGhYnB1FVyC5o0679wGJwCGm6d39s0Gw9y9GcS/esBXGF5wzb6ZkD0sEs1
V8IzXC6LohW6W4eLMW9Le18ESJPV5eG3Bo21wmzIjUwGPvmooe4nZ9W6Reg0BOru
c0Jo3Mh1bKqUrvuPgxYaWZigIpmFDNPYJX0k+S10UwljJWM/g7OKUKXsIuM/AE8d
L2XU5Q0MEl07AbKUZTlpz2j0JuKNPM96WXIU64WnTckl87jJaoREGDUuyN+xWy/R
VGq9VZkIKhVlosCfNOoYTM9MjbCltPPgmq/VdqlB0eLF1cTYWf+xRQIW18QbdEQ1
sBvJAwRsCjDnuHuop7/9TTVv+dbVNYuHpdEWak0euxvfUA8pKaPG1D7EiVY+xhrg
ku3I1d968pvjJgSERn7zyBy0N7Q1hitfmp52v02lvrVc2MkZsSaFahkM0UfAnAuj
4NuzcTTEQ7t8R9TodaY8ywqo7dl6LSsuWFU9fkUHbyPJa5n02KaI6dGYSQ7AFI6D
DFOKte+igGQdantgf/ydTeCAdkaGEG9BGx9cAFkgP5FrYnwyZTaY87elY2LkgIhP
EK6DX3jiSYBTjsQZ3MszJ5sfMohSOHxpxHAnwp155Haxg5mArDZirMz8R+qP5jY0
gB8OqoJ6z3yvbcbb7qdUMjMBClmgszkRhwcTIB4r+tqTApROTV8BMBcYKLSS07rW
EI8N6Jvad4HmBIHXYwFlaSjCrFtPYylvDpJ9DO+Z6C6CEQtr2cbahFGq5au3j8Gj
LdxPVLQwNFaoCLBjwpup6pICDb2hpPtifo7oM9JADhFgR6wBm6NPbijCM46X+xk1
AMi45ahwoH8bQ6/88THwpO7L4y12+Q6RdIylwys8jslH1DcSlkMOF4P77JbyvRYt
qKxCopEnbygI+oEuzG/TFyfF+32Hk4lY+UDC8F2EnE4BvgT1USXGDbyXa2ecydxA
jgcCra2l5XdVXmiEJgi9cmObNht8zBA1DGmZaFlPz9aGacvMBC2teVT246LHqGqc
dIOR9R9Ci58SMUtgvfVoHifQuiE6YSjQZM3c80Sd505HsDTUKvRc442RpOgEa/ov
Q1ZR1IBh8XTDFNhXngvVPwvE3bUawJj5vqmAb2vh/4AKxqcWKW4hDl/rh1CCz6MN
6Y8et6G7/5eJo/fnwGGnNDzL+GHHTnwNes0XQ6FmDBW4KuVFmi/wz0u0UGrvi0Da
frkrR7LJpY9oMmqy3bhcXkJ6MRtKz/qBmZCF7SxplYNXcxU8R2rvmtlvAvxAGTFP
4oKwo8bxHHKd/YBzIRZmHvW3yTdKbgzfW9ZaOZz/aQXR5Wg6hXvGA5Z2HtIUNOrs
uDf6Lz5TC+uGSVlx+oCFsCGZpBiClxZO0oRnnap1rWxOKEKUeNCenvjHNknvaR+J
mAscjKy6slA/mowRoiH70rOlucHuvhGkhHnp8P0IvKQkjG3IuKRHg/rSxGqbgQFb
t+B332BaVbrrdde9mWfEdmFl/PtJ1AitSTev5lPbkfsVPxRh9mi830y2cObUXpdN
RsBLvQDF7yz9IW8ORsJNgfwKPFdHRUAI4yHpzsUHN8+luQNEMWlkymqYgUJ3libd
GNqJEJN4lGq1xNyl+kcths2a071jCfjOgHMf+kvhf8aAVIKplX77fo0rrq3pkH9Y
7bkEp8C5G4dxmOh5eQeVJCW51RwNUB6MD8ltPtj0Tl4NfdcOICBbA7vmlkAenuLv
sSyFjMIqypZsE0y8jTC5J43a4tzzStVpBo3uDFjAKaJjlXImOrIylZ7Mvo7gQgSu
REoZvWrSCiS4JPrZbW6Ziwl+H/QY6hvOYEVH7HHcecJZu0x5iwkP8hfxC8bYg9sy
cKtAh0MkXU5ReB5SSgomldeQsHWfnmKGTeXN8p2lcPpoc2JRAZouCevuvvSZyb0t
flTFwSEnqEi2MYarTMPTiDsTVuZlThi6u6f/LxYFQzX+yMHzXwPT6sL5XMWBKBaF
eYHsi1sg3iagePbhZCucYxxTsh8x4H/L3al97jMj1+BaaeBHQxF2yypvIUNo+Npu
QShCS9x/NFnw87kioI+LP5yfB+wygyi+44AYKRHbrC6u9Qukzy02rwbXQLe+HaxH
oEz+CZD55xE8hp4cOARPKlAAbrHohGgkut/Od+cv7x/9ehdAZ5fV2kN5i6HQuzea
yqx/eHH65Z7XY2/dMrCd00/qRjHQFZfJWOmjNUA3QNieXx5Hih0NKdn8/lS4YYpj
sDEFzNjBPU8/QaqzR53cNE+o51TXjd6yrntjA3yiEnGcDTkNPKZyruKOKJAVyPim
Uay38UyMxipWHmWgYw2Qo8jihRXmv7KRsOqmzMEZvWqooGstWsg9EJZWn0nzdA74
/aKLqNR6NY+/rr79mZbRiT9+UljTM4DkCPiSN93qePn9EvIo9GReKQWmkoLp+YGr
W/bHobM03rKg2EAWKNjZhf/NhzmVBgHQ2IhHMBn/BhPfK1ESbWaw+Of4b19uKPcU
yqz+BT5z9KWLUBpLdATC+ADP7WIvzZipH3BfAZLfExV6eNCLDVDrw7WcBnLlc8K9
y5g6Fl+yGbJIyb6zcaHFlA4pPmJBlEMQGgA+L6tDxbEudPo3+kGgSe45gMA+aYBq
oDgVbeHYVAsuNsKPQfUrpIx+q3Vl9nKMHighGD1NYnVEMTIe1cxymuI+0wnlZFzV
N2QHia+OJsEcTked8IlFH9ZMBp0lEsag+OyBpcehkSSZ+jlmw+FyhMVBFcD1XWu0
M9vDgBd9OoG48I+LyDybaBoSJ6zXAs1J4WqVM3CNxgLyWFS2wuu1OaHhMZHaVJEP
CgVRb4gbGN3Gceb239qxYdknjJGeFkduprSFrya24uGKh3Pm2/hClX3js4NX63bi
qsbNGXmk3RJgf0vDiF8GBV5y0Ak7dhTrr9jp9POcJdHDnYxRXxXu7Uv9zenuzc6V
rLd+B98CZU9MDAi74uLm4Y662/VzcGDcUXNpZf2xUOznW2dk3j/zmaoAB77WBfNs
bo+nLojhjvgogtlHmaTwSzOyaGQw/a11OVryHNOxXVS+dW+WIX8GWTovVc+CKOpe
WtKh7Grsdqi6BSAh9nwGyK5VjRFT/GkorCNExfE7Mw44v7owoeLsk4MweeXOOWM8
FzyZnGLSPEjyCp9QXSxlbmr/ddal9VXjfMFhCTaleIcVPOMX92CPcA4MHwBUwYto
MmYRWIByv7MbEzBydxdz102XlZq5Gn+mxl5Torv4Kar7zRSslvrgocV0Uxp6eG2V
rPYKbl3FRwlRkJPxnXCeRrKLRgAFzTv6i+lq71VpA2t4WlwjIcozz5Ln5xD68ayY
AeQ0e4jl9aSfZUK2T1YRDUxM+/ft3W+T0ah2pZod+c6CwKREt4bBRV11eUou4M/S
e2dupbvkd80xuwUhjLAE85e8+I9gEqi323exe5nRXCif7wHb9Wd9fPaUjqdPbJdm
fcLI1MjsXh4ECfQobBTTc10dRSjMr/Vs0KxZVVS17+YF1sQ1gCR3m6b71LbG3NYV
YiCPg9eEoGxp52yB1/Qzvkoh2V3gdz2tzPH7x8HCZfTi2ErX3m4gCg0Gg4G4HWhn
1ZgavztCLa/8eDVctFxvPOoyG3G2i6HV62AsDeetWwoaaWFkXAC1SfXplt471h54
m0zlO8NxvQBs51iHtUFBAlgWrftqSsvOK0MrYG4yQTkn3BSxJ9ZCHcdsC3iNo8Uf
z03U6PYudenFlQsQPTCFjfvHZ1hVQaJvBhv+SGR9RbZNFNB5DAUEKuf9mypKmgeK
wDisOkNe4h/lv9NUJLvZk1CjIZRlBu5UnBLX+IIMX46eoMrIB+0vkbKizSGNZl09
SolXy8+nnKgFWr3EeJZeYGvR3xyP7hrjBa8NZ3H2jh8P9p/NnJylt8OCBMahWd70
K+zrV4WoTJNR401kqxrgevyNClLsv98GgqWpT7pQmt1Gw9HWwaIZGGEVokran2XP
ggr3JJx19khkEur1Cwioc8gDSl3G6ciAcfP4oTbbdkhOyoOdy/fFcWAKGPCZwsDy
llgyqHmteW7yNzHfK0egr3tCH+bIKPeF0oqjatXl8Z18nMAWSFtKR2T9lrQH9pUv
2Or3PK2aW7dBsFK2yFMyRFwoWk3lhuZhb/uqSuG+2xQ35/PUO2dMdLR+mJW0dYDt
kKG6Vjpb2aHDwTQj3smB2G+M+JBgqL5zraNqwjbz0cnZ8fFMnD99a2yZGq3f1L6z
JiOD203hihbOw8JFDbjjs1FPm0M3MjSVho4NeO4PPlRbABi4Ob9gQzqYEDPrAN5r
xgrJvxtR45EVh5uUO9Mk/5+ViQmukdLYBHnlsImn5prPmWRS4o0wic5xFxNHjWNo
9p8U9zwSvZ5rKdDGf4r9I2x+9oBZyfBcrClPp3JBN2ItM5AUfVK37kIC79FNuC4N
me9e1gr0J0eypVSKgWemG/g++edn+PjJ8KbZarJgdQll2k25jsiF8GoL46rUXHo2
XclzepmZ0y8H+pBzu1dopWvZVnLgbwKfpkxStESmithOu1NbcBFzNDS9B1de+Vf2
dIt5c9Cuc2M2O4ZinPOjv6Tezs11CdgJ96sC/y7urNgyTox7IbwYj3A9HLoDbM62
Ux7E9cSpZLtkeRjg7jjvC6VrrT0lRYlx5vQCkHZ8wTRQMobrbClTvI/0Bl/eFSst
ziYct5PWU7N1fKQQ+7x7tj8rE2rzFdkI//sne5dfuBVC8qHPp/z2bYKvZaQEZrx7
fwrmFwr0wvP7mpJHhli/rSwU7RpkAIE1uSDSQL7drvPWyVIir9touNVlxh0Zq0yl
iw1aOcz2UyzPYG2d3o/6xfbCm5nT37Nf9GJdG5s6sh1MTUzLVPkQRUJVjPu+9MsS
SONRnjD0tWL5NB8r8qGZqc/GRrib5JFYJKLRVzxTblGSYDPG/eN9mKKvz10sXHaS
FMAClkaGpe+KzxMjEinL8WWSTeLtqNuGjrS3mafcHVQgFZh8uvA9rLb/Vqdi0cmT
UMdNXwRPfQ0IDyD3NzlQvIkdBeQePQXz+EDo4x8trU+fP5ACFHnE7yD4Obqn7ddq
1asC7TPNn+MMepH6fEDWJ2cBg1EFzeFCIOsywfk9jzhHkxLRgDGkKZO6I/pgmEjZ
O0Ws3jSuXRc5IeDdl10R4QGfgQePTev21PH+EbsN1I/NBq2heGcSIu01WHdYJ258
UMjiuP1Od0GQB9gFp8reYxvOJe6Pt7Zkn+6NJI/uouv2D7jN9imvvaTcb1j30bzw
g6a1BlVK2SFdkfUZ6dgIZZcejAzLFi8s/ubibamHmfzg1fwiu9V26dTt57OD7OBs
xdEwe4tnGhmLIDROPw4GNuAFFiml50t89TkP+5PPaURGk5CRFYiyjjisPQJAl3r9
kS9rtrUbIIsI0Wy8rm4G6VqUBxOVsaSvvZaYcRQi/m/eyMbBIG60GFBm+pRqiFr9
cF0fSHYcI/2uakjRr123TjtRWd6gtH1IKxcZ9wAtok1Is4899sJ/szKzQhY++dQ/
4MxUKxIsTWcQmkVsxmTY8IITWLEyPstl31Juy4be9qTlSNPD5ri2dBub+wCfXZTH
0Tk6Hptk8GXETWSzFZYlgJQtucdDHA8I2xQ9zuhvFXNdQs4IRBqbzdSiE7QMrR3k
1nE9Un8RwKVyc6oBxU3DYSeXUcWCh7lZsmulrxuHdXmyKgZj+uqHfhRl4HkuTdDN
GXYDX+jC4wjX77R3heDxtDT8fHt1HvaFxH0nghtxcFDApxmHWGG2wnhL4B5LweO5
b7Zg89IEuTjaLMiC3v8MfbzRUyN4nGYBpuPrMry+xjqad6UXWxyg8NpSVOU1JCmZ
6MDd+uLDXKe0LaxsHOoFK4VU34YGRnuANuDqzBtkbLmrry4h1C6QqXkMHfdU/B06
N4a8IufqruC3c0WLwsprcyyfHW8LwcJS4R1jcQB8RJq1nucn2zMD8TSaT+hY7NUf
9se7qc7MBshOzf6kHxWRbQoJhmZ9U4eHDSbrCLzuHQ64A7+0DR/svpbUOeVhjIi3
3YvsekRak6cRxXqUlPSiAp83Gfudb/rHfsICMCUH4imEBctw50p+P7H0cdbOLQ9f
d0CCFFEPyrrwOn7fKmwTQ3oRgYNrupUHILQsIAB3dOROJSNKSrOtvls/7N9B06Nj
SldCvf7Qq2f8QTQ7O8mMLudW2XR0kZYXR4O0JsxLqZFqSdeJwoMN27I7x0BgcBRa
+zPj4O1PTKmKxuFf9TbolRSktegatD/gkPEZpZDSPBFgwRORIpLTA4Q0Yi+c8f6g
DbWAsbdJqO+SNvZsGpC/J86Q26nkEtRtnH/85hZvrYfBNGI5ri5o0XG30qbSAGuv
5yaRxmeU5m68Ca9G2KMRadzs88D3rlGIwLnds2kxJaetVPZDpDZSXycXWMWSX6UL
KLyiae0rCW6eydw5+pYuqckpOqN+y8L6Si0rCtt9eYW8xnuSWvBnXuEGPXjD+WXv
Li0sEh+yc0lNqs2hjlFclXt7TNdi63K/0Svq9HMpikrLcPYn7lywzaXca84vMOsj
7lYJg2UZ79JqJIpS4ICvG0xCiN8qp5lgjDfgshOfqpJvCngqx1vVmyg6HCFmgNNF
bQOhLRe+WqlH0vGPB4zuSTySCpOwAuZmXF4U2JPQDh1aavzRXBLb8QIx9GAZbDZE
wu5h2dW/GosQ1o0TpkGEmOiA+R67TEqqYKw6RTIJ74G2rWyPdJPjm+HnZjTF1Le+
EMVwAxNLqUNwQLe9bXvXkaK0hGosTm21y7QJhM6KMopSuRz8Pe51r0KjDQqSA6sl
9/2brfhi2f3Tu2LMcxo41vAJ86OGV69TWojx/pE4GsaThAETM7mNVM/d9Ku8U9MQ
o3YAFtdlmLW/lKXwhLleNrcExunyBOYIMr7Q/zb9uAtgqiadtv80cgSbkOUkrYMl
TI6/HOOwrwrCBTOi7xXFctZRlricE2Lakj5WL4xmDEvxSDnYkvvSP6b48cJ59n62
Ozk1lxwZm4xmA5yHhe/Lm00sgXNq/NE8Nm5sK4kPleD2i1nR5CVMNrxeiTOTqsK8
TEimqRNWCl4zxC6U+SlRZN4Yz7Oxm/yDlulsCbFANEjcWAFpX+Ysq3UbdAwzTP5r
OVTgd1siDVohSn9AR+ERtGeg3AOcXuUC8jeIT7AeiO10U20gi7xYr7qsSjAtPKEQ
JlT34Vnz4Ru+CLMdoQ2XS6A91mtL5L7ShInC5H0PeKsgaMN+cCeTb931ToO/nSzw
8MlgQ/T8Hb3jxlY/g4hgq4r7wb+YxfV2apkMG5vbBFiwcpK4LRKxeN96U63ilwTV
AMR24GgNc/iMjevn1P7le8PZWjFRHCns7emOWvM95ucpFNW3KlgfPBSM8Qj7IdDO
uTXOP2YpNbIwX82bcDfE4GVDKXPiyN5pxONeQT6WxJAN89kjMOPOf1pXdf0iW1fn
YMn4O9YGdA2y3I0jM9/uqiktG8xWu34+kT7ub49EfTrG7I61jI4HmfZtxb2wPjKf
o3tili+DGMLFC9ZtmQ4g0kvs6psMnF01RlIjLLXBvOBxXIpwLcpIhO3dbl48H2eT
6UhB0N2Qe+A9OS3ujLSQHhIu7gxMQUKqJVudF7jmd7DOoDeP/Bi93rogwAOM/mhK
qQ/kFXm+iIj+oUCbQEkMxtk8NWOtjKvnOicShBfJ2uwv0cEPYWdq18vscy477FI6
8UEYGB3QXtw1IuBVrPYewroJjKsDGo2bw2kGa2BD5TiAC/mk/zkYtNTarTBunO1m
WH7AJ0KYLczIgfjXTQtET/Nls//P3lnhd81mNIIwds4ubtySWtZp7AagF99wMMrK
Nj8JRzzgh8M4FswZW6yEFueidZjCkcRxMVAeYgMbFlIKjkVBAM1b4r/O7G7s/ktM
u7d02ADVlwxRDOnBvPiPjGgKzeEnCM3SuNHqZcHYq/LgyGx3rJtLCc4VabsetQdY
d1eGV3QHGkOsjFBVBRVUeEOWgkNgyZoTypQSFOy/AUCPI5IO8ctsaWGE8veQvtge
oAWiFCZU90sZJXAk5n3nEryNJV8bzsz+3W0vXuDB5Kw47uuZgPx3aMSw7w7Bqv/Z
FCLzPpQCkjsRLiF29hdQ8/1UGHNticvGXlyho9Q1aU+E9I0KV9KlRAMLAg6UZFQa
v1eRddFnc4b9wYHW3bGnKBKbndV/6NSM0khSXem5IUu4AmHseiC26+gdi71bfNNL
w3XGpwVRW5wwjRVtxveI5szwa00UGNqWnCo+qjoQAy0YDkDdRyryY4TMdxPpdJ1e
clA0RU8ykM4ImoLD+Rl89gQMjfDI4ZN5OrNQrw/tR4ycigSCNL1M/He/gAEyk9Eg
MTstQsW2CfcB8aVNO3Bn2nAG1q3kYFB3C6ulr6rF5fvOr2NSAxO3u8xF4NdhmMnZ
mRLcgLo1e5QVviMoccrP0ATYuuW+bnfgFP8+6lXuq4jd0UaET3tzwjB30mzD6K5K
IxCbgH+OaltBOMr1XkWuvlKDjcKDQXvmj6JYBxf2VhHBoua1D/wUsLzvGm/ZImIG
fi4vlrMW8SVD2Fb+9abTmhl/YX0tLjbCrQeEFtDl7KrWC76xA+izsQAIxXhGfL5E
Z27ZDD9byQVFfTiRc3TokCChW28OvLoQZHZqMRe1iB+1BqC+BUnXcZZm9h3Npg3Y
H0tTLaWe89n9xuSe2vU3U6gBRc+u77Vl8cwGYS3M41Rw02WWF3X+VAgL1hNdK7uK
oW7cEFj+PjGTCmPRu+psMQ4LJ8Xm1dDcA+k9pnc238vz/3CWDg0mYfYoYZOa/qKJ
lZZkKW9Y+b4q9AXll3xuzeED0bg7QgPGtk3/FT0YuIG6roqnLHuHstXa5fHLnb0n
7lAnLjz4/21HIbo8I5gWvjKyCarCI4zXg4sRXk+dtDlvV8Ny4258thlbxNp2VYnO
9WZlkh+MBEinfY0RetMoLS4daacvoBob6YbG5U1dYVp+aPD75uXXUuohsL25WQEj
Ik50UgSrWKpUT32ZyMDCNsxYPv9sHyLkaaJ+NH7rq/ofrbLzRZcjbZcqDI9WhloV
i6OLGhgCvXTzFsFiYrf19k2kQBK241zXsOYfhG0qHNeUWyFl+89g2aAQk2eEQ69u
IjHEkVAu1EK2A/M3gf7BOETjYdjcf9XIL1HVqpNSMNpJSwRHsHrCbtvZFvRrMuAp
HpTaqRX14FTxtkRr49edwpq9ZPdc1g5OV1LB3oB6Mxqn6e4J5IH+c4eTFrHvVMCu
zmiv+/ufFQUhikhsvx6oTvMVVTRHZd+mN/5ihJyvVUwSEoui/dWBDNbcwy3lGZTC
jTVXkKnoWIjUL0G46nKjD5FmVaOH+pD6aKT14WZDYo3zLQ2OVuGGq3ry5q9n5STW
EhtzyXPOpIaoOk2OXdKetjnApduL6mghzA627WZAKUIxBUESGIKejeT+U/8pGwo6
lwrEBYs4GTQyW/RgPxcF8EDCzFeyNrfTiw2HEDje51o3Dcj8M3oPTV/VWE7TxB54
b+MY8VIRLUqHmrfnPCiQUQoT+DAhjet7yv2wApbmdSmAb9ff+ZhYbXt+YmFiiMH8
HFDUPhYwRYjX+LqotTMlZJoypS5DgYki7XvFwvhIJIcuCkT3jok5DPlFOIiF+uLg
h1WaR1jNIYISpahVrIeEAkH/4U7gokXGUsJFs3/sfYfmHXNtgPuQKRYG6cQxT9Vo
a0sJW4cssW7l8/bAQc3UClxCJ7nAqlG7V/yqtOB9tjlrypaDPfgeeKelgOENDQaf
veJ3a3QxaIqw90HaA4lK+VF42q7peH0waxptxMTtosS1S1TkT2QVJMo7mwzHIcmS
tqA39ecCfyBh80FyJaU1bhiNNo/DtC3guRAbVQ2qk7hF5FcPlmc3i9kP/GO/Kzrb
teSSU/iAPH+h6AF8i/FmePBE2ZhoUDPiEX2PRdJ13LHJ/Z4U92jtrA/VuydJ3RYQ
t4q+rIo40DjrQ2PszpckYGSzsY9ZVdU6GBqFJaBH6k9+4HfqHZbzzKsaiYRiXwPC
CseGUhKDsYaj5kLOdBe7MYAk53CEsGtCl53p5Mz/9TRPHtVi/XYBkjLJsYzl/tU1
fzaIHLZwpLlta0bZpDN1EwcQ736YAlfPeC0BDxAdzoUT8ckqv+AMQfTdojPPIkAl
h/eSLdU3bI87TQYEffvkX6GOKHsd7iFFZS/NVq6dc6+1Zm8kJ2jhnm9aKCXhwVsj
vUUfkxnEDy5AZkCHdFQBGVSV2UuAryqYcjYxmx0Nh5fbTL+kVdR7+0Cc5XmpV7qe
P8f+QsZQI37wrhR9ZfT4O4oKUd9W2ybzhZYxdfpN6Q1YKCwXMEbH8dyUHPkWeN5D
xStbD0RjIJDQ5qGOxV98cEupx0q1etQ0H85h7Ha3q2n3zPRj8wLwPQdCtfzLAD1g
yNh+UW7/RyoCf5mxm9zgv+NvUjEXyi/3cp/Xyz6zONA/9H4tqkPTsy4isVFPC5/w
RbFEmGRkW4P+Tctf6unS1BWLbJx2zmNf+fgUtgKzkgwCeFJFm3RX49MV000BGc5P
2QSgAQQQs194CFjnlUlm3SKvU5BIwwETWBV3QItRGcyoyx12JGBF240pjqZtLa1l
gBjBujStuRpnI7UpKdaWNTIHSz68rSxSGhG5AMCgo6nNO2Q4WK52U6iETDjiEMBt
XcH48rTylmH1T2gMn6Up98lGke8hq6m3Nwv4uZFlOZ8XbioMLZ1clQrWReCvyzUS
T0mmYLK20oM6eRPXJj+UmbiD5/Z0FUQoONvAjqHIIqWRqG0oFBm5FgejPu9SNuxH
LrD+FeNaI187fXTgPlAU2xRClgEKN7u9KiCEiFSWf5W5T92D9y5Duhh3q7Baq9Aw
pIyBpgsL3H4B6/gPaPmJB37YCjDIGrHXuqXtMlj/boCVvhQHunnrwmFbDg5CdvdI
G/DqowIjrVGfwutKfi3W7opTUaGex2ufShTCekcLWRE3nIiwZysBkLCKkl0nQCjd
L2zhSBjJaZ35016nY8YID3d9qFdfhAaAcSOSObYPbB6c+MZMtVTLaJsXSvUpORm6
zv05S9nJQ6GBC26nuqS15LHOCs6kAL011sD0I3nogcb+ZFe0QFuh54F+8ussOWuN
Dmvil4UAxSvtwsitzURd4bS+5AxeqB+sgBosN1Po0FpgGbasGtkr1NQ1qffOpkhZ
oIDrYqhczZW543/McrzwV3VREB57FZn9KGhoUM8iMPVaBkiNc6HoWNxEW05w5sHU
XvsISfuwtAe9WZfe65D/Ypfg8HIhv++3cf+sYduhCA6asZKgrDjbwEsVk30rmUxP
BH71O78jtRbBRmt5GE29JXypMuYYEX6EmLgPYfhfYHvMk4PS03iCRQ6MXGMFO7a9
RXkdQ8/BYSoazJFObJYkj40mryN8cs6vUZP8q4qcj2cCkNwBNM8wpDF+3grOVu0c
IjCqOumOgitrcjHG6I7w792gmkcYHyJmSHeoBFSlp3V6lDcjwX/XM8EwOd7I6VRp
Ppp7yJQYE3PV82KRMgbtek6PFdhUO+iV8uTk7HlW5w8I24ytU+V/Z7as2G9DyBVy
tsL97oC5Oo8R1THyoXTSEGSjGXBbwXKBjdjOpAyipTPkvjS95zpgaEjk4b0SncFa
/CZzMO+A451ncTW5iMQfrxVdSLalSTMg9lvaF8bnGYvAfRkahZXlRtrxFFCbTHCg
yaqEFYcxDiGghDPbaQIcH0ekmkuCPYVeOPpwgZYRoW0OuZAIDrZoxNf3FgBcPw8N
rFko4RbgVr08ENOCrG0qkc3rJ9kEKBeEhcSCkDn+5u+GCXQvrP894bwqiifNu2Gm
igUWdIKRqhsNkhNeTrJiCZANmkaGFJgfsOdDiduqrDEFTtePnjxV8iuRX4KGELc6
wM1bZs1xKyaBKaYm8wQubiCzNUqO6V7vgvptcQ2m0Rpt0+BCxHtHicpZrS9B6cl5
wYqmU37u+kYkpR/dNnONKETfpLRreIloleHeep6SBentZiXJYF4hbTa6NMSAbiot
y+kPtm9FWZ6gOAucZxO6lZVBiB593Z3cshXXyr/KBtv5J0DlG9/uPumqVMO3Xy00
WKyUBq7WuvIIEzQvvwFg6wLcSlTlGOFVG4Ky2fR2YDcQVbgwrnX500HWqpWWb6sf
QfemhxBlXr5BKCQPbGN8C//c+3ZvGFLd72/WgpCuSMGhBrcHYm96FkEXAwl3Uh22
vQ6CKW6DyIf7wt94ZlaoHZw+mz1kfB6Brfk9PutjY0njlZK8kCkXYBvmbyvy7eQI
seggNFJTSWhO5/dD3+EP14GOaY2z1vxx8oSkRNzrE7IaOfhbcmuJZ8hjDUMdprrW
Xzc2jRkFUReAPw9G23X/OkdUDUZ1vJQrGrh3qD46ey7Ga+tyGGZ4M0DdumPx8ekY
UhV6ftfP523jGQ1CD1XGzEcJw0tH1qXlXf1yEpjx6H4e3TQb7xu6jkYik9IkrOtg
Ret273KejNuUVF1M9A7TnaWziaTMDHAzFX3zDx0bKglfm1doGqqQ0+//Is+VVECA
6KhsdjhwKUrZON95LdYyP/yhhaaTHp+cG7NAwJRSvfKi5GKIuAiTxY4hrQVxg+qn
F03CLWoznAiRV5lkDd0s6Z6RbGx2oGfKJf01uYYOxE6hDW+UbKRzvK++V2fzxdDx
O+bE6Zn36HWXwJFtpsWJlitLb4lEGqtX+jNnNGoTqtlD4ahN7cNkrNJURox4WMau
JMPwzo0T8Emu/YhXvJe+ZY5mKCg+8FFdX5MijiK6XsfBa2V9Eea7M065UGAZTgz9
Vo8H4XZmaekmyUm3Y0zuIN6rm9qnEBBfCzTUCDegboG3wtbo6AoCyPtKpFlgYYwK
IJKbq3A9x2VKyM/OtD+UcYUFXpMJAacNl766U2QoxPEVjnTFYv65imhhvgKMF63H
7uRXX4kP/PnUSQpyYHlw3ANcwrSpJzss5Nm+BVT43uTY90ZDBsGrh/CuOfDDNOnj
jxBv8ziIVFFmpCHVrdXgoW+ZCDhhICD4ZqhBO/8WNTVxhWtdcCgEVPm1QsSMrdPw
FosMmcswUWbm9RYn74mYlCZ/XzOlblfnLLZioVNtZayDsMpaWiSptmatiwYeyPLf
C0cs7/LQgiF5IimBJ+zETaj2o6waotbYWPfmo/MCIHeupoyfuzeZtzMiOAQQYrO/
1qXNT4wnyvS95KC+b1CYjikIhwRy9fm0UBYjwapPWHD+SRMMJd50b+IICuZAk18C
87cLlCo0U65s747LGko3uYAmJIjOlFAuO+QnCWMmvUFfB6xYY9GSeKhLbK3MJpes
s6OHOGRvBcD3d97i0qBQdKft46ZF5dtKTV9320eI/uQtn/QEq+EpAROz/6LSLxZ0
HE4rxYNiZYM/Vb6HHULSIXVahlWOv5u+/wED56ZDvo17sjZR7nc0AEB5X9cv+mHm
9KroHBDazKNErnpdPIANd6aNqUfBA5KOKKVLrHdF77QzuwtkD56YLXQcSTVsQUGB
PepZEz8WEwrjU1sDnR2yNuo5ClfQ1MsuvRhrE5ekJSjHdUSncJkoHVPHVDhvnF+n
QlsqUJu3WlQpUrCUdRLW2rWgTeuoxhnbQYbIOnz+ZG5l2JthDvV8pnHUOJlMKCUy
zFzeZOd2ALw+eZqx+PE1hHvzBLzewAO3zqPTcAZFKp5mVvZeaeA7+c+hu/bCu593
1YvwNwj9Tyu74EbSTwk6IYSNoMqYkLwtXKSOX7P9/GTPB+wvrRQl+yAfDVW0fTJH
AvJvqQgZHQb9DXMzKiyCc1h6emWcFHyXMgI7eSc5LU81PWKbXxY/7T2Sm5DqRe3T
97G/dqW0OgOALnDYJDrpItaxIgwGNeGhGMz80D+bTwwfJtQcmfghAy3ime3u/L3U
neIuppWQlpC3SjStFggLGWMyo1CbFbFXjLU2++mbmSh2PxhfTHBt54rmnHyp5jEK
ehUb9YSxX4eYSuUIfYWXRF17Ta/1oYpMWzM0wYs/wms5GYzaX+vrNP8A5T9sI1Gj
jMH51teEtanfXWN9QUOeq/8H9t2lWyw7dF8GojETUJQNUzjIx36UZwV+jUqYGK/P
fE6EUTA9yCf2xT7JcuLn8ZYDwpTOm/bzKBl8vUsTosQQByGwHTk3UTWIsdokpM+b
1cNIA6B6djHCYPKR1cEh7q6sIo6oD1xwtDq2a2GqaZwWftXX0hUXTdl6cpdul3XX
5VQkfvfsElxkeZHJ/84mTNqbt8MtpKu3u8qk9hmXeNkTiqmnxB9sVDOupTTX9/YZ
LoohbSolGA1c7DzaduO3k7XQC2SfClEPzNLvjdDkKC1xQOWsRMlbsyo05uxmrsv2
XVndvkIdo5fPJ9m37THn06kYbJqQ2HA04GQKuT5AGKrey9vT3jD1zAu/cOEGPFoP
aHxw3I9TkGiurJ1BsIDYXOl6oUbRB1ejEo4rsrN9IqgAv0KFEI/LPzzeBxvfWCO0
EGp40mclehvrwRP95p3XmPgs6x2NUWrAUpolSHwfWRDBNi1FVbkGz6pRXSpNcAGS
x5JvuRTpzcZtuBmXOXRecvghvWmwixwdwvEUoOzXccGGLteVq4jGIavhgGDYFt7E
wHM3eiLdsXoWjXLv5lm3EjrKYsKQ7uSv35/1xfwjPcjZSnLQCnl8Mdywb12gAuxA
MBEZZm3KqQgWNm/6gtsOLZ6t/CSryBcKZ5u2yafUYLjubT85DDRDQWYpUkw87XHj
C8k8RnLVJV20vT3U5sJq9dotJg5juuzdg263UePWKkjIStE0HFzChHmPnbxCJ768
t1ic+Fma4tb5StrV8nopWkbe5CE2k2vZANwYFklViu3dRB3V013rMsI1KQDfQqDV
TiKaa7RBMwKFUwib7rCLXX4dNlNai+n1cM3+WE65zXqjJPGgRHjFhfy9U9j0lYVO
MYHdX4/lhXzpxSLH1qigPX1i8pBzHAR64PuZU00qrAP/Lirv3YsgMZg9jdlLB8un
qWlPfHx/Kp8ftLbwPDu0/QVAncoWAUpb3QXAlfPphy6UOzze5gpJUKV13nwOuELq
7Akl07zTuowOJHwrYMwaRjKu3p2SDxyCVVHyoCoOICyK8jRoo5hf/ghV3Um053m8
odo+5LwUvDQa6SxZ9LMkCA8sLn7eFHI0ACQlCT/6OVhnaq1ocXp5gZT/dzW691fI
vwB7sqmOhgLSUUa3Ekvoxh6fKP02hFOc4fzkspyVe+vssPaSyqcNodB39RULSfR0
wEBrRq4HcgHXsUZI7Ar7mPeBgQ8iv67gegsnIMPymEbUMPTiOIdd0IhQkDgM3sOR
lFtYPIU/9WfvSTClaEZpjGqiBVfeCSzaQHPru+YxHDWMa0HrDCafuZ3EAKSjPdZe
qtSJ2vzzL22xpbVredbpG77Oh8BG/VIv3dpX+EhW4xYc1aqBTifeXJ7SnBnIoDfj
udw9gVYo5kEKYvFWZUV69HPoytK/bhQ1hhikjAdYxt1oS06jcBVjeD73xnL5J1t3
J4NCanbFU59UWgRsYYM9OLwWMG60OmQ98K5A2eZppZKkBHW2uCBXv4jNwtyAi5x3
rbzMEP5ytzTWmqKXMiCxiNUUE6FNrieeliiYEkmbrbQLfyhOUWUh6KfJ/CchyGK5
cqhAy2uUwqM1eb4FXNjo1bhqaQpHFjJ21WJDIOgcHTxsUDyoHdyQO9YbgFT4R1iN
9ad2E1ZtJtflRu1+LwbJPIwLgJIVeWdkosoITVCixcDbOfnO3JITSy4/WSbMToWS
5PC8fJ3uUS1IYB4SKjznH4VhYf6ROWhhoB1maQz6rJj8+fXiQ3qFHiGuEnj1zsuv
/bE5GDrFKP3tZ8YbLai3FmcTPPnqKazdgQ4nnugtsrYpeOo4c3juctIU94oPI22r
oQmLAWeGmBPXP3NiKaWY1fGvvPJDd/O4KMO2xMcvgUh0wk9fceEwJ8OVgSG6vj5Z
utK/XnKBSKJjyGXwemzUVE723EfZG+PmH4Y8eWwcM8NgTKQeHmufzlGnnTV6imks
mBE2Etrhh9gzu2n4j75SIGdWcKPeveOjYkMhrONNLc/spn+PPFH6S2/V7q1vMLWA
7GS6m+b6d7P9E4KUjQh68AnGIqM0totzAXzZuMT1KEvchj+2Tc3EeUzN9VD3vsx1
bUzAFjeuYHLKyHdV95ubw6GrQWnXKohSxUnlQdBuHdzEvkbyUTxAHegoM+c7JckU
bsh96JoiIhonFgE2tFuor0aPxyY54CpZZiHUk6zSDDi5/k/ulRqg0lIl8XK7ePE3
dUOOHWKfCsISKj02LaA48ABf3G9T7qEr/P9naOtc/u/JfOtZWD4Seba04WE2Je0E
o0rpD3PqIeSD6+bjicTKosDMdTAwLAb4TlPNEwxQnF+KV3MG5EszVN6/XVXFbcRr
J7jl9I9Ww/esbKnc/SLKL0cRr2TlNH7XNfD6+udOD3mAIyzIybv6raLE5y3teQNl
Finb+7yraSupzlJe70CeoxvLQocsKwc7KP9U/ZaSgZzI236dnoNb5uTr/t91aQkv
fCEERTvFVBu0NLXolwdHiWo/5+Q68ocgXbPpTmEvSwJlk8gHDX+FCmCuHHC01ycD
MGXJP2M0J/6X+2dWI+lszGXHh7eQWqV5DHgR7BaOuW2GGxl7Rbi7YjbsYKI2oAeH
D21HWAlFLGIWBxQJ+3cWnFhjukzplttZzgJDKVdnpCxU7VKv21VLmW8sZ9fqcGRJ
SxznoVQxMCug8goWVdZZtBQePTbm69byBhafY76k3Y9X6pet4MJThN8hGj2UgCbp
FHM3RBPt5BR3LIHmm7prdFlDYrg8SzGK+Ijm9W2awCNkE4XmUK21E+f2b4y4yOiF
nQAMsKCiGtpxyC+/Qc1zWf0qLTG8q+e9mXBZNWXD6PDElvu5LSDsr9fF9iDFN5AH
xQV093z8x0OtemDXuGKEWp5aC2p5zwnjah9QzWlKYnXd110rtCIEFXE41D8gm4IK
PPLW1mBCAJGMYnlvi0wkHgFEK28SdCOQ4szrtRZLAO3KmaahR1+niyU1U56JeAyE
kG4EQMbaJa0uzGe7re82AlTG+KmzcSxLNuzNdPbGuMElEF33RE8QuSDJfwGKMz0x
qiRk85DLJFMYLmD4dILGQ9RWZjCDMV92N9K5Y97BUHAXS3kTZoYqCDeCbr/Zy1tY
fj8c1RVJpZhZxXgE9UthI0Nz4nxA5owIyhx5sbJMadwUVwdFWm1WMHO6NEA8rRGX
tKsgCsjOsgUclsocBBBPKqqrD2OV4/KpDW/g6LDyxkdpFc7wYTLxo8n9N5WY8OtV
QZO+MPSnwWmKybOuIi583+HDbV4qNK2+FXfbkp2EMd5O/OTKqVBJhvr3bN9NOjMD
tm3kHGCBo/kvwYmYWZcfN+vpyTHD3tbLPGOtOutB8annatF9dFLE5Vy0aBnI5irA
VF3oCt18lqW3Z2gLBItJxeG9uAVIreSfP7mF+8ogjtRTWv67QjlkfB3j83VrfUsr
T91xwRNIHLRRAxZr83p/kYPBArtj4P/eq0Cer2ShTToViMEj8WkDmxA7SGLE82CU
b8dclUME2Fdo4gvpnh5Xg0/EBFjR9MLrXHaT5mDNxc0ugvh9HWnO3umUoJ3lLSse
tykZ4vRt7Ghb1Sw9BKlJW3kEhLULyeKO6KmMevWCzxwgcSB7gU3MDnJic5SkijZk
p7bxUJobeAu9yPuEhubNLkc4hYgzEa2eJROEvCeyzZNc7rKt6G5lARL/TbHt7BXZ
cqQqAhoYBH/w0ANJwb8mhOChaZ+vgJO0aleCY5UFr0mtn5hckzkqMd3hX8teZ/j8
5uZ5RkZgZB94o8vg7JLAadxPJ8V+aTp51FulLjJ1vj4J9GlipMAODiKIGJAk60D6
KV6a0DCu6rDgNfR3BSllTKKlAelDg7PIf+11woQYckZ2Zkwvgcz9wf3G9R09rxmD
0+nqBRmMKmD3fzdYLPLNX08qQZOClLjEv/JunjeYG9G3qioEDBCYCQ9sOUwRrgWf
YlO7KIfH4uAL4MSRggl/1sbyCmgQ+qZRz2x6Vbsf7b8hJj8FmCyT0/3e9WjgMn6q
2oFCFxZt80+G2bYFjMUFzF1U2zcjmWrTOn/XYIbS+gV/HpjtJa/dwOxkJ107v00C
b3nnW7h9tNGuga8S0Q/b6Ghi1CViee/3q6x1IIk2eNM+rSZHRuvIRqoAGj5RYSjG
n9gSE0X0Bvlh0cMv5D39IgttRYEqV7vBk2RmBALL47x3ccdQwkFawba2qmrnQfbO
sIG89dzeJRv+lYsR7EYP9bP5KUh4K2Y6oOgP4QJcJyAvtZT6+FUGbRlNsN5ZZxbK
O9QeBH2BAufso3BuyV8VRWfn8n2wuiz4EfIsFCOkK20eNTujvupAOeSWcFm+xjfK
kegl2RykWFyYiTRvE3+xOZQRlgMBdo9hn6+3FBLYzq5A2QVkzCrw9bM+FKyDTiYV
npB13cEww1hQ7Nz3zugWgxwHzjeQXCWQQsm+CDMxFYB28C6Gej4Ig4cbt1pSD+74
dCEMugmNZq7aZRdQZrmpPHsK8wRWQT6k8KWA+Zi+xCK73+2CdFLL54RKzonITVFW
IRqBisPXCv58Ujr9kYDWc1BtXJ7kNPpTQle05iLy1qLXoARbrDrbtCvmu4YOR3Ev
TMJaMVoVjiKsAOPqtVf0P65iW7bDyrnEPgkyHMx/TCS+RTai5P25nmmbZv6TOfmF
S2U4hjp4MLHg20MuNz+76RTQKhM+4IGDGbXnB7b/9O4F1Llwhutsam5ptBLKpviq
5IoCB3tKxnSyekcdboi2k+eDWT7ySg6vlBGgF7F2bkw93MiehqSYvMXGipCi1LBK
PDlSmguhI91zJAAeOmjAVBcrm/QupDRuePO1Vc0MP3+wXYOroC3MzDktGWTp7SIz
sGskMiMq9CXOcDMzUh/N39QSIDux5u7P1mPazg9+qK74uAQOQggb4Mz4/sZTPNeH
RiEN0puPi3jHZqF2j3V28eb4fb1Xu/9b7klwFbpTOfksTQ5KR1LsN9OZOmBBOEDW
0lzl6wj1FYWYA9xNzOsaa5MOx6ZJYw6SA7159FdlAzYhLGfjUzwLVdqVWUqnRlsW
kYbcclJ/P5Y0XakyY8m3FdtkcgOxjYPmuPcMj/rlrlVXRA5FgrcQC/GajQvLuWSh
duElkLAIL7qyiq+0KNawX07peXigSGnmf1MviMPfn4o7jTkHgDFX5debZS4OrfyT
3dtN6R4iIATCpvpZh7lsUdLaJYfvlGQpGr4lDZy95DNlAKjbltII2G0Pn8LeJESh
c6sQGYnYVhz5dYGk6ZahLA7vM6pOs1nhytzKgN/KR9zheR0FYg/oN+9oGhzQbpiU
grfXfWISJdElOCTfqEWB6huIbn9/t12XjKbdmt/Hv9EguBsc4fkDiSUcgwU3oCsI
KxpbYvcs0sPGdnW0OdCahPUABKchC35ApmEMVcF0SK7oERsQJyiBgmGD97NT5kQZ
Su4ER1vCKhRaTIRWdXvcFgnvAte4dyYiLR73pX0OONynTz84rXz9MagQuEtEsRfz
QOU/TGnqmrvxTf0s+HCEYuLPr1Ly6NlJ1ShD0aYem8889TznE82nopwriKNZr1v+
L7jPhJp+McCDXyUdUO5tQx9dDYeo1d2tRvbHE+Q0UNpkXH1H2SJ4Un42kq/VDAQF
AitPPVhEJWUmPlsLeZSuBxmi+92b9cLZypeux2gund+5OAxjhvuiqDcZgA1BikjR
/hGgKifK8sOfkjDAGOe3bHMrMrF7ktVx4rWiXwEdTqF5lveqi4+FFsLO0xTAWxxE
wSOFoCEjtKU6w7oe/Y/hjpZKu1trnjTylJsg8HsCA+GMEASLRIOmTIkQG7vmtZ8T
diJo6FAInfTfndkecal3sVyq6VsQXkTeXkI7g+9s2jmeU2Z5o5cB7+0olZQF3di0
7OTt9MCND/ngkL1vRYM18eKtPmmJrPcAcKZUiSJR3CKHE5XRjmuWYokThjNWDnQb
lDIMXmrVq/w2UrjQnFcu/ASVbXcQ+X79XlilsXbEfv9nZM8hj3WmOw5xbNiaek8Y
AuCM9vtnbLnuVZpITcFTOvw3RLbPMVQQPKTbK9wB//MmWCOG4DvJVEIZszh0o+ZL
+kg6gMoTxj+vbRhoC620y8I942yXmy3FE5D2LpGxhftRmFWkNICF+9T6Kqz+n07z
8dk+jDzub/gfE0XS0ulKvX+SZJ8zWihWHZ96c3ne35ObdEK2idP7ELJwqmHBjfL7
O5w0JHymLwO1rpg7779ocPrw6B/XaLuh1EMwe6esJuyjURORhm+NNfhiVvRoa58n
6awyD699gDd5/IFLXcPFXdTTepNK7sBbFWpMKu32Ai7kZjlrZdaKVH/nA2coEA/b
NDKiTwi9GJwKuVHkt+3gcRItwNOUr9/3VkWTRfnrVf/zpEhzpp65Z+FN3SQ7aFCU
ITpK0Bs2/rt/idx0ugJzMILcj4d8c0CSMl/vaWNHhINg2mqkF+llEhh/7nUwVsFQ
rfQ8qj1qGnFRq5+I/u8bKAtd8zrRe2vASBG8rbfcCiYWq5nHlIQJwKtK8nMv7fbp
sCqXwywAQzyQrISMHU6lQlWLrMb8ujh2J4d5Qjpxm2J5YMdbky7hQzhFmn+EFy7O
xNRLToNuEBdA+7aX07iMuB/7x3Qo0i51+dEbU5kKlwtd7gLVYCfepEStp9caGSM8
3EGPDSyd+kRS1v7jiE/hBbCHhsN22rLnV3yia6rRHKf6u6ei8130Q+D2E+A7t9Al
KJdamNTQtQ7YE+L/ED9/ZZawITm1r1BPERoYxdP3eGD6M5NC4JdQrkNzqe2E1bY9
+OT4ebpcqdmK/vx49iATA7P7toI/ULFel3fvM098X/25RfXL/j/d/8JapP8Z/ezz
c6z728uyBHMz7Hn92+S2btPIP15erWK4Ca1Jn7iFKpwLwesEsK1DbLtedddSuRB9
B9DcBXa2MK19wA5qO2NQ1bIittGtkeRgcVRuF2AJHGdNCxNtYATI1pPwDNbIQAGi
FYfgtWCy1zDp/PVedCA9My+yPqP6xP3OV1IMGZl7dxdM7ASTSJLquXnazlYuwL0h
d5tPDfoIrKZhgB+Jv4rGG+N28ZDT5zRBCmyADBkDw0wPtD8WQ1v5jP+QxN0lAoZn
XTplGWy5524W+Qe4UBHCSEs6ySEk4NZNf+WrBfFxuTIS6E+nm3Q3HDc80IChw0Nc
gVItrr+xP/Q6nW2lE0NwKF2jxSc5QVkd0OOuXUW5g4el0ozdrghqUJtbwibjrKAF
EE6Nd79v3A+/qNsLvojqVfMvJtWu6izTamNVO6VcjfH60X/b73AhQUNzNHJtiaPq
PD5C6FXsYZ58Kw390aewuzI0zLpgCshfjZbOUkd/oaIdhzn18H5dwQBM92avw8q0
v9m2t0s6EMATwEHCcyd9FrrPxs3xT7do1gQsAMMPPkNmID7FO4T9WGXKjYqsuj/B
2f8Ts9ooQDN4JoKPKu8MGTwQW3vVm3c2P76G9oVOZ1pUTTQ6iFyewRQzQQJtW+by
HGJd2eiIweo6SIHLQVINoiAJgfcYgtYn3d1ghxMy0JcnN+uMzMWAKzv56Twlz2Aj
fT5c0kfuy1FzbmWM/IOhhbVb89NjbcGijBBgs49LvTykpe5R/nB9/k/a0RP4WiWP
aZOopuDgd9MhNJt0VAGwzaSeqHfFGBc3XScRUpdHpW1IW6y3tH4qhyYe81r8eb9W
YtVXrWZ0XjM3uXsDvGx1Cqe6H9l5vmnPzCmHSKd7yxvVSaOaWXqr/KDbQau9LH20
kqbOQMwryBIDsy45VIVvkmM1XMOqAP3wrToNCAzSjm1NYfJMUiHtMsBYNS22PRQw
aAIsTMngbQ8Qq3tGUWjCnGmTQLCEwWNlwwT8GsvFr/CQxq7CIeKfeoDEHLQhrvsU
dKutNuXRqPcUaDRzXfF6CwjMavPmQB9il8OGOoS9zXN5aX5EWV0yxs9eTMTGxhnT
agUHdMlWRgZBHBhyoFlg5Yhb5SswEPi0rSC2qRAQKWkS4a0CoMZcMCuefY7d2n08
9XigVghGHmgrTBxbq1gVqta8O5MBMTY4uHLwJSFsEGNX59wnwub6EliNeCkqv8OT
sn0RjynkS4AA5o307NHhtpmk81bKewCRZAN6i+Tr7qsR/64o845qF8iBXn2izme+
UQojpl7Q30Sm6D+iusVsTQLrMw4sr8xQ4Yk7OnuOvFW17WGv7po8YeyYJWboxoPa
jTWZvkUILJTXgbd+2nHdhWO8QaRFKhCos/QsOhz3eg/xr8qMCZNzTBUD5GE4HF8y
QQKI9XBhfJ0QXNgWINJGuuUkyWGt9RqZrS/vfwm3+fHgdrNzjxkKxWBjQsaSCzH6
zwI121RXuPEyFZRSmPGQBDiBFjjBZekvFLN9xgSy1c39kZhd7hRNIPgOoeuUQhzS
8gi/GxfkKBhu6RV1i3L7xP2IfL5Ze+aQkjDoMtY/Rdb71ifdV96H06dDN3rr+3JE
7EVsF1T0Aqvbc3EoEqoKkg/ZOtIF9VyrbIXK+IXRLbyWi4jSsJ6qQ15zdrbp5uSn
Scg8XqVJbyVOhDyXGXieCeblkq5I+GqpwhyasiptJvQ+CoCya8MJUB1aA3ZinvCx
Fmd488DQUxT4Ae3PP5ffXbf8fDMf7BwzAMN8HMKkzUGAkHo/3RzympVrtewLmH+f
3uNOenFhBIQ6KjdOBVcYmVQR/l2n8ST1wZANNDkp6BGp/TztL2PlrOj/9M0BftFD
Dnn76WnSB44rXsGv6rzeatiHVOsRrvii6rTp+wzPfpBMos3yi4PVGPCuF5eg+c/Z
1VL6W9d+PDOEe1W1oda1vg7YcSxeV1loUyti7nBf2aW7TxTCSdFPVDm5pXVBrFdZ
Ef5Iv849FeZbf/rbK8KhrvSd/t4j5/sBs3qlSV6r06BU74v/WBMgJ3HLgl+r6low
Ai6o+yCxO2Chjy5ailljwKw3K/dqAv3BgzJGTGd2g/WILwU/kTNVfYkDIkrON5K9
NVCtVSryvgCti4EDhfH5JYbWF6NVnwVn+NpTYiRLZCoUtpwvLq//7uuQ4YRxMLZm
yK3tQPT2KYbcw3joUSeg9/kRIt2jIFBVw14Rin9wxA4xwZ/JObUr0DJqVTsbxpdP
6j2vpUGumt7t5rFrx422lshRR5uudjqE/6X+eK6/Tb4f2qVFX+8u0go6FFgVohFp
fliXvQflhLo/+QG2zxUsgEs/+RERsPpXCkTEyH5sVM4e+9qeGMTgbUm9bFSC4o9q
Zc+PdEUmDbsbEqBTOiGxjS0g32YKi55ZqGrlNO8qSuljS5fbZt8sKXO0qe9moDmr
WQ7KHJxztQJRprRrcWTMnXBBKANA87R2koDo6mGFEHHXoqZbSM87x1fMDRLJwj7y
0N3ofgGg/8zKeAyUIHqyBU18kKFALS6Qe5T+lyopKOrOw9Dvqfyx/SVETIxgv7M2
mI4z22UjbQlvBpv1wa1InALhTZpE6HtCKuh+1GzGePzxOy1rlR9x3NfORubv9q36
AQfgmkI4/T5SJFBN6r56KVrz5oye8RGS8sZ5Z9if3+i5IjpWwh4GS2uMDw7SOarK
zU01tu6CifciZBtp2GSwGg2ZQESbbYEhAisVE1XenWKz7NdCqs2otWtLSBycV8QY
++wCZLH3hqHjReF+HRfl0hicdLs451eZCWwjB19MCxsw9MDcCWkhtnvn6c/IYdR0
+uqI0o6eEZFAIHtpXeux6JPR4XORznLAx6NurqUQLjIXt4Z21bO2OrvdhANlqF4x
PjebQEj3vcCIzSBaS8rC7trNRGitxaf0gyWN8+CUHK3+Ui3LmsKYwXQdI3kpBh2e
9Ft8l2Qcw26Un50MA5SFdNV6h4okCX9NKXCtPzFPXKbK8ZjbGwkRqkdm8i28iF6O
KDX4rPPIisD1PX31bGuOY9qnLg+TrF3X+bU4lM074Yb+azpJZmB1RpHwA3cKgnIs
RdGHq6jskopWu3ZT17Q00phy4ApbZ8Rtmwtp9iwVTnvDQ/4Qq6z89VBmvHt8hWW/
cwzSYeibS87cYYlRVDCO+80/LSts2dR6o3UYvAz64bgqoanjj20FMkgPLF84LPs9
IrwnycHO3HzcxgwISJ69lLpGZCuXfXH4iqdCdxTaZaNM0JPEWRTbfXDX0OPW1FoP
deKnzRho5LYYjMhGtHpSZKNYAFAJjZfZCwbR5eOp+7fT4dQP36CqAVibfOrHnny6
2IKYFkiAvW9+BylEqRm7WVBQERJiuEsSbYpyDNQO+/UEFwWJfGoGWpbEQ8xmRTxV
08pCY6S+xS6tdY2RAZ+cqQug/MFuT5L0diIrxq6WA8l+aG5ScASY7vDiey7wZjnT
8FVy2LlQLM/1XQWncPScskpqongwmxBtkIVV8Dpu8dX+PvbirSMLxXxmX3hplY3V
ZusTneN3p3vn6RUKuw/6QqdkXhJX+FT5rIoXJ2IW8Ia9E5D/Vki5Wr791f30fQPz
et5ctws+21R0ad45VbKOrSd3tmkVwjNLdJxRO2WVIbsN52YtFX08PIVfD9dTaiEL
eKFQc9nQx5n61Das2jE5JfBXggg3g3CvJjSAuvy470fc48yFi1OT63u/adNggTDa
fLPScs1DamSx/Ivqk68m3dSKrhq7izs6JFF7drddJNtxMAA5VxQOjsF8d0Z8cmEY
/ywJch2ixkmgtiMeNOyN3aIh7WxRtV1yo7HOi/2ceV6GvuOMl7o6iQq7GjxCrmkC
fUgpY9ncI1ZHazD5lrE0NhwNyFk3/uEsnZzcitlhzHMP+1BWbUS8IEAZV+ikZgW7
ztNEMSCQd/SUbmcNBvz2f2mwCScwFdVsDIT1b2hVy+7fzHZLlRG29aBn2NFk8+xI
AcFdPn7APLoX1W1M4IIZJ9txpIranNLmNNVTKWkuE1AIGj6v04cRMuzwH44U/uMW
qsF5sGsOg4Jw+3G9Xx195NwO6jMWE4noLNYd2ICKZb48gjJQ1QCE62TEUIaGOr+x
lQVuPOT6nszbIDYDnoru5gM53T564MGMfZr4FVIvqgPsEpy+LQuE7ts1QxEoYkMW
VTq+D1bQejumgw3t7uuSbvFMXzdc8DBWyiYWB/xWPs18XEYDle9J+AyQFOOLnkOo
rE5DhP6m/VnBzeQJ/YsZP5tSHxP/k3267mW46Ql6IrHp4QbmOMroUihszWlwQ+b9
21XvTDmQUX/CpNedYin943JxuJ+HeZzdHvbalFwHZ984urj3hAyLfgEelhoa37Yy
cnAvDeXUGXjA0ze6fG0XyVfNflY+n9+gnOyfvgx8driIahQinQqm+2uIifrMi+Vv
R2fFzv64wnRTPghKtJIXnSs3p/ZKrQD/mh1+lUc7lmY+5IvB+OtPSEqaI99MEvjQ
6c9gQhOFjhSpn41ODmSQB2SiyQOp5McDwBOf9m4HczIBYC9eIBzvWNl9c7UdpXQ2
AEiUNeKqfgn1EEhdMS0Iws+ntiSZBudrhiMAvaMAPNq0F4wmIyDxHYG1cL+ZqRFh
JG1n900BFWyO6SQncTBhKbzJTegY9hoOwDtAMYEU1agZMqRP2p0D3nFB0ZObKaxp
xx2+z56p5tXdXezJJW7R+TUe33vBZWv3odHLYDB9R1AK8PTBmIwQE1d8K2dqW7ur
h57jdZOMkYzM/XQ8iV0UNJqoz1K/PNo6qGR3pewBt7Z8UTjvfTAq1lIL2VUgXGl4
loY830IOuHTf6ApbCYvdvk/XJBgrG/t4BWcW+/MCi0imfFsAV6pNTd9kdemgzqHE
tcXzB5jep/qqRv+lu6WlN/RDb1Q1OTmAmiDCHuhZdFs2ToMpVYhclI1qEoSzEvuz
B9S/bvszkTDLmR1vn+uO3Fl+5G+iVl2xZ6bdIfc5dpp21ZO3SXwUUSZZV82kqWEk
fn30Bbv5gwwLJHi+nmhy4JTHKJ6hqYODzagI8jFbJ9PKmcnOG41ro52VnKbNMG/J
VY29cqgwxwG/bqNrp20k38MxWlPS9l4xQJetXC290CN/R+dJcTabp2XZp6nOI4R2
G+Pyz4tCNznwmb7MlRRx945EzM7CmrC3KfDgk/+OvNmyCvla2quyDRqn4g5Wibdo
LR+rYsD5jQVJ9TyyMgD0QxqycLkhoy1DIshGngrTEfEDYSSngsgIgv7iegZ4jeTv
8TVo5fuhWeK/c2gPLKgGUP/NLqNtWQIyf3fmw131q7GKzaM/E3W5UyzM2wUDeDS4
bvjpoAPYqvzhN7qOTRE56O0OYYMuzdnSqsT8Z/zM0/PLP01ONE96KDlCajhhRisb
mGkrtdveFVC/9/G/4mpzS8Z2apTXozl2awZorfThlEoq2F5o+tCprOofpNlGv1Du
Z/3Mdhqvlee7826W6fsduesIAPnHNaRmB7Gk6+FyvoUaNGvW03YTR7j/MdD3hFSG
Gyo0jiiajTJyzNHZErKrBW6ht2tMdNqCvifJL1lbRrqU15qFWa6LUHxpDingsJLN
t5WRM/SX3UzXkWMZDG/0Q/dk2iNcG6xFy5vNm15jRfVtHG16azvqCZrVw4Y7uv5y
GZlUvEwyplqmhXSMZG+MhzIKFRcRUxpFVn2wyU4wDqBUzOc+UH8x7N61Haqb17Q9
emlZdEdK5yyRpNuiAeeYw6i+7UPe8w65fR8FcxVNO5vFA/tOz97oBl5U2IF6yYF4
3AdrB5UORK/nb1IgdlecH6Wy584JXgXYn0gNkvZLPnZEk8vyRZBPaDbL5lhpV8Zy
qZuFiCFGUYCR2CCL5SW6wUF7FnG6mbcbjaGkJlcIfipRkN+GBk50S5ZtJ1kR3yt2
7/HUiV1hDjbyZQYiSxIY/ZwIU8UDiz6opkeXppju+qQMoWiQty3UrIy1dXM6HG+f
iKDDQGbOk+PbNyE16XhdCW7L52xGTC4SPmGc800pHiW9N7lIT+Tm1S7k1yD4NL6N
sokVTawLssVJ1fz7VtaXYY7vTEv3XbZpiNVISMlgnwJApFQroBW19MqUfkwhidDo
UNlrizUvsLCxdXFrfEsB1jprgFh6r71hYPSb/UNRw66JW/WnLlAghstXFjGMeKed
u6CHvTcfvihzuV00cu2BkX7Lkf/lc9eHjVJQFlWuMNUYKu4IOppPImWMk9Wf9ZHr
cCHlE7RDTlWvOtqaYqE5XTeKi7I4mqpiH3CHz/2mUo8Cz8ahfY38kjLxe/qCgdOm
7FH+gHhnyN0YiPBntP4L2Aka6B5zae+Bq9azB6A64Q/UWacs8rl5KEt4/K04GYFM
RpsYwGOt5DpmQ0EZPbhRbB8zeUsHpPW6FEbTbSnms7TdtYFcuSZGSzujuATQF9p7
nZsKLidGjj3tsswXK6WCtyUfwAVlqFWop/WeXbcV1fVysw0ddQCv+jOwe7SpaIpD
ymY4yxR3S2e5Uhxio83TJTTgAL2iu8IwDz7uXTD6IOscZt92HJOCmbWBZqDcuxbq
GRqmVGWkBOYl9YRE9f7kCZdyRnmAjWEVq94A8846pPwjxZtc+KNJ2KYxhGE8Jahv
oWFUzDPfM+Di5/x37IT02sShzZa2SMC4l2VNE5ARvJvzJ3aJWPZrvKc1bJ0ZnVDj
w/jm4yuY8ScXYJrrgBb6RFqkNV7/tNt3rowYEANsfZzp/X7ytVYB8sig1POTD3yv
glKJ4J2POEdhaWtFpOlEJB0i79S9m4hyQMcR6ng+8vCfPc0V8gk71qiAVdbj7vLl
0mlr1BQ/kI7mhjx2CEf1292vnuSDXfoESBC0tGHS2z7x0WQN8yAg7SxleUu3T5b3
syEmsSP40G/fEsicw9HX0urMiWICjC/D53jY3CugaPOPRYff54bSBBJh6zD3bqsB
SfK2CSVMSrsU7+7Zdi6KrRg+vJq7vYIqzpD2I409DXHoTDqzZYQ0wdgvNIrCs5Je
4OXHhXq2kUvWfOrIGp7ZUcXN2QSPnxxtCnq+U5EJ34nai0JVsRHlSlXcwZJSaG41
KlzPg9Kl7bZFzLrpyKn3eWOS6G2rySODnUKZZ6W1G38pccx855J+5xEGTmUbx5Pi
KUNck+7T0ulYXoS7io8tpPWG0OfisA8GThARO/nvP87HMkPND5TUJO2Fvd+RrEmd
tnNFyVyvmHtArzKrleKQOPWLXqDITZDxm3U6Zsplm82FpjNvXAcarQuBe+OXyPWE
JA5Cmq9PRZr7k7WKby9PWe9YIwDl9Ln9DE76afidGhv/tkKtMzat+4XfWK9dEHtd
7EHG0HYi4aYxv46Q+MSvZD5CJhIe7lspWfJx4ChQs4NIgG6HuAHkMd3aWsgQ0Rvr
3iBq5R7gXXEt6jZiyIXxDeb3lwjkVzjq5+HYo0Mkiusc79VFs5Ygagy8w1jPCSNX
0rYrDnkGGX3VGWIaXVi+4kZYW9CyxTvbYHgfp7REerEsuonr+m3utIxT9QqQIUVb
mFUNWntykCBgimHyGBy+sg3wIm7SETqJNmGZ5/4g9DnH8hkboAlKU/at06Pmin4Q
Sm9XxH9poZ0MDaOb+esalhQd7ASsOruHwr5vVsapJiBKGluaF9pFK4SbwzyGxcBG
oZGmW215lLeHI2E47OPye4nKo4RALyIOvN3f9MkyWfhr6RwdDEJOp9yMxqwqtXlz
BTgb/rYf4cv6yDv+vaHWr8QL72K+dN0BOQGATbWnHzu11J3RRSdII8MiH8pb4zza
XohbeAIukc17/uafcZ1m78aGo7tSlIcKIfkkCCtI3aUm6ihs5u23dHSfanS2UFgn
RCbyn0kQ8YknrbYq/d2uTYHOVDtZj0D3xX/Pge5vU8HqqXXkcUuwAsrkJc/ijO3V
XIP9X/3u6h4J7th5RD0XLo0aJKq9IVtfVvodeCDF56lflox34ZJFVbA7tXBYwPPl
K9hcdO1X6dMPgAgXa7I8OC6uXtuNkMcYAOB+XzPz3UzjJkZXqGDJ/MgsJHZB/PG2
SV7QhqMFEhryu7GItj7cmVwAQOR4VgNuzFG2G8wrX0Ox87V0k5QVZ+0i3EOMOGXe
IMH8jQPV5ACI97uYjLqFJSx6JrEFNri9Fey1Woj0rM0FUKTluQ1WOQf1sDb4Lros
2smNiS3i3msPJTSmiR5OmJ9huzQSxDxepYGWKoTggIVoQ1JhWgd9xZrejOZBF3z3
3IimjKElJcLxNJ3LWQAlOTe0GcIlwWcJbHlNAPkokQa2k9mcLgZ7GB0Nn3XqOHwf
FXzxWP16GzY0jr/rADGI01YHga8krMR/TFFbzvdnYdvGz9Ny1EG/cEm2wjTsJhfU
F8am8OnkHZ7QtNKaUWGGOspeIioaQ8pPFl+QqvUG7l0CrWHUSOnZpeNI1E1U2o8a
l6EaOnpaSC5RIjsq7jIgSlOwvd9Raxgw7cVSge9An06XPgShL1jUl33PRzQBEQuq
idsbS2m55SGTiTwtj5VApgermXKoS7hms9cH58TbpQ0g6WXDorLPQT80qIERtYKP
H0S4OPg4uMDZvP0eZdnlsDeqeTXE3940FRDB0BYfONaVivf/pHsnvDFlLdkExhZ4
SOl4DfoCf9+A6ljGiMhS8XOomEDO7rL2Gsd9S+m2BguPuzn+VZ4M3/0XyWv4SE9i
BwzUiqxwORCIyGH33XorP4vlBwMRYtpaJTwqhwWAv7enyzmSt/laBTERmNaL/vMP
az46MS4rPrMW4uUdcGFbQp1U6YKcq0aWAZDYCJOu4ppFuwNbjJ4Aco38UJoNZxpQ
b5+NoO1xKLI8e+yqhmOldcpYBPJsut+ZLtYx7fowsHALQtJNo882wZ41xSg+xjwO
VpSrj3ouqfNNAixD0/oec3k3VwDAIzNqSS3hCU+8rSukapiFje2LVme0rg52G2aV
JRlqvoCA60S+fseL3ywFIM7ANpjXDNJH8531NLHjHyfUgj4OlpHPT7DwONBwewBt
XZtNT9Zy8P2INhO2O+kUMb+3cOOM6HT5juRIXl5yfaLU64rGrBTfsDcBDt5h34gU
ji+jCi9fK7G0UkNRLVJseKll8mR+zg1Svv7lIp5dPpLbxA7iAjkWWcsD/F3Dn2PR
7QP5V/eZxBlAtVYRbm0lmSMSC4j7ddvG0kCXqzC86ju02z2wkLOIk6hZ6eYzmPGL
dUX4UvKYhkmcYJdlfysjhGhTC9xMq7U+ZJ81wxiDyXBtxWKXPyihpklkz/hFlDo3
9JFdmWRs6MAFHpzu9ZHhPa646iGvWiayxDms3zfloUTq5QwCx5SDa7YcAEYcnYIR
BBxsca57PnAn8spwp44Fky4qf1g/AKFll6JzGs9b87cKv0re2EgsiREdk7KRqlpx
iYg+rhdeNpS03aiWJsB5H2wFqqwzweGdg7NmecKDImcF/d9qXpxynpZLQ64t3FaQ
Kn6KPnvFOOxAdf2x5V19gZIwIoRYOsXRnDerPtleI1rQJtm/QYgdXQ8D9SEChK/L
4M2qYoDCU04DZVxYyTfim1v/8wvYnB3Q7H4oDtbk0Jx2JTbSHX0MlDndXu9jDCzH
BmvRTwoDHcHaEXw74b529WurOxNfXFBOncM4EYssVJ70Di2uDCTBP0ds2s+HTZ3W
Hmyts53Mpy7EHDSD0IeejA8WBTg1P+SB5NcS42iMCC53TkTtxng8sEA3u1O+1vZ3
3R3au8tyk+XSwn/t6RNqguAxM7JiagH5oK1h0e1H0KnoOTGans9Lwgh2T7r4sjA7
PdeUSl7tQEn23fg3jH+HHZ+VfNWXv3g6cfRa93m7TITsx4DEbgE7z5FxZcOCTsun
e9KoigAt3GsUn0Uphu2f0JIa777r73OQPO4Qgc+fH7webNJZ06GNQ8aSVt23Wbes
9LWEWJ5SRejoeE7gBVq+MrLAegc2zMEOAOezsyrxQosbvxjmhbCazAaTSYGBm8vv
STcfhx9YpqEcQDCmTlz0/LuQGMTsu8IQRgG4wfTUwjf5r5QjWXZ87LaZKPRS82Wg
9xtaL17e/QJU2+dZ26Dj0BMr6pBw3ulFTDwZ0hoxFkcZodk7pxOmhyGYhBTE2uAG
/OQuvC8esyfJKHhpFn93jObhbGpDw/talXlvYmliKIyWPpMhh8YVML/7I8V4ZImN
NUggXLW5hHsaHfKi4pPXYPOcFBWY7NwkemOLAZbuoHS771Zr+8kUECNmm1YUhFwl
Qm5c88S0ohTCkrnal0iA6mHhfg0wfjdukTOufh/bmxD7xtVYiijk9foIyLuzjw6R
uS+rwKoFq/NqwPZcaJ7nzB5uTjxi7s6Jo85qIcof62yymneWaVX1Om+6nVJMNqEU
lcboljbLtrnmd6QYoAmrnikD7M47bKA+Qr0Xo3fG1H8jaIvYvwKv4iNbYrc55yj2
DJpxJgutmbnCRJSfzmJlbtTaCD1RUoXLvlqwI2EM9SsEQdr/ck6r0Kfg1T81FY/q
CiMoK996+X/9frGrHxrnLYC4r8IUs8seTz72Y/p4w9Yp8O87G51XJ4KA6UnLBcCh
M3ozf8z2U4bGmDRNlF/0T5hnE50YBy+hDfSwrfdLma9xmm3iO2gJVzlQwj2dQRl3
ChM8KyFLR9AgHiA0lWDmchBt+ngIKpvleIMo4V1JHp7sxGQqPnO6gCxDXOcA1lEF
A09AJZseOzSDT9tqUKpoYbcut3Qr0eebZb4bPz69cC6tCn8yUZiCSfUtSLWIExH0
7gusRO/IjcLkU5INYXXKTJizdFwvrBRATr0mxCd56q91gCi53CepLmehMkCnpRhZ
A6x/9eI1BOag9fp8ncNS/Oi/sZKemfd5jJY6RgRSpzXQZ7XwoGoiYVco+y8UNWe1
9iJ/69Ektw19rArb/m0OYnnfVpnoz1KyRS/+L5PT3BSvfORjwWNASdHw1dqdnuDN
CEOLrqde6MPm2uoQo9T0t/Ujkq7je8q/30wPKwNYCzYx1FOpr9vOjW33ZxLc8VPV
4k/W+989dLgA3sr3WLTmbi61g9HHd4iWSbKN8QTV+zDUFd3+bT7JAOko6O4IXosP
LAEASmoolVT1qNc8Z5cA2tdYa9vTOsmrMzVKA9TzRnrqB3H3xurd97eZBU8ehE4x
qXZIwQdn7SuVR6tXvwCLyKQR4OCF+wX72FvX5Ur0G+f4qXyToaoHS6HaHbzF8zip
5nNtfKndsFJnJatF7mbOb7tQwm/gnIqKjysPGS5bQldGJBXO8ykP+y90fDq4IggS
e/VvjbGkm5RI0OwDpMrsbVDOjr67j1o74vcz4xnJj6z1p2sRU1Z3TRLcWfnK/MhG
d/8HuIRYz2hzcf6dmjQ5vLGdpKCcc6y8wmm2gV85UJvrNAaFS+Q8zFtLig/41xeb
yjjxLxe+lNEMfOfhaWLbnbioBYK+l7pbedRG782338xhHMcciDFbCNYQ5ZbU/fxK
roo4WP4wJaV24D7HRlrQ7kjAolLpFv7e7scav+MAkKfmHZvO1b4VupAvUpZYhKQr
L1tzmpmvKRaCbJT5RRB4wLPngs1fZ/mEMQcmJeAd+gHF+x2kFN1yn4Zg9HEXr15+
r+hUaYncVmV/0nbM9DMw1EWcYydbDoEueTqQ61fYW3n+pR0hEY4Mb0U98zp0GWQO
aVKPYqxsiDVHN8FfwTUOPeJCzns+osAsdOja5LrQhD+QQLZFR0/LEDzgSstrELxG
Z3nVVM33N6Y99sgDrDBi793v4R9ZAsVG/FafdXYYzg737C/Au7/uksIdMzLWIqsu
1hzIdnQ0E6jZpXmPI0vIlsFtF53nwotiICJGvzI2F1oQ47sacYfutPxMV52jsObu
Qwga9onr8D8CpoY9d6W6p3qG60FkBnUZFQcwleiL6nCErWOAUboKClRREh7QeyYI
VcYys0YHJaLZ5eAIrhDgIZeLy7Slkx0GkOkS2RrpbYmnPV29lVc1mxm79bph5jXC
x+bia5E2uNzHoFRvnGMr3FAbEPOSk4/X4BlvsO5pCCAULHmdvqITs+vzB52YfDac
KDVFRq5/Es9gIeOsMEpQ+Fdc4j9fbZQmfl01rXXC802OEGD+6di/YZ4jbf1ZVlnI
I8/v5CglfstubiCtAi2zo3pb8bYM+BqDUHsVe9I6l3fuhGg6TFUAtHTWf508L9kv
5ZSWWjjy09Qu0On2TFF6MawmraXSzVc7MJpC7NCRGXR5vuHmdj+yLwvJVnEoU/f7
yFqZ6dqth8euIQJ23GJVyXJ3hc32f29jk2ic7/4+xuGL6K4an9FyhxAs5PfMRVCV
7I5rmNX5k+xTheZptrl5nM2XXqmZcevx1MOK65LXu8bEgfWtCInk/aTCOIPE+epj
hh/owMUkU9Zy//djxAjsHsknIycByVq4R1vmw3X3dj/pohTJtBbF85JecujsiV2R
8WwgeykKwkbSzW6c9U8ZpOqXAmLdr2X+nZGPggBnm/FLDnXZfS1fgbxWy7lPyIMT
7P/FUyQmIfLgxjAUhUwK8ubVFawu6DlcSwa25DQMPq09/n6PI3iuaX8KZZisGlIU
Ju3WyIk2MV6QPrpUMt263GEvq7EiegG+KSoG7BAsgEoNs8Y1hm4uWo/wnbPBL61I
BNDCAL7LV+05R46+hQa/b28yyxLlL+/aEpIe4gZSfdqDX4FTDSZs/4aCetmEZyOq
IFCVKtC5d2oP1qFHWr6wYKasFMXC4Z4GRYO3TNLA4esYEolMp9Kv6IPCnN5r6eEW
LuV0uJ4VbreVu2J8R5iBs0P14I0dfUugFMBWNAkv8XeZ8xCOOFbwmN1Yw4Y0hhjR
VT8qRnrh5Ai1OAizGYgVyx0jF2RYqUGmjxIg+pAGC1EC8dX/Jv4PHGzQ3dNhFpq5
c2TFqVQfPOXwAns5N9O8h2CSebelPZoZbtcDbR1LbwuzVAdXYd+ISDtsxjGcFzcz
UE8JppREk6b+lJRiC3YC3GMh9BF645wQan1TsWDdfoS+PDK+qngH7hzkJWzZFK82
RPD0LRLW7VEewM/Az9fvcamieArTrCE0Am4meCrgsupw1UnfoYJ3RACzbWYoGWaj
rswE9FJ0h0KQWPoyKBp5eed6zVSWxUSiY70+yVaIv0yFFynsCO9LTW2LEhzUhnB5
myw4//ntFKjr3C3V3yR5sEtm04xrTMPvhesTr5tUCsU0QmI/5eoeZS8W//fJ7eyJ
sORLEmBTjVRVAWcxd3QhGggzmFIf7N5CODHrW8cKvOOq9jLSNdnQXbC3hCqKywwt
yKp8iOKnf3/aIlpDsu0ZePRrEET4p5kDipHg/ZgYk6NpQ6olvjdJlP6t0BQoMaPx
yuG7/xFTy4aQ3b9J5lsIoKtXMEK7BN6T5kCbkb7yT5TdK8vIT9sdsqWUmhTAGXI5
Ddh345aZv5bveT7h2t5CJyWKa41P6Qq+UBLtxFvb+y5WjWplhDjsXjqOdTrrnMfY
r/4RM+9sQ/nuguRXeexS3UEmu0l8MC30CucLE63epDkLSqE9k7MWl0UVhTGwwxzl
I652mEQTGciKTyH3zHbO3WqzZ5uf2DMHCfnOl5r30zZMMyk2BkptJA1XQM8tMR+r
1V4W3UXjSsfrptWI7jIgLs9LXBFcORo79abdSypuPeUDiMusaVtyXLdSuzlaGvEu
gkO1pjkmr3ONIPnCXgT05coqlg8F8pOGcH0a2PnrqgRcC2Qt3WUd2u2OWV12DhXp
hkDggJOvjaTY15TgF7TRACT5zDbdKAvVWFwEbod00thJzDbxEWnTBZtDTrFOoizS
3LdY0RGwJj42vqjOAxeLa4eE2/7Wa62LqgPAl0YpEnIVi3PeWAMZKMDYR7y7JuBp
obyNjpM+4M8AsjALJKky94iIWgK+NFULyj0gm5XJWS1JgN6+GbnxFiRZX0Dh45WM
lC8apHV6G5aVsvyUNyOkoiXRx3O3Qj8CoEnpz72H+Z+iFu4xFFFtOdjzzp1GROSX
qL3WKCHzhxc+JqCksRtUhMnuY7ywqY+4Ba98AxhxOqh4KyaHfIKvoLBwCRbI/w2o
Yx4B8F56HOxDQYVAJk8PI8b2aYiIfqU9zLkLq88R+CHw7+TfHTl09lEWxa1RsBjq
ZULzGRpKN6UgiR5rVBUj+7w/X5/LaQS+GN1RNxcuvAQAPcqUi6+p/VbvSJo1144n
QvMOOHg64xmvTyHQp7jBA+AwKRyur41WNy2P7vLrr54EyMp0NRYgSvkZFvKmwD1c
9Xeo7/ByfXKMIqzepqLGA4j9GXAEs03sLJveVE73y3xIMUJF/eSAmf58USQMC8r+
kWi/hcpmhAFonRqBxYi/fL+O9s+I4iZN7HIKXGrncoi0u1pgccP+VbrcbIhcNfJh
j0w+zQunzx6M56ZhVvWC0jmyG8Qc07YOYM5V6CoazDzGSinHrwhmKllSF44w4bPC
CyL0zsj/cfwH7eOvuxcm2s4BOVyn1QgS/od1HLzLzAht/gsre/Gg5i+/jgM4oNng
gn28AW6TFVZBtqECcfn4Vz/x+d1gQFF4u/dpA5ZigUSCGxnlWi7lc0FA82kRJbmQ
+UcsLWLxT3rOBT7xj2d6CFPfaIhBBxETSeMWB0LrDPQp5idxPjAa8/uediDruO8I
XXeDipn6fTyiqvqpVAC36/svLCreQsakl7My7uHB7/ZWmgD1n/GoWJLQX10efjq0
mBjB4s9jEImFiYmS1J9BpUZTH0ZqSp5v2lvBv6LzxFbKtVOmYXqF3OnC/EFLGfme
AVAKkwdk8l57IR9wiztJ5nmLEN+8H7DsJt6ahhMckUSLcxha3K16COgimoCcRzFK
91bEM/ps1Hpf9WVShD+LR1BfTgW+yTeRPrxZ5RuBGw+Cv+jyLTYIxOelhVhzvLhM
BLkPbvXllwcSDMQKTcIbWtrgVUJJWxNPbKr4xPddTZFSJem5yx52fJFHUYzYqK6d
tGFd4+0eejB+EXSuTsTy/MKOPE61i7e2HGKXOJwvbzrheEYDNmESnAbneMuga1JD
KSGy/a1qjjsKrSntwny8ECt1mxU4oH8Krz6TbClt6dqjiVNiI8CT6aSSxfiPZ7X6
BOXgCmwqwPoolF0aSMUF3GeKeYaIGo/VNQQJ0rUUENuWm02jeyCQS93ofKrbBe7t
oW/VHoWlth9XBNTO+wdWtPQ/y8wKJROuZq7jST3U+STyUrtDWjqcSXfZuS/MQKaY
MadiErd53phJCAVzOmx1Vy1M1/nKQ4nFEP7quD6Ql6FhiorR6+lBgt7TQTRzVCnM
cpma255SOa87UM+TvO7LIjdrBr3Ew0M4uEtc90yfGgBzrpJejBdqS4fXfHfK/+0p
GDOWmdhQBTj+lAqsYkwaBFDPrsRh5C96Vgu81+cKzUHNj6J+32ToymRdSTBuEe0M
wasBRrrFEIHRpmMnMyHZd8rZ27xv36vTadR3RPj77in7gTCuTBbhsknwAZFCMElK
bIXxZL05qMvy9Qy6PSnAqTVE2yEK0cxHlSMEnc6UieE9WwYTjRmpo1pcFH0QiIOi
y8IG+ah9tir2ugbiP1nK1QaXieNeqWYXfQby5dsgzCm5U5XOFfcyjQmCSMrs759J
OgmYYxJjNzO4B84j/7R+VkAshzrEk5/5UfXbUQAt3l39YfOR7L0T3hqaYgiJLAmd
gn/i7nPT3QSdRYGq9VkZIHkU/NXtpZgZETH4XcqjPcK0aoEpyZWL7+i+XkoH+BUw
TEFUZ4pIzkfz8CJh2BVJescehD6zzSWt0fDDUF6sZsTEWTryqndAQjG4sZZLtjGw
KFiasfzoduWRmASQnCtcbPinIMxVdYSo1chgO/uoYdxKcQghNU9ymNZD//VYxU5i
oFJAnQ4qcd1MMAc1AKdXYgOAjmDh5It7Hztvsf9/r1a7L224F3ECYYuF450KJQ+n
TtCv8K9XnGNlL232TsE+BUsPKD41aZRshol7eywYxFk3ygBZxzdZRi6og88SZMgs
7yBj1hSLMlEJEfjY8Rqx4gAXvxlQW89/h/uMP4HsGlNZPo8Yxxzb5LnOYBgjhPz0
5qz/Sz19HYLtt7oZdUFaUXf0+dJQ0NPHbXtk1lDcUQjKVjdazyWtQZjqxxW2BtLE
vtOx+cm1a2fxOmwvOjR95autRYbqkmS2Ajgl2BhTqHJZGx9QDdytYZf7Dmv+4b90
5bt+LOFTmMU6TogW3oFlFo0PPud/bb93rk68IFWSOW+QAoHTO1X/rPmNHfRF+ReY
4L5ep1a8vIkMCS1yRSwoHW5LB/DQgzuZlDPisdhn+aAq8i5742DlHElmgunLCLPo
d24JFyJipaW+Xrmbf5PoSHtjPdfRItd03bJIFo2Cq7HKJY+mA4zxfAFJbT6AL3/6
MJTJ1evoY2VkeGblj5KIxyCDZ4wZ+IkzvI3HvyxDFpO6zTqDE9m75c8+hW29arq8
v3/MIhbYo7gLXX5TG6DIU+53JHy9W8Sn3O9P2QT3ajGRU0TiXnZ2jQAqHZQpj9Oc
qGIZVLTaXs7UFx3ixT3ps8NHBycuddyAjsKzNHtRu1eWPWHt/FBkk0SbhRjCJeE8
ReWGc28IpfvS0gmrRKSiHCKK1aEHB0Jgkqyu1TyJThaA4PF+wDK/t8iAXselTGKy
cJdBkPBMARos690evv76+EZea7rfMGkuA4uVUb+lU0PMKVrZOSH8OkYkDBIJW/DB
mDGAa0pcj06jCXImgHpux8YjvsBIYJGo9tLln8xWH1R8RCGzuhKqMJrFgKbyRc9Q
fvNA2/RX0eftso7wWeJKRGOy+yDhYZ927T3JKp4dhmYARI0O0TairmtbtRL7fW8G
z9im4xoMkRnxBANGJwbQu12UHtJQVuT7kR8Do+GSsIVVTeYIw+UNdY2twcm1hxe7
ye7ZptF/EtvH1DKBNkZAW7EoSqw2Gj9pKupQWtQpRidoXDfgOHSjmISjCdfdKMRS
jQeJkGYt0wnnqrxVPfVA6nPkv4DGizU/afAq8sAz8KY684vHpEuAetnl9NBfQA3F
2QdjuRYpD50ejl/8NN6CmoPYxB2AINUP2lQrDLb23mbvtCE5e2K2+QHgri1dv5Ih
U1gAzsismCGaf6NUcPURsjeZneTouUn4WR7aXjJxYKeqcbVVnXYQCOlHNj3Nvh2U
33wegdlvwMW5k/y52L8Y4F4ZdjQ2cF6XeWQjIKhG5T3nP1sLyvhN540t0jmxn5k4
0w/7eDq+nxe1dCcvW41j959kNVQimrgrqB3fKJR8rk7SmwA/wFx3Rt/+zUMMD5/3

`pragma protect end_protected
