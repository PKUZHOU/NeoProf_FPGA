// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
QyouH3JS01/K98MynRiaLpYz5e6E343vhC2rTPyC8LcanoVlWE9d5bNU2bKYaLZL
aeYoTLmX/pgMxDfhJ1DID5+qOnslDQzSIokh6LifQZTp3K/bS2dyMXgCC/crRLvU
TSUjS9FyIhReO91204tuh54mgetJDdByNpBssazg7VM=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 7824 )
`pragma protect data_block
3CwkNw2GrkwH/SaELG1s8/YxmKT8UeMGirGsfH1+ZLsRpZAeTNOr8Dgy/7Z03vBY
ey+neZJBJoExNPceT87p4N7hq0/7YUOyQN4EwDM3grKiPfpr2Ws/SlCCEyIKpURb
S1nZ1cS/LOPnEUM8uvRyLpz9k1zsx0PZZRiQfVycfhrR3vXfg3u1k1PDfqc1lhsy
aoNeWdx0c9IJZPelf0zJu23eoe3soYV67YDKLgs/G7bdeyZgQ6MAkLoHvpU4+qVx
jfF9LzJP1dw42yEXnf5oNi+cQ4a9xK5pj7LRUiJ/JPZTC9/Xk5guvxlKKljNzzqh
WnKfwM03kvu3N1J3p8AAU5txRztZkYLINDp4ZH7nAT022MFs+OQK9JPEgDOcnymA
qXN38wZNxa0oAyOwXOOzXk+YKpLeOn9taI13+mXfTeK0QsT47Oby25O+2dC+9njt
J6flexbnYVx6GZcvm/KsNeyWiSZ07hZjh4xkvsPEwZuO40DF6QVPhdthaZcD1NGn
oVCIdwm3hhpS7TslIagCIgUcvecObgxXfFNAcxd2xDZUl9IJql40rvhrzv/x6KRn
RrTAzNt4KCoiPsTL0/Dv/K7LFldvBmaM4W8X7DGm8FmL6ZcRhyXoAsDxxiY6i40U
SHq8tH3BMOGSpeer5AFuhUEFdNT5h9XhlfesPvMzUvy+HS2z3bYQStuS+rJWaQTd
ecQVFTsfC522WhOlWkK5BNy1M34mPQ4s8OT6xuN3lfbuZm0ic8nMLBGedL0sv5ri
UaonO3z5FY/Iy++gOFcvmjOrNVq9zgz87EWUmQH/3lV0qxoFxGVymiH3T3ePR/ob
6WsZsrtfTUoO/YUO55arwVAKtjCz3E0jMreqXHzDrapWIJg9/r0SJapMgBDPiq5D
7wfi+HFpMWSUYSu/u3Hw199A2vOZ/H1AlOvfLoVK4+IPR6rUvmDrTggoFBwyz8jZ
Uu8Tsa/q0jP5pI/gl/v1p0ZlCqL1w5ux5t/5Lw/iFLtGtnWyOz56Sp2HDP2z8/xW
HeyyU4a4o0u2phQ0jJDYH38x1fTz3vVyz65oNlcAo9WoyUC0Y3pLMwUt2BcFFk7b
wHAmhkedzcrP7XKfTZ0Cuc4hxVIMarwm9W1tN9Mqbxj6+ZwgOWzrAGcD59Dlo4o6
Bj0bsZzSU+B0vYAtzEPnGmPN0pkKA148hzKjzIMH0tQnT37fPKxrCHgjHIkko4wu
/7W+NbzaqxsmV0Vg22ABc5aDdcWO8DKPE8Hh7Aqrmgk6xanPLhAIOwCqJfyKUx/A
DEhorlvBsPB6jxjJ+lkDsmTCny6WcdJ+xqDjfRTGaeGhLaGUMaZvCj23r+Ju458D
F7hutmYz57t2u2qC8V0YfBCFcrJ7aE4ST3IOrTYj51nQ0ebBb+wLBmCfaGxhStOL
tpGW05aWR5FfbH9ZIHspMGvFkb2JIP8tIP/wj0+sMGMcLepyRf4nJCofuRJuHu/+
G+gI7vZ4Mri2X4KjsGmyRAKtRPABUsMunuld5nxlgW7X/+OKPvH+fScvSLkMdq0O
hQBPlbF4Hnzy0F4TCI8YHGA63a82RnovIwmQDgOncD9ZEbVY8BnLLEOyH9ueUpNo
AFW1x4WFiYrq6FxMw55X4g/vlo+xoLPgXcwzCnU6Vz/EO1/xwcDGhoSSPW3Sp0BN
rA8AgHSqGh/VBnJIWN4PZ2R6DGA0d14YydKur6hbbxjPeVX6PRIYxZ4wka8rLr96
55sUFaAtYA8ISZvgsgpbGV0YIz+1dk/S6YmcOA6wAoDeKYi9V/IBXdxGySzBpfU5
wMgqEdO5WprFmDa10fjHu031rjFvW7xFqQ+q4WSdg6tHKbRZ3wXDScZU2sBE8ljF
pTW+ODD5EoHPRNB8UQ6GQvoeaVrxvdkUruYdY1i2YMNeyAy5I3z0dsuIhmd7WQVB
nToL57R1r6NpnJcjHEtTGNzckHtlYk6gTGxJA7WE8/mHe8FJtzGOVN8IbBvP+C2R
ymaQBB2+4uGRm3gQkdPnFbkoyfBLB1rkG5wGwz9S3SJdLktdfHP2axZ6g9vuWnd4
sq/kkSgZ4SJ4gZy4tPBWXL1cOR55Sw6+ZWTaUAzYg5Zr5yxPko1F0+eKcsMaDdN5
CsOqAHIW0/0WXEPJU7K1eDvSvsgr5EfQBBR2PZhNXUNo5Hv+ALmOiVfnZjoq+rIl
VzAB30czGuX/EuiwDtgpwJ1IW2SCsak56y04S/ew6k/xUI5oYpM8TiJS/6lbgWjd
ASAmswr25nxWAKODS5VqKNVk1V4efLkBYSgyBSy3pLFYS3Alb3mhbWvT0W2Ch/fB
8IQ9c+PpDgYSlmRb0+iG8pB+Zay/oKakGVwdw211QFOforzNN0ZK9CxPKbAAxBQG
dSNUVGi+vOhoaK6LC5HERyDFn0rDlJLe1UN/YxgN/Bl5+dVnN3pWK1gyddG5VnVc
mzkYvDVs2+0dDp4SUWwXMXN2oJTP74Z2WUbG9UDO7VQLXTh7PWRkGLw3WxKd2Q8r
JvrnI+2FZBfj9BcvMI9yBOTw7hxWgKwJEaqCriFMqCOx6IbiTcwCeHZgbsfNO2XA
A/3yw15lus2lW/bHnTUOJKMci0fIP6Y9BLsTCK+tGruNBXomzDnmbwx9TCpPHWvi
l5EbwMShd56j/Muo+yUev319eXXiB0w9RhoOGPZfVue8HlChvFKclW4zK2EL7KEG
yKPtB5SFo0BPh8gj8Eq1FjhdXaKxsBJvU2ucXTzSgBA+zU2IzyUH5JC/BWEKK6pB
3D3VThFMnCKT80mLu9qaZOj3zdZ9qOOZwrxyl9jkF7aJYqqsV4134OFNnLR3NB9A
jdxJhqLgENdoO5LzehVvIUu5GWySZDtMvkulN3YfsRJx0f51mcM4JA9x82sJTuZU
/KXv0Vfk3zqbrzmnWocx/iETJfcLIwHWUr69Y1McG8MqnOBLRoQsku8Ah362YXS7
0/5QD1B7if7wBtwnCePKg7GCvGOc90zpHHLShxAtlE1Eodv8vQklT+xVhjCZ+yvG
CAaWODAvlJonVLw2rSUe8tOwTgGN1C7laEAkXVOLSU1UBdfzOZxEdZhBEj8kGnTp
2wxGih5EwKjCdH4JX8MYSX0ni2fx73NSFy5dgk+gEgvB/t26lOgN+EXGUKTY6hrQ
ub7zieXkwIWvH6JHQAI6z0YUL7r4SIrPE08mUcNyewVT8nHHRtax/hKtrLHAIXq/
0IPFBgKbzHZHrCAc77OKT5LamMhKWw96CX+aKAAjWohipCSck1tqSBhfvP2IemSs
9BExQD7OwERtknrLnwhklWalky7aH+xoXAkNjOSHkbYsmwj07f7eGcdeJsSwOAhN
8T7RUCy9FSaAs7m6wDIH2166ZI8lWVL992Shaf16V6rLowU9FZJuOE+flkhRWfii
Q6s0XnFsmBOb7zU2WHw9/KSZNWK+ghHLE9KgoPcTNRQbmYTQvzPG7NdOz3tLeXVj
ovJQbijHLkSASzQBOn3CR9h4P6VIelnUFwypXHBof+rSNnuc8uiQUvCHOG42EjdZ
YodZnG4Yju7AcYOJX2lxrjoH+PBtPWPF0HmL1d9DjmTdkWu3Cti6kKmmdwF/e1R4
mpkyhaQj3P4sRuOn00uVfNJ9A8ZZ2Dyg6GmKi3ASqmyi/lJbTLOZ8qgLfnI2I7dS
eewdwNb+m9Db+82xxHHtuMVj8mrwp2Cwk2EuG+30bOJ4nFUIp7u9HgEigI9J+yJI
NrBKQz1AJm46ssd0Dz1/XBdQc0IqH1ijgIW2uK98LkdVPfEp0vzOfxXUjCvUMGY7
edw01ReiBPBo86q3rsyIbxoHvTSNH0OsKtmBjYshnJ6c4FyDB1PgbjR8Gr8sc4mM
vY9SiZ+bcUq7KE2yPRGVNeEtEXB17sN8qv+8t5ZaSnrGQH1MwTJ7wCnNgL6DVnCC
kZU+F0Fu3Xga4aC4/SgMscLZPCGQavoJARuu3iphZHD2K8P5TJ9DuR6ypXmZRm9Z
Ad+P7F0Ol0zqeMsbXOicNtckrhUtD3cdd9RCFxl/wn1ak48hbF8sOUiTaRoF5z1v
0bdbqAPGA+CHPE6U2v5a0YqU2rZitL+XR7hCfs/+fNWyp/c07mgZ9REBkzP6T+zO
wEXlOMVGiSzNzz+GkqWZTqflL81r/AH/T9gBfhYy83KL+4b5Nip2lj42J6OPSeTB
vJTTepaCnpySMf08W3tLyQeORBBeay17B78JazPYh/Avr48xCZMSSO3UEX12rpHf
yYoVdtYWREL9rDNdcA66qVYhoRYzrstVtY/e+4f7bBgNyEcDfpDy8RFXa7Xbr2lo
/nrdV9klD5EjH00rEUiaT+6b/MnhwbZP3+EEAyLxKzMGt9lYan9TvjaR2eD4MUrP
lPiMHR01Uu+czKhCleJBDK2HqzEyk0QwwC2NBoMFwdDa7SYqPORoiJ/SnlH7gqMM
oSHOj18FtPDOu5kNKEC9J2WEhfGcL7rvuThIVcl7PsP80yVARZyJX3RLpUYRNa4t
fyVHg4XrAjdSDpyYeZBBXuXkT8ObNJTiS8+gY8KhQG0dvVtJbsMU7z4qDPHcLara
BskDcSbDk93W5pF93UviKZU7/zn6jIGYK5/LUsnW+64kX+vz6bJwi+WFVvYnFWko
SwWfwOnLyQ3BTp/OUiFy5vFmbaupxTaa6tFTBfAwo9iXDXTIXCKnH3ejZrDMoNh7
Eld/z2btddie3L1gwiLgxNb0BpFKD5oo5pHhY5lc16z+vf2kz+MkLn27pGGAfhOK
Z6452nzhdRoZpLaJMHnLWHGPW8Hpm1fNvFmdMRM3UHg5p3dbVQNDQcrM22uBo4te
ym0FAk9/gk0cAgRtyV2NkvvLpvNf0tLLMwwIX+VhtlJDH42dNGmStqSCLY2P8pKQ
KGATilPOiJ5uifG+F9/GldhM7Uhkn0QlqwLeEZe8u2F9VSdUlPKepM7M0MQ65VTL
LensAyMGOrvMo56agTKre8N+AgfXmezsH5MUHGtB1ek3X+5qU6CHjygN7pGiWZI2
pfV/y6+apNnPjQH1AgA8LomTiTwBg5g/SD5h8sZzEDEBQK7Sg9ojcO26ExiFT0FN
W7v1tR1AQBdzaAGB5lw0Ct07r4Qb9O0HsorQj6pWEIK6+49TkfdlH7v1/CxlTQfu
BHVsWo1NfNuNobJluvgEbvWyhkfhchmg3leKd9z8NkZvqdnWkLweNmyBd3gVVGbj
YI1ZVXUGTV7VXzr64XWoijcux/zP1McIMONXclpENuxAaFEoRrrBqzdkJc7eaTQ5
/9drWYqvg8n5Q1kI/npcMZPYvNJhRAEcJjTXwpc8ONORS66lVhFVvw5uUj4pUiJZ
e0+AMtqdRJPiWff8ZLM4IQM06QbxPtxZri6vBVYgu+CUrUQjiMXeHLXdn2GwhYQO
jU74lQZzwnl4XVLZ0b9LlRvav9iSOMApq7gnNvAj9pElJ+UKn+om+QcM29cILa2D
i0YuNP26ik7g/J9Y92FVjlUckTgB4FcA+UG0d5vvS5ujLbwnMTugLijzYWJMXjxD
mknXcCpXdJO1bTho1c4K6afu9pu+j59Bg4y9uZc0o9MR+drpa5ksOGGHQh8Ir9D2
X1LjBwcSAy5PfWyVeLtCmFb9/TljdVItL1Giuq1DGylWkuCn/qyOrTVkx1S4MRa2
xnnbpgsPEJuFmYDV7+ZNBF+19bETpI4BgxIIKd+p5NEijijDhWoan3dgGbPUoIVT
sLmBDDDnraproYwoi7xUhAPdZwuO4j7F4sTP95OD++AEgh2fwChfwMXKaI1Zp8eG
MYjHjiVIc11/dEGv3dzI6jXtaaqxqwpQOtDm0reQ5nyFe/KxUtBtVdXbbkPdwrPu
WLPcLyUcL/jNvbl79dJqk+EsdDLh1RYrY0uiTMmVoxyhtdixxaPMssig3ElCfcy/
JmFn6FEri7FFYHgX2qd6uN2I1AO2S79Xgy5QkShjz9QS/F+/zmQnEBQ9s96C7YLV
ZLSaMAvpyj1jPe7KvY+PhTx0JGXKJCqXOLwMQTIJth6oK3lMVwwE2I+t1ia++4sN
biXBUisfkCIUZ3PxcgRun4iHrnQDspyWEfwj1cj+2uxNiRsufc+1qdq3S5JYUPDT
J3vmhy+7+bFbZOmMf4AD+SJM0kXGgwoI+HJ9C0j2wRstDTiQ+q0MhVOvQ3fPO+Px
EC6bYyfsJYI32dWkq9LBhYI61V/IAcgfVc1wnNnrV2evhB9sCqp+xWObsSnAKB4T
2yewP4ZPLU/4XA3AdYPHM86W0fna2iutAFmI52JPuzect0UK6S1LFIsg6wBbPI/H
pi6Cl00Pt9pK01DW5sPrzGDcOrFeamaOevv4h3Ml9fL3uUpYGDTvXxLu1vaC/1L6
+ZW4HAlox4iDcHEwvLBRQ8gV0L0VaPo/KQlxS642SByWSCztCTxMpFYsbcRI0yAR
ZHOJ3EFYsoJn3UJyaudSRLz5GVBOHHUfULkg/qqoZnQlUDHxS/xl7LMh2yTfebXc
0UjDjISlJTEos84Q+DqI8BV84OLGbFvo+TeDor5R9RPGOwkUtTQuCn2T0yo+XXcQ
fIFEUwz9NHjA25vnDxNPTpjoaKC1GN8qapRreIsck0XBNyTd6+fukNvaZGdqgB/M
GEthderrvH/ZvfaOMmrvjiEi5QAmjt8dvNZ0XAOJZQgQLjUVbTj0Y/2YlHVB1qwG
GFr+7ekKzKmCoqeedMJFy4OPCBhkAzXqhjev/FSXdZSJhxZAWLgUV5UVyXWKizkR
V+zxa4MSEjUQaGuBvQfk1D2eBO2Br/sjpCqyGRj8rYzvQsx5H5BCpci0AIl7Rf3Z
Z6vWDsIF0xNmuBE7Zh+/xldkFH4Ng/pOnrKv7jwD76UuQ2IuX1cwyY6YmK5pUXFq
IyVnnw80HTOXups4zaxFLSwcTBfU0HTOcub1XZk6wcldaQmaQMU94Qo+PMLjuNuV
DVQ5A41AA9lpp1U7ik18k1aw7HABEqJKR+jAsvwOpnVIR4q5JEraPV6yZ2oQK7tz
+bvVVtWbHDdqgM6/JKDFpPiszY6VGBHwWuOZbGdkABOuOeXcRpbri8qlECj5qRAx
x7P03EnVW//c6QUIDeLI/t0/FyPst9cmbxxuNPLm8xK934HyU/1DgMeLcYTeuMGL
Ps0cMPXwDMQB6rTq2oU2d1XUtx6i3Rx3JPePu0zB1xlEnCu0mVfZawcYGvAGqjGv
6f3ESEP1vu0QYHCGxWqXBdlXIxfzZxgZVL6eUNFvTURXlhcR2VAWusONoaFY3YLj
t8Cv4mgFLMULp+6u4k1JqJM4fj4HlAaFHmsmFTDdQdM3lPUI50IVtnDC1A/hFQDs
zbagHf0SMmM4tMjjWHracpaylEKzQ8YyvvwbXX941YE7zVLlnwPj3tyYLldfDcRv
z9NNeEBWyJ48BWs7bb77wL7n1QF9lbB2DNZhUZtxCSbPCzEWQ3fuPKhdTZWuoR8+
h4ZIhwFHxAKpAUzTrSZ0i0K/lANfXlQQpIVGW9oi4mLww0ZbXkZbKh2t57oHv1Rn
ql1L8qmsy6et9tCtp5enwbd73+jLpLV4VBN7GEAtUPLkJDChm3gLdv5mK35Mh363
V0jaN8XM+TXdcVq2T73DMG7uKeXVL3Z255dP1j+EXbO9bx3b24qHIW14soKfofs9
h8+/xEtS+WKbui2Gz+UOX6ucM7QNTkBGzvBjvc0RAk0pKcx6f1dJG487KE8AfRR8
EdOG7wTS198CPmMLldPLIcjQRbdfjqHjHlJjvLdwbBIc6h4Bjf2TsHOCEGVF0XzL
s26BhU6yDESMqQ4CpAM2zxu9/CA0FrLjJG7bkYK9+AhJDXs9+XqKisICLkZ+1K4+
+zr0hWMTP1Hj9Xte8XPpwYofyO4zhBr4I9UZpptMCtLI4rMGYGWJE3OUVpwRGIZW
nKWvqsrEx9lNT4Isw35D9Cta5cilVAWkTYq8mrQ9ZBaNUI/nTcG62fAnjHZ4Xme1
7iHxEeXRp8xalLFQuO86/yGOReC6c6+LMHSH7mCSOepBib5z+/6nFGYH7QK+Q+ju
uNoFyGNq4aBzSrJBKOIkrg5oAtFo9PFE3frCWLm6bSp0RhCMd/KbsdtHbEurVXkq
03occf1Mc8rhOnQlXpG0UPcpx3XwY3151BjfhT+iKqOmTUPKjcrhbLFQqm9cwJDb
Eur16JQtKOGrLowd3n7Vo408Q0/AaxW/JgLY23rrV3+xMb5qmZWksXZ5kdckaIfv
rzdlBa4tZRknjr0J7urzlGK10AhjFyhbDl8+d8Ymk9qpNO2jhWka5ckanClNcZWj
fbwlp1wKucsT+RVpkAdzGE/ubwJvhcMW7dURaF6fTVcoomFeQeAaBzJj4NSVmo72
wxng4nSHB7YgjIg3AGIO7TLPVgMbhVngYiaqUOOmwT/lGWTfjlXr3B6Qr/8a/9Kx
xL4c6IMuSlzURLsv9TZz5lWgSDyrh8as/VV0glJKjjVW0I5zvlHib+oj1dygzvjU
vXwsqwtcne4KPARvRiQ8t97VFEgf0XvtlQfnQ5Im7r9o7JTZRbk8i04QgTzfSQtp
OuNG3DtixCeXDR8iDajrmJcvUKrozvMxqbQgU+e7+flSLfHPDT+hcP77njF0xt5/
iWSTbjPlj2NKJoy2jNksHbmDJxhIj8+1w53r4cwmnr0GkjuKA+zSZOIrThbdyqhr
swsWmgMMS20Hsur/CUmcAjEhUpbawKZEj9Gtpymq6kcxbP6tgOKzz0Lnw2V4TI++
Vg306sWvU4Eq1oqhU3t9i76lD45WID75JL1xuJodCj/sbnocxveu55PTX/oacGVS
BLy+EmkeO3tLZegHvaC4J73WvpyR8SfHf+KAUpEmSDW4uws3q7SIOXDMEMUw19br
qoBVFfbYFvSSlNEfiAR2Pml3UD+j+gdZJjwGNDJ9rMJeXf76IW+HUHD5eDRu2G77
VAFBLtzBAI++rMXwWTQv/wqyhmfyKG4kRWKvmVyp9a8DjvXvC+2yvJYzooN7ID1A
s0Z+PvbkLm+CjGWF74X83jC+xykTysT6Yf5DMnu0n+JdWG5NtMWG6CIIapAApZ+r
9Vurbex0V/nAe8ywapycC3WzyNtTo3WN/y9eMLCsZHtF9wy545uAh1dEVEbLyb4d
5roXlhIm4yzUrV4w7FGYpUEJIX+vT8daNLWEH9nRMetAoyvjYnvGvJCSGRNmONjj
8se+P9aZZvnGpBrKlGLj4aLIq+E0O4huRS+NYCO3BL/6F9PttQYfWYqJDIHhCell
FXkffAGjSrddhcIyS/AxxA3gL8wrDi6WbIlyAeLoYIkgAUvGM/d9BKjD1WoiFXse
JkI1bm0KvOn7pPlVK42qSNC6uPJyT9Z1bfHKqqPUbtt/UW3GWLi42sKKKKZ9O8VJ
7Vs2Ncph1We2JsuxQRAz47/rRnYTRbeeTXAHgaXoiop7+WPhfXzhZUBrUpwphofJ
pXXixjelN+qDPAFTErEKVSfGhniaRy7GihPQIwYqdbV0UJ1J+hz/Ep4abOWmifZg
5PkHJgKfLUb5S84icrGIz9skNMf8L/fuYMz8/IeNn6wRKjhisJVFfYpsuc9kkp04
956tPvfXGYs0NSP9Ku6MmqwGej6ZAs3Jod1me2OLQ0wn4kIFCzEL+s1NbcNluYK7
LnHvD9qbcDAY2LUBIyRpMnhL/vCpj1OJ8AE+9/RStDXTvbFucUy47BdUjXHq9lA9
KKKYLLGRjolxsiH9KWRls/L8oxKdveNyxHjfiPeSixO/XAgxTnCWZRiNP7tbF1cA
4jYQyGduwBYUpuJPmHX0+azzalBSAIteHp5NJgYTbnVlXJbD74SX09NIHyYqAywR
Q3xhJQWHTFep8y0561VdotnqAxySR6xyubnNk/TXsThsJHwuvcKtn/xF8U69jDr6
6Dl68DHg7LUJNiViqp4tKHnQY36VZ0EwAkwnFQPRiwBfzvqwLupu9g4/Ej684OQ/
3Xo6Xxm/O1tPVzd9n2sw12ks2XXQWPlUeLAEfUXRR+dmBt2oF6nMRJw83VtLujNi
TarNO9ibh2X/gS829r06Q6KCWVU8plTNPDwKP22TJDS8OvSpNYm+il/oT13mJMDk
trjWe+/+dyK1Oa73KQpcHM29RQ95feSGoYTBdmKgRPZhK38G+nMJHj6CbO/8QUGH
qHF+k3VRdU9HV10IaaBKmwwSrKLQjzeE4Qr8bRMP0MC/WILp1EJIPFWiaTveWZoa
vhbiWXVokMNo7c1vIrnmvIB92pM7D+gNyCcB8sBIC2pWJnd8rwdCiVsn90mS3/vQ
peTK3vCqRSd6QS3iFjZXv3J/Dj7STgSfzqoAnkNlzhHfAgL2iG/VdC6dSK63tzzq
tHnXn9ZXgJ1zPRot4gbQOzog9i6yQGM7b5/1D71dvrUR4/Nk493A99vSxNHJ+gLW
pk+M8NQCb4Qf4u46G7GfvMTrgS7rgPeChy9Ve7BjpTtFsTX4ha40fXcGunqhcvwn

`pragma protect end_protected
