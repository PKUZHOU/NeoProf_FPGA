// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
dTLfWMLnhycp5cTqZwNw4LpHL9ckeFuRo2qWfAJHuJOp8mKQPqruEJNXn5mtTVqY
CD1pOdXeHBtHOPHJ3pJr+wGrhzzG6x0DgxuWFor1rn9SX4RMYQKgHXrcP3H5/Jgv
lsQ7wOKUsO+RGTZ9+FWJW0hDPZETKjqV7zJC5rYjX6s=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 417936 )
`pragma protect data_block
SxpJFENjiWQWRzoj3+2M2U0Lz9/cEFPa76dvEb07CG3m5dvQh2yNkQko4KvYEQ7l
2h9g4mkg2JF0/2iBiYyRcUwOI8lbwp6jTfrSsXdB63xvXFvyaXaq6vjGRY6xMSfP
OpfX1nsU8w+L3VPaPwQQdet0EW+6toyV/z5RgWR0yByo4NJoW/0LYPtuvhiCu1Nz
psgriJNQocSA+u68tnQJoU2+7fZTrboVygjuXjOU8FERIGFwqeLnOOtBn9Hp2pce
SUFegUpwDlD3YCzvzSDfPlpB+i06+FaTx07AQENEW/74HtGo1aEJgI0QFH21hb9J
JGA0meEPbsltqzoOBlth3X4QyaFyI5VlHep8UGOA9+sK7uqOUimpzJ/iUpFyOtkK
pwbFZL8LXS6l8/NZv31Rw76FTX9iKrhmfdUAoDtb/blCrUG1htLeFdDS9mZCj2tk
6E1MUJEji5xoLt8oMrB+1xynZGt/jtseMYwqTerNvE5gAhX9NEyDp645OTYR2YrR
HaGzCJXuwhryUs9/WGhuEBXoe1VuPXqViwRwa+iriLpaeNl24E3pwDBQficTIphY
bm/vwDLSkrLZcZmILdluWq7ZARJiy25kAT9GGQpt7QRt5ATm0Bv9SlaaSB1cnnzu
7zTwAqbLH5C8Z2bprIsRh9RX4USjSoe7FVeXWh5wlaPug6fstWeA0t76fKuYQorK
miD0dFFjkhhwHe7S0K1pxpExYE15h0fi0l7XYLR5PZVZVhZ5OfOo12pkPzNPXXo3
40K37dgzdR64lC5xjsob/hUjhufzF7G1JjCT0XLBjEKaleTdjlqZaFdQ7YeuuflU
4aFgVxQDM+rGCn/+jLZXPnA6c/D5Q/ixnF+SIOLx6Vol9F6Z7VpNpZJ4G+S2VhHI
DIvk9QSxnN6E35VtUktf9oP/Z90QvW/Edu7prMo5SeI2EhoaYV8mfp4gCtSDErJE
PKG/pCHADBh73zZAr9BwhiThk5q8Z98gBbRQZYvHCBU5ChTrSajnIibI0Ej+sDnY
/YSadnureasMFZuT7qNnNka7otFL5lN+fS7n6z+EUkYWhznR1xTYkG75exGwqkXQ
x/jwVqnItzmcCuJBZ0wtNwBG36MPVTXt3tGUj6QIIizVj23+teNtSRKEwyw7Z4dy
TEOtNLCsavIuuuMWaJJg09bksmc8lDB5ctrSOUl8sQHVt7C0y2U0Fr4V6BEjWp97
zVQ6cDU94o7E3vYZtlDiFFK9VIfrD7sQpkXa5nBlqKYLd3H+vn84S+lblOG6p1tG
epKl14nC2RkCVPUcBESrFN5JMGsMA3OMvXgIjNOJ8+4Admiybam9mWa0t92Jceq6
ZtnRZQ3zys7qO6Zr2r+VOcjdqTf0KcOceEHOVqjxfVb316jwCf7PBqQG5APShlAP
CjWoh26SFA8y3wvls7CNn8udTMztudYIrb83ZAy8iJyKvAWCHvRBgPogtG4bkCbm
t+FbDAXfkidQmG5vLnpoSIMaw0nJ0gXYDVckrmA2JKk+MeRbaTp0146SOJF5dnop
g57Po1Qm0fq2YS46O8CXnogMBoX2V5YbKQ7IkeoqSbtXYq84KWQLJyI3s4I+5vdu
uS0MSmgfzIMrALxMIaXmZrQZzPPTZdqn6WtmuOlr5Xy01URusw567ji0IceQI+mV
KT5Ydxf2ssS6Lz9NSQKMv2+LKhnbG3CmdR8fZk4ohrlrS/Gh2NH4WsfBISxYysXs
v9DhbL9cydvGDQTl63CXyPlPyf/kqktLuLIbIw4HGHvkl69zsJBjhiJeRH9ewb0q
woeIgn55bfFTq2CDO4n4Lv+Th9mFIF+HnBeAzeikBuiS4addkmal7uTdfmBy7QND
Lp/yYDP+4ABTjPQMlC0qD2oi8UsftB1MKVNNKaO0m4EAr9QoK1+/K8Mm9Zg6OUwj
IlsLRCe/m0hB5LzuV+zs+PtM6gQU0iaPLDQTI3nusbi3rTt++VsmImScwwwIIb2x
0lxgPSl3E64k75VC0g1xFcS+elVfkAiasLtffwae6u9dZm8INA/SNpbq+mDvff3w
FH4xb8IQJMt+LNXXEqaQXRBijFzZQ0GHxM/ty6+XIKHQIKeEj42T6Z1y3mrJ+hBa
iSxstZD7c0to5A5W5taYw1bhX+nrUSLEwMPbOB6xoYQflR1aT9dnpi1DZw1QLRuN
EoXFc6/h8A2YeSfCsTqUxr1mVkTNfn4WmYCoSVu8yEAEArGrnXhir8rzO5hskmqX
99ifECDry87Q8XsOSoqOz5yT85flwL4v0UoJJP8u1dmesBFiDCHwhKKbGkUcPVMR
f6kuTGWjfEIH/P4KlEf5GMf1qlqjDXhjRaNBsWoDkl6+/yIXgoMbGZf9DJ6KaK3u
v9f7FABDECGmflgvXkCokO1YY4IQke7uu4JflU4cpdInN+xGr7FZ0Ir5Hxi5SOKj
3AoOhtiEYDt8HN/wyLgmY1/e78G7LBeZYNQZvJVq1i4v4H6eRIgeNBp425Ma9kAb
AGMHlVtJYo3pB1naP3PcSdThAik2uZN3878mXdkxIQP1p0Erh5Ry2zazkZ1QkLzx
0ma6rGrsrACi/ojqRzRGORpzXbFJ7bw/e8t5HAWTaeRqdMrjP7ml9lzBwsfddDzC
PoIYMokB0suI+F25gb2Smci5pww3pbqfda5JsEcUlwxrtALi37/++pzaoBWmZhFv
6YyMAV0T2Xr6R9Av0aVZqkAIF6yCtS6wMl/61O0skDeT6YNbvU2f7hJuWqygkFkG
RnHh+cRPXrEdFhSoScCnOmvedccJnHqIB0i/BPuPFB7UQvbe5VhhBS9JFWNVI/i3
HfsHtjFip9u4n7o/3bINQ9Zfz1pKyX76S0brPpGdaapYZhZsTcC/OLTopaC31rsN
5jZKhwHMy91Vhv82dKW6lUELlllafzVvOiwQvKQ6vdvNziGtI+N6fixK/RL1K/bz
ecFzkAAB/IhK/M1MCwlgIvf3I90AHq9xAhx92ET0isG+DFCx7SRLoPoZ/XM76QAN
i723YF1n69ZxNAAhqxVyqwJtrh+LYmHTzf9s1j1OOwku7iristnaM1/4vh32mwuY
kxsrdxUp8inE5xFTWHP9Ex6rN1PkUWWW5zANxVBrphwfZFGl1p1mdfFzSAe1cnzA
N/CbrIU21N3hxs/PRvs0jDyfa5arOFhEfNEX1Y2FTlYCFFIvo+xC+i4rnMx2GnZv
TP0MGEBF8ix20VFNRUmZnUa4oslEO3c5NUIqL0ySG9fGlFXu5wn6umIuxCfqXnsb
xTrKV5ZoZHcl7GHj2GLFZniV/MaXlvn+KhL5HUuze+yt7TwVDhQOUBUzWktksLSb
B3wnue4tmN42+G+smibkELrlyx5KCUzIR+X9dJj0CPktvgyxA3V9u1dg8swU8I6R
xmN73MwTojVIrdmDW7Qgey4Zd9Y5dd/o8d9XLDyPvVaPLt9xf0xbU77zbWCNVstc
IRjimroWJZQoEic3TqS0pNxAnImAWEnkENQf8/vTq+ahbD4Vj6tDQh1BgkRUFqQy
sec9f2UStaD6ExyBF42YdO2GTvVJiYQmDbUSAe7dm+IYZbkWWdfvwwzlnDRM9JJT
4gj70H2e2SQZpn9u7OU88hKzW5Cu3FuOPyGSVHeT2BIAhbZbWC8R0z60Ylc8hJbZ
nsswwdaMua7u/W6LwOtLNR6GICNoj9udYrWF8PTPzEFTpT2b2psH24zJzDCc86FS
96np/jqebCtXQKLuR/frolQ8/JT71KFwnl+bttrwt15BHE53b6T31AnvszRcnSbz
p0bimLkFDIWrvgAh7eCTzp2LjMQNyTxKfst0f5pJ7M8bnEplzCGX9qaZkP0cCsQb
RcZfghauC2v0LqG43sG2HQQvAwHtP2j4hYM4fwkLfic7lqkwfVGRXgHOeGUaiwf8
mEuAvYc6ENHIJnU4ADXh7obZ2PDTyHj3g+hfSNQXxEckYBJNQCgKa32/yJ0Wkwx/
m5QizJHp0luee3+gei62YaRqWjUubBOZNMjJKx8GxnIdwrdLcu/UbxOZScqtWZrn
q5PIqpbp/a3y6rsV6zxsC+/MU4ELi/HwhyUAPJ7xj3vnXUBPmZfGrilV8Lphr1XA
53sJ8nsH9ClqUF7QwubAtaNMxT2xP4xShQYiB6m0pe+i+jA85bk2O9mcu6VMeuVm
vyG3nAdU0sJCv7QWpRgbNDJ5LaumkKFi/4oWg0qauieR+Hoztc5yVMTsK0UF8XTa
TfnDBa8JF1pdVJt2POvvDa/94u8UHWwcDQOZigFixL88g70xRSR6WNJ6fjYSxdyF
cvs4vrIHXop/bRxrYBEcUdnukzVXaP8/9htSUocKtBBc51/R0l6GJjh4Kd+/ExCZ
BYUFcNwRttBV6uc2bSvJNDCVgBPYpQ3z44TZjvwDYWaYTpP+wghgBj6tnUDGyhzs
3q8TMxRUcjg2jlEelIWYJ9yKZGm1SXYHnal69yO9RPne26Zq6eEBDRmtwzZ+/Qt+
V6I82aD2qyxZB62ThF/Uzf1s91fRK69WxBEHqMM9nh1LPKaGqw6KDPLrD1VovhSO
o8WwrO59EogUKdJY5Bb7bEEaYu6YdrF4HUguJimScL8sOP28t6/6EraiiQuCqeCj
FaXmAcBo+IWuHw58QXCYMU4UXVhhnXa96lqa5Y/zi63I/nTagiGzI4cogvZvQXuI
vzOR6eTNPCkt8MPSE7NiThmMSq6vE2biCCAduCs6Rqk7m/da04jEex1S2ZRvIZga
ZW8aID3asXm+n2JW7dubFeqC+Z/xRdVEcIQD2V6P0PH4hD0X1lkioxiUgiuty2rz
36zK/PP2QazAeZ7R8sU3W85mnDbgK7cLMu0Zo9jJ5BGNq70tX1U31niodeZ1hVMH
EdWkciOc62xp74wc7LwVlHCpT28O8hbnmEfCbX+099jTyfnd/A0s/NzKY/f0ULgZ
eILx+KJibVqjJb1oUCkLPWy/yQJLr43p9W/Qdd8bk5Vlk0WlCV4LroWWMQGnRjDe
hoa4YP8ZU6l5mstgBnosU9McJVsl84weGCUEuREro6J6lqv0uiXj4CH55c7R84R6
UlOxHp8rJ8YNXtR9DIkGTEcEDVWxzY/A2vLQL8Hx567HNZb7ALWpQaEV7GDjd2e+
76wL7MZ8vmzse4K4q9e0M61IqtHOs19PP0n48VT3d1z1O/V2nTc8C4F2SPXZ+Sqd
G0ONP7jCN+lGtye7jJHlmdxqRxoyCC46R2yROyazlcrMm/Cwxw71696XhCuUVTYv
XaC5F82jDR6vi1Piwz14DE9DoXi97/DyuNbyefmv7BgBEo2KDZE16kzQyzDSakWM
GnIt9iFtljL9t7SKB7Xu2FXLG2KWuWUH1IIzi5PbJ9xPmOCXovw4ctMKWFoZB/dt
POztbobrvMffyT+HQ3ihmQJSy3gHZU2R3eXeQO0MZ6yWVwSUxIAVdRjKSn59lXu7
s4vA6TCMLCXhK+YAvDyAoD5eCD390rK5ZdWLAyd+dXI6vyssXk4RibwR8CkYlk7n
teiL1b6of3NxBbkvYP08ArPHbB4SL0qNIAS+mkHmqeMkEjqU/nTNI8khzezAx4st
c4AgtSmHtSByOZcHe441umng4IDoOL1PzisEwQZjfat3QKJgfonaXbSVhSoccmbt
nAnu8eegeLuyRGK8VUQex2UGcGOi3eTmvENbJKVvH4VdOdhoPcBqklphtvKxcbtQ
c+RhlPqLdPo42c1bGigkWRkOgUR23GJwNIqmlZ8MD2rnC4ZmZhyzIKZhkMr6YsyX
idF/Zkk2g7YefSiUYe67IxWV5qNOlFe/OH2CUCrQA2RIQEYUViQLiVHSS1Ixlrs5
7iYy7sdwF1Nmyr7JX7izhEbyBhfBgxZvI9KEZFxyVpA4PNi8hMICNJlU87FAV56F
0nF3/ZQiMuCQT0HkzTh2u+JNy7fZ2FyOeSg4lT1hhB3XNDGJ3HeXHQ5vs2DGFQ7Z
fGnLzG6jTSjkHDInaCtvHeJh5A6w21cxZDcnOMXo8VhmqrCBUIJ19YitWEYMQySh
7CY5GrSTwMBUDnXaQIMokseH4Lr7OtsNm3CRCu/ep5iuwng5KUNyUdTcMTcyKnsW
EvzRTzbBUolBs5iOBxW+nDVzR983wQSHRAcEnJfzjizddB6zewMJqz9oNV/Lf/ot
oIYddQhvlY865KUAPyKtceiPpGPKFkeLyyRPZJAjnL3qGKKvh40Hmh5V05gX2cZM
Uc8vN5ajK4ml5pom87wwsVxLZChazR+A74ujGzpwKnHlY34bZ4P0giuLCe5Hj9QW
EALKDeMBbdKYHe6QRIGxii7zbliDGAtQW1cI6bv+Sbi2c8qgBCT6HKk2+APgpfIT
JIvJgbWGEtkmLHiQqgtpu6UpUdviMRs+cdVbzmyuxb9GQ6OzHZIprHSt0PqCEkwT
TBLmO33avdwtDKh85EWJpTXI68gmMBtfDCVuwlmC9NXvJGojeO4hXSHkD9Z/dbuH
+bW298qyb6RwiivKHAua1MRZ09TsJTbH/StaDPzijsytr9gOG8GVqltHiw4zprzu
SsqpqzoCJmJxOnVjj5BxHcxVqCo02jXpzOf1gxgxcsMjmBUkgHqr5WikUTY9ODTt
OXiaT+/b6Aww4VXwC+5pn3aXIjD6Symmsk9T8ItYxH/uSJ2QDuGGJgBKHhdsUdW/
uVby+950uAPR8vcY/9K5ukOJApvvXHuvP6I2PWj9IoBr6vLifBgrt96Hbvta5O3S
Z5BvG4Q9QOUANYjXe1Y95aikj/I2eKS527pYQBR6AuTYqpQrWAborFwxYreqATg6
aj+21tIiMBBDb8Wd9YJSRsKDkB/5f/cQjhYGMrGVUjJvKDe/SIdHonT5pHpNKNPF
X998ZsyzZcbSDncMZ4R6ZtVzxzLZR3AAI6cZGQy7sGKZw0c1dvsrlqHkmxOJff0e
j674gB55Rh98ZqUqCc7n5ZE03iZ+uBnaom4t0NKMnY6Dill+lnVA09lpefbaAeES
aMJDoH3/byW6sqAjbncHTvsGewNa6tpeOE4uvNPZcLi0JK+mq8sFmEN0IrkezlS0
1C54zESrNmnvaK1hrjen6hSC+Fd/J6LbaYd7dH/IVpv+jl2HpVkH2YTdjJs6QEfF
Nwel5PXWsfs02hAANpx/TB4QdekWB5sQY2QamShY1grFMf0sOevl+XOSip13yTj3
OS8aLzoMS6hp7qESUoMBLIYf6k798gydWcNBw94YEtSJZBarWjuw3b8Jf9ZIcfmH
eRCSQgDowFC2UXWmmgfw/pksC4g6Yy3j5WIYzn2cwJyAk3jeKgsk7FHCRJAX6DUL
NOBrToMX7TcOBtA8RZGacNjYtkqhQQ4ATUigWWsW3MLEQ3pKe5i1hgsuNzJBPd7A
lqLB88uaC9e75vZQ9raXf7JolHWoxpkhbbRsik4XJhnX/6xli6q1L0dY+Tfoownl
+Pe4S77AKhiyGGdjrWmZLl8H4krDzN7VT2pYEetahOWzmR4YsSzelnES8ydY1wya
1o9KtrCBSAL0oKROzoBj3AR7IrLeTqXME3Y3xpN3Um3XgpGfJQPEhort/yiTf1fN
HlJq6/kul+FgFlgAp6OGJIHq4mZu0smyA+woX6+5elwmr2zcBTBgWpJ/iEjAJOSm
S48B3oxycjOzo1j7Ru1tqQcn+W10irNL0p5DKFfyC2lebNo8jBRef42W5nGkkTk8
RNKl2XpyunY16v5FizwWNgP+IVceQ8t3ZB2kLu3E5D4XAWaetUYHmv+y5DXiIY1P
23M/gEFVmFI26pyh4hPeI32Q6i5gSw6LG0HO6VF4VMm5abGwCcJe5TwAJVsT/VhS
sT9nvBPjAM7sQUubSvW6lg46mkwtgh5Kli91a+qEz7OneFQBvhhfCJKUJw9rNR/b
wsI/SHVYYpwqkhwlm6Cjqxa+2JhRNwHJ+bdsp1t/Xl97BKBJ63GNeBkkjfOZ2pMY
yDadFCK4/8gmuf9l6XFvLTrmXpfFnMHyy5dG4DK+JyqyOys8eB3N06NzVC+jgIyI
gD8dNUegVWAH+O1+gffQJag5M0MtJrg6Nd3ZPvzkTu/EDHp9byZ2wKJ5knguVNDh
RlxKVuWNhGkVUU+eB+dGjRKXTeezSFtDRgW8WOlz4gWbKtScnPMHGmFjDhIHUS9H
hH/Xlep5K5OPyTcl2W2h5ncxdUyc/rBm7F2BM4Gorjlu2WC8XBqrIbI+Z62Zogqr
yWt/bQc3FpG2zyrTD/5kFWozH9kgNKzR2ALcv7HZyU2IFtgtrpU+yuaI/Rzzoh8y
8GwwduxtEhQyaskN7LdpEVlR0vr80xPGkqnfpmXDAk+37qLLSKMx9KRxvJqdXevE
xfazmxJOPMadTIpQ7F6YeE5UUyMcZEe9YI0A434prok3n2a85Y3aXQZYvdEXhjzc
1fEprJ5pd79CAtjQLGfvbDmNt+TK6zw6RvqEBiYYcbleMicgAUppJQvXfMJD16ER
oPwaWxPETxDEV8ChfirW/9pwCcKBLDPU60YfnCN+hY8REDEf1CwqI8z7MvwD5gLq
OiSiTYgZhFecnqs2HkLy9irolvNsTpBkF8/a/BRjPBP0yOPI1IIl1NmHvrQ/uSmg
y4IcdiA9hTp2fROYDzje5oQgDUH469duuxgArKR9KYdyFDczuGE/i9dv1OjPJJl/
ciCA23jPtd7vqgWQSYE+/rXbIvr7Xo1PPWXDjvRrmv+QRP4F5syJpotEYBAh9ij3
6y2lWAvUSOMB66/CbhKOr4Yf4La7PL7TsQtq912NzFbeH7LbmwSG48TZ5sjf/RRC
kqoA4s5lJnYgr9sL90USSe23E+gzdtrWsgvokCOB9doCQs52VY2W2A4OpY/iBfKP
dY259aGza+jyZhZQaae0iA4ic3YgkDia819n8ig/rTZIY8eEqZZPwB0dxz8ZDKsF
uhwC5UCwgcCOmm3PaxtmL51jXM25kFITQyZI8toBNRy1u+Gv8ZPFYfavfq/UlR0D
+bxnS7LM9TxDfmuJqb9tsKvHo1On+yKp/ezsZjzYbn/Snuyf0sJn0YoYjUxEhCIW
YLT3odP6LbPU5PFykCfifTwHgiHyScJ9QuFJny54+psjAtLsrJ56oeI7pvfkiinj
K7n6J5kcVSneLMifTNtbvMfCyLafA95qtaqfEITn4louXD3JDsjKbL/gOb5BGXUX
NZLRycfoHOEgms3Zy0UHLo6xHm91OvGoNUjTgZ2OJyC9Kuj82bslttihtlg25dNr
HtF3CyC7lP5JDLXdUqdJzQqwOUMHe7mPXUzkJMOw9yPdFnXTqI3ZWAfWv8Yf8BFU
m25TOMfL8odtmqbuHP5C1Jj220g5wAGwkfECC1KFLvNufG/EOvlPgm883MOuIi8j
dp0yGSyTrujVKcijXuFJ1lDiJPdj6sWWL33qgUc0/+INXyQUawuZEqXgBUgT202E
nXNKESNjIl4wTZkyJk5WQE6ag4tXznkwCQs6PMkLAlW+2Vwi9oChQIXqr/+rhLsZ
H1N+bj/9pCw1W5x3zg2Y3OKYdCnsr3fwtuM7z5d9plmV8bvBTaEslRwg3ROmmB+4
gckTZ+TyKnp1XI3fGEeI+R0hX9RnSdmKuoPzInb+WGpD396GIvgdDK6tyXT3eFOO
F7eMoFKfB/ImKDAuTOp+4D+qnNXIm/gRjlRgZuBmqSSLPeV8uXL5iggHeW9YQaYH
souEhxCV+JkhaAmpHwuOKkCcSacW/ROAzAU7NO48CeiyvKIdTm43N4SleKtw3DBS
5pDPDa1CIXsO9hO1gc6ed3xWrUo5rADFyKi+UbvTX/qkHil7J5rnK6dPQNRvq5UH
7v0aZraPJTcT1DPcFah2q4bHAw2fi6EoXlF36C/OYMeX2cCZtRUVnUwBz6z+VhOG
98cZzSMCkW25S9FAKeF7CTfLcM6OfMSEzM8pcLVpvTs+5liCttEN2AQ2pw7HLNkg
l+fR5xo+EMTWJRInNxQvEhEaby0e4FkOVYRvh/9Airv8mx73y/2mEtVqm4KRZOt3
mC3SGuR3JzdNRiz9SxIQBVL0kzO2HVit0EqqW8gU06xr6qXgWSB64qFGmjEGrsmv
0JdSaRpjOBHAzmgHntpZYcrsh77hhAlH0Ez9VuVRGWfqdyjfc7Z7dJTPUru5KBZf
bNZB8Vb4BZ4HZRdG6WjyJI7E3htx94ZdfEYql9w2CEoo7/A9T+H/T7TGFba6iFPu
nab5I1DKvqtLmwfa+5gABSOUQo4BH6KfHRVaF1yy60s9HusYNMgTJ49mEfFYEt0J
rNunPf817tfXKYKyvWnfcKZ51+fM1KWDRPw17utWM7F1R1+mCkVf75hnfMBe9Dow
59/J52lQmZcaHcum2BmrXdYqnrEdmL9V1AI04cQHwpHhRdZe6te+ZaRBuGN0uwuB
H0UVbAMc9jta1z4foa6MmbOLgHscV3b6Eq1DHkZVs0Iz6T1NaBL6rvHY43LpPR0Q
nLJAmLRQN/fsUuvELOWSUrFAiqJG2ijD235uoQ9XjQs3IyeJR2R1Mjjx4HD8lcQq
QTxEYr7VoFPqAfaj9UoHpe3UMrRYP1wYMVn7TDyt93buOyRGqrbIJCb+omUuywk5
zYWaN/jiffuUNrx6i2rm4uJGsIoVznajxCYClriZZCQU7UytAgIdvIXIdLYMFi6S
s0QLcdMGuMcS7jHll4DzfEJ1ZXec0451xVjpFsl1BK3wDQxJ5at7QbDKXSiZR9vm
0dpH+yWVoEs9c1fwToDv8cWF+6JwmoEO/hyLchrEQh+l6Q8p+31wX3rO7IOfhuYQ
XiiXjY+xon8zWPzJ9n1Btnr/V8Gy12i8XptRICSPsrbjako+f8SFQhFUpPb6Edxb
BlycS3MVzhMNPnO3bl0CJJOP461x9aZGjEZRaXFxoM77IcKxTEp/ZwtChLwKq1zN
9RJpCv3Drq6LPN2PSJ4aZEaSYa0n7NamObwUMuJDsaulnCg+YyGz9OEYdX5yuspA
L4YlLrNPk5NUWUwOrVMU7rcKmoiISUk50qJPiYawzo6qHZDsC0Z81/au2cw1oytM
5+DZONpZSHRfRa314/FMO0q4mfsvwlCKHVjdl4bSQsJqA9tRnfUWaMJ/ZqvPi/9H
nPe64R3cykcmIFMhA/NeJ3UFqSfm11cAFmatCDNvZGH94FRU8Rv+pEJ37hjZitwa
cyBhL8WkFXqwov8UuDZX7yd8Xh2UBuWQIQ9pQz3dii/lb9JU4laZRdjiRs5diJBi
GbOoLwYMnZveq9SyigS5CG7YFr0YCvVlMDPNGQbF6pa+wXA9cCp2cP1xdPY3/bzr
fXtrKo5uTAHTryhObnXtS+sZLtG4v0e2+QzsN9T+MJqFYyYJ+xmqEMN0mKNqoc0Q
cQsBdppjUFobHaffYs6CjOpdq9pjSbKyzBVEX2MLZr0D2q3E8oJpNr7JZ/ZxAf+s
FiERKg+OzkTIsatn2ufQuAqd/5U6zUnJ7OtUOnrG5nfq9Yj2tntnDZQOp1GZRjU2
L9BCQ1tNzlntU+43RAhQc3Lapz9cZVHHHg90bmP/LyCv57vbloRHPZhNwJmUb0+J
nZcRpt/ZPuqresSAI6jHhTMWDdEPJ9sqcUHCDng1086P5H6VhzTJYz4PxrEysrAO
EdCIM/uwvD3GwAYCClyzfTOq5ZWwCySDtA8UERPRQ5JYl+uKoSQG7vHvXataW8ky
U+Nv31lqPaPK2eMoq7MqnbDpuWOyBM1BY6o7pR7lwcWhytxvekzOzqXHxAEBjcyK
8SPFtgY+p2OJLtLUoYUmbvAhL4Qcjl1ZqpNTxHnCkEf0ZrWTIyEKRocjIiD+OgL5
OBcA2PBDlwzzID7BBBdmqIBejp9cozVUvEHQhnwEJsAlfiKIOM1iqHqagVA+MgBo
20qy+81eYIv41aRBnDHDXbACkU808JodUpQ0csdRRPXRuCeor0ikpCxL/lwQ/jvd
rDZQGHFNZbikPa9MfdCk8fULApP3vRUH4IAsSEOXdx88GI9WE+VYTgo3FwVk1KTF
wODbPubNOzZ0biOReSxI9aRrcpADxyql12rxyXIvcFoV9xjKOm8dHoxZgn9MKroV
Og476U6yPojhYstE1qOL0nsfI3eemDK65WeUP8KtiwlFJM2RRBNTWrNmLXXfbGPV
kQZE6pRFu1ylhdNxSYk1GOE03Xq/Gn8a0JZgo43o1LXnplWyNhr4pLV2zrFHAmV1
SMzpLSbaBkHARxz6vqUo/WBZ8FcbP6FoBMps749PmwYHRNn6WGE5erTVKQ3ysH0H
g//GWN8iN9GIq1xCQ08SXpN/qc1n7TVuRA6ACIVPL0mX6SfSleX0/FtlIonsJZHs
OGlxydI51F+4tPVzLU/2uPKYWUAjHIMIc89r4MdUuwnHBVjn696krVpeoK++NASa
Hkt2vyPWtQiiwxz7NuKCcjN4irmN2m3xgMKMiJ+tjdj0OSlEz6YPrIZeoG/FZekq
HS/O3Bq9gjNuRnm6PECMSQS46mdLw8+njiF0bjIn6nAXTtR1Aszz79L+zkvxAgyw
tt1E+U8m+1eT2DKmrq3Kor2PKAlPY77dXdUpXfuTrWiehptuMg6jadm+ME9KFHy9
7Mt9BfD4ohpjJ60+gV5ALdLvmlEU3eHRRjOLOlDLS9Bjx0ldZ3GgMSPLlLfwJsCZ
DwMvGYdTosMqgHwOiuS256nRLU3VuAxvahwKn4tITwL7vwzvem1bXz40E6sPMwhz
u4k4UGn3SIKc6NNIqbKseiF08ct2Pco7SXeBX2kqBa0f8VBbATEiMfCPak4GbEl+
CcGTQEt6CR5NBYfpR9Mo6jWCLBzh9LJcJRRAUOQ/aT23wGTdO246w/urVwF4E+t+
qaU7GwdzhNQ/X9P8AfahMQBuCbCUamcg+bflDO+/Ygfx9wem/3XoSJ1YarGHXpDP
dSOJ3KSOVEds8Q/TKScCZa+4m19NowTKvSEJT46nU0K9JdoPY/gSO6B/RPIbMqZB
7iN+8U5OHTbtTEBoiQzMiRnnHRwrW7LWpqjKEgBGdECw3qAcp9pjVBVOrpSrQcKH
ozgUHxTzi+S7PJmnS55Q9ZWmcZonSQNRVmJufRlTs6um2xpGTDnu61mRvzA5UyCc
gH/tuuXAb/sjLuAMdtRxs4ZC5SqU0vozIWrEY03ZZwfpX+Ua82WLwtWNPKh55fht
cPfVjqLBNgZnb4CtMNK/cKM3B0KyQUPOrDDoLTruA8nNi4ZgfdNWL93y3x2KsRR8
LY+sfFuISUl/Db6JyTMo1qT6vbXwUHd9cF9JruT31L6J77WWy+P+3Os0HeG+soBP
yXMCVZpWSszxFBeISGejQ+qlBaF63LeYT1qoV8w7xm6YQkZMqi4ND1/QHJwxNBR2
uw3YdWE7uZBq2Ai4CdYJgHuLybFTaYSICr0Fbp7CMKx6JlB/wwK7KErHOTFMO4hJ
Hq6deI065f8VTd5AfAjRKYw4kBFvotzP9GjdKMgBWz5twWpj8LcygC8cOJ3F3Tra
7eqZ5IkLHBUOu+stx0VK8r3gyvpUQ7OGx61T3ovRuZQc3H+bNZYzIZ6SObyJwT1M
NIJBXV5MOMzW82Ye4ke5PWGDHlV04gL4Fxksx/CAIKGxp7eLf/kzA72xAFUNBFxQ
hHoVGafbDcudQvEs7+fhFtOCHepjU47JbhnG7U2dOX9WQVGO7HGmKHIfQDngfW+m
4R4DEQSdpina2N13KAaDAaH0mhlexgbTbSCFUMo8EF7qxv4Qhy18xsNRolQ6YDRz
b2rKufbyi6lIKMwQGXZoQZbvQz+GZG/unJwTVjKEO5TWEalSfIk6yAPXCR2F2Kun
iPNmKDvifF7QiDgsfd9AAvGBRhSHokjRxDtCWb7RSOB6NBjifKa03A2N+aXeIVCm
61BltTu53d52/cBr9eVzmfi61qXQhIgswIRyiYx0KsWR9U6x19o4Kmdm9Mzgq+CM
/73Ge0TUp59k1f53ZZk6Gw+Dae7RjaXhNJ34QMp3+05VrncTmfsBG8eULBuOPCn+
sYWoyCmAsaqWFHJklDzzWm0jB8mzWVcT0BJETy35cBKzPhJjZFlt4zEuuvFVX9Pm
AzB6EP95WCp+WNqfzFYJHhYpztdVDCVZV0XI5qrAnwdOmlljOzkRJF9bwo5vMz33
tyhSDuxiJkAcxwdK48EH3aRpJ7daq+BUSg9DR0jfgv5NdGG7y3r/LRZ1GAbwF1II
ckYj80qeTVzgs7U+RLcGpeTK0AqNP7hiCWKCU08KsuTjt9tJMNROYLzpNWxerUvH
Vd7OU4o6kgpeUb2P1chZ5cC7Z+t8PeHT4qxdIkX0AKxzGKqrO29cynC944snT1kG
9NjuJOChgo/UuoYhuVbmN6hNXVabL+Kfc4Nk/Dhgis+Smq6IwsSkxpRKiZTISbmB
FOEOuMIf3YC+O/3NUY4ys1tIJ57jzMn4cxJwOTTwwdAiEAD7ud8VS7GwWbtZh6yW
xud9/y/nZtFLP5N50LmaZ/pghCSoHOD2QBD51glwfxsxBqDqe58d0QcnbtUCvfJD
ZIJ4hKoTxgk2EghpT2p4SiDDPMOOTmF4jRIMQIdWHFJ41ycTmUKXcFA4jU8QlFCY
DM+OFufApa4pFOR0gn+rfBqlmv+f16Y51kvrpI1NaLfqnBEACnAmhiZvEVWxTSNa
oqccHVIgDAszPef0qVRDcrfpF/0iJYgvyqAT+ACUBmvVs76x3NXPPE5oSMxqDHOG
RyVh3YDnddLNutbvEMJzFmyHKu/4236nlvCsXbxjk/W9XfE/se5aPJbE3yezqDVy
4zDJbLg0xtyreVQ7H9oCvQpottjIaNFKCrs2AVfNg6MJkezbRQc65QNL5iS1nRgh
uH2EYH7wC5Rzh+RojdT7mZjhThfaLKI2ALkzDEh31Pt+uxhs1yG5cGMdbovH9+tm
4C1nyAyTz/d0i+tWQIdmMmZtYmmpLzl87zgEs7kOAQgM1nHNus3S+Z3YARdUxncM
H0ZHAGOelqellguUjxNsmoTIDk4PzkoRNM4/UT5b+JpWLHR4/37HGIA1PW8oDhrZ
0QtldD09n3JA86+YAXOe5HA9P8Y43f5fqNElKOQ7QfuFN5RmwpJ52XBJrpopPPKb
OI+NPzOnHuwPHH9m6XVHcOm6kNtfp9k9+y4BnhYuLpbl4keV2068vuBxDANYcom4
Fh+pw2keyrwSU7YgEITd/lWdToZYjV3s38rIjgkaAosXVaQR79n9lLoGL/3WzFnu
sDW7kUlJ9+bVIxEAb6AWt2NYSkZ23OcMDd8fGGIc5hh8amK0gCejVx8DOyrkmhXj
kSqaYSm+oQG3DN3WvmucyFa3gND4VYPjw0vBai5cgC2oLcIta+jZ3bEj0oKzwev9
vBnTCbe9tgS4bb4dzV0IBecbMBitH2LAl/jdvkFBkghy+zAXMxsNbF07Hdv8FAYI
82L7fDendxa22dD/PNjIo2fVBr8sF9OYcrNhoV9hn3jCS44APfWrs6ctHmD0MsEs
WJuThQCTvYeDWXLgdJXXzAH/58cgyH+nC+M3SxRIhecjQofcQJd2l7JmKyNubU23
+SGRQ9lwjybTpZqbsx0YuEX/BUxcEpw0LnlCFljMntzH6cY8QRy99IlOM3Y6F6Us
VJB4FOcDER9lFmWyAj5qI8UkHFRazDfSXD7RfXNRE2D7knU2NOTfxDYcxv9QGcii
gXiDWKzQtTiQNnwwMpX+jCfM1+KVC2kC/AUIPpmVXO/QG4bGprpl888BHPuQ3Wp0
0co+nZLYkotroGSyLk+k2XJp0slB1JVsRRFUZ/ziioIZo35II0lNedvO7Ltrv2q9
coBqHi7fzr7NxRwlV9HoWkk2A4dqhJa5Bnr5N8sB8qjOBrB2gbVBgkm7ZegmTssz
18CqRW6bmjnhI/kAwsyJuMGoVhSo/00JFBGv7+jDYousUatJYzgFmobJqjolmywR
JimLRnr7cg5JY4/bCLW3P0dnwqD1mXCl3zD8loy3K+cGNLSGlNieOtkOPW7z/dmX
yzrfQPvjrM4nBAJc/dxzuscO+zBM7Uh/EVic4U04KFcktC0j/PereeUUPjQTj56e
faLkWcWYC0Z+fZcTnjhC5+DKVcxdGvaU3ns5d/K71uyXl8F4daxKUN6sLheXwiU3
P6uZkdO4cw+0cFSsuq2/vPR1YBucS/GVDuXKMgwPmX1V34jmuQ/qJ/CuW6ooEKK7
QBwoSZOYYZaG81Qm9vV/Eah/VkvT3jzF6H5xmMPaf8Xf5T1ul5/FMQJoe1D28EPJ
HrnBjzbbfR5OLYnUuSTTYLGthwBPxtkzRJ6qHqKswyLkG1NOuduiZ3v27fce3fDG
fR61XSktPIQAiaeeJXTfzuOprOVYhAbAbja8sDZwt+bUptBgIQVo15ez4RdfFtiy
mqJALu3F9wAUtigphexXCKOHyZtMICmP+IRRnxPz5ooScAebwNRbXH5eQIYUnxpX
fo6LvusO5SZ21EG54UYMWPbeH+5FCibARdGmA6y0gI4La8fh6m3JswvVgDbFEh1J
dT/LaTf6RtaJWi/9yuamHmpGkBLaYk18ji/BhysbocLJB5KJgW7IBgJlvqXx3CTM
ClcnfFWxabOv3GSH86WKf5YZykFJOKCeaB2QqLriBE9A0jDai449NvcI3O8vU23v
UCDkBYfQAteyfbKmqcllI4TY7QgQ/m7TEhxadcNCkhxpuTDAaJum1V5VgVeUaE14
Zynt8VggNzxoJSi+13AEqTdnqOdt4KhdlkQuKZT90V9WN5l2bgL6jRH4XGpT7t9x
hluIwNcktFsdeHlBzCtm9BWzqtSy8xbXj5wsz+AL0J+3rVqTTXFcIA2mSjI0enfF
gsQghe6GSd17zH1l4jdKJGA3+hf58Ymy7Rk0j+WpQ7lGioxRhasqnaf6IEWcjgi6
C195ofBVn2Px1iZwJQKEcqG22VAVUb+izZeF/f9THprcJIhjDGtzL5yXyhEXHsJl
3B7oSHNzVXyDVgcXRarzhVL/1u/GcgpWoZIYh3nfelKw6xM/frBUymwncHLhlh1n
sRPOZdx72jGJmEIRRpFdOUEIU0jyQq+wz0vOBQbvAlR8vRtcvpvMDPcNsCh01+VE
1BLH1Vj1eG9GuqmUqa0jh7On3cerrZpHP/uynB80BgFwsW3Nj5BLyaC/3he9PgPv
feXCpLfWmmjellXZUyaOA31YApLW4gg/cRXbpvktuoy4yTajBFvOyAwlvW/seHXd
O4BCAgogf0vC8lDb+xxsCd1HYWl2FmeeBls3l3MlVhkJLik0vE/5NsTXJLJpmGBJ
5pfC29B5u3WmEtK551E/qLVXa6YkPwTzBR1quMuhU2fCUtMgJuz8kEb9gNAUxyZ+
R/xh9avX5u9GrZJUpuNjF4vMqkxZgYvqLBw/m1+qpy6vs1olYrJK1N2o0hU6qMWn
4Hwev3bOSodhYVIbwNQ+PlLUc0Df2XCbOhXzooHWTB2KyV0bOpViA1DdqjS5wwnH
7LAzWrMVrYb5urP5gL96D0KZnpEORXmfHHRC5sIoAa9HjMs6bWrOgjHsKKugNENt
TvSc1yQiKoIZ9LSI3K8NUKfZHZmTCpmuyL8fvpkgawF/WazRFHBIZQi/+Qk8jT14
d42bAdqviiW40MrJYsMRCRpsDxrBmWb1tyR0+NUb3ifzx3iW/d0GsdHb7qb2YONf
ML/TICn3y0I7VslOuFut7ZejBPUaDR+b4MV5fvw2b5LSiCW9rbIA7cf0A9/aEE/9
uhEGSgq3L+ubXLUTm9ZBLZRpcZrnk2mSQlVGUggrT7BsVtjdB0cFn/Xuob/pn4t2
2wmTtG0kH245ZsqszsJQHMOyQAUbGRLkS/V/4YblND157XLf9WsoNg5YXOitLkVw
i3xo8E/2KmLY9kWn8QDUakjwZ9a2vwaBexXe8rFHftad6YGsSt+4meytngmABZ/5
QZzxDQMgPuGjdeIBQ/Ejl757UGbYqsZF78TItD3e5kbPV5g/wUUAr0MQruu9jn3b
lqsaZGfEYZj2ejLARyhVZ8VusHArbSPvf24AKh+doY68m5I7b1PpIGbY9QHOqHxV
ADVnbEOOgygiAoRixtwqN5lrYQTzEvm9ka+XDMiYdFdEhd0qGdlLMd4gi6ZlcjD7
KV7Bqrj5k/IpYarbCvr8jz48pTW7PixTbcmTtXRd5PSmJI6fIIHVB22VxbUg+FTg
10utE0sGQoQEUKIKGzCEBB4tEABq9FUq/A2NDWHs2rFbaNX9bcFDH1ZDOWWXqUzg
Vid+/LtWWTsRP5/ONRXlvMxeoC1IHUJJHGNmGDbgAhCWXSbfHoHDT+KYzEFQsfDA
gG1IX+uwtO0ckidCYSljdD68CqaXDysetuom/9nRx3MCdESOx51V0Ne6QirW7IZf
J3dre/sGupoUrME5SzqTTsHMtiKYm1tLkycqsoIVDOypx55cUyeJ/7piOMnCkykh
w8bnFCFRCIN6mteEQvDCCW7SLYTs3aFOIVPA2xGz8kjkUgV4ByIaC6K41eUz9s7N
4sLaWzMvCRRqjlYqZ9cruRHEmTBDDa0sYlSBpM0IyooSSQZf+L+TUsrtuC4nX3e6
/JvMtelC3veJDXVAyY6NqCTQ4PM3eNqsRpKbln1vmWJnsFsUGBaHDjy7eX1oMbKf
SwzlZEqsolrrEMQArKfyCPamdX913us/VFnFvjj44r8d6MnoSUhkGNVg84deUndy
uLM54z50eo5BQ5ESTVAkuTRYv4kuj+gk1cVBmgC88lKcqyDzXxnwUtAeWG5gT9RP
0CR+8MDP3odrSnNQv5KHXhtJPDh4AryyjL7w7PWjLJU9OkhQWU4eMqoxRoACZ8SR
voqPnrLjpJwxxInG5ZojVceauK47XJJhkaK+aAYmFhvP2weOAR5Px7ED5BMtCrE2
FYRPV4+MjaI3MCyEX+e5lhnUtI16RsYiDPvCwDnWSkuuiAebyjPsFMdEggTnvLwL
b7ewRjsctI1HUcbXFYKs4G23TkC/M1NdMZDdzuqQJGRSQzZv2J7GFbNU48t0usjE
FOvoAYUF2xkmEGQA96Bymg7lAm3i0HguhRLDVKw6RKjNOGlUU7MQ9xiinb7usXaD
OVcYkSe/ZCk1ZJ2Hw0VT2rzGJwVOjYz2SNRiNaArJHRR4LkjMljhqBDlSBQnJQPF
7Bm6avdMNvwDeQMCbTEIlJetQSfJty4B0TA1nMYkPQKHazUpojUreZl4CtQiKyj+
XU8Ij37JvDMjSts9x97keovUUrL7n9gjeuLfJzMr1GSf+Byzf04S2nnN91MRKvUw
1D/xvuYg2WWChLVJVu/lF0SU/fvBDIxHVzwyjfoAOC9b08qM/6ok9A3LoS2IMBIc
tS/IfgzcPT3XdQ6ZLKWRZBcv3Xgt+kKvnpDqZeVdSKukGKcDqCFYqGuTqInokyIS
hHhakJ3qn2vlPxWg6eRh7OcxjFTbeQYiWzAaykXPb7ErGjE4qK5YLdkAlsERE8Gq
TYrVHDD+1XF+yBiq4xXM1zRidUnoXy2Ysm2EsOvyEOrAb/RcKptIxEJhi+iUsT9+
s0iVwr9Uo1gIBYKMWZpR4HWKz9+NJV1w+4DeXKWHsr9tvkdSjQ4W3qNbsL+0wr4/
E7sH5EjMUM5pWkLf6nv/DnucTLr37bQokw+tAByUGbPngu1vDgQHglNsJI6JJfjx
UQ3rUuevIVFrpkesK8HxGxabxdzBpj92ghyDvf3CQf0tWmw6CZj5T/ENvf7OdXso
8b92DFdGrpKXKogl8I5xpu0pTICdFNBMrerJQeUQNe0pW27EaqzeTtVQ9DWNkW5C
cuVVqaJLunRP+pnJDp6vxbSCAu5w83J7yYck46QwuoGeHfUTPYzrrw56anYIEdAq
BW2CHDot2OJymEio7KFnpsD5VBNzS2AVI2JBtLjZAAVy/8aHiNXXqbzWgNUXRz+R
yoi2/VFSooU41t8t9ThWK8bmWtFwFxgWuLPREF/AhYGWJcSmg6yxSSZ0/VnPKIOI
Noj72kD66JUns7rq7UYvaxWe6NV/2lfDK2OUKmg6zm2UJ2wBfFmZKLvrKDDxYBdM
tfFPQHqmr8QBQEECO+NJDBCa9NNfjY8XmHL/oUfrmbnYYn7PUH146EmaVz2xwSl+
QF8NZXPTUeXQTiiIJ19oQDLkCaqkDvjNzPgfGHAizH43cNGn2yrDZwyx7q7B//tl
vr9AEujt2xTTbWPfPT+Qe42XJlVC/RxA+XT4fReFuPuXjNa/YPUo7pExVM8CEOzk
Uy1Fgwn9SkF5wFDVjX6bqwyGxjqU3rSqhp3NVy44/U0JCs0NwN8UrLpsybKjR/fO
RIUSP60s2GjP+fq/cEau3+S2aL5E3a8WDfMbzHqchx/ADsW5VJ3nj7WRnFwRMe/R
CqNNwS3W9Hjl3+8oSOXoUM57Dd1pG24tuydBmEhgfu+TRLeM0TZImK58v38M0W++
r5hhNZC6zwA6LP73QKJ06FAxflTH81f3ZjeA+RzAq0dxP7d9jC1eQFd0FLv+EMD/
iVyygCFuniKeUQ4IwN7uwT5Drb4rkVtkWRK38oucdzIO7aHLjpwgjHGe8CmhyA/W
EkmlgNmt0//vKfne8a5KTqm+nneTuNvYajnKRX+nVdVnWz5n5kHIQn1+mCnFzbkN
pz50vTPAX7Z63XMJehI/N7HyXCTsXUvnnbrsWcOOYTzG1KTBVPf9aaLMbusakVu7
sk1CCgXfJpBUPAE6hMe1tIXmSoLh+mMaJssOoKUPd5EC00KOgN1RqTAyrTYxuc1q
q9WrHl+YQujPPCBNIM68GqhXcKuq7PcjVtP9zX8c51x4jjbvGXTugtemKvSQSbTb
k3J19PZoXWDx0EgTc90ayCT/oIsvAw9vOGtPQ58ypq70kc5vLiNnZXm8a0MJV88+
qLtnW4DfzU4a/rhSWbO/gGUJ5Mlt93k9LYloETR9yUbPDSMq9E6iqbCTuA34F5wg
Nuhh7F+iygvsc5AnqhEH3oBVYkD1/exzVVJPAmb9Y1A1H+0rX/yls/xsRyMMOxPP
rSB7hHJa3mJV+HfwolfNd7bhNjUCoPWWibetSHhoUVaf9I7VdNY+fjdipErArZCH
KMzUSeZEveuQ66dEJR1zQkPwlbr2t2tg7ZgzQnRau5KPEGEdBk5ujAdZijro53wQ
qbZTSzeeU2iH33Mjb7m/QOix03xR5UA244ZVSwagKAd3U08oLpAXADYMCjv7EhKO
Z0txNuYsnDAqLR0iP3rAIxyqlhGBl8esrEFO8k9CJ5rOZqgcAN8rIUPhoNhse2O2
QEUcUpNcq8spvsKFHf4ypKLn3JO0I8jdFGUiOkVovB3uigzkAa5Qdu4SH+yxCELo
5jrf63zvpppbyOaTr490agxsixYEoqLpkmT+ItdB8/QXBTof/3LnMHl5No2Z1iNP
Mm93SPF0TeI5CSUaAzFGTsw2nC1cTQgzv24ldnXe/cKk9KcrA7nVaDk15Ow8HgKT
agj32iX3pns/+euMJGu5A2oXJXV3QwMN11UszcJR9ex2hxryGwMj6kjr6zlVXqS1
v7/4TMJyGvWPX5Fn1Y9lrKj5p2ZvYIOT9fw70bnIKo72hQ2eBefkslLrB//zsI3F
mll5EsZNu8FdsBplAbiGppTc+0az2L5E54tDjRvKxogmL57q+cL5Pzy8wOLeoq5h
7dezEgZvdhL+DNn7llbWJWptZJNA8Ezb/G3iDd/5AkwHNUi5AiKz8AXGi1ZAI++T
O6nCJ1qoYhpw/I4PStZiuLFdqcS6qiKT6VMDxBfoA5rn7+azQyCAJ5ptCo/DKQ6j
fC+p8HL2PnCmmLMbBLVVBCjWdZPQ32OBB3mdY3LlkZGUeXnCcoI8jqIEirdFSnQp
MHqFzHvjbLCzQ1t5wGDDN3vrHy1Js6cpeDGz5U5XguR1+FSJ/dL+3Av39XWlBRaF
qwUB/VrgW78lF5nbbXqz7RPJ6OwDe4FNDNIsODg18pJdOUOwVcUNpJqBXYNs82AW
4+BgYGyStTw3EKfmv4AjyXTOrpzQqOb0ETbMbrNrCj7aN9HC/O6YOmsPWkrffGLt
j4SI7VL0otWHGnC3sbHMy/EXSfD0/Gb7UISCOrJYY9ZutQmBxLo8cOkoYWv0HYac
JZW/sU/yPriKPD5jNYgWVHAOdcH3CHhyfJrDe9Xw6tdrhcUr3DCCtHze0J2QZOlK
UfVT9SMpHrBdhUxaBb+vxygmGCw9FBwZB2ndGPhlDd7E1WcqFKGZtccrZceUrrGs
ZVbbtTRG5QK4rGEowwduqI1OULXp0loYZtSXZoMZm2Xrab5o/oAPhbyDpYW1cQgG
YSVNPOUxN8HyNPonwnnOW6F+aMXKEyrjaEagZUQYBBVgvEiOeQP+J1NIl/sigsnB
OqahSfguS1vD9NNqkzeCHA08tqOjRkbEVew/+IOWtLPKMv6BZiU16hQK6MbQ9gH1
aexcZzj+99U8t6jyvGtV1/LQWrapL/Ty5N4DrkjtmwOqPZjQmOLI2vZQK1GdVfLT
ae/QRql9H6J8hhBCQxo/sfRyifj3GMqK+xNJfvV0qLt5D16u4/mF0Hv0bNhyZPcb
nrwjEibhQ6ujVpK8pC5MPGgzkfN0GA5VxOa2jocnrXLdm1Af1OyNr3Z4n47rYHd+
4I0oQHfFHP1FRfQqJag1zL23bBU+NxX39ljOCebWpwWQfGMESNpYaBIM4CrdEXGs
C7fTImjt3TGHzj442JP/FNS4j7kRDfsR5LB2pxEwv2xJJP7PBazalu9XFiurRxOT
JEYqc1TtxaQ0WTujgF2oX2q1byV7NTxNQMoiKOqbVLh+81nmR563UApn73va12uZ
9OAsR64m0Hi4E3Mr1Er3fhewItKaDsABMfBFXv9XD0QJbmip6LaXWiVzUjAuvCXl
W/5ZcNW1fxlgPKM/v2iBaKglbse+6tXtFeT5+3jjE0RRDU7aIukZcRK6sirJaTK+
WdVhHbOmJSiaLfCteTL9gMo8PZCU73lMTaPKnuHaVXwANXAvJ4Kboa9krYZcaX05
aV0N7zysr0tdhSTNg5Qh5GyqJGGUk+Hjaxc+Q4GK/SrloeM8STa56uG0qcjEtV+q
5IP/E3e/PtD5W4lu8L6W8mLzrPnFq24BZNG99TNNgRYZIfmmGCz3azgQcUiLtJvU
vW+4KH6EEtUQ9x4Qqn63J0LUMlFhdJu4in1TLZdjfndpZtCB4eSwz54ya6oYrGEn
qPtgo52Y30fSLkgrKChi6ItYiwjnASG4gU4Aqr0eRtgcf7I+0m4OJ+el4e0xeEzh
mXPtnBor2EdGBzNLB09tzRlnG4E7EmltCvbT1W/e8tx8rc+67ZQUMgnLPrdsKyJb
C9xTixmX/1PME4AB8/2iCddySysI6SUSxY7pJbXae10InXHcoyw9iuiIrsLg436M
GfDlXUd0HBnoCjaDbiStGwCbP+csIFmS1vthQKEu04oYO20V1910d2xaHr6Fbwnz
0gqjw1z/tPthw/xH+h0Pd+vn9ahuaHQrfAs6fBZkxarpJyZF/WX97KeLeCpZCOWC
M83gEQWXtqcF0E84WsdmOuF0OCyV8zdP5DWihBuRjNJdG2aC3kTXkVkdk9YLF5E7
xx8DhuQQkn45+ysyQ5EUsRVAcv/P/S/Cq2IZFDqwoA5YTQKBmAVt760yqJR3yFVn
4HLWxIvrWQM7u2mKIXKKYmeQZD1OSTnyIj1hHkZmmOsnHtnQlRM9+SZbC+3oHYlh
vAv5nQOXPUWoBJHMgEqeTSaV81WuESeHcG+dv4poMpDcUD99h/jit/zzPJAMv3vh
3JzUWWXYuJQ+dgc3Ra1S5/BU9/oqXu3oY67IU5qbN3DwXk5egg92K2lYibe4fKVW
DL/LPBVacS/YtTRGdhA28xXJJBHl10h9gFRyb7eHFKbMNafmQq2y4e6vbSdudpEL
UfG7pji53VOP3XKQfNyzNfoMIFcIc6p5H2wgbUvQ6Hayprhd89A8715xOM33gOmU
ozdPktoNvrCTCIuH3CT1nr0H+ZWpuvfNbZh8rHJAVO3RxbzOdgdwENapGVkGUghk
FHQSlwqkJ241QAFh2B+VKzvGgj/Tqy6kML5Vm/wehq+EWJ0yHH2GMNPKZ9CFpeoe
Pec4X6hROjYdGc9lHCUh++09IIW63SJIxEFZBfGqtzdK9Er0b5OF7Etnbi72+FY+
Ydpmwn8QwbxIrkLk0jqIipizV2At1YsJv3yDH6YieFvuHd197rfXBj/fsHepyyR1
+ntJmYUefTRCat3P6Ai6F9+BJ0oNXadNJEAyP3HWYThMpbK2mMt6VKdxYugIhcuH
YfTBl7NWqqGz9CBQSLbRdhhk6KFxIDko3xCvTCwUHoN1mWMWmsXHPN0noPOk/XYz
ipFPi+4dGDaLRGmPo1NLyohEj13EM1QIlZCD8bcOqt1bQAicX7/f2RXJXBlmNEs/
NeisMTBFabnIGBslFx7iQShLR+hxA1f1FXdhrQed9TZf0gMsmiRKVoOU67128EDJ
yFdG54BGS0GUtvoQh1vez5mg144NN3LktdpsBRy8zIeZG/yTD92sj/BUI3ryJTfV
eETDVllDr9cMV9bLX21uX0pRQX8RLdUSM3tLPz125Au+hfxspgjKvPQNn5YGUN9q
gvc2vq0Xn3VSsxE7X8Q/yIEZ5C+R8ffxYorvT6EQ+R/n+8clVCsAH7dXWZWDWIJR
hl7xlsZN9q6xKcGt2POKm3O68ICI+bkii4CpvZ1Cq5CAuOf2Umn/6/GrnLSJES/v
nm3OwSsHFfj//l4/MQFGSMDpKbo5YbhghKMiYJbTFfBEjMFITdRfDNAOyOVlKb/1
7b5ygaAQSldwd5KZa7l4ERVj85j9L9D527V280zduXED1qQpkUCo/tuyRNJBpP98
b7ZAo7wpM+CsKpIs66BFf44zh3O1PD/YMV+bUSUlznmJ5ixuN1NlzxX1RhYlqCKm
T1OdDZc4A97u4lcjU57I5dVNsDUToxVgh/hYGEO7i2y5RZ72X+Boyl5vyyAc7rCt
Ad/yjt8d9UL0yJHGjtGyASJ7aNwxyZupfSDt5TqKdFcphthRript1KBBfXEDcucE
UB74LOIeAKbCsqcvbWnucArKlP6J+fjw5uckg6xvnOzw18mT/sPVcicRgHe4qO5P
4uLRHZE9iyE5JYhRHc2iOBJQ4Caksi6cABU1DBY3Ik62uFVQ5SBSFKdjenHuKR6R
oHK7tIsPE9ckMMaQlG0ibv7D4YP1oo9eRpqc91HkfUPJgTgftsHVEeeH9S2CO5nN
e1UKvfPKIFZTrvsABPmVSkaPU7TKdBeOnd3qGQ+JmDe379xJI/wPbyOed/TnMgE2
2izBF5P7iEHm/MBuv6rnMGG7ZWdCtVCqsxc5ZculZ02kesdsCisa4JKFM3ch27f7
a4x0Uh776EtI92Me7XkvrWZy6xNsW0poQmK09sgc9SWRsJ0VMxPCFtLigzL7mp9y
zF4A68F6y/ttoQH3sMByRQxDNqPLrCoa8xcmFVy1DIlHM3HpEM+XUpuH3Ra7YvPx
Tz6jn0WrffIKx27BF/BaN0CL6NsUiBmtDWuPcEduONq/S7wOYwRlCCo5WeP1D+GV
EUPNr2baF3u8Lzb4H0VrsZ32dno1lMSYxgUCgmlRDq1kPSvwol+SVSaA9WR0u2hX
k775E+NQMZAm/ekO3x/ozSxpHNPtM59ahivU3b+SchyzYVuTXZsZasNDyD8FriVy
Z3HpJEhu4vmJzsxntSyd6qiiLnG/OK1Vb9KbjYHIVJ5vjJ8zzQRhxGaLb3ndwYpu
45QYqeRMFrpVE5GhlCJOFOpQR3JrSIXieZdptCZ/C/jXW5hE8F2KAPbkV6brp9rT
H4kgl1+cRkiYxFCJLEiMIZEHoSMPzDuMTO0BOZ1wIqTBf92v9EN0PFlXm6jyy0/k
FVrY9InZl4kCV2swRRgC98f8INSS4D7qmq9kreA30O2npC9FWYvTNrvHQpGuR5nM
ZWLrpludY+UJFbBHhauYcskr4CaI6Oey+MeJ7I/YoT9BRX8I6X8fEo0k1Rqss6y/
PSUnIBx3qv0PaepVzNlMefOQl2RQy3aue6Hdwz9jFpf3XtslQVvNSxAlrOJiOCld
y0EPYSZlGxbfVs0jyFnG4yGMvml96fJnUZ2k2gS3JPmznIAhIqCeJ+4o805iQrFd
jGu2Ese08uVcgDwuPuaXuLRBWJ3najr6aTEcM+6T9+fk1aHqJDnJV5cJ9jFxXMoY
h2htNZkI3psMgDqPBQNA0QKk9wJAvpsesyCTXba305UoS5jayjnS6bXfRAc7EuSw
V0eu6sUcpRBuckFc+Z1gvACHIfWOMMGauNdzSJ3P21cIxAxk4UBZybJ89prTvW+J
c40bFqZ+YTjjzZm+begRPl7EdCuVhZfNad31TdmWK4aB4cJZBEjuYhfwRoihOXO4
Pcbl+Xz4GcaUoQbyZVkLLGeQM9MoCz8FU4yPN45OgEyedR19k8OX7CntckOHqxhR
QGQ0jprO8a8BAYbgSUHkNojLe/muhNKXhcZAVF17M4ypn479+ABCUL6SHyv7fau3
SAf2LQWAMumrGYTyLO3qQAxzsh0ajTxIgwkkHMYO6zW9EYZ074F/BTeRv6vE0n5f
nkQyi/d+V9KlMjs29ZI5RbH9crgkqg7YQEpdAZ6Pz8F43WEJYSUtYU/lc9RbBkNV
o0nXAjCculIUUmeRthxL2kpUzMNBt4Ply4lB6jrasjVCqM/FCyrS5xovMk3/xMMl
HCNdUKNNAV4Qw1kgdrZGfPDtR6gJnRQV4/zZiUoUkSCPWHy6agcgmtdxvQQBZHD1
Wg/kr2NWRrvtXJGiTHtkoP3oX643BqOZ0eNaRdJZ4reLCSoHrVk5/Pl1fFNcKVjZ
AmbKzZcmI/uhnSrDSimJHMeaUy4Wdd6+3ncuK7GI+7SM2+AQEy02GkSIgnEiHMI2
s3WZgZ+CiM2wuK80AKqN6p7riy7s+RgPwIcqbEEfh05F90GRzuzgXL6cJdxNyeRW
19qNYIke0Ni73kcJxYxGZQJ9ORc2FXJKaGMrP9jcIIUbYLIhwao7sagPyBXRbPPT
8L1H4VNPIcwV8GGH+iuPvmqk+LHFbdQHbtJrGkZRGH8Euujwh9wl4/ibfKhsttst
O6g14c8apcS+NJzHn1g7jYOIxuSBlGct9UuK7J7SiEgaXnlYpQc7gHYeEw9mHUC/
ie2sTG5YFRHUkJmVIvSIx/y/0l2SFp9WBgYqdoYF16r7HcYZGq+MdKtVnMbY5Rtv
7C/ok6h3YupNxZpa/FWDuu3j6xkEUE/sfpRBQ3N3SFRfLBThS0/1d9PbfzEjMlRz
nrZTlOxyusj2HZ44NCxZIWKxlXlhmkUd7IP7DVaFKYhhpq2NNixggm07MCULye7Z
oNxEVBlbjDUPMQc3knAh7ZW8QZWlS0dsu+dlp+dSG/a0FS9f99i0XuH1RZrP5Cib
UfBTDTgwYmvy8tXiiV5gUT8hsMUs2Gsu0RQfkBRtuWy5DZMCr7DXbbK4P+A0dntw
Sw2OXPxLF5K0GEDXcB4k9ZQ7+FsqReIzOqlP3CKQwfo9mOJmd9AdNynAe1gIpx90
cZq6ZBMpEVXEASFwxLV8TCRS1flQPXNmKhWgPzedZX0r96vqBCeXz653V99g5TD1
X1n2B+lpLmy0IOn96ccZ4UYEJ7regtl/3ECt1IZDZRcwj3R/bsBjgwZtW1r7Zl4G
y8TUL10R21CeEK7NkyjdCaR6z79k58MEIPZhrqQ2izGpHF4lWeS7asCWsZJNA59p
CAfsE7S2bi6yJXT9005v1jlc6XIno7KokeEw/YlTatuCph1bTaWSvG/H8iPp1ev5
bH02hKTH4saahPe+hVzDZ+LdkFzh/Ke7BJSiLfFDjrz7b3oET9C074Z+IVA0590a
qqLVEDeddT7RvE7TJh9pxvA4x5dC/ttLunp95j54LcG8Vu2Y1HuCTh03cb12+4Ad
oy2iM25JkfIQwd9sxMuHeMbe/wbiCeoZANnKIerx+EMZZjZBbHK01v8DyLkpc+uO
r7QGMlaUQ3BjLV/8ACA4Pb3/i2dAz0exUF/b56SKMlOKeR3OpxnB4yNLi2k2u5Gh
Ieq+xSDLOK0LVz20OM+fglEndJsTmv7i7IbeyXfYoL8YHtFQcTSt9yYblq/OQ6VF
egX9R7aBZCAOKAeC7giZ0lidrj9z++QOaMHuAR34OPSTZbNWTE785Lrd+ShLLCPF
BYVK9r3gtCvii+YAqxLB6lb8LBjsBHwlbvBgW4i/abNomkBXL6XTt7DTL5x7AVAi
6Zz89+fZk8NehcpyYMdsRprFHWG9owWYvOkB0uJKlXeNePwS2advTrO63j0VQq61
/1JPu0sV/yM9+qwqXge8HO0OnW9jdQ1UwYXZOPuVIowqfXr3wKl9Vm43lLDoi1CO
nHOcu/pxvon30oLWqLK9B/5DVjE+XdXDlr2AdD1CD5oVH3yfW9HxSoi5ZAmHrrBl
I6Of5fQr0ruiTCWqhpWw5FGgSHPq4wSywYMrLXW6Pexf/RrTYeSaB06rCh0Ug07c
2axZW4NbDbbErhytK/oF/lYtTGRU4TJHzAuldhq86ml8trXYGADcRAdI7eEBGYhe
j/zbJ0KKRkLQqSEvQFJoWDlxQ6XFJQWm0MTj7cLNn5CAAXldqKz2o4jy28SPJpBr
/PntK/fe0LC6ZLYMytSZcQrPy1aL1rec5zemBBNJZUXA0cqpIXc45SavyQmEZ+mV
qyCZWZgOKjE7AxUknmsCTI9RL+SDCq5xvgfdzKF+w1g7NHFvNSupYIA6ub9hciWr
WNmOdjRQPEg7jf1lmn+ztnSnq/ltWIvbz+KJkYm+JYbcqxxi9q2mvFN6+uMZsAjw
55YCkrAhQhdXPKtMVXkdNz/N5HLFEjRBA+jMGb9T01B9BiY5melSpAeCKPUcyAMt
KotcB0w6tzRm8KWrkUPnCP1VE+BNYIXx5UB94dh5Dp57Odb9LkdC6PnQKttpz5cy
OScHByOL/7QNE8Z8aZcB0c03QklyugvXhURciCci+YuYbO7VjMCKiJVr72KgquOS
VPfvNttG1S4FgnibxmECrKGyko9+RUtPOpQO3J8A24Fzl7PpSQsBWUmjG1ZDXDLN
Oit6rJ8UoesLVuhj9YPpahJy0q1fhBvQKjRjjD7BvS2hS7RcJEs+myaS+QrD+hYK
MvwVRcMQ2vz1BjfamRI0+MibDa8rDjdpcrXW7NKR4FrnDKsziOoo7Uq/5GSGrkGt
zBMrrP7fdl+cJKVJcP94aRNnm2Zqt/riSBT53gqET9eiLUBF4OxJvv+TU/2fd0Qk
iR5ikt/dorop5VQ75Pc4at7j1AuOTcsWTgYKHXQHGgXHk4CuXH2AkLx/Zoz4J6Bx
kJxLYd03Oh1a8r55CDc9xQB/UJzNCRhtM5taf7BASchdqLrXE7SJpbqqO0xJot5/
mRd7a302VZygnnQQx8hQN1+qkE6yD/9ytcHNhLhn3/Ts4vdqM5+JJhwqMAKW8Myq
YF4DSIk6Ezzo3k4HJ7Jyj5znFWk5qzWHedosDYOZn9tcxbJoqjUGMB0HesC45BZ6
j/bAs+Uz48NZFI7bW53cig5/ZT/H5kzTqWs54Z2aITwZgZ/lrSr56tJAQFFEpbqE
wdJZxF00mIlmhcotVeV9xqD16+Kx+NBXh9cf1TXJLRhMmuxL0h9XmSdXlQtQslGO
DVrBNaOxGn3ltnvkK6tlToQwSaRMBxrXpjEPCVaan+UXFnptlD48TUyDU/z8bL4S
8SbHNKmi9JAyNBjzJTwithekOFCX0/TAsHgMhRC8lcsqPKD7f4sNb4yGG1oJ+tQd
a9Qca+4PABjf8ZEU9rpEI3o0XJzLEuqiqzaq+Kdd2Hx5GWPBSwG2kBHFhNBR6Wfa
0mcYYN1hnw50hkkdeVOuVc3jHrNhXpEuvGVJxB3YRzfJaC3kR8Y2J6dMitSJlrx8
DNv+womMVCSMDhm3V2ng5UxMbcTX+uVTXPYyUG3KHp2HtCcn7bPGmYqBT10sMIDE
fZjr8oUoCLxTngfB/0z0nRgVhSxZ5cAjAFsYzHh/+VGDpiUC2U+HBF3rZud5YEae
Prfr3Me//79SRrj2u+/WJG+u/lrpSNhs+JXTntpgMjxr9j+5jaJunPwF+lTkI/nz
xq4baIuxWuGYAN1+b7QsYl8st6Tve7Y1xRQJLPLQ8s0prKHq9uTZryiPXKF6BhlZ
B64NCkCUrYuGURMhYBF/bq7S06zXSiTUUzGDTGkEHV3xn8KOkrJErSxkU0rNaK/t
lbVB8841J4fRChNNzE4ce93M1VVXFIkIZ3t7csRXciPfVv4mlvQYsNZdHOojOxV8
VIrYaLQYFQuvpDNc+lElEPTZeY/dm65ujquBYNPdsJHklBWlYh0QguEf990K/Xbw
ZFmGgLr0ikZPYOXwpsnziZg9TmqyT5ebZspbt3hLdAKYJ43401IE+8jCZwE0J8pK
mZwy8o/cLDwWYtPScR9l9zY01GnJkDTQ07FGYBbJBExe/GLcVI+4cKaB1A2Guz9l
UXA3aDGrq8fJkOTV7fmu7J/PNFTsDxuE/0VjMwiDrrNv4aaPn7+XxgTokDLExXVb
/Pc1mSz5z+8+LNETG8ecAAFu+43PUaCKomeHIu5zYlGRwPYRHeJhmLb74wGVhm93
s08LLoVbF+yF4Ic0vLkSIAtFrZ2WQpTvz1D7TrZ0wpX2TMQtfJpxm+kLRrb01cZe
Kw/f8b9vuMFmFcDoGqeZXOrbJ12BiSGZPRv+AMvaOvJBkHT9RPbpNmPX7O3TIStb
p+VNNKU9OngyXqWOUuf4g8x/KGABqkCyqUbDhyLk4/FGXg/+CqCS/hTRu2u1xwFu
1ut8Ksme4OZy26oEUn7nC6d78CypyB3D8gVespYGN4Iqi3Fx1UllHlbmgGRj+Iib
7dof9S7ItHTK6KnKfhSQkB7ssl1XrLCgwCJuXJfrzS4y9xj+zqGGwAxGZGF2UxGm
HiY8x+mV4vOc4Od7knTpKuYLlLnlh/gygKpnl0001/Yvqt/CrDkWUroLJT5NqRxU
bdj2BEsVyMYj9PGCil79oN69CE634XQEpJlVPCBv6RySAQA3amLn9pMZ6NEg7GYH
wL4bUNdMq+vVB7Y9PizseSxzvwECWIeDFcr6oQQ/yfgqo13cteSiupittdeQLuSs
by3TyPj+vu2xuxR6B63IK/uNnF6a6T+DeG/+nHXXqH34Hnpauvqak1EUfibXIA6r
i7KFa6421ru0LazqGwU7f6KwU6XMLXOtYd5Zh+p2MKG/rBbc1Cp2GlM8lTPcT/92
sjqluh1IXbwnpeLGE/A9tiqcsUU1FRdj7kf5Wc17x9TtsWqWvnXydTx/jYT8DivC
bSOSkkhFNgsf3/J/Gr/e4Nq3pbmuIapNBp/JW1UDBXPQpG9+y0E+dznsm5zLtAn+
Av6/CCG+iK6w6K8duXD3hjFOWlfu8GDWQG+0OS3bbOuC8hX23NkjXts7tz+xq9IQ
m5AAl6Lgd1ZO3+ei3ubzjnZ1/qmKV7kVwXXoqfP/BZV52Qo6QEEeSONLb/4hirIg
eJxVxXUiofwUPkkL99XzHsAcfXu/AHYClJZ+7ZmjxNCkMMOUsFD4si+2tsccbaf6
B5Vbk2ggzVAE6to/3NouVYA5hlNpNB/WPeIn/Svkk3w/EeyTtqmLA3NbxjcUVrl8
4kxkw7i7v9ck4dXpYMDBaT0qQSP+g+GA6Txni0Li8Ih62SsB9EWv9s4pQ0SAC4BP
1M6bCN1AGGR2/i+0zxRF0ScGB20a5p8BU629sp8lD6qEAk0opukVs4sFC0uHiz1X
Xlkc4MWl+YsyYh4Er/kUX7cxBTE9AU7Es5quda8f1sIB4dfTtgpbLAIa2L6KTPD3
TpY9aRZ21sJA5fjkH8TzpOAOw//8MbCK6GbH+Olb7Wv5y4Ig8Jisntq/03u0+uQf
MrC6uHyjEIcX/Tj14iFCzhL7HAwhBZW/8lNCsHslr/Iw607wWvRhmTqELqjFmaZU
cDBdzUjhCfzFm5jUMMCzYTURc63zzXiW1SEk1+hq47aE94mGzuTm9f4NNOii3LkZ
zA8Q9Y9JzYn6KEs7HTO2fQaeHVOW/1xpjoQH8/U+crsfBcWZ3CEvBI27PT8QlfQ7
ac9XqguLcc1WteG5cHCY3FYguSkhlDRoH+cZBk19MZg2roVtWd5pc+88q8crzM+v
C/3Wj+DC16SQNg+XXWjiRFKlclIIfYFS9sgl2hB5ue4VWTC2VKDjQsbs+HAEMRhg
n3fJu1Kucq/I5wwV57nRUBATYcJR5II8xCZdL0K/ZhyJzHgC+ip3mVr1K8r2Eu1t
wQ97PPCMYaN8BQhs8awks4pgTu8VtfLF1pMyZ59b3CJUOkFL8dvDacoeXKOTt2Pl
P/OgTy8qnSHgK79PI3n4qVoXwZ8n9CzESofy4Ym5bLNmIW3HVjfv3xm3oA7y0Uvp
eBqF2YPWAy17Vd2aWsKNxNywJFHQdhbdF8KaJ01xe5rf2QF/+22wasOyqGFWqFwo
7ToqKGfiX/0knpRear7dHdl2lOyLrMbZJdzjAo6zJCFnJcUaJpEbSSJM3PMtgGYx
84vo91Ga845y7ygVTDX/jqeKJUKlc2g7lS02qqiGSVfWx86+IdacW1TUkva+bX4u
C1s3QQW7muSlSzOJ8IRzTlMQVTJYJLEPLr4p2nRRbxEGEyhYyqWQQJNI25C3fSLf
+BBLJeqyspnhCwexiAaBq4MZIzk5B6Vn4tJnK+UPiWbFHjXsullAupkNUj6Uy4eZ
4wojxhPtvHyehZyTDgZB2eIYCWLHgHrxQWLnIGhIlb6EmSh26tHGEbTl+S5RJfwy
FSOQUPGTJtsoO3cfk8F1j0AdSCV7kgWtDW97KZpe+sSicGGGphQRTPcu2yb80QWn
cnP9NVLR6z5RmqiChhP8ETZYdIsn7/eOLJ/q+X9KPD6a5TYU1SWPO4XjkSHzZ3pC
4wIB1naMvFKrYzPNWDy4rCSVSxUIxnbiZdH75wAoeoC3iSOqwknTnrXPO999A2C6
odEEMe+mG5+6ZrSAVe+TZYM4RVbBdKHcxSBadkAqoumnbT2DJdCl/lWAPztd8VzA
wzsMNHfxg5OVUBhIg86kJ1rkdJ7pv3h9n2N2jgx5eCt0QpmIuVz2mYFk56xLVCK4
3S5rOHush+BgYPXKNZHdeVSPWKZEmMElctt1TjXzIrw6srqNvp24/65PM06tRELe
47aE+ZTEjTbzFuCa6vbmtZ6HW+Dp42v3MenGhZgHb9cerRGoPld2M+C08IRkymAL
txwVAI6zw/Llq6T5PMc/oQHfhy/U7T6EeflaksiYYgDY67wy4xEgd0ynaNsfva1b
X5GZxiUSFlmmqPtHwjkoqAK8hzHtee+sJ4yLbgheiWRvH6JuVjvwYAvAhKdxq+pp
nfwYbuh1dvbfZ8at6Trg8AAY9NgLCddBM/fPWLseGEpFb55Oc5OJk1AJkBHN5iQo
a9fhYLdskYYxI+KPWN+rSjRDvg3790Dev+xapgWCIdM+fAQAQpj4/RlWLq3Fgig8
85JahjRA4SCPy745OSfDPPLhMmWJcsgNsohcq7mDR2+9zZ5y+FNHtBFTGuSwOFp2
xmlHygT7eHN+HH6pnNpvJ/+rREqr+IKP9bMfpS8l8sDDPrhgBhDUJXT5afC+eYaU
aRd8IVVxXGn/h7QZNPUOKnfzKFMzrurfclU19GDDd6UIq4N2Bs1HcudpHEMqaZEX
/ZpYCe7Y8501On2npjzO0+w84RHoHZe7NRIaAVxoMfXbc9ii2ZBKnIFJ0WyPxpSB
oR8TFl/DmDLJbAsiAcV5iO7IG+/qFXFo3ZZKvdpfYysGmk/fyJOnyNHu7Py5403Y
an46lVp6QDtyUJB5NOjayRrpoaPd1zODJNMdMEWowhJbsBgc3s/U9I76j26OXs5Y
vwPrahimmR1hRroGtivgGgtC4P77cMJE2EcAGb+mmDa8AWGwytA7GvVfXapZGIYj
rlAOf1QFi2gndK09rO5mTSoo9mnxM7eteImUMOQV5gh8UHH2Y+wxhVrDNPDIXUNf
ICeqNw32grfeTnCryZXGIHocxLOOJvu+2ynpmMHJVyzL2AvY+bA6Dz8BgTiYVDmI
TJAKiE8PGppp5Eu056ju2m6ja3RvrBrBT7rXgUS0ePMKTxOoNcNEKpa59MFFao5l
0Prke3QE4D9XxUmYYt0HGe1x6jHIpFyeO5/WYbhVI3XQwf6ihaGdjAYE9TETcUIm
hNfhdL2WhKJGSJVIeOZA3IJH61us7ZoK1BCjI1+egpfI9WR4gW9otOUUyz2tDV+T
5GU2qPc/NjMEGZhK449TlcR+EEE0NMF6QrVJ3slZeMPJHxdoNomXIX3nXrS2EGR7
AlrybBdQDfbUSS5nEh5Wu849ozSlPxRycMo/WOR43yeiBrrcshjxQA/sG+SUdheG
HnuNfsRO1xw6vRY6isubVZ4oeSAlvyEFhLPvbKNHoIkVpTmlssAZoOMDlJ9nJHj7
9DnxBe+Ld1AY8m7MAj4HqUcmvOdRstOAy+5E1/LUvc/uxx9OAswSP85etEyTroDE
JJtG1PyypFkmou7ijBlMVY0QErS9o+0N8SVmuu2mziChhfSNqTrlTtzfGxHGGguQ
YCguRGNBnWb8+JS1nWLxozKB+0kkrWldcJica+Inb7e/T/MySrk7Z8BT1D4Tq+HY
9xqEg/Pha0jqws5fL+xdgggYq0joAk/TIJcXNEu3YhyuiWY1RjQqCUgjW3zHHWEZ
0D/JTq5XU7bqqyH1FHKIJASR7KP+6jiBkOmjLmxvsVeQOUceelEtSz1wX3afUF7E
jQfS4recaLthZR78wCZwXB4Awf0OV2sdhj7t7ioVUBnIIeNUD7ZQHC+TRDns+bxH
IiML2M8/gxQfKr1SN3zB0bW0/J6UmNtg3y/eEm5KtLBQpF+4vUAmpeyeF5k9+zJj
8xALlNM0UC2nHjUe/e2TQHXtr1ussjO9i+jKXaW+j3WNKHWS3DrXbp6IQZbjaLJK
k8KIo0OwUZ3tnzjoLCeVc9v3GenO0j2xz67MHY/OCH1PPAP7bw6vQ5LUhfSTKckg
lv1zsbiVJpHScGclE74Zd0ZbHHVo8KV3sU0SXxJLI4+MFzc5bbPV5abwTHY8WN7r
n8P7BefulaavwoPpkjUc2UDI5r/cD49S61AegElH9PHaJSevPwB4BR2hNLGsjiAy
weeUTVyaHEiMQ5wXj0xdlt7QhWtBahu+IdDm3s2NDk/T7Yqnzo5KLGQJCzaaiqRZ
ha9UONaVDPHBlsmLDPpMmFt80oyTUMTbdYJt6pDrzd5vEvSUDS85ynRnODZUv0jK
unv6bU8m7ZEjEQflcRDyiMAn3tRWuP21ZQh5+yF1tL+gyKphx8z7e6IddtA3iBSi
ZEZyUPubk1AozR9FD+FIYHh+vrsHyC02cA2PBIK+KqwJLWXgmxwcUdY0KO2qEYfA
YPN4d1mxBMpDAemGTH5H9uQ898QNKZ+TIDQ4vr/UYJnR1PJuzcFo4CigQJ+WeIpk
W9dIKC6BOz7wCZWkMYHSNJsawarMjzvfxp2b5dOzAjOHnUcGenvvs67I0jyKwtVr
JJbkEF4HYSY0UoRKPjzQg25EDpSEJxaWF1FqjiAdZphYHNYNWh81tRO17W+P1U0z
+KlhBH7xHjSOj9CGAtAL/zHDP7xB1d9rAuN+I3Qd6QlIm9NqhvcVdelHebBdOEC7
10wZ8jC/MSo8pNzRqeOmTbgvltHrq7ni5J+PjawmJng4tNZ6tUPxw8CH3XQHRFz0
o2dIeyq87ONUFpEOMdaLRcYK0P4EUh6OgyLCyCkmkXCXkMx3O7v2N2PDLXoP/eS2
8tHOUAWAVGD3OcfwVxvxvp9m9kv8Rji0rJHuBT9NztO71+UycRyUmqlvsURCmuWQ
whKQzFnX03znInDMrNWxq0Cmhrl+FnBLSfg4MU0PrG2W/lxI1cwdaFwNzW63hegS
peV1ZGSB3+15RDBqOkByMNnyS0d+sACy78RDQx6lG9wiCgdUgkTKj7tj9qEW0J5v
UQNZDK54LJuvZL764x6xdMaMCvdMtS9kJwXKWvJSjAHPbJUtVrUYrQEdGG6RSUyZ
fCO1L8lJz0bh9SzkOvuPjD1RDFknk175SyIwZlwBQTvCgJEG7sUI+EYqCB0MuSs3
lxs5K2cK1QKT3JSMRdQk1FypPe6shG0vOPm5uM5IYU+0+Zlu9GYBDUkfZcU6rgcc
HkqMEWH8dKCewVwCFmFtmDZ/a0Co6CoyzUa18bDBK3h+nhOPcgTtCsdJ+IgetiXT
eQNi1bKJZ5HZ8v17rPR28dDtcXslR+N+aEHvUJtQqCDxVbacjFQf9AZrRZuwhOmt
Wre1MT9NNwIUtSQ044ahYPqCEPU1Bddl9/vQPD74G4sD6mo7o746TMdKabf1lWka
rcyLUFC9Au9Op5G4zbEP74i70HcDdf/uqSzDFGjgrzxIaBjq5+pMvY1zCSlsVjMN
5K+kFMt+Mgyi01iB5rRgDjDhfFt9+Ib5tvyycqWts1++1R2qwk+bjXHGNCipYwTS
2PUcGOqcCehOXPPNRW4iFpRX6llt3V/uE0XQsuFKvhm327Kg62VbaQq2p2Boc2QT
HNe9O4ecDztpaqntC2ZeuoPZbIW/W0VjVioKZeAkUkIRes7o5yYRmjXjW1w1oqx/
FpXrLu8/afCi8BWGXACs14JbveFNzNMYWacMDq6pvKXnjLvcv+0gBxCyqvXpTUJv
/MzKjfAFIijCIthQ0LhJriNtVfm7gx3H7qzS1VOQODUblwjicpI/FJh3w6glBt7C
2AVWkxWev5GtWfWNNYHKwaM9A7f3mfirbPZT8QRsy0MY9cQBNvDxrhAeE5WvMQM0
ezsqh9j23p9/f4XEDiMx7R9Mhly4Iq+mNoAFpmUrbR386xwQI6ZAnC8D1bmgjqpX
EWSXcIRDBWuWCd4aJ3od9j6mX6x05UPi4J42jLt3jrkYNCncpOAAs20PkzJb3i1n
vPrBvpjL6x+h2EA+VaFwAtBmhPETf82iVrQMghIA2T/dAT3Zd7jHNQ4Emcq0sj55
jF6g/mDI/CVuCs/d0uuSORUaPr18j8iiK/Yo/k08/WOoj8+y+sfGhou97UOqDV1w
WgVvmHB82vGxN2E98WlIb8VsbkKPzNA0VLVuN8JdxoaPqwqOFPHLT6xg3UfyAdux
1+lu8GAMULxOFDEES2wlQxubwBzhJuN6QMMsOKceE4TpeLnmS8R8SAy4yQvq6o8B
Nbjuu7Y6juBKv2TCJxTVhquY1OjelZNcHZcij3ET8alPwPKlrz5AhdGOAO9HmMaf
Br/X+CieQJq11LNtHjNUZrgvaH9FR5PNwMrjPTHEqTlQ4fABNGiZNJ6Zefzk+PMC
xQZMvEun1fX15NhDwyOPT7YIsCwc4fPA0vL5UKY0uMUFFHo/q7fedbV5SKaSgvjc
95Vywx0nffZIlkXFVjCD2h+fgh4i1dfJuQ0EBUeIXQ0a81Qe3rogNobp6bPNiXNO
ZqInFFoW9j+1rjExLuLYkdk+mBedttmuuIYlxoobpH2ifpVQULFw2N2XHRUL1I3k
9dZKKCInF0FlJ+rOivdzvcnD7wQoDy73HLHvyRcWFN2l8LwRE/iowyfGlBvivxsz
StcZTRp7gDbsNZSygi0mh/K15lGyG6iM6EoN8qmT1FMfNFfC+EgElEihEJK9AxPX
Sk0nlWTGb8ck3Cyp81ZQG2emC284SEGE0zoo/S0Tc97oVQiNZONLRX/M5rlGh/+p
5wI/hoVm4ED3Isc1T5kelDoWcWiCPz3c1hUMJMZZAPEiL+KVIBN6onN5jpcroyi7
lVt5BFrHf/zxEiIhvZdtKgGsq3jwdil8a3tcLoU6T89BepZUdmUxpOASqifj+0AU
nN4d33pdJD6I2RjkKLRxMG1wnIU/J3/HMaorRfnzPEYjOFRIO7IvFQfulWpICOd5
+ToSQ5JeVCQmE7H5vPqqOqMKUX8nd1MIOLoeVsoCGC4gPzwmitD/GOdEQt2mIOZh
9W+Zxybu6/rwvo++u4Kix/S83voFCrUmg/NeQSVnX/hb2aflURgj3nHNySKqDXt8
gOk5WVbiBuOXi5ngnrALqmhp5cJ/MRZTWXDPGO/LZ2emJC6aBm2Vb8ZMtJCg6p51
cyJ7ZBkvKGgjK2xDGxID57fubLEiEiuuGKyk+ScqybyRuTJEjFjKI3BWOVjSNekE
jg/ik/uGT3adEU0fCe0Ak7ksnHilqw2G6toZJAuDHjvbG8Pibr9u4LsEYZ5ktinV
72pKvyagsBOH9UDLc4SgrW32fqd+Ftw7IXLImS1tk8JUsPo41hcvZj36ko7hb8Qy
sQ+cmSBbvdlpz2SmkmFxUXklPFrMe+omQRss/iDevEjgu18wjvwTJWXkpj/BQqMJ
Ng1j1slTDxXPvsK2rnuycg6Uc6gCr5agteZnWL8UsiZaVg0tvDT0dAMkwmMpYPrd
vfXPnl5pkrlFoIzeZxlCTvICuNaXNqyFNPUsyplScVhkTG3ioE6QhhpMoMLP9DXu
u00YB5w7+sCqaw41Yz5g06OnUpyfUQ/hhiZddt3ZwjUJ6R+gOrCW8hIXWculjvkC
c2EwrkC/Mj5yGZRCxCvQC5bhLfYu5lG/3BnDT/Yj1eXpOz+0E3C8xpCjpjY0CpSp
XNj1GNX9XxxovIBJwDWUqW5uq86VsfwoOR7Fa8iylIhe16di+QHuCuwsozRZjk0P
iBJ91IDmtFtXV0M1B5DfPAFlsrKUkh6z4znXg+BLtrh4COiJX87oNfgHAJq7zqyQ
1NAA/gQr/YxLmnjH9jGe8Zeg2QxPc0G8f+pAXipFgUdSSL7X1DXJLHruBSDkrCOy
9iGar1m3EOcHRsNih+LxZ9+535CzmiOFJ1+gmUXWk2pwWUcp8YnMz26fk+38wreu
lhqkU3nBLeejOqNxPJ/TXOr8t0bx+U+2uXzD5S8bp2vEZV7MYkeAb1qHzVz8rowD
KjEasK46Ou91geR/xOkp6vcnbmffIbgrY+EauR29mUzJKC2EyRQbW8zM7GGeVMim
GVrP41BI5Vwb8cTWWHXBA3dLFvOTsaxp1+l/V94BZckzzVjxsozFTZmkoXavWV6N
TfzJTLOlxsW5myE/rKj1c9ArWD2GtBd+uNjyyhoCpJURjcNJW2ZJK0RnWvyHyR+W
vUlvIKQGQP4JL4rdEuQeJoyZc5cpdpmmQTaqCOz7sm1vURIyIenC+oClbtSkIgpO
ThOKA1xyMSl/HtFOVbPiVfCO2wVtmsKSbmH8Tk3PpcPtYsKUQ+TGu4HfmkEC+m+K
0l1/KZrghQUam0naZlG8vKAU/mx6gvjkER2cCdkUAfu5kCqe5Gau0mMNFc9smkFj
WzxWLa/bRIkDT1jVq0MVoHUi+xx1M47dtGs65bDdTIc3j7swLVcpzzDCFBAF5+IC
6qY57TUSN5dPTEgMkj/WzsVfrf1hYzaYYn+GF2UV0Un58r+e4QicQ6OVxSjRajet
x/oX6rgOkW8EpHKDMMw14rFlGGBn2unIwm4ZxSM2Hfo5Okptg4O2XjEkaFz+/SDq
ygOsseJ5XZacSVIxnXYUUJwpJsckwKJB+BsCvaJDHDvfoDRkLc5KKMrqIlud62tr
6k4R/eVsbTdrUI0yeL5AGHsiS0lIBMoMetzIVNKXZ398gqup7W6yjcWvfBlcSuLY
LzeD7zLj3rT7Sf/o2JdcPyKv+QWoc1oQ9GLBDvDSb2xYiBxcTOTK+gdM0LGeJQN2
JkyMAJpIezfyhOV6GrhfmURWzDOGjy+nqf6KIlMNELwuw2sa14m/HxWbEdh8Z+rQ
q76QHxN1NTLExGPxDOiibBFvwkB5h2nJr1fHsMJfqMpjpi8nmTF5nR8ojS0rQQlT
FaCpeeb/jqhLb2e0xSCqHG8SbQbCjFZht2Dth60nnYVI/weR5RkV4Av7GVWlbrvK
OLZrsLoWS7GvU++VrqFYrB2RVhxFRFzZSHiv30GxDqtbQTaQ4SUcZ8Gpje3kqCSJ
HF1uAXyTX/Njgvor5sx+mD9wAJGJIWdm12yfQ/Y7VRtwcYJdGb8ZkqMd8hWMMw5k
NJZrbPvTrSobskSR9YsK5hpTEw6p9F8SuKuGCvCNd48QMOWF9eR0Ryt3aSUKGlN4
yM29u5kaFf0JeWKqKMdlr+dhsHtpLh7BuR2xqp30176sLnA5Yv05HTB+uSIUUmpp
qEYncoC1qEf3sxc61F3A8Jr1NLK7fEqG5sJTnUNKnQBI1pKAzIJkfk8tr/6LBn5J
KHSdN70KyWj9wqKVLgpzKD17hmPNVzWCCgGv4yxMYsICgLbDrsZTPRNApTGzqd3l
JbzO5v0WZqbUJBCZUNPkjZIaqrJywpD19vGprl9RXHs/VYRXnBrvUmPd0fhbbxQl
Nf+IvpQr6TMpt+BkcbNiKMXnHQQ8R4fY8vMDzk+PVjHnsRjrTvV6pNXkPtwSqytQ
eiWy/xuC1Mp10Qkl+mOq6zbdySS0adEMnDbB5KdIkS2YVejA0z2TRR/VnPzCrSwk
Vxk0HzC7voz7IQbrjlMKLjDNUhNHxIQUNF04MvfYuFUSJlOQJBFuqtjWfrgBF4D5
YAu4Hag/m37x2bp5TiWFqep/UPDIlDK5uWykcCAVOM9Oapq29vPp7Fg87GZWEDIN
8uvVmHJ6K6oX6SXe0vLk0atZ/PdMiseqPIN9WJ5lEdFUvl3JQ8U6ks5ZhYfHPF5k
fRMO89bbsn1QZ4eCW1TvQUDhDqw+6hpeq+gcSW/NDufDnUnSwW9UAqtDqTQksWFl
2bXYEtxnGgOx5Khf29TAFvjYqryh4D31ERE27B6l/Veqcp8F/aiF9C7OpdvIiWD0
CkwCst6TFkpOkkqjbiMoGAi/b6ce2irEzygHN7xdHKyKY2A6YJu5BfW/7lPj/WUp
ilt+JsQN2Pf4AQEkx80dMx6vgnITFmuEhcJ2KUZxiYVvRBbu5ilOOd1w6zto9wr0
z7NY8zI1KXCxSF7mimo2Qe+hAtwsfyyLjoYGVgI6kor02rHepNPy59HgBVtqTL56
QPxwQIRHDbEoialHTgF6sTT0uCAglJ2aWbO47xS6+c5n50JBLa6UjVxznlVL3Aeb
ILEgzII4I3/TJ3QRYdtMjBSmKH4fNEJiFjDjb5w3Gw7zW9X/cKO/gM2/y5alwEGD
Hvhwi9OtNd8pZBWJtcVEGAfusvrYjIpsoMYeSrNR0Yflp8ytKwdDyblW14uB9t/r
bs9gbaN1/3B1zB4Tw0bNpuNU9Rgtjj+VeJq/YbUwG2IEqbpZDmNslw5pqLnVfkr0
MO0TQmqobhHA4Ers/FYI9WyNWTzaKDEV1akLKUodwyMOTN5c/ENa2mt42PXNF2xe
h6+mE+C79cnBFQxM5HhPvA0ztiluL+9JGDEPcwmGccyzuEy3pfFCxp+2i4heEWN8
PU0N5Qf7LL4l3wWmekCo988uyDB19O2z6Ti0S53vnusizg55hxA4zWAfHLzhZm3f
w9NBAqOecBJyNlxwCVip6+5p4ThUeF4fOxneB2VGyZX8lfUrzDLCMQh4E6x2UiEa
+8NbxBJI+ZzNNXz4KKZ0jjbHyvpIMD6/+DbL5tr6oGpIGwP3TmfoX2x0VMJlObD0
pfIv5FV5tjjg6GvhEr/WTbGzdsLh5kpGw9SpcFLeCChm+aBdZnWm8yVmRcpk+G6p
NLDaasqFCPu+/JY8/vCLRlnHoNSBbM013o29vC2BgeJDT+bflBaJWcJ//z6fUdY5
b+iR/iKSvsmv63RERZYN6OrpyF92h86XMTuyc33zveSikTs4iM89ng0lZxw4RiDV
9hQYeApmLZpTSD1tpgoVbqmSDLUB/Yl+OtuwJHhmTnawdNiHPBTjlxlfyP6VzJZo
Gr7zeq8gFz1e5gTbZc07g41c/VWicYmTw8hAUoGpSJF774cwh5ovkVsEBdNlTcHK
J3aSt5XLg2NcVQDhcU8vaolcZmSp7vVv54BhMyZvQkzlAZAx9oU13Z7ClZ8p2lW7
ODI9SXQUKERxFdEPTGgdGU/l3nOzIrGIOzWnMKIwXe896Kxpo4tIQUIxqoFjiC46
A9G7QLNAIwoU/LX4q7B9SgadS9oojxFFo7tC/h6o9t7oASABvjJ8zf6cvdcU730O
FG2kBIrKHWnBqnQTS5pFiGMMlK9oChgnWsWz+YjRYdTNtk40+UIh/aYE6aQl6NSr
n09PaAFTrGXabEeoqZeYJq0sKbDVvoncXUbam5TiqDwlEqsc3lK8qvxcLSj+EL+2
0KSIV6AwPOsSHP3JEthf704vrn34kglXaN9bLVucEKpgL4Vq8s1aSd6JgDNBKRjF
P8HroacGh5HxjHKk99g6dBnFvtR7Y9XFHsbEM1omQC38i7glD4oj/m9u3B9VylXN
zMcJX3f3XOjb//8Yo8bBris4sPSQnxRI6Esti4EcB1HWKv4Erpv72dMBJ/MLAyjH
IK59vaQAAjCy+lMXtM+a6ERc7IK50Tbkx9PTzmtjgzx4LbFsCDow+8e1wiuqxSqr
O64RrBLLyoDtJSsp+cjt38bYyH9Yw19lRK55y7MGvnsyB6DLW5aCWsU8k1g1RXwJ
d3wy6agzHgHmj9xnD/OlVUVNPR+orXePVaAeP4ZAYs6hDWWuhNwkJLE2rT/OWA9G
14UjQFSpsL2ydDK1DicbbG8c1GtFYNZqF/G4fCo7RlxwdSAlWPNzL5KvW7dtM4e/
iDdiSqTr+KbuhQnQLY/H6YX2QLEWzbu8B36gb1CfBy7czsX57rPetw9HQ5OQ7Kmx
MEPnkuBUs8zpPGxR5xTWMt9PwyofYRqwqvYOXUjSWn2+UYhgWioJ4CWLMp0Q9oy3
yVrbKX8gWKpIX7ev4lKktq6jvWTSL4NBLLnUKRPluNC4LG+mEnxjsj+FLIyzAe65
3mb0z6GqZoXaYU2nYOv+V5PQgu2egHzb5h83EN82AJooRGOcw6njbPO28JZypZnY
//rkjwtwbupvgV7FjpP/abbRmCmlcOUPNE3P4gV93d+vAHZLqEl/IGujs+wqz4j9
WdUAPHQPqhP6UXYZQi7SDYTdyWx1HPuV6AFkIFL1Eu2chv407vRMnT6q6d0g67ZL
imGAq0OQPbkEbXC/aCm4iaMLAIhBrRz8WACu3reJLRtBwv1GE6Lvs7/TQUjq15u3
Stf0jRXkFrNbg0sfc5vsSsA3HWM54lZtIXSd8wHH3b8EF5EkV2MvK8VMPSm68KOX
sDemui5tOBcXwYruRZupLbSMlzPrL9aU4ukWV4E7kkVGX0JCoIUV5FrjNRADUTlX
BNWHtancthLwQJawF6pfhu6ibhRCR4zu00+i9VgqKcI8uZoWKK+r/W4+iEFlDIx/
iG+6NYC3P07PWGnEvusEWy2BTHl4+mYD4Hr48yClZnTM2C0sVAlSnsqHjzuekh9i
T88wsGlWngvrxkCy16LLj5h7JO/brFvdV8xp5FOEswbz7biU6JDWJJmCXd4rfLDi
rZAdxnhbYS7aK26Xof1vp91eUgOlPNL4UpDCFxCGP5KjljrXmoAScZQzgeZhYK1d
VPm7Ml1jfXq6N0sylODoO8qCU6as9GurwVR5hf7hsDzWJI3n1+jzb6alEo6GDpdJ
VgsYm/xjHI/J4wmr6qZUz7C0T9a5Ac5ocnmbS2xVtdoyvPa7WP7GXr2B5OJ8BBCT
fOadOkgxpjztg2FKaZqdCaJYnuTa2hdfbY4bzTCDY4/oKyt945GLgFNWSxsujoZE
xHprD376M+6eR9NYStq4QuYlU6kJdFEQEd3VimT5jqsjoNhCDHUmQ80p6JS0DifK
kXBK1YFL/BRzzgIc9dVQeNGl61s0rPfnaHZWQ4YKks+Em3Bj310w8+GftQbuv5on
TlsJC1AV4Av+hF0WYLQxD4S0ECcciYqISinbKrcJKH+2w+yqo9ATw4FPlStzgGhs
fPnQ9mqjfHoj65I5f9uyejM779Bdii8C19kvQm0njy1pUJKpSbbhrEVCKYepH/C+
bXxjRySVk5wkK5r4IZoVKrs1WyYxC+OXKaPc4gyEporwqVGDRrcr2UpkxmvAK5t4
CsLJa+1wjdv8AgePjoovzL2GQA4aUrSytYv/pHd9Po7s+YnJP5dIrK2ZixXUCsb3
f5cf8m5sUvMIc53Eb57eUoLbUKTmPS2i4PxyHhYQonyiK4t8hmoU1ApYCdXwDcy0
WgGaIVHhUYfbmELkTHNMBzQQPTLhqVc3aJy2UdvdUVVi+uK8vkWRH4F2PUgCScVY
YXSN6WdY5AKgvF1qfzuHlszD65BzNkAeBPGin9Gsn8i4hpyE5YhN8mr8N3coju9/
24L9aiA+4cbdA6qWcmWciBjVth/KeFhCI7AEH7cWVY1f6NdItOLNM5+awm76Sc7F
tbjWgTl01YOTeRwRYsvhzzytrdBVO4+z5OrJlnGi8G3OFqnkHaQhypCq8v25W/Pm
pCtWM3S2yKuI7MF4+z70AZui26ou1nNnRAvktYBOQhMiyVSHfZsRz1byUmd89z5t
WIEZTLCMUY2LnrrfYUNDXvZ4/dWZIT6essXcLwjc+QVlh3g1NGvI0OakubPnMfF4
BFanll+xmq7pYKyxnLDWEhLjr05Gi1mCM/wCgXi+rI4rJi4GI1KIqwxdGZaV+rZw
sgTs7z7spscrrJ3xDsruQ9zz4hPdtcK0y8CR8v8PK4lNkutcouWRMAPDi+kyceHr
n+uLQ/94A/Do2ImZA+KVGe2KnFSGOJ2oFWK8lw13TJWSV/m8JXZeJpQr1wPEKLW+
3OmwlK1/xFTfZ3SxwO8oictKmdrmBk/l6gXV9AYqhtAcPZb8wWM0JAHyfpZ6QtPa
yHvW/M9fwlwje6xc7d4htneQrzbNPIRzMKBHD5xMIlEaMNhOKA0b1G2c8spS85t2
QPzXaAGu9s1Btqi5vxviSLNuYBHl3kys0c3igiFc3zh5zoYVpuCg7yHxAyz9BbHX
rYSVrgj9gFxPdy99atefShmqqMp5QJIP17CdyEQw/nZ7LpZlVBgchaGE7kwPMqdf
e3kArxv7xQcWbgY+LiLAffOKtCeB4czi/NaCIAfnhz9MdW04K7UBkOek1DMWk3y7
EMg0O6Dt7eFT2HBsQLjih0zQuKTfYCsR4kP2pUPHa1o/mQpfKeTt+b9xv2VWWXiN
4Lf4Oa1b9lfOHdRjA1kzOHgoQr+ydgyfrZEgw7qoGaaxx6R2jWGpq7R1slCH+GJr
1V1n2YFlKdt1Mq4zPR9Yt+H9k2wlcNgf54LIaoxn+W4rB8q+4GGbJJzFCXUjdeWW
gcYoOVXuQonkAZwm1AZE+uf0yVaneMxhN5wb2IVMzTRiyvQEBDF7nzdMGsl79jI1
xyLrRN50IIwfaq10VAmSqD6l0rhNDF9TpYwhzjXYRKu6umOPPzuKx6TMz3qfK0eO
ZPtKJZZnOOsYIBII5CGeirjUADJyvnttoyUU+qEnRPWjEaI6NIIs7A7Jv9EyT3+o
+giSpcdd3Bvv0GdPWsR0XdF2sRBvmiRvZVohE6iqH8LR6Xto+Ku7EyWu2hSjNcM1
KVkwXedfGi2tnhNXbYPfJUvtReYySfhtTLpJErofwo2QyReKE/AcqdCXw9CZxISQ
ziJf82xh6Xj1oxVZJ+zAvUJiJVLeG62lmHk/iYAyC8gM6HxH0Vrd020M+pqjq1a+
noDbXQmIxGYy4JAqebcZXO19rz4kcCcpf9aQQYj1y0moxNGinNa70hJXogR9V7H8
obl/DVrGg4Xp7HtqOz9tsYWNnq1cIKX3saYzA72j1eEbF6iT3UZxLXmBshvsE/IG
YbMehKGBT9PImtLdCMjGEtJ0dRhDarQrtaXALOub1qLFsbeNMHkF7YtuBLQLWGs/
f0qghBWauwX1FvIBIFpbzjjAwD/dIj98txoLe6X4TctjT5z68XRBJ9xjOwBwptoH
fKgrXPL6csJzb5odSovGowjoomfNYaiJgGqK1AFO4dNrmaE2GLDMWbIt5+NdgGrm
jJuJaR1lg7YvjcgzXwZtyKwCjsbiB9FbraI72o/NqeWIQrR5C2aeJ8/4Wr8NHRrc
BlR9IaOhQCBq0ig/Buod2UlEwFFeR1oApvb5QKHNNoBCWn5Y+qsaaRa0VJR5N5w1
S3uyC68b+ga1W8DQVfK+LAsRnEZEt1LeR8uvwpqxVwqB13hrVOiHuJPjTLdBNT0I
eUY2Od1581Piy6P4+otn+d1jL1gedIl2qsaouTuZKHjNZkfWJLNP+Xc2g626iBCC
ZWcoblahy4JWMZRjImLMeM2CiPpPO8msm9Hq/+tJGogW5iueFFTEg7Ql4mTbpx1H
gVXpEw6N6JXuMpsVv6cCrY+WZvj5P15yBdcPB2fFwRt254BuNPdIplZZF/kyK7vd
BgzSqUDoRxP5AE8PG3amh7btRMlvflY5MXmzdw4oMMj2VOgPKNfy3uZI+H6JzjIA
71JNQWghGmlTxHXqTRec/ZkSgIIPvenpy46CFo4hX0hQdAkXbI6yu9zOFoEH3uwI
pQRSdrUThYYG0glylKDYZGvYW/I+2SXkjGZ8j2fqUArvcNB3fbF5qxGpAxWH4vJG
nNGnYxjfP5bJy2fuUpOd2uBpqARmzZ8fGmH68I+kpxuSNds5qnR1/EqVkIuiTtuy
InrejMlhZvag6OWJ461+hBjKoFNbwgR+LQfqX2luAczhlchl6mVpmkmmpfy09YbU
52m5yRVA/9XXad022qyAC3jZ67fTJFDhzZdufUH5/MdBUZ87E71tloUZHh+yavKr
BXbNILDosfwMsoFGs0AMdk5zM58Y2DOa0XxHKOKCDA6L7hMYKhM4gqxb2X8XAJFf
fwDbovJpJobRt6phh8mzGreOjJsEUOMoW9eRvZ8Sso0u+d7sjzHs6ExX4EzjR6rv
z+JiWlQdbHoJaPti5rwp+Y/JwTXNbyMaTP8GL2H0gHPtfdlyQcxj/J6AASLoNvig
bcDNPNunwjpZ9q7IorzxaAhhm5Jiv347jx+ohkzK39veMcQq3vUlvRis/3S5JFMJ
0nx7A4fSSk07ELAStI7aagDWCFMgEaXzEeM6Q4SGORRCZdiQGmWPuYkZjkozg9bm
tAWsPUkWZ9Rhaidutfzwz2rufcXaGTtTpjgCvRZ+mhtPDKIP7jyof1r80ONWcstO
TfNd9irEjKupxeQEgmAE0L8O8sFHVNHCl0ZpqqYPmrBGDNdr7x9+6xMBfN/crp3V
aVqEll/nQs+59Wu+CmK3L21TzJW4b79wq3Wwcxzuf5QRP1pH3+UfWIHElKpFhfVz
LPSFJPVoE0Bcu/rA6gRFMIXXWQMfUbbkArs4Hsxf9Jleemqzgx73O0LD2jrMPuFl
hKLQIx8Fk9+HTB7R5AjR5rUuyetBisZwALEK4cEgs3WzOoVjpMEYoYKTq6MkTEfU
Yg+ccWrfliInz2L2+ItiXYaHk5XKikW/rlI6NW/5Tt2/jI3FyzB5hly8MliZzgIt
8JAZsy5CS9szfPXTzpQqEsQ/Xe0x4CujfWlEA7EY5/legpKf+iiABNVZA1h7L36y
dvJHTQ7P5O2kJd9i8G39OeiWfTmB8vR9YCKyeasXSabTf76JJHuhAWymK6jD6gOi
+0uMenGfMy3PsUOg2YtYzwd9lD5wMwINWasUtSrZQRZlXXNPqf5hMe+My7yY9Xxl
virqBoneDDWsBA4LkUp7uh3X4AvuyaghQFGZ5wGaDKrd6S3ui1rZG3Z0J6OweRcl
TKEdDQHz826p3OvedJgLJjv+wqqrG+fhNzou0cAwQREZPjBHYn8JFfN/JqRWVVMN
AdYqV8Ceh+IQvDpNOxjGKetr61XWHcAKic3z3K8gSjh84s4tHyzWE22sBJ42J6/Z
4GOqhT84xfy/n1A5qlmG/XCyVXg3HL74SMQVFJw8VJfKGEji1rFLczqYhEHFRh4F
1GxTE3M+3y/nUBqZFqhLp3dYt52N4OkjGTK+Okyifz9VFiwzvxYYzY02l/KchQNH
nsPZBVecdQ+YcpMf9X4MHzBjBISrSFKLxbRjNLPISmbZVAKu8Pe522r+Zxqf3qc3
2uigUmnaQe3mE02a9z5Xnm5+VhGWGCxRsxikcS5XhGE64coOMuoWxQaCexqtJ47P
t2khgloYx3x4VKTTzwNm1LQE3ATVllD5xRNflWZzZRed9aYEywE1P9fim2hyDD/R
zgkEILHGyiMDEQSj1C3e0HLbii4YVU9ixDNzLcglnGd0QYI8a4P/S8ZJxE+2zlk3
rM4ipWhFaunTlyxpsmAnjGgodmbBPk+B60ORsl5EZ+3cR7teBfedIlv80wxu8PM0
JnaH5hY1PhelMnm6ndevzhvL4ovaGtOeh/QcBSNkAl97ciChvHQfgEHzLYCv/H8h
zchKYzfpISV+YiqrSrAnAChD+X48SKho3Gw9nrsGXfNSmAbiQSL2M12SnSSmUMxD
KrW4zDvr1A4zzwuAR60NmDhmMfeSubuKTd8gCaC3kXcc0+HKaKLS7NPMT9sNwlRS
XOcGC/MmM5c5iRHnOX81/lR1SFdRupHu5xkwhYgy9GQ0Xq2nj+dVt29+u8t1UuJC
SMwbYUWvKXkhs12de8htHlszaHk+JgXZPrslMLuF8qRmWp/BHLlFhjhb/KKQT8qO
Gt0zM0+Tq3cLZTYe3slR6smKxZZplU61U3bhzMNrw8+g7oTB8HUt44j7LutPvIsT
AQNTKpjeAI0LlIVKOGEVOvCkYJEUvXKRTZ9oKlSNVM/wpEw7kM94pplErBKBeBaO
A11PT39WqYS8O9eRo9hLRa6LIp/8QlUi0u3TQzIQR8p+WMu0AOkf0m+ghkkpjC65
vHIXLdqi6h4QC5Hc2b76aM6SnJ96CZaumZrbIr9x8WXjtDBmXl9OG3cD55fmp/RR
D3iWkbVjZhbgaWbLdTG/I6r9JHLHBg8y7XqylAIxfWQrpuWqMl1teMX4PolFk/+8
Jayzr+K+hsrtj2PinzAr4qMI29nWlKak5aCiGS69XF32Q13UTr7R/NG1B+f+0UVX
eQejRwZwjZu/PQvdwPpegwB2KUCrEpkmK9vMP3XBOv6tLYm2/vaUR9JYkHY1+MsE
0JDfWScuFouGpu1QYCwx6/g7YnGMh3EHmHkh1YiBu1dFdhRudmfF03fb/aL5NPlW
14lEHE/1+VOibvVLup2yJtWikqxY4ILFcaWh8WAiu+kwsr+8UAQV47hhvuprZHVM
sZDJnyTV0E46lz3GpP9vOiHMCSo0TA50nfRLBpj9oJ3ywOcd8ZVjoQh7rCn5EfpT
IFTpCNRQO8kH2LDwshPBn0Me/gNiYxNNc2KTSuK+HugSej6P/WdQc0niQYHkland
x1XfVXN6sBv7IPXfRFNpOWO72mfw3BxkUEJ5mqzaUQ0LgQ+Ussxf1VsyfiUN1PXQ
pF9mFQQejKeBucOk2OLnBoAGEaZk2hw0Yx8Z9W2xPijOpyVrIuKKncxWDopuGln9
RDHCkuHEPBFYoGG4JrNDhJQWitjODRz/FskqFV3Ou+0uh33IbZWWspDQ5DQURfgG
2Wa/XksZeloEa6Lfahgx7KH2OXn/HMt05vs1mHvL5Ejc5L1jeUt3k1EtnEjudMM5
RderFkjiQNir9ZL7sZ5ndOTrPl0OkNi9NWIhKbJQa0NP+oEkHOY7089qWA6y7Gxf
xx7R7Wzg9ojrKXhjT4L4xcyp6m+EeX7PDSvxumkL5cYz2/qsyzQfq4ZiyKIQFmQk
P7lYhXCuFM8gkJYxLltX3yLcMbA3DWTb35aJv/DsmWWdWixck2jJpuE6MCzeKxkC
cKmawLZrxiuXkl+A3ecmUpnHpE+Ri6RUfUuO4jFbu8qzUH+utjJGf8XKEdwv7fMb
8ceGhBl1fMW0fPwM/3qvxxo680Ec53DpkIMeEPqkgTQeK26X10hJHbM9eKPgU35x
074yEoCQGZAA2NDhXL8Vch5mNPemN3+0dLirFwjF1U2c8gAB+8DNzUM4t4MCndSU
KbJqNDlRlGcAEaVy+zs0hetcRpw08NPVRpytjC6AjYs8gK2kJPMOzpxyzsHcryjL
KYtdS2IvZSDqFfqyz0T1lr1vYU4Sy1zWzunBZS6Adk1HpbfrEOBGurCJ008DrRRJ
up+sGbwyolPp4ePilzQuN9x7/dm22CVuNCviI33donW4ITcve8tL1HKH/0LrGulU
5DCQRJHKhgUqentDoS/sCuxOO9ySwDQLKKiYsJRN8FakHPS6HgtDwZu54dY6RXWT
1Nv7K8Es0OpL1e2KBWmqbq5YvraVd9wP6jTLZ6a79GpYVHZDZ+CPeLrKihCJkM9m
WYX0NPel4PtFC6VDOhKcoax/vFVQEQ2zTfEO1lopN0Z6V4q/jVHrwORa60QHZje4
tcu+ZSSmmEeua6z13KpvXOvSDdVR+f3ql9QBc2OmXc0zAbp1o/Dxko3HxXD0jxRu
PVaXNgDSML1J1hRl0LUmf5ySdbPwDifkJueeBiDFBaHt520SwdosxJS4pnD6bVy2
ghCo+dzkALw6JZlc/KKqq9LwPoKx2YUGAOPErLKDYkE6m7qgu3e+jg2voFiOs1+o
4M7kM+qIHFqrLs9pSYyBGLFQBY+ld8v8VnYWooER+wdV6jU5SdOIiwEfWsNOsRZe
7I6c3kcySkih0ug1wWS35LTweAkYhXzrg4YV6Qm+w3QUbSRCje14o73qi5I7JnwL
Kg3r4Br7WczOua/7bwDpXgayZvy6hnAgJOLqj0+gGvNLWPaw7bdUz0Dc5DUVikUo
slbBF0rMo0dOVMNtNR8VA3kA8rJma08Nr95sGDsC5hE1hhRiig2G8iUUm7M2Q7zh
FNaBDu0yXFEHETo1ThFZlSGxwFQraVTBjsGsjDUx3E06oI0gtsDRNNhUBjtHLjWQ
sXdrOYQ2QrVl70KigcVD+5NlfNzsRZ/X5cYgfpgwHSKvFYldwK4gZ/LDIR7iAIPN
Y7J9uQYIJaQUqPjLXa5s0pa0cI/ki1Nfxu/YzoPn1VXH5rBCP2ED0R45B/lrMidA
f73cN9g1CulmxbfLOpazw9agjac0h0x+vmDDyj2tFAKB6CqoOznGiEhc9UrZff4v
O3+gu9qvBk8yeVopc3+zogR/KJDzV0b+9gUt0s+dGmiSn/OYJxY0oDUh59/Gvteo
w38UC0ozaWERba/l06fKiNGwMXgUvHnPS0y81tQJhwSc5inq0G64fgYo8Oic9mQF
KHsP88SrOAomXjAUF3SsultNGwx3xMNH/8MON5kqMWndJP+urGu1EFq+V0Zs+fic
OiEMqHiBtpqD3V1IAQWIRzrgSE30xPFjeW5XYJLzMGrOf1ZBK4w9LbPPBV8XDQUr
ZWTzhijlYWhmRY60OhDw/chtoO9NkjgonjOqYnPXazimwiRtp1YLVPg0Ndo0aUh/
Skl2NFqcR/xykNkTSFWfWJpWsyNqNNXYKV9GETB0Te9ljOM7kZLK/71ADWMmIds+
ljKzNcWVHY3x0hVHOotykV7HvsP+sR8D5dL4lsKYUfqqt7vJuqquo+qh3ViZok+i
GfqqQHKt/lRlabExrex8qLkErI4Jwd4BptXDCAfsOr7Lak9QOkgMfnrqZGK2qEuz
yrYVM/e8Bb35ccEehd7FhKk4+B9uzmlSQsoIveXOF2PA08DdNwvVTaVYfFcarJI2
yR/UjVgEuj4ohMrCU3UDH2icKF4kohiLpDdYxrJqOBe0pPt8t0YQhr9MvHj3M6k/
H7j9H+lr4CnFqaOdcXBXi1gwrlstB3kEiDPQO1QvJDYIV4WRTngeyaYakECuQ+fB
5/lTk83p0VgfJxOB3+zPkdANrm8TG1IgBf71ffHM3+BMwirN+NS5JmFWmIquXsbl
pIZOqcl7PPCbNML6cJuQYRR0rH9clF44B2iiGIpVOaxL86F6I5dbAAepIgHqHL0S
3sMsF/JaXLPl+NR6OXyksa5A3+c+efXv5Q2LXYQ4SgFRKLQnQMO/sizP/xHQfX45
jnEhGL2xnMHKrZ6tI6Kt/e57cf876HKa24wzqtArMfeMMX6wkBW74LvhN4PN48gG
VLVpr5ni6gd1jY3yG+UAmQbZxk/mWIiNXbI+sWiUFzFdfHp66vRKuembvY+RXgCI
PC+6CFcRJghJSjFKPRspirbBJxGY9CD3qy6SL9pnYNuneO6QnO65FQs3qJjO6MHV
kXUENTB9YTO0VwjgG56Va3IAfVsiEUbcYNgRQNsfbxy6I0jxNB1q2aWi08yQqRp7
tzElp+ce4+fqaPiIIR2TJ+JzVrHMHEsjen2WVSvv4GI/47uxSyyImgdeCrT7qla1
mr9sXdLJdL4MmTZ8WTOB9tOB4HZrO67cRxZ0Ev6vVJrjFGjN94in6ecarZgwjIeH
ee6oxntG0ZPjUGTGQzyuNzWLNLTR4lG/WxQ1pijvPXwGOe8LUVSyvZrJn1q8Dq0K
tKLca4KUheKPuoS2/wrBf+zsR77MLOV/kuPhMWUmOzN7fN6kuOjWmC8Op/F/sUwZ
LYLZ2WtEXlHZBAwFjuztRT5/Hx7ndRZrh9sH2LuTyeTX/BNPILknjS6Tvyb4GCr5
6+ufBvtSd79ByYg75eVrhKue+euOwJyJI1Sq0nYYXkv1Gzc9KecuWekjj9EvS1Jf
Le3qEBdO7YclSwmHrRdg1yfG37/jtBjYWnNnIzemMLh6HWwu2WVEROUnfoPfWiYJ
UTlkHpKQGJhbRnrJdMR7uXOSAMTKNHPRYYiiiRtVNTFkDfBnddoqqm7NnYqfikCB
O5NhuA/5rzzFxtltfZAaMtoz2RGsMjYduefkyk99J30ltPiSWatspvitIf5Owvtj
c1JjRlF93hbPwwxbqUYjYWe91p1p8HW8YgpmPCU1VVD9sthPvziTJ3Z/9q6Olgyq
0XkjPc6fTev3c8YxdRY4cp00WTuLwavNUQONrG6cWtaVO0nx1Q+Ru01G74vNAFNB
FbHGQ3761Md+xA4L+5tggLTCTCnt9Otdcb8EVP82BBaFoiPZnseh0NXc/il1sEZY
3E6C/mmb/e28AuVWFfHIxJTXLN10K4/HH4evcxAd3+qZ+oEYZpgeZEVU1LJJYmcq
WRuGer1WjVghX81fcCpm4z4aB4BaftQdVtL8KuFJYA8monKB5/EERxFA5gZPS/9x
A0Aq3zyt0KrXtpjNXp+osmkQ33WCVxdEQZ6S4MLeelQ1j8EIEdf2MacV21a7KLsu
40GUzErZyaexZ31bhbKEMpg7GfaiHQwxss4UwsuVwJuxucL+jpqMRvJm/hoktBgQ
U0bSNfCCOv5WvGubOFKj3QSUupgzRtv9dnSVaSGzOCxrWr5Nn11FQOq7HEXOnHK6
oK/bUiqAYLKbbufNSuzSIV8FfgtX0bEY9dDmgmqbfDQQr8YoMc/LPxHT5qr3LqMe
AvjGMY+qDrsfd6xCl9DsgG4gYhIEPCzh9H9aiYRQY1cNDWkoqTYjwgiLz5p1sNRc
nt6ypzBb5lOcwaLeTKfgs2I9dYAX7YTfNwaVP97GXGVTTzQMy82x7x5cJI7N9NAn
uDPSsY8onMybTIdsgHX1OwwlT5TvCDhNNh2Q3zCU3xoQgxCfc9rW7Jv9ImsoRqLA
wSrKxQeYk6+E4LyJmGL6eCdbMo5qwRPGMDBrt5rdEgKbON9gaQs1c0iv9VydxpuZ
YT5uFo1zJ7HFAinFesJbxC0h0FPO5ADAlOo0VcaGK6qKImi+wuqCXFnAym6nZ47p
QUrmFocattSm2hmIcxp2ifDkCvj045OI5RchCsod6wtNaE+STSlXInnzYw9WUHFf
d78vzwIsVyPsgNPYNiGHiWOzFqQe/Z8KwCXGjRszCzWQZJQ5aj5h/TPd1i0KzZI6
nUFzjNBm1MmGo7JsrWxr/nz4jdZ8+VtgNLk//RP+lwHDDcSvyeARDMSOm78LzkJV
Y5R5Mo1ZUOJpJot8aQcXX7T4BmYK6rz2Hp5a51s15axE7vhcopoK2OdGsJ5i7HBd
8uAwN+iqVpMYtwqLxkcayoowIu/mWpYkYHY6Osepuq+uxoZpFhaDtNDGKXC4Rtf/
IPMpD1LvNM2FYbIv2gzZ9qEDsbUX/uKG0vcvHxigXIah3oXxVJx7st3cyXliWMII
TQQfrZ5wzxoG0tlOqtdiJAQbURbboEr3wxuRLFigMEeD0Rr/ha1TgclT014a7rZo
jxJKnlqP+Ze0QHma5YasUSpWRNo6qn0yXVKQrH+oKdBf0Uy2eFpFY/F0SY5SJ54O
3f29XzAP5s6CBIKRHsJ1Zos8b/0kZYzFsxYAoFCvISVz5GQ6m+ultAkP8L0iVK+L
NSs3vbowuk/59pVbl6Ci+Rl/uQi2E4ogxlOPkDQ4lPuPrRlNtOO+EsWc+H217wAi
65EUYnOlRsvbQ61HwZEhqmsXW3Z7zGX61TuU9twZi2P/IC34hbcrMXnewX1Nv39X
7+xEkUT491hZ481Do/X22vdvhPH1Uhq5ijTKE0YmnclQx17LBbgq6Nq99bWnahPc
mRp64nY4vaX32jINMwXfopJWp5lDFCQcfiI+FBNQzl4Si+xGzXPqa2AKGnytrxBt
5tVBZ1NEy/Rzhg+we5ndjnu0dy3lZ26eZ8F69ZG4AQb5dQ1VgTGF2gLYc58lg80n
pcWi4M6IIOxbVEI2Dvcjw9ND+fNrlu8BS58tse2QAgmKzTRrPVTvbAVCAE4tlO/a
rwxjF7RCcKk0JrAJRsTMtLPA7vFvwo0O1TlRGdRIum+R5I4P814ReXlFPpdw/FAb
hteTuprMlzOI03H/KkVrATNzugwcabIGh4l9LYpLurg9OTo2Y6Vze1ekuPyAlh3U
ygZH+PlTByBYa59+mzewz+PH3ZP6HTS0H63Oog+5w15ohiqM2NpX+roGxTeVf3dk
/N2aAtVZjhib09IkAryoPx1i5ab2g6I4BM9e6m37+B/dqGPNp6heslDaGkXOsREK
UQkwY1w1s+6r204Ld1bYbwrwpL+VBwv69em2sfGVoeFAjPQuPTwlQJnTKUSakURg
kGhgMdiPv9s7LH/9l2G2XGyNmcf83Af6D/jC/w4kHKGpu56O4R1bG6oqDX5S67Gj
LF+1lXWruBCOOcEcf6RqMsPOsU+pP/WtvltiAMThCSV34xK8RoR+2f3ZY+eknzGK
g7wKsEZ4xIkz/IsvaPWz2eQbppIDorCimS0j6urvbaTxoahVWW0lzCEfyhXQKxHx
0xWx/gfx1Jjh3E6ixwMV963t+4gkcINn2Bhu5LLZJlVpRptJIY/4WlAwh0Qkbb09
YwWr00T/ISRx8t8Ne/wGZ92ttnjerVSsIxNekuO67ZeB8mEyaj63LqoQy/CIRDsg
Ob48DYNK7Q5uzrNyrVuRhnyKlFUGNv+mSObVI/rEaD7RUkR5FKvy/WH0xbcI/GPa
8Mz3DFJR27sP1DuVM3HMFOIrJjSvfPSONZ1eHjYjK2STlzRxNXQtUSXbBdyuCVD1
Y2833uqcYtIBL3qXt7d6GpBzpgcDp+8A7qXkA66Dw53rijIDXOVRk86d7IqdCly4
ytkLuRNNf0m9oP2onIW6ZYglZuCHzZEmyBGpK17xkXlrPTD2SXB0VRIQcl1UKgE5
7+WmL3g1RBpdRJhkGQFSJCOK4dz+cSY8Vk73Y+6KqxhIXNZI4hDl0SltXxI7r3D+
AmYmr1DV3Ff7dWf/zslJbMICeFtKkhWpAia3bzOZ3xyfx4vb+EQpt8tSgmNQbw6x
SikFDoymA3c8n5XB4frpCPQsB8up76jJRlb4g+kifUyiyMsf27by+BVB32KMqwsX
sTyPttPWtG2YapFl5zMAFm7SbiXc/chTAufbtFrbQqhRd23LL62cn/KanrjHA/6t
JSjSOX/Ti81GLa7mEk+gwiwKHyTwpL9gUjHVHmLnoKWLM8vm+hrmSO0NST9BNmyF
8UelT7QUjqqBm8Nms8qfj+1Phqebsj+ySHlFnaGbK4F9xttZdY/XzVhLhM+qkE7B
qKBh/sbbKnQlkAmE6xlTyFqb6JKw/16KTMdIJKIsE6kzXY5ioz3T836a5UwE7gbe
/5oYH5HNcy2tWi0OVma8VlkRZGLEIsZMbh4ZnOA6BdDuoSK4WyLQvRyh+aIpLIsU
hUrKKC1sxqt2CoEAd2saPDSj+c/tSxGEGoESBJWSbPThu3ptDWNenhnGkH1G1bV3
gMosHSdKd5EDIzg8SYQfYAYNgUlpRe3HuaA0zyDrPFF3UVjQh8EUgJPkXatzE9gW
fZhlDPXWv6SPVkEIX8XSw1rP6t70VeF2X3Byj/J+Go6n/pNdzOaEHqhiHy9yJC22
F0r6itr4//ZOhIXVWxBN4+gHzL42ZrBXaIoO9pUEYeAtuOTWvlfW7ZXGSokyz5O8
HUEbwIsfuuYvqz75n0JmAAOl/meJL1sotyATFgHy2WL1pEZfeXHfDga0t2406gY0
RDbkZ3MU5EFx3u/unKbWleN4UszeWX3XOfl+nratK87hqcqvLBkR31GwyktJOSSU
vnrbhr/MPKO2mipHhVLWuDXCZGsK/XiCML81B+nTndeXzn9uy9TJJPdc0p6TFW2I
RFsqA0xmWUobCn37okPIf9DJ1dPgFLt5wi3HF1WwhMcWu2y9LBEtIAg4HFB5tqsz
9dNdGNggGfaDAck8BxncbwGNYjC4qmUOUYRzX8V7Xg7Ojf9QPvmKPMir6Aws4vOq
ER4r/yA9e0L++N+mmtzIehI6StCYPQPs/8uO+MKFo+PWp9KGnULVbvim7de/+0l6
fVtrYzPYoYxUa3eBdgK0h/1G2TopkEZx+Ik9hd2Sh9Y+KO9G1NroEE1L2fyu5iQs
80VndGzVO9SeeOpYLZN1c1qAx/TENvNEzd456hD0WZ/MLRCmB3C/N2Hh3G93AHAI
tVVjkHZvWYuLmbqi0rs0pOeDvAroo/816K99IHPIGNcU1a9Q7FbAOrtjL8Mx0NAm
ZV/0rHwuuHlZpTFQqnoBt9T4y5JXwZOa+LL3ReTmeOAlsPgc25i+cMPONQdoORPa
vZ/OoEZ2Z5aIWuvizvNuGBAOmG/UbnIcaIAcIxTv54EEnhvRVTvqW914ipPtsL3m
+F4/mD4B+YOBhYjTt/caaheTAajVuzgN2VmmGp4TGfHUJhuk70NhwJ+F+u0sDRyg
JuiyqPwIFIWA703KHJdAvtYYWmtCJ+XGf6WTmc/CDcFlHj7x68RMaW3X7Sw5pUZF
YAAkQn1mR9f8K15c2LaGnx10DQgzLTZkQeUymK+r3aaycAVOaYjPWKiSDXlHz5kL
+Gexb1QUqlq6xSeTij16L8sSpdRQMMfg2lOpehgS5R1x8sSz6SmOMlwEyfMzwj7a
J0v/ZQgRyWgsR9bgQWEmijJ48VwHFZHf15392JjvY6VEKmOVDzTCXgTYP5cKHCkW
+L3SEA2HXdIhgq6w2YfOxr5YytmgVw2olzv5cE7uqDURtqFEDmQxueBHzxXVpe1R
nN1Yd5skopp3n/x0b2fvFOuaPXpRivXRJpFt6OlGuiMfVG28N58ktQtXXdRK02xT
pRCEkrBf5Kk3/oYa9Cjx2l/J9+bcQlzl6VJG4qmPX7ViZDpBCwKVU1owGzxFm6zO
UCIDTJdLoBH4rRBt8X3nd+pNWYajLNmpz8gxsDadiI9Zf9zu76wHBPOqDL2WvUBT
2vbOCPlcUM+sXcXA3sXasQP5kCnLw4td0anxA4mWDXwXLA6ntKfD+aHu7jUdo9B0
zrQ0LvkNMIefRT6KYnFxz4SyhvUtdIVfsLrW152V0WyJlOuK4ZVmaHhp/z9omu7Q
OGzZFFWT8QtuO4ms2idvJA+5cKANBiH7Aev7YlPYdrEHOdqUhYkXiGGsK3QS+xZf
6/L9UuAJ67WuX1xSUqGAk10lximqD+jdzY/ahWRgAH58bqRiZ3Fx76/Rar9EZAzg
2HIdmyO+3iMbY0syJVmbpOs1IejGBbR+i2BGi7hlwz+NrhkurPuRyDUKYKj7pRm8
AE4dSezquigN/1Je7Z2K50lD7rz2nuISNhgcWn+EoKsgY4FFNrHw9p6D6drxhyAG
t47qcDDa4Ks7mxOZsIOl27w9WC8hT7xPT2ZvNizLzCSMR9c/mCKz4MzO10Z/KmM0
oWjFA1pGgm8eN+WzxBqXs+KqyaDWOEH803Py9IeqqEGzb5S0Yn/O45myrTiTBtpU
9NyNGUBSJv4/EtTSb4zbZR6VINle5cvbh/2SeLcTlVwBSfOQe+rbjSpMlzpUlSzx
s4v4mLizXcQLpDoHgVkN4zjn4WxbICtdCr3EeNrk6+O2Nyf4+oIF9oaIfa3CRGDv
KrbAJfVH7HgMXiK4bnEO7MwxAWFDwnx8p04jE7sLTodJfsvg87O2fhIQofIdWa9B
DsZz4NlVnzJu88gxNj3A+u8HoPNMDc2hgRvEIjRbMomv6GLMU1HpbWuZAIjFWG7x
ZE20bGKnzKXsPuPsk6/JpPFftVQEc8XdRpfOJ/hONWGGzdq9LiqHrcMcW6uiaCkh
tGyYGGvBo9AAaH1fYy/yW8T9OW2jXynM6l6vpY02BybaBcNvrlsKOVfie1jatXtS
Roy4Ue8dM76+fj1N8URcMUdP8rWh6JITHVkG078qGPwOa0Regp20o938YQRp7Xim
hm1mILWKt14yGzBODuEnFWpagg+A817JB3vaVQtXIrXG+3vxTo4Xga3Ci8usaM5f
pIq638QehlMVrzvYRetjMJLJubWDbNlXMC7VTd2VWYTG9wxuayEQmSREScmNMRdw
MHw0AXaZrZZy+YcdAtbyg6t2D4w9i6+KqkC1V0ajlgBrGLuzMhUanqLmqEO2swsl
mT8gvZ2s3l6RypymP2mU/v84eoJx1lESAirmtA7Zhfks0FePBIP4u9hcQbme9v5w
F1uV3rX7cmdevRSQ4CUm/hsrzxGcm70qAQlGAM3J4DMTm7I5zIKFngwIZdDwThAb
hsP1ZDoJa4MiSVrwZEdtoT5GDP83mcv7lFLfn4TciCbkoQPtm/76j4e9/d1siA4P
xc6jEQ7zNTVRX62YUf1TzJQidOp+7XH8AQKw8sNBdKp/J1aukjRzF04o2WVYFdsj
GszHlMgCnLLGlpCbzjB2M43gNu/l2MXWQ6jU2xw46pMLCZ2TrTFKoWkqMiJYRa+j
TNTNN7p9l4pP9yOG3CW6qh6ka72qeaccrH6B2/00jyBg6E1vHaUCyHzlwy80qFJg
H1gtaUlJGgCDBMjLVsU5i5QOUJQXd6bcAkStEBMq3KA9aocI+vEAvBU9oRURby89
UoWil/svVB7YYB8GHExEhcDUfO16oCLdTCQe4+Qg0EAkLG/iNOpPeCvLBqW7+ZiR
4jihjzHYB6NMnwq43bwhQKo/S8oO6AmA8S//qhXOAnTdkvuXGGqG+Ev2eA7L3PEh
VPw01a4Y+M+Bv3IB0JOSlgghmdXbXmLGcCiHhbks+A+dVddhsCWTIILVEnXYbt2/
UGRm4ai1ghUvvDCl7ikKHKKwCnW/ZX3VpIMIUvILhHXCk1VGoT4jpdmmhsZAxbmD
K/JZG2fM6JcrWILKe3R9D96SDdBFHFH1ApUOaNrf49z/ovg/rCGsdj/lrFFSlYmU
Ajlh4ThzRQC0Wj+S3gtHUmO31Nqk9WdMWBpw27dTAC4dk0zqDl13Hg1k+L6QJVeC
foEAgdO7fXZJJRCbseJ9xMDULScQsadErMsjy0dH9A851+4jqXgZW+CmCQ6H0RSh
tdCqIWBAqLT5u9XH5uwoaNpMq9nUy1rVww2n42jB6PbdypsXGgOJIvvBa4xLr9Si
A+MKtK9m7npO5/YLJH3OOMdCYBgK2RrJulULokWm/1azPoLMAf29HcBUhhnOBckM
5urYRwsJvTAUOP5JydR2V1Ir2DnI1ofmSdc1YoNIoagmh8Hd7MpOAX++DfwL8Es3
p5MxzprWapjJo9karhffhzISvB5Kabsus78jSjFmw7GnL5+JYWAZ+o+pBc9OPj7D
gdWEJUwOQLXIKMmZMQRSIkUBibCBHJjHLukZDLu49uoPhcPEyXo8ZFq0Q0tYONaO
yocIYyYYM08QvvAH25yPaahkioiFeRHpBznS5Al55pnjdFxjATEhnhN1cKpwmDJo
H5iRIXaCt/Ksi+kQhpWqDCS8Z+DhSddhbOz27a63jvLC72lhZlSXeqcTyp/enAhF
qsS2M/tDYYofRjFypxP2h9YBtuRKkaLHQW82aj5CobnGdg7q5CL5OXa5/Y0G3XO1
yL8rZKKvxp6uiZqiFgfsbUvPxByp/Y6NZ7DvOarZu0FYw//P4Qre/8VU1kaFPBMW
kFjJ7GZJS50GlW6DGJ72VidzDEI+aNfYyuG2pNLgIIMFWVb8DKdXOXPIZsiVsKSG
lNXA8NOIxG0yd0eRr2DfYfQMbzoGu08rVBQSvnH2bjDsGwef5eDaTJJ6SXYMMaXk
H2+6n+4pNfCEl/yQl9M/njqIdkk/sQaWg/YGVX2u7haV6pY4uIBMy1Nmcg8pI1c5
Fka1wujuYWK/beO9DIiLA4ZbctUQ0b44/VpVQ3eUseBiKBCs3XG07GMfUI/dVv2o
VC6VZaE+DlSHwzK5UsDHNymqP2zjkbVzusv4Adzj+HZAjKdWVCOc0o952GMOIl8m
OA6tsnPS2XuVvgWeo1xhto2VT+OCGHem7B9v7F89ffnq6cEYLlIcP5kZfXO2pUZl
qIt7rTO5/nXfp9Pbc9SS6qMmSdgAUsxy6I5VY/cQvhebjGV0BBAJyZz4R6ik4Ks9
SkqkyA2XOruQqWBVORGy5zqxPMldZ2zAxzgMhjYw5e3+CL3o5KlQMxweJGVvLy8Q
Mewe+sFH7OpllMjq30acp5Cy2mP3Uk5yPyQOVAMNs0ClaId4ilYjhnopaGoPZodC
uJ5TvC3vNBZnsYQGkfPiVuylthfZyRJzLTIlGHO8ibgukM19HGFxzOkrCcl+ZSvA
LqreU38R2hWV6lBdJOP8FHD1SrdB+b251qRXwdzIBLaN1wzEF6LdYtRW2cf0gL3W
gZBtOD+4NNtyzSvCW9Vs2vcd064Py7vtgTo3yT7IeGcnOjVFjRQXQBfoLcoOBXQw
z9ZO3BTqDShCNBwLr68Cicrrc8Oq+HKbtqMtNtiRXFEF37axc1t07Oq1WtwU8mBg
UDvA39ZcBhQdncuue9JcFzdOXuxI5edPnNQLUjbRWLuCLHudUUQJuiixifPDlPjb
YfUbBpyDBV89NUDJPi83JU9l1pebWZhSLEtMS2D9cfAbYSVoRBrrulDxG1aL5FIM
fPZdSlVPjaTdrDft5yLgnhumC+MiKEgnAxefZEGDHEpHj/oPY1qYPdGissXFEoiJ
JprIoUXdSOljXSIrhp9N/hCcTPMt11wi7h9xJz0ZCwl3q/BCc3YN36umFrCM4iL/
p0n1GRQFnwOT9oVokxaVifp+I485CQ4Bg7s0KUjSiw+DiEziu0C+gtq0YeJD76yh
+TrVN+9jtI66T+vvZQZs38q49o/0Qop0juvDaQluMAvwEPEcwXBSREqa+savjRnc
cY7WgC6PwuDrsWeDIhHmWHFNVj+sUf2DHstgehJfyfO9sFqRL6k74QsIdLETNRa0
PuKs1AOtxrvM+yFqaz4OrNkPlrXkecmyKdp2jT/iQ/5Zd+kKjwzIxe1qxzIDRKJx
BEiHeVsf0WAZvi7t+B+y59c3QHE8vhk8Zyva8BqALbnrNJlUeLEMEAFTjaxqBBYd
tQYOijI+U0qkRct3nqwl6BGc0wa+8DBloa/5+ufdvADSH4YeElK/RrSXLA12DyUL
ucwflSuUgQT6kYuqQ1gjp/lnXOfpAuhqH2xwxkDOyNF1r00vxFr6qI1LFQwkhELa
LYtEr70XYAsd3GZELbUzqqDEOuhPqHjtL2H71b5rZisLxljVc75XgkyTAc87c1/+
KyDB82MhUxkYJ+YOj7dXow0UiMTmpG9TRvqJ8sp2dXP6wZKttEUJ6JVmCvgs1mi8
3MaPhjxbcSZdp9hWXZvjszkyvZLWPPMy/HYu5V3ckJL4bQBOcuLXhNoP+3016Puu
YOirY6GsMekKQuv9saLsMDwG1D5iQBnIsLPZ/6pjwrrfyfAAPr5KtbdcmV8oe2x3
6Axb2uv7NRtKRPCqP51kWPJnxeyR7QG+tcVglWYEXRM2JDugfM8a1TYuxLCx30iG
vqOnPHwl/cJSrMFaG8trIc7FK4gdZMKA04II0AqFbaeUxCeGTV0r7C88KBXrqPVV
N63eLKv37wRUfJXKHUgL7r+TpoFLbXGmiixuShdf5JyWH2mG1wQvlzBG4zAaIxB1
2tCzjwqyzrffHHKAPl/L1/uMFaOpAg6L0w43kmA/P92ApWTfHD7Hjn+rZ7X+hUAu
H/FqTbbC3wdfukCnihQjiYnzBNwIhKwyrM7HryADoI8DiZj+sHyNBNkvdGdz4m++
PZJOLa3fg0ietXiQyzZ2TaLubFzAcaSf+iCspx3iWJeDIcxu4iptSKCkj6+r+Bsb
cwLHLWqSoF6doHWB8scNoCrVfAirZ4vhvng+iUjSm5mQCjQWEhMz0GV4Cor0Agu5
RLQZ71XN2Lk9Y2J6F9vEIQMoINqCVdEBWlZjwlu/gJRdF7WfohULHns8vEcW6bo+
SBH3BTArPR3HkQhHalmK+Xcd8iweQc4zOz1cAWvtyptR0gPm/TxbE28BEH7XqKAy
zT1pAyKedVjcrI/wqG+GMWuSkLfAanrNmWAbar/VcqxuGxnp4IajYagBfBxsKEGY
i1GKF2SWjqiKx0D4RwyjW6rJph0mEgWbnmiGdQwGoYJvh8uR3Uq1KtQ0ncy1Gxgb
kDt8GoHExuINs0+mXnTVEvPG4rh1dZxDAs2ntFWCBH+pidydovZt2VXOzDwmTkvG
LB+MiAQYwnS4FYxVVlOzcSB5bsgDJYJoTQ2Ioj0kxe54yJ6G97Y9uL4YJv2lFlrh
Ekl3Q3JMXHdZaNPI3/942ek/92TXnWWvOCMx4jMYv8z4bLnJAN9I53e5aKgzqHRH
CKNPuMlFBNeQP2NmETgw/Jnoou16EMC70kfayR8MX+VWVoBGwk+eyD/gF98UOidP
BDCS0FKvIYRZHda3NZnCXw9ym6Jgmy+LF5Tw6rTJUrq4NIO/A7sk3c5ayzgjmK3c
k/H8Cz+pfwJt7kCq8HhVFN9w2vvGwzXCnZSwZEFFbC0UxM+RDDhFCKVs8N656ibO
9ca0RWfnw5cJRr7TyMQ6we8twGuxSqnJrfw3IMVtBVkvF/2royRtAZDCjyzUXsD8
ia7AFrsXTGWFyn5f59WS5A/DQ8LucH8epBc61rl1uR7rQ00cNngWnwdbJ2SXdywR
vY1CITxPbzoSmBPb065bZIwnM3SKXmmWlU7oBvjXD0vw2yEzrxCWgfCyB4cAxLgB
alWYnie3O2Wtb/UX8XTUnSbwUe9/wZk8U6k+K2eT4Wp9Gn5e+m5QTAtdEfLa42LP
Kd5fe6Eksgd0VYCHKynt7vEIDAXCqZEiU714h8rLKmxhNqOP4qJRtiVK/DQ/E3JH
3NSHNwWLIkDVlErvKzn8+KWnZWgrEaHR2LDuyn25foM4uCch+0IJQckKGkflYv/R
UnVLDJ6atQZLs+mVZv6MPfH1Q8+Bse4bgJIK3lmyax3PFbCsb49GVTx2mF/4Sf+M
zGQTcgULg5AIZkymmnuzvBpwGcSCBumsBxoyP3cv+23SVtV/MvAk/rgCrrFcdV3n
7F8lvYD34tgJ9OzleSs098W7UK3DW8CBPA84PAeMdbeXOz8KzAT/hNLv7WSo+tHz
l90wsaem0kEGgxDRfbti/Ylpsgy5nCdR70niXV3K/gSDWoyzBFPYiM3spi7wMvjd
dSqXGIH7mMmFijWSAg3mWmVFe/BMraq15ggHoWvnrv2EciBI+cukboR27LYSmA2O
fFtlvAimQY8swZpIdm+gESlQrBS8zHcL85VA7B7SuUlyn4igfTNbS689nSFQRC63
2hAVDumbkNXnJ8VzJsApHscaA/DtLVYyMYnfcWfE0pO0Qs/wb5QV0+wjkha8qoUW
WW2/4Dqh1kKaf8X0NZmsOLcH2cdn4iRir0IYPswFoR0DhXiAfzuM8qoT6TRWLNu5
XRpIh6oTmmAKnZ3KtSDMH7AGzIm7Sv1KapEDGRmhcdwyElDGpA6IjPav8J3NgaQy
5yRsxNti6/HWoryQQB6q6UTSnt4S7fXENxrmJZ0V+UCzPtwNn8RxyvIgTXuyYVQA
Tpgtz4IMw0VG/VzAFGMB5Hzv46esWayQ2FZG3rnDM+f84bA7LS2NcYjyaTXmVaMk
CufAlzvM1Ad0MaUhB7rAJ5sV2gkdF0MtEmC2kORp2NLXSQTeLOn1hiVf7BXzsKSF
EdOz2ojUVmsZeJvK+CH8Rxqg99sFO48BDye+BkCw6Nxy/GL1F7E8v4uueFUoMJN+
GUwsqBw/Esp60U4MUhO35W15Ij9rEDTSPeHhpUQSfKoma7gi4KM39hUNMHrQ5J5x
PPz7sd1INma4lT68/FLjhO1XfiQOaK2VPMZHky7kdC/6tInWltOwZgpkd+tI3Ep2
A6p3ZtjdL4TU3ZN4rfmo8OPpJjnY2hqUfWrsJHYU1CZkq26mChVTwifZSS5XzjGf
Gf9o+VjdRb30qv5rbXF1gY6J7ENt0SfNXFHwF/QijZRUhS7mmkRnNEOdtcsQPOWl
EBlYK3oc9DMHszUCftyBnYVJY3pvQmJqdhP9/mmBwR54hio2xr2cqg9apDxkMlGp
qjeB0sIBy2txBiD9dbiysFO/ZF9ucfWVL8/HUc0Jf7qq3yvgc6SdTIaVfLnjFV68
AjFkl1f7UDhU/HaZtgpVMoHZ4QZRqlV6kPkpCZIWLTTFaddgSQRQeP0viSi9fnM9
ymkkDl4UvDEM9QbpCIROMB69aiphPK1/W0+MWEPTc7MTHPRa9O4WIovZ4y+lGcuz
PBRUmkmvZsk2/fiuuvwH3lvnw9GD1rYP1UEL2bmEKYVtlYNrSQ85LlMZRqXG6jdy
t75/USZH0jQgu9R494vG4UzRZIk/tDDOJ/GlMcuOTBTcGSXS4HPBumleoCr1tODF
xNPdgcR6Pz+ZYKhQRw3VcCA0GSmf+tqNwOvgRb/SzlHEgk6bX1LExPZ6YEEaZidH
WJQAkkEDEMiYTQrVhGpddra9mCO9z6i6C81IS5qtTa1/IviJ4YZg08SehZYBQb7U
ri4SqmRcoEn6V8Hq205aBHDFIp1cw4dno7wTpKWpftkhtjeUORo9kI29cbAFNWal
paqsIH9rAsl6l9LwyuwADW4ddr3B+uBTXgv1BqvkWIlbXuPAmG+1wIkUPlX5KCDw
7IlRk1uqk7yz50zTRQy0n1u+R//dU5+6RfQZNmYek/S++36jPI78V0/tdpUxMyhd
FRXC4CSPGz2RhMA2dEG0IDhK6Z1Pt0jl16rgCcBjshlJWHMIJ0bDZvo3vPaCa2MJ
DBMT0OIXWSdWpJllnZ7A+P2O1VxYoDysZM7iraI3JLd6KsxbHDWFVUqAfmA1nmvT
kRpIDs7A8CUmVNNm5KifTPr7eH4E4rdnfED6bgCc26Uxt7egBzK9ddCVvaMJe9nN
BHxSmOEIXTrNcQHpztE5CRcmcazK04NGoNf3FOsZ6oTYaoOy74oWiFEhSB9c6Wa5
AngLh8ttAzzmXwcCo5BnQbYmsytWM5737oQ6146ZqyDp1U51YH0kGJXX4XZ7KZ+g
2XZDfX5YWZRJ+HOJSjQop+xL7Kpfaitsxu0xVV2moAEpoyBz/ZcLEUkjhJFiI+g5
ieR0PmCYLYChatE9Xn/4+3B38f4mjT8lsjyVOChc5+QaJwdywcWCgZC+79nfNemC
lrxj5bRlYfPODvXaWSGygzfswkWr1fP/8EcrczAhVreggSv9JF/cOarWUM2lAc1n
0YihYOxDTVFQsmPYqKJOTXKApgqzwhTdWeujpmHuZ6p4uJw0ZeWpwQFxNSdUwB6H
gabzQQZ8vVUiTfRWfrWc33akCRMl7bsrtefKBGZyl5t5ML0H2onr7dgqLedxul53
ZM5OyTbhflHrrSQrhzg+S7Yd5Dc2S/3yV+f1sHEDBGiZzsjHnRbxkWZdq9z7QNvF
1qqe1XrZRqGjBLfVt6MZ8M9P9iCoqhj14aWvZPli8aqhquK7yw/sB0gGQSJ3UPlu
13Hi8uL975VB5uFKlXwvP7aJ2h5ycoCUSo3N6c1l6loShbMFwZ/y5Tnu41kJdafY
WnWsE1tbebIV13uQrzkfMQKe3vkAbddRB+FRJna7kh+n6zbhAZop0WFXAhg0UMrJ
oAoflDWR9uQqaKLLEbDuV58dfMXAsLpkOaLiZ7WAhE9dCiJrOtRiRpKkROFYxDhr
LWdquDwaK6obVaCtbRxnaNCKPlM0+d1Rl9e8nNYQ+yzqogOUWciHte/guCKK2tLa
TQ2JAWxpisZLkW14eTKEzktmL4Ci8gYrpsSRk/6VSYTDu3JYAwcSNcCLJvuWjq9/
ZGzOA+wAfnKhTCVxJsMKko1ZteN1Rskrl8pJNmt15J/l+L+JyKgXMkfU7E9yjkx6
PrXB+dNecOcUxuBmdZw4Rv9qr4LH1d9IqZtZqSQb/ThD7Ah9SdlSlR3HiJVIcdz2
5ZKVlInr1vcThcEf0SzoKtIBXQlfX8MmnRrot5EdMq1Uza8oAKm9MqXic87XVxep
BQYH6yPExQQelYwRsJWZVfpKLKI+prrEfirmbSeiUxv8+M02oYhkznHNy6JBJKWe
CsAYxmdlvekoTekUf6872T+dhAAy+OMbj42lftWGC22MyUZNHQc59WI6NxJ2+XwX
ctsHOp4tea20MVBTqlbojAbj8x8YUl4aPrN98WAgyCUwR8TNVRhrFUmTOXwRRkoi
7qinom/IUoEAbLh0DGtB9C/4zrISMbSHsJQ2nbpEczpsaJ1wz7HpnliriFIIHKqN
9n8wAAZSQRlNvUZn28QruDVqUGGi6TQW5Mht6K/nDGazSJrXIeo6owYob0c60etk
AGZ8Ie2X62x+3V7VqGwJfqyboZczQ8vKFoUQ/MLqMfVbt9xHm9osYvEhCoem0WYP
x+LKaKNV5uxlRGxj+XAKPKKSz9iX8pV3eiVbKjkLkMK5cf1qbaMQJOEkzGhIBUkV
haBVrboYz9Ecr3nFofEo3mDjNipc4K82XmfrEdfUPHDPR9E+N2beb9Bb+a1Dk6BS
kTDcdwrFKdtx/PtNooEz7L9u25Fb1E+/Vni2uk30Swd+DQjYMn21NU9bzHxIecq9
2uIVNd3Oh+MiSZTventLA0pNBxHK6uXG60jP3zq09fImhbFmrUAmPCSt6vwJuWEs
Xj77Stwwkv0Sd424eolRUbVo5ZmWVXeCtD2Z2uqanEBdfX/ro5EXRFEWm7odb/p8
qDV9/huxwNFKd82X7wILBVldv+PmzQzP2/BSR81EKWprxNvusOwO2KzEVR7H6c/T
g+vnJ4bb+Q3nO7/41Iar63FTaGyTBqCwjkGEkBKgW632ru4H/Swr9PsAAeO1jP0F
6zFGbrjgG5gDS687p9TyUw5wYn0rlpQcqLNsKNAzeq+3qnf+0cEiAnIc/GFPBxYa
TQfJDx1G40QkzsyosRIJYeus9j1/ZuuvSGWI3y6bn6Uy6Qjl1uexH3KD5TCM2weO
M3LKCo5K75MVzyPXYHNbCRU8RUvuSStADF73XgAYdApRUF/qnfuV+/9kDWdLFcHw
1dLUfSU0SWUm+NaG+t+3kwHTut4Ems91vpi3KJyrVZg18WZmkoxoAGOoTQecWhXL
mvIx69i9VRX6oJDR1aQBHE+DLqrZn7P2tBYm6ESWnTSbKZGz6eTjS23a19Nt0fbd
ywW8atWNXA5KOLZot/ZlJwSqv9IPlJ+XmXAdJgfagcAvEgZ4lC2nSHmGjftfNsev
cf1ZULaaDo2hND7J5eu1ZFDt2tJH1fOdPQASBN+Eo8kqO1RHYnwe8W9ZRQ3/iKm5
XWgnGS3jA/mVQYHG3vRjDrXU+PWgjuf5B7B8qJ0dPpTrpJPFaf0sB5s/Dnsy5z5Y
+riGjxs1xCekDo6zNMPpVAyEL9njaSc7A43h/DSCn/skY2AeoDvCKEry8s9hnOE3
U3zmzl8BkHehF2KbEYVbaa8bOAm/fdqMNXt7j5UBEPtqaIcHfVra2OSlijxE8V1Q
4A1/ByKHvqXlpSOYcnb9aGZncshNUpabWvFpktCx4fz5wqVr0iEsNt6O2kRnKE8D
YoRHeVPkYgJHZiOV9Itigd4/GlWDPtH4NA/JcKrgDbsKbGi54bbsYant/imvd18r
lYPIyPuKT9QfhlcVFfSJb34M4Vkojy15Y22PlXDZhB7wl4JzjRBQwV1xkcUatQ89
FULt0mJw0DRG/lVaP2XMkNWQyWD5EBeDBL//Sgk25u02WqXCdRw7TaVcQKqtLbLJ
mRyxfvFaE5+kwvUZ5VcNtWZYEls2HREUbmX1EULUW/0NBdLrd1VXBf13RgOtmAZK
/ZylWV3zXdnsxfUM/jvQ6HJmzEg35XJLzCiymTO8hbGnIXYRHASlFMiTOx1Kx1dy
1jFn5RMKoYhupXdArsxL3WiM1hDtABCkCTs/FZ9b6CNP54MyKeu6O4RYA7RHv6xV
xQZ0WNJ+3QcBDPvs+ILXurnKTM3x+/SDHLaYNkfjHtk9sQ7TMshSSIXD5gkKdMbk
USS+e0hBWJxWaXjgHCrB3IbLCBIZkE2eUr7RMRBI6uyani8xMemJzZX3jG75vuTD
nxWnHac8ioF1oNVXrQYoTV2fLrYwa91HqWhq/ZJ/fjVJPd20eZzJdxKs7+wm7Z92
E2PswmOgb41FueiWZCyMQFdto1Nsexh38LhyEJ5Os2htSxg2gZ9yse8lPArmKpu0
44lfTJU4qdnnw+hORCKDZr537ZaLx41Os/HFPy7RNAQBjcMp02Hh+ohPXOXffv0Y
Y+iCshDARpfXs73MozSP0zIyM4161jYV0KRldQcd+f4ku0KxMYK6d4uZcAZjlGRX
6/bRA/JhtCN04sDYVfH7Cx5zw1rOBt7oGOrl3+LZit3n+7Ol6r8KFeyP69wTbP+j
hl5xeicfsTaldiLvidwZ+sEKST4F5MPVhgqdiYVHUGmrfKyiG2n5wRjdYFnNg7TA
kDxo6N0YpHobjQglKL0fCvAUrwZUk1exwZLAkBoWVMgqog7TUywiEMD8/8L1I1wR
7KQH6WpiyhSQ0o8uZlR4mIodmJ+NByVdug4DG9o2jdp5wdu7HJpkfWcKCCpf9fwl
Qrq1yOQeIINaXbCxEnkcTj+2mCioqb3z9WE9LMrRTCvq+xFcUDxGpkWh16KILXww
z7LQt4vHl2opnFweotC/vJ0jr3Hf4SUED0q5nlt8qACINLtxdsPiW1rfu8n0OEru
IMy6rVFtH71lh8gFhORcFQAFm7FFwczEjfki2Tvy0lDl2Zbufn9+8mkGHJeKcrfd
WwMZue0huWfvTf4K90rFtVshEwDhN9oHAnSwxcuxXvNUM9/DynhWkd+cvWjcwJsU
JDW/o+6clCQVyfU8F40FOcSyvYcSynFwy29GrHjwSO8shVyJb6ICUeTRo8kqMCL5
I//00G4vh6/8u8ltYX4CBPturebvOo7paEjRW9IshIkK/K43aoy7igUtRiBokAjx
e+ezqZz15fQ9O/XEfpnFf4wMKc/3JKxOeG1liF4SICJX8xm08K1Gd/j6vpmgjzmj
reepT3kc3EFP+/YBuNkoT4r2no8OuNyVtW/hpQTMWdAkixmUkF/XHqzFj23bHhhq
fBW3++KFqu0AOsBWYiBs8b3YQHQGpWr4EL9IcUP5nhzmBOJ352/j3CbNh8b1uNdg
4Mdrd03xcwWz6EpGk2jSUSFpKXSW1sHiqfI0YATEc2Z9U8C+jPM+cK0zlC9Ttyu1
HxDKXVXt0LDvJi2/QmQDbudqO0HlcnssWhO7/+JRs1U5cijQ194T6g4QfiDzP1mK
2Cm5axDSiJfwg4HhJ6CaF7XhUsjE7NlWlLKj8cF47o0BqzsV/WtidibfuNb9IHoq
LgwdA6Nh5dsJiFDOOHoPyKemhLbQjp0EwHwu1UX4s0qXpzRpsfU3FZSkCr2KhLnc
SoZ7rKXdKqJmaSEL87t/wvtjT2T8iH/nMcDEYBYjdLuIot9UUUYQ3ke7sl2vI+PY
FPd4x1FbX1Xd+Dz5eFEFYqZzok5WKolKfV3wWs4ubrMPDESoJdGjmIHlnAieetfM
kpGMPZJOTc+yvUSmZSQ3PI8PGlrpfLoazVOMWTXfojx5wwjVqCgGOMetx836AKvw
lzYq+DoIV2qgdzHgcourwXq6fgp0SU+bZ02aJw2qlQ8fHLYmSmEZ02bA7MJSsHFr
egSjEmcq0/3CmOy4FA1mK3ypIQc+4LDsP+4h40tlAHtimCaQlY0j2amVuXSQ59HU
FpjKJ778dbtOdCFgtRATr2+c3txo9+r0eV8wey7cZwO9M8RLZYihv3BH69px0dbE
ygEoGe4g13+qO/fWsaH74yg79D1/N5C6Q+CluY1X1BIlIvF62/xxAJ486Z3+77m5
9N3hqSW4Sy5rkZh6olDONbZChFQXb1nOO7kKkTfQrY7I6IepWNpU2NP24Wiv0XcT
Mpf0s/7Q+R9noin5HwkZIuMKZ5WrtzNeoxnbRUzIzyTLBBvs/Our0aPe7FXbRHzS
u/XLi+HUwADYA/h3hNyIpoI7rvctM3c2gi1EEgHBe0TzDNaflWGwgmf3m7naPSgJ
lbxpe6rJWoxcFFb5uAjhO4T/FQdk/QYp5aYzvuR38LQYTuEj4hbzK4YCPyZXjsSA
Uq4+WzUEmpzcJb8+c5esSqaTMeiAHunpcqvS7pk1QgXSvCJ9hvMG/Ngf7OqOKbym
lkj/MTJq2s0l2nRDoAilWrB3I8tH8DU/nf+E6QohvAdrlHx47bdhZuAAf90Cndon
siu+UcPVFCtGZxwLPt5Jy6Ow+sYfTSmTw1Fj9UZZovqdXZQ8SGk5XKJ/SdzNSqt3
mPPzX1Vd1cCefqDE2kmz2GtGoNmgynDp2ma1PC6RvOvl6EGD2O4tO1XkgmU9t91R
DtGAnWEIDzJUm+anDpNZlebls3RqG6sCfev8Pr8wvKwcCmZJxDafdpQ9tgQoMUXX
8DEF71pzlh5IloWk60TUtt3rXvBnBbh2jMob8YLqeeF1jqTxrney3Qriv875lQNZ
d8+ydAZ5c9sm1LiK1NyWsISw2IrY3fPdBFQNBKGw6HO5mv1HT85eFlPQiwMAKpH+
cWxj0RZsDaQyCqrshABZTs5Btwxn4fOS4XyI+9LQGpRkpN3Q1KbNHyD0KGJuBKHu
MHwvGbestdYkp9T5QI1JxQexXUd8J6OzyhMwVBfD/ItQ4ypz17MhF+MP9m70UeVk
zf/GSJZrFTJmKgCiO+NIixQuzXHNwq3J8Ia2k6TsD5LnH7srGe64EUYcOUT0C50N
AmfHsp8X/33FzOG0EZ3z7H8wCvhxtUCrwSVvU9ikKBIjYbdr5E7HoRJCrzDmEmUv
G2RWrbR35cUGjSX8+wkkhkeM5Cxmdhe+hrcF2LSyZBUTknTYXJpA6vIpKcStYYf2
WNgQBdV9f07Ezkvhhw+Rshb4ukVpYwe+iw5yG5segYQLLJ89GbH9PuMHSMZF375w
7V5vvTuEEzQ+SXvtJq2kG0wfHfW21qs9sP/OpmURmMCN0LQfhkZUCFrBLRLjreW9
g/yJXeDD76lJm+rk+W8CpS512tdN3n90jYu3TluUYOP3mJmliW4b+dEvn3wldJpI
th1NeRv2+nDannlnZ2048vayWnB3WDr/108Krs5mxNDEDsWoN0koZ9sS72dK/Xc2
JecEf+5efUY2pR5lukpesKSnF9LNl1mDsUPn449HyEqfxKYr4fRYuDrhqAOLusuo
qyThAWMbOKNhj+keu4aKjLJXbJqcuEtr/fgTCa2Bee7dVOHkEJkkzqto8o36Gooj
ottLjrrbopEXznZK7duDAG1oURijMjvJycp5U0sOVd2JTatOHvur9h/ZxXgDE3bc
LCqsrvIyUg5oS9m3TrySz1ohQKnkl2HvpmzgFIzOMu9mUiBLZuMopMnJKvRVXWLw
4hUMKpp00sKHJFzc+tHQhK3Mv0I5KENJzNRV4MIMwEVbt6PV5pTQgBlM7u2PIZjL
oZDsFEvmx3Y60zZazDDc4ifNOwH14XAw41Gt0My/Np42OoPDFkg8h1RKUMUiEE6J
p1BhpOC/MhTvDeRXuuaI0BcJ/3HPDexJUgpwYMJIL7pbiO/fS2H6+yzD2rmLyM5Q
lohO5DB+G5tXcJ0+inr0pJ15QfyKK0yLmuoWXLxvQn7GsE8KwCevZ1uxW6tZ2dWi
UesoQk6TTlUyYJoCn0mzaoFzWwKjjuUFAvmoeX6lUGTtd8acZNhfoxQBWfwMsSob
DtF1LrMByT2D6vhpV4hOMV7KDKKBzBuEpqnf7AvBFvZ0f5nnVSbY1xo1qv/huddC
5a7h1Z5fCXB74GHzoMTkdeOEo75Yq92QgyYBBZw8y0KiBBGcJavYytM1i3TUZzc2
RbTOLD6p8jWrUKA464GRGLMwg9Ec7xFMHyDgV2b1vU8N+mengmytnxpiU3fPfUjf
3PyIoogNxkuzBIv/PtIKvg1TfH7AhJzoqkkXyXYBH3r2IDicy35KZ8rWmXSiivVs
4W38hvoDxdKHsV9pEWBQodqoo+YHHykfJsPX4zZOMpjhPCnQTFy5lfAy+/XKZq9u
fXnvB4IMfSmhYb4VaLiMJG+2C9YSmljOBmr3bbIGZMV4/uPcESididjIOfxC7gfc
OyNkMvzXKdJS5TZxz562lJT6gCcLtV75F96L20ZZ7+/wgD+lBlcCEhvp8VfxaOTf
y9IyjPRlS9aKL2vyeUl898H7wqvSg9u4FOa2AyU4zGuh1FIsRZPqskFcosIseSIW
7S3Y4whEkstKo1s88a2zx/JeKdGscVe/ijlGVVhWc/2+C3ezAI/EdxcEt6R+PcHx
lQFaTiq1GEKkE4U/JEu3mLyRW/EHxOR0qWJqNdQiPARd/DTKdnYCA75G7TTzv6ld
7+D3rdnSaEfmS9WXGSQwzKtaBOp2TgpWG2gyY7BziU/6hiRMD6qMBiHu6c1pqIfM
3KgiQLK2kFuwwqVZrpKWrUSVB4MrmEj+PqsrD0iiB8Ux6dzIFt900WS2AQvWva05
xIqbGUYw16whhBKOTkAlQ7v5S0UCv6gpZ7y8r84l4R9zRzQ9v6EEwuypMr4BYPR1
blQrTiL9NLzTS1BIbeFQPEmbB5J8vBfYibeqhVyvxka3F7zySYJF1854jwOB6Yrb
sEpdrq5M2UNUy0pkhTnZ8AaLrNUjrmfmtgHokF5Yvsnt5o9y6JF/G4HEkHkK0n5o
C7NijFhMbo2bYv5LCgc71XUnbHQwxGI/P3sKpttiG378Am0MmyBzip/NsB66/gfM
afduSTiJDIgDszg1NE9leKGsZNAmPlrDYxd0C3qTTezGh2Tkn9d8CP9DJljH5tuS
ShQFe3KBzSePSd7GtQ2Bh/Jzh12K3hBQYGbvb5PypV6LNrIa0resT4f8AxR1OunN
OjDnc8qHksH8HoEpzlLT/XXuRtp4hbZkpzC+Hdw0AKbuceO+JOZL9WPSE7a1ajm8
tHyUjAeI3b2qYBnpGKk+3HoiRJ9jcatbNQtQi16/J74z6VEq3V27N8ICalx0VCAL
x8yYNeJv+lBUAYwkogXOwY8Eh1LXp8OQ3Jd5uFJp4W3c7SD/FPUhJjM9W+3Kx0KS
2yBrRf+rNv6UhdX5f4Gr6bh18K/XezO1tWtyrR0ZxUPnxtqWtJosAcXZmDYutOUD
1tHI5W0iyefDjTaPUvZWWfM8YwJUfVbILzBVr+1+FXlxwjp7QO05nhP/T1dMk7Cy
ti6ydK2mpYXHiCEg6e7+QhXDiLu9Eqs1XhZmWwv6aczXwWm/E0DmTpK3OwrR7idB
2VNG21OR8Q34jpv10tEScMG6nCbScaAQbxzCsHlHcUfFxii4hofAK/AiXUZmwv/M
FR/2TMgQXHJTB7YhsRkxjXWfYadfWoUSKbbvwmbpHKsUsA2LZ0FBIioRwtz2eJ3W
U2p3fDiQH6pWn7d1LPRoJdwprl+MjczTaW/RXM19qabRum8c1wCRQULEc1TOcFE+
5Fhw0CKySdJu0GVfLmTC2/dMsgtNA7wHFo1GI6/M2mzvinmh19Ha/C4+SKKA4m7q
wX+w7NgX8xcNwQYE61Lb+h8kDRQbrYBgE9d5rqBCafGctHHvde9RN+mtzLsMIPCc
n2TJxl8kDNxmL6ZBJ+qKNKB5uaiog8sK1MvFPmXg/8k5LCmJ4L3Uadht8IZvazeM
RP9lyoJ2eeoebSJY124a0z/q9Ke6+XA46WDWFMFuZgKtK8cs23kvBeQMwzeu5h3+
H4dAyWH+Cdlq38SejyM6ii2ZF02HN2Hjv6uzsyxgoK795z5qM5cOdrzJ78fgJbDG
cxXl1w3i3XHW+YFaihB2CP/nYdL6dll1lU5wLJWVXOgmpayfDrdcco9w0V7Rv4Lb
CQCcVQl5j9D+D4ChpLiV6+gNGJ6OK5LUVzMSSlEnhPSJW6jnubxK6JLEzeYqv6KT
9k7TBw+wj+pWDUD7h3I5XqFf0Lh4O0w6eTrK3uI2lXRpvG1qzQ9skj10jsqc/98d
Fze1ZAZbGjZJaAMEumj0Te1dyNGYGoIIeg5dIf9Kunai2JGa3HJLjsaO2dNJJk2n
aA7l8XhEcVh4+7WB8UY1rtD1Ly7eGkoAaOaP5Z1uxrhAB8xWYd/gmF6TORjtN252
Pfge3H7Q7EfGRZ7ed+bSfSj64EIycdENLUce4tvDr8CTBbeAHSrXhZKWC89f9mum
xBCfZ+QVEeYbdqoCWBchYc2coIOGMz61iS5gUI4FvSQi+DR1PkP8wXM/Jceh1crD
iPyBNq+O1qaMJwEgMBcZTVpgNiQUUpv3sVBQxXjblJxauhfsSdYQ+GKBbVmPPmed
0axtY2RZ6O4C8pH+Ia/JUoaUo6XSVY+MBKy7cszICevepDRDBGadu8jGHgvGmXKk
1TppdbVsw8ZjP62vcgtrz2DkeptJUrF9JkII5eYBorLodjmu76d3D0s8HfuKfhwS
OmFlPh6o4fgy/v9dwNhsM115bdGTjRm1vy9mavDdzyrsRD0LSFzbhm0/yMVT8nrr
tWM2HVsPyPHR7ZAaC56+xpt27DmKwEC68pARPYQZvzzFzbxQIiMOvCMBgL8Kd3QV
cGNJllCyBX3K3FvLNzlhHkp8doligXeNGM9XyKyw0sGGhTRUs4v+k/3zHySioRD6
efz273tOjbfvETd3ak0R+eiS6lvU33siBDH3F+aO/Za1EIxHXNOZGn4yDCanq4F4
COTZgwJjUP0SNQZTqXeWBLFZGvWL1F7jYjml9XklV1TwsBB08S6dE+y75My4jWK4
1GrmupD0s+Ly+cMIaxKCTMaflHuA+CJm/F+oelCcsIZaa6tRm0ZYxbxd4+9pxdu7
rMl5x4C4UsiCHkmJzfb/SK87ipZ0iIIYF2Kpqrr/rkS119G2i0+afO9AHJJpILqY
rjuKSAccAwmOpFGZiuAK/h8ZN7feuwEMDmLPLd+X4DbqNjZMwKwInfjeuqxYIqls
vp4sMkNu7+IP4kZduyYoJLkNRfgSTd6IDT10AzvdsMkzkHdpoMEuwu0PPwrUU5Gh
0OJ6qGkrx10TwFKI5MG/H/IJ/i2P36uoagcvItTPBku1Ywnaqtmi1SryFVctMQzy
X2U+qmViWKBCo1v2a6/PY0MUj1526VjGiUzNSjF1Gxc5Hq3l9jv5qWDDkPhNalBP
EXq7er0iwpTnKxZQIO/91MG7qFuu2LkFXpem8LKjdDvnmhTj2UJRFSvu+FUlzJ+g
bD7sBOMw8Oqm+SiiLiVuZQPaphQW5ZorbhW4p5vXwlcPAz4BY+pJt+Ie1CR4zGU/
GK7kmYs1KAUgJEXDx35YUUw71o17+yasxecPyzl0pvSZ+j45zmi7Sr1G5VIrJ6il
K5On6V2ILts0BahuqnmyQpJsI0DZ3oV1pztsNwcWQAejwNNRJs6pMh0BC5frsPrG
z1HI8MHJ/CmqIaFmS2c3BY4kw1ysdb4xtS+is8zjR88J959HLFMGbRpGU4CWMppW
uYgsmK0ZKHyNjGWLYoHrEc/juYd4CNsLlMX7+eGdZ2fksTf53EBRv1z2KDXeCe8K
r3lYxOiEiYCnzLmu+J/R7kG8QNmK2JEkK0khTUWNxPfh5fNAVELuOQCxH1mgRP4Y
SBivuAgedY4nHm02eBoXOdnFgGRvq+G6jjpukk8e7sE6Ro3ZuKxkWHbcElR8WlVg
DWY33mDkMc6pkI6J6qnoG1u8pJ72DCCrImG9f2vN2v0mCjZzjPkJ0rGhFQeulfnH
fGzmQb8j8WwDyAme+tTzYYHmq9nJmbPbBTlLVivuKQE1fFwa0LLnoQ3PMYYtxoQ1
tvicpBmW4/53JScc6WVcFc1vu2t7BG8AMsgoEx6B4gRfHxVnOPfPxns/IWPdVRc3
bEeMK2ceka53UxKAUiR/ceNOafTjOp2UNI08Ph9EifUz8wFv3Yft7WSFbvKAe/mn
eqf1HRASq4xhemdiRJnc6MvufH2TOTXaRT9efVK20bs97aTvD4XwHQWnRoUNrQQu
qXyrApKkAh9IA06MG7MUjNMTMR3JM313M/ZNvyEUSouKAFOcJmJppE+ZLH4BoNh9
FQINA5viEahUIXSe3uUGugK6iEgX3e2QnXKC5i6j6t2tv62IKS1lxdLJihC/3Nul
cy9rOfQOqwBW1TptcsjvNBOujrTUcItanvJXuqx2+cSIObc5zMvWyJOi4sryxErj
vgMcG26Dcd+zqDZe6V3HECJyqcbNMfmldTierU4m0CRl/jLO4vEXJ31LCLEBOTag
gWFRxOUddT8LRGxai1J3nlvs21+f7ZcSgogtH4FHIXlPvvnx6tCYSvAsYBRAFo7R
CgmEkyQ18GyXHCu31pC9s/ZZJ7RzISGZhvKXmaVUNHV0oN7c/fIkLoeWpxQP+R9g
2OduHqcEuqnwerPhgMy54sKkeHchFd01Ng1gPBqNPGt/CJntnK2hawg1V+AeEkov
QAJVtgf7bSwhYYGGLj3VwSheTKQS2wQy7scsnsUPFin9aOAd5vWwQSpZNGNtnxI0
/L2qp0PbHSwlS5iM7KNdD4Vh9fEEOJtVZkHrKr5FghEAHT0Tg4VNwdTpWyNJx5bW
GNAnZ88uQqXzwgqVQdPEONSXbB3myQEuJHdxSID7zIN3IYLNeTgYSB/HBqFTPiHe
XffxQbPG4f5uEqfjllwJ/eSRkkkcBFDywhl7Z3FWpRB1VTMIwBV/kcVESunAZVA4
TvJvb7tCDXkGAcBKliqN6BtZYOfdKs36waHgZXhIIKeKJT7Hv4xUOPr2YTQxROpR
YoN0f04OQa5GwxAXkgBInw+2BixtUOJteRb3W/3tczHyl5ChaG6gmQAakDhZ1t0c
9m2acdqZjPZP42gMj9VeIAFBkmdiAGjmas7UR+K/6Y6o9vHTBLtMu22A3ZRFV04z
hkNSztMSX65jlc5yOjvoxgLA/evSs5vk82PpTrsTsBcrUru29cQ7mocd7E045uJC
JfJWDbdoC6nDIVDvtxGXA2L8mZ9j1juWj60MDLz7DiJqTLbTamYCu8MKVNCRX5vq
umd92fWY/nVgnCdiaDNV1Xe2eUuA3fCRKjpMpW/HCeMqngpZ6KoxDpygB98W+AHb
3fSXy4GTIOsMGib4Pk5gGxHs1PEYet8emQK9EU3ss/L4eNdxOHbyfh6Cb5bc7q4F
A6KNsPAOvl/VXCBkNqWGnxOKXn0YxxeFn5RkkHETE/iR4A2BR009sJlxQi5Vz8Eg
bjbcpGpJTHPyO3h72PJ3246KQcb84sy9lM4Z81VYx0naFAhWZp58c9VyKaBJPZYf
0Npg0uPFUAkcHZkCkqorPmogLHZOcO0TAAh80pPNEBBVbXZTUU2PWfwSvQM/tf6O
pga8QNlgrCZk/cXQi2uP0mMuZINrlQavIu//6EI+caXvgRs/WZv18AzcPwfegHFJ
ONFO3QurvJ3pOJ1Q1Habey+esYQ3VP4kQXTBpqLGP7vVMbRaI0IXZid3Hbd/SE9J
YHCsufGC0fiufpIDKvdElmfVkhV6nZPXn9fAaeI3+fj6P9Js2m2IpkmzsFja1ghe
9i5yOwooTOj+jvONgFrRWFb0bs12mMLyvggDuYkYdus6GY5eJc5SvSzzkVywFVxI
GAomCpwNgskq2BPIoUKFyw36X1eV3JusYXOTMQlMMVyUddjcpcfAb5VnZcouC9El
tMiZUoY3d/3X95wSEzKO77pIlXbEY09cP7OVOO/ASKSAxoAvxd55My93SI+2TLvg
LZYTjYal27P0ZS0I47Se+HutRLcbgMLkOROi2kOxTWTDIoP2yqh1LuF04qyBBDdF
DfboPPhhYrC5IVsI5ksevwJcX2tnBfyH4uM70BgzYfF06UkOHyxzZ0XTOSnsgPRF
CT9ywbsOyVEm0YhEqD3oKvX1lKP/SRIyRXA6k5gySpJwb+e11qfwUlP+iPzjcwJh
xU3jT4dm2smY2ZTQWscUEMae4JlfTv9obV7vdFDqtehhzxhr2jwDKUSjmz1geqJ4
e1mcagMlA8CWoZynqbNwN88sPZ52yxjK9GNHrUwtxjE8RCfWkibkb8l5plp2REMJ
TFbKt9q8h+yfOLYv9bWMNGmFdUX1O2DfZGBJKXA0aOLHCto7P5nN2Qtt70CeTMFg
f9qt6ewk62dfWyUQYBg4YfYP2tqu3qCcq4lNKMXHr5+xMUj/GBiK97Tye9BlCMs0
zzU9M2IPpYuMNlLrA8zdrZSlxNC9CQPDvcIDP2PuHQj/LWpqRv194FfNesqm3bVr
hT8mzkSl3I10Ngb1FDBeOePB60OrcUPFaGJx2G+zHr9kDhMjQ122CCJXvTyluv5l
jHrMGredEptjGTSbFCaUZykxI17ea18MKWVukN+6bBoeVFD+ADjFyq8QaDDIxgqD
aRy3mkwJA77OWiUV0RfqjIm0RLttFe4iBTcuf1evU6ITf4NgVKgZ/ZanFhdmXmqq
lRBVyCY8BMCoQyqxnw5TrWBu1yYjJytIwzQYCgHBE1MWn7wKULsbwgkura8VaBsY
SJAfrGSVmZUMXutX6+UCzvcezvSkLkkghNULjH0B0iX3YMuaCDxqMutsWE7HrSWe
wv4wc0t/DkiP0qcZMi87qG/VyzLasYKwN1j8Tea0wnATJa9LUNWR4uuC8VJgrYoJ
+HCVZ8IuJbnzul0ue58Kf7NxWFiAXgCXFqQhwffVuxvN1k2uOWhdXKaHX5QsIZWd
banmiAc3rIGcctGEWC1EsAaQWFV5ZuJYp6duRoiTjVI8gdfSkrppPBeTyoVqylov
++NIoSrtWqK+GUM3gc8X3sDaf77KELE8Azi32ryhSr8ORgbZ8ftt7HZjFg1b7HiE
n3rVyNlDbJn2S1OfqXBBQ4dOUKVq14UsS56mXxOcRnLclAIYPSumhxtIl1Id326X
EtcLvk4wpPCzuIz3mxyu4qg5AAJvuC3WW6KyPdJ6sCbUVqabzMzbsxEl8CwQzhJV
yy0EGhFointRO5TpJ4ZGZ0nPwSdmrl/BxVAZ1CN03mPVe0LIKCsB978ZbHohD4TH
fXuVEspDL9HeQO9sly6uJOlhtwpErZKd0WFn5E/G3+mQ6QE4pDp6vRI/FfBd6PXQ
0QrahN+MEDCLvUZN3OG4XaY6HExECK7yl3Tto4qohlYfSaCL5U7Xq2kD+9CB+mx4
wY49Sa3dimrY3MCIRh0aWvJAklKRrN8Nq3ets4E9bPWyU8WYH/rztFHZf9O+M4T5
vDr5y1OWLiq4xeS9PzswrBq44Ahgm9iZweyw0YrYMTsWHwKNV+E4/TDUkIBqhAuI
Fr91szQ6aqOFpz4sQrRPmHY3bkx7C7iNELsJlQfLajGfiuuZwZLXRXd03yhm3Ntk
K27mXpQwsWIMkrvPfP9JbBF6xB/LMwoq3Uf5hzZaCqxl36WFJ+eUasb4+1QgKL2i
CjzCzsPCUOrb93VH6m6rnnSHUeKLjfDWyWkGU6KL1BHUtxsb2l0fo3Qp2dcKY9jc
XVrBnjV7Y0XWkgO+pFC7TxIPqpEYDH6Yy/6lVU8J6Y/xW6iiL9Fm8cxh3Au1FHp6
eBr5K0YYEZZluD79Z0zENsukQ1UeAUsZjpLDj2ehGMJTtcclcnSjdDYVh++xRfNB
9I4xzGwE2/stusi9BU07yDCPTvj7ywGs12akPhxKDY1OS7S+7ARlOdRIeJxYg3/G
K0aEUAo8pOMHphp+eKyJ/6vPQq32DmZrEwZME3K9Ti0o0hVsecQhNVtNqlIrKMS+
iwzJYaI7j/CLQl0sL3lWV/SxB5WOMVvxgtDXRIYFaConKZEMU1pg8IS/mT5Mwq+y
FxjKUhaR1sXityACvk4IDOaqRNhn2qoTtsmhPLRiMQopoMqLH0saTL99Kg7yZrT7
xegNT7qKuOwvgnzHAsx5ysO3rcVWZc9aUXig3dwDHDjS8alyNzbYy4TtBrFpnCyL
k/h85IGgtabEifgdCtJb3DSmIJhad+TUCmNNYVlBZ89rScwTPL69D457AxeaqT2E
SClYhrMOWtShRzBytQQmMhU6KtvWqdoEtnCSxYHsUSIrdQdAg8jNVH/64xIL8odU
qq7TBxEqSy6tE51oYvMY4a98oYArB6Vi3Gt/+4/kt9PrT1O2HyNJsKuPAFIN2VLb
NaCaboKr16DQ5W1pWr22p7KFJMmhKDXejOvcogU9yO5sk/MLUPr7DNvIAVJIZ+BZ
/eEVAmGusyO9op5KZpAHPSnsEftWTFmyeGO4gE8wnyrq1ATAFfgOYlwTvuVjtLOR
wndLSRwwUlG62HIqfGHbgfYB1aeIOuBgyPCPdCbdjuHIBSXZ62QyGF/mnYd6tb2z
OTVKfZCMlTVMu6TiUZmQP41X7eEqWxAeEw9w9DPgVDvtXIYwwjwsT/b7bbaBhoW9
9zkLj8sM46IANIfwzvBXKiK9iaIFcngm78NE/MP49l4BpEn4WpgqkK7olkJ33hZ4
O0u6Gpi+Ghb1jpY+pLhnd+z3IfXrTl8cOOyUCjIPxCs+XroYkkPXI6pLQnpXLHJB
1zBdpEE25v7JnewwHQ2EQdHA3wE8Aq4BZVUD75zSS4mPu0hIpUvd0HT+BSaWwbqS
Un85sv/C41/uGTpsmoEUJ96442o3HgwHnl18c1pVKvPK5weK728PWBpcEf/n1UyP
93DB8wesyraYxWQA63UwyjxR2DOXaYfE8P++Uim0pvcr8R+XeEc4A2QtCinUxmXm
2+GVJyBku/8uDAD8jPWYnhCoNr5ATIOF31UH0jzYHCgyPB/hnX6kHg6GOUnYLrNU
h0wh7yofGswJFzcux3j73JmPbuZ92/C9lmb2ieVnll5da2iO9Chv7oltsmO3h4zS
xY/IVKDIQYXUID0jVCdxIqOHmm8VPTPGB0XtslAuqLcSlLdjS42y4wnKHAbXoGEQ
lUEGQdmk0FL/XVNzkuWvd9NkqrCTMdKhoDhUHLf5z9Jho6kFweIm42B0Cs0QTGH/
46xPI4DcEBdWDXrQKQrWZdPWhzwfeh1t/GyLTKQe0EPjMtQYUX0oU7huEHaTApWx
smawTxOvIf9jHKItY8mp0kWHFBtgHVE8iaQb6KwrWjlYXugTezu0Yy7rLWlCfE/u
CFHNVZwWkVzWl1Lxm7ZENtvsiaMcMRBeFHMn5a918uyByDWw0PPLQFKtAxcXWEBt
fAFtj/mhmdNjAZ9NPWJyGhqhwZ9SrLF9sw+07Kl/AcYlnwqv+ji2r5iiEJUYG/j/
Ps3t5MQ9ZEpOxdBKoDBmiZ+dBLnEiG0BH+fLWJm2iQi8WTZVVPCgd/+/7G+9FV8Q
9O4y2G5pYF8ngwAXq+IehaV+F+rwRlcd1hOQamhnmTH/lF3zuBTGNCL5B8pykxjM
IgWQMx97get19UmueNXmG4dCDiN7fgNRxlNlhxvzj+VaqhSJGJrMkOhWnz09Qxd6
KKZ1OcFAHW7+FdDPb1gwgDGoU2opeyZvKfrAI/NykjmgigA4z5QdIsPGQ4hClr5k
d73Ks1/39rAEA0f5guNXvQvQNBj8pbLlKVk/h1RljdsXra+3xhDZW33Yk2jIhR4Y
eQUJGnhRW5t/rNnza15zGRsmBp9MKFZ+IsIFPokqRMRFaN2Dhf3OvIQy4CJLeGpD
JUCbXWGG9B/BGjF8Nka3b5huHRsZx2wTMQep1Qrd+XqUEkmDq7NWq19HH0Egs1iB
bi75RPNtjqPWKfhfVVfTkvEaL4pdgpMX4rdnXjy14m1FgNiYmkdYWAzQR12cFOhQ
Ggs91ZT2xPb/Wpktxu/XNgDYPUikddC4vSkPuaS4JW/W2lD+jIAQRnbNJbEQmay8
VaTjlPM+BTksLR/Tdk/X8Swhm5pYYdsTYcH3quoP53KHiW5mmD1DgHrffnCyqRpy
lf9Vhy+mMzNc7hxkKcp2WUUyylzJI+FL6yNzog6Rz23XTE7gVy2ozO715SAbJl9G
WPAmER+DEWIVewVkuHGgon/BCYtPQ6aL8O736/CTVKYs/lJMVY6G63W+clMcyaGl
pM/T5bQef155z0yEgBm+rQfpmjjTMKnbU6D5Lp71hoR7L32rfPIQsEowhGqb5Hbk
eqqfQ8QKTjZk/3UttYD7jtT6QatHHzXlhonbKd5q5bOBZCzVMgZECkaq5sdchSWk
pmgq8WTjYNRd27LhQqTtbDjQ5+lh0eixrvfc14QBsyc1sHQMmhp6w2phpSCYPQrp
p7a5syj7iKvGxUo2v/9cHFmMXgeAISCX4qslWwwPbKNiflbv3QXXInqrjh9GQi3U
TaoHbbKCBfy/Xy8WP2kHLObXespvn4CB1uXLfFB5A4zsHe0v3VkZ0DBmFqaSWfJm
iYQRIC1ZnoXidOZqE2lX0yiiuID3iWfww6FC+7/tABdEhbdo8UndPz8HDvtv6aaK
qOCC2mD9MSb0V46r3JIxAfGRmIHileJ6xA0BOjL300AqszuavWcJyXjv1CtHK7uZ
1EjMB/x+3nn3hWGLqz8prUcYC1SGFJ5rxFO/n5EBIKB89eUX/PVoSM6OxFfUBNX9
dACD1tHGD1SK7KlODBXnNzwIrD+0Mqpox6KE8wFB6no4H2exPIiWjZV5ZB8CrJaL
1RPUyHCmeojyy00+4ePT7qgDYZdi8pC4WJq5t7UE1zysWgOvUuBVq6bW5pe55RUo
QK6mIjmlMtWFyfFqQjxPs2n10eSqONS4SHdyebX553sAV/h7Fj+oYK+se71R5Ayb
RVlpNnza+NKu0qg0q3EW1tub+i+GG1jVSDEZcDxbLjgqauniTV6lOpyHh6UjbIFK
D8wQyIOwtJtEOAcnUI1k3XNM0yCuQo3bnxsl96IwEjHpROjBzsFpv5AmymmuVkok
nFaoEuP7fjSdv3NtGUMGPNdt8qNh1Dmr/O2/RK9Nz/xq1RZNFb1GcPQZjQkSVqWs
n8UVO7M55pA6LbQrTDkRHTaRvzdW5W4GeH3cEB2I/dOFV3NUb2A/A44u7U//RfT/
O+xN+FGH8eJV/VEwqcQ09uYaI7m99cXAmt9hmYYx24m40VCi8aIkmBM4C3149N5I
c1kBKQyNyfJnFMRcVTbhN63EdQkhs5+okvo6mYveY2Xbtg/o4tHciX0khnOolRXR
OApiDsqE6DVDqIWzMS8ilBmPKATN9QDS4H9akpnavuv/nk3Nf1InNVWqoUyGlhGK
wcaRG/FXGZ1aqpFf7mVBSwJGK/p3IbxOZYWCLkn2ase4vpDYRFrky8k3LSvhd1ql
cUeQZ8ta7MF5rge+xWqKFt0FVf3n+jH9yJs1+M8QqXCTuh5L2pgFGbpEbLJ4YO/9
JwwJAKvMbK37RSLyD0FdGMqz8MXUnZsxuxTN2iE+wUKU96GMIkLvYm+T6CF0XDez
O40ip6DQMKY/K1m3FEv3xvOoKibPxEUN7+MDLyE7UP4DIp5wncvgf4xnS4gEcwvu
EPf4XniGmlYOx4qvKk0PRf4ZmlJQ/Qyv7oigTlvaIl0T0wNm38n2sAN5KgQs5BzH
D04AhZ7tcbwM6otPuNCvHRopNKyf4t4FA9zt/0B7ge0rXg4gKpxlDHVrgYWfxMad
A7S01TzoEELjs/bc2UiLMOvBp2iydCs16uL8nGurYU4ils7AMHoN0gD7sus6HAfz
1AeGtm/ReD5cXUhDUKMfEk38tT2gjVyvCyfTCMcRAhpcSYmTx4AGMI1tafcoepjG
+fmcpaPXPouwNYVpVU3uJF//o4D7R214isoINwXXwTwONjyCToKXgTFLqd3Uo/WF
Jkima6WZH/MJJg+mxTihcHHO8Q8dCNVrGVey+4pH9m1q9tz57t+4TYsvoHf5KVQ5
Qx2pqbYFfaEhNzgvMgcwC2AYvnPh9Fv5ELe2ilyBtHmwHaUH6fuDt+xSMlKq5a/Q
bj+7e/iQ2rap7hTLvL6EEoWBKA7hzCZUELEOZyl0FSWJ5xyDWG6P6On3sWd6vgKL
tY0H0w2j7zmDYPyimeVHl0JjFnMdwnigJg8yFrbHl3/63wY8EmssRhT6L4ACr1nZ
42taMdxsld5Kp9MCGG5UL87xweh6juIr2Vh8PcSYW2iUzf+h2BcxyJrwDHEmD6Cc
6if2+AEPdWnCsg5KG3w/d+NQQ9BTSEGDbFitvwydXAvlzb35SHqRq4pWzFBN0N89
mVG4mghaqFx6R6J7KrmfvInGyGddCgwouQI+kDxhm2+pHARZ8rzm7OWI8s7WEvKB
+HefB7ORt0r31YCgVOyCnB5DcKTRLdRCfzdPjhSSbxYv/GwAXne7ogNGxda7ruBu
lQMYp4nfnrjAdJFjLXW/heIX3WKOjZHOPDfNsuOtlGOxnl3j/nZH8/y87MSjS4q0
TxUNMlgWwqPc3Ac1+d/KhMCCc3nBpOGr0gZCndP0kUI8fWCfCUCkgKfzexhgWKi2
G6je/e0AUG5VzLw4K4agSlxBWi45X0lSWE4zr24rv9HJ/RG44RwouuoupBnTCzKw
7k8Sdc2wK/JJg9Mo0w8YOq8zOpHhw1lmnt0SayB8vytj2j3OeSjIQSmGqD9bP0oV
x3KquZqRDDB+gCuUSmGv2MKEbIiAFQZW+Vparo5smWgpw+eHwjSgK5yhMJFcEJ1E
Fv4f2uwMJ7Fg+QFzV7AOHKqUsadvI4sA3pt38K84iYdQUYbfFxeQHLj44WxQ+qLQ
fL8tV6imJ9SZrJFEdDItcl2jWLGxGX/oLM1IbAoyWb2hHy6dmUuUO7x6FLaf5I58
RfLK86DdcLasv7dMm3BfbsHtmQzwXA2w2QkblCthGzswA9yHin5Ch0I7QDKTszMj
4uD5/+m5ThTMsdzSnCUw7t1Utx6TbUjQlDz/udcO4+79de3bKztNdu0RrwomdIHZ
jDsUuYMLHsZe6CfgFf6zShXkUAGZ1GifshfZILj2Nil1IAXIZne/BPjYYzl3euAi
LSvkmyENrq570GXjd/gQNloefFQJLEHDtem7/ivmJTQjC1GPw5T5iXoLoPuAOLm/
HqW8VCxd8AW1oOiUAi/MTiMrBzjgsZ8ZG00L0iWM31TB8UcxJJfK54gg8udD3r+4
Ndxj61L7n2bwiAsONOOlq8+Zgyy+CvuYZfDI84yesK4qHn26wF21mT74uyrBNAwU
O19QdLlZNNEZmlsz2bc+A1d1YqnoVss5QJMytxjxIgAqY0qOKZJUXj5CpIt6IYsT
D8SmIqqDXwyUE0GLtlpu0AtHDE4J3WUT8ZxIwieMRPSXmEhz1J4g1fUJDYnpSMBc
VTNHsSuIVqGRAC7lXhvoGmXQar+zsCQRnppe04vbPPNkaXegmhwLKbjkn9q0fwEw
EOIM/nKeXz32RPlNezY4KoVkGmQlDd0GaY+pgeMKj0B2yYm+Wl6i17HxgXGrVhdX
vra7xmTsX/7qIjkh03zvPtpVx8EqcLN4Sfo5+w3gOCsjm/9zyS4+ARmLd6eOKk+/
JIgCx8w5iTbfYnKHl5RIuCtSY/Pg4z3Nc3HtZMEfdFr2ZUPNhjJsCqoOg8Pbf0OC
ufbnjYbwUcPF8jP+OmOIsS4VllWr4RDywHngHAaLHyIr4IDmOPsPQRSDO1RsFzno
naIN9+71J92Icwh8HTO4AwqeHj/hoi2f+N2u1IizW8aeB4Roaf+zVTFqnZt7GKdE
LILr1XV9S51fUn8vVBBNq6iyVtsA9O7LHBaU/Eji2/EnEPvq849vVLEX3egwhInD
L7ExM5q00SbMNpT0RdphXyAEtqiOmGWCXqVYVPbCvg7eURktc+crPWvutHTJvvJ+
/dmnoV8BAOdTYuwLuL8VZT7oBR90yxHgV3jgeiM/j18hUzLDQcQNCopzJjE+srmm
g4tf2X7OCo++0sDuBE9ws2BOCzvOfBAffZNYnsDVMsKE5q7tUfErdkW09G7OzLxp
byWzeYJYmnHh2v13DvQqgpcqjoGgTwI1qdDn8vfJSEg38FXqC80a0jdb10/9JXFE
KtYlLvpsojriM1LsS3I+jhFWp7PVbssT+E75ijIYA/b7+QgDmoxxQMysSO/gPEgx
3nunu0ap0BUuy4BC8EFsQhzEtl1QhUQccwfnn3kzkiyj9saUnX4+ZaIAS1V9l+0c
h+0l4JiEoClpQqTeht1PUK6FC/UvvF5t6d7zSEUgrpVqJJpzoWekzkETqX4PgwjC
fQnUKjVz8WYdxPNEbjJhR/LazcTLvLbOmllH3G1RzpWUs9a9kMIILnvZe2MSWwwU
D/mM90talWlcuWseAbHpyRzXTdF+CyNKkPKrEonynf2UZQjMW0NdYmiBm3GNxpnX
OJpGBYUv1UYQDTD3eOWIe1Fib0Rqq6hVVnxt5S3G3H78QZAt8u6z++jbrFpKIIr4
w7tCxwx5DjtkXUac+mCrx3oAYLrUf5//37LGgsyJnhsEtE0q6/mhL10wywngVMcx
BWyykOEATud1cAnTfFG0pxiEk/6lLDE/tr9PXUO6UtdD+mpEO2/ESYHywfZyqxJG
gaAwQvmA3q6PSlEAVWG6f8ZwAXwjqSAXfGpngAH2mraQvuxKy5mToRR28N4NL+uZ
hzEAdE5cb4QZFC4Gs7zQZxRC1NV3+93Ax7vt8PdHv5h6Ssy3FV7ex0esYRrDjnqW
wvamBN+ik/+hxpARj6FFbryDIKcAr4aR0lcsK3ACZ3ifxpYUP9c3Oz4PPSUaQlp3
ByhhuliyYf3BsqbjpFCStJBHn4PLRqa5N0+rLDxpL2PWZzie3svqI8xDj9WAvE0j
2CIgjTpiMRXtHowprKJMuftcMtgZ/CiusPNnGwmeB5jOerGtPSnRMBOCRreq4ubx
EDZBw82095RdEmnirkHUPI1SZjSxsEP5vAllGC3EpSD/bwzqCllRRIx9Kumid2vg
QimPq8Ln8bGDRNwZ/Z8a5pNMxCGZkZFAIEfq0QIQNgZzCE2YfUREgKmuX/CaEAor
A72SlIIklAFv/QT7Zr+f/yGIvHgJzXw1s4jWKe8W7OCAbXLhdrWH3XUOA7eI7Pii
CYvb/bC7mVjmXXwwQOf1RUw9jhKMSGlkmJROcBBwQJxWyrdw5HmC5MO2Xr+7SmqM
QREeewUG67GdGI/1EszzQMXXR8b/P9eFaHQaEZd7O2umzRrFP5WPfV/t5DZ/KHN5
bVRvhCrKp2xAeYr3KaDjjDZqwFFFn3aWY1B/89ySzwJgwLlPC2Mr40PtWRjTiXxC
sds5y5/ksMJO74TolyJcwjDPpvpbM4NjtIl32Pu8OysHOZaDZAEOBYFj1Y8NgGfB
abUdtFDLqCOpXQwFTkmL6E4dfuEZ1tTaRy8b/BH4DM7dWjvbFmgJPNIJWbFvPo/R
NBB9T/mQBGDWPdq9LBwiHjYPQJv76FQ9VC3oqTergJKFO3tclLnFvJiv7Pxby/f1
CStk7jw6Lx58XZN0I4LMKOHBwO+VQXsSqH8Vwh4/wFPlyFid/5X4e80aUK8JQY0h
oknBPh4GnSwyHta9PesP5DPt4hJBJQZU7mFH1p0Gedrvu08h0pUWCC9NKc8HrB14
W2KuQknRR/8r7x/GDocxllIClEuptIWwLkUZNZbR+WqEV4g1wzsi5FAg9kKfzbCe
6YAoW6lwXXgizdqpzKpdKyyNxvs+atarDrJHmfigLdtq9orND2dsMMhW/2NzKZD9
9ETy3fKKxkSm7PtchPoyXgvFml0YhAlfrcD/N+uQilrW7mnDxrXM+yPjSprto/3b
8RIDYj1d2s68jFUQgFpa458FE56UuRa8X72qIu1Ip5T3CbNayUYZk0OU55A94XBN
9AYCZiwubY5ojhrlMEXBC8qI9uOBHMsiAGCrnJk0SSP6Mt7voy++Lfc/6XY7UNGC
GwRqsT4iKNTgDBHaISbGHzrOPvK7gs5zLUciTYJp3VL1lkx1agmSXqZu/mGaVmRl
qQhITQoBdG1mpdwyEKjiDxu24s6N1a2TvqKW4jTB/t1nQz9gP0tzMlmBVjue4xiB
2inWBevyqXQG1AtKuUAV1jnlWaNxQrMMEw3u8PCpMm1RHR8LKbLFabk1GUfCnQLH
YDwE7zYMmkSVWq5yLBmAZjvEkFPzieuoXYU5lBbyeJM6t7NiSVM7FbaGRGN8lEg0
Blze02WX7KDvzsnIli2e7/EEwN2wKPE/9+/3tB1/ebSA364ezvh1thtahk3frqhv
kchYuorFJZeg/Slfw/VU8hriOLNqdaA0sWBabXdBXdKyfLOZZUFCAHmKu/nBgDM7
qA6Y9jDKixLUFaOACE1exdc0zSAONMA70PN/jWdT6K3nmhNd6NUfOpCR9pZEGqpw
S3j4uXb2jedWLDdzoIvbjLJeguAcyCU8lDOy9CCLqbbsZ6x3FIznK0BRD8nf+oaH
wsng0ZkkjH8eq66LdPTy9oTiflNDW3QCLG0U8xzusvYlQTWLykr9AHUcGyx6cTNB
PJ1vPnatf4BZxCjCApWncUHpZHDzZAfB+8DUfZJA/djZZFklGllEbFHS3yLBGe7l
EPLR8NI9G4JqgV2MgSjZB6T9wQr5IeYiw6pf0We/PoMgi43oFVu4bX3dbNBlxCqL
BxoHg9yIwi7j8ItMZKEMrHQCVn1jvLGXubNGC0/whvRiEtaqiG6RswyXoGienyBa
N2k4qHfCZengNKL5c2Hpq9lZpVCQQI/8B9Uoj04ZqY9mH9ceCKE5vMaSfDN0v/In
c8xWj7ulCZFJRo59ObLJDHjkx+IEk2y8aU+qIcLV7CzXbxaFWZkGewls0jtpIPPi
y1yo6dI2glVgePK8JJ/ubO6VXjLum9saer/SZxbeKc+xnBh2qq6kn0FVmMMn1cPx
by6rYp7KGaHq8D6ee7hXu5oYJRzhwXkh0ySqv6KEOc4/2Fg85zjXBlmcdA2f0Kei
Ti3xJWfmqsfOcIHnXr5ruyK08qwzRocLz8dUq9XTotd1Bwmv+yhBp29oHbBNiJ/H
Pj2JBrGSv/NFI+4wzwHI529N4HH2yOSFKOw8lTsuUYCNLcqBA1VnyDjolaSiROPp
ajpTEweAjEYrkXKmPKgtlnnH8KJsrCtssjYaOw2iFyMkNh3zqz+kmC9112qxFeXt
Nmo9lDvu8Zov6NI2CabyRF3O5GCiIszTej1gTWWtqZajBjywAbdv4iK9481Qxmj3
JPB7NkYicBt55xyJ2PNQkoJtHcEuqatZPRdSjQX31krCqVpzr2XlkywGTX1t6le8
TzUfT5vcsGeeVS5HvlUvi/BRAtWKsfifg0O8okf25uKyjSZmKtVhASFCeYhkC3uK
2p1WdxFiuj6lhEghaYYP9ucqL9uCvTEq2EXonCHLohcI9OdBXc2lxrHjWUrnp/8Y
xTJFV76S/3OvC02cG1i2DDiUaXW5OMfH37Aq2a5veaPs/VnqktpflVBLgyfV+Lst
SbedDnBlD3w+BSs2wonibEwWJVt6wAnKEwdtAylZX2uSmw6NWLdnzbfzUTcB1O5Z
Njz4SO/h7Y+yKCm/o0eSLYTAlJxD1Ie/KcX1ZOeJFaMZe5qsEUTApyLv95uervxf
NXy8lMCdYJzqBKoVGCzY1MCjsOzuc6G6sXX4qyottEULuTO9VDl/vp9JaI90NRW0
z4WxmxUSddLsfJDb/XzLI4QMNBP73ZNl8uR5S26Oa3q2azYhaDHhoVeSgTnjjZQZ
zIBZYtHk4yj7ZLKHPbnwl0OTZPE2Y4K9ODBIW7t9JIgFQcpyh8ZLI0rkl2i09lhN
Cm7CON2lrTc7oi26C3OACS54cJNQHssTlqwgHE99zhCW3qYqbJ6I2D44ME1T4zSt
KS0x+446wpwtmaMsAoUy0QBQrk9awTARW9Mk8G6KWhqT+Tp1aN9x3WZ0AgzN5GsO
9akWSygw/FLc+e1HD3YsyPrcqlB0mf/rC/eyAVpRBHssARdhED5kMG1g0wYBTd9w
K3ysYqnNo8EdzbUe7osRSUOjlUWN+H2biE21pQedPp6ue7g3Dv+sIhDwWPeocQwm
Qhvj6oNPff0j4PP1I+8yvEoTsjhwpR9hQq3QPBsM1Dv6ACfc6U1VA+q0iP49fyW9
zgeRaI+iLyxfPYpXAXRaJaCCc4wNokmfDMks8u0pGLDtR9rXynh0d/AXpLGGQn9s
zIzF/vvHeKET3EJiQp/GeGLVm2VZEpVKogem9OgYmn6lWx/qPdpqQJqw1zbcJB7l
OpqHnyXTQjyJAsVcwDgwMNYghZUr0iaesBoP6kb/HteWvC62hlz/+tGM/DZNTD3g
ooPycY/bnBkSw+mWJrFG1LGab8nraQqVTsmrYDidGgeb/phAATMGxMRk3VS9FCkr
ZsDcYHXoqo7ikQVu56JF7x7fdu1u81KzO57QS9V+M8B3IC8j3dU/iL+TqmTl2I8Y
Mw8u5k/1+8GPAFMz3GaHHpfqPNozK/n/xP8bwqBuDBDaSh1qnVrxas7ZNFYcumER
qEPVCFJ8WPtJpDdkqWXH+z0geGBbuYBKL67YGi+aEieY4Oyc1cK6fngwya3VYxQw
+m0RNl/QTGHwCXDLRzgzZ8dBzkXgkniyS09uhFa3wNuPfmFYfJw0KGsUbS/Yi/9a
Z78Q5Kha1/ST9RvaRt1N+iEhp75lO1eL3hnYONYkwzgymAYI+Ho3H+7sY/O1pxOw
xAqH6dZY7cN6GUkp5w4a9LyhPDGhNFjrQzuwhr5lcLbkIzlQvbpEOYfRZ+Zf0TUb
rL7/6/829DjY0yGbG/TRiK0wZ+ZREpSq5pZBGy0n6xQt95cNPWJuDK1Y7f3QlxT6
9fQvC4Sulq+3kM/culGnIRhGnoCEYTOjBOHnCF0XeqoGaXMfE5+JLBGkfwfdatJP
OUT+kcuKPsOMxJgowpJcjnapmPIXYr0oDVCLU2kd3Us78McsRX+IFxuj+Gu7QeBI
5gHfRbEQMq2xssxa+M2NSX2vcUX0L8o+amLk2HHOLvxRBmZK/L8crzX3GuSG+cnA
vGfP0n4tVwihWwvV3Jf/P7uuhAEE3Li4hJC4t8JHWg5TuX1RzZExLqz2d0hu+YRb
+DSELhpND54ri92VtqwTvWbLyppzts3FK6k8HZH2/eAEQ1BkyY7iUv556Z+33BKQ
yIi9Gj0giKv9N1W8T4IPzuzi8oN1RnrZRl2hS8+gJzIqoSlQ3trPJCWWDplYo1+k
LAncArrMV5KjRUHemyX0qa95ehjjZNWOlyhJQxE1QznkgDj/GWD4d1Svo6EVkYpg
vWriaScO5mkLAHJNYhFJlBgReGY5sHRbdqz4TIg/69aiFvbt2bcO0B9eOpt1Zfay
Jy0n6kQm2h5NviJqeZS0bL+6PX2wSLbEho+EfIjP5Uv3xwWk1zAOp8fH9YC1NteX
9UTxYgRdvgDVFhZ3eeZCDeDde8bn8tWhpPuHVPza3I24ht1BFyS+f9R90o13Wl81
0IFnL+iEmo39KrTk76dJaqjOIzteJZC9zFnMiPhVlJXX3Rksb6Zns2QA0qRbfsQ+
eiG+woYOMNuQUwd0g06L2UMBg9UBoPeYVmtDvg5Rc3yJ5Urk0s+Yk7aLlHMMvbAy
OwcTisfETRGPgaZYWKRcOCl22PHXaM4P/XIW/PpPcvflbZJDMJIlkqKnAPMpROlb
DvpO8jKp9Zf5mHbwRk4UZaE1rfNO/zgUUwIgQ8t8owiPIYV235pcGOGtwrBG8lM7
ephatvFfBTPmiEF/4Z9Q21YbdyYMYdAvOoq22GLrebbBshpnYFy+phcTm7gA81R/
WEoXVUpMXR2kW6s2siv0dsq4SjEN7QZqtjdkN/YJgXwKvsOa7WauiTt60dcK2saf
gvLP/OAdvLM0ve00L3VWWuBZG//cEeaVn7zcvXVPgub1ir+/YLt9y/Y/7OfacARt
4WYGadsLL1hqSXWyU7sRMCqB0/hOClxlZ2pGu3lYf7LiTgI8bmL2UOplVKeFd44l
QAVFB+5YrPKpJ9fBRTvNdjsKazJHdmQzlvjdR1y72nHnsYhDzzR8Goz1fUkFBDsG
UP4PzyseJIcxqp5wXvuxw9Q6q2+MPZvUNHmiQOwRZrau7SjpHyPeB0e/TLzJu3h1
91uoTQFMzX2lOZj8xvg+tXnK3k2yi4CAef4/lm3/3LbBue1y3d1IZU7gSoygL6fL
YA20GO9p9blsdlZxNAg6X7S+dlSg25l84o/ZEBM3oOHqZYOxQGULpFYiYACMOmDJ
qZiCus6kvyTfne76zs2R/PI2OIpmr1gK/++J5VgO/Dq4a6oXl7n3kqxaEDQND+cX
/nlqZcXPlryCvMFD59sg4LSzveYzg5ZcSobd1Ky61vyWi7LiT/M3ytscY2qUfbV9
/EKmaxBQMYZgLJWzLx/ZBBzfCnDWf+hBAn+nQbosu6f04aQTOaCE748XIS+QKc8e
nK4Z++RBHd8F9TV0lQP+OgKsDpV2jiOTgZeMB4C6GmsAVWqYi/Ud48Ic2sELHqgc
SClTF7dTAY8xM/WHh9oahZA8oOOTIi63iERFyd4y7BXKnXyovyk1zxDF5t4jhIjE
rvYscdHrYL1lmbCdiXlBKVxCso+5+waIIJJMmi4pCuiB9EbRo/JZpR4QDqxHBqfB
bygEXQUoeC+jFJAJ96NUzzqFebPAHjv+ZOKhm5fSNUYcWY0dUuXUnwvifeFOm5rG
z7jo2l22L0kxHiAPh+K49MkA94h3rdSDzCbBg5JThZqPieCodI5eYmOROcJ4y0rl
c+29XGkSrGVtgwSZUy8XuTLxGCBL6UzUrsCE4gx2jGK7l6UVZlmMBGDJRCMJ5xET
2qtaBWSqpfBqpYprsUifOdXwi0j3rhoT6mFiV8QeV/pyphWdEFS8W1u1zGEGiPB2
kTqPy+bLOJltBzDwZRTE18MQPHjodq/AYQ+uClLt+YmrcZUilQIyUuI9sywYd1CV
NjQoB2HbB/4YdeO1FYwNwzhqowuE6QIEHC7UrFmQIVOgHlPCuoGl58hRyJiDcPWh
5pDshmV9hwoVlhvSQ8+msM5NrqCqeAAUAB407HkCIfWJN97C6vZBta5x9lvRTW+Y
L8Abo0wLecrXOi/i2B1CnuDcSetnM/Yoa4muiSE45w+e+pqOjXsnr/VcPTRXQzmi
nOUWGcytBonh2MyRpHhUU6DSatgwLevUcp4oX311Zbqk0K1Xn9ERmLQDsrkk40fM
rQC2JCZSNA4ox3eKHSyUJ1REVaWBczAey4CdbDsOzk6TbhT2DVdXH5N6rdJ0AeZr
Rnjs5RYvMKqXTF5kUUGvy6Fv9IQ4ScOnSx9VXY2sgUyeP8VzIt5DHAto76ljwN7W
y7glxbxYy7Op/1O5w+c26mxgMenOV1jsP5hO7OkXTmsdXzap5opUWtO+YE2CiyJY
mcZGnden0uWpDWr7jU6qmkPx4or4OniHQFpxxtkqRCZaMfHevLvemPtKs8rxb98Q
FvpF/R+mnNWShi1hK3yeuZu47sVZht+rmRJLx4TjCcWgFKcXIwK1zx2CyH0jfJqD
UicHka+umSiQF0AA8C2ihTOqJ24ldt2Ujn+RVsHT945EWuXf71QphJwN5lrh545T
tJX5zPDkIwfb01WuK1kcEJ8sRfrcu4IHx/VuqqgvFSXEo1n7M58CTb98TxMo8oVW
cNfe5KeXFzN+jm9dqZj2eRR3t1IBEcR7bK8c02Mrkl76VJ9pl9Ov38pVgAEdRwtX
nxP8j/qmUAG+8C/przv9HlxP3xTEoeoUI3yUOCSjznpOf7dfB7YO6cJujPXUP1tc
kDmnVhF9s9V8EgtmkQTgIpiGjAz3DS3bBbaljmOBk/gHIh8hdg3ynNHDWqn7pDcR
bFEj4gVRIXl+LYuMb03vUK4NF79cXr1tM2AoCMJWp2O9yi2G83JWCCLQocgoHFBu
8G/X801H/r9YNT2WdxjqkWni3189djhAoThJjmOnPVk3Xwv61VC1MdzVGsYPsQIp
Kaq56JOmsFx+7iMxDppgQLAY3DxKTmuJtynkghzviBnQwZTKjADLgiTjykplNGos
eN5zA24Dl+vzrvoQLiKR9xDEs+l/p88Mqd8+EH2RtitwUotWEmCOp4JEmhYzPRQz
jsLPdzYaA9c693m5OgHJbMD52ulZcRyQceT6JU+veabifWc4FzEx6z2n1hPl/2w6
Uja7dIOg0pbBoBrOxAuYRM44Wo8C5dG15L0tzwUE5672MUe3qq+pjEmlkGPbk74L
iZOFVs5pUI3SvgUXxq32sPf9OY4OUtybyNUp7CugJcj4t66yfD/KFTw5xKLq9/qA
qgoX/n2J8+0Bvlq9Dkd9Gt4OfV2XMypOm54f/LCwie6EeNwtscXiZJ8tBxaPq6oU
2LgCCC8Z+yHTCHyQdtSQJYeOe2XEy27k7c5SEa37WKkPFt12ro4+N7zsagAkpEKZ
nHGWHmdDGPgEFZfMb7lyjXZOYTEfrj8k+K4cw7VklDIDcwT1Eu2YHk3n4HU0CVlV
E8lmJk8iEiS17d4hvzOzkmr7HBGh3roeGpI4DR8qatjz4ZK5senTLj1pFR1h9tLL
fJ/YKhpAJpBz7HKw5YkCKpAu39ImSmU/lG4IMRrWfUsGl3vhNl7K0PFP9d9COPcj
8jB3cRIST5IBHW6wKriPNkoHq5YdbW+FrINny022aeUvZsmdZWWO+idLQLO6hrnl
kbttc1A70V/iouk3w5QHIotFN+ymSoVKju75T5gQIF/ma3oNoZU+77/L9fgktLKB
pGc4dygQ6MwnIoJFU3cHScCEmJrOhtS/rZld/jcDXVQElnYALCtR2VaTe07Jr39N
og4c4WYf74EyPG0quXGsT6jWplfcasRZu7oNnbVmgS6XNZ+7gnN1Hg0R5Wg7Z4YF
aWWzb5Reieezt5IFdxyhsztr4Eft2ygLggfFwrLz4+yiEj6FY1uI9MYNdiZvoqDC
xF6bW8aFWbJpfiCBAoQmZyPG1Vm8qQmC7pA11W/lHAvl4hgHe+gCSEJirxvIV3V4
LXql3KDNHr4ygMA/5KxmjQboWgltJbf6xYu8snBQP5sQT9JmQsHRmmRvhEwCxQCG
mTqf4Q0t2EWCiZVLRUXRDm037nme14+osUzvkdG4/Bxm8SouQMCEfpSXGPNaoT2/
VLPkhi9qRzh/dpy7Uz1a3vZ/Ht+fFTcNdrueW5Ko8I4Deio6rEFoy+NzuvesGYhq
9cydkx2UTLKpG7Ey9t4N8JCW+pjUlVprOvc9NZpZEw9328kRqVDDIfLOsLNRx71+
owZ37OIxH8iv1VNE//EsiN6gDbkF5pHOemE53ifBu4yXi4l7K4FtpEaNUncxWFNJ
DwwB5fKeUHxgn6ADjC9TmcTKT1mm7kuguOPXsuKOzZl3jteh/j9YpJTF1EE2UYzh
jkvYG575vgETx4YfjMxZHBsCq0TqRICY/WgvAAOCKdNew2z7Lot5RsctB5l+gvJm
5dTH0xj6bNuz9fBdV56WLqOx17eI+JK/Wl5ov7hQjL8fcIkDNW0l5MPl/gIjhwkV
3qwEHc5eOqiF1D/Vc//Db1cPvUw2SEroGpvWHbtPMhOs0keRmdFMwyBgE4fzjoXU
oubxYOMWV5TfVUF5AOtes2ziqrpGJNz5TutGzANnhjZncaZuc6IOb8eIpHgtScFb
W3kjuOqUtrQ6cSVMtf5v2GvKO6l4NXOuOZ5Zv70462gOAezJLr+yTNwJYV0Cl9U8
YPTfVVogSIdhA2Y2Vv9Hp6MK56TanVvFJIHO5kA5f0tFrb5mJebuJcJq+Ynr3Bpr
ZQyCgzG3rU6vqjYxBN30Bogj14RnInK1OKFzfiymelwreFYZkyBsqlBoVD4hKAWj
g8PbFM05BauIICSKbyB08DNb84EGgNLaU16NLvKjkwD6221C1hvXBvUXaqYT9IAd
KUuUu3GJhG687MuBfZsqyhJxWTysQMbICB5qBkgAoWkDTP+cbJGAXSGljh/XnLGP
3PLDzwIijdvS5MNszhTt1cti2H5okBlj9DxLWou9mqKGu3/s4br3ZI8yDUD4wkUO
A3AVDcFx3HwW4GYxgu9lQu/jTPR43NKO2QFpciH4bPOZbHxVl4ndBCjxqA7QLANM
LHifxj1HcBkl93ZOkSAcqHOsah4bUlz2YdFzzPk7XasYJddRe+fXEHOlqjH1vvQ3
AzJcno4A8MXzf6FuRvGo/CYQhDbMgBJan0eWFff5wn9u0qVAhaPvErt98KoM5Erh
o25713KbX/xT/bctCy88/04WzUmmhIfFHiPft0yHMbClNleNJY3whHxZaMXZYY0i
shj7i+st4FGafszcROAwuG0MegoMZ0MrQSjFhSyD55wAUO/Jvp3Ma7dq8RnTaCe8
wft3ss8cl7mqaQNSW1oKHq45c8qDKt6sj9Th+Gul9C8bd/UnUYfrojdkZOB1Xdla
msR5rr3HU4zxrXs5L4rQkk8qVyNufo/X/0wBXaVlBofAXVmadz/AFwqp9WkP/vCv
lm4hJ1LoRLAjT/9bJwfdwQyqp74OWDWI4QHrbBSPeGc0n06ACuSI7bH8Hi0R1jdD
9iwajvdMo9IbpVY+MNmOmqRkFsd8t2ZbWs/Ik60qIJcx16AdwQFpEmwiSQgZYH0l
ihhD7JDyM2uUycmsqm1AtZpVdJJy8Zd24ZeUmYvF6JJ9Dapk8Pruygu9cUGKmyx1
TwNr+JYz3uv0EbyYTnuOTbeTxPHeECPiypm7zhLMsVT3U1d7nU8/uf8BvmQBPDea
v/rDJ0v/zd+5QMMHaJHqq3puL5VusJukVYSF/1UKipkSWpFBTyaYpgUKIGuhT8Ne
8YzB45tajq751NJemi75TAfp412WPWTd+FJpL/mZ5w6Jk4wNmO1sQKRfnNlAXOaY
MXoE3EMnHSfqYVNIt6nWi+EdNqzl4wG+sMftVPR6g/+U0jFx/dKl2OYZSxaB/fg3
th31Vkr/ZtoX6hPIXQ3rPb8ZwHgTA8QTPdbomteS+lxLbtyVAJ6tnLWFI4fdxiu0
cLyAxsC47NN7XuWRBYk3bcFD7HCoCto5WuniCWNuq9M71NeVaukEoYe7zp3weOA1
zjsGOSkwlzsfGDm+FKcBJUAqS19V3oRUBH5zLtRPpr6vv5R/P1ZgV5nI8qrp532Y
C3PonPoZLJXkIIhrXHuQ8HV4FRHw/QsVL6l7T5fzsQ3n+oMAZMBypkzR2hX/gh1F
7DjwzvOS88ZiFuMAKdWV5hO+LiYGQCy99Zp0fcW1DWHLHQeue34yBrnj8EsTAGmT
5NGDXalqN19D3H9xkZ/wUPiyxyfm9qtztm1tBlKyzC/ZY8u4UzIgR20/o6jjbC7U
1r6nMS7KkPSUnnEH4kkIs+5r1bpxuCXGg5LPR08CJ+f3hUSBy2Bc3CQTWQnMspJ2
A2P1RWw3NigzIVMbOW1X1xCYTzH0n3asXAOXN0hYMlIVRLuN++2pD/le9k3Mk3by
TTxN0HPcDp7Mze/TiBkPPekVtcQZp5bMp83RxhX/QYgrWF16MxDysSCnZmOc+t1f
FVKBv+mFX6kNA1TulJ/1Es/W8/dMzrNPjPilq57qehmz+AdphmbwgDfn6OKw5wk8
90ZQIFUJ9YG/cqc2YJ4f/47bwar7V7+MdiD41VF3RyvZ6BiXV+pJ87I322Nrt70K
BTDpRcNoIcX29pCpgq2DjcRNy/Zf6Owy6y6jRq8bPLZhoLPiyXlvur1BuMkwI7ar
y0DzsLbFRurljmozlI27QAhcWBOxv0LOd3mpYTvY7DdyQkwkACA8tJdZAXsVtDJ8
5CUJPhzegz8uJpfQjVshzLKohxYdVrf/ziUaLcli7POcjA4WE2FixDSy9ePg1xcI
kmqhA8G0i7w0QF2sTW5/xgxrAKYAuY5+4zItGJ9qDki1rnRHdUa/tzorkyZ2rIcJ
ReGH5Hfa81jDE0P/2J5DHt9gi0ciAKwhWDIU/IJkeJ3asSNK3xaa1VUf16DmBMHg
bGZFZxOHfCdjx/v1/D+9WIJtiyJZLLHT5Z3z97H3JtzcCEmd1/nZGPUHeqPGEO/Z
hv/VEs0yH4x5JMYWJj+0cJpNZE8WD/1g3PON3Zz/TYwQh5ypVmSoN3oy/ECBTk4L
RYCP/YZ3Q36WMyFEfDfX59oXsDVv/2ZEDlISHh+VcglSXfiXIj7wwVyNYm2tvkkX
aOuzq1jQMq0PyZ4ASNrK4vBbM9+YLefQ/H3JVgxtAuahkfQIQJPx5u8N5S0bRc5a
W8d5sxGEtWbnXKpBOKO6gtLaS97J05/8Xi8EwV8BMBDofnWpWEiChOEfg+FQ4l6O
6f7ptWIVTdV3e1IILQk2Fm7txNHQ5kElF+jZX+pXaXJjjlzrlhFUF59mdiSc3bMa
UJoKQnPfvQgWwszeL7jYQz5JqR7DB+X2cY7eK6ZyeEVfdsLTxsJEX0ZpW6SBWOVy
ucsXDbmfzbLZ//7CFQY1uvUnOdQXwB42G8VV9siqas7Z6QZqQREH1/Zbzhh4g7tl
vfuW0jt7wyazSWIf3cexRcdcuBrUF6Lrpke87aol7vU1ScHQTPFUjvxI5GctqFJo
VU1WZRR2qPT5URO/gIf5zQf5dIxoe97DveeAI+GxakOBUAgPcH7kPivxwystqqxU
58LIMOAX3dXm5zmxjlf24jNMI+1YwUuHNesgM6bLOTZirf9HXaUhGMZf/r3vcFKR
JMvME5dcB2T/i83gbSQtzSj5WhVIC8dzVOFN3VkkfJ7XJmmujp0Ivk/OpX3yNJJ7
olo7oAvJHojKHUBt5IaF3kEgl8LHS87L9SB4Xcnw8SyXylhnv0nme4rkxpyVLtHa
S/G7OkQ1LmtTH3kFnL8eFOXp8aw8YFJDV69dJntylj3Mw4/PpipupUuLPvM2dGQ4
LYbeZTbaZkZXkeTGLu+flR5dbvl0qfaC7MUvPViJ+CH2WtbJlF/8efmJ9UzETRbg
rXTkXSb04Gn6jC28fuEO1DULTUTGePoKWBxWZ0SNn0fFjFDFX3la8yr0WeulPpax
oPeLd9MkNWstWgBiGHZLZoORQRvmQTlEk6Pa5JZ9sfikpHlGoQSGaxaBhUGXdUtH
+E/uX0RHIxXPxx/Q3HsQohGy9lESRu3QWxyC3dzNgR6jQog0qYRClrY5zLKFGsDr
uTpH20BWRnE3aYoPncj01iplBQMApdSV7xkFPNRMfkznOC40B2mOniaHsQbtvNOk
zcPK8v9BnHATVqS9lY/G4u/Ehy329crad72g2OENX2D9P1/8JpuzLW+g62n85A3v
8GgWjKIQ0HuF1TjDpbXBNPNlACLPIpAnueGevzd/PElat2WHj0KL+t/84RRXhnnu
sitXrMkf2iIkt8LHJYZrTRN5M5fwOOgQWZsgrOngp5Y1huxpA/EYYbOa+qTo4na7
LzGMJkdJ25Nq041z+ooa+QSrBqCrDwcTcB83PSIKH5u5ouqdpWvkAfmkppy05oCO
LBC94C/o0EXZtuZGkgw95kJEvwzBoP/XC16LeeeYuRsXJD/a+d2wTyUjUTlRU64q
gNHM773F+HJ2E9SPWjs2Py8zbxLHvObjr1fIhYyeeDgXsnikw6Lm90ZxQOEFJEgy
Qc3loYoxEleWLhRQL+mN8Q3UuwjikEwEGroSts5Zi0rqrG9gJN/ISp2MoORXEmmA
KfAgEB46TeUtjzI3vZkSSfHgvennfuCAINGS0gDCtLb0yoczSPWsEM28vh0xVbRH
ddO6G7i76jOBAjrBgXQelReIg6/6zoqY5xJaOOvCDy9grOMC55p5vv5FuyJvpj3o
B11Pu+uizfjt0FTc0wCseNXEdKpqzF/kB6NOAjXWLpr9KNf+J9VUhL/wy+F5CIil
9JjuLOGSoED5ptNdlzMK37tg4pPNJPfY7clLyAh386YqyFGZAN5C5lyOJznkjNNs
1sX9ZIMF4tcjo9nEVA19nOlocHIRR3AMZsTKAKLvocp9iESunVRTgkl47VcZIvd2
2+1ohPVg44PuWkspYd5BbsWEyhdGJm+pLkwhr0qj3V0nWi4GpR3pwHtRyAW6s9Pq
Q9spPEtrMU5MMi4lKSpdMMqJtdtyGf6RaQE972Rm61czq5kASfQvVMBkAam9onaP
Up/BUsZV99cIR596QWvKDZjneMa45SlQ7jfvOvhJP9DP3Qd0eGRG4HEx4h6ATe7R
GHsrUVUHP/fOQdeVXvkvV8Ngje0+8sV5oYPofQ7j7qOKYpIzasLeZkp5nwd2hloH
G3W6XJMQ1IMcKtLZk+FVOHbr0Lx1f9iOzyPYOX7Jq9AQGCCHANOx0awf3K5JFt8R
QTqgYH4lvZFimOa05xbibz8uujLnT8a9ATDhwYnr1iRskZGpLQv9Ybj4fmieSsgd
rwtfSYh9Yj4tDecJaNC+6FkRyEdPiC6bI1S+R80t2uzE/SSETtccV3HOZf5LUpfL
KtAFghnlKeOzhfvrcJ4HXc2TOtjhnQvp8QPMiI8FLgWVA3JBdU4nLV+grGPupr4N
hl802KKv1jUSXVzTQ2BOcVL7lmf5TmBSThdEmBOn20rz+xkvVdiD8QpXtq+mle3a
rsFExi5/Tgej/YByBu1AGsUa/5XUW0hhd1uWOwiUTbPQ+d+zw8TQV0liwqd3sfjY
QcwyPGOQAo3ul7uADXUgn5xHQ6EBQ1kfV8TbpNnzVK4Z/oGxWIC1bXQtFqoOHIgm
3tcH/qbfjwExByGPGH7/f0pCDB0OelBHWKzJLOjDUPr9XUZP4+Nn12I4954k9frf
hBy6JO7nfoJhLz5NnYDTrPpCNR0tRi1WEg4Tu2aZa57W3cyQ4cZmZBUobOdcC8Ug
7tFXR4Ggc1/4+enYHNel9G4gtA1nFlBev+EX7rqshHPMr05HPpB7eJXixtaUOJg5
gsapky3b2zIMbZnJSl1XxT/s6oRparL5JrX6cSU6TfkrHU1Yno6OqGSJYca2u7lc
U7FVYac35MuG1Yb3j5YNxrUzv9cmWKOyvQ+F9Mkw6sFQOjJfvDu3Mrjq5qi7/ZKY
lARimIQqWmsmEwghaYJpIWWq1ieBDz+9z94u1qUt4Lg7xTnXuJB3IeSDBTHMeF8U
85l4+gTrSc50avmh0CEIT25MMuZw7BAVpWFDNdk7OVb/nLQSzQlRmiOEhkAgcSfW
yN3LUI16KQ3f5qu2H1U2RLOKy6eZ/+/VtPKv+tmgiFN+bT7694SrCSlnCjSPxHAA
r7LiwqdpoWvEjqgNVNYHbN7UypZjnXck2QZhqbxl5aD0k7g0Tq1xBvRhbSPGUDY1
vs54rWuNmsFkHFZJL+Vp2cPM1iFzRGsISfapTC/xJX6jl4fAx2U49vJe1CVSNImN
BrS9zmkpaQ2U7rwZuHcXLjotn0d8eiUa8vjftdJk5zhBSjvm96ckBmUDUP5JF7h/
Yl5Y8e3crJdB3S2VgWcQhYBt7/6mCQnbssJSMvrf8XS4i/3LbuEcLSpNZG5w4HmA
cWfCpR/mq9KCSvRVBrUkNmX0C3kjr00y0OPmUkQR3qntlVGjvDf+W8M4GwZRTiA3
PNZkbgYrmzjF7lwSabzj51HJM1RYYitl8Qf/EZWSRCvME41QpEJmG5Yhg2YThxgk
V1oSDAyPJ5DvbQChV++xrPWtTim55DTG00VtCDJNlB0F+H4t8cZr6/6IvvjOBUop
0XnlcqhN9yqa2oTvd0NTIOrBrtkABuhV17ux43sV7CF6wKRJ9phSaVTHJfofze1H
vkJjMFdZ8nH7r7bDBQRPxfEEfHh6VAe9gPHcOYlqtkx4RUq0UwA/9+//b2HrIfg5
ZyEk4VFeN0huQO5Y5LJqiiIkvnAA1AEodyOIfw0LKImJhfD7d5/OycA5fVyp6RNO
aIb/qBvrOs5JDrNsfwC5NpUJIGOhEUXwxD8Qgq+5seCJTne6JUoHsK3+p1RTXgMi
9x7AMsq6PNBm6azw8auItP7A3cW3+bcfzM0sFDNB2hNRCAxeHbXUak7NJTTgpz6l
PopXnMZSQEmv/Csyo4MrAVo4D1o6atLuptUxfz4LwMkk4CB2V69sokRAaNyzy9ar
E0qSKQI7cygQm0Cjzvrm/06X6n3dXMZVnG6vQNd/QVCEEu8v0DKuSslbRljS9vJ1
pR89Poxr83415lRCETokQVPtxs9zNaJi1jKX3ByugeEGgNtBerCfQR2VfYfdoVHu
odf9hfnRl1WjHX6WpiXsK/1Dv184LF/vWmzGqWwTEzyWXVlBRHwAn3tUKd53g/a0
2QI1Dbscx0vt5v7uEKFtag6CiVVXBQKoqcQeYEO5heJEsgV4a34e2hz4NIz4Vwi+
j2H6R6mvRsfpEup+b9oG7mCVQIZYWqk7K0cb8zYMBuKSlM7v3IGqs2A14HAm3eYJ
mcp2ieEuYcOwbeBgN5/EXAx4UqTFzpprqqx2ew+X0UZq/U+vTCDNrX7U5oByzkh2
LWAl/6c+LzHje24rlDjcHBDwqwSY1Rk0mIFDb8P7W2e+Nk2/itbCKK/q4gPmqGgk
nFPMvj9q93EQTEoUkLImBNAOYJ4fXx5hjN0d9OGzX3m4jkjhQPpXizu/x1vGlILQ
aZ5tyyldMQxh1xiB1T5f0B7szd9v1uR3/hENa9dE+BY7wo0SdpkwDysEbhV8Mgiu
5FJxs+vdi9wSDVhkcJ6IVWRkczwyFRj/RNF2Qcga7jX73dsJtqYPN26HCWiBYc47
uDLJFGNmQ6RPN0UN1/zmnVYJU6/qGvVIyGZstVrCukVzHb1aNbO53899d7FvYNmn
yh3HGeyBIfsBvSiTUP5v4T3EYEYrz7VUOnk3FqetrCib+eKwB13FOIKI8B1uOyUF
/wM2Fpe6Biev/SmaweklnsqShqeCjny5uvLeq71oER+wAm5Jcpan6F/vgn27cp76
wKuzyKitTuZyLW/Ce9VU4G4QUEF3/7YcYGu7XBUFvVR5SD7BBSJKmYKCepFZL2Sj
Tkg1mlDO0ZY5jBb5LoX4zQBbCouzP62KWpwFzIp8qeAR4YlSxoNUoXfO0sS1o+k8
xlks+PxPj5t2VVmrPjmB+mJDeeGyCYIKcOM/Mt/92t+OHfTBxZt3QlTGudWJun4T
OmJhBcOmhAcy9N0jJiPJnYhDCVzVW2FxNqroSNU7dAV/06yf7/2TaN7rFF8QNFZe
O79/Id6uznN96+aFQ5DowCOhr4OeOpa/ZddhhjKIirU5EmWg5p2cYpaNw8x0uOiC
/hI4Pv133Hvl2BIq0T73pMmyW2mhjDuNf9THiNQlUdXB2q17eJAV3BDJE/JQ+DaX
ifQYmmrf+FkjBkJecREQGdekTg98DRGiGvbEkR25zXqmu7Zj3p5c4zvafzLxMmfL
eUk7wNgjaEWx0cWTjdXZkP/elVza1vmroXRlF8NoZJ8PDwvp30lmHihU0gHc+1in
U9QUIf6UjybtzJ8wTnhqWYuXe6lZYyjx8j/J9+EwTZSVcCUP6WxfSHrKnSPT0/Za
GmsBJ4+PZIpvcNgRPCzCpw9KLmJxd/+ayhVdQAF4jRwUydZW5JPNvmkz3II2Vn4R
Cue2SkdR5OehW9VP2ZkpBDool9LYPhKDNkxkSKjWvdLVn8tOHkA0jFmmaSgltp4H
D9HkdPaI0YSaXl5rIu8ZSyOwVNSdpjRY/Rqn1Nnu6sQGbtMsvreDI7/M5dA5RRhJ
9aW7zZUjRQlZXGT6HiFX+KVt/qw9UyJILEduylz/pJN5a5F6gNEqfuZBwlKcuq6m
UvSYTd8NbPkMDDu5BvIlwpl8dRyUtN+5QqxXT5yQL6qj2drAbRzP10ls9+q45l+j
fPhQUMlvjD5oKwQ68gxMuPuiBn/uLC72bX/8K7LwQfqZYdQgU3gCdrG48rmh7VNo
z6eE10WZRgg/T806iX5GPsRd9IzPU45ZhSv7mC0ap4fSJ7ISSTwmtVHuzajv/PZI
R4bekVmD0Oj9CtHN25hPLNxIFBCdGCBgNdx78mEzxNJp17bME/TMiEwWN4OFE8Ww
du0G+QqGGFX0hv8u6giO7cF5URLc/w7ecPG/+dfKDynTwf2LFDMtBOYhIh7d1WMo
z/4pErF9zCsWrOB2OAapSRPs1Uw/igo/E5Pq0HvufNtFAquaaNdNz4mnldex8/rC
1zq4S1FO5PLcLmUzSOb5gAQr+j5LZH9w0s5mj9S6dV/ohf1qn7n1WOZ9HlBK3QCg
3BVOR32CClm2T+CrSO7L55whtgHzYnKXa3FPc9PwLI3YDgHufc3rf9wPFB6ucox0
1E9iUIkto76iL8jPDPYPG0sN6sY8XNAN5nMLahDSlYO8ScjAb3sJJgES+x+f2wPB
0qnoR5/YDbcJGJ6a0yMTgbIHVl1hH6DSkGA3sy/rZBvxCxyrZroYyMyt/jycPfj7
XKi5jNTYnhzWXZZW+U5/e/Y0U5jEeGBbCHD9R3gjdju/Lz9XB/jDnFJZGh6AOMIH
wiV0zNX/2M40JWzRYLgLOI1YG0UeP66/qfiS26or5VZi0EQyiSuQduRsn9Ji/9g2
Zx94rFEgg3kQEt25EuifcBD2y2WP97jpIGTJXpVNhKswEwb/aAXev5My7XfgS3DR
D8A+/uxnodrpyGyxEEssh4Z6K8H1rvOXNu4udW7AxnWrlEujsDUHOazgJChH1YwP
cpeRuQLGmCCPj5xcKJrEDaRiYWgQfYgHhCzM+jbecz3AjRnhsEwms91Xl9+Cc4kd
dGdNg3gT+OxsUPzHKyBfze7c4is69rBTfFNoXoagFoXEASh5i1qhaA7RAyzaStMV
7fJszMcqWcRUpvqFltMrUmDwHFfskyirC2RjS966dGkSlOMsLZhR3qeQHOKb09yj
id9fJAA6RcfWXgHAIethMcYnecqlbDA44l2BAiWW8r3x9Kywly2JV38quVHUfV3+
0O9MwR7cjNxvJ3nQyZLhuEV0WiHhCDyTO/y4uHO+oeJKvn92MIGAkr2HX2Xjy0T2
oklOjmLpiIxQBnWUAsGhHeoETG+McGxYkPojHZyhkqNOtSQag9X4Q7F90MsiLTup
uBh4lR6X3Yn8mR+KJIcVt1m8OivnLgieEmlvu0aMvz/DNI5bCJbOOMuz3x8XZI/6
9uYvgxt0yaDKBGLuPoQtS/CzCUd7NrDvd77bdFuCiYwBgrn2E16JhxXIXHwwHE1s
LzHJo0coK6ORbD8ANQfIaiwofWgE3fUaTEVwnZe5o5d7a5NdVck1e/Q+QerbaJrf
o7ASGLcWElVKl7ZJZGcJo1b1xFz+lSBktCHYqCFEXAqtxLNPseqoiB9BCLK27/Sm
HJNrmweRiBaX67KehM5AfJbvYyGqZmzK66S31FHOyLT6pu9gozL6vaGV96a7VdR8
0m7TqSPL95tpGMFkBg7hnXXKQyiwTNgJeXpxI26wUxDBysgAnzWEhBZtl2wCb3he
QAu27MCsX9rMTvxazJI+HTHVltjQeh4pEkXHlW6fubl5dayDo/eypq22RdodAxDL
yL0a+k3s8UPrY8a+u7NHa03p+r4PFRc5GEr0Frfa4xhQhiyc3RLF9QBcBWmxxp1z
Yiy7W4l0SXgsEQF+Qaf/NU5w3SVzGoA6uqSLzKxQH967DtWIn5BaQ596Q1x0S8/3
TIl1qBXkp5+j12QiJ5aftYNlinPaPiuMUn6v9gII+N4UxWs/hqMQF5OeFDWPDj4X
aJUGxYMEjZlXmyp7nVTq82/1OyOBVQ06V1B1crR8QFgsEpuj8x2pX0JPYNpwaSCn
Lu3JmPc09g2dsPlhWtVijaBgs3E6DgbnKUVcioRSarE6wSBwhcuQ3erzeOuKZatx
iOWetlSHjGlhilfdasVmydUZO0gmASsiPXEcQGoc7ED4irVMNeGV3UPJNuHpMrgG
+oF9kDu4OBIvOYy2pv8va7Lf4QjxeUjx+TJz+OiO3/nyb/fZlrDo+cYm2JIkMxAR
6cm9a6XIsJrL6jDOMIh8tdVFvd2kiySY2fRZ4hTCM90mLulfAtKQlctuNtKz1aj1
dRQirIFfEuxvqy8dwfemLvCNgPncBDYJ+/fDLft/aziNSvtoOVhR2iox5ONn5gK6
4xvO0DNdOYUvtmBZ3ZMN7ISEslUKqAzA98W6dy1vJ+epHqIpojiL+AyDyu1su0nP
z11W8mJrq/iey7q5zvWg0/R5u7j7ZdL+CVLHZypmz/UaGRYhEXqggv3MyFb4foeS
RKY7Gio3LJDcRkfPnCLvRytLuQNYUe5MKfJuLzBh673/4UsfO/rre5rs7dXMM353
jfLrP7Kjm1ckqEbT3Dk5eGHjcFdpdUB3EkEmvO1TL/kgum5PtI1hp2mMWtgXNs66
rWdBtAlI3VR42+AWLZQgkGiqKHn/JXmpiFiWP4qJwYjuS3ZogCqBJAgqCWo3s+Z8
TlLhKlRj+JIAa4ALkYMsNN318cnTtpvk4K0foeiaUCH8SOCJPJ0VvNnJh6gWcTID
AUdu5HEjRA1LLr8Deas7tPJpzDrWKygJd/DOHTs29WS3S/b/Ije+eFfWNF7+gFQn
uNgVuwF345dl7f52BwVIs3hI4Qke37m2LuQhnJtN0itzr5PzADbNmuu4L1+kAxcS
twEJZjNh23glYPiRuJ6PZ5OsViLhwySIOeyby7rcH+4CljsSqZguM3GnQuxJwvFP
Y1ybSkkWZf4Z16iTX857ZhT8SiA+kKuHzmHs+l/W+auPR3l6Z2QYgESi7EzPtJp1
IIalfWTxXKd69BZMctsqG+Wsvom/5vQr2UDbUFncX15wPV+VZmeBg2oNVoPEpRM0
1CZd780CgrMlpw9g1tC/7pZA9bwWBPmCyF/vZPTmh+0ppeL9yjIGwDfpeZ08O8oD
DfATnx6vjYhPudVwQa1wTRMQ+GrNl8bxYGHyMISN5d7I5kDTJWZkrQ0NMVJIw9K5
jijxp9Y4FXACiPa/nmEFv18kxEmCF/VnZ/Y221jNWNyrx9tDBGl+k4JZdJXGVkJB
TkdfAZyxQf5XZs1tsXLSAqCX1q0bGt91JDj2kbX09+MENE02nO64b9CJoxbO9fYZ
izmFUtIFct7clY5cg/mBKL0HJ8omxkZmuDRMLMEFn64XPMGdScHHbEtjL9zBg/P8
VJOLNXbmOF8hGwt1/ZtGY2UvD7xbFpCHy3hcwiLkrXBc7sAWg+5KEAjxVP5jS6iT
GsRq9z/WmkIYOngHs5WU0qrLM7Op+V50HtXtjBoCoCZnyatqG1dB4CU4PFwTHsRN
rZDfxxu8fxwU1/U4z2geKx27nL7N0cndrKihoq49NSxcpAv9zVzdhA6fOmXHIhpD
oMDgxzP52oTpb8zrn2FI9i7ybnjrNksAeOd3a6dU+FTYN3/FWF9LYwRq67VqTKnH
hbudn9BEZjtUnVOYCK3u++fw8zQaD6lhFtDmt27FMOBrB7rJbz0frhskgLXXUJwe
9GDUKmtUuVPJ2rlt+CJLFt8QBcQMWgetC8Oq/9mBdFcJWlVv3sNeGxIvkWGLUybO
e2oybEqMdYxwy3TKqB+xR9iqumFFO1/toDdzkmoeYg5Rif7iL57Aon9WOWRYxcLD
DH1NCKZwrcCkPnExS/2U97+lFh0h2/jgF5pKGIoSuK+GFLhNuzT5nxrTsdBpLCvJ
1T33pv2+iS4pFKm5tUByzwjg8ZV521ay20hVn9rmDL/QNRKARSSNQR3f2KyKldfR
4Srb49Y32G1yHHmtV7etAc6ivNVH45UkV7uwBSB5+qHCjHsw8CKKizNp1vhRLqI7
9sSqiBEcMWYIinO36jnkaGsRMwlzlb4wH45mLGrPmzkS5f2WecjwFqN3oBAYTi9A
Vp/SjFrE19MhNx6gTj5Hiqag23v8uRG4/g6mR8AaMh7tVUt9ZJrsr9krKpqmOX1L
/DfG9SWcb54Vm/Bxus+0qBgwZNOBhgG+e925IwewuQtCzQnJqQbmC9HkxIXe+Lor
+eCerb6HIrjYYiLAs3gXMGi6KQXxYjLmKklFX3zWGkcp1RvTHDpZC6qz7Vxg2She
cuckPC612dLRrNoZyHqUmDodNCJA+ISFa1MRsG83n2YEy/3r/mN0cHb4MDqCGSpe
Z/p3TohqyWnptNfpsxFzGC6+ZG9i9MZPsFnZpI0gBYhn5Sgr5HLdYnf97+WfGlgh
iD5aIBzQ9iThLaURiMuabrM6zOIGx2NrmM/wKO/JvQhAMeEYViX7dJ+qsv5qgujJ
xLmh86ReADYNpIIDMIcROTfxKhRoUe0FRiVRnYanI+7mtQ4PqXoUDvDYQV9BbMe8
B7Oj7jrhij3AizlX6rTZSaWsEHQQpqRbxQJeG4HmeHxpGNOvA/0/Nh0JoSXrNzyl
E5k6saGbZO1NBJIWVR7atq0dxkLuixOvD7Zv6CnpgdubPwjN6koLL9Ofl1ifdImJ
L7q70O57fURn8ycLYi9xngNR4zl0oHMO+nBnY30NGzvo3r3+kQsGUNP0BLt/o7dI
MhLwn+4F9UxbeHrJC8Z8q2tQ/Uky0cwlKZ+iXjEMKNmkybeSiPkjTs7erz7MxiCH
jnEpiL4ErqWUaNTRTy2uEMrCEAaShaKXEq3cVP4JULFxzxALH1YPTVA9u4/UfOKn
i90lIs7/B55H7gyVWQnjRl93svjGNGq1YqAKM9l1xlNQ/S0lJtTcygshW6y1aM4Q
x9sYov93ZsJYJNwmNo4HBaWH/fMpItdFW49gFUEF+SyQ9iVjPvhEM133pxcJARHh
6N4Ks0dccz2iF5Z7nmxxbWGWpsyqmCPsFj7oiGd1u8JI+ThHAAoyn4ijr4jDHNp+
qJS3ZWfgNv6soooDxghU4YX0a2aVzclzC3QkJBhYCOm/cu+LFyO4kO30qSD8f1bM
+quMxeyrejUCiFkx2xXCbkO5ECnHevtzP7mGcFaKDKu9Rzoq2B+OrDL0gLjCWtcy
DoSVINbcpX69liGXT5F+NDVlI8I8Ouk/gKhqw0jff8IHu1iBw3s4Mx+oJ/bpDnvq
4cBbVaS7eU6RMbQqE3YivoBC3yk92kh5lnH64l6tFwXiPDW1ISbUR1uyFqApRnm8
jDSF44vcpnT5lHgdCQFByZGgC3Zx8/Rv3kZE2B9m7k3b9q/SlpJN2IzZ/oKtk7HG
R4/pkYzzIg+rcvJ7zSp1Q7CkrN2Oz4VjnbEH7CLi+7HR48CTVM/WMbpR0+AjQwsj
fYLF8WldoTHpOhITULLqQxf3gJGbCPi0WFAqw63k7XgbZX5INMOsIvRKiiZhriBl
Kvv+HsSeAkuCQjKZS8i1TcLHOsBhG0aJ69lfEA1eH9ELGfs0rSP05NES40mcGIWm
RkOBB0OgpWrdqK0DL+cRRbRs9HZQwmUN45p0Wpw8TM1rhwa7HH5TbT2IHgglIc+O
8LPCPYu+MEJSfJFPOfIbU1KVgH5OcLEoDtsrqMxq2YHqmMvAOvUAeRBbHpj+KKTh
FX8gS0rLxBmQoz1yjkQ8I6pdXaQp70F92w5rYSVAhyVzZwvBXnpU56dD2ENLQPUG
pbSG2L3wd6UUaL63WqlEMIk1gfb+8Fs2nnS+Uz5EaycPktM86SydnCYUaEwW2Gl+
3HgYmIedpgtoypMZrF39o+p7ERslfH8YtcnGyK7lJ5PiM934tqCm5MUz3l2y/5Fl
foKzkgEYx+NJJOSyF+m0H4wICCW7txjAn13MBThrNwDtYDXf2TitM7i6QGBFbIF5
Iqv//8vAOq0yC572rthPnL/PYyB3UDV0C17exAmR6LJcEgXimqQ6xh1EYX2m2T7c
3mkpO4P6lCR0QcWWhxoqhRkWnUVPtm0tD4HUOU+dz92XM+ww//ZuClw0h+llCzLW
F+pD/5lLUCdoNmAUvz4mi4qhEWHmuOaO4Z/gFq2X0S0c8DjBhWzSTtQ0ByPwvTzU
4khEdbBUQiPcYx2QNwVLH0lg5f3XUxMeXc1ZufDAq9SccYVds0BS6b8VadoGO8Dj
9SmxmOMXcjIFoOH+3kQak/mD9iFjcixWOs72NBX7XPBBRiePH62TVJlrmQn/wKCZ
wk/7FnVqOy/1LBezp+bEqSdQMYKgsoHq3dGrHJ8UZy7BbPvCTjIZ40DnkGwYY24L
BAJvxEusa9geuAKJf1VlxxdHLhnRpgqlP8xbWYNZfleb0AxqWBYSccC8UhWaR2TQ
H6qzo9xUvIoDOxxuO+d4rRdDdWl2uu4A7ioJmH90e6FTDmocN8EHou5rK6Pk6qwZ
RkLVjr0JPOUWySGPkloJtDnehdtUSfaTnsvSpkSRYTTmoQSzonhEtXMKGdy3O6h3
f3RwOfD40vTaHR+aTDEbD6p+ct5d04brh4v+KGYoB3CC6gL86PYHNubeFBgqXbjq
OznTPqoQNLhrcQQ1mQAHfhgkr+uupB5/29ALRJ6FfMsJknRH6sU3dh7jTtCrtO7X
Bc46HKZ0L1SonFegarHOswi2Bnt8RSdiDOFeyySsYiQIpN6EbqKMIFNCmEO1CRny
bTnOiTfo/kEOzL9dQzzGdqxcW+0lsL85hIFcd8dfG2Kw2ZM3wwV3kMGNUW8IimMY
VH2bKPDF76XS1xro0YADB+9xprNw+ZHLhVouynPbZn0eSHUnomCcB3bVECSxrpvt
cKouuvDbXEfeoJAm9QudD+Gv65pmJ3zWxzJ/5HS+1cjp/f4mKUqVqU7Wp1hHZAPw
Gf4++aSgHLo4Ynnvr0rJuE1U0YXQpJXhgqUABoI7QlFYB035fkYYrHxG98b0qxc+
MUVikNaNvGgxVO0j+hgJ69MGK9Wy3vo7uvssTXz3zPaMmRuPHJexL5sYBZOTsJAW
AbrGZ5E0HzhB4eysBxRML5RCnAoTRZjOAWlmKtAT6MoDjyqeO1Zi7Mz/QtxE84mG
jPpJ5+V+9/Yo89YujcxJyZFexAXbE9HEDuyj11nwiZLVZ8HPTUNwk+0gz7wiXp08
7+56FlNAJXLyMF9jHHj172NOmNmS7UIr0eN3AswJ9/ty2nrlcrszgLD/bFkug9dx
olpdD7OdiILdv/NOH8d1bPSwI7QI4IU9IEVtWUUZe81fDtlaH/L2E18XRWrzsy60
iIU5G/2Y1NrGNVuZCQPojrUnQC3Ka7eG/c3IwaroQHKaCv3fiY8go2UH6Mk5qK0o
Mau2aGJwcINbmJA5eo4wKKmbulANp9cOZOcgKiMhG1RrhAUztAqqQnkxCH522E7Q
BDlYzrJtQWIIWK7K/QqAnc3OS+BCUXQ1M+MSvN8R/GGFN2XX1FLmRmQNF8yvmRBu
fJ0zXb7uCkWJ2ch4kUECaTs66wM1VFeFcw571pbrwHF020jjBd+hJhFfFeNahBL7
7/lslK+8ShKCub1jnk4BvRME7s5dR2A+HqINUy467N4ashJ5Sd2TmIUHoxqg2K6U
CaWYpOiJHtYYIvxRi5ICF1dgO6l2zSqloDLmQhvVe0bPrny1yEGWwAz+AU6K1BE3
El5O3b40ohWiMu4VOhJCdEu0a2DBeke4NDoljPQR6FjeikRVUWnfde+QPjNgjDIS
b1SnUnzDof+0InaaPYoP6LeZWHEiCOEN3rdXHGzPMo/3oOOdEe0cxrGzyWX1G7NR
/ZHd46YHjr6AfEGfsyR+nRiZLiU2M9Z6X5HD+QP71fwhetJIs6f5L1Of3Ux/MNx5
ABWSvEvM/gVeSXqwBuS0HhIYdU+dXb54aPGdQrxu454QVbzhR2NpQ5aqV3K7olrj
G/lzXD5GjuuL55BlcvcEJJHBdYEGaLVoxpppUVZUGu5tGyBIYkkc7nvejxNNJTYb
wp5Eag6V/ERIwG8TwOAznKNP9NGqAsw3LA+WI3Td0iKQbnIJL7YcxdOcqhtFMwuQ
LeWjJv5P7kd0Xv1AK/qKxXRX8fiWAjlGtzL7/pHITJv3hV0gzLNX78UaKuV+wqLT
p8BqI+ofWa6vhHhyesEcxlClT+h3nrpx9kit90ABPV5LKHbSPWFRSzEUH3EjoIDc
ABE9Hj08tj2cjKUQGYfksOZxTHZDZyoNscnX3leu/fHRORyaBKL8e5ytQL9gua+M
J+Y7Cb4fyyBDnfGNlKOgvBwT6cqlz0P4PumHKHJGccRQfpLBlfOuCJ7qu37Cy3dW
fvR9cEVZXd6URGB7PDZPJ/k3FZjgFQIin5BtYHG8H8rRwrEKSPg2rNpp2OdR7pwZ
ANcq3Wg3/mDun5sIzT9+nv4gwzV0iPbfUjGuX1ZwTdT9EiS0cpQPnsMg+NGuvRTw
z+fxFbTMqw/Le2GRyrtplo0jstoIcfbc3abobRC1WyBfW8raFnIUB99cfzipbPgE
AjqumT5Hq54kzFHD2W6VYjNQUtCNiSvGbZD+84OYSAzS4aCjwvIDVOm9iHJ3uQWi
dVqW0xAL/tHLBEbm4epHcFW+YaMqq/2HJbrSTvOHiL1aiaKnu7iszw7OeHV8nlbi
niL8+im0uEer292LMsVdxak29Hpbegjs3q94sCDnhaT3ATAN87VrrUiKNYAIDfo9
U3lRAgbgaH45yCESvyvmKir8pqURcN6RUJto1HNIm2gZKHbmhkdbm9LcsaZTkMke
jwuarYmdUiIH7mZUOTJ3r42KMWdxhqOoPGODblHBfHwpancG4bH5lCDHZ+fKpECY
V/61a/9XTZ5TGA+H+tEMI4+wCaVsDKw/2nt2Ld/zsnUxWF+0sYq/NYCY5TSCZBgC
IQ9EYlOZ9wqYovvCAxUPxQyW0bIGd/PuRTxs4ETWilGYdGGVBxKs31eyTan5omak
SqrZ5NcUAMC6CVimNtW8g7pkgC4HBoelQb9SHEzOmyWrAkdWSFnU6DS1cKQVZ+ri
+MQ9looef/rGgy1qNyQ/gBE4UW0nuGCAh68Xj6m6LVt+Lpke31ANjYJhO3HZaFu2
3yZ61v8nxrDaftDvdUE4mGlrhCFlylXdTmgadCBGCCTG46kp77O8bhhfmskaT0Pk
9xfeJqHTv2ZTgiMVawYrJu75K+zcxDZVDpdZzvCW99jAM2brTOaprcuJCQXsIUnx
H7nwyW6qHLYIefNGMdGob6JmlUFkaQxo8JYny7jiFBCtMZOX4OEsJw9ybFVz/tAo
v9r4lMpK33u3uNwquDgYcV2c9pTXyXR4i/Tl/BeMavOyIl8rmwEb6GCpxQhIdnmR
TYKl17j6clDb7g3L7oTYdT1NzN27I3z8g5+Yc3Y47NnkCPbJEeHj//jWTGI9SLiw
hntj6mo79nAlGr26SHwbOY3pUkTiKOw2Tclf83TEUPAyGa4exMyMnedZNXL7muUs
vi1rCmORhHtoungoeQ9EWsKj3v6/5sbgRRayd4UW6OEw0SwStCX532+bNspa0s4j
Qe7yONwylJy7PlZx/NLXX4kwI99IWk69SAMb0XnliyjIAPPjMHCA25GKdseos/nO
OYWAHyTS3LcidF8rSQnnATvHmXF71BdQYoq1KKai5myO25qs37Qxr1focZATP5g1
f37HV/5S9QWt+9Qx7ItAppyRzHsN2sPCB/tcEh2yysDp9rmwcV9Z4Bu+9YoHIozM
ZO9h4gHOhpbzoaJpqNy9LGfl04W0iqEsYgkZH/og+IpaxhIU8txa2GQW4R5HZdE+
bjortedAosKGTnkuAnXIt+EEvaTgdyk4MtVZv4A97mYYkFMe8pabnD+uYy2IM+G6
sco2Cg8FXkgy1b3T7HuZdvVi4j3+062KFjXNHLhmX6T85XyQH2AAyWiPInnLoSSG
exmNqPzLUI5wC5vpT0OkY2UxaHK+5ki5ksXGR+qUFFXmrxl0CaXqFdnMFUh4zN8w
RgiDKnm1pqPV2JH+CUI/+Qo0FwWeCtJg6+jP00ZyK7zn9BkuaOfwbK9nrsR3ep+d
3Y7YbcE5/DHEI//U5h0rUUWkOJUPJ1W7Dn6gW1CrJfpIindAZCvq+riQ3DU691Ca
z35f9UQIpJ9T6XLNtc+LK9VDRF3+G7j01vFmSCMMGYik4Qnkp3Ua0xwBkSp76kQW
cDP8VC5oBy9ZrdhRHdpzaJsKnwXB3QtxhJ6NaIpX/oM2Ij1rSPiCoCYSwxcKYSVS
3LZyFXd2GDYPYXJJd7/tvZjFuXHjovGrqXcDcT5S5zTa5/DXwEGpEyL6jGU3cqYf
NVsob15nfBn76Fxwrdk3YLEIjOuno58pvTuGcd8Cmy3agvHQAACUEMFooNk9VjVO
bhUr1c3RcARIqLaf7HWayZXwrioV7qh2kSvWxHDZ0tEjjLwK5Phn+NazwsmvsCVJ
eHkFiNaXC4Hpz7UATcN4Id2S7pZcNsVAjz9Px2HYzHgFjCUunKsaFZLG59FcBvNk
8Xre+OxfWwhKpWDC4q24sxp3bxJo5E1/CWc3U44SaQR19K2nqxEUj65i42fikUbp
eaZqXPDu3M487UOwi5Lolswd+tfHbuYBclRLqTkooeHf3CHPWcKvzdkooUxPmIZo
VajFKFurSymZxJeOHBokedOliWJU9PNXMDVxETPBmuoWc1r3oYEgzkPJ5eQQGXIU
FjZB02AXxt/QidiWOFcj0R0K1NPlG7Ivt+mGyWaOZPP58faQpt5OSUpNUi1s6U05
za7/K5JraB1adJ28GfyEeHMKdPU7CUkZOnyBOP6eIQqDAwN8FQGVXdvEYgTuxNoE
UUI9U74g0WnIt8YCGjD4M6lviWuGXP5ndtSGI78IAmuQomBM0edNBzJjkyFf4T7o
qfWGNP6to35Djt0De8d44943dliTv/MHymuahyfF0Hut4Ou8fjrOgsWkaeiVQPJB
xxT0mleglt2iIfFxtqeB7Hhtq5bi7HIDVWCV1WSBRR9dw8GjwIN58d14FdnWLQUS
v8Tntetdu99SM38e6e8k3i2z07qFQ7mDQYSBABcCoaYYajysNcU0aaivxjTVblKV
IjY5r+flr/xsjyfg3oFE7+49PE84l7gDyIULb0ToeTG+dT9+d6aBI09FBB+rAcfQ
vP3URMMQNYnqjCeKICZUX0rMjNCsXafichuidYXuE5dcvsXW94YG2cPjtCTL0mPm
Lw8XUST50vMOHVptCsJim9bXYEx3guaWWc5ETNw47DOvNLw/ylEm1/giVKDhaXAA
Meij+1e1BaWEdyWyIhABQQHCHp8vysFLhrazHdBMkxqZj9x41ury5YobBdNoTZXC
kQV2q1ZDwTn6f80EG8+jK81M3d8CN6ePdr+3uauPpGo8cNK4YNzLmzY7lXOdaXwa
AKHeAZSHyFapRiq+Oaay/ObZ7PGLvXQLaHeCijsdl4MG8Yzt62FX42VDH5V/Mso/
UAMszImsAAdd0pHSpJ7fcpxWwKBkHR/xNajl4rUaoBmPbB04jiHEOnSkt2Hzq/Nu
s3y8Im5hI6igIe9P4E/m+yU36OV/zVCjBZ+SxTAqIEorhdJckHthaToWBsTEnZLi
GL/vRwRSUb3ZXaUSQkmdSjYFfj1bK6p1P2xwB2lsNTzPskwz30Yq65D+8OMI/rBO
9D8/UTNtBfp/Ucp+NwYcgThc9XKE4Ck2ftOIhzrbbwv49jlzNKrJ7aed7S0aQqar
FyBMUG4BO23sFUrmondhZkkCg+TmdbszQCxBRGuYefSFR9pw/NGdmCXnJueOVzUw
0wp8g/fTN9hTOlt+AIX8TlWF3I7IQIBpcAke8J5djNWQ5UAbBENorI4Oem3FToKa
/j3aacXAMm1Hf8JkVdRakfkHNQx59C6hGlsFNwiyV3lE/Ufsp1YycwmIOlqPN8N1
In+ECE1zFXam29qu5reG8A0JFGs6GEh9U1P6l3Cu9bqzSFWSmXgEbXsPgSh6D5tf
En3356w7qiXmUJ4eC+/wPm5RnfE1xekZ7hvW74eqsLFLZUbrvvIF0aB97VB6R0eF
vBsokb/5p2P5NWKGf+EoI5CJJbd43+zTuVke0V4iiS67H+FoxPzIL51NGDFSXci7
sWvt0mhyOyA0mWXdKU8Ikag80il8ONt8bYhOmKG4WalA0OzFFsXXfhiDkoJhFrEV
TpSsBBiX9BbDec9Ua4IsP6Rv8+LYWYb0ycbe74ptLhmmlL45I5txL4npBPzMF5iW
ESCiTif5GUt0eiXx9luJPbJSd9XV02j97jK0vrMwtq2w4P+ZPbaGfj/7Vy9Sm32Z
7VwLPUIOjOQ4yWTShW6aryt+g6y86LEIcz3NJmh42OHHJo3TapksLRhApl/Q7uWo
gZ9VmiR1XYuSyzHfla0fzqCdgHHTzeHq6vm77Y0hRLBG5XUZaV7kd3bVwjhT6S+P
MCb0w9dAX3n5Z1hLGECotjGH4cFiQ7nkaYxlhYSNfwBvV0l0jpGfXt4thxEhej6V
0sYyRtiW8v1m0H+mIZ9JCA+auO930YZPQlIRHnz4wAAwA0RLm6TkDEtWKKyC1zU8
PmhnsEF2ezuoXchxRUKYOt4z6/IsPW9P7j21NcUgVzgF92ECDRZUuXMPYUzaT66h
n1gjh8GuksNtDx9xtwqwJzZtj8O3CviElLGxJUUVHpUetR2oYMXZz3r1/dqoC/mp
Vr4hhoS81p3V5xdk/PoIe/XoSF6gbIoAvLpNF7fjZ3nU9Zzjbmi3KTUsNPbOzZYE
NxqcHvVO4Qn6m/pE6CH51anf9EPOQZmUREl/NmTz/Z6Ax4m3YgaHpQoRxBKy1C9S
knJiC4ZcVHAuOqmwayfvJLN+HUW7NFk/evtltvCmC26jlVi7tSRzOeBt6Y7kvpzv
+5ySflwc5m+Y7Kb14nk9nw58kuRTf9cc9ndqjha5iAH/ser9p6wdIQLHuzDK3+Ik
ifHvWC7MCvP2OXxOzDtLMD73uSEZcrxfHXjmA0RJ3qfl3hQyk+CiBiFYCpUV0wC7
sYXfkK+dKjtuMRSP8kACRltDQULK93GRGfcBPulZjOyFoOSeU2OfODWQgKMGAj0F
eCRRgrSuwEqefRiSNInZ/Y2fW9OBPkQvhSe1o14grc2K60uiCmaOohiXO9myW7yl
DORagj2wPqTuQxOd28so82Kae9rvtV4vF/My1oDUQjpM4T0azGiMlluGirwdiiJl
19HHSFePYM9MXtpjPzyAnV8vkbyMtvXyfmVE6znbYaFRi7qBajFo84F6g9Bcf4bx
U1WhoF/XbR+DNrBk8IimjygH30giCp8hfywcC0vApQNHIzHovjZN7oqghPjjj4YO
u7V7B875QAYrIax0ywSmoJNk1svQ6yHoa7yzQsXYwh+AzQqPOZK5QMW4009krs+p
LEOkEUKMj8S680LN03pA4rFqjlH3M1Nd6aECC/Iz9NAEVCxLvtGlq724aODA2LNe
tr1W9H63UqUWVzvtYYF1fc3qZ084Co2/N+om3/WVH3iIF4Kbxp7UA5mxGmaFhtJl
jYW8S135caF3LucZf3uP+bNdm1dg5N9+qnf2UsmkaOR9MylMVlPmgd7CQTnogoEF
Y7PvYVW2eqNm0uBToLG3RPKPNgCp+tTj5xyhx1Iyg11MqUWbXpd4KEBjDkUxAPJd
bYAzHqkAghJYouOZh+M+dpo5hMewpc6I7gYN5dJiWVelGcNFUkCJn/M210SWEVNu
hiXERjtOsu6NN86MSyHc+8IotoLlqqwWEnWv8RPCsHkharuMj/UbrCwAUBIN3Sf6
g1ftTFp10QB7TCRUfeU8W1nrqP4NMHPoYYdO/qYsTbWipXeYEQHSgirryNKVo7j6
c+FPamR8/4rFXp4Zk0kRCo8S4ZZ6wZXrV9xu4y8e85qp1tXpCLgZQt6agkCPUJ7T
tcSebggRQvEQSg5rdBphusl0LsOx44ve/rZw1V9rt7S7VKZcCySBCf2kgTiLbefx
9OpkodrcKMfQu6wf0EAGzMo+kMcp2M7HOHNwuwx8FBSd9gsbhNPNryqW2SJP48Uk
e3gwv5A9SJ/0f/yzIVxgJHDEUjUP0S8QaYOQsEC2Ga2ru8nJSTNePr4s1ln8hkoS
gMtPG4aqTYFu3RBgGB1Xg8EOl2ofMgnCCdvfxFa9fCDCUFxJ8F9ik+g31oYTPnyQ
hcJFs9L7N1xKOC+sylTjp2nZUIcBJ2ibTn+4xh5nAVYvKMqifw2SYm89oQA97w81
NYNPMIpGiptmLEvQZrBDT8zJBi62Mg+rxqFp9Zbq58Ngde4mol0jybyymtIY4MB4
mCN+8TNo2LE1dlhCttm3o39LBxy/xkfOLCxWbKB2Q/m3Tsq5Y0CCr6KwExIEnfUo
cdw5ZysVPPSs+baK543ng91MOEsdQl4LTTlc4Lto6abNuCzcdyLqmZJGPJK+fi/D
FDHrj6cI9rKApWAyJ1VcweCN/mifjxzvRL/w/9nAYn4urhzWbw9CFmaj9hX7V/4D
CGLOSWg578161gOufsyNUoCjLgO88yXp5JI3htHRPMPDBWQWO7TAoelX6irvss4g
A5i7mlvxulpAHFlUv5Z3ikqjV/BmwOLALUocfEmzdLa4UpDqeCyH+Au+VcJJnNWM
5Ol2I1cpLLGiepGtwVjc76jAhLvyIJ5jWyglFmZ2gu2kT+5I+I35D2QVGNaxszkv
Y1J6O7yh9sjwl4cnkMaJhP348RMv7x/h2ospjSjZPh0SWJlV/QVbKygNAfX0bDIK
+xJQU6tu8B6D9Ya/cDgDhZvpOVMm/9F7FXMhfm15CmBIy5ASj+qMdEkkAHBqws/g
I8uDiUjYsOdA+Twu9Zvh/NIWy0+juPTOBNkCBpkAMijtCvSFFlQLc2D3Eh8oe6Vq
v8Ypx3vHdLKTODElJFNiYtHvjR/kCUq9YYbh9cZqZDZPsS13/8O2OJcCAdxTPbpl
0QKw9SvKGV/UsW6P7pVn0YxkZvldxEgoAfNWfuf5OMO7YgQFgAYaYUVCIN6ioV/W
VOE/AcYQ3r0OIzojEf/d4BWlAuzMCz6VF7XFJ8olMaNv1Y86QWLD6YXaZfrc9Ztz
qBlK32aAcjla1Wvj3wZuJ4rXkLdXZgZdsaN3+JMDmltHwTE2tyc78M0nx/ea+Zmp
Jd9+cM0blqn1fIotq/Wr4A32hxtQbW5xdK3Fl/FkvgjbuSWuMBJ3fPGKLcjjwlVG
6UzIEJ7IcpM7rAs2L+N1SJoBD7pbp1CY9s66a9YAFZDDqeolcHF12yjOjNEApIfi
A9Fx/v56DI/OfOGWQjraYt8OEWMbQAz5+r2CSxjGZ2/et/48pIG8KVKRDkFNNahI
Zf2AJxtP9SsyZy5TmC2Zek2vTuPKcPuvpG22VNloIzfajgddjxEh20atREJwaq91
7shrWrBJBhQycqb0L1i0Q25W1P2FHvVgYUIPPbUTvVal0Z5TWKAkcGwKSPG2x+8f
2bx1eejG+MRQfS/JcwY1mHZ/xKDdg06vPudBYEqyOzZIZA+ahlB07762KwRLglpe
U32AbnaBD0++sVoh/juVm0YuY6+vnUnHCtjqU0Q1CQf/xYuMzCjqsmfxGJq78/T4
CwEF9eL33VJ6YQROMP7TRBHoB6P11kb1/ECNQ2vtkKBY/avUa39sbTWMTDJgnrBs
nOPch3QF7Cs4e6iURahayHBSiV2GA3/3Uol8Xm/RNKWUYzK71YQ2rG0WuhwvMFF0
bkiY8c66vsMzApBfFxI+RGx1iq29fPa4CB2J34hRynpWZShdRxJiK9STnrqVGey3
6RCOpwvr3bu9UsXSKIlmkHLY97tlHa6kdJDsYY6zz2yzgMNLFQCMc8a9NeKuMCDF
RNw/VRM4dmW5Dsfflo9hNEOMnV2QZeztU8JmDePeoO8CXp3mLs+/JM6L77aGC05B
bocK4Csbc3Y+wc/yKoh2VKKY69qFScLHRod/K6w0udCKBX9QnjQ6cltPXJNL+Apy
n701vwOTxeJLM2oNYKvqNp7hTz0+Uzz2tvk7RvHF5EV4mFmVeVCxVxfWqv3Xw/rb
WL3RElc+cedpVcjX2+zHLbmaPhzjh0wycL702ysrvSxZDXQWL5mAKlca79nIyEk9
sizjUWUNajD/pJnyMzHsXtDUpdTYao2Bx1oTawOEc9R7vxOURM4ixAHck43HcJSa
9TfwJ78gc23lI9epQ+1DEbmn6dq9GL6ODpBxyuN72fRQcpplURPI5OprXIU/wFmz
r5FAox+m58PCUiwF8yQKPLecKz/hfi/D65Z7sOOAJxBWBgS2yv+zIqCQjrLSj1LC
uAAq4WWtaPFPnqszP3q3ciFyGwZ5cFX1LL95QXQ3uqoVkoaa65XC/6MWcfOT5h2A
bGePS/kUtxMPk8/+DFfdPmusCxvWTz+Mg36vgPWclWldSKwEb9aiM4xOYjkrUiN4
fC6+IVWt7CPkXo9vYioEQNsDF4lU44t80CdYh0W4q67eaorQZjL8q5Sa3KFoSWP/
/oUtVHtNNA+tPqH+0+52oZOFDmQSU/gkGsPxkTbLochoqxfILjBEceiZ+E3uL1hs
XFFEmTXx/lSo4McNyPnE9bu94NWPIoMXi/fSuR7IH2tkwIUWysm57+Ii9pd3OETb
9UpcTTi8Bu+o22Z1SUFlYoLkATeWjJmZTt46pEnWfYzduoM5/Iw33OXKK1kU++DM
Cn9HB5CJbMxcRB+tv0FJRJNSxCigB5M5dhtbB8DOqURYy2bO2pE32p4WJ7cv7flN
nBr+nIjvHfPAvOSrKSZJuWsE882/HPdb2vRkMwNE3/FqWqu0MUERegvNTcNvXiLm
lO4eFEOolsjbRA+osP5iyK4j+nKsptg60wMlk0XjzuBDqcWq8x+6cz69D9HXwvC0
sGbK+4BYMXBBoTo73bOkmPOAqef8RmNlxdnWwHAP6lNt6ee92XCJaytzPfM9ulpN
94dtK763k/TiHwcMiM/NS/nnNbh4a8o+gooYmulo+LkTE4VIZvEPECLvV2EBqbYo
eplSMVOPNBIKFkdXzbEqn5mKMeHepkODJJ5eUDJMQ0YZslK4qMeC3IJGwc1t/Ae2
93oBOJuz30O1opaqwAQhbuIHqZzI7JvdaYjGWVbEDui01ega3ebfpgd5LSnWf2JW
lWMFkeGt4BYjrDDwubLjtDbR2s/jaO3vVszrBw8utTtUhixULseiRM8w1KU/XgsZ
L7zQ3Z750NlDrcB0jxLVAxnvB3CXGv6KqJpFgsNXQsvx51Hb4i7AFvt84uZ4gywc
r/3dgQIwvCQ4+xOxtKplI2Y6W/9LFrlWaddlC6aDR8L+7EQkMGXqephGA/EWhTds
2NrRhWmzcUL6biFA8U8GnY6K4vwjBb2HmoQHUNgBDgeOWlxc9Ey74JcpuASk/81c
/QFA4iH+FnzK263BL6A/CCilpaCktWU/axZsMX7UoZFI8pMX0vNws1AYKU0u3ssW
WpnPy8pWZcTS11Yv/PCH/Pox5MDyBtiqO/YexwTKj7r4wigUtL012rqNjWykBBM2
fNKr4PAWFmqXiFq2cYq5SuGzszCT5sHCLcgkCMUGkzi/ZttOhkx1hnHKAx1x00TA
UwIZi/bru7+8qPblE6CJuGu+mI1hT1zTiok0qTEjIHKa/6dnWMpKZDaq2M5lWWnm
xWJ8GAk/C/mv4Itzd++k6m1MOid1ZNknjDOxe7mUVTzgcO7lags5H3UZ8DmyWLwB
qvOVtAs6D2IsOrQwfkD/zWz/RdafIZF0n4CymQmMzvpsO/UY0OOyYtcWr6BOwJmD
wicik7Q6xXnejuURse5SvtYZfoY3jBJgrrK5to5D/cX4LZAV8YorcC+Uk+J6eri8
M5E7s58JXYdKYeV5FWkZ9j64sG0HbPnK/J+sm449BITceElRs7CXq7xCU8Iwmtef
8exvs8XYSnyJv3YLS+FgpxclQ4j6HqE0igxjGYf1ETojchvhF9027z+veU9k6EUl
cd2eWIAzicGWRUOOvCmExntHqYInhEz6eF6c66sUZuQxWDo+q5BQeWKEs3Zl+78C
CVbVR4O7BKXPPb80jkqxcCNJBUYoGJEwKDsEbUCOpx87palkCRXF5QyFK87cai+J
s5LFHFnON0E36AOS4L2+phza7MMIJG9L9qFjCw/yj0tpyyXGm+gQcKDbmCTdiRZW
GYza0KULe/f/jxN9FVfqbOwAMwSfHhsjnYmh2PnD3Gh1YGDjKrP529x/IpL808ui
/hkVvx4Lf7kWMZtkcqH0SdDoyfdzRL3ZiPt6MSI8M5/ynrARtNGhRIO5nHkFkgji
7YtDEoKA429d6Z75ttrNRTialSqKiApijE51lIx83oC802MAWFA7UUVtZrzaeB2N
Ly9HG6+4KybAi/L8B64IcJyOpbRiiaQPunCuTQSiu7vDKeCWTVomWWz7zZpW5DxQ
etdAxrRH7zF3qSJsYLU59d4n9F7/766y2YegD0jcoNTHHLOdXPl7DZ7ROxVTrAa1
W+fcpLV8eKuHxLO9vgUZVVawBWG4LHmiVnAQIlVubj936m7sygWNT6fFW2lhqDI3
vNGivEcTqg+nAETulcYTK6Ay4nNwZE4Ji4az1ehRw/EEdm0mTzC8p9FSv4RP6gzb
wmKcBrxuXG1AJKGrXSkugPUfDtTxapEDGZUOPI0yMWR4hPR3zq46krzV23HXN4zc
nZXS5asU1Ye0hrCHftPg67W2zQxUTJbKEdYwal1vQpjmrhmlpvxW5Z8ABlR8NjJC
7TWOG2xsMBcjpCQ3vO1mnfUseMT43+V61tF7KVANEXvHUI4MDPna8Gc6jYoX4PQL
wJxKfmu1oSu1Xk4AE6zuhYs6+u+kkcnSS5KZQfu8BQK95J8/plybGPc8llRyo3U3
ksR6N7kow95UBNf5cUnvBIyOQQZ5Rv8iVokG4zHdjxTMmTgjr4LyaMd8o+jIDjxg
8EpEfkXsHjzjyf/mlwYHarhnv5pkChBpnQ2R9zbTtkSNgF9VXW9tHvXEtNr40i5G
e3Lxl7n6MLmzxPOBmSyzT6vTE0d3HgLq3rk6lZnJSuBZfEU7gUC6UjL8cYm9o2Ng
or9oA8uGdKpLetAx3L3STDzNlSBCL8FEje2hPcVCFJnynrCvTSmzH4Zwe7bR3n4b
T8sBfPh2vnhL/gQ5HwDTKyrwfbUJyZ3SkB29uajAERMb1FPe+dPsgo7uBnF38HUm
4h+OkNVlXgMim8eF7txANZhY1v+yvr8C3mEYVtuB86S8gietOx1ZLT6kGxs+mxxn
A3ViFYFRyy0a/7gyvnWB+K3RP/gYf7ZVNZ6yQKU0v1ccb2xHljkSZYf1zpwqtSg3
o3KjHw8h2NK1/AW118bYBztuhx2d8OqBa1zL2n6//q+2ln+ZV4oiKAiuwGv/++2l
tnFACGeBeeVDJsO38X43ofQAkT4LUL62kfAREktQL/WsawHaIAnICOl/v+WkVE2X
SYC6gVC01PbFuwrcmG2OhtGfXYaeIZnkt+S1y8mJgauJKKhXbjkXqiUCe7TF48IC
8fTe2UH31eHbjRnexM/PBSRRN+ZE4P+jRsS/kaIo/qRgmQ2jhr4rG9VMbRn0RmOD
pnYINJt+if7GJl3KCKnz6P6ANsz4DF4Ssp7BvzTEBPhFkJvwutYsG9MQW58gex/M
UXRzSdvSEy8sQFoXk671ktU+7IQ+WqRRyq+nkNwLLplnMSOXQpCsrx0Q3wucA0ul
a8o90ETCOuBSWkhYAaB8P2Yi6oZGiFxEv9I+ZjIWonWbdfJZOMvVUHsl1KolMgkC
j+mEZXVEIwUtjGVDADMLPQ8sQQXB6WGx6fIbBJmQRzbXyYSda6HRw9tT8A5zQhx3
J9KMruMuZNiOyRywV9rMoN6Qq8YbSyEem5PIlxMkZaT0NU+yYr2K0rrSfe0Jz3D0
J2Gj7o36mluSZvpagMWrumYVHUcW8uLUPZX3k0VTnO/u+9uMnXlPXkXowA8HvBW7
aVpavJhFhxhnifAh3TyL45maUnG4T7BPChYw1AzgUGEfbH+AwzWhbFven6yCxCuJ
z3cIGeoNYe/sLceD1hwRipj4zPGyZT3nkzBNT5FVvIAQpELbOu6vmAxJ3jr6YoVW
GkEgHJgVPRI/7XjPEwif7R9H266j8cOgbBq1s/tAOFcxYn0UjXx9ucIWKi7Cj+Yp
gYUjt4jWTQ7OpuqClaa9F3Dz/Y5aEp2AeUvmZaXzv4D34QpeWKjl4Cw8PpzH4c0C
p7vdnGs75qRTYDqQKg9I3s7LWvF/aadgCQuRo0G1Hl06Jd5dfH+5OH9aOOuDruq1
Vuw4fCYA7S8axsHRbe2TsOqOXYQFQbzqRtR8G/fYCidXNZXNjO0eolNzqohOogYc
6wPJc5DdQhILg/qul2/n+wCug3dhjS7+g0J1lbULbOCgw9Sn6PcVdKUIVvkmmVaG
mJen/GK/mb7v6qwmP/rdWE6YexoOfPY+4JDiggW7WCGYs1Xikf5OOGjMAfRJ7yjk
/6xQv7iIyGeo2Bm5t7DlA93ZTcQkt1NxhWm1MNXW+EicIr2E4pY4vdHdtazir+9Z
SXMrUUK6USQVsGlDIzEfHDbC5eylvCcPxr7JT5SonvOWzRCnvOA0zWYC5HJWSSz1
bhrnUUnmmgTTRZJxS9Ba7zjG4DolkNLz3BP0dnRFIwtReh6q4D3WHka1aEAxjlEF
X7D4WGwYuCY4jZKno0LpNacka4E1fLwY+8cf+sZ7Pvau7+8tIgCovf456Ki7ymOZ
L3KqgOGInxuJf0kcL2bCbCWStZDRUbeOoE8uGpR0BJwVpZYvWxnnC4EKeL6Iysar
3Z2CD+GOkKJm8bJ0xK2IUCc1fzdG/hfBfIVnxtkrn96R5IFGcymYoQ9xNp+y0AAT
GnA4Ydoroe6BA987h40k50/q2PptX6+ryq6AK/4STzpzoLA8jECN7JplosX/Zc/9
bc0ZZoVf+TGYxF6wQqBiZVIn62gZRNtXL3mnTukMkX0Rf9WJZAyDEdBQ8Zwhuydi
eY3ctA0yYs/5q1+De/6rtVqwJyecnisyEdv9r3riLUHNiavUxCmHet1Lk5GtPavl
mCsqUONzSH7n4ViWwxpVxCzPht3HdGDaHLmAwGkXBJ9VcNHIPGq/fyFILsQBsAr5
vcsO7roIZ7m57yirpghgs5QvdMhjaTteqEm8WM/UnSbe7IJbfsehU6/4RwYf+kcf
GX7fNZ8vD/zvfaotiJZM1p8VWN3oVFc53waZUzeZr0f8Z3XAiBWbPPnwElSTgMAL
DeEMOabiOdoU27HCuPQ4ZrdOzMu/wtL6YFDG1yscGDZZwRjaTRnU5yzMUCwERDu7
11TrIf52fo3hmgSc6l305ahpot+ylXqJkMyBdsLB2DmARLsoxilgQPw6GoRSJwcV
EThgNSp3aMqDiByeRPgMYR4lSSwqAH2dM/gS8U8zEnSBgtPn55QU1rFcjYRApaEw
KmGsUA19EM9H671I0vmEx5ENy+SMWnvI7tTZOLLLdEsdpJhZKUQzsShspNcc5Lxj
GXg2CBJ8zX4cOorVdORufXxzgUuXekHMpXaYhL+n0axjh62yuraxcsrZxs16NzyL
ZjHmyP1ui4ocUW55tjQjyNM64S12LjKrnFxC5XFtTsjebgcJ3yF1u7wwrcG2gSJZ
y0u94buiPGRVdoj+YTPy5ccJADx7MuZTqMTNAZlh3iRFqXP8idU2ZYpM7XnvRabJ
sH2yqRXQjDQ2bjskaosZmwHmBSeHBhBs6t8tQIDl4LwRfm+2G2Ey0EiWBnILkAbH
lM72aZAjX2T+11tuZpcWxacSJILFsLip+BBD/JD2/HbgrnZmNGEGTCHqxBNekRkk
Ov6aXExi9Zlt8KurLJZ2Plwqw2cbDDytAG6NtkziVfBiR/ZxBTeVfLrY4QpOCkA0
zLN8qj7iJ+dAl8vNEEdJbBvtGHFoMof3n374u7X/Um3fSmV7pxuwoBS2wWUU3USd
D8G7KnucVZLjsfAr3lV5DpKJXcexo3mUgMn5SYYNVZ8yjnOuaoWEOjXCx4zRLzk2
csKWTL9JRjgsbalIZa/gqnGPHAFL898VZH630wES3BrLqDMIsThYc/JOrFF8Rv6n
aemGBUzVoC+eg/Jxa6o9XmxEPJVO25OaylHT72ON9pku5DzxnnnI77BDvl4UzdUF
42ZhguGZyXG07GBB7IJRjREVOI/26hoT2XAVNkA3SFnuz0s4buvidVsaJrcGBfcX
j0RUKx8XUF9NII/Q1IHornq++9dbqnClni8849KgS665tYzbHU0s6xLXH3omRyZ0
r3GQzVK8Tp3JUzGrjcv5ae/3imU3yonO3vLmrlGnAFyZeThd4wFBnVCFz5esB6IU
JOM7n3RnfpHbsuF14EX3BlhKDANGIj1cn6Lg9sTpaebjtfvoUvXLvhP2dPJMolcw
sZ03GHUvq3JeuOpjRSp36ZlDrCxMIvLqHxjTNgqjAEx5GkQcPdDodhJleto0UQBm
tcw25IW/c9yP/no0OiiMfJhNRbHN8FOj/BFPfvoJ+h/3tuaIdLOa1Ulr6yTIR2po
znig/erXv+sr4XesRO9NjIxvHpi9TQ/XzuJfiot8j2X5yj/JvAOBdUrNIydvmgLb
gt9RwfIHdEiW1duSHCIjV7iQ7EHy/kjGcz8/mjO0Fvfiul8afZN21p0Gq+aPy0t/
MAIB/+wnWivjRRsD+E20CypMSXNIJvYqA4O04k2auwVpXefZDE81hnDdvBCrtCjY
lF/fBxveNjF28xaOHG0+5D5X9z/LoRvJLLjMo22cusxzhJhbjHhMoDF+LNBGt/2Q
gCru2RQxldqc3o0bHaXj25Fily4gCOW7eHqmTPGWUVlrwNL7cLFre90CzYeHd0q5
QVyfJ5HmFylbAs8vAUIgsXKR1oA48Cd8+PyQfu53n5Rnj9k74UzsB1SdyCly2tti
0XxSo5AEBBfpGUB0rPqzCPnxS5qjKmygtP6DqpF52CP0BMU38DBfLwZ+t2iGmrYZ
pYFdgNd8WnRphi9JUmGMV9r/dlYVBw9nCpJp1NIWlhc2Ye/AIq5Gfa3MekqItTVA
0uxUCKwuXx1BGtNhhns3YJZuHMWbkb2PrWoSs9LH48KBhb81ykIV6b6ExDo0tdN6
xMXZWH97qzyWlNsTZvEcHrJh2gIp0jxYk4OC9h7ZwD3fvxBGQlHeMtP1wCu7HWA/
zboPBVcRcSufttp80NeQkw9v53yKZXmdeV8DmT51x4GuN+rXk5TDSSPpG+rrwc3l
T5Z4dMsyIIakk3elPKSuUbLCIQyzPEGlPSNxf1GsiaErkhVlczTUYGpn1pzHmGVN
d3zoH/WZ8+RXgMv66uTVCPoygWjHE/25zI8GxYqKPquUj+OpUmqWw1wZOhpLxS7F
f8nP7ijtwn4Fl+gJOOqKFqmzRlZ5Q/M+tDONSsnmlejuTpkYIScN2fYFYshHewEv
4glXTR3OkEgj7Zet6Cc77rOf/8uGk8nuyQfAL944THKMvVMhuxta2BPCJ9CkuSGh
VpbHNynycbkTHqBt93eCQPjJns3P2s8HQIhlsCYGZPfCBCzgUev+ALe3b95007zF
6TWeT1qeUIIPX1N7Mg5DP2kwmq+6kpk6OFa4EWQ/gJm/6e/2J5UbDa5FNLONxt0/
6FJzscMtqkdQ3tKBdZlvxV5OSSmeWPkCJ8QZsWAUOYufFPhC4t+K6Vi1oTjN3qvO
pMJHW+fCyaUdDLQwN0xnserMw2dxq+NDr/Kovq07rrcJbEF1N9+e/GfPLJ+uYKc8
WhEfN0ubgcn6oO8YCrn8Tqsa8JrNjEV2AREhLKoj80DuF5G1aKmCVhbSzrIvduRl
e6PD0Pzy0gUtz9ao8qDlba+EGIW9kqK5/gBXjv1c6JvDputbsX795r5f/r3y24u5
wSTeNHJuF7M6pW+qlEPqu4833sglD3Fk2AaO7F7SLkLvduII3b+Bk6bY3yD/cw1L
0tFroVERrc41Pmfc69KPGDZaXav+8jV/kqb3LGAQDYGcUa60M1jTOyFV2m3lt9ET
WnPeNViFnKxzU+cg3gf0C3WrpjzpjDwNyHabgGFMPgNiIZGLML/6X+PL+XezNvBE
N14abC4LNld+ePhnQ0pk0SiHOJ+EXeLtp24S7egKnyKEVC1c4zyGhDxFcs8rrpKj
ynEa0Gqtjj8Wyd6v2LH+jGqskVW2HYvki2weOd+y91sMUfVsGXUQrivobUGQBrob
jATTgr7u2ius7uIZKyqhRsemFt9osK60WO6Xmw2lkRwQMHiqQDNeFgPaxpoK6T1w
NfgOrFqfzNpgFjJUPrpxCDsCOV7/FGE0GO97FcQWqzaMnMLAt7r1Fuxcs/KbKVG4
j0UYdoEL6fyV/Q/3MzLYoCW3WXIiTvaTfVWf68nVc0GaS4ng91xCuxIKLlARy8zO
cWOmcrRmvqhmBSwIYx8c+nZNE6CWCvVTXl+zFAbFCEAJO4rtEZYgU3QaQHaIkoLF
3m/q/610PFkt+ZCWlVcAPFUBZBQ03dgY0ZAGUqxY0XHaNRBDn8OCdsXjkZb9ziea
l9iqi5sn4osJMtFXCl7UPTBSSnjSf0xpYicNUYWMFArm3Z/YnPYlh+zEdTL4qwhj
9+wlhTvtFKzYVX3F3KHdPQ4NO304L5IVeRQRRvNJYdU0n6g1abVaX1tKO23BC/Ln
mzuxi6GkwoXJqpMdJ+8ckrW2Y8zmzaobfwryG2KwvpW4EmOloEcA5/ZvWV+6oDLu
nYnErzDhL24VittR/DXe7GHFQqf5IQtp1f1tzRoe6a2WT66a4Pah6UUXT0hom2ey
l1voC6XBZOQj9kWYxTJdVy/YrB/FSNoAZ2ZHZExd1mJtnPR5xCu9xDr6GUdTZUqU
suMyf1+5yUhA0ZBCydTwFndO5OYLd/bALSxaj4kopmXRuEwPE5FiIr6CJ8f7MdxE
VtIzSKSlI1z3mRsK1Ran2kLLk6to1Sgei/gw5xhDapNso3umbaZ6e+wtJgebQtHr
MdsZSdhoEQkhB+UP0dxpUCfxeRGHsr2aNoTJTBrCB34Burao2C+wfvqG2J1HEUDg
05WOXtep8ekbTkgZVo/iweF5Mq1GO9ArRPeqNnNGQrzHHhbcOmqGCFD7fq+MtQLl
qOkIHLo1dEXemcfzVt8v7zH8WBhGsDEhdRArixW+/2BwE8GjAvQEpUP7frXlwitN
aFtnRl4xhlxLl7fZRFczwbq1mwHhHHZBr993S4bl3AY2b2KoU7k81MgKxFjuDzk7
Ug8wdwoHFyzYROkNwOdYmXmd9ofedFllAEF/ldNFEyiJpNNwxV08il7gkJLs+820
w9t0pCr/K77MDEwkeFvuYfIjh+/zGY34aLyahQj/ECE9mRyVhs+b/kT876hu6oyp
lzU4dZLSoQW+yjw61rOk58PllFZEm76ry4Jf8y1gP1LLWc39Y2AEiwwmb6wM3Irp
6pg4J93XMAM2JNp0WstUZApc7msAS/6WoCV/PdWXb1VMkcu2WQ4sZCSNZ86jmgFh
t+MvLtoGBssEtRS97SbcfLOjEpELdYeWdx+7e2C1lMgZ9Lp5QrkqE4zDpiu7hmY0
MSVVnseJ1OtnpUP5BMiJ+T4giTbL4l60PshzWlxw+jHv79W0pwYq3ugx1ET0DPYY
JaIzntjUQZNCTeWywAHST4MoLFzTPor9FP91hc4v1mnyHsJMWIUgtTxz/Y62CXkV
oTjxLQ8RQRcsZgGHzwI21e0YrX/tiJVnC9UlDGMI6KxWZynTVLDODbhcDuyaHKke
L1NClNdJ3PtkmkctJgpw37Z8Mqy/bEMh/vJusItEJfqQrwIJVJu67yTy96c3S5Pd
6lsTL3Vy19bUE9QvzwCSoPLLQJnRRZEPzdJ4ut3T3obQ1DDaobCUDEEzH4HnJBmA
VPZkYOqfcCmLnHUJdPHAi+FazpLLJ5lgvU2isC431B2pVPZjagwTw5ACuzNxAlYi
gprfe0wHMmU/b8PM8AI58G4ehG6e1K6Yo15alvLyUcQGVlfzMnTM/A9XtqY8fbpv
RkN07QsFgiN6WJMRpQaTTgA/HXu/WDH7DVcoI1qjMJYjgnreNbvz5ylaVSPw0Fle
AbbQS6DLzqiZewkyjvUimZJASlQig2JEEwE0DoSwTUDNQvhG6yen71Iyr1d/66S2
E2ZiQsyb66eXsVfTQTr5xkwmZ6yDtwMZyDytOnShcmTyi77l5NuUMN2oba3Ipo46
ww9NTnfkmbnn1KYymaGFDDRgLHGPGeYb4s2qpf5oa5JkmAUbWddtCVtcm+84Tpmi
c+NL6SArjRjkUYToQTF22daKjG2xG0+CI0MtWl1FYZWOaVG8c77xiFkUZ88tMNLC
zhgK6b+/v+WbRbAgRoI5+WOoU/fueW5ISFe9W9TQC/bT8/ZwpzDklEXJ9/nQ6Meu
JX6NMojz4hP9eY7nZem0LEAlDRE9nZkuWInCkAY+T9rSmgtT54B3LfvGh0VpKHDH
mWzBIl94LnMOPIwtKnCx9CcyebKMVK+X2QbPMy/B+QKBgDFp2R7neuexiv3jCul4
iKC1/Acr5VWwfHvFllMVIZHKaPTfRyy/Je0FiiIh/M71nIUZpq5fIZO2WZIz4SgD
P4Sizi6nXPum5EmbJW/bFY7WfJIFKUcBKfOFYfD+qWSbQmLcYu/zB0fSK1nQ9Mn/
KdnNBbmDZKOMz+HNXhxIhjS3uDVpKGuJqRGkBmy7WTghE6Jl6bSFIwqU30/bpkch
6Fso1K8BcyLI7sZ8A5oUACVKPZiGl60k0AY59p0Z3p224FSSVk1Fn2nQ2+PNDoSj
d4f0PMRYLbgXjS813zXlU+a+894lIL4/rNdv1VJquNZUGiGyolcCUi8yzuKQHTRG
xuN7MiKzw+nLkw2QLcbC7SYpuS9tCCqHX8vWsTjHgjBYq3wH4JFDQlYS/pJ1edEW
lnpDvSsxgZlYNpnqPvSGY3RXB3yW5QZO9Fpr1a65Zp3fRhEdbXpQNXnqHQRYCCC+
HakH+w5zxaEuUMqMQTIeigzKz+24ScBA5ZZEhsYIxaSzIFl+afKwKKUtkjg28+mx
SNqzhrhfpYAB7vEFz5nWP0PIpelR6BfczV4GgjsFyMUyAGEEsAsLINO/v8HZh/l2
k4JDqS0UDVB4eKFC49dEpkCa2iTpBDJstyNY/LtSZezrRtGKYoNp5b7MXkwHyRbB
LANE4WHi9I/SNXpt04ldCnwMtMYNr4HOp0RwUBSBrSiiWjnSYi2S8MwXgLyxh+ok
0ScHuAdMJpVgGGATt5DshDMRCopmHvEGnq9PEmt2B2DQKxM5HL9hgX+xRN+EH5Ny
6DYQrC27gK3bZ5++r+m/CJvsbX9YVGGUoOnKPxpHuDQ0Qc9AOtZvmzxLadio/Xkh
NbhwSE25W4YCVWBN2aRM2+GWNtBZ94iDT7i/DnvjFUuHoYWMec/TtS/KG+jbgHAH
wIQl1+/1fIIi8t8dzET8AwmbdCvSZgRrabkI2t/qooT2c6lGXfk4SW26vuRbOzh3
rAI4hpZi5SGO+v4g9FeJtiR+OJeMshMs3y0qX7Wx68a1Rx+wx8MsCtD5rqgfz5T5
Q4GggLRSrNH5QUP0J7kcmfOKW1MrM53zQxIw1up8CYcGTdhdtRJSd2B6m/lNDppj
veyQYlDBexZ5BaNfHmBp5IfA8rYTc3/Xx7gsDehNPSJsXKe5SLdRykvJG4eaNXww
NaEbBXniEiCqpVXsmMEckp8MVUAQmGbgPEg5ABaZfCDeoLfP6y7hQNTscb4NHjGf
7q0fAgUE2mkisfsUOH86PhelM0gOerlggyhVq2O8E/s+Ad5qGMcaC1gUziJM6xLD
uEKKOtw9+c3e04qNPdtnP1aZ2N8VSn0vubgbfwxp1stBKRhkISepG4ymWf5uWFXn
7FK4HSs112QFischQDGOeSiibh1X9KZCAksof6wOtRvQuCi0VpKWsw3CmSwzfby7
HxIXKVuBHzxAKRmqZ1HoRR5v1TS0Vl3r2V2rLuu/2jwVnTBsKLw0WdoJIEQY6GVR
Oq45N/PM/9e/Amljc4vm2E9jAytcTmR2/lzqgtVd1MmYgFp8FcW9530wXOBOqnZQ
SZATmLRmbFlh397PUc6OjhAZWMnKZGwm2sq1HTNsU6WPWe2ckRKta9J4HY66rRbJ
xp7stIG4Vw3ITTZ9vtKhNw/60+WrpNVM8QBROB7o6sE8efUrtVQe0/E64khX8f1Z
hR5RTEMn9OuQROTuRvjrX2skVagWhRNTob/kpayx0zEvqiCdYTguD43Ff5Qgh3sr
iUY721Aiq6A7H3ZO6VQhix/5p+CBH3Yu+FxgPKfPoDvTTYqle3reLXHDowSJkxoG
VQ/W1wosFrKZz1wTc38DG9bteCxQlrVXehawjqeyeBH1AzFP3j4hXys4vJClq1MW
kyIPLI3kg/0nD+Z9btRrLdNgDXuYOr/DSqyzvbWde2gDMlxdj1AIQQ3RH+ahGgFP
CujOflyISeJ0Ky2BmO0OwaS/xBaa24/lrlL5gZM8eAmD+YKAdWbRRI7snGALrdF+
00fPj2s5fpaTC0Al3LPx5rxmNX/RUQpjvUWIeD4vXy4GKyhQANgsGEKnf1mFTVZl
zyQMYqd2oyvU1rl67CdyRbk4zf7D3uLn8ZduN1vAQ9jv7iwH49E9pbN2/5Pr7Lp4
4rcc5z1Mc4ozPMUZi/AEcZ+rI9+9mbEmQRF5b7Jb6zUSSj12vNKWOCBBXXomzQkf
cNZB2EVJCbS9nte72BJ2VUSkFzVM712tmWK5hd6bwO1Yb9tRXIc/ABDNLEfL2/kd
5wonRM2NRKyTWlgZoOx1jn0zLFg5AS6QwZtnEAzraQtJygQXVBTPuc79CvwuW9xU
OU2RdnQasNFbFpDFVg5POxNfkugtY1a+ntIOcwe5EAhjAbDV71UtZaJOlXz7yhNh
r0CJcyiZ0dLVntS9M6utpr6FcJ+C3OX+OwA2jpMhsq0g8BVRl+kGqJQuvbaWpvMv
VgHQL23814EdE3Flii8/0+W9GUxdnim31deoH537EDo6sXczlEl2CVrgE2G/rkor
JWwUwCp0jq3+54mC9dLBS2j0zQiw802x4Lx2QD7+gRUIeYKZWqWKHt1DVL1RuIs2
FMD3uj/cW+0orUy7eqJtwLYoL2GxjCe/gq0e0W/rpiJ/oA9VngUJIDvk20DA+mBN
Q5FZsoxrI6H58WbWFZIUxfHglqi7tB+SeofJgfpU5j0L9P9FRCtqnjBwElCTbJw0
AifqS7h1YS+Cnad7p0EKV77fz2nqdDAqPMgOI7kzdB6a9zAPNAPNyEU5n+uGm1xx
ddnVVoL9xXdAEGMrsezBPzIxfVjuAn3CbzkWhIlTYtH6914kaHD3YP2DS62uJG+4
7RZ2AstLJAfsf8EoKd5PIe65LI5rQhbl+EunFyBelZPQPo0McD6KoiBmbx7GQS4m
XAj2/HqyZBpkhUQYJVte2gtiaQaYMBSW90HIBpvVleKGA80CZXSBUa1P2+bCZ8ga
Uh/mn2fsdTQVbegXvoDPFaKlUA7K5bDH8Ls1SZGrbwGTq1iPhAiTrDmOZu72eh91
7cujZaS25mB/n4RN8Ep0110mXxpN/bvzRYgS7eKLlmhrHUhwXrdZBIo52fYOMJ6T
fw7JUIlQVnvVQI6jpWmGrO8dfYAUuw3Uan/D3dMpUCz3JIAOqfKC3JijDNnRDzYX
w6O2AkPS3fScdE8Rqs4LSDSeqEKxwlLZtpfqnAMGZ2oKoE+wNyaBtT90TgFNeWJ3
P6Xn2UHmjxnXRo7HeuIfgZVTDkgPTy68TSzif+NFBngkRVh1hUqpk1RKjfbdWjoi
FZHugivDKT5DkWtqRDzmgpAQWug9J5N7vbnmz4akXnJ6oYoX6Q3e1mvBXWG72f31
mdyQb6NoiMySFIC2vX2lkoicOTVmJcOJRGVigiUwg+2Yds4bWp3IUCD5Gip8OCE3
kOSSFOTSYjwf55axInpHN57ExAu64SKU8miS2CJWxz9TCLf7q/a5LtZw1MLSzn9e
HOgzKuOi7kj3eqpU9atB+PQbj2o8XrzHJgiQQxmgLZd4jiHNzQigiEkgv2kayp1O
FmvxRXNfhmd7ts+RkHRxOW0Cp53C8jfCtU1fNh2kB3hHHtAXojasgvFgwJwfK3Kh
jj/AjvLMQC59i0v/cnb0rmTNSoSDg2C2CPVYzOhedzQLD/+I/caJSti93HiRqyyQ
RAE2ShiB+y2PJRctnqv4ul2BGdOJqCl5rYYmzzhCDoB1xAz3mObkOu0IeyC5Uerh
nKopJQqG1H3/5B+Sq36/12PzK3+JMVfSnzNBR59a/oX0SL7Og4epd80+LZUC/31J
fRG5Vfi+gkHT1d5PWbd5/1FJVAugwDuRvFxy4otvBIzwfuj3lLGmjG1Q1XssTp/h
iNwPjeN6V15W6PCLmr9JY5TU5IuZeB9VH8avoT6lxyf8k2l5rv2Yq2d6fOfrE1r5
csZzCy6krRLxCJDYBr/j0ZyTRit2WcEN8qJXhcA2Oq7n4VDmr4n8DueSb20M/r+s
NVKnfSN+peCjWDP2T6JBKi76aSr96nfb3QXr7vfV40a37JFqv59N/08ZdpSn4I/k
OfswPAwSH5A76o07nu+r7dCbl2TiIdk6C0ok/pcfbi4zAssvt1nzRmWksdW7i2Sh
tPhl28zu6o/zZC0js8QauyFv9UOZWe6MWIBSTJycLG3tPiiICYFvStISdylUestd
JFXC4+yxn3shovof5+mUGWduKsaXndzTRn2BFSkzwcw9feO3Ofeaeo1BiIKryDq9
AXz+eYrU1JrrRw7VBLxg4RVpF7EU8wLolEivYseDvsR8Qs9Lf412Xh5USOKV5hPs
Ab8TlHGRt9WpuNjAx5hRwh/vUAAdhTBbi/lE1NyAYnm9Dw08z9vZ4/fAQQDgHtnX
P0GSjTKSdhGvCDK5U46ZgfQ38uPlH6WtKBa56x3s59Q1Q5q+mUbRzmKTLFM/Nobc
e/46az4Xa5EtFKqzYB3TgJgOpc1s+b83SPqOuNwke5QazLI8WD4ZSATz+Msd8z2i
VK5G+97rwr2CroNNn1ehS4OWRRv+VP4E4HYj84u9SSNFGQ8ndcg1SWnfcCHGtK39
GpiR/wcjONucpYAS5PMtWuya0/KlHPceqsoNwF/xXe/sXxJLxGKzofs2i30sL/JM
2hR4vOUdO94T1ZKpEhfLiM9RgNo0XdVE4SIk9iyl1R+sPBtQYoWV9P17kCfNHsDX
BSztUsHQTeTS4xeSuJ3Imup98JA3SxoqqTg8BxT9bZEIxL5382735IMHKvil0GYf
bdHEo0KLFNQsoJhLTIqRiDDV38JRlFDhZEQGL98BnXoMgLR2oiB3SdYPRNdgytj3
ovJcvaDNVPqerYRMsjaCEjMRQ4cjQc29NXwrz2k4b0YZjoryHZ/9AEegPWU0qofS
B95BRW04IEJBz85ky9y52Xvp4gkmqfwD2vSM7Y4ISW98USUijUfk+S2LiLsG4RPO
pMNTXnObdJ5lTyKEB6wGOnQR8mqzPp8AdBX9hXepeyjh6iTkqVK+t/rvnBcn7huf
9xgFi2NLPRYf7kqrm3nzNSKmdnbjBNp9cpopj1yGyrlSuCXVOyu1vnB1ShkxnhYW
dLsDUIqJmN+PjwwHvFdojBoNyjBkI5ixvRfC1xO7w1zaIxGwtYA35gpsrebr1291
qmO8JHEl3/6ozzNSsd+ucdxY6g1KO8fDKs5KWTL4H4sQFCWZGBhMJ8eS1itK/xvh
sNV/dJEx3RL86o0fYyrxMz3BmUy+GdOR1md92w856igrgu/OFYv4VOFgRFZyzYAG
1YXO6/PBZsGmyGTj7maZzID+apzTj2J24uCCyd/o6dadfibH3hEzmQ9KuwagPpwA
MbyjwDIqOgMThkOnykjMb8hcR+RNqLG7+f+Rxzy9IhYARvcksTDbS5O18wdV4mJi
eOPV7eqNGERUAYqK9TAJZEtEeWIumOhkEOI7xh7W/iAjFjcVOF8VRiMRF/kU+ORp
Gb0D2f0TOecmis2BoMtjUYfTv3NJoClVVsCkMzadm/utSc/xMWSSXfklLm/qfRvF
MU60gZjXMjc6fGyQQd/kj8YSBGGNhMgE/l0D0ZMmRiCQbGuLlj8nWQ3l2XrOD07q
6n0HXkQSi6JlokuIOexJ829V87uq2QUzMb2XozPgCe0aIr1EE8HOZ9lRmKLNJUmx
E2PAbC90H2NWBAp8oFzzS4oVnrkNiN1S4vW+bMPvM72Yk7G8iFaGAf2gsiAHjsaA
cUvEwt6NKHdGtXaoN/Er/rgycbr9090pswZ6QRVu++2FOG3wG78olThRyxKm16yi
8LrDwxZMCHq6gE/mBIQyrJMsqrO955wdY/4YZW90GwGN5HEBE5jDG1+wx5lYoFWh
qzf8seKrDbMyCK6evVI1k4hLxBd4MecN4hEKJYajAcvtszkwcv4mmKuiDZG00HLt
w7fONd0eotN5lgBCyDX7jICij0qIJ/BqYJVAv3PC0Qisi9K6RI0goKHjJMWnY+8/
4CSvaEpeeun5jewuzy0wEHQBA4pOAtch19Gd8ZTgoosZHb009uAydedHWdrwkKko
5VrQGJUnpZhRY6h72el/lYNXKdbBDkcBDvd3++uH99JIcbg5gFw+ygyZZh78ha8H
Fa0Vjrv4fHhPaf+l56b80y5yrtzvABu/EqOu/14qBuIvrcOU4HaVHykOkrzDiUch
lVPQ1eavgQymIcVPe44U6rtAkZ30Pjwo4PTGjG5yV7yypUqrzA9yIhKqR/D/Wmm3
mhvp5VkCC3jyV2EPksfdmT0iL4h72sb4WAML6K5DpFS7c2Yho8XD0DMf/SU3GC3i
zpdFtqy0KtNeF7VIWbdMu69aMuGsyNOgzZN6Fv/wzsLI8DbtYDmQdjzOE+EfQTxG
OyBYDmlWwMSygcaSlP7iycSS/4PZuY6zZfOEj5ENA8gp9FROey1K5O+323XvzM3r
dsmNBOt2xfgfmOzOizsa8zQQD+KjjjoQ1IGJYG0vd5k2Nf+S8mt0UP5WtM/dz8Bd
tUc5/ETj/RCkGeVrCZ4mug6qARv2n5OTFgxslKKgLzBob/pxiM2avUkhvjd/V1H5
9Og5Lw12YffgbTE2CfU6dh/xEdNE5WJeyQbSiAyX8rXOaM6jWcBOAUFI/DCgU/PA
7+mKYNolNnyaSnK54bVPo6SMixfQ7/+L5kP0oL1qS4MeznSvGXX/MWq4pRZ0eV6G
jwCckdRAJrQIHDwYlO/Hj6vXeAhy2tCLPc7uio9WE7VgBAgdW9TLvPNrvOSU0S9M
a6sOQxYfHeEevlLTFXUo6mrRIGZShLHteKTqkQNWDByxss8chIXtiaNR47L4/OdE
rBtZnrMSsI1F32Mo2PIHFECjfmMmZRRHRYyJXX5YHIm2fDoQoLBr3qZNQZ8iYpM+
f9dhP0BbIbD7QIUrTVK6EIMw1jZwVQKv0ugVFqhs813fSEp9R2vxr6dUfsbCE5jB
mJ5c5ocom04Vs6y2Zpw0HZ+OnN83JrRfXBranZ9vQLSaXkCQeOJxzYnljM+5mCBr
2pmOWPsvc7UQtgjyCmh1rFaauuRlJJ6ibkLVVcc2YtFlGnFXZ+9RZrrNJQ/NRuPV
BLpdwSLAXNvtmA9q7PJYCi84EVC8+CbsiM1RVy5paBIuHtfdM/igVk2WmdpIIIOG
38C0wFnHMt/qyHv7j8OAbjf12W+P/enGbfra6G4ir0e3QqR2DELfBjS7S42lTloF
BN43/Ay0I9bTsy9065DLGTJ4/wCqIqNHqp2rxrU3vCVNrDp/m/lvduHAo3QLDpSm
T32LiiS2yFYhoGJtzLli6C1YRQrBBjvoz82/rAy5I3LtYwIuZwhPK5uQ4bBYIfSn
9eI4vHS1lAE6mgIxM+AAAqaUXY+RB/souK5hdF82PCRH++k4DTKa29kIrMfqs/Gm
cqTwyOAkP/a7uc3C2SdaQLzOo4a/94z0UgBsegCqwU+yYpA6RUAlKVoZdYZSoGdW
lYy/gI2De6edelFKvJkszhri/fQ5P6Szc3BICSNrI1yotfSINM7pCxSgLbowwfPI
Z4XcHsNNTsO01qndtQd98IKBBsFZu28mTXbRH+PxqmHdOIUkYXEMvdRaHMrDIK0K
Bxb6KWhIutLwT6fSM2SQFkH3PvW/l4KrG8bho8DznlIvroWSV3vUORXEmF3GacOa
fVQPaDg51ent7FFQyK2e37JiDgxGI1e+Ayc9YhaSy4/ANGmUc04609uLQKR0nmtl
OkLUZFVlL9lh3Hpvj/p5ZL9wphEYSB4fQSJxvd7vUfVPEmS9FoWGafOB3GkbRzJj
TXcCcuQGsf01jYSp7/Z9tUFc+X9o9ThWr4W5IMYx42LMYmkZ/ZCFfir0w7GcbP3K
iFQaYFJfyMlsaILGjz1WnX6eVe7mUm/Jl5xa9r0AmtMUD1QwLP5qlllaSNQWvfd3
u1pVfnhTdyIFa6XpD/hTApy7Qi+39tQDqA0tHrBhJctGEvouC+3uSwhV1ug85Hvp
0VfcwrgSsdPw4r0u+3xFMnF35wW2FXuTJx9AkH9ElY/qm0owDlZkSBz3q9gQIN3W
D+nLfXFM7rHrHl1LtRMYzpemfnEXkAJt3flZWI8oYe4Hk+ePlrEbpTzzkaUpeqMw
0nedjSAXGl1nTfg2SmTDauEL+xx3g7e+Kofta8bk0tgW+kK0SoFeeHIT7PDzF5mW
mITG+XM2CmXg+VLkYePXTQobW1HNm15Fp9zwYeDujH88FgcpVmnthUUIJJTT6S37
VUqQMVl4/JuC+btwfVN08PDnN2lo4rceeNZXIYZGmFHz4r9Z6D5X2gksgpslUYWt
LDmeVXwBtskDydiZdZ2OZFptYbC3pD6hKo8sI4lcoxmTCm7sas8hCcnzW0J5GVLw
Kquo2yXlh0jv5iCR79P1M38jnsuXPAuycV3xOfVkD95l1VOqqOsHfFEVLWCHo9Tn
6A1qYphSiHHNV3fSQr7dKnrAE6mM3BsAbK0jLPV2g40KlVoSLnm6YYH/S/ZH01jl
wOH6ZPyWVKOPpbRlPwiI3Q56Z52ekFMICcL4RZ1gYb4Vtse5gfC7mUIJAMmw7XKp
DyXYcdgLcVfl4G9hecV7idCEwMCQk9w2HMBmQ9fy+aBSqoGS8wuCzj0QpfWEbAdk
+0xYDhuwpWc683VnZl2ci2jLky9mlENK5FsHkSwxuj0mgQAHEwpoZ5Zmni6r/MPl
Gx+voLEC5ANt9p295LV+v6vlO8EdHiI94bjcJDXxivwOa32Rt5/X+uf/SLfqD1YA
HDH0oP83sy5A+R4xcEPfSFls/ekEXniVKpqCIVY5WMbXYgQ/Ng99Wtix5/ty3CJT
5DGRKoAxthBxQOt/y6pT/GM6P4s9yaFsHSpkbt7voxASE660dIJLwIpbDWooDFH3
tUALhWJYSUE9SsH3nloCAVVLKAk4+XVwHxa0RRUMrec4u/IlqdJn2ldLDlZQRXhk
a5Dn0IVsaRMOqBzjBUsmopTKh+lGbQe8L566z+8FZwawVyHCX/loaR03LQEUN5u/
Yic0V1fPRqn0slYq9iylndfaTq1wkG2meOlWgq9Hc481MO74GYuF1KTKkyXiECfm
agOhfVwo33gj23rOEx78O9aOAb4D1NOyqPlAAl4Xv36L060meoTzGKScW0OryWnY
GLCQAUE8ugpr3SC/4rcX92PJzzbqDnacbxTSyaKxuKkszJ21iXFqmLVGdrScIM5x
qUU4tul4EDWfdV1P2bDyQf2f2mvs7+p8dI+f6z//ZZTIgV9j6sOibKMxERio1N+T
wfPwDS/q1m68mmOjQSCCHi1sQq+yQoXeq8UNCzo2K5se0dH44TvIprk8F3x90CGV
doe6XG2HSvgC6OE7MQZyd5IQaMZHz4jqVDL5refGTwZ69P+Sp2ZvtG5OUKSWOfZf
etv95TwfC0X7k4qt0P5bjM8tewg1agE1zeNaMMffzk4LCDtRF7aROMA4/mRcUZFl
ZKnhscfnHy9r+pw/Jb+9BTR7WvrlB+XLWgp9gUZsUrd14FVpjyiWJXt1dtV/Bao6
JFsRj/RvTQSryvTamPuYSUdQXGKU1mY/hAhHA95w8aPs1Ihvkbkc4vYKzguzxBoA
bSD7+rl6otP6DTspT2stf97RX3rDvIiZ5Aj0JVDlnMNxlthV4az0YrSixgHvsTyw
si33lLAHncBp9TPOc0xsGb8PvVW5nGLl44iY6naehtqZF8mka5q2meHh/INv7el8
sgPuC/vH+4OL+qj4T1dsrUyyYneQOxeT/eMBpEeae8cajKw5A35b0OWf6sp7k7Vv
1FdEfLqXydtc7Kh2+qGzsHmm28cE6mMUbPobCAEOagiNAtfw4N13R2XZFNMOMI7j
4oFz/i+404ZrsqmQW91jT6xige9G3pbJd+EJt/MMyrM9dP0iS9wv6Wjj2eabSwWd
cCohP0fxrYy7YfxqOGPi8XZQXVk7l5ypZK/2PAd/eYXdT20gHKDBhmEFNuv6C835
wz7PJl5yHPKQIW49Sv/WqHei9nnEXOpZQeFRtXCDoJP0AJIsrJQwaRoZjF3yibzI
N6Kx/M2JQMhzA9lgoEVaou09R9FPivGrNcgyApJmHYAkJUWxN6L0IddoskUs21Ev
knSG2kmZuWKJdcBzSxm64kyK3AfKvwAkyEXf4/pUg4a16wcfjFlCj3CKGqiIBoSK
7yPzNHxdu7GxBKTlMY9vxkiwlmFLtpsSJq+XVzaBzC2Mn8PoReSfTr4oFFg0DSMs
IpaAf1cUuGodAn7Hj7h6wXct74TMr8c35WYoa4Rtq3CBdRh0RgIrJFzP6fS1g+Il
mGfmlQ5Y6KgFPpkk+cZafp8zGK8I1HD2OTLfhTvaZZsxWb3NiBQdlLBWxgoL/zLg
ADgIPOz+JxyFGVSB567s/y5R/en/Es25cGLvQ1YFvbQ+O8n63YpE0/Yom6Hdcpef
VjJqsUZyP06TNLiZKZKO4NEZLyyn1mEika0QdnlofMCspxxZrdyILrVwXLjRt4Tb
lccUVvJ7CORK5DwDyDKcmCzluPkCIjdxHOvyRIl6ZrBUV9K3wXMO1uxZOZMuEs8W
u5pf6x6k2bLVC1hF/wdgR+UiYvZJHpDiw0dYWqOqy5cQ0KIr2S7Z/w/pQJMfXsRt
GAjfQLjt8uRr39P0GXND4ltWIgZTSsSNak++Wf66+EG5uVsigli19A10V+VApBSV
SofY9zXrJU7JQ9oBMae0u2rLqS5dBMwsm2bRDncJmARxKCxCTvtLGDXpVi4ynAVq
D6gWrQZXqTIMzYSr+ZOAouWaMjP/CHqYETIGsH/AvjQIh5kT0UecwzOI49LXVeKb
bxShd+JOEs1ERSLoqLhkLq6wcxG76OiZCwFt4s/h6hAnw5rnPiALfo+TK0mvjf+j
nZIYmN9CY9b/6TDYyp4PhQsJHxVPZ3uIwPUxlT8Rkq6JPOayQCaAyzIm1aLI6Sl9
9L9GEeZLW7bG7vIP9pMhBv+f2I6C6Q7NWjv2U4YpET0S19lvHwdk5HemycBYl5k0
MksGoiNAvPa8/sxBlWBaq3RP5PUiE4CZOkWfZM3PijxU6sm4ju771aLEW2kyZcGk
Vy6jw537uqDu5JwRTv+NALwdItiCIvd6Z09pMrSATgshMYdjGRjiI1wrO/VvxNHn
0mTvsV7h1zE01fm8Nqaj/eXa+MgyihMHJHqk0F9gguPGpBceJ3aWLNfvCpSr8E7W
BnTccAA/bl3EXF4L/35MhX1ByqE/78vjXKLtSWF7UPLow02uxANcmRJ1rbEO8hl9
6i89Jleus4SXQoTxLhHHRNtfJuSLpG+DpU4wREnijIMmuRP+ffH2Pp8Qi9NuUF+x
hKkT1J0vJ7prjigfQLCgi5ySMLq2lvACMsG+cHsIru6vyFIZOssiLEGDdGpuZB4o
l0MDoLXLtWDOpTZlVuCAenz/U9c2ddXh35nH4QFv6nkKjUd0KyBkDwe0AptDdvNA
dXvPE0UZO2ApDBJNabScBNI7v+PDBa2SZWQekFm3aIx/6OoU2vhnNyaEtaSUqd1k
0vGs+llDpclDIHJdYC0tZiiYxfNZoEkplJ8d0dJ4XxieMYNzJU3+nXpCpTmkEM25
I046nKqEvG02BPH3B+1Tw5m05FgiQh7cKWSL8YlX5MJXIjv6UTACQnqB1RUnxIQA
cYFhdKxv61pWsUtDLx3ear8PFqCzGalA4Vd2buVZ3gRXR6yoyjcVKWB2hKA8Ldjx
f7AUIDvB5w0KG3Ghod1LDtT66yIAn1Pr0iAOchSCfQuE1BtGH1hVq1rZfvdneGVX
haZej6+vY8qd7sBWapF5hzp15KDObP2HLeHTUV7IEJzDBS2NjmC73jK+I5gxNgVV
/bOUkS4HHFqM8sgsKjEsq3Bi0UHq+l3oZWmtW7hSUMjYGndakIr6CWuUouvbXsc6
MCk1RThD3i65hyTEjy9j1ZAIGbUalmVUD5NJo5FaVivfkRnugBtqGo/QdutT+Y0L
ioufBntKbKWvqLIUevPEeoHdHxQ+cqpsPd6EsUIbXpf67cwlYnynOUHsxdCaASQB
MOA4W2lgyf9MWxMYpzEQnyWJo49EGXEbX6BlOtEaxpYXJvIb1a4r9bSWd5IxDbP2
y/DUsCHdqBd8Ow31jfC2herSiPxTIorQTU360sY+3IaOw6Vt4cnrcg2cde4fjT2p
1gT72cbq12197ZAd35uvnnW/7RjhtR/bcvj0jDbs8paaJyzbAw038lRYMTiOpkk5
P29BcBdML0qDcAX9MOSxKc6XQHxtX0iNot5BxSf1yZOJ/9awk5XnYfg6UzUiQPjr
7W9XzCYAcy3JtgVmRt2lV3aIAyPwLDANQnumRukYWt3DcLjXN850drh+u58aSC3s
ZV6nNLKzepXV9FwGAxiwbgv0nzKWVyMkUjJzmoWry2KiHWY7aYpaSIZw+Rmm09b6
lCQhNRGJ6GfV511WiPdmdHZz019YwvEBP3KVXBpUvHj46FXDEbqjizMdeW8y2TsW
G9oF7RU4QVWNRoQX6sIgbFdgBUIS+CbJA2i63H7pBhmL/0GcxQAV3OOHdLG9cjGl
vbBJ0CmoiX4twgPPcOQU5wh3KbKNaXXJapbGPvgtw5vb2mBiYE5utRv6RaoB0f2b
g7/YOq6H+r9VUzejMLEQ+Z+LytvVPzaD7iJninKOKUGr0nUC/yGdZuw3eqpe/VQs
0kw1oeFbXq8XZYimv72aM+SimZaSuazIN5rFiz3IrNcrlIXlAFXqv/8Kuj9F+oUb
e2ow/7yIyghIo52FJvH5XBYsI3/kFziRWTLp2iijGxSCeBdil5SXqf81gQ5sV5P8
aj/YdMwSWGd76471nAD/MHfBnvhje9G3WOf0ypWr5wglVzv9Lrgp2lEFOCsFOaN0
LKmScoA1c9Bkkz/en9lbOuSp+YfCpXV/JjKb11HxHBp8noqe9vrFD0J1ZG2mb07w
YO7sP1h1SB752HQHkdXtlWPB7k5Ba4aC8SrPIyB59+8vtSy+se0vY0LU7Uy5gAxL
BJO5fq7vF64c82BZtnv+F3p4pHMVI4xGAyRFPjSRm0kmNB0mXqbochNbNmf+yEuL
DBQjNDuVKrhIQ/OKw1sAKhfSuG4RYpgEdH4mDta/O2T57+xXbH2AL4B2P+VILfLs
X928WqzG81QKwjrIPqebE1C4doXkcF2OXSGd9/E3o9x4ST2LaJd3UYkDvtcLKs3U
bZFgi91LSl6SftnB4btypFjbw7K8yZymtSk7xeq7tk4c8QelZ+d4t96IB1u3AzId
zNUVV81suZ5i3AGajlLRKqWAoKzvHUZLkdR9GdmOoVh/6+cSM6j7dkubkH1bjbTg
OW9Sfi4S1YtYoVqMsw4BzfPUTZbr2frzlmJv5SJHKWti0MyzqUupgXdrBwx8qImY
Wn/BR2r7JjoSiHIpNcpYhjCnobtfZJOXHNAn4ftTyFKBhQyaL+eNa89Eyi9EvcB/
TFvGE1AQZ5mDTB1WTn+Eg452ewtI3RBQGVqIBiclEFUm9S088Vbwz/1T7ZEe12W+
HsMISYLNxH+CKmkQtKfJvC9zUZev3SiEi0e80F9dSv0g94D9NbVF1tf2xrkYhCDk
Dkj5m0uNhAGKeSncKU1AEduLV9MA+hqHN38kzblrylxMuNeefhpbzVxDdhtMgC5a
Q8JEo2YcBIg6ghK2J2JMJtwRTuX8YcS+tbjjaxERbtHkE9oGHaakEtuK/MdWcvc3
PsMjgJF4+ARxh0mwo0r1yhcpFXfUAqBB+5KLqqPSYsgTHkZxtjiz1l5xn9JyiJof
blE1wSPO6H1XtLuWucD2S97LOfhD1eMYHFbtzYYvfpmvS8vD3KOQj8RRrjyThTJ/
gDZD2Lm44jjkOKceQS2lId3rlG5ZDQo/dI1rPVot8p25jKEIynbXg7r13kBigfu6
un6Wyz/1CuCqUT5KUrWGjHkwhzfJxsMXw0Q6Ws3QxBD0VPsdkn5ooXdu7xTc0Dz8
9cukWY2t+EQns3zqLkVDqgjtKcfz5YbTJ4CELcTznuX4mQMHYOmaO//Oc0LqcjVc
2oX40lAflrv9DUjsPb171KqhLI+0GZTwCisZx4tOaJqAZSsRhoS+n9NytF18+zz6
3y7o58Ii98nOjyK1o0fXYtNjPJeB+thj3aqiWIoDNKRT5dl+KUj9nHx3xohDN666
wcft0CdF6Qv31OZIuf73V1X+SyZd0i4pUYVOjs2N16G+h//Wp290+FZdHX8y6vIj
wMwWUbAxKa9RVVMGys0XCSfWPTJjb2dTCbeSWnMA54jSog4hg+zC1zOMzNDoHsHZ
LVsYt0lVZrUHJfbckUOZsZlI8AWr47tNurchE04sfeC8Ty4f1v05Qfet2tr4GfV1
muIXZbQA5L5ol9PnL4abiP3l3pv4uLTKVxNJuRwRAcpp5Lp8FlDkjApVr+HNfmuc
+McHvuSTuWvIgylBCI6NdA7KRqRSXu2zsIh7It4uWZOrQldXGXrvvYF7DMUPwOWP
x9TsEcZBdftc2HlOAJLxFjHYCx7Ax0hFMGUrYCSt/PlHFx6KeiqIuOF9Qy9F9NV9
N4idclcGeBgIdcky8N4/cz1j4CGR3rVynvVoIQR3D4vTyiFgprkc0CBXjSvlssta
4bA0VNdDCWLvYFY+JHSLIadJgFIzmSmGuVIQuzunW9RwVCyyQIs6HyeH6ZxKg16u
Cot8CcOKoPxTUcV1chU9UKMwGR1kOzKX5JtEpxiq/BQHTsIqdiHoDFKLAiUlGAIu
5X/UtzRAZtzvqebcQ5U31UBOOWl0O5WzhRDdy/vngFUFzZm1Pi6QeHKk3DPKaI3E
qSLDQec6WVWDn6P7tklPR9Y9qiCsqwN5OEtIScf5Pm9CNuDgqTGXcO90Z1o2n/wq
6Q3ftAlx9MbmIcDIQNr/S+Py7idMtjVRsIOqkeO8pzH6QkevQ9hIw/O0ds9AP2F2
2X8rJVs8ct6AdHQj8aegLmo264kh+B89NkJHZjYVKCHdS7pDWtpJycJSUwx3xniy
Y4adTK2iKA17F7Pma+oZfxrOiPEsqxWmNOmUDb0Bh1S9+/R3kXls3l+cfnDzNJma
xkR095PkcFDsWPDw/1WfaQVdgVIdFaRZpkUr7AQip1OuXc+g+s4FcMWcmb+S50j0
wD+pB5c/1p5rDltzkyFLdEzKN8nuEDvNKK8+k8GmUlJnW9RRbILMEc9PU7ZYELE3
7AES0kiMK8utl5Ibx3DQ6dIZe10tPeZ2UnubHQUdMibUbKWbViU43KM7CdEBBpTO
no6HTlGagUUmMYWQWKchPEU6kqk4VuxWbyymAVW8i6wOsRhIDyBgJkbwfF/QdwPh
DD3fcKp2iWrubHmrMYIjFJY5ogBYvTNUC4lcE9JP6/T+/0IZcZT/bGNca1lyMQ6M
GfIEgy7byxqovFrMCx1RcJFpvGt69lD9f8UzQajEkxTIiNNbZ2e+5ILfSQ3xRA5K
GtpKArASc0yK8lKRUbwYjfbm1cyxDxhSfFcCZmARWLKVLbvTLd5cRjcbr+p+VveZ
wzVJqrqikrzjYKdzLnnH4YOIcAfhzerhduzLoT0XZlwg01GC+rotUzKMkHjqZAFR
3GnegJVECL9pBNIt4JlleQTQ7+N/RBFHuzVgzKpvEo1X7h1PkqAx/mtnaxPBfMyu
8/ZtbBsCo7hks7lAIvAdPvRekOgtf7kH4VCNzOTdsQYue/vLUx5pR3+Un8JrGnsz
BuqhvhgpEy1ESlO6+HovAeQNggtEw90GDjWpYvFc6cG9Kv53xz99q1hnn+gk2vGc
sSufA94lwZd5JLBh07y+sHFUm1PqgFIsrMRwFx0rw1PM2A9LLhtiPS3RjksUdLGR
plplO4ERkUG3EUWbZ0xdCKK106Z7KEpiVMNYi+tqX2wJYLKyyjJV8QlHWOQhyESr
F9ArT/L5LWA9dqHLq9wKFd+NcofE0wjc/uAvPj4/L1vk0xCPGHXMkRvmPmsup9LP
OiSEMkBN9frrpJ7iA8IL4+YMzmfpKCSog61aKTsLcpf2cVw1WHigUjWMXlt/5ELf
9OY/VCkIV0qBqngoEnfuQkn3kQGzicKqfI/TW2W3jfyyYiZ4uWap2xQy40jluTwj
dQnqDqmifrBn+ehkK1HO3AUCU6JujyktBrp4P/RO0yZeCTauZDr3tAmY5kZdWVpV
5CtYuy1f2zPDl2uGznV+IB/PNTnLIMWLcay1j6JXD1Kdl9KNafeiKz7ZcYO1B81l
aavVhzwpyQXO98QaBCnZSLEst/8nAMyvuOJL/9mEo1lZN/IiGvrKTjkbjEJ2hHBF
TwMy2VAjvyClwa5+nFiNpIr2ior1arpA5ROVHlJvFuG6Z5mVNZK1YXw4cgwzDSMg
PAc83xbNg5duU72WEVeP47efHZzgzzBqABcgxOV4vzc0C+cEdxrR0oVXZL4HwxA0
fDSyLLAKskaNfHKpAaB2sIY2V2os2DZ/K/euKM4SVKuXS7aoIc8BeH9gKkNLtMZn
VWsifidedVn3xTtFo3AuXVEpw7I2SCB/tjQO9ld8D6DOE6dRYg1k2lseJNX85noF
ExhrAUS3d3n4qXqU21GQhv3BclGrl1UrqQMOGZPmmdB7EI9ChHxel1xCTBcmVoPe
WcXoiP6OPAH0MMxeEfKKoBCPhr5yHGO4DsmxIwcRcw2fRZFX49PUEhancY2X/sA2
VY8S69gXUU2MRdmCwdcyqnkJyW59/Gy2P046L/LAGQL0j8j1159vyBl/m0vYydE7
5E9rTACnczIYIw9cUCvNuIbTulxDYhEIjw7vWJ/vmUrfZtDqk4VJnX6/2IKvcXqB
4QzzOHQa/1VRk+5OmWTqliQ5ha01Hhl8uk3BICCHfb/1RxU76M1kAE4OaAmMPq2a
WmX5CiXWuuwkLKIrKWXPJF2Fs7XV2z7gB9oTTbcul3PVAlhzIfoEV6dL10RZrlPQ
vl9/UHGmtaqgdbLtSoebnJOZbLymUiha/bBh3eO1TXGAYI8bQMiIsIz8Ds1qqZHR
l5XiwEiHiivv9vBvL4OO0lIZ7+qD6UQe2+Bb1FRFrmSTJPu5AmWg9alQmamVtYKx
3ptIUgXHfRSGUtVhRczWV6shhVmwYuEHNitsJjtfeoa+heg8sqQBgBwxXvgOziW+
mXTUgjGj5yjzQVo4MktjayXUYfW5jf/+sJclCnOG1ek55zzd9s/hyyAld7PGWcSL
inIwwu52lOhAx/QP5nSswMhUUWXDqWCHpDnNdv9jAd18WfMYXYfWnG74eKn79PbG
9aKuA0Xoq8yjP+V2o8aCxhtK0/ZmX6VvixS5XK+NbQP03JExSdQHBTCKSfNYT/bj
GjjnphNFFO+7flEU0O8UCiB3klVKVo9X6uCjfW8mGfSng/FOxyyhLRtfBhKL9MTQ
nQ0GqPC5wJcn8c83TBQU/Rm0/8OdGu/zKNiMbYYlOseo9dtduy7Aolp4aEhZVnW1
7RNMuE2z8GGSwj5htilM4ukxrbBDHMm7alBi5MKxHyzyBTGOMUrlIrpPQQcPiIDc
7+SWhhHjZRa9RTWpJF+R8hj2A+1b2wAdMjGCTW9O8HHxE1cKVMk7eJslJDvQJQ45
mJxMvxoKC8DNrCoE28lrCseCuVPbx1bcHffTz2/jpuJ0s/imGVQxfU9aS1coeaNv
zw4Yqc9uqDFFz9aKj1vclZ53HNMsQBX1QVfJgGLVLe0VDJ7agxmCl7mjniGg1ehu
8LHwut4DnWV+sepm3wWy9EZQ8cIGOXZ/fULz8zK8IA1wIVze8c22huBcBJN5jZZJ
cF07ouYlGx/fjgEoIm17BdGDyedQUPSjQlnoUqzLGQXygtZUsRPevFciux8SEG5q
A4NMZaDDj2e6zRixr/APTiiwkwTzuElOyKRKukdQKi+4Y5Nyn9Bfud1KruB/7byG
qHeEyfOP6PDvZyoKtCBRLF0J6E9u5B9oUGvLmVxmF66X3NupS99u4TDrInF/JuaY
bAarvEqTzxazKrkc1DfooQVwdxq8p5sNAQmfEDmsS+21vrT5ZRAN9BHWhTv5UmVU
mvnanZK2NNAntChbqHbCZkOltMvlhDyGsylywQOthSrm1mRmgpmASQYT/evmgwlb
XcxPybzBGeptjScNBD82j6bLcOOMkMNuWr+s3+MmzlTVKDepG4KZqJtiQHDxHClO
u+dO3Di+vY0e7BpPVXQxyCDaVX2yws73lbt6mb8U4Buz2KtVjYXOQTDbQng78/TD
8EIUGQjBr3CVB8LeAxRzvvR4DVU0KDEMAMabE4iqWoRKc2GzPPePXOVZgM/1nw7Q
wuZsFOvsyBdGfEbdJ8IeoS6HIAGUbi0SEu6m++DwCFq3Z0AaX0z9PkfOq+Wn2NMH
tsFlyJXrWWSq/IZmZi6GqDulx8H8+RscKxR8zEHYuwpRiL+uX2AoHu97yQueykgG
sB5yQXSxbkYSupVi5Z27pRPLjmj0I+9C4PsOlDW07MTzN3HuegflixPPUd8S1cKq
YSQtwpKLc+huftf9fUPxf3m8JOXrgN4w+IyDVOzOYirwm5/FRuN7oPODdMjcyZvf
5IkD3EUq/JdFqMo6b0R3Lf4OGjO4USH/XQ+S08naDVSVUl/Ci8cI39NQFjHfMrMm
8T9TniM/YIQL6bliZX+KTX7q1rfwweYwyjvimPWKrNGmkG/oU896ZKHSyc8C0+Or
vSdwF0adYzQLfh66Ioqr3x8w86qW2rrnVlVafUtkLtOw9p3+W57UQi/KEvBemnu0
9xiq+r51TZtD1FlIK5TPFG9BQBqfzoNma5fCNF8a1EJ1Q+4o04sl0xiTQIJjRClJ
cEz45h5/7t5wXMaW2Yl3gA9pYYx+Nmirj5AP9KFm94gUv/piLIR7lepkCpvPghne
FrHzkYKdabkjNTS/0hm/sHbZTsyIJ+eK5hhtOptSD/odXg2WkivxBTgUc1WsuXVB
2epjKR6NrNOmWzHRCacirQKp+gVRnM3kjYF9k3r0WgHvZisUM/jSgRpcrGU6lMOz
Lb7JoVQ+r6/CNrDroBkbGDCXp1gVVqVVumutz3Sj1HTr0swYBzfhQk5d0LhbaqZq
WsQh/hHvOAyv9mtb1OQ8UqE3+1CYIToyHci75hJ1wX9qpyIgBlMqINb7m0xZRi3Q
rcHv85gMTQlwZiLsG95th/fsUb8xtKIogyo42AZRibUMO9N8hY5P+fKC2PhQ2mR6
QPcpsh6yTMPluh/WSouGYMlrbIANHnAtPwoBGjqlEpN/EMkFnXAFqcpWpUis4Gdy
ryOfHrBEs9clRt6TzJZXR5IE7OaVgqybqcRXCP+LRdthmPdN0NLU6du8UGWql4bI
kPxZQHsjspQBJpQQQBfTKAXp5oISpG9VuX0xi9orFm07CLucwgkhVswMjuFpTkb6
JoC0ZZlgTCbgVv1yMe1C4SiMvfplK2CGVm3Y32bFOu1htAVOJUJ7UcI4o0bgBZ3o
pg0dpsPZV1wTHfiEAaiKDBB981IF3fnUvqsxR5KVqISU59bv+GZE6wrpfLE45Eps
QfqMpzB5u0n8yF47d7L/bWmbRLAnkZ++kfvhpTKKDpVuGP7MftoFreeBloAeZM2b
VgL5GO3Z2IEQabUMx1i6wTYi1Jd4cieHu/7ToDC0cArSW1oFwH4Mb/2kMfc9W3WC
RXypss4DfKpfmBn95islzjpJPlKnHE3za/6SQLlVfP1mk42aa7vsLf/aLtgWat33
SWwhI7VzCUTXf//6Fq6XJ2RGENGFus/weemDgz2Kg7UaIb9+Fld6IQwVOstxusPa
pUiUdtKhGfDSGlaTbuZudRwmbb3EbANIH9a3jS2CKvEUM4+Yaw43SAGMBVGlBAew
c1pjHNqVRGGKDLOWun6pqOdDcHgIk3BUBmhzfVBfvd2YMW5rEMDSP3sYWO6Yowv3
85DuEg/aqbYPmCxxosA7LFDzgVHtkXpBTub1jjKreDiW7hEbBnMOyOywmWm7AlIr
+8lPngCuOS7Wokd4Nwit910plmEB9c/RXsbgwlLHhwXBber6jwbLjx0ZI8QaO49r
+Hm/oX8QBOjpXbsjrqkzVvXO2W1eiChsBC5Y8k5WZxkPVk4zyhHKdaZF+lP7A3rI
n82m7/0BiLp0Okox0xGz9RmaOuATMLD8JkzBbCO48XI/UdZZigPVDOm3wc2Vsk1u
eNijSIph7qvVwTfDPq6b+gHX+oKIKsG29YRTUxfDuaTZXdqyUAX5G3CyVsy8B10C
JU+0rjwzt2/G4mw2qadv0eyZPxPUSY2pSbSFZrxKioFRU2lJATF+mwgkcbbmQig/
s6T3QE93/oEviMVelN6brHG2m7p8KUjEsXBNMYKz4x8PHaaz6Zdv0Cj0HX1/e3+f
oOtJZIZ0hH4yjmeujvq/asxBLVQMiypZ0fgGkoH4QMkFIhGPO4y77M6Qx1zMPNEJ
nWzVftJr78nX0wpGLz8MtDANomeaZig5GTxJWIcKApPwdaOctkqaiezPvJ7iAD5X
7QGP62nPaQXGWHKGsmLET8WrMCzy6JadiSemJ/FbCzd0rfoPTBjBlCNI0Pyc9ucD
vWqVatB+U0y0Sdz1m93JtbcoSJCf7DTZMgBNDT0aVsTiItPbiovjN5UR7V5VY2MO
oHcp22BZoiiMBDOzAl4XSszP9Ohjq7RIUQsQSwXnkBAITjuJmY44QOrqsblRJYXA
bRIzncEcJkp5+1N3/ktqMSNV4u8EFaBCvmKRtSUqEwgLBzlMexYbJtdo0Wc+dr6p
4qdBQC58m7Esir1GHQQ3UZARQJrC4ngOFcYlZpzECz7UDPpl2zzJ7EZuLghGAsGz
lQsUSdWp3RhiFi0/ruVW8o5BO8LKasZU+di29LHVi+1fbfd60zrYaHJR+1nFO/dl
NvPJbZ1Vx6XVFdJIbmbUSRq3SeUHvDLm9wpZ0b40tmSkbgUzcFcvnk2cibhZ7CX8
tqGJWcBX4mocPoB4Mg6hPOvKwiZa2hyMH3Lzq+wLSqleJSlR1z9IFvHo2kz3J9Zz
+TbIehU/dCRqxRBgdnfUF9QJCNW0F8aiUG/pbmLaLbPBgQyWgxZh7+WE89k4LM+l
wjy3ePDpuZOySRGdVGGxzWJsTBR8aV6TOOG+BzSmcVrQ7NTSiYzHROlVAGGYp0C8
7mJbnX1xrti32y6oeJTCZxSeUZg3G5VLjCrPuwHARoVfrBPsoDCkTy7dDgRD7uHZ
6BymSbPvcKuvzH3p9Hp3pXfmDjxwjtYUA4m13wtcnCuO7XvAzPLvwKW1avtScAMD
00G/AuWSdMl+Q0wERJfFuIvc23fYUzQlkFg0raPoQ+y6UOT4cTMfapLK2jmiCi89
0ugR8jm9D5L86scoUA4TxJyQlGlHmwPi8j3lJMYx72lxgTDjVOPR7ZZ4JtiBr16b
pON07ymVHnBvBEX7ZzY1zlrinmCx/61jx3TmO4mXMA8IMxd/RQC4755cDaJ74a83
sMpbUpcqn/JxKs9fbVShoYFXHXg39ada85kYejUEhbLh8jhk70S9DUCjlDavwoiz
rvv40KEojoazanX80FBBSiRmXZnNa8cFYtyQ0bBbzENqZsXXlv/rDwCcxJaOhAzJ
e187S8xavlQdsVsu+eZ+BcD0CvhvyzBO5QsThp7dzLTeXKrLdpOYEiBtKU8WrIh6
JjPJm3otefYS8NW7l/zn45Lmz1gE6mT2zwfDcldBl3aFuk8BxEQ7EGP7JAHeFVj+
L6uEj4tVO8NuL7pjLQid4UF4aJ8T6Cf+qvuYn7j8L4JRVWvUQWKaiLV8xusdIb44
YofvBn2w+dQPS/5GS9oFRI+P2uDK+DX5ekSqDU4i3n50Wg5m4HeRLHVnYTZf4q3/
WhCLg9tItpH09OckExHme0dik6W8ACYz/6M+9uVKziUYgNDXXBwnIIVeNjH/+mTS
DIQE3mjZs/mfyDnfYL1+vuHRIq4kbc9mHlPTl2am1KeuB6SjlhlP1kd45n+w/xWR
gy/+xF81O7xCT69EvdKR6u0DAA0CyduqY4sIyguOWOKSwN5FbhTTWIozDEXEyvbj
z0TVDqpuXW3C42nalEixAGH6sCu9+lY8+qL7QxdqUlZGy+RZzbXdCNKZVyjH8adD
SG6AUaMf4PjpEKSRQGGOX1VgZor8PtnFQ+hH4dr9i01BQn976/WrFaPQybJfZDCB
ZVjEf0XFMobSDD5Vpp/INtwP0d6GP0Vdk+aGCnYRJEZC0xYFkVrdiKc0yeQ2WPQi
ir1Q48AcnfgZ7YCkwkFmVFBQ0mSaGV7mxGlwVK6DhKzGgCB7VEWH8jUlo9LAX69S
/kR/9WnEmeapF4rZZJLF2iPvhfFUviN1ja92A8+rvjwPnPji39vDZ/3L/a+AX4UU
ZYfdhdxQgMOCAGYREzisUdEgiz6jTFrFzWUnouj2Em1M5qTQEYQLdd3LRTTFvLyd
PgWnS1bknI7HgEyjODNBGhGh4Ayp/io9dQrUT9TR5ymlUCeY/iI63G8HhpDu6JzW
frBIi8XUGqaTXDVEbsS+S7ZGqk0AZwyUNjHI/x5mWOkiesGXva9cI6NH/8Yya0B0
BkB794MQXKHbbAZxjajNS5ARI7FbBxI8Gx6r8w8gAmsur+V6xmD5ehvmT18YKFRY
iNPk+6LfFzDrcoFPuqF9yPeFCWgd8CgFwVOLaiPXCc5wYVZhKoy3cxvMvBqMuJyk
8SWuk2q3x5vH1eNBT4AKnC8nZMNUFdnOfXZ1LADeJW9R5blb3lqoKlmE0U5XyL/e
G/ME9myBrGyQgWQ7eidCGt7gS4d8YGAFC38oUDseC1G0wZtw/cxgV23JYoSZsB8O
0QLjYudmOpOJgV+ZnJw2iAYJPfq832w3WHTTP5Em7PejkXo9eVEb1oiroosxHnJ+
0jubIwAfNp0gsgPu9UTbyVD0npVnbegMzp9LUJApRD6TUNl1eokdww4qSA77XcOy
xZrm55Oj7l+3Y87wfpXTLUj3kKOMJNyw46nFoF3IDHIdKNx6nnfLOQlMKDOm5y0/
X5H2ps7uVlmdGnJebKh0/zrkOsAQHrlb2s+I8bOsWwao/Ifd9sGOjdPu9JhSB9kw
+ixCiAIJ+VJualTu9EZXhHGAwwE5yRyvOfX6V0m3M61e1c9+YTJahIRlmVz+vjUn
XPc8Pi0f8RP+65SYn/mHH0jxsQBot8HGOiQupoW+EpZMSo/sHUfAgHtsfQP6HGwm
z/uUDEPI1ZP2mTPeOez9OxR56ET2GTU51CB7p7HdDND/0DpBDc1xoYfszmT3c0Ey
sYt5V8Y+0wt5LEqscMjJ53G2C/gtmRqEeUv2hIRG7p+O6CGdCE05uHIrRRaU6fPn
CzyQMHJFFKXiz0bQZiugWMaZ8Umg5T4d61vwdDK8qshWn33PjH1QHdKyplkmwnjL
yDQZXUMOfccyzK5RrAZY8J7SY+4WSoWbn+C0kEEhx+W7Q2dw9StPa82Zijf6qnki
6IOeZPMbWQ3H5x7gRpLFWsejwIPSyamX0hh+e80xPPzvc+ltYMDIlOi2TOomb/yo
gv6Bk+W1Rx3/viyH2aaQS27QsHduK6xlxsYqnIg6XkxxeU+K4NNzmdVifeOGKpqJ
i4humnVWSgqcGsSNDiBxrPFGM2kjspNvAHgLEReieax0t+5+mEtW1RYtFZMtFtoe
0xzOmJxyx5JLw5isNXWQWDMnYO0+F9AcyVjn77qo0lP99Huq2OnCY5VNSv4rOfku
jCKCZTEDhvv9ruLlw9/i4NObv9rGCXogQbqN1CI/dhOXHQJrK3ltQik89kfWOVL/
syXnjmn9Y7MGjk7+Wn5i7DMvR3+A2AAN9stfgie7pXu2u7OIwJr6bUz5g279GTJm
m6LLIJzzg7n/MTa+NJEVrWzDyLo7QNG74ly9l1CWA+FN6hxhTK9Q27QIXN4r8wiX
lRb9jeBPxPpuW3yGMaJZpr4s4Ta/EUSM/jZLp91gjxTm+B+god4gYVHwuQoSh856
5EBMc64RZSK3DoFBZW1hELH/6rg16C5AxtS7tgQtDe+8h0pKB8hD8eo3RHrQIQa9
Z7r3Zq/d8vQcKtWzb3dQZuoYdJMaCLLEQOxhi+u9ubK4muYddelRr+/U492emdhb
WKBRj0qPuPl5nArrthEEpQvE2e2NygBQmVQicEFqa+WoJgHDKI76jdYbHC3NvNHq
otlBwLQmte4JdfyURPnhboXq3SS4W/oDGSpHWVPdSboSnmMpOxfYY6vzSPt/WlVG
IC8ibIuL7kPaEal4SKi2wF7LedVW0LXOOXmo3EAPMeJA/LN27NvsVZA/cJbnFfjy
stnWc6pLlR9cq5PZx3Svlnv3eLVV/wcoGFbRjeNBf43090NTf6mFH4bXDrbo8IBV
bJHvUZrUfowbil0vPU6TJbrEO4pqO+OLpD4rch4TucomXFkIwvdTxz7rjKAmNo4x
zfhNTuCRH3sthRNwQZOm5s/vzvhfA0ldNSFPp8D7OT3dgiJ1KSIWVgSL7Pq5osu7
2n01TgDDmkEmudK8VvNhClP/XiX8N7eZfe3i0dbK6lGA/TLq8EABVUc967DMse/n
ad5IsEji+gsRXOVCtNXdZ7TQXt7S2i3VpiMw3Jo89u/xMNPRUNDb5mVyFsvSR4wZ
JwdvFn3ssL7rtL0okzdjCQCzeZX1DtXHzBCAScp86l32cUEuM4VNxPoLG+TXOlzz
mGmekm7ZHOPjKkl7A+1FHh7yX2ODGd311EGxLTU1yUIvIvioxX39/WN0JJvnezPi
tN9zq1EfEvGX4aUxBtmMRZQSW7SjH7/KrCG5a++gExXb8ve/vdvhul1kXY+crf2b
hp3FTm/JMZ4K23gwwabwv/wDoVzy+p+ic+u0Qh47hsNQVOBrxAvlERATC4vOx5Xx
q0UiCG+tPm20RBgJjqU0xPr0S+3kggb5IyRTEfrBtSQ7Xxqu4u/slkHC4TNPGRsi
SBRGatz2GfeSbNGBoSEsE1HLJE9GcGwK1aFwqndMrppoSCH6ar9Ncz6o+TCMoiaP
+f7QEP5pB9tum5xt6FwoceuKPLF/3bzI/t13yB/7pwFS+RWChDUFUQBt86JnXdZZ
oBKEU/k/x7tkCQ8tdeSklVj6EhT3HMuKxOWkbBxrDzaPQpsl93ng+GDDqwwfPLeV
v7+krst3AEZZArsnbrop76BAQC+NwZWN8PFd+vcL/5xU8LdBx3BilNb0JlIMXmGp
05Cwtz71khllWgoHcH8DWP61waAMBExIdtbkkack1AflYHBogLdoE1TDxB85Gx9A
1VKz2paTdZVEGC2nC7tglr1AK78giEx0LqP4ZeYl/NSx4dHQp2UNjh082kl5XhJm
yHRYm9i8vUSlyjUB8ppfUgelpxoioLmtrvz8qZFeAL4/L7iTIIPX98CK/JBw0LCS
PJOAQh3392GQ6VRDQn1/g29yzGl9NaksBBtiol7O5M3ApEeW9sZu8gJq13aF21Ro
miV5QMEPCYUX0YPKtB0ZGKqTYTx4HL0LpmEki6MWN9Ji+EwCZTz12hmUfqwooe2K
w4lCppg0pV9yX7mCrG+5qsyFXNrimjglAzQnOPr/rIo2IUOopwBaEH3NUZVF5IJT
jzZJNZqxmUEhgYLkJ7M/wnWrJU4ATbyU+mjYfb0w669k0NeDO6HodmOoVm1EFlTI
RHT3QQ+a5aq/z3yOmrSKLutK8si/Uz6+waAzmiBWTsoWTPnSoUl2vdBUjb+Ne66O
TbTX1t22BOc3Ve9qZ8Way7BOZiN2boPlIQ/Stf0PbLXROjjGqRaJXhtbYT2SlIKo
uEbn1f9C8KzunsH/aaWe7zeDQLKaYBhk+QebqCm09SmwWTKyNsffSgDa4Mg9RkxU
tQUH1fWMXbsid3CnOzSM6YWtFt7w1j22eIMR/pOpwFVeeEqkEq9IIZk+QGwgjOAM
skANapdjRmw5e5LOGaQmkY/Z3eE2U/7cl56+7lwHpZsCaav9YVpscZDwbDVKoKQ8
3vMQX/szvnkPK8eshCs5TJlWchGClUYWP0lU/WZK0oMzpBeFe5MlLa8V0FN+r2dh
a5GYid+dFRZBTaY9MZio8w5Hf+RuoPLa6wvWFYXBZSrnUYq3s4XmK8LIZY1RiyPj
ugLNLC1UPPkoVfN47gnrd9Kgjaqstyd0COp1KhLSv7RIXW30YnbrYIYkHxwt3YkW
TNdo9BU1fQKTxWfVRsJrLr3BBX1jwjVT16jj6G3TMo4+xhBV6xK4R41IljM6mAki
8tVkHz4aA5MMl+YT3nTBUpVaPGOiG8z8hArDxgntI9m6pgjLiSbii+OGHpK6gdkm
d0KVcr7YoLlbjPc+WRpxB8R+36bK1S69/bSFRJaiSFpdX6VcGZdnqeGa7E6ayvXe
ERGTU7wddxS2zydJN7LjBQqc2dynwe/Oes5UUIikJH0FYYNqXleUYewgPPC7qIud
bwqq8Njey/s/ukjRJz/rYtUnmzPr/0OG5k7idggZ0aX+dCXDTTtHf+bn2sKOqZ/N
7sDLBjDCvlc+HovhelBh6uvFgp9MoBiHwAACzYI9mKGGF+WqrT0zDRpG7EGbmr15
ivKHbAKdi0/Pwmd+9E3jCEVhmlZJYHUolH4GCLXsvuIogXzwOhVaeqHGgNHOrBW2
gsiICp2H+6O+2XWBCjZZRWa6Cux9gzE6ERA6jGRj5AtF9AszgD6rCy7hZjmjMjtn
wn9rnrM3oABezKAkbhu+9O1LwkfR88so64e3fEGPro45SPgvL0VnBGzRg6UcYf0C
CEWZA7Tmhv+2I0J7v7+vq0w1cQgUtl7wmOY4rr9aJ1tfBC3UZe2vtlzMwtT1rPEk
yqHxmzkF9lBpnBu4WuD/jArB2EeiLJ9d/zIIJzgYSvmjY7ZKVg2xa49vaFfJ/YGD
ydIoLo0f+7/UWyA3xyHdlYnkMwfbAcZ+/cqy3oRfdJT6eA12Li5hRdPVx2aQKZqF
tiAPUjHNgHnwwZkh8w1EVk6Q1LPmO9dn0mAV3jyZR8WkxncwR6Bf6SEKTTI3EH1K
6/aQxM3BYN1AgViBWj6qZo/+DHhQdQSeqCPRHBK4YyQEKwyJ3GZjKOe+TSLZ73lZ
lDlLTlT9l5v2SLllc3pfY3gSjv55nC0UBApGo4U7VvqTdHHeq5xFumN7YHLRHGNp
EtPUQEFMdfQzBjDb0cl7HnjZwU2JGaBklUi58DPmgKXSAVzcI5ctPXEKVevjApfu
FGEcNZ3YdRO7Syjznrp47XLI45+vXuCX/zYADHBSx/giTjIRrNdq0QQbtumJ534k
gnwzm55WJD3ZN2Z43UFKU/HC13h1lJeXEX03zlx1xLaXhTe97K7Ez6PZxZ427qiB
GgXpgd5qfPyjlq2iWiT2RiNAqc8N3KPvW64zsreqSrLXT+prnfz8+dNh2m3RA1XA
IPMLktep+mrUswC+DZQppzzgPv+fMMOYd4vlikJVmMcXeK8AcGpckSMm5ltnlr5f
6viKALoPx1L2GlbT4/2Kduwfo9IcGLSwX7Zu/2htIyV9zTZ//ilKoe4u20iYyz8c
AfOCj9oYrdYRzbBvuuBQCkViPJt/AGoftTzLMAwT2TLOZNky+s9t7W62RM5di/Fc
c20551Msuz58PtbgGJGhYU+Dq4hA0AVLZnr9EOliXFMKlVscsyI5QH0CGPtxysqq
oQ+fzZdcUrmSCDnYU2Pa3hbCH4CckMzcmCaLaAilHUZhOuaw1kLelOmz6C3W81SU
ljbuykt9VTnvkjY/1BvlEDjsCpvFLVsk4kDxc/laxW6S6w1fdY5qrZbuhnnRirhf
z5tHaYN8nMYRm7TgQu8WUFiJ1j8OZb1ZQNwJkfsEr23nBjksAuVI/lKiaZhM79Sf
gZECYolsdjeNdwWiljWO2/+0xVxDaz3YZXncD74pOaCvDghiHrZUEB3PtCuQPe7/
dQiLOVIXY+ZnccMXOX8bsJfoQvQu4dT8qD+ObX22zA3+N/S/wiF0QACkaBbPd90a
kHNleP5GMQS0zzzusrR/4UJe58h4N2tS49DaswPrzkaqG7/kY1r7zp+jpNjHmStA
Y+m0qjxG3kShftRmi9fRZQbDrv+H0MDZuYGmG/4LJRsmtstlG+6ZE0248Xgq+GLA
krpI8N30sCd9pwHilmu93w61Ylx9HgmZbIHcykbChRfhvzDG8PMt/iUQmN2vdcln
owSrB7vWU8OZF3r12PlgaxGITrj1XISJI46LbdfGBgasSpOLFjixAcoA5+niZwSo
sgk2gqtJK1OJXRI/Sy2TcrxN+Z89jAbDk7aj8PKR95xJiwLfpd4OeFnz9hV8esC+
7CyfmJ4O/2UzD9e4QcRBwmHuMyiLIAO6TgvkHRFKd96h1zCtr+iKK2H8oWh74I/o
x2qNKZDSHyFhtKEVczVMdAa82fnw9gHIq7ExkvM6X6VWFAA2iUlT+gWQsR48dl9C
s7gPkrhocv18kBtISlvCPayreWgMIvGFqZcLb1JHN2RNAeNoTVCmor5vHiM2kS7F
r3FpNVfzVOT/mJtI817rfy4VkA6B9gWeiVGJJ41UUR9SfjD2/YVYZpC/Ts9TbJuK
Dmg9mowJuCFhpNkrySNM+KRjqu610h42dSDKTb+YSCNYXeAoHWX+zZjAR89DVhqm
RHaGD5zQut95QnWYVpZbM4r752oKtiL0uP55bGtx+bP16PpEcUrnJWFU23egWWds
50ukAwp4+oamMIj4SLXQJ2h++4mfN8hz6m9hiBUfPY6T1a5ZxMXJMNIODLH4dh9m
7RpwkHCRqYMndAQWqzfcNyJvJaOS9L6pB00XRXUVOMYQXRFgCd4v+kI97zRn7JgJ
vmT+tT77IoUCkl8nfh6stFG4lE/3ILSGF1RcAXhP1XwpLQQrMZ9zepwwIiGgnzXi
Vo1w4HytEt7i3+o78OXJ37juEliYTdozX5p7JXIShcbGHDn1xfM078vnXdXT8Peo
gccL4+ln69Rvd6perRaC57tr3xU0kpdgp9wY6QDEAYwmpWs5wnvZ2RCyYHyqedHy
IEgXAJ7gq2kV/nRDG/8N0I1mTj2/3C9YlxrRnfMw2kkJIxdtvwkzvGC2Gi/34lSi
EtveORynz9Tm4/gVyPWYLjDrgpEj6E1etoiSBOkSX/7RMWLJNAhlwIuyqKoN0iDZ
xuE/b/Wx/iJnoi1WcA+NtI87Bo1BIOPcoyZ4kYfkFHbWCMIcuK7w7bi0IkJEdDeu
sfWnecDrTZNUkU/3oKy19wEMkbKXSSMGxFyDA0eI1Bn/V3tJdFvqTStIKp9Ruz4N
AMfo8rzuyb7ZUCqwwvt6APiR97YzNXQaRlytF7sZIuxQdFd7UPJ2WK8lOpewYWg4
4g7a/Jt4mxAQPfYeh2i+8RFms/VpL8q0SjzJrhtjynigWPi4qck7K2s0C5KMOu/5
yBMMNltTvqyNymcPoXR4qnTilwOpgEFPwJJZegGHP3ZoX7k7IfjbLGWkjkLeNire
SxUmJffMW0ts8yy5UHKi8GDfwr5NAiHo2p+2jC6zJkocZzFtakIehYUBUZwGUl4e
537NM4r35KqPSyrcTYLCxakahoBELH5ylkoF5qrHR3IoBzJkBFp8Py0ms7QTltrA
s5SXb1FhPoTZbC/aISyi9UjD2PoILReRfu5PKT61ysFV1L4p0kzaa51GfFAeqYTo
RaRt2o0rTIfUN9Wq0mq/SDFEiQtNu4edhSQEFpGC2RqDUCndLPQK2OaIaNw9SFbk
DuaUbD3VIRUBnNmibfQ9g31vlI/V94p8OJYlkOkxu6S0bamTFrNs7PUDJ43wEv1p
8Da934C5eiImVcktPjJlxdQPXel9JVzprneoQdPLevoC1aZitt1rImtGGhAdYV35
tFmMQpZ4txEyloZIq9lETugnvZ0rtDilDWZOem25kAZLzJEjCUp63ir0nU5SSsdm
f91mZ1guusDi9HyKT7/XHJdNv6CVblZdx4+p9uI6me/QPJxO1gqI2uNfIJc/d+Y9
qvseuAe/UGCOWBd72gfUTrLW+aA0L6GYznyRld1Yh/6/UDEs42WqzSWrcTtRJZ2w
i7WT8M6IXA9HPbRP9au67QlZzQZXTBBrtJFwAG1iVd6hfEMwbdsy1+kgWag2obfG
GtVQC+fPbIqdgH/KBl9e+Temnv36bONVshzokln+GRX+HwHzI+Liq3Qy9QI8HNp7
H1OEJqMqqrP/s5VWUdGJIDt6ZynA4eewk0h8/5Mk/zBzGHehd38dJSfp9nG3NlL3
+DSAyhTg0Aze0kb+B4Qx533yLW14A9B+35oQHnTGW8/VsbGBMlC9UYQQkEsB4Yi7
T/ehyA/lDtED3m8uMY2lYx9u2gLnMy+rLf3oPS4FOeN8cLsWmra3NV/B/PRXNHZr
d0/d/WAVaFjK0qmTQDpyoaIo84Mj1v3KEQD370uQTEiMolqhI+BMVcf9oebgi1W0
h4Yik7yZHCFjpglwV0mndO1W9aMw/V7/mxKle87RQOf0mVwt0o6tsbL6FZOqFHWO
M5ozmUkrxWq2zxVE2xHoFVrn40Q1Sxq0ct7A64writhdvXI2+etbOsv5dmNLSmb3
fACkFveSBw0gll+vRogK93SIQ5RLrCis3flFT6ln/4ZDMHGTraoAq17QHfvjFRMl
gscC8N4ltTXJZ8keYQkw1DDcspTm5CunZ4zVir9lIGhFhOTjinXNSSemQn5KD3qY
GAp4eXyvJO/+WT2bLnCNt59/AC4TL2lChPEj5edOX9k7iM9qdSpzo117jnW6PMy2
GwBprTNBPOdt50EhjfHBJpy7JVWjIku9c6/A/RIrPYcXGjhsbWFZwXfbWQReLhYp
A0vKDdyGeMhWulCTClQm77oDaGiv9Z3XDS7G2Z4J+XKBSlJFJQiFZrGbehh6LzZp
GabcSEQpb4IR+BXj9gqM1iU3ivyhmjxfeg5ZVcyRY/BykFtOcpTtWQ0mVFs/iGLW
ycx6dR7MqelTFe/o1FD4fzJRetI9dmD2bE0N1APfap5QaZex3bLGiNxA+ZEyfr/x
/1in+bwC6nACjPd0pzuER64oathQ/VzLctNSRVBxcoqvdBiMy9tHmSb8YQgUZCrv
GbsABq0NPaczK6uHQO0JIscHm/zWGC5FvdZqacAxbDkQ7/bJl0CfFOfFKzvmGMjc
KfAUrstbRmg3FC0Zz1UR+wcsaGmoMsUOoYhqrBVQqgZQnOrbDxXrKOzakuoRP2wc
sHTqI89mj3fHV+8CdIRX8/bk54xTjvuEqBW1UA14X9evRLXGrMEVqaRiK5FDLNzS
CDpdhxV6hLulgC41T0djYqFyhhddpLH1hI8w4o3CCpsBX3HmAHUhj+9gQ5Ik6Hrx
JbmJiui5lDW9KQybWtanSZmTnwtR3l5HCAXTFjxtKopy/orHFU6PUsyvvibyhcVK
ww9sVi3u6rMXwxqgIn5qDnpoemNFxNVjlAyn9u/mEwI2SuS+Ku2HF8FC8LkYTq47
Mo63ii2uQPeZQnFIwtkN4NbFxsHt5fDQzBtBzoMPBT1609uQFpdWMChoge8jxIr/
sNk/mnS23InC5NDflChmdSGwB8nUefUoRMfDBar7NMeN9cTeI80R4tjCZiFK8w1i
uDHJd8UvE1WtBQ4HY31/bxhpMw42YU++ZiU+n/hdYMmhB7kOM51tB2mqcHOdWshn
U2FwvPmqF1q2Aw+PQe9pq1R8rMsRadOwYfE5U1+n2Jj+3q1jLiwlNC9D+b6mZf9L
BIfkZ2N8HszvXI/x4TIy+g1cWAOuPenF8gcQWK7JWdZrbK2QUmmrsm4I1RR5oWsh
PzW5M/Y01IrJX5eVLq0FfVr/OVPQv8Lkj3kGKRlmaGM3DC5CCEYGL0DLF4zgUlJJ
vNUm9+evCbOclqvjIegmSOp39GJe3EFAJroCA0w9ZEFrnTkX12N18pychKtV4/9/
ych5hTW8LMmoIGa+ASIh2A7a/N5/FlpE8W8Pxl4Vy8DNbBrpOePj0vul1zMbSul/
CX2+9k+DvyJvyBbqRYqFW2FpdAectgxIFYUofN+c21tuemYMiUVTmHkglpZR4aD8
T+9RIdG2wX18lPI7Lasu26e3MS6j5PXHNcuvN0esYoVgDUVLvuBt3UDoLjeeoXzG
N+fySJS22BnqOhsdOT3lSk+Qg4xCjZjEWS8dk5dv/lrMbRoErExNLlRGSXTYE7Wo
8hNb1q2zEBU3/GPrGuB7tR4YzFEC833XesfR4d6V6haX6fbDPgSxDCOJxKF4VhEU
h7sWMJ/2JJwbJo7iGj9/y3Wbb1Jib1BL2uHkif+hijwpRr1gw4uwTFVidiZggiBU
8v23YDT1xeLmg/UMBsxEBr/jcH11tF67fNvkKTGbEbs0G2Owdbk3Pza4ilFC83SJ
OmKESiyMIYu/AvKA4rxVolEpB3dYi4QF+HlQwzkUWqjERDOiAQcTlO0+jr/6B8Wb
OkK9aigU63aLv2HLxdQSGvTT83JFFb+vY6lWq9BE2dUDLhPcx+BUvGY6by+zx0g5
8FnGQvlE8NqU37j1fK2mLGMxenDG1q2u7PG5tnfNNnN2idZFIIpN1d0fPHUKQiMB
7geD4Xi9d7/RkNLwNkldLECDoVZT90G1vIhNLfiTq0FESDJicQW0be8QAo4O9vWI
bJ9tEaWTI/jou0EiB04ZcQm5P8rlgX36FatgfmzJY2hdM0a5ErXpm7P1LqulX9vS
TDfD7AfHPaj92YOa3rCs6grUJshoC9kbepyMQ83s1FPJ6UhC9p3lH7HufnfCT1j9
1QwkHYA8v5CoikFfeDbAqEMCFXiCEKWgOkCE8te6dGfcQ7+uYZkXsWkh3l/uzQkK
zVLC7PXqUe1vPW4srimjVfBcI80BYE/8yCnJZSrT/QfoEEoWSOdaFXxhQeFlbKLJ
ZeML6RbTJImoimqWWt52Q9RHQB7HVpzwkXf/YISEPtq1sgDmmYuK6ctyDwkQNhVt
B1PPCN7faMcLCGafI2BNKugKkYL+t8xoHpvc/Gij+FRO3x3F/86C3/fWh/h7svcl
zeSo3Y5w3Tu8RSEH9kWt45T6yNpeyaPtSuZAuG9unMOaFGdcPT/4EIhQXjckcSzP
AsD9UhP2vTS+cyHJVnchZ+MRTKcJpSAzB9YNDllVTtjvN6ltJKzB8doXg4H5Ljcj
zrixp1ZzOnR4lLyk5J23KzMqA7tPLrxiWoha/dJQYINY800Q8f6cnCJxp1pezxeY
dXZcTU/INSNgHkLRQE2NJqs5+6ckxyhKsEfbPja01JQqT8rGlubuv+4oGe1maIh+
+K42TII5xXaIRcy+5RVesBDM6I3Swbe4PAtyaHRon/8//ZScWOxZCChHDyRpx5b5
Ut5wOluGzIVsB5Vu40XrC+rKEFEnRx30WIOzTTMRW1tLX7/n49zaV2wQ5WWmArmo
piJKdFLYcd3QY6xq1h+se0wjdfDO99g/YXff+kdI5hocKnDE8CafsO5KQr3ahBPq
qkSX1San6hBk9hKhuAV+fN9L2saie6WGUXfG7cF8zdYNzeSsIMTL0QYjSXvnAtnA
/QTNIp7L0NhFNFqel1IiKjFtMVYghkhE9BlXYjZO0l9KkocuxvQnBTst1ajhFUtN
/bIFuUzuPpoGg4CSTD2hm+hu1yJJZCS60aTOBtrIF6U/4xtV//Gsx+Ryb0B6bWq9
39sDWyyb5cU6RC9xar0f2ZuGFp0iavLm39nEm52n3ciojStGcRN7pEvv36VzdIYX
GKxiJYA30hp6yq/g4T3L4mdn4UIII7lR8KQn4QYGAYaSBmrv6PJZzvFeUQGl0SZK
K2XhgVVL4ulr6TWFjwyioUqbKMkWoe/lrvxjLU2UEx/NwhCJ3VAiMWgibcpaXJF5
EfE+QRCYva/hzdiqPhNGDnIIfj1wu/x707sjvegIXR5KL4HAy41ou72SgWz4WIIf
gnasisf32BCN1RVQlZhY96dSoZJSxCEZdaYlQ3QZNIzMKF2fID765xt/8WNzeFC9
nyuq1W+j5TNYYqpq4wRpGjnXQU+C2f5lr0wBKE0n32CWPxOUY270elhVddWn3c2r
5UlIVDOwc0BUAW1r5t63H2R1lajKiDMsrN7WBX5VEHRJOzWm1VIkydmN7AGvWemV
Yx4EP+eoriin3PgCOVLBORx5ZUTNTYrKEiwS9vLWryoOnF22viXDZfAHsPUca/b/
cz9D0YfTuCy8kqhFoUWSDccoUF4lfnxns1cSSbTJp/FAyP1Vk/6AW/cD/sRx2+uK
6r8GR1J77ZE2St6RDGoW7oHUKLh4RF02RqdTIhEI2fTVav2USxe3dJFLCBcPI1sk
7m1UYbZVA50D+HzJWVQbkOLQlf5ItlH3rS6xqJlp5nBN4mGXA0yNKX6gyWZCQSO9
AIpziIB4912L2yPPxUcL9pCISxgofq9gIuyUSAE1UnnYnKDfxBL83yLPTP3V1rRx
UkFHf7DoA5prElhwLRoBkmXEsyaaPehjCvB227Qjq0Ce1Hj/OKFeaGCb9Yr9DMPZ
rMjYSavaG/mDOvFsXnuqaIZV4qJSqxr97yJ42OlItrKP12yVf8oMKKhlMrxCiGTh
yUVLdkUoAdUxCtWZJhpZyYQXBAxRS6L//CN3RUASY1NYJlHpMrigBeBgWHDld4K/
QymZ5PbDbAkxA0wsMoOxXBVndpzjYN3OZocl/XLLItO9dXulQ2i1zLz72bZbF+HI
OHbvzoN/9zgDm4ERThiZkpLRnhZ9mSH1wUVZzWkLFiGCZkjViaaijGfnJhIeabaq
xUGXhtRQhxSngjDcZV7yHiMfuNqCkVmba0+rFdpozoZ1YkOlzYcEfHDsTFMpauSM
cc7b4d4jW3gqk5W5zZPjOTCRO29DjcQiUpgz1IQSzsp8AMWo5Oa42HAOQHekUK2r
6Rb07cXogxFTAG0W4IynFwyoLkdH7V26vp+zd3ujnV0cqVv331QKSU9lzzVqre8B
K8QNnfqy6xQUFcCZD+1rGw++JB4qSRicwhHJIbdrAjrDiBete0GI8sNyol/YhqkU
3OKFoBbC+mwsDzLOj37cqWXrb5TpkbMSEfzH1XHvURc5Z1D4mXEVjMvynEMWMeqh
DL/rTWbw5qxaqZh46SQ5BUNnR/afKjZ3LQC+XFfVkNDMixbhS5Y5fIQhaY+88Ik7
d8wU47HC/MfwXzpI89mVuk+ErhHFBh0mzkH8bQmgP0JFjMl+JKBbOhgltduJMmc/
AtfY+SMJ/tCBQJ04vr9pO3Lft9HWlRy/STcfFiyI++r3ZQmkzSN1Rv4AuliY9OK1
9olPGsukzU1EIRJIL92UGmHIuuQih9dhQCHO3i/QMLH09tyh2qM34HloC1lcpMqs
fIzn8OcMIVv+gmnSNFN2ow6fA2spCXZt1zu0EwI0CumDBsv/9YKRFx/JSrRGeLUC
+j7kHDSzZrBJgQp+10hdtteQmb3wgHM3oq06O82OgjwndEj3/mYxubbJg1RgkgBW
2fjIxHc6M8JaEU0W2CRA81Ts2Q1oGKFrF3rZhw5Zg4atcsK7Vfc/jbVYNAb4o3D/
d8/j3UNoUS/RUDXPyWr6E2UJc9nTXToQUFTNjpFeSsmxnjXW3Gkv/5M03FlZekVx
uSWNTouukGjmnoCK+uyZSSu95z5busuVHt3le5c31oVsvqQTp1GLc/NZL/yzpzPf
vMW8yp+KFpcN+SPt50GmKiHi4XMwoH7QeWRVzA+yzV7l72GNvN62ApsRsMjcTQNb
Oeoz5r1ottp+puQ3LTA+o5++jmjL5cf6mVlQf1ecT+COIM2tr1DlJpbluogTtW8P
qD71lFBNdXdrsca92goUodbuTDJp3k9fCk0VudwHFhzTzskjfhPIDKbsJPyrYrqz
njjJ08lxnJVB3Y5gdD/j+E4kht2qZO+YtyqATrumcZveWdzTfFSRwGGdFk76Fckv
iksiTU5Z7HHHhLf2F0kMviG3ttXm3okekU8hV5Hhl+j14NZgk9mowvLKnsusHqvA
FlXhmKnlyDS+7OjgYWwZwA/tuSrQsZIL60ZGT30nesnpCOaLZDLvC/jIU3JqGN/A
lOrtIVGVW3tdYq2tMq6geLx/Tors3WUc/wVp+r2b2Km2E1+b3RqzbRtICVqJkHUp
bhLxaoV9SHTAenpWJR/7ndrEDm0Rf21q5ui8DTDdIKjWOyVckryBoKYnjAGiIYnP
86j+MjsWRZ430xQ7slDJeYmSntdS9LX8gJrPLQBr1F+cmyPOpmS6nFloELnY+nbE
DVW5+9I+OmvpsM5ruMN9vE91YQdO55vfrqgjdbe+mBIU2AYDF7QBLhQ9pUlEYFA6
lL3gAyXk1B/FBRYUVWx8fg/MAy9NJRX/W2cJ1AUDCrG6q/58IdSSXPOT3jXoGayu
8CKxjVQK4MG50KMxwNmunvsVFHpaWom22QM3RyueuNRA+FK0I0t03b2GSxapAIGU
jxd1iuBGsISWp5Jw9D01Up3t6i1oZJAiSyr32Srf7J8vtKZf+C+jBuHreNOMTvyn
y/pBRvt86T8S2YjR8CG96KFODx0Ra4UR+3/lu+0s8wYwkdrPv+uSiMBwWe45v+cj
AY5kKyuymTazjsu+vRotZXL2wBe8L2PcsuRy/r5ffHd0GVHEMSYV5HloTYwSG2nH
Cus802KgdTLQJnu1ugYSArEy646F674cIgfVDbUGN2G3jt1nbjIdt7qjaBieqM15
Gs7OSMqCy1a9D8GTiajdSINmv6qEJJDsLA7DJnwEEBo2ugXqbiFB0HVdAOEW4GAH
DiHsjoSVhO9/dMyQwBwY88/WUCikTZIdy/I/Is+fPaQpTcRXJWVLYyZ+EZ+AUO8/
v+gblpapdL7izi1P+BExaVup+XVxJmPhmRqopuRx3qGwUpVTazRQH4IW3K8hPV6R
FithNkmGMR9DeEMYy9q+oUDeC0C20UbQlSbD73ERqSUyhYGboDR75doWCViFWWK7
ZsEEFm51iIg3BbSfJvtfkF2NEz3knFVd4kFgsum+0f6E3PKBmvNDFN254gLtV4Fh
hLXmUzWvkyoHANDnatyo0WmOYjW5fsYx4/arWbgH7Q76N/N0H9JCvTBnIqs9lyPc
IWgGluifMOcACSwj7azHuQadHjHajvbJOb9tXj8uElOgmrSVJlRVahV+ArUp4Ity
P1t0h6LwEwVXb+f66prEVD2mR4nsnIDEQqAYCTe6zxqPUIv8/rSaOBvFgNhJvgmO
SeaSuLrYn5l7/9CxwvWtQmfw1Hh7RU0FtJq2OgGMN8/XHaF3qVzzkMhZcL/C1NID
fZJPGFTLt3Nf/mCzSJhMbr8UpZg+PlNzJODfroj97Z1epEzdLXfbjB00EvebhMzU
8NA2Z+Ijgh24vP2061/h7OWgWDusHjwzrehSF3Dk/44lYP0mecMuBKjVvjdHizdk
5lUTSANFLmp10s0HVijV+g8H/cL+i0M9YGqDP2GOjNloGoH948rGxlCmSyworaH9
oMwDlV3RrVyR1jIlj19KOQNdffibIff3VR0gIogI/Js4q9IOmzuyT93tVwpf465A
Kga3FpM435eOs/fclstb184xx7P9Q+/7UOxWeMJFqVdt4Ly0Z2/fn4zLAs/dsnHi
0FaOKYG+MiOG+CRpavsGuLSQ8bwCTbrF5gZDIRg8MhajKGG8JnoQ39WjTgTlELCU
7Lso5O20YxpnCjn470AhrztFiYZX6JvR/VjV/KOIT3blqbbyU1jdXUiJQDvEEDR/
4BPO0P+la3OqQ2OjmpKGV3+D9UvT4x+1hp6lApWdXoEAZ8EeZGDsyccWCNCRB+pJ
YegN6npFrlNqHRAdWE2ygWKrzeoFomoLArPreD5Yz4+jenMiIwfDWdu+vhVoP+sM
6cQHeUPgnYE4us/3NI6kqgoqEscnHayCx8HQI8ps5sTwp9Af1cn4YcDU3DgYlzhh
oDwffkjA4ooHBMz0FeFl5++cNOZIcwxKJheotcy7+RFVA0YlnOpF5+KYYWNS8CvN
R3G8MgDvcSYiPNt4MJgwfIPm6Fb9hM6HemffMerMm0dbGg1p9EP7jCVXd1fMM7/F
RiPTud1BwuSu9zWXUrYJbXGxphMSHUDonCMAPkhR0qEy6UxGwvf2bEQyuqjBdt11
pyISf7NP6Z4bL6w7NASQW1U6sB1DpNaV2rGMizyE3O8Ri4pkEQCBDJLPDIm6YEqt
J5nnJ6/HRP6zSUkiR/NTUZoBlHUSjl+Aw8YN999gIqambA7dyTdp1H4j7AJeUz+V
xcfoS6MrdDbiUyMPbAbdDqSNXSkgFR/ozdKsx5CXT/LU+lcci39C8mLAJl0+Ip06
9q/4nmskqFs54EZbgTVY/Zpbc4QmxUdHQQj7Dhu6G7vVx5/Au+bhNvnOeKuFoIhp
6olJBXn7TaTdk+RLG5vu9zfjjNybSfsnmYFkyAD5vDHp1fPJyNUYz2sKs/4G8BLf
/RZnRceP8FY+boF2kKovr9y367KFYyIrDOjJLxBG9fEjD/mIrtVOcONPulGcZXvu
6ZtgtZYgUwbO/qhTdKbJoWSYTXBYskknxuL8pikYPZ8Ox2ChwtNlk+v+jsQ6pXhN
F9QUEzKFieTHeJfOdpAGiQ3w7lA2F0vSYfI+zGA9O+/XITl3uv1natxMoN2Vd3kj
7sYqTxhHpeWuOU33i5+DrlcSYKurO6KPHlzvNKHsK5vWY/81eDOS32B4f0VlTRJY
44WeXf1c3TEj+MQaN5agLpn0RlegekAB10vq7SSihyYJyIr8l3A8NdcbdF3CM/wm
wzbesUZCt7SEVZ0GAraUimyKyon7ZzLeSTPksRSnum4Qa3hXzsbShAldznHdSM/g
RxOE3ZEQDnIJC9ETUmvl9tpFghG5C5/Ah/inFGdSHyWRGA7O52Fo9JOcLTyyu9bS
D9qgd3LSvShdfw7Y0q3nIjxmU4HDoKElnw59ba4WONpRKHGtv4NDENGUgxYOZGDU
ox55FBuJw5l3op4IEksAF2Nim33tw5b68JTq+usAgYcf5v7MohLCYW4QRQjx59YF
eR5G/7WW5hNYLYRGai9ABp03oNRHeuqw+Jk9Y4c/jNxUTs9iPdpMx9CvVwLLInEU
ILos/RVqQnbcpUsxfPQnuVVxKwikvA4gLgsughWx7UzSnKSbI7RIVIee/GK6VeGs
jD4h9Yt7FONrYrVUk3RrGjV/0+zQRbwiQOmbHZ/SORRH9LNdqNyIwk8M1qDL1JFT
C1PFihrlxCtoS1LQ72q6gFabxCs34txoeXE7TAlepJH8U74zGkifm3TbPdfrNaab
pvK6nS3LoOcFs2hhJHkgTs0imhC7y+JPk2TkcsLOWPWwe2IInVfbZRK0y9gz2z4z
EEz8BlMXZrrERlSOL/dYctZDGPRMVz0M9MAvQoSEPwImKsz5norJt719UtBQ+zE1
oyH3qiainFrqK7a3pwGBruktL9ApdnS5GHfp5Le4nzv6R44c1Z0m/ioHepUiyZoC
mUKK7uw0qIMGEV7mYGtJ9Oom/qiUap29lgch82F8scaljRQlU4Q3qx/poTaJy+XS
aAzUvVMjt2sqso6yeGjOUe4aRP5a5OKXJTNHvBt5NsCtm5AV79xYf2g13dzMERqw
he1dcDnv46iMbGWc8cGKkNJ+e5chl+ZSYV328jmld8plYB85P+WF/7ePJPyLSP7/
PTtHugh8Iwwj6V+9lH8Is0fG8Toes6ZvUy2FIrAUGXk0NykXG/N/xw0lofvCaAUl
q46xi4MKlKdMGebp/FLG0m/FFMOey1nLzgCp7mQGZaFlFoQSz/EiGHJVxH208ngc
4h5HJs6L2gvbXz55/epFOWTkgV5TLSdbpNSvU1jWoGjX8eEFjQNR5sKaG+aDBQIl
Xq89uzefF+VZ4GI8I4vZjSgyahkZA8MT6Lfpi9NSg7HQt5kqHfyfPAxj3RDp36ba
uZOqZQWf0J/5w5HP97p6M9GB/7nhV2jp2G5F05eKfx6eBGrw6U/SB6z1VA1+9Oc3
tmVfxi0QSXEMsZyrLOJGUKb3fdBC7AeG6sw1t9L7M5BDUpHWjyOIEh8D4m+9JmGP
eXgyuwvShM4ZTgXF7zD03O+GH9EocJ+8YM94hjzoldVze9/cb9xxyq39h6vRNQ4P
zIYvFA71GjUin2hO0ygyC972Q0YBVejAciByhXougQJbvgXINKJriXMYhfppEmzp
Qy25mFugzLxIoVpTZI4EbapuNTySRVn+RvdKSmCykKU1JcSAHvBfUTso6Y2hBGHn
dgiJSwVcasPw1EL9pn49bKrSBqw1IrUjyiS7ENbB6VOFr969rwgdXwl/iAB6523I
J4vr1zjdAsBxlmFZOkq+wJCMrTU1TySbrREhaqbVemdcW9OOa87rwemTD5O5O6T4
XbtUIZHwV5B/QI1urLDT0ksU+LYaWTo6wK9YHC4zctk5P7O+CLfuAqY+z865Cu23
g4Qk1Eh3urCt/2E5RUJ+aerMf/9WaciiWm4ULiV0keZBqPd+yR2pv7ClcrqgSV+O
UyxQfB5luyPxudvLr5zKuMdX5x3NFAzQME/SnbSkUlvh83d9pKQ+lMV99UyqtVLs
ICa58BbSAtsBTh/3t1uflUOBcBBMb4eZ15A51MtzOUD98eGndPtz3QUPbLK3uThE
QAMNUIZ7K8m4jL0TTRHZs3is7vpiFBCShWDGO45waxTblSbilupkIRGM9Q4GSH04
JU/eTMVTU2CMfF28unFFsCQ7WhcDSqevkSMzqEUM6AkvTYZdZEkMGFfepsHl4EiY
EXao4GXM9Xgy4v/tr8CZQ5qrQLtC9C3vjVVpKQAnsvucLoL5fzO+ZpszYboRaifi
l/EMemDtZ7CYyrz8U96TxbFWBHSeo3s/r4oflUhXFlXG8HNfls0FPr4DSOuYBHnN
MyWShr//e2dpu3RvTZLf6DkWXW7uou9RO19k30tEMjFSmdVLmPVrUpsNklCxBctN
fdXefcQ8Qn33jyDwXDA3W84/gOxM675ESnzcfsl4skbKHmcsLFXAC3Vvwe3nZKUa
mdQkSUCRqzqBs7VoR/wB6VqnWtttECpyvYIbjmsqua5fZ5BcVBK88ff39t2IHD1G
cnkGHk7OosLbjeRy7N6/dLH7/vJrJR0g6BC61+lHJOSOW5WkO4E404Uo10bmw3+6
Scb0bCOEJcuoSLXNDwkLBzWO+GK4iRQu3DuPbwQQL1LNkYNJ7c2w4U1eoY8E2YS0
zBACOouUb/4qjf4GDQmf6/N6vNCWo1EftiPSSqXDpdLLAOrGxGMFBTKdeph+3AIV
L6aLHAcsGUfJpyC5BQAjfHMVbH3zp/X9Y3v0/3PA1pvha61odq1mePgOTYxKivm/
FY61O93O3GOCDuK63A3ntoDtlWv6RT8CZO8W8etT3/S8RT3qtS8T8AWW/po30oTO
I9Yzx+kTMWuWGl4mUntVG77pNOVwWnqzcGxSZRfFaV3IEMTQidN5Gs76C7yjfNln
ptsqX+b8FNY4WQuGu+2yimkYtC+rg//PVT0M7w4e7eVN3t7ZGdCYKkjKw99qGSr6
wYWagL+Es5YUnri0ZXnC0shpIkSlH6ii4OosV7ANUrgeYQLUDk3dkrRO0KvqIwTu
zvzrQ+vdvWuGQIl4IzR+Q/bEZZUkoJRV26fEgvHMLvpAX5fKEoxQLJJFLXIgqb0m
zLKwvawZnlsxMTLA/Gz3NTM6otElLoC4CpHAjfsZFiUwoOMobfiQE0jcXzFN1iZA
UdDsqB7dx99FZdR4JXzMEM602ZNNRpUjFvjL25Ht1I6iRde7YW/x38qyxqOWwd+i
VGbeOtQcy3gfWf+yynLLfDlPOhr/xZQiDsQ1Zp7U2B8d+4qLvEGvZUKQt2ShZ5sc
LQHzeO4e+UCx9b6zgw8UTiHQObOrPumBPzFpKKLZ4lG74Kl0JnIgu5nH5GsPFrES
KRXK+Qtuio6ZFlHvi359MtY7UHoG7bme1TrQmrEYb/2A89BJFS/6I2OU7bV8fldj
NhLuJfu/YyMqLpQVWUyxvPf8TQ3qC0CcewSk4Wx/Cg78mrLPp7us2adH3c4FZ9Eh
i+RuGkzDypUOQ2U3veY0DKSMWJm5Z9DL7w9Pd3a5uNfih38Nc+XLmFDDsk9dHZfO
6q8GjBrbpC5sz6c1q/aOHVMJtredkoi4UV42QGLpih6zY8p2qQs7EOPAMhOphWzF
kM4Ue+X20m0eyShe0nxaiiTlIU9c3h+JXX0ut9dYLuJlv2kxt+NMU8p6RrJewdE1
M8J+agn7eagWUnwtD4wrGp1WoGYocyVJTDSDoZomrTa20/7JJ1/E7xKJFobexz0c
FNFENaPXtV8eK5QzCGLAwILbj0WIOTCKwP2tY1bpygXMcM85wNcO7ojdeWBFbyTY
9ep4RHrAXuI8toy4B/U00x61Q04VYvF2xEGb2+eYd00tQ3K8NS4MSco9ZqKL3eWG
ORYIs0XiA0PBKgH5k5KtFHRaMBPL0gQ/g3CywMcX2+ZsrFfYO9J+X1FT5LeH7W5k
p4hfOi9CRjrF/LD2hjNoBLkkKuFP+hb9XNGWW0zXKzIdqFZq5kzRgm0wVq9R+auE
MpDGJnt2GPoSx3lhyK0RtDEvmytoLGY6M9cMs1dTMc1xl6JlwF8E7KWlYQ1LPG3v
KTmJt85PJL3PrrK5YLXoNjEa1nmirg/R55atQQh3lLwzz2HEVx1c3CnkxKuQEQam
xV5EPl7baF52M82cvbqNMiOilcCph0GQ8qPZtCL5WC6bHtOmkY/Uv1NnjNpHXghi
elPbALis6oYTX1yk1r7pQUkWvW1qIqpxHzyxy/RQnumnOyfpNOxVDMWwW5X74jHt
a5ueS6XW3tyGnt5oagKStM1RFoenFU4K07mxbpehp9KULWZwCkjJHCBmKGrDukdj
kX9wMY9YMdlv7BG6Blu8Figg2foTTPOqKMroHPqkS+D9t5Uj1V6jaB86+2V+kln+
3otWKsnEq1Xn0Uhga2e1Y0CUCreBwWEd683w2fJ8DdDBdn8zopLN2EDwnRzl1b0t
0ln85QW1xu0JuBhok4pL3TynsEbSlHwC0JgzVU3De4JJd+biBwr2j0TQ7Nuaxfln
9OVaIf9YvI1hpLYSneVdwxF2At3VFLk9KQA2FgA3BIOEc+auj04T/XzD85YW2QQK
SMojpgxS4boOZcJ22g6OuKE+6zGckjSipPMyc/zZH/YdANbTX3pIHBwVU0st72XN
jGr0l/1heBKLsNTfQOp4Of6pCMpMsRer1HSrQNYDO1zKGplvrOnom/WCcjXu6mCp
pUHgams0yMFxmpIKXQZE+HF9S+YpM830d6fohEWVStFBGqP0XLEY6AkSCd1zGcQz
hnZw1OIuI+4wk3V8EsO8gZUktW9Tnbq/sw8SIWKNfJMq8Q3UsxsSvYfK5ezIAcNe
w8AFhz8F+5Da1CEKb4yU4LGyMZjmrxnJTAKBfBME5EFPHVfevaxSYX85wUtM1q3E
biuHIxIpBmBWv3ABIJU5Kk2u7uq4E1is3SyJmGIoD6+DKDhg8hOYuHemdhm7zmJV
fhPwMQsHxwN4210mfdR6ZE81qfaDGOkLmdvq8DsF9dJaC9ocurB06jp4HoYaikLX
CgvQSj92uH+xlIBXRyw0NbayuHLVnVaZNA7OnpT+B+PegLbBZaPAuR+T9f+YageJ
J1/XcV2grN9PPXH5CPtSeWBI7pahHAU8iGLtlyLHlZxLjZHTIUKQkHTC2XPJbXD0
FbKoPWvE83mCkc6VdhxrGT8DXrmURirVbAnaNRm5w8NAD2GU3d7ZNckLNOZo63Tj
lDrefqa0gWNtXHjCBXyViGWjZE8JVDlZRBVGtlKdTAyDB6+rOgaorXHtfhb05k5n
anqAsA7CkA2JDlp72um5A7nORMI+xVqTXwaq0TOHNmx2wWZW3GqJXS/WcLUiMRZp
PnfjL+XOyTRiavNaZ2jh+yzw2dch0WkKYFLqctT+RfyX4RioMxbHbgQyONCLpwsC
RaxKjG4k434suWpDg6zfFJFRI96OuUYonPkchYH1tld04IAoQSM4a0O7F6jACE8v
iZagUIjbPewvz9iZTthXBWrB12kya3NTOv5ZfYvZ+SFjUOxhWXWjTTDtxexhzE4c
SccNYtK+6+EBYz656n/LohJvQW7tiSycnGdF0//Zwok1JR70okwo+rPUDlCX2Gbt
8wFB6ygcZLS4MR+fSRdhyNmxUWPGauT30OwQKhkQIcRW64gTqWb6sCJGlhKPG57V
OYwgKoTsFsrTPBcjVAxuYnACE2xOGqDjeVRrs0ZbxExUbms5du5mKw1iL2eTr9Pb
nC0/HSAMaycFEAsJrwkiAAM/FBYIpbcn0uEp7XZfNNlEZmhESz+XPu10mA0KLbWz
IRX4c5lGwab3YPeEyXsC8SpeVW9MZXIXbuDtFI8C9C7OL5Z3cn1NiW5yjzYoGc/I
sbc5feQJk8pRww6btLUG68a89sJ66gtviOwR863KFfQ3IMMbtohlvdQ3zKrBzsCc
K81pHUS+Ok6+fE+pEyx50/R1doEfufKjQnCQzgsnsUH9yS6hgDdohfhVoPTVFzZc
GQooilgbm7Z6EeSfVTrCT51oqwxGzJgpKxuiKZyWrnAIW37K/AVFDZLsLR/9AgGq
q/rEDavoDR1SpagkjA49ZwcWU03y76t4DL4uPbQAqXkDRczUWuwOt7K2dshvsM8L
zkBDac5+pmzEFDNhXi2p5hLamFaqEVWZZsc0/kh7Fz47Va31dypU0+fuTgEXjVdO
/5R3b05HTQsnMnhv0pua2EN2L+WgHJun1FWPWdAEAZLcOJCp8mLhKedNcRh9enWM
6bwr4+Q63UMfAbG4K2bY64uI17NAk/9EsP3r3aGShUBHLC5fG3YtvKeYQmJXbGDv
o9KfDytgXXnCaf0XEtuavsD6jER9IIYUDGHSy6Cp0AeXSOaIe2myCf+0O4/ogpFM
PQ0Vfwkzz0VSVO9Geir7MBQqhtvy2NpqQ0acvbDeE+1elFBYJdvOUqVj657EG6zM
SVzBnAx6xV+kMrYpzFNYjA0VhfIrPYE2Lh7+J3fsepCjCHuNM6nkIRfyrnDyByoH
afDFjEV8FYJc3d3kAmjAj32Yjo2FonXOxIng50ZxX8z9acvUP2xEHG9RQ5Bk6YzW
B1FfuKZUAuJ+sRTYLl1YZqmsQer8taMkXouG/Lyle7SJvC9Ib1K/eUp88aGQp3Kt
ZpmNj7FCfbEo+C/3sUtN3p0dzXkdAVG+PQy+Nj13R5gf/W0Q8sXkWj8pJaARF5pN
+u/Qm1sgJ1AKx1FrIYpYQweBUG8irrrPtqHHEBZxju6dmM+8/lZb6TpaNnoMGcxd
t7/tW89fMR/ObesmgNtSUr5uldgTA6yg4EgxTYLAXsJMxhKTnMNRMryc/YOMan+0
cdOS6KQ6FhwuuAvnSqhB81UGhR57qjddc0zArjks6uEltAsxrMWq6TKDqzAuhbi7
9E5rt0xmlPalmyOGhK6c9XPSU3W3qXxBm8yIVCyNC0h5dRI3lj902sLFevX5Nlnj
+uHofXOzvcWlKcj3+MOo39l/A9TXqmsBduxSejE7thJfWT+7gCp0j/VEpLD7oZlM
ifC4p0Dr3KTEl4kpA1aaElv/DqopPW1JvQbeKsNl3h3dDbyKFCBcqmup5dhnw8as
5nuFviAgei181UcPWeXIJuHuPG9YwXkV4iMX3nQ1ZyRl7QobHFQun/2J+2WejmSs
1d+h4wrDxT4D3/XIZFO6n/a/7hQfI3+U8cbp0u2jrT8IrtJN4MlwJjKxkyRe/INS
EnctMODx/1lTcvNEMhxcoYOon9xcXysizCDulR8Wn7SgmQXm+cNzdnt6+uaCGKtz
IiFpOd8wYiY0VIKWRXET2b9goB56rw/VX78KA3kU46rZnoMfPbyeSQs6HsP6qLWU
u/AfVsvmg9keiMX3BpQ5VHyunXeakbnMZrYiPFYEW66CI0TgkAFb4/Oy42wM0sWT
yxucaBoGHsBSjQ8aP1DXqtizYu4O1q7dIH2ZpTJXXlf4Ul3v5jJI7V8sLc6wUXOT
GrBtWjPgiCRE0822sL42tDdpmIESkPrYR0WYgd/shPgks2HTx8i9xyR8evodwXeR
6b5mpFr/B3jbPppPMEMpxHDX3WMnJTIa1bZqDjCOqrQmlF45+qIYhYvQMhMJ0RYC
VBtuAOa4FX7mMXMTnJw+VkoIMJRJSo0Je3tO1DtVrZWJRE5HWIjhI4DTBCZ0xUi8
VzH1CbNMvS1wfkLsJFK4Y2ssqt2Av79uocgC/kdHgdCFTXF3TRGnHYIiWEBm1uXe
ZIoXY2Xp9u3wccMn6LbAmm/PP9UOwJJZ6exO/OJM7RiiI9JrUU9koAjtgcLQkswU
r+xrEL0xAK5h2F1cKNPdgzSzyAOWq57zyGKeVaQzsb6AW3CXdFhe4CEr3J1zogxi
qGUMMxsp6a2NlIQqPv20iumwY8IyDH0mloiYQkKJZhYOCexmQH+xwBB9D1QNCi4y
BiD6fCJ6l/hRipZ+jPBfMdgXRQR7ESkGu3x7BlKKypAHZ34M7ouY8S2fJiYQBgux
ezPawuJGnH3HtKXIU2ZlIpZJEiwAITUQrxKI/HO+qUe7Is8baDWbqb9Q9EavxNc3
b61Er4SG1AKXLLb6l38YtWdnGCcvimgLWT8v4iK3edmnWPHoh6s7FeyoD2/kQ4+M
a5DJ4AkpatGFL3ieazqtEBHCl5juUKpqOkbmYxYBgYcJDBqo7bD94JbkQVTaFFNQ
3j6KNIm0ke0AqPeJyP23Uhg0GsSf5Mnzcf3AVfPjVxlqHzM3opEOhWey0MSxp8T2
Xak40sl2y/6fr0rjK/cxLcHHrYVG85NtnOXyeUe6eWe4P1bL92YOjUAv2iVb7/jY
QeXNB3wUnNDL78dg4lJK2WODj1osJcEuCyV5JLXGEzyWrkCttI8U3VxpuxWRBF91
k2u6sWMaFTUsNRosjMU/TZajpkYZBgSbfQHDC1MNKDAd0U23+2ya7OpDS9v7I7Fb
uVm441Ty68XQcnvdwo1/UAv8bck1ngQmGReeraeJHNK+oNVJdov+RDCQND6/NpsF
RxuuDS0F6n/EASwvYb9R57hqrXEGWg7Bu7v5ZoO5nbR3Akq+bpi+UBNG6AyMhfay
hqMdBdpJtHTj/xJ56jYPWFCVKYP/rOuD+39azYTZbU2+YuRuM1L1j1JURag3AIVB
CUXT5X78jQD4M3w9QaW0O40fR8ox38ya4CG/X+ogp3a2JTnP0z3KKj5oK/M45yHH
nSu/5wRh9MTrn5mQI0blwWFO18RFqP+SNDk22SDkrVT2gWMJiXsMPHMc1zCPchK/
Z/jOVhBlX3qlhNznZ8P21rlVK3xhWLwcHIin5uWDdgNdo4OEThaL2Xpsx+EvCEhI
AjFcE3u2tr8R1QH26Xclz20WLx/7l3H4ig4NQp3TXGcCx9VBo+ianx5qSXmrnAwZ
IciBFQZpOo513GTCrXNcDTF+ttIlRsmxydpkDPmuHHM2WjXyLEsvjb9aZGDQjCJg
+cMmaO/4eg8yr+Dx3wLY9AkmxafeB22ME1qNL6i0OqI1i5d2XxLmxwARBO1LPbt/
M94JV1N1cdwvj3/AZKtQeg72Am5C+xgJ2IHGmNtuz/jZeuukJ4MST/ZADgLhq47W
NSErkQ/hgNkhJPzJwDEN/u7BH2e0fu9l3t8eKIb45Gv22qfhHOGZi39SwPsh2Z7I
5LeEdc5OIP65lrTsDj+jlcOwvVjiFeBlJZuwupi1CfHZlRhACgrycadSrWQNstWH
1ZbYQQVp4jBVL7DEnGXWij/FHz+gGlySTvjEM/xBnDgbisS8odYaBMkPcIzaLjJA
dU1tMW8nJvS3dVAhQjtX19WemI2u+tgXUP2ZWos+oj2YU3BD739hxYDASLwgDz1C
KeKx1dNMkWrhXRcdvo7k6COKc632pRdIl9Kkfe/NoAlF2q9V4XOWEGTzNtLwV4Mm
ep5vkug+l3AYDz+2OfzBnERXmVm+TL11ZplCLUquEFMeqZ52Y4zXICKdwK7FjZV/
2fTvqhFhmAx+sm27gfC7PHfbk/LCGli8UjLgVhBAVLQk8/eh4/BvvjDGglhVCJmJ
ktdRH33C/On1VmiiOY+3X/7lpnfI/W8tNkaXrxfIDeZvAcd9dHhl8GB3pPwXgtfE
P9PATJKPQr4RXD+w68m5VO9gmKC5xsqZs2WE7Hl5gIhytXLHo/WWQrLFz0JLBWct
ojUQ8od9gTTv3fh6Bw/y/k6bGLE5y+GnLUD3Zt4tJdh9sKM9ow2leZPyIz7WEj3C
RE22WUe6w46A3ShyFV8hTVFWVi+vHTZqoGMvpcqR+uQdVYkrCn9xMS/K1LlF8MOM
bTTYBLJkGvKuuQ6gnY2TLGB6Cy2UFX6Z2V8xl0gB3DaAIhDCqKa48SM4RPM4V+iG
Nhy1FS3sRyqQXi5fVQDVLUTfdfDWPuNotGuYXwuLQx9XcviSDHB9JuJ3v5lCkgh9
rcO+GRFUrmMPYfD6oupRftzmPCIsuXy0vA1AGHPtyJZRWtoxSE5h1aiAx8pD6E9B
/zadevSpsuY4J41Eg/eSipJ1DqI/w9eJpsBxvAJ28j0/0QIoMlnsB8mZ5WiBO3+F
KoezJ4iuU/bmjE6HYZf4X76BW02rk2CctcsuXhg40GngrJc/Cgd/25mEy8kVPwUB
GsxOc4ZAj2BeuKVjevSYSts25DYmXB/ooyj7BB7zFmICSbHfj5ZYXO7ALsbs9HZM
hdsQD3IirFdSG84z+OLqUkD99uzS54TZoJ0tGOub+d7iZmQVtkCtG/56caPQlMsZ
vbEsFhd/CNdLsaiF8wg3/AgMpxvYoMI4L5CW4BDNfu1OoL35c82Y6UyYeTv90P+L
fzvZ+HglDzWvgH0OyaMzsOxOajBoRl+8NGnmAuQQ26LvT6cvV6p9czDlGbKEvjpV
0gi9Pxq/DkGLFzn2RjrXsQYu+v+6h03pEWBpfaof7oPnMFUaCLrRO0UwX9QGCjGX
tfiqCnBL6xcUiJVj3Jrv52LdbkjDPCVVGTPbi7wi4dBrbfNjxFWDsuPOCXzLPp5d
q5EJ5euAfq7sQ7C4zCI6Nu/FHMBwiDL1MU+8QpIpX94mV9+DFwHXWGwoV1FbLVFC
VMzlqYMTceTMQudvPsX7HsN5NUHNUstxqkE9s0j5oOpk8iz5M5NfUC7pGge3Mopl
0q+7DZ10wVQ15OetUIVxUV+R7qkvh82wFD3Ppe28xOLy7AvMvmiZ4CYX21Sgnsk5
tcIMGPg8orrd1PRXL078HmYiDWtvY9DUWIy9Y9NwirF4GMFdoZzIHDHwVCqTLpen
6ZsHOVi0Mn0zSWj0OjvVM0gx31whq2FBu9SY4HZVVjurpXTH9/W0gwR84/gIPx4u
MaF6C1rM25Jc5ha8UTQNd2hgzPGJgG1FSpY/fM7BzyyE6HBsAUMCLWmZ5UivvvC9
+bsTT3g50SV4/PycnHRZPYOmVg16UroKTnV5M3mlTkRYhrv8TbVoFYmd5Kpr4uB6
jptFdiHCtIzzdrbqPBve2D8+k3pH3bgsAyhhyK+sgM9np1cpNB1b8+8lEotW80PW
i0B6MFJGrgA6CzthtSdJJxVLrRdVyIuj758i5clhBv18ISuC+G5q1zgH78a8lhHR
ic/w4iNoMXrDVzwEN3rDRHGtnH3hGQE2NcBjzCdBwuI4cYlgsgTDMls5uOlf3PYr
s3y0zlxZxU+Kyl8dRU2jfTxsfwveXtNF84RCamTt1y5YNvmkJdYmAzqzqOt/HWth
2qfbaUaJru1spqNQURZtu3DwRIZCOkvRLBDXkid58HgAezp5/0iQ41dBevXaw/ZM
xNWAc/Hf13Uce/88bp/p74OLsQup9FJ03BUqVmKofdKnxKlL4QW8ZNYeh948N43Q
12fi3Jy+FSPE7CIvT54SEr57CMBFHvggU55hIYvydqHBftA/EiwzrVwjsZ53/Ycv
N33lVp5O+vwB6T2CnUJ2JhRbLxNaZsROcTwB3WFoOn2Gz+5kvJmRfI96yJKg/3n8
QysUBjzqVJMTzmVc61t9eZdSFJBi/rB71NgzqPO0vDHmWHOfbpgbw3XCbUElYQPD
MbAsPCZ+G9gbBzAioQDoU+sogd9Ugz22TBaTCWQRzO2Ulzexejn3clNlojEv6VEx
/DVcDdjDQz2K+RkPSED7S0mJNY2/JTuIuhM6csq9a8MwC7gY8fYSTk2l9vY4l1H4
FSjg1VFdDTLjRv7i99wts//T2XxfoMVTTKPQs8NxWADN+udKMltW0rucpAT4RkT0
poirv65ORdAH+6+Xv4zHsJiy+6GYsNoiD0fT6aF/nWvpPUlEdkPM80QnwbKD9vmt
VjJ9baY5s1jbXzFRljxHt2TtGh0DYU5+OMgQz07f5APD5WXu9Y9md/9tSAulkmJV
Q3Bjx6IH4XbDCKVhRHmt74SKCV857fwUUOLxKmSI+m4hh1wKTPoguhrK1c+UIzoT
lFjnVnyPzEokwwmZxwinK634LpVYABmKFvLILZQOqG3Md2PpFDmN0dbPnvkFugn4
3yBa3vWgS90xoEGH3jPpMo7V2Gx8iJj9iolf/kGBk88HoiQxW4YHk0zA+XXVUz/a
cIJllZKmokNNRKkwL7HkGGvcfY5iFyL8Zr3+con/Ev6kCT8JVj87Kimndilp/hy4
Zys7kLoaCQTqSTv24fXPkqtIiVhlkuTKiFQkgSkvMTyi6Af4yA3GV8di3DFUf/3R
eHVda5qGxfkmTyfK2XES/Q9lu7egOHlyOzkkiqUCMfhwQonLIS6CZErHeQRv1auQ
+WLAE84EdydKWkwzf2cBwpNUqZ3KcXkzEaaU3EJxlC2wjOiEWJmuWPaXapHC9/Zc
zsG/NEFmclpGDnOWsO5D9v/El7kE4VN8kwl9zsI9kvUV6ghj6HXapi90i2KyIE+z
hPAgwatbPLafBxJjxnmgIpjLZPMAL/kVrx+FaWH8Og+5sfvGRGC7EO+jU+XOMMLI
LjzKNxTa1O208Pp2Ra1c3WTo6meU8HkchvcUTpfqJ5M0b5V1NfqcTqEpiFKRnl7k
vRqqeWTaeTquZFgig/ZohX5TM7dTLlC/CsK2etgIc8ZDKatOT3FO2z0oaT5GOzpa
g5NffazrC+A+hR/K1Dw8IMpqSM/+ygy7R2Km79TGv6sd/xqWGRSQLXi8Zwwb9VjJ
ZA0tLJ7f9p6iV9vCNnKTOtq1ZJawP6//xU4k7kpdKXfXn0VbdzCMnDtWViyA9jjD
vNDLsYgO+aEyqh4jJ/L0f45MwTbBYhUJd0kej0sTkLL2VPCKv3pD2l/niy1UK2bf
L06pvC5UmafZk+uZyqClvZW+iYFRAbHiQ9X3/9SNw1Yrs0vxaCmYsFMBSYxX+9l2
djJ9r+WMHDFr26iDlncXz2AgaG9FNVFKvpF7n7n34x95IYsX3/IoA/9wL1wUmKkx
m/7hPErmPxt4YCOca6H4AZlNXEVQipJSdt8b9RKS5D8Z5B3mzAwF2Lfnd4jjI3NB
0P7ya8+5v/o2p53yOsxFDCTWEqtN2x9IeRXdw0xm5hefNXGCS0fwCnhJPNFPyp6Y
IdGDoaCaMNEFR06VliQT62fgO45ScrUBoLexhZdTddnaIlBHWbeCuWuXTTzLwmMu
FDub4zEIxZYOyZo4DnxDr53d0WFcZp0lZDAO3hbt3kOPRL+iHLgkpL/L/kdqp/iM
Yi8QFQpyO0OuNaGhgNvHvK8gUxkfXS7lKQRpP9CcAGUIHK74avgXeQJhaWwEH0wI
t71CR8tHND314fLgN4tzjxE3OYusW4CRRiHddt+wkH/6s7k1RMQURFy65lMjnU/S
h6ZoJIosfZlcnHz09EdbOn5bPC9OAcM1RCgfaI9kxUFYEeQpVlVNaGAJHDOHiewR
EHraHHMvn28zjxwWDP3Rc1AJQchoL6lDkTq6YcWrAtWNjETxtGml+l4X2zdt5Np4
POLXoAOLhbKQIpKgWYecKodtVOZmJa4uy5NZ72njEG76h7m7rXep37K/xvNKKt69
q9miEdziFkdDDJhG3YxoYOJFPGzMqT4up2YNE26IYw9l4OPlpdCArv1jlzP/kirS
V2PpB7QJ91dcLUK1J3+NgNnBqsBoa0rmHzhoMt7oNbOWLG5RuKeWUPhanqeXj/G2
FL+arwrG6z0vd/VEunCi/2+A1yhrQIslIHCrsPD54w1SQHJQZKy9xo3yQPCfHu7i
4/UW+cuSL9VQwRRPasbX3dQZflzSWKpL2ReQKi1rDZoaHnlVoCSXegdGN8iN8Vnz
jmnOeDHyqBYtfk/r6xqju9dqyV9jsKYvAhMmTMtYBUkrt3U8leqWvyu1gQfhtDwr
3Kbs4q8B6exzRDyn2pXQ3Mcegs4lWBa3btQVrjxWWPLG1GOKQ+dQFhVu6hwTQL7E
EdDF5DpfHP8c0k1qVjXKarCpiWIn1mqQqtepzOwBZ9H4uPSSo3cyyy6IJjL481+U
v+YQE5G5OaSbdeR6SIvF4j7QeFKSYippLDAH//P8uQqOKkUk41+RLlBEROLUkTf3
IRTOQXl3/oMZstJjp5V6hpRQ/my0SgNpbmvEVeA4ay+llIOFn0LA7nOB03yRcmS5
GHSA9EYmjQ/PrQIxgwSR4cMcVcbDouIEF9XtUYWSc7CdGUG4hnE+/s4xImh1wT53
nupooYnyLgZAw7ywvibeKePh4iCpwNuhmjI7C1IipEZj/l0rMaXA612syy3vNF2I
O8TKDlCZyy8l+zfUMbZCmGzYu1KOZF3TCZ3Xr9f4JnxmY7gdgC2OBWjB6GhmOzWd
CeMDWfOFdR4xS4U05NE3RFjhV2OXtYhExpPVFiMjVU2devYofiHG/uBTPbiA5W08
ll4E+mJMWwqxGru4R/VRNtOdgrkcFvn5eMJ4GuNiMgDZXKrTibPGGCRUvRiMxZxT
P3Z1n8aFDxxDR8AguVq+xJ94vGOT8kUU0+G1JC+GuZ1YwuIy7PBa0fSVcUVgeeJy
VrPe2HV9CnlmbA0O9AKgdWteEDIbT1Gb1DF3fjuZddwebemfNFQH+57WeQFeBM4/
XhI79aX2pdjOmXNP3DIMiLZ+lv8ScSFn62Csccqm1eGQKjsPVFCBsiywsq/NMtZH
Ahn+bzBZwnJtV0ZbwKnuMjDIVNq4xIYNvI94fZfB/7prRV5CGoALH4Jo3qA6jaiE
aKNZ0Tl9sGw7/w5ku9fI/AnOtFEgHcI0j+sPS6BmfTIZuv+v7RNi2zTpkvmnhxdg
QMpeNLSfT8NCjujI++TuHiuk96AtWmymX79Q9VNrH2RzR11sDzSgPinHCQqczkGy
M3ZPe9uuWJGl4kjJkTY4YqqaRkWsFjUkc/n6riDSYjO5VpJ2Q28uincgqE5/bRZH
AubIbI8qVG8WBYTdfNkNI36M14Kzey9LHYJUUaL37w0umEcWzrRThDQkOQu6dm8N
g14xj1gj0zQC7FvzVBnuhx7prhh/ZOrgV37ZpWcvmamFMOOR9vos0D7GflDK8bof
0A7xgRaqz+dF8NZC6dxT4vh8Nv4WrALFUzIb+DccL7+7/H6bajg8D5dMQiNIIez1
WNtKyjeasa1Abb+IzkKXcw+RIzQG1A7D13LA3r2q5kg8Eyc63N6NgFxD/4T8atwf
N26xKC2W+LMfpUyIbQdA2PzwA32kG2ev6VgYhpX40I6bPe4jHpPD0uIXBQvISeLl
pdq20hPj4x8uqRn4K6kiC4dqOSV7ZrMN0vGzYtp4N60lBHdrydY7B8N6zsz+7joM
TejnJGmw/tA6SEirienD4+dgS6SPOCVHboaggyt8LwLif9ddBhlI8R2clcWHiKTK
wperAY0kz7jPxtAwKcR3spIiTQvfWobyPvfjt8IOogjfFn1DWq6oyGn95ids2qeL
EfBYt7IhavLLPJWSPEN9h98G1rD0xMhPQXsncTqg1QMlrfcrG2suxYa93UJ+Alu/
KzbS42S9+G9wzPm7Rm7RJrSCvDnQmMxrTS3KBf3eRhg5sukfurG0hayp6l3973Md
NlwSA34wMlaBUHp1Z1h2z5JQhE/cIA0/j6k1IMntrPE647t8TeJCTY9U9hwE/xBR
DHkmT5o48q4b/+J/4sshnFHoJ79LDChQYLs5OOIoqzbImfe6osZq+WJGzPiJ8RWp
Ryk2V8SvW0k2iOrY0l8FBW6iyDB6t6fLceO9XDwcH1OsjQgoesaU3Ntd1Px/Ql0p
nBFpaTLINbxnTG6u2wJ4FZ+aI7gunTdt8vXpWlzv/zKBcqS8F3rZNUmwOZJyL46G
R5qAD78pPoscAhZnn2+IeZqLusr8GeunmGRmtLkQgR9Jk25zX6R7d9xyk4/Wy7sg
2tgwh+qNyDaEUUX0FSp2soGVD2V2XR/rcSj+j4+cutA8m2RzHv0SrcuyEmCSPzM5
VTVAgKp/A0BNytus5jLnYs1m7QWKf7GIoVAxHFc8+ewteqDKbX8RW1eiBNdpBURa
TMtc85d2Tt5zkiUElNbQ6rlpYXBxjoYC/5UZZKmGkpfoI1GjIv4r6yUinGS6GjJh
LBQjrWDrblo99Aqepv8p/V2t/ogT91SmMq1k9UvviXaN+LBo+1Wbd6axkWbZVzKP
E4Ao8A9by+KJ4FtVQoLFNpXalAJVqEn1CfLoW82RfgjbqNIyklKqUydxNGpjhkyh
k2lj1yAQebB9Y84y3Bzmvt4NhxYQfQcm9xZ41aAkd5saD/JATZC58O3xd89VMXBS
MGyG6LJHRMzCiaC26bTkdOijNMDab4ILuZl7V0k6q4Vt3Q8fH19DhDGzwK65UAzL
VHelv5//DIx8NhEFXqVg4sjcoA5pAtC8uEx8Rl+Kp/yv8Q+hELYJlz0AX1DFBtTz
F1KCieEHiIBEKNZA8XUXcjJrVHrWUFHHqXx+1avth3fHiH8iGesl92i+1AEe3vf0
Ze5JtFxhN6GSBQs4ob61eDT63LV3Cx+u9UJWIFZQ2y6UiD5JyF6JtTQh+b+BQSYN
Z6kvJENK3NWEandN9gx0Y0dbcr423p1vwE0H4odBp4mOBUvJ+DosrbjGJfLA7UZh
H4cRC6SHDB6fHXpfwwpE1ZoI84rmt4kGx5/7k3IDHiWNQ52RE2nfZyOg3JuSw9PQ
cMa60EC/c20PuV5Jo6EyK0zbI+brhpASzUKyjuX++d6ldQUuSIpd6vCnxEZVsCpX
pUV4HlJ4puizhJ2v+TDpOMnD/oTJJV8kAgWgO36z7h+25PHi0DiBdKxzKAJe5JMx
S9HdACVDeKblcJakuPFD2ue11xNw0UifaD/t/RTcHp3lPZKBv9aMZbOuW4Sa/BZm
blmnYLxA/pQXFSLlf88TAFxGmub+xRB+PpbjG27b9Gjb9qKNHaoEsQTAyhICGuCx
S+BDyYWJaEA2b2pYnkUwTvOsF1gWeYHlswqjQiadivBR+yc/dNFAchCG58AQ/1BZ
nnfLBaRdyEG0o7KYbWr9O58yBgiZnkoCSJWBUlvsbWYu/3da6JoR6Wrdbedmor0M
HeoVVokfoTR21AoUGvV8n7FFXzz2ZmZdjPctpa3t5bySkxtdlKJseBszL0cpXney
2QDp9dLVFBWYVYJ+spPKSdZjyXuoneWbSvh3STigKdSMgBuBp2OyRPeiHP7o0Wa9
FZ3o/cCAaJDVgk52AyUnk+jr8F7Jzp+9V5y/YKzW+PyeaDYorhYY33Klks+khKfL
gfZr9I1ldcG/P0O/5lUKngzR+ZsjHB71CrlXOjIfxcDfHOemBFOCcIu/L7O6ohPx
aS6PqRMO7W+t1L2oael8RVQzA+igTTEWzTzXnOInZfYsf2EvjdIQWJc51rtA7kqH
nHmy2SPBh9dmpZp6TtUiPedQvs16sTxGKRmPfOFlbktK8uaNnOjHmN6ePkpZrQdQ
OSKwEDM6I6jCURxW9Ui0cPZ83onrcR0gR/KBshgPfRQFJBRUodekTt++KtvWzQaY
WGlKZS0l/+SrYOvkpwQw6onM3jBqd+EwjGJ99ylBpzZU2bT6q0xEfn8W9m7+PLnx
dH9HZY4xqPX7MFn4l3loHb/Swj9j8xeIHxE+iIw7voMH0f4lDmyKL6s3+9D+COhj
nTkkKfrgtGmI22xkNlMrrYo+HWA1BnHm1VMqEsyYGf0AxDcKREusK4nxlW1DqSoB
r9Dej7ColQXmvChtE02IPgQwTsevPT92WrimPQ8MYy9HC9oLTgZaAWrcYsZkmffB
f79IJHygR0FuaiQteS56uA6vLqqRF4WNfsIUkxCam/gzTf08LWQATRRtkA6BWiOq
vFfxZ0Jd8oBcTH/vsUQNLXMn7hjKOwzNXbjkVz4hB1ZCNKU3lYu+elIsVGXFDr6w
hWUsQpmM3pKCvA3rr77cP+TpOnzLDAPu4ezqCQAPMSiXu6akxQGBm32BjKFpxCdB
KqOjLkZToS2Wzh0DPcUURUasXeexlXsoVDaHApuX1sBVozPT3hYVd5D/crH90SR9
26s00u3YM2icgcmzSmzXfX9kxPiBil5m+O4To5lNZUVYhvE7vTpyFsGjqA/suPcn
LAc+uRVoliXI4ZRVkh7h7ENz4eCJYiQVz7iMLbbg4FyNUoKiCX0o+s2fi93G52dZ
tUu99VxhWVmpW5ehSXxRrYKvbEYOV9lYVnhTyJGXAhoJhqwRFTwSYo/uSGjKhfRn
cD3YX0n7YEsHUQxYF1R6TQ6+LP4K8TcWkdTt883OJaDNEU03NxZjMf7MEAuF59b1
NWwYjBf2ikaEBSB2yn/KySrHdSWq4YJCJYAfTUny/JzT06GpQ2mpXA5Vp0+FijeS
ts9bQ3y5KMCfs48Abt2RGMMR0R00BDTqjNtOxVXj/z/BMwxUj38+dd6B6j7ZhUn4
DyhnBjMZGSkyaFBvBcn6W5HO6WFNfjJ0g88bv2Soqb6I6YV4P3Cm1C89AFlil89R
VVUUA9ukf3g5pzS6DDGyYeu0VY5LBfv0PQRhCbpPG/jVUhlqfXua7SLrtuClGMrg
5pqOHmZPHBHao9oS9R9fZpoi1zlFL26Uss9eQcFdnyUrexKacM1rMAbt9iXVbdaQ
CiktZGNGhwOXlirBJKrwc8SST6De+Tw0fgxqobgB7+JL1tLWglcUW+WsH+UbWtor
NrBcovaPklAiqtJIijiRhko3/6eVLyODQVKOjDIJmjPwigBu63awaNZg97Iu5/tZ
ztt/cTWnQL9AeOe+pPcvt5cokBfZIrdnrkp5hUjFsQd32OV/KG+qsjaOLhQIWtDz
nRhJ58g1IabFDm7D9usX7310Je0C1JEBgA355mRIKmnt8H2U0+BGxHQRxz7DgGT5
A2B3L+bAlfcQ7xL+bWrbEH/6HjJaNkGhb6ILRCRGno/X3L77QUe1YRRvwgNkuRco
3JxTg92XeM65huiwX09KjGEauDqs4pjnrhqod31oFaLvUWywpMlKEKyjGivs/F7m
XM88AnaTv6KdYIrvM5QPyza118BZ27wdVblWIXHU3I8pNnpvd0DS763mtblBZDUr
V1po14nrUYgWHFOCypm53y4WdJdGmNgfnYErNBK3ZtPBiT5FXiROuLxKuVYazFPl
vVKrSPH6YIMlnjaAy0d5MiAkyAjbgdqc7y0yyq/MnMT1dExLEBlQSCDv0slk7AdO
IxNPPLEI4ayac4DqEjf6RJM2qnKFpPJAsWFrIvkxABcMML6yqMe2rpqIiJKj4D7f
SAI2vkQczzZUbdXol9pzoeuql221cCZ5eupaO8foARncy1DUMmBrETJOJACkB8qp
xapHdPNtFJCgGXRmtMdHfMGopkYkzth2TMa5qpBI+Syt5ZiWpSSOTOSPCJZ9r4ij
Q02ii9p63VWZLzR338UlW7pUtj+ZR29o3S5zwppaG74aAjjzhZV0aUZHxKyjRrfC
vfSdyZQ7dVeqPKPotwFYjkPlN7WUQMAA7RepbLt/o0COea+IMJaw2riXxVEX1YYW
YZk8z2Oj3vGkDjcXm5cNj/FixUzCQQv3ZWMpWLp3PkVVLY5SpnhOsl40Ye4l1my5
nj2rDvzumfmyYOFXG11X9IWY/mX+xJ/rtggChBnw1EB5omdUNgIxCPLjgpuTcoIB
J0bswrFncsvPyapdnRdnJB/gScOx+kh8dpAbgu5N35k5OggWmZG9fWCe7md+xBD+
8RvUj0R8Xj3RFEjJZh8dYIPlRFmcRzdrOTqwX068La3dBqY/IqISgaEt75zvbLXo
JQZYMbbFQNhSvjQxfhOI6oEJ3u5McPcQpHTZvjTBckfmGbDidxk93s9JgTrv0ScX
b5x99Vj79l3tJs0tVq6y2pzgYU7FpeZK1bn3Lg20bDYIGatWXP2s3/VprMjU9bGK
lRiEWl+rhAYlLTdaGYYhoCfGX7sdoOYytbsluC1+2BnnSc+sQVzoeRSxiWSwoqDR
esY8HCf4t6rrSjVO1IpQfDZy8Tms8B9D8dxQl1gZcwZ1fyW2NT2Fdc3tfs9Ct++E
4+5K1AsCeF97QZ3jjUIYnb+BkbseTN1Gn3QcDazn3xu5r7Lrf5/dYbUUwwEr5FMh
zF8NXXkXlyzm05smV9+a6+nuUgL1GWy2ry3nP24C3C3oUeCdDbF6yO9msQ3Jdc18
jxyzYBuFEwy15a9YRY/uoz/JF+auPZgExZDbGVDC/NkH6kvKOarxV8CXDnorSed9
wt0ll8niAnyjXfPdDGgRf0n23l2dOLhgz/cYJDfOcfWCOTEOf91FT6qZr+OrAKsz
0KwO0NXpM+Pmsr9aPjnQMgtv5CiDnrIefKjYZBuxn0gKcb+KkGHgK7mupjfti3OJ
MQFUw0NqZXW6+6Y5l1ap3Dy43lzhYnbmPK+LYEf7R7yKb4Dpt1YOI5VfpY43Vmp+
9JffAThEgcJeUVose8RrdnTRnBP+j2XSkPKX90pvHOOICriR7AzX1nfL7xhzgIo9
V6mzE4GkNC0AMKA4gXWGurPi3Da61jVHOrtqhKRP+DKT7UsFu5UnpJ+g/kk+HWv+
o9nmOrmvmlu61DFNp1/ZpQMDLM6/WckeahaQP95CmK0zwPBEcbiPtyuT63iwx2C+
eJ/T5Ws32fr+3wetRy2J1knIR93hoggWMzWbuJzt1WPCu7pQ6rDU4s2ucWU4R59H
Xgije03U8/qxScrdYzW4HzxN8vvcKzwKkVilJxRV/ohurDdf2dJ4qfSWHDDPvpoO
/08t8kWCZ1ddZ3ZGt3WwrbbCfprm2mwVpLxRBsy1rz5grZ6ngQ6dMkVvNLOdn/3l
dFflaEU9t6iANek0G6B28CwIUB0GFYHTXSb7uzkbKUDtmm1EiUZK6nBRc61h1Bo0
rgFB+AEdvG+8tqM1lSvbRorMCRmkSMD68zelCmXAhk1epa1Km4daVZFDiJC2j8CL
nBy9RPCjfDD9PvvKIrkICXazQLu901SNwYz3YbNKfjo0SS0jkssZIW2POO9vUSvO
vloQVRJFSsp/3GVCqRHo7RxUOeVa4i93TrWmmLfQqe44Osv2Jry7w51U0CDNM/nw
LczKeNRSobGK8o/d+nBftQ42xqMIVEaGINVJ52dx4aXcVIzVLPDhr88Txc1VCvaZ
k7J/y25X6OFbLqxqJY4s54BBmqUlsAfHNA/QeFIEMurmvrJiGuUv6AV7/jCHBmGg
BbfRAdAw1zlTjnWrcH+oqYB6FeNh+pt7D1S6NdM4li3jUduGBEFK2cKRqAlGtJqO
A9pCQIcIOIJRfyCxIDxb9oqHyg5bbsC1OTDdADEUmN/2obJiOsv2jf9rwg2oFqga
RarKbV5ZRnBEzEAP8UaLYXzcXTpivlAUHvSI7xMlg4htKq7XvJFq3uKe1QCTrsWW
GUvDGLVa4pFcpdisJZVC0aPJbgL8PneJns6BZ1QYOhwlWM3R2k9AtWw8JxnJqzwv
Pyh0kt6xJjTpV0UxA//5OWemxecl+fdqevZ+4IYpJUaDbZul+jXoK2hv61c16UpU
DT6a1WhWKxUs94ibZjNEgjVYRzf7teFH3nt1CN9Ty6qwkXiK5129wLs0KlZyo/3g
QWl9RoOeIaMFJ7QBm1PgqeJScwoXcmk4cJC7ZIHs+3lhwaAy0HXSVK6vVFhIDtr0
zD+m0Bacpo8EhGxe6l59+0eFCwjKvGnvF9Wt1oFBAPk5J2WKtY4bjg9/u+UyogEP
LX5TWuagJg8rAmjIRRWy8M94INgzMcZ0migtUngkKXC7P74QTrcKclKr4oQhPcSZ
mhZqccvfmPeR7qUqr8kiYUezG1v0xVr2LQLADI0VOBHT4sQRMdSpgM9Tb6aAfoK4
kuhGYxq+KunXN7l+mr13WpVxOVG6SpAuRjAMlfQes+lzBDYe4T71gkKmXsuOrLXe
+rydYlDUeOr9ZcSSjaAdK+76IBfk00P7eq3YFi/ox6Sf90C9x2l/8akhrEHqobSS
uDNdbo4sqge7Ox7P8KY30Gp35Y5wlkYSkuwV/dtJYoh6F7OIWys+CYEI4BIkC5qy
q/Be9Wa6pBdOzA957o25pVfuzHbGHn4ayqr9myvZ3BTbloM44CAbmiEUkdts3K7z
HKwpGOmVC5CLEjS8xKhvi2mvHkVx7GUWRVd9G3NWvJuPNjEt2u1rxK23O7GqKQsN
ftrHdY1T6qRgv715kyuqw8LPbm0QDj2X7qUD9Kvw8MUEjRwW9wlPCMWLlYIn5+3u
W+2d9ddWy7jx0/s4/xAyk6nfQ+69hvlt+q6Z8j6Sn49NpmDIOU4PJII8Dc604JsD
5Fi8Feo411CxeNOLXdgFIUVPGlCexB/OzNQkkrzi+s2L5FmGhi0hF7zTvkDnmeXy
taxWAsp3KpNM8c62p/WYpTnEEetykbeaZK9wghCC2FyM5qTp7R1sAWFAnSI88MAy
crE5ntGfwyfLQAQZh1kVItxENAcBCBRO+yMoCS4fvhB5xx2eDhj5vQ4CtJXCB10q
S/UNE9RdQgOLruB6Z4a6O4orjNYOJgFX8CKHHoCCWrkBEzvfn7TYkzgrDYAtD/ps
+FGos4NwdAyA9tzkz5JOLylBJquUMyoEm5wi1H5BfV1cdNqR7p/WFNcklFPTtFTI
cn3Jwtl6V7Uj4Ki/nTGZWZX4v7v8yH7vH50OBgoZczIIdxehfHu16DMJNfyLXxS1
fjSOmdMxZp7UuvmdwIkUaTZuqVXnQb1KKrNKZVmk+QZV59Br8Qd2JxLuafvfj11k
T66ksUkPAjOfr6Uo1WN29wB14zmYEaAvyxz5rBFwgGNapplbVrhm+EWZ42uoKxme
gG9sOhBIgRrcelsc4k6tfSIBjgWE1xJZpwssR4MS4ayB1rUgXR6IbYaU4PmQWpjA
Q2l4NCEPnMsaD8mP5KTweisSyiv2GzVizTqYKapUkAiFDhTVWO6Cvn1aR/0DYdR4
DHxpNrBV7zWwhhJzEEP8nAtPXNZ9ATKbSgQtFVuX6wUdacCm2iYRZzGSm9kyPYqB
ds4pcEovv5D56SKPLydJ7t41sfoOOYpdR6CiQUFuzasQGBAsTK5TxOK++uw56aA4
dBe7M0sSSVNqFcfBhM4+dB+ggGGtaiHmETyOTGCxCwJC4Y0lrCWM0dBf3PJr0SVv
rJg3qg5L2YhKPUImIz6OFDoflVZ//IO3NcBIVilIZKwJ9LqRJTFl8wmAT+td9DZl
R9mLyqaDGkAu9rlqHLy+xQCe+N71MEcw68nY001530vlvJo25hAtZnm5qYVkbHub
E1YFYjwAdqA4lx68xASaP/6dcrLQ1e4KNwBKQYbqv6Xao9wfNXLsRdS7KSu/b9Pg
iBzITeIxm++crU7Sr5KcT+2ebjOnosJm9qd6eToMLIP2vu0e1lgdjrqNQPD7YRel
cW4bO95BlYw+4TlUHhu+ueopIoUFaA0q3/w+ZZUPCnPYgHiSAok4MytiyJGKTEhs
WR2AZITH3MKbHTovoqZIsuqGPhYXjt4lKWiBCSVKviYP1FhejGB/pDqjmu1GJKiP
iPnASey3S/NCPiWjVX7mvtMtlXSznr/mDf7fhZm+DXef6THEJ1M5KV1ER9QvPWG3
Zr0wolgdsZJja+MObEh5nzoA6BgjE0FinoQP3Fa0/aGk565Oy0I7yL/bDR/A/BbI
Q5yjEuUxidGdj13LmghlBV5iaZuzy850Ruhb31YYRBdqVJ27zAo38HzJsQoue03w
qWByigP8sfaAmKdlkKhCgFKbQ48vhYwA2rFKHa9L/T+4eet04xedBm3vnM5SwpW+
CqAK0fFG/7xp/Qd9FBFchxMoep1I0b5J60cFfhtsi6hxBLsYt7g81Ya2eZy15yga
7ygQL95EEUKqNBtwkRdPhKZhff8lViri6utxoU04sHy46Qh6Dvt2qGQeguLeG5vk
dYh52oXiIupqmj1izmQkOtqamzQds4rCY9ZbmNQau3cY3IH1Cw6friM07Gimi+u5
5UwmfU4lXx51B1nKVe8bIm9xnGRjQInrL29RLYlZD7pAKU1ffGO3NKWPW1T2TFjw
t8goYW8b96WDlJtyD4NARU4NHoKFxX+sx3l9JEBFpcijt/S3az9cO2dUuBjAPVpg
gv/v/t8AudSUmw7B6dtKDeYjN1raP6b5u9RChLEhEVDg2gUsUeIRGHiZYHYOt6Ue
cfLPXcZ7l+fSTSy2nJUp08iv1+RzA7851nFeZKTn+eAI54YSYuxcqhKGSUMjp9v3
9XeVF6xIpSEtzVU1Sz25Eo939hVt5q9FEqWXW58ErOZsjDjfNpwcqImhhnkHg2jF
6DdM+cALIHoINZMz+BN+Uo248YAM3aK7rh4tnMxF5U/XS6taqZLdhq273itXXDxj
vqhVgRwTBEyzFSac1FjuNwsVzkuwUUF2XEdU+26Wjz4eB8eJ4lBxPRp3zUnUFSsX
hM2ImvcWleiYyACNsoDsfjS0aJW7/Zuhd4Gr1ZntWj7NornfYhks9Nw/BTBxuyz3
qqgHiupnzRR7blNCKESkjTxyRJwWySVqWrCbhsixm7cptzjdoKbXIJ8vbi8Yt1Rd
CNbfscgWlWV7Tri+QM1g1tbN28mBlp6GGacXZEqYBolWFSTblkCrOaMsXmGOUgkj
blSxT3z45uwHrEXKqijMj0Yu3cltwQpwbGuwhxDnbb3MM4vdMn1Ki0Qx33X3fUPU
FDBCesq4gdId1Wg+3nSCksPQCtjqestdRBCD1T8hwNS1yjAH8aWXQZ/WBTAeDopP
JhVSaWGEMEvmdP8GyYRqZSjWfrdeukcUbbGTkSrtCo+7arJUZjFjzkzugi02017V
B9J489tpqCEsA2rxDrokJzzOT9PFKFLjqmqQ1v6ZCztKJxMU2WlMZIjhgcz1Hpvm
/Zmp7C2uj9lphV5BWsPKhZPO136fWZIC3Xo4zGYFox1U9Dkl3FIExdMIf00iCPYa
4o9Xu7gxkbLfdjWWF3Pp0g7Pr2Ai94yH8UD1f0zVIznhIFjPmaNemJ/3NQx8xwlt
/Q5OYOAnAuos/5rJAGg8lO0o1vYCwl2AS6nne9QTFRciADhQ/kz8g1tR/YfpfMiD
Q6YLDt1SWRsPLwN1WG2unOejo3ieTltyWQRMMPXCcE8dY1xnUpqdYYgNl8LjaVh9
Tpagv/D5bt3T8/tKBBI91O3pTGEFNgrO1H8c7pKZphj1bI93S8+ma57WMZ8Jvmdn
MSsRRvZR4WVy2AlB90FwwgviEqwzXXI38QkyHXUE6ezpqjmwBS1attDF+nKEBncn
x1xlqlIo6mvn58p1APlScwCUS8zYTpU27vPZKoG+nkQXSZ1jPt4i/bFxtPbtAD27
ffZOFVQd3AjQ+01fsCURHz1fd91zn99qc8WoncMfoXVvuPOfT3sLUiPVGzAiSMo1
LEFPx1JTuXVXSJDxYCRK8tHYM+aAtQIrauk0DtM3qQYdVnqnbFPKSWutqwpD5qzI
nYDnK7yZ+t+sZQSfy9j/0FZ9rjbRsafcPYAulGd466T4Dmtk2oNzU9UCBwOKmKxB
gx95kTfis3h6GCK7DEJP6fBrwPjfHmilTqbr4kaFS9NrQOHmab14sKvgqtPL2D2H
2GSumgwC5q6Z8n0a1loKtimgYE+skzNVyrrhrw3MfeJQEORfDELnIppdhQVLcgC+
g3LsctD40vowcFD+cQAM/I4LeesAyvTl/3xRfB+0cqRuzXqiIAEgGmkodZXMA+SO
GSZQjHliWzRYTcsR21L5L5WkBWIVc4dtriDlipwSlhppuLtNaAsbLpWucBiQRa73
X3825ReEgB0DVKLuxJGntAl+5K/Xb0I+27TjSUGrDAwEo+fuIQnm9TCbcGQL9R4e
av9sLTJjc1BJvfgwwkTB5JKQIVviMSPfL5nRvaWZCQOF8I9SaaiZRHgW0IdcUfOH
nhzmiLm6eD5CPa8f083SMdkGF/0MB1Irg4qtnqDNoxzXPb9BllXUixB2qINZf9P9
aaZjiSJ6tPlDkJB9BKxBRVP2HRlYthqdQ+n7p2CAJ6VKptt/V22hT9qMES2wFL12
CDU1lTWKDEWBNQ/0kyGUufnOsiy4JIDljMF9jP7302TbZGKLvj79Im5tyFwKNj67
4XVkGLDCfo/qUny8t3Y1kkCWS3XJqua4IZX/AoZUPIDlGdvisuslohNxSsIL4JgV
ynLYLPFjLDy/csgighGiHzAErsAuLDCwfXLsDWUdZMwrntY1WxG0MidfaegrUE1D
bfjRpNQqa7Ef0baTlAZHgAxpkbksJOctuq08CWdRATIDENnPY2IQdH7+71iGvq9X
C+WCPLlQ2Yinrcp9SD3v+xAbVsQv+oBCrxnVZiPOvgSRFr3sLFuH3Jp35GAfa2JQ
eWMSLkuZAvts9i8U9TfjCi3O3LtVbgdumyipV5NRmToyYp5ifJixySjkf3TNgV0V
vFh38oHjKrOGc0IdHVfdcNOQ26RDK9pqe9CziPjb+AkdGoH/i1z3aNEt86IbWStT
tk8zlLeR8HPy+uBDF+AMzrkUekEkHXBT3BSaUATSHC3//HoE5/0ZgmxlAM0qliyB
XbcihWtbqCwpyZ5nKhLHs5RJr3Zfv5wGqcPfUmUacqW6uN2C5RSMWfIXK295N4hu
DMswdQV9uRZwkkOYhZYE4UFzlVZSNIkzHXCXb4EoLcfP3lgUn3T5OnvZH/sKvY3o
A6sR68blTLSY9Y6izGwyWxY4KVWpltzX4Aa7oO4HKDBKS1y2IC/qmKMQTAJK7iLV
9yDrgjUwHW0J1hXBlqY3gfE/trNSLJPbxpa1G3C9r44fSRpSJHPDfHc6Je1U2xt+
SC66bdJ8i4wa330vdpvUrEQtptNb5LKiksWNz6TyjF0xgOPr/CfKkIZuIWe7svmP
6/kJvjjJQBKgp39CFOmWumLt6aXRE64fUDq10VTBXGKbCYauUcljhdkopVGOY71n
SvVZhuZjBeTt1zn8wVOc2YgIiLYLpeRd32bLkd1Ghxpdt8zgO70FHEKcQOva2bpS
PyJeyK+KDjS1FEGI7OklWOwPOf/is4iGHWUQtvRzCMXgGwvb+uZ03N1nPHDVqiCx
+7Zo2nuam6lYU0Mdzuq8Dk0nXCOTOWv656L77oY3ET1uLxQcwKSdSm9bsIobv2xg
Jo0FFdP9qJFgR+oaArXtgbzNcLNvV+qg0Z7g6Zm2BoYLEh5a7HPWF3Rvz7KALQDY
faChZ1BGZVINV7FTzJ7qdWa85XqTj/l3vapWP2GL0IfXA2xA9nZ9If2/9ENNPsn0
X58mgWc9bs7bE5fDCDl0RJwkfnQohCmax1KLXDRTjKXfdb/YigCUf2W7ZQYfTwAC
QKddZN/H07cZzvKNeEkgLgCKQAjv2ankrBlzh8HXD70+6AF70mSnXa/Irblp3KKr
BHlGgakgGwH7N0TjLTqVlqlr4H8W0UeYrl2WbqHmmtuPTlupnou3VRezvSxAx6ln
ES5K3OxPwfA1YQblYx+UmYAH7FsY8Kmfinwf3BTghXkimF7NTs93ZcNNg9eVSQXM
OzYOiyubE1obWx0G1r2eq9xbS2uFnxzmmKCrJafKOdocAFN3zQ1cGvasVnKtN13w
Wa3y+w0nWMX9pRNq5MvJX/5LFt5FSO9FUNKABhW8wwGPC+f2O+l6fTKjVsVcknyT
rP2XFah9c2btEhEPqG2OR5D+YKFFji5XxhZ38LWmOXQ9vsSJfZaeI6qgHyP6+ma4
uF87Fak051yz4R8/kC8jHgVcU7QYifdOmXmToaDNDGAGWxyEfTi9EzfQTahFIY9x
mhy0xDCIbzEkPYs8Qyi4uJLEVAGEKOdgOxXA5eCHudwWvoDvElEdSXkGPUA3UFKI
/iYM4RlVlV5fZfMnCoA7MBImWv7POKdBEqCfimwcqIHT8+LLus77nRb5cB2f8NAM
CWf56gd5Qk+n2P+tQSMecj3w6Hjnmac3GwpJeZf1HH7Oqlx68D2f8vlLQJmdELkw
ylemWQs+pQKVEMO9nTmHnzFBYDs4t/Xq/l9pATP2Fe+6+jY77X3Ycpgv+BFsyn9G
vy+UIh2Slmc4bThPh4Y3Bu4HHMf3if/mzFKn++QFwbLfpS05+87TN8xVmuX7vswe
VZ/mjPCxAbLYD466uRCYmLdhCEXT6xzhRCl3E4jkO5A8RpVW3YKu0o3KRsjk9AQp
OZ3Fu1D2q1kA0odGOuixAigyMs1W9ibtV6eV5VBURcppexC9QfU/F8ClrgWS/vMt
t4gc90j4xFsX2lh57YGYyWRtWHADuNh6N2NAEkFnAvTTXMnc5dAoYGFV98UFcrzR
QFfA7ki9lfyqwnrNe8QGb+J7i/2Ubs6SpP43nUvqBIp4wl6ttxn4ksAfpalXpC2q
tX7kyTxnBprFj0pWYcPhKW7mfwhcFj8aOc40XGUhUxA37a7G5baVeXW7gV03or+5
tEK96p5vWBaO6tvgJhCalNh6jVZAP5DwkQ0+IugMKZ+vEUsXEw3MUG5Sbw7VNXaE
wkgQsqqutDmyxrn9ULYFZ2VaBoAM4Ib/eNM1nAmn95MejNvQuNua7bDpSQtsYJJ6
coJtOBsP4xDIvlqhrIJ3NshEzqaey4IiQ+ut8v2vEqWozYzCmUVTMTFf/O+R/IzN
Qxd1Ay2hw9Rf8NA+CDbefQIXr3jg37Px5BBqmoEWX8L5jrPxp7QBEZkCY91jbSHw
AziE8jJ1Z7JP6SqNCvNGYiicboAFk0/Vm1YpRTqRTS9GvPW0jlmk8vnJTNuYlJSA
Q380c4rnyAfxmT9Vv4giCUYYcRwhQCSdG+Eccu3ksfB5dJ5H0JGj4XjRpjzOVmXC
F6/go2aY6ju+4MrBV8KSz65gCNGFo3g+f2PIAOmk3Q0wpxQTfdwK27aYxEHXshWI
PLv+xTObg0V2RhYuXpNDS1mdtopG6AaZ7JHsSC1ad9ZMkuCnGpNwxEvRTKCSNzSp
OubDRWCTp4JzPEveevogPZhMuvBzamDZQXdmxui1vWtu9r0K1eTOLwoYeM65sTjX
VRDfTw47tV9jUfPJLaPAlxEeHMjtbXgOX0hZ+uC3Eurfbw/bq1NVVpCr8Z1jV3M4
jK2+bVbHpFgYvMM1vIlV5BX6Egg17Z7GBLKufQW36ke2Gu6uA3t+HXi6+Eoub34A
afm8zOb5Azy/u3jTGQcH6AYgHN9wY7LKLLbFS+sm31j3DNkU/aXeO3OyR5p0zMd8
3Lp/AnXAO28ddZM7/mQ6axP1EpjA/48h/+D25QvPtJcoQAFF0tIzHKiRhSlvnGjG
uRjvpLbWHP+zbIY86gPpokZ4mB1YMMztouWWqWiiMLNR7M9/HUPz0KB9nueP3HgV
l3GoFUCZcCkYg8x+SsGne6GWeKYMn3OHyhivtC2AKlXD0JOeffPBp/4dosj/C/wQ
sASBb0mdY0rRHMSzMrdR4R56ypzny+zYtTEdX+qFybsFE+dCKSHlAirZ7X69bWA8
MlB+3kGeXRTY1SBNVIHhw724GlDLdUBcLOfh+DtaxL5tWAkL2pCuA2Y8oGFqAbFp
RLCnAugofmrYpkT3Zk/NjURZg3ghApN5Aj1flbWCpkkfS8eph3E/VSg8jlWwP55z
DgtU41BeYF9QZ5wOXAjE4xAFnG0XLp55qMVkMTnTUaODeR95IbWcfcZAOK+LWe9N
D3w9H35MNXBybkp+KdMX/uKKYJ9yGz1efptIb+j9afCVsbKd3OBAjw+RjbvwcG77
Aljm0x8ib441HIP9TOgEeXe5cI8RhDnZDPwrrED1yWp8SnXUw2TePnHQ8z8RS7gi
pxvUhcFZCF7HbuwyJl7H3/bHYn10GcqBhCyMHXGBVQa3yYJUnuISZICZy3XkEYZK
rO8rMrsOvXs2eAiNEJF9TczOSFe+sg+f4UWp1kXtIiLHzH2cHKoZuwFfAcF9mRkZ
ejQDBaO4FA0QCZUnft8gBSDvWa7+UCM3SBkx8FoxA5wQisVdvWFQGq/Rg6cqidtV
aLOWdrpdFZbXUTu7WDxyMEHoTscGyHm7LX78IqtybCZd2W3AQga/UVp+2TkF6FpM
Vw3wqqXTjr4PyPtg8ygQ6shl0aZZLnacQxxSdrBL1AKXWTNsVx5D466+hPKRL/65
umlwL9pRe0CGZRnEfaxSf4icDYjbooaabvL871xUeKjcFLlwQnXkZz2KZkyPlNon
9WrhnQq1PyGgL/Xy52kCSpiD4zumrpviL37acVHnlUpOCubFofIAGcZkgAri2THx
MKw2AJ4qXU0nPqXd6hPtx6orT6DyIkNK/h14hc2zZgWneJ6KObExtwzz/CA4EJeH
JE+PO9uiMMrt/B/NoutwFpEROJpO2BTMVryjMXn2qNujVXqOzF0gCUr3el0Ym8ln
ImH8mEUH2lClsl3ovSd9DPKI7oglMV04HPgY9CsiYjix9q+PXnDEdBpQQ9N+GlMP
O0k6N8iM09fIegsd3ilg7nQxTGUF6UXtwG2ttMkKRkNT/8H2uwVovzB1kM/vCs2b
Xj1PVLK538Tgefxa60hcwfQVvL/rN8pfHQGqpaTGBHFKh3vKRjuoOMZvFdkJ6E/4
VQMGKMCazUf+oA+CvwRHQXk4YaGz3aOXU1dNSlfCpt7N/h7ral0GyX6HOvVB27NK
mYi1j2Di27lY6JiGy8EwdBboo/rzr6l6Hv6rd6LBQ8u9DeioUANrcMnq0pRSQjJn
6FgE6dK8nyUoerqK21awqQ9cvFLfBK2QUxcZ7y8xESqTjX1DzctsiGO80uTQbloP
hKeHfjIAx4UUXzJSZ1v5MMP964X4bEuvIUTpy3ceoZVPwBDgHgVTb6iflSi/r/nE
hcSwU78FQIeUG72Zz4tp0+KDW/qWHf6HOhJV7ZpyezxA82s2KtwrHtJ6KFd5371j
T0PrpIZu2Fe9jXA5uWOyb5wSYufT9aynv5fyMHhXvR1voUYdmGd0RdD9CHdWUhay
85kv0y0Q04V6rdIHRRdCz1I4IFftD3T7kLWcwbR3xp6cO5I42iYqmhfMNdpwBWjb
EGKA2FmNihKnpoWsDD/L/wA3bhcP7yi+aKgz7dJQv05Nugr1SnDF385tGjDz+hOI
VpiuTGFketiSGkkY+nMiMoYyCniMBIVlLZsVSjeBxVNP4NSZcJ7H0X+MAgGer2Qf
Jkx5lXNE2l6YcscJbu1UxQa/W2JLL4M6JaK30YrGyh7MvWE2Sh/OHHpgzKv+m3iL
rVMnvla6zD7eco6xiPszQGm6SKziCyTxBLwsHumSPSiiMK6P+GhIWoUtsdisMUtE
shKNN457B+Or062Z5CV40e9d7F4Wgo2C8jQKOfhX9aR3p5iDqGD7Uf8BE3sjMqCG
yBJCGXrvBa3oXu8+lktkA8Db5ZqBjm7LuhmRSyqBoOz5fd+RbLGGoKcRgPqU9Y6L
c9+nxIndwzc2I8d9xdtrdvkvj3MzznV+MxmqvN4QG9uor2xsqTen6sp3/F0uud18
xZ0SQi1p5Dt1G0e3KTKduUTEncdr2vH7SwdlSr/wCEsFtq4N/KQ8ROQIjfqJVELC
cTnoyIZm4fvwr4Yzl8zaUPt/aYrDS2RvCDGvePrslm6rngVcaEBCwSPOBpYv1pGq
MGdBQpDg0pb+v62UnSuQrHCvbc8edsKKzWYYXJn+7ciJWn5wWDwiNdT0n1lxSWdT
yU7//QGqud8a1Aq+2b8DHHwaviBOf0Yjxe3W9rBZOK+rxTkmhZ6MSlHORb+DXAlZ
5OV9mpMKtbQiPpT7d02Rs5WtXz72yZ82p+OW2/2IvGUaJC2SoPG1i2XJlET6zePt
XF2+BcyqqMNCEnxW9WHNQIKCxlqsznGSkEm8kWg2pcC/AvmJfgyM/gXyYlYF6tCh
s3Bs1GLiyTEfrziPkl1614S2LG38dg5YlpgMnp5Ub6bCFmo9z6e2eQSXL33IcFBQ
YAfL1EbkEjaUtcCc+So2klaQSleXM3w/0ERgwo8UdjqqUphdk/A/xqbqBDwOXNlM
ydUNb9ARmOFZQyXGeAqCrJN3iQenz+l9d7DbWG86j3NtEjtqs9Ga1Fx9AHUCa6wy
1pZNl7eEP8/EiXexsXD95/LuoholgegMvqRjV8NNPMz7j/QuP9hSf8thvWUxps60
Exsu6Y5FaDwu53XtIweGiFU1WfZNYd464WaxSl/YSYXYaz/qZs59ZM3kJHzJclNj
ZbPlk2A45XbMP0mjokw+LQThxpQrWfE4KXyixel1Fo+6Il6LUp3F2VbbLPU15eGQ
82Dgzo8iX0wV6T6GHJ0mHaBFRATTpo1g+FeZB8pCEhP53+/quBtfoyVsb9A+1KfC
qk0DYC4BVWSgNEmAAFvO1ceTR/X3fv8FpLVUOx4YyB3vpR32nY4ViLFfo74MJkkz
J97tQC5y/q2dTpQ4ihnHbzSML5zTV5p9uNuqkbvgYL1FvylTtX6DijR4SRySZVd9
e9FEqVa8GBNf1XimEE22yGyIp6ZWBiIGeAq/zqhOoN4BHJ42TQnagEC5obkG91Ls
rD8kL2R6q4yJ7BP1C3nVL/bOdeHQON8IefgQqpWqy2h0OE6nWMvGIVaxIAbVTzRR
OQS02cyNTGhUud0tuHjeIyQKz8fheLuQXGzGWfzClQdKNP5a6ahDXJQNPHPFKEva
/tqVc+YuiYn4XwmeeVCbcTK9oOfNsN24qoCK3lfo5u61M80uXSEMxQON6Y0A9GkQ
guqpr1s0c0uExLYwW3+A+IwuRf3afzZuOgR9wy9QXwGCZtRWoAfVA3qxERKsc4Wy
9TTp2LFNMvnQcXzRjgaSAqb1GcivTrPIDl31aPqGT+s+4g1ZgaHq7KUIVFds9Grt
KmrHUi19CpiEmtj1+gzNCXOhq2sheslgzH9hZa4vFza+ZQ36Q8zA66rPkKXE9fsm
s130a14yJWONnO7WilQQhYjnGk6J/0t/NjrQNkNKQF9h8sWZclumrdfp0ms8PHg0
GhjNpGwtFiUYCYDxIB67vu4fRmEs/d2i3x2/kiDEmFx7p3dB/aWG93EjbidMkv0d
jL8jDYgD7pWzHUO/0MkmKLP2z0qXlRz7jMXZS5414H/Y5t4BW7tCP9r3PN9qCuDp
l4HQJr1lXUCfoA5RgCwqXiE64POArHfE+M3XB0E/C9QYFFrJSdb34ffnkKcQP7TZ
PCZIliq6pGO3NTQS5OE61+2ENnCOPZWSb7NqvBacjsU2xZ7lsoxMkxmnwYTcRoOa
3EJvIKbokhrzCb5TipDXiG1eVKqKbLxfmj4VGgAn5l1WlPmZUOdJnIcapq4DTVky
8JUiILoITi5AmGexMAnGhacwoI1+5ZLXTeZHIxkDhgBlg+LDOjsK4cSOOAC7GDN3
Fko7QWUZdfSwTxBudrRCMoZRzsEyt9ROmCHOgDueXsz9pKrxtlYliwXtl0mKBvAf
yFnD06GnnDu7Jjv5h9bkyp0VZQnKUNAtPhQWVoVMXA/j4uxri/Gr79H1AZ3bE/yI
O0jSs+BhrOV2x6ACqThrO9DI2A/zXYEStPGh+DI2yWeno9TrzysURF3kLJuZDxb8
GGzHRSgi+Z6Aw5hR4kNY0K+5zPImrYOWG44ZRY3CfPHgSWqnTyEfOnMpT91h2tq+
D+xGOPJQkL4B/qZxkluDyq4FL0oJt/Iy5JtpV6k2i1O8BAHqMJyI8JXSZobc1MF9
EkWWL4iVMCyl1ILIzbtqGkXBfBYBEsx9GtVaeH+ptp/R9Nfiu9cmbi4b/WJpyK2Q
qz9CjBoCIZs+P/26buaYTb1oikHj5/wOJ6wR2M7GljPc1ZO4Eh+5n3NXsEw1og7K
l4XlyCMDwWlb/u+EPC2qKWv+qGMA3xvhpAdn8rbAQdo0zAqNmvlVM7QHZwlBHb3F
1rn2FC7OGpXq95wG9IaRzcYAkuC+JoldTD5RWEzqZ/ZGdwn4cx6RJ4VoKbIWPPb2
3KbAsUFHF5bUMv8KGysFLQ1xbtN7vNvISaw33/sAHOdTQU1p5F5BvWOtKxrRN/Sx
a4lY6xv0upIBwd4HnVwIF4fgVIRAO/ZDcwrxVm4pMg2GUtXmcJ66/fU5211z6y6g
AJOMwiGty9/wlSVlOmOzhfr0ZNM8bunmwGkk8lnSRLpqG77w5k4zhPHqtv/APoo0
pQhCzMmSn4qLjfXVtZnWgYOaQoZ0Fe7emtyP0+l5xia1MDfWotMQfv6dcj2e28FE
D7XN/i8Gd40LmWNbvv1hHQAdGwwZt4FZybrnQLoBo4c+zxMmrglzwN4LiG7tPoj+
820niuMXJi2WoMMCe08xhS5oVFVwo1JCXD6YCHZ6t5At4/wss2k3ASvLzlcEe0Hg
LcsUiB575z+d5RJPPIoP5XwlayiHpO0x0fDh7KqqOOfvdunMHLXWuy7P/vmqLErC
8FVLhTWuI4Y6rRYdIaWFx+ed2PPu+VmNzQKctRkEdAv2zKJVfmKroFgRHPjFxzv0
XmludCEtMODAFLN8wZV5+lG5mmfvb7i1gUwTkUov2CTGk4e7NPiPnK9WuHsh5oPU
KaRhVeNG3BNFMe6lbWLWOJhslW+oSNcF1oTKta0OOpSw3Ku8qUJz/vnazqgGITs+
ZbtxHcsiaFNs7mi4Ub0D2v1FIzrLYKR6YxGDJs9BFLC/XbJKwKzBlIXkKUqpXYJA
fp/OBxrhYeAj7xINEBA9mnXV8FuFMi7lNDo4fRdq5IFBTmGYblERCqCSZqnSI14N
kSxXQYioJEYwb3K+MtlZw0NlzcMfqWPvd5lMVf2Q95SX+Xv/1FaNJMFaCv1wXUeu
FqodzeCT4EKVlkHHSoxlLgIfHkqNw0q+a7vGJvy18WmOM8jW1m/ret4pJv8G6JCh
KCuhrl2RSEHowO2RwTewRPBoWgdgv32F2D5cDJmw6M7Z9yufqSaBzmsDmdwkGU6d
URnWzqbivu22lXbvTD+amy2/c7rdpyGScOSSDpPJfADdhV34P3GYSXj682SKdERQ
0/xh/3ZsKkpY0Mn+8cKPLpu8TswezloQ9tmB8FgNNjm7y5AXLb9e2kcwkiqox1UF
szxqPi75Wi0SfC6rcexI8ge3k7vGMtzHokgk2MXMjKP9I2ec47Qkyeng9lMrgHoK
E8N+xeWOal/bmkgzhhYutnSAIdtGoEQ0B1OvKVorZJTUmvGyqxQsZB4mo6kj8e7m
iWu9xQ+1XdYIxb0Y3TnNWwi7LVqfasiAj/KHnPaisqLziCfdnIfSPTm1cjOQ5Vi3
qM81HNMLxBgEDjuqhzHH62RKddcucGw3lSrY2sMvTFNO2+gvRkidB2aDBJMDSXuL
5rB6S81h/XN+nleyMp6+XQnhSg8TKGgv+Y8OP/KXUY9TYOambxp85DNNB09fYgqe
S4gywqGFyHvFYC1eXGoZKNyBJrfdAO+B+Jo5UsRLv1JkMlG0mqgHRsPQJ+fYz8/f
w9nxQsI/GmmkeKzqTSCa7gkVGHGZkya1cQyBZbkDVNQyxjYJadEFOvIiqYFAPW7J
QzQxBpFre9VnqeaPoiX27yANc04bU7j7fwhKc01XSDgVMklxYu9dETuFB2u0vLge
hJRw4c+rOm/HELCGiiW8JokYFNVmJoLsD1HbTRGrzKDQl/BQgBye788QArRwPEgG
Oti6Opp+8httX083FCTgvotN1RY6sFfGuJqtpz6lM+cqw/HOXjeP7ueVCEVILW1i
QjjIcv+Sf4hO51BEnJIJKiW6qc+bq743p23rxEG57YsPtfLek/5yFe9TpJqutahY
/J+CV3P7IwNAlqWMC+3dnlOpLA3FdvAz0ef5OywGoM2uTMKM30rfrrAGX/wOYnxb
nw7ma506FwLO/FmJluz/oGJU++0yCoIB0DV3is87qkVkWxyuJelMW3Mawvbv3vqR
lYtjf+QEKNV3SNJWsosoXetw7BA7sQgBFY1hL+tJh7rzkBPBTB3cFEBfqJ01frRS
jCBvZ/hYcZPigvGxRZk1h1qMjgDlE7xU09a4E6mvMcKi3BoClcEbQF6gOC5BFuiL
dhWZaBkicXWvDGkXUTD09PZFpUkkuIvXnsd6tzzZiZn2RXmormQ1LHkcTrkQxlyP
Hs9qJ5r297P1+jdIwN6Kx47roBxTp0ycNorsp7X/MFJt8Vm1YyeNQFX51hAZYvjV
+c0obhzikTj3YGLwsF1RTk+kzFZQLSqRnfqJdzFikP4JYsS4ohUxQQG9/dKE2JnW
VET4ofsMjcHgP/1C2Dod8oNyTRlxIkwdo9lsUg+7oDkLqEVFgJAapZJMMZD15YGQ
AOaTbE9epFhWU2qLmVeANZx3O4LO2YowyHPBDN1uPdlL1Qp5wBD1X2owaLIfKy1P
t+qVDvA93igRW4oykpbe+4P4kytyW2h8daYE7wl8dzBJDVKcVojSsbVxIRF1w8sq
ENDE51PO+D40IJujb9+xMZWIrCw598M0Gkxf1EgYk16IqNSxcYWQhK6zccPBvJK0
B+Ax7voDAbxKrHRqT0tN3RFslZkVwvj8mpD+Nrzhxh7GshMwDB1O5MHrVXan29m7
udaLdJ0D6K46o6MDm9bNoMQBattPtwfx41U1o+MzCY9wMnuTIqu1TDQtmPc89d62
PuXTL/4gXdARPAlS2xf1xG8JE5/MlWFQ/qOnfNhrtkE+iANx3M19SnQ4tABwsEQn
VCZgBQTPcek8QTHy9WZg6/HId102r8orJjFy2xF+WQPvWu5MdaE5pLMthE5K3Nhu
dAdNirZlqFDWyFrC5lO7Qec3TQf9xq9BwL12djYGM321rzsAB95AX5OR8QfW48E7
zUoprJTaxwjJOggv48p6P4CZLthUhz+OwJCuYJCv5J+eXgNzXGkLYwUQwVJB5G7x
MMC2Yun66F/la3f5VcAkTqFgj/vUMmE2AAyMo95B5dnr4ADf3w3j9TZydtBxUPt7
k5mK0KwGjaPhw4a6YGWx/23/ezCRthvEJ9StVVMarF8MXLfPDJ3txPNN4y8XthT2
sRKTI3t0chYvyaAIz49rpfKgTrO+fusAvafeOOujlclg0I0lF0bhwSX8fyhgBTMW
9aBm/6KjPm6NyXvQ1ZIdXWo62KUwRydy/3sw9NBpHYXNNNpqDtEAeEOIpWk/9w5u
8J1mNTYgHpO47GeofWJ0lMeNfXci64jXmRvpEQqG6BqoLgadDLomi22FwZRnGMxV
e77a8ABxOIO7k0Ud9aeQjyqE4zT7widxg9G75GTEwol+AeiqVz3F5q7RlY8572I3
qSmvf76YlbZ4Q5kF9RGaNmNFTqQLPLJ+Nqvamab+Y3Ob/86dLm22z7a7z5ujiuG+
r7Fce5ZLG3Mmgwc5YDfVhb1/SR1KDeAm4UlqTUAUpnHMTC5ekIveQKk/EPv48H09
PBpANw4XMHg0OJzVY4z2qhgDNoylIO8SxTsDRpuLcLzvf1WZAmaoMoBxk3bcWHS2
Pxdxc/KRCoMtf0Jn9gkp9vgRO0+On23GmMZVQOIyXC4MXiNeswJOCmV9a+9z6TS5
q9ZkU7qocWKoC+bFhoBmXyt0WbC+N0z5bhAKVcNPMIVWbgs7VjcwApvqvhcVSDvS
fdxsN15wlP9VgN+7VdBaJSVvOhLQMYhE2Xh9FOLGTPMBXz8a9bAAS2qvAo9xzYsG
LDUMRI5mq1OGcRlEkKfhzLdd4ENmSjBr3ed71+wVrCvWna+oMzurXeuWDtMQxCZ4
fmQHEaMwC3XCEOC8daqOEaBVNpen7uTyF3TkQ+5s22a5I5JQXey0m2K+b3mxLLQl
YOWncZDg3RKM9pKpDadlAbp7cVMpirNrSnt5Kbt93gLpXEIIU+0lmKJ3/yu7kRfr
IVE7XnzNJ/mLRV4JNAEk27tPRzAYagvxMxjiLzZ0As9Wez8QLMHianTOQowzpAdD
+jTxDZYk/cn79RwydfWpabrIblvUU/3LnsPmSiARaA7ZgsUgQ83IzxXACKqpSvxY
i8p4SE+rHjA3A5H7fT4s06NQuSWao1nL5siVao49+gwQotCkOTvt83biTBvA7Txf
CeK3EWkXBOMzGWH2z98OH0HbyLLVQ6CIElcREY+FLuQclrlq16D1pg5YvPvZVVo1
cp2e2bzuhYpaV2xuajI97vMpBPcSxb/gOMmn3Ga7L8f5syLbd0VogCj6wGE3BAc9
FP71cEcMK0DwWDhqx+nHVK8rIXRgWPJMEm/cTcIcbTsbDU46kLh5ymlue65Mn0Aq
7OImGA95CfbWWWam3oqKsOikgfq+0El5gtlrfWDCsL4AT+xweh3xpEKBXzbmnOpg
LUQGTpqx6EsMzHLQDIqw/gglZVn97tFZ9sC5z9+gQX9oOpnv5FzCgXcCjN81P8VO
DxWXJGTW0LXB/bdtl4zMBbtGcXBv3J//KE6ZHgpws23UICOANPxE/wTBvpkwZ8cA
71jfON0SBLsaCeRqG/326x0cW9Zjjw7+d3cyw56jeEIG8ZLw/WgQmNw6yiZEVQwX
hOJlAi/vabWuDui/dJsWZAB0dQGKGCms87iKp9K5Z/qMM8pC8A/W1vFeEkgs85dJ
F1a8sEQrHV3gEIdDDySphBPtL5L1FcgMiE6lIwUryRFJ/nrg4dhpwJsZAPDDKCTR
zgi8bmN2jr4RD10+WctFjRYHmOPvA26kv1vfLP3+bxOrIRhPDUVlZpRVr5CB6loQ
hG+FWYkLIZc1ddWEwRgT7c6Dc4DDbJ3im2kODdmVzEg97wKwG+K+ksnEqLDjBMq6
Ra8tZ5/8IvThOVMyvO4x64LtYPzaNnk0zNAF9nAhLa43xPYPhw1tZF5wcSsdZhn5
lOMbLYkuFHX4htEg8yI2nLBqJABFO7QFI7nFZnBQNhzITrXi7UTHgMbRi5s5wUwm
mAni3YQaYbT4WWwm4i0Ihe7TuNGTfCtzuofw7Xmr+e5PjO+rEtANjFlBKHbQ1wBN
xxuz+Jbka/HCY224BE+bJlPKn8kaX/asnOoezYHSKib3xsl6K8AQ6Xoh+stiJiJx
qOluLuiVo7Z6z3gMypMLgEkG6qzFOSgUD0PQm20hsGrGnbPDW8rvRtgKCR5mj9rZ
+DGUMC4E95mnKEs9UPGbHut6L+WDr8xul4tl/QwBxfcz1QNdYJ8dArsYMsx6wHgV
i2xhC9hnUMJs+uSNsTW7Xbv7G4LH45o8L8gmw605JOWVcjiMjkbfH8fbbsbKWi26
8wGp4E23b4DOmWQRZqZ0l7ab/4YTDDuA+5ngx9RZgYYVpy8NApl5f1VGjpZEdGko
w2KrD9zMG0ZLh7KZBkWOHRvcwDoz0OjgAIOOJ3TYK6RaMlHWCHctw91Jv243xX+1
UbHPNwylBdLrTC7U7/dS1lAuTvFudZxe/3zF3p9jGzHWD17hYRehAeC+dX945KDR
nSNtM1sNYUAshAv6ePkRVAqzgPNLVTdG9S1U+mu+K3UibnftPvHD+GMRVtdRtpyx
UyuKOxWhbHjCOKs89YwXK4InFo4tq2zOZtL7WU0YTqZ+UmFblRnl9lytmjLJdn+A
um8KakcEzjHVmGX+6bF4stfnnc0SmhZHgFhs6aspNBZhLn14HNszX9uQ66SS4wVw
J4pCIpkPe+SA6ualFyhb2/wVrxIB8HNamj4CTrcM3eS6ugcLuFxn8ZXCTpc8KVJZ
29D7ZbtZVmeL7ceoM/xW6ILzn+LZEgaDwYg+8RsLD0vA+HaZvPBNHuWVYm0zcdJh
3mGYELC4Nd0Zgi+gjZerrm/tmCZ4EyqDyn6CmtHGvB57Rdi7t0rbhmF7U/55WeWm
G7kT18B0+G5IfDJdQMYu1tNzmCt2g7e7WEa5rFMri3YdauRq3OfpF0/cYij8+47J
wNzIf3nyBGCoplNvQfY6sTxHmnphb1GgRQutB9daWPRHVeF8YTCxX+ojHE3vdJCt
3WGogezofZUVrbMxhemDHArh8IhJQmXnLszD/pc2Ps/quHqwGLU4FsWZmGzHqBwQ
JAI9jkU/9piEDqAOXTWvKWD16g0ea27f8+K3TKBmyfsL8O0A49i+3JEH1tgSctoQ
v8u/SdJagvVdE7nMlV3/SUJj7zgfRdCbmJY/z6cWeRaw/4C1R8UdtLc4pClKDlZP
+4JmyruGrtZ7ChRJ4plFen/aOrVVBLFQkY4BuY0R7EuBrs9ToTR76CHzcbtCVph4
d3KcdfdMcC9/K8Rt58XqdYMkBkguptdFWm12E9vHW2PiSa4kqakuQnGn8kRJEybR
nrEL/GIKdXpaXZNI9TaNzZBajetaTBf9yDf3kqtO/7eFqbtZoRxXr86qdHOtBJxv
JTjFIVBPndOlPI8X+uMF1hYmIpcnKhaHOBWz/vOWfKGAGFIkA+WkP0E+zexcfv/G
Ap93qJbJ/JnmUvqbSvhlBx1Q6bFONKCSt6snPjIkNhbmTFaRy+iQ8WdjQ4h4qamc
BZ5ekOuEn6NwQgPcXz4ZUF3SAbpSVa0bXFeWORGtVh0aK1t/dwTICEJy0HlaUFQ2
fkOy9JeT3TW07jnSgcTtdxTQCXNfGfFSu3wwwT3d/c29JEbGXlUii0RnfHK+zUBY
ITi8Hksy6fM2m0Y8oYh4IvxRlm+cEZ94TH5LbhSOHU+RjDn9zmIOE/VnKHWZzpro
/nSLaiqn2wlpLft4+/fN3IfcHnhTQ7gv5/Q+PTMnncjNc+76INp0F0IVavfM+tkD
8AG34BRxaa43Np5JGNqW20uiEn2GzN1uZYSyNj9AuNKyRmq/H/TmXH9upxe9KbFO
v1m9Ll0fjPDlGoHvjNQ+1YjeCGz5f7lcUhmBOb5GKdnhP63BByhVMLAeRnmECGgt
vLp0sbp/Fom3JBoE4td+/wvpOW39+mLPtiAX921TKjxW2PUnm0NAJETHbnY4YCYH
XL9r+3wtzf8FPW/E6UTWdQLOIq1bn2vAaPxNm2oJsydQYCdRXb2syQnDkht2kjV9
yo9yqD8KY9h3lI5IiwA0CRKbCUN+kZvHmlQoe66ZnO4JP5w55N9Xxk08efKupMsE
OH7KJnZzavjAsn790Md2XPKpNB8wKXqPW7K+TwnIt7VSLQnIk2y2/Cz7KiroYlxc
JjU68bxVm9YkvEGb5LTfVSUYXoUFtBZA5kU6gIayAxTicf7SLogWcZJovuCdbMs1
8RmnD4biqb6RxNIc2X7WNRVjJdaPO1D4Cf6C19PW8N5zpWDFwGqJjaVvUfmCkkHo
fY8+Z/oz9L0L/OFRdtdeeTh9BKaRqi9Abvbxs6+v5liQCHUr1T6UYkyMZGF2rVSY
ow915jizpz9ZR6XsjmsY9ZwdTqJwyFnm0XBaApe2WND1lKodYntxq8v9ywOx9v1h
ZX/RelbinnPWWSAr10BkdmbUnKk2XWAqXdS6dxyJZh1lrD6eQuH3HpIATarK1238
zF9lUpwV5TmRGWimYGJFPj4Drh2v0sRa4jauudstjx8R6eqLXdv3VRHANI+Upyo3
+YG7bB46VOxI3ZKAzcYzoiyXUQdzsHv1Qv5nGsK63RZuqCr7Kny4mrtS+H6OfkAJ
JYaWvfYDJ5pmVVWo2m5TOlJk9quJlCLVXPMeQLzwh6MktI+2EPprENZV7IJ/ze3P
XrCce3EehgfvHydwHLPf+wlMiRe5Tk17VGc47Fq1BOpZYbViyddn6SXcW+nkUhUy
mUFwNLGzDQ9LrWdYnq7jnbvANPgCOUYH1uQuTQjfz3lzCjT4KF/LaBL+wAbCs7Rp
lBxwD9372MQZ+C0VcnF2f3aWF/3YYpyBr/Gr7WSledaE9iAyL0RbKley8L5o6VhG
BLqSmUpn6GU/TxsYach1tIb5Dau4mZw1Lya5DDZwzLQwxWiOf3UzAo+nhZ7SF8yW
jbqlJb9a5ENlG1BfGND64ONY74KkN49x9H7Cqr34y21oW1kcghnxVOxismpUhem/
hv6J7Hd0+osXAe+TgtifQOEdgCHoNscW4XQYXy8+oKquL172mXb9QG771Ea0Qx+y
/6XcoFWYVZqebZcNQrod2Cqo7Q8cZKL8XqaP3/fHANLilmkB7wvJgI6s6P+1XMrJ
mWGDSRpBLmCt3uPUQ9u8h2pb6rb4uqBezQ5Aon+r3l8PfwXwHRvu/bIPZOu4qr/n
OcQiJi5bTL/vaOGEJbtXcqW01Wdksk44dqD/lIm/EW7qzKvykAItq+S25l+2v6Pr
vP1xNxe5kbh+HHyR1DfFph1q2nSqG2M6AGfejyATmDmzKBXuBD9VUIdxDbHOZzls
kxKbw2a5LS/CWG/benck8VtCubNGvczTLzRAykk0MDftsLt+Ll82k6bPx4+YnVAQ
WXoFQcraKRAxPOPqULp7mjk1fQEHDKZ8+fAvIRHvqlQKUYQ7NnqnXxHh+QCcU6BL
i3pqSRhcG65zEOwcSA3A4qNGSUa4rgSgbUN3ygli60mYN3FNx0YNpe1r2MiYPPYB
yqpdVeN1Nri+vshKY1SaU2TCMISs6r+m2HLd0a1G+rL8FMMtYadqQihna1kA/ONi
YTcoZgPYMH1/RnmsVqzMMgUN1bQjB0jiID0WhnPGyY/FKvT+TKOfoopo/nXly3NG
1+Uq2QXZeAvT5wGZjO+O4buUFW4XCSajDAxcZTY8h8XjJdqqNhVRSQAMYbOAT0q9
2QAECcXsrH2GmLGAxwpC85qpMAf3zKxVyLLKWk2SV/QebUwlBH4/5sEODP+wEAmz
miFTIb8rgBeO8C3qumyS9Y3TDUDWzI1iQ4CBVjHnEDlcrSN+aUmGxZXqQml79fn4
9CBJ0c+RvJ+GY4iqpTuQfjcKw3wSm0dCZ9fyFKpLTvQyGWUS4zj7P3+4B7lMRMkS
kSMiB9Gbj/NL23skdneER6gYfPXu/xM7nOuVlI4NdhhF/TciearjooA/FxlhCxuj
fIYC5hRy2UTCS9lAZBPQdv2MXk4+VN+xnKYONWNp6Vp8zAUVzyMrzXnlymdOYf2L
2ayJeQ28XYsGwKQTAEIgq05tkEFi6NVQEU+tFBOKTjQMk2vBDA8gjbeUF4aRqafD
Pf2ePLQlKzaj9ekk0lcOTVGKU8QuEIy5dGOC8MtioQsOF71hWFLhVa2Xj3U0CAxS
w6bKr6Tknx25RFc2Ry86Ykvyr1qbOrFu29RnOK2+evpC2JIfaa5JueHZdcf7kjVA
/htqV888T129R9eWXfG/oGPI/zJEPu5Yj7myHT50/DeuueBeEexSVW8tOCBM1KHI
u8UBiMq50VVAyP/bnrWBbm++Q/mwQHuoluKIWUf30qNY97OIDVk8JlgflnjFkeR4
rbYpb9iaLzCS0aGIjQzjXvgZUalZEtHzQaS3wh8rPOJd6PNiP24xpXj7RGLbJhZM
9AIXUdKfL2dCkfJr01Xs3UTbkcRyYbfdc5+Ca9/wRnyU1+9sDWT40gzNPp+ZNQnS
t4DxxKNBkKG5EPWHONVa39KK2gPH2oynO5xo54fKiwEnbQGOJvzRs2HpTvLVKgVx
NFyekhZB7nzvMK7BJ7xV599B6R3vRG6yYqp/ZxmZSlX0xdndpihmTZ+Qaizp3DFA
58qOJAz3Nq5AmyeT3G6yUkIBQZebA0XMq9CjBfHaNeydwavcvD93FWPaChQ/fYaK
GsSgIkhCRG+M6cnk6c0dUIKIYGp5EFYKIRlBhF0a0P/u1ugR++kWbFb3lmFfQUwT
aQMwyNCBidEqHuhkWHgFDMtex9ESG6c+x6792r5o8HzEKESK/wKw2PULzkQpRHfG
sX3L1treMzm50SBidstdFf2iczhq7T4QBgArvBFe/mwVdUCwUEPqMgacOqSUq56k
os56phtXz4OvPCqG3nWZli1b8NgNeOAvHJBrvjEXMdZH+o92bq4A/UKmZ5F5Soxf
EXBr2I1fClJlcB8USN9xweFYtUFUSQ72N0MUAD5lbj54+0Qj3EJyhmMRqQD4KjlK
sRuDUFg4RD+Ww3MACVi78liUpIQcp4XcEEfxVP2//CocBRsZ9nrDZnPRR7OcwCSn
Dog6Xb6Y0r0wY0dcFy895+xcENQAHrXcmEpM5cT+ftBBdW6tCGc26diVl1QfRs/V
2nPLkmP8su1TNl/QiIfa9g0GRgfAohizlDf9mVlmwsFexRWsWyiBdBPYYO788A0E
ZADpgHO7wj4QTwDOV7DrXRkdG1z4pAt+vzLak0qbjXLkYAU0iNfH8jZYcrmXT3Dn
5EkwP3z3/nq1jhRT9YDr0YofcRZo25Q4eGo3zhSNyl0nmrQClA/g8Io1tTPfRhzp
8E/2sOxlcYCzB92s7oCzj78Q2lEw8hdqB3LfvlJ+S0l7Tgrpb6BC9NkazyMciMlj
JNz5oxeUgaMMUzkM8gSJ40OYKu46RBM/WvhTPe+AiOMuUUvkVhauNNAr150eso0C
AaH9A1TRRLSKrvrzlZsjS+6PG21pwiSIXjbyyXHhfjJSd42Jm51VInTQi+kO04Vw
ZLmep4b/Zn08tePuwzpKbmcnTIMTytMb1uYjp/8QlR43Mab0fDWcIbNBQ6DDdsjm
+/YbiqYWIwqVv8LUfv8fx1HiaBUcYSkl+OFAhxE+WpkuhHIIG2daPEPF+BHTKYmj
/98+tcAz2bwLib3BJ0yrSWdzceRboqvXHVcNstA5U5k/whfHXfyaD6bhgv96JoUu
QoKzqLniWyqRj45tDJ5SOJc2MV8lgh2/Aoj+Gt95Lxw0oftdGi9m4J6O5WfOL49H
nRKzKLngvHDYpBkYIKf+V+ujaeL4/oQB+1OhactaQE/Hv4mVHzuCjlJTov3IdM8o
d946aOhxXHskRKd7e6BZ2VrfJ+IamsNG5exkbF2v1cRLK4WFTF5S7U+F7ZNLgOAF
tSPqJ0QbNvrjovxjARTSloHtwhYhOrLrrCPGL0E2xy+B2TsGec/CxlsDyWcdJf2z
HvrusWbCdyJ/yhhVQIew/RSMGBzgBrmy8RWNMjrhBrV+nNW8rTdD0YrEOuN4zZJC
zIgrmVWxKQ/M6OeBastGl14qQJOPDZu/MnMNTEeo4q8peQT02fPege/Rs+ViMjNh
h03zqZeus2uy1Fr+VtJDEnL854g7aLpGXfcs+ubnsRq4mb8coPF6LUkvjcdunhRp
KTrXz9JTRk3CfE1CsRUxSnpg+QHpfK24x9qXqv1lSp/PQpnzklpL+wbeqYykV0rR
0jenWSln/WJfgzX2udl3yIMrTL8h+Px+cFc8PVWQh4x5xr8z9yvF8dqqfsKYUE7z
NDch4wqWE2UdMIi0wcIyVButHQzZSjZo1KEEfg6uASq8mfWDbx4kk8Vz6uR/rzoD
gaSZO+AyKAPHZ8xxDfpZknyr+HhxzOmf7d/8RsS3y0UV+ch4F7NHP6vPhhlbBWrr
6yloQCWBKNjnc87ypFJyWcaSDv4USrIe0SyBulxsJ3ATU/G8r73hvgaTHURkH4uh
Bx2YCXlOHDs3eNeS7QmKvNdoTCHFedlYk7rjSfN0sSdcwksCIq9dDocN21SSeq5R
7uUyiXCbkVtWCl8uaDLE1J66A5el6q3gTQ5fGrmgZb557LYHigCaB3PXn8GhwBa2
mT35KGm13sgKpNrY1X6/VFPKutxJSyyjjo5B3x9PaO0fLE/zvLiR1Z8PqcfA/gBP
Eoh6XWqkzx5bm8rotFou+escZkkfEbH72GCQlwcxKidK2PTttJVzFMQwngGnBv30
+/8aJSUv5ewPfPgaANyFP5KCadRNFztCQ6CWLayLxOEHKAjM0Vwi38yjZNqwCb66
xWCZ2gzKNo+hyCKAAutVgBXoeKBsgLgmq1gVbTktYSEkEmFs4aLQDtvDZjf+cMFR
rNpUxrRkjlF+huhSmCg2rFAkG3LEwk+5woXaygvocRwKKzKQjbSsA7R/XuSFDLJA
F9av+UMDt2/I2UVA5+4W++qJwvgo50rmHZCGRZnlsEidObM2dYOKPv6RGqPGW4FW
qXgRwYOkqf2LgUTgQ0rjqPE0PwYYQXvgolO1v54ZCd2FXGPaBIdQXSXxSB+seeq5
Lgsdzj9zAl7xm7FyDIfGTn21Io+JMQb5RSW32TIWpBU8spfhGxD5+zYXE/IfMkL3
8qiOHTej+IXvGqPjNlvmbxtvSzsBlGKm6OI1s7y9UntuzeVW6UEMR0cev70tKPvD
N1Wiurq/anXkuUZLiiT3dGmM0atX2oT710zWdZRZ87lNW5FBBcwdMS7TNRW+3z8j
+0JaqYvmWS0e3pxBf2PBnkqKADTHTILLTlGnmjYOim62X0Kb7QIBzeavmCNKuRgU
2WLIW40bZsetrI4JlZLhulvXCTXNswqqiG8p6mzIYvi9h8gPEUxMpaiu6YozKoLr
iL7zoOtJYMoxQTS2ifgyZSNj/10KaVBUOyQ7smd79bIGNjRzuYJZvBSjitD44lIw
FSn+koop25dwnJEewsFpX4usBt3EJ5rHmqTLI9mRBl17mG8hcGeymov2rfi0K5fK
BaTUcQib7bq4+wkK0OvLn6puNdcE1uHe6BJLtMfzGO/rsEeDL9I/lb9CK/5A/zTn
EB8k4ds8jUTvO2ywUqVFUUUz0NrKf0SlUiWjnPyzpr9PdDBQapL+SQ1vefNfgCQF
uL8MTaUaHj0Ir0qLtN0NansEkBTvqdwtYLGp0xFjCrK1r2IkKEocHkqCPRz7eE5K
FkOsOYhJVwprwx1rvrE7sYD662QzGLpwQsolLAHU3y0V9xXy0ISCPbQPhH/T+dC8
g/IeotyBgdZvgCP+PMUf1s824lfnzPqyMPfRwSKpShguRs6XyYv/DwmKA60y1O4f
mGHbPC5ORGwUjqEmZ+QXPesU9ITMBo3JVfTAW67LLltqiN1tf7jrvKOFoSsIkqF8
wIxJPJ0KPgFahi53UdUysPyLu90h7Vd92yQvhOsL21x+86DjsBGkMwgkidS2pP1O
EGaUUl7hsATREgUJYTd2D3H/PSozB5X9fEiHqYdG4JN6uqLOkrlW8AE6iwxThA+B
DrMj9UTjI0nqb6WPXJDgThR0HcYfev0J44aoOGQkdLXTQU/z4DZEVDXl4EPnzsts
lHw9T3OCyBQUWSXcFWRzOoLbB6UCaOXrQTMhhM/eSEN3VSA/0EgcC+0XPUAeKW7S
xkItkNq0MGWwh+6OKdX2oYdwG6+a4ymlAUG/qMSGzaYPCafBuAio37OM/AsJ7QvA
ZlX39pp3egRDi2ys1uwM8pbhgCPvogkxVuJufGloFYGctgxGNN7f8SHUP8n48JrD
hSnUV4r6aySwS4te01gpAlgFYSu02eflpoTFZ/iCjSCNq9rsNxk3uJSoC+hMLofS
YCH/XrVNue7yaYVyeu9oIdGGTkMuYZV1bCOBnkGO7W8RTfBjrwlTR6Sk4Q7fTu2N
hy60jbNTLKYxj4D0WXRCjirQGAPYQYaoWzWFoyBP2/iwrVroF2t/EMZcplNiqLe6
3B8NZ3WuD/tRolVDD8lCrAcWE/iXloVmq4lkgb7FaZB0vPjHEnyaaPh0ZwRr2eW6
jIcOGfoVOQ6Ad/S2zQdSOLnKRFro3FeaFxIQbz80L2XhEXZ7K0wGuyBj5covht1X
XIaeC2T5Ka9WkCANZS0taJXFjmk2B4LHtM/EpWKyC5tTBfv5mixBO/qAGQBrDOyF
NJEPuVhl878ss5jPfAnceXnhZb9GEi0h+FGqFQvft1kQYrB2S1oZ5zug37r3oikB
Oo6TIVztemFZzBy5+0Ke/j+/1Xl30qYcyPbxI582iSA4roo9kdgHxA4kPrFbGA1K
OrUZWIroJKonGH2sEJTfB+yWC5pKXa09yOisuEAMMs8jOwQDT/EQUwmkyf5/vMI9
6vzfNA9vO1V9SIFs1xAna8lNgCTGbj5NnuxrFLWECJIE87nmykTChXqbdljqahtb
HokDi+fYBmgOcbvVN6BLKjTy9nXFUAdCI1HYs92C97mlhXbdxvJuI209P2+wAmVl
T3IMl3V5ihEyTz2Lavc2zPfwsvUnH+h05yBfHwZ57nKMzCjMYeZBJ6t5YvCIzSMn
u4440wnhUCPAaada5Hwgxp0FHm/M9Vl6+exKJBG3kvjBTy20iaEp7Wk9znF5v/AN
8jFtNOZd2NzR79F6v4IPLSfteI1JhXojyEemNO3yFrZfREMsN4cDnUJTx/fwcC0l
pykhWOa/gZRNv9SfFj9q6dtMy1vP3WvKnLwcGNhauhljUGeSo1DAI0oT3N9paBqU
brn91ihRrBjuu2PDap41hD+11Q0q8mtWLEY09wRdGjg1VQG9ee/s40O9qzFaRMnX
BrKuzP1d+dtM415pJoENpNcq5/ZN0qXKMG0gXEiChctJNHZnjruFgSWWD2yH7L8C
k77Da9hkaguqGRxwxcVh3YaarMa4AAs1rD15fx4fgXhLFyqy3xmhtiyga8B57irW
oH2dDKUn18CsWLYjJbiXFTT1QzS97L2qzbuwToc2W8M2MRQLIBp9aSwGcc4zUbyz
G4nFQfEWvVhVC76qkPhr4eIV80RSpdL8rGAaFryjruBOyCpr0bTu76YgX5qLspqa
10anw0aYIxLoDk5QyIMgJqlJZx0k7ErJ4K4uV1dk7qCvJ4tIQ6lrQ1fZHiR/g97w
xNyHei8ymIxEF9jN98X4e4+f94UoGwZeOL3Bvb6Pd0A0Q7N/nBzni2zggMXZSBjY
yQJrJoogtqnKYny5I00Y0JCGrVqcteXU/jei3k8pbWVgj6iwc4vOJx8ISGVLq32y
WSP/DWUevK89EjnFdOhRS5P9M3l2upQ3aPPI0ol1f6OoHPQBnmzGO7wM9Ayu7TZy
0QdlwJKXymyFpuqXA30WwlQ4g9hvOAhLY15XLB0boykfVfy17birb9a7/IHClrIb
HbZdExAaAsppqu1WCpr2Ie54+HjIhG1BW907FfA0IG9cn1RiMBPCuv8fH5Z3nVUA
pXw4g9/CCitExNymYymmHodEkLt2fq/fQAj7Iw62wtnjUT8svDuy6ejd6QlVQXlN
URnY9oF9VAeDiQSVYu/3XRnC/carsBsAfLOKDKXTgB/aNg3bYQBzljLJPY/qjPPN
UZOPVqbYei7Jb63oB7KR3IHVBOgwkNcR4lj1KfBzMYnPTqPV5LSyw0sGGOUGLCy7
pf0jh737bIZgZ93jJYGAzcOn1DrX3/ngF35jb8ejxeWNZWyShUHsNulsrEgSEPyo
xnljYds5azFF29sbUgA8DvLKpI+A7kkvs8GgoEoBgbtyfu2Z8dCSUgQJpyx4EQ9r
FdYOC78ztPZKPgMIwKAzRi3VxxyPQiWeLTwJbYCrLfNsiYfM4UT2fAINqsgiGG3C
qQYKX/z7Udjb5T1OsMMhUiAu4v4FTQueNdEbR3si4mIAcFdt4zWaLPsdRJAihaLV
Rik95AXqZuF2UTJl6AsDMtoK4OCpL6D0lIQ/7n+VsL5LCuBFqbVdZ9cncPY2Cu4j
PCVzJuGWfS+/o7EnHj70G2nweXnKjs8U7ITLlkRPWuJIBDsfTF3vXFPdulghXSrm
le3m9eQzc25XsWTL4I7NseMMyNQVPeFNXCMdltvSWAMmeTE7mNM1lnRPbSoYx7yN
EjGKe+9ztLOP0MJlORDUdFSD5xw0dKtMh3sZ1+o2kkQu0LDD7saM9IyXYU2qQTJk
z2ukkFTtk1LvQd/U757Jg8aWpWV5ACKF2B+21NPXdemKAd5Pv6raVkIYeJxy1SC/
ILwl42BB4rjBPYWRfsn+GEY8DNtDToVFOJTX5PDy7r+wOey1SvZ/a0XQqF8XO63l
Lr5YbPYzXc/MCgtuG5QAFmqRk6JaXEmCBjimJP+6mpjHrJfFg/fhmAR5x7RUwVP9
eyMzvZuVU1+f/WCXU9B6DYOLeKkNxLFobn5RfPSuV/Na+Ptriik9vhCd1X5Do3iC
/+hJ/lemP55CTfEa4wKGymcz+J8klrjy6L4CnBWRB9tdjb6MmSq2X74Ck6dCFM99
nZ7S9Dif0dr8NoqvKSaeLHSWAPx8571T+4EDMHIKHVGRPoT/QkG9CMsS/tnKGFda
QVWYfjxPpyZBrMUBua7tWx65mvkMdu2NernoIssMyJGt/duo8r/8k6M7kcIsttF2
j5kuexjc6SHXWLKTNwPH/IUoC+XNRHtUG2+psJSmmSrRQRmy3re0coweL+DVXUBx
TNE4usrGzGSH/Fd+mOoHC7P2YpPQT0hyz9diiHfTj0FfIkH7NT+DhAk2T6ZHT4o+
CQujZVJtjqqGcsNCxgYY+iDy8EN9OEbi5R8IlVBQrbudNfgr28xHmbE/bjsWtM7c
NPjXucY/YPcaqgVxK1sb/HJ6lpDwpvK843vFTKULqCqtvEnHImf1ZMK2PzWyEoNa
m/ARblmHQKHI3K0xY7onNToJYbZrNRuFi0iZi2e7b5uYH1ih61Q9OSqXroX0M4So
NtmlnSijJ6I2BbQi2cunhcP3+srDU8PdrLSmX5UCjNQskjMIpBToI5CYzE1uc8QH
cFrQZzOcaM+kQ7Xz2joP2IpYBldVq90BiJGGsZdPAPZ32LaIkDpe/WYnjtrfxRm5
bQ3oTFlyCnc90W2oo7qg/rTHrfYR0oWDjVAqjsSLvocbsokrQ/u5TWDkCNG47ezL
WT6+wVA36WsHsQ1mHQzEavfAXMPwYxpp5GJw8L/As2YxO2+sra7vrHbvXe31ObKr
3XCZS1lh3ZsNYGoCe98BdEALAVwnRfDvYuNSUn+S3lfMRvuJF039+PHcAVCuDnrh
udQtZxRrVj7wmnDRameEqiQ54Of45gyVW/it24HuhTR41PNRTpss/tKBJW0t+ndU
GcEsbncQPXPefj3RrD7KEdStm6Voe/uOd3TsqjyUEluLrEiL1QWFtA4o/vEGLNQ3
qO7sQBZ/J6PPDF0bNiUCaFws/ibukydA3ItJrBf7uuekdUtnZ3/RaQn7y4l62my0
ApG5+azeYSYe1QxUrmS2XBGWwDrHUFuWacuEYm+QmMjdGMT19ys8Wv7YwT/on2Uc
NohDNt8uxdrmbEpZefMAmXpNXCdf9gRxa2Cvn1Y8j2Kh8QyjMuRS1p491FapHf79
eZCW57ztVKcQJGXi1S7poNGmTfcONbJ4VYIaDiOjAVFwA4vgXCyQvhhHPxd59Igu
/gFBQj8XrSAmabtoMEJO8/a8XHRmgApSEx1EGzDxoDHvcC+ldwuYqzg2vq2kET9R
kRqjzcDud+/hF5OleMoXzLVviFKTzrw/3am78o/dx8QIWjO2yl3ZE2GUxQSC9gN2
tGirHyDx5Byv2DQRsXJ5CsyNAeC7kBwNfFihua7VzxB2eBYRdg9ylkp3B9z6/Ugr
947RBdV+TJ2RXWJJgDT1TpmJlWVBjw1iZTvd27xQcgP2+5vyDpUS5zO9ITUOT2Py
nV0BwRe26XkekUChbdkuXn1pbgnfEttVlczmrN/8jKIraUlBcO8ZW/+BhpM/zWfN
6FhJ5RYlTzVUS5kja+90phw4/CHmtch2Q9XxBIqyTeVxeOkfhK/KCt/VK49gjepr
QbCZwW0sARq08x6SPDwoLiS1hCk9y/griIud7L5MbKtN6vNymJecTl+fyPt032Az
NINOJ3NlibgCdeEb8FHM/fUWbTQcG70xMdUGoQdSGlfJIzvQmvjsCwWf2HPIkR4t
EBrwvqPBIDCfuz1/7GbqTJMayJVJOxCpcWshhOpiWJ0hq0CoPtfGys1tNGcMy5+n
L66eSu58R+cMsmFar1duHBkiNmCPBOsyQqTVG8jK7y1KRovejb2e4C9TOIUqxROV
z4rcP/jYZr4YYMWWKemncy8wpHfs00USmrObcp0OOdY5Nif0YnOupPxk8d45VkwE
th4sS7W3hkQMvbjsh7yVHHDQRlvlH3nUB9lyYwlEVQL3KQUhCfLbZKnqjoCfCoG+
t2NvikPBRjxeQbGS6lXuaEp6YA3ujO5wd1yWSus6ckA57xH0s5jtREj7Ta9/YlOY
RcTidGKCfhnPOcxPHhcaFcXEhA475y7zaamFtpRRxn9iuUrcfnhUA24wcurmL2pa
PWNmLjVwfV4fXX62ex9TgUTFyHiDoIwzDlJB4t4soiSU0H5GVbF7W5tZxd3oIF1C
yC1TMYtsPsTGj5QgCGCszp8/NZpkt2PDNIOdjjohP/7FCKL1HCfOvwonfNuFawc5
TXL2Vb8RUu+W/f3cZwc3PPIzqmBqyYCkLi6iDrpY+LK4s4xzKLgGKPbJdbPx43Pr
RhkH45YEQ3zlfryi5KHuKWwqQA5lNfbJprRt+lMZXuFJpkt1SatUzVaqFwcD58e3
Zrbj6mR4NxFwhyW7N6DVu+w7Ccs+Y+dc+N9Q6OtocOWk3988d0Z2gzKUK4WvfOT+
bxylfpruZXtFYR5Aig0V6ivzo6X4dwwk+BPwVkDRO3A0SNPXSYUFoGTxfevJm7b+
yRTNa5RCyPuSUXYqCpKk6Od/M39B985a6tW4rq4/bdMm3H0ds5Dat5Fi2BVCSg/w
B/ZRKhYu5icedMtP7uGnrIlEjiqx7jkctXnV5ZX+NjHLacJDAeNjPC787SEurRFf
t+PH5Ui9cGxut+XxYSG6O9jDTsBw7pk618Xbz3n5hjf5drW92K4MbICl5nV3FTBu
ZQAOeCn6biWGXTZ7mzNt8JcfbN4oNE8Aslj4HcQN8qcRmRNZU0fSCftQUSGjwJsE
HzH7VIt97RLIZ61JPOzpyS26CQvezbyKOo0ozoNPWdh/FeNMKSPAIHGBIdORVF0F
UI0UbMT3/OzwH2oMBnzf4dmy3MjEtDKm4fBT2pBuRJjGJVllwIDLpO5Ntj2Q+qww
47MFCw3gR3RMtXjh7tdw8qpYNl1I8J4O0u/dV89FZKKQVUvy7FldnZSXpanBok2U
3xZQQHJwX6XFyD3WrdyUKngmyKAX0iwcJhJD9d8fSNunXqYYwpQIaYbkJ+bM1eYp
wr80hG74dH4Ia4LGDhhXqgQJJP0hO0seLMnEe3ggXydF8ouxRO9PxFUPZXGCOXIW
J3NBuLlefW0LW8q3PTEGeCMYGV7foh2rRxaWWHhl//SCluZKBtezQckeIskT8Lfg
DuZLzbMOYfGTbcuPCEh38VFdlpAGathmI/7rzHKg0uym9iuJwCPAU4fJYKlzA1vc
lTX+LSFM5aQP/IsnxLVP7UHXNe++/N2uWqfRnPt5pqvg2aROEzrrKURLxy1vN8CU
psD2+ATgeD0a7UlBvEB8AggFKFx8Ac46S6uGwMfF5+sQv9PUjKXe5zUcmg59vgt0
yB1aD6Mb7zM7Ps1xyDlfLtjO31pYOjar9eNOroGEXTfh43LokMnCme7UZP3qgLeS
htsTby5GbhYHYAdj78hAwH9QAVC61Kv50SYG/0iDxSGdSKIFZs67IjWIc7Q6+wE3
3hJtf1Sidu/6mPpDklmJkx5HVtf4H/jddOHPMcgPr2OjB+k13kKkxi4CxrEIc28K
koHGUjgox3N0+PdPoFpfz6/VWCxXfG/ZyesnSbGHp8DuP9+RZmy509arGND8SWvl
ognaO1oGi10NPPl2vWyadavJmPTuSET+xTqA5FZAXWq76KmzFo7WaUg92kgMFwIC
zlIvzQHuUkNz/BxHpp91DGc6LOJmE/jHLM2mHbJYyoA53Ob2Do+oAMJRovtMViuY
OsBnJiVvpaBpJ06qoRP/BE3gu2Vqaws7cKQg50uG23QZ82Qj73pARWbKeD98cQ8z
yacvuHl7g+jFBPGOt5qO79xBhR9IDhOTMFoF8Iv4+XSri/oYFZGbhrFMHJ8bz87B
aIsKYi1UhNWLq3eKdPXE4y2Gw6R5r1jIRqqLjAhGjjtcQghwrEl+WgG6uV5upCQH
iFllv4TVN1tK66DWk9AxeRoxKsmY0c9V0C5JpP3Z8gPR3EMWyw+0o53QT0grT0jz
0H0xXFuQFLBGO9JJtXEgDgdUF8/YBBitkbnDsmbFslS6Nb6hpJFW8X6/ZcaYEUN/
gP8PZg1eCdJT6+MhHImaAXMYnipxEuNYnBcHbP91fXNYRskN6qFvPaYcimEF/Vde
z/w9MmFmEcNkntae84z/IcxHPbV53bten2+Yv3I9LV9LKUcpFsSaFt1ctvdwSCT1
6voIeudb5knaPc5EyaEfaykFBo0XNzviyEtWtTMdfH+004/bR5v0cR1gznDEYMze
oB11olTdcoDnPRB8+zjwj6CcHjZmqoF1jbh0S7eqbncCR2yAaL6aqunONcHnpf8Q
3TVzVSp9Dxt4n899mEmUyqO0wB+Z3X/I85az28OL/rRd96RUGlm7nPzbZr2tCneR
vX53gnrIvbdtppJAkuAVKBcR3LOamqiCIVHnMYEFDl5n6Nue5FMB7FIrsi/g5Pq+
VqD4H/3bvw6pdnlKipKX6uP+GiwHS/oCmcGOtseFSYcdnSDIQv9MAC/ZlQkLh/Mc
JbS2nim0N4jwdLDxIsEYMz0/87J8xeLf29kqegujJZWfH1sljAplv+ZUvLcOSk8F
m2qFyI31a4Ny62P9kIeN/S50WB54Fd/3Vu1JMjed37/MbeK/qo9uoNU4aA7Vuihb
6PeWxqL4iYMsDaAbImDbUAve7KohxiYNZM3s21oJu1XSMXOsLTR7JCtIcAHKESGO
syVzK3IyF7TsNNSJvwGgE+gpq8EwXkN22P0u1LwCs1kKCVW1a8ankOrmd9Tzw8wW
/IgPBP3e+t3wyCCb2uQdvZc0MKbJlqWxpkfLs4HGvrCyF3OAQNjZdeCg9uJZJt96
Op84hrwK0XslW/JdWNQjKyF1H4eAKgBin4qmxfcfZ0mdJx50gxQNo+kQxmB+mHtJ
1WWBAXrx5tzGGw6nsg4hHInq+ItTO/e1tuTNdxXFn/PjvaZ27r80SFEWw73d6VLv
H1FILCam/8cae/ABycOB8OBR8xw2yjo+s0MkDKgz91q+GSo2gANhAKtSPngIyNy4
eed+EJ9xsJpi0rLWU47I/ibcgM41ooEuopSPeXtDEopVri4TA6jKRWQDaLsq7M4w
pKNzx62jhgRDzW+I0IGidWcF/WWFzXYwuxLPv3TqjEPYYgZhfQtmDQpFfO31Kzj/
MtzRL9QguIQ1GvOc2Nwxf2f+fBD7BxrQ98O3Yvcwzp+oWs5twtBtrPbYMWceDzts
ITftFRZfLEy9j2TMtngxd0FJSi8x3gDP5uI5vqSvEZACDlTux677QMT3wCGg8qOb
RgANl0d6mPE2q/dNJzAKtpiVd9feSFPUmWUNeG6WXk0SGq1uVHDWszKupLTuJ+DE
8s/Mj6T1KFIJsq296tna05re4mtApcz3EzqZpNP1bb5h6HQyQbRhWEftw1tco0+e
rihHBkUDiwaFYkWoStWGAVCm6aHdhWnXy0uEFuVpCOMiwvmN8grBUjfe9+g2SR0S
g6zIm2H2YU1PP1s8nKa9JKyhOt2NZjWRqG0GR4jY0KuqfJqYQ7Bq22e0rlQy7UwX
NXnxkdcwyJPSr/frUrwyo3LaKnAblkc3MExngr8hGowLw5YYhkJdWf50xzgRZO2j
TJNdPDx+KPrwulkVkRAzWTRdDUmGloynU6JjWyNizSz1oseHrpwu2h+8ZqXvAa6P
9/y9w1lLxR/AJDe3AnqmoIQ5Ib0DXr9XNCikeSMtVDhZWyITBpmkd3sqKz/ZD+ZX
CM9JxzutiZjpe73cu/Ajqgr64fpYkDIX2zXmjcKCg8CPnNgK2LLxHU9hLSzcjQBU
kt83R67/pSo6nIaUNHfyqBAWtiAIRJkTaHQ9eHro4PGfpkBZ2HDRHnQG4aum9/7F
VDi0w2NdRVa2TBoZtuL3EaOz/xJTTPbcF5x0nruov16BCslE4zW1qlal8X/E5f9D
oInHH6AZQQvY2Z+esYhbcTjzwCSvlSrGqB2aPZ/ABXI7ivLWmqoxr5EsvOenAd3g
KOssp67LFoEB5KhV+WgfUaX+M9E5uBwyy7Y81aDv0LJ1wSJECy/u/iQmoO4GjHxI
2pAMhgTPE9Zj2qW7/PhTkQOX/oehLCP1ThjlgsBz+5hjN6EauudvM93C2I7UROFX
eqm8SJme5jHc/zfh5qzyK0bBCbTvm4UdrV6XdEVqPh/HJVzSCuYIAxrQIS1T0zLC
1L8z3Gx/dKfOPOrEPHXMLYuJd4clbecRKQDu6gIdP6GCsqLXW6wvMapqwGGziSZh
U4YJJEeoPQFduVpGMmiI+grnhdM4i6QTnvaXNEAUe7JpWbWGYn8xwzc9xOiVBqvV
Wipv3GNZdJRy8/pz6Ue5UuoZsUSKkdLfMb46tJWrj9uMdNTdGWGdZGeVRH7GOVr2
GIkKpIdDlFiaOhDxXW0WWsIMIVc3fgHlPrFQJjSlJVGew6rB5GIH1dOw2/ViExsI
M1ld/ojOOist1dbyxtWFdj1KxR27vMZy8cxU9E6IYhOwnTo6Z881RY59CCPKIuZB
IwEdSViqtsJginQqz1a/n8Z3jDl/uFidJnatW4qn4oxMrMw1O8fJL66HC8sO32iH
CnLqddG61iI8qBjmFtFQeeiACHJBErI8FvGeEwKmEejy6FrtPk3+rbgsovN7QLtb
FVxArJhX7Bjgdr8uOhQjoOwT8HHNaODSatiAYcKZkZaDfsfijcphyMsWxd/uovRd
HRPWJimgV5T7tyL5zmCH+rHmGi8uLlywEjfkynt+xVGKMSX9atmN9lY3p7H2UiZD
UculqLOEKT+GwAs7l3KARae/5FdchYBE/ZyFLJTAhuTcH5zyAyQYOYVmeGkPHr4q
O2hQyrxX09FdiO40eXk6TNs9pxXEg7t6jTOJzq8I9M6Wak2JqhF49jFvwlxIPGcB
hAMR8pRpim3FVfGvlUMDPlXUvEmmpA+/rATwVkUaRuF7jDxoYUvpSX8iwtLWve0i
FlcmdVkVPOgsgW0eJemZvEsXkaYOZB2IQt0ZqyIc/J3xrKm9gb4hl6f4vF57CoMJ
y0be5A0wIC4VX6/RR4WFdMGh6k2rxv0anlywn2k/LVOvHEOtUaFeRCBd7nbwN+fw
lZ1tMeNPEMRZQVSMLDelYMnJtDukBB0SCdv/IzEts4EznAu5SYRPBj8ZSRm+E5p4
1e+DFwhH2Jdo7IFuyvxQFftorotXeS9NgskkClvlziztfMppBQQGDA1R4GL0VEQM
XCXBGWYdXNIAC4s0I0DTjRchKzHN1iP0VNAaOqDQ9SobIieCRklHanIQTuJqdN5R
VPJERrlSgECdYaPvyjl2ZPkNmrJutL7cWPvGjMTF1ILuBd07g051abQDYjof+4Ks
ujl2yqtPGfaL1xI8gxfrzyJLhlIvD+CZQ+n6X0NL4GKNK2CozjR61r0/lpZKnRTn
lfHaSwHfV08IAo+TWHkESbf8XpRqMW7hHbN0Sf4GO23fEDhwhOY817uMaVV1mCA/
QFIWJXNMoz1mRel/n1xuO34H+MCU9mfuGbdvEfJEhkp3zDLmWDKwZDzRS1Ki+T6m
d8zPWoOWNDZvKZDpjACbbRS528NQEjRyMm/xM0hzm8g8OplhgDiPWWZByOWc+1xI
3l4XXrXwLFsWu7gItQ/Hv9YcPZhLLmqbEWAc60F8jXW+wEPCs8CnjFOFDoJi9ilo
MVJ5wxha5sNjU4F1EpE0Y5Pdsx+QYrSQQhbNntnQpwTSLpfmFwYOTfbcjH84mrw4
BnMlAZZpKmoL4jMBXejk/bLcu2ah9aXZjAaytRbcHsmGGWObkbTDDuRSVcDQs3Ja
n4dUss4P6IGoiR2yValu0GC3bcZ4RIaFKO25AYfZurSbIfzxuOemA0gF2YXZcywq
n0GG6gDX0bhyQJdOISq7E4CHlkvw2zV4O44BxHjHo5Q9cmNuzS3DLNGVXHBGE2z7
oD1PMlzUiF+aCJOO0aXk4NzOF4PGNHzHNntgwLZKRGlPSjps1URRQdpLlBflA7ww
KK2s4EXZL3uqvKfZratczKbAtrbR0PF/tfeNH9GVJKc7IflEXz180YTfkuCsGViZ
993GpJyw3UNYnRKSn/eJw2TDQKJtw3XbRshtsAaji7pXi8BNtzpf3bCRQGmQMYyH
Gh3qGg8sHQF5qFTjdV1P5+O2P57dLYGxfj2FMovBalq4a9/sofqqRdxE2tQI5eef
Z4QEzpjc766OzUdDZpwjffxXGVCiRM43647G6kLpHlHKFSCH4TNd4mFbSaV31tpH
+ctvh3aXFVBFb/B2r7NujaqCod+LmMulpwokFPNvneQXjENxoG3992e3buuTmbnm
iz/NCbpKUgALKIbakugRKk3V64o2fe5ev2oZ6czsFDwwyyGWjmCK45bjgDa2KLKw
UYoJqfeEWBhO1/CMu2+ptNJuNkkAl5rFiOL+ENG8IYYhMT9u06RZZumnrVdYU22n
HYQ4Wbd3kTnet5ctMcObPhQrX+1kZJ7IKtMLrrxC9YU1GKjcZYP+Y7iN285xPgZQ
xUrVWadVhG9DCZIujEkLLigQs93KJk+NaGKdXDirEMtZsM0AiFg9ucErxXlPfGmD
4EZ2HlqqSG0b5Jhz9yJedeun1FPimwgRgVsPoDgOknyspxaSUn2v0ZJYdI40P6eW
Xh0DdUId1IHYAHkd0KJkrAQ2BF3hTLSXOi99Jy7rK2ZoFVpgv8AlLAm8ZooUc6KS
PiVl7g9mD4swtavnzqq0vsk9iz5XasJo+T1dYChruifh3/mB2JnGpj5VzkXj8FZe
PylXRuYrp4uOK5AxF2l9B6Jv29siFQ+TA1n9+zU2CR3AabqyS4CpS8DnA3iyJ8zK
QptDNqqmf7YKxOv21ooCqQUp4mMuVxX4TIPYuwGaMpF42pWQoJOkXgQ/klBftnSW
2j2HFoUfSDPLHYhUDT5VE3dS27erBD4gvbGHDsomyyOdJrhs2seJnznLtf4VmdY6
Te+2CdO8E2dsbYq2DRAjcAMBsCQMORBCiiN56FvhCg+kp6xAKn5XZ+8tc627tB9Y
3+xNdSH/hv2xweADiRWyhCSl72W5pe3xUlQk5bIprRZM2BUOBVEsoIIA5lWK9vxt
N5WsqqMyl37fOvOvSGiSfd81wJpw0yyPUnfCmu4jb2aN+QZLFGUS7FwjDEx4QSh0
EbaNRIrlcbYGSavVzUo+a1qbMDBY9FOmbvu6BUKW4M97QgEsRmktwZhMK/nyDdTk
Msc1lS6P3bMJmM+7iGXb2utTpEKGQUn6qNVAWn/AcOo0CfmpyV2/4e3xIKHiS57i
ftgrJQurAmGjA5/qsdQFiJnPeA7xQejj5ig8QN1a0DReFJWnnA5KX41dvDHMdDa+
IWsOOU4+0AXU7CkDVQz5IR1eKcVyyGclkTRdYl29I7WUUHWPYMFuIk9ZgZ4tC1Vr
zpifsjDl45aG+pkjn3P3ZugY8IOIc6EEaSX5wwBH39TYUvq3pW8dNIcnMp2SHwAU
I/Qr6xkCk72CtOtEtBHQSpFiR2ZvP1CBN/hUpunQWfUhh7wXUwQxX6O6MFubLL+E
BiD4fO3jYky4gFWPiioDJ0D22APdw4tMr8ULNYFt3czi7RlUhYlz46CyQuZfW40b
slp3HtOV/SjKA0U1KkqSm+w2T/NIFVEcTj9rmq288+uJzojLU2MejHJo+YXBBlZG
3f4onrtL85r/o00m74rGWiE6UrPWIErDRAJtck2DT5LMT8n3OSHli6Yjem9098M+
zRLm68Cv/DMJUuw79oDce488qkoDp3Tm77D5RJsAfO5UotncGHwvheeVfjOsxhQq
KMYTxy9TJw/mpKTiS3Ha3EgqWy3yxwj16Db2go33BLGV4WzoueoSYx+H1juXCpZ3
9GJwrcYLd00So4ozWcF5sY2HsszNHfIRPnUC23yp7qEN2aQ0aKD4k6hKHL4J74Qq
ddcoqVG1uaZvwYp9Hs2P7OyV80JPn4GNFf08SxIqR9+2JQnzx9szl25Lt2Whj4OV
/7LvWp23kSSbhYG4Sv/9L28BclXTLKFvJzzWsvxlRIp2KigPreccmg2Q0Mpww85d
XmtTmP3D3+vfzIIo2Gcz1N6p9nMDXebA/Cq2+Ctf4tvpJnwxcATZ4F+1NMwROErM
XgtKZFnJdohnE8XudJuRG1sTFNqiaFuapRtKk68PoQ6j4WikEe+rXmJWSGLLPAX2
GaALtfjnvX0mUBeKmWBetILeYR4Lvy9Tzmtz4o4h4lFKHFm5nCFCocM8P9x9DHL5
SOVB1ifqdA9TuMdvCLnmehw1fXUE6NzTSdMPeK0P7HQq4l0njQ1wE6Dq2sdS277A
9Fb48shcx197LpRQ+PcEoXGyXpXL1xYK6d1aRK3KjCRsSULVvsl2P67wJTPPJ2iV
mDA1w1mwXpkjQ+tF1zqrB9RJHtADbc89FfzikpHWB5GYXZqIstSw/3tU3bWYY28T
wgYFthOqlq94d3+pxgID150gDFuar2sEx0Tl4Hs6CWCLp+lb4LGe677OAIRj7M1Y
9j3g10DOEpJ2Yz4oFLWzKAzl0SsYBRgsIYZPvzQDcXT1SXO/Aas9kcXDrtSdFi+6
5e1Mq6pB+uvUQmhFOISJy57rtrv8fy8R+31kKOiqE8YuX6kE7NZHAZxe49fqyI12
YEKonp0hJwu+A6dNbRf8Zg+vwiO/TEwvMhZ3rTiva7CqRzuU7lttx4oTBijowiUN
78QsqrdR3eiJ+BujuZbbvRJRcZQiUmZoOOR8mT3rQvD6qAzEMWGinNYf3OTFb/91
diCco+pWdi4gqODGaXXNdj6biLrs+JnHHPiEeGuH1z97NgEQVJQYJJ5ctxce4w9Q
GqjJiXXnzmc3cqlQajuTCNN4GLtHUmKy86HJ9+ywUHnZnMKTnH78J8k8RS4m+Z27
pvVfZyMDLXBPtypueRbQ03owNla2Rs37TlRJaFcD40OrWHZrgPQA318MiT2rPzyG
FQTfsW4/nAUIvujZg3u9pUN52jbK5ipIkkCPQVX3ONTQA0O7b3TSyErLqXgITlvE
A2psu8/o+J/kGiimsv7i0nU+vz4WMY5MYvDL3q0yt3tIG2urZ9BPTH0d7Z9ZrRg8
DgkaQEL5ZzCUNgW8zoWOUMuISCkiBIBPIkQjiNH7WUt7AuFOtj90iYb1lKRoVGo1
pDPtfE//k5SA8X6hFA7WiBo3icppx6QeKv5V6hFAgi4hbSIhxgGG1Fp9J+SZRLgs
VbbUbFhVi31lnAPuUrSKaWK/RJidIqR+aVGzcKsQvhC8VthvyztlHcKh+kv3Rd/Q
SujveWR2532UdvWIcy2Pf49eBas1w0B09jOnX3iHBtSe8uqXijgEtFlyum9A+Vb+
fVxCLmH8I9HVVZDnQoDVjZgjYd3ztcytKHHd/MkQKrTxEkAU95faih8HDEkWo4ov
jSopOKSPxNeKbgRgFpp59tOay5PeZL1NXqPlUJ4N5GHjj4lcLjaM9RQ/3sM5aekN
MOZcAtdgjXetN3Y9bSdh35hrv5dvtp+6j1iVWf/bnANpLmf205540cb8LIVNKsSK
ZGcoiXCQzLeNW+23mKCkzV+LCaNj9LWvueUm+En9pKZN6GqJNYnRj0nEeAa2Shso
yZk1XAwkmOV0BWZnopA6nyVgoSONgddaGfkKmLsdXjYuguYlCJKpNj4qFL+3332e
ouLAOSVsycnxCs0tmI39c4UxXdD4P2cuV6yq+MEY+exLpmH8y3KLwlUy6VZkMPft
JLeFRgA3tBF7cNYQF0ESsfERjB/LtuNZQp6GiI4z8MNefpMn3ZoyeyZO9OCWSFC+
1bdD5Yu5ecQlY+oi5/un/RAVX662D7QfyCMKh2LA02UNZCkeLxHAGTkr4hL3BKH3
FSk/ru2+98dT9FvQrl6/Xp20Xib0B23k9awX9MmE4CHLIUzn21b1vkiWBNh/kA/w
jffsfo+tef1ZNLrG44j50F4vzKGPjEc1AWu12hTfUjBkLeT/20BK/FvX7V/doVPl
aWprNjH+jn06NrDSpTcuSDGOCnPPQAzpC6CZcodjdiQBuGo7Q4osbS/rbF/WRLze
NCOdLj6y3FakljCKcG80YF0/lDi8WB2FgtAHacxfnqT2MfciFSIrVbvoc1X+bDAQ
UYIW2VIX0yGIBtBRAHCBWv/UP2iTg7cyJz8rXHQvx8g7GtvlOhudWCV7wl4u2/ag
SdR0d/J9SswfLtpqza69Z/VUbyJf29+TpzvLJl2ApwlZYQWvk6kW0avGtyDNA07h
X8yhZedi8bb/JkUkYWmZAJhVhs7+xJ4WBai6Z8EeJSgtnsDTmyTRCp9j91odQaur
fqDdb7ZytiQDF1mwY41QGjuxH0DN8moPBw5A6q4NkYGEiMqcNSmV6eB+UZ1qg0qp
zodvwRAimTV/5CQiizFn2Re6KViwwArclkukDjm76Gkr/YQVrSGc9n3611nsMZfu
5x3Xfsg+9kN2VQKDQ+t7iYopHLjRheBf3PhGY7n/4sw4UP2oYCGlEIek/tAVsM1T
q5ZS4rD5J83r4XknDB7u5/vwNYCfxfga53v6rzioYgJBMoL3+oIdqpw/nIdmT4hv
PyTeFm517o5wfTui3+o/g6u1SHWRoPzpFlXETg42vAZAvao08IvcJlaCZxXA6LHe
CU+6qVpI23E0SIjMiFj7ynsR7bGZRVxpPU6IoHeX7KqSI6TgPdRdi/w9azofw5EH
mAb+yDabq7cbVuXdgQyOFaZzBKAys876jrNOu3ySLYd0U+TB0V06uxeJWfZkt5bs
a2xnJ0NvBr6RWH+fbqaJRG/nrbXZC+WPNErRWk/9xGqfcdv/osPrZxGoj0w/AmMk
MnlrInGNUXuD/GgOP/AUPFDXIBpvZIkWr2YrVV/XsgE3tNSwnq2v+rGvdlgaaLbp
Qw4lt0MuVO24zdGH6x4oDwemMe2+cDGdHh/7wIn7OqY7eByqI558dw+AdXnYRSGP
HtQ8pmVQ2X4nIxaUBYg/tgDLs8osc3S41EOGApmecNQ1Hdx6pZhGDNxvQuAVffoE
ck0Q5+K1u5PmhuiqJoScNb1S7DMMNktoKXMFuCHiYCjfYgR7nBPZDRwM8EPvtLYb
pN/FPNBdoU2PEcInCOWXR6pMlYVFfDidESoN81NkW6A8gp4Wqz3wpB+63A4o5w4V
XKcvcjqSl2FB2+S42d6UvSMHngdHAmu323vByVSRSf9TO3PLp3UBfzGu0a5rOzrY
yvFS05CC+of8ikoPN8ELFXWVTXAG4BmyNo3ks6UylMY9niyVXxpy61F+Q2xtmEiw
De0z2msN9dcBoxi+RC/WnO3YD4Oy5moPa0xrSjXY2OKoNTZw2U33geAdBENpk1Jx
153v0TNHiYUhXiCW3zZE2VBMb6ufXu24+pq/aUyvQfcH+8aVAY8O/bxxGscFX2fc
OTVRskcNpt5s3J81GOBrTAyKhGvAYZZIbECEK1GVWykP0eADpu0SWYin0S1Z70PI
zc5f+GbyolkODMQvYNMdRp+KLocRJF9Tj+FozF07ZqzJ/gNUyX6dRVsSrjl6363c
0mDNPriI25fMuGZGowtiGf7YDe+4iq3Q96wulqJmzPH44gTst/bxpMIuy0HN5QMv
DudtchQZQlEO68KsmQhNdzXQzRl20GjUsatZHBmfRUtCH9NPHGmfD5+8y4u2v1Gv
h23RwFpACzxsZmqhwr1fR6Wp9GJGWxBHhmnvt9p8Z5PcZ6DmrNw14s+KT5GICR1G
Ty1s4fPq0pt2ycRVW6zWPxd2tDe7qt37rdlNZGm2NYEFcSqneEl5VX5sYEOeafuo
0wRwUk0/YDjz/+IgyEtu4KdJEQMUaPk4yGTJNUhCfO3ADOjMqW8werqu+w/+TOF/
TVzX/YhEvkoTnfD3R2aYJsbGyJ9vZOWaKEhWb4sWjF8ZB2ksAlxBJb0MM1m50inA
MR3cxe1F/7STtHE/k5s4JRFkWej+Ok7zvVBxv8vDgjyU09hOCh+kRa47gu4+u+He
1V9vlbKQaw2YzdpKoswuvKPVhm1s1HfS6gcYJnB1Ua06GW7Etw/CcQ3Pp8HqZyUM
b21vKaWAbA/Osx9pu59oRU8se18Pu7xvOCMb5+Q5b3JkC052RywsigzoZMJQmG71
J1buTZWWQIAqCx45yzvl/AQUDOMyT2fr9uuRt2Jz4Niblj2+YGIFn5KbXK68zW0e
A0wO/pTZ9PZOHTcK6Bs5gu0ggLLmBcMjnCxXh1dLX4fqJKsiAQ6c2g4V0kwT2Oyn
xqCnJVE/1XqM6EeIZvc1RGjofwVFlbZMvP+cIdSNf3db1LMC33lDhHoqOusDqX3r
RIfROcCjp1Hq7j4HSYJsm7PWXa+Cc1BG8SvR77yTrfDBFH8inF3Bg6c92WsEEylW
3tNEDQXMZYLLBoOk6DT5EXrkjGfCzEMV6BZgThT8Ug2oEKvDqNGMjNC6fLrNB0CJ
GMpyCiXMhLgPd7LslVctbkB26DivURWmMstyLlFEr7LNWxVnO8rNprSE6PLrktzN
oTuMvolnMeidZJRW5K9PMsNRyEymy9al8n1elYFQ7PGx+1gTofqX7M1CiK9tiCqY
Sr4mdymDeR4qeOCO8fITo7z6CQZgAT4WTh5pK6E0x2xcRF3CKR6RL3kccFAOuQUq
rNaNTTj2TxVsH3QZ620xDc/GowZxCQ8CFRyoCR79FTWyxjEfe/GlbkZKsaGyeSvt
sWcsW4yj1StppUDN2ml0Hv8AYCAkDaEVNUJmC44jCaZBugNxbgcRV3TQjrMsXy+s
lKlKVGNxYskL97209z2BeeZ/P3cczWA7n5hE9FmEI7lic3n4RJ6FyBbp93xavn8p
GCzSKWa10BiYlbo1ydsfqr8cdmXFWh+E8NTT8pe6QaC8DwfX8aRRKw890xTEmUmG
Zj+3Xk/HVVR8UIw/brs2xv4UHEktz/nck97/0Mo9yFf8e/R/u08vi6P7AfWeA/Ib
IVgeCEcSscbVmA6V3BJMlo9ahC4GjLc2Gf1kzHcw1mCtGcMy5doaMl9SNhTY/mwv
Vq41+4xpfpgFx65T7vtQxpDWVwOwCz37vUsB0NLUF3yZmozjSgP4nbE78tV3ATnx
qVGSMgKZEdYIDjABEDjuWCbwJo7Vbe890w/2Lc/Sn5V2OLV7U3E/rM8b9m4zs3j9
RSdNfwERPy7LpkqVUOrI9JRK+wjuXT48BlOt0ZN/IjSEeWCC66dVM0bpWfJd7Z8U
5UVeQ1ocL0DQvrSZTYMnZ78MD9ixiSv+OsUiG7vLwoaJZ/icDMIPY15r+SCOCnwT
B+P6o0vEHn9zJqwlE5wQTcDp1IC+YmAu75d7XFGzoyRQnJNNztEHtKLyL5X5pV++
RFsOxB9Ha4Yn1ab+LC/7kwGnMGX5anQsGpNkRWxI1QbVG1dz7nJJuh0McsHU3DMe
q1CbTQh6E1WRGRV1L3bpswQQZH3UJ6qhiYA5WLpIsVJHgU3oMnieCkFP0whOwZsr
/U0XrE0S2uRbD9Dl9x9KhLzBeQqAZJ27r9Z4K9P/T6zejWUV8OgQiGwtMAzIObt3
g9gdm2re7OtfCOgsT542KESlbBie402JcEQilN1+lyeLKsjeOKA5H3MSdvN/NzTj
v5zA5glLMA3CUoc40UITLWGB+1Jnw6FpebzW7aTQsAp3wsacBrYf2btbV8tYCfKq
sxvdJFC5wKBkhaVIamaV3eMmVN7bjmI/ZL2N2vLKR/PlQ5IseZN3/QucK7vrumR0
9c7kw5Wu/aIzhQHTAEL/GJgeFG0yAz0JPLoPtAh0wyl0lGmdGGJxmIObmR1yUSN2
Yt3smej5Zzg/Qdwv/7SPu+IVVzPTH1sv8pgF+hvnWoLTriW1WcDX1d7uyq5BKmpe
VJkCiZ43bwGBpIzSY1PBcjV7lhoNdQiw7hdL+rzP290xQ5cNi+Ul4ApDodnuQ1po
GHZRFyg27YkzG37IV6BetyTaJxXbvPlXiZv1rkXL+IK/PgX+67IKRLNxhmAhpnlL
eJNfAgAOQAkhKwPM5vTt90l6gwiNLmfq7wjcJQ8voekfYMeWLIJPxvL/po4iJA8b
+e1ek7l8TmGmUzvzRiMtxgo+UTaOgtlujOpGx+sRirAFd4WSPkLQ1dyWut53K4p1
p+gVHe+fLCVpe8mvhtYZOA4YAKIlEKMgDwD6jxH6iA7BwCzWm1z7vC8oTnyLeIW4
mmAapUgZPzTJe/3BZhM5hCb5rZgntYC50jusMcwBIli70ej7aM+8kLC572JO1xQq
++v03N6TdS7xVFPnspUBJgfWSt1Eg76S5Ti8PzUR4EPFeNz7AIAHRtYEcp4PICo9
VpfR1zT+1sKXxxPc3bBmdLeuZei3HT+f111XD57wEVo0VnZO4JvKl+iEdLred6qh
Wq4fg8aiLJOEQQ1cY/1qM6Xrir8ACYPXqvSFlCSVBG+/TNJ5zyI9+vC312NozcQf
gp4eqIn8qlkDf+40zESahqpwark8nwpnVdSketf+GFmt4338om7dVkle1/elWyWW
yiLuTj0Ifn4pIeWtfYV7lEuqvns0mWDJqwvRYcy8dWRmEKlTq7XdqaL8mazotI+A
NzweZuLx4zbtDompndnkw467aUpYIDr1H8hUR1c2CpCicfmqnk9XxbS9gFXkSbJb
RZ9PD1mrkWENSXnV0voRwUvJ+iCiZ7w+4lSGcA5moY7nVAzlXQg5HmEUHA24u+7w
dodxlKyUyKBD0DB535qCcctmdbv0ynBBXusMe4MpdyPn/vpTVD6WJ/VgUnGwAVCk
ElTOowqV+oakhBUyy/j/FWMVgbWr7eN4eTkynlsQNV+kUEtttcQluPjqeiBr4Jfw
8IfEVxIKQVXwk+6eoKkVJVijVziWYxM/kceobEkwu12zi6Pbs6VOU2VpK2kF7JRt
zih+Pbq9czh/YtJS3+J9hR4uXR3UzST0jyzgvADYZn3SZ+4hXPIckPNt9gXjCzty
eM7vUh7gC6iASykf28JAoYRx06jbU9qQt8vVIo57kFvkjaUPQ8xod0uaWejRloPJ
V4QYqRnuuDEzFFiU3jWb7Puev/7tyoRC9fMqolt+EIHGpvAJO++BXcdSTvHYKY2w
2iUKgIUAuNWBtvAhnB1xsA/guhbZnY4tFMjrHZuJwjOfDZyjNC6PdY57PJsaQeiH
wHcgeOQmVXv+DW3+Cw2lZj28jv/0atw3k3j5+Xvrd/vW/TKAU3a06LsxHrp/Tfzf
Clh77stJNXmtoi+d1dOMfzxt14dwK8GE5OWFSllNedq0RQ3pj3/s6HLt5oV3d2gm
WAujvR5reyVFXoaaP4Oq/HpgRUMyozQWXCcvX7XbUEMxL2w7pIfcohXBkP1kQ4zQ
bRPA3Pn6ryUoiEoiDj6Lkv5jOowAbP6lefIxkFFWnVNr3M6GPsRyuCXY6mYxuj3K
cKhlYR9ep02/6WCreXgQJ7s1xAhgx0FIm6j3rsIcrIQJiYxjY6Esag9NiqinPZKk
PK7kzD+rwe7qVpG7K3jcSTRmB9KAIgXFbKM9/233sw+e3+jg66O724dDLmCVwI42
LJJSkY+PZQiLlmMBlNA6rrZq8MsTRO4qa0/LC2d3UE7KNmRHtj4nANkcEALoWsiU
/RpnHcXvpnmFcksgCdsm2fNUv52ll1ZmlPGL/oHVLXjORNQEYr1ga+WVvOp7/q46
UT+0Yyq9xIGia6SB6F/7WGjmwJQzmxHdX20ew9QYywNKZMN+AOrz+3ysfUSP4BHD
EKWOjCLaaYEvHkMCwciAKwJK3JtlRnjVC+s3Sqah4jQaJjks5MvFTWeHFWV/sAKN
YNRtSouOgcRgd44BvPtUE+cZvg9sXTYMm45isBcrwxIe6KFUetgTl4hOMuyOKTpk
PHun5pAHs6q4KmFKifBdcRewQIIUk2U1zacIsjeMGEeVILedVF15Qsx3sp+gAsWs
aT4KmXzKh3pOWHDLDs8En1iTt6MbJZdM9q8jIR3HHgAJaenlzfT+lzcWTYqPFDgA
xuUE5wXD7ut7yOJPa8Auz1Uwj6oEwByoIFn+THrJfZXetur8u6GPD2FeBKH0qzgV
V+17nK1iywP/bcQo5ZzerLlN29vJ6nxZ0EXONdRcXGd6PvuyJ7Syws5E7B+7IWeH
WcOMtqUqQs/CEPtTdp1B50RfQf0SHJLbqcqFaQcUg/bV5HHuME0otFRhPYv6aJTb
bnmvXvci0PdNEo02iIdIzhDY6atk2HS1SyJEbXBJbAqkmUFGIhOLOrA9djHNa8vK
KMTHIoTgq/ydHoReYN1pgpYCnzDYxBI91lo0V49jMD4dLLXuYNBA8gHU/coGyQxe
4C8UAFu0XUFzS4cOIsubLoKY5NEtPPjDboPGvJ9hildiIuNlFePmvIUkL1KjezNT
Pj93PEoQhiL1q3DPYKLDtJuSpPQnT+tkq9THh3wuTSkVV/oSRtXXUG2XsHBTJLeN
Rs5WUWcQUPN03aUI3K4xCDxVa5sAlM8gPXGV7AKRJ+C/oMrXIvAoLGnpJON/d8OJ
H6z/wEy0govj2SFrxy4YTYZjRGc2BxPPvfTy/WvWIkM5od9RRBQvgtIuYEIZCNf8
c0Qq4/PMCaD3JGxMnUg7oB9x6lh5zEWqHJCDO7zNaezxOwBx/TiASnZbSdPhX0dB
T3zPv7k9LUik7bNIfMoz4XVdPC7DvxpowizhCbUQwyOUrcCYvsfo2Zarr0DjgKK6
Pt48QAy8PTGKMTBoGxdSiPyyvA+gHvyMQvLlGNjNHRMz64GElZV8MZvCyY5r6nuo
CVHmJSQkgrdvsxYf+L/kyDVlaLF3x2SRkAMAf/NX+ZtNSDRV7O3O6fHVqZ3TFwDE
WJ7cFzF3I8Fn2gdLygq1HML2/UxlXqnnWGpeArFujgL+AhkAkwP30YbW/8vh9O9L
72ZncSjEjNQhG13AC3sE7nz13CZMuwMZ2Ta5aRZL3sRh2iPKVBBHcgc4GRChl3Sw
lDDollf95vhxEe8VTDbOWNWhj+0qBVzK6sHW2vcKEKhb9XlbbIRWTeqvOcmUpc4e
EVCA+L44D/AHnBLPUOtS/1C1qs3ETbIb3BQCXucXrBz8RI8wBke36vuA8LYeoGym
iISwzTK3apFdQKsRQBZ6iL8ehPfW5truqHHmkV9qK5hMPCaDwdLenHZ0jHQILbI+
3UgifuVXAPNw2igHnMmg/HyiD3c0ICjfDlQMFNkTQuhGoyZvrfI65acCEk6BTq6U
YJ88RFarSgX/977zQs+M13fPZzz8bcFRjjudDtxlHu0t6VXojLvytQ5ZjAggMW3o
JDM73XQYziJJe1PumJr+bCKzlaPqvvaFfjY3MqfpVRiHXWsoJACzlNAMNuKQ4NJM
zM4pArmOsc8m19wP03LP9bqBT4kZGCm9iQ3ae72Q7waQQH7acvflLW7TCBUpQo8p
nVNPTG2AVJNY/buFLu7VbeE9hKKraaKQZr4SU4P43HK3+nxfijoCVQvy3PFel2ZE
p7V7kDkrAZBaie/tV2oehSty0SahAdoj5WCnDnWiyF8c1FQURzT9OZL+uHgoihih
C8wRPmosBgP0qgXxHYRwqUmeUuEkRav+dofIuY0WwO5udioSXW3af1mkvHP5+SoV
gi7C40cBY/1oAyvWzTwToKdEjL6wN1uDFBD1oYvXdron5evj2J/UKX23T7vPFWQW
rkgnxhPaNXNKBQvH7uHl4bxIZOhgbQoNRZPSBwaguUVlH9zffTNK+XtkgOp7YApE
KD6PgKRO5GdJ5vJIy4b+tN7YYwg44lLIwM4JLCkqN4eVP5/3D2+SeTxPkRSM4xiW
gpCeO8XvzXAxomKd7kqO6aKb0EOHeczqQxaNsy1jh5uXndhEhmptUPkK24Z87mLY
1fpeepskK+bX3gFKwfUH0mVciLieY8hlwyI86dnqQ8eKNSDdDSZhwP4Ysr2dw1tP
mG+Hxiu9v0+Lknedi36XXSUs+4ESsQPtolaHcxgIWoQwJTRdGvWe0ln+ViLXqAlc
4hQJSDL8+abGQlhnuD4x1m9GTMnuOS7CtOYDXcXLE8V1/Xi5oUiPUjbIShLQ74Rt
wLICV3PmwRvQVBZJTGrpI7l3iRGOddfsnRSZnWDGqXrK0okVAA15KRap3sBoMe/6
38XAIITn7i0AdB3qv37j2QdS1/pLuMuZUdUc3vKEsyd+F0W+6vWUZ34n+jhu6zaP
WoE4ba+Bsm/tCERba7mnlEGXv3A9tm+r0rWgeLmWLpZsMMYTkbuydrVEMxjpBkWS
+GBnS3JtPwAq7xJAMtZbQReSH0uCqxpNZC32TiKG0tAmz+9DZLNnuAAy1IPUk38+
3ZfR1/pkHoQeDY8vfCnaNvFvW+t9kRoYDm6kyYO3ICnkEKTFjgBrBt9jWUEnKk9M
5Fa2uwVRd9YvYdNUOlKHyP3grOTAvfzhLQRd1ID16o2IJpuYSRFvw9Vn024GBf1O
wt0n14g/niHn+5CGHfVLmP/Iw/kWcBzZkvKvzwyZle9VYmESBXW5S/+stGj12Mix
VC0WgEw96qhNfBTegX6vRKp9iybGpNpx6+bDFY9iD7lbkqjm9ukzQubQbi7Wp4CE
Gj6wvl+YYsIRtN9PAEk3wILdksAmmbZ1XeKCxvCO+3J4dgRi0KqEzAzd59qoivHk
oilZfPhYMfrrrTdqpqryc4ik7azqcncG5TShbKbY7DIMatjS8i/WSQUtPDIWQspm
nt//OEUq8w3EmSxrTMcZUxV0OGLSWSvuZdwPUlQbOPAjI8S+XyY05CDi1HuCYUdE
+KityQOUk/R5dA/nxmcaDbgeRo3/bfr5L0bV+/N9/d8kIjdBfYvdlXHnLCojPnyA
WzYsRCsPJvITWP+fqabow5Ut9/C4a5t7GrR8Heab0ZJMD2i6HrWJJuLd+l9yrtd3
1UJ9IcThlIOZhbJorUG0ctNXIi4S7osHcV1m4fPOBl/sPanuHByq/cjfHvEqER5A
TxjeDpRFD4nyUh0Nik9HI+yUS9tcZ9NAKtYLfTQkiYllO4JPweLG1oD/d0lPl5Z5
75Jjw4BkdSRrFyd3o644UeF41z2bDA6SXO13bW+A+/PsP0kkZkAdXCcSQozv1w+v
t73oG4h9mpbUcN3ysFuJkAQ744p4yOPoKft1A1hZBJMq83gHi0bbPisvyo4kFpUJ
2J9BinhcTgCDYkWAOmLp0BTaLBSMfN1m/JPJe2//Ki+QB51UyRx7C33a9IwtcIlm
wNwJkEh/aO04+sxe52hyvZluQBv/lfsH1Br/E65KRTc7T5VDSe84woOS4/PqDj6j
p+j3a4BOlaqOfJXiL6Fh6otzfG9GxvxJC/eHMGxds5xY0LUKU9+py0PIKh71LqEn
x99bo6v+qHUq5yJe9qZzwsK37078jjVL74GHu2/3mcoPJ5UjwXDpecpvfZJzTFq8
zzQiGoX8GodQ517ibPBKL8bXks3diNkCQ/e6FN4nRnSYQwHLl6tOwiVE1DSXuM78
q0/gXIu8bETHOzifMJ35gKTXPfIEKhmSRm4gAmOtLSZjsLRIvN3kVhlU38GhuoSE
OANEXWjdIANtcdwC0TRtjFxSfJYmPrKi1qvMh4OGfTglFDsWfT/ntiojcWRVdbRB
qkQVwxRDJ0qE4wcZU9Pswsi7ti31scWymM1C14KzAZW4Vh9aF1x8eelSmv65Rw4W
VFay+qwIIX+HAwd0DmcEcGADy/Gmd7rwERpQl3OqavgKwmvSqABMs/ljdgpPKjol
WtyuCX1afOEzd5pm6nhvLdGQj3ctAiRYmZ9mXUPztqQ1XeKEJXpSmwA65uycjaiQ
sg0OeT3vNN+w1zVlMOsFSOloh/oFq3kvhZ6CBN66Qc7wwr1LjX4mTBl+E7VdfoN+
FAy/Wr2dzlSsV3PXHU5JSgsaBYMs04Kdyq44Z74xRwN/XSnyai0iuarAv+GLGg2a
WnqligAYuvqCGH0UYb1lHWkGG4sdbTusCdxSUU8v/WvInivE3jcOCE6EllwwM0TR
/CQ+tLAqSUeNPd9JBR2BGCWyRjEEErCle1EyDWvagNod9nsz1sKQuwZiKUw7eCvN
4t64tfmCduHHHFGgbEnsVj3ih79zP3luNFefSpNTw531e1k8B9ZtEqgkBwVaO/gb
N6WteCdLf+HIq2N/NmGLuWVK6RFVgg9Q2efX0e/xwPdaLL1ExwfV40zhIyMm5PAb
TUqKJxMHjfMwRUPNQydAtmTsPNPiL/7DVxZod0E8LJgSF8p84WGR34DxxEMcVbyV
J4H8qI07yQNnoFV+vXTroIf02zDo8wWEPaAV6el8JGNOYss1h/RxepELGe/hnGvZ
dXOIq2dHbe/biIcdMgm6L/5ywcqXpUh5v+g0O3fVHq1h7KDuqdlB/s4+5BE8h0n+
B3fkMYdzoYH2ON+CbKQaYEYwmFqnFe84Yz6oFq/siofBYwBtb4zOnQcO3fGOltdX
vO0q/yCLzJ8EHjRtcjH+pkD9q/wZe/n6UiqigYbrSV+xcvrH1IAqLVTFLKhNurnb
tnuWBnPDVhZHU4VWwaNQ+vaI83MIWgpRs8kbGL9shk4ZfTTVEg1yY17gWOx62UFI
4P/aspKYHzxGuUyofOCUI5/gCVR/OaBfSBPwrctkiFL7hlS//vDf3Bjkao6mvU+z
K8oFEgJt4PHGj1QJG6HuR2RWBWDbA0+qtRd17y64IFRwaAhKbnCC3vcIeC6yK8E1
GRCSET1pHg1B1i+tCQPWCqf9gbyDa+nElGg+G/jms33Z1udPFtd+B/1Xd14vEMSa
+lcXcKEFEyHKBXSPbtBx608vyc841G2drF5HY9fVtKyxeMRJenrFsnQOzaTPlpCd
mylFJk7wlWvVGuXB65WFUfe0Ei+uIru42i4Wfv0YQSMCT5kzenlevsxnU8jQJZlK
mtwBFlsTDwRaWG4tHM9dJnjJAOltdnw85o5iEi0I0+9NtANTBUMiyiSkQoCzHdqp
RGshSyWROvn7Km1DVkfUnVCky7r1g3QeuZWHjxiyV8SrwJxJOukP+bcY+X9ylfm4
viVsCNsUqM2mcHQzOcW5/rHyP5zMVNDrHzzHPbtf8Kh/0PGqy/FcQG5+1HipY5C6
BEgRETb5XO2sIQ/RVZ8zUVBo+jWYyA5WmW4S8oUbbhX1p+t+92jo4SE85m1Q4lSX
eSApJYN6EtXhbSL6SdVXlzcd2ShZj7smDjfjD+7u0otljJRN7A07ikhiRZlzzWBx
PGKkauED/6ejBJfQSGF/4esVhx00w8sXbTKOM+MIWQA40XIVXUO13CzLoW8i0PnZ
DgIsqbLY5M9uHxSeeIdxGn+3eQX3B0HRhxIoaG2ookkyBoRcMy/ZZTIxljb3xlPZ
yCiGcRQ4ANHEtlvKzttQ31ZRbR72SJqHGHbCPqjWv0XVNqLO2aQVVGZ4FZnqNz3M
K8ZhMfzAnkkfhxf6qUzQZnscrnvboWk5iT3olj8YV1XPDRmMWrYvWer013gYwk/a
/Sf3A0ouVmfaPo8cNcAf9dN8FP6BVeUghprEgmwZAML8Yk1KErUbSJJ7l87GFyD5
feX+6vbdI1J7PJl+k0Qwi9Z3ROlQgtQWMC3aySwbvwjIYDZODpcOsWXmh3VE1sP/
1EQPtX6Lm6ChkZancN6CzTl5jB7xTze3ZUQX+UK/qBXB+aEndUX1/LXztKmBci1D
L88GoZsN32wN3fugxN11QWyFC33AAbFUPdt+3FJMquttnr0ZqswLBpE2X5eef6CG
Xy5DT5XsPSsJ7M0Wz1X322dLKCNsbdeJjyPy/NakhZp9YibM9Ug6g0g/IGqbaXWX
1OSO+9SomUJ2sYAMW1YS55etohtAc6vrPrpZKm1FHUS8cNqewwYBeH/TvvuxMswz
DWBZZEauB2eYfI7Gnx0LVg3cbBgXIvBYfI8uYWHy5bC44nWkq9SBPKpFo/CA9Plq
fNU/mRbDi0Wn4PUELHWn5iinHxmi3DsRlrYUtYW+P38TeUIGgRkviR+N2WASeeqs
1sGw9kIXD+OysWRi5JHSVarkLDKky9ml3NzgbODfdHgCtpG1BkxKf5Vf9WhX2fok
TZjjbk2PNKQFShSGWe1jQAm/BeM/0KMv93vx5vD6ZYGHhdhV2VViHkGY6Z3Ox4iL
SN5bpEnLunjvycJ2DCVvZmXqZLpkI8K6UfqwtXyH7B53pwVU/1252DSewtbehWss
u5Wx4/f9cICiucEv0sNiAYx8nEVbhG9dZ0P3dcF/2OsAoILgxw/7orzXDfBu8VBw
ThNhmDYPWnCcaPf3R3lpWroDyH/64p49+m37sbGegFm0oPUwUafBEOGC6Pmzlkhu
KWdDSF26LXc6dfxzKL8zODw3kEOfodcLfcBF3XjBoSwJfTfpWu2M1x3t3vflZP25
zQhO4LxORYyh8qisvxaEig8BKPr8g5NKvNGcAtZQrNx6lkHtvp/0+YkYQjXlVW73
SdT4egomUMSZfurtq1rewC8SQYL7pYnhodXgVQIco9X1vkwyTygz5vaIEr5VGkDw
Mb2kKxi/jQxSsIkN4ReSBJ4tqg9kv7Qm13tkeptA8MPJuo6221Hm4VNP+bzEPpO4
j6Ox5OTG+sFsrXpueOCQXNFH0Ll+oqs890Z4QWTEZr6Rl5pb39U4jXbd0Gj+W7fx
9S/Mt+srjTYoycQcjLWscQtoDxKjleumbSDSQbWNtvNZlumUAa9ZdxA3OTFsu1Fv
eJyYOEK/akgbHuf0pVfeW5O7DE3uO/izWueFLNLZHTytbNDkrl2KCVQ+Jwq50mn1
MVI1wDlArB886wjyUIRn6/rttSnWVvJInTGYrC0ccnO38i22YBM1w/1BdF70hsaS
U1n+J7n14WSKcENVWodgadX41U545EkW4w2FMLgd24RHD94lNmpFmXjtaePHYthk
/q/J4gw2DR3KCCyykFPXYKBDMGJvsPfX8HZv5husvWhzftrRTTWUONYTirzWZHex
Xe7HAPzWGNu8XAebs6C2DyHr28AMm8Dz8wXxUu2EJCH2+vKJlpdLwv7GBaeRBi11
xls5S6jBVegoZ7ZPIDsofcRbZI8NkHFQvzXy9zl6wQTSf4Ct2+3Y9km3wl/B/m8L
OhNTSwBLe04+A9GsAVMZyowRL3tLkU//Ec8SQhRF6nt6MjccfHqug6n7IRm43INT
ng3XWK/ptPUlF0/ydaEwhrSQ34BJB9Kukq5nAZuE0WUzqhLm4ojsR+4cBlghZRSd
/GCuSdX0eA63e1mpssCPJsbHuM8NMMYeYRSBaw6QXsqxngLo2lbtGW6hVwmwI9+p
CDnVn3OZPdeuaB6Yh24eb3DHC/wKaWNCJolY4SwnpMYJi7KP4ZT69u5244hhTEc8
D4gEbtbWIN/0tSMAy6TKcVXmcx8/dHx0pUTlr1bcyVABSSiLlRriEnFRtDJA0KNe
U4vMC9oPb+cFS+qA3sEWm6YEv+kzHDf392Xm63OTzxtHntAFhorwLEQCPM4WCxce
A7cI2bTxYanMQ0F5/IdXvWZ4vHMoVero7L0X0nUBM1miKwf578oUnCv9Ei/n3sdp
cKhdJz9WTdv/VfeLxMugS2TnqurCpDs5BVbxf9BRSxHCJ6P/NLbZHzcQQvRrq4aI
00pKkKjwfyuzVZu35cDVq1D7EypiEikIqqFFnLkR9Vw4WHiPQJeL8eOx9Zlu9H95
/VkbryfYPqMnz6nlQRKGMOUrb3lkpdSpPAcl0LalCxYaG8ycG9ZxqwdX+g4wkl5D
6jQlRa/T8jp+5bXL2SwAlDUngaGjkXiYEjK4U3jhs9PyGUTM0Ng9zTMjaEI9xnAc
KkmSJKoip86KV9xiH8MNOSoNRmgK7IfMkDtrnQmtY6trHfCoSfd/cacaa8caRNjn
RNAO9NiG4K/iTg+6RQ7crIVQw71FRrKrAE4YB/cMFHfHqFvPqaf9DCTh20LiEWTm
/+sx3Ya2dMzdDTRRqAQuWzejhinNCPp8oWY501t6YCdjwvcc/6yCTpJyIxYtRfWo
bVFWvmm+V24/HcFbh7ZiDPG1y6CrKCaxLyMaHUWk/eOSXcCfglKnFHX2EkJaEBa3
CdjPfnCxJPf4qsShqs45cgGY817hpwaKMkfgeG9ozurTXHenlja5LeURvchGTD12
scfEL/NoqiQ9j0Unnx+T5DTTB50LXw0XHLPwQBoA+lqA/f7ULW6EET4kYXjQHl8M
HUhvdma7sppqO983ejuO9f/OaN3HU3AfHKSXizWCkvoB4ieJO1uh+g1++pwPaltm
bkLF0nX7vXCsIhK8c5TDAbYdmoM/9vypeR/ZfwjfYeInhiNPY9ygEb8QhrO++Plk
m5kz6lvG5T/keD5sSfBR1o+3Lrfz4tAWMjGcOTAtB/Z3htF2k0R7OWI+qVlIZLXT
v7qUFAy9rWscvNXPkvIp4YEwKX6PHwB4jzFbvXrP9bILMl1jCfh6ex6hYQl+bdrW
z9A2i5hzF9K53Ack2ydT0ULcnVZcEynrXoLpisW6xBgwXDKuYGJuhbERxKVlOQa7
mjaYskp7CV1NDVz8eEG1E8lNWydtTUJjPZsWEPmXZelKBLLPxi4TpWR/CgL3Lw0W
tO358nGYjtL1P1LIVXDk3YSPpQUy+Alz8J0P6vYZfYTF37PW2PgZq7EhoLNj2wCi
4WVgGdXpOmbMnx2C1Nz07Zh6FrNf480NKS+tq/GN/W86hrKQHmFR58qriAxQe5Da
bnCRv1OLn+e0JckLt7AMnkCV1Le0s3S7nW5FptEfJG2p5fAyCakCiDyHijAQ+M1c
GMi2kXeuh9wvYM6UXUWym+Z1V+rFNEOHbkJMKRrC5H5tiExjedhEq3RrpynQ4ose
ISkLnf3vajcJxoPkAKUEoiL2iAmHmAw+wVJ944XgubY4He7ePypgj4OgFLEYxCDP
nqZIFa51sUk8Ke6tq2rU+4WJt2JT8GR5fI6eHx2POSyCAMoJiTMckWnXjXsX+rsZ
tQ2y4LAF2HqGeFWluO9btBP5X4lfu3INt8DEkajckFmkjjH2mHdV8X4NzUmwbKyB
nDspwaeST319BcaqWulcemqt2Sc7y7fFcuCP4t4SIW0xX8gb4DSbv0dJHGCIWNsh
VDA6H/tzOPX1SEJQf23h8oYDKmwrirrOtgmzCNUhsQyaXIuLXQk3hoQWXSEsXa3o
CCYgJE31kHaLzBYXI4cofApBPiWwHVN+wE/SlgCrrcUykiy9w6zMMBR8SKWr9YhV
KzZzanSHIab/JvjcpXefeHe68to0fO1k9C1QaWziY7GOwGm4VnBVBxi7dVA5CalB
Uq2cR7wB6g8eZ4ghvixupd71+YpdJ3O900ZJMxM3LbhfYirS8NRomnxNg9S96bF0
xHxArZxk7ZTYR5doMtY+5VFjgoBFobLnSabjyYQ34l37Ve9wWxxdraDwCNlx/EGO
owVilEA26QC28ZGSVDi2dSAoHDqL99me3q1E9o22AzhTEO/Lhc5mOpv8ANlXXW5c
yqnSf66AebG501ov4v0t/X91PAxMpO4BzMvsqJ995qkmGCi5lWW6TgSc9De/pmoL
hSUKo3e4KG1ikFItFLOIvCR9hKso6ylmZYj3IrvpjTicqJqu/KRD6Yvxbzubab4V
8WCudDxtVNQb7uob+w/MFNVSJHw2UUEKmR/ZtBRiS3VHIq2Ehxvvp5+iJYzlkUV+
90i4kytZ7SU1zmlKPICohRXgtBolNR7K+M3UFNP/CStmOfYIRSzTgoBEFEn7aEKP
rw2hbOuxpHb9qQ0WHH8gyUquRKtrtrGJHpw4BMLD1SztipUAVq7MwStQtBli73hn
AdGnDxz+mm9meuO6yEEYs1XHEKZTowGSXQkqKjV7qmCmFpYRoEh4cwSWTbcwq9ns
ZfXasPydaGwkVkdXPIEgLzeZZUjHYPVMbTjF5wLFz9JMHKXJAtsO2bzB8UsHOBBm
krkS1UAw6NqIY0KGxOl+fvu2vx7GgSd/Ou2jCqfW7aVxYvpub0n6G6/4iE72K+6e
yXqOZ+tBxgP/vLyB58lOBkq0PmA09WAhBfTxyeo7ReVnjDYCqKU/rPEXcbY46BkF
+XJSf7UlHn5Rj9NObUvonn/Tw41GCXaeFk57Y6vm1qebdDLv4w5bHEWFM7GeXruk
afaQh6dUF4L0h17cKv1wUwpD35dljiUQ8AdSof8O3RPchbFbl7S4Ig3eYyrMrQY9
xbCoLvuNc6uYo5toL3a3nWwdot7Rd5oaxGt0IHINXhE7fq5UVsAmSz8JGu2FivfV
5dSS0WN97Cbr0gIWpRO1KnKPT++DOjyWU+qQTqVSlAr8PHEQyrLuD+MqKo15NI7Y
tmWcYXHDCr3YiTXd59ybKhUsIDzg6U21UB+zP3QFxNWC+Wg3SaUFppPGuL2+LXTM
kZpYMajfTeGZkcMMXj/1rcN/q9obtcuPr3DE/IIG7Qt9eSmUMXMm4Q9FJ+q0GQ2O
lV5rtPrQ5DTLTb5QVRw8xdDRiQT81Kecrhu9hwVRvuUyunajc0wuHJNzeLRtqJfS
lpyy6X5Gm+edT1t8B/ZP36gwhNxAvJ7AItNApT8xYKoMrWSNT6vFnVDp8faSV9dk
+4N/mdojipzkNs4ox/kE9Q3J3HJ5PDnNMT56g6ys/jOafYK/lKmmsbIiZD+lNxkl
TUPBzmwR4ERDhx3mKzRQdjrxxYYka5QPkbQpxI5HCcJX+zLhvh6pqRSQIghguj4D
+q1CwnVlQyh08vk9DRYQQHbxR1spYbEk8/BbBJ/99hO2uNZBxJgO6TCLmeBcSP2V
RjEdArRuzMkKpTPBNm0EZNnnsK0mjie/m2NHCkRcjbnNTK2lsXHbc8T0Lqexw6Qt
Yqj2oop3XOy4QiC6jGODfxKpyHIs9TjYXJFVWTTxkXZ6y8nNccUpitZD3u1i+omy
ascilOcbqUnXjeWR/9oSedu8xvQWzTSioaBd2iDus4mWHm9wc1XlwCnLDu94hoKs
JA8QWnxvuNAlYAINYmD8W9D+5FtZseHnGSp09TQsyvuocx2h+xT09GqjOBx95DAE
zTtJjHD8jsk114yAd3aKH0XIm5vGcpYKy2yqybuQufAMIHxI2iag9/Jha7WGbIIP
1xsqxQLFIIb/g7+quXQ7DrEtBn1L/54+FLxulQU6V8+oXGFdK8EDlnUU3s8L0oi8
S6vv/HFLtoLeCa1pCG0hU8zObEjpg8kOnliB+xrgPgCA1hYVEPPzNH4ci9Vta/Zw
cfsIig/9Osqt7E7B3gCy6H4Qcs97TCbA/gHCNo1jfvn5IU8QHMRxd6nbRDdg3tAT
LcKdpUPVbjP4P6HE8hzWduNC5+Rk+VtprY2FWaym3K+sIBHDpS4uXLLwf779o0CA
JnKxcG4+VViLSQO37AJRqC7h0tAbnuw5HmoVCmO6tPZ4e4YvWoabCx/qv9ep8ydr
3VinPjNTX0HaS7ZSLcZHa6suJO7j/EQATm6puS8CsVR6aXdHeuwV5haYXBNpNDHC
2/liPs78cVYCXvq8nLYmL7WE68ju8W2kyueoBgJPTfgSFtPOHT+qRbx1T0KBbCNh
Sn87bxVhlNyVSbkweWazJZ2TVbXljbo/XKDq2qhjfwRT3cPcu4eO4RxN9EZdPRRg
EXav59zVja2snfP2jk71pO3opVYbUNLwNXcVSSWySHCnY4bpKkHcn9a4SeFZyGxd
23OGKXGgkg25pZ+elEb6ptM/Az98SlH0/ITzq2TRNbAsmtsIz4Rb6oeNjmo53+o6
UXqAWynJnKkEWavgMPbi6Zrlphu8ujB3aYN/HmVALivQRoYGwyCG5j6a+/Kmprw0
f5YwsGc8DwPAbAlxNPPj7NdbC3c7CmThJT9hJLpoC/HweSTOJrXO+4EUDtPLgm7q
9ZBnTgK3OQk+kDv+JeqaTh1+Z5+Vvs6vpVUXj0pN8KtUBZ1/XC5umuYiJgg1p5Re
BpoOk1oqAdbmafRyfxJtIqEYFRPF7KMozB8jOy0SnvuKiSAbi7AG6BUEpaakaRXB
8NG2hAZQIb3r5+4ane7fwz/Kp9G9AJszY1USSsTO//ZohC5xgupgEKFad8wZXEl3
LFWoxLABibCYtsWsAGRmPN7iaP7FVRFL9vCfc7lxMAeWQOPbb/To3XMNj87ODmfa
7C+1/aMmXsGT2wDM7Zu/KT6cISr73UwMFqySuuQl6xMZRNNa9Bs8uV8p5OCqRu8S
Y+PO47hnOqlilyLXAVEeFk1v4wdSaDBGo+xcjrTBwC/fjK5REJu5ChabiaD2tgfj
H08gcT7nZQjSMNygUMuRujIpevwMod/HPxPOKX3t3O/FCgE+Twuhg6iArG+/pkSE
TJwoESq4/dKfXgPvEzQO6iaUbKvtxyu/faLP6yofVro667DF0HsuO9u1jxUQdSmV
5uQmlFRoNKAqATv21KgxyrMI+ks76A6Du6AlAordRN2PaV80U743yUUvj/ImEyMJ
+cfJjEyMlHm1JXveblSpgi2nWAVHNbQmmkekyAuHKmx5LHbO09S6AgsaNyN39i37
1sV7906CG3CAuKNF/FpaZLGFUQh/xPN7bLWyxahu2d2rE050qQNrrhl/Y5GNh+PS
IwoS67OdqQT+1iR+2pU2xYeeC+QOcFIDr1CdxmBrS374Pngne/2YYtZxECJdSGS0
3Gdh/ID6XPEH26XZUhCZm2gR3Y7pvkN1wd39WaoS1xRhwdCBD9lR76niuJqEuiZp
IXUwHePNlIjCUY6EdhJkp9x15h21HmbnmeXgI2CCm3/2I58mQgujo6f4peCEMbG7
akk2PASGSV2gqXkQmIpFomjnLlpMtBhEMVSXQMdirfXxmC+Wqxs5ZzlbNGPlDQvl
FIGBz5VKpS8zYn+9ymjAPWcvC0NLLzqXsgzL8Hyn9m/6pCRlfwtWETIgggt9JhY8
ATp4i4ulC0VwOp2jrNj5zLn+LTY1lkTeFEpfltAI/nJAySjZX8yDx4RZKsABKAG8
Ry5w7GUJH8JxLfUNAs7kWHDvjFu7DuHMMlDlxgbB5HZtRnr/2Eyg5XOmInjwY/BG
1y2MY4h3nzW02+Z0SON6toUExqUhFCU5CPzBEtp25uIembcaBNb+elZBstWj2rdV
j3HPOq2VkA/SvRGYww/q+bemz4JY6N25PmmiM5e/j1Ek74ZxUzU2YS0bdYPvSPA7
lvbtt5fMkirFWPcjCXN8tZxHvw3hMV9xKzl0BZ+C02bqoRs6/GwwZ4FECFCj7LWp
SRSjDQ6wcjdPBj3SAzby2P1ryrxwyXJPLIGQyfzHQclXQx6feKQtSd7nKDz5FyHB
LcDKM4lxH2vegt6ZUobBRhIFwmyzkvuWHjjeSvsKqeSk8PMpObsKtVchFp5Ym+pW
sKz+jBgw1DjGJAa4qDxHHgvT1Pl/9U1jmM5htByhSbh/xGzSUfFpFsnEQEPNjtMt
WEMUdCBAvns6H1cubfiKUW30T6AcWx/1G4v/ez1ow628JgZUxGDv1579HWS1gAyh
kxSNzYrh2JOWrQ4OH4f1JywWxX9I/bq/PZQ4x9wMNCqWmOkwdOlgVMeCqvPX8OfM
a8HDSMjN/5DP0AJVxm6wRcNiND5+I8JXUTexf+s8Ao85850sZDF3pw5lLlBDhwFm
LBeI6fkS1ugnlZVEuUZ8nRPyewPzlRXOGql0z1mcP+9PaqkFR7cfj+TBP69h3KRm
LiXtXvg4D8696sXvZMidFWvSu+6h8FdwxNgAKlkVaDZV9jutt9T6vZCxDEGwU+0t
yeFj4SOC02GAQKPlywK1GwNi3lpLu2e+NpA4UNKv+HF5S29Ml7MFA3yNAPCCWh5A
rYn8JkLSyxgG8ZFO5BtHxIXc2PZ5vbJXCo+ZFEGtiOKCt7zrI8yP3QtvLI6ZW1Z8
ewEwEDzvc9GbE28bIQPycU/kvLxL/A/mD452itTRPn6XL+xi62Hprk2+81H8Q3QV
dezHC8t64QctzVhUseofUSP4xQ7Ei1hoKATI3MFy11aXYJbzzKlzhsmDyAiUvja4
hl2iVCT7QxTlnlpdW8EUgb/vy7FqbvhIk8wpWH3bYijIbX4O6wM1Vg7kT6VKGio6
nEolIjHEN0A71s7ba3dScn1qYCV+TxaV4gF1MW0H0UXEGNAwl3CiHflNbxvTjvOQ
S6if9zC6W71uvI7iNyDIB4J0kKcRhrEayGkEidkECtfjtAjAmJ7nt0vcTxXVnzF+
USuTMUFlUF5gC7PpL3yBRbvjwIkmQHP47By/QppJKOsnYDuajlHUwwoVZy5m1Hgk
Zjphecxvmqa+3R4BHXh2yb7x6RLjab851sinsZNdrKI5f7IQH64ikjIxiMFBZQ74
EyqWpEBhbUoGmN2lMemJh14Pyz7nQMHKH0k3OXKETB8PofQKwWFebw0WewajQkRD
XDHmJKj9/sZa/ptYkanKQQapdKJzDq7N1VtKSdR6Hg2GLxmsP8F9CRLK9HdhKgDs
koJRqZkZzr8MSlayM5twdGd7mdMdEXhKotgMbffCpi9qnFadJdA3+MRddJ8gyFYa
HpnjT2INo/Mhh14XDF1XYAQJaM3bzl7SnoJNQfuASlcOYv12X29VuBopegBYwvuf
OikqwstjF4ydreXB4qn/iq4v8ehAi4iNunu9iD9dE5wyp2mIYW8eXzPsaCIVmgFf
US9qd3PcnMn1PU/bZmoHdngGh1U2T27l4LGvRRrejBDZtOgtL2L4EF0+J+mG5QCm
13Y94Vv8O0ZottzQuKH0uYqtaj5CDXxlejTM0Sjo4HXICZyGnJ+4MMYdjMbEoMwb
++6dGr3U2L4d64RR7Q5huF6s3sikXm7CS37VLUNvvv7NFnwAOGBOxARJbEQctRS5
Cck0wgRxoVUF/dHNZkAEwm3MnAhEZlxctK0MN8AQA3gEwqIhjmEfntW3GAQIACCj
Ek9J66TvtI67X4QR2b6LEYPP7c5WmJ0HpHtBZjo5qMRB4hdE4KX9f4ep0FKEPZOZ
26VWgyABm1iCY8Udj+PZ25G4aCs7llehTCPGH2mN2Hgys1iBPDeGVoLjPGewVHaU
GZoISF0w0ATbBzabzHUmOUuGsXMJp0uaoT+R30flEXlL6pSmCZhNymenb7rqxAqu
NHNH6nGXQYjOlkhaQypMElyMsGJAv6hT3qYAmJfAdRloDg0Vq9d5gNCjUqKSU89L
TTt3s5jRVk4DwJI9EtcNjkZXRNqow1cmsAB3QqkfYa6X4WvWgP9UeGbFf91vEC3t
YZ4LDNypfzo9lle6ABGVLUcIHRXdhMinXc5lyFTG+AId/ii1XB1N1IDZDfdXd0Ya
BrIgMgBSA1el2umhXkqVsEMqUrTdSD2YVtzmfq6uJJspgSTP9Xd9yqJjIFB+ZSGG
D0tcM6NTVcQ+cptlr0mpvS5FKPcHXtdQvRbV59itRgehTcojWmw7Skjlxwud0ob7
bQJKcCQw1Hu2812EoaBiK+jlQBTi/+TLqQZu29sySEM/rULh8Pb37meLEc2Ru3MS
Sxf2hjjxDgEgPgPVsZ4EaoiveqEnDUFUdLZwfOEn+47Ss1SHGqEgWudRnC9hMld9
eKdMSVm11y3o6CiUo2QbX0LgabydKB70lNZtd2Tz43VVH1GmyFcVAZDG6t6Ptkfb
qDVSCxzMLL2yn3SRk2qT+iVXtNL3tFyHi61HuPugilfWpiPks2EPRbbdTAFqkD0t
FoRZVtBLKF5QeYmmf2yOqkQ5klMRh31laCIMGjYRcrkTDVncwfFTdHe4zJqR9azP
9vv5eRjnhEkRwwQzuGEJC6Cmq5JohRpezn50cLb+sKnhj7suu3c4UYJU2YgmSUr7
UxFNRtH+QFKf9U4z6dc9liuEkFtXmE7rJC9DNGANfDegMz5GoZcgXHWnW5cd+5SC
lyFCv8dX4fp6ZnnW/9/OIdkEqItsQVyrMfpVTmpDG1Vr9XA/jkFyks12EcYwgcTv
TntSDo3ZCu8HJ3ZXfYJCXVFhymvGF2kdUYyJc/WofiPWvIeyKJcCQp+gYVnET+Ij
4nbhuRp4rwmdjONEd4YE8byQIQO8/ZuRDM461Qo92smwOyKeN8XTVNs/JC67d8JR
y63vuFSP4a+yI/0r8cHubO/gKy9XxxwPr3FPrbtKgdgTwd1jsIhx1DJ0k6zztF4u
vL84oPgWyREx5TsdLH7iHr5qsPysIFCuNeJMGsC9GAV0xNNd2RxI89JKLt75WNr+
06q4ylwBdG2f8bc8yU7NXpknlPiJGpxBCa/w1bd+JevNYO9GFgxXY0oPLUVZnpp2
xDF6jdSL7/jHmU/5M8qtvS6zPMstne9HQ4WqEcfpEbRbnE3VFip2LqioyGcMcmJk
B9IVvGfzMxwYMcb/dRA4+dalSuFEAU1BFte8Habz2wE0Ec9/ZBIRvzQKrLyLG5HZ
SWO2lu6jMMKBkZrMQpx/0xlS0cjsdYRp5efkA6s3MF4eiezMzbyVBTk+AiASpFys
Dw+Z+dCTCtXj11MO9uadItkKpyNuI6+3i5wEBe3OcBSD3LNjgNVO+4jok855xX0g
Z98HVgxjDc/p6hHCooipkwZEF3F3hhLyVsQfumeiySGA/2HKXhgonIo762xX7CVK
3GU3EZ0Ym4Bcl++NcWzD3oD4E39LaLCYaTGWfj4n0ukrHWoVBUO7MyQVBqF99G/n
1BTblC3WoGwgOCVbJSzjDh+vCp5tmA3NBuePgyt7cwC/895a6YfKr5XrO0QJq5xA
rzA/fs1iB3pEsWKEAhVZfBOCUL9h40Jbu8UYBgdPbFeAqezSwF9OWSzl8D5piR2w
0IcF5bockjOkz0MvSGtxnm3s4/Mc2/gFQoixlL87Z+zIASFVYUPN4+zMMKPmlWWy
P/HzH/J3wr0atShLLf60gv0W++8N2eSI+TX6DowAPCXqVkt9ekpC8Iog3YWfgBzu
A+bqlhiJC/mepOuXGNC/xMYbDb5ftp6Efq3FjQlsFTiPKQX8XksK5fTnBktMqY89
cNc8gw5JlBxDI6YfK+rWPpUJWB+6rAjpqyn/brecGmr5DY9GwoEJQPM0u/Nvl6jt
5uqM106lkHhwcnWJp+rBnigXhf5/dtIHnmPcS1hqbVKSorKWKYWyJTTTDVqGeBlQ
5PMbi2EUfWQP9uvQ3MjuFyTIM2sgJH/ZwsusCc3l+ZK6sAsea9qc+P2z6PedtGh+
p0MHB+FvR90h6OoYZ2M61t6JKH0jQrX0DDirkXvIHYr0TCusDr8mdHx/tcuENoVx
eQtALlrRVLNfhGHHy0Q+/aBxjiI7Y7cAxFm9O/TwTs6Qr/uPKHNRszyjf3XJRZ5G
PhEfao8QIza21ARoaF5D2/g9sB3+ZaZa1zsY+tK8/MEUvtBBkbrB+rfvxEbcufXB
kSYFDKXwC1jifsH5plAjwSZHhihX93pMd77hyMIKI8Gh/lxsyZOe8Grr+P6EdBjq
V9VuCBIWIEggicVELUfto1Z8IRLzrWINk2B9p+86jyMU6HmeVT6dXx4E9L0ns3k7
aCG/N50H9qrsYLiXYsp+bNIRPTXsYFIJMjwZ+yMzp6Q2WyMpqWC5TNCSr5S/Fe0B
uNQm0k79aoqkSDFKeT8rgZOpfqebvWVuvd98OZofRz6FYUod+n2MHwy8OyHjyjvN
WPwy0z8xbdJn0Q1sPua0+9/UNtu8ECwJPfJ6woGZZpfzcLMBa5M0oLwQBI0MWquW
wN5aXNRmMl3QTeCVzCh0a/lunfMe4z0+oGk8rHd9T8OBoMf3oaTorQq61uW/pl2h
AA0u5UFCOcKbAmVvRvNlPYzdYX7ZWtPs2xUs+DOFnHrS1vpIjVOcijNKsz2z24Ec
kmRyhTCL44X6mpBdT286i06YIBaCnheHxRWhLvl2qZCoC0VKgJpxn/SdzfB0aZOW
p7gnZ1hvz7AgxU/UlMnobX4YxASMBMcG4EQwUZh5GBBfr+505ldFF3pWHG9DO/6+
veOws3OQX22mhPKVX0fqyRR7AZrwpYi3zROF25dn6JicBSvlDPPMlgowpy/8vI7M
LRQRKO/jrx6k4aGYJdquGNiiVOq54JH4h1AauSgPxuX7biZSnrvBAhthXcPrYsiq
ETBf9bfv288O8RYEvXsZ21h3HLwNLig1E7JTeWyaBnXqaiPMaBGs8PuWV96TltDf
WWZ11UV2NVYiHn/etfnO+gJKXZruLr4OKdzI/Bm320AsplZuRAV5nuo+4+q/7H46
Lfh8s8d4sON2OaRdbk9oNYbGEtjMur6CNgQfcGKAHQXfxW/2lWCREJQxh/fMYFiY
Q1ogXMtglCYmU+3ddz5CTR+CHi0YhoZu5bnKkERlUmAZcjy4FLwQvGXcFy0A6VVb
tvabSp8RPWZux18onCk4MM6HSdiP5oDt8eu8bnXvERKubEQ7vdAzqOc/7t3ILkJI
YV5eq1UHhHQAM7ecJfOjWGeLZxbb1Pu1mWJ8pj8foa81oPhDBkwIlKuLGN2DFajS
Y6O8n8qy91o93mg4R6RHd2rtLneIzEkr+bZ3SSrFqxBZNOVxV+Zaul7/fjR14kHg
0iGPpHmoxo8D+A7v0aGCMU+dy1TEUlMBGVbh4SwrdO1hMhzGFkPkE7hRngbLe96J
46iluy55fqAwceqMn3BZB2cV+UmLSE5S1NJDD/XxmIgDC0VgWB2UI3muHcrq5XHQ
w1EI3kzJAC0zztXyGKCNxYxEzvL5F6EsqZ4GNGu4qlxmw3FmZUmSN7LnUBgqulRT
gRpkLrChjO4Eb2AI8HUZcuHASctUxWknz0YXiIhAzfmDAJakxtoGiElKZSIAhoml
kUNpmCrMm6bYlvMOSRb+IABrzd7K/JsWK2tPGHS3QsjNjTJB9ENkqvOq5RSpZ9kR
eMcgZW5NQj2820UjK8/Hdwfzkj2ueBDqX/DcWfFlciPZ+/2486q5YbBtSoB/492V
I0omNdFTqntHqLTSJul/xriouaMOEe0xpxko8LtaVOMD8Nqyu9B6YEVAdTOqs20u
K+rfiLTuXcUquO25/zLHIjp4AHtP8TtkN8xzaqRfi//7JEhXdN4X79Rdv1DnqK0Q
Lk5OWmYC0BdEUEL1kHhQNlJCxNDVY7lgKC2wzqTIIjOIBCalDccYrL+EhA72rwTD
9sHGrq0sULAF9Hf7xkg/WyMgk4gAdgd+O9ULPyvk+j+ArsNtfAk1b3DHKHSuG0UX
W7d+BTurGvSyX0d39IWLq08uwD9JYciZSIWvlpQ0X2zv7CnmyfxdY26W3xjGjGjS
iAevcexNgqYx1TGlLrzLPIBtulAbMSP/upV3ZkhljcE9/FY4yeta2K+7RUKilZjr
sWnu0FTtYTW4NPyQce8fxvzVM+Iz8pe8WVtRlVUC2ai6fuFEqOnJBB93FvKmktHG
k4qlH2ZUEHLLHV20q10iRzFPRXmsAxW+nmxmRpz7dvE/qcwrmFfhtcd9bQcLH6Ll
jGAjeZBD9AJmqh662o3rcvC1EZdPA9R4djpN8HjnXblxVl6bdAxXs9BRYdCS4m90
IUh2D/QyIktefK9vZo+XxSv25cV3cez4Af9cnY2e+ZHSMN1wpZZ3cuTFzKOC+6ZF
omAEE+Ef6eTnogF2Uv3jKMnsM0I6eE9HdMgJ/1nscQM1CbqZc6LlBtNRMRD5VWCw
X1cVzMxRuA8kk9vs+nQCHkyH4zCVuvvAmmV9VJNO/HKgRr+leXbGAjD0PGUSkVV8
70GTAVNVGHvI+hDUWf4XEJSX0SnaOiPQMTjfzgifMp4TdiDIT8Qt46TEGEjRq+3A
pWY6RYMsWm3y1rjLQPLbgy4AK6kYFLsO2VRRoJDGKj6ufkmcwSFhF2p5x1rRTVLB
333rneIkGZq5wHQllo2SWy7o8HSjOUxUW7IHeQBPOMto7PzNU8in2w60+hBdCYSM
uvbanEIfxdJsSkUIT6PQkctsPX/Ifm+K6RQksMmQD4l+C41QPYu0iBY7XDjtQdkq
UdzKKpKyf6/GmZr4f2oYufAHVeezAI3fJzxDAN6sqRkFZDcCgXeK8kgpXoSL2PMz
Hu23Mkg6rYiC5gxZLGQq/4gPkv8/l0Xy2Wxn5MbjPlH5MJWecTTwMdOtGKihfXW+
OJDSHt1KWjJtMRc25ZgfXsM9aPxMzHtqiC5Ede4TF2lKpmvxqzwtgvjjsJCwya6L
iakvTKHPUUH43m18E+uqTyuWyWLbCb+ggrJvBVrCRe098Rv6mxt2nkK2Xaj+pJYK
d0Gmqy3W+syI6Pjf/au3GXn8QrCawp4SBs6LoCadmuDqh58R5oSnkaIl9QCVmUFD
kScwncFC9S/YkrVogF7pGpS809zoWd97yJGuTxBFGhgTD0AQtt2jUM/qrk3KRfes
vtCy1w8xAeYtj80ITfThquSjmpu//Vg1I2xvDK3Ot/MvFGt0dU5HS22LKbsfkbQx
ag06R4r1A0qbA/311jba7AOh4blge6LKxQ1SSixkZKtX3U+pdTgu5yBE99MpX44v
V7Od1xuFDFcCbN1fFCVxVQimykkztA1v0qAipP5uMjFR0DKiO2aYxMeHdBTe/hfB
WC9Pazm3CwsdsBPNIgblXP0IiQg7TJxg3fBvAGapKzgVl4llPSwMMmPCmWW7Yi99
208g8iKkEbO7RYio8X6RmHitnKqkVp+jVZu9Q7gmNc3LwZwloXIR9HEk46yCy6OH
+G/RhDLAkPXWoTC8hDbFgcZpRF+EIe+pstjsyMCb7TBBe4nyB/lWD1L22jPu0itU
/3z1nAvO6cBHlrzJ6dHRXRKFI4Zn7SGn6+uUQjdi6+Vs0S4wTq/wANXduUZjM1Hj
7+WQjm2hmpPKdpXLBK8YfZNPgnM9dAKqhNa+wVtc0BfPqCRJMOciY4BZxaT209AE
ocABW7RQU8Z2g16XDLwqxcqWBASHpn9FLUNcuIoPapPdAFV7PRyUaU511bSS9RuX
afBIvzexlrZaYG4JCCfWrb2LuQBLmOyY/fOOfA0on60f/MoDToLizExDNI3GS68L
O1MJhZZBevgh316jtqyTQt5c+J0apCsLLez8FC4GawvIxnrT9W/6hnbnn0IE92Db
C7AjAFbvaeUeyb1j53Zf03BlztLHUg6Pcc2MwDE03jxCGI8deCQ6nMUBuLgFxzwx
JNYaCek8k64Kbg52KT7ApC2SohqRcwMompQ7cHNLK5JZVt1inloMjWSOPvEc6i6C
lawQ8RpapTlrF/DCjxTzDk0cTSGjmTbepVbFaRLohaP61WuXC6GIbvF2BXTe0XvI
fb3GJi5LisiXf/nTmw9aMVWjOty8OiGFmk9BvevLItoZIME2R1Zs7h8Fb2y9x0kS
kuk0cul/zseyI+OQpDziVdrDq2RbNSs2nJPn2YQHxU04N2vLR+KmjVR+hAE0OY8q
EgP7m7IHPnoAXpxNTN4x8l0rVGSyqb0q0vnm6F211NgcobXLCA4gHmL85FmbHz80
DOVx3myPkvHPTaMBUZHloZX6qx3XNPhbwpFv0eeaZQxRA/CkU2et/hJog4jSDo0N
PpOD6aUVy5zLyVvSWulEvhaJvOxspSpHay9r/h1/XlktriwwNZQ8SfQ//8HZmnJs
y0KOM8tKQx//HvGdedhzBy9zIWr1noLClfFPyFq4dqMOgjQINsCTJx6zpT0t+YKl
EVSgAClUQxI8Aw17m0N0jCXLfMbQTWjtDLwiplxB9XmVB845vTWwQVeWbyOnb/48
thEaHaRAX7o+7h/EfsHg8AQW1edJtKcAi6gW+gZ1Nvhqv9WBRVIR1SfodksRmmf7
v7uZSIBqzCgRBhoIDAUTqaAY0uRBo5BjMPX8wexbwWQpRMcieIWkPk8qTWjgDQ6F
mNPcgTB0TUc40DFvNqM2ibTGRt3lTYW+1tqJapa1UF4X/imm6yadA07u2bLGVyVi
SPOZ78bf8SYsF86yXA1Oz+yF4YcdTdYoeeLw4s8qiKWQy71iFF2B7XqgskznoNCV
N5YOLu2semCWlcOTEhAS4Ax4OjmvK/bS2b1W39akTXZzMov7l244nMcFatSXjDzY
b3IGuzu1viIkO1veOFPIH8mw1WTU49F0+ViMqn03hi/qUnmcluwerZ08AYyzaUwg
zC9PGN+cW668mPD39NBfoiT9mOUnC+VGV8MViwLv2lLOvk0DLHa/R1TSh8gAUWRu
A811kzUjn2GhgJcy+j2KX2itn4aUQdZP1dD1JI3WAou9bd6Q5BrblYHYYiJPo0tb
NjZKePT5/7LWihEXjNWnfy008ZDVwqa2cz34DtfmXgrsL0MGzgyij061J8UIE6IA
mONuvq/JHu+abns8AtEUAeM6Jd7xIMmTbVpqMHjW+TKUwlOEaqVh51cslU1+ZAn3
a15Sr38P2OHatiIm4hG8+7wOI3xSGjUMaFO7ABF0mvlWcbkzbQhIZAGuspIlaEXw
3y4zrxZB14DmI/VWzXOcP27buW6/WzryGZ34X/65IxI3zM0b86f5gi+Nyx4kFAZp
vimUOvBpDdK8AEp2M6OeWRyj3KTaij+NA04hxnSzzzaECBPXZS3e0brbeRtgci3T
v4tugFsYI0JlT05YQJ5qY3w8qQhDnKh6SFJHwsi04SQwPkUClav2wN/M8ziLAm1q
Yr+NhwHhfFM6vSKX1jTp3OTba1devjFjrlKQJVHMryB9NopVsep3PuogKSiw8Hc3
2sGBW4c6FTr63ir9XLwkIv6KH6NmtwhnZexsD2BKYXB/Nn4sWO9YRit+tY7GKHFy
ltfB4b26ea1+D7+7fzESl3jOdWABRBAWcq3wdw7kJQxsxf0jW3DD6RzCIEXJRqYE
PRzgymvixelaDHgoQsdF6Vp98L1B5TMw/K6FxNsdfmQHolrPl4qsRwBEYQD8Jp+B
05cBijzJ3EbCAplEM/PJBR7PqiaHoGNepKxIvd7TXotT6uFqiBih2whPLczEFb19
Q/5r1d7cIycbdhtWFexceFiqRjnVbGeqcxSqrgBLHTKngmYSN5FUQlntrxDB7yoL
OP7H7qPTWfKamcT5Cw59UrzFXkVmYqDCyWrgq/9pBkpktkpiCmFuY9TC3q3aYhUa
2dEqyQy8rjQ570oWU/7b5HPVQl+z995AO8TD/YyQgB4a1P73aLTpTb+jkU53RbgO
QWEbse5W1pSHwHOzb/yUuL5wmdZt8CMwsTfyVSElB00pi5ZUhIXbBIBjb1Yh9APu
d+ok6NjXjF4hu20qD6K3F3Z6GcUUaKk+iYpI0AtMr33jK4Rfw//Giz2/WhHopRhA
SGDFvyRJs1Va/HVmUJnJz7smB08YkXAF4vOQC2wi1l5NJWgo3oO+M12I/4Yj0ab3
p98ShtzO4m4lcKZjGAo9mQ4yYGrQdS6uqDh/Un5HiB0oTPUDRyZ7M+OKWkFfLraw
FSgCxUsI5el6VlqRDE3xAHqzxwZF4mISiZdjkslunKZ4WEiqC76TT7a7kG51oFAX
TOD5tbaajKU4mUtMvukxKDn4xEUoc2e3hqqlePmw4lBkandPz2jCcnoHcWfdUA4z
pZMhVgQWIyNXCOI40CBGTRNaHBUI8Mpc7hxZd8X+Cd1no4h3TFzCSG8CldEuVMIi
yvNyJZo1VLmScEA8RXcBzIJ/tp+bxPv5URgmNxiFo82AA43rkKh3IotfCSEYWf2p
uBYhyij+uZ5G30Oi8nhDeebB48Wi+fuIFKFfinBTrw3cMC9/JesnTjJi8OX98QEd
bnsrknyO/MP0sKF6RLiOxssy8Zmh0w9Ct2+6/25Emd/DgjrqCq71zptSWX9jNX6e
2+r2eR4vMPChSfp9NKoBUutm11TRVXlI3j62tZRQxJFTYcW0uernK4vxvjvBT8SL
C7ObF4p29Phlj1H5j5R4sXdY/9/SDtUU02BorPzgpeBqx4cnfNIi1hlZG3rrpeqd
9BapGWEwEgOuZe7mfmB8p+z6UtwP/+hjL6cwf5faEahkPf5gUEdKwrrGzBYT4C8h
7zQasy3cNXYmnhB885+gs2BmQHSRrPH1cwjjpuypGECgev4GzHHIn6Twm0RIjsil
WFUjYfJQFHAOGDsIGcc+PXmJfKuo3Gwh3ZXCW5ZFrxQaX47FgFCv6nIqQuNlAdS4
cQZB63C2B3zmzEkN3YCiJB4Slly6yTYPz+mZpvTjiewjx9zqk2LsvLxMtunNnNSQ
9Ym5qKZr1V1Gm/9UvCHybYYFLxi5tT5rq9WyhXGQ9vdwBI6BO7Q9XDGtQZB6WZKM
xQzZUNhbUkUQCmektIwWsufgP7YIgqrE8IjfjHZSpnkDXVLjlJ7fUHdY4XYk6G4s
quORi351EduRhOsCe7vsi/4+TxoPQsE4FMHIv0ZJx521/Hkmjcj5EOFTVo6P4Y9U
asrXAOC3fQRR5nLLDt0oefJok59bBh/SlAn+6KHEXOSO7iZrDO/zeQ/eJC5ahWTo
JGYiVfpGUO1gPmCav21l8YP4rNOqWmTPOr4HjQwouuzOh4w0nm18gwgge5NIxDzw
fAWfiJUEW/DuDhSrnTC5leGOjJMKYAQqtgXz2+AkeltFEhlDW5qCRRdn7PXbPYma
MmHhBg6jAyPCMAbP6MT/CYkMlmp2ETtKApM7n1rzyX0wQBXCD3j60eUEJ4eRV4go
IOWc3Ycl02ualBU2NpxZpYRuOC0S83F0jnmp7Q7AMMHZ2t0DKsX6Ad76Tj8AAwVg
6O7c+T89aWcQMbkaFTuVvGU0a2Z3v1/1eyGat0DuscFTIN4mLfm2EJjfX7vRy4Y5
eft62V9xcVN6Mvf1D83o1iJ6isXmczFireQ7pMKHrZF5Gn6IRVGjB1sFWJh/zcqM
8ppt9j0LKovnswd9haDYht+YITWn2GEunnKZWm11QNHxc3AOF0n1mVKPjeObydFR
qwa1KW3twKgWl7Yq6KJQcd0Czh0IB3CeZsT33B3hyOYcxxl3ejsviUEkRLvoAtQX
7G4ZLbFGL57Ta0MbJUHVg+GZFMMMEUrDohrMJom/v+gGyDuUNd9dxjFPRPxHXtIU
AOBhBgfGdEh/CF4L8Vv9KHZtmv4b9YX2er2kBsVe0GdhRC1eCLCgDS4HR/n3AVHG
UOlw2loj42yfQsCVkygReS3AjjpLWJ2lc4ycOHszGYXFrisS/aGmkNYyEdWOjc/7
jhjBr0ybGDepUSmaOPbglMgQ138IcMCruXF5XaIeGfQEAGWg6U7zy2XvHyPHTzFi
u31XDIHY6XQIk1bdLnzJTGG5MB1lK/mhPJ8aYQiFh7PzGtdk8LmUA5nLxwMKT80g
stDpS8RdBGMbgVn0KaeQPaZ2jZQScU6Wq0WistmDe8uXlRqKWazozJdXSlFJJZtG
l6hQ1izI8PbET8ivLBQ2dcMzfd1z83b8pBsDx0c6CRtpOdvdn8Gplr4pbY/AAifk
GNVP2iOdG0/nkefMwW/JuBupMFoflvV3MwgXlethZKrTM1Upk4m9CorvljbvwJ31
RLr29s9OzzgvQ9Wqc6gpKMpsTouKyUbychi5xcp3eaod5hmtjO3GpwkDpFp9DKy4
4Yl3b60Bl8n3izemSKbkRV1BD8EdlWBjxkZMwQN1m+qJ7W5XtEW2z6OpASCvypDL
sTVnbTFDejN7XZeE8PR0Hy6mvsXVrP8rsSedB25qKrhXvuzdKMG1JIARsS4Tc2kQ
0HzmBGsYgBqBp0Sqb0uHcOsbY79B2BfcixCGok/xkTGYqTfmv8bghW846j3XalH1
4+tJBQsOvrMOgo465KqQRybc0a85C+KZzd1fBy1wIVJaACoxzU+6rUlq7LsrRvNo
unJiOlYVQAndyEb+Iucvo0U52p0yDxMcGaegMB+XClmbYE+CRdxZybmVJcSLm+y4
aMzeNs7L4aOGRE3/lVNLeC7ZZ7c9cq81URBHOZamh2NB3g4tq8v70HUL/984/DTL
X77/jh/T4Oi3Ef+ihm1fBpIoHbxaGnRwCXnh+UpkIfDmuyPyathXn5MImGuDYHEj
XfNboU6eNQd6sRRC2nYglc9LJli4vy7rec8+DHU+TPvUK5FfYeQKhYmTASjJYFiy
KTHVyniR9lfIBATx70bOrRHLz2+dYbNeMmzfAsAqUbYGK42nczTLmOEVCPrgGoZA
qJHrj6u9Ly/2B5zhiMbWMtu5+qYlcDiHpLigXKobTQr6Ps0hqRKrpKSXp7jTZqD5
6P8or3FTSkKaDtMRpVPtTDmKAiFIDuew+zAdud+ErBQ70f+/AFeOg70q33VH0pXX
IPj8DRXiJohBS7Afc9bJeXnr4JIi741Mth+6VHXy/V9XTePrlaGSO0Q4WApsyDdn
9qm0wXlHBHnjdthUXg7OAIgyoUCVgpjjbkuGHPOU9J0vshMc2ie5fRkaeZu6zK4l
cYfFnifoIkM/reuOI8HscsGr+G+KvtqG1GaXgA/xjRkZKJW+cUYgHmGSNeRibdZ2
Z5lsbn/kUHRxTDgvkIyPzKl50W2jOm/dRKWlxx1yRm7+ns9543ESZkSgALtuR0g6
UoSuCpqjvwTL1t5mtv9Yg0H2MvoupTOz9S5JtNlVRFcgi4dJsHmXcEUEF6l66Tx3
Rl8BUy6OqRTNxjZYhA5fFbVyIPFQZAB29IIcBYhGlg5c8dMfAcEArNZsyKyGgVnq
cCixBwAoXIZgD5FNhpyfEKJglUkVITuYwi9n6EFg+e2Fg2+t5iBet6iMRi14l/Ag
YOHqjrgzwApoXOVadZ863PP7zsTpQ+lHxCyMZJtfwgn/4p9H+TM71zhzLvJgr93B
K6/jujDXuo7ONbKoVuj5AND+cSGNP5eMDg1s47lToROT6iATDN6lkRvNdeqpPajA
7HoB4Yxv8lRBPLxS9ETedNtYwmdDcHr65TWenIvWycyLavfaaCohwQH6cpfQSs+7
JRqbjZcmBD/hAEDOZhmNBGNICRMYb4VYouyRerVDs984cZ5aWX8VxARl0YvuGe9s
bSNT2zxs4QpS+lUUE6IsjQkiRN9yxJplS10uB9GFnGZnUMn087ucYgPlwNyMpbBu
I0K/0Bpv11cUCpvTP9k/+6qjSwdpjraqFcFTEKY3QOunKsSClBcqJzrd8lPWflml
fw/BjXysNb/DiPFWsguKikFszAsCngxKkLRA/+BrnN8dEMqXU00MTnNRqTRthX1S
Awtt4ENi2YxPlPak2yocSfHrrz66MIXuy1/X94jRKKEnkCHzEvD0gqTiMRQh1tE0
dD9ekUu3UWyo7p6fJULUV+4GofNdIvnSfpkbUi/y9wOHvVD4BAyjli31SzFb4SOv
GzhdRtj7UCg6h43I/X6wAGnKCRAhIXpxCGuVNVzAZ0mIOeWTNrL2DXorrAbBpHEk
BxCqW/xLt8cOSbmPloRr0SDNwgwI2eFQkBlD4I1Qtsm/UsKK/pWMG+LzkoIUuzLV
3Js6DQBEfl+ljn8zskbrvSZ770uqi/7az5qA3E/v9RmPRyCTKnZRHJQBRWMZ3O3N
KZPAmuC5YQT2khecrTb/wj8dIbPnfqlquc4URDPPkEIUDItxRPmqbYipyVT4h4ar
tHVq35LFLu6vBI5W5VrMSSrziIPHQxsIIlI3vDhDcqwHhe9W0M1R2dyIri0o8d7n
m1HFtZcxSys7gLmamZsQSNjKWRLqk3/I7cx1FfjVjNozGKAO6oB/LNyx76OKtNFO
jVwF1lQdQRFMWwQaFu1kbZiQWJ9apXYkMdHMj9Lti/fr+RCXJ7m654bu5SP4+7Vw
uZHYGPZ44sf+E0n3YIUbyVKVdvWMBaRVWkbj6B7HqODxK4KXR7vcSMugpJyyAr+1
ID5fyXiTcTeQ/lF3WJIuqJTnaL9RUc145HBOI/JNcFyajuoVhXT+9kzNJuRXN96F
C9/lubzD5gtFyiIvbQ9nfW51lwFgkpxewA5bGfP5wjQ0TwoFaNtzCELtJUZX8NNc
R3HhLW5OJG/tS2KDW5sUlBTNDRNSPQe/OyoVCIySOSBdM0Q4OnxqprRPGoIcBx7m
03aM5+JhNN7M76yc7+Ba1pEKPwfgYaidFW1BcH4YfZgdXarn/fgs5ycMrvPZXUSv
km2iJ9B1CC/JcMa6U/XqZ1qrR0QSJu3nXr6QRoVaTKzWyvjjn4RYpEuM9WMc9ZjB
wu5utgK0X34lkA8pHYIxsIhkrdmvRSyj5a6owZ0KdeMtjD/s88INSHNI/b74WnwH
QA/P8t3YynZdztaBn9MN1qNy7eWzm9ueW7tS+Xt168oo197PUOkW2JI/GOyUwLPC
FsqHOyW66C8hK/72cj3QZkYOW+na0cfKXWcH63pMb7E+nfyAxDcRNRYkYCt3ygSn
MeCVOxXdwxSSZGe8PibgvGTnvvaOiSOWrUcJHvtDUAKF03UOFs+b70YdKGlM63bt
mVd6UmfX00YDiUuBZ8WMo6+Spd4h9xgKRlgquip4KN1x5RANNJAfyg0BiV8CxQDD
oVVm34yk3hIzANIAsOZu02UA5qBMc4XkvknHPSxUPGLSQqI1yI0tqIdzCn7FjfCx
wB4TWBKRX9Nh/3ZJMUw5dOvZ1UZgZyBQVovIXbxQ2zyobCbx/w5NPeC7iyDNI+sK
c038Fe1xLIc7SL16C8wIoGQ6/IxbAi6gYHxEJ5dEnUZTullqpAjE96Scuf21owtj
CaxKutK/4pwGA3qNQRu+t8tgU/RjCXivCiPviYXwQueUlK/SYcWKjsgHUL/g0AaU
y3i+vmz0BFb4w9/v9lhU0aBxCPBfSkDi2rZGD3AEPxU3xTTmGPD1PmIJJ5Pq6G1h
ItIep2LDSpQrBftz4TlkooPoiAclkQV3DCcHUxe6LwveIKhJUNBV8pJWn7Ns5b66
8Uqo6WwXGW/A7VA1AFIYX/LserNxMzbejud8UKnwxtF+XhGbw1E7KLCwbL+h1+ZF
O++5qcQaQYZeMacp5LvLALYqLwcZvpFV4OINVrvrLiLa6Du7OaIo7Zn1gAsXSR8V
//Cz6+/Ggh+ugVLNJSWUjx6404USFKAx1nydBHUCclm4UogGnuwjzKuuYD0dvcbD
UnDo+Kd8Mas1MZCpaKq5KL67zUtkTO7i0g7kf7GaduAJHP5FGqYrtExsRJ2tt+6a
M4ohqXCVhPZ8/r8Q2ZsG3I1smBl25TwCK6M1oNVC0FlrWWMZdBkSDVMuJnqJdlCY
ZasOkB7LmrO9I+BPv1sOcNnMmhpjLNLWxfYjjfOI4A90i+7eOUD7CiDke9TnbuiE
ozIjYtexTvMrz2LuasKh2vtKosXyBR8LFQQiLr0qgUdEWKxtj5rg722+j+1Wvavw
BupuxChUt2xn+/5V8BXgVLaajfyM5o9TM1BO7pKE4WExQEh2oz5OR0CV/QZPF6CT
5rFvu9DaA/d0or8PQPZAgmn1O1weIrn1ndhkpRbbJzU4edBr5BHF64ox5+HisoPV
kj4yqnfSoq+BIA0lkFJccy4YPxzwPUMlsuzkWld7Igb8/dxlLastQPDxFjvKP2A4
U7uKfdS4uDapgrnvoAc7cBMVFVnCz5wP4w0p4V+75h9IccSKaugpYCgzwm6ZSeFB
JEBJXHwqGk3h6Vop4xmCo8CfwwX/kt7c072Li1mq0+bIMBraeIdWQxCkG2YNIJ60
vgnDXWDq4GH4edsj5HVAa4MzQnJNiKEOKIg3m8Npxn0ikC0YhC/cgfpFb1kdkFbF
kOobvXpP+5Tivg5pc+Ug/108ZhvD/Pl0oAzlN06346k8fHnkbbovqjqLsOHw7hom
USG6PlENjW3ADgscpY0ahXdxvBAyDlGTIIsFEjhQFQUyu7D1VDcGd9YYZiBTud4j
zfka3/6QlUyLmYIQiu1+o2eepxQ2xGvxsnH6cO1OQA8JnmT1BAT8nrp3lWBdl3ae
xeFYzcB4e6czCilhOsO2va62gRZHqh9oxsp1DxL3ZcZ2tQd/U6J/K6NmL/hCNEvg
SsLnHzO/jCGgE60vwvn0hX41a9gNUu5TeWzQMYPPGsMHjBCDA/YGFnb/EgOT7RXd
kJRkjJoo1BJtkVev+XkwMrPuGzKd/QzgpS3zoU6icDk5WkkQW9qOZ+Hzj4pXZd3a
Jq+y5S9M4p0uViLIAMHWV794ZKMp/kDLEQ2ygHL0GEALNli8dGIl67MXYlZVvKhJ
OvqEPVw/8o6WhF3DrcDoXhA3RH+bU3LI1r1WdFxHawoY+RJV/vu2a/aLzIRiat3E
E79KuIHOZqKZ5bgb3lwd2K3r/tE/Tqu1HmjVADHDYj2qiH3f/Xpre9L0QfLTkJVK
MnqdkjWQ1GMsE1xodRje7tHDGv/sTU1/DJsEulgYkRMXAXpUm9+5Vg4CR44lOcGG
+RXmf1hnO3eoOUH71ZrZOpjEaCrSOGVBj2SwEsrmUckh3+hH+ZZWCADIk+JgFvVk
kQCHn3CIoWyAxRMExEtbHzJYZ8bgUk8vLI+dv0OhhkOlUq8l+7Yy7N/2eeSX9VK4
wTucOxNQs6I6AnklejHJK/5NYGZUIZT7jhE7hAGbfMo2JBy3PHJGHgc4oGjSzwPp
seFsAD6s6c6tOU8/jVc64aWt+X5MglQqb+/OYYaiB/pcSvWq3hHWZeGh3AtooKop
dfUbtYQiMQt/k1l216Rt9Nn6jWuzkywHWKs/sXLUWoQwRyagxu0vL0YBcmRMkuSd
N4BDo+ThM3PvsOKq51iYKUM98rJH7rCbkDmKZn/9E96lgJ/Zl/yJ7K86BuCAFjbA
yVG9fjOs1SF2BjVLTrV9IRZhaCngQNrkNWTjtvPZbUu+PeHFSYdSN7bosYRufez+
fBIA6Jno4ej/9UxQtDBcZn1BMnMgHbI0blF9yAfBPHg79q6WywlBGDBZPdSyGe0l
fbz9FA2uvquFQdu7u3RLvFfPbNVU1ChnK/kLAmWX6oXFy8mkr0Er+sBA5+YZLInX
SlFbZBAnzXNekyDu7VBGJa26CBzBJO0eEFFlcPXagISB1Udws9ixKo/P6Gs5M3BM
eJ7uLu3SNmcOFr+UFHFOpjLqrYnxhepJcEPo6cBNw3tS/eBx7C1346DTyBHTVXku
eqFKnnCZU8EOWgw0Gy+n3s1Tas3UBReHPBeZbJEZd/rV3va4pi8ACR/k0+ZxfnAP
1taLBpiS/Q5tMAnlr1cKry/huqk48oaoTbTnnpwiuA7YKhFGtWVpklKDd3zzKw2y
cTAG61k8WQdyXtmhpMrQbY0wj5TRdUBehtqlnh+Gxf11KVBm2gDlO6twDXIeZMHC
4Xci9UMlkv3tsYJGLVdw5iI4JsPbHbm7qqGSSL4lQEY8E3XNeuzQ3Hu73Bi8unPg
tXrNlwPFDNdi7jMELHZmDa6u9ion+uV1CH/MilN2dfRlBG1+FMaPZEiWR9XFQy77
Se85KQqFpkv438iqJWWYkNSy9c6niE+E4C0fl9+VxxpzMFBN51HWooIBsXHbJNru
qoLG22hYSEcGawApG8vs9HUWz32BR9eFeya0Y+c2sY00zaQ+PYTKlYXp89xBZokr
Il3yW8YcqT5ngYkm3DHlYCC84946hQfDYvqwul/szezuDm1fZV2BaK5CnJ72J2So
yiCiOAmDbeQnuSc8TVov/I6F/8bB3Q1SfgTdOb+IFAIxHdT5C8ocVXvzkVxlNPhz
jVK8xMSYbvZIoTsA87fE9arBu5+fEB7nJbr70+On3mUyjeEZ5PmnoRrqO3yili5l
5t35WrCzoLoSYnUirVfUU+KFQJMFtebotWYPk2/nEA8UXpnIzWoeLZc+PbRHuO4v
VXsRzbGZ4zHvyTZBsmp5fTDv8KBOeVGcm4lWepfSYm6AUXYSBI+bF8fTY3PIgEjN
HTLyvSRgjxSbP/lsH++z3PsdYNOHEfRftgp5msEeiwTNPwjuafr1c66HilXjvyLe
Ew/fXXLKtqnbAmlbGVJ4NNu5T0dHas0caX9lg61DxMeCQpb+6gJ5mVXyTsfPmFLJ
XU9pOWFnmKRNYh/NHr1EU2fsv0NH5SYyYF5Xo696x2cIv65mBI1ZciiROrF6CkQg
l/dwvM7T4tLMF54/EH4iqwUCUss0h/fURBD1ViCwgBtdTysWFT3E3UvqkulB4n4t
zdfHpYb5u8bqddAwaCXfet4MlAYzH6vbFT1Sck1VN3Svw9uik4UQjGTJEVK0eULX
k0tz9+rozby/9bgiHihOwFMrv/vc6gOdY+w2ZTBGfEb9TxEoBC6AHagerns8n8V3
6qP+FqLuvA/wyqEDULQArps2kzwwt4jh061DGDmB9Auo58Xfaax6lsLKTS/hxdUM
23zuTF0ib4Gro83fe+pHOH/Dv0V9Cq7+kwL0LtY0M2V2QTR5Dx7hC++qty14Rrbj
bifvcTddSwmMx2vlzpjJh1Q/E2wulJCny1SHLaq6YWSI3thoWclJBkmXPdTdbNlf
6DPlvOZbcfWDqj23SlJxlmPu401+0i9Bu5mL5YCSClfILeoHvo5BIKodnhPNdFXE
Dj3ezwdKI1jDjgH/PrWbx09YaRvmqql8FzFdO5iXWyO6yuyPwUMnKWjaP6Dbwx/f
HzlXahNEnEdO7Ihmwp+ngxKH5ZQ5c14LBspp/anDenFaCUBYebDRBnQwb2Nc50hQ
zms+rXnIE3K6NxXcsIIecJ+FhQ7kGu5cYaCdCKkjr9wsaLVz6DyNnHCXRT2xwokT
6DdC5Mp/QG0FDWlNWH3PUzESqLkpt+0tlVOoChZIRyFbuZYxw6L0YLI7LzdmeLqv
plT4pbc8U8DsMPw4W2W5frhhq8zr6Fi8jRmxUBioAtVf3S86RrOJFioNgbz18dp9
a62GpvZt7i3fExutzP96hP2JM3LtQ928aM+rx5A2qfdMN2gEuh/uq3NFTs1fDztR
sAzNwpjnNqIlSs4f2Ol5KkAThbXfFHS+NrIgXHkwlHOcvYHCq3mSgjzDYtFv8PHN
WJl7Qnphge0tmOaUNUZ5UfncPH+PEV1gBeX92Ee/QSh5zvcs59LfbvMKS81WpjFo
EVnfroRs8LOR+SEx6TnKXRhRbvT2Wi3zPZaeyhBWeOsAlQ7KuCN9chgjC+OR9hlf
eriIYtwFKxWD1WP70p2DVrgm5z1z97gfmPgcWtqpWtxiWxyMrBIPuZoREXu12T3C
/F7C2bfnAJI/yZ/FvyQw8PpXxq1wpfQZCfUesJkzzdgjI1NC9251lFTKruY1sv00
M14Z4RR5VV/mluvJDb2aN/F1CMAniqaU7DTmVmmyDxQuRb8uXI0qexoc22ql/pVj
qRGZWsQmLJwMOIVygg9Egz15Prhmz+72C6LCq4eZNrNprd/B/OCqiX+dEmc6ZwB5
Xb70AygMdemoXvZDzMRccVDkow4bA8gScfQTTdaA3yOPb5ZnLHXSe8V73kOuOvOC
pg88azYk8Ha0w/OqFjU6dugzbJxF9xkMdRGHnoSqjcQccDS/NpRBzJiiW+kZ++yI
NlE2zWWB5AMNzFnn9Y3lmpa0QEm4jTET3s5ZtyTpuyOhcN55O+m+nfqUNlmZDYui
F7wnpYy9grfo9d924rcJ3gL3/nG71D18RJG1cIGurynPNd2K2XD29QsQolzAJD8O
y7Ev13SSnPB7BlU/VmeoQ+Q1r9HfCN7TMXsw+nQRfIaNCOHxSsOc4VEZWHKwc/v4
RcC1Vfctj8b807vNjl6P/OjzOBC98AOcwmMSQ6Yf78cSro5+uhzlHKCJpx/+aHa/
zK1Y19jEiq5Vs3CP7+/iQRMGBOd3qTc+DMTXgYgvdpAYRng4ITSZDD2x6wDlrciO
GCCzHQIiNQUnf4N9Yt2iyRQ9ACQuLD6xHx0+4TiSzKPnl8C7kAclPm1WaeNQEFEH
7mR/970VizaADd6n4MEX5dj7xH6MGzz/Pjf1Y4GYT1quw1GfPAW/7V/3wq1WpBJo
6cRFEjn/Yx/MjyRcYa8WfTjGoDy0MgVPkQMwPDAmJ+QEK4noQU6qjBWBHbojQHcC
yu7XZRXxCAihHWO5iIVfVyoQeX/8/QnwhnXaVFKV7m5tefuJkb4oVbTPOTLQa3jV
HTNLqf72Rl4VdkjgR3xbpyQCFPWXC2NPj0vyKF1TLg567La4+Ns8HJzwcsbjJYNC
CtUvxGFT7xOYQEMMgNDroPOvru0bI+eUbCq645SuirGPyz7GYd7Y2fWhZz4FM/Hb
dK8qccd8a1JiHnYDMKAf+ibQO90yb0qaVJJ48iVMMswOB0j6oMX6ZSZ/zKq/eny2
nevaDrmYqKO8y0bDra5BvBSDrcKdvZRHADzlebwhGrYbmNDzovlp9DfKqP3/RfBv
4VyQxemLeXHvf1uaENvU7jchzpNqQZBD+wcCvrILuDs2+/a38GwSNUhysHcagOIW
7jqvfkGp93WOt+Ichvhf1pt34xwcG4GLBsXSgbSpUnI3oaC7Ka8Vyqo0nw5xp8L/
/91TjKwnOoKMntFwBsePVoZyf4BZTt7ScBKN4hZFqZcVEMVqxUkDY+xwdMD0lJnQ
oOW/yXaxTPiE0XEahCc3hUo5VSQMFyAuzfUT0MD1iN4/JBP1Pl1ZkOSRBjzm6AVi
z5uk5tfLk3wUYC+UoZbaMYkr8D7lhQdiXUKn3A+q8WyXSTDOD35hn4J9nwLEeXKA
MvSjKoRGbHPCMC03lhgonVhIlDyh4XTcQZcnQ3STglcCA96j1gLDW6adxtXyWSY1
Jpz0/PqgtaR5jcfPfAADO7zYXgpfyX28jLrMR00Hn5fon5wfmpvOcnuUng3PN0fl
f8NPLf4hzD+eQ5Jt5bP+gPHRTAubeP0n4d0tsupf8CSgpP8LqtE+o4axaFmoTE4O
QBo85rXqJome7vcQF4QV84sAnXYdw1d2u7rKdX6DbBsIg/R++pOO0BOfdpbCkSwY
uzSctmhuodJP/uhELyED/JqbDRpie4KEHArT61M65jZpF1OSFBdxSzWJhjl0oZV6
Rw2MGquXdGxbYvCXGvXcT9HQiSxYy7UGFQbkn7L6qtDGpkI09eFWakY4hHzHHlrS
2saPPHS+TYhn/ZHTGHdyzL4WwQnyV6Lk4lnyDDJBOE5kBIv+V0XCT2C/Hj4Cs9q9
nXts8+1rv6tdb7q2rU3lddxLEP0UB3nBY8eUo+TOg4JbD1AXKOet5blz5Rr9y931
XpIomHRpm0+m8kkHilgWJczLqYYqKULQlGPM+2jF36RKUNYLosiMoNTG1tEuNm68
IYTKuCLQpL3P9hw6MmOW5UE4fKYIIlobGc3VoQWcAURc0dl/s++Ylb5ZQHPg7JAM
kOFBWJ1G+4SYEIawv8yImt+pnsbRvwM2STXqUrzlU0McyGW4oFEE1Co6gClPdYK8
JrnmEBKJxDKelD6wsYVQieBhey/uqRAfuNlmKyHDfKGJjsC//gxOIcviOHDs/SXD
+61NyCOdWh4Fw+cnVFMEx/J3dZf4rJVfkl7ntppfbOxQybSLFL7OVVebaEnq/vYJ
PqQB7WQvlwKRXgGOlQ9yorh2a1vW3WSVmpu3LRfnHTHx8QngnMVM6bhbwbUUkFcY
4pv517DVSv7zNk5a+KJZAgjiW0eyL6ymBRZKwyd3e03OovOT0FqxMska5Bq3eWMV
n1Zbg0AOJrSgym/EORLJaaIRXM5XastRE0w7WozNmioFEUvHGoo1rMDhuwWNYVKA
o+QIgSz9h39+JPjLFNKhVl4xUoy4diru6wVM2ztuPmIWthdTysyeqCxldk/1KAF8
QGBt4nokHP6xbzrfRrSMbo9WBQMaqpoz4lR9X0rSg+eyOte25PJ9ZaFuvfrW9OvR
Z0w/E3H8SiWyCH6vuEC3T5RvDn2EfrPrhN6vVLUKf9qLysC0s2+nXqd/rIAnyURy
qWvZ3uwTrKCMDB2p1+x9U6XEhsRu5DsBzBVX1s7FEzA06SWKq0sax0o8Ko/0jfjv
zgfnbBLFCGzhlh7NiZqNWHGy/a40ALgo51OnpjE43uxc37MVmkvHuyaSi2FEQ5ls
8/lEtRvXI+aXK2ViCPMZK6g1eittJMBO+i1nFWGQxgb6qDz3Kjcn8IAdTtafReU1
g0P5AASEV3WpRTP6WpK7wlVhGTbn3QXscIkXIsN0OLCST/etLlQGJ6Xyz4rPP/qN
pLtD2Mr5MSQHB+eEFrQDBEtUFU0MdmMlHN7BBcsDGfTr4PPlXteUWPXgHwHKbYt3
R2wI1veBlOUjc4hVAnxZkOw7tt7a0WhaekuD2bf8BzmscRUgwxv7MYpkDrrKlAf9
GwY/Hzur6crf9BK/nOF595XoXhtWRSrDgNr5x4fIHKlDsuQTlsoNjlhV4tRrWK5p
pGmTq8NXQP7Rg/AjMfxG8FTxn8vPbxmualoXLHxG3KFq6lgTnhe4xqFaoaDINeFS
Z0oFEdvNG6Vl5kLv8GVgt1b6AGbP/NmwEdWtSES4/Lx24A2TnlFTEkMl+DpzUkUm
gdHF0wzBVqLvHV1wmy5RAahvzQLYvCejH0RZLEAOTfQnoQbkEx7xL5Xyj9xACJhr
G/sDfLhKAHdYWVdKGSrvN8wJfxmhffLsMRvIqG2gVJd8vpl/skx6Ud7y746w0RCM
5IqMB9HZSmJxQRqtp5preffjG5uZ2D4Zpzu7o3m7ehPuoJ37pNbVfBRTUIPr+vNs
92Jd1FB9E1Io5KnoPQGjvXDxlb0TR5BK5ZpYLrm1B4o4pjF0LG72Lirkp/rX8f2C
5ql3tNthATj+OKrzOyXGfDtudhlckn1wo0INB/S8ldZdLLsI7D6bAiKzwVTn2a7w
KXrYlHDTYU6BRPskxxDVejRzLXRtFtgPWfk1U1YlSyVk1YzvLHeBtqgta9wKsV1l
Q5rBJkqMlXPAY0t2NXAuzFUYnZ6JWFrUN0L5Vrx3RJxbV56U1eyUeRJkBpNWQa8H
v2YkTd1ISD6BNLUqqJPKNp9fquv0sWJRCjeNvaJrS3gw+Qr9XctRHy+odhLMUeuP
L+xbdVj2x4BPzd+A70YE7iW5E7hbC8OrMn4WnkeHOGYZNtWGOL50+56yqxQRxKdq
yJNg5K1hLCBlGDQkDjiJYyIvcLcK6uHDgNj45tLQ8sNnJ1JL/1iU9gaOVzcZhDdK
Z3i0f8wUJWdp7EGZy02zsx/yfW4xzeZT0ype74roKLwq6C4o1fc9Q3i7DqjlfesN
zSQCtkNorWUy/MOP4VvcavGRjVm0LQYT/DkbfxoXgEI+bLLjVCnUQ2EnHDnyUBRu
xxqpLf1pSm8ysYLiolY8DD1rrKBZ6UfhyWzKTviFMjVYzIYmfe9J2Grv7OiaKp7+
bPBx2EJDw8X/65eIWJPnHN8dTXsvDUaBlwyjYz74rStZb5Hl36ntEDPoTw1q0iO4
rsn15D+mOPARPEIPe5ZJ5yQsPT/3zkespQnhW2Goct7CyF+XRXmzIhBDG039xHZQ
6m4ZjkXZpZKr5CVzGFW8Dh1Oy2Z74i/0skjpsBZhTymYzxDWqPfiXGATW7+uXFh9
FCxKdwP3sqVhMBku5cohYz13WrZrG8kXQyL2me6EwwFJBAyvAE+WhOCBjaHkZ+iw
niAKQ5bH2KwwBEPAmB52rB5aZrfIaT3xYt/RJr2JPdHIeWuIlbXGKo48tPLbgtN7
XpIHm3UGKSnJM2B3xSrPoguSNeKtPo4ShpfGFX/vpFW9i68Kj3QNp6cjr5pI/juC
ncxwCHjADOYEno/AbUBhBYidn4LABTDzqXA3trraGdxFVNTYRp3zIy2xBJIuf1dz
QswyBXPyjqlWkrHgjaWm2sjz8JoRftO8coAca71pYVbsU0KGUKFXldjnn0wKazez
iQSQTugX1JqBtLU1pHzFlytmoVOnxu78VShFIhE71JwbeynMazv2woI0vC9tA0hx
wb/l/uHGLPXx2syOWaHaI71Yut0/VmS69g9/eVog1yya06UgzXU3DDOk8dnxdwNI
1hxmQ/FoSrwrH8WQMHnA0Sn7n0/6JqcP1U26y8f9ahI+gqisZNsPBnU7Eeric9n2
zVSmeeG9MNQb0/uvI8HbuCEvh8fySfV7b/52CbpogABuJOy25UGc3+zkrLk7ebRW
UXcHDQFnamVnuiGjP5avmV2GWP/S8VIHh5UYlygNbcS0bm5hdalN3+Psz9trR0zk
5CU0ppd+ycxjxCDi9EkPEsYwETxSx/mS5g/wKUYKYoqxSMRtvAPpup5+6iqsh0sz
8C5JJB1Wvke6tLvdu/2BaNfGOHf2IxW3VsDKIJYMTnQhFiakTuaNSw9lr+SyAHx8
EB01i9sCrh+68uUFaRN21LhO2VWdW7ElgyiArbH6P7+xbgbhezOZlb5UN3qRvG0e
nSr7GmhK+ycbLsL2bl7PRgsI1xRQFRMdCUsMlHI+UXxhyIODhacRw8xcdIZYCtl/
I+L036KzeZwEO0r+/V07r7k4cB1BUjrPXlskiIDlRfXHIKDwAeWKMc8bhDkfRoph
5LargLvhFv2t16NZ4INUKPFamaXJdpPe1UG/l0MAD2UYYvqBAsD0yx1Dr/Gvlqhk
yr2b5cicx8HznMTgVXKXULK4uReY7+ZlXFnqHeF2it3fZug4VXFJlnENM6ypEJRT
/p9oodoyO7IY1caw3rVKb+Qdx8Q/Cl9CyAeentpExr5lcFGpAUmG6AoondbwrsZG
DAcJF2TUAah5gASWURhYTmcCOCUvQGGkNidf8zqR/e34wAaGJcXoOiGWhykk/AjH
3k+7lakRH8EGmOF8RwpaehA0J26Vja73Ksm1uju7FpHi41YpSdUW8OHsgmVbCjjY
14PnkTq7AswYxalYGp5NB6pe9A4RVIyoUyxpPcTWjobe8Wv4D5crzEEmByJ+rCdM
V8v8PqVWf9j8/kX86UztIrtqIB6vPbquI+E9t/H6/yvMfZwnKeqj63ToAE4PND3c
78Z9PznnkPB3GUnZZ073vg6JSCupDmjInGuiRObWEzzlfKEe31GLvvibQGzmcoYs
KutCHxk2Exa4lUtr2f3/xHQWRvABHr1ANy+ySX76zW+onoq7SaV649fAAz66t7se
IaUFcHyQgmzaq0URh1x7JYxPICIju8LvzMMsZXvnmLp/H1UjiWASgmaI4G2T2nYC
Jmla4PRebUme5/BXHY7Rql2ZTbkSSBLB4lEX+jDuTQLjyqM1bWvPZNqBRwSAxwB8
UItKr6lOkZI7PvmnaYbaI6LjVCOECqtJbZcBs0YN5Psm26odLKCAwzBhCnm/qz/M
u+e95U4aRQaIJ3wB74Wkofh1jUczKpjFzJofLhm3UZsM4acV2PCde/AcV+z6BUYv
KoOtA22DbB3IMo2RQF1Ln0Se3p9jZMk+1e6g5f9JyfyULoVZMcONpf+z7B/Cs4Ss
v/nfhgUtLz0zr8z0GiMdFsuDGCPG61I7LDolkWy/BusBu8+jo8D15sWMZRlBQhWX
L1PhEwI/+DEjo75b9XkfaQ6mJIMqz2pegHEGQ/0Rjwpmjl5CT1AFJPyZuqzj1kad
0MYOgbkKp6qZy6nwImNWR7UI1wmhotFb9m3nipMzAJIEyq8nZJw3qAEcxElGI6qC
xzFjmMAXZ5PmbxuXwd1b8/uob1lF3+OFfJKgi8n8P0QDZWtnEt0bGxpBBI73OMjB
ao/KQiYPkfbnECwvPG2lbdhxA9NsDwXg8kLIhkEKnBMgVX5sWXXY9iS/tep0O9ZZ
Hmb+PuOmvcgMDkYYBk7ExDQmvf+yeyYaG7dHLLLUVBuVgwPgoq3UeSWiLiSt+YLD
R+JBp3sNGS2J9rhlkb8kwAmuV4Unhy0Nrlblo3AghQJptF6ADZxjWvegGdocvA2j
RCpSuIPzO0Er5Vo7b9XYG2+PefD/P+0P2X9BiYt1AIztPhOv3R0q4zyATpM1Db8u
PxMaudxTnnn9QLe0ifqm9lBiOodSNpjDNk9x511V2drNb80BbYxUwEIqDttplomj
3XT9eRX+7GTiIff2ikB3zprFzYpCk+AtARgWZ4/gDypTmkFYSsejqKBjtbqwHIYR
M20XtHgcOpN3V/TUpz6c8MakDdbcHG0LGv7uMTIEt37fbHUFxM78des64+tUl6qm
N+XhSH5gPZ8HpWwnoT8YduQgxfTF4fBE30aj0nefVJlDlbNxXqhJ29e05q1P3miP
Fc7jTSr7sLLdwajLnHl9/Jm3ZFgLUAjqNFZvlN2xRPCkczUJyfUgyOsvL351BGCk
xClr0c3URV6C9zTQlJKLrx2EeqAOq6Y6RyXAsvNPcTB+iDwt1qx1RXBHRlIpNFc6
8bh48x3SKIxVwA/4w5Xd962bvM8+ZNF8N25j38xVfn6l3JzvG4mT+UFtvEELlyT7
JzhzwhLIIoCp7iOex5PPjpcFIiNGMO+1itHX/Cisc6sEy4GBm8vuyaCaxLjHoc7Z
zdiILPFciSRFA7FrpTcR1WIluTuFSjYDARxL1viqknjZfNr+KlCcH4xxaeu2SikZ
/a/riBUFYDRuyP9eVvuQ1Th8u32gTLp4r/V4dg3oaDLtCO2VTKTjI1hIrdjkmttU
N2vkOAK6v+PiWZy9lN+8nsI3NH35KDTdKAvWRHRVBrt3gS09p4pLnQqNt16yHAPQ
I7Wluwwj3uAzRD9ODvMRLYETxJRFvDU5miT/H6J90TBTOvGMbRSZU3+DIWmPUcCR
mhvbDfG11n+X/7s3RfD1cjzMvtYH0pIU8QfToPozWouYq3oTwaUvD4vBQMHr4IaH
Ek1xfeJ6EZMY8NBaP197C9shMdQpvUjIXyVv658zA9767mLd6fKJ+CSL0P1mPCDn
n/Wht6H0oSKUUMRCBg7WiNAfqZvhx44zo//AeWzgXTwOmgIiqVCedHRPq//kcWq8
//kvjpk2B2xRCCRVysvbVpYnLz4x0fUupRpuWo8JrnpQgocOvU2tdbAer4N4UX8p
Ul0Ci2gp+K9G1xsstf174VsiFA1VGIQ992o3eThHWZ9K/7agIgEg8zuc6Dw/2rTV
sWWXfaIj+7dBOh0XTyUZJHHI8AfM/55gvZl3z2mki9ho92cUIgsJwBQwM8l90RZo
r48khWxJiFgeQ2c8lqcqv5wz+pRyR+x7YJttRF+cB3lK7eYKS5GNcpD8yRN2a21a
83Nxo1dkXcIZCFi4o74lgj4rfrseif+DY3tXcVdnWkhbgiY8jlsPUbog60VhMwlt
TC7CGhn8Pk7Vh90wn4xM4kUY4a18nseh6qbyIZCayoIDTQWuaObETrQq33NonPOK
pP3fNNXIO7aREUZ0A2AOoz5EKJZKtmORW02jy5ljh7OWVYxL/i/e/wyBl7UlrZwq
lf6V8JOEmvoD5/TQEZk0jcqZUWvdI6hu4L1vBkQVNpJ9gdz99he+oR8w3wYTOMR5
JPM1p9cEuqzB3Opyt7DfJIiS4AdTfXdkSMdEnsRktE3oMqxN/iT71s6CVyq0yiWP
PBmzAeKpDQ1qsZQLy89FMBoAiZb8W/8t2R0SMu1WoccNLkAFueKAm25mshqTG3Is
W3i4rBXZBBceRWiC1yZ7kKzaROp8cefjBMj93/8M2xk0CuLk8rrI24mf5MVyjqz6
zp0iqaSZEc9BvKstGBZHWrPBlP+dND545l/7aZ5MN4Wii5QNr7dQ3a3dQOECW1zz
raT7Cdj7qtfDGk2PNI+3TiuZeGEd55p0uApdA/z4ciOWUPiGCFDUwMLWG6cTxwZM
vLWWutELYpa696y4tJi3d9UYzwvL5DWeDcjXwNdb0EDkdjpovs1lOPGo5vAWca/f
07fuFqeSdGH3vgYHYIkHipIXbBIL3FJ88AMlU4phYXk3YJPTpyAv6o0DSpo7AAWu
RidbUJHeOkCQS6L+XPyn13C6NpCzPp0A7nriZVzfxiio/v0nyor7oWCKg5cLRTU3
/DTT/KyA0gnC16nuATJnKC0/BYIWOVn7m3O9I9d6PFV4MGmVziocW6cn2SJHErJq
Uh/2o/GNVygDN5+9oqNyC3FFOzzirPIZkXb4u66iEzidMdUfJvgkjNQepLLbGzpA
Di3mHK5ruukDQncRbfwbklOMERYwLleU2+3gunMWhElboQEShuMmHKC0+fl07IXL
HZc0v3hg2PHX7HdQdAplnir03rkapFQSjMKg1iBFhwrrLZ9Gm8rjJn73TlOoOOyW
3zEPdtWwVTJhyIGe5aTwAN8+hTTgXgw08JSYVabKoERb3cXWqgzZ2A59pwIrO2sY
w/guqsHmioYl2fznKHdjGiiHlhFAp+T+uSeDHHYj07njQ5rKBgT5y5IQCFCLHGKa
p/8vtxZvz7mdkEjqyFbafDA4inFohbnHd47mTDDHMy1SddfayfRMocgx6BQdn4IX
/m6mDdIiNRkrD0my6uORs+pOVJX0Vw2i6OZicpPL5h+Q/6hmhf1MbH0tQBQN1ntO
sSzMZS+LdxamNawABI75FdjXrlFbgP/dB0OpMjsheX1JeuTq/z/St0HRgWYUPcER
Br0LCR8PUCZ3Plbk5ZwltnRgSnVzVIovmLAeEaS4X7lslXFHD+VGoHNNfikItG4J
ofk/E7ixlpbJgUCspiW0cc6iFxmmh18OEdcDiYUNwJBI7e+n+/viRrt+WApHJ87o
Ml8fiwcK7uNbQ0aGBAmDVHsng5Zt0XfOxTE+vDiudN1W0+Qgp9h3J0VuVnNUE1sy
AeK0/fF2X/e1S14gv6LhvOFejJ6HxxZrSjUvoiVLMXQjgNDQLEQGRo7HdlLmEjxY
VTOVzPvdQ69xENUCH3vocXTUHybUbDRAj//HH69MQtQP3gr5V8/XFnMR/VcMLkYt
81oOiibjMNZP+8WMLjpRn8X1x+2Dpq3OlftslpSxuTOwZebwgJHdMBPhql8fIwyu
49ARpxOIrhF7XQC3kFybRQEoC0/lyh5YxRL5D1qcLlDx4V11DIU3loi1vPqC2vfq
T8cIbfewTPjMmqdI+7gV7aqRi/DaCRKILX/YglCFBto7Wzv06UhbtZBaD/ieujh4
DMrWm1Bz/4vyYJLVDKg+AJ6kJWKMcbbUV1+qoLA6BxidfixxidkAUaz21T8VWDIA
8Fo2Ku2WDWiXj7iwz9cHYJoXebuTKBbahFMtiOgBwEDWnoBKWh43VI9UO+owtkF7
yzVG+UTRuTRJnM70qYc96KkWCGo1rVa1iFQGtQIV3sFK6Jh6A8+K6fHraRsJnxyc
G/3VLRgZFeYpcwIt8Q70uQa2Gb1euikkonAOLXP0HYRHdXnWml0T6KT909jlnzOF
u4lwITD2KIOoEob9PYZYIVSZSxb5/A9eMeNJes+yS3J6l7uI7zOMdHi5B5hSVK6q
iCDkBN0n067bu341iZ4Mm/4m94qj1uAR/yqTqzXMTKGD2bkQy8xiwqG7hh9IgvNh
0JicOvPVMqJ7mW6BH8EoAKFHmzGwgytwl09iDLfOZF9aPdNXowYe/KodYcg7yV90
WyqnwRA6p4/QYtTBdZDOgHbREbjATul5ZVrZ0La7KKj+f2TpkdG7WX3fjyNrgohp
BapaTMaDWJ1x/2mOE11A6N2IUu8RkWaS9lO6WRE1VJQxdF67rNhU7DNABNsiT64Q
ePGGoJ4TGjg29p40u1Ksdk+OlHEqkc7eiAY7Ih2D8n7RsiZnfpAmTnrywDNzihoA
a3ADHqtVV/YDna0l/id+hF6owvl4Y3N2r2xTM4OcuxvZCjcVxP3WRU9V0E0FS5O4
Pe9OdHn392t8bfeayHB2MxVP6AWQCShclsk0Rya3SkkwgygSuczNEBX8qGzBq/Wp
7ccFE6p7uxUTUESDI7J2UHObJ8zgp3ell4hQd3z8i+hAEpNXvlLSZNhNpceUvWxR
287f50zNXUm7YRzX3+deV7Yh3QgZm51ldfNYyTTebQOR9QuW608WzlM4an/bhFn+
+8x6fHVbmj8jWrfc3DsIH8i0WgJ/rPaDPDFjzZgMDJ2Iza5vSvOVCvlvp9eg1R5B
NwFdNmnZO/0gPviWvw8B4IET+YgwjeMuXjwvEPuoTzG+G3SOcaa1LmMBP+r5DdEZ
wSldzHAdhyMEk8yWiiCQ4/kzbRa5WrZqaAzfvZG7cV/gWAeU0k4IGV6EPwlf8wF4
3gVtrVoTLxnScX+RhVMbfMc4lAfEAgSZ7U5XlUoXzm9lrtqGMiF26FDO+a9Ci5bg
4fryX17Grfw3NyjocNU3uvl734WptGHk2k1KiVJwNH1MVRDxUklMJTlsQOJqq3Db
FNyufcr9rLNusbKWcNNs1ry/NLe89lS4lod85UlwK6/KrXHAff9WvWSMeGeWNJIw
E0VPn4IcnDfkambWR7mNA9HZVfebhiyjCU3+o1Xilom0CQdUplaVKG5w5FMvUzr2
+xTQ16+2dGzZ/NiQxFT3H+XpIER5cQJStS9n7gkBqJ+je2uN22jYX1mPVjJx3PIO
NT+Uo3TuTP+f5tPG9P11QBPH7z3iZ/bDvcTz6j24eBtRxVMBNeHMD9VNQo5BVLFt
9driXqkbyHkdFeOUmTgwqJi7i0v7CNVsu+L46zUGzkJehBAEr9o3+LP58JKUpRn6
079Zl0BhsTnsD++yoxPJcA/tyzBnLvCi7tWYEmoA6PqUN1wOEXUzJZckQdeaAADW
u6xAefXhWAxkxy4OwwSLVcdABCSI0m9oTR0YcLL/ThctiyY7zmKHtVtcAnS8UgRE
UZU57uH+7OHAgUY54Y17SdE4rK1lz878LI2qyj7zit5iN97iZesKceRXP+uFNHxk
7OzraOmNxSDlhzE559POsWwpqIRXD4ZrGg9++3kE5SHBOnBlNOr0bIRPx/bWV2Zh
xBlKomDERIvWc6M+1L7LKJ5Y1FTJFonpwXxMGAZwMi2SzS2OiUWK+9tuO0GnxJMW
hLhkVHeqV92j66Wn0SgIgUnmwq1mzJQNPy+UfotmTJl/gyKse/f7GIp91PQNAIll
xTE9yF0bn1EbAJKz4SxfpEgkuCkZ7auYLpsdBkoFM1ssevQI00NylMuZrAFbfchL
tRoZb6V2OowKB7/c8SNAdH7VTHxUuYJ3Avp0Yr4zre/DDcD84zJdO5NN+EFPKcCU
6MnvrD1aLlwQ6oXu0OxpQBxMxCQe28D91Ryf7gZGNNBOFL1S/xJ/p+Y7NPxc6lgd
MxdEpIO1P3aUZuQoGRxFyshLRz9iPrS5tPCYUY6cCpuLqOpzNeQcx3IwCpkoVSTf
X9Q/UTF5+UQmTRNAcRns7FlIuumdOzXdzwU2obAuKKf1Owr7tJSwHoqnf2KUHTn4
UNEZUq11+Cf8ndXS33Ww919pKETMuIuDcSkCarXoGqfWUVXKv+ZDStCSbEp2vbn8
NypG0x0iozt0bhDnRaVkGJweJNXrblcNeTtXrf+tWo0djDMsWVMXGUxgpoNSBhK9
T9flIMvuH80fM4k3rAkQm1qe9S3fq7O/WuNFGfG7AOJaq6JB/PMuAK2aDbSESrw+
XkcI0xt4uk6rTHwN2ytTNjmuiu2gH7WP/pxGEni0rdJRrUPzCtyU0JwSvdLdUD4i
qy9sd6E0y6vK9L5ZMxAaFKpImFAYYhI9lUw1CgDlhDL/r2h2xKfzvOCdSak2l/BM
9izfAEGkpjX0RlrIA8BpsqrRshKHL2ovsU1DVHT9FC/uxOMLV+WU+YGa3gCQbSYz
RTd8qCftCoc8n9fBsLLv6AhYaJC1RtkHp9JK7k8ZnEqnVlvXOAs7R6YE0/+L8Lpd
qCq5n6vuisci0a3U/cfTMta/0nlNC0/o9yz4hwC/Vr7AgSsU02y81uJqHFQiMEap
DteChoCWsAWwsC2a9Z01bAvRc6rJkDryDQ6/WZSOP2bxrOfW2/XV1vSD0PdC/piP
sxa58n5admwMIsRqu1ocXlyejQzIMojjoyw7DndXiTxdRi5GIF9XK2iKQoj5oOay
peRFq7aLrdEqhcrF40LY2x5p8pkk++pFaNZZi5hgBIkugsy8F16wd62ePloqifh0
yHrqEdkRZ7N33vd4r1Oa/6ihj0gw7Nkzwp90a+kHiDDeWnet0mj53zDDbKU2rUE2
O1VCIw3+OsDgPYiwKjYZyksQ/ktYr+plGe/qJ3tbEPFiVYQ54qxntJS1h4iTVgKw
c2a63qsU3LxJOOlxwTeX8+Iska7eibMlpRENc/a6fL4Y/Emnz/ESK6HvK4goI6qj
g6TsbrRo+XFCaO9VMFa/afpfyQUIkOBnybddmZeiX4D2dFWCl2cMdsQiuwnv1XMU
thIa+hP490sd8Nr0L7W4ziiCnu2V1idrfSh3C5zUmzKoKSgDlVRNz68bxXtmVuTP
/syarmguYmPU43VMTURkNU62jfo+PLABhEWxDxfK5gscB1TODe5yKj5dVNowfVLQ
Qsr/IDGRQXQ7XiOJ47LcyKwhJmDuw8X8p5ZKG8LcDTU31VRajbkHo/SiiQ7xRjuj
xXg/HsuDTkyIigGVPiXzQlOGk+Cq3++LkD4kARgtrTKWvD+7RJUVcgnPLN2e8M5t
VCM5oHDK5tQZ9CmNADkeEg7i9aSGO+5QJiFwIA40KNletnYUlf2kB+epcb0U7j5f
l3iZyGCdm/QLgnL2z8QMD2zk+ri/s+6S9tBXdd3XH3CI4O+Wcuy4vyP70ZkI29DK
Uf67ynVa2UHO+OYZDvwrIeTirXG8D1vzJlBrPfGnooGqXRVinlY+cUA8ZRD5dXMm
TUUMV4X+o1ocdduCORNKIpx+2Vx7w9I0ACJwm37CMJxzfCAgOH4f7FsP4aAFtvE3
mUm/POKFyFdFEjsF0vqht/NEXN0abltcekSJj/2YCaYLL5rkN8roOEcTjWsg3EtP
ZsAwQP839I+/Khpy6k5wik57nVR1kdZOqBpHbXhkyiNUtMP46+zHvs1uqoxDoxCM
0g8jycAQucPcmWq6xYXvBjavXQsN22Hnsjeg2eTRCMRokPliJ23c6BSYPLLlFnx1
yaCuSKrrQLLLWpMpMvXVa5TTlBO/+OcZFHmBxsRbvYre7JLqDk6BbDramfaFHu8b
F4rO6gqVu4iM01t5FrvoyN4PMv2UD7pBaH9tdxnqMPR4JmIGTTSLdzhx9uCksZoF
+agULmzAohAXc4hZ3WoVRu6wc1jvGtkCRPuqSbJWWRb0hOoSbJN19Pw3eFoEKedO
2JTXo2q5dRoOChIzK8B3shObZRBbEZ0gdrr6noFeU6KNVcIedA4MJaCik8WKCADE
EyQjrM7hmW6qzCI5yPUAbhdMYcXktL6dq5hVARdCkwou3p4g57hYwM4c6OLTt3vR
c1BqzdaKiv1KymhrHCJljvyRDpY/wihhedXQZFmuAes7YzAswtVAU1Jqv263vbwr
WGbKBOC9mk9hid/IQemL7/ciw7gibPDMTCxa42n9lsxuersKPeneNkJgGq9j+zyL
iZRTSwyhHINxULM/I292JqjIOO++OTaV2t3uy1Oj3fmefRiVEqj1XkGURZrbkanH
ZCliqZRhOIFr32wyMo50zZyi4MBfWpjLzruU4n3uiXj3iqGCQIwp7uH817pwsjD0
6FMPCJkbwVb5okZMT47eraU8uKKmMHzRU2QCg/y+1lw6akBv8UijnRGMetn4vaka
mRvVvGDS+ewqqfHMyvYi0QHGbDE7TpcNslDamaGZ5N441ntRszHlSmnxScYoNs2j
Otif/6pxVb+md8xvrY+293bTNYz/M8FOy4OzR+Pw2Ir0if1i55j661w+VEhMDZAu
ihpUCCGepOKrohs71fQ/kG4PEfdlL91DN8nCVvoLSfInfaLkDStSjckcfnvy0syq
Pd/5O3Prwkt2JFo4xH9fFkVgFJYg+uhgBIWi0EKdg/Zv4Zq4Gv7797yiC7IHPNZf
kerN8rWlpdLMnGrKU0LP4/Dw0bfOpFkFx2nq606APOAlEZ1imEoAnmLwaoBcmQdH
x3WsNL3FrnNC8kDgH0CR4t/8ePUxPCsMwiGh20Lucd141KY+7igogeLm7GXDGPKz
9v/osCh4xq51+kpmDAF9QJXPGNDZGRBmEmeo6rLGxOgSV+8I8aPPOAMDV9zLX9IZ
LAcegwM0tGYtGLXW1DMVKNuLXWlx3QDFma0oR3hZytQwvkimTFzwVf0F0o8XHcvC
Z0gDaqtZBLsHGYEe/Nr1UlCTwaXkfW31TzKEZAAp3fu3RABCaNO36vatz/Eb8Rye
eWCjKIO49d1PgdLBxE/3mpo2y5+6y3AxVNWDl5dsP6nZMU9O2aViIkwu4EY2jvGQ
iZqwEyw+Oz26n8lwOQOEeq/LpWG7SGc37ktqswaEbqetWOkqrGcu8/BgilnK3DHt
HXHrRoJwfIVSc7gbkHCk+gSj/ghQM+pXi5mqZHKyaNF/HgugCvf4RDBhuiJuT5NS
pHdL+AJ58BbvL5MH61Z9N2/1aWPKF164sxt3n9g0mrKB23sE/DRBYnNAJTlCGkW5
VkxIOG6i+lMtVKBLzbgJPisDfNRoHv0Sp+q3zIW9Z+LnqjGqE0pGgG1tKPMis2yn
tTegnhxqc2E0/kA80T6Z7Pco0COb8hwUWckckTQCwd5Unv0Yg8PKY0fayu6ppiXe
6Nl+/IGIxDL8RbeJ8LTgYa+KrOGD2s0pc+4MA08/N3sLRvQN3oDMLZnqtXFlKet9
CBzNm0aAPDPpvA+Gy/UbIyUHS2uZpgsHfY+NwqH9kRke6qEow5R2RmuxzbPIDgTQ
CfvCnTPWHGVkmrvIL09iAWMJ/arVqilHqrrt8O+E+Z5/v3ANq9kT3JmhJdKGmWrt
oBqnviRD4LrSLfD23nRWpfG+HtAoEv9VArkt6iCctBptzRYnSjQ++2psB1/pNIut
dKISlH28m2FDI+AN3Cw7f6kN9nLjbPepGR7mLX0+MFiPScxw+xjAc08Qi7Je/Cv9
s5cmIoko62X272uAVCvu+KKX8g3l7WyPGLtHFyC/o1Kw0muw70hnPbmki/blsqaK
BzEQdCTmr4WF0GJmsOF1+U8S1icpgdXeTuFfP/Jpeeq0jL7OmUDDQjZiiPxNXVCI
8xHHsL5xR/qmC6Rsf1O3Uq4Df+U7IJZmRrkQf9fWdO+Ze3dOgPF/dyPxmQc4l0ax
NPOGkQNokb6pqQiB22gjBAxMejrCBmT2Hu4I5/AGD+f2icCDC8bRRLjXaEYbsGCq
ynmcKRLz/0aMsQ6ccIr9qMygpdvd/NzWA5N+yRgr3OX5XakA2EtPgDOKmggifFMU
56oGC0QiPMpFu/AwyjvKl0sAedqkjSnQJXAiN5e6ot99pyVOZ+MQCeoVqPoJDQC9
Cd2qgBK7elVAXrJeS1mQ88ZpgGEnsB0/4HRnLnyHnY0XaFVYLYQaEbJXzOO8+XSe
OMgX51tYv35BVsvQlfHJiWpzTtofH99Tm8CQQVKXCjRi6ef5kL9aWGsuuLkrwpOq
7Ah3TAtzI0+SXyinPTks1tEjHFJPwlc5mYn0EZBzCu6a2HstBWTXtlvQu0uTNGOM
fwpbj+k6jWi9trSxDgPKzR8ntwcLfKRosT1hSGh/NVX8oSpdWqO2ftW+JPnQB73u
Ifar5/NbDBwK+uw/DJ6OdiJsBIx+OtRYeuHjqg+89KOAyrqrZJ1u2t8QWh3UwYA3
kkznpOklA7SeALW+3IyK539+0MFVXsQATklH8OfF3/dIZtSbivw2KpkChrjOt2V1
MfQOmvsXYKEYwA6uCLok23qdKqEszgwPz+w5u3OpBjSo1/ejLKwK9MhqH1vGLD7Y
Tj1fc8Y4BHmsxMv67MtbsBP6BeWQZo1ibMhtQDOmt+CDo11H2M1nQXuaq2sKsL0K
cqlgGGA0vb1RGh8TxQmZM+BDtzZxZMg6uCmcrZO3/FfCreGoMB3e1hCpDCDVC8WZ
vhw3RXhhWQONBY+XbTkyMb9W00jJYTtc14lVf0ddHDhQf2SgpkJGUOTS83QnWw/i
VrldFaHQS6Fcn//SJaSOZAw8txlUqzUWfchBFh7/Uaf9LW5850kC7rWo5dsty5bh
/G9504gZvCAMikTmoxhCkQi+LMn9WxTXnvWPggHwPEit3yHToqBX+YUBuO+ya9Tw
xXN0EcGmIDKlRxG5my1lnuMoLl81KyCDQkB7KY6SeyJxTgREf4SV2X5B3kVXntfP
SjVL46o3juA0itfW4g+euEdlZz+zVbmxgv0jNW78GRl4d++aZJS9NjQpMZgSxx4r
sALilQtX5pbu4VKqCJCHRM2bDTQAIpfOdu4YyI7TG2TDnBVOwIe0TahUZ0e6SvKs
oKt+vCC/KAYf88c5srcbfIt3vzyP6+e0JoKU6mPzrUw+6SdX51kkgHPOoMoP1O9t
FhOltODCC9B74G73rlwN6scYeCDpOzlnOSkyXoTvhM0inHyWM2voijIfyHtMvuN5
RuMJVGtuIZeQO4WN1c7JTpeUJOc/xNJwe3Jf+I2dJbHJp4uQ48wZqgSx2aidtPSc
7wSe3uO3yQnrpR/CU0yCbJLHx7HrTC1sT8sDUFOcbhMc2Jy2MwykvTmxDaKnB02W
K+7k7h/tLHaA9JOhAmhnncq98d2K5hjZtokqPJwWou3kFhcYFJWNcFC9Btb50F6Y
r2bCYqTT/5P3nbfbJLdIt0lrITL0wwgtc0SPNC0b9eBJmwNV7XHxkfakIVkkBrAC
PzC1/hKdNSe8b0LdJDeOsldP+4Zcdhqcx/bAZ7XHayvhRRC6Bs92dTAxF+kE4KHc
gLukKKCw3WuIKth4/Jnfk1vZY+rTZORcKtQ9P5Yy83Agi1cIqj0kGTHVKg6wGtez
CH4zeoti4zkIna8Neuq/QHyf6Ie07enr8p1DAVa0gBY8KK2a6kW/HJo0/B7aYE3c
oL4GsrGX0rmEjNuQ5U3ifsaCiFS36qcSQBeSPEPHpg+msDWhH5utgQCXLSxGvRR0
nzldCZ1BAcL8I89TGO5XZSqH6zsqvEUbumzNQoIbJggPeeyZyYJz/Kd9QZjcfbch
CvmkCqV4fStqaJ1FCUqA9KojZaLhZ6osrZnD8LTrJW21n8TtvF7Hc2NQwxPC6SAQ
SxUjDQBKFizcdMl+h+x+sTrsavzeJ/8jKiPf8lQ+qtS3LdJ8V9JyAZjxsLQSUTrt
UO0VHxn1splSjhRuQt2cu7bic6X/+krUK4EE5e1rFsIwXmvgAVGHEgVTcJJCzvfL
efNwhdCklWKDfEHk7vVjl+Tv6OcD4USTL4HLqvqNm73OO8fRaRKjYjUgD8LD9h2V
rsHL39/h9uS9FcqwY9JAO1m+FvcRdXe4nGu28J3Zhyb5TjAi0HpzDsc5F1cBYCgs
MdMp6FMOtj5knM5WMNbheyd5iwE1e0w41DhzZrh996Ofdx3X1XTcAQ0NZNuCf1iT
ghvcWmUbdUJ0KIHdPIHvNnXSbSFYfDvlvqulBpENnLqiG/4lWxfxHIFcZyYowAAQ
FO378wKIOB+8XMoTXahIwJeVnObB2xb3e2KPeKmKPONTk6IOO4UqpmpJqqJ294gG
99Kuu+juLheTms5Id6Ixhj3kBxnF4VWMdli0MY0Chgr+AhbEqsSmjMujF0P4C3GP
PgkoaPraVTOo8fyhLJ8e6aKPNzlXCiAAa+GkOyFZUExQtj1uDCg85rnEY1/2cW0g
rjm4C3S3wL5OfQBcImJeibotLpDQ1K4vkxaedAl7sGJlp/ICAJUR7M49s/RoUjgY
dyxGEdRDGk+uzuYCZe4rVS8PLT1cOq/vAUwprKwUX8x1NUtVZ0WDlEfXL57ByQ4s
+iICIRduGoOmZDR4gcJJmITaB19fvL5/7h3E9cbjGIWjUeuk78soZutCs4nUbqBs
0LXE+TmT+4dfWFeip7cB++xxSbmA0Rb5ZhiUp8gTG7940UjZVRA6KQg+J///XMkR
QtxZhH0JiHyx66xnZpPh26SbovHrKrBkafJxBBF86jUvIyURYoTv9AgBPvfedcoQ
20nSthRiJvc5yWgHYOFMBBm6sNRKk0q7rOOtIKlFWL84QD93nbTuOma8cMbnpnR8
kKMK+NYBV6mc/l+5TC8ivdtxymXYD3McN7hfiQakVlYcM8n6IpdRC6ftNlMnu1ei
MtWjY3Jys/OgQGPL6gu9rfatppoEpv+fYAXTx+KORT4DzVXAQhWKJzAEgKzbs4aB
+Q2manxaOk/4dJudkYVwoooambCWEToeBZr2lJL+SjKfTvlQXIzzBFWjkaWZgb5g
rUANEnpM0VuAWGldr5g3URM8Gi25KaxVl1gjPkozPB5/aNggslFcgW0XPvnzhSug
OE6w8MHu9kiV4uS2zsBgZV0UcUObQM9+SYtvlyr1H59JtqAHmBJK5GX11nWmf/0f
XVqCBftV/GOUkWVOVrTLWQRB8W4kaU7/LAvfnyPiNiEsTPYOtI52wqQyzAHW9wRG
HFOFXU8Ir4c/j7GfDQ9/H/BViHD5+/eEfNG45/IgyIuusSIerC8nuPXdML8TOK74
OLcHSN0EPJa1EEiMn0jyngK8MSNZQGzic6lRmPHrakh8CkegtAK3t1zTvoYthBVm
TT4gtfwIfnoNPKz6ETbRYTUtGZkKhSvw+t40oWyxO4HFxL8lsHae5mwvHYWvOggR
O+mm+G53NnUWDu8/dkcUa0VxCubcD27YVVTnHpx/1L13mYzOn2cs3lM3ejK6ndpQ
0N5c9kE7wLVLoPBxLvPyUz7Asneaj1mFL5hdD8bhUaq3Y33wv7D67nszSx+fpzpt
U3AS22odZGMkJcrgM28NZ+CE0/hrevrdxO088hcXMt4LeA99ZGqxABz27Qo4nI6E
bhJ0oOeGM6E2UT6H9UJZ3xiZS6ucxhBrIr2bVoymwpKU1v6FG6Vyzrah6AFawtsa
9tU6lmNtu6SU2Nd/a4HuyATNv29yM+0inBJVeVcHCPq6qDWp4Kybw+jDF1B0faer
0SiBj0UJSD7VVyrpIPpDHaymuP9PiWuGXQiUdb3hN1+ZMw4hoWzs+AGKcvT4EelH
de1ngLtt/BIjxCu33pqoXXFmW/7JNQDknfWChLjsWq/vnAFgA/7i0jIJBUw8Uz7V
Ws8WM0OYfA0GaEGLmQpmldRfzC5iynzmoYRQ9MtkPaOGqcfXYgChHGdCjsO9BpbJ
qek0DjwskmjHA7DKdzHEeCjowjXiU9eQ5UkCDjA87sBCpFz5709k7EWFcqyaJ7i3
KgoMklbSRMit4Zu6AULjDQzR6ZHOv3y2jhC2XTZ9o6jQolFRrGBg32yFe2MHe+wQ
vpqKBHKRGzWVQINYDT1/lrMW1zsTBBnA1+RQLEcPF25OKWr43dIwaQanz83HYKSS
FDXbR/AdWbJFi0o6E8zf1rFe97bKZhOpCkgYDAuFjqVPEC1OmNv8mPMScHRdOPzN
f7hwwgnGcK64CB2vTeyYlXY3+Tq92jQ6gyV0jr83bOmtGsc6SgmWAtxXIDf3e3KJ
RO0sbgrq0jIclJpdPAtQfGhSUMbWINfUPzMc+2hcsEuazExt05Dh9+eilcyBecRP
O5qFVADH2dVJVAMapFJIcFouORdxGccPs6e8kE/fYe4WSB5yyiGy6FdWAsYxEouc
5g/lbzSbNTCujgnlRypJ4QQqtM/1lXsT1JRnqg/u7aWMXvAQGfPkCwzAsxgPBfY/
O0x/Dnai+7+5S8K6Xc5lj6av1CW2RuCeD3A7/sMToZUVAC0Fie8YFHNbDNH+a5hm
GAyMrObDufq49kKA7v/jHfB9rK0/i2xUBoX4q6WZs0F77VkeAry1u/bAbKF93+3M
E/VVn6NLbltuKZ2pD30F9HWbKCc3SefixINYQyYDouigSfsRJKyTcF7DmhpuHnkX
Tc791az1/yccvN/0wH2PzMOtwwBAn33oBGSrgXTYzqGxwu3NlT6Hgyo3cgYwOQx1
mNMRuY4BdjKv8TcwUsjioIkxJIi0MdTtC63Y3M9t9u41fhKe/611zfkJJt1EGzms
BwoQlGdxYTtdCW9Jif2HypwHVTMYfJWpozrkgrL+sN7zqX+1gCGcSRP2PaJ5ypfi
88W84bwcsZAuGwrsxzmlONdHIiF0BEq+8Ne7N5/h9rBiaNOIXgEKARgD1UvMSGgT
xtVv9uBLHrZ64mFBg3V91S+2GdYhR+QTdIJF+snmU63mG6b6cRxuu19fXy9+Mikr
D/AxRPvBxbez9A5HgrY6zvTR9Lc1IPfil8cUiMRffsX0Np8mpKz0PzpIoeQcXgrm
ocuFXccc0uDdRMW/PdkeXsec9fo/UFwFQ2FDUESllaILTDPNpv0bJJSVUayH7NnH
/Q+/Gp/zrW1qjTImEgjNP4xpEHav5z0rrHL0w9pibSu2SbwbtLwuvUw2r1n2mtgF
SGAyrGl+IxRA17kfarSmYXV7kemkJ4vMApoBqzmVnWzeF2zPSEkea5BnnZMN/z6N
mORyi6kZ+RdWbd6HrO9ltrbLl8BKHGgWt4B4V0gj7QtkwAOKjv5TXvGsTnqytSo6
KqVDPy/SZAakrB28gNKDsGrwTPRn7FsFXgx1d2QuhHZxpiR5upSzJ4Nid9ZCuimH
kfc9E8zUGI8+/fyevU6hgao5E6sg1SsMNXVFPtEubvnsJQzH4taEwgi3B8GMY6aH
WoqU6Wb/Job9VJLSLfvjDAzXancBBxOSz2jzMS5ei74h0aREJgD9VpwNE3LB4qoB
2yznOTZ7jrzLAJXx5EMRS5pp03wnU0SjaHU2JJgg6HyERUf/mbUzronqD26xM3jc
4UKOKTEv02iB02MJ3oVPpEoidFS3mDL/LWBx0tKs5drR+Bai7qqpA22+/eQyJkPH
0nuUdMwjtSoYerQgVzDBmbA5nL+d2V9EoN02AjYoBUiRC7sE4U+AT9IvNqcn+YNp
31FnPpsQrj2ruT1c3Q8uQTq9KCpHPq3krpifMDx+j7OkN9mlwOpIJ8dEcY8xAzHP
S3xxG+Kj6UIEoyXQWsHtKYaznw14LROtl+6gZxYDgu0ybXZKUrNvSbK+ZGbVfKi3
TD3O6vULEYbmnfjfrfE73ZXBgktsx8P0ZkjeW2T9c0gnRfcPwyFlewe4rHRT7R/u
jms4h8z/2sEwfTEnsLOi45QANybM4MobE+1R2w9K0G2MBM6ochHMsGlNZdkUmye/
K61os7dv3Z32YUnuLMmCOGKxjewimg9voiP6OWmLoBVSxkP68gIjKNiouqitBCmN
SWW/lx3RKGlEOTKM/bfXtjB4Z/hdFF71et7LPmtkFZM0vwIDLLvQMNbY45qvlaaP
31lts6lOMAa+Jy7WofUbVloF671y55a4VkGcDJ2z+2g7hOTbDXfwRdHeg7UNlb9T
6SlPayW5fDF0vQcAo6U5IgV2qTot5vbjkPdYHMG3dzpaopoq1oqhbTM5mREtJBuD
OMyLjKKxGQXFaL1iTGG2L7Vnh22zZqv5QKGRwysK3dnctAdFJkGwKK799pzTom9K
n2rB2xoNUPPJPFQ7JBxHRVj3brzegm8PUPEuYujfuWCX+jplpRwTKMFE5rLQN4Gy
hmHO85K+GeVM4UlfEotGr5lGUK5MVgoL4koqbZHW0fh/5XUWPaUxU7MkTLl0haC1
0/j86hnrIZVBwH7P/D6uUDC2GcH8bdFICkbCinRztCij7ybV/DY5CBWdOxaEcHy+
cFTJ3jegGbF38wnfYq1fKPm0WMLC5lcopaDY8A+3YK7QbLeNzLtVtSCc+txS+7ua
vwW8Sf+/77I9s2q4txYJntmvb/o1EmSanQ5MiBVWPPN3sJA2E+kiwbBa+tfd7+5e
MTderd8aNRMCy61/t2/6b4ypHGyht5RttUb3fg8sRbq75gsH70/9EoQV7pn8ZvCt
1bk2xY7EyQvPRsTI75QmxA/d7FuvG769cIwRAfshZOcGLvZNRQUHiEOdHdAjjNBj
40qmNQ8uShpEEmvfiv8wQtT4VAULzeoFEW7fEmy3guJiDFJ1UZC1KPrLhJslZhRF
AAXW3nMhXqQgix1a5GqyOGwl7tqY3fWkAl2yCT5YeKduNo29vrC4ePdbdB5j5JW1
UzMUsQe6a0JonIW6drL7yg4FyUP7yx+10bD58vZ/IxbiNWZh7ccqSSyGug/zh2BI
yaP3V3dp/pbqSzFRSzGok8kt+jjds2MmZ90CuEe5WNJPgKKdyLB//uJ+iBEOdVxh
QzKWvuqst9JbksMMD+cP4vpG/hMtJnIvUrhCiT0trIeRLZ/3WWSsvpDw7HfkdJHg
URdfBdrzI8+HP3C4C3W1oaHGJvdXetSQaY9yqrWLXOVL6yW1bmsY11MPoCMtcx3E
w7VM8kCQZ1XjlpoDCvsBu3w12qnh77CpTOue7MKY7/2wyh422ueptcUGYd5es0K7
U7rF68LUQinFkDJz5aUrnvVpIS0pYFCZm71NZNM1n4mWKByKPwex4AfQVoym6bQu
7a0VCwqkwSfoUSyuK/hmnsElunUlP1L7gXacvqd4UQurJMLIOhyDrRWqUFxQMNBb
XH1oasrLLpIiwEmyurREovBAzvgPNICdHcMyQgVzLmY14dZ4ni6lkwKco/CcxeZQ
5IJwBLhKTKok29Skv/UK8jUHdJd4nddOK3FY3Bu0HHegR5MalyHzP27jaXOq4PaM
Qf0mdRzi7m3lamr90D+SVaOWAuDoo700miH9n1RekdEZjnSzVdRa72ns1Tb9sOJ3
/8mDBPFZoDlelL9tqmZ82T2OizHEjw1S7wtbD+yLFbEONC4ON8Qm4s6avvx2skNb
Eiq4W9a47Gh6n14HAVzq0VxsXLaPqGLbiuVJYpoRlzvG6HTNbeGITJwo+RwIO+vu
cQLJUqkPQB6tqOCPFAzoxCy1fTk/pSPZyPd+7mi8xu92sSpRyJfbRehJsOoWB9cC
YLZv6eEWEy65ys5pZaSE0bNo/09d30akW+iK+llbBa0eA/aE7IXDH8tNLcrIVnya
VY/h0JER+N8YSbGAG1ouVmuvNWUx68/jprkDykD1RTl47SCE+B7odCnyXR8R1qLR
20oG9r3aknhTcfxFa7m/jWbm+IMzPn+h3BSZjb04vtrxbvJLl3OUFcYnpkmD21lY
/uDFC9CN7Yae8U7kfUxtynWbnxdM3J/O3LTJehbSoSkvklJx63HfN2gV2TSajT0q
PFUC+MJ9v5XKYe58TIU5921hq1tStw0EduZ7lmrl7RghJy+fym/0JoYIG0iQXd5f
vKcI11Abc9b+plQEqSo/RhQN9TPqws6e0TSxmiE1x9g7yJpC/ar0R3MEqcbydVvC
m0i0Pcjo7X0A6CNBMnL1ctNsUQ54UVUJoD4XP5EaZ3xJrKUAXsyPiHxN5oDH+eE4
WLv2zSyjehoqdeDuf/p2t3KK6YD+uRfMJK2gu4pgrzodR4oBuTbiw8C1kl4WBqOe
Dt0JNM7FmLvby5NqYOdWawYtr0yBhOSpPDxIlKC+H9YknkVC4k6XkXdlGjHojz/x
ZNjwgLDV+obxaUfj1O+E49VLFz45bAd5H8mWJzOgXRL4PocwIHKKSVztSu0HVibN
ZdlcSgV+vw62LShhyI2FjnCGVi+OPZ1hGhBZNX+3CaKGgDj8DzpaD5x7dHV1dzRD
4WzUlAnXx7q/Fw+X/4M3LWjpyo5npmq2sQN6pz8LyPzNWTqhoCgjGyCyzoytlikP
4Aj0LVzEaIptwBTpgAsvSbASadqr5rPVwKDkfxcfHULiH0QmxKoXBGVJf8Iv//56
jxO4d/JFZwmVgEBt+aRM9jS8KRDOt2JsVQpitgFMpG4vCh8cKLa3rWNxEvw3+71Y
8G6zgZLogFgH2p+UelNYrqelY8KG3gLzCqCsk8wZQAvSBqRRdD4l4ajlE225B5LQ
IdYvAok6vEh6OK1om7ioKKTdTPjHNRVdZZIOBtlKXtslz3Pm1GB6bL4ARA+qqUSy
fo9CNQpmFzEDgtvrR7KbclgmkHsxzzf6j27p1EN0ubzbDrzl86jq/1OpSGDU4bdd
eSu2Nn3QE0rolul1aWb+JcoJdLEU+MsJcCmIaGlJKPpkR3tA4hBYXlevxlnBVXg5
djqipdHoQg7VKYKDWCPf6OylWgY8rt32zUUUdDMKVzWWLdRl1pQh15uAUJJRY5ec
6rWfj0EXlHpnYygfcC+9CQbKDR/JVeg0TOM0XxO6uwXzqMioo4/4LEjW1fxtnwGu
+9JCL4pPSnyxKTkohQy1oOeaq3mTFq2MKKNC1dCP6i6Tt0sxTDxN2y3wegS0gccD
7cyusS2LIbyhHRXLwC7juXT9/wkufUbLTkjZGtdJo0kwIWOcAfsFXc/IiV9cnYv5
ZboMdpJ1wWBB+Hwswn05FHWqBnXm/lFiUC1vLz+bT9d6TML2VojKS4B27AtWraoV
PUF9sjwGbIEMFOzdDt4VoUsMfxFecJSaTfkZ9gHt5wATsR1ytizm3s90rwKboJUs
F1EtQwnOApQVmlxzu+Dbpc+I8DMu2vDd0ZhpGj0YLZ9NLcPLVqjt0qConpLkJSYG
A7dIVUKUqPcC771GfOr6dmgtXnsNNcRzkMQiJzjoZCLkHrf0TK9JPahWVESCvvfN
rPZ889SC44lmEyqtYqD7Y1WpyfbM2TASL2hgpsitX8WKAcrEvLGuu50jnnli/atf
O8nXD8hXQqI8D2a1hN7ydQd9h19ON9aznWtv3SrrC3V0ZCgk79lG+ajrm19vJA8p
QwqggbYVzCyFt1fK9ma7NsNbnYBdCgitih1JpFShICg1kVztfulpJssnQKwXGRYr
wVoYiJsJmlxXzEdTe5v/BGI5R4bETK7CkKSzWjWC4qgMVM8TXRMYyqMMJk5Igl04
e08z38BUD31uGruMQlR7nSwATsxf11Wf0NUdTOfFGTCE0uUdWLd7B0GVTMW9fz0/
ngBw8BzB3kuCDWvk2feghVkLNmYxr26ZoyOMKQoauv3R+b0n3T4aCX228jyChJ2z
5aS3QF2bGB6Fg0vymnntTnJyvm3dMCxTlhBwMVupHV6jtbQBGnH+vU2t0cbcJ9oy
0g/jY5HikPJU3sNlLcGiSXLjUfwcbkSw2gS9JCXF25x6vhFmhRpop/uVE5ZvPEdb
CH8Q1/SMpSoIS0xQ5Q86ki3c9sIwclar5P46vQRef2nxn6e6G83M2kzY4EiRkcMN
5no8XV8w7z5GbACjr7kgVyBXmy+Awovnr9jqwFutG9T5UWXgH0UyUw5KUCeyyVSU
si+P3NZRlPP2bKiSBFTdLgjgEbRZBamy6GhOiXV9sQARH1jZs8SlpEptJLK3OLTf
w6rNl6P6su1M7KlMQ8gPyEbNCm5RvuiKXG4JDnLxAsBPX/528wpC7MP211uM0rB0
hSs6Z6MwiMdcJd8hL+0mwr88iH0AMpgqboZ4GqO0nm3Uf6TBtZvG42OC6hxoh0y3
xIW/nHtGrq4NX+6UrXal6+blJfNMA3ULGhPE2dPpYZhB6hpUDRVFVPsEsM7cnwwz
wHJJM6Z7cTKWBUd1/Yhc6MOSf5FmERZIoILwFwVCrr0UJLVGsHM3TacwbqSyMu6C
5j5N4e5fXaKJXG3dj3Tyl9eQ+BjRJxLZv9pvmiDdku9cF7vk41hqjfarDLfDfo1P
EWuk7JpJkqLkfGhh7OGPggRdKS/Dl/YbXtvkmrMpK5yjAnP12iBIVjOQyh6NMGbL
lZHGQGig1mUkHSqxrDjzNPktGn2TFnD9aFsofCUMN3AJMJYs3/joTMW5j1bKLkj1
Eqed9Lev+uBQTSa38QWghAKpewXaRg051xCtrRkYprlKWyAmWytnzQM1bX6D7cdk
TayblsT5OavwycHzfgcbKY1YFzdDa+Zv5wYo1rMs9ivkWgSlCNRFkztLu6vpMFsg
PsNSdoMnLheuvWlw+9MYxRF5K8fHo2sxA77IYyt9WKjwRWcOEB3v+p8ZwSG1WWBC
bwXQycD/6ikEDjtbEhPk7DRQX3suj2k9ijj7TYEK+TLo0YJH+yCpTfyRQQEWPq2S
j+xDXo7xQGrIchcV7sodZ58PPTzgIR+MI+KX2BFCEt8yGOtH15fibC6VtJbfLEyV
t7r2URlMnRAY6RzuNZeQsBoY5eYd7Ox3k9dEf6IHBxkSLrmDHHtqJkkCkb4CDCpR
eoPxs7UYAexmtCQWiZnDA6vnzX958WvbQrvWYJxoO9VIbIhqXnW++ZO+bQeym155
rm98qfIdHIL1TiJGMyKg02dmennCGBsrvZuD41TK6J0aGKqg+xN/khvKe8rMZfk4
coZlKmsaaLW+zzfA8MD7xBuI+PF644NydsBlnstwcY5julwWIIGirajMeXerUQjn
vw9O/BptCf/QQb4w4nU8Ue2tg0R5oe0/0M0Srpdp0bATR25crsqd2m5GrAT5IsS+
XYM/7sr3KgLbf1EXdCNJP9f6FthkbWhm/4cPwDpq23W9NaowOgWGnk3raI9mLQ0j
ql49t1moQywPFIfmeX+l0pFcrCCNnW/H/wjJOSkwLwlypeTZcff8JMWdM2YnvKtq
eiFlOFWgMgB37dgGyQBnvEFQSOLeG06mG9uCdYo3dpQUbusCE5SeVaVp4JOjaADm
87awZaFd2ObV3pR3l/WpXKShw/vc5+mmUNLdBx73QPKZhe3tb7ErtQ7Qb+pA00Th
4o7j6BfDuuMJEsj9hf4wlCkp2lSM33Ysh/HFZmUOSm9deAvk+64zoSqKIRQh9zZp
dwysItqIIHvYgNal1kXq/ApwvnxMggxAS36CAo5CzfxjlFq3ebu6964mLD1qN6jC
aDe+fCMVxOgfhHoZDhSgdHMfKBedcnIPTtuw4MXQ+6lWCJp4zlf5nqRVpNsCd13a
Bh/b4OT9bTnpmQtQWfYsT1ZH1aIjG0lvXecXc7yKRvnY6rE+z6oeCEafUzMPPAkH
Zwt5Z8Vvb6WXb+YMoXD5PD63joABXyOdW2lr3A4lzEOyhT3LqeEBdDlUbyZEWTsu
ZrQLie2cUIVoJEAMVOvXkmI3Fu9ibB6/eduYz+HtPf8hQCi6lJeH4P4ijgWtYFeV
oQNLZ/puMiFgacMCKitd0FF8Y0CmMvOnWQXVKOTwtK1rPemFCjwUHY4r0iQ9X7h6
2DpVhuKji0nnwtJTOzm7fYnsyfrLq7Rf+thaUj/3jjtKiKn0q5EokV3opgxuip0p
/UDIQNV70UKAhUgxKm7Iz6CN63Pb7yxVlVl3jq8ynrVNDWtqrwkiAkF8Hbb9s/GL
893thPiyUzK2OPi6KXrzc1f+LTtLhkwsqynMr5ZKndKfSetaVtiM5gX+Xh0x6bnF
obGH/5cQrhNOLmkmfwJ/PkILsUmONWDYELCd+Ap/5qMyXlTmmIQzXUx2QPTgn6+k
8u+Wucrs5fHAm+wkCqhrxiMV7osfDYTgKA4U+qoF8f8Sx5bxf30w14XBy/45dCzQ
52iCcnl7HjzyMJT2aO5kgBxvIIcP406npBcKnu+9jQsdfE5nWkA6UX5f1uAo4KrX
rYHEmCN07PaxlHBCKQUCtQQXTTd8gPMnMT+JWFKbii/xoGgOrvEDAU2RayiwfQHC
A55yLGoVDisj7+xkEviI5wuSN47OcmIxxAO8r6NOmlnslOU75szWhqVWvKBeUKY6
udm/lnvuwnlHQWjKZkHIRfridL75svDR7TP4lvM6zsmUnsDJwSnGxBmo5AfSmCb+
5yvm8ITIaJfbFQ2kmyLBsjFIHUcudlsSYbX1S8/WDNiKKcnjTd4IoLpMjGtu07Lx
13KibDFpcDsFm5YumZswG2Ib7MRMiHVuEV0heMol8vFVR2XnzAS15mOdkvf9aAD8
zH4ve4HX3EnUs8FsvEb7QuVReHxl2g3sghvTwFSW3UF/CcxC2mdit1+zAJC0ZcWv
LrR2UmRm6f/UAksT/I48Qq1ea5ikSFHPJNX0TfoKIdfV4Sly0ml4blf5JGWRaAiB
DNSDWYp1Q9BXx6NbI6tkeh0AxhOT4tyhsESVc8aZVrPuwtSZYACkgbCNAL20hmEg
qIQY0dOuo/F9xTlm1j1ps59cqdPb+Rpk0gdiqYlzOJ48nYkrwOryhEvJWrgrut+P
mnfgSh+5RqVNb0bt3fk9ZVdEH+O6z27m3wpUZkQ3PgtSnDyzB8xczESsLLsP9tWn
6LhRI1/YIw9tD1lDj69CpySw5iGVQsXJ0sTjJbkmbiSvP03FaRSNMtjUkC7Di0Wp
pRKHn8fs1BN+rNDJjkRIm9tC3OyLhnydLk5L79eLJTh5tX6SactTDtcKngvV2GbB
B7Nyt3TURs7/xJCe3fYjYj/sm72HIyzWE0oEkBgBKGRfod+1l5WedXzsAW1oZxiP
2nDAlM2JIQPtQdS77OOYIo187NbzRVehxOLM9nzjCJjsACgQOPhabP4DvDdCZ15Q
ZdMGQUl0S159arwpK/wXfeRay6LA/VJb9grs685J0AejwXgPqGnyA67yfVcwFyA5
fHoyEvtQGAX4OccnbsS43Ajk5aoQebEfIB1twhYG1rdA/sLYzX/ZH+5S15AHn18Z
aLtCT2kqwysocD8lxtNervltx6qyoOZ61PVE3N2HYc6duLI81F/+mhNP7WU/7yfL
ed1c4xwK8kabzdDJl2sARdDNrAuAMhPGTjXVSZf3k6kXVf1nMWYSwGje106zgn/o
DRI6J273r0Zwl9gq8oel/y7dU+EJfzKz7UnVLCOqefcRPLg42f2ybo+EHaMPRKyy
RlBGZfwWMCdq5LrXnt8l/flNPF99lYM/Xn3hpeenqMEh8xAJDGhUAku+JtF/DTMo
hNEp3RLUFKAfj9VQc6g6F7CUJiVM2FfGWObPyZui6qz0LtTJ86w0DKvjes3b3Gxa
PACv9Z9swqPpvRQ4Hb6u4UXlEzj4AQ9OiVoyYKEHcGm61GkuZyT19u4aEJqdJrll
La67uJHDS8uwPnh+9kJ+TMSN/91DpjE7ecazcrAhWc0klDacuuQRhf7bvNcqe6Ie
6Jk5iIKi1GWJQtzZ42NttQaptFUiK+wbdDawkIfU5KWRBC88wI6Z3SjS0nICLdib
1Emc4DmQi67vojfNEu+R1+nfM9Xm5bdY+HNFJcAt3s6lsg5mYalWmwD6TIXXwh56
6Fhbr2KD1BvjvznYUUnu5OQDt63LgZS6XG7GEnfm4x1jlgCU60IJayFUWI6Xli5F
qp5kvF9g8qICyGSZEkV4cxty9AOITGZRXTWN5VF4OUNYZS8FT8jyYHIGCTzVJLM3
LVy9lriG6gge8sImGl8iLckCSh4/GZ6navBVisk52zx9FyTOCjvpU/T6xgtECNTv
Y/LPHQuoboJeikRjAsGtKY3qaxmWV6iJP2PR3OKIQANzB+htI6jKq6J8HrnwkEZW
hqMzzclGUgNiVn0e2+BKrlIPEESI4smXkrPuov4xDeOE4OzJu8e6sV4nI43RTDWG
o8bA1mDJNKDEWRTBydAksgXpDEXsrYYyKEkUuaD8MXrrGCG4wEjuaof14CROmv/G
ieibsYjIKGx5Pb7/B9R4dhzV79A8RbQGz7nFNBUjSk0VzzWn6wJhRYVNJ51GwScy
l5ttrotyRr8zxF9J5HY2CM7rLSYOfxqzc6l20OLYvTUc3/Jjdi0wPxK0cl2ZjdCG
s4SEoTFMITIhqALMWX6qZvkUmILguUVtW9GUPwMo8JwR0RixpQAi6ZZEvSWzANwP
dv2pptjVIsfUlxIzgDhwAh7Yb0iIj59RHL3Nxd+kH9PN+OEBPA8JmoRTburJwEOm
GCyYPFkX3r5Z5w22lDjsr8aCvwsUQn/pvQoayBOB81V5Xwh1JSffap0n9g+GDxYq
BFYirYaK3eZO5+cEwzXvRIyrMdJWT9ik5aYSAiUSDDJXtrc667g/3ggu5fDwWQP1
qmBAkLMUJxiVAzTAUXKyxhuYCLCBvGkv8+i7G3S5W2AgcS6+EthnZ86SzQM1pS9t
nUM6lU0dQjd91KtTCon0RXTj6bWzDucXxWHX1wdldE9ayRr9p/M9puSsDwwGOqFJ
ri+eyKVY9JzuiD6aqgaX1M/xtrdBsMqPhqb6Cj1FGCi+gErQQgHtjPcMz2CWMWuS
dRHC1gsa7TbdEmVjVU02Lz4JzLh+yWO/6Waef8uBBoH1M9GJzs6dGP6l3KE25mZb
lBkMIh2rQD+0SW/G+aEv9vXOXrn7N37D8wNPMAp1C9sifZyf5XqPKCIG5iu+JzdV
rskQF8xTuFyrc/gsU8E0VLRpw0vLVLfRyOHU0RlH9XsuVdpFojPJvSxfVo5UqwQ4
PoKj/R6P0Ok7lgDU5BMpoOZqarmlrMtSdxdqZ4Hwbx5mxEpBHQSQlgBgNk79hoCE
BXsHCmpzwM7bdae60Fpy3Qvl77RuTgZFMAID1zXJkWVKkwMY6NhmxxyC7qfqZSfX
8ZZjg1KrJwvSYiwgA4NjsKJebt3klDT0o8NoWK6v//mqguHa+4exTAcck/lpFJCu
lIzySSjkEMPi18w1ESBvtUPxZq+zafsZKkQtuNL6z40F0/A+9IB4Y0d5Cfqkcymn
IvJCqmSYBgWajd96ul/C9AO7Ik5jGAriwGtwEr3bHSQkkXFGDoTWbOs/KBBj54uj
Agi64AFK/JfQOLS8jhEqPIlCFcFu13bQlPoFwctLqMBxdcaoBNKJg5ex5xxY2u/K
RPQtDSlhSMUaA8ySbWujOQsRN9xW6KyVjf9jyf4x4c/9lwx7JA64uKlb/Qr7g1Y8
8hue9yIP6yHMraRkPhJr9292yQWY3k2kHU4AHtkNirTuTsyPSe92CdJ7KZisrIfD
A7x30d46N+2Y6JeEKQpqWO+GEVdGiND/4++nk1QjfivMpub+tENrlOb6gkgaEPLy
k0YikDgnoHnph8DnNXdMXaXdKdDCq+mis17h61fXPOlTa/hy4XI04u9dJQe9Ib/E
q1iE65Lwm+HH3ms+dQsYwm2F7xlDcEwQ6Jt3FRmE/SmbB2QS4RWAwNq7/Eg9ZO+i
1Wyg+T818H5+o127+dkUmLHvPX8DMw91dAWTdGhEuupftAWMjHso1vUxgCJY9oCp
7LdJDFn8I8DAahrNMLDpvJYYBMNMZqZDVwJZAWhDwVk7i68ym6rXep2yoOImccoI
SYExk9iQA4y/6D+E3b34nN+qG+bTk2Wk1+pSKJj05B6UVvcuT2ufWVoQxhrsnZVQ
/xGxf+wvyNKJL9uXh1dof8GJuJBIhA9+sBmr+sfFmeIGr5T/de5wfo2A2BqtTSjg
oSYOELp5XCYRKh/2IjsVOL1li9hEmIbKawZbHX62uZ3kmjC/RH8EBFW+7OVdqMp7
ke9RI15cyRS8+ymmerD0p3DclbmALjMswpZOBqH2Z+2HIrMHzJNHYF8YkVIqnDQl
K0bQztQUv0XIWtCb/xq6lIwApkWLhLqivTiOYLZh2SATeGJA4UedljjkNCTdmNYj
cESfuHIe7wvuoDgrZ4SfRa8E14spQna/LB4DmJDPIPMjbHLEESQwSCwgOUdAILr9
D3Lz2qv+ch3BR5ptRq6eX7E+M9g20hL/rwCBDNqarjFuUFnAQ3h0h3AYItp4x7iK
kklu0Onx3lZ/4Oekw0cCmfKyNYxC4cjBnh9FoGCj0jfYAn9mjBJRpoevSnPeVu0/
2r8BW1TK/BXfHUfiH9IexfjlWkEhr5y3mInuXnOkD7dYqXqCP+lWM994a+rFLgBF
hcEwr5gxfdwyp9mSL4Pm6vvQt3JmD/OOO76Ojq7gFdTK7ug8VCzUHxzU5T3ZazWv
kTb2SFm9MMqLSZ3fjpzP9e26LHIUCR8aV7DJIsSCfqrVaIERj7Z/o30iGs8ufp6c
1rXCn92OOns8nGV1WWKsyaIGPWFXyEdrE/BdZh3I0OzH58xyHEf0aGLu76IbRVrz
ILGtc2gWnyvDF0fJ6X2yfQcxti1gqPFYvegdoqeTDyjGYmzvuUczkanTFhBNGPwT
MZ7OQavTSb3utMdCLkJisnhePv5CW9BMHaVYbPG6GSgdBjZMcnOf2KK4LKjk8Trw
dSKSfLX8txD6Me3gm/zqVehN9EmYdYuYcrwOqrCqd8haoQpYuabXs1cndOzgqhUI
t6vMGOmSwsneqoxNqlXFGe0oDLwpUc2RJIry3IzB71gx3nj7QJcvcDZqqrE7HDH2
kEF7QvGU3aujCpFSZFtaXAxePf1FcLfYGb0dpJOs6uMKCfP6wgbgmdbs0oEciQws
Hc7Xtjl/CFGQKEE58UjjjlYPP73lm2zvK2H2pMW1JWA0PMJmE0mmyoxltsYo05oC
1jbnkvIv8vIG/6EL13B7UHhmqXNEImweO1ZI75AIenWRE2VP1xjKuZv/7ounFt5i
gOmpwv01N4SkUxoPC2mTRVUBmcsk/scnZ0yKN2M6mw5xZ1NrbCvMdWZKU+OfVFzN
bfja7NueJmJzqepWpwLX5VIZChBaZqBH3Y9dqFPK1hjhVV0QK4q0SeiczpeZlRxC
z9TLO75K1rP7oUjJKykJwTIa9OXISARcDEfCW+o2XknQuYig6nqfCsT7B7GCr3HP
C86zzAb5AYcL1YW3yi5PHPrCGDqQLmIwmX6RiCXL+XwntbmXdn9t/lKS2Xcd08Jv
PrDXAPoSro4tzDXURTRZqqcj9MB/2SfA8e0XfZgbUktQpn6PTXzBLH2JPE7GJDPI
aTu0s32aK8sg8zALwQJOy3u76fJcbUKG6z0ioYaJjfL291Dr7ls10Q/+5KErP72P
3KOH5VPi5IOvPTE8aNpXQ51k/EstuZC33IROE/owbvt01xREt2qkJGEk3ybVOu8N
lkdJF+SFHRoHhUgjnWcbCByhQjATDxtW49xNYIqDtQrHrBYxiZ/qSmfivMSjFN75
TCtAcJj5CuGwIgsBQB0inN/at92BxTPPUW96/kH2wIUbm2+daPEScDF0yR2rdSWM
GdNM2dCDzpVzsALiyWlvyIEEhfZeVx7CJXAfm3VehJXtHnlKhlHy3vHyckOawAeL
YFuBIHj77yZawqwkwwRt/MQZX31iMSVPv4EX4kjE2n+WT9QrA89TekU+pEJAtGQT
RyzgKu0SZpXNEH/A0DLg8qG1FzC84qOicWG3M8rgVNpz9zIRr1x0+JSZ0W4wGsIN
cHyiiBhymo779mKkSu9cBEAROyeFckRtq7AqQMqK8xS1FIb2qOoPNHMOi/VzXB3z
fEDiZB8SIgwTI4wG3+i4XUagqGwAkRGTIeBrQegHP2XAaFygAUSxtiYjzMUjEFwF
fzEf3PDGkfy/AIUqxvUoaW2Laq0IYQiHWW89wkZh7OR2arv7AbHcQjj3rp7ds4Zw
wlp96Q49isAsFP16xE3c/3XOMLWs58y2ZHL654FIYBvvOR0TCqacCI8frGdl/1ti
moWwGGp5LL+FZMP1TMsFVcjyWiPDtkEFePMOJsb53ZQzpqXXpJdxp3kc8mgiAVNS
E6/ROV6RmXsKoVkGvqb1iQ+61b52NgyQP6O65/4pyiMN0UfK5jVvCumG5hH/j9hN
Bbj4jVseiVMmpO5bF1St9Nr2nk8vLVdzS9CeuOZjz+7FpHQsPuBuhunE1Od3GQmM
4iIsmRCmdwrKSYEsWRIdM9Gt/v/K3lh6uPt0HfjgFY+4AYCHltlmDNFDTDjMqd6F
MdsyNgTFj0NPZS+eMVU7XIgo2xkaqzZausizZFdVH6qs8rqsE6bODVz/WMMT1cno
8CuylQJ7wEv7ts4ry9sYsgkpBtlFpWPXSI4r5W1lRvwmIunKnGK6P55Xa8kx2qMh
3CZA+TSlzCIijduHF9DpNvmRqQ+WntgUk6F70HwXP9+dqUJ9q/gGh5syXbcAcYTF
yj3TaaUk6sP7N3NcIiVfs37HOdx3YtkJvFZ2aP/t8iSwnYQLWJdpAf3ldZr5/RC+
XpQH460aSv5xhspwD8kpoK7R7oLbBs4DwYeyxHpx2gbafUjGrlDTiuOnwKp/LNkE
u1uKDGC8BsbvnTRpNC3aSW6/4XugOYf6PIR0qHqMtG6D3gTrDCQWjvtlmpXIf+gU
OKXhAUpakk5pqQnmyoxP7kiMOPUl6CVeVffMX/H7aa3ac3cwQPfm8l61s5D+R11V
EgPEf1iXleRN+EqKqyCLKAaO24rmB6cI6eX6Khmc2u8jHljKyluh3eIflHfeFUUJ
LV5jgBvmb2BFdSzqkhnuVC+P5iFPrij8K2Rd5aJdvCFxm/BXebXY8sBrZwzfdO+h
YerUiBfajn7/l0daOqLE+9vcXbOXb13ZS84Qt03kgV9lOw7NZQA78zFus540d59V
68mK3n/1FhohNXTqH+JxylarrDbZpzpxvvottX5tNJ7G4ZCSF5K3a1ADWo/O5SoA
z+KXP/sVEFXiMYh/Dwh5YvelfD2sg66twgvQBQlZtzPnB9EtVDH3Ld015hg/ictg
IECn8Djc7j6j00bJecBtq6G34eU3QKzJwH6h/A0CB41ekcGn7NWpJUWdAn2RyvNj
6mscjw+gVSeyVvF6yHB7qok2o2VY+o/vVhp9LlLXCffSBCmbyAzE7MZklhf+LEYf
Qhcb4bj8mWk1/VTaxRG7t0RLDTivbc3I3AEIpas7DOr5g/iB4iPbXAIXYfOR6P/V
3/vWpD1AzS8bBgPW0zV/wkNq1b8za8fvVb7UZH7+HISt9qd9PoVD9+Tt8y21nTXr
DMkhMYqycurtiwAIK5UN5VFQZw7ErMD68V3Dj3MkRDA7NgACpo4EsdoqduNHEuRG
lsvW9wS2RHQRLNqHqbMr7DGpVlHUNEh7iw1DM91J4DCmqNZ9YWX8E8QmyTRd4NZW
rTK67v1/vSmAsb54hshSej0wF98vKxxc0LY9tcRSVLsjL4fOzWDRY0yl+GW2sjQP
jLDgX8O7oWrWUYlNgMe7IuKE/NGa1d2Mumdfv59+Ys2PpQCiwJoRIC8zibCZsmYl
GlWlfTfpmujwmMYX8gG+8ItvTabWPjPad7fee/IFfiI8TO4CiA/2K7s9qJEUDrEq
FS254J0d375JhZwNPk0+L0qbA978MHPuf7Q0VYgXpzFbPUYJYJ2gp0C5nFQfldQE
Q4wDmykSxkntFMurXCtHV+/swyGisbBpCd8yRHcIDzfjeay3YNu52n1hcwP9hI1x
gswsUV0u8BV7JEIwPe1j2HmX+MMxfvxxE7zeP05ck4tWH/vICgpcBJrdPNlRc06g
pjuN/1hhtOWllv2LTBb9WWa+QOe+S/UqjToNkdmF+wP/E6/Y3Qnn3quZu4lckOpF
upAkr8vwJ+LTZt81nlpbsl0Dtdd8UxIksUkmyUys+tvS4dECBJcvr05CGvL5tEmM
WzLXa3IVyL3G30irBNUdOiqv//ttqm8mo1XE7LJ6BeCKZQZabPM+JizhaqPc/1f1
nGAMaYSdYYusgLxXafnwBGMUae9MKSgmcK+/Hbz6t85qsslx//XZMCpMlBT6/pKl
NaP7icljiQ68MD5VccFu1oQIm3O655/gOvWP4hMFam8GFZ7hWLI2TwvtQPQfHSf1
lubpFmhrAHkTh6S7StkZ4nJ+3I7Ny+kdXrsE5y2Xbfh3nOAQ6iKOjFpmVw5cBZpR
IbyCxKPX9ioXXrMArGTFquO9pe5ZQbumAG6xNovviIkvzgsNCegkYg1OzbWzGGFI
KH7X81uYMwQ1CVtPmtwzCHTCSJaGYg0GH2Sud3dpvkJIFUlNLDT7JvIM3iKPszw9
7TxoK+wHsjypgI3ya3OvMdXK5GDmlOxKiH8I89xzqYksrZaXI+tlGBx6JNyZ/Z0m
B8LzxumqDyJI/fLz8Vt7RpgLsmaWugyoDrSmVZSyNPm3VDhG+gR6Qn/XRcdU+ngp
+D8PNUYbotTtix2dWfHJHB/+cvKy6AS/M6znnHN9XFjXiE1QaKuHcSot2xP7UETP
CE76sucTWyNplUwIl4njBC6H8vtl3576Z9ki9+87JC3EkPsE/PdGSqecRjlUGmJx
bEGpMbQTSC894EaQoIr6pOO5d7op2s6nT/RIUinePLlTcH+woHZz3uNV10Unna8B
aBl1UiTgu0jLRgSa4M/OlR8WFY+WvfMjQVZEkC9GWF+Nzsag2AYWuy9mTxMaOVHo
8BsQwF7CLZFYOAl5hnBTJGW2MPEUC8O/Dsynfepi4LjvTRdj7P5UaCunlU6Ol1dn
xvv3o+k114iWhESXtzk1On8yXmnVj+G0KIBli2S+p1moxnaq5K5lYcIJtADZ0XMz
dZw32yoR0nmr69zvgYSJPKIFmEOa2iuZCYxtn6avbmc5rUbDjHAkSykemaYMlqCa
OCFi4MOgF1s8ThcX3h93ZmAfMPWOqUeIPnm/KBqb953mINYObd6pK681fpywTTbL
aSwMvuyG2p/jOfb928rBaWs4EVRNaccf1QuT8YWsKJD0eMyJA1NCIA3JP84RKnN2
wt77YOQJbyTinORHeQHeop/GdpHCjaEnq649etQjAdsjESpLVXbNhWsIYwnpuL0m
6Emt/vMVogec3LuERLf8cuDRyBOo1BVBFLGURPFPh2fGbIS7Z/gk8qTJkPxDlwod
CXsHwtaYy6A0l8+PbI6Vkt708UkSg8inZeaZpASXR4++1aTb7NWMytG9+JkXUluH
SaBRxtfBLz3bYIxwPkyquUK0QazpTrF7qkFDpiylo/k1qynDa2VN1xnvIR8mruhC
NKRckPzMBHx1k6e8gEwhY1ehT9FC1s5IN0W+wEdysBOywZZLQi6NiWdv5fZKoLle
4H7HH3EQjcydukWeerrtSCQOJCyUcTaHStrUD86fZJqo5ikUvHt+cJxfhl6VGS0D
QWPdnTs983jDuzFxQEe/b7qw1qsI/IRz03x7UhOp4z48TcyO7/LhqHKuKDOhk3qv
3w56OFXVZDIQBPeeEnnnjB4KjjEBREf66DIaCErH5sFpPtTJod9h+JATuoMyq04T
7ozOCmjFvXJjyF+D5FzJg0HYb43auiKPdVP1tdUvdL0HwyIpxW93m+KIa6U84pNQ
JiL3UqNr7KBUrArsbgwQ1lUjcK+xNuYldARMKXo1To/VN0rQBMO2DJXNPKX4bizq
zWmNStmKmD00leOruZ/l1DMTkcFiyvt8/QB5iMXqP5NEKTNLkbBbikjO89WGtZm7
oeRizy1CA6AqqtRx66Dtu+mT8M+XaKRFhw0OSpiX7LHU8fUfugYtXRoSicMj2nWg
lOVAyxRM7IxuPUsV0AIZsg3VJkGr/4Z6XcNV6JNmREceldVaffKJNiBKocU1Kj3e
/8v2hP09x8FL2BfSD2OzFtbyDPHJSNZGgYmRgeZs6xRRhDCih6qUas+3EzpIDeb5
bHTVmlYTxTu5bxfMokF1ndv3lph15/GiRB/T83fi1kz0eVt1I8MKkMPTrQK7aSJ7
U0qsUwhiKdAKLNOrH8KhnQfNs/ixra5XZ8sNPBZiPtcH97bC/KYXScrMUlJ0JGhj
QVndLioR81m+iv6vaQAeO0XPIxaWxDYfEW5MSK4UvTPBz8SQUuuFeMVMJU7gPKB4
CxGfT4aUyv1IbiRIq0LwjhmkZbCcdMMIPmt4wGZ8hH23EC05wBFXTc/krOSTZj/K
TMNPNoKWRiXZ26Jx9mDQZ7C7jMtWQiWV4VJTks+Q99pmHhY6r+S+CBXhFp9dJHCN
Rtt9ix+bCtFZvZxV6WfnVwjZb4498VRMw9aHWKm5q6XHWulMSFSUdtFpZUtm88wH
fXTaHelRkgdn5DKGtwX342lgpLrMZQVYnSQwMt3ikZGT3eN/VrbEF0rqzm6VZvA9
0NoSh//6vfFnDX1wEpA4/8dLdVVtJ4qWSQisvMK/IyKKSI6P8YNqHYnXuSm1hrhv
jM2xCrTbrJk0PbfMT0kuyVKNmkfwYYFJOn0TcKpSz7T7vm1jI56dB5MlDbzO36Qp
USBNu/281/t1CfjpTVCuyo/T4e7LdIl+Y+Zm7pEB2NAJmtWmhJ71YEtgMVTB1NuD
cuwLqh7NStMYnRE4wDsjGcgdsrgRPcET7nbRXYezLhNLlJ2EwmQMcFRDjGGPxuPA
cMm8eHnlbJ4ev/OVGoNWKuv/vUyPA6eIus8ZGbps0tXxafpQlunX4JJqMnLLRiNY
K2yip8+c23P7fS3Zkw7cHYWhnDyCGjz/6zGH1sPmMRBTgnPhofyc3Yu9UFOhTA13
3HPWLeQ6p3QNWhoZqDXNvMazEcY5gSxaLrk5AyQXiLv32iajiiku7jhV6V+U0US+
gwCjzia/x11iHu2ztIbmbIB5JjjuWmbCOTR5BTg81U+sJCAozpsYaTH1FoiGJTYy
BPIOozu8GMdX53n62GVsA35P/iu+2iqcsvNY++Fj81gaPwBa9tu2iin5gIcHWXdn
TL85dhTlfVDODlltkxsHJIJ1VkDgS88Md+TwZ84izLjkrCyDf9x9j2fYvR1+5Svn
HwkKRZ2ScG8V7U8Cex92N7zRsWNB/XHI+c9GEWTkM0Ez/AXBys8j6u32gqcyjQnW
cpuYZdeKq+hzKSLZOyiQr5oSrriRK7ywzBblPT0Eg3R00jGlBcSpIl84C2piF6u8
s2GgmaiK57eeBP1t8pxddBVMWVkjYnxOhrxi/uUH10yGHLQKeIxd2TC2cwvBLWRX
MUe8R3A9O+dZkcGyQFFOp6IS0YfVBujgEe9o6kEYRuAVl/J/5Z3x/EKKQ6Sm16Oq
peiHIuJtgDrbnFigwgIEV5uVclZ2Pr1ChB0zDMhLWvjMsUxc9Nspc2O0nntalsi2
lo7D2+AmMmXgk1yo/rDk9gi0BqYaFBUHAZuWyoqxEmnzlxfNxCQsJ+DaJezer4ai
qJfqq88pvNmWSNF3hI6jiss0Mo/yll6ngWRr8M9W8FYg5fDuTdiQldYwg9JuhbGS
MxJPAI1FQ/VB0N1LrVIeQMvNZiJHYMvbEsGUtdRaSmllR3FS6D/y8rzUCzzX/Fmw
zNOoKfj/SYsyuZGcv6nDG0veLmWQlyRWVUwutzilaa5WjBJNEbYR87l1qVLSrhA4
gqh1wEPJ5S2NK+cGU3imJUcQn6CItYI6ZUuv/BMtgy25mdywYSG81U7eMQapA/K7
uRtqYvx3oz7eQ8LaaSboPBoYhd1FhkEUuulm2+AeeQvM9qMbNfohxG5JuzouAfzp
zzW1i93D44MduqcWyhMJWGa5lGAlSsFxo5/OVrKUi0z9xlLpKByTGpSV9fSBZ2P3
sbOcfuTYlB8vTit0dTqP3pFZC+PsDxNkdbLMdIYWA0r9Yb7J8p13Y6/ngbV1B9Wi
QJ4AGSTAEC4ULgfcLxPfsNcuirmEzNx/vpojeva1VSbn/ZscgSn7eujhNIyVd7Mo
udOy19I/+Cns5H/bXmAoT4ojpyKqdR843hPy0sutrN4Nlk2bMgBonOwsaV/JiOJP
CBVKoyql8K8XTm2KvbMljG3MlD6tuASGdfWO5IDUzAy7zl6xklWb4kPzuFpFea8h
M7/RCqSwExOB/C3e3eB/zUf4Lxd0iFHLIZz4lepullmPLPHoZctBrAUjx+oLroeU
EIdyw6Hr5SnXvBT7fSnMvG5kdFtbssCNjBEMzVfEx03dfjRF11HgjGGkybx52GuZ
xDp4QTIXF0Ovukz3JYxhSJQ37RGOGc7+ddt3p9UvxOl8o/EAOS6gDi0m5BZaxLVB
DNQA8xwwBhI9lLU6ZiMfJBP3T2BRKBKxvoxXCmb7dlwEXClOEFQX07SkrjVv0P3/
zuln4xYhroxXpEnA3Ecc4OJoImZCm6RrVDLofyUJpN8CKECiTNoiY9+gz3U+gblE
TOQvc8XKTdP5aNB8JVGfzVNo7AhH+4yhK+erKYtOi/0dsGqoALP4HsuLm0cqBb4p
1vsCIBw17o7EcQAyf23IXANA8qpSMIcDe7IEQ7UKpUdGcQgh5fKdZE7PslqdFIKe
nxHhtKJf5AY/+WqSeMkiXYa0atDAoaNTFG8BaaFJiihUXefIOC5TYY92if6nRlqR
WL3nzV/EN+VQHAL4nf+G6flmFeMDhybzn1+cfyvvJ2+EtamAEE2FUW7c1bXbFGme
/VHn0nza+zSv4QDwer6O4I8UEojSAIWeh2+RrBFpmBqzYjgrxrEB6WcfHcg2Rwbi
QQrdmmxHJua5buL0xNAFwvVmrDh21Nk0Yt/O38BgFvPBjtXC5G5kzvsiFL4/htT3
+1PAZW6BXrgJpHVM6aRhOyFpTh+3uV1sOHnrT37swkBvcte6kmcQ/a80wXd3MhlR
zA9wfDNHagjUtFFtVSEmLq9nWIT5BCrBs73nLFmAYUWQu4JxSj7MWJ+tck/fZZAf
R5qws2NCXCEwKmZQvlIPWhrYvdKulTl7D/5yF6d49p9Z+Dp/sbq6ZImjIXnPNxQ7
H0kTIQvH2N/PfXy9txaRL9EyHnp4bIhqH66tHbG70TsrMCwP5AJ/S36NvGbfhABk
Ww1CdknRRcZ0PjpmF3ORV1LIsQI8/qCs14jvN8+/zHK/3oVIoEQOw2YxAsE+FD77
Cx4Y4ueTy9L4Qz+iCVUQqyebNFYNEfgvfPA+4UswHpBgHXAmp1PSoFR6qWt/FJpW
+r3tMf3Oqi4SVAIFoyA+tJbr6ozTJ5BDEJd4Yx3k2EFmF4md/iLvhaxrZ597mHJN
ry9AvVYY8pIAcF1fYaggoVdRCJ5L/PLLtAL2cig5JMnhIaq9GVbyHkEyES6H2j8J
9S35oPnobEf0BzEJ6EX6jyS+9+eKN+4Bfuq8DyyZA8IjUkuhZZhEZa9hJ4L3Z47R
lUKe1Qp46vi2m/g6xLz9p0zh7DqWt7Ub15fQgrNzpG/Zze0o2YJdUNyv7ukqlNdX
jZ84pOQxVHgNlm9GF+XbfgIq3cH7HT1/UaTnzOQryrGhIFMI7jAWoDmyQmvoERZ+
ymgDaZLWbLdULo/qbxgLTZ+RCTtyAOdJeXPc38BPH2yJoN5u1g4DRBXh4uZwaXg6
tHYIzkyEa0hP8F8AO6HBgEviHz402bBvMOB+hRMkkrFt4aOV6aJ/YBylFN7alFyY
SwDI8hTPgJC4PGMi2BqI6Rk6nrI3I/iqUssRLaHw7vTP3SK+UC6Gj03mqrP9O54e
P6sSkwk1iVfzE7lUmnGmgr/4mAcO0LOr+8A0odU/JRmOVmcCDMohHaVRTwoN8t74
ZWBtNO6Y8cYxqRISFlud8Ay++h2+qYHZ2JzGSwx3FBhOz4Y4lM1zSmfWk1H3PLyo
esa7W9y+StnkRNOyLBDyGeQWat/V6+b9PSwLzASUezlpJYMpRboAltq43rYyW9Q8
KKscc/AYW314xEAhy6cj3bvQJDvM8DSXPXEjPsNX47Q2I2vuG9ekXkuW9mQc5cJq
YXuG/PhwuC3alzuEtt5rkE96VpQ/BPsXeAxaJ7GDp5YYLxUhm9TntFaPSnRrKEjb
Y5Frgs1P8ukwYe9rOtqwiOAN1fWjtwnmVpYeXypkiI4MU1xl26X9lYsc3hKqGIUk
uhFChyO7wpqIW04MAXwJwyBbZF4Ib6Xf8e4zJbxIBsUeEomk+qTFCs4++Ksx1dDs
TiruEnXcfRw3iFKyBFgOXh+hY9h8zmjOUZ2mub0YZmrTxZDXkrmwRlpoBmO8mkvi
9JuCX78RD36CXu9xQO9rhXi3LoCXfvU2fieQYjJSURcOH9Wjzn6BxICKJ+INVMZ2
GBx1JSlLYhmH8+MseljCDRtbZm4Aq23ad3PxZp181c+UxQty994PGf2RGA4eW6uq
D8QzKByR9s7mF0oeWLGplXsFGj1RF99oHdCDxlsgJeyJRG6aLjXysIv9pBj7pO0D
e3Hf2XKmdgzgZ7623udwa2xXDOEqkrsCdNFRKk5liXSs1HzlEuyqSMOqqD7lBs1c
wJAXEi2DsVlnOY3EvuJ5FzByyh+dThvn/OP4FAPxM2bzOcVsYw74ZsKZX3WKs4eE
Vs08gWVolBYjhY7RUuhN5GysPdXlZ7b4FxG1u+bhPFcyRFOwrOHvLqgF0PT+ZXlE
lmfV/ntMp4NriIXfg7z4WFSxyrEQI0KJSx89zytfpYUeNFBlCwib3fGRfOhO8C8R
YWMp8WgyKjIzewCS8ABnXnwfN72GbzVB0sEWobndix5r7scYDlGZ/Kn78DWV5T0n
0kYU+17qKQpV7D5tMZqID0i84R30nlAEY0x7gFSwATo6DG9rewRnSQU8YRug/1lc
kZEhmiPhQQSyzOSHjpaIyj+HsP/jVE0k8GGL5W1WTEcXbL0XivSk5m7ExwBTltS3
LtwKxq/H+D4KnEJ/+7+1zvMYDo8KgV0GyipME9MsyfXfzBSrD3cDFy2EfmOdwuK1
wTW/8ygvwzfUxJKvv2nPbSLOL9Wmmb7OR9wA9YJ/T6ZSWBLZg7Oj6t9E8yN+OOv3
nz2B2jKepaHAcitCpIavZkWgduhMls5/OUbi9BlW/4D733C08s2F/3dR1jMzLPLF
ogX58I2KNVS3poH5CJhQ2TTUAyFsZjbJ71lUG5AgdLs/pF0dLFpAwa8htAfzkljm
G14DL3o4P+3n879172ksoI1kUkaXYxPIcyHXVTr21MK0lS0uLVS1ZWpcs8gW02xe
VxjHsl7leTXgP6nEPZQ27+qVia1i6KNvSoa6nzOpn/olx1EJxL7+MCbXP3m43FiQ
P24bgYgQLRBQzThwumQ0A/RbQCKZimAD48GQyniH9NMtni8i2nqS1pSnRLWm3hHe
S/vVvKD39qLOR4/rsD9xw2RSJS85DDe3GkDf+z1h7PKMwFEfYuyepc7kjS/Etk3n
jsRQyzxfukBKSGktIcC4zxxymPaA/1/SbK1yhQ33E9SAbl57YBUt3K9pDhCnfSAN
9GdKJ3aKGH7ZYERNHGHKdt8718dgZv5Zm5ZvWkutb+zRhrR4g75XyPd8qljyhfzG
HbXHf1neL5nSrMjvntPokaj1AtP68D4NaNllIAgiG+XoHiz2Sz1BQLpqHJYO3Bly
cHmJOTIrc5m5lXmh2Q44EG7Q0gikL9XaxR+qhJPF/PA1KGoCZmkqg1S2kXxC6OlT
nGt3xuUrSPbHOzkWh7y5pt4SK0B4lqTqLzvpgkzociY2bzP7rnSyZuawwrSaiNFD
m+M1iFIe995WGLNI9WxL1zObyzqZT7Saw9K+5qqUUtC1bFEV+/qM1aG+77tHYIX2
Y6tTUZONP3/9awceGG/a4P5lgFoeI4DQFSCe5xr4bJjttvPfzHMdmetAM7txfoFO
aTKGf9IaZ3+bXlCdUay7mNRGuLE4bV/3BVJrYcZT06gLyz1dO4vFfnTO3QS2YVGp
ad+vJzdFPi//mAKtnC9CY9yuJt6wvNcMZXAJgXVxtddI9uCcXs7Pp/2V/I+O3mWT
ZbRySixl65JgC+81xapJr7MovzQZrHXfJunZ25quRZeZCfIWjvtYt+76VgxEJiwX
zqvQnvBPTS7bvhVwllWC5kkyfonau9PbjxItV/B9pRC4s0a3o3QhWpuhzKQc4arP
CLIW1OtGf2H4MfDxEoODZpJsAehgxcnGhUDuOBKASKDyk1qu8KkywiDBeDoPYa2X
yaKVjq9k4VGKgGNAOq5QM1vKfFUdpHtbTgZb07C/IliWtiIMYybCn7XmWPiR5x1z
gEFZYgrfRXda2mIr9R7o2RmLhCZ9F348J1ZFbAuh8DTtGvbIp1l+ghn36gFnOGwd
P7s5nvG59pf7Zge0KpVo+yZyezeQKvK493GTsCfNxZPgZBKcqukMg3jwKln19ouJ
+e0/Hk8vnSXpBf38MTnK0cCrxzNwCfPd9TFwQjgQbS6pXly4VWWnB9ZJQe8+gPow
7PehvHErpP74zavI2Y2pvcsvT43kXs371xPWfYZEhsn64lsIvx5g0ThX/uSNJw5L
D/rbRBpQOBCYwwGJTu2Qja8vLXV6OSn/+cSdOqTlaTWDqc4/teHLr7JhEcWQNdIu
fPBbb7FMvpXhO5iVXJ8PfDmSUvhG9eMb2E6wVdx80DeIu0kgtbM1QevUBD8ZofEE
y2VUFV5mITGO8f4f5LFYB0UHgJy/TcfTXD0bZ3qDkDLTamHIqorZC45uSe+stotl
KHHMawGjxgFmtMRtp75IM5Lwtb/eQAMdisPT/aP1tcPKeEQWOMUU5g+zJosCMtRZ
Ahpn4rSN8KWFgAc2Hyh0aYba6t1ZMpgwocvFum2dLkqFgXD2wOB6QDHR3+GxoOAi
CXPKU1AJBg4ocRNRpe2EVRYgGQ1ZznROjrlvhBkUisMpEKIcuEbGZMRzD289e+Z+
GQP8hRPc3LYqrGULYt7M5wiPUW8Lm3hSmExnuf4I9WeBuelLbsKyB7kIl9Z7VoDy
U9DpTqVvP0PM6jkuVE9ZppgRufUcExSEQw27AuV9FuGzZAc4o3GKNNSSpgZEADNS
oqDY9qGCEDlmtArx2w8QzFfAcelC+qpzVlQtNJ9d4Yi6/+sMO4Avb0TTHebnD86z
7hewpO0FluN1LvWiW7bo2zUlAh/P7mFQ4szcToijCB4kK2h716FZP1cH0Kkg9llt
DG2tDoxApzOm28A7iU5ML7knzepPSHhX7+Jcppl8CrpaPg7P5TZWH6pCZhUvEIod
WHPMLhyTd2EhAdeGWpU+MUZteeog2LILrQ+z/HskCi1fun0hZ3xbWiccfQZQBjfi
N05UF8Uyybvl6urEaVKhUiHc58MCN+jMZaXbWTD+M09yAKjoHn/hN2ppH4u7kUME
sgtxm8tiLoeKa3DeLmYsCs/InL5YjI40UzXpd9eF1LSPKobNbvKIEIw08vTFJjZ6
FIDHWO9oCUJX9e0lSlptiPZmeuBX+CwdS1iUbJ4gBkPagUJk2wUR4YfmcRZalFMJ
YPDf2Hs3s43u/jdms96s5KI/AdV3zWl1zJmeXYnBeqQqYC/8MBsEntbOhCLX2U1J
ldXTRsR9FqlAUjNEykDt5CD1tukMNlMTabd1QK2evIknnU/oBnoq2z39aNDo8ORN
htba4zg1cw8PZOzPbgc7qPtJXv712MespUeuB5uqOXIGUPUxhtie/f3voZKGhgF/
Sm6rbnGKNvRO2OILVHnnpoYBZRBy4uTtOZ+Qr5u5FMGX3exXfRoZUU4pOxGEhlVR
oVLCmuK7spEGbETDa6VuyXOBI7l77KArnm/XxAVJ+Q8er3b85Feqlt2PimKW7zau
JB457xHZsDv8+6mWsvujYiBfM2T/o6jCTK7sqcpt3ZI83qVYVRmKplOkHbAOOXIj
aCJPCyMw+OljWYvTTT+5Lsl5nRl2zmM56wKvRrh0cG+hl1HlN0BQgwiag5jvrUKi
hiZTgsOfnmLb6uKCqctb9tqpWx2/QfB1E5VVZOX9d72yTA50G/B4j46Z2UrfNeYz
YIzWf1xB0JdG/Gv5gFoazBLD61a6TmEM78aymyd4GpKwsMBVLyS635p9T4yJPhCG
uai6P+zhS2WE9yrBmj9+bj/qJp2fHWDvVapMkBrBerxxlsKhrPwyNwpO9ADlya/C
0jX0zyoz7GjwFXyorho3wAe3BuE27Ub6IVtob0h5JSDdtMfDYdEtJFdmVASAzbm0
2uyoxz8EydVNpcUzp4GAfjb/fBnXBJgq289dbJPgr4MpmJuL03nR5UQfw624sQp7
c61xYWk8o4sgvaj3H6N5i9hlYVfa7bONj6WgEKp2p9yMnS4Ktp3OwrA3+tPjmxtL
iiMVtORyB7TnHuzJHCL7310HbQtKVvDRXG8JFTyRjf+dhkuZ46xFbw6Y7Z//AmjD
oNZ/G1Vjqk6cAbnd19IvwJGKnAU3Of/Fb1M6UquwbNPDbaKtRNjlB2XRBeMxTN7M
S2RKl7u58pIxeJlG1ZWQWHgG765L7vCXV2Shhttk+7Z225FtoxoyJT72Gzj8Iklg
Wcwk7bMM7M6YmDEq8xAcvemL9hO+rY//aQPrrHCmm6AGaFXe0iRGMZ9pp2GsbGwm
AnJABTkOVtmJW9r8gL23nQZjcURCCSQ7XtcuDOJBwpRHJLk13WAcYDh++upNYV97
1bg91aN2KDsmrmKNDp4neyxb5G3ftc2NKhQbsUmOsgthvQ0GeLBD/ilKBZr0pXKY
5/B9nVYV3fHYrrzVxJxxa1DcwZwfrMD6VFMbTO+Wql76xy6iPqJHZ/7/uHAgIOn4
31SwPJkw+Mi4d+falPzzq6+5w/J4OfyFKWlIChmLnl/CssOY3ueiMF5WNvxB0Z7R
uHNSsF2mEbsIGt30YuBqiKu5+Cv+oxWe642BX/1doAlqc81lhMcBaBFMYMEINW4I
g3Wwe3g+rirAi7LSccADaNEFJNGczSXU+WwcYuVRL7XCHvym+u5kXSuy0MtTTCwf
pb/5OBMhYzRUraXkRk0Gq8Ck66+EDPVvmTHj19dpLgHDMlscJU+veUwK3mQRqxDH
Rxnmr45i+ZJKqVXb0LprXv66tmahn5n2snEYeQR1/+kdn3YD9SdAIOISjyyjhzjS
pAAO5NQaOoVbiBcQqSlc6D827AXEm2mmSFK47TveNPmTFY6hyGzaRBR06+s5euOr
HvQ2xyq6ZC9qyd/gTik0ulzNqyI31wMjLU04gBwJeYyElXgSh/VsPGZpVcLPxOcN
D/s8jf2WkTwN7g8b2R7ylkZwzNkYkqIhQkDAZmE8M1klUWYXxRndCCRENG2hlmA3
noqXs4OOD+2s8kmtHNKEZP237vP1sN8kmQ4H03gOMC0EMOFoJF6jjT6e2LMz47R+
vZZesy/YE4zdIk2EWntlF8Mi+QRDILyqXcHjItlbqaXSWPJdy6Vf01BtE6qPmZPj
IE5vk4zONyEdKXEp4L9bgUxlc6plI6nVIsBrqKEaHpU/OvKq8vmea6ZcRR06eTBY
Pk4FkePm+Hmm7CI0dMbMzTjGjSlDCSd5i+N2Rz5lBVS65B/O96o+2NPinMHqTMh4
jEhlYrJlqJv7lwZLhA4e3+XR5mOpazPTM58BsMdElvlg5CnkK7JxtIjCFncRscbP
O8FCxtuvQykc3bNZXmF6RSfxrcmN+XoGKbChp0ohv3LXQPonVTGs4BpxsRgZ1vRV
QROgsM1z4RKHl1Pnk4QaxzCderdVOkBkmHmJyHICl8iQo8rJ/Lh7JRpwrOBPI81Z
0nuI3O49Uy78KzoLk6pzt3K+5Ozdg94HF5+XTWqxkv9ijbps1PSi00TRHFNyas6M
EwQcXXUzcw98HW46QqNaOIYABe1/K4TQFTP4k1dKZrB2Dylz+dpAu5J3ccXgb4ZV
B+vr941bNabi/WGk2vmp3KQh6qP1LxQn3lne0Srgm9X9ZGBylqvZAfq2GlhmWTfa
DdB3oOquBG7WCPDraJ+3wUyorB5ReTL9z+mGuFNn/Tfs0D/KOSSXVjNtwUhJTEVe
QC5SYtUHMlkLirZ5g/h8B7zkCBFjd9resCnCbp81oQc9VMAO5tWMI3KKPSNlTjTC
hBayMO3dGuDTuZnHRlT5XIBR2/rIzLYO/8kI4RoJMI9y5YhnP0BdGsd30xGpiFrF
snAEkRpBNMdcbvIQrsltfwzPi8PwU90IWwq+xncQZyGTK6nudW4s9stzfvA0EOfS
2jTltshukt+UWEsHLJplSrfCn3ZhU2I9wzJwJIYD8Rjlvc26UWuxDegrALrp4323
1TKKO7fTA74X8Dtby6lF1/zoPyFOfZ1371/N9B5RyhBqQFzUg6y+32fowb6LHO6d
L+uN8FHHKP/88Z3mf7Lo5OB/9VF4jWSC0zbxzRgy5rWstKN92QwJ/D732Upm59Ly
SW0JL96/MOkMJls1utc1n+HeyucgCVINzhngBQ4liDRSwbe7B1G0uVNZ3cHGpyBv
uSMmtBRivQiuOC0Y4C48xWREwK2DE5E9nd9Ec2trJh/IXHaJ/67fWt/fysChNW5W
6Hhj40hQASbtPx1GR5AunSx1yMdV5hLzQkT5VGAXU8zlPG8QZDVmdd3VrJ+xN3ra
aG1W4vSDrAdWGYYZxRU07aBtK2lmY3s+kbQUBNrShludMLzJY0ttL3t/JH9icroo
KUcyDLLCVv/AP9M+f8LZc41Ar3YrejU6y/b/Hs+hJGSjmQhrz9PjX42iHjZlhGm2
EpORcKUu6Cxrkhr+LkjlYhKzChZrnBlX1yNVrkf58AxdoJfWMos9sAPOC4unTvqW
ZPnYr4Q256+H6HmkVbiYauwqf9HSSKbCpH/zkrYAqHxRJ0mWISrjV/C+1xabrYEA
aMytLT3d0GpP7rAUBy9YzPHQejyqoeKISAcB7KnTFmtef/tFCvajkfyQbat5DlqH
MsVa8LgoVyNcgaXrb2WMJy1ROK5/S6qlERyuE0M0s+XDI12GPA0mL6fY3a8RzHFa
nEfC4s1msFKRz4Og4YCv4z7gAZrPxv1fE6xenr5qSjlAVkD6ZQ8idluLfK/joNvO
NeNLw858EDMh5L2UyBT5P157AqhjBeSZQiaOJ3US9MU4goMnXkrUyJH+iDfPGrmZ
b2bY4DoSd1HefyWhYkKO1T9mvzqQuZ2zTo7B4VcQ507N+JvK/OV6CkrcY18eZH8A
M2Ot+7qGxex+t8ZrOFXrbGPTFWUKb/ZkKapDaGttNH34ljZcSMpj3DZEEEudaZPz
MBxpw5QLS8qFbtfwYxFdyLn1l2/ku6QIJibe/V9rkb8w7wTsW20pVGewltZVjSkv
me1lGa4+RIgoUlA7KpfwaTVVbFMqSTtwRb8e5HtowIssvYOJkRDdIOWovNghp4Te
fbvBfVMI5L338wHLqqEFkbfhgTAOD3yA7wcxIB1s50toCeMoXK6oyNl5apomQhrd
JBEAm0ywaIeEiPUK1wytZOGATMIKefIZzxpb53ZGIAYQSTqGI02tfn8w68JBKy0l
5k7wsK4J4qSQNSymjUGygImEGdQ5JdIgKE3bCoi5FVuGQVfqHKrz2NwysJB10+H4
kvC+338iKFL3tVs4l1k5uAlh1ZMYkMjArcfeUgTJURWAgLFE7+Bhoa6tuM3vJYUk
hWEd/7527n0kLSCDC3d4KxExqjo4Zt3OuUzQmKo2b8uoNERcxGaW482UqGBcsy9B
wYRQlX0bRsB35bVr7nsyGAHLC6hLigal+jzT2EtdUipkplUMuByhCnvhx/ihnM+m
zjz2lUifVS0Ey39pDPMixLwEu7pAtou1U+bijXyQNH3FRYwn3j6F8HNqXAZSzJGn
uWGdn4HXu1veTXprru8llKw+GM3PFK+5DTQniWWogw7xr9fZiqYbwyx0b6tw8KhN
HPVjl4dVlC1qKhllyIAfY4qXJ85VjHQRZ/yyebN3sXndv6ddzfgZTTrBqvCnune0
EoxIeTClxctvZM3EGq+HX1TcER6Ji28OCjcvHjT5cTWRUYnpvj6Ivv9qkP7HjcsW
xDrvrnfiDabZHW349K+/PldtIBnI3TtzYF+dWNZ7wrbVmS7gjKrTMGwg0F55NHU1
UiFdc98RzkGq7TdhoPiNNi9PmETpd4s85kbstArEY6hMS2aLmhO28f7BDKE05H+0
IT5PqYIYUGKDVMrJVCDRdmruEPhgSEfRAalZmWNRs8iqgCJi9lKOM9ob4AVafZ5U
bJHMNBljcMGtJcxCp6HwGIIljReMKXnqpxHm+bVMxoFfz17ykO9TarZMGNIiwk8c
H/vJfxF4e0i/vV4lH9FYATcxsIkp4GoSWzbUXpUjLDXISuUyI6OF/j9PYrLM4VBI
kr5SyWvjNazu4wPL7K8XPybaRuH7t6/tNZDabpQmZq48Pb7yXIUftxrO6ITn2Jpy
hXMyRBf7D1LXzzpoBHayFDlKQHbLFk1szauDjDiClbilxExZk5bVEXcIjQP5M2IX
eIlsyeMbdJIjNPsyC+Jk743bOCyug34xSaKdbCODVIHCHMcQHG3r/QGlhGEBIRWy
UGjtnluHnOYyp2QadfXoriigqcm+LZ5fOfix/pCd6413O7cyB4iZcyrp44Z3RjS9
5AiiYbyl2oeB41D0XIPgYA+aZgxrCWY+XhW3xsJQlK+dNiI+HeV74DzUwAeuA7B4
wYk8xmH6fKVBWkZ3zY7Ka45kTBEL46YbfkkpC1+HATYpuD8sZf7QuPKS/D2GpF5W
gSSRBPKNSKBphwgFlXQxY93MtXtBicPPuOpytm5CqhsnhPNLbL0AO98O6FM9XFaR
nQHOvmN9mEvpXyGeC6M7Rmdo+EZxkSvPb/jV+UdOsFa7VHSIt30cPEhHEEZoIIrD
oLTL2i/c9OnuwZRHQxClNT6JutvvLED2/RNHyhau412lwo4GdsPpmTyPTr/tuRtB
+Zrb902hDW1OKSpbJUaUMQ08yGRpelFL8zjNE7OsM8fv/KROD5WbF4RAVXPUvQcC
/NihUHrNQbSRzvGUnUmU3sK9CWBd0K7GRkW8Pi0G77U73hu/S2CCDqropyPHVRSy
pGm6tCzebtz9SQ1TZshec+yMMlV1WJnkUKQcXUJnnsmRPDaMk8RAbAL0g4k0HiSZ
6eVUhVNCmYBUJjV+SVOmzmaDy9Z7J4IvuUlgA2ccW7+P6/ZrgcODXP9Bdj/RGJHL
epdbnrTUVCg6ZIW1tPK9HY3UdVXQfKleH/mJWDW3DFj+X0PB+WoLe5fl+bg9vcHK
kNtQT1P2whvMYLZxWRJ81R0SswkqvwZs01pPDVSdILyGBSd/yZHjamd3RRP084gg
x4SO8Eu4qpEQpgK+gMlVl+AE+7rNIPYEWqpvJrxlPI4F7S8Topw+JwcrR9EWvQuP
g2UnL7hHQ4LDa0XUDlsPo8NVXROORixDHIzWvcQYPVMNuxJ7WzVoAoiN6fceDeIu
Wu2e7JzcnzRGq63ogPapr5VgZhiroR8NAkNsdzHeU589DiOmZdMDON12M3kngBN4
dYQbLayelME2q1bQVzq8zT7EJJaQJHwILpLoqrZGXQ65olUCKl9Vd3x36swxzSSt
/gMOJu9Ft3K2nP9x5TTx/pouOlKtqPl5PuKjC1ftGJcZUqWcpE4x/rpPk5NrmSQJ
iTyBIy58YnDIkaEG1+7a6LEmazbp7Uod4/RcBZ0S5OFFaHICrwkEno10LFbbsctQ
lLeHMxdz9hKlOKvWIXUbaLYs7mVt2PvkmeDUGqxD3D5fj8TfDAqMHL7l4nfSghiX
DybJPcSuesqXwoDFXUt5q02pLDaeotQ+lSsvTWMPqwUTZ+zRy8zrB4nkohcWt8Hh
0mWNSJ0ROD9+d/ilLDR9GXAyh6LF45NS/kc8qEIET5vlsGepNE4nm2DvOY3sh11D
JJZCpqDSV9+WPefuS4iN/6bZvKtqka1YVbBuGzM3CWXtigmj2WbT8TRNDoIbE587
OpfNWsy0m9WJtdSgMscPDMxdxnVKyLV7efYkDLRKvQxOVRfdlHj6CC8+/Fmf1eXo
4V5oJVesOSnZ9GTBz8Kuy+qRa8K8Ki8es/iBrfV9b+tYtVYEGSAecIEKbMk1Rzyo
Pycjkc7lzRW/TDcx0Rw5xqJGhxgSmWlT4P0Ao2RSBkWo3QUtQHOHuyWlHN9klsYU
JzJ+XevUwiWEe5sWVAHY8hC2Yp5uhMJVQD4DSmt4B9NREPgoJpXuUD9O6MSZnGJ+
ycxxN84fEx6YEjck1wYgxQBoNl6UH77059CS/49iPfSMkJVnvBa5yOzyQ2WKI4ao
AuW5lhaTu53vZqc77Yefe3MqjYpyEJikLa6O9AJrkZl2vvhJQHoKTxlPhjMrPdiH
xHWAj12hvRnuZD+A6UhK7P4HUjYTMeRWlKi1oj96AqJ5lAt2tl0cKOV0XhxTPH2w
iwyeWyofJfwL1yDp5qFE5NaDOJt7ky597w4EI7QsGILXPX0f5Kd92MwCDV3y+ncr
EKHXPt8gLBSeXG/ADacS7ZLlybnwDBxCenSQtZh2BhRCnyxkslwTISlDnsxccoyx
jDtbeX4TnL+CLWdVNaucv4fh/rtKQF73J15ZlzScsU6MBxaRtQDzYVEvvE1R/3FJ
LyvMpZ9z2xtrv2njLvX/r+VA54h4TPQFVTctMaPYB6E+h6lgGYgjL/0tBtN1uy6m
VKu51wIUwuynnwHwo8dnc49vKwjDIZm8p1wVP3yF0ZU+JtRScJ0viyxRQAtFrz+M
xHnuH2f3pIPicbX8gfz5ZyuE1ddtr9ksyQ5cOdLaPfIbvjY9Y8kPCkxXNJs/L+oN
ybhGi6kXdd7RZl53//DYsRt3mnA/Sc4MwfVOCuN5RSB9opDCZAe2clsm064A5yFP
LN1pmzeT0eXOk5AgzUxsd4fN2sjdt5dFeH+pL0qAxq6IQ8wm4YX0TfIc8dVobcmv
l6RxBkboog943pP11/cLQR3DNs3nHMpAqhXp76KoA6I/L+t9rfYweQcvSRlTHae/
iVT0G+Uku4TacnTEeL8GvT3x48hOfwleAgncZcI08Iie1FQFdEbUAZ5CRYIfbTEO
7yVi49z+uTNqPMjiOta/dy6cECenGFzWn0d+rPPhH75a3kLs7QeL8/w9t4vbDQrr
xeCNYrfYJFlWXbEqwDcfrGWwhykhJsC3SrgyTGz6BOsS2rZsyIYuFVnQJuw6+KSw
uDX40hrU+AMukqe8nfnBuRkk4X1qMs9Ma9Ow9yl72ODBB71nkglN2SjuYQIP1j9J
c2kjJHWx9GCp8p5sLSU8RMWdOI1NyrGWTPFOB0wIZ3qeyfDidZZuCNzzSe0F0Blr
Ld8tGn91JgURYC5ypR8wcBKdwE8BMXS7lbBMSi0w3Fc0BG65CXMgzxtgBSd9khGd
jbOw2UPoKwyGlKZOdzd33BVH2uV4ZsH67IBabAPTS2mpA1n9bjypXfgKk4Lh/aCc
+remmjndH3uwRP11KDot4B73k+g0T2Q/wJQCBIRwbm0uVdhibwFcS5dlZeOsl/MZ
gK9B9KZ/xvZkW2ZKVuCzOSiF7+HVrnqimYiZxJ4svWUe7I1HrjS6JGaTxdHg2aOG
TWQe+YadTxp8ddGj8M3I10H/h7QtlfacHgxa938SB9T1Y8K3FZ4u9y++y1894A1O
idRke8R7U4FTuGL7W0p26i1d5vY4T34X+gqoxBpwF1GDsO0g93qa1EIuddWlRPrw
rko3RYI6KOscN7MTStzoHneSYvSiQ3QrCrjRwm+UGcvWAlF7qytqmBdEpL81ztlT
jp3JTqQwHtWFEfMd4DRk++N7el6qLgBozjR3o3+DG0pwD5ur/bHy6ev+AGhSAnWh
52NcEwxJxgPhUU2kjqv5Jx8AKB1foLR9ETU9i2KTmAxNr0O1lCvUX4oW8nw1TOuz
hc4SEDd4eeghn6nsXT7EqsTec7inbbXedylmpzfH0kEd3xLMxZSbZjVwgAvWX6Yl
NgtrPWdFJOD4dwyVG8MwnLe9h/yTcJUX2nrg3ZO2JZksJwWrIujdEH9tllDElBmF
H4USmgU0B7tuB2BI665XTkJTtcl6NgjciUfKh7nQWdrF6ThP0JRuj5yWTYAIQzuM
8Wsgd51tQMOqmwGWuciS0kfK+rATMNnOK5uUdU0j4JPZfQkHrX4/SBqCvKdyRbxK
9X9gSerrpUfCSXeHyiZs1FhuCZRvISwLvcvn3fGlA6Ji2RPVcgM4qMGdgQysPzWz
BfIlX4X1jP+TsiMzgLngv7FTFreHmZGh6e3AWP0bCoYPOQU/+/zsUbcqY9lXFW8H
lTniIrg2Xt+dKJUedRF8CxfiuPJ96698KE5vUj4H0KLUBj5YMUHJkiSr6r/d9h+x
UfgQNA3WWqYUfJkUegciW0dDRMirNl6tUQDhYP+Y1kIB2iIxWx+eNTNoxUzbd+hP
fMJZ8+K8lDsq6gXhY4+k6Wfrbv42XAhRpcDtk3/xBGGGNc3s+6tyy39cDDy8wrwW
y8XeoZFVpkr3azfd7gPAvZMGa+a1nut9DrpXGCSkdCTMT14Y3J+4E6MFf//D5Tt+
o+s6JmoGOcTUsuW+rzp3uvcY3ej9dcoCPF6A68PW+AiaDdi+Gc3uu1nU5p4tlcTx
cUrwYm3iSXopSP4gE1/KeHfE+r3zbVgLStXOEz7tnnqOLgoqJKnXZttHB3vE2fXA
IP5FiwZMf4wgoblFyo5Xd9quxQoGJ+x2tQ0+dCn7Zz+Zxx3aqVyqxPyPaERopiX9
HQNcLDeYf8RR9aufFeIhW+JsBQRq7EbLqOv+RTP/s/QjQME9USzg8EoIzrYQuoFj
vkFiz4/mrlOX1ELXbBV2kIIOhP+Jx/Z5mDTHmdmJq/j+EMYCfsZUvJ5tNwmuWo0O
tkgJZd96JcuRTaKyYdZVRh1olH63eWVQ//sM/Y8JowQKr4gqQqKQS8UKqQQycMWC
dBcgSx/lk2rl+Gdp8cSZS7bLUx2jcvUKf9ifMsBEWrCRaBv73Zt6MgJTZeAkjkhy
1+pUrIYyNE3CNGlCWc3J2oJjhBK56e7yp52605LEB1TBV+mSIAURGACl03/waQYD
9uEHrv0qur9SU9iT4sWZwy0VXOJO5gW3ySlj/mraQ+hC9Dzsp8BULy2ErkmuYOsT
BfF6MG8n4Rp1TL7dATnyLLq1WeLY1SRmOXBuTwuUET7LJKTkWh1QhvrYkT0M6xZQ
v8G9wRjIeb/2neDcuQV50nNUcyUVUa95bynb/CyGVgVtW+WW/3c7RY31HpacDGEQ
do4Fk8kmHkiXwJfev79QMLmCNFTtkPPw2+EoL/Hiq9imoUGSxG891Aewf5dhIb4r
EE9w4f6cNgcb8MMeY25lxJ+M0azHV8vfbNNLA7BTf03G5J0ReKZglDW79OuHz7CO
7jex7rDry7ZARMMbFCsHUOXLduqMECCPXFnClPEoADQrHLibFZaYQQZ1xb7atr4F
zFW18NTw0DyFTBx6x4P5QSB0ER55HtPxcouXJyxyzLBLhGxRIGOT3BZERjWmlNzK
oGNshZc7GY9yIEyobw/IxBvAcheGtu/9VF9kN+E631WQXlPG88C+7XJ3gkQ7aW1e
4RvDJtofCQg90Pbtr8zsYy4fpuXKaxOAAkUSCW+lJYczGmefOWef2vuX0KzHlYNQ
GgIQsFVib3TEzs4uCa1Qc2gC7Cq0PvLqau7yYzqg3TavzZVtV85vpLIH+iVH2c4H
FUs/InO/d7a4oBM6lBiLGKQpQy4m0Hke2svZtGOZcUtvFxQeeS0KpEEnVT4FtAPG
IpZ/LC4a/FxE8WUDveGrYfArKXo8rxYADieBlMM65A5Xp2CgWqdWG456UB+XhBXL
9fOh0aOGtITOweknCLcsQ6PltAr4L8d01q+CP6cKRDkDcpjukSrxdj69I3pfo6ii
0DqEv7O0WnJLf1IpH/2ZYu1a3ZRk724J6kFJaJoF5RT96WM0nDZbJ1md6yniKYd1
E4I2tdX/MA0hCbtjD34JAd4VgbNEoCEjqO8GI/7iK4zPuoZirphIf8w22SdkHUqc
gba5jiHH9lOYD1xRi3qw4GTK3UchDgNxP9rBT28h1nCoNmZH5FiP2qm72ZMLXzZy
LPDMrj4+EpwD8evm6AT95N4jvvL4sOsldLSBF3MK7hP4besANPO+fpo/TzuGr0uL
+bnHJlwJ+xOffNXPdtL9iUYKhf4uto1eN6cwtirqkXEQLFl9b21olxAnPgqwCWK4
6A32LC+NWKFILzLmnVgIUWIxqgoCmlo+2yARXfzfktpWoS3K6152UDXejmPoqYIJ
IA/GX+z+KGJ9/FpAIznP4Pi7tGQs+TpBROC0TrGUky5SQ+nESVsD/KIYIKWyePkz
W25PX7pNbJeHLBEqpYQ7hhsP+69yqwjz8bnPsXq03FgeADVFhk9orkx4AOHqYIJT
aGAlVCDHe06WIrHGY2btDDUrpflfFkppoQAWWqa8RssTwFHoD1k+setZi0uVP3sw
xSu+CnXljNUKtuwxoNMiV7HRnP5oWT8g74KIwnTnp8vJStp9JfqwryRehV2nMH+K
MGdatQxNrPv94UHAJstau3wl6P3C4McNFDMvdQBpT6V6AztlUqSlCJR0TjsFvwKP
ZHYjIJYQrGWTi9RqJSpp/zsM4GFv+igcdTnXRXt3ZIBd7yIrfi8nb3+d33gZ4ciJ
Fx+I77yKpMeLP8OgTPvW0b0wY1KIwhlx9PTRA3vCSPNpE6bS3EONIzIjLIliJR7V
sXnJiCI0LIlFXHTBo3skSmJLtHwiODra2k1LIxqN1jrQPqy7TgJ1IL4QcvAGOHYQ
dpZb5oxCa+SpgtC2pQt8mUBaal8m7RnWEZitEgAAf06AiMNa6J+z8xTPJ6rV/9bU
M8KiBIEOMF4UmBQrltQBHinkIHdv8ufq/9tQompLPb9ASTqRLDnIniY5mJRC0pZ1
Lk6ORMd8i8PwY5ViHHuVSEvrbqX7VA+eo126NLH0EO7L1zqyhDhwHEu/NxjR9dJ1
xtIvh8M0gbHZ3B/D84carTW+ZVuuqOakkuqvmqJuKwCF7t6zXlq2Kehn8n7WcFmi
psozIt2/Cd1Seisd8jCTgVJoNKXEmxpW3aIk+RNajaxjJzDCmoEHhp4b3cpZrHg7
REZP+iWuCKCkl89Cq3kGuY4dyauw2nnqDep5faMs3QHkIb60/deUJKd/QBOr2qEA
nN8fbNlPJyF7vGW7T4diTiYQkSQjqFQPsbx7o6VIBc78w2ZafXojSEIjLP8ulBuH
p2L5vYDln69i4vcXKaOfBEz7HUvYzvkB8S1e5l7LoZRskAA2JOUe9pZ1uhkJmZ33
LuwLIMSqF3ApgVsvK6lqF+u967+m6oFqe0jq2F7YBEtaTZgv9BYjTMGT8ob80FKv
68DTxhhjmd7tnPGNADqJpeOqQ9EVEI6DN0QiqPvQp2oapoP7lH6t2CpBVtzUPrOZ
BS9ctznvUdJefmbarOb+TtleQdELk+hqtHzFlNcb45IC2Yg9jqbT8QIxVyc0Pfj5
+DkyDBgsuWD3kakJ9aLjXvMjMdx15HzJGXtDVUk/EmyVn2h/vGHMQMHFXqnPMpO9
9J5goSM7Ue71m1GUOQ+373fZ8pm9F3ofEPtFLeapIJOY0SMutmP/nn0Tr7KR4qNE
sHy3UF+AD8LWy05cymSlDImbWGixFi43ewzK8ZmeveuPYpw9JOV0MPHFDgcIG8Jm
lbvy3ARP8NE+6B3u5i0iKGGTtOoapPmnZ+2fNsiONgPgK5HkOObu0Mb5ZIMwl+Fh
8gjv39CLV7Y0T38CI/uQVlR+zcgmV/7LNWoNF9SbYjwHRRZgZXquURwz+LPWYVwB
GMRPHMXoz1u16ey3AyAMzakIjlyaoPPe8XpLsijBnOYlRKV0LLEmlkC1G8IC1tGQ
Bfhoho5lDbOKix8hlTYtg9FOeJTR6ZBGpnEtkZI9DXR6F9T+Gui3Lj+DFPuypaG/
hCHXp37wY52C2dcjsK18hZtz3D+DEUGACRN6fuiX5kAbac5C3OQcKFEKRrGA1xA+
92Ft5QAnpmm+ad9YA1kLFeOaTFJaIOvlAJ7r+T8z2RdMfTXsKsjPRy0Rlqm2Xj9M
p4TzbgmReair+HivrJ4Yq7lys68hXxtdZYpQg0+ofNNCckeP8/fStCNQCoW5SVPw
CWDTVsZgYJQCtvA1CoxgvKgTEHLN/xmK4lOSKjztr4/j3lbC2Fp+UuZ1W+oSe2kH
fquEYhS7UXx+M2PMy68pYyIxR76CkRZnMdIwTluG08ufMv5kzZnDRymSQQ9LE6+n
TaQAde63xrT6R32XhP0tiDI6v37mfaWypmOiBjiggavCm1yw2EEd0ys+StjD8dRC
pQZeN3XR+w0yMzZekDkWFKVyPiBZmJPof2LtLQaoj3X7h5ZEnUciY349QvjhBvz1
7p7bhD9sdFOoon9GXufg/UlAARisPAg54PsTEzK0GdA7HNJ0X12B3+wdS6wREbgR
L7tYUde9uaukY0OuWlpJRjF2psH5adjRLWLj6fHPZJmJSo5n7TQXjJhbv3Q1Caow
ZcKbWSJbkPBIrsL/pT+IuPKlWi58OEChxMzHAh9DZNedsP9KnlzkMOu9z8Wp9/dk
JMvKWuyqTVSxhNqOqdc+1m4Sr79FA9A17CUPofH+j8uw4koklmQ082IOHK61v9tn
G2fVZ4TJkyd0MlV7P30KxMBgwAMTry47W+yt+OTyc23ba0IIR9AXccW/N7oiPScw
997bGvyNBI4bFB6e97fOuTzizFLsilajRb0FQ+6nxuCjG8d5Z5yUOqdy2TFS+VNL
ILINIZq+9MU9nPixLM+dmEY4AHT/WHyrntdqEteCYxJ2AfMLtMYlydJ2RJAEVlO5
iDV920k5MXhle7ner3Ikv8jBoPk4HXdZ2y44ZzVy/YlKNcNFrdd/ZlKGrU575pgV
c78SaaHSrZItMrq4Bff/HA0fIOOH1dek8TaKYBQYqvS5lYrjTg1+wrLPiOwVXszV
6nPYhNb4pEnhZ9/bF2FRIZLeDDAaznp1uWC1xFqy4dThd7aBsOb3wTlqmo+2QV6d
h0KY55s6vDcHAXoy3iFT9OdQVovHWx9YLoYuGB8FlAfrcmk3ml7TGFSeE/Tk0O2v
XI1eLicDMi4XGTmaa28IVzMre2gCHP0A9msnDwWdWprFIuf5AHEj1vZjUI1NlECe
aGhaK1XEw+DPm/iR3J1DZDfrJO4bSaCTzL2CAcC9lW08Wl79QcdkZj8MYjz0r2Mw
81O8VUTcgGtnYp5CT78ioZC1GZy8RDhczRSbNP8wIEwLVYcTheJiCeyUmrYC85v5
9hvS/Go5xpOXGBPlpEMZaUZWoQtzueCfwsuI/i/koku2r/JpAch9Uc5FRP3ZS5aw
2V1TJF94+hwHle6Pbdo9Y/Kj9wLTFgwufQU4+1Df8QGrL7UtKrXfHnPTYUlNZjqE
a3HT62M+9FcbmK+LH6JhweXwph5JSMCYr/3BzQIX6Drta/QecLf1RS1Xs++brNyt
/kxpnb+BRC1z3hU/sg8F5MB+nMOYDaxMNjRoh9WyQb1fhoaKPSaTgl7Rimb40x9e
s1uw1Ggi46i+uIYX26QsEmJm8rgKYGwDsM8vJKJamgU31GvMqkvWsUEtdije6AB9
6SZLqqybOjTT0YrGJsVl+jSHxM//y9HfaPy2JQry8zqFQfRpAQ1/n6YHCkuPcR9P
1WDqqdnkEuMP5VMqMtDW5WxlHKLDBVpp9dRWT1cQz7vrWAvw9/juXsKZNgD1au2/
u/Ddste5WeGdk9bglN1fNbASe9XBKjkH019Va+nmsqTveTQfuEV1Umx2Vb8fnhtW
BL4fif9Y+IFapl3gCxmCdrira8y5Kj4EFdCiXe/pDnSuBtEt43eddzvKfWsxNUO7
j/3wTLITMP2H0p9qefQTEpSDexWNiMHfST16jSxPzYb1FvhFUEF9LxWAqbRHEDsF
ju6w0frw2nslXi0rVVeLh2W5Cb44LqY8hCefdXofwkfAWv0Fb+bMc6etVS54ZlAn
0QNkw6ns2hi/ZHkCOfLFmS107c+kOnayOctN2S0DyUgpsKckskzX1vM3g+DDf+3v
aINFDZvPBVpGwH4o4jNeUVTS9PdI/51vi93jIyTT5oAIMolMyV9BZZlzA3b+HtEW
uaTyEfQvvgcX1IqhQifzd2FwISUIzCWkO0xCRLYB0+TJz/u1Bkfy3oqZaPRro+YL
SxGOtB9smPssfuqBLP8pQNqLxqX5BSM8OgH3nznJ4n2VNkW6hhvYOXr3t4FTZvxv
xrYiOoodK9DBYCO3tzzuswiZo2z67QOoVUq7NwylOoU8CMevk3iUB0ta8xu9rcuc
nHNgSlwnDNJ9aoNtjxEf8ayEMnzfzqTVfnQW/cBuVi47yYDfGBBmKhOz/060eRgD
aMCH8HO9IKOzft86g5wMNaeudM/T4aKLniUnNdNsDGRjfYiz6Cz55X12RGk1Jbgl
vR+UH9+kjoWwQjk7ZchONUCpYvJ4NI2EjsXL72sqMBmyY8ItQj29DqPcuTarxyPU
dUB1/TsYMox42iV69OztErTeRNhuw64TVTqr5mxKVHnTpaAFpht6S28Uk/a0H1b9
j21f7ppuogGNBtotuBDCvGLiSFDqfU2leuRcwI8JDaBcaUKoTkZ3tvrpMGLu7Z+u
PFHgg7TWqwPI+4S/ENWvo+FFNSrhdsFRBIBcQ6TWmEH8PRR9SsddVEDAE6w7rR8/
OlrA/ALVORb/T8CRzHVNwUgqqPvBnxupSqHWY4IZgxHVHUPcA7aEhuITK/r+38zT
fW7AbuclnPYvZ/3Ir+ur9NGYXiCk5UvM4NUP1z+u4wvKwfrlqQvVI/4UYYHU7qTc
SqiHbbyO2Mvx19i7FHTQID+8QFxberAVRg7XXW3Xz71Vu4kKa5cxhsavv84RQ/VU
8+G0yWdDrJV0vxPvwr6pjGdg7zNrxw+mpe8QoPXRAcpoFEp5mJTLsWpjx6ZvLThq
a2fHimxGIyNJyH7WQTragHERW1Q1JZQ4Vva3CGTdwAWswaoN6AbbDiRG23ZtNSAD
TsVsPkUBHn90uA/wc4TFS2qIol/D0EZwHfh/1nHr7VM7B3Zi+L1WFbkf/YwixRQz
TPpYrthe5Iu6xcjh/Jv8gruX4nqPsRUBNaEhlr3hoHBwiSYh1gakXZWcIBUGsowN
bPEPIXvvcCRqmL2TrtZRo8X3/MWsnENzcaxLy3qcb0GkdlXab4noqqhULg2V4B28
/kPME6VUMBqhh0sCWNmnnD1Gz0MmbA29BdGKYOVL6TrO2IljkmLRBVGyYsHB3OsP
R5NfWN6FwbuMRDG99d5MUAcA73cM/B1lkcRtsyWp53HftnScx8cRLxq4+ICda/8C
cO8Zufz2fJYqmfwb1K9vIRmVxl6cBZq/6jsO69i1O15dhvKIvvyDWj/VSdyc3us7
4/X21feqysOVndDzNo6GBBO108cgO+MD/bTKyloV7x11lut5xgPf89erj4CRnl22
0lYAr9K3wxhrbu6aW0q2jqth6VEJ9ua6MvNcuwVmT9oFo8VUF6Lo4NQNJdnrWp+J
edaJPbS0+pgzkIsS0W03rkZeYf9AZn7via1SC2LKM9BjoyMobFcwS16rMdXP+inO
mWt/MT0v3iCvCiLftiCeXaGWtbVXGvtHy/vXRvc5SjEEnk86gDbJrRHFRDx1iaiG
e/2oB0mEqV98aDJ4xBqZyVK+OuagwsYrR99LxQCqrexipAhELKfsRiqaJ9VNECNt
NkdB7SczMtdY3Ap4GhiiKh2komL13zNn/Tpr1ReAFyjVj2vPkPvngiIaFMvCtweO
N6YFp2Z7qK8IdopdBZ+C100I3utO20UFAGrQ+EhjhERXlmQ3dFcQKv1CP67pRJiG
GM8e1Q/D3+Md6KV46p3+kaIEbRxAImf58sE0UvsMxPxOsZJkTCXpJCaeXxy+h1IE
/WJd+MaV244fSj5vg0dSFA0jkfGrZXCHU7fWdHWWbt6L7ZFhxyUTKWAHDK973z96
mMcBLYNsu5O2Obco9Y9puEQ2y7aTVsQDux6etMaUD2btoCqF1x84TfApjoI9wrqX
lpy2r5qB0+GfhspXRP3LkPQIgb3hxn7Zu4kbzFbIKOn+tEw1Nb2NjHGU1I8HVePo
uqOmFBiLJ3TRne/17UpuFexXa1dDSWO08xwWi6nw6b5sC4sZdS2KBj0ftEosPdcS
mx0Co8KRhmkigfYhfqMlT4HFlobiKMyuOfH4PcNJjyuM2iHXdqK4lNvDQrmELUsS
MRxiO4lMXQbJu6DI0sjxgQKMWHfUdHyJhCOMCmvILI9MQEnHo9o25mvpoB6C2WTY
qlJe96OMSan32cB7JPhF2GJmC1dRDNZ3PIwjXKJzjOcQSx4YMMt/D4v3Qbu/VmAO
3lXP0ef1Biwq90noQ60lf1iSituuIxIhEVWM1fAtrSCZfS9E1A8mTrg9jlc0VUz3
JedQJIQqdjTWgGo1ucq3DAY0sIqzCI/+cX1Ogz4bfNlyFBpysCZQ+KbhFYS/akOV
2gR8BUWVF8GIEiEOtX+e6CZ21hZ4a4M0AvIWMyPOeauSNr74V5I0zoAJcoWgJtCd
T7F7zCwux4swaRXwLVj8vhjoQb7+HbYLh6aqjUIWijCC+uY1cdoKDlNCos69z8D3
TR87kLWRr+OHSN2MFS633sthWOw4DnIUaaeFwOUlXONGq+9ERuuVAFNwkeI4v7ND
62x0kHxSB/KaiHp+ZuxZQnD+mGYI08+XgEvu95z+EZnUARfGKW6w9MEMWpd9L/QS
9tv5fE7yx6ASw3KY54YUSvFZ3e7jkPc7J56gb8KWZIzuW2jstYjyp71Xv0kTLwZ2
FdX4iu5nmPsulaNAarLUKX/1IORMQKNMsbpzl8bFt/RKp3029ECTDxFaR7xWiRql
NWtoAeY9xjHofjCNQj7yKTe5I15CoPKfAY7E1KWH129PJHNuKarL3/PJAE0RcLmG
XK71MBcwCPm/We7u+vwkUErYe88ZEbCtsoY3m/2jKLiVPkX+kbfXVeMk9SdTCEK6
jHi8Ze4uLc1Fq1KVe4K3MGWt6mfUgw+bsMNPAeeYcP8p/rZ7LkOR19UE/M2DMuGt
roidaechYWsXK8IYbuQfX1rwdoQjzC//d9ViymkMmQWVjJn1BwDHzdLAsH/9ovlr
0KwXyH9sGnACTFwDWZTB4wSpepPiH61qtZra0mBlcVY62jvcAFLPgkbrg6Jgo189
m0/BE8VL2Kn6naN5RK35qbiFkz2lf1l5fvOe9/k7qdcTiJW6DXiYlGSTuwdfH1Q8
jzbnIvynEmBACr4/SGeSB0Xs6AWhdiOEBPo/DDWq9gZS8kGd84Q3Yl/fUTKOO+fv
mlstRALQ+SfI83KDDodtgAuPTUJIXtK0qj2WIjmeCH+6ifatC7KSyQIRumL0Z77Y
WVwfNwtC0J+Kt7RFyP3CwHD4RHk3NwspHnHhQ1Ieg7zPgWw096da9S2osx4YvubC
eqHKJAwh5Qa6ZKcBjOnsEqlC5KTdGr1KtnqoxLG6uamcar/iWOTTJkX6OeLl8Fw1
vXinoKcVXRp2g5RCnqmW9fsnYGRqXXEXaUOYO/FI/J9LelpgmK6izYmIzDG0/bQI
p/oDRDi9Rai9Pk24yihZ9XA/X6ZINaoq8sZLDbdsFCFe5/aBuHw4lMsrDOhTHWvr
P1tHOhnVTrdXAHVCXCBT8omG0V20QcfTA8fuxujA7UoPMEN2+hpiOPL8DETwnCKh
cTOPSEGAuJfMQiO1dfJVnPVLBV5rg9Ad+/bMp21U3hoyeAuX07IZMqanc5i+uT/x
qAXfhtKv4+l7/p2lsKSVbPj/942AOBlpLmB4Ld2uBXdtHNLDEY0erIJXlTG8nbz1
DlgB0MrjPpyR4BospFi8KasfRnWjxY6inDf7xvR3UAArnc44G+eb198an83mXGqs
TEfzDsqYIq+Fx+QQbUR3CyZYQDLP92aVQIrscU/fOZLgxn9CGHcJnVhHh8J3Ob+F
m0rbfhqkmSH39bwNAQlQrT5nPDLKIKGScuuOhDvy+VI7fGAWlWqqGUU+lHeSrqxz
rlWzOneWkcyzQ4paQ6yRk55iwuf+IM1bp7J/HgXuLA8ARMKKCdNAjgXMui06bE4A
W1bnF310hM3wo+lgiqwUn5YcZ7DM1cymjWKvMVWb2giD66xRozNWH+fXrydF3yBw
tlTm9JuyKnXmLhRnmudkiZLKPicLjY5H6OLqOf09TXBcxS19hSwpNBUryMUVGh9b
fomv3dRazpoHozt5jcMW3NUrchfYLz5ULooVABEXc7RL3DKliigmbCxkcpF5sL/c
+syoeMd8It/QkceIA6CWPzggCqD4SyCkTEkXM4sprhlXRY19MFa/FV7Griaz5ilQ
7QtHxEgW4s9na8cZoK7H7YEy8+k5KP+rDP1ePXzpx6DVbRGz0dHiaOD6O7K/SGF/
7m1pVGs61rw6aYKgVSVA+DE2Q9/qwORk/YDyvEW74gl2a4R7YpOVxinuEkOBm5Lh
bzzoRY9RMbGhnu90qoowIKbB4Q8D5kCp7Jgd+ip48JIBeWWOuNs2ho0AIqhlTqel
r+gb96zfLLFksLdy1IXg+547e9aT1m9dBHijoL0feT83EVJV/U47mdJRuu9mj2Jd
NYFBMlRaP1l+6pXwEJCzmaT9v1kzvK5ZfoYNoWA+XV1IwOWxR2n2PU36Sh46O1Z9
VdVXo/hI2PNG1oSu9h8x5d59Ypb97Yj6hr124o8s59MqnraUaJsgijlDxpuQlQaz
Iek7y4pvubu5qy6W1XQaK5iHX7QLbY7Tsdm8UlzyJJw6ghsrQoLIdhdXByPIFqtB
jsKQUAy4BTVYzaDmGpldx5zSnNANKsI9oR0LOJmCZUNs9hfh83YHqQIwZlYtWS3t
T2xTc5ODdFHUpJudrLTgXsT6kQ9w/J5F36kq4AMLiJPPkxf5L2MKPoR4zjgihBv8
YiNWgjYZ3sPEINujMyIItp+ibsIXnf/JzSizki8BfMygaVs4UJqZPz/OWH5ISkn+
KUzRt6YR6AseB78GK3d0o9wnovo2945/GdpnvjchHrJ8KOMoDV1BaW74SaYknIKY
pzZxRvkVnuywuFCFKY1nlupT3luEeYmfTa/ATnanVNhd8bEheRYzIuanMN5hocGK
WiEN1OKDff658IyrTIHq3Vz7G6tO07gLNTrrwjrNGbCa/HKctC3g78aAM/2/WmPf
EEZGWrdWNBcH2e3JUlW6ldmUlTuyp8rlmTblN1mjtoR1q1lfEqgQiK0r3t4dAcSg
C6zndq9Ad18c6w0nQSvcTPYH0pZL9+ZcJnsVgph6qIWnH7XIqL4oRQe2X3r2Vc14
m5CVoFr+qqHHmGRGn9/3yj9jiXYicp/9kFXf430c+ibJ+zFVa5x26drGXBMoImhE
liJopna73Kl5snxDFcyZGJSNq/X7VRV20x3ERsCktLedOu2bRzLbGWkBwXOr4T6e
a/GyzRaEOnoQDer0pTd0Id6OeEguv2e+C+4dSgTVINQFgO2pEdUXDZrDYqqFvlPs
a7DsW/oWV3wJPGFg2RIbGWJd2kXO3E2vxYZoZ7B/l8fRCzI79NjcaDYUfsPDVYLF
+NtnJ5UN2SQnuMOWP/7tjtoKwoH91ZOELULM2hoNvfUhBB7ySiP9h0KJULa4gb8z
XEp2drdQu9SQ9/fvnoCpBlTDzGp8SOK4RXXdyNfFxYBf5uDIb7iKoSEkvgwggiLd
8bxH7mEiy97hzbV3g6dvrQu5icT/K2rDulc558d4ZWkSq6kXa1VH6mtvM/ilRt2r
292pw0QRaaWIsh5jwOprpxrmc0zieDNkaWO0prx9Ih21VU5omzneQI4a0G4R57qm
UnDbe1ns/eApSflGpN/Mo9XWZUlq/6n4Rc4FVBs6LL34GfSpz2IFHyGubiPPRnvp
gqcgryLrZmx5ocrDOLv7oYe1LTWRuX5/ayU6EMtJHdSZDfhXzXRD5FK1QBm0NwxH
TAHgsnTi0zgLEjrv/zAOu2mlm1CvrCJF56htp3k/pG2tyFVgylW+f9yMUQ2r3X7a
zzqglNOhT7P5B+TXNSPqxF4RFHDfWeZ6rZZxXl5rwxC3CW1QN1aELFesi3eWYXzc
hrjAyd000KFHDLJ1ZWjxi/bNhwfeuBY07LEWPMjZ83/idFLc2lrXKbaWjg3amXd/
zBHX6NfYzQiGU/K76MF+MwJQ2Z5KreNlmq/16RJKQp1KanUO6UXw0C5VPDhQcKAj
synNsNeT6VLQZkluYt/eigvh25SQTbATzE5WpJpYMA1bKnu5h52C+0TvL1puE2k7
/RpJ4zu+uPyUanPJivepywq6tmwGcBmeoLI9WCzrSZ43D2LBEOpDwxLdXkjPMJls
/cWQdjUWVui/C6EfN4tBzogUhWv/dgcryNW2N6iP3jpa2L3Ja04aYqmwwwYoPqoS
glCDw330fGJnDzyKeMjWGb3D3bH2nmNL8EtNf6sXPDUro16cr4nlnqNgVsLG0BeY
Y/I8J0AaJQRLg6BgV/qPemJXNf4+W/YPClj5G7bvwQaEKUNYjZawnJGCdWNFxcxQ
e8u9wd9BneR0KXxbPrgMys++yuGs9yMC7GE+AjfEG5t9jlIcHUCBJCkV4zar7UYi
mgvoPTUtuIwlotr+6TYztYo+RE9JzJ7W3aETvl4TG1n+ZaLyn+3A51qCBN3bezNy
G+XxjMWo5tcjQGRZXnd+IQ6Rr+sf408chqX3vcq2QGUtrcSugtEpzS5tu1H2ZWyA
I1NDaQziHg96vZiY+M0KlHfJh7kaRXZu3ZS8+Yoh4B+BqJXZGoDI5/Rq0+lLsgC4
P4BoKwabAyhHJQVy+CAM+2ivnBwsntRz27X44ZGrVOzOWqJVXIsV/KfTwGlPWTCY
6NtbE5wOwJof+FcCMBTSyWKa9qjvdp9fzFrHrjna6xTIneNn+Sj+YyFU2GtPldkq
FJBHP7fiJM4TTMRtZR3bZl4HfT988d3glAJxiPtQB4F65tocWoAyZ99UcRsdFqNE
0KKuxI5EUwMCd25pXtFCg2HUX6HQE4/+5v1XKTw7a4+JK2SNj2vGyS6qUrNo3fwz
TARj+IGVel8bFGxp93RfTNzXz9wVzAK7zIBtymdFBtj4y4uAKO3aP0VlohgNk0Rs
QoMf5IyFVOZxWxDhPJDO8MoY6rFyQSFeKD+7MWE+bbcOplBpzbRg5iJwknzIZDTK
HhXwTtNBId11TQXy4SS5o1jAyvOc6YjEIr2pUJV4VfTkltC0BEmCHBukKYeUmNrb
fcoN+rrXmW4TFIXZHoueCmIOr9vQVSbhbN2URGAsa1YMxuhmo8UWeTuvhk6sCuRT
R5lvu9DGHMx5vQ48LqJbq8uWIGIokZsKDmWN2NDlchgwfJ3ByYA1oZEwBvm+aL39
YgLhlvyB3EqgupMpm62Jqq1nWadnmUORW6UiNHee0NjX/P/nfP+kuSxFDZngtWF4
YlAL3zJfOg/CUTsJ285AU797MT/7VN5+rdXPbfKpPMGxacXEek8q45pmXo2/1yRp
S52FtGuighGu7kU1NMP+z//cnsJ33tK25ToaAS1QB47bTGzyj0BVKXm1wmtOsg0x
HuixlhwZjTDlZCZhtQgEhQesXpAyJjwGNap/JtmnwexxIGHDRWUGSysOdG2UeG/W
J4fBV+455NFJ1a5DdMrQyqUnqvGpqh+Z5gKpLXWukbiiV2KcJXgGqFT9VTo78P1c
aFoGmXxvCPYpaNa0UnxTk1LqqWRQvHViuOec2Heo9oX3C7oCPTVUBEryh+tnSozr
VFVwNqzDYmpJwJHYFMJpw0pE/fzvcAjD58bwJMXTmYesVwCJ1zOP6KsxYC3MavY3
NXCE/CxLvxcTb9JGnt8PJKgX7SWF85hvzwvu5PVcRterXbVZzNV5+/w1pOlHSdbi
/CoLdoQYYy97v38yhxckFA2qommTCxxmHO2rVlr8XIQ5v+c2wcCak37nEHTyCMVI
3O1UUFcDI6NTZbnHbpz1uvvUWfNrcDzE09BDNuf4ZyDFU+yK3Z9scPX1L16IXvw2
aXkNdEYgub6zpTHAkB42yPoRzn9tuVZJcVTgeHvU1mEFDLfkKNso/jQTJJ8SRofU
c0Oy8SimxvYxWjqwtCeAWMfC+wssnhH8q0IG0L/A3/paV+aVz6sEXCFSvnKY4C12
j/hKH8lK7g+mHsmB3RMIqa1cGsLW5CkagWC4sEu2H3bgt9jRa52dfpYdUzCIUNnd
XM7C9ndmxXEzQcOvFzA8oel03oXrr/HrQn7k26Mx0ck4u3Kmv8ONSpHW1o5XAEq8
RTGZGuHwAuf3ikc4G8LFpHV310alT/JhcfG1Z8EQ+RfO6D3rvRE/joJuyjZYFYZI
oA6e4AcG1Hs4J/I+01SD+XYloAWJJeXGlcFnfar+uVJb42MVlSE276vKqmllzIvo
55hu1WBah6WGm/plsdYOtpqmI5xD2V6rRAuaStWPtN7GU89U7IZVEpHfM8oJQ6Ch
aDS9yRMR4nmhB9UfjFdWTnYvfRRbfrHUR6lHnNomf+G7ZmQOI5qQDgmCG68S5glC
DYBkXWNOr81hDmu1JDq6/1aafq7lkH0M2PMLH2BsMprVcFYQMW2O6IvjpP5gcdkU
kXS6jUEEmtCmV1lfShPmUydymcI2t489o4xaP/oReMzrX04tlT90cRB3AYNtrjIv
3oWSbXRatVcbWb8YFCvE31PCeKxAIgD4DhlL4G6Bnbc539aA0WH8uCE6SwqWQSB4
fj+q9m2+ks18zaeW7u8LnF3JHSjKjbE16h3tQHfiN8kCuaTXrPf2ImJpeBdsrUCR
/pwk2sp9NdleqzqHZ+lk1CWEg1AvTo4vIF31dfK5qzr38Q2z6zg83xQbvE/kCIBl
XJVMWgj0QzXoRdZWY8cQrCFW2vU0jTnZGhpUajaG2mlyGF8mMRfIiNK4I2yuJAN7
SWWe3YXCZrzqwTLbaYDD5k1C9pwbbt7nzl/mD1RiBXT/c5knraKrBJv1H/qfu39d
Rb2w8oH6M87RL1uYmDZD0HOztp3YAgJNoiIovmBJ7ChiY692zJPHQhHsI5I2Z83o
m9kVWxCajnytZAHMEITXEOaZfd2osKHAcAov4fscF/sfICOnpQtbmwlWqSHI9Rry
tDzOLGvs007vOooc3EYyoD+7UVY0vmihIlPIwntrf/UCgoK8n+zyFEiihvoMzslC
h35CVthXEg9bvpn23iTQJO0sE4vZzhXT4EHuo1Obb8aW0qb/fwED3l6tIqlGxe7A
QKPykb/eyu0WTp3CftN0s6mOOR8sEtaAtv555XmtItDAGQxwo2mMZAZBi1HIJt9k
vKRvq8qRTg/ZwQI90MUJYmNnNnJK28lD6RrJ45LdaYjpX97oosy6I06wkWEBokrs
k2HXixRCJeEG701Pkf1r6C3adDGLMlUbceWfWQmlEFkCid3qSoFUTvDA18GIS4Zc
0tcr2G6Ysgi7dRxyP0xasNeipo08Fyb17jX4p6mnzWmgAfxP90jjzSgHXLaFI4+z
oUDLzXfb/oc2ATXjM7zDpWL5KEZU+28n9hLqUfxWCJUWU15uZkjB4kC8oT73+TOZ
UUpMOBDqcg9O1Xk4SML4v6O6X99rG9cfRJ1Ln3SjW30rmUU5bN9FErR4dvaksrEF
/xxwtyk/QkBg8nJ52fR/IODfMVMuJLwpeW/gq/XJpMTZHR/Iuzv6YbGP/z7bXDMB
gq58uhv34oL3ed0Sq3PzTizu4MDgaN4YUYYYtDJZZrDtrSODlBmLBiFzV3eTGbUx
gOoI9mV1L0/2x5JCKyISIV/QeJnB6c6bcS266UaT77VcbPvsx1ON5oxjbbZZl1rN
9Gh2mwg68LamOJOIfzvENxI1+BjZviHhode738oup+jMB5+zxUzTqLLxHPT1YSg2
X6QyiR1umdhTouA25PtpemvmHvDFjIvXg/KxYiUP5YtP7EvnqkiAhf3QuZKIjBSR
zpBl2Byp7GACI11zVxgCws+sXuxM9VMQiPHvE1cEZy+mh49T9CH5gPDKt9Sptnkz
aUBrXBgBxXgHTtzYtYpdX9+2kq2M2ScAU3hsKFyjYU33kEWTWZR5CgO7YSQRqBlL
1HVzClwlDQvrWucwU53ttqRgMrudrzqaLmiomePieBsCiUZPCYdUBVL18suNnZ1/
EA/rAbv91fA8CvUS+EtOeKbjrhx5oM9eKjt2LimCbunFTwGZQVAR/plXDpH1ra1M
rMulWPrvzpuqgGeDpoqrIeeOt2TYcQhwfAXYD7q7v1lkEDvJZmWSRHbPlIZWUFb2
N0jVMi/KC44eTe6l051AOiqo1nJFD9pc8wNUGuQ0NCm1i3VyyIzormPpOMJvYSis
EMIrB5rdmXWGt+N/SvmQyTAdEvCuSL2ic1+zfc8YVnJ30Zjrror0YVW5SskwhkmM
HTMx5UBbqqGP7weT5YOBXPfYlkVptIdLHgKIyaRU5x1Zau5wOT7GXcUPE6Pickqw
9R3pGxzc0OnkTvmpWPp28W//hYmIz7jn//WpkPN9MofKLdeDvUjyaoZTYGa+GVn0
mnN8PYwIj3Adl+i8qb6SpV5lGRXMHvaBCCO8hNEmc1uIGz6BjNhMjROxCjH7tnjt
EjbsZvZ2V5jt23yRA2GXUYybU9y56x+4HKj7TxfdZUI7Oc6afL/A9XvAff4DangU
ZWQcXcwmRBAvCu19/uv+kb0q2KPCLhFkW6Xu/SPD87ymGZ3Y+9GU+KPm6TQ5D5H3
gFFj2iNIzOOARavhox4VcWmF/gn7TlQdXcyXLPnWwPjGgW9X6P2Wu2UHqM4e/Vgl
OdlHPzuzN+8TYf17qrvDlAhTCbBgUMGqi8CSy3SiAseb5gfxxzTWJma5roAx2XIv
N+Xee+sYAUY/GDY/O4l6R7TCINnCju/a27X/lI7f9JWqr3L9gEu5uw8I6EDzdlFn
Q2x1+4k6fOx73j8v3r/DrZLAVjlH5wvwQQZl06D4y+rbHErMZGXBLLfEq8GbyyI5
goLnkZ4LREmrU4OJzmZUyPQFHKCxPzd2nRRHjWwfT4MJbCJmKXmPqOalvOVYAATu
tNurG3CgnVlz04Ei+sfn3p6a6jKlKw8DU+ZCta5EAr18UQDd51wxcxaTobf40BgY
ZVlmPseX3PRu7ScxGogdf53YBxZ6/+uMwNaf08PJ5vwYaC8aIZ3GtNo6vCN12cXo
Iv92e0msJjjaEAX3iKb8sFkeR6K6V0gNwBNu7q+FFFnQBc3OpVTWn7oAQcsJIL+b
Kp95ZCq+vYlMkHjw+jBA8FqEoE85DL8o5nR9jZHpeGpSLGBELUFJDXbMTtckzFbH
UnTSHB+Xs32pa+UMk4polKeLhEw39ViQsIlUHdmhbYe/ntgU2Tkr4DXWcQqD9e9V
1ky563aq9E2LzFGWZsX4QDm6AjjbigVb6mFmNHItJQCRB6Hk2uFEjn/1rNLBvnru
uUPfqb5xCP9F6qhreJE62z/vPDokS37dvosVEp93aBtLV98x6jBMldcvZywL4TOV
cmGhgqgwPU6TZXIZHPED7O0UoSbqtAp5TAcce5QPOCRsHeebO4VaJmC87hVNQXrc
BQAcK34xGnwSWs9Lla+Ymom0DMSb43X7bH63FObU3OWvE7PZr17aZ2q1fstRw130
/yVt2W4xuQo6DJJnh/PvaG+owYbhQoVfz55LUEv0/wg61PKLLAGYZETYS/pycDKF
zCpOgmI97iCa4yKJBVf5PhHnw7QrG/rlieIk9Namb861Xd4NV6YTDzAnQ3G6fRBQ
ytCu9BL4Y/bpUS27h+C//443H/Q7MFOvzcPFKsNgQfgEe7OB/3foIr12yxYGSjLu
v2XG/3Z/laO1TBIR1Sd71GCx3gAdX/FhK/viaN0TwYNs6HVH0AFDIJwx99MuthWe
IpWdr5s2utr/9GhwO3HoXxnmHPRxGa8M42OWRUgHdBR23/EviDSNdawf9+/BpgpE
3jsA6Wi7qTG+pXIXILbL+hRF/s2WgivTaXXKvktTifwrSGxQttuZ76U2PL/cWeco
CuO43EnKSX2WRpuW0jMq24iK+2iPzZMbtydkU21tIVb5n+8GmEtWOUplfcRTgYNa
4g+JrlHFNNKehjy1HcZHA2CaSaOx0fxdHwKEs2B4CRSNtSTs++sfDfYTNwsd0/XT
3rcvngjvpg2zPz1a28lC/tGzHHycVaCJ3vlQG0gaq9CzK3g0aCxqyGs+rJuHznQl
BKGXWsurz1MR17WJQPy0yIsi4hf/kjshrDUkunmYIhbINmRj6jdoCH9Uc8UH8aBi
xEfZozGWxGL1TSpFyqZRV5KzEqK2/UzynqkTNUOhtYrol8lfd/oP5bUdP+6uEQFf
NPAPkeLjSo6EnIo6dqCTNUjJ16E2/T7nYvbBkOsb2897jJylTqA3v4uR+Wmm9OyY
IfoPerGhWwantsWYei/woemjYptTgWj2lvsE136bmkQv3m7r9QnxL/AFs80IeCvO
eAMeAVcXyb/4/03a4JrFyrYleMjG4rz36MQ3VTRWsvDuxET4GrqcmCmVOZGK6DYb
JMpRJ0cL5tBQ+CVAevluSodRfg/0S0CYn3bY+oBIc1nK+0rY0iMlBGfqqn5fUXZw
WRPaAT/PHiuycn1ZRfvkSve1C2GA8iPPqiK/feEtFigbVvo+EfLXvkOJZo3UafjM
lgLHLO3+oKQpyU1pABWNQ9Rs1eSo1Z+hkR4Hn3yZTJDAKYym5tP314s0HnKeasqj
IKZUg+N1s7fpdMIsNG5RcQS6mYcctXYg3a4BAJ7HnTBBckWRvD1Eibt77oebYOCs
yurjdE3EnjhDOEN80HTvrPfQQOsjuf0uHqu6rVbWDAAxNcS0lAzlrzbEScH2h4mR
5kPiG4UaGeDt22QUD5UQ7DUxf5Ml3WSdQKrs/dmE4hlt+iJM7l5E0yl4zwZnwslC
6AxBR18dzNAwY4V+kz8+GewnrQ3EaYOLYBABAs8XbG7PMqmRYN1rNCT2IM/xNisq
xN8EHswkFZEwhzsY294LugIDmAbJdGk9JPkyjcSMKX9sfto47drib52Cpk5Mhtkr
OSrFi9ocPyRQwCi6R6UNINdB7xtCW2xr4z6u0PjXbz4CRPiVKRro+iteL+ld4GD8
4hyZn0tZlfP8VmFwGw4f6fMFgyLSgr1FDakscIytcz/C8cCKXQ0hO4pat/fdH4Qd
U1VR2AqVliU8zptHlF514hGoOLcrZVHcUqBhjH6vOiOOYmaGBNu5w7lZvbxDYMlD
Q+MX2mhs8w/DoiaGAc3M+Zwm3zGmUtn+2PBgRwUm4+JLJY9CM7AWMulZKeDZ7BUe
8TzZCCDj89a9I2yTLWeaCdFEbun4iBr86v4iqomm3PrR6EulUymtEnGd7ghHtQGv
Rwpr/zBKAKIE8RocVwPWw+QFzr/2MiX7yYrP7PT5gqBS5N+6mmN708ZQ8YfQa5Wg
emrUJlKz6mANhQx8NNZxJxlTYPSJ1zlVrryUq7jmKgjRLIjZyegrb1gaPKtpMyRM
W7kYdhmlyjy5Yh8E2aAaTbldKLmHOCeQTyvlC0w0Gjv5NByXun/RxPmK0DfHvtq1
jvBDGYiFwmpa6nSaJovcC437CreeHZ17DuSEU+yHxH/Af71dyb/I6wMboRk/Bdxi
h7WjVaZ8J/xZyGXjzemgyJshFub5d0wugHyPJY2vjT2Up9hG1Gvqyy+zwp6hXRHJ
JgcGrvhhNLpjc3rmU9n+Vh3gF7Mc67XZSOMsE4Nfvon7yWeAu2hRs7cg0ps+056+
QehBXKucTkEwbAxUJlzrNmkyfyfQp0Ab3HwYN2WujvbJkLGMI9dakxCCloYTZXcQ
J9aKTbh66lkwjF8tC1QGHZQy6BqWsvNBJFz71vKylNYJFk68OLz3t1ouBt4Xa4l3
2cHMka5T3L/K0Uu6Qe9N1yUvxTsLa8ZkwvKLoKEMuVBfHy5DcSIDHEptlhqkjPG9
BEqSoezyhfaoCUD9jRc5fomLwt7rCacDvb4+Kac3dyJ8/TGJ5RoCVN2VCTTV6TxP
+sTVkuAfHe6c446CNVGFVju3WntwatfKhDl7uxVi3C0CmPUaCWy/Wa8eSuq5wILF
o7Y8I2ev5dMeGARkbJVga/x+tcN9MF9R9KPQlyh6oN4EodONSOwlEAAhEnKNwjWC
3U6NJnyxhRcITwdeH+GuQO2d+5gsNjO5OZSpUni3VP+Wj9ub+enLz6caIbvU2lo4
OmeenK23KYVWDT2fDuQ/4XUlRi6O2h5BR4+Pe9hE3XL4bGnaBm6KL8ospEXTVj0U
feBLoPlHfCopUVNs+4Wg6wf19QFtazy24q0iJ7UPJnYY/xL2HqCZ3vg4VCVSWZ3s
w8f1XNEGBhfvzlizSfTqTxweg1XFweYi8nY2b5OyJBTPQUhEffOZJ6k7JO7NIU6s
RLkPeHbGM6Kbjc8++q/5miXBZ5GFJ8Mn0goGIJEEBQNRQ7vRsJgWjJffKMJObL7r
CeI9RP00M+j4JEgb9W84wD+ncDlYwwxWv+TG9JKf+L8WgUwjdlw3Sq0+PWh8zW1L
6s7P4jaSbjxF8cZ1IMdCgY5TdlwQcEcx4SQ6tbzTcXLRomn2is2zCgCarvKA/wj1
iSR6KJgW0/gBrlyNpP3vubRp3mZQ5La1P6Tezt1nn1f0+W0bKqcE6X0Wof8rb4EP
aYDDYaSDd/WjyvZtX6cUzqkLos9wzDhIeq6E4rZzpxj+PRYHY8Dqh4AWQoukzBDM
cTg7Z78DRCWymLPrzjuJCawOIMdP5TeaXHtKymtfwTvvTM1wWAOh0wLILMtFv6i7
/6J3hbFei0gkfqghrppdTrmGfgaVuZmHTlMSUW8GouRRX3qZ/4KxZKy4ESVqAjIz
gYvBc2+/QJO6rtRum7aK6nLXXE8N+GzOklmiVRvpgaadQ+fQj3/tsahFBEYSFCNp
/j8QqhofJBDax6JDvxJXRyH8rqa6eVWOE/xwSAy1/HpERPQVl+T7t8N3s9TjP2TS
ZIHDceUus6uyWUBZjp42g7zw6A7xLZ5LAsq27jcvAGDqjmQbHjaU7cp0ZzVzvbvy
uWpxP2w7UpnJLY9vx3B0FMiwyHgysOWK67b6jEkC6gMoEMzGxqNJFBlQXGqOS4aN
YXufWxI3K/YLcD0QykwFbTnahq3BTDlNr8bwe39Cs+HvGD+ld4Cp9/lDQTmoWLjK
eAI32rGvD2b30lshp1dQyzWUBDf1uuBR16vrFjWrQ98ntVEVEW87cY2S1Vcj2MU2
U4AzpV2vq3QL/7VAtQwOne9ATMcddg1+aEIIKYwCx9Etkk5KQ47SM5/Q7pr1Piu9
XaV9fi/qErZ4HmDVhBDn9GmlMN1AKi+LRHYLG4EcIFsXetJ2ha5DvKX+vAcCa7dr
sNL8NmWNle8aVeO6J6hhCfZPtg42I9s+/FzcBQvIAsekHCFjykVmIbM2e07PS4ik
DDyqSNefGx8UzeRHIbCa/tZm0MOtzHp+a4OeoS1zPmLnBnRTmadVxCku/L1SLAtq
s1WDovdMTCyr7o1fKxlHa6fpbo4f3tcz+OnGpSq4c612O3o0CUd+TmqaJY5kCr+r
CiktMzH88sqCew1AQS4PUjQBMuQidil8RtkPeTl74aHYmUstDw+7BgCcYofZ1lAY
/MW21dmW07k+znXCu7D0E3Ngl6iFYyjTXOY0qplRvqmz44ACupda3cCGcdNpf+cX
B0fsEpHy2riLHqbbsGlCgjyBi6tH5zjuTGhVF0mU9Tn3dShf3RNuWOa52ax8s8tB
eXkPXxJ2q7+tQ4Y3mZ1O/XV2pYwEyC2912z7CXfnTZXEng37vgY2vZhLuxZW8HqD
7lDlhr9D6QdkTaFKtr2VfHt4JayHN5+ggN8IDA+vIsJlQMKZ8wMspwyERrF5yKsg
4S3U6nhg9R/KPVy/5J7i9buQZB6pYyYxdXL++qrlbyS/WqfKTUras7bfl/eGR06F
bv0jshDtw+vT+/TyiB4lmuUCqXdJQ/wELit7nqKjDeplgfBKeib4zOiX/0cneHLN
cD/EJeP5I+aAkLmg5CCfbS5mb09WSYP0qxq5LlYeDWtzQ4CkpdHvu+2gp81CKGew
94I1QkDtZIM9fSax59JJ661LcEA9BYJ60dqcD/fivTAMiZHVM19+cyCfBUU43yGv
rMm+WoGDgOTKnt6ZYGlQ/T9D35uRUcalHKc2gWfvwKUPle//yS07iahyIYRA1KGg
tIR2weUK1ESRA9KJnWgYZgZdWUo5WygIYFJCVgSBJkrKTwGbrFyGCJJAxrAE2DFE
FDHPwqfneHuhlT9bxn1pS7s88K27ZpUkeC9pke6o0azjTwO2TzDxqc2lVNDzuhNW
ut4VDHtlENaszVVSUKNbDjPdoC9sWgerOsIb3pKYv3jmMtQu+LAli4jbJdhu9vy7
UJF2itCyiUopjPvxt/ppjswUL76yPU2K37TjM7oNDovoMm8TaUDchoW+fJM7pz15
1ONk6w+l42PyL2w4Z2o4Oc58UXiDghWoOmoNlCtUFLXJfoKxo33uxIEAg2qVtuur
m2LweSeuiusyyA+dJz5vyEtU2DQaAQoqdJb+cIqPpPqzS9L7v3qFureF6PcesQOj
Qg6MD43xmgyyEr9/nH1d8H8T5cBPgGFZ5tZHxouksuT9irvf5COEsRSEeLISwB66
s7quOttblHWTkvs6TvhYkU40cVN/iRaJ2woYpakxb/k0pFSUcLTfZob3tfjkceAO
foqA9Ghz8Fq8Q8UULbpDJFyaI3JZTG6Tr76gq1sGxA1pr3g8w0o0fYhAovgn1X+t
IY8fZ0/XZYguVR3OxByRrm8rJn4C+6Dln5gCvMYTxJCRA8gtn21Mq7Uc6JJxkeKR
kEdpP3VsusdiuuPV0PViiMFljwbO7n6HKNiHvuwH+4xeos85pxvQUY4fkGczvqf/
PpkU/s1XKc4nH3NZqaQ3paGPVcGsJvUHgmRVbk0eneifYoYocNMMVlUul4mzjHJ7
BLEFuIBPVo2fY0OILJpvPS5aymHH6cC/n/ssq/6wWCg4gvVEoMaQZAOTpUip+ZTd
ot4tguddK+qlQzkCf4QZVp1ZXg5ppFrfHuBL14gt74LD3cRmd0SToBBIUbfnWvbI
oFotjAcBaOHJ057hkjK4aSHwFMMz9QMq9EyUN9Qwraxdh5ROTFc7Y5bKlRbUK0CK
zSPyD417wM30FdqMfJULsPWfuutABuqYH+DC34prbo1uEqg0MrAX40jdFVruyrgq
ERtxgsVxRDHgvAXDCPs6VzwpgmEM7ICjKSLg9yedvj7lPpAbUlgcImmv+Tb1WqMF
FT6HZL2SgQSvJpYjdLksCok18twR21ky02ICu4dw1saK0LzRj+rBpB+J9F6I+p1y
IJuWd9fUC+wxfsB5Ddhw8dO2X2INH2+NaaFjLxLl6JdQr2bzTw6IY4dXYWynp5/D
5SK3M0alKCFrJCizQQ7ubM4zQQMMMGA8+kTO1lpHO/96cf3/hGN18cNu4ZIlVx7H
btAH8ybMqekIBYzgZd/Fdj7PDjI1ez6UIPh+eorL//RyOYzbL6Z8u+m4v3gBNwmE
ThntITRHsMQ6Xyyc900sE3bpV9xS3UR2mL70jLy4PntpUzzSVOHb22RlWYR4DSQX
3kRgaaXnDHERsY5PkBoVeeirFx85ZoHGv4uM7XRino/TbNGcSFj6bRpOwtHqkx87
M3qr85QqlFfhqKAUi/NMzCXGrsQOMGBZ6Fx3+N7MfF1pKY9NvCSU5MsBY/lw0ztP
9jubXDEsfFy9tc/f2+EVZYIAwZqRa6vnH5pmsfbyMpoLOwCTbdtkjL1L5n36SZaN
POJwuHXcqN4c5pNDrTxWwsdSyGCDBo+YrW27j9eDM1p6sSprDAsi3wa/5A+zH39Z
0taGR2YpEODODcH8R6ICYTRJkgiPDfdYC5oWbpTOh9Z64HsXFnvGIfT29b9D4rRy
7SVdRqfeIS3hxKjtE2oufEMH6Dkkc39OPLbYAzWpnFTO4yK7fsx5p79tg+vf+Vud
5PiQ0uHoOR/oCntBuYDtzRGpFJttvCTU28ORmgDO2OOeGoYYBp1XshNeEIIN0OVp
fiYsyGHaXi+M0mJOye7rg+iwzNmii9q3gruu73tPwZ5bH3YOEujTZhHHvlNgcJWd
8hKCVORLT47FAJUXtuJXEkRzutVd8sUONR8bMee/ZxqJoqpCnwsi1PnH4v7znaaX
Iwz4X5q8QSWVquyTv83fZwUGVY4kUDL4k2pO8//HbObx9gF7Bts0PIiSJuCvNpnJ
wtMQ/q9xSctikqnox+DKobQxUj7Uc2rGu0rfv+9YZVShwcSbCFM1+t1RZcczW6hB
C6ybjhMmF+/+Ep31xwfykmM5ZW3GXNGQEy7mkHp0RNGMjRCkUHVmWI5q4t2tjBrT
kW/DXA6WGTg+krZXbAwGbxojEmhR3FPSogkvJm2dvc+M0uUWeBWiZHovVxnE27xg
qt08hoOazEq5x4iaDVpT53LPeco1wlmGKMIJQhCk1zfImu9ftpqiAxNYLLbm75nw
P8FR5a/geTxwYT9qHXIkdluc7EGmO5xcq7OpCHwSL1ayznCd8KjVic2kn11FwTWO
kRbutqFSODbho+QZsqv17o3be8gi1GzJ4U9aPVkoOyLDVigEXCjP6ACxCnalOcSq
7fQDgjouMZbptYw+6nVOcxgOu3BnCLVQAIXa7nHpeptNAIqBhUT0oPBAfTunF1tz
Sks/gk64Ah53FCtaCCPcCMeoszZpQaeDE/KSOSCDc5YkLKh+IVSWpQB5Q8bJLBwB
xkZUOleP7W+XzRoe4UXqFndHByralBfEAbxTGTsheVq3O5BchhgObYGVmcus9JTH
UfuHy1n6o8Zz5NmEqZ5tY71N/ZhsJxvnl9ChVAXtjWsBsnNm7CbdbfYE7pQfPnBg
AIABAL+7KekfNzOXwsILuwa0Za3mKQ59ftMamyxDhVgOsxNJG0UMn0ghvgClVS5K
or0/OajQEzQKooehqpJcWxqpLIsArJDL4cVIw5uq0UU80b5//xihtF410bge4riL
5oqPXXxluA5nY+bGFxlH9cz7Oo5lyGTdoea95uJ1AGLl1IeBggK4gdunKokMcg5B
lOSAZUEn0uz76A4u03R+zNdJh6QpYI5yQIVXzBQzGt+2oCECkHYCsmzeud3uvxuO
wsAa4fWf4n9YnWJfh6tELwF5YJiZvWl+P1jueSDtIWoUom5mJYqlNQo+T4s8gvmJ
7+JfF8aHvOVQljADG4KCLoRHyFUGBlch2yj2b4zMsYE1SlVqxBrZQXMln98GLdvL
TL8L1SPcbMYheeUzona78Aa0Z/SYc2KyaCM1MZlSpwGT/0I7RYuT1ool91Di9xtY
x0ienjshfziNcPsDXUl7/PYdGBkf668pNrsEGcNo9hZizPQ5/bZxmT6+NLl/1l8Z
IJKf6OFQ1lqCuNRzNBt3rGbB3uY2f64dak0S50ae69byuJ4xjWej89V8ADEDhqpt
jOs+8GrHMYEIo7VnGEYdbl65z96wj0PqG8JLi0uLpUKVXTSxIh8xjCvqDuIQHQWt
v4RxOztoGcR1rwQi0KPPLUDRHUDnHfe53rjwany+qx9M1GjIfPmb5bREO/iIH2mw
CcKSJBSrVS6MB3YN4TsxArX/SO2m3bv9DZy1BZOcgawC//tSzzVVP+2ELknUH57+
ueDuxuARryWk315IfCDH05tYsIlpIz2Z8i++o69YXE/2NuOtPr65ftPRuWUt9RKR
WXPV6RaZUH4sdXfZexL+YSm/p3f5buNKJZf3ol+B8jAfRDy+8pNgufWOluSZ9637
elNhK7JXSdquEVNQlvJcOJ+Ek91coaeJa7u1ZiE7dqMj7VmQDEwtkoPDtao343/L
I19MuOs0nbj/doD7rbNS5Q0xNQdGRAfhDcIL3RxqpRjUyJy9dKW5+Xln8BPCf/d0
5mAhyumrE0T29Suj2x4JuFVstdVe0C/m8oHv+F5DosNN38psYAj6mxNVNtoy5D3U
ZztbeMwzcW2zBG1wZ4qSZc15BzPdp9qzl51ed5xu15aYVIM4Fm+A27ctP/p69Se+
bkd1Rym/Np+UssVxL8AiyuR7uLJXO4mCjk5rveqlwE5ujFaYDB0BBj8q3NCYrSH7
w3siqNmWzyv5PytkTYXPqQVcjdsT9AodI9EyJJeBYtTx0g2msbkQ0toSBKzO0oXW
lYhmFxfw5jqEm8zGae1Mc+vK+tZtflo9ACe5n4QdWFO5b1N1RaL67+b0FhYzm3fb
53nGyMnEaKdpl2l3UnQABv0FtTvoLoM1fsjXLzvqPuEi+DUIwXyX8H001ct/ZOZu
wkFdLBK8aKfortm7a61aG4vfuJWrlnL36fZRqYQV30Go0yR5l+RAX5qQWb4aQa7c
uPLafsVTUKsM7mC12ih4Iftk4v+OudY1TkscdGuNLyuzFe9dx+8DtgoYjQK5NFhM
QVERzFC4j5nNv0uKVs4ortxUD1xofzIHj1mSjVOaeCzCUwX+AGlJA/znF7HjYn5f
JMqTaSXJAd0hSCS2h0l+FzBkQ3ortMF5xCu/SmIqnYfNfo4h56VUhkFHyfU6OF4c
HJZbYX6cGtMWm1Z8xCrOH24sww50G0auwDVHparMfJ16eVrcGgmjNISKbY0iWwWl
HykhVr4nXp00O4vv/6gzY6kAflN+mRXisKqq40Cg0SMbhRmt969YAlrX3A2APOua
TSzFlUrQxwol/Vwe91C39dS/BOjay3+8FOC7b3tMqpWpA8fyIXg8x+PWQfA2g7Xu
FY3VMIJKyrElyJEIbpkaz7Ur4p0fM4+JjwzE1gyVwhDo6IJNwBvTly/MG6ks2sQn
pdZ54CqTSt+MThosoSXjwNank0NAH3A5UUC7unr1UovLtk9I/3NH8fvUaqYL0YK3
Yivc48Rlx1QfKut+hu4ICU16gxt5LoKthy9L5fwCsk8Pe409wBXcsV20BSiVlIcd
/xiPNpIMKyh1/vlOJ03Nb69vAxn7BBUpjjJBDxAN1RKdc4Xfo/IxftVTdiI+BrFp
SX/uc4+k4f39ECCdI1lC6+MEarg9AZ+X8B5GUSVADKnf6csW0y+tl6megpAXAc5D
uJupIPwVqL06+uEpul/d95ftLtXJ0AzTaTKIA/GPvc2tBCYPpf2HtoM3pP66tkuJ
PtU3fTblJWagYqDNatMwe7Qxw3GeinLmPWPgL7ZTMPARcI58FFgDvn/kY4+gCGqO
d0tFwAZOhWdqVdT22oNdV48cyjR5aZTYg7Y1OfQkunAfHxqsUd95EKLzuj+O8lpM
4HzZRNBin6pijcsCEOuu3bBXRTA/CYPN6nRCNWdYSYjiocaT5AIVYJtwS4cIcIsw
LLMGVIW1lp8GvDHI0MgYFivgTjVc4OY7URZgPOLctyc6vbK6XFjMAqC0MljsrDrJ
FQQhe2tYGHm2jfUnePxCczRexLTUUAvjW7NyRX0DT6dRE0dNNqwbT5zbFBzt9Vpq
W/Mg80NVRt0v9rVDCW4xNUvQxKRylXHI2ShiH91yMUevh8Mmt15pIf6tzePFHr07
FTMQqmdjP+wQfptGoj5ae+whGlwElYo6RDt8uuzq5fJDHV5wovIq01R5HafD9vSc
3fhY7N+2lHhnSaMUlIJUK/kbY4jVUibzcbRnWF6U8xxx537/omBRlWxDkCH0oJ6G
iSIbKq8FGX4c65oZKqWEOnp1+hhW1BiYxovK23JJ4qC0mtwEJsOPyX7gm8ospn5W
i5GEEIGfVxnjoae3mUxInkVSzT8wJcqBBX3gg+lIsT8p64YhvPBcZpp4GtarGX5q
0D621Qq2mhm1pwrAbSicmUz6Bc/FIkd8EcWOuCsyrfD9fAUCOXYeXQ5HkqwT94zP
Tnk+oZlvXE4+abeWjYcDGU4BtR7ipsPLk2SjnlWkiWHA6WJqqTHekXd/FIWJbcdB
+PmO9+S2v6zuk45ppyn/WMY5/+pUx4R4iroNlfI5ODlVfYJEPRLovZmdbH4yPGP1
Gf7TGsikU820CuC+CzJa7pXAeDqJIQwk8Tl5CXLG9M5zSUDlXH4wcxTQpfx/0S1e
PDRpPYWevRA3EmhZW5lcvbftDKcGFQ88TyWu9KAP4Xk183RaPtKuVnvFn1+nilB4
XMfHfZ4nDOOMxXcd6iTkep2zPShP1johRLbQ5NmaFpSC9neIt58bpgQWnwrTuiOB
3HftrzhSmBA1Dp64xgdg2IfO5TJqUCaiwx1RZQohgUvLttIcZGh8QOiyZ0N/sDbI
81NW/rRA2NmBSCUPsI0hqJGnsv34NXogJSoeKLgisr4gfLhvOpxDGGYY10pReZSm
rMSD3WRACA0q+s2JymBqooKDGspcyfLOs+WIHzfayWcGzKN3aawNLebrozbt77u0
DJr9j8e1ulqw6vyePEqsR+HKny+m4giT9h/trFau+KgXfUz5Y9rUiH/mGdJoPztg
iSOI+0DySByhqD1EBvzFW2WCwIbRTFpFmujTVFENhGN4LeQAoYol+b7SDZwXpYcU
p2n9IqwesSrCZf2/9V/ECz+qgPLw9YBsunBA4PI79+CGLez6ejwvWo1Fe48y9xEL
Cm2P/UxBo5rcH4J2LUKEKC405YNtxj2pyF9jEEJwlh/k5UIr6eBbKIO89zw5bZgB
owYCwUKGv29rV8e9FWhWgxZ4OEGq9xNEKMiitsHWS5mynx4PLnnh0wueqY+BV4K3
aLI4R7ghKA28n2DENOwSlkVynXhRERVLBU4uLq+hrOILcbX+RilCYTsMAdjY45fJ
K1lX29xw1/mNFX13Ro371zbpvbfZ9UEJbJqOFiAbdZh9xDuK6mOc3e6LS84BLI6x
RH5Bm46E1zMmMRjenkixjQiDnjZ8NU/iA7HCMs0NVOL7bEOrFGXj3EJfhu6RPtJz
59KeXT1Yx3geKVajRcxKUBKWjyxZiDAF69PM4VPpXqmqUucDoNZLnkFZPuBsYMRd
JGR0QisfmKdX7wWeE4KOf+MCn2bIqlg4Ip2kktxZm2xQ2F1YgRJIDz8OnAyTyy8e
LpJMzE1xDriTnfC5vT5R3gIUNoR1JHvKdPsYNJBVvJyiSreTPEo8mHh2B1IsR09L
YT1k8FI2cSQlabK8/6pl72EejuU+v2LW6NbFUl6bWTSFEq6TOHIO8vu1T9GWwJpT
EJ5GbxvkMIuXwgwxzEXvWpJB1hVfYvf59gvVwjyHX9V0NHvVq+SbPNDTV1wlQpSq
/eBiiG/gDj5G7PfuTekxZjp3kE46LfRsAkOlZZFAqiHkYRZx+JYdyAErkQkiI1j0
7QCwzyaDX1CFrAq7EZ6itqD9RgkZfr9EIVya3Mo/pxAfOkLkAgrvwkRiEjDAvtBL
9M7i9h7ATo688snNyv6m/yxfFLcFTP4cn8LjLeeV2N/OQYyG6KXqwQpMiH+hCcfL
dmrr5YNIPYj5x2o5b+6CEMr3+SbXMvXaubeN//opBXNuYzgHw1q8zYfQ+FjwRqtj
h1Av6NMQ3WDpRmC577UIyn25SYvKQMm6tCOOUpY7c8CzqLR39/jBYnWqWsXlD3Gh
QmqepXxhaT+E07HhxJ9n624oP9uaqHrFAoiDJc/rr1UsnXePjT/AY5D1tOE3TGtR
cx+ofLYWUogBgRhBM4ONHBqPR0ke2U6g1htIE4jIDgjNL/2hbZ6qBpCYptYn886G
RGyNdeB4EOGeAruyAfF/KCqLATNBzNsm9zONvJ32D1GwO3B95gSI+za3YfFASafu
nZRq6lkTw/c68WllM4jj9S7vzWmHUSBRvo1L56vyu0Ax8QKs9iJQsU67uuKhetgZ
FyHjIo8mQ9uPurssLn+aaPj/dqT8MbrdIyGPvi1dfobD9BSdeLC7Aog4jyD/m2e6
moHlgitkjdodjywSefu5lG6NbXQ+dhDZGjQM8OSIcBGNnT3Xcxzhh8Bq+WlbjlyU
d7xyevR9Jyincmmzd24pEvzrWRkQSvjk0HLCwcSzhjvnbYijVX19Ivbfo/sDhAGa
+tnsd8PbxtnxD4/ok8qUnl+mBWKfG72SHXjeNi1xVQNOpCY84dIh3rLaVz0shUmg
t5RhMA1mKrue3We8qZ0xNulaj21itffWBQAJID07NB2zsnySIRTViFVXMf8r7ilE
6/15S5VygfO9T3QDGPrr7GRp29L5+7MlakLhfZt28WpQm2/UVX3S7BZyZ97wlUe8
4JRXNw+lEHXH+qHZUdD3VHIOgFdY6vBvvYxDEVICpk7PKgcTs4tR5Jok72cIyaLf
A7eBHm0NKDvbrgMPVKX40fDAV7o9/iUsKysHiZoOBOrQ+fdx08EVvRVBokTgpnlz
tQB3sZ6n0M0CIwJSuFD2MRty8HZkHWcoSDiqFNHDnGyADaTmtwVZ2tN2EbekpLQ3
9c0dTRPlYLAl1KRYJ4sFB/2w+D98Eca+SGs2qI3rynb8nCAWyrJy0ObIX7dsRo92
BR1Kl3ti6O8Gd+3IvnNsAfrhH2kdiKc/xVjBg0tnHnwsNe4Rc0/cufDVA5pPbx5z
4zW3cjszCt7QLf4CtMUL7JD6CqDwfqywV7UJ41Fbawfe1z8VCKr2p990JmEwjg13
cZJ9N547sVNErKyU4Cf/Auv/nEZEpFY+lLEoYc3R6zl15mr+RKeCv3x59PxFnRl2
hSnqJjF9ID4SqRUCUf0Ixc+g9Nwh5hQMPuE1fLdm0fh7x3BwmLmf84AjG9CeOf+1
E/RkxlL6+MvBnUhP9mpj0f2iufhU6YkKGHbjqNqNWwnnEW4Vpu2fdMSmCRgisvEC
BqRrKwS/5Hsqk8gO19IcS9NTQ3gC0VoT6pIr6WF6/gMxs+N/pODRbxy3O51Bxp/z
UUf1Ckp997t9iQZ0ZQbyxYHwj7laNsjd7aumjcM36nzEv3l9r2uxunaBoWxVAZdJ
dCUvQ3v0XP9iK6qz3DnH99OK50d5blgLGQaFLy3lp7wl2y56lyfbAUNld6+VDPGn
Z0xSlSgiAaYnGFqDZ0MmUYutyNSbeHYPRIiBX9AsK+3rTx7qB7yQqokuQdtbFdA1
/11i7LNc6mbcFE4MccDkrpx3Ufes/U7qK1kkGtS/D1kOnT4Fd95x+UnWmdygwiXQ
+D59x4hN52rneJE3CfihxpDaHPALRhjDsQCvJAIhkQvaX1cpYYp66hMFVqLisiHp
hrWg2UFWxkll9nWtFWyK+X8xkQSqGXpws80ZElrQkA/jwNHJWpmipjUU6s49WRdy
HH6I53PpJvmfeByYFU4BiOiyA8s8wM2BycCMNfY/Di3HOEhebFLj+D4e3GHYG9YN
5rb6+tIfCBlij++CT5VZRMEO/0Sh5odimlTC3XCcd4Fzy8RtX9T9NeBng+LWBjHw
TMJxm0UC/2lo6U1j+4gNVmqOucwZMfp+OGGo9tpwiN7LgzWZu2EHZenTtl2zzzSP
d4zm59e8oUJ/qcG4UpP5mLiVJV+RDR8k3B5hFK1GUXEbp70GojlkM41rUNfMI71l
34BEJRVPgArJ1aRVZfk+BlYxi/OuRa6v0lfP/EsD2gKIBzyzaOXXufjD50ogtJos
nEOMtttDxgnj4CigSEUtLb0S+tsznpiQaAM72IcmTVxHOFNvKq0UppNHtOB+mX1p
4M3ExgaB98QPO7AyWx/JzGxTS4M7rURdSTpO/uAlDHmtKY3hwu3rc0ppN2Q4eweM
I1yvqDs+5CL+Myhc8zZ+OZPwoHThkG0Y/5WBUrM9JKhVTRp6VPfUmrB8RBxSUUCT
wy92xrTmEzrmXNKHe4epEtWvHCokWUWVlYpAzFOY+wZRol5HDoVQF6q+a3gIHY1T
2BhXHocyuo5nOM3CdZiW2LaXmgbfYuzVpEhwED0BVLnB/SzsUV7j2lkrUM609gVJ
CeXgWOdqR/iqeKVOIwUAEDidSpoJqru4NXc2Mnj9i6GHOx3VOtDPQj5QD5RVnen5
EfrYXIiYzs5EOP6pLBRgZpQ5GaLoyKJu3EHyK+REe51ekFFv0IPun9DkrfCNErNn
YCNQXPSAxIG08c5YTOvTXqMy4CrukTtaeeDS86z6lPojDNbXNtyjZaEl3IqD+Ndx
a2Y9FYKmJOssNTTwu4Dyain+05vPoVbuGfBLjve0H/Hhb+17f0zENdPNi99dZyBd
tIjdujBOQ5MKMwhaFShixP+eCfCIV/tFrJmqcvT8NN2wb1Bx+1O/VGj9OkXE2awP
KwnUiUedi5NdnT9wzUoVPnyTsv8uQjXnHDDOXF/44oHsFLf5QAS9NTP7iwuUmyCw
dDLatqJA1jrxcVFXBsfvBJMpeByI5MebdD8qnn8GYdU2n108AVcVuW9WuyPkSqaU
8sgq3WnWYHo4V6B09VRNzkhpdCjvEWcE6eCNYPAhd+BqqgVPYQFMSivE206Clqw2
ZSv/zrbrKVf+t1XC4uuaIatRb1da6NAWQo4hckfgxmlZJg7rY3ZkPmLq4o6u8E1U
lgnlrgez3zJHqCebYbkvix4VtjoEESONTPjIBSK7rkjv+wWcynem9hbCuH5+9N15
m/XOUnwhoDBEqFBFj1tOMOxJYbzTwkCEDOaUSyjpNi466FKhm2BDvJzWkX/Qi5bz
QdcLyRQglpAgkzK760KjDbVD2vejZob6b6r7xejkAcJhMATALdnFZkELAx5JB96O
zuIvSufCybXrO9HPvH2sSXcDGcs7pGW3LIbmTuiN1ZNpaU5YC0zcYE7ACmzOz8bj
2CVdCvi95ToOF14sEqK7tMactFCjFX2fy44Bzc1kZCpUlU904mFDGwwyEWZ+av9I
1bZgRUVaf77QmDCikhgdozXG19C5SZtOIwnbSWSXyxifpW4Bor35T5jmmcG0q9rf
v1HsORRH1TRgDyL2EkgnlV0ZWItnBJtc/l23/xPW33x1noz8rd5dOFWHK5Q0X/M/
GNR3my3+fKAWWt0YXGeFdyHNBMpPYims9K32KL45FLyKxoLWHlnwF1ShNJmnfstr
OsbGk260VXACCkTpN7VTITbjWd7WRAFXN8bAKOn3kUmB/6JhWeFLs0mBzjQCr3sd
Tkm0TC8vslXAm30Mw0NmypvutTrMYcvcjf1IsFsO7jmDkW6ttsz0UZ6stBBRtOv9
jVbKpp4zfKJKkHcyLF/SphZCUEQJcqUXMsSpHPiLWQ8KzqzE4CJAuYLpBNJosFYd
chzW0XROK8Gli3/CEnr+LykhILgrPPXFqP+1No5zcbEG9cvfHYAWgpoS8bK/knQO
aWnvZxkNFgm+4+Oy3XfsIh7gqX3hfWbRG0AQMLMPMEY3fSpVsh3pTRoRl2J/VF4D
jNVxFS4dbJZdVfTFc9zsIJfZPQLpQyTpliOkKoNwk2TAV1pfLiKeDaUUX5qzXt/Z
yOWgGqSQlVYGlR62fWN+eqWNsIPs0ImrqZwHHjT2UateEDXFJaX79Uft/4BpvkQK
mpjyOgJQCrK6mp7QM1l3HVy1MDe+3tzx5PlzlUd9aHJ+cLGQsqGCyfdLiDR+/f9I
1zI81hkcPfl/BFFLq67KWwZGPbbD5eeTUDq4XKzgfU4lXX54pNPPFEIj58H4c8Fk
dbZV7zvdbolsiTodG6mztH1L1KoU3SodLOZ+2buBMr5X0uKJqxS4vzecigLTaZYu
+rmPyUGutDX9NLMrgIXq7/eYoQeKv+fyFBhgro+UCHiIhi+PcF/hjCvCsFrR4UKb
CRfMiQsagBnFItyzu63ZgnGNZ6ilf+fUc3tYA8M7vHDAMm5/DaHVvUZfMRNB6azs
AitzCxm6M3KbObScHMVx4lH86rVwN39X+dcXUn78XTfcb+bqceMukEp92DlwN9YR
xAP5M5qZUHx+Nb5NQSF+pEhDth+d4ovSD6aefNNFlkwkDIYc7xzI1s/9PVZQqEW9
YT42GmDBrJRi2PB1QXlRyqhA/Fw7wUP5ag7/9ajf5Ffu/xdXHqgCFs2x5oIUcA+J
FPujpAuJFnrTsFw6+l7tMC8UNcCcuROWleeBvau5H77ueORntycWng9iJbsI31st
XQ2RR3Yu5tRUw3xEkx9HgCixPX/EQhQEO/ylyCxCY9eIR/op6/gwWmuaySUA7DQJ
SCubQ0cs23BvU5Aih6xQDcxPUPamRtf5id4KB5ZNyKMZMx26erTxazJdZ//wikE3
0kqJhNPkB28vxXxwTyzxnjm5L9SOZuQmeEMKEw9+C+2zMz59M0X65Eokt1JlSSJC
SuiyEnD2FTmiOI1EWl3EgzLbrbNiM4GMlz7DkTyOg5vul+dSvturHgLoGbDB5bKB
SNlhMiUpbCiMwnCBIJ6G0Q3f2GrM4/O2EQFzxDWy4j0ww9yqiGgo0pLlc3+5EZM4
slaLX8v0uQzKr6H1g5f65Cprdrwc3fAG3x5xJIx+Y0IQXTZpMHsokjlu5Rzk523n
Z4r5YOiuMWsaQMu58xNHiP1C/zWDTKfCnIgpKy+Hw8uOXFAUDd8UUmRRYJJ61BEw
6YFU89e+W7PkYdxK+5shgyG6X5cU3cuzFFbnpbb6c2SV2hHVfHeiF8jKBVKUb4r7
A+lRRI6GpV+lGYEF0tZYgS1IV+f5PWExhJYgYz0SRxPFXds6YieZ70Xx4e6StH9M
Cyvgp7usu0uW5p2OfE/lpFZ4MP6gnQYU+YmWbYolFFdTwYh/7zVvm5Wm6Y5iydzl
zk2vfirZEVtsGJue2YRMVn79gzArgthFOFyrsAAt4A9WC1qTLFXrAs5GCpgEg447
BVCnJ15eVhzq8XOBCkUTt3dufuJ8Tpwjq5o6joOwuSKb7xsurdFKPRdoOSiB3E1t
DCXWy55kU5c5lkGutHH7sCYx0RLKAiC7fZJB+HxhJRPI1Nd9UIUt5i+mhzzrEZKv
ONrPPOezLJ9KrTYPR7vxIXYsz3UAC88CO9sTmr0ND8HwUOOAmE7xYIPflO5hq5it
d/EtR6bGWrOhXfny0RQIKlcJGgI62oWtRvo4GxxaX2DvnhvbDap9g4Q2cy/G9T5L
i4NcuCg+JeYCAuTb+xaP5OG8tDsew5Uc+v6ZZv/eoL8sluAeAXw737IyspxcfTW4
U5NP4VZw94sLZVMG5LsTxtXMa7ECtEB8nsFIlzQPBFqSF3jrXI5urBhKyA+iHz0P
rqTUnzbxkd+DtJ3EYoWu4S6hzwEHn4E8X5qJuHALmXYSd5ZxozYzAkfSNN0F7WN+
/3XVon0ZZy105juQ2VzS5jEytT5CZWBuG1SYq5DP8TxEBqdoJCrgCZs6Z8qEQnhA
kwaCNlp2PVWQgySTu5Os7dmZMKU0nprmE1OLep0iHn1wFuDVFTDEkle9sa2R5h2J
/B8FecMZSubTk+ukN1mUGvThOeuZvY4MaFswwjBNzKbCTD1tMjOewLSK7ERgsj54
z0WxM/5YIz4ZEBetw+bB12ye+YbYIfX7C8Bnt1wCcRfF09Wogz3gx3/Ge08HPDc+
Tg0z282eMlXfcM1PKoNce7ks7hhf8y6WP9hMBKodlgFuqnjIEvL2rzO32qSnUFOR
RmXkcajxfKzRBJx+5rEwEy6zlKcBgOfeHKG0sU0PDnjQKYFI1PaI/3K7aMszsHZl
p75SSoeAg90LPj2Wl0VBLaBcj8kYqIL8LqB9gVuMrBwxBAI7EIegNCiAXfxIqVKJ
a8ore9EiqzoGSnSoxcPScPsznFte5Ss8iE1M8LnNiCIKi6wy9yCTb2QVl2kHp31A
nfEzCpooTkUURE9tCmrnH1qdcBRB3PGaL49vZewTC1hgAT7hzR4DEmXtmtoKeIC3
t3azTBOcpf16Emc0zJrOafhIkuqGagVR2yIGJWIAwdT6by60+7zKerYJcw5kNkGO
Fusz3RRkQdG6fqC6Y7TyuUFSkCQ8KxIINHMJZkVh2r7wpw/1u9lAuA8yAEGDWvMa
Bfqucv+BjVnKiBz3g6sUkrsYeVoqA6Lse2kBnZtJpfC6TEiwWS6G7xK+tyYXTh32
1BWtehOOudnT5FX8vuj307gKEDi9VTTAHvnQUm/31QSJpSb70VPyudVDzY4HaSsv
FYBdXx8XNP5mwPjXagrtWYddaCDzubIVvMRhroA2yw1fubqL6FUc6LppXtG9PnGM
kBH2ZS05E053gYFI3PHU/n4/FUvh8ag0hLHwx29aI2eM8xtdO+FKqLIRQG4AaTvG
BGnDF0hluZPA2XeO/qjp27MLELWzNauR5jFK5HyNR6AGEWMk1K076pjaO0aUnHJk
pHsXOW3pNu4X9vRwVzuWgkvcl7TkNpEuik5YHEtELik/w7QAhgc50oKi5j8ycfkJ
YtYIgnqhEtHUWN61kOhVHrvia7spiKOc7Kzj9BaB1Vb0UOk3OB0cmwKECIzvbmF4
96IOq7F1v3YLylFjC2waw7x7TkIilsx8ypPAyW3xwKX1txx5ayKrKBv04de5Ehkf
SD9UaP9BRqYXUYHvzPaAhhAJ56N7PzHBjtDS9BdzS7WfY3t50aYukrJl4pK4+dyd
RJ3Dg06QTzwG2Nah0UuHNy5bhoZltKgQ4tX9qg7meELCCG1yWFtG+zUr7dokoyCK
Q++RUmEa50HVGxT1LfLX9eXw6aF2v67LLoPkaKNFZEGhB9Z75tLq+RqA4uXKpH2g
FZhSW4BnWH6gArJ+K+CHHdNnYjHYeWNmppTI5ajUiYKJRlW6KGW8ny1q/iVHUXwr
C/M912IdadUGHnLPxSQWFbng9Wi74iVleXFrbrNcUaJkAYDJpJMYIe1UQUXpMq7v
A33FdRndbjh3ceR9tKg5wrQbGILGTsPw/WmMt1SEzfa5X84twSo8m+/DXIcBSKN4
CiaLncCj/57jDUSlcj3PY5F4HNWhtEezvMYuPUr/uspHWSxAHh3f2ZUEIpBXQbx2
Aj7KBh4WfwsCiHi+e2W19v1hgPtNkovgdtr+uh/iRgo+VRlTfbDQLQ5Um+2C4iTw
y/FhI8A4r2347vzQQpaaW1WfkV3z1gCAVTzYXM7duV2YSfOxj2KT8VJPcSvYRTfH
b1L36uIr1xNZbSbyu6tr00D1xsN0iuyGpjSCXE14LGPGYHTWVa8ThjPAUJVdA5HZ
Kb++PHC1gZNn8CeEnkvCxPrvkY3fscnBxKRmcfJvCl1LasK3d/klU3zmDAbjReIS
/1BqioSCrZTg/A5xJtpqm58p1381Melqy32g9Tkj8isduyHbbdWvgUo6m+ndOhSb
izlCTTDRGC+6ljoTQ3BAtsLCVqDSW2u+PTZOnPqEr+L7nVapQon4z5aFLjvbYVpY
9P8GoM24pUDjPNLKJwt1AMiZfW4LuAUvJyxvZJICYcUxOlHvLEDLNrjCjLHBfqY9
03t3LyyV9IkYEvkpTDMusk/BwkgOf0Y+Gtg1eIxdYxVkh+k6A+NnnentBRv8r+99
oacuikorNR0ZHyA8Yv1pWyDIqIM1LV65ghrgVpPcKaEf+bREuwDz5ACRZ9vMD5Rm
+3RqILMYJEIiG/HejGU7pj9VHySjShP+PvzlcEh5G3HZXgSAhggWC7AXDXy2lEKG
XXMk/cH0NT8jHfBlo5vsxXPG7/l4NMwYDX+/DC1YqM8lf78X1rkwx2ribI2O/RNz
LFVGGON5/Cc9g1OxBkhD53Kvw0bTR3RQnWz5Tl8dLC2VbNIgXC5Xa7K27Oll33Re
HsxgoEUULzHZj5HPl07RQDiNvfBblBfiTtEhUJ82YTaXS2tzJfj1TgmVVYrvWiEb
ZMWYKWLVbusoKl+OiAJT4XziLY2is9OHktOcKJOMkamu8Z5kvlss9TPLMxdPkfo5
J+Rq/6DHA85GHkIWitCfQqn0fYZephKOtU8kR/FEPy4w+bfn6yqDNkb9kKp9posT
a1oMgWnJS/pjtLiNgnWFeIZ0asoVrqu8VtEeG2YJCghlgDuWr7rgnLSaNyuykqqQ
KqQIT+bSknMd2qC3a8uzyHxTFy6Ou9WsvAusvF/pxVcxRcvP0ATBM2TvFEqrYlXw
zZX8GFZcaKs+tk6nyGcyikuqWPHy2UXko2Ay0fhDic4CirghTr2dnBm8pv8ISGcH
SYi7b6SeyX+aByB7jSyC+0b2TNnEL2DNFU3QyRqYZriLUhaG1mZ7eQ4gDeewkisu
E8rF1JkiigCF5g99NQp0gl6nA0HHJ7AQtEfYsGpcFgjagBg+1tfOXp6mtgp+XlZl
7ISw2CmbySocXgOh0u212kA5dedbaBuhBcl9KdM3IPEzW05b2S4LypY7VS0RU3SI
X5KfbKvkGD83Ta9t5xvLgxgEtc9V/tY9fKgldHdtUtvNX5RQFrVnx2Yo2kXzJyPS
5Ho6M8AI1q+FxQkmnrSKl39smKvj1TQBkjsZVPbwaEE5vSKSQ8jezl71rr5yX7mQ
7csg8tjxUeIZcB0oAfpy+a977yj43RFbjWOS6zDnEtQTERTt2wtWEl5Uuu8Su0HF
xXQZbQ+iB3eASfypsZ/wGCWaDyINf4C5rzMxF8rarC4/8VV40sM4ODJHBqkcI7nl
JVNJFaqwhFcMLi5vpmHIXsrBmnBmbvNTn7TXEzVN4+/JLcneJ8xVui1TxpzY98Rp
RqgB4bKiFyr5lPfj8uK4dfnUVImWyeHVoCBqYWm9YLLnAhyJuOM43/ObCOBI7UHf
/1SOVQ3mBjDP2T64y87exXq6jkzPdQDQXBevJJ7RYNQLNKCCyqVp0jC5WtcxyCoc
lzY8QR0A+ukbD4DXIwlhPmjlj5BR2IYL/fL4hP33RCNr06xpEEXaWjQqldsaxgRp
BhiLD7gQAaZwyb0UxHtojOhzONkgReJdHL2ykm7lnvWvBXIs0BQySM26obWe6SvQ
G8l14IyvOamMq+Hw7VF+QgGq6359EhcP/1n6e3sVax6sOFgo9ggnXmorFKlMwEKd
LuNGubUbSvO7jGpYZ2At9W5hLrzj/G7zJQtRsTpeztxL3nf/lUL25XDh9mdHU3sR
Bm3NxZCQapUpH4yzMUGiFHo9AL0GVqF//Cy7ZXPswUEyIwbS9EX6n7bm5Bwubss4
6Z6ctlenn+JcpysUg7ta9WJ/tSXRJDm6FcFwrdx9wfe1iccXuJlf63Md1tuDmCH2
j4ByRYvxTFoO3WtcqseBE0M0/PLzR6HQKeazqDzBC7Pw1nAzQMjaD3VlRWfSaqB/
zfiSfcvGWCtFg1Mejil7CA3b54bRrX95mhRn/epsiJkZD9y0xGdMzf+PPUS5M9Eu
J5b6jRStUwt0fXyk1BnGFPT01cudbXkojbBADds8TjpSWFWpNf8KqzknVR+kbzUO
eaAgEE3XshsASIMsHc7JHLVpORM3a2X7Wdqy9zLkna2ycVnUViEHlScaNqgIj0n0
WzRpqjRAZesFZ6WlFgW/V6Tyte6ZPEvnLc2tZDw/H9MCFaPYTt4jip7qMyz3zbTU
8j8Z9ow2sd65BogxQFeIQ45kxAp3S/RV4523w5z4ufBOhuYUtrUKODVqXfvFhwT9
XCZL3bnuXMr+ezysp5/bokqcN0FjkwUW3c3Diakfs/GvBiMIMtbGhvgZ9uBLm4uw
jgCjhZLh4J9aV4WK84mF1h1T/JVNn/vvtsrkScbynGHIu7kxEnZCnFXYW0GsfuGL
LhcIRP6QXMM5RwSxJNGEZm9qjeICVkddmF5Blz229NEUi7OFm3gpdHUZoO41LtqB
SLrD/M6VFVQb72CSUN4/C4V5RNLoOQkX9zM9VZCzS5N5yVFhe4TC+v2wr0oGU7qa
GGyi6tlAquKcgCBcDS0xB1rVpGQhHds6RzfVKTTBBWi2XVR4THUrW3Jt49jE5Jpz
dGnZAAhOcl+3AVhGB3pRDhT9Jb4pVjMeQcZ5CIM46ijP63oxpmIiJAV6JNC1BSBI
p8SkLrR1vHOA50SI4G5ehksDqKm/LEbbE3xnr1BamxN/kesGladT5ntZc6Js5iQj
pjawY3e2HPBwhbyyoFcf7sydqglD3ynXleKt2XNMPZvZN31Sda3jZK6QKdkvQL6t
TkZS9WlrJ4zYiSiNnbHq44uazRzqFF3DzCG/5Gd0Yc4fiqayc15NiH46eKKg/oTq
WNfmKD3GX2YnQBEJPg5CWlwzr1QX1xL7wn3055KeyCWn8R1EkpYDTrq1PMmYEJSt
6OZZFSKOk26TrpGsnjQErY/ihJl/cMvQYHJZ80T6kLjHe2iGI+gDAZQZ4XDP9lwL
OEfb2Qdb70tv1VHIwf+qQDtSrpRaVdCCWE5ZDuquSrjtX1X6RTdXOq8Dr/ktrJ8c
8cC5GgD/jkjqNoUcXAvo3Me4VJav4O4rcpD6JrxoE51+eCz4CsVQbQHLZpqvQW4Q
3mTa4DdnmRgBBwH9OO07tIFiZtaCbsSiF+qXyjKtKRzkPjlb5h0i1uISaJeso0KJ
KCZSkAEyrt9g9ndN3JgmoNRmU36J3N84mhztRmN0CGyFWH6zpW6I9ecKCSfprk60
bAmuMqwQB5BUCBYavY4ANDo/yUdY/Ytu1JnZjlQQqP4RYDhm7JVq4tUXS+9Z2Evs
3+eIrRs/kU1wPMDKdSzz6AqS+ToIMBsCmQnLGLqjh/jBhh8/4mBkVm9T0hzhOvCS
BQNKVn3oR9efPret0Id3HGtsyobLRuSdvPrY4wGCHP8GtQHGPOlD5jU9cdxQSpVw
YuS5r1cu+EGBX5IuzdQJwSndd9N3QqIiEU6580dnMYOuuRgsV38en/fI2SNbHjX0
XDG78wG+z8qNDtsv5I50In21Fs4IaVYsj1OA9ickYr4mJjHpyLI9x4ou83FU6m3R
4F00SFdke3xhNx3DG+NNsDJEkH9ew6nlu8O0/MTMT2OBGs8/BAyD2wBCgi+qZNma
R+K6lQHyc47lV0kDfMqBT+TyMDQKh54SxQXXqG0ztoF4pMtudUgd6eVpK7Rk8VIi
ctoI4S8EhqNYWl88DgrnP5fPxLCUV42Jm7sJPQcw20AnigulfFw0L5AR44CG/FyT
xm/PiXhmPdi/ZuyOYJ957E0QX8MhTmd98G++v3OkxowKwEKPfLichR5rzFocRjev
2CakJXbASAVCZyPW4dgTOwe3P8Mh0vT7P3jaa42YOsR3Bucj7LCt3GSdszMRHMx9
46g7OPRoN38rTMo+xoHpyKfRB3Wk4WQEoAPeJZC1GyldvNxYAnKbF90hkfAWllGJ
eMTpA3vgcOz4ybA+gApFENYZJf+xZ0TtmZXxe4fKBGiyN6o7ic0gLtqa6yB17jpK
X1WraXlUZsjtfkWKVlhhcNrH6pGwWrfuc29Hv/vQG3sN/UoyY+PGNAx/K+khp6AB
cKADGic0i5eO/wMjnEHk1je+lA9FqXjkA5X6ReqfVhz54Ep8KmPBeQKrU/zisYkb
waXli5enq88H9u0lFnTyNYUTXvf4ROfEt9nITwCFm2Q/rhdlXv7WwgglVw6oX3Bd
L0iU0BN9v/GQADSMy2vuT099dARna2S21Q1BqOzxAGgQ8pc1BpMpj/AjGp8dBbhn
vOJBnwkt7Qc+JMjTBBP8mxB0p1sZBEyYV6aluBF+MDht2CGgNTa8XUOZHnrE5m9B
VzrT0ja0VQ4dJYiTsZp0Epty9yLDpaQVkQaiucxwdFWrkhARtkuExSZRdvrtjiCy
qvULirRP1gFlW2w+3Z9wRksWGmwsh4BgXDRq+IXcVHRMO/bqu5+BHCwLE64UT1/1
tNSSsAWVFBNr9SfsAmztFqKo3Du1X+BpLN5bOw3q+fKn6eBMubZZ68SB+Rcq9QWh
Y0LeUulM1ckOQDq/J8qiV4yNYbtWE1CD/CrB0BeknoH58kXUZp9cD1sW8WKSbF1X
mP4aRUR+3uKS2quguJTomLE5QH2bfxRGbN9AJfOMvekBikPrIjZU6RP9xtEOq38K
vDsEOZ+tpb7yXU7AMzYmnMWX5LAf9zW2PyBGNbX2ouTBwj7vzsOkbXsUh8VeXY+2
QqEQixx4zhitJirczldhCsGVcHT2xmOB4H9j1z5zSKsxbIkKuVJ9bagFYjuxr6yq
pvvObBoVnWadZqpJAMrz4QJp3gcZrzaeYr47kGT3L6wnKz+NEgXBIID7jOacM811
wC/S2lVU6jWwl13bSzUBq041/0d93CGGAUOT+6enR3vc4EkTJYYoqCSB2WsSD7Up
kmuxe64S4mSYj5UssJur7jhirhu+yy22R4U+M9yZWZL+KDGimAElwj6OoD72134u
F9VlxETRua7jpSDZM9/8GlORzGUitpcieB3J3bLA8Npb981yiD7eIyD1lOvVVhtR
4funx2agEpZhefftS1Lk7aB8dGxzh5CoZS1bPnULdAIFtSvf2sdt3DIM9zK4aAon
CJiUANzMNvrvKJSNDtmk5OIuQwfsTNr+63Bz4/xFr08xke0LQqMo2Lb8NJAcR7WI
NWlkQYYMGnz8Mxgz42thp2n1N1gQ0Hg3v8/yqQJQcHSHVJ3hug9i5x7jnVntDYJD
W/op0ON37QbIglAaQJD34cT5HMpG1z6smEpIVj74iuqdpk04+xTAa2mNrpagr88h
6QpQf92fLUKtalwHXLBjcqVssFe+m5RGx2KSrWtt0C8hxew5OfaR4nvZs/BZ1xY1
SPFELrKpZlDKtbboZe44nlGla3zhxvqWMOqNWnrUNXvCjxA0q0xeMNWrjYd5c4/O
fMFzrjZ8ZldCEB0PDuUXR0CLZGE4PvZmGMZ29VhCfNVHSUA7tx0+oUZnMrt0fcfb
RKsBNmIxTf5bm9teJtTUuoOrE4piuGVuTpn2YnQROtNpJktnuMmGtaNYE/z9ZnJN
EdLybJc6zY1m60lzopb4fv4AWVyLZXF6FFETlz0RX124REm9Iydjlf2srLCHB1Hl
sg8e5lj3a3bXNUqaUCE5Gi5Ct8RcwJMyGfFFljiw2xtDnYR4niamEFEWNMs31DA8
05ghS5IY2Nn4SZkMqANZtEaW36W7XPAZsq9OND0CBvYpeJOXDC1IdCeZUEMI4dAu
FKjSUdsksms/k9RBK/QrMDp5BmuV0lFUujteIqJXDsYTV0OYoeBTPDLFiI+kW112
qzNTZiO1/+VJfRZ2dHwg9gZvGZeISuDkuHL9nAPZ36959ntoo/oXsg9o0OJJSgy1
EWS8k1IWR6OFVUNK7fwMBYCd7+UJA0HauetZoxkqXv3iorLu4iEupfXU1z1QAHIU
GO566Dvbzn+NDd/cBWpw3G3sjWHXac6noh6eTjnZnuULWQNc0fLUJnA7rh7TySke
YOrNz4AEElrvv8PRaCGF/8LXXKyy9pQHf0PXVUHKfueNsc4LpAQvFwsnBohQnoU9
8BXwOob2Fk66NmQZqcO/zHoIHBVCNgl00UAoyDVvPe1tUvKHLwIAjbi2TyXrORhV
02CX4fZ+DP+Qemidt1WM38o0ZmXcIcN55N1m8+ckuUg0Dh35rE3wkMfN+k+MATLh
wO/4ybYEDx7l49c/7hNsvWoN+8d6r0sF+zt3HUExtC4qXJZcEQXzb3nQ2YR+RYC2
ztz7eSLfHID2BPkaai4LcTNEPvrS9ewLI03A4BbrrjLUJN2p9ltXarTjXWFYnGZ9
uyMrMBZqL60JWOAwpD0WlHeE9AFaruTGZtJFE58j8a1t4lNLqEe5L5bbFvkzFo8E
2VVYaC8kb+E94/JUh35mvQDmhAPk21nR8DfOOTtDL6UErSWkJ0jaysSJa+u1fTMz
xK+ENRTPwz5G7vzFNnJMDXbpqM6Cxa5Uc/w6uxEx1g5eKyAl5hyqXVvXWcXuPBTU
49ornP6sy2yAFb+vkT7mNozux5PZSW67RTVLo/v8EBQib2j4Ss++vxxR4U9L/72k
aL0vnt+zJKf8idub8D7X3tsk5lsb9YcPoEdPYD8eUnc7OABYN1LLB/MNDgh0LSn1
lAxPLSH4Po0gZjKh8NqtJXrBJsjP25ZrNBeqK7VUdMUMnTDkVM8klHStu1F5QND2
g9XkerEENOmBsKt7GeofgwRI3mCZmOej56WqjRFFxWcPNqZBUOFOK4NgIhgfvrUq
+Szzj4r28muzWl0U71zJBd7QfSDXkfrWASg4M94R6/CXXZ3Tg9FOZsW3+87BXEKp
t+lmQ5wg0nM15po63fW/qTtqsJHRxL+2N9YDM/w75+yd7rycCLG+mqZF5cq5cNdV
Jmzn9jkMnJDnep7I4F092xAUTkIhp4RULAv03pHcO4P6+zj8pwxdyLifCBK+EHD3
0+1tPTHU/MDAJYy5dMebzHHpz8zEV0JAHrYdnZmgFaAgsVxjZAkeAkMLDiKiW8CA
DfBeE917xDEnAaiHPVbBch3QAuvtPwu96NJ3zfsCnLHlnAKK77zOOcMy7YIiVpPg
FRyfaB4QWldNips56tCernOO1kvX9fhzAHYzM0bBvXYoxcfPEq6dlfdFZohJvN3G
9u3P4ec1745+UBZjWqDvJ7OxMiNcrUShaxgPzpxpmxtD95sCEdYcDKpo3nxgorxQ
qLRl3YeC/dAPEv3GPXkv6UxSSHbp8AVAKrQrgvsaHPIVUm/BclGz5fo6+KmZewl2
+HqCSn98heLPd+9IWW3gT/2T+IdSXxX3GXH19d4iHE+KYWxn+nfhw33tqu9qydxU
Ly9iDEByFOX3EzSA1xzS4vPds7Nb8/ETtfLZSq6bD4csx1i8niQsVoh/6hD1yomA
hRyc4UiBaainhccJxa3Qyo/rp6de/NyvkrIxRgBtkN60k65YRbnkT2ODce+EUNBj
0xkOOSbWO3V4cXcc1d4zwyLnGwC/OPRXufEK29AF5yvYXcsAn74gXAF1wjrEBeYl
EapEtr/UBAGSytVnC4s8OuNUDWL9F4EtRM8cYEj9tLFkH59iSJHNShcWMSgMXbHN
+KjGaFspxpLFtk4/C014x2ew9ejW/qgb0iu8de0j9hDJxCM5d66kNrmFCKMyvThU
UA/51U71eswVx2LSoq3FhGQxV2kbVVw2V7ALrNx6fTR4BKDiaXnmjBN8xu2XjdWT
GnofHt0XJXtsOlDkwdTpueT0n/393GNYAceU8eTQC8hdFzyDjAwS3WQUkCON9UtT
NNDrGa+t/RG4otEQGMp2My7Vpl21g+O9KopF0Hv7m9C2Pch7X8NqCtPBAqlGt5B7
UTZ1OiTchqjrBsr5ZIHy/Xd45deu0bDLCSztjqeIQceRMhPEXJCRpJAOrFoujYiV
lK89dFVwrOsWksaWzrnDqZby2dUP19h6uZ5eY4olGre/7pE2+7QyLVgSNUArKSzj
nTc3428PTOSj5g5IKfOZqIpL7sSLBcqJs/Ydoh6UePkqe/IrCs1nXzJVBKjEtZw4
VCazsbLu+LiriKFjNr/37JjprdS6AhiIANNvFQO+b1gVZtOsYWvf48KNFzm+G9rk
dev2pipkVqyVt8IQ77nf6m6u81Tk+e/+j7KGeHxaj96y71YOzcKGSWAnEWqc9Z8G
cKgmYsX9wC1Qk9HOuFY/LEiedRQZ9dHJF8Gye3irDzqansLQz3Pqyzokh21y7Hbc
rOYfGK5KUBKPTpRWFLPADi/xEbLbo4cN30syOPXrp4rLq6GhikFvtaKuGowuHbha
x3MrRR0p1bdFWOoBOV9HDqAyT1ZlUt9PqbbBcytRYTyUlskiO3gVmF2DtdbfmeWo
hG9WhTzb8Jop0y2/HxdqU7ydEHB6ih7c6W+XraqPDtOyfSFXoLEwOHN+IafdPQFO
5mdLlpmP8q1ZQetGPyECJMNjMmk0JjTET01W9eW75uEvtozXT3prisniEqX9lpVL
zj7BUH/cIcMKbTYq+aK+89zpghNUavwtwNiJ1kNMXZc6QsCCEhktj4y02fPbOk8Z
j2ftjPojUvTVv3nSTHs8o09vy9L/zFUuRT9BC70blSR6S7m6A2mzNOR10I9R/Rsy
GzY9pabebQAGhq3ipiz3lneNxXLfOgHEr+oH/db+bR7bhItIo4AIk4HzpwbQGsBF
+LJz3bVYv+0UUbdzywInOxLcbXFlm7hNh2EQ2WJezJsA8ULUz31t5f2YglbdXE+v
PhrimSukvB394FY7O4d809WclnQ6AUzeVQBfdncUqrV6yOoEHaratId0YT/OTw5w
P+IoP1/fAd6OjyJ48A4F1gtGHdKr9+YrS6NOotHeZjEVjqerSyeQH3aygn78zWBD
ifG0vYizxJOGKSyHpXmN1Z/G0N+ShykXIS9tX5kNOv/F9wlmxM+Hqd/VAtM3KexH
5Tl+BwjGMDkzWisk42SZCk0X7BbiVYiUx3PXP8qx7Ko2MmSjK0bAx0g16W7aa5wb
TMYqBaIdzzeP1RnzKMLPk6x+Ti8HjT/eLQ0dfXt+KKByLzafa9rY9D05SZ3OOzzt
NGfFaVqVaYH5J2l52Vg64VviEbvV/Y6UhPP2xDbNAGYWERuCdqtp08Tuw2kND5XX
chAqqaUkMLFe/aHHnOr1fZpICd6QVqDpAVKxaUUt+H/qKpjXoOVte3JlXlDihlT8
OEnMULHSe/cmCm1DSa+BXNSXMdlnp2IhbqhX69aw5HBJPiD9O2726Azx/q+VEQ6C
806PwoIv6AbPacPISRJ0CTIPEy7opY1niQTgChLM35PKjkUndRWNKiFZLhMvd65h
oOOuzlVQ+kYigmzNnwzs1xvHKT/1DHGI3zZHvgPtjyZgH6i7UDITbpCOeTdmBKfA
L3VdYY4Uq5xCSB3EmlEtj25gHWgEv6TUot6tB3eYOHpCmayOL82cf3R6XhONL7ph
fwigK1QQ47sXr5ezBT7dpn4jIaTnCYJlBsFM5tbRhxPM8KFdBkLl0j8lEllQ93iP
+I/X/hSlgIdPCIA2e6RNEJbt5LY1WCEd60QEMaYtDQmaDdnGJOYdPWxaAPYNYT72
7U6XqjqADZMHeqPuJpKkGKba/YumlDIR89FvGKHBOOs/eAFzvjf/YaVfMIlNzmbJ
wj+EaJ1hcBXd2R2c8fGbnTUPGQv8hUnigJ3kwybcAjgSaWqj1/MFkp8J532Sw9Lg
pGPX1l9tZtQCPnAG07LcWEvlHzhSn2X3XjLP8Z85b2U+7qFHSVTw8QUSlZXSPxC5
ISFk3zSAmtWuMwGDCZXH0IlGnVXLDoFKmMqo1gaXJcjd/jlvBDZHieB/AFUNxidu
AcD0Ao+fKpOo3OYYizjSnw6smsgeTA7bh2r1/qTFZViKEBj2HRgduPnF0LCoO9iG
rj+emb0CtYrx0pnCgIKOxuLV6R9Lt/ZXGfV4VhNbKiHuHEXXZLNNfkpOJ/qyThTi
CmNJw7BGIbkh3u2VdPEcsCj3I/Loel8sXAUX2B4B0Nu3Dl59/zwDOodtfTjTwk4w
28Hh3CrDGbMwqEOMBmaB14sZAM7uP+1ju4xYnwa91xn2SucXuZtSSsuhdxKwXiW8
5FkAmQtHuGjzOO2/0lAkldxaMTtjtBkymQ5+sc/+rkuWn/Zqa3V/CQdVuvURWG7P
FYLMXShdDnZ8jJ2uZwh6vH9MB4opTTSbNrfn2kP8kjgnqT9gKaZ+0i+1x3mgMueH
YzcbMX9ESmZ4fsR5I/sg9/FoBztMk1huYBogsKpCZBrb72wBl+zHc/43cjc+KobQ
uwFXb/+PGjuHSrMiCXHalJg1s+euFDhvH/Kjy4ZwNvpPVjuJmHRYC9KJe0u3OWA4
eb5McYbBW5f6w5c6JuaVPKWKP95hV6tFuAJ0Iwr0pE0rLRtnrd9Xb2NRqvXLzls7
Xdx43JCdv9yy3Dzcp3P76bcA0qM5RNWT2ieJ5/fl+3h7BU0swXp6iFNz7R/MUftn
znXG62zTNOzcMqT/E5+Di+d9VjqM2NfoEfxFhSBR1qfUiopgXb732zwQSsZuyHMs
kKX3ThcsJUjBp2F0h3YMfoGUiJd3Wc1hT9vn8V09O1zatZpMKSwzG5CWG5A3pweq
k2XjKph6P5sNEwKhmsJQFCz8QuShlE47WhOCkSozMfRZQhsAz2BdPYTWvcBq5TkO
yo5lIxV4Le/c1V0pD9Eaa5/0PrE0iWDnf6DtrnipniDMNXClWETR+dsNqd2U7SMH
x1rrcpGPR/OghpOTXpJ3g/MSmtESJ5WW882j3NPSoOSdquhUVyNq1Y734X8nqWtN
1b0zaOVUVd5xjxRQsxFfMioLwQ81+9/7B5jFprOomZXMDRwlQqqYHXXxkoAdl/bJ
34LrUOYLKdhPbIEpdlJAMSA155KKrY8eTfHhpvVX8qqNwyIqrBIBmwOCwtFLbKpn
I1Gw8bQtQ0TvqlWtJtLIu5S42u0Z91YQGDlE/wfk9sthRTYa5FNvULIISXwbepXY
OFVUGWgiywpY8l2Y3MmgxKoxFZuDhRwZgYVDmc+/3fXsEkXrm6j292gA6dqo9AEa
2c5lU8ncAyLLgTO7PO9VkHF46yQFObAZGbqQgfMKlQyOjS4g792tJDqrQAzN/RXd
B2SBpmxqp6R1YOL+67ZP8v0hiIvSomDU6NgZKAmAaMCnQFBqRSJSfIjVIlYtHZRF
RrM4UC0C4jIAlldsUprnUcPNb1AxRuMR2a7F24CIBcUQzYCAws8tUogdeKAKb1VQ
vMOlZo0aN1eXFywi5Bf7rqAMDNUYrhcjJatLc57T1SN3Us3lZkN3xMZMrtPHznYu
si3xAMNaOfH/YtsuJ7ovWYAHRdo/5daqlpMHZFVQSCeZhXR/Ss9XIufuA4ILElxV
yd8O+gagFJfTxED19He0tOVVJTfnJ4mIMtu8cCkaksa/Hwty9wdoRLgEzgA5KImI
EWiADLwRYDkYrVk2gegNacvMnNrKLAJHFInxk/CNsjUQ4kU+H8lR5uhF27vq99OI
vmT8BBlOr5csBKsuz/F69puLgKmYWGHO+h7DLq9sgn5WQy8faxlF5uprueus+c1i
FlOrMZOqFgm/7L/po9g+g+UiZH4aBwRg/TIQVF80dRl3F1HeXHe5R8+nXpN+9jbc
3Sp5yZsszDKBpifj7FXi25PCnCxTScgY4i1GbyGiHOUG0wlCcUcUJVX5cTUnrKAk
uSrgRkwjrazc3sqWCPnjuLlSsewCxQseuWl0Tl0vFrY8LLopKatTY59EMgRa+SI2
kfTn3AIqn0ywLoQy9cVubE2JrWkBARCMTLY1iapbzcTI+wRGNSa0lUt6EbzYWAe7
7sqsVwICqCcs+kClPr00Ubyqh5bjy43dsrLWDpUm9qLkg6MLBl0Fec9JIiccc+ZF
wYouClJx7bnK7Kffl4gTWAaUDTYJIvBLf/GCjlKVUaljoQ5GprCDMNZhah/PYryE
h0+UYFgrE4GW/d090VPgdO3p7NY5Ll1wExIOgo+aylxkmtB/RBu5BmUDetxbRP8E
JsjCHKCZpcZFJFK+kHVnQ4/fY2esOxjd6LpqE1VKqWZPMEbf8rEESCiiuahma6Xz
4XV68wIwqkaUNdoTmyisthhdUmEHTECHQWCfunsVbETg9MkMUVYxxNGCLA9uw9cG
AtcfNrP66p1w0Jhb1QKgSDfiKLXzdzjXh0LwK2I/sXAbWziLsSXypZFBzcDz6K4k
x0dj+1s5GM2GAaQQ4WNhmch2WdpDpS4RawurERUOZhLvMCtNPtxhY8g+ooJnjO1B
3QHWBu2BP3B3uA+qca4ogLPgYv1muWMJHSnw+zU05YLUPTQhOp+MH95uLQklw/+m
7uG0YjBgmS7k60dDL/Y2kBS3GYzExTIFTrqkztaA+hCMsgx1wymDyUEOv4aN1zLf
qWhKsbgbxLlN2ArZRXOH+rAku2QJIn0rn4HDtMQadjK1nGHhlFCNq3/0dxtIk/2C
6QCV1upXHSaTTDC11dbRjrnVQBOJpQManpZTpacpZCqUDJeAAaLBvetl0e0Ud38S
66NhRJViMaZwrg4ONvuwKs/XdPCCy/b5Lnx/jmaJM+7rsPlb1OvTuETHTHyitZN0
P3qPf6AHHgY23H8afwfuJ1lRGmn19vGGzRxczqK2n6HJ4pQ72n/RUAoYDA5tzvD1
0ODukYoAZpA/tJ4ckGGVMyvmJYioKQibxcyKPHCDkDcz/mwEwONg2m44/pF3hzK2
gPbRHmOdy7vG8sw4pB1ufd8za7YdubFhlfBVw664Vl06om3qvNDFNvNvKCxAP4r6
RNIM2fDo0Rbmo9GE/0zwtRIZqwSkuJQUfN1TlcENHS2VbeDPhGTYdWkgOrzr6peO
1aoGZKnzbGyU2I7hz6yqqXwXWQHW5A1CZJlfymEvhfc2oDmzJ5oS0chSANz+qvt7
6ST5ZrQMVa+AOgT98muMx81EOBu/KavULYpij56WXAyelr5+6xFRuMx7PVwrrsR+
fq+tGutwX4xZuTYE4Udy4J+y+/UC8uwqW2Hg/hM2YL9EMYde/FgZLY8Nvw3vz5kk
V+dLWdby+Vw7LZ++rfse2bzPb7ckvu6KE+ajfpfDum9a17pIg5asrvzaeT7E1SLl
CNgrpohaUG3ktApjhRLqi+n07n7gn3ALOD23dJ/y8izK8nSitUWfJhV+vPivMv9j
qOJKrVjJsG/LYHVUvzWYnVsIH/vY1bBDZJR1/YQleTk98ej8hOuaLVFcHfEz4Spv
gaQykLAi4WunX56GwoXfVYxVH0+vRrje5bwtAohA05o0blSxm8XEmldCw17jITpy
sZCjRrEMLdDKM5oEfjZ8lTOki4iEqQpwGPfscmkuM2Z0TP6ftAGqqTg3ATiAheJ1
yD3OW1FpBNXXkFs7XyaG+WjFgpcut5k9DbDX0JzAwF41iWIWzOHu6rlndiOdJYVh
gIlIqS5v0aknkNiB3/9KzglKbTo4L0TRdda384JuwIfiCWrTkqBkAztzVwRqBKOV
SiicOI0rhkpASuHYjwcpy3CHvd2apgVvl1r3YFASkVsSYtIZECX+sNEAVUEvbLv/
iyzbnNCdHgLSMcCMzZAZY6jjzvWqq8YsN6pL9nmXHk7UdeB74RXpWcFoeMSIwj/W
7PTFdXg/c6Ljg1rxHu1cM6B5CldISUasD3J7x5Miz0pwZG2xPzaHFnxOngeBu9wo
gR/MC7yDRis6biYKQQNokRzIPXFKeGwudp5O5UGjmjI/wK6IjHTob9qOZk9bF1RP
/PSqFE+lTeUwB0T/gGDb46q+mNCLeoyU38GBhyS7GUM8K6vDz6bUflsdZkdBv1gc
HYPgZETLSFdEHRHYXjyq1oUkQi7R348IscIYulfnXQUb5MqEdgd2nwLRXOs7P+2H
snIceN6t8UxwlY/MZo4+P98XmdIfvBcWudXId4lEmrpscxwu4pq70HlGvitC8IKQ
V1DGTKLCY4LhAQnZtE2jfnQRkgvtG6atUxwB0rhaxPhfINvKhOWnL0LHTBq1HUZL
EORTgwJREgwKCPCqfKNJ9YXBDA54t4D4WCuLfoXLlM6V/CzlCday651XtwUd4B3Z
gcmTsGmbLkBIdhLz1oI14PWVEPxAppoYtQc1iXHvm9R9BwhMk9XHOePpkAdj8jKq
pB+iNLRwVANQnwuvTHHpGz+ksw1CiOVD2UO6H1nGea02InhVAlzBJxNg16DLMGLH
fSlmnfVjK8wJSxJYCXdxfDwIBFYmKEiHFaURaWj4DSf60/a1luFIne+Bw5NQmnKK
7QuuvDGRqWw+HzEx14mDSrmswoZwDTLspoO8gnulbqpf9MHbvJcxWsr21JPRaZuU
7ZbLTv8PJ4O5D325Yiudax2Px0ln4OsDYwnKUOdoYzKk+MqOcHTu39IBkXhPGFca
qxSHAw7fOmqzkfOBkxfvixKOxQCkPiaJ6cICYkOCmyx1XPE9YEsq9Jm7pdidvDX6
njQ1+zpAXF15soFDnbdrpeZ7Dco7NYrijpZtzd00baTWM24mWY+rBsSTlwkmSiPe
VkvjWgPU8SdlyGZNsC/dLVqvDNAoONVD8zcZ5WYSlwC0LMsGUwc9etpED5Bm33Qa
Et1YcqKMfgJfDAr+5uZjWtjBB1vB07wIJ94cci8Bz9I70BqO4V2xTlZ+rTm2gcOs
4vKRrE7VVLyImvQ7al7hbANAVZJkxUvO24+P+R2YL5Rl6hGLtht0vGiInrM4owmJ
taGewioMIXnb+Z5Tg2VCc/M5JR7lGJ/zzEMVrGaR2+/AewpEhlIQEPZLjT4ntZ22
8XrEWDYrGkBBPBR9I1+Hi1kMv+pIIxMs06FsmpXSbpsg1uPFuGlTfi4SZfeMouLg
Od85Bz7UqviP/J+SysloKorNm0a0MeY4EmkdywcNrCW9/41qDNDo7IB/S37hHSQ+
NEeP77Kgty2eaLRogjw314PhMlDwaosbx4oGju2iGZg7jUd/CycubGR+BYLGEuyh
C3pFTzmu6yTxN32W9YoCE/nbyQwndqp4t9t3ODp9dApij4ikxAXQ0h6v6zg/lLQ/
HScsSHwL0RfQEVbeNhhu+h9aW7hK99R6+pkWrLJhxNXqVO+gizdsT7yf0CBrkDZP
0HzZUQBHCzaKZsF01ATHc6/RWziq5qsuuZ8JQ6N9ssYcXPpr/6s5Y0464mxGksaZ
krYAyXnd5GtX/9r7/1B+3He9/0qjdaeVCUt43ILj+5EXF1JnkunA8+BCqm77Z+ym
Bc5isV4NdMhdtmzaxbHbavAq8utSqgat10528seRGUksxwbvYVjW7Dlk+3s77rH/
oEIvFtOySkrcneJRNKtGmHtvorjYFoQu82grpEg3pWo51jwnSPCdrq0pH4hyFtTm
7DQuPgrRLtwoqU8/nEvLF/e3FvdC0Me1Mta4vQf6+6XkZuttPyo9NKOCJcM95aPq
vuAm9dm/a1og6BEWCEKcbHNmYCyd46ZrQdkMNJ7l51X5IT+aYrkJfFb6yd2q6Uz9
SvtRlUNyVvyY2IdOIQSstjQ5MjyMW0UnBq1TK9cic1fNrS8gkFuLNjJEOyhtikdf
oBs34X/ojHYoL63x+HP6zupP073gZCCa7HmPMfKbqtuQW6/P/ykCysO8IvEYJtyt
loskcR02sX3fn1OxOeYPERKEd0ZPjQ5JFLS/s5T/xvwdCiOkJuPLKNxt5oMpgmQL
OO+irkbIDjuyYvc5SGzVbo3xArHNnZP3mbXGJ3ibXFb/PQ/Xr2VwlD/eyhpEj0FW
TK1uXgoU5COnkJqhzrRyoAgcqOg2s6P8R7xWTu3f3UBKYFmTl0XnaFb/mWosBRQq
KPwCIRwbh0jQehl9Z2QPzN5NjBnrLYfyfUYYdHlWza9EgnjtiSstaUwLIOxuMpe/
8v4QoQtVegBkG0nNFXzQTRSYGPdIHCNxDy2mcgPcKzdyrdey0kobt9zgieXHu1Fp
6cGCEzpAJ6F1dwe9qTVWZMwPfJNZr9vQWgeOi3mhIdZ6IvqoUl6PRyZsCb41oHOe
NSKQyRRFEtEmC006g6HtwCb6VM9LEc10kKLW2tx4wMFJYs2ARCqq8gvw3WWeYtea
dXVegCbXIYyiR+SuHeiHJCSZ5hHe2UyX08p5WLdSCs+Ecd/gzALYj9YnC18PIZRm
Y9AnTYHmJj9BKlG4Nzj4ArxhWFfnj03I6jONw0Mznft8DFCZtmpKOad/nTpZ45h+
VauL54yerqnJB6B34HSNG2FCZMjNiMUjdlaShdACBaz32O3fOxRUZ6/3GxsPgskt
duaUL/HhA2WLHW1Gs8gm0VkycfjUw9j79QPdWCvVnpcGmq5BMEalPFx9QoUHmvfa
EIkslRXPEdEsJIagoN7K/Ctr6KB8zzx14dcmegUg+XR+nVLdOG30Ec9WH6hjC3FR
+ujzEk3amCxMsUqLXAjVm3+xHeidP31DaFMFlAb3rCoyUu65mA8uOK5muES4o98M
S6/LIMkT+82kh5J/XRCHTKc6UhgpxSy11jcTpi2LMZkeOVGSWOunau8H5IBQul7n
yksEQfGwrFA+u4pzXgcfq78RGxrlkKvo4sMCGmUDP+XbN+roXtyeaQiSPcK14qzR
JMI+kZ0iPYB7LBqFJqlAblD7Y3muL2YCECcufYwX2lZkX6TW00EWLNwStxuBIZUG
yqLH0HzVXq51zFXGsxyvfgzn6wU5VMkmUoORVoiPK3mY04Ll5L+5/d74uhNibXIw
bYNh88s5Ol7F4PjV88Buoj+dWiAYRz5zw426AMOr60IW79NHtc4p7cav2IEJ9VE5
UFU2o1z9aOrWAv4qf1G+ns+thxBNLY30Ptq5wKQZdQJn08yWzyY84WZtLtZGot2F
negfpHcpjsGa5x4BhhZlXsvwVErp7Ra8GnxNa/3qtWS6xNoZWv7gk+M0HV7lA9oA
YWgKrY4oUvPyBVHerkL4m6ADzcWg2Gj2hy3EhDYfgEHOoinAyUyC92wbSxjc8JPJ
Vti0NlsOA8XLcyETJE/3NDm/FYuBMGaJ8yQYufELnt6QtmOAbPjZGqEae4mJt2Q9
7YWgbu9fp92y+DwtyZCC2gXvP62++yLyje03ff2N7wAnTCGQgCzdD8uHRHiPouwJ
KfnNg2asfWiOdDRCyvfHMmX4C4dCcE38eopDyUpNqtDdIeYJHW1s5pXGtrQnPBIt
Y5Y7iyRAFzXrW/VbVP61bF2pDMF04lyR3oqJJ+njFWWp5qT0ufrHdidG+qxhQo8Y
LTiTolFdxBiTn0NgHODVANb73t+YWV/1jwGfD71gwaNYVwn9bHtxGBFipvQbjkoJ
oIBazGzhZsHQw4AUkzVU6zR95NYNXcioO87XUMOWaXAd3nOh6ZEOo9ZaSIVnv+V+
AMhJgCL3ebEBYNnpa8Fwd4yfrfGbVw5FmKLP14IXXAKSmroSvw58gla+UB021xTP
SUZ9SpcDycQ3CnmpMYJ6MjbH29SqYPA0EwiKJ9UEPoi0bDUBP/kYUDNcIc7zwFLb
t0/z5gp8LZzP8IMjqqVn2PpfhDXYf0ZMmTsU4nMGut9nwL+6invCgrVc5iqq1xVE
Fi88QbqohF+NBSJzA5It+d5ksVYHU1MctceREWRzF8qoB5isqKZeUAwfUNeHz5Ax
FnE7aQ/G8YqrtR4k4q48G8jmQ7GymiHlWVYVVN5FxlNyMjdCJeodpJ945uMKfIh6
Pu8xqndcFo72xG3I96hoHX1/DNpBAcU4xYn6cVUqNTeZk/5wBooBkHnjHYvM1H5G
/yzbwuFC8DvZCcGzB0z2RdevfA2Wp89i+ZXkk/fmRQ7xeZc/aTcgxYFx8h0EgqXm
bMFff+ymHooTcIuOufAaq4YZvJQxOG0gw4kqIQaV9J5JezOXL+rirBewADISTV6i
tU2q6aKTaMUR00Ae+/jqLoLbpfYQNhNswxuOv2+f631Rx1HEG41Z1lkUkKkbgQzQ
RUjAWHFfJBwfngsjn9waI+FtEKO/TiF9ebg+Jtks4u42H65suh2aVObsvMsCfopu
9OKFciyL2TDteJQhnqd1xQbBBiISsLndvZ0YeKbpB1zJBTjokg52ffQaimZ8LemF
1Hfg+yyaODjwMfr4BC1OE2XjOujfb9IcxHkviK+CBxEhhOmkuptA6hzi/TcMHd9k
DeCuSoyUgcdP5zoK0GSvsu1Zq8gydMdcewUVrwB8j0COkHQlXBmVHgdbnSerlh8T
gyLdgzlJR4SWZ5iZJgoSQG6B+WdWkOHYi+IHy2f9KipEPO2zKv58tKbQEWAJB+AQ
V0Yr8jw+fXlmcxqVvUS/pquclNI/XB1b8hyLii7woBU985PMIcq+9JcFDytNzvIo
aVY3jFQlkZYROtzZlBO4z8Rnai0Uauq1xq7OFbbZetoKv9ab4ltWGpJKhdyz0wHn
XdJyx3/pVSrR/l0xjNgguhD6EjBzzlKBNuxWV+ehziwSLI1UmAjoG9IGaivI1e3X
2D1CaDdjzpNyy9jBY2ROf27cEw/btgp4/zX16BPp0GV/ao94HyzkZNEdXp8yc4t+
Tmko0jZ8w0i1hmOZFCTmNKZelV8iuCNpwhXYeaYFKrT69nlTSelQe45UMWPRL4pf
S0aMxDbN2t7gGhACrgVY4sDwCiRdOxLbXhuC5Baw1FH8QPj3T0OVT1uh7fwT6j4s
LD5W+3IVhLpnbs5fEc3k5JSSDcePGVgTs+JCjqh+u5kbYWTAjXtzrzCuaOtrdbmO
AxAknLb+OysJ1IKFHUqO/HliEY3diy1V6QWqagxcoDPNX89PzyS49PRSrrpFtYNu
quLCUQrM/m+23WEjeBPHkQ+ZbOJlyTmwOucben1iw8yvB/LDLF7oX+hyD59scC/I
z24VeA2EIgFjfVLDvmis30vTwq6HvvVO7M6OVM8G8nz+O2nppddgVhWSCqj0G4J5
BKMrRxRqBC5beWgOsX0QsVty9/r2Eh+KdRx8Dzsu7HteF0XWFPocbKWt8F4ScnAt
4/x+02wOFxdWG+a/DD56HDEcKDkmtq0OcR9nmNLsmvR3OUnTJ+QJ4D8s8gHjsNHZ
pEZO07wrf0C77HATyN4GzcxXjzdRFxQNyw+g02oBcq8kkAJWTRM4DSC7J/rSdvAJ
gZ+5FPfOy8g4OHXlvb/MIDg660ej7x1jDfes54KQqEHMRy6hwUDCD/k33zduGE6K
5BK6QHNdUeCHvFNevfbi50qhBiDnSTh5Y+0AksCFz4g0T+h9hmrywytkViPSfRHC
Gvs6SOoAHm6SPHFJL6UVoZZq6NPFy9gKz0XdG56PoRCxKdrSfNQ7SuJKtjesOJcw
c/VctnmwJhjy1K4puiO5W6mXKa0FIPpGcZ7CGGUy0/0yPdh1r9SEDXkvZm4ZC3sm
r239QHXhZmttaNXGl4aHPNZx41zrMwndv/GndLBmlDdF0j6tM2M0eJr//esBNY8i
bRCr8czXVyZCDikcOU14f2otb9FJKBmzM5peGzNq+j4Hv1jFfAUL8XHWsPK4xQTB
OoSiylzp5uiApAQCl8mdcvP/66AnmKZcas1icEPaurBefJ75KqGCSCj4IwAD6da7
Ucwcun8wR7667xieu37NYwPC5Tgsj4UCMuAyZFl9YDtpcy+K6Y5d4IBHAxZen8BA
Rk9RoJN1XLdHT17w1hDyl3EexCFcMGnQ+Wvu5UP6nNnWsVJ80KCQhC0yGXxPylnV
pERXBVDmEmQ6q/Y9CbSj9DH3dZy08U/IJOrOhAk59DA/WnxYrCgdblxz6L9CdOa8
fd+ZLzK4vWSyBg8RKsrVHn6A7x1cAM8NP/qZ9IpJuhVFHeiBQKmewXUK5YmhpJNK
Ky/9yF8mBFbEAk32zeV+PX+7vPPRho4s67vQiAUoPnlZUHuREtJfYVrXWL6rGxm2
rFwA19nx0l9CSgdBYIInhZB7ZtaugqMIybT8CPaDZ7YvsR3X76iVNrZLVSekhn6K
HLW7NSUviO6gM+kPdxTfJmcJyhQq0DYs9UXO9T3KZN4IDxn4+k6/OsqM6w46NQa+
wtlvsgF+SoHXUrK4Txo/WLQDcgAyIllVS1YXUrr3szaN9S5agUTYP5wgDU4LPTl8
vwECOKgVlh3c+VP5Yg0Fkzeaea4mS3m70okPAZe23sonpLD6TZENKmTrDUHaAhpL
pu1ARLS+PC2qKEA/otMJKj4nij1J8Vixmsqf9tOJXkgKQb0tgArp2/Hw9cu7Umv3
Bl9uWNpvmkJV6exWFqfzgAw+Ok3ImjfavCNMdxnkqf7FpOY8sHUusvNLyDC7wewW
eUUqv+qaLpyCs0RspGYxSgDU7p67FI8GHn6z90CdQ88uyvNjnCv4wKQ8qBdIjUVK
32uouZL0HTBcmCI0hQW/j2u9E/rwdFMW5rdGS57/j9dRZwQyTHvaRRKGgtvy8QIg
0+++u96Ps6DoH89N/bSzOqNjPTVAjJl/ljOfJaciow0qB2J12mSy09pqj9rQoE3x
JeXrMY8ccc9sqMOAVMegMoYcfnevG4TRQAy5UI5yVTS/9hxwvPamQOtjK1WKVEjK
SsETWjDroO+bR9hrw9qf5KbaUBVzG4JlEwmqkRDJXlntrqWvYPrs4vXlESDj22gC
AasHHaFwOcjAiuZc3odjKU8m01ruHy/7ufGiHjEmYzdQMQrQHqnrjSLk0wyAI0XT
Dxqxqw6FpR8V7QZ6yi8A+YVSvxLlIZ8m+Mitp5nrmtGPDBXoHNPutaWd+KCCL3+i
o/pMnJ9vhbI60W38rR0SdJTWJHFgOMoH+HAMdKMsmJDOj8uBB+FctsCe7ecy8dky
Dk5+1CVMzkcwREQz2qCoY+tz7jPU3uHfhLgjEpe2nyhmemSeB9Rg9aYsauGW5lLq
uFwDIBpJ+hKYUjlYN3B+/y1LhYPuiLiL+QgMfn8bIxJCF9ubwCz9S6oLHmQ4deWQ
HO2U2W/pVGmXe8+28MpVwGvlS0HoAplEGvNuLs6DxGcfOfBcLcL3Ali2ctu1FppI
Il84HCwDoQs1hLZue0f6U5TJwHmJJZ0pX7FP6UbEkJaMkeWhQVELf6Yjcs4Nl8cq
irevOwnX4cTHdOw+Ga7ZW/G9983A2uxXzzFjTmhToIrk3F4yaHeJmbs+oNNW66fZ
hl+fxodypkljEuqkouuKL+Jo3VeG9Evx578uQhzKzsBBw/gaMNUiEMOdZ10+1qEO
SZTtCLiz0jBcD3Ob5swVqRWYW09qtCu1ZU6RHLLqX/+c978l6T4pX1yJG9Ik1qie
UXETccQ9Ku5ZAGOU8wHrNnBmk2Y5a+OvBiGMdlMafvjE0d0uySdu8vf8r7ohQqEK
DWhoqoI1ms0ff79XvoIM4JAx8vMeCDV6mDeD40PumsX1lb3Jhge7k/ibQyxCHIHK
6iWS7034yYaCm4yyNbLSVLZatyKW6/yQ6jfYHs+IrAwV5vy4IXEsn/+JIylOVOVA
krwsvlHlKgJTXRx8czYsgkUFjRrTqtZJkjKEI7J9JaOj00WucgZluVkiVmHh2V0j
f0rGBrynjgcsDzaEWRLMmN44SGWINiXbwNdIKkcti9lSTzL6qlTBDxjPIWg3a+G/
UcwTLPorTb3I9LGkJMrWEEXdFjCRjfP0JgS/OyGbI5xhhMODThioeV+eBF614vBh
kdS+zVy/ihoaLlhzmP3mdlyywtpzLRY5TOxUzDMBOcoxuJwYiFzhbZEhjLPA0BFd
s0nR1Mbh4eh10EN1r1W0VRUJwYLCvlmctLe1dRIox+FTjVJvV0AAF5VC74B47TtI
j9xE8TAF6xw12xEeQMsL5/F6k/SXm4nheahdWC5FtgrCBq9R2snkfBsVr+Ka18PT
IWVEIeC0sMqFZT2MEsaoMh8ws/8Lz4MWtsN3yKNEe6LU0B/c+PTrPCKdpMqnfSIf
PMjOjKuOCdoHhYzkpkTgCIlbK80dFQw3ruRbSm30YMA5hvyOnxOrUyXwRxSc1UeW
skvIcOtupQoeLBKAilxIZ/JM7D3V+yf/2nmgj/97m+7lRLI5RJbeAKGyTWDsmCjd
fqPc9XINegTWBuPrrWDVUtTiSqjP2HRYdyPcSoptI8uVDHiXWkuxyT4Mv/MCD0t+
E4IymawxxIa6yZYNv8xGgiEMrBsLyJ/mO6rSmMCL74xic41AxPrcDtxZAwJx2fbh
5IjfCFWDlOx/O94HUdXX4VZWcXyk0gz25MujFGawoKAea1zuW5aAI8ESSpGd1tnJ
ksm4DjW5PU1IjnnkTHSOufrAdQQhcgdxbHO1gN73Zn1IKdDAFf+/fG1k62fqFgXK
aTe0QY9BLC+QmNKn13Vq37oMODnlzRQc6ed7XVMf8AzykEdWjGmMoosvXWGK5PHw
GU60iMlWmM9R1Fabgn2PgNV992w6UjtH6N/Fpz6sKk5x+WVyILLvpmpggTpovsoA
AMjR+d6RrxM+hAUcVuomGdPgTt8CjZ9kV/+raRSYy7MTYU9tu7BT2IPWjHKbsdsO
r1JnJ2CiPfCsVpidAKNVQiih8ky9DZAkcI5fRSdqKsSu51vZZwCtIjFPNYaIQl2P
5z6/lFmE+GHZhlFJ7wTJGTLPtcRspfmDq7ZJEzy3K5URdlAK+JoWgsEcNOBUzNAR
ojktpVIBBODTBLRYB6zZMYT6exIP0gjkBcOJZAR308CVwkPmpzyBeXFt6VReD/9b
e3YgVTF4T6RpCmoL6hUxpRiq5HbipwVamc0GorJbtqK04QrZ1B0YuPIaskYF6fQt
8POum2bzbJ/6BXfcYisyLzSCzqZnDhK1lB/izoRGB0FYVXa8lRUXw9N/YzltQlbO
azmrKA+tjKkUOkByBMSLaiJdM4Zu3aiTVw+0wjCqkSEf6Ki3la0UB4Q14SbxxSMP
dkLjmln7pJntC/6UpQcD1BTJfceP/EIIpvVcHEo4ZwNpdwScWuEgGXBkBKkNYyrN
i1lc4iXWUZFU0hsEQAr3yoL3/y1Kjb9FUgBFgRMNQIQCzeZSXWo8RmtVoD4d3GJV
B479Tyu1D23L8OluNb27n2knbLlgYxUzXBJeldND0fZyNhyNczrWHMQFZlniAGrA
RiYpy+htCcqCAU7X44V/ARzuQO0vWNL4O9KFDqLEfIOj43e39zFDghDUg7qIvpJn
SIXCdDvffepJyPmZyJ0ZGzyqRLZmhdsSi6GQpguHdi5EbgUEtEo8oFpr1euSnwzB
PC76uSdu2ZfbeXNPmv2zc0tX2z3aiPMdoHME4b7SWWPJhjezHfvMJVPTRDIhgtcl
zTeTVskqUg3QgE1/W2snI7Mr/PdNJUzXwiHLFGHAcvoAPUcAqvlvty410yr8xXiD
B7NLpXzjwqsxP2l9oE3RnYFsYXAZcMXLnG4lOz6Bt4siCeW2Tjrc1c+i2YXzqI8C
jtSXXVQkejD6f5IxjL133RMzs2GZyn+TkEZp4qF9RQ4lvNSYARhPHhbrm1bG/gmf
oF+nAmfl36JOoiVFJVgv5GIjPCPOEse1ek9xK2qwytit9PRnOgrFy7lCYWIL0DnW
LZ+jVKAmST0m1bv6787k3zPiJgACkXCo8nfdZsa0V/dvazQj/EcKyHllOZT95O9V
Y369AKCWlmFOgrdTlRB/PaZItdGico5JlgPTKZUR+YgvvFhhNTWIO13MbM1wHyUH
ODZF5R3JDVi2epZOkHpGykViZObpK3/pLQx3ALH0zeH9JguMv/4GrHaVRNCHZEwj
EI9S/+v5dIiEitWk7Jcw9XkvX41KbFvxuKgjjgVPFEg7tSWJvJSVSlU2S69map5x
umQ/tGsou7w1jQjvlCXmCoEyqrsZ1tQl5EcmznbdZgHFsRcOmfOgoS0HLotqOpI0
xD6uvDxzwI0FaEmTmbUqQ7vzRYOHAFtSAM2WLBc5jOu/PEGcWToP42QZmvdBhz8g
EcVgvOAkaqLQ9hBMkRoWhYy27lqJ3nZpaH+Bl4VLzLHKVZ7YL6KqvYpdbpyjxDgR
0zwqD5ZhTKHw6Q0cxLB4CyB9BqruY389pVHh/N2rvYhxh3vC9lscWq8NoECD6+Fd
4m9bzxZLRtnybaf2ZLaSrj34acCIkB+mX9DF1zwpVmhEAFH0GgEaXORJ22EMCBWC
1VAVu2AWR3pdSlLy0gdAD6WKJUKGAVQZfbp8MyyppGXK729BS9FPk9BXvcJdvdpX
/7CiT6wc0EguHkdxiNxA87otQ4Geb76P7Jl+ffdjEb5ErKqtAa0DoPYdpK8kQ7lW
45lavKuqEyGIRP30RID9u9ay6WPjaSinLHWRqHRhtfa7inZMWXDciLKsR3iSFot+
km2bZFY289l//hsvuwYAwLzYKjgWQq9OUKaGJaXi9cpW95lHRju5uf4qwP9Bm3mP
yS0EhgT5CZIAwjruHPuIUmHqpQHfNmXZnLq3Oi7yx+asYb0HPloyxdCxrrGgr4u7
+FwCwdL2Obs2WZodupDJT8SAx+kv3sskwSZIs/t6Dj8DcX06avbpwJF7flQOpUVs
HbUo5j8YnCzFpoEK8Xwn66Dr1oRMIIvH5ueF6HrEYC6z9cAmEgGEPWkrM64BNC/A
W71KLveW0G4xgS8yRf7UkBOZlaJDU7onq99ePWzla4X8Thi0IYA4jGb7n7U4leCe
uK41r7wn6vrWVMxST2nGo+rU0/CKlVyRlAtRFohexvs8ZTBhxl6HkejodhfskvRu
6rXMh+QVrDy+MgmNbv4yAE9smul0vQQqCpcyhlPQRSscD7ssHJ+iXZ6lfnJOdtlH
2omNUOdwq10eJvevD4619vZvF1Oldb2T6jP3OayeiM4fkzCQUxtmBLgu4WnlnaRv
CdVrF84kUeK3CGnZNAx4n5HiKYO5BhyDGO6H4kiBEdq47T62S8TGmp44887pFjzd
3FWIfRcrRA4XEDtxq2ptN2vDxqdDU7SsaHSvd2kWp8pL7hDnmacXpOiMrIkAGiaq
J765m0GbyMFyEsEcPedIABZq2O+veMDdGGz/P4BQEgS/zRjvuVQwuEQtVNQkQ4Xm
EkUUfOD8l+p819CnRG0zwPUV1+KSJWJGiz+aTxWXMVAqJpl0UkTIftk0hjOgpvPV
eE9oedo4mhHbzoJUddKk4y3ZpuPb1FshTkgH7VVh/oeC7njVG1aTmMpEaZPMN6iJ
IG5iOwOcPh6YpY0GAZ86e9QDK8YSMtcshCbKaxfs91yCjZ518IUdPy+RqwEfL6zl
DoVln09aQQPfpHoYBQypAHJZ+ciCqrg4Bo6sBvAdO+Kqw1qhiafcMCaT8oNikQwx
8ykGA6spfgWu+/B5o14XyLQE5+nTJM6+aEQfWrhN+5C+1w4Ti3CDGyi4gQmrIy8d
nxwRAEeU2n+uIkkEHZrE+feOpcsF6GVbiEnMtM0Qs81QhH7LXSSOk0J8/ZyGWNZD
PHBg3+JkWZqAem2kBSkMacBoiW1Y5ytbjXE1mRibx/eMFI912MN9eedeFMDGn9DP
H0rrauCxHYzBQlD/Vi+PUAbt4Sl2btly3AnT/Vilg7kHg5rM3ta+KJy9FZxqYYrV
65cBg20+AfDYaoaAvKJdFY3+sICiL2gJJm9p0/p5ePJc09kDVulUJ79pBDlA5kxl
BZzXOcGSXxcT1XAY41C+SexnWbZ/HqW/whVN4jt8xWR7zi8PXriui78dRBhKhKVu
PRjcjnUJC3sI2eR/HP6GfDuWbOdho1v3pq2JdCkFEfAkpffg0IbmlE/JuL6dchMR
kl7st2p1WzddEzWtaAGfyZfS8n2NGnyjEiUzZB1+XRmJct0ZeZrTYxK9W+hIAD5F
YPx+C4j9royIIv9j5I+EQP5J0mzbql+5oiEpk8sCaBkB+KJbXSCygp+rd0VM2FdI
1wrK9hoTgNv8HrKwyMSG7Rb6Z8qmLwg/OXg3803QDciYzXR4eMC00XEiH9ioAVTI
iOO5H9u2UTB79EsvicS/zjQWv+RGTZGB1LGZlndBePpZ7m7gBlE5zcNOMEOoXFAe
7+9xIqP3d2cNxnCvRzXG4nE40PnFluROxX+qGuE1P+19H6wE1Ady1q5MXehUQkWL
2GMEtzLng+5njlwyNvKbFHO1oEKXitzddI3ufQ0pLORt/hzEHgBFdjKcWSyNTzue
KGMuWAUKMfHNcTxvXwDWA7s8X8SUKKJYQIInRqFv0WjoCoMASlSjqNJERtjLKoOp
WNrnH5EhOVCdt1fIQ8DgBJAar/p6Ldq3MX8wl5AXYIeQ1SVr8s8lqLv+RZUC75rb
/Li6jwQ4/cnMg3eqioTgxOr0r9qTDPptGWWbfvxgG63HcYp0PoQ8AOrWEOCfXker
GPhq23v/LmsWKjeBGdA9royMqa71S/pNsulxrtbXo3pWcKnrgpqEz36/4jhJBvl6
R7/byd9dhLar/ZHokbiIaB4W8x8Sg2vq80gUeirZW2h7aqVRVowN1XRNun4RwQRk
TxAiJX+jCFDs74/Plb/2CyjCeGY3VHCbVCmSOcyM2hqBc/TxfJZxopNjxlu0PyvS
z3XvPxxqEvcwUU6+z5HIjehSS3y/lLpMJ0WoV0BDP7VYuTsXUyG0tN5kNzBmdu8G
o/UGANtAYCvWsYhZ0tMKTbHcLLiuHjgjdqUjakfS1NHscMaCfliF4PBUVb/RolZ4
9RaKsh8DHz493OOOXmt2rvuz8Jj8DbXFKj0mBFJcDN/fDY0rJHFjYOK7U5xCT8cp
Yj1DEX00US8Ris7XLYqGEKqreBn7PjHg75PNlizdpU8An7jkHB4ymHoqnxFdZTRx
VjmN26s4sqyXJI9+x3oIzNGX8GyaYlNSnS60v85eZoMa2O6vsMgFTlpOlLPeOdYf
GvS5Xgd8bBvwgNpufTaKZeu5zsJf6dI8tRbdMsIEEEEj5Za1IHsC+91JeKwD00ay
hj5QblpCApkmqmkmBqRCuHdF3zsgZ19JSexmKtYqulL/c7bniD6UgiaUij4yLxK4
TOHjH6bR3LDXMr7FywNDCgn1vMFA0h9pyCfQs0dax6x3NfHBM24V9gjbdva2K9wB
aaFzs47ML+beFa4ESbSliR21bJmMCmjZED/uopqMOsam/J29oPlGdWqfIrsyOi7s
fBiTK9Pd4axNcwpkWsWe+/fBmyr3146/Hoof8uuRrL1Q5Q/eONP3s41Es1mKP/go
b6P5HJMMN44F1Dj3NFZpBm+YZhMBie7J6/rOidY++z8DoeQwLbl/WvRyd6TBElTR
4pXcSfTiyUmDiQz2nhB8j4Lu5EfY7Pv53K0ZZtGNjFDzu2efhBr3qnmpu9VBBDHa
aFpaHJj5QFvaNATxTKpGwgU8kkDiOQoEjsQehEK4nCnIh2bdFmitrqVSPCDN5owO
UoFWJnhNMRDYrMgBrMIm964LG6SDN50Z2leTwb88IVDIpHU6UqMwlSRV0OH0No4q
ANU/noU0QzsxuOcPaA2Hfh6JQBWnCy5g9HfnM4M/kgyzRVGw53vpHpr8Z0PoXGKP
q2JDNmS1jOS1xB5DHJd+GyzinMQMI2Rwh1TfWFvbiOAwymKq0fmOnff60x92x4vv
KY5a+p2SDRg/XuVE132Yeo013ILpdCuMFHdoqK7Bt4pl/3PZp/mEyOkQjlH9gmhf
KmW5vvZMFdk34GhjZ3M9nfk/n2zN730Q8Qs0hGCpZ/F5oVrr4PmIhrJbxftLRlsF
EDnrHL0A1fgCbFzg0V80M8ZzRZogFi+zT5DkIeZ0QaTPaFhUhsr0JqrRQhHLnw1e
nEkJ+RmF1kthGyI04O3Ix+SSJrqRITkHLXtDGEmeAVKzlAP18ywBQ6t9EKcBEIZw
96L7alDhagnPg4QR4Bb5RebGf4ctGuxkIakpBmDOSGcYl/tnW72mBdi8dZyW1DjP
kh+WSg0fnJQszsqZktsnINb8LrW1e9owUmR+j3YLUGONtkseAg1woM16teS9hsN0
iOqZijV4DtoMDLxegkPLQkdV1Gmu7qq4FgxVHjBB2P8pfK5ZViqK30VHw3SxV9qI
W2QvmDjr8E6MkUH0iSFjwpOOI6NI+at80GJ8vnZEdmeGvGyGuFe6a6BAV6kyx9Vn
cwPFkfGEu5m0L3WRPzwdWRX8Xz4rqb9/QzhDffn67tyFgPwQHJX1BmVj55Vv05vS
+Jc7lyIlgipk3JKGzkbyVcRvauaywRjXOIVdONV1JEMVpvz5gWlg7IZ2Mv61NtzO
7L4BhLb2K4rirtKifDtLSl1b6wrORq+4k/KHl3NpR6c7HrIEgUaPG1ZDemaO8x0y
BIt2MwNcHSrFkfEtdtENYqJ3Llme/3l1MCHZDIMOaD/uHsVur3xL6cXTcizALPPT
GaKMyM+C6lWrOQ2lwgBkD0AdoH690NQHuWNMV0yU76els/l314Jh/6EuORy4OVfH
uMcB8eOQxpbCPS6x4yy+2kkDLTrjf4LrPQsRBWq+wuZn/MA2dPnNIXjyhM34UFUu
5Gvc0lfU+2e36mNnKlKW+56TUH66scS7f/XvqXEVfUWEOOKmiUEBX/GjMV++pQfT
z4Gvf7kzo4zMraxH0+SpXooT1dKCKNGq2+jO+JPhmJU80Ei2DGNQ3LG6kjBtsf2T
jKYscrkcjywUkhl0AYiNMJN01SDQxd3Wf2SbEt+C/+P8SWjKHPJEE1cFVDVn5oNK
L2Fl1CCqcEjlQKw0T/NHkNJ2P4HuDyEi3MS4uPgxiq99iFoHeFVxf3FmcdjUISxx
P+zWNxDra6pbsqi8nEr172I+Muu9itQPMtWBA94hS6zvVcxvCl9Cj7tdDatPeMOr
GSmLVcdidXUKEOJ5YrRoC+7mlgWEQPvG4DvsK+y/8UgPbEvsDDx1Ubp/Dr20x1Mx
yBahm5xTy2Azfh3zJuMOslcyzbKuM7XB8Ett+2rSobyRr7amQ1wNehzRC2k7L06p
4g8Qaxf/itvvEpyRbZmNqXoKhJqaTmgn7vXLy5Qek1L/mvE2blcKoOV3Q9ItcA70
E4rBamdz8AUjHKhZXWIKVwG/Xd3SIFQxYQP3//olDkoIPAAyhC5mzq+6Kzvsw0e3
9VlU4IB3u/BaZtyRncoeaAcFpk5x3H+QDN59dpL104m2qg09GUBGByDl2Y+WkVZU
S+UM1GQBAUgQM8X4ttBrDVQwY7w5ixR/xvxiW2HYlWS3wXYahwwHW/bDERa+m6FF
VeoB2OarQDMSaNB8E7LdBr4HdgLo/u5MAtJ39JrO7dI6a86ANDiRnKo+YOFkDD3K
L/wm/atTrKhNgJvRGsumAl3sHTYS/skFKpsD6jVHOSos9u4r3VvTqiqNLLSHylRD
ieuXIvmLHDlvXw8bfl+O+sRIPhNAH54EVH8g/4YrTxnmYLHZdFmPEkbafVfMUWgO
6GcWk0TtCn4HeMO+/BHsuasL9YTP2nt9xoQd7X2aAzR59Kxa9gF8lYGICwaWpQA/
9WtINy+PmAXY8J1n3qeB9Eckmk5i7P7/832pmiuvuK7sHlZ5QJzsy4Z7Tmc3lWCx
nre4FvK9IvQtp57TJHh85VTWYp1ozdo3S6CohhViR6w3Lh5zdnpBHN1ziLCIdgZL
ykOZxKf7moFnhbHV5jB0ZetMjehVN6rhekB3BRzGMJt3hdONAU0vmtk3hkexyUBH
1EoQUK3wpHLHaq2TrnnDno9ACXSXfF/tzm8L4y9yfh0aFwZrr4GVa5BwtiWfsbM+
kIK3Y5ou0U4V2vvJoAQt/I/TQ90lhCZCBJNhb3baqc3nYE2nUWfJnA0UwNDMnENb
iXvLpPdaHNKzZWmolPLX+/eb3UgOFrFGZdRgA+qpVL9Cheg56g/603p70EFHluhB
VPq96/XSzYRuk3eyoue3yEebZS90AapUcS8CMe8J866/I1p0K2J5FnFZlfQHFpfz
nWHLpFihE/PzKKaE556u8BxHxTdQS3wno4rvg+k6BzpFFVYaRpgIerX9WEnlbC/p
XWI1oBemKt+tM8p0llVsArbIIKFvQIKIvzHYEyYcq21ytx6MbMaSXbuWtZkB4qsB
EFhlF0Pte9yTDrdoLH/tk+S/QvWBCwi0rkvzaDYeyi+6TP18fBn2KEZHFbHA9/SM
31MKnQ6RiEDbqyTHdv35FYAqaLJ2YaNvqdnPufZcRCe/tzhQ3EAW0s5PU1Pylo3Z
y+EzT8T1Ma5Rzaq9ZBaMIJGkLnplmKy34W0u2/PtdR2HsCrey1+xn7SECwikGjD0
d8ib/8DYwovehVlopeOtERBjH8MjggFYav8Czqyv5709YXfjvR2azoGtNuwOhFdE
ZiC1jY6fA5QiBDZZCnNaTZStykJ/ftbfHG7Ns8zSI/tRnWe3stIxyY9HMBTSiPQc
YWNo3Hk6rH5E2lTAwluA7RsLMXtrY6BbOgfLHGWGInVwz29BCiqaJdHFq2zFFRrg
ZDZsJLEybVeQOMbWVRNUbW9hkueG6ulB7V0LyCKtjzTai5ZBauHm3nwrH/T6H9X8
SvwYPMC7K5gSpRD2/4goHTp4b9jg8IMTdzTQyU0j/NRyYV2jPB22ZyXMbXl4Kaf0
JA/tqC3a9/tDScnuqAhxaQ3+7CMgWVoagFo5F4Wu12YNlqvudKKA0G4/Js8djpwC
REwEwFd7Xm9hWWA6NoF15+GRG8/2SNh9Su1I0jIbD/Kyb4FLvUC7M0ItAhLj7n+F
/RUG9ZjoPYkrG4ePIG1EVVjgN6/7wPiJ1sWUA3UmulvRPw4hrWEBwtd5rqYYBVBz
tbzAUXRAnt1CJyj8KWaaTbl7J+buBeDznnEkxiBM0Y+obFKdRFI1xZxFCbuoCOtG
zbKPqX31u64mG4DiEK0h7LvjYI8lPEs4QDD3HSZDegclX/KwpK/bXWg0BHT5PIY3
9T+IVDpe1CvTd2QaX2vw2rUmZDxCDyNuxCmt2VZr1g4TVCxLqkbh4VoIZ7TWW3fF
lePdppbWv2V5rj/kPBnk2g2D+B0DUxnTZWTuj78yKDt4y5emLN4a0u824bypuSXl
JKbsIc9RXUJe7DsGCO46vus0QlVzI7pKkmiGev0pMR38qpPmvxYyd8e7fhlYYy7h
mOQpHIgUDHV8AXIrb5IZCHziarHmIm2jzU2R44sIPkzseUBvZHig+7zW1npoNWHT
VBqsqzRUZFFnKXoUe7qRL7cxZYpS2jWxV3K6p44BddiYTsPjzAJHt3kKtcHVqIDt
0tpPi7BhzTK2TTw4eM2uXXRluiu7E/AgeAJdpmoqniJ+hN6e+I5O+7SLm1CP904Q
F8dxml37eZgVsagmGk1UcaAcsCRAtogPO2mrifDARuHH7GHBuGHdj5CSP/1c0FUC
NiH9IbrVrC+0okPmnOPecjq1pc/Efmuai9bjTlyBD1q0roTj5JyOABgCosQG146X
e4oYpq9h7XLPt+4ckb70/xoIK+N6Xh6SQvA0BSvdzZztipqDCKQfaPCWVvlDNYFx
dG3+ORCWu3df8vWbdq9oQwPQ/7OLqHOTxlJ6zQYOvsr5LORXMdYzTEFvvviRo4KN
+mV6m+rSC3btca4zwJPeb7ICcZQrbPKIij2NrcnddtzFDU1USEudq/NnjV8l3S4M
KoQvMAk/iLAngBoZ+jjKre6vYawh0LUErzfMEu0mqHTDYnt5JP4L2FRtncVruX4a
8N4GmgR5aMcHrJbOT9afyI8SMaS6dmQQv/9euTgA1oJbhO2E0u/h2ftFuHDFuKfR
k1VwYX+IxaJhKu0EQsI6ZvJYatayroIcV15QUFCbnmXSaEareHH09r2f+4gbPg2l
ApgFQbiPffNRR2iJZgXuOzF9QiYBJm6PmB3+fyiQno51maNaKHiENxrWQwl/pr0W
4W3lpcQI1BH5mcmIBKlRn9sdL/T3fcivC7SHOKIyeMMtf5bpDLoeO9x/xG3LSFkM
xVvwYlGyFl2IUwUrc7a3bx/h32kJFben1mpkCLYoKA8Jutjbau6Jg8eXKZT/ngXt
IDhrZdLOhwxQArL+OPQb8DdUM0K+0nBy4f2TiB9tjZ1I4WaWBY0Fy5xs0XOt1hXJ
m2L7jZpVZYZ1vP7zvcxEiilIdXDjxpZFf71YrnGnGr7ZcLCwxZYQIFdRXsHXgdBN
KH9JueokQMEetcK2eiPO2y9jk9lVIZPd/xdJio0E5f9vnu/dK7/tUJ7flun1lzNs
2Dp7TaK23RiW2hoCRqjdMqHI7Y2qulOlTC/6H6BRgtHuQh4qIg0GAAS4z6appxrj
dupAFkq1OQe+XXn3a5GaE1ZDdv2yRtZqfOh6EWuZtYOQgfxJ41+GP2WiibQfx87z
F7iXJsOQAU9aUdnq09GPDyMfKL2VEzaQ8NcElQtOpdQvhVzomJxdjmKdjQJKjvfr
WT+pAB9Deijbbo4eDajrf+FJpz/yAU7cElYzMm+BgGUQ/EXRJBt5g4lxpV3gYzFh
Q/h2nEwIPBGtrKLjXXNItTv5g1qqNZH44TFCkyF9vXM8kK7xLcayZKGRsY6HQNic
WJCRjnFvNgVwPlWnCILkrDOaTH4FIVJoxLcAIg4ItrmqNjTkVH6TvxDboUtmrgM/
o8EkO4R1vA//30o8ysW03E7wXNfWDaLy4HqA0HXv32jAt4ZxDBh3GzhhXEOrc+E8
405VEeKPwvztEIq4muLpABikCx8SrPNVL6bW+1djZmGyAuUup1vocYRAyKkQRgZk
90TMJa/kPowJ998rEcJK3tMHDXz1L9x1TKTnZ5iXZpr9SEc7r1PTUvJGkvrSLdsv
d3NuaJ/rW6M27wkL/KJ2oE8jPaUfgfDE0YU7AcnfmA9jvXJPgJsTF7pfpdqu1wm7
Jh6MSKWRGVfdWJ/pIuRWQSBXUnm7Ywoy3CYEAC1XRX8S+ws15fnASuM74u25DM9K
fQq67b/gLbIyeKVUwIlrmrJDRE4w8kGUcGh7fq/UZz61dP/w6ApHmU4QEAXaFj2c
AprmerfijrwsK48pQYL2x9G9Z94WUFvZ4iV3XCFpHYW4mJkx2uzsekb7WfgDflqw
zVtFclSNazh3rVSBLYy1LrfCyZld3MDGaNvYs7JzJTCkIx878wIKw16oEDpYZmUS
C2Gke3c6T6H0j/ZptRds31GO3XW15SIDOFbs/cv1wQYS1BGWKrbjau5gA77YXrFg
UL987LB6U8oykcRb0EjvkpyCl3DW40qIB8f+gbDnMCwfZd268bB6dtw+qZHlydHR
WFJfhm9TPYAkWIELFlauJ2pVdq54ooOGRTEeTHA1yfjM2z0UsOfefbi/6Y+ySjiE
4bRuE5SIKmagsw/QNqzBJ6pgUf+BjyAMwQDsefzQS2DYu19S7rBWkpasu+4Lh7pi
pk9z9+fvlaT9A5WIs1bszTYJPWdfA5j5YOUElyoGwc0/sk88grMV1a/sZELKScWu
a/OVtZ99Ub2Fmr6LRxc3bPp+yQEtd2uN50/w65faaQUE4FkhHq5dBQccu4gfrePC
7nLNrVzD933zMmqZEsy4BHTYOTyJ3+vjkVQdDFoxTw46pgw01SOwxH2Q4ANqKtpT
jcYQ6IK4qdKsn7deygpKDj7bG+N4dBpXLjaXJOpklsaL+N9MtjL9VddrbR6KzlJ+
W+50kt7ySVcfSfxkaItBo224qhCamNoK7oAz7Wh+s8LyJftY+AFxODoiPj+atvlt
gACRXWOMXF+WPDQKR9CGB4YuThYKqfDsGCu8x56p6RKowV02XAmT/loffOu74lwH
dR93aJ3U6uWey8sCToTLFlBkunh48I5q+7t6bvkyoEk3zDpQVp0MHs4GiZc3mxnO
It8Cp6iQJeLq4yAn7lDgJxbnJWomhugtmP+Y80bsG7+vQ+KhtxGsi22O64H78Jpt
7/q293XUesSDX4tvmLXJVtEz6Bqj7TNEQ4H1J+4x8BKaNmHA8qWP1/8Xp1zWTlcX
dXK2LhCODtw9ozaGYDf5Tg54QJxNB2iJ+zFiv+5YctgUYOkBX+lprP46GzoSsh+e
TmUQvrJgNKwJujrGcDTUaoh5V6yCy3w1hSnX4sUn/WugJq7EzETn71DQ1HrtOnxx
KhWF9E5yjWf37SX6xuu1SX7IyVfJKYz4dpGqt6XsPZ0AtY1IiXM0mXGivkaRly19
ogUNcCaipIesedjZ1003lEbZuN5w8MgUCqF38uXJ4F7aeznnNjmBZnkve6PVgpTA
RqGP0h+F1cRku01mVtS3NOu7d8J3ezyS88Gpxc5yR17YDIxhHIb5j/83crtSfSlE
g2GbX8VEaHgwTwWO3Xk8eDVAJ0u/nWdrip07LZeBti8CeO9cegb2BGXR6kirvIe6
mlqXZHolRSZoTbSqrW7kM3mvxA1USlxi8g4QH8ZnuImN45vRrDVgmro9ztB4QdBY
Z2u0moLrCF5loI/82bv0aBj1AEMhpKtMl3SyQujpN0lk9SrJgoyd8DEJ8JL6k+dS
ZTmYHsBmKdbf53l+5EWjkKVoSfauDDy4016V6wMO1jNgERoxnZrFvxhPA5eC1aXF
29TC2eFuMXp0Oi2jE0i8xdr+o9cK/Jz1307YX97s0RFmVI/C8ixaZvYh3RJtFAo1
v8aJK6Njxgpmk7ByNskXrjtMpqbYNfzhcGamRqbfKc9opyxu4s2sbUfeeIQ2VmKK
1/GfE+2A7lWguHricVXaY4nld9J1hTzKeFFgi5vrmuFBtYo5jTT2QITT8zUlPjvm
6EKei6iAeQ1j5V24rAU5IC3CNZ8DqSZDMsPdnEKUnWMB4u9svVlerGVMeVNBzcTU
2HIIkPebigsCB8NLPR99UfHGlAeFzwDNzyRHt3j8FrOi8dGWng3aIkvrMJuDgYbm
70zON9evvBLycpnojJ4UJP88KmDQTks12XHRbkUUj2skAkO8wMaxuhlJZTQvcfAI
jK0fBSZq5EYHGZxYHMlrllfblZRJ/9fXao2QE/6ZxlG4kyuxV2HThdUPjLrVDSj5
Gf6ljtt5ysS/lR9orVd6X668E6wr3kKV0EQt9b6igvDObzHkY3xfE65SHPT3ZFN0
z9xwKHxJ0ixXQHVZQ48hZkNNHECL/QwzDo1MTfJidC8GfoH6OeN4P3MCGPonGKi5
5tMy+XIzJkXfgbXL8I+VKu9qQ/Ad7MP0NRxLQcowN24zmWPKQye01xPNmQtFMhyA
v0UN6OIwUkGGEhNTBvWz660U6MyPTJMtOZvq/YVXCuUhEZXLY9PBo2z5OxsCPoNo
Zcxw1OMhF1rYbeEIVeL46fn7zmItXfvd1/nqt9ijFDgMBwmyfefYsOrf2UhiX86U
eLY/1ZB3erAJx2tQgcCmIMZi/kcit18r9ZY9dOxfbPG+q7BcRWSm5epLXclZfcQY
CTpBrgDo3ngXw/mhuyU5VxoMNVqMHAdtiFgDxHylhDKm0815XKrQkwz6D1cgeow4
4mZUyaVpoffAyTyv0fBAt73RoA1eL8YJNC7DwO6XNW8Dai33mgjMppn1hNGu9EJV
VuiT/3HIfzATB1kEk+nNHTX0tCA78KJ2bcwrAWnjfANXxNcDYZstrLTI+GNoZCcA
bQdiBlWtyWCkKSIPDZ1dWZdCFShxkIOZgDONZhqjK0ruXDtCwb22JeUa2LZ3HKVQ
vDLOFnizsC8A0/un8pymt4xTUw+RW72RMFGSk4XjyTQ5ZnhUQfN9U3zOBDKRD2wC
FYeUdCYpjozAuRydIpHx/iyDYpcuSP+D7oKjCbMRwOiQZx21RgiZyTsD9e3F8wrH
2ubfBvQNG235CZxmeUncmth+JdRfyWyMNolbD3rQhujPHbM+W4Bzux2rHLj/mUhK
M7hx/KNHGJH51p5e2T3ryW5Ntl2oJNEasjeJgCbJLZEcNd+D6qcA/GL658ICtgON
m220LEoF0wVe7rcWAEYPCsRQVNPQgjAt3nd8UbnEB9y/7HctYo9LwMpn3jI6EKuw
tP7IrZJqmN3doA5ANt9b31M/3UZ413KU5w2dzjPfn2lyTpdRt8Cc5hIJPQegIuTw
TdE6xpCClP66aCOl6Owyx7wh8lfEB4MuMb9043pQGXY/G3M90qi2T7IYm9/VfkD7
ffpgtbuFu8cHsDADSdQaQw6iM8w/jAZU33dLw5kW47f84I7YqinKktRn3OLbKkEX
PTxwHOs7pF2NNyJr4nRohZow50j75zGgMmtfsySUFwmA+7P9HevwN1WnVLpt1kfu
rBF+EaAxpWzjb4oKyXjKpONarBRevyiTu6AR5YMDUahOZEfxQayxT3afSFJk/C50
UfhsPNZz9VsR86q5SYu4wNNqCR+G7yQGVj8XW9NkvD+RpvgE48ejKegvHUPmVA2U
4WWJZctnVquY5bQUsFsPheSvjBDRmWcKeGWhllRNqQLu7+xbUXzLw4x8X1LSzPsS
W9cbVYd5Nvos43rRSHQ4PrVLZHQGkYTs7ORBhaVlZpte1ejqFNFTStapGXPTOZD9
3s9rKtChg7phVTPJRaWtXSlq6tid3dtsohtooJ74yk8ZzOb/2ElE6zJ6DoOC75aP
c9ttYnHbEOf65g4SXPx+V46DOTNrq6LJmlKcyZyxp4DXmIspbcneSQt3C3elpwMO
DYVQ6WSDrbhMp5QpSBp54OUd8osNByHkJAba2EGApkYx2+7wThYprm5kLlxXCopb
WEINMq0y6i90PKgi67cH/x/0HQpABwXqMGMsIK7mfg6R+Spgj9aP5ZpXGhZSmTYl
JUjAPHIWbLTJ0XhEZ/SSPqhSIESxppVjPCCnjVVJJFm955ZG5NKDy6mu4nEl6xf7
6Nlt4CFjU2WiU2cC4Zv7Jt2I0RbBMmFCMbjB/uYAPaBzSqN71Y+rKs2Eg1vrIJ9j
wmj869S2z9L+XJA3yPYPSf6/j92XxQO9Tgcez8vnowMGKyYGZBxgzTMZABLLs3jp
8Ca4axielo0V+SFa7WwYcKG1P4ZuHDRP8LXycfM7iRI4pCXXiBnZ7h/xvcXCgCcu
FMrPKubg6Ff+10vxSGjxOUy9C2c2Zg4vOTxyyIBu1e6DSm196NUv1jFn7MIYulG0
L0JSwEJhyHB+m5fWLGNHMC7PVw5cQ6b/UP5koHX+Q7V7wdz/wqv1uo7kzEz8l0tO
9G4fdfXGIPQ6m6IQOkIpyrcW8jMbp4m3XugRhSWxzwxnWIoJIJA9ysEtRpvlOeoi
2N9VLb4ROAXFoMmKmIfwRFIjRQmdkcXsJX6vbttp3xsNPFCotpKRgIN1RKx30+zg
A43yNPqWiQ2jkxwuDGva333yGn9ejdpSLpel3z5elPt2zUKTrPwblNbSl/BfeO6z
CsY+bRyut4Cg0scDvHVn1yb+SVQxjnPrD4+uL1ZopJ5Iv6D0jN1FBs7qs+35VerY
HWFYcJouIsTFq2956Sa/d7OW94S6awRQAeMBNHx8g70vX47podA2wZJhChs4fYXS
Ebgh87nZ+W7dUh7rYwa3EBkmcfVXcUFx40uzaM1Q4ndDWs5XP+QgZirFkQmIcXZ3
6B+mfBYzr61NIKGZiehhlwQ656kXyy6mERYSJm78Bq/fEQPpXmToLkGN0aiUIWPt
CjcPgaUVX1Ud7bdBnQNxss0QMAk0gdsFcvD2FKodgq6NMRM1fI0vQM33Me3gMQBz
ACFF38mdK+MwiQ4zCBnk3HDehN1Gyue/IsyC/JoUvg9vLMPmmZtLKnuJ2CdLTrzs
Ns7aiwRLGaZMhJG4bfHnLgD3FdPdBwO3HTwXLvrQX65JJejUeQOZ49OUONSoFold
TQGllVUbcwFKbv1D3Qri62ExhyRMbEI5nBO+BuImS5PV3MQ6QZ+AnDpwNr051Z0Q
ZMUjTDccQe//xPzcDh3u8WpP/9oHDf21Rc4mpOIZ3XrZBs0VSVU51zKEayGQ15zz
tBbFKNyv5ehuq8TFuYZoVa2Fyn/kpPKv6c1iAskt50jJKfdSd1bXUJTXNoggw7ku
9wG/Ekb00SgZ4mfLyCdIqSKtAnSTS1OE61zsRCUo5dsBvUX7TBjKb95BDiWvC0EF
yT8Gpa2gX+EITP/Gnl3xYKFnXNAKPzTopdLiljto5b4SXya0kSHYsYoadeoU7wF5
QboXW9vvr9fTRBRkgPWnW6Z/TYIOKzs69hSr+2zu+znreBQDy+68i99O73p+vPcH
mjHyjqJE2CSbQgRlzwEDJP0WQm12rGQeGYDfqQeyJw7WxBMQMf7HPdC5LiA0dLqR
DxetekKpCOBAsz0+KdZ0ZXDj4pprq/myjOY05B1Cv91MYQgvmQcjwV7xj2EykjDY
fGFVVDSe9RtlkyMU06UtxrUlIVFRhjY3+j6ivHzfeAG8ch5WUQ97sXot8gX/8QMB
2OHWUeseaeNba2LxXO6jyRuqM6++Ub2BrTDAucjUw9xioa7j+7kW/4dmSBWoVi0p
NaU3npulmMM+u5r6hR3eMrmf1hpBiLM6LZYGGDQ0O5JurcjDFyeWrL5xQRRuDbJK
v/CXej6T7eTstfvbjQv8MVqpBb+YvRbgyt6NjqAtOKoh6A089nxrW3qbYPdW2+AG
EROSEA9ZM4pfqYFDNSI4msf1XJw6wPl4+UxGmCTLfNcPOHiCwTkNj5M+euUA9qVN
kltTMgbAlGi9sGsiKjSZLZC3k1uVDuq4z4Q0f4KmGJcf+X/G9b6zy22XAErN8r5Q
TICUdgcgjE0p/yeByJeaoGeAi2z9PV6pQy+UcR1eC0aV5B7oh4VKAPAd2T8+dTOG
P82c1EIOcGG5EBbks0be+26ShTFrgcaNDiMoT+AqCAB4fQLEO2MiYmBt/Wuy3Vz5
GuHGOGJIQt7AgM1JcqW9iuQILj789IdjP1hCRa5YB4yKwjbkaPn+odeokbJ59vWZ
bPRw6rD0MhG5J2/CYJQIwdHXt8QaTHfakS//BGCcoim2aK19CCkSsC7RZlJDg567
e3IZEWKrCk5jqDIVdCLFtX2bLl/++KowDW9rx7hALrjMu+6Dou3rnMMS62febWz4
mXIL96OLk849A6fg8+6sDgMaHkKJs6JpVnS2V+qnYOB6Pq/UrriMVmHzNBIX0OKg
wV6qkAJATl9wpUBo58lBWOcni5sFdtzV1+7xhJmZQhX37E5v/DGJXSDbtMigzMIY
MrImHOPBDIFCfkoJSpqgmJm/J4uKCZfR3If6Pfn3Rqp+greDo8v6glOoavLE4Z6h
kVPy3o9gjFFJGoXXt/+t6RDVyWa67+dz4VUfAQdNWPOG0aVveUSD+L8jj5QSWRY0
kCwj5LXRLv6aI19rVELrXlB1cn1AmVxCTZk6J+RyVWVpCvFbOAx2ul/VWqA4zlsw
vkn3Gnb+7Reh7KJq58vMdoL7Oo68eQM8wBiSDLZtj1Z9K6cRweHAM6+t+mmJ/Inf
CtyfnrnTXK75WxFnY7rvIzI1LQVrxko+1+FSPqgSuVCmhfaAsCxBn2gtCLfzp1WX
hFjtKjl06OOcW22hrXDobHFsYdXmjb+f5HhDLH1iHGS1CxgiZ/tBb+DKHNfFOT78
9lHJfcQ2gyL7GwLZK0VFNNIbLX8oqjb8LIjsaf8FJISCQwUHRPEELWi1G66lj61h
Sepma36XZCshWzQ5p/J+C6HkE0pc8T/K8yBpD74RylgvEZJN9TfD8HN34L1OOn8t
TxQ0tauxBD+9VFS/rkF57QWFswQq2b8qr7OIx6vI7TM9vhXgEpBjXZJN9cvQwF/f
ByoFgxbePC3hkf0ckJA2T4zqE71/M7YiXN2ZlwE8M8UEfIJxvHDW8mmkCha8nJlm
J5YxWAO2Je3VbNAoVeuIpybhafV8FnGnrA9ST5eVJRGqgnjaX5bVUtBcqlhMnbfl
C+GJBCaLANWAtKbhGpbTd11r4EEETsysxhS68lWcTfe4JRHmFV5gb69dceHIX9N2
+Mv7VNT6TISqAx46S7lmYY4pXFi+MJUnT8SrC//yKtVVz6coHMe5K8Yj27drhk1I
sCYvmsooc0Kpwx28RBHKwydX5CuVbcHVxgUFN2ynop1smkTUIZNHoraLvCv/XFD9
Jd2plV8gFeTl4wFDxfa5MKblET+pE9gFbAcCz+knSxcUbrIN7R1DFc+Umh7CVq7j
K0DdV9oFdJn0jmj2I9Mxz5bw38bAR8LHPyWTVOgyQzFj5B96d7JIjBlNxwCUkg6o
wEq21/gd69VUzxq6QaR40TkrdbIo4bR2y/lIvNkMjEpiNxSNJSnntr+V87IfI2hc
YsRlULz1Ej3WlnQ+Wbnj8WT6wxrM0gt5CpZF+PXG74KwqxVcJkTyTwv7R59QHpdX
YRlNzQVODvfpooAi+v+mgzeCVHc9Uqhn/XRl7v6ucWHjOmpzSMpFiBvLczSI17VH
eL4IfutOkQJuyFwJxwAYL8qHnuMzjtl/MY9SiHatu+0aboJoFpcQpL80/BBx8vzt
MsRZqXqvT5FFTVsRMIBBzwL7Yf4BykarCuZwKhoUfHVK/yNPBIClHAVLxcseiFWl
AysyC8u86zDCGAR0GMBhWHQToNGWPdqns43p801ij9+FSOC6RAe1ImYz6yK2PGSF
IXW9xmmuquOI26Untk2VNIOGrZSyQxHVKA6Z7AuYic5pz3mGtPS8MpPQA4SaZhDp
zZ0jj16IEX43svo27YLbDpeQ1raBiU6SAswRRqNonMPcxuUKwIwnqC6SiCTC+RKp
IMXmyIcAoVP088DJC4RJPRHidYqjJBWpjV0L79MAa4C4HMErRp20nZrBS1W7E7+l
M9lQ+7C6k58Km6sdc9eWPp2ycgGP6xXTMZFx3aA0i9XkSegGkBbYGeJboYQNAY5d
16K84JI4dzQMCBrr7YD5ch+J3vf1bnJpNQRTomwvLi9+anvfrXLLDFzwiZpKxWOw
41liLcTi7oDjeijU/MH+Se+ug5cSCK6wKJpJm+E7H8Fy+5SPnzRwTJMGWFVHCGoM
cgTr+oVnt4Fry9RJwxcIwNcyoPWaOb2aK6UpebMIzGeEH39WjThVhK74xbS7geyg
4e8H7Pwa6rCzDkgGDkMci1WeRwJaZi88+qTg5wFZAidgMcMVNO82CfdLf7DPXXhR
CREnGj8QY8MNTL6FK0pz5KRMDOgXjpMVF53tHcJQnKB8/qU2wOayqV04gP8pNaCm
LQnD+6c2HuuMmOFqTkxYgFy0xXlm1ewDYxMAQxeZzbqxUju8IsfTxzs11aDXDgcU
wiAbJeKNHymbqF03qbveH4uZDi9mnpsIry2Ve/itBex+k5mwKnn4NY46laY6eL75
YUgLzYVy/ohd89CS4boalQmvQfAyupSQtkJ6h2J50ZK9lkWTZWKRS/0cPAWjick9
okMz3kBd58kLBqTAHk+KbFLoE5kLxi+sV5h2/OyCDLQLj13ykMvxtbCLFa9vSDTn
nAPn1Sq/uwbBMPZUZ3iRQT0MaIpQ/5fwsUmZirwDBZUZJRum/IDqpTGZzot4V1gt
dDpPcwMJ3Mkk6FYtAn1EpwtK4QCJEao5/AU1X0a/MY58TcKRqxCgTkPSK5DIYLBJ
yhlNOPUQy9wwPAFMNqk/Amu/VK6uPYzlXTMTNf34GjWT9fbMTV6qTtuDYNyabpDV
6MZI7ckO0k8V74k7N9hBeX7sKQqAZzAwQUvwfOaP7+LVuOgWUbbARZTuXsMsdRCf
mfHJ1ijMkYCaNcrwknEgGgvJl7c8kXsktd4sQsTchp974qVEDgPAKd76FiqrQIdJ
EYTM7OtBTThs86pQTR0cBc0bd3bVg7463nP6gijg5dqC8dmwplALSDnNfoHgtnHF
/SoVd7yZf3/P0cQjo+HqkWZaU5QJknMWid2p3MTNPhh9rInxnpr66AU8Ah/X9DhG
0BzWi0T+iYb0t6yAJ7IGYswrf5Q94HCX43516H7RatsP0pVYQOzLHZWlEgDmIPsk
vUZCgUxY4po6Ob6F8d2WaUlE+riL+CMnc0fXplHZjc5FDrdYlBIlJaQJFkpVg5rn
jpBJ8id/mtKRHCGQAJhRJikrUwzR3A0EdXQUTl9d2Kzg5ri+mV37ScMVWDBQA0kN
2521KpHvMW2dsVwHCXvFKo0FZ2DjHAopbso+rRBa/UWVBPJ/C1XcrOo7ZCR4yI2Y
0QHC5zCuMufRi0yrUSsC+4egvRUrl4U/csDV9G8s2s57TPr8i+16tcHHRnLkQPfM
WbglObdXdklATIjVkN751Gb7ScrFMUSsb8QG5ke3yLHWtKAsuXn9kLbpHROPNySr
aFDgKJ/PiVLVZwyCiRI4hQQ+c8G9ivQvdFbD/ecxKUFZEjzwWS0OhShYdq4xaXSf
gEv7BEVPxblvr7cyfodiqEN6ih2ush6J5DuLZvCuJ5V7Y5SCCJxk8nNkEsWke8F0
alKnoAVeNAO2LWNUfAkZjuJJRTzwPYyEMy9bt05NHCZEWnS1F90WPjL5Ro3NY//m
n0cCDqVVwviWackMkOxP2j/of+xWHLjX+UatjRsnDmv+cV2W2fCygcBO+ymUT6qQ
1x11AvACTvVoWuIY9Hn894Q303Yz9eTmo3Ljb+gA0reCTv7GDUtQZ6p64nlRLHkO
OE1IELmzS/qtH7HjZYiuaC2fVQgXuMu+OTOdMbnYASgi+vhjQwOyoGe0oQzS4vNA
MNuYQRD1kI0Xqx40O67RQv5oj7fbHxDlJYAcvJxkomywqaHCYRNyulhwgk2Rg8N8
mpWH8DmZY952Udqc7ToZ76BM7JoCQy7FrD24brHYj7EPfwpjIEwPv85PMIWAJiBR
ymmNgR30+NXGz/Q5hGzy+lqJIebkGloqRRo8hG433SrBNRi40AhxYrmqmcindnQf
BZ5rYhc2SZisXkjrPqiVW93pZZqvg4xUCX03txJVTrK7KmuRlcFeOuK2KIAHRaVT
H3Tb67p+KH1hska+65Mo8jWD4/ocu94Exvi8/C0lzm9H1GYT9dE5iOMr4NL3tJAQ
eUZH8g3yjggc/Q7oJZesLso++EgAemu8YUI/4RQssCRGcsvvFxcbqAAKIJcAuvqi
7Bg9yLxKRkRVcH6ALAsGRUNZ7szCZYTN6h3hwati+PGnrSCebVTITrwdudG8+YAx
ZzT7HAmI1yrhnXarKnQ4BNGtQZM3xrt3iYscIMA5Wgb7BWDqd2zOwYqE711FbDtv
LJAbtbbflBl2ywiuf7vvYZSX/pIXAMRlxDLEzBwIJKwFBZHKKiNN6Rl5UqEb1vH0
3CDkcaowcc/6TzCbuX8yiWZhJLXEzjyw8yPS3HsSHLQIfYU8oCKcMxs2Ata8fzbq
zu05KqNfHP7gb0FlrQywHKj7sTBav0+HFKhPFPeh9WulEVQODkBklTKiaQW/rwEI
AjW4IJemRQhpHu2EcUNK0uSmLXFbuf/DPxPOFhYZUdjKdgq+NKXKgrKIWE1yheat
CkXQ6Wwb80FKXNiCoXNe401iNa0vLHh+ipAR0Z2CCekKx38fsX6W43aXIWy+GU+9
YKDwGrk1/TtodL27/MD79i2htTUHbI+tKC67tg/8ZsM34UQg3qfCT8IOpo7dUWfC
tqRyuhD6Q64SXglj1OPmZ+gzQOFaticuzZMlUK1DDQd1ZYuRJU/DCR+11uGjLnRy
oWrOyaSiv6lMULKeMDPO55ODIxOKw6hOATzomIyitDZXJZ23QFApJl5ptL1vXllL
qcUv8SG0Hh2bnC0ifzbvd6U9ENRBA/SDbnSdyrNBNSib5D/77z1tF0t6x5XFlPkW
FHlW4J2eD9xBSLIDnUftnbQQynUVeN9oqdd4yqzsCZ5f4uod0AU0jJ4x2Il/XFyW
J6yMen/JrolOh1TTGjcGif3S+JMUwPo+RacKtMyr+q6IIdy9GpqpjjjNUuo012yM
S4tY7NV/7F1oRmZ7n8vOvgyAzmGkSVBlB7RelG2eTQUzG+D7Hmb9XwMvM4GoKrql
/LSTlv0ecCZgYXWOgSVGv2PxS04zufjTA8Bc42aaf9PtZvuJuFNagSGYyLj1/w53
uZ4ezsO1f9jW8WNJR9Cfda2GvdtXIZdPJYe7k2fSvAV0IG/MM2KOys3JGB3BsF8I
+0XO3IsAwRpWuTNbAgGak5TyzTx5EQKqnEOr/Txe6l50G1DUaIYk0EYi7aLt4BJw
9/SCX1VWgEhnIEjYQo7RHYhg2T5+qHkr61fgk5/iBTBRdrDZXsAuCm6X8OvSu2Ef
mzd5XMnGClkjjH3Wvr0nMvgeNnenz/oKy9MUQdrBFS8LvqVQYglHCPbOyltzOdGc
vcIq4Fe4jli6klMeq/VC0BV2D+SVbGL3hLJY13kKKUjdrt+WsWKOB/MaqEW8N0fI
isN6PdN1+r7rHKW2CP1PkSoesG2pLjzG37kj4naiyyw9Z60lryJuJ0tOOie+T7EI
qbw2hTomTuyRZCs784sCJ+q897C7dbeXaDUK58weGNeNVHnTs3p/DThqaWXPHga+
o/yvTtAKoDDBUWVC+yxjM4slzNbnejr44BldsikFsm7GVehfW6Bq5rTNH7fhsP0s
z97pk7SpBcRfUA1Bzz408JlvTT9GyQP8yXwriw+A3Ql0rJ+D/LI1VIbo7yh8tvcO
jMgrGmzW6dDriNxthbwEcd7EAY51/7xoIQWxKHAOQfKwIP6T6Ls0wnALHkqnVnTb
Q7TxvKzQMHT53MK6NTHv3RLmzDfcyIFEvJeV5UcM3qvVfxuTa61/UwluCpHUBiRL
1vBbo+iMfF+jppMVSujEARLEr+OxYjdl6CxQymRAgy/ckzryA/KoHYGkTvWaeOoy
X4paCXClm79nhrf9XdNNEWDV0d/Tuz5C5Vi6i2AlRLsu32UdMy5BsraZihqSozrh
KC9BIuDU2SUrd0pGSByYtstjVFOoX8YYku19p9RhK0zKo4YJAW+E+Uswxi2YFv1o
7z6Lvd+kyulOojdhhQCmVvFcCNB0Tkp6dAEaa43lBCcFqjt4YFLRxAsAr51M3Tly
DgNRRZbmJvwdWvznWxa0Bs16hV8W83tloLoVP+wuYi1y4jzcNda/6wWeanf2EPAo
b6uW1j3+IJeSc0xNIW5aEM6AkW7Oa/8KtYbQZJsKhMW2HKv0Wl4glTp9hj1RG6Nj
9cKI82Z6B7kGuOcowoSu9GawKz0d4bTcw2OlR4ymABlQKhuiXQk9+V0NTFyHeg+0
jaHJq+qGWxNZbipreQUL0zxWU4hrLhms+WLn1Dwmu25+r2vbaaPET7It34eVEC0g
QgWoVUWBA6iJ5nsHEPabBa7+cSNtCY4YhqHlF2Q80cB7SEOS7FZ4lGlueBh0xINt
kYiaZ2rux8NBlbgkk+qpUqDN5CXRyFcGgV2mxUUCUAfC90JaT5m6xHJKOEKHZDcC
YxNXWg5aLRB9b2zxkkLXdGWMOMoNRGcdpkDYqxA5QPfXUrvtXUXg5SjBK6Nzw1wS
AouDvmf42Bbh4x90vjOtiwsxNHiav7uTsxlLaXXSNuyaonuPTwps0Ir7GjiiFNpC
r/aQ9TUi8vq87XK09/tIb/LIIj3EhEDwaEjVqKQNm/ibAEaT+PfN1YfmblxKgrW2
3xfspWlkObiqaounZp3lwY1SFX+qNVp6IFx1XC5eZ8yOwzekenJUDmE6esOtMBd/
uM4hXs5PnXLzQ5ubICxiQfJSpzNZp/ysGUQG3Dx+Hcb2L9pdOmLmLoUM32XurQCQ
xcxBLlyHupO2DNiTegwEc4Hq6beaVGJ7tFIKRQLRx9glh5yMPEUW0NOVL38MScg8
BmKn5bFJeikO/gFR54dJzaqeWX8jIm8zdbeKzZdUI0IkPZojJs2gd5rmPZ6iilfL
0H5MI69td4vfln/3PkoVHCJkJ7q/9+Kb4WLcJ2vOwtyEkZFmNXr3shSt4Ih+uQei
20VZH06e/7Ib6ov+r1ihm9BDM0HoEdStjFzGmO1AFyNJb1mflZV+cThi3Xj+GBmZ
OsIdf5S78gP3MESQEI4WQ2NF9xFQ8+2A84TR6h9GMcoys5Uz/AdPdSpvTXSG34fV
MvgugjuXGB6QuCpeyGg6CV36BC3idus2UMYQ9j5d58BHz48UU/zg8EEfSv0N1WW7
FZDrS8jWOPlOOVHeuWzokPwsaLvxALB7z7TE44pzcz2xONZITOd5k54RL8TLFKm5
+cF9q6kKHPl4mx0qU14LKgm7KsFWZyudPzbxB4AbnVuKawIyE19AbNQ0fk+uTGP6
5JeirQPHk8+MT78Y+KXlOs5vlGR8HhW3UXHMMnDduaAiL8neBmopcQp2PbLaMkcm
2FcsWJjP3zKwjvANcMkc6ovNtCIrkl6KhdOb2rCHJjGMzCSJsl77x+2qLYFzB70j
95Af7T20MGjc0NWnI0weiMWucmskoCppFGweDEZuzYmbKX3PRsoELHbsfhKmqlNO
M/Pxs5gSbjnAGydRuESm0KzCRM9sZcfZS3U6t6c4DSUwZRgBDChEsd/1aOu5R2OG
4y0Km4M6yM/0irRmOLU1UWT5rw/unfcn/Le6AzDhySPGjbQLujHmG8X2NnTR12nH
RomdDhazT+GORMYzXnwkIqBKvMJXXdD3VIM0LjW7lfWCh6pbRB3fxk5orhHthOB3
AjlC54ys2IScyK3ei3Anc+H/28nhH/sNtqbe2Bt+YumvfnNpU5p7zm8Trg38b6bq
XN6D6cJE5kIHHnLRsKrTYevymbpcim98/hbeiQHRutBDbWT3C77bu7UoZdtPSFaH
tzo+Kptup3huRQQnoW4poh7vu8bDw8nAlVRfnMfjFDpGZiKxfTfq4BlzXuLjGTSq
3oKjlffs4WQhxaA6MDum0jfLq8py3dwSI6GL/2DfUyF62IIT7uWgB8dqEV+GZWDA
ProLKKB2+B4XmdWR/xsEYLOZDBG6bUNUyk88szoPEu9VtTBbUXL9fXYioyVgvlys
0QfR+X+rbEtzuP8OBubU2ym+PQPK2JX3rA9SIWh3073A81NvDX1Nr/gyJn5q0yHv
e2icGgqcq+tvRx/yi5qqEn02pXTBbBAM367S+s4hGPogHK0OfHro6EUbxWYDv2Ui
XsLFZ/rxUjgEstY/+/3Lnven7uUetDn87aJ3itWFO2oO+7z5MDg00r2RMxuwFIPY
+7HqJ4+GQ8qA55MuY8jmKACHDUI1LINffRVxHwH2cMtf4BsxWr7SjWBozcwp0OMZ
qIBJZCT3OepnGJMUJSb6+WYCCmTZ1T1DOSXh5szTyNs85ffONFJLKhfQnkbjF994
eMKnsHaHUqKRt6eeK4H+Dtx76aN5Z6knBBvO/z2JGZ5XXLTl5Dd95IQhw6/7YP8H
ps1PQCLvdUDcfiDfde7oT5eYIMi+S1/9DNvy+p+g3YCMFlVQGqG01f/+/JYHdjfy
sO4E7oKcRWpWbFww0kVwqKNAy3bsjjRjyyD2cj9dy1adtZlIcYXui4/hbOLKo2PK
osLJoJbXpJ3l7sy5APRBSDQYpWn+HLhNtrvwqaiIfF1ZlYRftok5nFFtPRrxLXHu
/vERbUpsk6npsW8wSXIgWyA0oT77GdTajmaFZbonNUkFI2QCHJ0b3dp2/H2vs3cf
toI9rGHtD47FSV53LGtREaRWFYwGUfceBkucgbnJWbir/pEh+hY6eKlsT1Xk6yDI
ZCgc4/ErGlFu4p/smzOjtIAY/rhn/VsqKUAffYFzes1E48vRpKBNBSxBguKHjS+s
mmMbGVEJ7/IuT4yRS+UrrUmFB3X4JwHzeT8iHlCD48J1wPvysOQ0r1crfd+hncgY
RsNfJlpWRemD3AaNEKfmWD4msFgUf4s1oXzqM6TFDqF64AxtK0IThe1JZ3JuhYOl
Qd/9Co7LiMAg+hMvasGZs2OecJs9/Ky2D+Vosl/4FBNnfz552D0y7JksKvtRHghR
WEbX92Q5kwt9ozpGeQpcQADfEWev0joNhncJWeaLSNa/oh0dGKb+Q0GbOSRUbNku
I2A8wAt70c6hV2Mq719s7ankzX+j9pzlOB4WMAl/mpBaCG489SC2UVTR7LVJr/MM
6dLFal5wSr4xLAxVJPCsbHZHz4IT7x7Ng5TwYXvUMuYKA9OK85pOasvj5kl0I7aT
TwqIO0XUuR3A0UPqThv6bnK0xx8dnPun6dXvNxHNzgjGbv7SciRIA87SOUc4spZO
hBq4CW6N31gQMay9MramlOrvZaZB2RcuCu/P26L5NcxwTEuPDl9Ig+hswdL4aR29
iQwBJu+N3onFWTAzW8J/6a91dQ/GMUtIDievatcJvAeIAj/2WD5pQu9Yo3QEDsth
QWKX5s3lqA9KRs34Xb/g+mr2QspIXWg6cGPmsjajYMGtDUo/RkRGg6SO+tDLQy/6
6iBgHzE+CKTo6OQcSYAYY9CT1E3/ilY7koHmzyAqWWcaQ9hnbMgVtnNsEmnU+qYi
esTdGxGQmB9yYJIrDScSHKZkk+Qhoutncsx1LYnMnChaB2r5T3mVSb43v/2M/2B5
zk39OMzEmcTatq7Uhxv1xpFtU/t857y1sC+rd8lZeWBWBmFAPHGu33Y6FwrMJUNW
KoXwKpEPvADdS374qTa8M6Mjdhv5XlKi7DEcW+K+UvrkO4ycrDgn09P8aemj4iTJ
p7sSDFDxgrgFQGAol6ALAHSSL3gAr24BnCnEYYIUmXifizQe9VqP6z7rJFUH8fO2
DCqP9yEwMKhhF2ty+ofAW/8n/ibEO6AO5U3l9SOmS/5/RRZwZji5c85SjCLvS/Ia
b0EAouRtcJBXAciM8jU+9P1oKagdWc1yBYCefJlzcmAXAuoE3pKt6m3zFQnPdDXK
+VpTFk3ElBLCrfYk9yoYI08Sx5Ud20q7ZW5Wsygj082hm5Q7Fy3j3PI0wsHSfM0d
jfg+hI19RVPdyDFkYmdJ4HS9ppD7Zjuc/3jU571o5hdzS8Oz60cFE21vCVpyZL+V
2o6utkhOOpF99151yTqkaildu7XUdZCU8DX3vhQSQ0WIo6JTDfaNzSdPqYMjrwrC
+ruUuPum46YfMw0KfbAzqa9Q+Zqmq7H7DvZq2P2qGnOB8IYNgLvtmgIVUgh9R4x8
61InPqr/j7PBos4T6Uh75TEOeIC6orvak3dG3Ey0CCAKJxSSoFmW7J17dOJiFF4n
9Zso70JOJLFOtPzlrEqADoLVBY4QRCOea5TgLkI1TQatOYH9483tZ7ZYcW6yE12u
C4jC8Zn9YMI/DumqTda3pCqciSnHxY5RwUsYjaALdNeNetISXlxUu/6VJL+nSsaG
IV83raiPefeMaANMAnIqaQ4WRbVJloI571ksO8UZnFi5lbYE56NxIEBaWlEqXEZ4
dX3ggovfZQf9Pnl3uwJ5OtZfASJwFxzifzvq0P8uONqH4vzKOtE+Wqr97B/Oyxbj
vpcMiji4lsFJHIVWxQANQizh3wMmiMFhzJnBwCeIxHA9rZBJsZs5wCBbmOdMfMVr
VuHyOXnh/79AQyiJmQLA90kKjG4y3N8V6RYGDhVOp7K0WPR+QLvOBVfhpUi3dPsk
9mFdmf5x/4lVL+dr2yYe4S0mo2Wj4yue6Op9F7rxeExemq/GL6SUSr6kTXyWI3f6
M97lfNtff9IKn8TgAO8yyD0ptkPuJVpDg+wflLPHEIxn4Qvzic3svF2qsgSGTeuf
R4LStoPbaFu9rCKYxp5AC6c855DQg26o9pgM35lzqk0uB0u1HIjJI/Xjsp5eJSl9
NfTaf68hcpmjjoiBVhEXEYiZavxrtBtYySc6xzXx0LG572I+g/lHjeDD6aevQxbQ
16NhStEhCo8Smn56E4S+d++3s3/myi0Rs3goJRxtd3GZHnEEtCIpjQegebMKs0CA
FUnIRrxstgdq/cT2ESdkN7zkZ7CTWbjbRCJkC+dg+HFubIiOHnlItp13wCuihjm5
aDLorAG+wwa6mOiAx0bP++znt3wesVFO7Yg6UCKFmP6XqqgT6LGu7f+H7Hel/0fR
17RS3/FY467P8YWgkAJykqz5F095dn14OaOrt+Vi+c9KJf7PuCv+MBNZvflQBL+a
7qG5ukKPyQXI+ecLqBVjVl0f3NhD9SukJVbu06vUkeYgNrfknxM7PshZRYMopTzq
dOZZzBiGcsKBwjeNShgsenqKRuXkc0X/6MuBmq1rMbQTQby2dm0NWu49Sly0rJas
Z/5vH7beuQC6O4Z4LUJX5MadF6sVu9js4gEnFrdY4to+zSc25+T9iVwtf/Pzh+W8
aXBqk040Jljd+wVxpuZICNDS+dYKLv5kE7Xtln1uiiugKEJMCLz2K69nDFMscSoX
iE6OLxwC0ntf8A1YQIV0Ukyf1/3L3f+Cna2SY1m+VQ1ksufn6+bI3gt5Iw4d+c1j
fLljP4fCt/dxU+TRACg08lPZuRoMXfXcGx830oy+VqS0+wzHQYEm/WSomrGw88dm
/9RIQwJYNaBY5hONV443QjhgHdxaJ+xyeZlZC228oCdAWS9Qe1qmW+RScEB8NvrW
t9VYXfe7f+iPHJEsitjegh/jpnurrqSoXvkAgsRB1zULAKEtYzl0RLmqSbzyP306
L10hATBvIPKsfoWQzm92a8miZ8S+Ulsx2wsKR/9vjk/x9uuj1YKnn1y5HVScq4NM
oC+6QN1aB5HgAz8e3q5lw1plRLctaxWv80ztveDDb8yLWgVq0et6jGsl1Xxw40cv
wsFDhd3FkiZseEFX2aC10HjpBnqeyhhtwnvrmu10PqYmmsjwAwrTiKJHkrB8V7hE
e548JJsiuiByK21SuisZrfUcUoACR+lGo8LHxFYXN7E2MbncamZNYhZQTe5EhxuY
64zahCeJlYjZ7IDQHDQjBBejZwxitBJz5QKkrl5GiuAxgAlbUGO3oqPUsXu+hQcK
XMMXFGvsE32P4cqUtqJ0LSQ2tjz5JJHFbUgnYQPeyG4b+tLzRtwc2eWBvUKaEaVz
klBz9UZxkMToq6bkiPp0GUMpauJk5/3TeMNZJwY2877h2FmL9cn+MaqW5T4XhtdJ
3prD/V9ir5UkmUEOK7DYiRnwpEeIEzAeWe9PM3xB0n52Md+3dfi4aGtTnf3L2Wr5
kpPSfkYY1oKq6ON6/0UBKef29dUYmi7W7aaPkh414RZ25VGUa0V1NNg8GaGduaRd
iWAUpUUQlNhTuV9wckNxbm/33oqJ4EjBv3/sCC8n/NDtaZkpqzThrLsgdpGI4jXy
9GTcKIHwiNn6Ut/kqFck+9CLWXqaLOYehocP4WWvEDIFZFjjHUPSfOErs34G3wPO
cQdMb85olsFYE0LTdpKKIxPZyRXBWWFo/GZcALuLDUVMB/qUJXjK67QkWrMSqxMZ
3Vkkfky9m+jNPpiCoxqh7IZvHnxRrbFxD15PRMap7lmcdIf2di0VDLbLiMPMTStd
mA8vas2A2uYtCMYFzd44tjMkRrFIiqOzpWlLBDoQw8aeTtO2gh9ldX4kngL4Pqvi
WbGiRwPwSLQbyKIFVBKnKBDn4MZTUdVLXr9+IHfQMyGC3U2VzhS7VWRLVWLYAGPM
4O/5ukW3JVyL3YvwmaMwaqCVJdHCZBrYqzdHauDOw0Vx2UfWDBRqht3J4b+yocmo
aLJsV4qq0APITlLLFAgChHtQESK0d91c0aqzhL5eTBaMVgHbDdHlt1WqzxpA6R/T
EtMFWuh0MNtjS/EnFIvGlubqSDUx8n0HCpCTCspIWDtG1v6+VDkOr0GVBLDU1BsO
JISqjtYbwN42n/V9tZI+tU27NI0Uzp89nUKCSOR9XlaJNMqSNC2Ot/t9Lf2CWAAb
jsGZfR9UKj4eSlAHiaWGgYIdXUthcRtfwYhAqSQK6+ZmYMDfG5Ql7fpaEs3kF7ez
K/pnDsKuPokaivvGKA6STEb+QtzMSTSjHhuU/0AGyGmH53dseHbi6ZqqgCoSImTX
qrGD5j4rC9WaLTLH449coap61WpxKjBcL0AOnK0OCe+ToRZlRL6IbjNJoOxYrvXo
L7zVyWdHlJloQX499dOC2MSDIjxz/RJA975YaEaCRhrLqFPQ0Bg7Rvi9nB6BILdi
RmtSStKS4ME/38PYGUrNpM6cXvWLvcPbu/sGDbjIT6mCxKGuWF2f8W2V7zsxEk6I
xaMvLeoAwxnSPJh44BCJ+2gwhmPHMk2ucGKWxN+OD1BfTCt9WqKc4VAN7sadRY73
nns0+KO/SslGVQ5lgg4okjVHGQ+eNmcfoVMMKTVCEBmNYXL7ivNI5acbOKa4Tdk2
Hf069cqq2Z7qA5G/9RoHXb/S9BWNrRAr7RhKl60GLJSJRCpxucsRc+M0VxcI2zSO
AJlIfQjWojXKrjBjQu75rB0Ic7Bnc6qVk4Qqu1hV8BLo3gBOD7w7ccnOAEx1kgNW
DHgPLOGg745sR/zRa6TYHTqx9aHS0rXdofI2clNQcJiT6b0BA6mXKl6yRIN2a77e
gk1zDh+8Ce0GmPlVx95N5ZzjBrPH/u1aU9YadRsyl9CUbXWiqZjplhh0y6fZaAiA
vljxSVKgaE6/tFpNE8/TUIXZsvg+kPghDUbYJtrWkkUIidnweONKNPc16575js9s
y6J+xA7FPpxWjHEiJsmzS8uelUZshII3yRGAOdooMtp3vdLBvKfsjTtNggrwukqm
sUNxNLLcLUBl56a116KECf5D1d+Vpiu39WPg9vt3L8YlOX0Bis0AwoeuglXScsYT
EtlFlqvu98LOg19zjTiHiuJPWP2u6DmwiJGk4eRVwAEY5jolFcbx32gEwTn4bX9J
cOrjpo/Ie0O6peGcY1Xlov30vz4HZUPjZBIY6hMGYmZsWi5ZoxYE3IOn53w6FUO7
vIFQlQoIU+TPd4IRiS8DxLShQ20kUjUrjXv04UEde/G6Y4C9tKiJKBFMPX6h59/N
lEDwf4CmudI0WO1VLSyJlILQuwICqooO8IDznF4WVWmdfDGGKX9ElkmH3h0iOqHO
yiVFvsUFMGa0vuEp2e9yMbQkefhTraoJjCC/jcJI/zKCHd40pWr6+K2a04xCDkUf
ta9MU3JnU3AlNQOa5893C4R/hD02LmQX7KlWa1FrQIXWsBqiGxGKUFt8Sqx9IrmA
phEtgYvNv4u5zu8/OtehOmvSic6xXgfKnqP5tQDyq2fMCYJOU5ZVHslkqrT98p3T
ugnQwCrBb5XKAJ6+BzMHVvpQYoFtR11zszrw5KbMHtlnf3xzsYgXwFGRh0VAPZ4X
gbE9/5g/9qZwTTZGQzoCmB0SKQfyUDVccHaRtlrstJ79eD7l9f+U7v6qhWzIAUOA
vYByiFX0gwzlZEEubwqcUA67z+5NCMaIQEBxmKcnClpQUSQCGdsYWSWEudxlReYR
T9+n9TccY6RRNoSeo5l2VFwhCNOAU5II/Ih1OZSEMDrtsUe9KxLCRmMqXBKQRE9W
CGYB7gYXo6jbdc5Ip1XiB6UMqHZ2ozGdZlywGv9jqm1bJi8lBp/y5Ha21ZWFmzhK
GtQ8hN1HcA5EXe45H5CcGncdP0Ud6qJzoVegZ65NHHzorSaCksgAVckUldbcNe60
A5l2xPj5AsIdRj7vmFp4qSftDGo9oYryA78juqGSALMR+zYsl2aVoo3p5wRUD54W
2+iCbCBgExuwQ3iz8jRoA1FYnLDMWoG4D8Avpx8DrhbUZhITvy/kubH7h36lov1c
66ioQBz8v+trKJav0QZTKLVT7rwn+aJEYIGpIQ5cm9p0pozaEFNP2N5XXGHweEAI
BzG6cOmzp2PQz0ZrcuSi3RlQ6DeWSlzM9V7WoezE2bfkG/9XX18kIzFZreX135V3
gjEUMY7qebfulsRxVjcqM0zu6K4jeVWZK0pxDCXOqdBh7Rs31vW1UiKz7y9iN7Vf
TyH2T+Bhm2mp09zg+ExhOzWajzW/HiafvWGqq44jlI1Kdg55toyrGHw5eP1aEw10
CtWHhpmwq92wRhyeFuqgjy9S9O4OTwJGq8pfpSlKKzsJx62opeWa5cykCoQWvgdD
ElAbvuf7O/0GOLpp/rGrzbGwO4Qut/zc/AXIIRYCzufnwSgQbGMtSqgg5biXVZ/A
TaVVOEnikeqfXfdLi56B7vTPzNjfT88LI5cOXhuj26WtpVwEe7rRzXu3QmLmPzoB
AtpCkQ5E5DDX3whL42b1NJbWAf9jUx8HwT1LLYnbjhN0Ev1roD+WycGriX6Wzufj
igDxs7mfkNfHUItuzek9fCQduH1sTg37d4VwnxtPG3KExvUZ7DuA9xiQDaIuqAEP
NdcqQA1GO+L8FrCyYwRNulZzFS6Fq/kEb6OP6LZPt4HbgiMpkYMHQBfpkVX/piah
AkWwVxrgk2tiNZ39QqSK+XQLtAOMhcxXrhXUAl9flBql2ObPk5FqV4TMhb34bYPj
Hz/2mpxxJMD/7AACXlwHJNWxPt65YM4yEbQfOtbXHhYk/D4jfEA0fWf+L9d87oe/
BZBWjt8UQcqX5Gtsjl8lCDcNALlRBfKTlS9iYXG4PBPP8AlVHn9AS9TBKwAYEvsz
/rUIwxpHckiexrUBEfrBgC9Y19EGVJqDhbG8goOoU6r8i4ZybUE+JDZP2o/RCUMa
nIbfheTWpDFxMbDyCN3iTPDSVopzPKea4aNMiGdJqu9dUhwIbIRhznwX6zIfIPhm
FsSsyIh2lcR+xM4meO4djqryexJIAowusU47JKPrrHwvI8tRo16oqhg0WZ+G5fxq
ZGdRG7cnh1KDxDfIe4ZsPPm90tEu+eMPgStxIHgyvZbqtrJXcWXp+4nBRzX3IIAw
fYFGYzxzsbbMsud6TDOTrBUrqLDyjgFxK2tImipeZ92z1mnExxg+DdJOL+xbWAYn
u8gCIouQXPZeoyh2YiKpwVCTCS17+9vP7PcWR+AqX0CNan0UDQ+gaTM711P+LGWj
62ifp2h1pG6ueYY3nuDkMt5+EJIhGqlbxIjfhW2zDlIeo1cHHqX/1yaa6LhWhBEN
YM+bVofdMPJ8hOw+VVJVKX5pt9BYlMBYu2rFDiSgTfNoZ7Llv8vuqcI+T7Uoxhl8
h1EPM+NSHbcchDkTLPKNn1RAgDJ4u3RASFxT/IKtON0KXY3TJyiF0SEwHNDLPTZJ
N0OgCcjJH9XU/7X67g7AJdAKhk50f8QN7lcQDiSYQ7aVXB5X4Me49gqNMlVXGMGr
SGQEKSTdw3gM/+3y00aUJqkJTy4NP9dd8W3DmqqN5/8vZX4gWO1kxAFDCf9pzR4o
39r9RTttZLqtR3E7toCLX889P82Ox9+TF7fc7ddBqc7VH5VHeiQU/uHX3hEDOshI
eUs5m+HcEbWglryFJzHXe16FL96g+iOHdcgg3TwyiQTuWESmC8nJXLINgjtQ0EYp
uqBVaoX7OTMs/2sr3AJWDrvIIREIzXO5bAvw3vyW6MHKtwf0sTz8aTKmOmyjYx3Z
UL8z6vD77+5e5J21JkHtJfea6pYRiY57fDz0BWeUTq9bJO5+LMsniGcr0JMdatbz
ujnKr+Pyo7w7QJakzpMeSxGZSpXdb2IwcnDgzOjoenSlT3Y/Gqwc152wa28RArPN
FY/soA5DvBSPCyNx7IX+4g5PPsP1huI2SYJq2hudYurvtAvVrdSy1Y+XlV5ZpCin
nYlEEzJ7dYwSm/45KExwGFGPN8naoCGGZOcu2F9Ei+VOw/ohL8ev3iDiQ1tbLm50
l17sdVw6fNOWq6lqUkZIqiT7olTTvQ9F2YO3gTNtyDDmFRsMQyZEk/UcEBKtUCXn
eIgHMdt0CsNuugN/LO8D5qCZb4412ehdstTBqCOfSP4Xda71+lcgtDZZA8ypehIW
iGSYthSQNdxZdZKTezWxHsMozApBGFB+uCmFHg3WyDqfuBDMUdE+rk6fZ6SPiMyi
XHdTyL81UlhgJH/ja1+p8JXNKT1De7RbFFavRTKOPoo2iaUen0719kUCnlVkYqZs
CgoJud41c8k9c74fGedHNnfWnDFa9K55n18GpxbiqVDkjt0Yfr8gCv88NTTMnGJx
D53aQCeqyj9Uqe7L+glf0DiWqCCjnEOw0+7n5+Kk5ff4uZWKnEWwkJ0l6drUbury
RZEWBy+Va4wbyBSzVGaYWP8R+IqSz0ReSoHS1o2l1QHyem41/ARqEhAlPn2NDpkm
cLFmu16mtlBVCH7dy3TAjfcSujA/wAxpmMTrEbzPr2dI3knVFdxSq2JdEKwzHZgD
jsufDgW8zizkUwkAxswZm1XdbmCVzY0wAIXDzPd7B/cHougtv0YpW010oPa73mOG
kkve3G3BEajMW+8E/GGbuDGnTlosKKfOXspFe0j5Nuts456I7BaI4rwRIMcO7APS
WQm33aGN8cD8o2G1CKYEUaY8nLgXmpMEvEIRd+0XYz57PbjqPkg2I3SLHRAA8iq3
5uKUtzcdaxAdIQPy3XYfPYU0eQ8Lf9AMI+zn9vBDBybXpH07at1IqugR0OWJEon7
ho8leSa9pXklLqKWd8Zuzj3aeLPwqTCV8EiNvnwbE1UuajAmmaBNvPxbN79jBJee
J/ZAyCPBQy4aBXrp7kPyUOWASm9vLUK0eKCwHFzY/NVibEr/EbJzLQEJVRC9tned
/G8HzkRD/cdXfNJpZGGNj4/mM0tk8pJIq3jBFDf4B25t0uzgidI+VHL8tIXQuEjd
fg9VdAQCabaB4X8TR+FXI8ohklNltdUtcq0UBTo7DTgO8o1cxalDgkjOlVQTJk4x
AZC+Wj93mMv9TbeLYjD6gidnT4U9yNDN0oLuXmpjyS5JrN3ErcjUhU2sIYz8Gt60
AYvVmmJfwb71VQEGChyASPgw4czqmw1EDPd0qwe6bUPNl7FKaXYIM/TikCTTCZzA
JtI4b5btykEdby75kGzoVEWviBufOEcBWglfaLl2UxepxkgIfsC4Xs9jOkdFY7gZ
K3b5+2ZL1iUkLkKN+y+f4jJtX5trKjRBJgRe/pWOEtP5CLGKdLTvwigrGo7EbHQ8
ZNi111nzyNQ6DSz2R4bT4+8Zjf5OjYUNPazBnDwCWbQs0PRUypKe5w5KEScdvPsU
O9gDyBTu220IWf5OMkOsiZitSWpefTBrBwZ6+Twq2pbD3DfHG8A4TyMBpO5wV9dX
IHiNKKc5oftP1izmCABIR6NorZf+4NbSKtktUGELws6gJIQBFgiUFzHPdrrWzYk4
ZzWClHZuiLOmAho/Ta5SuhUsDHtUys7Ib8pMZ/pViSWMZdNiaYx201G4x3wQT1T2
mcS38vpepdE+9JMMQbBkFmVGwnF6NrDy5nPCq5rPf9McjUY4gSGl45n/ao/MaeKe
NGiMGSgBsvDk+x4kFZS6R/LM1JoXj2y6nsgKRscBHuUbY9y5tKpcgHowtN1k7X8c
PMDWejMix5lQHfI3FgjRezUzM54+c8enH1jiI/vuPP47f78GQUTS54RTAW1slAzR
MKVDTcrfJIIl+zWHBNRW5Y0UeP0LTR7+/TlFER+2MOqayticWeXabC7QhPkwCU54
SjGtdOaqzyqHHt5oy5akb66xosBUFT4cIVyEN3RZvbnPrI0a0v7HM4LrPjJy81tX
p4BJiWvk5byoZJ99q84kOQoJV54OoKpIN8jXNzSPFVGr7iuDKaWBqiXGxMcHK0UE
EIR7V2neQgYlDxT6MIkVM5eKacNuWKryIk57vejBl0o4o5/N1RHgSiWoww0Yqvbw
L7KpBG1rPWfbSj9khxsHRoG/SzgarFiSdeRVVzPe1F1oSZRps5qnKXNkQ29S6ysJ
keNe9wvf1H/uXrmrVMYDISLBYij/WDfpH0ge9bl5cDWrZb0j0z1iL+Uc6W6lyELF
gjcI2te8eUw0/bNVDTOv5Inp610diuO6u9s7iuCQqDgfNRGg4YrH6Ml1cF8AFP5/
4agFuyAs/AfZVzJ/MA7Rich4DNncS5MJ+hwVnUvAa0sYWal+9i5DnOT/pp4Y9f81
9+ZrUkFxShX+l0jJ4xfPOh0nDORKkgqTEcRXnUptrtWzCEkjQ8pt17GZ55th5i6W
yfQD1S8VN7H8jeh91CuFVP6T42GzhCZzWR9JJxouDlYWB4mEHyndLoq+6IOw8ge5
AjlWSDd620JqkvxqAtc65lgMp52nlxHeJBSBQ1QoslKuUN1RDOK6zUqbJ38+FZKS
vak4h3sewT3vtq5HDxizCp+cskWMSpYhUY/xVe4N1GdU2xYlFaGVvcrPUqKdtu4G
TJnZgLTEOil0YedR4PGTMcRuzMxdGLhLE4h0QJ51elwAJKaWr0nQDb1XZ9ykyORS
tqj+oXpzwJ7C3V+t7zLex7d3oMcPN/Z8rQTwCZQQIQd46FUK0kgRj7CZbyBdY7SQ
OHtBwjKetrst4XoxciU6+u6n5C/rnOECpyjjMMGtqwotgfa+mDABySYPssuLKwU3
DfEoQT7jabG8yHVHvGcEnppmTFZXhw9/+jaxvjzPfz5Bm4aZoUQqcigwNHXLW5kW
323X+Yne+9oPdWIoSK5wxjZS0cXTR8buMAcyGuKL4nuEPDrsrDFd3l8ZpaA2mQsx
SYjfXq45An8Q6zXyCpjKSau2cPctr6fSbVqPHTSOkdMr1arw8hrD52UagfC+a8c9
4ytDI54oiHv+oUoSt11lHvSwwVA1fmkh1qujOaW0XiKxQ2rSzt+1KUOeUeoEOLjs
lkRsxB14TrpdceGkcODbkRd70r3DUPtaQDFzGMsl2KqaJYzbRFW+8nX9Ea8CyAZd
8dj2ChoOju8KZ9Ru98n5aauRArllJYdeXyh+1ktHA2Ghi3xy6rGN5InjIDIcLmN4
2w/SkQw+uftTfmKjPUyuqTCTzEEcuvskGUDnKIItcX4ekBwxpkrpgpF3wOTXVwEq
ZrewAHr6fRIcHcn3xTsGeulZjI+ZVWiWZapoGhiGL22FcsXlYZEf6SitjJPzRGdK
zlLsix9iqejM+f3JUoSXzCAG7IFY1IeZib7jvDaCTPs3WSZWJO0NumAm8Hlz1UG5
52+jPha+F3Mx0Yc5NdABNMSNmnd1/WJPaBUd6L5sSeaPm2dfMy7ET5DLv8l9Jv3T
2EbPvceds0jC+LlT7/RK6Lk28zVfp3ECdh6uKiWtYxqnv1ojle3wWdJdbaIYrEei
jA8ilCF1PfTnGE0g4sKMDRRk3TiQ4N0ZBhUy4zFRdGPm66O5pia/tV/L7ryapSsE
0L+lIKaZW9wn+QwkBNZli4P7YQXdYIEmHrneRasvufeZy4YXGWfUXlY1cQmTOI91
6KCRccxMBh+/S8Cx+WDpeDvZoO5q/e0NoKUEph/5ZoagC+nme2B5SeNhgEXp1Ycn
bFSopi9A43JbE1XdZymGEJoJrKsiSV55m7JVAwim1I/uccq+/dd+ZJWEXUhJLc4W
7MBMW8ZMBXSN/rriTPzzWtqEV7qPppZRQliXVrS/jmA3cDSCqJzohiwS9k4ieNPr
aQ86zY7KAr0iW+wBHeH+h47QZXqUl56Pc4/JfHsmg4dRtPtdeFn2/T4FElXr1jij
NPIGr6doy2Jl1z7hpU90FahxztOAiNwFtD/gJOMX9w3w96TCkKirgmfOPYs2FD4L
BNngsNu2XwDeSm5gKmTbadtEplch7e/dj9Afv0HRAwIvMaEXtjOkGY7vasLtbgMr
WYPQDn7Pwlq02JyLlkkLD0abZrRLbYhAgKfI4dQRmkUAloQLgDQ5XIy4oa9kjmyL
tEvSOXI1+OO9CtHghob8qQH0xLuGTPdjmBxRJRyb427hPCA0tl+JBVpqrDJAOI8O
rnTqz2eZK34nQw9PCRgxqeR6OzRjTpB9CvUtTIUcUIC1pvDmOco1Rpat8xZmJ1C9
HJkCsvrfoZkAguIjwIHcraRLl1UbYZuXTugXKTdWenSPsDX7hDunkLYTV1w4DH6d
wc+s0cU1W0jf/IcZzLTSZ0y9VzK9DRKwj1VWIjKo4+WZ7Y3qTkCw2+oRQaTuM8z6
tHbvqoQg3JuAahOAwKC3z/OstNRXoGIClcueA2cHHoU0vVvSIUMxLvFYO804Sg8T
NJBBiR527QQ6ldgOYLRE92VDb1kmiXVkV15AL9KD2QoPDxdXMCJ5oxi2GaCfmhhQ
AVnhL2r+9aZEjcGnYiz4/Dou3iPH3juUZSWlKtu5BV6B31Js/Gm5fm9cgxwHTtOA
4jOkvO+X9bq0w0NqsqQQcxcTPlkaOxmKRrdxMFFxZKnfaKDVnQH7LG5jmqj6/NOH
JVt0ozkw/UKxCY2t5StuaMQ6wBFZ7JFk9mqdjnies5tGR1rluD6od35n0rKVaDc8
NHMSzbHEnoKpBu9sN+c61AhUNfrRYRaFGfvV+h8/tmklOJXHPS096cRi2dNciYuS
Oabng2ZZbDIrcdj83Az+Rk2EPUIjdDzzbxAap9Ue5JsFInZ1GQC3L//jbYpI4Zwz
EH6dbr9fvVtZ8xnqy0vW/34ZmM47pSGJVkwIrEJqIhP7dLHUlA2iYmjqesmJhbeO
GxXQFW2tyX3KGgRhUosx50zw5bPBq0+r7FuDEM50PXVm6rR6R9bF0XF9kFFvgjBU
szbf+JQ0LUEsBu8YDcI0SJJK4RK4JxFZFTce+v6bhFQOLiF6vR7Lhzma3wkBLdpY
vS4glFp5qkKINL+hiLRJaqftx3GBByCtPSPsgpkLVYlpDzSaANFP3TxEEED0LUK7
22qHc92Z64P8nlH1c6UWCb9+iCpycTdjNpdex9uMOPi1uEej/bR12voqKdSEa7Gl
PiQCKBtmpf8JtYk18GnQSqticvEgjSI74FVh1AZeAZQZ/OVew6w4ePsGFi+XzPbR
gUtF4FFAXhdMiQ75+QZV8XhR+WKBLMSGyJAiUBr7iqZCCiBP4k0X62jCEjvLPJid
W/gKh9jCMFJ4QZlzLVSNLHv6bMXYkX4VtZUyawlwV+tN8Yvq5P6UDOBc6EOgwGNw
s8cv93mDmf9y/Dx7orEhSQJZGEQeY3yr7WdF4NsFJPjTcApafwoGVxb71p4EJmgQ
LAE20JZ3YL+b3KI6PGpZDdifQo2OzquY1c3rKxLVxEvUdfTT6eQ27EOrDjzbENeQ
Nk4FYInpDClbkoDK2TKRDHNP4cVZXGOq56IVJihSTUgKiIadfldxuP41naaLV4S/
Uixl6A7h5LaREjJVpCBVMkAAcyOlxfaSMxW0bcEU4lWXQFJ8aDSXUVkhbD+Fxitw
DLpPS3gBY+Yrt4MWA72N/f2EwBnV+W8zMh/nBEcswSk3viLbFFyfiXWulVvTJOdp
Qpx7UdUSbduIQ2Kb6vl+5x8AZiCxH4dRV7GJYg23dHeZS08LZT4PZfTLh5QKkEg6
04fUAC0BuwDHmi2tLxLEg2/TSQKtKNF8g+HNRaG2YBWYmZmg07UsPXy+08kAFJ04
F7qL4byhwfrt4+fehLt7RvR8PIVeMC4WrQPxQYdBUyA1FQurgA0Kxgv7c+H8OGq4
OT9DBLjsYo7PuZ0I72vW7YoXc+ME8zDlX5vEzXyltC10FJytqn9p922D1KdJ0HnA
X3ZIdtYwxxxkfO4ZCDZQ3xVkbBJvCbRduyAQ2BHqW+KO2i7EaLEKRFAJ4cBEuRdJ
aKnyHVqCrOmGV5dSQTeYFs7H0L7CNQ5Dx3jPbA+5oHMj8fjNjETEpMpIKucME5sB
KK9q0SCthkpxjmdx8YG1aD2MH+eAjUVwVjfkQrIPd1iRDfY5l/+aA/TXpqRihF12
/b6C8IYIgr8lC8qVlnpYQDGKOTzHgru+UWebA+LVRYozhRF93I7KD1aI+Cg12ZNj
GLcbbAw3Z8lHfH1e83PPWqgRhxbYGu4iQq/Z7D0cacxyDhzZNBD32+9fggxnAd/w
FEDZGQZ0fSV1wwq5CpBvHvnN61A4fXKWk5EPMk52ajafNesnlXTPTKSOEYjkf4VZ
yuWnsFFy/8UbhyI3dEay0d2k1Jk7jyuz2bdXEwLipOdRAlg9gtOhhGp8+5rUAiE6
T8lP1OZzq6/io52m7F2MfGJNUhNBTRV+wb4oQG9ZwAQC9mH0KYN19z7TpbvXtmYW
HDW0XG0JDx6oh+vWHhi1Q85LoM64SFQh0+Vi0dtXoXhk/hFf1kkHCV3nZT6G/rT3
YOVZ6NXP5NAigM7HfTix0OXBl1gR1A3/nnHZBpTVTyPrb987CrMeJy/Xk7eC3gc/
7QqbWPb1TOlRGU3w+WBeLS6kX/Vfl0qcSSfSDtBwJAakFCmEudyfIEs94gLe1xjn
a/13ZvuKMmsYKdDMVYA5OuEHLFcE/H4r/fxu5+mMQ5ariGlE3LIPLzKczj286wgX
ShTFkOig0xh2wQC4h6v3rC+eaLgfeAeiKiMLWbx+uI23W829ndwT4rfmhLING4zN
i1P4uK5pod6oy2JloJmJhxWm4ITNLyGLis1TItwsuttIJUmxGSvjgZMCd56ZISjS
iO4yJjZsS4q2m3T+CQNtqjt8m3UzgVeV2w/ckRFsAFKkzRArAftXK9BzrDTpwoK2
Pwx4UCk9g/wiWIO34ZhD0Us73BLfbC0q5QU9RRHwgLJIHbbb1oCIJ9nnS/9c9Pap
ZYX1zzqlJNPZ3WD6ISdSCYICiHqEvugZBaHQFbX0JFJssm7YzXECbSE/PlPqZXlQ
hgW+j8kFlYDIawuS4ZnpZq2lOQ8E/OSz/wBDjI6YNfHK4Buzsr1ZsxDfQOL/Fobb
kWNH2gdLNP/NA5BoVv09BE07U/bMRETWaJ8ozAjou2LAC+7+mbaPj1sMx1FRzWsh
ju+PWa/mY2bBlztxpexs5erFYETKaxsX6GjEm80Vek7cgr5vhPEta7zjYn6Z9bbl
zqTGfJvSWGnEq2WlUcc6V74LAjnORmI6vJZJOeAKKRtACrQwcWQj4KNUBQiiFx1p
glnLs3JxmLGgkX0SnTFZKAHv0CLP9WzEpuOuXfxikq5TBvu2NrOb4Q4PVYNwq8hH
jTKOrApppcN1F7d5pVUrcb++iu5M0HcYOrUkrySQn7nSPyp1YKT/WWB2nKcwY7eQ
U1/Z8LtpLEY4j+xzh9PzDgBTn96oMJdQFrGD8ALbZ2b0qN6QD9mmyIbvFtaRqWiC
CR5WWoWymEv9WBeBhfRuOrNK2yNnboHlwEzb3rRrqUpxykqNCp7dgXL8kdmOR/fE
JomTpwUffrTsjIhsQzt8lXm/33IEe/6gtgk/1eUpVTgHqF2b54s2blEtl0Ti51O/
Xj/Bpvd9+LEFL7lcyWg8b8POympbwArMxz+wKGv9LvuYlcJ504T/lWSXA3tKzgwW
3EIvE3tmKNZw/Rht7e/ZdvcYWTr4L76SwnhaxQvOASgsWmBHVahOLDoszyz7DDHA
E+CF7jZaZnEMq1W0BGQZDgQV7rdCz3MQM61J/Xv24rWiMCYH84Y0cNPtnfdQ54TB
iCzFKJPUlK4687KY/JjZGb4E/lktvN/rYoZ94D0LcIVEmfVD0kJ9pud7GBTDnqwo
cyTMnDKS0b/5zEInSxh4q6z/GT/fnN9+FPPWUacw9EEC5IH1JF+FKmflbGCuDxhp
/LnwbQDbiXHLJSezBr8lyXemy6N9fUtz3v865IJbXWcBgIlZNOWWB4fE9qYLH417
giM72pFhMx6zao0uCSBsnKzRLaBMFR9p8w1dd4dO829v7S+N2Ylcw60r9WmfDtdT
zxakTiD+g/HfKBDQp++vkx9JYg6RFzq4Rh4OadKO4HNh5TrNFVdKYbZ/LRqrU9lM
KnOm6zudMIo4TcgUpky6RPsWbsrWQLhPMS0hcXuHYr9z5+e/4OqkNc6U/m5Iu9vc
c3wfjhwlw1IZpa6hf6/VKVOUXO7SFSnCr+xplzAt4+EtgdGiGPZClG25bn0UbE4d
baAdydCEX5kuuwOvOUMIssjicugqHDRTGXUp+8VLypboHLvy6SZPy1MOqk+W4VR7
xn9pEBAa+rfavcieIuF+2ITppqWHqk6ZNiDTNEO72VTtmGLZM/PKrEnnOqDiQSo0
sD0Kbx2+tb/Rqy1zZKDiJcCUQOSxs6pqVYZD5VdLdtBRuwm7H282xVAisV3LDjeQ
oq2kk0GlyctLAjuLH48/CaQ9nn+ah2QIxV410UzFJnmwhVKvuOShhydIX5OTh0Ye
TfpwTXPOwDFRhKFll0mn2HjjFVjU4bFPGjNnkpjHhd5DdFqaWLpUakavUwMftMPV
GZbJTqp93fBcRG3MO4UifYvG/2QaTOyhxk/XYujJBUBNUUcwznT45mahZVsm1r99
lqoxLSel6AY8HJZeAhCEdEhyEyY7oYTOmyydQ/YmRK38qoM1b58Lm0HbZTFxa1k4
u67yYDq6RheLHpe+sYjTP/91l8Zwnvyem3m8iqmXa/mdJI2JaK48ZrlmqvUo9tuz
oAkHBjhkuxj/Zjd/8UCgEailaJWwrxXZm6+qqaGbB6gl4PjxEpzDhWhIhf1x0KJd
RUngFe+yuksebQDSmTj++wVzzA4zFt7QsLl++fLF7vYdpzOAv4hStTintQbYXRji
Oviesu2F4KpOoeikQV3bZSgs80LDyWLyGGs17fyT+E5GmA7aAq259921bYSPNFhH
QCM+x2RxXbvXViQ8PJh9vF0qUgXJ1d6wkm/5FnGdSL5qvvyoq1OvQzJQcwjDZU3f
j3y8wWyZYoljgnTQ6I5WfwwO3L6X8nE0zZ2mfkuLzmjz2MFmdUWCuPtIHunHqEup
9XmKtxmFAXOKD4oEzhvdx7AuWz6lAd93wL6EPL4yd9ceTk8bVa4IrMZG2Xxcy803
3RwA5C6332maEXlWM3f9cfoeflHSyTl+GE3CE/D1f0tPxfGFcnspptoRBTduQrm6
TnfL2ttg2KQEtsS93EbHmZocUDXJsGz14EJLwaVWfAaSOULIFA9BOtXMnmdrQ2bn
QN6jbfkp9M5qHJslIH3yKZm/qWquxo6Dti1bT2YYq8KSSIKKswEc4jUxizJWTZ7A
FJFniN2hht+w/Y69LSdWUmBXIPZtFKlimfB4VZJ91rMQx9tAA6rCA5XAdq8j0ZgS
STPQIFAZrBpnaIc48stBBmenjZ7pqLFaLSdz/N2mo9P0mNDA8Ca2ejYMsqP0WyXE
ZL5lrXU9ixllriy3pESf4yXgteg3BQ7yys1R3p71op9GbA48p8KiA0vqm6SFBpGL
dDin7FptHp+3hkkC9sFt/lQ22I4FniB1OZxOsV9ydyMNiyFYWh2ohC+4AGdi4yVD
9EGxRKsM6gwmOJjB2XOuvhYXijZa7b1I9xpwMvhbB9CMk65OgmAl3EOah6nCqvUh
C4cAvvF4/EAz1kkZwKxpx9jljPJhAcM4fRFBmkLGQn71PQdgeVlRuGJjO0YEgPCS
2VOXSkrziu24yh5mxjlu/+hEX4XOUaMYJqtMXx218bNPd8fedTgGv9H5QQddCiK1
dvqUbrv8JhOf86/TWQ3o8Fh8dWEriIqoWs217FGqJH3If5GSp3k+Wif+Ba1FgH7A
g57El5F/lBWci5j8cG4a8ITTbp8s8uivE9WHKlSo3PjpRZXWTi0adWfO0L7/SBBN
Lj/khHH6yRBhwefcSty3AjFVhC9JngAp2QeIcj2KXWbPogQzKx7oKhlKW06vygVb
oGrv5OndBxHqbf5i/zk5XuWLy9+NiZRNAxjiJbEXiMF1PqTRp4l2zMbkeHMp+RBA
7oaZiZpIT2R6vDKdADlvPGVtZPU0PaWvCBjbhqbbkjEbvQJ4XdGK6eJtp3HmzCHP
U9YO1EvVgoHCzbq7yRJOCcp57/yom/cPTSZiuzHRApHETIaKeQx1LQRHJXYa4+Fh
pLnKeM3gjgJLFnO1yY9QZMvT3gcHwC9eRIWzdhJ4A83KG7jW/mCzhUwx2MA7HLgE
az4jh9G1WNBfPXF94GX/9q3Mm8MqzcE90BRDiF/w+v3I8X/0Gh23a59qmQzfzQxh
6/6cgdedMxia5WDFDFUzY8lNLtUY9/ApPWNqAHPhWmugaCf44qOyfWkOOJ/xES8H
UJ8Mn4uQNhGi0h8RIKzNZLpgNiBtzHrE8q/UPIAb8a6bJsyIbCqphsRXITeKtsG3
Z8V3o6WWnYO4xTHDzj2evaLiSC923TlzsXpsBspnq6fbViL56nCHzK4r9cnHaKn1
dY89rVPhV2Ukn9aMiv5Qvfhq4khcYYimBI2fZleznCBZpbj339bZxidwaWFUToIn
CurauCfekrruLJ2hQRfsygnNC4o5LIWPe2rZ+uuYMaaX7dA9+Ja/QULChQ12De5G
1oWA29eICly+T4vCBb1gQKE9Z6lvCJ9duFRiwK2zyNZBfFl0Urkju/FUALf5GhOu
kMh0GRzta9g0hVNLc5vHXif7stNdSQUqYkvhf54R6sqHEYsQFycwocmNAfqiaeev
2FJdQpozWYKQRN9CgU3lEO4GnnJp0aMiXFvRtgHYisYbKaFri4SQNB8z2Xx6KrIu
IgzHEDVx5W/VdPOzhq5r4MKKGeIW3HKB7D6JCA2SXrB4kTDiKsdH3MPPSGheSp2Y
MB3x507YkOaN+GRMCclIfzu6b7HWIldgOgVpP2wml9nSUN5x9XW3oJ2d5YVghE4w
RqtgSuaEPpLQU9XG76ZeaOnAdcnQAeB1qmCmZxJ0jvxy3rwkulCkhqIn/tO8jn3u
rNREhLpK1ZFCbcmb2J2MhfAhtNy5YiF+yny2D9QvdyAJMIlgnqXkwnAKAY+ANpL6
OCphJ1kNgBT3JiNynAklkdM8nCbxOCLKm/hBdM5G0g8Vtbj0iPTIUz0MRNA4tRXn
OEFcvvh7WX2VnjzDtAmqkcu+ORVSRVFfvy+6hNIy1HpT05Wmb8vZnbE1r5WqT0XN
86wo4Lld8z57B2hhiMIrSsGzGmcMmbELwFH6E71O5oTsMD4gvSi6yz1uX9ZPVicR
F0KumIKMbi9t/HA+cQA9+JHEFOZ1TNqlQPhKpAXnF9Pub3v1SdhV7taT8ouXxkKB
AxqGIoDwK2BRgP9dgqKHB/TKDg/YLkZOc7UqFdUw96fgg3vYeQuaYI+svyCgXV+S
FVQo714SHAHdlBkQi32hBti98Gyhy623GMbhurmpFhB2vTLLMsIgUel8/UPSo/uW
bOW83nXCv0tbvu+x0yqtu/Dq/LpMrUC1uBoJj6SnuaZ4DjJUcjopVpJCzmVbSSvc
krTmwkAb7qBTdENDLigdVfo/+KDkt6Q8juILrGnxA9cI9qK0BlLz32yN1+HO8DWv
MVWtTwIoPZv1q/qzy3y2MgUCwmccuhn8ixzMpZVAW1GrSWRlDildYpCKdEnrJsXS
79ceVWpEzHwKS9Kt2MziTpOpu90iC9O3zdvgUiDE7lI7/fyMF16RwncmqUjc7c4j
S7tsseXKMAlX4m5VmiC0CKKkMQMJeJeowEYJDXhY8WJ+NSNeSwzEMz3uI7f0Dfwp
EnmtaLLPn9a4YYN9JFpu2dZQKAaOHCCzoTFrYLBO5qSrdT32IUJHYlRe0BPovhQU
02l7QrxUXnGedU5wiHxyfMKSNInUjJ7XjtqtlFrrxXiEeteyFdon/0AOBRv6hmO6
LIHAuT8ykuQWzGUJ2bBPpmuBDISLwX7AU9bObEDinnDBOpnW/P613ztAfZwrIiYn
X6zD3oZathMtOusx6Kj49NT5l76AKI2eLVFmh64MC529kR/rodN3UqTZajZPPoJv
qQYQ8WBWlVjGgf4ZQSzhzeJVewM8HxcrsNjPXEja/h/QeGBJ3G2YFWZOkZNRcFnb
Q4Hl8oIK9hzOgjESjwoaMwWkcJ7UOEUXNCsVZgp826EEUEDjYE2s4c77/Sjfb83Z
tK49RkEnGmaqcGsFuVzXPsWnpmN8ClmZnH2bdTRfISqKky/aUulev2sK36kG8ZgB
VjBLrxyHFpJMkUvrgIv7l+/scam+0zAKv3qXgOSzx5mumKCz9QhPG7lQO/XoM+8B
xPKwRLocK3b1QTw10T6fZo3wulJImwaE/2wlBTHhbCa+9G1d2klCGCnN7uZh0THr
/c4npqIgKfuX3/KuKmsLwyH01ZQ8qFpsYOq8v2I7cZVo60iDvv6EBx4Zl6zSdbuF
D7BZJGLudF1D/4I/AWQuhEOf+F7mBSSmmI21Of0iH8cDNRMahSfGZznn6nrq2CGX
kQbTOHzd3S+UFOiHXS+IyBXVVxt/I/4TKemcoNr1ziyrr4pcrMI3snFR8ogcYtJU
SlwtW4EGAf6dRPHW8qr+wiVjlnqpAn7tnl1ot2BvlWPqiahvyVB24NW4V9iWbiKN
53xB6TXpX8SIImarLjOUaSa/AhZzqdIIEp3xJOVXFfRW7ej3SdgdeQBXLUIAFM4W
cAWca6SpKUTJKPus8dzo8Sfe5z21L4xkQ7vXP0XMMcMVI0EBx8pDHlPqzB/tQskZ
uce3uxOzIrqcOYjs9aRfiHb5+eEPUfR4FNH5BqPSgSjZi086EYGvDnLCesnmuMA9
6pvkEf4cL84Ue9cD+KWb06vjt7VJ+zD9tJ0Bigl5il0bIhazGUezlhIzTV2Y0F9a
aY7a1iKX1/gJ+j+mnwb+E1/YQf6sv9s4mYTfy3LekOj4V47TffVy4EDkvpH1OJN7
uBVqlAdG63wjXZKLkVi4Le9/BFDKIwt4fBqKlB3KKqbLrhrLsQu1O+2ZBQINvctQ
8okG+Mj2iNh8374ZbDlB0EjVwxpG7CDpjK5tCOJeiDNEr4I1/tcv3J/1Y2IP+EsM
Latfel3aa50cuqVDVTmL3IzAp4jJYhcL9gilCHLlvLaUeqbmt+PtpRZrta8Gg+Vn
yBYou7fF+dQbyXE354NuzqZtEbbxOh8qndrCaJyrYy9B6PNMvqdd6B+zZF3wlG9W
MNTqj19EHGiGqz7twNq7Hkww2mHvyG5oM73z6h2HUJEZ1tGMWCX5OF/rXEici9Q2
1kku8aWRz2WkVTDlv0PEUncEIYKt54f8YSrR4J/g/7B22RoCd/l553UdkH6JByJ7
D1ccfa+DEUP4jyH498lF6N5UHNa+X5FFVN9CWsrUKe55BKB6JBTLFapcvl0lIBC7
bWINZBAxlafgxDVXK/zbt/0TmeWpjoLXv6piowtj14BvzZmb0pK4f460eGIujzeL
tcY4g8KPj+J8lO6M/KzC5kcYKRW+9O3hOclwXCwCpNrMZNMFDWchp2bNXNOlWrTq
VjxVYkjZRWAh5NUbe3E5D94zM+Z5SRbEDfMw1cjkvMB92QILnCwkAK7OM6GHDVTP
QNqt8714Xl8Tr+nDb6OIYNh6irj29HTYuKAN/CPuQAIVDr/KQIxxIxXIFImnO8LO
4xFpafeU2+wpmFhyE/0mIHMur6OS49UhBmKggOjb/tQLuY8gAkRZQy01mGyuwK5D
EZQBFPrTW1CHJ6IJsXH1K7nxAsKrzXmWWufrn9CuMiOwQCMmhF2KRjcux8FGqUMk
u2qQQfvHVVFoXk7/rMnUgKeq3KR79tQfpSwCYpuPS3wqLgvWcGlln/+oavVGphpV
UyC2nKQ/74j0PjXy52KH0vEWJ8Mc4r5pMy+yy42z9yFK7pEL2d2fgZsb0JtEgXRg
C5Xp433C4CGnghPmQLVYgJ0fzP7BBtJ55XAwwVZ1BfUppj2u1EwpKRiWK5r8pPv5
XF7VNKAH5ysHKK61HqxSuLNFPlpfnU6K6czjscXHl6vL35jfY0ecKmcEA89UxnWg
QD9/nsoBn3Kf1PKnVG4K7ZWPQTV87YDRg7K/rk8jlcYwvRaI3k8YfaV0Iyy3/RNN
5kiGI2UyWk5tJYDuETOztpPDchY/LXm5wxWYcPoBu/SNBT/epmFXJRcJBzzoSZOk
bWXuxtWKz7bRPAgiXWO0XHSWbSP7w/EBTbXx/5XXp8Pd8+YvH9ps+PmTi085uSJN
0QbKlkUgJ2A8cRNMR0wBnFeLkg0zdXLinT+lvx6u/YQXFMWmXbIJp/9DH/K0ZTuY
Y2lGV1N/HRjbetCjHqWQalzn9DFdadp/X1PDbBYJ3Q1XDzz84lY9Y1JlMhSoXaWc
qfH0lmOUkQ5lGhmsCpc/bEr12M7DJCoXVOT41O5Glpolhag0VV6RSNuoG8lWNNhs
VXnbbvnNvX9k+EQG0SsXjG1twlyBEe1inynKbIDLXkCvbh3B9nBxYEW+yPirf3jH
d6fRgJyV1Hj+xhgcbg30PkQNO9PX8QL8+zpuesZ2VQl5RQhdNo9hz3dcG2VkCNQp
xJ1GwpE8w1zrTAXLO8a+IT9G6yxfFl8fIDDY3sfQ6zznF182ypuZTsjFlCamK08R
Gwzv1eGXq04VsVATT+6CN3s4FMgr9uZ/6bWsz50lis7t4/SzngRUiuNsB4pzDLbf
1tFKlTHU+vn/9wAHt2zP1DRLq5S9TPyeB84UwXStn/x1LP+jryBhHirEra5BjuaX
qX2YSGqcGGCCkQyjC0YbmzabzBV27CH7qmQ7socVAq0TQmz+VSMp0T/ZAMSUSFJZ
W7hhfKSmfCPtVHWsbZn+T0NYalNHe4LYuKc23gkXZKLly0dsk5Z4Eh6Wa9wExsS/
Rbj5qxw4DeKKx0DQza45LdVqk4WHQmyo48pKoz5ugKA4BpUKSE7V4Gd/QEUo0Pjv
PuFQmEBArYIbvc4RKTtGr0Jswb/E9x/RfDTQ4BM7/K1q8zloYdvZG0yyExv2gKGR
x7FfsbHwyDsGfEPHjAsIkT6LSEiHCbOo0jxj92H0aY6O5jyyq1C5y2s0H7gPXeWG
n7mv2E7+FP1Q1B+8AlNATlq6aHLW7QMDo/MrqdlM6zW8aMVNtEIFyFE/8reERLUh
F3oFL5AImYjaQxU31OXZjuNH6t9r+eLpUoCvf6z7oplEFCprVVL/WzRMB+pzGoe4
iunx+TvhptDE9g7sladcVrcnWfTQzzhYF1xCGOSq7H1K30Q1dm37j4JA7l8aoNdj
zuRQbRANKN4FZGHUpJAW61wxrcPtzEhbymoG5mVNBOyAUdLRSW/0lGiQZ4dg4FzV
iLQn3g2uPPB6XhU9Zw6wnvJGqFJKhgRPbL4tNgjg84NO9tgC1W/bdMdYUQbnhRmO
30XsRSv9gMJbUk7xzNd9UsKxFaXsH5IELjIBg7s0rixUqH6exxaIC2XEEPl+mdMo
EblDMUbsQ/IN0xuz7DRId6I3P98Xg31ZBKlNySUNWlRSJWftzHddk54745Gy3pMv
sTIk/+lZRNXa6EU4/xg/iuYFPcfux0JBlqFCqcW0ooBVwYI2hpFC0c1VpziIj6HF
WUupbOutyU8CeddVunkX9YBt5x81L4VYVm2xyngvOcCl7WzlnhMxwLwocxxNNZiT
HlBhmQQ5gWuiMv893lcJ3EsXhAE/JIJZ74xkOLfisgv8S07DEI6yKyX2NRLe93uE
7kBUM4cXkLbFEPZ27YXvpyuWFPk+tiOF+ABL9qoRIcg1067UUuGGZfH/97Mwuttj
dsxz0UlAvGvA935Og7Jq1YHGYTgfX6EUWNY/yWdzIEYgw0SDNZNpuUvwOZURVHlG
qXg/ePCT59Z+hVcqUQ09XicmSQ/jbO7yUCTTwjWK2OyzMwTaNJit0vh7e4xs35EA
N7oWUHC+qAVmNClGBiZbEdumZYnJOq5C8h0GVNZj5BJLXxIa87xPRMGyxgX4fJZz
i7ML7cl4Fh+yIQkMtwJyIIRJ/s8HLQO8hQ+pso6jMTA2EonhYa8EuppSuY1qRbuh
THYc57qSnGmTUAIaMtG9LL06cgWkJ+2vJ1d6ySkK9u1Zr7qN7nwQzdRGyACiVUUh
XaqoGELKLB2Q2szRpOMc0zZeZpqod/KVCD6zKvLat5rFtAdhsnsYGWjjmh2pmmmV
RqyaRG0wZkMNt0ysMaWg23X1XMG2Fov+kd/VASqQE7fThVgrrgscztpmdx44AniZ
BSwcwFb8DoeByzDhyRcas3KRlGP+3dyQNGA1WtBb3rkoJMiyX+CtX74HwNxEacYd
jK9hRVVE4m7hyEuJDqNz7yQRMMA0H0X9Xue/M+Cq21waIipTQEXIwihoA7Daz1pj
7sk7Y2oonUMzhqvpXfU1cxuk8kqSE8UFV7+8dkLCV3uDeAZaWYJH7uGRmyqhxhL+
/F33REOaszvpCaSQ6jjD8DisLTFA2X6AGJXvsDfbYOXiiQgaCeNdbM9ckuJJrFhf
TpU/WL3oiKTxySn8a2LbeEOWfMFfk0UX1GM+td1OPkixIryLBOPw3oTgktyZgZc2
1YOwrds4MP7W4DlGTB6GGsq5bVlXOHbDg5gBuEl1LzlsYYmYySYeyxWABpyOuCIa
QTPbp/gsU1DGlAUVN6UAnRVMj1tzK9KBfyZRWtAoKoVwcqR2Dq73wWdLGbrUQmRK
+KDFxT91LKKjDtZLImWys5H204qEAxMn0zZwRPYt3sF8my/w++DCUxFsbkW6IpkN
fKDuwcvuOfXFh+o0COc4IDocdF4hoxDOkucmfP1lsmu4CeZoEZWQfggO/njx0g8Q
IrTE07qrXY5WJo0QTdkqdBCy59kESByV/GeY/Q6RPrHk4ecEOoJ4/JzxSrUHTX0s
izsDsXkz+dgo3Ik5vhMjZyX1ZcUgpgi6Mw7nyBi+rnLswNnnDISGW3v8jcbzd3+v
bjg4IkGvC8h+f/Aov6qGIca3+85HS2IRkfEDEwk3dJuVHPCTOQj3Xa0ULslInUkO
ya0yqo094YFuHUxwp4T/7WBdgyoX5vDxm9dx39p+2Vo441xUC121EEBvVJ89ogoj
1eX3BIKtzqRO7FefQZnkJTLQ4rZoauixUFkSvxjsMx2/khoidQWyISWMcFb9urA9
GbMQp/tOicRmuUdRLh5zpdS9ZvUCZdv7JnrMue1gjpQzMpgsFg/38wT3FgGwFUf1
DcVgS5iSqDJao5hUzjuZyca9sLrWoli0n2XLE5/GBilWCGd9SHM6XiK8MZN4Gdoc
qFgOrFBoRfC6Jro7FhxGEACDJNPIEI7bW2yMf2Rd94KDDyHp4Sn1N5LeMNXdApQW
bdSCcKKrnXfdXVMl3PmJRDzsmpRAKud36NNJQTQuD+V1rCTWoSj7IY1lVqAnj3lw
IUPxrzjU0HFm2J8RuMCTevrqYMMoF4SEawcfFB7WOhBD/kCxbx0i0eExgl9jMhIp
7vrxDbB6JhnPXwE83wRfZ90JHJkssy70etM7PNSUMRsW4Xm5HDNwYcGOBPIjetT4
s2wIFmpXyjtQjc4cjhLN2/D+idWppsrF0P5sJnwDPvrv0urA4q1E4PiveMlqoApx
eJLhA2SMdAK0FskG2Hqz44q+xJhbsy2LSQtBm6zhgD54SERjCb3SwFCdvLPWIsrG
UxGE+HB3HHhBCWHyDs0g7Luo4sl2YkL6xT3Pj4l0ncK8zGMCW0D06/spyxH4D6Cc
HMYXQYf5BXvYvcaxROUvayDhsB3xpvVkO0XU5w4IaqKoWHSSFUS0HhvGdYgIRzAE
OKjKD8GxQvYc7jATnbC0Z1PhLNqwtOUf4PIjdWWmj6WGyb22tiIGRL4YMdcbED4U
j9oJF3wnynXKhx8xHp6nQE3B/2YG9U6kN+ok+p+zEcGfocXOmX26lSsl/UED0/jI
R1vUSvUNMSuc00tc6BLv518VBZ3Fg/j6oLj2QdjZQ309q+uYAM0LhXLj/gAxGAAw
00blL3hMGURsrac4Xo5gbPgE2JENyD+l1h/fEEt+uRzt/77qRv9Y5JKOIVDTTTLF
4ajnxSSO0WCStZze730+FqvPL9uf0aQYCUuQypSb35MX6A8y+dX+1J6fD+yH3hhn
xxbI0ag1XCDpjJa/5+78hoC8KQHpx3NKhUbH0vCv2ALrnEk5v4MCuLC/3PRPc5i7
/ocQDhvDXFysR9/gld8KSZmOl3fDyCFL8XFXYKW9UefDYzdEYqGS26G26CbYW1bd
M3vz9AP64jTSCtYfq+/ZWuj/xGW/dRkCKzYAbRE1scjlRUYOWZdX6E49Q93W/Poe
Il4iASEgwLD5I8/dPxwr/hKd87V+4STZSyfUjH6JsxGOMbVrtpkdRzFtUdb9mRtE
Y4ShCauvZ/eTeNgs8pPUMdY5F105GJ06GaEwqmdiB1uPNxpd2BZagzVLnk7NYeNh
Y/qnAGGtvL+Rew38YwS/b1A+RlbJNJQFlsceixwIadtpxX/X1/XfPEFHodHzZX/z
nj9S7uDWzr6kKXSbuGaZEUT4wr9WMJxhBSHaolSfBE+ND8qSlCTJ4c/PfgqQ/kQi
xpnlxrDtGUAM1/ZxHLucPLGLjiiIE9eIutgPI4SNW5Kb8pkZ40ByI4oe4oRJbkG0
hFgZ0DT5IV5xy00IUFw9iMKTL9wIUygpzRdjJ0e8k8idYeC3eU34zGhzXIurOwTf
V3I00ZWVsSrmxDQZ5+W+LZAw9VNyl1x1ABAioN1DnKxaPPCd018stOOBbcsYEkTt
/bdBNjJbw1dsMhcFFWsw0g5DbasvEF4gqHOJKZpdNh1ldgUYyBV7IgyuBcVletLc
8OHu15DXnT3xTx027Xp6Sbr1o4punkEo+2Nr5/I0gQz/EORYfZQqEBSQb7CqDRt3
zr19r0/8EA607GUNT+YaG3O75iR8GY78e0QDxrGWqhyZy0Fb2OgXlLhNrZ/zcmfe
K/WhLwaGC/hvCOkB3V3CAHn4uWadfrdmpuVvHrEYKnV6jLXnPY9GLuMHB9RCece5
B2/DMB+AOnfMPjBrbAkap2CQsrW8QBxg65eoDhhyWCL5C00FFHr/+Uj+P/dNQr/8
MiCJLE+7Q12EPhanJmdLItdFmy518F9mlUg2FVu5DQ3hYy0aH1qU3s/ButACxJ4B
pB19puGImeprmAtL4SjtoiCw0OtzEo0mwSx6Z+Hnvs0hzIGytE1KibYQxUq+G/S1
MXOCjx0DNpfEwSMpAtHJdYu4bWDj/i6+TmLVtY6tk/s57HEIHMF0oM8XkKg/++mH
Ed5tN1nygxADG7kDQo62litoFqyW9Lga36uUE9IJPxWviOtlC6kP8PNQMF+fZFIq
buHacVdfVZkwp1MjaV6gE8kKXJU6H+PAH2FhuM2IB3Nfh9E6Leme9SKIn6oYJpZT
WtKN1iGrCDjktimVR002ViaIEoDkyXhgoUQHGC6rT6EkGt9+4LLZTWiSQomdhfeX
K7D+oNeibxl9/GlRtSqdF94Q+hxU568ez2rmgC9MuBB5kFfxZUFf0Z1VhN6Ti6c2
Y6/aNgxvah1vK2d4pgCL34JeMmv10o/2YynCt4PiQ1hiTLag+0bH+17lncjJV6NZ
hbsa+27JANyPGedULkxsPLlhobJfQcgtknkE68U6ByHSsZOSaiQQfo+kFHVTksnI
B3fYo8+eENARSywBvU56Fi3k7JFJPMb8SpZhT4iAyX4xyUrz2I//TNt8J/racDcC
ljT3tMgFWhIZuYY6WAPUBUvwMfXdCkse18MRvV1mgaD4q9TjSNTJstkV9QoRZLZx
wCyKdbX3qjB3jZLGZjJMac/Dq7hOCq5jg7O/LHIGfGEdkkNdjsiRfuXZFGKwtHQN
+T2OheRg4AIr5nlecrJZNZ3YsLuD8L8HBgzJG64ISx+kyIVeuG9m7TAoDNOfLUU/
ma1udu60Zriy9+UR3aYs8N4Hv94xr4lrBFPKZXbRSwMqZFcrJVXSsIrtEMSll5KT
fNg79kbVO3SHbZA0GBMCJ7v2FCvGqRsxMhBCQQKHd7csyHDt7Y3sENlCeel3GRmd
T+sridOReqblBJMA3lfk03h4M6fve08Hbq1QHqLf+lG0baQlSrxTjG5QE35oOZti
P3/Q4oRCqphnjxxdHSt+z7oiuuUxMYKBWybJ5EH7NToZ/d7naDkMY/0wZ/M28Ia7
2SioLzBvs4FSeixDovCrqTymNXduGpGw3XOfxGyTh4ytlS0c5M1brpOqUYNrlSD1
Aq9RicHEwjnjqcuiVtwe+OGJ1epat5i9oHD88yU+Q7kPl5BsIhaeKrBP1AirOwTD
8DKHwHKofxEQXvMuWSY2yepa7hLWr1ianrrVeSvQX/Fj879g5JKCTdbyKlKf3d/A
9Vd7aTdDj+Dzb6Gsyg9Ge5h/lMmpTFUg4BT+rHiTrjLZ4Eo4xEy4EPWPdtIw+fzT
XxXnD9YiFuwkNpSmTlDzAbMJqJdN7nFOwLlSSx2ahzioFcRlzy5WmHFS8VJr/LvG
RelDCR58MjJn/6WUVI3GdKX0YWBk2mFs7N3tdCfwbWi/3Bx/H/o/t+b3EWgF+MEA
tXPAj6BD4JOj+s+mnM66cTo0TKwZi9/BWItruDpp4+aHmmzz9lCqqXfl7ouCW6ZK
i+4jpCVtDkR4ljNGwSPLm5ovf4ICRb+JVGvrw/jSG0yaG8CCLI1VbPejUNi3DUG/
1nma5PQnkJIBPBFzHY526ibkNeMTF3YcAsx6+EGbbRrSXiPpBM02pgfg07LcF1tg
tl4dPrUXl36SNKmsfFvu1nrqt3JY014uzbMhmLI2CnvnOpcBwiaDG08FBJQpmB6/
vnZkbUsya0WpOv803ws3LO2iCfIiCyx/QiPlmJnhJK97rCKq8XzaMaIv6mpOCtOQ
B70kFHi29RoAepK/CBNWHeFyLkwUfs5+1mpbZuZEOZaIfANaJPzW0fzuSeIoYuKb
Pa4hXPqGZ2weN972pyXExeQvK4o9LAHt1aPn6euBbrWM3KFWrLj3faXmXXn05T9M
sB87cmn4ehiucYFFDccbTl7hXYAfkkCfsmSKSKDUSAlcl41CIqvhObfKaC7OQzGl
8TEVESfy3p7TYQpPsvb2a3WVwAcq0VPoOYDRYO8l33/5df2Yw17smv2RWLzrZORz
6BrrdyA5qipMGeHGgyK9gBz912dLEXyIDNqgsMZBzN5TOZcdkTG3uetPV8hyKqWG
8g7YoXY6ZmTzzi5ah6IuQAhMVTzUCyeSXaKGKpuugRaBm7MMxQmN23cnSgyj6Ol/
3N+2Tn1ZiDzJuBaXjCbtnMU60i2b/T9pNea+NbaNfTWon9uKlupaM0iRBdBd349C
i8oSmZwXooAlM7CrR6KULrLIJTvcJI8Ya9iimFcBWtEUH2VYsoC+xiPqQEjJefRv
m8i669TXkV1tPgoHP9M8gtwQrASam+sbRDmelVijVswEfo3z5feJoTDEkrt+l6gF
n7g8Kxh9uCbUC0VdMJVV7uJ5k5bFhtUV+gJiQziyfTXpRWOmnaHtyBg8ZMOkIla7
2/eDja7XgzpfZczKNihVOySdtGdW1oemQyt0HT2Hs+kOOlyhSzqhaKx0K8RbugEc
hjtAA7f7YEJVzQbOSvWGbUpRelmf6OmayGJSlVdl+WbXJr3G7stbKSAazXI7DWbA
k7c2OM8q5a99KlxJAkFZlbHIqfLNcmhusxbpIk0YnvXVm8CgbdjQTpQW1FsMF99S
9nM/fpfOofX2Z3YHkDMwaKAO6f0Un8cAa3vlWEJkyz3s8ZrXkXS4wxoUR4NKt8De
kbfArkJ6r6Z2eTl1LHLjuUsa4CFV8q1Ijwh53in1PL7BiigEuz5TWCdjx4JZFVAO
z0nZfnzhcZpTF76ZS9KvV7iDcRn8jUSAovV7nrVPq0AUANzGiienj4XKIdRFae3Y
fxau5tTG1UxucO4SZU63ceTlPHCINKwfrEfhVy9Lz2ln5oxeqe1AM5YyVeIKY2qv
y3ug6P0Vjud8uNEE4o12JeP+qryazFGBVzcJNMZ9gedAvENErd0Onlu2lBpzFJfg
PitjUXOWXuFSRkK0KqKlvQLNJmlFzvqAZVyI75gu0/SykgLzpYfxi2Yqe8/CFxaG
h0cP2T4xMZ502zAsPx/elf9+Y8yiAAQ1hMKtryAH5fTeqpyrhbNOtxXtssudEtDC
+CoeBtzZ2eVrShkDxYSXgEYnv1DIHeRcU14Hr5ez3WgoCHs4vEdBjaafHBs2gvyL
7zupZJ51koeB08U0u5xPOV6jzR8DdzHpbJr/7tmR5Nn29DSeqNMG5XCdG/7k2a3X
TRjBIRwZQl6TFdOW7oZDQwhT2YKOwUSD8tKF7bVAwonjfK5+6D59XVHVlp2O9Ugd
C48AZkDXCd/+fgvom1dhO59eM8tIWcNID26cgka/8SChq1M6uKxEXUWDXImQCwIi
6VRovCmwm8NuOs0By2djAjEZDHbRY2C6q687lWvg6DUMUuNweB8NisqlOYD0brVt
wv1lRIKn23iv+CgO8IijEeKATNYUi0Ahi4U/TuhZV4g21jJaoFX2+uOBha8dfd+N
6mJ6EZtR+hFVTR7+egXfXLVuXF2ssp6WT0nImOOO/EuwaZlaDbefZXppSguK4eZJ
j+LFfzA7r0aH8aoy7dHdl1I0/y+Rc3pNDSyDwsobEbcDfYqFNP74mjkcqx0NzwTY
5vLKQ4+2liyZIyFHPBARQ+yC1iOe0cxfqO4G+LkG/hvpVb9SbbTuySpE7FqQp2MA
eIP5XPQ3/zePgy+PpkRnSRZOhPTfqznr8b96A4jJlr8OoFDw+b2XR42ODnF2FKxl
vRBF83ZQUCCyjQQ1urGX8YhX8KhdqzgxDi6UXF1YMIyfUSqUlYbEgG/q8eB2CpnH
Ptlj8F5fMEDeUNS0pOFcmB7bJ2PmLIZ+0wPo8mSOO3pa77WlzgEpPXO6A5it23kd
T5O5zeph4PExdgtJzS82OZxznvJFo1qR0JL8iUPqCRJQujDD9vgLKtNanfkB+47i
zYnm6HFHbsg2Epjdw4kn4OwrzI/Yk/od8tOt1wbYFEsf7qZ//sRVNsIERb3SSoq0
Hqj+G6dRAY1hp4pK0v3TQk7s0BLXLifrIBRLG8kVo0rxdfgC0juShkHXnPski9D4
s5ohqPoRZkvaqCIoySkbOpJjaHTureKQABg9SCiW4ZA8yGgpetEviyh4NJuhH9QR
+p8LZZFIH73OcunNhdLzhPp5XBiJWv6ZEd9P6sM0UmdCRO9bsq+cyj18qi2racfm
H9ur16cr7GPm5EVnV/k6H6MpH4scT2ZGSZ66RCp4b3+qp2Bsq/ye86nGbZdLyLRo
CNV/+i8KWScqqpE4GZhHgbb0zUgUcuOy5bgfbtFfnqJcP+q6WMzM2hXhFCkZCZT3
1ibuTBUgVmm+dusxEftMeDN5oXOQ1ZC6+X1q5G0EoJbGixVh4W9nHMw2Re1q3LOv
5KePUiOPcynDG1+pcG7lEIMjAE+Qz+auDEVYN8y2M3Wf729g92RnvaNR3mwr1gHE
qiIVzkdjeLrJvg//IdIgVvaNMndrOMriy5zVBeFgXBdNmpYzrQ5h3Yz6hAencwg5
clLBeqZxC2B6IWaBxAmPLewuT/JLxbKM+kzsFXFtnWubbiIB634Fbf7QJbxdwd80
2l9cdnetNi0ivpS7RXrp5TzV8mx3Q6niNLfKICy4BTbTOc/aDTMFHf5XPoMTs+uB
Tso4ZBMFxSAX4KBO8K2le9W3XNKBraUnVe6UjnfXNzWQeeqC7bTOi9nxI7f7Siq4
2HZuInp0xmw1XAPLEiWw4OAbTOpdzM4Hb9phL2+dhr70EfrCc6SYD5OZN1VQjtvw
EBtsb+emKRrbIZ4I9mQpV1PKy1lIrtsAGXy7zimJ+rBsR31m/BELlt2LN9Ovw0sc
uF4wzT9pVkibFcO4XmbGSASsxa4Da9cbVk5+bW8u/oGREPXgXp8tHOXuYqdlcadh
/oRQk5QB3xrSTR5WZyzz8X4Qz9qc6Xem8rhxB1UVbl/bi+JWej1t8Adf68O/EJFh
c3FE8OrT8Kod3cIIYz/vctBw70vudJKpx+1O6NPtYgMUeMp2u6uoIALrBgQk9O0s
QJvREE2doFdTD9bve/5Ivtbv5Nv/GfZVAVV5O4y7ceiW6Hz//f/roirDnidsyVGS
t8xzIMtoAHJm2zxWppq8r73NjfmWvKvS3e7Xr6zmF2hB25Mf8I6j1EHhuPYUyubb
IaXNimt+1Dh8bf+0AhmpsqsmwWHuWw3htJpPT7HQztQa1kig0GCIwI9eCmXNT3GD
T8L0tikua7hvq6FIp7q3OLsczz+HXBTMgJ8LJdCoK00HP/WG2iV0cvRoPC1pxnS2
FjtmhyYRbOTQLYJpCdh1/mYsxWC0boz46Dd7fflFRrAx1jaOFzLDHuwjh4bW3pf9
6fjVxOON5bfSgcOCE5Ui1yPTdvKRH7i1mIXe2m6s20FadlidjaiwdFwRiuSBnP+P
LmOv7UfftH59JMAu/GIddYEwsXRnQmkJK26AcMDrvqscEZOi3pJe2WD4TCgYHhrB
ut81QdF6P/I1kIjNE64y37WXsnNINGH5TvVn/ZWL2LQG82NwAaZaJnNhn41P/s/V
IFaQkdn3nhKCJpTY17TnIfl/odnYcdcgY4vb6rPxSm5BxZT0BBjfBJoHw+dCJUMy
ODB5xuk2OHh7LejFegfAi34ZzhVlVUtwCP7dDvP8d2tH2it5gezrWvv3nXOoSFNR
R4gRre6qEeNAKQYpYhhoAG8EzMVSQhmg+K0ajxJLDh2Yt43uAOAAkGvRI36Oaz6H
/OjZZ6Kc/OnSEMHBZP3vMtjvWSnsLqmgDOCpTlSmoXQHssyZvCgbbGb/H64fqAE0
EuJ4j9O1+MCquYp06Nl/4P2Afa2REsUIrwlab1o7PqkryT2ZOr99/2VOj4NAhXT9
mCnj6uwOwJTNE+kj4K/Hzp0xz+pLB2exx3TA4oyM/DoknQvraprKcHrQOfC8LEbw
+LpO5fFlNkCYvLVVqtGqisDhmpvU+Bdm87sBtQ870JG9Zy95vRJgJzk4g8A2wtjl
TiGbizvKMFPeFmJpK45TsVt363HPVhsF/XlAWXRYMT8BqsOmK+A9hBiF6FNXQRNY
7Qus5mMgxlXd66aRqIfJGaBdE2J26xOZtC4AJCwvO/Ov5SQTX70FBYKO4nb6Q5Z3
fM2dvNDuVcdRblA5uEk6aknRwwDwA+HHGvMUcr5dwdzWHMJUkEsuOF0QesB/mZpN
uPvGatm9cSeOmuajNQ1DyoStJS5+D25mmzO97erUCNgJwNBqzG1tVPoyoA8V23Cw
BjpDSftz2z6ZVHXNyqmA6+63oLzDhvuXUL3eYWWW0Q8nFyEET8XIZmjpM6vYbShn
tKXowMAE2Dh4aE4Ge8mU+C6Wjip1qkXKGzDEUqEZGlg1usVYMPRSzbsWoWTtHF9O
pchiCW2EIBky55LnQJ8e+1wxPekNdkcgFENs8u6rQM71uBlRiDFrPa3nG+C0K8yV
foQQWxXjvQNhKK/w6pKY/EbUuTsg/TxkQF9FUox3VBpQZ4DTPYbllVuEYv3p6Tey
bHovGtx6YukW3eycMd4kyBTUD9jkHSW6xfRkA7B1mvg4MaC/dcsG/Qtwx/FgJWpu
xgqImpcqDPxi0l7qH4Ax9GCpWPuMmvKFwEooVZbz+qlrtvD4qA7NsL8tElCoHmKf
BQ6qB88PNWzpIqxOmoR7pCURhPJp5v/EsiOg63VhP9cpycowSSuCLJyal7qP95S2
gyjLvR+RiUCVwoBnYp7okYigv9i4jLXbLN0xFt46izKtlE2FeG9chhTkxrtZtQtP
7L6bh7tPWC7Tk2skkTpM/Pxf2YC6fMZy6kl+2POqyzfjS8IYPU7dfFdJlA7pHdvd
w2i/G2ZnSnNHcbx6WmREnqsdZjy7kO0IR1e5wpTbXRGPXOiQneH40CTqURUSc9wy
ora8uOOLBU2xljWbpEORKKhHSaOgTpHHJvSf8HGAtlV4do/5nRZMo5E4nU9UagtI
HCfZTquh5x2sQ+wIKMVyCc0UukYnkSGBOE+Kg1oodd29l4bUcH4s/Eo5GoWY5qMh
587O/fwXUHWIZ5+/C7bYIXeUwmNxTP31B9yLXKNIBBuNaIbFm/2MyhRpvArIFSF2
GKBgsFGm3yH3b8z+eo5hJ8RUras9cR2gwsEySvhBEIRX3lb4Ty8IleLOKqiJMhHD
Ni9H+WE1rGnxIiexlrQJlHntTbMtE5TTwTzy79i9zD+9GOUFSQXnpjHieAmzbdWR
P0FCb5hUshiiUDIaLvVNRrLoteHeTv52mQSSjl7eHZrJi2AlXPdxsEv+169FKzVr
gOl106JygU+d/JBlxjszqnp641HcAjMkkx4wNW4AFfzXjb0IWIfW67EZ9YlW6bLt
Aocgxi5TIcUlm7S6PTmz4S7HuwkJlpD/qowp3JGLHi6Unc62XZjF9ssrli/jAlBv
zgQCfsaR+wks12KWYUdZmhe5EKIKHIc0eUB1eKMg4yn+r+Apk+3R/E9IkI4OQzi7
NZ3hwpeyWZNcmVyIJ+Dki2s47zSAnIYJr6URLxwdtnNJjCDZCvyXLJ+yRa/MSt9D
YFlWmlPwai9kIWCq4ztBP7c6FbdAM15BX7O2ypTUg1s4VabaHoNNreW3WYiL0tV+
3fTYL4suf3W8iJTK3dV/lBZVvgd3AhSNTt9wJzVf/aQik61RS50+Fs/9c5X4PNuG
sKuC1xRTpkqau9+MxHZSFkyfzntuLK0Rh6c76K22XZTkPTkQmJ95Bd8etg3+N7JS
juACUwCDYTltsPDHHVlOIOajOxzrYBRjnr3yk5U3pZ+eHTzWjHPBd9rNZ7I8sfz3
kr8qc8EH3kVr4BlgGOrwHey71Slyhvovzb/9T4ejlWHU7m6E5m9/Tkjz+z6Uop1V
jzzhv8u9HQUAmqdWWW6ueBuGrcPQ0PlqSnOVDkabF3rS3TAKM/MTNr/RqzBZoAne
7/KcjoEqmTgKXyB0QhOmPZxWswoExeBSTGIpnXcpyZWijsFV9khF+AKxer+BRbwI
3QFbZsj8wKNLBHJn2r53weWqVEjFYbn/L8AgIABA2vr6VdxyKaUPXuMMeIpfEs1B
jtQ9GBs+U9rpn5lX0bk1hFeAKiDJyt4fMmfvcxrfVh61z42IpJT7oyJoRaQzUDrR
vAaHoC76yXdBnYBSao530DnRuqdAHMvYJh3u2vVsjiypk9wPgCskdr8OhWERKko2
L12OxrAvrtASBkUOCHqSky1wdz606j3BC3GYH6RrLVCxs/6ZS4jajHLmc8lAib2h
4b5CHAsx81trfCoFpJqOFGgVJEvn4gfcv8keg1oP/OCjEz8ezPgNaXo7aG8GCi8A
GBQtKlLcCpsXTsEQKe+pv+Q9mOcuZ+HhQmjxk6DzPwawkAbe30t9Lc4oZ5pTCq6i
fuu27HYdqCGvc2xWt+6Yl5QRS/LFftULP0WY3Gqf5oH6tNaf45fvhHeNpR+InMU0
EX38jZ2BcahFPFqGoW4LTFbWOnIp7fVYAY0C8pxOVEI2hR4kzuARWY+L7454XDD7
LF0w8IyUHmLH12zslig8vtqnqLsTTxtv7gyVd3bmxCmZmj55ILqQbHIRjqYg0+Ha
DyBuhP3Soqyy0PGwNbGyI4vFhDwuj8XJuLDuJmIX5O8U1iL1pqqCMWX+O+0kwVNY
Qa2jyhmjzqNk4a+y/kk/bGjaAIFOaPspT0gdr/3ENCtoBdjyUUF9KIxNoniNR/Mf
sTCuJUzBWPJZEcvf5XNKbuJXwzT3ptsntNPEFjcM8jNouAJJWp/Odi84LLQpE+hG
TTzpNbf07UhUIgEHrsREludC60G1BFSHL/MjOKW3O00iJiuCaxba1h4Vq2ZVxcBE
S40FPNyQ37I8GuJkG3yiM3MbzdmeS60Xw1dtW8iACNQOD0SsmahdtkOjy8PtICkS
JvCt+JsAoYKRw6EO4KB7zi8hEKHI+Jqc7d3HiiriHF3qSv6Ll4tF77zdxkXliFED
D9PKZaP6G5CwgcvVPkRJB/yZjh3KR+jYx3WUmKwfOtwvagvTWxxjGhqwWcC3yFZy
b9fOMBxoJsWy4+USyq3lELIk4W/C7Zz/h4xai0oxOP+aCvyhm71jR/zTR4rhYJtJ
PAibkUK7sAmqFYTEs0f7czUbX6rBjKv9k5qPlcNySXHzwaXRjR2vC5Ag7R6gRb2B
qxqjPnPDVl9KnJFKvrcpGP/tuGM9wyvAEKB+9rCCdBJ17VAVRb73DkUcftUdq819
b3po0B+atIhyLl+idcOKwj6LgDTuJCHND2tQWMz5CUyHdbDbuJsXPDkbDUVv3w44
TL1azR2Aay9cj1838/KDibF/XG59XGsDbP9558/+qdfK0sPRrMQ4bCqEv4mXjMLz
whJ6YevU6ymfTgDCgWUrSjgqJpd3fUK/Z6IulB3jlZ+uq17UMyEFw68CfXwe7orc
iBHwEBf3HtzYG3HRMMejVFxS9+QdXf5DiyEtvMgWtrbHX8VcP1npjXJ7z8Huvwso
6buGAtLcqW0VzgZLlz1ZYNIvdjUPzjni8jlKIPd38mFj0z6gxgBxGyzCC5LWOvb3
gzmC2x0+TUrPt0E95ZEwK/g5s0u7mhTVGrm2GNAVPbekCrCLlKvH4Z64JRcYYjX0
k0GMCN69OuzLhKG4PKmKJv2ZBM3uq/F+fIapgwj2rtxuHj4rF6gKDtxS1glnIXSC
EGJS/B3pbqaN319Ns2AjwjXQH7ZcXHpSuu8AQreff8ROdr0diR7z7hTV/3WpO4oc
8K13knBvEOeC7Kv2RBYlp9D8egyVP2HTVhFiY/qHiWV2mzYkub8SZvJjv8zSFbAD
tqEyuMqAK8IimppfRLFyum13bDXy1u8pMGQ83jzP34dH+qxBCtPvSPEIjFDL2EPh
jUNiQBmRFnHIDzdsmTvJcVWERz3bpbD2K21CylVJ+1KoiK/m5K7+6mzGmzEMk1Kr
ULcp6gAt1gbh5JBjbfVNLarbQJHThVhjtub+TecsFqRRXgCWZsnS8tl3D+VEhRqN
TX5P+Eg5LbwDus6JENO64m8NKBk2KOBbCqyfblTVjlivu2VsPyzPJY1lmmloPPCG
cYP9rNaHDUbKDAz4zoR5SlCD1041bOhTUG/u+V7PCBDKPuLINiENsgm0wnat3EBQ
2OHczzKy6ly8V7EKnWo7MSGNi3j50QL5aZljQq2AdpK7JLc23eJ+3Pdm7gdhT9v8
Swpyk7iO+WFLWu398B+exMp4mOIhkFPUfi55458UcrlUrFHZfb3Rnb98TBwAmHd4
PrOTS4FEX3e0QgJ1X2wLFCYrdf1yZF8S0SJy77hVxhUeZ6ccWLO2XhWvhbMEDyJp
jqWibeBSDkB2dZWwnh4zlMJ+Kw/ISxFr25sSzZ6A2wsUWKgP/p63bLV4LqmQYTpE
iaiSSEke7ZmamwIEvYCypYlh0SKKX7cnYWclp5AxQ4fFv5Qok2jPfJ+0oE9HSmP/
c8RtGBdvF9vqBPAlBD7Nc6C9UtBEdgQ/gKOM6eIlU4P/hMNdA7T9oV9RrRseHyiN
G/CjEOGCiAu62dqWSN8nLHp7sLDCR2bk+seqwR3UK0o9hNyU9Kp4T9ZolH0gCRHf
CwtxbhRABpK8y6jsqNWy2bMmJJrHuqDWxACA/3qUdaYByHIjFnNRIVVTbpRnATWj
cif0+FKUWV5f2qszfXPsLHNPXyFNzYi7LbGSdVGYIp8wqVTN2VYiEHh0/OrFPlB6
cmGYJ2FQdH1oZiJgx1n0+EEMWWoUiJh+O1zKNqisgAMwhCyaCVkBc6cZI9GHHUCQ
2EsAs0KgG1TWPHPojPBoKE6A3Ze1RUn/cD3XUH/COZ+WYog5LWdKiMw7/w701imP
vYtzNl2m/VBbsYy1Us8retu7/kQfeUcQymOOUWK7A1i7XakTh/j3UAItEXfJ0r9t
Zd3jxPeDiSgOSyFKQKtDF9EeBhGla3NJBiiA8cgWGtcXRqBgXxXs54cxk30IRWjc
t8xl3ytSSXsENIDS1TbtPj6gpzJR0D6uqDJbWk7mjvAadINNrHYk7o62swKfubgk
0ZnWI6zocL88eUEuBQ7x545cB9Kp2R4HsvmlYu8Aa5NPGP3gMPwXte/zUGXnIOGB
YPyi3/hqFcuv45ibmevWVPlZ8DrYKs7jl0wO/1atGzQ67XG3Bz/J/nBazKx2WcWL
FdlAyIcstUlnE+ibUAUxt1ac0BgEUkIqKTgqlPXWAKVvf2U2yA85e1V5BmczVEyT
JSg6fIXqUTyY32kv2pw3kwhpayjQQfxoGhaTCSzs3zFIVHiO1NCHpJxMOXONmKAp
j3mXXEaRmcaHoUKJnQ4dNcKt+yhRjxlBHjm/BwGqtFHl3djItAqSOoPMvdT+WjzB
N40ZRrw2wTY7u5dT3CXm2g+7xEv/qTEnCGanT263aVWJvIxRliS57MvIT5Fld5ei
4YUMLhd5PVi5dqglsRAH/jHkXADRbs/ryKwy/FhzBiz1btEfnSyA/eGtwCBO7SuJ
DFG61ACCbTNh1x7ClUnPkqm1u83AdcpA9n29fWXS0JqIQKZaJLC8uuwHRwvNFEdi
COruLB+iIzOkbDg716a3DPOSF6bL2smqMkaXotM1X46vLq5cveiTw6yK0O9NArWa
5+oltC6ueuxB68ODg/T2n3+CTul2ET5TKLzMzmu/4Jv5uMave+nMCZIIYKcltsjJ
GsGg2ck+BaeyH8MfQxUzjvWcolYhmnsXQaUknOOESrt45hW6SN7z6A4xmjp6gRcM
ODVfaNhDACnkXEr0rolFmv5uzG8uufae2BP8Bhc1+5rM9OeK24/tB9Zx+lBSNu0X
vQItVo0Y/RjlvYpyzbFTci1cF8ATG5Z+fwCCWt8pz/WL8t1HMIMdKpR5KY9UGmCN
x0AxZv6Pew9zW0xqZbKpo+13Lpz4U9y4Bq7CqGhBUi5D1R7Dh+3zNxA/qw0M3UGu
AK29/RxYk0W7iACF+Q+yqhZetUB24lRARjNYdGS/j4e3Peh5F0H9XJdjNK6/Np1h
+JWxXF8yi58IAo0DZm2sypDf2aNdv8lqCN1JWZxip76cjhFf4wpQk0pvNhiod8yC
YOFVgSQ0tIumgLqoyaxncsB2hURTOBXDcxCJFA0C7AqFCJCtJLYXKMCjaBhK33RQ
MEgHszKsPkqk78hEJoDBz/H+3IoBZZpAuLJYHPtxvCWDAMNf46MQDxGq0fbyrMCN
344bEXerugVO/4eI6Rl5uM9Y1y5lMIIQH+z8sF5wZxgSYEJ3viGWnmFV/rmCTWC5
eKmL3nIvLlWCrRqtQP4W1/vIjJKHaJLvqfH8zxoV9ZWnK+h1b1k538ucT3UGL1dp
FN7096gKgWlFCzUuncwnqp15VnzsJGSq5MPZ47friZpmeMHaHDgREVEIv2nYpHms
v1+7TBN+hsKapG0UWRRXwz5WrfnikllojABF8VnlDv/L2madRF8xLVzbd4E3Lu+G
9ORa1GSalLZaBihYdeq6Bq/FlyA/GOcub9Hdx2KPz2d401g7J7koHH1+I/qwI6il
aKEcAc78LfPX64MazABKVu/JL6/jjEPGucvahMdJWJgpJbksdO5mwYjaxKeRh6Uw
s5nxobHfg60Hi2EuSnKFIXz9vh3SRRmZmCUhA0QrHgB7qV8VdWt9MFFv9FSBPEoZ
QT2Azxx8/DvkGHvQG/Hrc8mKGtGIyxOQ9NWfO1gblEm/lf8xx/hNaFHRzAjlC6l/
IEulwyily4B/JnbUQ40Gf00oqgbF6/l4BrfcFDJ3BZOt9Yl/k4m5mr4MAnW+w0Q0
lwkHDBsl6updHc7KWboUHaQ5+bbfWu7ns4vJGqZvCvfR6HvXF4HvHTmmuLDMctIZ
0ip5vexJ02jC0ikCKoCt3mblsUw7boVV4OlXfXjEh0dmGJNNZ0ENY7YiDFAdpS6F
sKjDW/lXFFumMGlP1S8cJ3lhc4pyzypgHcDkfHg88RxHixR3Dsjdp38vz6suyxnO
AwJk9xXbcBhYv3UAAnF5Rk6oTXvUzh0XeBZwesRWDpeFfx4WQdA3eFjvD2k0K5UN
qWieJxeQDDYAeGl0BeJxsEI+2IxcCYQLUV1I1ihwgJBVxTRrRHIacEYlUxY6AsoS
q98WuBsjx0j9yMsad95EuS0GcgFJSWD8T/BaDFDUsw7c2D8bUgHllufp99HhYybi
+SjoVNS2WHrl2nJpL8zD4ON+O+a/MyGWi851mlzAILoT48pnk3cbRuFiRfSEkyPt
cT5rUlItgzvABRXm7P9N+kWDH4RRUD4YZoFCpQhIYoE8Ll1uEEg7BVbjfo3YO9vh
HzxEmKYjJBlbpFdNmm5KRuCVlyPCd6KHmcf+tKuqBkPzD1n3eeUsdmZ8Yf4kfOEf
I3R94dWVUG64M1/BiQJiLb4T5YOdx7ehUyw2cW5D74jMdTPlqzTyEm8nseoSAlkE
Hl6KwolEbmvhJuYSdaMLwma3ft2V/XAJsiXt55uaNb06n/GQmy9yfep25bif7/Zk
kX25aNclhycWEHVdX2o7n/cVnLA3LaGOru4gitKLzC/6q77c5ISurnPx4JugTcso
iZOnyi/v6Qn5pGLPRxNHUgld3SktGYYtrZMJ8XLIb3cqQmDqqzUygHXjboAxtMwn
kwVGt58aydUtD/Ft/jqAY+4/3U5soldfK0B5ukkWJMtYtsDXbaNuczQEcgft7ope
WCHqvIwit7Hi8AwZrolpH8BqgKmcdRNGjzKwKTo+ZIHOyjwpPhDHJlyg2tdC2IDh
GFAx2z9HwnT5mCWRVUWENViJxCV8/Y+pEK/9PHZTYA1QQkiHKbY3NmOsSevGyd1Q
cELaw20k0eyXVwKdfDoYY/qbwoGLzeNRjgHgcbDez9i2pXNcflYeE+b0uVUrpVBm
515xVMdYaPD3RF+k0x3oMqGMnqOuL5BVVTqbX0dUIWYw6IzRsZhy7WXwJNUPtqzK
4aajtPQw0SNWKJD2wZKVP/29azfFng4YVjsCnjp8J7ryI1wv/pt4k0VRX0aQ5DTW
HfdP2S5SINW7EpQabf5xbAi7N0txSLsFLdyItBeCcuGtl8TXmzdZS1C5ats66dZa
zrPWRbFT5fs/pVDwvjCCu6VSO2IyH7i9NZm8EmhP4XOXWsIh40AlLjNoij9iqv9/
wD1nHIWnTfF1qCB94+lSRQwfRTzv2LyN1Ak7DxewNaUcGtnJ0H29X5xPlIin+V0B
Uh/06HDS9VH3ptkPFzqlpJgA8pO3BJveq9iaV/N341TTKcf0cZU8Eq3SRn0G9S1j
6jcoJVw1asC/P5xArjKUCPnjdp7xrTRsuDZTHTNsq+rMZ/BWwMkc2rW+f84hVZzU
YjXMxaHZ5RDiyQOeT3sH7Hzd6Kv2kFE6+i0De8Eb8Hhhzj1gSyQ305RvRrW9Hn8F
aCoKqK3uf2QmqU3PIj42W3CJGEMqhHVEoW+nu4vt104eF9AFwui/JnJS6Fcf/7C6
0a1DYhfKH9O/ylGiu21863g6IG5kMhPHjTCXrArNPAmH5PkMFSDw85AolSo9grCe
j7oChUcgPTNsb5ILdov+lzhZ0nXIqMhTwuA0WYhL8hAYtggV+AIKHewRjHPsx2TK
wMkMlGYVHz8u4aOxStwxUfTUWFAYOu5g4TnNKhoLCMbl8rO13CC1duHbE4DEP4+t
Ht0/lGoN67MjE8+o/fYg57O0n3iGifpkMmbRgUhbt/lCakWyi0qwmOs+1w3nT/8P
OFDlSLV7XRRHGqSrZoesZNekdwjggyo0oitHQhRrlJ1Mc3u/F9lB9jVv9cIr5T/n
EnZlhhYwtyRYQsoP8yF/+7JAORUohiv/K1FhakWZHyYourVR8AhPxWLLsF23wKkk
n4qVALX00DQ5W8Bzgr+kZoh0GukW6MzDAweMx124AeuQFUR5VG1EVMTqUHgCrRro
m9zDvbKbvYAcaTViiBEG79KAbqDl6WkL31Ts3kCYc6yOWe9R1Ba4ts99NVd9ZRT0
ZjOAxY/k7jjQb5jUZ4oHN/TazevH9D2KAnFPht6g/grTxAPkjcW8Fw6cBWgpWyCk
HEhsWRvDzK7hLtxQDK8yMCuIo0vy6MqQtJxxYC4ZDtOwdVIU7VUoZQ8n8u3Xt2gL
1NVcq9aEI1TWXuPVm5qHbpEAlG92ebFPla1i5iaPPowIOPbQMTh6gEwijp2cqXIa
lxbFm/GO9YwIE7dOkbzTUVA0CxQlQjg+OuBedfPiC+z5SUP9becUzirsdvOcdSo4
qbp3yIPKUIbN1jVgAFbHoyP2LPpGuVnf+elKoHHiEVS76BbpDPWXeWA8GvLZdwo2
Qzq9SS779KQoXWaNKNkSM2xvcwvXs0gmLPchztlwCgLmyKKfcWG1Stl1o+v3MFHI
GJOOPpL3Ct5CYV8Vn9xLeoRA7YIwcZXMaCm4GZpZdRgQo1YsnZ4ZkAOdbBo60z6f
XKGuI4kPXmdt5xSMVTkJWpCTKmMx+KDn0abjbtMGixm/CYARLDvWUoGVHCz3oTuW
nACkMCIZlxSEtwGQHmGCT1GxXNRN9mUm5KXPWeXZpWQFRRtM+BQOEt1Cog+fzoVS
9/hQsMnJBKLVRI7h/X/KD4MWjRC2AOVRFr+4Uyg2CfqdMIeEAXFWcuEPc38xFmMS
iboLimTNUkvUbTBi/nwFDRc/D8cyj72VsygMqm6+hBzNoXB7cJyK8VcyBphGLXsQ
IuZqGWgrzV7WENi/kPd4YezGLL+sC/GCiwf56XcS07OR99D34pBcJFzSFevvb0k8
FKHdDT2kTbLpB9kNQhPe1Hl5mUvtIDNoMtK+yoe6gNrf4Duq/NJlrjnfMQLEUUyU
M4bnI5TYGtuURQvGLia9D+aEMX0uxWRnfqNNaJmDXhw7Gg6omHYG28fMPWFJlI1O
ihznmb5FSnoB9KsyPf7LsY9ZG0h/6Ia6S+SpBzMN85vY16XePaAcDRFufPSy/Geu
irvicrW3upsREHNdT+v/CEb3eyfsqEfl9xwRb0Jn0HS4UMrWOv6C4EjBnqIF23HW
zHmN3g3lCdaEoN+VEZBYjPXrUYjY2iOvdv9g0AFSa83t8PfwNi//dem/5kPw3d2L
5994XgIYo25nx6QEPQBlfTaxG7eeYyAftqoIMDEC5S84GsTT1b2GNLq9UPcoy4vZ
V2LL6Kr6k1Zb67i0LLOIOujTRi5y6PEmcEy7qBO284GO40teT6uxcOQ+072oMZRQ
vmqIds9p0jXkDVVMduMHjjWeOm+uNBnRjfxAQK8+YMZXVz91WHk9aZar3svi6um5
2OhuOkarOWoew8EX4n8SALiLrmDe230lcLHh1mx92mVywHc8SIQ7evQBgejD5z0l
3dCXetlxH/aICxME/Jltqdf6llmZlUjNm1tKMAmCm8EQ9KTwc2yT1aFG7pFxbRTv
A5Ohi/oxbI9mSQl4nTWB8fztKL/Jjdv4JeyOkRxsLqyEjKZn94OrXEnYnr8Xeopy
DozmDK2UxO1G88zBlFZ2RsrsUXUpOY3Cbo1sE+o/hGzIfRHehbOQtiKahgaluiDZ
F5s17yor4Gyo2NOO1ZwKKcks+wLcOLcfWoLHYlc5WIuRc6A3Evr+vvZsKliRz86M
rHVTu1gk11ls2zjGS0mJAxa0TrFP+FXm+PUjxweYwthbMiNH4VZBELaOnTXQZNWL
MSK+vY9fJTPSReHMiEkDoHKfOLi+m98AAdcDJkL8Vu+n3oUCIg9lzaW2N2njnryQ
2hoWWpxLejB73BVHa/hdGX1lUH2TJQuRkrFq5dEjbCPJWSIsTpeiVsHVsmCsNmSH
KWLju4A//nv2ZkPY7xa9nuUDCigsNBsdX3DQPe/va3iH45FVmFvVurmDzY8EO2Kb
Nb+afFDm1fXw0CqhNqXDHK6K+xOn3MGCEe/rO7+bchz0oVnG7riHhcBzrc9yvq4G
oBpI4WVcK14pl1aJKEM3flQu6lSdrYGtOf1uK2blJ0V5dYaRWiYzkUzB9ckl3TLE
vCtvIqPz+YWZzgXK6Cqb2KOwk5SRzX0i4FcT7d7BGQSdQkcilX6Ozy2KeL8TegQE
JpJdT1ad55jzhGs6YET6t2hc2aJDzjm2rGNb1GnDWkrBnLus6H9R4ekBRjrW8z3Q
5Q4cB68tcA9I0Wt9OxvkAM+cbGjl7SYn7vBrXRPId4VErQU8FxKmmwkow6rYTHxf
OrwUqW0KEZqD2y588o+wQOJo9ksSqwCd+q7odaCI0aoLdYvX3MS6zIbt+BioDnIu
ZmIB330367bDtHeIMrbqododSFSQS3oTF2m0eQsBzEgT8LiWx446pKugaQ0P/Hyp
4CnJ9M6XSulFpDSVxf/BZgJ3TbGqhFqXmuaiixu73wCvpI/OvRG2DGKd3/sZ2j2J
+ax0QqFFyvjnwFw7CxJAdaIy8aDBFensaKB8Sd+HWFXV0Q8Z/rWKfoqMVMc4y0Lm
bf8xcWASECJYq1ABDnLh/TZu32YsHngXWs8zXKwnpOROPsxGSrfVIvhRPNG5t8nz
mnWu49KteYU0Sm5IfyGuztVbGSRmZdQcNUNMyNeq1g/l9gncLU+s8A4N4T3ekL0U
+ANabaLdNcQa2nKBJfoyGSwyGykgxxqNIAsIR82F9mYqRCbCVOO9fIsurf+VZSQu
VtiLxfwxTqHGUhmpMClComYZ3KBuhova8QJOX2gD9S7Yc4RQy5uKXJHZwj28RGmI
LtWitA4b1tmCqYHl1umdN7j6WeuoUTZja7z7ZHup5cQjkyuVXiVpN/juWyQrG39v
GOEfDRDGGHRk5UV+CfqAF81rXsU6i04HKOHsVy/JH/tfryYPoWQvZSplo0jGFqug
oNN5JHsko0lIcbE4Sf0QUQh/cl6NkivHNiHjVm3zH0c6RvxT6J5s9Tv0qYFoTJyq
8X6iBLJwjR11oolNvUl662gyJ0fWYFX6AWoopJhrmtSl4OJ3iVQIWzrb1S0M+tyZ
+EypZR9t1UQLZ0u9GXJlJeEYbR15KdvfwGKp4cqED7BzC/GOJm1W3cu6rXpcO55a
UsGB3Ijt7pnfOYQcHejDQM2kzYXRwO0l+DlBzhHOMX0dYDt/pttzzZwjAaiBNMD8
9yGZbESJCG8ZGFZ/4Lh61LYs6yokAfRbgOEmIPxWN/qmt8XcKG1riY4WfOe7p0rO
AE72M2e4NFCrRPfrVqKcOjHXgzZXZyGYgjUcLxI4AfWaTxO6m1cvJiPHTiuFIZ1a
GSwljD6Lxjk3VtoXZrg0eeqE7lUfBYhcSqg4Mp+Mu1jRjo3xUNtiw3RftJNFQdeA
xgqMlxTTHcqjVSC3MDBW4LhWM3LI0wtqnNnvLPuFJjo26WZbSyOJAkQ3xER20Y1o
jM1A5PWqochHH/ccl1XtMhlP4djBRTSakaqIRl+7hgCZ54i4TraxJDNoZm85uSrt
CWqJYHei/GfBOAhLsh0Q7v8Gid8mb3u1XenIGwYBys50ePg/RR/InLiqXn1QIvjh
Z/Wx1UNkzujELu1v3SSpX7T6GYMZ0QXZfkNLIXjh96cP/rPyRwTJHmtnKoZMknic
Lc0btdRoG5rKGY3q5jOuef/fC2Al/TxLH8VY9sv5SG/XtdsItscytgENroLCpRHQ
3MOw2stjwgTW0RlHmhqJq7EZKFnwFT7UiHBb3Sjsl59Lag8Z1xvVDZJanOrzUe1/
4jFzuSz5YDmqSx/6fe/TM6kZCBzY1I/DV409riyH0d3pSR98CwYcZfzdQk7CMnuq
I5KvQnzirnQJ881tEs2t6noSX+D58sqVDtyiAjUQpsO4vMExM8sNOFsJEeGEk42n
VCjSF9hxnWw2vNXe6oBQ44sk8dmifMKmsUVVXrWUyzAW4NJ5/vHPUsCzNYsOu8HO
GC7wOb5l1N5ZvtGK6gY76EPnZ/4ML5l/W8Jq8OYfDNcNZIcmDlwQUBvbC8Hx699B
Ku6y9Gcf7GYA+nMHB6TAszi/Wnp4fp7/HPEXmaTiJVFI7To5mDLVCLqXrTp3S4o5
Z0VpsRwT5Fl3bxqxdIiw++jZ2vlanMwjZ/6zzTpE73bXgmQj8OY7ojcYf23Ln1Ad
awcAiH4yqsWoApYyroBhFaBiJlSB31LMlP39IW6s+BvwuoAiBPmEdvKM5Cvno/ol
fUuhxmW4aUdIWUL/xkCh3l2wXhfdRQ9z6uDhI+cqi4ufPhnUnFeNN20JWeN2XX2Y
2v4l2Wm4vVsYEd+E7GLydxdWAOF7eEIxSDP6uYh53ipRZK8djURv8gI6NfRyecr3
IAaUiYWPtOvBFeERvZvuK0MgUw1oryfa6frUYQpuGO3cnYBWbJw0COpY2GlYSVWA
ENV5I/leazWI0VpgvY7kQlWjaQ8CNjQPF81OVucUG3c5lyriCJlYHM1imRaf1zsy
eHTbILwy6duS6/ut0GwxIP2zjgSyOLSJRabeslyz2ztBg6ve1TeP1hw5j2Gz93DT
aXF1u/hcC9dw1J7Z9qbe3uc+6VphZl6YoOmXAB1chccrgB9sTfiwxEB35O5HWYco
s4ZBhZvB8iiMCsrUYMKnvGtBf0j8jtc/t/7uk0Jph15jzkHDj/UNI7wcOFi5fYGW
UW8/Y1lOnrmwZjtqzsBqZldaySfo2ILJvVgbYVBC9aJdvfZoZsgp/T4Us1S1+iRu
Q42buyeCb829DNOxhRg1isFKDNf1GSfFymHSPUWcS4yXPy1jF8nIDpR9wmzJw4sx
3TJkLXVpYZp9XnImW/DQDXDAOXDEbSvmsfFFkxImO67yDNZPgTS+O4p1dRFBBxy4
BtDQicg3Qm0B11FKCkU5DCtL+5/BwObhTIq+TqxO9puXdXiUFwK4McztfaSL5qUY
Kd1kAiMl1MN2E59m91EfIJrmcIkp32Hr1xgxcBrSV5ZRcLDs+h0HKrF4bQbXzYwv
ky9c3/jJzIh6TfQsWxlU8C5dgXMrXGSEgw3S8AtSgBSB6jy07Vt9Dkk+7akVUlkx
FK81e8zgIJnfu8QWYmbcMGRvBTnbEe+1qx7fCmoxoyxUAGMzhp4GStb6TDH2aQvF
aDdm8UxPoylt5Y8bpH6n9iy3uLBvI98066J7V56FokFNFKTg1vlkT0bGQzpkdz6o
QU1kl/7XyXVt4a7LSqL+Bn/u+NZVHbrnZ4HbIJu6q8Et4BJhJUbnBu5ID6qRZ81l
JO3E9DOBJWEV0WKgLF+m7/W5D0kttBbIaQsabT9gAoiHg9DJqq3+ZOQZH0NQni8Y
iNGtBeqYyDgS/t8ZXXC3sxvETF0fBzdkbZJw2RKXNPqjHhTGTdXJ2bVbgxFNxB1H
IXOQUkoLKj8rlBtbekBMJq1/sXrjRBJAUvJNUwNTKudvAKqCeIWB2fWdQhegiWBl
TTevxaU9psRF20IilBmPv6hdSeHEvXujGicmPHiEqW6DxO+gSpXZOXdRpqcTyyvV
posfBmo7BaaWWKNReG2EBh0/BxiLMe02OwBwXutCWPS9sKPUWUqw6qBx5wBO7o8w
fNwNUYPNJNVxwiJpbLAOeuKqZqo5WZ9zFEaeqkIPwEYO61HbYjr1NXXR2nnth4Yc
1zO9fS3RNrHYv7dHOUOn5WTX1f5tbEdh0eCsCYsALerAKXN2aEfZqwbe6W+4GHvH
zmQeWB8ouwmsj1PkPa9yvTIWuD2XYPZglSmcibsLIAXLwVp1PLtvYJW9GyXddwtb
PNq7CQ1KZTjt3okCE4cOSMN5SGylJ2LBmb7reu8szmB0AM8Hs8g+63NPSTPPsAYs
LB+Truiq7MRYnWt/LyI7cSgz6Vc/ITW3Nfyh+z56afYBan6sKuEzTGvLflm0NMtp
CsBsuB4yJZzHBjLdXx4VlaZXVBFJZsbcXX9iee2zyRFj6TeGryQuh/38hftyG0Og
lRcJbXrcC5+Ul6hAUE37VNic2755ay9/3NmpPuRs0JXwLOLF4BH9b+xkOfwBtDV4
TSTNO7xPfSvVdhgdB1EaR/VmVDeP1exh/pl18/t8uBQk+ZAusNMOlBP1xzsQ7yfC
5Q+hoCaI7z0kiIm5++FJ6jfhMET1m7rA0cr+mNkldYyxJIroUHwdPLpKCsjB+iFB
QTGZiE8Oo5IT1h8mk7vBwv0/Rksds9VDIgDLVVWuWA7JbZOHkbhL+/7QrlcKzvPK
S1f6bzoTiTYUOnrGavUuNh5QWwlhAgNy2SlO5z/mgvU0eqjxi2b89y/3xhxQK3M/
jXO/8IS+4umtMQdzpQxoUMs5fslRqEYKzL6zEILNG6TzD74DBoidfkr6Rn395ShQ
nmcAsmWrxHWIlZe1Cw3nmNS9wROqksCtl2oMlxcpff0JHC3lXTFJCQKvJYxiVuE0
X++hv5PdqHPVNdGyZA9R4IVznD7ld1dwmR6YqKNNHTy16hw0JI22+9w+rJBK86sK
OTo2gaRsV6s7cuvksnUhsRtoBTYSYxR1FgRMKkfNM2QY1UGAi1zRLJ/K/B+m1N9i
SYhcuKPwQ/C8ZnZ+AmP4abQ62UO/OyWrcuKB66gLgeMr3QZ4N8Nq9UHOXgtlpXdy
ynSYVc+jS8ZitjThP9S+i/chfOgnoQ/X6Wc3eRpQ9ASLIAQsSsaUPzvjlhkE2bGf
Ie1+e5plC/XShZiVWx/KdfRTFPdNY4QhJ0ElMLdKh1FUeI5eVz2CAmIu684N22Ux
jf6qLMka94UQZ2gmfMDOUESgALDKJglUCItqUwDhhPrKi0PyVYWgxSKSKZKK4k2b
+Wd7bqHFw3RfHWyg8yrq0LbGQ216cLp9rp8ktdyICi6hXSHs77pOC4s7QYTM5KlA
yzu3OWk2gvC7kbSHeiFJ9yIOjZWAF+7/UV17OvP+1MuMO4jGNMtjJa8F7g3Azxgp
kKVTjd8f9HZNKrA56OjJcvPIFzKJSxelHZmrGzLXhRUW/bq+vB1le5mQRfHbp+3g
sumYw4CLq0dZ8FSd5IaTyh3apwNHEmJcYO14Pum5q6EHTOaIyHL/2J0qvmLA6Eee
2SKPDtddWJwfPIBVz1LTeujISxVzvAsa/ec/7TT0K2x0Kp0qGWyv3hUDKOKy8QRG
Gayco5gKS/Q0/UOIsJ28/H6UykQCM7LRAksULBaLLdLz6bZf675GN86vcoDUgLSM
StvF2fqmp8sA7+EGTL9aMVk5zX6NidJR406mNnBaVmDjmYZbPYQfj5hjbaMFQFUL
LcglOFnFF3vw89dws32zd+43i8dJMtwuBuU5mJT7um1JxQ/B87PEFJN1dQ18yJd3
OlwYcbU/QKFnVTSVd+UycV6CB4hjBc20Ez4jSNmUNMsxLgw8CfqPxuclchd8sA9Z
wbQEdwoIehAhPn8uoe6K+dGV6JiVNIjBnl0Vva85x2V7D5VKpvcBaG0c8BOyAgbw
qKOjWFQknzt8lp3Y/ZR9kO/zPGQw1DaHHpQnyYCHW0AyYyj+NXyBHMznhXfzR38p
GAcQSAokmkW10NACEEgC52iQKFC506ZpGZQX0+zL6qZuWfG0qVvwVeLKVFBrzkoV
4nGw87mD/1NwPbY68Bc3CBcKB7rwlWLZWUZqD6ezzpcBWJwlJVTsIEByr/BaJ4eX
ZJOAPIxydwORaf/GEInALwZWJN2tDiGtffDCjE2qefbWwhq/csfBtYNwCS3uUnEE
qp//xRl2nKevyUkF8H7/LVAIOdD2FA7Yo/fkNpGDM6fTpdrqkPJINpK2YNYfhpSL
TUARtRafAKIV2BPQldUHyEXqbnraFr557tGGk6MdfuiQKzTqQy6Zx8u1EBbbb62t
8wUx7LbnS3ZDpDavz41bUbvH1lytdZt5ICE4prz+jHPoPkUmKRv5tjryGc4IRgEp
8PfABiHIXPxzJbqUZogeOVhwrLeBzaaObgNjdC61iairkEOjfnjvJ0X5H7uFrDzY
6NmmJ/TfdYyTFRiAuG+dNR2cMeEk/Nvf7m7lkOdjJrk+N9us07zEzRuWI0EtAqET
QhKNvt3da0/32c61fhyRssGxF9AjyGt2HWpX/9tDfvGRhDdRgB6vHSyLwswS9vyf
kKQ08VyUadOPdrFIBpXBjbwkmoR3bBoQ/XGcO6Ux2vd5W9QYoil2Dp+w8aCBI5pX
OPps7EKkJeT0H3PS20K5pF1w2LuJoLm+9DnODsFhRTP3E1aB1BbSZnzxkaQyGkvv
zat2o2ixmOK2i2smzB7Zm+FbtRQMw3E7dCGvwegz1Guo2qSLVu6gyQgXVIJme4Oh
KRfTFBNTh/Sg6c5RTJgIQfRq8ELSz3xcR2UusKut2h1TMVgyD7DfI24BqJMcEyEZ
/BZMuWRUcy2EcbYKH0eHZmmau/roKINTUR7mvNUSTarjF+TORCCKcLvzpw2uPtyH
2Z1RoNdn5cU/UZFh6uNr2eHFQ6z7udo2n4w5Mw0ETrAm1KUnBs0y4E2/G7a79yyY
LGCTPWsBguvcUMp4HUIiJxGDBvkEHG8uX0D6FBgLgUc6FiJsxICMMd8C0N8SlxB4
pQ2wWIwfr9dHSbTIXcIxcMCJ4yelefwQ7/9kgM9bh0Z/p+SFhrQ+5RE1/lB90ASA
NkDt0zR2UC1B2qBytTih0pzfAvnm0cp9gLkSGIW/5XVhiqMbcHbG34g0Qq892uwg
71DuGkwOj/R/O9ESybZtT2hMZFWpusSIZuoJzy7/kKwAD2yicB+7rRp3hiMK6xVr
2kBILA7euPwPgfEuLHlcsBdOt2EbFh2MD18449VZPf9wF0FmA0O8uHIEuQTcyi2x
JNVRGL8DVL0DAZjWdH4N489lMb5stYx3HyYOWvfiPgkBZgp11VTB3oQjmrK9xT2b
dOBgClOVfv999iMKMTqgZOV84MQmTTZJEe/VlyL+yot7YH1Wa8KtEr3MCrkto/W5
RSA77tTyZplf+ClXdf8elAf8NJx+d5KWzRv8k/9o4glX/nkswgUYul3j+Zxoe+A+
2/XPZkEqRA+bNZH3xHodBRSEXuhm24ajklqvuTq3WvwGHO+n6kuDi7eKJEfuXEvE
O/mkWB07g1qQb1oPfDS+pX2Co3JCGXywQIrldvPSv2EFIXBrJcgd3nTRn7JhCtbp
0UiyMn2j/mKzIdw3jFR8lnGfg4zSte/h426jc86Cf/9t03eHBBFSAASICYPB2w2w
yMv0wfgU9hSQYMWC9zCh+VT0iROKayiuE7EFg18O4BhF3LOc+surstDTjiWEyHlx
oLuDgeHoqhv2a/0DMgnW20ZPjB3idV+5r8IchWd0xuH6TkpjQYnkaLHDTaaYXUBj
ACG6LkzuwL8YpFzkhq8AOy52o4uLlM+gsk008kNPa5tr/YrHEj2AQCusVzw4Lpoe
OLeS5Y7biLcQXeJSkfiauCvoz/Az4V0yCa/A8qU1RXp3PiEpWQ1hr2EAaOv4SE5C
xLiKwv3kpA+gwZJh9n2/dMfnrdgyBkrSZjhfDkEm8COSp5G0BF1GcQv7/iM7iFYD
JV6tYiPdJ0GGzKtbLV0VcdURQkcoB5f1Y5w84NtAf/0gyKp24ocU4wQmpAI4mkyg
wziEanmUYKEZEplrReY+ppRpaWSUPfukX0MHdroyH/oUudSfBW77AzlWFyg8S+5N
0HU3JRb45/1CwUco8ofRG/NFh7XfwTc6quyzhFaXx3cwUn5FugICGhHMxA9NkXmJ
SSbjueKTtguJhUXC2coTvfkuUMYF+AJinKdAMPK0rzQdhDEmIyvnjIPi1+Qr+jJ5
Q+nh6Yo0659n1KacJ/b/WCjgT1AMSWOJI13jJlBC0VXrQ5E70rSZcqsCo8l44QWq
QbHs7xEwRHbF3en7C9sEYeyuYGHyEE8B0tVtGNYrcAuwutJ1cbavjBozd4+Q8/OI
mQL9VP3iLcUQgJihIRW+2Nl8DWKQfx4vxDJmpQmpegHQPCGrMksCg/wWHbZ2/P1j
XPyDRFWe63nqQRaC80S3+/KQWjY9N5/ei0nV9BzlATJ9uGEexzDrNM+AK5VUj29z
VRRF3GclONBsNhelYz0mzyiYRyIxpoVLvkyYVgGDl4SFR8Tsi/XADHGT1A9LAUsG
LXpFcba8VRdStYTlBAN5y1Z42p0abFdM2siHX6PA2lSY1NCjUcoEUNltWarwesAx
qPWtuzJTQYFWkfFv8nBXTMMAR4igR5sYJCJgiaH6w3tpLioLf67q66OYbmmYhufu
huzJWvEnUiia3NncEMYQm0Wh3P2r2dJJm1fkgsGiiWcfcU5i3lmZ/imNt5diIxEF
GdVIdKx8UO3hoBKEaJbDoONnsq8TQRSfHpezkxQuIQK7hGcS0+y4KviVmkgfnZ1i
0IVfvF1RICGOMEP/YwiXjSok9ZUZl6Tu+J6d3sqyD+I0CxwJxAiDoFDZ1PQcrHNz
cRKq7dcE9BP/IlB2p9V6dGcmbjED+hYfUup6MTgu3GWJERUZaLWwqZ7fDxZPR2jF
V0XBm9H1us2wj56vewFkoFTSvbahuIaqQk8MYljXCUBzvil8whdXovopdjClQh3l
/coylVXAooHZCkhzkHX7Gb4xdT1d7B5rZs1z/lvkLUDtrp6Wjj1lPKdR4XVTGcYe
JuVXadObslXbI3j59mEQgoswtqtmUUIIn4QpTBsBgyfqLDZp0R4oK6Asu//zbGi3
vJ+Qk0V8tPQ3EreW4EVzS/xrPypPK4vUt2E0oYMpXpu7w/09a4oTXKcVyEPtJOID
1flT3au94hYlWh15ey37umRWYONB6ZMmEiD6qDoKCkWNr3L5cpGCOAUVHE7jq5B7
Bg8mP1CXiUrIwsRZ5XZ6+jCiZ5+63QL9KGlcZs7YaZhn6egveSqBNdOfBaupNBXo
XvQG9k9mnviVqQ/LKbRLXcqpuArEmo0vQ4/4PumRcJQU4gIxtGJ52Mq5EnxAw0Ws
6bfSyb9sySYeVoYfWWpWRkueH9kEqrqo1r825KsPE70wogWTJX5rfvcSuCHMShhB
RC20MAG6ExyypmUbuT4ImogRl/MT4hRPHxmrLtall4Ug0+yRHMvNXoc4mPw0+Rak
YdLqUYY231R7RTury04yQI8xDNxNWQFTaesE3fP0anp1wp6dZS7K+domBS0DQWYs
7oNjYU+2vfiWAsy28UUmLaf6ORAyZ5UT9gS09qiSJ39YgtTHAvAOU9WyIUFlA2Vh
klP0HmTDrZHfJEeGkfjI6KSqPxI1ZbnE4i722+RwNuhdCmndX7w1Ljit1wsWujsM
TFEMTbyMnqtoTJTskQzFQl4tarIGur4WR7LIOVXiqBdfSoJilGJTkdwm/OjbgyID
KJdXu3ZJ4bRPAUBzVBpTsTKdzcvywg1YCVUaxJEqPqj7Pxbhrs9DR1oyp81YYC4v
v4jB4Bqn7prME4i3B8/RJYL9LAz//vugzC7Oa72lbRRLSFkl/x036Z0KSnViEMqu
grSjPs3KTm+to1TDNU8gMHmwyn0cKw0LFeVCCn6Uv2WgtZIgkOX9lBDzbcYAiBgz
MH8635OfU4FT5MCGZzRbenYrx+CwiOoOcUW2X2Iv1EsPmjy8QKjuod3PTcy2n6/D
qSDU01YDRl716LSSJzUBsGezmDZ2KIRvJmy6E9YnIcSDQ8IKh1dGpTmJfByQAu31
mcPxmK1BdoBtzRitczwcvXrYQsJjUMvswvB/ixmNdaqsADCrRjyj7nq7anwatLfG
aiQh/Zxpnn7XqPumT95C8LhD72T0HkWTS28BQVcyIY6+LJojZOBndqyHrk55DGlr
dW1+L8ahBMnG/sEGBBgmPNGvNf59K/GuYka0OWY8IZoCLAXdfaL2KKRC6BfZGJfU
GdAbHFFWSsoTQRwlwv6XdPj6yQc5yuZJS1f3CFW2LeueonFRKk4Rr6eIPOApJ7tO
JDhK8/wUqft7Dmx20hwjXhK6IqmKQxHHxOP24fKvL2dkKRUZvPJOkv5u8MwqXTo1
Myor4i9FDdh2C/uA5hJrlx0C59D0zzIG1C43Oa1DrJ0OLE8+Xa92031sW1U3e6WS
FOQtU+qYzS1cn3hIVzO3lxdbxuCvCyO6gqVFgOCiGg59ddrnoQq1eKvhrjoXQ8om
nLWjxdwheLOWwg89HUiZwTmIgiUNLlQVuo726ZtnB7MOAQGLruKF968O/dLen4f5
4gFGUI1QzrLM/NOktYLNx6pkfS3m45LYfb6h50t9jIjKkAk7XQJR+J44z7GL2NIW
AcRyT/RYd2a/hAzH8Jws2rI2TgLgehpmsV8Ye5F7y/ubJ8bjWGEHB6yUal+Q453R
6noYrfqTD0LcJkrL3IrdFuUpP2oo8Lc2vmldjCDSF6hI80bhLimednFxHDHBj/My
AvoMgnk5D3P5XsTJkGn582QXnBl95O7qj0xnh/+7igIFZOGDaGZi4EmIk131UwZO
iegKJmzUeJwv+kJJ/LBnxns/XBeXB2c0eRndn7Z+yl6nKVI4853GONiFWDjkZGf6
PrMF9SJDgovZuRRpWPjKxHzSAwH0n8D6+RpACurRyTzbfB57V+55deej5UJ6QYOO
bqZ7D0DhWMdrZ1rQbVU49zSdrnq+Jguqi3tV0Sca3Kw0Nird0pQw71LTtd1jIaFZ
NAyyTLpbm79sE/jO0wr3wjMbbHuFsg8pcoGR+57NXuTHrEYKFT6qQAmpgfyFkNMW
P9p3HvbIBnj/8x0RHbBFe+6hjrYt4xpCo3qDOn0Zs/bbJ62rGntXYyMtmF9S8Rke
QkLUaJncmTBhfD4yYOLbyvS6tB8WB9fws9ojmbLiabGlwFIAG0g29dQl032kFHIf
4hzeiARR6mALl0fC+71rABIUb2MWPe6Zf7P3wxp6j+FM2lC6f9XIs4f4TAIBDjtV
2JfmoF2JFc6GHj9bglv9uQmIoVMRZAATpzdZwUngIEIfQkNVGu8FMP26CmsKBToI
q8o/7PDHz/Fw48vH97A5ieKe6Ool9SG1zKs0YHWUsfWlonUUYxBgRO+wxYrdUBRW
Ocgg46ImZ4IJ35ELYvn4p31zNTi59wjrq/Z1yHpy62eKi4Poo/9CckuCiGxXjAnu
h0fDxOpx/pcy0tzMO7Ytdtk/TTefeVv/C5SXqUKZjT1ak6g5WkE+yYwbfg42fNOo
SEKzCwiUWBSVjczntOABdvJY7zXvaou2VmQrCOpk5b0yzQKh2YZ7a0c0wx6QW3+L
GpnNLgZTgZHQzb5/B5qcyPUS3OWponB723L2oNQ1MJrxF8/gnIrRpAYElhPBCKC8
JHs9r5QMZj5XAE/KWo6QrEPrUE2I6qxLr3mg39UUDa9oWLV8DCku5yNlqTb42KVl
2ZW7CEDjEbyo2U2qPg+a/fjWIcjdiiAsaZGWE2AJfPpbE81hlju1jo/ia4Od8cEb
VmVcCG3pBhLRU0ppKIN8uNei52ET1MIOThITaZpYaZbTqMYw1x4u4Ma9Focq+eZt
gI2Rg+C21WLqc4WDO74kZrbAXW9EZRjI/wvffAfnGbavfnwLc+6BclETCzmOv+n+
zys0fbRdRR9q/wPNW0mLuSaTyqnxiXOft2VCJBa5HYKl81q3hsUVYGL67bmmCRmC
B5M0l6dtHp6qGcVOagMTL8TARQYqyJiI/TNplOgomvzwW4NIZ9nyVZgGB/+eI0UF
gZJRcGbL/fT7Xg4R8maBxoI3nlR++VmjdFuosG74Mal8/YAie2L7Y4/zz8AJI4UY
RIgxIF1grU5KLePIo38uhb6M61yUMNCrbYYAcHIXlfX0SMvib922EfTLwSwMpzUq
w4cbDl+U40HtpcAInIJJdbEPQLsLiKffRUZS2VkPtEpVZ7Wz7LTV2AhRfdyE98aY
B+BNQXqisdDAjFfhIuQHlP3nYwceh64k0xNtIDWXgzwlwwSUF2lH7ALV29t8KEov
A80Q3AgaKB85f6OsvwOwwoBK++6G6WxJ560531x6U+tLBbZDbJ+gWs5FA8xrtJy4
GaIPoMkIMeP+22sp6K5rlcteoH9oCmlneQ/gYHpaua3F1SshgQr5I/HQhySY5Xq6
U/1n/NzWAjGMr8Ak7CmTYNm4Ywm9Hfr6eHeTQcTwY5iGgWIL5bwPk/x3jfI/ae8s
9ddqKcFSOlQsg1WQ3qQjNKGq/cDkDy74jcFR2ZSzknGgUoPHySl3mNOCJAcyQuV/
Ms5Y/2HgmQ5qTLAV82CZVrrF22GIa6F1a3J5BxOE9NFUeM9zby3/ikMpCi9RqI0d
p3sH184v5AZzA8Z+H7wRzxGniZPn13Rcnuudf2yJ8m2/X92Mxi5CEiilt/X2jKDo
bVU1hjDNuePdMkzoJqo9/1bW6BcbY8MimV97G3VZj0FvnVQ6SwFbyCzAw2lGetdQ
VTWZ6V06X9u8DU+LF+JWKdU20XISthBLrp1M4o3eew5Mmg5t7uqQoslefgrxp6U5
UfR9yiSl1D4SO9KZEodoomdSeZsgcEdYrnRzAtTuKo3nqRjrUnA4B0TVFq6+xtUE
eM2rgA6K0w+1xIA9e7Fr1RguU5Vrfxc3o8pf5Lqb9bv4MAQYQfTkmUd6TXWZx69a
2QH74DUjH6W+Rq106Uf8Pny2utujz4rWVLJg70jfKhwPdcrVtzG2ArhDt8wgXXPV
KE/E8X2nKf8QLWDp2PVVCVmWVv8rAfbGXrIKljZBrWXCQYfi84091pZ/i6UJcoZ5
H+SRWFv9mXYXfuZ/5VkcSdMNogxEVDo3QXt39qs9YmtFCM2QTuapKOZ8WRbPCRRm
C8FYnQJ8Kwkj6f2VObgxS8EZYMVuKb2JOrwlVpHpeNa3YiwJ+LZN+p9gSI08PN6e
b9W/nlu+2ft+NPl83EJ7hlOwd7mFrQKhMjEuKtNT5kyq+Xd1ag+aWpEkaHpRIJmi
wmPBr6/beFu2EshBSAzs8UZjGsn0iNx6yZJxu2GMD/TduXryFOnGH3IYMWC2l/2l
Wf4Ix943XDQt+I8PJlv2V8VG3bxwNqy1QlKqYXWV+hQceGZPB3/J75uDynrETKc+
qMug05wFeXp81FKgZ/0mvmLIQVU5Map0u3NY43w50unaO5rdQ3NOiOt1uFtjqPRu
YoryQGxuBOMCNNfWbuxAr5thz2Lca9sbYJlOlB/+OtHnp4C0jbVtfrWgCsPt2ODz
khsx3NCZ0TpdYnNpFNdX4Zn8nEmwXpetl4UA4Kw9k8Hdb6nokZfEHw7EaNVOEhyQ
zP4+EKoN2dVeJzHvIAHL8EllznULCgOkT2HoIoaCmAFaSV2GadQ/GEvJzYnjpl0+
STBgHJDLZXlo4IXwqwlSE1JglpzGCY2UHD3YR/avZADvm1ET1mxotPc5jRh1tTXN
N5TuU3R/fYOkFgN6hA4YzjxA5M+bR8knZgVwK0Qxi1Ol+W0v539VKAV3jkHdDFJJ
R29mrYRma57xPa4PvZpIPurRtN0xn/sLOqdJ50fiOke61iaFlo2mPmxIoU3q2IIL
jQwfm4v+u1UJ4XNBbgHQk1MZsJGqPScuE6IsuKfH8CxrNNfT4kjp8D56U4kIzcC0
sVDFT8HXtbaDSYbrpjWOrtWc/o71IZCeIkf4WeVya8ZqG9BnmjKTc1quKJ7DcoaU
C37mkFGEB4IT2+34UGNRnm2+32huUwI3Ck1C41HBHmNDHLX2pPCVaQ2o0En9Jhn4
rNd1+7SFNmfZ77393/afrb4vbXKCITVs3ddoYHWz0zlaYJVXkW1Zv5KBdvEFx7f7
ZUgJyUFQkKMnvfVAMidDYBdSNyU6qBWFO7SrCAUBAXT5l6/LJI0yzB+zce9zSPHq
eahIiq/oAI4XNBKLcvoCFcxl0gSTxhhvQE5KwSv0RaNo5EGnoJru4hDIhKm6VNMc
furzjTdP0788vA8J1QXDWU0cx90QLbxMTzrbW48wmulaKFR4OMxxz7Wh9V5A8zDH
T9B3mBlnZgVVkvkkwpY1dTpDYgzj/kymQENIK2CnNcYUF9yeIL5oyHwI1n9px0xj
q2H3x2Ge7/Ze/Jc1FAvUT5h7ZLMKOMc8HfLarvTBGan/cHjRJQukIgt850HmrVf5
SFX8t1/NRgrps7jQ+gjq04IL76y7BNcRrLifi3g4fHW2ZVZAr/4F0mcGeAJNM3yB
UDBhW9F4X4IywFrvsSBN5yvF80vrZY3/59dY9FkeW5yNpLViRqeO+0qBYYuSTS/L
fUAXsmev6kbJuGz6eKKAOzvTsw1FnEV4K0YhSPOtMQZkGcWdD7IKp0O6/bkEoQY5
5C06teDTr4IG4J58Wmv6ILp+va/rpet6sItjKVvFx7GiBeAIKIARh58FANH0Dzcy
tJ83IHdDKpir/uaLnJ425Z+9DjCSdZDa5hgtMwNmM3cCQhGwvPi69VAj+tqKDlRS
HjOj2GtoBIxsPmL77+DPmNRK2JWfU+EaYZMJRUNIBYFfnUZ8+HREhRQKDBk6iJ+u
efLVnpaOu4+8VXwIEhJqVN4mUGXk4KY/aCr6XEdv7PQh1daWHZ3whg70/yxunwcj
KXQ+6gYpZdeEWAi8snWJqp+KITp3LXJfaCcK6s+9obREkcI7l1B9cC3IydncvtfJ
azaOLsw2wP7NgvleisZpCC8jmKrG0Na5zD8stTw6ntG3Q/H306fKNKNhWIDUvN/Z
EGvgmQNdyqYgPc4rnUtD1Xk14DRvfLcq4J3o9AoEM0yt/EQRym4qv4w1ES7Ca0zS
nA3TA68ZVajY560MYr2skaDSG6MhgmKFtYNoY9LfP1PnMnVxvn/Uhwe9khAzzkZe
DqEtdMwi1JMVWE5Z6mjFmyGdXFsxA0O4t9A7xVNjYs6foDkPBVKnAw99dfSG1uWe
EIdHbmOVGjjp+tT6E3hoWTMEAKJwEMyTTBVnJNzbz5AhzM6CZ8eJiWJaGDZCWldK
jllYxWdKDLVfM6VstHXEva8CqqSglaXIJISAWzPw5gZGY/RAAgHfLAhqpi3dbWw2
dL0r1irozGKjwU/DiIzNXqFd+mpb8fjiFsPmZz1m0BLJMJeCVDzCxL/M60oCLtuB
a0M45n7TjwRsLAtymV/Fgf4fo6hfhCfsaewVIEEQ57AFY5rdLfA5tfv4fpDU/jKz
SVXO6OCtqQWGFgP4WBOusnFwS/+WLu9oSA8ZOnchFcuJCUIjsoHleYC0trMRGBXG
hT6dfihhUwVud43IhjjvuawxMBmW/88MIPKG7MslG0RotjJfonjk7gvUtJcrqBpO
7ym0dnrpcMblC4CQlPh8egDMaXrWqDtI5Z86NI1HRT0xZORpxE9TUPPPeoAVmvyM
h9xwkN3ye+Ee3DzHHgAzXRWMmwABLJN9m4ZekggHTHNvybn6jY3BX2EM501cs2Ff
rqJPeSFwHqbkulL8IG+npXVOn+jNACPq8fY1450HjfeNJ0JIsoHCO/dfLa+Sbbsj
i30SieEhVIbAobmp2Tiu9w4sVsIReULS+BL2QssfIrVpBEJccWYU61IEFFp4Y0Fj
ZhN2tV/8+RGJj+IhvSrRa/sx6U5KgmCs0KG4bNuL4YoYdkVltL9f4Q+btJP3GIcg
LmYjZHI9LbVstzbuzIjTY6mu0TTyKZHphKGsSYO6ziaVRX1EbBD4I78IY6BHLWie
OVrggYfzV1Vy2Hn/yP/KPYNlEJq9zSb4gcI2Xo9MSphaS8+Eua67X/vWSphGVUUB
qv1K7yaqDaaAkFinQ2IGAmdOeyWDoivS/KTo0OCT3l1ea2SlzIcJZe+Su8LqGNhj
dSKvNBz+XUeBalOk9F675sZnxd3z/CUQ16HrYdsyXnwUnmm7hZPHTJ0zIg3eOC3T
f0sNsXp6wrG7EVxuCmZ2EKrcSkmpicOhoJOy1/vIaDulWgW57sH+HENPsuxNSAOY
/mLSLLz0RC/5kuDMW43Im/k3hMGklhXHoDPiIHdZnQc8fjxR1+ShQ7iStuMd8alI
LP40crXHo5Lu0IsoXEFUZbB4iQB29/ZgBWW1rG7KC4/QyYJDajQE6amIzxu83e99
0cET3MNdsR+Hfpfz34/dd31tpNbtSyXhB6hMRFg855olSG41ruJFjJxMbS75eRbE
13ZzCi7+4DhzEmS8Hud5y1T3h2MdugSf1+cL5d+m2uramqbyHzCmXmHcU6JW/FiM
xqvilhpP5daCgOqrcrcp576xx9Q0AaoO+TalZb5Z7ONAZBxih4h9HpBr9nzQPKE7
jRUV4zC/pK2jbW51tf+8RIU+Vf0GEP7Q5AYMlYTXEzc7/NPn3q84eEpjFJHv7yr6
pxFUIHSfQ+72Ax8QlioF3zG5w0izfs6IUkUhcP7xo1SbDg9mCVsbuEwJorKenddg
BlJdMYhYRdV4hVj497LLTdCYHhESltRThXpmU59yN2mcrI+9lvxpTN+TElJaUFVt
5Sb1S406+SCiujT26alYxzzA7rV8xJBqxQH0BqXwsdkm8HZs0Tx0wVPk8y2SNQlO
3i1e2qdvHL9s1ynFfEmvDoyGKsg4O3eKMZG8oBepevCPZkLRXghFToRVwTXgQDYb
ThW2Xsb0RnI6ec+kHo9hXiWaYb4ALKe5nhjAMBdri34HdRlgXTd28CnLoj4V9h1Q
KVJfB2bQFz1IC5m4Bha5UFedzJYJDzCIn8Kg+6Ltjedc4Bfrc6q8aweV1xpebRqJ
UULAkSNxAV5ouiPdyU1KKqWUOKaL41YIhlqReasy8iomxFgmyt6nIXnvK5WvSxTx
r4cqRDc7gaqaFcKSuVV4lxuO7HMukIKFeONAcgkiUffdLkKTcmjwzOJzsXY12kxz
6kpF4O1c8PUs+F8cD8nSvGzU+YPISHVjCN8ecbnrFJn2pGBWjYJi0WRnGI4rZQiF
aZ2v9SvQDOO5gwfyjbpCt17NGDVjTrt8SE6BZIkVjNkLANndPFL77Du+Ip/BBow2
+Pb2nBo45ziZClASBKf0JrVgfdvrMi6rBBz6IZ/S0VL7CQfq9lD4v7UjxQSPJ3RR
aRqSWSOF4SyXbSNT/clwU4omY5W9XT4pudKw9CHUXBYdrU5++gmlm9MlCRcZUnvk
07KlWCtX6CLqOVtZERphLINMjRUYdWNKiCJ+jb/z6BWDBZ270eTy5a3olDWJNljm
E6p9Zic39vI6xUbUZ8IyZlr+omdOofPgac1GDVcikuRkl/tiPCEz3VjVdhvyWQq2
ucGD6lNSUa7nZgT8sis606v67NaSRETOdhcv0OseMxshOZQYJWLr/N9Ary1ol1qC
gjkg3UNxq2ubulpfu59Vwci1rKNOT+4jCexEGNJcb+riDqHojjZYQbeQ8TKpAf7Y
6xXxsDT2cOpa1dcaaeUyv3vLqSlRqgS7f7PCFMcN8w4jfDcvbZHUh+j9Ljqx3L4C
lge//YKk89Bpigxq547hJllTqBOPskI2MWNqqDEX+HQkR5h6JIA4l1WuCWCwwa9/
S8dPr4UsrVf21DTSmSoRk3WJDW7sx3LS3X0cI95s5PtEGZNatnHlHiT50/hLtPV4
chfwOqJxwEgXUeYww/5uG+TbYO8I+KKApua+pjq7TVuOvzgAcARsVPRVGUeqWFOY
ECpOorKXsZ7txZYpVDKfslBSpwA1qo8+F5AzKzpwKaobzN2+oPhJBDUzOSf23ui6
HmhN9XIaw9bmZyj0lC1SH1GV9Hw4+UOEorJRaa6h6Z9t8K03nweYS/FSXEwOJR9I
U0GNy3iHb+EXTnmtHmK+HtpnVE2XDheoFS4h/zVjftVnYH0NxqafewnrleTrMvy5
lipsEGLEMfOBThGfs70fSkliALyX3wvtZuXwbKzFyPNfVrdhgAL1ZvnMXuOSr1yL
pSTyAHTLG9ECpCYLk+/QABv43fBCpNmL105tcM/7Il50fTzvko2hCZNK3Qxi6k6c
LvsQRrSgxIOJTFNouvm/k5p01sNoCriwWsXD5fTrzz7Tzh2k+dFla7CnWmJKaPLK
9inoLQZIiYC06DUn6mAlGolBCPB9GTRnE61Q04M7iVbOZJO8f9CGqH7G75ALHIM8
VOx13IM+fH4Y3B7Xombh4fNXzppI4FycsSK7Z2RCQs5MCmcElQXmZ4c4nTMNGdzB
/SEHIUC6yp8E2+m8tCoS5ubPBbnbwP8qIBdEcZhSs6M0ZZ/atkAdwLd4xCWVtIm/
wxMFQigmLG8Y84GG7R3cvZy5VObogt6X+OWX6TeGBToSOjob3lhMzEYGQml/dvHu
/6I/RXD8iU5qEdSXBwfw33QeqmMGNI8dDhg7srUkS/i5RcKjPDaH0RDWqniwrZ9E
USa/3pcOvfJpalp/+tNsgmkHlr/+PwMPHVj+PEaKQ0UARqiy6yodwQtt0IoZLAmX
liU5gC2NHtr9cTEgZS/3ConiDXS72IpO7QgtHuoZYMl266rCtPvwWMQRBvVhqKrJ
IhEjurEw3WaPGR+6ftnK+bdlNsbGVee6J5rwrl9W7W0d/J/MP0dA7NdV5uQwKAlU
Y09qxXj8tG+3rHkVj/ALZaOFEuMae4ZcQ064jCWc24tXl3uQyP6nqsUUpf7qUq3D
PZP1tAK5otWREnJa9m9HDlaNyFtBAxGTChJMZFvHQspyvxgrWYS6SwHThr3DMbSQ
1WJa+Bf2WTlgfYhb32iJxvKBKhGA19T5NxILHNphPz2rH63rTi+1PXpokf2u+kuV
W2ze40BadXKzS87/cLriWO2r1BWwvuR+56EEHjdQSV3bVubbqTiPqMOuWEzvEkq6
i7LaGrK+NONK6d1VyuhpcmWUphkDZYW31RyHEseLeLI40005gaQU8U5cMkz2hLE4
3QQ9sVz9qW/bCFPBQKw5q/riPXzwTDz35As6qltYA5kJ1GyAYOlKKNUBZXv2ioVV
b/A3INeTcZ9nMGqVtQOhLWDy1yCqMjzEifMg2KxlFxHPICQKc3fNot/1yvnMmwTs
ukyI6F+42o5neour+cwtmluNmianyj4d1tMiSCoVO5hKKEZZra+eTPM0cv07Z4VO
TjAQfgmJgz2/k86M5ZDLlOMPqLnvzIR5qVkYFvbZQ22W1+K8JwTujUqz/vtzcWty
xe+vCrGWlY8zgN2TU/weRS5C2/QyIkF+6ZKXf3w8FV1hVk4sB/PVPNrYZwertTZQ
wzrUuEbE/Yg9aW2xsangVFKbf/r5jeuv5fAPazjcV16aVgY1Y/uF6D2MZYrZPryO
6E4+N7x2KgqJENkgU8sr7K1ZY/Xp5hwQyR9Uyo+8xH6bOUxpANjz1rWXxc6dThA7
hQXx+cxr8l6PZBlKSSDvtFNDIuci/Q1qQXHgG7OrLW0zV2OB6oL2uEPkCvvtjG4o
MAcAPtTm/i2bkSxcZJvZXkKVJhzeAbYG/Hyzae851XrFrk8y6npPgm9WSpngfY0f
ewEUlpKfDVUEAAo239ia9C3Twr21KLk3+rnPq4AMe5iQe43TdACpi04GCCRH5xnS
Cc1xL8y9P5ObzcYnL2gS/6J3OKGZbAwI7r3H4QvNOmIhl6Q6a7/myzmViSu260Yn
CkRrY0vNqyUcEe6NXLHbU/+FwgVEuqoffUIpbo2a+8ryh45a96SdFoSR+No79zL/
xa1HRR4vMHoRQL6NLL6X+RWapP9V6yJ4NwMaKMk+MZnf3JIWviQg2ieGNoNVY7eh
CJWnzoO3RNBaxtHS3mxBV867AVhO433DxAvxG9Oj4Fk/2t3w1A3aAJxxONOMLNKY
ccrH4uWIRMr3eO2v9U1LBVIiSLRjjD88ikX48BfjMBlg8/N4MzWjcb3jIcShKZAz
Rv/X2+392EdW8X3eurmLM9dqwgLRWRmDkwCsjZNndshoh6G1bmkOeRv1sg4ZSBtl
jzPg6uP5ZPyddcT90+HP/09MA9JoNfisWtycB5B+u2E0cAdrqkZea7XzjA7LytkE
/WNq+XOF1yUyybOBRrnbVDqOpMXHp210yE3FNasaswx1O3VmKy8slDWOkeY5pufJ
uCGCthFXytt7B5+LMg0SfowK21XTXI6rnPkMwAGLAA7iBe4FczjSrQXZ66q08N/z
Nd58AF8KQ+Dur3ZiW0na3dwRuJ7HdMI36OcFKxJVvgBoHaeXIwqzJ6AFTTpmVlUm
lh8xk1nJx9esFH4a2p6y5NUiNft5hdUwdjXgy+L1gOBK7kf6rMTdx5cAD/DEwEfP
t45B82FHYMPrKT2v2EInzgo5Fwiid4cfadl2uqrE8svUQ6eMzYcUz2d39rOWSSDU
U6uul2ekWsJUBy7INyTwNYqPZa+dSwGhxrqdNY1igGxB/apuVMj5T18blwjRK096
T/p9NO/fdJsl7wY4a1DvQMVe4gwn+f2UhSvM9fFv5fiJ90ONlEvhUid65u/ZrLpA
yXuqC3PIXcCaI4JDcrQiLEEQmbyfTp7b8Lb/Mn/EnCe19veKJiyI9Xc8qbZSiWvq
evW8VbEehBkqd7fO5P5cT71EgCE2hWNDs0fOkkbIDSOWneP3Y2ZawZVOVeLtMGxU
hYwkC2gNfg4KrtgnrLCLZaMiFF6KbKpiTc/0Mud7xajzqeGi/0pARUInqWG1pIOc
8wlBSzX+hxMdx3eGhl5+pbBCXXeH9GTEjYNbsRO0WXg63nVxAQEkrwhvU+kX/fGX
S1maLGXXQAO1QkmqQqIP6vNL3DMNGQLPYDVx7YuZ8Tih0pYiFb/UN1LxulK3ABr4
aXbs5rPU12TvjW1fSGcsG3Ez0Zvl3Tky4X2NmULTyT7pFW5xLrbxiyuVMuDfuEOZ
meWJ826xFoB1HSl+zye+RDMs3FPgIEmKyTo9XDM57rMMYFg358AzeE9k7hRili/X
NVBS+Q83F2JA1nQhh+OGY/qPITjGmqYEv5S1yEWKPhMkuRe57qA+KYiTTZ717TUc
Y15m3I1jJUn16Xxir3+dIIbNz3gLSW4lvganN7+GlKA6XOF9LZrDu0Mh1g7srYTZ
z4BLJVNZDrXyDdO+dtfOjCSECNVixnQxzEgC4yBIr37rHq6W4j7MM77if+YQFpJ4
6jSK+/DbOIYkDDwA75bErVmEH/dlZEfpmto9zw1OFnWyImbo/PSJOTpnvLbWSXRV
iGaeNH8GTlKnBo8ScrrI/pFWI6XQQc/yyZyB/4bpcKl2ReBSMvQNc+Es899yyoU3
yc2U0AVXWIutniazFqcASNAnX1hf5WqrhF8bZgTLLSBmBciNJruX5QJbLytGVu0h
ruO5CA+3EB7OS4AGJe4xYNDe1Rm27qubLtb3ClA6h9KdKPAKwt6iDGJiL3GSqTen
yuIrHr3sdu6Wd0BYOSF1XJT360P6MLl5azh0XOsLn0FAcI7nZTBK2I9kJ0Xl6iBR
FuZuuPC5u4rq7gbADm41FJqqqr9VYJy4JelhqXfJEhUZBkWcwAKqyZg+6N6IYtuy
W1ERSETUOGctmQt+NR/C1Xz1l2/XOmDklS8QbqLnvCP2r8eXEbsMbF5dumvnZ1IG
bjC78i1dr1T2bTH19Nz65E6FprhhNZIWp43wolDNgix93zYHziKVcxYPbeEsiz31
DRzgT30DqdYX0FlcvdyYi5bI9XGSUKeMKa7vkJydl7/fijVm3GxAWV9PqL8NoJ5c
R2f6o34b6PAe7nDCLfZjQNeP6p05bY0dtDcHgS4Iy8B+lfDIX1h9jlB0xQIGImSI
MXxT54lNhcDmP1AFlJd95ePdkhkaYdn0SPMwndOWd3VaaU8swWxxbP9pUKRdjGwq
wI90yTth2h65SvvIY5F/0M1+5tktLDiMpTwS1ZxEgzXLFyiBiK/K6BKpobVlUmUR
C2ui4ZbylVVaiz903RS4FMOLUFDT2mGJpd3GUmsdVsefwwsgpNsd+LrbEeOZkJIk
SYsvlF7TEnOseRJdruP21nMQG3rgcA5ufAns3p2x2kjwYUJLR825RSMXs6KupBrt
q6HJLGx5nCP1k+QlmtIC/C2dNrDkns0mzOO037kJLGg1s9lz4GOp25OAw5bSaw67
hfyiRwHlCYoW+MNV7BtQSqcdQz6EzdFXc6YjXGZzfGANgD+PovYVVtl4a0bWu8Ap
fT89xSQRpacnR/ya3wsPOlyZ9ev/+rvMsqovv95DeUA6VJKVHkufOZCP63ROHPrL
SGNrC9ePtoLPKtTF+XS0BYbGWnvnULCKAf3YAGRjdH+36a2AuVSOAookN6wdSqkc
P/4m0RXpbqwNCwiMSd8UCy9g/EqvTjAp9lX+0pWb1fsJJ7PP5zhFercZpyxRqKFI
sndSG0rEcYp69nx67DmDu8QoDglgiQQ+sXxBRoKcy1VDjsW0H3F5EdhDmRgwyTeL
NPaHcm/4YXYsPcEjeEuhe4pHUBQM+uStOylwg5+fOiH7Et+uJjP86WFJFUqmvX7p
DdVwz1r3D1gUPoaInBUglcMdWw6cPYIUB16ndfmlAfbUTGFWahOj92OJRBYavVub
o3g3cSL+24gWrZWybBTYjLRU8WB/E7MjmlD7naE8H4QIiMmCLIiT/za3oHt0ugFm
G4JwUQz3OLVcVd3MtKL/A2IW3aUxBtbEIT6CyMnxV8pRP1HqkJcE+V/wkRH62QlQ
xEJR5ETqaQw9P3qAA0NarmwsiD1kdYP/d5GivLdnOLbSny0nL21qhvBITuCwdT/p
nXyWL9MFMfQdB6CmFKaZL4aYwhY/hQt6a2QYR5Toosex8Tj3UXs6XRXQ6xec5zL8
IQHaMNmqpdFl/Oh1+QhWtw0Gvy6usN2xsy0cTqx52/BAzfbJMSA5pt4nZwromYmP
9WlXLUZEyLCMJhtAQTwZijc6m5MAMUpWc+XsVmUhZjvW7qsqEIpvw2LcM/4Mit15
CDrJ9JO/vD6E/r39OHjOcBdOKlGNZGN5NojJI8tbgfjZ4UhSZ8iZRMiUzdVAbc36
pdrO69q4R4zo9sKio6NOatzqYDq6OM5Sgmrt0+EgifwwB0j7C6Pr7l9hRdWEHKLL
37+/AfTru5tbALGPBsdbToOXoVBmXRbAu7Om3GVpyxWXTvy16BEn9EwRZ8fymiR2
d8DJyv3f9UMHg0sCVz/raELuhEeWC7P2Lmtua9sMR+bNDMW9s77p9yM4Ao8eCYtl
ssJP8RmGyG5fJ0gB9T5953KmBOH/Dgc/ZIl9zs6gF4akJBE6A9IpGOpfLukNT7J8
JfWsbuPIoCQgAyHSzwjNRQ49yCmBgfLp5n3nHpVRDZMOTtmYb8mgx+xZWMcz6Ia1
kW5qW9yKDQis68Sb8t+yKqnBD7z5t1bWLVxdkDhzv0YY69LnLSJgeY7pQYavSGdD
5n9Ok5jdLjnlTRT/Kk2oPCtSi8YM3VJXnoOOB33PDgs8KGi6riSIgmGZarf1ZSAc
Mrr5LCZXYfFevV0WNyg/uB47JSHRWw8OAhljbquvm6NSBbSflLyJvF+xeTq8UIbW
dmhqe7a2FlSpFZqXZ5gEEY2cq6hpcmVTrhZzUv4D7cXUTiJ62iHNWgyhXXPBwGOJ
YCvdwYCEDtFINBvB8xGIYbWW5cLFSpxwP0qvNH8Ja3w1jHuXuetbKhJjXWMZ7rbS
6o3ZeZcWkKe7iPJcflD6kE8hPb5KForlvgCyU4oWev8pr2l1DhjWSjJPZwungiFc
Dv3ZuTFXdlYmDX+zUV+SpgRa8F9Db5UQogiY/0Q2GwPysHmWkQJYI2XANupGhlVt
KvUT0pa4ottGHvLgKkFaPqHk5QfK77oYhvxwaVWbeBjqMF4wzeC6SfMkT6HbODzd
j0wWV1LnAKQuZOUtiaOcgPylXACsPM4Udj4HfXm4tzyA8OalkoTFmfqctVHoFO0S
nqAFh5TrGmZu701bpukaZ9W1ZUoX5/e9D1SxiXg1+IS5GmKf3BnfiDlrwoth7Dux
zezF+eZ4vOrJ7MHREciuUuOSZIhB7pSfZ+zyjouXgvLw+4aB/iJUqKlDHVqSWVsR
gaZKrdcjkUb5eoonRj1eQ0aty/ZDeSsACZd8H8X+gCqJYFZIESdkZMd9msj7fksp
gmGVKkhWHG9kt8OLkgs4BsikRnPKIfdsu7S6dVbnvF+2mQkgA3WVmGN5yvUqHgNd
Wg9aalDRobj2t3qw9gh49RfcHwR9Rv8AHzsgswToEjvwf8CmyQb1AEF9xPnKya3Q
vQRWKa8E4BSmF4Iq5bbrnkDI5bcee+76X3PmDavodrUKshof7S0/1e9nCGztnrQD
tn9Q2GOA/87p1RZZI8ccqsFVXNDHmjiFb4q2NeDN3FpYN9PxGT2nhX57TKDUotqI
97vFYpiJIDw75tPtKmFJ4x6dyPVf5/YAX9UlKeUEpBzHcJWGCRWMGnl7r2DoX8DJ
pxajoP80pUDok/v70MZsW365jMDfMH+P2yz4tL/6IGUC4HQoEHBJveEvuf++jCzY
N5BMO8LHbG5KaboqAyJ0A8gO2pqh9cF9NN3qOTQYZ69h6RnDbci0G/eCNHttKaln
grcQOXZWswLPoN6qiined6oqXW8hJR97hdQ7zoPWQev1CegLdbIH1KiHbzdFb6jf
xBN9tWHv6qSj56DADgyP+qC7skIlQdwiAyy5Z7HYnaPzVxY2v/pSudAhoSWxI3ao
ggFY2qhHlZW6RYLc03cDPxa9OHd6eQBZWW7/uUa+XxO8h1Hcypy7i21td+t6LCwi
oj5et4Qc2vRHjnJ7RjZIGRhm981+HOE1QVdh1ebakpHWh4Tzp39qHAAfcmTn7pMD
5C4+NDhTkp1qZvZkhfYaqPOrcL/dLe1AjM3UgAI4jgZbTf3hLau+wNDiwZlBDuCe
o+wR92NuuMZouO9uxS/9kv+w7CNSyHKLpYjmsRyolAlg5lOdN0+xvrCN5ORG/6gp
wJbEf1w+1a+5WPHMOeBtZ+72RjYam+ZjsoMj+cQNUZjERjWcWj/z3jASh7JXDp8j
RvGIOVJJ3waf73vG7L1Yiwtnu070kEcfM0y1AuXt70tS2kwXjqyUCpsNDM1/doMJ
zs7gM8SkHrErkOOxev4BkjrmbvNYr16eMW2o03KBh4odevR9AzSzPGXWXQldJZD4
V3fH9Mvo4egzIpmb+VnuGkos7us1cXCov+NprwDbQxqP0o6aqtx2gHriWaoogo34
+IKKWoezUKY7kyF1tMZli2BQl/0DKTbwMhmwlKshtXuSeJgrVV2c+E0Qoxr4vNEG
PXhu7FLK26iq5849xvtZaAUdXCZa5uuNK3tEPyWJ2nj1NrecQat+fZj9WY/Ma+O2
vS/ioCSvzIeEUEdGFx4FkGkdzD5SoJRZEtp7ltu7T8C4kg8y4liAOJN9Kj3RYdGy
BrBToOA7Fsu6gsxQSOGFrTGS0Tu36IGA/YUZlmKiuUHvnDretCfEMpgP520VKMQt
mLKh+/tBeqylYm0JgKxqfTVzHo4Y53+ZV+Z8iRX3ue2LEh/pXg1ejkIeT556j+Gu
ieNV/t5jf3p2KsmoNb+EHH4SheLcOMAsI2U23eFSvgKlwfctelPM8hPo5RvWqsaZ
DsQwY9Esv23nn3DXAGfnoEDRePSFf7O31NsmX3kiP6EMhxf/911XjsvkUH1iJaOn
5or3XlJj6cHajvd1faRPG0p8/UJaVj5hS5t0YoxmmLlqTr38xkLwwRvNQir0kCDA
n4pz7KB1/BC4EpUpsLUXqEomiZkxmhpw/uF4467//iwSrnhOqj0w+lySnoeI6ojl
O0w8oxizKCwj4zdFWpimVCcfef00wfBuNeZv2xz1gjCUAES3JA/TfEzX6E43MnA/
w5LlK4UXvDpnFr6v1hhIWGXxCIJVSsjMsoJXsVaN2YhV2zW/PGlZlCVAMQG8A3z9
BaKB7maQ/QXOlmxMr+aAVALgU3oPyReUV5yidbfr2iv0RNNao6Mmqtn7cdDn2Gny
JzEfAzvwAooavOWH0wIcv7Zqfimdfvx+DwQOK5yExdav53o5YqVxoGUkxRzlimSm
Ka4LgdUyEAxg4GiE6wA2ivk3Mq79vTHCpnc7MpbFR0/mIqFc8UnVPW+2Xa8QmbkB
3Q3tQMubGFagpf+u2zZkPhatn/my8pr853GumJuQAIwWlxDmb3A9NMEot1HLv56L
5xkyqh3OeCTpy/fA0T78Tip6SqN+cO/ns82cYPo9H054qgtjWEoDAW7/02EMAd+o
4VKR3zi0tX77NzmsMrq7/DwaVTqzdvqURwbWFv17HKDt1BTBrcOy9okhNHNgPLZO
4QcXK3bkAxYqNcfA6iRpumI9qDkz1qveR3PFmWq/zUtV2QpRHjFV26e6YevOUnQ9
lBZUlKtA5SjzQrBJwtu9r+uFgfMlv5qFI8fVFGYIrTv0KcOdvOwuX+6wt85DWJcb
ykPuvFbrHQ0Tap0O+aMpwX//Vy5xBjtKUAArr3eKe1AaojGyA7nrXA0rxnShaxJ/
w97B8iNWG85s8CRBxtr/0OFG1/4SI+FeVgo9D1DSqSkhPksGtk29lRz9834pWLsx
yIia2gKpWMar5TNG/dXZh2XMa5O2zK58vC7kC1Ugb8OW8Bc42jYszh//rK+wctF+
obzSuozqSWHnk/9PvqaSm+T+7hQjT+jWsFLWZiYv8377gFz2fJsAtZkOUn652hG4
Z8Bo0n1S9V1UTmFcUzu1HtZyA9a0qVhxWsNzTycSr4f6p2GyrxjD7u2La9SlgZYn
EIgGkIE+0J+iuXdV8hm90N3jcKduW6x39Gx1qzg9TFX+MtiKFcFvc9k0qUYHVhqk
2rzPKI+MGaMoDoEVcD3ApDYxzK3i03ZID+AuWwN5e7S+BTSffWY1nUd1asoU6LZ+
gfojc8eKnPZ3aC4QYVnxPuZYB9EnUvMXb4UIpD2o5bTrDy+m/Oa6Qtk2emqQTqLc
1Saj8lpnVI698JMSuXdg797mM5n3T1DWUfJUJnLixcf+OjuT9lQ46YqEIVaTka0b
650FPtvxb1PGIrJLo7R/m9WinFBs7DpwzLD0Yy3Wa9QBaTw7RjUjpDBGBQ6NuHHs
yI4K2BojBjtu3wpeLpXZCkzMuG/GEcuyyad1dM+fhJ8uQYWMFY9PudhjG4ET1d5j
qHPl1uyDuwIo3sj0CSfqiW5vuhI+BBvV+0RHHHNlpnISbi+Ru8Tpc5TTdvTP7VqC
Zt2M85KWw+XrhGNic4f4bnrlBMcyYLO/ec0vh4n+cNR3dyiC7yPkdXrRV3pUzEBL
27nYZi41lliPHwS4n+Ra7bnEeRl1MAg/kBo2j5MsY7Nsia8Ij9hnjNpll5FO8Qkx
vS4JNcROgCPAgrxyCDIK2JCahbdYasvcryjr7XaFbMMn2/fqZzauAQz35Is3wxyF
Kc0a0QCHfIiYy3sS3m4DwEPQLdmKAWmcqFlgqLAq6vNa68Y5XVh+7c/QkVvQUV24
kmjHNgqznKQTuP8YN1pujlbVbGD2j5hwQtgGOBORK/cK/6rN88bGH0biPSNAZHSA
8CU3rHMuVOh9WvT8kj2UmBsC7t0KA6cFm1/V93WMrGGavpk5O0AlnWrP5IzGr4FR
qWAC+F+6bNCE6MUKNu8M03S1JCBi9S0hDfiWS99JnIde+oohhWB10sp+aEPbdo1q
4EME9z2agHoeZ0X6K34qDiOlgNAgnoDXUD768Dtlgi7uA+dKBFXYcuWNmdWgnAHB
UqIxom54kVelvbmRIj3jxeEf1rOE6k+7tLKJO91eBaFHu3XS8RFiRzGF5yAHad2E
yORBttTQGQ2vyhFmz8hnm0LEwCQApBuHfqW9I83rkY33UafyArxeZgZvgA8v5h7l
d1jaQC5acChIHCVKvE19rABI/efOBPjQdywPkeDUK2BQm2tcfeFovFRkYxorIBai
TIgPZjMX96IuVnONNCjUHoWs+dbmFaMAd1KWsMfeETBjXhiy0Ad4u4NllAlyKwn0
SPcbnZvs1SJUUG2Osr33L7PpiN0WiOcljcesU+KgmShPelz5dRWplw7m7xdNr5tt
ZpBnkGasrtD3krUwChRrcEh2APh9UM05JJ1kCYYe7+IP+4r4Ii3hs3HAlAETsqHd
z+Km8i0HUkgaOMKhaoKkryF40tZObFXUTf2bzaNR073yYGTi2KKtX7n13mIC98Ui
YR5cQwU3jqHaYra1Vy1wWEv7E3+ibJ7HiDiSU/Uijv1AUFYMTFKh17KHrQ1aUOd9
U5JjSt30VRpON/dTscPkUmNkJ366Rb9EbWcl7C3CtnWomtdniP55lwJk2d8aEHXH
9FBJS6s3eWdEmPeqCqkqVOAbzOb2mPaZLHhEBC8u8On36wWQtRlddbCiv/I7Z7JV
xoWzpYiVfogpe77T4e6JJylPK+y/b6V0zS4JdiuGdrIaycNYTkg//ZrMUKIRHD03
xIj7S6vGdEhexf/yEa+mVRlgp8ZZ/gchn3tvc2taIpwDgGxMpYw4kXOrn6NaiaP7
RMFjyUQuSN/vam2rF7gM8QEpXJNyavoESrESlMtvL8yQnjcU6E2bZlQimUwe2BQ9
CWvFcMIAGhmRpz4snZYMPRmok+AaoWkG9NAi96iM2GMtsinYUrmTseCiLvtnak8c
TKfbKfDbMBtnl4bCNvUuupqF1qE3K6sqT3+LZTk8aqzxiAZ73qyG1cD0LqBOEqwz
6YZaFsxNcOTTglNGDPu9/WUfPAAbjPpvqpjumXIgJ/io1cj0YeFwxFr2pbKKe6Xb
wrIgj+mJkaSGWZqbDDuks5ZD19+l5NBZFdC0H6CCRXOeq5O4ytU+4skkeAevCGy7
aanqdu0kQn4s635o0sYy6POxqu6Jb0wo8qAun7yHilIz6SyY9BVRpoOp+DiDTbVT
kB1C53ey7neGt664p8ixGQ3hNpleJDSLB8oxtwvEm+jXrfSzku4NvmePcXNHuM54
MaLDoWwEyLDEsp/84iU4IdREiryWdcK5M/QEDVYwItStxuvdQrAd2g6w7Us8McAV
cA4dqxQ3AGm+580eNZ/D1N+xIEiIWPXUbCrRm7UniXinnbR6whFR8UYCRuvuQNsT
YyRkSFFObgnnRP4L90Zt0iv4JiSp2DbavOjrArRFvQ1yhj96vz4SG+2favVFX4Ix
Qhs6wdB1nMp9hG08Gf1TKdeVZTSNi2ybXMOlNnXuLTMewu/qiMBoRzlXlQet3v9q
G+t5RtTyWPM7bEcS/ahfdOyKKV6cQniVmahZo8wqXkqFgY4zimuRY1mhFLLO6ono
cMmtSVQslwXNhqjjlSxDQluZamz9kjGInMdA3oJfLQwbhNdP5SQATtEmJ7Ytto2K
IUQ9lfFXRz3boG/C0XurQc8qt0Aq7suMeCGfFT79gHw+yN05kEaV9JP/KZRgx1Zz
k3XHRO2JNyEdRLhFwpej1wJMDYhLUGfOSrvHa3+CEFJtrcx45dM3ABvzOhtMxuFO
/VpSAl9nQ8S4pXDfjyZLJ+jb1eObIU1oWirC4qbNjOUbnzvaVsAp1DKF+XHIPSOr
JRXKdOMULsweXqO2xaiLBk4i99wTn+i1fyYN+Q0J6T3nz/Fak8HldFAdtdz3fTtI
2Pta9POcyQt7qi1w4Xy26/bfsw1wJKNrmlQtfvxKCDYex6+5b4ebwQvkV0uDadAt
t0fd4Y10f6V+DUCR03j/baGtr+ggyy4obhGJCS25vsVxfUkaF0/ZoZMRxzMMJQnc
DdYFja49cf/ZKFHzkHMdW9iKeEAdEu317j1xHGNKI7NJ4HQ3mP+LE43jk3fKtxYE
Gi2r6DNFav5ZyIAMPQ3pCH1OhKl2XkgZ8zTeO6EnUjlFiKDpgBxDCGHOPwYRL0T/
GASx0TT+G0qM+sZMiy96YOUneiSZcE4H5GIlZwayiea5SweI2K8Adkj0TNTJUM9i
tBX30lr1BNCH9nYx9TL/yAooTN9SUHnsGqXeichzD+QVYFtRCfB6Cqd5ipyzm+iV
yDVRCorRRiK8+Quybkqagou5Z9/EGPw/KiYlCC+IDK+nx8krnYQYuQ8S+ylI5D3B
cfdfBJ4pvQh+KnoMYk1QHfk2Lp86UCVZMB2mhnU6TdvHJISv+m6+qykokoXPibpD
QS4P5Rcaca/hEXVI9fka6TJUvBGpHQCgj/xbviTESchJ9ktuBUr5HMuodMF9m244
eJbVnozzTMIgATjf8rnFE+hoHx8oEUvEzFtH2p3KTVYjPSAfAYBeHtQcjQySL6ld
z29L81LjD+W4XUobLv1Sv5Qiwq+6zRH4wmTDZkvfmDGjh/GFnODQHNxhAt+wkIDu
8Zm0W+WqwgCYWpFHJoimT2tjsBLdu2UUUy8QY/Trx6fRX7awGswwK7LDShVFKcjq
of9lloOdvkbnK9xXU5pUrg5Qv1Pp3O4MNrHOO9NxY5hVzGrd3lEI2sAU9bsfD36u
XLU6wjhJQuQgUJ1Hn1WcOb2o2fGcRsd6oT3qsKWOEMLG1KevAsyLnBEhg2GKpKmk
9uxwlYcC8f5j9+a9o9dsmnJ/Gns7v2Qn3I4PLy1FkeLStU4esatzhHlReDVjXHop
iA2OahY+Z+dkDFLgkxiOl54vtldWzUuznKdYEXcrcop9ZGDKMEqbWms/2lMufw35
fpIIw5RqfkJ0eRGdOwObqEZbiQcmVkuvoE091sVmO1WE2GrLKremVnrcIR/AKaoX
I7GX4psOFf0zT0uKvEXEaeDaF1LAPw/+HmMPxuPoBOlXc39qUJ/rF+ZG9fVPMXvd
SSXZ+YqDCv1nS44z3bNaQVv+mFfoO3dr/Ha08WVDorPqS41oQXUUFEvtSOHTdolz
bKwSxA8NjyhKuEhr7Y3j7LDa7fia5YQ9LqQlHHCKAsMIaqy8NdV/QCFwR7DvShEx
4wugSDHj7XtSRjk9b0YaqAqSSx/xtv7nW1xFGrqIyFa2zaUKlseWRMqkTW4NxwXr
FJ24yJgpeQgc77T5CfCYz1tviCSxtCqojf18VZgP9PbWyKVOITceadaqMhrL3dTg
v4VrPzBqvCNwpUTKQBmV1p7YT/BFtkWwsNtwpkBnhTuu3PzVMd2EG6Ug7CfYZ3+R
N45SDuV1f2oVbLswRaUMKiPPgSU5c4VRlITRRja8oFTDzGrPSCiNgFGDZmaq2/EW
PSIWIKn+2ADqhfOW0Shwr7wje9V6g31YS1JHFd4Kc10nNkH9HACglxQP+s1ZTPpX
jHTo/UgCE99ttqzqqzRsdhtL+0zOUtQrv4qZzBmyuYeQFXnkyaohMXzxCn03eGy+
k0ywle6oD6imlCOvGaX45U5DXhx63YxtsBxf3x5LoblU4lz+8c8gF5Lz/ZJ5ItA/
j3kSso40zhzDRJtPS321gkp6oVh0GlKyyON8J8w4df0GPdOC3MVCfKF3BJIOFETA
R79eMQ7+pZG6AwLZIz3p0eh/4InKbzL7fSRnPwGxxw8dKuQUrRcxnjk8XSY7Phdk
fR9B9zS0VXmR4jz0I9hIvVwoDZHuylOssaabFMcfEAtfxADa1bkhA1AdXyMYj6rq
+DiLfmGp1Yi1P/ic92HAgUnpbTYuhzTihpg4L3SzOY4iiVQqKnBG68HcrY00Ai4c
tjP3mniSgdxLEg8n8F1TtQG/L7+nDvyuRmfXLo8+sm+QCN8VVbCGg3EI1H3lOFEv
VrdFzardZz1RjvIty+aWYp/SrJMb7dfIwO0q2iqp8Hpp4WHcT/VBJlzZY+cusnpI
Se0mlreqfmdTBbFd5gbEeUSnoQnBOcnP4gjLXUAbkfSNGzCTIrv7x2DHXKGQIW61
YTpvOLoNZDl2Lz3QTEjFs8WWNKFc2mmw8I/BU1jcREVQWJN/bS0e+ZO3gpTOxMI2
QORy3Bpi7ow8HkeQIM0966brsH+t3x65S3yCm8j3Z1XgbfnXvjJe7/A3GQNoaosR
HGvR33XkKqjrMqTrLoQhi9GohJ+Re8Kgzs4NQgqaCL8O4OIsz8Th76047YqrUok6
KtSlQ6wocHyEAqiCPn6mJMhF3WolO+auULg6JFoz6gXi7EBQrkDkWYzxwbpfYPnx
ROshjS8Po5oAjQ1bVgRgK+88C7IWN0PmljWFrGAsx5Mn9P2RE5RXbjTmBy16ZDky
7E/n1jb98LLkBiYCK48rkntedBuOhXYXzSkFNOJdjwkdafffNJg5AHpAVvpyCbXr
NgVucI7SuBIRCqPy7BNgeOaNxYGD8PoJV2u6RLr48j9zi0u/grJSGmLlDWiQreIb
eezf4nUPxG/3iTMiwilEKK3DGF5TprtVB/EiMzmSeqI9X32UmxiCauk3BOKJeABz
4bo5haoj0GS1RBbMrXck2cPJndFyfFfSIGWRdUdtG4O8TlKzcgse0YFLbQ3ThEy5
l/mCyHp+UuYO5EjXmn79ORIODPjbMWI4ylaU+si1WO+JuzlJByjktaAVss44BpUV
EQVSE3D4UFqzTEw5/bcvTWR9T8cbhO7Y6ZXHicKgSorEeblXt7yDR4aEiLFx//5B
CG8ZsbwXGvQdoYUHJIoNTSOwJjfSydw+GDBCrEztnCD+LIgq4XMquGi9cJXxnEjW
VQ5NJ9c3I/f8K3516PnbgH52uDMLSYXQnekxcg8EtDk0bW5EyQq5CRy67rSqOGb3
37GqgZ+G/+3EEQSa+i7XzbdZYX3tZMYtyqY6l5G2H7RRPlHaFO255n+kWi4avMrS
79wIpmEkWwe8rHlyxm0tUA/+ApHbVjIoMUFgKpOO/qtIWY3J5uEzUs5xNko3I/D/
IE6X58vtaEZvjv0WTYHOTh3ze+ZoWO6i6Mp4jU9S+0Ay2Ci+Do7QHAmgcHAZNncT
t7fkL6dYGhhGPJRLNxQfNNMOJZJfB8kxnOgPFSWjamfWILDX9ujlpW4MJFv4+NVR
K8KaV+N1F2x8l8reId6lQyA49cpm6vON0UrmahjHX/dfI31bOYZg4/lCf14IGy+6
Dgxf8169wDeJsFks2DrlfqMfYjPkYJfzRPTBzGCsHagklewLDFTcldPWqIF98ctB
Nh3Co50Kph/JwqLYWquluhTS9b5wxW+9W04QLzqqUp6Mev90ph+gdoFOU/61f+c9
nVfDfigRzfpEkEUFIl/KFP2+DBQTsBiwJ2C2gX2yNoixhtYLqwOxqsTDhf2FhBJY
aJiTN32antoVPZaaWHVedPzgTTL4ZhqGNZ/sdBi9b6kYXjilJf+Xi08sspWZUYBS
6S8QYjQYMOLg4m6TrBzMYVK58mgVK7RkGsgoHrOCOjutYd5Tdq6QxlZJt97HE07P
QSHNzWkNmtirGAFdJGQudMaJnVpK0+R5wUBizFXy3P63C88OeP+feZ4efgetBvXS
KGSXsILwWoGKhwVCYwi+J201fDrQk96qoGdNpB7SPkn9IqyxXOUHY+H4POKMF1kW
vVsFIl6rFBRah/WKfaTZcjpIBwENwWXQfdbDeNnMDXGRNkCZj0YwY/qDeo4bLsnm
VZZLOBbRdjkraFC4FoP+SieBZgwKK3HDhB7Zo9icS5qwNV5MSGFb/31W9xyp3Rmp
V379UUF7AZ++U/bnP6VGDO7J2KyWy5usyKMDZXqRUddw0i0rDjNUv+NBY3Szddny
vqy8B0jVJkse+/xBXmCSMq4siqEuLieppcc+0cDddWaaCnZL3w2JT17exJbDrGld
VC0eKJ3rOSnGV132pPHm05burc/ALi4L+nyW+lA3mhGt5F16uITtCNwWQfBsJ3cm
O9TClej/waR8DQuwrarFYKPIzcx99U8/45ZEZE8AxYTOhHggwEgwdK9XIWbc1iay
Cna6CsyoCcleRfbzAj2fHcWO6hDuDUyPluqTVm9RXZRpboV7SylO540QS+Lxyo9k
ogA8geXx5sY8hgcU82ElJpNsdd7u+JncCoDdAs50Ydvr7Gzbs+O2aWssLm31iSF9
KjZaajf3fbGTMEm7H042fbLLVto3vcdmTnpiBC4uxOeHyOw9MYBB97ha9paEhNM+
5bKKJ0FdONQpjkqEraW2ln88MexHlvNQu7wVVpSCcZ8sa7g9gU0KZEXYa/JD2Bcs
NTeuioaBcHgjXNCCxqTjITiDXLqYg8T7zetqMqnzShrh/YWxhc/0+ANa7Gwx+OW5
CyfUmdKDPYUVAm1xsrRPFes0oaWORlN6r/QZfWfz0G+4W28Ipi++6BbIghAStkGR
w5OmdPAWLIQ1QguRXWQoX4sVz6xMMgm3CcVJvs4Ps3i1DtN1vQfcp53xjC2NlHwa
tAhONDXw86kPDmDA1Wjl9YGNg0CdLKHWrFP5pYnDpWMLYMSM/smpjgdXPIY5t/jC
8sqqxJlxH+B6KjdANYnSXmKoJ+I/PUJXcZx9p0wrhoZbm+4r9N/c8mdloWzoso1X
8EjG4z0xNIaafLqQf6ybBO4BnCl+2tgfZkhEWaG8ofh6Pkbien9hcfNLpxUdvmKv
pUifUwhMecEVmTs5LOxJxbBDV+H5N58O3r/plaOJCYP+JpciK+mkOhLzStpW/yKZ
Y9+iekubpvEZwl9xDAYs3585jyX4bLJ7X8pMYOzTcoB5Rurd/GStq8r7qlVtbcEg
ULq6bgkM2MFNR0YfCqo6P1atQSYDMoi7m10frcLyQED2D6w560WuXbUWvZRD9vwW
E6hdswe1HOIbzpIWOsP2RZ+hzhnrFzUQDUMCtejTJwpPkZ345z837hzJkgCCINj8
LBoUA/aUenma58ZciPiUGwtkYeXg4Q4Ahyi9zq0V75GnVWEh2yCSxfD57IHs6MQw
HzWFRL/5qWS6CCXjXXcU9c3M6Nb3f6y48vSoA+3jr6VG+vXXUnOqXWS2311LL6f/
BZVo9AZGwZIweKGWSe86QN3IBzX9EOI+fZCZKXgciY/eeDpWcaXMxvC/h05/rwkS
VjIHyH8X29Z52CSN9TE0WpeR5rF4vJibKDRXN8xzRLu8JpZPlpLkd9fKZSkjcsxm
U2RQkDhJsHufrn6x+yOf+0zopmAegzMNFqMAJV60KNtMFnvZODVyaOzVQxidx7Yv
EigKe6F9ABjUe4LXCsCN2JPmUJSLXwE+g2O0fIAyhsyunbqIz3MwQ9Pe03opslg1
WvWJ/qq9rdO597cLhnZpzLEiusv4kIGGxyLFl+7RkjhfUfRlbFYWc771Vg38uUDS
wcaOitxq0kQvXLeyaC23NgjV1DYzBKIOmbcsKVWHVbp6vwcKNipl2+y7HLq4KehZ
1YlNe042+XeaBl2OmylHrltbB5VgLrloNZN6OLQ5uQIjZiUU/C7YkpYPr/1jcRRs
pMYw2bXBPwz4r/SvA9T0DbmgnItlCjUTRxtiljKHomDPntFc6VpGQbrxaBOlo2rw
KKJfz2bFGbMycWy6isLhleEu3/3CVJ/xnh6hnjkdox5rTTBcKKOGFlSmF9ltmu83
qTGTM9htnXDEz4Q6ydlHnKG24gzoQYg+QZyhac44Sb6xUtB3duSg9CLGEKCCTJc5
zC0WG1dj8mDKabRupN+Uz353nAPnbnSpMsRf71mcaxq3Q0FKlDUownd/4YcqTK+M
gt7+jcdFe23/7AU9psw06XxoLOsteG6GfCOIeeGbs5N7Ntp5GtoifH1aq9N3CyuV
zVqYW+I0sTyFfFtbowSbwfRlIDZOqpxMIKwN3TalpnvneWdeKXAMDpkWpUVmbGhV
/g2XgXVdAkJxJ3Ty7UK7JZzd1Wha0BNX6KYDW8JeVeE0B+O8jIjLbKrEBfZAXoOX
XPMDqxIt081hmeJHHsKEzmUScmWOmznbNky91fQDz/aULoA1yo/mpT1kRps+b2p1
DE661CWHWZv5NkwMk9frN2Ssk/uaeoq+Z4ZFxcqDVzVnWtuen+ITaEUC1IcW5cmN
2sYoOgO1QsfjqjdMZZJGwats1k/eM3PIML7TgV2hz+VWCGvyQ07SE3wVYl1F3v1A
AV6/lDd5hwynKr0HEMH/TpQpeS1RcOVmfEpFjA1jnpCFujhXe4VDcd2dotpndN86
RscVA1+Jpl8L1OpoOw8FdA4MVLEuAfSeF+OXsikoipT5nYW25DaY+HVuJxYBKtb9
ePPn3ESyYAj8Hykam8cjPlI8MZls+71uzeiBmLbGzqvzCd/z7TtaV5i8m6zTampW
X7Vzde29FzFBD57g2dtF6+VxU1FTIzgliAEDIAv0uloN5a3azXNQvw9rLRLdqpl/
7puONLFxWw0NXYZrI8eX5zwY0OHy6lZ8t8VqnqGWphMVUm5Wxp82qN5uHZGA4BJx
+59scy6McvLTXM5/eaewfB68K6Sq5UPsqEruKNBa/hm6c1dyXs5CQgjJ80x11y7h
wZiUjJpTrbm6YiT9abk3N3wqpLCs2hSmkZaikX7fhayclAYeIksOToU2LLF9wt6m
qtFaBZL+hzm1v4r2ebpARth5rO8HCFshc/uEJkxTZ87er1EvXCFxI7gTW2ksRIgy
c61mhVgr2t9I+roD+OhUpEkjHXgoorWyeKQXnvk5tSCa3hgUscQU6tbvJ7ULT7Uq
Q5aMi3jnWmiriI0T8XmVhjut6aPug5sVy43IDkp47wDeIJyTdNKawI0SmGOTcFkh
/T0PphrCkHpuWX34AnDRDfktW9W1idYSVseWes8um0XW+/4ArwBgH/qy2an7WGpu
JBemxVuYydj0C9/qGx7/xOig+y4Q4yJQnIGioZLnffk/ABPdbgFXFci1OuynrUO5
BciSUpOT2y/KvY+1ip/bZ3M/8iXetlyIZ2FCg4ZkkEGbakE7gCEKk5z+2RpShfVt
6xDPsxhl5viXw7TPaa3wdaslDQdL//rES0q2UFVFfInVFrOGNno9okJDYZ9SdVQG
NyOQFt4uBq3wDsHwk5khdVSOZPlig2ya2IbC/XyagGGdiyAYTztWxJ8Xncx9TGJD
OwMHMJkTHoGlcox0QsubJwImq60ACBXdJ8oZ2t35zji2XQs0/gzfuO35/tDjqfW5
uFCpDRAPEovWZGD1rJHEL/1ujlotvmefVI3rLEZ9yQ21Jb6N5MDnUr7ukhF3UEJS
qp8ryUTQZyYfVvcxNwbNfwLMYTE22Fq0ANll6uU3wsbNX2TrieO7igvl7Yvfuv6t
B6qGMQotXI6lupeVnEyaTkMYlgmQIG8TmXlxPiWeUJrWab3x2QoZKi86oM7vJILr
yTXASEXL+U+uo6Pb/bRDjUyO0p77f4olxsXU1IPfhjwpZZD14CrMpOGz/Y04jCBw
qYqthBTsv225C91bzxGTCqDBqC+Svrj8MGE9i+YbCElUarC+FzTHY4196vNS2CZj
EylwnuIbY6CbBtywFEqWPxMmcQaz1E0QO1vGut/P2OPYSG1PlxZN3Y7W+spzkJXV
De6H/G+esyyn7cDzOPsm3hj3awhUmYckcpYb8bEZ4SwaPfyRJv83BrX7/eLbIMYc
efbBvWvURUuIEUk4yObGjAUhs56PorDgHyYD6x/J9GUuSDMqxmCm8cp7AQrt+q4O
7l+40BTLvusIDc928zt1MntaFYvDA5o39LAiuJHig/XT+jMu3hdtI2tnnGvYeHr9
SB6haFhR8c4AfltKNEh6+UIuIdgCY36Rz94EuXmivmAJNKwxgT6XGdaLqBXRclrh
7j5M2NY+PNYILo6oALPMYZRAtdJmQ2WbdJekLSXS6bkEZDut6SatrX/kjbB4mr6u
ATBGZZhQLTrB9QDKh3QEM+RRWqrppF/Ge2arz8XLii3AMW7GwIqI/SSuNIFtcRWJ
7ATjVmzggHtQ6gAV2O5SDmSaC/LuHjIn2HYomN3nZOeu31KG4v+ZXz9RZACkCfL1
PseHAVGU/QT8wX3cMM8IGMwmgX9S76OrhVhU7KrEt6o3BIzEA8EKGpp9ynmXXkCY
OzW5ne+JKOKtk4a6Ya3GsWfJ9f7xt/gWGpqvXafMF4edvzqUlzcTr+KB3L5j/RKB
8Mm3dvW4UmZ2ebsYvqP2K7kg3ASva4/hKTKQ9cZVD/Q4kU0tJEWJIdIHavFySMYE
c+5hTmuirfAflgcveQDf6byLiDaO7P5mf/JW7HLFvVwXalmj1nbE7psXLB9IydQY
+M/LpxFZ7HPe/0Sm/HNuGKgblyLJhLGc3Rb7A2T28n/pNgV2OjRiT/hWWWT+qtpE
3/FJeEft7CdHGfdUNCPgff7C/cWKzvdYsSfbocjLne4mOTDC5GUmbDaYKGdYp/yG
Rx0WSbScsnCBp+MVTDF79TZQ8k6xW39NnRacBpED69GS5KEgfyJiTYvnqLJrgOGQ
BCGmNjB2lF93namD3lXNSi0ggNdmE3urC2YCWEpvS7wVom39TjmR3OjZ0LVY8CNm
M3IxiVC2pOMgAnCV3CxM3eGBJ75PrwbzH1MEHH3Sb7Db1pQj7r6TSlKdkZkU6VnE
XxSDp3nROKAk7WweSARkwVv9x9rN5iBFk/gou6+HY0rLFfAniQw+O2bIRpoYeUbk
2Zs8OXh6fpro3dvZyamjXyhc/XPorl9KkMurFRHBtsHze7qSnEYAuTsz+AS6eANP
gTQTJg/Gqs7G8XO2jxmtos63YLgOfmWl7Tt+zYz5FwwOxIGEbuC9f0tZVLOg0g6r
Y/gsCX7rhTYJUn2MhIOcnlVgelkov+d1neVS2dEEZ1Er+h74O+jm2c0cgbS/KmqE
sbkKhpQ5Fd+Vxq26uFonSBdL87MxfOborGLEQyz2fbiQbThcpQQJwuqZIj5xvvzZ
OTOIAnlEClAc2og4Qn6WNvQTYZfkQe4UnHLqgZVGC66Fs/XM/gmeURo0epYqkNq4
6/JAkpC/4RhXVQhQoqOEpPQwgxtWvtMoaPP1K22gprLBomZ04v3MynIjug0JpRDP
vwl/tDCUIiEIQfYMROUg3F5RmEdesD+fe8tzO9EiVqQAEsmr++okk1Tg+Ybv+8mR
6C3GipU7G7aqlZUhY6vPc7NSXeaOoyaR/0dW+TZ5JfQJLgwSI36WT3pxSoKHGuJ2
Ce3yQY2IIMP8Nyp00ecZEEYOZLWHSOZt+QXtzYNYkDSQZ6M+NYRv9CSXs07Sqs/c
X37JMzY2z+nLBTCngxhFgiekjE1iB5hQAFtD76SvR7MDebay6tIc7MOtYudYRrKW
n1Y5ORpCwy0UdQ/yT5McHZ08wMuWWM9/1J4Q5dITVfAkO2OjjoOpomdA1vGol28E
iwoYYUIhG+BvijkXqvs3Zm5KtHr6W58GeHxSP6rvBOwuoMmxoId84tDaYxJ9bgBg
OxN1x+VcG3Gn03CxaeIf0Hmyo3s6U9YMZJaMrRdiC9zUvzBXt6J0KROO9YHH/WCG
2E2ObD52/4xhcN7z8KrVw6GQlbhUheatXU+jNIrB8OsHDXPE8U1btz21K8qtT7rH
hf4pe24h9OatG0ZQOMEH+ptEBWuFGvXxqcDD8jDTyYQ0fkFUMonJd6C6T1azYBNS
fbXCb+xmVVXHub42ZUAtBlFEHUFAlN0Z7LT5Xtpxq8Ev+Aam7OFiXBjJMjVKqfxO
4N1nvBpKhzspRD64ZkjwoBq9HliKcDGJCzS9vkPn/CcnzC2AN3TqASR6IJbWCScq
mEtnq5LiFCrtFJ091HIdS/2eFSltRvfYpyoyK2m+ZN86n1aQPaLjkC2ZM4Q5j0Ye
YnQeNqOkFpMAW3jwMszuELB3D/qgle3kVFILBvcI2MZkPKs+v7SspqXyfjq4dj0u
usm/90vX5v75qZvpDLRT70zd9/m7VcD2BU7H8r7HrNwymdFxx2mP4IfGHjN/KUeP
CWWLDrhge3yKxwJtLCyS+qhzZToYcN7+ptcaRQ9l7Zi4tEao1u/UCTwk36+hvTjy
bDpYXDdgwOHNjt2LuPPBwW4xwd5CSo7yYi86MdvR93sYJw/wtn/l1Qd2hebbK0m8
nvogp5b8oBEsB3I1tBb6ZpU5bl/BSRJprS/aSQQC9laUhecjzRdtoWluQjHbbLwU
s6bcR2vJizkUel3cXh72eacWnZkOQCe1hRNc7ixDoOXnw8aaoJ3Q0vf9PCsB2i3Y
SJCtnb/sb+LVwS7gW9h4KvUWe0kdbdOfsi4HcHCHjXfp8xyyS3gLIZAiul3Bwme1
1HeiVBqF6Hh9JEEOIk0bYVapQEjxElE3nkKXLLoOpcR3yP/ARzm76Yf6WuFo/8AB
pE/kB88ukg2/IpOXDY13t5azJZ/4nNmeRwNnm3xGfh9XJcjseuQuSCV0n1ylRq8p
14EMH+DO1228UcliaNf/kKT8Oz6JN+bmWsfSi49b4yUcZtntqilCmD2EAL2iz5/3
emlP01hScYdKlyc4wnIReUhrHAb6Pkul4mHrSsfPJXOMN07+ox+ZmZ86gvrTx6VX
LYAN8dXDb1pS7J2qat0U5q5MXKJEmnlvBgN9PZtBDkar2i1+QYHOCFSsqdSpPykI
t5E/pj6damjmDfbPJjZpkrBDvcbmSE6pZ68SfrQpZGAPs8QfDRSDxWAWOKrxToxM
RmmuAxb7TR5shK4DWqf77zQ+aV+z0rzVMsDN9tKpJHbrADPRI3r+zHbG2rC6wI0k
usj7FYg6waJALTPHt1JFtepqNdBux762afbXJ61kZFcIg20Y39kNGPeNlfuQQRGY
CNTp0zhG0Z3ipZMKZx4gcS027HQuRWXVey/H9oCctbMc/b3G/wTlzDGkJfIw6JYH
gi4X3NEeVMOz0A7oF94sWdewqFbXE26QnhNlorV0OJJl+vCrvU3EC6i+mMbBTlNz
jf7mxFbQOzO4qs7dec9SSsPESKplZMRo5hn9MDAvD3BMCYsxGGwpQvSdJhzjcS48
PeG5Bz5/WzOOVidfgjI2OK6i2JpgeorZVAEjeXOvbqSgFhemwgNT6a6FuXdWKvDP
kMB/Hn5+q35im1vEMAP20ePLrmmAooMk0N4n/6y4crrRLBXb0pOHlGDUvdDNPJhU
zKQc/7LOvJ5z0eecl7ki8pMpEJ4loGJfx6tyebN0cTID5V1rrCFgWn9Asl1T/btc
/v518FcGV7SK0mxfZi3Zvtrb1HrCn9cBUYNT8PHCBbGTaMD3I6txt7iEGSgZbihV
jfWTIcuvcL0R9oxFZPUoCh3VdJ1+Qwr85PL8t1lWSfynWsRnwpddIKfKCnzwugy1
dUY2ry3OBSpsosAX3Y9AXEDA/7+9jcXasl2Uy/eL3/+8m9eXH5dWIKTC30V2mPoS
XLSNclehYKgYaY/Ck1PB54KQU+P6n6UlIc/fd9ixG8R/BspJuNUPUmqMJ79szxqq
yS4QuJkgAF/bUsPFD0wrfwwrug27/scXu/FftxwQpjohtjLAJ4IGYK6MsMNMYfBn
oK0KbX5m9dviOIqg+VVMpVjgTv0NvmIe1bArq+FnKRz526jGhX5M7i5XQet0aS/f
s0SCPapkgqhtVm3XTZQ2b+BZ/rRCriWf4WRl3J5HfzHl/+qlKpejMIMJq9Pf3nZ0
GqsLusLDzZbc/5ZWafxmsuZGheRrvBCjjehI367fMevLQzibckC4HJGvTBiiBYHn
KAzh0H4mBAMdfazFAMK8JHrJs6P9eCCaBnMF375fEg2gy6mRDn0vUcwdfSF+SUi1
iYhjlspVxuMJtLWQzpvMCZWBXjoBMy3FKsa4uJIesMKeLrQcXiywEWUF2nGCR82/
2TTNsSiqJuTYfQPXglcamrrIlaPz0+47b3l0ZgRhG9X4CaJ5ImhA5NK6iser4vcL
AheyVSmgXXuGPAxYoawAs5Pj9rKpf2nVNBp7p1Y9oJe/ds3xKNkGd8QFgtloO0Gr
jcxmozQtC5WsAOMtYDba+h9WeAcZROZwx9jpljK92jwgwMjWBwXsW1CZLrENplsY
4hZ2eUi/i9rvfFgNlyhtp5zuR8QudzJbx0Dbkq4wGaj82zh0/kMjnC836po6iPn1
v9FiaXfDGOpMozWULK4t2Wsl2gxaHus89bAAklkzfLD2FCSsOXjbJpHnNDWgPsXB
Txkvh9z4UpfSjt08eSYNCBEQzmG127API3THdXhw4j3C4smrs2ousJhfQmRb9RIp
Jt3lzyINuWmXVTTeYwXmUAwzj/OXXbZ2ig+vXRqNgwCAT5Iv11vQB7PyIK9aMzIj
EgLOaNEoRVZkCnKv2kU1WlQ4s0TOdSWDQttys3+OGCXsCzlo3mMy7sqynh+DiAB4
iikQ2rDv8k7iQOZf4HAzSfXvuVn8STnZW6iq9KF1GBz6WaAzdcFnlsfkp3m2LCgt
a/dAf1VUcXflji1lkFcDWT9bGYwRvmErBJQDrg/tUS+bqYaSrll8eJcZyKEKrzMP
c9hpfWNFYWNVYEEPmr0lBVxOZ2L8FgdKmSE6ZLRaTC6N4aS9uYX74SGI01oVajFM
dsDPNsVAIdPeIJe31kL3v2t69o8Qfu04vBGgSj0artSlj7OW2hJYab0iJV5w3d0H
6c6ti9ByUToGbPj0DpQqtGZ7QavKjZQdqLuizHiUn/S85wwgv+DpnGr+gwYC1Y4U
J9lsC0aSj9epUcxuP7hSHA+w9OdMbzbyG7/3kuQ8uQhQF5WC5NjuhID9JquQwiWT
Nhy3GDV5gAQpp9oPcvxw0lqtXPQ5fyWUdMYLYhqT4cvwhtKRx5wZYsB+19foekR9
3gZ8LrRrUZ+0EBmaUOiT2Q8YHlAKerJGzddBJOrY7utfrVhSX5VlvDhKb1dytQwj
j4rh7CKC+CmS+ZtSQWrAfMWlrDbvBo5ixNpdrsoDIB9v+JAVprBSsC760UQLR/Vv
Oz3t6ofA8IHRLNfzxrXyvE2idbmc66E6PNn51FylUcga886bu3lo6ETRr8SPeDXN
5plDPW+o0JkAX9WckTE6+fP96KCKr7U7SvJ5ew3XvgeLoMcF5n2RATOvlj8fE6LN
PR1Z9wGA/Wcm2eKHIJ6pIX4w3cKPbwyqbd6UwufJIBYgz+wzLpaprWEzojlB592H
I3JfMMkOrqLy0dVEALh8yb98aGSaFpqLEqFi/dOCc31sMeJDhMQ5FeBVCTFMK7zL
ATM1tKYzykqMM3tVLYaaHAMGaroLFL7KRe08L4B9O2z9XkNvkVgljQcP1CbsvF7V
Mn4ub3A700cjiKe9RQzfpepbY7Lak65yjp/bxpKijiFT/23j4KkNUx3rlL2gZBTI
sNExN+CV9w8Z0CcN+hOFLPlK8kO4Eo++tKtupZsqaNuybBCJdb9B8PvguO/iXNym
YktBB0adDSYintVG053Omu9JugjpAe640AICiCeTJiyrVrsLKq4tTBxYlnSGZtMs
PccYuqKNYNmO6Eezy04JgFMzj6MBVLvHh8Rcb8ou4W/O3o3Qr78Y1FW707i7ZiIW
WMHLVaSWMANU41NfU/XykoHlgV9FF5jf3QmTl2XXX/CRgXXfSKWfCmvTEmDSQ0LY
g4t/LP8csyd2f9DBry662t0V8Go2O1knuhG0JTkMV1sZVW5DE1zxdm/wgizlJx4o
bKv4pWZNV7PUuoWk5212N8UyHeH8aZp/mCz5aHi4gtQiDSOIKIxyhKXd6GlBKToX
z4trnbJ9ZhwjC9FwdPB3sVe/vGMc3v2Lk8rWHOnMQvWv4Qqf+7iyjOGvsc6R5RI6
0yODF1qBSs8+Nr0XbVUCXmIPDizSMI87Cu5vQt6Np+nBN37cDkPYX0o7h5PEJoUl
EQtuyOoTCRvyND/rhvHfdQqAb4BEwKk6gPnUPqJbfHzwBaFMlme1yqaFAFEqDPVY
G2uBo8o8Gl+1Vg665xTrOcSrAUto9gRSAntGIuEuuAutD2FnXAm5XLRn3mTDSMMb
d9MUzyRvm3XvFrBg80ZA1n+hZUmA9WWPxHcBf1aPuDCqN3BGOtUzqTJewCpz/Po7
99zPcU2KOur/W5skmaGuUC4Lkwo9q6BM40ahL8FEtwj4Bu973dKNoso+sXxxZQXG
GiSg2Z7HwBHnET1fFLrHDLJ2Hzpp+02ew9hpwxgWkYJfhLz/zL7z5le3wnhzTw+k
ZjBWnoPjDwYyiH0UpGUrPyKhn/tUmmOiAg/ZpRgMHcCBh4+L/oBjARKy6fYN01yt
XSTMnLV+xrA7eX82rcM0leEIiViEVf9tjAu5jRrecyYnpC6OTtDxpo16hudbWk/M
Fc9BVWqwELrHiE0HwWGHQ4BpysJGgPPrimXoVW3/98L4HPBk27+mevo/26KQ7OSd
3GOAEeixcVCvzfCkr0HlNJeawL1Rdoj6x5cA8VSwn6KW/JDkjc/lI5KKcHrB+fu3
I2EMEXz++Fv1ijENKpn+TO5otApgvvAN/lJ06R4z89NHzOUoSrWahAEUJydC70rK
9BRodnmnkdQ4pZTLVeXf+6iFbVExBRBYmSMMTsqy1vhn8nPAXgRaVZLqYsbvbsgz
S29dLc5wF/Z0zYl9YKBTpM2RiNCksWMyJ0d7F8m+PxPToIC8cX1TOIm1E3ohEyzh
riCf18EA5ROKBtNVS0IHlLUmHOvgrROG2KMWSvd0hYfyltfzx6nKBVB2VVL6Rong
Q7T4PUemeIk83Bl6O5X7Ts7R1eOtE1m3NgMf2lQbv/XtAu0BFUHX/hArDC7820R9
NqU1I+s2ZzseXr6dujzwtbaO2oKnWjE6lg4YM1JmbciXYmHUHWljeut6qwFQ0PTw
Z1sy/MuZDPkw0Zoue0RH9QAAa1q/kIAj4JkAkMkTKB4OEwjQLO1OKMW1eHfxZQ8z
zn/8Ce0GN1fqNt/V7zFwzK0Uqo//gWOO8bnq2BaUMEzOkXiNUcNdRM8UOAQ4zu0+
48nFOw/o3Ftu0bgU9yj02AWZLmn32aay7yDI7GBQCvEaUfdDhZ6OtQQ5h/DMQi0W
+yJVzvs9kZqFWHvndMJr86W1yqDm9bEvFD0IVSRzi1z3PBNCOnMPCRlzpLALcZHt
dzKweXZBVyptQLoHC5GW3ZxtenXS1YWh3elM+mjk8fLv7B1fne9/TCM/nFpDKRh7
Rb8ra2Mc8AEf6b34QUQuGPm5zE1SJwkzokwgO/7UvupNjw/JJLrAayFv11VyP/w7
WxObLcGnM2AOBOTtQgJVioM0gwl64tyr7kHaXk4pmejdYf2pvuc6d/ZlGJgIqcmD
7+Jsoy/nnjtEEw4BFj0im3IXfmeDeRBJdzPO8QA994nSM+kGYcG+2LqKGqbKH2Od
kr4gEFTgqjuLviCQElDPMOVvYHKwq1lA87hnHw/Mw2njJZ3chnN34J02i2LVbaCo
qLKkr6I7/YOpvxzY0ttbcvPM8YD5GAdzFokGeMaIXhaDJ5gYJC5EJ5a+AROTH47K
PMsX0tgF0bGij0EXEYKUHpJFo3zPUuRghFnREN94vPbBsCPViE6ak50u09vR8r4e
VIHA53/08y+x3z3L4Fqni5doOl67opUiwLni8vtHuF/wCxfItwPJHseOTKFma83h
Y+NDTMiUGtqSPetpPURb2inMUdSlni9/9DKG88/RLdZvA3Cja7Lf+E9XNNYi1/HV
YEJ95vS1f9fvvEZSnXhnVqlF7EVVx+0Kt6IhFtUneEKfsMNt6Yr38de9DNjuybdH
fTToTuAN0EYKOk2VKoLL0HbxZ1d9W0nhEt5WWtO4P06NKOYXwW3irHc61uNQEK9I
HPPHdeBWlJ5MWoecv9FuPV6rGARRUHj/p9+uWnW/DLA0CoGFkh9aU92u9+OUDmDu
gvyFwddvsNIef5/d/vDLOd9camtAWPbURFrx755jC7gs8moBdzfJtEfU2xT7tVA8
qIYJsLv5f89p6JNpai+og6x8keb9smweGKQtCYRR4wuZUGc7kqheKy4AhROTnSvi
KG9HsrePwvwfadVyCZ0QWmdD6HauctsZcFFce72Ofit6jIWEMGqXojg4cC9KdMXQ
2R4qfaM7gg0aucvFuz+qvAscEFO79h9pO+Isy6RrhzXZg6C3Y0quJUQ6WOs2WxlZ
44l9yricJaI9CPkH2Hxc8KXaxQUnoB3d6FOiWJ99bMNc+xzrfldJpwX1He6dOVvt
23QjuaOmSzSoXzUdTVqPdLSVOYwEscMrtX5t85tcW/j+K7FHeaVTC9Zgano30Hmw
1oUh/F7oDifr0wGl/Zd/6AnEUgNBaTMfA5qlRUh6yeyC6doPI5heNTHnsetge8Ij
1qz5PMBjybHrYxURP19SeDAX/nNhhPwlWdST4eg91qViUcb1GCT+++EkgoLAnaVo
Y67TKLl5U8XmZH9Vb3046eLIp4Iw0XMenLdcZR6EEKV7awWkUfhgq8G2x2SMZORd
h82AyFyjUo76B2k6OP10jvtdWBaEPd0dLjqWPvovR0KTonGv4O1HbhKskLu3Xp/h
/1YQ0ObGp/m8OQ+Fn5Oh0L3zNiG8PbZuXCnZxLWwEnOwKtywdLC5Ec8SfvWK3WwF
y3WOBRhZZ98yw6IYpkpwzjyO9DcTmy2NhFjWrxFOFV3FJds80wWLkuSo/yBHNbAu
I94Sy1E8bqjGHuyY3EQQM0PJ3k/jfTi6tirV8L2aRAp75lD2SHiOUkz6ifuVmYiK
2RNwsSus7nXsPeQXDcLRIFwteIKiqqFbJdtmRbwoTHXmRFmSQCjet/eY6R4xMtAm
C2mg/OXri0Qlb9OomyAsptHLkEcqeYn7UbUwIwFpoHpXhZZUgE6PFu1Vw2EkyRAx
/ns2lUyucydAX4akPVPexXPy9lmId2HNURabZJ3xPGCq5TxNpzM/eWIKshMscrRu
yNgRJM2i0/obiDdQyCDofH2IaPcqC9IgQv28gArPqZZb96dXTmT+k1/YpmZcokq/
ZSQ0k83HcQSm066FePaSD6cW5E1HVIUR8C5PGAQlc46UyEMmapqAWGGK+qbn/hZS
RvzWAtBKC5U5cYo46ibgL1zfthPwfcj/B4ykWwZwXcYYE5AuBtDd5cc9CpadqAWx
/vJfgZz/C22eNT7M76JNq3T85EJyGU4uqM4CBMk2MDB6CA/Is420ykpoQYEZmGQ6
poz0IepG9xMjsLhJBu0rGUx+ikOB6Vo1MAg8/uUd6QdjPiVUFPHmajY2H1hfZY+1
eVbh6iAaFQxk48pOv21WUFujKAV+/qtC7yHboK9KkqXZrWXvUKUtTh6tIkt1MfBE
8aTYXtVeOM1b42bdCwo9iSBk8O9P4HG0VwyI3gRJdmceokbL/LolXXW4VracvEec
ewrQMjfa9XheWJx6pwaHMOWoy8PohmC54VedGy6xBnsWObpifITopUkav8x+3DaK
uJFeJusWPq6eVsRxEU2dqvVeHQonyQ8pP9IHIjqlqEjTllfm8R+WHQHmugHSdJBK
A29hmsNOHlIfRHZUapmCaZslb27hH1wQaDUSxwekDCLF88J8DGDc0joqzeOqGksf
RTLvZOZZjMwbQYLh3wz1vhnYP//PHX3bgiQkXSwVwRcU/w169MY35O2Z127yL356
prhFF0S4dDIx8VLnp7EBDhNFSV6NlYyvpwGIDX5F4tW6KK5+mqbzKTuw1eGh64lR
h/FarzNYsRuvsQFbBwQafPPklvuT97SuTUM8vAuIBoSc06Zn6wiCxoV5eFjrmNWQ
pDiKs0blRD33g071QaQBej3AEaRUpKW0kWanyCP2onH/Af/6BAwo+jL34SazcG0u
eD4cLeHE9Az6WjBuQA+OrtwmtdjuOwOvOUntxbpEb1ekucyn0w4hOitUb1b2g/sA
nF3SdJlUmrPwXKvdN7seRGoWF/tuikcKQHWIhUoFmSYYND0JY2M6JDSU9ZaIxOBk
hGl1rnA2+8BpSHbrehU6hKUFsdspVYxusoxeMpmZ3QOE/hw7mGoZV2mPyPhEa/wy
8rxWKqN14ajD8yMdLRjaNd+0D7QoAWNBT3aGrVjqVKdIaRXdViM4uJk/lrMJ6l/U
oDHK4vAWTEFDV9zgDlnMFEDt2xCaJWPzJ32iUeqA6+PmrTGV1tdr+Yss56Lh7n0f
KzL3kVexF4sWH6V43AF1NiZY21sFdG5QllgJR5kqDo9OtOQviBjtFjGR7TIY8zKx
KmIQCA/yNXzSByda8vM6L7VluFNh1Bw4qHsBrwXS8SCxzovHRvYaAZUcWOTUDmyy
hRdYE9v040q++DDOaDGPj1RoZzJV+9bTrcY2bA6AwbqRfVSykxdTWKWvtlzHxXdJ
x6jDgyAjee+VOconL7Ppl9YMqK7Dgc8PJSr9K3Y8pTNJf36Xdlp+nL2jmnHN6UKa
BhRPZMqXXXT1DZibtEy4UGW/fkp3oGKgjSBmmpfqO2CIpHrNUDltv8ppNC4cMhG3
hviMUXEwGAW+AedUHnndXFtEIIvBev0q9xmjIQwJ/3lFoBBv6hPfV60yJZ5bi6DX
emLJY+WwpA8eEIoJ/QZIUJDPPJehvcRQd1b7cStvLqrynF0/AFaPdhaflnQQIJ7O
Ec2RuX6hK3MaK/HDmL9d6Ph+L48nDuU1nfvmcLUaogQ6gxrLTEZfbPCFOnoVS66D
X725FEzeszd07W/Sse950fuuaVRzLn8qlW3zCIEIbZR97F2LHu84bT6ZN8TaPHSj
WprKG2Epl+FGO2ar4fxK/8Hax17X9nx/ASgSIWxFw4HkiLqNxz00wcYFqYWHIo57
M+YzqoPcoLAvqIFycw7bZP4cBJyi6poYpnlHwwHO/HS6Ggg0uZMmaXb+2wkXg0NN
414PBxiSgJDZlXqYtVtL+f+2UpwaMfCC33COqhagN3R2aeVXj7TvRsoh7oHNAOtF
QEZSPF3BOed4K4/WTL8KTXN5U4y8DmXdNDR0v9m69l+qcfTbrqOiICLKgPbGy1fL
HarXxzOcSq+UDHMn+CZNuahqceofc0hInCRpOA7JZzVxCZ6AzG6l3FfqMWqjJ2lo
QFWI1TjxkPi6SL+j9GcEaFaHXfaLb92EQz4/N/phEKAUipRFDBLO1g7siexUC4Cl
r7uFPLWOvcJIkPFuvLm/Z9+8U0SHhZ5FVZc7Ae1XqClgfltXE0Pe4CtnYG/7jrYf
0e/lruBWv4l0pvcxlTPjT5aQmWjt70EdaeqBEPraVY6qmNwO9cPnsPLwxIx/TMYl
S/fEJgBKNdmU1TtmcMQY6etVM1PDcoQ0zkHp0pxpISrRbHfcJfN1eOmNibbaV4Dk
JsIxyUHuwV3Wcp/FgiELA08uDTrMKaYbj472D0UNQEryiXae077jKULLmGcwqM0U
D+jPEaeuSh7935aOQgluQGns+tp8clfB374+nBTx1dB1t4uwJWf0ia9RZ1+uoATG
TeRFR6StHcXvb/obN4aMDFOvmQTPuXZ/vkFDJGVO89riZzQANUZAWRkKbi0iIU3F
dSeLYjxptbMb6h4oJfc3mu6ReYT7JgvY5J7r+AeLap+jGSmvrZQgkIBdHCpuzLcw
UHbsm7w87g5Aa168RnWTLQkejcecdmQnQos5rpomK1fCuAHoHexUkD8zKItUv1cR
NyMKVTe5wntXjOLsZnAGAzOldE8B+6SnnFrzkVCDpGSm0VzBEyuBIyk5p7oP/VE6
uhcnrxZkkPBlg2Edne1nB/YjQMLIsid3BAM+vCtpJqjixXtLUHvbGnHUQvDoHGWX
gpJiWH4LFV91YRGlD/b2KltnBAy7641Vy2gpHa8uC9iUD9sNKU0cBjBHYB5BwlR4
7PVy+MfTRYHv98PD7uksKMp/h16x4ZFyRQGYLmSiyW+o64IZ0BWIqvKAj/dOwgAT
sSaSL9Z11d6P9gszoAIHi0tCx+ILXRhtVLqphggw6DDGx+dOXTQgBnVWsjagF77x
cUxqVmcOHUr8P5KxrMJYTFQDJfTmWoXyyozVXoK5x0wPd/xoYJZNAuh4YDcDtzfN
CSmXespL8SQYL+wK8XnZKLmYu1durQIiAfN6+RoJoda35WaDitADpOdbNvxHJARO
xxxhS7swQGBAgtkvsmFcYPnr3lnZU/RqSBgTyB9FxkKqBmS5sQA2AZ1uyWH12Bc2
SwBR5GTkXOmTECzt6D4+wvnk3E9+b9LO5al5i0uowPd2Wd21TwsP1bmuFUGiIzHH
0czfDyzsjBpgBe3/lpdtg0DghiK43gz5mHUzE7ZhOZjV7oQH6PbBlk1oopFjEKDe
q3fWlElrf+wNi5AtRfg3TIdCihHbjguvnwpX7mZMmnlr3DPlhVB7jPUasa4XBAMc
hTGuaSl/QaN/BJrHSEWgnWO9g7GQgjODrpZNXqHz6lbMkKQQ614hj9b7i9ijYGWX
3JHhKYvz/aby6iGv3jh3B4VPTKUHsQkwztSU0ZZ1gdUG8Za6Jj0XaJi1bKQ6ZOXt
1ZWZ0lIYssUGxH6SLb5MTjhXHuU+iQ8jL0y9AUdZv1oYvx7/rOzOUqAXZgG5AxN5
XnIPmgVoIqhQmB4L39yQMQv9YH2k2iNrqLeaRTUXKGCiNvpnFVrZUL1mcDgo9BC9
G1vLrYDpe/SQynkh5XP3E1Azc/HJUZudWLcAgO3xszVeE8eaTTfbKKjpA/nyNHWr
2fvjIR4ZXkMO5Mi1Me5sZ7wCvH+nMt94CNgYXO/EjYWBtAOWTh2gnTaNPFEKDcEa
ifOIxkXnqKm9ZdKjPfQe0LhXKBfkmX3i8Lp2JT/WIQja6DDDvu1GS8786coBbCjf
emNQ+06aFYPSdh47bNjOodxF+I6eat6WQxY5zEK5vL+1HZmWDrjzSIVC44ZcffZN
O1pow6JJvj9tuS+QY8j5uvst090V688JouqA/wYs2WJvggSSbbfCaj2/X3ZMJrAw
zP83Yg6jaOf6yjIZBaF1pBtOXSXhWH23diIPiKpf5F8SSZFf6dSl4bDhtQWIOAHP
TbtmAaUxyEUO4hKZYm5R4ejbdW5QxLPYqiSWXmY4mYJ9gZFTnp0ipibc2IVUW80X
rEkTxiTsrxP9PVX4y4x4M+4ujFbhT1bGldYuxsuYvjgnudkBB5nv+Uk3mXaktLX/
KUvVHMXZdu8wlao0UJb9VeCQHMBr7r+2ut1BIj1t5uL45puXz4+kfJwfA2FLzyXL
GQDVgNnsBIpSvaCsAxrODf0XTqhMFkJ9/g8hAfA1k/KU89iUpofiLw5kODeuUXtf
7/nE47kOSVxRaj4kzhGp0tsIAFjtGmCpcIL445svvMhKWhXWKk/TyzVoc7IhODhu
s6S5Pzxgz0f4dSnxhYVZgu5Y5POYXNapxI8/Y4b4GWH2C3ilXVhYrKZEURVtnmcG
FPnEOdoqiov7RDn3MK7BVXbVeMmlFCvxHZilE65AmvPM+e21MfTCG5Fz6mpdShyf
pauCVlZAaHX+NreFBg4sG+HflAGkkhwbMTZ9Q5T7HW0BefbAF3L/Jm90dkoRMWfu
bsVG1D06fM13+gOMWH5ciiKKMCiJNCiFctOkzdkNzBhfxlFBW6AFuTPd5JTx8ir1
/YViIG6IdJjlTQuBAuOSDH+L2v1ZySy6+qQU/rHhWnxSm9HF960TEo19yFx5Hd06
J1iNOp3k0RLVhHzzD23YQizAZHlrl3R5LoE9Ee2QUGCVoq6CE/hQMKS3BEodVCcf
U9VE/WrsfmofREM9eHcSMF14+9UOzAY+5wQuNA0C+upZM1WCzZfGH2jjbO5yhgvt
qdGbHji21n0XBL82rrKyZHzr9G3LJggZ0JXUICvLoxIxv+Zso6ZXnMLlwY9M41yl
inpFSgMgyhZU1RZrIxT5XLCSnoFXNp+lnxcypDdq/lo4i/y8CqjZahA1VDuDFbu/
pF4F+YTH21jf7vFULAa0FsCqhmhKVA2fYDTZ7jyfstaa/YbUZaEdreAEbKNNFYol
l/xybmz8kq2lArHb4+NmzD3OSmSjgwyd/C3vKzREa/UG6lIyRMgK6PDUFTgHdOrM
NC1uDDFhIEsmEUCmJgIq36I3rmOXm/BDcZa4sA134gdSErVRu+Bg1WVzQsRJ7v5U
PptTSySF61QGMMIHegFDIVVO5Jjbbg87XyjVy/C+AXhA13vL3E2gZF1jfJEOVjbs
ldWUlaM98kSlIU7dfJj5TI+/WU/i6lw9d7io8aF6JHZYtqbIiQ+y+U4yk03+e+Sk
2PQCdeKjbWIjNP4AM9gtQ0iFw6kdic5LXZxuSMeNNS73jCWMrd3GIp1qUL2uHpxD
hVF8hHa7HrlJp10yu4Q4jQgVZrzOvqjHdEY9qkij2kfUJBU3BMGyL8UXXWm5Q6Eh
wog5fW06WWTbFBjx0zsAyYQ5Oj6BmYFPYsDgppU+mLMgKsG+S+OBnJp5z4NBgI4z
I9gQrKk11SgUMtMNowu6ZxBR5lOdeOAUiPfUsbsbkefcsyYF0bnMPy4af0IhPxlt
N+jScnBgss96+6ACYGkQpnLNUdvve9qqJbo5kZVArL1C20c+VjiZ9GofzCIYV4f9
dIwtBhrevZbhQjXHUwfN7gFqLF6NicLPkYS1gzUs4SyLNolDu3EVTrlKssLwRLug
qSdU0RCWaJO8kYr/LoJGKiuvh9vb2zu3BQj5NV5681ibitj5GqW7I367YdJys7oH
hZga5rTp9ze8ZT5lfSkTa35wh8mWQBrYXglgQa3XTfr0wGQpjhHooJlmcuKlsVZX
L/ihqMM1Faq+3ApqsXGyCgTLpuzsl45g3gAT67OIB7KuqnxH0Q1I5G6GG6x8l9Dr
MNQ0y/z1XM16pfBHvPgGju344N+0qv9kCBgK3S1FDGSwCQQB0Zj798KZNVk6TeG0
ZK+2bKtLqmZ0O/5+RlBQDxqtdpZyVxfSg1s0asyRlk6iW8nIkr0z2EYOoEu7Com/
swNMvYz0l1H+ASxw0HmHp6wy7WdE3XAQvEUc5/HVAGaiJ1QmZtv2N2ep9InGnGY/
AgXBHZaplFtYGgZ3x9qJenNsgWk5TnW4frsj6DScx+I3tP9/F08bHsEpIm2gyzgy
ezayvKhWE1gg1iFVsDYNfylqjPbwVDgHLHU6+cl9kb8vHbLQo9b20SYpxEQynnw4
kf+6fm0lVKYxkRF2H8+dg8SVy7wxDt7ntn3pX2pIMB/9iG5UoT8e5RoM90nN9hMD
I75j8CUU6U/o+IwcuzYkCQKG8G5OtCL8ZBzaBxFrkAs6OlcLX8LZ/x5W0U0ZPPL7
YT6mieuTPI0qlKfbxio2013ADieGncXgb83fc3YIYYppIkzA9w4ujQhnG0xYJJAl
Y92b9gNjvyGPkqEqf+CgB/yO9fkjp1rpT8fV+wmqVg1NHOrVegbdEMwYJm7Crb4S
HgHH0zay+wPYioFxv3YffVzvip1fHrxR7PnSkM7fwtr/Tt71BosGuKHPFy5cDFB0
2DweQzScokDm5qRAxAzqFM6bxCQo3hZOtFXPX7YbBIS7TWrrTKw1LdDPbWUetzUR
F/2gG7+qEsBwgrJNS4lgxVlSizlCWJ/yf0bjkwLViNrIj/E40KuMWaZCX6IKbsnE
40VSIpTYGUrLWbiseVyCQnDziKkJfD9RIDNPIIqMY35qTdwXy66NdBklpw+sBoaz
zHjTHJXNhMo0xv8ppvEvN0I4pvFDvy9DlX7rlH1E+QMY64QWGzM3U/hxPJKUtUPn
YJsLm3D/bq9QeZqV5j2eIGfwgib3/4NccpBgt/odlXzk989ICGojhyepMyPCb651
SiPvkYGKRKiEwQ/5Tmx+sr/Le9RHlzO7L6BZOT5Z/JSK8HD4jdFVMGqyHl/FwwI4
cZCkziQB4GX6/02KH9sNU01QUOlIeoxSEYXcBpjFOJAJCBbC9rl3J81K+KecY1ep
qAO3NUP5OImDc5ZTYokbvQnMeBO+gdTAGIP1kHpyK+idEtNjruV0uTf4HqoONF7S
wG37RJ0yET4eeU4cOklsgb6ssWEnToRowvXIfNAhhEYzLSLzh8hcfqmA60O2eGbf
AcqO8Z8YgkH17EO9qqZHw0BYswWVzv/aiHgNqmteLlP2Bdgr2rbjo+8cMOi3k8bs
FIZ+TSRFtO6ptVIzWZgqU71MhLJyFujLu08vQfy002VfMgZvw9HLxSARcsy5CmF5
eRcgiSTZ8HjfEueTqzQR6vEBURZGntdwomJRumkEZehjRL4tT8WqfLJorrYLl10O
PSMzjqNyK8cwenBYIh6mQtASZSJw+sTxb2RaPHlbfirk5nKHy4Svb4+qUNyjOjBa
ujMMmDsr+NPt7Kqc83LGopedRNQiPv1Z5hwXY/jWuVWb8YpxxoEm8K/HeLGa2KfK
YaPs8zioMU4qS5H5ePbCRk4f3tRK65RS9zxplOb6kkEtWQTHTOAnt3yq24E/9fwr
9vn8MO17xBCzdI/2L9HNQjuBZKdSzSkYmWXHDMSYqm7aJmjDsT0qEqKXJ0uZ/1Wq
aAHdDIq8iQf7LGBAIVBKWlNJbnUG8a417RrIjKAbhmRJx4wnNmpl1ZScS9a2SFka
i022mLnRv1uk7B3GMn4uHSlMoSMav9OFLr3nFMXZ+4nGJ/RkkIqnCmWZC38X7U8k
yZ29zrP8qRWRH2vJgvuZrgxS4bJnAIWmgc2XuzGIcSuSJ0yBXcklqu1+b2ReNtiB
tKCYBk+fxnvaKnIZMu1/Xu13N/kmXrIvLxEwBvDhTJcg+SjHi5FvS4WI+pxBUtow
9QW43c6y6KSOklrBq+vflyGNBNMWBxbeGAh9LhJhOZefd20PwrYbawzlzHb/MrQa
4kzeF0X0UWpa/UlgDwuRfReBUK3CEHT3S0qPYaTJNolHgA2nUOMldNNU895gdUpq
fnV4lBq0QYXOpPNBC/PPs7HO5y6DcVwBKSsWlOJLcD6Uh9D6yZ2eLEAo0J7c78o5
Juppa+in8tls/CiOi66WJlW16SrZCUcqUE8K0iXqgF+UHjJ6rZimAfDIWZCE8LEZ
imZk16iJwQ0/0WMc+JI9sKmlwpyvmmFtgcjWHqprMxmk/+Pd8KxKl7GMNrIryquZ
Ggm0NEHX2bUEgOEcbiQVXZbK55vkTmVXFEpP/w0IlmTRcbEAh5IXyGx7wKUW0uJQ
61ze3EE0LZtbgry+jkBvCRCHPw+eRxrBFffPhKvfzSraeTyN5THimipjWAZ9Jt07
Ek3FDfGXG7tcoMqkopv241PMwKD7Btp1yX6xcvw8n7fk7a9OS0kHGfste1WEIlNN
ykHtUuLOtEWRzNGde8n2ooVa8b+3iS4OM0fDIfRiLepmfPrHzVse9nv9ymzgPFdL
QbfhpK5YgKuWjIvmttQtiXC5UYDfKj2qnLO3LaUzaE2TMzB+rUYPHhkkq+TONTYj
vbhA19JE2eusJ/vykoEJwc+VVLmYaWH2GSFEeFiUvmk+KrEDvzOYCUBwS6D3Y+5V
Zv698KIeNFAHakdA/fi+OKTK3Dn/bouq3rxhz4pZK0ulwBJBDZu59lV45wUxhj5b
kIqtINnC5OjIyZNy1DkeYRYj1tEWcVWzZF/EK+F+V5xFIq9RKmM4wD0XGqJlltyM
Ev8Hjbv7unLWMgfnZ+7SgBsGEfVuVkWnO7I3pJT3O4i1QJrLcnLvQ0UsX9n25Ybg
IwROdiJSJwoVrJQGOK/QsObxhx7k9voCMg6kP4qsSxl0LbCjtgl+DLDwG4O8kpl3
/1nI7C1A5ozrHl5Ap2eRrbP+eFASrOCkoA/4jBJ/zgO+MJG+pdWLvnZ/y5rPaUfx
NQ9Jw1lpICRZ0jGGeDNXJJ7Pz8f1/ojpA1hi/U5J5BTM8gI4sPMhcj90gIkOWbPU
X7YTel5uj1ojZWRX2XcKBTtz/Qb1hmiiRcKXwTlS8h7maWmOPol/InEM+qD5ckWf
n8HZXrjy0DHLimV/jorLbuknjMNKcQAw4gw0JkdUnYBtPOUlYxkpimTUeJkdIXWk
0ICNmQCvQp7gjq5+yMAX1h8jeSPr9vDSdf2ogDPwipTgrjULvFoydTumzQG1eAfE
KZbuphCj0FqMdjkV+hRlm5Ia2HvBCJN44fn3vfhhL33xFQD5k6QrGfwvLCoAe8WJ
rlGOcvQt644DaNisH9l9Q88Je1SE6wGGE8ZfU9kbU4K1STgn6oRmWAbWgJzd4+Ls
IX01oL5MbEDeiPpkKb1xjzCpl/FVvGKMGUd6kmo50PfEioAnMAZwhHpkmnom660t
BcTw6Oi168RDClI0O43S4muqH1a01GpnvfMA0yGJwC691V73uqalEhjt6Pwb7m5P
R5XFg3WnnvInLQofX9fdXkSKmQ2+UcA0LfzGz0Om/FHTGjx65JMihdhOCh87dNC3
xzAduTnunWSdc7k+9P20WKvDIYYFJXpG1Upx41+8qXOD8qgJEygmgqL/A3sPCrIO
Ls4HmASAM9D7VT5loeBA7Skrdc+GHOdGMqJ7LnAzJk51+BjKNJ3TNF7vWvyVeiBS
En45NIGqcZf7WISDZl1gyVxJeroXWxkb2n0bA5VM7eBqMa/cUUxzKWWoaAd0VE3w
qOetcp2l1srDVllTETSc62yJsBq2Xybtubd2B4bOVJbSwDx8T7J9dk/wDyotoCpE
ilA0NEy4bzA0IWsF0cD3Y2VpUogySyevmcv/1wSYrBWJ9WhavYRkXbFpOWM1spD4
vWujqsqr5Ofp2w2QF5c1B9N3YAleswy461Ug6ychB4UqfZvt+EZDCaToSYFq14uW
KzUAuSiYBovqD7J8JjMGP/5n8YppxIsvEQBr+LBiy5tre1uJAnkYRRFsGVwfE83B
69W9aXfeqgeC1r5FVaUcsj9hGAaxgOYDJQqaJ9s9WjFlP5XddzH+bDyk3URnG4K6
O4CBd5OA7aShnzjpV51aB72OZ/nfYeB/+ERP8GExe6SIFGVhu8AoXue2C4281rgR
Xlr2sSQysuovoQ4JYsQbp2vyrl/co37Cp4cFXs0OV08XHEredutpV7FyavyOnSUb
XPDA317a+oND7rf6l36WYr8/45xeHoS/u+AqiJ+vBYVYYRah3lOXpE/ttWk6U5Ye
h5dRCYexKukNUM722R7Stc+BZMft/es/a/2IpfYWAccrcnKut9oGnFd9mOQ2qDiv
tKx2fv2zBJaSun8/ZVqzNcfeFETN6CQ3WUECiD9aCNyHHRHjVyplOnyFDqDcQdtx
5L87SejkXDiXmJyRxaRXA7iSOwaOkR6Uul//IZVPKPcyvfvsfjogUKUZLrzN0110
RfdSDOphymvpnnfjiBGHYbkpPivGm63C+lzaZGeP6Lonc46zyyCU9UIfuhZnlnFY
vdKVI7Ma1/OgXvZ/WU2WkpVjxNCu8YOcazAfrXsVUp79KIOcFI+EP8xBlQYeup9u
JlEwZt93a/R2Uw5BJKSWmqfeC4NRLJ8POO7ePHrzrUkRGHk1H81KELPtkNNRDqB6
VdeNTC8nyNMWAwDtxtUch5SfDU+xO3k7SG7Dg34EiDGzZ5F1w1tBkEnUOZWYq9zO
s2/0XA6NqT5aG4SiYjV7P0TPxUPSkQ1fYCDChAXPrtZPP/rwU9y288gLBovk3Ype
Zi5JULURgfFKFl0bDD7ty/Elmq7VSQS835yTLfwebXEJIEUeqtgNJrHXrhqx25L0
fGJFkUQHzf3JXNWs0LdP0KWBOBopSj6eIOz05DwL0S+x1v8pLT9SIyXO/g+xqvRo
Z10KFWyL/fbE4M4GqrmsWur3VLvziI+rA0eC/3Pd0CyhMAu5QSEoiGiE+3Kmjokq
pH1yt+pnZZG3cvWBZbpGEuaLMODI5nQ+5BWXYLJZxBhND00xTsZEvlQSKrh9KnoZ
VHaDP5LmiVcjgdLY9J5gNYNK3YpM11/vUkFFeLnKK6BRa8gkBsotlRye5Kb2YaK/
kMJLLCudAo0eiDzSOFtYe0Rt1eTYqma8KOnwVObGWywAKQUErgaPV/CovNuua5Sp
XfVAtrC2RRqfGN/jg8gbdAcuGa85GR+VBfxHxwp8rdYr9/BC2d36vWe93nnVYQ83
2ETC0ZCAivsREo5Gb/ifAvSSfQI8ZEXMYSwLtvlHVdRQBQmjdpUY5dGEdJL15pAu
4dBKxJu2izj2S1D3r6ilUWm3Z1q/jMO9/+vOnPC1quRFWRbCWgg+Pdh1d43h3VFq
GhiOJTeYnBaJ7cyIPYFu4xVZzDAJy63MB81CDH7St++aooKHajm1ZH4kMDDPWjb7
oNrDA/5tLxgbphZzTvssAzJTw68YkMUvEhYeJvXwgwUgrecKwILukj1TSzcmd4lP
ecOFxtm33iU5QdbgTH0FgUMZCoUD1Ao9QwTKGWRjDWm6x8VBZDbQKWRZPtLj+6qg
hPGe6x7HzhSxUWNoGZ3mFfvBMUNn4ikepDLjxuo3vbzeTqbnlmOqFY/Dwf2uO9J1
irAbxpfG8R7yxxmNYYnMAW8WyWVRDoVZxtrPm93/2Ib6N3EgMusFLOZl3l/bns0A
K4XwZyf6atfTzh9J/KPpOdmzSqx2npm/oLFsebgR+w4fQS0YyzOISkNQNokMIbVL
4qRk/05n42elwXQNg3ECUiVce7EXbu9Z3rBk3L/861aKrYHmm8J9Ll+tqa2AdmRq
mTDtRVXZ8Bd7ZerwN92SoMjmwMCjk5B7mQEiS1TlLyl+TFoKqytmDxruj6yW03AN
aOT/ViQxvyl2X0ezcPEw6LpTp0+naZgmy4wcKybOfoG0zjk5GIAa9fx3mPzNfOPL
oC+PnhZgiK84AD7+LPsfImXXfK6A1QJpRw9Jv9MBlAlQigRYKB6QmP+O1LcJnORV
VaMNIonoz3dkj693CxAIyd3LdyDW2XW9uLvgrGuz6FJl0s0TWzBG6MrcjFUCURzq
TtxgQ+/THrEwClwLcjtbieerU+mYiQcDM0RfHiieJMjoHw058HK2cNEEVvkht6t2
DnrS1T+ERHQIX39Mau6l3OUmhYmz4W/Pl9XSQlDL6lvof70Uy4CivAuvNawc7zvM
d0Rup+ZfIXc47cETI1ew/C0Uka8o7j9rJfMAXwfKBrSZ/s2pm6qK64L/vytjFwaO
l84Cq1mZ9K1VQZxqff+kpvQWlRgCBFWQvIMKmTwlN4uecAWLHfY36UM+P8nXsend
eZUUgBuSbU+V9vDP8Ifd5Z0TzYZdrc5/9Ey2o/T6t4i+Hi6qJP08abuCc2ieclfZ
PO9k14wmf46pGk+iuuxI+/2diQ5RhATmvOSt61TgRRJgz0JNbTIq5+NFim1nDGur
jmaGP4w9PJdCh5XZ8W5WV5JAYygy1N7hGYamrsAtMG18E0FB6N3brKWMRcNQ8TNu
Cg7tbpRE1UgNvFAR6Cr7c8XGzgL5PtenmqrwEKjsTjyPv4dcgGlHxJuUOD3byYJN
VS8eMVbRn2L4H9lWeGdilGKnsPDwAYDsC0Sr2Y8VZyK1+5ZGhxra2ZH/cp2OY2Ce
OhLWDbYviOr8yu/fVdOPSSyMu5t6I+AET9wjbY9ZdM6R2j0zIa+wvpOYhGWF2Pck
GhSKgkk3+G0ERt5tML6YWP7oep1iwPuLVXRRynqG4WgYnHU3tqSA6yuKv3HHFljF
jgEzGsOk6t4wbYiKpBad/1tU7nWk241h5axT9HRtFchMMSll6FO8CsfMxuJOXEQV
EVyzF2TWW/QMqNf4pVJinE7HcvbEQzfJ4ZGvC9qGL0dJ6W/+t83wK9oRRpnqq3po
m9gA32gBYHlEnLHlK3ZEFJhdAFFUujKGahlDfpI/nojTVo0oC92byL0WkC3TKpy1
jfes3CY2RnVjzmxnU9J56hW9BQK9QPVCSDyTwHjNAovDII5FC3mtjDtNV7akrKD2
2jt7Z/Wq8MeJUItqV0aqJewGttPZOCH9D0FLy7fUetoZ7CMGGYq83+mKmeGCVEdi
nQkuFuU7Bo6oSmxrJBNWP3A4xojykPSf4T9CpFn7XDgVIv7zsLz9D3Hb0uJRKArD
M2EHLNT0YTW4npZf3d5gTCBqsKTbAGUUPorCnGViYisVY1WdS7dBpju3SHkqHkGO
3tezb/B4idaB319w7qWQq5oYJLcKJRavI3pBLhJrekmIob4EqjTZXS0j2AGtxFCc
Pl6rEfRF+M86h3NEu5MN87lFlo9kKxu6F1HOSuw6sgBMttVUq8EACOBUxfJ0TG9d
/qKuMdLG1jQ+YFwxoNFA1L8+3SQyPNbrdwyD02eNCGhQ1guo0o2mDRLxKrzw9w1U
C7GWvNI1AcMrf1No7Wcku8E757yTUZbT71ep9tkTOEObA8ydTJVQQJJ7OKC8Rbh/
ykTqIR73GXIa9OcxVWbFK/oYgt7hw0Tz2vHeDNZ8ZQwdI2O+bcsnSCHfw9gsV97S
RI4+s2AyyWbqyRgr0ihWKyR5q9NB9Tolrujp/lPL3gBH1vykwNtSYBEtYoIwIqLp
VaBgx+6tsHq5lhlTuotWXCwZVSDFLJ7i5THWMUcANZftgF0V69W+Hga6Sulbrhha
FnHkL/UBInxMasq8eKCsN0B+foFwjiNLxHlq4CIr8qXgv0Ge9l1n8Kdmc8lib5YP
/fZ0vppJZA+VZxRLux2KKXz2wnGW6KMxzugBmnlM2H8EQ3yBlswEdXVNNCJuA5uu
CYOSbdMVXsRlAEZX0/HtlDPmdzu5i+w9GdRUk9SyaFHaA8I1syll9qxjzXS5e9bW
+WpAyJzb5ZUHquzXy1YAi2CQWxzoo3tBBNf3JRuNWza1mZBwvWrByUl0OCDLYbOx
92W6osZZgSdlHuTumMlCOYegUBe5rj2NeYzI3UVF7yGNuBQb/8AU27U7b2NtrDbo
6fEmDrHEPMXJ7iHcHYVrrnKjc+hyxdajwh9DMR6kPIdTJ5PepsG11LPZMpr0JWhO
JVCcwVGf0xUpAFrHB4g7wunPrU5Rt2Ay22dNGnm5PJSP/l7sAbSvQEldkHTZ7yjo
SzC+zo29mf7Q6AGnE05BnNINM6k9N8wCsgcFyMpDTX16ga8btIiAeiCl7PSwrRoC
RQn7RMclH5RoVZIoyHO3ePW+ibte/OfZ80S/Q6qdWdjT+DGnWNzstuXKkE9ayDvL
g4YTsuF34EAauZOg1lf+Sz4aDBpw2vytSoquRBvDj0YlUAnbVhxbN9JQz+HKQJUd
AJIfJGe84xsmPaYkFX4YhTo4gM0ggMazawrH/hRk3UPX/UCV7pk7JNFCBn62Pw0z
guU4YuT59znJYCWr6Nc1eD/6p/zfb3Sh3fXUZbiFortB5ZhRBTttIEJaEuGRjkUS
FXCDUPxVK2eGOxK+dZLpGkCq/j3y5PvbW9lVSJ/rnYn2/QqTizEHiBT1mGDjCmXe
IvSUH/yfAe9A5fEJ85ryIPbzBrlv93IAN33OnsrdZdqyeSRAD0hdW8dQW3SlBAPf
p4KkRarwOTu8036xrkyTiIJr6Em/3NTnFykDjuIQvp6t93tufDH6l46cw2If8jv2
ZSdUyQ09S6J1lyKpSESV2HOYcrP4IFWp3VCfP5ngNTV0wgnCWJx4CiPMAIDOykSs
jN1W3JSRfiVpF9pahbIp9F1LNaoJ7I9i+FyZ/dLmI5/gGn2lS6Nv5HrKUtjqOfL6
NWyYEYDY3OvrXvM3UAfsAdwNf6bhqA65+QR8pQoGpA1QfH1QYASHtbwskseG0Wof
7KGL7OZLbgMNLVd2COsllpn58h5uUm4d9R9Xj8sAlwzQ2ynEFBSDAox2rybQZHfX
ZOC03UMQ1X681vk5/RxHgSSSiFugg1YY35nurB8y2h7VlwSo4ktsBdUOO0YCJyVz
itjlHQ8oxi8E4ZvLD1BpM9QuJfy7u39bYcgP8Xg7xBZ3Gsph8BDQXdBBdatGQ4ND
zloSMthnubWNpp76VYlEPeOVaHApoH8VaEfrFL42711IgA5jLVhCgk0waml4kX5r
ao+q7Vnt0Lq7vsK4Y5COg+QOttqbsdkalCJNUnC5NNif2f/2IiXtim24YAIdEFI9
I9dCWpxNugZoO/U1AsCEMqVyeHAv9mabCTiOJGAJvQpF9cX2ZtlUY0wE8CKjFOjQ
t1w9HH1P1TI9THJRakjR1WNg7aa18NAzCWBLQQdVNMVz3c6CRJtbewGlunEAVmeT
JGPtxrofu/hsQ7sUqpPOdMNGte5jlqCBiHcto4DoiFb6DC3tDilbbHvTco/SiO8B
dcjA3KPweijTjWBJM7gvqOdzKL2m2YEp+v/e5f7vRRyWRzK/4gMCl1hdfCdqejg6
CDufsW2qp2xshUts5KVJvGQGFOpEOnAuNPScuV8IL1HkgHu4fMTDErbG/LYsVR/f
RfrwS3ftVQzES8JtNplxWyqNd8TIUYX1K2PhBqZmYnOTCFI6yXhwNNf5KmGn9635
uy2Lk01YqOkfFijGQwwl5tKw4dw50yQG3oZU1PCWOwT4TcQ3wkdwqj8d0YJPFn/+
PY6UwVv6GVf8IT7AllNNwiycy2EerCd7CiqvbkmaIuFqGvK+xMopCzwrlkKVlQn4
W+/VhJDrfrESXx9v5aVL8zEVbIKJpB0bh+e/HscLCqBHmQl1h6+YvqCNdlag9Mrs
Xghr5EKKxyWW26E3kiuHX/wdvu4Xgfwg7vHQ1T3bddKvLOjug20timZqSYma5w9E
GUodpF+wghrU1A+q33WeXlZKOu76z8RCyYc770qunCTePgOk1QwHEchbQgvfCNsG
n1vdK9fpmpuQZjA4EijdjSHzDuiEEmQVY7W1Sv510wIkRnCn1FOv8CfvM6qaL74k
wIUgtWxJqPrpD2SBXN2BkqG6VT0twTsYYJU4u5KVsvJBmOL/L+vUvbNAqD9Cl6bG
G7fDspSIjhqzGHSLPenpABp4qGc01zXPyDFE1zpLSB30lZNBDfn3uI1hlLxXEOFn
OlN5xY5Bt2GLPvnWTQekx1rVf95rW2cwU5aOW7yLPyKKuJp2IyjMAjYD2iHbCfo5
fp61ZZ59edgMbUZ2jcKKX3641Ol2FLhtLUCIujpEiqQagOcAvQTO6ZSQXLhmCcYp
m/Gykg5Z6HnXrsIxypZw/VK5FX3DU/zapHNJhRlYO5DBKn040BjjpUOjY/IQ7fb/
s2trlS51zLCGG+csuEpP0mQOZHlE82AdJPTo8+PGPELjH52aq8/OC/vN0xpF3jed
o4Gk4epvnMaHsFLkyFifeFBXQ2u6VjSC1mD1bew+8lxR+CukjEfLHCgBjSqwwmJC
iDCJfqjznWTfgKbxB+aBWRqA6KSz67sHnNUqZFYpSE/MPEXPk2E6GrQ6HohGUI5g
noMfeIWJZaZzMKytWVJjFwrbPrr39I4MXDjaJhOqfUfNdiPIQYshRU/CR9HwUxl0
1IVckkFw3VVx0mTuqS9LT4Bxg1HPnkR3WmrluO8q5vqu6S50nHZpbKAzsPLQ5QU7
4wAgkVQU3MzpmEL9xVFQkoxB2bgcfuxl4x6qRKAZhkTWSpMXAoRLYxd+ehNe22ew
KuczqGC6GwuhudiBfMZBYkKVdxzLuEID3X2eFMpJ/hfczoWL6Li4JbpRYUtUrAX2
3JQv5BhMSAojuDlmXMaBl8tHnUyTcQKl+E+zpOHOLxG8BT3V+RQDLr+tUXTelHQ1
B2hMA2o6M0PLu2WC5cVf85hHM4w9Zv/7SRf0dFJWWsB0TF3PyO2X/QRiQ2r/lk4K
LhGnGJgWcP51n+phbvLp8836GmX4NxLZBIOtGO++d2bReUoruhIW/Vna+AdngJCG
9b+DB+WletQraEwtT/eHhEKz36bEJg/ZBs0UabSgdlorPeRzktyFmb0xdX/0XgTu
vDLw+LiRI1r0NPd6oOmWZNW5NlPtU3s+znsIuITF/6rKANl34hbQomPtBbFXXtgO
dxkn1l9m9JGG3lfi3Z4UNxzAiOTaQo5dVRJgOrzSSiMlht4dBUrxEHaQASc+CLkC
7sfcQ0GJye29m8sfV/Hmi0z0sFRyazTOzF6DbH0f88mBIHSvnRr8bjZOqgFtdkvQ
Lo7btxomdx2Ux97fbTbOU6JL6vAMlXe7Wcc7LSL9hKvVveoKdJp5zLEe7paImTho
ERwnO5ZW190/ckYaG7qkjsCYyBSaiT2i5JaAOhzsOrKU53HRBtjYaVXJdW0hl5qW
Y4G8KpTwYpCYRHBiN01IcnMhDZCZ5hFdKmdashXukB87ErTFn5UoSMQKzU9dA3cu
uJ4vNH992LWnbSwzyR+R9b6FWcnj41qVC2M8zGKVurl49btq/URVxCNYkdINP9mP
E4C+aYzAo6kOgHT+XXY31Rw1LYUeZIi/rcnfYfhRJPTqji7pcdzG38mZqnJ/g4hL
X1lE2CSEyiorAetx/biXtdu4pItcnon828ESlzzxh6r481YCRdwoQH0fsATtJTAF
mjZS9DEiuzl+qfG5lxedcysPMm4ol+QQXqR8GzdPEP9nyOgIwzZ4dPrrXRfFOpry
XizIniFtO4KMLgCKDIo2zQCMLmt9MvARVVnTGGFkaYXYbyWP+yyLJxqkEUXcLVm9
ZRG+KjHSB7eoMSFKDcywwwSTWSB4LooAZ5++CowYyFn0XrUDXM97Mya5ailgpKKW
8CpwDNobAE5W7dutWN4zC6GrZkIL7lWvwnJNuKmYUKXEqbqtIjT9K/GshphTF20+
zHpLqCboQpiKqYQd+42sWQLAzt+A+fei0lGQ86vmY0yGzGHK5OuJGJTH2uzH4DSy
V7ysyt5rR9WKrqt2zYp7SUVPqmyX4s4D8+9vAMMzvHoxWHbk11vU316l9E3Zjw8F
+bkkcsIqCjNAQTcofMpaTu59yMLHb0f9mxBQpsT4hdFZFZmCXzYpngYjnvvCNVyR
YucYr3k2ah0VbvYJmuIFb2qCUpQn8HKUHxyfbA1f45pH5gTAWNu9LOkmYtHYSKso
c+D3kHG4LrAfhBVfhyZW22rEpirYuXR9z2bHUYi2a80DfPUGPDp16mlLRk6pNJol
2rUhIJr25NbOpsStyEKaFGd853++eNfVv9fwY1W8QMDc46qRK92W3bROh8Uspx6j
eKV3tSNQ1a/pqjv9hFJKEjlqHlENyLj4TOP2sxjYSjHQ5IH8e7hkPuOA327gGYGZ
cWcksMswyGSo8BLU+JvdBM2MCK8xsLtgsvA8Gj/CAIyC25QcYOKAmvZ276TgguGd
GHw4Esc2MNqFHXiRfQ8brjU4yY54GTHZGYxCX1LngxiAtM5bsvn1HLIM4sr94d1d
O1K9fr9Tptq8ld/8pi9DyVbRHHbKkaVOE3zNpMUFRJ6fB0Wk5wM/IzLoAgJRIEvL
OhWOMwR7KDv157rZ7NEFQ6cri3zK3JbUmTv/L5t12JQy854nqVMEG7ApZEhBmesM
cHsp53UsFu7F2uiXDKZ879ZbMl2Z7Q2r6EZVwexKRYiMhJpebwwPxuwThR9YZmJq
NddqOfAnXYJS/O2LSOELcVh9FP8c2oRSTrEsh52oKfrnBd9Yqm4+OHNresz2JTQs
xiYouAqQGVWflwu1ZImWejexHGjngV5TlPumjaaHnduC0u9CpDdKXoMT0HdX6WxM
CV1m65Bl0KVsZdTo4gvYUsfsy1b6yAaMC+vzuDRYkhvCv/K6BFw7R5e0ooYkqa1F
o0NCvw1dsLYlIwhAbwNOiPaT0jyvm06khhvZlyoCrVf0gDF5gFEPOGcDHQY3ILrd
jZi1IfE+HDmPZQWqz9WoAxPWpfMBq0Uxdrt+m7HPWg+1e4+853IQpiuJKwT1L/HV
9YtxN4J9FdA71jKOGnQ5r5kYGDXFCkCBsff2yrK74Bffvh28eYWWNJ/BFhhfijFZ
0B4itZNBmBCSqTOkZUjNSf90ANQrMmU2SwT9tNdlzn3J2okFRunHRNfousHBHMSJ
vhrTM0/mAZOHaHXVQER2G+U4taCAZvjxkoKxOGDUrz5K7mZaYi0bM/ghlY9ZdTCV
zfzeakO6sUmono4wGOpiElwL9A7jGLgqPD+94QJFimGEZIBWbFpg728TO1juv0pc
FxR46T+pX+ZAcUEg26rucO8S7qPJH0rGt8g80ljVc3Nh0fKJoBqGD9d3UtvQvlVH
G6v0vb79LtfKVdMp9/OrEVy7eV1A4ZorcwNY6Sqh8yGN7E7wFzaXEpjkklqEL6gF
7ZOgwjh/JkKoIRrxfobiUmUt9HjJ2rH6bRfSvc7xm/YX50ghKe0DG46koCvsAEmr
+7dlSwrKQ0sZop6xioQa3H96LiYAamAHwghTagjqFxBQM5VD0+RhSMdnJsL/Y/BR
5fhCoTQKMjfcoc6vTZT+yYt2cRV4D/oeXLDanVzKb8izVrzF+b/5cl+bpRpMABua
6fGBClN4w2PMa6AFiYfCWqU6AgI1/ZjWllk54rYsgRRzKnV2FLEir+Go3a17CjWZ
fvqpLgjvUo8kfgCVKSvI6U+PO5WxisF5dVwWRJGtzv7QISZOHvw4El3TjGFiWt5I
X5rSZLhvTjHgypWaY66jC20EnkTLuRLyOHU4thKDAzTcbnOpYU7FHk8+hnYcWm93
zZOshi9TGbFwU6P26BPxV9fCUXXPXT91F7ttp5SS9lGJj1dlar3yk1hbXS93Z3iA
hagx6wdgKbwApvZv42OveDCku5lH3dHltd+lylzB7d/LA2IElVw652luHeKBW/BZ
I7wo7jNwV1Jnum8462sj3moWhCRd6Sep+nLxhS64oFZRFaStiyBIq6xmEOQWm80P
h0hiYJX1hEEoHg3Xofbeim1rAEERic/hh3uaDVUjGaEnWLb/Kpei7e/PbmX0dAQD
ZOw130usteXSfqkYuWhY8FoEeXC2+BP32qnkLdKBV3bnjiwhNnZb80Uv7u8Y1MNv
iwHPnq98B6AhDrNkdL5EQlutJJcIObpZBPUnz/82qif0emuYCBuShwVmr+nhvc3/
yMMQC+aQUenT7HBwsEWrZEPkNqbHTPCcg4JwwejzrqFwm1bniOPxsEKe18Xrld4D
kfd67MdIxNLXlrxzqm7JMEs+xPdVa5m8lSWPabq2CP9XeddVYF9SkQLv1SPF6uF0
aRJflIafmDuSmKrDfo1z+cVCsnzCFbrgOccOgFDDef9YiNUNRDcAtMNsl0wKo+xx
Z89+7zRoVLSPu6llr0CnyGeEySftZphKee8etctUF0srpfSIpkW34EjzcEkxDRjw
70QhpW9f3Ce/GF3VmEjPG76M/rBu7ok59UzyE4N8GBBkQY5xzyHDAPu6pCp/FRhY
1+xvQqtb9abxrgl+GmQGzihbL/Q4+pzKK6UqwJC2IvMUF+sZB+JQi82jOBXKSdt9
qp3/+QzKD/9rfJKU2idGVjY1+4dqQuJ9Y8tZ0PMWmjhztOmCTKFkoC7dynwoOadA
6vRlH796IXk/Fk0SzWs2fqwwWpEXwPOPW5YUzoXsJ7RvfXXD1E3ADweCgKJ+/oJo
AJtxaAWCHzoUTR/6DD+ngaArL4oWLX3j2121co13+H46/qEFOk/eGCzoABTSQ1OG
cw0xcDsTk6zNa6o4o7re7msfg3dg5xxVtX3s3qO8hEWZnZ+NP5P1XwkYw/FkZnvM
pf/UyqDTU7zW9XbqyFaBd9S3zuAT+7VMvV+CG/UnJP8zSItcHgyVDeRyhhJ2II8N
LSH+ghf0fn56QOKJbuBWe7sWZj4WhmzrKWj4JTp2Uf6nUHYdtWxGG73F0Qw+0E+D
IzOZnHGgjXbLry83xYQIbAYv02GtbG8dnwSlfIClDrcNFGM/ytpkGs42wer6QVSV
g4rxTSVQTktt2cdh7b8lxFpwCyy2b49v1LZYS7e+qL9Lfn7QGc/xZzpvb+TfU7Vk
1ynG6y7ebTSEx8azNpV3v/chc1IvTaQDUpGJuc+NdO2Vt7d8aAVXfsqZfGUNWUg/
ABQSKoyJs3z85RqJmzbF1vYv5jekMN4UQkZVvKL6pzf0zdcn3BMAinDIH8LqXbZ1
dCYXIAcPki6sLq2GWnKLRfHTc0ihfwqFzdgpvQEYV3+TlXepBb8PcBQ/py1XR6Wx
gcoTDrVIdqIBm5VIMdap6xr5mNHAgHK+10m5qGQcXZ/7tiaS7cSgc5rJTHFs+Jkm
YnAwPN6NkcXrAgr4m8IDVS6AxnLnanxi1ZH5YzHGs2+Ll6QlqVGRI57i3QURwPrM
qhgE3hKGFWFRV8ghH+SmPhXANWtjRfzR1ZMP9JgPyxentwMSH/dLo6PhGrROsh90
3rtm4cb3epzG/kBU82j0SoCKPsl2jIqyvVHmZFLASVFGGh0y4PudU6x9cgUgc4xm
ztIpInckDCl/738t4werqDXI//zr03IB1wk3Yt3DSZP60m4ILeQlbWyKsOniTn6F
jHaGpGUQxi3Z1y7DP1yur4ydFQcPRBLoEXY07ix4NC5gZ0DcG9ydcFTRW5KTERPd
7+8lG0oLwIBwBIJ+5UV9GNFhLlcRH18ovE2r2GFMKX0CyTnb1IiqgWCuKQPcy3F+
EpiEaBi8MWcBWDy8lGYfPwLIHER2X3i+EY1m/CCeBsmrrQEC6G2BERHf53TAL0Qr
VhIX0jYRAtGfsamUQA/Iw2Y8+eqiqxsqB0Rucuf+hjbwMSqpI6A/Nkm40hiQQOW/
F9JpGd+BRtqrREF/Acrx5H4XK7sQ3H2WzAek7LvLslHtQbMRH5h7ZKqN8S/GSMlc
IomYUE8riBVgzI7xgsciPo5PK1u6a+tcjcg/I2mRDjdhp9BRghdfIS2NhmusZf7i
lAYQnA7+YHk0oloCH5uBIEqT7i8MnaN/Kp2PuGidyFi+fXlNVpoBgI6LpLf7h7xA
q+74jqhX4omTnyAdoIYrRNAH2X2kpHqmqfDHlnVaoC1JUFTM0IRYGOc8icIQTjKR
qqVSs7kEWDGU4mn+OA6+aUyrzxy4/9WSDKWveo8JLy3wx07VP8GE9YrX+RVYhhnL
Qvp1A2BAmsLwD4CrGKH4Sjl9HEj/BavzJreaT8MWS71XFsqYmDAQZ/eKkjXlK01I
kAegyOOF05l4ZZNyAIjozoCxwGW1CpFippWOCOHYU0jadnDGuRAlQ3VRs6inYWxM
FfSyuXxN/2MRe4HhIdZoIva19pI0Ck/lamp95gSIHBBtfecNjnE9M0lsVpmiaagb
56PVb54s9vJR6AM9RIfsgl8vCTbrR37CssYUop2ljHau8iYdCkFp3Q32fnsA8+ho
kKSc4lqTyrIXhJU88K2ySLMtFeosUvofCLAJVwH0yqBMAt+KeghS3ng+lNgUNUMJ
GZm3HYChgxhrHsORHvWGxUsjysBdNoCa/ToPmVCxU4W0fqDLb0eF7CaaCHlgSpDK
lccVEWqFZt1CSmwIDqpZpqlPTBPlENWAofQphydh+J63mkjFYApDmcQufGV7tcRS
MLwU7sxA+SS7ykimEq3INd324F/m9ym6oA7nSrD5WaXv5eDHtSlq9eH1Q82abtAz
DZD0QozvUDw5ZOeKNHlOaRZRRr96vsF/6rnJ39uYX98kU8gF0/HP3Y8cpOL7q7Ss
XkZz7Z7ucI9EfxkVNEJvZU8uvG45M5VGJOGXL+8mKftP4MJItYGHrU2Vf1oMGIrD
VdtgOpUm+WGYuD288qTgdNykardGco+LUriU+cpbZIATGbguulGVkWB2ZBfJfq/a
SNvDbmCuoNVT6uV2t7uMAfJ7Q483WoYgn8GPmzCSxdo0O5Ycyt06149QrP7ycVXJ
e/ZepYV0KfNagz3lWiV3GySPsskskHJmnaWN2xw1UV/s1ULq0DJkD7aTNv+O8/+2
BDPxs1YiG2u1n55VIeU5qL+2bm0+Fi6xqgOD/WK7y2UIThvesSLq7pMgyOMDP1/O
QWdcYcUabapb+wknWpljLmbW60wlpYer1caJxwqdXk6Jfn+oxRicqp1vc5Ciz0g3
lhG/mgJJtUdvY2VhwBe/Ey9RHqCyl3jmT8tKjav2X03iLY/kJ+IciJXDas4vQJiB
kTWLs7QRCy0ix2LqYrwe6lW9wa+h2KKyYqFmGXIoYbgZXTMhKPVeRi5tuEUUyHss
A4tIQrLQcY0WyHPz4h1TKQtQIEZUPvhoMFpsPn7sEkIeKME88tPdwmuZOZa2Pvwf
s4LAoMZ61PC97W2TPhwHp58fEMv9DWpv6XMHmbYozW3ccBHbFOGqFwH4Myz3b00R
V5HvFksaXaSYd+s/kvbsdcB5QNc3t6o+fNHi+QaVtUUhrfe/Wun3RnjR5ZAoSVIL
qWqwa1tqOeQ4893rGNZ/5yMz4WuZbVbJOfPfaRv3VmEoj3FXYpJyhbLf5AxRbTfF
rqcINLOoCIy0R7e0zStRylMHAG4fuajxBvH7WSVAaCxzkCVOqAi4S9aCJyaHtRfa
lKUFK+d28AjWdRQBcBkDgwqjDj4GZ3Ge/nHuoavFOQvFuGh07Geo3wevyP3wKW24
0/cMXT2YcVt7VDKYFndmJmnGme1c7Pl5wPj/mZpnd/62QHAfxelXpljnoOE0Yybb
h8M89afVuwTuYBimClmH+roHekH+8xLH3q7Xk4iKCz5FwK51z1DlYWizoco7MIz7
hZAqxDLjcQg59ActgZW0VeKyQ/MD6R72ur3WIQLDRecOzgKJaFZuxtZwEPHYNodu
NQKT3zpZWJwrQXw34+0AwCD2FzeBgC1xUg89/2z+15Xf/Q2fwgHImRxJCOsQdP6v
2wIKUStcqlIcyxMmR95WoQWZZLa7lMROLxQAXdsR7ynV9EDcqHjVd56vzMMrWlTF
r6X49idkpPwdFinymHdIGpXjBlnsb2Xjk4ELsNv6zOQPrW72J448lNeRVOUcOY/a
Y3p7E04DP2UemIDpg/G5C042gyOmttT4YihRyBJmuUB7zVhbl7RI9d5T7FCZ5pZ+
aHdWt1rREayY2DA4sbXv4zWZ1Svdm0LoGUMJ2Dax24ouxtDpaQjQGX6Hkhy9rxZ/
K+1it8c3fr5Z8jJwqpIRYmC0Et0Ncp9JNkCjkAP8uXG9QWXy+yccDVSmtDE2/ZKe
Qb54VetIEhP5ZQ71O4yva2oxO9zPRXkCkCpuwcH/DKb249yBePmhUa6VIxI88/G7
RN/XhOVfVAu9xMxYHWt+Jt+yWa4AuNLNIUvv2uiMlDrCFOsCQ+klZnzUfGN3OjAQ
pSQyc5sBmKxkJMFTMC6YCH1dmZ49skFr1c20fhaRGj8xSDj/ivzyV/MLF7iadnD6
qtjqfKJiZYCo5Nv6FLZelVnp/P9lu05sYPzXZcywCA/KC+FBZDaPOBu6n8wwi1wY
hCrLaMFzovHO6l1aNzQCwVNXRCTp7oNHcExOImy7JDwRtTuYv65Ym2t3STQbGOxa
5997QGhvJGiRwdQxoKl0mPUdzvkxhNsdCDJniqXhga1UOZEJenO1sQH+qpOLcEJ2
cxre0sp4rOWcPVAUuGFrbi1eKltV8pOsqvp873rwoh7pDcdswz+h0xF9A0cgpAXc
APiKvUdwzeJWgmqgX8bGr3o4hXwIsC29gDDazIN/DKidZSIHGzdp11wysJUusHy8
xt244vJs1xZ8o8od1Xq2qB4DBC6JqGcWsj/vQ+CQNT3a92NBwJCj7RYt3aRjioLb
S+zpIYIxQtflU6RnxPi7N7dgo3BWiNHs8qnR5x5MrH5fFqA01zNBO8hovf+Rc91w
S1gwQQoJ61Zl0sDZ/jHM3CqrF20dGXI+ddkrzTPObDi5cXxjUnlcbkVP+87Y2b8F
wQ+649eKkBQDIXqa3Y5jdISUW0zAR3UBI8LMGyStjM0Fyrz66XlLJ2Dto+GsZNyK
zty+3c4qpeDUFFL4AEDdITz9W0fHQQN6zISTFxRgce7L1MrIgZPLfYzYbx3u94ak
acpAMpWn9GgCPvQBu3C+JmRRe55BUXAqaCVCWmLQJTN9+yIe7yG/HoBehP5SqyFv
hN8yQIRQJqIIz2KV/UvXOip/rvWWEMo9jV3K4EWOSeSjL83wS8eoyhBbVHuakxD/
krNC5Tx7egmYpD2Ukbz1ryJ4G2A0J+uxwG4N691sy3z2bvsafLaWdc+4BVy2e+tV
cZb72P2eJJnTA2ApdHBevl7Zfz2I9q/ex2xmaq7Zo0edQL8C5Sb6x9uR6A4qqa47
uBXEIerpj8T2YeGuhTn4yXIZXQLpD0Wq25ccp/lFY5IweIM9jikN07yLB45ugfbj
wRd652XtTMuAm514VIw9NWkowmq+3VT7Y+Na5x/eM9mjEzuhLi98GG7IpbKOCnEw
qLeHbb+rJfxerMXb2WBDGgABckYrDw3/ZhHwosVgigIoLTtMRTixNGcLx9m7lpB2
Jk0mptVK8E0IIf0dnRJlQ3rwiKFKJXhDmU46CfW/CgSCpMLfO6MCfT6Vr3BTYNy8
6MLALznG7rvBWueOVJ2h9uVptuKd4adEAAw3R8gJKTL+oGdVi5S/jWgq8rPNaRCE
U2J+/CUB/S+JFhI+SCqs4KFv4aF+cKmNx4TycAruVSJO57d25WHdWgfY6Bc9F4SC
JPMr1q8MaCuFYA83qWfhqTyVsAkqI8lmrxDGWLNdHr303TNbYFb0HQvMIQUcCJfw
7lvlGIRDzdHK57lBwAhdULx7JDnLYXPA8SBdn4p8oB6vLFGLLs2eAjXUPEklQ+E8
DVRwA9d+KjmYkOaQOpgrnzCU0eWznPCcMgOA/K5xvokF5fWLMRHjlE+5/w06G0+Z
MUFpIHIhBpXO/R15Or76qgn79Rl9Bq+bnrmPT0zsEYZQaocRkei+Z2dQA/pgVitT
KtkXZw9JLJ/6Qgcm8663bzep/bsDw6eaER3v5W1dOIYY5VTqhvGhelivja3P0Cdf
iaiQx5lhNWy5x9/p6GOejQZE9v54rsgcEsreH3DvzolevH3FzYZM9/uyDXwHtCfN
cqY4kqtyqYglyFw7I4dY0etQEbyXeqiOltmW1+EwExbMOproDyA+LDkYbcNJtsfz
4q0JNX/hssyNNAI/e5frfIc87U00nSNNpamMiavr5jARHeBlLykE6NCG9QFo1mXo
idbUKfXQT2phQsLLfP37dU0I6BR6l/pR7ReO2ucU7Y9/J6sqPAo8DOBDEW15t5I0
oSK93ByzENAxHf0T4IM5jl7VV25rIlsbuEKmN+Sxw5VgBLmmXywoNEa2Qf+FVuXa
Zziyp3M0CKaJ+xau4L0fgO1fUPQHoWuGc7h/LqTaj0dOMvjVf49CjVmwWMtmmBNE
/RRhqVZBGp8YeJCWGJHEcNCVgSs1uSJpkK7z1JLSTG7jqoiF7oZ8jRkXNnRCQcw7
H1ALnsdh+7KpnxyqZiEjH5PVEFjYVG+3l//nEvFeNiHL+AKHQhzBXE8kC/czv90L
tSUTfxmrsZBw5DCHMzPdLUyoG2KjGHr3oaqjKJiQbyJwWG9TPgYOhO/m08h2Y1da
pWOMnYzTA4Sl111/E03kfnA+zfFhOCi1Hl19ZMma0Y9OXUglMNYwtPkUuuSSMk05
jN+dFamuCWpN7xfEJJq12dlyqZHTaYh/EOi620FxYYFAoJzkniZ/p5DHkyxIkC+p
JcAJMv4A50mNB9OAHopT16ZkJEtLCGfwZ101fRTzzsF6c37YdfqkVpbiiTEAH32d
GlrODwly3rw+y50Hs66fanLget7grOUbBnUVI9sfUijk1lNf8HK4in6C/ii73/sO
WARNxLeFu1JdIl7D20oOt/hxpyXj2MeIGUUJrhTrkwFP5Dtya59Q2C9v2qVy4He+
KXtXvbVM2ppvNcG/CIJWuaCqPvGqcI5DfC6s6MnlSgTEtErSXrkIMG89m1vGHXye
tSbgyCd05oc/cCW8Fb92GhDx7yGcThUtmENyW8kIlHwnwhiAcYIm5tY/cWZoOP1Y
HwiYNkfnRjFqYkbHaAUOs3xqDicwDKAriOO/UWTTm56k6buC2oFkUrYU1Ax+qw8J
Q4XB6ditDzBImpxwugCGuo8459wGGbXkMoAjsEOhkvpyXHUPXNkVTwUcaSgh+Pqe
Hmlx+BPkmHdjvw04UvVfp83pLYG7ppwFg82pVScsitWtbNlvfkIdET+KKCXDDM+S
VFhN6Pb92yTHXzC8ddMxez2Wx2Be9++u9+If+thm3sTZLwqeLsCpbRbNr+Kw7UrT
dH4MxSqiB3wXdnHKJBTP1Ekhg2Id2q8NZGp9S9I9Q9rniGGIv6XBQ1T+UTFylHmU
Cw0SWdWaW+RNGq3TljMM/MJorr2rMGemHxxumYKk9U3DjN6r/wJFwWewRhZ2jFVc
yR0QKYw1rYP/AYYHFBxmOeFCRb/EmB7xleGsxW+NTvOPkzCw0P494i17TW28e5le
dNMHI4lg6qK1r28+UtEMBk2cgb13fUXP2L2+lzvW2xl5uH/4jcpJ/01dImLtsGsR
J5qWoOX/1R/+7mtHdqbnIKaZDvGOYDOEm72pnH/mSyDJyJ/STbY7N03quA0ICrwL
QZ664x8lZiWfNL/an35BrUjWxhHLtkGGfIiFJPq1EV6ZKQO99b8FnDQTcZA/2m0T
qh/3Uq0fcmrt1eljBAbwEwjqHx+MgRC0QR5ecG5Qxk9kSMvrcHicYmrj6EY8V63k
xZCWbtZ4ouP7TDKpz9FB+tLbMKZ1MTgdFXpWjxxCn6zlDUA/WvnlOeTG2mb7H9Bz
Mlt8yYKYLq2JbK/qI2Q1MOdl8c1Z709PE9pSbcq6yX6GAxTA+TwaOMSwvq+TKg6z
w4dN2mP2diRtQBD6UWjyCLo99EIDKJymmYF7GLy5xl5DyQeNFuPOFpcHqGptpeDC
eTAXaT3u0N1ujgYnNIfZqwVeGEkzTuPHhbrfCl1oQL3/m1YJ623YrKYbojuOBqbR
JHzDahSKCkjOZSpGL1hqiYCqJ6tKk4X0SsPuFlGVxu2dx7SiB3qmW80uPG/4iLBN
oNc8Mi5pX7tu8No9NcAvzeB4G7qeB3kczonl2+qeMHshzrauWAAAJJuN/0b+doWY
0qqmg0t78MINUjkC9B50nfTEkG6YSsqWnpuXLpGc3rbNpvYElGbMBVAFFf8x4bk4
tISd6qMA700EcVl0X9iVLCWNjE5l8rgMi7/a4FDaF2PkOYbNt5zAJ7sOxD9cfmi7
MDN0xsB6nQezHKDUj/rgzzx+dpNcsdIa4OAldEx6vbdhwxhejQZ62pWlwbc6g5nW
Ro0uFjprs/atDSkwHy04OoCurrW28C8dzKXWxGpH4Y2unAUs7gmRTIEWk9fTAFqK
0fZfXuIIzspdph5dynQy6Gj1dBkcn8aLUkoLMPeHKQ8dmvy3J29wGPAjcyi0/ISZ
WN3b7ISk8iZynf+YdYUdWMnF+75ZIs/NpoBALhDpqWPHgEfv/00vlA8RigIuHDQb
c3chtVfHSISv9blCGBtQTKwXrBspgb9xZAyq2UXvwBRiGgIAZn36K7B4SLC5Uf1T
1RpqnRR20+lGL9/fEn/rAzh2ui0CRR6XOpzjvlauFafaruvUTfYkWtH2SI3nCF8w
mHJY7ov7A15h9+FAhsHxZmjM1syV1Iph+b2GztiF/lXf1KkwcjoY/tHblbA2OMl2
OOAW/35wew3lKe25sOFkrHRsqyk7nieCb/+4id7UbZb3LhV8mT67F5zMnAU4zJzS
yMKPtF4lh3B0j+CQ1yqIqwmZ/Wh7nRoAlqcM/diFvTZYcg8AryQ2kRxBzoHWCY+L
38Jki7/mjGTFmW9tA+t+PJ+U1ufWiZNhLAQTrV1MTL79Yq7UWNOZ7SnmM1v5mbK3
DAFojflIwzENig1eBTeR7kuD4h2LTgIhMjRyHQR6jGfSztRjlt3cA/cZeuNyRgM+
fybNI+HRB1k3FPMKsjk1mbWR+nMKSBNfEYIYIbbIVX4Eaxlwbl7JjWNdY6pSIy9f
ITi9f1rIj4cHcqlnexIcw3A/0z/2m6RHpccC3arVpNaUbLDPbCkSXWKfntAVN8I8
sOR+gqephg2co6zEopTxIh0ypewlXW2pdsebzd9bWi/S+iYYMyamolRWkSazeWMi
ePneTCQy9KetqXWMeCXMCVy/Se0jnk7TpvQnZ8st9x7Zk1K4m6Yi1M8Yrc/U8uAG
ClbV63mn1LfQpjqifQQTdt7UDXAZfcLvrCQ+U11O+d27uP3aoO+SYmNFQjmku8KM
KHAa5mBkSabcH7CRMdd48BTt5BAa3RoB1QWDKvUmOfEPPIJH39Q0lcs/KpqwJldB
c/qzpgU8RpJBPMQncsWjE57dw3CmOmr9+DRYs5+0DiiPEaF3gHQFW4o+lpDZpdiB
KCQlR3uQwWtZPmUer7wqYubR1TlEG+t/GDfszDz+9whNrAWhlCWZO4CFyO09Gyjg
Co3q5k8FJveDKtguklm/i1kTWZ9aEisKfKuc9zRGMg537mGsvRzIB5/iorZuZ9RM
RfSZ/KmN3V6bCvH/+zRNf/bfVHOX5Zc6VCtfsG2vWWFyoGOeP6t14afYOP0YzXJl
a7P4depx+iT4M4b9SN8GKotnUfyNMyfqAMK1Qwzjt3R6SAkuc0tttv3kFmGxhEeD
/SzuMUReU4gxHA4wsD+DNqvJC38o+zZ/pWZLfxSiFmIiIvMPXiqxX3tPzDJT5RBg
O9sQTcR0qTI/oNZAHIGNQ43E0v6W9PMX2KFxBP7nkcejGu1Z6cNtGR4WXzDJvZ2Y
JeSVkXLEsp2/fPosKdAvYcPVVT2+9wRGsvzjzdzX/yWrU086ii4Aj9AIEbRESwEZ
3RmSLdQridw8quEILl/FbIOLpM1ox+OwS00LWUqKnEp7LpuL4selBocXvuwZ3Glw
cLUvVOiKukQFEH1DFMgAEzIbSQRg8RVTZHpJK0sNL5265s2K0a75ayoZjoHXUuHA
MfhLbPg+ZxaAzzAocA4UB5KBebckk+G1r9wgoIcIR17+8udbIi60Gh8NKwAMk5yJ
mXRWntGSzbFsRdNMz6HckCFEz0GhZJmyFWYtCt08zkOONO/PaD9ae2EWA7Jo8xXv
m45Xic05DsofdOsyJfi4+C6G6KBMfTOPZD+yUa7d8sCauRMx90XrTw09DKRG8BIY
mVbudFKszZSrqJyNinKyXj97sO/tzGyowowK4pk14rV/HTUe4oB/6xiq52X8Z7Tn
hJij3l0pngO5hKhb3Wci7aBokwnQr33djoqDP35q0xEdqshwwR5ZLqmJXfgoD2Sq
gjczIwGgWHrSK7K5pirl32FmlZrkRxOsNF+EcaeiV9pVIuBDt0z5lWxUbYqnUyxz
uv73GkHK86gmfLYVWoLBjre0Jk0Gyl/zhf0+WIgcozk5+wVo/RBe4x8paoTms/ca
FOdfEo/niW64B4lmtq9XkxOIiijXOgMTfrILITaOdC4LJ55F2chkzwarA50F0td1
PLO2iZ+G0bb9L/e9kGZQcDZwSrygFSUCUUqRBupIXVJFDuAPVC3PKGsTJjk4akLY
AAZuyFQo4CwBF1BMPl421aW0OCaqQ+/S4yoeXbhYuYjh4XLAhW6/Bgem9el8G/t8
DU/ncwKK091B522/gGUCUUx2qNY8NnN41uW5e5F7NvxYp4Gt04aybgqtjUa2p0/D
HQaW4hzbuGuERz9eTo5j9oGBh3kEr2V8RvX6sQ/+fbsOKizgLDNZumWArrjGR8wU
Gp5BnqLED8zPspgZ7lV+U36aIcn3RTsbyc3CCwRcstWiERF4U2FXRkAzj4jCfSGr
w2tnXPllI7HvZWLp423Sj0drw5UkBS9Oif9srlN+e0qQ0M6R9BV5MFAXa8Hhfih6
4yde6r7C3XQxYTFP4forTam9g+qCRlJuyW5V9VcBDXPWEoghC4WY51rUrpJq2Py8
942Ln0CeC4rJPwNtZVf2Y7wOrWR19jyTaSfIQxbiHvMdxfVr9nMy9IufGmO8TSwN
aQZU3h512EUFfx/6yv/tQPAsRLUGblu2qNJlw6wEoRri5Raa1n2YUdzmRKoR93WT
ISlqwa6fNb2JMC0SNvW+/9lEBEL7OgID+NgCibQNw5pjrGJpowOZyp3W19XDz8Ml
XmC6d0kLHzD+B0GHHVtx66+9yySqqLUZt91OW341WRZH0nTc/HJNP5uetDE5QgZf
uqAViEefmaMkdiJt6/kWlZV4c43FZIVp7CZ1oBvESa8KwdilpuPtfyYpE6/V96ny
8gezWez5m/DcNMG1BoOd1seaeY7swZ1K0SQq+X6vBDGE/r/UI8BoTc2kePbLfsTP
mpkjeiIHsX2YS8u5RQDabLVu0qIDC42RnJwnFidGYydP9aV6heVcBb+yGKzudPZ8
JKzLe9zaiQK3jsGRYaoJDcPDdg9F6GC+LgdKPtD3q3ZFRLehgD9sdXkl9OsnqtU0
+b43tx1AfmFwgwK7GS+GDvM7y4Zcv8qvhvRyXijwYpHE1b8wdwwQYgpa+PJZD7X5
ilnKm1M8SncF04np4BpQYT3hOMiMleGs4+WaWLztJ4wkrC5qPaZexW48rBlQHCX+
gbKNLOrC3NO2zXAtOnZIp9yaJSooXdxCrC1WARclZRiZOF1gKbSqZfWndo19peiU
IsrRsmcu1eRMRyuF0K1qlsIWgBTXfyhA6PjFjVIp27cKOO+vQVah1ZqBSUQz9npR
W8mxzDvASEWYnsaRKJT1od/xKQntOg5ArYa5wdHb75LfFZAkiGeOohyR3J6oPsoT
lk8IhYqB0pzzUTCuhXqDl3vNKTZumciOlZKJd+eTizMQlV6V9r8i26/2Yf0uhRIQ
s1gyff9EYe4NuV5olZiXmH4mFT36tPrze4WPfcmrzI4Gu713Sh7iIPjP4v9RvvP0
8fnECAs95cJR9O8t4J8hqpH5qUB2jj4+F9+X3ZU8sORUCpMTbZTW/UNM3lPeEvfS
C1QjSiaYdztc3pnGpNwRZVgwJT134BPP6U0IF0ndOuVfgdOndM4hkChQRJ0bd09X
wgxQs1dDJuVGI+oNhvAliImHN4DiGRuP8+u8TQMJ4ohiiAOBbDnS9C4Ja41uHfO6
CmUdj11Fuvdw0dhgurzydPrplGQjv4xruW5ADHHIqyCpe2yDgMp9E0i4alZ0KTkG
qme/glwUKftBMiZSOwqkwPzrTMPG2hIuHNW2Sr6MsfafxERCzylQD7hqI2cB8QiU
wLzU9i6hYBqs7h7NOsAn1l1vnABxO00ON+c44CHAK+k/sYs7pC4S83R4d3snqkF2
MFj2iuQM9YojFHNbRMiEIceAUl6E7moLl98BdXEeTejzlWse4gEU8Z4knvA9CxyS
edeTeTCYQc1a/mO8kXHYXfwaWnY/32QzIRGkZwwg+mTbAShlDlhtZd8r9woElduh
dBvapQ9h6H4SW9ImodDEZe7uUykEaojgqD34owuv24ria9CM0ypXrMmeJ3L/0+2F
HT1bD9o5PGmFHgqltuu/3chWaVJMzU/QLGr3vZLH6Ue2otBTAxW6TgDDWUznEn5b
SWEvKZDUh3eWIKrHe0qZIUCqCyd6MVAJhM6mxvE2EzW7ZqjHTbuDwq72hZTaWJGG
359Hc7SGqTZgS/4dDXD3p492vOuBf7L0Ih9l1zepNxWJWlj2gnU28RZ+XM1pLNsr
AhMuoeE8ZWVn3CDuEF9WErPn0Q7Vnz1yRoRmNAX2IY9GPWr6bIWSbh3dQbGA2yrt
HHnVg4DtGD33BALkLEWIc8w1ZIPC0HuYfzSVxLD5pp6mzpDwBgqE5F/ig87uvXri
ZTN/0vipTg0jEW4rmNWQe9BUVx6xMOT2uvUC32eaF7+SBZG+qzrAGx1CTqjAuBA4
dXucroc0hVTLsIuQZFfXUiLYXdsEHdKez22rgc4NKhHpMEs0mnHu2anjrQ5FDg8o
z/OJaClcteVUDgyFt13NWs0bAw9j/ml23v3+IRjGNojgM61FJ7dKnY1D5yzOPoSr
oSTwyMIv9U3JuSUVGmchVerF2arSJmemoSyU22Pzp82Z3Rdj1dDUmBHs+sA4J+Ch
azsMXr3khuXvw7SYEEvVPX8Y8QOmBCqExKd0EHdnvHpRi4F3lQ645WhMo+B35wYS
wzqyLbQa31n4buJWDzKgC7LxnIun+6EJ1IPnq1nP60MLj3O/8Idqg/6yKURg1Ykz
8Kz7YhlKKzrRpErygLWqpbZ77+UJGkzdU0dnhwLc1Tjw6bFU2AvxoQ1GYgmhAmMq
TcoEbm67ZboQ8yVJ7ODmPqDySwciiapxvNpCV1qwkJa13t7wBuQrtS47XGLiOe7R
YZp5EVp3PKNFbmqYdO/UTUgRUkOPyhfmgzw+vD52GarshXX1Z6WBIhzD7quXe1wn
yeHEp2UWZVxI5PWnDYs+UPTngC6nHzY8d3i+ONMdO58ItQBpwEDBkQMXsFgj1201
2VOJVpJ3/nFdm2LKLDdOgF84vOX4ncYF/n2Ps8zGJ5CMF/XEGRl6+dfQWrIJLZzB
k4pxEqw5a/QDYdwVs42fPAVtpkTsRYxkkgB7Hnzjhw6cYFsumsZb47pQCkIgDwEq
2VNa1iPKAQpGn2xJRO2ZhV6p77OjzMOB2E0JY5IAQCK6olIdSClqcOAEHuJmRone
bQ5Jwo4OcnvcTG9EXuBxA59ZVaWq8xOhCZeS/Qb8TPdQYWz1iURkPLEq5IITy3vz
2b9vZwMgzNF7gEc29MrtlVf8GKOPUneTUmGmlG/hSCLnfLVxJt/xX3xb3Kbam45g
rpUCHg5Lwi6I1DUGhvk5LLd1hnNhoDzrw801iWywnVONlyAm75hS31S+eBRWcnkS
41Rn9iV5SHsCf1UZmupSTP7SRAXi9WvSyBdOBBHksl2iAxB4fhBEuMejmydtt2c/
7gQFBb+LzAyiewHE1LA/LfJLVxFEUl19qHCAqpHdii8uHR31JrA3Az1eVaSm3ifY
ljm01zzQSo2f6Vc9YrsuxbuOkFMDq1FjyWtSxXzahetgeuSCGTsDpLd6rJyet4LT
G+53eIj2h173DVNoVwNZdEl9IG1CRM12ce0Lxxeep+h+gq9BO+C0z/yz0PhwVKxM
3M8xSW96+fachyPje5p4kPgJhDQWCEgp/aN0a0Fv/JNBAbuyTO7e3GXsr7PRC+WK
HGGjyHgG8mXPquFGY9KgHBhQLoUiuX9tpJJGpVtKEriJLvq7XZJXmy5UMNZuXsto
n0i8Uj3Gg2wSGBPJVYI9gH5rw2iCWtbwF9l/lQA8Y9gc8yxAE/8A0VI8ivRYZ86b
cQdmfD0aGfjwCku23q9WmOMcabffX0gS2ZTA+bcLaibzz68TdAIoBk/HX7IITrDj
gnwjTWae3ezqZRNyHrzOpWAISPFRkKd4WzlSD7yswVXmlGuX1prEMtybQBn7/kXn
Y+eRfjOr0R7jRjRZy8MfOTVwtkUrJCsxykXP+gGZEXbaLxFQG6zOAm1xUy7lqN4J
e8ywIkcQV10utQpFQvFUkCAcml5slLA9bZyyeHo11ZVAXrrCeqK2CgEOtzwDXvpE
iFH94vwAoUgGXccas3DOob7SbtDM8XoubvPa9B8qeML6Ip0uAr4Pl96AIqi8jkY6
GtML38MF30YO4OxeX7tFYDh0yCyvq5NxRdikg5rYRYvNrp2RnV0BoHxJW/oBQLe7
kIbnePlP+1VS7nYUV58lavcjm1GogSc0fMO10lyEb/p6zlPCepG4QbxJ1yo6T5/G
gwfrXhSAurHRQYNyRfjihok5jmffzxwa5T2PHB/ZTJfPYKeWBi/sLpdbhUX89P4r
RPIsZQmtSs+3icp2bxhZ9C0VgC3AX/y/KeOLlz+Va6kvHOIcNvjH1EoJHMUitIiM
IaWXRHeBeqt/1IZ5zKnnjLiKG3LtcKeaigYRbLfkyLFnyaj+rgYK2uuRbkXCKqn9
/X4ec2fQFYK5upQXndOS3yJ7VnUQd31uILf0qPyYlYfeVY9zCE1kCNQozirSVxYC
HOX4eXyB5tLcHjBv6DKuPVbw0GmGglJ7vcCORcArYM9v1fQ4+RHZKQ3XCiKVf2uI
fstOOlWr1HxxoIMtJcmsSAP4t3cmgfRsq6/JngqW4dHacHQ1qFBpKaemH/iPNlgQ
3BaVJYby0s1BwQIRvG7yJVUz2dOlRky7fbSLVsK8YLSRz0lVndDK/8eVjm0kffQ2
Ll9yt9wQ1psBM/luxFVvU+LdBKy3KQUFhUb0mY5I+SDAw96a0mRI/Mjtl7NvtkIU
58sOWe8X6N+io4BeDlbVuTz6T5qE7JW2MogVur/B5NgPTqjNiE+JcRRKOConx7Ao
SbydAXFl7lzkQ/i6aylsFyARSt7YygfwDZbycSnW8L+ttI/27FFvjF3DdJoMIeLk
f9e5oeddzEv55RgqYKkk8KUh26NJAKKrrcPqrus75b63kPkcSFDq+sD/qJ8SoB/w
b9sw8WhZrBOGQGxEQtCgTD+iopBW7QFiQRAVrsD1Cz5ZMT8ViVhUqm403/RwJYfu
kSgPS6z1W0/d08iguFWvHnDAJG2w1WBVzOh6vNnze3W5lOXYFPiTmGdbvnPjccEX
0BcdoqmjCQF9+n30yHOXsUEA8RAc/vA9d4BqAaUa3t0E+kqoBJb0JHEoVfDt1euU
EekNSPhDuRgt8B2AKC1AYOZnmKLYDqpqWvEnVleyNkgo6iEgXbl9MTl1pASOCupz
Nnb98as63q3tYs210+xcQ/w8FjqULmkdEibaImvOtFhIQ2RVFLzS5tsOSwFhkO2O
fxymh/QA8/Gr1WFcVdNik8vupeppMLfInnKOiKyTiPtOP/W2UzMt0pU/3ilOZr9V
Nx2e+Jh08K5T3r25bL+uWyHmK38VvBynQ1ICHBG6Oc0mGwhfXCEw3uLctbxjQmtB
ulBt/41aHsq+tDJVrFGs+eBggncu1zM5lf26kFD+c4zPRMhdqvgV0dgnEA779Zhv
ywpdYtHUC77a8fjAMw97ZZgz7Q2Dnl/zQDQouA+gSHGqkW3VwVeRjeVb1cf4Rk8f
iD6Letm3aencHXRd5PKbrJ9FbZQfxU9l0X2PmjSS6OdZlWd1WoBGO7rGOfo7tfWB
jchrKR62Ffhl5+ii8HGdjnxGPCrfkmzMJUwdWdWo/lV4nWUkBhQ3dBa01v3DBkxG
9jt/maK+H8XqjgVtNp5iJHxFCoONTLzGlg66XA74XJsxdrWOFHkYsqO/6wP7t9K0
O3YrEemS8nNUZYGcZS8I+ZsLT+rAT3mkNhoIrN0OiFgJ4VKl+jR8oh0541piBY9e
ZvbH1ya7LWSPW3DoWyBem7WHVb1QLj0KDQzEophEkYCez3xtiVAiVloOUYehbF7W
XjR+90CS9f2fnbYT8hI61hvaC8X8WjFzcjJLfZAN3CnXXf3TUvgQ24/mIZqTy7AX
VRNGC8N7cffVd+E4UPBW7qEp8tjYISPuQicvlDNzVihR/UxwMhYyM8RjkYaNJi2y
ZXhixqVt9VnZ76Y2TS5A+fCniPW2SRtHhl0P/+XT1PhqHUi1XA6+X5U7lyGxcaCz
4HPVH+0OSR5bvBD4Q6nkEO4XX4HH83Nb2r2AkUkDL45wBhwBWaQhunj0JAq5urLM
IYcTFWYic354SBKAucIoBssuyyY0cJq7kCGdVvUDKKiEK6Ku8r+VnHi+XdPv3zwe
tcCA2FlmcE4s1TSc94IsldKNfhaMwuu5BO/QXbEwq/0tuVxzfkqIcDLYvbPJ9JNb
AE5dszg0GRgZTxxXnJjmPtK32WGzjqGWrGCTQiOUCU+cGcjf8hnc4kMjeOu9JtPA
8gR3RznX0S8DaJnSsdC3U7SK5naBYEXyM7OWRWCgkjQWhzf3OrmcH7/l5Ssvo0ok
DOgs0JP4VCwvP4OD6spHmqe3AHqt0hZjtQG//Y70tsMTPnxYKdUeHN6JqqgwvVto
unstXZ4+6viCh0wYl+IWHegk88snKiPfTPnioygGAmHoKeKHYVDbRfB5ibh9hVZs
4nYhhFivF503M4HngcWWWxECmjGdEoWNNKMVIyh+10o70TM5wq7Srf8XfincKgkA
d44var9YYVv7sNSeDgPYSRs4GZlwJo6GXlUagF4TkXL36VPiw0WgpPiH1v/0NPNS
LHfKikMXb0DAUNHhb666nRTV2AR1v8o++dAn5cgje4YSvw9PX30BcA9NcMzuTW3/
pS5elIC320IjGEkL4lSiN0ofkPP4PZdnG4v625GFSi227CHxqi6WkW2QYGmIRmo+
9hDISnD4Be0vWfdloKH4M4jx9ImdTWUGV/PIf1GtskY9IjLlZ6JOLSQTN1cyCEbp
sPD8sVVSiXQx8tYYx/qyQZ2R7u+00qiZqyviuMgLPr/Wcf7/eyaUugaCbkQ9khqf
L6C7w4mIYp66XylgOPswPYS4Ej6eLfic93AbS45idMol/qEr2wTHQRMPeLLUlPcK
ScBk9WTawlAYz82qdXM0fZ+QlLP/KUNLtVlXosL92YgVLhTq96gzDlNbxUxnfzp8
kT+ES3QI53OLL45tuZ9oZ1Zvw8aPt7IrCjBflEiJ0ZLsKEyIwHrcogXRzZoxVj66
2A2GPYxfeXWhCv4qloNERlKDYC1E8/Ri3YrguvTemzsw1wzRXJnoaaPg7YVgGpd1
06ozeTdHKHx5crmLYDeAip/IFowpjOblQk2pv+MOkpnWG9P7ZsYDIW8KXrc7YGIZ
aDv2IeOGFfo8xCaQTg+4wTp1Vol4is7H87JfYCjgBF312JPl0dkqIonVLMetqGuH
xc7gQrzJsm0R6nZzWHn+gK1kXFwxfw5cGvlhbFqZxojKmaf5omlVub2xjd4gku8P
TBjEBgRLkBgRa1+qmT61jaRAE0U9/BcHgRVDGf2yh+m25cxz9HGuwHlvnWCcs+nt
NvgWAN1L2W0c9s3Yq1fybtu8ozb5EU1kGLT2D8EecAwbsL5Y3sTqgdSj+cY2TtKW
++nv74z11VEZDvtyLmr34ZwpYqjHaP1a+atYieIIDeQPrRuBHgHuPvbVzFQpRxMF
+4QU44TBtfMrM4u2DnlXpO/ruTfv51vKeaKIg+AbQm/I5QAbWQKqr9wrsZoTasyG
VcFSNFOhRFmekqnCGnRH/IMIWn9g1oQ3oGpuDXXHnmFaeN3FE7tbo6G9cTcvNBiX
1i0UWAFKL6pEcmJVUBfGpvDKSOFYdxqBD8ckOhBhyrWsyt76+erlK3MhuJ76ECBQ
MzWymoYC6O1wcr/QIkTs3vlYPCy4/18IRzdTT6X4P6m8JoUdufum04Y0/ifD9Akr
tz1K0Ybj2hFYWCgQ8C7ooRgPrUhMEYa7Bs81RpyesN7uOYS6NKX+P3MFFW0PGJXJ
bKa2kawHP/UYFa7qfvN0/OJ9wT++tYbytN8MZyrYyEbwcHMhWOyBOMzeq4osDDPf
ZeuI1kChgALfyoiSw8tYzmai5g2OzZZWbKjZKcdGZoXJwEBY1CW7V/gcXWjkJuQl
/+G7BAByd15ezJF8R+CQ1TRkL1jvvrD/PMuprg9AtkrPhUj7L8yv4SVpa3ZjREgy
BwHv9A03KQm9o7TtASuiQFiIZQi2rFcImk38f/xVM7KfBh4qJ8uBIhNj9X74Fqdr
pOJc9HTS97yY88YwqwscNjxlzbXEdxjSDZBnfVZ/IdSwxwYPfoC+kjeQcyEOBeoN
VtaL49cC8FuM/Y+MAzTu7Iq2hSpkrV+Qk/UB31jFIwJhkILDxc8copBclyKP48NY
apZBxD8fx/6HiafXHA+LGSfjiHTOraBInlzlxrMuPEc7eNxp1hBVUld0djaQGnCa
YGjw/cxFEQapx6R/M2Jajf/qLVJiMan4N2WCxUlCmgMiqO6VZUg6hE2S0lmQZ96a
RwB+kpxbpuUcV2fY7ydxmgA5Ics/HPIRnwJxPrayU0sj87Gzf2zADiaW4OLcVOqH
2m68Yxvamj625+lpRniyHY6JqytRdYAZBybwlZTQDPlt29ksjLROLBl4n7V7gy3q
U5BsIL2e/K7H21gHHDp2tHLPICPbP1KHJEDAGKs6CsKd8C9sj7SB2ANK5hPeXtpc
AQJcmfDBJn2zh9qyzSDFzQ3xNqcQACh6bDX2KHecqyeCdGxkUFHISl+KO8BDGvLF
xIrpeNwjWkypn0Ibd2y1RXpHz8ahSrq5encvk1gkoUMEadm1gTwp7iP9h+d/T90i
+Bjy2uTm5+C/AuzQuOE7lghnvyjz/cfxadgvsReZPNQn327fRHe0JxfitFQPxHdX
M6gQi/KSzvDXq+QC/eTPuasmQvXFS020JZa/VbvfqgVKwM/QeOZ0qErKmOVR2rmR
gPtk9d5HTlUvvloia7wcf+7MMfnpTJtvtiLfT37LgBQYLASSsbkXPGElcSjb3nyP
eI0nG1Kn+x/1jX4aqfPywKu6K0aDb9g/wqmfeWIr5U4FNLBNQDDZ9RtmNieyaei9
lMGjQwWbaxcBWI8ciUKgZXpJyec9imWkSnyZg0LOhXkVWvSOVqHw5kdPPXnvQoh6
I8SxRcRPFNJ56Wk33KqLu0bkr6phfH47qeNZ39X6Z0tsBoAP+qdg3fIbYvV8XTQP
LR3Pm6aU2rVuSsmtTcEaTp2S8Idi4BZuUXlHv8CsAxrzrrI01vrdN41xjjxKEr6E
fewlv/BTmAWEveqRapUWeto8UVl/cp6NxhJh8brfRoYVeY9QWti5r4ASVhbynC/Q
UsiwkZ3cCwSW2y1JoW/+NRlm5GJ2JfQcGUjeWXU5fhzTIzSauEnF5vUzSzh98TKY
FFZljlpugawt5DD11E4Zk+JUYlduY/B5dCjPyNWVlbIMuqAi93f8H8UDouHMBAKP
BlyxjXYs9CGJwEnum16P2eCR6OTGigN5xsDZ8D4TCFz7EFaEuw0Rd/HNBSjwfC3w
Jza7qu8UfhVOVr3YEdJKcN++dAYrDivUL6a07nCkwVPWevksDYPcZMQwhDEdHHm4
N3ZNHEauGlM3qgX+43EJ7kHFXCRGzW1zq5+aFfRXIs4bkb4KCiNOl86ztfhbpC7v
C2stJwpnw4APUbUsseHnP8oNOZAKIge7ixWOtnP9H1EME33TQ8r5ZHdSwS0AjZIX
1m+AtTSDhTL965caJqntn6V5UGcTbguvSpvPrXJnrozLZHFLkjq533T+lDtZJTWa
Bn2eFv/zB36o+TsUaUyt8kbHgAMU4tK/sWzBpnSqHuZ+QTk9V8mUmB69nipkeRX7
uuwDpl9R6LGH/Ur0X5Om8Sd2rF7Opha4FUkWk1iSxMrgB+YRhtXhxhjjSR2nlJxR
XsRjXejVp0hEQUhmNjT6Gu36ZOYplBHk6/sl+HeqQtifK6iLF8KrUf+wXDumc0Po
SYDJo5QD7+phvoXe8a5PQUqQp4I9VXGve1KVqa1Ne5doJmrGfIXrGNEdMIX6pRpa
j8L/T2sSrm2/+2+pky8GudEvkCgrtgiCH4olejJD9eUKiqvSehY2Hvj6lzp27Oby
sIYDstxGSsMbmK+wQSpo+jJQIdBbp9ieveyzGEU75MX2Q4hM+6JtAWe3VKMmbehd
dqM9/n0CozCC+8A9ctvHcTXYepnr9bmHuaS1D/7x4PoCelwIY2I7KdRnfnSKNNj/
ZVWlBizVuZ8Yy7yxwlxOtspL3D8+vacfFvKxvykpfaszad9wn2zyc7p2bqdu0Pzu
2GABUO3OWqwCr/KK7HkVtcQnDIKMHPaA4XzFMmpIxzCWSxJJrlCRIkUOTxr8Z1uv
Ws/1eHGsDfm6dvfnEIHDbHqmiAJyZZ3/kfpPH/GnFJ8XITId44vcZUqSygZmdvo6
E87QI8hxr2fl3oVpIdnHUbibqrjgtcOKmXrAz6CuEgzp5kI5txolqLWse72IZ5i6
X1lW2baZubJitWCJC8UvsjZoPEQYeZELkDrq62i54rIrsIflmtn008TUr+XnfK37
eSYroaul+G0xxZvOz3vTB6OAachITzmymRHEvMWiyX/377J0X0G+hRW+ICwwxiMx
Rr/n2OeurTdX50H2s5K64G9NiTBxgcSXKGdU0htyEi8IOOB07vAcojHlid2RuPyt
quEn4Ki7hKGaZiSh9+uS4zQkf/Sm9Gj3Ht1c9C445thD7/5eb1EBb/3rhx0vJZF5
dW89c7Ae0P3j+PbacOfTLcjXE0e8eg55o7rAnopoIspCt4S/ZitTgzJXKI6uVNny
QoBdv/ORi/WA6MXw1UGbf8Pk8FRIb2ESJP0JRryR9A8iIdQ6oCUVPjMfkPdTyJ5Y
BcV2pwWrzECIKXWhYuzryyekgHBb5/6UZo9SK6ZlZFTGh4MRo8vmKRjdnLv0Avvj
b21+QYm+kbTj/oX9g3fav97ONd3HirC6oHEByotTjz8JWJf35IJU+egpmXyekOuc
UMq4DeIsIrEVT0S4h+W5z9qd+ltVjEvCTxY1DMDoBZP0pJoFbmuDu7TNg1l03xLD
ol4ReooVPXkR620OuQXEXwMbE/I4ZxsCgQiq1BkekmN46zjIo7htpWLElzFbEwPL
2s9rTivSSAByBiFqFj6VA7V0TvW8yiiWDSXYbLZv4yXq8tuxaONTLFUxQY976b/5
Qz0jKOOfrwXIG2ma7r9LJhnZJrR+uzoXNR8y1Jynh+jxg1BojBaSXabm25b5BcS4
Yt1nH9QwfUjoXBsJCQc2bzmIk6mmJ8bH4pBHeQ3KBM2Wr0og6ZxE3A6WTajfcK46
pn9NVXda40Z+I6TOR14u/XUK1MuyknaS7Yu66CZgdnin6iU6CGdLDgzeSUyCP7ZY
67jAoKGdLOqkMDxRnBe/8SxcuoMKEvqm1EshUP6uNA0MEuvu8tsVnGaP9jbr1uBx
v57O61ruCBplbpkLprpt4vYRvPijeW4bIyTzr0bt7ZQA+d86a2yDDyjBmE4Mozat
0fUXYPFwWPMcp/fuPSp7cojwk3mPNIIQJIyA2BCIas3QBt5OHqR6hp0aN04REqiV
H4NNUTA0EY7bxVyqA80aY9poAFc7QbSwJh7dmkpAurMzImFEem18b0UZS8ON6qoy
/Mytf/7WAp5qMnHPB9iGV8GRAj6fzHEgYWTpn4nwP5vW+pFm/IiRha5rW8n9jULO
hPmUjsUjpEC+W2C144xkZAAsK/3eykMZxxcr0N/a4Mvh6lO6pGbU2BTpS6qLK8TS
TMbkt+Ur8aTv2UXK6QPN41a2Qt4w939ybcJPLbFwJYK9rhXi5CCGonMCezHwYMiP
INdLokDbYSTQCDJNXG8whwTFELRTba2RbI9tqcYcrXm2ViiTKA0T2abguIO7FKFD
ZZuSA8xO/MJKxZTGcFc8ArBZIPc4crpULESQp52bHYzID/T0HpKs12dYN+rvKcw/
hGz8dGfvfF1tnSR7Sl9E5KQkuiid0Jp8H95fz+5UA7NBv1HzqKF+gPgCUV0TsPqu
vW6mju/UBIZPC/R/QXoC5n7mcqRSnD2tHi/WsBb/JTmiMuo2ovSXMH3WnfQhZ9xF
SGar/L+Zuva/UjyzkKWjWtUV977nQG8QUvffdbamPrJprzBPBh9GZ9B8jSu9+GnN
Z2AV34+ascyCGAnJR/KOmDYlHyiI7v06l0PT1OGQluSBWu0F4Tzw8heWzSYYEFw4
oeYUaan/ibJG0+YEf9bxtS0U/1vwGQIb61+k31arCK8IpGa55GO8Jb2q4zqXB9BR
f3vUPiyAMuAgxyGrWml3HPA1VyEi5OF4CewbMnu+ILu5HPo4wNxCNMgJhC4Jf1th
ph08qcBhVtlIV/Qp/1LZGzZLxaU05ekmaeSHkN67oy8uTlHZkE8/RGkheznL2+z+
gLMcrtCHtlJ3XvZvVRq/F1IyaRwnuxA8/3uB+oTU3pfSsqyXZYQmAJk3AaJ18KQ3
+8HPhxaF5pRfEC0a1a8cfDnfLp7lfgqq6S2Ma9M5dMIY/uXHAMFFhwePHElIQFQ7
z/w5fYnuyfNqKLkKsSGpM1/X68VxggVISUcfQVGY9NR5YDnpaA+BauRTGNGmuweJ
dK9N5BM/3RezNCDVvM5DXr5OOaV2HToaMY5WdTWgOdLg4syQ9bvRUg3nyDtIbEav
dGpn4FvafqeADkwrxI79Oi+K6xrfT9cVmZ5hLqxqwVriUAUSh2G3hyCb4xNOiq+T
MS1soXlsQclXjQLE3nisbICoD1zhI1sTQnsRPCqsCro3dTTTTALMa6x4ZZ5Iuv4w
31xvAL6txdXMLpwzdIOgKQD3FrXz8yNewux5Y7rmJrOWw3/qUQ3FkCis93M0voI6
G96j4Lh0D1/Wgmu4hN8ihwztfIgT0+oz+NsLRUCwK0nFIvAQPkDKfwb4YCA2AfY+
/Cs4GTgpfSQA8uk8ZaaNYc3B6gkdjZDPXxoleYk5kZmaQd5HH1J/WJ+GCHBGl6LA
07xwy/qKmSyZjp3ePVHq/SusOpsolFpi9M1iwLmOykD7rSd01PS8DGjbklA4YucR
Z+HndtWnMLbCYsgP6gjUPj60eDLcifptf6XTxisgkzeMhur/omsaNZ7SrpnOw/sg
7M4UBaOswnP+TTJKnsHRqNAkYsdxFoZVAixtjwL3y/opKcOx9w1wsWkc0lJUqjfM
7OWXIHy0i+xKCyISzKt5oTrmfzdoGFQYBXT0SztNR2pBBcfCxN2VSwi91V3ganXT
yKX1tsazfrtg/s/TXk20dKN/w6wyF6D6nH+pZoYIK8Vx4GREiSAdtFnu6cZe3I5p
4TZK2RrMMDyKVEZyWDH2iUUc1hc8nbiJER0qx7fV6VIm6GBirrGp4q2hSwk1ced9
Z4GWk95WWOU4NeqU6mAFCethBIRK8i3RvlWHkS1X2/oxoY5WgPW47vVkbYjh/V72
pOB0fj7Aag+I2pv5pWMIbiP1p5Ormwcz8gDzsedpdQVG9BpbcOl6r8P+18I+5ufv
aYumvQeiaMB2hEkR24yWU0cqn5SwAB3IB5vVgrOK5ZoMJ8lbGyG61dILtbiw2vPN
F8hRoj7fmZcsVD3PBWUv+y+RXpIlt18x0Xtq/l3M0zqgMhFnBSJV6N0T9n6YB/9g
UNOU+uyQrZLLzrsdyHuAJFF3cLQd78q+U8gjIY/D0nSKICL0F/LE3Ne+VX1zmv3Z
AX/rVEMvNDXI7Oa6geeqKamEUoQtGekWTpVVSU7/kV+cKNFzyVsmEvz2IP2+fEwg
6mJvilp7kYMvhnIekXJJ/A360+827WE87bChgqJIkZvmyAN6EaMQqXZUX6dDITYv
sttKv418Bucvy6+F/7PSDHifwn6EkUH9GzjxFpHz6W/nqvBwB1J71TpUPRD6R0cA
ixOZ3fBdpnsrBQezbUlrwvyIlmIWVY5HjbcHu65dlUV28PysuuCA8bJ6/gEIV/ZM
7NjoNzP7L7hl+0Ocf3zZfj6eiEDKG7fy36Fpv3qIiUERbeIYJcID3T7LT5RN0pVF
b88TpCV4U8WhNbNmjRjZ0jZgfzwLeybQciUT8oAqUUdhT5gmHGMfDaRYgM153sEn
Z1KOxV4p4F1U4nUhj/M5WPH+y4pooOgbBto77ghBn2MKqxfwN0hXcF3/KGRZC9N7
4SqHgVFiUhfxssVw5T+/YOIVvx1+ej3rAilN4oFweNZFIdgdNlu9EwGkl3uo4Dk/
q3JGHJemZD2NZugzr02sEIgSRF/HhyvBvRZ3V+kkeLKjyZ5ovrFCij/JEgJ7dJCO
xa6zfsU+flg9u9a4NawJqBTyXYjnCyXm+6TdEq04SASvinZyhLocJTPJt1W67LyA
WN9JWH0IQjzf/fKeb+fLR/XQaRaVwc5014OCOUA4G19VQVfSBcmYhzaFCAhVPZ4h
KXA4ujPTZX2qrqR76CIrQcaeQgqgiUiKAF+5WLZdJag4sdZjj/kvsecfs5QX1O9C
fWL45F51dT/wXgyCR5OwTJAdnFqT+3E9hHqr33T5Rbs4tOGHS93k1HwCCobIFvx0
9PrklLwHSLuEyrVSQLYK1c7k54yf2+m3Dkz1kKfd7J6Edc7027LrhxLJz7xX/q6X
SCA2FoJuNoh1KKSTCM/8/SAuljH2XnBAXGretuv31y+Te7dEgTFEo+5/8kxWbU1K
kUXGyfhqxVqrbJSYZVburFoIvSNw9knF6s0GgJg0LJCIWfi+s1iR6+SE8bSpkGnM
azaWXw4cp9CMVg1velWP4OmNsTcXWVANuBkdR0hijt1eTcqO0yGmTw6HKP78bVsI
WhUtc7BwwzUH7X6WOOTPihbYlHGAUX5ZMcx93lI/Ecgvx6KspklATH2IKq8grASe
/nfdEzzIqTpaiibcDx/VEd7aXYW9tIFLxmVSqATlBCuy8et+m3O9dyB/dg2BKSwB
2KSrwu1dXzMn2TgNiZBreuKx45oSc/6l0TbO7ejFS1K2diax2uPMlfmfj8LC1POq
GH/fq8Q3VglTJdH2u3xueKQfP6vIOsb1rDS2ZJ9YP3LEgNM+Jkacs9zaTAhPs4jI
19kfD9ZADKc/XgrbUxvvSV8QfRomEykTXaEIg1dW+trK+706uHmuxQyEGFQM6aGQ
NsN4JPb2XMqKpDMUJo8PFMPyz2sbkbc4zKeaoREmR6dTblWEoT6oN+mK6+WKhrTM
UltZHzwObSf7IFuJHyodhAE4Mp/FXZ8wDCQHC4a4gFONwpxUdnUQE42Aszyk8RTt
7Ih2FFBqCACj3Gg8IKFtb1qljLHlFoALIs2sSyMWGDPuVWgM0+TcpkWWUEdujHXV
D5iQEp3OdnroNqUOxXPej+Jy0iOC07BNrxbx0PMhqzEjnSsYSs9K61YLVObGS8G2
ZApXGTCnj3BH1MBQhpdLg5503Q8CSMnCJWKjH5t9Zp+jLnpLKFiSLmyQTKdJ3Q3s
jFZyZHnk8KjM8l8cGJ8wzKdrpqr8XtfphA242v0pjPIceSXbMQ/+4oyn4cSBpf2p
9vyqskfzYOMzuV6DzDYkg7uSdYO+oS27Ixq7d10/cEg6mS7Ca3rk6e8300UEbYKp
KDj4fbkeMaofRWfurS+E5G10o/dBgrKqZkyDEuA4Moq9HXhFUG0nWOzOUpKjJf3y
CEiiOQhLGZfi0P+MoO7LXzURFC/BuikmoWnNIVpA8aw1xTACx8yad0hQYOu1cNLX
CpkyJnpYiZ3WN6UUPHMXlh8usM6mkJOB9/lSorjhdQ3O1vVfudt2QS4FW50H/dYy
X7nre/l8LOoIsiELckHM0cFXkJl3thSbJKvQEebV1hBaB6zA97Z20J1lGEcydb7C
27mbD8rjj3ILJ8+en4S3lcxgzTVx/qtbtCcSn9YUJAcusWvzLUklEkkIK7eRPtu8
eaFVbmjj6mmNNG6SF9lJ8sCSHacfyKOkk6ph010Q7Pi5k1In9/jhb61Jb7QWL4fr
1wA8k0QLfKzUDO4q28+nKyYJhztf87jXzHnGIcrQ0xxD7z4e/vXG204HUFFXt8Yc
hCnqkQJG/kymXbHWERDg2AdflMrBzfzlHkLHDzt1axKgCAB97At7y8qkthrFIGRY
OLeMJgxcUf0AKq6Ru9I9aZPPRKvYB24IclNwMzm4ESr9xzuugQH5+5wr/c8j5GpK
5plKOnK+IH4yPzmmbW9Rr1ZaAQ7P+zC5nIUrYJvrXpHwgHYrXLGAaySrCNaYTM5d
OgNdBHjB7SW7KR61AkZAzr25oocxQTr1upXI9OkLfxclr+Lr3filJztyQmQJ2oxs
JSFScvXwqfE8C1QCRnavmAg/x0B9kwX67a6loZJ6h+HVH8YvIYLWgreUOgC14V4E
ILnG02Z8KkFyf7hnVyYdhRayn8U4ZMaTkOjKS7WsylDB+E2lDziJCUOpam7PxlrL
2HHjNjkUl9lO/K33vpmYsXC4N3rfXPfaM0AKVUEBjc/UMfq2dj7u5fsO3b2+UWKw
PzA0AIQSSq1gD0zbDcAMnq4awUX6uBtEa1+oZGiZhRBleUgjp1EtUUZ+Iy9z5sRc
WnI+EVomURYCjNQy4eBIhkvMGmTegPCdjrP9d4SmXqIsGEUWnGj5IDTvSmLpYPxQ
r8AsrnMEpC5zQzvvPEngV0bUWLwf2RURcvXQmA35g1JgK88iRfcT8ZDooBAErbA7
kv3pAdRuAn8McVcqMwjA844FKG9+4L3u6QPspihC5o5i7If31wrcChnMxtJakh1j
UFGMAspQQZ0W3MwshKxdqbGx6WcpxNadL6CVvbwLnLzgXH82FO6KkVW2nBQ7kF8b
beWq2VmqaSetR0/ORmmZ4bl14+alERHmhVqUfFWlUMWJ4JJsZ28FykB+jAW+tRCS
ghLx4qka764rb2e7d6WKAu5ILBc3yaVNVAHrRtxc2CcKT3oWj5TPu5qj4etPc8jP
bbs+ohRkm7iUXLsgsytWUECalHL2ldKwmXWpsMrG89FYURqrXAKVxhQh2pP3NC/y
UUagVtl4QDsnaDmkHPwJs06crtpIWWCqOH20uw+hm7VkVBvSTqhiFZ2OJ2nwTUOt
rXqG6a/XAYGxT+5+EY3kBfjRStCljeEsLyeZczcOYK7JB0dP15io4qv2uDQr5+mQ
TNuhoivklQ8rks27wFmiwscOaPJb3FdqYde7jwl1iQpJA9MlOg7dBl0UPRFj0PVG
2S4KsrzEjOHfPB3XO3RjYh+b3CoEuLGqoNk7NxMl3WP0NsIZN7s/q4RyRmJ+9q0j
muoshb/oB/gT0fTe8F7k6ndllnlAlkFqcKMwXwRiGavTPNWpghDak/Ebhlrit3EZ
qicA2DtCqRNu0Bom+SD+9w+qh4bygCxyK8JBrWksfKfc5Qzhe0UMbKMxO4jTEZu4
w4OSnUXE3pzgj4aduTyTcdgh/BgIFmUtJSuS0rORa2CHZm47LxlSOqranx0x8vsu
2TIvAK/vL8O85eg4M79X4hJY5oLujHtfZMXxcW4rzMq4ZGFo0OuxFo3tjoUipMVr
9nw7iJ/KTZoxaRXbcKe7OOK+Kp1tiVYDzDPF7b4cDx5jDr1sZ/jjWLvP3jz9Oc5B
54u3ygrLZRCUX0W8cUsIxTPYl+KW+MFg+U7rMVqs3f6dX4SVZr0T2ER6WYIk2Eoj
HcebdhheSiaVY6NZADr6j8CP7BgXrST+EfHYlEEZJ9GuxPsxVY+9Z3yDnB2Kcwfl
C+U/wKjn+6ADSCM5h5ccnby3cdKJfy7ENCDGBseVJXpmStEowxk8zWtt2SlJw5mJ
svCY1PTlfUT+S0haih+dwGCdJb96xHL+Q0enuS/wrZFahClVV8KwNg2qJXh1hJ62
FhXxUlg4Q9V34u4G4KvKxjGDOiNITOexnqwNZc6R8jiMw4Z6yrcqH4wmN++s7T3x
RQpNbTzYdnsTgt1atCZ7VbWdAl0nl484Q2L/GKkyddY0rrgyoj4mjFtEtS1P5oHL
qNwe3l/K1P+WQR2KHDPTbxWKbRsXme0ObCKElHW/8xEm6HqPwj+wVGELz8cYMF5C
5Xl8qHYsZe+p6d688Y7zUu5tVtfqFTkVT2vVAGnQh5gLp8XXweA4argUbA1V8oxP
X0OwYPnjSAL/OJVw21vBU8J+590ZGKpK7Z9ksuyr+UUDG6qhLGwRWDjYthDt6Wk1
xL9P6cMeIceR/vKzQk419fH6ErX7lnk7BpmcD2i63jaDndeeJvQiCSyZD8S524JH
gE5mdC0EpO3OM5JcRXLJyLcTxxcojfoitGExmo1hQkN5lE1E3lvjsz1t4Ds7Dlp+
crtDB7e+ymXK9KZhvWmTTC1vvBZCkkQpc3+eg0zhUV3CvWDlj7hty9BT11NvCCxH
lKKvDRx2GwvoFsdQIYXGWyU9A3lXtg/qorw/0aorCMGQQYhv9bpH2Os+vqZ1WtOa
LdPVQe7pG2eBwoxMlDlMGnLdNeXySEO1O+atr8ncwMTxgxGIlsIzIYDimG7YqNKM
BTd6WPVLrYBQB4TYfoN6fb0hmMFTv7VDU3pN7phJ/5dprlKULZfH1qIonjgVSAyp
O5nQci5LNyPyFzDA3yPmcmvF9Pz7hay6Gj2ZZtGraH/AOXgcGgrk/fAp4077K0TL
ixAsJEXFTcc4/Ld8GnUl2O3OLgs/kjh/IQtE2MOtA5Q0g+E1E+YjrF0GqpH4lHNu
jE9003zHnSzohWvSrpyFTv/JAlK6eFYYA74+OpRdI2Ydd+SPv8TJO7ZRzy6RXRpX
QILO6azzNwlNLGlFI1sIjAnYOeFAZ+Mq6VE1nbB/Qf6tsHL0OuZiTZ+b5J0VPgDi
Zd/1Pik+5ZmFntoanrMrMJt59v7LvpT4AMg1s1gssVyAU1pnJZXjNFnwDpzgCKLe
3kOzqdsNZfgqPZ8478JvbVWdacRkHbI6yFmsVEmYu1M3J6zhpGJ35KvCc9PyBAg4
rAN2gG5+u81a7ug00SSZaa+Q1yn6wASWQ8p9T8p1ghBa9SJx4XK83avXPMx4vV61
fygzIHXhlkArPRG4EP8r81QmychPsHG/A4BstBvhYNdHDRhXeXk5A8zEjISdpWVo
j60DQ/zC60u9AXOu+6uwXhVUrIeC6a5jHPT/A85v/sW+euCZeQvIgpPWh/LLgJbj
rL8tkKxb9BdlzcbsgvKJFsYM5zXC560EamfOt0NEc/eZa5kVW2Mu37FyYj6pGr/5
IppV2l5LemvZ7klTH+fmgTbK7WExsOI/Eh1AJa9Xis7uTKeIiWAcvKEMmpS6QyM2
QuEPcClhL1slfBHZdGLc8lFjuBhn4LsKiad3vF+GcyJs7le/PT2s14ecwmga7QpW
nUIEoLY19bqPzSgNrKQvX4eUFtXeQI3Vb5NgS+M47yIgWpmG9K4XvAhH0l0RSfAk
jJHBRWAvwBT/hD9rYfhodaAxlMqiwc1bHZokjgGHxYXpcT1VZbjzInEf05FVkcGA
oqqZeBWI+ZQKVJNNQLdH6kcNjgR3boQ4YLwESoh2eqjDPLJRc2EU2JBfvd33Wsxh
f6sYYVnWgT5ZtVTSMna2OXoeyiYN5HsyJevyBG8u7HttY1E/i+GUHyC7vZXyuRLd
HgjGVHu/SddwuZjarWKp5iODg9mC7BIzzN3+aySXSuiSrQYvQpf/c6djKuTli8Fo
B641RFfWykPFB3ANiyzuE4wVYf9po3Sd7o5l7vUtKhwkZcDATHhjKqCCvKobMG0a
T968/BBqS4SGLxPYmTaqg9rRAW4Goiv3aTwV82nFOBtpywtQWyVhWTehJts+Om5G
LRmBkeN4BX1TRSE1Dc78oYJwOFgeuvwFCdFmqbHT8noH7BcBuxGgqvwr/YWCU5in
V6Xu2+iVszxAmdoBCtxGpuqGFZEBnpf5ZCMup98qeamb8GVbTsRbsPBHBls2+CVk
rz1cN+V54jo5WQB3oTKCgdHCLi1HuubRZO1Bfr0f0Wxvt/z5FDB9/zNV/7ZzqjzP
of3GtViuvrhKELzW38ceUxfVLdXSGXZtge27PlxEM6H9v6q/czF2fjT61YpnvCi1
KMG9A49jSzKhVPZ3sj5AwBzS9PLd03R6oW+GBLFfDhymU0A2zPd5qemP6KwEbkT3
AOwy3WUlh1+fXtWZE8LMnB7eC3E2lUgMRiL0mV542/9UeUSJvY3JxldAsmQNbuAs
m6Ozhu931uoDFLCYVwSWTs5ZdvxinqH00mwliCxxHNp3spw6C1po1B+93ognWqKM
Qmpk7xUcakHsUeZBSNta/Dct0T9WQ1Uz9bX+qr0G22rGaOlh35BPJBVlKdc9nHhv
Xh3mDUkR1xvB132TafapelQGbM/q+1GzmTxmPc7e4jwg0RqdZkx+vfPmcC96IeM3
4SvJ1jPI+QVC+waFn8oFiqH2WzWUf3pm3qVoRnk99E3pXvuguIt0Tv1kpLfxiE+Y
SKasyb8LRszMwaDv/eKRU8KKbJu+r+wqfXgYkTyUegKwTphjFnETpAnd+B/CwgeV
5f/T7/oyEulJ275BXly3ot6fj+1NXAk3GZumVEFtqU90L2GHp+E66ts96lG4Nfma
PkL5HCxWK4hkOx0sh1Se4eKG5CqzYCh3pBEaVnz8qi2iup2RpfBhxpoh0r3X6FzP
49SHtKA2BgreXXiFgU/qyspn5S0WZ2+vonra4ZNuC6jIllZelJjhurpZHJuC/PTC
m6KsKZpWTYFojPbutHUm/FgYHo7ZBzb97nRrm68gfwWpePyPo2K8p6Wqre5w+MFm
D0Hk6Xyx7+bemh6iLCFrBMiqgRCj1AFlhUGw1zI67UUrN8AoAElD0UAQRCm5R7SV
wkbIco6tSpkqejt6H4UHzZ3o0AsAjs4xuSfQcOD1VcrBKjAtUnUaAiQQ+1AIbSmF
rK3m5t48bfm5uNhGJEHajkwKdTTfJDYMVJ4/Ff1wq9M9U1yJIwq9sTnLXbNJu0Yq
pq9Atzk8KYANvB5BJPAG7MAqVYIelWkfkTvMBZ97e2VKXo5GM+5fnFNAyd8UMc2/
nejRdMlXmllqu3kTUzcST26Zou6hgmnb6Dtg5ubsKTLLf29c7jid3b+PYwqfsEPo
fjym6OtdiTMC5OTw6L+FRwPjhEfGP2VZ/RWZ9HFmiFK+WqFT6dODWM3xGfsVPYEL
g3GMM5iUto0Yj3xDTFKaKPDyk0tXKXXlRTA5jjXPe6jw3gwVe/BozkkB/2skh/fa
TWIdnsEhe0no8iscCohAFZ3Si7yPsDkqTrsEZ1trEaPVO8havjzg58fwuUjJ3o5P
WWToc1qGkT+W+zf60OUd87wDQ4K+P6GuVdDIb+kqJYZ3aTzvBB/J+vvJG1E6w5cE
ve6gqiYIBxNVmUvHHnezCUH+qSMtq7Lu3+7iJ6EBuyoAsjmME1idRpabfWrp8JF8
rFQur4CDz1uY8bM6H8QrHcbe0gKuYseL+e5xyrCsP0qu/RD9rpcQ+C5AX/oHDsmz
ddKEH3OCAjM8fFMMuamBlenpp8jvX6OR5nXdHcIQWIt/RN46votW9IGVPDWw5P9N
NVwtIb3kYpNRPVYnFDrx1kulC4l3uk2XmlKwUpmR+y0HRS2s+HyMOZijdWAbBOUR
/g9FIyaVfPQLBHdO2OiOh5estSwtDbuogrv/+bx+8A4gcyf/jCziqpGxroQJKyFw
DsqEa25Ep319/KFY8er/+Nbwkg1PJq9zb23FME0ZckGcnfmzmn+vgy2V2H0GkVJ1
VE7TBGdIlOAThquaZFGoBWzUJENls1pXPIhi7xxABh0O3WnUi/gKPytyJF1t+KI4
258fjDyqdZ7FVHfKs8XPT4W2C19hWzy4RB1dEuch3tOEvROue4HiQ9DF1deqJYEE
MYdipnGzg0a1F5ahJxmI1m9Gb+MhFZE7MrP3L/7F2gBtJgVHSpgNKglOpsQAgvGO
a+vTVmJd6Bu9uA72bi8QhYI0gOzHN1cROe4Y3H4xnrBvJGMFU4TPsuq2LUm5Q2Q6
NH+qtEQPLzsm31bJgv6/cyFBYQtjVrGSH6A5S+RjrMCLkwvAI7G22q8ruUqqbFVV
FAguHwxEKqTKUfZMuo/tRTPs4szGteAnXRZFd89XblxwhTybTFKRm23NX1L9CWHr
RFVFz3Bsyzd5OjC6KZUWTmy4ZSaftBQjxtBRF9Fp/sGpWHwjaZc2zgzg4OKw+N5E
E7o3GVdX8NXbyGHxpEW/X16UapP/7yvz2GRMTXIYw16p0hiK+xvxrQ1wCQJA7j4m
OtEqkOL+U93jMG1fzWfm/9t7Ew27mCv9ExOW9vR+ss+JHVn4gu0OKrfoslFVujQR
maeJFBNDXTEO6LwmpTlsZa5ldO1/VYfjnRYSNKbb/lFBM4Yqb+8EhHtAw6X+fEwz
5YQK6NOdr2I0obavIb8bAwohPlifONV1oKwS7R92Q3A2YuiTcYSMw00soa7QtRPT
oubV39hfSRmJUoAA1aGkuYeTZcl4OmeAqi79CwtOXpKKs/jstzOYAJyajDd6yArV
rQkTcpZvv62gdFBk94G6BNcCb93eSG7+/Xs+hs5gSaHOfn4g1NY4wAPzvC5F/lpo
L6uHZNGTxKBlkiuQev6E3pM4ojk81zDoVTBQKfp0nGbBoBsg9gXfuqsB38/qpFnQ
zWE5wdIVlKtiZm3cO11IVup12W+Ggo0bswXd2SDNqXGRRpMJhLKoOuCoySK09+Uz
9XNV50rOXwZRsd3zTrlCYFsyf3GGljgziiNSodiiN1tux1p2n0Rc3LX9HKr18VHN
MNv5amSv8T63LrXqDv06U0wTsQTnJBJIeW5BlywYU0eTgkPuXkLXMJ3hI0sxVkKc
dejBe6wO0LIwhPWtSexzY3fMC4npBjut9tvj14YXcFIwxQ2/0xAdfG0eOODbc0KZ
X0uT6RuHKGzPy1v3lXpsg6tDEa6PAvUtCOlPEnKeD89+icyjqdkxyIARCPqic418
se6cl1lH2oED/eUtoull1Sd6WfHBrkJtHdTYIKpOZjBYcgzNY90vWf2FOlbnS7oM
glvknstWsumXqkMf+/AtTBC9R9W9U0kKp74GOetC63opcYeaCGpQLWigZR8lYUaD
GYWxvO2aTGKNOz6Rlm1pbwhFt+Un7s4siR6MdHuRHSBoGsQhsZuLxU01+zYMU1I4
6xSR26HfWzjEy5bRmI99oocYJjrGDRx7PI+LauPo8tEevtXuoxbBYOgdkeGQvgk/
k06UDfouMoF97zbJjCm0hvY3LV7MWpV6PhP2raZsktogOC7Md94pm71USxftkuPt
lTZwjJXK+oHgMMNDKV9fZiXbn3TOWp068wm+124OQGfjeBbWOYafCR0mGjje8uhs
P1ZDYhMqKCJHz8YbAuuuFjZUMJNT126YADFQW30+tuNNVXLzIhQsXcsZ0Yl4HkXN
97pWR839KZuzr4WFdtbD5v9FP1+3fzm5Jlbhtwuv3l/oYQ/YagivKJRBm9iGizxp
n1+phCK0zapNacb+h2pf5BvAnoi+oTOpwEu1Dh3380AEkxqaL5sieQJ2HCFOZD58
WDcXEphWbwUg3Gzn8Tco1CS0UNVOoXCFvuIkMFZ1LsEhwBChH1P3dGQuIylfmT47
2qsdqU9obJw7ue0+ynv8ndcaCTXTR0ZAlj4hHwWmQqu8itV8FS1mTm8Ris+vvGGf
GaTdZs5q8BIx4QgxhhR2zOjWKiESETNplajXbDEmMal68dXBRMTkB5VFN36YukmP
BuI7dZ2rEN6OJRAI8749y62tTWVbH2OynqR/FsMSxdAmmHtCvBciaDT8lUxI8a0j
cQzNy8SasvkiKbLowmRbioR+S/f8YRkfJexv/RBOl8w/MigSlPj3IrVxA3hIhtjU
tC6kenEqh7qvxh695Q0yUNQxkHk+JkEb606REx+qNnnK6SxBWZNExw0HeFH/vggX
j/MpHKbiLJfnRiH2wLjINsaPAtqALaPSVPvX86I0UoLVYNdgtbb33g1mc7HYGeMh
0tWAh7NB9BgiCegZQarY7c8+EKaKGRC4YXMyE28RGahqcwVQplYOxi7jId3mQbq/
JCRsNnGA+nrz1WpaS10Jbya+Yae1GFEcNVnTjzITSw3tFihqfA9U2vZKiYzwHlFn
JUgcVKoIj52Z3eyz0Tvk6Yrbirl/7m5iHSheIn8jd3jjVOztrOM6oA9UcU5+n8mk
Us64Zt8y1uu1XWi9gwJ+2IioHqdQnbkxovbtz2daSjeK8Fu2Xk0ixl/xPzAZEL/p
tdYk23AVJKkybe6Cknt60rrPILFpoLIWqcguC2WSVfsKQBdODC4+JULqjuw5Wtjv
GSWoSSlxBpePUEX+JB1L0GHrxlwnQtmoVvWAk9rl4dDgYg91ya3xswFbVp8xwqZ0
LsoaFdXdEuzubBJnhIUxK9yru/1lmqQVCdIAySKGeK5HpTCk+YnBs83228+qRpfV
1IE0Pry4pe48bHpVvyanzd6gdJo6JHDSTa9YwJ8/JzOEPdkQgEB7C20vRbMZeMYm
BB8RhyMI+5wvvkeOA94b9e4/6P6NsDU+/ZtsMDCVGJ4u3i3GWz6rfeJsGl4b1k10
oABJRnfHUBhvztM9WxhqO0RDRwCvsKXW/teFFivT8IEaiy0fmnfc/dEG4OFkm5t+
qwdxWJW7mcjdRXw6PxmtQ3/Gz44FdyA08nJ81Sv7sf0Fpiq23wi86CtXCJw3p8Ro
8Gff4gLvRp6+H6h4+75u05dW29kEW7ytOT5u2gksrdrLxhdA3RxvQvF76R8pS2oJ
gWtVNWRdjnzpcJDC6BRJvmFbJTn4Wn0ibd0k79pTruGMR7QpgaRuF4tDUPYK9oUI
8BRMNnRtEZJMcDL3F9OB2Hdk7hUKjyTBQQiVI1+gU0k1z4ogmZRhArdUcumtbRMI
3StbSt67Iw8wumG6Od/nOPry96oHbpIW7AROcXLqyihFo+15ostpI6ZofdBrohEB
yJaroHLNvQWuOPyrt/kPGRwI1PGkrj+MWH0xFLyQRcy60DgvkskwKmMrT9BuisLa
yUzCwxZM7jcKTPJf+mkPLvTzhGDQLwifGwTouPcYeO4JARrynsBJ0FZcylWdZxKb
yCxghAQ+OfbbEPLhZa2xAEFG1M5GxUFV95jCYWsfEFrv13n6Q6Vpqa0LUt+e1oZ6
EPPMIUp9yrbl3PTwLiJ1Ze1r8KY8sYWzN/eqWRHgPZxmQuW5xxLHokIl+kUYsSwY
Ko/+i0HYfei/ymulsoOUkMXC+7qgx1DhWJ9j/tQjvO9kXswAn+oumr52teiFfD+v
7CSInuH4mWG/g+jb/FqJYHvygNdXjtFj18J2Rm4eQCeVVX3LSoRxp4SbRKKF0BII
5KpwSDbtVFYW53dOPREEIyNikiGktE+VZa0LocM5kCeiu83Pl22eGTsk6Oe+quml
iyNnxW9hBvsB0rBLEV6+jcyEJOFe8m7rbEW+ztZS3u2n95SPEQXRKbRQGEtXtvuu
FjIkJCEufpT6Z2rDeut9LZ7Q85rSRkw9K/m/hCSzPP03K7Zp3/nJmmMxvJ4mW0Rf
IQX5W+YmPVfHw4ubeOWOnSWrploKu9xzHYlVSqs0u+2kW+JoUeQgQ4V7Ns9VkkM6
SVx2QugnTRPS0N4mb3TRS3dBgt2xy0kTtthySGPdqvruxW4AATzpS35ut/LBsROI
3A5myHcs0OEaYO/dRuyaswiE74ZEC4eTgBZF3R58eH3W1zlaOqd1uIjQcJhE25wM
lKwOaLzbraRXNQ1jQFAsUXQpK2qlBnqg/BnnWl6iVchfKRY5F0mw3Gqe8fkp2mDt
vhfRYc0+ns/YkiiySOyVXXmxRhKLRUp7cYcNgjSIlD8WAdT5XZGl7rg+E+mauC7b
Kobq/QLxG66LATiGGrGqiPZBEpSJjH6OupGnmWgUOFVJqSdMHX0StsXAt4px2EAQ
M6Elr2r8HzEiR7DBFgiz+r5ircs/QFbbooOVIVcIhYCsboYb/WwZvMyh6lm/75Pc
KUqZRRVqwZ3i+LMTlN8EdKzfRBYQBh/6mAWB3ib1EfHDPGAU5aINvRJwlRXY9kgr
qKNrVYAXl+W+ttQKy5i4o1+klXCr8OyetFyb1SaQ3EZc2+NJiu4xl+0GVVsngiAg
sVcrUm3fzrbUPVYE1wonKETnojnC/3pDyav4/UlL/AUmat1u3dW30fLVSWH9W75U
uD++ekvb+Tb0cUWali5SelX1CscGS2ZIfpdlY1Uz+ZExkDyqXTEuwmLbGf5VvsgS
AUSN2Z5Zz5PJOs3urL17KDxv3FL/cQA938RdRTjaKiOdUzmyATb5h9G6dy3lD4kW
LUro1Rc2BVx66VJj5/SFew+DH8FYkb9uB2ZqTX1VMuEEGOwb7XTeA88RdCqV8qVY
US7NESlEoTMhXkVn1+6ZUAueDe8WqIHf1rYXkOqhiZ6x0qBwQtauEaRrNFDDJxPl
D20d7Otg4NWTjMYk78gwCF0mnnXbnmvyIjiXwpOxlBXtUAuNvbEpwKgZmi9R+0ke
fCw6Z92I/wwqI8bZ1jWWsPm2IWx03/jDx2laLsyTCzY+LYioSXy0iXcWbR5h0d8h
DxHC50uJB8ElRva54kwVk9LT2AKfVBroVIhp0BGJ0pFwYLi8X8LmxES4J8ONKRre
G9a3EZclOHk5xIU1qPXVsScH7xOcCWzZjAkbaPx+y8jRs5WRLOO9MZjEQc1s2vQQ
ESd6Q/0M51CwHwcdDTqiKNW8+hZq2rEwhD1WsGD7+UYO30tkDyEa0/qTrmmPNSjY
2q8dkwUPcNPxrhu/QHoX4V/KPVE+GQjMLFgkUq0r3FbfnYcXd5l9064qFWCcqRbs
Lz/houAtAmymeyP9hgFnMPHJ5Y8O0+i+UxMH4UQemCdq+QwQ8t9SWWAsi9a/GFVX
cNVmOrJjtp5XjEA9KuH0fZzveI0sqjCNKuNsd9JqqXOO1NbD8NyJVdEBXTzOqMdv
LttGyz3ZcwFvfY6fJkxXQu/lpnLv9enMnGgBhzk6iCEOTe4cs8MuoucMqmkrlcR3
miyKOEzKa/8n9nC7poirqCZCjHtIHjJWS+h2zTdNeWs1CFgGSlJzm0fXUUjgMij5
AIdRI86x6yDaEVM33ZbsW6Ls5udtY/us2kEasyeLZ1QhOsPmXIuTEf0etfIKBtno
hEf4vxhEtsRYZtJohV78RplMaVp8xxqGM7u14GdeZrjEFcABKFMbxMuu9KEC/rVg
WxAqMySiPdM07RRLIqMxQhqsUolPr6zd/vKDyV4expnSOFmN4w/CckmSdL716KgV
7A8LEY0Wo+plupBKXH8OswD7p28JIG3XMBBeJCdJPbP5O/IwkMKNOhzmn5XVGoLM
gXogWxmhkdwz6Cyv+AlS0nuxkoJ+GteKsVPdv4jV+cnwa/2Uh6pKgLAnVpr5oKxj
39XIggxJNSKhHa8LIgBXX/TxBm48X3qGHYaYCD0F+3OB/0zSiBlE4463VF18pfRD
PiS6DKPLXU94nEwjzICqkOVeZv3pSR+Dr1GxxwSrQjDiVgOf+qQiloC9t0oFoyTt
S2zHppDIowbf8lmguO+pit3qiNOGTx7jIooXuvDAtPgXEagC5wJztAvQCJFLsr7T
yKXrhqLjcf1E4aKvpEemrW/xrVgc4WKiDeShTA/BgHlW3MdwkheQJKbs37ccq/hS
LhpyVNiopzEGfZ5tDcdck04OdiFeJF2+Uqk07ry417eJxflO2B/VYlAgtRNQbOk2
k9zg0R6jWUG6pFkfDrlBZ1qRetO3P20nRj7WjRAbTZxg8ac5qH9E/y2CP2QhLBbZ
ks/ypgwljlQPV0Q+QR1iqpRyff8SbUSwAGWycIA+0I0nhaw8XXq+7+4SCL2AxSjq
WTzUXMV/H9WFWzA2cnVka/x8cxkZ+CCVPc86aWTg7Fi3qOFUKzfOoKBanEp/32X4
zY6MLUMo/7hTO7mWN/VkgXl1FfuDagWD9/G+uKwkODcYiLE8JRPkdyeie7iajMae
FDhWz+jYVK/vS6o51czF9N5gg1Mki/lscbKvU2BtrOqp62HapvGX6b6Sh/Q1ViyE
5wkNESpb97hChndQhPvghU8yIDokQehHc6Hz6yQEcqMt1soUczhs4RTy67y48YB4
Y0SEvJ/K/y0lEx/sK1BSd3l91K7c8rG+ncKMhV7IdzeNNIRBuVpF0m7gEYzblDFN
0qb3020TGs1vyf2FH7GMfOpky2l9n3E1igjivnqo7nYCIOHX0uKsj7OSz2xq8X1k
gsDWdOYfh0KYtbq6CLuHnJEe1Xu353WL1VV1gOBqV04xNgZJ7sG0IJAt2LMUcVQF
jphsBmsfksMDkejKTRQIYpmoy4qBLK1pxwbkrR0U0ybM4n5qMrbcRzMKRR/L/cfB
kjVkVWBaLHxENgwDVEQoC0sCHbAVi6dPpSE4M0Wr30Nvh0mUWs3Vt3A9rJKasWfZ
WuoO8joy6yQ5Aor0RekUq2NX31sxbhcvOZNNYrodqj3RZOT1lhT2LXpQXtBI1yg3
OCxyeI+ZzPTVM5pGBPeEX6pd/D3Vv70Atp8b6rcaey0ji/lM0dxRuc3V2HHB5o/5
iIch0Xwdl1SfDTgrPaU0blOwq1bArgqayDaeF8pKlObTdplFnOBnOPqxJkNv20yt
C/AFB99tP2oaqgP/Ky4Freq6+T7mML9T10dhu8nUBrLMA/dR2Db8Et6O/KhRwxOA
XZCbMeRNgfN4BJ5hiAGx0HZrSv2GNrpCrAbXxnXBB09B+SwRPspHGC+6F3A/rRGI
0UUp/UKcywZGQLKDFR8lAdG02Rfe/sDr1uvinqlvGiiWqXbZOrbzwR3WMWV2TIQf
11zk44/9eMaUsqHa7oJ6mQRGXD6ICiA9m1/q+/dyz603urT4xaRxAqFOaxla1vq5
2JCMDngbg+AGQxS1OgPecItRcYo5hNc49mC74erNoEVMXk6ttzNCMUOdrgTM9+1w
3qvJoM2w2B9x9Q9d4pYZ2902dsNQ04RtmUgbOePhgER6A82Udv/EfnFi+/jAgssF
yJwIkVePM6LdT5zdqprz3I+5IKj3kjEHu+tF/4WtOSNiTOI9iICgjEB1iQmuRRBT
uSBfmh960skMORmxrsoiMRTYBxvBIS1xwoSSbgku5Mb+ar3JdIFrWxgAH1yDgeZt
vYyGYB3rKBXo1yEMAFlOmMm3gZTdNJLhqTUGJsazJF1AT8rBJcPQIB2LqVqJMOBO
UWaBPmoc8TtvIc0b6WSsAf6v9Sw50l93B4pHAiThTNvHYmYXEN9yAeKCDnObngAU
OJ3aZ9ClAWizBtzQ3lX0ttg8tpt2iJtBk8BBX9rGMJ3HS2i40bCqE1Hzq8fNezfC
mQWnjDWTI2EqM3MTK9zmdhvl3ZnY230RwNlcFWTPxrsrswVjQoNO360ArPCcz1B9
evrNGsx3DW15eHx65c4ES2a3ucCzz9iNM+ljSvGg0SVCnqT12oBM7M3qn+syouql
nKnQ71KaWUFvgnekKB5Mtj2wfIjgWl8iRyWAMrnRnL4cAICkcKaLSqpovZ3tueZw
kOAY5idqUzNauEi55lCl1CXUs/YMLGnKKoM5t3HNScuuM4FL6lOr+adHS83pnH7r
te07vV77BE/FwWIPTHOyrX2hHfYDsKK03+7SuHd33vk6f1wezaQIfgLB3mil0wAv
FPQOT7FyfuHfyVXRzNJMuSNehA+fh1hdwKRgSVn5aylBdLfYPpyJfl7GaCHD8dMs
97V2BEk1ZsJpm6azeRKj6TJsukTKY6HCVFKVwaqwV5+npCo4/MTeStfpV6NFjDKh
1I+uHxluxTfEpVh0HPMOSdriO2kIKIt/q28lopq55W4KsY67fC49xC+6alkYfsgr
NOukS3i0Zpjq9sR4ZLBNGVrYkXBKyh3EWm/ftDFLk4PShIh/b139ulAKpkh28Aix
GFr7v0Bs0nmpdpSWvKM89epTsgYPVedief0dTYWT0A0sf7mmsZCZbS3vXU2b8tMR
lPzAc0PdQw7M1cL6WR8D1BQXyN/YQApFXvnqVmJi5kzjKtd4+3N6EmkcNlFcwF/E
wN6jilClkrvsIKQ/rFasxPKJch3kzlSETsxZI/MWiubswohP0oFRDLKTPWriZMEi
Uq9ICdGMD/WNhYfGbrcRoka+0/IbseFmX098pPWX3akh+Xq6axvoSRkZN34t4hCk
N0xkHbPQGIMMcPwIClE4B2+7jf8qo4OgXhJolKpQKkLnGIrlHfqPyBszjCyKpHCC
KZcnDWzUUa9IRb3rMgpIwSMll2r+SWCWOvENKqw20ABaeppC8ZnqoFX35576blVw
nAqFLEsD9mpi1mzJNLgYuNe9RTz0bc5TLl8rSh2/3kCELQf1cgSdsZlf1NgevXkm
6Sow3qXW8FBfYNOD2wjIdWxn0E13zMrYxrv4/YHbea8jt2za/1STEpxEWR3ux00v
hwSVMyGC5bR5HPXZKoEgL24Pseu3VDX6LA6YRoSHNUGZlxXHcx4ueYUvbKgituHc
5IOsU/M7UCSStOtSLP2jE7P3u+Uw3S2nFnjmNfgfpaKXrGQSucznvDcEXoDG0Wgf
DmoS5lpJ20+CpeZBuTVfVfbd7zjd5YA3J6celeNrdxgZyeErq91auDxES31LnwmM
b91+HTpVPv0ifJoTmpn0X65er5UCe8FcKrbmp26DmmWooop6pokmc9V3QR+xPFl7
snwsPGGF2QpxySUkS1fM40KYjpFnKP2bZyCQlVA+Ihwp3SW2heLAgqUKccIqa0pL
q7xUpyowe9CUt1QTm90gZ1BaigVuWsIsFX1/OaNdWVbAvvjwoSeN8kFWuJBoP66W
+Zq6vVSXUR1FMH17usUGkaKO5fROnYAXFx2d31Jd/VJiafXfycFmHjtwbS/qZ0Di
AWF5V8k0fzo+uemPsyJm1PV+Qcr4ZJGTbAM+J+Mt7zX6lCKyhaaUMTs/R6aCLk4i
NfjL7dNWabusF6WTK1QNU5gy9lupNMj6dU+6a6DEua10wckq0DQuoOtSP7Y1vwQ/
wstQsj/z9BmzWRgu96jjTPC8VCgkACzmssCUfE8cnASFLWfmqhLWcCIGpxFMLMhc
qYlcFjBNnP/8xRx/1FsU5bqesoIA4FKyRYRPQVyJCy2nkkq86KI4VVh/cK5YZqVZ
1t6KxRwQUQkbtUXhMCnlBKfIaauFIctMN1gjetRAk/lcTamtmcNQRfBLrqqzb8lf
72ePVbSEFFl9LQoP9sYJoO96qcWunL5VuqGjBUZG2MZmbKeTroXzNLxEBM8d4ljw
PAp0YOUaN5f1M6bK4s+gSCU/ndWBpQv3muJ5ZfSCgATbTFsI8+dic42va5sZ8ijp
G1gy48FqDwPMV2NPMBTQHfHfAaSfCE/FBGW8BNUxJFmwHhO2LlJ0ue/vDxp7kGO7
PMCHpM2Eh05s2zIixIXeA7whz2ovu+KpjJJCAhibXfqWqzR6WhHqY5DnGd08zQdo
2jvzDVTSAADNzdhV2AEyR6L4KfGxJK5SikFukyXbGnCdoeeTX1V+S51uh1K66YtJ
cO1mPzNCUm4v5IrdVnsvCLqnXlhqxmwZ7PDYs2eJAGfjTxOnVeAW86G3EXwVOAwa
MCBTQWiNKGSTWIx2zWZp6fMTCWQ0U8RwikfGmZTqxO1um3Zne6tVIUs3i3rvuOgb
wX0x4hzkzyTS4JINqdjZ0uvMw/UWdIo9dUpNdYSIJWCZB/JaMm4lFnQ9OCoCXmNZ
HFn0YDbxVXRw0b42XpZVbXtxP9XrXLv6VE4eVGNh0qg/tx23qmExb5tuxS4II55k
Js0oah71DcRPpnJQbDulPs6HWuZTKza7C3AKWQ8EpesI1OKkjNQ6F7rV/MKThJoH
5EezRNOupuIAZL5cBkGYhjflqGWwNw5HFEjQ7szPrTn0f5YWizzDB0V55fOlb1Q1
MH85iG6tUmcF/cyrtjlAjQdttbvYvCdlBYFD71b3xCGnWcOQcNYuf6SJ7k2edZjA
Ga+sksHrIaY/npPb0D9dieIWQ1DKJkGhziZgBy6EuCAwarz5GjQNSNezrBlLlXiI
OP/noYLw6Qj8Gb8k8O2Ta1kyAuvKv6AB0Qc9g3LHN0J6MdP6BmOQm6a1eXVUTzuE
r/cRwYCDHL5J/2x463VLfifgSYlDW16TCrtEtLqDkLMv2sjFNmbpOsGW8/FK0Zju

`pragma protect end_protected
