// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
bLNF8fvtTko+h1l+OI/OmQcpvFE3FdJyCTvXBDaMxx61M4IhmtJh9ePkBff7
XXYT2OlZf9DHbTolmXZGTuigSLowchK9r7ADE+vqYPML7LW6mr9rF6eg5W9m
yKEOnCNysHe5nDWTAF2RkZb+LoO4zwgL25TdnbrfNcbWwOIYLS3TBDpAXQKR
tB4hn3bP+iW6DFO96c/PYlzSyFenEaOJ9TGbgELZXXrjCu2fPC/8+UUxmZU8
K0PSorU+qsshTKYyS+Lx4Lmm/77lYWKbzaQntByGy5fKyQOPZH+IrEzk0yfJ
FuvwcfRgpTdcmKaXo/NEI+RlbsE3AVYDDeMZ0Ngfyw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
qbo+nsBfddx07z9c+RVnHJCD8RkD6bZukcHb1UR6JuWEqkaMW+KI1z9stYR4
7abc7MXU62jJAx8t1nz7gYGXiSy/3l8YSlMTDJD7uzAsi/DA9TuSPLeA6OLf
LuA16bEktjDHAoQReKX6mgsAz3IxlGKaZFHTKj7ni6VaH407N98MXxguYya2
vzLboCLERRaUGguG4wXz1gHdi1qx3KKiu/Dk/PpvIkDYV8YnEmsEb2yzx73F
04+ozSLHYTTS7kaCpNck+0HD7+3U1foHm3+zE+KaPYQewlxILl8ICvjn4F86
aNOluHSA9IHwYsvHsNeRLibq+L0elM/HmsYJjVHmlA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
l2Jw0fBic8SoT9ey/Do/8EfXZErhuDwQSzQgFE+cY0yK+ydbPedLfxKXaKuk
WPI21Y5A12kgokKBt5JTwVjqNDXwbvHDAstolwMqDtOdgfkvZSrb+hCBRZ1v
Mpc1C09RhJjJxsnp5NIdPo0N6JxSqWMsEa1k/B8LvC8ikq/oqiUWihFxNOtv
AQKUOpL1PCRNuGgXdgywBf8hhlyg/11j0CU4B/52MusE8s+D0Z/2eMYz0cUe
LsEq2uTS7C8IPaKTbId5KDj36pVY0FPs/FXHtttIxdkkBc2dlG573EcQL+ZS
tu70919kpVVzWaOsWqUCU6K1oB0Vt3Wu9S7pOyBh1g==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
P+pWzmUmm4rK2MDjLKkeaiTzuJm9OZ0MdG/7YP232gqbcLv2HJWbNCfJ2oRP
Nv90FxXkn+bMCGRzx0Se8C59/1zKg9j+W49AkYuruRwP3o6BTfaldCdAt6Ll
WPiGjkyzVfaezR0Py9uXUbBBNwHj6EgTw40YxlKMyyBTo/z8V50=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
M4C9sLKJz4heW8O+4od8bNbXMd86NaCCSoS1s1Kvkt++TfVa7QFUmJie/SFm
BbToKvclHDZZCNQz/vcZ0U2mMz/95CNlak5Xt/AnW1PcGzIoWI7IUaXWjq5q
8rAdPdeM+Y07a4ag4XLDLu89NRZbIle316pGSdnU+K6qnFL+1dATge7fPL46
UQuz4zQoRDeJ+sYBPP0o3t6UCurJ3agbqUnXW4VoObUv6x5LPh2YhMyzXUgZ
sR7/nFxMSgsmEXNcpmvxdHHaTawK/MrQhOGjfPxHy6D/LM0xrTt0BZ4531QA
eaEMt/blNdgsQXHFcj/wlHEMPKvv+E8Jg+w+KWsid2xk4XMPUPDQUO9aiAig
wdW+VhSKQdXQOmcpZIRrFXX0yp2vJaojjinmnIoskALy+K5i4ZR1MsMf5Zfk
7Xb95Yse4yncNPP1Gf+QdyZzQTqE2emL03DM9x/71E9W8BRLrOqrWWg3EZlE
864GMzyRoAlEuAFZ6I1aXetGExG9byfm


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
uWNxXcdUrQgKBdLA7iWaTuIf/Wcrv+QFz+OY6BaRhFGJruZyc0jUhggTAeMa
MhQiXFbkHYfkzKo0wgYNqP3cBuGxU7uOY9JukiXyldqrG+mI/IE0OvBFwLyD
XGyimTq62OgQdhyk9GUhagBxMxt4jXwX8WFSTWWC04dA0IrEHX0=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
N+c41LsbS49V3LoKqbrJBoq+ZUJF1/RyUYNHhwHdZ7dDjGOoMZ2u4Mr5rk8J
zXuA7k3mSUp6gUR5gsKe7c9sBzuP8vLzL2pNVD8My6yDp6dntF7NJmfuxUBt
KsZo5XA/v3wRKxBrJYzyR0wIAQ1i5OQb7vhtBawHbHGuQSwHq6Q=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 72000)
`pragma protect data_block
cSVDKBIgFymI+WV1XAjq0kag6MtaMCj6p/1AAyUA9vgAfk0GkPapvO5So0SM
RVBGtasjzcp39WA8ovWm7xjPYYNPipEukLy/c42p3eJBJBM2sAEn9g0M2gS5
YTzd6B1T8DMSUL71jU+DhLgLeQxQwcD8VRYFpc0azHtWVe6OYQPDZZQUbgjS
mCa7LGUL6i0GFCz3gQvHR/2JHqUyR0gI+seEABRiUpW65umD0P0Fcyl6GC+O
0kV8NCWl9POO/FZlc/pgAgWL8aNgOtGKPl883VKzEAp90TbGzLCnxlekAY/9
HZrkDkQmd6zFrThmgwsBXuN8HN0sRFQ9/FXtj4v18YrtmuJvmQdhvYmITDlq
EVOGFt4nJ1rK4v36ZXpYfb98d90+vZrgwBHf3n1ge5YSQfp/1HSjdz2Reqfi
20esBpo9ZaEecRWlv74noJ4NU4xQJtuwM0D2vB7MvPoQuNuyFB3U3Lfq81VB
Ku6Tu9fN8YOfsuDjPp+uQwollnSy8FroRukB6ELWo2egan0UsF+adX76Axra
60wjvLf62juApdoa03rfKWB6l74J7dGElHn8JcOBqEY1pkX3q0Pja+gvIxFK
DqR08uZBMZ53Im9Ak3B73l1J68Ho2nTQsfd19BHJLdLJmsz8rDmMFlPuFKhn
UpJfKYJhTaqBZ+gP5PCFBjDS/utXb8RR1jt369dpRUdApS+H+4Y2fn2lzpW1
3eHA9hrhk0eaGqXpaQMDtXhnC9jlsHVDbm7ecI3+HC6XPbh5SkeOJmEAkJBk
9l5M6kcyCvnQdGyInlf2bLx7QLUJCtzarIfd/LqnYqA8SWdO8RpBCj1aKsU2
iDEJPuq4KB1/vgO7+DWjZ/LH4OqPIuVQvxMsOgD/lVlmv8UhVUoeNj1fQxa9
epyXhI9J+ZgVg718CMEmwt6I413ZVm/3/y5o6mTOWCYHYfym2jEX2hnT5reH
w3//Oefs5cgt2tjd6O3BuTwFUaMkWnqdGpNSe2YXUHWal91zV2a3evOwAEbi
eKFMosj11m9uuly/0zNOvgudqPl4m+6rxETGnF9MuWrlAOnca7cM6XfmelQ0
PkgJ8SphPN32sd40i+asLW2WdHYWe2NMzBKUK8P9AzSfRKMPgTj9ruiX9MY0
K/YBjiodssGexepbwK0PioXi8NNUOUK0l5i6zCz0fetKKaYsHbsaOhJNOIdX
SlPnV/djaY7HxMv1O9Js6urUPmDs5UDD1yVlANVNgCnHUtOUASJpSWdzJonm
gO/bFvyerr8WpIUM3JChEOimkZTvVXMQO7E7coxaXq9YpP0HjrtDJZMpXcUV
+kd1aGUxq7pvRzA5zTOTd1N8fX4x1z2A061IXPj1aATi5GAxhVIJzn7A0zJ3
wgsjDuFaFv1WjEqvtjZbbyKf1druel84eNzh3h+SX3+j9zX74I+GRWiKtLxl
LF5dGYRrdMo++DaVUVgaW14jH9WLK3cfwQ21CQc6vQiBm71PGoEjxBCBuQke
jy/M5672oGHjLUI9k/cz8fkN1fOxomFCroXdLe2HeZYZjUouPxMlGdVjjyH0
1AWMWI7ZsY55fhgVwkl+iyW6Hj+SRAUWRakLG3VHT65G7/wm696ijocg3jaR
Yt095GUpRlng3udosQLfdiz45FpQAWCR4DZsxEhtdlydp2L1kVYzemdmdFGt
gPX1o3nBmxo1rEwWzFikG72S6syKLQjRbscOuTC2t9TLMC7nl8WRuB2OyyIQ
6EvE0LoBr39dEn+GGNBhwjohVFt6AVbU/SBuli8yTQetxggIAO8Az6ZJhuYf
Yxjh7RubTftGxtawBFz/7jC6GTiFzfZAo/4oT/8crFE30Z1P2FB06zVRsigo
PZLdRBrj8P6dUvsuqjdpy+XhsEBD1FtVJFlb+xElC7cmdPAnlJv0VnBC9qKv
bjPyrQfDl9MPG3dQh6X6/pUugQ6mlPvOrN4ziSvINd+651zkC3H6U6K+/qDL
EpMB9NR1tiWbm30tPf3y/TaGpyfCSBiPHb/wNE/6JOSsBFaIVZY9WyXgh1hS
haUs5bomH5eRsxHxI8DRgB5Kr6TsqVhuQEd2IlTXok68Sz8O8wG0NWfyLd2l
Up/l8FuYO56sospoayr5cTUDgcVLS0C/NOTyO3lO3nHpiN1FNp6km/i+hIHM
53qe+lqFc1DkxxzwG/EQGQvG/2tnRuqWStV/HYb+GSZWiCGrecA5ODruKFam
hPDyx0bc3veHLlhDCjj+ReitRPGL0IgTVB9psLXXULRZOaIhAkl2sSt2v4is
fY289oqPzEfVXRYrnnpEZYSOisHDGs+xyscoR6ZR5sy7fZgyXC+tlYecyMyV
8jCoIUCGQgA72POuYr1KOfLOeORflBqK3DJnIexOaI6zVrO3UGF64YiTCo3f
69lIGo0LE4idEKsG5EMalQ7hH49WuLvgd45Wmqjlp/cqhXYSsqBzpHxS5iMc
ewpUpI8L4wU9yv7Hul2IboHGxLQjZJA5E30ipMzofb7j6tmvRpMnCTmetY6p
BVYtFRyrUSYlqSKTgwiefni04R/ribWwF7bSPh1ZeElb7kCCpKiEgF7HN6OR
EiKJHGoVbTJs2/mIfnOhfBme6QCbfE5kv5D5Vx4dIgOPX8J3KWwvoFPd16Fp
a4s5LiESE+DZs0ksV6o+9dVD8cgUudQbhBkF+XcKYYkQaaUXI3FGpbtvv7j3
gwNmpkXHCkUjKme5pABie/PUWzon60Rimkuviefwx8K84EPRkylqRmOMAySx
gDCetDUv5JH/FZ3QCxH+P14VYvNyJwgn0fAwumGPmozS2Ha2iRBw2Acx99lj
EOx+TvZBo9HWAY0+tIYXg0VFeJ38X2JdAKh46asZ76S13D9or7OEtFwbbqBx
aWMe1qacX5g594BqlKUWOF/vPpQTYiJUaaZ7U+BOmGcIyUhb6Wb/B+3zq4Uo
+WNTtg9sduaDsNoM2YWsqymg9Hoib50I9ShWHEw7KRtwlexMsYadFV1OT0RP
l/1iGY6BcLFFf27jJzoulvS1gMmwkg0DIPjwU4xX8xMxevT8VuAHPP25Kadi
AjlJJU4KWYYFjlaGGPL49I56yK/sBdDPc3ooUt4M5ZyU8j6iyyIUgolid79V
HithCvmPq6YI2hzUkYwaZHURKQPRIOEAUOKFfu/2e5H3pp3XsjMz9AqdK88y
oNmJxXb0Wyk3C7Ng6YUOsqjvGWaPqfyMtmAiFj9gypT3yiMyOsViXIIoboDt
hmCSnTf3ExuKwVdRdmZmMXLEjRrcIJVSSdLrFW+OQ1t2OoTGaf0s6G27bjZQ
nJVUu9oibaTFF7HetGFlzoq9J96b2Gy6gAxxZuuG08JXZWvlz8tzEMKjdlfs
PisAy9Lbn0M+3nCv+b4XQBNyXe1GHSHqnhhCPsKek4a8VkkDrdJ+vrJlA5DA
DYfZf7mVZXZ24iWYWRJT2LQqTzL/YfPLYCApiej8annNlJSE47Gv+QIPhYRX
TqSEw5SDe08p3CXsYYTEQ6aJbRjtMmJ2Bz2KztC4j5jKKp5ejjNXa72cBEuU
MheWJtUumQcj/NQeyzZVKdBX6LwAww0kGa4hzPZuJD6kj2c0X0JAtesdrLU6
o9gWoKob6oDOFcEpqGQ3bfb/jmiNWgh6PIOguMjWYTJd0g1/2OxqBInnEfmx
Hhe1jny81mxXYhhN5csg9Cq0UkeuCYsvEixmv1/bPa39/9kAg5z2vV1+7ATC
XwzKehg5f/qjgaacIRyuzltT6ICqnJCy+3nge73/2fkeuNvTBenZU6GfQM+t
Btj+lrUgyaFL3cWXMtzCRm4e7E9qng+XzWQJ0sI8oeRBP03MzaeUBaNVoLTN
KmtN9erThmy5ftaxwapaFqMx08nmYLpYd0pfqQTOy1OpeMhcWS4kXATkY8J1
R1AjNH3KBScm0JTmK01SbsMS/7rJtbPi3mkM26n+gykkRsUHu/pvONP0zvFZ
YhDlTV3/nGGOf/zO1Wufiaj7OSXB3o5Hgsipi5jbuGfF9CxWsHSot0VxyZ5G
IiKPKR+jjnvDvIymiPmWWg3VM5mv/X7rcXbe9T+rSdV7lHpQlSGZqyLQ+P/S
eOrZOiXBiAFHYs2487spy/Pza2pCDJO6zHsoD4yEdxCTlHYVZqzBHuTiJbO2
pWVyNyybDgXiRU/gPtxSksl4E7NPDjn489fds48a87YTleNR490Nos3ClG5P
7rT+5/nvzrHGTHtYyVac0dG+RdNVtXYvYBwVT94BEBTTLX8+RaDMHuoPEcix
ZfMSZg7WQEl3iZwcBBam83kpMNIxB9oMNTxWzvCdXo4qY9jV0WtkF5AAFtnf
MVazMc64Zj4q46oloSD2iGEqY66x/Ctb6TBLRRibuapYCssH9w9qfEwHpCCp
Iw4m7Z0mKYOgtMBAvidWA8ILCWxsaguO7+a6SK5YY6+k/dk63Pl/idZBly3D
aidGSz/Lqy196z1ptjZ/VJZ99wcvKQfZRC2IjsPpVvc2McbhB83MUFosx2Zm
nXW8wGebltxq24v7mLZUOz92O3IdG2eLbOsAm93geDuC1GE1/8cCMA3qrwF7
i4NIOH5bEKFs33TKaCVxwxeJYQ6hTrLDfZ9odTe0KhaGSPlimqXM0YdZVcud
g9BSDhQn1sFt9arHOcyMQfWiBsMI0/2q0tV3ZKdlrZ+Q2UhgKLQod9AfL3Ek
RcCFc5ybcF1QwL8O3T7EGzyZcAPL2cdnIxmjPJDe/GxIwh0kv/3Y3RQDKDF4
etEw+kIXGsVbfWecjeDnUony/QyPEO85bvG3RwLjQ0usAzCL31AyNZMjUmPM
hcJy20N5rSdiqTO9mH02USbjT/Dn/IEuGiAtetq5LRip8eQDcntSnfFHCnkj
rMhE7lgzBlan4YLkppGHWqWuYnD2/p01sR2t4vP8d9LWbxFNJdzCOPYArHEw
eD/Jpq0YTU+yQWeusharLltcXhJTOjz/hrtPJNO95deVGHNybClNsdM3/4wp
S4xMseBrYURsMFtY9yCTpa6KmZxEKEcVCyYzzCiHJx2Cja5J+AtDFrdGB4Q5
2BNLHVZjZGPCzLDyYY4ThQw4/3F9QWirTmrdzvRFMXI0M2T7ghXlZT//mN3U
YBvPn5c0k203hxX9zSRP9/beeO0PXoJO7yv2ydrEH8E70ov0W3tXrG0Xmoji
myxaCY8AzSGI/ga0mFTBHGX4vLIdwHITYZPJdEXJudylOJksOLL0Kys39Rts
GuxhKMew3IjJo2QmjZ9ahllIvCgANyezvhxlVVlJR8X4iajVZ2fn3lLbtFiO
W4qeCiMkZsJMyzy9NpNyoWTJT3cZRs1uCEfGOltjhlF/8uEiBU5M8qAlic6S
Pdlw2PEv+LLku4TMlPm5cK8dXVftlQxHDciCJK0nMDEC3DaSHeZ2n3fqg0qG
72IQaQOEqM5nK1NSdqzx9BIorMXuLIXBPNE+c/h44eBf3ja/r8zopzSsxl+2
8IgpwiIBRtV3JeaYZjqaMtHBidKlPa8xYIO4t3BKrvGVuiUBOlbPXr0TevmE
gW9WSs+nzZBGftCxU7Q9axXW0TRjoAr2e86oITQkJ8w/FPUnT/0ms5J139TV
pGxjToAiD5AyxUOpgxSJ+oT7MTG9SU9mwDUt7MWJpQh9OCqmAuXmAK5Dot5+
6mY7FKTLDGrOj0TPLLKOLleZjMq0UunxNPpXxyj7pnWpV57b0i0Mq2MnxY16
AY4Y2nfrYb63829gmu4m2m4nsG1IkFQsINTqodSQVEbuoc05eGjR51Sg2Mw+
z7EdAtLGGYFoMyxQdNfZCk2/WUXkIUg6uk1U2apYi9ybxOcllLWEhyz302VL
O+82O6COlwyjldpvyahAxcOO6DPy8M/oH47vr6gZG7ZpFPUffPsaMABp0+jq
zqOVWJJtapMTB91CRf7HNjo2SNo8S4xYstp+jK/+AoTJEsmxYIAzJV2Ab3gR
Il5Wl1o3YyMHrU4oX6x1Y+O2mZSfSIhYxmhn1XsH2rRYGoSwfc71faVP3Ecj
YmZcWiOC7AlCp0veD0XxXB9BOqy+n8NQKwdwY8cgiN1cwaMbg8v/J+KI902E
DT1RK1hxDNKVDmVGA7s91Wsub4ULs44/OZjLf4lTVvKWNHhbNg6ewTdvL65x
LD5GSRqFr+fY7xZAShOKpMyh+iy/NotZLYwVfl/r5kiGxgzae0rnCtKI3kfa
pD/Uf1g1wES0CPHPmYlpZJ96jD+ArRnxeoBjEkpREoebQfqJeHRK/+TfPu83
MJ58O9Sh/ViUPRT84X++wlIC6B7vvY5cfauMkgVTOZnUq/gwRF0AxhyrVvy/
vJMBzSCxzc1R6tSUSqgGgCPMhNRPqaR/UCGk/9eGtx9bYjs83giD7a/+uwsZ
HtU/6SkvY7v+nXawP2VI/kGH/wwn1HzONni26nkCBa4JWtr6TBmFO/Lsuniu
F8Mwyjf1GgVRCoSnh2Xf+RIgFPYjQyZJFLiAioDIIxEOln9ht7XEGHBzzmPm
Sa9VzsrAeN0QtHPiLKHaOxsfo2/xgjSXMfRdRC+mKzIlG+P/kdJUY/22HdoL
I6ckvE6noaf7ZnHsryzIC3eYLJWC1ndgtkrsntgajdukl0tVLA4ci7EhJcbO
gRgtg3+2x9rH4SyOYQ42ScFelmqioQrOYq3VZqj3AdDw/IXkFfN4CWeVz7SZ
OQedpYiuFyipMoulP4TSYFj/oCVZDhbcwFqOvcNjsVMklRHfHQyqFjqY1nhu
jq325w3FuM8lxww/3B5cW4M9GoArXMVnq24ExvV6RQe7UDKeMaNPdeCwSNT5
q011gYW1bV9OfSzzIX597M5ON71IcWZFSxj74PIeclN24/y+H/iLTg549K88
r2oXYrhTqrgbCNYbNv3OITbHAvbpxdfbd9aqKSzDtHeLbwFLu91Ril9G8ROI
S00E7ubcDQB6NP1Om6+LhvMyDNjNQ/l6I5mn7FLzuwGuk9GO1zOINtvHMG5F
5yqyZkZXPFp+IAqZOypG108CaCtfFkQ8iSAxXilVNr82Qlq+YVT3ppxO46hR
qR6TMFVSAJKF7wUNpeW3Swi+B1EqHJDd+H61s33bJpWAQItmyBiQIL+2NQSU
mKtCLvSWlZCvmIjseKaYwAzzHX22KIQ1g3pehM9eJCRgwZy4g5UOeIPgc3o9
3ognBsin72c9wXhrylBg1l4Nme+6TOJpw2INH/OqanntC6f6iw9jiRYbnnIh
kTn35gOFrIyJuE0NMkv7/ouNxAzo/JrYxW7nydjkqwd9v/EO1OIzYQIvxHyF
cwSMeiXEJdoqcC1m0ABSZ+IV/LrX2cC1F9LTMQqoXInaYjwy7n8AG99YZnSq
nVm82fSR5vIAJ12pVih15uov7EYsITB4H9WmaVsxATRdoaIf3YhGaNnuDYO9
o4kgQ3Eg71duvdgqXgR/2MPjGmAXBFPgWzXtLAAOYHKtKjCVRhuB3osUhgI0
l5EiQT3ZZ2CSmmCg+64kiyqsyzSLmVCeyFeKmraIwmpJWy+6oitHYVhV9ay9
ZHoz6SXnC5oz7vlFr6tMYl8kSeNEOqeia8u63v3RiJPuaZhtPNr+Q9gadPF3
8sxZ5XwWzQtNPklBps1GSLUkGNGRbXN6LP8DulWzsNGOojBINe5/agY3HQCQ
7YsirtfWB/1Hw6iKASrtObIu6DUfAOAkIM8+sn0jzAmC/4NtZnl9iWj1cO1p
y8I/iwnUQYwkkcnkg60tLQwPArqadEKpNhYPHAHHuhuEZDmFVFWM9R691LXe
J6imh+lwivN5Di1nWtQyNJn49D5giv4PotxcLP/q0eceQk3wuNZrGguG3mWG
EUWhwNDEyHmtf1Fr8Nx2bMTGVrzlYYIR9q2/JfexiZf+yXRmRJ0l+SPlwvpj
wBMgpBr3FyGmm/bqph5FEDttLMvPcNqIPW+aCVerU6tEJkxp/O5agBkkkpAQ
8WWLHznUExaecHH6wJSuOqde3jazrI1Xs7dKvTNglAhXlwDAHFqRaMbwQ+FZ
YfHKG6StEGdnRuW+adKP7zb6QilpuILssTgwe/gQWQdWuoNQPOcj3j+u/NUE
SlE8R++KkZXh+y7K2OiViH70R+FqGFVsnqIH4xi1XTyVk6Wd3QJcYOdG5vqP
wOk5X7H1ABz47Y61ke1HSvGrvP5aAK1OQpRa5og1xJQ8aDBYyDlIn3zr7Y1/
IwVz+aLLxIVCk4vx8z+LUvk+sGrs1lWOEWNsqeJlDPd2McWQoHMldz9nDjU9
jFp3lCrw3gneGGCEkrJXwQCgogHg00/RVyRdRrARvqLCGm6RbLeBLSfNXfS6
IpRMIEnRHl7v7iHfgvAO3xfHTPod6hcn/nHBnaC6ZjF36nH9GjmDRhAfg5v/
hYFWjY1OgJikG5o0iRHX9642+/0ZffuUcqG02y09J1yzJuNQx7aJdvhjMl0t
d+jtDP2M/Oc6ybsm22GoezPPpzti4AykyfNQdRPBKZ7u5l4KMQri9h927FgW
teaaw/K/dIuKg1LwatXg8CGodGv3+Xxz/4mLoCaXl82cJvqJO9WbH0cRYepA
6SeMM8/NNNCmrEBr4kV9bY+aWwqxthuX2JEFxWEJMLFUvZMrihTS/ScB09aI
i1A8huCiE7HVFECmOxg2iIIy3Q0AvGYxEDiZJx/xFzOyFoT3WTjlwJ2jeHMQ
PabL4Wx/HYuR5LXo6pbIiSdlxxgJkKmE0Ga/472c2eWPJUD4rVMqMZqgzZHd
vgbQNlPnL9d3XvfwB6ZIarbEGLv9hMvRhAsBTIxHYqb2EYXCXeLcKJmr45tx
s5ZcwcWCEQ7zDLRpU892ed3Uq4tsHrawdQbMgM7Zn8tk3T/SoIxiMdCoGNaF
Bdy0FJFNWFn9iTIlA8L3WW+bzhKYxboUE3WbP2NKivYNuYZutor01ShQOUJb
Ms7jRoRTHm7MNnNdCdXhV8B+MNX9HI7Mhg4U4oH1OUvvwpFPJKbY3DRc4eg5
aKdqBpqsMM25wSv5+YQdHqnZJ4aJy/z/833if0feRYYlKgBhDt3xejaY15J3
yqLHzE6Ztm8cQopa3i3aAKcTP18vstxhxaxJmh8KPXlEyl9wyOkgGL94W/Ar
dWJQTNIMpJad2LOUryhbh3HZwmWyJ4erJ3GVj+5dL4H8q3kzQ7nxGN1m9LgQ
+76x4wNuIQl8vbPup7Taz6vSwRpDq871XIV8OMowVUSKdgEgJ0BT2hL4Zvue
/P7D8yFPtjqQG9pcuVVvIVTl4eN+yGI5e8JJyPf6oANMXW9VUT38s6yFqcDU
KvKQOktDU82vFY/cjwYpVC8Yt0Y/SXzhz71FRPp7TRT8NrwXy9yymfhBCNFT
rjWkka4xvbVf/jswgMe5bapsRpETWOR/4fCgXpT3pph/D4/1PiBJwxwVkwdU
Vl2ADs0r/ZW7lgPkyV8EOf7foib4ndppUVB5cnv395aRzKnjBeK2gVQcZAlV
IMYY/ftcZTbFld7TtKMU7ffOacU/SfKpxb2KJnWbdgy5emC2o8S1JtZcmIkl
0rsycRbJlnEMoP80McABBaTpA7UbmhRMh4PEp38W456kUYXJ5tl0b5AiNdLd
QimznfGsya7OGhTDcHsjKkiWyI6PRZwq+ynHJbdDLwe1Vri0ufwbKk/zVVB+
2+j9vR+uuNGYkxzGb9oozUZVRLNtiMrgjeaJY848JOt+KTHY4YoB6Bw4H8qA
Y1Rsj3v7LPHkrWnsvThr7lXk8cXbEOx7mpkhUCAJWXGXhpNaec9UNG8q3FsR
bc9l/DWzXYgr4W8Tq8D1v9anQvFVsltn3mg3xynEUPOVHj3SZucRYtwB0lZ5
yiyL2eOflKBEpg45zVN4N3gD4RDgYtelSqNV2Khk2ZjojMXqaKoHGmY9igyj
4ffjrpmZH0uMk2w6E+V7WeEv4ZgCniCouOMJ/gSmEkCxEcC4IwUxzRTebrzL
cM1mK6wjSeaTnu3c+2aZ3qCl8ezHwzbxoC4uWxnhyGYCoZYHgEnP8WYRubjD
KzA34XyEyQlUKER8dGsBcbA29XYpzu4cDAJNiIYiFUqr1H1EK7fwVI/5jv9E
64EJv6TEuE/PowISgxudLzfWK51/TNOpq8Jl+T4zZ6R72mBVRBIfrpKoEsNb
lggEhWbZy2zqyYlKxh95XJ7Ts0psZbREicrMkCBVpZJTPMlVPNhIwxLlvk7W
7dOdvt6N78oMz/pjIz2RE/qbqbkPabie1uVTLpkLdnvm2fYjAutp+G+rU2UZ
XO77+eHQEV0QoCZnxb9g7fWnCy1z3WJCALIGqvC6jrwDlJV3WGdBsXCHp47D
sWwZcXPcwt6PEfihp9FRuI/T4onApYKJQo5scASYZy6eEm07w03lltQ6dx2X
+tFXN/qQkP8VjMNOQD/3D1Vbi/E5kC52AP8+cPgffqu8c9GLKkevAx1W4zmP
QjsQifb2jMWFawOmBb80tqGOPRo0AkwsEzhNUmjb3P60ukRo97tgIukF1VQY
+RFfIZpC2kZT4hV9tPsJoNduqLl4q+JcsBYPzh6HI/p15Qiob8ZEJ7BPHC8h
K/YZ4Jw6OH0I/S7JC0OTK9dsqwciSUIY/Sjf1wzZDTZFD15ieE1nuveQ37g5
anXfOa16ShmaUIseESVwIfgByFT5RFdKS9LLW63lHFsKMFp5HEnGkAUwzFNz
q2DY3orN0hzzLiBS9bXj3dz35dTvkzLsIRh95ws+O+q4QJSXPGVI4UPpcsin
sr/ih71HlDQ0rZxSrKvo3tpXbgpzD48XsRaO9LwmiHEQLNf8nMRYpVHsaHBS
tLSavfjPFh+a72wDvbvyemNGn51+1Sl/hjtUCXRCjP4kxv1idivWfde4ke84
2kGDO65vEJMUjmASPlCUokmLFww6xL+j24q7rhTy7EaZtO2soG0pUe/IYJW0
49rRuavB3l1UCRf0WZ39ISG7zR0CPDs4fjUvsLsUui8kkBNmu7aY1wNcfp3W
40K5K/Rv728qIcAQ+JhMzOQTxeQ/23Xxljei0kPH8UGTrbyqpM4OyfIZO85N
CWstgsykwXeqDPrqP0Ne/kc6IpV4450GA67/+T1cV6ChIJJOy65P2jV5I8aH
hUbAfYoJrzAnO5TSvNQ5CDnJyCLTu9KDsbQTtCn/4Th8j4fGHpE1mNbS60Ad
9k39MdfiktTu+f90LeJ4TNZy8/m2NrVNAzl7yQuhMfJf1xW7de2L2T/zivzQ
XXbcjZxb1KP1EPOQjdwSt36fmHH6iecjv6agHnFnNDtmtXFO9MPj0ZRcp2Ah
AQ8eRfX4DhEW6ArKlJMyEv4BVy31IkS83Xmb9Ae68wi769zAlgfB58l3Evwd
7zVnAU2Ug9rGn1vwTtmkqSJTdlP7tScvZfjF3/Dqlr8QvYCiZPFXQxvhiLrG
fcAIMB0Bmd7xMo54+LidzpWUUdhS9QMn0TYt+w8NfLzq7d2BQ517L62uAFSJ
yp0JFyJw/J6RSyAF4gpFw4DVdeOTZaEQIiM5BfztgQmqDq37hdFC45zpzyf0
qYNnoGH/EWXZdRC3vaTnk2dUTvB4pyetsxy0dxH/eAyYMPCG4Q/FVQmyQW6c
6VTFJElb1vh95+gBFuVioEf1OhneCzjZirySJebK5l0F/JrXk6RCud8UqoS7
Ei66082jhB04KWwOGvRJbfJadO2b5Fsb9YcQPRgk73fJIbHSMFpGjUJJm1kV
2IlBRzzTH4nn74Ge3HkPD5ol/2wLgRpZtYGkJzaS3eK+2FlDTgu5XPk3opD+
zG9EBJw5Ne+AkGfHAaLpxMEMSVMWsDwp0bqClcKKt9rG21HZlPp3dOMx8lWx
F6Btgqx5EthtYT1nZfA0ftK+TfilBxms53nav0xYW8EurvNDmCMyUl7Xh63t
mlTPvuM0mgmeFgB5EwDFYI66KiALZ5BQhOSfMfMSIQx9wAi+VrjbpZrrX2fR
qlsROBHWD4ZIWMEXi2ogDJRw7RJwLux4YmaB09SC/1rblDkZlp6TuWcp/Kvv
U4uNDLhYk4Me5BxhCQfBtZVgCcm9Txbd0xQ94I4AN9I5BH+KUAMUR8Q+qdYl
9AMrNRkEvrRHAGsDsSjrCBrkTDe1U1fWFj+jOhchjEZQCxzqTaC6LQqqbwQH
KWci57m7ZleGnBa5A301Amh8fmjGyHzptaSuverfzSMZLvAVD03E3YDSmGab
ydDAMVRdyLD6RJwnheehnI3GnPLQP1IJB+mmA0hTx/0I5qaJA5DLxgnEKaw+
8AcX1Go44x5kI4Szr+7R81jinyb4z7x2fihjEpYtd79zFRYi/qYnEw7q34yS
dea14l97xc3VddZdZI0eO43qAdldrTMbGnPDaV+bEpzN98JYR98UjbOcBUm8
I7OJZkLLPadCL8MMjFleJzFbFiP5ROw1C/yzqIUWHvuLajB8pb/Qdc6BtYwS
wOJiI1ZhiqsSWL2pDfEkTVjq0lw62wCJJ1yjezmSwnkfJQiiEVifTXRmGhjw
uuv9maha1PKLmQrpAufRMgWHowypB9pgW9aw3MAuSbx+pigw+pyaLnmt4ZW2
hOzI6SNBmCa5pmo2WCR+LDyMGdzkMJ7cvaQLKLNn/RHHHfORNIaVxnxqKyL6
92y1xKhcVZfOcU6wPgY3oK+KK4DxdKm4tL3370COa1gklc3hKgQkeAbiVd4j
p6OXofh0SxLHTjD9WaL7d2BHJL1/Jlv1EtzAiLKgetpWJlL5D4Rsoefzyq4B
fZzyNEMpwX4AqlLNwqCFG2BQe3Pl2sZ1EsRId3NtzLehr4CUI46nGH6UXEeu
db5XtB3PlIpSoyQBKXznpbdz3QqWiiIVzHsUNlAq8QJ7QOn5Z+XG97w7/7NU
IFqYnka7+nIWdhSh8/BRZRAf8ogNQqE9Cy5eOel0380IGlwvOpg7FytIDRFG
/zOnxS3PGNfEurBGTVH4JO/H0a5OYpUG9R2DV94tsIdZk2IfIEhnFWCtraQA
ImZaNQJpfPgd5IXzf3wTpOoyziBg3VRGlN6Gp4Qc86crgzUfxm8ffHBMgR/p
P0yGKpqTUhUJxuzBjBlKiX3Cpnwqoe19qYeIW6/YoVeizKCBA6mUR0aCS79E
ohD9I6Yw0VCCZoLyVUxqQx7G9jpK1utJDfhhDW70GSjKsh1BzBcpKBnwTjzs
2g61U69YawvdRkrNLtlMyH0+TvPX75FBOJHIcn8EY8xuG/h8oT9elVa3dVsA
6yROPWOyl5+9qr1rgn0/pgXYlD4058e6GmMKK1tqcUH2B2c2fhSu37UF9sE3
J95pnpvFu/rTVt50KgUgfIFPZoJcpx70rtn4YlEax1xC6nSp21mzUqySPK//
p/C6i/tbcgDGB91cFK1NzvFm/ddouCaVYaTAjhRXLB2j7Gz2wcNf8kdAXQwu
Dm+iu0J12l1DOam0KhHXQNOdOhGPcWJvCS04441Oy0hsMj9Bipv2Tmi+A6No
h6PBnUjLKBtsLzZjCUHbiBBJHTJRakT4pQMAU30rGuuLDFE+DiF0ljsT28eD
9jyvQ1/6dAOZzouLlSLRINFMiHoqlvSFQAPoY3MphLawL8PPAIZtGiJVY6Lr
cY0KwjDpQVYpze0x0lk7tcRFOa6IX9Y2FTj0RHq/a3tn84RVUYxBjVoVfTl7
wQyAC4hyrIR/9ZSidOgsERpYZIgJnrsZlpjrbyQOzAFCbijnVmOM7S/OTdzo
SgXqQXJT75JHka8vxBUI9VtaFPNgG5k9tqQ8gQdxyNaE+gFHwlEOKnRvspfr
EWedR4n7mGFQZlJuYLn+jvo5tevuRDuWGMn7dPTllO34v4OQRu6zGbsrG4u7
cD3LDwKcE53E6Xg5aJuthoKhtWsybbcVpqqfuOAMyjSM/XkM0m2N1z1vg1V0
6cR0w32glfIgSD8mZoIctN2NqZ+FNFR0KdoNrqwXuPEfIp2BeqyP6sPCEZ8Y
g0gAbS7wOZu97BG8uyXOyPRM5NEHCbl/kr0zZRiUTAElRJijHwipYk2sCHVh
L9FiMK0DnTxzuIJx7t4hMoenyhBDgR+zIivn3QcBnfbdWxc+NUlP98CbANeE
OyOwE+DKvHx194iw42htlqXLFSAxOPesNwpId6l7ENtc47TElNF8iGRgu/c4
VIpOzWM7pcoMKJSWIeYIOaHvRGz0O9UwQwVMf/+Fwz8gTrV1b3aV+k7TeZGH
9l1ITK5Wtuy9Ic8H6dxTzync75DVZDNqyKlyV+zmu0IqreAcVzAcL5vp3q/8
CSVFbChdB4aqVV7BIL7snyEiKLMyfGs8PqskQihHijNh4Db0nAo4r00/ZDS+
rSf1wcVuqPsFqW4Cnmsswxtc9nk5O2B8fCdPNZJ39LNNeU+lWxucn8L45qtP
9w865rKVOnqwB+lYNPq6oItY2uhJTPFCaoqQr4oQz/MCsGI1lSVOgq1+gYAl
aN770Mfao4v1C7QO4ddw6uwvJDqM2V/8MuhfBNpZy/Jyh3hyco3ZwW1ntVaY
mPKXjLU9Go3xPO1EChJC2m+yT7+xCNmrHylDLsiCig/iRT10wZNJ+cOI825h
S2mlR8rrEehUeAnDsPwN4Ngyc6p3i9VzLj36s8qS9VA2jO+J7xDr26jPmn7g
1nlr9mBLkdYAyQcP3t64gHDloXJCMGEEdpZtuKqqdrpzX8kiIlOiDj8e3sZy
nvaUvs6v8az7YAARKyKeW3odbSG80RykiX1iUZu/b3bSH60FAJyyWsYtr6TT
p2ZQvGWkz34M4lyDer+BIl3Ncd0M9GsYOAxFc8W9yBN2GZC24Cy5GvFObCJ7
yeCO66JOv6uVwJBcHxw8eXuXHweG+/GayVq/jSbqlo5C3ujC1GRb7DYBSPx9
pAQoP8awnCyuvtkyXnd3XXbsN5IioD9e7XFVr5PVa1zxVNsh/O3C17QBBPu4
FENV0hrR9ujYdXARlx8nWRIXxwyzT7+FYY67GohN8sroOySabHLg0iEtWaEI
7RUt5iDrDCq1QRMJUb2azk70r9tMHgFQY5Wd73zoRo1w07sNXBtZtH8m8dIP
ALkyvbELzp7ofnFi3p5zerZ/TiuYAqRj/5Exz8jPvPgsxoGaAQrqp+vXIYi+
w/J3r9sWWqa5WUZuEiXM5/WZqPOehUBzmBQRFw3qlzaxYiJpWNth3vLk8EIk
HQ0x5VB0mF8yOhoxhxzxjeaAkKWa6voL1qQ0iV7xchMN5gSK4q84PwNpAW7h
CkL4UrA/96HjAMSTvPTdElC/fz4PB1jK1AtmlSCxaD6pxEp7RGw3UJ/m+gR3
CGu94X29BIzU0hrHYBLmaiw0wBaUqKknMYMF2o1ZpJqkypFgvqXgrrf6FPYO
6V8D8FyeZGMV4FXIXe3QyS/3t7sOzxPLhj9pDhDuMtGS/JPi6cY/QPEmKIX7
l6ImKxNCNuYcNVM2cENfbMV/gFb3X5ntoZ0ldZ8n0J801Y0eAER0OK2Maa8a
sH//mNFqYtrhJVdpVK8Ed5RZjXiDKVpPNTs59gf/8lRrBhLmZgnzXEyWZg4b
/NzNUrr8jtDtpUJqlMm50afv7IRvdxjR3S799Ze9UVKraXmMHYeU6DAdvgAF
cCwdp5wexKSSVFAkciSDntI15ihlPZ5m1rQuHtBZ/xEDAdPvXaG4rQVPoDq4
sWmcm1m/qrjdC2RPg7TH0qXcCF1Pe/X8sDH43bsWUx9hsPkspauzBM84KahE
RE894xecXOG/ngGvG1rmMJri8NPNTZ+oVg6UBk0Kh1Qkr03XY5yqhU7oVIn3
pB10I2BjJujIwIxQfQ0UeVWiF6Yg/XJYdbV/ASn+t6RlRIiMdJufqshi86zQ
4AEX083VMxeUJ42er1pAWz5oicAFRfAoJX8IQ45At+LhlftfweWIN8wkR+I9
wJaq6GqNyfUN+xichHKy9ClnEQwuN3fZnp8wbn6Y2cqjl2ZwI5Y6S6UbNmeu
qsZaFR+OqXpVisBmcb2E05WIdtI4BKzEeznhnjo8lDjPtXYxMBKGr4G8dFXh
+GHl1nnQFhwyPr8ZYDgaaZdfQuthRpHw2ve5gZP6RpsRlrlCLWOSIhY8GyEo
PB526Uyuwql0GzAoCeT0GDtqA66YZFNU/NKG3bPmwEZOKNp7Jnj3Cgpz09Ol
KfRTMsGIllihJRu6Uk9etnmxLNKF5vZ298DUIiOZ+hEjap0Wl46V2mNqLRSw
Ht85Eq542NMyZY+KMa/o5ocVxafuI0jbf3FyLS6wr794+d3pkpzZLBlRRAOk
WGXZ1h0o4U4ZeOqtmfEB4DOOijRdeZ9CL9YTrnrv91/8aj7kv2Az5xelCZVJ
ruPWkdOf9yccpQw4gRvygoFZjK0rLIjeq0d7jFloZXKcbvgkw3dJAFjdCMG5
zuoh0dnQCcm81GTYCgJvn8d6teaMxAjDDs5pcSNR8cjpE52KIvm0I5knGM4s
aaVMBsPNYvBDq7StwrpOnAdORI/jHgh5kelu6xfy+vsJ7HnDqCor+YCQ2DD8
e24iJjS1TOc0pmv9Rm3wyGvgFXb+tmWarf5cSpjVMYkLrf2M+VK/96/ExAOX
0/SHitCiaOjVgfekkAibkoH1NuPmK7XG0Rv0izdY0tuzavqjbOnbzFPjVLGi
L7PLCkigR8SDtH2bcF5Wxa6qKSbg3mgnVXhkX6RjbL6sE/HuNlXul2iWt6yf
yGRoc7ALMd9ZbN1xQPYqitck/KxwElvRy2ZIxbhhoqK0rDCjFQ6yUBkUPkAU
JXew8kOKzSSJtYHU5uhqx1MJ1rg3atifptCujxkCO8XIHOMRJ/Tz5L6om/CB
az4wzxtbHG839CAAP9K8ugtUEIdHyPZMTLOvDlnYP1VipfCxmQ9LWZ8HAhxA
VnPhnW02MiA/Flo6diqm1/PRL5GwoUfu0+3debJFaWLkzTqjSCdXTfXkFKOZ
LU8uBJ3ACoGSxdh9OQt1ykNnlESc5KW14h/oRN+M8VPGp8UsuB9e8AjA/X/W
JGwecr6irJa3L11BXj3JCXe4uuWXhaCZ1nPwMvFhLvf2AoFxyTcBWOLYSI/k
IEDR7pyvy9yXiZDUNcxAjSZnP6K89v1WYUiIAr8xQLJK8ZpCJnKC+iOCCowK
3LoAi/CAWYp1DlrbK+KuqQXHBUo4RSU9P1mGXWmR4f21EuykL8meZYSjwdjs
hXMFg3hIfwX0dZumwRIrYUkn/AoHOgOMSB852MPjHuSnDiiX73lQKfl78zhJ
j1iH82QRGa2KXl+nrDjYYe0IXQKSyjVW1pu+3GQPMAvGJPsXTltmQY6z+f2g
oUJJz2B06J/6bsLecVWrQJU5B2u6SjRXi2iJA/ArZWCVj0ZKu72RH7ETJ1X2
HiBh1473N41N+h0oONEeaUUxBkhA4l4VuqNha5cmi9tp98K2XAnqP0lM0tsQ
7rur27UKWsz09h3rbijnnNz5xzXFe1wwnJWz74SNnIhecMhzPB/c6v5P2fsS
bt9VE6URN5Ik476acfLJpOmTsviRnpmYahCiKzw1aFBTbvedW092frP4svyi
DUk2jurDf731+5sHbK2oYOKWNxYpYxeOKBdFFNrQYJv2U8p4se8wdeiirC9H
4KD1BCaGfvVTaNm7emh+JrGSkV1OqVHc8FQWH2fDcD1XrrDffNXnzqN1p+VY
VnWosWFy5j2wvjy0hZlw1DGpj/6m3vRTDoWNDLc3B3uaPZp6DOCTBwCsbRKU
ZByvFgFwSl+0IrSqIcxU/+JflKIu4sraDd1BgckP6PAU6fbDlUK2ZDeSsBOK
Drnqzy+0alHGxMNYe3tcnEO/s+LKSewUa056T3URj7qrAhK2Dc28k/C0XaC0
20IAcuKywZ1jJwraYdGo1YIem+dk6UkcJvyyUuwZksFgI0EQ4Cx6Ol+ffg7v
dol9qhyugSLTvOi18cDvAC43bJeNIx0jWHaOu9vwFpj6ldQ8kWNmQ1ZnbJSo
AfeyHXJYfVAXB+1YXaolQggqTpFLzXPyUDQ2nqffUu54KJBOuZcdvfEZByua
ZVKuGIAgqqTv6p//BvIYDkyKnkR0BKAFw1Q3zYlcAjoGTuYBF/S1xiZEXM4q
6HvpGgyosNJDDIZjyv9ZtCzWZMjBidbCYD+/kOZ8GsnDxmkre5xopPbMZLTp
fiBlDPkGhYzTQZZBAo5VlHIHC9f5A2PcwKyus4frh254c1PsTGo4ghhqh/14
Mw/n8KAPu7+YZtyH5JJQIWnbuHBLLFObnceKIyzePT/RvREr6Zz6VhHiZTXz
sxnSMi7jKTbXyUNRby5gWi6qDLuBltbX2r8ZV/e1juVueforJIQpBrLzglqH
VTr56Eom86VDWr8RSLLPzYClN7OTPelhE/Ne7dUsvSrhcVzVdyCIzl0/mmDd
aWlJeY1XlLhKeadmzwwKKjdS08fhJ6+JvHW/CyWt2VRUNivxnSxk252KYj1w
rD8spC7Jk3b6my7CKRKQLufdPUaF79k1txiTqh2FWM7FlpkVjlj8eNqpMOUL
cZ6NM7XnBqLPP4KUErB4hLGyqOCvXWxKWZci7DfXzpUP2fi5g7YgS/lt+wHV
r8vOTTkxoWRirgPpvpUe8OoLCT91SqecVajH1tBvP6y99kCtMCLIoBlUnyFA
/iv+Nx+foqiVHzbI3p+NKCxGkX2YpIJrF7E96oVh3W1VWwH+wHIdCv6lu6rP
BEkEN9GyaL4OPUvxqLXFzxgtvq8Qt4RqRhpeTliMaYUnB5eLtuefbtLK3tAB
YcKC3BwAzQoBpcSRsxdEvWsD3EVwRaPle2KDJu/owxrNmesbDeSAfYiq4bjm
ekq8b8HIEeqyBX84GQaUNkoVIQQoXGweNUsBmEweYDRcoZ3jx4f/fY8/OEJI
IOEarEVTUJ4YZ1NVHN9SWbGOU7Jh04wLJuX0Sh7n/16crGGxE6DC+LskgEs0
+jeACgm6qi+nTBJKWAM84J4lMO/ruXrYYXlvFR0kWVtv9FDmKjoJQ/usfpvF
KRRjZCSzqum3WoceU+2TPPlOZB9ZVbM2R0FkW/PEGd3zIVYEHhhCOJPOu7Md
F6VhwCgbZNDg6elZx4aAmFSNpg6VSQ9SZheONJjHFbvKlpN3UB0kLrLorqFU
Vrx9Z47yhr9uv9UwOT8QhaBzNsXaMpe47Z/xPYoN7G4FIt6PRIreO7l2D8S0
txpC2Nv3KW3A493uId38t6NYA6gymqj1mASY+J6KlHs3SMmP2kYC5oYzkiyT
37c+UJXnyKE+wWJhbkKkqe+QgWWNVDq6QgRHZk2l/7nlOFoWU/9bdZ858E4Y
vFTkmbYAXcGlh+t4v8HaQPvD6Hx3DqjC/FGz0TkwcpJW75pP2CFhP7rLdZYH
IiTcPoNkjnSIIj388ngwejoIdTDOM5NWzpxB6V+vl4ichdHvdjpqvS4T+Pbf
dqoh1StCQmal0rtWmZFQBt719DHYXNboxFF2mp3DQyhW5WjMINawCV48nuoq
+UfBYpACRQC5qlgzF97oavvNpxm16Fc20RXQGmosUlUVrBhguLrkkXgO9Rjz
lv/ToWlidSXcJm0fIsZEX0idMIX5LeWkY/qkdWcufMA7INrCEzGvI1xGGcs6
So0cMqpVwRlA1XQxIj08dA9EZSt3z8C4DwtT2WE6jtOMclAqbvUGHzGAM6uw
8B4ZzDAOxe7g2qhxJhEJNlznayO2rw40VbB4rP7eXlGTwidGniAwkq+awTGg
4IzNrK7Ns/oGSDUAdLAh5l4e0LJvJSHcwQR3By+Xmji9ijRS0tiGAUfPWw/6
4p61zT6psu/Ro1DuoaInrmSP8IBabhyErks/AibjlecidlNkIUaOWV+3LGyr
PZBAwQpHEuDXhIqb8uVtR7+sNGVOfPPUsRpWFnK4eZOIFzZ43v7BaZIedQ2b
eeGRKzqy5d538AYtthnB72Vcrf6HhUArdSaA4HcLCvJS/ikB8MWGvUO6+PUA
vMSnNK8ncVVM1o4dIbWofHmRcNsqMPMcjnYtTRlyDbJ+EAWGVxDCVjxh7cod
u8/aBD7my6M69acsRFZp5TY75X/A96Ck6qL/znB4E+8LPur0NvfNfwuHXqrv
lqdyKqYba/lvTDzP6x/QBE2byjbG+8aAErJhXkw1xx9YYDk6mmFsWS6WPOeO
rP9JBQrXHrPYhl0g280VEgcXhRsr8yMlgFOMZJZiU2qS9ixRvpbKOqJQCndR
QDpCZZjmSzN6laSu0xtECJy7ejIZxjBxZle949tgb+zJfXlle2l8HM4e86KY
Aw6DCe3oys9dCEp5UAR5L577toUltOiljgpB7wPcdQ/l1dPx8kjCy5fOBYHK
R7EEYd0eeIXTrPN3UkZC5tYAe2I0hdrSyobya3czm6L405IQH3HB2/v5Qhne
+4zesOqVQPFWepLiuKd02voe1xWfMS4FEd0I7YxK1Vgg1jDNOlbmoebs8FaS
WAVpJiu8t3Sy/M01Uey11hLZF1/ODA0/rK4kiRZEKhwHEBqmSM6kTomTwdqC
LglhRi/PDZc4Nnp8o7yQE6l0yfQTYMrDpP3tiWQ1Zm2Bj7q+NfFhtvAGfUYK
CnQ0FDziWClUhMn7/ffMFzwVzF5Vl20WUJSsYWukdwSaUYleShQ+eXFB/LkQ
t8Y55PYoi04kgS0LO0y5ND81SQnwvXAavDfd/1Ti+z8Uk4AQyod1NzC+kldM
vKeVNKH09PM/wJLf+3IFBnlCu7T1SEpfSDvEBIQOJP4X8cbiKYT5pnDT5MPV
Ta3VjTncq6IX2HCbc9N/H+IUREERkKrB53HHWcW2mhgKs92l/uOMww+4Wvqo
ObWGkdfkOQ/YX/ZavdRTAL1PXHowgTbmJhac1+dDHY2r6kD6XrVoIGfhyvl9
ClIQAiEu2/HuheniRZ3yly993VL+2NT8sbBHoFw9d0no6Ap19Tdq3DSNvRiX
pbpn+gvuyxz+1v6WSzG8sgI7GXcYm66wfS3vzrfQI638gbjHSQxwUbZs4Izv
CcWQGLxttOpRfISxARApQapvwl209+K77r4etcb2YD8qCTXG4Ip8rMzGRb3O
aXKF4lL8Yrx4j8vwInV9lieeYvHEf3zFUuFtwuQQT4/Ts+zibY8s1Vpb5YOO
JitahqXbIzcwXF8DBF1+YQqlHsZOEBn2/NTwtxkTsGehksa+WfkjjZAQg02O
p3xYQ6j+JhvNv6HQIRhlSw3adly5J1keoyBXqWOPHK+DJwZC3Iq1jXKe4fbx
VpVPIEK4d/XNNaZZpLsSSQrpCePChl7IAD3rGowhfLoz8c1dSEGBH147o93P
dljedoAX6Txs7/CinapB1TY0KCxinBhDj8BFb9ozmMYv7PQ7B66c2YLTg+L+
q9HrcKM9tNpAAstF0VH0vLJdbwNgzJw+E3AJ1Ej6IlqyW3dfIU+GVzv6PWwG
hGseoNbIxQe9D4waTHO20p/jUThp0Avhr3UNytRquZbE7tBipDsrMSKkakVk
iPKyiflekzSztdd5bjGjkJkfzJnWeZNhdy2iurTf6h0w1PoCSweHe0tQVJLp
oQDw+7SHRxnk7hhBWHXvR7LZRy+6TplGe7l7GB138QzlGUWBM59zS69INQyq
7E1+px0C09KcvMPYYCl7d/jDRCrgspfq2EpGYCba8JGz48Q8cXsLTCDN5g5T
z2cfK+Ci7R6WjBwF9z2g45NZr6C5iGLREnCGslxv/YxS3cXzthH1ly4CLZs8
t1OD99Yodqig4zPJkpVYDcgchh2VUzOlb/uA8ybAk9N0IiiwO9iH0vtJsEUu
5WV8sLKfVKnNJwCJgbrSQWTT8NdvUxhHXYcH+4OpGp+0klu3GUynDHYrvbki
AVI/E+NcoQeCfmdyGAatoaG4I5Ky5uT/UYoN5PaaxFaFz+ZkvbsVFdKzpc4q
bnhyIlJcbQWiMJU3S/bzGD8n1uSwhWXM5ogv0d3MY86HW8qEg5z+1SuO4kLl
sCGr1fx0vbSXu8zGc0Z5loxLANSJiIya57tmOa94s6GS7CYMEhtCBXyCOSce
t8eoccU2C1E2/aNjKBsdANY364zCBwfzRF6QNky/rh/wWBDwcBIW5t8J7zfZ
XzKEciR7b6Pw2e1LLYDAdu8duc2fu6k+E9DuIxcUbaZaifCY7Ixs2Gi8zjIP
cgCTnos+9Em81C6tOEvU2eh+40Bpf4l1ZDb4dwwRGyhfbR9J3nlHaC9vlGtF
debRW+OdXVq6OzwmWvUm7l1ZSG5DSVJWUo72fJP03Ffqydm+8cyfhrqrBSXr
LQjrOfojemIevD6v2JK7NFUjFpKX8qxTIilSo9Iz0DdtGd/BjlT+DgVdtbMG
gqpAo4l6qK9QyRVLQ2nC/hjASUDWLncSUMnegz/Na86aHrBZRWMvT6STsDyC
Y9QlspSrPwWITqNliJ1eT6RQU2oYB6jF88nPqUgM9Co8P5Gq7tR0UUkGaGk6
wmuUMIEFwkyigS4Xo6JNE8RHlPeOu5rbgK5sm9tAG7BHLBwCE0YDYIgLwBPg
qmdhUDyKimFKEPcQJMqg/HioeHMGoFuEwWxttzj4JWCkadABEAoS33YfhzG4
7heR0cemsjBGaC1o7wboTpQ8nOVgzj4bCQ7V4ARW9KHujggVq+zSJ/QONHYY
bNJ+TUTPjcC0Asdyol0zy/XyreDzl/9gJfIpk1rVrhbpfdnDAkOWg2aGHNDx
T5aBmoWEZCZsdgJdisTJbv+sge+T5tmgSgiehMkaGOEa5ph6zOtXMc5aO3Vu
OmaTyhwikVYOeQkzQAJnXZzls/3SIT1Ux3VI+Olsfs9+hXvlFq8l3ECSIX2B
URlEcflbZSaHxvMZVGxRbevOpuYDxTzeViIEbOrzVcIF5pUdlRavrgOwS0x9
pna0xQ/3Jije8hHZ1jrtNhS9z4hV/eR3q3dVUxMFVtWcUr7ZU4GvFhbe5Fm7
AnDAY1TcaPOQY8KXRAmTUFiLdn/IIKg4bCtKK7/dqwCqoxP1voUvHFmfOYZu
RnAKUKStmut+YI0khnSYcyMFSc5vvCiWR+frsTS9DOU6gFpvMl1jSALgqn9C
sVQLOmY+w8c0KFQp62RXvO0ZHt6ykG28It98HnINjPMQYCzthNUcF/RDO0YG
Ka1mW5KY43JP1iLZVfvJ++Pgh8XD1JELVo/b1Z+f257c5Ckb8RVZXkD3KzUb
m/kJ9Mz2VCmt6ncAiYm6JnSQZrUec15hsWvIXAtlCpUHrzYSvQYyp3WOGS6t
uHfajCYuDvfTz44aulmQvQKDp738JazoZOy0qsdf2s+Dq+tb61Kw9RNWW0uh
2BPA1CApdEI6Bqokc7mTWq6qiXorJ/CMHR55WN7zhcYLvwvGwv8RUDKKcqFt
UQBBSitcCnC9rK5TS8ls6YrTOtkXprCNVC7jshVljaJwrJ4Nsn5RyWeFajCK
qgSVqoGPXPNMSaRk6Wm765S7V63bGskCgZL2TPIb31oOw47DiFpaDtSH53bA
EHX4NaABBIhIh8k/OunMZUROFtRrxuxyxlq8Z120D+1ZDZC725bWwIKryOzZ
BK1ObbdMbJ5014LpAOtN/33RnExhWkGEktZd57hG1gLCVoUs0GB+2worGGFf
dr9ejCgGoUGZbH9a+VmxTlglx+Q7IrAlLVxeFNDnVcsYbxgQFE/M6aht2bOD
uIBqyo63cqD7q5WQlkzn8OwtLR2+xfapDKqUFVao32F/Ww+p0nKEJtlnBt5r
/TQ277ECuj8WZovOdvzOCrEHE2Faqa714KxaBna6XIv7U01EJ4P0ImHaKLEK
G22cxHDvW3+/LRZXjkQEKeXeTUF8PGQkbLic+whxiBCSXGd4lMmeX1RIxbnj
V/vYvY7p0liRZ/Vb8a1W9Pzig/aDYvx9FL4EipIvYR4y599T2dW7R8bFhAEy
m+2TSFoDIDPB8cNvbMV/n4Oe4ulhGVq1swCtDplVr50ayGSaXYW44W4OBMoF
BYNlsP0463N7Buy7xhiDg8YBuDgCdP4f/6wWGnqKWMUOGiXP6weQiLBo0Dv7
JfLGfRH0ramIGhr2/T455eH7rN0Qv514dwLFG6rX6Q6utcsFzRWri48vxw+/
TNbM2JE/Tko8lcbArosk9QtEd6N7BsQEVqrN8oF5bu8tRfG5M3U83In91nxx
0+OE3xQ4AR6ObiACR41l9KAy3avnuppLNqUZDHI144K1RHtVA4siSjKqotZZ
W7l6Efv+FkIcJFRppaQx8MnysndKHbXtioGP3KbZBfB0MXEWJPR60JA5eCDo
sawUC6KlS9QNhhkVeW7kvNFmI8sTaZbOHZ7gclcAgQfH0fvFVThAaManmVY5
SLQuhL0zGACcYmU92cF6A5ngtB+cBYUiceyL+y1iZqPPjcIyZlZKR0K3cgbm
KfTf1B5dED3U83OwlfT750Kxb4Tz+fMenFwfY6TplNnLZAtpSaY5bhawtDYG
8zvommTCbhmhyrXHteFf/t+rpZVnhUPCk9ceh/9UdfSZmQrZvJDLV7PAv2nD
Ny/0eGjLySkmY3SO/tQ9fbNuYPDXru23KXAN5H3DFlG3Vf0hKq3qWjFFsYnh
68oEP9W/Qi109AbpyfTqHEf1uBYhVw2uyMtdc74v3oEyOXZZiS7OpeeyqR11
jVerLOwgRXgp/b1rhBU1nZCwWzI0icMWeqLUhNQMaRmg75Ku2bvwGub/L1p2
8lTo8us6WluHe0S+mh3nG4MJ9TnRehSmmlvhZLAnZbrzxOo1vUif7mC7B7FB
Xu6iZfm+2i5O8PSzQek7M0cshYUthUEtihHUKnx0S8VZ8f4W5ZmjSWDc5eV0
549x8Hw6B8/zzzv8UOOvdOeMaI5MAWBrE6A83sgM61CUif14+gza31+TH5Sj
N+jghyOkPdXF9NVKpK93wmSqE312okC6NGEm67xwevxmDhjep28XQtog+h91
rUvspyXW+ToCwP3KZsON/rR8EF4IkokrRxf1RmK4X06NtIU8D03jcqmJJNAr
eoNfG9Iqc982C/TaIAAXpqxK1IATTkTO+LBxJ6VL4HQQYF0l0bQZn9SA8U4K
ktexNI/pG2aaxcViWeRzw87vpCtE11xgDJqy3Ejr+J7tMpE8ZZtYiQVn6zt4
XAxK/qDfSkS0r0J9vcJZRamE/bUQ6Cdme8sWRvPPf7Thk9Drd9fVhmASd4iJ
y4ipovn2EgEkw+rJCEJeglqJioNGsDizCh/WZ6TLYafDdxyCfvk8Yy+sm6DS
ewJXJ+H9LSu93WEEX/VLwLak8PCc71s1C/LSMR5dVyTxHmsc5s7FkZUw5mGm
0iL06buAbm/ImPk6tgO3uEmmmBg6fqb8US2+qxpMTv1fr26NGYZxkeEGfjfT
RMyNaRvpqZz9s8o2pDrHhP8TqkiRKHjc5+lAiIL+Bn9OWGATQs0FSANcr/4v
nCxzlY+IgQupynKYfexZLSW3a9X98kpTBArdhbMEff6JS5HbO2ufMtknyKUw
okWlmXMA5KvVrsYeXQ7//zXHMhzHLM+PF7Aa7GZN/8ZNuFrPxCSKua39EKjZ
Xm3+qYv83PqclBvR+dt47U42K+Eq2ESMvp8s3p3KSedk8DkJO5ln0LtkF8BQ
xRLLXh0sHEmbrdCelG5061ctrwXDnoX8otq/6iNpMmX1xrVkwIsbIIa87QoW
Us2c21Pmo54Psvv7o7tfFe5hYWZUe59dwG+c/drQn/Zz+bwyix56CnumaFuC
vOySuZs1Lw4e2PyD64OuvtOB5e/2WWJ4P5k5n9pgF4UXHmT22XXnFxr+9xem
uy7QwmJzln2bPH1rBP/4yizTElaEG1bP1p1kD0Ianh4QYUsdLPs9Waz6ksi3
UT+i3dkfGDyEtG7axICMp/mASgePUzke5Kzwt0N6MipxKiZfHU0UQWCUA+od
T3XJiYl9tPaU3z/88t3HvCfwbfYmx1L+6S2zLdciwOKToqu6Q+wCfG37nIQG
nY2oDqpaW6VstKwLi0UpbklHN7yEGgdLbW3LDUD21in48NNBZWh1AhzxDVPi
3ER0/fgJHr4jDzwKZCjcTiB0dqGUU9mt7ZxOV9SprftYfAoItg5iGW5z4445
4psGbOlzZGxK2yMRrv4zKCKwUZHUCbb+jlPCzkluMwhd1ZnSbenFu86HEjo6
I0xQFv5F23sdpWL1TM5xnUXZBN3vHv+5n1jhwQIVJohIYLFkT8ovY3IHh25F
NzHp7zv/3BR7aJ1HM3TKDglgwOTZw1fdV7FTD1VXfY9m6lpO+EZRr/hiLEsF
H3IsQm5QiA+sKZtfnNZb78VoakzG13Vspf1KkSCkHZvjM7l/MR7tppKa0oqx
/TU9kVZ1Xd+u7Gtf0U/Pz5W7IIyO82z38i9KW8/9NqsWOpnyLHljGk6UX3ZU
bHeKwpU5fhQkGKzHnfkxkEZe++Y27e3DqwkD+MOWF6JWYy/Uv15uZ96k2lO+
AwjnMD6Yq3+HDoJtw4LmE4XRzoSnInuO8mGpmEYuraS1WnKhQqbOEhYPV9c3
ldZ3oaynblbigBI2h/dzIksMRsUvgVGDqBN3seTzhhO+nUlhvbkybCX04At8
/uAXOF8WgX18WK4HWswA2vQ0/dpWG5UQltecM1bd2Mu3OV4mF7H0blytBU5S
dlLzocJWwO3uT9Pl1OiE8GSIyCsA/pV24ZQpbg+DRt5a690P4AlbZQlIv0IM
gNZo4Elibr5df31dLXbLxvIGNUwjGxhuB0q0BnIGTAyURCd0YTvVFzMlRJal
XZ9JtFwoWVKiI2IOKDQtGXFGDFCDZNW/o80cbA4THusgf5E4ArSaobRJHThA
N02td/UJ6GUSCyWqQ6hrbLi2moJySD6TKoG56IeUc4JupEW2rdrH3Qa5PMTW
GK36BOGm+GTUbkE2wpr9GBpEzwK831MHVqTMXPPbGBpyeWkeQKSkekSnqzug
SrrNEkAvFzhZ6txgil1XPdE4GxpllTt+PFeHanTi9pfEG4vBrTOm9ubFWWOP
XdqITjgvqFEOaztFiGvjhYmcQ/p391HVL+EdrDaAo52x+CPIeVj1JvBb8NuO
o2nF/cZdqoV177w/mV5V/m7em5EULYifs2jRHSC6eQF/ICaqPxSOo3W9vLAF
oYavK2veNWtQk+am6mIEkYI/KzRqlbjRV4eRiH+45memTgDSHtrZ8UDIQSXQ
wuWeFIVOf7GlnhEhLDmguaOztIkVWJn321kvrbjiHHNHrMuLxuHgAJzncDLa
paHWRusDzXRsNFjrjTyR97Dm2yyy6EplFo5z8JT94A3Hu65bd4e8CYCqujed
liB18x5aDBAPoalodyVUmAM6IOltDORqjqcy2e+adadAkrAL1s04we99Uh7s
EoCXaRNqnAlc1J2n0OL3sz4RvIFjoKPVdKMTX3oaSVyv+p1GjT9GJHmLyORA
RRj1mLclWQWTn/wJ2djxnr08X+crI7tQm1ArpBCCfp48jHIZ4rzq7ZgyNgZ/
I0lURiE2W/PoDYBB168gX3XsLsFTkXFRQZp6QfEW5yEGFgn8/OBfJy0Myhik
Dc3GKCbf0kRnU6iRKDQRVQ4F0crTwFa40kYHImycpq0Gb9kcR5UKS3k9rCVG
nfVI6YYRr1xirJ/XB/I/z03ATagFJfph75CG77JTE1tAlgAQu6vP1XsBred7
Kjhyq3U+nSYF12UjrzkW+zKC5S+lXF7UMmqQnbgleVTeEQI2kBqBtrMovHWh
aZ3u+Di55lYE0mRS+hMXwUzYUzOeaVtvhjq8db62aaaopt2nSPFKFxgTmc0S
J/hRI3Ud4yKhiZy/uv5XyDx8sSXzKGPFenNw1B17Bl0bQaKobuCRaviE+gfk
/X8L5QYZtcqSXQ9zXQRMUpQGWA6kDjsZ9hP85Yx/B4mGtE3jj02lZHWvPOMo
bbkUdAy2/roJoZzG2YdcdiJ9I1xwJoSmChzmQFQNCzftKFbna6KWGF+Uw1rC
qgfgiAjYHbmydxkJzxmjiPXEgiwEBx6BIpliGj/9Q5E8h4Y3NsqiJheQgO0E
qwZTwghhcwSDqGjVPUq087wnxl9BvbMCiRwzrIET8H71+bcGQUkf1owHBGn0
xZTAADNsU/0r9cz182pjujLemPZ4Lz/etqeXtHmO/W+3T3/ln3KCrN+B4GZE
DeZdfWZZrlsPAMXs4byE/BFsySuZjzYCfImkrzXC6U74fomiWL+pFnoHu1nO
wxLGqFJgzBhbcL82VaSrJqS0MyQNQPgrrIkuPvrUk9AwVjTpAA6PQ3i729RL
OSJpxFETMEBn44L5bala/sqcbeRBoBEZvzra3NUCIf0imC+PPH7ounvSWrIk
q1ewfPBd4Q87eNIzQqLu+AsHN0lMuNOZwXhe2chLMvRonrnVd9n4OUAbw2zP
YoIzhn8UyFNZcHS6mXmuNe/GFiRUyYxoPuwS+roeR7/tZhfg7Z/S4oJXUteu
ELaPcl4L32ia7OTkBqgYWmfn+RHRB1ZPO5PsHWTv7nJqczT3unJqqvO7BIjU
K2sGPRx/V8FyVWffi/WKtUWNqsZeHulVG9T7tvm11Q1Gkar7lsZBxng3DbA1
38SW+IyGg7wQwu7bixoLqla86TQq1zAVGRlj/JAi3lUTJB5jN7yP8UxdwrYk
uc+Yhce3ELwPaOcjkUuQ+S652PPSpxoHqi0ETz14fQH2Ct1Ke6a7a3lLhOq4
0pv2sT0ML+q6xg+30SILTBf25tMYXPBzRitTWk5rMVb+/zSuEQvosXKk6P3g
ua3Z6lwlAogjsOMogl/FI6rA+D+CRGOs5/jv7+ILO4BwGMijj1dWace7nn33
X/U3m0SEXIDMUejpQ/MMC6Tj57AXpCgZqpQ2+XmE84ekC4u1iBNP3ZU7iBWz
kKRrJHroTpodw3L4NQwvf+uoe+htm23pnyxRGKZcpMlW60xxE1Xqp6PXjoc/
VHUmp0KaHjAbns8YtRDDns31fBoleK0ik0NDCs2s+vOof7Gre09uZG5B9fkQ
YUTL5DHqxMITLUXLDF1WT4PC53OvIT3tAkXeZqr/CliZDjEekEC+XmDtxgTU
InfoBsxAt+YUGmLUnLdDgR2w6y4/U6PIRuOoJ6FC3tdNUxSbHnGgsJ/TVJQp
xocRzSIW56FPZA+As302DocnaQA9OPXwgeOk7MknT6Z8zNYN9KxG2II94Szq
1sLJe1JhYR8fb3phQ/M+Tt6M5MMP55zHhe5FAFdqYjQ+qYWi1E/to0KgcFG7
wxvmRyGYa9Ih1eLEapvh5ZlK5mypcAh6vb+j+Ao1ntMux1UFQK6jSaG+WYFF
WhEDyf62SxiUIXNJBrQRQGphj9H8PN/WQLf3uVsWNqoogAjt7n+LXdaualDU
F3/ZL8qV24/oFSCjbBDxv6bJY+UFObgMCcSyb+OveVsa5s9GLL81B9ip0UpO
YWfLfR9XS0UOVDotSXnMMmy/fQ33ED8NO4p9nf1fL1OxrMSOxgnM1qv/ClDw
flR34WLZNc49nUuEbh0ON8o40VrucZRI+mP2gwWk8oEWFtQGJUC1tGbusRlc
dO8QR4ngeiymtbvVNTYg675A/cEvm+bqztjzJS5t273bDpiESC49Nvuzs++n
M6H9vsp5AW0naFuc3g/TQ60C/RKyHvFKkneyaFkSYk1OOeVJw8Wo2b7bfDka
QDcygAvl29JE7QDhsRAoJcKx1vJ/I8DdgPaGscClQL/qX6HsPhxyiIIDdhNS
08Dn2+si3JGlg2P0wIs2veVTx3mIuguuOypmH+9ExPXcTKtse/Y3srWekY+O
l92BcbTOKOnv6n9S7pdj0LAUqjy7z8gmLSwZT4v9Z72yoYRG3AE6So1vzCOX
T9Ty5rsBUKjS5tZeUQ+zUzDXTQT2PEmXrALbpR1chWFLGSqpoyhPUe63GXDy
x1TgStSaYyfevYxVRNcOtOGPuEAQHs6UXl5lBt0H+znR/EsOgy9zjHqApJlO
5zoAqR6kvqTzk6ikA+FVsn/8NpuMUeEQpyyd0jHILcHh6z6u6V6bXNpvqKJ8
L3veVJLSJ9OWKktVHWmjq5bTkKRDWC8HSy+jEpbR2oHj/0GosduyBQjKO01a
H/XyfQpYJgTLPU4gnRqzax0u9Vx1gWCOZpwXNBjxsTW8TZyAM95rJZQL+3DJ
GCWTg0OBn2+M6fh867VjcL7hVneTxdXjxA+73lgMI1jhmXvPKUGWmde9qdqm
cA2VL1dxK47lqujmAfx6eOQY3Jfxj9ql2LXe1vFGEMIFGWgNqCBXKBhXI+2G
JjmcmZX3yUGru1DP227sl5mOcCCOG9IVU2wvO7hIbFJou6AWWmPR28BNWIG5
31BieFZPyZTlFUSSnUdiLpb7svPDIjZJk4B8AOVN+uuoGzKWXDBEOPtogkxA
kMerCwhG4NKcZlRA0unoYDcLV234ZW8r9aoWXv5FKT7zI3zqmVsSEYeW+8GX
nvvzrxW2UwyrGDqhJOopJd3io2x3he3bBNtC3UTtJr+byqekej4B/amNFAU9
tpKYvstkrOOWu8lthql5+4iUpBDJMDlJV7S+N/z93TGNo3JxK2OvrA2u+w6B
l7Y+DO6V4IqXdNPweHuHnO9opDi72yVj8FFaGXUkgcdu637GFupNTyzS8gb6
53ZxrIgndafuin0Mm48nk/7fW27983QZVXOIZBk6VFsjYEpy/PJTvGFHOhh2
sPzqg6jagPZixCjREcaMd0lZNVeNqVcc21ahs1ZRyA4p/pPBRMS85uBcXVsm
IvhT9jDjS2MDXsr8GqmfA01uOhfLvXtsSlBB7gbKhR5jnhIZuWT1QDm9VTLs
wcXiyzcR84CjleflCPJr+4BEpXK9VD/TEZENkiaZH0zH49WAFTMz4rAVf2ql
xGK1dpECboPml8n+xyWjrCD6cNownSCTO8Wn2EOE8QYr83z5KXNHSccxW489
omWrCnWszP/0mqP9bT9Z4iSA9nHe5ffCjTn06FUJQtyrB/UpISPLFwcNxB5M
9AmNYtqnsVoZo+bDa/O7QhlrCypDbQ76TDuqKGxFgFXqe1DIpaU2KKxrJ0mI
fMozn81/Z4nFyusN3DA5JkZ/ei+fb5hxDtJ7RbxC253BULZVduzgbYbzo63e
fUGJKC32bJIh7RkvjlsaqFWTGOdlZaaVz97ooX+j7/qOkE/PeYG4r0UOdI4K
sfbEbbMqnj7sXt8rYi8nyqiMhjsVtqNlUduvIyJGc5ekmdBbglxxd6IvnRS1
TFqV+s98sFJuEG8QbxxnajGQasNZqdg1p+1rRftNHv3SA1mCns8vxv4U2IfN
Ly5xCiTfL2QgpRYzgU0ol7JnNr/zLh1BUh+pV8V0hzXKHUqsEPTqFvFRmrGO
O8wSApEmKsspF63Xa6enFGN7jssdqOrdBouU+35O6CPXzTLrCQgLaZE1SIR2
7TnzHJkRgD8Ikb3iiOLGxWA91Da2aknlgIOKZ7ePsbIhb1RfhIO0jwdGebn3
nSPk/MlhfJCeJkVbEoBGcz0vL326/f3Jps5ayo+WSTfr7NdRxkX8nmH8QCS8
d7MahiVxTQtua6nIrJCrRyiKW2rfEYcEdJMB43nxM6itOyqftK86kH/wO0o8
JR6q167W6YT+/eKNFZe84k2RpN7IWkH08TBmppTOV2+RBhAFDz8/bFbpQCwK
/SG1VUoXTreJrlD14C24QTn/oi+BXB9I7i4z7w6NkjtMT3ggSV/6PtBW8qZp
aZkoGDzxkXjgLKsZ0CvWbT2ooTcC2UbBInkyT0IXE5V+8K68iwqBnVuXnRoP
u6uqnIcwkdZHPkHQtCfXHu5ATDAfC+3awRBcopCIE4MSTOfdfOovwBWLhA0z
21VPPJrf9msosf1haoC4gatUNkhe5AoMOQ/0vTS8/oNsXKg7UZwTVgDGTlQm
Hb4BNhkYIB6D5WXCy+i9bs/UXbUI+VtE/yDkNy80skNfxnHn2+Yd7ZRIu4PS
bdv0ued+EldkOx0sO7kzmnHpyj3nb3uFGNzx4x9rIgwMmO9qy2f2XUU4ULnY
RQRha3VVXmVYausGWthPnCaDeIPzwU/GLod60qev5+J512lzqBZ65WL4ekeG
CQjSMhXBubPyH1O6U+eAQBg4gKRpEfDYybWoe/bCAMVD5tsRXgSMiTO82e5b
UvXiaF1Pv3JmhFHaycQTdpoTC3toBO0CjPr3e1bcZD9hTjn5EZrUavU7PqkS
JM+tKoG/bF2jcdcuhVzmwXCTGkAHdIrtFwj7+R4nsg7yckiOJwW9a0JG4HRW
djcPcMCDRq79gaJUNX+LbyQud1Xcqx+SUoXnLCkZAY+sKskV8Xt98grA6mtI
1AuO61Q6G79afvBzM0JLXu9fn4lmHtSlrGZqlHm78BtZtN+8tqHbu7C/kKs3
DWWsyzFR+mNnbKPlvoK5FFVeRxny6YXR2gR6FJkyjVwtO17ARYff0bFDrv75
+m25QCkLuEuMMQDgGgBCHuVbGL6a7zIPv4x/3b1tW68vik0UFvQJB/ZqcKfD
8y6h5KKLJNBHvtU4ZhGt3mpjgYKnC0oqRm96Hi6QVGPpss5H0PQ7rUvBfBhN
lNXjYywN40bd1krFkPY/VPu3LVmM8wx72Ahs5WRRxYJyCbv7k/thPimTGL/P
YlKribdbUbF5rUYvmrc2GGOwbQN0ObJ/7cfUOpdmxDnAv1fP+2T2y2G/DieD
HW7VLJxikFQCxz7dK1HJ+HotYNOiLy0kz+dL6ISZUcnflbElSoMJD92sQG4r
IQE9bcSb00uyt8HczKGyFJ4UjEXaNvmyLAoBg4wejzqJLRvVBVUySiOmzsEK
NQpe1ZJuaDDWOpF5xMnWwQhiL5Daq8qjhrFi3SRvg/apBOsixLAuVg/laejJ
9TVp4K9ag6uVa7fhVXUn8ha8QRc38KLPyDzqcQbJ3bBho8LRjm6xMXdH2oSM
hI8YFT8i98dx8vlbLmJcA4PRF2nF2Qi/niod35szikWEPk6BIM2EORgOu05I
NJaViHsjWXKqE/JLmMJXdt3WDpb4o5qF0yNCYp7E7xNWe0MCc5ct5Xs9ziyR
/Ocv8umpkFhkR22sCUevecI1MY6o2L78a2c+TrJqPlsDVWS3uc0U01DMxS4w
PP8x03SjiNcSvYKkZkDEOYdX2IQiaCmmireE05UyqiBde3x+EZOqt3u6eJxO
dA9pesjwySJDtFVf6R9UTQXpBomy47rVIx+P81QWBzIsGuMXoyx82hUwXbFI
5oJf1vp7k+zbQ471tKHzMIKG/E473GPBLs9gq2gTGCmNHWvisn+1IGpmAbqL
cso1zotKgqNeVfYbJq1WssIsYSWyQeIvafeXjJ+mkc1f7z9rqx1usq4NdUd6
51dJKo1LKtl5kgvBOJn0/eP8L9zaqKRDHeCXF6b5i2dD1LKdKgxOjWY5dRte
Mq82MpRxALAzOBpc5vrbqQpEb+OqfB8Ovtkg1GR37d5BZXOMbEaXch4UyAUV
fuZmtaDuuRo1L3T5sYzIIqjoQ5TfWhL+dEJor1wH70d13bf71jxhDXjkLEVy
f6eKd12zo/gjXHkl91vql0qmbLHDJRtzYgzayeB7CgnqosTsOhlkjyWFFXFf
DBDtqZpKujnspZEd+44FJNR99fxI9XGFJZhZ4e9giwSo2Vgqc0yv4s+o6Hcu
FE/+Yi8cpVLlDpZZ1p43SN5fXPaVNoL3KqVvmg/q8hC2s58DndND/Mwo3Pua
/Pd7wL++o/Glwl3HtLhjLtUnBT5CcUuDusV+NjPumZTQL7b6avyIKx7rfBjK
iag7CbKeE6c5wh4VQ5DzsmEWaNUhM5ct4KxIyVbyn5P94uUbWURdJKPFQaWq
s7ibECLYeKqk7+mGlqEjSDqEHQaDCgjErhnojtyCkjNPHnSL5wjAKF+T6wnb
PSFH4bYvtuuO8cbMmYXE6+8oW1rRxPry3nVt2ZxNXiHs20k15jG5d0EpzWMt
UkCX8nqQrZeyPz5HHn2RPIfoFsvtR+3yrCzThoJ/Zg4R+G16dJde3Zq/QxPV
NYFfJ3wj0RCO4VqCAv1tfg41TrpzCtIY6CRIlOaNNukRh9/O2E5DqbwHsDti
Afw3JtPeHDHmAfz2farsmkBg0K1uu8uwzEV/EjEYbPkuZjLJ/P/knXAirrIn
VAXV3cXv7BtF45eTWUMzZ84xDBsQ7dyUVMWZhodgoJZ/mSQKcXtvsBtZmIBf
+mmeCSlPqkz4ZZ7IqCvdcCourLZOmqQz0J4OXgfy+M9bze0CEgPnKTY0T/3s
EdvZ1zjzUfmYaRyh8sbYYDGYG3g2CaP2/9848mrNd7ZUpezosZMpZWvcfovM
eMxsNPamX45bouwRUTEK5QGb4Q++Urc7KIG9l19QcS7sj8aNY3d5nbLH407X
xA6pyg25Qdf/qw5qHAr9n12f6usB3o9RPORfSA4E0M/v/t/c8o09hVMoulPm
IADF5v0ww2Rb/a/eh1CbTHVJeQhmEduPq3mcxNNpcSqC2tGpqBsgLDRpP0f1
PKANKeNmq5ryRDEHdvSKXszX3oJV71qoGeXbWMkhZfZj+EWvz5qFDKADgwP8
OjYE4FT8Vl/v3sA9DeYbWKrTXkgy5CwQ12gpowXTbOZBETnuqRhCQ+uayQVQ
ghuAYXUp2ZDHHZRoBfumDLGvGR6KC4632ASEi2p2xxTViWlMgfgBVGnWFyIM
K5QYvEB3T3JDpsI6hjCakOh8ItnVIPjkOB6MX9iwOybvBEkV7kJYgyQVO2Ds
s7bbgOove3/9MGwbKYSyEg6M/QEnoRxoo4JC6B0BJEesOB5YK4YSNEb2SiK6
CG8+CefzuRF6HFN/aqf9tlQnZd1MxN09d7/dYqCjsQPMG07j7a7A3yIuFW24
51zO9Q6GOdNtQFPpmuG0xHr5dN8Lk9HIARRsCdRHfGfMneE85uMatpmGXqyM
4VVGyZV5wfa9xM67exXSuUt2jCC89AIhAs2vFEztlvlLeF3JNWlLLIebcxnB
bRjxPWy81onZ66p3je4YkL0FMS2BberVnvpMdRidR1UURsNYmX6ouio/rXRB
Fe2bYS9NenR/S3UCemBt5gsPDnQ7mDP11TSPFc+Hufmjw+IpjUo/5bVryXRE
X8A+lkfRvGi+JNnGELmJBO6V2+Oc2Xwdu7W4d9Zqr3ITEgmN2ArZl+e927dp
AftMVVQlQx5YRjSJhQ+tzNK/dJeZDwokflB12Bo63KSTY/GJWyDlU7MhrqYE
3ghVvmKZMlHnAbDVv+jrSu97LbtFJgBydjghDLeZ+U0BOT9PEfK3jtM13oyL
HNz6VFLRH1vBeHG0QFabuYcRbmMoO4J2pRrYCbw50etFoKUQ107wKQBLWl1r
lJFy+BVUbTujTVu6g/EkpEZo67BDoNKNGikAXKLLCC1sb7eDySfiHRP9ggPy
qMRFu7p8bJXePxr/38lYfPgqNIqXTlMH9UnEy55QrBe+oCu9ilK/fVWSR9G+
sBXH/MQM2qnbk0KDF7ZeyggGS1xSQ2gh4pglagZEvPY1qLnoREBqWwwy5UCm
rtqNFfhfM+Jg3gI6qv+XBPE0OD+MNZO3tiexAA1Dm8mNbqpU+xN7/XTt9P2G
r7tK56CJN0VPWAR+fF9sI3FTUUI3sLxnxTSLOsrJf3Ru0+XxuVv8N6c3xFG2
w5HyFIBtXb2J3kcWB+JC6I9N4ztE1gZLne7M6cNK/wNKp6Y4mXKdlWp1mp+M
KFhd1Yw9kUKTMdwaYPX96Jzcy0KPPB/T0pqjcK0mp1hfPZCisB93uvF1adw/
dmkOnD0H30l3szelOKyKYXS0WIn/XQHhIjNIMJvY6XBXF/MDaDwxqMEiygW+
/EOwtfiMdzidTz6MfJTD2UKDJZwO9BGY6ftXb/TbeA7auv2jaYzASCe3a8Fz
SVL8fpR0Utlj1DaanN0ON/805WyB/CJxHbykAaSNv8wfhAiT3IvROc/bl7w5
nrrzPkoJ4Xsy8TsVALcN+AkjPB1OPKsrd+SaDwgSn/BMBA/mLau1eVVBWdbZ
gz1oJOiFNs+esql1P8KOETQwvfWRUCFrk+e3KFGaGsQPoUUNnOwNqLql7ftJ
NDpaTkOBNpXTowZg08iodmpxYboSXIE0X8b4lcIhyELEqER4sE0Zdo0NgTx/
OXI3Vqgp6tpczh/NlDfQQJ0LsW69eoYCfzOGbxLVGglnvOeozSxP+QumFZ8H
flBJ1UXMAkcjrW78ZEFtWeq2gKiW92ih4TcG9sDXX5hTHrSe6No8OMQ/GhAq
rswxe0aBZOFgeVbuxW+gGhVbiTNJeiClNuTxi0nwXUCx66iBpepTzRnEtsQo
MhQ/ZBBGHAQBgSz0HY1JDgGrDu4ICkq40vschwsaFA3ner/mUlHHhxBIVefI
PHbccChLlbJlOnfuQrtDcrwr7Tt8yKP2oWgeAwaHpsufK7xpgqgtE9GmSEbZ
ZiARz8/pqJUQwk8pqZrrxALcFYKpPyVBrlsBv4G3VAgjwGD19A9frooHGslG
S9el4n57tqeyJ3T4kjxCJqF0M3eMIJ3ksBPN10wENptIcmAKUkJNTo1X8htk
fJycBo4vHY8rQuEXM2X9515L8a4N9A63aX5QirPCFmYP8fyPoE1puJ8IoWFc
FAb5LoB743ym9WD8PwrGMtJw23naH/2TE/tRYUVMF4q8/0Dh0zhxLiZb8P8E
611AqEWTdRIxM4cI8zXEAROOHSjMNBmKAaxL5p5cooFTgZiDsEBtjmipZ5ae
V8jLdl3Bu8SiNuTZYEGhrNU/3gYVttfMPwCU/f3TGlMKMMkHHbpVTgKF4dj0
PNwYjXS8Emh5QRq2xrgYL5fVu3CrCsNxrcLAYcUVJ5y5N4Kc3oheq58ZYtfU
W4W+oCjr8We3aJ+Y0J3ngqNpSMExiq87p5pRlC0LWTOl3bEd4lo1iFL9RVrU
o0yn1rDX1Ue9zeH100SnY8EnU1sAVH+tM0btObNy0J4RyMGRuVtcUvPVQJHc
wjeWCvHZaloTHeukx2MmKd+8qCZCg+npK8kHIrtvSikjWlHfZIZRZAlLbj5V
cgg77WDHV5RMd0ofUCzQwBQBs8FtnTa90s3QcstyfxjEQ5thWyEM4DkuDKn6
9X65uMkMSH5CNm708Wijk/cHwv6PRp9HQFt3aZbNnhgzsuJHaE+W1vwSkvHx
O/CaNvJwYKqpL0kcx6fZXfAcOMoph5jLXrIpaIxIXxn8s7wfYTT/hZgMzblL
f19LHMwPD9MU6vlom2Fi3D+DkdIWoQe2BH0rinKg1s7vdn1/F40O0N/UTQHM
/cTBYCJ6tehqXgOTypjlOv81YArD9PjehevKHXGtLvvzEfYf16vw5bjht1jO
8rxSI/etYY3ysNnuF0zSfX7BX3o/f0RJXtnRBhFUAflfRoNcImhRSdW2fTXB
bJhPl9viMETJ9TmM3Qg9AoOQKtvZH1lxELm2FcwFSO5ab6lm5YmWQyWoDE8k
vpH+B+q3xHL9Ra4s65oLnIFUYYzJmKPXaOVOhu20eIPcrs75CSvlwGAYNsih
iCnMoJ8UXS4tWQic/IERpzHgRMBR61GGbnNAaskI6Otd9jIdjmDvtCFY5Qrb
BqYZbiWUt5N3EEikSd9Meop7doiH6X2/kTSOk9LddbEtbtxQPf/OYckA3zx+
ahN7YHk97SqlMPS9GEEiE1vPVPwgzHMIKxCzuB2F17ovz8Spv7W2y7SjuIsf
+/7f0i2IjHtr4zp+iSx27KQgy5WTD0eO8iF+VrCAWxpiAL86q9DQPP/ceTMx
nXgtZxQJy1HQdKr8SkwkaYWZGDi2txT+DC/0xNFxl19oF2J5lD3dXxDEmB5e
ngbpoq7ZeJJ6TjoJZnteOBE3eEqrqqYnN++rpe4cvhU/EkisqTyVscVu1Upl
nGN3O9/PfDi5JTG2CXuJ7UnU863Cb85gIqWNT2i+InO6RGU15IydF6y8+GK+
TiJePVNClTnq7mF2t1TlFMgCtE/PTq+LRhktvuBvphJwpbX3HrutuEf0r56x
e14tvNdOK91eoxdBqkp838GKXoPB5kLdwyqUTrVDoJk00a3H0b4sWJuw4UVr
2/nMBdmLuHis1PPWTkjXb3OlPcEIUeLrgNIDGnkdwa3yjp2ez1hqxrt8xHwi
awnvmdsmT/Ey70fjvHPAaXd1I94WxEsQ4fKLhXd3wh0rfliXmdZivp65ekX3
dhdoFftoKuiUmT2rfaf8EzwrUlprOqVmuYoD/twVnSLE5EV0fgZ2Hvbpy7j4
l2/htSiumjjrTqMK5TYN6KPYSXVHiYNFSWZlvlVmDPoO5hTZT5nzd/K58B2e
8tdw3Pkcc+5n0+my7a3ECLXQCfH49CvJXGAyBHChcib3XokAHSf6zdobEcWH
e5kWTmALyhfP4/nn6RM6KJTKsxQ3K8bYLrIIiY15pfSa1zThB8oSzsE7gxAd
Kx95140EyUg5oeNV9rUe9fB2VyzLeZhRHj22UqcIX3Kz2DYBVLYxkONwOppR
SyyL/nK1NxbGDxZKxBvXRm59sCoNPSW8pcQeCllKuThXhAARP9BsqDZCkAFq
ieLSf862mXjklDdE/zy1wrLFt4NY5JtOcEEAWtNe8ojq1mlIuo/VqOJyimmW
lAptD3wKZv4J6lmPQrXuw+OTudQIFIUVak5y4cG/dAEg3RVH5vEyJeEC847n
qMcfNg7QRRBWTS+8WPk5AxSMrGoloxwcninMSu2KKjFoOs3/quNckHA+jng/
yt4fsv58116FV5PIMI7+UyGY4tITwzMPpYKEuHbdkn9C+NXuTLNxlLkUItRz
4Hx8BWyEMREzQJzqE6mBMcHfLY1it3nXGK0KBWN8vj4H9sdv2rtADnpRjB8G
epHz/hlSOj+iOLUhtxaAgw6Q95Z6PMbz9JmfwxXLGOw8ju28PXZKGKCIvIKb
ONANKZwgnuwpdsT6NYbOXFeDdZVQJuxMBQBaYgkyHZwK3vt9MiTmxoiT2k6R
JK3+CeeufMvtBxfpfmA8zP+4/C354ZSATEL+BiOFGnlWhE9xn4srMYagIZT9
ftWizNBbYE3A5DlUUe8Uu8J+Z2uj2N3bg/4taFKXtumiU+oVUAbOKxd/gk79
51cbeIYbYldEkPuupSRDym+q/PQejQ0JpQZ40gw6PNN9EtzmwmTB7yLAu6EW
10sXMZc3sQV5og69FSEHo+qO1qG2ww0eRvj13ocCHuOJ3DTcxLceIyVveqt2
4ZjS+QM8C3m+cO7rt0MimZhyFd3GJV+FiM9DqK57rJ3EweJlt3Ez5aDjUnig
utRRE1ysPEQlKTp9uqwTable2iwSzuwYE7SFhjdmGfxcMOxXQyO5ciEClsqY
EyL/PRb0v+UmpHkD4B7Lg74l/mvMaC0HFuvS4TEisIIaVvE3j8ZEyUwa7gj1
lu2I/Mn//yap1Md+h+AmaEkN6OgYGcXrFTzecPSvMsrhllNjaRdycZiQuAIL
3Dc/iwzbyHeQXymKcPB9UV5wiyCezjKNhFpIB0j6Z5ZbN0LEtgfAyHnSLjdP
hRb59B0LGjN3Jujx9G99U20Qs/oYPLGNv89irK/89JC49lq+4Y650LLwPeq9
QW9Qz8WIAoMkDJuHj3fRBezIt1Tdx0yoXE/Kr/M1OtxohzxgFS59jsltUvU5
HEwtRDWdQWcgGboXWmxjjw5KD2X0klGEwGQXwd8J+auyMtcTsUhn87KHzTYF
fUImVcGYd1VM7wuRaY0KZDvSZj6Nh7KfdZq4s08ZMsYMOVqmPpRGAj5lA6ZT
AEBtBPofjts38NONvc36rM5rm6MQ0x5PM0f+nWqtFaSc9KbYPmkhUH5412N6
DhJ6fDd05pW5JsvPTHCvxOjn3uFFUuTGVzqQ489sT8JpUzVbov7HML4TK8l6
uhqNMFoL6M0OWOeplZoQX16C+UYaSBz6/2yxt8L0KueqZ1nvi6/rJnJz+Jf0
lwFo79PVDKhH/pnsOD16ru3PDVoCJamK4RsqCCu0ZLjonBqyvvFHGNwipb8D
VJwunXECOvmLVI2Pg06KryziRjXfXsmWd9IRlElXQmUbS9+j/1Ud0JiKyZ65
XZVYTxnEGy/MO4/R+ddvI0DQ8IwqkHNhxf0eoMf71TJRflWkfZtetnTe1eW8
n+QKr5BhxIN4bCADkhqmVzctiSfeDqpjEAj8rdZ/RqIfXyBniCPn937t7tf3
YRGia9nuNpGvjk7Ucvv9MUYsVTwYpzEuqsTLl0yHTzLZbo4mgmxQus4Ft9/0
+DvD3/NlbD6BqLgg3ZFEB2xOeQ4a4DCtsV8Ac3eI/1Ha8lqC4nyk/OsyXrNn
wGYyDMiWiV7/L1hhmxSYm2B5QB2KAFiLp0LUVZA/DGeN6yw4HSil3+p1FAxT
9zmkjOKiSNeOh8srOEHxHqSjd5evqH9QN2JBs+PPIcSUVVYrPSx7b6XIgM9C
BsLLqqDKzQ2mWS1JvDaHzre0hc8EuCMY2bblGiqgsix0IcJrTNLbp2I4um/2
+e0iNXOycdFfdgHetTnCDYJBDbSNl49Hwj0csaDqkQ5zaXyRtVz/RLMqxV4W
yvHcsUdCv19mpF+R8nSeqnAqGx6O1D2f+QCRlA8ihy/6wsoP6qepyBnzuBUl
p5+pFpL29+RiCaFUDr8bJWLdNaGy8kFw2JgrwDJx1tSkHHm3BJTM/JZJA9l4
ldyeZ+1BdmWmWpPvtrViVT4t+RiDX659JHuFNMJB60Kk+3Y/d9Cxf6BCcD06
c5/U5krSpg6LItq++5g4a6x3nbhkLS0qtjf4B50+1QGgdTR2D+Q9MiDThE5f
S1hzizIcAFEaQXX0XsCf3eqCKoOae+kNZFVnyMB2VyLe1jwevUJ9GzlrTp3N
l75OBFvykhvGRQe83NfQOISwx+JLqFYn68EsylHXSKi+11auqWPEUvGIe8sW
2N1kt8tLSj9C8OeQx2Dy4id6ShUHHuWKsnpQE5ifUid300roQXtSOXieoL4F
ihB+VFa8StPTMbxbgtF7hYQreDCxLS6f68mne0UnYn+Tdd/h3k9hhMCtSCZd
IiaDt1Q4njNGJ6GPB7lkzX3FOVt2tPGnnz1RST/Jblia3OZ/FCJfyov0+7Z6
ncZKUnjkrcu0wNm81eX32uFTT3ZYygta76GjoyXpuVJjQQAl8q44iDEwGkEF
e5oFubf59sBPpKWiXwuvC4+Z1EfVX8ySkIMKTiK6JP+pa8hASJQ5yrHggu4k
PhrWyDBzZkmrVreuhl/iX8fVdNgGjmIVM/PX97GMD18oM4DGhNMCYuNdiZLx
rplTo8pzQJMxBOqLzJ8IEj5RHej7LTcA2pBwUkGBqb3J/+wumXSE6HLU2ZlP
Ua+XUb1Q6nMnqJJ+ynErosn5+S3CqAAqZqn9o+BCu3mxnSIUoLeca5z0ObX+
ibFLd6S00Foczn7BY9mHcEXdA7s5IocSaijE9eiIomkQoilW/Ak/hbKOr7i7
KFd9XgJhv2FQKU0gWnV47BXlvjloI/3ceXNLV4fz3yRDXEjWuNloFnABStk4
emIWLEawb8+vp9j6rhBFUU8mYCOcNpFR9GLeXqDYBoaJicAn9It48hb97MeJ
QtZQ4yxmpverLtKPYOi3VgCXhqcxpQZlV+AvMPFs4SEPIyRs4+lQ4UOvzbqt
PUbtepwmV1zNlmmfEjj9yQsRlkuDhJY1Z9NBlzATGcqIrzXLOVZeZA+qo3Jn
g7r9M6oAoDNU0CGWh6LDalL05REPnkm7QRKvzt5stPKD/IrWErwOVO+0ujI1
+QuwA+y8xoqIsp5sMd0YZrcsCJmsVQ/fXBYAmmDeHI7tjebzcUzFF4C4TJQB
y6fJC3ErD7m2fYrG4MWb9wEgii4EyWNyfgzUsx4KxgGWQpZFxodoq+dr58GX
lt9cG8yb2WDJiKBu0L+xirLlRdi/9RIT3NBAY1SjRYSOAPuxpxGpDPWJD4ro
avncxGW9CraTnFubfyhmzgSPJliF9vQpTLlPBahwKL+GjaQfXqtyKjJDZfAR
oBhQZJAlmuAICdrSYjveOxUBp43LFNLpZ9t5Kh5fGyQhowJmbEzC40XkXuJC
bHnw0Qc6oxCDrAALmYV1s/Q03drd4zVlMeQvJGscJVN+d+ajuLSWqVBOXYO5
2ss/ZkhNj1rwWjsMK5Aoj93sVhOWUsEu0OljajMnKXUUQTU289sn0RjOA78v
S0VotFbOkyhd9r62HbFuKroH8c8eQ2y9dxgl+1yqZzJmDR6RvShCxs+vQ11R
K2g9fAYUi6dc3PvXC867GS51YIEDPM6AELanNyj3hyVuG9Ns2Y3vCO0fe7wr
6LvBEXZU0LZsQyAJFSem97qT+nKb4lu5yvfBenBKxXERUzNgEIePBDXb8BEd
p5Gz5xks2pXc3ILxscaKBIKKXawC4tc/8+NLiEDEhMqtIBOdJzTh5icPkniy
yhsEdsOfMxbVs3VIrM8eUJ3d4LdtO53tnaGRMCQKLMnO71i8kJgvkihOFn1b
Avfvp44Rnnm+qKm3lOZDYwTN3ix6ad24Ah2nfsDfgtjRzECYUblDYVo4rWF/
wAEKM0QbJXixIhFOYTi6CG9ZjYEUA8F0437Zc41bBjO7ekYA4ZkmB/Odes90
if59dIuDg5lApznc+jxHwb2z4hvXBrXaodN7uwPwxmBvkPapFg7sv2qL6SLl
oN4gmvQ8vjXRgcGekHCuHXco8RqJPsw+8e7oOzw1eHDEndsxSJLgLq3/0cUd
TvyK+Vxx1RmrDrPvbvBAf8KyYtNZHzUXn9Jzd4CHdARVTytoaytbb30z5ih1
40mX4kpaG0sYnzLrVOlpUZi2M46VGoiKybGpOxPxiT1vIdUafyOC6A4Wwna0
KtxU2pNpfZV1zUv2fe/c3n8X/DS9CwYHXTdf/7bJfN52oTK7X3SVjF9Xv/ZK
qLRD6aS1mdqEGKs0m/Uff/llfy7Ca3ou5MQGYLUfet7Yi2LOW5yjOaXLsHbW
9YoT09MX6j33fb6F0AZyftWth99Vw07mD1IrCImDpgQL1uIpp9XsH3dTix94
u/b19xasGThVQi7MOcZgBX0csGV0d1HnQfJndwGY5B/CwWJI0J+Gre6Bnf/7
T8FI5PQYTYDTJlMz4ZNJ2ICIMZG1aaTxoAvrGiD5VAcaq+do3bV70hY16IC8
kZ9IADWWLx/qEOEAa4C6Ve+B96jkntCL5yD3+8idMpRPRsTv+gn5Rc3vz7yM
XmcwUXWaop8+6huEE25Zd+DJmlQHjmm85aEKnrhvKBPEADowl+SlGf9kLfmK
9CXjzdKlMzkKA2ZHTUk7kpCuLL/ybywLjga/J0Dts1DSmrL0zwCM8j+2U/9T
Puyb6PAoDH81iFDCPElwhM/4Eh4zzqToByfF5la9BuTePDQrchLuCKTHWApd
B7qqZK79tv6EC1FBDxusUIWv2zOXbsNXKzArV7dKA11OZae2EaxudUQ802MD
zis1g+LZEF9wIl0yEhd0E72PAevY5mHwV7CAoziGsuAENMk4RjTBdE+CC7lT
BCY0H7vSH1FfisomYtKP+RdFhdFcapvkjLsckrQrM9XCsq/ftN5DmgCuRPzI
RDsV19so+RLaXAWTOJ1+b5hVihTomDJiida1iuwZn8ILco2O5p2zlWydQB98
8SsBiKtjIpBAcYAf9kF+aPqmrjCmc70alocg7BVX7/Do6gC8f0gyOSim9DuX
LC0e1U8z9RPbyPMSDI96fxGI7c+pb5Pqiq3/d4cG7GAyTythOlBtI8o+gllB
7ZWs1Mujg/8RQW4LpiWmKQaidE/ikIxS/T8G5wzafjerfZRUPoDPT9XyvL4/
qSGzXoYIHmeSfA9tSp0Tvhl/ltLel8iI6VGRXCOvk5R/5mLUePuTjk02ntdC
twmKs1qwyll7SAHs1pNtQu4+TR+Nx9nJOwYcapCw8ABsEqHSfAUlVic13f1j
4b+DKcGwrYtxqbOw2fb0RfY5Q7Le2U1gelU1XxMAoKX0AylDo4F+kzXbf1kQ
OWBuiOQ5djhYRnptvD1bHUZs6WZPZo1MnzhSk1BBgnxJuSumkfWfytfupx6L
/MSh2I0/EoS1I48tkFwQzy20LuT/jbLkcHTGSb8ZW5roq/+/lIAGFckFB0zI
0NcDEbSmpEtqbwYOFrmkG554nQBQC2ge1b1EI7gwMdzIsuZixhs1rAnOcKTP
RKe9rSXqpe4cPUUQytoNfV8xlzRDVc3xWQbn6KlS+4DNOPv80Rzn1zuxIZXu
ZzirR2xfJsDksCPtNHmWDOJLJsC9h8DwiZz+cU57Bj+pnMQTtWehBKvY84KS
zb27dfe4RUoc3bZ4KPkYuNbb20SwGMLzYFenagwW51D8b+qaROHq8DTmZV/q
3PvrmZOHkcM1QPq7jVeYWtqJBJZ0ARqAkFk9djQLYxXh8x08GsXQQFYWjhk2
8F9igi89zJpatIQQdyqsMiTI/uRqqr+RQPx4zDDPbh7Hlo0jzRwpdf7zrn1/
IxfBoHwOuHRsIRWutNpGtfLqiYaWd98GbK0oAIxS3jZWv58pMV73kXcXm5UW
5ZzQ4PwbkqRrjn6ILTLoyP7cSv1lSsvqxBEhyQElK/mQnx/7KIP/+au6MIgO
Yi5lbLH2fI7nkBiAVzsg+wmBPzChgj9RvxO78byaUhx3FjoiEVtrLNZQLDdP
zL1mxgm+4oEEk2mit1cNsIxgSTQyLECN1HeD0CITI7M5+FC/OOWpk9PIKQgh
kyrVYE74vJAaI9cGlxaH9XsK0MjmlHZ/jZ9bjk7P34xvxT75ebVf2+2ET3/3
LWy/1/MKP7MgryBZtdmspxmw9AHTt+ifFuDPXvVF228OS6+cWJpKIV+5JReq
1vsWbGOMSu90YnLp3yOBiC8DJupfOHzOlIJhwfYdFUO+XpbpHAU9GC1RGDKx
UUZx8BrlMvFHg+c4+s90d9urXINlsiye9Ak0qNEIb9nXxrPl584xii/or5mo
36ifXzg2FUUclJhfbaGYv61DV1XGfIeSCtm1BfEp15VJvVnc10JvTNGqcENu
Q7Q+7+sH2UZgo1CkMgakgFeVShEig72We+yoF6C83TXNGAlDYXpggzPFRMZO
1DRBT9qTrI2WpQygtOhH7rpTLLxdKLwG7FtnMw8w7lxiTJ9sV8trad3wjMMO
U4Sl1hSKqfuOFd1KRiv7gmCITcm1CMXSvlbL7sQQWzltHGsx3vxgl9BfA14/
K26LKVKxSdvTrePTF8cGfOtsEGEmxQegT8ZaiNnUb5tlNpVOYU1Nn9Aop0Qd
cnFVUDPodBvEHZ9FHGFOb60mGas2qcSnyesylF1JAyTBHuaQ9WNqJn9XBmHZ
yj8qB+eoC8328FHvvkApNNL81jxfHltDM3kBvVzDOBCg7S9hl3cCa/tDXSnm
vsRn34ssa53WcjUGVNF0Uk5Q73Ovrp0Y47ouK/ItdQv8sF5+GXnHBpKhlxjI
h07E8TBROQUscxifSlZeXuVLWe8EiPXuAnzal+lwnu2Qn5sVIcjJ2C0aGpCD
eLz/34iaiODuWIw5R5IVrDtPO2J0zNXwrIuEX+Y+kz3dPRxgbu3GB+LMOQsE
QlzP91JspMArJzhbPGbMJ+B6UfyaAih2I26aMoPpricwo3exXGLfkLZJLcA9
NjWs3Vqs8lqc4oq2JGuODfAjSE7a08kMzuXrqjMuztLWJsRyw5fBXiYalz+P
qnPi4eg2ULEeebhYXen/elh9kF4qWBBx/vQKKtSTPObrkiJ/SAVW3uPeVSd1
oZqmtOb7PXKHuIHq256W4AVr74tt3P/utzCXQWyWS3g7DwNrQnwTrS3qoBrm
E+2wQjEm+UzucE+a+mPinhshrQFq7s6+4zsxKSFtt+cnrntp/EGy6/M/2hiY
PeNhPhZuFmTaIT0yim+UWDtHk3+n4vEunvwOtS/PicUs8A+zgxKD4fA37BBY
KwD7Tz1Wr8cy0TsTcrCXD2WQ9DquPI5LGQ8UUVVyzR0/mt5ca7T8tVdKDs9o
MSfKtKYQXpsbFEuxercStAA01ZfQ6kDF9pSGlu/JwdS8N/DGkcI35t/jqYMy
dEfMMIka2t8JIvDercFUn2f7iFBwIgNODvfKmyFUz0KS+L7EsZ4wT+fzVNp0
au00JIr/MBfgk20FoNt5COWqw8RbKYas+KwpizGANe+OsmuGR1xXs4N3/4Nn
GfSYITOQDR57XqGcPKLs3WTv5bSvAAYAUkhcP8auEWJ/jhokou6ofB2G+X8y
ZJSnumXHOjiYdjPaudw/Gqej9Xq7L82GfLgB2pdeyvPGvOV4t+i28pqtf9Df
vEFtwVOyvVe3QA65n0Z/oZqqQz5CsOy83LDd1Drx0/qrHawERg+SInWPc93k
YU2eNmYxekjfasQoCWeV0xyfMXL2gdNIc91ZO3N58SA9ssdKBqXe661wIDtO
5ZzAU+3MAsm0Od0r61NEiGNCUcWJm/r67V+g/JFtA4+nvlOhpfEmuDAhpZWb
tezTA0pcJCKcBHhKa7MrdN+pDeMFARfXR6WDn45YghNddq4zRt9ZgqTi73dV
qYX18+IoCiRe6jk24P5p5y1mgyFuR6VkOCDm92nnjc5iT+3611zVHQQZpRGN
KJ9t7MsytL4Qz/1d1tknjgLzF6DcvKG1jCggU5MXSOCTzes6eF8zA2GctLgd
47fXFqxjL89YYj5psngL+fW201dVGcNrCuChPcn7kba/9bq+vgRVfJLiXWfS
iSQQe1m0DuFuQN4Qc1jB33RZFJPEUP62XLl2D/vQjlQ5/VYqlLdEHOChb/oK
76QQO8xIbKLqtJKKPfed1fTPPwPoju5Po4cwoASQFmETLoLMtOfBIHpX2qAq
J+qJcn51m3GV1PDVZ0RGlx2iroLzqfkncMHniuokrcIwXxDVwJ0qAXzaXpJa
odS4FKFIeG/4OallT9RrWi8f6zUdXeMKHMZzHeiyP0MQbiehBYvHRPXKVqne
gOV+2aDBXQZ2BNCnJpMfpA9d9QMETMXdlrQv6l92MnwuTNZ1Q/ppb9OjYXat
Vdn6FGVNs91Ex8i+6Dkf5brlHQTxOkjUX+ntmCD7f95dxCJBadoId2yxoJbr
Xe9UidG0lrJDuANJO/2w/5rhc4lM3wZsQfTB54wysDLCW3FgHTZeaMez6p9k
pCkBqNTCa04ybVOOOM4GqlDQreB6+pKaEYheOVp4mT6a8MK2LlL/Af8TpH0j
ts4KJWTy3+1yvbavuGR//SWzUj9wI79cnzit+aQbsU3ndwIWYGkusG3Rx8ZU
f3MGYgY2WwWLR9pdwHx1ov8JAoHrZVD+HbPUoeoEpqoYG0iryUSC+MCi6+xv
+wFP1PVNwzvO3Xh2YTeFfqsbdUX0ATs6q/8/63IC641dCmI2GAuCLIfXSWKk
RJxXWLVoDS8VLMbebu4qHxfmoLrpsSt2emvp3lv+/XFywHE9F3GRQ0sRj6dc
wfGefcvxk8aygFxvhgoKEykT33LGIcJayLzjaAGs6tP9+/aSGfa4+XPq1aTJ
zmipxFkT/jBplF+v5zekFM9kg6oi/rXzzlqUI0Wvprn6ELWMweTkTF3+SCLe
Y3Z5SlyZUngqmaxOwf7zzGkrfFNzBHNPcDTDfNo97u0iEJsSiJZ1SKlizHTq
otwF20zVml75GFkiMaJt2EjsdeTGYMeDHjRy4ZtOBKsn7h8MPVp3+OHTgbQI
TtdR80bS8SerZQQnndPed6DlROgHIeSyrrWfmmhmzibWLWrjRMd2jmtEnL+x
oD3DAkfD+LH3AkRtC1x6O4lzSglvFW8MLuaQcf6Zbw+J6KDJcR/Jau+WzR95
rpP97NXeIviXFxx6/im4IKZt3Old9gBAdJSyDUfHbYJShlibOFouP6P6DQpx
Q89YFVwFQPzT1mq+gwCW4rx3DNZPiqgqoQEUBmX1wtdC9vWG4COS3Ctqk5nL
FvcNKlEz9FSaNMRni/eYQMK95CA5nZJE1ZgWaMUre3/LxK4Oo2cCp/cWorFX
jajktkZHpNTR3HDlYvEg5cX9k7pCel1PeC2fzvdBxw6QaDqnYMo4cXZ52FDk
rO3iqeSs0RlyGXavLkrxNunYGVkS1eBOQ/HvPp9v6MAn57m9nRLpHHRhoOwO
Kymf7Jtu9Qkg62qBWLnPw0igY5e5nzoAahOE9dB30rFtkoKXL7e6Fyq7FDlq
RGYsP/DLx16TTPyydWJwnEoQMLAoLvP++EhUizBCHYHXs50uxETGCOZbZX4w
yDIa4TeZ7Cfl+U2Htz7tZstkg787wyyaAc66KQAa15C/1gaDUetts6kGoPI6
Dl3OrDTwFlyfOywinUeZswVMBNX43KzNwQV+pmATcrP/QcHVhHHs5H5lQRxO
MnIqKbnzjOh5nuVFxT6uZPokTx5TykPSrHHKAOjf9FADJeQPIfUshdZ6geon
y1enCqD4lSGfCqNphCjHtHjKaNV1dr1Ap1NPLuBh/CiGGCM8YNZl0bYDNkw7
k608aHIgw6+ouQxEdkdOMGQXEYCjmse2QrkGz2PQPPDLkXLuE8LLXhsan/2l
u35LYw9T3AVHORfXBUelzYxws+pqx8DYRuqK3wv7hyvx1MS4/h1UFXsgcLTa
HCAxjgul0pmD9jwwtHy3X5lZnk8NT+pfH+pMVSurF0vq44TudPlbAPdjPD9p
F2QuQes6B38D8J1Dxk7CgrQFYhRVEDHt1kGqFYlGDkqI6ykjBw3TZOSbwo6p
RHevE0Hymo0QJjLzgIltQf0Cqe3ebjcJ4M6mRJ9pgJ2r6wSiSJI60JDx+/e9
mT8o/PQIhBWcQJ/ZZfGuaJD7GA/4+isLFvl40o3s5SH4kIH60UfxfOdP+lmM
yMYLT3IxQR1Jdfc+Hal19M+dGpzLx5GQMTplDFb4AGwTUyTIO45cwSnPw17F
lydmPQ/kwywlLOB/GbKH8aA0MXG78RbcOjGKeoBjFw5mmKphTGF90/JdON6j
qRgU8LvLkvjs2XXXzwW/SoFPxoEE2JROcLifmfXnqhm+u14VJi1cvpfoIS4x
9knPD0aPrwg61gLgb4GjgYLTgRNSbN9LxcXETEJUu5n5UGakHkJnMHR983av
/h/H97Wvl0HLXEKUZB5h+9kntOeV+D6WvH4tkyD3CtKXlWjf/p4XxvjwtjFD
HPXmHkdyIzGRPh4pmwgqGpnIlUiIiLunaSBnQtnoYBNk+3YSkmlGf6LEbHik
+jllY+YrEgEhyE4DM1jlqwKhNjaQyQihOm376XlgMUB2TIiwb96hjItebov6
4BDTJP3B3FkBeh6Q6VSQIMdFdx4xvouCo5+peqdzLch4mgUFGnbfe9CU3fMh
yh2OOLS0/HMXkfeYN3MYrpJT+WJYlD/ZWi+0pCCK8tEW12YWyXgLQJZQKXyd
uoC1+rVZg8WHBO54daKrhZWtceM9SDqp6p7QBqz2Ip8wfwyIHwMOatCkjNrn
iVpSCD7kBiouZcd07wsu6c094ili4GthipCoEBdntLOPMDxfVDCLj1jc5NB7
1kuCY53JG/+gohERDopCa++xz0bR61xTz8jkac0kTFHb18X3FInICovARc/v
qBaXtzecLrf5t6YflTbJVknsKvj5cNFRzmS1UR43WwE5Eo6CgYWqcmiLp/RE
Y5nS9rvXqbs2YjvwjYq0fVNpkJ+zcWduE/U50W3UzFZu5UiaWXT9yj+DvtYT
CCNlyFCnH2aGakhswDrUDOb3UXN1DGKFui31/RpRKwHMnRg4mtn8vgGFFg9g
09hTeyu7zmTiVfAewbuNxydE/FItdyaGxXVxJodAYZ2+8XajgpIVCDAuENl8
M3AGa0ut9k+VVtuJH2fHRqQhXN5PP/Q7MstEqXUYUJIWcF/Zzrv4ZcOGX6C5
IGZBAilPXpYh2SD906gOh0vJGgf6hFKfz3gyC+5lWzqZMcpNjd+mML2RfkEk
S1KH+BqmjoF8isNlKMAmc5JZr3idMxpj8Ttlr658De5jYWwJcOEmBHsABIMi
IcG3PGeAFw0Ps2D0jOu5a3Xe6NJrFwh105cnZQu08evIAZ1MFaOS7AOiyLxB
gaZwRHSs/mtApmtYM5NzdWxZWxcYTsuukt0vCxbKdAg2qhGGU/VqNbSKmwW9
Ouqx/BJ9Kr+82wypJgLqHtQ572WVwsN3d6Ex49VRE/aiFkojSChzhG7Q02F1
yLQEOLshQDCeYTN9T58EOrxrlrFKZYpoCybAdgMG5XJzKUVo25EI0gOgHOJ6
Y07iUF2cyJyrtmpmTvt47ClkfER8e5u4kEcp05YlaUrlw4D1tBA50SZp2QOR
tlCSJ5QLR/7giVebFIG47XLOMUYIvgYGjN9eSTuKuPqGmKsXd7ClBE/tnvRx
6G/mdgdQ0liU4xwsOLpqFvuyh0NEIvx1/I5ZwdSMrc49lPBy6pF1xozAAEfY
qn4bcWl7F059POuIQuhb+9im6+YEiO4OrPj6O800X/qLIk0URsSgYTlF+uXH
wdBMZOTO5YWE08v4f84i4XCPYOun7o7Guaw3/WByyKgPMdL6qCaQcF0hiNnG
bbX5Z/DniDvC7JDkeUH7NDVu7z5HRtDJL1kcJ4xl4u4MYXXPa/bTBSDdTA4b
nHHdvnbDrnNTjUYlK3DWQ81Td92OXt9KVJfgKlHB9IUpQi99N7+FM+6+j2sG
Iud02EK5UjwtEzcarpF9nxHkPGGz8Yxz4ctRea3BExCE8X/dI3ZILXaNz7q9
lNypnt9u8imVbfN6loLc6SqiFodF14+L3H/dvPU3NDKlBbICLA77XGt7DMcm
9z3XJw/Q2v0E34YPLH2qHm6U6hIVlkc2uR8UGQGgukhqJX5ugRY3d7QWSru8
XKRbgobHNTQ72WPbFL56UTPdyN+BUx2dSUYFXTvfolLsmcU9zmm9tgX2gQnc
jbMazzM+moLiTUFnZs2Ui94j27PhXIFksAPpgoHstcuhFaaVvLCwmNdchDtr
rlmd6bd6Or2AOle/5RVgOOAMEmJ4zT6736XBsqQAxT4EUUlYw9CcMXhogZ2P
BOh2kl+kOnH3FfJDFTwX9zKtxqIWy4YHvFvgx2QRntC/NHoC14NCr9mdFbzC
RSafioa4YcURGSudK8MLKewr0LfcnE3jJHoSNVzdimT490cEZWQxNnuExMZm
eAaBiMCNazHMAkdewQN78ttdv6dIQd7zf645SbI9Uz0TfVDQaxhaMY/SG+fn
R0jEiB/CyqT+ynht613jQq8VizVezd3t9mSYHl3hu9pCq0Vw0KaG6sy25z/p
f6PZD6qJwfNrrMkoiYsFdaeMU7QeqkpOSUna0AvjjzI7PNTPwaSNAnsf+jTv
1L5xfRhLP04ZY3rAK4FgoCKr5kc3AfsHd8FWbO6y3a0bmHE+6fmec4Y13Dxe
Nfv1S2V1hVYVn5zjX/8W0okpL9TCsxjT5YmtxUfycEUTZXEw9gP2IgbugXcH
n82CXYWoCNzxJNdx00COnaiE7QE08v1Ldh/09+thafGMxfmoVgIatS23wOCj
swJq3DiJJCmT22Ki/TEYk8DkpTkwylJ7Vcnd4dxCL5i9ilPlxlFcUMj6k3FI
IgNtFa2bGfR/bXFGSv02KSBQuPswyKO+7r3+HAyZgTbb+zGNZ6tevsximiZZ
1CGsIg4RM3LITacauThtK48OSWwuOgW6jadSQR7H7jeozbTtIphTd9PwZjWk
ffXJATzvtF/l4ocT+L7b6MaHWKBA4FarlLbzQnHM8FuUXcVXHPQnAyE8bMTI
8iRPqyl8DPXF9MXKpLczMyMKG2Qi0Vqn2DbdQEdJQw5orghrKj+0H/Ld5ssx
XZ9pVuVbM2hR58/F97k8Krh5mEGNSvaL/5FrN9jq3JbrtUiBfnwiOqEfdSYG
cViBjYMbp4G0O6bnXpkJuk3dYnOv8mUx82jhrwA2/n1K9fZRot7S2XBkMoBg
xSbFDb6q7hiPaLfIto1/TJmgSf1SEaKMeE9jvfUlxdA9eddP2ToQbKNU0dBv
CYFHoMf9oQ9DLCEJj4wxEwiYIgMdpBCJAsFGMc88R/1VWg6Ol09u4d4BVH46
2NTF1fieiHIzeUftwRh/V+7eVOrnFaRR79ZG+8DTbMUF+Vg/oXLMQYBmTYkv
Gm99noO5ZgIAx0jZDDT4eOHMDM6OZ/Ra811++EzrhvHL7e9LI21NjRjkLfH9
XAj8KIhFHW7hOr8zXNRVp3po7h/xpqb/+oTBSnE7YqCRQ6NGA6HcvK/6wNut
AfZcU0r6AvelEb6JobI4NYDGQZNR28lgg773FyPU8pW9G6MQU1v/bLxPBD56
cgBtbuIxYY1mAbtJu3t9GXM+MLk4BT+0csqyCEhNlXB4v8N0PJu+5nVmUJaX
hB6K+bHMDMK4JfXDkLgZnppHL+EQVEaJSCQ0f7s8lVAkKrD7IztWCDBjDB1q
1x8R3uA+9FWCvriEtv9TXf/IiTzl20s+onwVK2wCTN2SCbzBQDUIAMnYfAWE
yC/khCN6foqjP/cOQ0LPPJKvSngmWWthKRKkoK9c3YXO3oXT+nTD5BP5cRMX
8To4Yosz9svdsIulAiLemismO0Kxch6bx6k2HMfdS31wot+uL32Ag0XCbJ3d
plLveEu4stxOoG4rbDGF3NnS9gx0EjhkW6U1GeVjSdE63Nf/QZeUqaDVFr+G
epLLWfd+xzTDtmdShuPH/Bn7wG0y3DIYUy7oVbg4RTnLqkURq3cyVn1zxt8f
w8FFfNcVbXLHdrm+CNi+eJWR9YQRo3i99YKczngRQLFbQv3Stl3iV4oBKgpf
Q9LvO6WdiHEOmZMRhLPTxlWQdAcONY52ml4mKcvcXBUgO3m4tq3gNMxj5Y4Y
VXvd7J8HvBLJoon45IQgRtEJS0cRX5L0Bpc+uG9mHteiUt2jAka/12RZ02JY
i/c9ydomT0R7z2BkLqIvbdUJ73pz2RJJOErHqeCNxLXynqm3AgpDgH84sHGl
SpQ9ZEa1sNK2mC/MMxtPvCeru5lZvAbrCzPalEO22EJZfMZsSvcTiRCAsHdY
cJJ9a8T81inVzTn6HqtX9YEncQDQRsuI5T1vmPmy4XaR6i8oXeS41xZnVxsJ
m8cEeMEUy1BipCbKCWt0z8pVw+88kiMeeZn47xeqv3aumfK+4Rlgk2a677YF
1690MYegAv5yKh3MNuiHuh77Ko0dWJ8likzhxPVTFNETxxxmgL6bWwyRSwGg
FhnNgvQj88nPfskFM4CpyGstrJggU9/dcFD58dpMQPa9A/1DHRVS4QEN6h3n
H410BkhUpC3Z62pcQux5oliK3i7E/07KqOlqY8KW7S0onOah4phVVwMBocCm
6dyqEn4cM7IJxD2kl1yRNqPR3znRmU+X67Qwqv7YeGzrcu+lkHjUDdgTt2nD
QkWbkSVPezM8OxFOqji+qozmxL+akjnc28uLbFVqodFgPeaAR+H4FdvMkYlJ
zma7ky226v0VWAH5I9iM2DHCqQlLQLb2ACk0f/BeYWN9x4j3IOOjosK2iDPK
mSr0e4X5AWUdid6LUemO3ohrblN3lWV/gPnE8qiOJl+NN2jsNdCeLW9Fl9w0
CUMuohuGGUUEpoXDMU0tcwg85F2BBjnA+IBodD9lE5q7wkKxGR3cM3goA2CR
Jjeyk35KO9M2FIu2D0GiCeupZPCaR+lgDHJXi1S6hPUeNy8uEJ/fFm4jigWB
zIwcp311dIDL8le4RqxTNXj8O4pfQESTTcr9/r467Z2SHUp7X+pcI34ly7ZK
/rTktu9RyQ6RKGM/aCqd2CY1L3g5j1AvmK2kXFcrB9lS9hJNgxrc/MUIAv/M
2LkTJM8BQp39e8UcCVS3RsNbNz90KBQd6UB3T7XR/I5vNmf2NK68EUGJ2A0A
KdWgpKUgcYIg3+bRFUww1z9VGNxn2Eo8jLk/34x37x0bEAZ38COgbLiGcsAU
Erzghi7EuvhFoQIbN77n5/rt9QtNjUqjJY/HcgdcgYbt3KcyLPzD5iaTN+Z2
AGxm2cRVd2UT348YE9GPFxR24Z60DfdYc5mVBiqBHoQhcY9mqBdZPT1TS+IU
77amcQdOCUDGyS6k5xEnKPJ18eVH8/hbMNZlQOSL/uvwkYUC0XEYDs88UHGc
DFJN6UcbClTV9asyk9/4FgQuqW9pr7jhtWgKg8Q69iVFcZSzDrtjguA7e1PJ
tV7Kw8rf/8bK6e5fCIjV4komeOCp4FeNcYyan398QuosQHHQ9Pzj6FNjhenu
EDNFcW1VA6Ltg+9Oe+0HjUqB/Iwpyecnwazsprw2cYVX3kSbfjU3f2OzHN8U
BFXW4hfmGq6qTKx12WvJKrbSDimHjnFVYDZhNikEL3UOwLbCOEBEudWsVclq
yVzrvRCA7ecNbCiF+S06PwXxnAVSK6lFAG8vn1VG1KaPKOn2pSZvMqPmcBwR
trEdeplyIqvUIeS9WOvX1W3lUSIFDU2pQpqEd1FEMpntq4P1QuvhYicK6Q7f
r1Zs/qFVEFMLNLOx/V4a1may5ZhOq7uO4w5fBeDUTcOhF2flNdJuhADIEEuz
UzM6COyKxsPAOD/UFK6i6OcEA4Ml6l/uPP/UJF322+AiixRJCI3iLvDGXWdB
Geqm47pUUq+XjbyEUHXUgOlbb2OxxSY2OCkRN08vvGVgzSCNvOq8cFGwFh/h
nxiadtyuOkCLfvqTWZpYoINd/XA+y0mvTempofN7uxNCJEwFYU7ddy80el42
w37tqxc79Qz7aPyjRzzmkJ0CEI9TyXALI76jrZZNbA2TXTu3pa81nWxkKr1g
5dhmSG0OaWHmVbY+oCxKFCMDIfPKXIfN+AQHYffwCu9byAZo8JfQmeLCq7Nt
tHcbKUQTCcZoDA3uH+T44XFQdt39pPd3LXAgIL/OyLwLf8OSJFpGj0GDX1Eo
s5RYqo3zqXmnPDlAMTcjq4piv2GeYehO+pulg7QJVjyXFxW8+P/0gCFkeSXe
plMsvCpUilyFmiwTTIwzkeXBk4MQ+YGVeO4ztrxP/mF0borZUiW02vKUxW79
yLRQsRz0etSm9LcImkGO1lujqSSM3owopeogdKFac19f2mdM8FkIHzRwsXgn
0iPrsc8gcZsX9ajUxPRBP2WhPS0hvKHRBazYlVJFzo0IFUlI1rpw0WTWemNF
YNZX14xLnrdn/QdmbM+j4HiGa5IlSWMGPbaakl27xs5gMSphmqeWTcmJOH/L
wQgI8HS9hW0pAcLVY2SnTzWqNmWZJ5tq2hO2mYIf5FaJjhaO/6qeM17IEXLE
YyS7BPq+3Uv4GsKNRPjjpVFHfhy05zdmaJp97/2WjfEeehoWxPwuD6JQGKz7
ID3DXuca8ZVCeRFqhP+npNL/ZoEOCVwKtBoQ0NEcTQkOU9KfDLAnZR2Kvr/i
uaUKUoxeHRZSEn84kWRZbk24UGzYnoBPB14QlD/MQ8UsCU+ymbBmKAvapiSW
ysh6Na30vYYfeMSFO/XBNocCIdpmO1AYUepq6Kx11vOB8rEWBps1x3NtzJlJ
Z9aEMo2Uubp6ExIMBU/BqO0vM4mgSV6FNcH8b994+3lUntUw0RBGQlmOPeXb
JM5tCuiUqzrAtQmbmsTuv/5F6v4G4wc+uDYYv56HSnxwyZCxw5RAug8YVkYT
EOuJ74ovOvaxGvhbF8rQd7cGZueBmjjJUiQua/dH1j/pF5UMc+N+NknuGI4k
ygVoGkYX74yLRVsRgLsFTHlvLpTjrmnL0DN1VNEFs2XxeM8bvMMwBaHMomSI
UxyWqNIC7lrMEaUX/uG3lWpJyn8kicDrAe61JMFxvk7mZDoqwWP8NawDGL62
xTfFtmG4n9knN35fjBRFuv9h2+cA2akoNSq8CSSIB5koKLEWK2BJCR8+yPtu
ygStCbDNO172Yk22acsEQJJCuxikpir7Ot51MgOmzGr4zjo4zaSqZHwsVWEO
2XnzN3nOklQFwnaxFyayIUOdFpZpHy3rSjDASlvnGubZsqCXZydh55G+dmeb
jfX/tllqY9xw84poOuXkg4cLMkBTenC9l04P0BSVn2V6KfLnWEP4PkwThqjW
7r15B9Yt1LvR6nIMtbsYqYEYYAEYWCvSR24qTdxddqmYD409iKDDLYvkRRxT
ddyZSnxNO7VyRhh1CXtWziZeFl7pwyZt7v8ZoX2GCLc8++Z71K+KlnbddxtQ
Oxasb9jySn7upEzUVgEQlC5YJcRh9680HJDysxkAgfxQBCmlH85Kr3HWFTQY
pHT/j2ttAng42A5bC8aWt6zFmJywFS2z+AGlA2NRZeDCPOayE7sWmkuUn3hn
g9EN+LCMaEM4FBZsgJXDw7gSYGeop+hax88+3p8ItdJy4S+MbAKXjyI5gJgZ
J9GLcELuC7pE8qpvBdNxxPKqaEwQYiYuSQhabxSSE7+qpUScYI1p9NTsQFLa
zPsnYdkFZlvIzEZ6kMJJEQ37c1YWlbBocpO0RPCic0hYWPKE2gctNKiNo4er
h6zgZr9MqWmb0z9no8T6rQAi9SBduBkBNdoD43mH/mrOuEN3ujm7cN4g/GjR
q6MN/0MtlmbOSKJTTCGPgSN5s0lmj/TFsHwnWsAYqJ5xVr339ilIVlYn6XTd
xlHuyhHJGVNyHS3dE1+3bREaHJuPTPSWMv6UOLXCP73roRCOrKKKDwKih65c
Ys5p/JXiqI5Po6R97thrL+OP/w6zHOeF2MSSUNzBPFmMDmHP+B/UnvYoVEDf
XJBLoNdd6GTPYmGtHhrOkFmMOBjfyjahljNgZWUSd6iok6ynl7/d7WTMy7vc
YcSN74FBKJw6qinK5KExUhwvE+v93R5tnLuPo1qiQSIsoyvPk4+1IGPwOnaY
Brc+NqSejYHbMsvY6xWpVVTUL07D1tko20sXkiMmoJW7R3enGN8yidQDI410
DDNlrn3vmpHs8DdHw/am9ErxIGrE6gMxeVWVkF1dc6p7EKZPowmPc7a+99r+
efdnDL0GxtlbYCv2tyaQhR57LjiTPv+3I2AfNtCxJxkGqAx9lTWqcXy8foCL
qkC0tCYkL/oO46z4hwbXKb5T6rzijRKQ11rsepVkNQEvraPD1HTpvnkAWlpY
sRC9RljOJgI9ePPr0OLUy2vdUaL+D4yL2fuQMhs8U4oj1CpdsNlOUKLlm2fT
4OxU52kQPR5oNMOVkFtFV7tpBKyJCVJASIgVP/c+PbfWS+V7loySPTPI0cgx
22e24NFkb89hGU5BBCJ0WpVxCueUhJs0gJokRB6taSN7NBUsEP3EOoOg4AjM
HbhHAw1zZH31ytzfbek/OhjzfROqchhBd5iSaqIrkS1OhyqcQztU6cSm4T78
U4GmjkKS4fvRxTZiMK+W2fhSscmIn35gJq5NUwmO2JM7terj/OP4CsK+T/pj
ZU3nwCb9cmNXwCTYzXHR2VnBg4rpb3//W5Y08xv2jWgwYx8AuozqHnLIVuGL
RYbUf01LWPpeuOowSmbCNnio5A9Rf0o35DhKOINfx63Nbm+MjiSB3BY/O3V+
DCiW/LTPITu7DuRqMEl0hguG6vkg9gGDlV5czuW1Js02pE+WptdtgaDuv6+/
7FcsGSqTrfZXrrAqkg9g7dYh5jqkqRwv0DsCBX3uKYJL/ib9fQ5tgako1nKb
QOwQpnfMJZacCNbCh51LLMFbUISZMfjQHn2REUUQ4nhB6EnK1zdFED8HQQe1
9gI/GV2PR6xbxvO6S4gpwJ+4/DZpIpVAhgNXbzR0FionYOk0I/dMwvovf1p1
wwUqaE4W9Tn31P/+cYWi7D/ofKZi8kgxVigMfPaX7iHvmKp8CZjEjaWthEEr
mhFLuqUC3zEF/ZUcnVGRWl4c/KzSGGIK3UHMlKDvZuHdAg3AG6dMJM4vbtWg
BGHWCavI6z4v+8Qt0YAMWRGLKbs1HoKeWT2FMn9xHy13rs/dPHzpD7xGMv7b
+juRLV4qiFvBOEkU3sYUN6I82d3UrVQWiYpxK7ygzAb0SE68T4WLyebIdrMZ
K4p3ezn8uUmQebVXVYLXrM8NoRMlMpv0HjNSnCopkgI7Ls5ugCbS/ZTWmKT2
v4noi7NhL7DFNCNKMmZIldy9TQNTM4/qkZfPtOWoMDTAF8rXUDkNHGczTUmE
uaVXRXdt6hrUW0WnfRtMi2RHSWmmqAaT2uUb7sqXCx2uz5KP2EJLnQi46I4o
vWNr8uQTjlNOlmfZ9qNJaDXBrjMSxirAdd3dHgFGmpWUgw5NyiwDm5YFxOv9
u/7SPZOXSChKNxryUcwqjWHWcsG09Jfy4KfgMN26Sd+cMbwKU2PoM6lUWcFj
4lXwKJ47U+hRpO1HUoeiusz+fYA8PizubEV53ZEtfRm/jpBFNiEtxmYUcyys
WfDY2awwsRh9UMuLYeLGqdboOohhDRE5f6uQQxKFnIv+cD2FSD/6G/ICLc5O
S6An5R4W1BZQtNUI8jMwS2TF3U60NRqKwRvvKpO301kmVsqPWD9L1gAyFBgd
zOjGjRbytynfW38MAVbjWoWybaT1Y8KGsY7fphiOblD1/qlNDUAVBYj/Bekf
5uEp+j4QrKB9fQ0pFt3dlPtbiWUNm8APlATRzqFmn51d1wMjodCeAfq5NPe6
ARDZNfGYJbNBrswjYq2VcpMvUvShjcDNoaS/harhOMNEFbf4wf+cs6D0+bGt
KXmKclMZ2Xpdmvvt4TPQ0EB8TdQnbmiDFSqrGLtf4QfRugxuKjWAZXNg0trR
cJSlq8Q6FqSXJ4CzDQPnP5qA4Lii9jd2met/In45fx681PebgXvTnF9X1I9U
VLqTmI3vt437j1ploTE0P+hQDwA6V5s8W3LXFRDGZ4ZpQKgWXTi/vXNI25Nn
ZVRpGy63hEu1uaPS1lRMR8z6W5p+ogte2nyIVum4OfPPugOtg+1rXems257K
f2VjMo1rjLrZCAa83YdwboYXCTZpvo5NCApyUO9lMHqRPToAM/CGUIbX7bSJ
DzusWVouASUEjZD2k/a02snjCscip1bTfAy35Lp0vL7Qrwd0cRYyfx5eeHte
wl9gU+39nQv9hYoSLqK+sd3HzHJI8OEZy/16sHkqm+QNF20Q5xXW+slBwM2x
jU71Eze3FkABXojT7jDOM0myBxaRJyiEYH3fMKADoRsDBhBFmvG5pmfcwd65
nSYpOQfhcq9bqeNgzQEXKHTRqmBGFuRKhmqMk2483/uBzfms3qo75lPYJocn
NkTIaOLQ5dRpVmilG/5BV81+xC6MBPswrEUqBqtYoURmABh8ZSVSe12H1VZA
+zMY7VHGyylUstX3TH0YbQb9+dg+ISenmXQT72V+OY2Vtdtna9GFsoZFe8ep
fMOygpx/CnKpe2sny46mtwHKhE7Uecs7Pn8JFQovFNOpYsHYmmvvSsPP0cqj
KD/dgraUMn0OOFCukJzpV9efWK1iJi1RJc0P7ZAqnQywYj/UgX2vZtbaS0Lj
hWJjNj5to4Ywjo/d0BMiCxN65KBz43DtftjCpFnvaNWpvr1hM0myMrkgEcr5
fwMqpJ/TAFNsPR/0TZHhGRVhnb+A//p51PXioZ6jlYu1TkPck4Z66jZCNm9z
yCxP8RJNBD3eSP+fFfteJihn//02sf2ZGcjvXe7YyBY0PCIzfi5QyPBHC+Du
HRLWANuvJYFTWDv0uilT5cf0v3j3haMluNLq2mA8cWsffJdVEp8aG4G/30xy
auQW36qbEwZap0mNYEWTue4AiR+YrDcEWbPX1HjdnT8LayyqSbzUd9KNidIN
ayFvMLls7CPeCwaRtkTDM2H6cBfZAFc7ZQfZYn4WerES3pFIp1gt/v33Wuj0
3kZobfeADmowAXnFUPuy5i67z5iKCgTy0WVtGBJ/aNkOKq86NqmpFQRP+HB9
fiiFbtHobPeHhD81QEzM6zXGCrUmUfgGtPy7zfYMLJMoLi6Uv7c9PdMANERr
AxhVvrFB2OJvkz1pkXC5OdggKijS5KjfESO64A8J5/dqzA59zG4+FFx3E66q
Notna0FzEBTTa5bpOtrW/bdT8YWAQBUXyZwJY1qnR5GH6vGvnzTWfuv/mbvp
+B/SrG3eybYodB/vCbGPKBAYoI8YVFDxkqqZdeBk+ly7k04Xz4BC/cpUUbWv
i5uTxdwJTo/t3l3PseDz4pmB2rVuQUgcBaUJyDiVREDYVdzvAgqi2tZvaGPk
uNGFJkGNMvN9l0XWfTk1qXWF88shunAN5CwM8kg1lbPSW9zVvoA+i/vCguO3
W7xyENxNkeuqNhT64hm4S+HAtCESWcsM3zOpemDRHCC3DSFXqHyOMKJrbnqO
QXKk3/aM8brwvFHlI65AnTiSDYIFlOJFNBfRBxPthebTs2dQ7VbryXAFzzVR
Ph/Mq87Q7v88aj4QRLGvExVmdoaLpAVJOqrlYIXzl0ZHOklqxxp9YFgkv0TZ
Y4wUAeWtFdVIVvj2V7X5SxjrI7NCdh/YtGSNq/U34kjacBPL6DVIHgH4N89a
M81JpTfwYL+ufwoS8Oq/DzxkxIBVazHVEXmzaEic3SxLzRsceSrrPuquU4FT
PkfxtnjrackFbRrECvYJ1WvM4Qd1HVni/4WS2poHhHoLVtfMsPp+z4AnYii+
W1NmcQAUp9mY3qS07YVLjwrrpcCDWizOJKw5UKVYXNt7sl9mIO9sN5d2awPB
Cg8JcJtqiHCVcy0loIB+q1sUUNr+RBx/VOq9rxxJP2iv44yMsJ1cznhcROIg
jb2mhfPnN6QAId7Tr6pfd1QOPBqBvmkUxJCRka9E9GcYB0OzDKUcyeNeDnKw
W/26qQPPIAAY40U2ibEKXHbsH4RErDR3FQ/ZLX7lxxEtbuztKEdRtHier4nd
FDzq1y3BmJfdHDwk3TiUY5NcVELab5J7yFKLkaKHDk6c1tADC1Jb+dsULAHD
msmBxrvEoie2IZG+6hO2bL2fPPUPVlakBbl+140yy0QMQvQBySGSTcqm+YM7
u2mgGpTV5vEAMFGgmnhvlCvWlF/EmQ958CCivh360fJNjmyIHUEp6wjRncNT
ohgbq+BRmC7oPJxgZ/2Kq9q7i48CJvc7zvrVKTuXwZZo75Ub/uGw7WOY3ioZ
fTBks0A1NY5rVlWmBtVPOcNFVxuIKgy+6OyH39WyOMxsTQeDq/6bMxoQnwYG
do6KekC3WJnssLDgEa2oyK+pUFbcel19RyJBk9ZML417RmZQwEmusex60twx
w5Z863EcV0ZK8f4+AR2pBon6RQQxMJcLhiSGJ4Rhv4iF8iE0Tm2UhCHGuJ5/
Ayr+7mEvkOijzUJoOYmPdCQQP2iKtQYC/CgfuGQbEjEw851N+Gi74LCZ7F8X
18IErIgizY6xoZ2vFj+ns0aSea+LWvvv1mMnVnP1D5/qT+f7YieKzJB1tl1r
xl59YKdYTz7I+E/qDL9N12cj6XNtzYl1+3KD6su4kzcQHiNcWQwYBH4stW1l
YE9N3QPCW0hiRE5G4En5L8uaj7KldP1OTbHMRwDi20YB02UQRL6n5nU+iF4p
Oe7iaZC6r2W7UDUdb8yrSe3wffUdL+Q7MyWFxbmXoJ+krL+DwL3BiqyF0fri
hfJAxsBAMF8D3z6bA5mexxZ3jFtkB5wbFdam1vqVpaU3E/Ot07kfaFPqfgnn
B0QhhJ9c6nh7JNvSxkuchuHjVRnD0qba1ezUYKP/kda5CN0HRuEIEJTSjnxG
uoIM/rbZlH0Lua2k9wUuH99922qFr0f3chfjJn2ThyxcQrwkQMvF6KsihYK7
jMocmIcz6YDdfvsY4M908HlWc2edKk5Hq1RlrxBrtkUmFus9981h0V2+umHv
fjA6MIyzs/Rdl3L3NUsszjiMf8Ltx0gt1hGjmeZgTYiqcKVkGNtatzzl3Din
FLMkF1Vl+smtaNZTKR9q08eAzvVLNqTWWOYChjfVzYX+nJY2G/sWfZREn3es
GgGo+AoQsZL7XR3eq8lMIRZUKeOyxJFp1Xuw6Xb1R+gjQYwq7L9jak0JBS8L
ocQaOBfcgNwWNXaqFOxTJpgsn27DpWQZWLYJELYyuU1opfjgWLfG5SFk1EF2
Bhx4y1DXMkNWICZCX/jfejYzIp/XV6DTa5NVn7jDopxTlWsnbrPWQ/S//UBJ
pGWadZlMT/hXXCsBCR7Omsn74LCXEwb+0ObLOTvRsxtEEOXFOD6xr4AFAVCh
JGaWBSy/54EgsMjt8Zx3KUsSObz2pegsKfdkFT5oxrrjlqQZ6N4jJB/LiHMC
mqjI0mPdSeBB0BBIJw5T3/fPPHxBhxa4uYyuRpxZEDnmyjXxB/5gUe7rf103
0g63WtpJzTWHy23JpqRnHlW/DtNXknl+1GTGyKakMIzm5xALvLptFE8QmpHp
FBhucs2eusLCkr5Fyub+53ScCw8x9qaIK+0AW0vb39xgQfP9GKtBpRKesJx6
FzTMmiAXqxaKHY8AOzLIkVR9Nt9wBuD8s/kkBHRxapHLGiutiE9MA66OERa2
b9Rjo0f19bZO6OYgHpG7UBp/gFqeH3wcrhKOUrKvfjwLAxWkxG7cv439J+Ru
hCLai8NfmWb1qQd0wjJlTi/iCXROyNgunpZ6Cqt5HO037/qu0gw0Lm7ASPiA
WkMvDgZJXrExdCAZDaGh8LpKdTV/83Wls+WKH5vHBTOKNhZ1bk4Q/DvuQVtJ
GagjMlEjxuZzZYlYH8Z4TF4wBRxHnFA3hlNCnnlmI4hOwjibI+wAOSmbDG7a
ir02GIMiaM82MNjKBghc+uEkk1RdE/iOhG+GmkmE+POGFCbvD/li4uchnmCE
eweiFaEf1BLTzDilVgyBUuNy+/2/qLLSiFhlFxXWjamTm62X3M5t64ldAUj1
AAsLjmAXSkKJ13/40NOp5T7ypIMfVQqxx+gWAOdJU7FTtZloWK/n+VqCR2LT
ixtXJ9g8zmU+p0g31SX63xZMugkHHPGV3V/ijz1lKtRWYFIbzGIZhui/hd8/
I4zMgbkzRfFiRqPY6MieLY0Tsl88hs/ki/k7/rg6XarmCLq2B0THcNtzAlvq
gZ+LCN/8UKj8GDv0GfcBUMmJt9a0UR4Ke/mdiMgLvg0z2bqiuYwUPT6SAxwB
x6gHDyUDEz60+cgsK6eSu0gKD5rpzgq3gBD0ZQIFT8eTWvMQHkaN/hO22QR0
7mI7tuQJElx2TdnPtPLCCE+2GlT7YXY0adTnO9cVT5v7p6VsgbAprMj0nU2j
6qJCu9UYarlpN/SY4+UGvuIrpRgdifLKynjR2vWrVeJXydAJVxkMUVwUhu4D
4X5wDrzlxx8/fRP105qUFMOvWkxzNFdB3P/D8X70M8VtrrhLw9VcC3Vvco7Q
SMb8WtxFomCT0prlk8duwHj7OZ6fBHzx6Z3WIta4apdSMGzC87oy2ZQaHEsc
0On4jRzAjlGvvj7WNSZcBCkZGuuYE7cBKdbk5CrFCGFVKxCNlR9n1vTd24GW
WAqclEyyfP6iB/32FjY4qJvo1EBwCBVULEVLcUtNGRcOyuxfxsFd4WLoDINY
R03WwrgmMmiEHUXAZbm9s6UsxymLeNFGckSLKtMMjWNaYlAszP9G+2bwubyc
3iSmRMUH/90xEYLHKB7FEXpcUg86ivC6ffGfOJUA03aboD50wvjRIr/ggXHq
Zxggji3TEfAuY4NsWfW8BJw06eNhMUtrzfoVz1xIqzAdrQ1qTDaGdBU/J+3U
BR5Pam6OTJ3me5pwfqW48r8N8qlC0odWLDz7q+cgf7A0oZVnpdLpauKXfniD
8x5s11CvIKtT2HUSZm1MqkBV1C86/iBWSkY6BBnsN0x+atA5McZjmHcfeeCK
YP3RBjVhK6NT3qBIg8aPZLwFJAnHrPIVEatH6NyaJi1gTiHVe9os4g9Cz/4B
AONhJlFuyQzzKxb4bLYKM3kUlXycB6m2alX/3kXKxz6lqJCQhLWHH7w22cNm
/HX2ybaAv2VeWYPjOgDinYEp0bDm8E0DxHnIWl6lHeI7DrgfweN5ykRS2Gpa
hff5t1BXVUe56BEqUQt+S48O6ROXkk18WyGJHIMtNXLWwB0uRnoH60qsoww8
AHAl1niw2DfOpkilX8FWL8uD8SrUdXHAj2bydeovl1tb6QLdujeeFmMYjXOl
ge4SJviGGKSnVS2lGJF9BBrgXbG3QsVG3BxQvqMN+kRVvWP8Ocy++FFD/mmy
Nm0VgClVy2jpuIQWaCIFigfNgYkdPcKHg6kwMTHZ48C3F4kSf2bZ+pZtuRrh
qWAHrL5VRXo2EyQ58jzjmkfnYM7bOo4CanoYi+NiNk8aoXjdb52ehRHNtHTw
k3zsHcn/g9YtGc46SDlTKCyTKYmTRg50QSsugL1d68X1bNHZotqArNkVaKaP
K1MZZPtw8wjWOXUxdyd0ro/JtODDmoah1r0cRCUO4x05EzFCU6IODIuIZfda
hGFrFYQGFwIJUHBp90KrCVMWTbJ7aO/l7XhYfEG7x5HnFmfyfYH5xLShWTPv
5ydEqSctdiMtjWMqQ87XP8TVPdRTSZm//ljjzDTnoFbHZKfVLaTLv71wGnKf
2h0rlId9ArM+xk7rZV5gVyd/0oVoejk6z/zRzyfyOQlGvzchfMrfH/8Tb7a8
6NdDtWzPdohMnKvW9uizbJ6nc4MS+Sm1rvyQf5Qp050+1Ej5vgqbw8rdt2cS
x9fs8oV1wskFWmeIbslkkXBlT0+xXIw/X/QiAHOjInGd6o+bksSb4FLoszN+
uCnsvESZmtMRLmJ/VgalZukd+AJmaK9p4+1KLZ0tRyPnju+C9tmRcZy42Wvc
6t17j/lo3sgjaDasLAE3uSBMfXcG3bgKZeX6mgLhESpeFUibIEoqGCbPDI2f
ivWV1d4AzNddEjIt6QanR8+CY/ajueqs4l2SfOpHrRnRpWr9Z0cxkYcpWAGb
mxn4s6v6CWtTuTDw/4He2P8AGtsatuJhZyVy3BA4i87UkzXsAmofA8whw9fz
DziY8f0e6A/0aA1thyXSFiSzBickqgqbcalgHmLIGnIb185u2wx5GjvO7UO4
zdTY4FP93u6iEUyRJrxTn+h7XB8wg85J/DkDHUJ7YJvWuUoTaGlk3/X4YHZz
N/ajZg72EqDWYFiPr4qMC65Liien4TA59bFMqubZEZfihDd2tZRMZwrTFwAb
/D7hJc9a8dNV1Ore6KTE1Ey59bEF5aLwZZzxGgB/nzmwvGV0uiStarIoNdKd
B5dIvWMemCyDVfBvODac+7kHWl0/NxLtXSfxIGY2UDt+AZPR91HyIqfFBcZm
SK2TXdzJrOLCZwOvtxT1JsZ15oJeL2V/Q4b+8p8icv4zKdXT6NMwWEZ02ujJ
qHheIEX9cf4RQBf0AZh5a9uqJ0WkUl3kRK+dF0VxIz5F/g5hBUg7UMGb6EwR
rcUj8Jld7Q5aQ/IlY50VdOpssKSYW13eokJtHAMDy89N05roOKd8dNvPYStT
LwdVDk61m5dAxtW94rSpmNgszJ6QUO/IDa+fKYdqm7HaxMslV+FYQYxEjvvQ
tt/ttSozm8UBeocNUm9/FaoNW0gjg9qFjBy1QnVONXeVHk7IABpuAGXoCEOm
FSCQ07tESF8lAnSELKU8eX4EmxLP3Bpb5vecJi30Q8dJ93hpm+GODGJxCiXQ
p07KGh+ydJ0GhdPe+tiiBmGzAdbC5ex+CiaGQJO5vyPPapeWgRjg5CujBMIU
b6xC/Veb9Ofhop61qdT23DWwGE7ANVg/dMSDBEKKR7POgTGlPFuHWUobAalT
Q1Ig09/EloJQnqNcXWYeDHgrOFcazjrCHa6Zl2Ya/jSo6w64qLJA+cZdJFlm
oKicfWV7H5TN+EKcy/iUcKTMSQPpInk5U6vCG67X8UNk3VCnaKA5lME1zwEt
TVCSRF4FiUjDKpCJMPAyhY0y5JL1IlxmFg3AZ8wfJ3wRbZc0zxrY9uZRwXhp
xipC9zojuPMrhl6sL0+TZK7anGNwFvWguOOOfclJ9x4O6CpMkfR0J+H8rAi2
6aDtkz59/ucAtJKqwIO+pk6GtQoUVWBREPZ/NNWOQlhywMcqY+ldQeWouexL
Jj/FOAasyP4YdjpCGRZW+1J+Wa/EhI8147R8TGchzXs2U5H+Ebn+hddgnbzK
Hsi9WwI/3clZMJ8Zv6lA1S7U6a8Wy3G+DEWsLYNs1ZNsnAeFl6HhmDobCWIf
o6CJghXE3hNN66h+r3Tqa++ipNma9Dv9mplyk3BwphTgsQTK3rOPnUp+mj1R
a5Kp13Jv2rRUERaF/LnVtGNPh0o7+BhVZDQJF4SwbxCnfT1KKOlpheuHRcSZ
xCA4yDEjknTfQ50r5wrVaxVDNCWOW1mLtaBmzGtihyJJn6fd+3DupE/PZAmz
nr8y1x9G2Kfy1gmYPc/lzxzVH3xKKCLDR88expfsQLUaxLVhaSCdMpgjGPRn
Mq6GsPdDhpNNqxpw3cBVwYpRvIPJFvytBjDeD1RhxJba+6sGrVlETT3jldxU
c4yQvk0ie2RA8z/M3TK43H2q6ZFOAZAfkzEbNQIcHrJEa3QJ6hfGAcOFDXEL
80woDvvRfqFhJikmiqgQB1SjDv3tM3N+gCq1aJSOK+R8mXwQ4T7V+pkTVSEV
f/A2M2y9Y5Pd7cRCQ2IVNYmuIbsgNDcoU4H7NnUlsGjReK0tJo6bmaUTmLU7
jUlFTVT3sa6RU0RBLsbIA1yWJ9gqGXSphMlXwsFbtS/eXEn8ioVFMvskANwj
n6bpQvUKVycdjRTUeeCpa8niLlcrj75x8LZhGUUzZ9HAoqOscs2LFWzRhlT+
SxKnrd5olDuUeuwUTCt8Ta3R2f2hByB91xISKd+pcb0oUR6TjjnT42Wj3M/H
M5YtsJAvDt2n75o596aVfUYSkpIjs2fkX8tZgIxA35/EwBZopvWZpwHbxMsB
C3py8I7XvoZPdFtEfuz/kM+mMKf9MBAX4aG0oYeJVvCeEEObgRRAwDXUgpKq
x9m5UBM6qkEjNI1tS/j4WeAkHf+B14us442Swbmri7Cl1mclfOxom1GJgKLG
PfGSCs8n1CDz4MEUeOA03rojtVHZGdVdC8YyK4valxslxlsNR25xGuhAakTt
OXwXE9MfnKdo8aCrNnE4WkDJP1SMBnIsW+mlqz/Y85kj/6pifcahaLpezxyf
XsC7NtyrnLFQuPZdZy/qN0cVE3woEYbIHfn3rypWB5g8+Wmon2+V3EJ+Isuz
tuRSQ6u7AjoqDMUn4pZlZxuMqhC9G4+mHjNa/7fcqR21/7EZjKQKWlUM4Loj
bsctx4J8cgTPINnh8YF3v5e1ormeXT/7vGp5gQudYQe27BJcoYSO78ggC7/Y
dtkLAPVlthxcII6Y3lUT+VLyL3NtkcU3DQrbkT0WGNxNy0rbJ6uTAW1yVNqs
yFgkjVZZoZII8CJudR8CWmTGggSvEJwL17makYgIItYKuOS1dWiv2RcWksOa
tQtvfFGsapbtWjqsv9D9GRCzrTFfLTZQ2DFuqZoaGKO0nDxSVM64lK4NKumw
UHe5Zivnt7BT3REfyVvTb7O/DK3+K2eq3vIi0Zz4zPME48hH99aH5mJybfhd
cXkwwhQMj+wPpiBUX/I51CK9C+cidjX4fA1U4Hj8mQFdZzc8F5ouT2sFaKs5
Vf36rW4UyJyZh3dEgmDAz53NEFKAjIbBL0P6uaLcJij+ZdM3STrEezm+Nbz3
RC5koQclWogZzKPIvEq2EyK0c94YUxQ0DxIKenMHtik5rlKvTozg3Ty4rRNX
ALFDfGzrxHMHW6gpJdX2ETyIMLLaaChtnbcuMVToGvFZkdzklr4xLetg9Hg/
HbKsDCUSiS1BnQjG5qUKRx8k6qx9FKrWKHqY+mXvd+koV+l4mDqgeMFrYy/7
vDfA6tWZnRsNpxLgSjXnOQVHhTjsuqZB2NYj0ewfwm8wlFb4XexRVORC9/fh
mMMH+02jbgYVLCn5FexG93q110ouA8SMEsQZp8dlhPBZYqKyCldqXjzffU6Y
tHaOg/MRqarB5kJdv55OhbQXaASrJieLxaeQ3PMJQA90jBKsMqovCE+fSSnd
PDFPICHaQAFZHuwjpn2KGkpKTw3A4LLu2/b06kSG5fs6WdsBK3uuTPRMeb/i
uj4w//g3MmMvXECuNUnb8+UOl4b9R/Th14pX0p3SrXGrwQ0tWp6Nn/VFHjz6
DdJxAuHsb7sqI8kRIWsLZXg0UMZ0oG/Bs/o14y17WI+g/bAhyVa1948yZ7PA
oapl8bu/09iFjzXJTBQHwrz4tIzm0d5xO1k1os6JDSqbl+be/IMWbqddjMK0
MTRAMZmqgUUSvP5PeoDKs+wMJa3LunYLYjFbHPG6nGpP+BetbNbqoz1yh+Rb
9oLyofviiYpor+cDshiJqCuhplXwz/kOWRvuFU48jkxRibHcSe5jycx0xidv
RTwWJ4UuIliRgehIr+H2jP0Ub1Rwjb6vc0kpI3LYoQdO4fQBsXXL9MSbbSnM
nnHAXkAGM82zHLx2IEGM3WtHJgPRmGfdHQjeKR76gV2HzSPVTRCTdDGCumIT
PBf4hTLXWdDhTtbjD7enDUPTbpe2Y0lTjGl95kwwVYczWxDAEkCwgn1xrIzc
swQN9aWjva50xpm50Zrl6jVq1YQuaG3wvTzusKmgSxOs1U05yHlGnjKvkHTV
ePZrXzEPAX2V5kq3xgbi+min5E2zon7vaV5SeJovSJTSFi/m3OSzyvEoXCEi
6bjeMi5/LdlR73PLmhUPnLOZDgE37FFdDYTgP5uI5KcZb0PL5EU7P2awf0J0
O5o8LvXhcwxvjEKuKUPInrKeu5lcYlloZvVmwxfilT6uqo1uGMWg5Csay98j
QidOP6kMpnLhQ2CPZi63KIA9+fbf5zO/Yq1jXC6oPasakQ33RV8bpAtQORBO
90j2WYVe1kBLimthH3PTRy35eIJXrfCmQMrJynAOc2gpwbrgbgwsU9FlTTUd
/cI5IrN97XtWTE2pj197oyiaoIN8y9Nf9ED+Y8quwDffLtznwmOdtP8QqL5U
mwXxzx47LYJAfGsrDHpfEaC2fIpw/JbfCxIx6aDZC1WjoSjKabHMEgY0TFtt
Br8EYHBdZRzWre8mhrEHl6aNFT80ZkOv6vxOELEI1dQXndUmPFxXAZsQgJz8
S/7Z4WlDb8pwbDcyVNhEtjVX3DZxX4vCy7Tsmudxy6qTXXDCQJsD1HSnMv5y
ps9BmslcgLzwpHQ9RryWaDRFk7M1fPDqJ21av5pcXNstqQvaHe9SIZFpI12D
MjVkLiZ/Q2IVjIo6r2fy4D8KyeMrsRR6dNqX9vSWyFi4ASz6Oq084v77suxi
eykVCynOQetxwS5apx0vE0ByzAP4HwuQddcqFPBfELvR3DKXnRNxYlEqNxsA
A5FvZ61C0ALDXG5WLQ8emo7bHLAETZVWfsA7vRHhGSeTosxhwwsmyDf+fb28
Ag4meaYXipzfD33wgj6fmY6rYEs5AFhFSjPe/1FB95NBM4I4iQMfKqpFGOm6
a/Vc6xyJ0aMdxcEppFB5SqjK2RSgAOcheDTvRpzr5bxa1X6rBndnTOF/88b0
wlrRrUgkhsp1O1czVgIjQ87uW21QEDEHUl1lkh4xAV+3xt0goEpvp2NsH56i
CA4ZsZWGShcW3JBntM8YYI2YqZMv70lq6+Idm3iQI/oEtYhoqWEOrf9I57lt
EKPFGuOtkL/OBuHg+ccumTur7uB1hWGaFTHA5dPMMrw2/jgp6JegeOayIQJG
4N/m3i5XDoYRJKD9e0PXtxOQ/4mQHY3G7aowR+GEQq4X++9agJmy7djVM0ru
VFUCKx0d/puyaeZUHprbHQ1S20VNLMOcE9mwo0XKW41B+4Q2c/O77oK17mXY
+GUSS8vLeUvhNz7/9fJjeenpmCPULk4ZoluIffc4TY66d+nYBmjZLmW4MqxS
C9B4NyV51EYNrZrVuQhpnx28/ZpXNbyuj2y2IO2lAuz9JLlPcHf2DGt1Ucp2
Jsj3DAB7Qc75hsrmfcTZ2UDffbFNMcGFCJd8cINVQqMhC9XdYHyEGApaq/71
32SwBMz3b47dHTbR2MuZN4uPuQL3BsV4W7usv6z08Wg35Uzfn1p2hoYOgozx
0PxajhaAKYIH9kwpgPr1YBvtenCnou7ANqs/VssgynxVaA+AsR7uludJPbki
OYSqkObsW/RRwHl3ZV5YCCUkNUBNqzMQjE1kS9mpTiMiO9zUC4dX56uOdBmd
HMmByTolVu+kw/wGkeDEAZOwHqRF36EjfjuXWOOvA2T9nH1NPO6MyKhnq0xN
00gBrvPj89+C/9relpGKVzupIeW3Vd6a6TbdoKZmFpZfdzF/wnUPxd86GwPC
Uq3Ah2APPmJg81k0rKXBsrjxHvrrAhhIEAl15evvMpY32SyQkAx+XusNOt5q
nZlzoLJRZERxMqhXorPgDWYOTKPirpku/5cP3ZIScvFaG2AYPLn6SesyE928
CFbl4nWO1hlUXHB8DA8ZMH+RzqZgwSOrnvBTAzVsa97L2llaZ+9lX3c95zhz
MntQubuie0uWJ77wFs/L0jE9eK0uE1vfIBaXFESjjZV7K4H+/al4v00WI7bQ
YP39wANP4sR6nyCotP7XG400ViDjEkvQpbrJEewV8KVpU3tGQfpWzCK/u2kJ
6unmqLwT03V0ppeTWWf7RFJysXWGOZb8HN5r1H7JEqDwVhwT4Ru11jYw9WQc
/STO3gkYbYmDAsPoo7skIUMi7iHCxxbIUuyMtflgfvKafwpnfbZozGB63fYG
JlNZiDo/+Jpbylwje8IcCg3pYCpbEhtZENOc/Milce1U2hT7ez58JbqzEL0b
2CrGdJP5YzcCrUdec9Ua0OcqTvdVvSCQJlRAUn55Ha5nLEBRAqif8JfkfCh/
UNn11JreBtRIHAS5t9Zd4Y7k/S0B/CkMAE8Eo6XKcRm/k9x+syEcAt4V7wYp
HnOSbUbU68mD+geQ8OIx25sC381qdd+OhiiK0hfqScjnYNPlzS13wgDb+yFO
83i0Cg+3AeTaI7k0kAmWwHBHZi+ZTqojXcVkqO+OQTAry4ixMGN26DLbNvVB
kEYRDt0GXiDoYsds/z/3Hjy+3MJS8HG3RbZxRw1qvxsCDyGHct6dvZI3HWPH
cSnUVcUVJrfWZ2/vdUQaf+qg9JY0VMlB+MZhyWKYZWARQaS4pk3PcNncToZ3
XodysZwLYI9D30lgYEbD5v4Uq9XS7mem8qVX0t+S47x8fH8GzynnEsXZkh1h
p81kTj1WRpVLbOdvbwsrX5/PqlWsqDgxmxXOvc4MsDBjitkO6XgwdsSWqK2a
Rs+7c40uZdhV0IaM1wmE/f0EFHAkMtlFhKc7U+HlNnkF/4UwJ7UGkvSujPZE
CnJRLKK/rXRwUvdznaBgItDQ0CTXHjIYUHrZ24fPewsm+1pKolRmVjfgf6cY
liKwLDL4iNkP9SyGHYv06h7yNcwM0rQM8aDLdX8zvSjG361VQv3R1GKidiEL
ygTxey/o74cfD83udw7aWDA59Zju0frl1T8OF/cefOZJjzs+V+6ZxmMXH35h
ZvMp8GLPJvRb3bEaNUY0TlN05NuCMVJTGpZ0+63X0WRbXw1mGAlZfOcSQV/+
yixFf8/u3KAxhr5uBm3LZsMLgHh8vvzC7vVpXJbJ0KY8Yv/V+/TwrC3BZac6
U3+f1yxj1UWRKvgLr6HZWI5h4dHrnffvc0PiUi70O7jlE2Ny2kAplT5tG+YO
rGIj1KEWhwlj77j842orOHKUorsWjeMwUg8ERKW6nMWQEoMt8uoGHjKIqZEb
MbAkuXGHEqTIhgIZ6pmWv7rlz08Yx2lugrSiSiU43d0ZJh+6ab/zgJy/O4MN
eSQoneSVTw6rcQQShSNg4fbyGtpZLt6sMmK8PSZRYcBJyCb1gT4diOm6KzbL
QzAeGEfLBGhatAmDLKfz+93ccVMK5eCjYkeg0B3gidoev0fe8tPxFTz1vqtU
V9sex2fVCaRC5z/Vg0og19M1uzKzYfl8gVEk9hHGqJjBnG3+u8DEzxCeRxre
SJmJa2kcd+wmpZ9gNYUZ9nwX1H7VfANs3kHl1na04pq2YE52HqnzliT3f8Mq
pO6mnkaSkB0NKMtpDrLf1dtDyd8ABZ9I62RElmGUhbR0vbpsb6dfU7DYgNL/
9zH+Zth2gaMruXD6V6RNB9k/wt6KXoSTT9bs3f+tFbJSAMDK4XxXl+XfKmAq
NZdIL3brRD2QF+4kq8yJG1gbuH5H1kJQ7qq81zOqCfnWfWBKSQl8jOwrG2nF
BQqpLC6s5o34IHv3CeYw9DheO/q/0U8QgjnHvrliWRsp7/noW7/N+AhNARX2
HgRqtX50mLdQGWCEH5Tt9PqCq2xYJ/HR53IFEOg+by6m5HMIhmGXtSaQuik6
oawhly/0jSdQc6OVIaiRRiOERemE4n3H/OwHvL6XxOhCY4O0TI/Z8P+9ILEf
vxcvNkd4cuQo6jAGSckpWRKSt36VndZLEvrAXSUPdP6EhWGoqC9nW4OLwtAk
tYryhRfAARR4hWuEPGSzfrGQCLsjZ9kwDbryorGFq1hwq+RW9hNu/xQFB9hO
1BmIVm3bX0Np6BScoYysLI4nKXMf3NZB5vfg8zX6Xl0nXdQqQo5kiyi5Ad2E
d3BYl3iZqFqJuwJrU8Ju2EtZkr78Pc7G9EAvMQWn9np9+4JLp3ti6N6miAXX
QKhwV1cv09lo+CGSybaWIWZ7/KtqyarV55HPUifygx13PPED9yeP13dpJ1e4
yhNwC9s2qSOFw2D1fEQe/Yn8oOSgA6cmZyNcCb9+2zsTYXScJ/g2h2NB1aq5
tGAhR1SQfHr/LoxCKlnc1PsN9pHum0pTcOZL4DzYys8yQl9hzhYNV/gzCXXZ
zyyqEWYgREHYTeMCns2JI0q9qHmrh7igAHoVhqhQx7IBNEMJgN8ZXUjjcBgV
MiKtEu5qanlkwuDhWgBDHqNtS3V3+rHVcN+lmu73qO8LJGlPhB7FKK0n5KLk
u1mK4yMh55DjGW9ywBineiFggDMPe2nTaoHS3/2oHGs/PHiFqYdTIkSFChvu
xZuhAOhFuHiXvtuDgdsU2dSEKdHMQWYgwkssCS+5ch5m295//Jy6l7QgelHl
9S7BkWqk28KiGlhtbtekv3OquhRYnMO3K9ztSaVMU6yzWo5mrvdW8Y20RWTL
IwDa/N/Z6TUQLf6Po6e+Gukb9G2Kqk0PM0+1r2Elpt56meWnAS8hj1mwePq5
XLP50pK0sJ4q4+1BKnl9I7yzdDOkw+hTSk2DJcNWWutnQs7J0va2h5/+xVO4
4yubPKgUh2/Q56FdanYZH2WyUb3d4eat67Y1DZW/m7JY1LrSxns6Tz+kaP81
QyPkrmjKMtLtDBpuc10nju6hyjhDzN3wpJbW6Gx9Se9l+/DXdUKGjg6ZLd93
AAKwwTqxAThx+Z0gQMzgs3jlsxQIohiWUBMBKybO9+GP8Jyiv6hm3R2DaYcK
Dmh7XQqCspBqgZfliOEGswxYCR4IGmSsapoJp3COQ5125FUDKM8oNBmQdEtp
5Ka5DOP7pSItiHpOCq0VLIi9scU7rjPKWT4CL5XbzXDqnNOut/94SQKbeRH8
cxMYopFESCJ6zFhDWGe3o6KvSVW1hwUJTxI1Vp2tl8oiwf31oLWE1UyYMp7b
ppk3gZWnSbaj1PDxjKLOel38dRsPgOdaKdLLRTnPPECbxSBp/+FAZhKvcTHt
UVLcXFaCcoufLAGD06vH8YNHDAoxK+Pg1vbuqDZmTV8SYMDuqXXoaR/EQP91
4fi/5BHmMAEuwilFj/mK6je0WL0QsfJIrQ2xEVnI6C7E/CngkAlXNZjq9/5W
KIdslaUyiXM5x5puRWtUXiK8LUF1MJZW3YXBJ5K63juL31MtU/83TD4QP+gq
LE6Ok/swGaMgJGiXAg6Zgep1B+JMgPi+2rX57wnwNJmOeRh3B0GPbKjsGfi5
WR5armCltwkRJhnB2NzePGXmQml5BQZ4etfwRgo5OzKoTprzCXFblKfTWdo0
+24RuM7WhSOcQ1S3c1zqd3gDiD2MOCCAVhAJt+QxphzGncao+eeZzkk2Ohhz
tOAVBmusRAJJk8F/mbzaOZ/obdmfXB1slPBkI5j14mupxhiMFzXF7PfSl7Rc
Rf7WjRc21i/HuBi1SbFIwLlXUKkkIFyhzrJhJgJvhrsWNkFUi8zIgowv1S4w
p/VLlLpakHmZ3p24y1pSWDFnrRjbnaAd4U/nS2CgEXQ/6ZfcBqO1KjHZs1Yg
NC6vZvPVAj98WyB0dJfBGaPyKeVkPObOUN4Wbq5WQRSbvu8JmXRY6SYdQMJw
uksRzeoFX2gLoQghIpH+zdg4vZ1mvmMbEvMaKE+yKMKJ/nY/Crs2Oz7JzzsH
meAkcqiCVwejl2ODubb1rQ8ww89GG7WP3klp1f80eONM0hml+jRYKpnV7pRC
BpuXeRg+t5QVQJhXErBfI5409ZMk5vSNTV2ZT2ajykAUXLfdMvXMBLnxxXYc
ad0rD0+S3rdYxYOh9nS9k+dUtfR9JvxjKAz395NhVVkccDyXMGbxT24x51p3
Oq12RwTiRnh1ziD55eVB8KWZcrpvXpI04E9f58Wbrb2UZ9a29AYlLrZixBDy
OtDLiW2HuTDueNtJ3psRp1uNYpaUnsxv/4hn3GDih6Hd3uPc7kHt/1KdVT9X
LTRdZM3N0tcJPODSYwtf7V3J76vpAtoclqIKVPNqcCizfnOYwYxIWbaZHWc3
M9T6tn6gZ4WMa4DVRD94qAQ/yoQaJ82c6SJE6FMQhJ4/r3K7v9sWc4qVKHiT
DBvL/HUwffFULzhASqe7bPj1j758mouKAGatNpaPxLUevrQtM7NRCd8nBfC5
a17aRRuj5C0XH5EQKp2r2etruck8k3t1yT4tM567bzzHa+XSkrvzhAsuf56s
HF99gdJDN8WxXm5fmpL3BmVIxLPaFrewA93Qtdd+ly1rCQVRBbzQlXEFCflo
a6zl+p0rgDmwtDUhGuQ73Be+j0/UDU1+fn9gCzu1pgTKQ39u0Eo2+SHoZIh7
id6nhlrVucz5ivvw/Onzn4O7OYX9KTijO+coB7T1VOaCP3/p90hKA3MBTsxo
htwpLyYabMuObvw2otkZwVyOPtsPl9+4zNyQxA9SndMA/CuJIKpJmDlpQNMp
01T9bLYIv7Pg59L0pBBlr8R++Z955Q51mmJI+S/21Vgc2IzjUzxElL4rastj
CrA7J6cTC+655kuoFwC2vPC/T/M9ToLugGNReRmR5Jna+uL/gepT6r+I3eJS
Sp2wgekUuR1rok/u2Ixny65PYLzhRKq4oWJ1I2UBAPckEjE0ix/gBcwVaCH7
4xFNUNs+SEtAWlY12atnp3mwamMd04sMJQl35oP8cC8xwWTHYwMbiCgoAtfO
oqBgwH4lzcZJSnD3BcgJu1mdH8uG3ym/HcYpkoSJQgI8wB96kiQ3ykxBnA0T
Xy03tqdDOIR8inZOj84R7KKryyBp/xF69YVhA+6Y/JOm2g3a8acU0nfqiFfK
ZaU+9lHWw89KTcsw1Yz1V9li2AqrTI+RRYxLgFOH9X/FMbVyH2BFkesgFrG9
YX4HmyXxzaf0uK97z/4Z+ajIvKM9BiQiUjNCjyFjV/mELIn0prizlEjMCbpr
lCPMHnv+3dNZcKhMFp2/iXSOojrPQ1z6dPC5ouypTR60iBo3oOJchTV5bDbJ
NzmGTUxl0QmPIJ5EMwpyXSclYh9kdQd+bBtp4I784HAy7M07QHnkDx20d37q
cS1JGAZGXFqggTp+rGr5fGUur0PiBigkpwR4ZewNyikx8pCXpLiHuLquWzN6
nx9SSgv7aHmAVgbKEV1U3uNw/jBCzMSxKqzwuU0ZmyVBf+SLHnmS5vRMtG9n
1nGCacqbWXsUKpSZnMqojHFpNM/gFfEXqTXLj51K3KvwQVDSlEUFoHQycN6X
qG+U7cNfmd0b2Bcei75G5UvhqDXpxATVSR5xorqtqNRBzqlMSuqq+8WB+pb2
u4vBFSVzNlaoWtRG3VOZAg2p4CwGEpBlUcWQzDPRk3a5zxIoe0UOFco6E1Uw
A4Xf4Bv3chya+Rtl2QI/7VSYh0x4tY8UMRqW6aGR0B9/KnEK57NhDkOl4fRi
B2L0GulNh8kBBkmN+HSkmafq2PIlq02SJlokYMKwUVX1TtGGWqRKfYbk4pDx
rfgXtuo0wKeQVvk7dBzoWWH7xPgbsLc3W6sM2F40E91gJ4F5F5LzrKISpQTc
BzdjtJllcb0q6m7Va7TkGJgQF+1cdPUOU2K2RHMi/eKEUayKaiqEV9F47RVH
mJTDwCqZ7GyBhtwTARhaS8p3t2+17rwKdykaf57pxRETCOpjQJnfb9odRMpG
n2ZN7cbfYacPQ/t0JTwcJlXApG08nnjuMCf6M+xdZY1rIlY1RolZnGw55+kQ
79T62yjUbw29cOPIrON/tIIQMk2m+VHax86XPPQxWAQ7fbGe3jeGB1wSqaas
lFGhu820oo7TjsK8UObQT3Hjpf7aBn2IpRzHg44EwfYTm5h+TjrHiHm0tfZJ
sdf4FSbLzENVeuByuTy/JN//pL+YL28LDRwz6dWW+LqWfHHvz9smRMUehmEF
QAjptOY8qqhFCZGI05cQAH9ymTzZpuSJ2c5G53Q2wGA8yZwyxiRjzAwHKV9Y
q/X1lzgWYN+JzO4Pef7pDVCzWs4L5h/mRFFxKro08fxhU8wRGTponB6oOZH3
E75DrdL2Kl43ZKvj0A9VTYin20sVh+GfkQnRRstRHEBEH+qBhuvVRiTrZvBr
f7TTa/MsolGvQV1zAeAMxSFzH9VprsLK/Hi0t51buyzfqCLo8f25BS4R84BH
IhB+GFT+wSSdtGy0ZkBSQQgKwJAsAI6debVEtDpN7SKY5w+ecUVBGz+LsGS6
QdtCqo6YarcNxtm+lRyPqe+RUaLdY77rDJdPqd8BgDkIpSpixhhSm87JuZRI
UknkFf4Qp3fajSwJHHYr3PaIf4BIcXY0X0IaMP90Ep1ZwwNybUA/2tvjRSX0
jNQy0n4xQlJCeUiXwOAOzKmKsnVKmqWOIximppYpekhTYbsVKLvvZtNZNhCz
UmPGi6BMD7QQg2HksrlqbpntjmgBevP6xKDI4AmFIutieOkCuwApCHOi8jnU
C2SL6je6tisK+sBN3nDy8C4NKj14eJIkVBWa6we2p+mmMeuhcBSFhTG5491f
L1XCId2CFOC+wP3Q0xypwqkjnFcCeh60EuaeQ40w2fR1X/uD5WrLldZGnf4y
X/+wBOz9JbDmH5LkWupnTF/w1butRvTVEj+f+Vzh/msVe0huu9CL1u1yHZ+B
RYBm5gScqBylz5DD0tDEfWZNYrKNotHmEGH+OkpgvOblAAiJK+q0UmAHg9Tz
IArFhh9krT6xDYtTxI1zr3KgD2kzz3SW8kR4ybjb+uznawJlFK4Bg0E8ye0X
PNk5GVKwS8fNABo67Qp0NrUh75CBtyZdDReflipsMxYtcCS5zVWahZqriizi
NJu9NUwaC6Hx9yb6MAOQl5pcqMpHaCtv+63W2EwPB1Zbj2pj9jk8uyrDuFvc
rDm6qRVThBTeiLE0hird8Mr2t+n7enIDO2A+JLuSkK+duwoxaPbu8NNUlrOK
PguAbdFgSrpgYo/nYr5KfyoB8CzBD0bh4R5FbxX461bJ9Xk9vgaPB9OZnVyf
DeZeNhe5YgQ1O3AI7eVhzhO6iKmNbgItmpZsS0vjHyu0JCMqgJ39lJbBeX7q
g+g3IO5cUvZdI+9WXEzJeda+bXZikuKM18C2EUTPPcRjlPUqtMz3OC1X1tRw
M39xT5VprQ4ftysG3EPifG0IW7v+nuCoeR+9kY3WFwPKOtGiHkXo8+eoRTuB
reVEMFRFhknR7p+WHfGJxTopNJmR9ye1TkU9El3C69pqcD0bEhMnl/kBVnqW
q53jLNA81Z5KcPYTZFnk/mO2LMGMIshJxWdSKbkABQvAFlhHwA3kALKMtECD
eRyqMNhgaDVPJqcl+oLc02gB9SI16kyWn4VkOB/5jmiNuoguK5nF9A3vJGEm
ei3NaIOy4TG4q+nHz2nI7i5A2qUb4RbmTxxb0elPU8HmsBjAnKZIFNHMbqAI
W2HlNDQ5mQC+54Tzj8mmFXcKAOF6mXfBeNL4smk8FJ33E/icjpeaHXhFTYKJ
AfCpnIyT/DXkm1SopNYUuIiZuRsijx37oqdi489V0oUzLVE72hozy49BNc9R
Os6+o62zq6SyXQllaUk9YjRt9Q4N6JHhgb5qt3ZEKam27797bJ6nJejy9DYR
HDfX3GnM6grQa6hY0ziRWTcUAgPkNnFXbQuSl28Y9onWsld/t4fK9Q+10NTY
rZzf/XpSxao61fC+fMI97PI064IkWvMNbGR9gnw7vnMK0M0zbmA0m4u7WrJz
lmsI4qGCViLOxwOe3qGvMgiPiZ5wGCgfBNP0Dma8ZEK/08r12OJJmpzi3PUj
M86734RoTlrsjLSDe/AnsePiDoQ+8Et2F5iluYQKeQEm+TsbhcH6BzYRac6A
UxJsnliBUsfkpcLQasfOz66zIUCcJWot9lBrLf0HWAunvpMPwkAGF2bbqmbe
0o3DWLYL8bEeAsblyK5QyVDQj6g4Q8VSbCFhER7wP0IKYCmXzYwFfzlrCBEW
jHQ/ZtIl4XBa3S8TqHnVFGXejCczXjO/HfvmZ0lEUUiO33E3vuxu39cG2o3+
0jyfVqoXryujPE+FgbkTQL9MlJvUMXa3kRBqB8/3HHf2Am0jtIvX1FRA/714
8/2GVR3b5eX4iQJSPy1dtkkorrv/jeJp/wrdu0ryXblV8c90undAEO4ahsPw
wXUIT+ciEidGrVygvsaoU4ggSwgmRcQ95ptvPhnleT4af4QZAYuy3piytHiK
66QZmAUkuCq7ZNTE1SH/6lTmvhOxqZFqtEPDNbz5ssXX/mk04fxMMXIxUX7X
W3/RwNUS+pAbEpwpo/5MJwmQn0i8G6GMQNT32U3yom6ffl8xRFv7/EuOx5Ei
CWJDrOoxmvvjjLlvU+pBIKtlObvQiJA8p0Uwt0pzYiPo6tlbD5oYaabVRBIl
NLc6KTIOxXF3Q4/tc4db42cOgyEBB7T0BzfzFJGOFlBOHwx4SDggE+51M+ue
0hLsPUwseT+LQneq7xeWjqG7MGE+v5LNGEWKikvoFcJKrRakp03amdMd2fRj
RdBoiMn5Afs4WElWWq90f2Zs5o9RXqN3UhQIffKe4nRvaeO5SkneZXneJA+7
ZtPekhnpTzxRALU2FpJ5GLaVUJHgsOxxUMZ4qsqH1OdoCUAXMghmBB4QJX07
NTGDEW5LHWF2GR8OWKCzX+i/UNbw0TpQ2RIo1iTE0cUZfigQTJ0EMXtrCplm
fCqmtkoQKzpK55gss2bHDjSt1cQuduwe6a32JTsJgvCbkXebF5+dRoisZjw/
AQWrfm9hFPWrs0VWxvACm8++dxNzwWvJD1lRfQvcvHn57kBelxlErZltx/AI
G9X2zuAtkWEmOVs2OcR0dlC/lWu2nrAp0/rttPA5HYT3xctvXIlKEnPSUiof
k5VEVJlCVV0+9K+149dtx+Eqmrr7GXiK9R+wI/Kpznwfun2RkapNDDufit5V
qz2R+2pcCAVDCENPKGCcYOjTD8nqREhfJBU0UH0kTpzf2BDwSCes2WVp760k
5FtOmYUig88rXRd3MqUgOVakLUZeW7cbD2xfuRRv+3moWvMKF+UWY98sgIVD
d4bRrwzBAOv/Ato0ijs+M8Ny+wkWGDKXHZM0Rw9fTSJWMt1HXrMA9HRUMEy8
BeA+Smg8w5mXx5cTROEM5HmFMBwcjnGVwekZyIk4lZP8h1+X/Vodmz9yUgi1
oEOg372WjM8gSTqQHIjWLQ/ilOigQAMlMx0MP+G31PwZczw4o+4mJJi22E0l
qHqRnn3Zwfk1ONqmZT88SttVdGY7zoEdwHCQhu09Ccx0Huibtzg8TJk/E7Nk
VfU8BHqNpXnGY2aSQMXqGquMEabR1JyljkG2AW91lODGm7HObrNqsDTRW7V0
LLHZxwnR/JRYrapKOZUlh/39chiiPSzwLOm9XPTM4pl0D9+4roa7cungvcf4
kqSpBIvl0f+aogFmXOEc+YyCZw0XrFX9O4jGufXvCgwqu6wcQOxChUk+17WQ
DKaKQtFeQ8lyUcgQoULfA+cNuTBMXqFQCDuHFG8I/cjstgpSIQocB2Z1GzvB
7D2kKx54Kmpv4hDuzI2ipUJpknpvXHK3jVz6zvopnCiOPh4sI5KkV4JgNheE
GIkXbMEnwhu4yjMD0MsmxesAKfp45oA4OJs/ndU6mNNgEzrsrsK92rW9DDJt
3iCz1HbUQ0bmET4QD96rVVEVmlZJ2iglXsCQKvRLLcR09sdEMjbMW/Ige0kK
WVQX5w18Ko7DjSujKc9SYZn1564N9JXka2aqVO9TY7q7gQ3OXcXnVjMN0EgP
UV31extuS3lBEZ/VHq52tjpp/uVNGg7/jvLHhFzU22h/REptl3xskHpYgS1B
RD/R51XunF3Co1eIqGCVfs+MD10DZbtkr3Z3f0rf7DZ9hdGenM5WiTMTUN4M
IRJmmAsfxLv4GGBYEkmoYqIHdofG41SzX81kw6OgMISPdJbf7jihKYQ2ySin
WkVKtDDHCujHiRzNLnOV2Oypf4imw4OKaxPzrAR5ppdKUt4A8V578fqSzfEq
pvH/h1yATdgTgkqnFd4gboYiGoluy9ZX7Ve3cxmC2Cx6wrg6m5LFBYWRkfzO
IiEJi11qLGVAos8Eu09cyh6CgQkpNoERNvJtTSwyImEaNKwQVEa8i84pYCJy
KdDsSTXJHEPg8KL13HAbTuffsSdwSBhV+0UeuZ/BgiOKwQ6Lc+UjRmxpBUYc
wy+9khuDsSiLQ2yKTfX0MwxM47bVNvQEJncYDqGVGbLFccM+vv5b2mKSjBvS
3i7zXJd9FkSyruB6sx5Nje1gIE3i6RFYVoTAStA7XncypSBFG88BWlv2bfrE
i0NSWXLPQkoHYuMWZh7P6MH94aw42L7UrUS47HROl7PsJa8Y/XR8RnjJvLJe
0QcU9F2mbihsoch4eWKWStAeT1H52krVFt6zHpsPKcSWTZ1LaKM+d6ExRZ2C
QaV8AjA+G9yYtJxepxngllqgwtGLk9DMU0uObxxACOkI8O/3Lj12k0DoQcz9
OpAhSCF0YPR5MBr3uiTszk1e/AKjZpHWUkFvuQuUUgejawNonscMecDhl+0m
mtZyUWkTTOwLfVdwwS+SPjqEsZ2VNDikb1SorAIKuWS6R+VNqA8IRb3aCXW0
HjRL1iG9NiLLF2dE2PEv8k+2xPIK1r0cuLiiJiIR++kCH/C1xJUymyPPG6M0
0XAtw8UL5TQjOHzJpaZuOGluLfdmELGXZ8YNhlVJRn3PwRbmsW7qCjciiGX2
AhGOao77JMwsBDJnVIWzFTsWjA6b2fH8vgY0cwk7kA7ip7bHHjYIuDunJsOv
VWaR9ivBdgwHtPK1Az0KoAODODUIdkDXguL1VBRxHcYK2v4zH/es6vFXiUPH
KxVOMZRsT4eTTnQmCRlOnEwkZv2QDTe269w0YLMOX2H5smWHfhFz+xiQ9ACH
4s9oGst3ljqF8jRSOEFzKWPNp7qAfwV+EsN+3WWu4DefCfyYkc2Sq70ZHGRL
snq/kce3yYb0Ncv3dNafivzEO6KvFW7RPKn9xUod7RtUfl+61ykBF/Iml64x
+an/wABkWhHBMQaOVpd/kK4W/s47w30Nnbml6MObqbQkwZ4UeLJXaN9fYPFm
N7QVyZnCrxiQe5/FHKJweWxfL9nf78lFP6F/qIkmNaPGePKWTozQJLh0TgwD
o8MU6mXpA6qkBrSENL9jgPtEMzGxRbmYwa3tdWyDo2ptCLDd894Ud2vbZUHV
fBq522kBx9HOX0i2ywLnhb/hsNvmOJbRRCXUlXn+QgTA5K+L76nRdi+HMIha
ZfSewh5iu62sxdMssKvNYxqAdqqxqpxKfDrcEXgk8Ffnp5a4beoivwmXvdMQ
vsn8x+oEESJkP5NPA5uzYxocGZuB7KV7pFVXPtaFcH/L3Ut2UCiHh3eH1XOH
cy6F66AFKJbGbMPZWy0Iiwq3Ruj1w9HGzF9KydPk/VaBIDovYOyYznjjuQLf
pFpjUeuEyYqYNEHmI5hL/2srilSdlur8jhyVginv3rZCEUxTokGe8oTMSPPV
6TnU1fmMBdtF6ORmBWD17P1Phsm+igdP7IrhBFE1ULb4wL2o/I4DiXPFCGxh
zjiaL+5lUBWfb/KIxA8K6/RsR9t6NuRdavVWkBTtUSrhhbMtp1rCf8CNiFdX
LhzJkhpJWUuGR+ijWIZwcaKxsxf1KIY2AZal+xZAY5DJzmAkpXvFRY1nEd+1
FfItD3cUi7+D+6uENL/C9HMgc5PtWdsvwQOUbjxO9BODgTowdQjXn9PGdUqs
YhCKUlvChWIeOihBNuUxdnEETWWMV+FW991iUIDWHf87B+zP5vI4IEOCNnDB
wRblKGI/+PZBK4h5n9HSUrSm3XJsjWzjQT/0cLpYTLEniO4+JJPKamcgad75
9FkO0X8FwRLfY/o4K/SDDGciMkhyXxUOmJQzPU2mI+FFQ2Fm9vGc0+fYYkAL
QzTk4piBN6sM3dVIrtINNoDl6ZcKStTeziikXjbWXqKrf9NdfFHM9ay9Fhbj
SZgbY2yFRQWU1pggS9aPLBlOw5Av0z+Q4gEVRO5ytaKeGSS6cKHmJnSFPA0D
84CKwU10OFweXRr55sOHDPYSxe3x6Ru7Gji37j+Sdq5hxSJo+g5/VEb5lw8h
5AE1QMJz6jBrlAeKEslhamq0w83E6xXLK1qSSmZlcmPlzj+Yr7aKQeuuN3L7
QHKd+LmV1zHCru/N9f9QrLm8c0L6T3mNmxU9EKS/kjUEIvXw18tx+W00/7z8
N+OpIHdKUVGWaHesbKanX7evQ3KwG9oTPJ8/OjIN+Ajw8hLX05FalrpXedCz
bRgoQGf/0/kP8huhyqsCNMMY4Q4Q6vHNdSMYfgdfhEJWxp+npXlp3M/MK/ZW
OBQHsczk9eXPJA2HyswkuQQ5nHo96pdm+GWq+v4wIJOC6iNGpP8u6RB9sqB6
Pzn3Q5n1j5VFbOUlkVVbAGsUMMOy+QcrwB7IhtoP+4gn0Xx2o29uofbiYvTp
Yb9t3mNGUWjv0ZCt7sjDHCE2/FkelzBC97H8oNpsVCrWZBGpkp7yPt7IG98r
/+NFEyPnFvccpBfZSg3GOTD8vdn6X2rUIwmuluzoPzXIikyUbn6ivoFKbh98
yfu+T5CSm1zPQllvYV1Tv05ovjoD+HWWia+Fan9MfabA1VIdrgvF+RegZgim
R9cM8M1g5sRvRHea5wSfM6absdgkI6DFF4dDIBaO2uPTHbBkNeU0YYlX0kjv
pgcAEL9MjI+04Uuu3yIRFSbrtq8Ah8M/cEVzgFihrydYHjL413bs0K0PBlCP
tuR0qIly2AWs69ujgZujR01uuxWfHXZpXT2W+pSnXK7ZXQcv528Vnyns5KlK
7xYzPPMV3XOYLfw5LUcwl9KSmI5k9saJK/GgHnecEHaxYYJPOxkDFQ2tqo/n
5/BwYGkDNY1cIRyrQw5CnBY7yv+skA08sR5K15t1aKvICswAwzgO+Fq5wyNO
rQM8jI+a2pyNCwUu0Rdb9U6Dg+SmgAp0NSvtD27LHKgQ4rbZvmfcpZKTMM56
hEEP5VyIycFjTlA3TaVTaUdD1qKw7V6dU0wl6b4Reva7diBABKKE541Pmxka
RTV9ZrywcUkwysBSQTnm83I0p/oL/Lm9xN1mpawQ15nUNOspONtqeKvhb/Oa
EckIm47chlTjkyGNpn0i7/xHaQnZ7YH6LJIidO3BiQO+NSOj2G97i/sGwFDH
6LxRM3DExSnD190SDCfm85HVg831JCbOk6QUGbuIgJ8qj5PzLBhl53kRgaYM
fqxSqQQoNK1fR7VHD7WpLRmojB0NvopEx2A3zNsJM218ZSX77noMEJfzWhXE
FxOSfBRaMO5LwDNpJ28q8SPsxwtIC4G8hr3nB7dtVR6/RCL9EVWzG0ueCDW7
qpgGQkWQclZD4sfJlrvcgsb6qEOlPegja9yyYqo7YRDZFWADyJ7pgA9iV943
T0kAkf+Y2v722Y5oabsR+bZQyun2ufCeMIOkaCWjuyh6M7E8TS3xLj8GdGC1
SRInKOz723TmSW6zLQMOhaUfbCOYB3rQfPruB5ha73/nKaJD9a+220ausXvU
ih0CyqJq6Rc6cL/7n45FkYE/7GZy6TL7h5IoiHd8MtZPkFMF2itX8S2llRaA
TtE2iffMWwVOeIcppcG5tLqhLo29iv/w+0dtMLXTVAK+sw/MJBVmr1O6tWdt
WUSlR92ell8LAjcbLyHLO39zaS+wviDnzcWthu7zTHKdIN6TQ3hQAqD+YR3z
x3ydNxJku4g305MNtj9qjwZCDa8ZyLZ87duVG68ZYH1rTAL5g48ITvaAKMY5
CG5jQ1TNlURYTDfRhdDU+kU5Te8GzA02E0xVFkvMQqqYn5WyGc/LGj7PoSz+
Dqni7o+yZVDRea9qqTBL6ID8LD/lEt2nfdjdzX+Q4V97aMhcU+hcOSVqd7Yd
z92oR1xWpxNr/aU9qgJze1r1zncUQkHP3inU28dul2Jg3N/+JV+rNABj0fsx
b4wisQ2pRZVpTBO6XRstkk+EHebHF3xirouHM9sWs29+5HBmJHj/CIfCwLKt
Jx+7k3Tw2QvgkK8GaOIY8bTUavsa67ll44J1rhun84VG2//py1tsYDUiG+Jb
Nd+8Sc4Dc0SrhjisFRsqpwmZx8yJgAnvAcUvtEvFK8C+HHAQq7UzOklnC5Yx
0tALGC1hymo7LKPYTEnj/MH2In5bwaNx6gSN4FPekFJXVtZNZjpdei9sQ7SU
gDgk+F8dc+dEnnGRumkXuKaz9rd6O7GmAKozH1XQz2Ia2oak3OCCamjerK/V
74GdHN1Jvj11RM5B5YD7a8LLs2vTl0A4fQDxE1+xbw5mMtGd9gIfTArENrMj
5V17yJohprU6Tsk0icU/Vldv+x7qoUKnc0whd4UlFoL6TDJaRmw9Uydh6AIF
bb/NuowN1csMKyHk0ZXxZudI7TJ7F1neQr2jde6Pey5R6KBPc/2X89O/nOPz
PD/x7/kcQ+1PNctCZOTcUMX5JtpjBHgDyxJx31Vu7KxFtfq08GbCTHjyR2v4
pxPxRV3E3tGA3BDpIVd/ykkWkzPTyRIPfmARoXoRI0+hLBckaLbCHZAF80VH
4iMGLSLOc0s0UCIUEW+r4OZoMzXMG4yUcnr8v2yoguNm7bp2LG8OKbMPD8Cm
900lF00ISypAGp/v76whqM0scM/S69kk35mve39r8NAqrII2TaJHWXZpbo1l
134wcP3b0TF375NY6FiOzzi6hH11YW7l3JMANQI7YBhsmlcHGyFNxCmAtqpa
xiltxpnaI/L2NalJqmqfgiPgOLkWtEgw8ne3QjzJ/2QHQGZQbfOHaU9xUTCT
OW3Gp56qJ/DB6mllJZ742BAGxcsia7BWsILS1jx3sRx+VP24N18AG7/8Kgin
kRQVh58GERjKDhvJJNBpWFFI/0Pl6LLmOLsoT1hr77DWaI8r+3KL/z1Kx53a
xoZ0JG6WXHoo6LS1hvl88EA7JUKNK8sImiEBui0ghYWwbh80idgyAvm14SIw
EAfhXmFkbTrAQm/XlxInqQ1YPSYhX82X9vVpTFTiwN+QW3hIE6d3qWgPqSpM
QetEmrKEHVy3eDMQrUaotxFGfnfwu94e8jCxtke9IuzAPLI4Oy2WQyqghTA/
Uso/TqxeEzta/wn1Jeg//ecchCuTx294+bDltHeAdEbSLh2bVCa+qrsKnhAV
tFoerzFkooyDzvtjc1c+6uMeHaEQxRicc9rcIK5G3fXSrhqKP3vLogvHwDL2
+stSy0/mF37HFYXW+xL16Ud3NNzbE+pHgUdaCwk1rdNTi664Q0mRQIZhIq1k
Z3a6EbizUX0hcDpy4E3LNSzUitk+wkSadXNZrnjXy0JPWk6k/QWlMojmzttP
h5zYLGVtiwlkJSxZ+gzBnA1FCdjv3tDx8RDiAz449LTHlKBheA87g+6fuWym
IlvhpfQYFR03NAzxw0N/vieOSPsmnHMCWxcQbtnETnqeX/FG+9jgvvAbNmHV
Ie7MVmZW2p8QPNXrh3UGAQHqQQpu+aLXFnjY7UvsmLmKxKPaQOCafiVCTKrX
qcZsNxuth8Gmt4Rz3i/2IFRf5q+KX4M00tHPLlF4lNUACAOY3FPuMU1dxg+U
8d/7YDJN+5/ajRPNrOy+uRU9B+btR3ECHzhnDn8cAcXzAywyo5L45xPBXTi7
mw0Ddrkz2BZKdZub65KYziTfcQDr3PcQvv7R9VRDWGjz81i4gXKcL/eDn1O0
bQ1MVVgQ5YDn+qHSjufNn78UmryrBHWM7jeqzdYw28ciwbxbWjkVCpQlSRhd
sW5vIIqQs4YvQ9/6YvKmAwCswRf7sflhb9fSQ2c87coMtsUME5MTk8vMoOJg
dlhwPBUN2i1vdVAfOj60eBxNgDaR7dMoR8Y1gCzB+/zyQLCBP1C781SOoKUI
usekhlcAWZm/i91stv2TA3Mrf/DV/nRTSeYoi2+zwaOmly/WG+OGolcp+VzM
ZsfNDqEoq3wzx3wc7FwkfokxSTLuGP2IN+vrK+UVArMyWmh9z2KAAH/5TUF8
YJxFp5LGJztozlOpYjKuyM2kvAelU9M0kmh22EW81j/q2RA7wdmGzhfwjus4
l227QEWVyLy1IpBHu4NOGG58pDEIFNz3DJzVfrWRkZ226whtsdeIu95MRPq8
dzpzTaAzCI4umNtbeOvNfHY+xwxUTOLo8SIW42NWe+F2g56pOd5NjoghVRf/
epIpBdnmJZrvgseOrrjQ9O7SytWS8v3fEDzySUEMQpKUYQsE9/oD9B6DIHNT
QfxCSNW3bGbmJEf6iQ52vdJykCV+svQXxJh+b8FNjXqJJwQKLuftecgxbmZt
w1ck0nBNThbcvPQw5YCkkhHSVYEDqQHZzz5vD9+qVJRPej5PrrED5u24WLss
06DEKx7Vtuw5BtJQYlpu5wJAhZJEEzIU612Ck1he0R10Hmj7/xTlHYOqtt1Q
WTMaYypu5pZ4bXNbJZptJMzKjgS2AVQ3EsuZjjAV8d0noHzwSyl2tIP2egQ+
R9ZS5ev3dcAhH2isX9h7HwWLy3reEEqkJOP8TTCpuFQfNqZjBhxXpDtbZvdp
Gc64Ew/VJ3HJ9YUX51VBh8ASN6QY6CUAAM2jZv3fiB2lo90seC5rkBnc+2dZ
EdxE+7j7oHqjz3M4HmRYFWjt8T9Qda7zAE8P2JyFPj6QyL8X1lfV3QC8oZc5
ekM8kfv7nUD8LMeG8bT01UxnK2fr5bGeQJSjR3ruY45RYu6errVvcSBmGePL
GTpJY6TlVyM5ibLG6yxUSlbOJUlDDchnS3uOYMKCDuT17N8DkpgpVFAUcF0w
jR3fw8xDGNZCa9Q0pNmHnCQTQ3YBjgbgBGOffJfoIRopDD+8jCr4vFWo3rMM
SolefZtIJXkNSYatKEUFMYvnpUtfUbFNHeqxAGu7ftuC6sT5pCTr5r2rQMNA
EUciiLV1lSWl6KzUhVdc9B97QTwIaVMKPATqaFtChmnh9AE/gjs51HPHvaPm
B1OXq2+2lCrLNG2zddCrRoSGWlS39D2qx+oJpKxtovn+OIil7Q0XbyPg/n3M
BarErTUIIPzfN9/eyakr+1P9nxUn2kajosnflKYCTQHx7i8a3T6Pt4Qo1EIJ
J+eekoZ9gpRRcqnBRCS80fGwttEvCiCRMqCclUvyZzlUplIekl6gaS1kP4Mk
Rp9YeQUA7nCro5Ij93Wekrbw1NDt6lyPks6tWG565KsAGXf7ijjP2h34OT/b
SgO3tHJ1FE/NpUG8ZOK/WcsrveFhyiK2szUHDJ3pDUzF7J7Z8f0Rbwv8xXRY
83qYdcN11rgIeJo6Ckyq6FyNGW4YSUsWzCHrWDEj6odrq5ufFAFwQdsbQqoq
pjj4Ffi5H66pxNWoUZQmq7OvIwhpM31bKp6fK0DFFAOQATcUi7/hD1IjEcfL
StGd5Set5T+sZvDhXBh11ckVghpak4eVjFp/BMy+xdA2qbvCq7cWlQfVe84Z
BjugDX1LjQhycFOz9KbeW7jbrN1V5CYuS/Y3Z5hcZ79KHNL8i39zGPcl7bG9
z5+Srv5zzwbMr4cSmDcKMESUHy7vJBz/vjMxzBijzVZAMphXs1xOVg1EC1Oj
+l7RnysKtYFensg40g0k4kEzCzoA2v0/WxHdR/ZfggHQtabW8ModnYzhOmo9
EHXnhdVnDwSt6RrP+8LNPI0Y+M2MaMDwSCGn+FavEaBPvqi1lwXDmyjQw/uD
fSh08vuA62mIjYrSvbI0TsP9B1mxosc8LBh/JnGEabDAemehNQuKEsrF2h33
3XVVjIcYPF0xINNjrdB46oRdnTv+IB03jvnuGTZJT3NUkkckZPE2amZUXsq8
MKgTtE2bTXplHgX4hBzEaq0hHM46EsLTq33mB302RfOzAM7W/+gyTIwpreCd
QPFlrbqH+EOQBr5Ir3VIwtUoTgp9MpMA/e0jKfApxh8eOGqqUs/lAE7h9Rm0
A3c6p40nAA5tsDoIrSHP9BB7RUkx7QrDGF/K2/Y0cvqPA8WaJi7HHWY+qQ/6
KYjQvt/rN12LaamKBkbWbWJQ6bBU0W4pajgmxY9cLPj5oSkI5JjpUrLjCTQa
ZYoDXsiVsA6nSeBCZm4axa1B02ExdhdTFcYZ9b3w24tGfReoNKY7mWQ7s3Vj
ga8stID51kg2+gw+7Tqqhn/vJgFMWHrqpUD7jFY/+CZMfqWiq29IlvMyFsyA
9ZEh5hiJMLSzYs316463wPRp+272oy9X8aPAjXfZoeRvMxHCWJ4vN/SydE/9
Fv/TV2IPvU5uKw+8sFYQsPq91spFWkJjexrtxDteXI2gTG0QO1LaaIila7+7
D/AT7YxjW64NGhIl8dRvGb5V6RnrcgADYlIOb0cNZu3G34sxta70BpZZogcN
wiv2EUF+A1G2ZSlpQVykwaT8fqIAPwFL9YWAP/r2VWPzSMd4aBDRMUAZp4pz
fnhSCdIU38+to4iD7NnutysCj/DLQgbt6JQ40q7EvZlX8UnquyG2OuqRHgZ+
N26oliHKxYESwbV/EFM7zRxpgcxD68ahIyID+F+cvrMww2uXaB9Y1d+Dilmy
RHcDowJjFUEC/z2JCci7dUwLFIIk+SjR6YCbKpwQl9CUOfLpZqBzqVRKZBnJ
A9MSVQAqbSLUYuSqTOyqeTfmoVnQ7pmI7qQdVqKGi2XZFtN7pmzOfXchN0vH
6H85bI1rdI4aFtn3LVtf+SWEioF/04hV5R0ANVjfzCH6ia6msi9lyF7VzCF9
05XqaSbzl6OIsdxf3vVs+hbLg/CKCn46UQhsm77CxahKVw5/JcmONUyCemfG
uHHFvIWAQ2p2sjnwfI6Dg5UUCnRrHdBOdQW4WsiSAtvrdk7/ioWdSj5fXryC
kAxxxk4H9+z2jBJQ4ko9ymWTzGrbavdd35jrInlZiqZYvR5YTp7o2mH+VrzU
QgbSfy4ifiA4FZl21wQ/P/KKfgfybjyJvhiu6he+i+m7gDhVbs8q4L7iwE4f
Gn44Jh4NYfljj03uSLmxiGEUjsDPn4Vnun5DtbHECzX7ZLeyhgntops74Xwb
gDY5OsF3RnYp9H7hNgUFddZ2MEZhV+DUCFBxymvU2jjS8VThMkW9qZ9QEw94
bSS5BpRCgMvjpNvI+DulPozlPIkcEikbt1px6Oc2J8OHyzdSsmH7AYbL6jHP
xW/h8j99h5WgshXGsgDp39ZnlnbTfugC1jE1yQysWzo8VVo6Btn68OoTimzr
6eCZXWtpun5fxjb16q/SY1THabUHFEuQqawK+WDvHmRBSB2uRmrm1kaX2ifr
MIa5iFu1+FLvaVDDCKot4Oh4OBhRqPeGR2rNzUUXUs374pa2lCQ9GTMsW0WE
Xp0iICX/PL8lC8bojprMhVdjTlrgXApSDFDvS4DdbR36aF+KKEw9BbVG3HOz
vpwzX9iuJ59N/kbDwRft/0mjietK7r1ppSI52mHXNf7kjFDcPeDJPBP2p5up
gizlV96eHJODs+zrjhfwWfGTD7cLCmiD+Jf7nzIgNwW3pQtgay5+KIJ6IEds
V6LQMwEB6UM1isExfqTXofNz9CruYE9iM3tEfZjsR86uzJDyfZBbI95H9HY5
hqJ4lIj2DA9PRf2PHwIdRrOXuIDMf7eyE8JEK1/1rKzFmC/6B47qZPoNnGRC
lhX5n9nX04FACpn7Y87VB2QVxv57wVu51FkS7/q/y5VaovEbhe/cPOEm5dAE
sBZJAd3y76E2m3g3FdK3ySs4Abzb/oNl1zWRGRiyhqqMki7+68tY/Ck5ZTPh
b241yA7jaLbIR4HzHq1+dVWs5BiH9WF6uKNxqj5iIRg176F2PTedttOyevxy
mY2WvnAvWPag9QRvrs7ErpON7kRWeYTdEEy9sNfx2SVW/UozwbOzWCxRak1O
5KXP2Fj8r6vPrwdrvulH2klu/Xdx8Yc6pcmlMOv4OFiRs4HS0FmsMSUm92Ul
Obtnr+G/yV8Gk2R36uMeaxNNgYz4MS5ln+rbGesJ+P08iuFkMl3oZU/l0SfS
ycNd3dA/kpoJoXsq6Tg2ldyxpjtwRSgwXdEx/MqTzv4nxOFRb+uBV/2Hj+f2
hCqv+Kpkivlu6Dxn3wS2uyDkNl0XVEzh7dejm1zHlekTjgYq3AdASzKa6qwB
qalHP5WOJD4bnPo8K3nXcLDTyVS8s+ZtDw2Qr7Nv4LQtKI/gjmzoHanfJSEx
74Ne5VKeeeFt8WlHSGgAyOGVSPX4Lns6lhloj82Iwa56TNZfBY3kx1LOUi7g
P+YBgafHMIDu7ZTuSnOB9eC4q0DSitowMeQxcf15r2iQ9r/K/250hIySdRv/
UbN3+F4wrmjmi23bIgK9LfBLh1pATaoUhEg6SXueJBkrvxeuCpnYazb8i4eW
O8RY5uW1sphW3LRXn3MwzQnB0eq5sVxYySL+m/s0SNQ/oJmcH1Oi/2WR7xtB
5N/cBrJoAVkQxSYolbxMDfzYdsbIb44DcimjOGUHBLR+FZuEOqR3ArId46xj
2SO2/+r6pBObDlt5TNCN9cn+15C3Qu2WI4WHdHUgCn6Oa7hk8TwxEaApPdgb
pT3/WWszitRs8jxgc2D3a7uEONgqZAGL4hIvVe9Bh90i/hLHdnUem81rtJvC
ZVUs1rd8RN9OUjH10VTMiYcbQOYDKzmo0WvfAbOQ2y1fsiKHHQumw1lXBHqd
1Sqf+p8QbiW49NMGpEKEcl9Myzh9CDcPtKaOkkTi9aiM3vTabVIWmfObUzmq
JRn9hmpHsZ7MBaQIVp6yn4Qt6niRiAB5PCy0BY6CMkP9MAn+3j/098u6zVK0
UVECuDr4F5mPxETtRE+gV5WYgJ2ubpaZp/2/91akvVof6/Pcg3H6gzrjO+xl
5ykSjkcImPsoT/wGSoMUdU/XDTNpWajvMeggcCbeL8xXmZqV0NAmICbsFdwk
UFCD8+4BLl5CvbWm+Gd5jomu4VpwH8bfGMy++tyETJhMBwPXdQ0pEundsguN
zqvCShBrOTvpA4SthO3OQSThDp4eKG4FGUp5ONdWza70m9PuXjCjTGjReW5T
Bdo8jny1wGUwZ/7t6UKaC+ijUrL+xsIRA1hQw+OJBzPRRUzaKUqNWjRmaZrT
5Z1s4+6nWiPzbx+A02l4jgOLaaoymi+C96OazFbKOKmZQ79CCpp9JklbY3vy
9u5oSsaO9PXOS/f767UM3vdDBUd5KpannMJl8GZYb/qQykeIcOPRJSNqS6ZZ
qpImPNXoSZFNruSUh8MMGsL+1ddIxVhv0bDZ/8Zk3iNLWnVbHNGqCmFi9AFG
xISVBvCIcmdyeEy+nIxs817c+iJpS9dpm4ZAsao+QV88FVZKnOp9DNuABClG
nbRiitq9oRUopisxsUr7fiBHuxwvli4aMFDh5ySca4YoPiNwkmVQWDThRVY7
HUKrGDFH4CrNnG7Z2okotItKdn3pZwQo3Sx9sKuidG7CRYPWYowhlUh7hUpE
b/L2GI4E/W30weJFaos7hQmpcn60myp5N8iXiFBDIYCcpxd2IKcja88v0lSa
oh8SaJ+vIB34T/Dlx8W2idY+f6XYyMPvVd3BuyVTBjGtSui5MGnKpK3yfpGs
Dv6ruZd+j0pa3rS6OjxHuFDKCffOTIav1iMbvvVAkvH93Dlnu4Uy0e7rDYPb
lI57w8fW3wzGc7cCu+E8HQZTul5m+lGhbPFEV4Xpv61BtGUmd2hJOvM+avUZ
oXts+o/r8NkwZuaJq+aCG2vFuqPZfadb/wmm+f3q44wfYBp3oY9gJBou8Csp
v/MdgeodK8txflz81m6aqkphWm82NNNF+1AyKF5nXeFza8/0ipE/QV9qXRDt
oTHyF6SeuLP9xsMfXMm6Z0Pexr9qcYwsF8LIAgh8KDEXd7RiuojB3dvr8zju
TzawXGeXvQ2cjfNJmMWQYW9UuXeecJoKvrPExueMy1U47ubbArkBzQ/kql5F
xR0i2AXVo9milWBADR82NU2hhsBMCWu8sj+VprJDw6ZmvskqyOaDJhtN6Ctq
pKYbntqWq63EDj7FASpKm5vHtvFxbHQJny2sPwqMqeCXvYjN6ihaC8VsmDTk
EctMQOho71uwO50ugVOviPeWY0meXhI/Cuds2NJOe0e90V3GpeeC5e6O+n2G
uCmCE41FvADhwr7hN4tVQFs7rDLzTNN4984USWKsPjVoLSDkl4apLv72Mk48
/rkt7kHaKXT0qojw4C42f+2gFL8Lr4lwYG1KEtN891nQzvIIhwe2+muW5JDL
UY4CXRis+QdOWHgbvvplNIjDWTqWRyNgKsyutwlEGDkzlNrel0IxXR29kULY
rwiOtbsOFL/k0vUr9oou12rRzHAELITuoKJMDURROnbcntQ+NCmSfKZ+QzrB
NdlAh6sGJgBFf8ELag4gPLf3K5vin1Sdio6YaR75VsXSvz/RIqm3JubhIDMk
2KzpZDQL8sZ80dAJIdp/mAvyLBPa43weUiZSWBzTyo2GMokaDCAsBNmg6PAD
FUWBu1wcNj3WZYSKbIPgRB+7vnneZD2LUjLBC9kCMnnAkUR8Sd60vL/fYMsN
5sCE6sBfEteAQWXgf7MCuTjsZiT09gIVyjjJzBHKCp4eveGTa4+6S+mXUrum
PckkAIa/mGKqshhDxTtbGE6TsQkcATA9k7QjEbAVj7zR087k+OduK6SC3h1V
hHAxWhMIwNw10NVIPacevkUc9HlZ3kGc1x5JhAoSELrBx0W9e8y/mT4QYVXp
zBUACVD3IcZiHuAPPSrOMPTiUqKHaHxz1BS6jIvv4XMd96BPL6exlGUEuVzs
krPCeiI5Q9OqUgtSbw5XJiXAUkn8pWnISou72+7YCL88EeaK1H/hPy87KTaX
UnOgCSY2mzRU2LWJh9AGm8W3rhek5BHAgAMy+ynTG0zQaWeivOqrHlQ7pD/u
LqYv+mwP3P0XHJoP750aAVy+NZ9HUJzTIjwR/12k1tTU3Y+2ArzAyn9zUVyx
4lCmmc9wbW6Tf60tcpRd9FYWx4eUCALgf4smU7iA0Lr4qJqI/5+6bR2aCK0E
xD+fGv5GYHskCopxZlFOoBgzdbaH5BKxoFOqld3SLC0CXDzMXuqJpANpBe+U
VV5HcaoUKWtueYNVmhNkE21mg14VAQqbG19gZJTSpmV6Z5M3h2lQWebAV20G
VAjt/E8wEEJakL5iN2LPcYGBd6Ttmoee4qI6YJLsKioeBhJysrqqacUKEIxo
LEgcWKwEnFav3JZfnSiNfOngc9L56uewG7AUNZzUwAajQWq/byUzmD5witNm
QBhp3GZFou82m27wxDYIAwkhn08Jyd4UU5FqROEVMehj8DIR5TwUu71an88Y
DCnF4if/aGsCRLZ23CNhxOlRH/usyLUltlcWO4o87zDorhXEKIfY/MbbaCXL
Wx8ZkPw+PmoHxI+y360AeTpmvJQ4hfCOhPizMLVz6xmQ3verc4U3KM9tU2y1
5QLrmC4IjuXb9FJpncNjHJpDEfBjs+iGKaGzGKwqqO8J5tSoSlgBWdHTv388
ijo0DDMndwbQN1PEq9tNU4vWAhCH6uNCz4+Qsyb5lY/xTM8Ws/M4dQwZGPOP
f7I9CcOrnchyen0k6634fXG9B3pUMH18kdsvOqPYam/OhJtW2tH/rqTeLFNA
MjjTKSa49GhrO5uKAwhvDHwV66/uYKehZF/86QbTv32j0UQc+VKR00wLTBVu
QydufQSwGCI961eFtnnp60xSmNyb2UwOd3yH62bp9fKH68WXztw3bfIOhICF
7lP/rIbdgebpVgOp+FOvWRSSZE3Jb+LXIIkN+gwjMongB50trMponitdViN9
KDHcrP0Z8L7B6j3xjSkbvKetTABj8thqj8iRWMZTyg488GbLP0WJiHVaa82r
hAE6iEMGd4EisaSgwVi4L3RgmO2wcskMZBjm83EnsFU6ywaTiZP5xuLC2q0C
HFBDa5HotFqtB8SxY6nrm6pPXvzD841MSvhKGamZuSGpCS9rA5viUAzNpb8c
pT3NJdjyfi1vQV2jw5GRQfD+r7BoZyNZLQHcBJz6kh7hNgtTPDwO3hZ2gMdN
NUVZMHactOl4dgxwkpOwrQdWHDJNaCDMxG+gZP8458HEHUjAnDE4/Z4iXFkd
9uOKArg2ka3E8jN5ds+KFagGQkdL1O66rQxUg5zbwH0q83bG10k2ApgCnAgc
tG7yOuZUMeYd3QmQRfEoz+kUfTqXmMiDttyuCvmTovLyKbEqb04CCWTmAi5A
kRGSMcBI1CQyQTZhtNoD28784fJY8J9xEwnl17o8YgVoqZMG3sPXwGzTDRQQ
nHNIXTpMt23CHPOM0iqQuWE/6MHR9NH+UZZkUy34+Hx5KPcBcgs6yCmZVH8E
v6REgsreZ5qvlXxawobCp78bJx8hlpeXZCEhzCFMKi+2YA0l5pGnVKUe2O94
QOp7eFVq+bW9XtSCzYHHTP3vq4sCX7q0yH/i0outQ7k/8ali9edALdeW/psr
4cusXT2FnCh1LUynupN8CH8c3g+yIeo2VRpfIfROX7Oo30t1V1+9mAsDMYvU
faOcsQE43mRv7SRS4FhplUwpCCJRjupGKeX7Z7b7GDSaezBNK6OPOsudzqk5
UEp0cdzA+e5kFF8a+q+0BgLrkANzmMj4yL+tGH/ecaByZ+mH7VuyCuFgG2V5
/yiWI6+7UVvDOKO0If7a9Nm43gOIK+CFPPOqGe5+6AiUeS5CKiCHiUXDGg/b
we0t59MQRgNSaP9YENsGbX50myQu6Bm93SAmjQmowCpvOPT29X6s8NKKFcW3
IAjAbMmnVz6KMQp/e52v+PuqopEL6qjEyPYUFMJ9pVOCnyuy4mcY8Czh7tAO
QTEO+xEbJaWpVgyJZXaVolt2zPB1nyvrkjArt/rfmxKUVogHx3Ebrt6bS5Qu
cAEdEwvyQ+u2xU5Pca9WenNmIQk2MQSEZVrOay8IxCe12EgRRJnV44pJb7PZ
LPp13hHMFgAP1+TvS9ysuDxJMxKJeuhx1vvZMwJNzgsiBHZAacAlvV9i2fYP
W65aTZ6BZtagreNvBYWeM3ChTY0gfwuqd+q1t1jF2NURJv7H02v6Oa8Mg1sd
7qJQ+2oBLDhOR9Ux+V86xHUvKsHKHbjV+qID7RM1yiR2NER7Uzq7WHtkSl4/
AEnvVuO/lgx1UT5QvbZXnusZ4IL5gQzqVCmtQ5Al1zEqqMRcYvhrXvxijFj0
viOPF/1TPZL6l33D9tem5tqRGxbzQCXYXqloMbhA53d5SeWkrBZKVrcDlBwi
41ehsCIluP2KaeVitvpjS/zlFNTex+y8SJHKbVf/mIil9AJHFXv8xF+MeFTv
aiRflo/IqWKlTzEIf72jnAGb6aOqS0fNGXrJUS52FtYmy8SDf3cKhwQnezFB
s7nLPQ58XtLU/X9VOg0ENy+xhMfARstQvQn9gu582VwSfSGotTv4NA6P6UBr
Vf9xxiF0NZfmCZVUINnVyIOgsYuz5DVGDRgOxISXcMdYwhXPmlTNg5r9gQKG
eRYnInK7AgIXK4WbXlVKXTL/jEf337ZNn6BPFeNoGiz2DJ1Jx/9XXwiomKK1
kEtLZLs1+/h4fmWr2RCvEFc1m44jpvMphhovKGOijYqhw9Ps7GS8YeAmACPs
z4t3+wqRD5WjZ3oBx7tFXxFvJMAxI/6PRKo+H+EkEFVy6Soi+Ia7tClujjow
lUx7BPadWVl7q1u6agJ61lPCYz4xqgrhlBCdtptWVsdThrfcRzTvWMCdZ3nE
U7Gowa298DS/vpwvh5FarTNxq3ynGShLcRBNaYCD6HnYDRoCGKFPao2PK8lO
ZL3PQuo0eeOn8k8zmnguSidL4H7/NEyNC1TyHhfti+4nVaJo4vxFiRIEo0uQ
KVVfCaFfzyZZXLT4DOyg/U07w2EGeW9bUAUJqn/1mAStUEuUOarbBf+rbK9x
NMPbHEfQba7g9akzoc4+wDffQrAXvPFw/49MsDg06KzLrsmN1SVjTKrhopZ4
8NWNCURRbZ9qf9ZdQMnnXCYG9zOvsJFavTxnpeR49aeLMjsmIBppBRy189Pe

`pragma protect end_protected
