`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
NQFnKZSngLUKcY46LbhCyIkmlwTME8HPzFEtdOtWdIyMEygAvztMIgooDlmNBGLE
bY/UH7oYuUa7yEx3YtfxXwly3sK9KIoSBH46Eanfd9pfDske3p+ilTCJrcjStWxI
11pz6s0AKzcgYv2OOQCt9HIrf9azMV35z/HAijPOfJY=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 11360), data_block
oG8h55XhsTjAgbJiypbXT7TkG5WoTYn5qrMgjtEpmha4qWWg90q9Bhvnhw11jBL9
qyO//UmmRIF3p2T1pHD08OYWdr9NVB/XNjVFCm8Sh75eWM3KRs/4Dvez8QNoIJgv
5ZUYObdzUhRA8LrnrOXWlj7zWwW+H9XDNWz6R8fs8TnhluEIDs3iXP3nfPtLOtOa
SnsRV04p2DBrybkHxqYPcTP8iOCKB8IjoyX0piLadQoZB9qlnzyjUXKZDzrtp63u
sFonVddcbOqRuu14zw0SAU/b1MaaKjV6dD1nbjuvfPB4NJq5KXQqSix8TFY2W+p0
SwWNjgmBkg1U+cTI+5rRW/Gw6iCDJ+rOKk4TsT1lLbbJJTu2rDCDn4Vdkti2aAkb
HGTpPGLPM+ZoNbFcQBeJIXNY0PIPtkjI4JgDzVwA8FFpU1fFJZe412hH3t3s08j0
RK+LGK/RLFw/ly6x804ragZyPbaUwmSdY97A/VTtYExmULTo7Ljr93cnAeN/Q/uz
HV1FVlAhLYNJ8DpyzC776+dlutx0ay57hoXmL18JwjNe91YLppPHW1t3cqx7oMsm
cTCeuClVRz7Hsw59CpOY8gEQfY2T7j8I9DKeY4Bncd1ABG3QqiXCkrqTlKeCpLPb
0A8r1SgOsVQBHnHXYxyOVdMcozzlXGStDMh5n/DjxT6Kg8KjT4uYHDodIs5hpSwa
VVuTiPXbbK3kJhxHnusKt6d8KlKkxQZdxUFsz5/SOgMGj86BP32e0uQctkLUtQXa
3hKSjtYGXpvH7PNZACL0MslJ5aVPVRPrO+uHKdhEtzOZF7QIem9j/CjURH5CPmLB
NRaaQnRHMX0csLEyLw/lhtk6Ud6gtmHnCoIjQMd4+MlNiV2kPGZhzWnyMzDUS8Q/
Mq99elMX9GpfPRnGXSZpLfquWXTHMMsVwB5F5rsyPCwCYQuodKmh4p+muMjbQeQm
aefYTtEen3sNhuVFFgAGeaF2t3GrHwYBe5hGGGIhGbmJsMrrfXfNWQkUKVrXfeIL
DYg5kpRxiQCcFCW+cGXL1SbevvlG7/YrEtPcZveRVpu3f3ogUNo/p3Jp1zkYE+pW
SZcBT6F1tJ3xSxsE5dJVzE8C2hIoT0L4gUZGHrMc0d+WPhBJD8bntN54L0AkwTV1
CBvwJCyIN1IO+97tKZ+h2BHOdlpd1HYve7WN9Ff9AEGZCHuTic3YBmoEZd29vC1t
SdgZFmuvUR/8I/NE5nCjAOYsrIBKLXh/eU37nKAqUJQ/Cs8106+j9zMiJaI7LBhf
AnZDVhTzZvOAbVbJjKLCHfPQyySpu+zSdlpbLUM9XNkZ0Xu2QV0K0wkWfrlMBdQm
n8VVRhLp4oPAuaMar1rkK9BqHO1weOt8VNc/LLAvvsuW+U6/QMTxq4Om/9WOSVh7
db7m4ElwZ55Qq3tDb9y8RxP4dGx/0fjyKbpsL1ztz/pFk3KHZaraBIEx3K8Vdt2E
btgyobaRyJjKEFzGVYmnaHxtlUTCEurbM/cQJGouj93gpU52nLqsjs6d6/ee4Efd
/1QuswnUIJpDcTA/nnsPSegZ/TeH4BiDWznl07Lg4KrsvJ/RkUCWB5BMIlE/NuZZ
R128+dTG6cY6+YWlV+VN+WPBYTaLadKbXIk2ccp/NE/32NuoWpWpkE3FAsdk4bU+
1tJfMmr7MrAGZgevdqUzo/CNsqEZM6xQEw45OLLdqdk48yMcUfKvJd95HKzkPuEv
6nxmD1oauhWb8Vge6eazKhvJfvF2RQdrN9YfKGRUAOXtGF0a2+lFHl9BVRxLxynI
3UyYK2LOG3m23wEK/r9QmFWuH6kKxDqZtBEO8xh7mkFxOMOApauD76DdIa1SnOBX
OGiaiqexnjWXktk3GjD58DnY0N6nwYLYf6v1uneQ5s/8nGPiV/PmwS209Sx9EUbf
lHE79znG/bIIVV2TmbjP7usEWX0AQcWLITgHKNYPwrQFrzLyqq4Jm3isVvvFbHsN
VerhV5nbNwWf9nybtVAYsD+jZ+ua3kOoCJmgDSjx/4g1s+tmE1EPyPk9DPaGGp5I
prrg1tplO+YgySC/Pu0HBtYpLJpJhbfj82kehYzXCEHqHahKlu0YGgYjATQ/87uL
QZQyjmddAHrisSBjKDzm/YFZAayefX1HTyppXncRJO9sdgtv0i9JA/MMFG7slet4
nPlwGHfeXq1UxY61Jt6eKTGTYWjiorgo/oeVVFjwcGHPC6l5aThwSmQ2sif4MYK3
dqlxDQsFjnoowwJIxlFN55OpSCG+3W0631PbBt51kz93SviapDzC5mowGpBtDiT8
ISzTTIgem2ExPFBaAMt6fkt7FD22E4XGM/x/0hykMEipTmyFY8/Ww0+owXFFy7Xk
toGm2jog9nrJ2hHojZIzKDm/1jdTm1esaaHE9ulkObfYD4AJqdrqTezezdcfK//v
D3VD/wIq9Wv2PJcOEy7RRkIpGShnvsQuzJvqNUS2kOVC8FK89dymOJnkvJzCAj9x
AcyB0e4YOGd49p67p9IrsJFHMvSZKl28HDSgAbxGfl9DpgCNEp/P16vgQ41g9b03
vS+AF+R5BCDFPHyalYt0tHA+QYOi2M4Y5tXjtIRtNDUKd3dUxMXumZ6w9XwyKfK1
hunB3nhM1M+oHTxoXXXFqvmwwLR71OpT1IgY9phyMljaHaqe8xNcCzY/q4Z2jHJN
JO6Hu37hhIk13LpWKnJzmudaYX1YpuvZkSwbevKreJNbSzTc4L2NTympXsbyaA/R
qhYURgjaHbRmfbJvrboM0mLj+ibLH1vnq1P4miALye98z8oX4gmZAIj+dV110MTX
HIPHCuE6WXjGj7TyBvkS0G7TO5r2aLbOIne0BwglzWNw6b8z3eZ1J7drqdxpTbzl
hjaqiSYCaBmt7ZnvkEL7WjCAnd56NeepOOEfuyM4p81TMsO0eHI4M+yz7jcdOtnu
7QKaMyB7uGhGIOE+JFFtB0YPZ1UiPCSE332RrNnWA9Adg7YxG6yoQRrPS8P76i7U
Fu/zdg8OL1lY4AxSPRMbGx+QN0D6lHxdeWbUYrXezDSgFszYzgBG800HVVfifH1H
Hn4rTM1LwtWxdteMH8FrL94o6ooSPXU3PrReScNbTFSfGq8ucXMXp44yAuFMZZMK
B5gFFoxKn3+cmlhvofZhEBHV69/X/NKYkN5G/Nt+7N8GtVHqhr9KyucOyIReY+jx
gus77pMKilexwwio/T4fjqajbCKWP0jebgVNMMkY2KeOws7vGwu1Vu9rRnU7CCqo
b6mcFov4Aa58Eb/6Xaoi9mdWnBcyqHnV/DfiFaz1pm/3vwWQ6FWZSFJw6xw2LCOa
WqOHPF23Pc1RAeySFXzmOpZLLAtVEiRvD4w2lCk1gyMBasuLePdR50B8rym+hF4O
bvaRZ7k5gQJWNWDf+sWO1ghNLYZnl5K9rfegd1x2sYsEY4C3uMx24AGvPPHGX/8U
WGh5VB3ASvClvqxPhA2yB7+Q0anWHBXzcoL2FjMNvhkwzpMncwXAqOq95qP20sAd
sr/SfdnMxBk79CbvlD5VckmcPoflcCC2/Fvh6vzRU+/nsL+BEaMLUq/mQeaeTeam
Do0vISMylP3jUkaN+8UKg3UC7qhD1BeF9+JwTBb2bOVbUDiJrB7YHNzBMe+1wERY
i+lfr0SAhmD9zGnTNNJwQLArR60Tx9wilhk29UNRUMhgbVb0Lrn+f4DtzD8SSAG7
a8rzs2Ab8yHGb/8pxxM9RSF7tgt1OkC3L67cvacRgbQ37+ZyDcrXSY45o5usDVXG
qvX/G7BLKBYNWQs+xu09w193kpKSZYlDoRyH1M1311SqT0Nn52CQxAIEWECA8fVA
nmAY9kWPobaaLY2AIWCeheCW5H+4xF/s8ISQfh+6NqgfFqSZbwR0uUmafgF1BJb7
PmmNxzePe7SFgX0l9w/IaEq3hj49TZAl3ZYJv3/Nd8qXTxUrmpvE4uBdj7kGWqfe
ILEvnDTi4X1shld4KsmJmleKDfn6HesHvHPXuSFD/Pr0xTWoD5z6Ab8r4ax/af8O
fbMbCNV2pBxCPujBvfL/uPv2OMcTZ4h0k5HXEPEaW8M3A81eE9+kXo5Wio0sh8KH
rnR9C3vlQo6N/RwSdJHWNBepCIbQOMw+S6fH/c1LNpUiacSEBG8509cIE3rI38/c
v05vdEZmDo+OrfNy6KvmtDz8kAAzLUDqxUO261sAKLhZvLgh2Q/lyu49KaZ0tyyF
y4Im4hMNaJx+CFS6umfUJNbkhQvU4x3PpJogiDrFCYmToVY87r1l6tmmB2Y3zCWn
vRFzhgWwAStMv4xqL11LIVT/CRXUBJL+N0o3jUIt7LHpzcboUJ4u5xWt4DCDAdr7
WgI570qmq1rzpxsdixV3w/b+HXjYKoy6WHRalriX18ZiNJv2NIWXl6+oXfZprPtF
JNCG8Qmed6xd7pc7+n9PnARJAym+9g2OcyaR6bwcsDK+JBKyPFEUvyaLV64WVReA
VUmBKRxJiSzr/HBv5D3D8a9Ny7rODyWbLy26GshN0VSA4f8aOvbUVvlW+ArVRZc4
nKDg3HjqQcbqsBGLQOu1J8tkMcxHAXhKzEOqp1ac4c8/VyPYCSEl6ZGd+p9ItZ8w
prnxXIidFx9NbdStfrfKf2O2pQsVFHligOkD4Fa6m3Abn7QXazF1IfM0xPljWxWd
rcj3ycJ8IpsAUgAUj/IVnqdPsfX7j502xMCweZt6lQcBgzxadD0IXHL0qrJ7RiV9
cGnR4012olQ2OshPJWaJ2oti+VkFsff2hDLd5gT8FsH5hcrNtfhV3ayGLXSj9ILI
9Dkn2oi4ynsrmno+UIJcuwvBTFct/XgswIW/iTushMYiO2IMYftwVFGOeCOXxjhJ
dmHYjikHoeatBFa/nrVGu6H2O419NJ8j8Ed1sg+PZNDQYkO0wlNytY5nAm84M3w3
FVXSXSesZqyITknW5N+Zm1hIeODbNAl7lH7ihZGYFFeUCTX3T4lUvEBbHY/Q91EK
Ww3hV4yobXtdQp2kKeku3dugJRtHPKvugflCMfpKcyFoymBJ65P31uO5lSW6YstI
F6br2ovF7diX3Vqs0M8XVVjld2NhpTYwYjeADldUfv17zZPtG2M6x9NYDkGxop9F
RqfOMoVPUl2nBdG5hgstoqKBp67gWGVgVbLDI8Y2Fk5U//qrwpFStpQ34EiUxQ44
369HARSpoYpcDFt3aQu/X4ys6N0schgKrZDM1cQLe58dkgzTUm9bjym5x+boi/FE
hNdhF0Afk9YQOHP08K+IzOWKg+WPKdex+57DqFfypaGJssyjJGFN5LRrN1+sl3Dv
2bQC+TDAhJNeEIYJRRTr+421Q4WJiL8zSpsMRsTeMtcSnp1zBNflYr1Erxb3M8n9
aWV88ROtseaxc618OJq3f6S/817I1n61htFobg8tXjzNQfhByGOARvR6nZqf7Z8y
NeeYHEq1AhqhtPt9ze6A11oWpGv0K+pc7sGCpP8MCxg40+5TXhhpz2Rw3/INO9Wu
X7XHzeOZswTsHqKQjozHEft/ZiEonKMz3/xwtdIoa75sDDYvM0bNlM7qRm3Iv0/S
POkFFbanCC1rj+BpmaiXgcLl8L6FQj4Bbp7TXBDdPacL4XB0Oye5D9klbQcP/qik
1pFZFEa5rqo4ADGSYHDMkQ1pCjbUrrlVJS9g45RBAQqEATp9+KESlESoZZL/G/+p
g/9Y9lskYuvm33DNoOqkgnwnMGiyncv2s2K2fdw8LopQihvb5jre8XxzFkkVi3Ly
rksIzYEE5iDFHJgF8bCFXMW+3Kp2i9/g837pQbvji3D8F72Rwo0ktTudaEzLjTuH
WikV+iWf7CxWcINzV5jprZDhFlS5LG0Bkq0v3e7BmHuRI1EUU2G53ak2LnDZ5mZ3
nunoPiLDDlh89IkokSrukdTHCerEsTZBS3ysCz0ZwVdZvIqJIhbQbgVYKURuJL2M
lbap5t4CISbMrGzzvk3nER2XCiqyi6lwWT2cG2JUoCU6endttxdRdkREAn3Flq7V
KOLLpuAJH6vG/RVLaTJ/5m+ZCVBV2n0FIkUL79DTNOl0Ds3hSmnvjlMgVPXnDOAP
9r04yFybk8GKfAqLqunVm/h6aJMn9pq2SoiC/wbogdr/aG4Obx8gDWOP5LGFUqsH
Jk/bWXr7bGiT6pHhh+beV+Y4NfjXszPqg75OWUSoOqphGluEc7SCRjYY7bjCeuNE
S2RerM/nDC3gwJDHBJXyoPoxBpT0u0SGJ3g5kmRegONvOilddomlV1tgPTc0Xm5G
MxbkdYxl416YoqsS0KhebHgZacmx+jCb5x2dueKpqpH0y0riIP+jSKyL5kBI7lQ1
Afo7OpT6M4v5KK0Nb4wzp+OzMcZnYHmYB3IQa3DwG/pozqd6L/X5X8mIpXM3Dw0C
lZ7v7RlA7QLcSmRePsjYbPsnU+QFm/ofxaqeVF5X1O0Ao+GKBcxacFBYW15ym6XI
kOPYvQ8bB9Qzdee/1Ni3R0eIEfM0FYuo0bzaUuCG+IQAm3q0yVW2wIv3jGJb17rV
5THSc+cq2esScTOhzTmh/eRzUbGxawz+90SH6GBMQtVMjhOv9rAkwLWtl5+ozDTL
nGX7Nni91CQu0t8JMo7IHu38oQzMhkt8b/QaoRA1OkwlGfASb3AhxsdeSuzOr5xC
PEsB9EH3H3I319y9yTbwE6o0zqq2whqL7cIw0fsg9lY21phg84HGamcvZU95/ADh
1I2syHCbKTHjnFVgykA0Du44TIgILihWtfdQS2cQMbXmjBovrcozHGbHaJzBzfGV
OLufYoJzm1/1Agysa3pWdhGYsvLxr1T2LzgABX0y3QxcbhvT0EWDszM9uhIDm/Sn
9kG3imkreBAZTPHMPJMvLBXS1v82g+WdiKrK1mQLhpcBgvNx10gcjoZApTAfPE9c
iuEqIn5QSF0YnJgqNwgrem+kiIr9CPuKVeBuy9/NqP3bHIVUMRO3Pb0XIFFi9szM
6zbbT0VelucNhAUXezF1vN/0KNRXVJ+CXSEO/cMAhNoCwcMBUo/ac8/k2jFmxAWv
dY2z5KBGr200hxPd+bCvJ8YwzHH9heNd6anJ3aOL+FGBhocLqW9RFYfV8y+rl0Tw
CGIlr6LYvEKE9WCoYnS5aJ8Pxfj2oc/V6XUIxENlkA3ic4yA3/WAAsax5EAMRmYA
41uEk0iXhA0bqJVlRXG89AQGnQB5ewNNzsjGfVpeNrWMJxX5U6+rpNke4BiZzBdr
Kf6+D1FZN2bJ+GMUYd/B/gjfFvomiOSxWlQxoaKxYMDYBJUySTyCSVyrUMXFDXt4
3pm4KELB3ST6ZuY3h271NoyEwSJq6jHQhs9BGAvnhr0DCPa6yrAtT/1L/cb8bPaY
VP0mndP3C/f1y5idiioHldPF4q1H8k4WMX1V+a87RS9l7+5VhRJgUoD+WHuEhcd8
7zqhy524UxIF+Juine4ISA8S31UTXvnWWwQnCY1EX+LRDbGdjkJhqXYmzK82TKBq
FIB/E+wO359NdUUajceSpWUjWqkzMANPEpzU8ob5cH8nB/hc34gZt4qvu++r8PDV
zNaXj2+/35vG6yXn2mtYz2Vv5kWmT0lnAQAIZijW1BK91AIF1e4z3ODxHvKl8QFg
UHch1We+Gn74UAaUVQI+Vqa88FMUDSBVqtz2MBCnpYgfZuZYT5w4Cpl6jfwaDcCA
ZaNef1ZlaWp534d6Eu3FuPQeyhjsXg+pEH8Bgq7mnBZnZ5z5X4wiRZvMPio8q7Ul
CJu2dY2vpd3ucRQHSFE6PiaouoEnu2AGRiRF8BlCFtnKilDj9orEoXAXPEkzVvYN
EZ+41GWjKez4GMFz0NJps8e7tzT35mRTAwa5gY9ap2llTElyQX4iUoVuYPsjhqFM
UPoaGewia7eGZi4D4gGOg8e19AwuOb3ga7GW4UWLctsw6ukGNFzUwV2dYo8y3rSc
UjEF9UlvjFuW32vQTu9KaVLvkJpZSXSIvC3WzweSS0PMGGTrz5BlytjEeF7F7S0E
Z6rFMX/fhD78x+f/pKJHssTQAH3vVTXGDbXOClbd0AmYMI5tz6oYFSgObsTEVVhs
BrbAlg0PxMX+xUGzU91/dHowZvc9pnbsSWnaYdvUMxQyZQUFUX00llD41swEppQh
16qZbMkTjoQfQNAwwWRFSehVNy5auX/6Mw6WNVS9L69ykDebHKSfdCnprd4m95b9
AXPXMC0L8avfYY/YT8Za/tnwkirzrroYI7hUjdkuSQK5rFSd+Bn3OlwGZA0NVzfB
JHQDTw9JXUsb+gLLyrZTOTTG7n5JPijUnpkCgy+VOgio2I/y725hhdvXOclK/qOk
xMP4q0lh5VeDV3SCA9+LCEDCrqXR9oYEnxwR828uIxgU+DRqJ0uI67Ei3gV+o5+r
cSEZ8YNC3lwWK9c1SYvsMskHu3qER8IfV+CRi8BNbTS7ac7elGxqItLbU7ZxSOxW
m88fSGZCE0PdNAxhst/daw1BQMIww4GfFh7qsrywCS/YWztZWa3laGyWMci5K1CM
9ckuqjU7h8lPYjqbWORAycMU/9Rv2geERBmaFzJmNLhRpwFaM5uypIJlkrwBGWGO
vDmEd6JL4DgTe+QpaS8yKx06k0KSI9W37JchLTpDt1lQMediFOjnXuqoaOyx9Dc3
LI8UwZ9gKLZ033EYwNQb1oNCcEuH/cOW3nj+srOC/uf25g8ZyIdCug9w8Md+8anX
BhH2lfDFnlrOFYasAcvsMNXxy5SSTE0mQWKztsNY9Ewi3bCT4vqjgz4F9mMFYOk6
R4ek7+sxM5vmCGhK2OLEHGpSwZS5gZ1lYaY5bfY0bhpMVeFfTUtipYnbEMyG7Bes
afg3o4zIIQ0aXOOuNOUlVBNxYISMnRKYXtdieki++aBgS4NSZUxmzPbiTHlRhKKX
nK0ScijjiS9D376qEkbMSshm58O7eOjIbabpzb6miNQZdyXdIpOIJTfpaCy0VGtO
+h9exjlvMJohaxnakMGHa8puwnH1xZGjaZO3sKs9JBvR8s6ufJ7mZjRxflTtihn1
4FpZT2uL9SgKBS3JlhCn4b3F/cJe30fIUwhe0uPUSpNIStV1SQ3CTBSdG8ozWrOK
eA62wJP+PtvIBE1+TBQPBsDNm74spZCCdl3n4nkH8m2cSz2d+1dbFExECSWNLeqM
8RdEx+IvmDwq05oAqaYyeUFuZkyAf8e8WeHgrhyngGujbIcG5uRiPhFlMw05aGVL
vejfp6dV+0Yh/PKiJJbsYybWZDoDrvsY8/b8ppGH9JSTZuex08LisU674Acb9Ux+
J9Hbxp2oebv0tSSyMqPP9jRS5z451+knFXWAK9AkZR8NeoW6vnGdwsPRZHcfIhTD
iIXUpQ/umC41+63KZB3c+H9hQZfpyQF+5UIxyRnrfH46pk1J0UVfgZ7lAe19KcOo
4D3RzhpL/BuripJ0nxD5IRA5w9Y+zaL+p81gqxtc0e68211oLHVaV/yScEsUsvzy
7vhEstfkWlkJ0evuCSpTm9FOJJrUkCkiBbbQ9ab/c5k2uMeZcinKK59XF2/t1xO5
7QElA6uQnNPUpR9JVuw0T9Gy9SGgCO91OH8jqpZtiAThkIa+5omjAI1hjpOrwUnU
DHtlez49mQv36VHaZWowAiNRzafmEfZJZAE4YRyTJ5B79aV99CLOo5bzsXRNp2Mq
FDE9gaZQLzgsQAe+DHKtGFK7ZQIYgdYiFJ4fQ8VDN/pLgdF3TiweN4NoAJjlM3DI
WS599qLsroTYvalzijDbLlgPcPIFOiquefW/coxMPmI7Cq2+06uPwsP2lgpVK4rS
+y98LQPog5MB+021G7Ey7qZyIKL+KYLRGRERXwIBxRi2ctIS5GRmtKpOciKW+Cr9
3Ugn07vMlzyLYM8YLtxnl18R3KxrbATaiw5P3l/HyBmHOfYhKn9tb8w4Qq4nHadE
5nGffHUO+F7vQhj02Er56PzG0MXo9mNQxxtiaNtwQ1xS8xU9TAUfNlEXCdhfim6p
PYbgFGCTGRp7AsgtYY6vjl9qa481WXMohOaMNCJ7ZUL+w1J4TxS2Y9YJ99c0AaG2
UKfn4QnktGi09urJnH5LRLGwkruBzV0DdAg/hGYg/+VzOGI045+B7DCsfBlYcg25
F7tP98K8pwf1MgvJ8B/YyGPVCaQXyDziB1Zp2cEThrEAxEINYyDdU6W1GzS2YPSP
2Yi8ZhZt7/6OBc+FGrLbrRYRjV8GrS/48U+rACoTkrCLZH8CPd6HzjMHldhEZiLS
mCSgXd0CzKcGJq52mHJOst9g69zDZR+WmqJ4aJt1CggMABMvGl2wMdGGwYDZIsxe
JXXf1gmqGTUtGB1afBOr2Hny6A0S570PLJLAxDRmY5UKaHT557vErmX10DxZlJSe
cFOkW2F2GMD4V4DrkG7fn1dZ3wEwjoNjS0lc5HWSbtboA8nErvTExME032cYU2gO
/6bE/QqpyXdUchiMtafWE+jCYZmiTmaDTDeUfmjPjivRBM9IUHqLBkWnojtBROEV
/HsqkcLyOrPYi5Vn1+7F9lH5G+K8I7YSnBf49u5deyj9UzusCGx52uiuB5eGC0mH
FWpX8KX8yZdbcRwPKs3G/X9+1fGDoMASWsiic8XnNZ5WCr5D9smLVDyk0PuVIH4b
uu1VBTvICHAJZ/AfajKb4dqiz7iHs5EPHHl76mMas0VSkYHfOr1pCoa/TI+PDWRj
gWmyJkUvEfneh1DYaJcwYQB5B3jOlSbu93lgqA2ZFIo3YnMKg99Cv+3poXi1g88u
X/jaoOWxjHb/ezgJaHlyxH2MvCSBBXaH3UKYul6o8cZp+3nxbE0S+ebXzczqBIl1
29hpqcAOvu6gh+rw9Hb0o8I/4phDO4FTyRXc0lY79U85TgveP/dIIMd1cMGeOOyS
EDmO7hMnu4zsNYv8MP4L3hSEc+QmBg8sNHAp5bmmsU4QfGtFCnxWBeV6oASg9VvI
eqSJVITJTHRyEvVA17D5thA74l7JFfVuPYI/7rUZHD8ZIZqkQZNT6uNwFAMbiTFO
jwFX4GUJ1o/5qM+i40sMYNC2CS1mjFoUkwOMP5gky6S2DxO6zq8hgjGKdjd9DVZM
mVRNn2+1l4iFPC0JBgodNaCF/viYMD/NQ6RGWLoNHDFC0124MF99/Omi8EVlOI12
rr338svktOw/aacIoCvMjtUvl52IpgF+6nosC2Hnq5c2FTCXSwMf2YiMZ+zSAd+h
TJECBfFeHefx7JROi76obTAzfnsvlrrAkPhYIG3nTxkcTOHL0nO60cDjEkP8NSfy
hZHueFdMP4LaIzv3oUa1HXZEL4T7kpGQeZ9oUAvcIfpcp5QrVbMQtmX6GzxkBKka
ahEIt6H2ErJCn3/P+pzhd6Gpli8j+ZdSJR4GiTR39QnO8BddMpUtuTvkAifhPnAM
EQneqFDcSIIbV12s13p8cd5Bn6j0DVpsiTZQObVPc/AEDF7bh8HZeJYcL8k2fnA5
yUJge0hqA+vCRcRKIJwDRN6L8ndz3njNOuc3PZJzWZwQQT7DcbfvyGaKo3ZohxMP
/uf1pL4kVDrNNiOu0LAkD/hxQPv5ooATk6IiNtUqjvQ9lh0r5N2TP7TEL22hGwfb
vkFjnlayySK9fsz+Mf3nJfq1quvGbh7+kSmpNHBaMtbXfWS5yL6grEn69oFcyVbl
Mke9pbHGKXukwOdbNHsX+9/93PFmOnInUBJmXmyMSTFGVbDbOOItJ38Fkyb02of5
i4XZ42Gw+f79n/NEh1EEjfrZt3igBJFhAUYjVwGWqk8xUkPVdUmisn9bxnI4PQXm
aK20CLmED3KD8/Jf4sdxSsYthjUSe2hrLZjNwaECem9aTG2NNMi4Jm8wMjvZ7M4g
SZmK4cUp9omiYK1GMvhUNocaZFtr2ZuA1boXXn3s2VaR+qq9FQJqnzNXzPTxl8qk
Ho1lH4HulOdJOrvwuzZg32wbzgHbiaCY0zaQ6lRclrwk+oq2hrvsYOycUrAo5S0l
ddMWjggYKwhjZvpuo2vhJcf4kO8QQqh/AY+FRA3l8hImE92q27IdSEeo5PAXAIik
gXXtKjufFOhEjjj3kJfoBARHMP9WJOOkTUUayR3P2d2ybXuMzxkbM/h7wr+K35dm
IUmUXEGpCq6IrpyjPoev6RO2WW6Jy7/LcyrjjWV5hQODRJDzvOg0Pwke4xLcgibs
cWJL2TqpaI14PnDWDDVZH0GyztUG6sOwtKe3rg4cL5Gn4BTr7GjMlbHrjEsS+mAj
g4oaOrI3S/dBF09gXWiGSFkhgLI/885JIN0Nk7gfH4sUj28mJphu8qSKZLLD0IXr
p2F2VHvi/KQKlgk90e9B9hQUctNYloZoijgcY8oO32nh37+gfUOo+fU7Opd8/rlc
Z97hINMdvaBd0CFp8SXO685e/264u2yHWHO7KMBYaoaciA0PYAN7u6sw2WH+fP/C
CWxGkChQr1GZFPbah7WZoeumZyxqiYoMLoVqBN2RG6mdNVHUHeKMaBxFEu8tnQN+
SZs+7N8z2+6Q4HcuwETTbHElgjKmeqIvpM+0JsOMPw4+1ljxDeuEeZIe/Zid8BS+
VFBtHprSrBy+tsSwod2C9ZIspDqZmSmuNJt6s6aIYdQxgNchh9IRBSMT6IbgmUiy
XWRGBdXyRuHL30LWyJYPJJ+HlzXyT/AQAQILoBEFzjxF4ooTwrDzlpdJuU03ZHGG
Lbte3h+TuFhIkFWU37tI3qIb05hGTGys+isDClcqcN9nub+PfVB4nUz96sO6nsYg
y0xyISBpNvBZadiJXB2gWSuceqrWcPfUPmT5GizqBesD3yJV0RDC8p6fKzOAH2SI
ChE/lM4ocOOGawQcno2sWsMgLGEAFc+E+ufqAMRub5IvbfWiTb9sGNLGYk3sY9Px
2tqCfVRUNqadGuM5TY45DdSbbqcuWYDuAeMiZ0jEaX2BDjpnQzjZRTU3aJCvutGE
My4WRc+yj1dA4A8wffvx6lXwZyHn/RhN0P3Vf7/WkNtp6iqq8MoeyZCkx1EqPhdb
Wqwwf/6u7QrKD0d45D8L5VEs8lhLrjm3ZJH9spXKYHCI6wTphuhCvKFYIcapQxLp
zfEJLT3FTgDzXIPE96y31W6Md+GvFB8ZJR0o3txIkhZzKzcWiV/CGC8LiiDPtJPr
+/g8Iwalq2smgO9djOd8y+3DVm58+MIk0poWsztxYxFKLO6gzjwaOvR4srsYCMJY
LkHle8dmw+HHSC7224f6DZ69m8+JMYl3kVl4Wefm7uFtO5pzbgzA0hIF54UmcfVM
xiEBXf6Q7PQlS1wsSdroF9gIZU9624xcicOq7tf7d9z6J6JqFa7OfPrGJhZs6b7q
7ASkje/7OQCiUeL3gLaKLSY8QW+Juk522iHNRlvQGwidYfgiXodKcDwAggMAV/cZ
fO4BjOSUPDQL0Fvwp/rpxNzZ3DvwNePEMTJBCXK/hD/MjwTSqfZ07QVWJzDKTgBY
IfA6PIj/BwmM5L6Lwwv3fcX+fDPz1B+UCVCOEGjsG8Aox3/JkqEiEHGlRagKytcy
3KozbNuF+s/G3hqUMPmVtQJfLoovFYuxuoBjsZR46OvmFiVqElaZfTlKTwKFpgE6
D0fJx5AckX4NA0Hl8uWpgxYaSAmT+6yO235swlHPOE2SQ4VRIdDwEpZJ4BFojBDR
+Kif8TEsHxRKzOIlpWoaFRow3OWjyQcQduvFxdP6TBN3jJuOb3FdPow2K3fpM98X
iiVvrFY93nBuvx0n+fIsXf16JVbYnuqbw8ZJPS3irJIi4q3q8j2bRDwmzwMnnnqO
X/Hg3+DTX643E7OXcBjgtHy1jFsjlJ6JOw6F2oUQiLEnphMFfuBLucSRgkZAScwl
UP5cVCl5v/Y06wtgnuHzctTTjLoS7b54et0prc8PZHyohCnTckgUEl7myhAWgywP
FBngTVPMLPPeiC4fdhLMNActOoMMCm/D0AyBUavL+wF82zW89VBfuUVHFp8wLB84
VINRWiuK06q7penL74tj5Sy0vYovHj0StQb/JCn8H0tEz/R0y29ky3eGE2wwmf7P
PFFKm/UhRBOAWlUdXtxSyy1QBsVjYn7OnX5hTn7IbOIm91Sp0Hp3/tDBTpYm2jg+
EDdu+47fA+m+T5oLbDcsdCg4MzTBTOzO7PK6XOvAZPQ9rcKZIN2vThuN6D3K1wsV
DJbuBAnnEBum3zziYYOgVLyNDFL5Av/grr5Z+rxRnVKABFohJ75wy1gDVlJAJ7Io
i5RrMfZsRjL4CyGg+4lXk0yvJ3ridQINzt2gxeKM/iBIr/lK7QcKJ2j+DKCtbKOz
TENzYsZlK6f2oHPjVM5kHf19Sbocdjyft91Dtxixj7GRnkHXkggEeNmL1Xa+YvK0
DVYhF6qFgFsdQ1Tqrn8RJvPyZ25cYwUAS+Np/nPiigWwalH3D786gwkExxm4VpaB
F1D7qE6RSFHFnmxY9umjzuED5RQRZu+feODxPYOnNCBlu84UROIVbHFesVqB803B
LLg+Mju3LmbjyIPGwEx7DEX0RwrKpu4t/6nVIDsORJASDaq//JZ8l3kcqIkuWvge
0vWchoL6Dsacdq8wc2mGgP++tJ+DsEyYWFBSS68jQocNYHc2l0kp87raGFXwLxxT
qMKlDoUNJOqHrkNj3g+QwgABnbv1Qx7vQM8K/970QNh4tcru1NCkhMgSrq0UsGAy
64eBxQdRyiaRCEBNzJ4FQW3/6TnwQuhvRZYLYo4zes9XzlBiyEOJIUm7UqRitLkR
Jagz4eJYO8sQ9tDwSj86o6+mUsAyJdIe4PAUJIHILsfiGjGfaqPrz3r/R3XOZe/J
clwKST+zaiRQAGtKJU1jkiXVtKEKVoOUgO/3CzF/LpXFO39ABxGfok7WnrUFxeOG
SGw0cG6KbaxdVoA3EwJMGT6FBVZwyh6Pm+4boWF8SGxIS20SjQe9nshrRCmxsONO
yqq+ULmQtXQs0Z4dcCj6xN/SoWD/xot3raaPDMF9M8VeFm6q565nRtCmhbfe169K
+Ylm9FwE19fj6wg6BAw+tVajlCjCN4m28V+Je0nZspJUXfsiqDRMdIurswKxQtN8
QdJdurqqfj7I28Zb7psQwEHyvEHMjtX2vXJ8QbJkIC7599B7X69W7I8EzBcVviTO
ojntZftiR42a/WvBp4KifA80/mZLT/SuU21BiB1hD+s=
`pragma protect end_protected
