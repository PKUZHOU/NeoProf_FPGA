// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
WVfZgzXCyCHLIsjgibaM0kBzhFQSywhGTQwDezpe2bJVXky21Pfsac8JATqK
uTv86ctUL0EXW6WPJYJhVhmUrLB7MgH7r4iHCb8iQg1pyJ/9DC4p7p6/jfvj
R6VSbGM36fP2WXiN+KXz3L4l+ksHcCOsGSvFVwbb9SB93KeMV58oEeHUhWVC
ikmifXCqfCDqNvSMxvgzXOqWQF8lKqnLXUIqvtdVv7JT5kaBCXXbQRupRvv4
1ZNkbxoIoTy3eRquQiQdbDopyYU4fmUhY2tPaJD47NEPVXbQq5doOb1o77tt
SiD2pKXAWNPsXfl85RkkFJ5VMt6JLoW4LJKidBWmgQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
W9MAJhvbddvgpOimrMk8J6X8ddCDaR2x7MZK1QbrQBxM0A9MJkyegJyEh0of
IAn9xDcWIcrZXGPJuHAgTG9oZLLPzuhCsP6C8DFx6I8GeVbvKOMpsnWrRjXq
i3IBySEttdVIk7RgK8u2/yeXXgNTiICqTocq58/SAwM/on/evJ3VhDxoJ9h2
c+YJPDvdLB4gwiDMDj8QBxxJeS0TxCpqoUc/POls1ouWVkYaQyh15NYKtBLA
ebIAAaodsvVB4tEKu8hVZg4ILsW96vnwGskGYqTGqkhtTVvxlFgg9twub+gk
I+P/hDKcKanFxKqAITTKAVdlXA/pEG+1+wMuPg05Dw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
AQReJY0GWJ8wmrHs5RB0L2h6QEx3k9a+xGV/wkcIUUpF9jbwDGcUQEkhGp8l
V2tQEMvSmti5+XevTJdjD/YCA2k2K6NWqhq3ofbkZeB7EDh+vjd32DNOySlF
Rg7NJblx3mmmqaGcVsZf5cl6cKkYY6IRTr9jgtscz0zLU9zEs0246eEPeQQO
3noM7vcMgjkS+iJ8vacntpYGEw81zbf7Eh3R6G9mXfCtKBnvSxjVQHWt7oWI
TCdIZu+X2SDo26c6FtK8vJfpRAYhsasq0Qq+PAjNqYpNtlIrCtA0sWVh26hQ
ychsawtOgV3K59CPdWhsYjBUZ49MULH8hT4r+jDK6g==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
FGoHDNHZjtBRipYRx2HdQBg0Ylqg2Lr7idRVJwqV78kc36eRL9C3gjkSahBJ
eOFv9JpnrldZdp+MElGL2M7v1Ghmsdw8iKvkHn+Y4Fhm9aoaj8zOzf2hlgzW
j3E9df1BFo+osHEy6ikkKAon2Sxn1wPccfoTOZh/ikJRksyCbaI=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
NpApG2rvlME+Q6UIViCDTCfyu0eYhvqsLTVyRK8QqPIbyZBRDdJJYHPNAAYS
Xz0ZO8gKpEvvE4rqpP64HhBoHrfKnspoBeiegps2cCjedp8NvxoKPwkiDuRX
ag+UhHvS6R6zNIcDmYDoeQa/uU8jQIbFEWbiTpB9WisUNF0YrfvH9pUABof4
XmQn8KZYMH5CBxumREVRmz9I42ehwTCYj5JeJQEDC6tP6zVR5adarEpSIpSa
+LegMItU3xP3AhxsBCLXqz5UgmoCmvuPZDqRgZIS6QWUfgG/psxDLKnreFFa
Z3JcoY2dSXH2VKHg67OtM190KHbpZBnDZRgpIoZWwIzifWsOpuVDfFUVYy/0
CMMWgNJQ3wFjz4vuGuKVKTwFRL0reJyG2ba/M5msh+87uqlWbtxzAtxNzHZV
s6IVh2vDhFAHp8n6FL9jAznf3496NX/qNZkaF4CazxYCLty2xc88I54Bwj6P
H1bXipOIgjbAPavf2JlAxcw0L5/MFhc/


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
pBL6TW/nOgxDbj6xQp1j2yE1qsM4+UQcSqsMAWHDgRZy20+7kfYfBUctCCAj
MNKljwpaxTfMscM53Sg93FNGsLPTGCEAbc+5SCw4z6xGVFXcajeAH75MFvJf
oircYVyV4L+A6lGgNbC2hLfuL13VLTtB6SSLve0gbnTMxGCilVA=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
nFQRubJa9HauEl06yH6vy0W9lwhXkhPT9WgCiX7y7A1L9lGt4V2BVCZHL+/J
xhQRgnoMkWwETONJnDCgYAKwKbbTrqrgEVG1rXj33qzKBWEY2ASzkwDo0/1b
t8TbBA62Gdix8aOo7i6idiiZUXIvkxpcE5Htz26ZU1IqINiO/Nk=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 12528)
`pragma protect data_block
sK2RHjIz5MQLnwtdpJTMERWhO67V22zOTlgK35Xgi/uHwCYVAZr4Ryg7xG8s
ywIUA3RMN817LGHu1Lmixq5I5KCFpqORa8CAWUosrbPXekhB8UCXdIHnfqVr
JzLcKoUN8I2uw6HMgyhvhkUeAttg6tyLIkHz2JYZ8tn9V1FE+NlExWThMbFc
fd4zRnUrERsAoygo3ZX8Un9o8EiZWrFJb0kRyfo3wznRaT00GYS7JkfeVqNZ
OBo6x/ajqw68yGlIfhZQK3dnDd2cH8B3IIySyC1cuTChX/zVz6bg/Qg9wBwq
ZkZeiOU9R7QIKgEdkMoBgQywMhxuM3x04kXMJviyT3e3e6g5CKPB9vqO4xwL
eYiS/NdMyG3mQ83/NluYkHaPQ4fmd05Y7KdbhQ7/lw2YIvUbaLFhRRkOjrVQ
APGRyS4RgE9rA46nq0y8xa02BaPnLah6SF//P52hFcekVoJ8BEg7GRdy0t/h
bCJ/1RqVLS9TK1ORnyIeOEwwkKUdCbUoooeTV1b5zbmGxgXqzi2HnV38AFVG
1RYKE6gV7C8TtZl0wgRYg9VJmY0/UTnD6kJbvBcxcUKEMS+WXqWNlK6iXzR0
fDYsGH5GArEHrmWnavk/ZvapQ22lsGh8Z35aR1CZpF9FB3nf2PqAPUoQ7Rwf
uA5hYi3Tb6j/i/m0Bqd7Fw6NGgX8cS15SLy0n++WDr7H8YJ/2EocFEhKNJgE
HFwPUmk/rmflfaD6VCjpBbfmp85RVhduIyjtmGPfuhsrac+t0+YFa8n/l8Z1
gmL9gndZ506luwywt9vppyuVsqPI1PPZ5ecGY8oeCD8G1MZS1OxHGW+mIkbx
IizaugXV2cLKI1ldl/bbGq+GcQD5W6K/hLHVajOfe9UT4OVvnkQesPZzX3lH
acS1keKmAuXgJukeyueVRFcgUPFOWHZBS45pj4ks56nVVbpW9YEBDHT3DDIW
WVS0DRZspaWe4fiPW95uk9dDejRPB8PNQcO2d0U+RQwfD9QPS5YgzpgYeT5J
VaynVYMvwqOcKrkIgU2pV/xkAWQk0o3WrZihQ/u5AfGQHBOsPW4XYExf/9B0
/vtE3utxuLUipnLPCF0uZdYs+L7Uikmv2O/pt1yVSiYC/dXtbROt72Y4ewEA
YSa3u6T+r8E2EHQtP4Vd+a5/D8ETRrodjwGRr7JNCyKuJdDj/bM9GvMZOX6l
Qq1rBNpnJTrhwxDea4BoYX+n+WTyhI7RwQgTK4sHroodN0Hvv29Ysr5EgeiY
B6Pmm729XekEZuoe0hi5y52BI/mPUSyMH7NiSdX+gGCty0gF2JT0ZX+egQeE
MQMi/jOQHh9ukjUaqsyk8bSdtY3K7tF7UXHFm2cf2QiCYtoNFccK0BxTt3jM
+PQfYKE1SS/Va/hdd3dBJceE6347rpdLkbqjf/RTvC7MXibB5MSrvXA7P8BA
Q0ViUP9W7E6av0MTiO9CYCAzg1WtQiNyQgdzvBaYOeYWX2wxj+vUxgBZemHR
XyHMJs+She58jyzXx1KXc8Y5dScBaznDc1JahxfQ/M08e1sWGcCZ0OMqkXBL
Khh8pvN3uHQmAq1wZ84KqC5NiV7YO27ZzvYR5bW96LRiri3wGhvVNVI56MFJ
usbhZFdAWafiyP3qwg11emE/yY+bttO+q+sSXDZcCkQy2ZhzPgp7LKPh+sbT
uIz9zDgC+J3ZBJJ57t8BwCmrBhm/3dk1rjB7G3Tfb3JvkF8HfP3KHvUkBOmB
ms4g+MSKhAjmHAGuCWz0Ua+9mCrOhlG/Z/t4Be33fdqwEw2SVH7rFKlEFwGI
iB3E8vY8GCTRiAGBEsf7qWskZYwOTU5q2RVMuiAwaOwOiqGK0d8p425tjbrk
24ZBPgfL2ZWuQRSA+ZTeDpLufdCViLvzfdLoVTc8UXY3U3cHlcsXb3MzVleD
8Cl5ahji7rjhaN5Aej0bk3WVFDNU8cAvKj8cpw4F262d9G7WFXAR/TWfw9q4
9Z5Yy18kiBb1Tm+Rj5nUT79d3qQrprIsYngOY7DCsHVxfX30tzdYUmgihaDK
gmPdAIo4Pxyyf/refBa2cj2YNOGo5TNYkOAWDdK1JKK5wA9jtRGddEmPF7Rs
gujJ2V/6QuYoB7RJeef4/4Yb8Bp8p7TcZY1oGoo5Gc2bBg5t7siW/JU1hSyv
FCN3vyM1RO2wVgJxO/lbxiO3IkH7XGUKA6H/2i2Y8rm/BQ0A+D9q2/SDJel8
Wo7oVyxgD+06+NqiEwtwY+2+VFDzjFbzDKBBvw+lG0xWaJG4NgXaFOHsw7bO
QZlLEcr1A+SuV+uXNZWXUghFliIOQWI2npX6lsnhYShyDaHgVQsLY+RZgfdD
J1IIcLDNChSE7NGFlMwv5MhkWmWG3kCBLjaOOyDXYQGoMkAPpUtd04uAmhlF
cGNhiVAFFUU+2MIPkKg1nTSems5kmx539XrKG7lqkRIKPf8/EKHtRTgTQY86
sHCLUB3ZFQe+ZlrjoeOUX13/OPsd8WYHjNuORjbh4OrSnIvV+NseGvDOfVdR
VlHWHXa82QljDpbDbfwxxctqnJ3Dw+fDdlaEX4corL5Rm0eDiJqoZRj35JDb
tRnmn2wvYPQXTwCv0Jrx9zeBE1KVVQtoiaYWs9jWoSqk4wrcR2Bf4QlOoS0b
FUoMxBm2VQ7dcy/SvpBxmLHi4+tUoPevBS8vtMVPwDcgLZ3//WCzYmIRmT1g
ndmA7q8yHfL6Hq31wie60E7e2byPGSfq5iMyeFWDCPkRDvRFF3x41nr6VXkR
JJRRlbdaMkUlCvarfPTQOc2+T7kQ1jEjflyLbvc0V1lYvqXknKY9Oo2Ey+Xx
iiMZMF7yxzf9OEEkzYl53XdSCaVsaMGoTMu7c3N9DPv++9AAi4w4tITZbAU7
T32BAsAPQnVcI8GFje/uTuhJ8kD4RmfCSChtNnsfZbRf02u092yEQSVVKBXN
CoQrnY4JsJEtqNLsI9zi8oCEhK4OrA8W6Y2RaAj7QbBsNg2Pnc30G3Xa/Ps7
FGhpsI9La6OyHheJO0bfnrFxVWyH1gCdn17fwkLuGkYkcy6DyO6RUyLFw/Ee
eVGn/j2g/isK8eswarYTe5DK5CKBFdCb+IASL0cQOgOvO1YdMyoU8xXi8G3v
imIJE5f36uM/Ci8kuAId+yzNxqfYOc/wu3T6m0uCQqlRy98ojxLCOwMmZdEC
TdchMefxRgZodI5tyM4KGh8ex8yixh216uHFFCa5Yp142BEAlmeNn+fgV/Xe
RZdnV2++8erMX/8ywvBof4Ds8P3MsrCmJv7srO2t9r+b/V/f2xYLKyalnGxf
XoKwyaEUuiIhvXLGRbWs5aoWZVWWZFVrHhWbZr0hpml90SzdPJhZAr3AUkvY
Zp8BZWCU374/ksvPSbscFEpci/gBWDMeOK6M2ECA4dsIi09jmBJCVSNatmDs
/7/LdvT6qFI5QiIA124BxDRg6nhGhgG7utHXsW7splhFoOx57abs6xN0X2zd
FBe45UYLl36cOxz+q9CYBo5A7cLOQDfVPFdhZ2+ZWCV5fPFb9rbz+NsJ4XlF
pMql0rlKDmLSiNpSuiAGp8/FY+8iQ8VuMCVgd4cDPBvRM2QeoILJdnx+xgAb
m89KPj9eQrc9jPWf7OvyY3/z2tckgTVyhH3N0+Z+wE3X+7+lxvQCVm5vvxwY
Xn3a/rRNQNFLmTFo6RJXuBieOahe2/bsaURVlHrThLvzCBsVAUOzcCKr+q5L
pxI3vcrohJ9MT5W6GXxgBkGzZqBpoCkw6/vCy7aIDAyf+RKkxgV2lDb+i5D1
b2aX5ioq4OqwzFSMlvN+5eOQgtXX8PAtcFC/TVIv1+W2K8qv17Hf6m/Jz0SW
iWslBYlgXDvRkYk0EwWQfI5M3yvmOE2aMX76w4lKKOB90qZRpQZYmvjvAD8a
VdtPCpYboZVTOybV+XcutalJ4QU3TQULFO+WFcxFy1Y5gNb3Y+NN2L6XxxYQ
p4fwpOULmWxOQwWwCoL6CNdh7On4Ggc//X2cx7xzgd2AqnlVfGk0xrv3cIAm
DfMiqSTZP9pxyaRIcHezYchSxV76S1afE/F023Mpyg9Rhyr6qVDcI+kAQR5I
YtsZgT8MjGYeZxFAccAdmPH0+da7hU1+LxLejSd7l8OoDjmFvTMcDMJLxcwM
FYJ/kBrd/LEsX0dB/2rDSGQ0ONqooQZiYxwYJ8VuMMRICmDiejtzfehuMecv
U4zxpWG4LBlO7+CN92cjqJg8ndDIz3jkE5dsHRlyIpUG516iOh84vKvsLiLX
qEVX5vXATW0XnHnjdt15yBVvvLuNnfIvkuUtc1BLq2Eb82OZxBdT6Gc2Ksci
xPfiE4T3I4rLPwEPJeBoOfgB2xhuw4xKWjSQYUYVSPnDc61L8ql+27l7OJw8
IxNbLmH5Du1w2KvMr43EX4ZCzX9K3t+hrwfsX7z+8/QWO17kGA/Vyxm/a5zl
sTHpETgebBGsP6XHkBnXmfoZxyhb66yiJtRpYAdzAiNxFokxD+nqRYluvWQB
EaFQL2E7nr1wD2kO64XeexD/Cgl0TgEowr2eqV7O2qBR11oKK5Sx3epCbUtI
bQCxTVBQwOLb+VcW3E/6qrSOOj9gKWlxVl8EZDDvcP8PkzhAWeIt7wBu16/t
nCYwqMODYyvBgVG1MhWP3CzVdDeEDlW1b7jGAOeUc/1pSd8QVzOPJEGrehYx
MMBg/D+O0ri2XzMIbILZwP8sGSB7HMVWNZjOdpUjvc/KPFEk0QHjbfFzs83z
s0KmwBqp0M5FXiINikUZ3JDgYVKFRCCOvHpRFIDlGJOW+Siv3dJc/73JNpMv
xAZCLMUy1PF8QM8MtUs2mMawApRi5ME3LWup1mhronLCor5TLI/krYrDvWbz
tfbHkDWzROxhoSK8Ay8xNtYeNKI0wLf1ZfW6vJgtWKfEUTVq4l4R7/wsSe1U
4O6lcA4gbHda3Dsz0Nd5+wwqzoxh7yNGhrmoZ9T1ZbhmTO7apNjE4wSMQzt5
Auh5JyuA8kk9ZvjTwVEdnnkotE8aSvYxwvoOM5QcER/xA5EoI3NKlU5WDh7A
uvDs51OZa5fWamujr/aBr1yTxiMwE7G6NYAnVU/M0RASPjQMMDS/iY/1FpdV
RurqQO/x4axBtCkjXoieccf7cKnd7dHk5xJSLzhYemRjZ33Xp0ms/sHOJjxV
1yzUaYV1Hg5Zrh/Jf0l7o1aOEhh/GrCIi0z5k/U0JnEMAN1aKnCO5V7ssKMq
LETnQejePwD+05DM/gI3qDxhq1q38QqVOG/HiFg1Qn0JIji9FUGRq1uH3Zhx
1x9eFX+rDkJ8ADwmF+kvp36YkntiVk/rIdkTctVIqFSxCZ7CvxIn0Si7tutr
6jRakvPtLkrheSfVaJCQGTy6a0Az9KW01mvgqHsyAanYcgT75VvyxQJqYt5F
Qr0ZIFQQGZJ2WRZ5Jnw5X37BO1OqygdbCiMrtfY08dFdhpS1DdxNqmNufOk4
ieAcR7OSkc/dsHyHh/laQKA2B7tWiiBTGSrV8tN1LB3UeWYH3QgUyvgWF1CK
1Bcp7XfHYJb0QaoS8iKlfK1pGE3SOrJA4sXxS3EVvAie+ORwAc8bn0oJXvqZ
GLznVjL34psS9ohTPFryGBGqhg9Ijjtx34dwRrDc6An0+1G9oyv2HYfyMMhL
ExqBZNfR63V2ZERJow3eK6m3m6ABdbgDuZ7fJGTKrOohjHCR9ESrv4vcjRrX
j9QDNrplObeNd8qcIxp3B50xISq25m8hlEoR7VCQMAxeb8a2+nkBSl6fS4eh
JDtnG96SkKv4Rw/q8XJDfEbhx3LmiTWwvsBwdY3C4N6pKkLLgatH12kcAXlO
DmV/aryRA8SR1jqy5lYK1hF9HSh6P+RvAgyoqfsjIilieCQbbx2m/60xqogZ
i+M63gtMB4Nvcou5fF+u7iswODXCumW0bIWfH/62dV4LPgq2uVm+8rwkkg4F
n6bGPuW/DGcC9Z+Lu3y1BMgEECe3vdIt0wtRzE3EadFrpFW4sq8iZofCgCL2
7dONc9E5GQnfgw8vZVGKzoqwAhs5svT4Gn3i/y4kck+ov23enKHw0cR4zsXZ
zgPX/TU+yesDVH0wWainXbSNzmQwLzov2inj+EtFFpG/X4ETvToT2Bta+X8k
IiX9E1/cbyeShkneBeK5DHEmiF8IoWCYQHuRwmtmwsgs6efB6iLNjljsnVfB
CSip+pGl851BWBXIn7QpWykVdpfhc8EBzHgR+yaL7OGLNUzXyYiPqqAQDJDW
JgWGFI66qnvDPKzBOZdC4kPFsUI2Nq0Me1XM8YwvJiZE4Iehp+nKbX+B78l7
dGhHHzOTJ4J9GNzQXTQhwAQWCbRBYy669W4QAyuXCHK9XiFeFNurdIgK8VjF
ZrggNnGniL86x1CkshqrzPuGzGImdLUZT0oByctdorSquXBRF5NGX12nBy2y
OOYPex9kFN//ACHQ6czi/wOjbdxbQQwe+PN/3bKIQ6NFaC35koRIG/S+xcxj
IagO0t9nwFyF/uro2+w/E12Jubth70jp7aVNEHd7vvDoO8z0xicbIJgixkfC
CDEfBZMgVHUF4u2yF06A7ffdSkN/xmTF/mccMO0FExnDty8OnQtDGvxnQAan
HzQIzzyxk5dnJYB0U6i9K0/EeWltSSYTroVcvl88dKtM4KazdNtEgNcAyNYO
VTftRUC/d2kkJODoILnEh+bDL96ZktLqsQkJhXkNF/oQWBTxMeWFwqHcZgMK
Heyh8fpv0/ts7uLFL9U/88AZYPxT3ql8UlWuJ1W4J5T15bzoHuu3He/9I9+p
WnyBIHOUYUnIL8dkmEnd6XjLyfJiycTXERbm1JnM7m6TQ80EeyYx4wtopwZg
OnlECr4HkGvtHEfysveXnyO6qBoN1qtNpWSnKXGgWiTgq0o9sFoePvAd2u1f
aln+nTMicPWpEwV4WVcnc5uax55s57OPIFRA/etFNF0+cnfzIfKbfwZfrVnA
D+v2GCrqTeLbNFwrzPNTXE9PK+4Je0JYgKNu7eGEZOpf+pXxmE3xt3xCF0Wk
uGznRE2+/dnvYmc9+4p9gaQS49fDRsqBEfnHsp7wzd18wD+y4m4zVvnC+wUL
y5UH+YvZb/2bg1UMEpMQgmG1ujtJBsLSojSCpuAHxzSr6jIDeU+RFTsYAMa7
fxnR3d0V5Ii1Ahjg5nY37EQpn2pfDCrRqLQMOec3quoKiOQfrNkca9kqBNJb
H3//tE/3TRpFr9nBAqUA2DvxfefvH21p4rs4Xw9xzII5Jn/+O22O1MUFi4Ew
BknGRi89sgoWB5em974cAVkJA3NrpSYR1VwZQXkwY4AZzF5WXOVn1z4hxMSa
Q/fBUHbyj6TsTAiNkAqALeuZTrxnlTEPFbOBadX6AAw19RjZ40iQzYdblJzm
2qrmUe9U6Hx1NCn7BdvC4Mrsf74t/KnebsR7KtLijgCv8yfWGSgb+zvfWzte
kZ2I7sUy1X2D8Iitx8m3/QBuP+rb6YyIzhnbWmrWQl68w0PQwVNO7bhiU42x
6eerE/oUSKEfA8SFon1bpkN5hbOp5sCnL2DUFCCGLHJ1LGzvNWJu/o8XwQ2Y
EMWuRYmY8lpXz3fHCJg+yxeGDs642dNp5iXhdOW1ratRQ67TjcoEFrb/GyoU
ieu2OtmkOF8b2ByZ+b5XM3x4y8BY1ujMS2tay12+j8lka3N4GEvWj513D0bJ
2Gw/GFaXEh78m+a07SiZIpZJHVp8fVQabnFqMDwK0wUXoabN05FrmbrwMrh6
9LaacAXeKSe2+aMWhjXjZ+nnv+SjjNQngWEo8jIgtHIQOOVnrBzUxSC2Wjph
XwWV+dm+gO1VAsXoqAWdopRCerW4VJ15Ory8APNLzpxRYhxjOzcFM2qT+2E5
WQOgH+ZtLI0NjGrtD69KSs9oFFvIq+twideDa9TBVEpePHxSSUD4a/yQeBw7
xRExj6sNi3qZhZFMsafZ0uCQca23NFK6epzhx/D9qRBAUKIy33ckI0NLzLJZ
Q0Uoi2+85dGmTByTvbAEbDEhDW+lPwMvl+4lEbHBuJnlA4Sx0OuvLHD9CqoC
k/LwvaiNkLIL22XuliQWfQRZTFEk6lBld7w6oz8IjV7vzsYPti+ctbVGd7TJ
kJ0XhQFBfcPfFxqIoF9hfmUNsUZFi1t1uRO0wUBgW3Z1/sp4B4zAQZeX+Dkv
Q1xajWy5hXpvPN0JmjCcUv2898f4ifCRc3bBO6AdqirMHSROxhASMQVOVK6I
3C1fMlcbNf+4lzNZKXnwkxkpsIqHSc2Oi1WbS0NLgCuRKNXnXlc2Zg1iCxLx
+OCtKNm/9pi0A0vZmtH47MmaDmMb2jv4FeNswMtGLste+ncbRaGMRRBnSFH+
0CHF2sYUBiG/T+kvJLeOoS2mvsbyuO5ctJkjbaFWiMTlKolSl2hl72Y04MVC
bh9HrqOgCmRbsmBagc8sEcSoDslnpKfYnxq92yhqvX2EQmv57zPbSVuq6HZH
Z1jNUywGfMT5k4Ny6bTiV7ng9e437PpnmOB/O0jIvJawcCJlBZQukXCngAfh
LQbKBA76oUFORhrkTEFsBRsiQ/m8wFisfH3+4NGBsvCXSMZzv5YNX/p6QDjr
Szww4IjvFuCtusHrrHNK3FekcI1kNsb4h1UKo0NJOyFcl5XWopTqIwk85YtU
k3tVZcK0Y1P3KzZlLtwMJV5vCTnCKLxNiNuzgKuRH/uejf5HleioC56FGgza
YRMHDU0ni3HJvQroWnk8a1Z5y0liZNScW3Cci8iqdgxqeWX/DHS3nW3JKEdc
NZldFHo38z5nj6/13WlykHquexAWevLh1klTXLmfle6GEW4oxvDI27X0BAHo
l1kMUIGWBQ1s7CATuzMyCc55/EsqWBGN+LOk5I5T/DGTLvvu2tm1pzn+vxs2
/gRI+dA0+lJchnjZLGFkiDyeQkCNEyzYfFCPaHAc8UANM1At6+Q/vWS+63jl
/fw+B/TrS6aa8B2cHCdPy3akq+/pjmkHUEH3zAm+56FdDdJDXHoM1au24VR1
e8tnnoHlbzPsbVOBI2e19lCQEUks071KPtLEelVaL/Tv1ftjZlQRCGDCB3xZ
gZ1FgNbYzktiJEoMxWZyyODZiz9tk2//2a6OB5bdD1//pSeQOI6k6frVN/En
FJtA7TAYvYD0xmvNnXPR1gogIwMiXLdSWzp0k5MxPhTrbevx4ZdtxfqRY+ZH
GPWubCtyPStDj558FOtxjdJIcbyiA8HrjqLFHe4WCBteS/65effr713HTAzk
BP4X+T+2SPaA+/03//Mnpg45E2j1ly1hYGAWMNBsq8SrC2/MxuWYzeQ1Fivc
Wdn1h2x9tj9/lp4Cx25WpOVWwZBU1JHArWY7dsBORnKbZJwW7lr4rDo7A5r0
Cvnwclae+JZLW6BDnQzSJFXDGjyHxHnmJuuNVrNO4HKYExO9U/fIN6mJx7Uu
H3KXpg4RvrwwSKOS7Ei2DWSIW0fdT+yKpGk2SnAySbt9pv1qV3OZmE6Rk+Nx
g2ZrKQGOK0c9bgrb9Djr3IWdQpIwqEgN7DjIgim92gB2fMGp/GiqShpQDydA
PdyPK8LTBNP8Oj0rc7a1Ay9G7wtmwhRgs+uY3asr4y0jna/9FCZcQXWICB7X
HiyCPfw19Pj+16tcHInLKBpA+SZu+Qbpm0LfkzUYx6Hl2bvXt/SLmQ4K5tFG
JmrsTHL/Y55acpI8T2jXMPvAfoDvnSbWvpC7YyLY55oIuZRQjUBd7jO/sfml
3xI1JPYuK2vdD2eEjWi0B2zMsWKTaWIV9jB/3H5i/t3YQkXNvt2s52qo2zB2
Kn+dA9nGXKoEjFtEfdW5ikIZ/pxYw8UY7/fhkJu04bkPX9iK6qzLp6f9SL6Y
zU4dt9R9XhAIC1xDh6tIFu8t92yA2lvKp1UdeDfbL+CvK1gTKXOqht3SVloI
Cfl5Iz87hqK+afyjuEM76+cW01/jacjqOn8Qkovda2Pcv89QS2KYjEF03Dt6
uxnJY52J5QQ78IalcHVEPyHmFbVV22HgELoleEwaB2PR5tVHDGJIc6rGbAco
hNYYhpnP6hSklBaQzNdCYcBscbyoxixsix9obdl4KzcJe4hWn4k7ntGM2/0Z
kdGcn6ioVq2Qg6fmURlRJokSfbeVwRtERKRVMasitkj1uEcncYslP4F/+nvJ
cqEAGcfCX01rsXekpIryI8J+9+Fh10IYYDOvHbKNAUQEKAU/2ZOnoaNMNYvb
t8zUfcrOS3+RpDLJW32nrrUdD2TfJ9IwgVIqlb1Rr+CN6+8QQZLw4vqnc/49
vTzClIXmuKYj2PxXXwkXQGVzaCQmNQ1nJgbhZ71acat94V1Ca9lfq5kdqCGU
jOOJW13mboNqG7GpG9J9ATSgZ44AHcu+UIgX0KSD4P0cx2n3Lz1UJYcdk/W+
Z5VQMHAMcFQKCRxux5XVLv2i/L4ElobSw0gcS5Dj+6Hpz52pi2qYml3ocDDN
UtZ3v7NiBeJcejwYQOv+jZb1Vyjreyp8hk5fH+JJTD0uikiIaIxwYyzWHCb3
ZmA3Yj1YPNwSrcPbgkO8U+F1dq+j8mqMHZoFrWNgoLv68ZvQEaqTf6LpDRz1
ebKRf44LNJxMgh9pLDJjjxRpex/8uc7SXrlv+TkXFfID/Q2Uud+j+kwfkejB
VyiNXLWoviBBv5qgx6rmI8Sm7V8J4WFv/vGQYfmxcwQ+I9D7H7IcZheL81sF
1U2Nb6eg0JMzk8vD2BV5u9NzDYM/tGNLv8PllCv8nPuR2gIIsDnRTf8NmHdX
JjlERXn8bJvyeTUXJ1j0MUdK4uJSkisilgea5UxHwVcds9tBL6jq9403RH9G
Lt4G7bTW2MqirC3846k6JT54tphqQW/nXaPdq0j/L7aJmedXM2bO1RNzEJz0
78tNNjkexD/Yn12ZTSOfIxekQGx+aDbgkq3UMOQNRJfwKcGH5ZXm1bvixDcZ
MTyg/BxbKAw/nFWjIj4eFqmE+YaQXt2kJSdPNKMyKWY2VW4O/knWIcYaLVAL
WMewlP+MFpNpI6xIyS5wjqEbC2gz3yUKG+VBaGAL+GKk6ZsEZ2uaaPE2YhYt
lHU0To7GfgYWIzcO2Px7aVI29G4eQ91Whilzl1BQWa9H4MIhl3ZSGYo76b5Z
xjHB9NzgH1oQUmPhKG63HMJgjdIHaNMRhKF9EgZgWvuZijAUKz/DO4Cd1KVv
tZWObGovKLEAwhvky9rOKA2LzdXic3+q/FrYfX4tRfIbX3DD6gx5RnVM3PfN
JD2Kr2U5jM5LhzwFyZzGnv8wxTHXxmIdBswg5r3UiuPLP7Jn4eKQtyu7CScw
6wyBkFYJaE0wId1NaIw0jh6uw6FaXn83nlGbhAToutmWsd1upp1h+nLwQQ2D
b7DLyN7U1ozfcrRC9af8vXmXA8gq+brRfiRF3/ibkhDErQHnp1HLnQta4LHm
4vnr7nyFauMMYVnYGC6u7KjfeXhiTzBgKrhYPcO2Oz4QZO5CTkZiRfMnxTLl
dd1maocTFBQDfYB4cv8Cr3NWcMr7Gnzpk5TUFM6FbQtixWbLzzBS4yzBvSOE
tvgK6usYXhcm0KRVEKoe34Q+hvI8OP2Ep5f2eZICObdaSeiqs9poWq+TFjn5
DKJ02JGm1fA3CkofHH1NEh9qoLkjyL6m838z+ug9NF9y9EwiXkpHaayP9WbW
/uCeWYLm/f/jVxRQOkZZaZ6xatSroJZ5aAOCmkxr9aT7S+c/7ldKdYcqQzgF
DGvDqhdKJvjC1QVC8OY8skHFpeGvUxYwP/kTrJXNH1qV382K8FQxVaSa3rLf
gVjBrc5eka9Am4nksH7CyLibuRVcljCBBG2gBwIGwX+bH8ShM36GCXg4FEGp
8zrHAITEATqQNiPU88PZXlrtqQFO217JIQcrksWXMRm2TzqOpwee1R3LH67l
RU2oIXD2WlIE47uehqE9ufGQuJojozfRedJiDl72A/OCjHWVHMjdG0MOJt5c
MRpAaW8Likh0otlPDcFPq1UPd5JJFFexSBu0ZT79x7ygafsYY1et9oxdgLuf
6YYumHpnNg238wv/SOGYqCRvANNrmk5j++7qLbqnTg1sywUfqKs9RmtH3BM2
fMWZCKrQ7acXQ6WrpjWJ3RVm1kFx7LC6FnmmA0RT5Dfv0Y0wu0hI3jlZs/JP
KRkbHwPbqKFCRnug11mlTYLhBbWGOosOBZl1PWC0u7j3ttKNcH15Wk82heKo
Ix4sSmxw4vVH2q72/1SSQ87wSl6lXx4JKmVoaM+wLE9QFJglloyjFANMiyQL
yXfHuwEsNWuirj6BQG2TnEpxpeccbbxYgk896LrrVEScxa2U64hGjRSAHX7l
tDyHaR1IyYRBz766YMOCQ0hxhkSzKqf/zn40ZlvdRlGI9A1571uGI2d07BMs
6nTIM6Fein7+FGGq3uVf/JVs7S7X/KV4idDf0cmjGGpCDTdxXWEhG1VKYmJy
RnsGcQEu3+4s+88mvjwIFdf8ZimA6S3KZsI7NMPo4kqV8BEOJyhEpmo+kn7E
qeq95sE4RTZ7mUOlq8fNctNXXFZSs4dkAQ3uIVgOFtQTNh3qHGkDKLZDLfot
HC7n+ZGQEeVJU8zjxyDH6NRtbftYCpX/YbW3EwgulSrWxWPXRz2hjznJKu+E
/tDKGZY3CK9UNSd8j+Rau/crlIkyw5ZhF5wxEkEK6iZ4L1qZXyjbdVm5sQqk
Kv4s5zWl+QCMYR17bYSdC9bol6/1iPmWNlybQcVfK6ihETPIX8CM3Flt0tYW
PRhRQLMt/v8gbDzyXrMxu1qDZTR28tmo066jZFBaVu87SnS7TcFbhpWr+kRV
hfQDd7ntSL4Oy3iKJSYR887SbE3T4pW2FyGr0p90U2kN15I8FNFMp3+p2TgV
jFDfJgfQbIIlxrz5H62k/Fp1dtMwbFcvZhwuSjeyjU7Je1R9f3SnCYtSawFA
FRMYb1Ej+xpFZx9SolFrmh+wUXJfkeDtlk8fiaixcYKGxtUJH9X1DGBnIePK
IuTloGLyIqBltKWY67ZHoZtQr/8Z3q9N9cZWhzgw5bC/Qc/2kanb4B5bQWc8
2X037VgYnAI3ktpAt/trOJM7bkR9DCsVw8uFQcrjvrEAaSJ/0HNsBPZUxrOG
tjcX6a2oSJ1SaLdCDp1dO2+hwWpxRVKQ9NMdviVpnealxYQdMeQNbcjD0i38
xIkwInfnUyAfCtfL+b0LepcCRp5mW7fRZz0fLYFJJQ+db/t8I21pBm/yuERH
KW8UWzfHJFdrKzGRyCBLthdj3vUOqGqd+aU4xSjR6XZFlUWYt5RsVGtHSN1w
lE8CA3Dbk5ggMqlJsH6GpS2SFwf6xskA3+e9FB0Itk/Y9T2rfqFe/cDXXc6y
O6QJ9+34IrNbAHY7s11jlu9fUwibKkx43nqBKqY8BQqTj8ltbg7jRSOQVZfj
KFnrXdw4CgQGNkoKd2jdI8pgGbXriv8xkFk7O1DRvxl5sAvD35A2znGFwIcb
1r3TPjUlaHqVv23NEd/RIKBgYfN8ainQ3DDL8Eq2KgxNjZEYtpg6hIA+ameB
aPGIORf4wpfg3GGBMANUBLnJrVMtEo1fvUJrsdBnixSHMAaZLz4TKZmJYXkx
MVOcLsuNJz6Wnm/7VU1/U2O+z3AKDLw0wmqcs9z+J3Z53zhCYVYvlEKe6rj1
yxEGR4RxvXeXUadEBenqn+kJamENnMSW2JQjvXK/3gAXu/ZiuMdOmQpoDW7q
4p6S4mtIU1HUeOmbqbkEzZMx3Npz5jbKUQOJd90qb42IF99BxEhbY5LUpkjK
ShYApEI0+8hS7AGXkNMTtVCGMpqh2Kl1YpyPZSsYBrgFl+26Iwx/8qLfpo2p
DerI3SaHWtmZ9JZ2eL9il5u/dDS7/XasP+jlmE9qII6wfeG41LiILR3fhbOM
cJ+xXcURj1nv6x0pDk+7ZPjgua+OGS/OciNxWvHefN+boXIomYuqOG88/rEe
h8fRz5dazEKIeBdExNZ03IsSbpK5PcaJNY3C1z/vWWAzy+J2oZy7VHgWc+28
VfSYInvO0m4uLx2FUkIoXoK+8gzDlcnX7iGJe3HabD06bfuZXvWafaseYXQ5
+qSOake8r4Tstv2/p5WYBot+L1LmwW/Mi2evOBMOq8h25XdNhqE8bf6920j5
CH1cRsunqqlOaQ44qLfR+mTkjxdBCaLfuPPh5zdvkHZa7f+POMq7/9SAGXwS
JtRorbmhRlosRVd47ms4KwEyCazgG9xmVqnj3ujlAolgTmnDlghu4MYClndG
J1M9F8QBLTZF+hIUsCr/Gj7FmurLjps9GiEBWtc1SaryP9oVe2NpCZv3fwVA
ECejFAbYF4kxDlOd96SkVtMXTRCrg6imOVCpbLmy7kDfyaRDwf68z42RoiXN
DUFLyr+4pbW9CandcNW0K/SZf4jRhmzm9tVag8NpzrMQoJYyESUxZkqDf5wL
9c6M2abDZrKz3lnGDIvF26HKyF893JLPXKWHtTL0gm8sR8CaV9Vk4G3wqDFt
k490s3e5WQ1YAEuH4rNw3GFquj5DooaVw1P4+42FBRFb5K/Qb1PVy2W/bw3E
w/QGtVASLDt4+cppDsk1OHKzYSKeEgeSe/MpUxIJ1qGRSxEFYF8jBbsLtc/Z
kxE5pcpXjPm2Z0Ny6COVp9swR2itNwDDwDVAZ2ZkCjIliCkxaQsV+7QDzmG0
CKRRz+TL87KQHlKsEMOLeH8tyQJD0271gcrJBg3ijcg2r244KAr+pBDTcmKt
SPEDuYlgh08k8qlGvY+dLArit2SCvajduNMuiiyfDtDQaLRovh3yFt321yEY
RfDXGaO4QS04O48I/r0+80vlXkwCnzgGVnCMCfSi9E4KcSjHtsGz0m6QTORN
3AU8fBYw9F69ll6yzGfYMqo6oXJgIrUkhzUq4Iw++s9O2n7RBcn8Rxp2Ucao
93QaV9U0ibkDNP4KL3e4QndftUjTe0LAkA3hCZI1ElSVsyCdBls8tGc5zBBS
FK168dOWyaIMLaxDkDT0GIxOfwKq+wF9RJzoV4+0NFXczcHsZPFbm6FYpfX4
hziR6L6qWA8TnswQcSuRG0Yq1l4Dk11E0JrF95Hb/ogQdvVs0pwcWpmqXT7Z
FEixgOetx+gm45N6Blqx8UFtMRlpERfK/MGQg7mszW24ZDbXmPrHwXnA9uA7
OSqHB9K2IEEOGKt5u3RtqC32P1UeV20ImmfM5sN22g91ougR0iTs4spUI+QE
0DE+WzCU1426tCRvZSfY3DHAHCTtan8DIJxrqKIym2ilbdnmOQDoiqLir/D/
Hp1Voej8HobRrLKo3kVoRV2/dVkvvVeAfIGuY7Nbn8e6Oe4tDVlUofv61Dhk
QRUgrNeUK1eD4XZ3WxChLMSrge8WXwlDX6h1nM1Rn6S25sDcoF+5ldROGcv3
auwH9Bm2kZQ6zuIRAS4jhnBq9QtOm5DP6byUgsSJo+WP/uZ0egbPaSh5kFkk
cMxG26adxVObOPZEzqJKlDQB0mfCFLeou1dc6GBlAdKDMoNmUQf7WqFK+NE0
Qe8jYV30WOtPkBZNC8nZv5hl0DskSyPMe1BGtQ1zsMSk1H5KVIPozqV5bLzQ
C6XQ+9JK0XSk+82Hp6dLJkqFftUR1OBFpQM5fvmFY7i8jrdflEhGIskAEMfr
eIuWIAmBkvjFWRVSJehY9V6h/89TmrHmSXHLsyAI7QJH0BJH8gxnxEhjqIBM
VxO9UZNDtrLFenkGVdeoZ72XmfFlRfKXKd7CKq08guC0nE6rvVAQyp8wdXvi
5x+bQyxIgE6aKM9uekL0+JQI00Rue9wLqOqkJxot4FQw8QOK6DenfQ5IumOw
WuLHAFjQLpdmrlNYwyfHkW0UxQLZ0CYF8ycbN4qjqUpl2SOJzRUJnzty8OkN
jia9C2v9teY4lBmDoPZny6WBnR3nhInXmIuKpu+m5Hx/s9dfGonNcw80MkTi
lYUP7CnScHPAgD61xDf2kqauY5lHPPB0seUdM7yq+mVztlnoUt8niVjt9XGs
/RlIP6ZK/I7SLqdTx7eP8xmykLO+6jgzbSWgerbFSZT+pY3UsDC09Mx843vG
zgP5LFBl26opxVdpjVL3/5tfTDJyqz1CgSyjPmYtG4TlzUhxitkisLG8Mxi+
rSuxIPJSWHQpoD2hK3BekJIVD6Qp0TAYgbcU1BSs8B+c147JK/TVhNHXxysC
gSnFb4bDg7HITfYeUdg2sM7811bsJEuw9d6laeSm/yq1ymtx7zaqMPGtFMo3
lxivCDHB0v3/w592t6zyr/H9ImhfUiXMfwljbbXd27u593uszzLsEkB4qwpO
dj+S6bhuxr8POdw62x69yPcZGewr6Ge1dlsYx5c91kHLHuFQxNDxG670vtkK
pdogQDZgR3+Vgwn8VR0hXTryFmj1q89JsZapbekfw30alqWvorzFn7nVlj9v
VRPOJdnAcjJpyiRFh5FIyHnS1HwTDkhwD3DxOVU2C2v4e/zjX67DfB98tURZ
k6/mIas8DjLcfrnEdvZsMIeFKGynA3OVvpk2DOjo7AwXE3cEQpnQT0D9o0FB
thLRzjhqncsx43xbJu+DZkAt8989IoLRYjzigq6GK7kogxAvbZooURbWZAgd
xafmtsw96q7LgBK4ppvK8yGjxgwkTr9V7RvDYU6oLuXl1OyXjMe6uucoEKEG
6d7Cn1kowgB+59hgmRxPtqsPtM0f7mKDNUxphNa4VZUFTenc19lpoI598MPN
oO8wgSDFv3owrVrIpk+eeyzE

`pragma protect end_protected
