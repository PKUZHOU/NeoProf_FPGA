// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
AaEmOUS1yuqGItFM/zehqhidMTzm/Y0hklp4wW2sr6uaIG1b1oy5isMeOHwv
ZQAi5Q6H/FbEeROmiW1B4ONpjzM1eTDssrcCiZg2bKJ9WxaicTOwqQG9nrjb
wmMIwyb+YtnUzsSO9EkbahRbYxTEeYEzneKl69z4FEskKygvV1dgXpm3Bx2r
wGbq9jOEJI2t1e+uAVOIRgIklP+XEGO0l+Z12M35MxEJ7y3L6oQKwRehM0rj
f9HUjepMqH2Y/TungnNCghLt6yeW7qMVfxRpFSkYtVKrw29l0GuW38pdxqHx
KYRuI0QBUH9bn/1Wb8rNAjXmygUQkZk/vpgIT3ecoA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
DdetC7vQxRz0chM1nvP504R71H/cprisf3Pos4w6znMSPaggNP/PZUJ7R2Fm
x4AKuRLSmjYVScJQ+enz7kpsdMVjZ13aNQ7P31vdE6+rgKRefDEVUR8V18ET
oDlN6S4VeldOK51dg9AvSZO57qzh50Kgfm5LcsYyK+qmPOTPO5GnueIXBNHS
MejJbTieB0drJglSjL+joyN7526+4Le/U7IFNg4ikZurCVRIslbr5H4yZOa8
jSZ5dAU80DpJoF4IIqrA69GBFrf1jf1/CRVoc0X5sXF+G9d3LYKfYpOXABqY
ozsr/Wz45mwdJXTUVE/3z4eMxNv/NIhTxVRUW1xmhg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
YfZWHnTbFi0ptshSIo86jWobLAoTdpG1A3OMUVriJhTpMN8KZ6JGEuaT4tLr
b6uYdqnUxmIkgRtdZc43MrOJT31XGBUJqt2oFdvZNViZrsg1oNpfEYBX25R4
wUUK1Ur3yzLUrns7SxjYGnAuO5IU7c7YgfxZZyUGkmOH6D9mE81pg8MsPKH1
wd5ANXGdu+WUQqV0i4zJ5LJYsu53T9vdKOCRtuIYOo9DVpJ+Y5RCHkRNRUza
nWsRWJzmslBebdPcYLyZ29bLtCabXX8UOG/lFGBQejOUHnlXHheh4SroR0vu
F5MHKfSYT6HziIkg4AbhKCiwphCY2wU5LTlZurpGNQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
JwrGDEeUTU+1EpW/xENTQ/rlF0HEEufhSbQzmLDHInhP5WEki+abxxcl7oZ6
Q2GRKsECxv6TsdQdRku70gdk2CTbHRqIeCCz0BuE120FmWI4zwiyNZdFhZbk
5vmFUNv/JJOoItGXCnX0dN8MBNP7I9UH2OqsoIbJ8Nl+/sjOXNo=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
n7RgGM9vYy3zZMkjw+KTtLUQSMI7o/l5LqxULtbQJf7zX2TVUB4HkrFFjPUP
mg8TSS+sf9JzY07NUt080OOYg+3oPadmAqj2fJSgKMXXizEu6TVFdEvhDFPr
RJtl9nUK1hYPhmuYDKhj8RTUYmzLJiLz+zPCB2VZd/11qQzTCQrunMaO8IqJ
ckOmcHqjbYV2jp+BTSsLLITgE55OK91Dv8TJtODTpjIk8sMujBuiVm54UBFr
vTXX4qrhUAf/aHXdpIezfl99UTiqG7Kq0oXEzac6UZuXTJFNm65rgg5iV6s7
9yABJ8jj2Q5rM5ne7yC3dMlMvUG8GVRu5u1UZh1m6VHa8BNKh47Rk8NAigYI
7UKwOg8jl26+7xQqxLbBy+jObmF7zZJWMt5+uAB46PfigoNXzEvkDFuaRtzf
W6Vhdni0zBH/5vVrpiaFD/0XN1osaDt1ZcLlMy7ObZgYLLjBuxUKoo4szBaZ
cn4yc2HBZq7pdAOnETfJQ8RZN0MExoDK


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
IwSnO/qiSzZLT5okj4ZOjixFEpt5AVlvmoOJXEgwfjhVaSjz3YgAXcT7vbWY
hAKI9kTzqimGBE4DJQrHwtclRZXFuS28RLquVtrFN6Z+wZ7bufOZ6MKWhl2y
DVxV8KmyxmxKcbjAA4p6dumocL1d2fdcvdP7q+7BN01ne1ek5l4=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
tcwo5cKO7/8IU9XgoDLs4rdCkqB1S/yf3TCeQk57HhlFl8mrv7jN/0/dYyBX
vtolzERD8sO21at/VwXgyESxBKnOjLw8LjncC0JnFieQsYwldL9dr2taYdt3
lbUkLV3oiMR+GH00VT7jDy5KQ4WPAJkiVB4UmCTRXCmqmydEg+k=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 2576)
`pragma protect data_block
EL5PaIgGku4tvonqMVBUvjvMUOuEpksBNHqeHi+UXnSWJ9ic6CLZOMzqCYFh
H/DmJqtVbbqmz3Pli8Y8ufQ8oovKlPFO9uGHUlj/5dDIQOQt7upvn9OWofc/
aHFjuNRhUo+s3C7Sq95q9S2r1lnyU9eKGR8HVH+yuf/ZCxYVFv1Q5YLWgXz+
pVUwPBeYEQr9s+rTik6LCXgxV7mMJEyvvAxo3AglR4Oddc6Gdb95mdbxwW1I
AouGCXNk3tUHA6A1ehPFKLQocxBajYJq87Jc//nZ9UMMQQH4u35/slOnenyr
1Zv+LVO3cHRHFZUxDxx38p7da6/qpi5tn3bsLzpL2H+e1LCBhya9284L7OA8
afbpJXqBfTi+/j+y/SCxThH6IAkqSNGKOrhySVFrk2UgR0OyPYJlX7oAfrkc
ipI4esGtZpAtUrTrFAc4fCIbDv3S06boz5FNV/MBaIzncBGzpEu3Lq929n7S
kLamYbMjiWCkBBA+xtM92Tr7s8etOQFH8u3fLnscGODnbx2GOBK2NXnHPx4y
vKrbmQ6I+qPZpDApGOoECKN/6E2Urpc6i8GdEpsIYqZXE1dw54+1+j2J1w8o
vy3oQdfv56UIf01wp/PWNaZs5vpeoxZ7+j2V6XZfgXsuf82fLOuBspK27StL
4cmV8Z0gidg680d0PWs3lB7ly+bBxo9aMW/FfkqK9dmipAWi4FPIiV4kmDVH
U020BdjNP8MSq0Uj/6Hvn4g1oNM6zRQPBjr2lZ/kftOPR3uX6ZXsN+WgSbsf
oH1NiJtoWHMh7/JzcIFqVFbH936RhhpxBmEOipM9aIam3lx4b2h3/cbC91bZ
b8bf8KmCfcvHoVeBK9jL6r5R1Gw6H8mx0WJIVua0Iq+riFgjnXTR7KCQSeZY
Yg4hO5uYvboM6dxSVf1zNKS6kp6NHnjAoFfsr+FfNKsTjkgJux3YlMZsahzh
GCium78qoQ3xu007WtALWdokdU3bF0DVg7dIt+Dw6kGuqSa9vLQ3cSCSVcwv
LRg/sEopeR2LbqlCwxaiLDL8gRtVseZa2s5PvQJE0eVEU9Cso1KJDwPbHzSI
W74U8wdIW9iHDShoQP6PiWUhJ4JXtYrojjNUHyTXLI0s0CrZLF9SsQvOFUr3
Bpjir4/Byjmzzap8+uwOfsQOHojstxj4ExDHEBEpbF9dvv3ROdzTyVIxUA2N
viI95o16NoMsa9igCzmsYFw6eunFqtJGLL8Voxucr3scC+aJ7rSi3EqCEXiV
3I056dNnd6J9nF5eCmz/rGVTaNFj5Ihmzo4W7SUVDNu+t1Ho3i4RNFsET4Zd
8maMUh/MCudOrmvk30UbRAp+XMp6L94S2lyxPBH7jHlQTZuPTeNzS9/OSMGO
i82xyK34VQ4qbq3H+lRXpaKkYa5FNd/jJQYvGHmJ44qQQV19tUBbIpXCE2ip
RBC6K/Aq82aQvS+mJkmeNXWw7YxB+QmbALhqdd1ELY7TqOiypiNAMGU+eCjM
r1kVI2Ly/G9Uxumy0o1hAF5M3Xa3Kc/iDQ9NfMluD93MbFKNvgc6PLxs595T
bbpUagPzFjSNuqT+WokU8ZX53E5uJ5S3yam9FZCWXbaIkqo4Ax/f5uFjLnhR
+JolnvidpdN2MK27cr3kjVn0K4lt0H7Jj3sMQTvmSJeX66nqjYdWDZFsNGxQ
sRM27CWAKzcIWeA5sEOoOl96gs/kpAZsfOFAytgSNv5nVOdQHqhARwm4X02C
V59vcUct1fHf2zMGfYHybCuFWCubPpUtBE0A6kkR9PxpSClfLgur9nJpNynU
gT+AUDDJJXNLRPk3LIo8VnrIRRWhHi0MEoOtyAHiX7IvKM0/QJkwK9MwcSod
NLBwAX2YVE2cuR3Cih9S4PfN3TBcR925T6D3Gn97QJqlGx6EJusKy/JEHmIy
FRH6sDB36w3xe8op2uvmQ9R248FuC4pkPMMJ8rOn27PsOtYUrqlGcBxcAH9T
9B7zIlRM1uGmZIAvQpvNMyvyCwT5vy3mxQJSjlsjTw0GKzVD1nunoserTr1k
+7kDrppWyDXXyDDaNkJzvKXYe0VNRG9CDgJpCAk3P8z7Ld2XrpndlL04nrB8
Mm2kc4yEiUhnluzIEsKXzdoelQcUaRQl5c6rtVu/MAgRPCBPeajWGTocf4g2
0tJVONJmF/8y5M9EsaB3qqWTGVueTG/syZ56JunKQ/CuAdgGy4UoXs6dIpPn
7hI9opN84JVScwd6Z4qDG4ovrM9B/q2Tiuc6GxwuXC70Bgcce/maRE1T7l0c
GOM3bVSxh8TCejUsmy1rih/xsl71xTL8hdiU4WdBwdBB/YA5SveyHnFzloFq
0VTfugl0lLjuSFX42aRGhU8q46kTn/vtyskZngFSi7hlbS9uFY3c5gGzV2VY
gb+98NVWm5QvzMb4M2Lx40aVMM+jr4U2JjFRPYvwha1VhvGwDF+aB3dSWRiL
4KFKG+zykmQDLstAzdf7gGA3MFC6eVnwH3f4445jdL9GCY7JeH90FontL/fD
SS6u9OpJoQ70C+b9Qlk/778CQ0OnKl6iM2dnUA29vEGzwOVkxUn4zIlvAHWg
3YGZ5I2wr+1aLw8YYW5z7zJ1U3r4lh0O8lRDSqqnK4IyEN1XucSUQSF1Wi0C
poZ320eQS5eLywooEg/zhAehkSk7iexojfQ9WEC2BTSFxs1/YszYQB2fOOie
brjjmAAHJjADS6GHyFuRd2tY+Xe5ec4mf0BbbUM3IaN9hJIANx76PLWs4Ld5
Hb0Z4pWnyv3w7i2i8a4uYqGstYvvPUCCs8FPEcP91iSfrPw5AEaVbOBdop52
f40bYCKMXLkIO/ImYepDXQP4d+icRnnGuru1v6HdAnSqZ8Y4VhIJ8X4oQa7t
4cNmSn/hyR55uXeT95xZrHnl/j4FoFZYCqL6jYogq3Z+yKi8Bi6KwnqBOt0A
jckyIX+tPv/8NFQpzdiNj09OkF16GJUL6LSw75VubZ5g3koIiV0MpkXx8B0N
e52sG0qeVnYQAVP2TEPEcT2WwYrff9Qx/Ne88jCIk4jibA/tTb+eb7EA1mVO
ZgokUY+0nf0NY3IjlBFfRlTJp8D2rIDC3+VanEwSpgvxxAkuU1056q5p/6Ce
+wR795maVZvvvXTYOt5mRVOOPP396C1ybXlJUi187H1USCNcaAhbVc513qE+
F2oQJ2ipzB43gBojDFL9fXERWlyhux/UhX6CizDOzp/FbD6abfAT9cBgpaOD
MnA8kEOSKThta8O1VlSVqn3lG/yqqHA5wd0sGSEaiPjwPCc92yqjZ7/ecNr0
WQ1jWL6LkRBjpNsajRc2nhgn2HNC6EKDcSWl+vz0neAwD7UCCLYBabUaCJJh
mz1CYZsb8mcLCpWP9LRYV76/EKb5uI0kJeIV18OzMKe0WPvmehrOeUfcljgY
Wnm6uruze9cG3Og=

`pragma protect end_protected
