// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
vC1IyTrdfRRI3DBUeRTt3NPI2nYjvBigNuwqGN1a03dCEeaYf9A6N3IC62vkU9Rp
SeLEg9PAGuK4v0I8b/vn4/A7CIWUM1d4Ky8M+BRTNkQbu9+nxjn0cVtYpze+88GU
WzJLLpaTrIIN/xFzZHsEYk4IMvWE1AjmWuENNRJsXJdiMD2CegqRSg==
//pragma protect end_key_block
//pragma protect digest_block
vTzep7aPBrDyJaYAuc2dI3J+RjQ=
//pragma protect end_digest_block
//pragma protect data_block
S1p3nnKkl0LYZwl8r9V4ghfCAFFYVfW6EvrzOywcCgIIjhh5K9bywBXKDZi0yIiU
0efLjlDjpBT1KNb6YBAJlc+/a51jyqRzOysthCGyk5PNbbQ7DHttLyJQuqqZPCle
2cvXhZGsWMh3kVb85F6AJRdnLS/5n0+4UnUIhAK6ajcFZjkh6QSzC/CLj4huAuf6
A8lUHaUN/VyCfkpdU2PCE1Opym6tIFGgPOAKBI6dG14Og+hkaiko8HKvbYTIr8ku
NQz3yYUUH11yPiCruMLJ99xJLZAByBJDYf00Md3fS65yBBo0oAmlyvLM8E6SiLD4
dvEc+6x2forlmBEOiyscYbITqpQKPzbA2F98U/h/qqBrKafhldadgkqs6jEDEc/j
27zUsa1cBglaYf/HbTRjNYKLcGWULZ7MYRpXuCvTKe138AJe8ZK3sHbe6ax4whSL
aAvSxRqot/Aph5G7c3xiYSX7it7LO5mNBFxmiBNUkwcmQGUwp90+mm3FeIBdkDFL
3wMDel5zmTiHBytSbBWQ46sQfh2mGpw8vqXWtiEsZBF2s4r6zjbc2atP9ZQ75JXu
05hVXkI+iPsKKN2swoEA5eJLP6VIzYrleaJj+E7wtTd0x3vZDioU2hKgVfA5K8UC
VnAK3ZaPL1dmfQWk0lqzTfha4iw3J3F9RBCifcyXq+9ySJvpw7xcanXsLYKZxE4c
b7WQ3y8FVfQYx8qTF5tENZGpMP5KfwXE85RYcGDERJUK7VykL9f32HQxtroN16r2
67yg/D0aM0ERm2AvALGR1B4AstC9cQ3eNmGcWF6AJN3Y2YZ3bZPGvRiIYgTCONyp
2jkvtb9fz75DpAMhI8Xj1X5clSEKHKHgyCn/wE4CoT/1gv+BY3JR0AQ4CSg4CBT/
IxB81608UJrKBwWSxbIm3n0RLPBYsHKtl6wFUmwIR+6sN29GVseah1WfgdFtG4Sd
HAbBnPNKB7ObHX0euIBVZGbrj7RNhrhSozW34MZaKni0MBzbBTCV3yhzlEQWsCB2
L4mFR3pvD/ymofISsZjzzxv1KjS0ZNd46YLNSJU7ukWl3SzKPrALO1WmV2Bw12P0
5o+B80gs7a0iHF1ECS7I3KHAINUmXuZvf/fjTBt54V1HmAm+EFtsGu+GX67huM0G
36bVT1qgn3fHLGsXl99FfnpLDuCx5Ql4qQ5eG3g9tCsEllN5xrMricBM85K3rVuX
iVEXRU7ls39v2JDhRMVq8GPjv8BlZfknQjZM3GRAo9vHDV7fVLGhQKhs0ANht6HK
KMyiY36yTgK/wLuUyOItSh7W22YJgNGfnBtbQApbvozqCE47l1+hTo7wl/Z2cEzD
TQhzqyXirWKF9/gWU8hzHjA40hmyaQ+GkVt5vyMAANqG70//cqbARifJf8LFTT2U
zs4WPrIWECAqW8sbP8E3jF7zQ12X/hPRnlIkUyk7VOcnuEOBVH9K4UcQ1Jq3qesi
CeUUxiqb3kYQLkljx+X6aCDdAKjFjx+Bw5fDussv9Wo1U4QXJ0dHnZD22pKM6a4p
3n6GA2LwTVv1cO6bAPL8qPhx1CNldZkd1aN0mEsxJBlCagiFOVoit93pZjsMkhF1
P9wS4U8FiIrXjhKHyAahhWVhexAL0iinkfpAVhivYQR713WTbaXilYiKwKL4wo4P
UwBvhcR7NtSkH7mukzSzI6EZiLfBTH8gM3kKyYyJmm/1Vxv6udNpf1+m8Ygrv9+9
5gti0zXwwgOzKrKmJsohdsaZPCfghHbJSAqPddHL6rnk0CLK1qCAp4/qcqQBVoB1
e/7HkBQPDvjGrqe/FjILGqJasYrY6h4FkGykODTaM9m17B8sBzFi9xQUUE7DXs2/
w4uGwIxZSOPqG31QcXFUdb9GDoLO65A57jmqvQuFFxF5IAtY8JJ+GgeVIoKQcsqV
ipkKwBqI8rluysy3jli6n5ckCW6GZdqU5oXlesxFbiuQk6EYk3728absZqjkMlNE
qcQSuUg3z4ax5V36L2J5xPWgXeoLU1z8ePxGD7l+A4i7jMza2SQInSc2zk9av8G1
vsmlQZ2Tw9R0Wp7X6PE768iRogRfpSes2leiHaOS/UglmPFJgwgfSjJESt+o/Jzf
n2U//imPIPTE8M0y3X95wXLSfhvvEDxIzVOK2RkTrvMH1EZmib2HAE2ymgxD05QJ
IJ7Wp+D9NFSFRMGWxvLLDOeqMiyG2LJCjUVlR3nhpZI685lkXdl4DZylBKP1ihbb
tErzAfn2wl9bEjo5D0yGpvAtJUzhfGuIKHXQ3tezsO2Pu+SCLZBVsx3ulbR1/kb7
ZZC9V/yT0/TFYSFk89FOspqJhv/Kaqyo6Mr716hMvC1bLhGrAzeSW5d8yTq7P7T3
CR6zfLRli6eXaxrn8yiWM4vvuAfIVk/nF+AJmiT3U+sYHVocVQNsNwEhPb6RWgeh
gqfFdj0MGgBXW//lyNla9ksgMFBY94dE/MRiFo931kzoaQW6AaDfWjaO02FCrcoq
8NsiJ4tPXghUspHCAQmAMafz/01wybXbEZ+LAVuoZpNNOrvuhGe2nApd0yWOtDQl
Pkk9P2BLH9Xw+XRRDd4xQjgGPkmjBJeJWdIC/wZtDcUA69UfI8X4thqLwgIY6Ncv
OMQuwjyTGKS4GZuogXmCVVR1PgwaZv3t3wyq+Tbts+0M6JmB0n9xA5qwOfDsqbyu
acXlLjbJ440HkkkvIhVSD3hjAL7+84wPfF7YWVl+37otm1odQvZmzOQ81vcL13fF
zn9Tg4gaXKlqIp4DwIAP6aNvGDgIGGmZZH2dKt4DWQsZaF7F9eDs3I3w1j0myptC
L/a+lHsIJ+Mmkk40DaiKS9Br86h+I30qqTYC8oVtqdQnThHWV5dCxHWj0NxV1G4p
Y1D0p2dMydzdQL/B2Oldu1hTR5hBmqAN+DchQIbGLRYPZ3/Y4iqoVZCIr+itPSNW
W48s+7mRkQlm9Ya7gpbeu2L0RzcrXJfAXswdMS54ibfvj2m1NLE0zu8xPpdd97kj
VFvUHvwl2EEsXzt286cJmsFKl6UpJZhLjlHmmFyd3FuQYD+CNGFk5drUO8BdZlqJ
CqMCdyaQo7bVZb/hfGUs50SoZ0cvTTCBwz/Fm+JCJcesmBjZ7vwE+jLJcrXQLQ/8
ll0Io85g3ifBXM1x6jAorM77+E4mMAfKXYgpG1OCZiCW7rS1TfP16Fmuc3sIr4LE
pMoMYFkMzGf4vs/agxAxuvA7IXOJSuDfxcIg7BS/VNoLZIq6n5fe6s1vYq/5CPSa
MIqd2oWWd4PV1IuGyfIupmWADoo+7qPBa4DonwQ5vgb3d7a4sOGCSEaPKxSUxHiq
CyvLgl6Nu8PYgn/VcKFqKG0EPuEVptN0Yr0jdDcMu0hebnxBqHG9nBbKx70RgAGw
hd4xFuE7R0crVwInry8inG9QpPgDiYUOSL1Oy+BflyfDQRs+rZICmbkx5BYpRlT1
h8UGm8+hgGVc066XqphEEganPIe8lGLHCubmRFRaVq4cLvstexFR2aMJGgN9lXVP
4//Mj0kEIL8HUiqrWhpQ81UAlSMXzwm9YpwPF0YCdSBplLcYa4UAiUOoKLaVCJz0
5q9DjjvZ7hauGt6swwTHjjG1nZBlZAvHFD8g9eTjFmP5K1mjxsUb9efx6O9w0EJw
H9mNzVKmx0emFMa/8HHvWwbJJt82hpl9P9qtWYgfifBswCfMXLbshPTVhteeJhYX
mmisoZRMzWvTOwcXW1EXq8AqmBFokwjXtDmjdtXSg/PjjIEo7BUErJg/564Evpsk
2sSgJiMa9MJJN7z3ngX9Bj9ZAlcm3l4taRPmfjUu90pSJ6VRANJaNKLmjloVRrM4
VYxnfvpUcvTOLL6bS3eGOZAXM5Iy6zbhnjLrVxl+ghgyPRqf6aROEJkmgaarWgOJ
IAtq+lsYODV0sB9FysiZPf8qT0xphiEXQvC0v214gPH5fYRxlXCavkH7QgnR9xQj
ZckGzdY7LZF3vVUuZ03/BpUHMG/UdAy01uaVCzhSMggwTlnZxgHJ0AaPZJcRB2tP
jFD7BMzuStP6g7z90aEOQZYhAsS7Q5kN37/WD56UVNQP57IyojAJhFxks9VRxiqI
Nwb2KvZB16bPa67mbw/2XY+ClTST+jQfv7y5z5/ONP1VWQGhU7LUSvjNQVJTMCTf
mdtgTGm/hniQ2OJstI1s+rKjvOujBCPUdYulSBZWqRwpfkApW45b3YruP1nCDHRg
fT0a7eN4IpeL1TKFgerT5LQwFRZpyH++EOU0menrNLKcVToYYEyoWK07GdsxLoFH
CREiZKgacKH1lG6mBKK3Buzl+480XgsbJDCgmSvP3w4aqqj3pJyc9sYSNukREgrD
4kbg1oruenLvZ3hnsgQRisHvMo7NtgjR2fASmL6wDJE8HQqcIBSd/uboBkbdT0Ah
6AWbTcFfgZxC1DzJVVTtyUKW4ITuIZiQDCPohiRLEOWMyRu16n58CWj3PC0Aj7s+
4s8RcMnXcmENF5uS5Ze1qrUn4ajxXurUMA2d/91IQQ2i9UzNGOg4PDjr9hC6h2P0
TioHkOOjKkm6gqAVg9NPiPmfzyuj+l5ls6TLFNMM7M6PoB9kusNDfbhclgKJHgVk
5G9Afj54SXKBlBq1fHGr7ZhtRhNOvkbN02yy8p3bEGXlA9WKBKRMq2q1v/F1zwWa
H8h7/731ZJ9KT/hU9aZfESg0PPKhs5/8PCBd1YzVzId0XxSrHC2u77Uu84fWuomn
y5b1hfOKwrcSR+puZ6CrhlibmqqvkW+0U4TpAtN4OMWBXTyH1gBsYBBvUj4YtziB
FYOfhllloY0Zb6j/pFPn5m9i4q9hCWz5lngKfrwr8HuMLCszwfLPLmlh1bS9jKn2
Z9ZXYAJZ6MjtDgmbvD+y2SHxjZNDEf5KdxXc+1VnzqSi1pzG91LFw8jXxapyVkY7
X4P4inF2Isd5jnjPCSYwLjxpV9zvi9QvXHvAU7ssAnCdBibw5vZsph13v2YdxcSG
HSJC82RJY9oJe4YAWu8V7474TywLEJkCXrWs288pNDzn/DtKf2OHfs8V0pv2iMZO
IDXwgu4SGhwceB7QEIZU8w00kmqBmYmvXCypfPkn9jljPv+t+aSQy1Qczd27X57P
wFAlQZMwm83xI0mmo2kuGlrCNfcVi8z4pToglsedvK09bHEEN04xpPL4Sb4WBD8i
wEI4uzQGYx4T9tlCNTwoNPROQS2gmBPz882k1BrJn8rmzkyO+UXoMRvXipmkl8kc
qp2TsAbjplMSlF3gFNHwvs91+33jb5ShZJn0zvxzItXsNaDGYp+twKIou9atbt/G
a95zQ9n0VMrkaTiRiVglsZjnEVbjZxdjeaDkkAcuKoUhjgvJYC2XVMKceHShAtv4
bA6oWa2UlTZw3txPGaDcRb1zyMUfr6MZxW3zJxHLupg4LzDI1uMI06hYHhNU6Jfw
sSc0ormgDFRZ2/hQC9+MrycVTk+yAJz/SUskRfElKAoSOh0M6/6nO0rKTe3mLGgd
xSathHc5wU58Ksyjm7fVyL45PBpyyiT306Hw5MEmnvbVd04F3H1FqbqILGiTWDzN
cKwil9mGt0Rxqtz8dhpda+/mfP+0zVGGDB45fEBoKAn727UBFkZJFXARqHab4JpP
9xUb85yDCUXO49fhKNjX1o8xIR0SXULkCqLLzC2yhbxcNHDDquD+GMgpEOpes2b4
bpcqmJJHnIDecQOmK35oHkTeUDdhLaRGI6RFDS9Cgi9Wuho+OIYdFdcVsXtqBm5c
iT0lRAEBixbFTHB4NmBbGiOHhjP/3lL/5ucC8FVVC78lzzD9BLUm/SB9U3Nssgzm
+dN53Ix8nYxpcC9HJghzKL8q+Fc4wFK798H5J3FiXcT2ZKQlUtNr5Dhs2+2HV7Pz
qITwnJhMEr3ZknVFh6QJTpds4+osI5MTG3kR10tw+y0X6QHergcJSjvFQ4pSaAA/
C+GPluEWhFVAo7EszkUOTrqSW760+2f03mcshAvApSieEk7pgApkm5hiUsXXe4/+
3eoWQjyvCfmFsmuidzojP41n2tck3Y+XXWVLaXG8ROOKSyqbshPoOj2poy+eCYmc
9Y0+PJ/IYciEkJIPKjDBaR2JOjBqp+cUl9eJQ+Orf+I+1PcJKZBZ1CNWFHI3iAPh
1t/CyHyLEMyDrZqRgcEuY+2NDMyvNpbhcyivQxQ5keWFcQUMXS3EzjiemOJo9N1J
C7T44vtK7DRmByhMwqsTPqA6cRXZaUyKL9ew3lwNuXbAoSjVwlCbtHy1SLJeDJxS
l8UWDZDl5lPSOUjlwekpENFSmKLSjQm1UsMdNqA2gBOzdYVVgV3A2BeOCr2kk6mY
incROG+z8YyjBFsb61TYVl14jzxJ0sjmfTylb0naGXniXck4s5lqtJzjN6XhSkxK
+ZEBfKAeokOdzrrq+8IUyObc7SaGTJzb8AN8wRHbcSH2ZbshALokPenC29zI+0Yx
ZTNdTiKUQkv3VN/ZA0TpGqMcEJWBz4l/nsYiqUJDwXer6irWVcqZifLgW5flRlww
iWHT4I9qInGKjko+Lp7oUD+1JkmUqhpqQ1P7nB825aT+Pl1V1a5xJcZ80cbGUP61
JzGvK1j8o/eBmYGwQ9CZjw6UErqGLgwQHzeyiXqAq2likeLMAJbVTT7PGd9l3usM
w/XoQrRshh7Xe8nw8OrHf+xnfOdHhY4soiuTgIzsa35TpVSVIDlSAxT8GmGZmmwE
JDwABzbtdpZdmhq29jYOCDkEak3WszTD2GGpYGS7LtNsQ+Bco681ZKuOw7+wa+2Z
30rtjGLUtOO2Cskg0+/baNblrcMVuFpiVESEWkW4yni47Y8GicP1nJxYAg0/cRVp
hHfS43Vmlp5VUYMdk4dDuf6g6AMYat/BZclSpgGhjSC0A3nFEj0WgtanFD9nfjZH
23IeGNRg9J+cD+c1nQ592FLvw/YnaP6Y/V2lWmMms0hO6V2N0pZwW9DrhNlZHSwV
wjpNulFgOQYsJRTejKrkpidpx9SojGhkwf1+el6+cRbiIveeUM3aKT3xf09h4z34
uLGB26pqMw9rmvllJNXubJMmnLzY7dbU6BUYlGNqfyVnktFlsU817NAao+GSJ0eI
yVt2M/1FLDz9UUR4JMzEUIvk80zUf0KGqZURPaYygSYC9+dfEEcSbiJq2PgT+och
TubeAqjNGdePRcZuM1HbF9/Sp3bSxWBLIFZS2/9WeyU+dX4+q2evwb+WpvJqDaXR
+6zpCtU7FANUtYFXRS2ulyR15tyhfKzUBW0Ylrp4jp2XrVECb69HYszttaqDYPSl
NIkfN8JIrSymRwXxdDdLOjk9v+HeUGkCeISKzttpEwExfsot7a5rGABi2hAs1o1K
kEUS0SxCGow46xN1TWKUA+oubR+KJbS/2vIMVmZQB7NMYCtHzpy7k+z6QvHnDYi5
0nGzSWM+4REZcD1wqphzo5C5rD0Y9n6cNJ6iPdsYAu8QCnTvQKoP6ehJnZ2mpnmy
l29ZLCTky0IcgsaXEhdICWRKuJPAwRZbXaSFQGuoaFBLJMikjAJ85JMSSFtPjHnO
RaA+helkT4QYlKq+jV0WP7+56u0ofNmX17ACt21ocZQd/PTv7Em1QNAFyQFsaxYL
mvHIKrCZHh+dkjkCjYxAdKmO0iIBM3dv5OX6828qwNwmFKNRtP5cwtPT7CD2B0fR
k8xFeYhfd7thFNNhc7erME5dghtXID2EzlBawmB2Y3ZUmZklgIP5xfBoxU3OZe3l
IAMiRa/VvEvm8lOcyqD/mgApCpbRDh2pIUIPS3UTpNjl75LV2JawpEA2jNqDpfZp
jLZgCTHLiDksQmChQZ2OlutPJPzh79VuYPy5+vZ4nyychioD25jR/qQOasIcYf52
cCqUCXq95L7hy2gGNUqwKacpj1oAB3jl8GPgw36KXoeND4XMyA2ijGdZ0pPDoikX
kCkeoGimHaTL20ouIGHEao/GfXgxQBUnlujDbQ48MVMe9DN4ouDy8KAZEWanVoxu
cVd8K5bv0e/L0EcHyOu3qGqfugtg3jQETyTlpcniWZPkR9693OZAUZQmxoZoa26E
+uzNjUN1l37LRyiw+uT6tMblBuyEoGQwn61bUwm509gavviEIaA6jcM5ISMQ+xUO
o7pK3pcJr+krEz8qLZYDS8/EWBlwB1YKq12+W6fR9QJKOfxLQSwzLTUu0Fel9g8x
ysuh1sPAPwaMJ6F0zOX9EbUAx58N/9yZjOJDecB1W8eLwwc2K4GLz5rldkN8K5Xy
keiWXW6r9HUxrS9sWgWPb4EnLckt9T6NYk6nbAzTdhmu401Yq0bG9dvyE4zVSKyL
OpmnUPakthWNHgAV6V0VcPKlcxNasXf60/KqTkQxE6gQEXRZ8nI/CftFdmlLQsts
ANIqaMfoEzxaTA17awgdTutcJxcjs9FVdS6eZunOCltBzpiMYM11nkxe0z1Trbiy
5QFbhCSjN6APwcjHhe55WhzMxdhT7M17B8cc6tSMAmvU7bqjnsW4YwEzhlGlJSmH
bc+Nh+pm42fSYyPHfhFkqdwTuYyOvpWwdtFt+bwRyUvs5skp+7d6dJnVt+7Mciuj
Y6IW7sWHdAoCaFaglsDe6uWcTGHfhAQ70pzz7KliSJeTbHnO06eAhmsgJ4HOQqV2
7nJUdicbD1pSbXqLZyZWw58lvlGCfEjsHW0Swpg/nRNpwstzQekJfQUvb4VgAZAk
0Lhzl/3s0zE+hnyhu0+RNnymx6V1RkVY3HeKbSykjPRn3+PFLHkg+f2gZaJDNJEm
SaqBW6MeKyT5FznkkvC3jvdyKvd8Cag7XdkEgSnaGcRJ81OsMW6rrlMvcZl8ziuz
LaThEvAwejtYYEYF2vpWGKfQrmlsulNJXOXCIlheMx0fQVVK6NLs8aHaIvqQWsbr
45oBM8LKAWRLWPRet4NFBMsalS+3Gz3GqdOezO2btcSJZdgVTLcKdcqiPPq8S5nW
1csnI3MefPL9FzTWaPVDHyTN/KRW9Z0/dLC6zGD7QrwbBINDEu4SsXsYe76lKz6H
afLyEG2PRQprEn4Ya+6kma7JR/m6SF2UbVUKhQIWR1WmPlvTaMzRC2GH673JYoMd
beURBZM+ybFHvZDYiAm1LEGQUnED95OnqTwwW+yUXqMQewMIyiKrpYiCwdEx6My3
SlGrN376Va3NNoF6C/Qn7pY4/UJbTWRdbDSp/vehcFA8t6N7c8+V7ZGPw5XiwEup
eW8BvUgUtYkkk/YbUIcsuDZvLkkALqWmKacIRuBNaCriQnbhutgpO1KmTAxtZJhL
u5AQVHRLKWNZ7IKwtV2JaXxYKc44bblS/Tbswh8Mz/CUBEM7RkTiasOE5YU1vC1W
2nDSD3DBlH8XBLJrY3qgXEkYUQXdhtai2l7AbiTpbLcbX49p75qswko+/r7foUcL
46epvUcfJWV5ZFnjDdYcmFpqI/GVMcLrghCcAYbg2ZXUoR+316chD0t3dCryjPmL
GX03SheDUNSQjstAQBtZGPYuHhAOGWqb99HtxROpeg4ZL0YCqFMjG0kewyIq9qDA
aqNcs0BbHENInT0HY1gioS/ODSu5Z/42dTNnWC62UeH64CMCVnhcg2evNGiEtWH2
rNf/OFFjst+Ubq8yHT2IRMbXRC4hZ1HluprBRCvpQXalGX6eASh/VtTY/KSXC/Im
db1fcWehrjWlnrciiSgwQ6FZG3qGUodyUljexVRz+eapx+YHhO8Su7W0xrnKApYz
rTWhs+S3N5TTigfHtYtLT0AtWIOZnnlv6IPoRtcsaa3ZN/WEH9ZAzk4XkfoXa+Uq
S/aCCum+61oPKXEjqAS9cMpjHT0bDjUi5c7D6suUHVFmhio4Cybyh0MFwSecioNK
BQ1Ch79M7Q0CsMlgW5qT1+UWuNkb+vnTdDlPlLOyMmvdvpi83/LqNVVFw4YfNHWp
KJgN1jlL8tZ59GJxZ+vEzCsdyp7NRAWu0ckfbst6HIyR7JXu9Ccf6oUPH0HkGpCs
mBvufqDf5EWYOwJLwcjsP89B6ei4ADUZxIeTPa+DCtif4BK78oxmUJmaw4K4Bagt
6PpfKw4Po/XnhnM7AwoJJYFx16t6nMkQ62knIC1eRKlZs3fW3ZrDGROzPmnW3cve
W41f1pSgdvGVgALs2u2LG+F1/HoVrrF0eN859W863dh3xAqvygDKb97+NolNDuGw
e/gUAjLp3lDL5c01OA35fYlkoDbun4W1B5Ht6lESfSxyXhd5TNMGf7l1NzZpBVac
7+/RrFnLm4zZZq/t/n2wRkebH+hMwVd4QyN7cxxa4bUI4lSMts1KK+eJ26doafJK
SASVAxaELmc7jBhTTT/ZZCxYFlG7K8HdtUkCKCCSnOjkfN05KbFyQ53gDb5xNS/W
795JgQYg0TFzfo9Z2w6Tw9Hp/5ha8uB5ZrFi2wboRKLKmqm3nmbqXIh9UjfuM1nl
gPtVExR/Fu4kVWqiS0oD0KqjCkcPdIrkExAoVAtfnxZAGmVDvJJW1tOHarwRPx8h
x6fCNtlUFoPzKd8b1Ft1NR7agSkIz8GX5k8CW+wAE4FFGzg7+A9jnih7v8JaBfAd
1ewGrLNFOXDCyCJuf9y+BKWgV7IhCdYCTViMBvQvqs+nLuOB/nB33BylK8TUFwgo
YJaDn2fT1wImM759YifUz+PjQynH16y2VtxGPIoI/by2ATEjUif1ZEq59lEx+TBD
Pp4ChlEmRur2FSTVdzVTn629yU/P9h9BqS0lbSKhEut4BcD19AxTJW+aRm7KGgBM
NCN2AEuD2+YwFmBVu/EFyNdICWeT9khLkcEYIJPjmBXqysLRujTll9jPOs9mz3Xg
oQ8Eyn4BjsrfRZoBIwG3r9SAivEWnqBQ2cHOBPXyo78PXjBCj8/CRpTTpqh58iHq
nNSt3YYLJxHM9yiMEGes80OpBfero6jx9xej3BUBfu3vYUsN5GD4RZhcBl6fQYTH
8SDV2v71RuqWQkoMJrXMkmzspHzLocM4T6JhsXQ83cSbyhyXcFGcdcChTdRtw+yf
Dx+LrxbLondlC2ss3c2wGKcdyKXEpFcW6UOz7YoKr5l4/Ydc1NLe0CHuh6DDwSO+
pU3XmXLg/Y5iH/kAG2VyGTFlEY/+Vn6toGdxUjsT89Yla+s8EUE+7cajtfxaSTGw
10B+vC8JwTVmnV5wEowuWpVVKsyyExDsaf5PNBxOdPDYKOSyM+t7nVSNJqocZj4j
Dm81gjMTrLeL0DB8++lohMRV5RhN/vyOYiWUbnToWs1xuNvGJMxMvkaK62G9dzPz
xiJMNVg/7KueNewGnNb1qypZAEmrd5rSWE56LZsmERyxW804nw1+FEv86OJF7JWN
WI0h7hjdq/m8raG1dDPSzggzZAvBKaat2P/hb2xsrjM5D/FD88p2BSJtQMj78tcQ
PfvPquWFaunvAO6LTWoI2sH1P5dyBgfBTI2AZGu2JVQ7yvrHUcQmPETjUXbF+/fG
WjyuYOjcHvKaT2DGGgD67xkb+IYrCfaNdd7L8FbXjddRFdlgD49bC7u7LT4ImXJd
iGX6g7sh1Tt57gnwORcjGz4YARnxUS/GEvZp0GpzA9uAkZoqyO8NcmRNbu4A+vSx
9hq20hRi2BtFt/W4Ssxw2cJF515iQ3beCxv+GHJ5W26O6/BXw6Mt7HF14bvxXaYW
eXMq8hWwn+KoM/eXCY5dqt4Bb5XJO1Byn26u0KkbVC07pmtC51LpqG383F2Kh9cF
uu9DjQtapp6dfqy6H0RuEH+awG+xwRRohF1GXm1rdFalipzgxK8q0Df7awHF0nVw
myE5YL+p2eDZsbO4hNpwSNX6GogUZUvxBgd9zidBLz0wriMTHC0Pe1yFLqg3mnMl
4lX1ZEGchoZmOWTJtiifeVQYqLbjUTOSv5YFpJsvnp7Lo+zAcZqrjbQYLb9vqChx
n8q9kGKlaaypKiH1FHoS2xpVcnWQ/ZDJ1SVbOmnV3pOG6wHaK3bss7W8a5XslMIM
7h9rT+/9RXmsXE/dca0dUadrDD+x3KOrEnQ4tvkr2cz5N8nqlyZu7SkvAdTqx7kn
RdEe849CrsBNXL/+OnEVgHIh21n+XoKGCwxY9hE6vtmI1xBxUbN5Luvv7QFzZTce
lm8XVWoRefuYEfDdQCn5c3gCHgLZtmezMoboLYg1S80mikQU1pwYrxGq3Hr+0jgn
CC5Ansrx3NWvwone7lef0F5Ml30WRU5g/qqnWddIVe9GbwL2uynqWvG4w6R/asIK
pE6+COJUFxm/FoowBfgS91ksBCQSFKO+rhHNjgHCOd/TLnGGyJ9KUc4ihWHa0mpc
p0KDardtA3Ba20AW9y0hkOtz1Fcsg8yJpvmL7Zj4tOr2EWxY5wO1OU893nwsSTd7
zZ8VoQupWmSgYTDHN+ERSGyLnqZKAabkTtJ7ggb5mE7kdkENEPRXPI9due4OBlOa
0mblzagmQpWVlF8TtsKF213MeH80zB+jXfnWhvcW4kJMT0YwCKbMxp0Tw0hT7Fb0
YWXl58HmTk44oACshZ5ttApwov98wuFWHnj7KNV+kCBHowrjOBGNzK1TDU5bBXT8
3qygQ5i9GxMrDC+A5zO6qOzU9UJBCL50+w+mS4vEKgGipQ7yhVoWEHDWWtyv4zXt
vkN7QGXsvrRi0Omf1tWQ4yJ76+yXcMT9z3fmeLsVmTyGhgGLSXxTN70M2BTG/ogl
vX3TkxuNNuf4k7PiAJhAepZl++26W7A/jMYFSbm2ecw5gcd236WPzqBFjbp85VrC
80fKhTf5f9CKL7XJ0FYaoS++Pn0KczTlZ86OSNxL4YZh0FpB+MruH6d9GX3LS6fo
GftFrJkyd8FQtqgBeGSCP5x17gs4IAh3VQapJYvPww0FWSfGfenn6LPdkYbI72aI
8F0EPWhoXqCryvHugOEzaSEebm8AV+11Tzf56Tqd5CJ6pbJjWyAWlMEItVoasZBY
7dlZlOOUuwtQO2nmbGbMp5SUNez30KV2TfyAs4vhXmjO2n7MQYgzE3a5WX+iFnWd
mxPGzUjgJ/aJv5zJPTr0fg0yOrckJVcfyVHXY/7dh/sIatZA7JW5zK3A/3/VPEby
wSzsflP/dQCbP+MrvwNVpFyNbpMdzjQXNpmJtSAJHXFKc67QwqwaVTtwjWoiywVm
5XUQHJN7WDRXnOM/CTAl1+zztxdMQeVVJwQzO3VhDP+qGnT2nJjT86vm9+a/aBeM
hloIFi2B1psExUeAuC9MWfyn1PgTXT76SD/s95yRXfdFDYrVsHPwRoSQ05Y8aR08
LpJQORpewuw+7wVpboaw34NNYceYFZVHN4VHBugLmlBC1G21cfpy4s+sv1c1vxzX
Ub6rYRZNl1HH8X9NXOx/bEUbEqI28mqUz8Epqo2tL+xX/q88pbboUR8Cm/z00XCl
0rkTdy8BEyLSnV/RaUuoiExx8ntKD7Nwj59Ojgock2dXT4UqOJJKtSUim4IpMAgj
qf2LXsYxRRfNHCOWxQsN+rXf4FQbs+DY0NE9rQAsxysPyuraMU5flBiCRii82Z7B
xcCX1b1fmJ02AWWpWAcqcVOb4dUwFBQwKgTfbQ2FhRGbrvZIrQaQsDjCP+CHaqyK
vIXC8A0+57p+FnTOPEIWrSkykEeyJK5ASMFlo+QDprm6BtylqjJWOjk4LabqM41f
HGpN8f1I6+tn9RYdznbdd2LdiMTmtZ9rTgRcsvEniZ9rEDrEOzHEphfuW2t0CF3a
gTN43kZjEqbymNxLizBQBELapq5tXHvYzs1dyF+3SIpjU3LIknG0+ym1BqkdyFLC
4+rYYBZu1JW93532Bikl5GR+vcPu9m3fsQwomXdOhhmMMhlKqMUB3ZOpfUiohgDD
EkVihrpn9I4AIzsAIDXE1XTFafXMNincHg1qBD2x2+LHV5aiiGR0krogWg3yzxwt
vrB4H7hp/JNWwTKnMQOydyEhKPlN3buvZeMQ9zNtPSxxU6qecVmu7+0mQY7l3ieE
JuegTppUCNFi5htw4wW8Yqmnwv2kGDIHeIbkxsifxiqUeuHvTnxDYFjNmVOIMMBI
LTznDkKnUIBDrXpIq/tq26Hr/V6UPFLMubaL7ThXWqKBz4n8WWzGvBA226EIR8m+
nED3c8kDMf0sWqxC78Ai4EfnWPMmc467JEroQhLW03okdJmAoOc9ymgiVdt5yMYT
TJPCU+PTBNjY8CY91k1fgcNhXW6//+OL1xI2qF1KGk3R/iPtXHyW+wayNoqEY5/m
zsTMuv0pLT5zF5/dSUkATygVXrP0htkO0l24qScqJwSw9hCqXpdGBx2nMW7ktVwX
do5kZxySfSt8aHY1w1QJfN/v9z3RJ6L8g+6T+CNagboJvRs+jA4TdV+GzlbQtnKF
/X1LtMw3ouQyM7nzYq+6rGTcOOpj1zOmlv2NZwZRzolXmSzaf++Vl80ZPz0qVk98
4tj/j69aHIo8kx3AGHiA6EXfP8ffDjmiNMqDqUTZ/hXLYieFJ7CerQ04A3Py1MAB
3fUBUEI77mAwW8TkatMCqTgcLhObBLFhUJw+QY5e4T2ti0sKd59bUrdkcL8dlVhW
jzbPDAIWJmpRF1u/xkK/Dls6dqbrfhWYglPBlpErpZ4fp/Ko2Vs8Mz5ijJNlf9ib
NhYo1b7nlZ3/0p5UcKB4MmlHrl7TTBkHKZMxObtrNTTPWEX3/3KEJ6MfXQfTKK4D
+OmVVLGqhuFQc4kuWYU2L34qm6Vh3616FKxf26nccZAGY9FN9/4UDAfhVpsgwiwT
ydwGn/b4RAq14bdN+NZxhp2BEkdwpbk3TwPNF0XPLjSR4mibCbMkR/NSGYraymYq
nSfQTVYY7rBQGnMbenTz/Wg5UG8u38riBaJHbf/ZFnk4erj82Uo1ZAs0htExgHcP
Y54H4FsnVDJVV6CSHoglW1rq4FHk6z3ROok8v4PBjDb5cmwbkpA4K9shlIBqbt/0
jLfjjt67QrsqksTR12f/6BptgsjPp6kdnImj1Bee2RgOKHd0XJrmdvEz0lRAEgSz
gcBpcd3cqdkuRXAXEsrRlD7KiVRlXzi/yaWuvvGeba3jSlOw/3/xI/95Ncch4B5K
jTSwAyIIKO7B9DGrUHwZQlT2TtoxgY7yVFBawCzdq49rf8/x7e9Le13X9JWBxDfP
0w1tRSjtCT9sGtpGX4fglLmgHVHLl3NVQTaX8nWEhp1/Ui0obpORfwK2Uoh/1OVP
J0V8z/L+50M+emngzwUrqWPpR1A0xhMxP54NfcmxR43teOggs2nr7F9kxx/XNZLT
dSghW2UbAYDIp96/C6fX5Div2ED2A9O+im2CRzeLxvcjEKIlvElROLpGqz7GhYpy
tTyKRLJKoJXMQiX+g/y7YAkc11QLseL657N/y1J1oYo=
//pragma protect end_data_block
//pragma protect digest_block
79rjDsJytL64pj/Srtdi1/667oE=
//pragma protect end_digest_block
//pragma protect end_protected
