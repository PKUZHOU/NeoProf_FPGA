// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
Cjcq0JeZEq4zS9CDVgHwvtmSlC15u3toJXau1k+GE5m7ocpanv0AOI7AfqESB6gJ
bO1WDSJtaYJkATMUrw0/eP+s7SDI8KKsT8CqPt95xujOP5QLT3kLaE9YSN5ahY2N
J0DTOdzPQwhwkpGBlBtOumLhF1y4dcmw36bmmTF4yRY=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 11120 )
`pragma protect data_block
c49CD5ciFL6dxFvylXCe+mj63JhXb7gTlhFm/Gf8pPPy9yjnXOFWtTmDqG68cidm
XDMFadqcmIpMMa80z+6K0lrPCU9sBalnPzDVxNzQ1r9KYpKwj5vCCcYxgQ2Z2p0L
XxEczT0KEtiAXtpHZIz9CdedbSyhl1xO3H3A/8L/XtY9IY9vOq9f/ylcUQTpz0Tw
zy47xQ93eNkcUY+8gSEp9NhSHlRo4ny4rWlhEZ+yXBuoxE0vmtq3meLonC2JvAph
MgbJMhdkj96dzQlQuse9qxekyz/E4WV2nZMR+qaeyNP8MUFoujKaZjtWn1et3s7h
Z0emlzjeNTZvjow/fZBbOQizVRoJzrfehH9T75MF+z1OI5dZzqwFvo5bj5IDlo2L
gcBttNawaaw7UPOXutkjx1YtdDT5QIyWfyW6gw2iMSdDHPCEVCLLX0qw4sP2WKS/
obcJmjX67P04DhgbTC0+y2ZNBCvEp+p3WFlOjmHH/kMtpN7O6xw0cs3NFWQ3gTFK
yf3MZqqpIp39gdkttQNSoc9Op0GNDZgSvJYD33g5KyS+0hDsd4lFcqi2nDfVOWKy
ciyTcynBYvoL4ovtZ3Mlwz9OKOWnJjr7UKmJRbBVHR6c5lBCUlpDXw9InxZ5Xy+v
F/GNsOQ/ommhJr+0fn7o9kPphRN6XkwNsIHEU2jycObUFwOl1I/BSiY66dnlyBw2
unqfvNRXGnKN9DrIZ0hNW0S782Zq2NfmjlmhB6P8hFlJffPSQ8WtLww+rBNDjiC4
yW1iG5y4N8KXXj2lt/0v8erxt46fVqYc2/72146bpIx6OeJVcBps56DyYbFQYTc2
wSY0QRwOTexN3afYXmgHbKc9c0NZIHuoSlR3Yzp981pmEN0olABkIG0OgWIzI00l
IMwbvnJ/I0fev3U2PIr8TtEI3d294aaoh/UubmHNExewGHBbP93fADEo+i/w4JXu
BYe9kvizGxck8IrPheVmesKWKMUYHhi9HBfPnK2yhspyCruw4F+naCBe9cgKddeM
WMK6sTB6nu6nUI9OrjAl+0EYFwoxFAFAAULMqcZ2Id9bEhfn/UEP34Z9JDe4tQUA
/cTBlyMy9HMoji6PoKntxBh4rmxtqtgtxZWesKAV4NRpdRxFGXiuxBBWc8BguCYH
TyGHRnvVKrOeabS/CeEPof/z+k3RBjZR7437+4XuzD0TGGStlz7C66IMNhX4klq8
9MBQiVTVnaVr1uKRmzjiW85FqA65JY+5P8FzpdWe7mjJN4XfKmcdyjn2BbgcCoD+
i8beeYwy3skQUwGZoBHCYS6vGfMmYj3Yjy+RvvOSroRVd8FosEcAjyVqfpm+woVl
E0CJABDedV1XXxH5kRnuTrssdPOngeUXrhEpFyaB22yminmSOIwWrB+0fqXlgQhY
iX1tYL39GGmd4LeB5NxLBSuUFdN2XzrWKefK6jVO+9iTtC72lSl2jpnenyYmAgzn
8F0I9nguuMTNw3AMWkNGX9luWQNn4/qf4fS5aZxLYk2e7KswvJkDt3kalPMEoXVY
RXumkFCzNHyqRtXiYRkKvw9WOoE0vtkLMN/Xupr1XeLUVo+rizPisUeWnyG8do9P
Fvp1zlbbpiqu+asiqpfuV23h+EHW9JFvBpG8fKi459ghkwV8sukhsYB3JiCIxidG
vgvwsDWnwx42dq0TmUl2XH+4+FwcQGsat8uPqwCLm5x3HWDM3MxU89ZD2gsH+4mG
cbz+HKhzG7ApzgRr3KRfb5Ot0oJzP60SGyPtP/ZplBLTiPVT3lxLMXYqCNKqe9ZU
Qv8vrPfrCvjeJYXTgffaxt8Prg017+aXfcpaSvwzBwvjOigP2It3ce9KUzVoxDaC
ntux8wJ1IRJKtrgDu4HEDJf9sM3NuF5rKYUg4Km0/IPBvab4rI4Q2q7lmjiIUeia
GETX1rnZVneZrcWPW+2sAoK0KkqhlUmwNV2S/hXXzd5WIIVHy/yn45gpb8GUwQWo
GHzhA78wr1rPFczvLec58esIGs4Ufjo3+36cprLjtqCFbbeDaUDIqA4OMttAwE6k
xeJvAzIAiMWC6LD24vD/Pb3wLZZIWYTLgeltVhtkbgVrh5+vvxLhDOvc12uc23xK
FaUkLPceXDgJqCfloOgOXdCKSc3rrZff7pMtXm6te0MyxXOW1wRA0BoegdJkzdX4
BvGQc8qaS6N0t0nl6Fg364AKoIrfa8fN9tJ+eyrEleDypigO23j4g/NRUCPF2Eun
QGhxTnm+Z7wZdZLYO7KVLT7vcMgTWV4ZoFzPUJYmRN3RVRIMkB2ROsUHkNf3794U
ObexPQmJq23b/o/nqWTMFbeuX1vhhW/Y36pj3ahZhfiGCHkcRDy0W97k259fDyx3
mq4bii8fmABxPxlz6eQ7xF39HyxbMZunGweYFZnGukyRTiZfV1V7mbUD5ZX132Jt
z6dz/ujcxM1AawEWIrK/HoxrlnWlGyykwgVpWGENU81jALy/6LDIZSEsuvVIuJDE
jb5x7WJIOIX+5SlkqOoPsf1IXO5I3xu1vM/WDkV5+i3Tr0rBnIRAY4zpeROUKChq
zODX6J8snaN/XlXYw7AypUntAbyD1YfN1ZlzYjoCxU7Cz1SDbmXsDGKeAIAy464O
0Q15g+4oOaWNiio4HNBB64+y88iNX2nZt38LhBXgpSS072kPdSzKat1+zxmTA5qx
B46pRjcjbWHcaU5DZL2EMeOFK7mnthQDqFwPDLEMIExOttP3sYh4kx41Yul1Shu9
N++ZEwD6lhkzz3Iidq/8HRc9M4zT0uZo7GbnSfLGcF8ATurOXhBoOTFSmfhidlBh
7klcMO7CZ+VBTDKeywb36ynffiRmznk9UL1+6PcHSeoT0666jc6O0+HE291sMpuA
qDSgnpuPnqyg7JFJGJR4Lxw0IhkO3xTo7isAPshwCFm1Rsv5FxAxJkUJ73LQHwmV
vNacFTXSJ9UZhQY9J5apfTZry/rWvHpt4N9k1Szva/sg2hU3jr7kdC9OOLluS2v/
t/A06WYx9Hey/1AnjWwiJfzLwyUYrQQSUTlB8UrUVtl/UhbvZay1yxsIk6cT/C9I
eszPVYBTuDQncqrc6ZQrO9gz2QmEjpLEn5OK3Y4eO0kXp2SrYl/9s4gq4iNx60cj
TLva9crkUAXFAolciQvftbvBml0d33EXT2hujD0HaOHKfnXcSZSO0u8Caq7kWx2C
N6CxSKlZ0/E/5ftoJcOnS3ayZCBw53sSvjt5coo+f89dFx8qICaZyYd0ntlvma1A
Lwig3IyXvptUAJbK8APWqOTfb0f6bcYjAPIUd6Y/JiCBTEn+1pmZ5Ja0fx+xLi1o
E3u0RlZr64/txxjFq+hSgyGT2/bn0K31TgE0kWbOAeO19wwoqskz2YEJJj12HtHF
f2dWste7eI6C+42P4vB3l0SiwVsH0OVcmkTKJrRLANQsmMgaKcQzUgyHDuL4yZXO
KcjxovZGd3+MrRBOxuLkotxWJrLKG6Z0GsYAHGr2XFrJ+Z969hyJPpz9k87iJKo8
fNGMgcULXypiscIHySAwxFbdznvdTM5KFoxuxsl49XhDo8ByPxT+GWE3amG715ST
2Ghzn2rK5vTB17ZJb5sTNUtxYZCf6wJD9VDvIokPkhQUyQovnGw9UkVYqQw9saGA
k2k9n1F1Iqe3n9cYfDWkPDhw7cKWi+JKuY+cTZMiDjZLEQrsrpHSUoFP1neDx1Bd
UjXA7YNg4PA6ZgTO5y3c3AXU96AQDdIkRMFM5DMfus3ysNGl/vm08Wetbc7GNNyR
zYK8wJmv435LrYslsap72PuJso+LdFFOT6owv5HibB86dOCGUw6/y/SAED0z/X3i
HwJuSfcsnkgsuBSNZqWCj06oB1edHxfgu9Rqr0W77AUgyHJ8tVG+qSpBI5Y8n0tl
OrrUstmWWSmQPz621NAn/qbzORHE2k01WE65HmQDnAx6jbRHl+uOe5nRN2a9j2/r
odgQrwYkNP5bn4f2zgywzbZUAhgTgyUvKr4do9FdSAdNqHYxE3iTLCRabDDIXhHi
iPcryIXJvAMF2Y4H661YGE/PdW0DlDPL5hHxq8GaxDENUlgpKO6Kk1pDgvEXC4Sv
NFSMSxgG8KDMHzaJpO8yYlEfFJGbM98jPGodO3wgtmwDxjfd5AIhC5gpmkusua0M
CyQWnqu5BLxqMTvML6Sy8z9ydpwySSuQas0pRQD1xBZRMCuEdTRl2/VZColUUlVO
15ZCLxrzkoItQvsQ3raZkCCb1riwIDZOFdIAygKrsW4l62NAoaTwHAXAXHfQ/J4u
IOO4it8s+JX7YXVFUKrDJ+gp4wFqgnq0ArC4ug18PUmtWh+4EBzwZgBRSGBm8oE5
miC4B7iVj8MsgWjSfBuTKuBCMuiymMlHtJFyy7XF85bKHHbf5ba+xamU3poz4dah
mVnR0I9aOStaBDDwZAzbgE1vCb7OtMh5hYNfLpgsl2cnbfjhQqp8dCf1x+NCeGlk
KJ4XOsZA+mvGzLwXz4xf8hx1jt7xTAGzsl+s6TgwHViLIMluH/f8sYGnu10V0TiU
l7JsKiJnPVCk3nemPKsRwkdIMll1/8zSRsZ3gbQDWpWbW3jmOFarmuGsueeECyvU
NyToGRAs+YfWuCfAhUD62YpoVgQwgQgZQXwX9kmZq7B4ksQy4BtwQ7Ffv0nlgsX2
JySsWXSLkzxPVh3zvmocaPkPyezdsy+uimm2mq6Nwm3iSns/+sRpCFS8WmajEhwh
qRB/hASlu/mf6//WHGvwbiOYVGD42PQGJIVShVMunTiSEbaFd+bAmur2j7BYy7ay
RxNFyR3eYzjrxeXUfER0TzWs7LYN08KJxc9T1HjDD0IrfF0D/IeKeZ6zq3Hm7X7n
/vKfZg+Mw97hB4WU1CpvUxW0hPxQ0tOPvBh6gjLGs6RZIGSdeQnyuqOXPvGE/ZBw
dFCykigX8hq91AZIADN/OcW2Bc0/QwHjK1C39oVa8INL06ZECpyNkTkQZ6bbq44Y
S+tNRvbuRtajcR991nbWXUGqTzJyHcSQxQDLYtZz91txEh9Ox/gh5L4uATe3G1gW
2Jxd3Eom5F7uMgGfprN6FKCKuZdcBs2sdj+84sr4BnreW89SWhNXfUW8UZMzNAp2
nldcu8eZoL5zEgG+saFDjGFtxoK3dkyT/NhFZX0XvR3mi6dMDj+qm3BdVfsC9JwB
WezKmgGt9JCLXLuZkOW1WJdWoAFvlPTeJYzozMoyPm7H3+M3V1dw00uX4AolhKN6
ZCUL7RAHvkZlPYG0XbgiN04fE6DzCtp1j4HWIKd3cdmNdKGX8z7+7aQWcnvY1IxY
TU+bMWLZ9mWkQcUkH4GIw3WDXfj+WkORLcco+eQ0EBdZF/PMZZMjZaF9HL+3U4+3
VvHTfwntgOMMB51GQlT3Fn5mFXuVDDhHoILReTvFHPbsna8ZTFeiqPIvzlsDWg3M
jJLJLhDd4R5AF/guUWercaRLqKo++4ZB83V7t75hQozLS7eYtnLo9T/Dv4YHPXpW
2j1k6gK203ONVzgH82DZNgcyKkCMiIHdWWTuPIixyBmsiAI6pFHZmjjYuauLWiyf
EHj0mXrf7qpqXMjrqFQs+s2gffGXeC+3W/8NAWmO25WJs39QkH9DZGXsBIykZ9df
d4s02NeDh6cQKSzR54esV2w7WkE6w0cU9Agky1G6Cn7bp4N4CktCMH1BbSGwqpVj
abPFrCsqbINHzkN0S6l6oi9s6Jab+LYI4Ed+Wl37tyVNXMJ4rkxHigAYwtkmQVQh
Kt/NyDgrrvrubgq27CZOzHK0yowagI+FsilGwLzemOOHYekYHEmLH5Kopjd7YEWb
nJLvrpBtp/hZuhYzWoJ5gcXCyYft9KyuPrrublRREBuz3+zj7Oa831+8nbo2qCm9
0gkvLqUJ/QdUkbCalAKhwnAhbDC1Bg2m4p5CzCCIufp4Lfn8mO2Arbc1AY2QX5JP
JHbHeatCcvPnZm6BaSqi0dzPAF9k9lDD822UAlYq5X9FQAqMZrlWaRllSiHouD71
Gk/RPw8Ero7Xj+GymifLEDsjTZTFe/KS/zzCXK7y1UwCyXmxElBvoP2f4RwlCf1d
u/y8GweJ2BDhoT4s59hPBDwPeDioecfbrCA12Cp2nQSvK8uNJrmHCEKro8Ucq1H+
HhwofHA9rVlpjMcneFHsK7KuYPYXDuIGT80RhTN0UO+11YKUjracWOagPKyRiaLu
SCZIn2UZ/SSIPNMuuiLgEaXipJkYxRjyjyWNvTKwfK+BkAA23EzvoWBac+ndQjwF
yBnw9DRSCg7gvJVN4YtspgoSg78BVMNq7BYY93Wscmkad8iN+68ttkfLZV0+gPIF
RvQ7xahg1rMpSQIm0ohOpIdPL7f2XINSVUtV8M0Qs7KBRWKIsmOOldIasLDVKb5x
AycBbXE6oJ/13O+MR5Wy68vY7brAn8CfEzqGfv3CHKb9TvRBXhYOENJFS/1itYrd
odD2gry8Ii1SMMpEZSu5XAl6uVGUxfTuNm9n5si8MLn9jDhXiAeWhtnZi7GTZoxD
GuTjZ+HZNvosN31YMf2sEeUxvD/pwthgPhIn0JZNkEH3JA3jwWBdzHM1YbW7R5u7
IliuAQQMhC3MVLS1N7Mnii5+nWnbuEoGu3E8qgF8fXUjttYx2Fa0VeBWFIfAz69v
roux/v9CacyWrbfSRedHVqD+W48mOiIWjHxB0SqkpqIME0v9Zfvk06S/B1NZjlcn
ozkuYYR2avvvDqOcevI5DEvCr+wFP443EW1Q7n0DHWucPVtvOWdsS74PbQT6ob8q
DrV9GundQmhGdHznVZtncqOPrtSOFRLXjhT/jxwnWc5jK4aaBYH7H4REmUh7NwY8
IqFf758afqKQeV8uCmU9mm5IJI4gqeSLrbwIaAqBwEcWqTjEG8xjsTgygp1rJuwK
BI3zIAJhmt63GcCmjmYztiYcsklsgnIk313pyIqJf2v9O6xBGqS4FsJQQsTPmaXN
zKH2hnDbsyCWU07LD6V/x/VaWrS9BNfVJJxvKGBKhWn1KZnabngU+9o2EfwVBt+x
H9yyvzLctldjaUtSfL/9f53R7HK89zcqXr9/RMA/WEwzwBUciV8SkoY5bkWPReWr
5O9TNrco8WXZNM2048Y7jESR8ow/lsu6PDUa2nq+COiBgBlFDkTVXpMpYKY07VyD
2xlfO2COSC5fM4eiFLFL64E8EwwSly3K0dpKP1AlEkMeYaGDUDO9v04oLNo2+RVS
2zIpGQjvSdS1p0OQ86tB01ECmhQJM+QDSMUBujpLqCKk0qSqPxmvLidxtvp9P2Wj
VRc+TrA8p+V/iDtVKKsKxeRfDE4eeU6+sM9MGjaP8bkKK/LJohKxJzQIqU+DLwlD
EG2RGIKDNvzS4boTQ36wWH7ekGjZI0j05JYXKMqX6eRpImFW7pOfgwEmHufqZtty
v11UeRLbR7w0n+ikolIM3CfFEvvsCN5rNXYOFebpk0eodMWqYm+0lbCE8Qa2KvJs
M/MVNc/hl26tLBJpV7Yk0xM/Kxa7T8Vy3dXtj7im1CLH1O7hWdsDxSulSzCOGzvF
Zfj4/rr99yiawC2PnaE5FHKfWoQDAbj8AYiG1G/n5f2cJz+oDZsDTGFCkHF1HioD
ynek1fXeXLWt71cvLFJoxCxIM/Q7eBslSDwT49ue0XGJ23SHVgY3gaasTvRDUfqa
Vk6kU6dl0xl5BFKOiyPStHzydb9KYLuYjFKYJ0BkjTT8CoEegt/33ZaAlpJ52ud3
DejrFgNOOG11w1oSVNk1Lfe0S9h0Fp8LJIsKEvmZXsx3IhVVA7XGjuA/uWPxWKwk
W6iWKXfaAUK1GlcjAFYIOgXqirVem8BuAaSWs4oYSgCb4z4wKI6znsKOZkrYcIrE
s6wkcPHMd6cE+TxhVfSUEuis2FSgYp7otvkkpKY700O78IG1argG9h7vzhQycobY
heaSfcxczURqA6VqsJTUJX7ESq+ixBSAHsjmgH4ceSXLUc6xWJXe+bpivKRYCIzZ
AFZ5qwRwRMMWCb7qqUDErFmMJBHrBm/nLGCkPIs1tL+UlBPWwnGXO8JLjPjkDVRd
h4RF2MNPYYgo8o7xqhUVsH8CqsBGdg/Z8Prf4DjcDFQj4WT5bpFN9cEZaWq9p/NL
s9opQmdZWR9u1gDb50cUZhj+W2LZB4RG20iWQs3ArniuoUFQgVv99ykjIZlEaUZ+
5Z9u4RPZmpl85llNbaSowIhqnZAo2xTEZ83cRVZULin6GAmL0Rud+gRCX3+psKYs
nuB8GwjdfjjJTuJMxSoIUukIq66t9S+q+BbZs98NlxMkKOMIA72erpmx7PCOVCha
hHJCr0pCyjOdWCwHz5KLovsZchl4/I6O7Y4EV6vUSHAz3eT8mpQe5sS11fZxt6Ap
lJL/4X4jTqYxK57a+7h7BXkd7TJU5Im04kNz1hEHTxOFnuttc7o7KUON27NNZVK1
zdDiw5RA0l+8ptL2B1UhZlNW0MM155XHPlZpfbUb1GJsZM6kjkOq8Lv40Bdq7WrX
ni38TAflh1frMSpsgkPvnOaN2Qpc3G3pEYoeN7+rjmYceEmnUUVX9ucfqQ082www
KcKO6qJXJIdOnONE4BGcBA/hqhWlGtKmNeCH1RK7YRHS+IgKjZxNJm/rbyit5C5d
xQbXVCmrmbzlX3Iyqnuf5YDH9/EUj3RNpGr2sLkraE4akPwn0uacViuPKr0b2TEE
3L781maEIQoKiSQ6zMj/JfdUkyAW5OncGls6S2UXsXOBLbboxTTKx6pESZZvHXyH
E8aSkWHV3elzhVGEka3uwNbNLXntTK0pocY71ruDdAK3JaqzQUPP+IYw0c73CGfe
tHEdgH67OysTD79hFib8sfELu1WTOtDu1/2WoFzzTIyXDUT+yCVynzmzs8zzgSvF
GqK6elmPB8oWACgmpPalT1SdPXJDj5g0ttA9h0WUzQK61aDJhXGn5sJBf177l8+n
JGC2hLAr67Mbom+8tWDn3g4SAXarhN8gt80E8TlbpiMM2iQ4LWPsWI//zEfmGBzy
rkF1swhiJCKER2Olg0dBI1ppUFb30LChyTmW2Q2jh1bzP9lFLKzOSGU0YhRsb5oi
LRSnb5cQhgvcgQG7bJBUJLmy0zBpp2zBtnaaDd7q7WIEvVEdh7CieOHmz7nljrnY
LMJxTf8iuP47kV6qd3NHtOhMcwUAQRl06IoaatatxANvxGU+tISKDJodmmpHddkf
zAPgy5/+Ib5mhAdJt/QqzKSv4wJG2dLCewlzSMq1HLoLialQ2rEL3Oy9W20OCoKY
i+oLRI8tnKbTy0m2SkVggWQ8zVG+rZhOT20b3dpeqHaVEnkw8dhfvXe9/faogZfg
1OSXPLVgAaQfFcEMCeO8Lz1nDPioQzV1bUnQOg5Uk3JD3GJ4dzeUvl72Wrtbc2dK
dcrrfxoS/SBV4HBqJm7oHU0VHcJ5IzLWPedlF09VEFjyQXGMpo/L3KUrumerle3V
dhaQbUjMATkmx4y+FD9QWh2ZGRJ4bmCIwkWZXUOgzBwHcMc06Hg8BgwHdttZkWn4
vt9zX9lBzvqJyILYOht0XNzj3/7At64+fMt5BVn/ndofCNjTqcpiZUeJBza3xh9s
UvjNV/qxDbrq46QRXWTLvZxTX+mbbG3sQ+LTwxtOvv+BHcbejav0ywn66Ctyo3oY
uPhyqP9RzNeahzI5uyJku45EwFROQvpMZFLYtp4VJAZoatRLjZtuHQZ/+jKGc5lh
fbNtjCYJEVumpviv7c92oLN0wT3qxe4UKopV8BkGI+frKfqS5mCCTelwQMpDREIn
JmbXsi0LJZE1niTIN+uPHOxBUc8fUfjkMIb4Oqgrn/mWeOlXWLMCsZbgF3fUi47l
zvF34tWXXcqRFTMuZYe71rhVZz8t3aTXbYU/BF6lAjY2znYeGdXSGMv0JCOhmgst
s6wW4gkdT7Igv8QL59XWKNYNIxilidJ4GCcogBEODTMu3g1eyAqg7ieN+ta3gViW
IGiU5TrVKiUGSXFpaajic2VnX4i/+Wo/YXO8e13o5vBNY/WjPEW02ArcdQ2Q7BZg
3qdRgAzVjQIZERnVwmAijpE1FRMtXGsaS9bL8zpqygj9EXstaVifM+oB+VT0Bb2C
vyycyql3mMcj1FhwtFNwHzFgmfZLrGVi6eWIy8BiKvBuEQt7CzozY438gk8syDWC
XmRjrWLTU++qhIslQbRJfBQgW1pb1yPTEWcnEB0wScQsRNuU/MwUuWUNM4A2w6Hv
il58PKl9c0beIUGprnbsc1S3x0AWtlMBzsv4ARjsOWHi5zqShU6IbcY3Jm32yvTo
PrQCzRRKm+KiBfPTpQi/iwp4bqsoNEomHDFXjbKVoDpFEW3KD5DD+3Wm7aRDUOOD
fHl5VJqnCQR8ttIpbk42DKchht6Ih1jGInys/iOV+SWC5ioLLRpaGq+2/ZC6u4O9
o3AMKjECSaTsvMz9Debc/hg0inDBCCYkkNtXAaoJhMlXbpzGrb4K4Zx0Sc+1vOru
ZwpI0jKEdguQuAEcBs/3e5VgRhxKShryf/DO07fxRyDTF65dF/dMxYm5/IJl/HJG
3OkUWFVYT5GbXWbi+VHnqdpj3IDQ32R+eLEoJEogClf8CNuAb1EmSSoPx91bc2Gf
4rygK0pOm8aYdkD5ebXXCG0+SMp8LmmexAEkEylEIdX5//H2ZqGGccDpX4no64xB
gxKFnia45Xc7J5JRR0lKfgjj/l/NiLlgF9rt/bpSX+o2U65nAQtZsgUd8+afSH2u
XaLH9GYR/G5yQXXAWcdp4qWd1TW1hOlMo7oI0qEWzNbnz2dJUTmZsAsBej7AREJY
3zF3rg2DE4MD+32n1rZkfDSJc52GA/KJIly8dmSvu4+lXzNEMCdUIQc94Srbr7+R
mgDn2Nova1RwL98Y3bjW0LMEu4xJpiqt6CXe3lPE6fmUfqQW/+a6L8oTCmPvwuwW
++xC+UIABYO2b/7Zqh+aMt4FD6lszFNt1WOhBExnI+3IwuFepGdSoFthpkkgbEUC
/fqucJx2Z5PtEvGJDaNfXJ9PyPa7VqJjpfEmjOqwuLxtE2Rmuxly6Y9n8gJH3gmf
7EeDrzbVaLRkTKFYDOOuseEJV79wuiMdtpftctOBAqgw82GZx1p2F95Wzx9NV0DT
CmPhHXCy3kLIYiWi6B76j6tVMiODCIu6RRWO5gqVZAP3/IaMzSmg34R7sxUUuVXT
WnMjQ2BCnL1xOR6cvK+GxofVg7fN4K9/5MRhXMdgm7EZWpaJbGu3b98EJDy1765B
GwKTTgvxBo4h/ugnfw+HUtv6tr9DNTW4mWL3v/jEebVNiVW9MH92VRPnDEAwZ2PV
jbmh8AtR6CptsfmKpK8zBprEgSNLuA7r/gYIiUA2LWAnCXD6FNA9eKjOCWVIr9eQ
SrPfmkPBoTOjFEUA87JGHfZq0jHUSf10lBlISWZQTBstvH/bkAGnCqBRX0QjSLmO
CKhTNq5sarHv+7Kmd9nw1LB8pN5MUCdqLODrqSLpTdbXGhdRAwk/ZqTRIjcl0k1S
YMuZfPifGO00xDo1LqcPWcVo6yzOxsOO930u1jJK5BED+ay3vPKXXZ9v56D/gysS
I6k/dJBDszE7snJCyGINUjUIyO5NcuNK58LDVxoei+NjgREX/FtzIur/DokgWZzt
ilPCg9LKMtEy3ANGsCrqRM+kmZBhwFAd9QdUdq5OApINEccA9JqRav9+KVQCeePg
Kc/EBFOzzWLVsRilF8oCq9Bom+lpZH8Fs35dRCimrrrISVu2vx3T7Zywq1zYmKhH
iaSBUyrmPSn6nsjEeCtUFZQUExt7nWNfM2Zddjnv3Ia8oJfPK+G9TJ9PUqKflCla
v7jS5z9mr7V7h/JfZ0yChW6M9GhF0byzOjGp2a0/O+ZAmGIZvvDt4N18yR0f3CK5
uCQDzvZHeWNhaYued3kAuAGOZafilX5RzON8BjWRbRiawhu5e2hhiDkHLC7C3U1u
ulJN5+KRur030nnFoEtZ9gDQUXWtYMNg6KQ1x2Fg2oADVa5459MHZUCWSQIWxBCZ
NgN596obGtbb9VO76iF6pP7rhu79L97kZVhA12HwVhZ9GBPcLeTTqaet/xYOv3wA
Cd2VzthpJQ2feDj8kvfhEbUisk5FTAkB+C27h751KsX46ZO7w573OGQDXTM3NI/i
CuUHprWb+oKxOWtg/jIYVnsAKoNd5exu+vNN0RTUL3rmuu78e/1kDwXOE6IxjtBG
8N6mfNrmaXioX69ruLbFXEvd4b0N6DtzNz0yezh8wPyOTMmmW0Ypoxrf6RlC9jed
mbcvsdvDRvEtnQNOlQkMkZViP7dxL453yUnuDIriEObqTWocVkx5Vyexawzf3Y2T
TzJPX5zsuZcXJbo4+813FG5nT0oMqJvKNIdiei8sQhtEWRMxgZ0UjDskMvJNKDAU
96CG2uYRhx4l0UQBlCl84YIuhB4+S+xoJkyOTallPfa4KgxDu+L2X/f48GX9W4g4
MnqCjx2AlVKMOW25YALtVbDlBYkFvcgE/aaC055xfks/eFeTFzO2VBKk8rvh+Gui
EhCwK0wO1QZqED+uvKj1NebrxCLRWRdLlS4sgMQ761/uy1cH5HN+k1z4VBX3BNDg
ANnOEDi5ZT6wte6956x22eYtQDmble4SE1TdV3L/Pyv5R8x5IonIBa0zImy7pXTp
pWujyOgnZOwpRAiHLTykatVpcVfLeNxfp4cvpXNnEw6V99JUJ+bH6nOhGQGOHHui
kqCBuuz4uo5LxdU5wbeG9loRZmxzRKVenZIUzRkG9jYtI/GH/BQmBypj1yL4StR5
0j/CYewQCOevo+5HZVi/yRXbSonbvTDMQTAROYKJc0xgS8kL3YFJYxWALKyV8feN
YsHQnxRQV6WD80Y7lUQ8agnAkOGyQlA526kSn7Nb6E0ux3JSkCAEYJB87xsZRk8N
GVHLp0PNWuvC/blwZS8hUBmWKE07wT3HWA/6aLahnIcZH82otwPtVqnTcfApO1/Z
tk0WxNVv920/0AUmEmthAK+WegQdSXdWYQ8aY/RoBDYtyxa7qCrSNkVcK/2ezeaR
a6NxYlekaJzPH7rBovQ/rM7o9ErZEA9z6pNJPmIuSago3MhGwDzbnGxXV/x5u+Zq
ip15w++YZTh8/lLJvmDqLZklLn0LkGc4PfeGwvBdSgMrdyCnMM8voQtgkNkVCeP4
lPfB+4DB5GPJlMyPq4kvMURWb9d1jl25Kvlsi6OGq3qYLEp6mFSUY17QhW1frPcY
0DAYRZ7uaR6nxCh7jFzoKI/CsQFPaO/QhjONuEmhobhi2QAOcvIPwwlO3fbyjvi3
yQGA+Wfe9yF+i7ZtUFmBU6tLnv8FatQeUFXtFT9fb313CPftGhJHeNtvmFlx2CTJ
/+lkm5958ALCaEXH8br830UMvxq8zhfWrhJhXAjuPg+SUTA5oyKQIGbD7JnV3EXZ
HDmQNkTu3GIGc/5heSS6/ewLeMsEa4+s5xChYVSjm8IcAOk6y9j9fdRssLMhQDJL
64EzOe7deE+G5lOVR9WJbZX27i9Kj/1OYrETUoHIFDmYfmTnJBCeC/nocGpSSpSD
M72XN395w8YcwT+1U3CGKAIT2zqjojBRpS68y6r7eecPOHe5ud/r+aaucpaTZgf/
i3jCfuZil3lpPUbdt3XZYxrtefH0bD8iuJSRc0dwX6/nJpK7ssI+DZ9Jw8JcbcrA
g40T5ebr1xc0pnCvAaQGctbSFElKoWkicWyqKgSUjD3mKS1wOGzn0ig6hGM8hInd
XaPmtYyOkzNVXXfoEh084PakKZAn7A2LZS8xOWuwxedGBLZ0OfC0znLARe4Azj6h
cwZ793LuE8+uJKsUW6JRQNZm55JRqsWix9FqXexEOabVtNJy7PGuwZUL78l5u91T
5QJWN7t0KgK04S1zg66sI2+D8IeyzN61Kd2a48H2E45a4LtdUYjb6mf4UrCJ1Lsz
kDICAMCCVy3zZdJcocwl8ol5yOEA3LhJHgeuF3Qfqcs3JIjB8C/di5vHrW9pc4S8
JJlQ8QRFZkr4IVck02PDaOR/KLTSJ2DmqAT1t3H6DqeN0dKYrEtKI5NVjsXl0tYJ
YXN62MYJ7d0NCTgdQydzFHL2yWTXyGRRJM0B7yh8Us47LGP+mgSUvQ3VfOZXnFSd
OZNTzMC917qRY53Cjp/3C6wI5q/Ix3V2mQVrLmlyS2ezOH1ZNuGTgDJXlBRUTmDF
nIPh5XQU6wzGPKPLbfvWeEgErxOlL3SG7plOtR0NFYaI/oJ5Mr/NM2kYPUcQYmsE
LpN0arCRroTuAvqWIZzDAETqhWo0PgDDhV3mMAqxEu6PSi0l85nYLoFGeoWOq+Mw
dG6aLB5ZWLXfjaWZAxImuT1DWswCk0VOY+3LAOL22joAgLKAOzDQbBGyh0hLjx2K
+xmj7uTXiq+PwDqETru+ES/9IpuYnYGWd9fUIRuALtGspBaPDqmYJnRiBZ5GaKwK
7+qrewvBD6dQsMTwqeHJGoyVh9WjvYvYn0Jua8J4jmRPdGxE2ADbjj7TABUq/6Zv
kpbD+/8Yv5vWwO+LY1qpHeBYa3tSwv4dvbQkSaGhO9XgbWG0Hpn1U9zilCpiIOK0
RLkHt4DiItV8Ezeqn2JVET2T4DB6tDpNznB+kMov1Mdst3uAcZlVnW5Q0+qShrwl
cbezPhYjBKzvtlUc7Rz4Wt44cSnfk+guustouD8GJcaNkFMjibymYj0hqjh2VcFM
n8jHtnHVXMpojs1PsAg4lytwqrh+GqJBeZMxcJUejznX0ulOuqCzdwR9Xmft9X+Y
6Zru2U1wWketYAqEsQ/tGZHkwR2wqxoNQioxiw6V0Ds=

`pragma protect end_protected
