// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
yrUcuWlrX5YcZ9qocRLpzkjZDiYbU8zBWyhcEsmDfAM93oI8Ma7SJE+gRAMY
hWdDAj+KWEjL8PQzQ2xedfHewJONVSW63uZFDnxFroyX5/sGv0FdNV/wxL7S
dDdpmGfRnm31iFBLQZNjYcElzK5H2vZwBzABBFMyIC3xjo0xCkHbxxpFzemR
6LJ33CV6Nswkd7ug8fqrsYfzGul50jklqXi6JLqjW3p4/fAYkJowW0KNYqS1
RQCVo3dsTzfc4lDrqQBEvoWBKJ/lamEmCn+4s5ekoGd+0fyrAvqO2gx1jid4
xYJEnoEdI3EZR/OEinsJqvzy3A0ycA8Qsa37LQBDMw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
pIQqzeQ6Sx502ZdWsj6mgaOwx8wVBc+8WTN2iBWDZsgU5jyiIccMAQM/46GS
c5BIKLh3+5tsANd5zQxhJq71My4tXTZUHieOARJjeQWpw9eu4nP051Lpcqt/
eOrDqBzh12Xfhb5KukYl94l5NjFcARbWxCKFejnGrRTobsdUuljVUBOUz2kV
ThMZ9tru0AFBi+J19RZ8aoGNnjLgJ8HbRfNggkOjNldLvQCZBzwHbfV7gO7o
dQEDe1R39ug1B+IGtC0KS43zr5tnOq/quIQrbFLnQi1dWXUqZKKa09lvLrru
wt708hmYGbgpVGMP0MeTkIl5JcaIp+vRymW41wmRjQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
GTENINuaZ1XGnCbtugE4QuwqEUxTNT7yHjsm/0qbhKCm6ZnlnRfKwpKNWo28
gtQVHQ1ozgu2WLjOI1PkeumGYK1r4SbtzfWJIc8PiJUxvi88qkyIA0gHxB1a
/MDOXKuO2fjxolfEPShCrSjS0rJwJPZYleo5j/FNV93HhZo0mOisibQmR6Lx
kRA8PY4O1BjCbum/INDGvtR9dHYtIAOrTw+Q/5fsYXBJM5Pgx8cTFItFIKS2
zA1B9durgARIpiOGis8PNvk9BSk2q2an8bHR9F8V9GyMG1g03uoOSmVVDWa+
m1rjkLsgDf0XCtPqlhMJ40biKEnS9lLvoUcNNgNTMQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
lN7E2axHhnLQBlNFFmAuPfeb/t8vPQbn2H6q33EITBLUjZTkzWOfpeXME7NC
Hi4Z2Si+qrdsP/EgbcQrbLeD1eAcxfjm66/1CmDBEI4K+X/r+eSSG6u64RHn
H08MBKbxVF6huUMdA6DSLFaNNycJXqTGAqUAz5NfvdWpoBKHI1w=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
cYMgfH4X5e6Xagq1pTW9Dj63RLFFX9yIlzpWfuejhxk5AgW48DNkvNtIRrzB
GEOiQ+yB1lISsNGy71F9un5pWfjEDiCgpfnN+Z1jzRm4d5Td6O6WZg4s+//E
hjlLqtR1tO8PpwMRESQVUbLEp9wEUy0kV/fb63adRfa0sxdGdfQS8NUHckRf
beVZIwridbUQEViJgWkT3u858pqghlIYHluwSXvaKGIYX+2WEdOHlT7subMK
WzmC1nyJkViMRCFMTAbZyK+JvCptCahdyYXamB/26cQvN0FN+CewkEbPVTVR
5hqcjax3hP2gp47O97wmjj8J5pYNcq55qUy86UBA8z7qdbaz3iepfus9ZDBY
Is7K1yPoOMIfCsVviyW1Rlnpci3pAqLXFkH9O9QFYhEJl36aEEwqgGVqQ3la
XQeURTBfq5+XW6FGHBFvF3/VG7eD6hV55rwBrpgOZTleLvHfVHVUIZGfggcC
XF1Vwrd0eY/CaS2wVnqtRMOmMGYSDywz


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
JMP0egd2VB9L/MImRuomGktmnlPiNl6hg1Ia43OMElMOYGjfptNJvAjd7Lmu
sL5ShDaM2srxD8/MHFJvIhPd6lvqjpGB9JGDaq1toryrBzaF2bd+6lTRcg15
zd0Py4CmrY/p/cgrIwx9dVJist4lqwGq3w6qANBoaSZGVSsGNak=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
hXnblQj5BqSempoKmj/sCjt4xpJ7baN9o+RyUfSD2JOoWRj7beSNZegcIHjM
aqZ7uec6sVlsxUdc4QeqI20EroRaLCxTVR5QCaudYp8tngsV/t6SocAKbQ35
AXLRHMBwOa8PHOGBACNva6W43VzzLv30fvjwIr3WZQoqb9cRXwY=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 9584)
`pragma protect data_block
CFqIOCFgDipvnC3vOhlq2q954WtwKs2+OL6OSOhFzjZMU5hSpOrVMiOf215v
qSLGthXHQr5+gbaivQ1SCclVHfi9NBHRN7EkO4NGYZaDGDa9McsWq6eHkVzr
Xc3ou2swu4retEBR8/Brw8IwmGjm+uAIvHX+x6+MwsgSSv4UgHR9DXA7JDV9
4whJlk/Taob1tqPhJNMgyiZ7lGYWnfFdY0X0HY01MJKIcp4ASFSqBh5Dwh7r
GFDtj20o2EauC2UauCvnRu5jNbOQCp/32A+aXSC45UA9QbKSVWGZARjKP7+c
8f/KTvITM+VeoNHw+h+v4AfSJ0ZZ4sN9ukAnj+OCFbSZoji0cCwQuZc4w/Yd
M1uHX+gzk+xz8fTujy22mFAC9u+L3SxjKpQpbVwWc0OWiz27e6zZ/YbtiJM9
lLeu3pBYJnIWfd6ykZucAJEUq1EWCQo6qxPFc4WvoMtOGBMRH903a7GART9w
US/8hjq844/FNgJ9dRtK6XBOXkDdSmhQgsGaKZ2brw8JTNPmtClYPoyxlxLB
KjVdCYHoHQN1Guh/v6vUo3GyAnU1c2LbYWFztENxNg+Wc5r2VCY27BSeOBry
wQcvBcZS+T8BHE1G2dPtoaCtqPhV339WulGRRJfC0xoSEmHspvOoxTtUPeL6
5ONH4zEQNihJlTvlsBWZ3b0Pa6enjyvSDk0YsHPDJ9+b/dUeLJjZ2HIjsEjU
AW04yAM/q+vw45ipfRN99bmtzmfmvxpil6cKv3tki4UMb2Du6Mk4+ovHGNwV
JukpjsbyxiXEyfskJhVV6oQbMC325EHNIpudN1+yQ6c6qiAjnJCkdpWMFzwb
Tu4WAjc+C+bicgEGNOfPb2NLTZTblCW69HZLHmNa4IZDuHpt+DJ1YTSLbPUz
LO7xNQzt4EQVoUmzTSA6aiu7k7GFSeXZBba21XPMDTxP7+HF64freT1x6DAO
1NXvBRYU4zE7FRgvBw4zRafOnCwRsbnY6dZ3d/uNHkka9OGMjcQIdSkANNub
h893YUEXpxDZN7jPmcr18VqXRBQHCnuP6kD0rWZn4rofeJ13tMa2AEMNnk9p
sftnKuxLsMawPGfJO0wlsJqGYGzvgWBiyMIueyXe3kL4JR5RDk+4w9DXHoC7
OerJOLQsVbWDV2knFpee7eDVbXDk603nv8ZE4wt8jUi5L3tB9SBJ2JAQQp2w
2EpnW6VXo76Vlr+YFCG5JzROfqyBHobGtfnaBxfywOzxI+1Czt3gTHIUozqA
tFlfNqjgTUSIFrBTPqLr6Mu2NKgw2UZ8ZxADCzDZ6gJiwD40dd/4GTCxbD1P
expR5EByEr+q3ZsEKcp+Te36cjyPIFFyq1dSycxG7VzwSL0U9lca8S+QK8QP
+IdsQ0imSbikY+4e8DNLEiaCVMFTSZV9ixeCTeVkyEMEKEwiQvasNRF4juCW
4bTU2TvyUl6cg5TLjfCxc0a/Zn110gCboAfFMwooc67XHOqWSgOld4SJXL/K
HBXAe9GymkAeEkZ8pkV2XqpJm08qfgijq8bYacPFZQeSfgyL3HaWc+VxDA8o
RCmNh8caCJMzChJ9GiBPWyPxi3qnnPYoZsZXdfmO2jItKrmRsVVgUyfXErte
SgZHuwWpvCnP4+sr2T/nxhkTj3PlT3sPv2N382W6jwJlDgHTkL3Do1/Q2tHA
Xs9SaOBC9cC2Z+z+V4dwF0qW89NpJM4mHhTNKzozDozhYYG9JKj9dW5OfOtP
wn/uqhPWFwIgOYrMJtB6UiJ9TUytMXlm/Ab6M5ILFuwWeFpOVjs/jIXALueK
BLZ2Cuyh98H+ea/z4bs0UByPNCyimNxCuOn8xqkfkCyNfr/X7jgFvixCWojz
fMArRywFB5bIsyZZPFqRMaSObbsjPg/hYwWYcG4t9ets3VWuwQ0aSUURrgJ0
JL9IzoS3fiAI8bdtHgElu0XJKcDBwOzQ6PZaMQKAdTlZaH2d+58ELR7RS/C5
5yZfy7ovOWfu56i4Vg2ukC/TfJro4cxqxdNb/6NvP+1Qar3e4O0EMwQJI24B
iajhrNhAVbCivOdXhT/QVOW9m2Ld4KalhqciJEGM/wtXWgWg7Jsq0icMadE4
COSpaeZNojblmEuZWzRi+ggcltFpqzuKoPK+nUN7SD7MU2dRtuLVoh6ej95e
Fa1H1iI4BdDEan6HESOPwbeDs3UvlCFzTX3Fe4x0Mg//LYLwj2U7H9XuOBYK
CEcu761seV8itW7h5HWlFzK+gFmeZFHk4GNeT0I/YB7wQLaZLlUceJmSbJ9u
Pf0tU2tH2To62T2mXqw3iT0TBOAgtf8RAIvhCOdAo/Hk0CvOXnlZ7ezcXe8m
s9/BJ4bTXQEh3qNRDSV7MgKTBEG536MPy8NaYJ7s6GPUVG1VOSL+3f76r3Al
dv4VsG3qSHA3JeQ6cqQTcwEF8ZZF9DxD0NGJGsgg/ne9D/jnmAZH1Y17ZlwZ
8p4qR+UmXDkYsjGiHLJ1Fbv5AZdujQZElcafwRd5bSdz7Azv11dQMYgeKE2G
vIYZnSaD9t8RVS2chfWZHcTHkdIc/Yj+ukHBCwkCjVSO39kaCOrzpNAGETte
WSGY+VD8G2GibY0+VjTzs2wZ75vKZZliuFlH4nk1RsNEcDpvN0aNH+wn7Hwk
/Rq92emFUP/2qhGvBkAKprKKfDUQjETSz77BQa7tRvzPB5G3sqN1rX/1e/tB
/cUJ9+XwO0rWWFTmV++rmRpJ5RNElzFyZcp14HrsoNaaxP74vF6T8V0X7IAQ
lHSMRSAr12W2aC0t4F0B7ViCYeVtC5i0FJTzEIa8UIUN1VJzp34Vonb5GxRs
OKiMI5CindTPXWhvr8OXnK7gklDi6qh/5dhG9XBTSe2W0he8/USP4aBkEIbt
IrZvb8JBUjFEgp3QLZ4U7YZErYZnHvtMtiJAe5v0r+LztmnAadq6q9t5zS9T
WdrqylJxEiTWmO+m9By/vULe03340aQcZKOU1HWu40gOH+DbX1ExmYK41aZV
5bNZBN2QEBsJ5wP40mkVbBWsK04cPLWmjnhHI1BY8Wr23IHt7QRIt6ep5HSg
/QUAec5oi+ZbWzXy61FzmZAaOVrgcTSaMuedy6ywI6G+u7TCHA75+b3y63sq
YNPS5oW/E5bSvJgnFUmay173bPIaS0qYdSo/h3KAkz++Gh5sDyRjSk7+k0oj
NnjkmdO/ty6lHMT/YZCiZ5Iva3rRItqjfnfqHZDvw7RJoVUW5j3sWiJCIC4u
+RsZnee3uFiKWzETioLYgaXYaIOaE7PZldtuqDL2VhLwm44EZhFAAVZc+LpH
1I6a3iar/cMpYIWJvXIQdZevk7pZN3QukhgLmNiPTNB1FoSjY4hiPmmHx7bJ
x7lkRFNfYKEVbUIfuVNFqbm3EzELeeVVVCqYAbYvtM9X79wmfamjtB9uuQpS
FK9dBqqd0vGqY2JHjr4Z5LYqqm89PiAXzMiREFJnyN1VJMcx/XM/E5OcoZmk
8TmXK7G+JiBwmEMhFV3gW/oEsxuo2AF9G7x9o4CnGw4++DYvwGLaU5hToyOP
1HNnF6tyAAXpY5JSvQ8ebYzZDElR6N3Y41pir3Do0ENgysvaIqc81SyLw1w1
4WEBGHHYnYKfyasEPOT/y/3RPtFFv2yGbw2VYesqCG3IwFe91hof5MDEbA9Z
ThXXB4Mzs707gp+9QfymP1I3S+ZPRux7cNJezpTwTgwheLUhjkENCENIyfmc
/AZa279uvnk7DWRoxpLrHWtF/4N6J4KBe+8FZ4Z/yy1j4JUHvlI9F1Ro6LEG
72Mca95vu78d45sUJc+PhUoY/mZJ0XjE7nIQsyhiULyAnhRtubq5B08o2I0X
Tw2TBoyjK5bg7z9ZEGxbuqFiTiXitRlLgdygWi76j57LPOSsWGBAP2Fz2ox+
drQDAJIS+flQJOkd+Z/eeHvDw2OUEVOX2/JUujJj2UwIvlHiJgHVj7MKOv/X
hikfgNA6HElgKED0BzmXoiPQgysBRR5c3jHrIRx6ibMw+unS1U817xX1XZqy
jO699lLNUbSEb8mucSXu6daVmYJBaIEQQEGlqAdbE6DebsoRMwAu1uvoFONv
QqYtA94I427R6JJN0mWlsJgcO/x0YSx8dlDN9jK1MHuXxLcQoL3ZNXZxaykQ
y/KyVQUN74bLdsoYjqQeje5NebGcVbXMo2UTqg1F5WgxH8QIIEfE01TaGGzk
/AD9utXJUqLOAlupl56HrC8NgJBHyROdYx+cg2jG4TypOy0IaGniRObygGBo
sB3LRpz7F9jR7iMdqAcDw3d5FKU5Z5dfq5CMlO3TpJ4bjJJMqYpyeuXsKAoo
kRmNQtNok4mwiiP+5MtlQ0koErrOQFNSJL60/229Z5NQzmOZ/AW20/Uuaiqj
bjzIafWgAtMyWpbcBr/HwMqaclePyERnw2Bu/3kL/E6bSqu1+Bx8bBgVQcAy
ZsbzBit4K0xKCGLPQ4KxrQh574ONjcmmGfmtNIg/lpRweyC2zQjRrDU7WAM0
eVQy8FuLu5SW7tZyxuIu00lQ/tbVnMOHC/hYHrJRSiM7VFAEz7IA8uFw/MUb
yrV96xakVhaEBW2EuBvtTVCCkcy/85O3yzUq3UotwGaO3eQHQm54ft1HKGxm
nIDEmozo+nj+aENIeHChqww4jr6cAFdWZpdUD1Flr4ow2wpC6LkSKqixBYeP
rL/D3wUT7CQvwVDTYVf9F+n79IZJVudIoieoApjZlHEUsHsFD+70d/f+34OW
FbAxAHyVM/VXBEw0A62zcX/pTHLm59jFQzn5xQlQ/0HBSWdBAjkdwjRGdx5P
3UhyzQHubeqyUyuSt7rhpkqEejX9mBzxLCAF/yGLFNaS0kn1xa382ysBHKcc
pXN5LAVwmStbx+Br3R39GKHGlT/YbQ/5eQv3oKVoXl+tOQ9EolDyre4buHTw
Y4m8KxjuUxa5VlJ7xhkAqrjTQ4jIap/8yas4sdJBRFOpcskCssN1LUh2gRdB
N5l2DAIJrBn2D9wGdtWSAX6Ci5qfFlw+KOaG9HJb1Yyfbt1PgEOtOsZzxaqZ
dOp3J7plHL+wUptdU5qhTCxfiyhTlRJr2tCWbx4/Sk7sQPP+ZjBqKAFiJHKY
Yqr7oznuwoUoWoaGXWZBRadRqLgKvXS6VJdmF3eOhhqfatH5aq0WdhqvfrZa
f8WBuuQ/UAuPp91tKEcgKGzOnxjHo/96FPGrXBUiqCtF7oRrfYYafTd2ILr7
JoR/RJ9iuOUi2AfD0hQzk0WOkK31xnEmk3w6ia+UPtrz3GHC3+4EwtmnFe7T
t0SRWDMSSAoIpW/zEnGLIE5nK10dk7YYhy/uYkUDmyoV6CfaibqaYoi5wwmI
ZhcaYxtWnp1VCDbmI5gHjPkRx6jHHsl3sz6Bxj2esT8m9jxwuCrRoX8ffm2n
ErA1yB3+K8gQlPU76Oi0qahdfWcT/tZYMj78mmrwGPc7JdZplAsHyBwcFl6L
TVNag3PYUuyQbNOb1+kB5wEYVnJGb7Dz2LeZpEATKr5tL83obzyl86uKyv/Z
stcB28VoJvFGH5/8i6WdTv3yw6zL2w/vtRBKVdeu6vMIDbH4a65ISDU0HJzf
fNzVWnuegC9uhWsmPrnyRh702MzCPpn1VdC8kRcWfpyJ2tX9LoBM/JvKxTbQ
Vw6duFvBM1OyYsgskYPIbCalEpLQgfROte83kGwS+4ujejUdExD+Dr6afTZf
Kp/pZ7J1DNAI06vtoZjYXbBpzJEX6sTlD/VJEdHYr7qG55YKiWokkwR1zthb
0Nol0e7/b4uv4EOR4n+BSk8DBrVVC+CyHEcu550crHp7jQ/FfCgmBMGqG7lM
Lm0L0yUbzToeMc18EWcIXI2eTyUzLGwwdIJB98pld1jcsQQ6dKO373j5zAme
nGKDz+k4ZIOLH1lgd61iCFnLxcyrN/xghZygByDIXhhTulcX1zOIg5KzqTmI
4Et56rQ2S4FnOotgFcmKGlBp89PdlZk8nFQXQk5x19xWFBG8Efl92b9qaoVY
A+jBkvfHMnriZiaBggPOnA7WCKjytBQA1q0ETidlXyiVeLiWBRfG+SZtwn79
/ODRBlvczpZUGSW3WPmm1QGbsfEC+lv8a/Y+h98gEWIgmI+yDnOjSdWY+kuT
0lfLkmD3abWY2aCUMImSkf78HpmroLMF/4NWYDMP19gG0q0Q1gARMj67ulQP
k4c++H+92Pn0LRYjvS5Bm+C8XVoOPqpJAOgubyd7wPGBzlgWHO+cQFkx1hX3
W9gtenUn+MetrciI5DqW05+wZ2fe9wdrCITGmcKEgHsgPfdb2zUSBzvvQobi
jc7fa4KkwEE0BLk2v33bNvAJpG8SeYBEOWlNLOkZDC+aRWUpoFjHi3zhGjS9
CuLJfjWPCRRtnKPHq7T/yPQILhiHTNxotE1XQWCrYJH3UWcpyTME0irQ8Rfp
NU43EqTJmEafKkaBaGhGznwVZjc3Z7QyRGI4hSO9YmluuzGiirzXjOOgu25i
oS3Z0TM6oXXJLbi7qiXzhm9tUTuGyLCO695yaYLCk30a2h3I55ffXtICRInt
UQZcL7FazuSWM9fngLY8Wr8+YG3EJ9paSGXoK/h7R4CpZa1eibvs1Vb6eB78
1yAgeOZzAKUMDsBoLgpXr8nkEi5zFyJGQhyU4KmJs/mqetrI5x5UxZqGUoCR
ONhVJmLgu3na/S0VyUS83n/09NqoQf1a3T5fftUujXLNCo4HmXPQZ0CkASVO
T9JOX4+Il3yHLOImi6TMy2nphW8JjNrVw3oZf2N/1+qM7h851cFqzhWO7Uz+
OWytRWWhxAZJoLstEHUWcFfSqrEsxa213sjah2s2KUPRLgPZEPatS+zqcmcE
QZNC2OYUjcEqplYSPhdXpD5qgoD7NXBXYkrIEmuSXv5+mACywLPMprz6icUw
xXIlF9hnQEpypK395nbcPK10j5Nc323weHW/AEpBgs30gFFXftJmgvaMndoV
fg4kcUqqNyRUaBT8AsqUrFzLFZmLyBGu03Eva4WuUN/h8jdXGmxAD5SUoEgy
Eo3/+BnzhdAQN1QTKXbaep/+np90bGx8rZcxgyHDqVH/V+8N18nmuOJNsgGi
sIqIJRttrkc3Y2d33EnaxeapiF9A9zsjOys08cQqHl6x/k47l3Dzs5O+KBFv
PbcAjoFLIY+t5RZEaponsETxmCvz9IEXMAueu8Fj/LZqRJ++vEpGzeBTixwm
chPShPq71o97+hS69BgJPZ4G0FlELYGU0czrWCSlgGg9PXo7YMz+36K3mZ3S
4dquoirA53KjhBP3TaStKauA4Qy83H7RVTCDVJ+azlz4v84/5WNPeOrU+8Cn
bO9FgoTdHuvyqA7IH+7VUt5BNQGHFvkGVO+5FKLyHHBp1jEcEFa1dsHVX/rB
G5rmNF7pEePlkEvc2R4KNvXzHzQ4HzcYk00xC7p8a42ivzGskCAd0/8l1PuJ
LA2vMxuTTdLYn7NOyFaM2PHhjAP64uiWqQogNJEEqzVAsiSdjXQ/dN9gZEf1
Ek9imZOt8oWenFlXGcZNhcTuntw8nQNzsIwBByNue+NwC33NGJ2LzhkaybDk
C0Rt2sUnE28ATHNcXsmpcW/L6jbYTrAB9WEvu+SPy59NCS1Z3HYb3Pr/hN/Y
QbcSz6fcU/iBH2dQ+HDqYEOyRpkjaLmvfwJYowwfLDSwUYxFB3WlgKNjdw9y
AK+TpfIUGFUo5z2B75zfTaNdXHC5caLyqfSHp/pnKT0tKAoOtidP3VBinfyR
p1RQ8sh5VwgiH6lOPFLS8P36l/jlOM5QbD5G6BU6m84iH0cZcfJW8mTRUR3Y
MnjpHhlHl0PyrlX8ZF1lkDTbZWOBY4kw0kGK8PU+aH8UN2ERjAINQ+XDNkxn
lnXkChM4w79CJQ5u6V3GW66gFHfs/irJ0mtzTkB5blyT+GkCSdZC5mCFzY2E
HHDk1WpbqqSizmjjzJiT+82StNpYJQtzpUekUeLgbFLJjONkb5Ll2f2qsgFm
z3vbT4QPrvpyxjJUwYplsyDtSpYZch3fFJaUCYrZczxMb3pEIczFBoFnAFpo
nljH5jGoOZYsIOhlJMuHBtOf1KDvISYHf3WRk2F0jYWQrY1QSwQ92/EPQxzK
TMTpW5rs5d0BONPxI2O5MoSJ8vQ+0g5+ajg18pyYhY5dhyyUbL6fYh7QQrPn
fRHVD5yvr1vEEuM3muo6uGlY5kBUlrjqNKgH1vt9bEG4EzPDcOYQiQxkI6WW
IKjP6SvbJmPEb5AD0xQuI3fdsiydb3lpXt20VxtqqaOSqZtZZz8ZxPAwYBvO
CSgBB3XP97DP1Osd7DWgN7o/WvbuxDmVNX2Mvmd6VX52S5vIPlzFJPzhNg8O
0Qt+Plh9CW7VnBLcBYD3YlKMnRTmTZKrF3kvJWGxHebOEh+mcVw8ovRF3c2Y
hc4GZyIfhGcymbWsLbTeYF3iVNVzhDV9inAE6KB3tQ7paicj+ZDRLlwVDZKO
nJut1EJUCGaea+8lSnO9rJ0hk/v5m4QoSJbL2q8NYMDjY574DrANnoUHiOLZ
yTkQh54IBv3cqxQofKqJuVau2JGucOkGq5nAnAJrYmKAldZfyRySjhWXGzyr
zDvR2WsLC+JNLub1HJXQY881swBUavlj2U0/GS6/gSi9RHdpQMzuq9qmycBQ
g63wmEfwfmjlqVDuBcfKCEto+ospkQMJQXjhKYpZKSuw0dYORTjYfo3l0omA
nK76nba90VevUJJ+UsDtke3qf5gGK9IJTKaKQqHA7/pWabv/zAMIy5iWvQA1
gX0KmZ5FlJJTFAEwZQVTy7NRe07ULQXfV8oFPfJBx+MrW5Zzdzt1/AGj1vJt
i6Xx1fFk0zkoLEYvD9jyY30nxcAykOAgHdWP075wrJtGkfI0d+MUolYYlLLp
nwsGMLX678Kh9SOqagqAeth0a10T4quQBt+F/zIs7Gj1QZjzxEyGTDbaMWHf
ARcAnRPOvEaUiK6m9y7mDsB9IX0/yd302/KXVofOqqvF8vg8CPkRDzP2mxzm
k5PAqRoi7lfRaH6p91Unhj1MYQ37/vg39foY2ewZ9r/2h57dYhIs/r3LDl1I
efS2xVP50k/uU4nauM7TK7pHimqjnBwkGHLEJaEPNQHcEgQFsgd/Ih06eNXM
Fj40RM+BP3127OOj9iYpPlihoy47wKrteWieLIgYJW2AfSvGNwp5MCAC0CGh
0bHjzlr1LU4PkqvmTsirXurvYc/OLHt+cG3J7U7bCymdxdRB25IFtmR/QZUI
/s9Qg8kl3UhR1v8CB6my4KCvLsU1joxAkaI4tcLpnrpoh9pK1X4qog/qPw2K
fjRbd61gKOidimFUvD8+WxL+J57eciNdgYa0rrndG0kgK19xoaRRVaxszwn+
pkAKkcQDfKAnPyBgMCEogAJPSewJBOmmXsSTZ1ZhDxBailfh6r4+fga1RASh
PoAfeGJg7KMy2NBKtlS80OAmo26RXU97aN7Jx6QyN6SdmCzZhg4PkkenbrH2
VZ+2D4ITog7qZZXOpvx9Vb5ZYAL+ZWvdKFQGYvIa/CiXUNsg/8DcaXsVmyrW
Yr86ckqxFCqTJYGieIT8yWfyplb3ntz0yfXa7ucqM7r/ZawiFE45Ny+4d+mi
W4/vPkZBWaQVmtYePL4pJqaoQ9/L87BudVvKZQXbqg+o1OS64/zBKG7J2xgG
dAp+wHd+8b/ONSet4o21MBAwHQMEHKefa+45C7USBwsQLKn+WD500x+2B0qv
iftfIXmFoJ5fLRrXGmbggTgQuMByiL+aBOtyXLnp9AA1QklLYK+hqKLPL6GS
hvJyucsY19Ac7syspyydHtcQEz8dSi+NLDOXqIBsgkqZ7M8DN08R0G4+LaQd
PE4FAsAt8+ADaArlgYyPRIinWQrhj4q8PpfqaNMEcRcNPtBeuKRfJ8CRPY6/
HGm+5el8hEBYI+f3nOT5h4z0QBPH/EirLx9yFz8rxlSTviSSv2OTnJkeJ6IQ
G/Cru6GE/naRKhQ9FXcvjgelUkg0lMVLyQZZ1GvGkGIlgDa/f+SkDcxi11OC
lJVyK98exEBsPLWZgBSDMjp3lxKGKABLi9DwVEEqUGbEOfupJDigSUL4/EFg
clPHGZbW/uhnAswGHTVWbW9VtmvgNtN5b5OLVvj5bJsWqm4hrSX9SmyZIW55
JYzQ9gFqip3yXmgnij4kKNgfz1F8BW2OrvOweiCb+GsZkBjNMArHYpaXlH2G
z+61Uq5501ch4d2l8798FrdlyyTjbiFtE7BtpxAY6YaYEZ64FYvWk/Bw/GjE
AbIWhUp1lWwMxKmFiAhNVjL8yDYYzv30c/dbXYeQsH1h7kkwFcRWgFBLlaSh
bwG1M9FksjFYR1kvw453khhnVBWbaA43K4/pWtlljrjo+npmQI7a2/bC5e5X
GGmHLDyQbVPi5z7sHercHIRlqM6n0cq5W4+166giewHQ7iaHdBN+/4J1w7wg
6vDo8XIOF3TkqGexmRgEBQjGO/tgoeU+FQQcSRAcGtVutdPvaWBzsgzSNMTE
Ojmz3ur5PoGxoVVcjNL1IkkeHprrxgIjJvdyuavwX+Zge2jZ6WUFiXggEQxQ
8DGCQqz5obHIFX78Hiv74O2WP7cF5/r7LgpV2+si4fx894tFvo+leXr/a+BR
7E0xP6JdnMHllRGg50Z4GvBUDJUnQKowN94K7DfkO4HnMqr/CGGNr5u3ok0t
hXhIXQcyvVg+Yzuoouo8L/UngAhDZJpa957+K+wC0bSZX4bZ/ZEFI17rNTe2
9d9TVhB1PAtDDFHybCmmqm5+uKyYGPgtN2mwhCqpv3lY2eh3WIPg3ZmEEJsW
e8A6qota/ElR5Sm85d+8jq7ZGuyVA355rGDV8WlntSXZFUFCebPP6QbD/5ND
rkHIMkCe1ICeC/6+vYGF1+j1Z3Rypt8/A1pA5CKR7EFpL/UKKLl52gUugXyY
4rP+V3GQq5hX/pedVsydH9hAPwggfQ51oCaGLsXcIyks2mGpWLG/WJTFkEw8
v7Kjoi+Uy6TchsfLR/0YZ8V+EbLeOC1zaPNB7Vwx8xfl3OddISET07xLEu4F
xouPwcPMaqNnHGa4QihIMGM97DtFC2l9Ap4x4wnczPOHv6Wu65KPJKw4bdYv
CxqOdAT74aDhZAfwiHGvuzBu4Vrfwjl1WOh+2g9+E/g6+7RE2nGx9+qm5BVK
fWoJ9GQJIfyBR9TvibGLVQByfPn7UjUoGo0DtphE1T3eswWGi3Ol6xx76wm1
FNQ0fMJxF+BXCwlJpIvl97cw1MS3phZD5iDL9R+Ov28if5g0ffBs1l2jFVCO
VtqHDdrbLsvLfsYytvCBYDTVfqb/Kz9Qn+mngjrOKdWkr//O2IVYc4IeM26V
Hd9xbK9dji2P8XyOuTJxFsWpY9YtieHaY5LFw5RKl7xLN8iP0GjVLu008OK4
+VfE4R4BqHTtjPOvhnikrjL2BjxXaSBXhEM9aG5utJwthKnxjrB5HpfzXq1q
cKFuAEHPXJnElgX3DjZwTnOpNPLeiy9vDfWfStiuYETbfLjTLGyfaOH1MSm6
p14rCt6brYog+TZxCveXxVe3jsoQKYQz/9fUV7nuLGKJkhXuopQ8gus9w/2u
3kfb0ZLZevrs/TLgSwFmpJzoIyRiIoqomIUC5TtFunEMCsYp9AjWPKFfGwu/
5VicuP4HETRXXaSVjJlkG5WQxOlH/8m9FvMjkAXCCXExLwSOJKbIXCRsiJNI
bH5647RicVSFqUNj+w/5+SQtKwqrzqyZb5i9PKhyFT5nLMUsDQrPLx8jBsG6
ZLH394GhlOSOYAyBN+nQ1SrvC5oEN1fSqfc+cOORSOQ5u6ZA1MPQCi2CXrdG
Vfn/6bERZN9J+KXT+0ymXkCfdZJ0J2wqLYsTdxE98JT42vz/Ar7BSukzGAJ5
VrFn6NPxkNNySXeb0BuMZIZywHX8X586AXi6wmTF3T90RYMypion1wgXY6rL
/sVT8F44tXIB/3jPAFG6I60IIHmvmkIToXVB77lMlCDB9xm5v6iuYLdoA1kC
KrRyfgt/gOyrUJNF7lqacg4UazsohZbl4rWhbIyVjbMKreL1UFuRgDCBoYYc
WaWHbA0cUdmtt1EuSXPxhJgjDi9PdCNnkQPkcMJsABDyDHPEC31iV1n4yhEL
yqDifw2xinFAx7CHiqZTPHMREMPbQFPSG+ofh8y0qQpVNkrz9SlR/7YCbMz3
WcyYmTTpdFdTnKEuXJONIopJxkmps/dyUT1no7FPSPwG0gjKeqqWBO7AwRrn
qo4oSgiHbCvVG4OFN6/PYTs2NnejNvAOo2LatybMAdeFXlv8I+Ov2R96gAlX
LcPhsWcX+I9wasILyMCO8rFgSlVxYC0/x0WBV8NDwP0GPAoROHr7Hl2WPkTx
7js4ZTsRtKScEI6get7qa9bo8JtzlI4gHgJVycL5EiewC+AWAuZA6tU5a3/y
zVxpg3Iq25SzFDrPypezQK3Ad9ZAldfJAKjifFGI7LTaSsFsrqYgdlPp63co
zpsqVQqPeZQSIZoABp1CCIMDh7nJ46zau2eBO6r2lwXaZ8Ih8ZVyuBcRJsTX
5/M4FQf8Kv37Bkp4thFWiUdk2nG6n4+kAMutjbJ9jZ0q/KHdDJhMm1chrYdO
1DPP6TVDsTjzQNvEiiBeNvOnqB0mxFucbP09OlEFBIh9xjU2jtQ+ixEGwtJz
pD+/wOC3uk0yWndPTojkEReJNFIjdWsAg2zAYelV7kEz5ThMovkbC+BgojLF
ZZitAKloqdlDeXmbDzxpoDOShsgTwDgidN+lqhBfRIk6oibVJfs0UPT6KnA=

`pragma protect end_protected
