// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
rn8tv5fQuwq1IcVVPFudCFCcfgicdSy9pYEL+w13lJc7ZOjK8w4Usj3DwZ8du4oZo9BdND8/vKba
1Cp7MVAOgJ6S8CkGkZrwuyYbpzfXEguO7QCnx0JtMhZ+cwUdFrR5e4dcvHW+DaA0XyINIvqad81r
qQGNso/3Ey7GiscjRh3HvF+6jj3vSnPArMsWEYWShcRArk6xqzZjZzDGtZQ7qw+zBJTqVSQ8Dcbb
40Hjv2S3w6UP8UTP23bM0VDgJjHoUgLho0fuYY3RIIwaRBAqMS68CyP+2IkTPBlYiAYp4BKm44MP
jMXCISR/EGFVB+c4D13RRfEk7sEZKPtd+/G2MQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 10000)
zu8CfyudU/4Vne8MPS8HPQygERNflFwvSZPl9U79RNRhd7aVFKP544Avp+UBruPpog/O9MY11oQ5
g8DQbLhmI9MtzcYLV1B+XCqImRlyj/53FpxzhcRwxXWdrnBtPcEIoR4ggqsmeVvl67xbpy1BRmvc
9cFttvtTo6fCF//sU+bCQhiZBePmik+x9Q/R2Zv3C5vNr5ABGirBT5ru/56VJSIXYaAk5JNlimO0
YnLmJWXG/THx1eZZFcsVz4CM/GqsasBXva8W/K2sG9nNT/G0HwJtjs5HaJdrLzELTD+Tm1rNULzF
Ajr+efF+hLIpDSX8N2heaLo7ZnLHFG3UIRmNZnTLWDtCFZgWzzV+sqolEFZIiOI0fgqvADian6dK
E8UI6jL2Mqd/fZs6dsY0LpdAbVoNN1QXA8oyHYcVCVWsr266p19oy+lQ5l54wddIa4Bs0p9gEUYn
57upyefPh0OT1J00CT3wBkNusgMECIx8BYdfZxjEjlgMg8oEkoCgnDZOJsLlgOFZhEt8Fm8JOwFJ
texB22lX91MLYc2+TbZ5/ZSk5+p8QmmgdrHjf+8nf+TDt5MF7ZGsx73of4AZFXxaGuLCwWabHTtT
NdZd/1THZgJgu7jvKwOv3J2ctppXavVUNgY+PueI6yXUu3oAvfemBax6B913rvFB9d6/jiD11RCu
peIc0w9THd8jIS46AMkmZqTU6IiEKdyEHiIK5iRo5xW04gEiqMaPnqv/ouelNinE9mSXa1Uiwki2
lGn1UOoLsJ+R5kyD8AwR7MjgGeM8SWK2vtfCry+tlVVfXauZ6h6rdkJC61RLYAWhi5uaGO6Xc7l3
Bc0a+2tyLQKD9i4OKhT54xhgTuh30a3uC4pHRsOJq0itPZm4mTuW4c37taRK4lJgEbaYDYnjlxlk
iG87DGWsGYsHzkv0ElLB7m2ZDtv4DzxPOhXTnq5CZ8eSJtfG3yXRblB2bPVvLNrDyuFvi98hN3Gj
UDuDTDBH1arD25DbTPWdOMgQ4PcGUk5zLBZ551VGnFVwnVkiOEL7ECiXm69wQPClfRjK97E/oPod
bWgERzxweEjqK8zKuHruMx0XOoIFgregYIYVjLEAoVZfP74ER4DEPixuMTM3oMm59NuInFhfuoUr
gdruOZPtOj4L46KOksmzbzuM/VhPr15yHiNUY1iMWiFIdDfldB3KUPNOKB+N0h2bn1Zrs8kl8YjR
a6JP+iNsF2UZggI6cu8/nVPmHU9E3D+qaRDhkuM3YM2sSvPp/bR1BbB3ltzAxKHI0jAu66pFt21W
UPJNqhmW7Nuphf34fgXxY9kcf5YP3MEEY5+dyEnGyaox3YD/BBEWbvBG8OzM7b8WTclw/xxqtn0o
Co1NRIGqcYdA7gJkWr+4mSGsTKFOX9x30WbZJCGIQkEPLlU9Vm/NglXlphvrDvQkh1j/9AgvMILt
wrGC3kXn3URKgXFcSI6VRN8qGVHBLoFHNc0ndJNqvYSBSc9uwE1WLYGcpOs2po9oYfymIbT8AZAQ
Qhij0Peea6dybbSBd1A3Z5VIvU8bM7aJ2QxE49DxKo4Dlu9yT2CHYMs6v9DZETixJiwSYeyWXOWc
Uvgpg9BsbwtVWWqxXVKGF9CM85HKjdiVVS604jCWDuy4sgqwu1OqqJQ3Jekb5/XPKUQr5zcV67Rw
JOoFKSoW1eqZFoDUDO50Ck8rjsNXq7fyw3meQznh0hs9MtKKe8t5EEOmSrBBHYYaXbPEPwgvivlJ
8Op+Zt+YnPW/U5MxMGThHfZNEPGH0Onqg1W90zGXkIe/5cc4pj8hTSEMSa7KTzwBIvtJQFdL/J0O
suXlHCL0r5QLhPD27wCuTWRkPTV0qm9F3BC8HtTLxZfbfDIwwhFBxS+g+Ngu0hXdx5ncJeNU2nGB
UIjuImipesVZDBchOw0YGEXiHKO86etbcABahkoR5Tpl1MT/Y/BKI0e7+rdde6rwLaUrMIH7+QrX
8FaiTNb/DMtWV7inPPKCfMjKJBkGzOwhkqsCMB83HMHTG5bwAqnA0eGyfRt3u4nflU8iq8WJjf4Z
HDJ+y3PRykp6FvCfBoC1XtsfIxtxJPvuKi1tGzrAVRB+tsJkGpPcNpn1ku1X4PUFOW/bGp9cj4SH
zoqpfAKMLZbQ4rBdiUZOOu2KbW93b9zMHwud2ccWSZqpEEQVu9R7JtIsEt/QVutJRz2vXNX4vd3i
vDSoHNe3BraRP4TUTA5VZ2fxiokH3c/IPQv0/0uKMEKiHYgnnxxiuBn638zfoTXPeN+g3K2Z9u2U
SuQujw1vqdklLSOdwNhBc7/kj3IkPWKJS2HD+rGg5edYXi/zL3Qznu4OIZxt9OqlNCB0caaes9Q0
rzqEUtYnYzpvfI5ryMOR5qvYe+c4b4dd+sDy0pMzn3rhjk+XNm1PH+CtWj4oqYMPT4Fe54C5AXBB
v4sWLze8oyoiB3kv+iCHHvo4AdiI8ZrG6XY4CenfhCdrVxaY/1d+yxy6uq+p2EEIk62Ibvdm93CC
6ueIDiqt/nxMtElNFaOSOUcOvWXqSzK4JEZ0ceN66UxQFXfRB7unbEoAAs0Ixa8yl7LDpXXU2R7g
Md3ih32x/AzGNICtD2CQK9+uGvyVJ3lHEsVpw+T3mXf/2QiTsVre+co7pMJovcbIWSvKjChgHo5p
Xnj6EHnhkyvTp2ukbLyWeJkd/PX6FvhpXsH8OjDaXFtr6ftThwltJY0ywHwe/Uw79X+oAo9Pqtai
T1iuLpkf7G7G/cXwEjG0TE8IrNaH80gQsphIvd9s9wld6biqX3VS5WHxM7Kw0uZEK/ueD954YfcK
CDxoTSn0PKWorM3Cg+NyWnOgEsCFfj5qRX52dpl61IS1Rpbih5dC2gMh3suzazsvxyeSeVDGbdBO
RieRYY3HO6bQUaQ3GsXFeb1QNJJGt0QrOacaKFjMZKlDLyHU+Or3f9SdYHlOX3F1HmTak6AKBi7Y
oisFJorO0Sh1WfXXzEfTb9iG/rJaADq8nZPyIr1Cniv4E/HuLcSA6AwJHT+cjKPGF+DdM4+/yMRN
zFqh66kvSRHTxSx/NfmlGRHHf6Bc5QBr4Krmyfw7vqaqGk2DhUlpombstYXhtIPBgybEpsy8eM6r
RiNw+7pO4a9quJ+eRpWLm/k/ubKU3PNDgBBL3soq8OkGrzepTrUolkeNq4ByPS6m9uaG4+fLCqfi
dEjoVfFdu3uGVxIluUU1SYdyh4svth8SrbXl4bgRuJBIDio6x2JRJEs/LhOaSI0C6uaiaS50W262
o10T3y8aUpAmPWU6O/ATY83YKFh5Ux3FpJ3zup5xlHg47EbUqQ9oaPJrbSHAUWKsQ/1qzQouCRKD
auQguzx+en+8ywbRl69AyNwKf48V+qte9A9+txPeIlW/lsXNfb2TTgwB6V54WfaAj/LefbQSzizi
73Is8Q0Fi0wY127V2ExsH4Lzht7q60l6nf+oeY0VgeHotxpBvDUolVBrN7OXR6guw7SkvMaHpEry
P9M8+us3CmOoexdPjVYLufU9OMkLdTVQ9URFxlnwnxKSZxep/m5AYz4FEi73Fe1Xeo8thjxH1g9f
JVeEISFhjPYr78iZ5xcrJ0gujpDZmL3fX3GmwBYM6x8pTiFY33C/BZFr6zQO3Yow+qEoY/5orlRK
5pxr01tCyH8HMzp5iMj+Luewc66DTMdFgeq+vsy4N3iXJVplWoHEbt0OVeymhyfWNTA1BfSmFz2R
D6XUfiZ3KzD9H/jKwhmxv8CxDgrGUkMswPJ9WrUDzwhiVgL/hOsSW1BIzSdvxADVrTaYZWvrTaed
jtOzhhfofxzudK0r5KXrusljyzvzMQJ2rhbxpygwMEIaeXyX7hO+ehYXURH8YP7KpQXNjZn5S91p
k/Frhe65rRdPJQV10TnCDKnRjzDVjD2VSvFsMq3hAavN5KT0QmVLZ3m/Nxtqw9M6+eRU60rXu0zI
5HuK3LEhh1vER0K9AILNuzVGfZgUeCZvGtz7iUKJKc6kPd/tpj9zhMcKZycV0qVUfbvQcQWeSg7h
18TnGYO7+UMtNX7JSBQV+71wglx5OygOpBHovj5fU1xN+Cwt7GMnmuFsfJNawpnGIivXELcSfLUs
1Y55YLgYiqSoh1Gkn8BDRx2K2WMKooCIc4Na5q7AFgTGLhkUtoqJTdiTnFT4r45ft2sycdpvb60E
ScpFeggU8P5ZLbBuuMBGXQraV30gMoe0NFaSICxtdujrVaY8GKNnVV99GLSGaLBnumS1TU9tlnRV
LKxUN4E9bLuNWJxQdLK4bKcwQCO7OE1CWXmgu/JJqqp9OAN5gSHQdmbH5oafcTwCa9DT8m2sU7Nj
ocRpzHYRnnYPuCfAnlAt4+BdinOKpvP9LaZDT5N0OazPt1xxaxJRAU596eIAse792vsYKAEidCvK
XlfVy/ebsCChhqx8whazcbyvl4AppQ2mcpOg/0kSyLPQxBP8KPiUfM92LkfwJ6JikoMfNAC4I2P+
FkodT7pjBHpEraDWSE4UjWgpvyxLZupeUxC93kAuGt+Qv+PT+Y1kMShABtBpbA0qbzujfEV1vR1O
sQ2slh7mxy+7bvYZO0kaM9fMWBvN/ZtuL5Ca0f/97i8+MWcyk54XfhvGbv5/bQNEZO2FHHjjGZM2
LrOyTeNZXoEfeVsvFHYbr3N+MB8JZ3Zjt6ZEbsJS30vMUf0ITKEQznElLJGvB8bY2Kiejkt4i7KA
8zvHPpcqAsFVW66K/tuJZ5B/B+l7csaB6TuEumBXllRYB1flsjh/EkR8ONtgKmGy3ik2XIz3JCAO
OF5uUyYjTb8g6v7sYqWO7zMpm/52rQDtd4N2NKj+wWiOUyHrSxtqJ27/EAC2sEqJ1001Bi7uWoi2
yFtlvhclvEaBxzwKFAKppKfrHKHWkyyOJlAPf8zOA6ifyd8rsnQT6+JPeNtIpIPzOwUFnslehdSW
cg7a3tLgaMtfPY2PleZUzWkALpZCh/kvasvvfQ4Z00gOXfB56Dwlvgz726BJdAi3/6dHSDYbc/FH
y+xs5dMFZLs/vt14kD7uCUqrrOd1ULzJv1kY9BWnsK90354xaPmLfP+bOp7XOAOhsYASnrI6dQKn
UVmpoiMP69O2fiq7wyvf/4dUj1uJdRGrSI4dCS6LmacD18zfDJA/EYhaYFJ6aE/cf5VLqOU4l2bD
/QiReYhannZ6HC1k5JUa9V3XJbmJFGpLA22KC4bjQK1Y7H9ittDLt4XISguuM+gk9WCU0lg2NQzO
r+XccbbmyN/w9eTRw8bTSJ71PdyEJaPG/mooBfAv1FZq2s5+h2miJ/j+LQODjYDy65D24lMqrYuh
Dvj5FPSiuOWSCcrY48o560d57JOnvavPWuaObz2uVNSuYAUVCM134iFS0RLf1Km2qFDvcxBH5mpq
7VFOExlFyuwStIGIrzU8A7t0B6oRmmZelbq/H0kIf8ptZE47MxSaVl8lvJu3dR/sXro3r9rqqKUo
7iojHAhwOAA6yRIrM2NENYuStFIvyTP+911yoTIBiGwKE5iEnqppGua3/qV2hl+0jRgXwWjtU1nx
VfD0z7qMFEUub4krYSayL+EYWQsupJzu1mwBLQr8+GDB05He2q2dxo3Gw9MQJ28GRzq3o6MbCReY
QQX1xM4mz0lSXCw8MGK4k1VjnFzIQHiOxJeYmJFeC8vkHhB128miPUVNZiCqR/mVaNkvx2TfL3Ek
hzgLmM7b0K+DNn9h9DhVsJ1Hu/pJ3da+lWWxGVcU/iD9/3xrmQ4hf3IIAZVhvpvaymEpSxJiABEV
yqxUXO0hx5SgD3DnxVHpHx6xNCONZm05YiHeFih41c1AqP4ZynDoDxHaGZuKo3Vd+4qVB/0f3m2o
wIEXswgOav5Pay5ZQcNQgNXkvj1W7+o6lBv94KL+krOePKqaYVlfIKHHq6fElrOgRAhuUEDOmRmE
CrxeuHoVu1TL9wCjkoXZPDlkGDN9tzR0U6nFBm2ZXLCgZfAGhl13s1rxTU7n0uLRgkS+gfQlcrJj
LuNwxBPzaZY5BbBBeGNUM20LFSoshEEfvWbYGLt/qBRQxvJUITBHj5FqJlb6P5Nwv+us8+lSgaot
hQcX0UZbKXkByuejK54S1tyBXCDE0OW6TFQMGl9MExUFx7rB0CccK2jddbO1YMLh4yJ9vV1yUKL+
NRN3dZpjPeoyOF0goWNBLfK0aDS8BimJAEyONJuwQVal2Pw58BHkfiE/izCetWkdYRVE4mrNaRpX
3MaPqMwrjWRPcbGX49Ew/xp+fvdx9nV/PL500kvj0mF8kXHn0EdkHNr9Bgm+4MeVEMW8PAtFXSNn
GSuPRZvIVbg9003vqBfUl9CsLEVPJkYsPooo0f0MP+3mDBLQD8GTW9R5rHylFDAcPs6k79yKaTsd
LdjBkh0M5DgaLcvkeK92yM3OH6olx4d+OTGd5o2C4vXn1gt9qyzPdbBRl8BvrHDg/5Z9J09MQf+A
UAEISAS0IGoFO8T6lUDaRAUtzmcPCP2qKS8VbRpckwnnC2FlwHj/glQB8rtNXGby6VWICtiFQ2NZ
IiaP5D4RfDbyoHymsJVAbbwKv7ruLzTRXB7FTiBT0v+NFHwZ9HqZqcCaRuNA1DQ6ho0wJkR05A9p
KzaIXf0RvTHlcA+VSIYxoH4kRDSb4PGCcAEJa5dnxYdMJmy0ctjn38F26Y13PQCWkGYY8v+hxcOO
FGxmhZ03kNJuHNHDoS0CK2uU+kfIlaAdBPBBJevT7K/6DKnpcpQiFuTTVy2geK82jejhXzS6ENA2
EgDkGxkXlDFk6QQmccirrzvz+2AvB7o0vkQcmamNFfOMc/AfGGDYXtej4QcgPUzhbRG/VUURNOFq
4zO/SKifbJSHWuknHFN0WmDe5MDRp/gz3bMayeXrn3qSQrq8Zu3KZyN9Ki1Hv4570wNGbSaiouVn
QdmkiOjCfQUEu858jdf69nqXU61YHHKeO4CXW0NNP48RH2sPu6M84WIMiUFOHABdIVOINwvC9gz4
Al0d1w9BTV8SEiuD3kZtP2PX7Ff9fCwlkg98a1Yz+vVDvQReOnuVfT5kK28L7TXrLCbHAVp6aqhj
PvRNgutxYM/AeAj4LHF2Xq9+PrZM5Z4btZloNl48ZQCYw+11tl1cYJtBa7lLHALs9W9dzUS7SH/P
0WcAAT1JL6SYqBU7leB22Dlf3f2zFFzpzGBB1lA7L5YUaU/e4y1Nfw7ZMInJEFVj0pBiAAhHCD5q
sQQLHNRijrtJ1/0xuF+fp7/ktzYQ2RECW+dGvZIBP/m7UhZQv9bsunaPbeFmk66THaa9ik8X8Tgn
11VE103g0O2BmHQcSeJOBbzobmca4bgF77hb+Bhg8N9AQ+VePM03UQrcCOCZQ3xAkx2NGEUWJ+0M
GPNQ+HpL48AoqpPIbAkwkRt7rsKYJ86ooAN0GKM0EIYAEJwr9Xd+579wui/ek+e5IGaVWxJ4RBHw
NHHQqITpVBQ3OHYa+1Wf0EuIDyEDx5/17Gft/40O2B0Dv4z7PZONJ/g4vu+hVcLAebQSKRHJjBnp
OsGBgqst+nSjlcDbA2k8aYbuuV0tjVK+0AbHosPsI/A6Cur6dDwABZHYzwPbWPfyIm30IzuhMZsZ
VEtWdL9E1ubX0SPhoOZQcfF1/9AvSLSdE6C7nw4gMJ+hd4HjmQTYPsIgO302oR3pjEcZaGBpzq0O
dYA/aCuYQ5PZ3By1sdLaeWJZx5D3XoNuq3uCq6+DLdn/WcJ2bTSZ4azGjLUaHLqB//6GH1Yi3qiG
OL4sm/PEhxJkty6Q/RB8SmSe9eMe148/4ihRzKcbAFpTSrkSADPSrTByugj35eMkHzSszSEDnFm8
gay7GzmuLCH7s3R+nhXRyTGD5XZWStWSyJTCZth50CNNzglXbCFnOUyHF05yyrcyTrATX397wBwO
AWJOikPPjpz8BgUg8ZA5jsscK8KtMYe8gJzDDXT3901nTRLpnHI/0I8oeLXoKVUmLjUOB0WaQf/+
TuJjA/EwiLqivglrjywDeHPFvZzW0tC9ocBh51eat1wlXu5+7pV7g+kVfORfWPuI84CN7GLkIivp
eQvo7VnYpVvmdGMcLQ1vXgKxsUGtQcGyJZxmK1sMcxma/tL62LItsc2CHgY4WtszlAABdU4CvYkB
9wkMWcIDvVkuquBHTbVmLVJrppmyGYZjLAUZJUWqwy5m5ugtUULodWw7oto5AWrKmRL2JQ7vi4CW
E9ntQNfHUmRwY/qS2nu/d64THZj4Sq4KPdHhgZHPqM6qQkAUz2uzIHbbpZ6e4eF386aQMf10skrR
sSPom5vXIiou6bi6tfDrFGXHAFbblW+2DrlMvEBLLYHoYbkwKnblDI3Usi5AGFMUgdXLnVrmlvkS
09N+6n+ZhPqmy3BZUdD/UzgeNCLVUZ8Wk5zwvqRZE5+TRl9uqulL2jFXMqLrHDUBwYkcKbguq/jh
ql6pSvGdGyHlZFum8zTMrCxXDm7p8+4sTW1ah4tPEv9HKtPZXbmSO88M+Oq9kHCXfAOKsxxkb2W3
qA3LOTPUI/5ILK5rMMS7UzFvvzEtWBqRzUKTokHDZfqc8S8sD9RjqPX23AeNoLdVsbQTV/jFd7Qu
qJhoFVLMdOEjmtXvYzesJ42HiiDwpFpu6xlx0r0H5QSK58ruxdSqd6bUwpItZaI0tkSWkdurL/ln
sv74aISjzyuxNZ7YeCqYGHYm7mCj6cI91jCk/AAqVh4hdKqonukg5Zl4K2N4CyEJxzNdc1fjKwK1
KzaukyXXIeU/NMtoNa36MfvRg+OEc2CMEIeaNp4aDdXUYyBNF/dDHj6SZRJ71TjZMf2IvFFPSHzV
0MlwiXWDQkNdRPUhdYHpnHwxuEXD8TWxLpJSjKmGzalksTnGkkJwfpnWNi0E897oCeDvqh1rkVq0
bCGkbtrpWrEaIM4OGSqkex2bQ66a2CaKG3k5NahboCFZTRpndfWkuemdtMs+Mr+Yqm1+lykLpqHk
yB/1U/PFQC5peDtVjcnMeIh/VE4yRBbvmgS0h04593Q1SB+SzoHart2pqgeJ3KTqlLozaYSarQjy
KF5CwFcG11T0OHb2WT/di8V8hGfgD/go857STxVUxwsFfPci4Nnf/0fnaVuzAhS1opCcSIBOEOeL
eKA8z63IgzXyDIg+i0ct/XysjVhil4imZ6ZwXCFE9YGOgloYob4yg5VJXhcUaVq1p9D8Z3SbubZ9
wr9h3Kpkd/1vKGiwSFgnlkijE9HBmuqrNbtF1+oXrlx+YbZXnaS7tyDyZyqpdE4uN2c9SHcuSRLz
0voO9/1UPXayhCJmQBKSniSRhrF0lZNdmiYNCJe/WGHNmJEeUrm4O8yQdfg1/G9Hxir2gALOFER5
J28FrDysNp3NFRGhGazvl9+ILILKPhYEjlPbM0b5kDdQVucnefMEIUOrEeanX1lR3gW1TUy/O8Wj
2ETGrBI7JpVJddQpBNz9z0XL1R9OO5sTW29Z3btbg++kmQHw8no5hgajuS6lUeS5Jo+d1QrLpNYq
jN+Mss2ndE10VmIWbHOlyw436H1sLW05zPVM/09pkLhcGsSP+jaKD8hC2nlhpAjJFLO8xlMbDwQd
GsEkOjU+3Xk0Kl/ddPJIp6cgcSxd9Z6XvT4vxhlTswbvez3AiZ6wiCGctHE/FF2oc9BIDryk/0Id
f+dBEoQuq1ShzWVO4JDBxOIDPlq8Q20FWLL4HhMM/51QdIjBQvlY4t/DvHU3gffnrhrvEVZaTvKt
+GkJ5n7Wh14FqChQO210EpxIvddaQZ/ICAxy7GMOJOnQrnZ0mXT3xypm1MeBL97LKbiKtBD57W73
IET3ZTuERt5SR4Irqt2iiSzwE4q1fJQFWN7hy9MmVDI7A6z6jizqPLhdil1G12Se/LOP4d/Tr0DG
nyqAjNu9W+UvuBsE73c1K8evQmnNRI3Mj+4Kiwvk4tORe1kyryqs5ZtcCkEOCyCAk+UTk17QKw0k
6eTH6Q0FQscRrz55KnqUlxLXotgQfw7qD7BlblIGSLP3Z0tSJCfKfSgqoynAZyhmZFAAPwfAbAjX
7bK2wCnVum1rRwt+j5UES0ETSlqSm4S+TqFHZC4D2wKWx56UzSXQ7SgaxwIDwcXlvHQT9TOZHMg8
cFh1K9U5vzHG8xM7RyYGcYt+NcAYxGjmf3sVfTIrUjWf1JfZZYya/IvKZmzO0BBpxjA9XSd3XdpU
WkSBLMAGFiqw/PFoSWzMR5blLa2CSDDA7oaGNKbWmP1sIc1criCChc2TFxgelYK6Ld+B0fcVAylI
MKhYOMKvnCZQP9sQWCkUNs/UA58dHxqzZdCAqiXF39TBGhEmZQnhaJoZfn9T6I8tomvT6XL62VR7
auq/yHxVGbai3Uo/VJ5rJrGd/YFIbuFWET7WfAc/2zEKVSnY2lgSWda5sn/iA9EXRpW8EDixsDkf
zL3CmzkU0r1di5W4e1lEiP50wTYJR0ygEw5GMvEhwS1tOwEgRqJDskH1/DNV88vzVmO/GH8YWYFu
igOdZ8MlOYWX1PpdoMFpRSXIEapWneVx9AAYqkrQN2E9h8JsrrNOitMUNt9pO3ZgnTcLQMwTKItQ
S2+cTFOIfHQJ/Ptma0RWhN8+O9bYj70wz5gyljojoPefCHucPHnQ7SGTdpPbIWjdTUZO7sbGZn8R
WGn6SClUM9LuRSz80w9oPNTaIZ/iGDezWNmdSFnTxtLIoQj7Pv8Vk/fDHjXALQ0pSCU7P34qVqzB
pPZtpkYfwdyomRyiO39Kxh/HqTh3HCpilZ5ZCRKi9A0PqGpYvCXuDjbftCqZlb1nWYcNWGxFay5j
OqvJL/o2WWEHKfQmFs0Ey+Y1f7KTUR6pEbUWN83BwdZbMUN0/wtwGDGqPbXusojU6rvKctGB0cSW
ahvly8/+zPoTtbS7fI/NioOMgAqm7GPOJYuDK+CBN9M8JMtvqjwcmp2m4SkMIsgDij5f8WWoqpZc
DfqywBGYKd/v7ZJKEJwAHK280rEWYPxpin01cEEgyTZt9KCC6j10O4I7cH0KBym1gFBOUpaoRDgZ
6BWD5SDA92EqHh7q2x1dCY6trsG32dKhVGGBgIp1hDXQQt+2OQjUC+0thZ9a2gOBtI8s7pl0J9Z3
m7klURQTNUI349OjNrdi0Hp4jRcNSUqiRdaPrD6ahUIsklWMpqGFvfnms7VHOcqyXSY7ipKG+U5R
vcwmHI5GAqDDGgo0tjgukiO0JgKTrznIXaxBYWYRfZ1F2CLbg1xggQ+U/QAcHv4lGnRQaLGcDvbr
VXBQ2ozSWG3VdgnBqi/h+4bIbKPYlqVcK+GofXCHQQKszBxT1GyiOz6HdwCQejKS9Lr3KAbh4FCZ
UvwI2q/7QpWLEsM44K/raEAu3UgekbmRU849OKibIuoe1BiAixyumjwgquFFW3e4iuGvlcC0qAbU
AqipCCq/4QyRasGGNiyNbSpkib+pyBQ/zmQYE5XYEtICM5lnWJLmesKQC742DlBTVNI1NaCSRGQ8
xtNDF3lowoYLZF5kO/goYfhS5me3sdkwt0Gd3aP3s9FZ6w0hN3W56c8dfSBIDB4CtP2/Q9U5Z5Aa
QExz1TQEEoe+1UX/5NlvSPcEHrZVlY6OnGhHpxsjXGcX+d4yZt6Ze6rsJrM33otlwGDCwOy5J01J
mt9TWirviIk+zzYs1X9DojJCvllOwRNHTp+bRfj+mPGa9acu5JQPnibH60kie6dOJ5VVcLYKJN3Q
hfYGOmYZHjMfFHcGdFwBLkkSyTcvVu1gbjuOAnMc0LqaGnUGIyFBIC/6N1rYEktfBxl43JbrhZtc
AvgYHzBYyzvyiHw76LwO6F2v8iFvJ+BbgUTFda6n5/qoD5xcfv1plGlSuFpwRrFwdhIsU66cR6ne
O03C1NbEP5k1NcVIpcN6pva5xumvYX7Cxd4p43Uf+5eBxqgYe6+BGb11fpCunyH+sqrtg9yWS7Sl
1A1QelAm8E+5CPbAN5aoNn0yKff2OsPjSOfhY5FUmNVEO8MoNsQ7T479Qsx31IrHTvyRLMj0V3FX
B45dslrj7TNbeeZCl7SBLsnqR7i6P0NoMUAC8GhFcbbxjCxJQzVX9Kp+y1w2kQyI1ueQEbHpYF/T
f0ZtHJPJ7IoxppdnwhnTPWF7ffcIl+qxiHfws4y905Og7hFiQFVQxiPWdUEpkJGFO5BM+eD5W4/D
Cge1BHMLIZO35PGhQX98u1VldWiqpiRgdMw0soTeKFkkCX1XOUjBOYZeJsM2WkPVM0WFQhgm2YJH
Om1E/p+HIauVPWu/Ag6GgsR1taIhpbkApa7QMngJxXuh0RvG1bFnyJ/zewVkitFsbgXcJpMnshqd
xD3DRIcgdsk77PnAbimfZJh8IlxJDMji2TIEqz7v3NLJErO1LOU6y1dZj/TAO0X59dVmbsfS/H9E
tBp03HQnSw831DT7nBaBx5Wlm7jcC3UEI3OBHgvtbN0joEB9At6NnSYoQZxhJa5/1nUoYUOODpyc
ulbDOaeIq7NHC+zRtsRNBWUEny691OapMHWm6g+UUvZTKLaVr5+wcYwbd7z2l9fngkRpi+KgoDjq
HBNCPe2libtEdStq0F293fQcRA8OBdt2sPpOZGYgc+cxtpfpD/Toj92zKK3HpPixa8jj2mwZQRHs
IJJwnlf7SRpr1qu+aGEXHwHUyRUZTBHuTAhFHnVNYeXhN3oa9su4t9fwdfJjN6RoworoCW4QRC57
4dMq9vhL9UkUPrD4iIyyG88l5dVV+/gZxM2m/VJiIhEROpa9cxDMwu4IXvyA499uLBEjXzqZjPsC
41KeOFSEbdTjMuT7JNv9rQUulqTeFvua50BhhIFtq2112GP3ToUPHkdHZDqudRftT4s/CE8rwWcE
YNj0smdlJ+riskgLDbp6BO95lcUejZWgqpMsvpVg2GOgwViFp1151HPYiinxd2cDB42Pz+RaCpg2
Rc+CDZ+GKCb/OJJF9s/qKtxQz8OlIx79C1BEcuKwoxf0eVZBS9ErqK8QiLxcvzXHWfMl6zI1HVA4
6BY1qvAAEd72Drzp6+sBciTvgLEdcRKBdpPQ7vgWKk07FQBMyxVMQwZDNLRY1PH9dyB7a15q5sbs
8lw6TX+dzIAiuHi70gcSjbBkmnhsH0OKGAhz6C2fBo2LHfaskk+NcOgVcY0wJZSj1SGx/U1EZBi5
9foawbVQuPy4piWgs1d2w0enQ9SRsUKzn5t7OT9hYuNw8UgpkMfH5CudP5AE/n+GYoMp79auA+5A
eBnFNdY14Ziqnn+AJCjM4dy7goy2kRv8HjmKuQBl32U3Lpj9jcu2Uk5Y8GnA3vXNM23JRq7fdBFP
LZtpOUphzke2yHuBfHbCBM3hEQARIDgfYw==
`pragma protect end_protected
