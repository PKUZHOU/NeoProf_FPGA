// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
os5PeKtmP59uqtFdLJip1SFvsJFgi4x4D4NntqGY3auyuTdsXlr1bVkvKJquKg1D
nuSvI3szRfYnpgTRwOXHRYJ/ZYuTqQSg84mw5IHaM6PYUvmY3RTWQyBnSSmxrCkY
FLEqUzKYh0TaEygDi6sYt11Fv7zL6I9kaFuLzVn/P9iha/hC4KUj+A==
//pragma protect end_key_block
//pragma protect digest_block
IG09vV2J9m/DM1hPBD9BOyH5DBM=
//pragma protect end_digest_block
//pragma protect data_block
REo1DedvE6tRj5TK4yB+TpSdfexnun69lcgLy31oOi6keGpT7vjwAmQVDcJmHbAy
U/L4cA3HFbJ46awivoGCdchzI2CCbcF+jQ6H5EuC2aZfGfMM7ePgZEE9Am9mpWdb
TMichOnYnRv1gu1ZsRbWsgmLV7qqTM8NA59Wm4jyIdqrPDCl7ol6rPR9J+GH1bht
zaNCq0qcemGpol66MKBDHWmYoocAs3OzFn1sx4xz3k08yo2HiC8c2GqYubDvsl83
oG52uFyn92Z4eBfARJaYKUUNmbGIy2KUk2EQJ0naEc8Khr8q5OL+V3Y7/Sm3DyJX
VENtXJKpl8eLGJMOaipKOtiePds2PsVBzkmWkV+ODd7/e1hLndcS/m7zFJeS5w8L
eNFojQg2KLLkhdIQ0foK/kF37/ANQ9kyIaq7Zc/WUGBnlG/kjFgfRQ9D3yWhWAT7
3Zx/A253NlTrt3KmoZgalHj4z2pPLWykTF66bYxWCyOS9l2oDGKXuBTlh66iqU19
o8Sn2ic2kZeINlbdjbbIK7F5fNxbcS+cS/dJhoNjOavNplV/9LanU2/eMXL4i3Uf
xdAnyjL31PffHEb2JyNYwE0k2JssZ9TfJ+Fx8O/kUANEI4pFAFcKJclk/LZhGxmm
7NihXqlvfIe0YEfU4ykVnXB36ZFhhaNjVFz1O15qq/f6tXzGK7xc1pm++B8HBOX+
qpnlz/S4kYDI9cghUHqfHWAaVA283I8QVbVae/rW7edEeWrk1/jdiejrbS632tmn
q6IPey9hsY6dtqlvvCugQiCYyPAcEqa4439eaTSZfdNbFozXYVbNSJrIKdncYn+C
hs/EPbPBmQ84ufwM4b0VjmytfzXE7pY9UxkonX927ukVza8m9QAy1K7f6jgWECmT
IjDXLMxaIJjjyFkEclcyU62oTkLsmMIZ2WrY40AJlaB4RatC6EQ8tMpUWcU+zE/9
qhlOpwP9vT3QRbmzHbCA4bh9rhb9mjIOO6wbnk9uN+I6XnhI/qqfQoYSRzhFmQ5T
XSXNn7PWiiAHchf3eIuXQMFIr3N4HfV6AFWT7Bbwz61wI8a45aaVKepahDO9muhT
lh8F0Ky2WNnNNQ6PV4iyNZlUjLCW4MJvNNOlet1SzSe5mRCqkhbYJUeBvnlIu0s3
4pzPU23OdNt9PiEAUNIk2eiNWDdnBqCK9fOqFdO6DolLPQ4EiJz4qkGTBT+NB/en
5/dufHRh6/q2alwwh8bKKHel/IUHsCbqoHR4zh5NpN6VTXEvvZf6Z3SKmxMljIAU
xbST48wFHUh0mA/6K7ZsPc6e2jvjuy/MME3j9nDOviPKSagjYZiraC/rDq1StYjp
2pp/joivGYbNMP5tLc4RpI/XZ0ZFEFZwFvngCVdhoSo8JlApKB6jSESOrYM0z2Wg
LjD0LtIyD9VRZGkybPeVq7rebLJcaSY2ZunSoalo6BsBw46vppTidjlPq5rjY5vg
LqQZjaKlqvRwIIDQsEteTw28uGAnFvcWv0HxfA47q2aTC2nvBmDRLit9ZfG/092x
eCWwXpYkvDBBM6eZBk9SDBwMxfcuf6jsaKuYvzXBiqGVvIjrHcWxxLjqR0wkdcVz
fS7TjowpWQSiyVuxuknnXKAuiRImreG/g5QogPWKvRdaSNEhCcWs8/89XdgENiwu
91kXw/+HeT07cbV6XhrPOitlLRpO293zcYttTsCk0IM5r8VOoSg6H30WKcdYl0Hn
NdYUtcwbOU2UHUgsCEZ0IzXhzk6swBvFePopQxuE+WM3rrrjaWPyA+SKWlVkbmmX
r2+vNZDGTXjVpmyNNt6w6ThzeI9dV6qDCnehtfbkcDQsCsT7iwnHgLo2xRJftQ3X
LCT/FeOhU+o9u9Gow3ye4NJZ1lyCOr06Wnn2bgRwSYcH9XxxBypYCh85Dm6asMuj
rVMDyYXZQtTG+y2jHzWAzj++FLdzyZcoACvr+fK63AZSQ1kbTI3sCAh9wcrYwhyS
A9s88+farifocS4w/K/HECujzgwI+0c3AnLIEliiDD1Aw/OGRk4NG2h9FmRi6QG/
15Yx45gFgiq7igFaqdxPyAgRmw7YMaR9P/AWuF1misyaXOe5uwquFL4yutb3Jqjj
uPl5sSSscVNKGtwo+QJCEhip5HmJOEjh1IWj3KCSV/0K2zFFqDyHPBFiVPNbQRWS
D9MkusIWkjblJNOEAomtjuMUzPwdC5S48CzNYpH7jgS2gozPAnFriW1GZfM3Abs5
PXIjRdD19elKIpGwRsoz4rTpqoNDqKT4QS/y6pK8fvLovXCSPLhsioXGeq4TPCM3
9HoXUVYAwhqDUNkyMbA7EvW4Z5eRBZRASoQL6hVFwyVL2YaxtHj4/3KrZcoNvFP9
DD6QTLuy9HpSlwOFsF7EBr0ilrJd36SF/QL7x+aq5vzg/8B76bYjGPBlyATX0dQ6
4a/DmisPpt3M2Ds1uVYPU+B+F0CtYZWGxuvPAUYLckDOtWBAkvZjGKqXZxw335VQ
nJzf4IOtUnWKE97+qCyPZO1JIYry2Lq7hHtvPrtRZPCeTYAoU19UFGdISNNFdKeo
+YJI7h1a4BMKPsY5Wyg/Wg3PY/YlgiO+uF+aAyTHHHy4goNV+55lKdniU9pizPoj
YcDPy2tiuV6KaZW7DXEM2z6N/2yWqRymFSsU5AUaBv5pk491Jq8O8cVM9m0dtp7p
+4oj20RU2mmvkKeDcFji1GgN5eZzSsq/SL4dtysSTRvjdeyAsGbrOGCjk6/t6C34
/uqhtYuQpQe3rlyAL9Z7az7m39fqtc6gar5FQ1sdX1ghtFKv6Plc09WWN4/ceIRE
NLNUtUorRZHQO+e9o1UlD8FjHiKkNyYx9dgykGlSWGTQDIXggi2idWsKG+zc9sdo
7J9nDCGEzsA7Aq9+y0uG5nO53VLAHNyiUtNb+BjRk+idjucEVkNv/cxXKFSQprIf
9Izzh2sf/8qqTgoTfYyvnPfOEu43e90Tm9ikvxifw9szfr4QVsMP1OB8q/Ebe7CL
ONLjHEqcBJtfsSdiyZah6vRPlLrRWx241T8y/5Izw6eTvobtkl/3jprdXt/1f8n7
gTtV9Twca+kxf+4wORlx6Ly4VnP+n+j9Q66XEy/ZgLZUXwfRWjAKzvObigrbdpBe
gVwy1YhAuC1DkYqgo4uySzAXgL7txOt5f+rlOFC1CB9UAb3AvDH4T//XTmKHJfV7
FM4EFPH/EIeHhbrj1FmDt4de3cQsyt1717NgvLkRZsE8pw9SObaJiNNK2K7Ol40l
0sO+PZJOyiWzmihmp4gPCnakvYd/q+t++ZI2eu9i+It6wA1yypyyw22WSm2Rjvjk
yjmw3pMtWPslpZKBBsU4Zg5xK6ANBWNIv66CAMDvfyvXkKE3QTTpAYy3g/ADcheB
tFVXlUtGJEEQxuyQlpMM7oASl9phlCwKVigXNercRvJPgUSql3dMeruKHzCFK/Rp
zENAXU/cfjV+6XSa0C8s05H/9RFgmzsciMZ4uPIZ8S2NDC2c/l8cxtEBMPccs/vc
A3EYgIwui75YbhI14bKzRvswKbK4oFJF4UYssFOuECQyedyio31lC4LXpVLdri8/
5CV/YSYjV1R+HD5R8lw1pHUIcMBVrjnmSfWDX5cFCScTpfOkb1Tb0R2fYKfJ5LvD
QGHWg63pTRFhzW5F454N6KuMLrdDTJYHF2mfAdNTfgKlGvXNOnsxKIJaiFJMV2Dc
eA1Xy0MSqVElnwgEMr5t4GYQU4ajMeByBLu5FqALnwlAxd34+XeLhhR1nQLllzgP
8KAIFqOugAMAm9Sc43OtXQET1j/nW6+RJ7usq5s4IXkVjb5AwPpbnkJGAttfjDUP
4HQwBXTVNYFjNZhVRdKgXRX2KLIJC76G/34jXPcG3PAvBkC/LmyrREEUHZgoKZ7s
UqMATCaY6vyQeSJm+z7UzL8U8XeDmgo9dyYDNackBOyIBfBHLmWLuTr1TpvM+kro
MatvZFmMUTMoE7FbbEKIfl0Orrdlz2WszF+K/3L7WYxkPeHmktvFzbxsBpDVVQV/
6RSpVzVahgF+DxFtlZQfZtuSGXFRxdT1Z3OhYubR3yHZaKFtqU0juVZJKONOMOcD
Ko/aI58X8btCFBe57zW2vi0wTJFOefVw0URAJ+NKEU8S36C+JAJVIcxo9NkhWqWY
e2HRqvWwS9YRk7/89qm0EqpQye4MeqodRbTZ198YpJhx4FTqxrTpQQ89XxjB1rxr
bUekxZ4at/tLuBFXbhj3iXbXV6+o/LyVWryaAi826KSjTrAaajEoRp2wq1EG1DaG
hnI5Ar88oVZ4crGpSzAf3WMbaMQj0v1f7Bea2iknX+qwh0KPiUQuzC/9naSkp2HJ
mXlKUEnfv0BxtW6e1a62et95SEjDuD16N8esuTqlFKTzbybEED9Khsm2jFa8BYTI
I8jI5JTNLGUjBuX+1aO9MGe4ANU8A4Ei1ACIvD7xV8u8fsbAg7IfKRRfy7HpUC6S
a6XREaG6RfhBsOFaWUMHZQ6LIgR+Qtip5xfmRdCXU5pIcRVFpdOoHUzej0GfxB1S
0ABCea8mU3xORf0IsCBJawis/xeraWRe06L1yqN7wqDxxLM3E2ePPgkVZFujJmAY
UqE8r12xlMNCiahUmmGldiF1NNETAjmTIHtGGZGkq+64UsOtDBFHXwU0d8VN9AYH
AUZJqjShcD8uKcJPGDNKJ/Q0mVl8n86gSgu2IapUvpe9LTJeX/mYZMVWGgdXLKxs
dRMkRFVYiGvCcN0pJ2wvIiXe3UCv4Sw87p3Xu8kw6LsrD0g8Uou7vakTtfCt4M28
L1nqkUpGNg9D3hfsLgkzCMn0Q3a2kmoomrbmv7vRt9hU00VdjDYhr8ZoMOnNT/0K
wMnM0YuqKGqmLr683/47xWzqav316FT62TCW7iVLIOjZQYp6BwTbNWt1DHwtS3cj
r02lhm4ZQ0NRIORwSiYDvpzeawB+C31rLUtR7sJk/mSuNfuqKKpCd64dKRt8LIn1
cxw+ipCLZ2ZjAv8lSkW1D3EBPzHxbm4ZJQ2lx/jS0KO3yMRBHNOf4ae5+sX5Aka5
/EaZIGKsFFnhclEol7QFVKwDeqHARjg0RP3WUKbfbxi0CNXjwHyUnJxg3o4jG+WU
Hy3CWbtKQ5NjEhbKxDbvPzpoXMSGtPdVNKNjgqWaU/tWHqKbL2Df48mQpUP4UyUw
GH2me7l4IOFaxGDqKnBM+pecLhJhqsp1/mu7y/DRXiid12co7CldTLOEQi7p8nyz
d9zh0gNUZvipcZSepTgF9pEfdN7TerPyTmKD1Jipj+Lkk6nnpFn6Ej7X10Txn5lf
ZHOy8UGsz9eoZNVjBJmZZK8mT8lNhKqCsLXz46P6Bc2by6aCQg7in8z2XITmBXH5
0O5N/SyBeK7/cd2r6GHhoQl6tNLLmEzvBTh9KXqDIeTEslTi2jY51v98cUKNR6Xh
4KQHOZlkP+AaLIsPGFb6gpZ0eLObvaB/KMf5NsAAPztwK/RKmheLzp1B/Ffos2Ix
VIy+ghyEBnbtssqLUInZKzzHwyr86Qye7a3dkgfJ27BlOFqkSgHgIQ8plW9VZ3Ua
niPl+Kz4NCmwlWbI7xPbkj/GX35dTmX1CDKhtGqX8EnA/YVFAFpTuh9jZxO2H0uS
/u/0ciKuNdN95Uf25UqU5se7tGi0owXoLjVY2I02ukSv/e5hSO50fVAb/uHvZlvl
ztOX2ZfiM73CU2sO9kQvSd7TypowvRn7sQG/dWcfGMOtgIQM8jk0NYqdg7OM7faw
IZ57V9XuBfIWpWZ4W4x+AJMOcYw7fC63679lpo7fatpwO9RFK9884gbuqKHE2//w
aSqx/XnF/EDYf1NwytHSfPa9i6NX+oMBJS+yWGQ5r4NQUczUPPIHmGZraiqMsALa
UAkZtPjf3BLHHqNrs0PJ8NbbFmSEnsQBZCQcv9N6Qwu098xVhaFAJc6C0Ts0qAoZ
jmCULTEe+2a/2xvfNGnErgaFH+bzOnMIPF1rFLk/NJONRBC4Gz2A6IKOVfpyh2+p
/c2Cqws8tXiz/CGaGwZlRNZTxpD/KNPZRNIbvXYtOjlpQl1hHlCIYeN5o9jtqZjR
u/2rdlca31x3MmoX9IjPjf2tKsDCo8D9gl0OmnCH3mc7Go3ZMiI0+5DSEp+WoeDF
AWkEuLNtUZgUPM45uTR/kCL1bteCGOo8F3ZJnYnNG7DIKJTenZscW48mx44N0lOk
otqFGV8iQRhWKRwgBsZnWQajekp+2ukeh5PWv5I2/emzXJnrJy529APcBHuE8Vtc
GrXS52a043lda65FoiywJJTxmagtLNooUbMqItKXuOBM3ey84jopEDqO5DxYNVhG
+nUZQLHSTKeAuMPhEJvTulaG3yffp0gb6czEAUGrh7uqccJsRbnxMKgoe/5LCDCe
qt5kOJB5wFMeZCzwfGFTpKH6j3jFJCZWDF21vxnFQCNP7wb/4+xNEtwiSOkkfrzC
fLcSYSAnpTQJDmB7Y1mzuSk6vNcToXdB8evJuc8VfGQZ+8WIQLlY3tsqlYzqmHvu
9qgx7Y3Mqjiey9f0a/rBXvGx9/UQLVoDPA1AawMQU8cR6LNxXzUNIW8h23bRz7DJ
8s60ZgKRihH3bwyrsYS8+I9OPsl1RP5N7njOQ2CwWMwrhQJh+DR/oP34+7y8rAJg
g7AWcvB8Z1HeR5wvBLiS50XdimmBhjq6HAnPgqFCba/oBUgFLV6FkCavG+/tu3a4
aXyniRW6T+LLz+JlPdkT11f7ybVlZV4c4d7HOn8V/OIUyzR2Arp+QwO5x0x5H6dP
uQUb7Y/ekJMiwQFekrEdkeWP8Yx1NhUqh5qskPPe9kjrNNqZFNeqz91QAkW/mSAy
rbQMpRNXrMClgnaqLVQWvkejgc8IcF9vlCz0NuB4ifIi1S5xNK4UYejpXxmGlMi3
7hCyp58UQsRLMtj4oiyC6I1GBT4mqMSy/meP9Mi4CYsuQjYaA00F94JBY9GRZa0v
pgUdwT8dKV86vf0OYHsQxQlifztJPcPcURECe+XQPNskCqdHR6kSWVuxtbXVI36q
OGe7UDHPWMYCyq9d/ycHqXHu8jf06P2ojzNkrEbP/05A4dF/pC7s9r8HFYkiOFth
M3VyxgCns9KOZxOWg+t+EKMD0C9Zv35VPi2A3X2mqhfehbpyodvaGOccR4+VLntG
RdctA5IPGGuKcuLk7ZtaMIkbvKWFVLEtaARpyU3H5BzIpfOkJtmYTGd5pJNHFAPj
kCK7V7aT9YXbITt51hoGXlAVt/BtVT0WZ5EsL8LAp5XrFnzyZfPlOFT1Ro++J6i/
ojFFtg02XU3tt0ylB8v6IGRyE0oTiH0XCa5scGs6JhH3t9lmdYgz1XFijh5EPitS
wCaGiYoJOVO8T4CsdVaY6vjfxhdkTVt4DhMPRKs1WTcO3F15b4bg3U0qh+GbEQHa
61FJyLG21DV8fN/ut/+3GqS2FmTQlwrGvmgNXCTsYI8akIvudQk4WUQcqXYBlRNl
oPEd4MK0u4i5A+OifTLmw3ggk90MwBk1nZhhHnZ5mAYUFy4l/shekNeAczH73wDp
zbgBOwjbWVLu1H2ihxci71IakvvfHEWHja0vz2PXizB8Al9LJ2YopnVK6y7np61R
BVHoX9r7JdLL4gptGtKkHhsjrKNz1kjeY3qKp9bzArpr4b1y3+IGaIiKV33hhU/Y
ft8B5i352ztubhTo6yalzQXmHEr/FtNm1gubyscXp9lk744Ec53GliyC8rBtu8Wz
NXu0j42l02EXlWFA9A5G/gFIK5w0nJUFx/ehVtleIB//oa3OfCA7Xc+qZMc261zV
cOcsR43Vjy9np5nXahegu8BH5egbRX4tHTxnMZcu0ntoWWDaMMP6l9pmPKWey4oK
BtS6f8DgLlSoDjNLWzXdH7oEqNl+Oar2E5u0VG8e9ts+Pi8N/ccvUJHfl9YMBjM4
kKSpSpaw0PC3BJ6YbfuDoHoa3NGdlQywHMkyBErp7jo9Coyo5+FLQLVFZlKlsDFn
aQePzqmrXu5boKV4Lxq9FTVPeK4WbS2SeaLOeaXBg8SJ5QqKHjY3fL8vIpY6tWiZ
/g7MnmBcAzwFV6q/yLWdok4GYsX0xwc2JlQAHeue70NR9WaRV7BSxx999p6QTld1
LgvtMZmV1d5HOQ300FIQVt1rJtuLnT6gPycIdZvWlCKl6hqhmWzXUJ50OXA+zrk9
R5emHHDXElAHCyUBJUILi9S+Jk9b9panDyVN/awiAhUGnXBBauhfewHMNUS25HvM
CdVnJ79tsvxcexXMW4B7aPP7Z4MaunpZyE4Pppa/UiTotKS5JTZ6Oku18MQkJf+f
nzCGUWs7ohRjJWGnj7nqZ00viQ9rUoS0M0jp4D/9WVQGXwf6lzElVjDMZnfteuwG
xe2KZjEASylawDItb5E8XIv6NuH7NUhavMbyy4XmaKJFO59jMdyERNey2AR3Mqe+
V3d9lSg/2DaYVA/rdvVTRl/t/YxNa0BA+b11HpwlgWfMkEL0DZEuQ+5092w2BHhA
6XJK5pXL1No2JhmcmkeAPQcgjLzcAlLNsC++Ou+PELmYJLUnpaHh5m9d0taxrISp
/NtOQ9Sg+BFGEUDwNFfYoM9vcHoDlDAVrQyG8MP01p+p+SHKEXeDStbci3cA3KTJ
qtxKRWrJ/sKU89HiHWQsIa1LDHV+zSTnzWl9IEMuEClUwT5/U6A2Wq68PPo7Bs3W
qDXk74HVAgHY5cwcLueXmrEH25h1iC/vCBEiiQv3JaUrkMWpTdJcqN/87berK9SW
kvnm1YFFQoDZXXF84ct392MZ30QVovMsUbiTTYyyfhynKUoGNOha73aI21nGBGzF
PjqXpaQobYcflGG4yKTo5kjjMvfnhNOxdI5/O9+yqAswdrNAbe9tvfBozwqNGIyx
/EPApKQVXDmNrY1q1AzHQKtpVpvM50y8TFAL6OyZnGj/xfK+dhHVHta9vxLpoLDf
s2A/ialONkQpOT93/PbYTiUfkDDNBoscsH02MZSQZPuESzpvYvyIa2cxumJWwGCz
GvWsoDbWPWwSNcAiUlm19+RLHKoGM18XiB+AUgdy6qMO4m20LcEgFslVH+xKjZVP
sRDYg0+6J3u1BmONhykbvDm6jKp/4GAlXHYANPx8JLggJQrKg8JWA3S1z/WQz5RH
yCkP274mhha50gEDROaZvT3SOxGL5UDO/lOPd5iKS+MWMURwynrmk6vQZGkPKyYs
0bFCjBYmCODyqmIAq4zpiymE9ETMvk9uJw29Ex7NKLo7YvcfiCvooHyaIKi6EG/F
FAaoja5zPT/XFISKkA5EE+JkyLnv1FJDGY5x2UR3bkh0rbhLLBdcWsy9VqztlYkh
bWYWAzPZOb32brq1THf+OJ86oJHVJe12XOgKojc8nLbMtWFsFmL7FPJ7aTrUdBIG
eb/I1NPmySubzT4o9ETWIGWxVyv9SuNge3G1vN2iZzDnz56twbFFlLGnwS78S5db
v/scCORRbDwNMHUSroo4rdMrkTHApgDrhq6BGcxFAwc8GFzHbsxkDMfyFABHDT9a
ypq2IClXQBzcjq1uNhDhbjYgQ62rfUyrGLkKuepeSZlAUNWfjkgqdc+Xo4g+zGdv
tIUECkVTGmuIomIrPAloClrOJC6vV0P2+34vNMdxbGbUzP1k+W8MnpUMgTwpL+ZE
7MEdrQG1wiVH6180XF8ES7I1T3tTmLAQ2X9w1ovtoP/NVh8l2u5GFiuYgs93jpRP
7iHj4iMZcoV+fbiza0WO2fHJcEQQT8tAuCbc7hqwGiCNXk7r4BdmFXfoeLiSoOXQ
7UPaAx2fQsZZYxdru/ByGJ0hYLAirOj7qx3WE49M0O2CgGhoz97EHVTm6xevnXs0
QSdndtbO0QUNHF36rQyQ6nR25pOv5zmYJLB3pOKse+453FoFMasLrwyKKv09q2L0
sZ/eNiYNW7un0pAp8w+eEaIGrF0p0rVMhKHotTjGsaRc9WJEplFaXxFzre+jCXhn
xW0uIzrUmjVrUue2OKRf+uXtLu3iBH9GxvxHRf2i2Bhat6tHx2JADYfKfkcaZMYJ
hApjvVp0REGL8ge3z+a/OEzlpfFdSfdctBZoviMRgqkULRloPeBWd4g4RNWxF/ll
iyNowRa01Nu678HohQmIFBt1gDH5g5odPPoxPs+lQaz6gw1ITSIzVKAYWTN4BDkX
IglgxzIItLr3xp/S3MW1tzKkEeAafnpCHFQbgqI42yR4KrGXsB4SJLhKI6QNXe5l
oKWngo/GBjhqYfbjsS0A5FrWCd1BNGT4LkM8uLVr/mItRV5MjtXddHJ7Y/1cqMAI
rbxce2axvcKlu8i7WhC9QShwXAsr3+/lqRdH+ItJBjX4UjkM8EYUmK6ZZ/D+orrv
dY5hu6Wyz3MF5zhYj2HGa1d1N4RdczCyaBEOb9MRq5JyTj/nXOpT3S+o7BxngI9C
4pXt0q1ZB+hsEKCzFIx80llJ8yOSFlOpbwOtXOE6/3PKin7jEcNQvzB7vV75IjHH
c90gRyVzOHEB+bQ00SWHAK7uM2h4yEq5bRrG4toNoS1dd7il1hzu+fQ7HbLP/anO
z1N5NGASzmJbSER3ep0PPty102dbdAPgg6eTlQw5LIRrlK212m6Qba/VAX4EhbGo
n0n9G+ffyBt4o10lP0t2y2ouLFgYPGs7wpUbZDQdBIOvwuqILa/CySnWe/h7Kh21
9opFc2DwZzoBtL/unK3XwmUECy4QPdZdJKee+XL8mXyZ7ekZlQHdHiToyL6fKKhv
2kAE4dKrZDSnWhvwM97jgXZt/rNaEBmI4wjHCqghz1yTfysV87HVu0pof7ngOiOF
D70BFnpx0/Ti1B3cDfIPDdigLH+CBi0RusIfrmc/IfwcuBq/KE1bqONswI+1Ylh1
lBdZ1uUozKI5jsvH45mzGJAc/z1BI0bBKprAtzLhxhykVCXLD/UP0dTXMgQwww2V
PmfSamE71BqrjeNNa+v1okM43kyXaJ/1T/cb+GA9saSTCu28vLCJz5sjQCh6yucc
z+ySo/ElTaqOaNJXl4NmCLM8iKuNNJeCKGEcrm0XurHixEhWI3BB2J6WRvJlqgun
f7pbNBU53DDr6QKXd646JW7IEiG9u/jfyHl+FovpnNo6prkz9MJfNNNVyG0hg9Ii
AVDexnYql4Z+GmfKvihHbp4c+S3Ws7a5ZrRfxX4QNfI9QSDPeJwSSZyhwIioJnV+
TaLKs2G2Kw2MrhvoBkddmLpH3Trmsg59729OaorO3MOOleK40NRIczFlnEWAwJOc
b5GJniOr68TJm3vaSlMPLuWB7wuANM6slBuxy7dUzQYarxjgdg8k5p1S3Opf4ZyO
9TkZ2ybKGyAl4VapNbS1yHcq+yiBnajUOj9NrPfazNhO1mHxDOj/pJvwUY9AdzKZ
ouxOw6YPq52r3jFCQ8psbtSKz4wNlaH60W/OuYaBoqY+rF/KvrVp1x1t9QB2kpbp
3LrCdF2BLv/b1F8gJ0DIz3O1QEEVaLlFdPSv31farDlyHJUFUK/CsQmtQCRj+Hb9
sP4W5/IKejZzwC7CElERAeli/nQRBTA7JSyXK7r0k+UWekD4xN+Jrp1pp+lSdPDW
VBvqD2OzyAkozQ9FiHhZbK/Fd4bX+kYFrjr32cKW3ZQR5sdfIeTmCe0/L1lTqVTH
RKojECm4Vbp6spkZ13r8OBcfDpVXXRiJyf1ZKUidFguY2Un7eaYA8GTAgyNzsqJb
ODZH/jry09ElFKpoTKmM/bUNNLzInywzOOGx5LjOzethcvB860UJV4hg9KEMEWnD
8qTUU4l5X4qV7VghXaW5vxGgXSpAmHaZFrvrhJMiWWJnVJJ7/1TRaasKYv2O1Zxn
kY7DvehKQWSORmk+2qF2tMY7jzQ8YIsrZEGt+MnXPYc28hH8BvcVs+2b49IdCm0I
YC3mdglNOWDN7f+4fTHu91BHPrdhEo8OnUntkXXKPtA8UOomZA0g4Sq9wrZNXEac
Gm4Lx0xWWf+xIWkyYs9jsZ4tjelxsi8oaota1grWVpacZKHceUO6iLgM30QUkH+/
du57t0oI372Q8NXY4AcL6endj8GUz7DlriNfNvcwI6jPqlE7TNtPNSM3JD14Jj72
UXSW6AvUhDPY1rPc8GgISet0k3OrT+9gLYCBrbtMHGvc/M70f1y2DoQB19/dIxuE
TDqmYLYslaRsSK08JzNaqEUIGmhXDWEQ/NscG+zwbs0R0KJ1vQBObf4Abb3EoU0I
6xnrMH6YJg7JmC09NjvW7lRU66F0XWU8jU3iIKI4RyXxakwXMZ0P0D+Pjn/JZKTV
f3zxqr14QCAGEuAbqGFjkLBicxkUPG+shGuEm1wSZ+iYwV0d8jdTf969AN1kDSZt
0ZiuzxoYBeIVBtkVThlZEjWec2Sa5qrygDO5ETlNDljYsgd2Ik5/kAq3XlAEnJrB
Hk/jn4vf1aG0deMfzpZkh8/ROcroglIynkJqm+1xa+bAtyNWcTUqenKgTRD4Smvu
BjtjhfSHXHU8XQYN/+yCmjbwpiGjamanZohq7/UFux0kEqtoVRF++LsyMPFTy+E3
2VGYEcKnAx97jWF82AK33oDGhbbDDxNyn1sgOTWvXB4kpiaHzygz6LGxkr/r14Lp
LLBvdfeN7MTHY3lyilQt/a76nAuETz7H9PqLoNjPjWdlaIUGu9vZ9ilXWJlqvJZV
pXMcn/IBykz/WN1bgZyVtjcqM+t5L7u5r1cJrzVH/vvF9adoA+cGFnpN4x7bVW1q
k66l5ZioqRJ4e6HS4tYZV/0V0sT3r/ukkusugvKIp7Ig9brVGmb/ot+0lkhPmwwN
Pg8/q8Mfs2RaVjtfOIOTDDkuA9lVKlgLodHanBHZ0yiSzTDTVjsrAek86EnvvB+S
pWKv7mrhWQmoXyfY6KpIqeeUnQMXBMMs8QiyXubbji3o2im5Q3AsFFg2IZop3Uot
alPtO44Cb01qQKc+QvvXyM99dRmcM3Yt9cuy2P8wVf/NdqbqxLZyByNpJfBbx0HE
2L2bnoxRQ/0zKWVYZBS1OUztoO2tPR6DnEhvFqHatOGVT8vFvB5G8IiGd2lH+QzE
FfZ18z926cMqh8jGFefL2zV1hvVPW3y52aYF6Lo/GH0yBU5nyEhlxSABbefc6hTj

//pragma protect end_data_block
//pragma protect digest_block
D+yHl79goV+bswYbLLsOdWliEAY=
//pragma protect end_digest_block
//pragma protect end_protected
