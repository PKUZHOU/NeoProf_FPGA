// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
JeBwA/RjCzHLxRs1YiIbASrqbH4iMMzh7FF3z2KTH9KDYmqaqrpdtzyu09eQbcDceJeSxlOnBmm0
NJZS72854GDSN61v1lRie/jZp4ziYQUKyW23nCWcwtMXryYPL4UiSM06/dKSNY/YsbVLuY1+tEfM
AQEaiINANyWqE4fnLtqpaBzxiVM2+lcfitTnPWLnLVwgb7oXiP7m3Xm+piXyDLTwXqLrkd80nJeF
rrX65ub3pc4D0RJxkCx99werCGML8+RzQjFpHWzBqmsno7lpehjjXoc2o1BKmWvWHOgWp0VxHih2
QATg9xlu1wcY04LxxrtmzkoSLpNX1S0llAEG/Q==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 30944)
K1eJI7kmQfUa93DgJW2yP5BinUBGKwy82Li/i3nD3wvIbLZ/nf7EkYrFeAskAHD+fI90XyJ2Ht4J
9Cye+rl5pqjYtKgOdaLMgfSSqtBs6mkGiNNhAfB05oRsHdS5oDXdUkU4tf1rwaoJSwvQF4rFfC7x
00lLXVhRh5vnjH0NYaAnzaWe7p0WkUedYrfpJHNXuctFwwqeHKrl5f7qRVCmAfwHyMcYZIgAVW5C
i7/EvkflHgNACTVeo3mEkraNS2Qe42V4BZ350H7FBz06j+vWfbdSCe1KuaAg0XMUmC2ySb1p5nnv
1JbrDTr307l5DFYxg81SixCx9cpKAjxmIvDKbrzWQmFjg75ZwM//mmHMpwo1R2+yObt9cTnIVAOq
RWRe1Hssxt0N647XIDeKZwIlGY4A6JERoSESuRF37KckOY1vrhf3GrH+5WrtH/CQfsdnN3uK7N52
VQufzklIK0y6cEqz0PkkaiMzLg9ptQYejz8VcpM7u2ixwag8GeWtLY0Uw45V+UJnDA3YpQW3OsQ+
peWnMGsHLljBzyY/FLYYSfYDY3gYDWEZbqe/AEgZJHBUecY6NErbJpHm8C2lMMQE+khPhTN+cDVc
vQeoCnJJ13Zpu6Lvba8FVsoH7+/hLvEtld46LNBlkgyt2744KGjeYnQ8K9jGsGE2AS/lA5fD0Vji
/DGo34fSrPkp9ixsL0YVMrItPqD09o22YztFHxJp1scOZSi0hLFmzj2pZ7IaLypEw0sUllWAZpCO
E3e1Tp83F7cwX/G4E11aTLipi+ma+PDVgJ7F99x3dlN7fO/ptiIOYXKgvhooppsRvmIuUszsX/MJ
fG/lZnmra1voyQzw7YJbFUhz0fruVf7LOiZPmET0PLRyAsSym26Rwco0frmzDucH09/Gpao7NwnU
Oz5FMrcxEZ3mF7ZejvsFMlc5O8LqiL2vFboUFcaKQkrXnxK1yzPd8ZQOqxuMzHJoczpaf/ZQNl14
OBDWhrYDeF41YOVh8E/GsiZa5oTcQlgG3/1UHtuJXc2bWrRxjO93leJ2xgIfKsqjG9yi2ATLYZ0Y
kilMUmGxdsXH5NsQobpEMhMCiLb8IdH26gYlwa8W88yzV4MwJKNmGQfV68CIKavZ84GCo+yXOIxE
Ny0FRbatLDXdxN1PMbx87MoTteefgTucvf21jcL7dYdVejLcq1OWOuvd3/slQn3/BD7xEZqrgjIj
KiDzfl3IiJHxWFOYTE9tGKbqOf1lE12DBNfSFJeBgOQcO3Bno/Lb1tAS0JbRifGjFoFWLzdG9XQw
InuFdYvLYgOGb2UKKTqkWU7rrnu3OLZaw7Px+d8yw4VD2iReVatvGAeneXrb3YI73MiRAo0Oceuw
7S3R/pjhS88ZfpG8LBjEDHoq0rRlzxzKWz/r6DTJtbF2M/CbuZJEjTgQyqriAiaGE/JcdMLLFfZ6
th+E7iIwANoJlkPPU7VEde8VvQtRWd+CzWrACJ4Yp80u/MxEZVUSgUI+PJ5MyOJENJIUJRGiqHiW
fbQmbVxVioPdYl3wi48Gv9Dl9q7aWNyZCANxlPSHujBn5Cwzg0iK3/Sl8REoA12UhNPyulx1nfNY
HZAU1eGN6EYtuoOvpty0EkO0hdnI1XTszA+zh9MJad7FF8RVyH4XBWeBPvitMPKT1QtfBgHZFKgp
oPufx5KZK61xQxrwLDMZwWPu8hSbKdJbn9ixLmxub5CPKa7Fml4a2seRLdLnv6ECWp4goKZAJ9aI
Tf61XQ+JJHwuT+ASkGBp/Lnm9EFGDudabLil+Zu56NQ09IJjYoMLqKaarpcKnCBYTyemW10v1vRD
eHQM0kgX3W2robPhoPk0Bs/N2t9LUDnxKRmIBe5S8xkx2Fmjh/lXNlOC6DCMEznMGKMYWwKB/Xcb
XOevflJ60ZY2iWeiTtEpWE0bIUACP1zOIXLyIIGh2EpRFewXsoE03R9Ffk9LPh/ij8yPnJhCjfTf
jIheWxKqhMvb53/A1BXX2nE1wGqLdZmQ6kB8EA7t1Cjhsx5ORQC4wCrXYC3djvSOLGBuoy0vIv3w
J/+gpffNf9tKKVjAcfQ23xM0zKbI/Mi1mTrv+4s/cxA47uG8dL5ByUL6OQ1lSZr2qMOGlXJVVfuh
ex7EPenqduFtNiB/2EJKqhYD6FucoEBA/n6YHytpyDaZJJWeSd4Mu/rtJaN/4KT6nfLSyzeWFc9J
a9dV6uHqRYSSpfGR/48+LknqU/2yY6LKgoaH/vbBkbWBctxsR09xJoB92t3INBXyzppAlR4mi3in
J2rTAlCAPtKu9U7OL3c437aTXSYKI2x+egWXdrCgDo+yP8SjNBwrjEpw4TZuCndVTg0deHPO2sPe
28JpmHr9XzTxRPZzUeQIKhfcqrs1RDU9lBCLYs1k3z9Ut67Zpa0dYT4tPRxmVlc28EEQ3rmYjmOo
LpQWe1oicjzlWpThIk5jeeEOZN6IODvYKJdIOhq8jS6RzRCHNKXrB8LnpSr0yKWwtX1/x2ywVYTx
K978ap6DYmzEj81fVtY08NrTqxla49YVYazmHFZYIgf1iCjj24CLWn4udxd8p72PIDSOR+11kiRH
of4NdsOmX5jg459A2eMUgPHUeq6mQBnnllcxMYXNHq0g+23vmxbFlLGQJlRk9WvxwaBLycXagLdB
hmLb9rOP2tfC3tXIS8mbc45Ni93afEYuh+tl4FrIGLuzo0qlfhWcsJqHZv9Q+PaYM/UlUqyDGMkA
09NVwo8xe/ABBP6BLrsypHHbEeDCSt7JyFv3mLl6AvB/tvQDYSNfP/UEPNxyxUpZeNYoTMi2qTMM
kgVCYJGoLIOKfrpvQZ8R8AyVOw6IF0L+ASq97DzHDacze/IngQlEaU8mvTN3R3eBoEcdnBmKnwUt
bJmh7nWa6WSvvQ2Wv1E3+DUhsXcx8WRwmDCv2zGqj99hHYKzShAQkl8STcRbX/RUe60UIVyCyNZp
wksTmHKqzXd0+OVqsMEB1P3+GFflWVDzrE4PiT8VqVTsYBTm07w0XdXIRI49ZMvnXCRTs4SGuYFN
MzAxzCIm1ZJJaBruLiZr6f8PuT/C6oV19k/787QcCNIBAocqK4Z78/3vRaqKnqcEGhfEvzvyGpJA
zZTQQ+2ogKV1q9kvte3CH6MqEemu9hkNODYZZAgCr+CpZCU0bZZ11rjX4TDRes/owM11ErikS+XI
xft3mOYVkpoZlIfn3y28l8AVk/+5ZSJgJFG9zYjtCXpCAilpjKT0qfmn1wbSykT0i8yLmYJXzJIM
SVBeh+N447HoeqDCuE4/fnfVCNrtNbwnYlmvsrjMpAlcU2/oivd1xtGY0xlSxRpJcp5UgaQOc7xT
y2ix0X7dFENDR6VoKRz6q1Z+XlekZ4ElLJ1lrT3h8XuJsVBCspUTvAeQ0UXW/0KBlKnDxTUxpWvo
n7p+QrcVJw+xTdyv38Gnq1e4cwCnSQgEpkqWIACjr/QdOe9K33d41ngvJ3YWvCShYEEhggnfrRz3
ulPdxlnU7KUTOr0UxX+wcRoYlqt9CD8GQbBxEKUuFr9AXrYEXAV6Hu177UR4QLuLK1VW2m6M1jVN
y8VP15il6j5jBZGxeZc44Ont/118KzpodGUiSRCCYtrtmNrSY+f34FFE0J/GxCb7sPGeNbx3ZL9o
l8L/9vTSn0WVCcuLcZaWkDIcU2wAv+jVSYDqTqsfD2gdCBBYS5yKk6+geH4pRIluqGhKvZ9xXQQ+
7hcuP/P2E6ybHonfIs/yeeK/eBqaPw6kO8jXZGqjd/k5KBx841LO1GxPzatpM1YZ5TwVpA6iWtGZ
AnQggHy2vV8nnmJo1ED5FhnTp0NfpSZ0uAmvw6V6zNGb+XmgE9gR/ic4YONk8dYmOmIqqnYau8ka
E+ROgtL5Veuhc+9UEFCPfuNPXOjj4sCQanul8RSLFLgxFKsA613KiM8QVlJJ8i2lh37O+LoxS/6v
lUNuV1mwBAPKXEjMoUG262mNt05b/7cuyqnoU4gix8/SePckMi/YCRytYKGOoPGXI2Y+fS6C+7NV
CIYfHWPFFwmonVzw1c1W7p3HAfhCnoCaiyrxO2It1mi+9IDTYo53uKzF7QbhE0J9b+Tj94QszcJE
x44ZNYlLwRi5MJNGdUi6HDoZPzB5h8pKbKs0OQM1wgojy6AXM7Ucl451KX8+RwisjERIHelI6UCA
efoEhJqMtNBbZ94ewiL1liF9sR6FZ5+FAIzhN4EwG5ipmZsGfxMyctfDwHuGNhsNHmDw1FBbui78
gAMDIje5f1I72ym4EjOqHr9kmiTOh3eWCHC4kbce7WbO7mLipuTiuId47kzS7gXdYXgWBX1mOZnT
QlymCYa9OGaAmAoDq+L08ivfRrOHYtoEwQb6C+wJDigYzRaIlCjLShMneIGErdg40v4UDNaZuUXd
/rA5G4czf/J6uLwcbynLZikB73An0JvMbnGTUHoi8wBTjBJoF/tX6WiQ34zeAs4jePvUkosYixv5
EuA+d7rI8QuKdFW2W6Z9pcl+GletomU4Yd9yNgKdLiQ+0oHqTiDkDhib8AyAyJE/Ak/g0KcULsis
r3kd5h1mQxCyivrDjJbns3NYmTq/LrabQ/8gOX/Pghl+Fw/7eQk/8BkGmQlrkDDt83s8DTt4zn5d
bH6PmIWw+qraoj4y05yD4utkLMX59a5d4I/A39ciWVaru1i3Ed9ke3QhQQsfdrLoHZwqSx8cnA0P
YWRsR7PuzNSPQrl/T5BezXPlY3xvgwarTbGL/3i+BoCMdCNMoJXMEHoQgq5vRccSRWotxmjG1y9n
ygzFRX+cWyr5jLdLx3TTtN8WjbNTJIuJB/DtJSAzKwB4wV6+D1a4tf/GMGyec4EiyT0OI9f84/HY
2LbxTDkWW+3d2+Ho9qX55XnM5l5cjsBlSbHDtJimG7OQT2qaKpnL0kyOpKYfbD5wd6i7l6NkMUnV
KWIPcn10P8o0g780vEWyoR5x7yFD91wbHJKXitZg9qy5dlDm4qXdg6QelZ6qH/3qOFDhbUZU0JTQ
Y7jVp73qzP3GPRSsNERqjPRTwoBwsxvOeQQ2nH17wVo2+Wok4szh+xIodb4USe3IOIfUZFU346zX
5pOVEJ9lSZ/uQNNbo/T0uz4XGeImtDEqdQqtVOmg/fL8/vm9HjlgUdnIlYxJSialvs0EaW63n3kr
wReTcyLaDdC5Armo1EX5mF5hxwQ6fWggn3f8x7U+XOMLQXrVzqX4ZZab0W3MIWyhbY0ukt+j0r3o
k6+SLOMrjdlf30i0kflmNpspksyjqwnXPddaOD8wF2jzCiVvmhYRyVqF+0MxEeFZWvQKHgbvWRZD
ryXbtHoot4LbVvX3QO87xbB1h0LGJnIsNMY117eAQrC0NJ3dEkT7PQza/Q7SeydnSKvbWdMW1eg5
utZb68lqNsE1aP/TK0WQOYnQ+8Y4S+b5gaU+VCr1oQ2R9Y8O2engizEqvFwXrNJphIs9jQUbKv3u
ByxlEN0D+iT6LhAABAupocFf+gMjDLxmzsDQ/vIpsLOLcAG+HzvG6zgKasx48oHPhYmqlOX8MjhR
eiDfng+bueZ6DquJuSvqNUfDvAAmZNMNee7Q1oNkYFL74db9HoBbG7nr/Qut5HDDwNdN8l64kEt4
pDxXmoYOj1bDf4/Y8ZNCP3xVFbSXlKvR6XaGJU/hSQvviniPK4s72MUBeUgxamzgWCpiKcZpD984
deaqM71PaIKQRjdvNcj+ej/kSN1t7ajXz2cvEAfJOCeJ2K6A4qB7vZpRaCDG9v5eq1qMnyGnzZ99
jqEaiobl/WUA/aw3+gHj/+R9ohAgy3SaKMcVrrWzLJcORCbtqTjvuzGnH6pAyfyXwOcprEofTOj5
Juj0g3VDyuBPNpOXnl0NGLS6NCZlD6QKGgHJGJaET0ZQpRrRKz6Yof3C7kgEPuZNScF+tsCb3iXq
AX9V1NW9E+V7EADS+il1C0CiGsQWXL2YbJekjxEAFIuo3tpyq8L3VaN6bRPfXwmRMkYN1Olqvsz5
NmqjDoTefn3fdgrI4HazD5MYH8PmD32gSa+ZsMJ3mznhyaGQnRwsE+ezdfYGsHsNqCJ5SiazcxbH
AekHd7YY3vXFYs2/JuifQ9oPRObBhHtrHBy3a42llMK6vrluPV29FHw04/IJz98jiaXISkaNGhsh
0Fy7sjfXeoqzl7UYx3IsJRnu9eIJlv1AltcEheJrpHdlHXjA8ewMvTIHZAtiiu8bUdvMfzvpTTza
ZET5HzkQw4tsumFN5f6zwQ5hoW0xCXM9k8JUr79X33CUnF66vONYx2pFzV3whW4h0+qsfzf15y2O
f1oHzJXrR3Id5D0KKKdLQm91ssdWCG/sPK/1GBOk4aFC8SCDq6tWRRBqrDZHjl+FDdu1Gy/790D/
jy9BxzU+Fjwd3o9XACDGrO9hhLAO/fHxJcb6PeVNepWgWHPQy5qpOYqGAS2/EICFKozwcSqLbhJE
jBaHnUB8alJrEqOWQi6tPM/1xoxbmJd9c9uvglGOA+VlWSW40rF9dZ/ne8VUtN7+DF3dhn/61Acy
fe9PlxwcnuAaTLjFH0rz45QACAHUlcIJ6bjHjrqJXgm1RajpTY9CEXfJy8g5sA85FzUQLGHz7o/w
WMcy2GzozErnz+IP7kAKUhVgiwjfewn2AiAOMbm5BIV6TLmITuhKrx0OqNBv17r5vYwnjpPnaAIB
HLO2SVyOI6eUzuLTBbObJkht/gDSvHgueGwSW9lL/UGVZ0OvEt6srG+OlkcRNhTIMlnsw5AbZ+NK
w8vxJHt68E2oUCVqHFDrEKpt0ygHcr6Wkhwj6/tGykqg6XC4HZ0RnPS6L5NFHEGb6dsis4qxHsCw
r/KZKR49OXw4npEYcPmHKcAq0GFAiLqx+Q3z4EY/avn6RqZQiu9XFQgw/+Z0dbknT0TWqlZtVNvr
zeO0FzxIG/OUSf2wV7Dvl/EqYJMTga4Ml7YmzG80ocRZijOyIQ8l5A9Zkm9gk3pIsbu9xqrVI3cP
ugDKuSvYP0RCfQMc5mAQmMrrqCgI706ypkzhksbbY2tsKStC0yJO8RD7PG3a0HKoYdYXfZHQPsaM
YdJD0IjYB4iuqkQIBJW52azxh1hzDXmt1COThWDCpiRM4/8koJns5ymvvwvFNZ6nV4XPyi0K4p4H
6vkaylQ0V7bqmEEFlBtdAm0aYQuwTCIs+JoetesF552cN+mksZ/SYTxCDeKQ2/1ZWE/28Ei85o4x
hR3bYDJGbzjkUdfAu15FKMCvnwlBDOsZGRRR6ZytxGFtaULY9iAP//BKUAWk1kmdGUBrnqdFPJkc
Q1NObTEO/KGmYJVSlS/EyoVQU/VJU9qZqtrQZlv0AQqUs6lizeqeLnQU95hf5KCKJQ6i0xJBKbo9
G8lEepfVjGQZqXwA2jS/+SS32j+mFPwtmZz7qZ/2aIBjcNuIpQaPVUFnqqwo7gzfuZaPp5JHWGlK
hFO/30M2jCcSp8IRBme9gjDlxhMN1Q3hceEyLo5B2VqDZJqERHQ3VU2oRp+DQzDrK+OByzc3lb/b
MnJkf8LUeslm8D7IKbmPrWJ45T1yn4wjbtHRcNME6eGw4cbw1Cejbwzd/7h1Q6lJs8QMb6lSlChB
lLVVqfQpjbAvl/6wOnMq1o5I4+dy+lFEY19Fuc37bHG/NT1BJuZL1rI9VhOQOQamOfxFU/GQQRVm
To2kQxrHaW56LSGHufNSoRY7Fy1UgNdPFZGV6eVrKdrzBf1zgSx507BfQ89paREn8tuNV/81n0Hs
WGYHZf6DpM67rEBXIbm7fQngKfSo6WknwdMOBBY3+UDh2ZQjkrPqaodYbjPU61v+FmDnA8rdjrpf
BYjOClylyfVx+2FLvtkebuKrzoX+884sLyW8l/vmQxpw+NqffWUSHdUvMXKDOTL5mfbswfTSZoDt
6N4femZ+ZdI1VDvemzJXzYKuxB/hFGoO8veCS6rIcttNHodiAXP2U0zHbE7Mmbw7EKvrAHBn2Qov
Of41dzQ8lgNnZ+9J0zjyiDOVlGv2YLFQRczP7H5AAIae2ice7zIDp/4i2EmApN4cQmLmXnManlPk
DPks9ZgeNDxZ/jjON0A5x3PtWGFSwq9lLS0rPlWWV4YZLqFjn4hPCH3UILP0uHwUK1LEjvEgS7yx
bxJwx1ZpZfl1B5o8fDYmX6Y0e2wBcSTVY5kt1yVtasV4qITOnaSogh4/fITRRmxoRwnzmsjeFR6R
eQkocUrMBdDX5AtUyUU7zT2s8yO5upYiVNKxTELvlNFkvmvol+nE6Wtx37kGUUIZJrSxfNga6ztF
2Sj4DJLd73H4TtiRK2ba8v2eHQJZtZFwB9gcxfr3qCkBL2kZuC0OMP0DOeVjJI8ZHrWM3VUTKQqs
dgja9uR70FADIRdoLxu5LruZzWQ+s4yioTyBEB6LuTruFFkDyzIY5Bt4gRdAkqHXGcICYig+U6oy
QKSH3xtIDUd2Ro1GdqeveiZCVGdAFfok0UPr0FM2hkC5Pgp0f9iMQTBF51z2diXI4bUmcn0Tn2gT
pEPqG4GdR+HuBJy06iKbUgW17iU35qbD7gT1HVPK0NM4yt1vPXINObxZOUMzJj7uBw1kf6Gp7rbA
rSrRffmDLS4ETtuzRmsK/WlZM6uX+ibbWzzXy+Ivv5zseBFJs33SgD4wh6qlxGLEvqnU+2dBXQwE
DtzGHAuDy0TfMgw0SmSyNX1/4uERmip9BAUi/oIEj7i8UknJzKpYH5gfD2wHtVR/qIhhC8Fl68Nz
fGNFDyqmLgVgP12le6MSV8Aq01Ok4oQzL92UUsHIPx6irNG1MQPjs0V0TMGJZjZ9448wOUrTf1RT
sVuuqQ8D9Mw3roUMc5b6waOrkaHW+RYfOsSaa31okH66VVJ8ioIIFTncL1irf2vAGbNH+4RzGwdB
rFO6BLUCjYnZ1JvbNtk/iXzem5jy9x1IC0NqIbiSVgGfVAotQDvkQECklM5VxSuf8GyJsrg+woTS
mB8R1kFrL3B0trke0miz0BuIy/fFiQTVcWPnRWPkR5sv6nF2vs/jVamotOAtBegmCNec14+y1OgH
LGybzTH8SHsp/dnq4/nisle01VOGHtN/4qDHO7s478yJnCEtyj8im2iS1IFoidfEUxWq9Xr7rawD
84+G6MtbdpJLl1abbt9ZvLUQP6VVoM2H9gk2VYlbUXtWjeR2QQuqS+aiF8zrM84hiq6sMpxbFM9N
mfWlJYJx8oOgd5FNswYZ0uZHsgRHoFRec2CJ+M/T0EDc5Olx9QykBQ3vhBEkF7SCbT7sifOpJqzg
xMzAWIDdDja7Zx4eUILYmiA+wWBd1O22PL5aHdqKhYSsm7JVxz+whIYSxoeFMzsiGoM+mACw1UD4
B9KAS9GLV7Ug5UEzjaHCz5z7Htk5WMN81jsCqO9ptYxF10K8MMdt/4UxhTzVYXigkuzpquD3z5Zi
+xGUuOQJjAvic1dZX7U3Zc9edqQ/ABokHS+T7/FEF7mEqo7ZcHbJ9eyeM/RDGqG+EEIYFWcRBEmB
mOohgurdD41fNcvvspI5kVg0dUO/NOPOiXKSWupWjg8h0s0+O2xKcJHxW2iigH7hTgqAinLExFqt
4Df71OqzzA/q5sfTUkpYzSH5f9IrfHrJmZF8qNPCCxggwQS8RnSq1gpMORkMqQ+pbC/tfpD82BmB
15htun4NFicgTe9qjws4D0D8r2zySwON1R25lO9m/sp+WH6CQL5WTy1h47QntAgJBFwD47u++Q0C
hsFAbeT+Zq4VmC4iM5vIeXPlQKQn2WLXPuMLWpO6viox+kEqKAoIGLaXsLSNskpkne2wMM0q9dLr
Rn0L5fODhK7FfL78KL6Hv5ljs5+0VKNrGBUUoeOZHlLl17VcTvZPHx9UsfVXS2EXkgia1mG7pENi
t18DvOENTrZCsQsey2VruUuwsY1rEzSE3aOhBVtiZ9zHdihSKYjAvHrwNBMkneHvhC6Yra1b7XsM
vIdStYYBj64UJyreq4u7/XF6o4wxrp0igfoWy2ipqq4pxWWqk4t4BHDUpQl6NFQjON/t/2DFWZz6
wg8Rz8J1TaSYoyJ6Qk5yxYY513XBb3PrJnsLImy6NhPvOes0MlHAl5N0VSacHM0kiBwRa57h0b9k
gpy6ReYmpO1/TAw9SLkt3cXtpAwlSgfWdOLKabwQaOE/XCFz41vbcncAgM2tbcv8R+PttqBZL41D
/41mqWk0FYsKuYAgdtoCnBR19iGHsKhdyAqAtAfImzYSDZAJ+ZXwxLcy50sqVy4/OcGoj1FX4gm9
u+PQDk/ZNxehZyIvcdLdSfJGn2tFUvyn3wyUkM9DOttkLyaiOcKGE4QPBayLqFrKe6gxp59bRCOf
4/1SuvPVfvohxPcI7ZX401WcnzTYdua9BfzKlc4l7NpuJ/UkBfJkbUahJtRpTYe/cJdCtZcrNmo4
/8ywke84eQk/FaT2IeMWw7s6fzT20ZzI5iiT2bkXFVKmrPu3dRAEpnQy0MH/DASGb54NC/i+FIS/
Mcb0EQ3JD6dmIFr7OgTygf15+SqQRc4fvlqbIsbUYj0rVaIv5+3hLDFhtAp5Lt/mqyAWqFD1EAXj
cDhjFnpcnxixwI4fuQl/aTjhoCNwpLtg8EKrd5XSzbAQaxZUFNoeDQUfUFC47IJng84UcNk80e1z
Shzu7mcBskPu4B3MbF+4nPjjJX3m3qPTe3RF+dlo5RegVWu9hTYQlIygHB/fKE07mbT4dvBiufQ+
/6i+yYoUqrg4FZyEuVIXpNUelDdCDalislOQUERGZ33Jd/FEFw1oPDnMZBa4S6d84y0WX1C1YCyy
ngkMB6MrB+NHsfZxiq2+nKn4rLUwnYlgJVulEn3nJur4AQROnh0YLoGNoR8x1kniyd093MrnQSDJ
aZqBBJcv9FdCsnYYJp91UPktAJGhcJ2uR+qjUDj709ONnR0ETAXwOw0U2HBF4p6gbq9437JqfHjN
OGco0Xu8Hz+/7Y8DF41Bu+7HwAWUaUj3It9bvrjxT2558y8y70sq4oaSpS73GAlWODNBPbYKAc7O
wuBCyNweGTh4U60Ct/dRslI7QyT49thSspgtn2ovjGBcy67sHkGXZzCmH6WwQqtwDknw8inJCdXR
HT/ZfkWXLSzAuIet/ttCuywb1+RdKmxSxksmb437uqO4dnU/RrJgGlS8dh/Sr98tW4A00TbMVW15
+kSXVcxftpSydGBnqJf1cFXcFRWA9V94FoErkFmZ1ZN9ip5DMesZg57u0vnjCOyjM+0K0gO1nBVx
k15tb49AIT5B/NVt1V4OzuuBYSNHF7c+zu/jdYWyF0esH46knnTYvVzDhnduEpmYnT2lt6oDHVEd
KgpVIhrLR5XiW2uKd+Pg3UBbbeVH3JVQfu/hSaSHRpCWmji/ZVJ+/PywH0pjXEgQ4rKa5SBiw2hA
jVZK/E4FCH2SppVN0vz5lsIHbMJQyM36H4mDf6h1qnqdo6hBxKhdOSndPczZqGPKpDJpnYE6A9Ck
u9+2Pb2uYLUza1K3ckyAfn9favk3G92mUEnkA3ub0yawO7UQpozZEE0zQvEVokRh5k9rd0VERy/W
e+CDImgI3rq3GHxHSk7x4suDFmEQWhFBrAiE1NHNAzxbWUgl7hkFp5DntJiAP+EybaWUAA2yZeoB
TguQxuAECmmpZi9fj+lrlIlE5EsaBwhOjR6V+5vYz0U9XZ7ytW/NvUdprjRmIY8DlqLf0qNJp52r
MlyB7GEgobvsUbfD4YCbC23JUXTaVb783IVdxljuKeK7CZT5AGu66nwxWzwaG/SLL3Tvj0/GHDoh
Ja45JcpEKsqoFmzaG21HD6EvypdLa7JaD2EZuknENTTORdpeOZ+Z7umv+GhEFxsKqTlaLsnYwh1o
D+TcDSj1VJkW8L9LDTNpXIwhFUk9FST3wJobE/SEm/QSCdcuYqGpfhOzRnv7C9atBcFvF51QhUcf
SFaaPk8B2l0rZWPs0JQmbt1gGsCaK2FxJLirpsCYwzWbjhXfzTuLvjJEgxV2u9+KLC3EQ7pavKgI
HyxqC+CA51TFuCvykL4oe8Kv6gtqUzVQLuNiKwEi5H0+dBJ5dLm/ySnTDVvuXziHvkSBzBw2GDH5
sU1+WK2JNsZWR9jSq+xxJMbEZgyaAkfZG1pbHLAW8FcHheO644hogcSmiLRqCPnGQuM0+sW6KGZz
os5BFrIMdOzpwT3Ryb5QsztiziSbrna+fddc7KIJg7e7XERxb256x4QIEHgURrf9YDNUyiwHYpGp
4qEXwK0as/ChxYnmkNvh8opqpHNvCvBv99X8wAh05j+BbDMMKXAcJuUNEW+MK30CDZw4DpWhBTub
5UbEzD0Pf0prNrZ6l7Pkrl2IMeUBgfn3G8bfKmUPuM5lvUVrMWKrZxGpRGyEJyVN+WUQaDiTmBfW
VQNt0VmRe0TckpWekRjqJG3p0MZpr7y6oue03uys8U5oxvK46QvhERV6fS2sPZRnJl+cDKK1Rqaa
mzXC/sQ/FK6mHxMpJWg+YPfLSt1lMMZ33pJ9n9HqN/s8gVU6b5a9mhDwrUhlIX9KOxCsfHefK+Dk
3yKhG7Z56+HPfhrdImGXIYkbOmigzQQIlZ7vQoMSVR7Ukp0zVx9f9RLwCz+WYTLm5mFDcrlwTLzf
SYYm1Wirw1Fr9dJboerD/zcvys1g36XGRoL0iO262lqO8GS3SFxoKo1pTiM2TCoDxq7jDaRE0tDl
uz8tWdBEAKJiH651GVvSkuI6NzKHBv46EKZKWqpdIXBiVv7o9reJY9dOBJ/hPwc5+wJyas32wEDE
DITQzyKTT9AKZ4vaGH9IrfogUmzRmYN2FK45fhryKdxnlvUJdzhqyUXm7m42+Y8oSKzsZbrEp9JX
r/g6fM+1qhrutUFUbJgdFXQ9D5vZeOEBQpPpN4qJivqcNNhx/EFf2hoWWP3lINDii8QrYKAvOQ9v
OIAeq2KWgrr5CtsWJUQOD4yTWJjIB8vfwYwkEci3gbugOjM8aLoaO+0mljjx0Ssbzmphg75y5RiH
h9xjCWpd/ksef4/aLwg7ymN/OFYJ02lII2ukx8dP8YVnIaUrkgdSynGaOJ7qu3BSHK5TW+r5QcDn
w/+kjsOgz4ijCrkk+2fj88V8qaWgz2Ej+3NTHTdNoCzAM2Que0AwvOMJz0vhqxHz2Dipfzgb7nrV
7dlPFzY2uxGFZC5G40TSCUnZ9CbHQVb0KbgvcAj8Rj3h5+G2pX+vbc26we2KqXsxbPMGwTxqpTw1
wDAzuUbsLQrrJrK+QynAJWLy1NoihqRQ9h+bNi196ZOmn2fEcYJ2wJOJAEp67zXC/fcj9aWXIYIy
xJX04WCmm69ZpnXubZyguNclVPvYRYsmiTMxxgDJjYV9PLZgyYZ6Wvr+ZIyrFuEB9p4wjp1HnpZZ
+kigbW0YUYAhZVwlEtnLFUiFt6Ci//wtK5reOWQB9XZ2uOXSSoM7qCzT06gIKdYiqKMAZvwzJR+5
LJ8ZcWcAkQcOCThtJRucHiHGpLkgVbFrPQEPUNR8nVX1cduS1pkSNh2k9eJjQjEFISW/ou4/2B5n
9h+kt9VnPQmNVV35m7kF9x4L7+76wGkj/mBqYRPh9lO0yL+//2fiSrWehbov+ro+r9gmu6QcdQRw
3WFZKcOn9FF45hjQUSMyWZRcfBxK7rPjqIigsdFATeX7hg2MCuD5/V6H/mZ4UFhwb0BHki2asZRT
mFn7JMUC5DAkzHDLdoQ0RX3SMIW2BLAfk795zaIH82+TzLxphEZv/NcAHCJ2RZNHRawB8/My475c
EoJBWXo8DHNt+LcvqTPxRxaUtP9gAi2ot0zoim6/5acIdgqTLFYjwyixdztRlYeOlg+ixNzBZFLd
0qQxVKJC6tTmm3eQ7qFb46StXs13RRxDK0lUyjFL/a8EI65hVGIGQAEpUSXRrq+UJxGAuOOwO1lp
WJcuBBl2NLsvrYVqjA4k0CSt4/2G8mrUB7qUu+D+DTgnvYLQdduenuCdot/0/OhrqBuRnmSRnfor
y1VzhXfKHaWFQfZj5JdrFXp6N6AVCDLCj4tfSl/tAsYlcpe8pHEJpG+YOsVNbhub/jB7RU/tlLiS
BunDOTYM2lhkT06ARAq46vNDeXM8ybEDiT30vPs4fJAvQavty19HKNLz5eZ9lNpPsnOfDeVKKCgG
dRiaNe+Ij/8E9RTMPXV/39eZzwJQTRP/4EuZiqrH5FJT/WOiXMuakIceyX7HwqF//mm8eKWrOuks
3ajkipLES4GlU9gNOtCSB43pfmyYdypWEHf5I4c6J/iDa1sTaqo/kI0XaSQjy8iyYfFt/mB33YSa
3UGXWf3z3bAtG2ZMpsVpSuLQmqaRPixsqb2mcOdUj6YodemPYDsl/mT10BC1joUOtZiSryfprMqq
pmTO9bWBZJ1EycfAhglz1yTaESwC3RJ8PZH+SzTraZxgSkil1/D9CCH/ekLFOdAl9LuAoBPOZrmH
fjp44IwCDvlSgqB/L9XeZfuhcxM1IKkKF8glALckI68gtjcDv7FLxvkmHJvDc5KShDiz7UWN5BcO
6lsU0pCU0Gu/mNzlyisKNLLPCy0BEykWa98mDDN30CXjU0ZLP3rngX4X+4EorWgdlXUpV67siGzw
vuW98Kh+P28Xqiy/TKwFGKp4rS9hfiejByjl8MOhawIwtBTMp58HyKXEkHqQc/keDfWSpsi4T8yN
peLMYPME5OaFHcFrnYtQSQb9ZhiGCVTSCacEF+rctGiz1I4QRYtK+jizUV/rXngCok0+XK+KmljF
37uKKOfl9/JbRkbxJ51DYF0qaeDs+j6ZKY5HTPY3R3d/dL7sqTvT2TOqDOr9COQztlWlsVxtNF/4
rZ6MeiC3QzC6qsplMJHNHjHu/lcfsBHSuCkL8urxJ/2j9a3vMiWKCTjZEvj6N20wTvNkLSZCTlWT
ECjO6ItfVb4ss7ZO96OHtB1Gcertt+P97j7jBedKG/onftm155ZJH65MJ/dYi0mT77xOVM0cy+Iq
DYk5IJwYglDLLXlbJiJoFD/cyOG0hTU1+JrpQ9L5h5QRkraRPtX3198qjB41slcmOK7x0EIT+2Im
Q3bXJTQtq9UZo1X22mLf9w2v/MmC/QhZc3SQQR468DwEs/UDeJDy29mHdb/8+RwgBStWI0QMtuDB
9xL91HurfbycCn9Q/ON4IYc8jU95CJOXwu5TNEaexKokMNA5/tEasn7CTlwu4d77hq1Vq4d+F+qX
G9D2WI59LRxhCEsEmeMezl7D++slVT4McqrqZFgFD+67evGA1f4cAwGaoLZWU2U24E7vjOfwHNPM
ypjnSErS43TVG45SJdb2NR0mDfCVaFtkfkZ7Qxx4L/WjCX2CynDiTWilwrh20p/D40wm6As+bm+P
kqEcHHwUW8J+AktOe4YuKWE3wxG04P8mcyeuk6/gP53NyJAIhyUpGUCJyn4wm+uZZ/EVE6aEB16x
9u61aOkoxiyHRsAIz34jFM+OLetC/kXPgl+W95f2UWCoiaitptW1Dl4KrGyFa46JdWnzKYfkkPWj
2UQV0rOtsDv7s8Iv6pJYCQh14xoqOP4fL7XY5PWVO1fHde5ZkrFTBtGJHYveiWc/7yk6hV01JuVw
TBgzwWmm3GXVwFVlxkfRpvFLSJCEZjzoa5ygEWjPvYKjCzc4IkI5T183+EMGtHuXwFRfQebJtzGZ
KYpDpZ8BCmeyrzhOIXefqborg/e4GpijpwrB/VanpcQTaxK/4y9pQ+6TZhM4g+LgAl+GIzt06mO6
j0jWnzv8+RJg2bndVg9qmn8gFdPixgkWJiVK543N7QyEeg4e2Bqn1Qgo7wSoxGgglc7nmfhrZ6Rd
q6DdVMNmeaWEEBeX6ZVcL2a2/DMKRluIDHtiSwHHG2ozVQ+hfRWWowVjdpl3010bXEs8q2LXiqRc
NWWEBhCg4bAKmaajnFY3MbsTHIs2bsZBBimji0tRVn9mrIGG9ThN6vvrcBTz3YqB5JvREoz5xfEn
ahPwKnkZJgFOYaJrlK2gHMvyEJHeJ3nJ49MiB+R0++p1TfW10XsstoByC85T3JTIqUMLiOvKINic
13JNPfIJlJE+UWLaa6ddo6Uj89jSHF2qjTlCpKKrUZayE2i9xUjxKJ8Ea9nNAkGIZNjg+y7N8Stk
3rH+Wy+tH0ct0bkxCuS1NHgICT8tq6poECkcm/x8+zjSVfrTikzOavZnkXAh2Qn5qvxDWN+EcZiE
JjQoI/tWqEyCbmSFCr/7/q8uRBCG8w8v44VVQYz+g9C3riEzG9nPJLxfTE1Z0AgfKR7LFdZ96PI1
4u8P/SaT/YN6ysmjWqtpe/yGRNjh5fQlNbqtXzGGEIlapVZ0UJy6Z8o0RNZ2ftMEAQQS11bFvob6
dS80PjCDc7TqYFk4qeEjSTgTubfxe6I4LPl8jwecOwQBMIbt3zE17338/PCjEFHYylCragNuPSdK
l9PqSmd2A0IBwaXJuLOH5TnzovbCADqoZ4ccDrnHcbv0vEk8+AKSVcxwQECeIjCOsv+cj0WeWql2
Bmz5ZmE+urtiIf/f1H8EzdO/t5RsqOwY+mZt/ubagsc93hTCubXR54ul747VrH84v00Lgu0kh9Lp
X58d0yW48MVlQPW+7y/0k9ks5P0UL2H4CS9nwo0DMUH6ORR8s+IUH2rw9XsXqwhtuEUD4iusYJA2
YEfP/Y/mGychhN/GBWTdZR+Dme68FL6FYPaqCFRpCQweML1hU20JWpJjfzFO9z3JRI/SDvJTSoMQ
TPiSRwuVHL9M4pIRpadxz0Qgkzm/g0Y2nheI0W71oSdMlLZm+qiASb34L4BY08I5f30j3LxYvDCd
XhrP8hQt/StV1b5GEeGY41s0m0/1eIDmVbEmB7RkPKqRo5/wIHJkDHXDtb1GVsw26/mC/PHYuZ6w
feCajKDEn0m0oOHCYn07lhK+239rfKJvM1KdHafZetw6wVK/SbUfKAvzxeArU2tGSE43lzv4A9TC
vnRqYYS2DrBX/MBS30AgS8JSpnTlDfvHTZvj0dFORaL5gpClbI/dasnKMgs0+d3L7/I9QjLLqVPF
BzpSnZEp1syfnnK84TZ8iACF5Dh+2/UPSeogrReEQ9qOt4Gb/qnAF/TEQcPpYlNGDPB8jJhFmnUp
WnfYvOKvxvRchn/Rqd+qXK/kF18EwwLwMj8PWl7y1wOmYqjR0YGiCxavZB+/3L6iZ7My4BTWFg9C
vGJhPYoxGSjDTKjDyCbghBoJDpqv4bfWUy+lSxsrhWVpIhVv69nF/bJswTtr4dguEAhWLJRPCgF0
jVPm8c8In06MJQX/QR213qoo5//Vo4xHnqCBcb1uXzAj7sWUpbYMtN6WAsgjV3u4of3t8XyI4byo
btQ4JwBFwURLZwxzaK7Dnk6hMzWg64Xx2uUYO0WXRKxJtI+E04bdZSGXxxA3XzQO1fxQSC9JlAm4
E0E6FKbiyERJhK84h0EFe+XM6eQQdkYo9yv2kY+5rdKJyc3Am6gjQrH4RPle+U2RgD+XlqK6T6iV
T9nEt+4meoW9zwxVj5yMvhXZyVyP5mbRDu18Ea4tJ3CDBTK1LjJQNUo4R3PAKohiodqesR72n2Zd
I0RE0ODVoj3qdes0QzjqFwYBI8RiX4N5cNE0zUjhDPfAERVP+ZQAZnopZOicEzrIWEzQ2Op+ypw/
fTz7GFx09jThDl1JVwmtcnL+5In+Hpjy6QrZyEUqiEVqxaUZpG8+kV0Z2OVSXk3hlsSPoItqTieN
S09StB8fVEnwG4fCvYgBpTHUGS/r+Kv/YCJcoW71hD1KMM5dD7frLoLji9fVq0F50J3oLB6L9SWB
ZS3NjjMLAw2g3fFWxyXeRaE7nXbL4RJHjazhWDc0OlQ7U/Fmv5KePnVbBvxvdl7gjEWeIMVL1D5g
w9mkh8Z9LTmjQmiCGpZAE7ZWapPCIGAsFHBVEi8bX4P4F+XTNm4R9inUHafG+vo3CpUCCIOLXVgE
e2CIjjuu98zt1Ux6IKIVddqZlQRts958DJwysVxZly66G4ekhnUZGoYEr6nZQIP+BMIQJxc/NM0Z
2eM03jzbKdD0LHJnYfWLDKasiNf0P2IrUj3JC8dx15rJAiLToTPDEBVJng49OVN23VfcM2Xh5Z2R
lEsEyBUCBqrFKKWKcurHi4myZC9WV6cOZLpLiIzDDRTCwQ7w+yLqozZOP1jbbPTdE9AQzIgbyUzJ
26fGC46IhjT/zTPMXJqSWDQDTR6AYieE2SSZHh0/FwsWphD2WRB+rj0No2+73Zvoqlwwn7i0RWVe
PSDjxYcFxlscIce0BbUC71tH3sNqtfhe2QneMPH28X7LGEocMpztoOP28Z3WkLXQJSF8DZk6ISBU
kDL4uExHGvCxJUnka9iR873qiTJHA792Ua/LtHC90H0dcYU/sQ0x7egN6uNiw0XzTnIM1bmcvfxE
TbXR/Jyv+HbOy9wlDvbpy61rDpujjqEf8F5jI3e+i68+fUNNR3vmBFgqC1Ouu8YeS3UzGcdnk7Zw
I3eFyaX9XSDGN2/gln5W7RgdVwBiyBMfn6W11idEMiccMAbxXKkRixLHS5IaBcl0YHCaIGG+Utg2
gTh72qhqNOBHprp0oEB58S/2r+FPkAkBQyg5tce2arpDmLKQW2+/1/YijJ1hIr0izjiexchDiizP
K6CenNTUlqNLv+2+Jg37j89MAxxoQts7zbiXeJcZMWvYjxpYZbKg7Ph5ogeWyDNRRFcErbT+9qq8
D4ZeadaQpiNhUEHDF5YCSwuL3QaM+fAn5viEi3BPT4+kfiNsOAXA2mbzJ7G3rih8jXLrLr+PfZtn
4uS5mobNJ0Lfzx8oSdwZymEUZnWLvXOehNOQheaM4EjwcaAlCwYEhYtxGHMbnQiK6in3+8EdPjA1
+skdR8r6/gdKoyzb040qtSiHLytwMMN53/vjZR80fKNewLOdZy8QoaB3mY5mH0FbOwYLShX6uJmH
GXLW4DKAr1itNKI8BuQsk6ATsWejnagNyH+exmBugrZ9tMXjiYh0XtFXVjai0LIbna8FXOZdSFLw
pC9ivYJpSEXkwo2h/Lwer0yDo6nWO43XG8aQOX2J9P+jRMod2xtNczMnkuG8xOLFQ9VSBAR7waTl
gsv/mRSQycLMDN5s4XEt3i4DOqqKwYs6N7VkQfkXdVt0eyImbwktBL40j+A4+X1JeHK4gyi4b3gO
WskZcPaTiPpAOGRJez/5EB1bo7F+a/lNOe2ZtJhVmPbE9Uh2dZ9U0XZ01IDYQFpazDzFcUk5Zizp
cImpMAsB3Ws1PDDf8bPC4LhHXJ7naJ4V3KVvXfw1jHqB6psHMQMtrTehKDAnW009dqm7a+od0Cgz
17WgPpwtwQkfO2WtthDTStVZ+Sous/UvRAcHIXKE7OXRB/JVqHOJedsVCGgbCyDXMy70DzCPSOGp
037uFDryET40A9GmkG2Gl3zZrT9vD4+2tdN8aGNgUCVjgeN1fo1C6lbwAk6gnfrIG70ZAN6xUeEW
5ECygUimkT3HMhxjlR136Icbifw1BVjlO6T6FFuseSvC0mhRSGSKBZc2N8jEJ5AWbROq/G7wg1rB
STJ+fUgZyrVcYnwlUUKIErke1Rhl7YTxRKzpjfdHtzGDTFMYkXK81OdHBpB5bimlvB0cqmrC55Up
zpcVUVb12qKLSlF3hTKkS+n03G42fnT+/UFq3NaJcj8JsFlHEMm2jMbaBETD45FNNmUo3A/Cbkm9
WPujJA0YFn3kLraLkd4kw+sCVwzxBUX/pqBV54iDDg/akVDw3a90FZAJavQxxSBoLJyr9JnWwahU
WHG6LRhHWvTDUWptsPqFcHAYVnNRzNyxa2b+4cDBf/g3r4mKYxvzJJ75EttDh3bkTAzA6knlVlME
QIZLIhsEtSCSXeL5PbZ9rqBM/qNZilFwlMHD3bNrORkiwNV/PbF4IBgxBZ8s/HgO8InLS5eqWOXl
JOEZR3y4pU/grnS2nDPL+mMlIlJ+JB9CpyjleV42BcwRHlhzsiyke+JwyrILiofSqtIWYFMvdmvf
voOiheVXEVn9yK1O3w7pkOqrPhmLHGT+2HgB1TBe/+q458pXkh58840xsucmie7DO8SeY4e77E9P
+ni26EHUgE18LgtAr7GuFXxgYVB/yPwr0mVsm0NQDXLL+ZpauLEKAvkqkyC9IM4xnKSR1aDnKqbE
6sRO22stVgFoeDswAdVq/ZzkR7q3OLMsqIPshtF7tZye6j9R/LGLW6n6MJdYuI7evaHitk6vv6Fx
gf6nnFUzjPSl6orNnjetFbQ/T6l4rmEEhKhhIJJdoJrHpnHgrhBVq2T/3DI7C3bYePjGS4VTCgD/
EqqSJbnr+/vvv3IRc7DydtzvExd24yPWIHhuxGWFosC1rIfH7BACF368fp3qXkDB/aDCUup7y6Jn
j8NFQBqjRB3ZGZbg0XqUbaZxx36YNnd2w8GOsPC3kNoKkSsvVO9WV6FXQdqNKc7wDU0GLpQU274K
rzHggrfK0V8P5gPsg+2cHHnx/xZ+RBi/rZGvv1kdgDSNM6qh3usQjCo8vb9PpU6bbHXLyw2V3rsc
0Ghvb2rHXL1AQYBvOmOH9/wBsXs/2ZgBVu4IGON/j8mO66GY4Mek2ska13ejOY7cnb14JOw+UORy
FWwx3DiIi4dqhKZZVEGCzFdx+adzrvGyBivY1Qes3fip+H6pHtR+rm90NU5lpBVT3Nfp+TDof3rd
Hq3GFEuQnYabpRwdMTFz+BURPhOocEB6nJQv//BGXnxTvspXdY+W/BRktUOIOVpRxvf/NIPFZp4R
RVlklw0YWb6cA35lv5omqFAnwk0yobRuTUCHOw1s/uD7rtDAwHgknoLwEywHFGcek22CQy9PViJ8
X3/Ff5j/pTWjNViyfAK5iSGLOisk4wBbjrjvuhpSCB19Zj4+OxjNc8LrSNXUmRVi7SQLyvUm8KrG
3fdE9cskIpR6xyZi7HFCDO0msA59N2k+l7zkQp7sJEFUtAr9wk1AZtzi+f1TP7G2WBMNVlG/miwA
jPl1m8CQelbvl2YAUxDcDiXEYXkSgzCqHfXMrBd32+9JZTgVD0m7WzGp34asFI1erLyoKLrt8HFh
UGhugQBOvlWmsj7sueFs/WdQQ3aikcdLNus1Zya2kiuFxK9RA//jYDgchD5XqT1K4ZV6PRBUeH5u
Kx1KTOVlPIsZU67b57U3EMMq/8srgmpLsCwxBZOCWXsVPSzH5BqFwQHdAKtX0MTqRPkZDi67fjv2
zpdT4qn4XBQsp5y9im4rzYkD/BmabitMtaV4d0T0qvnVXkVF+PpYRovJ1Qq90SmiWb8Kvx6/C8Ia
1oWMzFaDgRXbcYtzLq5GGJrN8UW1zL64qUueW/yvJDdqQj2LqEq3aExBXB0U8gC6Y60fWwUDSAZr
2vpyJUTCCQteux+4Go94M0InaGl4BsX5ot76Jupz7ttG9qrLH30bGrelt2P2+GPPBy1CB/6JmroU
9tJzBzNQSc1sJvDvF5JU0z3Y64aX9KEeYOmqENQkjGMWeVPj4viZDUgWnC3mKVYjVZc2PkeAW3p4
PcnQBfwpSwf3nLdn0njsOVokSMOh9CAHWJUTuNWl4EhRbRsOdWNfhULeBBbhsyOfHqfxyqx29pDP
NFxRskiVLb4vefnoDIs+yNkFHS0qpO6VhWkGEgsd2cC3YrUQNuh0dPxiSZ3IcSdfqCwrrU9QAZB3
W5Q1wg1u1L9kLqNEnbPKHWDJ/WmBwcPkgjAm06k4AsvtcsU5ZBa5dI8Vo0r91/pE1UgAmLGiT/nn
QZTUqgOgVyDmqlbPZlJvB8ihAoPkRNvuYUC1qBb2mmkLJDD6yyEECeJj/1QJ5F9lrCU4jucB2Bk7
WHvuFidG0NDDyyJvoStZWQGE0DsLWqpI20Yhfq/Fnm4ZcfEKiyTucRnSEnm7+wuB5oBiLsTbbQjZ
uDrRM2GSWbkHUVaPLrLhPJY3Yz2dWvfK/kXHCa505xhoCeBe5F/CKH3OeJfwE2axHx8P960Y0EtN
UjiBwO6C126lIe38xGnGF63UX066Lk8luvP3nfUWZxpkVVs4fZEkJDBhecph8m54FmD42BNhPTwA
I4ukCebCAxBK2kl2fZOS1Xksmu/KJntuOIF8e/O2rTb4CYwIHgi0El6vxGkK8HSvDM26SFfICjC3
y5gsCXsAAAypUyzgpMuAhGuBrLQj8GQKi+hr62y1XXbn78YS+g/IFPJ2Tmj8zb24krsVQAHPaBLs
Ibt4Ew7FyqAQWV6USIE9mstvUjeHuWohJpvthcnjD99gfIq7BFyk2KD7+2Vk81dMTcdT8WoVTTI9
Dg0KbE5SmjJgGgYCbg2znctE8FZdpk+7ffsGWP4G0hIMYaP6k41TG0bTZl1X7UkTydhkvzXjbqF+
Ob7U2mJVvT3NDW3IW4kYvSlLB5IdLgDga96Gfm//d0mAyq4SciyKyL5JCbTuCmbmvbJSi0PwZSma
dFZxd2EsQpvs61uzExO+zfZBATO7yK1Cf6jeTV2KRgsYm8qeaKlrffpJ0v3u+iA9dOt2ntLRD1fc
S4+A1LgCUVnssWsryZxHOmF98xTfRAWPHqbuc4PzRzkB6WlgnWn9JRZN5qmwDwScuOfiHeHzpAWX
UHeXjZ/DCSkospw3H22kP0efJ8jlh3lnu7EP5YXyTbzs2URlgJadZ17ImtD2eyCMeu0pZ9eNLABK
gZeNHd0rzKST1egwG/y8RSNyiDJu1XNHCtdmF72EPeogbWX0SDR6BUi+qmHxwI+t0ziYyQdvso5n
J7G+iveHXg6lKILWNZZ+EZBhJpfzG5aClt5yk9+sHZ2PUFfJgpYjFRzzjXPLM6aOvUjbY5FJ/70P
mfTn99egLoRXqQs8lr7vkoosBwpPICqIc9oVAPnQiWnU6X2lmeOD4P8iqoiZMOowjtSdFeAkNv67
MDOqmXaZ7cdO/DzbZT/rV+s4JPzikx4N5B0HSLalqaMSc5qLFopEbwgnq1Y+xeJjQug+I/1UshSa
IIcMAsD5ngZDM6GlIw5UGyE9kSr+aoP69k9uIjJXexUbjI9kQA1XVya5nD665xW+wc+dE5L/387t
mTsaofU7MEf4+6kfqCyraQrmZUug1EynJoCzJi+NPLQy3jfBquTxp/DXlg2YVbPVf+9l2hsfZirv
g/ERI5b8DMiEQgjMz8+bQQRizamEGigHk9mdZG74jaBYbA9421chYloyr8clNquyloJaQzJzLZxi
X/O05QANvdbl/I7nz+a/V0Yn4WCPwJxzhsjUjitIPng3zFc/Jc4pzx10pXhhQwEAUG+anvIUREkC
EBamil7Z3RwnM+QNb8RmjD0K0bjm/MhD+O53W9QwfSZ5Yie5S9OQjrK5mJs+QMEvyYJl76gM3q5d
T364GkiZEqKc7iKSaRnhNBt9b7uLpiQjVFDagpFEYarIf86+FOd1/QUUveyMSCp2ztQGeNPKj8aR
odgN9Xn1T/CK3O0YDMpUYN1GZK/F74MxzMkQnOZZbIcrTmZ4E7wZp9nOmLhGjOtaooQfvQbanGxj
P58Dttsu6JaMdfbP0KgW3qIq9O1S2LpGcU2M6qTgCGSvLJC3Vn1dg89npkLuB3nqrebBRlhuPKVk
zjaPRmJntIm84CNG8uW2Ga4UOAropAHYcZD6h121a8D6Hc2PFJOA2lUxWt6nkXRharEfmFOcLkcz
7w9G8w9B8EgBlfSj4oPXIZWkuZWBpqfAhvPxNGPm7YXu2Sl4RPwvHqFwiClAv3iRW6TlAzO3YwI0
RRhBBTxdTmo+y8L6r2RFVr1I2jjTuL3Zxrizcz195c9pYYMwjHblj/YrOkus430NVXGN668+exG1
Vy8uql8q0X4v7DTopnlzruxeeqMCQ1d/ttXqKhQWvEQZTUdLTociDsa/91vARGtrZIQDVMZ/xXtA
W8JRHzcYHlXm6MG4mhKoFMSAPMBffRWd7PguMLtw8upiPegdhmglowtDt3dYugn6EG9oB2P2HaFH
RURW9brgpJ9E7paEdK+MZJpVwRHwmWt14vvlRMUU+u8LHYlvZvbwx/tYnSbqs17wdPUuIaxO/oTt
WXF/OoSkYRt9TaTF0yoZHd7qc+v6QWt7KH0EhzqESFSxjeh4O8nIrb9G/dV38WbePLyP0F07wx2H
goVjwgEDDAVlYiy+eyju6088ZRgs/8hnz13R+Lo/vZc2m75IZTs1tmfA+py7UhZK7YzxDuuTjAsi
78Su3Fa2HR4GIjRF6R0hNl7bOmmTCJtELF5tYHCquxAKg1QjLTFvLhwFVL8U/Gv4OT1hyl7EwAcn
zTyZMRmu0lXEFYPIRfq6FZs0vMGD1i/bSpRtyz/zI6KCbMlTAxSNfi2XcGthNTudTBe4uqjgdzDf
cGPEKDf4Pn+aZ0NsQlJ+B/AY5EkMtBNpQGiIFdsx+enFmH+k9Mj+xRd+iQUYt1fPGBuL9JPSVGfj
oPc7lXYfootr5WMdNffu9Ifv6aqCKROPIhWbo5aqTasnS4xbWBY+Rxhp2nsQF+piuQu9dtenn/Nq
BXpvQvwQgB8S2s/0RBxJDCkVRW1tBJ1xhh3Pz3nVYFdrJfMOdYgo5TRUDmu9sxVxcd6f+j3DOxm2
JCFNw/uy9PLO9KBlVv2y45rn5yAgjf1EcxITzx+WNdaXgO6Mgk+m24vl0FvKFMtXRGqD3VN+gs+o
QaJmzfWBZyY7Ej2Q7cKy+HkzDxryNkQIEP8iJatBN9zggUTcXOoyuHvcLukGa/E8b6VYP9woQxWm
2irJ92WY15qt8YlelYVqnPNfvBziuGsFqZv9P2tZEWeIoxgK9m5oSLPL6PYiHBgzDoJc1RsiHZlu
2noQmrBGdP1NPDL8+de0rRjBtcupmJ6fTRzsTAVvQSjq8gQ3X+BGCZo9Vze6N+TbH91y1QNRPEa0
qSAdPO+Ku39gnxwLK8pGKHo+5n7zEhTpcXYuZd5qX2AetKkeKetDTLAy8lI8iXKKm7gk716yqIDT
6R2kleN9HA5ub77QxDZ8DzcVGfgwTL06cT5xz8Wh8WcMObQXcjQIfqVpt+AWebqperfLBTxWH91j
yYDYBWsx7USYCIx1IbRiIZLTzbOGWNc+klRm9W6qW1IJ6ktStCD+q5JYsCyUS5kFwl3iU+uTjl3Z
kHiUTSnMqib+OaHc9xu8g8aSpVzM9MuLjvU2aJXYbSyFt8sq/rko/CGuWFpSSK8Oek7pnqO8CPaH
mF42zvxWnEHTj7SZGt2JdnHfDOS2WxtryDWUB+8+1Z/ArJT+8YQgCtuVBUe5BzcNEma79ha1eFft
bjGJV/yC4w32TJ9AWQZY4Hrfphbeds0m7O7nwZkjb0Se1XoqNRni+mrDb8jdLWjCp25Vcn6acjr1
Xmk0gwsmvIbxpNNGX7JieBLVAqG0+iuh8bu6MP29UfEMKMr6b5VpH8doH+gSGRRad+0lAMG7fnQe
id3eWxqVYaG7WK24/mwoDvToN8gy5Uo2lZaFPNvHUG2HPCMWhgKdTGjpiUAoamXj298DdbagJStw
9XejT+8QGEFJOWDJfPssFzRU9UEqrDCtaXJRHACrCJipW8g7ojEvHJbWrW9VXN7DqF7vbqiS8NMq
zzngY+2QHzxmKz/p/islBXBFoaa8edtkJbVCixyFWaV4exBMtQxz1Fjjn1rk7jW6TVz3hV7oD1Po
YmRvwO0/7lzsBTsg0FMffIunv1+bcrpJHgHjTK1d2BaKRR/1ZiiaS1IOJOfryPuMqIxBZZOfldbr
b5Bpvsv7gDTPraaR3f/2Argg+jAFA5PHKK6SeUVBfKu1Hs1MQ8fxVsqfZnMZrtsNqlXtEjVfN+Wb
M5sdCPOfoGPsQRaqcVDuU7WmvIUMqNS3sP4HXMI8nORFq5XAhUOgpXyeTfchBmkqCw4y58M9jE/L
SPCJdtodxdJXtEAUWWYTivK9i2ihq8Lg+5/YJzyUonwTyAwt83YVrmpEbIc6ToiUTnvIRy+pmZe5
ZfZV54XyVFn7aXVbIQ93kCkDJDP7ZHsV1qYH+UKEEVuUBNhhJYa/4fsclpqVzYVqfQsGeyTFmiSP
M52PtfC9bZTfJzmsOkT/okjtPFcuJVXoO47Y3WbrgkmPXcTVh6V+D+nZnQoplSHzMO4BtKcFVVAp
4zo8XWw2BAbsrj6Or0PolitvkAFccREXhnKxMStciTdAxsJHbjfdliJRrqWNA8CTdBBXuIzaIHzY
s5Q+yiUHw7P20rgcuv2Lsuqh6nMYU8C/e5FFDhMuV31u+iRwwQN814p/wjoe57wOykap0IqK5t0S
nM9jTuMj+9tj3u0kU+UpNhRfwGC8De55NFpd9j4w5xOCT9pQr9grObn+QI1WfEbYpSVCqttfFC/T
LTRc5xu7Hv7dEkvzwxFPaym3Nm83UteB1s6LJVczBdZ51/08w0HTBR0Ky33hdqJXgxtq01OR+tlZ
oEVrbhOTR/H+jLuTVmJy+6u3CCYlo7SIsOARC04ARWzFcJiVZSN+iIes5hqsY4mzILqJwR45fHVh
QN180zDt3TTrAEe8vpvbYwDapjWpXEqLSf1i3/JTsHm4PNDSTLzjpkEXnY9P9MFaSAWXCQnWinNy
xptzMxcCj63yFaoNEhYTHrMhbwHxJg6kK/XP5r9onHjPDGAjLuGp264Qbc/Nx6KnJ8W4AxeaUJKX
W2T9WjLG3DD3wt+TE84VIp+cGJ+4gZYyGs7YqAc1Dz0MJY+uCzGXcipDaI/uc8lV+dmH0sVWZy4M
LjYefjbQ4rLWKOzxpoXSoGZKJPutdXyqMNY4c64zijK+SzfP845pgHZ/0ZJtX46NE9NRYYtr33om
XvAQGX+UrLOp7cU1w6jOfi8LApZ4mazSjDq+PZsi/g3gjSRA71aGhp3YGQwoXbZe10cRH28KYq1m
QzLRY27QaWoBSF9I+Y2M6GDzI2Sx6nGYcC1xyJp+/4eYjt5TEEtfliCEk32II5pjfNHr4O0e4Lxd
1kVj9M45a6PdtE8ds9V65uCIuz3TaN0kM36iMp0F3T3S3N8Lx8vHFPmbELym+qinjiribJM7PfMy
mdy2fe/+p1X3NTnbMzBcJ/XoaqlF5dRjmSA8aHEAUl0yan/pjm5GXo65O+s3s32EB7VO3NYefD2k
xI37GOWWG86HvN6c5qYWyI0VhiEtAm1VZ5qFt7NI2zJtNBSehF6R9Oih2f3IGnZJ+nCxHumnxJ1O
lw3zksJPjHXADcd2ZYgyNWx0PDqtL53AajPPStePX1BX8kc56U1Hm2VNavsOEiaEz9lxBrkBzvSK
drhP9qb5naIb59r8hVBhgk+S5dPYPA5G1PVJPA9OyWML1BXFUIKdGFqZLXXqhAORhSh99NSHo5f5
PjTM5Qdf4sHJb0krTA72e79w85N+m8OzAfqYKBId/RDSlYSL+94cIpKdp8MML1gJURFImBW/n2Fq
D7AB8fwMRjCQm1I/6Z1Y6p4Il2isnI1c+x/iz/5cPmUlyZ1rbDoVgLYwzAj38eXlkhPjPaagg37b
icNg7ez7iRzpEYQDA9hRJglRHBS5vvdVHqpfzBDrnoqDQWhlJlrLS67sqJreqcy49cgxoP7iB5Ki
lnfypdgZgHPg+tepgw0uO/faBKvr0JWUtu8HarlRJQt7WHN8LaADSGGR/+o+tqQCKYRHgEW4vhnx
hkb9vYXQhNkVWUJKwSo5eh5hUaHrqnyvsHjTOsgLVthP1Uei9jTAI9KO9j/59WoPDuOX3WrxDFZ5
QQEQDSgH3FSkDvoBtArGTqeiLAKad3Z8HB9+AKL85DZLkobOHGDEdXdWnGv5HkBxzODxCgD6Zp/x
gu3oKENz8JbzC92UeXDgC9w80rGV7SR5e3uOYk84q9QvdOCU4ZjnFq6s84H0R42C8TcPJkGgYjVr
B2c/VYOjHmnPB+FN5ikfFqwYU8aFYjdTAnhKy3BNxga21UXfiU5FoHeJQc5mLFRwSK3IRRBBx9NW
AjQVfw50X48V61yMgggckPAPIMCX/SZys6FA3jro8KaUEOjC6SQSM5RND1MT6lUzUvnpfwKQNG0p
5LxnFv7Lxpvo4/WrlodBklBAhFkmMnex8hsEkd6Zs1HDy6xizB6DApTmYp87J24CqcB0nD3VhOvk
mXb3g2EP0v6NiTwtoMu8/jI6q5RCUsEJDeI9eGhijEn4FAIMjLeVw9oR8pZTr2DgYJjt+4t88W98
gFjqgL2/qat0qDsu/SL4tB7JpAe7JFRnP4HSEm8d2Bgf2v792sO4R+0KE3XcBRxgITULBbtsxtuE
wWcWsWUH5eOv9k8XwtWZI+RBBICTtWxAyRYi45Me4oqruXtTewUEnKldDwBYWtXxqn0eT2qQJ/v0
IS7Qg4J2JClJxxP6sRg8eGfJOpkQj31PiFsjYHk4W1WfBXCoqeb7TdC4zIQJ5+pTW7HORgOT9Iu/
qovYORsp1Ig7CA1o7d8AnTXyoTXJFRyGFwnQXYvUmnHiXUf7G0h2oJyVxacFn+HrgJLD+DBjk/+d
aeKbXNZBA9QiLC4L659eZeZOAxb/R9xPUr9p/ZPPQxk62XhM6V3rFAWiwonwSM34+6zKa6BlP7zI
l4qZHbnTf3HPXJm2kqhMP32TgSRrIqEp6PjKzDaGulUMiAXjUzzW0Nj+BU6zugzmP8MIdLHFK0XP
xW/QFfOwivWFQ46yL51N+a7Iqu32vsmGRtZjdkmBeoKjs2siTICgmpZ7CnlrpRDN8GRtXuQ1azmR
IYtIZbW+9kfpjTETk6GKzRxpXUktFYIaRiXgYoR8VQrh4OVBWYANMGc2IX0NfZKRrpH3u2ALp2Kl
ZN039MxyquSA4f3IVssgm2onSmf1kjLsa1cTeFjtNjhkPk3yJEnXQz60YYTAGcWbTENDnAZnqKdo
8qOJT/sjFDEWLSkbsyEIKbKLqHRiXwqXBjVMP2uAZefV8UhLAq8DlmGZW0zoPmH7LL+4Js8xN0Dx
S8uOFZF/8iUQAYwcD40QwUjDQzxy2aj3FhDkLfsaVJ2KyQUUQK3dQJc64/Y9X4bmv8WIj6QK+zeQ
4rMhr5+hvLTr1Y36jscdnNIR3/AC8C8SOB2+2dL9D4rgUlixR4GQOY7q0UmgvdOtnPRCc7ugwFxn
OF71d0c+DswZzeOrh6W6HPomwuHrztXyrIaHi3J5Dzk3AjSfO5WrmBvKQ7oHT4c71HR7hetSsn2i
+O9MP3ayPNmxAhuWU47C4z1Ow5LlFuoHwZecLG4tiMTUt7igWtt4diU7i7nEueC6bn3/5qKpqU44
/y8700nXSFaH9cnvnQgeW0vYk8KWeGZ0YSFscHcMPtObDI4mOkyvLcqVjUynB/qFGOGhBM+fEeLC
I7OLz+0Lru/PhAeMD3B0TIFsKfUgEB9ZibwT1gypv4kTfKp0FQjy2HGtxP7KbA/2i2NV4HtjY47c
nw2hPR49HP42EvUiFgsXWvuUlOpQhmB6ensjAunRyNN+IakPMGdFAfCkhqbpMpyOMYizxT0KDWfx
nUblYpEa5Ce8oGbhjhoCy6fY1p/b0RYZbsmLzbBOHxUUtEih1VqtDd6MgN2ntcfRc3PrYP4w7q/8
SORNMiE1cVniPg03fRSloteF7LN6G4aPZUhqlam3j2ce9SzBqtqD5LtqSOKL4oROp0OVB61Kg0pu
Tu/T7kpb4uV+bFhBZzudJXE2HdapLX4cmGoI59H2v5EfbfsvD1Yvja89eEv+agBi6FA+hRYzkBqZ
Fvws59xUFij/mtKhnFg/g0x0tSvNSZ9A2umaGH4yoF3deHPLVJ0VpvRhiyk1RlPeBQHRhRgMu3Dw
Z53CC2NytAhAh6K3D2PXfqrKB2Yqh77Q9EI8QsINeFpSYbU/8SLN2GP6xDeTQGYhW5KxonBNye/j
6Ufpr+cX2e3JJGlZg1vGKFKpT+ko4il18tV708xGRihIn2BDxr3aXDEVH2j49XTAd+Xi4eFTMGDq
2ekF87Q9qb6kw3WNuea1so4xPIg96YYMNLs4rk1VAJA/jhxlrvwo64fJvb2huL/ywno9BNLY0Kmr
tnjpfb0lf/wNFDEKcwKv1KKMTyZ06E/Y3Y63s4Xl+BBNICRxWpEHFZ1J2mFmXLRblwXtNp5tbFe1
HJz8dgE3X5Dc0Qz8XiZ6vl4GJuz+Feip8DZvSCA93DVIz6es2SuGY8KWGeH3907kQ3FXCnVWRbiu
tPLHTSauphuilNI3m7iwgmAFcHMS13noQNN6J9FHV0CeP0DFo7gfpdxqB9g8KbdkQGadSKn/WVrs
xzJXpmlkXJWsWgtZm2LXpveepidcX3aH6RnYmi3vzwiXguc1W0JbEhnYddRCqhk9YMBNrLRXW7Hb
/9MpBs99Ax6AleG1BgzjqVr1m7H+mFckszhRuMEvaDvKJbrfyHImS8NDb+ZM0HwKqSLqm/3T6zOR
6F/sY+bGqkTw0CiNBk9kCUTR3RbYYOUk3ytAMHqseAY1RqMVtSX7l7+XZXLTJRduwtAAL9MqS/4w
jwtKHM4VMZYp6ifF/KZ9K360SwOCWlJBXmfyR16dGgtm7wuu2MJhvDfyWzsNSJGPVXPrFBlxOtR6
2kjuLbGzmwtxQ0HMzXbtyimM7e/nqlgDD9Za/jEhD29PKvW50TJnxjE4DyLpt8atbqGeF06jAUn/
t6XP2AIx5DCnsobIoLGcxokJYuMifpL+7m3Mv+SaQpjjhcpeQlqA8T3ktmxMeCuZ0M1HLcTcQa/c
uKHmB0MjHOewIBNhY9qjdc9gZRQo6mWe1IbqKVX0DFH9sBJgDa77Tqn3EpBY83vUm4pNr8yoFVwt
oOSGpGbyWjULssEOp3nlHdndKdcI6B6Q5SU4T8H3Yfdod9YX7d5V9gg1nAkUiog9K6J50UWFRB3W
R8XSmKoBxX+Mss+8klY2fIvES64t6VLiaDZ3ydrX1pOCZP2FuZnPfvwWqPCL4mRuGCdINMiOxGD7
wmJsPNslJXlzxucpr3HiCazcMv1xwpJ+ytdo4ZC7DUpURrR+gVXlWkBgrOm/muU/u88tgfTBLGd1
plZgB6WfnX3OpgSehcUQwpcq3ksPfuEOCPvBs7vHQv+ldLRzgkQie6mrzSMEYyINOfMey3DcQ5P3
uHciuyhbNY4r0Xx8ceqEDLDVna4uzP0jU7d7BAMTh9zGTVhg8BkU4pUyueqZ0PmUjpoVJ8GOjtkK
wPD2OZo3QpqGFAqnuixrXTOyOnEgyZIGWgaNioW3PyTGYpfOwCVTQKqH4E3aSOU7pv0icGZ8Bvke
eEHdrntRj1C8ww4tuFuRTZBxHmYHV9gU+6S1kQ9Cz7bdpY6v3krI+Z9Q7tHiF/RV0iD9/cSJbSa6
4IJ4P4o8H9flazVYFNDuQNPWypbe1dgq/ICIZ+rBbutfL2YOrFAEOwseVjkc1R+GHu7qoLw1nSua
ZVG1Fuh+MKVmfExEApuMjoz59BXIQWMthiZEnjybCt9tiZ2eUANDi0v6hv0Zhk/U/cyJKVA9gFIj
Dkb4Hkuw9XVuy/NF6Gi+IvHg3FiT2A824N7bYpY+SLBaPe2Fq8hc62MW/ZmM96n5m6l3yPGelLBu
xI/sip1/+EMN48o/ju3snAHnwCzgG0gYOJQmmZd8aV2YgToc0CEwfk3mLZxkw8jc+TQufFJoSn+v
Vz51btt6Ulzmh4uS2R5S5Vir1XPhWT0c1j1psycb5EgI2/Ej8QWYgNBIXMivkHuM2M3oMbEtv2xg
J3vfpPkRKG0OTbBfIqFBiwqlK7fpNf0x/Q/7isVWAb2WflBBK41tBYnb1Qt8Wber4qWUtD41TLB2
PyIHtRGdY7ulO+lOe9KmAaT305ElUI4b8n8UV/pxbGL0rldCQ2JwCrJZyy/Rbb96fEYJgG326zTy
31JJb57guI91lacnqrx5zqkdo/XqZ68+1JS+8hOprkhBbvkFmqVP7LUJ2ZwfJxi33QYwyoHW6R/r
U3Veg+/2OhrRgwlgiiq6LclJbWB70wUkd33TGkFahPSqSUMsvWLxslXJ8EfixAUOx71xW5dAdXxI
ZaT/7rAVehWZLXXbxOij8liCgb3uKMNIcIQX/N5PVDs7EorvbD8Zep71WaXNpFDQlndQoD4Av9IM
KSavKP92YSNRlyGgF9txEZ4uPqg3zqWGQO/VpCRS2JzVyWz51I1QTSWfowFaviswJhLbgbBDdnY9
Mydxng9yhWcuhFV4TzLDmMxL4retfwex/K3fBxoXwGZx2ILGMmrUWsZjtgmGmKd6cr+tdCout6vn
Ao7UgMn8OEcPY+CwyE74K9Cxfi4E6Pbff+F7Xmhs6wqsp5X6ZQtqWG0PI0czvZK4IclEnoVG6UyJ
MsTSH59UAZz5sBRb8zPvSKIii28jhopykEfHgqBh313XFvjevJAfNqF805ckPUFxUNoLWwPD0/uN
rOMnLL030AJ971AxnziXEuz4L6c4JQwQF+mOkTpYxppRQ/ObVO/s1Gp0OWS8jrbNUCdfFMG6ERQI
2xA+A/dcAIXSQCnZHUSVEavrLqhz7evOjfwyO/3K3Wkog2fatB2HRYJulDRKRW7iaktI/0xT8neY
xrpVclOPy6S45yvulfr61XzDaItC9st/4ARkplWNFhLMeDq/LH6UhVRWxjtjlHJ+92GfQMTJouGZ
jjY3zybUedpLg2k7g8qRpUuRD0wkCbgnE4RWWfZELpstOmq1nbzE/fhtX4Zbs45bnYXVhpb5JxcA
yH/oHcE7TiI1Gw1Myr67kSrzjQrxoMBKa6N9M7c6QbMNGC4ZRlaERZm5OBFqsa97+O3YSTj45f3p
4kCqZvozJxJwRmhuCgEcw1GGO1IfwXrXSrcoExWln4/QPOMbJImYTt7WGlRviUBW6Il8ypRZhrax
FBNHMkF9ro5XPJbtHcz+EJ2BhEzucW63o37GW9uEo1AN+hPoCDtJ1mDtUvTQF8F9YYzPcZ+/caQ2
peAtdR44gfIQEELtlnJ1vXj+0HVp8aN0NO2bntJYyf15oWwQFtAHHjiupp8rV1LY6tIPj7AxKxMA
zKMWoyYg157xkPUnKLdV5weqd43BU2rtyiyY1ukAHDBcroXpI1UyJesa06ldRfTwohEtU68k8nqx
SF1mYS5BWaqkhrk8sZNa3TJlmrDP7mzUooNdC4UHoVuv333oTbPFWb5+KxZwWJs7JfdpB8iqDPYo
O+kaumBMhIQt0v6W6WQ75lxEfnSvhvodpk/nq/74nuSGQJ68mqgkqzHbalaSPmYbNoN+mgLsQVUp
X1UysE8F96CclYttJaRKOh9/hd35DH/ArMTtrARymUc2cwCHEMOnUUrqeg4rC8TF6ShQ/Fwjlata
AS4CKQmPQJ+w/L5EBPluZQr8xqk24QV0e7KxZ5k5ttO4Mk1td3rsRSKSVAGX5kF0H7LIsR8fx8B4
JmQ+lyX1+gHGJNL/7LQCO30t7MkJU5DIaVvKwgpeAst8uRZLAgSLIqDU25pab31ASk960B6rqFiR
Pi5Kt1zBkn/8ktooFMPvLeu3MF7KyO9Xytke76VnsnzNTVU7wbc4QAvc668dVV9f7mt0AX3oAAlA
qsMYNWQhXs9Ofc5HfJvZbG1cpIaC1Q6t3+OWDJBF0I+CqjbgX17KtBQwOEBex80nVkrA0RcpD9lB
xkQrpFPVZ1aPyWgqWUWVEwCg/o38OOCCKFpL8DPHO3ka4gMM+v8Fl/pH+moIm9c3CeaZY5UWq/Du
915nIp9n3YKwMhUXgIc7S5NA2OMcMftrg6YwtLBaW6DU1C025kmPb5ewa0p5ccww0WCWOqH9bWrp
FREzQ2G3zsTxYMpgHF/gBosYtbvM0EsVAzqEtkPpMIymjaF+Gwg8YDLEHQx8Fr7DVsViOEw4pnUH
f5FcDjJfu9lQHCvye6s0xoQc/yRAXL9f9D2UWOgdm/2YDLTSuRCWYwEBu/pkFwgHQyC6APvqpuXy
YLs1panDTLRKSVGWdukOHTh3UHaTychlNPEOpa836m+s6iugHdbScdjJTEKEuDN/lasovfzql23E
g6Z5DuPUaZpcURzFzhGhBljdt3fCXhlLKqltl7dM0lFOHLsDhVHTnUUd3wJY4Kh9xtcIbQgnuRL4
A60AhFLTZ5KH49jI1UEl2eC6M9lCumMLeyCkt8DMMeJ+7umVfgvMzSjzQVp2cDlm/Db1C26tXUeb
jFL2J5C+Iu+gGrQOnWAUvFOVLCUU99S7YBu2xoQ0wAqnjebb1BZc2JR9dSyq5qmC7oCk+3r7iCk9
1qe6HWq5JwMZeMTbQZCI+1fTMYoMmLGUk4emb2sgrV7ZupI5IKNez5LrUOuNutQs9iOT5oSZTlaU
u1/0QZoJCYFBiCtlAmSOrfV161LX3RUnVQ7Ict50JZGGhc3qkJY+0+KIJuS6N+UJZK552IrGoWTi
8EX2vjSnS+yX+qRWZCTRBMFYuvAlCqf41JddaAf+R+3tkUw04W/jUUjoPAq9gU4z0FcL5a2YkMm/
WvNzvYirGPxG1Ik6QsT/nxkk1cIySEouOV6qdFB0ptmZCoRTDFYseNsywzM9ql2Af4S6Vqkxk5z0
rB0K2jrEgeSGQVoEvFT8kN0jE1Z50NgRPcOnCbmk0PoI/6dvY6Nal7EKrKvdKL0NhmpQvSZmhZk1
gGN9Nsf9GGYKO2wQmZB/5t3eZO6L6DAhRpsj6aW7toP1BLBgQkJMgVSdPJEU8p4dihCS2u8pOAnd
udvDABYv9iEtndJRCdcJpunHg/LkXeXDA5vAEcY9/p8Niea+81D3G1r0U0Zfkw53XnNtMphmATf5
yjbnIGEyP6SXn8EmlK6g5+iLNnWKgEVaPIlM5y+uK7kt45IkTb/oQ2qi5e3kctCotq/JqZoiNH7N
rv3kgR9w3Hfe4Ix0YRDQQbR1CGW01HjCO6R0srHLESogIqAirgLVw03jpMCU8Jvt36CIoFatVM/K
9cvtrEKobNY8NqxN9O4Wo3YA71clKNVpOmFLAR3sTKmOJWx7ORZtjH2LvB79dZ51l03Q/WY2YVyN
Kja+TzRrYAZgHqlpDwrc2q9nR9tmOOH8RxQCE1rh+N4QcheKWRUaVwtABMFslQPW1ZjmX24wwlj2
gxZUsA2bin9nI7OIJrf00OTtun0hMW438xmOV70FRWZ6Mitgk1+pz0DXuaTC545VKYUjUFAfAcFm
6IumltOY5MSd4V+M1Nvzzo6isnYJaBHfcMGTdTh3mM/Qpw/ZNANtALk26PTFcSe2OQX4ZgTehvAT
le5vkJmIXUybiR8hi2Dgt5llxySANArKbhUhkZTUPBHU7M49S7Bug61h6r1SaBB8PFTNy9E4lJX9
h1q2qgtKgpICNsSER263YseVTPbikwrhUwUYlT9pYTUNpPShpg8k6CBztZsegOI/lu1grqwhCnVs
lE5AK44OA8nzXQMqalrdavj6CMrh4bgVZNJYz9P6Myvv+qgWseqWkkI7I+qEG6Smn0eVrk8SOzZs
Zcg6+nbA4gesVkckUHOaGJAQOnEVw7lFOFPxlXJirRXHJGv4cs7MWhXBq5+e+dOruk76rm9bhQYv
b2rV0lROnor9xEhSQ8KdsAgIAH+z5IO7/qPD7CGnZMpnDbtbHFdnYVYRTGVz0bOp2XZWSE1bJbE7
EytmUUStMr4wW0e1hd3pddEaXK5SY2iiTJvODe3ESKQn4uvElggZbIK2Gi1fNRKvX+CnNRPacZWk
yHbmezre9OtHLQOYhSVT+9CgmYxZGB2CSFI31bdytHDwuJU7PdC9a06HMcy7ci/JAziEKG9JrihX
40KV1MvmDTdn0f6qSUmKNe+eQ3tuoFgMf+pIwgtFvaBt3IVGcd6Mi50st/2KIhlTRgHIqNS5iuA9
bOAxDU1qrAOMujSOBNnm2+pm2HCdDBQpdoe8fxzRwKWyUE20v6COYhHrjHPD+FLQDNifyC7P1spR
XSWwtbEY4dXXc/E4zL3I2dS5x4VBrP9H8chbthHAkJUDzPs4EibioGRNobZkA2CdVCwTb/BNzHbp
qYFXXbUo4QYbg7D+s5EATgynElg1qi92PEO9pMQlxfwb1i6Nn5/b270Rhtg/QW13pEhMA1Y8BFe3
YTMEJsyhnB0UCJIOFcx18xgXzxjbTjdK3GfQqudT1yMrYxr702dPNPyUJJiJeSTsWzxYCUSKV7J3
lMyJgvFPmTUDJExpdVkLwiYAu9HwT3IG4VizAYzsKtskXC4oUqVd5Yv6jHbEULUlkSV1HbjFfies
kySTQlsphFt47lrsfu46wSUF/UwrYP+wSg/+VhC9sakleiRCPdW7P9vWATEl9wKqoWgKmk5wNlCQ
oxghTQ3bQ2qIcasvCKILz8ln1ztSMFJ/Ku//9wzuC9AaPyUpXA444u0Lha5M+3rECD94MROqp87n
x4Cz2Hs80NnvL7WKO3NEVjAGdM8/kdjMX1A/wTVRRYQP1a1dkBm2fLsNL76j+Bkkhm9aykkDTWn4
o51MqXWz9D1PkMWeC6ZH7Q1iszdxDa/wHIxCBnF1QAsTHzOqbkifodMMmHZrXWJUFv4vjldWEwIi
7k9lRYrndfRlMIK4tW8UNWx3yqHry/Z4mYv2LAtdTvAYvv4Jdwk0WcFurSm1EwJb+UcqXlp+2mFs
mXJB4s1wqkg1xlny2RusQtOtTfFzVDnaJnerl2P16EZs12NcxcuLahWKwP/DVsWi4ZOqiKyg20K+
RMp34PPAG0BuBKGXQ2xC26e301iQXwcqtx9BjTPAlQLTJtHUJyKrnARfu/xtPrmwT0ESmFDW8U7R
bKrSkKr+yz1+DszP2xE7u8HjkPOjEGtAyiuszlAtQH1za/EyTuXT6ygDUXjgS3pyvIE691GBsHox
CRxXv1Wd165fS+oQhzCXZoXkT3GzD0s/MRo7zF0N12n25UyZeoDEUZ2pOOgGzli0s55tZ+KGmtM8
POIV+/Bq5P7b6JhEqbeQ+ZVW/AAmgTlWxHmqup3H6V/VIZcuvYHM2c3BW6Q7qkWWqMVfK9OISMm6
S3XL9hjZ1H2h9X9sd3BHEv8d97CLDRIaQ0IPDBw5TiGx7qExd1rGdovWkflhCQYwCQjZf1lUTkA9
M11f5M+dI6imC/OpdPf4aqUY2D6EStVDVHlmqx2O/6oC8aI9AMVQhuP3JKJdYL8IQjsh21B1FR3N
qZqN+E9qT9CqnUFHViZjObhn1325Uz6RFHzRhlj/1BH8jeHSq5mnfaGbx6SgXxKRMcKHRqH/SSeb
M46fa02yqs3qSERAHEpznhGLWl2LgBncgNjwpYnwgGhGylII4sQ7Opyqms9HTw0VLEbKojTg2h0A
/zUGmpz6Bbf27xTuJY9PIV4Z/GffExqQIFLn19rxQQlJDjpiFGBWygGlFyhdmn8KAHRMoVIJcG0I
l/RjLnQYaG7tFelx0v2wyt6py/3oKaxMESb70L8ZRXOnxv50JOI+8PULcirW1fWZcv1Ix+so7H7A
T+ZAIGtDb9MKtes1hp3IeSZn5DZ+bJr52LWM5Jz5nKILGzPyLynLvcFybuCI9BUtiT4benl2GKd0
t9PPykUToLn0lkAmeTnceokbB9Zmo5qwU0+4AsCgcQJmwBcCC3G+cTN1ugyX7OaXxKgGDntXYOJD
pZjo7yniosgzLjN+1q1ow9b0Ti24GmCybD+WYnOgAxLjLeGtyNViMjeOje6O7kDybn6tCZtWBWMp
EPG33pi67Z4NJ+9i0AnEawUhe7owK17rOQova8RyPEjcqQOlxmtTyuMfYCceqtaOR8aJnjcEeXVX
a9WMCyjEwbCZ8H++7Dx55gl61fHBrTew6kJmmvv/6wmQlno6BYoB1SaGv9xSIC/e0gY8urqcBj3c
Q9kwjU0n4ucMQki9lMzZK2EJtzvFtEcDiduXsWvS8s4rUK6HWtpYF9IM5l8IPzOrqWKc3LA0o9uc
x4HE34s6GgKPt8e5KkLpuKDtIrKKOO3sYEZx5e6EDAjiN6fvNPg49EXfC8VTW+0yeOiytu5HpFMU
bhJYShubJyl1kvUN8iW2FbaSYRBugyuqdDNP0Mx0oU1Em+ZOHPrH4AIyZBg2nt34+l9YXGjtq6Jx
+WnBYP5iYipoP36eIZ9eOd0MfIAOmjgWH51hOHMq0Odvq9b4vm9faHs0+EhLIVj1s5yTdGx86tUv
ttRbDWuzvi0Kx/gzP+4SkaIVu13eSlGzsdPsOytUf8RJ36bebWCKVnWmt177YnevW1fd2JCwBd0w
iXefjsl3QAZeRDA7jxd2Ri7zozX98Bmmdv14/wTR1rAWl7bhX/TsDsFhHs3vrHOusRSYN2s3SrWo
smOKEkGBJFAJmyyMOYhrbkuSAvWVmhtZRRGmlUvNDUKljePJpufvbo7HBJdhqX4igI8ZVOl3V9UP
1zXFLmHb2n1Wd4HLQF01A5rUJB9xNf5f3w0bsqo8KteQ9hBo67rgBZF4iACGALLptfvnr1aN0vLu
+LfViEmHEdoxbFPrhMxmal/w0ym1YQ7OE5QGLbjtgHOlNdUWpvQu9fMAh52XWsBuD47RE1OrwnoQ
aajn2yux8UF1r7dRqSlxsTinozwdFF+u0MeBcChFkwxOROlDXaUWOOk1GZkzHo71ZUXJ2939ei7I
+MIzhkRbMczHCaxzunF9wiM9est6MlmnC+mayBFxxDcV3/T0WLuyn4AQjsWS/UAcg1iw8fO9KdRy
D29UQ4kMt2M3uixoykn3wyQvDKVKAqDh6im7jEVpWXgkmZj5imvYJ8wuXAE33TkkxeCs6AiJoS24
kWGvjucZ/bXZWV00RKH0arjyRnILQDvVHFR3DyxqZm+AFfW+eo8wsxf9IoA7575WEM7bjvFJfV16
V+H97PlVyIAaTgwzx5K6g7IKVj8qUhc0NWzmaaE/LR2UisLJixEGRcRjHL9MEOLHefr6Z/gDGnNz
/m3RhHFSgbRbIwxlYpGBC2kdvhBfE5k2sj5oTk7WalzvcslRAhB7jTHXxEDyARzlBBSx0AYLzsUe
S3tVcZiuX+jIiyAgfBfDHt/SS1wPKxdMBi/OXOJXcAXCw6H18f3FmKi24jRIDAqQnribUpJjm0g5
bKA9XhtdznX6jS7GUJ0+4hjj1qhqMMY5DFdm9KcNuQY7ptewjJF0L7sWnAlJI6mgyUKlelVAVeFE
J84gQUtEG6C7b4q+9yJylVMM4vY0sjATTp5WkjWK0sYIby6wFDx5ybKWzwSo3r/Y41a3k3enX+fB
8hwLLBgM0Qn8SqByp0ZrE/rerZt+UgMoDXOH6ogCKS+cSdivmqMWqPUKMbWkzU5qrfYMG+3PaimL
Tq4Y3scIHtVxE59nP97mZKcNZJ98lMN5nxDtgu/KodxSOwjvhEvSPRR00CphpYqu8vqfX8HRoEqZ
dLE+Azcl3RUkf0Mx9f9hHMNHBdskaq4bUkPs7tpnw2L+NqfXBo81Tz++24Op1rK/9muyGKNdmMOP
NXtwQjaytrQLjiwf41LhHIZ1E0iT5sX/3n7MZ/0juKvbp4Ykoj/5tye/hFA5JfH9CPP3dhyu3zug
7gksVftkEcaMg2VcT6wfT2kwEkLjhAKLpiC3oWz4FNNRClEKUQF0ySS1fg74GLXjHrIjZZmQMBm+
sYRGQ19uHwKtMhYCp7zlmjjfD8NkmZEP//3edWN1s4IqkD8N+XWsmFkY0dF5RIJlimYM+kwCOk4c
2Zm0TkeDacdOoc8ZoALH/CpAN1Z8rr0o9IA6Zyn521E6USepRPFcfwm3/m2xgyIjI6VjIMguyOJl
PQODPYGW83EpIRSK5HUsOYjM1tSM074iEcLl8uhXVd/uP9hqqnOJ0HivnfYgFkMjQuSvvoodNThg
0xHhlsi4mTIF1/9Fs/fqbb7WdF57PPbX8olc8FfpJiZ6s1KK/WnQLuBFEj37q3g9sQbIty18VaF3
L8c9MUuz3KLVipZdZhG6q2ze92I0hwGbHA1nPHGlfDNK9xiuWsKu89aTB9RkGqt4avYKCnyqP5sv
JCxJlGlY9R/VF6/eNWHE1lnEiyLnUhOME2mPWdN+fkokr8NYiNQXF3Gn7+Y4+ZT5C/Cnm+zcz6kD
naA28fmf7tnwJpRLeVY/knrM5ltJY3M5lAWw70G/R0ecRZbDmTF/tINqaS7fZPA9sxt/FaQmZIOD
S/gwW9CNTn5moBxx0n+PX0Fu41tzMuZiDh5LoP+Ddn8RQTEzRdX8unTaR8YuOrWwhuVh7i6UI6wa
td7qaN7TZiS3OzkcMK6H1HRJOEm7erpOdWfsLVH0HSYKEn27oL821gyBQj++Zjv2KKLNDcxtNt1/
KNtIdQgfltjRQ2Wri9OrYUr1IdokmPNGIcP0fd9YUNu63tXs4aecrhxMuc3SGPazOGIAtNXZ/NWz
pZ6E1ShTWP9+ThOSEu8/Y3v8ygGZsLC0by8f01Z15gcycvTlsfqzmMjUqbVLlQwzGc67OGxMCWyx
a5ljD+rlC+vndponRB4y8ZFSoJZRbrVYKO6pEUpDtdGXdM+f/OT5+znLioagt5gST8s11B7pyIZ0
nCRty7d26eI/38J7ELhIO+C4iuiF7wQ18HUXivhCaMzKa+HjTaM4Mo1yS8GfVEYKoh3F7Iqie9C7
NmkFnjKeRVYHdKPNsfsb4LGcEgDfHWJzCR3hOPHBazhIRNxkBs8Kse5coFMxmOI3AOWUgdaq3Oi/
Zb+cms7onnyH7CNiTbm0457ok9M1YchZkrjfH5Ag2m75BQECqMinWz+4MVV8kDY09aDF8fjRcOVd
nfQzW9btmRsAxuEuiagGgkjkX8IZm1UdbWITzjsVWEtzEDWOX8f4rvXBFGS6AcS9hv76c/bSoD6L
2HjGAZ76qHeZhVEK/9+ooAgMbjlEkI6xiH95fK1QLpNhJpMPqZ8v+3GORlKxSxBocz4TJxyaUWvS
n9zN9hPUjK3Od++Il6jAR3wH5cwmvgPKPVL4q0/mVZNLod9vBnZbQVPJyX6E+afTLMJzx2qdv2Sp
czYG76z2c20RtZ0U7Z8bp3WsrME4qoCr+1fccjh9VymbXrtiVgSkQxMCClIVPKTiCYvEnxFODa0M
zS6jH5ZPzxhVkWd23LPez+BxiqN5OsCCMga6P7tH2cU/G8ETdGjj+IvVA5hGgBOo94zZijtA7x4e
MQKzIi/gAsRqZCZ8Q0orEKIRd7lLoGr60ga7u89nW8MjlYbbmE0BwK4e0ehGdnd0Q6v8gRL4WyN0
8gMlhwssPWIv4FLnN9G6/8LnP2LM2dUpJWSbTfZJe2CHKvMEjI4Q3A9GKQJE3W6dcUqqCGveyQQO
ihJjucYb9um+Q7r2futbCnwyWMdBqagR6jIM+XdQh9cxvJFmd/l0WYd/QY+NfiTLmpHSiMl7McAj
+3vqu8QRDPqYEbojKUlIHJ7YODTLn/v7LvIj/Yi9AI1cOqLp3h6bzfgzXAjjVMZBON4=
`pragma protect end_protected
