// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
d+vlu0yPV/0vroTf2jHL6TdzCHEEgimpNArqdWuPYNVz6Y+1wvI120UHYikIwWUOmR9cQyNHU6OV
pxb4Z0LINBqffDd7QWImRJ/BJ2rDKQ4C49BXV0RkdCvoGgHCmOHcV4n6Bz7oL1lQI1zU6HQDopyJ
wAD5nPHDcBLtkpYz9FyDV9A9YKqv7+SOVHcFSUNGs3zuQGUVu5kHZweZdC9x0bbBmhEitcaM1+BP
E3tu7xPFoqPORqTGFv5/J2CxmRSH/G1+ss3kJIEcBXry1htFV5hv8ruB/8u3q8x9ycLuxQfxt6lQ
M09jt1UDQFa7Lx7StJfJO+3l5BLszeyRwTfH7g==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 4064)
mfWfLj3qof0Rnzs2qoAfHY1t9aU4BUBgXQSQLcsVHwM250KPKDi6z9lFhm4sSSa+jwe+pyquFIFy
fkfpYZA51bH3s+L2hau5S/ZjT53gEMV61zy5lK1bOzMGNqofIxfgvdGttcygMmSyC7H42gdjrmAC
+I2JJPyz19eJg8nsXYExCGqs+3u1c1+id6YRNCZ0gB1X9pSPr4Y4Os71xTWRIMF52dhVOk8QO+dR
RtJLZ9ldvaOEaURRmt6I4dBbplIt6dao7lF0kn3Y3My4uehEfR5xWgkkq7wdRayevjT69WKFaVBq
J+C90wB15R73vMuE/KMPxL7mnAHj6LGvpiLU1jUCtGU5ljEXBk47fmANTRnRSm1SpXOsZlYQ09Al
dfSWNe11k225rLm6P8bC3hMRDb+VrWZH6kQ0RKiuYcnr+FTUBKqlgdzsgVQbInnJYcYhwPyORZM0
ji21vwIvkZfYDIgnozxYJ8PMdScQ2A3Dc2V1bK4GXeqH1MifvcoqMXn5nbV9A4x7+qXjZNzULw91
EglzD/IbWG+lC2lncSVufIR4uxf7XhEWn7GICvrzvdPpQrtEn5+yET2K+w+/mNF9egPhnjkcRRJU
vhz567zZF4cn4ZfdRgUeQfEu6vciH97g0RZAjP90c1ob6gnMEGG5lLn6yhWK2ziRSGNYrmD18ga4
K5TzIGBhMYLd7b5swDif1OUCfr+jvLga5pAlvmSXjUrpKxHwMl0Ny0ufIRhqO/evLENcWRBxwFGT
k/0BYJQB037D4U/UcobpMKSISRd+6+PiISPMXBDbiNz8ZSi3Taf0koOTblzmjG0J9Q0GzzFVqI5G
HaTzNk7sRgubbyW3xYUHXVUurkII+xGXkXvqbzQsnKwQvX9PcQKSFCdilGieXiiSr68YfRccPyyQ
SYEHZPAW5ei+Hig4ABMLLGT5hRd8w5bkeImNSsElevCiZlb59YFrsfXvcE/pG1IKPhxWTHFnqxj0
+xLYOTcv4Igph02b5dKGbJLM7D6uXi1i/1dnjHHr+E1d5wvAzNROdewGsq1qynAbXMjP4OfScIiI
y96NkncEZDGnhuOIKo2y21c7B5cBbs13NB+McfGx0BwZFPhTVTd3moa15URVZjE5WpxorHcSGFVj
LmjgoHwhKqeFHMb7Jb3SjbM2huWN1M7/GVZPhpLtZQoNXbifypI3GHWZT046oTKuGvCJDtzO6Xy1
us4TTS0H9eUvVUimldNW7LtUD3pxzuknD+g7gjPEs7JeeTQUKOX5XuobTEtfVnqr/urImiLKhpki
Ms6790FAwOue5p4tGbwUO3iPETR4bKADMOZty5kLdSZqw3wIPBJPHVJnRH3K/LiXyMVL2u5JTEf2
+KauxHcAirir5D6nMDUt1QI+b6qfmVmas0p4UZ4V0WvLJLXgSNlRM2dUl6n0wFOaw6+W78b3hqhw
EZ+hQ8Rgjw1mb1iowjvqxRyUgxhHlha6zubGrLcmd8JG9j+WudiO7oqiZnJdrVdbGe7Z6c7CwCjk
TqYP4BtnQHLFY0BEzZJjudc4CRsecFvSam6ue19CaMafruLGW4DcGNo0itdP3mSYoXNpSbNawitH
Cz5nvGc3ORCgVokpIf6rC6+JFpDsZRtgYK5ry73qNOLZGgMnblozuXiXgqGU1OXiyolu2BSZ3tGW
p//tuRyOa3eZyCo9IGkF9NCyHi6YEyaX6zGXY8QeLQGIvqJM/vR88EwVhBF53BYG7pnGYvRAjtZ5
17dpE+WLw8zM1P8Ar2g2oiN5BNWbvNdJZM/FD7jF7JQqUmPSOmviucMfVtJqXRkOKiyTCmri+9im
kr9k/P7KUR2S9VAeVV/i5j7ar1d3tJ/Gm6zBgcYHiuyveqnyUtA3eHXt8MqAdYiuttIdclUBa9LI
9+GBZgW9Ba0ty7rbT32uZWGDia+G6BwAhDyfqlZrV9x5xYmuUjcCULuPExxvhxnWqTEsQbOxRHvy
6ps1/udJYMxc2tMeEZ8AejEzbRivaJfs5sY4J0VN4IWCd7mKicFztwtgxCQYTo/olnnsRfA/S6lT
y8af7SzahfaoB53Xv+P6DND2teFzWCevrexWTqVuUdgFlpjfiofmeQg7GidG+G0gyXSN3G0uy/3T
zGk8IIN6nb6UqVJMuP8zLjN5Pundea28VyM53AKfVIRDjIY9AEKuFzWzghtm521hEbSAl+7FU6mw
zc2FL8aI/JJH+NCyjbVn4PNeb7u2z607J2eCOlzVJa4FjMBZUDkDQHkuHdgcDDDD2MCEYk5KIEa6
uvyqcE+fP6jH8EAOsqOemrwkcS5AwEEsZrz3cTui6Wv5E6XNqi+PUD/lHMDPFp0EIUno77WTTOPQ
d+aprW8hoYR2WvoluUl+wdcISL6LQwQMaLfdNQxZqf4n0YopapxJCBftnSwATjwjzdJph5jE3qee
0DoU60Rb0LsUCS6fgiC+079u5GRPnykDXcf/oWBXPMX9OXTV7Ph/zuFEwGWAkU1oOoY3Po7+iJYx
VbMjIcQGxpMDMnGUJRYmC9u81V2eqU8Ca9TxvVAgsAY7bazqS1cbMHVWb9z1A5WILNMa50pXHHDD
/BoYScLGTS3GufcKM7fs3zvkLEQxUlleM3ixs5q+MieAOhpq8ZgfCND3kD+hfDKQcIYvbFLE6l8G
CPP1Eq4evCJWUvvJM32dRx+Wt8mJIHJfIvwCGCOi5dhygNzGd8lSUpzep949zgY/HCWZWvQmNgKx
wVh5CLn172PMZlDoOXKhlw6LY98nDKhrtQOUwoWarE55A92urHBMbzdRMJvwllwzq1ICSkn/Gd+z
fFC7Mkqj776Jxfq0MZRlArd9vtK9Sx8dDNp5+7e/jwGxGKF00/LT3E6PA3PmfwR85HqMCAIMsWZu
COLbB/ZDJwlot6jWE4o4wr8F8qQc8nBEuR9nDUTE4hRhpC8KV66YC/hMPW4Lzswlp3jf9hNUNhBn
1P7uvO0kOy+IJqXAW5e+kklQ5kySEja3fupwzYA3UVP0ujLHv3ejBh/iZuYgCoUQlVWDSzY6rUj4
FolgQTn8xETPiCTwu5ba4DPPA6WXsySTFskwA4Maejg+8Y6kj5MxlYnf2Z8eeUEwgL0O6N8mnjeB
/SBYvd+g2Jh6AE922TWDe6PQsnRiamJW9g6cbPXM0M1kds8YFDEh9bAlev2PlQUADnHg/PkdfvXx
UpDjm2gI3FjtwauzNSnwQGXlVutHHLPyU71O8zwmIvPZINd/890VDBmACGedMWtzZzGOLkqyKghg
1yZTDxdk/c73t2+qhwX+Skz3hq8+tyfJDI7Q4Th26dl2qOIJ7lakhcv39tVlnEp/iYdCK8quNOXK
lP2PAByp1/hP2ZIg9LgMaAG6mED0z/cZQ4vNjttDZrf13+40pwC95FP+f7R0o1LplTQE3SH5E7TH
HWFYS/IkM5HX/yGfl88rjfWSFxMJvRdZRt2ZUWzim/Z4bsoazPn+96LQXlByB1b0civeK66dxtTT
+3mUXh0XBhQjtcxtDUagF0z1DW7T4/nf+x4PVxIsM+eHqbOC9U63M1oF2haOvTGetOuA2GhJaaPa
HOTODHpApDFdQa8z+v0h4sv6l6qH1opuKlvagCY5VspvrU12BsnsMxRM3pnHcbQXvUrdnscvZzY0
yuqp3Q7ceCCqn0XvLibBf/C02krM10QKrs4S9rYwQdYGrt6PJqCxrEfnI2xnaVgKWS/yhNyj5q+s
3DFI/4ZeGORrh0J6ah6nti59xvtFBUperRstVPbsU6qZFQBo/YOf2Bxpc/f49gWCFVxvZ+Ca9M1z
7B6OZUA+r8INxp8pvOUFLWiwZXafAytPiqgo5+Ai19zXti0ps5sB+xcdX/DUXksV3FzUVhxWO1/j
/wKytmMTHUKGfGTA4XHWSEgKSuKu4ptp9HO0doY6EJ7U5tG0U6ftNXClV9O346VdJ1zdy3sc7CX7
O7R9nvZHdkJHXE+lNHUrwWn5EHc21Die4HC+aue7Th7Udci1MrXW27ixbPrTmybgfVhxCIQQtQXX
PrWRx+/Ef456auLbp+LrN4dYFj2mjlY9+hhkNVVuIthAU4p25gXdlGxrAYL7Yc9VwzPypdOp3t5e
1oJqRPp4YRx+H5ayICVvaIpM517iDEw523A4Z4S2dinyDpFMAgndzK3tnvzVOiKCk99H0xisAGvK
8GSDBEg4DxrUApp6unrZ9hCleULzoAlTYBWL+mwbHvneBbkHBxw42IyTotdR0/J8oHo0AYdrN52P
6xlQM3tMYKsoWBQveI3agS7nfBWSRUC1GLAmacJLvQYCgAqqpwTAu6Q5W8lLQQ+Z/04cA60eLh2r
iL1OM0LqVtWpLTnVBh2ggBrkbfu++moAGZul4YBcy6ry5Ur/YmzlFlrdyY3A/0Ms3sqRBVjG6gcT
M3+fu3pPscV8BB850S7/jlR0uOTXkswR2oYhIAHrJ11yhgBFQPVpeBPoGwuTxuSP4dAt0osigvM5
Fcl6Ye4qcE8SkrtlF/AJZZfM10c9S34fHmMydYykr8teXWxoVvSkSGv+JnLI/5t/rxgCLKcm5IHA
KsCxLuy3M+qB7yTo8qHvC0OCJyA9WeDktdDcRHLGXq10GupPVzZuEuAX2MBJuzJzfqoRxzSdLw3v
XiyRuELVBGWmcvQ+BXzDcHO/RCEFjneK77mxstlpfHsUUj0ELzRrOR7EolkmxYx14/tH9P66FIz8
61AX/1BSPOPPOU6GiHJuY89XKDjZJC/ww8zqg9VgrPNUykzDsY9f6oAa8Sr/bsGkX97wpT926D14
8OJljQcK6+2xWjQKitRQhT1tZJDlsdit4wsArZzApvIoblVxHXf5VCZig6JBnCjERQlRr1Ii1a6a
sJserJ7UgyuBJNmAZ3GQqhoTxCgvSZm8z2ebZUJTb3TSOrR3ldKGU2F5mLvOXgr8hrQ48FZRaZlQ
vuyYsfK0hjZhPLMzLP3BG6KZbLhNs+DFBebF07t5Qpl35M0rs2rPxiwk6uCd6zoKHZLzqItODMar
B8AgN/Jmnr7/tm2yQTibCflYo61BH5myzH0fR0t90ik7/LlYGAG7O2V8er70bw5tuCN3wAbrSCKS
IYjlNjYGKphotwEUcuDUJ6rZzyzjEf8emeqUuM9NOAAaUqKN7/U9jAga7GpesJhsgroJiHVpj7Gt
iCySJ4KacR2zLoxgh6jUf4jG5BBGnm1hTfe+cvN/IBEDr58e8I8QOL6pzhtfidmA71oHTR8G9MYV
xqY4Bff4QbYInjCYGfxuB4jdAemAVdX3Y2NtdQpQLTIzXh3AsoCZ0UBktJzYj6DAPBWtAt1zHDDp
ZVKh+DzCIzCE6WuZDbcQz0sg1V+uSTWEZG6+eqEOKRO98pbarzh7EuOAOt3t+eTHq920O74w5Ul/
d+palABzLqWIecHVvGyCFsM=
`pragma protect end_protected
