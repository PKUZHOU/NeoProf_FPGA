// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
BcMybMafv0TnReki3icq8+kPUxqE7grYU3AeTiPF75uUfEcuh1tFJj5X8A0h
t4/HtVQ3P8Bz97aWv7UiNoTlK4jGlM86jSqm6nqFvSepMt7YfuBsQTwWXHea
hJBOd1zKSU26H5+zFgVNK1auJXE96x6nMtTrByZ5AImAHt9iMjgDAOlm66yB
Pic3nVX51ClTtxN/celrZE1Eo0qEtpkSR5t87aYOmSqxwyIDHXN6XdSlgUuT
fqtvfcukHSD5urtFwCPZM6PDvg+j0ZRRfHfytwwJfpb8tCdVTkqaf9z36VAG
ZqVmsXaaSUg1AIrni8J8sTp96cfeSMjGIJQHNqgSHQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
iR4FCorNixAZjsElQLsOl/AjZskCnZ4IVursNR3AFtjGVwLAystSkI5kbKDS
DtcM2G46ytgMrmjjo/Xd6aqz7k1YtGp0tnyijMhvt67rnRr0yXdVkUMfPFOz
wIXkCqqcXf2vZcZ9uOW3TlZZa9aTQn1QFIpOLEtEXGr/fLifTcDQYuvFoz1C
UqaEWWwNMiqmp+FyGw0G6kFSltXibM/AJB6s6K8tgyMjWMoOD8zF+ezuhMR4
9DoVesdxM8REf9hVd5xrkPX2hVYcsrXveGrtwK0kaCEUYy3fqkcBFGqBIGRr
O2ZHgHEBskKl9dPf0cL9gyG5fbK9vcu7SyX/JD/hwA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
PiE9NKAZiCUFS0IEoR66GXuG7iJNJDp5EJVEH1V97vsxJ7yElDSPpXtdbkig
CbzBU2N7Sjg8hP/g8eRKq2an40tyvrWVwsXb6FL+ab/vta9Xz14yTN50xwVH
8x7fAp8eREAWtxaAv6MiWVw5AkaGQz9huXHa9apcSXqauWe5jmk9yv5QQsdS
3C4pAoQUF3GdOgsRCQIvJY0ccqEo/Gq6UiEBf7qsopky/ES239BSzqBStVKW
xDbiyFrP+GTqJRt7lDFHohcMFx9xgnLMqsYvr7+fSf9+pAJO74Rs0uMzQHpX
NXXwZl0XtLU+fHKif3kPUe3ACW7991wxE1Mk8BdKnA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
s07/31tG2WyPGDQL9J1WYepXEWleB2CGGzLWIlk8qg4LWqho2mo4GwOfbIv0
+v8yYUgn68Dx/SCrhq4EZ8HCb+DDb/Pjtgw4hTPzJ7dm2yjBprniszYI0GtT
CLpJyktNjmxpsUpVM9SO7evumaXEVqQrAI5eg3On2DivSiOvN94=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
pv+H19FhclLfjPg3kZgfVV28ytF/fARBBN77pd6hwj1yDj2neQ8zzVykVe2a
iCAad+zzMIxUFdVs8l3vO5PlfhkmYQ1hMMCEbrwYz7M6qhn1mHkW33u48DWj
KBQizI7P8pzkr7ZCyG7X5+2deHLqm/z73nUAhfK4dcmfL0IBMO6wBuLZa1j7
VskuQXETaiIm5OxjMVkSTTcCoZVu/lcDVhfARK1+DfGipozyg65cwE1idktF
VuEEx43avf+ZT4jpYyxruW0+J3KhI2OseUPtGGGlunZuYS1tA6XhfthpzEg7
HNyhzPN+p7jbktuNkwKpssK4/WvIFpdLhJI1ZIyM3bGTYfKFCbfUrcwQNq+q
pMTroIUV3fcWn6qLVnKHtF/8eY58/rDmceHoeoMMu0VC1tO1dAAVJczT2yhN
pkcNrjwvqOxkeJcUAOs0rJ1v8Aq3awMnArrzZ4sIYmQdMP3KCyUl6IC/u/tz
/IV6jrHg7b4phXDNRF/suaWBArGAjWJn


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
jAqWpQUMQ1STNq7HtCDMnqS8bOAlZfC976gQldLAgyyes7prvMpK7DKx7yh4
+H0N87eRVuqABPzCTZjsHl9WQzxCgCTGhkE0GlBExxk6kNCorK1AQiCigrBA
JjUECkRKucFqrTK369TbWcoWSoJsAat+OhkwMKgv4oKGNiytkrQ=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Je9hp6m6LMhCS5OT2a4mHkYuLMVM6mK07xdgwaBuUeh0z34a2GQVOt5J8V8n
PEhir2FEnuE1GJRa+RcD78WBh0j6FxHLjEYMr6MkQr9L29IaV4xKWZqvJcRP
E/lgKfa1x5tyQEtHEamrrAZSMX0lCQovyGvPt9/KDmViIjmfYfI=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 63728)
`pragma protect data_block
fJajffekN5kMJpZmDMPR8HtweV4uriqPNVGs5tawmtapN21SiskkbX4cA3Rg
2MavFEaY+4rgOEVafxAq7ITVu2p/SDmbwqFCnIlDm/sE23+UzL2nz1RBzvhr
tQQO51i8n26jW1Lwgei9yCYZ10kKEOk/3+Q97UND1mwEaQOLPILD+V2xPrMy
l17ohTIzd346uw+G3IqvAKbC5AINgzZ8Y7Tp1UT1jndA3/UP+zaOgObq08jg
9Pa/AD5bSPGr4MlqnfYlJaALDPizYJBIbocIMUEuezWwVvWklB0fus/PO/Ur
eYQpVIUPM2oDtkvA8Vo2MfMK2H53MzhG0XB5lEwwgITpRogwl4d+c3wz3nNV
wsEHd921bdBrBGq88mctT4hywzSshKe9vKdposz4nTdR0Wxlw8opdcPzdvx/
4eNpK5fIQdirsFaHmk8JRxD8eXSSJFaZt4nbMyNGqlLSexFiq/KPmiF2eifG
olwdhJyurfPaIpW9nrC4w/WA/SYiPy1y5eDIxqy4DFHQvqMP08axR8T8IFvZ
3+pMCFE04QGpTKzPDjqRlWVIR5DWhlIaC02IXnNsFfJ8cmfA2VAis6HF7a89
3Ybc/vpxJziEXuQpOPFo0brX/zesk3P7x3ufTPIbpPfuD0fRtgeNIWe7KU2F
KOqADFrO8a6RxLItw3KB/ISWETQyWY/MDpWBb8KRdbU2nuN/OlWzSwCveoMd
Xnk76VxWXOSqeosLHvd4znApZBBrYBornKPwbCbXto3sfLPmyU4KnSISkVoO
0T4L+8KqpLRCjCKnKtyf/xW1KGsO9ZIsmtykW6IDcyScKYMjSb2I+fehOVNV
PBbxtGn5cePnRtG8RwPSVEofDXIAxXS5LXqAZaXgUQeY48/tmLLhUYj1xegX
xfgAgcPej2PAgWnLcxS9CLnn93/yXD2CtEcR7l/eQtwYjj1VgEpTXILYnNax
oSYViQ08JN0+C1wjbAjlza2FnABA4bc42vTmtzg8SOMibfaNwQ2grOejXfsC
MwLp8Bg3YsCxL2F3gmkyb8nROID7UYK2r2Y75FiJHkU4FPZCTONZHJsYdDEZ
w40s6VatSDnQXXqxM2libSKZJBSXRES9WP6Vsz6L9pjDajuUERjPMu3RvqLF
j4qrRztrmFiIKCE/0rLjpF/Wm9GGhnupjrtFVTiMGMhjr4TG+hzxzrSUst8x
Ka562vIq3IBJ0L4uqA7coMP1WI6OgOGQQli+2FwGrzwJaRcJuvC8U75FeogK
rgZbdSSUHt2+xXd7ETzbObCNxV2ukfI/11u6BcZ6at8i/wr7GQHQ8FZtj7hK
mEFc9SyhF+iOnVwknIZnh2WcGKcm/njVGbC69CCeJgwFGB7yMTBwvDgjojDD
6kOAfbTBuUT08v/HOp+8d2CPV2ZKgIghkZnrjl5/1QsnDPxhghH/0OMxMiOE
maKcD/WkuSL9Maq+S5WlkcNL4sMG6pV+mmCjjc2DfzCzZ9KfejwQpYqmVDFb
xaYPannW+DhquY4ednkfoF4GnozF+oIiCQvklR+uuVGQi2OeTGxCqfl/rEIO
66RtedFu2yvsqx+K9y2tC2GqDfOE1eHQxJM6Ge5i/gvFN5hb6h7pYONIHPo5
b6zh1EnD/0hjPRpiIkZ+3Uugy/URyIwNuvze1lilUeon77mK15TYZpYgIloJ
uUKyT3x3d8mZrN5Yb8FR5H+xAKKsBoSZPT1vu8enz5JYq8VJ8o5EinesU+M+
S39KYUwn1S/XtW7fHsA2Y16gImgmFCV2z9zbXkAq5q07I5aIsqUh14diFFVW
5Yg04a4Yk2Ze9PCrX/5hYwmVrAdVlsKJIristxhklnRaxIIp3zv/fY0csoKo
KKAy0GLVoEjtPqt03aKRlJkdRBmQP+j7sGhteLKmxyhI2Itk49fkG9cV+tZQ
+595lpAw/17HubUh7T1b5402GRTiFi2IPGTpEbGwldATQwsdrYlX5z/2cgym
F+tAvwIZb4VIXvQ/6lO9+5ysLU/4c6VyZdkUjYPP2BuyHh/Aact/dqQgAZGl
g/9T5Da/yu/MkOcflDL9z1PKxvTjGeqE+6VaxIxJ+iY0asJ+0jO8XW38xzZ/
ErVJKLB/9inOo/YEdpT61dyEK4Q8wjLyGSB1EkMv4vSXHVzZObB6sr5iiPHK
3HFlYeVHxdVWU8mzrS5f895dBvHHRk2rux04K7E4lQisdZHRbLHCwmHoCqJ3
tU9gq7OHFVFfEowCxkc/JpDcj3IoyOOYlCyBeFmiY7K+2/KtdgJ/EQujOCNM
SV8cKZfpF+WJKZlloZqFkPQJtKSbkQpuEE2dJzCZdc7J97Qrd5G3iJGqxeRT
faooeN+Wc3uiC5gTPYFEV2jL80wn/9JDVmFcILdQK6scN/aJtFao1nVx+kZt
HnK9eQKgxIHFdETbAJUmhQ0bZ11W3avfYcFK0KAOJlFOeE25Jv/lnZXOCdqa
S4ZrJbqzCUFx1TVlxBNfSbJ6V2HmcaiKH38Svy2DVYjCbeAB56wkQznZhz3t
3RUE+hM2eOmGiZWsjbqnf8N7s9P36k938fElxkkG/6KajLug/NxPyHLLnp7m
pQfZS5JYsqbugHQWttHM0Kr4tc+x2arOpI+2KXI1SPqP19buGevcPk5sUDGr
SdXwwJ4jeEhPSGzNPflL0+REuYfy4S4I4ebBA64jlskIGB6gUYLxo02gpeXE
NYZion0MT+5TOmrTRn6825pwZ32+BmbgNHDqJjsNVfK246jyFbwGSgBAS7p2
LqoNu9meOIpCbvzttzbW8bS7iq+TK1xHjNMaQquFe/jZQ7ZXkrOw25dVf5Dn
fV5UxQf/E53AHU1Sa3HJqXa8/QcCfhOwQsxLriZVnuksOj2q73G6UIfC4Tys
nr89zAREAkFsxxpYXZA0ysBBNz1Zas57m2c9e925kk8fG9E1sQIcx9DRxhcT
1bCX0UkeWbXVEEEz/x3LwX+JRtZIqXhl/cHX44S4aJqnlJRVdbOH6+2YXLNf
6YoIMXsqJuJZW/jReikuyTGzRtRf++wTSEhuof37+TCPdAUEb9/sGWsfNoaN
T9GdG9wiuiTG19iiZbPRY1YkSSgWaE4K9IXKNHYFGLRi3ggm4IzNsh3LIPEE
Fb+X0gA4XqbMSUP/UNLdI7EGXafSp4wwe/IXVCl5n6Plzq1uassQYt+Ka/tG
41VyQkwGxxp1q5Z+hmLlYkxEROYFN1KBw6y2lBagPX1na3G4NfSDNSPzmyaH
m1OdgbhKQaPZn1D5IT+VkQvYxueB9NVQQdurxhuOXryxZ+1kTkeIS53Q9R0x
aGAr8X5KmIusxLzEy0Q2IJKFKPmTEBcN+HY9cleicqunaBM/ZkvCnw/6p7Or
VZT44XOcg/jVhVmonRm2IYtU4n9CfHA6NWPq7yuvUcGBcwaJBMJ2R13vosqB
g5Tl4frEHQQ4bkW/Z6sDYkGq3D8W3k68P2XR4kU/deaKS3Jbf75HxBfpx0EM
6IU6d/61MQIESa7zPL2srtklWSCNmvZkDTp9n3MX/3B7CcuZ/sdqgdZOYYLh
AtmqsxJfGkjnI14rLUwbGuAUcf4WoUsnAEJzQwO4SA413icDCscAf9ZUGcoO
ppMFNuQVHOz1y0ksaUoijmVrPPvn5T4Dw1SE1VR8KzfTLclskOEWqmYqYfnD
YnpYDTM7eEM7gfg/Z5n3tsGhKfjjqTOhlrl56kDfB70Qvl7l7WKS3dDF8Lkm
TtzSchV+nES4yhCf5+pjmhN9YqP+cHwfXXi/vEPlZLpx9EG4+u0Z8B7OH4fU
Umu4ju3lHhEThKI+v2ZvNHX3hpkhJWJG6prL0M69ZZ6Y3LTSJX2Ws0y6M0fo
2jB8Jn+0yM3ITWCqF7SVcOXKfKI97GO7jwCzSh86cQKo/a4eggTkajelpmAN
HYcGo7F4eMU7QV1bJLs42/t/5wj+JdjRPdw0bq1hYfnmC8h5v4szdI+sM8qh
1niMjUQBKO08Q2wQU+c5cfT3IaU+Hnmt8QCgq+9QBJgxwrzjtbvqbHuRdQ6v
bQ0sYjvVqTr2x/oE/D2UtkdD6sooU0mfOFrfhQv+RrBB4NWZeOEKJJHPahw3
Hf0wVuRCciclvjARwTyMtTshdwLj1sm3ZSXyz+4izq2ZHBuJ8/OQwcwqkc7q
DOKRUSMV7+0pJWO0TOyCpQMj7x5pdjQabQS4Amivp7TFNw2fmOibn+ZSKi6S
UgX7WXVI/HYd+SLKRPdSRZArQ3wTzKJgIYpC46G+Rerl4wcp5C2raQog2fIO
iw05u1cA6zQ3b0JgaETJ7M/VzErGj6+IMC8QdY/f6QyBr4+n8JAkr0ObLMga
cinvuCiA7HorDwLpL75SGd2QyRiNhzK2japn5qefUBg3gBfpsPIEBM4GepfL
xK8JRQ71DsiNTKo43bRK9f9Nmgvf2Z7rPQ0qSIaL4xLG2ZAZZJ24XG0TIDsw
dh6Z/kPQvkePAm7avsaSP2aloxXvJkQFoO4KVRIgE8arz/X9Sfw1KT4GiQck
NCwS/UAPVzJG7+4/XwlJ3ERRLlr2KLJeRQFhnpMfri9vwXuVPqN2wJeriSCh
+tTGbLJ/E4mt+KGxCPqbPLJVIr+EMBQb9rdeVUjqza6rGb1j8WOqE55E3/mC
2GyVkaqLGXidoGXgVFHBjuWC9Z6Q/YU4rSaA97L5+WGBn2T/aiI23CAblt9t
/mkDK1Q4/oNFX65gil2pcWGPaXIFjwZpdAY4nd0QiwsrDQ6JQj4/uTw97AvW
Wgu+1OhHMGyxyOHV7lStsEDcpYGxIWngG8kieS147fPyl3O4cEEProRj3sK4
wFdP9zWhSrlFBvUASV14E3grhZV+dvgqE5D27TAJJRQOODx+gpLJrRXd27H1
5GiSr/GfUM7INgOkxMxCrEbi8F3zEb0q8BtbxRkpP8oRv08Xx4+zvJM7pXYY
lki8GqjvquCSzBoCSQ0sZ4klfwAN7nK4W1DOEwQkRICHqlJDG30z08r2wsWf
kJLBD7aof8PXfhCqY4rT8hb4D/Qjeky3nH32zrDE0t0S0qz6dGe9Oq6bnKz/
iRx7C658QdRRbtkXQ+kqCfq/hzbYjIxy0X+eVJBazcvhs/oyjpmzqbsGlrok
UAA0tSA/y8qneO0aaWDJNAsp/RAXrfRdTY/GGXWQtHFZ/hofnhZxXvLhyIaA
sAfPPQB2jwXUtVGsmBMEBeyYsIS5g040dhLSjNrWlzl87RbRMAtULlpZnvyz
Pe+R88+dnTzuV3fG0JLocw9JuLegW4uE27CwGXOvDIa/iOMCHvPSKM2i/h5h
rhmVXCJtGPY0pcHB249QbMcaFJytvdDKHQFjFRKGxEVt1fbCOUCLLHvYZ6dw
sYzJ0MquWPs1MPq11TabP6rYMg+ZvY3Oq5uxHQmNC1MfxFZN8tPS+rmXKesX
ybZzhVwyxy0zeamAos415GnUNyrEupw4A3PBaLrUQ0lB7Rjs95daaDeCnnGF
uZfW/pIe5cM8+nZ00+fT68l97J43mjs1KsNsX7NwWexgVlSCc09gL3e3FJsZ
D2RDu4iznYmn0dSYkB36UglvWTmFf0/sy6b6e295IrSHUnv0YyH3ue5RKXA5
wgfXggXuljLRBr9rWlv2xG4oHw9eJD+Ul07bLx9ls3b3Zrq0FH8Nx/3GxYCh
fxqqyfdYkMJV/GQL0quG50Te5NnnMc4HWmL/TiSkl01st96rEP+HxS574SSi
4hLOdZy05ckrvMFFReHFv8SrOyooJqPC7vunjk+T5p2AHGjfPtzkEkqId/3T
vKRnHTt5wbRtRn07mtqQGne8JYROA0WHS+N34xJhQgmD0/76qSvhAZNuk1F+
Xyi4vEd+qiJ2ovyzagNVGPz2MwJ+5ftnnc6Qhqy8gTF21o8HmhbDMKKZl5v4
X1qQBIqdRIRFuk2dZrnURK7ve10xO6LoL+MtpXI0hecIyYBNw8M92inw0gEv
h+Aoj/kcy4+pSDh8UJlnUQFxzBqN3d/ekdLKor8x4xdV+TwjNnrtmXOecXcu
LKHlHoJOnxbuc/+ty2TkgbPSuRPGOuJHTZ2BzaJwVKLu3mpFGNbr8/yz3CSa
uiVzpTvMyhzAMMsk7eGbd3vxIp40n/4a44f/MMXkSOMNkhFqRGJH+IL4bzJv
NY4PWZ8O95Sa/o3Yrl2Ru0zIMhbhLlDs+tWzOpeuCPneErlJPym89t04Kfq9
tz3QRCzaNBQfrGWIZ7OiWXwRwqEX37YwDPfTV6H6dBtgJIDC9jwOSsYhf6Xz
C3FEpjv+htgnoaaE3I6sDJWLaUo5IOq/tf7wuIfqLepiHaHjth00Z+DsQ/HI
U64tPzlBmaTf4u1ew5AMRGw8lBM0tkEHNcP4pQugWq6Au0c5/amTAjdRVITa
g4CrcPYbwPLZT9BDZOy1E7qe7sJNM6raUQkRpciXNRb0sLtRWzwlHQqnndwI
jPxwV8VQG2CJTE3+Kom+kM3czY1UrykpG+xvCrqY6I7oN1ukzI6HcmRHzFhQ
OZ6GV1LRLnX1hA227ZSYAH5nlwwbYDp+O7zbiYdnj44WhNNWADZjvk7Lclgh
DZunDyHveRTsdC1AggsS8XKl60+YbNKeXpnwWYib4JAjN9zBM73vY0LLav6u
FoM+3RarzCSUjtg3icZ+eqLokEOMmMmSoqhI3yvYSIibTU6+sMbuFnqRWX9B
uNnx0Iuu67wwp/kdR7T7H7JgkAqOxHp07b85qxug/brBVoZaLf7LeUNp2pRb
haveGmQjyBcyxP1Q4xLogKTBl+HlflnpWlVz06Gw0Q3N0YfguiaHcixADpyW
zEPgvl+r5U3Wd2URBXUw52vLx3NhJorkbHd4HHN8OPdQXKftt0fGV/+wTtTr
XERARgAJWli6bnJ/mgC+1obcNI6geu6ERGBh5zldisEyMuoZyHIaMIXBZ3Mx
S8kF7s/9+D2jrVj0PLy5MQ/GB5mk2IuMHsZQBJiUO2YDoP7uZM2Wpo6sl+ow
1jF0MjhygKEBTlDtv+ur70KOcN3RgrFwWqcWeSv4zZ/ejPX5Jpf54w1mZRd3
oe2yEWafJTb9OKerXkQN02JxcvJN9cPa3ghyv3AEmlYe3tGgFKcZt6OWrWDy
N7ujBhEgFZ7/IrVwsGNaW6RF4NaaDxMET75DVvwmLBX/qS6/OPRcZwxNhfZ1
sjpHQEZEAoqmVHFcfUIlZIkA9o1MSJLa0WBQCxsWMr/t7KD2qEYEug+5IGef
+ahCqWt9QhgKV1aSMWZh0RgnmD3UJtPyHSKs1EPupTOQTOcd2VbNJsU73v7N
izvQxz9giGuUf1Eyt6dfUS/ebAmg5dWZ1/xrOj5hPQkVn8Wh0y3L7LBPLVdJ
X4Ij8copwAfKT//AK9HvJNVX81ehu0etSMiCbQiBjar2jo4tYza+lRM7htIS
5TevdlPlI2JKFjIR7Mha7i7e1WiAY5T81K0RKYUyWYPo0wcE7lERnFqhN5Bo
saVBrjQGK8F8sCiannnnQ9ngl3gDmrMd/wX2ObLx6iYC2hNHxd5VMGZ09JL4
RiPg8tPTb7Ye0tUyS4gMQ6igMnHtsZiivuxk9Qhe3bCBOjiDDhTkkKdK9dKD
+Smo9+wPE91uQiOIemhBVQ4++j4AkTWmsVPL+qxqPtAX0JAv5iIVzu/h1DQ2
6Ej6XL9kVvmz6gurw6YuqSyVgpBsY1lUxiPqnidkLKYjZcFcVe3UGut20dLe
T3xLzt8I3tYBVGSn+2b4aW7aAgsQeYzHWbm6C/6r8Z6SWr2CiJbdmaMU1r8K
d7BQWSB97+1Zmjn0v/TWVV1noCecL3OELPIoVyuZuz4wuejVR43XtVFL1iw0
grnYVr5ZaaFxX8iI1C3YHCKepHJt7MaCHRT3cIt6gNF6KvUUjCsOroQkHWhs
wbYdhPcW6ydObqp858LTG0zbDsW1qZywKxV0wG2+tD83dziA5GJb9t0pKy7y
a5StHy2TN+DUIBNAj4K3uk3PEfmfEOr6ki6JFTqjpGQYyzBBvQ2CmTOI2ecr
dsb8z8RRtI6gNOayaMAvot5Ba0yXeS0NFQsZ+1x8x5Rh3dHmoWjtAQO3MCUz
DnReX6dBUM+aSXRIU7aEm4g2NRuMR9FWUhcVbkp+q3wdbxL2ZTAjCelRKu5B
jLOgPPin6rKnkyy7xYnlWmpfu9pWbZoeWarlj5COrs7QtdZao5IiKBbH92Vz
prevb2ktFBeXHvNT0CgChRTmVbmgizQVSC4wIAjj2FCUwE8TFa72j08C/SHo
EyKi+UUnq/cjiJ13oz/BKzvHciip6zUOEcdHRR2DEA0cE0BOZmi91d0/hSGg
F8TzEzUqsomwbzz9YWiQg3F2wAodAqekLfqUcqLZZhWrGRFf6lt62M4LPNWt
UBlD7915KnlsK9nEgHS+g//8073zA2d83quqv+LkbM0flgDLI1vgRQ/1a6mb
DVR+DGACuKLxXvc8XgNrvsk5H++OiLGBICy9ZCJ46QPJxPhKRgviEhcbaXLz
5zJFTfewipBEtM5qlLKcPEwsIKCzh0AY0fyX40kYT3gdMqulTk/g9PU5TZhg
032/ARKZI1r5TK3U9IBDGddDEQQSwZY/ULWFLgbUFZrDeDzLThr2tO/7lrDQ
+CKArpfQGN73MOc0kRRvfth3ZD7CGoB2ONfGU/mGgtd92w66LZQMbtUZdST5
2GlQZpY1xLYT9RaOaRYtl17E0mZyyUphEArzBcMK+Jhy8qt/TjkPtzxoyDpX
4xL+TEVlR3mN7wJAdE+AoAif7aWJ/VC+A/ZQHlemMqp5uZB0N5Dke4aqH9xG
DCVdv/0HgWvXLvb1TxfYbVKVWNM7t5g6JTOtPpEZPTmenKa2xdu3M/ZBDu3+
rm0FD+XHEUInsAzg+SLMWc5Gl5/zQS9HJtOGtfxW6Dto/XNuvZavGR43yR8z
RBkLOvNG8C/SceA54MajRjtHsGnOP1VuhVRG84gy63w49kZ5EFdW0Z9OFFJ8
pOtBpdv/LTKvolAVQ4QAKaj6WWHDda3l5lW6EZs/vgqWTroK6AeseWgX3Xkg
U8B3FjSK3kvjmEsv29HDJ1sHHogbdWDdtmWx6rJW7jmsvgLUOc+tf3qPVDVe
hGzwMRdZmQ4VqpFkQFLk7wvIicdU4DQlPXa5GJ/EncF1C3mvjt9x5j9ULs1U
CNvFXSERKxiI4NaXqKNzfzuXFNpA5CeIw0cYFmQEA3xbujNpZYyLjUaQoGtX
3iRwntlrKWRJRxsAk9Nn2uEzhx9VXqHs45zDngc0c5OsPR3n4GMMHCkPU34B
ocwMLkr2gLSDQIS7rfZHpUx15Iu4XAAZSbUGqKz2QFErOICrTGvjketFDfFI
KufsPN5/h2AkDOTiU9grxo7E1C3X3biVpKet3iGyREa4P3DrhSkFGIhKqYVW
F1Vu7bwOZM9+b91S7kl64xMktcFCjG0MydXRuQo4E1Tk5d6u4oYFVivOi7X5
EKVL74bcdJOb6WCNB44usEyFlikwVGC68Zjj5VPyTNcXRkQhwgrJQtzlOL+1
LNq/ihHGmv0btJxroBn9rQB9+G3NCLWl0ASAJ6KG59EjiXseUKtBfHVbWaAF
N5XIZppuvnmN15DLl+LZbwA2DtLf9R6Dg/X6ippdZxNI+EuDtjT3QEAIkft/
aLJ45AwSZ9l7DucqXSqcE/Xy6ylgK0ahf8SaFTJ+H4OThyzTk1sg15NK2M0E
eRoOZ7rc4av4z8DH0Qb96Y1WD2Gw8Yki50N09raEFNh/lgcF2dR5K4HgPlvr
2UwYGFEBFPX7gNzco0whL9wI7lj90891cY6vavs7oyJFPZJc2tCAig1tELGz
7CtPSc70kK+1/YS/ntST0epr1JvZJi2Qj6AVXKvPmFDfxmjp19ebA62i3tSY
x9xLARUi0kx9TRBs46h8kxjR9seMm/QojUkPYEK9eTN4WqykHDuS7qp3YQ+s
DeRR6imgcCEyJCmmDv3TBt/4BlBmI+acvm+KgTsLTKC1fqlxgBfvMjn66CWF
3/lrI9dFpTEeckESZcc8lUIOeDDcsAX1lmpoq56FY5WjxjTEk3bIiejHnwho
sv9e/jpOebwcT7l0QPngpBFEzQPBd8ygMT8q7kMuAEpAiZkWYaeBLXv77Fev
GIOsEv7PcTknHOtM8yvTQE6m9Oymhcg5XV0o+xJQmWGaHwOz6WJzOr2gxWxq
faDpUXaxrS08GLFT8uvA+mEWnB18rXe/DmvxMPW0Okp2kH9RWxKNMCvVBml2
WsaQuxn+6lbGRSQUHtkYoMzWWZiXFBsT7vxWyjFn0Q+cX4l2Ji8itWtOWOrw
u2Bq1wyIDqlm/ku3UlfJgE5z7SQzsK5UJ1fIqUO83XLj0OxsIwyj0YSdVH7p
hgV8wVnVwKmpg0qSM9TopP/BnxZEn/mwhntYAd6QjCsTCTe+ATL8UXCCQxTa
un+W5U4sD/4/Fp5RpXXYwpalAk+hBpnvlCIHwG7cHszPqpTySCnoK7skcjaf
AGK41ZOGVuCa8TjarFeMuW8FR8E069Q8EZSoZ1iHTvO9DDitzv0voY3jZy8W
2CW1Iok4gO14uY0W/uP6dwR/RGPWinlg1Dyc8MBbKwSpaRm7PMAkHN0NL2fD
KvZNRyRshp+rLPnT5Y0aWqmJGPpn4H1iOoxXVLHQt5mHWilhh9s6fhoiaIxG
YAmhr8I922gVegqmOjvtcIVVKmyYfqtOihYnWWbPmun/Ba+NgPpnvN1DqtSW
z7Cz+qwgpZSYvPJDsh8f+F0y+n+xDb3+ussOhKnKoLHrgGnJLxiL/NH88rDY
aXqWpfb7g/xt8aQo5CEvqsfz4VnA3uovV7LvdTtg5RbNJHJn6U07qOK9PXWh
iVBE/vFcu18ljr1rawxHVmmGwsHaVo+/CuMhrT43ZQ6IhC8+odEg55DdCuw+
niQp+TMThi8z5+tXV9EtegQFy7iAQ77rikuNWESSUTTM4bl7s9ncRkqQbSHf
iaw9uCScCXUt6ddDwlxwMQ8Np526lvw/724XrcHQsRor6wrsAlLnZuUudimk
JEw93kfeMqj5EQkk5qhWaK2bcy9g3FpaFtjGpQn/VLeEnWduYvisEWtWjX2W
k0GmvILrTUlaJ4H71rPuKEUhaaianXqSIIPSIJnN5GGqNJHwHAK2hnlZW4ez
1ihsnFK8+0ZsFjK5KniTXq4rVHXJNne8OJauEypa9YVCysgb+CXs2hX68xUA
FQsPMIsWyJ8G9zRZFYqS0HxrWdwpPdJQhoSL7+P/aB1nNhxeF1vCbF5rn3Lg
hjCb7dKtJyH0zEzA7uOAeevdKV2WOfh5FJVBiSw+TdX55htB8IE9U/CYYk1b
+R5nKoEtQ7jIKJOrR4X2Rc6QoPM0wKeUBEaBu7WidwscjvcbnYVu7UUxt8hW
vRpIBg71WpzQ96rERm5IoUgS85am0wlLp7xctDnWFHfUQZ+rA0J4SVDAKKtw
H35pMS29gMN7YA3NK8mC4FDO7Skdmgh2bTiYRL9XwOUxgoPfrKuKoEHVoO9o
IB7ZiP36uRHe3RSyTlTP31CInZEe2St0St4D8CXXvkydGBBHFBuBJ2ZUT6yv
PGiU/hOkBN9NQD+YRCUsvt7JW41QqRmTChzt4Wcvxuru5ZYE+RENrHagtBRj
hjc4Uqc3zrTs99FIjS4qpQwaVrOYMbgxaVNooEZQdMYG35kESPkuqxu+67VJ
KO6ts5dQrMXr4KtEy9VdcIARMfTv/kLrgNnOtOJ2teOe5iLzn8lvK89JvOpF
unEih49xHg00adCksoZ5F4OJxhfG7noLRFirY1bwaeLzbFBCOmJ0ZwNORsqj
AP4DtrEc4HHZY5Vg1+4g2nNm9M6dNRvAzuhXeujkAGCF/VMtUb1XpZI/qZMS
fskyDwqbhHK0LZj31+2seNjGPP6q6VBRZx3p0HIouKGirEI9qUAIEzjs20SI
7WQj5gOJK+qKP3J7PYYgbPCbO7N2AU1KO+E1mHOaAX/twpd+MZxZ7vtQj9LW
msm3Bfu0ddl8vciXLzLMFRNAkbMLDt+Wt4z6Bc5CH/ccml9p14426kFZ0HrR
hFiTq43Vwlh92oaXAL+/KNyTuiIrjeaDbzWv7seNGbQfn30UuXZ2USwID0GO
W9STRSZoTn5SvwBXJmkWwOvVC2f01pDwT2j5YKd5U4d/lVqlj63yECwoZZK4
NSt9VkAiv5LXEITshfs10GeIijhgYiebhNSnKqyiFwQtm7ZS1vUaK8nugsG9
IsoN8HktQ5SHbg/dtgPTD4Nd2qWY7qHC+4Q5XTbr86XrtrofOTRNxKZNqAdd
7wPLhgGsXoys2+7G8Ig7B45yNYizbXYtNuQeecEXXC4D8MVFs8EeOCb3UAz3
DEI5vO8njeb3Ivq9GPjhxS+E9/rAByJTJ2vrsuYz2E/42a2X3AbPqGZ8iisd
81R4k9uyxY9aN9mD0RALu07u0+K++wsmGCWzlm4o4ohVoRWkzAoGswsOq5o8
VyUW+S+BxcsM2cibp5mDkABP8nSLXHy3+JCCSEfRfwICuT5VgcpkMFmY84yv
4XmcSNkaoRG0Hz/Vz2PDU2gvfknK+0LyIRL/8HjJQ06qhhppAzoLBs/Mql+x
pk+Byi3wByLpmCBi3jSknBuRhL8LL8lSIgA7rBWhCrdFrUK7H7paL5qHJApq
fYvTDD6HqIHyvaLpX+elegEujpjtv20DCEtszNuIZYuQFxbDpcEsSdhsU/xD
aNM3V2ZzXKD1ajmr05y07C+uGgLle06/1vq/Jn7xBg0ho75wNnTeOukirRgY
Nbrw8Oa70266p9OYBDR7afa6eMza353p5S5BKlvYVfC+gY7fRsSSnMuMBG5b
iyam4RwgD6tSXEgNfgFNys7X35qrpIME7qe2V7/L6V2WN5OYyszULqwzXTWE
hLHDrWPbWTEdzgmhABTWrjtgHSjtZaYdr2TgvgpPYBeZHI/NaidK1sxKO7qO
+5Rd2Z1KilwhEC9A8d0spgiRk916r34s7lT4bee6qj2s+lbev5e//0KzHFEK
k/PxCJuoh6p67+oYX44GZAGxkyCILzejQyKYR7oXyP91lj9xx1hHEwwE1Q3B
n2x+WZ8IaRD11oy3qAraQNjHWD0clkLLBFDgCLnyEdlwljJgMvUQtA6uctoV
7YJtn5Gv2ysliU1tzrK3MOKLzYdB0loeicXBoIpnI/sp/Dk52LXxrIXMGEGz
xa4xyMPBmN3Vryve7+QAFXOzr434R6G5LkuzLPZgBFaSiUqTYh1jGKxLFop1
TGyKEvAdWp8X/clsML1v+MCq0RH67YEUwZBTp4ODaJmC0I+RfAr/AM0V502z
auSk75sVN6nfXI9iwjeOQGQkQmUQpSKXa4KKIRhwu8Gj1+5X8isdvbGibAaX
aHRIdwP3ChH8QhBz6ishzdvfR/eZxuAIWLyfoqnn8pQndX1aJwDMKbOn3Uld
jhEY9hgfW7S8fjykwkjdxi1pgoxa821FbxZix2XEqItuU6m0xRTvd+EwouoI
+EKE72LFuk0H/+m/P9/fe6mqJiBIgjXfNSwnxDldojejwcLDcEEPJkBMoDJY
B/kQwYU5qK18mNfOtbXAXvrjbekcZaaiuGFLwmEw+8q6hrZiKvI26h1Dc/Hd
HsbZ4jot8XSVyvEokXQmljKgTI6yuNjT4652zw8srSKz6FQ/S8NKEKVobvPQ
kHn9uweXhUDMP17uVYYlZouhWWz59+4p8xDwBhWbbpquztnEkuMKuPKt4Pzw
jnjxWOeejhZp6SLNfbdecsprBEoxnJt1drN4+xseAoy0sZNKGnFgQsnukZwc
ZZKT+tgDYDvqKm0FdIpE/UPO6a3fuxFibhdJXdBnkVVlXrGJtbz7Hs8mvMWj
u3cS3eYSGP0tlElxBYJaW5UZ6vH/Pt8eD0DA8rQRG53fKFZbh5PFnUHt0U4/
gRkF75NI+fRU8fnT6NCKDXJFaumP2dxvLOKq2pWj+jxNswDPNPfnfsmvKpZ6
6acY/E7wDJSXeyQQJlu1eyY9GJBBGIUH1UYWCe6+QRSIlecDQ2/j9zl1kJ/E
wf1yopktnZa369QGpNzCPd5SP2qcgWJjVkICFC9/PD20PGLJDCwTvvd5vrZu
RHAdZDSttE0wLRol1z3H0U1azSbbkIe7iunGhrp55bNB+/Z10EEJPA6tm5vt
7IJaHsmlCD1bV2z+CgEIdTTxJTl7Q1EV5tVFDPDKUk+nXJUsZ16FUovlFN21
nXvCPKnXMup2Rmg+ULVFLYGSEP+msArh/9qqn3zjlqrYa2kwGP3A1lerOVat
6PTbTw2AfN0gwLNo/XG7I+KQEP2j8h8oA4ncunKzIVcelpS0Ai5a6HyVtbkF
oqmYuNMYlgMF95+sVcFdBWRua9b89Caz+mSpaNbfvkdPKbKtlmPvT8sIW4Rk
w39+yPiWcV/R6+Sc5Rf9n364rK6AakvJt+gzaEEYoBf8Qm5O9gxSmgeX09tX
juA/6CJNseZ2/pvhXyQX07l87u5OdP/1WukuwxDFYlxHWw11LWVHRMEE0vuv
taIAehT6sFMD/6o9HTheIi/pK61R0oDLParC5et1AEh56NtaHKwkHQOtg9O/
TgWxKKg27LK0QcI6x1ikySzNShrtvGO+v53aZsjNeKA9MoQqQnF77uO3bdaH
VVTbvZ4fJQXDnbehfUT5en+EiKVpSgUcMh3ZXDhnHevhdt6+1pkjp4DjldAl
Zg1HgV7cXNcQeu5lDkqh+eQ1elGfpLVGIBtc8kDGnNxuZ/hqqGbKAdYB1c3y
xKEzAKawu4gUGZCp0no0fMlwhvGJav36ZrCBJThOGIVpbOko3h4ZaO12rVxH
NYAbesdNis8Lx5eLMc2BETesUU5R54Km6/L/EmW/Ne0xzmt0WDmA3LShjbfl
q15Lu1FQ5fBiNZW0aJRnowxOZvsn0PMO1naDmocCjmFTpsHCdq24cwX6qLhp
g1KBBm4zfEN0MorHzZFYMTijqEcrw7S6OCoFVzOpGXPmwGJAfr74nIfL5Jtx
UovcXUEXg/xBDNJdAu/tKnU+lln8QUEzFufwu78ZUP68YbCYWi36hCJTihQD
HnBMGq1X/SUNOwdr2+TKeQzHeEdhbsYH9W/YIrp0lg0k2yuSMOAZx0P7KVKs
Z+v/iUUxo5s2W8xInI4zESFigvNTdH1ZMpKPqZG+9Q2L1EQS7K+miQWgrWPT
1wazHVmZx0yGXRSfxy0V93uC/pQTjUJTNTD/SDzc4QhKeJ60zWd9LIqI0qOf
AupsL9BBzY9Ws4dR76+oRI02C272xlp8Fm4B8a6qK+j62nu2nO58TG8vNw7j
o2QFQFtJAbYqnrLbkBOfdPZN8HgY/oUHAic8kiQGX+M2w4JkP/8ttdITTdT5
0X3ZdkwleK//boxvPMXkscqXAkYe8Dk2osUrMNqtEjVJ/2S4nMg4GVBP3v4V
4EPJN9Vbx6KQtrLlTtGH6EkOAdz8stnGGblWmyNGOm0eb0nkKkjpLWe3+JFc
uj0+wvam8gwLwf2UEaJpYzEY7Su8TsQpzL3cvgm4JTYOiTUvoPRmoClpYjzz
GCJhYF6XgTPPU2aTXruKv+SRMVaVj2Rb7Aakg/cSkNggpvCrlmVYaffBTbUd
1SLDkKOv1WodwLkeAO3qRUPMVE0cLCwL6T2/g3hgx4WMoJg3plXcC0fWER8n
QIERbvY4T5EKfzzc2OY0AwUFpHzjRUw+vHH1g3rqW8s0EWckeMRD+m9qJiG+
x2rNM7JPmYglSBNIflXRoVot8Y3goB2U9/F33XpchEqgYFom4XLgRKms5EpK
lVsc//Xu3GcsxAoh4ohmG8DeI/W3YGmnG79aQOKoi2ciNO9DIGdfCr+mqBp4
XYGzX2S1qLT9R5dvR1p7i+1OmdbPAb4dczG1oSSwFsfkr9FHFpwgcnoUbTG8
IXSKgAn4mgkVwIxa0W+R1RGtLF7Jz2VRbARyIxZ28T2ZG1ijhxHFf7ngWI2s
GJi5qE3II+fRMizqCfhlTnSgV3kQtYiZCBO7dTvRj/sMDe7L2uYM423peDyA
tjAlFqHC+rn9OvDJi10fjTxoISmuttUXw1p4Ie95qmdpegPjx9Rie/2uJWpz
pfJBsig3f28FXvi6Jq9fqaG5I1+g4+ABY6wlPtlqGIhP2HulTHvY3pnfVn1C
VldD7ObYrWloSmQYcVVdA7Jyc+Ija+Dj2UYW0oClnVU7oOfSQkAUbCwSR80Q
z6CQqP2/viZuPPcMncO+AeDSIzSFzaAvYy78hwk5WHKLzqSSBVIXExx8VNYm
KaSbQRssYE+FPPTmDWfhyyePJIGTMxiQ3UULFig4ipQbCXwPL0SsCJsZl2Za
4cz9Is6o5luUOt0JF1hM/bzIAjlq5SiZNHAPvye4LBnIW018iEwTIcj+0oso
VKY7f+i1dggxc3cnDa5owKEon9LSxfVzoJ0XLGln3+0eqskdmfyN/B4Gs5u1
hgDHJDynh3qyuS3tUHRr6L2UarcU/knrWVamRgt0oLIEsn+Jd6mLh+VpEECd
CAHbocnYB5h/0Z90Q22TnqE92UpmulBLmjK3qYB5eHc1oUb9QqmdNOGkG7DK
mc321I6BwlMXIdJhqpD1RIT2APSkqMNuuTnvPx3s+T2lU+ADL1WnAZPJzkj9
BJNNzS5QIudl56gRBtlz/BBJMUVTUHcz19mQY17XzSlKYv6gYpcgSFWO3GbS
yqsc7xY/OREHRWjmm3hbc1vqDykfi1tT+TSaz1lLglglmjbjhGEtKKOSa6uj
BDzl5HBx3U5JQ1IX1jCMKVpAEZqCF32zne5KaM2yR85qPApBUy8kG7K7xlsp
d0xKER2/1TY6fKe8noK9mhvw/PgCu45UOMtgpj+JgVUYaeo2eGgICMPk28nN
CdElQd+lh0/HwIjoc6SlyHlR0nUqnZvTb/QzqXXUqPNm1MKvMGw4sDgY7iYY
QETwNrxo55luWbmS4iXHe0A+LbJZgihqD0t68B6AOfDUERWDbtkdx01A55w/
11FGqC+mbArC4l8vkqBSlvQz3PJm9Dn5c10uKkC32d5U5Rj30a4hSTceAh8M
d3qtvdjFUdSFPkZM+hf4IpcBuC92YlBl+dnIm5go0VL2tAst3k2HRwKxwWAw
lGb24UJ1RLXm+CY4AYt9wlHAiCsbZmOGEuabDwzqj6noLvsvnoc98X7kgMKn
wymuM1+WMbZ5baoTFzCqxs4R2diNx7PeGJA4uOekxRd1CaJ79OdEhEOBSiSG
mux6Wjjb8n4A6DZRhxbxDZDq2y+xIOYPMDGEs0CKg8AH4Ohn1KbIznnvlDRS
+W7rUqpr3n0J3Wh5zjFg/bjtZmCuhVdSFzfClQUpJhnvYrsBblXv9yetSQgo
s790qVLmCabFG0lkhC+V1d3b4iJrwYVuSx2LC7L28lrpCQIPLmhwbv5pWsgp
GWoZ5KnBnl+ujP/Q6MsVa5ywDTZVp/uCsT/ppfM0pCEXRTSWvVqYWQY9j9+W
POwCzxy1JWfaOY1PKQATFGSo6kMdXF7/pYYgmb+BAeYEb0TMFLJqz1rpZXVC
76t0W9eQSaeghJVIw8FLQsWm8frWZsUdjN8eqcFU82tTQPqCQalGLFkvr+bX
j/T7GjAnXl7xD0l6W9Wns98HOPqFSAs7a/TZz8Sb+s/BFm6vFl9JNCSzuWpE
d3MukKOoiRP95XkYHeSi4RMVjfbnkTHrTq1bkbRreLPjmfA0D/huRKDTYuCF
aCy/lNph21vJxVwjHPmXR5JmYUfTSj/DJoeJDBaGYeU0fbqmgTqaqCAw8eUo
PccqhVbPjtmM25gFjWidx4ah9HNuZu9bz6c05KV8laOC6vDctx4T1CdUQAwd
xhTHT9ClOgwLNLfq4Yi7vUkRy5/fvkrIQhKz9eN+8j3uNxavYanNtsRyvaEa
vUrDCdKfslXQzIkl/TFaBK3kTUehXcjjfS7ooqutfDUu+Nf91+OBEZaGLvlu
VclNyGEa7sBzJrgm9VF9MEvc1VT0zxLPIJ1Au+heOMSfB0/QyflXW8MYv6m7
gAUmFBRlTHop1FoAPvfLizHlfH3ImRUTtqpLaWY2nOUjsh8udvkM6P+rA6Yk
tpnV9vCnu+chSLb6FRfoLGxqRcUYKUDBQ2Yj5vEQoKvtTc6WbJ+2+PilqrDL
/Q/UWl9OfLt2A9Le9zemYmL0tpSOuvyXO9G+QR6dWVF+SlOAP6zsylY35eMl
HaV2ysz5pfN/8YA0HbjeQVl9lZskzmIgufQ0rbVF3DWKx3mem1cS1Hvx50fs
Q0yUCi+a7alYbJMn8jYeYBJ1jthbQfZi2T99RrFPu+VSk/KzlqHicfnvmm7i
ebOWxHtpgExqcRS6AA+lVawQIj+oVpBq8oVYJNzCgeaporbnnzJPCe3rsNaq
J/6PhV2sF2LtEGF3GEKLvnlS64E8z4ta3aQ9JmIN5vgih6t21nQfjragJxiA
0koTnpGJ+cxyETTDgSkQL0lyUNUduMAMi/68EBmLuELEAcK+bWzcSbWX/QrV
az2zWNj5ORXHwx/zETYNSnkH/GCB3SJZi2ZHFOtdHPqlSZK4LPHxT66R78mu
ph900n9B7HBR1vJX1w74JjOWpmsYqbqjV8QF80E/Gh4sqS1P9US++6vqOqrS
Kfc37qTeAd+k6F+tGkoV3paDEPfmrWVPS2a3da+3VY+bLE7T1Ok3BwNXLWD8
nZkGUoZY4V4LEO/GgFEuQAQggo4o3A7KeeFn8pSBEQbskZfaUjq5mSSpxncd
v05p0a0uue9r/L1pvh8YMQV9AZF2guVx6S8JvFviZLBBI11kmfFAYtvjDSDz
GKxJVQdVTP39SqwGyuLBDW+3glCQ9osXCDy32+GpQouoyiq7X7TeEV5xIuOh
LdweRAo86v0sP2F8ggwqqwOfHtr5BZH/wWNDo4BJKEWFHukzIav7ji63Pcwx
+EH0gI5raE+ELC+WeCSl9xseDyIwa7Q6rvAU7jt89/EMR09+EwB05Od71pQn
PlgnAt1oSF6yBqlSArhEGQECqwjOEsUPbD7WHoTnVvIr/nondyh7ybzmGUmw
3r3EGmif5LIejuAkRWEYcWr/WDDnM2ieFnEoDQRwXgGLKrk3p2h0JnMY7BEs
Q3xrA/G9f+DvmmGoHrZYiYjG9hpD0aMzVR5i1Q5QAGOgjt8Sbp+neSFV9TiC
eziH2DRf7WpOvral7AsJFTXyNdjxAh/qKhSzNB4yDVAZJFKqSTzq5EwLx9hk
WTHdrNDGz2a+yrlK4yuJHOqil8HQ2prBGPvJgnosZ6XFMHPw7ewBYhPzf6Xj
IEtiba6r4+WYgRi4BqJ1cx/45qjPjeajZHHX00xqzw6/rS7HpbY1J+azlmua
mBel6D5bZyAxl/ZccwsYZHQmzuv/4zNy7h0A3Q5jpQWCqx0bYwVdYwhUPVOH
q4BpuXsYOaGzVbQgNq9oLVKQpAWebsowWuJbr4k1NweznamYnLy8UVYVSmFQ
CC3wLw1XeaiLbsSfIv3cSyfK2x24qoWOq9jKDyHUpBdyGampSP32lkCxK0hv
P6WgP9DBe8D73eJfw4yGftHRagO4/OGeftcC5kkfytdo7DpnxA0F8tCp7Nze
3PWDsvf+Q5z1EBSfVSA3zFLqEcP86DNJ5A+WHzCyVd73ffKSqGNhZEANeksT
e3ao70vQFXxkInhE9RiEyI9BrVISSMs03qRP5mCR71AWS4LnEgRKr7j9yTiI
U+mgpD5wJIhCkoHrYMNPgOJ+nW5ZDLaVvcNI0np7QBaxYuIc6r3qfeZAc3MY
XmvtKClmk3dfwGuAHwW5YzJIw4UHEsVrDmem9m0c6WtPih6MXf9pBfZRy6+Z
FoRoSohWw5BfOnLTjYR/aEX92esYX0xDbl01VmA3U02IuWvq+55JwvDtaXNA
XRnwTxadbB7bPzNOt/+fST6Wbr/5Owy6AMkDCdRObP7soIXEUqveI6U53OYr
NfAPnrnBko4J0O3gsR5MwiHuo764HQJ5sondMgKOXm2K8oRIYhoyD4hlaNTT
yJr0AtFH8g5riSmDsplY1O1zwU2ogbo/jvS3gQBQv4Vwp3JF4AgKHF3mtR5X
MpcPKYtF1a8+IZtGLQQh1po6hq0iiiMSabuq13hr+vJ72ITtO2LNbKC8zUDV
bk+7aukCOJJIfedkNcA/ZzE6H5+1BAqGlu8Jkq635SaL10zxA5AgwtIIhwrj
aUfuTE2WcVIYPdy5FLDB29/ovzH9M4yRSji49Ocv0BH3NmmxyFwAx181a0SR
xXPAVutl4af4jazBRoaNZthxvsKjoNLf5m3TfoA/i81qGU16/r1w0jPtwOBP
9VIuevBVGPOqNMjRhonX+/n9Kz6ZdIoepjWtNWnnItBYTUDEAphSpZsA8pgX
MInQPs5x3pJ3rtk45G+yk1TL4xz9WhJAUdf7/+iC2oZg8n7YpbmTMganSAUK
susRaCHY+HI2vVp0FhGIPZ0UxzTlezoOQZj9+miFO3SV/gQAuzCfQOMNCCiJ
y99AQIBImniL8F+pfivAyUtN77zD4WXlPHk0U7L1ZD4Pdk8j1aVkUax0qsYu
iVveJ5Z0tbBmPGeWvS9teLDJRmJo7P1iSgCxj2ljd3Pe7fTr+tmM/s212klF
2Pn1yHMkD6q4TFqOnOq/bFTBXX0i9aXHRECN23UyXUin5rHbrUYubePmqa4Z
FXY9ZEAF3oHnlKKGDPXYSdTBexsYWfjqIipgSfSW7n7R6wmt+izPu5cDngdf
7TfADovmR+T7RAwkHHbHOv7yGKkWM9IUH9KYWpnQWXOalvtebKznksGJfrVa
E6ObJ6erxISO0BSNgdxpuqeXpbEPpZ+27EjZ1FAi9PiAnbkqjt2ZuAO4gD+D
eJ5xN2uv4sSdttSC8ITr1xkdUKp3WBJy0NT+k0Gt5QixJ9ySeZAivLpsQh9F
xnJs/OWEz+M6NOpVHZWdVtneqSc/lwxAMyoCMOJl4W4Ib3o5QHIedZK+TyW3
jmsPG0TYoLCPVVmZCMcipj8taj8eZcTQWS91/ZXjmG04Q243l/wbv/LuN9JM
AJQvooA+l9usNGEiKZ25RIdOgL66+DIm0Q6WM6g/+6dJl0Gykj6P6cfiPQ5Z
BbUmeObY2O6sb/br8r3+/ZnJK26yJ1V+IMv2pb2tVmnxodTX9iOCNYz2bosk
ag1EKzbNZdABuLzIzS9KqaUOjT3s47JaRp5aaCZTULF0jUNVtaFyptb6pvKw
cavm48Y6vVgmKHmoawiiDa/Kxmv+uWGypWJbfXp/PE/3YJJOzvTHohPeIdXU
14n1X1RI0CK1gviDimzNwoI7q9fQvllMeJu15PeYTyZ4kHjLgbHB8BReL51E
Bzjs349uE/XG7w8JV5vsBqz2ZKILXMxZLwxqxauwtFLm5HN35CZ358kkFHPb
1QXKORcg1eIC4GSXHY6Z9ttRTLG8LjCS87uKGdHZi8pTXScGUb3NpmROppRV
48c6FzwWyZyVBYPeRH2kqN+StnXXJH7gp9VeKWb70nikgwCamI/OPGkz3OSJ
F5+b05Hog8PEvBlJHBV8C3s8SUaS/3lbMzS381eFcG/g2YkM4zEPoseTUuik
TfEraGywp6wNQnyhTCjls6GKbpyjxJafjLtQMPpGE/2K2nJooxwLdv/WTLZL
PuHfXezl5aXjLKtrqyLZ45M5vg90MRVu/OPcmI6USyoBwGrDd07PTKdNlHSX
YGxNihNHVirRQPhY9C01c8KgU82y023A8A/qlCWZrHQxBtA/AcjyTbW2rC1K
WHsrImvkyKuPZt5n61J+RrD+fZLrJDtxxdvAAgvZJpBdl/BdRXSJskOlv76Y
i2Xagmi6vba1885tBStZlNhmYMZ0WsgoXEl36nehuT0RUaA+sQfiwVaOZMiz
b3K304kGt1qEHBW6ocQTPlU1m6qs6SRd346bwpYCrwzveYFvSNyZQLsvhgRa
KvlBx75S2ivaBoKbCvY+Nmnk2Ybe0syXR8/+XAgSMmlZYPbmevymYqTIgoW1
I3tNQORypcwgzefzsiTtuFvmA9YSpIYx/KTKxW4K3jcumMRcP7jcZfCJYMOQ
GZkEwEB86XBmZX0DHcsJKCvnJY6bH03SvYcFqvU9TAIM4lzM7Uzv3C2PDUM2
HwaMU83r8k9JSl9bFoWx2anEnzBxKNEDWG0EGw1rOGcrVgLXt/SqPpyeBVoJ
RtCnZaNFVk21F4n1pGTr665rRQ/5XY7fnmDT4nDNUj5mv+XlbVjcWjqMWIjh
/p/GQ7DWHyCTQL6/CKQ7yOBBmah8Fb2RAElQey0V6sq+4likMA7FpblkzCv/
5MhBSkfX3rgTLiz/ljc7C7ohFQUJgOoSlAt9Nxhk4c5STmFY2Tiin3OYeIfB
1587mM3UE8c48hkyMDb8ChSiowhO9Tz+wu3+2vgxvL5ttMkN4TpT6FIoF2cl
FH5l2klIiLwHwehQ6zxuLKZoAibJN9gCEJvfWuyxmyFKmKTRNFMVY+Ne95HV
lSe49ZQ3sABiynY5QgP3rSCgd1qgUL5gXZdlm7wZHLmhrj2DcoxsXNQKA2GR
ncBcfpJ3g9FlzYdGpyvPAudgJIhFG43jyrGChUWjqWs4grlCS41uKb6JXoUn
SKc6UpwmtF5C1FTaR34HqkUwwxqbdAId/RZlR71615oosGgrBS5JlEYg+usf
Fi3290t51fPTvrXsE2mdyP+V7Vm6roaNkEcoofLmMGr50ieJvRnu6x6bOn1k
tNByXLZr7xhGK3QQMV9pN+Ip1pUO4oeTKowqu5Y3IwL/0byz7DDTLDBNstpU
BntkoiDWAS++umVmiSb4R0LC9mmUPbOVf3PHP6oyZePRXEyfQytNLRT8wihu
Y8tsMMG+UnlskvW9Fd2yC4Ua8R4Z+BIesxck1BVgSx3/5yINlzSPAbYZk31q
vAdP+hdFVqv5pdH2XYFQixIh+TLncQdA+qbMmXepb6HuKM77q1KsaqivZudy
mteV3M1/6sWFIWf/QsUWFTGb9hM1ppMGf5v28uF5IkZc5QB1oiMZud3iP3ha
y7PWkOibdDQrHj6/ka1ayG/kdQSp35zRQAacAC1nQbL5HlW6cWYmPL0GmnxZ
nK35HsekuE8WGtyHwzUFGKeLsXl+IBKjVPifratHqyyK+XbvgK5ZxtbuiK5p
BivoBeUg3RNvDHSuUApDmr1bFRMUzT0ETsYnQvYUFLmD6AsQiyhGQ3x6yBgt
JXGhJ1lwlKi9a/EidD4V1S2B1P8Y5H9iCV6i6OZldNQxB4iedKAp/fQe4Mmj
NRcZfPHInf8KAY3Jx7vWSAIU91dxFM3UwfRIMae1ckuCxCaZ1noyiPZMSF3d
0NuvcXdkX5+hDTTJhDo8zxHMxwE5IF6Lz4sxTmhJs7kBMVqOU1BlldOGBO3d
mFTyBPX9GdI1qX8TIoP4vbYUa8oWGMQamBi+8Zf56M0W3O/tTbm+LRlo+EhQ
T+GsYhjR9dwMupeOyYwZZIxBioRNV1pxk0yCbwi4tYXiyQaPflx+7p9E3yCR
fXBZkeZoU5kjY5HyDoKqvTUPXz0EsXL3HF4MOyXnZmxxiydCCtWaRVYhsEyu
GqPAcvcKVX1wRFUQc6j19WdBBv81Z5sFVargC4A+qIGaNSmkslZkaCqEt39h
WUNDdhHjWd4E+kFiWMtJdUx1InFuulW2pMe1KJLKjj8syvumPXb+3Qvtr5k1
dTuqwLe8z+a1w5og88XXZABJK1mfewY4w04b60jonvJEd0na0YCbKF8MX7RD
ZcoRSwDYJi9AYt99bj4Pw3llgCOidhpf7NNHYyktrEotxEjC6IaJIMd7qAWm
NCQmrt5Y+6QslQYZ3PmwQGhnRFuz+BBMKegXzlqZg3F/7Hcc3x5OmQlVGWiV
9MezK4HaxzG1RHcH43fx6HSbwsQo7+3WoDoKUNdpFXSCyDDGaOQeIwb0hn0g
DDTJDmUQhMT+CYyEe4SoMf8Ioq7/IxJDnOwjYBMhTelhNGaEOhrUCm6HOlif
RzS5epkXzkIMZU4dYdkzgQwadFtcvmSKodp21MYij0a41lcY005DQnJcXawV
gDrOBKpSVSaUwABRgopDQWBNIoVnpLINSvRzOY1ehcHcYLQF2QB2yACz4I1s
fg3u6WzfmsxRrzDGgIjIp9XodL11kAPwnbLP18JW2/yLGqif1Q5I9KRe2TkS
mZfWZp/Onvm1cpGqIlVeZxw3ErPKJlrSbJjyAkB/9bCfyWaUtiRI5w7EqA2Z
RkanSELt2hQKLZefQVd5pugdLIUrxPwwA9UXKw5isUZbfP7G2fqk6gXqjjqH
W9AmvMdi+cOIotdZLuk1wvCGrIObzcWlhq1NARjtYYQi9DyT4zqjFYg+7/L0
Te3p3X+EGmnnYeWqx59+vnrdPCsh8onzJGGK6ttU06K7qMuhR2adXuLgZYV9
11tg8I/fI7RSdoQK02sCDIxyQIyb6VF/IaWYpzs8mkcSlRevDHldD3P2n68i
VfvwQAVDnmFUIUBBhTSY4k18WLSiqxaMJP5M1Fnsaiu71qLlrx8Ut5mZz+RY
R/Ke/IVrsWdNs49RMS0LT1uPX8ow+BEQFzxm9hBNJEUlzNv3b1c6AHb90Xe9
CR7YLP0dcSYFBSd0044cIjgHt9ITFcCMCOo+LhfIU9WY+kw0Wu98BMgCA86I
PAMYs3EUuqpDKtnZPeb0qdcOh1iI91BPHs7TWHm9PSE0IQuzq6A3Ie5JkClp
F26fyrdqjNAUVl80rR5zB5y5Ls3W8lNxINs7FRHMiZgcVz+7VqNbze8ebOaE
QeHv82sioOAFfusyEBifkU6yc66kUGBVcci281nRGFww6+7N9Ua88rdlA0Ss
rX5gtx71vRn5PB53xhUVVPtK0heqTOJEaPi5yKqSFGxqqVX3oxvbfsVqhfu8
2qs5Zvovlthjl+Jmj/SgyNJeJfH5B6XmoFsPZHHT7n0fW5cq8Ye57Sh/o6aU
xzqXy5Q4tpKhDzL1Q8XAD+JsXqgS8mPu/8NgDJMfI2+67qRBFNz2RCThh7wV
vveRxDUfisVyoARsX/pJEKLmlTl1SRPy6RZcrPxHrZPwdLFP6jI+hDIagbTU
pGVo0Pl3/ACgvYvu+EXh79NYvJ3LkvNlfNj1v/hNe3/1jYbPHc9EQCaVpxnx
OBYX32c5Z1KofFcRK4wInDsM82Uhy2P8oFjIJqrPSBEstBLc3y5BKhLrk8Zu
t7OKJ/5iW18rza9bd0k7SlMX8t20D1LPWucEwG9ue9koYoylumwsRSvxvQVg
oCbu/y/3qtyPj4ZyrhiFJEFDLSDqrvJJthGxfu0GBE0VbMMgDA9BxhI4hvzS
Y4seifpGRvXfwDa8JSQ6iiW43fsyAW3SCKkIbLnoUVpybGdFsxRfZl45wXMZ
0WbPa1yxBiJOxMIhuM4WrlE4LGN3iuc3/RjwlRfVI9ZVGjPf3+OkW4gJrjaU
m8Frd3RUUzopRAv/vl/k6JG7aOnuAEPox+1RkZHcEBp0TpXUMCByibpE5k/0
qT8RYyDi+yWg7KyulUHMek57bhUG9QUGqx718p7aV0fjEEaYDaQigqINJbuD
i9WhuMR2RfAWIBSvLniv93hwf68uD89b+kDKnAtRaTP/XSLw1JihSVJaTVvI
BqMepo9vTgXUZAUm0o++d0SGmx4nO6Pr2umnAGORYTdJe1Af555nQuhgdSw0
EUNTU1h3xs/fls+XJhYwqGXDUrLKf+EsVSz9YR/iHsbnbSSjVxRK2Prj2cPV
dfdOsx2fQm7MMUcmkMTYPJhcdWjhuJAKpYT/9OkU4ooJ2askWLgZkrMCIhZr
3ON4Jj2TohQP6fv5c3H9Qu+T6QtcDnHDEFXDmSUi/rRPIBelRGN1wiVaAPkp
jJrcKbUaKzA6dQYRlEWINrlMF+3UaDk3z1O5EAmosZ/ZvSsFRFC4uGov8jz/
K1HlBc2P0RgO/DLEus3c+JKfJ2C8H7fEV+bI8BBoHnovVSkre2STO832scBI
LBNKDRBTEV50I6nvJSMEkz2rsEbWseVYCSmP9CUrTNr4wrm0Djvy5xY6RW5n
xOnLMYcsGBBYszv8N7nE1kbuLz8Jh8D0bXKN/A/tkGpA8Sy6OdAhtsVR5F+1
SEeU7pCuOpPRtM6W0/vllt3OtXCvltScgKLBjrjmjDvhlEN5S/TU2t9B/Z0T
Q8oYIrMXQMfmqBjYMiwuK+qpinszKyT8Ty5vaYn6LkxzXLBrpn3ToV497UAo
Ent8ROa340/jpSEQMT3dN5v2jNeGPDSxa1l0TOLDDDXf/TTXNq5A6mR91BVH
icS46UdkM4eYrSHN/cCGoA/Y1LSDeRH7ZEQ/8a7VkW/Fup1q0iLjcBESA3Wg
Z7kWSiFRzqvto4mA75VscDmJLoE+KxjhUUIrUeMgJ6L2Bpi6lRbqJsmkuxsX
X6gwDHWQ+5MmxNkyAgXO4D+60y2tiw5WocXHLv/QLDUCgCC5Vtp/XFnc7ZDl
ppCjhF3DdujBAXBJbv/eixJf8p9CGXED5A1XWoEIdIb+ilZMsR9pVQLpmGWH
WmV9ftD2gV7j0MTejQD652upUUKgbRR+quRXL4DecwMnjhmGWsAdnkHIrP/9
CqI7eVmXeQKzyrcST/QJpWLUQ2iPCOb/rYBvD173N7+O3D9mbTO5+j6SzQfT
u2LDIt/INpTQOA9+0LxcKrbsE0+RJcywehOaPPg5kGYROl7+WnyvkSddgNga
qGWmIUnUB3lLI9XN2m5/Qz72v+smc2SbN8aLOwjINauxtVOcpKwLNFPZMXea
e50DtjkXEsY/2twhFfLImyKI2IBEQgheIwptrbFDUsdk1e05RlTpTeuffc+1
n+t72pZ2wFg6d8GODW0pM5jZG3XxP50w/8tASWBLM+la8ZaYFMs7FhXOMPSP
p9EvYdedUIiHhCuskaZrOeAkDQzw0SG6XGL9whqBepHxfpLMxFgRZqug2po1
DfPdjtIRupOlU4hFig14YnlkeQbL1iA1SEwh690BSBRnHB3Lfa5u4z1G7sEo
I5PeC3Cr00mBIiS/PmVBNAsFmjIpravDOB5y5v3UQlarFsOQ7ZfG2Ql+TMe6
/4cdMNciXefquPanG/VNXZZGTXNXJvV2IudahQJ3X999EirJwuLutOBTzFH3
QuLWJNIzWBgr665SoJLkmTfYLLfyWZlL3Ef7nsROh6Z5hjppLRBS7RnkJjqP
UEMUUCg2bzapZPZWI/csa4PN/araxzv/xCDb1rewChxx2qZ4+moqPAa/B3r9
sJXHGSAQm+APr+cAICoqsxjcxeegRPxipt8OUAhkckDngL3eDvw/myX+rFpA
+OHlWcR0uKbv6JOsvA93QM21awud3lE7ZE/6Sr8xRZfGJ58E13qVuaZUqZPn
nFPZojylaToYo849wZcOti6IWjjCgKvpwkbAn0UjbOly3geDIUXydXL2bVt5
m14NYcpvPvcZaqzhR0YHRojl+/bOJRzQ/ukhfa47eOiRs1MhqICUWN0dIyma
Za/3jhiSF3gmtlFDrT07Z328jg6G0uuvxa8WVyzTFiNCBrZBSCw+3W+a9e1G
J35V05tGfgM2KgubtP99mkEknkDvccf5H2VKwyj17jl8hfvKj/c659RfR536
wdj9XOk5uTQEsxk+jS+muB6nWm+G5P9d+Ip222iTSKZJhP1F6LoGaPxhAD4C
6MA9GaX8+Gp8+7aVsfVV2NKldOQgYcJ8DVIqFn5iDMLE+GbekbPjf3SIP0uL
/XbqFTjAA4YGjCm1CyGCJy0KlKfJ83R9iZKMLTci3ZYguearwYCX8jTc1BFy
rqg0OT+j6eipKr2KSevMH4hqzfrT1GKL1lz4cKoO6MI9fXExcYXh67ny3gLb
WFj95Hlga2uZ25ZK5cdnW38ziF6VaOLCfkicoUu1z22jd96EGH9YLafluDQ3
BKXvzn1wM9llAI+0zmXecjanZqD+Q9Bqz2BSEZsRAG6TgKG90qX97MiPYqDK
PYimOsG7ueLqoMaVnKtaRJDqCbSjlRwAQiqqGSfHYlIRwfNtTQuZ32XvoG0I
GVENWwFVDlv1mdbiZZ7ehMgxrXiQR+XgcLQ/LUJUqpJ//bwdRc3xOtuojGDR
EfmlEWU53PTLpemxUdBRVaVG7JN6gN5Bco7OxnI73pTpAeulai5FlmHCa5G0
Kv50FYfZNvql/6ObaLfn+HTSxuktWDxGsoRExlGfW5SfmEoNCkaDz0YIJm/0
vNnXJzH+0Rm7LuvHUapuUzP8bFpY7RAENjOuoyedMbMUwZn1Msq8OeYoozaJ
2ybihq6ROaw/viehSJIMu9KUvWe07G98plPUgHy7VRn9Re3fPvZYWyiJXhnH
Wev4TIGW/+suSRYSXreEJpTVwnye9OEBM1ejW+x7GGmfsZDIoK4lJ30Wvcgb
WSUZz1txzv2oXCk6yQTVFkfmrGkamnuGGILnM2UQbq5AdELsnMkYuH9kx+ZS
vLMcIlOz5C57V+3HtLet97y5oBnlglAgJo5NNigkhFuIxBfPpN3ZjPrmmoAK
CYuImLCcgxSyIyFOg5lqIPLgkKTcU7xUk/a1SzdoBDab7RJn4HWRsykCbZ/U
dZjYP4sSvwDp+FVrplImXqVBo3mS+T5TpLuntgZY02ZqNfBt9jSL0ORVmfBv
I5yTF8XHqEevFTGvGxfrY5LJBRRXPHdA/HbJJ7u8s0igSMe4dFVJX4iQ/B7F
PUIGRHWeLcq73dKErhgk5q1nQOwukIdscNcg8ewxkQjtsHF2rMvqK95mHbho
zx9uvFc9CpQemWwla69bGvYWOqR6if5mgPRjnB/oDUsT9UMVmKrY8pIxu4IJ
DDeDw3TpqwsqW9Fo4pUpbn9+Im03Gsiad6JQ8HPw8IUBamcQdJru+qXb4hhM
696G18b0BlUlsrpnkW/U/eE/F/CjijcvlXptRQ+DTCIM7u5/Azl6ZfJZTcDu
54BSec5RyAulclxGicXU8XdeuEESH9SvQmSLjh1Zbbm9Ue8lzCAqa7QVPaqx
q8aCUyXVkqMP2yj+Mj3q7gADU5ZEqXzA1FTy6frBoqIJvyPbB8OoR+ngCaCe
IdR8mjfvv5x2pyiWKah/LYWY1okmXQGVaGTjzoAo7VsNJja7P1Bcqyti9m7I
hHiK4UvXkaj14BV3SedNXBTvyINoYGI8fJ3zSWT6JqAJkeIl04ePlv6Azsy6
6gXKGfius5sorOvbRh6WoWavAX9ZYWcTakmIC+shqtOcnmesMXOOy7oaMBf0
aIawD1jKP7eS4s9VDhkjvaJWM0CnlVcZoPR/PULdxZKDxKz4hdS4P5dM1OPv
eCmE7n9Uo1QB6oVjhwc/3J6pOVTJExXst7YyhylJqFSMfmxd7QHXyAYdpoQJ
P3zSkHcb7rGKqkQ5/0+HDSd7yMJKBbKIfObRp7CyFR5kLOlcxx9aWfvNmnuQ
ZKb5qX6bUxcdxNtwo5SgD4/qlZKb1jnFGr9Pr+l09UyYPjGkMNEp8m8CntIM
+snT35R0pjbcMakaPlZkPFyjhbcMyyf/Q537rL4+07kZz1G3xr6rdFl9bwHg
RHLi3Xdx7rMX7T4BmQhQKbLa9QTxlC4nnIl8JtTHY++0d5dCrXjUYgqJTTWP
aDRmA08zjF1eqq+fK/2mqKy4WXEKO5uccQTcxV1Jk7Evc0LzkZwYBMEHbni3
1bLC5smtfRPS6V0doyXsxdsLE0EOmVqpJ7rFHiNdyfGg8dW602gDEcsDxOVP
qAw6M2sotdgvtGacGiEN/OEWclQCfAMYYkaakXa2C+82Y7n2gnBdSXXi3+Xp
6yAnkEd1CH8ZY0dgsDOck6GwLXA/xGRmpQtNGxctIwKxJX+TbhzSoE9iFBKr
1qnks4gMUfs6ue1Rt+MhEOsJH4Ey/tfeqSSBE3jbaYrjb31FBFgSGqwJXmo9
8A4I5UGa6pL+yslUoqnBpBDDvs3MG0X4s4fgoXsDfO6c+Rsk5VMFV39Y8wJ/
CJTT/l1VFzh+PKr8F3/poOAbAGD8AYBRyalew4C+UvAa/mGqcERQ99rhK6+a
DAb4KTECxohTHIfcycc6CmP5hf3BY195Io0tkN2HNn7RLIYv9rtmeR2V3hn6
RH8ibmx8i11DT6TJxAink5kdNcV1eHYLCUo1n/qFENrjcn/iu1EbR4GxfbXo
ScQnw4HLAM258EPkq4yQ87Xeh5tacPFVYR+cYaFuEURdUSvhC5b0AdlNuGSn
WZaOl/6GJwOnJ6Oc0e8iNDHmXfcMEMXW0QzpZ7B8XN7Gq7JW3RIoFLF11PUs
jn/cDxOT7LPpi4FLTi4N6EcknvWV/Wooz7gU+rw2W3JFxgCSY0+5pPrV5XqI
X3u8XQj57VaxIU5+GU6ZdQ4ghsdBeJoWZ7CZKE/hTgv0JALNZRERy2zVx2I3
7G9rDA3WachoN7rAvxVAQ5lVOTBq/PctkTUA7CC59Ek/oGJyS2IHSMr00fbz
1R0fi+WNWccokt7tLFb1wTI55gL/tIkOEmVlxNvVMT4OlT9AWF76youB8kqH
SnUNGW08/ZwYG2rvPr4jEFqHV9dBW2r27bxzdmzjSDoI99By5onOPEasBWms
k6DL0bz58xC+H8ztPfYw5nh5h1tfNCdc53QgOH1/QTpJyWacNuaBcJhRuSzG
k7PdwrEQrs5RU07YET2Wyg5JLtrQzEawOCJ2VKykjcYybB3Vn723G0Xu7TpE
r1fv+C5STapFS3FeQmmi+dCCO49w8uJnpCsZXccz61Dip+J7JA+35NyoR4py
+9u2qK7ufD4XQFtDDj3lgClSkXlreJ9TOwaCyq5WruuntYZYNHQh0o0SOPk/
SpXIvR5i4Yn7ATCyI0xu5EcH6x+5zhSTWXm1M0mKGVBLsUyFttq8qFo6CsMn
RnQKN6UW+LfWBZRHWoWDUrr5KZtJ2KWFIFc2bGMEkfY9xr/e72ymauatNjow
pZuKBUFcB97RK2WsrD2hPsxyEFKe8Md7S9VqOYXPQvWmuFREeT6vvvqMcM0p
X1CJs6xB7/u24mKmPeNXJRQ5f2DpV29UC6t8Q4OMU/57HjZwjqAFMtDMERMq
TWf6OmP2E4yzS/voBYstBmm3K1yh1rnXPqPHyTYIQi7FYfHCVIQ9d3pixy7I
SEMPpETOTY1OoUU9ggJMw0xnYYIGzrr6IBMqYQpOde4MKezNlg4q6LKiQ1F2
ghzLf+FT3ilmuNEt3QbBvb5ll5Su1u+1dA0pRIodMXaP5k9/8vYIdBS0Qbik
wublZgtUkXOaCCTq5HjbqnUJidFDy3uDtKqHZIwEFasa7WjOVsXMJMPdocsZ
TFrmo6nJxbd3w6d3+6dYKSfneKUhyd8OHIkOwF+THYVu9u/amP7SMRmQPa95
7weEzgQCMZDqdoZDGgu6xt0MEtgXj8XZ3Uzy4KlOVIcwUIrBMBiK3ghiRuNt
rBRvLxUsiwU34kKcq/xUyaqVayViscspmLNAfPG3Gki+NlmFVxFMeLmcuNTv
6u6hCWkWHhN4L9roSSRCxEI17cfksE/HAVXdX304YHFaGZGAcwZqYkQmTsCl
ppDezDczJ5JEQvB4LiDfTGhOa3YgV0IUNUw/iucAO5JSH7iEh2zqkNnJwtw+
pp/b8h+sGFrd7srh1/WMfpsbiaDOwLJwjmeZH+lt36T7k4wopld0bXoqika8
x8fEgSYs1OHegG/BtCAOMGGwNi9ROVkZZuZQzu33eVaKMgpxfWuB5BfHlI1C
8zgPOp9ZBVJMzpjBS4/TBlyOksNBquG0BTixV/xoj+Yz7qerpCDvmswXntZf
H+VPn6bu2eUZFruOk/DVYrrb6H9+BYvND1xlZIvNjQt9hJlqDlgX6giKBSWQ
lyCs3FgNlD/lF0fc1O8Uva+qeVRx1nifAzNTMKm7as/qXWwzSzrtwSsfU7fd
4wWzKjuKlfzkOQ9dDSxppgcMZiy8fAlutXLaJ21i4iyqj1ZWeBrgzSIRebG0
8d7R9v3JSOqpS+aPvqsk0d9GC+5CB9uTQIVG0+wTLzESBUbyFXlsE2YNftMy
jAW288kAsLSR4Hb4BtBFJkUCNFv5vHxCIp4eIuwLMLUE72FlaONg8Qg7Pj3u
5zFwWlWybeiTnmogmoGCp+pfokupf8vWupIJf7N5VFrdTTN3zO3Scc+U9QYz
AeceCVo4MZL58FwBNz9Zeye79RbO+5qh6TqApPbWc5nhnyaUsOc6u26pb9yh
PR8AncorxV2vOfBORKOJdf+3LsyWAkYikkh8OumYDhPAlVNP/b9P9Iwx4HzW
QlFEFvJSaJsXrMpixJgC1iE432Xrd2VPjIGtnwI4DqZ5hRlctGOnDDKJb8Gg
de8v2to8zbwjpm8MmaWQtOx99L9nAjonz+YM0u8tGnURG8Pz2D2m0aN0rWQ0
1z+fMcVdmFefO2c0JNZUY5c/IDzIGRrp+RmuFSIUJarn8IUU6VCs2f3BUIIV
/UqM2sKiRj5UmZt6iihuTg2nnTXbRxBGwRBU+vcwtSWVN7h64EEU0yUYmEVF
OxB4lwM/qzaMifXP3LGR5eqpjA4MyAXH2pKevPB0pUJPFt638dTCIKL6tC1F
KTVtyjHkXxz8SCh5Wr+ReYAPv2JCJe6ASnflsQ6+5cHZ0JWcDp8ZWP6cSsa4
hKl+Ps8u1CfIaRP/yga08TGTDKjzrVgVXVfqrejDK+A7mwt57Z0xoH7Ocgax
qThzTJA6SLuTclaR+mc3VL5FXyWIs2bPjoflbdXQM98Uwd5fgzmsbeT6KpDE
jHrHQy/kylb7uuvJwri/4mxe9oTZunmorZk3BGr913aDZLJZGq/o/6TYM8fq
6oh1NKMdTqbKx92lPbGt0NpZuUNNi2hn6wrII6nDBYv3y7TfMcc/fa92Vcuq
93ddBhS+Rpv6ZDzpjvxCgI84dHphxm7GQ39up34UHcJVUv9IbqY3+x4Etxws
LWLVfDHVapJ1ix1kAJXfIlJSUMqK0YZ7tKiUUKUbLy3N8EX4pdOnuBRUv8v7
Ks+dnP+gn3SSqElLlsObVkzP5f6FfZnxm5ZS8rl9r95pc/yyw+ixE++Y6QFk
XGJvjWcyiACA5YZFE95Iclt/GSOxMdPrG+9BszQ5nnxS9xOorRKCeh3Baf7q
iUvL2+eidLZtVv4yOPM2zJrt/bhZKZ7AZzspkfS6Cwl2XKjHjcmm4VwEZ745
5jIe6zR7aP/4jB5MJLa0N9h2ImemuktE6n+M784/aVse6JPyjyHUcLOJpLcW
CEP0RULYWBKsuwd8RS95HDo+s4fbbaL1yzSWR2mFBOj9EmDO2q++gxndodb3
bjRJGFVlom+vgthuek6JnAqBZGcqHXYLIq21F7gTTKFwR2NEm5pdKW/kWi3W
0+KR/DHEnJKRIJFepDQH5U6rNvRwnD5jM8EKa0NWeEbYGmnUXMR+GpdGgacv
vYHfvyVIfiv3PjElZq9989OdlD7QWXQ1DfXPA8Dw+Bo6CypWuqOfVi73Irav
rWOx4f8we0LJKn/9u2J5Jg4MTXejhOmdkOYseTqegcmYAxekphgZ/D/3m8ed
36sYPhxtWZ+6INCND8lWZMZIE+U2NHTJbAuqSDUtK+p5qNZfpKQeaA+EEyce
IB7BQy8tb817NLnuTbRlloUuiwdG9b5fxDbkhmQtnjDAKTsvX6/A0vKVWY/Z
51TWJem7aLZUjCH4molPW9q4V247cnu6ySTOtHEBs3B17/PGpIKtUJaMEBMk
Ea5TkFopmt81Ku43WpEtuibHspDnKRD3vq3VE+OIdJsFMJaNfKc7izc5t9mV
sUHGKh991t589yGQ/tpONmzVwpm28sZ/rXt2O+H+qlQLI4qT43M7nFgI3NG+
Lnf0h79aL9Z8Kk1BTZxLTppdR6EHWUzAMJTvwXBcNx1VZg1BAmR+iengBgOl
j3P3pz+Jj0pQCsm3sFrYs2mV/NZ6+QoP4qF2I90NdvKi0lSY7vspRgp+8t+/
1ifKwiVexzGS9bRWYuw5dD7eWO7cY+Z5tZ5rI1UO9QYdjH65TwaBMZ6PBsVg
H/s0nybWQlfmhc54/6c0y80+17e7KWpSfMYseWRkYPCjTf0EvRR5v/8fcVSX
pnlCvHIsBuZ2leh39PxlsvP0c/rpg/apPZ3OqHdU55UHncD7smBCPFRHXYXX
lfbXvzXHC6IRzhQ/MCplYAateU6u1eOwWMcdjqN90hDWh4nFUAIGfSvgKuuU
rFMMJNkaJ0V5NCYOG5NPKjsB8P3d3S2k95pTquHWqmwOAnXyuQFqj+Dqtj9K
wbbQ9Ukr1K6FdfAoGc0wzBaVFycMqvr04+Dhhrq7LMWIuzX6Uzo6JcFPfjTh
3jB1qcEv1Hwp16o9d3QNvFkif0yyKMBQTDIYBeW2OxdmAXmrF3wVWyO9nnFs
E553rpYqdKJ/rl67aKH6zhwnYF14B+6hz/x/fTrEGtunkbVJt1Jx8q11R2kU
Tn4dal1OoyPdS/AQ0EPgDLwqzLEneH21Tf19QstDnvA15htEsZIflOct5Fj3
mKu6xvBbGvsJx9jacH2rNuzqp59kgle+HCTchFeX762Dhqwx483DHHStw1lx
x/jJqXPe8nyl/ANG3kNseLXrg4dPdUxRr9IGkw6rrpfncAphClqLvkI4Kpkz
ZEtCR49f3VBCYmtlJvAeFs7K0UtfPUO4BBMtoo/U/X9c7MzpPe9gqElTzQJe
hZiTxK1fnbNT8KTFQS1a3lUpx5JOjBgJgPfLWIWoI6ctne9Wv7QyDHNvRzKH
QIR9aZTXSVHmNg8sO1ZUTaZsH+velVUFuKWTXsbTTiVs+yJ+JBoaUoBBbQ9Q
PwyangkgET5a1BASXzook1y2RTXNEl6+rqY6jmijUQsLd3qtWDMNdJTIDwoc
1CdKPcxAHTgui+yhCcGe0Cx3eEh8oE82/7PidjEtaCKHTuKoN9Al7BqN12sd
IvgCVPtEfIurVH2riEscAXDU8wrOTy6fb3BtyQNnvuve0K3w2OEJ6MZJS70J
JbVq5d7J/IDUhM9poQlh6MF5sPn/UphMh9xj+PRY1VJqLSOB2kylx7+4r191
HrUCcyjV2hF873iU4fDmh+pjhuQEEb0yfCWwlTe+zxmz3OEAThe1DXiJ4KER
lac2SzJ+HU3+RWjxosDctk4OOn+FQJRRT5vVq/vfU5v1DcooY34DbD1RtXAA
LXBExeNxDYu19b32OyRT1ObNmdDzyRJLA48Dm1QtMssYN3+lj/QqGD5Dmng7
1CrCApb0uATPOGqcegFY3zpEMUfIa/jX9DKl2Af07SrijX7KqqKyornVyEmO
Oq9VdukEZXiL/FOoJ/SV227fM1ZTQpq6YDnjHADHYPjbGobCP8mETB0CFABz
+pc74T/0qhzrKcbzJczIbwQwK99DoeQtxjGYuxY1N1xJY11Lg48S7yg2oYRK
n7sFvgB7JLKz3Fu2tSJJkswLeccHfnb7IZUSGpP8fK067VnJVwa3LeGDHxf+
1Lia6lMKXbDqFffZl0SX55NcPCXhKgFiFzn6APYeJWt38oB4sAfhJn/nhIxn
tvF/QEOX+SBbzmj7wm2D8c0A/UPW9SYLas4AwfLgmwmkeEdt33amSeHbfoee
/+l6fZFSRsDQLZ50nA2b06bG+3fkjZ+DAxNh7yJp201fUOD39RPEPiyg+qU8
HLG7Iak/Ks9KZnLFIKTCwz0ym3R7CeZzf/1jwOxsLGQGe827Cs71Da5GH/n3
BDZ4buQwjt6PZr4mnailBnKMXbGZ93gyHyOnUOEWpQMcbcH6Iym09rLsc+WT
/OFTRihltMkqWjvjB3/WpVnIJ6tql+GZ3lz0otJKhS4IWJCP6MI6mS+1MH3m
Jy60nXvZ8ezc70mcflgVllJWvWokvTxR0YgfZsESMiMFfWfTxKTCSfXhKWkb
Ky5g69Rbu1vfPlB/XT5mDXaa0dGSJZYZdCfvaRtH1qEvVEbB302cL9TAEMIl
o+imv878lbhNVc0wEjL/u4zXJ9WKCt16XT+Z/ZK/H8sdFr+oJCkuZjTiKwtR
UhATFJdEsB0YFtgkedYpBPJHdKO3ApRW2z27hzaqvVijeoGPVrZeVFWoQjJE
dVSQTFNxEeyz1Gl5Exs0nJG88LRKI4/sZ6btwM+DYW/Atk22Q1lrRmzSwjyv
Itqhju7CJWaC0p+UCtfBX6Ke/KroWSVSqtQw0tZHLgJTmtR2nobaiZ6WgZ2S
Q3SwES814PjSnt7sXYhvJZpsk7NoA3DlelFZvD+yUOrv5BxUecA23t/I3dTo
afwVVOWxYWSnPR88i358+PYZQo8/iW2NOCK3dpi+S/wuIO3r9YC4i/ub6Sgb
yVlYfhTZVTV2l9llQF7dNhfd9kpXyzKZqtHPvwvhyABu3MYadD09O+tpcYee
7beTbD+EDwosQOu6hgO8ByMIt52MDbUy0kjs+quG2tUV7B7Rl4H6mMaSFZgL
WH6YPGK1YEmG1GUSvN/jWEqvP3VdUCppUofINaInNUsb2DQ4+KsTJq7AMSZV
byF9TpEB9lzAABKaQ9AAuV6+sPVJkvglhjAZVbtqvqtnGw5lIAFkonR2vpOX
+7pMfqBIPKZch9Hqsx+1+tU5nPWA6TkYv3FxqYE7lpH5Epz4JNF/Rvw2hhk5
9C4Exl8xlzl2JFzcPozuwzXkq+cVUh+8yLwp5YXa9JtjhehcNOixxviyNrRk
xDjuModLgymBux9sataTpvtN6FoAaSgoMfYjKD46Y0gdJ9h4v4Kmrkb98JJB
wuEM91cl9zkZnxUzOnJaGkmarzivE+LDM+ulk9H+HOL1D9auLLgPpl9TaVQJ
dS5I9INiFBQyD585FhJJNi9286uBPEBzymfEuWZeQ1/w8ZEfPs2DYyDSxUlk
2JRpuds7NrIPL4qNmQ4rweZ4V5IztmS7fyasuz/OO5tZuiv2dRGhsNDGTo8F
6eUPPzzgWHwYJpRXqvcx3/wWvuklF1fw2s0ilkRLWTeSm/Z0uro5DVdXTOzi
xYmYeAKVkVlAN1zTgtb1RbgfBMpy+x/SPOZdxRQhk6EnuyU4C227WAUD+0M3
WCcaycfNJLjP/dHbl3jBE5teZWChBp0p3bP2nvyk85+6e04IQZSxsP2l//ux
2d9zGnad+pD2gxlL0FNI7D5lIv9wZWmn8PtOIhso54sB9HRwCoOSL+ZR2Fgl
UfTdDO+ZUh+ETtV4+E2R6rnmlmHCRvzBZdVMS6CqlZlVS+nNyIulsN416U3a
D6ud6ek78Q2NAtBtYUy4DjkjMdOi1gefEwPfFTzoGDHwi/5NOyFrY6xRrFr4
/4YFqVrZ5ZOKYLxSplPrgeoV6OJPEGjNgX6b1R3wA+5QFMpv6L/mAEXHfWLO
5AXuGVxSTOvCPBe0liGiNdqkLSzbpR6C2mLbf3oWeWnF6SyAiU+ZYO6LZWG1
9IILF/LOSYd7JpX1X/4Thq4GjlYEFShw5FM54mDDQL3YI4h2elfyTJG5VCsT
0/6jZt2eTq/gDn8D/OCPBGgE1GfMM07PzCQm8aUbPl/TA1tEv+ruFq5bpIwn
6yYCe58kMTPgfzL9kAuBUV9aXcX+Ru9XThHyAQ4vhIrM+p8qdIeNwWEznJtb
1zWprLdYGqmTHE/GxAIdgs0DmjS7OcdpEfC9+CBR5saqbqvSQ3Q1D1XU4q8A
/03SxXL6dQsyKHSqaSTeLXlZIqqvaEBeqILhLe8paZphp/VvGgR4zZVNxIDN
L+BaC6Vz5q4qwEzC7UJRId5OlgHxMU6kWx5lwU/Zi0JUUy9cIIjzZNmYAYl6
EhYnuCwUAqcY+tu18QLxvyHd2WR1bk5sJ/8kRnEtgK7YdB+EUudTsqq3gxhH
I7ZI7Bz2rtnwnOpjPQsBIKUekCzNio7dVWC8BdX6V2HLSY0hvity/qzv5WNn
npGdJH/C8rv1sK9V6g+h8y5HZOSuGzZqPCXmzwqLWBkRw8X5YzPXBf97FhtG
Lih9OTfjuxjNogL9hI6Wt8BOl04YeuP+XIuwgT4PDOTLxvwE+9KZnWEwxeyJ
UaXYwGEiT1+CfLNgYW0iP7Uo7xOZQw6jzyLy5LaiwGE6YfPRm1CTTT3tF06/
N7xz0We09XLfhhHwvDh4BRKREplWZftwmXSdhHvBqeje5V9OvksczGLGgYo0
QFcwLfzHW5m+rYql+IlkLjwUWyErV6u+X+19jG31eYlRK7jHUvPN7Mg/LjzB
HWtxZjdP9/A+psl7KWV5hRbgripftOelM4pnVaX5sxotDNy+Akdxu0/2vwWW
rz/PI06rCSZCdCL4BzwXwX6WxFnwkxvAH39LkMeecD4DxZbXB4sss7FAXRLc
c97IvPGWb0GDMCYy3GYT9o0gf57Mvd8Ihgf35Geq/kDZwUFOPVLAUeolAwBf
i1gBNFtxHo6V73GHfSgD1omwuULkMhjDIq/OpZPL7dimh7ckrfvdx9WPKsJj
6wTl8hW2mWOR9ahfi6ILFlzCH+1j6/cgZWXhFRZlv/xBI5QHlpcjicmZnNZA
feOFcScq2FdMXxOVlT9WUdoLRKWfh8o/Va8icp/TOA7lEc9ZlhUuRybWqJPP
B6XzLMRyVXNI8sK9/3I3Ua9n8oufe0fzn8sOmqAOJzOkbEwqLt2dro5zkYGS
FJOefTzFhzCXoEFV7H9qTNCb9o+56zmmNEc7ueZXNT9H0UMK5QSMkrNvF8hL
Fj/RX1UR1YF86WE0CVZoI4Pyi690JbCjlUYi4SKIM9SNzqzPctNfQHcdP2m1
jdzfY68flk4ZxprMU7ck450erFg4g/UA59/jLoZYE5Hm8XDKgWVmLUw8QvnJ
EkkOMBbt/TuSTDioRNFG6SlLL03rLrF9tNzbbzUsgbAAr4lDIRzNvryWL2Fu
w3VihORRE3eNCDAwCZOJLmpzBN/UaIWdmTdyJUeJPGyFA6ZGuHaFlSKAf6sB
ck0es0SBOoa/0wS3BIxr4Xmuk1xh3O64SGAv/IAOfzEAYYkacoSlr9PHOOLL
f9unFLZ0CDiG8N78rSRLwPfDv8p0umIZDKqvglWdpcuf9OggcTj7BYc0sG8F
sr5z5qZOH9t+oRCm5Kngp1R9ndtYRfArD6A3LQl7b0ZljLFI++quCt1UWBJl
9t5y6j8k4Rnz7QD3MNG0vXcquvnP1we6ZQXAMgKsMcv5f6iiqh8LGXy8zYip
oV0HhZsWnUq5qp3nCz+1hRnRDEb0d+ItUCIeX7QrC+lW660Z71TdYtPpOQed
JI1DfQ2Szwrr+2iLqtJ5j8LlSx/uBgDyEJlYVN9av+RNUzpwrhL8foYAFx00
MV6oI1Aib8cEewnwndI7A875DeCKRQlUXwZsIxVlfsSJfAjtXGL3Gc2vZxnQ
ydg3GgOtE7XPWz+CHPfCvJEuuyTt61iMCmfAIfBoFzcv9zw7YPLpPXyzGp+z
Pgjpd/+9RcMq/1vLKdGdfxEkwXamw5lVeOtYKTgWGiPlzeF9i10wboaH+4+H
FhJ3zGw8zkyLlOUmXk2tZs6GnTfyHMONf80YgkBnbAFOeyMpSfEG4jGsjHC2
oNl4hHKnsbdTMPWEsr7H5lJWkiiKO/XIDH2HFc3FkvIL8fztw4C3WlhhiwgB
Xix3KGzWuMAvhgaawVGE9kLqm2spytoZPWRkpS5/8iJZsnF3dt9Bjf8AiHdX
Qdp/uhEsRNHysbbZv+6ztRII/8dbdYy0HE4oVKhOwW9E6PLOK9+ZB+X5b8HO
5oaQr2NYkctdfPJ1hP4olLE9uXKO8YFBQD8wUoVI8VU9WtxyRzG2LI0QXLwH
1V24XwcEr0+crefNndfQCh3bm0oMlUBQymfRYPYhato/NyzyxZEoWyFQXO7X
JpgDCZSgLQ7A+QIY2dpL3EeXwluGW6hJrWZcn3Sn8w1V5YmtLSKCqsAdlIZb
Li7eTa//TVZ1Gn0GLftdCIWMy40BopLMkU5XFvDK0ujVAmBbQ4o/fnR3YAey
QvODBM9rWALnwHVxFtVaE8f5LNwKPvi+gTDc9N8j0/xmRWBn/NEYluQmTYvK
SytYajf1S935JNOolEwsoBcnoDeMNOPeSbw0iecUdpSS/xQJRxTAsKNyOX4j
eNFwny+sYJWhYYyOtGEZ1uANO59P9MhO4R+wHn+0dzc8FGxcMlw3CEQ3izX3
tlTkulWDfO4lOPRbJLlEYXiZayfB0zQkDovT2I1jPYmgrtXzOZE7uFLMDrgb
uDDNQ5X5/DJSwOedxES+5PwP+eqxdn1pzVWufpOsiDvl1bxHjTqItcWyn3Ay
MRjXEaylxgPWseGnUklnemNgy73LAOxh//tvbVX5VgrdXsWKS8GxHMy2JZu0
oFWSWXfroYkiKUU66R0A4JdXp+fe18onAMhV8RFzFXoetjOZvphY0azmZepI
EMPPf0kgfgRvt2/8b4KWekGydjjFtLsOe+CQMooGXJCiPU8TCP5OwQJXMbYd
Iw9vkB8Z9bgQlnnGn2qHYGvytgMXWxSi7BOr452zxw5JlwWwqzuTgk+Sso83
IrGkcQmaq6RVijVnSTQVdQ22zuATTqR3Pl6zGOSnuTJFpUrJ5j3ibWGNfAyj
f07F7wl96eeJwTp80jtd93D1llekHlc+M9mu5f2GLTnuZL7YQm4AFbV0fBdo
YbBUr/Vixc1bhxN/PhWS9WkMvmtpCYFkQV3pM1G+dols8enMVaSeqqjb73O6
tmEV9V09jAnjN+Yhe+b5DH6s0PCXDbrSBPmqU4Pz9qLiKRSXrLLVbuknnJCz
1BqhRBBrZR0EWZaeVJV0zpLthwsTqe8aFygHhHC7mGf49mR+kz9b8USjG69c
YFaQPq6mwm+JzXBa1pzFWDnZ4UhELivFA5PnH3d0/4bvp0O2y47KNN9RhPdz
LkAPx+pnvIb5UFeootkKYoHCnyV30Ty3m8UFEpDFruS+u4ODEDUrF2SPbyPN
0X6ic6iYLExSj0vn2hveyLaTgm/WsxYRSYUIwTWaGcmlYY4d2f0vL8XHN547
brBIvGzg8EMfmf+xnhKS7fFDpOAAVv28JhFIyWpkURm6riuV3BNE7hAbQDCY
cKJMYmQm0O3xGnG/q7/HG54KsSvw+1r9uABQkADNkBRJ68xIhlsVZ2HYgTZj
1yz/V1fo27IUPqtdpCoPYkuJrHhvojo7gh54nA+Zxg8Hdixsdl9FH+yPV61E
VsPzAg4k1nw5wSR2ZXzB+Kyo+EoLUTRm7CzM/PosurAcUvchzF8fkApLyMnv
LXvbvDDHyjXpo/BX/dTNPIqaXMeHtg9WrY2tvEEO364/E3NIWsDnlRfrbpmd
3FAGDDwbSLKuhd8PQxjMVx0140X/ZmqjZh8slEitkK64yY5oHKQAu2yTHDmM
7zYLHpJeCDjeZjL1wKhfLDiGcB3cPpquEJl00fUUrruS8VDD9viXPVvXM/OX
6YVNSaeMKKAqEaFJyKjUrm3W/AFuL1jeiKjsDjDoncRBS7ZmTyKzPhzWjEoV
I2SxyXnqHBiasxRLCZEjiVMrpHAuh5uNniUQxw3+OeEZlEH37leRpLhDDySv
KI0Jc+NINBAB5Y3ormDSh6666nkUJTNdUSznJ/Qxa7lWiEN/QaBzk2s0/gqp
NwodMP2K0N3LMRMJ16z+4fzUDL8IqRjpzFjNAlDXmfs6lEHwrXJ2grcwyFYn
5yGgLnbCncGSeuj0VJhidleAo1yyzG751pFhMA/sJxrP9nC5vLbTUvgskjv4
xSzUFg2j+Tm+qxBb12Avu66+8k38z2iQ94W/oAFvDL9GvsU9IHSqmGHwXXF0
P0e8hgxHOG2pgJivwW+/tgMs7EUpU1WWtAwbG5fLfkjpgakk3o+PnxULFG9C
BZkTycTdz25XQz3BEhjwkpkw1PRlEqKffUiWjWTwyg0cGjR3RJj31jafXD1O
k3Ap8BPqllm66ofe1UGEEyyiDRSSgq03EJnPrBHxFwKLvzmZkdUp/CpiT3RE
rne2ARyPSzZ8SNCeZJEPjXBYER6Z7FDlTgseRK/NYDoY6fcs3ZPv7BHfVJJW
nP5p3UzDrbZGYu4b79iovnUfp7meP6UUkDBGCdh8ssMcwmhd+XQfgmj9hsfB
YjZd+iSOdygV2UCC0iUGWA9hbE0SNJo1jPMKUu5XVlgsoh8f3YzJdROrrUrm
ZnyPdCg1Qh4SMbAQ9s172Xth0KMS8NW0om+zr6mZE1cil3m5zkLMQ2EnZRhO
XXsdz0cGz1AfxGDu9T4pRMT9+MI89Q9rC17V4JrtW6Beluvrt1A5RNpj7jZ7
tnKYplvMTnEIpYqZVXBwrdMxTroMAIvSeYNgVxS0ENkA1LT5dLdASSd2W5qM
njwefaXXOV1Nwt1FCd4XOHHiXEB8DZ4c2WS3hl+EGe7N7Pi5q46ToRucpZm+
xhCUvUezdNVhX+DQOEq1FpWYAKWGRxqyvSO+IqpGfaKcA1BonaWTCkiwguEb
W9CYyxso2Albyug3LG3VDUUAZFUSBmWgtYslzEPoze619vjYceyRCI5d2ug+
h7PbLFWfOGSF3crL8k270uMXt9a7OIpjWssfaZtzQtvKSUSdzCsYIsxNLmcH
YFZwiwkc5UOZWf72ramg5GX7eJ0ADuadq/WW+bqISuficyaGRZZrokjXKwL2
TFkzi/tydAZ1GgbCbm2jBXT9JpVu412+QD50M87PSCgEoRDBzOGuvzWUUlLB
tSBD+SEYGqAJE/tSWXnO9mK+lWrOEna+IhLXKv2l6deRa4+nqknwnnCzJuR4
8ndZ5bWr0cNu21Masx9Bdr+CLzGjbt3yPzjwkwWZMw0zsdXNrRrdvYZDajEE
wgdtcBJcj5RmwElz9VOkscLIZBHd/AlczN5A6NOrIAMudyABhdDySGTscGmu
3vhc5rN7UcJIAb6sRmMQpdSKzzPk1Eti+s6YDFtKI7EwxutIh75PMsozy09d
hkG4GwSGlVYzTebsr86uIWUBNKRhYfKH8SYPp7DN+Ccp51kvDB8YSIbCoEDl
/bZfxcdg4zpf3r/FpS8zaqSUuktCV+Do68MoU+zCu4tuSrCojJqFikJu77Ub
3BsGqc1esVe8/ZSXyfe3zirOvw7SE+Uhh2GvuFFSfgdfDXRgRYO/AF6TFxFc
GrHuuhKYg7G0vA0jX+R1oqM6Gp3GyrKQCcQ8TKW29Njvd2k2vYU8j3EQqR5W
xlf+X1Os5uT8lAHeTxkueCvwzECHpl95i8VCCYJV0YLPJfXF90NTAjxxmQ9F
z+/VYaMPlhihZd+jZBogKXXAd5mcAD185OKg282qgxfxKVYxDBVtHdCbi3En
igDpgGy9KFtI0wAdaXq/RDnYSRHF/XaqQoIn6wX/PqQGuraRWZNTflHd1gf4
NQz/gUIRBZ5quaF3zsqNxQPL8WVCofGQAz/9jyNmrMau6sSOs9DdQixxvetg
NV094lRlhrh9XXrcOh0BG9n1saumrGsMB4sSGESIKphdTZz6d2UezrTv+x0Y
GfzVUqJJhcddWlHcLDXPcZAkXmt1Xgzoui8sZWln9UaUIv/BZPRYGit409Wf
C2lc/XSnLSVusIbLFrA09op91hAC/0T7lU22vvFvJIpe4DRK5Ntd93nSYGXg
wTY6UCS2xoyVyoPuHm0R3/tirNEqqBl4cx5qjlfFyYfn0lMTzqtR8Gd7RTX6
igvpHvF7LQFNxxJA6LBEf1J957fy1skTRpGtijjk0ywrxe+1oh5bIhc7gUNP
EByG126y0D9LYAu6lBiaUMlbQanYTytX4rcqHD63/i0cVeWlcI1wfzUeEMPO
CuiRQIj7kW0pSV2Hkp69XFQJJ55hF1u+ro0FnQQFpjWZ1YLbBT12q8y+MwVL
V3m4SMWuR7nerYLsga9+TmYR9iKmPJPeYUV+eHWA8KwS8GWzK8p5cw1/Ep3P
Q2s0CKh+V15pBSMP3Blqosg3bbwOR+NCDU8OxYkbGrDAElcJLBSE+tSUyY5a
0lowplv7rQf+sMYYnd0dgrL96jkz8Gq/ESPrfD+j9qntQyMzLUZwQpY3OX3k
XYJZswhnB7KOIZ0U3OQgRULDdjFp4yzsoXAfEp910zPKpR85A0pNPbrfLoAG
3MKuykREcb74sjYkYn2oQZqvJovAvuAKCelVhvWIXqTVaM0DBxnKOsZXYxFm
K+Dc9rIW7u8JEVvUX+9DeXCmdv+s4Dh4NU46UWZtVK7c7ZZTUuSi8Aht1yjT
EQfGoRduhAtsJe4RHOgw2pcm/c0u9QM1mw+zXOm1MoUjG/U3jpqhTKyzymRj
rvgo61hEvt8wZ4kLbxOGMvAX6mWT/c30qECLTY0tEOhls+PQg4ISGZsvA8ja
rBkshhrdhgYlXW5WUmKNAoPUL2ms/O9TyCgPMWbv2RcX/LcJCGYmU6YkMhFP
yo2DeHSalyEBiilcLADlHXP0lzoSso5pqBxqLrhg6/hO9xaWxZ1vwhoIcqqw
MM/eE+lpawm3YMdL+qRnp099I70qLCNRPyQ926WkjQvbPzMcsMidwo9yAUl5
lAN1fdEHy0mCrIerteanHLT4QUSzuwSXGcwtQ25eRNBIxrkkP9JZIDUtaaJ6
Wv7kHIdFaOeXkclChpHWotu72B0PErBGO9Yv7S66AkWTXVCwvoiFge0Zeftw
O4QMugSkSbBNe9IHMnmSFVrSejpQzgZEByW8UgVlbSfWloFKq3ot7fl+YjyC
v6UVDK1EEeyBuSDCKgXOrbdxD/VCWCjCykK8OhE3Su+xbc/wLQJbQeVXwAit
H+zzpI0tHTmmjdSe0AeK7BOwfxHpIDbxn6x0MPk0+/EuVVowlH8/bo5TNimu
AhRJ1AYSZD0/dal443yeVaFtCABVMiNBxouGhdFX0kUmLJvzi/jAYKm/E8e4
isJXPNh2iuFbs741xzLY5vYjAQnLzdaY5DFp9bShNROjWCYtHdgpdMpY5KQZ
PPsnYbzyHuut2HscCkbce4Geo5OVwUMHRLLE09jIXy02AweWJhgRHASf4SPo
V0ql7Bp1fmk8E1TFlOKM8j+dEtpKqjsGDowjdoJHFuqB+HmfUY4nQ+fij0SN
xfaRS4Nfyf1iwMDYI1hZqWfP6tkyFF9/b6rfhobBT8VwDG4t2OtKcNdr4XvQ
dCZGrwzmL2ZORE4wZbq9dby3+tYaZeQtxQN24Om5PbQT7sLosdhxolzcXNMf
PRpjnpZ2uWsQv72G/xDVJUrzUC0ThutUPJZZmHFPGdbsumu5fKXPCRkvwH90
mRpCcIXFT9aLCX1tHTlkvYH3Kzx0b4nSyrvsBBUp8NfwTRG4TKtlkVAb8nTV
jcIzvBTLA+HGjENlJXYo0PSUMBJo2V2mAYzTjvav9XcieRbque7ANpIgi225
m/e3XhpKZljqd422Z+y/gRp9/L0aNKii2bGKnNjFtWwBXTiyjGjQqPXveY6A
QjXhjHZXDbEy11arH9MpEbf5u99gOAF52CwS61g/zEtWrobm9xPGJVQvjhXO
kKo/KGEwDsnCLBzcyIe0gS2kjjItt6biUmHyidlvYAMpf3qSfkDd43YJ6qbA
c5kQdzj6RWIyvtxltHPYxHrTBI+WBPBnQQ72RBjl7wbt/z3V7GSgndYoDdcb
jHDSZkA+HUCMgG9m//lgVhuhCnjbxpTTAMdA+jGKCzW8hEyD+VjhSBup1N+w
6VPE//Ynj3ms+xr2G/Jo3chOEv37vrKcFuUis1/gHTrOCcjefYhVfCvjHoFP
JNto3gUQjTbokDM0q5//KrhrOyM7hmlWymi09SWhKymX4bm2IgSEiC3M+ZPF
VX/nnkBxmCF2mcAGiiNod8Rcpm/+NWCklVu18g/PEnPcbE5OuSkFqdwaVTvK
Pdz743yPnNONDlNcVFbA7YTCdPooDoFb39+ajT1v4IjHuC8G+zhOD0oAjz3+
9pikaMMjHQJaw7UZ+gj9i2XDcq6KGZuW+wcflz/xswCk/6mGyqbe3dq9emw5
J/gweZ4sFB5U9wYP5F5kR8t/+7jX/lIPlDGlG7bHehtmpp9RBkYvYcOY6b7q
LoU02OPtA/6RP6cuucyUccX2v/tMx/+oYMNzWLG0BS5aWn9mKhd4vnZTJCWR
nfofeOnmqoKszHj2yKo7XkhO4RSaVjFc81ZIihEi+LGKCUG62+jCqm6eflsj
W+QuKcC+5lKzdec/YnOVixIl56xuxcnit7sX+nUJF0jTfXxypM98ExLJkv1E
/v2BkZcqLhWBrIvb3atsqlstMabPYOrHW19yNHvyKg5VHfj8jHVXX4ctSSl7
KEG/1iGZkMozj+hj5DFlYlx2Rt05oac2c5sMWN7zgTM7NKAVq2ilkCcxQmy5
H67W2DE+52etBMPQpllGX8gwhvKlxJ75b1RCNpwzf0PuGEe6n27zP20zuCpT
1sHEHvkoyux1fUUOi1QOTC0He+t0D/OKNJVV9Fiie1cSCK3ncqsJSZcGDE4Z
Ed8RXVYIT5xCElR2BWS7tYM3dbBf5tYXFpyZBN9gQe2dywiwbLEec5KTO3IW
2lJkmHGmac1r92nfdKJZ6hzvnBPazXbOf1/e1bMsZsG+qQ8pT2llvbOjJP0P
nwIYbXg0c4758w7CPXjSPom33W8pPF0ebbF+RQOqfmbTOWmknceDkiT134E2
5cMX0PF4227ovXXE0dpCI/pBP6jMQcbpifYPw124sGVYSICO74nYQxE5io2d
XbXNQelI9aVBkonsniYqLXxNvZyYWwTjpkG/EMIU1l+ytdie3SqWf+tGvWNq
Q4EoYyDLPBoVp1g9u38Yxi9Kfu0O43eUCFwxx67DeVuhIRQuYcOX+qosusBz
xN4ZH2dDnY2/acxhIg71g8DBWVjvnzltCEc5XuiQepj39tphqIYzYUfF9MHQ
/o5CvbhL6Uq4F6mxWtPD7Fw9d2V42GRQWqNA99W3nOVk95f2qqJV4OmUArmm
R7rR9bPyg28fiG1FuTSeuFIlobADwItIOJ7K4ZC7XNp/57X/GM+FuiOYPSXZ
s72P9hqwpEIBRYRINejNVNz/jlwa4+nWP8Q+BU5U/5LxEX9rbS3mWNP12EnV
3dy0sWWCksEKH5fRlNok/11hubwIJ4L3lWuiiIlH2HzdkD8x1Cy6EOROzrS7
xZAW5yIUOJWkRShURTLdnXXwZ+2PW7GkFh46twsaH+a+F22XJETb2PnvjLB/
uLOcXo70LS5euahstXH9/Hfg/1W1GjiZcQa/10LWcJuryLKkJVJ3xR2S8WH9
xNPqOCrZT1F69OwjceW1cBmXGa4Nal1QWo1XtrxRlGvKTdJTcokCgNnMwFyt
en2E2y0TLxEzoQFptD1NUGp1L5XYiKqb5GyUjXW5m0nqhShNjSd9gjX3OGfV
qlX1KcDreHtHc4Fp9imCgSYs7uK1Xl8VwKPhajUGs0fONRgDn+PB1EHmLSeH
Gblycz0EeEdlJWCIFixtAgmizIlWYS+CUsM8J9WiHRWQ3/GfZxywxccqWEmi
rxmDznjoIeMRa2WciEQb47iOtS8nogHDfLvQzinU3j76RIGPiNSy29mBCij0
ANlxLZTtH32OPe06gXh6ydWlN4GkTzyEm/Z7YThEdLY9a9AYynCzXrIz9aCM
5z3gVsmYhsDQqvamdjBZNbKADxjlhKD/wvzLkVHfFr47xX/0ChHPUk8EJLl6
oHwNB0J0YxK/X3XABDDdo67qH5lPeaUzPY3DxAV0YcaSRra0VhcE7FTZOIP0
JkO6DumaWKqzZe69k3On3Pk/Y3/7/e77g4Lkq+bNbI+21t4Nc96tNpnFg99m
U0oNFhSJsK8z7c2awGpDhoXJug5rZFPntZ58YSZTVPiLzP/0MWFCb+6qmjt3
rIwAhBAIRlhxpvJ4ScJWYF//dxmM1mf2PTAXEedXq8NTsExxtKK7G5ylcP6i
9+vBV+T7yvTekUIAZBIHiHO3jIs+S/J/aM8D4IDOypQYxlewAp5rkvEovLy2
inDh3Js9U843YhfxpQFvlFHe2s4aN3COAYZ9ZrI+ajlx+UW0qeSQXpQIIjdP
lbcyiKuS4aGp5053FSwR1+Rehg05dFMsqbAc7WlqndgBeU89HsoTAcdlskJB
9ULNnhie6/caOpQgDFwJtn5YP4ag/MyDM77Fwcp7mUjoXonh+Io1pLCJGhyT
J/ZjWrjq8iKqIXj5KF8DCbKHZJJfeQgdu/v+oZIjQUUWla/Fb5MBOBGUqXqP
51c4Kx1D6LgAkPhCnAJDWwbugykM3J0Z60ljFzfGR19P7efqTGD76Q8IwgEI
WFkieDeihGmqPJT+MzcgAcWz5c521JYAZPINDntT4MLqsvo/PMONjxBUQkPF
7NUdoewJDDTiltSsbJRQG/QLzwOlO3K66uqICGM4mrbav5FGOZWxsHuSP4tn
trAc3mBgJdlLx22eipbwsI9bFmdueRnBXOw73qka8Mf5NsHbPJhmkJoouSbQ
z1BRAcD6aftfcuPCnGRi4QxrYpz6xD46/kxkTtzNJbG6tasuD3Nh3iWq8i5n
6qkQK+8r7iZUZqT7HiA8zRVHy/aIN9C7fj2IBYBM7bRkEHCvSi2sqeL/nKlS
j1C5VpkzoqYQqhNonDmWDVQ7Qr3f8QuLZ0EWquNUuT8iRBnTD0DYAs0Qd1ux
mQqRC26w+HiAC1dMkCoOHp0cS8ipa7OZxS5LAy42vET0E8SV7tTsXAR6JwON
qcfjH76aE1glSd4FxToMz4BZW1dnn+lUyl+jw/IbBlJaadd8oCzyy8gJUVpH
Rpy4Nh7ZZex6wq6frkwJiwSkXuxFq3nH77jtQzsCN0p9+yo3PPn3t99+o03a
uZkr3mdQPr92gIcK2kIivvuMqrZZTywztDM6xfzy4J0KBL+Q2aVHggxd+DKb
XO8GIS8ngEgrQyklPhjnLdmhnWsQ4ieKRRcLRPBHManegIb7/XA+dlZn4jH6
sTN13dPfY1KSVc415kPty/iuFyn1f9WjghmK2f2clKI3LXVkxbR4623gweSc
Rxd5ZksduWG7DZGSLOO5GHuYLa/GQvMAw5ynOFLeTAGXQcoJpLmt6RNai+Cz
YDp4dJ17JtFFkmEiyxBcH2679brDzIXugnHsv8k+RjjI7AVF7gFeFMo7pp8y
n0XeAGYkt5Je7aXVTwUVxfA0Hm5Sznd7QzNy66Lfe215vPzJr9mtTCg1Gv8H
A5dQVj9lTL9jv1PjWr/tdPuw/RC4Pk1UmxfWScjEKxgamH2cBG7QVQJfwzHE
FAmoIasBIvHD9OTyg62luf0B8I7+i/Kpy2JdJa8Ewde0kt3DxAtX/KA3sqrv
+XWEDbFeklUcV8d+1eLmZ686MlcCb4WtMb9M6g7pWrvAHlOMJvE95GYX6HAv
BnI7udLrnMmM31J/hOPmNInvE4YP9oX8PjhiDP6ZclRj8+W57fEot+btH13X
Rw/ocw95G4/OfxGy15hNVJM8usKOnTYh3QtcITTPdoA2HSjgfMdVwF2rg07T
KwG3fzw2Rwdw4I3CrIbE0uy3pf+n1xJ2mrZZCq/9ffYnWepzcpxs258mHOJu
Be/I9VwKEjp2Kug9rhLPtZ1VgHNCLD8pny8nHcbCV95JZ3hH80x5iuJhEjlY
mPvUK0zXtz4PUXCKfkEyTyvBmbLq0VNrJt2Xc18qDqfX2Qpr4yftCwqymknf
eJpEc2Tc1Oquul4rfj51HWtEC/ykPWo79/wgovphG8meS4hmIp1Co7875Gzo
tvosLzNZLXbdd8IrbcEz3rgoVc2UlvDBTiCcOgzUyNLsEfpcbQLksA4KaVS1
WUwkOlb/XJmMuXH1NOyHqm09yHJllxWJLlDYSgk7nBDkocjBz0Ma8gmB3HbU
GQJGTSLr+ilvrjoSeKpSE/HwWUpSZ0pcPPqxGaMoC0/vKuNWRTvRbey5IGcy
NWHZT5wRBYbTSMMWmr6HKwjpkxilEOMyVgfs3Aw7+91D3Kp+g3OYJQ7rboS5
KTKY5xOz/Kgsk3slMNlgJs708LQrP35sjM0RFrtdBWqhv7DJOo2v6J7P6hTe
k9ZbqHFj88asAEONvl6ZNr88RYRa0CMfLrdYHAoXsmCCJaRlIm3+OeeNyPfp
sUBwzoy8fZCLEmN6l+ZinBkUi/Yxw7W+pbLcuXmySOlT+VXfaXwCV5jJ6hIn
7A7S25HsdyBqDw6tzyCwEtHFMK7VyrZUd2i/sBa5aDbLhQEgwa3wLPxtWJW4
zd4AJBJOPB68dY3ZpljXySm3xYsY/DtvKBcCOsNuI+aut4Bjlf6BGQnjB+DO
YrhyxINc1oeIUoWp1VY9AEktcqA/e6yEitggEjHakeT/meCkp/T12wrJ/Enr
Uy/EP4iZdS+HCKV1BGvwnVqw1M7a0C2ZvlQxYEcNxAg+1hNI/G9X7QGLXina
QR952xIocTg31vmQAjhyUhwLcEopagTA1FksuP1EWMCXhwbVculYbG9k1fEQ
FjnvpPOMcbJZel+A3brS4mgSOFi3CfT94saWYIZPTtWqsJ3Ml+M5FdhJyVtt
Y6vunCUn4FuXfqJbLo00IMUGxABZoVVeJw1c6X1EW8SboYcy+8NE+TFHollk
LuUHPE7dzAP2hQZr9GmUzsSumk+rvB5B43LIIlixETkrjit/CU+IBCpvsBl9
CTRdBaky0wkBNXLRcMsCQ/eK28fou8TvXyS0JHnd9YjEeUCUZvLTM3i6G5eV
6gWJlqYxcEhqiRFpvvTd/4B/iWeGVe9Fm9FNFFHNXhp08Czg32InZGc8QZ3q
92KUc9XbixMXN46bdvgHp1D7Vvv1oZepPziEZxrmqlhtxA7Cy6kfIYzMqYD9
NCm1mx6GldNUpSkg6lrIdZtMoOyN52x6KhkLM1QZSXdw3r5007U9+hpVderH
8SLTovfQ3hAzp7JQ59jsCgl63tJuSsQzQpfCkJIxfIHcmmBS9anB+f+O02ty
Vsv1RVxeoGwg4NGMWpf2P/AapKvUw5uRTimP5ZocstfRz4nzM9Smo/E5f+kG
MjD2tUPhW3IWYJ3mjHztBA4+Wv+LZt7TW5bMQuAuzK4XK8fSL4GBvcYdgLkK
q92YI16KbyxtMO1HhDxfwUNZz54z0x25qTNGK3d5EgtDnFHQXIQxLfjwPeWX
xdZYJbr6SMjk4JzLBhBJY9FuXjVdTGF/Ahgf6MzLD1+9N1gSCXRWymbrhyNb
48sf+l3wQIHoPwkBfm0SE948N7yGvnR+Nyug87BA7lb96uGlnh3LCG+HP0vj
/p7/8kxFq94jP1aREtTO0KXuQDWoNeTFRniUS3k2yYrtArgN27qcccjOTDTK
SS3FGa+dtiVx/56KXZ1utXHOcKSY+5Ro+JSckojXogOzOMCHdd/Rzj+EvGo4
T+CFsEj/y6lDwNqNmbBpurRI/tPhAXCczBY+Y/PSHIOp1RsOY0niqSeh23nV
xfiOBV9tBPee4NF6Ho2R6c0DEm+zpFzQ6xXZFFr73q9q0wqj1gDm83HUd+D9
SDiPg7IKGDkWiYCFCDfnyO4DSESXF4BTu8uiwtRHiLggPoYNSqyBjVNURd4Q
2GqObhS4vh1Q6jCTR5WikaQuq6jiXFC9m/6M2AT0+DRl4OYVv19LDVb7i8ca
apI5oPV0KKKB1baJ7GXOWY4lvbGiVn3Oa3N0S8jLhbu14dZjenMoRMUcgO5I
hscQVx3Hg8LVYfRtzsXoYZoEAzV83fIy9jSqLaiDo6+JJl/7CnkH2+OCIWsU
2Xq4SI+A0T3sHw9MejytNqSPFZXrQHT/fDG3M/VzmzPY/HF3mZGbQ7Yiu4jP
T8d9qTnMPJXGqUYJQcsgz3JybOiqBcsKW0j+oO97wbhe6u15Hp0NHzQ4C61I
+Xo01msWLByS2ukxg4VkmdQpspSMLNf/cYyA5W0QGb/bWmG4b+8s0qJyJUZm
BITKkZXbRaJs4gX1J9syIOFP/WSDKpvCk8U0zQYYsP68gaSScePKGa0Ee8E7
n3bjlYRAVljT7ndn3qOPZjVWRxwiw9w7TNHnkJjjWQ6DJe8qFNbwHVdce4ek
+oI8FQbRPnlCv9C+boeyaocMstUf/wPWndnYd0Mwn9xm+WNKtG//levUe7lw
s1iQYkDfdYkhJVOBR92H1VvDlaPWA5BWyLRQQ9ZLA3YphwbrXe5ENQRMGJEu
BPI8ibK+LEH6Rs3tiqltkSlTNWzO3n0KCZIWInqw4wx+mvipb3j552lzCXV2
XHBhqVSJAUaNz7jI0+DuV2BS7nSamN1PY4yydSo3WdJwh5YaCBy2tUYN1Cyp
lpd0lRXRLW3wT/MD1v9srmBqR7HIcaNwV0j1Q31123jWYGG5BMYu7KYboo97
XevRdF0dfACh2RIZPouhTdMzCkMbIL2v0JDake7/FPxXEZHu+T0bpXWUf+so
Fu1qFy8NWtwbHI2zNMNNxedxl+5HsiGvVKLK0cFRKUi8E432LVQPCVnV6yIn
MJmiolqRNmvznmCk73ydkCSvlpuCALG7wy5JoJZgG7YGk+vshPUyD1T1SNM8
7qQ7ahlxnODz+V50GMsduuGAdPvJFvLpQ+iRqk0PnegFLjEgUqzwI49prgEo
IXuJNF2/sN6WKcPDcciHAUjsTHCFhX0B/pF9diUsjytY3ZBW4XpnyQ01Scus
Wdq38KvE0MmfDo3EJvvScCJ5Tv0G/FCh5SukhXNTdh7bMJY7LC3VKT3Z6ZQ9
JEoryb0z7eyhHoH6WsBVd16Mlck4A80WP134hT0njKw53UzSuCwD7bof+OIG
CWRiLJnRAfoK2Say0K3gflm81bmALWxQ/jLmAXH9yNlmKbwADtAMC2SR7ljF
tO3/9lnzgN0nYEOyXQxjh1jWo75R+7tFdpb6Kj/ixJgpzb5HnCM0ExugdM3x
YwjcmzX6khPtL80/TJMZYkHF1RM0NUSBaQlBpyjQBj+AZjX1/s1d7ma9TON0
uQBj4uP3w1TKA5A2TvoL36Rd8gQr4idEQFXM9xAvEKTsVvHbWB+0eawXztvc
+yGkqXMrnGGKYOUGcsEVMBvriv01pJmb85id8DG+iBhUZJi/yGiI9FyUu1e4
faHmXSZnRYUuK2Xb7xiVlS3u8keGVmenUMhTJY6XvzjOwRs0fiaPolzRPkI5
LqL0rBxPk7RyYuCMtHVyGOkvAAQj0BJRC/PSp35bvTLQ8quy49mMw7agPgNA
sBVtWVYZ6neOlBdGModJom4Ms/Oqh8h68pQi8sq+j6a5uKWuMR/fBAMAWAm9
xTL82F+HqV81CkQTKeZ89RMp6f0AUuuAR9PzH/4iTDZ6WhwLXK05kZjLk/VE
BnLS037Hl5Ppoj8Wxk692JgymaeT0iqE7v+GAymWkvuzrO+deiW7cF8Zw9/U
jdCtDgxSRc/hzessdtIBmj9786dBcJtm6hz9vSBn8npYPIM90sEUJ32Tblr2
uFAzJPyz9hvUTcYEP8eG6ao/qSdbWIhKC0CqWhTVfACr7tvexv2FyBGFPzsG
9g1mFhHKZmJ7wkNrCUR/Bg7oPKAafKk9Q6l1/5Uho57ltOZ553cYNt6a3y4H
1vI5lU1a1kRZf8LpwurXM+iOpkqeV6kZpYBbdnZvgDn6QBLnz/wUfu4VTq3X
sskdL2Aupm1gH0M9btYDpVx5YvD7xKpbnX3eA2OmJJK4sPhByTmDu78ZlUnF
FMuvD9C6bD2xKuMZspPxS8KMYD/qbivBLbk4QUjPkUmRQX9co+FmdjMAkgTE
cctJGod+6fdHRc56wUFyQpPY4l+lh6TaiJdMP8p+NdpulOG4+ELgzgM7tDaJ
mXMipFZLvy9Bv6ZuHy1spBU9PxVJrrsbyCRKW0/QnRnEh2WDuParwVbzgin6
lGUspoUfzeBdl+QnKwYbzl5tQXxBB7iINnObAQW0bkWdlLwFZdMR8QGRz9Vy
zkOxMwzuTCr8MD4bKKOnyyHUgJ0LLJxk0rbVKr6nBg4/BqAQJl2W3Fxw+5gZ
7AmpsT9l0jDh3K4mZyqumapjd4D7ePlOw/Qs5pj+DwsCD7IHOjxl8QXLDZu1
wEEquZQ1OqOJr1AtSPQTjsC0ZIO5eBfjLM0sj27SFHfjqohIM7yTfrZJZQo6
100sMe1Op7gXAN+Cowe9+SJhMoK7xtb4SBpeD5xD1r+LrtNzFNEpNZk0Bw2W
Z2Sak3ghlNxskrUpbEDLU6RZ9clB42rWTBuI+fGNNaM+o/Gxe3fPdEU/03qQ
k2VycNPTfFlSW6ekOzSqSphWqNbDEpPCk7lhKEYrcEbqvJ9+yh1nDYCF0vBQ
ZosoFUnO+V6DnESELHPzyKhJOKViTzD64K1wc4rIxh5g0zb8g4Rff5+UcK8c
PC4Sb+OvNDRcb8jZgRTCm7eNMfX8n5E/BpfUJWOdDdN3JOBv2nJtWOflMs5X
DZ3RQc/UCFaGuL+ctvV7XahMQNe9JiCoB2DCK98Upt5Y7rGoxmGDaT0Rq3ln
vD5pCH2Gs7etOsJg3aeIuXkFdyD5ezEVrWkHMCvwc+lBDvYfleybqDYL4XQa
aSxnWm7n+VsDZ7IVtkuK82EMvhC76eHcj/kZFqnuuRmAOH++uIaYlglqTqXp
6JwtI8aWMOydGPCa2Q21gyDcoFUxcONjxnbkZ+eaMRxgsr6tmFCZwdMeR6dp
WzFNGZawJu0y2cy3EW6lkzroN0Z3ur4XezstCBhrQ/6ZYXPtNc9txyqWrKoM
IoBi4hZKPB4/oeist/suoTt6t843D9OFY7PUPLM8KxO7aOzrXqQC6OQ/f6od
Ep0dd9LSNOMi/P8ty1I2zQWHIkyTriLOu9zmgIeW4P2yqi0uLwbk1BuQUuTK
WJTJb7JYw6Fz4XDqBYHxsZqOEA+fh6udtKYSEx/Z0pXlfXlN49hvQR2ULBWH
5sYr4qFQBKxfogutAI8iwrBIMWD+3VZhGZ61INVrYULGwXX57wtbniUY+WGc
TVZrsfifNcci39l+SwEWp8FhV2nUKjtA46MO72xE3mO2QY/MuWWidBGBAGH1
Eyqni1pXWYh0CE2zDKtg6xH+mL/2JYVe14YXLtOD7/j4h8hCAPhRg+rztX8q
oDJ5xFSHAo7TPHgBZnaTT+y7/6CnYZV8uJskt4UHjhlR/l2LvoNDlRv7CGaT
VAFGsPYCqsATBM3YSfPFPge98a+B4CdyEq4b+Dp2dC372I1FVhy/0QcJpn/k
opW2m8uX7ZCPEU0My+mxW2cz+L7UyAh555AmgRKo6yPTP5DbAB0A9MO7VMW+
hZKb/Vs3OlpTXEQ1dbugjzE7K32kDPs8HRfXehKDsbRdyIzi/M4JMkHQhUQS
31whSOYquVkJUc1Jnw1a0ikNbWm7bpn8SVNT1EjRur3m4CDEVTSGtKZMuzue
8ey3FrMkUVuarM4zEoDhUPmahiWxe53NrwMjReQP6OPzPESvDmbFz4NhyfiK
oVoJcmeXh+P8T2XxilFgnGuBy+mU/UMlda5+8oGAtG+bsF4QTFbuIyC4o0AE
ESH5FKwaDYznrb43tjpK4mUV1aiLaUqaCtkhpOuKHHtiUeXebpQKob7NB4qX
s2Jnmb5pUmsInxq/AH9Six3Elnzr9psldScsDh/tPUYKVXpO0yhk6carbzDm
BCvqATQfhuUx6KAPg3FEggi+/H/koxDWU0Kmb0xiwC55Rt4mp9+791Qbf1ys
yaKdvotFOQCbu0k7ItAeIDgmeR1sRRNpOu171BmBYqpgB+qzoOtaE5kD8u+X
4l2CLgK5xHahp9TBqO2ttptPlMIXW8qQTx4g97JIeRM+OaRUdkrFHKE2Gs9s
KhykEF8TtB/eBIXG3ujwvsbNxaJTuXTx72RM/2ptXVZQAS3phLaAkuZkJx2P
n4zxQ7RP20f1Ni33aaHqX/c9I7hWbJRntGKrv4AZ5ePzuwgcSNz2FF6nRXBr
8ElSDteYfR8fBKfKjkxvztSssrAgWBjKS0Uxa1Bo/4tmOxxm+aEJ1f2mZ1yj
HmFNkjc/o8IC4+388CfyOpr0kXio1vpPDwYq9npCSJuMJW1keXLfeKvffueg
p+BWiN6SjWqsVa+kpLa7zQ8MiOx4zux3dXOYSADGP78D7D9vggwI6uN/Edgd
uAZ0ZsBP9+fFvDh2rCF+CYylBs0KMToAX2Ol1Yv1mrxBTZeyjifccImu2r9f
tJM80nIk/zvsZQE6drLi1v6OpmDv5SPw57Unme0e8LeTg1RcURgTgccDhSOf
ZlkRt0wYJFzSiTrk74/KTo+7wtgPYXeKMcLeWO96R1EN7Q4hvSIR9vVCIpah
WsyzIcJFD4G0n3ww+aH0gW83TnT7UwCB7OojEQI8E/GfFowxEundTnA6P7Fg
+GmBc66ZBCwMncgsXj7nW3efLCUaXak4tPoY2e1IAZ1ykV3H6HckMzuIomrl
tlYHf6r5r7slH+UKaSZR1U3WFOzxePHJgDt1nGZ9meLXqOTOmJVn6T7Oj9Gs
AkWGd+cIeVo+/7+3lA6Z0UYUbJjsoGywfP0YeZM7l/Qs+tg1o8ea1A4FUHmx
5cVxh6YukmSeBo9EL72bDS13WobBSBQ4Xf4J3XVKsCnhW5vuBw/biQWOdNPo
11QdwmzRQGY8aLAIuSqeFl+RPl/EeOT5BnWDEhADACUZj9cwhV7Sj60Jp5b1
R54s2o7eIBd+xot9YO0jQObOkOU2AZqeWSrOH84s5GMzJYDLDOyq4l1SWwBL
RLg6OfMRr62V/N9IXvJxxov9PVGn8Exrw7gIbSCDK08mTdFyYPn5GBbQwR1s
s624jFaZQjCghgGbvVELA/s8wmuvRt51YSnCvmu49wm10xqxJSESW5gQBySs
YQiIA1TiWMt0SC5BsiJpLQBgSrsZ2UsZXXoqpYRWyJVx0j3lDp300n+uyDmG
Ibix2ddi8DZlzh+8poG8ppfn8FgvCHs5oXJHlGlMYBkJgsO5jlVxSYIF/Tf6
Ar64EYldrB6vt0ejWtLHAeR/CuwFC7q1Xx2qL5A+F8HFtSGLVgo6E9Fvc+om
M3h+bCbWsyoJJOCR32ZzrjmqkZRWm4KKOx9JE5b21DECaUJ2kbQoLjfGwM8c
07qVRp2X2FaF5Gi/0mXpfFRTbR/F7APAJh+MmpXLQZm4RA308X2cgYNNLNEb
3chNIT2QCF3rKDlkndEnuiIZbJmo2ubl35CRZFFhgbnq0lXppsK86HHQLt6x
jywh27YY+K7FQHAG3s4+4PnoYNaTELMoDS6owCRADim+eTiyroJzyCj1b3aT
wCcYA/UxKy734ioKL5glW38RKrB4PaNfO66h/ZrRrSc/7QrUzQyTGoR1djz3
MDLoYB6eneZlrxK+0hfh7ZSEEgzIHVZr04Hc0pIHNUzkjFGb6UtC+TOmyHw8
QMF17Mmpaow3k6pcf6Ki9pFCz44gBPJchBfkCmAp3J73xPIvMkaVb23wa/af
xWYgbbPifFKvep22Vkzd35GYbXdjlqOhJm9VhjMMZOxivH/qbLlIszRQ9Kfq
oTYsUanBG7/Tb7/oKQc3h0uqOSaKJ6JPRVxKIDs501hd5PwzBlsJOzMIOY6l
E3oWuJoMZmr1mSSUtAnb7/r2UW+J3TlR8MHc1J+bIx7FuBGw+Q3wC3Vtdjuq
niG7RrcOwAX0Vx2GgodPoWnU7ZGTspGLTKIIGuWYXDaRc8YpAlHw9S2qlL5k
nKXX7fkgYd7i8vAH82jVQKhJmbbVF8HAcK5JFRqekDfNygwRXpbkSPcBu4kp
x1Tp1ApKTrBNggbSTDtRDlw4+yANjEAhGNKBscvnwbOf3Obhfhi/rzv2Lg6O
SwrqUhbqyldSXcCPLHhtd0LqkywAjP3XIL6lLj0zzhBEP15fvNwEluq3Qc39
4N21g7kW+KQ4i1NVwsA5Tzn2TweDv0Fq40i4/vjhkjKGB8BYvEhhWCSa5Onj
4UYQ8CWwLNrGR3PTiF0zG4QlqowP7hLl0HBIfympAyDG2homheOUj8qTGFXP
LeIIzHnT5L4AlfdOB3D8DYJJXRyZgnBqQiZoth1Zq3qheXCVZIty5Ky1kZSs
QQ6U+z1gpvaCP5ydSBDl0BPfMf4MG+nb3QCL0sSxfCE+zf11vNF2ES4o1wjg
3E6piTQX1gBPzw8QZUjD45WqvEG2ISDzuQWyZCKzHWwtj1uHUpqFS/wsoRMv
6w3/Ky8h68APNe69RHrabz0SsjZ9GBl8s4K5ZvCFgdXmOtugDZxCLGbjdCgO
Kl8g/ROK24dKSR9jSgi/72Z8Go4r7L1qMEApG23ISuG65hJKYt56mmF8G8O2
CtzHkhr+NIeY9KZ4t5IG6N4GQaS5GqYbGfxJ0SnnT4QTQXKTA5d7BWZiiFRJ
07Tse0yiHP+qycVzTWUuQSE98wuJEjyxADoK1jzYyn+nxeMhHGc7Y5BvqbJ/
HTeNROczdma6XIDY9f+1VD+siV/T2IQ0d73Tn+Uv3Ac+EnTLxEpy+SnmjM0o
oEhemHn3e6s2vojdvgSEZTFBV3W68eSEy4M3Ycjrp7U8EboNmwGpJn2hOCmK
wIwTEpiGLuYtkt+udySPIwrsXyRVvSarbxHIi70oP8iF9IBGbqkdnvlI99Cp
H68Wie540VmNXIzoAuSoWzK+i4wIjJP6snpNdHhFx7oU4bzsjqvk/awvkfyN
Cxm/CBQUkmsPqn/tPzNz+X45zQZ6kBxaDkJiZTR5bzbhhLDn+0anusqRhEB/
tfxb50XWdolD7DX4zjB7HY/OhvAw7xol8p5xCJhTWktyCFDUS1I/gvpfmEAB
Jy1y5IkUgZV9N3miB4/VTuysL/Cm+veKCk+zQCNxK6UOLZpAWnvs1o9pkSVE
cM/0hfS3/XVPZNUsiDC92gMoEm8qzuM7hdBPGuz3+oTgzVtSepqTJYl3gQfD
A+kObSalWSwaQ4Sv5DCj8TB+vPI3k3qF4nyWxWvALe8gdbTnrElctJCFkOtF
wONowqWFtGew3oHmugo1RY3dS7cao2eUtquL7gnDr+zsZlSRF0YcA7LYdsvn
P+Nc7ocWNFp/E4ZAlhnZ9myQVtID2cPoEa0pVbUBS61wd8gmhMCzYC14ECm0
A/yZMG8xbxJXuq28/V3tvzjhe02Vx2fWVKdVWSWFh8ZxCylq5rubjTtm1pdH
v3vwJf8J0QsjGma0mDfBETRSX5VmBRADUbPuaFxZSRGtm08HguwcGyo5cKTK
objd6ODius65TT8OneZTpQUCNvXfIdZnC5c9u8EeKblQGs52eJFizB2cO90F
1v+zf/1b8RnUx0ggnEfBZ4irn6vx0mXnGya3DoT3LtrbLY8mZghu7WjFPrWB
9n3bvDZCWCBXpcg0jhs1xxR+sAmWCiEe/63WYEAcmP+X7Us48H90r7mXPqKy
9Mv0z7Wzw9knFAUZR5dQIG9SLfLbgf/5ejZaptMeP9PZVYNzWL9BSEW/qkl0
CxfPb7+wAaJCFk8/vf2O4hjvHgfvnnd7BOVGPF7/JoGS5NLMFyfIQsl7bn36
rXR+EAFrpMI0iZw4ZNTRnvh9DsSrwOhZHhdCWMPCXjTJHGWfkbF0OblEbbUc
XfCHQdkGMQ97fNf/KBqt3NJMzJmASo7sROzQJu6t7gZpM+NFfbFXH76hpzYU
A7+N2sFSpu7IMh6ofJ5tJDbU+o9I9ZYJLQ7E58DUOmug0/4NiRfvvWyKqwxs
xPqrykJYOKPSGNGu74LbGDco8dZHhlOzqmcVHayRiQl+Vr2LEKOBbvSvXJOO
E9oqBYVQgPGZHDJwNGQiB5MmFqAEtkVKJurtVq07eH0cP5MYvzQtTsR4BfCH
KYIvUUX7h8RTH9PAfOmGW4dk6js+aP+ylZUWJi2oIvKRja8rh1kzyhA9wtK5
TzpogTWcRQEU7JWJ2b6tIu+lmYnrccmW6+yVrpGpEWGLNAb6uPuJbXEx0Nqx
jnsRc7UHLpAxtooiEbnNaTzxb9pXkSvHyUTrjzBW6rXXGinIEPdeOJxIJbe9
IDCaOz10UX2/waGNSA+05ijvgiXqj7QHqfD3d7VmtM5UUnq3PcPbxAjG0ooU
qfd3vcoyYi1VMPsMbR1CeRuCU3Gis6XqUyPbu3IEDDg1Vjd5ksLSVRfK/0nV
Kylepppl8DuP98nChmHiqAWUfF/gJjoUP6eIQ7AKnEFrerKlopgXweO8/nfM
JXzaDZdi6fA+8EzysVFbTuJt6vALg9BoO1bwTmVSUP0qasQzEyASsKulIvLj
2bKkgTugHA+NFJeuZY3C3BX3Yx6JIuf6kZQQwE3aCca6Y13HZVHMTjg1kv5K
S0PkHTLOv1VJQoHChUxpSphM+swmXXKF59a0b2LuUwiSor057IdlXViH9nUq
B/J3TahxjhKc4I9t3h+d5sn+ti2WAX0N5WUpe/3XqZzsm7n+/kD8bzLer3Ht
WTVkYzmcpSPldihlbxVRv/R39+zoQe+E96aagIz6g4Jc0jxtsDq8sGwhuCq+
qbKNaL3RCy+YirBOCS1SRaqJ+xT5O2T2H7Nh/jv/rc8P9n20sBQzHYXw4dlc
o9nh5AiO7CQo+Q0vEOT4l9IPVJjBddYInRD5tdBP7/orpxtTcDX/bl6KGK9f
o26bRY1Tu+UROpAgB98N02PJBzU/MZEjsE1nEiSC6eJvFM6pQdPsEL2lzmxU
hmLWkTD7C+IU2hkPSUu7ydTNTq5h+u9FuA4nuMtfiRRa0QsXjaH9+ODsXiX5
J7RWRqPBydZNk/DT0s0Bbnem5rbI3Rp7AE/evculvvCUAXvQ7zPYHzp31PO+
mVFp/KAMcaD6zn84c7ZKjUdfH4vyZr3xudvgQun4+r6yLYJJazCfczQ/yuTL
CHOi36j5TrtekXKcBRvl07nIb/sDGtCL/mpu4Qsn1yeqB80EJ/VhdSao46uL
iBGijY+OAKJoJdEBOYwS0+3JNUawIZSUo1wWO/ixj9O8lh37fxb/n4Szue/h
4b2qTkO4dtWd5ilIZEU7j84AzJdOIq+1T9mV247dGbxjSUT+19mMe4L2eqp6
UznjtvZEd1E3KUVZ4M11wl5cwFup4+rBlL0zBJiKdyNUthHqEuIpujy7QVt4
+7Lz92gYVXrhtolh7ZVQoQ1Rd0rAZwhCUsoNlVBnpv5y/uRHiRUWErCinCdV
knCXXSajQvm2AoaCuP2zspz4tU3LTOnBrAbLVooXZ3wYyTBfV3uSizZYvziY
NerJsMCTGpEpCfzHvaR7NgVpS3bjxq8kXUtB+/1ybrNo+Kf0TBf77hZds2RP
jsGvU/uI8evK5k+G6uoLHAzkXCejemNPS7aDQ6WvsEFxQSZN8I1vjD8SRY06
6RASmFd3LK2bVTC3oRG4EMypgmK3VfAxSGhDJ44eZn8abAw5IA5knQRgZh1A
szSpx7DBgYZqB53BQISyHbKXU6Q7J6QYZGg/f960E57/UGzpYCcDbRTKiM4o
9fPwtEUmX4yW9C7eRCJ0fwEv56IDZvkskduCYFbSNITgdzVnx6yRdNtEyI41
9V7hFmig9hyjSGlT5we9XCn+EDjkC0QpEZpDx3NQup8imCXUajPXmC1AN3Km
XRqdUFj+qp+idXqJ81P045yWmxDnXe3EvOky8vAuOzSZJO6ERun3bQPANte7
S6egzb5MROTvtsdNiQgK+s12XTzmwlYxiQVjf2eKdAEy93aE5uTefvFy9OGu
kZvo+9a3jYccTAJ+jeSzwMxZ8vAY/A4AFSBE4Fn/qElHmSVsEjsYVJblrN87
U3Q3ykcQ4pLJ0+UtxuNKZnvp7be5F9jfzLXdGIgyh70febDky3M5H2fdTbo6
x3GpeDSn0DQ73j6+rjB2LyYzj3U/l6/vc+dZwmHWCElmDadeMm5syT1gewVI
WhAmpKORjZAQRmwns0nI0xOjYVhFt08j1MfZjJWylaJa6D7NYeiJUQqheOMd
mMxRKgo2jkBNwzLF18f7cvc1653ttx8rnJ+9rGOnZQP59FmQ0KQKPuq7J1Un
i7icVgTbjqA7ZLaJIsGKTDuMPRxc096YbmdUDFHs8+z41YRdvDsLWRapJnvG
dc/yQurXCSBVN2sd6goZSQEBBwvTWm4G7U6wvSnCC8BX44VRXETdrlLKvsh9
UK2V+RZhC7rGmwIg+IIpPRdYXrsuWPwiS+wZ2d6vsi0AKfIJonaxXCuevwCW
gAbALRnFt1yu7FA7lkuZ7OSjaYEhB+ptaBJm6Ik3XWvbMTkSoKc8A4E9apyI
bwKp2yZKDarbYeRu2/rlVcK0lEBjGrA6AkP5PFoVF/Wq43XMsKFVTP5Nf1ZS
rW7Jgp8zMlB6LHIOM8yeW4IbWCZ1WuvLvOAAi4C9hQ5mX4ongMlN4+q/XlsV
F5ojNHJ8ozAxhi++Jl8R4x3LMyEQNqL8i/1qJhJW4E/7lkY3IavNz9/wLDpM
y8Tot0qnls8Othr3b2U6GkYYlolqBQYZuj/GDr4zcRQKyIsrjlEM45vaHHaA
FX2ksimVftRHhhnrnLotYid6rMD2rSS40N5GbpVJ+ENOnEVQxnp8NXn8VmXJ
/z87gMtiYbrWMRReJHwRe3VsYYjLfeAKwsqaHj4LzPeIwlwOn7UFKCxQmeo8
l8AUfPBt5+lBhsNAU4LtQQaHuTFQgTxk8S+g61zKKtWP037/d8xEdrwTvXoP
Osa80/DU+WjFft9ggwYx5cbnqMn9wLylJbWrfTZkj+7r0Mq7gBPbVOsGDD6a
6S8Grd1k2/qqOt3GAdZ0h5aYLWIxDAtLWoyYsSg6aDN995m0qfGIzbt7oqBY
7Y6H5NIlaF4TqefPnHa0ABT/tIg0b5vOJRUpHeBXBNQUFt9QK6b4+UpYPl/H
mzHTLxKLi3SfwSvYaEdbg3RfLF5wSS9pxg1s3IE9yeq8ij1A7YoMUyNm0dwt
UrMVcKvsoatZTboUqXmV0bKySMJJcwChJIEUAyf7J/mAGLsk6VvRhVidd0gX
CCR2m+GuaAq0zDX5Uzqu6u92e0oJfWsCLq6ito9rUP0goowJu5RD6CCUijEC
fxX8Pgihhu50/B0iFybI0RX+MGgh8zIYGOGDwftWlqHNKb0JP9ki2wM+4nrB
bxDNQKcffSnU7EOT2DggHEMURhFB3PQ26LEZNbtygSKCf6D2NsQU4tSn5jg0
XK4X1xlDncI/LYB4pHGPASsRxlqNGFiUodBPjpos0OzsR8pTRM1G32yc5eNr
X9xN0L/5FN6tAqUuY+MQHxOiWB/wI4+ZugBjL+BI1c3Yd0vQeSVLM4pYIxQy
Z1rIFzBUboJ5S2DgNFxySZiKxqPQnot4xM+O1Hv+IbvW/heuroTDyI2yz6TO
W/cqd2aYH+5ZbJ0unfBc1UY6nsNGNuouvIR2OZYz5Zy4MX+qIss2KWl72pdP
FuMv5HbGF5t8LfP7z53stLr1nPW+gCuIFX01xyDay9xrxxHqDzy/4lBDSCvc
LgsmNaJmTviMBbXhuBCvgIzl4HsvucMitsqCoDGQo0fe+U1fRybXndmqF4Lw
YmSIh9bB0BaNSZlybfmCkKxFGMwjMZPPOqf9B1bya81j5EVmBT2GIdbQPMk+
UljTdqSMLQLtu5DSu0ctho3wFMeJ/vn4RxcwgoD65oG9uIEytZal/u/3OwVS
iHgRj0aLp9KZfVDfx+mKjBHMz7Mji7RE/Kp+Pkk85XlRvKcITmxhjsnlZBid
9xXxW7VPWl47sTLEHjoQ7SE0HdRc2QGddELkBKu0amrRP+W3DplJaIzqMdO0
3ZQynYRj7N80Fh5uZWSKmjuargFrazAdyx8ghiYBaZlRVVYYUqkb77gVh/Up
PL0boioSEMzO2g3y/qfgdVQg3J04NuMyCCVQhZ0wAdS+KDP2Vndc2pX9m8gs
09MWpU8YclWDTaVRuzSNQ0/C0ErEh4+Rh39t29KUK3tJX6xuKWLMutpUXpy2
nS0rAZvHAUonha0VwynQOAPz+ycytmlWvqtp+EkeaUVXYltVzZAspIqTdKW/
YSwc4UamkvTpZgoHTlDrdfVCuL/K+RWrQH3wGFhbgWsPfTnoYRb9U8C5+zBZ
872I0HU07FkrdaBb85Pjer/XpSejnORhHJhK3SQXVCtnEhx2JiJYgkq/kljt
DACJvU4lEmAnLR8wel6s9kmDWSwN0MSrMFEFmBQJjoExK4iZUlyRsi3t6eIb
G5ciPL25itbb4HiVyzHOem5bmjH3zOhK/lQEaX/SxEoXh1v30o08/LU8qm2A
HD1NQWPwQjpv+DyXgvObVcpPp3hdpRweIEa++NN67alVO1TCjqHndqJfyUAW
zV0I2l7lSnLGHFfzxdYpYVSA5w70pMcwu/7DLucngAf8/Bby/mkGrvLsFe6d
xvfhPCPnz3ZNd4HUKIBTummJH5DbGqTy6v9b59iBntIdT6dxL7TRtJhk7eO6
FA1WUqmi7qxDxkTO3vBNhqs8EpoDFVdO5Rlya31wPe0MOoy8+C97B8lSfmMt
QoYHxmi0nB9lfJrQN8kJVThK1gZntVGziofuGncpqNaPXgE+Gj//x1DnsYmF
ROY4jdV2GXfXntTdNbnYu3yoZLQG8EuCQpIBJZAB0pb7gqoobU7FLpuTM5eS
+TLVFUxss7w2be8GyvBNTTly1QRYMgTYszYBJ214fXSemuXgV1pFUUkMFL6m
6itUNzK61b374NP+NJoyDlWPBBeDoXfGnssBj/xv/+1rAFSFU2KTQowby/tK
HMQP2gOoZlCqy89pSkuVLUeYfL9F8fJ6XJ9xVyqf6zSVZz2z28VOVN+JiunT
Lck1yukpFbWNYhkYUBh3pTYU01M8HSHzbG6r8AONvJWviJwoZsP/Vd989z+S
0p66u8baXqoG3VeWgtgC9TnJ1WhrOk/tUiQcBA/ZpyjsbfNvzzzymfVmdJFN
8ByvrubBtTUn3bXKBlPDFVz4Cs1lVzZT3wc1QAcALK0l75PyrASmB4zeqlPc
2klTSdK5aG33sPc8y3zUJKCAN8UmezoJhwV4DfKWE3eIyx9Z0NH9FhkKnfKc
RSEWwAFQStUtUst8ktLsg5Lv9oY5mBarl8meDRxxpBhSN4U3Vbbg+dbvs7wd
aoMSBy4r9ll4ZoAwVKO7/r/GasyQ8XirhMUsTENHYJ/YnGkTFfsLYkrYR4l8
Sp7TgblNYmzDtUH1ksSVnk2jDunvm+Jv8ceQ+mg/ZLnn/USBHuqlo4x/o8mF
iL9VdX8rQ3Kmhst7BNEZXywNRydD9+ed2qZbuIrT0B0ZNYcmY7OSpvDZ/pNb
5Bhd2fWfo1nJKAq/67TgWXj00qY8h7b5YeTtdAU6i9oY3p5bgGbhFnZE8jfg
TApMn7R1/IMsilomiqrULxqWHfyZiBIxIVqXXD3dYF504BgIEeHseJdMt/jA
gAL8m5sJ0FGi0a+hPPwKvnBc62M8NlN1r/IVrmNX7i7ByYD+QVztVL5CGgb4
aW1sqXSkNZuqt6qQy+mD1WFWb3hXgNovw2bfFMsLIjCUvUsVCX78ImV6hVj4
YKNKKQAnWFgGdwaUUErXzTCV1SqALgVTFR3Pl7bZ4YL8y0rUWjG7RHjrySRu
cxkLHWmBqLexHM/b8bTgnIoMzQ9a2v3RpU5qqZOQrTekilZQ4JPBuxW3oRoG
u/6E+GuTsFoBEZOzgLaMYniQcXhvPRLinEal+FLvpcmEzsQJ+C8ahwn7Tplg
vE75B1HsIC15qtmqM9FXS2a4XQ3CO5cf9HsqPxz/ovpwcpPCJie91Er6L+w1
YSRDLKxINvnhjADVrixi3pDGms9diNg7DyywKkTkkrSzdzvDMNXSoGci0ULc
0gkZVTjkvznAjBSmOQev4iXOyjFCKivtRS7ta3KY4MC1uZGXiCv6hqaEFgLu
oIUSC8VQ4hsksJpu6Uc4/TUKseubX9C/spENmibq//vvtO9AaIkF7qwdrmls
ktjUz7fCj0lIpHJyrvr6p6PAr5GpRPp/IyS+sNcWc/CdsfhSAgmZqIGnr1YU
ghuBNl/7dFdqOocL5KTkCpk+43svqSMjY9vB2c0E/8zB+wf4AonKKPo3QDPQ
0HsJMud85Wg1s9q/arkmEKLYR+UkU4hdyJCoGYKAJDPraSRJcJNTjY3QWMK7
bi6Ng8SNfsokK4rmsnLAkt+9bvaI5DGwj0bnE8PpclJKGAVarkliN+AuWKDh
1VWYPO3ppvcoeR1NUZh00U13KYwp0a3WAZ4FQgc0KtK9Ga0Ltf+BQKDjdPBk
PvHvLdC/REwICPVZ+sgle/M+5CKjIWC5uOghe02tv52Dwg/EkukSPBVJd/7p
cVweZxoyQJLN+nZgDnzjiMmvozPDfm481+vrEEOoGygbsonmKzs1t/exD3uD
AJUts8/4imt1Dch+RaLhY+T0yAUUU/j7iCNl7Z9zHBlsLLLIkJNcOfiy6NXw
YFVR2A30/EzwH4q2hfnplyP7ZuB7mowVkbymamyFweIjxd7kqagdjxnqzHvF
LbRQsao4j3IAT1kkOndNaHCH4BjtSqmOSY2sXlN44LeomhfhBKTEG+tWvTt7
qQjeOHHsl+6iJ2hAGJTJ8na1wKL1LEcz+Ipj/n+erGkZMpJ0pm9Wt4DFhP0R
7Vh/sTvtBvnE1sG3SOc+1fKOLSXbXl1qIWjTHhw6fGPFad1PSh0DnSnMofZO
f+gw7OVuyC4MZssTDtibTZmndR49gCVU+fsrT1L8Y2xgd0HNpcqKIzdBsMqO
oPsyVLDW/xLO0+h4jRPWAJY+lyjVo0+c4FgJj9NQMjo7pN22p/r2KPBhOcck
wD5QY/7ai6OhHiVRzeSSLyA4Nd/Btq4TmK7PciyZRd+iuzbQZy6rCEDUJIEf
vpL2DbYLmO4NtOz0EYYCbWdiW2295FhEJZQLzuQftEz8/ZF3cpqD3hsAAcTW
jCebeL5EssWh7GK21ndtztbBZv57oxc3pykEHNy+5CCIL42CXt6lKiK3Xdl7
7G24lrh3G4EMTVfIDCYrQKBzJsLunaZTDwtEcinbi3Tyf+ExW7Q6L3Imt4HV
r03m0ySaqtzYELOjhiL50Ef6xKqB8JE7PkG4fcOa9Gr9OlvgEFko+O7eebpc
LJilEYhcVcRzJ7Lxb22lFB0jDlpDxJ3w81SER27OQUqR6o7IbaOdFdK4gnIm
RKEuVqyZwIK+O7u028pFjkLjTXWBD03xRvOSr2oCIEUcq7S8M76OBZI+Bjoa
QUnTujapiFoFqR8+ag2h3wC9RNkn4FOI6B2Vr46Hg2Yrml/096w018PUSFE3
yGwoGN1HYGr/UTHE0DISsjuQobSp1BNF4dBuLXfUOFtqd3N7xjI4I24L8wMN
BXKGmPVKHxiEYM36PCxYzc6YqWWszAs5ZPDltafUfBgg5WCICd9JJG4P0dhD
Nh2FD90EVgZPqtGmduUVFAhCNCS0nuSJpTKNFjcrvl6PMu6zH5Y+Vd6QGbiF
jX+628tHkDb6raEl0J/vH+lY9k0KBwCyeIveFE7t0eo4bJ9lgJjU2U2eIjaP
1OW7MDh+yc2NXuNi2jwgauG+/wK8/F/gx3dUuFdTpDIvZaF2UV+Wenkk6Yrr
DP1wAIR2OcOX0oWNqChOr4/ncDZmTMCQaz5NXsH3pNaFf6rR+1ViOIs1/iXt
vf+SkYnTnvo+9U/TGa1v5eoIJilSMVGgmPTErhfNh/RWz1s41S2nHZf1sp+9
ATggZ/A2NqzWDQrQhKYxZn5hvbmlK7u9Z6uhl1m/741fX1++buEoNYyjpZzr
Zk7wZQlM3gJ4GG8wWuDQucqEaFflj+p6y2Z2dACCV67tNqqz6A8umPG6Ojht
D7TeAWihYU9HeDzAdYU/sGEOXiav1qa/ecCVSKCe5Cw3O/vD5N2nNJTScESB
t2XbLQbfE5hEtFBfS7w991gjZXtNNrjJUBPOJu2h6Olfh6N4xeRMWTrTUaJv
Wr4wimpJepAe5tjvDhx49+4dWmJX4iGJ7H3pu4cWayPnlCKa2YHa6jvMcQUU
89CgLWViK5zGEtfZd9JRbkL1r1zpdm5DFtx/NnFnxIJr6OqlRviQcF/hnDQ6
v0pJctsKpVApVw/F/MTSZKBnFkkX3uwZqzJh1cFA+Rs2nD+fmSBXwp9WFMWM
vmx06R70L4HE5Iiqr6XP7H/OZEx14BttIPbgCwoW22ml67851G1xAZpJu4Jw
mMfjY17XFwxG6G9f1mqC7Tddgx8KtJpJba96fPzExOWoCLBZpj8Bt0uG39yc
QxMTzpJACSq2abGkEEWvgllHrbR+v6bzeUFj24LXq48geWFGoayAuK8arlOi
R1t2Pz9EcvwfQ0zAx2WFPAFteS9RO+G/aJYqsbNEaqTaZQwtVrsSCcQt1gcY
3XSGk/qaLdJNFN5mp7NfSZXp9Rhe0BacBcbKvqC6RJq3F2b+QuquyRJub7Xq
rT4Sk9gGI6yvNR6xuuvg1tc2IRk7U3dXKmiDqk4qzjAruCr0yB0TlJ3gK3NC
aGvQDyW2GFK7pZFUeZOm6NtT/JYtXKoKoruSn73zJFigkfJbGXtU49WUxscU
Q+3yV5g5CCeHzxuscVxf0tBlaLvgFbG5YaQo8jMQS/P0/VfsO2xYJ5EH6o3z
15IuZLo/mKg+0gaZzDg7cGcffFFZKz3fj+JFKyWVvpiF8nxqLgGTiVYcu0mB
AKDs6TvV0gMqooC0dH6We72n+Zy1KRs4zB0CMXzXoAMrOFVQfzz5/CtQm6+V
KOJv/hftcPFrXhNbVPLbWI9TfV0wOxAQbTTLUmFrlDTnGaJuwlc+rkGWbecZ
v9v9dLvHRg8I06PzMTlaq0WilUCaqZBcJr9xIUUlB13o7mt9G6gCLlO9eB1z
ItuU5YHORglgptU1FFVZH/WnYjEcBU8PF4HFvtWuS6TFHW+9KMVFbQbP3Rog
aePkap+2ag68RUCC8wnL4k98s+mDs88YQgknXKSTNempJfCbyEQ0iGPnJRCa
Orukw0Sceo1yULiWJtSmLdTULGptXWd6N2UiOSxRTOHG97BNG7hXpQddRrxN
0Tqz7RaAMAH0yzXRgnm0BsxGsDtZXkyLrQkP3u6ZM7CwvcIBp8F46K8YwmbT
pO5phrQpRSXFyBhQKPkIFzsYR3qKeacjZW8RSB0Y4Nl7uCXETBwDmzEyRBwY
a5I5Ps0CQWTQu5iaxJkpw3aEw4Yu5PjBGLg14aBPaJVH7e0y+GlPJUQw76Ta
fMqmRXI2BZEnLq3FZjqx8BE6tO9LjxOhbyFqAJ2lhzM6T2OdmQhmUnXaGGJU
MUBCQPIlPcIeBwGG26n++igYFXalqveYuVZjCDvniLk5AqC/Vkg3OyWwjfKE
qcnVDGSA01XFL6R66kJUEIaZSzCeoDN5dttucn72QAW++LjOgNd1cvF1oK8r
I6UxGm2oA5koOVwfQ60LmvwXQZRpl/ZtOR8WzRJ76JsbfUhk6NZhYZ6Xu1sn
tO6x7PTXC6qfOX5NWV2Wmz5iX1ZkrR4MJ88ywLg1tjHyzbL1eFuM05MHooPl
gliGPHb+lDvEaKJJRbyYnpWZ+7Wb15DjVnEai54H47WaiBcS8cShJoXVHk3G
ZWQMCfdbmI9nYX5y2FGtVA8UeWLYu09Vglxai7bNFGCrFVjkvlOZFktGtXfF
Jxf46tpZ7LY9wrsOf9mcLszK0auTYJ+kA5eXjGg3DnYIToeR/GRkBKSqZi1t
YChMwrXQeZ45rIorDH95q3fcqJnnBOqa+sKZZ4/x/Bk25zqSdWRVS95k8dUe
Rxj2M4GA8hocAJPU9AJq/BwSvJuL7hyBzr9xAO6ClBpe9KlKPfdWmGp3iRiF
V4elfBTP5TEeNXrYl5mOIo5TZsrXxVFgj5EvFU6E0MW5R8m4DxnZTwejmdrR
NTPs6LJINtV8mBEn1URYbqDmNkK8zmDiacLARIk6JvPmAeb+5Ql0hb1mAgQO
MgCqZeQ4Da5Q9vSaqrFBDFVKxElVcHe28XQeU/LaPsaPMJCr+NYneLG83gsB
0ojHfXIouX/pce/lvT/GPHJVw5YaJVy5yglsQ//G7mguMi1G2kfXRvNT9/rY
rj1Idj88Eaj83Y8FTcIspNeHvQi2oeNfCsCNuWALAutt6UZUXFNN9NA2sKtI
gACbYSekZRZL0uzojtLgCUS/rqsu6QRoELZGwODByAhn8EQrfKhHooJL6+0T
GIzVpULIezUKvxSGCo5FT4E/Xow52d+/tm/zffxlwFQcrSt27ImQ9o+rhK0q
ujCHctFIR+nphWJEKnhxR3mhNmVI6TZzPJXhg/0AvbYfaAPuxMogLNitqenl
T6DYFXfKvkLNQ3evYG638XMF8ZtqYWMLb2cTc/lOpH7G2Y377UKLhAy1VXrj
BR2Bzxm1v5I2prym2eStUQQ/puEoY78FVm+5kXWNn677FteWdotw98hJW8+O
bEyZQNmFms6Qlbqi0Rb8z/Fs/R+he4iYlV5O09P0M6IvfHc/oPeo3nzI3Bgf
cgvWtI26KBvEj2o3eIzmKjXTWcgdVHdizZDctI+HSosD7iVSnqX2uNd1PIe+
eB33QBsklRcJ83JlsdxB3cTTZQbg8Q4vrZB+ROQoO3Ayuex/ZJVYp8e2Ic0t
jfhhDU4YmDhTXgP8Gv/5DO6b6a6ico/SqZ+quUnrFzGR/2vv1vkTsJZAAse0
xzklsVa+7Ek3ts8GV+JProRdvSEJofd5AHHTQ8T6NvqYipNsBeaaK0K1nvx4
uU220ejAZINTRdgGZT9mXfwp6t5e1svee1P2LrhknbU0wKyyOy/SPphOkP7t
9hlU6LH17C5jCTGGi/I1VUERq8joZWepxBe1ebW0ZiMI8VkBq6mEiUDP6A6V
oWBhyugLDy7jVuzvW7q7up5D3D31QFSQOwTIgjDs+ALsacy26OjcMDQ9pHPy
RYwzWo+mXFnh37251j/uCl5vL3i+2scSbAwETQGYec02Jw0c3/TTZRtzcSZh
MP4ptshYwX68Yn96d5+fBvHJcvKuCIzqFCsylGFey2GAequQMb9bo6zSD6TW
L1Ec7Lucx4xTXcQLRpZ0kDIlgW1ceZPG04mhZIecoHJmAXtK0mEc8dkpovzY
/b0e7/B/zWNc9jhDheouykbs1qXNOv7FLs0aN7/8plSizjSW52vrDgPgqsf7
axqxn3878wm9rV+cVjmr1S7TZlCKU0Q+JQtZ4PwpEPfix1CydOXuOHwMyXC8
7w8/zaXYtRTdFUq73crZqlgaHgSZuyCJFRBy1LIYUMiYeHUaAZad+k4zpjyV
ORtFUKomn1u/DhvKzNVsKpLnLT+4FhD/vXRPaUHpjxH/uxsp7ChrtuqTYoWd
mnSiWfreHMyEoqaNMMG923hTi8WcFKfgWnk+xZdKLi2IYp2Ff5w2BFEkUOHo
iG2hxCGK1hH7EkE2UfOjBQ4MIlMA5Xs1svymqemwDjSCMRtjuhfJ0QhPLweB
yFisBa363Gk1XlZosU1sEedecodDpQ7Ttw9kQVuINbUmy+wdDZw6qqVw8TlB
5z3hPMiaQHu/NGhCjVLWByzyaI2UOa3tXzj1bkNd1jvue5fIq+4xzsiXISXT
ODhqX7WwgdCwlIG+/LPWG8kNMq4KTFZvf6J5k36hx6B9uwreP/X/NIgzIDRE
LJWkEFN0abfJ9IPeSgofJ3xuv4KwiphqYyYLWRcOtMd8rekytLd90aTIKLzt
lPS6ffmflmU4TSa76zoM8O09wXWznrQV47G9nPEWTzqCUGozB3spNaijuzab
91BK5jkoQGsnhTYdGCwRiycDgfhR+prwXRJk/dT8JvWjmMKnKmHfPvyBM9WD
iIy35ZxYpTeinTR2cfHnkl68BYXOZb7IgdcLSqYj8PfqWrdpaHYX8hWcO6Dg
d5/dsmz6O/muKWVURwR5BF3Fok88BxIGCBB0W7zCZg7+UJH2PWDraQi0b45m
wnwsRzHIyL13j+OVWdGsNe4TYMoR/GK/edDZm+XmgsktFjsYcnl9MkFDJHT5
hpiePJo50DrxyyDt7nc96BITy0ZLTNGmZ8j19Ksl0ZhsPwxTQlbsneh8ETif
pKJOXrBQz1s4I080MpVz9uKgPudpr3Vj/pRLQmUZq57hRYDBA7CUUgd9Aw4f
+LWOzLDHxiDFd7DwWSBl9OSl7OXfWJY2gYIUCwnjJKfY+NPXHupoACar6YKg
KvJliVd/I10uC3efqTLC7dFLPj9GaNqS8mCcKHbzGPeH/JbkmYtPJqmOPMcW
MSE9TNZz3el89K4fUNTEA0Ooq43zVdEEB4PxsE+g0jVOgBKYumIUYefeCVOb
SeyAyc00Fv5nUCyOXfCNLggf4jmXUMF8La0mew0EmxyiI8FZSYJw3vpaHTys
oCJz1ERmFzI//8Vg9gwA/m6VkfaxOQNBczGmBQkB6NAcPtIZ7sNzX4zxPNIK
2DKbHvEMVNTZ60bFz8LLWXaMgYqOSE+LDZO41GJjsevZBLChEVrGbOyzk+Ka
3me8Ee14wMXLDS8iFBdYOiJc41E0AkukJbIKndhSP0vCPZ+KvugPERLQpYmg
Yzn2y0ycocQ0G2faPYq4D1wJBVKhLrQbCrSdQha94yu1GUz+7QsbKoJNdlYC
VshAY/zkqUdiiRRGwso9INmNq1FE8KWeYT5Z2tLazfIDaqNeWFRi/L20CKSX
RdrcYQ6kWAdnHLjurhQ+9/HukA6Z/jgXgitD0i4TDuxpltnStg7hOn5ibxZA
u0LNFCNqu2M/TneL/ahgAEeA8l51DE4pqKKahXnGKctroIccr3x1wN0/R51e
gMReVD+kOejyX1BG2m2g25ORM1T7ZbYyvIkNXHvDG4u5FnZHSXOflllZWdxe
rZhqBIux1lepoVmZKB4BZfeVkbJtKYpYLZOplCqqQ5H3JU9SiETpajL+a4vl
SKd7L526HqjDi493RKKNyqiK+a8/Ohl3tuoJRCe+9LiXkEXrm48bHSQti/S4
nurDDnM0QNnj8fUMMTP73jYnt4VDhCZ9mtLXp/u/vcPR0nUHpYzdlDdhSpMD
bq2PM5tJvITGtEFZaaALjYNNDtZc3qBr1icY57DHrIDYR831Rt9uCX1DEyhT
fY2qLZ3t1jNBUQNYV/MrNORGw0r2xvqW6QwDOV5LxuJ3AEJEYnxFCPkVyboj
MEFPehYXSOZU35mw20LJ8YMDc8T6R17qzbpfpA6J609njQIdfHkNuXM6tNXm
K6X3+jUnyFtUFCL+8ynC3vT70l3Zgu737YQPdrQ7zS2oNat2Fm3EC48ABSrU
/Yu5uIVRhB0C0qYF6ACQhPdGkTLBa5iNZ3xj+hQFG/bC6JB0PcC5feoE8rFV
eHDqEbyPvBzqyV/3BrxlZvM+W2RRjVLO/kpx4AZNvO+v4CIRXQF1LZwlKYLP
5vFqKXRCo72dmNM2cH34L8bH0wtrNc8aCwvBWbiAbuIcomPIlOG7t5RNfkas
3xcN5PbWKuztjAuYKVs+OG41gHUz8kWQ45FL3Mqawof0Mlh3O5HfbOdTyG2M
5VdIsU7FmqntA4LzvrTj+F0um2eSIiSR7nVzJxI3vItmLHEHTOxeBHVN7gMn
L8Ah7nEQSK5Hxi+NDA/M5SOBRbINWS9mlqcwrxEHGhoerkW91ni6WOMrM5HQ
SmfwGtAGQVlKtzmgLSO+mm44feBb/JqNXIqWDifm3tiFULLy6zGo/Rh8/M6/
9UWwQkjow1P8jXEbu7fM3dpyxaaxn+fnRZqUePSYDwwp7UBuBHA9CY4/yVhq
EqJ/RWlcx74BtWoPceAdEK35q/rlnoaaxaj+wmEp+kn2iMMxCEQZ3JvQaBtf
1++30EswPsddAxab7qaL4WDPpARL9TjHXZXoZeqJz4SutoXLArTkBkz2T/sl
UsipLm3IiKfbWvr5TlpeDxQdCpr7kWcuT0XFn3zOAMGJ+G52MCogKJHJhcAl
qzciwZ7A7vKA6QzFs9cNqVBGYW5DVDhv2m3F6vpQhf10a6V/j9Jn6Zo4M6/p
Q6PGyS8K5bdr7FeZO4WixQ2Xsmc4EhvWnqvcY8lgX0/g56IMnm48Vekqr8Uq
I9x4W4wO9MBoBqg7wpb4v9yixa830WgsrJLZPGQcg6lVwSay1sVNukcI4vta
v1wGZTEJiIhZEP2CjFQVQbqQ0grfzlp8rO6OQQ5inRXVknZorndCw2YGxKak
qZPAtLlhOeRksxmA80MZMM+Bvn3K7WtA040z2l3XGB78aYw25mV8Z6SEAQTz
JR9aNWQDyEOmfAxOhD9nEVjAnU5fvXL2wbtkRXleoLpxopuyf/PB0JWIds+C
bmfG4/lAVVgKHXq6InHLq/E+rSA6G+qySRmI+HWG9S0Jii3wSFGa79TuANRU
qsB+vZsfAi9QNz2H5AbB7OKz7vjvXJhn2Dr9qWRfXo/Ij5XKnhAHweXVI106
CIyONYLc+3srTdq1NTaVxL4HMBbNmY6178k0ip3+5T/gVgCPIk0Z2aNq/EQE
j9bht02EKVNPT++2NIcRP/suS8zSlq8aI0lqGhU6dNfnMkEy9RJaMTn0yRU9
5Y3RnK58/2DHp4MkzykyCCfiY+o5sOleWpO7mxjj+Xof+jaEq4u+xyiXwWkI
9dEUqYr7WoDJylZE/xzs33u4hrWRpvkWmCCNllAtQkNFTw2dkY+459Qbp/N8
NMU6i5agMpYCV9y7fUSezIJIO8OobgEGpy5V+87CVRMIGFoy8ixCfJaDSJVr
2dcbbmdBFpVfm+VASgzB4l97fH3qlrsZoGFSdup2//lJYtAaZ9ucK4uuqUuu
Wi9lsTiPJwb7YMjMnmWr8ABNz5o7/8XBtQb3odFxAPgKT1mc+ZLAinLwjdYU
SmFTh1fzYzPcyUXUjoUCeO3rXDSJ+juTvN/tqhK4txZvz8n+vzHImNUO+ZXv
WmjWClHPFkeZxwV8GhPO6WXjX60yVEWM7+wUe/shiu7D7WX/wKmA7u7aEMoK
bpvkbZ0Jl5Tv4T9riffe5SJab+8RsSxOHTd/JtKW6oIGEY5AslNXXlFwhpmA
+s86cwdiuVYAGjRsJp8PuuXDOvi7iSMXM4OB52W9WYRXw0MK59aEHBaP5Hlb
xw4hLPAHaTX26Pe06DTfRyrZxDr3hOoYDPI2ENVlY13UPOAustaFQazzI89d
HsnHJwCOFRTcPhfDkFbakhJAjr0D+kxhsxYoAx7Qi7nJatDdC4lhcJHnFhds
skSn6KGEzZuPjbg3JFxuyZNs4NGdZ+sRVKWcouP5vUWr8SZT+yBdWdNHqfQI
kY9FJUSMj/6EdYblswfX1HtNnE0K7ISDAKQ6UJ/cWFYtO39pWgsG6WpMNo+R
Is40k0+6x9b526ZyBz60PqY3ENbRg+hbo2FA1p43Wx3ekunekKt0DGx/EOXW
mQiLu88LFLHmZvj6LIb8cDjQ8XWmQqPS81a52WOjqAERu+nCi7T1Dyp4eSyz
uK6tu9J8QL9Q07NmTOi3rXruKsQjUxhsCU+1eXw1JJKKCYof0iOEbPyiCmr3
FQVxkGLxqELud810bjNheJacjYFTyMkpv8RZoSr1b22ejWanzKRAvgFkEs5i
wPcF+Y7o3jNl1jGc3JS5dYqFBznbt+sSpowOAzBkOXCCkVhaCHfqefYUrVsF
vFJ7qWJVIRD3LML3DF5jICthMO7/rWBI/VG4bBBZYmFJbKnaL6oIh7jrnbNv
D+qAPjNlHsUFtDpeJVPXwSr/9Dy9Ng0UzAnS5RpeLaTsRJx2OydEKKcfBC5C
1nd0i6bPp3ShPqb0fgqmLwCX/W5HNVeTF1a3RpdBdjGNHUW/h6UsvG7ONIGd
OOKoy0N9nGKkY60JlfLWUbv9KU1gjNqnP1w7HD4b6Vw377cadP+V+hTN91NH
QlANrPK+h+t19yTrcFpMFSNni+E7nOKFYUZU2Gb8zpoubtbp36imb6pTV6YS
1L+2PamGZs42LZ0u7faPnYaeYyUULZvF3RoORMcLvgH11OfDAsKCVd/ZQba6
10Px2UcHcjDHtAdVs27Jg3b9LLUuUQmbRwRIiegdWrxAAOK1wQ3/Y1AIHfd7
aGd2lgIiENyQezHWTWowDyzCoxSh4ALj3O6Ot7i+wOtCU7udAglnQiKCX6uZ
ILHRlrq5hgCZbTKKoHpQcQAkWkL4Pk2vrHY3k/DaSwBuEXjI4rAOXdBVahlN
Ue7dFRSCdr3p0sgryUhY6NWt8GVqLPI+vax5TzD4+D7RCswNjLhANceFX+Dz
1OUZay+xoGqlYfZ1EC5gFULcMkeUwzMtPKSpUiyfqPBZqfiD3Ptj50oiBy6f
fitXDT2XSwzfPkwon0ukWENWLVYKl6DIXZFS0IduJcGo/Qm7Wipc9tmVNtm8
FO/e4tSUzY7pdqlcQOp1rl5/2ktHCH+rRgsiZYOpUOW4pAOKXrSn9OJ2GopW
m0CuhthXrppNqKivzXk++G5iWNSITv5Y+0OahdqyQWHED7gconk8QGxeEGAf
yDgbiCHXkUGuhwAzw0Rqm+62J4sDykmu77KdghUJarGgp5+MvMUUxTIMsvo6
2OZoNI4PIJ0LAdi3Kl8t1Gv6mfACpONSobMXAXS3d89DxP//df13G9UP9zGk
OrdqMncXH1dbCpUe4W9F3yTTu7MaDJ4e/KtwFcRe4B67j/aieFi002qZfmg6
DhWXtN9k0qBMdO1CfJ+YPUrj+XpK5Rg2soxoTJx+tPwdD9C2V0qLWAIGNBuH
Oxg6y57tz90LhBPeAN3KbG2zkIGNZjVBykgX4OVkJyx8rX1OMy+yPzSWrj/S
6xZMyv71yJTFEK1UBB6coSRmkrIzGchgJCyPDmDbFrrw8vVqYiXeMBP7XVlP
uvqlQYrKF9icbbqaefIoCRDWhkR5T/k1kOY+Jh59IILkzi2RA1rygvsUkQIq
nILJkCccgLHxlSyMAhv6rogezZcRcGzoc/hz+PrKtUEkkNKNhCeFd4OzXjEL
0ws1CLEhjQBsTxZP5iVuuZQN7ydwgeys+ViKIuAMVDyIeGs7+YiUA9HaCwpe
xeCzUmULi4YEmjieUUcVcLCHjfNxvhe0zoiwl3BuVmqZZ4hHgL1YP6VqLQbO
IKw8fdjO+RQozYwhocFdNdSghEDyz+DB4HJHjWRpuZL6y9hWVl3EylMlxsh9
TOsHQpyaPadRH4ucEhPWE6cddg75BN3keR/RqHpDmChPDqw72BCb9sSMrDw3
s4NDRUSfu/LvGxFiQuC0rymOVj0KMustS976VwXp4wwHdgP/uY6DGXzqWAH0
tyst7vchuYZs4nBJqZbwX7j4I9+WuRzcHC03jqGCPc4J9PBK96dOBMXIQqqg
HW5ApOOX+ZxcxZaus09SryCho+BkEu1Z3X089VqLyBGgGvKezehs6ZZBcL4c
NGVvmjnW59IFIUPPSubpeXi10HE/ry9kMM4c8JI1ra13TPvjDrLPZ5YMcxrG
fzFIkRE4q+i8WKJi7BoK7gxa1gmMCVT3+bdiqsM7NSSOxXEyhE5wxW2wxC3r
LURjrxJNFWK4TC/NW1pDYdEGHEyIO2XehGry5ytXuq3SdYQk6ja9SILQ/bsw
vGD3wE78LdbRdQ/KiKlvlBSpusscuvPnhkdu8ua9nuyk3vOEdMlWIrk9ZWvP
edDRujYuiypoAbIlg0Eluiw0hx44bXdQVtidZDCYAPDeT+b6uKI9WZZw/n9T
PW5Kd7KVYaxUXeEEXUY/2NtqgFdbwKqrE0/mxJIMwvw0V4BKTcIgcbQZB8c+
CITzTQviZ8UULTJzeCJEYKLTVZt1olSpQ2e7yeMV4hw0MVtAVtwk7dCbJPHU
HqIMRjVNTsEoPDgTGs2dFvBq9iXO0dyyez2VZjJeEY1VJ/2Bwg0CBedX5Cm2
awoDQdOGdnEAoiH7hpHC7lrWuIyBNFdvI0wjdB2qCU6R28jsBOzdXk4ei4Vi
IdbiIQIOkvXETfUD0UTtrjWCWYeHC7KXOyP+XMy1+uMojDJLPU01T50KkrHf
+CVhdra3oM5R36mNWWjwkhdY43wH7Mr0TYgwoEuK61V8QAFA8g5XD54t9+X1
zIMwcZInHh49T4xc8yjHw5ruqNMxsFGkVpZbn6uwuHKWXHrnfGRufMm+Bp8b
fHu4aMvipl4KxT8Kre+yy3o0WTBt0YifjJxUDAOnHhU4HWdJX61EA87QU9zM
ju/U84qWzdVRm+pS4WT9WjuAMtR4DcoGYNTiqcdKkELQ/4/oX8VUVK5gFORi
0vT6vpxw0v4Rkf47l9GvIqfPX9YbDSLYMXsUm4kWKTLWIu5EYNnVqmXO2SQ+
wyQp3StFiXBCK/1KYVb1yzhtmnm37dp1XnjuwhSIKjuzjLQf7uCX7k7TzofC
OEH3+WhUyhjGYR/GTQLYhUdv/8KFbl37TxAHXAnEUk/NeYhCC7h0DxIbj+0w
ZjvdanEb7w9Q9r+ipKEdWjWzlqJAhiY8pT4HCEJ2oK0PP4d5PDiT2h7UsuZh
FExqpmhPlSwiU6hrW91ysMpj2FHpf2Gqr922wNOs+yPSpvyXq3MC8KgIY0u0
FbHUBogjBmKnHBJ9nCcyoPKDoLKpGRshTVIZ4wp1djJXc+IMIXVYc2ZT0Dzu
2ag8KGp985KUar0BRNWkaP45MGp6B8XrLk2P4qEqX1OcnGvCMpXMVeD5Qf4M
xWcpicqIFRbp1u6MkdBPHgOToWvyZRzly7d8/c8pUScLbxE2N8gaIEC0DCjD
yhHyuJjrPBFGsmRDiGYU6YS5yjlCTXxbVkQci9XtBamMehg0mtLl2O5EePPK
KOK5+Hjzh8nRh49F0xgEwY2S04XgeUl9hU0+bYWtyIkGMQQTWRL6cp0zJ2RU
iNzb3DYIdYxDpr6g7oUV0/iDBlRucip1mAgSdh0kXRKta1vpMUBOPGm9iFov
1Sge4pF4mrMqMAdVZG1HW1T/w8j+3X8jHSc/YeJnqd4XmyUYY477ZzB/kQw6
qzGsc7aOjdN+4NcBhpiEpMaoVS8C2JwV5lXiyuOBsYpk5v+yeUqbwL/512Rs
Jzfye7GlbBEcLO2pRc8vh0fyhbQnFSTs7LcuMX8xJ6BjKMtAVCXoV0SdYGN3
u0UvnHYFcYrJRg/RE1iQkLY4t/TsB/CbdiGNgOkSeX/8JZ+cpZBhuo+byee/
AYC8jjShXmZ09ImGG6wWGF/yha7F8HmmH1sgY17ZLhikdo9ZRQTrYlWy5Tqe
HISbc7nxTMj1Sx2oMH1sK+PwafhtHD+wfiPKey0jtwg0iaepyfDh5rONn0Ew
xUwJX4stqubin8eBPXWerQ0XZaeF4W9TQ7lap+5QepMUz4cazOdClBog8GaK
Eu/H7ouPDPKmvrWbsw99jF1otWzd++7K4sFxq4n5n/EpdLvfL48TuBJbdDoW
J4YjA9THO37EjLEGSTw1M2jwyHyaRtihNvVFYXvg+2SXuLyyQryKjQhl8ueM
+7WjqQB6Q1AyN7QCzO2BjtpkfR+jp92C3xGEZ+OeBJS9nbsKpUmVtYEh74qv
iRh1NMiShgVYXo4H5MY1dQIPwOZGyELaeCMys6T6+vFuiv3NFcimVCZVWEXN
BxotMX3mTC8CqrpBkPFUGnQFT+NTVGC1D0Av0TKPo68IlELDbkFvhVVlnCB6
v25m8ZMOXM/OwZuRe4SxcGlzZ8ISiOXMJbZaOmMe23fTt+jPI2H1e51L7mXs
CEPF14FPRU0X1NohcTQe+DURIL1ShXg7f4rR3vVnDIXRDWQElEQ3Rg2IiYQJ
Qxp89DglTuv4vlvShIZjWl9kWSpmUhk04P8ZtvL5yIjDwPAfu8EuOZxktkcA
xqmfz70oRDPnfodDtfVJvDmZWyqmJLHQ1ErjoCFw4217NOZ0R1BLLBSMBmD/
EO+Xmm6vyS0qSv7XSTFtdlalZl880J1xIRHtZvYzJ7+pcMqWzrVKvPNITnxb
xxsW3nDgRsQJs8mgmFsHceFeaHrDpMCCJVAg5d1INQvxpS7whg3XA/umdlON
zy7SIdSezDgtHKHzSlr91Wzz1h93xT7sNtIp/ftxS567bCAu7qV2Yak3/GyD
WrYQ708cZklXPwBTT6MMfOlbMiOXt457eshq1jz8HnulDfWxnhDQKndn5h10
CKorS3UQvO0+wbkRW3p6CDLXiX7HrABoEJ+Z2Tluozh2eaFzAcWqhl5Zd+P+
NiBQmr1HJmBssri5g5ZdV0x0UHZ1s3aR4L2yTP10zE0K6ZlGCr7DUyHkQDoQ
6RnPW7PY2lJ+c7IX7/Y8d/hsLm4YntdhQg1BPE9ER2B9p967PdOkTAvDy1/B
oKMd6zwwJ4FcfD8QlsUv3isBQ6xPVRnWJrMPzaMAxtbInmPtHUZVqZPPXGEb
0BTSpUZhjFKp58Z25afNNHIo9h8X27ryhkDYpRKn7rHuVXou+RvBMDD4H3An
/JfmuuT3RUS6Nr4kgjsfIFMrjNraJqalFdPiRK5g79yEVN0XRLe3x6TMlife
c28SllsCT39J0yQ/YfHvFT6pm0MvfkxPg2nAbPTFFdA9tah0YZEOGpGzCDKv
bVMuntrfJDFtB5fJnvMQ4PYB6m3ycOuiQ6FMKSPgLJBMHHRzistNzaZBvjYt
NJk6oFv8bzlQwFUJhWfVKQo3lvTZzXnhBYrFFTt3Sfpj45Tl0cqVnAWlMX+7
6t/nDSzw8CmKCl1ExB8teuQeDfSDZ7GCN1UR0jUVUU/RwQtgX7KHzFyhIDxw
6f1mK4pT3StTF8H2QMiUHMcqTuwR9A5rIOiCm1UTwW7Ew7ZVrotTG+WsWdZL
nNLQUtuRJAykJzzk+aiul82KuH/mMlYY2aXLVvIrdb+kd67wbVcyaMqmLCsz
oDGwXM5NqM02z6B8sNfaOUESOJ22Of9no8LN+UKnWvtarrPvfB3ffj2xkV30
aPsh5X8FhHfOYGNzNeBSR7xdEdWuWNYP/uLZeUaCzCTKOtZWmTEJJrzN9xL/
QiCkTkbcG575afa+0ekGOS8Hqh+Da5mDowsiHkabadftkjM7GmzPuUsGxxzT
8O/Ban5NtDduBeWe/WLKKRsst2ZL9+ko6uFKYnZuf9b3f0bMI3cWhBbKCke5
h524wK8k+xw4J7Y8pnc/x44cdLUF1QQf4T43xKHasgDGRLv9bV6sufDXFS8s
R5coU6pMz6Yian51OC3PHXO7X+WO5MafD7rqSwAn60gxR2EmR1u7YlQDhRV+
jKr19XqDIqAI2mRdb1nAqJji4KXyLnUbY+C4tVfgYvFTmQAKUyt5WbQ2CLnu
J/j18t+i55YGaXvZGQ1Gccr5l+dS1ni5xooS0V3s8cPwbHtE7zi5ZPTzUOAU
D2/nWWq4VgFPYft7Bh8S17Z4gxRgM6FybmWzh0x6+Qf1Pw6dVVNiidLxaH/0
DbK5to8hvwcjvy1rC+dXtL3cdEkz5QriCCPhEoWt08tynJAKaqUT402xscR/
l4x0xQq2Z4sJ7/CpcEwcvvBu7MKoPG944r9GclA75+yn/WWDmZ6vIe4IN52v
CJs8PsTzjEvnJbrGt2nSNAPLvYvWzgOXxfji9n8gKi3axCEePUrS20cFD3CR
PRvx6zLBAlz75H8VXZxzM6Okx8SBVwtBJ4hHiHCC/4cynZwSypLjEwQdDn48
gqjYfurE4+MlKsRbhLgkcaBbVPMf/39W5UQmu6aFZdMt1c0A2nj64wX/D4K0
bU0lOZS+AEKdEUUf+4ozsQKo70sCVNBiKxfpgJRHli0ahV9GFCDGtSLc9pts
dEAFQBdp0VUO+dgKUwpNL32etmRiuWddkizgt0gjt7tDJ95+ULUw/EAZWm8J
KzclKU6nk2NJAvnnvVCeDSgtEaSf9VdqMUzzmyUUMZoGJh9OvqWtDZPeuk04
KEa6eVXcjtfE54L6BqerNscScjY+gWTktWa3W5HCrXdRpJ9x5voK570oOQw4
H4Ggg/YuD2DuSWQm7eyVWw0MCACBSpxam5TaDzgC9blR2HLPbnfUBTf/RJz/
qVc/fAfgxfD1IaleIVszCUZBUjk6NH6ZyOLDVwA6L2WBzIS/wKJalNd77n6n
iA9iUNc2H7V+U9miIZAJm25cwUm2LQOwxrkjuAT8TJTqIPHGPM9JuX67Cp+Y
JoJHFyvV4etkWKrZSYn43hQydPsTM8DZhpk8Yme/D5QkFCs3cYcPG0eOStlC
lfa/x159GFaf2oG9u30br6eHPpLSP2ttcC2DDd+aYukRdupIuSqBrSoVsUFH
o/l3pbwYkzkgWjeYV+nvzzlJmpdN48GirP/RGh8qd1+yEjYZzpUqxR3ltUZF
Tjb+q+2J39cnLsKPFourYtTQuvW9YcFl/p3luDetX1b28+lW89DKbi3WcKaP
MWQdgX6gW+53NBs41E1/oH7VVqoY+n8qa93NkRlr6BwSxeI6xuekMtfVXxwl
Q6CMXF29xD8gOCTWR/wtgIRv3ysbUYBasIv5NJx/I3NqDuRMsu0xzfXfwDFx
n2N4tBlOxXRBKyhHsmdJvMTUOjvXpJkM3HtPTIDvRCur4Xz727k7yEqstxOU
y1GOcWWQrxeBAuCLKWTQbbxLTkFKWmCqzczD+1UOFSt5usbEPNn4G74hQ/nN
kV2R1u1a/qDipMIKmxe6+v2oafhuTBBODKCciEzVsmg59mrNXlPcxNgZw/8k
KaB36btJQ1TBoxI1jZuF0YOUSR1kIO4/r2ZKTAnlrnR8hiaM/SPfMiBwUK+o
SWmtHciOcErDGAJm313Nklao0iA4As1qkl2FRtGN/ZrrRDYFUZtCcOMjxlPT
iLi2gUoQXVdFN6PkSAFqugCWfhjcuL7yic6IHbvRvFnz4HWEH81N3oWBnxYv
IWGZlEVtYd7LLcQx2P8Q5gM5huZ0w+rvxAEcdX9hArlynZ3n/SQCZe/jbo9X
FUJRY2riGwcuuEGPvFPsFf91lk/4BC81OQU3m5MXL2vemMQj8Fhz5ERQOLac
+XSLiR6ZTfbnHYN4JNrhNXfQ/r2ShjW7Dyjic9NDRZ9cpTzweGy3mHt6i74H
kYxGQ6S+SMkX4ZoWBsEKAfAhjyAvVjkpsMrpUCZOxT1GYYe06b6ITrM+XoMG
N7f9eyaXWG6MJ4nsFRyIiv79j5ovPrBeBbRVweLnV/42XY6EdswWQC1PTQbi
O4fmpVcxE9ABW4fr+RktXhXNOGp+9qGpyxjq37zOrPxUkZB/qLP4zpHln9Mo
nlXO/f4IlWsnDTCKgSGi6F3ZMJ+qY/97Ozq4twBDAStFBSccjh04rW3bgjLu
ynKlRJbwnMvgJP6HwuF5qH4lGhwxJK/IKCbD8t1ynryJCOCa39rhZzGBTH7E
Ko28cg1WoVzKq98qwyUL6rLd/QCNlZmRMqNbMDlzLs/UY1OQ3WYqrRgJIDJP
hOAzq8SRcMPQV/9Fj/cH+pFeUcGOxsmV8fwc2mWmEtD7KNPePtmB/zKd18tw
bwNJXDkcs8HinoI5j4+rQjBmOQKd3H6tTBTX0lg33nHD38Wk5JCpQUi0/r7i
IflWpxaq0/roLPtce3kETsTplVtvGVz8eC26rFuNp7nxXh+l7XSOs6/UZXaj
pqZnms4uzQe2Axm/jZFkA6rYavpZ/juEWOsxQFISxO+yE7vjy5lgSVOsSdsF
GS9z3WmxbfxbvVnkze6f+kN/fROAzC+MXoqLTmWanAJ1v/6gJ8QV01JzJAZW
a8Xk2TbKnKCO3yWKWZKDABRPPfHIo5pG0Fs6VK6ko+ByN1VAFDr7BQ/Bh2IJ
uunXWyvV6wue9gfrVixBSo8v7n+fLpRTLAI1YbhxvR/YZTjy7yMQs6hhE75+
BPprxCG35yeqAl+madn/zTqPoMf+jokK/ZQp2FNWiLkbkkieCziiP0+X1aRm
9D24djwrqrtfH3/Ww3m5kEc8OHrmwl85eaWiwGlFS+ZsxzX4GgWKF2JGiS35
oSIv3wpgEVkOcn+OXa+y9FQS4fN2w+BAy2DmbxRn0G0gnvjIvfSFkcVu8+Yq
eXZCuuybv+d9/lHF0CLJLlGrz5mrJusry9G2jw7mQwHJQnPRMcUmufBsdVfO
hPFHcFdzFyOnHIMvvb+/KPzxdcGRDacObIZM8o6jvjAAHfLqJg5oV2xxvMkA
jsNxVaWtmczp/8uof35GVZgbHlprUrTqUFr9QrzPuz5+LQwYcFMfuoL9blHT
p/hlbHgPau8ha8crqOoQH1HlWBg4OLszYwjYR/Pfcx4bb0LNLjU8jVgKpde0
W0g+okzqQnEvq5yOqZdWjZt8x912nmAo60PbK+NiPMkkxNwzIbwMjOMeXz8D
0HweQfGkDYfsmx52nCHQ4NYQu6HStiXfBveLng+PscpNdgfk3szz1CS0n/7B
wBpBHHXmbvJiNm3TTWId8s5iPu96406SBI16eRMSH4F65HA0IBNdO29g3vni
QOpnkBv6VdXKiz4x8J5B3ibs96o/RjTO20afHBCG5efYL5iau1dgx1pM3mWO
mkXBU9ksl0r57F5467dQLk7l0CErsWjSFmXKglf02D6CkbKCk5go2Eaton5r
/kgXkOxn2/5+o7/sVwNnQLy37/a673j6KS+/CI2cRFO/lbs4F79PW1NNS+mP
SuFJ/uw71zz58viOmotAlFl/VMOuafwzmqe7/1/Smty3r9lCcgtT1fDJW6W9
89ZO2sRiP6Kx9LVL+glIGwSw0ph1WwvnvkNr4KMezTyR4ysy+NrIPkRRWNEM
bNyqiGVw5lxhUPkodPiseH68npKjABa+6uqCqnLHiLqz4/+hs8PluJVFnH7r
6+ZFln+242a2t0xgd/IENdptbZy+vGc85louZ3aqEoLauvYV9RSEk2cF73bi
5om/pjlqkQ3rRlQ7ohAa4TByYnLDCA9dCdJzNXvNPf+B5hWl7Ak+T0XDf+5F
Q8eWjQlWJTIjoMIqtXeW5VW7X1Kb2Kg44axDO5/nLHib1LGCy5SapgytMqBb
EdJhtzU4MD5ToAoLpse9OKMoObt825x3abuKIh2tk3DynFxdhb3zzpdMeNmy
IpukCWbvTXKJVVf40XGMZwDP5kgrLib+u5TkbZNjVBxjhtZI1SyD3YY2/ExR
tAMAC7ePdP0V1zt4lkA+s6h7vGHwtzLtEoyHBKUDnlQvhLm9DB5QjWBWSzcG
RPyzkF+Z2H6h6jKQtK/28zSoeSHUjqHOGNcmgh0PitX5OKyLo4B4q5qJQnAL
DBH/MJ4pI+ayMopXZnkDeTyTTZrQ5I2N2yDMQkrzEKnGvIZWl547LZ4Bz7Ib
wdxZcS/tya9ieiihWnFFQmqlm9+yw4eWGj2Fpb4gAxiBqJDZ0ef1zq1/L9Oh
oa++gctK4mLbCJN0FgncjiLgy3kW8VuMffsC4l2TE19RJrFDcDZwWU7Hn0Ff
ldqVNBIDEIZBro19jek3eyHdvNVIwTUIl3F6XmHTsTA1p1v7pNNFF/nvZkPr
GCFzXD077W/8WHrwIuNGq/W/wvv+knE/oco6sBU4BsKPjcyDwYlN1NoTYCbq
Tin9KhST/ctTy3q+N9lN/JFeWL6lSuUWlKimO0LPS0eiYMGUW3d/6UfoQYkY
m6gxkVRKa9eC8/89buwWKjR+JUZd34tnrWyGqqzoGHFFfglklWoAuwYQjm4X
/hoYs6HlGp60/O67TwAGAV4V2CGZr/0HTVgT5CpWqtDLxrH7Gn6sJZGhNvrS
M5pNvEuBLGs=

`pragma protect end_protected
