// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
VLMtkFrIUoKkeIOqNNxk7P/CxxXMwRlEI+ln73epgouUfx4oFEo2BHwhj2dM
N7MOG5ilExUDEn/337i+qzq5g5nd95ys3/TGZO20ERmtDxKpny4qnpcllgYG
ZtkDL+Yi+D+PTfOzTWPe/jCmf5m5LH8ssKiVgVUMGvtL5SXV8Ya9vr/bb3ky
DmQb1t87wswWo5DiqouknuWGD1gPowLhxfHmLRHE6DfJuPYwq3eqpc1Bq9Zy
ctwrF6XqtwgIaj+RpqtwfWMYNJqVkR9OtnnW8MXb93GVOmlWS/EzzZEOsQQ2
0k/09eOmq8uJjt3mZimm9QioMHMI7vly7fL+c+MWFA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
fjUgsHqP7ModHcodCRX5PEa/0i/3d27Z5DYceWzbOz5YVqSLYyGrwXBWFeRV
XlXvD0tVyUiFtVNYii8vx15wLRqUK/vwUz2nbN8m4qlS0LJnEdWT0/O8hVhw
RAfi0NE9NZIV7ABVl96ajeIVtYRxFkWK511lO/7ure8g7DIs+h1zfW5xS0DW
jieJzABRWZcRErBHQAJ8Oo2RHnapsaxPI2mAGQdbHP5cNakGeTWKiUHDW8Ob
zA86QicZ/wXI2ZZXrxHcn5K+zq4MZkxmQfDHan8sHdewiwY561tmz4cL8a/z
kaCcyePVC1MEefjKk6/wOdoc6Yph43RLm1WXHs6+EQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
KsqHxl8OTJblnN/SXwgb/Q+AMm8KQpoj1SHW0W3BVS2KH4WDC/XhRZmB6qL3
dZdzmb2yXd4nvQtE+dGwmlQ8tyqb1FtEI+4WeCbWe8+Di5QrWI2DlscGADpH
1jKt67DRcVORSaO6Jduj/5+JMH7og3+AUXHy/RDy89gK5JOz4QqYn4mI+Etz
0SLDZ1tXj46lSkhFu9EFoA79aOB7EpiX9WywkSA2EhFQw6qGik+5bvVg+mIx
UE1/3gv1aOMKpdeuqWvQD+5EvZlKvYpYKKc0T5P3c51s8Ft/v8gfeuP1mF2y
q3VbuO1n3lZQdBNWXbhSOkvfYkzyYhgxNICc9AiEVA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
eeroYHGOvUY42vIcjOwVrp7lSGl3DXIO8MBxILa0PJRUworfo7RCivDH1Bwc
CcR5oUrmDM9RYTFSxsW6EG0lVjX57BaR9/u/WokKdjqI0sLX/pHys58zrG22
sTc+qkbgiccs3ORbG/ANFwuLXB/7LToQslgiCk61ynGtWRxa5oM=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
RyTHgaNNjY1NnHIXAxlo4STh07HTU6s8YPz9YQA7yfbLXP86GReSKx8dDjMQ
Nmv3X7PN8G6J9ddwWJxr4LvtGifAUOQARYaQnmxjNsb4GHasqOwVN+d9z9W+
4lyYgNMLhz/krUQYghj8atYkg9RHnJrBQFmdf73OFW0le11G628eq1u6Yamb
Fhloq1zFNJDR35xxuAoUdqzBaq3wbUZTBAiLGZ0jsKOOUvzMFGYDsbAZ+3oG
5t0o+cbQAz2CjXhI3vm9dD0EaXHMTAZyn8wpV+PrrRrrWzoqcIxWGtThcB1m
VeTHap+Tg4RT1ZRew6cvf/akINluzho/uDpXDO1tP/dn9gzxe+beqV9KzdxB
yfS5v+5gkK2rLGhMzNDksz8QAXQEbrezwPqiC3Slk83/1Ic/ySGy2W9R9uu/
aLNHppbReT4ySvNnBIF5t8o+0dP3uK/OF0deWpfP7BPYrD5Mwu6II30gqPTO
6dczXUoNHp92k1/yUDvOGCjAg2Stv7fY


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
A/iuvB/ivBnhbpUcb+Sa2Dl23DSI/dgbRh/UupWEZjNkt9eZv+phFASc2MqH
uv0da8wbpS61W6oQSMg1rnISVuzkFfy4rFaaRYIsMtlusqKkgu7lo0nWHVX9
PikbBYUeP89XkQJsJCE4pnN5AlLri64vP2y93wYrGiZVm9V5aYg=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
VoELoJcEy4/I/CyHGhHIlP7rhinCCnqRfskmR09aUPYYkn6qjdlfTbQCGIBs
70fij43TTqWmJhMkNcbkvxf9PcX03aIPk72bgAiRVNRbK8Dtupr6W6Xyje1p
ASG4Tm4Ry+7ckxFGde6uIM4edVlrCLOXHhZMxbygcpCNMGZTVtI=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 6096)
`pragma protect data_block
s0KE4/cWKoSBMcBXuCg2P6kYcUdcEh3S3FGOcoLH1HOqXtNuAVcFWgYGhLhs
bTYekrVDpC6v0oJEbf7IXra0cHpn+oITpKm4dGIn/D81rhUQQeyI7KRWjJTJ
PUTnI7PUYtR7kBjEiDjdmyaCUkf4YNuUQxWdAdaedSbjEZuox55UUJ+rdqP9
limc6Gem5cSafNwh89sY595O/eBQWnugpMJcYBWFKe+RmPj8pKQyRUint86F
BnNUFFr4Z5YFuIMb0NOuE5hF0oWi89ZLiEIdkqGtW3SHcCcQNMqqsA0qQOLl
K3GN3d+MFs6SFJY6UT655PH41Ie6bLwL7ktBZ+/KxvIxNpQxnCPRix8N7/Pr
xPEgN7IL2fcW+XVsiyJvAFa9mNKG3W85NlfaZIzjhmKg6YcabhqzNsmNJbEf
6c/u0TsFf5Ip///ddBwC/XuP0LAWo48RPwYA+cS28m/qqrh0hKUTmJBqxJDi
7MQvjP8vUC5nICyMBkni05HUMUfEepAjd0oYmsirWshJA+84ro9R3zHDXWxW
x12OvQZQIT9Br/D3DZbTb9+jCP23u6g4KJqoF5gHxmq6PLzG1/NY/pdWk/pM
hO9KxRWB1UA532dRdDNIqpCn2bpeq+00jT1PC/Acx+QwWKNzMTgV3SSFWfzs
SR4L29+sWYPIm/Pktc+KKbTiKH2KSKfA6JT/rSJVYrq/DUEPXT+plKLyz/iW
n056+LSGQFWIX1iwadjdRDaCSQWBI7la+nObD004Z7m2cFymO09ihvFILzEp
aIaKe2UE1sPnyGDrkzt1TVt3gbN2meN/j//wbX6imrZ0eoXYfBPs0KqxEuGH
2wj1pZgypPHxNW4pJIrWtxrAsAO/rUaIGPF9otADuXLFK34gYU9I/rpRNI2e
3QmxZUnxL35yPpCB3+33hbfFSvEBBwoF9r15zhsotPVF3DTaVnvvPu1WuF8d
s8pQXHNaIJ+lDjSr/dt50EcJ2OTdp7kmBDvNUDuILwl/AUTZ0XWoIBktGm/I
LBLQlfxWLCCRp+kA/LNa4BMhsr/hrhoF6ZH4AbUfWO1UvGVjvwqbOsSkYfoi
zW2tSum1Kt+G/m1wFri2gxwb0nkgcc3GACOn0GfuCWPEi+piTcIsE61C+IQa
NDqXrny31FUUltWW7BpAVfwyo9lftwnKrEdiZSAwhb3Pz0bD1dKNu3mwVcSj
eCPrNLbJAK8yCAVHDBhERyXeHufQrL5l092ilGxXZDI3Q4qmzP16AGbM95KE
CHpH9MrE8gVOgl0OrNIaxQ8S+DJmx0ORZp9+ayHuN7aznhHNLR8HStPXDeWF
ZVq+doi6AdnmozEVHSy2ZDpfY0ey+oMmpd5Rr3+5XSDDtkHLOKcI+G3e7GjN
yv88gCl2Ov2FYH9nxpZXdgXwMaLmBWxel3BflxISV84GHz3gihJGcxyo44vk
DSAH3Xk5EQgvfWn2ihkyI/U3t+Lep+FgXaTs2sfhnE7gNySRbcLhQ0tk2fbJ
J2w6HhRV4FJG/sGmdkBplCEiLufOyXkQWZ4PvW4A/jnKCkkGXT4fZGjb2x2h
rdsV38T/Zej/Diu742LyAthgQifj6vayR/maWw+lOCiaI+LeH6mmwyzfCx7z
uvw7FCgZSAX3cdfKWM8n7tBHXFfch6go+T76/HRlWhKhGNSDiwu68iGVI7RJ
vNtxz51JstqbGkH7DeUk+sxK6e2WX5chJT5uOs4O2oWabmj8YFr7Tb6C6jdM
njdkYWOfBjBaoV9xYfYD8VwoVUlwUaiHWi975jASOYpWboQj8jSF4grJJLwG
aYoUpzjmL2arQkO6q2SqJiHDziJEy4T66w6G0pAfNQkgSvSjgMi/ctMoFNUg
GhRdLaXDvgT+uGXTZh5oUx+SvlMFriC7UPZScioPf0sLVVprTHoNac42sWnx
AG1R41I/F46lAmK1a9DxQar8Hgb3T2UBmh1Kof2xQePUi7dzCjfe1rnaLkEo
f5/vhRD/L/uo58jMdbgjbiKaqm1y/igenqKKxEd2iZ8Cpkm6ALjvC9yi5UcR
HbQjE/dE/2NSHE7dixspZmESCIL0hnMjwqEWv0/vDeLQOiskd1Tqj3dDZqyt
EdXO6M2dVwSpk9WIenZrRqrO33ixOkVPuMgk3SlwGAe9eLyhMTeTB2cpX3pI
fswbUxXKVbUzthjOOPxhnR6wGfKwZN8Xvl2Oq9/YRBj8gE4w70U7HkyDUUeZ
YOFOtsyvjvNMSRWxEnsm+5DDa56KdY201HYdhrZ2yOa0qLY0juI9Vm8gFerN
b5Il/hY5YdcXP7mRe9AftHAw/7JiQFGQwfrhK/D9Yc5hTycRM5aihJS0XJmp
XT0uHwPiph1Zo5SkFRuV0+V9plw/D+hSfAaUBF5wsHHuAWveILnQWaOuxNXm
duqU4SQD1RVXr8M+ikVraZFdO+T0R43/aMJS0aRxtv9wo8fg7QYIzuYHjSGo
vJ0FtcuoYfFt4Si/fdkTy2GNOYZ0fubB+lCp5qyO6/gyDWe/dwWhuBQ3UX08
64bbJyywh3aSA1SE67UwSPVUU+S1TJuvUX3/XMMR30ipdUWPyC+2ku06nk/c
LPb37JhgzInvkG8SqxvXptjbg4JCKnSs4bbo7FmZfy16S40TxP0K2/NtrhLk
VyJnwrVvmQs1oZ8MPQkM9ESKmDqb7YccUGYsOrTqY66jdQSyciatFRlWZ/FC
Q+8BitLLyaUfoT76VEmR7lOpqG0nd3vtQM7m67HUKZ/zlyzjN2/ivnFf1K+1
KhGXRX4l3TMicvysstnuiXSxZ9GCqQ3GhPoz56M1SVNayAdlU0yg8yZExnvW
BfbXmvQcW+4qbSd56cXNzYUzyifoJ5aH1Khi+Se/DWTL5PHZegqswt3Xn+lA
S163mjXKJnQsUebGXUcaaWms2dMqivzlePkL2VRaaKYJmxQeFVfQGmqggxDS
tXMkSekhX2EJLySnXM27TmztcpfaSr0T+8zkqmspORthIKGOKvAkilCvs/Bd
WRrlJyXo9dXrqJe5d5cLFS9kVEp3DzzD51dLeQv42061ZrANHPleott1lOci
EB1gLjrjAE35KUJu10PBtSdstgIBtWOTJV9Zg1pjOR7Zewre15FhNnQ0EL4a
uoGj15pDcauP29qEhdRVJapjUiWi0hOVCB3GDbRFXpD3ydw95TCJO8cqlCEn
/AGDhVpbfLuhSJ+HshANFef9cOrx8xUo469B2IIDjfL89ZJ3IW2oEK8BmQRz
ihZGYDhPvLat7BZ6xOY6QyQLHP0xjOLmy7aLpjGHYjDd3xGiB7ifFtvN4Cdy
lqDibsEJ07iSK9RF6t9WzPNyUe+/lVC04oqxp0ail+QXfun5L6eLhS+W4Srw
AYs0s+IY62sc/lWrrac6MnWeNUlkvS2urwEx5HdYjqqLp0wHk7hWmae2N8gp
WEXqaMeAU43aX+gYkE/lYmhsunv6V9Fh826kC44MRPWOTuYEddkmokAY60Y4
v0xCPDNI0cvxkUIiK6tH0M/XmP05BVBZ7P+mYrG5uGIK43ZWCxsyIYb5Qbsv
1Bi3+JtQHZwRsVhPk1kf4R1sXswJa+7M0m4ycldm9QCU09T/DYwxymMmLpGf
zIQbbKeTKxraUJdLnhdeCCJ3CtGSYLEwRLOIjrTdb+TvgmWm67XjXwtFpKAG
EIinmxQBtn6u53UwiGJsIvE+MLZhXcaVDPz2orBaOWPa23XcprI3Aobs+xkg
h9p/W5qx4zoV8KuBjRKhL/p40otIoRWl5lOfGRnu29eM5paJoRWLvdiaIyBu
uBKZW0D8I7QAfUgq7eKeTB/en+GTQW67oSl2PhEt2CIlOCnRqDUZdXZyW2OG
e8lkHck/UnvVvX0pmfVI/VIC3tVrCOUPywIEjI+zPatyH9YdirSBuechxA2L
Mj9TjS/sabZ6Xu+/tnKbOI0dbKJTEls1UAedRYU9Q0rqfUJcMV8AXPsLghJn
39ui1gi5vcPIOtQFrH5zDtUvi3Xv/Qr/D6EuIHqmaD+5FGa5HXGh50PIWUdb
ct/Mo6H9QPD7fkeWu7MAOPV0H/lNVJ//QDTNnyMWLBAuoMwOMSXJ4XUI8eeN
dnSCAmXjj9JlsEFdSD8eODC2R5aDk2ctXtrDckxON/611LKKbWHddDFKLC4B
qmFMDG4IYyb3e1NOVR34lRD5vivnQbxcNauQxpxLX5ZnhLY8oV6DkuBmNEsZ
9FBWFqQ5+Ki9AF1s2m6GhcpNWuXS6QiO23rf7d8j3OOCyJPaFgM/w5cVZGwo
6OUOMqYGbjAx/1c5SAUZaMbYAkChbgsjypkPYmtd+5HIqXSoj/+2WesaPSR5
XfZGZPwbGN0RemBBrHIVgpmcmwGyMCFoOPwj1gdGEoBiX4YdaLYX36qqBEH1
ZwOTOu4EZA96j6bU6HN+PZgdV1MsZWXk4C/43F2XY4GaxNdNKZ5QRKabyctr
nOHOBm3JT3s9xAEFJguyTn/xgGRJW8BrukQe+dOSe94mmwfk96VlikOW0VJd
3+9tjblzvr4a+H6Kev/TKBPZJjbH3JEZhU83PDlCVG9GYrKY5DoYwO0Sohi/
QLPqMbMHX1ovx6biaaCAOZDh6Q3cXpIoSXNW2ip/PuC5RqCJ3I2Yy3utXe7G
OOvfdaRQHj6aQpcm/zdcyP8MXCGgUbSHMPLunH7vjKFn0LnE6WX87mxypHix
UwHKLpD+SFke9BTcJUkrqXLTZ8RQ3Tv1tGjmH8bzbX3ihsIoBiPEiiPnvsh5
rhj5tBsG2zHD3M7jmPbjlJpYpLeHfBZU132f88QZZ7rE1WxC70xVQYfiA1rb
5lHrvmT7DyfHwZJHB3DfFNxa2GEIfPmDXuUDvkgxMAJhgqMdxUt8WIltJiUk
8kowmkzQGHVgHCAg3xZtmWFiTKAERVrDEe0Jv7oDC4yKofwuzuWtVGPclIBB
Nmj1U3E5KV7ct7dPE9YAIdmQLPt3VbnIkJEEBqPwSEPFMjMqFTP6crpPMIB/
HNiAwZgCLKVKmCsFqtB+SB/s5oNKgitDoSl3COzLwwmbmCqvp+PPGc8w2C+U
j/sdiiM8zoougKshW0RBj8gcUcdvQH7OYKCerr0Xj9V/JYPyOcAMECyBvKnA
VQsiwJR5cTR9swZgW7gN/xP8xO0yP0oHTP/epn5ZuSs9t5dxIIAC+ScDrxKX
5mIl9riGEsZB3/sbs970VA58PkKrywIlQV379SS9W/FPGNDk2cNoZBLtrbc2
HT8RfkMHm6XxK9ivVLPE0dz+UnLt4THw70XTztLdvH3MVGX5i9jD/9lOydeV
DDDPSPr85NlGvFbKNz+3XMQIIQZa8/SrZq3Z8qaSHCXHaDPitN6lwUlSlDje
vuwlMPQ8LO8zUmqoB3uqvmDeSFVqzuvVeY0JTfwM4masukskWQeJq8gsC49Z
Ep2W70V9xdKdVuyCFz+02WY46E3XNGYljdSgH2XQXp26jgOnC6wjYuDPrejm
7YPIYezFKL9VZwxH14frOGwKwjl/zZhm0f3rcDPTn2FB+QjOItz52Pgctyfm
EkSSplTDk6WDJzPQIiMcVAgsJ6O/ak+q7p71ryRbSgG4om+1MJrk3seK7Trh
My/7SZ3kqCu5I2zmMmQny6+m9+MzwxUgGjWfEuZeIiGlQc6+eHToqzvq4d4K
XPvfPRmW91i8reI6vxYGO76uS8pJp+6QQ1l/uFGt7DEY01gE9Db8sncw2Hbo
bVdJ9BqygMZUozIjnfOu/OaxY/y88DLd436afzAdjTD+daxOtlqPfP5UmC3q
NBvaEYyrN4J9WKDz3nJM8KGqayaQnMy7Ti5cB2zgg6CDKhcimc7wXK8lF7Su
4PKz/RmGuEsSrBwG8/uq+DYunardek1woqe8etKnmE68AY4t0sJOVNgq7Lbo
g1hfONEbkG5gtyzZDxXSgdiqNi751BdtWYvZ3osr5Z41ox+0mx31th+N1I2i
Uuuwwm62sa0OGqqmmlcCDohITH+c9nKhB5s3YgvuK8dZbrDZxViG7AyZj7gu
5mNIMBL4BfdYcTMUjgU3nkgIa1FKpTIv3dZOmdbjYakuuObaKdTEOQtFDvrE
B/sIiGqpX6nSPNzFMqhxcr+HBgwkUFhM0cT9KqrSODOdqgFCLCEChs1Aupwr
GrzpOPKumRiGTHbUXTy4t+LW0dVA9ajchGI5XTXJj5Qlte/ZIRBx84UoAzYR
yBNHDs0QfF7weTJ5wub59WL8J2M6s5vDPn+Sk80fsQmUYr/VUd5AUd871r9D
SuRQQidvfJyJ5DqsTt2d306jY2fOPY38HxHR4Kp+rf9tt05AK9oObtS/EWqP
mh9cdUrsuYcOndVE3D9Q/G7vA7h6nLVma+TFhr4UGCr/YFUKOdFJalOkDyXO
cKyFBnhfk4eZOWHGQc0Esv12Z+uh0gSv5ro2RctkDRdNdJ4Yy2vz/RQlMTTj
fCmFAqJCgQgW8TRTjdZPdSyXzfNgSjEm+l17MpxulswPQ091X9c1qNeKHNL9
NU4WmHTMYv0mRgnNhgxaZwwzYjBa2e/mhGPxP8VDoSe2DUL818oSqAmM6Rz5
ZsYpNapUuRLDJr/YBefQUmSnA/sFnAig05CEtWFf7SkVMwZ4ijsmV7ZaMTEb
U0IaycVWHAxRxje4SJmD+V4RcoGHpFoSdoN0Xy0hxNyYrDY/Bh7zX9Q3pDZk
Mhl/gUSDioXNwvyOtIb3i4dg+sQM6MruxoRTRkVV/67pjmFST/81TV+JAS3G
xFDbjnw27M8xEyQh9xxoCNotZdCFzEVuZXWAIuhBU+VveUWrXXjK/8/7UOfN
+W3WSS6yYdXBx7IMM3BnOXW9r/34G8+vX1BK0WU6oy7VFnj8yn08Ihcbhyzl
w0lnhzDDRTkxplRRLpbRdS9EJKvr4Wmsxuu6uszuW9aQbSgMcVD1Fmm9Ie7J
H0Vf5WWaa74gQ557p7cLhljHo8xXD204lzshreRO3woDPeTZGDQ+6jQhS+QC
xa9W/oPKnhR3Co1u3NmIEeNu/taucbKOmzm78PgifazYi5s4FxRNuwvZ5V+j
rXdNiCgPLJ1/UzU1lWgMJVxGK8fNwYhbDj9dUbxM4cy6Sr1Bp79V+4YyPibL
04mMy5T3hglKbrOuVgwuJAp6t1cZvocBiu+DqDXI/7pnx7j3PG0L98627Hw2
X3pojZ+b8rAG6xNeu+ujE9h2cx4EbXBnXQeMYrs8z6n26N5VTSL1+CARgWsR
joZh5ovwqd76e8J8WmrFY6Qm3A7dGPuXLhKEJcsFoHYpOdw50nBcBB7TR/l/
mM3lF6lR3oCqcLPiKebvCX+O0pbJj0kTSwJpCjx4EH/ZaNhm9Uw75w0X+Bx8
vvGrMZFKx1hQjNdLxwdUUWF/DSGPSOiMaRabuP6nbGdVEiwO5lKnFjgeAURR
J3EH60BSYRhFTYeImtX7n9nTOcp39eELsqFKxBhS04wIfThH6AZlr3c4lXaf
Pk/AjElbp4ORELeCI0/3VXPOuVHDEh7fH/H0ty0LyI9ojtfZ7E5Wi7h8XgRm
WmE607b4UpGYECyDuFaPUEV+W9EmAlChvrdiHVA6jIx6jnRA8RPWLx5OD66c
64kPR3COf/j1YgIGkndT/SWhZijk9ETGJnIGzM1St6YWeaUY4ZJlW/SKrH3Q
ponT+PocvUf0oU3sBXzTuGc2d0jWjHsonGC/aCflmLXVauxdm1+wFPWu5XZX
IuxTUce+5P18KTsehV6N/iyJImubZWuRXbGkTdY4iKdCtnAopayzrzBoLXqa
sxtX/d2RlIl7KUnHjwU/nRQzNuBPXTuooC/vcdeiL55xxluPJFSGC4mqR+ZF
Q9u11vt4YTOUkyPoBaqfeXsK/GASaNAf8kk8Hpz0V+XcrSB8C+GLLFtKvA0z
mJb+qhtWJ7HDBnbfNwlaLtz1i5t4l0FFY8942NVZsokvPmnP8wIbcTGFd6DP
UXKr0V8kfwOhYWMS3wc0Dw++ifuK73v0uzHumDV4NxIJ9ZRaw92W8gDqL6fH
39QvXJJxRgBTNMEsgpwlsvlXM+fazj2lBges6mpKzjVOtzQ+qwkPhuqNeSZB
KimRhQ50Ao4HspCtE05T8xSLU6KlZyevubs8UWI5reIIu6FtN7vU+AsGdY5r
kpo8Jj5oi7uLk8HaxTzwuflmVIfq

`pragma protect end_protected
