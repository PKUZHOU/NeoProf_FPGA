// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
OOAzhb1Tcz3QoZ0pEHkxTUzK2eCqqGB/MFZFSGyK88yOP1wunZPct9yFxPcmo9JV
uo6bYu2FV5mFHtmvDhEGt13PTP9cviVS1nbhAxGs3PmnvQyg8PBYyypzPMyJWGgY
ndggk2vR/xnZrW3e3ZRLCTgcUYaN45cehfoE5LfjZ4E=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 2272 )
`pragma protect data_block
FeGl4tQbPuQ53QpLHZN7HC/2lNFxi38CZhZE/mTXZuC8WSEIdrPJYDAc1BcSb1BL
MRUdbIIK0AKnhBUwnsMD8OFZqwxqteobMmx56NLagF+9Cw41xnhmBv3vIeD5cQoT
QVGWsa3AABfed2wR0gOPjKnH9sa4M/+xd7rGRyGjkIgcJdBOfENiTGPQYhOu03/B
ed1N9WmDzn4tYZgZ7gBcxFddfINlanIybvcfyzs2qTrqlliPz0QYBbrua2ZTtZ/v
MWke5YFf2LZal5t2MVl0v8uiRMzhZA2WjqWYyprI45CKjppA+ijgD6pw9ckXI5c9
fX+jIyUfIMhsKDEbGdgcf08cxCIsvyRL/3cOFJ5Pr4dLpqT/AXqZdGDt7S+2+k1O
XFSGUDcBeTlAyaJBQekmOtyvR0zI0qDsP04dcE1kvRStn7ijxtwWKs6LAFWK207U
+PcYSY4OOotnTI3UnPcCMpazRXp5zw1jGOgKNn1NBdTGm4/ui/z3sVh8In6BAEsO
TZ2pMvmOu5nmPcUau5WiL4WmjYPX5GOKGZlhyY8nIT9e6zfPj5QyPDxgtx1sVyIl
WgP7xYJTJy0Hs9hq/2nOEBqEjAg3OQOHb4mnEUSNLmzL2258o52GpIzdAf9XiBLQ
Fxi6VlIoQgbdHABYZV9esOf5KH3LzuYRxRYBePNdfOcF5+e5iom9QGaf8LiAPI6m
eOuRSUhJk0JQLOl5MroKoIEjUJj+ozWry8GulBetWLKGJABLo+o7PPhbKkLrGJ3e
z4oqmCkrYReTQxouh8BQI/630y6lw8nbvREuQ0G09n0IWBz2WNGmeZUn1NMryZOB
Jh6OKMVqkpCkPEMld/aic5xO8qU7vUNevvAaELOJNF/XFDqz2zg5+TLqByoHB8/+
wULvQVtcvBVZehz2xCm6aSLYnb0uKi9KN2pOe7Kyfm1igZ7Iwu1vz4a/9nlZo/hA
AzrTPLwCw6sTtBnn/bdZ/EaQPIcBmWTszmA2ztGRx92xxtMcqRTCNRPtT9z/Hhiz
oYy4Hm/QvD3ZmU8bRey8mYfqlKbAzIQr6aU+ENeRciZ0z7Q7FlFuHn4JTygGoaKX
ZKtnZ0W1ZIASztjTaaSoemlFTGg0jNKgRRVMLixB99UIcpbmHKLMLtMAp5IP5xrp
wx0/Eo/LJsYHlXcXCJICF7ZKyukDrGeTajSqlNrnrVE8KR5fmF0dxHJ/JHmNqGPe
WjrJUznJCl9DDo7qXBxaiTQ1+2w1tOOePPhNmVJ854ZbnV1iFV44RHFByMrZIhpJ
D2rIaEroolPklwP+Mi8YLTft+BfMslpIBYd8Z456n708/hLRmqy3bzSKNdKbHJGa
8D5PeESaNOWCZZuumoLaAHNwmGATEMcr+0hHUvOogM8QOWiy4rGN8eFo4yNuFQAm
j1cqCNdazOro6TITFkkrqHrJmzQvduQMmC+KKNc2jov0iJkJ3XC1fjpSC1ymuKR3
s2nk/ffTYie/5jro0uudkH4weCF78OpwA60Elz7MYHXn2lgxtggCiktSeUpsgvBp
NlWGM5jocQeo/s6mM5OCpHJgIc+5WIRmUuTrG0iWkd7eDp4Sx083u82OTzEYb2qL
kRsMt5VA0HLUcOzCjo7cGbwLuoNbe5Xr4aBVW4Ij11sE+IL17mLutA1ikJzUQtiJ
pmeNgC1NmVH4c6rxvzG9Qw6DAF9dcHKVt2woxeKegJu8xX5bLeth/InrP6CSIZK2
G179D5aSPy2YoF5VXnuZgapyu7+uPtudinQX4vFwnjOgUAizwhY0wgmULuLiPHg+
Fj3Fcch0B5VUAyEkvluZdXqnz1LqxL817lfiVu9zbW/+HrMQ3fw2lHEcl112pAhe
JAaY/F/NBRmQtrGZ8qtybrXg0YzaVl+lIU+k3pCt3RgaSLzoAxlsZ4NxHPNz3E0/
ru8ZvhE1pWz9cl4C8xq+L3jdjiK/hbO6NZerzZzR0fuCvThVWzF0JNhd6Tr65i8Y
N2Lf80IYRjqRTccWlvJIft+JwMK4G2TbZoiJCSFXn50fXHJiuV9BwwB+Yky5sngG
+0mSaiNZhnygoORimdtQlcw+4AqmA+fPfs3iWp6JSRbEg6fX9dB4GClfVmcJZuLu
zfrv7cpPTg5guhzhrbIe8v+/cnBz/1Afd2bSnFtRmx3G4M/rWkn3EyF1j7t3i9np
j/oJkNZzu7w+pxTppOdXFMJyBsELmi2ST8bwCRsfVsHx6TLnfEJYdVPlmg3iNX2b
tJZyLga6rG6/KI2yvDfSl1QXtpaPuQxhlJlL5xnESMuleLhGGrJjMGvHcNd314ad
Lj6YhmN+pmeM/Zt3qTqFxUFs5UsD3tYHGejiZEOwoyX06uXxlsoj01MJ3I7INvO1
m1v5243abXOe/wSz46LKwl7/HzAcu+qQ04YW7QcfZs1hxeWFmnhLtCzsQ0oWZnyK
kGgPrQTyGM0Z8I98429UATbUMpEG8Ul5BZUx61wJSqZlWiu7bJVFBmFmKVDk9TIs
wD6KpNin9sAmvzP4Z7AVBwk1hF0SxTax/aTq4LzahyZWbXkCr+e4Rf5Niuus7ZmE
f8ddkMHWfD0sJC+64X8+TmW12AoAwUhtHYMU8uD5oEwNgLx2RbO6/AajWZA0mTAf
EZtrNumDjx2WbjKA/V1/ZIvVSPH1YFT/6rA3gj/2EgBW57lB35ecuRCwBLDIJEuG
oinBIKAMZ3otRYNWzfeS8ELPBCvNmK21Yz53UDIrnqk3xZivV4DBeSWqw6ogVFwc
hHdZJmKpCrLnnJYOgSQaeajZQaFjhhLmnE8ceg2/XnV6ykGdRuCs8lBQBA5e2nB5
mGQvdn0eIBXAnBPexzDgjNTGa1Cvka/xNzNczOUQ3g/NTGt7c/q6CKDlcNDEfNSs
CNgdenZuH/P8N70eFGWZ/RDxrZj5JsNJuhA9rKXqSbmJefBfpnco2Ff8s1r3ycey
ZwVgSyuZEy+X+2UkSyV6Ty8K/agkkurtcwhJkXs7DvWM47rQNeWTQ+5JtnBU4Za0
uKzDz4TfFFF5Tdo1SccLZA==

`pragma protect end_protected
