// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
IcBax9mpAJaV2gZXsLsgAYjxrrVUdZByJgFPhJyfru6rfM44VgnR28E7cMlI
u10XQ8gnBQPy6g0wegzM3lFWytp7Azsk8bXyJY/YF4K/t4NZLQlEx8QHtkqG
Rxhah+WXxm4bT7LzuukfQdJzlLMpmiBA5G/UIOwyaOoTTdvFXq2VueOHX2vt
6LdVw7aA4PVHY3Ac0io7EaMZi/Bhvv0Um+Ni9rRBIb2eClNF6wGsau3b+osP
xTvlS6CXlilFFKfWfZSDib3ss/wg6TyP/KewukREtpvdCnLACyDGtRMbSOTL
EqlfY9wjeChGPwFQI3Cf4go8jg5yGek3wRsUth3hzA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
cGvnppWzkB6tnKTcazt71O3ql2nkOdXIwfmCNz3vKMjs10PdVOqjbFRXQkzA
MGM8Ia17P6RcPNe/1Plpl70PW17VKNnfKtRIcdjFqWi3yIJOVuXvMMhUTUlz
nCrpUVD+AaRf8P9mSfW2VE/wxy0bOl+fnUuvr1Q3XmUmaeKbTGPAgGbpNcAJ
lLVCjVBpYKMbb7HaJUsXm46+JVzVANlSma6tej2OdXkmxyxFFQsyeluGqJ7k
PLdHApDRdWt79JDfK/M7v5506yUYi+aGMSARmieHR0SxImva2pHinuEpoKJH
0diqpE1B1kQlYzysx8wS38KElj3uF6XQf8GepvFqyg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
pdOCnrW5jbW4cSEiPgp5vI2TFoEuUZDFVD2z1gW7Th+HPcCIwZVAGVKAIqfW
i2YcckOPEfxY/8Xa4BP430Q6hi178rLIY4OYMX9kxlH595VhLalDr5MbO91t
7oxAmpOOt3MITMopGO42M1us9+9+c4UDrNiwN3SnT1Baw0iwBJgD6paNFNNn
nwVXHqyiCkQH1oV+13iNDLVqRJqxMkh+/S7AG8nfT/aSBrBg9jAxwuPy+b+A
97VaRvGJUVMJhG29+QDDz4nF7sAkmibE2o63Ov+L96gTWUrBFte+MhShvyRI
PHYiPPphR4ozgA3eIJzLZvRXML4vDcMRNrj56+nsdg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
PN60Bme3LFUJZFq/m43khoCCBfTtF8K8Qqonw+leJ/0q/WHiPB830u8mhRsU
k3CrrA5ljuqDQVlhBniSB8qNZ14YQFik/RSIK1CKYv4pdjBHE6IshIV/2237
5pEEx10LGeP03cSIANzYyM0K1DMdHr3FBcZidiwhmlhlyFvWuqo=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
yKrU9hFJXEosU09KlGlA91T53lFMeWraj6C511Svo0h+CRPw+nkPmQ8wkDjn
YsYHFppB+AWiTmQeBYyvtHrJzMeLefZJ3lnR5Ahv+SoarwBCyUVyXE+RwIHx
hyOrhIveEEMK7X/h6gfxLviL6YzUVDmihwYyp0TXFDcegS16HrtHL7dI6vIf
2ID4lCYNHfdP00CITxAlGz2rUO2EuqRK9RZefifMkc7hxRFgqMGYGcLTmXph
pLvgrq58KHBRoZqwjoliXc2XPqXBSuqnYo2oUrfjP56fY1/piCznKOpa4P83
3fPx6YMu+ExIxczbGnXOsJIDxWuMLaWjAfJdOKz8ezzd+wD+0c5VOGeaDRK7
Iw+ckJn8PcB58+ReLF1D4vhaAsrZvMjKRFqhn1z3vTxrvYDUU5NNG2cKXe23
pPfGNNTSF9GPG6eWwCl8PiAMdNfFrwIUDBWobQiC4fr1kSIsyf/mv17DZ4TI
Ch8Cf6Ea4JLWRFsMZkpau4BJmonAH2/t


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
cNiAi54UbV08h71JU+HoUBNFORQineh5BHCVi9KmpS7Xo9X7W2bH1Xd0qa9H
BpS5IWisd7Z+Yvjz8F10KTmPSYNuFgeoOqb6G8REhvJttQLYk4t3QceESc8n
8g6XO7h0XzzH+ie+G9G9lQYtzSHHXzHI9RoCy4Jvqr6jZvOzYp4=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
kWbgKpby9Myp4MKy6C0aCmLJJtDeuZZrJpHzXLYVYvacbNZPN2yklgyNzIO2
Z80OGoe1ih59uIXDX9Q7gFZ/54NxwncxwXrIQ2U3Ht6BZ3q9L6Fxn0M+wHFS
RQkclMdb2btYJls3eEpKTl2CIHxG8Z22fP/pyD2Xvx2n4HtkbhY=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 281168)
`pragma protect data_block
GeaMsqjUqhhqdZVl5Y5VvbxON1W7gNT6918YGSjUV1F7D1QdPkQJ2rb7zIRR
UCGMszdvN0Fcv2CdE9mvZCa0+Qbb4aNFdkxZdvMeV6rwa4wwNKASnOyXd5ko
7CWypNjcUJ2M3VagET3J/tvPVZfwAFSA7Y9NF7FgdGWdApapARhm/b8+X6EF
3ZBaOeRWDpLR59YMJwlFRELe/Y+0WpBxzfLr7Sj+AIOujc/+Spm3C95I8+Qa
ujVbc31lksdaStCD0fSacC+Dz/hU/BF0vn9yOfGG4z5FTRHG7f7NCBiTyAkH
H+eQFid1bK4ZFZxcixTZTgaV7xuTG2LUk4NwMSzgAtDy2bf2qx6WLSoProef
LME2vn4Zj822Uur4FFzm6Nbj+RYaZZvyiA+D0W+uCE3ixnd7KSiKpumZuTS7
RFoSlsChTS2nyBh/kfXjaihFmyTSacX3oivccCRkUXkqiva1bHJ8XEi+Mc1B
N0j7e1u5v8upeSW2hVyFZlDYqNcEvDKpvWtBKNNgpz7rCzB3GTlZDCrO6rpo
Gl3PIhABkejH8TNiDdA9jTxiCfk24NLqCBgHrbMqM424Xf9tE+owx1VDgGbI
PWv3UT9CLHdQ21O1QTbrFKthslWrnpKePQ6a8xY3k/nhYbZD/Ufk5Qz56t++
3hpNtT8uTFz29URvWhlaz2AJIHtgzcHBlcgB2uvemS0kjSIS7ikYjTuVY2EG
4OKBmg93URRN9m8kZTcJMRPZthlXPtOOUUv59M31W6TUp1iWV8aBUDHObgq0
sebGP0vPWctxZ1MKzDDagTbVLihtiy2pc0XLB2KyscNVM147lz7xtQ31vzBM
tlaP99XvQiXbr+ZTwb8jRhGBPOb5X3+B4tr1/rnhXznNbFtqoO+o2B3YS6qb
F0BwmtyiVNqd5EWA2BxqJvVxq0IVwdv5o6W/Z9YMLmuEA7tSJKBJc4oO2htj
ozCLgMdP9ebYWE16n/5NoSG8eOEbCacSN0UKEPg1oo0yiPT0fhylgLFMBthw
YU3wro8Q/25wtxwMtwNzuXpVYPZ4K8OMJDEurInBh+FX98DErZPZRXqz2Qch
fa6RIPFE8otN1rhOAH50P78G1DL5Hg9T/m3FsZUz7M6QlbAGkrRLkTfvoieS
JMhqOA++YAXuQN6FqtQwhwnhYLOGaH2zLAWa2OCT70TfmjiveaO4i7aBUgUY
183HEunnZvXr2GgZkecIcP+v2aodyxdRqVGcndBzArlQGLW6G0GgYtkeOYwp
yv2kW3Gd28MEFmXKMsKLG8qZXiE712gaFS5G3+PML2iuPw4u/5Y72AsqaddS
nOCvzr9Of3RBtpQp11Zhyhmbz9KmNccL21kuinvV4dMGMThBSH1KVSeBdI4U
o+PWvS5bUgMENAEK2TthuyUxF3YeZzA567cRyZG85pzTtCt1Ak6+nMq2tDaq
qmv5m2plNh79S2SI5zcBhlQYAmgY+mj4yGtMd5aYJMdCAiRhE+zUhhekECu7
J9iv77Xzzx0VrSO/uHBWXJeQLxUylf/BVS63scz3CpoF0NQC+rq4oa/+/uOj
RBbaNYXvoioVEc8tJ7IRAzfjzJiHoGH372XF63LkNWe6xGGgrVRnAIcQf+ea
U6JYoLWcbM97+q0PBcp8z0cspSmvvpc8iwoxUZrmekIo6FlFza5WuJjAoCKN
uROzHziT2Wk4bR9bFn/BD1s6zK7ToDooXnbrOkpjFqfXMxuIhS6xD1cDEHla
MKrBCJ3kunZCPx5il39reWP01IX8WnQQ1BomB+T4xzzdxDM8TrHTgzSO++86
vvNNTfaUwGhjgF8MFO3xmNADePQoVbDAXdA6Qrr6LBY5KzCtInY3OZXy4B9f
KMEY2Kzk3B1HTiD3t7d9/HAai41I2PBtv6sUp1sDkEGFDehuMWQ5C5GcS0I8
+u8wnw5TY0Hc48kZx3NUQQ8se2DoKYNwX1btPavObzo0kl0SdRy893dqBIQ6
ptNXXKpUSql1OKlDWoJ5aginbIFYAGxKmcRMDTxlMM3/z/qU3SpJuCqRmdVM
rTE5/jwc78wSjnrg11bRZgFq/5waH0t/phWoOOiY5xnhngZz+WVzUMghlWkL
gu1/PyntUY+CIueo0U5q9X62dcuzHeYdFuIDwqhD5uQzgXRYZHDZhJcC3b9+
KMk4MYYKuVxWwQ7VZX2cimyvJMtrMkRJoqbsIomrU5+j7Zu4sx+cDWJsYz0K
rD2FGVWgXt3H1T/55agBnBPjF6Re7hXHgIS9EdIc5gztGbCoN1i8xwZHT7hN
YC7aNKO0n27itzc9S1ZcZ7FD4euFcYI58vBwl9ekSzH4/pk5Gq7lByP8L7Qs
8N3uPK22PlHFKGsdE2BNWNTKvwO5OGF2F9pjRKULquBTdYGtcFTUTYIgYvzF
fpOL2WTigYRA5WNwsxgxAbR7d6uAUA5wQ004/YE1VdHRqVDOz3XOX3nmO6SU
5a7jB4gLydK4lORMoodhxX+r8s+PiWRDmOJWATj09b7zz9uIEsDplYXgT8yH
p3vjzOnLgLQ0uLydzlTacZHGi5yOBoYgWNHUjF5w1wJJwyPq51U4GOSAlXBQ
GgUpQ3mtHVUyTBdkCc2jBCzu5m6bsNK2Mp69yf6Y4N1a+frZ10eDYq6KkKfN
MbjuUEQZOaFL567InpDK3bBP5o8i9SyUDiefNCR1aWxxjC414H63xAjL45AI
eD3VZG1Dz5Avuep08UIfm4YNa+IyCSnom4C5D+4x0MS1r09wYbRY2C28dUjV
dMU507ERd8kgriUcV+lrOSEXYv4nzIwJltLkeuuM12eOF4zy2HMDCkgg1axc
dY/B5VbBm6Lrwih7iLnwCu1PifIRMm4ebGHVD1qmFqJXPu84+uS5AlVr20yd
8OR1WvVW/WX/rDy0Q/hJnloW5PvizE3OXCLtPIH1xD/dStqxGESYl7cylcsu
J9+/22uiCbzmpug391I9Mbs0cH/Bsp+rlcAM2q6R41cU8vvdT2fVA/8UJJyw
JqfYfx6+HUlbddNEwCtyQ9SK9Lac3wTrC7Wl0hoBNFyvpgjtyPPKBnM9HJgz
nFsPQjmmOc4IhyUVXkE557dGfDKWka8v30h1FSN+50nQqo9KP+XJt6FirRK1
4w+mI+1cnetAYAK97wSw/pYdXe9Wwd6mIBH715wFe6WGmcEYX0a1peTZDmTB
pIgDw2gNendEv4FNL9wUMeWjDHZ3wo6UvrOHwu/6vK5Z0lhZeGdVY95sMf9B
YI6WFx9YLXbzxjm+9WMIE8NEXE9TjBEg/LnqigelJ+sgfaYgogtYeygjNhVs
T+lfb9iWZ3mt7SiXx0Fy3DGEw8itISxnCmlySm5XDSFX73kqMzKo1BkkcnWA
lQ50EXElr3/28WyZCJjG8deoSGZqfEiCI2gRUSl69tkAdzUGnWNxuoN0aFsZ
UdMsKQ86iyEBwB6lZ3Dz2uKJ/izCcTQMseRrfU4Zm39KHDMlB9SXVrfOjGP3
msNPAy2vsw7sAzUE5hMhqjmj4zSR7tyBCYuoD+qjNsnFRIzYe/EQMUVC7Xsl
FrLtRLeVHlQLXsXzCI4GILsPvcNFsQ8ErNQbC8UP8hcDXbZZUqm3dwgbICKW
skHYf66gPiTRJG62qBxe/J6KCcttttTcv40tvu4h8KQxN0adq51nD0318sRC
hUbzus2tdOcSmYitRroqa2XhXRwovLmme4L/RK9sJO1NI1nlsyRAu9cH4b7C
H6G4jALydSO9b4GwNIrVTwo456AW1xHoLhS81N5dX1CeaEC+nKzi75Na2ZhG
8gvPxuDjWVLkKWK83ItfveGxhDuZEmLP/WiIVNS6lstEdXio/LnSj1+Lq3HS
lfASCfmIquxpy5VwSfObIK15G3cIvHUC0FU69rUFa2QjCvFkmicmsyTILoRs
xzOywlnJZGsn6heWgoEP+E8a6xw+xBx9Pnm9nrbuUH1s4rayyV64+hFqTNW/
H8YExZBXn4/QNlWvvf3tsQ4YjxW/5/QKywvwGgGuQie5SKZvc2qthU04CUCo
czHuaKTCE3gTQVEOsiw5I+7RFeSzAvdWbE2l2P7lpy6x/n2UkemZ+nO/O3cv
r0sut6ImB9ooAFzUo++ERrU5eF6mkHPPQEQFhbSpXes9a7VdqsROXSxWPB77
ww3FJm84OTIzBAcSpNExyDq325LLn6MfP62Uz2dfSSn6G2MQQ4SEOKD+Q9zP
K0EMJSIdb8H8MJOzy3lC5feqJALzFrvAwaFhY2ij9Yq5tcxf+es49Nn3/Mca
C4LJLwd4VenphXK3KnWH7Zj0gqB4uTLh6Pj9xZBTwyM4Os7Jv3y+MRUfI0aH
s/CFNtUGj5/KHKpVJrji4/uTQp/itYeSBXSh/eMMHHa3OLfSlf2Nbb9s2hzZ
D5tpF5EnAEmfEHxupbwfpsrYMaBNM0+BV1Pjo4gJVN4vhYVi5geeG4VJTuah
1J8EDGgNB2OmaQLoYbg+Rc5ENLxwfA8yTcqNmEnVmT20nnEQE857fkwdmpMT
3hB109CkEhRVZZtvUr71vHwZ52lyWL/fXT6RyvGrn9BHW593sIUDqG/OS/KI
MaJ5GD0GAlsrBt3tdhR1GJjkXoL+ibWa5tIAWv9Ijkd4DBiJE8bkWA1lkg9n
xuE1RbBgsOmqmv92BlCF+mdXmbXBeXDcFJhwaZLusUZ0gXirDHs1Gd4O7qO0
dq6mz+iuzGdZNwBMrRP1R0zOtPWN36aFv5a0/5k+7z1hRlyxF+DGJ3p4KQTI
V27AZlvc1X2M8kdV7906eRxntCDxzxvhOlA5fmgWJ9ErX7WEAiT1tyOJ9KCg
bgPcmV8ECS/chK47/NQGGM8x6gZQYVUHmjsiSywoHfYG0dSz6VqCzFOnlJwu
HEPgmKtXCf7Rk7IU69PpgRs+p3gYnEsQDbD6Cww1QuBPNmm9H/229ECTlib9
jjEmuXwcHlvVrWVkd2wEEUt1b/dS1KTx1BvBiiYCU2GL9IIzDfKngxTx66py
0cpxOHm3L6FAV0/Jfc2KakDi9vei9IKhTkQJEFP+/68jlbPCU6B5732cX/c+
d4/QK0tXbi1uajA06vcUmGSTb+bnjrz1LDwMxvDhVPNxwJAzacPLkL9WKao5
gYJeUVkBSfZXsZ8+LzAP9SKiJmFHYJ3Cij6yPZVe5JaIvM4dbRJrv8T29mMq
EFJDwTpIBRRVxAlnFfls+2nZD2gI63sfmhrEqXg9DPnwOzcLRPTj9t8hS6DU
0+1xsRWs7934DWQnB8jjU9eLY6snmnOtNOb2os+f/n0zYARSis15cim/LsM5
wJ2+OPLa9TC8mT4f+bX/R+KSI2vMBqaHhY/GB5ewvx1KwPc4jbvFOpxdd3eS
XjDAH/XtH5dqo6mUTXwDDjuYCZRX9GaS5PIGeV5GlsvO99s9AF+aGWCVs2R3
bn9LK1uK1a7qQEbaR7FuEDT4JSP/0KGox/0K6ijyofP+Zmuvmhp4eq+2G1am
zn8InOPbdbPGojB0k8fsvld5/FU+kVWuH9eBBjCAt1W5oKkNIfPOt8e4IDuR
ZYLUmTtkcVfyC2Z5o/zAtaQjElJF94+GkU1xV25vK6evLiJjJvQeVfsfCPFD
ERyj88UbVAFag0gZ1xN4r8rVzUPMhKV9TN4pHwrDUwS/mde1Iuqt3HFLX9+B
CvejxAZwAgW7BuB7BX85I/FDCVsZGnFCzoa9DIxOifivxZPOgnWEicAQgWBZ
TDGlcwOouJjtM65j4YpoEoTjfpdfmfCcubmI1vpu7w56e7sdN35X8RHRZb0b
ps1QnmtF1HgRSqgfSieggFOC7nVPWJqbT+zoArnayV7ToF9JJhsbYOUIvsAd
C8kpFQTjBrACXjtWA/GOi9Si0LKV32FN7ZO3FxXNL0JQ7XJe7JOEykMZu5oy
lfdedlMYDaSfKcPx0KBw4BIc+A3XJVnKoejJJZrYaLkO+5dW2KePnvzUJNhb
lV9pzieSaXHshBvvyj4W3GRY45OQatM02X5yqumIJq5AkMFAyEV5rw3L7Owk
RZJZsa53BIjX1LZp8O+NbTnA1MzzOH9R0j47SQ0pd8ScsY1osnK0Ndf+5xlU
V5E9+w6VAd9uXttih/C515mfiopEGBJjOurJ3Mdx0oiVyRJ7BRBUTZrtEKbY
Bpw79NGjsi1Pn/Ok4TvNAb6FLEWW5t7lFbZ7E13jwPayeljz+LxfMUprIaFU
LK1OE6lGOO1lY/1OCdDuq4z/JIT2lVTohYsySh5SVnRP40QU2jXYxNM7l7Me
EJVECddwtD3q8ZwFoAZ0YMsRd17r/mNW9HgLzmCQ4f0FX/j03xeuBGj51GEK
tKeFaxj+YyQErRq27aDqlvAh28c3HhkxRka0WiqUTbo9SIo3bNdxNA/fXgTQ
lfCuX6DP1tyxboKS/Bof6E5oZnyyKjomrx1iMefajds/sn0UE7qIykG/6Fuk
A0uEavvdVeISbFTHEG88xA2Ze0OgyRt5eQZQX2OE11cxObEwh9x0Bq7aYsWw
7hZxT6lUf2QKvMmN/EUrWUoFWU8PEfS6iOx+e8F7ZF11W+NK0kXYg8gxkNnI
8Csdi1ENO7MGDRoM02ri9pkeE2YgMDvifazg1Q4pFLrf9F4s1fPMF0+2aGoz
80qv01anY9BiPGgYa1VNaVPi1yzFs0OTeFe/IMQVfnrMXlcrFJFbG42tR35+
CqgUPafa4lOelZkk/TJep5GxAQfEhbG9KX4vIrEVy2AVbKAqfiaZB9YWIGxu
6/iqLzF+OOpyIwfebcR7jww/7v4oowQz9yCdBccK4NUuCPbJtDKButbMpBhV
03K7kxl3sxDYg0ZV1BnUO+tDvkt/PfK3hyROUxg8ZDH7FFP1NR4KriJKkVY2
3IavBUIIxPJx3AkGDCYMYgsq7D3nLraJHM01hL2ektnMCzSc7xf3CLl8BckB
ws6k3tq4iSewFrVhWDuAkTVCvsx7hwzXDYktCRirQAWtWQ+VyVPL8ufCQgdj
PRDwWsZhwxnVuHuFrQW5GVzZhhPDRayYtujW72aL/F08Q/WHX/o2eKEQsTzm
VYyjiCFmd0l5lw/INeAkHf6TPp7asvf5fmOTVflcZIT2zWbFxWLsBa2MuW56
+zfDEmh6Za6JwryN8YdD0ecI2NAiTPk1UGHznKp+iq+QrB0YO0KWWJCStDr1
EUY3nTopKJjQ5LhCAxdd0IzJ0G9hwCSgwJGwMRTIJX6bBETchngCl1onnP0M
BQPPDZlD0YhhjluRnsUcOZKbfRygj4Lrhaysal+cSxdXY6D+ZyZhmJOmq1mi
eHo2K2tWsgmxWtrDZ67s0dGmYhA3nXeY9/gzIcYs3kXEEWntqOcs7rMarR+E
uxz3sEKPOckJwPHFHWRyFNb4mNpLlJHekgu4IcjNI3/QaJKeRz68Bb4lwrJI
N0V5vjsNPy+9s9o+ywU4T8s+2zAYJ3hMyfMlIavcRxz6h9Pni+0UjXgft7Ex
tGUM6MCdc6KV/shWw4mmk6sFW/K6KSNKul4CV3hgJynSD1VoFCvHpANBXnP3
JvFlUuWsOlNpYP1FLnFiuJowB1xGscdc7hIO49Ds7l0jX+422ENHJFSf9Dca
sBhHPkenNgbHI91p3FmqNLg2JVomy4Sbm6jvjxrG0o260Wg0VPaXgJZ3JBZT
AfcOPHZxj4xH9cl0cUNbLMxB3d6b6S84vEZrs3WTst8YiYBpAzaR8lpGuGNB
EnVyeWvfxMDwEpGVroePPws18xIvP18xD8JyU95bp6ahabbkOIeS2quae7/X
FGRPY/X0osHgVEr+jLx5FsryrA56nFNq8LmC+l0709wBjw+kutAyZb5om9Vj
0FO6O6CC/BhChOjfdWb9C12qyHy+DYoo6lXihpAMIzhPtEvJhOIRCPv1R/q8
bryYE34axuul6O2oXTdsDdweB8dU2XWF9gc2WBCDOqcShEfOqWsxkEo8ZSap
fbBxdPUJVq1nPsGmMW9Mw27edAVKeFF6fh/Z2iQKa9vyyw25EoDlVoct+8oR
NVwU1zJFQiJq9dkU6jwG/kssjOVCxbTgn7sBzohGYt7POIcUWjmAs4U2qa6V
A73VA1ZJwCJBCzuwibvJG5F8fa4JXjFGPl3wUUQNFnBP+ybHw/pJpnfFehdV
9G3MbZFURp65XHB6dMEqgigmF5zPt5bWlpXDNdmORiTIXL8HZg2JwDszD7m/
B+2BJRG6LubCCjDth+XwxgwwxPq/FCFwxKhT4O47bgaOCEmX+2AjKmMyrs+/
DsL/P4vAlNnSfO2BVZpLcioM4Muwk7z1mG/yZ6s/pFp7qv283VYWsBCS/Rwc
Krcub3Tg+HrUljAUxFMKVnz2bwarOo8VJaFM2avuq8Qtef6FhejlIwkZfKas
0oH/UJppd3+GOZH0DoTxKMsqa0xQrbTvHzJEgXFHb1RnfVIogqWCUHOcW3A8
6Fo1sH1iI54Rg2glaMVUJFV9i1Gx2+LrKkYdJTWuGT7xnYjfBDRqc3OBystL
o6vbop5BvH1rv4wvGOqYncwsLwlxNKlmtLhCb02jv1pakH2ix7GQ4NnhoPGe
I+kwwCQvocS+OIw9HAnFpEk4u0ac7ME6sF1BQKTLgO47LrSXYhD6UNR+9xFF
D+0YW6pvI61ZUbjrRm0bBTEy/DwFVDv7Qosdth3B5rAq8DAT83gGY9Dj+9KV
Ka7V9bYTfsNvVFH7WYSixI0Zi4M3DrxurSLKOnbi7gIBc5QtZ8oSI3SUmh88
vurTY2x39yz7UwBk3xSIcxjzjBJedj8kc/SSDt5tisZuzU/R1AvztRdWRjN3
wncNFPPD3t/fpzD3dKyZw725nM/LQSKtillHxwfSGBCEMpAMKYQWJ59V0LXp
BiW5rqqKBuh+l83COTkpmK8etX3WQ3S4/1eRlk9zlpkko2073ghdegoOiJYq
9kWL7tjr1vDtBSGQRfOZBvqYUf0U+lOAjb91J/DPBW8Oas/+MS1ADYdlJ9YP
W5plnvFY9HJkLrpZGZRQNnMowiPJlaRAw7kWfKnjxVovW4wfqIecVB40gswc
7khL2267E9Gkj4qPsj4k5cDX5L7rKMAvcFm646n4g8QfCLw80cafZsYNHMKj
059httA4548lKkrl4tYVP84ohgDihskpmlAwvs7pEkWMt0gxENCg8vun5rUV
ppVDSWZGTnVcSeV8HJkY6sEERUIRiCix77gqi8awabU+sL4Utc6StU+D/w/V
7i18zNMLUq72RacVRq8BFshsA7bQ6PmtzGy7Shfk71BNjXJlr8QuLBTPv50k
4P69kFAbx6ouanamshCIb6DqwP+Yp2XJLOD8b+Xmii2uBaixfMKyclMZWcJ1
yijh5SLD6Jbx2VVtzxLooy+PKE6AW119A3FOabUotsUY5kmoLUyas1THFELU
kf5XrqNZpPjwBpsPzGu0DVcByoKMqjgYLGWIJSrDHLYhYfEMuVSVVCoRjs5Z
L9hEyPPrN2Bzlh3rFSChfpDBzUYAL3MQnS8tDlwk69c0uAiRtjDmUdCjcojT
mcNUU4a+zVo3oadgJ8dUH07zonJrqg813C7PgLD5h8tx9mGTEs13zRH1eoyA
VI4P4QWqKXpQ7/FWdxzQ18nqXJ3/NscVOFVmZJQlHuMz8rA0/R2+SVmc3hrW
kC0ZhNKq5cJMk7yKY4o56UQW6sQqGLo3atxs7SD2DJjDyz/cT8OCSDZHzkNd
tvsVFQkv0mRzXvSxSVHiUXhCHrGNB+j3lJRBbBkw10RQXQ27X1i19TmpjYju
ivkX6A0lV/9M7gVTSDKxX/Qghb9F8/db8vFKT5r6/EDGJmR8qlHFo5lahHC9
xt/6b61sbGPIeTQ9Yc5QsfnC/Wea0hxRTjHPk0YVaUv9X25N+lvM5q2EB3Wp
nCvNDANGbrWxVOQU/YDPyoYvhZphQ4TB3Bac0xkX9BwEaBUfUpEFLD4OseNL
7qiV8iy2d7nWnIkDd3c2RrQ0acuGCG+ECZZBa9tJvALFU6j8hR+uZvuARqY/
NTs3H9oauP4xQ75QiiQV8NRTM5xl8bf8sNOYXxozTBGxma09Vhoa9qQ6pfhL
wlx+Ei19Wr2lJjOBsZ82Fy5k+2B0GmGAaqvE9bQ05HAqnjwL7RIAzrkUoSLq
dK4T6OgW9Hlp41ASFQWtB7reB9Rhu/sRxhYCuTSmfCn/tqM7JY04JE7JhZjv
nJvNKs2iuQ8+5cyG/1ka0m78rvYIK/A3v7uSihtZ0ixCD++FvYZHN5Bjdkw+
vO0aQYqS5Alz34yCbLiPJB9+Yx0Zfo4LRe/Fv1sa3dD0lR/XyDnNV7EHN/rl
LctH0w8dfFAYqaqAbt4wT3LuYanXoZdi7o49VfZLtCyhRpyPHmjdmFePkhsO
YXUt6NMFc0htZfxAbrSeggLP2YrfOAv7YvGxqEUb8nHNvRECAdJIn7/StO7i
ddERFAydFHSwPlpnb3jcZMeT7qeC03J3AvQK2r59HSETyvBZNlmhFCggdVDF
lqzj6e/UNpiw10Uz4QFpg8hbULd2qToSo3i5ryyItuYpmJxbYpssnia60Gp/
1PMgPmijb4IJNsY/CRRB59FQtPSmI2CWxHQttUWE0mRun40SogRlxNiHanC2
JPXc0zErRsf0L+9+MxNYh6k5eXtP4KApy2I+z67GzFFRFxikxVkiPYpJEqIi
7V1TF0vFJqLuMmwYXNc9t350P5kaT8tgKBmgspMtOopzs1r99sPBNmDDGqkV
Tx8ZqHTYiW37EQybY/aqaxK7ZqFPuLbmGthQMW4WWWExGh+WqyNBSHhq8lC7
V+l7oNPv0FLoLoz/kFPeYI+3+NtzIHFghMI6pK2Js6MQbmbRDhBeUCXxpd23
Fogx8iJKCylKIJSLX4HkgdH2Oau76cAjgUGV/JZb0TQkVw4xNbWzPFeBjejl
RG5O+8tLf7goaLvFgtnvZyH3MtGwAfYXIroqclHuWoxT678n7xOy93gL0cMx
swIA/YUnl8G5T13cr151JkD5iMlG59PAhoRhRUTq33TAJihgyOpNDCHfRwxa
8y6KVaRg8Jquo/IijkyBwgTeVWIzlFedxqy5eJLnE6n1OVB7j6JhMexia+Iq
Ik1nkbuffdU0iF5/VlHfYVne21uyaXtyJCwO3UZPOLCtupo5xY6nBr8917Gh
dMMUA2gJgVw7OLdOPxC1yHjGtiQfxL/ZmhUxWTeZ7cTaNVphfDsOI26SvJzp
vy8bAdSP9aYvvrPfo+0XI7S8xiD+Bq0DytZO0PhOjLBdsS0Ir75BEbZIKIfd
UcmDciKmBbjL8pP6VXbvUeNdXcWeC0h2BAlF/KEhR3cP8o+f77sxlnNOca8T
R+NJ1vu+cgwzbQBKqyR8pBIBwyfq8BnK2ScIZJTOcSsZDVMz0+wrT3xFPL7P
LwRWeHXFPsuFO9lHCj4fKNZHVhGHw7WMfwOcslo1L7TE9m+i/7v/t3H1xiJi
idQG469d49wHekfXvzZnBcotkF94mtOBy8Tzg5iKry+35b2lG8cCr4C3N4OL
hSD466CotOdAhraoChqqpHbeMh9YKDp0K9id3G9VZ3Wm8upcdtj19kFKg6L8
dhfLA2589F1u3oSPOohTGg8cfGTrIPMytVxNFVJQAAVE49q/1VYvr1P6q/1w
J2kcOmVxhEmH2+0O7+Fds1fgZhn+uyTTrbNcf7DLP3luWxxqv6n9WRSY0wVO
mx0G/8ic6Z0DjZAksgQ4++QPFFaHHwCjiYjKpk5KpVMlt/m8NpCWXG8WOCDi
kMIkqWdmkKsetKXqyqYmbXWF6kKqYOdriN/VQK+cJndk7uT1l5z5g/YgOQPr
F9gWh1QUOb62ro64FJf+ljUxAsLmvRt/j/TEZOLxiWQbJCU/risMRk4MUVjw
EXMZYTTb8lSzgnoMSb2QqYOXTENzt/10xd4ZWFKxxQDtpE3Yr/iINTj/+0yG
QPTZqh1U0xWas9nVmNER2ITOhnLROcYAyVr9k12YkoaMC9vyiF6lK/c396Vv
uO28hgxfwFMuJZm1nJt4D0tu5gBDG6HCWYAsTfiLck/YyVDvo87m0LLN9sa1
DM9lMaFi1ovpp1CMXoiVr0Yr5cYyGLuXweMx7pkIY/hV5aM0RAwe1UnlPPlm
c55HC7F+VwokhC654YtRwelEQTPgwYKok38Vf9sf/eEO1sgokJY0BGorIV2H
RF0gwLrJlfIPFiVp3jS/ov3M7XZ3+AZ1yeVcwWbr6aH24fwHGPcUueoKE4tt
DY30HZdCa00da5f9OKgCnGWYNoqVvkamuAqNub+IrRGBddPvOKH5FDXfooAR
Cw9gobfY/VHLY5DP5hUqeEJrQXqZZlyb5TeQJXZqnYsdF3LuykvqnUnspENy
GcSG7s6XJYK9jI/JMuBM/ZmmXEHm0b776ru4XNWzOYwtt42cGMbfT9u9+K4C
Hu2L7B/zG2HAA7kA2o5XqcguWHSTBPQCUqnRxezRwmaw5CwmEVCAqOOY4hqX
/oZdPI+SQL5cI0Onb0CcB44f28EIWwjQjVJXZ8vJRViTq8AvmJm4PO34t/MR
TqCDfxKz6oqBKExTiqua5Or2S/Bj7nShCKWH/zxxCHU02KPGBRczn6sMzKdg
ZOlNlNxBR/nUeOFrH9UTMOKSlilbSFOpvRV2I8xsF41QKo9dsg1ujEOf7+By
CRSG8b6bTygiONK1TQomYrvOc44PLmioVDtt1M6cmjMwmB2gT3ERMO7nRs9c
u9naX5AfC4OuHwYnNH6RPQfO1/OCBQ/TxkLCyMxMDB4tPgquc853X+eko9nO
TMlUK2H41hoz7v8sjEe7qm1y33peDhNiVQZhT9ezLdEBEOlYq/FEzJT5EW2M
NAZ65S6a6+AhXs+y7M/V+FxATtYmO/mY8QSHJWXqE9sxpZBN9xH3EabVW0xn
/KzMEN8QrvFkgeSh3E8CN0yi2OzWQ6VFfgMyLF5icUeRExzQPkPvwJ8LptfU
E0sbRcWvRcEhFPITujPMUWL+EVWd6Z3DO0Ab8ytHw9+hUfgl5Um/C3hhei/X
Z+q0tD+1okxadFGx1PhyAldK+KEEq5m1vj3XLuFKmJWa2CCyk2Wr3IgWYu83
RpGHhi+r/1XwJtooqjhKSjoy0pUdM6LKDBioO74Kdoe8kx9VS7VhlzdhCOp+
LmJ/7bm7HqJPvQ3BlGJPD88WC30xB191+OQ0zqDrnnDWqVZT7w0U67ngpO5T
dc7qLpPQVgl1hyGEF6rYhRwkTd5rFwN57w4+vqynCfi1IxzfKhYu3oxTCjMR
3UbmvxNYB8wJAI/eKZRVEZzs7tTf8dlgxSmCqD7ldQnWh8fYBYuVwZWlY6D/
2a6xUfZ7Fo4QzExsv8f+wVRZu6lEj3Bp7TdyOsgqiaqH6jcfv5eX1DoC856h
bTWBdplpwq0ynNgwJB8CVNHBDJT441wzRPyGBUpMCReQ7xFcvhagHzVYpr4L
7O6JbHE+MpuMdqU6QnUNPET7gB8nMT4ONzbKvxJBSI2SPWd6d7Eg4vu9O8PG
l6sGW9041OCqNQVJR/nsvJhcS/BvXRu31ndVrzeUl8yJxCGybpbxrYcWMaUD
nwkNXMYN9xj8ATaJEkGvZ6cwPGvqcLmkpSBCi3UNUru1xV7D3+BqV4YJiYui
zi8DON8k+oVkGrPlyqbD9PTOLDSgJgpIDYK8wvFfbTI25zttn/VAHd32RRxP
HWzdqg8bgFfQU7H8+xRMZI+pI8kDNp7rgp0Fakh5i17fv2h2psUi0TpkmiCY
JTAFsjdQ5XkmhflAE7BDmVJLEA2Z79i7HYnv6hwJu97XnrQU6x9LYRmnP62f
pYfHXZdmg3MX5tdRL6Ip1qPbijS33Uc7QX9mq6jGEwwY04+JEp27DNwrUlOO
KYT8sQudvVcLxBkIjYkfxYI6/pLDVE+i7YRoQw0MwioDZvUGD6ptqmOcGGfA
sZjLBC1aiJzT4iUxbQYanjjx/TrXSIYXPt0huUgMy8BdXvBLYRmWqM4IthjS
SdcTDjniLCOXE872vUUloJcuRHeiRst2xhaLmQKDltC380M9zQLRCKt5vmCi
4NyhpAzs5BAxO70uoQHoxSXMhQJ4gmfNomqilvQMPKXX1USGziBzUTf9d/iq
4VEck4AosMZ1QIMOGzqBzznWoSOoiVIfW1bKZe18Gklng+wpNuZ3CQHYNLo6
7327lGsSYiWZVlZ6YTNlwbSAtFRC7yxoSh+f6CI5vhpF6DScgSQx/dqLwGLD
YoAv1qVcopgEtXv8SJx8RIUKCEClUSySL2sDevf5wyNVDQGolJ+2rtKdJfAh
2kGdY3AbINgbP4XSbIIAQYRd1foJv5zgXuRCsLMV1kAicAiPqFsl2HU0vJjm
MfR+MWN4mEEU7qbrbGg39xozc4MTTDVEm5DKtmop1mErymfKSlj/U57WwXVE
q+mwwPL/6M/UgZqcFaZYTSz16eGMtkoicJxmzXyXXMNhz7AxtaAKQ6cLH80w
c4vNZoGtd1w60CWYmi9AW+2yE1fBb7ROo4Mm6yT/EGJiYLOtCNkQ/uJg2Ju1
PdkqvtYOvdu1NIlhBgc2pRjPMwa0/lqvxcAncxzav3nq2d38JlHisMzK8hiu
oLLNJey7x5nTSP3MUdJvsyWuGZO8hJFlJPbNXwG/6jXEzcEF8aYmY4h7k9g1
9ZQdeeG+lwC5nKNAaQaCpoxfgB2ikh2YlmDUS1QhjuzJEbaiDNdAG+KP66DQ
smZQLeUQkzdmr4iC5s9zAT2eC1WGt6sHojUAeKSr081sC+2c8gFPUlPhTLRm
1KXp6FGPxQig204/k+J8R68Ef617hGtQaLzMDhUENMgDWBS9N+NYDjxJaOOK
X6xiLzludV91CbaPUBhTgezghZHpAIUOgqiNQYyyPUITNY7FlFJknH6Zccz7
gV6v9RLFuzBIfTosWqqsqAAlkkO35V8s2DAE4YkoxWQaywoK5KWptNAzTKHR
RRINCHhriADDOxvfqfXS+xdrBEuApGMJ4/fYSy2+pb/ir2UHhvKngI8tXQ6l
akhZLUsKqjglBOTIsJCtIQRAOUzeMYZuMSLJg9750PVKRuUlNhjW+DMNnv61
uY67ZZX6MQZJSluO/MpyFQIqWoggG0Fl9W9nuBxuDhrkomu1F5oNgZPPZdzs
5nKQT96+glgcDwJk4rByOEcF2TQriaANzNtRw4Ec70lEXmvkwAh6peIKY0bS
/K4S9Mpv5FiiZDGTIIvTdu2XKscPF+cQAMPy+I8yxfxM9vv7cum5968xXzux
hEmrplz2vuk+mfj2/+tdUbOd7HZ6Vlyn0Zdwff3bN+yqvEc1QRwPDQERkI1F
iJVN+uD6mfLCg/80jTSuJDNqXWOe4TcyU5pw0vhUa6ZjCSuAD+5Cw4DaR67Q
HMm+LpHX/UOywLxuUAxMN8MrMDT/uL4QPKHN/536r5RhSkWuK1H51ON2HXY8
ojTJytdue76MCYahJhTKN5dPCy6iNcJ+WmUiZtBwKFcP3SR6/0QWVKr2Fws2
eS926DsQ6xoni86r5mOkaG+hH85iEy4UM8cfk4gPWz7xiBCSva65tSZuTnw4
vgtDee8wteERouiZM7MIqdi0NTNJSCEAp/dl4VwXPnkznjVCcN5EBEieqdMm
90BsFDkyP0vUNofeD5n7UKgaZZ3D/XgpyRKTYveyMsXp4GwlLdp9Gilh8Tdb
tmgY8v9qDjedhgmTAnFFxkIjwC1MjjyAeuo9uvM3dUUL9rARRF9RrVcQVAyx
mQnpttAmJUL8bgfPrx/piwQ+aAa4uqqBTzcfKE0kawXAfzczg8Mw+sTYhz7X
IGwDcQPFiaWTAIwmdTzD40bFq8/Ign0lYxhdw+bxctUeYyqzUl94dn4jkUK3
I/cllxK3oH9ssZgDLcMWiTZMy//ndk8lYKpdluL5q8sAkKdWQFXkueHNZboK
pIU4tW+Uwl9mCufSKcgav72rM4mQPfv3OSgacDUmkK7VhyIT70t6ZjqXmjjk
i6uvO2HQQUJBqf5MCETGYDbEFetYa5VwmmzoGa1BUn9KciEMCwW8xomLe+dd
d4W3ZtMStSefUILgpYS9uOTc41Ab5fXIuZorE5OOgjtmuBbMV7RgrltxTwRS
aZEtJcEVNbbiWxu/H61wCnyRny1aRQbBsR8598xR+k6IZeG6RzVpMu9p9Rgk
G3mnq3uqLabNdk6+aoGqja2v0UDOdWl0rkjnQYWyxtIyMNtPej+KSe4VWluV
i8ut+jbyjdCHYqkRN875M6XIBcsHws9sanJgTA+p2VJtCSvJ3PZRg28N8W4Y
0tnyZiZCgw34j8Dj7EzEYOcKwTyedlbevEw6VKvynHBcnqw/PhN98l2wTDVR
YkxJNagiuyMPCzYb+BWBKjlKLtIzm0EuFZGpm9zJmVRKiLFzKXwdGQKaRNev
zi0Wi2uNoVJOzMczeDz0aFVgl6QKgPzg3VpZpSNiQl+FbaMePHeQ21bs9jml
f32kamiSHNDkyB+ZbEoWVpkbM8vlhMz88N7X6nBk995GfBvETVVcf9Ka6ZAc
3/9nERF0zdE7c1O3pj2/ErZB2hpjjPMy/zHeRfYk06GdcePkSeF+QOa7rgQw
7N6XOxWRhnUvVtzcYUR/MLeT09Q53UzxYIqFg41dcmTASDq8uZ/YTesJqoXw
MIbNFMA3DQQcXFXuIJrYMhMhQyw0m64tHFuUQ7AyxvZpZGB5klHkPOkl2kS5
ZcB/9MV6u4Wil8YUvFFp80Qz//U83BjXG+dE6MDNm1PFHeljrJjlBBiaxbuP
vu+af70UQtizBkrGUul/hMTqK5dA7Ie6zprDj3R6lYsvJHIGGncGICIOS+0U
f63NuILBkYpP8hlW6oDBJ6o/pmgSTbYqvLCSKQv6+Is0J2uaw8aQL5q+p1iS
NKEyYVW9LLSiNya9j+usd+C75NNcaNjU/XtT2NZOitUp8GLr2Ho9NAtqIFcV
+xlTnIUc+ASFMD+dbrxNbRKBQhaH03WlFcpuvqzka0QBuFv/TnD8BVranYjD
V/E0ysUSukL/7ihyBdndaMZNGbneOJh8Piq+t//KaIW8pz0XWwuup3CiYfzA
iTX4wjVoo/S3o0x3TIgBeGkZuukpilVNUr96bZzQ860J2HVoH9Ggfvd3A75C
P0vSmJuUPqYXHyxWVR0wgAS0xYj5hV4i+BiVLJmUFMVZGZWIxBVnqNL5ElKS
9NCYWebOzyG2/KfBy0O3lAutzjTb52543q11PCITvhWr4YcZwffYeIwobe7t
0XSwcg/mlZJw9yrq/S2QhYK/uReAUsv9PJEZyck9ZSwcyUEjmQVx4Af2gZoA
gCKNVOk50qhxa36O9F7i+Yw276lcpiOqLQY5SP5n+SFF5cZy115M/s6bPtsF
PjEOI3qv1Fk2lsjn4eoV3VrNBnqm1+qGrntnNzoQaOZ3UC9uBKhy/Ggeq37U
yPWrCCYIrXWt8tXds3gImH76qbaXk2Y3yIHMk/eiMmIDgTAg5Wb3nNBoRLY1
m2Ku13yxr03FJPpWpJQxvpY/CYHo9o+Tr96kx0KaV5U+yuZ3pVl8LI9s4Pg/
FLLqCerk2B0pLImjOAhOhLbUwow6Qy4dWSpKOQ3NzdCP+0GtwYDPRgZk+mjY
fx0Df7DatpvEye2cT285/V+jVAC5z+4KVBxQKpWN/IfH27Y72UwZh3ppMKkJ
k2hhDP4UwQaurD2CpPXfhCnx4zykaBbJ82lEGtXx0Y9XZD9W6mkrn8KlrFgt
i/Ju2COrMOwuk9I8etkINAfW0/g16p2G0kV1DSQ0iSvYlvxUH2c02taOwcDZ
l9oKTePmO9tZYo/63lITR/9po6mcNfLQDfydGR7q2ScnDCOuYdh1zeg2vf8w
RZQkR51cgrR40TQzfi18XCyEV002FUXMAmbTYsd4mhi24wu5P+wYZgdxXZr5
e0Hw5YGyWMJwCp9aEmZhvD9VJNDR8dxNohoUpm2JTLJPtM01/Cbt2xBXllTt
DbvYOSdo3M1aDBZqKSYaGEmWwf4mPrkYxWOGK3U/d6FM+2iHoRqM43mM+CRh
Ivv1IWTGQ9EduuvT1a2e+zJJKBsNsBdhJI6I2WD4M7GZLv7EDQpsomYvDw47
iZREaDC2i+1ex7R9zFZTEbX7ql286/9GFYgA2uHtLny2DRQxcGMKnVFBITlJ
nFkmfWQVKLQJMuNQDRMq7/ehIprK7G1A96DwYtmobJJ1Ldp8v4QrkVQuzblx
aoStgCQ3fed0Eu8Ba6uYa9M7mBn4nTx7ktcsXvKQHrTvx19ARFb3HYunWHmR
Wx11S+VQO2TCizfJzoypDt1lmOgL+4KZCYq8wdxqMnwbXAv0P0BKmxc+PivY
4lBoQJtoTsEtJanrlWG1xneqcZHhMfASVRj9Ffa+n1sngax8UN8gEfjQ3ure
CHJumP2qnYpOcX+oK1LhHB0hO8rhGGrZO6Sn/TezUMuxYNhWqyHwSAeH7RMo
KoP2rkbnal+u/18Pb+6MLrJG5BXs6aXDY+3e6fjrxgTn8MXXWzpYHbzumcN2
g/5TpUKk95DcnPSaSRz2cj/2PEX7BrGcxL1RNXH1I8eoiyKdSzNYfLPvUUG+
Hg30CEB4QhlHeKGAG07eB341B5dIYI9V0b/LjDRcjTJNEngZrvTOD0jZMG12
zhg//iCfnUScUfbfcytL/a07pHMQ1VNu4baqsESwzlnFAHtmy8BLwGp7SeAL
vRz5DDwV3cydfqlOfrc5K33KW+QaqpLGHZ62AVQmvlJ/dxX5KNCb0QfarEdQ
WhNQDvdAjzPQAV37G6YjA0joivii04YmCK5RGWZPfm1KrJy0ZF4GnacmGJoc
CDEt7PtiCsTq/fU6skoydX0KSueCUH9bs0YXLSQXFRaCltWEw0PKsXZ46Rmg
EAt6Lf6x1iCuxQTe14QvAz8Buydr/d5y/TFAoyXFN3lOhlFMwxNfhan6CZEm
4T/5pXYMj0Yzklk+cS/rqhrmh4tKrgxCgeAjcN/AaQc+WocedsCCA8k4k4u0
Z6ag1yJl2iMX1P8SqB295FgkmhIdVrPjshxw4RYEQEETfNCninP2BOPeZBa1
Cyr3sOHZuT182gqArRiy7mhjMDMK17mcvUR/IsoRU6Wrzsu3CFJ1kGX17UN1
tienzXPnJ1ksIJ38IaCtjVODYdzDBti50gKHdpn7lj1HAd6+BLS/owyHfkSI
TQo3b7Jiqj46wEwxlZm1y0Yw5g8vnFBtoeP1n88nVklibx5GQu02hyDy+578
VnRlqsg9qcNrZCGLAx7Iss3DzAB6RmhzvL9SR31xOI0r0IpcPZ7lUE8FZwaa
VTXx7F1CHiNW7z7a1js4OhlwTDTPSPXJV3x/IzfvGYidipHRX5lf4BEDQ3az
lWhz1o9R7i3r6eXdJH9RP3k+eh/xvqaT1a2KenlGAe00MJE13VG0SZOt09y+
EM95n7ve9MOV3/8wBNpVse1cnkp4jxQ5ErORAg5MLpRvQ9k82dPZGtmZ7yNF
t6GDrEhJdkxx1ZCYdGw2a6YnoRFEWMFUeACphO5FIFI+lSxdS4wHg4IxyUFl
ICFcoQJ/gFwxTJWy3K5F+W7036hPXGfyevFbYWst+SUC5vfUxr1FNxbktqxR
QZNWQ1ZHV3e7IgcbMyLT1XCVI+rI+WBw8LucYcpGZ4FBcjspeuHIAJo+H5fF
GrGblN+Bl/RVr5RVgx/k2oaAZHtbv6nxNeFXSSvF76FVgPpvQY/mXLKsR8MF
7So0CRxMMLaw6Uii5h1iF6TgbaWcej1eK+L9Bjn2ghv10dxEf1HLhL6Syw2X
xHQzUoUzcdEuZpB7cF7mw6JrMzEqOLWKVmEYHKOGqcCzpKMcQK33UDUaLKb/
SlId+dQBY7bhNW/eMf97wVenLGAQb7gJ00koAJWFYrR3GZNc8OqY/qfMza60
/Sh7GRtxXJ6jRpRZ52rSrROcVWZJ5gg0w+DMV+TPT1SZlZnSEbXEgQp2kzvd
eltMDWwLtKdqqnYHmClOw+BLx+Gu1r2rrCDndIQAFEgBPpZoDQqu3pfyI8R/
ns3B2kwpSYSCTONp+J5i2CsEnuMr/LAcG0QY06f6U1ZCV5LEXEuKh2LvnhNB
qSRXpLWMYC8fjZkVoUhI/QcUBQgmnwy1EmsUmFvraWMd8Zrb9TBJwu8s2GMt
5BbhLZEz1GnaYC2xPK/RKuzm6TNR3Z1FCzP6+kKkAEDxurAcLui0DwjGFaGu
G9ds5hJHMclKAFCV9SRY8IgZDujyOfqXkG6/zXbnNFKt6kVI/wY654NA1PQq
7bjjbWym+35m0poNQY454aB/3etCx2BpZ6mrUd6dOZub9yvgdECGgoyWhqyv
qfNcWmRub0WCdir0OCpv/W3ur5xN/4sTdLBiUX4tvXpHchayuVvcNYVHefGt
d0R6mHcbCu7nhuzLkfXIISqJGdn8V2WKA96KAYEB7h6dU9wSnljWNOB1HZ2y
QCBoJwOterwr8HYrYLIEKSmosNukQ/299ZvPCQXDJEPkHSeTR3+QNwXp4ozs
jR2pfxAwdrdHuhLM+QPZ/m881Tj6fvaMUDK0filwYWlHy4fd1HnJg/dRkH9L
Z7lVnPnED1mZXytRzrnpWMlG29P0EZQ/KEzNmrbR10bWzGqYuo9edYod1o6C
TibnxahKoBD03RmUfgnUei/lH/XG/ArimskN1kkVk4RMA70KOROb1VXDUvMT
qgKMfIOU3Mt2IqZrmThSLyUGtw3/Z8OMkXFNjA2HvxUZcRLGfHJlccdS+shT
L4yQG71QELhCqvTveHCRiFHnSA9ggCsNKK0tUxAih4VecTQHoUSBNblCLK9W
FsCVwVTC8XdJeZKhVCXbviC+1Ndx/Rug0oyeyjzOnv2ksKVwotbD7SNpNWMA
3N4nicqNdvrZYoym9doPv4t3LhkyKtgTQZa5YU6rJOU6gCzClhyTw1xm5VbV
8LQarDDiwszm4JtuzaL/tVkHf9OWS3ksoGFaz5gt6k6dGvH5OUvS7wvQi0Rt
HvpwNfpGWSDZ9kcYaTBZzdFsWCUvqdvoLo9+Xag38ZVMPlBb+gl9hTnvljeX
LMMMmB21UTSUCve6kOKz7IprPy39efbIyN35ERBVBa8I3xTFxPNRukVw3h8N
1wRm4mhX+g59UJiBERMd3aiil+Q4I5kpvd/11lnPafBvU9DZG4UJSjZYw813
SFjSoKXwnp5qFNkAUjtWggjRz8llOS3UEFSrmqcvNJGtZE6yFlN1Ed3SWQqq
ugz2Lgo5uJEsG9DiadfrR33dvsMa0ccsJY0I/krkOkl1+VQoJwHFS3IKOYlr
wKGnPBlRsabBDyZ8126MBtkSJaQoT2+XWUIHFV2BFVClO05WJYanFfhl8S+g
QSHAH8BM4S7tzWC04Gawo3lf58SoKQlboRh+lzzUMJUEA//LCW8K5Z3ddJtW
I1lsJAUMUH61FKBw+kg979adsX7EXByM/UCGPs8sEzkA6jhvObiYqRlwyGKO
bF1kICHf8yuwDxQ0ojmloCWYnhQwl2vayEycLgojHXX8xv9NRlXscei0olbH
h7QQmZA01rq1cit7U7vwq0qr9WvwUqqOChcewEasLdQZHlKCjlM6wwev+F0J
GmvOik/jgeFEii3f2t6ZjsKfnAzC4mgc5DzUUam0urGWuNZX6wClQxmgtaNI
cADxoJROUfOKcAZL5ra3WmKV9r5KpPHEecejTzyolXxPJybZyKL2wjnXaG+8
0C+gpKJ52YpnnPC9Zv9vByRgw6hKEYOw5IIRJGEfXti2+utPeHa/gr4PRoqX
BVov4zgONYldJckDla2AVnR3dL1HknWGC2TVNYBNC4Kc7HPjeW5wquzyD0tE
PU/DYj3OU1n9sYPFzdAWy9zIywNMa/Qmaoa0BctxCYCApagaJYj9lwtdyiNC
xbj2sJU+paN9JwwzNPw6ln3kKYtXqopeLIHkipIrhZrOlrpRjXLkQp6r2L9V
NmcP6AIadoxYk13y8VUtoNNxtl7VYHslnmdyVpJu/dB77eByJ2yFD/zFXFsX
dpdIgQNtHbpEkFy6VolEwzYky1FmZ/WcRp2hpaK5i1euVnNGQJTAG/aAxEnp
pY9Tf+zxdIrl9icxiYniA9VOmRRuhryaarFEQkfmkGjWehRpc9Z9Xb+rFYVI
wJDjsC4lFuWbCf0gnYHo084ILVOX2NHvcQq2WR8BuqPYhviQlcRburLFnCUZ
Bk8B9236eLOCm5qpPnDf9pBNaqChV+EA4d12Kg9PNCNXFqybS8kF6aHbS57L
ERHMQmnwqjIIpKwHeOsJnePyRETay0I9UemErwYmvUdZbacQV9gNjjCEwd88
wBIA5Zfstg0gGb7kaVYCrgxKCbh/HuTcLnl6RZ95JMK2/Jc2n1reI+iEIjva
w0cIgOZi8bInRwWYFPU4bEKGecjK+Q+klv7y5CFsD+lboBtNpIN0wbpcvzgo
JIOmtZYb+U1yyL5L/airIB65tNaoMj7KggKhSlhTDEM7TVfJ7yP9sJ5PyOIb
kXDujZdUrcqEsX/MOa8vM27UHkyLecKhP2OAyq0C3foc+8h/LltZEyD6sMtl
jTJaUE7z0FgAi70mHR4+jntTtpP4hWp6bm3dPvEne2K2OdsrUoVKQf3in66b
ddoORKnhqME2cteEW6WWV7rQHM4mMRyjAdGtr9Fe9Kdhwuyf4cjqhM6PQSg+
Y0/fDXMK7JnQzQiCjafnrSUSWuFo/7AI9rbp1biHZ6Uglfnv7MboRaMWua6j
6H1z3MqhDwldbYGiko8L41kIj4gfbX2EqtumIg7fqezjIqa+Ox78ak/wM9gA
lK8AtF1CynZDOowIlw/dXz+pwGgBzLnqfg/HisVSphmplE5gzTEogFsq2UTT
6o10wCfNuy6YTVmwq8znbX8K7swe/2wi9IzEDmZaaSPD8cb8nQvPUWBRjgyA
cOR9U2k7FUZTsLbjmzzRFWDsM4azvFug93ubNs5spISeIKPGWlJuJdVKkR8d
z1awQCEWEphxxuwD68vggyA69kY6cPw1IxgU2khPzBoTqvt2zePqv32pWHX5
W0QGGbUktoxfKgUFMQREqh9M+bKgcWA5lpgwsQw+yj+cKwuJGD+ZQeZ39mn+
J7qh0bI6RQtOYjb8WmANNP6v2mY74h+Dh52IVycflbfKNKyPGPt+gA3Jzg9j
tejQn7bc6POUUpcM1icaMa1WBq7WulLBe1LN89Mv1TlDk1/N8d0OrlPd00fV
87bVM413RsiwOEihTcj586It4rrC+OQ7WFdDu0vJDL6R47izzqbLRIxQ7N2o
vNL1VZtT0hWKoYaFOzjyv7U4EMcu4zKo0FJrN7/9jZRIbQwDvQIJ9XLdyQEa
IdPtr4pPA8sToVBdz1SewzOd239ygas7kfaWl3PX7EzLHtX7uwVDl75aPiH9
GRS11ZtxtngPOBC35HSJgh1zRY4Mcr9KCzTuvcf/oBOsI4bFhgRb+NoGnqsp
uxwvVyJtRF2ckGYn6fLcdMBqvYPa1dFL1kkVN+YxCINTzf/+AT/gBww0WmTd
DEgooalEhGCpBYnOBUdjTSUqIjfmWdeDCshBk87x3nb7RwSWumUbU7meL0nR
HDJTCJGV4ZyxdUGlAPUn3Fs3Itsjo1iPGKcyWP1Zj/VzHH2dSR90mXc4NiE3
O2iS+mfjtJywlE83IpWaUEBIHBWipIOcNWU4PiNLRUu/pKq0Hclzopxmxksg
t1K51X6EXx5EK8Ye9KqmsObUaGg2TTWCPsrMJNhZmYHtXL14/8WLz6XCcucb
up5I+A8q2lEXFTzuOB1eEGLE1NIGqPYGmlvalItY+FtrM6WyVJq4AZiLlU+c
XZYVxRUAFbWVjRoZ1AqDkZi+dnOvXg+/TiHSb2SlJqw5cjJqDMMe0kzpgpdH
eP8vOrOqKq78eOHrRluZ+p0RfhfHTWZYn03D1Dqch9nmz2qFqcWB9iWUmNlW
c7Nuqs2w+emiYk6ScLICtEpj2sUmiroi1zRSDoQCLjRH9RpuS6Tty5EJwt/d
j8gdaoceRpbR952XHIg1mhZECchmwu1h0pjUxeNpoYsM4CS+Fwuo4EvZvtyQ
oSW4UbjdkA+e4emO8HaAQVcEhJhQRwAHoptuRGqI6oVdeTazMNzo8xFeTrlf
N3flzFs9taEL/5vQ2n78WhHtBZSjGmCEGyJmEnnBf0St6qCH8XH6w8LpeB7t
JqDDt7LkLefnqSszaEqGcuPorTEZy/aMW7jsfbQ8cbAIFJ9W/dhRibvBFhh5
X5FSNOGpPItPafs3HAiDhU9E2kZi/YIMBHBR9/AT9RMvNxj7M0rGi2HX8381
klV8Cj8hbm6TGVX3Qwsgc008orym2P9wT5mQstz5dOaVffGFFokNKXIk8Vsk
fJd3aapTPJq49LPPqcqKxMj9IfH9wrVsz1cPYPdLDY5tRGPnYJKoINIbfKc8
KsI0+rgev9Jn2fLo2a3l983oN8Gn1IuZzRfbouLP5b8qP1uynPSk8ZNzGFTb
DdKEV5WDwFOPzZcNqvnUSmrYmjz7shhU+HaE3VI5C208f3/eZ2kZHxc1Liq4
p1Q3BVMyiKrdW7bwqw+rMVOTEe5cTo/ebIXJCXWPcdYX2VBqj1KPI8x6cVwE
Ry0Qlm6ff+COZdthimRyETUm5Kk0B70tsHKPdNhTUFFMjzDumhc4fVOePECh
ODw9uuc1BD5lWa0NKcBuJG8al4WU9csVDGtkUAmLYBquZWdIz62BIQCxNaCr
75c9CvMFen2sNsHzji1IBfsZp0m64AhIsj4UvPRpECe/D45KKHAILXI0e+Jl
jCklpxA8O0JlQiz/V1on8b7zXiGPa8v/KS+yq5tiwU+2Th9A/dqkBlRDPuuU
nGK/i37VMa+Oi0fg5aouWCp69fbt5KAgrny66kTQfIzMYvrbh197NA5NKIul
+fQ+kvaNjp1XKNDKrZCOaimy2/gPBD051xr1TLGsVVZttaXHQcB4BcsqVlvh
6W2BHexGUu//niKdn/mOWGbMMgGhcxfABZqnZ5VRRj9zFwtE5vCZ82KlEUdJ
sTcFn8VK5LgYxqqUKcFCxwhqg9xHez+JotSN1QCC0k/h5P94yB5sibe/Ta4G
7v1FDwRbpgM3kyHXK+obSoQ+y/pp/pFb63YROki7c++ANfgg+NH4PqvNJT92
wR0E72wfKEQLR5Kc3Vo2TKIbVXZEdeJSHXMmBmkuX1fgGIYvlzSMiUJiNm3L
Dpus3A3IbC/uryeCVW0w7pdH5tSs99W4+uNHr/Kc6BSAKueVL0cNqcMSCAXf
vg5y1KCA0gP1fVH2jWkWQSO9E4HInruDiU//GgA9t2duDMI8oTktflJmFrJT
0/oXf/nHYGTzbtmTRiXdTvg3wjoN5nGp6i72Zn0aSL9akpkPp/K8Crb01bW+
OZK4nJo4yZ8hXk5wcV5fDnG0a66i0FfV7YmYr5wf4mhLPtGPx+IwD+fQmOg7
4KhYa4+iC72pksxhx3cI9UEiVQ+VNyhjxVMo7CMm86wTm9eufiSygAP8UOJQ
n83i2BnEn/usDcET82JZraMEupDnBmC3ml1kG0z7MbNhateARRSPeoPqk5Iu
BXH3ed47cNhiTkLtNLJmHS9f6UfvdAMH3NSn5xMqbPnHqnRilDoiBKeMfIwX
X3LOz4LhxFVS7RX2DrD6HT4FKsnK/hOtiBsCL9Amk1+JX1Zn7If6R1eYD5nB
sL8Ll9Zw965WdKCsZjaWRcPq+T6HiFnGxeGhiGCYZWwGdu1PHD01iuAIPDtW
cyeWgc5sNpjAvTmI/mFpLaKobJ6WnurK5cD9Ww0uOk+SIDntRVycxV8RVGue
20vyO9R7O/i3+Dnus/R5c18AMiyVU2zZwACP06hUpYMTebfWJWMPsFAvnHrs
vKPFKajpEQwxNuMQ4hChsC1p7H6Yh97fm82LBZsT04inhkAPqhXBTufMQfpT
/R6G0+JFKelz+kVkV9sj2n4mqV2D/CmdNGpkOC0VGve2uc+LVSlJl9s2kbsy
l8X3LOmsOhjCyCcXIwXzjQsnQO7mxx6BGy/38ILqAvUzbPW0BVI31QxR1WTt
lpRlDYXIsehe2z8lhTXa5UQrN8RPdLkPHLzkzz8/JQQUrIic/9Ilct73+Mdj
VVJRi/iBlhT3BIoGXbF8KqlxWja2RjVHkRjE7b/1iuFvWaImqfMNMz9KpDtI
hn7veh5AmUqj/ggFDa3bYkVb0EeU3ylLpj53dwmnrhLnmOd8+6CBJ3aSD7lL
sZzwdYy1rKIa/SzNcVx3OQZj5SIdH81PnGjRA5y3IjTk03Nf7ByQc6+I8Daj
2T9sc0tHDUHvvu1MtI5U7ZS66fVdRBF3Em8JTCyT+W3ycqGjgr2+scAran4a
gXH+D7c3ix1aMGKelUg0c12nxGFmN33IVDwdDrr0m3cPdgQU1hGwNk4d5DZe
5tHCdQ54GbPYdER/bWyKdVionQl9Xtb5eBj5Dutb/wrjvupIHDmx5gFsz4qW
WMyh01LlP+5t96MqA+rzOrcDx6kI11zP5Erhk6ynOTTMgws5FS1hJzILO9+i
CXhW8Ij1+SsnjG4kBtvv+DtI76jVofEy9eAHI2f7OaJ7UGPiWerHy/BulShE
UrdeCA+0SvTtunFmQMU8lkJU1JRtwHvcL+o9IwUF76m9XskdK0X94TVm0iiT
pzqJpTi8zVnR9TsWOMpLiUK4M55zI0q0wc0I25UY9gNT4FmzwRj++HNMm8MT
WTqMuxph7ER20c3+dUFLosDXl+aBPGwgcblAg4JymE9L30tVTXcxLMBxQwfF
+6NXWz2VFG3b+BqaumI1SBclSpw6mqcadd1Qq4WP7DmKcxpP3+0b+OYj5WZI
shC7tpDLoopejz/uYzj0IxtnBqlgxS4mtc6H/GjFz+8ahrZcLsHi3pgc45Y3
0/V4kVdMLEv9q58DVua0/hNDlBuHWAMAHp1gpw/JhibxvsXtXLlB/J7E8qqX
8P/aCz0PT/IhKYvR90VTX0eR6jSVX8S/8A1uXbqHQFh9rQAAlzFtnW+jgZiL
H9jGbJHg459/b8TlUs3+1dkSPA0IcQsjiSTYYcwdblMU6SLkIGQDHY9j9eHZ
4JZ7CL0YB8Ou9EnzzIVVuQ2B2s8DW1RoqbKslfAh561TzrAhxX9RlSvZv/4c
KATfrM7ili31kM3lpm3GWa63LZdfkWdrTEOBCr/XCF2xKGKz/Rj8I1NejFzK
BRbSy4xxbXci0Fp091tTxe4rtgO48ea07dbdYQLdTVIKGdSIGeASo2RFSK04
mPqLFza5SDcOS0jVDkhjC2zOCdviF9om0oqy61NuUa5iEDXki9B6ykIzGyTU
qZw7M6+Xm/+dSqf4W/UgzgTHZ+p7h+LRNIfI4j2gb/shb22WAmg+RdNgORxg
5v5bkiPjC/3WHkq8qSb0WKKdR7T8Hd5vS2ZxkoUx+BoQa02UImxbErgfZPzD
0g3BA0CUbV/nobvAqOyCyo6GPbkE0rJi5RW+uTWE9oK7eDPtGkDSFHRz0Gtf
TF4p5hDw0WCcN+L8gIFEhq75HSi+CPGF95O+bYS0votT5KWSEDLqdSeHhXR0
LMQUL+1hFD+tSDCHixtV1XIwO98w7Y/v1leP9xEiJdigVI8T7IfxZJZTPL2s
MFUVi5mWoDzUa+ZQa0NykeEKALRNKFdsktaexNjvmnp5+5zRVknm8mnj9ipj
1juZTN/Yt25wmrYaXwooboL5OMuZ3Zt6wgGadt+e2faZTXvDLNA8lXoK9EwK
zrve3dWrp2454Z/Rn/eS+y2Q6uHU8Zw8c9f6cO6ikMBWvDDjgKDtx67WAzLE
9BsbfxBRx+Vxgf5NYIHLhh3vSjC3Y7oVQOok8vQXB+vOZFtclIDCGMN4mY+D
OdawwLSziTAwvGXiYF9ANXdtpT0m/UUsF2vpYuXIf/y8H+ZnX+Fa7d+clgR7
FAiSBaNRfFVR2gcfmcWCT+tUt0DFAeWZ0Ctl4vjq5OU1hs+LVLt/tbyA6alH
HsPC9TgfT4bNi4S3nkdRMu68bsr1gJfDKOC/zErIki+iFdRuwevmlGAl1+mO
909targgvBpvhlazcJPX2JItxI8/LcC1ex2xtl4vNic8HafRTNUi9o38Uf2m
ZH068OrnFnzHHBnrenbBUBNd5AkvMkkES9QZ8BD871uiiSfbPQkcpvnVRsEh
PBkk5/zssfb6j+RqH5uTdGkVs4ysJLWHzOIUl+hbI1boMNBzGBt+Owau5FKb
UxDi1LzsF6CxM5A4rdT/puDhZmdpdmVM9UPh72lQN9i6ylKVI15udeXJiYk0
LzynFSU/DDAfrJK4pu4wafs4BNmFeSotnz2GDi/UCFGjDbdCnrRDM3z3bb/T
OviowE/sihoNiIyPisAMN+1tEMUIcIfZHGWPsslDA7kT3VnXX/k/19KRghen
kplPX+fwBrFYjzjaa/KsB46P/vlOdlEIYh+EERQWdJgPRXU27bax1+xzPxxL
3oqLyOvCN8kOyMp9zG/iSdo2E0l3mwTmPzY/YOL3yb+FJrU3OhFfoew9zTgP
vdmHM7nDioYQieSGsz+pqHMFvuNKFC/BKmnfDlQ3NIb9ArehfwZyvtm/kz9U
+3Esh8Coi7c4PelFWp9UiIu/j+aUrrRj+fTAHvmnHLRVC6FP/Kb83RPaYkyU
Yy/KVt8q0/XZy43vguotrlbsRKnDZGiw0bp0c5XvcYP2ZXDmfV2IL1BcnL3l
sKDqzZtiGbk6oSeBQiowTE9mOsxEnHO+3CC2IWhqNbR/ATTOqBF3ThgEM0HW
HcR0vMKqMe1Qo6HYBSUlBBPajWL1F5mRE90FMboscmi2GQEQBIFErl2oR2P8
tEubJyLLFyiSWerMuNBs6Ia7L9NkmdvjM0yhKXlflL7BNetPWLyAv6lGdi6k
FiE+R04bKQoJkLkabckI8VKn5Y1gSSXmxj630dNB29TbZdOoeyhi08VLNy1h
MiHa4VJmUKHI9IQDW1i9vr/eLeKsPdasOTn/QEJOCSUHBqkMiisYxh/3VC4s
bot896DFVBQpmF7r8dontaiUaMDMp24sXJ+6roKr4KXiGfasGsZU589QbE7Z
7SDZwQ2y7pIZpeK6n1cCpsN4oFtgt7XvvuzFQWwJUnv/bPu+nwtoPqJtcbbu
n3Rd6kY2ppXdzEpMRn/DqQ++ykVpzKl98UnGjivKzjBjjqzEI/ObunulFgxp
h1/kNjy88DgBkYxg7MuH7kl4rap90UOYPA5wvkqv74inX29j2BuuvUxuh4TO
KSUoWmKJGkDOSdRR746U+PKTGgmxJPHaWXrxeriGBbYymHMnvBALuFsF8/AL
o5dEY/k7V6LwzXQid9FHvppFmPP1xaFwCnzb6vXf5yH0faRLjvbNdNW1EUaM
AxM3Cn7TLfQ89f334/f84OHqeHiL5b3IoT6dV6UVA/80pKo2zhYmYKvyJ8As
2NtjRAyrW0suUESmW+8e3y4+LvNXPJTrwDBmA5ZAWRgzd9l1x3kd5IV1k98C
D3wsFih5uox3XDH3kqXIV5lHT9/IC5ec8GnMEiaRq5Y+sQY8ZNsP5DGNf3x4
kBe3zqteu/8sU3FGEVSeX+V2YOZetgISo3Qi98VtIjOj9HbEVY9PY5kQEKeu
mFCRxsJi3rD++IbdH6P7HlWIHA6OnS//MM672lWFX/kF0/3McQ6p096q6a9j
U4NqbRgdvI+BhOOhnDPkCyCkPzW/lujHu+dGRN2Rp3XBrpqi+6+vp2dH5UDK
bK5Dd1SFpfLgqEiar/qkSmgISIHH3mhl2qedeTU35Fja/Tg9xvsMgchOqsW4
HtsZfXCdtltEIvvu+RSiIdGxD7TXOyIj2wG4AP9a0Zn7KVwEDR6naUsjJe3i
saSjQpKowndiSmSnFZo4SjqkhKKePNbqaQV+retkIJ/BTo1spmh/+gdlBJrW
f7jLjvnbSLr/YfRY3lBXFFeCyRrgrKU+zienhL/Gq24k5Oph3Ck/ymYA/l1x
ao1OZgK+V1Ukm+uJGxh5cPKu+GfeAJqHN8MNZlSqmhqpabBUHMA1CFJLiOPJ
PPywoSkuPJi4IFGS6uAXilXPlj/QroYpiVmZvEQ/n/f90M9d0Y5omJ2yLZH6
gGDDGbtmWd4Nxg9FK82QmYtnjoqA3wcUARkt6no6VnliGFeWM5enK1NyRXk6
7jIdhsKcZ8mMbEXWDOxZVphcxlUM/CfADa6OpvJMpEYWGXdFdNp/jeHeogl4
dUc9DZuT9/26biSQeZhU460MEulQmFYVV/Y2bU9TbMQL4LbMw+CwEYgi+wQ1
zY/xCsqHDwd1sn+Nt0rI7Bo1r3rm4jRLv2ytK8FHQ3QvWo6ydnTZGqNh5Dkf
Mu2Gbn6NnsLdFonzd7RgVRduZmc1XwOI02bLouqv62HgJTOXrbFQtU2iqL8R
L0R7K+ZxF2vpk9/KBy1LMVd40ifZw9AK2AtBk1a1K/S8aiVBFXdUgnEeqJh1
IZPqYrKBFwEvV/bHe77pmLT+142GIekhFNU/vA6kuHtbAj7rabg50HLZDac8
4qwFHHVh3G/Tma4uZD4INveJSyWBIeY2ugAY33v1cHmOn2aoIkfNvYfpDaQY
sFC2Aa9R/bhSN3aqV2XzyA2lPHpsAOyoqXMTGmCbc5I2hoJ7m2au6NwxcXYD
6w2CJs83lj8Cuni7sJWsev8ItjnXspIkQpEHbZygift6Qb/2SPEk8WuqZfPV
R6Fi4+QpVbF5D6K1tVWOIeqog0FZVtQSgxAT5NBtdNUlsTnQv9htvKoK0bEu
DQbaBMVFdC6VrMrKFglDecR3hL02B+nYTno81HYrIudM0+snov/2gzE03n7p
FTQRovXtcVyn/w0yeiT4WDJx6NhdfLR7490KXubtTlhEf+LopMbheeZCcwOl
wbfIILfJk0OPhLR2ml2YOUzztT+k4I2K0r2Qhh+fUr5bWiTzEvb2B62HtIv1
3o4VMOueoYOXq0ptVdKX0lbYn8osxOJoigjM4pc8ydxHkL7zYY99bQhfJ7Vf
FbQ3q65zN+awY0tRP4TZ8pZdGbfY2tB5PtQ2YTmEUPYGTq0Fu+R7Kzc1Z/Tn
Iq4ZT9dSVKtlVk7jt2RTi9d+MFpPMwxn3nBWTwjm17Y9wlIM52fARW+vMK2g
h6pMMLFiVmF2+UvHOGNriXS5V4kbKaXlrog8zcK9jDDtcdSLq3yxUVv0yDRy
uHGhkGI6JrXp/pkg+yzxI8xH6DFRmdF2MThtjL2ITLA2bGDsH0sb3GRbUsZe
WJGkxjbyoDcJCcvHArposWQXTI+B1XAFh7fd1Tu7rP7mnGo+LoX1+N9lhaXv
NKklODsTrdGhrfws1r/8+FCbT+/rUXRnzr1JO149KQBMxuAPT2TbNpIlBPa9
pBCPeL47sJVfO6zblt7W8+TBJdWtymrqAk5/RwqN5J2p1YvGjBSJ4qPtwJ92
9dVzhNum+VYJ1pYpPIMzfFeoKIazennEtKG5qhqxTlpt80l7EJ0hBtASKoUt
aCouXb7aSTUuSwaDfwV8hHvPrT7ckQwP7IQK09r9qA1bwV8QBaFZHO7tfZud
XK8QZD63FJvVFw78D2BAcGuEuI1WpDFevhtYhlkDYU1xec4QKRwgvOwPB7l0
g/KwWG0HEAyg+ew802etDphZBFmql3jNHKhRcrt900/K0Hi2FjzyKOyZTlvz
0RakxqpNQ+3X4l5TzMo9ZfLNx/w8x+cRgWbLoIcGBr9QUUjz/haTXGilZUj4
sWge7KtHK8CRHquPg0xeUuF98HzlIlR9d6XLsCERNyFaPkhifl+d0n/W7mrr
IYi6XRmusCBOCDCB8jDEftHKsMHfEC8PNuOzl5bBt992X/3hgYifkj4wc4I9
IbeFJ93zuUocuOJlosWGP0LpIAKrVugdI1RkkFLAg9zLZvUB4lznuUD2lyBB
gI5FhSDiaF7KWTUONe7CxlelT8ZIh/VqX4oTZ0Et2X5KVUdb7s3t9gvq/hml
h/S+MUbxL4KpoB7TsYjyTbyG1OE0b12w8Ixhv4lJYD6XJJfUoQv3DhxR7mS0
XIe4GTKj/vb53s9BVZGe2nFhBEzDSigDpIY7dV9+Xy9fAnZ5G9MBJFodvc6b
SGm0s56r9kfM4sidhlqVbcJ0EXbx7z8JSBJHzSX7f3XNtpfr42NNJJV7PMyZ
cRPY0xtnE+b1C0p3Zg7NpDICSOBILqlu0ShcmImVhiImOqdFHxND78Di/j2b
c+1TX3RNRaCE+YdMphJE7z5uAMor5+kbUbAERBRJnTJrzUHt0uGrFl6espyq
ideSOe78Wsm01GlILzD55jDV/A75vYKYImKgGvon9r+0ftPQaldjJKQrIBUR
Oyd/2jLiJ6bML2/WaMKjI0KxYxA3fhnrKIh9/0VdDuq3YLTNMKQ4s1Oya71D
hQiScy/kNz65Vq8mbHNNWOHmvEDB3tEcHNHLTVFVn9AbZNy7iHx6GDOuoqVk
lqRtQ3hUryUuHTj0i8WqO4XNhr5DdbmE5g/t0fMtSKXNS0IgB4nQzgmG4o5T
J8OzXDgdMUZOxy3UrZ57iKBSGBnVkP9An53UoT36AHuzA7XYaoEaBaYf67h1
lb48c7G5OxmuqgBk6wjnHmprTl1KRlbEc8AD5ibtg+qHPRRgweX0Z2QS5UA3
vyNi5lkPFgd3yxEmg2D66bv86LY6Wj420loY609eeOGgpLCos40rtzVVVNJD
tsaSY87unxRyepNzuK7BNf+NmS44WIp8loIC5/6uaj7QiAkyz145DaMe+Yhw
v1hX3qiK0eaNs0EOHgvDRBbp/EhxQbaOBLdot1IzHQe66eRMYGm1uUZYlllJ
83QsUTIIDShIJYBOojf5OyaY92i8uW7wg09VkmEHUSFsCJRVGsJGh/xbs3Yz
rv+F8ms5q6iHA3eZ+k1a27V5eGD6ae98aJ6eh2A7ZqtKUoG60E24l0mI4dQU
1oZyHyvtP0ZFS6O/GLNyjHXlcbJBwIx36hMXo2ECNlssietgyozmajTYi5uT
PD76RxzgFG3RxcP7jTJvxBGK9dsSfUZZ7fsuh+6WySAWhvds2azIIg2u8M1D
eSOs40dav4mN9Fjj2UD3fOuis11cPu8IbSvbSdz05rWSKpB9sEOw3uH1oXqV
GSTRN9d8snV5OPlbp7X4YO8kxIlN6viWstFJxeEBK3kBvz1BrKFicwvs/wT6
jbnfS7r3o2wES+YGi7erDkOew3UF6h07oIJn2qChUUHD7E2eATmEoFQg/VbE
Dtadw6sjAnXHGT15/BEC9Zyxrr6nu3ogGkohnKhcCi+ymEsFJtIu//H/DnPr
L9kURKAwI2ayJFtbunflmUb9uQz7KbBtuVrePjDPPQJZKyKXZWoLdBs/OIWI
kGJsksRzK1cPDxenPYoXOVUlRbXFfrkb163EmIr8L0aV5zvYQkHvusI6TfeL
8wru8G4wqZckeEuPy2rUAiM+rvJc952N0QBhnYd28aJB4MisQ5wvKHJob/GK
Nr63Kjxl4FdpfYKSrQlj/1mYjV9R+Q2lwHf447pHEQKtEVn5JLAEaLxNzb+6
JhgHroDnYMLgmdA3flXdNllQZVCefKWTEdPOK2ai7kXsk99I+CY7EHxjig9F
ZzqvRXJz9gkFh5ZjmTWgwE1n+hkrx2ed5Wwi33YPXnnqhj7eu7AVxwKNLK4u
GQQR/Y2TztNfDvnhtkTKMX8nXb9szqy23jSAgDGp1Iw9zr1angR64STBWHWm
yY/QEHABWb5x+LiHfpnR3fGjesizxaKFH532T5J6EstEEGCXf6viWiVvS2hK
1K6LuF8+IkBDhdZWtRecmGscYtysMtVkz5/eOX4vQ6hsjj63t8j+vkLuZWsj
+CdgKTIiqhjN5FB9wz+BQhVAIZgFTzj7kBywIJ9anGNWXCNFtJ1Z1kJVAA6E
4oMiT1N6r/8HLvVsGNIMwr0PxvYa+DkMKuAdixu7nQl1wfTKLnEDeFG2jrWA
EQSyAPeyfB9sViqlyOrXdkC10xv9fVZ52jfH9iOQR3d1j58GDzjH8pNQotfj
yce9056ZCgZRL1tLo0eudi/ScVQOnQG5wH8LGnvpB00Cq5v9QyzDClBBAAZP
Dc1MoTro18aAN6OSxXdnDQpFGV8ue+m9thPihnfyen44DsJu7Gh+tx3dVAnT
8v3mGllajo515MFMww3DBY44FHXQonwuneT61nkBcF0n4Fg2g8G7RAm4NtCD
XARfNZ6GxtUayYWAnQkmfhubqAF2KXgA9oMRNGqoXOWzJHob5u7e2vDHLS22
wMf0qb2Pn++MvlKGYipxYNF2SO1tba9F6Z51KRhVEO8DieU85E4Cw6dLM51n
+TqRHeUDdNKTjLzl4wrjRsUdrepyymaHyMvpljgF0g88zGiOy6kC0vvFJapq
j7rnF/B2ClLSWPrCWM4tS8kbPHwoZDcwMoe1BSwfaz8MM3sednOzAmQFTEou
uzDjGlvdBC6sckwI7JxCuAK7vQWlLtnjpNw4SyLMjALRIhVGPO4Ww4OO6huP
4mZPKsbs6FQzZBzq1/55T6krJPdxaMk2LdsC0088dBU77e/7trDgpsUa5UcN
RaN63sW4BR17et5kVmvxosR1tBg5W+8ZlW2GW6G5+NCYhwJmtPURO22pwZY6
oca+cJxvWqSm3Xyi2zQI0CpwmDL13kRmHFuPLLGi4ifmcoB5mUNey6WL3F42
xvyWl0SJuke+xbxULkjcRlQ0W3Osnecp6BpqxKrDo1W+G3a/lx+O4cT/4/Nm
PzFfBdon+6us+LnCOr5vwa3R/C2BiNqEh0lspjJJbb3rI6MsPkTx7c/l6G+v
4UpJ073L8YBBjod3UJDWHj0dYDHFdgEwvir5O8UX53jaPySV+SkKdVhYvBEq
kkIk8BMVDDdX5q45WsylOPTXEzxQdit5z/mUmDRUGW6zBN4JSRm50mnsfVnG
dY1SqAGrkEnmZAt1CmgES12y6Uf3JDQDNzPVUaQInM1j57zr5Fxwhm7Tlqfz
qnUZ4HSa5t7sWEVO4GaMv3DmbgrD2LRx1yWNqjzVHgrPqHEEKs3iB72R+jgM
HP+6fvjPQXybV38KIcIzDakP9ryC0yNrXWdeTpQ1qR0x9TF5EIol7xezvkPK
d/NRAuKxQxHanaluzTtOnXCJyR1vTZs7BtrU8gW9xKRP7Zgpawwvtw3bnyzn
ECDiSs3DJ/ANmRtbvNgz0g3KWQiSemrQeMbzXpn48bGaddqsa7tNJQvQs6SX
BMiZz9gTsEi2bLedmEFmxVkcWzoVTXf38glRB+gyjruTKOKibVYGt1kkg8xb
/0AqPCSD235p82AhlI85ev2Y1D40jLvTTsut4e+dBdnPSV3y5YweJdp6kJkZ
aBo7Djwrbs6nslwL/y0Cb1aJzQrOOns3PbxxarG7uIi43JSKta4ELAcj+RdD
PAN5sV3uE+r0QfrVwf8SWtRo9jKhHdeh/Bfp2F2JKtdbiWE7KdloqVujUtWY
5kRCsQ4t/cdbpLKNbvUwo/gi7pFEM5a2ExGkHsBm4Qt1vDI5qtoZHZSFCoin
w2a4e0SfE2C/giaxq6dZx1IEFVVhsBLmOoOQNU1iaMqheW8YqDwIiwm8kS/t
KtFHtBAkM6FFKPjUehmcKU94fG6+lgz8IC0acj5rgzc+l0gMrZhil0lRB6Di
LUUzAEg3N3YPdMLfu3PuU4YMGK9UvCgqRSx7zyipbd0cvZedBSlWvo6jkSuw
4HrM5r9kcm32ykhzC5g9vAaf20bqFsn2IthbcUCfx+BgjNfh4V/xtpPXPrDR
YGollWrxN5s00ikMbOGHYCM87BvqpYMByBA9Y8PelJYgChErUCuz/8chouo/
kLJxbQlMBRmiO5rejjorTXeLeabGWIBTQMp5CG9XRoAhOOtYKOiT7JeJ43ts
HSX3Afe9M8/P0DdFPBVwJZdliyR6aqywyC3IY5lzV35rjuC4JM1hFMe6NjAA
JPYlnRBCIk9P5v+jH8WIY0WaXOOgN3sPVI1OL/shH4p9PvRTTmt3OJXE5jrf
7wR8GfNwdJLeans7Ka/xWUe6/AWMSh9K1Ij96bz75ouwGbk06kbz55ovS+WN
wz4YeeYZ0AseoQXFpywiOmSNPLQEIm44+tyCmpimNQ+Bz3jB0s4n8F9h9pr/
7cQ6OkhXNel3xUIlQ4tgwSd8cEIR+4cdRjd8An/GE7pDv0TBlV4yABjROuOd
89qq72D5gDe02x/Ig+py7ZAFBACGfh3Scf8LDNr2fITkYHpS53yf8IsltHRK
I5pmGsJUQRncvEJdKdqik2DO0C4HFZ2GvvcWu+Cd/TT2/b2/qgPrjBUD+Olr
meT/o3lI7Y6xqS3ML6VJICY9mN4XI+v1GGwK0oOIpQegvvLU4gUqHD8Q0vXW
XNb5DvzI580p9dbEYx/3yqtyr5zFjjzBdZdM4SLKGIYMNO2bKUqBqPBAIHjH
iPU4Q2Sf0ipVBSwYKfWPyoVpwNpws/9svDMfrWK+tE4lGZa2OJElwy//dSy5
g21eF7/8Ptq25fa/K0Z7ox6WpYmL8n/ZNx+2chZRLRr0n9322Oof4NRVFMvc
9HoJDz/8t6fFWAiRqHkf/fMmKz3RQoBd+YzYMax7NdQoK4pwtUQYlt7x6rM1
6RqRALwr2RBNnMtzVnGozdFsE4WybiJhTFHMrUvSFNlEkjy4lW2yuPGKQpIg
xAGTVLXncNZXYWEPMFMQehqbWpj/0S6gxvlQTeusBeQZPkbbZYhAkydqckGk
SMfKP/z2A7i8gR5efUapGYZ5DIHfpeuhaKGtBKtxBfST4gYdHYBvEh4Vz3EP
ZbclGEOho5LiJd7EU0zNoTMoFDAdyMNmrojr9MRU/t1TCAWQBTuhxENmPJ9Q
xlGSletNRULwRINqELsAbMe4CDO/VAtvBSRXmpn5XewuxN18bvMjAUl0nDeC
+4ZMCTi1r8MYN4MJxvh7AIRbr7TZjJ9XRrCRK8KGbLAq2NZGfP975gH6cXkj
cwIqBWXenutrMAcuuN7nijyCtdteLRyIRAqRvM5gzYLJrD/RU1ps/gi1LviI
1o0I8l7vX3sSfs0vKOnYuwjQtfhMu0EScpJfQgU5ammZ9RXGiDPI0nKxi+xJ
ZAXBHxwmS9uXNYuoZdGQ/qQEVXosa9DkGnpOoP7HCL9UTwNFnxAtsq3GicCi
LWt0luzisaYpl4J7MTtEj1Qje63uipFWgylO5bABE4ZxAUMEpfZKz+/cgQ1l
2SXQWZGM3CPyzIBiM9a34oPDNESJY9blFBXa2PFM+Ys+GhpJ6nFXMNB6ahJo
wmr/digqxCFF6JcxLdZmPg3GzarYFxYlwR9v2NCW3UmUZWYRwfh/bu78eohQ
OEzpFAGJJp+6ZBbciyDZumtVk4CPYHfMgFmRX8UpMIY+JgtTDlFBV7LpX48/
oOnMylHtdK08pPfYWR8IHFkFPy82dLkTkLGgUrD1hjvk1H7vhP9NNIUtsylS
HRMGbUPxy+Rd3E74Nrbd4Dy+yR2WmuxuOXK1Tw4DRxRtd1v3j43eFz9ALZrl
V1ADjyWVS61g5YizlZEG3jd5aMTZsvNdFXQR4zx1KsiRESGXj6hx82WI+jHC
lyd6CxgSCC8gscPwXI34iBKJRihBUb4BDTbiECt57AT1E9/Dww87pu9KlWL5
WpRDjXBFMud+cMDbOl2Va1EluQRX0L1a3dXiaqCusUKRdV80m9OfTXfn2CJR
gUTqGf4/7og5EqTFVlGy8ATB4eTStvo11cfGXJhZJ231CGXUEZGpjA6dPpo7
/QN5crhAF4tnXe5Y/5WgIjyWZl7zquulMCQHlGs5WN5Nj2tIc3rVsgxUc5vf
ERjS+k4offYihoC/5c8Epo6sTyhK8qvY5GbaODMA2YmVXNzr3G5k9uUepa+x
ruZkQfO98uumvnSYdQMUxJFLA7jfeS5wvQMRXWtpQLPmh7KpMu1SRb4YJ2g/
syeZsKjLx5Nxuy96vuw579PPxJOl9trZAE48FspwdQZOIIhIS3D5zkwMGnOH
hr9LCdZ3V6HcL//3Ioyze3d35mZ1SUJUvAhNAZeimpaXkYER28jPaFFh6MEi
bkYdfKS95+WmCeLRdBNiYOlMCZP+znoaquNcGWnamiVe73NnthCj4jarE28C
ST/s/ciL/QYR5kFEa8sCyj+rizA56rk21sSBuWs+sFkgl9NpNJgv1NV+m8DP
CyYl2ny3RB6VcfOevACwnkPqVhraRID9HIW0zZjV0A4EJYWliUFVkbRJKjNr
1sTg9dj2vtC19Ks4uPDSwuMaPRHmilPBi8WVk40BO9e7qWgZ+hjdH4pnF7JF
ss4zXSd4pUeQLndOBBo+8JjV2IfJFdiG8nBfMC9D8OAa48TJCV171Y34YntL
kir+NWx3c2rGkzmrBQjxkFfR95k3niluyUx5fzOGKSuhxaIrQ4dEaoOrdIYx
XU/FogqynZvdm8IkMUiPf4PKEZP8Rh7PIjtHpLObyBSskVEXskJlKW58U7rs
2PoHcsYnO+RMNk8J2guuzk6JgKjzpJ3eHAir5gmv193S7wFOdiyUlOtrKvlP
KQpX4BDkYnaRaXbrekK9OYKvJVbWXSe9SbSST7w5zyo+79zvbxELXMVXyADF
XRWRNWNneIi2uYYTHrU+PeyBv0UOJ74SC2TX/b5KozfLSNPmB5mX3HA3zM2E
nFHuHa76d1umIpWZwN8/2JPRsZkY3VG6h2puUW5dADOvOPwc2DLi0umpYO2X
AcniKPDFLICsInheoQATVpyxgjm9FpRoEQvJDBSjhYy50/l5h4QhyBDCDZxo
VmyMiOgpWIxg2c+VZux2X9T2XW1UmmKeMpKfkQWFoZw/rE+Hd82iTXoOpzmE
MGxYOd6m7zv/tGC+vqyle+D/ksezcDOJvlhDWM3R3q6zHcdEotfMWyyOdKeU
789u6ircq58sKD0p+Iyw1WmKZHAAYP+Le4+0+aSJMCxsmB5vYvk1pIV6uM4e
XJ+oVgq7ycmXULXvGm2Oo95ydWfsZk58j300qw7+hKnx0VbFroErqUsrlImR
9QBmWhypMcDZs5AmlTVO+DKkSEOm41d3d0USr4qo1EkY1GAkRRSwq38JlVHX
rypNso7hiV80rUEj9OrguKOuIlFo4QHXXI0DSo/HL3Z8XOVBlA0QEPOw6QhD
rup55FjlcaUWIX9tX9llsOuoWVG2xQOA+v1gpS2CioTTnalKnJnurVo9VDyr
n96BJxeGQAQ/cQcEdSJDsVnEQh1Gp1WD6mmDc0/n5043c/yUq6ApcKQppmY0
puCLh+6i2npVMN/f8Q8uxrWVtkc2t35luZZhJGN/xhZwAjiCQR74kVE/mb8S
YtwUKfT1K71zmCcMqSuwAvW7zzHTTjvW1xqdQpd3GjFFArpBnd8SOpTKl5Jh
jhb2n8aYvmDhs90WoItapZXvcWn7GluMvx8ZMEHDMfG0ZRfgzjbXOb/2RySL
SWZ+AXK+qrc6G2kMsjDcw1ftWaFRhVw+7hcbM33aRyTYmoz2tMSJ6b69JPJA
H7Zt6iQyu3eM25+KvHOlaKAxZGX51IphZ7kxS9qxqimrktgLg75Ox3Ey4tJO
pODj/zyMmIX9id3PRtVDSZvX6jy32bHuVO1lrRMipGqGnj8szjTqddJjNYHE
o2tzhC5aBHWj3eJ94CfTzanKW/UY43iuwjquH7gZ9S+upVtxBnVfXdLV0Iqq
ugBbJf7Gwmb1hetSJnEZy/YpHbYhinkN3IcTwsmitNPHWXqozPmVlxVyz9DU
JoKeZOryFj0APEbYRzMHzxvtWjs3RvKaoVqQGRHVRuUYosfUZgJAGVFnPmKB
c39bFIGDjw+xADXWPpKWLL42hDsffS13ErCbRrZU4Z7LvB+dK+gxWAYWrp/K
GyChazonrU0xL3V4jUdHB+ChMQ6GmDQOUgmdDo7EZATaVYAtGnueW/sUrQYL
QmSh5F4mL0lTCU9O0J4Iffoc+CjiWV16iRdumtAAe8tj6eVmE5WY2+bqYwOb
V2wsaB1Vw3DY71lsRW9mxCLGbGXyNJcgQvP2iAoGy6mYYaB5IoZSEArBGaPU
FBDGTWFYpFNiriTs5xLq+owvcl6hXk+oGisY3ytf0beA4XdwGyalzdWtCM8r
ExzSXnQMfD+C/RIDxdsTXAeNn4aGmz1VZ/aD1qwSwb9atwpfx4obg5l7FH3m
GKNSEQKS0QlC7Ady74PYqELyPyTkQl7n0+9m+lfu70lWcyyoFN1q79rIYRfn
h/EMA9XUC3Lp9UzkJ6bo/8SX4bUm1AUwKwusNTcTqrsN1T9aeB9t+buVOs3P
0FZT6St2cuw/J4bVt2EBjUIam0Da3P+pauuHHta9YmboPFtmp1G4fiZa55jO
2DVPJ0T2bD3fOVypl6eoO8GS5FSCDGWi+3wC/ffxiyuXSJLSaAHzfJujZmi5
zbqHCBPGoLaxZIC31euNZReybUeDsjtvDImfyxTKshfquOILVzRjBqkAl2JO
cVB5gs5UL9RJDyLhXiFrUg8WjlNAy675tiiSJBwFNvs1s9pfsKi1T1UcizMQ
sOFhmshNsOI6xIRJF0L8RpIr8zlYx9bHRhkLtrPQQw8laxFHpudDb7J68YMc
MrZANYJjpZX+rbx0bDNR1bTEC34+6kZmEVU8de3at46hIzMXt/UjO48uSF/j
Z4AGQRBCqIXBCBz/Bb7u42BcjUmT+i2V6Mn7x+ABO2iSRSUiC+bjszI0MoAl
JW8XSxG4iKXG/dPQZeiuW8pNpjUtkNxVJfqGWDgVurFfsgD3x6GhE2CTlcLR
mhhC5blOywxfnqHhnK6w3Er4QEZpVDhcu6fJl3MRigu3173khuUUGigdnQMa
WFP6QXAb5+sMX73Rf6UE+cXtsjlVXEdsWrZKsfJ0AolV4DjHwqsbxm8wHEZD
/7V2LYHiOQHx4KA7hdawtN4Kft8aQ9nmxAl4wHiY8DBL7TNMq5Jn+0IcJEPr
8Owf1o8MHV4Ln2FUy+kZ7EQdH5AgmwLwvkd5FnVe1pGJESv2ltesdWu4qNm1
2kv5GqYPmXEU1prPeZL/IJpJLc17SJZ6ROqyJ63qLjdoWCLwy0G+cG0RLrE8
I4iRtKzXMIrv+QjgoNTnVwud7kO3H+JXVjpWNhxRTu1ID8dC7OF19qzIVIhe
vmZUTTsDuH2DlpPiI1GH4ciJJbyON3tyZLdXHjgJrVtCQepGlhPCIWz6/P+1
zoI47cIyxp5load2UtdrTi264xAJXJis3KiCQ1U0v7VeAv4Dz8OJ2+z/c9UC
n9JD5uY4uBUw7inuu0YegLjTcrFqm5PWIRb0KcSvGWizpO2g4uUMgSzzFLvc
wx8rjycvqj13od7Lo4zFLwCxpp1JrTf2+HeXJj12dFajhKJInR4MFATWaez+
nkEZMlH2q9p7rZPsmZaKR6J7fM/XbbQC3TKyXIKuJMUr7DjGmXCwC6sSbeE6
SWFjPb9zQl9gmC8eP4RXev6LxGnEGA91IrZxtqz+Cu7r5PhtV3BYCk1qpFS9
yoWhjfjPyPzIIoDJWet3nI6VXFgPmJu9vAcmXxWx1yvjU3g7j9MjdCkasI41
Dx/M28XITQcJC73vFpteM97duA6Sn3/8c7vfzOktdb2mHaQkmkPz55FqPbtj
1vm6OvPWeXiZTzKwIZxJX3frISSO1H3rvuyXc/V9qCAx0buJXyNWWdhys2jy
OPLH/tzMOdZmytHHDsfJ56O/PPlU0/UvAB5VNeZInBp51fh9vf9aN1MV3/H3
wNWjWBAt/5Qs27UcC5U9YHE0EX+anIeWAk3ALUSh5y8doHOrcSosL4h8CsG9
lFbeW7pD26W/BSk2oYb3tOcz20TN3ZefQSbX8G6XwQK/Ui5hP7vrxU2wVpYs
/qPDgwwJkeOg+y4c0LnxyU9pSM1vf2uSGpd3BgKFiaDKRGA9qslcfUcM1809
BWs4LraiYMNaeXbsdEt4WI8Hc3aCTP3GWCpagf6YyDyAIvjjI1mqEkXjQzFn
2itDibctMBeluJRVBcv8yRpqTpauHkQDcZnwS7Z1RPztB1tnoVbs1RlMHajG
pLtvC232/96mfVES5TxkVpBEtmMGx7kxhYWCZRnkiNUALIW78/Fsi821kkVp
mZAoZ9GLkhvqRUeTgW1SxQoz/4klewWtwnSBjOCkPNMWgUeFhqK5B10G9a8k
Gu1lxnjNIAMiDbocXi/OhN0PcWzYKoVUsJ62rHdUz8kFBmWysqNg2r83O2z5
uy9ASxnd9ij7bVUaZTWULittvnV0347xmH+rxIWY2QsbQviaoOs24BMdPIiO
tvdWNCXFTy0FlYlgN2CvzklLDC6AvflsB2KNLPVxG1bTNFwSLYYyS9wr76gV
MCeqeTfeuTcMiH8CNbuXNTvs4pWMOMjdby9T8+sJLvf+boCIyHwCDZg2Kyyz
02lTgnHto+lZHxVSYH3Ux0ecmpMT0lBQAfbHkjnIPJFqTaetxYJhP+gqDNYX
DElHV+PpNmlV+3QHKLbD+NkbnjHpRQD8Wib3p7igjJXh8UnX9uLD8TjIuzbn
ljCoji72qPWog1+TWlwDwuA/fHTq658k5nACCxNOjib6PvNMBICpCdPF4w5n
P83ClkQc4NZjimuskcRA8FC4Z8uE5dyqK3j2pH/q870uS8Qcv5GHFo19iC75
8WARHUCKIT2KwCVfRecEuTNYXExo99LjphNDYhirrlFIgGt6WsKpZyjAr/CY
4fEtPMlpXQswFj99V+5CpGcyow8HCcFVpztZL/tQtPUsAZksOoINasV+CnER
UE/b9YqhU780sXfgjQafd89vYn7Kr+J6BO0vIFJq/9qF7VLYYZQhGpDlSek5
PtCtv+UQPMJfYENVu1KCxZzKEpTOA8bKnkEg5WkSV/QXOOHFEmFUaYMo+jeI
3FkhBV7/LYtO8YOAiJ2JnvpyEFYiUWAE4MShFY0QccKl71VzUWnonmI7Z1C/
YLA41jBivPPu5Dqn7rNVuR0OemB55r5SgEB9cnl4/Lr8CR/Zw5kRw2HCUj8N
QgrWePp6WYvPL2rmYyUX3T0rXZ9RD/FWClYHhHSd1en/yvJH8j/+zZrFpG7x
RBF61nvJpG9QjsoEhbld2F03qm8cMDtjtSBkM8wAfneJ4zcIh4N4YVipBe+R
2yEaKoqnmw8nUpPSKBdg7LXZxtv7R1135qi2X8xMDUyBB4N67HsYZNPJ3ju0
HuvSWiPz7ayZsO7i9/aAjEeiaeug1mvVFP+ScnWog6+ziA/cCND4MYuar3U/
fvgZ2I3/i3LtDkcQvbPdJ98W4GOuA2sKAeaz9MDVaq3Eh0T3Yr6VhlRreRHe
dlVw2bqCPTCeziNG2GGPBzcq/M9L1/SD7mnCQ6k5JHtOap49y2QlAeen5o5V
zRg/isRZqsOYP0i4eVNh1JF6RsoLTL9MtrFFTkMiUiMFskEpBkhbJyisdRGa
hYXU7LOMtwNvRvguXsU300BKWQZmlRulWGwu/oQs5SkRT0tQIIIQuWNinA+I
pBG5/fwM6RQA7OO0PnnjYbcAKPc7Ab+miK4btFvtJ15vEczzQ755eNbLqfZ/
Ldezh8FJYr6yLUVpCYMi+XizF0nWqKkruZSblHckMeIugXGGGT8nV6eLARtZ
d1lq6XzRupy0KOHwMUCC6yKUhCJ9eFNLJMM9eVsIjvTdIjPdL0pYBMJOcMMI
JwDbOp0b6Ns8U2mF8reKoTttzJ3nfgsZQqnlXEzINQhLO35lJCvBxByTPQJV
iQE6XQ6xwX0MZGZNoRm/XfHdUZhI6gR/16G/c4R8PYEazGsW0pZXzzoIpddC
dXCG/dEm3/G18dyQK20ngYdnqOC17i6WkmKYgJ/UqZibGpX2r/hxwwydfR/A
zY3SVNsn0JVlDkFR73Wn7X7F2nvMdwHOKARWvS1/YN/LvVGPo3f/VhzDhAM9
aB0iK7eJQ14zagalBaCaoVRpZ/rApMQWfIS2LkeBwfjMvK88VCwkurEX/MDW
DpA2NXr3LAOiDGwSOswCOh1PdGZRtHlgCRb57caCW+2hpXj1mcZgN+U7yr/L
UzwWJHIK5X4UYUYJoojfEia0J2VLxkcc6S6jNj55Ib+eTmTyTUuUfQCzA5DZ
aeXkG7sKeLO/TZoueJGi+5C+XpF7T/D2jn7htBW4Y/4TqBXrwS0/wJYLi3LJ
uY7vcKOYs2H3/b1w6ft4L8Me7RheMuF5vMCfjLfG7JUJKsZtwPkkw4Aj4dQo
kw8txGemrKtvZRL6GBJPr7pI2FukOY82tJRcDBHbVDPpuLzvwSnjqKMmt2It
q+BCHMLjROhlOolKvMB6iDAxCueX4CRLwhGV01X1SfYQWkvUv2ApDm6uANsq
HLcK7k+GoAd3lALyShnk6JVAf7++Q63HF+6uai7XANwPRhKjA7osHSu8xKaF
XwVsu0X3PcIihPDg6Vm3H0JMRhSJ/ZIYCjWZLzxnS6R3sXOJD1JnoDv6uMf3
1OtCF/pTV2ikD1mEn3AThhZNVlEZEjsuvXeZe85aPMF1BcDTpJ0M2fQKbj5A
4hhfIXHr/rYEm5ifF1f5LyU6P6UrY7zrueOKHHj+TtLP+3Aga+4m8qBzJM5Q
tigDQ40VBswYNya0VcMq64Zddpm+iPQQZtrK1FrXe47sOYCOzfz7/X5CQSFS
SEya869sCd+Iis/G4gbki3Ye3IaS42nwfq1JXiu3VZbgPgo8mehDDuuvn65E
x7STl+xXN61EIe2BdATIbABmM30QyTcib2EvZP3n1tKoVdR4fUg1FuDFC8Pr
9krE6xCGuU3wIQ9uLzO/4nZ6sMzgOa4bICHrBOfFZye+yRTIMg7tl9us2v7X
8ltP9+wwTXvaVbQRciBimtKM9ztIVe2q8qwH8ar+iqftwW7DczB2C+PJ1CT3
m1NUDrGwBH2cssmbSkZOngadHqbWoeq+niSXuM3F0TfT6AWWdH3fEKR4DJUC
KXvatZaKbslfNnCYFYzxbLjnoJxwYGdGEaXgYhhR+KuyV0Zt5klwd1VbH5Yk
juDyHNRiKutVmNzXXDvO7op77kdsnZdnlAtX35JOv4jhKVwZa9trmgvHYjoy
Hc/btXj1bO0VE1K+ZJniOVMUk7VVGxMT+XpwBJRLjm1/oSh5VPtcSwaswnDS
LoaFJzveaB2Wl/BOxFKg3Y7MQbEJ/g6TeEsXTBdddx+TvGqDss9LFlODKpK1
wgNeo0HGI4iG1usxFHmKEq86MSHKZCsgdzZLRYLJHIGIHCiDXfJdNm6hg9rD
FOQKQ+Z85NqRG6XlwPDtqrD0NdAhcf7mxc+dC+Vi5ROGlXRXnnN8d/9dLUl1
3LwPwxRtwiFOVYo8zHmKlpK6HxksZ/K1pUU7c/Qon3rtbfKhMGyTvdNPVgbT
5tBOSJz4vzcoZdV8uyxcQO42AjOUd2UoZMaLo5KgGlbeyrc0OvVGT2zi5bFT
7TcViP9ii8CL7iPTRaT4arD8ty++Yb70s7uRAf/aWWviCA0dE+cNuzkbQC8P
WJegmQxMGPXOypWh/ThTBpMuGnz9ip/rVzhXK0g2aC6mBtrwjhUfPEs2Mncc
npubmlR3s+32hSEgZHn496xOmd6GWjovj9w0lBu2kOEdqZsKZM9edqZEVX90
HVnLLinKTymFkLHrTHJhOy+y12yDj4Mb4O7BhQ8Kp8xojjgVOmrXpRYZ3W/P
YI2Yb2Wu3Y037hjRVqhW7xLKkh0Hk7rXTndsrMrZDxn4oZ6wl5mFpRb6BNYx
FUSKELeCPPHXfrmnaCQg1rwGZ5kcqmq9cb7KUsObBuAPzat6fXx9jdsmMs6k
GDn234jtGlljCcWACBfzcTzL0EsMIMB0i1ODaAJPP/STaOSr5ee6luzSWwQh
JpZatRv8FQhvLs2xqVR51jfvr5Wga/u17H8GgG4O7vnFobUB9KDR9XJbT1Jy
sQDINn5AixgQnE1oSNR5TLH0ULZFShsYJzugsKPpwE2ZPAJSeu54iS6HPqGr
uz62DamCojVQcp6b188mFzafeUNXmT7hJOrYZMSDSHoT40FoBmRpXmRaPgci
PwyqxfbRy3vILn7yRvo1ZYTo3OiKN8lzM2U/qo0R675DgtHhO6Gwwnjz9MeJ
5DIA7V07sDAIG1IRPaRP7UyqaucM0x4vfmqBzHpfhvW4uum7xxNgur8rYF+c
0CflDVXCbuFP+PQ2OGClC0mDcEpQfPx3sgFJGN2/3zpeArgbQwRx2Jw9ZqWT
bVG9fBtJqTpojMyE7fFkLbYklXS2N789kbAey+0uBpIKnCeyOQDODgvh2zkz
uT0pa29d3S+1ya+9t9JQb6MUKng55nFDhx04CorjfBC+CjoKiZ9f4JnqFpLd
cygatfAMWk9ZHSoX2nfn451sj2lVfc4qSKJeUeE1fxugm6/JPHcDOwD1NRwU
cPnt+AItN85W9alQ2KInW/V5K8LxyyaCeq0LI3bFrUbcKk2Hfg9p2aBBxQtq
44GThAX1dCz2bL75x9N5g2THkvPylphfAq2WKeDhRDoDNtAt6JWTSVLusEfj
HYPQUzjiir4PSXbZB424yxwmQmrefVILNJ5KQqkDPZy29BbATGx/qZs3Ir/d
9Ri2d6mJAWylbuoLXq2swvo44NB0/bkHWktlRW2GThBjkcjCP9C1jjG1X0VD
ahGhVr3sgmajaEBG3h9OZkiETYaRRygUBGN2KfwzJYu5EspVzBDAT1+5XCm5
VnHtPhYpiDJdx5+5XPKe1thz/QwOgnYJ3W08Ib8zE59g4FAm785PPw1r3VWK
GXl3ymBc8bIpe1WrRJliXDAwcbw6C4atrq6wRr+AHYOnpOd6RtE8Rfd3dARZ
eVOwEtgUkGw+fxvPh1yVawdJC9jN5Q6n+4LIFuefQaPD+2aYZbtOuxbAoNCO
VsyYYsly8XIhejV67MQDDiR25BlvWOOaEEPvfiWj+EIwyVYR4zlgaEM2ksCj
btXk/9J/m5yJxWOkkVMQN7kukPj0vR9Fw/Q3vMMflBR43EevZFXTXIM1ZFPk
K60wTGvDTxK+ut1/zi/0WNk7Q8XWs4BQXiQp1F1Mr/J4wZS5Eg9rVtr8mTmK
rK0vxcu5sWeDK/iHCQtm9CmTGLDAtr/lUL427YFwpWzCyG6Gsf67cw7l2yCy
4aX/L+fA0fO/iIefKnQjQsa7ParnvgoUNXOgDCYQdhed8MBdeeu8WRyFf2ca
EaRprkz6Xi0EJ//1tsk8XdddR1YsPWZkFjyKPs5xLYqeDE4HZT3dNZZZj4Uk
Bl0H/81ZF8Anb1rm+aeqcnopOGnHAdi8khuXboBjw/p+pOhYowkflPGsFG1T
tdu4yQbsxQdzHuzjYG9tW6OaZnm/AlekgxMZn04W0d85l1nHCoVkf7RS7grA
OisjggJmQV8m/PI4AwR0GrIFUP9+4nUJtY93S8APOGBe6/xCJ+ZVmySVTn1V
k2pfkJEIk1n2H3baXg+uDqNgQK7KMw4UkbpHBPuwD/WwaigTfFuIjXS5Zzlh
MideSYjA8F+fMy5xBjb23w22PDJ+vbBAwMP6G3CTtcEY5xmd/6xWITS3WNqi
4h4aXMaE5xBxJ250pSLpY61q1syT1INK4w2O4iWP5oharzTl3pFeiWymxtTE
lPay1GwJ9+Sxkw8m3r6UU3cYAYncCoH0NTULnl+Fy3LYUosbnU7UAJyc8yW6
t2cfiLokPYitDyQfWxPQwZ0clTb4y3BoYp22OEwKgw9xizGcwbOYt+SM98wi
ib18WeyJ/REU9yxD7uDyfZxwP5hJ2WbxQGmU4duUlT/G43sPfC3SPHetokq9
cocuNKdXzPUQD8Cq+F2TA6y+w69ZiO/49WqMKj46MwHUzopglCZsa41LsWEO
Bd+whieEmeye5vf1wpZz0dDVuPDNhzcDPXVAyL7dqeeGcwIG7yGl1AhhqHnC
VK38VCTBPgIn+f9Lip5BENpI/FYYp3GsmxX0XVxT2LM93KoXF+nBxs+JpQ2x
1un9h4fZEkHPtBbPhCsUuf0wynXgJtyIhDBYPNn/JKUxqdAQ3SGrgIrfZDLN
aD3QNBgX4bOwstmR06PNGCFq+17kr76g/fvTB134dNqqF7rkwoAxyOoVa3tV
9Kvwh5L67lz7wJwYKQiTsEx/MMwrVnUhIYRxCZzHBmH/DN6XHJPKlz7hvlcn
qRxq1a5u4I5VRbk44D/lf3ifBhph1xm19QWoMdlNKm/1d6fTcUP2noZpHbYb
MJnLLKSYkPvWAqqyTIKy3EMyRj7LpSnFCcblMBEBvMm5kJedvZjqZxv6OKBW
WYNSSREQQefVJIRXxqLtZd/rUANiy5zLePsE2lR4pl9WS0qGemV4vmEQHfRl
MaezPhQTftesuvrMWIxKOpP3CVUL3w7hfCRumsLlVQJpal/BGn1hK1mgCMoc
0anc5kR6wGXtd22fvGY8mTWnvSh9SKgaZx0M700f9HJAG40ycBxeRLEeohv/
fUQjcwlYo7yV1nAFpwJfnhBT5avo9aAXrzovAPGVTDtP72M5QroRPNF/4dNN
cZyu379CiFpR+tvKokioHZIG9uqJcpa+Ore2Apt1zVPjEHuf0Zja9kXiGf+c
uv0D7qEIncP0SIdpdeW6YHHVul03+DcRjatW861moFMj9nDgvQsMOte0y0Dh
+6UudeX5YAOjSZe5lzE9P/EXjtmZ1oLmsgJ5tV+1Asw2Eeg8gDRMzALzEpkm
U/SL/gs/ekyTdYtOn71Su4hD+yr9DOc9T847cbydZa+Skuv+MqToW9YH35QT
w6GajqN3A3y7gHkbPwX2zXogoGonNKkyAllAPrjnxJIv95BNIG0likNuYDU+
4dtux1awaofIUFglW5yZ2V8T8du2ZEzMre2uc+iT0sjjI3KNd7T1g4WZGZYX
YnxyxN7w//0IxIQHqC+bC74xdVKyBYY7WMM6bc31i5M3Q9eFk0PNW4OS7015
QGkeNOBWs5RaOeXWn+zzOOBo3waV/gYb1PcSsNBdRK08ybf/Ngq8oGY7s51S
lIVpEnvI4ZqAoqCyimEY9BBLLTeSq6b/zvI1dq4JAS8Ep59ORzkpfgXSnIR2
S7QFTKwAq81UG1JbqrMy66dIiV6Ghx6JttAcwEQWO/gUe4ETpLM4AGvxbFDw
/e97bj2IHSH+ncvtRlT1qdj2qFdJU8SfmnUxd5nl9JxNwBC2Mw+XXJIMPeWr
TxRWH3CjLxlLFOVBj/uWLITGXLxrB6RhXn8seMmZriMP/oHiuqykyqKVvwWJ
5gONg9XU4kEpysqzU4afyXEVjx9OXQAyn5uVS8k9/8BaDuSRMR/YmAWTndDf
J7/B3ZiA0znU2PMkdpd8ftwep+juXnelyI5sn3Gr+6PLC0PhVPTIFvq5Xkze
GybVk1Nic9SB5WMRYQq+1Zp4Synt61gFQtj3YTjlEoSU4oGXZTk2B+HGQnzk
sjiM89uVpS3DxA+BFO6P5sSflDsbmaCkiYkMSXFU3CGv/k6pBeTeLSH0C8Iw
NgRtMj0dy4RT7kHdL2AmY5cGTzYXHXolLMeiz4eyPYCveT9nQzRwjRnI80vH
afs6G3a34xAK1GMr+uY8tzV4kk4wwywoLe+ZnMQbO1TDznnaVvcR7wdJtHOV
iDYnBI6XoqIMQlSvTZZxTTs+o0Uxvn8a4XQ88Bzb/B6XQhRGEOAf35XLwajs
AhACcAE3blBPuBc/4LZFzDqyAAMm3W8xG7y60yzSusJC9nZSsO1LuzqEtuV3
tn+hD5U5qGz+04yVvn2P5PKJ1d74XlEnDMmaBx5amHvm0HHfRcwNA7rX1yNy
2uh8Rt8Bob76gGV4QaHhaZoau+CKLvHxV0MOs/ToLgEZgfV8KiTiQIA5EMf8
sa1Y3fpShyD56IDYGHrFu6NAb+y53/5L5RzSBJdOTf4WSU9p7OPZj96HsJCp
gVdF8rxZvNIPvh+PLzwDXCR9xfcg3egMSSolxatMTztWDHGGP4HPqKMMyOM2
WyHDRkFlwRdWdUghN4TFVwDrN/5YFwmlCAkBWQA5SX5eAAuouRpyHajM48Az
dQ2MAZE/DZn0ua/+k5vmH5xG0ZwHteFDlSsMFcwq4ezfWupUvE2c/bWT+vwC
AjVk/dg3qp/m+xfhXclOkb0Rm7TH8zsm/gF6diit9lpnmQ46ZdQeYlHQW5p3
+RnQVOJDGl23nIwaJHAGNfy3PXjnT/XHSzCXwuhMZ6LPw6Wjq3B+GPefXcwo
VndMy8VNeS4LTuVhMV5zwEH2AGrvd5jtXV5TCcdNAJQE8f+OMNNJfQ4M25+M
LxtEh0raWkT/4AtCL79T69bGm1bVtS4J1bgz2Y+eBWMOzm3ATL2s+8tlKnJG
kcppXFiftzsVr3UnAALhtLiPpq08U9x2HuX+QKh9UszOAZybeQVqcSggApA3
NoOehs0PaNXc4ffygYxY8a+IwXq2BP+ALIfL1hJpI8zDnPPKxwGP+4oleaT2
Jzkwf3pJHaONinpC28xifIFrp9ESpSkMDSElaSQKaG66WqPR65qNC/pQ26wv
GNjH/+nu1HG6FeKenIDqvry8TDBYD/2n8FUZJ8vw7As+3ttzCM52bbrRpG9P
wnlsiL4J+SjiaKKwL4duz9Tia/xCsoyspHCe2TxqQ8Adq8qCi4rXaDdrDKep
6AbyR9yTx1LaZlyEk6P/p6xUdiP/DkDnujSInCg9milbXta6lqh/+zLmUoWP
OZzMYX+rqJ7Ymn3ngZZTNyjf90UHR3gu+qScFmT/d7r/QDQAapC7Lcpwp/KJ
X86WZe2WkdaYKPJPxJ4+BI4tUFfJnntQ6bF0ynl0KQLXgi2SH5xADUW7aSrB
CET8tAzR+sM8MfP9dXuRz2Fb9qmrXk26rLEw248tcuEwSluoVMyUZkR7/HO/
UT2DXx3/UNNQtjvuUz7y9dc9HeNE76GSYZ6acbLnVrfqbxFUomW9xsDMItnw
/ufe3u/qcJlQmQ7Ln/YfALKTkbPZmIDhKCcu+WBQBJ1gnMrvU9ORrP1+bTCQ
zre9f44BujFAv7Umcty4l3DHGIsSpilI6ubjayrCntI6JeHQlYNoqHyS59A8
xEqvvrWCUrCc+rUHDGejPj/+JPhSSKw1jze1atDCZnlHE99wu305CYHYMQea
MFaTTqpMNQzJpcgSmiDyDs5uqo+eWZmSWu/H4oLWFbiB9Cxzf8wzrGHSm5hU
y6CMiYa+N/PgtsDxGfsU4tZ6ywIarcss+rlGNvphA/rb/6/Lvv+LaKq4xi74
cVqnJZsgXrldshta3dl9Mkon1wZZ1oFJthjTBMZ4B2pwOcyd17vS0z7/vPtS
tdP0tJmmDmkSLji3sbVOZspCVJRES3AafjjiHM+gzxHM2D2MJMfZrmdJ7urr
UJENkElsxKSTanofmzSExOhFyRsBFq2IJy0aJaDFtYT/qaGJgVht3zgXx7pN
JqPwFS5ZETSg8hLngPr9it6Cu6SAThZxRl9zHrBHwq5MBfZ5owR20Gchsg9W
zbl8iasC6YzrNp86d0meM8G0hJaqU2e2YtQ1J4Vlr16BRrzl5RiHuVed7RSC
98z+Cz2H1PvfbMKyULSnTsOpepWWnHHS9Yk2PJGynEEHqV0+ifd2QFVPsXYC
iaAErzWQveEt37DoOkb8c4RV6naCXj4hXrpNzPUT9uqVCM7tjJqww2B1RJJY
EHzjkcj4ktcPVVdj85PubgUzx2fodhguQR5g9wnUGFtvud3t/JwKta9g5Kru
F6yZ6IoKTqvvsqB3w/grEh0a4iCU/0jcSmv3EDNyWfNVEaLL/7qrzQ3qdP1A
5QOyRxMTiHN0uA0A0nFBuW0Z4DEBR/AURRUQE6bJ9UzDe4i1vSCAQGTT0oaA
epCUj90v0BCBbO0uw2VZUF0s14t/2oGV7MWBWVwM6HYV48DnF8g0+QOtd2Wg
iUdhUHTBLdM9Hn9QSiPWAX99O5JZJ9RLqaJTHAWywL3+i73SQFLMiIwb+reM
dm4aQ0O7ISSfqfcbdFM85kNXyEHaW5NVXiJNDkSKzZsJ+5yyVahLmXCROZSo
7bRu5Bhg2TF5km4G63TqEkOdL6OSJQFqIYJ2IyvnvNYppuwghzzt4qBrk9tC
xtF32bckm13xDSpXMA9KmWZ4vCVYg3tYdsC9XwLeOm1u7IVmhCjpjcYlH290
+xp/aGUwBF8o/UwtOlhCCd8NIvHmMvg62SnMWso9O4yjs3XzX0ZMTw98rg7p
jVD9bbtIKb+iL8zu6E0Z/CpdPovW9ss1KiOHB3faIyJqRBQewhsAk5hi68bY
3pJsc40V0D3Ki+8vZ06cVQZ6BnM/f9c9NbGinoVbIhazmv0po3XEJX+/z5Ln
gFzKjKmLtxCR9oNblXz0kN3ALBPnd9YW6+irXlx79VhficVxjsV1uNxPB74K
pp9QHwo5iyUclsgKAIv2k3D3wZJU+YSac/B6LVwOVgZp7UVHADalzxyvtSdn
llT6qKjSKr6oWsy3ksdRml/tuONqTL+ZIZOmQnVBAV9JeyKJmHG89jqS0rFp
2nZ1rdjwPIU9fpTUfOoOppBXHABWqdSO7rE0MpLSQgTet0yZzwx/37Dl+IYW
zU29DXDz7f1H0BVykQZxLsd7rSdeNVKSpzoVQEUi1d6/CozKeWYFUwg47gHq
21KLlxXvmROFVe8RLaUiOW2tZRF4uzS6oOscx/uaYqmPW1UeToDd9psbVs0d
RXEsRuqd2rHudpY8XHMeE2xOCXFJYjBzAP/lZaxGz8jlHaqOlnhTLrZsHkIr
r0PZ7vkJMm7xaSGNt9NaAwAXz1YiBDam1P+hK8yyK5mDiyEKnDQUZS65jqCY
QBw4W1LWgsVcInvjNbO4H+h7t5H4IOaVjNh3o28rJyUk317UoT3dVbsbyum5
VuVt4UT3hU6v3cEAsS456DuEfSYjY1yfTlXfCX2KqzMnNXU1lntbt5tZvgw9
rFQrG/VUsVKAO/zCMmIKyRSCOwhaKcvUsw8nfYnpGEaSJb7yDMg5iwg1jG4R
C3Ia9JDpS7haxcZRWBqgBIGq+WqNvg6gEVO+KBEqFahu+jEtXvhppO+t/zAS
XRwoIMzk/E5biqdczVe8V6sSFtt6XCDDAeml5UrlEErBR9WVjzIV+A6SkRll
SWitfjsO+ij67USD6LDU5e3lPeKvw6kvi6mBHWZMXa0M0V3g3/pScZKiM256
oEsX2K/UN/VBlR8ByO3KqCZaxpceiM/X/9eDI75AtpcXSD+lEKiik0RUptlY
paX9s0vh8ezJW4n3/nciHnUU98YtJXCLfdaMn1cwY0ioq6jejpDU5aWhmvY8
ryAEN/On8pLuaXYq3A2iy5+NBM7bbslYs2cbBcpMxqkeemZ/XFYJPFrR6by2
5w5gW8WmCt1sNhsXlxfkN4z50OpA2LPt4HQTO+ktH/4JaUUwQ3XUP4L5WPeb
r7bKIbKW7Y34KQIvgokO6hBKpkCUHJWgN1JsxkGx42UVclv6mgR1KRvw6QkX
8DqUBpdyIO0NTZxe4pc4umFhWQZ7jGIuLDYaR0n1q80XFDt6OtpDB2Y6sici
OdSahrHiAFwWl9+DS5QINTXVZMwaLfcyBJZCoIE/kJr0H4ycSrPQ+tAkFhQh
8ylMlhdYvO8qCNFsHlI5RQ/jn0GPDFDcgSb1Gq3GtPb2S+TdcQxvqtKXMVjt
DT1d2F4o1KGiPcJ3xIYDX0Ys610DyFkUNbZdocKBDM+YjjcwRjHKHxMI1o/q
KLho8ud5tMYi36KuAXkgMdf0XlQVHP+O9RVU9DZn1bFAKVUpGkhVTm+kNALK
F2Ues3c9yDeLVK46vJMYaBdliDKV0Q3lwr9YpO0Qs4s0FQG1HlEUzigy6cNM
ck07ScUYDyZ/b0gXVMG2s3F1rSMog0T/CPR5phKOs9+oSj0MaSrrkD+QYIyS
dvDd3A4pP42dw/aBUaBcQDgQnhEyFvM5oGcvgjDYfTF8xHZutDHqCfUUlL8S
frPydEVFM6jfQdhNYmoaxE2CRXufeHMCK7HmkupqJLAqzkxDGHWRfy0mjKjU
Y6SmZAmRjHnBR0UCkSbzuiBU8Vw2jFjKwTdVKr2vYBtgwJtapvit6AIavu41
4vsaCBWG5479sF5Dr+gAqHoAYHeorQiciZPPOPgJ6sP/2cbZTQNFT2JePV7u
cwJhcan8QZ2KKOohkQ5hi8ORaXoSKew4StktYXEsTYaQL7BdejOQl/kEt6z5
GDsMRMHj6nrg4psZalfxFKArNbYqA0bKb/R+OYNhMIwmYd00lpqk0Xz11BLH
LZYOhLHz6hl8SOLTZa09XOURcTce1maPbkTcpLNvuoVP3Wsjj3TpCw+TxjjV
NKO+I8W64LUgo3njLOqGu82SlHBcjAwsj1XK/m4zuIEPbmLQOBlqbyqkCS2W
KdhzYgAuMG3lOELcPE2gT1M1juofKKcVpPxN9w717g8+TkXBauGovW176by6
CUFP9i48kMvFxYkSu7umLZYDBvUYXQwcjR6yBk3X4IAd/LbmX4KVZOh5h9t+
Yalt+fi+kLYk56upyU8IxYUq9sxxluwFoHweXdtyqhRLxxa2if1hZWqdmVte
VIlUN5DqbqjyFaRbyYszq2ypudYYy360LDG5ciPZn8WGwxATqVk87IZFEU6K
BpT3YRl+EhXqkL1l2ATWZ43y4XTgcDtyRSC/Exp1bc9MRWn3eTWPXhCK2XSH
SoIfjHkxxarW/T+1ulF2tyGA8+6a/Y5R3YZyp+CKsmhRSUtJ9KdSvHKKTt9Y
9qF87GXOLdKArJKO8OHS2qeW+nRUs7dlQRo2C46pg6gTgOendYNuTZOSL2Qp
/B+I0NIBTr8tIYkUFwcFLpakfHNv+boY1CkOLMHBjZIC+CBQkQVXjThqEQvF
EjKDZPIez9cHrRABdhNmKFB/q4AW/b3QjlUu7n+oprfjprAEhHV6NqP8MET9
xH7YGTEea8mxjRWBqQjjgQCYTRohOnuNTuSwIqsbPA+YChqAM44LcTOyM06M
o+rU+eDq4Wn7h4rZ50UuFRr6m9AaorLD4aW04ofKF+lylp8qzvrWfD6IiIXc
f8OMQaVJzwYSfy/kIisMQT8npSzP8KTv/cqHB2KRPD5xup8OFTe+2hOqLKqU
1U6DrJfZDC398jtKHaQT1rsFIn+Q5dxcSYzQzwY6K/OkjFS0xJIKRG48bgG1
EgeGi2rogWKYWbIW4osq4iGIcodskWwqHNZIfJlTJyaw1UEM0qzMV6DfSH4v
M/klRkPTuQQlWzwv/GMK+KcZTPl/Ta+zzvztYPDZdsOUwplaAMgnTIrmNkBE
HqOZt5voQsJLRUnBMHH+L2buHxhKVBdgoJLtNwoJVw+UVrNrviHDyt3UZgSh
I1TsmNd4hf3sj9R65P1cUGZD+b2i87TXhDwuQZFEp16c4EXROguAbpCyhwN/
QQlXK2jeNYJ7K/nByGNEsmo1lCBtSDoheOCoMpQti17uc4hWAL9xckrCcg5U
u7rrefDgm0wQ26v4ggjcGKxa2gjLIK17jBlzoh9ORsTZ9us0WoOGPUiRPDKu
Z4vTKJcELuBumXXm+glwkM553IOmmP6m4dIQCggaQE0pasyp7NfKiAq1m5MD
TtPZmNwRG+W6kq+/J9uAB4Q5OYiSobsFmrIFhsZWIPbMwClsF0INJVjQCQbD
UD8FygqU99tONFNlLHQm7sHWPANnzvAM+arIN4DJa9eaisuMLj5nLh2gBREZ
ibFqZd6QW9NNkRk+FISzjCzzYT1ESB/3HmoYw6MvD3ApkdmPi3s8gZnWN4Ck
h3Q2R6cbhgN20XdRszjQGHYnv7UXJ6XQIYAZbVwxD75LViA3ZWkAqaEBbENR
p/1qiah8NZSFF5UVRR+/6ChxtUPboGgpsZSOFoEeAub6grUvQTe3ryitq8FK
lW9fL8G+4R4kaIKGwmQXkYdOoSUNcX4GNomxRdLZry1+G9evR8teSEWFlIlo
63DxoIG0cyexwJ+6KBgd7tMv93QbWpStMfUPMyGqdQddCqE4Oi9e8H/LssQb
+n5GFymApuPCeV1OYidvWyPD1pvU5vGYJ5BeXb0l7f7WuXDDDuDv2RVxCHZ2
UuZVW9ec50iMcDna6Ne9UCEyy+lnbh3G+BjY6geY4VH+wRxpFiJDBD5bHrmy
E3Vkn+1z7U/bquzS+QWrbzV1RrcZGbxx+fUL3dFgaDa4nWFcNYF/KAeZl+0j
VbwLP/uamdMOFRNU1yputHl9UtizsdeQzIk4lj3DUKkob9GAcAYQn05RNM8B
7vRBS82iMtFOyujvVf84lYg7fMyRVlDHEId6HuKo7TaykCITxpzQl+lqK7OL
mnFo6m4+5QJ6EJI9VxYYP9reKwVWqcSLLyb617nyTzSkPqYeARBoQgEJLHsU
NnYwltxxT+eRUY260Mxqmt0oeWiJbzJy0F8jrht4Bp/TMxx6qMeshD24aAet
kbYfkKaHpaRua4fL0iXMCAdLq0rxr0g2ma1qpquzAWB+MtmjX/0ex3RRW5RF
CU4I18vr1YH9ygIDHfPeTo+jC/v8MKg8pPG1k6jXmZrzkIZm3ira+0EgkxUX
FFTXU4LValx2hWk3qlC4Rx7abdfLNWUruMVlQXnxuK6qKsuhJ4K+OFhnEicZ
BJhvtthwteb+3+LuC8BAmyx2M+URqLcvV+UESWZ1Z21n8VluXVOV8Uc5XBCO
qxEb13ciVUH9iiy3t3oZPo2oPMp33Gvfs9P1EJ4u+BMbb+Th/oPkipM+YQYv
9/bmZzMdfRLSebBrhtfGCKcZ/8WPzxdLNp3apmabs+F/1QIFqcQ9rHgSfddI
C4z6hcoW+7xipwBSASipeepymY5oX6Q8WuFsFOpKWVg+mYP6OJhcE5t8h3sP
B4Pr0brhsptfcxkBZmecOnpT7p+ZvJmjsX4yAC3bkaqnOwMgSKjW95Agaldg
7Z63JO/1gIP8jLKN1DfRowTzlIxEW+oQSKy+aMKzHnh5tewjpQ0KcEmg4CPc
rwKobij9X3dUYjm1S2fo+4TniWatrdxZ0m1e3CZIFZ6wD4LQn+zBApODHx2U
BHE99XupNWW6D/JTTmwa8X4B+xizH+MBVi0UIi5oOaTXqTf1f8Ced5vt7vIy
WbZ0+uV0DKYtfv3G6IFwMi9JJKN0RjF/StcKm8ZtCwhQwdCtIFuaRUVaRhVH
BbYFCt5mi1b3eniCQCwDflp74rUiv+6Uxfx4g56JUBL88zcZHq830qrAa6Nd
y36S11oWrgW4UVk9WzRN9SKqWOT17+Atla1uOTIE0uWRFhJKMRXih3VVpvFt
OL0J/g7rulk1V2Ja3/BxNO2o5PxyN0TYDsJNl+Mt24jdi0QClJYAGVr26cKc
jvcec6a2D6qDa5v/qO8u4whvGB/QX3NA9lm2/FNrty8FZZzHPwTJckPGnAkc
gr3L4HnvRN2d6RH09CQNCMtYXqIWVZzTzzY0B0GLYGIx9Hv6b7bTMpzBge8g
XG9/uvRn2CPAD7J9SuMcvsclKVQ1KPh3DxdyxFYzZQsxSqgLNuQrtEOtOq6O
TkrUqA7eHj8jdTHq2B7JbSKnwiM+0mKpr/nQGmmpakWx9rnfzw5BoV1EHt5R
0bS69Wsthqm0deMlKnbBpU0HRO+YRoeHIeWBsqe8rmqahr+KChqZXvYQ0zg6
ATGfxEDMLO7Bg7u/BHFIdNGWFPpUnrrqFtp3zMLD7E5+z2RCuZXcnZUeGjl5
n3XGm+Ud//ebUWWkp5GoSRb+EEsEahNWgf/LIeDtq4XTKDJPBGNwo5UhXxDi
1rVe7srvsWqY6RTzA8lcZL4hhargcZHIS4PNdN2/L7BbGs/Whfi4t65a93Zs
uO29BzR0JiKqoqO85A+Xq+7hg7BFjuEgva5EC9kNjxZN8MU0/MlINIMxyNG0
tuZLJUMFbwR8iSB0LM1rRzRBhbUYILZjXwymMm4QTKyVtL6kKJRu85QUWf0c
sgffvAQ36jCXBL0h+n/Xn6p76HfrsSATkHZe9FMhrSmWxZOBLLaE7NBJ68RA
n9cASiqENpT/n0nudRovmCToqq1br/eCWtoWBV/YSdPE/cKA8JgiEDGG+h4j
gWLulGIBfMbkYmmH90AauhvKeDZmSbRv6h+qN/JBeiTbWo2KplFXqZbtAUP/
m6zKRByjC+x4vaum3lvIBxA+BIcSrQhf5U01WapljyWi6RTOK3k284qHREnV
MBo70+pwQPKDFKBjAj2CqVx+/b2pKAvrHrMg7NkKTyCmHf+4dFClUzair7st
4O7mwxe8y5dWp1K6LEkpCXNm9JSJP2dpyX+kBpiYU7NintwLfwjN344dSgzZ
uaNyyNckBLFxOtXWKIabrmmAOcIGM+Rt8L7mE3lud7It5n6dRXAQmVZEE60G
Mc6L7qK0jABjBuK0PEbqTLVyftL84KU2AkUHVQ0AI6K4z5CSk3unsT14cQLT
6HahG5YoxbzR3YRQ0Q1wc7FVrvmOBYpTr/ORQ6iXeAjG24uIEy8sPnCihCpG
meVW5LuS2kS9Rjs+2AkBXhJ7LXvxr3AXa7zargz7DyVMSjvUWf9idVPFUGy0
2UPzmiTRRmx3qfGaZ8wjvcBxJRq/frOWmzSj4YUMP6Zey7aFnO5jsKcquij1
ducbwQQoiiEh9mJst95CKvrEw3/wQE3qTA/qRGJwJ7y7ADcmF1aLp1luH24w
4Z9JaBNEx6lBmd+1NOc9HJ6r/v+iDxjjZ0rC3uidl/02fnTB/OnR0vu4Q+i+
3/CFAxOwqnRzt3uOvDI7e71UFSII89AUEuvlglGsMk+AGKgNLQtg+UOILfsf
NrGZaELDyk2a/xM3xvMVgWYwWhe8jmMpug13uJWIW1yBV7jC1JdE4/9dZXe9
KwsJV/PLoyTzf3CPTHBgkEdRc6rx8D8bYamElNXww5SmtjxLQ4KLEdP61rAP
G6Kx0XH37OYs0hqMS3iCNrv6uV45EnbcRk9us1YV/zCSmvy8NYf+9cLAUDhS
7uV3YFe0PrOAHtjl29JWj8kDcP/vN0uhdN490ZjXRVOAjZ7cpJ3MjJRp/ceP
vSqcjKRwb+qmAL084eec5eaC/eRthtbZZYXDMsYIPojwHzwBd6fRAdkbUc6K
TYXFgoXtPKvlyMhxz3LsraIfCH1HBhyZbKu0jnIJuEoTFhK8xkHL9NkgWwl8
G+bGGBejMdUqI6WkQbjy+a96AUQtOwD6Ew4PS4cv2yLQnlK8z/YsGUei89Zc
j/RfZCy5DEjBXtXcfShdSPJ7i/8zR6sdbWVK9a5vvPAhCer+dCDok3uBgSTl
R8MP2oAGbVxci7CdssSoldHsHDfRpvNZbK/bcHA2HAOTDu1gXsoGZZQ18C4B
C2+3qVw39nO99NkxFwBStTwr5vVd8oMobDOtJGNLiHBnNnu0ahG7qs7Nl/2M
3jv1Xu5fSnF4VotsC/RMAo3z3pdlzWj2wjm2PXKGq5tgdBV+XGlhU3+2gevE
TlVfrkm/1tjd+0fQwwirm2wcAJc3HhbwLKd69pOtLFvuvT2SS9AI147ljQw6
sW4vq/AK5TzqOimD4vyRAlTDnqbhfQnnjOQADTgKv9fJE2D2sMt/bMLeRhrK
v4/PSLB6Kc2nyIwEwzUSFp+gGlhGgw6meEYHytUJIDxDbKSs/qABGF4yG/kM
JOORurhJpkQO8idwpZuSIKIk0ihM3n+S2fxOjHSHOnk1y6inN6ly88usni2q
u2wwC12t6lfIBhAIQkvwzUgFEAFtrwu0EEHO1wo4urJUVGDpLZapZuUNKHTX
1k1JHtbDjh9+a3g9oBUnErX9QHJapfLYlfTfYFGAkLmK/EWH+Rkyx6R7JgJK
s42v/68X3/qBGUEtCT6O1R5+gbm9nQezaqGAkfkYoUqvwMvgHHYZ0HXpTTW5
R0lhltFt8vadYfFQER1X1qNlLgbReDIWL1pTpJfBlMRHvvjJC4fz9HbITb75
Fwxe94Mj6CJKJC1bvDsK9ooXWlRSucWry6XjR4Z1izRjWA+VTvkcbaHbHJ22
pxndfA33wzqVklpB/WU3ccxKkVnI8W6PFdr0CW7imbdPM6Gq2R2Hy7tRZJ1P
JRJz92skRV02sHWPiWqBTdU0fOhPAu1i3O2/87rY/auq4Ag5xLhlw3JM2VIp
56NAefb6l3AlD6rvarq4mV4T/Ew5ShwBN+9HAZ+t1PF4laUrv8BZtUhtnf99
6orA1ZT2IEWPa8SDMM6h3o2UI1TxC/UDWs6/ttMD1Q6B81v8vyMvx+DQvAep
X8gY4PIXd6jp9OkLJVqnkJ0zclSiCUl+5wf2KDE1e7KOaLkxG5tFsXA3anFA
Xb7MXoCl0CuXA8edNuxEh/i1d+PC98KB21QGP/sfu51IfvZgYgk8CLEiNlP6
vzQToc/pAr+fwQWuqNXBxOefpeLXota3CbpXS9gCAHa7VyYmfisfiX7KSvU5
EPRJ3/+/nW7zF7DqG/Ij192RKrXYKlCxJrWg//lTXJlb6Ky7RoUvq5jYdopX
yRzYnFlLaGrFxoAxd9PqImSNGTe+LAidPym/zotAzxPLxWTYA5+L8NfAk/vb
TGykWqcl9Z14kwP/Gwv9XIm2SNBYiyennL0qHFuUpks8twP5OD5tHsgoggzm
s3j/ZotAOC/MzV5d7sIcz1OFGLJVRqAYdfLl+dYn6l0HMRUAY+6QmboFH3jk
FyT6ULYJbymt6+u3ZgglqiAG/Gj+j8c3gIyQJ0C6KLa9beM0cGAR7TH6leGO
GD1LxGsib1xUlJ7rcqcVWQwz9AMn5s4jslFSQXfIJKC59cX3+yRWtCHD+R0U
daLaE6mXIjguk//JjKu6S3ZYiJAqB339x7kZUObBp/jTp3xd9A/HX7sYPXbI
+jKNMasmyqHrxwOoseov/PF/Fdj9697nNTtXwK/NOzEcGfaHD675QjztONVs
vUldp7gTy+PWw2o8tA4JmeR8UVTKh12cp/2yYJnb5rMGZbQdMxHrdzHLOvNP
VuGhOLLai63SFlUsbrQyjYWMS7xgPhYYQU26PM/kIJGDaoluOh52Ik4uH98C
DY4IQMJFinNYfw67EFnoxuh2dGFCDcnG93zncVeqpdDZdEuyeN+0flpXBpIv
PpA70pDAa2R1RAFSRFX2hc6S6VFsIzGJDfEtWTHKezdMBoJLzXMEg8JqBS+c
uxLTd0wa3b9zjd/Q7jsVA5GM74HvmtTVDZqg5hFcCJcvK47nT5NX6mtoIoKm
MvDAaqX2uKXvzEQnMCvC64UAjxkntPLwLYnR06ue43PaPBPpMQWcUc7+OAWU
lzcXT3HFnJW6I0E1ltcWQVmvqsL8MjRiVjFICpxO732OEbm3ul2Mp6gUleOW
gd8lXnfWyYMDRs4H7ebDrz2VNdUux8IoHvAlgNwzkk1Y0ae37kECFnpN/BlV
a2+GNjwkYxGt9xXJImu7PoqRTMrSJUe/Z1IgPW5iQRUrywDi6yqWYaQPiyBs
8rEUpTsKTDb3I0GWU9992qXXu2tSBfwmZfoQM5Z9bNGT0I+ZEhXzZhHksZs2
KVV2woQpwjvWIVMIiXZeeyrl0wUI9wfXwCbADwJikaVdBKgtS4dbOCqrwdNE
Tk9vQvxwvWp6LNvXog1UBgm/qiH5ok/jDe7JUtoDQ78i45ttZ9mRy2zbTDr4
zepx5FHYYSpO14LJJyk4z82FsUlAE+SrO9JijGT+JPnF4Jvc2qt6ZdxwcM6C
WIvo6T5v7YLx+//IL3D07f9IR5Gd2HesQHxy6i5hNOp1UQ039gmc6tdMlMjE
3+bE3w8n5AOvTj+5l4hMoZp/D5BOZi5OjOoHiQKTyuuZqn515kiabWPleJQ5
25I7JzyveuEelw2h3VCZy2nUE1UfdqNpNuF1jVpAfvPBXG5ab1QrVkElMjnb
eYzl4gKKrwqwJbwsdQr4JxeCMK87RvPl2d7OLokien0XCo6h1HM9Hbz4Ez7a
PRpSi5d7/elpLMPEUi4lXyyvtNwn7Ec5YdVZIUKakEislCmglwbyz/Abtf0u
VY+uO/zUvZqtC5fr3dOHSzEc7MqreMF5hfS6sKYPPCTmY1II2w1CBrgOEap8
P6oZLEKCjHvdyNZg46Nqy4IHEAFuZ9yAFT7kE3tGG7IjYtYGMDL4ZXG4z9UE
b45Raz133pX4PUhRGOiCCEP7x1neQPDSMsJkYoBffOE3tGS1kmZnjreOWBGy
R0YtUnKx8KYobaycU4HKjizlP68bvI9nFN846Gzhqm9DsDfqQICsNxKsnsZY
eDjtl2qwqRRLYNn5KpHbZjWB3GINJ/5aqQ/pWHYfr/82OZRFH/sbV7iBfvV/
Nk67DLLTJ5dr0ORAFmdbocGorlKibs07PqhjdksjLBXawGJ/zrribOVluGiS
ktPkWwJF+vYuASUOb29beDQP33YUjjg6gByNm+A7ypm3WpxqLPG1dv173tsz
nVRcITgszf20uH1UYQBns7X2l0EgGa4B8WlL9XJ+6+Ywfr1JJRzumqE4Z4Jb
nJ8qVupOHhzl1/rtgQj2jMwVfVI+hJ1nURP/nIonyXJi7OXfSDjjq5oaU8dl
9rEcWg57kZ5J/yi6g3wZt70xqkCibFEhojeL/Uzv0LQd5Gi4Tk0C0OvxFRcn
n9idg/BGCuNkW3tOIEkd3oup83dsCP2wDqSBauSZNy1T6w8/yUQBLD285WiF
Y6nDYB/2II0BCKycpgVdZHiiqqAEDTRczQrTzUJx79d/65xb/cf2ltozeQ7m
h2mcx97e8Uoa9u3Jerf6oIVXHcmVlMm6TqDA+vhFkNFw5NZNZuFQiFtnRbro
CPgtqGtvM4kQmGCq4xFB3EubN2KJv9kR4sC2dqzvYWHUPU/Wx+wJYrlpZ5Or
qAsrWKBPyKQS2GDjQeWgwGGyJe8XUqqpiLa8MNbJvevDZxOTnSaRd+FLD7o2
8qqoPJYKtIZ+67w6TOoyiQqc/oWmI7P6HsY4bz+WJ7fHVdaJdj11xawU4PFW
LN/3/PXarz+4w071Y9czp1Lh2B0ZDg6TfHWX6p3XTKe3jNLsP4rlCUKrzJBk
Mi+qA0O5tzseigDjajm6GBhxu7t9ZZiIjeIvg/BF3H8jrYCJbR8hCm7zls6E
v58AkRs9iBNWwfacA3xgMNRp/Y4DmUFdwIIKLerfw29uKQspP66AlqP/PC8c
b5xMV95UfWSWjZoBrkW2P7Q1HQtMuiWDtlKoBu+OHkn7jMgF3UdTsGGOBb+1
zGV0/PKsz6TmyqpCNJYZl89MGh2N7grGK+AN6lrkHqkYHXVfWabqPsBiRvTY
LKh7Lcq455SZv4zD8ke6gHQbmyRBvm3Ja8YtR67dTw0V9qVd7tFQVzqLwnrI
bZXz+1sJbQni0PPfwqXTL7HLU7Tltqi48aR0eIt2N10Rn4hWn4iXKcLPm2RL
NF5Nfx6LrgjTq+h4lmBQLVohL1W3b1wp19zdq+GMd+QLVI+yWneGCuR1LBzJ
GcQSIbMmq8TIt9jnZYGx59nUWe9UnYuDuW2jTWZHXADLIB6BImXsMtq/CdXE
t5b/8ZC1R7/jKGeMPcScaVJbttn72YyHjbV9tBYbCUBr4KlAOK9Whu3rYPDl
tpRv9CUVkc4rJuJ1kzuqZSRzWyySDjEmcDYcRJPNVCJ9V77N36AGrXJ0W3MG
uOhWiVhfz5IcEbJ6l3RVAy64iSWryZol8QnvbEUsv23/l2SXioxLKzk9+QvA
uyrWDk5gAHj1dSMKP6tMgyPx0Yr2GtfdNGJLZhdP4CFjtWqLNSgm3l4WcT0i
w0tUcHEJ+2Edsi0o4dcktBRFHjOAAkfFYcktrWECCbB3fZE08Usig8Dv1kZK
FJpXFtfQ1ch6CGm1azfDSu3mi5AfzvY7GBREWAmKuterEDsLwXhMB5tYp6Ti
fvt/oSHk8Y85BgB8XjU4VhOf5nV2hfA89qv4SmhH+k0faCj8fxzqht9THwgO
8rYYP7CblX6wKtFozA6kXPZf+DHvrW0+zrxJ+St+huLRBCSFHV0d0Enx/8AB
U7O9AWGYI7uqPu7vx6s3s6cswGrFc4wNmjld9g3uBfl1nFlXTChrqgZ5z8xA
wIqY1JQddAjUPP2pjnfQGxulEwCA2T1QXJ5jyRV8xnjrEjNsg0rXPZQjBBQC
7FFm7nmONFJL6c16OOZ1iAIz+4ZoRDRZKRh2UIisGwxwqyDOY01i8uwqRoSn
E8z4FhGGFCyIjA7IOb6HblGtCHWuV72yGZ1Rr/NhZ0i9PuZkSny7EiNzK7gp
zgSFvlvvVJzcPBDjnOECZoHa+UhXw6ecwP03KA33s7Yd8nLL96gIvoL+ERC+
SsyyH1pLQhULB+c2LLczexEbqbNtf8yJPcHbUFDuN2EFtyVSVQoaKqJ0K1hO
D9Co/rF67gPsL8ZCFubAyQz1hi7FIQNd9aKMqkNmnl8nmlDgTIi+JCa1GHfw
JRHISObenXIILDHd7bRMUwZofNyrKhEj8DzpHrgQJ7WMmw5tuG1D8c2KSNKL
tUVJQ4WSqAbr6NoNT75XdZXN82Tipk/Q3HYJFE1SzSsuzSPeKc8hljwIxSGX
Izu2y1NNxfXT+DV7vvZmCERCwryuTVI5D78j1UpdI/JyZlStT19KVWuB1sX3
tY/cukVFOKfPkozJ3V+2gHdG8nCg4MzecOC31P3atjBVFwksNmkGV0TL4Qa+
ExAhK62dsXN8E9b1j5I/QNTSiu9hEVi8qVWOEDCyG0Z4YtFUTGvRvB1pzCMM
WJLPXRM9uLaGLZynsltF/JW12lcs3JJrtmuUnlHQIpqf7uK3fCEOJd7YIIuW
hRHxQZuorbobhS8pxWpwTd7zaUkG7LGym8ijh9OnxwQIpapo6E1sxHyxyZUj
m2dVFCimVM6m2VURsMzLNrKf5LJwgTfNHuHEj3Gd6lQ1K7/ggwtUarCHCm1j
cf9TjJK6d6/ptScFkCS1gIO8h9aGMCKpNC8XwjFCcQVI8XSg18eJUUd7yXE4
kMedACPinHrSTUENfPSs82WUaTvXYJrz6NM3RKKLlSiQo6BN/UDqmgyru9f4
QMmyZQ8gSmRASpHslNll0xOGiqrIM5Nd+8FKZn2mtDBNcxdauswDUoPET6ep
iXQ3C8h3+FKWNBVXDe4ShOBcnjlL6sD8X+eefnpHhYRw3z4RtfY1/SyE/eW/
1J6kAZd1xDXmU40pOfgH78u3jUYNDjLy377G0goJe+Towzj6DBgYQGrsbgOK
1ClT2HzUF3LD7JfAZXIgTdb/V6E2tlafSSt0Uik1P7nFJjbsOnWoSOnIi2lG
eaInn5cWMSMMQOTgEryFnvdyQ+AZatAkcxhxBrMyKWdiWp8a7fjvneFHuwzk
Ht0TxRYUm92ecMsfsZWJR7CqX0md/10tuZX4TYGiuzchHOGKj3qlFo7Hz3/+
pGlCNSg4D6G7S508wAtRsSTdsTucrSNtj5Kwyv/eyZFfFqueDn4DISeRBtIX
EuLyltMC6bdgvqit6B7uSNf2Gygd6C2eq3MumejuRrV6DMETXVgo+pjksAZF
M48CxS/O0mMIMYBt1rALUa2BU/XQtcXeb4AyA+kANJbkABnCeKNZSuOmrPwb
WbBSyxvxdiKVeiOR6CqlWq/KmhORSEXRr6QmHKlgA/AxBuEC1wKO08+HorFy
i4NwRmQZJl2szjxMF+SPtF161egdmwG//D5gxKFh5eHbCOz+qpfkhjyw/V+b
bwdN0DG58odXR16D0HZQlBQpLX65p46bGrfPwtjqDIhMhXULFo4MSo8K7ajy
ldKL2TAbn5RWji3Xr3wdUkMydK+2nRV1wQrvXv5W5EzEXdD0SHJm906J11/A
c6ZQ/vf0FSptuPuIXQO9k/DvsxfY8wM/nSmGYy4NmxNsa+z8ihKuL7inrvQK
RPxFViMUf+TC3c5u0EyPRilhRWbvL6xCFF+ZGstejiGmc4NVEQUUtCRhkE2W
QYXWljhnDbPy95aFX6oD1RSteJhkygi24szmHUtkksojHBoD360F6bEybCqj
Kvb7MJZ8B2TSfK2Ujr8/SJAGH+coVrKMAd0ZcEDF0b0G4w1IJIGMXtZ0bQVw
y2N3lZ8emQw7iQx1wioL79X6DtouhloYrI/HPtSgf02LeLV4Q5mnwLT+tf1I
pGx3ePAoMqreomAa+Ij5/jeNuYqXniDfSFK+uIQ3O5xBaGjr650DAVZqSvkZ
UFlPdekEieHy1BXk18xw9zF+h//RmdfgH/tMykYr75ykriMyyOMoA2NdMzGD
xO/lsifd7xGZBUb75P4maCFXaaSiwQ3TQROeOMxx/dkh75T4JVBKsutJ0byp
G/20xXwFmRajVYIYyrzFGDZg29aJXsf/hsQrk+2PGfSh8CkDmUR4z3tg4gl3
nyvlgYElz6C7krnHKPcEQk/QehQDBev8YxL7T0HMaivxRtZZEFgI1N+CaUj8
3bDMmoEvsdzFBx1WwGgeE9luM7L7nm20pUcZNIjlh/q+94vFtFPcg7bGvE/Y
VG5MMfbHHu+WPHS+T2Gsvv+MfTAc4eJOxzBE3oDT0tiTwMv4f6EUGy5B1xzj
IqkF/SBYw5nSemvceowsR0zY8KjOLex13+ifnG1dGnQq34UM0219N0xkvwrK
C60apgDEZvOIG+sEBmaXeAgp1bKLgNTRluZ19R5c6KTLvzgyUm14dFiBwf17
zkJIDEgbje3iWQzyYTwqj+jTUyvMkLE4IbJ64jzLTeCx/lE258ajMSQogoJD
BsHv/yqsD3wFTatLSQAvnjgX9GgaN6WTd0+/ccfQjtBeGnwQOAtehW9mK89y
5mlxELdFHR35uua89ysgjSpPK/VX5mxT2JZQDc8pVLqjs4JCNLFX65m2QHb6
BkTkLIMCgHHsegXZ91R9zmJwhhzRL9UBpHFx5rN4CvkjkvqWx7U7T1h9k7H5
y9cRCvGcQiuf9w+Fp6bJKLB/iLZiRuxXIVKQ6zKUH5YrIrgmkE5CaNdaVyR3
6CYvngwsFYnPqoAxAuUaxKYfakSvd91Rs83o+chKQPGHK+7xmqT8YMyJlo+W
mkNAmE3T7BoRUUyq/4dXDQ5lVwlatnXK13tQUnqb3pFutfT9BsIu+xSJ5H+e
11p+d72DkruzSgbn13L4TzWtrpmFVBdRTfavrczPGTqG5ifJS6YLv3T8/1oK
xYi8KgGXvCCBj1o2cTbjNpWDdPeIHrRJmL8QM9MKO65BL9vh3qUufqL1hzr1
Dfjtk7iVY4gtQY+YRqcwUiTDJ66GzHZQqMRiIPggYY5gQ34IkI0jfgfkS8ul
Z6aI8VhdgPh3FXSJfVTm+PIvgW9G48XLx4AUyRdDJU4Zlk9wsqQ+T46OjfrN
eLPgGv/3hB0YevvfwJ2W95p2wKFmcnc5adkNtfHoIVDIMjkaDQOPZAR+N7nF
/6R0ujtrASLGGAK5aOSpzBnEUU/H99gHhZtjetgPWvAbYXlTuyk1Gm5vEmyK
2tcrpcqWXRuNjINh6Y5ustqxRK0U3tMzlsLw7b4j5aGh967bi7oqQcVQ1bBi
iH0t7LUV1/lghhxTGoHeAHmPsm7cUWEgjGDptmoBmvMj1VEBemNG7f/16FTM
lNzXHVXhf46XJfs0sizOqYoaTt2W/AJ9URJydiqYP/WF/jYGRFEAJADtWre6
GuAF7E+pa+8weJ3wWSSRZ4t6/nw9kasBOAoDdxHXE0Wq547RzbMxlzfgvN1O
uNqbOj/Cuo8Ve5lV+RpivJnr5/rFhok3fN3KL/h0TZOyOJ1w1g7XFc2OJLoe
8j2DM+L39SGGTE3EeI5is2EuhhXRUT6u9GPmoFqUDJEB7xIiLiSPCMCcM2kR
KPKSpuFTAb6y5b3sYsnbUcZXFpZUMy8UA6rVNpNXEcIoSfoHw1vCvNZ1Z9xB
vKDDCqdK1p0msHzyVKnF0IcNZ6ShCFfNtyS30wkZ3hf5avRJ5ehdPW0L0UKP
sKXvSu+jkbCsqR7Sls3nUwFOcB49yfkilqXrGkEnvPjLBLCguPhcO2g7g9nV
d+ct5uMFS4oU1G6esXn1yx5ULNPsdBBFMLgHlKXhduZXUdDxudZdsAPbGxEe
xbxyl50aawMv4WTdRQSRgKhHBQv2unCrY0uLM5YA7EutzqKwV1bm/C46QiPv
86mUclIv4SDjRhwIBuOxUGb8Fqt8/YPOUXGqGI3BrsOo4W5+A1X/tq9t4ZVK
BLEkkCiFvcJxMc8X95z4IpUx/GgPzKZqKy8ujhuQv6fc+NNMwMylrH/rvpgG
50F4O4PPAAyiFsK7f+Ahulox0vchp1hIZnAKWp2VnPgvoyRbU7Fpm3pmMTCW
ueFSSOou4lO5Y9AptTqdauDgtRHEzWLapi0ebyM7OsONCyl9HRyUE16gZcqA
iW5kwWooiA6rYDwxwVogysEF+1rzi8/ksIkNNfH3F97aM/1qISLp7TiPJj3F
m6JdpPV6TB5FsIkH3fMlktW2qaMrbrRRqOOMNz+IHeU3gNe4a17aTtm0jQ+Y
J9rYADRqwzqBAFL2CAQmg9v00pAr4aS3FrdQiXM9FI2vOF5gohY9y9O7fr2i
w2QuO3oPDDuhRLDNBUGWk8WN7h5phxOkn1OQN955Ge2IQLVb7kgpbG6nR4W8
IZLxqUmD+Drw/J8M92MBsGdrsNUaPr45obU/t+4lNM3GoKd2DYihHDNANuQX
AXNh6/Z3CctuCiVzwvtF0O0+nBuRL7bZzET7tmz0LkUC5sss0kzNBFXi3uJF
Ud9QXjT8GFJj1+4s0x5VWyPs96D2+Rg1J1a9Z6bqkTxNkogOEClYFjrJxUn8
GM2KoPVnVsFVjhNRX2phKResdYRI8QjcpHIbV8+GT3HLsQY2DpXLODxTEz9/
Y3zBCM1WX7QmNMY7SrqhXZPduu+8XbARfhAZVDowihl0slit81LkIVV92QIT
AzT3sDoxsmdle+VPPxeI34ljPSKZM1ueEQ/CN/FAS3vr6yLlEjgHK9z81B0I
D/WyCp8jDsljId/xZWH0pzNCv/+jn6Y4+8i+CF/a6bRoSUcUmMd7yuSyFKCl
dn5uduGWFEeU/KTjCr5JED6eRYKisGHa0Nl5CDS4j9tGw0NTJlALyYD2uuCl
tX0Jvt5MKUgQIpm9aMDzbCWidJK5z0IwLFQySbNbR4kxtUAxIgc3oVsnzUP/
+qcLAXTw7QBDatlNZ07/vvXZatIuTd1GAA8pSfOMYcJpNCDylSMTit18BeiI
1LevqqQ0L4V0zDnGVoYlFR7ewgTxIsRDt/syycWixZBIncJBhIavmLgmK7qG
DhrRIlWRo/4JHE1UfwDy4OSuB7UWIjt7139hZwGR2cGM90t+zLSBlCsReeLn
NZrhf9S99fM6bOdab5cF83nrMgQsuUivotF0ftLWdIZkYBQyAoTuJP+31z1x
p1I6w8HXf1QAD/dWBBxaXX5CsTzYjd9ohCR5bzfUFqhVrBD3gPFpvu2Mmmh1
XuVB8+MYn97bxQMJQvysptz+0uvEADGJ61i1Eqz/bnuMsC3yhj9s3b2iQadL
aEUK15w8lzD1v/qAu1hFeruv5Vgl074bOvTzGsnmWUc2vGlTqu1yfxIUDjLo
uAVCPScQGGrjx8dzG+7jtAssPldyMFsDJ7V2LGVPb7H335J0IM2dWqzDhfS7
P4KPbjHBWn3tQGQnlt+EM55TQzLG/lLgk/kB68QsjKXLW+gzh3VLUFB1M+wH
56xVxWU2jJnUaf3UgqwFW3L60fK2WK2nZEMjd+POsWcaHYaN70NBJ4fxgZ6d
ZWLMN5rYmduWRU1kPXy7Z9leKAGuS1F7lx9t7Jce8inSo1KxPP58TP6oXD1f
nWDxKySzvb1BaqKURUCPdDtMFvcGNu7ljYckHr/aCxDv/4PYhfmXTwvZVY/+
wtZyn7jnSYEsoz+4Z272r3J9hu/fwCqBby6w6tS8wmqh6WhTnZqxa9O7bSbx
QMuysD895CKGQ3UCqWov2TQMu/pb/KbJmxdCVC7zVvjjWOm5iLxKz7Ofrysd
JkZWLfri8puiMt63s5g9Hr8vzOFL7U2/qYvP3uH9miShzdZbx3fJMN79Udl2
ApPceGgbRkOum0XB6fUeNTeSCt8/ovh58tqSY0K2WIU5uGmSUSxntIxjU2jG
HmZIpdYkw34n5swMEF86Uwas0QE6aOJn8j2tVzUfiGsEeZ6ezjoKMAABxuMJ
g2VIOPGsu/HqVbopnb4ACyfaD7/bel4x9ahe84CVO/G6pWM/2fYr36GEpRrI
mtkMLyEQY7ySWh9edMmBzLwMWjMvBrcFK8KONMSYJPGtH0CO2zYLogUcxDLo
1J69Dj6qvV01NqASC4L+PXvohzG819ujcIJWiC9bDfaTnVF04z/7PkR6ZrHZ
334ZLyNeALTAmbqm+Cf7lITEKiX2vjXOPOR7oFVouU8lwukRtH9o1T+maPTr
TPlKw5K8LQ376dCs6VYiTaHMBq1DO8wh4WkH+RahQET/gudgYKcRH9tTqtG0
1SwP7XzwosP0SPfOoGW2vJoPET3y+GFF9RD6H6/AzWMPB5ZMYAAdEtuZznvM
/G6mhmKsy/sl1hSaX+qSuKhxqWWAeo1m/uBveiBBmycoaxYO5MfgG1XjtSnu
YZN6J7uNj9KQpjqqIHZAcInFy8F4kYA/ByLIOlnzTHcRLjxfFkkiw2/s12tp
E6CfG0CCXQd9sPIp9+PKYbXHSPLXEoUS0RSsHtBqAlEtR2J0tGKtr6/xWEMh
rWPJNuQA+IxVHm1TpEvO5t06CvIFNxKkAnZcyfPo2Ly4BT1nZjsZr0NtK/bM
s1NffWXLsylYhDyiHQKmbwQrKZb09CAmKHFpYdMwfcqW4+eRxlFs3MEr/s+G
8b4MNs8QzYc+ZewcuZRX0duiIQgDbuwTML5bPa1PCPbFrSNVdHNFRinvAZFe
jdMMvJlFxkwU1x85v907bjn7kpJZxClU6hYBedpkw0ozWC1CZVNNNqM9rDiA
/m2ilIFBjh4/nc94Ozua63u4tx6ablqgcnjCno5YjRMK8Q+UDOFiGqjvCU32
yWOGWThuFRdzYdMgWJ5axLJAqIQGIkstkPt3pYJwUxrbhtOraUMMt6FDkRBK
//E3HWO4ar3Q1iisNAmwgNWJoC12cYya7pbw+ZMc8//8l6BMOTW1et4w9YMI
ofSLixOeQG4Crcgx1A07A5e1MeH3W0ZS9y0HqAFvviklm6XKxBj5QUmUs0it
FB/g3XjzRqEo7EyfLLAFGKnR/7Dg7ZQET+1rNgByOGS+ZvmsbVEXXQaOzSKA
Yma2fOXwbz+Btc28kPREex6/LxpBCjXR5i3BWXsJXz8Rp5Y5e2XZBGH7O9cQ
ac8HhyEqDBPCmVA6iwLBhYJHl7NbjibE6JpuMBlh38UWpN8yCofn1ILH3NWa
O2RxBkTGOmRVwzTcp/IsUrBzTTW4VgXIgPDB+fGCNLaWbI6olSlxDWPhCmp/
NdJ/cLc54WUGPRbay166uvtHWeT7oOgsl15nfzkhTMy7mzpaXtHRH9pSfDoQ
HbFOIt8VkXU4Peqq5LpxyK2pAjAqLoaQQvwNBkoZZMr9rmK4zL5q/oWbaQGl
Dtej9LCAqVOAFdcEu2gQ8JGwlMUazJ6idKCl7I6if2nRfeG3IAT9zPK7F/9e
97MczFu4dORAoHL8cXXSj/PS+5nlcmTBJx+RmpGYnhT0RpRMBDLCMutuz3wi
Njfskk6YDPy0quT/ZPfTukhqaWopUr+rVoVjNR3AJY6dxNnhBa10zL/S1/33
ntFBZUwDuxcyseCyNUIiQptTmranrV84THYuwDU+hHHQQbiz4PkNe/yx3m/d
AF9WykZwwQ09Fw7LeWRSc+DIqjpzLMtCBd0mCix1AOUn0ft2MJPsJEWvcozl
Pmbab9upkIE0SyOkHVYO/QwqBhi4fVdOkRrP/IjrR81ubDzYU1GoUTBKIdst
Oi5nB4I4/HObpkiHmcC8Ery+/wM9CzI1iiiJwK6XhuLXdz339TxSuHL0FRXT
hwoP6HPYCJwwUap3178bRDlOWwncSCosR/NMsUlm3I3BRQdvacZLtxSPxYpB
f1jfI7dW1qCHc8KS0dNdvPPVIer2Q/CiF3pkWuheTaW8dH1o3ddNPNEI4Fau
aqjEzKRYT6znrZrqc9nODUhw0k6kuooUUJReBdfPGwMuDOfcAPYOrBPqAxjd
ZTpumCtbc/HEObRJDA/hsJtppwhhVEi6XkgriU9rz5R0hwBh8al0eG1LoVqL
YqNRZubmW/oK/J6tpp6KvsfKHTo+KVSVaFicQ4JzPMY4W7cYei1/OViZeGfs
bu5jYJLjWUrowif5xmkFdjZs6bbrWARno1j0fBrHqdHmZMI7Bbk+7pfHrgW8
Cir8qYo9nxG3Qyn5WGfV8UKNxFhXoT+FQdFm/ZZlRZLDHi8HvHvBV0RftUgT
y1aI1e1FsjyOURsH2cC1GWu6n6WUBjzUfSeK5yUa4X98ih4SX4wIVMjQLNbC
gTgOMgTh2ohy+rTRw/Qk+Ngjo8T3VNSDttE9N+lSM/DQftH6gh/Lz1fIyuok
HSS8/oLJJpdWXHzmDoBA58aM0JgEeleDSHtPxCkix17Y13kNqkZdPWJxq3iH
+DdMaTsGDUdhJQmlbAvxubUqKFW1Qii+VaY2YdmyhzspVruey/pTVbzrYA7S
c1OGy8n4YDE7LhprmX34FST8Ehfb4cjELE3TX3dFaK+MFofdoR9f8npq+J+b
/pITjNtfyV3V1pR//icZm3Ut0q6Lgxwd7NnLih32H8Ai16DyTWEYH7/83t8w
yntQ4wsMFzH7E+VTuoHYt6NocdcyHtc86JUC3BGMqulv8qyPvAIeXCc0i8QY
ybmM6TABVNiTphJyFwMzemPpq4X5HOggJI5PmBWz+JkvWuzTwiyXqvT8NYTg
pHrt8cbiNMBt+u1xQblJWmBB4eoObyp/BKb4Dvk2tz8TLNGP2DTmHDz5IPEH
ic4Y3xLGKJj9zwpXEKX+2behev7ont5JxhOgucrIVVAO527biEvxsjFWrS45
sUeVtW4Z6gFiJL8gNgZnb9iUOCHdWFoRTuEWeXgWz2SB/suGin849Ly+eBcH
FWXxe5F3Yh7etRWHe5G9tmoahI5ralTWwbe1Eu22HL39+wqL3yf4xcTo2osY
y/4S2iJMVkkAwS63GJsPWTjtJGBt0CK+RkU01Xp6794qJnDuiMn2YvUHLBS6
ECYZpUk3bTLHDxMH/Q1eP9R1Dgy47DVKNChNxbeCL834M5RNy1QkEC7syq/s
B4YBAA/3EmU3L32Ryv/YWmxUmrQsIsHCNj7jMakWQwsUdZ/6UZs/PqDGIo8I
xgobRS5gwTOeKnmLBrF7iW1FMkNUgVWtDZ7J55JuMRtIoh+pwXahRJ2ToELw
f0hVVOJF9S6h8v8D9ngTDct9mapRkCpztEzzqUffvY5VzdOwQyKkGI27EL0C
+At7dBOJxgYOaOTEGhMwgV/cmXbhqkDQ/W3CrelmevMqELUw2aFB3eUiFpoq
mt8Q41djV4gmnSJh2Z2OQjx55H+/Gd5aWuN3LcShOV7QFOB04THlw/8ga/zp
xXMVpC6BtzwWDQvPy2+mXM/Da1Ke83VF16nVHSec3HPVlIE/G0HWff0EUUcb
LJIpDobEkBEmSOT+1S6bWzgHleAnnJuKAQYYJiZFE/iyJ123zCDhT5r8sApD
KyK11qXtgbCMYS6Cu6pFbtG9rv7Tu/1ILtaZXs4X3R4AVVTSGq4v1y/WlAsf
bh/cpqWTamul7IyeZNlRLyP4lMAJw2aM5hrxc7INQJxFzCuMlsOCi+HkHv7Q
TJz9OPMwy2Vf6PnX9JvRTZ0osKovfOMYjBgN0lJNK3HU17WQzm/d69y8bP8D
WCLDdqTrv/l9STkA2qScRvYy20yJ5HkossunAyTsSN0Y5r6a/gBEE/ATFkuY
bhHSEQJxEJt/I1yJSOG345V2HcN/KwVy1q+pe3OU4tqSLNprjNg0RLJ4Pg26
TiMqWqOiCC3yh4UCkRfjpwUc4jIHUr/AGq+f7RbpId+ciQD6nnjerK0zwCil
n2VfFAZwcLgQ+nUlul/ov80lpSs1hNmlytYF7eIYBZAN4H2nLFuWhQy81CXZ
N2OTRdDW8KjMqcKraFuCV02MVwMs3S4KdW9zi3cKQcr2CNj4Vu50416ZeDUr
tzy1m8Ls3RuK96WaALtXDteqZ4gqpiWNG3VLUDzr/0cR+PmLBgfcemEhccXe
4KqDPoIZIp3ZaNImkKy9cG2b2hWBvUnFz8gnCbfqsfHEAlcU4sP5DGts6h20
RL6BwP2RsbEHdwJzAYhPcWalg96kBjBoWxCHcXWFjDO7G+topQ6Oh1zG585/
4gpMR/eKy2dJQ/mZUZ23XsHNDVM1NDDXx7cUIfxaqV3bBMWfg2TRLH3xjziE
e3s4ogJaoP582kA0c17PmlDQHo218NrodN1RniJFl8xVDBsUvIy+Ic6FEClD
G8qccbqVlu8KHfUUG7uzTgwY4Y+LmTLx26iJLJOmLMbCAWNcMBXgfxjZzCXu
YMMohFns9vUAMSlNZbk5S+x/YNygn4sZoYh34kVWkUe5il+4O3wJcaSkuFdo
7+yBnnrc0YIeQ7wZ/h1ZGjMjwVBrCc1QdnvOaZGbUONam7tYa6U7ywPdKj34
aCgC6JoU5sGv+wRuPv877LK5aq4smjsEmxcVG2oW9bIgqZPWWabrqZHpRaHz
QssDNfqs7emeyrqDa+dmLVHNLwaUq16dxtgMxrdcAodZGJa+U83iIx+SFI2n
zRRgkHkJkPAyXTQwUCWeRt2VYpg/2pWsXrKbvul1UYT7eSOmt8oTtzBnvonT
Dhn9UoSiiO4SB1ojJ5S2+3CQeJcBoaqq4Q13BKPznXBL/x4gMNyuE0iBho+l
NIFPeR81uCR9ZZozJhIcHsKn3Q8bS5E+SBfRKpJe+AU8OWZE5expuSWuDI7I
kiAiX9HCztqTM2If2I2Nhp/kfsgNEnPUzit4+aKmb/78Q/NjkXMN//CPXJcR
1nowioe0heJ4IT71rmCwcTl4pX94lAPsydnRiAVbZw74FACQhXAvYlgEHJdM
DmqgGeVv8TK2b9e3N+lYUGX5l2HlldvmsfVjOQvNHcNTrYG3C1MJLETzRpsG
rrnLTiZQCW11APStozWqM52LLeCJqIpRLFzLqvTmE+tnUv0TuswniM1QnEw8
X7NKrOQ4R3s2uRTiTdoXrV1SqmcIA4xlRq2H5xMpj2bxOxNBH8lWi6FvS+Jp
C/x3IOnshyaMtdIT5BTpLTf70+6wmZ1tIcMxUkU7JXhkY5ai7ozILieAzRZF
gtKw5E6uVVdn+eh5bhGbFEWOOsaB+LWQOTAxWsQ6pi+3fnV9KaWg3ej7R+yV
7f+JNYvD+5RrBVtlBRrK6L+8qv9bLig07p1ey9ugYXVIFu1HMmMwDC8MBu5h
xyz5XlzL6sk18H8YKot2mIe2GTF0XxjeZGn0WvvQ/e6bqzKkhU6ZzlAzI6n8
5xAstKpavYRCMaBFKxqZ2mwSePpP1lZRxW7kBOJ8osmgxTi6Jl7ET/blYVla
qWPJJ5uXHkyuaN4L4u5ir8hCfzwCnXRhjHiy96pqrsL8vYEserxBZPC4hJWU
Phh+myIM1NB9xmF6Fvfx0LXwJHZmzWqCS8eQ5fG2MUBlglG31dS0HKTq4wXc
HNH7YG7zfLdDfIh1I0Qjb0qavbIQUpEG57hopMOtYyr4K5j+6XqXbC4S94cJ
KwabSeZonAHzAc0AzB/LAjPdFP5csEygKrxme01Acb9CUxVvekOm8uvXbj4J
VgbD9R82QRgrr+9MbTH9LnFTJM51kmYVLDNCN//7bHniYVCGly30CUKRB8kT
NuH6fO9sdIdp2Sm2yQ+127ujDE18IfxesD7mdea5FlxJoYDjw5zUsN86sy+8
QF7R6vAatSFZWeJ/vw/eTedNYLGd7YvTAktVxfmmZ4yPZ1PVFcGWW4xrImAw
kD4+pxexzrhFMiNmAcliL32v07F/8cqZYn+5KurRJQO5cw+Ru+AXcsDWKqQL
glQIWrDLOcva+N+iLpB5aPnHL/RIsD6SGTT0yaKSaeVOLa3R3DgMZLU/zeHq
PQAYxlKnMu7Yz3jqCSdSyLe6Oq+4xlObz3o5be7qhX3Kpvqng48v9ede3K1G
3D1wXqQMn1tGZw0sDm0tEwU1TLsKlUdFkZh5dJkSZ1fx1tjWAN1M32RRAPOY
Cfum2iNtLzLYhhpstI5mQxH2sJYdcuD8s6aSzZeAk9WWVShzTyv7BNUWBmm8
mbVOv5oN65qUGMAhGc/AtqrfRFUdau44/ctKixlaVsLyjUX9lAsAjgdMEqgr
nFnMef3BfvjEw5CcA25MWjGjPiP633uD9SVRQKAxjLpOZ93YcVxczjP/Igwb
j4ZY4Sxygkzl55oQ5MDxHmNMN9Ml/J2O0S3Uk0rKo+27L9X/yn7ZPeZeisBL
zWpY0X1e5ELBll0ci0yJ3GM1/IOQxic9dK2+Bv/irXYJljarOAofcbRXS286
7lckQRRgw/QSzu1Q2Rx3iyYvqbZEpRoU+u9DeOvJ6rGxKyTZFSpkZDchPUhj
r9+hDx2ZNDMZClibasMSdUL5r6nu13BX75K234kH2QSkyDVkmpvENe23sqwn
T5cyPPSb15GJjsfM7IrW7M960BA8gb3JzbVJvusutPkbDa0dYJ7I0A9O5mtG
rmsTqghenmERaBTaDGGcCrRv2qObTLvBXYFLHeH4fSxzNBBTSQ7cwuncizbB
pwgr/Iogk7h0ypVLgiyBpH1xp902iej4gGQ9e0nduykzhXtAGe1gzAmIIMJ5
mL1jmCFT4CR2S5z2l8S8MEWp5Xohx72oahcROKX+SLeXOA4eNkceXLQbNDLS
NXBJbD4KlRls4lBhVyjcMewXJU7mkEikyBtHlhk6Gy0yBcFzNdi2Jm52YsjM
eDasV3xlPYaMuL0MHLyf0TVMed5Xvo8unRXUxTM2p/mU5ApoLN5qGdXctSyz
9ayHNcDnVSO51BHyHe5I7bI3AGDAzku1E/kEVP+WwsFGK0fpY0kvXSnM+bsp
SzO30BQV+nMFAayMDc4uurGZJYM78UKXTZuwK2Jl9xn61GA1KesPv6TWc/mi
BGDH8NvVPzSB0qdMP+LyB6phgeWd74BkyrwwQz41fF9wGXjD+DVxDcVLRvDE
K1NfXRB9Deo8NmjYKgZWwtNYtAkCYG5HLt6mn8BzsnSkSqXgVcOFR2Obgk0s
VJeSsaO2fr/EmOcD2BNcrVj+jAH4LVLEFvyXMDcGjgdeQXYqRJvjEwFOkJEk
PO+tCP45+Kl9gAXvo9zzQDpM7SWJmLzvThId7SbkA7P3OgHuRWX6yTie8RYV
OynIjsbcjrufsWSQn3iIjvlMIWl9Skb8Ssg8IlgiJiVFTxMEa8hARxOyyeH0
LogDMFDtkRDVchB2t0y865A5qk1E2D2AlEUazDfYlZeCTSlQvL+qdL+nM3+q
Od6HwETe+/aikDGt2qpoXnRL/STbFHH58hPXlLz2bTD8EG/PNWdgCoa38vSR
yQmHflY+U5YT/C1erpo6mCv3WuQsYBdka5uyrBkSoh+QlE+VDPbrJZm2FOWB
p1ffR2d9OZn+Gvj1R1V65PAkVfDRqwiG1JOrkkd/8m3Li58D0P7vgqP1g1X6
T2/Uv/nlKtOHG2+iSaKZRpHGeZE/ZhxDmp4OROxzXdjwDJCiy1c4uaMVNpxO
mirvXS2HKHWSGGbXiOILg70yDsA9ervGfYPjWljrdFE8QhtJhHuJeJ6GxWdO
L5Aiu+6Zg8TdZCEwsjM8aG2kFirQ4lR7Z6B+gAf9TcDl7mGEhOA+XhCUoy+K
RHWbbkD8BXo15dCYmZLItmdJc+4i1Pnqz1G7WpVd4xgtiQJxw0w7IsQ14XxU
MAnmIRbcRdUUpiPLP0hpe/bV9Iu1YgHr1h/HKOADTMenHBNomsZ6QAlK8eCu
yuLDTS6+/+hPkVUJXumFf/lRMuLjyairPkcLwvpLEiFIqmlSLgtW2sJFg6Z0
AcLNiqgE6cFFD+syjTuLnYNXjG65kJXvcjA7lSkOFNsSjhAL4zbUQmaBygvF
qtOVUvDSSU4MwHdc67ptjjKb6JDWmQuFnYQx+Rk/wluVSKy67U/jWvdGXL72
6lZxvHov9PvrJPoUQRyNxN7KKUejbhCKgoFZAOtCqaV0qTCAJQWSclhUcbYv
UP0STfVH0DI9ST9y2IBPuwUxiPQadfZfKPfycpHiXczzOyvSCP1HubEeuo91
z23zAWk2YUcpLJEJwyZcRcEbcyJVYsTjfksOLIxr0WcKDOKs/oNVXbdAJn6a
0lmH7DdMPcOUlec1KGOzOl+IRdjNPXMDskA7CSe+nrZV5ISz++jvI7XP3x86
EerKXs5hA38zl2q0eKjAV/hRmuFK3GQITrv1lh+3eOatDOJQnX+OtbH1q7sT
19ylile3o9USiJtxBlahFVJxVELmx1q5V4xwbY/AN0AV4sk62BGAPfhhOgUw
PNlMjuPRBIlB2bjRIjfEJU/RVoM1o/1lswJ1G/hHeJM0NCHLbo6y1jdr5LFw
2KRYF7oPufhK9XsUOG01QBfZmzUz/xsMXhBOuKMYB0fb7mC/ElU1+Ib2AHT1
+brS+7asJyou70Q5GNnGV4sqeDbniRbFVMSMtTg72l/GRKfp9ncLmVE4TcNS
pdzMHPLpFvM7FPuHmP/XXuPqeDj9eR10GhX4b0sb+9vk/2NoKO1t1ZUGCR/S
ZtUoOBuhUiEFaVGKvPUswKXogL0cuNBrIZzyB8MBqLW0cGaK9fa8mmbaQgIt
ecBH0dZPiJbFFEshtstqjq9D8Sxc0FEr6g14TxCPQH5HMF3lQZX5oRGGZyk7
syBZhyuS6Hx8fyn2fyweWCkbZAUC/EHzQ43BYheJhsj2IhHA7PWBSHZftYTK
NoSSO2sGC6cTUl5DM6slmqXNo+PL+hV6uYReZk1HgwxbF/iKpxYEz12zbZX1
wcNiL3fRlbPBt8fo2neFiTlBH7GISByw/64ySn+Ee8iReyirvHGmmzZ+qnDb
fhETwoV/Dj86UWMkix5tOboZmB+z+TcDFQC/JkpTM5Bal8nmwQ7d7G5CmyUz
MzmAmjfZY0g2Q9w+b9pZcPXY52L1B6pRplARqMJKA748QPGxmSL7GL8OKA5o
FSK9l98AT58PwQtKF5VIQge9hzF/+mtTqjDpqFM1CkmQmM1qe4a0pGAmh1Hh
XUwFjtFCVmHtNW+DpMfG+uKRSBBq8EKJ0SgTgqZc3h+DC2c2V/ngIHFIu5Gk
mz4PS5RJDcq0c65TqE/9bvTcqcLUzZ18hy10t+I89SGT9PgJHwojcxJfiXiE
bn6gueUNUPNlbyOyKM0xopt8pjKr6MgYqvB6/CVQxq7R5WrojLpvYdxzeM+N
6lXdcn6dVWVcbCGOgKtJ3vPre8JcFiv+W1eqiTXxM9XZKJ/Umgix3pGuvPzs
KyRl8YajO6MsAqFF9nRn7L8xRv5g1bJ1p68pclXIdm/sA707/nLrgjVuj5lP
x4Iu1K7VpFZmxsZO6xQqSGrK1Du/20rH52jCEWH6GewzHzZKlAjxBE43P38I
1MDtL/5K7LreVo5v+fmzw9N23lBseK2/TL/5+muZi/B7awwBinpgexl6M46d
L/JLogk2EDsiFFV87VU9v3RNw9qsOs/z68yOoNKRNolsWiYj+nFaKx2BHwEO
um2E2RciVOQ/CThEm1AyVUFWyU0/+R2nR3MApwFNIBQa9RYGMJ5i7LmGoMB7
Rn6WLfJHAjcpJ2Z4vDEhPqtmbX7gNW9sMM4lV3HVI+WuxS982ha6LFgjNR6+
rzmQN65MY+Bw1fKVy5D5jUVOYdEekAVGxc2gsDRrKiumCrNijmMGuGIBWW3R
fsSic00x6LSd/YogCj+PDdWwiHuUHJeTHTRn/t5I8p4cEFsEfaJ8BdoFPBDY
QcMZYICzv8WFEbtrNvZUi5AUmTNw7tJwoz9P7ecVBMcdRENz8p+e4tnYkovb
Roe7TfSMxDMKI1ehRVhY04CFbxYhSqoTjIzQ+MYt/t44FjfhDebO4SE6E5mg
1N/IKnbnIIcLYOpw7FVPAY6fshdU9ZuDf2ElK6utsJnP13OU0+yzeNGB3PRJ
YOOv/BEqFld7ayYD1nEeQTNxlwoCMp9g++lFAOY3YODLn9GhoF1wCpFu4Lcw
xV3e3UsQcbvB//02rTsXtCWTLxnyn+2k31DIMDYnPQpPWFkqddoJmRXDM06D
27skrRhkZBVwODuiUk15xWLiExia0zjvJBjsZw2wglXl3S2mtztuX+evMLSW
wFwFxiD/85pURRGdeuLQACH0Ojz4c4Vs+GQPPlVoW1jXWTRnuXSauq6R/XNJ
ClwAFfWsmBRy/EMAT9y0kYDR7YQL0ASo6M6DVdloKQFDGrCHjpMwnj1YCJCp
LzfF+IccfL+/Xo7FDVuqMH1ytn/3oGYvZ1YDXTaCloG48K1V9z43Yj+eZfKJ
i8XdUrPN5PTBUBNERZiTDgLKUuTyGikr8scIV2SuwHuyOBTVgQvSXwKADzQk
KNl3pDbWciPFmge0dOJlUVLHw7enp8jY3gOV0oT3ju0MnRyUPnmqgmLJiAhj
Zlr8KRymEuMKnw3SWWM2MikxuyybVgMRwRKX72raoHSImPP7C0iJaFCoO6LN
ShbCtZdOyXfrBCLHPN1cmZ1vyWzk8Djo4r/Ri62+q7qoFTBALS+CWq1MCG9W
WeLDPeo1wImgPy/lAREmhbDSQ6d0dqyRRyauS+tPGaWfb515LSdarhPDsqMb
jFB867UmZhMHZ9Da811QTLZUv7KQ8fwZfATs6boUkwZnXkNSpKM8qzXfsDXz
W9aVGirWaP6UwUahmZOMVvP7GIcbpf0U/eIcb8UwLCKGcUKI/sO69AfyXvbY
h/JmsEWa/GHVyNerif2f8mza8qcTDb0WpYnwuIcX64xf2549YrFXSZbo/PXZ
RzmUKDQLaCUKyIz7Wys/vQfflKkZgWfpbQqJCq3sz0+d+SJxeHaGzemYj0eh
esVAQxX0lwYcF5jUVEhLTtv7FK2wQcTDW0kZMpLHPGhm/HE0oZCuboOVOrki
7Yo+Icc464IGIk2lFN1aL6Ye28ps38R49ous+4g0I1ObEqpfrUFS8hT7cM4n
UN2znOyKHY34Rg2QrC+DMJGHK2Kij/OAvsSg72uJVM50+liA5/F50ag5kLaK
YFfMsgxRL/goHIW62WJFmiFzWJ+kPzwQirzrgyJaKeOn/SJHtpA4YiN1Z0dC
wkVUezfcfxXEZICkDe4LGK6+QEMwUuJ7VU18209uUc545lRv7l/JNy6sOWKt
mx0IMkl8BN5zuo4hf4xPzzM0wc6A0U6Dbq83RsiheKPvzQP9gJvRLfJnVlig
qDerXBugH3SbCkMdPyU6FsnOb0Ooi1LYU6S5t2/PwxsgSnGjXKrhNJTzQKrV
iexCXwzJHSOTtiEdoU9K/cvT2Nr1oMWPjNdmCeaxrQUU0CFXzsSB+lhzD9er
9btLKag8hTJ0bUnpZONOrw6QpZMa/+RSe5uGhG536aAL1o0OT6H/2ASzOdFD
hgTyitLBHagQ5TwMquNML2MZRNFocRyuvdEXpSeI0H73oz63EyrW6tqy7Sws
Ui/w2EycOt+0nMyRbX33GQn2KcEXU4LrhfL0DXBQDdaB2A8vmqjWGjXnE87I
gDsCWW4bwoVUut/R0tvmazESblWKufuy96ZNuu85zx/WBTiAXJ/Ey+HI3Wf9
x7wTYGSGooFof20wNqT8QG5FEDzEHDOhRibjTzG6wzPU9wtI2MBR2dT/7kfD
KW82UY+4n+Nq6LRcfNdJrwT3t2r/MLfFfMxPzrvCwotEQK1QX8MAQy2tih4p
RTfCxB8xKP/QzIvmPUV6IhjM9aHhqm2PhO8KlsthEa9gPo+6SYjJiOBuJGJg
4B0YXQWvfHlVACSy+En7EXHeU/61BoYtc9CYgu/7671VJalXxi/M6K2FJhKW
gVjluSOSgaNb1fwAAGdTGM8+NtyRDKvglIus20Y2Xl9JsLHYeqHdfxqP7QDR
V6xu8kCflmFFc0z/oeNKt0xoqQtFN7O74mAlalLbNIg6VHio/GdmIunbjkHP
4g1gWEzgzTdge7NcIxkYszD9Py9A98yjkBGCnhQ9jcV3KhqRqB2d/E5lduHL
ftHWYLnryKjRLykynBDpLvZD0UfDPJMaHtDiCmcRHir4Y55TxaSKYd61LxYS
ABcnBbB5g+d/C5Ud4OY+1SRVfoIPl3WxHaN+nqeRm0KKNnN1fo48sBlS5vm8
Ia/BdVLFtrJwAtNKhZhb0AtxqoezKspqoivFVPl0J0+EepfvbFftFh8r6hgX
1oIpv7RkkCwBoJKgGwbDIhDn6DR5Nd8jOKzeSYo+mKjWXVywsXCmDT8mWnwa
UyolqrdkUCkWd+8Fq9PtIdzEvdlj1YHvdNnZtaBzol6fWFcKBQ4LmTqNJUUH
vI+iu8TCvyzF4IhgJEPRtGYIZrrjlI0JWB99YCo23fmqE2H/F6fdG1K0H+1w
BycIDDLbwLGCOxucskZDLthcKXvWkNYs1oChzpu/iT40pRmiS/4iEy4rpkx5
3xDreCk2So/xjpmsVD/8D9oHrcq/9T6DC9kkpRPjjvp7ElYKYHNdaS9wPNym
FrDTdu7W7/FoE8IqTA+AiMWg7jR++gPf2wIrqFHlc+M5eXbgQnzSHGvufcUb
I1n9yXfO7+FxkGQUphPVglU6Xep5feMXAeiio/2cBJhT7wQU/JuRROCPnDFw
3K0kjHECUyQKm3bJZ1dPa6oKg6ZiwkzmVvaL2OhKBYoPXXh7kjlCuvdVGo7C
QHS8UWEYWW2XQGi2zOqyakpmzImSOzyslynfAGr95Gi3qDTdg5Qjvy/X73HF
wEIpkCVcNs0mOMNb8e5u3k3YO2Dc3az9+xzfPWuzpdGVQceeGwForyB791xg
ia4cC0a+kO2r6kKewTrgYhvYEwm/sYi0XjaZODV3cuaJqfC6wHnCkhg05gwy
3NRbTFtOzJ4uHjBp62fO76J3Qk16Y3b8i2YVnsQLrJ+BU1jgPWWZmdSf2Crl
kGj6E726ipMmWamBKESp7zaG/RUUbytnVTMSnkMPubwbsZZMzIt6krdjQpEm
BU+/iBr1j9XIdFgYhxaQBPCrIjJ3Hm+bQ1ydXSNLpg4LJcWZ9GO+JlggYsvN
cqNr7m8UTNXJbVqPoAyD98pq37gZRpIH0l2/Nvw5NodROQe81+fymDss5DUi
9MvGmctsxr0qT1+BNs2Sl+NBBk/SCapegL2A8wT2XeSBGaJUgsgO6H7SuJ5b
gc8uz0+9NLJyPyXtqYXrN2FlO3kunTIQGxm58bvsW6fVvaYX4q3pEWurwQqz
O6N/iUBjlr4H0jxGu9gAPED9VQ++D1LinYUhEkHFH7IogBzjnFIQlMXXiFNE
m/ztS2NRV5/jxeVSKzl4azB3ByqflZFMclBUI1X2OLhbbWGHniVCAWmCSLLe
N7Z9QX5Jmzlmd5b2UAFSUIh83ogDkwz7SN2DVC6uOoZo5yzI45GVOyloIJ0Z
eVK6pSWJwUlSoXbr9GtNaH2ou4C3WRPH3NWcs7G5kL9SqmcXu9WDTLqQa6Zk
LEZR4BGt4YdtDEyCWTFuf+FASlBxdiO98mgr/HEHVER1t+a9tQR7/QcKHnJX
Onul9PebW3gbgMnyaQAnCz3gWijBEeakL2RnBF+Yex6Bg4vCBkr/B0zmoVCK
+OCaFK5R7U+5E2o5JxFlmBlOq5nrVtmLHX5OzxZhY4nAEiqdRURaI2Lxwa/Q
ev/Lr6RjTiHPxkLRbTf2OU1E+KgV9WYvI4dUzgMj73V8I6pGRkeFGOhGR8cg
OjQ6+IEnOf2fyfE/dMzGCr20OJGF4OhgcTql97US4E31iDNCfH/dNE2K9k2H
aPwVjSzam484xKQ7leEXtVqRNT/2vqGg2FQl8ndkxHErAHFK2d2VkTWV2nbu
nBcaxM6KuV6I1JZET/GSG8FpQWGBv+WhAckmv+TAZFHpeGHRl0p3lJXVdzjU
s4vN3cTusotC1BiLz1htqom5B5Iwv6LwKxBf3GZP0wesWPDrEGXcv0U3ZI4l
jY22RGWVQYuH04bolt1+cg15YzDMFTQqvyHtSf29cqbgkB8N4mQLMJivapfD
ggdDsjCFobM5NrOW8TcPIusDbFKMcjCf+jFWw169awtjZB8G9/saHNU//SEi
We8ZhQ/DyrLIpVcjXJynqmTlHKXN7LSjamXjMjkP6HGJolg0qszDLKqIDSEk
7mxb4amFC+1l5I99H6LOIjrFg59iR+O6dwgDnhWvkiMOyWcY5ST3pTPjum7y
xLRsaXtjV0ZMhqskpgLDw6OYNCCthVAg88GWBTrWYgY9M3BQh6Ss4b00ZELk
43cMSjPILLyTXKYBsL2CGr4hkP3nJXz/b0DwdSLFvuCSq7RL+qTYyQaSL+o1
3eDJRnB0YtBciVtCEzd4cubfqivgeZGDxdWte6QjthRY91k/N9zpWC3Hw3W7
QXjcR2YmpUU8SVREhI0yWmNF46wcQ43fwL9oNAnSqKBErOWSwtAoqhW0735X
23+fJYOIhv4R9P2dikG7ADYb0Ym2F4+gtVtYaxMNFTPjLMdSVRpprD0pd1hI
PGfN7Tl5mQehgJcGXvn0sjs7126+3c3XmT6NpTFU0s5ZN74oTKYd6TYhW3np
ibqSDv2YdC0WbkMFCrscAr56wqX5Lnqp2z/laVaB/aXRf44/HrWFADbOFCZS
grpeFBdt8xhu4NPH/FCOJLZjQZAIcwGVUdjFFcKipfaI8FjoZQ2L6tp3LUlp
OwZr7oTqcslcLqN0Bkbwe9Csrom5T9sAcbGi+9eRshf2t+N2PMbHKEuERJhd
G9II6tBqfcs8Lbu425RMegfrmo2BK09ZknFnpik8FRgGDJMtAKyZ6sZkemVR
5Fo5HebMtH/Kl4j7hfguIpC3/v8tcS8hH/SXu7DUZ9yMQcxiVqPA6jaH3uHe
tSzElLjpSCOtf38e5iLlaE92vFpi4rf9X7KvKyqYnxl+sApz8Ouc5wfhEajt
z16ahV5kj+GVSRH3KiV0L31zJ+PCzS0vtFVhCCF3npEO/FSsRw2aoBlGAQ9p
uFk4saLmtZO8WUI2hkd+U4iowm4Kc41pGEfMtG0LyVcS7gIcJ1vvCYRN6r1H
HyKmUvNOGDKyw8i9oxvzJLDXLztf4/7dDgy37ZYv/euX7og+DmHMiTb/aRZ2
SIXJCD8vQm6t6HKvQsplsC2zsxH5c95mIWDyZlZewx1l7WBxTz6lq8xMrWZS
DTJCcGkwwQ8wD4C8Ox5LoXSvAh4o3twiK1vnMleo4+EBs/+u0pWp5RGOGhGg
cwYUPdaHV40EJPEfhj951zuTTojNFweO2ybYvRZ8zIuu7MsOsKZWiwfN7XCK
+Kp97CJgP9+Kxl7D6bwTwgHXi2voVCBAchpVQxHzQB55XFQLTVSPrDxYVFpa
p4NiJw+4mRfxFztfweA19UkKZuFXTFdmPtgeT+QLMywU2TpTfLllHFf7+vHt
ntirYWUwNLHjZKFI9oWbiOufrUt6jI+TXIPR0/XYlA9kl2nRxXK3z1QxiKYx
luKGp4pEt/6AyjvtNDHkdmlSLo37Fim00Hp3cw9Xo3FpxphWuWC2SwMNIUhQ
VXgDW+KFhUoSWkVaEh8zubyXJOzj8Bu+bge7Gzr7AQ0yiEeQwMHpYLc1u9fa
Cbcc9A1/k/o/X0FkFhl0zd1e/9eq7GQ3kyqiSRrfz8dmHcHZkie4spPtqXvZ
13p7eaOWePg2s2+99w5UQ8ATitWuKribjekN305EoelPysIUMTsYaIHabXHN
4Q1zJMmhV+xuHwaKQzRSB/xUnkoE4+GLWpmlSCuEcJgV9i0UTRHb0jZ4elkx
xPtJbbaA/BFBiRMSvsD+ETBNfZtB3RccoRpM+MRSu3r7UPWxNl/h0tCFDpH3
exPzVp1HogVtZ+sMjVGYixnqUulG4rpR7e5VZWhQSxP15t+H1caAH1xM6a9j
qYlp3dAL34PWvbcUAlYBiNXlRfHslX7y5DkhhMR0l5mblhjAPOixeJ6DmTVD
S7t63IHgEaTQTimcqFrp/BRRo39dIXaxwxcRGORjj0KpNCcns1TyKyjqQAFn
GX+6mihRmZ9fWLonguwZrGeFYyBObQInLgasoB+5wxJfjpWZlXXk4nAzHpyV
1bgkcTKq02+/3nKvcnYHevNyrcD5T8XTfdYYABhhSOqgVV3591FIIyl46y1I
BjqLRv4xxzl1/AUv6sBBtcZusZqiXVPOQLtO7K9kYXQfjsO0z3Ba0cLafkKT
kfZ6UqvmC/gfawMNnXXNdQgxL3Fg+26o43ZxLliC7gV0nCr8rL0By91GPFuN
Cx2O9XO5ZrSw80PMUYes1GGbqkdMBRHs+4il0DBn31cYiS9u8TlgKZ+KdARq
+5uAOGbwBn+pivtUBq7dJe1P13Fv0B8fw7CRd2/CvAAj8kAak/S0CT+f7reN
GEBdeleaybdh838XI4WupnAq59ug4utxF4FZecPOKCkQv6ladCpgeu5sU0Ju
QmFvqtlntcY/+o6Pk8CwzNa4yI2PLP2Bp0JKeoBQYDWyn9OMT/gYJfZoaG2V
1lov/I6lfEhbJmWUgKcafC4ThRXzLxlWVLY7BgwVSc7ZLhXwOeYQW5Yo9O9m
bQ1S8NP2tGETONUeyv1cisyxUe2mm5YNI7Bx1UM7Auhb+lIMxF6im7HvGNTz
3v6vcrT6MNxWtl+RkFJ8oMU7CT8a0neVPkRbZYFdmnPx2h5cnzHfExgGtmiQ
p+ib7pUrtEYTzpPEkvYA1AK3D5pYd2CuXNdoW6M9tKQUxzYd6AJqXgewlCiX
lBLwvXxebs7bx6L84R5pNBOCMwq2NInL8/J5UiEgvhdfEsJQnJIGolXtoQGR
sHCDaYntIbGv42qsBUcTNiiRXhRhw2WTO+dgUPa7RlAIKznq8C/iLJgcQV8p
natuU+6uhwGjn8jSymSlcsePjGuq13XRBFIIBsSFbISuv1c/+IWtn3itMCCt
kNBhIUv3a/8RskgNmcFipzRM28RdLaGcenRNvxa2AYLVVzIouNACSq/dV1wW
D9uUG9H0IVLRe+sF7AyZnwFU6XG1xi0evRpMK3rYJ5xfV6UZSaAxAAUE1erz
YTdVEPNu+0l9rz6JhWJAwIOXNQeumr4H7E7yMPbHxS/VWRjLRxcUh2J95Imz
VGGpT837gKqtju8TJIIQGmSitFd22ZjjWx2GaPJXR5xg9jiRyIBje4h2XsP1
tb3x5JmXbB/hiM1RHDk32RL8OQDg9oRk3H4adHrahjTrF3MOi+EnA+ku3Khg
q94a7DihZ8YwCIVGLo29iPuTU/QUYOMGIz4+7+Iikx00BSiC8DTi6HGo0D0g
OMCRzcRcm/iau1gGvgPDwuJyVWtuyZn556rrsT2oUmsLLAle7ApJ/KV7shYP
Q/BIqhCnDIqFpY2a8E4UQAG+hnIq7FtGSOmZCGnnisXk9KPUd9LVfpJF9PIy
8HcHPCkwSrqwe1kN3cV+2e3XsmW9+iGyPsRRInEoh61QD7du6I8SWjTJgqRE
d/VzJp0wVWSTyd69w8eav2u2ce2GHrIA0O1oCASlxZ60Tl365A+NMcdHikm/
+B1AzOnR87d6qjI9uoroNIwfxSxtW+N03B30nsfMfzfq5Cs2ipgnz+NetSYs
+dqBysgbidr9wLZ2tnWCn50gp0k1a2bnFz3VIVs3GAIc+iaYb5yrBQEE9Euo
T7HH1YmSzifZkDpRsQzdZNaw5gAfXI4mZfIETNP3TYDCuFYY12g495dIaPle
QIo4lKMPTEUw0tzEOLawLZ22raEqLZtFpt09ph/8Lkdz0gqZph2ctFt8rJkb
7l/aON9IDbh1AHftNwl76CZn8m5XIil2bfin1WnCxVDicGYfwj8UFIdRXPkv
W6F578FXinr7zbzR9Zs64PY7ToezXhCo3/W+Y7ybrzFRuwZMwbwc7PySuP0T
jPhE1RD579zNjYfH9VSGkkDLiw+UbijHZSKWdZEvHZQ1K/gUIJs2tAigqYYB
XCKtszbvoJatTD6HjWzYzQXGZ7Bxtb6/oB7BP6Cnn4hcvebgH1JH3Z7ak+qp
U/I1n0OyFgJMPwGNVg1TlF73xyqS9+0v7L7K2JzqVK6p9g0ZwGVHot+D9eIG
kzbh44KKov2/JCCTWiI0ze78tZhxX969IyNLuwpKJ97AEpq8zuIRTPHwm/Xi
DKfrZOyda5CvUTnsjjwhZDCLiaEUTFBd7Wre3YdoJHK/f1U1x36xiRPUa5kI
4obhHCPq0SWGpJZ8oQrhoqcCYR6bEEr7O/L+3Xt7JICtkcbUrjELh3PqvM26
Smm53O5qMi7AQf70LbpqJP+yfgvf0U+RDNyE7ZfOfgNEFxDwKTyhWPRHkZij
Z/Mc0M0NWjTbJGtBcf1PDWJE9Hk24LeX1kqWpgBMgz5uBMaYUi+Sara6r+7H
oJ7Lp5qAtI7P7ESLqx/j9ZEeV/HPi6T/QuCOS1pK7VcTebDtRwYiy52p29SF
zNuFWjQbo+RWm9O+guuzyP5TM5bmhME2hHAsGnjHs+18jyn5lJ3b+T/N+mec
cHy4mXQ+eINVAjN5XVZoIfBhoFFbjM4xBg5VTNUIhizPp9c2YWk8r1INg4ZE
6FmehRv4csTRZLowM8blsszzaA05vh8LZ8KICExwNYPepYlS7l9ZLpuuG4el
1Nkh6/gfNmoa7u1cOSG1BhYBVEFhai+npWq+G+QnKyDC25QohG9x8eqUGHxx
v9w5fgmyqYr6tYcAE+UyE3w8Pc3t3q/Ohr8uohY3Z9ovduvZzSQAPHtVnhf0
tny6uOlN19UvNgwzE9n+stV3xI2YNg6p4OpjpOrWiLqw/1FpTsGs0IrEBaHf
e2Xtlqc4PeZpWZKuCcdQyfgSrS7wQGbqNYDNH88PXWS2+tbnodv/LaMbOlT9
Px51Zd5onS/lunGueC3hiw+haAYLZNBL7BAUT4d4aFKPXyjf7AaYcRXk9FbV
oeXdQQfemSSguyFMOJtSAYz199xyjmUEjoyXjETvFV+ha1tChSowSslP9L1h
LTI06Akgz+YeaVIHT0M+8yZadZKk/H+cO5tdylaZEcRk8e+xlDfwM7v5/Faw
508A+Mwwl1nbffAL4afDh+ySzO8ZiVhDH9/Fs+XyoQ8Bfs6ET5ODVcQ2ex5u
S4ap0v00STAEluqykAFCz0P0T9OeRXqzLkKqUSyjpqWgsTRW5C/Od5TJYIL+
YIoVZ/QrrRWBmbj73wddT1WT9mj2XMIzRQnML7xBUISF4C+0N+c5b+JfpJY+
yczbZ05PnUEmIAAKlNa4abin5tkUketw35S0pZAK2KXKxcMYgXGe6J+inmvz
T2oIIj8AGyZzfMuWErhxVxJwj+OgVlUhFDy85PUG4jAWv7AngwjvJbNdss6Z
ECHO7HuO7ifmMZjT1gREDpvusfar4gDoAt+fdEtJE5uGXZMAYlgNoii+bzQW
0fulETMt4744zSQxBCFgB4KXYlzJ/GTbWCJSmWGAZzNQ6GRC2Rlo7cUbSd2U
0in6X7awWJ43ig9KpsBI6xnAJH+HbHEVXR2zzv3bc+ZIlbvZTibIyEUscgVF
IOl1/W40s9xu90t96/mGVrUlUhADOd7ant3evXNAiV179bj/pQOTWmAI9T9U
MKh4yIsa1NWgOC+bc3QUBqaSL+Tl9E9hSKG0LmkZnb5uBsmMt4Wn9LMiD58r
YFO2O076xMhVqlrx1Vu2ASKtW59kNc8IS6nEYDAClg8lfTWDNtxYLRjg5vwY
vrG8YyOYzrbn/pD4jhJwYaj7YhtVEKYjIKC4pwwYr0dtJblqowhdi78xHhX0
P6QfV2+QgeNi4qfDdSk96Ewa3o+XRpuULyFviwTZmaJ8X/wlriTPoPaWT8Hr
OYHBUm+w4OL3Yk09qef4pOTk+1w1w2lYQQMviFCiPYe//u3mAivPtPsurSPr
A1Sn9N6Wt3PhJb0Y2YwdvZrSR7glxUis/cXMEnDX+8qv9rSitc3QMD+blJx1
ME4n9nqOHipMDWUZGyLl04sT5VT57lKBMKKL7gvXTe6QWexKZc/Qtcek4e/x
RgZYkMP5I0IjCFhbBh+1Tkk/1wFSAS+KAO75skxY6qHimZxZuwP2bpsuELd8
RcFs5seZ6SokZ0pq6YKE+XHJwPzYoj1kmME2XU6XPL4J4d0jqGyU6W4tgqlX
HoEkGyul6nQekOsTkPsyv+6yOia25zt/zR46UfW+jx1yCaGhk7FOZFC49pD9
Sc7hamy3hh1mKdvwsExRvcXexaz2ZGznOOAx3Crr1QFYIsGtVshahvfr7p0g
2IzI9BVEiH94vWYCccw//h4/T44JlIUQRCVPCq+wGqjn64ZwFugmLbcla+A8
EEcSy8ymGPTf9HtUFAuvhBmFgIHtjzO+fbYYfCDTXobTXfVokkcG/CXZE54X
3M1SlSYCmEE9eIZov8eJ2DILppD0GLzGEgSYYd0xWhSFnA8bkKs/ohiLDicY
Bh2UhWmEfmDNqATAFTABlhSCmYDMf+aTgn+SAoCHc9N+iKWMCQBwIsbyJ1UZ
x5D0xndp4J/R66AX/BcignyezNHJkdMcie4wjpIJJjxdiucMMbcCpLF/Fkfm
q+HsEIIdDogOA3+s21AKICjXEfpB1OEx0fLe/jHaZwxBexS9iyXX6txUFOOd
XKL/eohvOQPLG1kZw/brMNke6VgMgthrE/4TBgUn0mWap9IBINVrl8iE6mLC
Da7RL2ZT48enLeXBdmFnrpgplnnN0k/Js3yhKKLmQL9SpNxuJ7XQoVHbq0rv
U8L1OEZOFknSFg/rs4ipGaz/NIAuV/Z1/K8HY28WFU0jr+ORnvC8Qq14ckDB
bGlsSTcBTtiEYzjWv6+qLIItJ+s8OO6Z7aL6phlKI0CxqT0S2EfIczm/up+a
YAEOEuDCVBjlISh+nFNv5H/1a4Ra0PTYf5ZK4VKG0BF9k5vKnCR+/scbsrow
inDQbsxGrfIwBU7mH7ZtrWfyDq9vtdppQtzfWtrvbHck+f9NkbqgSRHPrXNi
QWTsyZN+iGLqncZwJRSHpFx0KhoJmRO62lUVZ9M/NzCoNRh/llZUhZxdeC1c
Lv4PL1fK2p6WDfiMqn64xdYe79+zZ69eZvBsTs/rCGRBGQWwUzSjMk7SPfFJ
h5j3euqdDTADAugSeNHTyLHufBXWK2Td08UH8E2JvFlO/be5ecVxcObdWTfN
zVhjTfd8Z34RaTpX3TKNh3ASEoEgEz8PVhebTYO0ujPFpUfq3MfA5R4AvH9p
exnL+r9hfURIdwdXGDtTriRR4VEioqQnHfMQwLdbvvFk7unIqa9Jc0leHZ8v
hw8DA1AJq6t25kehG2t4VSNfyxgYbU/2Ck8JKDm0RBVLPXuqlmgknkkSbEwl
bVtxcQQqQJHX9qeevbeJgIIuu0CEoLFi4yFYWUblXMW3HU5wZNe9Rgrf8b+8
wZHJGrOipHO9M6u1imhNrv0boxCJeEGoGVZNm4cqNjxZ/EuX8cnm0icebAb9
zE2+Pq6+VDYw22YoL8VduovCHTat7pxo7D4TBsfabjyF0ZdqhrEHbYsDoy4e
udJAP9q71uRaqgzxKprrepOkHttNlvBb59ghzw5lTcb2HG+r9HRdVtJm4mIW
+Kia1e2CG68VnsnzAWCNhx1jffJLTH+b4MKvcH4XbtP+v4s74lTF1Lalzrd1
Jfg9mq+d+GTsZDDRMXVx95bem35+5sF43NO0AKWHTrQ0GzCC67aei3Jh6zoB
gxEu4kYif7TnAxyoic1qVGoPS+sAwPQZ/Z9N4dql/EXjYF7tVlc0/JHeY5pk
Cnjz8Nt4p8tuo/JMn5iD79A8YKQqZt3ioRW0wcPgxaC314KJWWRyE0FeahNU
Ag2ExDY/gsxwGCT4+1Kulr8iYDmmDVYDNgH1RKa6wNDtGpc0R/yb9F+eYqZA
9+HBx2UFzVY1PvDrHwDMTEWCpoJk8FCs+wVjX/r9wHzY/a0m/8uaua2/gM5w
1pzM4MqstAaqhRfQHV47ZupOaLDZLNZwbfaZiUf/LImGY1X0ZLw2KKyi5sTR
iFFdU6olTrb7YApGvGPQf5yk6rdKtyFAgyXNuN6rEcYyoj5ZNUSU4DJiNmdL
APa5aqdazPnkTS9RT0dcmGsne0eYCmc+7TBw0ArDDcusrG30KwBE6tkU1wp3
0eagGrCeJMHk+uKwgrg1Beq3KSU8mQCCf/v3BZ1ZoRomUQe44v31NQHIEbRm
k7PN6K2bUbWpWQsC8vtuew68LvbC0OweGfKVv8pKXk8DmuM1V2o2ONJUR/Q7
pdTmX2mOySoQQP7GLqHKQmz9GZjdxpYweellZOKaNRqmbUQgFSQ0flN+cOfM
2QklxkAJd9A01CzMAmdCNbzn+6mCu3R6989VplqAwH65LWbIlUM4/+hNZ6qv
luoy09taPcp/BU7CQp76qC16z5XbMTU6P7TBaFkHtluK5BElP/46MtWejX0N
6ZGM+n5KXhzAw6AWXWm+OqqQ0bABWAw3Kj86OySQKhsis32TC3IjDeGq5Jxa
wQQt0TzSKN+Wz0oC7dGgeFMfz075c4sC6L87X7gtwnm1LRmVRS0hqHEqb0fs
CwoO3F4KnHXll+y6J8cRNj5mrBS/UsMr8D+qTXS5WysTEnB8y1Yo/ax18dIY
xcoQqiMvuMUEm4VVSpIErmuK42slGkVdKbrIVd+Le0rFHeqmMyQfbjjdMbWP
uFF1/Tcia/R1Y2IaIqKy1lsWdSOTC5LWTy/p1pugzIkA1sk318pxlgXTWsbe
Ps4eTRCQAK7A/VVPKBFpFMjDyRLKyTLTecyMig5vn4HNHkA+Svcym3eLzwpL
EGKmwkVnmHA8sgBIf6VsuTK+4skWpirPXEVKGtBPEhn4Hg0lNcg//hEuudW3
o2YyUFFrKLrayQjDDtB10mg6bypjYF15mml3coNq3UVcgjUEkCJD9ycyw7Nm
efcHxxEVNui0SYb0RgHcQ8jrN4/GSUZ1i4h8UTVUzpWGOnwIqdijNMkZVugR
IoRQ6py9lCtbN0mnJXlamDO6kRyx6JJ6f8GWgRYvwI7Myn5TTk91ewR5LoyQ
5i40VHIypHqKxqogys7NYgfDYssq0Fk+oQqrQ7eUy9BlqE1HFB9q14930nZ3
z0K5OmUJhMTeyU1EpT+7wri3/3N8aDW4cS1EdrUiDQpv1VQiDVTKpmoYPGDg
pQ4PrGY+4N3LsEFWCTujiF6MuWyllDndSQfQDvrxFlTxMKcPIezy7QCAJxgV
Ey+JT9WDCSENncqSOLz2r8azsaejz/7Xv39QhyfjTHwWrwJAc2hnuv/hDxf+
GoN3uoXRcaCGkiwpjTCmsxKDpWoi5j4hOpLhcgV8s82bfyHbaxSZqS6CGNF3
zE55I2oS5RoVMEO0S3EQUejC47DgMT2O/j7lEpH3ClBneEAC+LDfupj+6Zll
ucswPww3zo6EP2hSe+z4DnvWIB0jyse7ZXiV1mXT4dgsiiZ5Bj2OO6Ed2P5Z
32ejw2i2NYDPsNfke3h78soL74beG1W1JSCoNyH8gQ07lnovYLO8V4O7SN9Z
gXVrjKS/g+LFHSeNN8OHOSCyrv/+7YY+6uZJiu5oRf0CE7FKlZafiiu1PjUp
0aCoT+IbvFznan+8H6PuH3TlXJuMLYdqkPdi7EU8agU/eix31FaEchiDl+3U
VLDQl0LkKeohQtWpx1hAtPbwfOmyUrB9KuBrDGumtunux/nHynNTt9WOLRXp
VSlvK+m+PL1wgL4jWkgizJyxwqdNPdgIO/0H9oMRmCjtgPq1hoMHlGb9SMhC
2l/4QFWh0bZt0sfIF7COExhjBiLf+6eO9X0ZkJx6Iu59305Pous1kvd15LK5
AYGxh64LTJx5f7kT0wC2u/T4PROh80K9swAAM7D1sH0q2qRQhKcF4Nsk4N35
XEqzqEnHrqnxdU+hsbErIqoeM//AYFQLsfeEyBwrxhR8X+jUw02ReE6+WqC+
xGHIaqR+g/0w5XY02Pkcv29SPYgfoxmKNBSpxYFz1RdHGhLdJxjls3jCwpJV
coA6AEywRhnG/6G503bq1xk588a6qd7yeMTmQJ53Bjyeyl7Jj0ArNSpUkiGV
tXvZBOhkLb7dgpGVIJ/43Dn7fIWYs6zZ4MOAtp8+yZGG50vi51WlQCvTGtsg
IpUzxbdaA151qkLhMmI7xeBewE7zTx9jNQzWuVdh8LPnV0/Aw5nIfjxDun1f
IY6NyPGvvakS1jyrkoBg9gINp7Cqb9tP2Cgh20q3+MMX72zMFGOBvxVTf/L+
RqvUmmCwHDIigGTpZYITEYm1luvbCy4dbxu5q7gmfpNfU8s7JpEg+6oea9lj
yyDjY6pak7ocWbyKB1IoJ3o8DKHXnE2u9JRSVbH8ZkWc3O7c3lhiyoL5k22O
b7DSVJrlS31O6TCT7lQ819mV8yPpqzlanYJP1HdaXnEyVSNKChr+3naUTlbB
QtVGZPoitNFf9GCPOtHI9J/3BA22NMTGEmtSwQgmEv7uKPwDcdje8to0kmGH
cWflJrKpfuYBK3mxctQdxbPj90WA5gq4iDTHa7SrwG3KaI+VWuvMYqbHJH5P
42Mt74Oolm1pUHFLeTVe5apQ9ctnia/i/bw0Jp5hC4nATPyX1fbbkuOaWJfD
sEOrfxsfCrnM/BsJHay/XvkL0Yoo3yZIsQK8Vq3WLbeNXsyl1KHnWPcZTi6H
chrNU/Bk7JTdC1RTdA6GAr/5x5+dd/1M2qbc3+LyWn8h+GlR6PqVriZYuMBo
rKdyHxGp739umEZCLHeI0h7uGR+Ncs8FJUd9U0j7u4LIqXsvMXcNWa/bL4P4
z9aoNXN0ZZKvstJzA+cepR31WoNGntDlT7Sl4wDnoZNajt/haC0iYn7AV8TV
EbLvIxqyMrejlarAUZRNaP4ehbqnt0X6mq1+UpJaBAFRZVxEdzIzKHhycrb5
Iq/6dCGAazbaF6Flkyly1j1seGyCrgIpE6CHdG5Q0uxJDMh4dgPlDM7+VnIR
g+SqlFlGa4pXHN9ELmSbnPamkCrXG9dhUl2DMdObnZCYPfbY6ss8hY0diSxA
mFa5IZWRX2LYTsYbLXiKhhRxGrxCrn94hb/GywpT5QWadEnPVl9F8X3YkZuG
Mb8EZegpi404xKAY5ohbUeLq7h3xaU9jwfaD/VQLguEPYne0gELog6MvtE7I
+LWglPYS/m5hwOg72RNelnr7USPgcQhBFFv69Nlulb4A1npuqVvqF4CqzKCt
rqVkAW8hxOGOznvdPZJrDB9CsAm7fnefZQeMAVo7wIhnAYN7aUZrmdnjag3a
U3A31QzdE2rfUJq+yAfnyzOqePh7Tek4jtd9lEKEK1T8foNh0XbKo49F+jpV
Bfb0AC1QFSnaqjcS6lH9xiAsUfcwcnv+BBts5ZaYRFFv++VcTxUDfM0S4DIR
H6QIZb4YUVHOBLuIPvkQLFkzEy3a4vB51p21VjZ95nsKPo7No15c7trhK768
e4/3ge2mlF6VGfxKrQog8+px46OIQgceLY7N0IjaqMniJj13AXUABmnJYnvV
9DGTQ4LM9XAwYLHXFqRfQn1C5l8N4baQY2SZCvevQaJdxerLpangV5nzQAEp
l0SAtuyOvv0Akkja3z2J0m2ay+wOn32oOYD0U8XM8ZZJh8xOejF3++tIHP1E
X4sT4ia4Z54YpDQCYFquQUle4RckHQswZ7W5jSQE0fH+OCTd9KqCBXe7mVll
uV/r1cdBWtuuBjyfLOxL24wpPmWXuoxr7/Qgiybidk1C2B6plxXsVVtX4MsA
BPvdMU1fB4x+S/C2sN7lzsZksHXM+HQRz4IW0QUo35Msb9bxMAdR2Hw4IPAp
xsJR2DDO5yIJKGOskK7dD2Ql4Z1ncjJm5ZtmteyUJWjLt55EXv+PcJ4nd03h
fQUFcD8ifVwsHA7rW3B7MSwsP4r/lne1JlAwr4K9n7YD0oQG1qcKKOJG+Uqr
MQ2pXqcEDIQHjN63aTeL4dOVz4w3M+V1cJhFQe+zNTHUB4gSNoORGGOUhBF+
1haLSRI+iwcfMb3UY3nT2mHfco5kSkHyVUome05h3Fq/nDSZf90ec1Uy6Auk
frw0zPXW087g8k5rNMiB39p5HKVVowl90K1mV+sgaprnRSkaiFSywFeYg0aV
bb6jdMnDiKg8XV8junn7FpOemATjbrbr9YIjGgfkGzrRBs2GZ7hLS861X3Bv
XpsYeuJksW1tDzANfUaWuOCB3sJcSwVa41OpKUKofli1bPEqzwpD/8SLPgNX
Pc3kxQumKfXFvhe4Qyn6EqznIF/FZAcoFczqOvUkxWAK2unljomtZRYvCHSq
eWbGepZJGvv5g6OcVTJMwNLFcb1Ex6PML819+2gxiP/SRF9sSaW9Q7iBI/GJ
msbhCfR+UeUMURNm83gMVFKkPQMPiPSmYvE2GQllFoZo30aD0m2BIEO2G8af
rXGBnGYsXwZEiu+ryJUAuByiZOZRMPgPogNCBeQ+psS/k4X87QtnGV+QmgFr
ZvKidxaVemonxeIFiv6vI+mGHwjcsxrJeqUHLX5iNFAt407D3WxIPMaiGBrG
Mh+Tqg7lbTN2ZVucSRqJMyU9fPDvG/Q1zc9y5Ok4cysAelKofnRCpVkmcL1R
cQyDzJQRrw91UI7Qmso4FqZpQrN3teFQh7GzYoIsc82hVNfqhnRzNWz/qwin
XuvY9beO+1uGpKlIwAhQDu2HWisoipMrjio54ta7NEi0yw/lmbaf654C5zAs
cYjx6iIyTdwrPdTZaewgtaDieuMB4nhiYLj8YahFRwHI9Nz8ofKlLChcy4Q1
Nc/Hni2uvuiHTO1vu8qtFloicQQz+PiO/eKAiKFoEAfaL8MA/wjkNueDEFzf
O/pO+lq80v5KbVcmE1222IIq6HnA6YBtDmHy0XaJ9fYhERpzRr91BTF0Cpqj
D9vTeYYRW44X/oKhGVn7AKDLUYtfY8gm7nzIPR0s5XTUbQwxDA0MRp3uodCL
MptD6NY5mnzXKwwPD56Z+H5LfjvdfHrkODB740vQ4bCLVDxB09DgiK8cxGqe
PZ5VV/5v1gL3PyWKIFoM7uaOmqKQ02ZHi7s9/LOCt+aeEz4f65KSK1AnWTB5
y2QajUjV8wWIhMsE7kuZtS2ZeAAA8Lf0tBxMvYTxdaghq+GDy7YbuPgZfx4I
4UbC2ehcmLW4ehSDvDwTuRigmiPBMD0P57Yn+xQBy6MLR3ZEedI8nAlsIV4y
qYz9OtP2eSUphQjMm8esey78M8YOzxiopNTsY849a/CbX+WR+jLZS9QL4A8G
kQV82+J75NBF8vmkSKrfkJmpFmzvm7fghk5itbji7I7HaFluVg34BPNdNpvJ
5V9UAM0gPH//mbGhlrjRZ2jMviKIoLjJYQDfxRe4plaea4rAx2vvp+yKYGta
IYus3FwF3aR9Gm+Q68ygN2Nfsr4mHuxvZc6892sBybl6RtTxs2LiZGzlX40o
0KV3RnUhxPAZcXYL/QfRbkMOMHVSip4uy1/+2FWZ07xBjlEIk2x+XFsIT/rA
4sy0Os/67tNO+FSKAyV2yLzdjPvQ2kqwEG6MypTPxzlpZGH+LfOQVIZkj7eV
qr8z26eDEPdWsekxemB4LYNJd/xO8qbLKytX3RxLpe7gApmRJQtRy6fErrxw
puvRd6pkdtpoV3GyaB4CXmNb8MXgBKnbYktQHOfiPq+TkxQ+U3no42g0ttL9
wQ7+owM9C3Ozzir4g0Uowna3SZvf2/WbIvDe5EVSQ6qn8Rrf4PVkq1E0aEbp
JjPowqRLMeDw3up4oi7bKNwdYUfZ+Z925eKb4IU1OV3gxUmrt21Texu+lHly
nC7gxswt7MV+BnKhHn+5uA3csr1c+9dlaUiVZjkE12UsKU2mYW2fkm7BFPnX
iimWRthBPowB49n04y/xyE/uzAG0GLJnUDTrbPxH29KtSq0YXPATRhZWzK3n
p6+51b43r3gI2BrUfMbisnR6DGpVBfjKyNtYJWDJ8RTI4SGCABxn5tCK5hjB
kNesrxGxt9BNg1z8OkdpDA26yFTGDLYTeHghEXEdcpgP0nJwKrFddrryrstm
5915by58XszbOOHTPOjwpx/phJOqOVD79SL1E8GgIE/Og3muTAnls0wNn49y
gSaQxNCX1GyoJbQixQtd0KR45TFha9aIs/SoLPLNkAux7E5cemEV5H/77Zn3
Q/G4/BFoBWPcWttfIgWOsmM9oFydaB+OLqWHT6BHRky+/WFciH2LvDKpPshL
27OstvNBZ+Vha10t0mO93Tk4Ud05rVoC9gg7eagtBhHteTg8FYBlRIc2Elw2
UvicXkRtnxYpUFF9z7CJxOxaWm/iYg1riL8DHoUPZqRFQSp4dSBcpGCUGhlD
dzRTjm5+QtXiae2WS/iHsCqm9gbZDTgKAzojEYj/14uFOxWz8HWy/1z2QxsN
u9cqfYTdCCQ3ouZM2hw0mstadNnM1Zz3EXlJcrMX7LXYiFBMgRC/X2tEttnK
YjtGfn58LywuXk0qR/QkRzFbJSxURBq6Gj82cM2vCowb4MXfzIZvBcCSlOu/
MWwJZLtbmIAvts9uNHTta44GarIGJl0qu8NvwMcu7gx/sOBX8ye7iJH9CPFQ
FM483uvMOK/QvF/FbAG7AkiRmkf7h9N7zOXOmMQzVaQspFuOtXAbBgX1Rp/x
wUGilhlRm31Mdj+RG1JgezI0fvLb3gjRPjxs5cIkqHe5hfWZiUGhp25aPQZN
A/++12OOCuKUmDel/vHGX9YzRTSkda+e6WIcL0964xa4fp6tiXH/k7pR1zfD
xZ7ldqVvL3mIy/YeuQqmS35QoH0pBZsDuaO9mBIGeiKKqk/WLBRrjEOsF0AL
p2urQ245rvHyiIZ2+T11ctfx4kbh4utgE/QBo20UIHcJmHDl2DyRxgcGwMWd
ewyAZHLEEToWr7gNchfcHHx+kEh/kCsz68G7h/1+Z+EMQqzBiE97xYycYX21
PU4J1+B9M+WRCMahiknVj1A1CFA0t579EJ0lrVhArhGzqKd+sicSsSiJxLBN
BFlj4KPsQ9/9gVjDOZuqoM3sFHxYMdYa+rqvR9MpfbH2KgW24vVziuwtn587
thAgh8xNJF1BzazHQrPYuRyQI6jZ4/+HTA6Uh0PRHfDrW4UGLrn/dHR6jY0o
fqX+wBq1VPRFLf54GDX/YGChoRXBqzlsHYnYlhcJL/JQzldDyXh3GQcVKb6c
0fHdep4Pp+SmvZL91yeLP2tn6kP3OPRDTkUm4LMmOnUTnBTKsnPl82M8q1CI
fJ6KTtPanBtReaBzTRuG6MrXbIxIkuXrk9pHq8aS17THcn/Ec2KbcEvqRUU6
ThKy6MQL4Wa6YbqxKoCeDANAkKS3gUHt2Ra5JONjN7SPety21D2CSO8TVwSg
fpO9A1RmfME7KoH/MOrokrSAzWikh/l1OpB9dE3ewxJ4cGfSYbfPk7Ab7jyo
8Vy/+fcAFNvtWWyYTKy1Ytm9rApJ1RCv1pskOJNZe388Eo2cK6wvmkAhm+Zb
HYRl5Us66kacOtsxdk6iw7AOsA4g231ifietc/KyX/+jnUiWz0DCt/S9+tJ2
1tyiyEr17NtpSKWBqswxe6HIQmvxtGiKNhxJ8IxzVebItnoJxezenLJ5T6T2
eu6+8/I8NL33GdwL7vQyYRncigp20MYc18Vn0Y9VkjbRITjiumzezlAfSemO
DOC+MW+/8sZ99EH3+p0X/ToiKohVTL/7zZnnfqFHbrodV+lC+fHiDF5QKka1
rHren1A4LoLRaBxgSNhicsNrWyxYNHcT+5tDfVa0vDqUqu2AVWWtF3A86Kpj
LkzkHJAKwfTA1J4S/SUqz2fRqAyIlDhrWZrsDmDfgxy88I/GQfuFyoq1jG5G
VseB5qnwQc5Pi5G0CasTW0CYwibN9IhX+ZsmIRh0SURDYDw6WJIWMUKGxzSx
0FOgwFpfJeV7KoNwq1ozqyElMpi3o4+aFG5le2PQyS/J4or6VuTzJYR/hmiA
zDsaqrRadivG/5E6Q9xfXZ7RhzB/i+D9Sx9pL/73SKZeTJAMqQkzIr40gYGs
gNbCQKVwh/fZgZGn8lwY6z37B5NrMnwWACs7uEivRAoBJnIk//zvc8yzYBXN
2+JFDJNelr3gDcDbHNM+Pt5qSU8ImFMKfKdCLO8YZjXGJGdZWRFd0CJIEY7l
aAEe8kupU7rDg2gerQ3pznoHWGizR6WGcYn5M0XdkTsi/Kom/omGfmCvl1Rr
uPAtDAOy8WeFNFCOmoQinD/8y3ywV9Pu29wBegZUU7b9/I9Qrpz9tNavc9Ho
wwAvFpt2oXs/mXYIQVdnDNR7IlG5u+4qxIhdo7urU/wpiFm9EN/jzaD0GC+e
WdDyYslbcWbsA+w4cW829ZuwfEwqOucy0XC9RKgO9wVRKtvID4h1s0w3unnH
+FLwkwlTJ/WnYUCiLJqoS9fhEiS0Mc3bSRlGcReH3zlJ1Y+cBVeMggUrAYT2
naFdS1hk6wzoBiEph78coH/knr3AObGU/Znilf/sRmiwkyeEsDKodJjyiZXK
Fw+8zIrDqCXcXyGTVqOp0waFgDYtubTj3f1hxxRHlOPgI3bLiPN30JnbuFwx
/EbTJ7evcIaARaejTmegX9qlnqfpwi8JwzaXMNhmFjjn8PlBMCiA2uy+C+V1
brO05S1sPe3oAdxOchmaYf7xgmD7Deqgz+sgcJYHnJ+SNoQEgtNlHmO0u1Yp
3T5jSVafcWu1xC0VXQDslfEndbMPgoUIZhPomQV4T9MiPEc8GdKipid4gwCb
/h7PYLw1S2VQnZUBN6VF+b/bNdPjdFUPFvnkG6kSfTdz+BPkgXxImDIl/Dlb
RQYi+0Ead6I9LXJuD6veLA1dbDCqfZxUZbCZw9oPX2+m1JU7gOnDhTZekmin
0+jnXwCQ9mafbO4afk3JxfQEZzw0M+/IzbuyBJEjMnZfXk5Gqa9vteBHDDmF
Fev2IXXFvjty9uxVFMPomKdp30MbAsSeXHKTtxpJnyQJ98ZnfH4/ARHjfZv3
kAsH/U/krzuvfTzMxGSXzK6VmN3t+yYtTlikplpC+a9RrimOGSTA748ofVQv
LrgF3cJcyigejezq5+dZ/ZR8et5MzFR7FPRVRnmYL9T5JBz7xn8puWB+YS6o
HPX5gq3b97TuP4I0pD3ToWz3q5wOMosYsbBCIh0g7d/nWdhPaqVRz92vRlTH
WhrPh3+wgWu31ggdYyonqWPY0Bnl0mM0nQBYnzhhw1MDBTQhal4cRVtRXr7a
YstMRaYMeekY346Puq4xBaLLsDtwD0sQkcdi9Hya/lS9wxyw04b5Ljqx5jHE
qwEJnfCzessK5q7UdFA+1WTyoU5Md6/fFeGKDFI0XD41U+M1/ljq5En9FJoh
N4Ei/xoedBgEh+xqiqbYiFYWWEd7Dfxm3wJa82lQ9t6BVrNr63vaJfpJixim
8MWo4vazcM9ynO1IEUjhzViwKlPBr9y/iDEjTKPM6hjPSBgeioc886Rlbt23
sYVZqMX3uw9eG5iq6GhZF6ay+p3ArL+V9t9zQUfJflCZRiffqXEC2Gd7dIVw
enSgfLf/xe+uZY5Fyoq6b4uyRiqkBX/Yffn/bllD9pKsSV6hr1Et+U5A2kKS
/zJKcTH51SsgLoenxlZRIiuHkhYy2/VGTVoSgVtBLO7PgVgnC7T6LDtaLGB8
tlml8P5Pdt5MYtb2ounqw4HfEv1D6Sb9E9hVp2InQnVbrpbyTDDCnGa+pXrp
uSBVBPbeTFaOzJtRGkF+h0cS1TuJsmkKcW/jlQbE4UXXCC9Xwz8vESZUmmjq
Qshmud89zFvd2fHt/7Br9q6L8iKaNWni+vLs+FOZzBYwLOt2dQW00bpjb7uW
4I2jOEWyWCjE448OlT1t8VhOYUfIzZrWqtzmKa8A/Ye/Rc5DMYVLZ2W/G1ON
GrP9ne/5WWSarau+U4YhrTcmH+bX3nCBtJE904bJQy3HL1Te6iEa69O/eC6l
B2SWdJKVeBx+nC9Qmr2XKdmj4vGEgiORfkdaQlcwa4NGE/uiApYvM+gY+YAC
ncm135sJ9ADyY3/Nh48Hkx4aAj05Tz+PyJmTS2WZJ0pMBA97+lrdPxuUbkEo
l1cH1oZ2jz6W0ggm55rTpIWwJ1EtAD/Ht1Xx2Bi61XdpHRL8ygbieRBdC+mS
D6xAzU4suPyw+BK0WzZ8RDoA6dd8yQruRZ4VWcon6/fCRVeqS0AXII6swHOX
tN0CuTuBdUy/GOy3lPJoE/1MjDLQ5eGsV704IdRnGD0tkcun6Ql0kBH2fZ70
QajkdkFDcLocesFXULURdRPwJjNn9qb03+ukx/uOuyVg4XJH0CA9+34JczTT
hY4BxEXxOMtL/PVuCAciW0O0CQirnMvB8MWfChH/08TKzFLKGmXw37F6XaWO
dZmpBlWe5QXmftkq8T/VornFHfyqBur3qeuImI+NFdoIDwwFu0MCVJ0P+Y39
kGaEmLJD5sq+HqLqvxuG/hCfbXyvNAbovG0h+O9u6KDwTI60IHD4x8XZgaXN
/sDa7EeJB1hmPtxsWykobcw1/zWJk2kCjOESNwD0bmojwgazxBvd8PUs30H5
7O/AYcg70514k6LNU/jA2M2UHv+Hv24oFp9q69g9jT0F833WuD55rYvHBbPO
1/ymms9I6ezpOa/3uTgxMM404cK7RgbVOPBqbly6x6b6XM1YYLk9KsbmTqy+
x5XpeOjbY+pAvJLU0ULYiN5H7Rvf9MCU+WeGyigIPaUdlDTW1QIctszM3XNm
lTk8nBTuqaKmbtkEwu/ZtVrE5lQlLLunzONUsPKko0Qjd6+EbRWrxwPODpb6
xvLq36YXxQg8oxTC1oAiB8cIgnR5ZZZNTHwlbTnYsfq5Fe/YSm/1qnHKqqwB
8benWQbsIOniVc1XdtqOvYYkDrRl2yQbX1RzaZLrTgV+KAHTbw4fwdA6hbRD
kGCsoBbHQF+awn2/h3wD8uFooCylOcJfJaCYWvXrgIV1/Xmn8AXresTpxeTv
biXB0/yKxST8P4u0KV5uwqlQExjTz0T5+3aTiwBdkgNpZrnPbHEfpK4HL1Fp
YVlinkjpkCIUNFiNgk2FnDw4frHL3io7SgWcgrg4emKULl/ZMqjCGfMg8y0A
7d6LzuRKN9n5DRrV8ChfmV+Ls4LN2sqzxEAV/cE7RCT6aj/yFHNX0tvyY+Mg
6FbJ/Vuh+1xlXjYOY4WsCeihp3PQ99NUaJAo1xHPlTar/N174ndMkR1fTKYp
lCAfZMAmRGOK2TqVOzavDOcb0jy79r8Ya/BQYit6SKSulEWXF+5xsbo9Tqvs
2CVzsstWsD/rcoklGfVlUSonJd0SKn+mkvfgsc2ErO77pSdeijXYkK9qoB+M
+qxNHnI8CXBhwvvDq+U23PIhh9EFZBfDPnYCXEj4mRkyfzHOBQklP9dFQrCU
dEVNf6c/X8292IxWEYLCriipz5ZnCRg3cZ7Oc/w7AAhMSyILINx1Z74pPMO6
RIWYixmivvlinraHCThM6RN2hXbPQWHOEo0tCvX4omhSbi1L2ooM67A9d9Xs
sffQSP5qC5Au/i9HLUCbO3yTxQK6C6b+1Vy7o+xJwk0eUQa9ojzWzHrwFk3z
szPwtiNms7TAgUwhV+xUIu5IbZllMSDBP3Y+Hc0x7PNsDNscQd05z2UEI8zO
hFRJcUZb36QJT/Du9Qah00bXvtnQ9Jf+BIv7GElEFotDElGcJjradHLNQDWV
tQPMQyxAu/i6S0BtXqzpQzPCsHooTRriKZHX62O8Uu25Xe9125qMwoBOdH+D
uXjrcn2vp40jdgwtIHwbjix8G8myaC0PjYMKEoo1ibCcNcm/RjPcNn9faGdB
bBhe12Zr1QNqCVT7ZWoJ7TH98zpvnjsZWUgIMSstOm3LdBWWXuWYEbT6m5cu
Q3xBpbXcPji5SM78sY5aIyJejp/mFHn2pX696Up90dJqDPQEqPpYqxRqruOR
XeNJNYshviedpW6UeB0w/fltTRa+ntn45GVk3axn2r8BEkWE0EowIxq6NKaC
9McDU8szI3ZMkQz8C5SOdWDAuJNzM25OBEZtV9r5rOvE3BrkPT6/2nUOVw6i
k5WnCpUeeYnLDV27MTPhxSk8Y2Xlw1sHS9yiMV5ASjj7pA0bvG/PciDjRXXA
djqTeZzIAiZwmH0I2KFSbr1d+1UhPKZZcUk1YAH9Wa5HwFWB1cuevOHQnKW8
9uupD72hkmJo23qsGYX4SGWcg/FrMnarO6E6ZzALPnjJfzeSknCClTxptEAu
I7M8mi969cMI/i+GyVlvvrqrOcvlN+zTWtHGC6HtCjP3RHTYozqYi+mDG2hA
Dq3WyvU1H0xx4ViZ/ltGmtlYqXV51UpzCUrJ6GkbzJ3L9NDtleYqehV2s7CC
TyPAvCYbj4EgFCL+MbgK2/X9T7quXMdshgWYE0ysW0xU9CLIpsjMi0c7ie0W
ZWrhaIPaBhbjDPjF5CRsfFVYEgUeOAkKAKrMVRk6D4PiIPxep2HMHrVUcHdr
ikDw7Oxw5dLJkjGYxRsYVRC215TJf5lhnh8z2N4UfH9TgbKia6PI56ioLRhU
EwLDPBGzERSfGRu9pV3Z3Jc+mEDcq5fOFey45EsqUCp4rDIo4c2kqzo6h9iB
PVjbO5eE+nhPhfnRJJpFRdjyYTpo0aKg7HUutQBoh2ln3MRVmZQpJBDJ3g0k
j6Pc/n04iqzQS0FyTPvl5FgKsBNJIp9+CkEceYYaH2ODaJJYokD1N9CJQ4gM
BjslLrhqaSi6tKXsfY0SEW7BKTqDSuREejHVO5ZnIQbwenk04HrRedObIwFu
Q+oY8dtWcIL6/BgFzEHsZwVccRXyG9rJJvlyIedFDCTvZRH5mfSM6+AGM0Lt
Qi8IzKeUZdvhAL3XWIKW47tAYVXpSq4lwyGolzBeztuNapw5aof8c2sGF20D
GyJJJ77k7oHMKa5Yrc+pbssYwVt/1sk3P/5j97ciRszDQntUHcRseYFOW0Gm
ecIgRnz0NOw9SXhrUWC/QWqFLMyTKMsOW7yDuDX2Pxy+hP3/3CGwDAJkiFcn
IJlfNSJ7mVnJSzMel8NzJz/0cBcuU/WRTCr7cvgInxqGfLIiNWLdY35Bm0KM
g27k/k5YGknQm3b+FMBFzJAQOkBHYcZL+obmV3unSTmuzoY2c06KDk7vfRnl
mOjgqXHYz5JQAUh59mXWhV5ZRx0pHWVB8Vr45fnfoAJLH/HVqSb2zaojjeRV
0uP0nb+JjtDTwBVPhVgaUlfXYsuu0VEYAKgeh2AEBvOGATg0VsYaG6WBQ1Zh
eQylZQobFue2ZEajpR43ATIrzbG53ecM4pD+Yfx/FRb1W2MlTYLIHx0k0e0Q
KwN4R2oMfl89VPm1GmXUhFnbEy1HX70hLmVK+jrVQBG8pvL/cO9d9k0VnkUr
Bfj3S9Pzd1CVxF7HQKE7mDg7FQLaOo03AxUr8xLi3ckFR3Sm8PLFxR1HNvOg
GAB9/NrcJkPXtcxVxrFDLb3k9BmxE5kCramv++6PaNRhRvidl/nVISbVyR0E
rSvvbLYJaQKA6lxJCQJzkYxUL7c7m1DPs+6rEoZ4ywnDQK4qCfSutpbPmRsV
uy8kH62stUwWiaKxMy+Qxs+S7v9TZIcqX/3mByQnntu26z+fw+7WHwEERCPf
AQzrroribnW6jE4H+cnZeXcTPME2y91P+RfAoqA8DbuMvJ7k5J3Bx/iyuy3X
P67c7YUlPxb/+YoefhQ9jEvNo7oY/yPVGmkYQulb3nIWIlFofcgzsQvSWbwY
jpHgg9sN0tF3MOmUeLfagZ9YzpyHUTSlBLyTiDJTv7tJPon/RmGuEj2jXdgO
Rc7D8HN5nQtnC/3Jl7/3tKxGeYDP7zdMsehCpB9Jq893ids/dWTxWNd1YBpZ
Y+WkYO1xWx3aIQz1YYDhDGbp6yATn+ramGKkCOJKrWH3SlMzkvYvA5Uhv3vi
ksFysyKhRey0MAPm2c5AE/JXZEa6VjuGsZVFOHFsCSvHrbBEcLPff1W1p98D
IUOQcrCC7j8leHOKSJCg6jBlN6pwvu5b4e6kywZ8bsrWE0U7EhoyOkkx97gd
DSEMT8cndApIzDGOCB/GaGQL788XcFgmcdkCcmLZiOrQ99D014jaj3jQ1f2L
qEzh03n+wvol9NEN7p9zDzloRzb5EOEYLjplAwzIsnynySuVQs9W7MLza4UG
cCaIs6KW6t3bYamxLCShFAMR+og+MOzHEBEu6QFaH2KBmNPsZYBFhsiEgrpI
NEX7HoSnz9cPZnDQ6dK+w/qa5JdypaHaV3EQBdi+UheIbNXgXQ42ZSp3XxZD
GGJu896WzQi1Ax2SrUXG/33G/r5AxloON/Tc7yK6MeEwX0T5yybrL0VZzSd0
IvD6PzZE65PH9BKrUzo3iyoFbm0UV6CjBDDt6z9ow9OB6KMay1ZPrzlvncW2
KkR/+y7bnShdjP8vWZsnJ+UntIsC4R+4owrVvckkyULqbcgCW1gOEy8Y1N6e
yuIVeGuidOCFMRMDgmZT7+svgtwXyFvOshZF8F9jHdXSrXStljsz33N4pwVE
FcmEj51ZANghTRfR94M1IcJEENycpCT8gVfAAo2OV6xrrPUH7yaRrhQn3E8e
OR+aOYC+Ske1d9MtyLJ2k9Ghno34GhFsSqvEkBCnCHMP2qLorYB1a3MCjyg2
Zx/p8kyshJO2DffeECy/j0sTfN40rBmgA/VUPZ2mop2O+fiq8erfLGTxIw6E
HuaZjsMMjIs5ym0AzWa3ugGy38GVqWuDrG6NIff2SUZSwOE2KYuQVGMjTUbE
9xMleSrWed9juWrLQIst0mIIlnwC2cukHXI6UPhGs4as7X7bSZd1RZYiB6Dq
UjwRjMdYIuigEeTypo3AyAx/Igw5OWHIrSM/B3WcHBp/9fZqWXvUazIrcJUa
WAB+zxgncn1dAs1ts4Ei0gG0vDaurt3Xr6ChqmqBKEe5rPThlXR5rD8lsrQd
+l7IV4RamQw307A1H87zOstN4wVw2XOIuSN5RicMjrDBSusvfTcF+LUfs+ft
WHU3xu9hWkxFLtjugW4fY0pCnC8KQrOmq+bOrv/V+Bcl5JIgUCU025zK8lo4
Q4j2jg25S3L+DDn5AEmyEuWvCKXPKOxXDXeeMI77WM4RpG3mO6FR6bZK1vt4
yV8CU492DuyeJq/vx0dHwPArTjZDS0ldgmM3ZgH+UZjC1V2mn6azPUNRaEB2
XbbovsHv8YZKiBrqF+tWat2ZUlBP+BvUWZ6WA3ChKRI2vOPNkrPBmcWNoIXn
QZqdiA7pUjKmqFoKIM0BiLUwAnH7dsPyIyKV41u+e4ddO4Ex/fAndA5j1Xx4
0Y7MAXklPC309+KRjSMmd+ZBxJVF+TZefo6+4AFxexRWkaNkfYNGB+2dpGyj
bsYwPow01JMayIPwrHSNV2oi83H3/nMcoYq9QvlFEnTMPuW83Y4wvDkUsckn
CoMwEBqUgKcC4M+uZ2ySOpeoNvB8boqB7R2CMW7APynjeiS0ls7+b6m84v8Y
1WePhMzOKonbpBpfKiRTRyc6sTaUx74GMTCyg3b3SCaW11UPubpm0wYUZDG/
iDudz8S21a16BqqwyO8Mla8nmj18uyG9t8Z/GPEFXynnon62PJTJ6SoESuR6
bFpAayv6I2bVvn5Y1/Jl8XPLp+A/AUavXbOcL3stHMWfepKH4Ic5ITUkBtSq
caPXL6jbas50NUhPhwN6O8yka8c+0TeyB66LnbHsF61WiDllch4snGpUhBlk
D8tKTo7Ea8Kmkgmgu9IGlA0YJ8SmI2EglIRij/bsJcKv19wYL1r1BGGCaQHv
6RasdEohiMVNfGUA+LCY4bXnrX0QuNajHGk5+SiUz7hiZsyQXhlxR6xtKWmA
LGIOzl9BPwsUGt8mKG1oP+fWFdhbzpgoQu90cWNRqwqTn4yk4RRrIOn53PpP
PPSktiTpbAFgnHAgAzkA8KBZIwI3iCt9uW1tAX9zhgBumMiUfWWQ6dmRheso
/LAibjqhOJ7lxDhgtGCZ0b7qSPnnL3OAb25Z8wSm1VLbTkF7KrNMdvolBL7g
fbAalsKKGKVeAQZf7KH8LFbOKnw3qnOqO4lGOcOhu+/KjZ6pEph1UIru1I65
2T62bUvwEm6Tpl7U4DO9dZVEfvvkpMlqM9DCwjdjgdysZvpfIg6km3nUCRja
nj9iwwIm6+akWnL4xrw5ABugxkNyA3xfvhFRgtAuUqIhgzu19GjI+Fj3vsI6
AczvRcVVNa4zPxij5/ZHn7WR42f0C3ITKYBkhs37lyOCXLjYlqNFjwkBeSXk
GgeWTz66jrjqzf4DDTXFr519lRIHlx4QNoJ1IcVHHRYKJ0DjSiY9H+yfVOc6
IZo2u8NrQGYtHfIumm5EC+roMBk/PY0XtZiZq1s+d4iS+x5NKCj4+g+/Lf4V
qPo1x73oU3x3QmzDk++D5Y8y9l9pgDvhnGoRZhP4G/+Quc4sNnY2pEQKHxlq
NA+FDDve8kmrUBVF1tpMJP9636DYNtf4wpJZuesGkklPR0lg1RNaQdkHjreH
xOTuPSZsKbDFAXfLCZXhPtV0gR2nK2AOVJOdkIi7Kxt8IqNhZfothJ9f6BwZ
K3Q5n9NaKJ3IPmGnLEpAeya2Xy0n4jrdpzcCIWZ4Zh2Mkh7C612hY0BFRZyy
4HIZUbCou3QE/uneS2gBviKS9Y240sr8cP20obUgIphomZSuq10AW66QNeBa
/AH9ScTiSgvV5Jgd1rT+9Ga07X7eOMlHANaAIELk/0DdOl+/gt7pm/EbNdW8
6LCTIfqxkX5uCkv0OZivXVj0YVRkAA3oov7GFEKlU6WHeLv7KbpsNeBfNpo1
4ynXvFH0zraqwb1XOXupQL8TpgU1xaGahSMSO+Ueg+bo5LqdBCe2QRQyLGpj
zzH4iJb9Pd4tsjO90PNcM48TCK0WfDjJjVPgoIOO0/ouP10fszivxYyXriR3
4B6pXMhBI3q5a3X82SXdMBBqZGR5C+/8utKfo3reYCjyoKTJr8cfWhwN+0l4
7tao/8fmZ1dMm3zyHYva9kAO0Er469ICuHEtIhDZmblICp7lA/BTH5qn/W4J
vZeUHvVXj/78VjnuMMAgKRKGgVBm/THv8HTAOAY1OLVtU40Qa2f4V7muUaAb
n3DwPX3yKUwIkWXmOraTnUqTWeaF+l11UvlLl7lIDnoGk4unds7HWhD5wupW
rDJd+xx/SmMx5rx7XsopKHd+p2gk6yUGy/sj1qydexbY3wF93lnq5vVwxvWo
+TqMePWY/79yJBnjBd7lqwikzqif58ztiIEgC9sq63tZRI30URw7ZauHUiUS
Uh7uJ2xnsVy2AmtHCwAg798LelEpmm+AwFy4uaSiRUnuqNe9o6wnHcPqz2cr
zYCZXBagTYr+WxTHZPK7uE8a+BzR5M7JVARX5f5B3pl38NsfBQ6Oi2DyTYKt
AjZpeV/08riJ6lZbp8GdGLzkP1tYKMOGCng6SXZHpgLJqtXGp24I8dFkGI73
ZwJElhbWra8eQO2EbLyd4wB6pVoTWMIlQhi+VyZl4/2Grt2+4oGEJlLNlDoE
SrkR0N+u4oSOhdOJpzmVEyWizymOvoL5L2l/+BAW9s0rXcVrwCbraNdTINHC
UhDN6virsKSmlOTScOBMH/mA7VlIDYT7qBCZE+t3FPpsKX1bDq4ndmjZnTlA
weUGJ2kZwVddqABk0hRGIrBqvRbMH96yYll40DJqKruNsW7NTJYOOe379JfL
Zyj5SBfdlWeEEBu57Ji8V38YkBCo32koAb6Gdiu0g/+uICEJ7CoyTdi6W4YR
TGeJLp4mfI/t0KwH5572eBibnicoqpfmH6YEi6etPjlEGo9I1OyIBxbbDaCM
W2StqXvLIYyFAuyisbISxwpZnwAMSg23iSsK6rMUeLW8usrpHrVA/+wU0nys
TMXyxZcbkPzcaiQAXWFuLSd6rltHfS2H95zMlD7i07vXIwef/AKWFLNBFqff
06belCi2or3XHKFqN6ZCzVzOR1vbDbtNtewdDtljLfsGSqk9YxAz3F43kq9K
VMEuOb/uauijRQjyuoz/s6Ywk+r3PKoDlcUW7sZabjSZC6w6cKlmEGYBUnmd
KhJ0mOqrYJJIfRFumDUV9hppJLGYKj2FPMrJIXhiMBIKtKXvTUPkVhein3Ri
WmYHwkvlTV6ocy0Lkq6buhS7bfJrMLjTY+qzFk7ahzI2Tf0cz53iW1to+26X
LA2R+Rk9hhWmYV9KbS9fdl5TQZl0/MMXz7Pi7Jls1ht5ZUxBeby/bvkE2iN5
KpkjJTLoXxiTkdrAj1zkBV76VyG4tdE+1b9k3S0y38pj1dnsodSzmgmfTorb
P/Yq2+oDdlQtmS5p+QjsaHs+pSCoyTvd32VrEtve/sUf2hSJY8e9u1/nfBwk
MRwDjvAILoNYXJaY6oPN1AQXpjF2zqVLKYekXCFWh0AWVImzYhQOQu7ePfyR
eLnIzT8V4oLohTqmdEjaZ1vbtAsqaTjWSMX8pOxZo9yLibAP7QoeRxec4y7P
BnbKA5bes4iR/ZUWOXJ+ejF+bSqhBuuBz3a4CMEj5sTdLUxvA7ZzrkSBrqCd
cGDwOoQEwH01fWfWe5rIZrsOBZxEjdBthJv9i1P9edhHjhLbfceW3mlPa/6s
bqzDKUmaETywWQLRfjuhFzc5aBXCiCmG3eF9l/2KKV75YQF4XwUhvrpYIRez
Ed7rvP5v/8lovF8GGX1SnK6n3BV7YqltTIInqjGaxL0QDeqz5VYqr/irCZ5G
hs8JeGefPJigQJzB9cVdsTdy/ufKnhGKHkZWZIIuynk2J/iTphW1TzgKgKi2
ka7n7u0RDPVZrs2uqnb/zrq3EMDHLlB2e73g2sHbf7EQmjCeYSq1i0XzvADs
CYdz94TKvog500zCFQx1bcSigCpkFNolA6uW/fOIfvC3k/Wy4R4nC2yjjGar
95UNV8oj2HAJw4VBaVCNy8KDLGCKS3rCk/kcDw8LX1coe9sONmqj1zHu3RbT
6EUt0G01r1A4n0j/oC8tvHnwCBmUOo6XXkUj1qOGi14DFdQUnvOWxFdIOClW
GhMJ634FQL6lz53r7kiBPPx/EeNQWLBVaXLI4FuOY/qfEEK8b5kEdBgCY/Yd
0d/eUMvwKMGAnEHa3kCaRbD4RbEyJmE4MUkWdfxgevBzwjyK46ckCjF68xmD
foc3lpNX2o0GXs1qP60vpusgZWo2XM27sTPn3u6T9ngELiu4bACciKtO2t0M
b6hWr8XLQwpik0UUPTKPsbMkbmrozFIWozlhGxDDz/pOp5TD1xc741EbdzNa
Xw0LhFxI04vpU++Fe0qgfCcc32F1haIjrd+40tr5oNNmRZAdFVLlowflaw2V
jLoX/sZf8+zzHcmJZwCBwP3e4RTbd11XjBcagc/vSs1fHWfX7oM5zNWOd0DH
F3dBdvB2UAbcsBefhvkc58IQ628/tDqFi9zKbBITb2xODwJF3VPEX3oE8vqe
coMSCEdsNQPGGYDS3jR0gU506bc62nhDUfN/iKb/T5czh3qMcYuIp96w4NGg
l+knKxhqpJADSBdfb6iVI5BwNOi5JWw0Qb+GWrn6AmmQtQ+2ot6RnXlTeNgP
+O3pxcHeDYZDPlB/8UMdLSUdAfA4pSkakrLbSSbuNPo+UzZuqsQmtrSdIT0R
NiikXKMa98/GSzI8P6DpU9hxWX5Z/Uch6jk/IgV8MuTW4mXKSBOYT1KnSaqG
fAqN7O6e+G2NO3MNohnSJDN2N6KJPhGQpanIyrCgKe8BBQLgOkXOAmGwagUJ
yoq9gcFUkYKJ89X2ThpGfBmjDxSS7ipQOAbw8/UqVmJadRNmEKaSCvrSWc6X
Hr8+HJPTL4MEcUTEXCTSH8Q/1uMUWqkSpHtC1VbATCjXqbSYD58dLstVhgSn
+WEtix1+0yDenRn/fMySRwDf+nBuXAyBsP8+2urlQ3R4XPwvdIANrTI/KrjZ
kNbEFpDLPdIqWe9fPF8rNgSzU9IRJtQuKMo2aBE5PDfbvEoGGULxLfWrjs6D
KbBNfbI9ZUOiTEzGw9Dlmm+qIb7Rmwhu+uOJ6BGCnyQNqjkfaw0Yg/C7fndM
eDGnek9ji3QieJXjoD99vmKryLi8CMd7eh4yyxHVOMr0L4VVThAB8UWWXfzu
tPRV8cfhGPN6Thit9G4lFbSa+qc43moEbvyv/rhPZ7SQMVmFh34KiDKt7whc
aDL8kJk2BMZPORi3yGtfg0v5mRvs7Jz+C9bMJ2iW5Cxwg0ZBHIvQYyEFFwQZ
HsRfxGOhMRmhArTB3xmmEj/qVHlw3rjJFVQfwg5+7QEFbo127VIhGPeiHY3J
gkL2ISQcgN6a482m8Ypiwrbdjc0Lx6lkzMpPcMEXKprmhnIw5+NJF3t3pn84
KNdPNLp4M5j4IoylGclgOBmUTnJof51K6So3EylX6BwBSFWKChX4Q3U0bpTA
doky+rFhuH99GC0iPm2wfcR0/iREEVifF3Z4kZwL4zjblDiahrGBfEwqQ9JL
XTPsaxV75myUg1cIMkxEvDI+7IC5hre60avX7qsfOSOdBiD766/7khwTt7Le
Qh5OSsLgzVJR6hrA5xuA2HDzgYRIfHJsLuiEJV1xYuBzCqrokfq4JcUBlDPA
FuL0N3VyBabl9sWHtdcxSRJQX7EsPiClAOtMce6cdT8ntOwm8QKjOJW7WyHC
KCQSm0k74RfQuT8B5JplIUaA5MeZ9YvKCeMFaQlNX/+uWPAiTpybnI91Cwv0
+IJFFp5kWvjf59qCfRhcMSWisv2DXeRq+SK5+Puck/hOr3lmcz4Q7O65gTx/
7mIQQqr0+fRhtbtWtNgDFHWZ9T2hcxAuP3yMlus8qnC2/0Acl2JnRjbj+Ux8
fnH3ohG001QYOhTIiTLYGVUSRsez4sHjjup4i6CIiQ3gn21gsl/DrtWISCWj
D9jYXScp/ltMu+R8HiQSavjD3F/vDIFUQzFmsz7dP7mpdUKzNHprxinQvKeC
jlyFG6LEE5nO/r4mLL1hypkLuQ/1Z2OD3KSnFuzykpwGzMCpTwobh1xhNrfP
rwt/rNWa7LLzi6x5Ir70hcxW0681TngYgNsri/o5/FWNDZxQXMNkwDySLLV7
hktU96ABaS+IeM/wcNNwwwJRw111VHrcoYDCMfC1G9SXO2yp99OX7I3aXPKI
aHq8eCnLSUwd8fFp2p7BJP2UZm/e2YkDFi1gfPL0AwqmB52hoWWmZoYheeTx
P/0tiEF95iGtzwOOu86zvWIUmqCKw9hOd0XBtI+qjjxExizM9L5QGJsx8iZ/
W5O3ojicOqCEpiPhKz9cas/UpUn/WiaL7+9kRlRyPwnPCzKE2QEjvyDWn/U+
Jvzg9/qvry9oVCTtW6bdnFPuMRHduyrzzRxgpbjnC+HUk5LNn2t39ehkdRup
r9VcCxbJl7NOTtUgo0UhxQOsjHmV2rduUitBe8Kg9NzteI4nFPr+peWkyhS7
AEZfrUu9U4adkqzEEBcioldUf7SQ73oROPVRm0olx2lhp9ajYMEu2mcJ0FLk
gSHqJtrYRfdqp/Q9ySlKTx2f0eKNPhRp1hQ0jqpGtGAxShJpNaef110psJYZ
A/OUyNlUwReIW+XKhdQ8OiwaYTMhFw4x0TwiaZ+uORPd2iO0Nr3mAkCx2Rz+
20PNxM6diGU5JbyfyYHBw4Y3V7l8vcK2lzrkx6XXOUajjtjOweOSv/t3WDg2
0JrG/qgRnBppD3jjXgRxLWolwwGIMxGW0709x23RTOpXO5XEDETwbBAzbGKr
T08bL9WkUEwT5125ouH0fgkEQDdu/Cu+hNbdmsG0PxqDBN0r/a8D/Gh/wFNe
YCDWkWAGVCpEDQlkBuC7L7TuKQJCM+Y2IYNQKd9ZLlXKgGcxBSY7yjvEQauO
oflZumeFF3/yLUGdNYMLzvyS0ZO+vh8M5EvbPxhiObB36lBSdArVbzTywQZP
ofgx1UB6tLjZn30XsafaW8UydwBAdig9rLzL1c247tAc1XZNikZB04EJcXxs
Ga34cCG4nExoJFOaM3OEguvSVzlARv8cHd9lv+a6+i5W5nWZR6h3rkZsPHth
+DIj79dVVp3kiY3e8VV1f+JhNm1J6T5Om3zAYrjiDrsZ9rFQjkTzWMMbr01K
EhCK9R+1l6EP2/Lez2gpgNn+acLOtmpAZ0BqFOWi5AEo2lMka1SvkLM5zO8S
zl/2UuzW/jRurfLPS3nItnwfR4pYy80zaHF9vKx4FFHQ0Zi/9DNTn7yNYYzg
JxFY0do9pJEyolL66NZ4wAauBgB4FdH9hneGiyeoou9DIeK1RQ6TR4cnK7sV
8wPeyudqa01T3ywKMo9cfqmJxdaU9kbX++hS2x7DhvW+32hc/ahWZVtEn6x+
NEcVhwv7dt+C5B5mEVqyAjMU66/w2ED8FgEE63Jat+IyF9SlKtc7uYKXrV8/
RH+AHBbRojKqB5akCG5v5xBYmmmbRSgjRNlMnkNikpn+46dWhcXE83PLoPyJ
jpUn03Sa032Iu0gdP9xAg/3djf158fMalqkjJP5uJJE1RAdAuN7ozHt+/2N9
Yiz6/J5kjjfI2u+UrutTMtk2pAbqqnzrk6MIYXeopgIBbnn70vtZBGNO+NSf
/jWocuJc+3CumD9t6bt3FYJKrkdbffrulL1jefBnxP7VKlyHEKgv/R0a5uX6
u0PWSGK4d8llLXXZr1Kc3i3dwYiXm1P9oBVcDfc87Z3MF+476VCY6JrcgExg
cLqggkdZERDwIstFY1Qi1LWTIYpHSBNP370fOY9uMy1gAxXJ/mBWfJMgihfM
2skAAzOpNoN9Q8hwkaaaQOAJ3S5ABv/iAVtnhaTle5UGjtMeLWTEPIFLZIqP
6ZIKjpn15CgZ+4K8AGBHvWuJ6U/j6zn2yPWZ/clBKHuCApXsPMonbztcz5JM
hQ/1YeK1S+5dlZd/jTBR9DOrrpqhvN+N+6/nB4eQNPpNUYZzFaeWoCsYD+Bu
B1ql/Gm964TeDSqWOnqHnFoymXlan4TU0RowlVtqBgpNoAekRj0ojZ6E76g2
dVWUAnH1dM7mETkfy+O139FAsUkdcznt7EG4+mss9Ybumn/G/Gu1zo58GO6O
2VDD1v4vzE0UyxMhAo6C9s0+rdEbERCihoLGskQPMY2bdDsqteyQS8bX8B/u
Z4tNSlDpjjBjyYYmt0cMt/7gBmeFN5hqkQnqhossMvk8R6L/CitI7TUcfeP1
WlZkd0a/2AgBmXMZtwzRK3gF5SokLsCJoai/2THrsTZTJth0u6shZhXWyqPO
WytHIm4ABz/jv4rqusddjLYmuqVFF3/0x6srn5kgvbz3xesZzzqpxSsKatTR
5wYMQrjJxi/9ERPHWAX3GW5cgWwjWURapurZIXcglACwudGDotXI7jRK8PqF
iXA0F+V4G7XhYiQtzwWRchoFFFqJZNuod+6K3d+NOgMvb4C0NkH1xH4lxCDA
o76sf8Y4zKCnPJJ1Y3RfrCzT2lfAI3tJ4xit0eE3UkLBV+3lOTHfDBFrxGis
lMUKx8W/lLcjBPJvBlNedeVsAYlKXk9Hxh8hadz4rCe95QPg7v03hH6Kghji
he35P66DTNdgaV3aJ6DCiNr9hx33LtC8SnoD739TpoY7rZXXPe1zjEZoAFw4
wn8M9AiMWcmPU5GUfLUi9QMmNl/91ARod+5NG8miXgKNO8XW24eJFETBgcS1
8+q1Tr0lGwajQva/2lFgq8jEqDyuiCRF/UT4ebmFLJVKkHBlU9pMo4+cZBok
JYTZMTewL6G8b5uUomxj+EiPckY/fELdKntPEjY277usTMhgM12cK3UQX9bv
cp9nheeOv2Xek9/Tm8gT26Bh/MiXCVWIitqeAOsQRwr3MsLS956VNnvRt4Im
RmU0LdbajhSIugV8U2TpJuXiWR+abOW3TaEJQqptnsGSgHmEQ12zsEhMr5UI
nYrzi2ySN38PyUjg9uuGRDoLDkAO12KcXG0cEQxG0SE3XYrYRyfCt369sYpB
8TQCuboiDtPEDwC2ejxdxX94RKzy28QB+tuaKaY38rHpwK03v+v/aaKRMTXD
S3SoXtQb8LXrRBt5ebw8Gw8ORx0bPW+j9rv9BC0UV8CXNpEVaMjp24WPHln7
4qHorJLPyqiiTPJ8r7HW7ylpRkogsOiH4OSpzI7RYfIkPepwDn4qPHmiIctk
6agPEICF62BDQhKhcyWMsbZHh07ZBvVBAcryBuPCLHwtohtENEhpO6u99i+u
Gu6ez+9MqLhqfd7MJOBx1RkTC1y8s7vyXplsle6eGuJLdwyUjOKQdjelD9pT
J/Ge5jkh9h7TA2e9hkhxQH6PGFEKKuuub/A1+5Ffva5P+STZXxjqH/QkAw4R
GybhI/YEwt4fCCs4Cd8u/+voNmzncJNAkvT5Y7rsu0fydNJ1crexaJHRkD7h
Cid+1xVNKMBYlCLZDNcE8LZFuyW5WYxROTYyTg4w0fhNeX0SQ6i1OCpjUGVg
qpnUfxhR3ksW0POQAASKZiiSN8A2grZvis7HYP0XA7ldBjS9TyPSGfunSJ+U
o/818ONt5AopNMpTJfmaXc4wylivkQ5u0LSwH47ORAwDSeUNdhnZLgzIYEua
4KaSjBWglyKXDVXoz/4lXs3GfWD1X+xiZUnzi5oKdcEEi5cJ+35Pru6c2vR0
FgNeDKzW3nhl6R2kG3/c6bpIIryhxxVvTf6762sQJVffFt2YBvXFA3panSio
j1E3HDuaTR2rw1L8NJGx8sqLH/Fp3i0ST3ewTNpknwL8ysvLTGMF3GSxM7mO
jl7UpMB/B/I6y8cme3rdEoH+TLhMxdjzQxrM35ClgzwVCy/+ufsJFIxdMbvp
8d31n9pXc+TgHWUN9uJ92iP8oWIdmcdW6ysj/B0q1hMFhvNy2Ln9jnbUnYAs
+01yOwr5sRBPTi3kqXTezzfMDZwdsoPjkOFp0lQX2NluiasNE/RvzXWAZfZQ
z+wZrnQzkfM5jrT1t1ncm7krKaZrCl41kPNEh1TuDvM5hD4TShb01fBZnAx4
wOQe3q8fLiHMFXckGttvLOFYsLmUJqA74EC/kNBssninJyWJKBwUipY8Ye/U
lFjINfi4LpD1Sfsi3O3BFQGoJcTEfdWJKzP2Uq/gTH/MC67eWSZvM17Y3Agc
TQRrHyWC5GPymquqaukjGwJH8GzfRWuRGusySmp4mh5/eAh3KPS0UOqKIs+3
/L0pZMv2zNDhi4Eflj4KZxksi9QHYHLD39S1RdjnmIXD10V25D4mAKUZM98J
Fwn3pVpgDruypoNfUobfNGffS/BWCIkt0+5nnfh0dDNOvLZvwsdpxfgMT3aQ
J3jaQ3yj0fuadLctn29OD0VcmbJGLQwUwoZUzoxccX8aLqSNR9nuH0XExHiq
GsSZOa6hE4ZFT71UMTEloDnbpcajebfnvz88PcYyNbkmYv25D5xpvUBgp/fM
sM29Q7Do5xUARup5NLxByy1/sflqlMPoxClMcPqnchtMWacRyZ23wVLcvMH3
jSRmVt3aFTSh2jwl6Rj3FGmVPApSrqhUy90wZbpWY6qcXp+FCYk4MK52/Num
Rwevg+yJWCcbqcLZJCRpzfSCO2XP5CGdPxNNnay55KXChbm4y1zdh2hhp2R8
PLj24NFXN02Xo+3gu0qNgJU3Y4SFcGiCRIi33eLWaiXDiB5A/ZYJXL7I4brr
mPiCyh5Dhqn/bAMyL5anUrFBiNxEkvfDSBHFHe1gmRlKeHp6dryFXRaoGQ7N
CgtkmKMO6rUr59VgNaP6s8m/vrzcOmayEGI0e/syghO1+IMQVZrNkU7DgQ6L
zhS4r3CzZoRYge2gCLsTm5BJJrkJ8Avojb1aYF5LAOfulFx2sQAZ5UTyKBnT
5a6E/G1+8MrA0QyMwT8J7pMTFuaqp473fWinScfXRQRAw8/hDZmdd9j6ouwD
L46Yg/OD1aC4n2aPuDhlSHsmz/GRKQHSQam0v94H5cMatc9PV7T3sZ+EiOif
25gAyVI9Fyf8dgNj8aegVowA34QZ50SiuSNuXnb9jKjXRbqJD2Z95Qtg6fzc
OJUF8/XyPCKIgsP5plhxo9QnQ5SAM9P5lm8qzrsckIM0YvOddup6ZHq0MNjW
YipYoT3S/qruu0oiUXt/VBVeXtq0zi3vqsLoBU+QzlYzGISAloHyxe3DDjpH
8h5u7HqjdXonO6PrKhnWxjp8+Y08AbTEVgBuDKtbTo7P1kfqVP6NhJPTxxMb
hNwr0FFcV+2yiPxIaen+u14loo6g0TiO4UqEtUTswNlzMKgo9M9UeOEjp7Ek
65sBKnUlyBpu1Ixsx5+i/zG4KbXm28wMKSNAu6r/vvCOuItafQcybc4+SYDa
Pwlemxt5Ar7HQufii6y0BZ7xu0R21CP+vdLnV4xHzk2p4SvazIpahN0UkHjF
RpZtxVnyXAZr/R0gW/dFUVO34m7FJRBTr3v0kzvAFWE+ypEFdCF4tG2tPtkV
xk4yklhR7Ds8g7NrZKXXcCcus6CLxAQ8EglT8AgokR49srNqT0KpOX6ObsJ3
8S7PkugtIKAjkO9ikqiq0d0fncEOMWFwxPoR8UkYmQrJ8ajiZnSZFfONcuBO
SnuaUHWVdSItSvIjaoS2gN9axifBNqLlnCSLtQHvn5CKWl+jh1mZXtayxtHZ
jcqsyVYwrlVCbOi5trIwdZlMFxMO7N3fAWpvyRECUMLl8rXA2BTAQn9Q776h
3rivQrkGWVJ7O11wpLcTLywRXL1e2KkDXpreyYwRmETQGyspGLuiFA8sry/y
Hz9UlJvJHeh+3zjMq5l4m7bwe7R72/cDEm7fuRQkURBIu9JvUSHG96btAK3D
81JnvpxMYP0ze0gev1UiEbe0edcBZHt4SEHJ+KJZ+UyUtX7235I3xJPwwx4v
R5TN5VYu1L5tfRS4MfyuMoT5HEeU5jIt+J7C5RCFoS04ZeuBTrj70p9Jnn57
NIHgkM/v5URKqk3bJKX0Bj5rrjyAxZcFpVpiBbGziZAgQQDEDE57SaC0knNk
qKK16rukfGkKvgjFZjc2jjCh88k26JR1yROYyYDZaIiiMhtHplembJZJdpqX
Un53QmHCtc0cClc88e5+GoP3lny5K0T+SA7ZjW5wgDwvPkVatJAlmYK7oN9U
uWT/Tq1/+pG/naFvMsXpbD9XAV5nY42ITAVbJubYmEfxbxa4OAUKr3/PSW2s
go0bYehb+TbWKsQ01SNDC4nKQHkPj316IpHGvhEzX48jLcG2Q+etltt2HLra
4ZfOog1o+umNp+47rj0uQNfwqJhCOfBotN8z/atRp0PUC5vwopRKkBLNo3nm
xcX200ewIh1p68u8T333e0JGtaJDoqJky+c44BFF+QEGKCTkpYzYgBu7kx4/
F8O+CZ2QWxYFEd/4thqdrumjmkxnawLhVJLTHPWHeqFTnSswlm/i8npkY4uf
LKtsZkh77Bl0WBcKlvnQbBF0HrN0zRgD2RCXKhbLD5BrcI7MAlCOxiHnd9HQ
ewxW91S9vVqmcXJKh74zZgvTQk2UEY9u0icnOSPDTox1FTvNrUtJLp3VZe+L
wupIeXZrlFZG2W6Kn78GcHYwWxK5BrQ7dYkMrFHyKyUn6ENJdpEtAO0E+/pt
j0j8sqCtwwPJqlCB3f3utklmYmTTqZESR6CA4udX2RDDV0jPc3Ki/BBmI9SJ
vM65+e0BrdEEcTjNphx2YHgeYVTs72a43KrkF4w+ATENHk+DM28IWfI3PTES
4pwop9/oE4+XytTK6DnSfGOngzFN/DZWjQwUrAeWk0Ju5Uux62Y6QXAsYHB+
tId62YLW4J7FLXolTS8EcAPY1/TrI1jLCIX0v3BXVoV/G2x3HHlOtEKbk15q
78mvJ81wE1YZUqc81M66CYB8lmQ76buu/wHnC1ony8Ft/a/UbY1CJUKwG4+D
pRH9Nm1M9c7Q6N0Vqw8dE1PWMpGgbpYZfLLMtvZYdEUivKlPMZLrlEkes6Fw
z8HpUIBmwMFBur7fLCRwJ4q5qA9TmGHDFC21WCiuTfdQP5MaqIU+gVS5imjD
HF2G3t34r7aGWDUPptQ4pYFRYllWMF4uX5FlIJhC4tUIos4oOJttLUDl3FvD
eMRmrMrT5zSRSX7vzNhzbt4yPpFLdIm5ZQjFTVVxEUFW3ItH/zWArgYUbwL5
bW8mD9tmZFQ5mBaE4M8UwKO9zHu+SCEPRGICa8QaTDdYVGkYQAEEE0LO0I3b
T+kBXUg06OiQDWrqG//sMEAGpLP/7x3XIxDhDdEDgysjrCS3kBza6WKY9cjW
YyYIaWLZGRbdbUWMMG1/Lm7y6GDd70CJrT8iWeV/39AOp2jgJ711uhgyQzXS
cMCuUrEXrHUN3je3/ZBYd/xk45JAGlkuJfBk67ZeqpKmEQlfdKcUsqp/3dUv
ySXznLbjfsdO0wbbq0zaFT0LBr1XB0NJDr6rSCpyw5eJjfaPNjN6pWVj4dze
l9/M286WzP4XkvMmfMi4H3EeCCVchG7xFAyAakUizZ4TvmLzunJ3BYKuI/Ug
Fs0W7CB9zIYJB7ioFdhStCNMaD4nwNIAtCanSxmZ65r9fFJ24qJ1um+KZoUN
jYnphtccUb7iWd/ny0QcM/0BFncQRn/djiVt5f1LqLWQJlmxtCT3ct34ljza
AY1N1L5IF9ekeKOVpetfWf2ysW7tOyMwTTn/6nFrchmQeB0fEZfCHFhECKQ8
RYNAAl8Xk5oju6fLpWzZxYiRv8Z6R22F1ac4/gLVLyhlMGSwiPLH2kXX+H+v
ipkxkCJW5zwGElAt+MMzzm2k00BrOADFgoetScrkLIIBNXQ5Rzrabu4HDUev
n0mdn/wOvxahE1oNFFO+XJ6OATWLwmsVK12+Tx8V2Oed7T1J/Wra5UnIqzcq
SBM0huObesljSkWk9lMiKTxEBWJCLOBBA9frNm/b7u6AZWzxZPLaO02ilJfl
qHUQJl/Zw98rfvhbXHxfwtjvoR9C0ZhFffe7/jTbCreGm4SwQnzyKiQ9VLVY
Oh9izmk9Sig6NIPatP0FVQJwen6trycesBFhkhHCElj2nmUplIo1ZVjkfkrx
cH0aQsQLEJKf5eXxSRUykyJMPp67JBUHoA2j0qf9muOL8kE3F0d/3RzhsfZn
lrBIJTdojNC6GjOyFxX066UN80AXCfTs5I4aW7coJmGlYsFVxm8khUFkTx47
cxBvK0xJVcyHYjRTpesZnG0P1F4XEss3YID5MelepfIfjUE7PK0s2xRvCM8y
DdjMp9+OsZI1qYJke8TQy0WJCeeAdWwlGyYSxh4vzMk2oNx8ZbMWX4j1j+9q
3/0w2HlFm9BMQU2BeemgL2RJ71vkXy0r/xG8d0dSWgtZCHj+7zkfVNJP89TT
tsXtDLTtg3Qetuv11tJiZ/zi9kyYHQCro3gau0JPgcr/ASUct+fLUNkrcoLM
nWjxnUP4BfhU2N5G6nqtD4c4epqmqWkoJJvGkKSlOLMBRN0gU+SzLahZ6rNR
u1buN4zOAH2i/RHmQhshh+3U8PnrPL/YcxjkmtDOtSrakybZhL2MoSuX0cTT
SyIuHsMo83oo5nDW8QIYtMNuH9AQKi7J9HdYV0C7OLczbstaUnEz+NuHlP6/
Lqm/MWdsz+FjRAyiL+9+HzIsGq0r7paZcr1KYGvbcJ72ZAc9w5JJcfSnSXK3
VOIT/LfLU4QS5VeCrsMUAxBAV3furSOZZWF9GjCRb9VDrUg7ciGnoqi95//g
uJETTtGM8mnZ2EeGHFcXVqnglfY8UZNHgnT5VtG2EitOID1s9D263GPrPd9B
TyvmJx2ryr63VpYHyqAGndIK5hvwTGi5rUcP7Rl2DUg2kmzlRgO5BoIRNNWY
ZX/3221GYAUe1O2yk/Fse5UX6X/bbQwxKfJSNhCuHswqLmbQK9RNteipMEG9
chMLXJ265fpGx8r+SKRB6Fz7xiVQMzOPfIqBZMkUVLUr5l6ztpitUEVspGQ/
KLK8HAog9OIECkwC4g22plwRbEbaHxVZlzmA5Abac4pnWPwn4bnqmHhdQi8x
JqXCTGtnik+ngsm3KUvNo8Ltb1TKvpcJm/PvJfOF0/RkbL3RzRmssTMzNAPH
nmsKiFj2tjM95lIuy/IAx70LUXj9Ny7C00qUUiNvUPrreflUsVwMNPSxvhkC
gdrMD8kbIoW+tjIscgazHnpymk9f18H/nyL5TIov0nN0Tv4mPoSxryUk7TaV
N7ttbqQlUkwaq1865+tVZxAZOkvgtmEONNhX2nYnms7xjOk/+5vHcBbCeC6w
Xo7XYwIw0PTZ6KRc+yVifUXs5EA8Ru2E0yo/IW09CwTPGRvRnOrBYn1t7T9T
Tys/TU4JxHm0u9hTERjYifNMWZ5SI45HBmQWG4Xc5Y4PHwoU4Sf/1j8Eni8U
/8vmedD/9OyHbeTPCVnRIkfi1GnSi64qmZrcgJoy9lFzWGOhY/CYqJU6stCM
mO6sLKfqNfMlRGwNkEcFYBg29AZdBOHYeQ7ohveETV0xW83BzJ8YVqc/J7Ff
PGfI58pg1cfm4YCfNJUHti0UWE7tgkev7R4K8SmkHuYHI8Pdhk4pTqPaJeWK
rg1hS/rGXIEebuDg2YpnQe61XiXcFAiHKfJuX3bFvcEZU3JsiCP59skqznGW
XdT+hmpzmncPG1kxQouRp5O0CuLEflnZU0caWx6XVp3JJq0+HLrADe4sYMv5
jpypmS7yemWo4UIKbugAy0CwOE+8jAyQnRjgyxt5BD/Dw1oIZnAq4GFP7GcM
AcX0mc/5w8PB6xx+pWyo2Ih0STq8bI0cR1VFjQ4BqTVd94P5RuamHbGO2c00
XVjuj9pHna4rScnF+kP8UkVyI1f7ZtkoVy5BEoYZD9UKH5MhRJ8VqMpvxmFq
sL4SW1SVtS/PjUdCvuWkT4whUf5AxRwSC4s+jh2cPXIHHdmw+eGgALPNfOQV
GjRBINXCMA+1MZvt/UA2+magrwhi/Faczzloob9TmtAz7CzUFSIJR2Hdr/Fz
BECtR9TWFOykBfHVqhaDCWJilgVbF1W924MJ+fmzEqNFk/XVvVkIsN92VEIH
D2wEtHrZDy66y+I+6NOPns88Kqsotjd1DBfjGNmtddJBswvxBRMA/O5lIIe6
SS7z3PS/gJ4hyCt1xg/h7T1NN6vrArqtOwVUl7aMrarXJ8BsWg6nHEYWEJS1
2joGymU9AxdQEyXwKCFwJFKrAuJaQ7SB+opQGpfggV+GOIYsTIxJ0Lh03Sx1
dFOoap0sp2R+4C8zUT37ndwrIx5tWFEnS6lLLxj+B1R3qmLfkKp4rW8xLdBe
TfReXNHEKPbdDdUZb6ZCPB1RxsZEteVW+wGx7c2DKmLr9k5Wx94ryI/NOLxw
H2wGg9moTSns1BnJgxAnV5+x0RU5TxqnGZkoDKvPJd1RjaRVmDMJexqPOrLs
sLU5m4UwAOrOn41/ItUxxuLJ8mCwvyopkkzp2nL4exEBLwmOCZPTXfXfGDYV
kCk8P06iUmHVPGoKuOG4FGYW2JBf/dULPWmlApWClw503pXtHtgJp90X5QQx
YKFSdWzKJeegSP9kV5puTnRaaYCipvNG/sclSGO+oDWEXspLiAm+s6Nmo5aZ
0VSPHTvWXU2MmeptqvdzKfbDi+JnWCQUut6bWXRBNOrYLEIX4iu+IdS1exjx
17/vkGWS/km3me0ethgde0mhKWojctC0FKw5DKzC5pcPoHF8IxtHUsT+5pHZ
wPtdgScEpyp0N/25XwH93NKmlbhwYmOmNd/27f085vCrWBIzkUK6zPU5VyNU
xevJC5KI5Jg+R2urTudYGFttV/cpIZIWvnUkjsMQQtNnpSVFcMMa2tcfIoUF
TIHNgADnQCd9eQ3O9E3YIK6/D3UJoPW8MImm1Ek8bPCvRzY6NAiuCJsnLlS9
9l7UfohzrlRFWkM86CYBWm6EXgf8JUtCDE5kh7qJ2aARBM1ReriD5F1DAQtH
r6gzBTflnPxJGAw2wy4l45zRY5GyeWg45L8jGaIZbjxL82+ZIAdrWjVUD3n7
1K2AYyNxc4NnwrplPifR0tTuFGCkI7a64DnmcbqSJjdyY+5/PqUhmH2Vfosr
NiblqVXl6TTeTPUbHxgXrxkecy3X6n108VwXnEgTTVpI1y4Rgc1/lrnTBta7
GBC8qNJi8wJqrpoeh9HNUfdWIVstFbAUomJ1xHlzfBvlVzMUhCn6IdWTsHg9
CV48iXE2sfr/h1oX9bx3PLty+diEmynOIfRd6Vo5Aj9gGZwXqPvj9geDKr7Y
8vGarPospCVJBxpILCxKkWv2/772zB6aKuN++EWbIogyqCfXoH7i6WatQ9IH
ODXBg7FIzWkQ6W/EOuj043KG0hCa9Njybp4ASmQr4sY3sbcvvGuDNooteDev
NetFRAKxO7Bh1gyzpLJVhdNS3mj+MECwi92WrJ+5i76GhLKbmgac6vJJieUp
RcRBxgG61JiDtVlUqnhBb7lZ3uD66+p5mU1wUyQi30Uk+qrbH47KQ5GpVeXH
+NmAgvA5k9E1xZbfIEtb0oRIRH08twHbDfP7KI0BJA7cQyBGnP52mULY97Jn
nLj1oQrHht//NHU37JU2pGl47sD7+BlDYm2cZisLuneVoztewaLPqwGroDuJ
Ta0X7rzM+FLDu6T8vJZMSHt+7sMkLTy7A7K50DloEMTEZg8KVg3EiXnwkw2l
CVnPkt+tKM8qZgh5ySGeT5xrtqCoBHtYuyVqOq8d0WzwQsTZgjKLmBS0EL1o
BIVkpmQJ46/ROdZpyuGFz7W8BmJiaeUv0Kzing7D2hEfOxxF8P8cJm0uNE3M
NZ3p9ohSU50cH7aXY94mqr+q76Qv1KQ09XFzfj7fS2s913DdggLe+y+XCWcN
dcqiGhbWi/m53xSQrImO8xsm/p32/xlOdvxw/QKw9UZdzxuzfRW7aOhtBWdr
mcOrEgxz4kaBeWCYaqsebaBM5Oj4I8o2F6/4Eg9oQvZic+hoapp/MNFO5XqX
UyuRRTQKk9DJpd/dhKKMRl7tnPZxhtsFVv39Ax7RGlTnX0fnqdWIfLXpopFN
1wjwwnVgMNOm2rqw9JBY1JZl2cIxfgEM0QG8isHfK1BRzEVRK1k1c+hHkU8L
8QDyrYPQGa4EtQJmsfzWPqnhBZhqXN4pkyS+B1Z6EM3biWXqrKb6KWuTXTX5
bsQctNXBGbcDuGqkmCKQVstxV04K2y0/LyJe7LH+8xI81jxAyKV6lJSyMRiQ
4taffxeDqPyqbnwFlE8e8Kkv+016oWkR7zHFL0tPUbGloAR0YI8enoLtOmVX
t2kYVibVEzWjwyqZFKEmciEMIOpRNhrKb8Ss7NIWUAoK7poV6+ARHycmuiPD
ELxaGlKFSfszNbsIHXxJo4yxFlLiP2c7kLwZZ4EaxspRrpyGCzXvNtOX4z2t
jkiYdWBL5SsGZ7hdNC6jfj9+yP8xR1lHidSZQKhI/Dze6orybroRzztPrxfF
3kWkNQLEECEOSuj+8C9+H2LzTlavXgQ/xN3hh9vUjEfJgeIWbvPSkmhpqKx/
mUknMQmJzwtyAvMfbrpj97d0Q9gIoF/75dpx3M9Kxh30VaUdexoW69Q5Y/ew
N1hn+4eEkpFzFU6aYrFKnSddYsvE2JFkaV+MR/5towZn+TnHP6UYjeA3vuwR
Ku7U8n+7nuh66vx9tvH3iPQYn5t2cTtuWWJiDrP1DE1wsvlZZ3aqdiU5PC7Q
9SsMuLYuRIWicD2+O0RsOpwnFQOTA6weQ9Ik55o3PIM1X0IKBELyiuvj1QHQ
TBvwElaW/801Zh3vyA7SH09kY//Fo08UaElk5hneczUhKXDmztj4mZbb7sV0
ntBL2Mt/sO5kMgMKY29Q7RmIzzaEyrYwn9beup0ehVRcnrMSkGGgU4c+gTAm
8b4itEN+F0XS06j8zVywa95/FRyvEMD1UzxP+zMu9ZYoREkchidjvxzflZSM
WLmBxkc2zcv7atf3bFa2C4PnMVzPjE5aEzK2T9oFImMyZo1xwbH7zOB1YWGc
VmWLh26p4m/31pbZ11UdBMkkjgMotNETCpZvZkc8uaKPH/NxDdTXiLP/ZvbF
iypaoqH/F4eokfelmNJD+kxy4XxkwxhBy9SSLKVr7pFCr3UZXdkiF15saJOt
4hQq6f/uQiMVTztOa6cEzubcbNUe0dNA5PwpG0CqXp5NmqA9KGUPTkdVwqI4
htikFtGtkv1PMPyEt3f3/7eYOlvACRdzDrqmB2NhADnRLbtehypT1u7wF82+
ZCQenyPNmzdhOZBwojMFtFfmITHadOiO2wChyE8XWBOyKcTYrQxoO/PoEyPc
ODsN5bLTWnTHZex9XKGAG0onj6hE3YYTZyWg/M+hv2ZIpwXFYQtsUHdIfn5Q
heh7fLLfp/NPkznase2r4K6e7Y3pJZaJw5nQ7veMw8sXPhBEr8cp1BtXipDl
NjFHyxiE3uV736Yxb+axXa1RFjCUzB3luaGMlfUZN6tIl2RqEEgH8SntJtRd
Lrb5bcqO9jAETI80S3J0rJJSB3RphUgrsyCJ+bRRQJSKH6jkUTL+nL8eUmv7
Qs4jUmXpfzGSZw39am6fZJdRsu+k0EjD+tjQjSeWFjPWFSy6GsU48utzMQmC
ez/Wqa8I55ZX2B7XkG3N/0fUYdARYPEcFtKSBNUkJ9Sr4647UBdvsdXRCs3v
CGZ/h8TzUYLKdH3nHXyCRULqn2CH375bbU22bVuAKEaMnVGnnMrFf6KzPGB7
HTTFqzfih6ISD82XS+YoA9h5SdwQXab3/FimrHbgQ7DSNoyaAuLoX9Keo7A6
LK7RGBMNQ3SIn/NV06WqUNP6dk6nOf04KkKAbX62l+0uqIhGGU8pogI+k3/7
Oj+c57b21vFHnWJ+hPssXe1TTxtKyBFvcRjcVaYarkPP/rkZjcZx9y5BzJj9
qcACE8nZpR6Brrsg4LJO7NqcUyTXdlSkE6+rlJY6WQnbFX0wUQf/efB6etcN
t87Ew8XTx0mlA+LmyfiWcS6jYiQM5K8UXNwecjrWnyZr0tq/ktKwiCHTtLdW
nMVA+3gg/SiKz33dbjoACD7yCybkUS0lJ8ouP6T05tQLKWKConxJDZGAJhR/
wpgj6oVDGLKfSCHbRJSfRzDl0/bB/eoqbqJfN3xK6rAgoB3t84fGntjeE7YX
UOdcFjOSOTy6U7TGdyUfp90607ylGO198QB/0fLkKSYt/sHSunu3TWnIobC9
7d+wXGpDyehvxe6iYkX5IGIFyRqNR7i5U8CPsb9xOud+hTwh6Pg1WNfw3ymi
DsPA/HxE7fovQfmZYG+KkoMw8Z81ocpTWLoFG5nJhprRbtAjW5ZOGuuMrvhn
CuWaGY5mdauq9Jw9cBOUPWMPiHe2/RhNSPreP1LkVC2/L7qRrcNP17Y1Z4eL
xMlnEPIr7JgWlsKxveII83oeE9Th3hV8v/pLJRCxuZHBbHVu5XwataPSWuUg
qNxPWZOzPvBoFKIlapnaIlSKbXL7ezoMdWQS9eJVMFQX4Jxshoqb53kzclap
yFXSpFmb6rbPiglATgJ1dPChmk3P0CWhizJG+ZHlL+mp6opT6NAWpaazJYcF
WpCWau6KoQvLwE0x1/yZJ78XPkZbhkQVFaRrSjGpV0CVmKs6axFwtGAqIdQZ
u8br2RmV3i90iqoKISdSfM5ws3KRTZezM2Qj98qIbNaC/qGTBQrgbWRVZpQS
pD53rDknIKBkXjY7TL2MXmffmdGelIisUGAgFMxX5BLF/lQWYioEKQ3/1SsV
FZyx8bXq9rfkcQIlQb1YOtaF4d2ZxFVAX/cbV8Dalvxk1hiST4MbEtj4oxQg
uO4vvOsvrCrcNzx1mK4dVvX8hJGvy9A8CHYH4zRt3GkxpCBvCZNUWLHlOPTL
HoSNDZ1Y6P1WN90BCkQ+ZW3fNWn6GWgophvtZ6qXB7Q08JkINVgPW9+0QYPD
zDvALoEy+THvx2fAaRCDL/DH0Bt0rllefjqKXkIDb/8lO86GkasJLk9Q5UkA
gGpal29NeiEpukDt3Trm9NuVD0aDm8hPt9uFm0AI7dyE8NMTuGfj5GbWfW/n
QlaBu/ikqM8pK1zr9TiFmNpFckpenIJNfcPJEP79grIHmVB8KSrI5HaMobAq
HQMJuDZbIzjreE1AovBgpAhEMaCthwYNdlXeVGYIE4tn/OM8ItmL54T1WJpp
1VzrnsDLt0FJ8k8lJPOwOhKeWUH+uFqqgAW7o7nS/W/7now5XtmA7UwMMG3h
fHrmHFJD4+e2gyPgE/MOJhsBFtKo9X2iIOGiLZKweKPXrLXehXaWJh0F2l2H
CKWXjqxeA+yzJrB8A8rkEfu0wbMJ0pI9GyWgT1SakXISKP0w8oY6kFEF6Wm7
jLYyAaPgt91O9ya7OQ7PlAFzXLGl16MLvTcOtHJMdbRDBZ/y6eoOfu3WTDHv
5TbGJ70ORuXCNrI/GR2CY1TDpv0wrb6RiH5iaI1P44qi9tIhmWuxMUzPKl5d
2KuQSlWE6zt9Mkinm3FF7SfuMXbrJGu7C8iwQCNW3bKICo94+hV412ZeErX0
uXgZ3sJzU5bCWhjcKPKmpYrfi/sPErUZ2MzOVV7R2Fa5seCgPm0ZLrNd3kIt
C8CeSVvKe+6S11SgoVrq6vedpHZGNC9v5XRkwv0JqQUXR1uOD0gQ0kN1DlPX
+d8l+9iJ48tmHNwBXpoAE5OJh/S5x3SEeHr1sYLais09IThHGqYIwZV6kBCh
CBz6tG3s3gFLucPNX4YMYV2HzGejyhYRVpgxD3W26HVia6si84h+vY2TfDLy
No5aaQzeDLai8fd07hBO7Pr3G/AWAYH3LcnR5NLljd6bBD6BE/HA+N2+ofer
aN3hhS1qKF5ilLKWrXHRVREgi5+VGXTb2+pPXCYy5NFOdLHLdXmEBtPe0LfE
phl+7cCXbU2usRwAeAk9MR/Q6eKvCKvhOmoDUkVH3K3ZLwHmjuWjoO0uqECJ
na/k312NrhOJMlgQ1rO2Fkb7qZmRoQ+b2Z6JFswSfmp2UMbJ2tINCsb92d7k
UN3ZetTiQja3CkQgdJZMolJa19uovQiRH2+nk2cQsErVNeLraydCeoJ0SP5G
QrYNS8Tq9U7GXCMf5tPlGY2Y6DsZkL7okWqbJ3dqhsM3xPq0bGpoMopjEN3K
sDomdu13mUd/ElPznoRRhbw08oICOFYVpwUT10z2tg8D5so9KbzBe6pqFsGd
JJ3N2ocZWxxFJiCZjwRrptdjn3YLIqXkSKJS39ZERHmmSJl5y854ezQUjXjw
6ny0p2i1UncMDW5++K/02PhfftlrNrxUaq17hPWWtNsmR+vYjmY27zTI4Mwe
X6WuJBaXGlbAGLqMPODVyZs2bCGvUMan9mO3wAtzmpkqC+L1RzwnOxH6cAuT
rR+Dt3Uuplvcjbam9JuKE7Mp62lkWTC6ELxNy1RKud3lMh/KMlsq2pEaDSGL
mERU0OpxFolWRi/3Vql6GriRwVjZA68MXQ31JvE3Snoum/JDx4aGLQE7UYhL
BPM0gXzHJRnzjN1Z38IqaceKHjJtZWXjEoqS4IFk2h0xjptwUfdX81G6z8bQ
rTHkG/EuSd/jMobfQl6j4i5/92mNjZ6BCdJU9ODyuYnpkU44RdPscZQ/TvlJ
o174ellKwVv4EFetPf63QTdtPQlJS18lpcfc2bMuBtAuj/kfooz9p8RiMQvg
X5T2MV4NBR4AXe7nh9AuVg/VvLlRkZc4II1lGG/xkqv9yRdXJgyp08kPZb8p
xxa0QSbw3rpdFrPhIuxs9P2jxVY/0KorX+zpXmiGBAbutvD+XVqK7Uae0m4/
orwoKzMbWLAbXq491IXK3ZbJ1dG9BO1VTcjinVTWvB2NKq2Cbpx67VO//f6u
h3T0oy9/l/jVA6WDFsJ+GGhqzaMLzLz2kvlyPCcg4MksfRNt9NMOusoy2WjH
GOdGTAvFw88n3TUETCjevflHNswz+I89gP1X9C+L2ZSOVMwWZL/jCe8Z34/h
UAoiJwz+Pd2uu1Bh8cQKVaHNkGgGD5vewcttXzhE7U8aNKq8rOs0VpUIjEzv
P7oJ8DmJUg08LKXl3tIs3d05se15jO/SCS+JhrugsV4A85s6Nzbqrh1RkGB9
njTbByG/bh1tPIPHXPuXvAEeufgviUVUW/Nc6KIZZ5DVjg5RXR82fRU4+Z8Z
h4vMQ1WDG9ATIz4sphTAN51BZDYnC3uNggAFE+DDbFHMxSN/OFvK2e6wipmb
0j7dc3lsh/c1efpjrXZcxsxmegIjObbCw0u0NJTn6TRWRfRlcOE/vzWfZtyv
g6FUOA9CEeYIFkAm4rIasTCPzjJ2VvC1zZw78TLD9m6LL7R3irI3HhUC8Su0
XqRQtjMA46wDIZSo8qpu6PFJlwVEE+CerhZyMdIBbBOG03YPZJxctxqezeOB
znkDAXvohqY/Ei11biXTyPFka2kN+dl+jENbGC0iNF2m8ExYlXGZif2hJqo/
vEpVTFPD8cwBlGvtpCOa/iSAAYrk8oZQ8UuIemL7XiYCQAeQo5XgDD6mj4h8
Q23C3lcvPZz0o7bHVy/PU77TamekAw+2f54vr8apaHtShSsTf8lf80tJ8C8+
V/BH5fbRIHdAHNuhboclxNAzBhq+WOkhWYYWkyEOBHYVlI4vewKRw7OuNs4q
reg+ZqGnLrHmXX2ft7D1HZNdPX+2dyrrR+cZXOXiyt0PuazHjnEt2Ql/oZ8p
mWo5FgEXqFxkiD/ZFrYWUcXCkRDdlrKRyk5+Ny8+58nMW63Qoy/7mGbqWLib
ypGy0pam5lnYE8PQuf0OghsMEB9UBYt6tAZnbSgA9GVB+yG806tDL7XIBHhD
ZUrsvbks/4JhmwPp875fRk8U+EMwcQvyRRbWSO+BWVTernWPWzZ9RXh9HUaC
0pWXPzQ2Q7ac0EN/aBzFiUzpJQNBW9e2gBidGpLJZaweBgOTNa65c+dgQ59j
11SR0m4J6NUpsuhuL/zFvCIVA8kRdig7r9K1Wpjg1rkzQf0Kqb0UXQL8TFUy
yTKV4mCllgAHi3EdT0AveOa1/iNLTjjfezjgH66RRnA+5z1qOhcb2S8exjQS
EyNVo3WAcQsDdnpgz2xTv+hxrQIkhlzAGvQSAS7RVPhyJTafw8jCmvys3O1R
2XozBm0BIlEuWwPEdAbj0PSfgEpLfDWhiYh5tby3IXLWjeIlxvlVVHVGb67U
NDrZedoaH5+SwdHLRbvpLRH6fG//UbOZJ/+jOCfhMYkhjrMG7zCiidFN9qq9
H6fmmJy+Z7ovm6aevC1rGEDslyOza1Q3N99o+SD/WyP5ykPBDY9FavKYWbON
yfyFQHo/cV/3vdHtTwDA1Nq/9GFOOwLmQd8RIELMvGLTet/EepzCqjQ/jV8P
yJUkpP2Dfnw8Gy55Uw68Zx2GzRpLflYPm7z38KsmT2i7pvHzNRQYqcm9mvTq
ToNd/GGMLkio+WO15vzsBpPZJ3sjN8tH65flXMTb+a545l41rYJ9LE7mmNGY
NEtbA8hFJMWsUNyXSwpL5lz1aBhE39EBamrHHJjhRi8eC94Yb5fDPN0PXB/v
rxneJmFjlND5jQTtW8AODrPTJ/uo6VY5Xko0nISDu41B+ReUcKKO8v0QG/A8
fZjm6jVs/88QoBTQ0PD2HL+TOYxcjGY4CJCEKIaX5EH3qKNzHHnmj9lnVudm
C7xmTcp3vbJ9MNHlHkCtPlOaPN8+LApN3J+jO8dAWkEYTFIWoq6EjXDR96YZ
86zeYAs/Lndm2iociAb+VuXrlNTPgs0Qci1ZoWguGuJD3vO7Bl/RCUJbz1LK
6610iMMmWZnz8FmziKYHn/ToIvIoDO7dtXUCoPLuijgRZVEvkSEFNerHKlPn
RjEkUuFc/JhciNU7a/Qb/6ApXwepr7d8arHKRaQOc21Zm0826/ez6/93UBPJ
xK9lBBSqSYgXLD/B64VUggd5fIRu60PSlfAMU86JZEGGrK4xKUHKYxEpjy41
S37OSUfucRzq6C8hef2ZsNLsduoD77JwJBpJIVmfdOyudMFiKU8jYcep1Cg1
sUjSxoh+NiUMuSty+5VpoCTWeGLOeG6MPhKOasD6CmovK+9Ilbyamsw4i6TB
+Wx3g9rzA0kjTf/9/gCDX2fwpCsg4Juhr6PpzOCd+FG2AwkQIpWa90P1vC38
UuTkiqu+YgKo9j+39tmE5Q2t7MfrGdOYe5Z7b3cLpZMpXI2Z2w1cbdiEStOk
RHle/KiQqwMLn3TX1qRo8Zb/0RfSsURwZnKvFqoizblfHp+6p2DIFIfo8FCh
bOcigAEY4OAhe266Bza+KMDyHgJ84p3/MRofItWj7GtCpTeouZsrtzWFqYsU
eGgZ2oTTCVmSaFBjMCcXyXM6YroJDZWCRPnuokdpUiL6gz58uXWt63xeIe3/
aZ7JGUVY/Ll98gWa5NhI/c3a9IKHNY+KNWt9533p+Z4yGs3jjgrVBktsoI1Y
JRAbM39fCEsO+fc1nABvj4BAFrKUDd6Bp2CSENVVNhVkWyA/JuwlyoJr+8Zh
iYUtIjLVjU1v1T4EHcGOOJsC+D9DDFs7z/edeQ5hevgllpSBxB0PKQFyiWe4
vofS0UxNYgcj4ULjnvNqqw/GAYfMKIgFItMgWRS0u/WU7UHBYR0ThKPmOago
988e3KsoLsZV1T16Vv7NWKBoQaG5BTT/ZvylelRLyXHuK9nVW012AJ+6UkDD
DJvqqJkO4fCzN7BmYRE8eNs359I8YV9hNNl4MOYaCQvFuiTdNiom0140HVWI
aHnObrwAEQI5m/gxpnBZz0xYTJY4tAie0iGrosYSYhFeQN5cAv5WktTj+Tfz
y2iQDJ0uTfWSDAoBMvAiaZHlcbp6JHcTpswKLtCqLae9umUoZ8EoaDGtW/lW
jhhXxwT+mYU9S2B2EDtsq+5b1BhPDtbZizDP6Hs8KKeF+aqAJNXMitmoCq/c
2xymdziIVY9JPtAKgiyEW7lX41bUn38nP7RG37iaWzKzJ6B2936ad0us9OPT
7/nNJTOfSxGhersjJ9KvrnhhhMSrT/jfR/gShLMg7RzcnAFtr9ZqHVlcCLc9
S/dZrjf7NHN6iM9UIPza983CzHfHT8lsljvjIEKAHxBzAujPC3D2A7v5XwBJ
+QgQP3unnA3dlDhByfBZ0AYN6k74xRQWFWeEGVmlKLZZXVvsxbxbARsn1TI/
4fupPYzCXqtaDK2mCAz+duZHNUtg3EXwAFqDMNdOa/rWex8dphj2uPNePjJK
MoTE4YYx0PUFT2EHyU3Twznd0sOutogUa+Jm4yz6jKxSH988/O8ovLHce4Pd
c1Xb0seTOrl+6JHIKsz2MeuFKDa1T/Wep6jqkrERkoUOXp5zLCF9oI8CVw30
aJM3ob4XXILeMQqfJfVFJbus6IBCshuSoSfeXxYkeVuqdTuh4I2KEpMI6otg
/Y/U8Rhm/ohD8oSj2l47ea6LcgB6qxp2MbbdwtKQZ8qacyRUObzqQsqsC4tv
8zYDuZygb6DILoV8lvjQUGWILkYKA4YLpsTWeHHAPwghmOs4GZwcBxtkNf5U
nqoCYEl3bJXUX4wfkdbGIFCg61ft3ylLFTwuD3oUAvBpZVfgUcy3xziLGNuU
MburVGLJCT/6aY5P5A+zKaKpDzlMbEhEH42kBQM9riLVUuoUFNybZYaNzsXR
NBV/Gq6S8Z37MZ8LMnbqxm/J382Y1tEJZsdc7TMJjZihPGOlyWxw6ZpkxIc3
twEKOfem3iUcAEh/3ZAy42LXDac7R5Kw/7Gthu7iQU9L7S4Db3Ib+CHLm1Pg
RQfV/ifAOQx/ay0G7mcXvalmiTPcZrRdH+cqJl4dtKPieZ7qzxwB+JcFkIPF
AriAUnbnyfWDap7NhrEbtfMFJFromrcXcuy19aLmIMiwDqsThn2TYEZxeurh
3uu9aBsY899JTL/8xn7Hmq1Yg3gmSt5zOct5bFaAYMI2nlY8NZvdNUCss7iR
ppeJQJlvyzKwX4bF5ZtMi+z8ovI9jxzjaQU0/KdmHzDCLaWu5lHHVEWuXOjj
Rlpv5+X+w8LAJmi3+I/DFdsR1wImbfAWgMfVuFNWgzZ3UUSIqICRUc1i3/lY
AXTy1BR51xitHXirT06EOzqt/ujI3/PZTiOj6pNaOfhp53RK22Oje5jaP/AH
ziMU+mn1xxEI0Gha04+CgIenDGtAa4ItsoirKD9gSJdjp4OnKrn1z3FQJeJp
Hp4CIeUBoWJeK3mDRiI1/gpeGOQ0TdkdYpsC2XpwOnxJaf5/9x7Em8Kb1gNu
5CpzsZ1mYz69YbOZTsB5/Hg9qhumbA5h798DLGAcfQnbsvkiiknJ1IHkCVpL
laBmuS497fHJyMv0LcdOCXbXjEEgxnpnyAZprQ75pBO/o8YkTNyINSf97DMe
nDB+TKEwIqzL52S/WV72ea5Pp44wdNkEFYXis7CWr4DOaQPPHUcrwrgtC/M1
pDvocxAre/OnPKiMBOkd8YKN5dWCGBz5zKHQGxby4FAzT1P5pPZh6Ubhbfjw
jA6wPHvcZGTenBwi3vKc6L5n+IgDu0lugkmbjN+4FOADMcEsVjtf2jKq6PW2
EYGZOBugimOtSQRgG2AWIq6fWodf3J0Qbb6UGzZdUgLq8t5ovb1PywFs6gOF
R3O/cTWuK0UIbc572IMBwmffIZjE6cGVuN1tX8FHuqxkcLVmHRCZwxOmnsCA
tSbpOKVNsmQUWkqfnqJdQjQ+pqnjbQkkHZ/jIGfvmaKxeqDKPUF3I6bKxcUV
f+9Yh90TdhOrYjz5XfOoS/diiJGVGCRM/hkTqEWmIvGyG6xe/hi8VpDtUZt6
Hx1fn/ChaJ+TIWDI7h+23B/oVozdaMgVKvUBzExQqf+VPpUyBYJSjtU2OOrL
VXV9ZaSWDB6hJivzBOLVKpjPXq0WgihNE8acWg9gOadYHfLQz+VkfwulTjun
QJ40i1sezqHk/n8XzBlwV12Hn+/m8xi0eeQQYyZT9mGYkazQQkp5H51vqtpx
37wAwsRC00kcm1DbRi/RGLjdpbaYkoWYBClMu2r6F4dOOxcKTBwF3Xrf3C55
w3j8s7/MMeiOU4oFO0vOqQdR2R7vhtFCy2oMPqMPaXApuThxJKhAU7nh2F0g
5p/HC2J22aevTRBMkpIhQpwpIvW1FtVVO5RR/LvIKYQXcCNgdMiQSemXZWBL
o0F/uVowuiRWPZPHyrXp2YeoVT5lhWD26DLEVuoJRDJMHp60h8THNEC/GSw3
MyCPbJVEnkkV/qZ6dqGrywC4UCxAQeyiebokZBYeE8aJYYNOT7aZEjSy+3kW
Sip8J/CR6Q1pX4Cvr6v7tvh3+jnLd41CBgGGJg+rI2Aju8DFOD/W453f8lfA
sODQ83WBqu9KfWRPkPn+mV5f+iyBjMBBZysKE/R9SwPvKzFhXHV+EKWGEPBF
2eQZyMnqMdOkU8epCMYVHJxFx8a9/2yzZaAD/VCqgPz6k6pH3au6AvxcXcjb
lniwjlu6JLfBdONE9RXlTPxJ9UNjlf6t8esGxK5eLN+UiDCj4ppouVXkIOAh
f0FAFD78XKELZfOJjgqZHR2VDIpFzwL+QRGSwdvx8KmqxW+9Qf6GnMqlGWnJ
Nz1HM2gBvrewaktGFIZjkKzGP1P+DXYnh09gOfyti7h24mkrD/m//HtAOr9N
9sEWxVHVIvGMdbnCOVaEHs9bvppbl+/4e3qDBE6p81ioUq+B4XMyVg4bzJKp
yshfB9umzdPiMUe8hneAqWGNyp9neHogyORPN0MjwdnpBC/3CuSBmNQA2vzJ
VxiDGqe6wRfNQ87/fFY/68jflaW4JmRh03InMgSCK8Z86S6dB0NE1CiDfesZ
0Zq0HaRdM1GcXw2ZYpSkYLTYMd+181y6ymH7lCkWk0Kq5jpa1eOdM+unU0Ev
Bv6UppW491IeEWGXEj8LnjN+QbfbJ4iJLeq8OXKJbSP1SewEKH/6/ZY9Dj4s
GeIhmRc6ELpy7leBqboTgFG/yk2S3fwhS+IVoFU1i18ySyOXhy/qgjBzl3Z+
cmb1xfyfNITjMHWDK1IU/bF1rXzgVWJiYw5p0zmwDTTfdq0GtZ8sNIV8/a0K
pmin0P6clvxhRTrKls0LozzUF+SEhShcvtdJIOWxX0nwuTUEEUyhw0awfzp4
TFM0cmUDBIGkHa/Bpp72pCAKYk4EoWVyBDGzKLXjD1dKxFKg7a+Mrvl922Jh
Sn0/kxMBZx/46Gc7EVwMN6N6nbMQv1yuxketGVeNTYNBPhCxFoqnceHTEq82
/U/f3ArUjcAnduQ5k012EGCQhYPpImcUsGk4BPc4UdHr07dfYu7kTwhlJyQx
Aym/x1u6WBswV4fql94YIQHuwE1APJxJd/L1uIXoj2R1ru2m3ksI7lx07a+7
xgQfxZSxQDoKX960jihI3ws+WhCliYzlEi9o2D2CbfyB/4UKupFPp9SKxWGE
KLyHbu9juuisovcWz0lC31NpD005At7P1vVtQxNJroc/NYuknqC/4n8GNdMA
QaeVzzLO1H1HJBAXJU7S3lJfNTyraOHD8MOES6pmCCUlm2LBZolPtDTmENml
Vbhx/qLEQJzxGblVJ9qBiawP6yS5TK/YmVP571iPPsrAU4U7YyRyji+JqTmb
VmIFGMNxHz/O2Qksq1S00SgixQWzL33yHsLyCtQY7IwOHuQsChVzMoyIp5qj
JjeI0hCOcUPN/AvE4ubucH6kAvG3BQBlwSIJTNslfGl5D2yuhGqHSGHu2oqC
E2k3AAyIm6aPAv2ljYpQk0PZqH62vt96AxbxwjAcvFuCmgLLthjWsJ18UFnW
qQbYz6X4OuyevDYX5BdDJEdv3cOWN0zufVrIOV3tlZ8tMLe9+f53FtUiIPIE
qXmTmN5HrSw2q2tAOA/hD/kMmC1ZrbxPS9berldp6gKxFkwHvWAelLq0097M
ZcIc9iOPZrIxxs9EpSUk1b6T/IxmIPu15XxMnp05Hzh5BDxVbGkPbSZyQlXh
d6T/FV1FRkyu6QUAxKvTbM+0vxOt9DlejK5G+8moEsZbd+kx7KcTqxqyHxOm
Ezy37mQ5Q4RsafB/uj4hKNp18Kph1X8uJMJX088bpYRZrzLFVkNvK1dw9ctp
xOzmdBHdLvFxnQO8UTmYqtyvDYggUcXYadettWv2eg1w2o075FIfV7bukQCF
Ae6qSbSFo2E/DIQhe4irJNtQ7Wh6hv2+F3LHfKhCrIhaIj/5UeE5zy6ffDud
1NMXkPMhobmJqltZWK7+fNcxQ8Ov6Vo97vDBPxf3t4kfHh56m9A9JY0sy/DX
LjEBzihVuCoGzVPQIsCk8ah4Eidqw3u7+06SNoDwmJBlZS0JnsfNhLBsjN4+
INAP0Qz9D33MEMZE7kvd89jqghuGqsKF1tS5gE2mAb0kmH9UcCszfJBiPF7t
gV2IKMG/Z1rv+YrTf9jIWmLsYTDU6Kj7XjS+zROwLjk5aAkE/AmdF4inZz8S
QisxSpgzK+0oxJISWtuvDrZGA767bWET69peoTy4aRbiGcRUj9v2WJ//aKxr
oVhQX0wv9GftIVdT01syma38R4+zAX2kbdEpp49ELzuvSyJOCqHVkR8VUm7W
A6pqp9he/m0t3Nd4pWqzPvHqVZ+TdTV9fG/lOtQZiAiXRgPQoJmt/xvJ5iST
k1Xd5/R2vIm/xA8IfFLr9U/TAFhCgzXgHSwcTl0b25rwAKPgzmH5EAtTcqE1
4iVQmpLC5jmVt5f7avkT78dMWH4iu27vv/1aXyBjU4c6SoWV43jxuNiensjk
AWLFELuq5dmwJJiA6kgpNotkO7YAVV9+NYRWxJnw+W/SIyRcDD+CafaCSHUP
eqMimYm5/lQRg9h5EJHfeqClasbg4EtbXxh50fKgQYVUCAGI1rAiJ8FJNFzw
j5yxr6mZ4CEUSnWSKD76AqjI9dG7BKLCar5ItKKRtIFZ0QKcTyv6f4OXO1JP
S3q46vCOw3IbJLW5UEiSikKb9nrZQYBypkPfJMRB3M0b6F+JK8Yj0KJ1v0PH
GDU+tOeuo5OzIHASA0ItDotVp5W0mtIvesh9o1yKykVW6HgkVUs5zJd/3fjO
Aqbt9dMu5V1Wf/2fOmjxKr6w9LgFljsgd92eHf1WrOh6MwZGjsFTAGEVQiO7
eEn+f8n6qa2lBtfsHhDFd4j9WJLf3RTbfoJetFR+hZVUXWUsRvby6yB277dA
Xd1rIPT8rtPP5JjPKqLM0agtpzzs4Mm2iFHXT5dJ8fWVuwocIzDwPYDCEHHS
mj68TIIPG24js3k1/g9gxMffOvwIAW2eAll9hOF9lb/ctlLTFAtS85rxPM0m
NFFidQDlSneD8O9wIZeExtC2CQDLO6PMbtMCKSkNRMhiFulEUyInL/4yM74s
2uwgDWrN1/RGzPm9OAx0K/sJ9vDSfkcuk7y7vSH6v/tOVjA/Mg4tqgdzZNfg
R00f2gAaqyqJCPtCbQ85frPezG8YEpcX0QbLRthDhW6zddL+gCPNPs0THG1I
W+G30XK9rvlY8d74MfBjS8Rk8oPzzH+S0AKDwLGPGQZGjvES++NtTW4t8rRd
x7BI4RSEeSAUPkkDW5PshtLohWWu9GDD1so5Vf1ye1B5n5dSUfV6cANQWA+W
FifKJ+fiWf5/aYbKGcnmGF2j31Th/Kdob2D4Z3rApfCNPD9JoeBBjo+0Yh9V
JgcYHCSXaGpotrnOFLV6PDeWt8yQ1fVftQjUelgA0R82z7buYn8kocSVpJNC
+lVesqCi7qKEZYyPOYZZbQWRzRzqd0ywCInkwUGQyNErrCwSE6eeZszVSxfd
bHnJ3jDtfCp1ipCKIUv7wMJOth4Xid2zCOPeE0e/NVSZaII/62BV4ewWa+1s
iUqeiK2xGB7PCBmVF+UmtqHEUa5+mTx52EJt8GXk/mq0sXDOW6GDkgzSKhbX
7aYJnxs5JewBUNAUJR2HpgSbQFIvsl2KoJIxL0jjoK97hBEeFVSfJhmAZTeB
VuLzSCCTw99ocxcogMrG0R4uSGSizMAopLjbJ0p3UjXS8dmA7pziJNcHQfq2
xTTM+nM1xGZJaJnoZzZozbTU3RDzGQuZUzznwJpGTGonfzAWx2A9j3K4Gwyn
3BE06I9Y5SKz+f/qzp3ZfPuR0lC3Xyq1HmyEBS/BR6JcimfaXsb6PU9d1/ke
RWMg3E1+ftxE4MieFvlj0clAJaZw76+k8SuWJ3yzFEJxgLtFWHW2CRoeHFVy
A6cu/kD6GMvajQtyqw4FJu2RlneKWbdasxwr3hn84TwgkSKL4IfkCJ34GvaM
yWYgnJiQ1W2UPzEjNW8bLuKrIU+EIu+IX7AlkSIfxYJKIHVRfJ8ysNv+SxyI
I81Ia4oLMVpbkZzFMTYeqQvfHgsfCC/hc6crtKCjeS8LZa9YYl4c+EJg/CHB
Zr2Rlp0JqJjNRQ7TD5Fwur8skcM3JRV0wxMdLLKs0r/dXiRDfe0uQmdYuLtZ
uTwbEJo8aEgB0AN0fmEwzoYH1y38X3y1TXTbUdesYCf1YhhKSayYa7loZD3r
tGErMaRO6dkFi3JGBxnc/GozxGTNsZbPFkd93dacql2me1L8Gd7X9LEV3+U0
cRS+4fTwQY3siRaUyFb2ucA6+me6yusJ0xz53Yue+ydNJRZjW1xBKrmGCujj
nVJDMwDYsSKXh5eeFwglZ5gcu3yUPE4HhTmwbSrlQSBXVDF2+nLKvJWBQOaJ
48yiKP2snN74hlqSd4jjn9Pn5neZAOOWI4GjsVdtKmmyAcKZJ8czC+M0WJY8
njsoNgOhSHmXER8yx4iiI7YUwkwsmuPf9XMTOQSNZZc8IGVukshuXTt7KalX
DyiI4T1suc91rud7CMjkUcDw67jNs/sC3pqSDnWo745CnvDP1itqaBO+XxhX
Iz+HzurqNSUFf04wn5HHZrU6P+7FS188EUPc6enMrXnipHxtiFa+a/8ApNQk
DD1n4gKMI9CqustQM3g/f291qsy+5KTmHiGvn5r3DUZRHfWbobGnt0+baWxH
nXVAoqvPgtja29h8ZXG0D70nlvVuEinmw4XQtF382yaw/6bUIW2vQtrOgSfb
t4GgjMx5R+YoGDBNygv3AjIZxo8IzPJ3GE698H2C0T637RPb9/tXycgH0vfp
yC0XF2BqgHq3BDdeLNUngd9P0Do/wbm/GNuVRnHFl6pSbkNQHf6Do+xEzW6e
ooUESZ3ma7fN+hWc6CWY948KzpXUWxL44Vd0xJPMVbSWdCe1GBZLWIfsdx0d
6YdbWXAgIqi7m/Bkzo1YyrhI6KaxUcrbtP9EZ6YK1EzAhD0GQVUzjqGdm7Qf
v3n7Yhxkyzkyehkup49e/XKgQl0MBs94aqtZvbS6EtxVL6CKs/aDldTSgU3E
wotxLL3wPsZ0b9FokSBvW1hYC+mquAF2tqFD24R8Y4jYpHPAIYlG54qjyDLK
a5gsFctbuJePu7IAGu/nXDRPZ8npfQ+174sN3IpSoyKuSyIL5skhDH3Jenyy
r+RgHEHo9aRxqijqZdXtzGoOkWVx7YhMahxiFjdw22ll3fxHOUJYBqrZBZZc
fbH8gWkhwhaXsgKDTwEPfirFr/EgMmhJJS2kLtzcQIEzx5alFS4yG2ffr/X6
sb0pim7dJjCapVrK5eRU3uimMOw7Z6Cp7RENNBGPcDrAI+MwApyHr9HOB2ph
dz8FzSHjebcbAafkYEvGB1+77HnOe6K8Xw3PYjSosfRFdKeBSsFv/ZTYrDDU
+t+g2OwRq6/fYEdewyIypWoQBaoiS4kjJWkhjSnA7qz8ldE7DRLrR/TY1IwR
eXkZe60M15uFMQHj6lyYCGxuWSslRm6mHUMGk51fb1gEoJr9tNSruLxqWrX9
4OMBW8R2FhQd2JPg/mTFz6sho8rIRqxm1GikwqRqbx8IXTKMrnPhDFd9ZIn/
yfyMrq+IVLq6qq0mnDJqoJAo5wk/0o5SaX/lwmVdjAM80cjg8AhzGbmFYPgN
vCBJnwe+Oo50faiRsB5hhlj8mAsns1FX65NI8+DHctfPkuJlHZq5B+uA1kEV
oYhe0NG+NYteLs6lGJUHZrNRiFuGrLEdbJBpr6apt+D/SAwOU5ZzX2TibZuk
FcJFRxxZUisJqz0cPO5QJVx9USOL7vLCrzW5JFJw6CjtKBWLtAI93VGJSdti
sPtSgofPtqj0Ue5J2i6NMzFePCm2gBUOjXNHZijgtgsNRHZmXLPXgASyOLxw
aP9VH0cxgWp9s+s4LY1Ox1c8w5WwZMDbnBhhEiwkCefy5oauBKhA6GEEIqtV
LyNMIDyn6WhYAVA4+UnbHLB2xViG00BV//tuTaOhnuCo/SX8jSxhFZts02qu
dU3tXWUNXKdU1ndZONYUvpTQy8+3fXIoR6XzJkiEovANNoU1B3JAY7qtz2i5
XViKkEWa/In3fPh6UaMtpg4OEPtDfgxe4yYZk6q98k88Hv7RtdF/c6/7bT+F
i9gDr3i/BquAKFTJqP5IsgKpwTpjagl9ymAP9jvzPfUbZl0t6a7chHQM1Oyp
3mBy7ObG+O/+TMzPjVY4LlIbsaiogUtxeVCCDaHt2nhkKgXZBEQx3QEda2Qj
Rf0Xq3X96+k09fMgKEMJre4MJD1L0YvnxWxX+N16AE3XclrGjRiu2E0DayCc
0fsBefWjvW6jliv3FZtdf9J4QGAFg0BSWdieaFh0pN0p73JDQ5b073K3NGZk
EYcoyR1iur7+2UcGWA/GQceLygI8a9YCa07dcsOQ+7tPOiup4bOGuTySNMW2
G2VSaaTgOBBCo0aJpZbNQuEI3ZBVMppB3m3TlI4GdUP//K7bKP2Q1B8yXOuu
EFQ/OfGiPRbGZ35YOYSpatvNe+4hdIWFhY3WvTlycLO3kgpyk2gYoH2R3c3U
UTAwrwuTThib0PCirn8X89O/mwuEADSQ4xo3V2PSRTwulMyh9kVfxB73smWz
/y78oEX5XD3Wej2fTabKXBwC+7YiROk0ORPDTBgdgjBlLjFvrRu6wgLVB1zU
bSacN/Ha/0b6iQ0AqPaQ+1/f2TiJCwdm+9iDHIRIVHz6+9lmTO4qv6l9WmQX
wkUJgm7P+5JdEbswXC2HYkY0tBOjDEHYIGmnEsBA7zrfVlv+T4saFXYrFA7L
dvV8eMSTmueaaPd2F+nlby32S5+nuDFHrEhWAtd19yqbw72xZEXY6BiWtm1+
/zxl7D2wrA24h6+akpk2scu1lvXfJhrgtb7c7nQt8un9JXHgnjUlSS9tUxpY
x1xpxtjXhzonFk8iipUDn2YTPBnzyU346UmlFDtx7m2//UipqP0QxITqLaBw
LEwdxzCB/CN94KTxwsGAcD1WJ2pSISkq/PLlP5VVk3pvuhZa7nv8w8shibRC
qJSTdNNV+SqXZ6FxoiNzk0urNR+tUq+1dV5WMB1mh7fDZ5xb5akqfvpoFKu2
R+bwQ2EcfIyHtnVwg3qKPj0Va6Aq60XF1gcvMp5T9LNqJW00gQBhtR327pcA
VStRRRBDO8aI7fWfPT5QiOzlMdBraW6QxJ9OdCkWNctkQnEs7jmk21wC6Myd
bdy6j2TKytAG966IFzoYTLXC0MjnyAGmDrMeZAr1eudraceWKFhoOwfv4WTr
sLLW0CRamkPr7I7C6CvYcwu97NTSnVANQFd74u44iD0Z+SW43i3yRE/cibSB
2XkxBal9eDzQDRp4j3ZEV/1yRsFSyF9AdAPP152q1XwxxwCwXHHWxsyE1Ezx
sf195blxhTHd6qwbpZ7TKquK5FXIPuys/eZ069Q/SNoyHD0qAAnUJZ5PboSr
CPKOg0juYdcEa61xrsdEvScTX1M/WhHp499FHT+v8WbRYS4AA7kZLNsKmhz0
Refb/+lIVjJXyqfZOqoGr+9Jyq0C/nILPtYlgtjeBpn8jNPMHCOV5IMnnB+u
HrW7lJHTPArXIsc347kx1ZRAX8qWnr7NhRu40rm+EZkfqB4Ec1ZydtM/12FA
rDL0pNFNkO3vMUF816nO028Mpp9fAxWYXVjzCtY8ar59O1qrSGWQUZds/6sy
f3IKxa+UI9Vzk110m6mPeZlu2RVGny05MlmN7b5FJPvLBpDkYko1B93pax8B
1gNTkj05oTvWxFy52d7lKXkyodcBzZkIp1Wswwt8j2ujiCmt5uRGK1jyFIRs
vIQyQyCuEWWWE98b2YQkqcTmj3+RMJrjiPsVDfSeZiQR4ddrvM0THYsUUzs7
LKhc3c2omxg6CPE7DFo5HHJxA8C49xn3kf2Lm1pqkwElzAmNuDVsfaUhA4jS
3QAYytqGrVcetNCuui3s7tRanI45ThMRXcgMr8haTv9IRe+953aVR0+zmc/n
KlxB8Dat/Y4apmjJBQ6BPG0PUdogyvKFsvyKSVuHMVf75CMWC2u9/v3gJeKx
o0bt0anlStKfF3Tz89A7HbXsOhFakpnsFn0K9N4+juAYAAfR1kkNna/d2jTO
ZAp0c//GsVrmEs0D8vKPOMiJeT4wb4nnlutlEezS7+Yytr3pp6ptaOYKZJTU
6yOdqV3sTlRtPts4+4m2gqW7KNQ3gaZnqbWEXQl2eBlNC1X8kX2CmEUayPnh
Pk8T8fmybESTcDyBmxCz4FkfpByeGk1RW/0NCv26Bn0HrnVuvftv3/y0dn45
Qz8yv7x65DjnJpNPuamjy+AGVhC7Jn2L4ao+4YzupL9ARZuwZqaYEPcjI9Z6
eQwNNrfWm5m/o5rlBsFp9f7O33zDFk02nBnHQY4WWlFCObA7C9x6jAMJybW4
k1XIUTJphnxh48H+ULa6g2+rfe2dAMi5TmdlLuLEZMVqR1ohj4gfnsLRV8Dd
YB7xKiyg946afoQJ1IL/28dkg6BiTQGFtr09DiLxejVZ8sRtvPwoKCKz/s2P
h7ycCtU8CKp1o8ulfy2WNbqOy2IvaGYADiNhz8CywqJ0JIUkNFt619P5viZM
mV5ohLFAjfqzZNDmEahDi0vGGkb3vctjXBuXyYMC/CePjGJucCdyxI4X9uDW
XT6VEUBkuKmDzwUKa9MrxoxKImSSQIcKDuQ+u0jyRfurXN5wqn7TXw6MSFt5
kxIseKFFjv9zvpXNjobMjXDFigYIQC51+NqeNN0Cde9fdWhJhLn7/X9C9HUg
UJasfdFsvENjoMeycJHL8u/hEaC0y8olhWE3c/l2p41EL9g0d7IsaZD0CIit
uRBiSTHGEJJlNA9AHL3r775GgC6Y7x8bESP9rw0Q2OpRk08LJC48Q78FvbKK
q6SljSKmVoac4fUFWW0AQKu1thauGHQI6j0rAOHLLHaYLXe+4FNI/PUvtfSw
yTLlslqZdhEO+M5OWrpGbXVWxTUPptje6xkSQJYsxahA5eEYbjCr97h0OLQG
Dlc0AkoR6hPxc7oRKY+CSCwqyBmtFlEqPkP41CEqTSj11GptHPB/7XwUy5Wn
6F+3o2SViv62eoXK1Yk0SKMJV+TVPp+yCNbuGyjgmSafwzWvUDPIXvZyI2Q1
XvBMWoE+mr6o4a3HovKStK7R9zGLJNemLMbYnQ2YuUCZ1co2hwFyCYUOPK6m
sJBt4snkzXVogVlSUQMwuYe4zbKtNj93jYObVck4ZOioa+RYv/uVRIND5m78
89DTQWklVKX49aAZk1L53og0QAeJNesm1Fsijug3fcZ9lpd1KHD1Bz2HZzze
BsGy3Fj/JXiHt8EUxq9sraCJytJYx+mpGN3oPw39EmtwvOkMQf83zqsd9BZR
Sz+DQlNeOvgUpUY2LSiFp2S0265arTMennPpPpkdbObtxhx4mjJ/FpxtuCLx
BJS35SROW1eWKFV8P9asynMM76yS3G1PHxsEMCMkIjdRZCpnWCBOz7bripv2
paqkEHXyzhP9AxyMBFTgD1QN8FEuuCmNLLGd3UPmU6r5aSs3XOwTMqcnWqo2
gWXfqnEuFMi+G99Zl0tQpK20kouQ+AutXGSxbKHoUvOOdGqdVMC7TdnwwJN+
UdWc5TEMpMFliEMlCFZM0PbAsg+OFfnYo0aI9Y9dEU9buI2xmecA4pOb+GqM
C0RWe1urHnnGfSHwoZl15hymf1f9n64u1yHcsebuoGq2QU6QcTync4KsrtG5
6UFN95XbNlriPszji7uq+7gkI0KpWa+3tVdmbuav37T3eMbWkLb8mLNW5Eex
0jLp26IqqbYlSjnr/yOzIFqasUHItph+X6X0gMG0mqfMhkw2RbAREuqtyQ2U
QE1D6h3vsJLicqImNmcgQWuObnakR5MbbSQxIMed7im7lrnZSRiEolhoRCWU
KFpZYXhmmUHiqr8a+Gi+4d3JdbKg/L92p0crbRnzHan80h9e4Hu3KuM24EKK
NaZqTK5w+xBQRe1Aw69stdOEKN/6QhAc7V+mHP2j3T9V+eI1GI9Ihpz/hpKG
W2+AmPVshkdhrLwscDqObuvixvAIXI9i43ECIg9NtWLGmvhXL13esEzjO7qo
Ft9M72LRY/5/1XuX29L/h3tTenB6snR/4mxuim8TrQjnlztNT2r4SlG73D7T
fxsVxpZqFBh3Dx6IwMfrHJsS607Ban37D9jmCubJeXDSoL1MaVwjc3WDqQhE
2txKstjf9lEG1saWtca4dvAy2YFW/U5xwu/4io5xOulf9g/aczI9laK++XAx
5YkFS5t93t5j87J6l8zNEVLhSV6Zm2XvyVUjwa0YXi6BQxl4660HfTFs3Aii
6++kH5uBR9IVgwiQUgtx1gfGoEH01AGq4KNQfBlmsq2mrY9libu69IysiV0d
eQFq21zH2hvtNiauCh+RdCrUg9W9nsuxm+H5XHWnR80pOaD2Uph8x4yCxgQl
bSO9e0KGVTuaAuvFXqlIrgaT3zj0mFuFIt5tgEeg5x2VFS19shO182VjE2GX
h29OyunOaTr3caPsK+DnNqH2WvwYXrknC3NhEGk17yYeG6IeqlUo8oCvbL05
hfjyA4yf9tsiij7OIEcorrntdp4hvucYsF3FuAeqUoURU3x5kMkeo2lbz2tm
RFKj+CrllGBzfDNcnRY+0neuaFMeYOp1jktiEw5BU91BWSockgsV8Rnsj6cH
rxgJKR89R7Dgi6vaEGVLlyco0pYtS2V/YcvolTSnfDfyVLAkA6T8bu8GDRmP
bAwKHjxQKg1OlQolIJAnxSrHrdMKrXg0csOZGSKBRqOXFRTlHESuZbd8GA7v
f3ax1TF9M/ORzw52T1seUaEBFKEXC9ddtYRtkgnL74AWKjnIQWUyopXH3tvK
tWsyBw3nNUPMa42fdH4ulpTyONCGSlTlx37SJz3d1BjegM+jUDtDaVWb5OAc
bnKBXgGwcQne9268PBdyrbfY8Q40k7O4pdDs2BeVHx5z+KHOzC+u5CNdF9xw
ocvfEUyxA4dW6DY7gpq3jf0omU6cIgBx6HQ+bko1KpcX84zEPxt2t3mrYMDh
4ffMEZ+T6lyJU+b/hs8SmM29kuyFS2yhQAeYZWkiodJQVKzdZT5QWizhyK1g
BKNjDZqv6SxcQzqVhwnVx2Ng+XwdRnFKha2Krt2aG0wL0JHQdmUJLtPdyjlY
Pz6bHOo9YaWtg5EHo28t1iEv1k0Tl2V2sjRoIE+ZnXixdI2nldaaOiNvtq8B
caDCo49W1Y9AgHbfyfdlrCrAHaJzPchdpJXi4UPpBQ/aPtxWmo9Ar6EHFyN4
1hIWl1dIDd+ObQ/aFiBCIrF90fWPNY0SiKkq61OQ4bkvGHZbdpscwzW/zf7X
zlZZTGjgQQ6WtrthxiZ+YeEAbs9HbTaGZsVRU4u8NeDGOpb58Fd39ynv+IpP
m054KzPP6Nl1SnBR5Se0Py5HdP7wB77XtiXxftWrQKa/mhekYTh862twaqef
v2p8KbT+/8/AXq3LSex7neGE5fljUitAjfDrdVFKFH6Sf4bar+O3TDNiS3Ka
DJQtFBvDu3nL/uornCMLr2tNoXKTBr8g9YUXlVS02AWOWB0ifn9EVX/3G5Ux
mPr92/Tcck0TUqJwF0TWCfS47igwfWq1N0kT1OoRVoky/fQ34LTPo6KOF/ik
fxC8ExJMXHuWgLZFNmpf46gcG4KadIPYoJi3g7RwEw9BJbuLXgfBWPG6G6EQ
iw8kBribj/hPZTHzMC2OMBpW+KzjrlWp5pP66OIVlS0DCNfsoo6WLMlFZYK/
gEBrjqAk2/EwEBMJGljPNDHcHk+j3dGJKekYaDdFvAgnYc9Qx3V8e1hBTLGh
ZIMsYziofSiQ9GpiHm4a4l+3bUYmsQhOBGkNAyUq/vbdnE4mgmAFHgNiPNgF
GbEYCZ1ncWSMiz2JKd3wRpBKs76r3EsDx2JIIsjlyytJA9mj54y+WAZRG/dI
a7VKTpD+qR9rnfRKdaB9IRfx69UNraf3T0OWd7skYhhI+iXgCy2/bHPFjpRJ
TYGaOx+ttpWsBE5SBZZgFQuRas3TI7l4jIm55J4UYdQs3mpf3cfriRBi5T+b
2SCUwky1dVKyVGnr3PRp6kZCBBJ/1Uq1QO1pCvJaB1V65fjSY8YsoIoeQbwJ
4MKZZXvViplt04xlUBaYORNMTLw6bnws5MyRImyc4Wql005VQ206hYv7VCCy
gOWl7evBp95475sxi2RDBKQj6PMeECLxF5iDjd0SU/fLv/toAA6VV/PaFx0z
AE1tBQfy0md9bhpB8Qhwad68ZSOd5pzE3nYTsK+Ahu6B859Z0KpXOK7C3iwi
NL+GNccEPDdgZ6xgI/GtAyy+MXPDqZrwDwtmFjlNKUEgMXZj1FDGAUFSgeh/
JOjWUxp46NOUNWtWMEZJHECm6GwmvX2YznfvNrIRjPBjEPtBVbXy18yuRS/K
WQCUO3TnJ83sTSnOSSGjd/meWohBBC1+ZcRuZckaMV/YTkOOShNwnXon+EEn
uK7EJinUhcAsiK7lJ0NzmKzc4fNtrDDCf8lYwiz090rNuRCiA9o+wktYfmcp
z9gKl5XcKh9fefA7BvmqwBSFwJr1BIit9eA/ubcsCgMTlyeL9HakENKHhe8K
KxPPn2cZHdxRgPsXChfEK2mVu0Ld7TBX6hF5eBAN7YKnDICuz4uKUsdFayix
iNIF4ZNnJrWfsusoHYQsFWnY7glreuZT4lM2CJM5UVGfRjrP1LJtGK2lNMTI
D30LTHGTNcuUi+euET+nlYeNufrWbV1cIqjojbsfDgAAIHVyedYWBcO0Zl7M
Uf+lg0OlySLYx0XIfS5ufIQVmZaA2hgSCJVx/gdWfVdCOoDOwjykgB0eKCcx
cwrBhZwQnSOyePwdvk//c+RNqZoX2FtoCJwgOmt48+Q2BvYwqic8WDjhUsjI
OryunKxq4GKWrg8AY0mxvJWGCF8uKRTpcdy79T+qtmYrVIoiBDJekLajRaGs
shoQqONF0KU69YfkpI2yldNuuApXtuR9s+Dx3dCl53UaI72zRNUmB2NzOLHM
+q7YPL7P9SNeLtRTRrYIsf2L2O/WvqRAWs30Yfu0U4SF6Xt3eiSKmmUdge24
5ZDUoEpdtBbUFET4AMHrKJ8u8//c9JbJjIrq+0VSAmfyftnizWZJUyxXGn1D
Rwve5kqjQzdqFfJNgif9TWze/0zuaadv0vBZUjd5sNB8KN/FnXrxCASg6yju
PrF50ixmCq3mZjmibobHMmOgOpsxEZ944AhX0B/jZRstgodeNVi9t7rji9Fi
bDhWOgYiOTsjhfl2NpWeKOTgoL6SRX0BGTdMzNdpHmhe4U2OERmNxAOV0t3B
wuIMR/pMd09Ina3JyqQhy3uxIYjmWnAMXzq5jntNX5b/sNdsS9CXeSH7xGYr
ARLZbMuD1Rg18kGygKyZaMdbbBscpdtrHxjRwGYt6+omZsRSlkdWuBSuqltK
NwS7Wkvt+/VKs8TgCrWF0vBhYQJNPwtLtEmp4vzhKEtjN8eefdAsCwmvt3Lp
yFVF4YVXWH0wLrjQ1fwgMmvlcxXv1nR6FvHxs3GbtjxhScPoXO7Xl8pZJGUC
cMEIgl3Ti6KnNQpksH6iuWTe1xs9v+02zLjVU5I4u6R/00J80ByWDY5oB279
2VlL1Jt0+UPxHYTPNP+uT4vIUCF/zEFNqYXWkdST4We36qmfAGx0AJ7wKeXb
4AMe8jCYvF7PSzQ5bT+WajPCccFYWvfbAdIrRx47rv19VcqV7iEUNHN0XlTy
zIFAywyr6HRKzvrf3AyvDdpBE80JqOOQYYCcRpEFfBnWED2TsuYN/u0mhOtJ
RnGGdyRbivcMNBPu6Vj4EVg1/jgzLGdRmWHFiBDDhCojpQSaF7/QTqLIfLmz
KKRZ6wNM+gFiEL4oVkNzrWjBRKC4+hQG9CH72TVzG4CBswYz5UODWz9sKYJp
a7TopFbyS3UR97Kc913kNTKOm4GaU6+V30dXc0mbAmgv8foazlpxBhaKcql3
/AH2JMF6Vb8rvJ/nl4Bgg+YkdEZih/NHkg9YbGfqNzUzeTGU1GNORubmw+U4
ROXYfXxGnamOG5or0zj8aNxjAxJztqMR3wdAAbCTFA44Gm3DdTrVA+dg/3hV
hjZzNhijyGmXuc7Gua8HyGjJxzRVYZXJaFGAbRF9ZM22B4hAtI+L+aKqSzPv
fcExRAK8ppV1lRr/ipz6mDdKkMIAxBhklTbiX/WanvaqA1h1bkesbfDcsQPU
DnX2snZJI2CSlUogGcdgUad0VVZZEz2wW1tN4KmiRDAiZtDulihIzGjM1P7t
2RHbTHxaI8v1Sm2096bomOB7kB2RHdVXpfk4ORqch8/EJ8dP4D22Rel78acf
yyVZyOu12YQ10w0Uhe2KMQPnK6jnkETcbHEIgoZ7/YX8kPZzaCe8MagOm+2T
U4LoYj2ye8JDC6NH5BONlY12sshbrMpFHAZgZcF24bq2LmOcKyUO3SAk6obg
f14D56bgVuJzYsJ6h9H/A0rFS6TtvQmmPbuwmQyNUOXJ44518xyNclzXIyAL
ElWge1zaMsEMr4wKRUSkjADg+aOhWRoP5SIbvp3w5cRBz0SL/UDp4Bjz9Ffk
0wYuhPRAG+PEGb6tgMu6iAqQSGxkZgngyDh/ZOu88NXviruNm/5BHeMDPe50
ONvmS7T9Nj08r9psKBx+ySSSfprnb7mLA1k/QjAMuhHkhxuJciCj8g/zKPkI
EDG96NnPBXQI51JmV+QvaGwl3Z4XekdWyGuCkRq/9+F3pCWMCfsoxs7M53jb
nH8A+zFChB0Z07ktbZhbpo/JPBF7hFNjwHp8dTHWAKDH9VEZqzsZqVCmjCud
Fc/kuUTr3Iwq1O7Bbl8TriOtHMuzXr06JOep8o6+ZBCZYFaInsOEBVgEzr8b
wBxVtJejRiQJM6JrVxpJKeUAUyzgF1QwulvZBXjms4aCz3bAVcwmtCWlt/fn
F+EE4r0duEjLba6vD8pUif0kYjTrqQO0XJlSiKBj2E2UareENpqbecueqIOq
ip/E0bWNHMRCVBGgckfmmWWYmLPHWT8hmiN1mMWr3S0xWVxZyjUlSy1W3xqA
Xsvo1k5yzqznQnjw6e+uPy3yuJRdgRQnVhXTPQcGdkEZqFgHAZI4JOiqjFEl
0l+83JN10JB5zMBcHFSeFqDLmqqfMeAobp957ZSrMuLBCN3287JDA2jH9IHC
KtsdKK9OxwW4QnbQMsWFzqUc4GB2mXuRdWAN6+SwMvb6iC/kVjWt1qtU07zJ
YOtFRBepkeABILpEgM1Jbbq40V5RL2jPU8eayCuhv2SlKScmEOJuuy3klSGI
rxkBMHr6v3m9f+JxPEi0SXoM2U5B9kKs6OiEc5Ee9gUdIz3olqmfieI23tit
E6T0KSM3u6ttcrDTVhC3kK9aRITV12jxdaVvWYbQvurQ6lH+Xe3Oj1fsnu5E
Y5mAkQvX0hHD35Ni4rqKNGvvYtljXcz3n0FDz7QVxK3P2Y7iDEFP6T5Y3k/3
SYdT5rNMnnZM6Q784ZwIPQSWTTBZQ0+rBtiIOzr7hwL2tAY0IClFuefPilYo
XBgTvC+YuK4jnZJpci9s9Di9flvlkFEXOSlsQHegZLDwkvBgoq9ReH245Dy9
fulq0RKLKfHlMvhiuR2fDkJDjf4ZuH1VzCgJ64lRmSOYZGL2OSGHDj36gsVk
J+FJWDXgfQBIvcueh97lkvUV6lZeIvm1AeLI0d7Wt794T/9kQq/wL1m106Op
fGzoCQBc29YdWA/lbE3zH7vh4rThSF67Rl73FmtuvkTJOI11ERatd+gbg/wo
N0lUjClJjilgMSvwysnR8LT/pAFwtIOMohvSlESqiFk+K4yoRjna+pvSnSF6
omxnyydp4seaXJA09Cqk7L/9aTyrQsmHH/cuDE1PLESVQvvxcWXSNHzmiD/U
t1wH3f8toTRqjV+uKCgkMnwts6X53PXv3oLtLSn9wbzC9QZhSZ819vjnt3cF
J617ybuJJP+hhaXj/S3pHqLtgtVsoLLoVVNFqA1+T2vzTSj9b5HxoM5dQ4CB
R2P7OrjKla3b5mmaCWMAG9jtKDUzNez+PrDS/o4BsnzRMRQ4lAPiPOb5/nZ6
r0Z13dJ93wfFpMakZJ7cgbkwauimOIaBYpnAo+4N2CJ9WhYfXVSINvyzEkL9
w+5rz+Jnvs2pufKf3LRWcv0PZG/4hOwxomlluA2TR/8Hs5v2PNTK2JDrqHko
a47NcFt8qpxey1gEudhb88Rxc3NSPClAXQO1nLydoQdME4cl9RmuKSPRFt2U
f5iHE/qjpZz3/qo5PbPybbDyPuQEgRhzHbNs9qSC8pCe+voH6IIGkFzktrWm
MhWYq03Iyj4xdAeS8+S3U+c4BmZf2CbR5Qv8hBxtZyvoZL6Loup6bj4V26qt
3iQxnWN5rLJIcmcmukZtjl/nVSVRQxvhcDB7Er64zKsF/tmJzkezdnb8Z8aB
EnhZXc+/KDgZjDAUMDc3an78c0H4nH4sm/4/uGcBrCIKcF4ctHqJR4pcNQOH
OAvxjY6SMD84M1OBkEZhJ0YtiZBtENCN6v01GJq4pf6Rolpzighi8B//iFks
aU92TvJNfoXOVyX1SoAgFkQPPoFrFA58PpZXUPMFU+AStvFsJ8e2/MJxzacg
yHPZsd89YipUYPRdoQ8xDOJLa0vgHIIJpUxHhFkQ4R7/sFdhY4UZgOC+hn+0
Of++0jGx3YZgV+lWBCMERoRoEGJwbzGKKFfArlb8Oglk581BFVe7c47IWv+T
0lwneE05HNo+UFNds10BXOGIVvMlflPdPH20F5N2Z5JPjIfc9YLLC2SrvwvA
Ja0ISzqnzqVYHqyQL+HCL38PBZnC24LOoQR6krEmbvZG0f/aD6LRnYAw9zYN
0cgf1RAYQXczhsHORqY4E+vocny47kAAo7boAR1Ha4cY6jNYb/lDwQWlJYB1
Q1UNPDG9k2sDPzjikQsN7rvm/z+4aZlEgCageU3lgrw/o166vJ5nJzn+XW0V
dfc+xgyRSy2mIW1tYRwCuFztTTijMPNspWaVE9QDiAp6GLx04pS/wU4PUaHS
LsMpHowpVXy9UQOzjDp9f2AqeZxhqYTa5/rxZcxhC1npoltNDHiVUWRLmvBB
p5ztoFi80o09Znezs0Kf4PSvhHrS1gFullURsojKfEafrnwPYkd90utTVv3b
xHbmB6SKAlByTH/6SNy0kC88nW8ZOjhJtYgT+cXAward04oghzbeQxULgg0s
pA4lA4Lt+26Y8i4qYhEYuBiSfqbPXRaOQW3Cv/KFmm0ck5q1TO//HxwCMoZM
7sSiAX9DHBTV7gB6di3TiOiTtzFoBw7uJhDVYGb8B0tJ9o3Utww/5wDVLIVN
buxP5tljE1Ud7Aeer5oi8xjKsij85e5Rq3LGl+xRaUglxD7k1SvaGFzX5IDm
aT5IXuvoFrDqKJva+aFcObxWT0nZ1jqUXg+DQTIXtiJDb9JWcNADczl3ekxP
ozi/wYhXHtjGGSBojUdwdju7a/Y5ykoRY2AEHbRnuC/kxSLnrBLllIFNE/IX
uY/nl++hIka8dXeqSjVeIQx44xQIwKXWda+qMJvq0aKkAhGtEpmuiG6w6wNL
iQ1xZYY4oQqci5GHDBiL2not6l4MaMwwATBjkliGrI1Edwrdi+rNB3sfWnEj
xeAJ9zjHC/vLZjbIIh51z2mHvuFwRpkI0nhHygOe5mNmCWBmSRne1Wsh0n/X
78FE3qWoEi/ZLjjeqvws/M1BhKSb+Mkg7TLxFE7fUNAcxN77gWDscmf/kp9f
XNG67TU5PoeRvrLZG1Mwo+Ku6W35H+Ib1X5195dUZ7VvmOzd67Nh75Lit2Zj
3gsho6mfCtBT/7r/X45oIyCSvWPo60/ZTCCptHIn5Rw5mYDGs1I3VIaOwrjl
Z6M6qdG3z0dq6SY7VhFXXN3Yh6ZZA9im1DZfqSlKLyCjQZpErrVMLpIOpHNk
jrmrnBK3lo/2KV9dqv1I1uWAm9FID0tpC6lM/NUuVM4+bj0Q5IVeF9f54+cy
UqzLHc0QnbGzrWfTKPx5Ypc/p8f/XR6cGAa6PNSSz1upyai/vmW+9es6cHcd
Mlo+I71wGgGN9xviD1DXY8GDiu+ZArTHDMq2LCz7scZ09DEfAj/rO3JamMUQ
ZUGdaYN3t92s0EiMbkAkzrSL1SJKu+tCqSJjE8qGb14sdUAVmBlKldtSnY5l
Cme7v+NVllrTjDfkqdehMK9Ata7rAzXD/3MUXxsLy9Ou6mO8EO3vbitwqukc
VxDSUYMZoqOH0KwHA8k4JGDEF6qeERePo1W12jaUTR1Y+rTeX0ppKjGtAMmA
DNHq2/TFMQhSDWEZy72PFNPUye8lALc5p9hLzI6aPIKUMgYRQ1NivcgYnZ7e
8T4R3+oJ+CodIMfozJbh03n6M3UNh+7SdJDMkz0m7b4IRUG+dzYP9zKxSrsr
6afPYGPoFAzNAMmOHmnAzS9NlDn8LbTnz1mlu4/oA7U8Cbr4pfNMR/KdTNWs
kkb/r890FEnQlppGhUXfzqbA6JglbYwfyxX35WHYPiQorwayBj8irGF2bQKH
xQf+P1zyIrMaJRJTN9AoTdY2wjRtZbiWHRqe/ed26fozHGtHEV+r7RyZKNbP
cOh22pnxbucKxi/y0GfuojrFrBhXKyuHC7bfehJKcLd4ZqIZBd7Hd41RdRoO
2396MRSjovqw7HlMBfZOc97QrWwUgvP4PzKayeqc857KM1v+aCWsBx7WWipN
jSoL2iaqE5ZJNtw3vz6mKqG8+SCDHwO4CRJQIMVH5KTu0zasb0RJ9MAGUZ7N
rNclkXXMndUar47i4qpH1ah74bUa/TdCwvTweVPRaGYIw+5MSotefCfoNySD
ZqgkE6xcD1+ofDnjtzoxXNutM/Vkn8KRP/OP6lxHdaz91z6L/8feVHac2aHg
RZEO1LbTVuRv5iVAlfL5qZjNFrMJhLvBplcUVJdZM1wy3HretNCAaHasGUen
h+G+Tu+YyLc4X+QP9kaExI/G75pSS6IsHHV2UfOME1VO4ThFYtcokgjkj50L
IDtcv5QFM+K+loyX1CpVEF0tuzrQEn0oPny2kI7FaCMXTpMAtFpHwvYgGES5
esnonTQOuEuXEbT7nB1uMKD/rhCXfD4Y+d411PrYIraUc/gLE8Xjp1NvXFqs
+suA5WXpQIekcQuQ4p+0LxLOXeNjnwZ1pDHhm+L/fE9HTCmMnK0prsxfaMSK
OWnqJaBtqcVFb5OywlX6kAtSAa49qNRTXX9oM6kR7XcLqiwhlFq2zWnY8kBh
lHdmmXHuX/oCwyL5JiOCgMZp4HOLi31K0Wa9J9DCEQswPXEOnBeQG+HGNkjC
e1oGDhW81yKgEju20bveA/Xh+hdkBLFchLI71hDXPymgGrcQCl3XA3vkZY4G
TfaSJzoplkV3wJoZc9QJ+bXJNuMeP+8OcDnWII5vqZbL78n9i7vjHNJS71jP
i24NR3LtIkC2IHUuFquM7Eo7LAUFjFWYaOTPIrlTLY5XSS8hiGTUmScFaM1E
Ig7NghMEU5v9psPQ+CdVM5SBXI2PUQwtjNElADM8UOxHlUKIhyXrFj1Yis1z
p4d8lfMu4Ug61RFYWGaUm/oFdeDbMrFIT/OCwWPgaqsXqe+lQbX6qvYoSLPT
CNDuqNYFBf2gAQd4OWYcVTHUFA2QM6uEbvYF26X09l1wXtFFLUDUqK0sLyGI
gLW7gUZ581D0neToBg2nxlMbsChYiCnVQU/ACmi0vIJOOnNb1iw/QccF4wiF
+e5EQ4Bg9e4r8uf0nQ/jPmOQOdE8GDAjnrPZWv8X0utXYonEE2rxkteUSHY6
aCDabHxpet+24nulx4HU2iHWHrnlMnlmRCcTAUvPzqAvSneYqLPMT1MX3adP
2mW8oxgDRN3nONGn/vc0I33bcTNvSGrn8DfHaEA1IkwAewL7+cfuMc6fI+hq
OWvxqPPQ8+kxiCDI0SyDaup99SMe/2Fa1FLIOIz+nbAW2VXXp/15IOjjuQSR
ZJQxlhbMuf9/02zxstpUpB3K9cve8nKz88yFqPuV2sK+n1IQNZjlkoCdl4cM
5sVV+NGqazQzDanO/pB5QPiGdA7LBAe0zr8Xf4viROaY0o8La9yZ/CBoYIVI
SvpYh2u+8HXXEcFmfSa0Hzr7H9AkrHVzLyLvu/5ZKPIH7nNpPC7K+3DUP40h
1mNQANTUVogBfd7x55MstEsyBGx0BZUR+3b2ZpfD3tpf0t2LBHzPVIWL4uX9
hhWRGOVAQx5wG8DKTrcHadlEz5lk4BngMl8zRvEhPrMUtc8oKPsLr0TrQzwN
JhF9Wz6a/rG6kAj5NvYDSLy9TdHfFdygEMSKqOZzGV6OSwB9aJNhl+Zycqx6
JzwdDizpUawVZY6i7Y3fcRDZSLC21TlJ/E9thpW4cqlL3Wzdn0mvUKxFsFmX
7btRDyhQJVb7U7W0QWYRyhsB05ivF1mP4syNMFGMVKGs3raenHYNGI/mhy5G
qQmWGBTqDK7gRL6JiNtgaWiVLo7RQ6eGKE7SbSIZbDMbG2E2FJBs7vJLR7jL
rDpaPrwiLpTTT24Tvb9kofjolJuB+i/qQEG295wVl0T0iUq+zZhg/R3/afcd
GmKNEhZaw+qS3vPq+DuW+bH0S3OEcPP3qXjz22Kp8EOVb7DfjH6SBE9Hm0R2
zCGk529PN3ldktAn71LYzMSCicuWgB+HDnIfM22c79W4/G30cAr4sT5LQ7eE
johnzLtKPZeKtu2OZjIZRcP5QIJBsv6+VoNBkulldIQoLXc+N8yogWwYsKyB
Uxh9C4DNvmpj31jd3v+zBX5QxqTRZ1JSANfQDwuBjs24ty1WxP7aQEbYP5wI
lsIUvihUbQTrZi6aJuWAQVuyl/oXCnB+GpNU2mgn5z9U0ZXR40hzVRaRewoI
z1irPs4ZSGSSS1pCucQUO79e5XWEAqY/uUru0I/tLPfDSCgacch3MB1Kk05V
1FDKVuXryyAsBqvYzIXJys4yEXLc0R1VBQYG40NytyjGmg+7SwmQf/yv2OK9
4sd5IUHTz94lSDSoGkJ6Tk6vqAzGAtiHT21C2k8ut2rEmmCXi5uegRi0t09d
VdahYsvoR6eUUMf591N7EDE6LHrqz3HKX7GuvmDHlRSgLyxPxvwLU4lzoY6F
FKNcYx/K5Rx1a6xvqOP1zGGhDz8Az/C17hMIcHEU/Jss85Xc57EAgS02fJ5f
pBengjLnx9gTRSvKTuLCEw8F10srVsAk3vYS+Z7V1cEargf/1TOE5TQQBgNo
N4+62m/22cm4/Hi7XcilASFpHwdE8HfDIUrTFituufqVRqZXDKziUioWgwh4
PinHR3ic38fyvcU06ICxU4uNCcC2icb4mc+wP8DKvbSOsFvYJ9i566mB//tU
yvVjMmAI7ppqQALmCzBZC3YK13zqFYZa1ROvLp4tdUl0GTUKBvvcno/gPk2L
9F6L0s7BHcsIf2pybhGyxMgRGNRpitsgjqfq68j4uoamC+gpeK8APxI4D+E0
SQzkXIdhg9tSihpon9MV+4PATJeOAy0Z0UsspBQmHmQrCxtuCk8PT+MzIp1j
KfSZOzCiNJWT5HUpxXZLLbMXvhjvVLJZLzXOW9OaMOOG2cqzFkVUj2vVl9d0
u26jIRXMzKTA7pC3XlED0ok9x6AGHzNm71XyVY9v/G0Bbbcu6JBGvGOKR9Ry
KOXyFrwzqXXbbLtzHR2TDGfEgJTkAx+4LwEXD4qCBNoikJWmBVWDyw68ek70
lYOMvVoiEuH450snC+JykPL+kfDW1L0/NA8/WTZnoFUdj9iQkTdN+nrmxYxg
ct4sn5CF55gVUpdJ7hM3y8YgTt7umkoS4PG3xMdyTAMFf0/MCZHRrY9SPeIZ
t4XQrUp72Pr6s3AAR6UzxuEGGzHqR3kNgsN4n9ZsiEbaOhTxGkYMslP8eeDL
2gPbUke9areruR2eGystWcdQgDk8pcKwtnk53KCB3u614DsKCOd6qoCT233e
sedr16qWUILYeBFTm6nUsRh/IOnzpjVw4s1htJJWHicGz8Z36LkwSNeYt04V
9aFUAn2Vby/7UHOmcvsDqspDo4HB144ox/eGJB3kQ4hkU3pMlcHY1NyXB9nH
S7/lsWWi8TUiWGEzeLti+JweW2SBTzuT6ZIXYlgxnM/L4ylWYsDdp4AHkiIF
xBZVaPQe65EnJBBNDmkpTvH8WFedsgL94csdap0lBdDu3zMtdRy6eIsc52BT
UMqdQ4EK7mVTRiPuLGup12zngEGMbiSykawTGHVKf37tfS0yIm3TTCL1lgwL
sUZGQwljhhEPLAn0yVvk5XcTluT3UvY6oPJ2lJMixTYcqXmx9Nmj7P1LflzX
2a29s1g0Ke4Co834/8XI7SpGzNxQGUI9lHLAUgc30iXdo0W6bcHSJHPCxOnQ
l29OzQ5ZUS0RkBJ7DAbSVTofY9cbsj1/t7oWKcODH3TEJwRDaQw387kTb8Qd
4xMXQ2GMXrWioC85t8y3ghOoGpMrVVaBLJIPe6frhCYQc1dsgUaNvqvSmtT8
wHDJfScPRhf2IUclEHccKKSAZcy6ICrwo6xTafvujFol9/a1uagELK94UDZf
c58Y+zp4ReoLniE7+iHKc22ETlAujlIHj1FjmJPJSEaqjTYTvacqrkbSPBGN
bY2xFCxhmdTxfknEGBOm0JVzyi7pJwU90HSPuIRZ4w3QnzZRCwD9upkHGZ0O
41gDyXXcHZFcJE3wuZmF5AW1CYfmcS5MsN29H64olavXTf5a+aZ4ZONHQM31
d15hsb7JBC9iJjs3vVPZ2bUlulturStOwawu3fG93UMEjq8dFQiY7tMJyaMi
fkcdFQ0GtNoDYiyPrmyp2xgcTSAsgyjuSsp/cKTNA4d0I2OSHqnuCDbIyLiO
pDfFpzjKHbRDzptfgYFwmycU96tK4guDJu/gCZnhrxVqer00suri+IFHfgNP
zG2j4ZXVbtLSHFBTc4MSYEYK9pdOrByIEzcwKzwe45R88xh5GKAQiSYrtb4p
aanSttmPKxsUDGCvNxKF+OyqF9ke67GZsFoVknYEXXkErk5s8wNTeXGUDZm6
I60hyc38a/M33v3NSg+Yl36NfnyGqgvYUGoHwMZkiP+E4ls0guziAjMtGINV
ietC7S8AkD0dGBTr43IRRPPlLzPqlPbLb1SLnOsJtL12H9gPO4cEgNO5irwP
N1Hq3uC8dTkXHRbCWZpTG5lzUSuDJNi7YXgWWZO6o5f0G9IyEs+ldrIlSAVH
w3aYDs1wBENtVZGKIWd6Rggr3YAW1ZOQ7okRPDfCqEJZXM5c3riXg7VNnTrh
R69Sbk9na9/xu4zgnI9v19msexfk20toFp0M5VC7oUa5Zt/uQoSsnxOOrUwf
Lfr9cBMn+hBo/4ADIfaghsXyBYNDTk+yPFwMkiB6gGw6kT5hvCEs+tmOD5+x
6u0uOHlrHxf0YA/f23I2Wjyvq7D2Y+ad5cDjtllzccTWGDFkt/TyBhxhJyxG
HzmEZFlXIed49phnIi9RKZi7j3qnLdsV6YonT1ldWOS3Kdzw3bepiFuaS7C6
HtqEl3KrK4KxJLhyYTur5FD7CMxysSMcihoQCM8Up2rbtFZ+xlGZ8uyiOp3N
7B6ynDO3pWLs1tNAC2SqTAn+RsTbZ2Co+OcyWwLbXnbfUGHbSn2L4oOwQD6P
rQZcBAsHCxouwBazQjIy09YXUtkZZLaGzhTFvJKHHP6YbH7zg67ry5z6s/x5
TQMttX+KmW7gn3BNtJDJsY3UHlN6kSw8SV63txwbw0P605bfgGEy76j5DfR2
Mjtpu6yjFMucSi6Eigfn9lb2XNMWzrLej+iproz+euV5Ta0yzZEdxoBNe4Yb
zV5YbaXLBCAOxPit4zlExOzFWKz3Px3YRFAzUNYGCtJDIgncjlqKOH1P3NFa
VbcyR4BGTX6pSvZPCSONjJ3zqA80Lk3dDGDaMp4ZpeKfF3oI/uQdLSFguPt3
q1dRHbbC8jxsRWgtR/24LRUaXVazgtCrLbIVH+a/Sn5zZP96EGgp3RxhhnOo
jOjWOX8ucBYgIbVCLC/jbxvN82B9aDq7SKpJ1B4Xkeg5i8K8BJh6L+ccE7Hq
pihMmpSHjRLBhhnFqqf5Zy44W/dDMFchuQPKJojAy3HsLX15jnczSvOurROk
geiIeOjcdw3FHcD03hQ8rcQspm7c/O5jehEG0aUIxyQT8paSLtfzoXUTiEgw
nq/ZbpKqtTRoBC5GGlXqsWdDwSwdyRsFhTmbPBagtZDEgscVpRqlLMwv/6vh
Z8OmA6lC52gX/fo8g7TEnk5cl0Yysv3hxcXB4OXxreMcRhvoEj3VtQNjsGD6
gsprEKNTIQhCTPFR9rycjXp9SsTsgj7bG/bus2ndBIo+EwoYK2R5BJJiyTZ0
ZpeHVtmGOpz5QiLKpIZk5gyLegeL4tCCWOpN5iKuiDXGeDuAUj9++w5nC1oW
6M+d13T7dOZAUpNZI+q2SnyHy7Lr5h6cYftm2hjRpSWU4ril+kB7N60Fg3T5
aJmfo5kUIB1SNhgmPrvI4Tc4mvYPDVEwGQDtp/J3Cr9c2A50U9cC2Fcj0rQF
srYsVUwpDsD0tgyQkGgWX1LpJHy8JRB3NQl1q9U0ce3quX8saXFcAyfjVroA
9QimovRVM0oeaqnkpCEdLaGeZIx7RV8j4xmfLLcnnfOhLxY6LFryXM4g/Uhz
WQ/hRjy+xRgRZpNkuQkZro8YHlwDTlj4eCbfOjYTTXCzKejdXh9Oq7fmpSqx
RjJQiTKvqZRLfKOxdfXqHy9P8tVA2m7gbejZSvFPLHeHRVSV4l3YKwwMf7Ph
aNU+EsSmnjqV41clLmd4rnaQXkGbXeOAXK0B0nR9YZh5vF+j5Z1TN/jcBUu5
oIk9tc3PLRCGXj+Z+LRddtCCRgnxf+npdaDhHUV00dMo0IzQlM2dTViVPK++
zuwCRZb+Aygj277JVjs4QwYTWHWQFF3B7FDdomRmRiEN1ugOtBNm2T8dG66u
SkDf5gzBTx9SezCh3+/Kw/v1gj9PHq0b5knXeLaFIydtfttRMar0ZmwOP9F/
h6QFtqWq/02hv3vYk7Rg9AtQRNqv5/57o6nGi/lcNHvePaKCPO1hq3FMmGkF
lecG3ctev0/8cWerpYjBaqsop+TuxZ7+9JxlDicFk9FZSdam1tjOTOWMZRcv
Of/VpiTjMoTVJ9JP/ubrZoCm82qH2IrT/fGGn0eFr0H9Xeaf9AANzOPUzwFa
jKAU0zXQCGOnT+NLKYOtJfsfbsHEbejCQaV01GeKalPlgZ5G+wGaOSw3ZpY3
/Zpnc2TolUVh5UZHEGyFJ/J0m7k6sbrA2hCEeLS0DXfTD6t18mx0k+PnE87Y
h4xAP6gv+OD9s/D2u/GP/DXuM6vajQn//K5Xvwuw56ChpaUzasg3WxS/Irie
UxsiKtmQlsTbNzsIWfVEM7yUM815OX047PXurY93XVAdItFKT90vG3jVVEzl
9GIjucKwuPDLhinnTz37l+TxLAwgeWdng8JbRCKC6OgBaNnlujVehWuT4Ace
4oCk/PuUp5Rm9NXxCltP73kWKsmZzH35BR5/v15gHjvw5nYH1qQ/eSBAB2Ze
CrNCcC9g4BnJb1a9qP39ZHrhWB4BpiL3gGFBi9G8AEuKWlrC5MT70XiiaAv1
zvNEL8oY6ZwrSysMLODQEvLyIc7vRNQbEhqKCQ1Aag8ZhX90XIRxyxul/SrF
L18kmFz550pON2Ee1vBJrOFhV3YOmOzeZgMxswuNhFlcSjE/xLr4SnbPO3f0
wmf8M/VNYaveNm/nFJW2/1I7dH8pxC/WmFC05JjUQlccd4eP5/MX7vZZrnP+
JLQCWXCOphG/PVXV9BbotbAmW+Q554g4ptri2JBTLa53Gasn833971KcsHaO
xT0WNlQ9xjG04k9hr3rd24flsitQZREIminlLbnims9UXnzG1hP5wg+A5frI
D8O0hxt4T+5KE28WhCc8oCjCj/NgQaUq/GMBEMPdupPU53JyjTXR1OlID2s0
+PvSbxbFtUGGOKBnLNLnKdCV5TmOJmlpWysZ//rzRK5kEtashTaYVrHt06Yy
D1ASQdH4cS/lBqDh1EPhrPdrdldZPwgP3t3EEP7/3CsAYzDl8jb97cCHNtOE
t1UerCes5WMbcsyYHcAox5m2hBKr54YWLNcGDyj2iDh8VfUGiAchw+G63nYr
oXuljZvSlwV0+tV06uAn/ptbO1xv4YpCQVRxIEYGDDYlOBWbGdKwnCw/Clyc
I4YXt2pcU6cIZZZgh5wzh25cdwBgQ648qEfmyWcFQLHi93v5FSJHDpPSFfHs
ioPDV59RMuxtujCnCnbWF6BlN94WOJmQLQpaktUqXcbjU+6StwFYyURh/faa
fgPIvdvavywsCI+sPJmrt2XNwTakgVWhkAaOUEW42h9FQSP7DD756Jnivd4K
JYedzyeU4ynufYgWGGuvf3TDpWYKHyyMktkNDvOGJczvL3u96jdEgsWB9kgA
t2QXUHoAl4xIgSiU5T3q7Xd/YvuZZRMVe0ngwizTdG18kPdH0uE5kyk1tl4m
Ul2q20InM/6Vkx1yQt3KPGslgc06gJNvfdiyowjueAgXlfxEvsLPZHlWfh99
bqbKIrCnyAQGHe4z9m3VGfCHDBgerU+R4IstiJ+IlrAi+RthFH9Vgv33x3+W
mBcOoJszVfXJuazBUHjpC861W40Q+mEWRaTU6UkGtTYMOsdgPKGFv/ZfH7Z/
g1GYRfdPwc8T9X6ncyUu6rK+XcZF+h6SyTxiZfLhn1ynqLHAZ8OJ6yA6vvy9
qyfytgdJUsVbFWv3xa9TppbfLwx6OGTe2If6Aifkn2Ymer6s0RQVc/Y7srFE
tsJ7cbRi2YRyKwK+JPKLx6wSpM2675O4ZeNUzWDjcNCVoxTJjVtKrijsCXW9
herIH1VI6GMWPAyIXxKK7+UNJd5WlVyaSHoNvohu2UpyogwEeH6sbOgdNDm/
i+p9nZBdzPsafON8kOjQDHTb086JXxEbM1Sg/imKsBivlu1hdEfzv+2NXJa1
fwrvtoiEgI0jW4OVu/hCza4BzXgs7C4b7h8EpM4zI7lNa+mCcUNHzSskGrZz
aQzpBJR5isWecTpX6Lj6DhJifWHTVdVpADaMWjL1VsIwQoNJGEjdxJjP4tix
44iMEfO8K2BvMAehRrPYnIUNG9wxSxKOG078Nc37Zz1/8LkjUSKziV3+wL2b
BcKf4dOh8fL3xSmy206UFvFxDBJw70KszBb31zSo7hovaJD07voz5i029WgR
8+kxPlcsiTuGUNysH9SDfKaBmGBp6fOtV3TTk3Nfp71oI8Had0uN3tlPOEpX
TxstOHvrvvj7pkKoo7kPWrT5XMWJfpRboC/Vk8E3g6MOfG1H/OrcWlqIfRVQ
OauWiKQLHNQcNsppDZ8Hz9nFlsBbq7xCC05cqvxXt+cXxqPyNgeHRm/oYA0Y
4JvCbUrRnPWLHyAtAydulygjV/P/0zsctkmbPE2J5qitBo/CuSWiuOUjxiKP
Dekj3LqvbkI7lME2Pf9UUP5zIhk5ykC9Tp7p0lyd3dvyKXR23v8QZ2y8C3IJ
eLw1GKwRMVe7P2IYeuHyoxyWTsC97gRBSIK/KFI18BHgLlDDwPRvpWkbrUt1
Eut9AFe49ioS8lnlWC7crFP0MlVypst2/aAf13XkRKGVzcSDBIq7EnIHqCjL
UHwJQOMBLU1xQTutx24+OmmHcChpMFxGgqCNkn17fTSo+gWVQ1I3cg1HL816
OOILioi6TsURWgYWacMDw1bx+y6uZ9KI8eaxhQTpboa7lrml1UCGLcGxavdS
RYxdHQedtjcBvPHRy5Jia0Z0XxorvD/8MhTmCdKdmiZOixpZ0BuhbF3GqOdx
piq7w/1cbwh/GwNogNvfWWO9pBzUCPfmFc2fCRI2pslepo6t+TdG05D6sRRs
cL0spEG3ZH86OX+U1ss4VsTc+9ojL1aA+ny9t0kioZjsHKnxNzG9KuXKJmQG
9+UzgLXegmX69P9iPNFX03dh1gnNbTOJ/V0bcb5jWAbRzwUwc7voGe9y76yJ
0wp8G+kn6giMJdihtybMZFhuG+4CQhli4i92gPFQO4FNmsz5XVvwmuh1CdWK
oQuXnjhbamld1cJjXiF8bxzN2ymwEzVEKHAQd1v6+XiiT3ZUsI0G1gcFcCjv
3nseQsEzfVgwNOmsGht1B1YRQ/aaDEbWDfU2+cVu9v+VhEEsce3OZOPf6P6n
isOzMBHkB61uo5pgJ07LpkOgbSZW9epOeKq2blybn5ftxwqdJ3CRNk6FOeqz
1Zf9/UYP6oeBTRdfcxpO1VeWKCTy7Enuwtw6Q2EyT8d0Gbk8biglDmbBjgJA
3EURyd/EsLRFgVCI7uKfCKBOP1tdSIaiUXbfEpNsOkXHxQTjuXqtUjsFN6Mq
tdtGojKQug828LXJyhOfyniPAl0V3FV0V19AaHP3NFJDcHjaC4TFFcjrEC7z
FP8u45To5oyDEpNy6uu+Ywum0lzOVSakk7QJNkyhyMk5JYWXHvvOy10oE5QY
zUf3NP2NULbsPnI5OhbuhUMlO6KdIRIZiSc/4mQoo5t0ANF+vIYN/HUHP0Nt
291+NxXkyuOiC2v0h0FWdpAQ6c/qnrJEViYZN6bE4g8ydJPud017+d7YklHG
+Mtl4+ZLcPcUunPGips6Rg3KbNkT4DJnPvIgd/i+lK+DkDzZyyw96gdPifVU
m+yiDIlp7x9EYRIOyNnBafR+2p28FLRpWHQjEe5NECnraTypno1qUs2IXZFc
UhCG5YGr5qTtLjfqyF8gNukloGxG8FUSam3lmRfXixvzS5jdw2QR4OQlJVM7
MNFs0bW+7HZ0SPm07vofVfDfCVbLpyOcEjMWF2eLjMkoPJ+QgeQPvcSfOTWS
TLs5+4+4UY3wPpviZsiff3dR63GvHoqJtQdRWnh3pIwWIs+bMqIDokuwlgKZ
r4jtvAl2mLkLIh4nEiXHRr9SzNk6iNNht0LNOMv3juxqVbfLB72/0hH7q57h
JeMm1U5+DhbVkWh4Fnl7uDPZRGlgxRKrKEOI7HLdRttiM7xq6IZnqJgA6zAq
t0z+sBqTAIrVtOaNS9rsgrJf/piaLtwTFEf4eworHR2hmw9zMrutmhB1wL/j
PRf5NOuwLgsYUgWA1H8fokOSoRqPf6GiRA9X+2g2PNUtq4OGlsh7WOv3fnkm
pnQAr7+WDKPrsZdcR3IJe6x5sfCKH6zV198gn/DEdF41i4dimgo4CsKHWeIV
iZ1Zh7LH0XHcdqlobRXg8foeDZY+/JvmMR0sRVXhVGIsWgKUZ++glvgS7mR5
VIk0hC3TDHqgLmoxMz+QvSgrmlkjDmpiPEJ8GZMYPerQosL8+dQ6Zi2qns3t
mxLHRI5V6xjxgshYDXe/HI5otIk2zdEn66rF1nxGAWO87HGEDywosyah1w3y
+slyeG06PIyCiwIjXmHlVHx5OiWlSvU7GG83qKw1yIncqqMmk8rvu38uvm62
agqhq5cw32urNscK7ZQE3XxTd0i5WwsW6FOHT2o8y+4MVT8BNQ/0z8EWP0tH
OKUH8LRi1z3pzwW5+7xGwyMxIKEgQgU2iHLR1ZJ3AAfdXPQ464ejkEzwJKF/
fR66X38w2dinHefoFEVBl7vZZROVXDJ6RtorjQNIseabytPZ2TCvcUeG4VPr
IrJ6U8O0s6jDG9TFr0sFssVQbvWzjkGTidpU2Qq9bgoua7u2fo2dU1iWY0Om
IiQYP8AiFdBj1diWpHNpmm6KDU1qqW7J/nXUcIk7a1y5h1gXVthmtdCcHdsF
CoORJ3+r4WuYhgUFfqmxDjb7JnFAqvjBGwOfyUcS4k2D3Wxbhpno1/sgOQ3A
33xZo31+cZhCAq4FZOZHOQLNptUUCcecD60UD5Sw1ltn3tvO07g2HnTzaOu+
MwQxb9liq2K8M1k/TS6sDbTs9hp33DCvReV1bkP9Jyou8FTeVyMoVkEfS5ob
Q7AG2ZtSKs7dXmyTbaOtG/4xPo82AMMd7ZHII36usk7WMRwbPacE5k/Hd/5j
QeVh3yMWmiAO7LpCFOfmSZ0BE2zUVSCUUVZ8iEBZNKhOvqjJ7TNXcVSQd8UN
Jg/37zrFfHRWpgIuxosL/Heb5Yg6E1/p/Nyo7a6KRhDSTSrR8HOygk4m6s/z
CykhxHkwFoQ35ddqNK4Z6he5gO0rlWBRYlypioL79xTU16DY+R1TcXXjRSrJ
GL25h5fXiiRfdM6yhLDpBgpsoLC0gSkMQQM3OcX+Qo3+Q/ftKoVQquKovw4R
H/y3gpSFn+VdB/OlVCIHnouEmyver0kvXGz+kWO1k6QhUiZi7kYKNEtFnPgz
cUjp4sRfpDBhdxRlI13YBSubTCgwBcDLO+QmebmC/05UNCOurnw2QWCCdHVK
H8zmZcUpb6GlOd74kvFYdlbK8ueVX/tlSEnq2f8D0BeoSiFFkPdxNKZUYhHg
HDTmYZPzam98rXSMvcNQNOM5X4W3zIBkrEbxFWUVFD0eRCEDQDuHnb+WcLLh
q57SR8bN1ItktxaUFFfBDNvqfVavZHPMgYKZp0uqrjQQawfiwQ0YDk8XZbu8
e6XG5hfMQ+ym+c7cl6RVlNcwNxo2XfltZawV9KHZJWwlpQG0Rd1ZE7CZN9UT
rj4AcfsqgNB17bQdkPD47MjeG37dAu2VB3aRHsFb302Ln2lcJWgFto41HcF+
LLhTLQPD1r9xN/x0gZVM1pD9HcjvjxqM5RuGE+bNhCFbLlFI4feTJPLPOrBq
z51rMhY36+awrdV3vXGy1Lm1hYIpzNJhGOdH364C9EsXzZgq7ZbEARK82y5+
7OfDvmXLVSryLDpEMLrTcWoK+L60CSrdRSa8OARonAaeGyEj3R0+DYzNnAXU
h7ha+EiT4iqvCaOO8UhRsoPyVVMU62cLiH/zII0GTpx3bj52UG1c2mHUl8C2
Km/V5mDR9FMhUe9sPib3StpvusxNmPgY1cMPfVcHllKn0UuB6vapmTJ10UR2
JdN54bj2zw57KZMthTVJSk+1TzGeuvPpwSjY7x5J0fFYn359OT/Ej+JVWFlT
9oodUU+QMglPqcA51psAdCvSq17P0JtDi4QY5mwrnsBUGWsyPNBvlWzTPpQ8
59PymEgk9jnFIxMLoybK9pKmfrmbTpqPtZmqLPg1Ht+6iitom+motWfKI45D
QnN59EqY2bvZm677ziIPr3TJKMnM978gSZm+B+Wm2fHIEAiS7ecnqPPjzWrp
yfCSxg8f8L2T6Vvrhwll3m791KtdMby4vy8KIS/Qd8Vm6rsb4V6Sz8R7tSzN
z8cMigNah14v8KjuoCb57XhNa2gpzQgNZTFyF6GoLbf3rYkAEzo7JnGqCaC8
pMphyWktB0nGBcbH6+4ToSAs6vNLovQ0/OiQu46pCk37+zwbovF+S7LCm9xv
twYqcoJkrdR7AfonYlAcX9kY9SSgti8peaigloNji4AwGBy6RF3YLAgJk7m6
b81V56mWkRdenbLVteGnu3YZ2IPXaTmxbiSeFZsdhYgqbx17l0iGOf58hxAp
ofByCp019F6odDjBGqpKjG0DyCtJYmfQOT14pWjDarIR4JJFxzic0GCOpa60
5bckxyT0+6fWhe+HP7c/4ReJcHWzdovqkJksh/ZPVu/Y2Yg/IMbvlQ/d94pZ
zQCreQaVwRVsuJiibVtjbLexyU2Zw8Xut+UITzrali7GpcEHAEHFEYIp20Rz
FTWZayJRJuqtlRXMdWxQ6JN7pBdqA6Mfl7zkXtOcGW/3Ocd8FNBdiMmqNrcq
B+W2xk9aspTPW/9gNaHZ4H6j0rBRkqWz7TdPEYN0CMY8qI0ABMfPo6K56Ues
JODcs6FgDHRDgypmbPNw0hhheraWEMekANcStUK++l7ptD4/hNlkJnQj44Ya
wWrA99eLWvDApGbn5CwvsJojWhtV62B8FdOEJVOFpjgtbBhk6ma8NWa8Sir6
lPvu9x8oS3VIzaK7Tb74dBYf5EAp8mqzOxVEBrKkQMcJO1l38dHDQXJpWGoB
Mg7zq1cP0HndjaQQu1E1IMVvyjatkPOVM9GpI4EosG3g50elNHEZQWkvvVEF
pr26w+pe4XlHWuyCGsnzI/VaKDV/zG2l8/7nVRiSTJSZfdCV/f6lPWZFefCi
Du0xs2E8fCG0SPVxNnuLSQYLZrQis7lGkRQYGGGL4/fbHwgnMyH8xCytFmf2
u9dYZ2fJgmErfZgeeN30EPlWHkcXT0O0KkL++RtOdDkVI4wIreZkJlnVryfl
bNDGTRSeCOpBaiAusMC730IRoy8Eq1MXo21ujOUIZKQYJcgQA5nS6byKZB51
5G+vXwr9VyNOowZYYvfR3uEn0JfTXUwSpPhtjyIMDDXTDnLX7hfD44oim4Yw
Aeb1xGw349WqSBkbL4PUuWMA3tSACabczvMj/ALn40DosGPQrh9NAtEu5mlq
x74lpmg6RwmybPiUqfhUjSudQ0vIv7gY45UIRbsXZJ8qsUju+iz77C1g1M9o
mlkJEmkIbFI4IjuFINib04ny5MtbSQu+nEqBT9X68GQPcarIKqGeJgMVV4ys
1mclw9X2J8OrE0NOblaKKAY/CAPIfUVz03tqoF1HrhoWPhijcI8FAyDKtaJk
KTIVAam268HM404fwtwO18nZpSWaEshNS+hfPQkuYicH1bfLH1cBwrEOQ35A
pIUGnAGsrATkcEeYgKaySPbWV6BAmg/4loi6ns53UkBiVaNOw9Pkj0raSbPh
vcZLbH6Io54rmM/z/fAx8QX6wbBFQ6mqiceLivVPaqEJl3PG6MhttdFH2Dm3
NJLeuGO2xq/5QmDEJI8Bve+hpyAap8L+D6JpMOmyapBNLiFj69324KPpYdBu
u7/JSWoR/guurHVf4IV9dXSmesbSg6CN4TiuSGjg24dp/0gV4VWI+KJIAnaz
3F/2E591Fz57tVdN/gJ7yV9wDWTD81kX82IUtQcHuICylF4PElkR9PAQBmsN
O9sK2yDfuZDs8WmLEe8JEMdrI5t19GFsiUyIJi5X9ZFizEmLK79JKZnnqfs7
MCzUzjWBOtnZeFvXu2Qo0D1rR/nM3FofgW0/FQzytAJtyyt5ZRztHQKIaX8u
jAgFzx4ucjeH5cFEBccXsfbC8OXFPJ4em/XF+5RoTYOERdwpwAmz2eM4PN/y
Rz2qgkuDfSCiLSOWlDxUN7UqyNAFuoxTnDZIXd9ysWB1xFl5TQzcWXnrm2Hg
fv5OzXBh2HhY+DwJ1Cv4b0JYLcDMKxhRn1e+jzGo9I1RIyBCTyYUsnyusa6V
CzKc9Yyq4gCBxMbOYKYIIyd0kHzs93KqqEl95Js7uRcragVEkWVYME2zEqU6
BRO173V/ShF1BetTITGvr0dkrMtJR0Z8Y+SqhERRil7iCIoOC2o83lwPytU0
uowJw6dFo9l02a1tcYTJZfDPdwuC5LkBuAljnKHPwMdPV4eqDdftoeqwd/ld
Ok8OoL5jz5/jKguZ4PClNSvBckfTczj4PBrxWGxoQ6t786Roy5/+JTIeFze1
GaYg0eJxc4jpUFjQuR3kc4iNWRozS21pB2jcoBGPt5ML3Mi8tIlT/dafuKYa
bICYYHaCazU6Ba7srBTuRyj791ezAcKyfI9dQVi/Oik70EesVkOmP3epLYC7
JSC4t1rL+JhmYNmcYQ5qoDop+eGBD07QJZqYb3c9EYclVhXc0Xqxi8S/IFnw
w71ya1aEC0xW5IO3prqqmyQYctewxvFXzNLt6uzG15Z8gfvRaAVunVHkp6CT
pato4JVH/lW7IPOwUHt8Le4ymICPhNB11EAot0/ycWNkXfEySM7rykpEDWlh
k9enzcU5szpDFv2Gjo32CZ+fQR1LSi6ief087RTaj5fZCiis8JYkubhPJVv8
b/mjRrIlYD+YGRnQyFu4LfSF5G6VB6tbPdcD94UJ5gc2HZKCQf/T/m/ZfqGW
ixs2JPO2vnraBOVq9kc0/DuWoYQFu2nqSqY/N7eUa6YLXnDn+skrHK4nWHyy
2pXGKsvgM7U9DEzfn/3NpUYKeZQVbsdKTe8JRF3V/hbg+nJfEqqLM4/C69vo
n1CSe3S/B2o9QY9t3GStI9cwu4vfhGfciB4Cj6w6JDFDkbQjm9QmE5+0xL1S
SQPrs0+4fx+x4asVAcE9EOYEEea4kBrBNyIUfnonUbV/VE4njwwXuOz6Ixgu
EH5a7V4nRADmrvFvWsMcAd1ckUN5//XRmhNW22/aJaeRCac3xzRGKPkoVbR2
ZdUcNYzRlbilcUoVqDX0Ln3sV0+Ugsg5n1GmJwv4abcnapH5T6xpMt6YlY97
z+42CHWTMbfW5/i64Iq9W6G4FK4gAI/y0Hx9dQYTMvJCb8IdhQAaoHZNniwn
cBgSAq+lR5q4/A7si004+8bzMlaX7HRjSkdKCIbvauEEh8FR52kSbHj0WU8D
wTjGeKpdw9WyxIBCsMBR1LLYLpdNccvUJsxMOL+phdrNTXRcs8km6QwrmSLn
NjbzpE+7GWhwD5GUpiUMf9tWGnN0NRM2uBh+gCN2f90JmkfbI3ccp5OTTstE
9iIcfpe97S9ir6ji0VdtAtwPQBBHPkcv5Ek2wigkNxfCM2qO22Enlp5vFlJt
Sfr7jQ55+GZOMARUorw7ATHQ8U2NiuNo0vzpymZklg2XjOjMrEmkMb7AUGUK
3oGsOnFP+VHO+1xyILnmHjUigARC2N9ErjClkeyqlNS/+Wd5NcrlmXrUpXDV
XutN9SWzRrP5X0bbwU4l2BTY9dRVGJmdTUl2LmO0fKDuryLnuKu+9hg3zsoU
W6jb7lu+JeRXHGpYASbKWZgIR3EddqFRT4kye2z2FeH1sf3QOK9ZSLtYCCUw
UsmzSqRSUcP4c7jr8fS+HOP8+8snctDxtzw4CrJNqP55pvcqpCftTF5M5H9O
/m1TkPSPUrw+vOsTfKC12M7eHGv2nKJzo9LmMX7HFisjdZrMyFlJ2NmiINO2
7Q+AxJwOyuoVEVYHvj8WnR7JBIw+VwIwdBLU9OJskhVUZtA5ZcoL/z7eaxa+
9/OCclDYZcBoo+n2PzrjsHhCfSYEU7cKRc284XqmMySpEtLEvtR0+lYyMp1T
bwalXbllSlH21i/NjtXTkspi6unkzFTFYrRTEbgo/XKenMFvRIG7bwi548KV
zAGTIFxMO+Wtg3ijtJSLJ+IZYdPRE2nOFAsur9yzBJ5eQml4aysvG37CtdVq
kTVH/Ts0H/rAZdvQiiscWJX3fsjq2C/iiNAgJqI/fVj1F4psFuG91ImOgns/
1cMyMN8dX18C12j8g9JczlW98Prx7OltO4+jbRJnRJcTQlfcVzYXKMTxlDMX
jUk2BnpwjziDEZeQxTpCAtoDSsZgwFK0hOenpjWwiQzMxuTs8l9ZP6B7zX32
LNA/D4RKRFHNmXbE7mFxm985sIUaaCWcA4fZ/oFOIR7v/XV2lwj7vEUwDBIV
I84C9/UGeQQ7+HskJCqem3pgIeKXYb4O1SdvkzJL+ICq61Nmr3v6jXAqMKYp
tWSX/2mOjYWJw6L+dyb7NMxAEw7quUsJ3pc15DTxbFdaKtTMDNhWRoWbB1WP
yZKxteB+m0EAhDH8K7sYapZtDCwjNaFg8lmnBdNwKQuw6dxZcN9MfrG8V48E
LnliXLDzozfULp3WM7VHI5JLS6+7socEu5YrHAg1bQzO2CHPDeEHGXP0C4ZZ
8MA2RQHHOezvpePvvUHKZzMBOkUmGTa7/57xKwUKipUhEve6UPE+PT6gOkcc
YuOsXJNJ9Sr+cRmz5qp+c0in4HXwe/E0ylJhQpEfX9fVtCF8y9xxQa4KbH+i
P0pb3BTAFHTxX5S6JmhzH61GKV44D6zLjTN17aR3mVoHVJX5MuhxyxfV+C3I
F4oaL0Sb2kYJ2szG80dBesAhyOnaZPfJNv/JoWihWrH1PxniI7ppnxO7djDb
M4niLYIVYGQKJMGVk/jYpFul238A8TP9qLEveE2j52I7ul/QKDng/LKvoi4W
yJ+fRTg4dE2HOPugHmahLmsjqQaYUMy0zBBiDw9SXONo4ezAE0OtzEHhIsoS
1OCOpvqYCfufLHWLWzonZsX1XT2EL03y/UEEVT1wfm1oX0zR5DohPWaJ4JzH
YPAurI+k6GsDcnyC3I8JZxrL9qEuPuInZiym4LZNQJWjw5cndcgpX8lKRiXd
BrempBEiPoBskR9n05UqtVm+mAURBHLFgsqoifOtA4yiSdfHWJlX+cfHpBhP
aeZJUm+GlL7KNRBJwOrt0C8reCbKUNe6iqPDOMGfeQ3D989dq+/DYB7iZ0uQ
QM4k9+MCSDfVSPt281eyjWKuXT9qd2AATr1R/c4lEGWoVrbZAVtmUrCyyKQS
bXdbyxk4gSyBAl5bvtNiOFqNski5KDXDo9nSrp6W5zda3tTqxGm4pigjN/El
hCgELi+a8JsulkhTVRh/yal+QlBQnUxT52Es6T54r/Ef3lxc1CvwWaWksJq+
RLUKYzaj+6ACMBdjhrYRhWrM9ILRLSQXIIntt7Fn3Rc6BE7ehqtEYmCKMYcJ
9TT1LH/jRUGFs3BrERAalMvpDoyNruKpjGgMSX6uL6B4Ao1TkV+2dWt7Mhod
lwhs7fIVivqq1y/nGNPVZkuRgjuiakVyb+HN1KwYAAZ2xKervAjKYGVnf/li
SBMh1HKrQZawENo3Ctd7Y458Dvn7eY1COKN1BaqvkxGcbRPCdc1FrvErr6qs
ew0UR1azvrlX8l3loWv5S+MCzIrbQSNK4vNxtEg/IunvDNIOzZHQAcyZlnck
5L0z91T969vKzoE/k3UIcsZZDaeDPur/5sgwp7NaN9OjCHxBKY6n2BNj0NGN
JaV4b8sGtGlk5re0tTIM3r8xq0OlViACH+E9owpW2BA+Zld6KH455BC68fO9
LLjz1cSUe9c71kpTeJidERBtURrjpr9v1aCZOJFEDuCC36gwgtwfOamwxyYX
/ZQa7dHieNSgemiauSQfGIWvsE0akIg/xyeimU6ZLf6zLQ/tmlMwfHmLG7QK
zFjlQtII4j/ESTS/FrgBSX+2sOrHh/Z1wAtBwp/LaSeCyyILXBdp1mza7BAz
AufwWTK1lqyQ9zowiykgc4a783WkDb1GIiChaIWBnnVwjwlxrOyokQjVmwy1
c7XSBL2+YmbRtQidaZmVEK1YLPc47hRQT5KiTrIt3afqjXS9DPe9ZunYf9Ir
ErG2rrA/cLeaydrxy7urIZ/UH6pkUnuFJJZkFd8++5CppiQiKx8MV8IwLAI/
c7+4yDdToAcdgxm2ubNVWYkeJyfADaRSnBa9iav+uY7m2pfzRoZOJBLDfT1p
41nilKP/QTB7t15VYNYuLSrvT6rdMnRzCzJUxEof2uEJ+hPhh2RetWOo5LRP
uHvPyDk1FwyeL+YaQajkVvEYYDaoER+odAS8CCFDy47QCYVgwufI+7h2TU0d
kdHTMZDJQQdiljoThvXzL+JXKSZ6ttITIGIJCyaKlz0F1Ii43J6EihcGwyTp
kaPHlTqhRr2lBOT3DpucZLPJwtjXIPrQqWGzwWeBxKtdhHL2edU3thHp4E11
KrpWLCPU538rSe81HprqUsOXZgvjVJ71+xRTUAUEkiyXYzD7DFZkKNj2qg5S
57IHce6x7oUfU1aDfgctYWW8uBsOVwjXza4X1npGWoD5oPkxW/kkI+DF4WXa
Ne+/RXh1NcO3ns2T9Bop76bHRvQlNgXWj3b7W8r5FbKzgxMi5/bHyurDraES
CVV6P1SRqaPV0jSUHmLs9auU8WV2QI5mTFI4bo53SKGRAYrMwH9SsVzdaUPU
rBQI44BeO1r2FhZ94KDEAMh9WZ9i/i/bWgnXQ1OYBnw7Ezn/xsa7YiKrUgYT
OQ0Cpqj7APVFLKtzUGlDsP9yarmtzB/78rp3v3EeTo4xMAZP3mfItCq6ew0R
3KevsItxKvqhN6g3vc5j26WpVe4pzF9ilsP+fWvA0y9VGVxmGIXLGAqyoMpn
0Lj1ZDeIbnREmmL6Nciqy7KRkgXLGZhxReJDFO7fQzX/ntGPPpLn9+l98/nT
H7LF86nn2lR2z9a/Ce62ul7av1qOBJauKnTjJ7N2Q7dvS2N5W7l0H5hoWDoK
t9VA4eW5Sh6Cpb23CZqShL6OgcP/P8k6f3SX8tSxHVIgZLoBNwD5uSdg9WZ5
GDG8sEvqod8m6MZ89jWYg78Q62HtzPyg9lx0erph//XQQ3KspcOvbi4PtXF9
nevGNVYF5qKyNZE40mXIqjDEK0dJbyw4qxbWvrNFb9IEFYWFSsayU6NYQVy2
dafiG2Wr3VAkitXZfJTBJBUMJslOxynRMtCyOAYSaZkkB1YRfeAUkZJ1WRu9
zXlL3sUuCCoFl+mV4rPfDKkLMScogrXmeiY+teuRCTuIW0vTK+tNl00bQK9X
K2yi+wpO0CH7fdCwUTJsDrged0QS/TP5l/zM7Vk2m+SItfHGIsePqF89tjUV
pRcDLdOYTdQ1lRCX8/2aTDrTTadhkK7qVU9DrujxR1xQSCHkz3qKviQgXH32
F2RmrpC+Kb5eeVqlja9HP9k80J7hYdPPAWlAZeZXo6sHwfiJL0jxkcxMwN9Z
TJYbvaRwpL761VhtfOrgME6GJvT4G1jhrIRRFoe3bMwmuLoxOR98Kg8W+U4F
mUBlDHNKUm7eH5g32lSvBaUzFAFGHFpKTsSiJn+oytuBIFS5aGnAyI1giALK
B8dptwHmGnKvxdbQBi5cf5haUm/CoqKAJnm92yVke0X2U6e64DgbMm/Cw0hX
nKSs6wRLyuINKOd4ksfDEeFId7cciWTjZBlPbKMyKiwibjqNwxMRK7jRSHRr
rybt4jYwX+Z7qxj7mAlLvwgHuNrlaAXHe5vo7g/jQgwgrRvJfu5e+PTT+Idp
wTAI3hi6HTMSumNirC+ZlwVd0a1eAF4Zb4NglsCvp8Ml6wHnwo1RaCBZP0yT
2v8v1sk2g6C1cPRNJLsZptbIydBX+/m2BhUsEQUfQUagtN/jBFTZ3Lvpw4lx
BFrz5tAbZUVWGk2fe+I8GCWqJa1fAmsevYLtfNGL5rA+8806cIOh1+OnjPGg
WUV9cLJ76ubT2dADlQ7Q+3hAxG5sjjPsX16mIW+8EO9RYm6K9KvCgVnsCI7l
QLrzc+x0U5zh3xO5rBX3L9Ipzk4kkrmV1uJPM2PnrVPltb/ye2YvWOWsmhzB
xBhkDVvHSJ+7yPAKpRQJ9VnmJUAEuZ02shy1o+MdISYil3DdVDVEztx0PdXB
ZD54tfRyUgiUyPFgyKmdBAfLoayZs5KX3TJilHd1SKlnvccMVYK78HJFQ8yz
Vi/oxadggiEsCVmj9BoZZh0vQl2dUkp8hDyWkMx7+FXKACsD+w9lB7RWoXLE
fR1RuKMZQbmBMe7FqeUKYuc1Iz8CI+vNyL2aa2gcXDR4kTprs2RAHtSMeIop
a8kjqfd57TJun9vm3PW/Rey+CDh+dvRGOceIv3VO0vnp6G/icW3dXQ6gBeKn
3MPgT/ed1ltU6WEkEmalbibXETr+7/O1U3DIWGI1I7obSnP91sACJ4zke79v
LJdksKJKCCNdSZvIUmaKl/ymNEYmqu+pdEvdhvNtxIhrBvnbXrpE6dnlu6Kh
hOqc4KYnGJc2KOSsI9pLIcb/6bmTmjRKPnNUbu4YdjP9DCxqDBz9Do1nHmuj
FySbuJaVgZK+JNHG+HncyFJaY1hdJkslrV4/acSXhszpajVZHoxrClBhbdun
73G4/foqR0xj93Cndy4Rli0ym4Ll7ZR9zJqDO/fHx68koy64PUii3W71OqF0
4jg0J21w9XKqDrIhR0RAOirYDyWYkaTRwXMJc2Ac4n4GvL+VZ4nbHwOhcbs9
g8FJx4MVqNP9OOkgO2SIKSg0i6DrdIAik+t/zmNfbvg13YE7v16Pk0u2tcXb
g3jvQD41D/h5y/YUSoWbQGjynudp3pBfRUY2w+52cinV1OV7J7TbMKga5jGQ
XTk7iLmn488UB6nF6AZRMRDrHT+KCW8XRNYkeO5YGxuvXMZBlPyXH6WUcGNO
nv1OdgpkBC9bNvWFO7w53VeTfK2YObOUrYVYL0RfxT25n/FYLMPtvwfK2+P0
Htl3S0zgulvqgnQoGq3YQ2/VWTuQoKIuyBA/O+tLOpdBtmKbDYJsEtSq9qNB
I2faBTKkTn/cXYpHiW3BBntN7l9cFGSt+aNafUGGADhWXJ5d5sQzUk/FfNWN
BVQ3Zf1kwQyoAz1coW1fXkSWP3uhZVaEAIsNmedUduc7HpJMD5tmQPBPfEWA
r0Q1GVbP1sR6Ua1fJDBORZvOzqL/lAxoPxQ0nUAMh9VCCifPvs/2h1laE3Of
ONBrjFp4UHJrKHszftbBNDIw05CBBZd1qvSrXWrInOOApNDeDn9wnnPUVyVE
o+0R9VGCoNLAPMRor+eliLPezW/B2p/86553doU/fOtbZWJo+scu+qUGTG50
BG6ETp/cr2RnTtTUWk+kJ5/o9UmZ7Sp9xvBTd+Y25Q8gXZnfKIqY3DVj/1Oi
AsUahqYhHz4HOCoysN3VDFTz7nlLhtEvi7+e61Exomq1827obIyJd6eSQ4pP
+Ov6YRcgQinGePefhmyxQCl1pI5lsklvZbfytG0wkuf7OTx5PdB03FVzH06C
mpxV8EZV+3WFzYLcyPzmSlDSwTq1Uwgf4+5+56gFHMhWdIYvnOPonDzr9yS7
Y2SdD4qg26FT8w4wIhW8oGwInIwBJzAzoG9L8EejTUf0cbipRZ8TuuhRu8uq
beCk0voBzUYwx0qXBCnKMh+oeWXKpEnowoB/W6q8DgCGGMuRXLhbVHgkdm50
BBaGfIGjx3YvazWtcqTMXRbc1nm5GYmErvJS3tTFuu2rqDM9KnBR5IbLrkoG
TUxeMDuilTZ3zOehlRk8M3gHNDpz7GV/bSwVIMI8gsMDG1i+mOhKLP8kCW1s
Z19X/WWGYAry3LqhFNqEi804MbMw/br4MKxZWhmjCTb7vwFAfSdLkHLzf3Zc
499r2lwuBN92UTDqBF2qV50AepfzAhJc4Z82hLaQKTHAmxsnrj3AUnf6lb1F
N0MHH4LqoGfjVaTAHuLUWzmN2t7bgqBIQFUPS2xnCRFTwiJp6gR8fhMIj7NT
XlsdU5WZPbPlu6F5G7JbDAe5fBJJWFGtQrxmnqjwjV4aYWH3NlUj7+Iqzmc4
p6l4ARYQJAwyot3mSt+daRX4Kzrk8nVPns+qFlhJk5C/v7TCun2ITCBqi6lq
JS56mrdzBbbroD0BLhnOXhNwNKrv01jTWDB4ZjI3as9zCeG4cGJmVkUBS686
8b1edN//y4cgmLfWmLHGQYK+9A0Y+b06iC1/4MOzphdbeQQAtBP33twZcU8e
7I6A4Fqas9U+p5dz5qo6uo6WuPh9CxjRZ4e5NW0IHvhdwlakKWJxBAY0hytd
rigIz0oav9Gq5tBbX6y/Y0gg+aMHrzTxih+72i+XBP569NcoIqYMH/iid0Dt
iTR2Fcp3LHRHVzCcsLkcRdbpQhs8YV9su1HEW0BOap1kchpd0gX8WYSlLAVu
VPSyvInzRVWOTlKhvGNakpMUNy9VXtrhZAhjKt4B3R5mZgA34D4fHgeyz50t
3iphZLOu4s52MH4zuBjNBW2adx9aAChsd4YIugz+Rh4SiqBZK2ZWtAYe97mf
tlgOCl/JipsrN5dBBAhzh4+BuWBoXFcuZ84rNSoBzzz+EKpC+YdUqeRpNt8M
sKQECOKVW6KV3qXi7nzU3+xpp7QDNHVXVXBKxN1uuW2x9LUwE2zf0YyXS192
RgDizesszYRFfMSXZMQ/g37mlglhUURB44M73xclSs1WFy5NjvuMv/0HfLjP
l/fD9p2d/wLuPcTa7D+d61HHxuOQf5/yKANMUiqkiGoosk0WxS6YmWdrX6DT
hxGJVw4qWJrqSh9BBLcEKCkRy1i4pX0SS7Ioinw5F1zPAk+nC80gLTO/X8tz
w8nPryCoG6Cdo07KzWj5XPiugyjZhCslo6KV25gzzBFE2QzuJ9f0lOXEyC+4
bWF+01USQizxwZNtTyDUcquSVuLuHd15X2ygX1uvgFkFVeIibrtyG4O7b7i4
eV+KdBneLmLMTRJFXa5cwRVmwyCEH9DrNh8PWkCbxQ+tlEsJX/r6/oP11SkD
Dr3D9Qx61GX5hsnf8PIXtYTqNeRv3jXUlkapu9FiQvLG/n2xoB0jaTVhVmwK
pTRfWsmC7PZq31UeU8KeKwpvFUMJfpf5IbGvHpOeNQHuLBRE2yehyM+go9QV
Emm6+v7aIw9Spe+B6GncHUuQizLHH+UAmegGSBsu/LKE3jGXYTSAyLCrr+7Y
EUM0vvjPQcU+tWniPAUsVC9nZgGudEShZ+M0/LVpJ/6N+KQsw9h1A38trdKw
IAV8xGKXHCQ6Mm6zUJnFaY2bO4DxSbvfS+a2Sb5b565+ZAU6oIoT9bGSlozC
+YFNW5Rqt6k30AKj0W2uOlgAZcEXyoJ3rSHyImfwhJZrTnvL4VZaXglHgo97
2W9glmwmln1RDfdmpDI7pNyCZSTRKjHhRC0gH4tFBPmrTbZPArmbydtSsXue
R8RN7NP6FPVhSNijXfseuhC2NEdRJ4skqigHb87zbpApWSm96aV5IwSy5x1c
ESDaLTLRNTQa6RBo/qTeGmlLWJ7zMg1vFqhSKuGfVoWVInDHihyw7VH+99yd
JeJJBHAc62qiOY4XaR8LT2ihxcmqqAZCf5wZQhbKP9dnk9/R3VahZuOw+GKY
Y9442R358I/0b6m5UNjlMv78RouecxcYq/1RH+KL0l0YAMDOS+AgXJ9gPnYs
2xwSEVt7QEofad0ki9koQOSQsDcO3wCX03+evxCD9ffZs9Mk4YvgQVof5qv0
+Au7cnMivDH7mpJ91C17sbjfU2rV/ORfPwRMTpfewpBkgPuEFwMYEcqvv8fd
zTv/70vF1LcpAdsTdR6zmL/cpjJRD8Tx0sct0w1DVfR9nidmHagEIdfEnf1V
VIGaJX/rp9wcUP6Bpq++NMpeXpTMMwO1pj//HCS5Oqwrem9kijXnfSWKNbCt
nkiwBN3wWzZRflxsoKw9PRTInpHwZqwLCwuHq/ah70a7GAC4sXb1Vbefhvts
xS6nkvyfxM5jbKPzrZDmYU8x2Y8uXW4mjs5u2q/vzLTZ1FVvYfKXaHGQkuJL
cwOEYyDQ8laEmnRJPupkz0aVhNKQUjIsBnEwCdjFVnlES0pR3Z3U1scGM5rx
02htVVKPrPSDc6nRuvcQ1oZf/CfBliuNWIjP71VKmLo67aNcIbAMlP2Qs+ce
DBpEQwTkZWLk3JR9xkjZpQ6xI+eaDUxCFlOzGJ6lBpqLxAQpCiJ9q1YLxvq+
Jns4SYN/WBu4kTxMio7gvU/stDLbn0LGCN9T9mjdZyQgheKw6tThOR751qIR
bzcFKr6wgsTR8sc2lbaQgO/kqhgDJS9Qkn2Jb9caEzdT3dCKMUkf1RtFjFl8
JYsrp5kYT+5YACdnEVpDvdl3MAOzp+KwWaDHcmT/LgO9MRgVtrRVBDiVmkz2
nza/EKKBKiFCSAZKr1hyo8AQTkSuUTF/MuNtno1P09639eUBrOecoZIrXWKU
xUqkAnYUkQpqoBkAzKVlP7ueu7bViL5HQqAtwyt2Dz7T5N06bUFq2V2Mo7Sk
POxOhDBNvlBklNohd4VsNeD48VZ4M+uyNkto+WJHxjOqdjf51daFPjQbwL/t
xxoIt/KjxuBIvjoKFNE+jrBiNb6RNKEg0zvemD8wPKnqmDTVLnSNu3UEtlW4
rEFlS+tT6IvSjKcKus7Ov4KiCNMJ53T5cgsMxtD2y/ht5QyteO4tewv8EZWs
Izh7ghdWABwZ/P6k4RDWSP2RRv1mZJnRiAr98qPC7cUFK7c8bUX1qzr1043y
hg5JuPsivU03kKtebjC9JytcybvgYgBhrAMMb/7048/E/K0KOyJKJaH5gLf0
12mGwKdUtAFgyD8Xf0i5e47mvobmQmapfgecZAxUELnDmMciD5C3svWA/rOU
ZeY3y+ICBvxxFBVdAQwg4xLfHnj2HiXUaj+SckBjJatQ8DbGUJFWuw3O6V6X
PQA0h3e2CqmaBpokggeSyMNPZ9RUdV9avwHWC3JwcfgJJJzl5bQgG6Eh8MEi
GeP+Eu3Am73DyWrDTvZMrU/sk4KQLHxS3HYoY15oi2Dbq/8AjByvTsJQ/tFX
cshhVnQqbNTFi2lgeFa0y2Pe+MYzyH/2Lhm8HTyTSH+OJx6/3N4hwA7ThAVR
KBkZdxnop9dd/RSspI+rgsdyFTGyszZKmzMdUiIiG5snKbC/jAa4+lyhdEgr
dEpZ9UHojApgwFDnFZ+TAY6zZt+kVM+Uqj+gwJCVDOoB52TmzSnB0dH92qCW
2pJDgVN4yS9TFb8shOzLZpRALu37L7dbP3Zcj0gVniA1+RV9UAEhqAOzcDlg
k5K2cGQM00wIiwpGW29gIGHJBP6A1zDKT+kYNkZcrKZo2ok4a158M5vzm6KQ
z10DBE7qhgDVSRQOzYG86QjO3laENECnDQCyGd0VDfFRp8AdIa+lKgDaTSxY
/zJIjV72xwJAXuAJ6LPeGvFqyiCsEqmZVGZUZyK0a43lfEwbtXZ6jIP5V6Up
gdLSLj5Fxe8ppYD+qkESpqjqjm6cIjLuN0uBRhpYS3lhlPT0rRrjpLnNS9bB
cNPWpcRDZiBoP3YaxsAoRZFVLtKNRte0wNAeN6deWm00zhmTtjU7qmIolr6Y
mhlFIUzmqRyDiw3wkOZ1e2M3UU+ggb0nrmY6nREA85TSLzxow223hYt5jf0c
5g6dofZU9HmsJn3+n+iHS/ZP3mwTjl57mgHOi5hSStPuVHmv4E341hTVZAH+
0wVh3SiTnZdMaMDSEa3liH5rMaf/Zi3m5tt+43+1rFStPjOEOBDHWPux6bHX
bSm7XnBcNEJH274XoGfWkp3QpD+bwcDyCcNpPZmSwryEU2ohdP/ccZPKODZl
owFYfeX1pQJBDtk+2siNusyA8zy6YR1Wdkax749b6JmH1GRJGM+JSLtf+q/R
qZ9Dz5UVHOnz7j5931xuR5xn+cL2paj+pJZB1P1TKBwFtflx/ieNQctZ78i9
PGllmKEobwxdGU9+CIq/0S6670HfWOwRzmZ8aBero3rfreIZEQdwGnITSB8o
gsDB9zLO7tNr2VriFQvRJD4Ew5/Nbtib6aNidJ/ht7HyGzCwKsR9+0Okv4cY
kDnqZ/YU1WUEVoKcusWfVyX2sbRxlwmGkOCYvR86uRFJVkq4ehXvSQP7bmhZ
f6W4R9UplFdyIzC+3vxx9OXjMGRzNY/nelHworSZTwuQDQpQR0bbl8na9TTS
1y9/9EtwK0yN7JJTj594txKE43gUavTTFOcuTNSdv2qCYVSRSMu+HIGF+4fi
gNZPOMY9Q81VIo5l2VrpmZBjja6GyL4Q95tbf5KD/g0a0UaMzqnmEaupSUQT
zaBfdy3G9vgNvTawo+hyFCVuEXrs37LzvRMwWhvUrGLSrbsqFsRbJdD4vtOn
SLjEW8G0UoaP/KvPMUMmEq4dlFqR94kYaZBZ1VSpJVEVShYezXKUUl2bIggl
oWgznwbnSeO0ktFT7s7NvYVkXiGF/Lp1DBIRrdCwCZal0VKi0nPtTFYogXbo
axswcjrMuF6mEH3GEwTlavIezYU9LqXmdX3CpPks8ZN9pcC7jr+FFGPF9nUz
BlNzDGxbKJc4JsknpaUhFfQocRao1HOd829wHvo1aRNAv8xrr3cdAGg+O5j5
IerJX+GGhsRr2c8ExmL9ql3QepgdIhP+95ms6W+7nO+Ll9NKH7kKL6+FJSrO
gYQAKs7Jk8mXKtmq4asPA+HVI3IRbioCUlKCA5eM6Ud3Cy2ie6qhH9nP+lcQ
P07dBxM5Z4qZJPzTq7baPpqjghycVBBFuUoH2305AAXT9lUM/wC+ouw37+kG
QrLruSLNT5ggGZ/NjHrv90SqckTC0iipW901iTuEixId/4LLs3PpRZ4GMUuk
z60TGwuDuXcjLVjDxgxc4rP9Fqg3D6eiDd40qwy/5uD63nvehTCCkRd3OdFD
naPh8AUxdlLJwOqBPqAgaDyWXLyRqcDQOQXdkvEJAxT81QONWuzjry5CvHCK
eaFpBigSCQNFJpQW2SEmt4/uwGhO8y59h2yR2+Gw6cowrM8pj1r4Dxss48VF
6dYweQPZuyvP1sqDhNu+c5sclZSKc6INYVD7Zfnar9/F7QIpgB7J75o564ud
QP+K1qhlwMY/5yZgm1djEaCp+O8i6xfZ+yDtir+nLffk9SJ7Q3WYJEnfjKpf
X8WoruSf7euAicmSkhuBXnwKvgi5Avno/mWFLUP9FcR0y91GyrIE+SEdYFYU
53wa+X0iLY9f+lqecdwV61De+wLivZDx61G0gA1OWwVMRkDGZ8kPbQiUft7P
dT1pqJDKQ0yWOKeKcwsZm3atbi676doAPEp66el3nQtzr7ltU4uVDhnGH2cE
qtX6svXTyNAjNk4zRlRgCgp7UyJdpmrC5Gofi11pfPrxfwzbBpUlS10bE/iU
RTvjFbqzBiyUzD3LrKDfe6MBxSJ+3naZGGqABplKnD7+tJ0yY1mRojB6QIu8
hSlo8WIWTYDVaFeq9a40RtAniTdzWcHtBfSB7Vza6+ORsjfZP8Ht6AjvUaZ3
eCwF7KVC52TuDeUSrP9zSMlfVNkxMsKRslpg0VmIH9k/QyJUO7Gkp5HoqvVA
loovrsqVKfRy6itIjMlbgAi+yS9P0ErzeQ60WTnm9fKC+gEkt6Mf724EfnrS
Bm+XK73zgH8e5Lf8y/aKms+0eCJTLE0/EXgbRhTCPOcbQpxESCHfRxbpJCDb
ozK9rImLDJ0kT8Z3fZUyaSIwhiU432GJLDFZqx+BoIN6N9+g0IwANzRNYJNC
PGEFa0LAuOA/gxXf7SG5h4uNc2uV9tXp3P75h4g4/QLC+FfOECviYjH8APxo
EHGH0gcEzze1EXW6tvtW91VvyRjcbssZQckH3mQUo1ueKxQxf8cADZo61icn
NttoIeI1xQe4nml0ZbOHbxGra5Nl3Zb+A3dVr+tkJEH0NNgy/5nCIx8ImLdG
7/Enudf+WFjs7r9IEL+4SApXLyGhglwrzshqjAbNA80sF4gTYqvVQYWK+0KQ
9jFPtxu9Vdv+8Fw7Blu37VBrGFepyvu7GCPzfX+SxVkt8AECdElpzIXHO65K
CXWrJSB0hKP7RL/deUyDpLfEiEoZxWhCrGa1M14rpAI2Kg06jOX4MUcc5ZK9
Qb6lLay04F51mjci5epNe1GBB3O0RY2eZuMPa4GlFhyCfqH4RKsUceJP58/X
Jp7O2zm4W3iPWsv44SucoXTFWIompJnPsTT7Vv57Wh4JijrtV7RJJR3lRK5B
azPWv+KkxB99yTBJyB8CnekhcvT43jjD0nn1RSaAN+3PhAKKVGWs7WCeaxdG
cVKSTrYWC5FL4lOyh2vw8ZSf+tsNi+PDhZEKYkUcRhL5QpHK9WuQL2yCXPeT
9zbS9pWvvjPV5UM5+IonljxdCa9FcJCiygyWqzFlSCnnJHQttvvuFzGy/x/g
fYx2P7WYA5DAxWlky8FznGARkcoYZisJyeQkz7Gy0wDMX9RDBSbRQYVwUo8x
xQKZ7SfCYyc3eleURRMwnvrvC/KiSnq3tu/v0FLcN1tLFOJVTNjIggKjPqZo
dcEbh997t4QedapmrPWrMhAmTf1+IiFP8wCjT8UzP3sZu2v9xrPLvO2hIVDq
OZRcZx/E5rFNYIrK4eXw7qdlWEDY9zd5NneTF7Ebz8pnNjMo/kPp0GR7aaOs
29pZ1JUB+2L2jCyUDu4IFo/WCIYE7/DRjNVOhm37GBufcDopazUgJumad4VJ
5PyvfG2TD8TNWmOz2HaD7zyaweZ9iwcRYeF38d21wT8JfVoSZA7F4L8KyRa6
Myz0rDwexPpVAz2sCMSmRHvwRDIeAhmiQOk5u8F0htKCAiRLl+R3hq2hSMtX
ZDAjjNeyhP/XxeAnI7FAa9XgiZ9KZmD+ROS4IbDnAH3z9R3JZctVoJTv88Jz
hIjXjM/Sf4SVXumMKnCwx86lBStxZsnJd4wdZgvsK9uW/dEenCUzAnbQtBXE
Fm2/WwsPPIlx8eTmGHWSeENiyS0HHCiP/XzWtc5OcqsL/RvlB2tzeVvtf/7m
Oua9zub30E9XPFdcpWD7OMYAGoP/0Lzbo/02B38LkOoyTMPo530N6Xo1OYPf
n82hpOeZv0SH+EVr/BzqusvqbVmk7a7N2mA6UrA2GxSnd3WCHeJPXkrOJglm
CpTgAq7YODLekDVFCwbZC18NK6Fa6IxVJHljK6fA7OLVgUrw6AycXwqw1AMq
QXDrjowQ8CdD1n5xBS7Lj3pX5Q82dLygyAbVxvhZDsV2q21G4ohYV8f6VzuQ
Py2XwAWzMI7A6pG/huL6A/zwD2SY17p4n+GYkx/aGne1BsSz/cBsNk+2AIao
snKlRUU4n27W3AOTkpVBvBK355SjEKj7oahfkDVs5EsqkN0GUGArOZCYreNv
WzMY9AlMBAEaLpaUfBpicYkj7T1jiUnIdabWSvMGtduh+i2qICpi7zNNLNhM
4XoDFRTc+Airx8RrhfkxyZzikZjXGhR1ctQTBhAX2h/bWiFN2bymjOFuICnG
tZvDVDi+7ELr2SU/nsIgKRXrMk64ingfPvLaxM4WWER7ExCpk9m8TUrFZY6k
Dajvj+Kpg8riB+pmlX7ZgZ9+vb5eyAu3ltaITjLDNAHwTeMFruYsdm7Ahsot
gDMKLBV2nb8tXjXagS6x5hP5p42L3nFPt9vKwVamTuxFzd4VTR09aX5RJfgV
rku+E0HGXH80wTi/ZzaCK7mT3SxeW/c+Meg+KV6854tqmWTECfl9WayW0RL/
8Xx6HJpOhwqlrT4qTx6bMiQpbn9+vJRgms4ELwjjjb/rHU4QGsE5vGCp9lDh
3DKOMjiV+9X1DTujwtzIbSkyGix/7mzn1Ql/kPghX5rvU7lX5aOQQaPnde/O
HaVwsXRraZNDRXr43vbniW2ll5Zxh6XvjoDcCkAGkS1WnSPALeYDKnfRPSwZ
7A9uGEznY1pQv6O/BbpIxl47TvXOEvVQ0ZP2XtCpCUNZTr2cwDNbrBRSrkq1
n8mXr00VMOAKJvbW6dJYsgrl5fDAqGRP9TRRgroKY9PLgzbmzNON6wjgm00Z
EUxFxbqSyX+fMWkYIiUCYupWlrOqSN/GyPCtNvs7AR9CdMjrz2o7BLixsBeL
voQjE8aOKC+7oYaUA/Kj/ki33148mEDskjV2tIe6vHk0Moto246bkr3GxlgJ
B18xtKE2rznP34+sEBU9DJnz08xb93TX2Cnp96XqdJVaHdk9s0x2ZSeHAD4Z
yFZTBOp5QmW7Hl6YidRhI9ibP27lM4iQHxdnhxuEsD0Lca8ZQf9f9jpsSND4
q2dK2nCinEBXTj9X9fHRCnlWjO9R3ifx/43keUn48+KzhL+8xjcQuYH3z3xY
K4xmM0Hvv/9jjnFSiVq25gM9t3pYDb9Pz2HK7Bi5G7K3VOrb7OQy6AkY1aYx
kadG8JRwK4IFR+tohKzIhWVeOIbk+itNObTFnMqXm7ipW1sHk6ca9Uv42gZL
9Z7TqIGfM47IkeGRj7sZB9AsCK+/rqkJCN+8kYsxLE5O3xOWOAvhieyoPtHN
UrdgI7MBEPHg09fFxOZX4uzd4zkMCeifzj51xCRJG3Bsln1zX5DJBv8uZLTt
zRbKGikxV8o56yQckHbKNUadBXSbMujwKdLhIQcs7XJm7fvlHIvNAULdn3cy
5rcwpECwRfNcitFOOK1uBOjj/DM96t7Q9zGc0ThB0H1uM+f/1U1wlcrDT1H8
OvGOQJ4g6WYVAHYY4MyHFCcARKg60qx8Dvth1I6LtLS8VIyj/KZ8PrIjhb1u
I1YQQ0i11FbFuXQ/xrb2FoIOrcRRw235cHLby9ZXd2P+xYiF1xfoeHjV6SOT
dnVTwEVqha5jcu2kHqSmUI+nWaJf44Sqo2AhtIzSlcvLHdGn4YON3iuN1piN
GqzV/xLJfKCC8IP0I7qJSEmyPL/x5BiN03QneXfvLUPhvz7IqM38Tj12TX1p
zlbPnLpMlmC8MAt7fKLl6YS0PHJNpbncYTIgidkUo8zhoa0w3/ScL37tGNlS
DRNOoh0icShGgjCCSfEHC6V/xzOxzB61qsIiau0nWYZE9bfmFFKvmMC9GiFq
n/gqZ75MwwQku3So6ooNvrDwkuIbbwDVDZ1+xbtkXGz/h7EbGBxCKz2oy40a
pFmUhowb1q1JaLtkewYl0rUsJmm3PQzslO4v1S8g7PRDoVRpGAlbK8HH9t5V
zUNb2tgSSiwMRQyd5VhoXOqOmpjsb10SDJY166J3LknyewLoVq3WtexmdV+o
CNx7vjgtWPQToitmjDxjdhhFlQiQI8vqTPlw05VnD945/x6d+pCg7w9TGH91
M/tH97v+faqF88oCTCqHkKy0584Ym8mYKJN4MbPXu6ZVhdWTuZBzptKjVKTv
EC7rnRIQhz3k8Zr/9wXrwpWDYLOkRUsC+p1W4YyvaMSt7CF+Sq1DhnT6eAuG
BscJFFLFZg0xAcaz4OjiU+f483EpTPwJzU1JwN74xOpdK6V858uuC0/EcUsK
SWtstR5CjPttHgYOx4zbXbn21f5KiSvgkaxDKEhXHVpRqiyEkaHvIdwU3jVl
cfP/g6c0Gs3Uo41UOyNjt6MffGx8mQ9uv/E0kYOd2vFnVrAK4ek5xQFfieiW
2K+EOzFhjXfu0OriCGprDnAOzmR+3Shd1U2KtuQQCjqW/baZ/sLaQg0o2ikU
d2Jy19AmdXj6O54hPpDqub2zuwxUjjURbRvRL06sK2tvjQkvGrCIMSwpD4/n
3YMFmMe+7f0atI1hDCE9ngF29Mb3J/DYyYXe9C517exI9fyrDqzoKcLkAZmv
FL5d6H09H9jkSFqg5ZpnJGED/cf0RFJJpPM4aXDIb+HgteQPcFvXIqZgvLCA
3Szwj/xEgMJsUKH+f/TEgwYEcBEJyoACc8lNSFTtJuG0ZUXbRFKFo6ovUZap
8mdKzufh2XaxbYqkXRUx9D3mMyoaB6Yx625IKeDqjCdN6gP+lfTYljw7ZJ1x
cyjtJkNSVPy1vQPN7+UnWEaEvKj4clBCM9FqXbPz3HqXMJZdu9eCLzMIfhQZ
ykVDpvGpJEL1JnksDnKYzezqAhQthUdNW0EsR7BDZm1fD9ETjL+aZ+Fea/IO
FdWxsMODE8a92z8QAK2NzFQyZBHyx/onm1aGKbYV1VdEG2Dit7netG6A5odZ
vIuK9MoaGaZn2PdStGaIC5dSHFaJAS5UqSp5dwn4ZMbVIb647jz9CdPX8s4v
bTy0vrzZtwA7kkwH0NAZkgIEe7Y7nDXRMT/4hG/ivjxpPhKRonFvLwsCb4FD
yGBViwDgBif9rTg30LFe+PlluDrtcqa7EBrySaNbB3wJMdaNgXwCjBNzZPgR
W5dlZ2mxV0Zgf9PsR/mRWvTrjFvyavwMQL0vqzUnccUPqLxqmnLditGgpju0
EnxkwDWeiEZyp0IeGKZz6GO0FmwZ+ovWnjcpIgDHsCxWyz9vkZGahn+DK3gH
KOnY7++5VQkVdCrs9985bnKltpVEPH94yLsrRZes3cAnqGcU+Fjvw/wpHhCD
qu//KUY0CGVlY+0dzKPVH5l6tqq5zsQYjTpU5sSDn8kRvPtBe7zVRJXvhXps
sL9cOqksGmuxofcxXRHBahLCpc27p23zKcGeHe3QN3VCpce1qF9dAR3k/qth
IeGF1kOfWKasxiGD20OOnaHl4wJPM7w+aHn9Touf7kJ5bLNRGxx7ZcEHTuvk
+VfGV/sWNWsRT2KmVKwR2ykhd7mPXLlt/KH7U72A12EjpRusAgtfAuIF24zg
aYTirD/KiF0Ua4bROeT6EwhQphUiuZForEQJTQOr8U1VHMJij+CP/0EI8boy
QbHtsBJpQnAPk7c5Zl/5AtqpGyB5g5g4zcn59TQdYR1v8hBOvV72NxQNb9bs
LLLIp5YiLvB13DZ1sFMtzbYrzz5pVCNGpTVVrExOc1sPnoHzuXjXN0Q35ZD2
szwkihI/6jWMWQl4WMr9PbVHoEhC0pCtxPQ4vCr/QxV8Ok5vKC/kuklzZhhE
C6z7CPUDSxK0f5cUFTccz5TP/PybTO85W3++7p3rooyPea7g3gof686Oh54h
5upgiCI/whdYw0RtsNecMItoAFo3j9t4mA/uZmTx4S3Zp9nvP44WcFPs79It
LJrHcDUZqt3TQhvmq5zOGWRnZzgrp8lhy9/MVFXkdtZDJsNdMzhqt2fCoa/+
Nwg498kIYUmBictVENaVFHQV2EEhAeoxUuqnCMGU+k1chGkIyN5RkNZQ2eql
UCW1Cg8NIhtIhCWIMIm6f0BgkB+/ALNMNnHVAeYekmEq21G0K+iQCQo6lDCp
nkpLpTLZDga4I/V82IT+IcIOK+iKsu8KzT9SRTthD/ETLuiT7wr6NRI7Erlm
jSDUOWXeOAB6JncAebGTZNnuh1TR8y8QiNMgo0PwkjhHle5GC/XXxvwfzs7N
mGiSB1G6azyPtiPimuvqRbVz6KhQb69IETu4I7BhzB8LN/Dm0cuwcymTpoxI
1E5SXXiH7na/35Dju3BktstDktmgZG8+bOZBYZYczS7J0HPzi5Zm1PF1/ODz
Qb8jNbCAXDPXK2jgHZTbe0IV1e8ZTrY0OWlfUd+U+HWTc+fnPsGAOu+Ev+gf
BNMOE/sMjanl+IgSBj+5Y2LU9vbNpqNU9fSaoZLgQ4oIT73NnSAoMWwV4Mms
b+AzAYVaVGWpl8LD/UJocNCfsZ2S+OfdZ+7P3THyuefrVLX/qFQNWTfNpa6/
PVKgrPZGWyou93knHXrHYWS4/vryNQlrm16jQl0Wdvm2wC89/SZEMZ7izIjL
jW6DSL17MaotEKGwxY4xXDMSlnhG2X3uGCh6cFI96nYL3cEMp8NL14bI/fj0
1JPGeER8zMZwpqw02OO3MLroalcVE997Hrf3Ka3Y4yvqecXFCvY2asJ4bBRl
rUeJp/VkYWMZPGpjEB6kpOHRcfLWMCmzT/pIDOeNGhhWGCukM8GZ0att2kxJ
u62OBOSMG21eCDvQEny8yYWF8CGqJunFxW59oDnO5EDsbJkTIgk22PJXCHfy
jfLr3PTHO0oQzM4pPbyw4mmGFBM8qoembWff+rdjQCiqEvNWL2PBZctfeCKb
kDQ1NNNYvgYS52bYH/SUXSa4mwkb6R7hM0d5TcT5y+FxPTzj1v3HizyiAjkN
t/Grz4sCBiWBfr1Osr2fndSGa0SUgTQ6XiBe1cUDWswjTpJaD/s/+HJdMlQ/
co2WqMzFLoJRoNEU0ILT4UQmwTstaqW3TmSS0kRkpy8n+7CjQWYlIA+mosPX
iU6zQq1VU8M3mHuoDgpEAAnzfVxnmiv5aL3Xcw1mxPmM7WCvb/UiTaOlbKM0
ZSJgjqNWwTJbphFC8MRIqkbxiM88ENeFTxi/I/Qv/jALnhd+FIaqC4KhqQAN
DV4lRPMg+XAqCquaacLLTbSaUQZUMOTAzoiBSBO9DU0GIxiYaIS001AiHbok
L6N0DsGB8Nqr8tFUJhjDmcfi687ow9dpzS1mZGO3pk/8K4JgvdRvwfb5a7vS
oz2OXVojfMzdfRrU9cSAxzpz1dULEKB3e5UQiX3voErfRnKVp4gEwRdbJm91
txap9UQ5ETYqJgY0RacM0EMvQ5h1DMLJZ9quyfVzmJv/RpUYR9Hla93rKPPI
iRqwseN1rtZjD3j+6josfF2AwrwhcM4imXK95D7iSn+poMjVrHEqKzK4iSf0
ixp8x42FwBq2iPGUPBsKRvgJVjdliv56WjGwz0NyJ+4pYLYkv0FpC6uAiVAl
TaXre51ack9tqAi1+OU8/b2Sbg/jBc2fhl/6NlpTNb/WzX97TVsdackKQOs0
6+cKJSqkCOSTtL/dKgg3cd8jtmId484lqpvUJCfZikcOlKxb4/pG+ihO6IeR
67VRwtU0q2fdU/xAyp+SlaoLR7ri8hqWn9GwvpBlLneuecEV1Qp6mtV/fWPT
ZlOjex7nHccT6lXbgVVFrdsF21xE9fVZ7jfsF3FkUVaDgp2KV3gHQsOR1XKE
xUgYGwZnURVRaS8TclPtV9I9NTMunbKYyKgwsOKiVpSivh4VU+lRbhqtRrt9
DhoX4X/1CYahYwkif2XwqcAUDLp/EIr3QcHEFoajZcANgnPOUzUhe4EI90yH
rXosHdafn2NkNjfCz7s+LZaHy7DjMgw0It5NguNG0eTislDbOD7SsIToarGe
TMzpb7uQJjE+FbrOxgJvv2x1SXH+A7x+XOv0Ml+SzIQyssUQS0+olL/jJA+B
U4tLltGwxneNQLbvAPeGNNSeDtk1mJJqIDHngt8eGsQ2RqCo/5WB8F/f5zMY
ueLQd0GO95jMYOQMtuqhSg5PvIvWuyjwRuEwlHN0xhBoaQcMBa3615G6BE7y
PMDooiH1OEHcO+09AsBzf7HvfPmS3qPpV0b68QZSEHOs9CJQi5j8dkuNJncS
D0ar1d5a8fnL8pUFbotfiXNgJT8zOOcWLxKgsfxa2UnbNkgVY3WM/1VtGoxz
tLdpODZQ7O1liMXOvABgEityk6L3zf+XpyhrRFbOIwTyb6XmqYwx1zp5UO6g
U5d3GrWt8+HC//+k2bDURJb0Xn1SKRJfHRaPmsduLUK+9uDqcCZlI6h+CRI6
JGcwodMK8VbCmk9di4cmdM2I1+tQcF0tc2s8okjBSqMgjuAf79i8WImeLCZ1
YOsDZfWsAzCoPMiVBFXqIMVtfs8a62+BSvgz3Pa5q7/eiVRhmyHAiodqnCj3
YiMnhoEvhVZ13B3u8CF/pRwuLYh+nJPcCZL2HRtCIQWIktR50Ql1W9y3PJBH
hWQBkKWcd3prpT9xRD9f7SvBGNf3v57DFcvOTVYcpkwhJXPQmYNf/lwS0Em/
AHUfnBl7fE2UnLChQG5/btjcYcBEmnECGaVYGwUfRNfhX7a6XIV1/Bg35cIa
/+4xBPIH73Z2Q/UcyuQa8oSVX+mvpkhnK9js0Wn5Xyo4gMM53PGnMCG1YFKP
8yLgbkyIeIn7EqjDjeWES7WkqoHiE223kfeGeeprJhIOTJrWdKjXFS63rMQ6
F1IRhjTGuubxanyHeJYARrrAicZTYKeHnIfGVQwTDjcMMpQNzMv/Y+xrXKdl
KT2KSAIXGXYlJuyfIgFP50jbFR932V1pM1DmRB9T2B5zgcicRLaNMzPqwFpa
CJvED/cqLUZZYSlEPO+6U9c0BNeS5INEz57KTLgtwxge/fJLQz+BpE+Ra4nz
KrS8NOhgJTtO/aY1+WDxGMWJEsBzKAFN6t/HJNODFb7JU9Acza51OZVRwTog
a30+0XeWmXzPY1HKhSvulp9yYEXLzF7lSKJG+C2FHiHj2/NNfaXiHX3YRkoZ
b0I79gd4eW3IGdL+7lCdit2HE2+Ea8sielYsDNRax3LQGEMnqbQSMhAtWIst
+HiNcN99/tMcw2N9KNMphx+it6kTmtg5MpkLx5B77W6uTdLZZBViw1n7/SYU
YFgJFnbouP9YqcNWI7ajt/LPNvD/wo2C+U49bupoWDh7EMCqg8nSkf9XkfF9
fjU24cy1icTqVubdRCfE1Ncc/MwQrlkrR8fxazuaMPvRA5jVdSARSJ3QQ+nW
Q/mR5UCuRNQn/lyrVQnq9tJwGyGf3jIdwj6hCQF74irBvxtGhX8qf9fQVjpd
a/tk2QIwqHWFXKmDWGy+l3hftUzcl2nYWUcAg2lXwASAXbH8qWCmimSf0Qzx
q2CMi5brOdWuL3o4O0cWSPq+zVAbetHbMq8MqLxjXEYaxBdWXykk0y0rVz0V
bV1hbE0/t3oUpNAVOz73ahm+wBOpQIgXHhV5xFSHTBAojE9CqVN6Wx5XXKme
ut95e513VvKJnQq5BxVLJJ6dJxc35+o8ITdBgirBW0l40CQQkKh+OqGr0atj
PcUVUit+RXQNy2DSbMSkROZb6WISaEDxaIj5wZTRZE4e/Es7KFpyywKeRUms
uc6rH+InY77AmIUfQcaNaaoH5Eh4U6dF2plGq5RUYQkZWVC7RiBK+MyTxjNA
M/+SEqeFlIfSbVBflRfRzmdA7QBh72bJJWBqvMB8ULLHbb6kSOAf7i8LFjxP
F3l5UoAjOXHBWkYLLO/XvKKOZ1yPOQ1U0YZvaojRYKBcMc4ErASYJtfjKgWF
f85VqE808GbHmpCKLw7j6cw4bE5N/qA/QcEE2dhXHlwwroi6gXSSlxV2rOyz
rPVax8/8CyW0uwE/4razqyzvx0vjYFlwbjP3ags57fcXvPgZHVdTj5ZmCmI3
UUx8uM/gAFuSPmm4nyzftjGOb01URtxGOuAeqhRSHBnkGSeIMUrWHLpEtvMU
YB7n6PDWWLk3Kz0mYzijhmhgiC4lPYyGXMSzX8PfrFlF85YywCP8rBGklrHk
dIIaJRjc+jio7mcL4dEZonwLMpS94VyE/6uvR/flDMbSaO+9E6UwmwzInZiG
yqtide8IUEsfdl0zeI5RhrrY1/q+l6Kqn6oZsx5VQYVQZhfylnDEZLwpxRVa
AjbUekSRIkQYhFGV3JNtnmtVqBVT9HFZaqekgPc/SVcdexOYP3/b/vOXiKxM
/MF9A9wIsi2jQD+XQU0inosThpBwCDz2fTIuRtZmWkOt6xJ5gr1XO4jH+/Ss
jwL5bUsu1W442OwdEcjiQRRKb/F6u1wpYVZrJiewzPttMFQZWXNbDFj2OQWB
7pxeCa4d53B6aILO5ddX9uP6kTp3nWzNYEEDs5xuuP0RM6Andv0eo+JunIRX
fd2I+9bXQGfGls8CHaIMRYJ7RooyvWysv5mQuKS38H490lbD6beZe7n+IAVF
EoR0QvYXextx94ooYLBgaLC914112estcGcLoDE2/3+z89J9KUyyZPdbgyBX
MLvjT+UITadm52rwbzsRiwek6NeETmqj+JJxViX90ovkOUWmcA3PcizteSOS
lLYcnE1+n4CzeLDq/BF5Jap38yqbpIj92q233FiHI4u+3xNYGidbjL7nD0i7
cq7se5qvAnLEPaS8CCjtKnSTPW6wmvSUpimyD0Cf93UcQWjHSBYPV+qhBrT7
fBlAW5Mx34DVu5UWIcZG+SuHqNECTcgQgIf9VK4pWGs0TCFvEZQpj62NTAs+
vnfeBi2b6ajF4uPUGyxWk9fqywZQ7XYoYPUYetuE2SDuyMyWuzssvTO69GyP
iHKFa5WTkhIJiI4VcOsWD3auqe9aNPz5n6NM3ouv6OWmnVR6c9F9/OLnVZrC
Q2figPJPryMo1k1OleN94KsOcgeeIDcGdjG1HcHukpCSwTWZu5h5b/W8gyqR
ZRFejpPJ/0k99UUW4rbDhmMSV18rb0wSOM2RP7MJGX26vV3J+VjrsL+X/zGl
nbR93qeUews/21I+9DNXp1e8w16byLr0h7wtDz0+yVNjaBActPo5RPHjUQ2c
B/XOmYJK6WlA0BYGUxhQVzOkOGDkYytA99nfSbA6mL5YLvJO2SaZf/xjJ2lr
Gnt/k70eil3+3ADdIZFOHvOHbuqZsU3BOmchcUJhWstCegePuj4wof8bRimW
Sfp1U+/OxuYQ7ayDaqVC7p9wx69Pe++jq3k0cKKZYnc+Gc+KdC6o9+M8RhPv
9SG7aNZ63sUtN4pRRXP5SNDy/p2bEXlTNhyd2nIzsrvL4bb/6QwjJIgZsSRQ
eH/nRIpnKTwjlS1QqpUWrJU8jE+CH17vpzF1NNbwMyYWZRAkOVpsmI2grCoj
EJKtQcGo0fgJ/SA2IgVp53Sl9nC1b9Rh/V0OUuMTrGDN+uqW/QCpv2wRypfN
RnmmGTHsQ6SauIzso6nHSK4hQVrGJBfd753UDXxbpCj+chPoLGrHTItqWRcT
tzp9i079Q8I26X8jiK1VNuDgGTd/QRJbUoKLzm07I0j2uQtoDt8S6RhXEE+z
/sqUsGL7ICVBLM/4EJyMYbjPBq7jMRm6W2tY/AKpw9whaGG4+r3vhYU9CEHc
/s7GTfFZl93fAkBJ0rh5nMBVPx9Egu8tTwO8QB/+Lnb2F0SNPjnBTIEC9M5z
OK1uJrm80CJfhGG2pm4lCY6Ws3wpR1WWH6JmGvOz5d9L+eDLD69eIi4cT97H
Goi0Sw+32T+wrUDW4biXhw9uTDQQd/jHqMoGJMxZYzJCkhnLzjU3Dnd7qxao
mAqHjTQi2AldmGv8h6uoQIGjyD6s3RCbhTF//wBMs1etAATUsRmWiWQqHmhL
VyM5HO/mTb+FKq70E34L5Ic2uMDd0U8qtpU4fY7Qv4Cf1RHk82FZnx1+KbcE
9W7yhOo58tgD32bDkghizlBAywAsTCRfaAevhJ7ly/9JKcyvnfJHRh3tfU3j
L2ijbm0LkWXGMVI3RlpMaucAt4Kg/PC9eKMx2+6+Cd6JbYDjFbJVCvX+fMPz
daC6XozDtZ4X8KtzhwPxDfx+hRVQpROQi0PHMq5unogQchaS5mcRAC0tG316
JKqMNzt+wVD9/OUdrEBU8OeUMm+6HOmNjlb80quwnJkuGXOXu6SbaP9GFds5
lXAP+pSzQ0gFR+P5IjA1zZOxRc2iDx2bGGy5ugHDmMxhuKPoHkYiHON8sl0l
KK2xmARcozQizYw42NuALUXSANB0rk4Irh6ESgLpHoOMdQpMC9/J07tgC95a
Ugu8jJLjXIJ2S/y4yrovMZcEdJczn54Y7ycK9Bw6tjhYoWguRx4u3Vhl9L12
qz0HHu1SAkWUKstfk4gtAjvPu/5eqi3JSyNByEsKaFfctd7CP575briS+Ngi
XblfnEWuJ6igjwwA0Z4949aB0emvNUHu8ikAK//F6nC+Z5uU2aTG0FSB7Ls0
62hN+I7SlwIalqx/7LGr9PCDYhM7eYdjmgm+fmq4T1UYps3+PQa6SgIxMSHQ
ovFh7P1ZSztOqa3VG11Cib6M+VTc3PwP617N8D290Rie9Jn681YL+CcTafdM
mI/7G+ozZ6m1yA2oiM60x5yYJ2Aen9RzDChYNBBI5aJASQ4P1P+v8hUYaetX
igExvikAsvyeIh30oHhDZQFAfMcEBoBUorEenkpkyyiqw4UTP0x0u2Qh+ehS
cjOcM0R/d/2mxeilRR+bYi42oROVmbYtuCzEDMpKIQrJKjpUKYmXDWZAKmY6
YkRblWV7qwk+V54IPf6RNyjL51dHyx83NNk8J/6lq8iVfjYNY0YORKm3q7qv
H4khaO+5dQNN4nubAybNvqu4Jsa+d9kDFvoROKiStlYFwqXgn0jHMrnLIMOf
WPl5hnV3l1tH+X+/spIf4Le3t2WCvvL1q+mMwSJlxN98tazZYrSW2rXk2A6Q
mJvXTPJqWF90eYWKVicUh8pUYF2NCK+WMX/BmJG9XyKRaKdTR0t29ErRR79y
kAHZvtV9AOWPRSqQGgsc0CHTuRs2ri0t2YOayz6rEa+FjkkQqVc+LSBsY60D
zN/pyp0HjALRZ86PeEJ9I8t0cjxDWSTgzOSG9YkAmrFYLt9gzuw7fdBlq+Kw
7ckmPbCpCg/1pTfxkGwUzIcHNIkmJXiiHaSKmIRSk8mW4gmuHm7OLT1JB71z
N2L0j8BfODVg1zV6zriJxHwy9r9WpSEaSovV3aeeiWhZ0u5ZDm0XeihGNxme
GRNaD1AlDdfZ/L1Lp5C42zaOR9pUERgLEeMoCxk9rBHyJG9deWkEvFF+bsb7
GK+jTJXp21Fw8mVJK+r7YQyD4SFI3tn4dZd8pGhMH5J/GuD3OV75XWKWik5A
mTlugrSzdJSrbp3PmzNjPFjSpvlUKsn1WrodHCycmSTnPXbhI1Oq+cJO05Ui
49ByijzI7peAAOZEmy8MdQ19uXsMpY5O6Lmbg43Epn+iKs8xI3QyRrWRuFnp
/dkXntPiHvVNu+DmHhlIfNr91EdZkiSDsaNSW7jEpmQedvOkwQ6mdGAiRo84
wvjWsnB0xQu/yXsxQ/qKJe4FWJ5qpsIEXTnsdzlCoHLDCJBQKsL7TqStv8eP
nAtygaWEFce51C7a+nmzrqCkZ8T3DcRCtg1qov6WxN6aBlsPnAVh0T5G+FBL
7ClOW8XcYj2V+Bq7WOKCrlS7v4iI9UkftaQo5YMGEzAxtzHgRQdxZxoZuWUb
a3J8PNe2LMLTGDC78gLv2+rXt/MLGbp8LcmsquHXA24ZrFhxNdykiq8az1Zl
Hu7ZGK/zul7tH11GZGQpmftdRNC3KhM8rJfzY+6+XR/PjF2MsXW5ho6KAVho
kS5fXRyGAbpGKijlspOcQ9/PWsGURkKc1VShSuB+eG3Vk91y7b7Ho0TmU9W5
fJeGFUZpgAHleA6hWrGpGsP5RYGai4o4x04fGZttSSZH1zC/qxbQKC8JUQUG
JKWWO+hG+YbeuRg1cvkCfnTHKSScVUvpCfjosAlTONqHApnBGVQ4PYOTy3IA
1kh93IaP2m0JNovajCNwqywnlibtEMQWQJk7/mzvA7IdoR0QojrSkwChHdV6
+nXA+HYXHKyeU+g8XbbaFeVOall4gTZz94vTGRIRuZ7lardIAwJBxAhshgqb
SuPKQbYj3QTLxu3IMOuHrVMosUljNCzg5BRsLt1yxsFRI1s3SGfLbUFL1WM5
nte+T5o1kreYjB1c/9MJDCLRswHQTXsmj0OkgInzeRSnBypZMhJc9arQa5Qn
cry4z+d2qtJmQIVfdfvimh6VbDZWGE0u4CNtnjjc5sHXs137ZW58m/jRJmcz
YYzqUr+YbnkL2aUkN5z2BDeb1KFzZx2X96JYwYxjnvM5UyxHv8Mnm3IpnMPI
Ga/4UV2lNQft3TsVQZ/ejQkFuMh4ub0ARfsJY4snPxEefzl9MvUzqiH1EFls
o/wgof4JgISK0FV/J89t6dzDjfHtoj0+K8SlGc5CFsYtrgyRo3GuJb7SEIMJ
85ZN1FFxR8JRGeRrZa60zKf7IM49mtMSBoItqEvbe6fCb+/LNR/UnBXwZHLo
1nlY4cYXMUbrIOnr97Og3zkMGSQqcvFBg8xlEdKS5TIqTh53DuUh2+JBzI8m
C+jlCqek8xdyBymRoh81FbtfwiGkiX/bbMY4Y4LjLG1b2ffFYyhzalFvotW+
llFVGcC97ZU25XPha0VtYNG3FbeuemprNC7fqvQVJobuKAC2tm+T9gVxBKex
E9ln5RI7Gpf1cqQnpxNTmL3W27ZMKfVTjc8OAhPgj76UrKVH8/ELj1dPtHsy
lhc7XFSK/dtybGXTjcrgNSxIDHyhQTOiF5DEmgQlfnHVHMewFn9KyRfO/C+a
Buc2yWCMZopyQGDpm0D+aD1NnZp/kunYdLUJTCOqMLADJbH7nhExi6jHdZCO
54avFoqOLoMXiHmyhCxKp8LUAuNca0mkZC0NVsrHVLBjiSWHeGnucJvxMeEb
sHSbKS90Kftz9sZ2gyGNFzFpy7f+Je3YKk9Y4rzWW8kSDAxljKJXxK8irqR6
2QTzWgcMF1OtybLu8Y212hC77oiqIusHCTURLq2k3lYLSxctdsqFrm6Hm093
fjNfk5eibaLS0t56EpMrBap7kvNnma7Zg9VZBewWD415Nw6eMAYWotSEOkJJ
4VXfoVYqNbliqtCOqEV85Q9E7miem/p3rrlLykLQn0n7vW6cPpTHkOFmPgi2
Q08fYkKvlqjFCgK9vL5hNfBcfRNF642dpitgSBHWYt3uMN72e4CfzQ47mpJc
/PzPyctT8898XAanrpVjk87yC7lbl7LHe/MzilhEKV9YoloqaMXMqB7dzNA1
Z8jXXwhJpDg8+VlwqRRDqSipNii4ONposcLp480Jy/gMdRij/iVCyyMGcPaf
FkY1vEs/iGhPTgEqtddTyWC++GzuCDkAp05Kf5PtveivZiiwAzm+oNu6z2U3
Zht9Gre9jLOa/iSNa+g3UsY1cMqNrYrY+aB5Wlcp6mByOJcf4shV6JmQ9Dex
GLTA+GYRmVYWXe2waw8Wr0Xrh1hT0P3D6FP0WzF2BzsbrINow8+lOVejMihF
FjFVeGqUy0b6HinpncPN7CXM5W2B/l1sFH8Gxu7zh7KN/1g6lOJmeZO0cI7O
Mx8aIoGce0+iLHOqf6rhO1ooIQLbd9SBj734lWtfSoZp/WUxD2EdoUX903zB
IBxS4NhwpH9OCNgmW/LhEga25COoW4e2lOxddsie3IiYCovJrjp6cMo2P1+j
Y8wRve50bQMRxBMJgWnEKgnkTKuRlR41zzT+o3To1utoQPo8yQWm6K+OQCL5
a3unS+lMwnJQMaD+cWCNjC6r3Ajib1GMfnKWocEgzv91wloJfqT3aDcuc+0f
HW1M+jW9FYWnnTcxfzDpIeRHMPNm5mNhsSytF5RmDF0A054SGXwIPwc/QyMV
WPUz69Z/XWRtWNtlyIw9XFaVtyPqpsF9BcetDOm1r7TQ9RmVjaUOWd41I+xI
NuQLSB93ObyZ0HsEuxNX2ILhLqyAQHqN6kw6nyyhAyk1SwYL/I9+xvKeLPld
Il3TS7cmfG1zUKQd7zdEg1n5+sfzurLN5Fjv48nG2l0+cNrBok6V0jyet950
kCQN7ngcAJk/pZOtsJw7dGT4PaBWP46YOJzUI3/MHNGAqnFt5NuKwdGpi196
gu2SH/f/MjvPRvFxkoiQh3OZSpdBN+Gp5GqcyHA0+iI8ucWyyghXq+RIf6Dd
mfH66C5nrFsxBU30jrdvtneOVGdrNoDKDlFVBKLoGKmUNuy4hNrSQcV7VsQz
PcNj61L7fMXOFUFwG54nzwpps6IV0bh6rBZtcDJxYmHO636gUWMQh3KwhOw0
qjcbjtp7RfXGSQQnWN1jWdC+XROjlTmGGLRo5cofAHG+apoTlkNdmC/2qfmA
IlF4ZiIFQHKF06Zh+Piu9muoPhYG0a3oaB1S2pngdKXghl4RThTm+8qP4d+J
bBevjXDOIAyGZhb0o0vqomunQYdv0ezXOBfu+lXUbc+RmFCS+oMFGUMqSZPt
RMjQt01Y0yrJ9y1GMV7tROVuo7w0nM+G2hzTkScT+0/KgrCnayHV9jZQNylI
6P5E+PU0UlBn5nQcIjEkZTuqr82yVUyfTCBn/isgivZkILDHYzKOiqVlo4mM
wAeLZdwTiN00xdJFC7dlB+gZNpn9l4a7aszw7n4O+ZaklzQagwipyUMxCrQF
LUSo9i9iRwk6GGI9ZEGYta/p0NEuWmqgW01c5OVAFhWlWaNhMob/hB6ihtMI
heZ44rsMB6DZkwBZGq+3i+MVh5jp/G2eQRDRaWg9zcj6pJ1OKuOYCafUQpqx
5lhyNShpdxBKxKVwuFF65ntRiMB8J0T9bqPd7OBo8Gi/HZPdf2XgnikSBStd
RU1bqFSNJiRUh19Ml71iOREXQUc3KnOPx/RwXKJusTp25xB84siKKOPQkmCM
EXRBDqdhC9mCVy/BnINkopE89ATyCfZkc9njyXvVA08KzKAUQH9Nz8+qx3Zf
GUPI+7iMJnH6IbTrN171agPoUX8GEE3M1eyv5Rh/xUficcLpwXGMtsujl81q
H6uHCgTz7z0nsbfuB1rqhrgqrk8ZrkFcOv0MNxAK42BDuzLjZlVmiRgxfugM
/gV9gcRMyS7MxkDYcDxMwdqBiBl1uYC8QRlptG/vsdZfAMz8OdALvySldO99
kMN4M8ct74aFjC3ZwMWxFMVSL140aP0W9aEuSf9FeZuyLxV/gRfTyCpSeHsU
2EAzOqFMtrP45DZTkIKn0ec6E3T32rZ7jwvxkeMZZ7345wE9CRTImWxzlldP
gd29K9W7L7JyLpFxKFpYkIQpVb2rHJOgikBQ/iq5S9l+IcpVOJc7lkyWYisY
lB+acj7bWQkOJuo4QX47xMCUxEHnolJxHoG0b8gLNYZSDvkmvSI6LGtfHJu0
0O1CXpTsb89SC0MD8KwEmPgBCtMpqXBRdC9d6MhJz48pG7nlOObOl/NgeudT
VqWDHWKQCkXRf5pcacmQ9z0QO+BxlO/ae9l2PX8w0fUGWzO9LdAtr6UpG+yj
fEBvMHMHk6sdcsreEfxpsLNRFWV3dqgXedPLZFdP9bnYw/Bi9lu5Nnlra2R4
1CHNE8oxamR5D3gd9QgPjW9l9EZj4PwV8Fo0Bt1nvZ7jujsracFlZXMm3CrD
gF5QtE/7TvP+4s7eAzxdVqvaA4DOpdOnQqiVnX3sXgI8gmAvB2HaWW99EuUo
uOk6yFuuON60FYq8HprtWEpj1dsrhWXHyiuZe8A7+k2Mq1+LS2/RinnnF5Yo
ccoiryklKUqP16d2IrDvBrfVYYd6+s9mxC+IRCpTj3SGdP89pFPSB56jN1c9
4LfdoRy58Je4tdUPeDzpIK6eWj0cR0rxVsc/FXMvm8OE1s12tk8d68Ve6n+Z
Aw32o0d17XpK0Otm19f2W2IxBzkQ1UQx5j7wPbcgRtz+tcirk7JHK7CaDTWG
KRkoUgm2Ycrhq4XRlqeVIBBNlKVVYLvoEWigcvX1dy5C3GYd6UARJCn6g31m
H9OhWHsc9W9gkI8ALexd16u0NjZ1s4InKtkJR3WDtqiUbd64aZf7wSvct43F
IiImf1Mn2RtA1Ho1+o2osejsEsdkwlvTVdDdF8NSvAR7LrsZiiqNLEo6YvYQ
i6Ff5FIPpzkQQI8OYEr3X2NGpmr+GtVRxRinhDjftzEkITKgKJK9ZhXDrzIV
ZUSfMaxNXozogdC9CzDfptw2+fvcQK3gLXBg0wW6O7eysOIJkU31EnndtBGl
h+7Co64WKkSRKhdGIfW8ESKLVfwmYtih0OUeh6BWll7KLG71vO3i7tWVWCws
1oQtpb58gyr0zGWCa/Ff/BG98KmvaK7804MNPkJ84+KU1ts0TyIV+bNHHUj2
rfThGs7R0L+k+yytCngySnFO9FNiC7wcy961b658ayiIu+YJ79EwEQX+/LwX
vXbDQHSQOCatQMa1OPIqRqQ9DQ0K4FqN2mDftXK6SJxbJIOJWdaeOBGq0SqT
yuDzn52lpo6DZExBsaUccJvfM7DGrNP99byAEbKlmMt49gbb8mpvLeeX206X
lnPptSH4xAsHotH2ekmLCiAUUvLoYxN3KC9AZpDbgLrgmkfFmYhaBGFQ3bDV
uVQhvy00S7NucP+bsDDsBTL8wLEdXuMzp1Ys+NXG5Da734Sg51zJ3IxuM4Ig
Tj9UZ5NpYVlI0xDD+4YYBtCk8jQU6E6DEiLRcsAeRQbAWO1ePNP38JtbSljh
JvmQ/FQA99zQZFfyi5G1W+iuy72fh1yN42c6q1axQXmjLxZjZ94qpzGPTIw3
gw7965U6318t9kdQomUHGYSUBfHbM8l3lg0eBFQU5wIJ9IlF3K3nFgpqsQ6S
+CMg6RPglghvxw0PL+aBvZTgd9bhBXfygxEZ+mOrqWY9jpot0NyotG3NplYS
paZco9OmTABUy/r8sdaVcP2iE9bXmD+iunflH22bHqqFMEcaWEctyC5Ngv1X
RW/rry/W+6M2XKI7BUD8NY3zQmMxX+5V5f+FaSD28Wo9sLrjk2Ezy3hcC4LN
aqE3Z/a0L90yCmgTL+5hn6N/X9TTJqnCmrbgyU+ICrtFxICMGDXowcfPtaEw
CYBiWrtcqRJJHVNoSOELSIHgc0oohtn26wTVrBiJ7Gl9+PDGtSuSKEfpuM6K
AeaQcpMS9s3HNBO5xElJYb+BfrDtxRwtEEMjByRBIjOljTaDvBypd7yhyHU5
duz3JQX5LpsVXAa2ZLCntFNJlzUcVmXYsksC5Ihv8ztx4cWFl3YI4zeHOOlN
/odgeS1modLJht1jw+ECy561Dr+z5tTjpjf02WBnSQ48vzkZwkCbVNMp4L0I
fxqBPzfIZbQWBoJZeNAh7bWqPsQ7GUjluX8rlRYDz8/iqUmhsx6Zrze1VP9+
aguNbHkxmrqtBtIGJtXe6S+EN6QZHpzwE1Uv/N29c4VKbIpcAVkIIcnr3QFk
CV1BPDFik7K5oGxPTVQaXS0Egdy7s/0m785Zfg9KvYWqWkU+Zzp+uMOgn9L+
jQW376pZ1Fk0Ve+knaBAVNXE9iXIhYLJubpOYQjU+0yclk6nUkNv3JLHWO/e
dq0UQxjU00td08hIxhpREtehXXLMrJljKq1DE66EjixQzkAykRKeuIkrr6TZ
mCpSm+w3FyMLwM413VXhup/ar1htHTemIJM2qwXaMY/y2Auev4GZ7wl5HNXb
mkjpHo6wrfnMcPMQg35qCWUnomzp58lOumXfE6HiC4pUfx9iXvjcDyvp7wGc
1TtMbxsc2AUlet+R6xSb5/6kkEs93GrVB8WWe0L7yLCk8oA7Ptm+qUCOvYLF
8z2JjWzVH23+08ibTq/UoSvyvdz9RaZET2DSxHq7H0UAHxUrv9ZeEt73GpDA
3D14KM/A+skWlmnD+GdQoAQQuctTgSgYzmPzYkzhJmdIWUpuS/wJae10uoJv
lHRjiyr7iupKcttu8Ywt+wEK9x5upB9Lbg47BPduYPk/T6KE0p9qggjtCGcn
33EBhLRvgSx6kajqTNksjWG431ldOKJ4RRcgG72ks4EPrOo9Eh7QPxTEkDRD
rHh+Vlknd3hN4wdFxL3a6+VM/TQRbranMdzbzcMVJHmDmdByidBOPLimdXlj
6/K/7n+ophoQKGiFrdqlrvHDM/AGA6iif7Hjxf6fk3iO/lr3XBG4lDyj8bDe
GVZVRRCCqQ4IFqK2GDNzsp2mQnxiLXVWlF6FkQ6KrxNhicpow3hXj3nXawF6
YS3+1y0JvpZPI/Jd/vrMclHXHDBN9ZHs9ARDFtVShCl5NYRWFwPMgc6dOQ/Y
IX5mqj68iFP+VBfnh31+BdmDn2JKECwvVkOE5P5IfwEzEmtm2NkVtg8RYFT9
sK0Pl/Yo//4jYDL+2wR+rn9wzrJGcYHcNZdJlmuwMW+8UaQZOU6Neb0/m0Sw
zvZrtwJVC+2qhW2qpX6Z8FPziaikNTEZnYTp0DugJTCpSabkCIDOAxP9fUAb
k3fepEl7HazAAic/HkVva3DEAM01weVC6/A2m3UaIEPlXF8V9Q3lLmT6/Ef1
3fUrBDSTwguePwRhj4CzNA0MGtFpOdPPgMlzH8NPEfsW2HtB2JOFlLFhDZ0n
IdqlSYWJx3OAr+I7J/HRyBGlDTBw7Z9SEgjG1SC9PYuP6ggwJx31i7VhXBVw
Yks5mdNXfgdBughO/OeLOIfKAP00R12dkd/Wekdti9VtuBjlObHCZ9UxRIO/
vKBKkQIEIWOGK6JFu7GhZhlHlOghfLkipuitbCzI2mtZAjrBA4p80niF0EXW
ok6OCfSsSqQNANUP2aSY/ilRphOBwAQRWm6lYjLlUB1cNF4ykZSM1Sk12b+M
Z8tQtlg50LyE47I2IAeQpu2vAVoXMPQl8ljt7Jn/udODV86HgN4gZ6N1PfVw
5XnVJnSVWetDVoKuZ+LOjyx+1Zb7bgYWSJs2E+F7dmgSPpFcf0NI1CaIMY84
EW5ejmiwMByid3ljJGSnARQqQmBUVG8/D0nkQtckzq3IYZ4q0WMoBZi+q724
4xldLU/m1d+GdYsN//BiWWY2Zcs400graj5nD/5tb2qmQ1ZAgXEdECjRvP56
zpiW76nh8ymt55bAlhSPShjff2d0pHjJdazJBe38NwTUOjmtuxyeBAjduMct
QJQnNG5aOBVUd+LLEf3rC9JgKejsSfdmJNzcesA1FNed6vJIv8C74gx6PEY4
POeD9FPVujmXKHatMvwFmf01lVYp0XPQhKptKVSM9+ndXZWihzNoyAew/WaT
7zgYGrIZRHK35gGxFOYtJAH/y7rvKStnFI/hAFYUxAiYMGYdNvwFWMVVVeSj
PWIDvoVerWp4mPwaYQWiO7Uj0nKEggiHkWLstGwBp/pNg2HfMxBBc6/VO5N/
fXhNXsJNAGxxDNNO1uoFWivNBefVNpiIccCTAP/Bv5Ekzu3u9+nJS/y+5n1d
PZsvxCpU2KtwGNMWDXx5G1BjfQ+WaZ0Wn5p/DLL25fxPzQSBU5/7kmGpEG4K
qFrBiQdaJa7qBmjwxcY19eZITO49QJrJePIb5JNHh9lBmik2r5nw/eBGhv/W
xqa9lKko97bUP711Oo9fQnKwL/M/18WmjYqK5YHHUhGxWrHuPwdrVe9t4QFQ
nuwEB5HZx7uboGYJvYzx+IyhNGQMcE3Xz4e5U+WzZuwmLhz/o+XRSiXcibzd
3J/alJVfLAmaRYtCxQZ+Wp6SW/a4DW8cAgp3N4Yvtv3K9BvuMZnwVYDUaOZO
j8CQgB3bb6XMiBiru105P7e4wRJjXpZeHxjYA602DAQM8UiD2Ed0V2NkdKxi
uPmFDEBO7PRMcBiH3KStVME6XMsXUGkuxmpIC4ta7QA9Q8lNwx6Xa5I6Fi/7
NJLOr7JSC+QciW9ltRMAjFcX/gtN0tYCa1cBXSOg8HG+5NL3MoDCFozVN+B3
TUepJwX8KnxXOUEQatPuzuqXhMkLx8bdOszcAW37QV24I/8Sh/UQ9sN63s2+
IDO5GsTuUaitBWrKOdPM+ROahblbtdfJOO6NWMzrqzj/i/JJu6X6trVsnh3D
lpANCuQ0icr9egZKnxLfXjpeT7ioK+oNQjhGTTOxsZbnfXRiv88gGq5Tkvdp
kDLfVYj+49wOmGklxe7B33jTjumHDWfI7Jj4O3aHz36zYqaVhDDSkOB0yORo
ouxXTV0SG+p744Bn+AUxgi/Q66KnGKN+NLa248lr5rN/BE4nhhtYhsmpHqVx
FFzA08/0bg270BhEkEXbhOcPZ3VdQVc4Ki+tuaS3B4D2E+hjbnmPyotGLGFQ
R3k1KgRnRQ/bhjgyyhkq0GuqGmUB+F+y8VyZoQyqJR5CLMaVCXdHQLzXmbU4
xMhNtEodSt+huyITi7EgJbrCFA2rrKiB8ZwDIWbtw2eiCem0N2cm4SYraxWo
40XgRibecGQFprRgGU6sHMo7AwLIwR16/em7VhtieZOTvKMyiFRCDsdqyfNZ
kh85WbC5J9wyM8Dc0mxTnLoTdlSnEKVQ6/S7Bj83+1VjZ6YDz9A1fbGvwmhy
d53FnflsdxsCcOA6HNUpdO1nAlV6/YecPeb9j+GtrCtzGHPgvQxRmNvobrhR
8kAXM3CJv1FvyIh4o/oNpB9LuxHxlwxIFSnqCgygBXf14ZvCQl4flv9WXc38
2xkS1Rfc5pZhwJmKCkMl2Ykz28mXwSO367Rp/pPWUPB9uroFWQ+1dA+qVedk
8/TL8gmf3aWQlW/5vq507tjK7apQrwHDjfCZ1/ERinkcrd1tkM99NgCJ9LYQ
CuPEWeR9nHjMxUrp6mErPOo6/nLsm9QFgK/ppGJNdaGw1WFV3DinZfdNlkuO
gpVrRxiDgSVMzYEvcoj8BneM9QXjarp7whHq5hStCKxeHpK2cK11AZl1KPtL
W+Qfg4O+oMdA48Jz1Y/eTmTTSo806+TqwZL9QCIPC4ILWuBbeOv+dFfO0FhD
elfs1ygCk9XiC+rCpRRsFz18HDzO7d5GbYGXZC7473BLq71z5lexOh/KdF0w
hT+aQCVQ2NnuvNv8TuGjVaYlAcppwvYmFRXMPKUUG2MfT7KD23zMemQozdXK
pDzzPcQRSR96J4OkjatEAt0tcJ0GKZIwBAmKBGJrB6kHsB3vRPqVcImOkV16
hMYQSvDEoKMUs5V3wYGy+xPrX9XXQPxoCDOWBdpq6pJQVhOw8KUMPLMph83r
/2DzFRfXS0ZzWPvRP9MtQ+jVNtizRceNfmfQCxHw0t5P+m13aza158fe40Ov
QVW5NE14pVg93yXZXrv2qiHyoZxf0q8an19fz1BMfWbYiWnP2zhsjY/n3PkX
OPp79IjyqBZo84JUuYQCOXtfYeusMmTp1LJ3hVAXvTQqvQrw6pHivSqoFHLi
yaDyny1EpsmDkbVc3gybse9eKkbO2Dg7oefO/9ccRhA9t5hvsqI7u+46H7Uc
H4XtWJdiSRh/O81G4jGUfqG/oBCBMenoMaI1wA4SP6WZYY/MutDIFyKZlR+y
lD8yAc36NvBmEBfPDl6dm5tSHtVYJLI/brTQDjpr6xHenMbq8JjCCWdRYOwC
XeFBazxsZ9sDia0Bskv2He9X0B9eHl6oyAJ7mNylSsCXliUZIeYEwIBQaS7Q
xPeCl+/mkZzdi+/hDbqsEyM4RwISms1x53vrWzXBgVpW3SSzPPRhaedef25w
awqC1v4ORPdwWSZwnd4yojnwbeXBm2vv4dwc49MQ9VDsFbsgsS8holJjdC0y
eXey0Qr+wN5uxdmsSdXFPrFd+AreaBEiSsUabtSSgb9rn2EfxXbCJnGVBwlT
E4W1mx+N2S+KB8iX6qawUtaIG77LAuG9NkNFCa84bydJ1Y5tDbWaxM74R2jc
SJM7uzI3I9evSBCLwRURFLT590oQIPgR53GShEr62nMa/FaN8Hh6jJs2MQew
4MmmUMPE0k1XPaSbSH3AZmEBc9d7yszIg2bCooJPWphTzrOkxyqPoFRfryyh
vbJWm4Qo/UAOPsFLYs0ib3Z9eFwdMZxTKsJlI2Jrl2rw5EIfFdJtb4I2z6Bc
SsCE4ZXU5TVn4yB3tlKkqzJmc5EXitc18mJmMBpMHgDFgnAvLOrOb3qaoqZm
rei8A4sDB7Du+1rpXC+mjXaaTLwux9LZAAGnMYjx8mAUkxIYH59XQOE/MAdh
YnjqsQtf7ncA5cinCvoLy13czsS3SdYY/tePUBhOCOakP1ePeW9j2Yl0R/Ay
XnaVE93K2BNRfEr5nfC7Fwb3b9oV+WtcjTWc9IMrPXPhnIZS/0fpvstpYNoh
YHOuCb43mS0iWMdKYst+n+HtTLgUgBIHa9fFxu0EVD0A2Io97wK4yahCnxdJ
woG2SWteei86NJUP4nzbhsOT6D+0MSIQHdevKh6luEuJX82lD8MMATy+oU+A
Rzp2iuHTE14fn+seney0rEW7Jw16yq5PjA/BR/079uhNDgHmunaUIx3RtuJ5
9LCGr8IOX8YDcKOjeXIji613vSSevFRcfxHU+P8CDVv+J7A2ZIQ4Re+/PmaK
p/nTm0WX9OzWitqxnkpiSCnF4X+s2YdE3AZ+S8wPBX9t7lbBXYXcKqAGTokf
gijASfg+XgjXLSddnmycMNP4UvG0pJbSi0aVsxFL6ekeoH6wSNiF5yiRYqi4
uJ/fpAu1rTu7pQSPP1AAwdrpyf4g++AJaJbgUJofUf9Mp+WYt62e9HpTXdy7
0Js7PSNWGApM34M3YfkZ+jlQ7iYEYeSMqg98OmdWgHgOevB9l8oZ8bNdN2vW
RhMky54NmDuT/147P6MoZAnbNL48t8BlpjcMPuGlW1eq+GyvR2ehGBukL5wd
XhxvoRmIE/u7UP524qcUlQoGTzjbTloWEPbeeIf/ITq3Aakzv2WO0+BsVVFi
4niL7bXNF1ibUoYQ/QCzQDg00PqehCNU/hDisPXVRIyKKeOJSYWNNUybz3m4
JgpaT9phgJuLDA8v5F0Z+N2RFF1lqP1kcvy8RbKNV90zjTEmXRByGjgjt9nj
0hD9bPKQarU59KSok2JN7gsy1u8lDjvmJ6ote/AoISjJRqlbJS87Z3gmACiT
U51zVL0204NZQu5FGr5Jut3QfO9caltehVrrk27aJge6zY/iXzVczoEjM8IX
HrSupiRqngx/znHc/au/Q+/tnIy9yOq+wlQI40qN63cwZV43MtWfF1ymABCi
rQg3BiXekVOZ4i2zvHZjtQeEQ+fx19TuFu6TictkbQJ9gTpBH5szDgGY5VSX
G1nTKL+8uQhoGroslc9949oUN6DiQb5tJBMigbmruSP8PgeXMjsEdi7JJrAx
8jvwTJ9wzWKATLQgarGZPVvSQwbohM3BIsmq5KVYchcd+D+fvNGqS3XwaBKT
EldXkJXHTdm8LIkkdjWHCFtZp/QPjScjH5kEtG24UtymkeYYnzFyGytKIW5H
wI5W6DoTkFBAhJ5MeqecZ1f1gtL1hInjbtM8unCKDzKIeXxYRNmnEqBBrO8j
wBVvIW7LN6SH1LkuvxGfJW5qn9UiJRNtTy2BTstam+cNAHzCo1XJ2R6/bg5V
UPdy98h76JfkzeYHdF6xBBMQcSz7coWjFALMGWszO8gYrCASi4AdGM2iscQh
TKp/bsAWk0y7RaEkRg48S/mGMasCRO/GJWGIBJmefe+o3Y3dgPLLAjnnpNJf
IiLmRPjjhPJgq653LMbmA7nweKBGUPMhEA21OiVSNkZfTwgenW6kr3Ku5KZ4
Y9EFLYS9Edg9UiSRtwCyHi/lfdwolWzKK3hI+eL0Lby4fIRMRtn0/IfKBYyo
pv6781o/yxD8IN04/Q+w66gf4IJ+eUYHCTDhP7TOMO7N6nEqFltKymUKXwex
yQSZURYBQmaK9t6c3RmszgtSVptYh7nLIfhQzcnxA7HApC6f0vrw5DykBF2u
k8ylwEMcOO8/UQ3JexU/zJG8YF/Dy74pyYj2Qj5v9TVdgwhAu7PLrg02a/Gr
XLxpv0senONIBVsXj3XGggCwlKDjFCkASUJSL7UC1UR87ZFNCOTLwVDKcSxV
SlMUfUJthnpniuM2LzsKOq3L31LDEJjl6XGT9xxlTp1/XY+selMwN+JgMShc
6bWQ8sNJ9FwEP+aONXXwl0C+chx7vDe3dFLAOeg8BOsVubrt4YilYG8Q4ayg
Jr6GFI7153ZpM9QyKh3J60qKD1ebu3z9bp10B9obfNnDAG/Jg0u3NSCxhvpV
56tY1TXu7r8vDI4lVEruMxUmLAgDjBqIRpfzZ8D6kyJ/RHfhRWZA+FlP0vcZ
sigUpJjeUOGNCCY/g6w9cCvMMdf8p06s4LxHDmVs3QmTOYGRM9zk+TQWvpdZ
Nmid3tkoZgwvTjZnTt50qJ3N2sA6vB4xoX2uTl7OAYaikrrTkoSuoQw0RULi
51IIHIefU34VuTN8NUITKpYj8L85eHbaCSW4+sao/8nbxI/DWH3uK4BSfxRu
Djpw833GJEQQGRqklH4I+asRDoK0SGxXmYCEjyJ2AAePZtsrrL19ZKhNvqVC
rBpJ/N9M1YsExhVPKnEb+ggqWhijUk4jN1XymvN+wWP05Gqzlf/35WjP2iFi
zrptGavkhWa0kUB7C2TMa660R0XngvSKsdHxMY0FQmcNK/qIiYnYaY4Y0pVG
83HB21sUzfeGYE4CaLPboJWf8B2BH/pVD1ovst9ElPxlzeA1QAeqT3flDY1Y
PzsdkukC1Ze511O9I3/rr9ZD5mtgLXFgsiYLc3UKwiOqIofOr9ZPsbxwc/Kh
O7xpQhxLPtZ4pusVyUOCUkTBVSpAfCw3cye210Uon1RHMnGMopdLoZoQS2Mz
RyUK5ZzWwtSeGg5cPlvPxEOFd8asOswDJ7G4i8b/F4BMYi0AJuvWLD9Nil1V
XGSjK4f1k+hKv/NGcgWGFwInxd1PUUG8c4L52m+0dRHOvP7i3DNfP6R7gaqH
1ifADC71dvIB6EARsenl3jn/DxzMImt6XlUlxeX/oFWgHvhUZKS901Dmj6WO
4CfMH+DhQCc/1KLPgxqJe/NhLUyrQiA2dyDp1jXVhuIO+KgOiOcOCYXLBuml
0C3rLoqTTwO5luzYgueQFjHFIaoJHfiAl1e606G7UDscMG7ZC2JAqlbxdQR9
H22DxoTf7+90x/Q1p4Tv4f8Q7AakpOy7QPyY/9b3S9JEXXyfocb/7beJ4yhU
LPcODag4lHc5db/RI7vUwym5gl3PomGGbFH6JCcFsc3zZQQTtjtfK98rG8mh
G/byt3QDG5bCcjI+DnQ4K+ubWRwWjJHLr4AlnWWEX+aP2xw3bzCgbsC+2BvY
84+q46WcTsCYAhjCC/koP0lnYn8W7d6zkCmqXlNBqSy1GZZbQqzV9YPO3ZBw
nKVz6QHvopqHJeRNtm+MFuZzU97PaADG+/a7JZQOujipHXoJuajIIARwfGXZ
+/AgukFzZr4Rd7fDnHUQBSJZGXqhTygKwrqmf7wRUJHe5NNu8RvbY3lQbW2C
+ERcCG0ACi3iw6L7+MifHUTsGYuFi5He0eVlhpdTFgLCeMmTT1FNNr2xMKZY
MztgyJSnfop4UUmYrZ+mbYBqZa4hRMSD3CoF6b06UliDgPCbcFRcXk1OXroy
m8D8/KnI7LbHNom7HBLGZznkttluDygWZOpdXR06JEOoi/IVujsK8M1yF9pQ
iYbFnlWQ4e6ji8xzL/Zuuj6fv2MTTprUKg1bXm4rHfL1Semdz7o3BPcEWHzb
muwUkEWPRWFxNEJbBhm2rpp28ch7m8yzgl9vDAY7Sc0aS4IRtmqJc3GvR6SG
bq9YRh3oNyQOEtnfcbOol/VvwJuxw2PcLSj7VgXjGI9+fA+C0HMJNQr6yDSj
AVtjCxjzKwEnYG/B5FuT3U+YlnvddhQsd0n+owqSOk8nrt6QJBurjaOXcN8l
JhSKpcJyl5E31Iyr+5dNKg8XAFM96S8ODzAaZ89n1PAqtKTaoDevOjIaNNJI
ENhykADTgPzYh/MKoqZ8cLmpRuwwDexzKeAoKV3DcJnBvgE30+Fkz+m4phRT
wTN+r2J8Sv/Bf9dvyUVES0ISXSMJefrQmhehhJ8HeeMwBQYd69/1phZj0pFs
CxRxyCRtBpPyDPfYb/Tr8uUkYWhHYhi92NknAqH+R1bhhIySZYqMqmx99xcF
PI0Eh8plYK8V8WNlG7TmELueHMrpWFJAZCixFq5VfKt832XgH1ws4eLn8Du5
Q9oG9+eyVzC7Ra8wPCoJUlW4F91w4NsJsZm/AMJvD0Tn29xt4mUaWca82nA7
PLgqsxzF6RsXxGc4IE3tDOlSSelNxq0jGwq2Wo+wD+3oFn0thULY0h67oU5U
h7uIxKvLqDeTOixuZD4eDWySUY21ZY7FIq2whVxOw+T3ohRN410Xal7eGwDd
tTvr6pCDJO7bH/+8vI7q4SMDS/GwDtwOwPzSQJ1EAsWiUArzt7LoSY3KzZ27
i05pG6OiHa2jgesDGv6MlrfsbyKx37LU4MBSmu0SWlFoZgDqtHz+N/rVKItO
hvBSZW1OfPb6Q3LiONLAJVGVKmzza85L0tDdgcpKD/e8GquSJ0awEyBLnlFq
WF8o1+N19ENPFalYCzVNtZJQDhzSj3RcgyKxuza3DXkCbvSZ4qhfDI0HK2ij
PTWnr7pxHAI5GIFtSuyDVEergjSFlLdmzy4W801Q/6gLOPWp8hraMRFkUkcM
ElL5XZXrIZCl3EW/xxkgKjQXb3JOlChhAfoTZy1WYPXuIDva/rnPN31bZHqu
Sw8p0NJBCOfxA035OA7WPq6mEmcZA942+ORZtYXlhUGLkrXitxnPEyT3lR9Z
Oxtyl0a6+n12D7glYaQOJs8uaoY/wexoDOj/bvRn/IH77TLPVBYjJOCkAQxC
etRoggBBtdknFctX32M0hdEGyel6ALjtCLYDLPniljT0mNng24t+CErgMh4W
Rkf+60zwcZ3ua5pTgu2X0TgKIhNZLVVcMEfnpiF7x6gm7fixPWEbPJh2Ln0y
4VafgeRRGo/cMM1MMAwS7csejKJBIt8MIpACF6DReDTx2BiiEXkHlgrNbV8y
P+1tVCVCZserrjRstH8cDZnYEkH9QAidEolkFTjHnBiAUFvi/v1h9NDLlh31
ErYl+oZLkU0tdTnfBQ/xkBNnIkk1hh/jvZTGUlakzhaXKJTn+63oVEM0sY79
2Wi6JC+AlkFw7D1dVH/B571BGvHU1eyGxzVB8ZKhbC/yfNA+ajjGmEnr7/qD
1KfwzL5Yb6sP1iUNBDjhgoWd06RKtfKW/WErvjfhWwMcQHkuNco50Wye0cDd
rJkjKNPTecHMeEpsusOsH/cQMf5Ym2vJid+pHiTlWvqT8Xn9NBXjcnCBs5+i
rKK+xzRnlimgqWRctGFqgjKVxmwSFQTFfddrT3x/1VjQtkz5Ror69V3DryRV
qHoekZ8VK1oDWciEbzYrhssu7AymvKZvJ7uACqSzZ6G0XN9D/W2raHzosiHQ
8B3CkOipNlZ8MCZSnh9NBFGlfAbsPpVaRqtcUrnxvq0j0LargQ9Tia+xtjie
SFa+OJTng3oTT09uokmbz9zQ6GbMjvvVqE2loXnx2Y8dLHrqTqukucvvboHZ
2bQe+/0SBUEt6+8eHZjBuhpPFat4Eoz16EJa0fa9kF94f5j4yPphb8uLVhCl
//5vRn2yfLAyvwqq6BjPm3JctcNsrVMhTmKR7u9MSOtVdDdlbhhGhvqNYdqE
IKFN1KZ0xW6uNhS8u7zaKNnKXEEzpojZkn0fnua7s2Z8e2jaeM6Cc8eld5MI
IPKN2PslxE6lYMIPTcvCzzHn2Xh8q7OYOCBzk1WIsnRMN9uoFfrz84w6UrmH
xqVByQaNgdCpZlrlTD8ilWoaL8eDJe2COAhIXPhN47wK8in5ZfW7uDDsTOfC
GNxCMD+BrDymI+hxvWVrnwgXjGF2fBGhaHkvipfbSO5fgns6H+IckgcfM19x
zRKExoHwCSjY+dfiDgmUKjtnebJ5ANjfK4sk8DSfL2EDnsiSQI4beqxBJKe+
6migkOI4qfnWAj0fUkGnwEDt6SZU6V7+9/27wP9M1YQQ3V+SCCm9l4z1K7Ny
QN/ZHl1Jg3X5lHzQn/FwSdFfAR+LiyoVNbKNyOH474FZlRHJZHfLr6FpOCyf
3BErFc77jl7D2rogeIEQ0gv9LB7FSaFZepDtp3YvKB2DG/sSFhoLlxjUGsxT
pZFnt2GwPI3YB0vcwaxc8F3n95gcHyd+2NvDy91b+JkzdFGPWXTlKGen8Bfy
QFrRvq+6YzH1ljj3JpQC8IxCIp4kCAOFORJpC7Leo1Dlt8TpM9NlHRKFsmAf
iMUvkXVjK/C9iDXSA8qVrH9y8zEOWmhlUxtUfekxKx8iDvnbOkRstgIZq5ZK
Vm68OLskYLIDQVoidavBFX6fD75NENHhYm5MiWCeiIc2e/1GqUSJvOrHxWrd
5mcJ2y2ckWXdp0cBvAIywGoNdUaoRjifwEw8kUBHYrXoeJAN+f748Lws6V6s
wrc6NXNSmU3aVnm67clidIfcGUHYzYtpso6TQ1s/RpEkVE9bapVdQvvxi6tL
hh5rJiLdkOOVGeTsJryK2mqf02KJYOK3ueXAnFbEOXakvOOfPQoE7X5lQMUk
oukNVp5Fb3S189RJwKkQElhFTkbPky4+W3/SK0KD482nLUxm5hOi49DW9aob
0/noaEgY4wG+GPCgs1fA+rhCDtpHVDnDQdniXY+h/pX9uhYZjiHnt5jTagpJ
OnFCgwyaCwP7Hq+2ej5YcZzghiCpCt+mdwlNnDW/lKeGI9Ztw0PbaxYzxAnT
fXK/ZIzTdDAhvr++TEOb690D4KEo9HPmyBY0bPQAOh5Py1u5nUiiIqCxIzoF
G3zisJwlrwyHtsJWJ0kErscLX5gauhukb1YEF8lt+nfy4NDQqWqyW2+WC4AX
PeuNoLajEIp/PvW0Chi9dWR9iix4oQ5staTOhtvgR88zyLplTtaSfI9F0J2K
DEZo+arSyxhY6KGbx98e21kV+DO2WjvfVv6IJRHgwQjPII4hJz+CwWO1O/sy
090eqmWHbMrs72FjA47iWz7H8mcDdQxXnu+cLOajUYkEtcbmrlxWo/vqlJMt
WzB7e3XeJkS/Agn2wUBPrl+m0sD2PSBVSob2LDbscOnMIhG2zEIxCKR4Alfd
gBaCPBcm9IJXYp5KalK6iOpW6eSFe9pcNJtR7igrtx7MKhdyt/a9rt7f/WeF
1jYLPENnN20fLP7XQ3omhK/hf0XMofzs2pbiW85FMZ/xDBkpD48W4bBA0Y2k
uAkLoSvdUmYYV8hJVKsaJHPXUyIsFkj0FvTdD7D8OuiOAQ4uUiCaq4nMhr2G
Tpm53l9FZx32u9rtNBCu/oIpIjlVZqc3EXxIyJTSXIaCd5xFHKBksRj3q96k
p1wDp0ffgPeGoKt+sUjpiF+XkBrwuTaO0olO+Q4f+Lkr9ZPbBxX4EGx3AZnZ
ASyNIO8SMV0Qn78T+8MNOQLWrJKKPPqsHkeE94Ojf6vC3ukw/S1PzJFbluz1
XXzAkBMh37Ifj9luOxsboPHZsZEaTBd9fSVuhqvqPZ7IRCcrEY62h3ZDojSz
2n1Ymy0GX5deQA6Wkddeuf8YXbvIsCoP7yNXcg/NosfRhwvtX1ZSgkBm4FJV
z00ULPJFlaR34yf7x37G423HC0KX74EqsQ2X4S4pluFFZ3lyQFqleXcp2ThQ
xpZuLoSl7ENIlCtQm//2Lr13YqINHdJRMUSfO2MiBd30IkN9NxHQZnCfJVho
RwmajNuH58YZCz8wXZJpEtjDqSHz/BPdkAIqoPNrLqSNBGRmbcKD5lWQ0odG
DcBVGg56rC+/EOLQPiVtYMYH+8qgByjBX8ifvELshR36M4kvbuXou1mNvKWb
sc+NJ2VZXCL0BWEOwFoxp1ZcT1rbM3xuFcYr/8vt3MsRnSUWOnw7Z8Ohjkeb
vN7UjfbaAmIcHpi/Z67m1nRcLLNM3qSOyyGoYTxIgS4yB83eCZ9jk3LNpjKY
05H7KzZW6I8j7cnefV5sqHPUXgHGQ5ErAkABCe6K7Vwji9ymG1tNxxnWT6h4
GGSIvIPrJ4a2ALv3tA4UnRqvWoc/qXv0YqDMldXgr5j+MdlpZJ03XXku9WOl
3/lrAasf8HshxBVwgkFFkvbVCrvAWMMYRHMEAN3niicbLifoSxJiTKAW4eLu
xqB356ujBAOgK0KGUD/78g95yfA0GVh3Z8PkgFhJa+YuXLxFiKTT3PuQmNVO
3kmXGXZcnvF00Bt+gnjv5jlCQi+TdH5xFVfXM6d/QBwIHklMDZ+ARvifsYAB
TG5j+ZmjW0EkEdD45LsK83PHCz6F8dDBmYAQ3RKIlEAKT2Xx/wVgIoTkbfrJ
Gok1mOAMYcZ51ZYj1bHOYkQiCT2lMnUhZDpkI58jODlLGtG5cw4zGde5Yv1g
tn4Q/TD6o947c3oIZ+/T5GryjxMc8xuPtN1tY8y80mzx3kmW9Sf/rXCqFx+i
1JfWkv43h5vYNhACz/RtXIxeEce95W6Sf5yAq3H4AzC5DWe72lguqPX8J8c7
C3vopbFmupNE9rz7/hAYSsGAZzHxdWmqXVp9JhpGOkoNeNJGOyP7GoErDzaK
XaCSOEprqiYdhUkZgGp8tkgBelqHdqTa62zpFtMTDoNtnJ/HgatYmncI+EhG
Xv1ZvKQnO2NaBvX2JYzhRmto94j+o7xGT8r7Zck6/CD9x1kwUsb1aA9iwgmI
jYZYSWQWzlE0iVakZCqkn4KCLLT+7MRJgOS0qQGinGxDmASf2+a8/LLMF+HG
6WDQec+zKaQ9JrO11T72QP8nCStOJ3tEFnARaiFRfF4BuXIKP7n9IkwRvKfv
MAO2MUMIwLIY5C2OKwaVGkdoZ09Nrpqob6c1y2ugwpr3fpdjqrjGR3JT6Esj
80WaJoF4jcZ9R+mWTgonDNEqys6JFmLXU8lZQEfTt8nTSyMvlK0s/BdWQsRQ
oHk4/UuZ8h0nQx9HuMy/GmCAC9m4ExDBVK6NevmFdMGE0QK/ESr/HsC4oz4A
FWNyQJ944I5rLlAMkzLn+k8+ZvfmgXE5lnWlK3BfT5Ko1xwkcfRJhWnSboqn
4/QGPhEWItLQ9BzBdVA+ikxYHDOr4o1oGPGCDncOhPkZ4n1ruLypKfDFPwqx
l0gMFfDJy3oexXZ1/FJHyBJGFIN0drdzhucG93ZR7uJjhMhhHNjRdNY6Afl1
SUpHl7dWKpnQ8bJ+mV2SG4hGt0z7wZ1/kbao6VhoZg/1pyihbsBm2btzySZY
LaW8hqfYaoL8R1YHuQA5rZYOVhQWQrZucWt1S4NF/aOO3OEtpdITL4xGI/+L
2oKam/iw1r3uMjs3ZZdGcTmxppXYYOzxftu2iS98FRHzrQrc9MNgeT6SakSP
QxIysJi/8If6PLi/W0oE7uvnB3hl3rnFEdb9gkcGfqcBtXwAP2tezf/NlQZf
jp74AAXD7NM/9QpWbHMVhu+Ej/lNGxInjAvUH4zzU7YEVuIQiWyA0uS49LZ+
hy0a2YJFaHL/qQiKeC8tDGWFsSpKQ8YR7Zg5oVM/yjvQHN2QqzsrGZFQGtcW
IQ3t+wG4pl1w531JqDreFudExm/aStBzB8TdhbR4V72zKCFY5WsEdPNsFsbx
ZX3edNzJZnL9mUx9m6KYMNyeT9P07kElew3ej0aSQ9gEmWlXuUuRy6bTs/P6
t2jFOWTPcuuA7znDE9iuZDA+ZY189vVHnz8OemRZLqsGoJSPnu0SF3UUTxXz
7O6xVGCLaEOq7x4eRKkhC3uOs5fbdphXMDQmp0bJR8SUq8DbrSzCr23NSUX1
wlSqn2V3yM6t5vYwwkWO5IkbpqL8dCFh5TQ/CqV72iclW3iQfo52bjnnKSpo
uYqT9kZc/goBw2Ujz021HDRDlrJy4u8CfK/pUSt4eHeKrY92oSIi4RqsCRYe
ePatX0w7fFVc0pAr+E2tUgf2qIJDAOBAvLUdl7AJj6WNU0vjpVDErYgeoGtL
j4LX+ezGeMzc+k2xYrDWlctNRkPyOzNFReTTA4cAajVvd9L86VygFU0OwXvc
ftPh39bG+4ltBthDKEaqg4aIS7HK9cF/2/rXDroa/LD6Rke4A2FhGtMby8o4
vnAK3mXF9hpFDTszbR7oKbKXqR72dESoOnlmx9R1x2sW6olu99HSMM8SV92B
vKLhyZaocIvJ5kLcoJCqWQSPUZv5KHOR3fuAxa0AhRH70Ml2djjBuJlvD+VT
+9RlBnR8zpcC1aBh+ZpN6f823lc74GVgfGkZZzJbM6+C6m1UGF0N1me9Ibhn
7pqIiI97W8hG8iJpOUfuuQs2YqSaoMIHSNc81+oww0LyOtUiwfpaRob5Ai4W
UKhnavH5GiQJ3YzeOz4RKoWcuG/VrExfWtaEbbu6Nuuu2r9bfDOqi0R3jKrA
edA05Hm5aIz1PI8HVnOJb201C4tBIUs/aCSjLd5tk1iPBywaWOEdSeqJVlTh
xLPsr+PNwSMynLM8KWRmHmN+qCimGnyCbfJ/d35cI5zEyPfNpvQpIulftxlV
ht/RieFepI1V433cvESYsjo1t8r7xLWpE7ixJ7fvr1bZY658zUrWsdYCB1xD
Jfjfdxz0X+nZTskVtb/SL69SdzLbr7Bzt0LtbJCavlQ4zqSTK5M6ZTAdZzME
z6zASa/VV0UXov9bqAqoLRZmHact67gv4F8dt6u63xQkRJijALDCj9qsKu4T
XHCFmU3P6hdwZ7niXASBy2ET+h/ZI/WosOy/H8qbVmsm9xXcC1B+OXF4g4C5
c7RtvqHCOXTqM/rwigQbOyGY83Al0VWjw0dMZprW2XGRLZ8LkkcKXg2hG7mT
UxZGpNG2DCDkzr/9L7K6mtB6LiZxDkkjJ167QkVaog+J5bO951YWIE1/QnV1
QmD6MpqBbOkNSJT7aiRvLYqJjYbfbN3ctXGl/f2Pb6UcruUYpCjOQytYSwWh
fz2vFOw1p06uSjocvy7oyb1jeSjAgVppPp9LkZ1rFQRr9khMerk1vNc7XheI
+Qk8gKZf7UIbtXwDSFylQeMP9nfwLJcf/VmD0lLjidd/6sNbzhZ9F84cPNHl
yT7e/qDfCzaR50MhJtsDETGAuEfVDFwkZSwA3l1rFAxEwpXN3i+Y4pQw4iTD
313Ow20x7oWC/pJEJdid1UNcw2U/CmipxQztIagZWS7XPiOijg3fkLq62xVx
fFO64gbmttYrPDmtuRokXwvWtiH22HU5KLvkikeUqDy/2VJiYjRRjIeW7zgc
CXQZSRMimppAvGN/tpCKsnJhHQbyT4gpX6pJ/1OI24k8Y7C16H+5YAJ1KH+S
DmSxF1kYoWn0/pKDxi2/zB/9ShFlbjG5bfdMqQQgstRukElpuBtYTZZs1ec9
C/ehp8oACuYkjgB5a4DaxG99SdPszJcgG2BonrJ0jye86sP/OvRVX5DiNxd7
sIUKhQ8qhAOYh3MHdt7fNfxvfWULFH8mJwgACTdoOsY9L9+k0kawbtwQO0Ev
ykNL/t/xQfygwaT967yb30A6HcSkMwtuk79+d5Lb/UEVaWse4W4EoCXnyN9U
B4yyTvx545jhmrKGPdtbDFBc31IZ4xDMYoafP294bJIcJefGRHDkiZQXKirf
CO21TBuCRjRhbPmL5WHxk71cFczYNoh+8CGiyjOOtg55SuoKIva5/Y8E9F9/
8dNA9E49zpyz5eOzRYDMM6nPGTDCCizqckCjZxmp7yHp2crrLEpgPJoVG8vl
ackuzCKQMof27c2oVgofDRjEEX6ytbYmwc0LAzhXWGlPTu/jYdVeuZ0NNFeE
1xp75k0Hd1QaZ1thQLPQXUzTWbBFLrFkpCjcyKD7dCIgdk4hZPxHXottXxF/
7Gh79I2zOj33dXvZd2ooJW1dacTGidQhLCq38R2tzdbML8fozV6scc/sXEr+
1RSC29uJa2LeVOz22tK3jNh7Jc9p6maK+ifvbZ4IFU+2SVFZDoc8r3apovX4
+u1oFrLeTbvEPhC8NdyX7OwpS/0LZnXT0vJE0b+oSU4EdHywb4k2vs4H6XB7
Td+T0Q8iXrue5HcnP3cLhVuKcyEMstUXPgONGva5z0KLWh6gOUhV7UHMAvL/
T5T2zfYHAdUEKYC6j4FO5L4r0nOwm7ss4f1gvqggkDcd3fr6TKJV4vmUUGpS
xgLMHfaAfcBbX/YDP4eNomavwgXqwW+qw5xg//B6Aoc/2AaCqehJNsBcu+NY
8uCLLmhuPa0+aofE2CmXAuIrdITQIGak1H1fw7eedlHjwJcK5P/2wQv9+I08
NVDz3TezYtuGIywjFaJ4Z2oPWfMUrz5KR8dBoY7JGEvidbcAR1dv/XSn+gDX
J55yXmDlezybVfsCHUon1gV12qCnd3jXzIESP/JD0PJQahOrS91idrcyA0pt
4fPKTentK79YGSa1pDu24s4xe0LH8XlyTq3bNwgV0upuBhkKVZbqtn9S2WXk
u06s5wwCwlsCVD1ORQEHB4LiSukUbRl514oVEgeSrNCw4uxkmw+8JUQmqPcU
IY+uR/gBF34dzoJvOuNdmP2Z/jMo7r26d7xtT9x6fY0tgiW7bUP3dMRr7EoH
ZRYRCrAfca5ma19aZcI4Pco4k8uubxTQwNTLDFoyWrKFWIUXC4JRAvCFz5Se
IPQijBIfhtWFydp2zT0PykK7z6Z08GkYqpj56u+b0apqVB+PrJIPDtHrsiIm
M2vXmFQWwx54YMnrY4fOIDQYVsOJMsxsMqMGHPYo1zlWNuqhJrbv4TZofQbw
g0fW8aiF0qrs209pwFtz71vNz+lajojvOicsRPVkvgSpEc5imNnxTeXB0Sit
AD4Pd42xqPFWyG5uYcfl5Ie5sz4mywrR6YWv8T0nVXk4F+scoNybBn6zA3Dl
JB5naZ7bpM8WdCKQ/Ispx5Qi5hYjCsGxzz+zuId7NUDRiDJNcwCo4rf0D4jd
Zv3S3M1cu5lJ8+cmxNhLW2pzTgNitagMxxxdu0Ho1rSigGFt47lXRqfNCpUk
vIpijAtjZnSGmWk3GEq6HgmG0vt6tMJmlhfLBpjy9ABmNJ6ViU7MDryVrXzK
xqOVoZkQCWTLG/1b6bY/N8VJ4OF4krFx/08s8ef/vdxKWMToX2J+viyMBlMc
GaB58VtnMD1gDXuh0t6HOp+OGA4iHl7rPF5yAR16rx9JvnutvUCZNOc3EjpN
BW8waaQtvurZnt7xsgMksj4a5PJ5oRUlBX1Ka7FaC4wscaokre4ZyG5ryCdS
jAZMc2g1Qc5swdX/kigQlqdbbOdKyweWYowZJl/lwXN1CLgMV2mnECAu/EOs
v56c5SQQjOOw2tfkkLS3/n7ra/1ckLIqhg2TKNlap04syWb2I+TuD+dBdOxQ
oCt1+eLPLJgkxS5hdv3RH3CFDeCUoEyo9GFpzGLkZ6G5OeDD6VXiewbB3Av2
RkhxCoAz4G/Vf/1eban00QRN8CwGHyLOcGYJn/f1wY/fbSuMtNXfBZIxkw/q
wzBJvM/1dGkT9lDJzFLK0TWyTuTiDFvOqUkj37OXRgxNZXXzlxDbyAqyxNOR
P00plr+nLpR8ylr5BfQWUhhpd0qIC6kp6hPwktqG9OzdXSbGzXVl3QhvmNmP
N/DYfLVIza4QPYP/RDSCeJx28tdaMzzkq558DxtvXIXXCaSg5A8+g8ZlxJxj
I/vKKm+DlalOmvcTO00o9+danlSguB5hzdD6N05dbGnbOvv+dAjqCC4zBxUH
DBs1fwh7VmZsQ0OL4MdaQcRmJxjo6rRwwIxz6ChmjZ0Y8o0BqU5wj2/7gHBF
Q94cNRK5Sk6n3A92AKcG98tquaEYS7LL7C/aW0fs6lv2FOA8Ot5W968rhCn5
wvZFnNY7IFIBOlFt2sUKVfaBuIANJ+ou53C/u44e34h5tQhM++55oshJoYCd
g0GS8rtuHLGtsdrE+u+t6XwjbDa5HZCDYbM0i4ZcroDIofAFMvGM/rCHSQKZ
1cpDDP1qIHcHYNKglFPXnXoHi7Q8+ldVjNUbbgFs4x2t1XSJ7elTg0j2/Dsi
/0UJmW4rCIhSoJNw4bWsbdJpL0yKrzIjMsDHrtwtUJk24/a4keab6C0Ws7SI
s8LFUh3Tr7dZY+7a3BwnR+NQ1qRb8a4+riMCZP+Uk3E/0FGD14FK2n+wOAON
JsfLHl9x7WXcuC++mzShuglLTLZVT4mNCeGdXD2l3IXcdkZ0uV4yOlk8trmD
5z4DrZmOeHKidwP1Ze9wW+bX+YXJz1Z8Xvdbtn+DjIbGkHdvjqez7RhWYKdz
riojOjbA4DJfA1AkTgVb35Tchp9IGyjsgBbcmCRodfIS/myysdwdlvC8MlU5
8viqNBmBbIOGan/d+1ssK4b1PDuvzNSb4F9GuYAk1RU0n4ygBjQbUSddJpCx
C0qltSeUuQZOoWqNvWHmQpFyhN7fYT9i/p5dF9/GmLUqZhovX9YN1uWPUoVF
4/Fl0alaFIRPHDbNvLMKHuHILTw2YT+m7I662YH8GaLUDp+hOVQUszi7+7Br
xhKvd9M2SRd+8d1vr2oSIa0hlWRYcUY3Q9q+bB58AlUOWQDyRa2O24dwMW/Q
Ck9pIfJDgc9VYLCwVXS1ap5GRuaKjGoNwXnCDbPqJBUfyLO8o3vaAJgYgght
CWOG/ZWXBIRPUf0xEoTynqqT9ibE/UWVOAlU6GjmRkPN2O7j2jMZBmpyNq9p
0csSLjgw+Ncfw3WVKdBRj/+pp1rmKdZt/mgBkDFbk53sRAxqxgv39d0mlKEM
/+E28jEGqgUwS0dAd1gHvtOEpC3G9jT6Hd3dv3yqXEREbBvCDrJkWV9I02J9
K2LYNU5m6VvQ5VxQ1xxjToPlVX2WgRn1+nSsKHxYetsxk9y5UeesVhB/IfzB
13IvfQS25f3x0WHp/PFp3Z/Aol95bwNY80aMbBY1fN4E4hiJUc4Ui0vAMwyW
6WOeOV5zPNsSo1LxX990+gFcIOerKnKZgPDDp3+6GS6Jy8jiHmXXbIr69w1Y
C0ijrbjDxRwtIj5TCCrpcdMFuc+G3O3uzBsSDjWUSHBQI5t1XyUsMaPHHi+6
YicfZj9j7o2jmdeL8FSQ01emJA/R8RsxZYG0dd91Oq3OZr73Taox7inpSqaE
df35s9qdt1U3t9yswqeUmtd8DhQeIb91Ay+UdMO4Lvm4Q7tB0Ga+Scifara5
tCOP58zigX0ExZ06bnEewKey2PRL8EZUBSdFK/4dn9GiZHi8cukU3galC31+
V5oPPCaTr0CRZ4KFS8yjzsnDQ3pDjVXjF+vDWFWLFCrjzerrS+bdCD0k0O3e
PavTfRGl7jdViRXB215jrvL0C5dGDGsFKPQy8r84lWZagPRINJZJVgM9yeSL
RLkdE/GI6NFpMKJaCd6UcDptoDRyJJHVPdcKu++Vi5+d5iDNq0Ty+UNkAP1c
BZtUJr6Dj9IAi8glpGuPTuqm8KkPm+YRh7vLjgoK9F3u9N9p/ovD7ckdlUoy
Ft0lII0oi7cV6h9jdvR3Cqqz2IHlZUNkZegoBqH6WlosktSKOB3jLEEkxCGf
/r9Uaqxuc162m9z7/UKWv2FhZ6FcTg+aZWRkCbEmQiDk64Si7+VavKBJBKV+
eoFbd44Y/MBEwNLKqJPrPNrcuyIZXquB9bmW3WzmEhlu9f8vjVWTD2YbLF0E
EKEnFNWmCK06vkbkS7X0Fu+5YCsNFYlEcWHYjj1WOeCX1WvjvXts5hWr6d7L
DgpdwrHhlbCs6sYZLzNil2T6p49i72SFZZp8zLZn+1HCmbmRU8lXCaOxvaJ9
gq9UQ7hcXhrHbQafydXxSK6ZTalMOCvhB9xXgEKshQXD62sQmFJwZ9LjHcex
S2O7CNoZpPS7NNRzazMg3nbZc65S4SJaBJfjrkemvNP06zS1vDuaes6FYnFx
0mYR6fuWmKKesucqgtcTFWV+03NymkUV9KHYMFE1MtDeF30papQk3WIlgmmY
3EgzRxfmt0hAz5yjAC8BJSyYEuVWnH6GLoa90gtJ5/eWHJ/fhOXmewHs3eGI
K/9VB1BGPwkTVrZoACZ25/Nt2+gpBC+Womdj6K9J13XHX6NOL00BKICg9TRR
V0rfvLY9n62rwUdyHVIkRzPg+WW/y9mw93C3U96XA2sLOL3HA28XGQ11V860
yEJ1a8Z+I03eV2HKtaBr6RS0D0gy/+kGs+y2zwNyPd6cMOtPI6Mohm1Az4kB
7JYbvRehhKPsD3smcQ8Fwl+d4B5NN4O4+UE6Z6QOvjJ/CG9pGkYTj2TR9Yp/
GJQbIokBWU9zP94eKce24abLJuSvf7DE8RJVZOb0OMAX+OsreLnZ5cLZmMu1
MWhcyBm32vf3Tnt8uZNhemNyQ4PWeeyQEtp1aaLhBJDPuiQEIGVKAXCHkH1K
h83vEcziB1rwbL6X+593Ygj1AD1kmOyuxOL9OzAky4X+V7PfOlynRSDe+P3Z
nIDvKjTMPcDQH5gmeXEysFqzEBm5MpdJIb50J00eyrN8vFAzA6MH51MWY0T1
JTsqwpItFCYXJSCbpz74HTnSAVdHcbVNRGsJYqJWns3jXQMpUN14bHRql6D6
zySC6srDw4Yiftm7AyCA77cDmPwZlyUg4XDYBNgHgTl3GrEA0RFG+cvBtIj8
OMFaU7CtsnQ4Qrmas1OI0+w0SyHbjkWW+X7FXnQdJEh1tHZsYZVbjIpGT2CR
BVGoX5UPgNVuX8KK5oJyoJJ3sYbJ4l4O/giYuQ/xSisnr5WjGX6yckgRxYwv
ACMKQRzNIFW4ZhgEcKq4D/7qzcjrDqNBxlF7THvlZhY2f5qbT2/UxcMvbItc
XnvjG5YgQv2Rf43oaRGhXoEVwLFQjQewYOWMfwwRfaolIu1iWQ2B1XcbqINl
RvZf6HBNs7Hh10LSB+/pVtm+2HqyB1hB6uUI1y89Xebbtq5zBvprdfN78yMh
iJeYEmwVtkpSNMmMtbOzmrOvOnerDtoshQ9EGR8idfiDsGo7eMDaNHJLHMDu
fzxJX+XBI/eiSVOguRGvc+CIEXWaR5YVA9DcqbShVuVdxVRPWYyeSpYTd9eQ
SRo4yQtE6hJNcldn83flMyo/+ZqWPncsZqS8td8Pbx/CHMaMOa9T2U0Hxnxq
WzYw5puIa2A6N5566kzBGFpPcc15Fa9VSonDvJDXxZcgpF2zXfRFiVqXcJsY
BrkisNi5ezfsowyc6G7LqY2EqAuUZekc8554Y3Y6Yt+FKGKAg40pALQSvhgi
3Jz3wblDe1+3/xbmq9L1wBLPMvYvNq7rcfNXjjPROo5ipn9mqQpjd7AYY0Bk
qnu48J5UgN6CtSYNeV3tNxmZPEEd8bi3YSvmum6YGcLFqH7H2jNTiw01WpbU
jcorEXfPRJrGN5IZgRgUCi9H0+octxL81X7e5+mo6rjP/klzh+rA6FWWQFyt
ipIKYNtxXWznS/TzkY/SWztUsh6n7oRECby3ZoJEWnp+p8kO7cqs8p2VA22Y
vc8k6kzPknBrM2SlmklfTZRa7lvZzJup6CY/F2+smcj3s5UUfcjyqqB0+tgr
1ZZBBOeMTIITTwsdniRqpPIjuZV51h8YZtxNxIWUE8PUZ5HQIVk3CjoJVrvm
q/vBNAJX/8T+2pzv6wiXtdxytifR4lTKuBtNDJ/xynGPJeYlLHfrnbh3Xrl2
BCTbsgriFbYeGBwMoP8gdDt1RXcWO4ZBjXY96vGNCR/Eid/dCosZleoIB9W+
BK1zAY7UQ9G9HFUGZGrcbiYo9YLn0U/kGIA3YMRfm+dsqrkzevjMbnyd9ocz
zE7CL75qjVcVfkRY8uEqj22KzYNL8XwDKZ5gBo2wKNlnM5P4y5+IaWzPV6KF
4ihjjH/63LneJMqOHdRhBR9pkYdAaWAk/4uO36cOr0zp+iSej181LmiT7W07
4n2F0qOEP5a94Xp/jX1AtUGxcRnk819g6gOmbZbOcA6uu2p8MGGsJYj7jQNx
wZ9TJi3ikIIVVuZ/svBPACKHl0E/0st6itopL5WBW49OBk4tVJLrIlpSdGn/
B/6cevw0g/0X/XwhlPcUtI6pfDCxcuXHS/6SylU1wmHikzi2nxCDhWhjjcw6
RwKDK/cXbE4DPsFGFmVXYwtwYsU6Rqb8hMN3d1rDyQreDmjth4Kq8GBTpxuf
yB7qXszjDcaVJNMhnMkN2r8cIcvT2xDEJsbp8A3KM/mvJ1uyQCAScgHtcg04
sAh74OhOK9SnBIPkRKl0HRCt50VFsqmuyB/CB72NDg+1jDdN6lXQFt2kVvMM
BsFSkO+0ACgbgmQpegzOrZlMexp2CM0oCaWVihCsLMZDyGruv+Mzg+x0XNIm
WapZTLC5BWe3zUxAuieWTG1J19q+8cvfY9WYk3lMXM9Vb88BYfsZH0PryhCB
SKEYw3xJDmGEXXSipdaz/ZNS9WqGnh/POsnZ9TkJan+s0tDryi7aFm579iJk
2v5i5GFCTq4MsqWgRwzGxjkFAJueW5rYDVW6oMKd2C3pPfJKnKYauGNK4FKn
mL8rW0ApF5vNglWkxkBYlA36V9VHBFVT270l9YdOgVAiL5wj4vYUMbe9NBBd
/5XpbpxwM5Zapu2gl0nYHBZ3jn9stmwtFAqZXrFQ3pfFeesYs463a4VudUz0
X5EhgvjkIT/sIxP1OdHV0or8H9ZVL2LlmQdpm/B9HbKMihDOeqmhv8AF/DhT
PJFJPcfCDasnus8tXmiTOsTQx9qVEiuVp8ui2ocYepm6dKp9jSUkuQsFwEtG
CTbulaEafAE4qTk3RM1GYx4K1LakigTN+PrNSxcyxuSCE1836qRoAhklTrEh
paPg+O4k+NmNaXkyICL8O/HNXVfSl7zLeQjCw9Qay2u+OkC9Aaotw3Epxgz8
VSD7cpc+LuhusfJpkggpQGNhjRDWmrJuKbx/DxjFbtGZpkz7b0i57L94Z3EQ
OjvT8pToHHsEpGlfC67xAS6jQzYUsHyV94OiQwTYMU00akh21Ha+ZUOkOMEk
fpclz0Ub2KmFapi0klrXqGL+ftDG4klMmvhg+Kk3NAUD+sN3D1TxJFb6Pt8a
2gQT8w3ALIGjYYsFNd7DORc2tDQe+fNENX0HWzlF6U6//ApulHxzglxg3b27
yCaO9q4y6T/EFjdiFYWXSchJA/FNmtI8xKLUFTtC9DR+Me/H2LHgQ6lk1/Bv
gnoeo2qSNAuScnwY7i2/9IfVgS0DHMiR85EdN6Hw7ZXIea3UbV9Ee7Gg9UC0
/RSuP1XbxlcNu7mmmulNkSpBHw4g+2sDaAJyj43MnDXGtLZrkQGeQtdpuWv4
X21k8rQAWrO72SJh5FvANBch42m71RPhZyEZrDZ7X53isCV+t83JZHbvZndO
Z8Mhx8MPr/n9QT6B3sEhkq5rPAW2AriaTSlNXAzhp2732csMWlRa4JWXbPYz
rkbLbV07K5BlD6g22lZNonXWoekX6L1t6OI5YN+8bTHUa+Vl3RTU3gl9UbUv
2Ydhh2UwIQgsO8FO6kUhEoBWUsRkcMqFAjeSBjK/+p1/YMJaYf9mVCeEBYU9
4kTsqvrBVw8kRZNSypO4R27qczXEYAz9kbjDIYYLg5NJAdIb56UDcs+gQFmT
/otMmwf5v3eF2w1TirTXMNJ/xFsP02eUzrQYWrE7W41X6/RKUk1JAe82jbsk
hwnWJ9gHMAjQ8z8Lct4jt3b/IR/gdpXDsZL8F0CGGcIRMf7pq7hsVkQIGyjN
QSgviQEQdBXLmhe6izbX+TwrDCG4zrc5sCt0inqF183C8HHpb2hvOgwvB51x
iBKAhEUMpywfpciKhlogl6IttW2DMntzg2hOe+K745qnIaEbtuzdsj5Q+vYF
0CPVfZ/EIey508l7bT8Os47tZortf6gbDpCj3l5+XiEWYndG57Z+WZHvQzkL
j7pD01IkPEDySqsSt+xj4XbupNVOiIvk9cpxkO3PyDx0diFF3598UsTtqKx/
U5HdUhr34m2Z5BpRFOH0L2/uGU60vod7r3+9li+ku1IX6+HUwAaDyZh5UXiz
wdydEDQcAllK8MePRdQ8OA3aWqTzh18wD6M9VB4N8R9OVvgsE6VaGeC+wpRY
wC/vs1ShmejdB85EYfNolaDcsO9oBjFsqIzfTBsO8z6BIn6NtMGgz5pDv66k
uXWyAp6b8aLU8/4s0/f5CwzTjnkneJq4gZabXbFsLivc6btBhD2T8M37b34p
82ywn1aKEOcHlbguOzGF7W//pBVCXnUkQmJohRvypZ+uCuNrZjl9Jq4Jfmcy
1fYICfNY5VxGETCRk6FEVwZTz3daa8OaYb+pUQDmMqI5P9fhoEgYTBM8Ucwo
hsaVf+UToCeHua1Wkn7BkPp9POuF/z+SVVEXzwMdeYmcwXg+Hr1o15oIl/u6
gad3BKJk7v4iU3ii9ky5FHpkJFtxJ71Li8f+oTc9etj2XfYGj3jAD6wGBEPK
aLcIOraKflqd5xprG8EMIpmEa7tlmmd7v2/AN1Y7jU1U8OR2ddzKF+/50oeM
gCdcSvMzkfcJffPMQD/MqJlE6jRkcJkfJxWVJzTEVo7wrqHi/NcJ8B8Hjmo4
BAqEnmRsCpOmqiRMT3tIEj8kqshZQxFs6qt8b0kTPEZRgL4gTUuIJLH3em2M
1vX6cXfMYa0F7l3o1epcCiIjKSn8lEH+E6Xvp9qhtd44CCdxNErf+FKQxOPK
ulWUnhPMJW7e3FNnog/OdobeLAXt3fBmIQnzoCPbQtwhiqajq6Q1TdnAHsQD
uyydDXtRmV7xp3nLg7jjfSJx8/rqEYpXJrICLtXS4+VmHXH3f1n8JCk4nceQ
7XKxae3fcdw6PGeYMMG2LaxZoeEKuZ7F5qiLY6qv8B1bI3s5c96sbRdhEtAi
0EwIb9mAAxx35nxZ39IrGDrL0xlFPIAEIYTTzEtkrH53KQM50ULjl9PcdRE5
GdcDKKoqBT1imQkWVkf1EfmcBHLWzzjz885nXLBbnUdDpi5odsGCaEjbWYh3
8fzSIcLwL+Xs0SyksjxEOmOiXkhleLFs7ZKTj6YtWCIJImEUqaRmybVV22mT
apcvbwz3Z/MmoD61QuD1qHxrNXnE8I3kLnv+r3sWRoGAQ3mLgclZB1A04KuK
P8DIeciF3MIYi6wK1CycumVXd+EYDw/EEyFXGul0yDWDZS8hLN8OVEOcCy1N
HtMTBSlJqSheUw7mIwe60cDGG3gLBdL7o7zvOsWW6VWm67NZZLU0Ykuqv9J5
vEowxIhxq8kYA2A1juRkdiD2uI+hdIFfGdh/nr9YBGX0YDJc/iH3RwCk8Deg
7Bc2iTzainC0mZTjU/Jvbqo3WR2JPm0JGFOVCDnHrCPQUTmpw4i6/PjEyJym
Wfz3AkPn53ZfqdsJbXeQ5gLLrHrYcK+T6cKELFbfI5Y2gBIVzYdZChuhrobg
p5ogtmaZGZvKSzwkYde5BFQLB/4QrrNJNOZsdB50K4oyzzMzuBAsjwPMNuKf
F4pafWXHUHT85JA1bf3w5giTu5DjQ3wGwbrR/NF/A2YGpDQgjoF5FqbJEqLs
y/iBi5iPSfBRW3rHLVuhqAtldgZH28sKNUxxz86kP5pfHAp5nprhd7IYavNW
gXYuntpSLU3vYfPDcXTuXI/B7AZa3g1PvmzMrSEjQFA+7B0GHkvg7BhUH3aT
7Rm5cL3xxZkAppJ/VOmuzNXtWx4B/H4WN/uEjgANqP07LQSRFjhEb5X1IfDD
5g8oFyQlnP1uiTkC+qHmalUHpZ0AFNtMQEK/1FM5M+pHo2px4hXh3ouVNlpu
ZqY3jdC90arVe76NFsNH+zNp4Kaspyzll9n8nQyHYrmL2b1K4mJnCpPmaKcF
R/Afh2A2jS9zrOfmfgbX0z/AiKsFVzparg6cCmgVyvgmEh9J+VkgyUw0hHBg
A9s0S8wlPuqYAlEd4laGQphnISVlcAtKoJoGroYyzr2TdxAMlI/73zJt4iPk
DBcv69U8/2yA4VEkSc7Ewamy45rQl7D8TwjQft6EtKX3SbfoTMS5Pp20J24I
5XgGWpqPnk/sZvgO6V9HIhgipBcWVAXVYHVHJlgigkfCQApjbjZg93yu3rjT
bH7FL91gS/biaY8J4hzVqvGM1nbEb2HTy4mZmKpqGjJaz1tnz6p8PaTbRcnb
hFVxy7PogylY5z68HzYUqRXku9lMd1to7ZPRLUPdye6cQI3i1k4QtaCvZjTq
LeVz99B9a3gHMKKZghhQ3fSXfycmEyJMwkIBAS3caNTJDDlMi+Oet0ymfIfk
DCB3LXQv0lnItMpMBttLfiIdHuMDrda/2FCpb/KPdZ0Q18Z/z3KpzsuDcmbq
64l5/C2SKGhTLsdbyG/g6XiA2duPTdoa+cX0/jjFnS+cIAyBLZCHpxaXzQyt
MLbAIJLFzbb8CM5Ce6xjgx9CjKB7t3kmsFkHEjFVKzd1MCTGu+aZmxB6+Wxw
+EyNU/xBU8hNqpoOo0F7bQNHanDNGiTvu3VsMPNSWmmU3cIWNd8kWwfd2GcT
eOla7dNaJqgBKHJ8isELeKcIzzx9Qfb0PldSGzVB9apnMZUGAv3cE6VdgMzH
wjl6IK1Iy4PX/hFmmy9szgN3A9Q95m/eolo8/CRCICy3Mlhia8GtYCwucXFr
jpxx2mD+uFBjpwZMp+cwAKVBTClzhCd1f1Y8RHAAYG2hCVy3X0fHEgof8sdc
NMtf8uaHIoJinPCzxtH6OVSH9hLez5yoSfJciPcVVmjDB1ZIWJZaSPzgcOjH
ToDvKA8/PEx7yIo7XPnuYSOi753E4yyaoQ//0HJ8M+rER1Ms3l+bxHCTtFwq
r720vBKYsg/LcVGzrWcSkSEAe3hesjoJyQTptK7mI3rZUoTFWDruhNcaDmFh
bGQ136bM9h5KBbXOS4WofbAWjmUwcZJJXMEWtRcGg431Dec7yptIfpgupu81
pI92FXytECQzsb4w13QBmfUuSHabsAEQNIArvPRJpCAG30diucLMreP6KaD2
Z9rWvscULrVvyuBMoSzVYWam2wawDYNtWjlSW47hae/enKl2mhx5rUWqsBLN
u+Uw+8LVqTaPxgFFQK9ip55exzwaO1gv/3yEKtLU7naMFvhVBFi//H9gZXZD
2Q1sXQEJgELsglg+MXiTsjuA9eXicvFqbnxu5tqGpko6ZeZJTJVXz3kZgXgP
CKhqILFM3qDlSyazUF0jTZIKDYW2Plm1WcKfa56JKb52aV9Gs9r8lodnAgzh
GLclxSLyWxg67SAOI8MScpGgvPThVM0q6EOe/voV1OexWvYz2nkcSxo39aQl
JBqm1qUEUSnwfg2X2uMFoTrBZnAdp2b3k0nTLXngBIzFoGQ+NxdJIH5oSm4/
ytoOWlwkm+cbqVu2BUFRRmqlhq3LHnkOvKmNWuiEcjqmFF+VMP6CC3MoSOzb
89VdfPlfgq1keA77TyJz3cUXQAAN0cb2buVLf30AbaGIk2S3v+PQi3QAq6YX
7Ag6h6CWmg+GoecQQe8JLCmCMrCQjscN2w8FD4cFtHb9eahkvLT5DSb2rbef
sx+yQjh6FVhMFyouwH95D+PI3Jjsm/f2A0yTQP3rOhLFx5xNELGjnQAAwMpl
lOoR8WlEWrSbNpIwpE181k579rXIGRhsXoeNcNDGbcYuklUVJFBalrgGVm3g
lAiGs+L2HRXhp8I8QRq2TpkPImtS5X/iY2beHnIQjM4m5NVgG59kZPvpdhML
GUCH+m+HQws9WzcAshp2kuNGj4Il6eE+yQiVtPiAs6JmNDlRJ0KoeEPzaGl0
/furxTjWk+VtHosTvda2h4rDqF9qcYYmVRpT/pUPImd37zgkrgzCuVpkBiXN
ammAGgpD5rQjuYOMBHt5bcNv4w8+yfAbX8PqDs2uCfQyGATyB+BDUCEIsmON
ZxHjUBBJ6wtQpRu9bzuLg8x8FO1Z+MsAmdd+mVl5PUWi8Uws1lE8A0pyUY+t
xXJVlO1rXbLvkS1psbC8Mjg2NuE43gYI93N/ztJDXJFXCJlydxF1HruF29Pl
wOUILLyOjBj7gjHRBic2N0Qd3vw94Gf/HOqr5oOBYARzfpGfkFcY0C1XwO/C
7d9ACGVwHu1qV/V5DHwCjTPwz4NDsc5nXMj8JkIJsc8q146T5PYbcWAn9yBr
CDL7ZjsaGtAZOdc9UXpkASwIFZScocjXrNiVSqh77aZznO1/DSDdH8h9M/JL
gX7KgF2tbSSC765a1PWoGU+2l79kyoUKG/TMCttw+jaWcB+zefGIDxJTdvr4
jeE+hSELbWrv8kN54hDrMz1AuAcxSv612yX3QhNP653GxT3FbP9KA1zvUS14
iwVgvAR2XmKAZmInaVNFSaHDcMKp/O7dWmzAwRkUS6XCjO5HKEmqYIeeQJZ8
KO0why5yRig/wyO1CAj7yaUGmquqV0ZikoZryDZ7/sC5oIebib8Kld7tIvfa
hwd1Zo/yX8XzeLaGX87xPtfHYrH5EBC+rm/63AG8UY5xGg+2z0Ez2Lre8QRb
jEXfhY2+nw/T+auIbvPEizgoeibPwpTnWSDZnjFnLiUgzX4H+8gjP8zaAvLO
zpW5K5r7LhqpUbopEJu1hikuso57cRGfpvCjxCqsM/noGYxgnAF57TM8cZ6y
PXuKPz3EPinnPA8AxUuCdzr9ocbIhJwI7Yc/pasUsFWhfxvuBnmW8kjnwMEK
XYxnNJPv1HYHb4SQJrzQBv5R9lZI1xJldcYi8S8UysPKPACLXWdUdtSfh33w
90TUam51pDEQU7IdUNAd2j4NiFV87XYuNqjvq6+5gDxBFzISFuxF1esb6LGw
auWlSPp9+MXm/UPdmXSOqYAMJYx+RQrMDAtKmxdqaV8oV7rag42QPVFiXV3l
bp/RWgG05/Hgt+8JiCKT/2Q1u8dG5XKkjfayAdSVnAoiwf0I94v1IQn76WuN
otMhN08F75Hx1Ce7zWsQejPOggYRCy4Nrma2DHODWOXMqrCzL9pBCcJjnAwt
5WWtCaiFajKDhpBEjHHn7dIZKWzDY97FyuYTtjwyyD+k6SIRfxUVimebD+MQ
3ixerW3NHPr3v/Xww9Sg6F19PZIqXAKxdpqy6UPtsP/m1fPjwfE1S7eqiWRd
Y8VaLoAjW8HJszRoLDDIWafmeaIJdCK0LY5i8KDepG4x+ahMpV1wzf5EAUX+
cNgOn7aIg9fxSECZWTFReiAIjogEhk0EWGcmGZz8H5exlv+FggD73sp85HmW
imxw1S9tVwdJRRWv6bgYQFmla/hmoQVCrPJXgY8s0OFFIwXVS9APgsjdwU7L
/LcfcAaBNpUXLXxBmTa1MuDx4sp7DqR98tXae+MMlumPS8J5M8u0QH0rmVW9
0/KJuG4w24ZwJXpEh99IrYecUCttM0RGBEcu36jJ8aBeNuFMnmk5KniNBi0Q
r17biMMH1bLbIQ8zABgeG83U6GjWH1UYdbmkUTRmKtdWTgwCu1WbFmY6W/t9
luLWnKQbY/ubotAl95pNsTULay1aaHdto3ZQJ/GUgPgFgJtz8ayJg5f+Iegt
tv7IcCsMjPinYcCVCOBStCUD7wsAyBDdecqOOIVbkG5/55d84LnmSxmc3248
1w9xNXEQNmaWiC2KfTjdOKY53X99s+p/MlH/krPhUwFsQ+C7buYM8uP/cP0H
7xoNo2Iae7PMJ9lAo1hjslt5WznLrNWLiXB0FM1mjb+e8AWoTeSq5DsKhldI
zkLMP7hC+4wdSuPdz8M+VV4G5F+lPijs8FYfzufzrHutxmjb5P1DDqp8v39V
nfPwk5uxLIf+Gpiitp2/AWWo5Ov+kCA5rsATTa/Cu3m3JLMx7Jg5Hsk1p7+C
OAzVua1YmXaqGqSAA1UboiM7I8Jr0WxMVbNx2XQupIohYJuuoVYCJAcOj20S
Tb2HOwomkO4WZDpvhoYFvur248WKCvV2+jnaErYUfNJQWRHs2GM8UlZGdpyz
atQ5WfYAAYnAWLwl0YtnuYK8pwAboWyaifQDfXp2c/Ahw0BXwAk2ZT+2i3DF
rCFU4PgpNMeIZJqhcv17h1rgI5gQAFQbTC1jhPy1ChVPRfJmJ5/IEvsQapz4
NxZ9FY4IOEjAupgosOEvpeTix8s4iVxbsKDxmbDfGUWHg81ztysvChKEqx1T
+iJXbpyLwqQ2KieZFUbY6CWEAPxOE6/749cr3CVUbtizfJMU3/SKlu6b442q
38/YTOggcRtTKu43/SRpaUeUln7f/tvpK5LHoG5XR1MIlwYOiMWpg0guySce
Iovm691Vib6u4hU9vZ0rvsamUpGKguL96cUylUyOOcku1yzvno03zNUrpDkr
H1Vz0JMkTzFMJYytpS3G8eUa/gFSqLIl0+/X7FRJtpcG+UbwVNb+WnJGQjiV
W5cSqcDV4x7Ftu7DEvi4f8EXTy+Axlf/l0OGVMTNCSQ0dIv8BFdTs1haDnwD
jkn9A3djLS3XjjoOPxbMETNSWcYtKAvWK6vaUOG1NCqlDB3XDF8wVtT76EeH
uvLvQ9cBt+W6YR42P+w2swOWEkYCDlx82TP+eqOSoQuftMhqh0+o/NwKEAz2
bcdIKLKanB2+rj6HyEwGRW6z/ivMdlz3aVpGTKZIZjq4XhsVpZLeWaypuSx3
T1asxJsIGWHvt/8OjLLCRRlppAkOBa/5v6E5Hqk+QwJqW/EvwVx8aTiUfx+A
h3FIdYJdDZDwTFL2qdciGgu8I5IGTjH/3BMVG4oz9f+GWD2L/rPCtJ1MRg2I
JaMYN6IOqzT3gFeFVxqzzPMn9/di7dq9vPBJRnMSRdNLYMBRBZUDV5vbNIRw
pE502YNc1jk/lRDM8H+83iSLpEqUJewU2Qe8pjvDBROtkBQO3ttXKVnjkJXY
T9pulueu47OEVD0PskhY/Lvezb4hR2DGy1Fj/zrhYfo3aL3kWv7jUVf1gOku
I6lBzL6uMX7rD7k0Yv0fPhPbL6byPn6Q9Vu5OutWnwr4dxbuXW78p3nnGLcv
o/E+I1yMssSyfUxY7fnyDP8/f/BBxnj0RE8fTqoF9sqLs/uzv4WD6GGxe5kh
W7ZKeKomb3AZv39Xw9YjVui2eEuq0hYt4vqyBUBIyD5SJYxRJqOUf/1k4aOP
5Tiprf59h/QQJlodhjIJwNd8Un9gqvIqtHkQKfD4/BHzOumOjoQ1LnAktAMM
hwTSOmKbIpa7LCIeh1oq/BWI7nMhKTDG/6m33QwZAmQqCnhybka9oppYLncs
96Y/GNpO2ayVgOQKOSqlpr5KDiPa2KOCrX7POkLCu3OrvRorntkkHVfrDK75
xTBQg/H7alknHw/zVre+hq3B8lzcKt3ybLZubcCKJfwrAx2GuO+ou1gRPXOJ
4mfFImZnF+M/cvInlr5lc4ItzLAZqPrPaTd2yx9zqjamHxgv3m9wGc27/6f1
b8DivXqhzWMV59y7zl4bn3SZZLcwV9NGeQ8nOUdoYYypkdffJkZDBlCNVjej
IShbIxyfmSJVlJ1syp4ppkjFWaV0XJ0yFD4nbOLqUPY2yn3UKE70DMnE1qb1
WWgTb0rIp+h+EEeOibjO7Mh3snw/V12QBvnZdwAejDYLfssVFtnlABmklHjl
XC0HffAZTZczlDE+O4F/oY5sHmg+6aCvUUmXxHylirKtNMlg0m6ql4MpuQQb
qPvjiDq3Aa3tXSKuG5BYXFYHLRvvWznDg8cnfyUWSH1/8xgPViPoRWd2mA4R
IRY/UoS3U9m58tTcpZMuML/vyUPz2SM1bc5TOHdhK48HutvrEY2ILuEj1XM/
gl0aOCSAboDanZzaddKYMxhCR4ltlOzpZ8WsBeupwXo9P0W4y7vow37d8dnM
LZuLJictUSAhGHfBmhtteyif9r8z7bkWH3DYCc31f1Ra9UU4YDuZ4GhgIL5l
kEo3Iku9Fu+3yDzlMPJGbGyGaFyajKXDVJJSuOfcb3Z/OY2hNZ9grCdbjqBd
4QEoG/um8zCvUqfSwbLoPJKUvZp1+tGHqyEFrf/J2/MwEQcaAwW5KKWGd4Sc
Y9SdQFsANLFnWwyilirhWdL4BOAE0nLSlHwkHctaPEQUfbzmQowF2/IAk17C
1c9YjyCIL7mHcihlxd+nrh4XWnyUyO/S/QIX4U2j1k41q9v2749iQbbfcUky
KqTBknY9bFwv5OryO3PqK3ZYa85031dHNhVTqmfJH/PmqwPa9FTZbRIgOfQq
wYMs/8Z+TnOczmmxoANm9eK9KvdcmGpP7x0WMlONPdoyxeci00lwLiM7pzp+
FZ9Lw3Wh6k7SZD8TJbvq3qwoW79K4Xo1aYtFt3T6RWcGqFYbYi+jeFNeCxPc
nKi2Z0aPhCnOZvAlfXPgwl9/4mVDnO8/N4l/F/MfXu9TJT/p9Pmb/KveZx6S
WepirZKk2paOBJ4ZX9fDuEjBOO97To1v9Y412nyZWfMEtz+9mfjnhrZupFYE
6pHXKewcziR5/7/gzrIJtkrre5dd9b9zzb57zvOo/5+4WWkHjlqD3e+ZJVdb
PvS6zHV2IHSmP2ccS5cQkCKfBTSbHrOOhcudaV+RuE9JrUsqf6aa2LnPcRE9
TAJ//mqm/ACOjzMji9VJ761I0D1R/7WXOAhZMd5LCzAIB5EFDo2AVm91QWZp
REoYBm7u6FYSwfQIPw6Zka5oRgk6qxydwF+y6P7Q/azZQXJA8ofvPJQV43N/
PWC2ekpg51vOpJygXPrIfzW0Wck9g7NV6epOQMb/DsmNmVajuSnPWTiy6nJ1
RrzLRdpLwpF337JRDF3qSSrU2ArHbN7mA1tkNDg+VXBkGVn++NBgWwfsFJI4
R823C8jGurlu2IFdvDZMN+8cD616YuQaopSHB2hKf5UT3QaTZzeZ+ONi8osf
HogBdgfoaFHsPUaY7R98/fRYK2EZLNq3NifRg/sBgq/NS2358FLOA6l7FL+U
Rhh8I7paO4G919dQxDez4H32g9HNzVGg0mE7GSuIrvfqg5Fa+oyHR1Wq/dZh
NKaFCJVkOySnmdUwk1eEx73BsHHvzoz+xXWVIb6i4pamFU6nRM9VHZHYLwhH
vt8b36hs1I1nWnkS1NFbHF2f9MBRUBlWIfTSQBjh6cYIepPnufiHhM8WyI4h
1q7cK/JKFHAxY63LffuQMIbsG5L358yHyogQtGOlO39A5eTYyrQMPI7rwy40
ArqKVg3i93OWSKFwh33393xGTHSP/9VnJV7eealyMD6a397H1uhrMlyjfoH4
gCo6ISemV5dx4EaKrm+hz4YT1KI80N2sEwZNpGIKS4Eezf1lmL+JAB+HtgQT
sCp4Jq0xmRh30iqIFulW2xzi1ilo0YaevTCk1JU1xxfQhMbavC9WHbTKXknE
HWqhbEnsiLQjRP8JIAYNyL5sX8OfDhYdWhICSLqSSs0Yy/YHu+2XlZqAQ9dT
3AQ4mb6dqsXtuo6LG2LeWY8aXQWesGQoZ/if8yUKq7CWkoQf0nIP4c7p1a5Q
oTAfeav6EYbbxaOKA49N7SIVx1nYjZ0pTDSO9ah8E4AIoB7nUjPe2ucJcgmG
gQpjQetne29UGCE1jkuxAqKl4kNnCOzXQTGT4amgbgDo7N8lgz3fLo6n1e9i
7hxNpEmE3cNG8oh1q9pGlhEL11lFTnSUW5748r3VfpI4uIPjvJsntYSM5Sy8
QW2YlWeAt4UvjPWV38Px5GOrw5WZXeNQveTXVJDKYa62ph6X6cY3AO8tlPp+
H0KU+JgEPUVfnU3q98p4JsXaTxlQwjL/eceW+H75JOyGCQu9Zqre9xwQ0pHD
4F7fiF1xv2MnmzuqtnTR2MfD3zymEpX6fvSHBcsd851w5PKMUAXWVwPoc5rG
JbtkR4OemUxDQ6E0R3mrmyu3sZpicAom+hoM0f4kLWF68jDLddID3NEwAmGS
UTE01lWqEDQEHySgjPYf3NiIEo3BC++++MHcgvE2p1V38Th6sX3dyekaGIS0
2e/tdY271gejADfkBl0OHuWMvVHueuSM7cBz1IYIeboJk4jw/UsqC1Kvsa43
tm4Wj5METUpGOAXqsVn6n2cXhuwU58E5r5IlYfsYdvpRsCFsJUEwOdm0r6Rq
jDxqD8hmGvg4lmBf/aU6/0QjHt5e8AJxbSB2sOENVYAclweoJe4lrp2Bcc0/
+UM1dt/Y+7wt0B40T8/WCp8hL0nXnn/7+RnrfbM8rWxIXoKdigVklAsu0KHI
E7COSgX5vnDgdPm0nx/bUAnUl2rbtAT6nVTHr3o+Kmr+ni8XWR8xnnRApyje
LJtZ5OnMBXvV2gSVjxJUNQBKJLpiBQlPMy2ZmZWK3Zyh6ldzMAvFkFgU5v2k
LUjL0qH692hBtetX+ZonqTX5xjInbQVeRMT69hICp78pwKEYZplGIoZ+YZPf
r5eqdbGJt+5sGG/TlImrhUAPdl1odn2FhmDsgAG9pqblbQtImY+JMwcRkp2g
VBK/pnb00p37TF62jAbouYxRiM7X0jWOghrBPQIZN8Ktx6XZ70h6rvi7Umqd
JKmMMpJvXERST2J1wcI/jWUnG6yHYC6gugR7FfCq7/tykRxzdEQcfmbW7WeV
HoAYNeVP6c0jHfk/yhEdm0uytxEDqwsno6F9Jh3raO/yO+CUvNf/MfIW2ID1
6obokSkMBK4LL1WNT92gKHNLMbYfuq4L3MXtIqSh9L1MxA1N159P9t2H7Vsm
tjfKFUN6jRMPbpDCtnSGVrxz6nfpDv5722kbDT5hjBmDqlzYUoWCtd9bKpJb
YSUdYjSaOnlnnK+gKlMG4fN7BrLgVJxkz3F01ztOxEiBSOksne/G+W0/OXzM
eqXmKf1vS4oATUH+Hov13xJt0416pmegUvmPqitf+IzXF2YLbK2nIz2cQExq
/2ruq7vf25CdxPdgzHFyLOFIvVTzo/jZy5iEhHw4BDyGLUpfVAEci6vnTOmL
HGvUbw2j1RDxU0x0BfHSDumGKNVEOXZ9WkGTzme7uxLTMT3RJhMMPoSwzgGL
UtpIZZAo8buvC6VNgpaoRAhTnWaqJU1J9wo0ihdIyrZBjW+4XUvc7lnto+G2
JefM+DFMHNFvWMuhOGGf42iHZGdkFi7dSjboUteLwOsn98EEz1qE6MlV054T
x2cCmErZPprSoxs3Q95yNoInKi9ggzsOxvas7/U6xOOfuot6rJHS3/lyD8w7
0BxvwjJu+Ik3gxWzOgDOBc2/L87BwQEyZuPRepWIJcNWnITpVN9yfHCr49pj
v3lFX3MkRbJEks24k+ghYRWnMq3Bep+RmxuYbPTSouq88bHNDmIvw7h7Fdjv
vNLiv1jsIOLoOvkzJh6pI10iQOUGexXROM67N2q0j1i/xzHGr49Y3AfgABwt
oPSgdCFzf9R7yoX202/Dj68VppQIXuSHb0IN/dAgO4PrZbksgZ7sWKdURpzO
5888XBNlTOSE91ZaAUOlghU8HcUHlTi6UHdb8IA2p9tnQ2MBlq5uybMeu86z
LCz3OdWOtneiKfN+rzp/Kd11bL/lQVqDIiWhGNoHfoPSaKXc9X4wpNouznQM
KI3L18Y/TgbT238+YnMZVNajpeINyvQYb7jITyDrTTZ+8ha/2jHPpomHeIJR
rmMhIlP4zrPt6utHpY8OEdYv2jaCV4MTC3wQsa03P+wi/6gKiOsgMixKBqP7
Cce1BWAFwSRr3PR8vQDLFwytoPCYuiVslF/Mgvkt7lMH8DA7KLtwrMqPjOP8
IBaVWA0zIMdmOa9vtKWa2xDjbezlnRHlD8qq9dxaaHjcOago0hwkQLn7cxkh
6FS9J4aPx4FiCTR98hCf5CccuLV6vNwYkejhzgIxPRsiuHjzZYbnmNao/P2c
q+sM6hLVHgM5CCCJ+iSW+gp0vtUq5PetXOyVwhUP1gC/s+AKwPrG5BCE4ody
jDP9zmF/wJ71Ui45upmgO8+JfVdvZw4ndoMYBIyuRliKy3EH1axHly1alwFH
BFbF3A9Kk6ePIdHMqdWrzeOBuYtDZEE2LaQnAkLPkYMvV8FsMxlZg2IBulzo
WwMzo0JWsBpu/zOKzfzYEBZKU1+Lru1u7EdxW+TDfqOButy/BmDiNvaPkfhd
tTq0V+NWP+uLMwD0s1QxAZtefPY2iRyn7TA0L6iKWgFnEdvlOhuImxqFrDRy
2tQxKxOSzoJRadb6efrL04uoqCj8MnBetfzUbv9DuLLq9Qq89MY/XohV8EMd
+eEpzGUTHjkVdhzGOWbA+hzxM/tSrbzDxDp7UXeejifDZUij6FGz+PsZLqI4
4Y0aaMAbIlonZah67EYD9wTJxX1Qu9hZ4A2BfKursTGOsXnE2P03LraBvsfU
MUXPo1EBx5xgoZ91Gu5SKNnUNaBgObXqxpkiWROHZV0wXQyjEysiihJ3Qq+w
2PYysu0WI4nBAw3w5XpTq3VIj49BGpsik1OiSWp+4LWI3HCnSaGb7T8tiOxt
ZIdtMDsRVTaUPn3ZHhSldgZKrsQgSqgo+/49fpwHhRspmYt4oCk6wnUiTiiQ
aIacDd+/i4LE4z3G08ucK0QDzvvQH8KKqIPbhPZLre1ZtydaxBZSiojQpOKy
+5QAUEN1C4IQPaI+ZYdHt6XHjWZZNYJqV031FMrcruy8n0ynqL5qa3w5SzZI
0hbnvHnn4zGtOd5hqqWmYR9K9X0OaxoYAgwZM/nzmdS3jlEQ02IUw1F1O+8n
cbSAVn4zPAM7zx1V0RSiEdxvrOyeC9MhyF024r2zZUFr5GDXk6wiJuDu8DZC
5enm4D1tooViR4esRQl8Jjc6v9mA1u/lxOGj83/T7yWWgRTRq99DLKhEUold
aSv/ALn7yeSaliA72ft4AECMsI99DgqMW0WbHr70S6tRyvP4qBey93bNIcd5
X3HdbjCXPPGk9KqyzCAY3fdhyfLOzDr6slT/lBINCKyZ687UMYCZH4q4nVIX
dsuozz01y4qZpFwoGpdzma6ngNHfJdxE3mZrOONfmvIEIx+zkWVKcjTQT0Yr
zGVpwgwqFV5zr8WeCYwBF6AAy8rwSsRfHVydHSi2THOPlb/CMyvwkZm77toa
UtH0wH9+xlitnejUWwPs4MCvuV0GSoLC2cd7NVc5cIix5aLCyQFk3JB2gTEX
PI17SIiLJ+pvC253OOJt1k5mhfw6NJIrIYCl9CF75oVjeE+j8oKgxvSGZjS2
QsHAe9cJoSRfHOzwA2spg2UxVjU7qaNBd5u51P0PcvrS7ILkSR5a5rRHTIyw
r9Lzc71N/BPKyNSZhvBSQkAuVqNQcQ7XJnJssied0+lxg1OePiH5ZvylMg1D
BN/M7b8sSer8N178PlKZAlzgzeEBEioMzyE4GTGbNygx9ef9oeQrKB1zBIKA
ipYB8fXbSof+Qn9/s08BbTt7+hLmhqJtuhWS2DejqU5eZUC+78Zp5yfMEQVi
93CnfbSfJz6Yq/L2e4ev0NWu5mAo02RBAkPLR+kuR0Wl3ZTdRyi2fkJDub5F
2vRkb6YoaqvYn+Nc4aW5324ege+QFoFsvziTtI/qelDWOli1dZynNA4gxAWJ
QdSKLv5BOtntohKt7dX5yVjissR+JJ9gbZ/Y181lzGRi/CCsWFOQiDV1xycz
gMIkWHLk7uOdVu7HTFDK/4Lup507VJJdfewc9AttNBldmNFwr1Kh8Aopu6bY
z2ZIVjxPjZm6K2wN8/8kGpuwgq/ikEr09KcVIa0af5ayQQ7DgRW8yLZATPYe
DZXhnBB08AizFbdIevgpT40qR05pYCIJf1AdyOWtetdumJC4uUaOeLiAe784
TgaH8DH+4YxX1mW1JDWsHAUEH+1oY5hoKR1bo+anDSvUQYMhFBU58cXe801a
PsCFtZ2oPNMLTAsnf7XI4nbPHpD7H64PEDErE9AOsBkPSU+ODVdJh7PEUyH0
fNbUcWnyHpdcxTzcVMCLF3jmLysOULIRyihZtg0HFSAltT06hZKgGnaInctQ
mHCXuQ2G6akzyN9tejNdGLvA49vHEIsw4ivacIPKYVeMOujphRAvLlKl7vR1
93yTMiZDSS5j74/EYTS8/o54eoH3WVgwUM1s9qYujjfGNc9Z39dZZx72O+9G
BaSFDWOxXGntY9XD4/A3Y39mFwjyLhwX9xbfQ/pudy6qkoOKOJodWfy9G4zT
15rY/4FdkHYPUMpFTxl+XRhyQKwTQtDsY+xRSlPiVvviI89xBWc+z9rVxfY9
2aQtV4E2KQV8SKKiy+VxmmX5wrBaGWqlK3R/djimGVhKi+jodf15fpad639D
xl2RG6wAGcWBl3tag3ykUsErFPfSCKmtdTsueCQD43EH/7+5tVpafUz7Ip3c
lMkh672eYF5By9qLPIUCh3uPqJoYRFi6+9tW8JZQFW8UfVnmrI8GjUNYOP0O
BFEFaoC72v/XZwb/xnbgmlYBT+QyO8NJneh2IhQEeURI6NGvODLb8YYzY1z2
x6/zJNjdvsOUdBYKbBQvkvQ9wZNvCZkkIh8KlFeAbv2UBzcU6UaiU8zQOya+
9UEiaccub7viiA0ykzph1FGBGJJihRCTjfIvaKMRjRfhNt3DxGpJtDIpiNeK
AmDqLLcjeyG30JTjfVkesX9izr1Pya0bqs1BmETZ1tXeyBs4ABI9jd8n9Shs
GYyyKgO6/vafcCHjmAoZcr2n0jwtwLGU5ZOUZASbJbUhapHFUd/IpLapxWa4
gFtrCSOpL1caaDKYZeQF559H7PHN3aObbI/O1A5w8FPgxMeEdA0dUfN3spl8
FSCQGOuZ2Talp5JHZyO2Da9k05Lc/EkqFt0Lqt+8CEmOJVKL+5PGJp0ldv6Q
70MRcDn6++zmgsR7+ZrnXLUejgIqKfifz6aFTaWxKLYAb/NlNCNfrkPKqzxa
CXcwSyvUFIVre3pM2GteAdVtR9y9klxAV5z5BeijtaMoESiY2EECfCv8fr8M
H/V4waXi9RMA7MdItsYgrvyGfSc+16tGr3gemIkG0eal3scOmgFPTzZN334j
XW+TjkFojNEH4FQ18KUNU4VborGQ3ExbYcgVT4ULdUrr6ZjoHeov7fhx3FIz
R+V02DA/62i54rhyXaJ2erQv4XRWDOjaqJmBOVcxtJa11yyuukrryq9UFHyp
hYFzpL7EhdENgtTBERdVbBzDq3xYiKxM1fDkxgog6+iibXHZPUykhcUCP7XC
lodEi19g52tSP0c4rdUGeiEVyPyQT9NVcBchxTvJ6oHNJDszslas8oNywnYS
92mK5SFMwh6DOXMfFumTWRBGsuDI8NTP99hzuCcXvQilkoaQU6kg5/OFUyWf
JBLjxzhk/c69sVEuNc6Jq0YMqyCMoJ83bL4eaoIdqamSTYgUE+Iea7aJWAJP
WRSGE8CDSZ8MYAH89ZGO5iotcRHkwnEfjtVZu0WRyqdcdnb/bn4n51JfS2T2
/PVD7o0kWon0vygzVw67AdcOSVZOx7/CUe3yKWjuMYWIh+3SF8unVUr0J1NK
qlHz7lLn/VWt/g5OuQMkuFnk9JRmYNZJn6Iu8Y3KxMWrKNLK35Qkf6VLjHMJ
WYPRma8tYrU6Sl1PlXAHklncvWNLgb99dVk3CRMIh5hJT+GPcRrcvGl+FzoL
0N34gDWhMyTxz9dJHyZKSxWvQei4vEFcHPDsqkjO0wNSg8agcJWVqeoZ1UDE
PLn1faG2oTAhRk12YgUgPczJVoTp1JLZo8hv6EkirIDfrFH4C+0HoolHtnnB
MtmCNJHXr631yR5WI3xHlfBw9JALzkcpX880PvydsuYSDAr3fMKPKuubuYtb
Ya2PjYwwOBF6ar1+e9AxXBlNKLB1JxGpRRrghq1g4LfXmcYEm/wNApD57Npy
gg/3s1cVNKMbwS+f+YoaaJ3YnaxAgiExJxpwcBzI8Wt42+m9JTV9tv8o6N6M
GMislgtwdErE458kyIJqLV352ko8wLcwBnh2ZTxDazktc3SbJwiCDYLtxkBb
PlzCf2TsqvSZbSVd0dW1PrVCToBvBqSkHHqVKc9WQ2GJV6kFlBHiiCHriuz4
E056xmw6FM1adOK7kDTD2mRtSsg2RLFmGuatF/L/JXJfksetIpVlvf810SuR
+T5CW2BmwqdpNKYg4/AtthIX8Aq3FqxCqgLlISfAdwdMtqwQdO0gHbTR7NLe
wHQ7IpvoOKTZ0XbRtdGsi+ydYy10CUK6l1hxo1AtbB+MXqKcYmnLF/MScuzX
if3mm4a1/ZAhz1f0z2+eUqtI4trviqUPxAFeiNmUTCzdDQjlvpTihWLmqXGS
/uiDa8q2+8h8m7XehhabqLR+7WqtNF1B4oiq7IIINVlYoFbtJjuau6Osx2fX
oeRccy5zKCIfG6VFzqwdRBI8M3fzXM+8VJ5+g8Kdnv1xoYesvPoGbhFA5QWA
J8XYtzv8hWjkJziFckLwThlRS14FNTZ+5ufF+DzTvCQhzxDq+8HcBWRreWm2
1yo5CXCdU+8icmc7mBxuU4nx3d7j8T0448B1s9ARjonwOOXRxmXQ2W3uoUgi
2PzZXDPnVuX2oBiWaZZDDpJOunZI8JH8NoMH43tSduv23piR2FXxbRidznqu
fbXiYtOjaRML0E3kLL9UZdW/ovsN3WDo5wKzbnTqN4zs6cblhZ/Zui8Ay426
NqkeaPc2FgkLY/6MBeLeJSMkP/iYKfwFAYB6XO5K8bhfS6QtIMApwDWANvxp
I/3OitggHS2y+WcyqoYHMk+LZOvp1iy+dDrcs83tK3RfLnyranD8i7hws/5k
O8grkQRkngz6pQ79ZdhgGBLc2fy/8sEcuaZpG4ocVSHt6eI6H24LLjf5BSo1
7vRRgu2cYHQFzAT/DX36Vf+LV5I2reSOYgGYmVGtUJgLRCd8A92cITZaMpGN
wyBPFIMxa0HUhjUOtQ8Q3T/OpOGdcNcvU2/I2sAfAWtfrWGtZGFdWtGZJa1w
/2fzmKmzAHZThWlfXBi/tLJ1rdeD+/34fp2jMvJPYmyEK7P4SnZYAqDJPYEu
XFLo40Lf8BplJoRos7qZYxK7QvAOHq0tz/HkRQ26wMnjvqu0kXGlxF3qRkfS
XI5tFiCqoCGogf2+h2yG3Qr2oWxeDI/ZRDEE8OwYnq2+9JllKfN4feqYJrGo
4upnATb//ObybTpafXl/W2o/lIRxT0kqe2/+xmKWoHLRJD4zK0BAprz+1VyZ
cH42PKD4O4/6qTemLwxmCc6l7uEo119Eo7wSxV0h36yvFTzT9lzNrTtgxYY2
N6g1XmDByP55AZdn27Pi70FC5eFZFacL9wecEZ+hCL+tZwgLRT+D1/uEtIc/
RiBcR8QfV7lWJ1M1IVlmEFlfhLrhfRf/dL3Eg22LVKUX1gHRiMe4RP4tKhq3
IXBQdfONKq/6Aeakf0KWO47g8EejkhmUAivA5QMffsk/08l8UnEwQC9O+Mys
hNwoVCoyxixa81NexShAVRggIe+BzDAFa3oz1/2xh3GZRYgAEVqbOKWzeb2A
Q4cCIpxtBsBwL5W/x7Yh+0aNjkNtnXem/ff0f+q2tYxjdGeKgwasU6vC9fZT
J1iMPjKOeQGmMFI3KzcinCw60ELiKtwi1K7t6zUTeoFAa5PJNIxNzSpejFOd
H6/xgZUn1WBXT6iBDwvT/RnKrwNE/N4hh3X6bPIPO0oWRIUvgSnmcI7/3dIQ
xibbvN2n3V10yGseh2hIdjbnYoKl3vaqd7wST0/DJiP1UHyPnvzbc5tYb3Y1
h/akiulqOSYfNGYgFsNfJHpKJ4p8EJIuRQzx083qPX4xccC1YyWbSA1YPHSD
QKgV+AqItYhnHhPkwILFSTPUvJ8bnN/1JEm8a2oDCcIXoSjS9bU9zIYNhJrl
za0wQFm/2BjTi1LUQKxzoqEaa5cjKHe3XEyvM+EMpApdAbsy7xC/mr+/cBUD
cRELLAYcn41hiIQDFMWGV9kWDvidB2OIIXgyLYCvCUoWaUDTSEzanp7d4qKl
g2LkUyjWRhaYLYGNNFbFiblWqekHcB2+0zIRAO6X8kHQGVRiCypP128B4mYg
Fg0sEbwHQbJwIltETlzI+BMfs3uUmcboyX0rRuWsxeIXVMJFzr0HX8CEms4Z
QnQtBvhyeFDpkoHfk39NJS9LNsQF6UqFmXkMlAUUZPnHBvVxqPNl6w+8gEdE
IuQXrVGhlRB/gOFnTrbC4THYCAR+bz0WMd92LLQlgFOda2kaJXclM6afROFM
0PxmtODQ8ctF910QcragkW8N9mN1/Kj293VLFTc0qgGHoRGx7oWF9TOcBMEe
PuC31GpGFrGq+SGy3B6JcWFAUR2bPIFQVQvU/wiMZWFZIvRwYmt88Dpyd89x
PfDrwXtuWpvElj0PPr96Bbd0xjVZy2aEXAnMYsjRqtQzJzpUiKyMmYSb0hCC
mmnyjW8OrBURmCZ02dsn2CDrTuRTqjntuY1/BCdF/05lQN5NiDBlWSnYCw/V
LJ6z6cOeuyOXXpVwb07GF2sN9V/3mt5OK5Wox3oqjvCWEGJslqL83FRO5XLB
7Dj74MCHQsQQ0bMa7SU7hfOotasqSPIxiUovad6AvpUsAzWRsfyjjvehpy9g
QMFVI8RQi6SzWTM2x1GyysEHQttjjNA00ZWlwnO7VsyAcDHMsjiWJRsyTYo1
cMlx3CQRI2m/dqE3HfHP6Kk+GqZvXuTYmeSnpBdRsZc3R5IyLVgKbGv1jFm5
ve8Ifuv3QDuAYcL2mKSK1GgRh4eG3VKAA8u+/1UHayRA5V29Puz4QF27lvoW
2e2qPPt5lKMwtcY/IzvDqg/73wKrcg5toEf9x3zWsza1vkizEylLJu5oQ/ww
wPaVHIjJlYdj2BJ76dBqdP/xishWQRU8l+WQi4dq8uMDXSWHqBKHdlGYtWtF
qZ97AaWI3W+o92CcBcnK93OeVbwhV5OIOVaeTQw/UfuwKs8J+UHpyzAQQlvK
irzsb8lvRFmDzhQkEjMfEb4O861vcecA0Dov/0kry+ZQbdq2NqKSrVsdXHhf
GA/5JRBhhk49LnDjT82Aey9tqaCm8PG0F02WIY9Ev+LdI5yKC/h746gYb8V5
tK7ybatXc5x7ygFDP0ujhTtvDY0Z7z58kjLhoeh0BL/32JQCRHQYpCvpEiT7
0knQ1Juuwa2xfoJ/MVQGhWFXfJH31tfeIip3LwTvHNNYIlpGNKwQt4ClihJu
62gaSNf8PfvOEOsvWiZqdDWRgOEpu8UoJPwIh2Uc8EhOW9ZLPRTF//mjgZFi
9mHQXl8ONQ1uuTenoz7tivsz/AKhkyFaySOHv1NvXtqpXdXJtHcSrVVez5qs
07RXnT87pJ8uVrcuhtXjeRi2c8uFJYFJi5OjwP+VMnfj11RWKyjWMMCmNnI8
0X3tpXGGQ2mF3bAjz2k50BG87AKdaUpf/ceHGuavWYhScQeWWT2EjElxk9qc
lDSnvchyTbPC4r1ND/fsUBnwMdQZftkmD7tgGjmItXEE77uxKNM1GPMFiv/B
ic6X5drQIOrF24iO4Gs37LKlekEre3gjdSH4JCNiIi3qeyh0hqSZFruAhmJg
aDt0Mzjt0Rb59g1RoIBtmjlOmUztuSHFywrBz1jUnzCmz6nxNwhr+9NQfcRQ
Bap1czV5qP+ztVfWhFt/PGcLh7oGYypSEWBTI/iiy5yBGlX7cxR7/lPNstr6
/a2odYOhGD3PKeLiuWZApZGubdM2DkA8miADor4ghgSsdtnHjxabPHoQVUax
VghjeREkZGkhgD4JRY8qZrxbVSedzvsEbYAGJstpd3v+zDaUWaVHiBXn0nsR
iaE7UNy1sOAUZwN7ppwXOiFL9AhBRcsodqxSLKW5ErL6YSc76R2sDA+31cEv
KFbL/Opms8XJfjJODvPTtXVIZwURuvMjfSWY0Hn4vcPmleaKn8HolnH/8a+s
hvJ+jedNFsKsG9yYW37cVqUDC9TmfgsgzYru1o3mZQ6Z0kjIjFUG4UoMtAG+
IsEZfjgSg2SK+5haMpCUd1CuE8fbbR0qg4q6V1Qm9QfGcUqAU2ue7x0qOMx+
9NZIYL+wAO6x+jy19n0CPAeSBryuDj451c42dogvZGdONft016rDWJYcjKS1
U8YGXVrxISov4TiAa/wEZdT3czV9Y9PfbW7ZQPi1M6I6zhBYRz3WT6JQ3bjn
cJ5e8d+FKmyXZEnROkVTPmrGKvsgjWvCtqgP4cdAjZLz+pjNR6vCZOdjgvsp
o4JaKAkaAgVPJQWNvSBNuH1Mj8jzpVyCy+2g0cUtL5YGdvWv7ni0w1+A7nWz
ND24+ZrE1WBCkWAj3jxcFt9WKgLWEhWgL2VM46S2R5vbuT69R2E9veSDRqeD
r1G2RZxD2bHMY6y0qAQvrT37nTR0fruDUiW8plDE0TBMhPKUzcyh/rt1ZTXg
HiqcQ7orxvc2woT2PFea9IB2KCKY0iCuQAOjoKWEOzyvN/DctXP8NR+Db89m
09IQ4BLXuCv4lgewR/EE8cXTzDzEoW7jeg5vKRao3QfLxASajOYHO6ttzmJp
XxL7dBh8/4On7Yd+EcjILYmoZ3Q87Ggiy0z/yXl9G1dLYNILbFaSG4JiMRxE
EXMKB8lgu2+pLUcZ1W8x0B5/EsxweFSxPCaxXnvSki6N1rhQUaNliGIcZr9b
MMoABgOGX1Aakm7yXgsdrTAjVgk4syqSFE9pTOXs7lfb6h+heomT2eKVuZt4
9R1JSG6kEo+7xPuuIcWqMIwMDuFzElfuFTS5qjjs9XIRiH+Od9CunCikI6qT
1MT2nUFOc4qFpZCnr9hNGjUnnhYofw2LE0w10uZ1U9yEn0OYtFGF1itWg3Nc
HxaJ/onNV78VdtEx8yxMUv31W6kjzI0fHns8vBRosD+elFSRcTM8mD6RQyia
E6bH12JNyh0ENwlh+byqeLMSxLbCgaICcbjYD/auzrObLruSyUHBNcVfQwMs
Q2Iuu3dZuHsRrX1Nha/qXKqPlKKvanjreqLKOPnWfEkQM/HpYMlZBodVaqj0
dv3bGG/KMIFlvwQmKXwE4mY7rHQd6Uqd/eAUlhbrUL/PQ8drn/is2gLQo73z
xLKpoXsRHvYsTbDMe47msJFwPm3ZmbQ+gEplADJ1d7HEag6XrKN+0U8OatOa
VxWddmXiTmIsaz813IEbtoo5li9bhOMzqQlkftw2F9tGgB2/L8ktNt9hfUKI
VfPYvrjiwE2Pu6qiM6JeUyD+/TYdi/ExkwqbjQg6u1ehn0WNqMNWqKOPkEP8
Vodb3Ajk1tY/43CS+y5J0rdFh9GTWkFBFwfaPxjKDHIc6jo2eVtIiPLJgib2
KL0LEzcxyYYJqpDAG4z9Wm+EjuXG4oj5QKmDBTc4Zlv2qRmtqrPe0YLdRmak
0zm9JckBt4QVbyj4T4dAhybHkSl8bf35p3UW0ynV5lM6eh54wmvWTY+H9LUj
tm0D+JVDBOeQPccliuWAEJaFYRfGlAvig1UBaRcq+/0/s+FcuWSNNjvQHVkC
nDnkCtZVjbFDN2jCFjxDmDJhmit5DCzEVExypMdDEHgjEoG8tZM8TF3ptkK/
QDFb1WcxYgy65dN+ZyuoLsCfZdrR4zr1mL7QXzP5jvHVf/SMhb9liF7JIKTJ
85oeRuEYZZEDqEBPRntcIhBTdedF9Th80sPzEhpxRjVAW/TS82VBXeYaVEFy
PSKJaJgJDoYD6oJ7eFselJJGkL4ImdaoaVCm4/vFXUC3MXP6lmNLsOrlZ+8a
xm3Juv9w1HZKX6/0X1rRBB8+eDcBz2S8TbtlW+I9IGN7PkinlCWf1rgs01wk
cltFmLMuue+zkfrtdHp1fmDaHu1dsWRXGW4wHJdbuVhpHXOz7sQAwpbBmJf4
MxyAVKxLhGlTpiOzvoamJiD0RmyZtTSpIiSZno0Clsib5e/thkKliCYt3lCu
l+Cq1obqGVKBSFZFOkylwKHM36Fe1WE1aqWNstqgmz3kL4fhg/HNMIAZNCF6
V/ZqjjCBcZWVg6xCg1pGaX6KAwoQFwEpo4W0q+WeQjQs30+16Q8zbgcBH0WI
O+fpiIxkfvJULcNTa04pyfdudyeoXQ4NPLTXN+ojnrPEZ/e7jfS9en0puXTv
ntc9FN4Q4Pf2tKgqZDL5p5LIbHDLCZM5+KeVD/Mk4C58QI7DduQhVx6/R4fd
6gmQuCeEmsODcnNFUSjf/ULyMg9HD7r/LMJFMPPpsfljLP5uR3NE5crcv9MX
Y7l9tlCNQPXZm5b+EhjAE0hF1V9az6Zc4ko84Spx9TxGjJ7oS6R7mpeRffZs
aB4EdQgVtDaCPvWqlU9eLp/6xXOL+E5BvF9due0sRRX2puHp6P+iIjNMN/kQ
2PiaN/qv9ZZ3Y3Sxz5Z/vtymL6vsF/CgTv9+ln5ez29K6Q4ANv9cfwdwc1cZ
fzaaQJbBoHW4UeSXr6C3XNNXLuqvVgAH4afOZrLLe0ytF7XGgg0KI60sNiFm
xC5+QMt4hO/pyKrDsfjoJqX87B5E5YV5a+i7ITcT61CuwIcJV0RTMVdIDVvc
688wUd/0FPdbAKhA3expu8r5NVyc+adVYb+M1UghlXs5lwxc9ga4Z0wVqApf
fdykFha2XBhpxGbfr3D7AXeD+AXZrXgKtLxaoqupaCmiQ3H0BVN05xMssDFw
wbeWkwLgvQXCqExpUSUQzKniziztAterbL5O5SQUC7iOK+Y0DXl69HBmviIf
Pf8G7wiydePTUTHl7LMa4KQMpsvndmkofWPdpb1kVmM1rVE8+GeeIouvtfQ9
PQdi51wEyzC2v/YOCZh5GgDz65N2hIe17ASQjMYVOVuv6W6mN5MLFwPyr+wA
3z40v1LxHHywNQuh3ZpZADM2elBfJpN9LKDLQKHdQ7mXCihlTflbIRY3f7LO
C5UK/IxJBeWFfb88fyudXu+1L0RRJjUfi3Pg4jEEw5GHjKuNBVfJUkONJUiR
N8hJzLyrazSqVn6XU6Sh/yDotx9mYuCbOpcCjRG3mbwn116egOQF0ki4IR5P
K3JvZqgU3juu95jCbqbjH3rvcpT+RWNddOB1GAgHzxQvm9pxYtMDsiL0NpCo
KZPJdpCgarDEsd9rcranmtxqWn22vqWJnL/BqW2fKJIWv3l/dFECvsdw5cIq
1UxfHqZNkTA+0f8NRge1rVCqbr5SbQH7SyqIM4OYDJgYTY4Wt0qwTn7k5NnH
2KKkVO5Zd6QdUCo1NvOwS/TVMS4qL7uqTjpEDGVkaliSpGYj2VOOlK/F4vlN
Mjmq8G13lGmnRBHMeBmi4b/49/q6HrsnEVclTUaepBy3vojFggmbn4cLfhwv
cmB+l341dN25ffjfAvDBKLgB4FWdw2lZ/kMJzpYdsEm4RrM8lS8hkYYR5Dhh
AanQnuRGmX/xLBm2GQuCqW1Hxint2wjYeG5M3KQ26YnLSX69KpiMauF1kzdf
MS+S31bWQFe0gxXTRTiqQDNRxKTsH3L59+KdA7patXHQdd4IICvVRMG0GgRM
lUG3E/zqgM7qFeRUB8jv1NyVz23NBvF/kIw8vVhkFZBVxFM30p4c0n+RnVyG
VXSeeYOAUC1uxIVCzXDbfATXV3CUfvejf+SxDmq6O1cYhec/u37nf11SI7yN
4E5NvWj7T8Tep8HffbYAD9vQ2O+CbdO5OYQW2ZeCo8N3pdFIfyI1KYYYxeBi
ahrnLZH97CV7fE6CoQ6wKS2j1Mv1I4kWOQ3X9vEl44ND52e03dgE3yX0MYg6
l5FZluwOF+FNHBm4yBl/aS1Vfm0lUU1WJiTd1KMRk161YFHRr+JYWiKzXHpL
B8yxlOPvKeld8sh0LgS64vszAm0UJ63a/14lwCWPGByNzR/EZ87nRqa5T5sF
NzQA9ozdVzgX3gPf/Xjl4SLB48Cx+KcdRUiIBcP53wgKUArK7CGOrEmp2GS+
x1+S2WGcB8KdWwQRkSP2YjGDiAmKdpSMpkdVRbvVXyP6Is4Kks37RYm7ewX6
2hvJCCd1CijdBuKsDtgvP4AF7JZtxCPjixIkhd2T8tbvPZPmOrCwT21ccBDy
VQvsEVbTq3aR63/BSottOYw6r3MRBsyWRom1A0K7Qdrypjq26lpqMY0XBS0K
vTgXjCrYEEt7pm3G0CWUKt4uQPaWYAtWrhAGdGX4BdMp0Z0EJYWBFh8RFGvF
K1dF9urTDXmm3vmEggFpiTqUTJULAZEXqQSOrVgpbOVBXF91d/YETfiuF4Qv
ohNud2QkUHJPjZg2wMw5ODtrbj60RHursUuTi96UZ2oVqv7RrksCkkphGZki
U4qgGItNLdWkMtCFue5M4+rujtamOIJee7ZElda/EcBU/cdosJRNBUFY8Sa+
eWnJuqSZv0EJGrCv6xnFYdfl/2wYB78HfdSug/kO6faeygxMvoIgIpZUkxHv
CRlinakhyC5vZ5PQ7ZhPcCPXN6nbelvhi63bJco/rxr1qoG3DYJdq1DVUAUd
DoJ1CHrTeBVqFr0BfF6TAVV31jXe2rF60bmbjIIWQ7aR1NkXgWCmM5GdsgNw
HwlIF0UWZtqRWgK5kPCdeVkYBWwDJP0/IWhIQnbxUQXZO7Pv2mVTlH09AZna
3iSG7A67WG888Frtoa1Ky2qPaw6F4suV3O+g1E8HxzTB5kexurzQj5/WXEdK
gV8F2sLousm1szKViUiQWW5FSKHL83ht5T/e9cK6tY7d88Q1emTmj6gEMO8H
xAPoVNhXVW3w9lhGEPjyJhHTCN7uLAHFRwLHBx5Lp/rx0IgvruDDLjSVfiGw
IPC4vue8QkZ9KPmbtFmhiuAa033icJaxk6kXWcYvSzFTTeYw763kKidWf1Ml
xq4Olh1ofgcrFkS37ym6qkg7jTUdninXBF0OrWLTmEeTE3K1s3f42M6JBTl0
T837UAe6XylHyqrQbqH9gkWhWea5BYVcRAZEQVlGg9L8y5kii3xSRI5mliBK
HRX7iR0UOamEI2RtggQ+czzwxIojLuOUyPDfw4ZJaZ1bOwNpaHOGAB2COU26
bWT2zy/JJxLIVayjzVfgO1r9nYQ+Ro2AnNHzcMqNbUu5edZJ9JOUZjEuBU5D
wPb1vsn08uP+sT/yImxwZ216CWoU5nOrngKjul9OE+QnfV2Ii9yKZKo04fRx
HdAjA0L9PM9rdoBNoPHABrO9UTkDyFDlqeRBFQhpUrrTkMYeYVxISbLEEVkc
y5L59h0zd+4k7/rtvtIAbxh6O00sU43OMABltSFjVc0U7cdEIUTskY8slZ/c
aEpVdiLrnCH90mvNhWYkAPjXeLFeqgXls5nuC1bI9SFBCpByUnwhC5I4yPgI
O64oK/Qg4gRKydK30y/a6T4mlSRpIZu/1VrJeVMv1JRHTEPDh+VKjyUFP+6x
HKCCCMFZxpaO+Q/7IlmCskkiPDBx/1yFCBnZOlBefCXCBMuMJmHuUs72SMVj
5clMWDzi8y4hFt1qjvdZbzz6EjTuBj6/HC3XaUtKZcun2ZG7NklDHntO93FI
u/G/WZrguUTRazceNXwS8c9l2t2ODQo/6v/trAM4hMQjO1KCOabtcQWs64cS
S44tG1sYscYburAKMOXHwq4+Zhb/l3jmHRe7n/78oaJXdwMo/5F07UH8GowT
DJRPulc7QxGA2vmGU4Ede0AXmrzL5Z61/ZS88KtFGlTrtyWjhTh62xC1n4XN
+9DEewjeqmq1qRA1tmAX+4HPgYEvyldjI6+9GqzCA2big5dsEKs/0hM0ZmqG
14OXFiMVqvqZJK4h63ZqL1vLKH/i1kNfvrPNqI32/jWB7rOucqvvfEHRMheI
SQ1KL+C4V20lQThRzs1pf3jLHgXxt6m56Fkyp/EmTyEcX1QIZSM4POW9/KnH
boPSdN/Jw23VNBqxQnxZrNKPVoVkZTDG8cCaBw6tC6uzcfDk6/rszahXh9mO
tOFhrF1EST7dHnt+YA4xMlctw5gm7awNjUS466xfeenDu5aO1E8K6nOetqyI
mbcQn3TZPA2Zd1c+d1p2AxynjK73jQH6mCeOLMYhwvUIsfNJQEUnQBtkgGsh
WQRpuiBmi0vIqv6qXW3rNepwU161jajqDPWyp9bN3BCSgO7logmL3Duzisye
B9ht1BnqNs7QL6X9niozMZECbSfCuXQhWD1ITSpJbxf8s6MNsRRNRzsFfDSY
Tr/6ExP2vuZq1qhfufihiYx7IdtJEUYvxwLA3ibN+jxjiDIUxlcqoArFanhj
EK8z50Wqe0AUTE4O2W6BJpUGGepK1QlIzdTA1HUB6tUxlKMz1mKKZtJ2EV91
ntrbz2uN4vHtTGihQABWQD+xVfid8WgrVadOX4DG4Z6OuA4Za4MNa5Uox+Gw
HEG4+AKiMxEx99GL+hbSLMMoQIfhLTiHo7wqw32M6YmWAvEtzCn0EEDZOdFu
ix8xK7WmRfOQoHS23p+wwG/cYhG2qb24VlBuX2Uh1RRhlBKjF7/QbAtdU86j
YG9N1UfYOJho/mIrzd11zWEMGOlMqr/UOvjZHtJDpqigeIj8gEiMIxQuspfV
QZUbGqp2+32sISnimuk85pFnCTJmq5ET7YhICaxfKjwMOeKSBhYTJeoMz32P
+SFnXtUG98iFPOXp4GX37jtdSysnSHBlKlPqtOrbad+rrRv2+z1rylEccjML
HI3XoOMl+WKjlmbKZccgPtSoCkAQhjvlwNJLjXISBMey7/9BY42q6xlIaM3p
FXoifmC9w2bbhdGMWv6NvAKQtl6QZVoggWJhL0TVlu9hCnnpnWkNYkL7SrSX
uyuJ4SijxV+YN0WukTaktqNFnh0pm0QpS0yN4CEjYIaL0bvT6J2ZDn6mZxSH
6gAmRBl4FbjgdwbfTgOLqz5R1PWynSAxNPQnjO6uutGFCMblbte7iZ7Jb9fB
oAMgngHjBZ+Yi0vQd+lrIlfg02UNLTi9hX1SLxTaP8TiwUy74JqvoYcjBDmQ
vZ4jcTOfbi4CehmC7LzPSTim0vUxZnR2RMQj+b56H9/ne02WD8jBwmpdC4Ie
//9zIl6bB69+tDxFWgfSGyqhA9jW0q0cYoIWQEZOMaKM2vC+gfk9xNHM58bu
YDRlSlvaPxjyWEkiqpkyUqtUufJ1uyBxw1beHdsuSPGg9JJdSzXcpS0sJhII
GGZw6TOt+FmPF5XQ+AsrEcARWFryY0MU5SfUghPMaHaO9rnzhfePBWnu+bd+
VJM7huY7+J+T6oWewHdsdk5Y+AowGxlt0PE9R/thsUG496BNyhT4MuRfan5k
mNcxfajB2m/E1yPJECvleGSq7bluFR6uG8j17ksNJSTCVaBe6oKP/hV9x5xd
hI0DWJB11XEaKn4VLT2z+suf3y+4/k82xni/vYdsZQNIAQ7PqCa45uf3BqdW
RcGcMWbCe7Nj8ux3QdnFo9yZiSTo3SWkaOxZXWjrI0GVxCmytK6cFUfG3Ytc
td1BdEWbPleMm5G+20WMw7LSV6uPEIC+aT+XKTiFSWX3ope8rCOKB5hjVauy
XUipxRFUzDrszSjlF5ZxFQCr1CzOSt+eYGWy/Vzv1Ite7/w6OI2WAaHZRtcJ
7sIt3h22MQQmeFmHunFtfJm7i8toponCi7jAESwrB0wqvqFntlrLgE1D2KBZ
Dc+QumnRGPeY8ezFQAohEW+35Ph6M5rLUXAI/utZVkf35pBfD5ZQs8FqauXl
mxJNHRqslbfzZMxMYOic27CwOAq8VKbKmAahPikSSv9k6M64Z9TDj8H8wMr2
G1NHm/PGJNE+Z7I4lgWdEidoT5yQfEau8feyUDwvNlR5Co9J/y1VfYN9dZTw
jJIHIFy9ENIhtesiV0DMOPzhI/8e+PdtO4yAbPuei4uYMgVKtphrDXYShExi
HhMdVYBY5LlHCBk7ctMj8/PVg3rj6Ca9Z+1gbQTEu0ilwN1af2IHRwPJ6T8u
buflwZDQxLpCPCBxF4hgmQQh4RGBLEoKtXBCSjRWa2pjycGhbnVuNQEpLlc4
5haGmuARmPQuCtBHiBpR26g7vfWMWHoBU1DnsWYujcZLRkdVmwQsL0PgMSAR
6oIbRXgcSofYkVsCLpxMwP8736KKNEA8Fkv/5IU3sfZa7aMY+nszqBh2hnnT
76g9Yq1aeTk/HbBTbExUyztvWB+N/tMinhW7mCTSupTCuKl3nOEb9Mj+WGdU
fwqmvnBDJxuBsitJ07RqlhzzdJOr61kBDZayyK2Y2leEMRkZ1N6ZXXydxBe8
ROuzzEfsj3+xkFnAvOeALY8URjVoqFqAfQHrlcpSBvDxagSjPn3mViixKjUB
oWZL5CYRiIFHQuuWwSEKL4y3ijGZsW6AFp4zTNXX7N86KOXTPYBHUJGavETt
OdKGFprvCoyyVTYQ5mnBdaPCxV/OdYYFE+9cVAuS+3VWZKH3b2dnG5IfgJSQ
FZheycQxarFi2z5WG3Tgp6q+CYLQH5dD/Ah4H+qqKyYxpk0etIH3hshwB5vY
Mm4pnKa36zCI5EVrM5ZY/U664lzN/qBkkAF7dQeOFeODnZTZGKX2kolXBj8M
+/tro7X8K/1m6oELkpeJh3ckFtlE5RnZBKNpw/P5g5JKySoUBnzNmoyp4zLb
TFxYJ4Xzc0dYLvNxqoF1rErlx7bh2D8k2ViPZEDjoOlKxpKzfc83SPAZo5bu
hmKWZT7rZyi2u/FV18y/VhwWaX2DiBXyGYQB/1+X/xMBzjUB6Tyj46UdUcUV
9h2njQ3GOx7gqqnerT0A/1leeLNps0FWi0Pvu+ap/cZFPzrUSf96HDrhTB72
rfIOi+57MDIZc9wwbUftjkRXBP8D5iOlzbR9hOxSY5mTNBpnnHSDv8XFcZGK
Vkbm+yl/Er8VEyDL1J8pCdx3KNT7CPXqEJLQfPxKFbGq+JSpyLQxNqUYrKM1
V0gyUTriOiapse0ZikryI9m8WgO1BXvxS4qkr3CpYXCftDLCTsb6oQ4Xvn2Z
Fvt1kh8llvatlA3UsVan3G+HUupNS/mHl0FWOBdc4Gm+uEH3njsavwRkNERV
anEEoZu7ZuJdGUVCDFgblboRzl3ajPfpdjmioKUHOrcTKlyzAP6tqG359cSv
xuD2KRYU5+A+KTC+IRADKMkd4tstFyWPzxE+8X2zeYJsVhWmxo1SBlkZ+B2E
t+ONDHy2cVn/9hm5eFIJbKO2Wz3pCtVlqS5WDzgDbx/joQJlmGj71J7wSRJx
gNtEJwAwkLntGuao2xZh9KJUdYzbGvyUnMNtci5FEC9kiw3VsR/EniyLK3q+
JfRxs18qiZ29fLW0wuqdRGHCwSQZ2RBjB7Hvm/LUHbJCqFCx4jtEaP1tdW+H
9bmfTT+zPXG7irxoza1UTBMvGWJRY7n/3tdMeiVX+lMJW8Vv5WNV74bY4fVF
Z1R29bZiK/GFULSd9Y738vhlouLJsNeXq6GecscKxB6S1qrGd9UDiP+iDJ78
fL0mHstv4Xa5DhxCOB5sHMIxR5z3eP4x6yAq5CWkp4PP8YtZ2IqaWNBMk+05
2ygTCL1r48VjYjLkxU4IcUTspqfAxmJnk2sP7GmY1N+1o1eaDeLkD8yss+9k
oh5s7Sdhu2Jl2MGBSafOWgopiuUo3IZug/pEGrzkIO4n1nugGKvK5RXOOfT0
qc6l3qrwMtmqU5AtkLOr/sXpIwrv/QW4tcuX6DUTjbtAroFFJdxLnEKuDryr
1cvlnPUabNzN+5K0R/BtQGZfelGNeJtMndyWzYd8Pgb+wrgSxo17A5cm0YE3
koPwl3E3vIEtovjtV5GyDyPHqlf27qAevEbmsYAa4UehVQ/BvMwout6OGXVp
Pris+HDEoCg2Z8r9BB+IOGgSgBqDL6IErakeOQ3lUMKsCs2P8EVvoaHoFaTL
EsZWYnV+ObNyJHV7E1iVxnUZm/GCiJXlE3Ah8snBrGz/8KQbL0NN/Ay52R5u
JkkB7spD+CH6TZfiPWUuFuKh07Xj1KBhSCgP06Fnw09lkpyy8WmtA/s8uuoE
m8aNUchiLdc/254k6YmtAq+7G5Ec+fAjUAvWXfSk4EUmV8ysAWPO+0JbjZgA
rrmTe8Nauw/UtAtb0kagboaRWno7FmH++pfxOoE6PiThqtGg4JzUyopBIsIF
Gj76SF4rrYtN7InHzyim9hL/GjKWYqggk43mabx8sUW21eB2HNMuUzogLCnd
9hXH4+7+x/hvHOPXS6vocCHuFTCutUVmmgWj9RLQO1bbmAUyIWSL3YDb4+M4
3gflFW97tIXwkSGujRUPaA754cbszqghLwxg9OX14VCQPTzvAL5KUhGikJFc
zWDq9EFjBegNx4Gg2eYF+2qbwq3hpV8zObGThbGCi6NP/8f8IiD4bc+6vWYz
sXMIX+MbhCeu10kfOiNDBqknr59xOwSoEDssq86/GSHQ4nwFH79ab4d7m9cZ
yW2IJ87S25ufKPnTuHbq4e9iRyzgihzZld8h1uKz83Z3RzAMf7MHd6EtKJwe
zg3Qn9ZBH/ZuC0bQlUHKFtV1gq9rhyIeUeTnuxxBjNZeMfy7gibZ9f9sEg68
H6k659LJbLHnTaz/hNKn2KkGV2b1bwvlNreodhmZsPmBm0XZoaEE7NMMvFFh
FQgOGlk6Nm9vFdZNhTHX8uzTJPRUUDj7Ezds4SGkKBiINt46NYxky6eRS8sG
DAEK1iH1EPONZ1F/fTg7CJncB+EKE7DAmpHeYTQuT/PsLuCp0ZhSiWuWsnwj
qloRn8hI3zOKyiBmwCoQQwTBvZS7w7gATF8l3K1KJTf3X46j7nCdkuQ9FGpP
hK3G17jK9y8bgxb2ah0TNpPP3ndCdWMauwm5v9oB6RI5DsYiA9zeiZSxFTtI
L3yk+z1tAep036KKeDUjKtk1HBfs2rVFfQ/sULszZxP6za7Qaf51DFc+WPHH
3WTxaMTjFhIvAePyXumqPdpal6pTG5KMIPKIAInvuskWcQLdKOzExBdZA+os
VMKZcflN6uZXH9CbGOeWY7DtSCbni3LewpylP1NeLTVBYuKQEB9hx+O6Mq3X
zxgX6LROVceqgtRjdAaVrr0++HNPehcEG/qPK+C1grIjLZ+5M1PN5dl00DJb
qEeqAlN/2+X625EREzd5fzih3YdycVmRATRdGbe5RQjtYor4f6H/RxBoy8bq
bqN9OGSmwlzVkANWP+lp1zFZiCaXihrti/SyOzJzt+D0EcFC2Hh8GNe7AdIf
B8aHR8XJEeb8h8CXBEj5Mgjo2x1fvSISkcwpD/RKKoBJhkmMbbRUM2gzOmrl
RzJqyfyZARAPoJUgWZF1gPm3NRuOavWWMQCgNFySdfCdQA/TEMsdAlEG1Im/
TneBvSuFclWIgX87Xt8JC0+TmGbv82QGyEwmMaLcYG/AqYm/PQUTB8zvrcTh
GuFZp+Y3e8ftz4jSBPPFQ3vorg83KkK9+ayHRdXggCTNaetytfj2swkPHFhj
fan29dLfuOhq3duDl2b1dprEIwQZ6KOT1/I18WMI1LGaIwzZywuK2f3aK2hu
HytoquGNcI6pof+7EiWOX0KzXtkMvq6+5hs/whk5QYb+3II7pkulSYLhKV9j
hF4SKKY7Du/i23S8P8Hrr/uw2y4xdZ4xq1gqd4Itdf98NJyphsRz8mhhfqeO
qFQhjC5kloD6YDz+fAVM7Dp579JMS9pfD2LzFxYi3MDTk2g5KLVsTTXu4CJY
LF9VtfbgGGEDAEWHBcbX3I/leTY6/Apx3iHvrgSzgqf+ayWehpSSTRJJqkIs
iQbgg6r97+rS3A2dZ+tE5d14s2wyyG/RKQlfzd1BJYr3ONSPZg7RbM3rGybh
s6Qe30TATmizMRP7rKdhWePenw/y36nyp8ckLT//np8bhlkCVO5VR/BZ1Ig8
LRmCB0YODbb11jYK5bxVXegNODEjekZl0Y1as/QuRlye4w+OcUXihwzsfsU7
S116SDD/bwiGjbwrVJPhwVUlu/vNlwmg3AaSPamLJj0kaVgB1ceZFpsJY2dD
7KQDnaYa0TXa78T08Veh6sO1+34SOrX2/ogimzntGhRSHsMYUCHAFjF6PE6a
BQUnGTjzI7lmHkbxUYLqIbDhIgnDAVGyLet6M4ya6V60k2vNJKsFi6ooCkG0
ZRGPfoz9pQwv6es2DU0bFkYVJlS7mPsSPIwJ4ro51gHYgQksHc7ciiSi1Wu3
KN6pxp7iDKcXKR/fwTg2VsN57FCH6vWxgpLI5RUDuuLSzRWd5iGJ86cvleWx
ARF9kEeBP+7gDAoJ+3wMeJa8AcckRLB1CRRqBXicw/jRPleW+u8fDppmRuBj
dgVzsjIGPvsNG/ctFgX2U2qCciSy9npyFngZEKxSTacfdn3JB/hmqZispJuV
L3HKuxhwuXic7NWy7Q6okWz55MZbB60aMYRWI717mr/6PziLD2WFOW5sPesd
/VGVyoRUNtkWAfTfxkwQ5PVzsXAeQAGkJfyPbSHlSiRMirU9s7CY4CYQzNIT
U3Fpt+thtLRdVkTjbx2X8NtREBdGI4PvjxrROC+uffYzKBRFwSP0oyEFqSJ1
41x1QohG8kF7CptII61nHTIMz+eBWNH1gvyGSWdxery3iVdhv66usxC49v7G
kpKG1UCsXvVy4Jy8ed23sYQSv4+gCdYajZDWTHjjtD8XhqdFQX5ljwgjLnFc
NUVefNs4UOQybC6ZABDwKxj/2vvnJ7RctLXh122x7GOE+w8oQThleA2WGu/h
D5iVC23EOH21z3OGudP38wZHQ2r67b/I5rUqY4ZTJPrR99ASSTLgNZr11taV
uhQG/y/06c5eBFOJfek7zIEtLQ7pSj/s01gcWNnvHMNuLjS2mn9mEZOpKDsb
hGmAW4Swj/xzajLA7NCMjKgiUGJMqSHwD84z73SfbyBxvJLyvBnlBSxlFHaC
sqmVHf9ZxdmYpnpx66KY5U8MQmoBywU63zAqEtT6NH6cIpdoD8IVVoZDLJaT
corGvZUUnCairpP+odDhdaOibjBZzt9cidybSPrKAjzUlQPGq+AqHlgqqKbe
nsrKt9tCcUzEBKrF0BO+jMJg+DX2f3AsmHlFRuwAKj+Byr/WTQkAXd6IYSld
mSRPnwtSSR2d26a6J5TlS/oqgAAUkIhnF4IxUDGvnkHc7VirHM1dF5Nuo69m
LORNHq42Ujim6NsXm1qJWUgygr815EMrdadbe5hy8OQAknGPAg4hnVlhHSwu
p5ki6WMvfuEKrO8E4bzofRC5UQc1tnB4HYGJ6tIepdH8JIVoYIoSqQD6Pdh5
vxz/MmvYO52c0pkSvkWUDyxxrDzQhE4KnrsyrLeDRncJ3XdzQoI3woDN8GzY
n1Henq47QFb5DLNNh/j3pDPewzkVERT197dKHA8GRg16yQ3TeMGOW+X6wm48
sxllKPJolTs5fRaf6RSKz+o2jm6RtUx/HZg5DUVTyOBudnvO50xPocG/Ho9B
6cPNaeoGYbUeAoc7r2VylyOsWsIq5UAtu1WrFWSDIkl/n4e+LhNGmiROj4C3
oAwhx1trxTGKD897Ju8xH1IROvLz4IsMAkCslgdGvXJL6jkF5EZiGSbQ4RaO
C6uHrCfm+OTqB5tKa3btVWVHSc9j9KeU0qakvnOKq0uo29h+Dt5Y1r4SQn63
+SjXMi7AZR/BGV2wp3IZ0r73jrm3/y4TsjCVfRy8l5TnJvZNKArbc6t50Zrz
hMfmySKCkBmBENx94AecPvVhFMla85e+AwJ1qvor8jci3YiXV6noE7jyb0d8
7dIgASvc0zcKldtKNdR2+dsg9Wxhl/ovPC7Ejv2xIEx3CgmH6Pa6KEkb1kKG
rAuGHtIuZxgFA29isljB+GhTWBZVSl37PdDyToIgnH+wqUXRDtQmZ01SviHc
PUp72IOePl5HxdcS5I0h7FkFYWKw8cVKqroqDg/M8BEXnYosFwq+6nI+x9Rb
ZMsU2XnY6lDy1PHhy3W2vQRYIbhAdMT0E4fTWlRQBFMnRXuN4Ql1U1vFFe7x
eUWiGk57cPKNUiidCcmtGQc2vBCYuEN7dex4mVVYzq90Qu0wiflShZlarsbG
kcWqrU/uPPjHjq5U/mCj936zm5uiOzjVcGZ9DzIL0j1ns/sI6amIvfmNwGoC
yFyNBTm2VSU6RXW1kPSBf8q6lL5bX4rj48lBBECBqRgtCEu47bBfMOhT8SpF
KG5SFZbdbteiWDMwvv7XS5DR31aaQ7um0x7nPGmfZXMcXLicjBum91u38cvX
pVA2Yj7Gea07yb6ncYe4ztK4sH5LipttkDfHJzVDcol9oweuawvyZHtq5WOe
IAW1nUIvKUZILOjctvKLXMho5mBO/DqDdPlssEU0iVvPepOtO4kABfy6pxNL
I/uKdR/qlGmfDs3q5uCQ+5Ftg3D3f3d3XK1JprWTIzFkhF4rSsF9UYijR3X4
BVLPdlFoAzUd0X4hN+8iTAU7ht9CymhLYgNgiaRLpj/LkZ+v2J3nW1nGegyj
gwJsmmXVvga5kE4Q4Bhr39jfEFxpKSGbYhGeJ/gfSpS0IYw9u+XzLCQOPjzL
CG5/gYft4pDKJK1QGxSF3OBsTOHw2omZCgPAINSvUT4OxCCVqkxsbS3/vFPf
wyyG8zFy1pnWBAESRZHB3CaAvN03PqdVgO1NRVw77loIO9T9ZEcXwOb9LF6r
vM3Ny34qRi1bOIZTHah5Y1UVHxdGtRLx6lozXeGVH5BvBGYG5JuO1NYEHl3r
fjNYLBBe0wxHEIxcdXaL3RhjQ7rwha056qh4Ba9ENpxjiSUwUy4BHbD251Ny
4GxvzzeEFxEuD/jV4kJCLfkwodlbVHBkhIUAvF3c+YgsqxQkHbcGfRfsyvBD
v6E/JGWo1TYjvdNBeRufAj+QJdXTVx8attcioJGgcLDH3Ly8z+2KI7g1NZkO
NNCh73wzdvaveLYHdKvVuQ+qFftBLoikaZdISsRCeWjehu5Ml/nQzJ4OQbXU
sOUSJTDYGM0SeS45lTSyTHxvrlDEwuz8e0mccQmPALTjNTGlQfqgJD2Q2wSi
XAzp718oNItkZ4BsXWeMM3OiiyqE1Uh8KHkYL+11QC/Zj2u4RqFJ5JDH/VGQ
89oc+lvGStwTrXou7tIWSpk1t5WrAgM0ufYIzoZWBRat2QzcvVVEHUhIh8/r
TlypNL/6XW/ya5NyuV0sSav1gsSSIb1JEDO7QW9qyMbGWh5quGJ2EoH4Um5P
rnYIHKAOh385TWYL359F6ccQobkXcg6avf8Q7sK0ec50fdZWJ3/hjom5TzIJ
ctkW+BJz4qumr6aV6ALx3eGFQdTfVHwK/aE+IKEY2wyCyuFQ28Eq/sc4c3fx
f9ERVOJkN5IgEvvk+Uz1KLmYUuc9eaBlOnGD4rZ4CxGfelnCJWOliMDjiy1N
mu+/7+1+16o7bp72SH10VBxH+Tqgohiqk84JZ67G9UuysJpAUTniGHoPRe6V
D1CpyfF3c4ONYBWIO709QjlYlFLRaEtLCsrlwfjV0cAoGYWQkWcp94YC39Cd
tFz4+PClyeRk0eakPUg6SjJCEfIBth0UvZpLWlxon8+lU5mgh9MMrvv0sKia
OaRb2KYlIxGNSO1sZvY3KILKs54JZQ220TrER6xSo3M6h5npm09wAjCIM3iU
+UUE+e3TW1UV6aZRNFjqIs8WGGPBOd7Nf9aiwnuvyF0B7v6Z6UE2gfPFkpR9
r2RPflfuZpz0Gu+wkAnA5E6Ot0pWUY5XisahKYqhO0YjOhut04jfta+10gMG
S49Xn8CyJmBtdabqL6+pnV+UZ3orax8GXsnAO5a6+UqPt/VEnvDTfZQY0PxY
ertcTAVbyTK9jh+rSSoInpjGFj71RqJ5elqrcZ3LLmj4vSy+/4eDEvSPwz7y
tXAsGRGcryi1YWTLfHimXUxtNLuoxxUQddCblii86t1DvTbKACr/qNW60/qk
W9sg75CIH5Nkn3Bxbhst+EPlcTwWH/Bq+xfw9txRJKCxblvXdtrtnkqBpZw1
dQzQZs8SvQ9obN7kiwm0NyQZSqQih2d3A5dOP5MQnmn+MLxML0vasX1VEL1F
NnddpKqYIj6PvqKjzE8FCEsgoaBZjYWgY1/H8N4u2d2Jxf7m0TffXPNP8zdn
4CT9F0u6N1Byjye6PXZCfwRzb9FuFfc34/7Ae8lixggUgxJt27hIY5d/H+Ej
snorFluYhPIwvgw6kj4D/ZNCKFeIiGtRF7oJagV3KnW40BR3IYAbdpxS3d6o
X8V6R4o094t2L1XIBU4BWGeEiZ+EL9w/5w8iF+3SwTQD8hKXvIHQk50+xeYE
JpgpXxo54UEm2AnRB1GEBwKNMhB+rzuIh/MjdSKXpLw+UnY/PKKXbjQFpk1Z
PvA3r7BtVU23J/LFbdhi5/o4q5beC1HZVPyVplcgxPd4o7xOhmAqWzvdOJ53
AzORQEAwD4ZOOXTh4wrB9l5dnR8Uhc49U9q04gBW7g8UR6enxIpOZqHRrPHY
of3VAqWVBI0x8JVOm9DvTnce//0Vm7y0agSNcyR32GJHvQ7OY73vkVf1spBq
mEcCBLMDOchO26cq+NzbnEJEESa9rLOY+vEVELnkLA4t+QqmP8FlfvaUym1e
6rAVc5bqTveQTfPkxSqeQpPp2OGW1ZgivfVrtT/elUNyV32SdPTntNAlp08A
/X4p0s3LZ5XAt/jQ+nplhn+sk7dsFKJEiKeWDRO6iWsMZC3J86YzZoSGsCUe
TF5WzQoKXHAhJGykJACFdH1o2KbOpWBVb4KbUqCIPIMGZB9ungofF9dqt0uE
9wsSa6At9MngNGvHm3Bz9fCB22+YS2JzCcratDA2MdhEhs19WNkreK1VsedI
0ubdCYOX3bkKPnxsggthnyXtYNbRXlGmY0wI9QPOqcpL3ZMfczc/I/OgHb8v
4JKRWh6NhXUxRlFoDeAC702tNcBf0gJP8SQLQmI9YFbNcFtKOKoWe5ZKpEVp
yHaxCOVa6pKzovx40M2WQ50KYPtRRt4krxloV3yDd/itoHBeMqD5ZFl4w5px
dsE821eDKQpgGaKiOT2LW+9YorBWo1YCQbMrIpvwgfkJuyxUymhYRd26/lXm
JcC9HAfmdJ3x5dFN7BQc/wv3J2Wvl4QQZ1w/+3tbQBxd3LyYK7PJxSA53MGP
60rpgH2VEnJcJmguiYtXn+tfUdIz3Un/SuUl3Ewet5C7xrpDooHQ9+du+w3z
Kb3nPRPFERxJ7hUoVkczFU2QEh2sgcJ8r49WS37S5g5SFEuUIoDZCCnmjem0
ynLBQ8DZG6Eu1yiepUyyr923VdCx7MjNUtshh5X3H7R2rgQMdUDjfdlF2l+4
HHDzN3smscvfTzZvOkZ4Ht5ExI33WcCpIIztx3AhyuOjA0f34qBt0FB6n/w5
nQwHCjdsQkYCLxhbHKjz5/WrNH3OonfE40GbXwnB1ihPv3baLJTHP5TF3w51
db3H4CjlMBYfmj+mYQobjMG48gsKq3dXEZb9+dcTf3N4Zg6xncRNrlfAqCm2
BLWYHSeB59hkq5hCpgSaeEawkyI6OVsk6ACW4Hrg5/oXQXoC1eeuh3yJnlx9
6Say01pvLzSe1GdHOhvJszvJNNVd9dmQ+7OJoHs9qivV6CoVhjRFBaSToEP0
bCjyAjH7nc+HG+VOiUzUzsAvM+4tyL0uzSK6IrduGWweaIuSgudn8Vim/Vaj
5qIuwXe7mfyi7w71ySChzL7XyE9p0UUvBdQxgJXv9R47lzEHptgzmPR46rZW
1K6eGGMNfdlFWTH0GJRTlgiNqXvdbThVNOI2dtDPoJwHSzhX0nDlD1Iorckl
oqgmpz3VPhjlbTDLBLA3bhXYplSbbaendFwsAkEqA8VweTcisJxIXJRS+7t4
nNfqQuwVKheDGcY/wrFSQFnklf6JXp1b0QLQ6m81aIpUqIRccJO0pu7LhyrI
ti43QPcrMtT9UlM6UEWlL+J2vogrSGjh2XLDXmqzAbB815akHVtEmwWvkGoM
Iq5we4mD28likCVipPBncVips/Rm4C9lcOYsuRzQ/bFZgeL474l44vuXZnG+
8TLU3Tr86A/zMxxCw2Min2oN8W8uTn1Ts7HjvOH/WGkIkeq9MEhHLSeCnN6u
y00kGp59Q7D4vu5uQMBebQiNaOVZJhH+bySD/IIj4/09J2yZV2DX5/67uAW6
KKps9VzM2+39G06ccoCyIX/frAzdx7LziwXKSxj9CNl5GvudV6ooYjMxjE4c
yO0r3mC9au209FQqSyCCLPlp4aINApnSmrwtx7oo2HXQmieRGErae0rDsyUO
TyI4svAS7pD0jK93kFVNC8x2S3+q2rqgBNpwhU9MmhjCyuVCvrdEg6X2ERr3
O+247zg0VdLPNz26XLMRjoXAA1xSGLSn4Fytkr69hKTizc+xxgHYLji4t20p
YsBNQzSUpeMPHjEn5P3osM1QJB+KAtM8iCkke5U39KbWa6+xHcXHp1p3nLBf
gbJ+rFVxB82OxpAD+oEigBG+H6kLhUQnL7daMo+D1Wl4sG3OfLevpe3AOjHg
+fDAATAT+LFn/M21DyRPTf+HsbKAD/nOg13YrGA2xZHQG2AHZ97mU+WdzNGE
dXOeNEWBpGr+S2B05JPKrWSoemqasAL5+qP8UUvCfgBXnaFCHpP3LvIVkc3E
OAUFBGCF6xZJwfKQyn2qxdb+QI+MCtHpvXLrtFQJ8UrxJ/AQrpWm0SRUtQCx
upuAaGl4bSzdrfP9UserIKyR6EQ25Co3z3TS6p/f0tPEcXPKfYyC11PRDB56
pyc6yITbrZYm6nYDDisvKt2KsfIlbukYNnDdflaqynSFr9aKtIZJF0nhZFo4
95o5LbL80s0MdWxnwrkRzMm/ww6QZ33CxtcUbmA08l0ncRyORgikyV7yMIoc
Oe51K34SNrTUquHqzJ11D5ux45DRwEWY2gHGNlTHL6VOfb/oDh8qwicuNIUJ
MC4+m1ecoEPDb/SEWJhvX72ifEG1A7lR3RdRwZIUq6GM+gQ2CQdgJ7mBevr8
gfE1RfUNBlJ51TojexeEXhQKmLJfSzVG0/JqXobs0FQcu08PKz5nakQIkjG+
9hkTeX6j7JNP+zA86lUiDiIbtStFZb8asIdbL8F8nYD8o+ih8p5d615ROnwT
bXADugyeTFoKjm8EME2JDSzPfNAeenralnE7dUv60F2pvTnTJSxV/Q02WdgI
xJYfMrz8PVBQC1kAv8oYttIh4kjOrQk8ef+lwGkoQs74F+nQG/zxrupMGNP0
l9VZjf4LYJTlsAQweQrrJr1vg0sCYvEWpOZDJfyS2Kmk2ZwRJWM0sUcKubO2
XGxbRDWeD7EUSTmgF2UGrNL8i9kru7A5zY0F98zjCEeAhW6dSMES+cB1zlbi
N8JFCBs5QXO5NRznf7VFX8XR2bsr77ZGb1ckxcli7Ov/VVXkggjpbK0lCg6a
tUN7m6x7QBKwAeoIFYfK4RM9XTADJaZa0P+PN+Ev39edJJtuZJ1wfRU3Ia4N
c3nEot7+r+z7dg0hsslirp6v0hBBQbygSBgUpLiG+luYKm6HfIVNyCy4xvzU
EdPLExLQCYbtXwb8E97jVLDP3VKi52Xr9jJ0d3IiKUu3PLknvZc3HuHeef36
2Nkmgz9RRJWBkenhKxKS/0GOnEPBstcROhiuzTI1B2aLVtt+QiGxuNEdSyiw
7envyGtIMpnMRI0iCvVRB6sDLDhYF2e/imT8eoNGG2HCjES55yefUn4uvdq3
uUoek3XaNY+TV4DJGvFL6dRYmDcC0aeg5mQBRw7cI/dbysyolKC1MXRmW+M1
vfxOYZjHG9K4cCyiSm0CgkTtxJLI1PJemUmOJZt6txyZbbJRjzPbpeEINQU1
ZDne+pZ8IaYsBi0J4inK0liagrkH7NoFZqe1+CbJaDUevlrJVs00xdCaRQIP
ROK+me1IHokojonJuty4qmdwWSkJDNYwugDbfwmmQII6mHx224Mz6aMi6TT+
hPRxZfGhJvuC3xHmMcowrmBCVQiXO2pZfL4hudY6jHj8FLovj740Mp8RWaWY
8i4bcdeMvkLKx9AB8MFQjFh0Y5hkSVW8uCNM/fdYXhg+1U2tMPgkV/B6lEqY
jDtwcbeq1OxiGZ/cPOppXnoj1oNEk4t+VqUVlBg2V0/9Xyn/aJdUItCHOAjn
IDjzb2VpKikzh+FYpK802dYxrwKawQzd/JcA1ZMTy2f8sqUVgwQz3mI7Xa7r
dQYdOm/YeQr7eYIOorqlR9QnJxxVgimx+hseuuOffEfCieLUPAaOQn7hcRDO
222I3PXBSRQtpoXoG36P/XId+1y6H7+qGQe5ruGH7/dCb/m4kE+gawxT4LUI
puRHXXvruehTOKJrYtiodZFwukXXEJEhCfli/kdH/CY5M2Q5TPQiHsE1a4g/
fGYexAqmxyqyQo0Kcs+jYH1bIt7PCJTDzdwGKuu9ZOSqYh2Gd01njG/0W5AW
onRm/v1yxMfs56oNEEwIJ+gxsXV0vQdP8rIfVZYF7aHCPjqF6xHJ7XwHCjyO
lfuLp3wW3H1QxUE4HPngcYI3aSqFr2Zw1SIJ4XY5faHn+5RNtD8xDw4e/Jck
ji0kRQ/VzrW+S1GNFNxl9823T7eI9/DOGAzxfEK60wI6HzjC0P8ggE5TSGGW
fnh6Zg0zGMzHiLodB5K5B0LAmb+rMhtGVkESbN64Fv95JQA6alvM2vHAF/V3
D7LLqGfu+CdoKWC56hJqrcGiKROEnfhDmfv+5vrgJemdDITC+EEv1PZdXHYf
tE6KWwlAJAlTrhacbgfjK3AWC0b3euxdrkBpWJLxYKDMQRurVBjbRR5xaaLW
1NE0+AcqyF7ZjEQSgcRihJMeo1WDsA5HhcIZRkr3WZjxehC5ev5lEzu8pxKa
t6cSUHkmzmFALStALZrKMf3YOmY8HJT4l/1xcDYTwE784C+impTf8uUg0FY5
1gp4t+K4yex+WKw7n7W9SpmlnuuczLyhTkCChZhJywaBsVwtvDl1LZWz2nxI
8SkSnIBTu+0oUo+U8YfCxP0O8JZE1m2W/krr3S+IzJiBovZO7LebZApXQfMU
GS2lGxGpzbhcnLDbRISJVS7vxvIcJlUjRy5V+w5/yvBAsn9MRjEQwoBhHcqV
oKM+wqd4JQAwYGe0SZ2NZDZfI+Bf1VZA/8krx82dU2Eq83DJCc+EEClwYSbC
rc235pp/9lCM4JaOkUg0VXCiVzLuh25OBdD/IoHHt1PuQW6cmYI5koZCQZ2G
KKLG+1YrR4QMkCErZn4PTLosXtKoa/rZ/RG0M3DhhycsFhXlcdCyXSmG3EI5
M5Pkyxm4+W9JFi0IuVMZXbvocpRouXFajfjFFBhWEWs+v4S2wTf7Cf9nG0v1
ov/FsCkXiKGgqMJqf2M4mm4i0P4359P99ezKdVpgcpCCf+rpsGZ71qSSDbt7
UdoTxjD8BNvAks8rBJwlvtKB3rycPHVUlrFANQPEwsYICbrIxD6T0LsKdQeT
yYlK8GzaUuaIu6JYY9VlaIwb03dDm1cXxHFPmvx4scNzC51azZ/X/rtCJ9hG
QSDLqE4xIIjEpMgU/yn9nJ87tca1NDgaRUbnlUS7wMbYgf7BLSEP1vEctIsp
3vwsByKlfM6Xoyiic7iykYEmT41BhOT8BJ6jbNqvrrAlH6cGguatsxxTDkPr
921nMP7ES4Ac9w9/H9583DEGwAZeye92EukianOL775+Cmvcj+teRyjo1MBl
hqebpoJ3paJe7q9ZJy7C1HR+Xr/XVv30RF7F66D0VEdCBGDScu8vI1fXsFQe
+OaoNf02Cte2mNCFzFe4VbJ8lAV2HlG/iw3AEwk/FzpuL3WjjGxWqNjZgjXj
BVCZ4o0E4v4c3u3rIRA2NFHV0jv6fSmN3dovtq9ie643HALOb2ccKtBCChe6
aAK67tRQTWPYTnxGS9enzbZy5HFTBB7EH3bR578K2KB2KFUir+C7lr441ycv
9yMOsuCKmZ/hIA82CgUGi78dFHCus0tK2kWzTRW91Sf2lDKfFi1iwJQwjI/X
AyhZjoWHlr4AOrHsXuQ/XKbOD7albEfzhvcZEk0Dc5XLn8ED/qrxX5ZueZIB
SZX0hbIg7QnmlixKsOJ7rpCEi6u9qcwrfDACjWegP9BZITUDcDwTsmX65koG
FNJCfSYiT1bYBR2mbzyHpF7cXsJELBjTXybrqgkPqu7L4WyfoewvQYYk+mJC
I914h7Wu+LuHUCyzpHHPpzfws7783gAilIHDcsdLU3CCkYR0NNCZqif5koqH
U+dIAt44CveBdpl/TymA2O0jHyL+ZcUh+GH8RubjWZ7il8LqEyYNEqZzVrku
Y+xROeYNkufNVUuBZR58TLOo0wsYZ/iutug7RKm7KicZnNbE0hRMyPodDbqa
gu0s6D62PTdnIVPlAl5iKTHkl4u1LLxzv4JheuP1K8Svm+A1uLHdom73bbz7
2/+u6mAjfQx8D74UFLjPL6Nwckaz2nNH/EhLam8pFIbKFjuLKkyjgdG2PsA3
aD7n8atkEyHEWylAdxiHH1i7JP7MSqgoUC2fSukxtoqoI971Ytyl0q3xhE5H
N+fSTIAMFQikJsYE+BRcgbHuQB3hcSYHFZ5DXgpjIMI4o2uM8IokqR0Zkr/R
JWwilYfiQRl7De7bqa3flrFvieq0PPMALxoiNO7tYHXFJt5ooTm+UYzYdk51
LkTPsYptwaTtPVKD47lQdvB0YPacadMt2Kv/ccFXTyXJlOQ/+6W26CKnpCN9
n6cIANfAAo7U3VOsTsCN8X8X8snO+B2uhlIk9hmoAiP986G2S9suCm29+Fnr
J17Bxba6OO5LP8wLVDz3uws+OS03om0IDrIcNPaRpfcPvs0v0JfN8l1Ia+Me
bfZ8HXvqlXh4gq7IW9ha8xqDrhfQ9070PNq6UiFhtPSEXC6Q0P9UUkkoNPp/
1Nehb8bd0moGwdvrF47iCAt8NwQGwS2h2AeGXhXI0leNWIXur/CLO0V4HS1E
XA8M/Yk7By/Kt4uvTgF/pF+NQfKOpGIAhVE5IzKRt1FePPEXZBNdeUiZhIaz
CGACWPy0YI0ZwxbGIpUU3vhZEAa2BLxtuwCCZb/YiNWk7zX6ti/5XuKOHFpl
2ltEO+hlxIzPc1FqURJJ5Nk0GxWnHGRScz2di9H/xNbZwZtUJn79hjl5L54P
g9c4sn7rAUXPspAXPl0cG54f6nV8fL9XSdY+znFl5CfPumGMopSU3T3DxYh3
bZD1mAoNQ/Qd4cqJAjyxSSh8WFArHVG5z2mk4DMO7GtMvjgRXlt95khoQefx
fbkq4N7Iwx9CwIS7bkYVA8n80zW4eQe8yTBMkdpxw4W7Nn0yQ4qmaBH/RI+6
lXp1ETFZm6QPtUyp4nevUp0LB60fg5QtZYy9WjPLUdFbEwj8W+6/Ri3voWf0
EoaN3KAtM80S7x6yoQDEsM0OHad2ZYSmChWoHreOrj6ueyvIocXPJq6ef+K9
oFlnfMQKIjwX6+tHq20+idbyIfd7uiq4SEJTMGdlGt9W5i7iJweL1hCUiPIz
JVY+yrSu0Al6SRW8x9rlmiMg/hTCFwmCPvVbalGer6WqpmBzdXUq+YZA+Ckc
bH5CUwXlkTPXQ98Wm1gx/gXYiCQ/3jNPN43vlWFLDR0Ln5pwV6RRlJK4nE/o
SX4XobKd9LFTbCq3V1yEqwGEZvV+psonm/Q98YILPO5T4RF0ZA33oXlLHLG9
KmjAjDkFRdJjiJbH7i4GLBjZ573pUhZa6F8ipzHoE69aCIpvKISRI2jnY8D2
bXb+UsAC6IIE3aOsBuLITsmEyRX+05p6jeDWhvcr2XL2Kct+Jeslc8gXAKgI
DB35twGQJvZJ/wbhTzXoTrKtpRPVmfPBVXhhqyBHbhysw9MvG/PReqSXdxVz
wNGJwBhZ2uBV3IIuGek/ZyixFeprQpAfj8Lo/iDKKtoZZmigsWrsbR4/9ABA
Sf+JXFGWYV7oxmaZbznTMM0Ehln6YDpRv/3GxCCqxwwixqw2ItRjVNowREbj
zhYhePxSty97+hKgrB/V7VK9Hwmnv5/p/d30PsCydCPyQ96q4RkGGKU3h7qN
u3YbWZMm19ooOX9ekVjDTUBiy8MEqhBV8JB+xyUR7Qnamp2PsuhafB8aKa6N
z4bNAEg8TaJreWW9zqmb5D3Vu7kQ3GWQIcZAiOdpVKNrqBTF8RsK6qsKjn6f
MpfzcH3z6rapn8UyTkxP8rHjecu8aQkqCv0Qr7VqbZYZyllk3MacVu6p9MnX
VJjD7AOWxsS6QwkW84u9TiUxvcj3pa21Ha3Luf0VT6TMkeLkzBo99QT//+Zq
RItusFifEthn85aArxxoSW6AQxQYzUPy6EMEhX1JpM3faKboY16DiVXYNPOx
xIpMWMc9mNgfS2mFIVVx7/2wCACUCpH5C2qJcUhzCdat2bUQg6WupUfN5Sn5
8UpqSmjlimhVYSexieUp81tE+tpvfbJhRkz98XndI58Ey2mZSJZ7JJQg17Oe
cPqS22TB+op52x9YtUbkax5eANOwjJ06376VvXuGGweOlsNdkvodyQWUC3YI
KO+LmOZ0R3hqir8E7gR0mF/fMoGSon4Sf19CO6chanh2mI2cQ8bCO70VtEzG
CMbVWkKYDKrBrn8y5kkY3XKZXHovZ3MzLKbERRjUwjzUGj7T5hzPtV5n5KCs
ACXEUq//sOyrwTX6vegf34MYfr85ucGTutbWYleHc1IynRCbpC3DWxrAsKtD
nx4es/6trwMKPiiROZfMQIX1/YCRFvdhxExj7gGw79lhBeM2phZbpZHzNhZQ
c6c+0mvMAYqu8NN+Uhr0BARGCLvVk74DDs4irdFDDiY9FdzHtqORQZCT0Bz+
VvnfWP7/LoHIMPwgb2Iw4ZaDQVN3mHh+FIkhYnI1a8mPRI0JnwpFizVf4Bis
8XXz5Je0Rd+poveRxDWRo+37Ri8KvARfC8hm6jWMG6DwEwTLJFw4LivmUtIG
cjmweONZ+eqzmBrV70ZhW6jouresFMB9QxGnYXjxNAXBlLDo+0gMJvJ90+7r
iiQOda4Co/alahDQEIP+iGEUyQ9e1h9HlKeIAKVgIIRCO/7kqUIKePyPt958
VEB6mgGlQKtn2OL59Ab1yVn/sBzoIppDJt3Op+L5lwgRbKGCpp0N+qNNkB/a
0zY5BSOAtUq7isdSm22M3j1UeeJVnQrAbCb3GOm0jlanSNsDS66NvZoDuEfW
JJAPV7KhhU/ER4CnF4vdXvqrM/cGY89GFnzXOE4BBuxyptk/rJsG6aG9LIFW
AHF3OWw/56ypzrE7rfEmb3cQrX9TWX9GcHMuzYh2gdyZ0ucpT2smjhUFikSW
q+MHc3IOUyQHzKm0ghVVtSpTNSfdg7MTY0uE6P+nYD6fx7fMnQLBHsi8f5Lp
eYYUZBNwKUmyl/c1vSP2rSSzb5WPv6iC+J1n25xe8oA266beS53L7931XsMj
fXh0+eSCsv2mCzKQXr0eGm5BUAehRyvPATvLB1k4NliRUL7dKIREgrT8b4At
2BhbqQ3fbTsxMxdB7wA/XzhSy418hwa8H/+K5wO2Aiu81Wi1u0QuXG7XfzCM
SETPV/TgY650TYWBI+m06ePjQieqJK0tn6fjo0CvpVqkbMfInLzh+Nsg9LxD
4zHaOOxHYCpmKYVAfwQae/9dKlmfi5gxjOykhZxeEUW9/oY9AzjTBrDNTUdo
TGF/kZhJHGYhTtuSKnfPAbFVU3bJdJBPoVfJ+owhyqd0vn9sK0dLi50k8Jsy
SyVKi/P7LXGok2+WAOqd41CoUGRAF6fwcZKNnpSErezHzoy+YFBk5Jg43Qt/
HmPjgJFh4f4Ij+Gr/2VUpNEeX5yAYDz3A8YziIgT0T03iwJ4zOMlMqLZCyG5
bx7QN4bPdgPKj+DxSC29Z4POdV1HzqoB69+kHQ1wq69TmmeXWGaIDV/obvCq
1fNNi9+/ErX4tXSUwxz54/OJ2Olhk9V63kpph3Zsf+4X3bhFXS86nnnCAlq7
uy6FiYTx021zpLidtcX88Boxy610qakc+DFo4r9MhNzHxrE3B4A6Y+uxHZhc
5qmLOeXEZpqIcgV0dNBGPlrZn7jx4CcaXlPbYL4blmXWYp1vfeYMWYbtyVvR
N/X8b7cbdKCDecnFCj4O+U3A4Awyk4URWMcrXbbzmUP1pf/HRJ240SXj00TT
2OhDlrAYkPH9xcH6f0r8z5OlHVJHfih01I7LWD71dvXvEvXZUzDDiPe5/xfn
Bha0xrHApK3ObwEUtVA5OiKjD/27E3IPf7eMPly0e6CXSyjpVP6eeOtOuhGE
Rp0LAg+YgWBZh+d4FOcWvgjeHVW9rUoDVgExkUtzw/n+pdsV9MS+ZwM4sxAn
ak+XZhyMTFVd7KbiOq7KLV8xGNGKI5yqBQd0kXswBxLDbP2sUdSuIyJ8hxcs
20MbSFMyUQk+Up3UP9H/H2mgrHzLwmwAwG8XMU+AHGJnchbvXfDebfzZMvGN
pijYNoO7aauFwvIUKxKLIkfi6Ik3xiqKky76gZ651bViBCD/p/wAzauC2dIs
Cz405QXnsi5nR08cJYe0uwj4sL1GntxxLl8PIK5YauikFc9z9TEHG/SLLIIA
hwOyiiJfyv4Obu2iJ4B423EdEjkH4HPt6byyTh2ElMDaaIlx533A44eC+kWj
renrNNsD7qwf7g2BT3lUNvYQ7aC9/R555gyL8uM1u55H+tSatlmvhAyY6ma1
QGDBTTpzJ0zjgwlCGpLHLpP3sS7ZQn4g6Yd8Lo/xNtczHNpHnE9CvlEl2kQa
jVUDmznzLJYwxMX+39qfA+6gkHWvv7+9wjsYceKOtZTu09mcbwKRVPOmrBkq
nYprCrJ+Lf/X6ALy26JelMJ3WMJ2+wL3NYsDfJ8DX2K/lNKcfdLgJSkkkRFi
WMmuG/nF51P4lQGH9sl++3JtXQ+yF4WBZ73E388m47QsuwvHorpEsCLMiyQd
HUD52NOybOVjlTTOka5pz+VL4c1CMqicefDBANji2QbuK6sg8WPhTtmtxodt
XRTewXyztP3EXUXSSVIPlaEWArU1S0l0f8SjAzY0tj0SdHVH7xqwYDU3EikA
BBAC94fOk+RdRG7jFhuCNGmCDbwxiUkvCln/bblRxpAsGVchjJBYvte3JX+z
grwOLmf8juH/dzp1wSdtEr5OZYmuHZKXZd5IqnBF++TVTfBygWY3JXZuZ7KF
cHFfVwXUxlwZ0mUz/bSYczoBSh+4H6jqfFgtm52vRDde+9HrT+GU4DBcN1GH
J/H/Wu4Er95xFj8dw8yUJuIxjbUaVaJq0G4QToGscIvay3rVLgxeM/2NUHVq
C05tkIBFZoh7gjzmr9UdreXXzNb88MbH5ihmam4xU0HImGdxJWMiL4HQX7Ns
Ibs78NKtAlihydkrkv5+2Rd13xNsGiL6jrqyYwLbAAJN8189xSVcRizVSZEg
iQJCUKw75Ysfo15NeLfhAKvb5ca97qN0n738C2pT/05+l+iwm0RVhUChUgYy
GxLOm5gvGfrC8rsvpJ4aiplHJ3IaQDF37dxdGe16AD4XRyQwgAbs+AIg2psc
yHMaqU17IFaxex6HUlhcgeIq/czAQKI9b6HhOHEgPTTUg2aFq6nL2OXMGYDp
oZbwJCmjj2nI2MiZqT8UaSWHsnHi1KzOyM84I/pt6gRHQFHGhJOhop3VS2Dd
eOMT5t2Sm6QtUJgnZU0e0E87AxiuFdj1t9+fyW61H1qy/RXmkiKyiwgIAueR
/OREqB3EMAmkhDasIGlN3AqIPq6IKKLk15HGd/TjQJTcj7KGLQCCGbUaXgID
7J8OKtJ6eTBQnVduwac3zr7rkydy+YPkrL7RlISqu7G/0/5oYxglBAtyLN/U
lm7TnEy2OJSxayGgfU3ViMnN7vjZTmnk4njiF2dWswyCEuyNsaD0Otzz69Go
ou056EGq+hLiPMcwevP+bNMV1oPjeqPAzA0ogoMz+c3IcDrJxQ7gimdreo1K
sc+yUF0uZNMPgBs76qXPMT6I7XAjwPUbQyU87qCfpBGrGfIQLEx7siuD4q7g
Re2f4X/mjqOx8pqdaDMurAR3fTeZXotFJTBSZ+1PS/A2iwhEtFBTK1nHGxeP
f6r0wQca/sX1uRfqjYYjMeUVMOKw8ff4LPWn19edum9skWBXyPh5aedzYiv6
zQbC4vAVhNKyEtlDQ25xN1ARvWDvcOYjxEGazfNNCEqjRD6SOAk3zSuqGcV5
qaVDBUVQLNL+f9RyxAng3U8YKpVzQleCTXDo7845eduDDJ8+bjXpJ7hu6Tbi
m0kkGOgPDrf9t0nRpmPz/+xnT6E74Jl38lWG68PblnbJfy7/GncQeiWd06AZ
lUNah+NlWYaZZdxb9QBbimHb17PVc+mxyWdNkfWGkozhk3GfkE/rBdOfIxrO
lK3msH8L24lC8df6wVoQa0wsBn5ntMYOgRC6VAVwQnDCwUljwoJZWjnu9GGX
KVYz4qENW1/ySjacn0wqZ2VTLrFZMQSRVzcVsg1OykAm0n3rBmubVV8wqgwe
0Jz1lUXeSMQ9oN1EpsRjLwrf6kY93k/FsWRbhl+quSsQiOubIVXd56L0HOMG
+dEWhVI4KI81AdfQihyjix9aqhDk7rd30NPKRULrkpSDmLZYo5rp4O9muyTx
gRNEhZ/DY5RMOlI6hIRZu0LZ19PDCdjBzAV3dLJLTPTBdE7Uj5oqQGBa4myF
+iy7FleiiGZbhgj7tLwfFNIdimMejuDSETK+IKfHS/YIEIWIPNjUCnzssYbr
IeNp+sBvHf9hUw1Wc3024wGaPKANK9lY1HxL7Y2ImomGNQZQNnhXZWlZGrPs
XFa2FNzKheUoEkZshQbC7mjX5lTrdnNLlRFS/St8XhixVPZa4HKLs7ZPBvGm
P9dGXpDUj1QNrTGzgylAsE7dvbYTlZiwDu3zu4mD0mDW7vxrbA4eOsr6LRIP
AofaQnxlZvLazV5rkAUsTxAdk3OrCjscA0jm78PyOegsiVRpKPqNo5JvL7aG
Ga17N8q2V8yKHT0QFgNdQY2wN87y9ZYY+ee45ne1CWUDcHRIW/rp31sIzu1a
uupjl740d+FhoS+7exz7XE0ZzNlk6B1xiTjuQyoB6o5DjOS439PXvDodADRF
Ntpcbd3jMjjYA0DNpgJ4JF4kJ05cUUIZidOWGVWq5ZRXg7n9jFxYvXkHTEsh
hzCYNAj7u0i34SC7Noghd3mfvJrAFDEDDFj6teFAlnMNjNmPR2BSIONemxqB
IE8pgqie77DpXlx4J26oct6ScEAXABgLDb4tiCKp/PbbbLva+ddHPy79zGWI
3RF2ySDMmYonVv0X0YPijXf1ptOiocZgf1I0CBev944gf/sFrlxwSvXLqkMj
n7CxtYnSTxSqYjX59z4msNUS2LzTraLMcMmHF3+l3Q/iXz8cbwKEnzZcRnM/
Q7VNcwTk3ym00DQ2OkkiUHuyQe84opEf6WvWPWL4Tx+lyEOjSuV/8FY7SFt8
J778bS1upSwLuFUxjHyqzctblPT0Umypnd5sizqaiGxuvjOgSH1WnKxqWL53
8vhfFxzZAIDu1GJC6YvRPmhiDLk10OzYfcIZKyWxnrtx2ntNZQEUIoLZ6b+x
H+3ZYfEvkVpjxYi5Nz18k6oPq8IrIanB3fHOXtGWObfAyif+1lmqEcIKGYyZ
f6eathErA9WLgnYB57Lehxgds2risQ/F5+rIXYahgplcJfgSNBt5TdMj4Cqq
IeHpckx7QTGAD2T0is4/wjTxe9UB2xMviYcO0LruPvRWzsXMobEr9G22AgT1
eTSK4IVRJKkMs7rpugKpTl9llZ4F+c47dLDYVKpVsdTU/bLSvj7QLK35OpqQ
AMIoNxw7Q7E+KYNcj7Gtn0OMqwAklLvI/2aae9+oP8VIHOZQzY+UbysWh+6O
h4mFgqiK5aqI7q6q8UdSkC3gG+pHESVr5kzVJDReT2i9iT+DtPX7wTv/V3El
fyoZwjHmQ6VxFHzy3nODq7SDL7TLqvDc5nfw22Ce/pDI5kViEW7HR+IOR7cl
ps1te+DJUVzJ1f78KWAKbGuWguozrErZIQ/zYn2SNyF5tk0w8xxeMQbIqgfv
h7IX8JXow0FSX3Hlhx88c6MAZwIqgEonCDemplfz7MRkFV2cbM5InSC3cGAq
ZGYw1Z2XldAW8FRxKgE3nL5q01ZvmmtN/TgH0wbtQbfL3+C9xHRLjNAu+SN1
YsaNYYNAhmUcM56I8EI//dad0udUIqSSf2NEtq5W52Mh2v4/n12HSo9OaOHU
/JWix5gNvNasx7ZPZF17PnHJsqeG6/KLePv5rpm+zpOyRtntq3vRLIXMSvmg
Qd4pD5fRQuGCIjXmqLFveLfWZ12OfhnnQxdig6tf6WtlY+G+0aGt3gtqUmeo
OZCMt9lHvLwkBkMguMH9IR/+HTgcwbfhoKga+MVlH9WG5gk/nqD4mLy2o278
bGMOq4nfoOF9HPrtrKT3sFWIfIK9k/5Aexk7lD1+FhDJ23tnOUOqzmvppdiM
pywQmIKcFjl57cNyscZeoQD8yG9yVrTj6NXCxIOu/Zc8dzbMig5w6PAjgGwK
YriNCnfzPSuTFYUpw7Yud2seW5a4us/e2Hf9olNYdb5DB4w1W1ZM93xkrML8
GwX6dsOKCemBRpltWnKl6t2keLvO3FQGDEHS/AHTpmJCRgA73eajKdPkj+Bq
uvC+a7qui0aKWhTu0wKZjQUOJXkm8mIMA26zlwEGxsB5JzaWBAWzqN7nUILI
9sWERbjdHgLO10xhh0WM+DwxUsXb6oV2LU6ZhrpfRQcNaccnZhI2oUZ6/M1Y
rE2oa/3OzVXLht7Uz7xLjckOog8ho4Rw3svG+RbsUrk0hf+CcYwEvoYieOmW
/Dw03qkmsJIvXO5FS2ezsvAw1+ToR+YxdH+pMoEBKxsN3K90utO4E4cBMmvb
jj5RqEcnE5/gSDZYYIWreLa8PpGATFJqtwvsp4820dhvEu6QGTIxAgd4bxwA
1px3BtCLPL0IGxY45BIZoOavORMvXgzlXuqcyVQ5gz3WoVz5SRliA6Le+IzK
9kPV27f3e1lSftbDSUn541IG5iHNplCsFn7JqOkLtw1PBPEJPzFH0Ri1Y0ud
a6WOG43qBw05tESOSNnVSGshRPS5XzSSDmLF+F1yhYwNA5OYiQElKO+1WDHc
le/V9LV+cPaRgshTtRv5/SKrcHaDnCDPdBaiH0jPz3k/7iq/aHQZ7dPozy9n
K5/HNt3GkbULMD/ZD5fe5gSWmMCbBocM5ETuSd+scbLsnGQx2UbWqt7mKdWs
IWF/xoGWE/N8rIRxST+c0DurvbK5Jwb+G8oUCOrQ3mBngUN1xIWKt5RHdvmS
boAQT4FMre6Z9KfXIoPzhI3z2aD50vPXftCwxDo28GoYjPHhzzW1HMK85x/z
9U/MWHX4q0FfEky2cLR8bCr6bGER5cI1OWnWRVekHY2l6DRyUkIWbugrCyza
gArq4mhpbPPIrrINKvHEEhqF6j2rnKhFe42/FKCxO/DJRyiXiwwfaflAmcyX
u26PE+trkYwzKg7UGz+8GgVjbwiu7u8WlCPZ5JZHfyJfnyhkvKOxUYO8CPsL
3ruztzZohMQVJq7oGzE9m8mhAD531AC8oqI7HNjU+qNCtTPgTb6EumEIoFN+
HrP04BzlpBNk+mFg4xFB0+tvlP+aN7NEOJMElnT9orMwy8a0Z4hvKU3UY8z8
6bTsCrBpU7ZcSEd+MqQnl4YEKcv9A8KG07g3RFiHM3GhboazolhHoZKyym5r
8pZxeSFrP2V9SizubJ4NR/At2N2zx7VKv72wF43RmSJVnH3AUS49qR/cD4Ot
ESoO0evY748pllWg+txDgXx1hT4XcV6/KFV8ANyn881nkDK4oG5eaiPAevkp
eo2EaEQsHVY3w/GUqxY8QObXvmyLalbdVrDsvQaJ5ttCCV+0g9PDbR0mifbU
v/p/gn+P7IxoIYayNwveoYRL9daC/aK7AYcOVsGy9hx19auBYfm9sd9Emshy
pnPi6G1IEf3viiTPKn8o+Pd4w5vm5jayw2eolioJ4q0Jba3GSFk7RRHpvnBB
t7Ysxc0EVniHoqCZABGm250paYbo8uxgE+cwhv9+b6AdE7ikYQ212hicOSRp
qoOQrtgCsOG7Nnu5cfrnE0jCEgUkK/Bbm8piBHjlj5RP/79qHH7wucQBQC/N
q6c/wAvz5W6iVo0V5fpeWy7TNdP6NnY7GBooTkWqTe0tgHwqRxy9PHz5qP8D
Jmtuo6kwNniUwmnK4L4VW63vxrLIBVQMzfkPTRd67cz2ETLH+HHwjYYTVjXE
iCPDVNYBh7hZkdJxXtT7j8Ij4aZQ1PM48NJVznMPBhOxpebdaOwdsQSZF+jC
FlIIxuWMmnCKAFX4ST/eGKZ8NYudO/R8Vh5gWQeI116pUb3UUQMiZjeILCCp
x545UmjVLBqfSR1x1r43L5SEO9rQ21x8sX6D7ZW1s2lW6bEIukRc5LkGuaF+
LnZkiwMqnecnGZp/UegBCZxj56dVY0IfRp9Ak5hIg4F5plZEEGHe3RMQSQM5
rNuWwJMnTAuzQKsWOA20JbhR+sBd4URpNPfMBaaHaQ2KRvtMydn5AfrPpqkD
bXOpPJk5aRce0+cR1NgXNxY10LiAW7C4iKqTX9JrvZ2x/BLLiseNxUKyPBeY
gPEVmipXnUKyfitDW4sqVAJgP/BaK9Z0qaq4ZWXbEWc2drUCM1B9oe8XfWD8
07EWXZnmpDdXCp6DgrhXL2bOyACgXNYTrcNNlUJ3+P6VxsKHZG3PwJD3K69a
6/KE8aYTPjLFUsEGfzmEzgZ5MYN0m5qugUBdHSvek2tp0krTNOMMDnaTmipo
L0owl6mnn6BMwPrFxWTwVe4gXvIVSvEFPrn0y2xPUoXA2n/G9pMW7/jEHF4I
A9hTk0OzqHmklugGobhVRIbAlha9mlM5fLJDrt4zAw34SDS/Y6DhyzG3EyjG
JPEITVXw3P/GTKljk2sq7XrHlGiaXOF3IS46TaoSWlAin3HNCiR1j7z9j0vk
9V87T0fywE95x9raLVYZOqapAJwYsqNYlMkpplT4MAFih6TKQun4TH7bPuBe
qdrwP3SIS9I4awdPpgGT/gHToXw/U73zTHk2dIOnbnTyxNiqUkatBaUigJeb
jPI3cVQF26SynggnddPI2EkfYdGAP9145izOkfp5h04KER6P0K13ug1UDaFV
IZPaD9qj/pZsI3+L4+U7/kvl8EcbrMv+1nKyWoAb3+DhNSTFE3V+wIacthT4
I+ka13uLSSgAzxZqK4T71s1UhRK2HJ8UTCnFvITe68I1E9bXND6XcfoyXe58
xMVTIXIAnSO5CDWAG5bgsAsYEbhKI4nzwk7fy1hPa+HyXC7gws+tgIvRDU3a
bUpLAOySMuDNdny3Z1tPdsxQAZQGA4aXQnGA1Rnf53DqjwGYJPS/wYGq6lcv
IU/MflyzXJDJFSgMA7WYCEEdX21aBUDYT79p8dRoh7bxa4B/kmhlWSExDB+X
3BmgMECToEsV1A7DO3WmErU1qqZXRbIqOWwc8wO1RDpNzdLod71+f03hpI2y
6imepRBhJs6eI+5u12aPdctJg6YhfKCT/S48c/U2oTlX7RBurUhM1gXkBtOi
lec6mUKRjmL/UkBbZjQloGKHfEQQ7T0vC5oZyx1GlqPop/8yH8toDtw3Ttsl
q5I7ss3ysgi3v+vdRr2uq6lWCwQWdFLOXyTq41C+kOvxBF2IUyz8dUBJYwKK
yiag0L7bKxtKKqNL9471HRlUhaCeFRoyqMb/nhC78bazWQVeuWlAYH7dFfoW
BgisHBYwhtEaHNaTFZ5UbqIAaQkJfgXlhGb/7tBQzJIX0/WO49D6Ck7pDDfe
cUsfyyHrORh/pPcC/BIzsQYtYe+7offaZXILG9BvkFsSxrTH4zTq0otcl2Oq
y+c97Ebwb8X//UpS43YBeWZp7uJ1BX6DtKQFwnjCfEMLYBP1IeKK5zbIPiC2
/ahRXDSZAcqA+xZA6rjOrFZcp3sIMqSHIJ5y7CdLNo29cvfAKxfQsE0BgLVZ
ZnzdFBrlqQazXBCbskRbvPq4lP4XqOGhqV0dZCVz4q32CXQx301fud5ep9x7
hvr/vRhh8jzT84JU70PfUxPkJ8/LNB3kk5yksOPGb1K4NUJ4Xdx+H1TpOpH1
3R0/67+WzMYM7JU2QGfgufh0kYd8GgmpyiRrmiUu+7ZNqPUlY3uhDNBoBw6I
SaD8uyaaRZMgDmwuyFOYKho7cXRUmox6MzeZCxerx2p3DA9sAJhZOvoEndl8
B/VCvrDDSr/+eEFDugeWIQOTv8k9xdz9RCHhBUWf5OgJhH8TDmIiiSP6L3MP
raiMCZPbjSbVCLDeWjtAHluPFjaLLTe5EH1c7jGEGHHk9YhKq69mWHPaCY5I
a8pX9h9crw3HUy8N5hzSTocPt15arEccTjUUObnN2HQG82t5pcO3114V23Lc
UZYcGf0/jdTRHKq7zWY8MuuVYdhv2m1N8ry4Osyp4Q4hgLiM/aob6UXNQYbD
Up7/DdlCT0r5azuRCG8/iaG38k4UOnf7olLNe/k+2kTM6OEj07L9z6p0Zm7W
GTTMYRpJJohi7x4J5Hn79FVozTCG8zjV2jD0Y/4cP7Uj8Sc7tPRhMmbdrBPc
tD9ja6S6A13+yuaz1EbcxGTp0N+eb0A94Sv1wTQK6ZD2TpaozR6eai97SIre
xMQTzBz5IAUMDWOK9zyIwfBoLLJrJgAMoOEZeFi8k9Xk30WjHzkiKCkyEGiq
HrqeHbRWlc2FtM6b4dH+hGajNnTLwyPpAnMZ9dnaDWkL2FSn0BkuD10Tl3qY
3heW2Ctt9D8OE0IiwFNPRW9eByD8siMkULnkKQpMgqhC6ShpVFS7CZJaxVhH
UFGBacev5k/fYghlENsb77XXHpCLGxKwS9Db/aCro84QAZA1GorUvVSsjG2T
Nay+G+1p/G2sl+DQ1bjk17EKlzzQ5O2Yu9fz4/kJiGz1PmImbTcSQlqb2ffu
edEZpaWixdSMEdl8D/imaNMe9TzDwce4wyoYnO/FOE3uG4pYXvrMjupG8nxR
ooUoLy6Iz46Jv9Fx2iaFPo8AP3IxbT4PYyyXQ/XYecNF+ez7ji0beCsLpRxM
YZAnY2tABMgbNb7+RYSPvhzsXWhSvUSDV70DwWFEzsdmDuHy6jFTjBgAnpEb
Dn2vMVbWLr4CYYSCIjRXycUV2R7xGSfq8qEJWziQtdfge+A5lcnTFs1BiHSx
7iSAomEM19Ny9ghKfteF1SPe6kbX10iW3wfEOSalCQnI+rzcjJvZl1WJy/ZF
Zc9NjU+Jbk6Q4QTvBT9l+q/Uvpdim96nrbUsyMdci5k/78kOnVXf4Ngy+zA+
qjsNbkuZJQu++k77gHKkjrhalN/iuFzxwcGohmLdvUYeSQLSy8mYaExWb7l2
wLX9sAK86KhCJ8aL8VECAiSF2b8DXX729munfXcbU2kKvI4UJywL49qGYyTS
bVxFjbuWqw+RHzfAZ9A722NExkUjiFtv7+4Y9bzo/JRL6K1FWV748KSb0d+F
1leS2ysKLC3D4tMHkhlF+JPOWV1Gp3r+tA2zYaMXFXpy8zLcJbqThVbxWB1B
lwqY4h2ANpbPUjCDv3ojjNiT4Q+gi2UIiLsTlNaeDWe7jIPtSdwcncx3V+ss
0i0ZdAW1o+q4rqI2OCUIwhww1RgBlW+kt3evGCT67yC2ytA5nukZK5fQR8aX
W6qYAA2nj3B2QFhk3/LkCC/IXleZb+8Qo8p9ySReNMt7HKbhs01sk2lV9PKW
nbUokBUw/gnmyXbYwOkOjeEjhTtOD0caq8lstdoZ1lUyzGp8fzgBSPtlGw43
L/TFu9IjfXgths56PhQB9EyAsYWJjGMxzro1VR2U/91SkorbObmewVvg8ksX
e7ckRMdOGHHHuX0Wn7f7cscEW4JlK0zpb0HElb9QK9oGlwK2Navrbxxs7h5T
XxBaIkaLW7T4SJHiRZJYJ8SOdICSYoGPDmz11MubLiq2yVqoy/5//5PWyh23
A+fYl4xszyD24G3UcQqKNTcvrbc7kys7VX92n/pIM4RrbDSZFLNvSh2Pq77k
pLWI4cxAgW2jbRpOFr+wVuzYTKNIDjxTeUjQokF2rPwohWycGaI2JgAjn2Ag
GmTw1QOicn9/j9vCXl6siTbUh0WLfYI/mFqBQC5l/csTQOH5a8FBxeY/15WQ
aSdesq0pUWhDbPTonDM1AHR/rHie5U27S2earLvksHt7d4guMgoqmpyvOT5K
2c7TeJs4XzRjOiaFjkT/uyWAgTa65mjD71ZElDcbaIe1HUQUt16BMBgD9iZS
1Neg6DZZAyMaFvJboVmGTMF9kVe4AnERh9lrJ+UYCKD9aMbAljV44zjhwUOq
jjev5kwpAs1oq2iNIunvBtr4KWT9Z9nDl7+ToH4g+fsikE4zBqO+pSmG6yfu
fGIbq1peoZN6Ft4NBsj78ArjrTjX2z9dP+SlgONbPvlY6h3UHpM6M/ezsrEW
kk3VEBdJP499H8GunjS4Hhk51YUnBK0v5OwW97PHRTqi1WQAAnX2thKqhFPt
0FH5ND5TGbCu7HvCUAM4INYXz0cUO3KxtGD0Y93LM2GEBM1GKD8kJZBs+bo0
OMI8R7hYFLbkS9PrA8GeOESE5GiS1vrMSeud/tuzKbB2glINQHVLsdERCGcn
PqCGBAAj+IXC2RXH/c3RloJy6LMFzcxZIs24srFAtji4JLzEAWxQC/hi//8r
t8r80ZwNjQf/hKI18Ga7HlyeT33qA+MMYNVjIg50zJQe45/TmpU7bUdlUYAf
RnzB/aBMtCrxHlK6kAOC2RE/OVTURHnhcdzudxTpN7/lTLYkN122oKT1I5pi
fvf0F+hHQ+XaMSMw+FaEvbbfjje7qyRMVGdPRVwYs0qj9IZS6oiuDm/M2fEh
Ma1fZomaLuh/bLTjTovke4T0ihwasfgF+/cAJPFpwHqJm6MxYYsj0/M+FdYy
NwQA3AW2eTDtyu6iTTLyLuTzKtqKZVjK0ktYifcATAsJs/cAytCJDAhS63tk
/qnOXI4jvm8ElsyP/q7z6LzeanpozudaOb8HvRw7Fx55pHSirCsyN7yfGv2L
iDMkyPblJb8HgQXMMbrlyEoo0TJWUAmJD4HsAFUKzZRUstO1XnBZGoLVQuRB
JK8DURt4bKVMIk7nDI6RlG5ZmzSmYSpSWpGlBUMXdQtS5ePYVNQHhANsxjYx
9wUUYbO6aeeFueclO72GRU73nfIo53Hi2bXu14L91vRjvhYMzXcuR6kIKVjP
q0Jj5PEUUtsLxJyqKKtih9x07tW9OSMLFUxim/LbEV6fcRUMRiskPZ5IoGkM
bdwkUDrKT8dp7jzxu8hv/QVW0JRlhQw6YVOaXcoxvlKB0E2fz1Ypn0JSX8BY
UdaaO8ewxtFH/nB/SNKg4v2DKmlBZ/yZUyhFrurNFDzYpyoxuXtf/W8zK2qe
907QnG93InXInUr/YRLVl+u21TBY10CSO07L7K/gGMxkhl5pXEsYaNmOMzl4
oviXRZlsua6RMn6KkseX5ShVKrl1lOdnIuttTI8lwsltsNxxvpDvwbTNZHt3
3RzR9uDE/Q4vX2oGzAMmn4dDgKsNHEkOLeH3krC77x7DZycFdZ3EuLRZ4NUT
qncPBZKc8khGtJ0QVWXQTYljWxO5tAyn2EYQ8e9qEm/hKpb8ydKcwitKDlFC
PIzpIBAyCpJNSw5/wixW7wglD1dR87/STmUzyXm3wZ5VTQIFw2EfbfQJ4kPr
NNSX5xEmWbD8Dtw2AjURvxLVnhcKMXETqJTMHh6vsaicWzIQejKJIKN7ITnr
J/45ut1jojJye2vIzPaI8gnx9CagayMOjsYQG18cssXFublGT/ZcwjXWfIcD
HRFWR7IA1KIF1rHeR29KOZ1DyL7i6EY1OhQHxIvAqiSUYf3hWdOKCM1l6vue
SIOEg58hJJgZhglw6vzyeKGhj3veFnK1NiqL/rs09bqAyUv6kG+Pq5hYQPA3
vCStazzDp+f+7iTm4kSoH4kwtX/uVdyMK2Afp9mDEO5i0Cmwp9lyBxw/V7H1
uu1Lgrfoyo7OjUSC4i2Lusmvuj2JpzB3Ey+VV4PLZiGLTdoEVl7RUnQYMSmh
EuO7+zAJ1Zc8kQPg3SV/3u0JDadUzi5IxY7X3mhkCUSdI6IwDfc3TogkcPzI
LP0XQSAWI9zUYZaMR6JOCKP/R8Svt3ISFA17es6SN/JbsKw8S2Ih7mOg4Te4
EYD7PIpoyS8ILE8Tq5or4pkxrKdoudifsVKzfFBI7w0VM7QOk7//5vi6rxih
4V4xd0AIHU14aZyeeBMv6gdQSfTSmLliZp0kol41BNOQanB/cAQzyUdXiL8M
FAv0gxaqbUcyIzAOttWCNvVSPC8b3/2JqmAHikPPIZXH/c57jBZr3aZus92d
mpY7bZTiJyKSK2YiS50IvZ35ZlGRpPX5FR4PYcBkXCBeOxMmuMiQPHs2vFaN
HbyQFQiaikAbF4JfKRo1HyJxur9TOCZWBD/NQ74xoxxzy/Vdkxp1EBPDKS4O
IhjvK0fuclHB2g9yHj4v8f92r4zyBqXsKFR/wlbjIn4Ki4AWO4Oz37o6Aaay
9fAzaaeDErh1MHzqLsmqET6rP91DKPIoTx4o5+O5l1megK8xv45IIKfu9E+u
Sl7LRlhiZg0cLUv9lPOwcRyY57Al31Fo74kYyw1jNvelPtQAGHofH8rhJXIu
P5NT+FzruuX9LnQ/yVwVCecw+/ufDtHaKPFMnod2+C/72ZlxVAP+2Mol8E3c
kOqTu3UagsuySUj52wr/4jVkUNHj6kuoJDek2pWPj6G754+Ry1umBZszac8h
0rXm5LA9KBukhnVIVbuM6BDN3SruGQNYZJm3P8gIhzcaETz9dTFCUbosbojO
UOonJSpEcjQCGtcv3DVyZs1crIunhoHvns8PnreTjHObT70Du66xPFvDX+Cm
PN3jljMf1AgTW74LpGjx1Lpmx+dUx3do7GgJzLzE8+GvZUOq6A6CnFNNi2ge
dUMcWBzsOo5Z8JMzDgaTwRqNPm89TrO+/rKVTox7VqTusGsIjKAKqQ9Ak1rR
C148+m2Xdg1UPrAdNRndCuT/xEME7syCC7peEEmywNC5vLN/qt90mre0uxzV
NEO/Psbygv+azKiyBbGmL7RMzW2vKX8PhHBzclzHI692Z6hgQdCBvzJ8j0bZ
aKKpbyEtVnEY1Ea2cwdRcZd8fN444ptAP/wx+Xn0uP30DwpY/A1Zfs4jFdzI
RfwICh7j/60J3R485ALUvEgoZxcFRihL3Ii/PJB1iR/62+mLlAlSyIYkqcia
vVynLNeOJV4/X3CoRCxg8xt0u2rHuc9TSvf7cTndNxDwPixPgpO+cPX2dY1b
EAREWtAKciryd0UpSIP9X4BClyMhIrJWDBfWHlYytlaCjGsa/17lhGBAkEMb
J4iGSJtvNqXgbyWbUVtzZxkUi3IF1WPAM2pSKIgMwYpBhOLH5nd7GxWQ6sHO
2ZnM4XS/bvnFRGaPYu2k/nyRuOmUSxy4coPmkChv7hxa/pBUo+L1Srxfeh3D
iQnpA/meDbwn2RQI8htnlUZeOHzaxJHUJ11TDsujfmyCxE9DAtz69IBEjRfX
JXNWXW/oZdH+uCaYWN3q3xB567Z7dvTqQoA7e2hZob2KBxMTet/KJKKla3zy
/boiHDb1YUNe9h9HWq2RG/7Do+7wlzByQIi2xQW+OXp2kGuTHhsWgudNfS6v
+OilTxEMvJUOhv99+CmtHIw3S+osHcgU4kABFJ4GnDjXUn+7q+kCctWwtqhM
LsiATmfEPBxtrBqi8YGil2Y8ErV51xW9MIT7+7oqb60zQ39G+A4shc+1WsxH
1P5MQLky08UWqO+dRiJhvu0T4YcEraquMM5Ked399+zXatxQw2tRFhT9wmru
ZBg6qluPGWYvziYhdfpV2JuSAKQFjC3hD7eHlj/6RmfJdNF0Gm40THSdaYwb
URcw5qfZkdLiaqG9iIPJgvI9R8HBT0CtjkOL4jIfqe/aXIlHO0iUaGOFHE3I
pjG7F/gcPAXjWmizLrIV0yHyg++1h7DO+8vCd+Bph3GxyOcjUAkxpuNQ0NCQ
CjcOYlqWcauKY1fTzeUy4SoN0h0BD9PUGmJpxXe2GzLj/pc/rJbNy/5XVJUi
VOI4BZ3tPfXDqE9Zg0IYdfoZVsA1zbVCzkKbfVKDVkvhX0OSNKn8hm/FkxqX
o2t1Q1CSJJ41RKp9abtuJkktb5WKDx+Ecmm3PeqNhRrb4lH2Zt4ZS0BVEyhU
pnlORJ9NNDCrHLct2Z3ueGl9C9b+Ib9FFCeUxKwrfV6UaENlpMZQqdeY7V+7
Tz9nf/EwsedrfN1MRPN+0rcCtrkV4VU0YGlssVmSw2Rppcy13G2xHiswkpWH
57n4PmKMdRMpCkJkT32t4est4PvqSrLULPPVcJLTT2yOABPuKgl0wy5Xc4gO
S5GCJfIipfJFuYOgZ5rGATdW4q4gGkrubxGyggpp6+hAmr8QFbli8Psk5QVa
WQ0l33drP1v4+SLP9P0yGnH6r3ejZZFEd/Q17+z83VjVHlqWEC1SYGu8CLoo
yzDrslwmBieUo2egcE/+HfBaDLXVOZSe9haVMw33XY01fNqxpE+YMcAERjhw
Rrul1j/G+sBqEY+Vk5IlMp8jO3Ls9X8gVFKJGAzeSU4O7SL6TSc/nNzvPKbt
vzj4mya5qUpoTdn6Oy+TIv0etcBzAm2x2eoRQJUJ+FGQM17vn9foL83dYH8E
1nwoBXGp9pa+WkkwOqmQZ/3FT5DpeG35hKf3PRs1pmsCOGt8U57PlWI7F2Xm
+jsgIQxii6mxT0pvGCY8uFVwCDAa/OADTz9EtHBXisXAzmCBknLJubuJ/bv3
jHai8CZcIbuAcuQ7Z0b+edSKuEIiWgJRuU7Eru3v5icofZMhwOQ/AdYPdwCC
JpyDyx0NOv73+4EplEhk8USIpWQZ+7DXZ5s5PJLLk5/0fjeSK8tqZT/unh61
Douuj2B5hyhER9FIBfg7WIq1xb4N4BRXQCCSljB6EhMfr/DS57IVeju33BmJ
jl5+AkJQcktHoi7P9i3O5ThJP/bRSGzWQZ7uKgm/MtaKvXEK3uKKd0jgVrEp
7eGzvx59Kbn1jQw4JNSstyjTdUE4dtBAMxoB9z5U5sWjrK1hxopSJg3AFsbk
f1qSTi5GL8Wce6vTaDSAOFOqMNdRwnaWFtK6mIXrgJiGU/2K90a4b18u0SS3
E5uoZikCjylBtT3b6GI4z9vlD8r9PjaQPAsZHk/SimesQM/nylP2WTCEAp/D
eajYLne/ejAreB3H0uqKj0yo2AeqlWOAho+Cfm1eKLCjrh3+KKKTe5YuQWpl
LWVeC+BUaBBMRqnTbp6EkwwRKyK/PKoniAINH6w65popAAaEEDdP1hfBAey3
/CewBKm6mUgdu2VTBHoL2p1JbJNuKXxPCEvhAhLk6ne5fL6Cy28ZXU5PpmM/
N3ZYiWHPEjYx6hec+tafcZRXF9ob2E/7HwJzqrEv5N/UgT8+sfykW6/gScYu
GkJQDbNqiIN9lLjqG4mwV3N9IEjuCTkwvtitO18/6m3Ep9s0oORj7D9FFsw6
z/BsaVqaRFY9Q2EJ/8sJ+JJVDs30CLz5nVW8wxxnKdgoWTfMdNu7CiOkpWA2
YLb5DUqPw0Ncb9ohaoGTPz9Us2sPdjFV14IBlrdcW0n25lVv6Mq7Z9WyXUg6
vzorNV7r4OSS3wqxZppApFPyYWJKdOvPBhi1KlA9nx+BUQSWsXu7/E/0Aw6U
1s2A88o6l6TdXcqLnvBhpzMhYP+55BbslK9+3wAJxH3p+xHKnV7q2+yOD8dv
xl9uipEeqLZIVuNubjWHlvmvqZgXFC46O02aG6AyZIp5V4N2LXcFa+hdQPs9
fh5w/zfyijEv7t9Q7+eSr33clefhxCvTyeh6/eL9rbd9fcQlk+KPlpLVjJHw
x6W+HF5PzFpjlsOP/8nazuW1fpocwJkFP9eSM0nlYGZJwyrfOjqktsUMQeAd
v/nhiqRsJ7STj9ZWTOecQ3Fe5SedhJZVYXyzHgYRERBlqCVK0av02XokJTsv
wVKZpgRqB7z25/QcoEo9ROX0PDEAqljBoWziWKVu477WQXyUAX7puWNWjQGG
yng7PYewE27mBeeCb1cLBJLrAb5RWfqjLNBZDmN0IcXbVrQZEPBt0rr1c8bT
iLQXgehOD02Vl0Mzr45+CDd5G7wLnBpoi8bhJaxgr81sx5zJH89wQTr2MF20
CiFXLLCnyyWOU/oMyMACzcNrEmaSSDbnG5l5Z/wSeLvSdZ1sxG1XhhoBMmF6
dDN871MiY6wB34yBsnJ6KQUaGpVHMBzB1Hl2AVMZ8b2xk00IiiOh7aEeB+Zp
5/C4Evl0ykxcuaoVHsN7ti3KlrwtDXnqS3pVFqZvadM61ucclTm82QnBoUOV
jKtTokYaGWJeTU/8iPg3m2bcSWBJ+JcUMHUR+1g28iNCD46mhLWyTATkx0WX
7rd//5RvbgUuRXB0wEhfOzRbXoBXv5r8rIPRiumyR0qn/OQIwO2TJG/tkHDc
W9Xjdfhxct+ITdlDs3h3145K+NkzWCm7CwYVgAWNDMysg0EaK09JBFBazx4+
M77bpn7cQ8Z9ZZfWolWbX+VPA+dsMwqJq45QUgT1437ccVGBywhv+qLWmdk1
O44+mblqpwK60iqqewyip/FRFaOh0dxCAZCB7bHCIz6byjlw2AETfIKnXNDF
+1/IFdgiiqX09b4NjbGWJN9yCZzJW5SIbLURlDYr7ZekAkIhdBwdywWCeulT
zLFRlvT9SUeX3q+vtNpyu+jD28ukJqczvSSPNoDtCX/CisToCaUdwPhuyXSX
pEhSUu68J9mFOKhOWezKMqpLbFKPEb/d0iT/C3Fh2kEFJ8viWgxbq5sHZhXU
UnbukXO/cd59XIsp3NsGKFbGBu1ilY4Kdjqk3Nn2+XOPKEM86TahRl2vzEQ4
atP/1KubX9z6AATvDomYqVy7iv0gMbXxhtZI5Nf9PEZgh/m+i4iSUIZgnHqE
FJYEdhAYE0OkEAn0/1uBgLCRpYZwjbenHqIh2XvItgu3Z5a3JDyOhicgDIje
S0PBN0WBtlGwvV1anusNqRrXVnN+NiGs+gsAU1T4TtqWmKLxGwz2EowptOWj
nW/6M3wnnnX6noGGkfNH+wFC/ACQ1dfnriKld8+OamBFs3paRCCYiTCK4lmQ
UnX4LmJLY/Q753Xh3nljSjNy80Wkz+jQrH1ucmkGTPnoNqs6oFZ7m72+iOqZ
3ePTzAVbbuJl+OcqjUkXx2BfOiAE73Q0V3HNA56xa9iEcW5DhVe9+Ueqmp8W
wowgVaEiEjF3zDU1403GlP/ckqKQlSSZ7vRslO0AcurKZ0OpGSyAe1E71PI1
w7vwN1ZOTKAR3JXaqDJKWoqyUN+8jh7WqBq+XmRZNKUMdcdPD4lj4nGOIf6x
O+R/vLOaLl/xAhaNvmRh9+oOfQWCUp7W6lifFsIQzwuVfK5h6I48wuMjgcdP
rMAXpjmXVLz4L/Bsn+jQGhiOw9f+hm2ZwF3JU8oabPWR/fwHyGQoNeFVAn5a
kWukAId8x94JAyrM27r7nkpBLTcs2FRg03bzfKqNon4abhEVpAN/8xwiVTZK
WkX/e9e4khSVKoHbPTG4JmlBoZ+pSILeFiuR32b5Rg2iDmMUOQQNjVY2wfe9
jBsGfbYeMBFIv45PEDbioC6zk+DdFGEvzWjhRvoQ/Ha9ZQvAguvTaF0iyRGe
h7lwxvUvUFWutJuvs+mRTu0Gq+oWvaD1OBSvMjY7g1lh5IfVcO87HFl74snV
0nLIKotuqZLppT5lUgZea1q693ffUiJvcwvJGPbKzNcqPiyJLlodTOn6YPY9
LLiX6KKlYRmSR+t0R2BDtwPHH4ebsxbu8G9OuNL6VrjYbKX/ZAzbTQKbiCO0
gGprEs5IPzaVFMVq/AjzX2BU2t7+2AO0LLroPLiMcYbl5B9oUqig/4x2wdLA
iAEpjZOKiZocEfP8GMzk00d4Ur/AbwDpZDtWczLojmFKbQgzPxzHb5OJV8nL
RoHYDIsyZU9sske7S6Ey5Nv8tnvSeeyurCkl22TzQa5J5lQoSwqjR1L/J2Fv
pc2B8tMKw5kjbM86MavQk8aX5BbMjT+IP+Ys+ZLPAnYYQz0dhGZnE9x1fqS1
434QVAvbBqt/Pm3yVltrT39mIyrT5kF/5o/JhzEQOKHbPDan0/v+mBJ/vusi
qJAW3xXcPaMgpT5Ze4OivuFta7xp2NsdgpJI1tYI9vClzzeml08Wk2SsiMAj
xLPZeL6MXOElKYpuDaj0uJARQo2XzRnqNDuueBBTRHZYf0ejBW37xmdLc5iA
1njwFuipcaq/H266dNm2+ERvrXkMjUEYH0x7AcdndRS73FMQqlPrtU6lsRPE
2443d/yeqgL6jDEeM4wP015cFmk5avTTxzsBjaWxOjKnE8j3h8Ej8/yYGcmD
TSDvQIOR4wFzETXcwUCTxTfotLc092esYweEY3F6/ACAIvPv/oeLj5unE9n+
LUMoPt8ABj9K2hglcnFvCQTr7YexUsuB7a4uZrE1fjMCVu+UD00dDTqRONq2
3YyhNFT3N4L2ArWYvjAy9YeH+FotCuk3p+c9AfXyFONQRMY5UXKnzVNeitCr
Bkbmw58PlFZiteOyPI3vhSJPckYE5LEyJ7Gd5PUZmrezDSjkGHRW+EfA9IlR
LyY7X/aIh/Q1Whhf56Xzn6kELTHg54gKEtC83gULY1a91yjg3B3gifTwqK5A
L+9M4dp51moyUUvggk4J41G/9e9WLMKtzgGLmTr9a/SR6gpaIwCUkFDS8Ucy
6RC/t+GEBt/tEPMYn05XPxXhHOWAHkaGKBmZ49dIJMpzw+tE73/j8UeHExD4
yGV2TyNf2bXEaRT9shQJ6Grg1v8b9g2EIjQV/DRlBQkZJ6JhmuR9XH58Wj3F
zUu8h5x4op0uurNNMUirOocF3w+lYyVGcPfiiha9MAqjl/JdsfaeJscpAKFK
5AzYdBJPIR5Z39UKA7aU3sMQnZKgf0oykUp880Xnmh36YdIfmbQkEjmBlCzZ
Kxz3k22ErwkwkPLsDXlXao7bLBR28tJjUu1NbuZv1Qp8OX7fQ09NFGjUwC4u
IAL7ug9vMv+NS7ltwKuvKaZuksSfnSPcOP3//eQmA6Zl2XU5I2j4Y4C0vWgC
hNS06Fy/G+53GSLvwJqlgOenKXz+6iqJUhhPtA/3Iknzd0BysL3x8FKsS/9M
s5l3oR7XyM17l0HoiYcaTnXsDqZNMAlR8sdE4QeBnKU5o5UIaxOR0fhf6RZX
Mdn75NnKE60F3OD+uRbkdsUvodgOGHehiq1s/GlVdBfUXRqFLGraxKfNbFUF
tl6G2q88NkilLO98uCLrzfMvwDGArylN+korhksH6Rb62+TRb0bdR2r82w63
ChdARoib89og861/fkgmWn15zwxUcP3FipGjaoU/wXw/YRn0x8yEUf6YHlFo
kXpcxZKaYiX2wsfLrhrOLFwH8f6Olp+pZetGcJz3zPh15JTxB4hE6kVILMHD
1z3iWr8WSYpPYWdF+0hqiR+I4pHlGhkYpJySURMouKWMsy2jSDGILK7G/9bi
jZx4li9SoVBFPYI0drMbAhrghb0kMX3nr9k63aVpNyFYFwmIpYiQRBW0Q8vt
srpiieZpBAss8F+FRuF2B7ZIlBS4pqLLCy7s0quTyfIQDe4v30X/FIPZmCbB
UCCyTFyykKi9Xa1Fow1kJeN+TVAFIuCOGlMhwCqaOPSLaIWFGN9B1mqxReSQ
1YWZzb7pxG3gMBByiguNr0k0kAJvKKxNyl1i6xW7A7osVpXEGprA73lwV7xY
csDu2g/NIb/xxJrQ1HrvmYGgkUdFDifp1kMhOYNU8ITcdM+BF28XkBDmDzY4
9UP5XW+3RPfXveiJoPLcZUtsjodwI2BQO5mmy9F4egrqcAbsLw7PRJsoc5cH
zkXlf5wlhFW8Tzu9rg/84bTG/M/p34kKaG6AgIPTM3MSN8JLL5usitFJDtt0
jRuxJKDq7q6B53qoOMh+SYHn43ZaiwAmNdlaRY71eQV5NDcYYLvKRdH3tehU
UKjLe8HGFxdRFZbcJACcAaL+wNCcAIeHMDNGXp5/Qupe9UXhWzPDT6QUsiOl
jCP4WB3uoIXUdv58Ss6IeCdrnAJQHoo96SzBCqDSy1u+LTo/gZFSXgYmfdgJ
fReEZJcf3IKb2ntGc75D27abhIV/Fk9hoAhllHPIMMbzztHuDvF6o6hq3pud
esfU0DPg0YhkQwYdDmZYOQThOeShVx3hgnjHoSY78yMhywzUYGyJxvhvBUKV
Ts8MDOFnkZE6gGtTUorbm8iYRve1dchwcCCjJ1xykMuGDkXkuAn1gHYbQHue
E4Y9XayJ71yre453AT6yBgvuveCsqp6M27RoM9Npab1ATYB0n5VBtT2FwySA
wz5ddPLrZJkfqLs4uk7S/zSALpO4NA4MFD2zROIefd6G7o8YkGU7kug8xBGl
hnglfdRmzxpSEk4bp5lk4fmJ54vIErsBHiveB82SYxYrNNdWXqlbuEDlaNKU
sGFsns0KnYulg/vi/w35yF3Q6+2uxG3gU9hhxti87age1bjMzyyIvQjNHNBs
nRHmWk8ZV/GDzQYKoFQ6/eGwBOW6xTd3otos+TIEAI8A37g75NPeaYra7qmN
hrtCBPaer975GQ67UcE9NF+ipRV5tCTQ5aHbIKJG3M9OAhC2yHgDeZiwO3E4
UdCaA5Cy863ekBHxA0aaQEyRgM/+lG80uvHJujk/5BFaJIazCWwK7V8too7t
Vd2bNNvxEOI1ROUQDYpjhBPhI2CdOIMhGqbJVNth2MPn+cMp1gJVP+mvFKbx
bxBCNHnDq8tXBN08IKLVTKAD3TbYNY/L7bGS17PTKG0h1F9lU0SQ0ApG9XdK
L0cG6xCAErSd/auEhJEesitxr5VaDWv16lrgQPcOSvj1MbPb0zMmW9a4245q
KBUsgViKFAzudxe7XUu0J3fSkgON8MlBW94R5g1q+Nuoj4wJ/RNaI/VOW5eN
imIFbPMep6IWCr1iCsL53/+VKdqcuE/LumIf4vaJU6Izt3MOQRtwqMHcQQwj
AcSZhS1CycOwoB+wWz4ma67aYKxLLtgrfGxG8Ule8MpllZy9l9DgczLccAtM
uH1HkTMZi4LKN1aw7vtDNcWASB9tAQw1udvsD+IK2tThBLKZMyXq4IJknYt/
XbyfTWKPNjvWLa60m2++KrSh0KoI/H/UY0pAF8s7K7hXMGRekhpkEc4yRTuO
/bYs6y5bw8ksVKe6avtNCHtKqfmA+TAyjpUMo6ZsfL10pvFlE0UJsmsZnIEs
0aGn+CNPInVKUbTJsvayC+MoQW9sNOUrjK6ow6zltToRa3WTq8dUJq1Y1Uz+
MGxsI9TUpcuEFM+Ayq/L01ohDWtnqizl+LA7MpfeIY/8Xo9wzjy2iExje2M5
j3fkVutzf5nmKv0RzJCNuovlt5WsvaCYTJXAQJmx4E1l/PRmH+Dcqkcqpezh
daK06z3CAMZ22wR13QxHMOr+1XnVhd4jiA3syXU48beld4FJ0N2GeB5nr+/h
3uNwEb5Ds9yLVWsdq84geWDgDh3KDWOvPqJU4bnL+lG0hANbgpWuOuxPnOzA
XQyjs0RHiKabNTJApYTg+QSBUyNqsbRken1qkBelEQSMLTQNBkzUZMkZZ5i9
Ga0KwjpuJ2k0F6Imp554ShH3NNVKKsUQrdNMfrPTh9zygMOVAIJTvMccd7HH
RbCPzzTkkzaHpHkMgCgqrEuTfjkuLh0AJvKltK7VZqfzSHea/OYM3dJ9KLE7
6ZWbghq2Xuej3tN3TPHRpFTu/NWSPOZ/MDjkYNYJgJcZWLkzHsf1+OXhv7hj
eLyv2Jc8Q07j6mSkRcbRo0sc3EM/6nnwVemvDQcsbSWZ5GQnkOBmo2iKGdWy
iny/s3AGXQRFqgnduwPBe6PJQR6G7VMKbQCZZZC+maMNRFFcBeVdM6lkMUpv
gbvAjKtsZop68WEmQG00RVr9i9cpFQDgm329z07/RCjPFnMHr9nRXc5rNuqB
o0afLaD8NMtzEZXCxJ24oU/ckkcUzkSbXViV2yMv2Y9KFXRkXSocZPelf+jE
rwka/UW3B80TcSknkV3mdB6T2U1uKNxH8s/QkIuvlnqknAcEQYTYlBfLUOYB
cncFg4SjPX1oN58esc5KZIVeKdgXlq1Yu7aRSx7EaWndceY0igriOfJKmiIc
P0sxfMPjIxMPKPLkhgjspsBaGTZBKguj+3aT40JK9QZyx0Z7YaRlQSP7IIbI
+sE+Msa1V1/u1DVJwIYQKNkW05H3+K+C2YsPDd4hnjSoXtV34NIhCiIe1vK8
OkMOwhkLwdWFe84VKijSs9LZsIKRBbdFcd/9q5BqPE4nWBRCw9apiL5DuAMX
DQJQ13E/4Z62gqanNZmwXPSlbGiz6emVyXBZr2Scz3Fo5CuUTYERdQMSpNha
T6O7BvnZMHRk7Pc0ATF4vFC3Rmmil9QVZ1vsgd4ytiGuNCgO3SliiTfN2Juh
GMMwm1bDdLlBuM2f3H76jR0HqeoM5M276AFcAiNQsD1Ch8zQ8axfyE4+reC6
vnYDKkJ3PlaRSCRn+lHumOUixbrqCg5r+4f1BbSywXDc6T8DfZaWTybrlTZl
k9TohrtdzoT5qNcxD60B2447UxHH+x7kcZ5T7AK1iqJxNmoKQdoD9n2zLR5v
0ndmwQHZhIcpjxSEP9j72mSG8JNRuDm4sJU5bh4YqgZs6y+wAR3qF+NfuKCi
EUmNSYYIUxymFehUmTIFonPODANSlZMUWU+s+JvKvchruWjLJnlCIOxyDTZE
53hVEwgaQLJbUISR/GPTlgnaZWfydFJNI+CnQRNyftZf/r0pym7oZtMCVpin
PNnH4Vd2Qii0REJzNKeFueWZEh9WELJOI5m9YTVDOwTwLPR7qa0lKbI6Wwhb
Zjp0eqm0Ow5gxexZQxTDUqiF22ei+HmP0BirYldutTlrxkboNxj0jMXKWzqX
wO2hNTrJvbeTs7bYTeX3GeeZ91oTXNJo4cs0CawQ6felPmhQEWl+nhH5vknR
2aWbWqB9JPHjP4oEaJ+z6IbkPDR//KnX0jRw0PkU2iy418rYHgJwoHpBSiPz
svNCu5H8wLYCkfL1SiLXrrvOxPlmvFS+DnA7D8gG7r5etLJ4ZDYxyGwDrwDs
m2uikfVMdvYNfZNZ63WY4UW6dHS9lXJjCrdSL6Fkd6iTI2lkuJ52bh/Qa3Dc
B3ePd0mqEpEBZApDwT2mT5dN9eOE/raL95JZo29uagRsRMeiOgfHNAZsY8Bc
5mgL5dPBatE+G8XevbSSDew907LyboYnQp+/uDozCzWLXyX/pb4sR83O1UqN
XERckqUQuE+aymH1FuMCxv1f+Qi8wujNRhXLKwyEkY54ZS+KHmWypw51Kt6j
t9yLCTu9ENW3/zc/HgnDjtR67nMUfM7BZYPIhqSDD5s12pc7f5RQRWgNexN/
yYyUO6GaD7o0edgGJu6pn+qWM9rLCLUB4FsjAlPqb8TVMN4DKQFKPebjFykD
5OEQh33+UlBVUKLRlkOwB/yrcy1rVc8H+3NSNjdVMzldgUFDZJcrULFPi0zK
9SjLprdI1YaXa/AW1jZw9hgArzLmbWRONpP90AiCyJTSrOX48QJUUrrrnE8L
wBLWJxcKyJBpeY4eR7debgVBkMw44ZhJGH5nQsJmbKxr9n3wc+n8eEer4aVS
kGtmy/bO66+DVg3JQkWTh56rQ29g7VgdBYVCrqNAZos8m88jVHHI6ubWmIFb
VMSku2FKX684bQYfv7gmZOtj2VVnUqjLF3JfsO5e0XMVxis8jDPCPJE6J+4q
NCLbdFTfgj3rQevKNgvPwRU4uLcgMZ0TMbuN+P9d+4g8UiSQr5fhyoQjs14+
d3njwKZla/d0U20fdoWikljKS+X+1cs/21sUudIe7U6AiShrJjhFYaI/wodT
dnfwXKryigtaZuACzn9r+salcy5HRYcNxo8LZDFotCHorCdfGIkX1X01i6pk
Cjzz5L+JhXlBJp/Kg2IRl58IEmv8LxSSzFgJKo/dWIIoOaJzuVhlHrSFdHzl
oe2K8rXADJX/tv57Yzewts1jK9ENAxQ533Lg3YRVQ8wwGDFgEY0BbGKmA4ez
xROpAjsCHiBM8JFdUNe3+vS7HbZJPDs3ZPJKRmR40GfXfnjO23JrHXYkgS4r
6Yt+wWo5XjO/nz0/DP/ekutNZUSadm4t0ZoG1RYx8Rp5lPnMpzp8JLKEKoi8
gydNQ9K5fndqtqUlLC6chVm/hq0McK70fE5q9Un4NuA0stgNQQ3y5JiblOze
UXv6TrI2rrkjgWNq8nlWwpUAI1Usf4baESxxGkfK7BC6eQIRfNJQWNWkHQvT
SGA4JjUcdrFfk4xoxO5tKi9+b/p0FIRZtn76J/yut7330v+RT74pyV9p+rZG
x6Ef4G5CsRhYBuovOa0kXMwQ/9Xaa7h041e/qTKTmy0HitctBjyQdw42E32N
w85N3gdb9Lw+uz3R/r1ISUDhHrFBBnjVQj1sw74/QlaeH4Wx2VZCpS85n0Pe
Ox8bbYJAlad83iJBYg2T5I+dxBZb8aU42R/pYD+ysZ5XVi6XIEUu7tyEo0tQ
dTdi2E/38cejql6cP2sJkdzOlvJaRzQkXM8EXV5pU+0N4iqvCJadbVyQN2wi
8bkWv7rOoeHhPEWte7FDzZSLPz9EbbC77yFJrmgSZnZojSgf3NG9de6IdT+1
aXy+cE5a17JWwMsgGltj/f6lFrxrcN6iXQoUUzJwaBe145fgwW9LqANiDPh9
+jok4uuEqaMTC7FHoAVhKaB48S1QDLYx+F5R6GlR6PZzNawbdXm32hWuFwva
IRYVKJmzlhYSEBrJN0s7KWT9vErRa9lrE/LbiM8H9vU0Fl4tp3yoAJBMOqze
+k+EGq9iRCN4/Cr/gOv6jIM+uAwPqPvqciB/5qw4EZvAVu2dYgSkWuoDD0wf
2oLcx04rlk6tGx8eVprYgNNVtXMxWi+ueQM/7R9HT4KlBXOt9WEuFkvX369j
NvqB4z2boL08co6S7nXBEtl5omwmOd2/wDQQuFBMBgF0guYdcVnsNeaIzdwn
3mpdQCzlXbcTzM6DAKv/Ug6PEy7ty00pDUULNms0QOOMily0k6ezxoCBf9NP
BBDDh8HLRzbr1rd/OLni8nhLhbsXh393K0vlTiKnICsu9NIMCcVW+bkzFiNk
YdEiB9ixODSsU52LbOw6pplvlwAnIxMaklpJp5lzXadZdOc41NLR1oiCP++n
0Q1Daj2jSgVppfeLPG0mHOEzWYHS7LIDv8XzSSWd9rr/+ISEMr0F0IHzlyF2
m7XPRZMlNY/wHktFtE5PQq53X35NpTOaKAncJQGsugd9ANrfZaK+dy1LEWzV
1RCcPTurz6agLJBiUU10GNW0l6Rvwhvj64TqfyL9hmwptdGRC2qsc92REr0S
15l7XpWigRsA9ZJSs4KKz9/54MTCTLtJTBnirCCgTh8pakqUP0SOV3am+hrh
VggkqBFHWZlIFhct40gsWMP8IWsvZEw/CErbldddv8X29yZDBJ2rTOMnHNHE
aasgevRlbSqQO6vyY0puQdjQnonW+MecFeLj2O9iBjM7va/f0rgCtefMU0jP
HKmmm1VRBPrIdGR8VGoaWdTTnz0uhwHuwaEXeUb3kswXFhLQFQxaIBYR4kw8
ncRTph2ODGzggzb939iJ1hbOhIwbccYwvzCWDTLH2ZyWFzJsF/GJAZl9gybn
zNddHMHkcp3B6uVGYGYIJcyeJ7fDUAUh8MmGIxH9Ah1vrNFBlcTM2anD/DhG
pf1F3AxO1o/+Yq3MTurJY236uP87Le1OeFK61cml8vT3TQFcyBkGofRvQ+vZ
d16yS0GyF5IeR5zppuWp6SfHaOf2SamTDsvD2zjIDHNOg1nCU3siStwo4WW6
tg+iGQVtEncIjDTIgGD53tsD3Jy8yzPH1kS8N9H4ZrV3DvKLrnkVRwzybQbe
EzrYv6LG3LJnMZtKCtqWBPId9NbGvixt6gLHU5eDtHpfMCSOQs/iVgPa7dfd
qBclnD2zcDaXQS0+I7icYDqyFi3jF1B2qIwLPHzhrwLBeT0+i4AR3CnjIhDM
YheXx0HGjuZLEXTDBBfN2DV6EELJQ6BbWXNIokiw79iZoilXeTKi4Lhnw4Id
u5/TJTuf5+DfnDoEiLTCDEGLKUtPUwjQiwbJMjq66C4qGIdLJkFG9VAN/3fx
cyZ80RsYNHZJR9geg/Hch6qHFSssfdzbqsPje6gxLAHpW+8ld6d5GXTMfVI4
RRAMCpSYB6QHTlpV8+/+6B7Ck0A74L6fVOIpSieMYT2svAPQ7Ct9FSROjyG7
PtCmCbz3UwBwOdZ78scbRT8GrITV+iZietrVu7T7Ka6WBvPG9jFHgo7EZJXk
7THYTZKVqki6lWuiUyOysU+K/Z3iPY4sWvgrfW4E4yFJvY9vHhMS7Jq+K/XY
TdoOU3SZSgxejctmP10kmEVx5HNDlWjmXRepLcqqhoxPQs7qQLUF8nsz+E6u
n+mJHNZB52dTudwRSe3Hvbn8HvptVgFss5Eya9CqJfetaYEM/JfrGPlE2JFK
Dq6atZTrQvQ8koNGWBA2nLLE2+xfl+5XcUVO1bw1RYWKPoSmj4ZJ0ZnD1xpj
2pp8VlmDwcbb9vEFJoDwVkSgmJz6IMzu8c3/QfqtMO0Lrb74nGvw3L6QYGJD
ITIvJ+NA6lpi/FfDfkt2iGT9rrDO78uwBHmuW6s3K+DYpJ/9h3G0rz+i169h
ezM73CaI5eIkPNPb1Efkr4edFaHcC1rwhQB+ZbS1vat8L2IL9wB58VBGVVxa
RWduDhzHitp3Mtgn8lHmAJfDXTGLpPJuF1dGRdmsZN9yTLKNE5T1LNOycE+n
tsdVZcgK9mNC2EmzzwhHnV/i7JSbNLE1ZY6L0sQO9noc5tMc8YcD95nN3pqc
eA65PQ8oEzJ0OnXzsil2c0GHdqXfDcWoZoPswAFbQjwM62Ce+iAlLDfrqhHE
iEiLSFA5PLLsgUGVRS/pkp6iwQlkQrBRHM9RTmTDcRnWhwOupg7ThbD2hSEa
Z2qyX37syxG3WnMkojsnD9nZ1o1S0D09HBhz5CQb42KS4iC52cC+UhOlIbbh
nfb9VSxTKvKMe+0R+lmKIjK4JagFLB9g/jnqr1Lqy4bWt2v8z+h8vHWXc2R7
O+/qYNgutYrbSjDCUJBZ0K+KQbRtGJ92l9gOa61rjWBMtS6awpn9MeYHq5Ee
DXXWSJKTePZEVOcO6ifbUsvpnWM97A1v0lMw4DfcnUdPLxqb0eBEWIdSoX0f
3BbijF5CUqq+L9T8rE2mP/nXXkxHr71xTl8sJY0E5Bhi7WmTvd5Ls2/Y9O/A
ynKRoOQ9SLPJ8EdPDhG7Y+kGKBL5mIvw9u/EhYC2mLGy6qXUO93ZlGf+g72g
QDKRiSiAkuWEjUlVzEf6wEb3xwbPmOII5ATUO0f/zSThqeDNOoGT5f35qdFr
qjn+P6rJYvsmIaAai1Ln1sPV8SqsOXJk7gqCjTCnkWBDQJsjUApYSDUlolZe
OJDpAg6vcWxiAja8QJI3BCGYAAT3OBCaoQx7qBlyRq7OnDfPeZtw/PEnl1wn
k9Ldy0tlOoT8KkyYiVQB7ZlDXsl+9cTdjdSdeS/nyQHH7VAw4nGjMaKBdsoW
NjFsL+51Ok6FY+o9kttojVtZum3TCDVVLQFrGNTQaI1Ccv/iwn3Hs8PwhMho
jLnw/vmnW48y3/LeHJsqYXjFoIe9q/zSXaPc0f288HUuhyXXkVHoABbaexFP
dvsUncs8OFkKdKdm2Vw8Y5vQmk8bPNFxpXQ1f4XG/eAzF6uz2oMYwp1jLMob
EjaIsCveVRxBUj2bUooR+rFfab4AmAm2enKzi/npvg3CbBgn24YaEBbpQH8E
Rfi8h9EzFeftsh50IXkHWtgKwv7QjerUraIX/MuLc4+h1KqJXSNzpuj/mwzK
iRa3BqQq5OmxwL0J9zejVIkAN8DL9vhIG3B/lez/+gfmXrNGAbeKJbhdZKWa
usxnMklQdXMd0QJVp6PTHHlbm6UzbOSeKyRIohD/RbAKPa5lVQt8TkHKUEjl
sP9rvkVU9SbG6IiIvE+IUoNX3aHMivqWBDldO6UgLwkE2FuVtuej49xCJUlT
Rs34+RaeNjVJ8zmgM+q5U3U1XdAhekfIW9vOgaj5qbD/enFqhm4TksetPckS
QvAEFGY2xhwLTwRmylZXkLNVXMNYfLfZaWt1f9+MKfhyIYCkImHsUKN62sqP
/aH/ar/3yAW3SQASL3HTIuY2RDmcgZKnmKwLwJmJoFcOW40ZO1tk+3SCjiXA
cyND3iPltAI3/HBLqCE1U6LsFKOUb2kExksbsBkv3yhBb7+GLGB4kG5YlmsC
XFP1xg4SL7EXKyMq/VymL99R8wz5Xt1cz8ZaJoc83WCMoOD3dJFTv9Kj3j6D
JaTP7vedjB7WN/seJC7ztNaikiRosMPPAvmOqu40suSUYNnB0ifHNJe7yPLh
5tMz6rrYp2sE5p/c161H2n5/ji42FqIpq/nhHgjb/pCRzKe35L4Tnn0yK2SV
mvHN/AgT9sHBDRO8r0lm/fqx1lTOu0SNAy4hCZuX8UPA4fKU9Nwvgp8F9/+q
4SNygHut03xqJLpjfAlMZeFQ5f4PdcHP2ddpkGf8XtjaLCm9dzZzAXWtSp4D
q+0f8jZxijmqrLbfMHRCRomaKPqTeu+wR1SuoEDpCs6iRJp7zAG09l06gggz
cb4oLikFaovkdmLY7iWPwNG8Evb95SQeJVJy8kZwZNbFPaoqX0rpH2eUWCrz
bUqjeq+Ua/cKc2DD/a7HZBMthotDyMZ5+Nk2+qNiHNuyLE8FMaJCmqomJABv
ZNpvUxt3guwV2kODTnRqMDIlvMc/DSTwUz8RZKczbxAPvGI4pKH+/NDbgyXC
feVQUYTHBDsAk4iWu4skrkKlf1UvQmbhwlHblMTan/WkPsabxmTNcdqJ+KNB
dSakGTMnOHvbxSuQfO/zcHvPqfFu+r/pjvAwNNmqXoEDrHBD5GayqAYgtnXk
MN6kxJlAyKwscOgOqewdLx5WGf3zRW/E4NlggMe2bBp8qm74U020AuctUdGd
AupIcTYmrgG2+2xQ5hykcEOD1JegoHfSuRktdO7TK/H9TuoOvGpdLrgKPfcb
cOznxWe5ZVnOVdBvn6UHxb9i4tS+AABfGEwU3d8vdP/tQ1SeuFYVCGUABN7T
ctRxE5fUnUzudxRdsvms8jjxRttiPqdbvW2Z0GgLW78cne5wa0+yYu4+GSeB
ikP60bIKC8nomUJs0Cwib7HTzeSK3dRJyPluinBzUWisXwAybVnROa6SWZ+e
m0Punbj3nDZKHIFpfsOvYX5mw3Or/TcZhzl6DYUq7qHHWpqPO1f0VJtQWAZC
nKDcZWlJ4SR0Aod5bdgIVNr/LAd7TKbNEf/Ol7Xy/Bapc27Unv3pi3Lso8P5
imyvykQyoCDJb9ELs3WXLbvg9+kX9d0gzFkrX6VzeApEIWxNBqZHF6zHRQxS
QEEYabwO0QAN9YDUgZKFaY4YAio96OZwk1BlJvRElPRDRzLgkiKOlzrUYQxZ
O10dSlt26FWTecaPUuDxBwGDwm5Fc6mfd/UX1ykYj6O6cdaxpdG7AKlUdQAL
1t9PYz+HIA/mkgZKOSUvaDw5+3dO8prK8EPzyL9lcgABPEevEnppTi0DvpRc
1QqJJM7LV4CM8gn2MxdDCW/llTJgfeGvTkulepQWvKgiZ3JKQiIY7EsS+Six
+ioDKnI3pBbI4KGARiTjka16rFEv+yDBudni2zb9hSvMvhWwHN/tFilLRhho
uKXWLlCUxYXwXh+6ov/t8IeIL/fv+oUoXrfIXZzsXHujbqvBmHQdy9MqF38r
PsDXXpHIFo95eMNMr4AQErS7hipcM5zla/OcqMi36mATWGauPp+HzEnyevc0
Qk/KkREcHVguj5/JG1JYgbRiHi+8ZlSP/yvcQXUwBbqmjU+Zh5duOCtAl+GA
OJdyQeHXGeqQYO12riqsh6fAruaxUC134fGIzyz/ns0ZiDfpzyfBdqO1iqCB
ZxN0Ri8o7Dza38y5KHrQdp6KqtRZWB73POK7mIzDhb10Sb2FCWLCHcDMiXD2
vAfWSo22fg7NMBPN1hZRW0suhV3jwGWBmD1jC4pFLqhuxbOHwcWPNlhZeoSK
Jnuz9mdb0sh2Np7UOzksXp/4lhsJBaMijtyhg74+JwUyS+aaSIyPFna3FqBs
8JE/GCnR9ffqg8vpj3UxTiUmdgP2Duwi/aj+xAMe2iX7rOaGdNdkdXkILZdu
RjJg9pLhCjAePMPHW3xxvl/R1jXpYU1I2IsijPvZsTolXH7Y/0DAtvvrG8YP
1UOdFOJBQd6eSc8eh5bJ4EveZ+n9zujhONdXqQ463o4d145yqQuUfvUb0vRz
RPTvasMWsj99BEyVWsrB4gjmneZfc1Q9mP0TtTM+YpyxOYr+oVPCVPkDlFzI
z3uU2qLgFqFXRvr3AezHBPDCm66JLNwI9oz22fboZ7ZFzqaAB0OkW2meuiGV
XognPul+2/yAxY7etG6G9CMjxJUjeW1k5sPNfMpm4ND5KkGzwmuSHjxqAvX+
A9LptPwYidlLQ9GcGYL9CD5hMBv67RzsBP5XCjy+AmGuBdfqPLHHfq6iwLSn
XLV8onqsPT7IWiIKmRlOsddQbdh+jwtowZBoIKIkpfsnkCuqX5m28bZr1PVR
oCySjnHGf309LyItdCD463ALD3VsEGmewvLQPcy1tEhzKK2V6FKj2OjFGp7t
ovFrOYTtAWx+APfhN/qmtaWVnVxMjKXMfUbQhPLTxtSJ/t2YS26t0dDhQ2hX
5jD9MHsmlQvJXSJy0yvo4HzDdObD8aINjLIQzEaND4IObyspmVj/7btjBj1l
inIZP6tjGJ+TPIZdIu6wsgtHkYA/3esU0PKu+8XuSEEOwliHInOmm6D/mV5W
eJcXyoOcxT/hUFa8IMrj+6aKVzbF+8BjJWh1O5tOl6cgv66ndWNgubsoHcFn
mlHnvg1DLGB/VAG8EKvgIeVyh2bC/40UO/zEKDz1L+r4KlzPqesg9HqMwqsq
rTq0pclusgnX7DeuKHpThDNOCHSUdQDu5x91z/6xuJJ4b/X5thzLekwVMt0r
yUFlWm1/w26to3zwQRFmVHuH6V7YkxovvOh3Aru4Zu7af3LrzOA09Tkql30B
rF2PhnbgRu+x7sfFZqlLiDohQZT1hw7pQYHeqw0IoU+hOCt8WcE3xqKOSPaK
eQthXlYMZxLPBeRCE03yrh6n6BSNFo7rQr90244e3d6T18c4ua4Ct8s+gogK
dwKi4wLguxPJaoMNKjaOqaig4U/W4xKZak3iAGznFxStq65aSEwQ4EUxtzP7
sexqlLu7ctxfNt/WL3X9VUXwoX2At4IQhhDbJuv9OnpT0f9AzzvYBNdS7seH
bEleeuC3V3zvmify6pNqWHB3P8ZvJByXj2vZfGh0Smha3vfnA43uE6iKwpzY
BRT37zkGN4A7xrXIixlOhRCck2lGth7fruVGdmcomcWn9UPYg0ceQwqwoLwC
3yhpytaF3SlN05hdoNgESY8pjdpDbnOQq24zl/oBHHDYioPsl4SA1x0p3gn6
5imtlmdsPd6ith3O2/Kny52qvcuaQynAWfIXwKjy0lJchoirMmeijnz1Tv2u
LWz29ynAsE3Eur8/pTw/VKD1zp/JNlaM9pVk+u1xR+JJd3SiECRHXd1u3Rok
u/3ct0QTKNj41TSLhAZeDM3iYzOMxuK0U7TL3u11djM39SMzbOSc2zgkzuVk
Sqz3ubc9Zf43DPoES3OsTM0+UBx0446mdhNJcg8N/C0/JK2Jhr3VtGpTiRwo
1M17AJHq9s0D82PbZn5FayG0Wvu5dBC8Iez3wVJvE8cE+qilp11iSsGKwrAz
yAGdapM9/sN8fk7n8f4RIXWKzmdlAOF0I/VbBoumD+n7YrGoENoxc1rfaV+K
LRDe0FgSzTRALhduMPHubmN7yWnjbNmYg/q+0t5S7VWFH2khx6Xc2eAjbBb8
dITPHzRa9+KjgTnrROlbKIrfPhwzNVI0tp6ACxYLXy2JilVNqBg0pYs5vWx2
Vb8zt/sYGjG9R1TBL5eJvbKIXvT68k/65E415y7HcfnxUYA4PZjDYm/X9AHP
9aMecaqan+UnEnI/tPnWadr05in+VUVUgMhDrFELzG690H5az1LxtMhgpOw4
Uy9MzKrzXRNwqtiHerW9lPifaM5dC9CkCjBqB6fyB2TLiYXQ6K4d7w7twG3D
yp7UDBEZr7r+2wFZm8bLvB4MYcjU2pv4MR5Qw1hrf4bRk5jl+BbD2xAPGRQl
Yevo4cH9T4jA5FZmzDUjc37hQWvf7zNvIFNnbA0KRK26WQ8gKA5aOySIDMTZ
9yAII7gYn5fU8QF0ZdQzgkBKrnfhtOxyFIG9wNkfVBtR4apgpgq25IycR80b
xMdF9qma+iDE92qR7KWRi01pQSlnkvwmaDriDwyrK8ibXhXcEVmGFFLte8Sd
XHNWHlQEZAeDiD/n3daH/VzOqScAfVGGQKZJSaIca2/SGA3eewv6vWCuuYXn
tJvcax/cXn/ANa0eMVrSONsXXFsHddMjItUPFyVEeYhHKfOnS1bLI8fIVipW
+1jHVdRceNjgwCa0ehlz1N5mUi175kwsyjAv8CAmooftRqMM1Lx1COVQlTqm
WjAIivV9rfTBifTJcSrLVRB6EKv8jyNw25M6k9Hwg1OYrHmR5Y7VCQtljL8r
eyfe//0Zi3XUo5Kye4KAzpxPqE9C/0uYtsdIuXWPua/qHcJ+xOgKrnAFh3TG
+uL2WZ16seq+hn4v8xwCMUKdBmpM6VCfEM4ldUN6PXd970ESXUu+MTT8iGGj
32kwo0Enaqd34l9fOEeWopj7AZeHlymF0DIZlCpg2YSiv+ert3nQeqCdDDgx
03LFVPO4QoTBTj/frYmGIk3HbPJ7Fow5ZNzGYB7lG+OU9Sg1i9ZivAsnFEU/
OUF5IOGvD2oEDbiTlrkuhOKXf5g83Pd9/C5YjL1UEPf8wtTKmhKyTjE991r5
6I4IQSEOB1X3B8sD/3rzjF+m8P6GBfTSqnTWelgVydaKFdylXOvp5Z2cRYIk
xD9u4WQkb/b/PNmR/FoO0whSHs79wVY7mZYwLVdONSwsZowbn72BsuusL8jw
jgOYqzRUEE6LC2FO9+LG5LDTt2rQyohnOKC9AImb68ApfJK/tMMKBFnWTcsx
KELcbrc6HngmyMTwiyJqY4kjvNbj4knD4Sq9dRhbD4fX8Z0MgT/Bh0eKynzB
blQlXOhhVfMNA8CmzRhzW6k1okyCKOzogbCmK6qMiVGle8q52Sb3+J6d2r59
1nYHDYeHM+0sNbhm7owK+An5pZ8yiOmFY9+v1jWKDtUp/aKOmhbWJX8pOfUx
yiwbyyyA97x+3YugAePVr00/ztrxGPCzqvWmyf6DD/FaofhcBulvwTZANPLG
vB+zFxOq7C3pIb3lHDf6+79kmMfWUonBWEAdChv20WRluYUl1yGUzKKjdvJJ
TuK7OVR//EssgwITr08uKncD86YXJGc9hahSrv0yzWmFQV2hT4BZGmICPurF
ZX4tAx7UGxq6oSjof1UR9UYYbQPpaRtxPQmpc67d7gTZJSCB7fpsBu5pCaDe
lL1V6f+zUAHG53tfi4xXcofhvobO2ksJzeA8/7HfgugDpPKFIbxVmYeCu+l+
vbEq8NptlMtmfmfgbW9nno1E4eGHuGhiabMynzzCTDDl8ZEGQiWVwQPy2r+m
H9cT44j+uQOAGpByG0AgtUTW6ZdivqW2OoznYG3JmBW01NVZv+dJZ6KiI2Gd
YpBHs2zWulDkJr18mGT8RQ6vt9YjPXdiLsycsMvt3SsuWaNWS+/GWlJxXlgi
DArMKzAeHz5gw9f+znm042YcGSCiI5PTZh1t4qMcyWMwDZpObo2cAMefj5kE
FrdmyOkRCUWPTEXO3fkW7YXBapArTnQc+2CcSV/jOJkRgCdmu3Ezv+ABLBo0
jb517nqOwS91Roj0ppH3zwWKlR1F1oRip6pskKh9wxgZ1e/p18o0xK3jTJ31
DOlSmrXqjA7Ld1aLMNJepszL431fj//v2L4tDJpXMFVPPbrLaurFUXHwTrde
ch8lN2BXSwFyEG9QR4FC8YiIXGWPTSHIGIbZTFTg8xmpuM1gb6gwgEwp4W+d
lgsQR0RYu1C3D3J9tm3ncfy5lp04UHoQc0CFbxCbudjRG3wHvmD9uXNbivMz
6GspYbp5UisV05XLUzBv6txBGmbURDxR5O5ctYOv1S9NcCMACRGy3VHYRLmH
oTpwElhiS4QY00P3umdYeVx89LCUE88N/DgNroflRpmDeLFvjF5dmXc+yu1t
V+nf6eymXmHr5kPgwNRBQrFvHg8JgmpJi4vIWTXstafibjjcZC0F/2SehdGA
Rb4NfvSGEd4X3a4Sa2/hXJURCOqSTM/6D76mwkhf5fsRBXm34hJMmmp+RzE2
y1rBUq6uC/QChNlOZfSduA6WzxqTzz1uMYAflLpqbY1d3RyBfgGMjdoUHGb1
10NWRrkrcA8IUcw6x3E3yw/6EXhO+KjbN7Riw/1aDzqZAOnnYXI8MA0Y13Zb
gOMDEfdLoYmdDXIqxporlWTireVADHJ88p4mCoMK1nklnwnGX+Y6bALmHtg9
KhTPKsMLNKG34lLsSO3nGeI5YDDgQQ0K9apKTM0ktgiSB7BKfeuaUXSgpSi2
8PimvxnVa30103qXIVz7jB0BBEWhxoK4f7M4pneKiPrX072IKrBBWA9n1QYV
lF0X14MOKQb1DXUgZcjtnVztr86yVWRy808vK4Zfj2swZ7kUlRJ1CnjM9LXt
uBAVIUa0gkY1MgKKX7a20zl6wRyb14uggybSffGmuTg52z3pmygNWM9UDN0W
IA+RNA1Zxn6g0qwscZWUaVjtws2I5rjDBfiwn3QbvWUMqOjiJhgbiPgycIdj
OfQLc2k1yP23McraQmNZ9hMSxF6sbcteikgrlykTqITN+2cLyUJCECLM4e7r
miv5gwyXxAyCPbHDEg+ZS4WrNqTgXLhKHXN8iBOl+WbxZN78Y0Sw5D1xWKwi
6qv3TK5nhYT6v85LVi3J8qStE7Rjn0tQprkYofWxiOQgh/gCByvgqZuOM6at
FOs8t32fKeEGLp4XHbn4PEp8KrPZu0J6wE+v9NbpDFpLMfrLxjdaJYv2IS43
lRIANMqm852GibFV0DVXQ5H1sd/Wf+B8rrg8Pg8iuZJzdYN9jZDYfXyfIas/
28/qEkH4cUV0gON6k/vPnBxLrrdIDal9Tj7m8+2mvRrh6CRZ7BRDBv0gfp6A
ym+X1JsZCYm8ZmbVDWh04sLchS8sSXP6mrFYJgzeGdSk4y6R28sAGRMP5PBO
IxTjAzHjncABSImRMPdpd6cSBtuutsqBi1P9DYHJtyvEdqlZFaVvDcU3hwRB
FR3d71ZNgbvD+vNpgZ9iuBXBtFdzgyXq8EowzP6VYvlY6vHCd22ch8xBeQX0
WrGe8H0WPuQjBC74CP3pEzCip/jpIc0iJQMaDCsio90cErFy4iNKPPgAAi+y
lIQdzxYHwhQXJ0anoSAgupGsv4Y6xnthrA8+tTlS9iCaDKLBngBg6wHi+t9d
MLzzw2/zjtqC+UEsGSlAzoZ4w/j5q+ugq2hhJc3ohTLUiHdlUT+EKiID9JMu
3nCBDzErjcFjSyyUuJ1VrAJNfsrkJh+dGAFDTknl9oA5Kr+I90YrkiXH5ZoO
Rpxv04tB7lW06hnC6Fbro14vprU8zYGmWYl8j6tiQBxK6fmKCLqkFIVF0qiL
RuJnTGTnluaAHfmfSG1PnRqd53NBMirYAWSfe4qnYjvFIJLnzuQgWGN/c9UK
gCSVm137eSVlS0Og2v4/twqN1xD8hAm9xOy7M6NFLKrkgyzT6xb+bQ7sn6c5
fEp+jK/JBJ2DsULw2U6rYYXbRYcxlumuv32mCuerd5PW+vpYHHyRGxXgXsDt
ZBSw36qTEyDVQbA8dZvw9G7YgdMCBnWWQVY59/fjna4+5s0nn3BEGFUiYsxN
ld1o5p4yJC4ZcUzWEK6QChAdZ5AtP9nfOrrBWd8nlzI23LzZrSxxq0/UMfLg
AAbB9/11x+bzs+azgjsFmk/WIGwZM+7x2UVmz6WnQULm8yHJ+4kH+Yb1WwSh
mnREe1D20NUQHOl8y9fZqsW7jzrOKd7bFYVL9EHt8odlWOWjsO437TBOf6HI
KcFyj5/gwQz3uVhC1sOezHqFlZ8Y8bM02OGOBJ4cSam+nnRnesQ6Oiu27PWL
wYLq/yzGacwPQOWJQmrtwEQohjk+wFBFozKqJdZBT/zcO0rn1drf+mJvJIRw
T1B0bTj1frHZkzWeNLGxY03B/kjONrfpQAlgMqKTgrFY+A6UmFtEElHJYAZr
hIXOW4+uRRpRihr8lXhBVPrM35Jhogie9uYuET9r2tZAaRiEfgq0lIxPpyx8
NcAuyN72b9HP8wSphzWq23E2BANqXAyffSrU5iS2xY/vslbA67SvPLJkqnCL
HNkXuLAnxnElp4puAoDhMPFxzcLZlxKHhp4zNT3btT/5R91/+zPsFapHoS5X
wuWh7NIJcjK8UHFkU31Lbze7/LLVdKVaT/FTKntJMvLZQ5g+Dvt1MKEiReta
HMLYiMkASOjhTz9zaFebnhrHmnk/PIUNe8tFXJ/ymU8cyHkFIXEIKrVJw/tp
yWqvomG3UEPWdC1vwhyeiqIAaPovoWC61c1VAuKhJpwpbSAkxX1yd5IwjSMX
QGNGW6IS/mKrMW4COVrQ3XvZKHws/gblf8ry3gETY69ACo42/EJ3hByIeGug
QT/JoXafmGS1/3/oVW3gw5zTs1oupYq+/5YxHiTWw2Xpl5KmoOanUPnWNMHy
PJdRvVzSueAgBlEvV3slVHSunsQ1G1PVvTTjltqWMpgPu0U2uAQBnw1uZGoH
nJwv/dYsnFvCjX9OC+wd7NiN9Uk81RGJPWEOO6Dqnp61/qS34wxKXUd8gKeV
y9ISFrwp42S8IIb3aLWwmluNU3XdpdbbxY6QxpAXaZcGo67DiUIkWxpG46CM
+ZL80vqkQPiyIl9MHMpKmj3igD+V0lqwfj7kxecW//FUgwIMUpp/pITPYisl
1CQu2k9+ax+fDGOYW/9iTHi9y3NrB8gaXk8ly0mXXFK91XAACSCSK+L8KRGr
lgcTYaApr35LStQN1shcve0eEmthBVl5Fqlt24WMB9lkF6X0cHMpFec5uagm
FGuKxdh5S8BiXh2/hmWXFhtcZRiS+RcUUCsAENKRwUsnF00oe/LZRXdQ9SkR
kdmaFVNqU3ZpddNb04ThVzII8pavU+drOBc4bzh5mY3/sKjgts93HHB8nTxq
3NjLJVV6JaAMcZdTREjg5iYKsPzNr9Uilrv2h1yqzU+svNDvIHdUtibPIhmR
C/k3pYgjU0rmD0t5DOunWAQp5qf/IhCLVx0zZixdImCXSx8l86hpe65PopGW
ikEGD++jLJ0PbZdsIFtp/aZljX09nOlg3KvOvr2PS01s5eLufug/NuwxrkRk
litDyZwbwoC5zoHExHxJVdlcE2KV3vJRQcYjY2BpFhf4FAvNRXur/TBBe+UU
mmuJT79aM+xWMgOxBouSoyxaHtt9CHmmXVw/vfd24wLbroA8JHgNfY084bfj
6YcD2DRz0UVwOrXOozP8eEty4wk7h2ykpkhzbWQhbB0coT8SXY+4w9sI4SvJ
a/m8w3tNCzy+b8XCb8M0mRZkNtxaFEBoM4E8WPHCLyqbm7g23HXq+kvrvMhY
xAkNWNf9jhqFuTL9nIoT69NfpnlGaWAb3iL8d/IqQAJuqGUCb27Dvan8lUGs
8m11oifn6jFO2cYAkkmQBdc4wsoAwm5K+gsj4bz9P+FwpWx8B9aMbNymFQH3
f9Tq0A8G0paMOE9XA60zNRl3oEtaMHWbc02sktjrmrvSd+BGuEW5e+m4LJss
6g17ycvPtsasWNMVo91xqajmnzNPVKjHIiI0QoszSP2eY7kImvoN08Y0DqYz
nCJ+MVrX0sf0AMwcuFMmQk+E6zLX1oWjvxrsO1R7oNrHyZkgOLdHuIrEqVCr
1QfNavDpKy96s8ZSTW8B0QmpVCOemZtwWuBYpUafByuUB35IbnZlktLgx37A
Jbo3KisVybPGvQGbbWWObnn3x2LCs5SsenNGKKzN8Gti3oTBFP9mOdE/6eiz
ZA+xPBEkgZxwmHL6u4nksDxbVIPjnV0qrbWls6sb2Yj189It0FTrbSgZIgSm
8fR2PIwCq5SaSoUmV5eTum3PR9wqyiRHikYPpBGh1eScGioHgcTo2WnH1hP1
UpghOImQISUJf1pUmyfwgZRfYqzxEf/jGkqmHBj6lNfuN1NsTFm+sPqUsa+r
rBGC0NTgXAPdGsg2KRzQ8dsRoF1QquNFAjtEWqH26AGkQjTwhLT9LV20RX2G
wxJJ9hNxP6n8VFq5caaMZlEfW66uio6uam4HX7UKFVhSrgshDEKUyBOOt5Qw
X5XS1SKitIn8mtuVONiQvfSj+NZFBgBTwHliFdeYngy9ZTxlpJDkobKu/Mgf
lfMnB2amzI9TaBQvNQ31w6fJ0FT4UWUXuKCpQD7d6/Q6525rHbQXB11UoHrU
yJchKYPBoeFME8mJ/Aqxx6RnLRPQzMI9gys1+9dYYg2TgUQaJTWH/sbkm6tl
c8bqnq2k3E8yBQ3arwaDhi4Wf2pe/t5XoLsV7xJjESOeW5oOnr2T9cb+QqFc
Q/y1O2Y8o+gIuAyW0WgVv+sP5hrMxDP6WJsa/Czvp+HcYFrTXW9Dp/tljrU1
cqDnwW9E9QC4fQRWJM26a/GHaVcXeDLvyiuJULwvQ8I5r94BywmEEO4AzxPO
48tC/TaZ5ydOHBYbsn7yOaZxa66ji36zsO8RoPJzLyzcJqSTUAD36YnPcBx8
rbfd+e2l+vOJqXADpeO+I7BICvc4ArDgqhKBDWH4tCOgbKIFFS9P/9LhlDaW
gY0nfulqEO7yrPdRf/9udCzvz0vitd/E6P2v6nyiYyrtNEhWaqo38aLrwSjs
jAnzeQT/qmhZPiLSpDjHEHjCN4y5T1zb/de33XRI/BLFWKdFvUr2uWQr9CdR
V5D5ZFo6tMMUgSyra5nbgudVsQ7CCwoBb5ncVaSGSYyvyEvYCp5UocJYeOmR
Gi+tu5/Bor78edU16FdZqaw+ow2xKCi4ukzkhG5ihNaHz786Zwzwkb+95KkQ
1l62LiRA8CVhWXoB4nzL7x4pyTI+keXAXhbO3VVsWgXbjzbFh1cOMdwTey2V
6KpDaD1wWLLPXdE7i+jPySiiely3x+0+mHdvQubeidRkzHg5uv/GgQatwllw
fHQfTLPp4X2JSQ2kouxXnIS/fGr/l8UmGvQzHMekgv6MnLquHtpCkEQjmAFT
Wiv6XWx7rOTnzC2r4XluYB7bN2ZGIjmltsrnIjIFB1P9AvFh744A7Oz7oSnN
h8MksVtQrYM4ejPD14bYy5sxZcP/NlDXFbuEvRJIKhrnbOV9bhQfhuddsSOh
f/zL0pn4RuAxAOf0yQlWdZe4w0PLrt6TjRE9NlMkzZG0F95vjfI6740hBFAJ
khkh8elBAUQoxmeVfKxn+xv44Jp8L3wdxQv7WN/6v0oyU8zj+5QvqcvTpo9A
RsY/1pclc3dIPdisYdXj0S51Mqo2VoxBBo2By+sGpac6Z9ZzJCy0YT4oojEK
Ym098iGI36lU11F0YrUbdatTYdZsFhJCtMmQaeXdTXyv4iunADjzzNYlV3Vl
Xqxo3uvs5R6laGuVfEuLYTyGhS59kAzQzYZrADpumsmwJZxhBpevtKVxi0uX
EIY8EV8MtCJ3RsJGeBYQ5x1Wn9mcMr0iVSNrIe2nLL8R35K4VMHnA/NyW60a
0OtZMTPswO0fcems8DzQa4FkoIMAsmDXiCnZx0mxfiyUChyZHutNA/eWeG4X
Y42jfzYXZBnLfssUbQR59snRxOCheo5gQk6T0BxOh9LRgZ2UdnjCjy9nUX8x
qkCGKdti6+QQL4quqkHlWS0Z1diGUXMjwfyq6iwnUrrpiV4E/ob880GoxmMD
I3ndGOvqRJcnod78KxaTl7EDwfUWtaABW7tR/17jx0ZdFAsRy5e3uxgqM17y
qdndeKMB21YZcxY2nmwsNFFudoA4CmrKovQIAMP1/wOL5wosAvD3bz3+ledC
SN59az6Bqt4hnCejmeeOCQru1336ypE1WfiOhRtjPJjBGDYV+9M9z/wnA2Zd
IsDqVT0cDF4NPtI+dP8aZuPoRAqlcqiSyPE9dNE6PxGjytyq1/KAxj8+poJ0
+4tkK/Vi+noSK3bnx5FoFKUx4ZqJeyIVShNwCppjc2Clz1+2NTZenjsY8jJC
EwkJAP1GfOh1QcNoxb31xPMa3x9k4rfJ6EzFU4lauqo+u0CVN86/JZrGGHQU
sxLhv8OCey+NJMJOuthZtym0QpJV+qrW5LhL1Kx6N+o39anSYscma97orNly
kkI4/y69O++WXeeOKaXhLf+gp6JzFx8GQpzpX9E65MZbBoIJg9IbJvH2UWtt
ibakWqiphZ0g2VFlhJnqahQC93rTUxayqI5g3HhqW4FTS1YmfWMKMSkhp/zl
OHYts/CgalZ9ykcA57RsffuXdfvhwUTuuCpowqaXmf/5RLqdC1UhF1FtSxo7
GIhdV37EHY5qYVoMYaDQ1a+jhNw3boPl7e0n9eXrDsEn5kT8IP12Sh+fe+pD
OSXzr5fSDhrYU7h+vvEloG6nzGdlfL8cHYjOyAwAj7uRxfKNGnSCY1KOShuV
pNjyB1f9lCq82nwPfs/pSwqak6OK/+WgEt5hgwwj2oq+C2Pm1Nms6S+5ldzE
3renl+KQPtfsTrZ+yh+ZpLNzOcyLli1pHBu+dlivTR2yUV73RINAjX4zxKxs
weGCth3MSfUzxm7xnxyeTP89JXdsbZLcW3XtgAYWDUsA5lLpB7GIoNzCVyf6
3i8gOkq7Iwyk4LHfVFRw+AJizsGC6LYENLoTXMhqvhVIUOBJw/6TBWJBa/UY
j1iQ+kNPbnV0SDaNYG/Ecr4YMZo6yjsDlCb2AzETWDzLUZLjkv9QsDXGVCml
Rd6Vozcr3xEK0Y1MdV8qFZeNF8zD7vWk8YWYCqrYEtMMtiSAvOHjD29vK+xW
7iOeg1mblmIdxxL4CC3g8WUC9B79udvJ4gz96GV/NHa5iLg4jf2LmyGH5br4
Wdc4xrt+z/iKlukIwLtpRhFnjWN6vm6te4ga0AaP6vJVXlGk0mXDV1gx6/Nr
b0PsDxZglh7bZxdwLRKUQGK3vCdr91ysD2f1tV7goi9JHT2aSoXQh6epG5kt
NmHY2wYj/MBIZRY7YFa53Sq+cBywDYHrn0nyzDDss5XEsI5A71yIMRXE4zTj
URAFkZkXMQDiV9eAMa/VEkT6UC5UkjhcZs27ODORyOlfZT/GbCYx6bQnPYpM
jr/tfTlHqBZEENSG9vDzOgpBMhlHqhFC/zXCSKd3/E+O0Zu27twFNHgq6Pxd
C2ekbra6MN7MCQ1fNZvbfnmFctYmMPTOy3gRalVtyBZIuoixcL8qpxUAn2O5
qZE1xVfhCckeVnWakON5XFyrAwxQ7g96gxDYtJRgujHYVYctPi/rtDKX/umt
km64Ma6kHpjXP/JL4nPOYopXIWLQAmkQY0RdJHfGoK3TIynoQPGIh71VrY4c
R8qg2JMxCQDwA/EZCyGSxnV4K4taJMordw3DTqER3Ce0h7n6xK3vNeJoY8/T
/ubiNwC+WhcIbUYf8LKhkE5AfxN9rxufRIA65DRysUicjr8P38Qc3tkHcYRt
CLZ8YLeP71ESEd8YqJNkMxO5rUlhMp36Mswjr/Rn6kOHm7IpuF7djfoxTNXw
rMSfvpuXWdjJ5JLGobbv3BDk43fYTx8Qyw7NfFWLI4rTAop4QyL1ni/mLAUR
sjXD+xvEvU//2aXk2q3vyUQFqdGxhLNvJiA0gOuDZxX8EKj2EvlB17K+eyDx
vyhZNWy93tdbYitu1C+IC/lTGKpJMwBC/GEjYyFt9uZZE3i1iwIMhTahJPlo
u+gg/wp8aKrv/Ial9vRutcQS1LyN0J8UVt5NNvATDCrVSVMo1ViOoCsHHEW2
pSIk5sHqHkmbUOjdUamHqx25VFpEy3AgT7mS36KL4wmdMhQS7zovUmQtpCYk
Bw67MIbpE7wdG8I7E3zx/dgD3EpWmDc3rsme3gPy8/OZ3mhD85chDKSSnK4T
47gmFhCIiSSsqgtDjOxnIVtDx0khQ8oWanOTFfWfE50mN/bPaX0DYLX4dhTM
ciu6CHoUZY65t72YWKS6q7k8vbLt+4pVB2KQCkB6DJegfLX14uhu+9NosiQA
tGko8OhREhRLptwBegnzIdZgEF7ial8/yXc0jwWWFI4qzRAvkYK6epnL5tTG
zyhNcJP78LQJxN7Prj44HXeM/v6tlMI8uQI6169no/nz4EKj4m73X5p3HkRE
3x2x1KktJcxWL9sIzZR5FF0fPTY/1vvgccUTwTsx7Zda9SEAaxeBer+onm0U
u04pVzS9o9+cRdl2qhVn5aCX+gsYr05JzylWQ9je+xb/+YxLSG9Js7AgPS98
J6zi0nqOopubfA/qDdHp4zhiO7qVAwAKehMjGGraE22HL7n9OXOBjZySOTVJ
M8fGCyrHAnjw+XOTjl4KjB7pH13LSEjlgblDWY3fNF+4sLpsl2pi3imsXVlv
oTXsz0C4wFUUsRjO248oMeU3AF/kDNh6iaSYQ5gKZgkHWaZDLxnExKEs5Xkg
0/N5GSpbThzG3LFrSiKhuJKHunOMIFSELKosDea3jH/vF4E+EjT0+DG8xJY+
XPEDC17lFBcGYvdZT3XllDh+RcefU4Gah49jY5mgXB59nfHGz/Z/OHp33w7E
uN0bnEkMop1l1A6iqZyrdMRjkJieQrLI/xbVy1P/N+J+6M0jqlJgCcb39KnV
pUOWOL1YVzQf6aZiWVZHtujkDu+GW50yglopANeLJCIG1d99A0LkjPbGjo1B
yvHgdmg4YERyVOEuIbLxG7yw6r5wEUSqN2+N6yvhsuiEkZrXDSKIrvOmNujU
VXsoxPYqL5k64i8f+B35XfUEuDd0vyXpCMHfrSpi9hsVozsBTExzYa253SFA
WnBHB7VMTIJQayYzYjl801ABypkLp4ze9cwKD4J8GwZ3nKOJ26qy8DBeXMXh
o8svYu341jhUiG4ffL19Ot75c3wahtj0qp9+YGFSptEBF3/yhNjgqflauMCo
RxXvFxaUqCcYSzxwz15N3sh0qvHdOGFhrB+lOjInKAYLmaG6r+AXJRQySv1j
2JxRyMoctD2T97CgAwnIB6/SHOypLS60GPG3NVvaj/bfrOWmcGbqjVTXVjZ4
DFsLFLG90Er+xyT96E1dyaQe0gGJgHs78qjihac94DCSr4wdGOpHb1tADsGg
FpD2cU0zlVXElyPz3gh/ngalQeLHGAkvqgkeNXMMhigNa1cJOiAacDan9gZQ
SGz6GwaInMECi0WjgtS9W0nV2mVDEdSb1fVHVtme84rWisb0OLlUHUbhg11p
hpzBV01IVoW7z3SNRoHySuF5pgTCVQICJefeIHEG2hs5IkqIxlJ5U8aETSyo
hs4SH+EZE4RqM2fF72PDlFuvDZOELn7/yCUvSKtZwKLijchHhFrsMxMLIFf6
FSd0lFdGzp2tTfHtEb4uoX+ueDcdTly5ADQcIWWQzqGlgJ9UNHTL98X/rNL+
Y5fWxwp5JGr7Q5h7Thqey68kuLX39MNcQ7J4k/nE75I0/KUkULa6N5hHpEsu
YpDeXxIQMJnzKVB5cHTDDdxBKwVy79N8dMUQ3KeIS6yoE0jxidsiK2Cp9FWa
tcF8dR/ZydL8SeKXOF8oBWENieAVlH61DWFWzdJYyqDda7yY8DwJYcm7kVr9
Va9MCYYVILYDfzhjMVfYnvTOI0qO0oahbir/TKMcPolWleOycy4ElOMByZy7
5FJLstX/GzoqnyQUWEfr2DsmaSVP5eBl21di3X6BqubyeheWFUyIbxr/B+8u
nS2neJf4MELIWZ+csOAM86a3chvRVuky9eO23EZo8l+5T3fUHe8go7WLqe7C
CPgU9bHyREDdCf8SF4EkNilXHFRI06/pxU2Gjcz4Se8feVGBL0x/kWyz99qh
thk8h+aAMo5g1VKhELWiJ5zzK4pX5ISYaSHxAVHIS7BPBzGFUZiFJEWDOL9n
NXXeI6Aq74TmZe4XytwgNc1BBM9oKjncTI0d/IBhWxr8nHmhNXSOnrZ0B5wj
kW7lvcugVOsZDGexj/A2EFjAQO/E8vLSkLYvZk1uWUqoKhwp8VTYbyPybTjk
bLAyr01BTSfMGCjKogC3+iGNmak5mrvr70nGhXRUbfPgfw0YCC2V4e05483j
Wkuubt6VEwsn9wBI+nyxuDA6cecLJFDVI3U2Fd+sYARyIQ84YLOJXtM+yLLH
EUthuwrlOpJGPy1Gh427YAFTn0wr9E06VFxMjC2gLMRxai4Axxttq07ohXyD
Mqb7FltTZGPXvRfE+ZZvmy6RsMrjlJ7RZP62JyOFXb6tAQGJ0+919phgbcS9
EEKiU1qZgi4ZFsohkXOig7sB68r8g9GnDuQo/BaepXHTDBVwZQ0g6phXGowW
mdETGakNLdrm/5ZxJ+wmXRM9pFUYjrtqHN2t3pCmGuYCnIUH1aU+GrcO5Nmp
+lYcpLdtw+2jH3VBTvPuKJAlNKdrwOnexaNCK0YdqUNHZgFlUJwNPCciLdTk
h/sPhgygVRIHFZqWkQOlINut2cEJ66U+qlpzoJxowtLO3GRk3fB5Pv1fGGWv
zNnzupf/mlVlSxVWARw4wvd/sQQfdMNey/EAZ+rFL0O/OYqxTTYXdPRis8wZ
kRH9SBSDbhnO1LPd4J6krAQ5cN+brl45Csrn6Y90zGYZX02o2Un5Z0Rf89Un
XSkpIry9zw7ZWqeof5KE/7FVN0NHy8FwprjwpN4oGq868koxP1zewtw36Owh
hwE4cH7BRrfArFK3NZVPfyrTx0z98OCV3aMVZdGq2x8cldrXhO5WYhvqA5Vc
M8OVeC6hDZ/kMk8HiOTpPYoS96L3oLECGTYY9e2GIxKrGqy1PF2pTnkeKyat
VfEUHyZW8Ewx6iFwY3kqeRKATNcDPmeipeb17kVwjs9fbKmxl1RVjsm5y1OA
ktJd4kPKUa40x8TMuuSpfV4nCiKimuSOAlEZqlr2aieaJeJePhuLoQoyGqxX
XQM9DX4z0cfca7r4lL2phlWKu4NWZj5PtVu5hyqAduVd99x5ry+r/4fumCH1
C6UbOHeKJZFt+gojp4j0jE+67B4r2cRiXH1d/Ts5SRHtBBiS6S8/3QbilnDC
48aiPJVJOmlranvybI+xxqq2LgmzNum2A4qgbYBxY3AgbZQ3MdIqBjK/gDzj
Z2JpSSJnvKBl/PGjy19w9rqCa5yBVcI8DReiz8A9ah/X0oCDiSgR+/7ocGzE
rwCTZG68C3E8oneYJNOJjHFaVVjqxGbgljf07sLf+5jWzFwLP4FJV7WJc8cU
lvbAqLQUZIvmG+DsMZXzdRYzvS+77NYRWCNMG4/SNo91A5hhi8gMop2xK8UF
DGO/whICK5Msq+9sHco7uD9/WJ7mPPZsr4uW/mDm7PR/ZZRCfikKrSKQRYjM
uprk2si/d/vtbcTzWGQz9jrHQtxIGBJiPcHZluVPJowTezr+qGa6nMwvPlA1
mYcRFwq3i31lVQ0WvS2z8pgdeWwbsRsnhRBiwT3SjJfSsV5BdKw1r8V4xLoR
SfZU81d8m9BxJKN03X8AWtTTirKZ5UNdzxpw6uSQmW370Ogve8U8swd3jhdY
qDmAbvnGDJg1W1/hJURTSMQL6kk1NbvJfFheJZGFaRBNNXpmvVmro+nvnAxq
GfRkBfhY77NMqvDE1ZccWK2PIdx+nhRqy5DvBdkiwxa1QMCSBoQ4XAaePkFy
kZAgE+dVaC0eBth4J5EXJJXcEJLHVPHqqWpT7IoXs4SON55HdSAmWODjC9tU
0SSUxjqp/PfnjRlS4auIfWdFn0qIiAlliMU87bQ80u7/+4qjBquRg5YQJJ0K
B99cd0QBiOCIGVAiCG9cUBeRhcLNCHGIhHgjFU7r005KcBfMZ9iIlN7zSQFP
NU5ZM3oTbhIQeDNVUhtL1MisiqusdpAyoEspXcCgA4GU6CmF5/9sW81Pqo61
eMppgvdzHn7q6yeyXngM6o1Y9UrvZgp0fsyfPWYJA9XIYuM8nBy9Rm7SSprt
z6yXTTCV1WtOeqdDjY9CKyx4eKaPFrYNdooY3dKRDpkOrBTKiYwECDu7P8IK
6efzlKAflnuqSmX3XINy4FKUgIwkMHVzh8uv+Iin3bNderfz+4aHCBfT4KP2
cJ3P868cXxKlp6/KMdxDOIkH6Lc4TyEVnsUCTCbmM9VO3ekpboXX6yXz7QQt
wKTV3+EQHW00fhCoHEixYV0o+Ci3B9+E6DzEfekNNhSX//m1NRZtpd1B3TpL
R8d2kmd1ZR7zjn7Vnlnq1EWC9SNT9E4MsoviHm3CbBWZpUjl1K0hLlSLbMFO
GsYUoKY2YDbUfE2Rb2mTHB5oQhvDXDM/zYF5zqYAZr2xCNCbTao6ZPLs/5mZ
k1j19gomLNUnS7KPEyKsNIBx3WWYiEc6NVCwmRRr8k6VUyK3Tub2zpNliSBV
pQoDor2OU8Xm5K1JQJ+PKp55Ndw5wNj68Ve4nqV6g8cHrs0qFpzfVkMjfctX
SMoASm2NmhzOvW+x6vDROO96rpdQSLcVhA7Njq2UpiayJrqvYbA69tKN5yTW
fMEye6TCRBmfF+xL6EPA4xh2phzbc4jNlTUoNCnSf0f4ylqWrbderUSai+Kd
1G5h0U4wY1AmOPpm7BjsvzhidTuFs4gvkw9uqpTQHwNp8IO7BD5JY8ESFviq
G25noNrCres+35Apz1dxRcWF94rqKU2P7v4LEn93zGs9iGx7tNyyyKTHMTYK
/nbffw1g4xUY/u7twChKeKvon9Bk8qhiVKXcEmuly4oV0aVg/lIBDjdyFVcW
IU4aNQunvLWswLxqIDCG8FKiTEV8VPfiRa4IyE2TfTHBzro/OqojnqIl+9Cq
epwqNlokPgwcBJWbjUj9Er7sIkDVDJK78SDwEkzS0Jng1hvmhupuIlh86i7c
qek5n55HpwuxgsDdAMR0H79h5BxAlO4wSfJA2dLyOs7f28N/k6fEiGYWISTo
SfvSlP6bFoSh/fDsCkfReZ1Ryw4jnaNP0WjkRopJnSI7t7Jb41vlNJWzN3ID
GNIIal+F0ZWhf0c0DtsNopINnhCuwc54WtvU43A7MXjoenUioju/Udb7GIic
iR2RxWuj4t7HhqBGKOVNrrSveP23YoS20/SoFCrx2Pbv0QIz4ESazmbIfK0H
fySze+qQiuQ2Okv5RbI8gULLi4qbPOm8FuKZ6oI2hHFRdmFLpuxa4DGzxv0L
TDG9CDN6vL/qCYHhcsO67RobvEY9W4Q6hz/fxWetM03ewUf0eJOohkFrmOEq
ts47lALkrMHd3DLxxv1CI8X//ahMiVsAxkuGDDA7ADazTaJDYlX1iaz/V5vj
m/hXL3nssE2/YYh8IuAdT8AwnH8gfZosaCE/PIURlp0X4KgDRr9315OCbU9t
ZPborL+AHpvxMlhaN5FW+G084OPx19ixyANLgO10w2XQ60k3f47Y5+cMp4xJ
kyTPsib0Fl1JZSn7RcdpiCcxDKsYrihCp+TMuFCcHu8Pk6prJ1kiFoj1RbJ5
eTgL0xUenDYVaTZX1PzXwrAcv0plt6epMKnaK7UhRFeXUTmPK+UAb5yIJz/f
vyLzqY588JEaIMOTgc/QincNAOlaE5oyFFoKpZw5CylSlacJqUgMXZyf3sVD
OaYrvV9VDW/NEGoMLu5jiDNyQZn5PABsBrDbHlP65aZ0r4iyHlUFz12RMoNL
/nXjUf0a6LSIfaw9GL7a+SZ6hWOQPPn/vcZ0BQQgFow64Z2hdhG0Ro2zcQCl
7O85qD01Ywg7jLb413zCi3JrXUB8TafZgqPeCJonAp75p/Ejuwja2kGrf/7K
NQWNGmMO0oTPxJMY81ZSm12drXmPCmHbGmJ8VIzWl5imDsypoSM3gYeUYBDi
1xrcszSA0BHssSXdcsILp6EJPIUaBQ3zJvWX9eQ9O88H2ulO5LXBATVbtulf
fVjwbaAayMtUqVu4OkGkUtMWZ6/ayfDuu16xWM1cDW5vaekJoe/WB7AskP+F
Ugigz+5+9TRc3KVTqt8y2GUYcjXHIEWXb1IjCuh6pPj4oD2GtV3bUQ7mun/g
4jtUMb8PHXBxkyZkyxBOgMfEzMHrgSWb1DPmZCmHWV2Vwqcl9HRGwmUswGoW
xUCidXpP22PwkYqlgWvq/PYcru3+srH9IkYsqA+3HKNwP8hOkG29gKAw1CsX
0Sx4y3XHltUXD7EGXbCtjUjykk4ZiwnthWctmFzcYbrV6oGNQF8G4cXZLTl5
jzpCFsoqjiE99MNeVVbOKw0d4KMSFVBlUxsA9qigjh15bghMzAww/70vxFfn
GgUjDYRbOAyTVOGN0wZVhZk3LP+YUWpifK/zJKWXyFHPokPlV/uqSWOh9uF0
mJdGL4t96+Yt3L9o3i39pAjSNo2YNqvGJ1I4sk4khe+PpYYQMeXdaBS52XGG
qXAvZXUTe5kjnC4Gc2HGjrG1YMbPJOvgGa3BO6vv+oW5wmdLldMExYrAWqWA
oxRevIx4EuoIN8cm/ArHP8fg6MpYZ/43ODYAUZbR9qHnOQkURuefu92ajJfj
ZctjxYp93yVmdV6U7khYbakFww2BzcIecJjru2Kt6EtwvSDw7GGoSkRpMQNw
3LyowybvF5BaHiNbdzfFKSb1vNirF5URGK0jCkZTZGFyasvz/bAFpi4H+LmI
UktkALOab3u6YJjqowjTbaUZDVtbiNsCbl03j+EHUyCTCe34bZ908FznrV2L
naDD6k1D/psRij5/M/3nz7EBtYAefNvUpQYdWZ5XxT1AkqjDqzixp//Ohvms
66CW9uIvNWbkS3g9qPm343usWwMBDUdebrZ5L99Vaj8V/xE69PMGji6ICtb4
IA8NPBBT2/2sA+JQkqUV2nIC0NyBkhQJRgMlKG6RCGBV3iQGmIqUDSP4/lHl
pv4n6Dn25wb2beRRSLdoU2H0m6L1PChZTH6ILEraIA11+s21uLRoUelCNwYJ
UVzcdj7w3ceFc5ZA5s8QL2ZhhZ6E4oAJlNWKkVe02tee52+3EnhoK9cKAFoG
hS1cTz7kb8B5iRi1SRJPdLxrL59TsbHP1L6Kk2ypuOlG4hhWT8/CUws5ncMS
8hoOLd/7PYbwQnGVfVVpfzRsiGPrx/6jbXWx9r/3A0vemLAuttsqVM9XZBIC
+/mqEPCJjwFX1HSX1Z4yo29KLRrAZzhAOZ18E0aksRaIdAk2ZLvcUVRyGmNt
xK3fTKuVp1Wd4wvBQkNh5Pg0lg5wOjqMfVkiF8NPEKdabnWPsfC6kieLGe/X
/Sc2FE2naz6DOSHZUSIMn9V1LrR0A+gBKiGiVSA58Afbyvde5GOgOyiijmST
MeeA1jJ+lw0e2CSifhUxy5bpBhtH1B78ptuloApTrMZJvZqWOctjZsAteFcr
PCWeckm6v0xGV7L+E7SquV3jJAXQPQisIZjsR80AesddOxFLoHo3BwYefqOS
N9+P/euOr1H23wUi9X5HkO8XJVTpZGp5jqrqekt+VofzaJ88yunrB9UmpEzZ
mB7zAi3TegZCRVX810gbE0TRfDGHps421kWSF0ka8rjlX3Tv5oJXTTvAp2W2
BTtlTRt5TwwVlz2k+fQWzbCTDYYMYH4P5jUPuF0L043+h1P+XljEcTJFxz8t
KB13vqIdULtJThFZYgdIMABde3YylCcqrCTbZsXd5bYQeaemRX+xhpS6Vha6
vW2IdX7rRPWQifKDeUMn1ZxzhzGxnuZcXjjYaA1epleD6rnxOwpNskmfwt3D
jwsNvWRUuTTyh1dC42EnGPT5xY6q1aqUI6E0Fnn4oZuGVPoJ27KwCX5iPm/x
xu5MWLc6BG6WHm62ghrqCugr9b7e8X+amL34SrpwVCkqJy8bWFAsO5XgQXjM
JP2lBY8hAlzz43gTvgT/LhQHWG+XIpyTCctUaYczskGAXKgpsjLXoLVimK36
ZIgkGeWpAIcimVcUapScr/0nw7lL7Jk6QMBTeI4iEw5Vb7pV/AvQY7+IADtx
WxfzZS0Q97VaYN5Jr4yPwYDntoMwRuVpmf+MBxTSOp9Ozj/rMIzqHZ2QQ0Yj
maajKhn7PUyMNTr9HH9LH+46uIJ6OJlmz7pP8ANJPaiIgI61QfT5qNtGdKo4
QiXvPRD2WL73q/EpM4DM2EOwcps5F5o6ziWO0H+iQbdiAaF/OFBQxUekb0vp
BGE+DfthcmHh1iTO0pvFPJ/IoeuxAYgqAIesofXBOXaYQZJRRpSEs5lsAtED
YwCINO2feOUmkHCzuWpv0jpn8E/MHzRhafvhtomt+4XS0hq58Y3jXrzSVyHx
qo6o6nV8hz8qkEhr9yHIqOQMpcI+xRWdKXjMdCvMryZKnt58cgS3DC7QJyDU
zyU+AXwE6O3daY/rNZn9RLgjuxSzoeIxlwxYbmlkILTEwyy1ILvN4dJD/Ro6
8jPAE8cgR+O1Z6fwZxZm+G+oqBT3I2JVIWCvrYKBWdzEhF5BnuG2ULLQ73cO
vmCIqeHolL8IbJ2WHaWPfvY6yJX9clUTuv+1m0yPghfVVTYoMmtUlq+7hfLk
PD2pS4fjrcZ+0xVWRpFo6tNWAPlgh9RrSBx1O2RtanCAkUy5+bPza/HVUxOs
6tadZN3Ea9WW13H+SNo9ArirpxAYJClHHWmGhp+asYnS03scEZrgBn3pASxg
hvzzDRoRs+x8mWIXjl7J+CdwDqwkleWWLP8BmLoTYXXqjOVuYaendR4BVUhH
wH8hlJ92d2zWRWQxwQUFovKFXEwOeObVHsGgzCXW5ZIVuk6EWLUvrqbSHzNu
iiqjGszOsQfRGahZU1WXjiogSoy5Cf2FByhySaDSb/k+xyryvm6tje8+qtaY
fVna9riDaidV+LGMamuIFQl5mvzuxfTaG8lpdVWvBsMXFWdDk/rjNMB0YeQF
sQxWiVp93kxfCRq4AZXLS4q8vwugLZ5I7onKUjaGuAZ/831Ga4F5+FigscWW
yr1OWpnajnuFA2mMCvS2/Hn2Uh3tyvlhmfXHaT6K/yZyW262egU6G9AofZUW
AQgebo2ndfqLKbnct+iScBMSjZ0YjomZb8zoXNRrtZJrl4n3w4Bygspg2aT1
VasAd9hl88GJiPSzRYlX6fV5P2OwFao7pZ4NELO3MRfm6N0h3jffeugcF4RU
5UXIhk9cMD8H96fDUWW+Tq2OkKhWZIf9TXI48wbgEoDovlzQb9fDyCNk4HJo
g1e0dPvzMhtORKlu1Q6VCB4ruBgSYpa5JMZHD4nkC1KiBNn0seSjIZmG5Abr
0xxaqeCPfYeMXeqPNTm1kVzQjlhElIBj6rMgPEddsAHC6/EYALPyLb+/Plcr
y650Gy4rc94xGdWBEaMdmzgYhT3MqKFYAbcTb+fTCGubUML1RVq33Ohmrh/7
HFU7MAN8nxCaenVoJxvdx8io/gk9Wc3tv04aHqe7q/pNJLFyDQuw5FN6s2KP
oC1IZINC/rqmsyNZyODwvY+XqqhRmadXcBpcqNtJ1ygwRfvTtJcQ3g/UtjD+
n8DJIJiKumAfE2RlRTwYMh4Y3NvCHA1SrTxsnjyTjXeUJotlH2uJV/n2MrOx
AULv9MJmtKQZS6nXICqaAHJPZMYBLdXM6wUZYvoT78LhP+IFVXT5+skuKpYw
xZIhSS7l8sCHQ8jxXjNwhoyioVYTEuqOFhNR1FpDSwzRTk9ayh7pmk4MhR0z
RPcEMcqnaH9IuiHDiKcroAtDGcbG9QFaowmPdUy7vC4AEKmwQx0UDruI/ReJ
YHanfghnbHwyNaQ3bmW97IqGGrzjgzdgb9y9zRLUNd8cWlLhttEw1l/NvOvY
gnJeAgeKKi111N1VeWpBLj+KjMtrjdvTZRUKh7KvF/1ORDdmqAIEZ1WT0T/M
pjb/rXg54EUFsUg9zgs2v6SyCXtNO29VSYDL66/q+y/MwHGpUKyqtDaVtYU/
qYMRX4sfB11vqNRmsSqPWyWi2wn4wzULeJkiUgO+ONTPvY7Jcdd1yfloFjRn
dYIvkfXSJb9A2nOozAme1Gc0eC3CXggYtjiohIW6S9woQSiMsaI4WyplkLHo
zDfRXA3GE9ZsO6LhUge063emhTlrqzlyRMbIOE/rH1Q0hwJZzQRBo7KSjqs6
EhU6LxF2hbObk0Gg5daf9ismPHDNluxwc1tphuLB04L2BUyxfqB2oGL7ys3I
QeJSOBFDrsv3PqlZVIMzNloomUAG5FKH5EE3ETZft2Ln2G+qtUyhTvIcu3TE
KWQAbF/Q72z5vWfyngEIhurjZIy4LKjiW4O/cVEwjBD3UVIptn+Fu8qXa37s
WZLalkyQ5h6Sf0lCTW3ryjAk4l2O6CWwAmV4o74Tav0rAi9To0nXBq25PlNp
QMNWixR3LCkklUZpjh2HpuO/+jSNM3WFPq6fVD1BIf6vuvDQmwHnKybEervY
IgrwCrAKkv8BttE9A4qwHBba/LVhW1iHbsVzfpE3a604lXOdRjEPPA2nJy2e
zLdjmaOv19KkKSPik5gFJxTFGhcS3PgLx+PGMizZX8ra9N2spDXku3z1ePZQ
/BS/ePze7E6U32uT3aLYFMzsbPzNyNdQr7MBRubUiQ6g29o6Y/IQWwp3pA8X
zCZSzUJ0ymyyWHTy8NI5u3gmWaPM59ofx8M3inlPK6pxR8sWOTvceK7NCzVZ
YN2tEpISTqXVQL+M6GRY/AMD5QXY+I164UiEq6y9uRuyNGq1XpK1tPUhdWQX
qanDADCwRzdPuCMy5z5iQ8eL9DGWESuIzEidDAQksNXfT3347zvPUTtfufE6
uTur51A2e9UTU2ymZuVJpvKb9WRU08ni1lAIKppz81SyN8flSd38bhrIBuqJ
Y3zVgSBlW3yDJjod0WcLXqejbm1fNXgEVuoWnkqjElI89340bu4GulaYy0aw
+ohizheJIwXFl8Dea6oJdvXIrGF71caru4jB8Nqkq48rsL/lo+/SD5RMbT8r
xpWgmGv/Hay3RLigrupTqyDD5Q9z34Bzm6WcGPoNDCjg55bVrb+pocfmkbuD
EsXAXjmHLHPXW/x6bv/xZdZv5ybOHbR8Kr5Y93KnN9VFL3Rbg/OyO0uQ3xKo
byU3EPZcpkVbfwmycvaHyhTO5F4+W+up1hKaPC/4Tzpu/Foo8BFqSNJc7jjL
EcHmHLha1kxXTRM5EmbnHJFaPiWnGEM97Q/nRyc54CZbX1L8syC4HvzkwJGR
ilzA96pzVTkNRxaHRnViYCDrXv+FHkrd7rMnOwPH+sV1a3QMSXAHSCFXl1zs
dXOwKPWIMG2Y6emiqqT6QzWZ/KtVk+d6hv1uTK/ZgxXZkcrSLGUQOqNZ4khb
YkpMODFrhV5OHQ/Px0uCErivhSdEUBE4qNR0EJZm8viy/SGPUkO+HMfNArnj
DbZLeOy9cu/IaeLmm6qkq4S4WhO0W8BDy07eNLvSRQZWm+GYx3AVt7aoBeM9
oUz3h4/3bJnygRaHPdG15KkTHtiyzaxsA16qwjIv5BJS18Y6KfQh7Xzg3JI5
Lfy74u6k1r4fYaN6VBqf1rDWnv+eFAEHBMEsk1KtZR0nqfxFSULLHxeMfFfv
egbnigD5k9E7eKjwNim4cgb0yx71M5aDdrlC7VV8KsdztC/JyZAVeEDrnlLL
8B5Le7OalNB6gHG9A4UbwpIhKVppdf1CTX4YshgjmHFG/I0W8/QnlNqsxJwA
NipWRXI/1XyqBwiGVicZ3Kb7BdziFB38S3IP7X/BJikpEzmAopxT6M3ihiyA
Lcr6nURnttIzhSEw/aWQ/helWy6gWOGVqx/wg7rXFYHAhyQlk2V6MYHKpApp
dYq+6G0RZ/QPJ0OSXNhUO7wLJEwGrC+xR5+hrHQMSdwhJVtG7OS8tNqJIrsu
TnUiuPikbJpHHVl4wIO/kBs4d9q9B6YxCWrSJCOl079awix/hXqBRqadTHaQ
1IWSYuz9v8eM7sEVFyGNv49qs16RXvw5Dzzeaxht9y1nIOCxmR8NOuqD+l9v
MpZs4dp1y8Q5hPBRzr8OmlG9GOX5KzX+vR91Kf+ri4ayqOsIwL46HGwJVw1V
KuupYlWRN897QbYye6lvnsCkbE7o+fbxkhqltFlyc0mv4QR68DOwVRwy1VhV
J1QXZjZYfZ8UQFo94afznZJh8REk1+WbaM9oMFx5fUa5B05Oz6ihzk68WGet
QT2sTmlOpPijlufSTTA8H4L8M3o7vw2TiiW1G6UGIkWI+jDPjY+daH2HFnWy
g4Xo2Ln58G1juWxsOIEaVqHJc2koTwBPnQuHXyUSDjmd8HMtdVo12CxfFmrn
PmXmRbSNAoUu0zcRrXKDMHAiCkk1BEoEfuoC0vswoNBnhPsExkMmpPnjFCHy
yUM8knxWSuKvHzXGjbOSXNefQZZzl3WM/QbwEzl2vtyymOW/70vY2uakqTbZ
C+urVOiKmbqj2WVHZt4AT2CHUeF3eUdej0QTvwWEIiBVySK4bFIA/2V9//gn
N+LAmkEpLCeVal01k+fQ6lru01Yivu8pCx+lZvHfKkxR3E/cqyVjmZOZDf/E
P0106p/CMykv6pxNo8plzPl8VkEyzZu6Qfg/G5WeMOcDFljr2JOvo6PvmKLG
VbCtFvXU1IOFAONR5ewDqdNWsKx3EGnvyFXJunmRx3BU6I49s+L181sdq8Mi
C4HVYS9s6jlNMMl0DAnGvOOi+igQrlkP9D/Lazj2hscEIwtcZfDtmjsekPB9
7ux/3HHWujqNl2rm7FsIDBCwe1xZ1v68++z7B+4kHF5PuJT+U5pwcXmZ8apc
E7J9V+r2ntPsuTqoCzRHr/Dc/Tqfw3Nl4Go0r4WRvIDKk/grGtRtRUuiiZUt
m43HLDe6k1gfs4a4YzzbL405s/6tccOSoS3sNokp1RxiV4UZ9mSpZt0zIdeR
HcV4AzwklOrfNMTcRjpTiTz33p41b0mGBFLIZTmhUcjANHlFBXHwtA5mQ8+2
L/xFbALEXMTNLIXgk0u7a3+nsvyPk198X5eofHHeEnURAqv64VeC7av1LFVD
X8bjVIWCzGGSHyfx14F04WwknjZusYkoIXuL15BeaOrxuHEnupO0Z62UMIVr
u9i2hSmCrMaBb/hcnuGg/DMxPGvx6FAEbmE5L0PAI0SS4YQLxElTBPJeZqql
cjGq71HVn0rVoXiRxtrwCY6G0V+Pa0p7veISYb2c3i+kF1MG1Pwv40dVS/5V
G3TwMNhZldCVvG3ltwaTZt8r02955QA8yVSEVIYyLmu/utMUHTHIM5UV/M4C
yDH/LUtlmUm3U670pGPKY6VC5jlnPQrLfmnPAon0Nn2DiUBVUsHvyeYIyPZs
fWMTAie8vMPQvFpZ09eCJj8bJaAq84gl5O4KlD3rMkwg4HWaSu0QONXp6Q+9
J2f6rQpGkVOs3s1ugkv0X/8grkIYq23CKBMytvxzPiWiVtRSwKZkz0/1NRAE
9/Rlds5JruC98sr1z5yUe+GUnCL7U0fUPNMazLoSmYm0q41CTOsdQChGTpMo
TYiFeN/vxoPHxNhKPSedIPHcCDwXU9L/bIjhRYXFEFGMLDgoPbVndltqU2dG
+qIWqpw6nG9OzXCDIrqi0kz9a79GL5Gt0qJfm7A5KtAzImj08MFSnUpw7YGg
qAK6+WjMEWTLpw+t+VV+BJlSdYOtL235qh7RpgteKX3UKTxFPH5PD8jhNlZy
OTSDLyUC0SdD3QyYEkliJ8ZkN/22TTM0N4dUIr878XYAfNOhzJRMlYYIZpuj
xmzCfVT5KFKloscNQclB0KOlKCBBaS8CKKmd/fkc7be5mvtQ4IO7LPZhLh0Z
4avXU6HQbyHtoHpJsaPc6J6g3gHRfjSgHMmTPoFo13N4pDwDkemnRRf4krvR
OKbPbCmVUrmSRS2pzwTEUrRUrk/+UTnEOXOPdwKSYHxE9C7X4qDxSz7imYKi
VdmwX1R/ooh+892IIdi+cz0VCJqNuspYAAx8sdA9TBGLEs4uh0Jh2holXy9G
iWkbzv/S163INT8wCjAclQEuiIL111PGber5tRTKR3f8CW1Rd3dx2YoHsNWq
1skRjrv1tuA6NV0ePvHRi4BrUpetnxtXjis+9l82QVtuawuhml8e7QyBh8wF
CCFkO2YJPHfm8jt7X96o3YNnDk2lB9aqNFqPjSc+SOV18NxQY26nXF9lLeLM
hurS+XTPBugjvlsec/DAY8F3lZ2cM7ly2ya3u4TzyMYKlkwJ2NBqsVP3NyuQ
EQfF7eWSh/2DA7GwHCf+xnm2T7K03oO2jW+rjh9TmSj2nK+CE5ojXNfDYTe9
Nv4j9kzQMXO3onJRb0v+sLaWCxh2jYjmYAMz7/tYTSUC8G88HXUjgK/2KkNC
qx4fCyl5CyVhpwqa4X03bXvha2KDjpCphmf91tkE3SCp0VQOzh4IvkhaMzBM
gJP/rRspzGh1b1daZewhsaKLJ7RXjcPAXCpz8FCN1kTnnTlcZhx4Vwpr+IzB
tyXqC/4OW2FGvwsV3XsuzePj0MbXJOGh6gL/XpMdg6nyyE6oJ6ew66F2exJ/
f5AhpWwWCore6Tckqx0mrTMasalBwepRmHt9iTSjAI2kcTbEsRvMry08MkSR
dNK3kdK3ixWfZpbZ6iV89xG/Uurh4+sdEcJhHljIyIFHu6O/A+41qLoO/x6p
fNtSaI3RJ1urdhqNZpVJhvkZuGtHYVUYwXvL4IOCV6ljFjRkkJ6Jgpjc29H1
J/MAQwSw8aaQPW6TUtgRyzNOdrGbAIM1cy3WeDl8i0cWkALthN/BH0erlRsq
/ZF+/CluOF0rTSbfycHy2O4u6ZIUwyA/5F8NNUZCEqWu12jMsALN+YTkUDXy
E8772QdPP82JoqecWaEGMd1aYLklj3JPm3exK1rZ3DsuTGOifmjje7VhXjjE
+fLMzEVGd/4Olw1WxasDSLRJ9usmz51zogP1iooQ8YQ6no9Sjwy1Sq+j6zWN
jBXX6Ex91KAtCoP74aa9x6rUlleCI6v8U2EaPLerdsJn6oG471lxytGee4qX
tH2YrLY1UIDlp/OR7ixGk2CVR608mkS40VB3A2mUSR6l25wqwcBWl0kfw8HT
iyf1w/iOF6dyrOJyGiy4sBT/dcz8OXbmgwoUxA79HtWjXC3Oh9fRmyJfi4ps
f4VwweMvxEwnKx+rHxRs0LT30wGoYJ97LpsZCkFOfnjcAQgg/j9wyJkcKfp1
lM7ZQ3E0CRYgRrWq/aKSYoK3wuSndPBsDiw8eU55hJjNA7C6hfkaGhWSz5Kj
+/U9jj/R00t/6isfof5uDTZ7WwZ4lsRwGLpiIQ7dWnt8CdWHkVVGGKyqGrVX
IbQmQ/CGdxQl6kBPJHspO/rr27eSecuZgvX3JlXuzTT6ZZpWGXzPM96xH/dM
qiTwR8F1F9ttzPY8pCciPLGK1qKWZkZ6kAaBnBNpvY16fdYLVKUoRx1xlhON
xxsA0YKNYvKnocscMYrdbfjn0GD7wj0LUGdh2TjbZalBIhnWw+OL52XQKulL
TWeh8DIGEegU2Nf5As1hcMJFKOSZRBUk0a93z5AOuoQTyzJndLkDbmmy+P4L
xvlIn5XNi1KOiezldgq0GopCtYKkJyWL0YqzzKMP0ZMgWD2usOiJi24gCHzb
SYmTmFnBKE5SzoLNrH5hS/qMM+AjCZvPdP4lIhImA+o8wHGGwounGAO/BTzK
M3zi9wC+avqexy4GxbPjdptnrOHUtxrNGKxJvbIyrE4/A8bNznz2vvx9hc/f
BGaNEGkegFOOLEEeB7HKNCSYaJRcdLx1tAtP9Up7zc4APYWTOwr65Nss+RgZ
ag6mJGvl2SDiNkit86aFd2l/iPbTwQ2HYnKbedq3pJOb9xAkJeqmQ+rWilnP
a1XO00NoArYuJrqdO6aI+mudSJLP597j1NKrgCnqK8u7lKbl2jtbpLJXnudt
+7QnY/zUWV2n88nPaIeZzhz2R0/SVB8r04ojjkehqqyB7Cqlr/NgnzjX7xRt
fdohL7fRgaz3vVwottuRBUfXOr97RpRlCqjzoqJBu9WHjazyLDEefa3E4Mac
RcNhKGflCBwxXx2/G6wHVk5BotqoVuAE/IzGwD1jVSEC9L26uJHUhElZxWS6
36+rCRIPg9krSxlaSff0qfkWGzVgpTjt/ccwLXXHcCaZpMfhAZeA/lSlE/IC
mfnf1kboOWPt7N7zbJhovFcS5rGOmlIWhXvGzK+Y6Jo/hll/JDZR07AdU98D
J384YuGDW6jsoG3ZmHDlbSYgmgG9NpKQ2zqu5rue0nCGaIv+RPEtWlaIGgUe
q/Li6xGonuKuHCoHXnKh0SGUEfXixaRRKuQgfv8Nb9Iagk9OdUGdeFxUUDr/
D9Moy57RRnxvhk23j/rL5Q81CwIdr0ejBikGQtan4yMB6nVwQse8gd4zYrt2
kEFjbOEmEXs+lK9FkH/ZT2o7ZCpyAg8DLndiNlbaX/juPS/8eXCuSrqYJpem
DRo2i1vt7XSbyt/yfy810Cm3VyOYZEisjQpN55KUxkGKzsyoG9vskVVRW2r4
/dZF1u+H0zo6kFIgYHsABpsjUDBnzGi7zG24EZMFr6S966pvxAHBCNZ2RYv9
qHdiWyQeTtUN3t8FTrx3Flugr3owY0wVpk8Ae5dA9P74mdOOkLeentyUKyFm
SHf01LDKgkxnW7dk0pUbo1dtvGhDmDsmvNGuLp/w6TYCPIMX2eq69AC9G1xu
Ewj6NOQ3hWjeOQKVJk5pY9UWKbYDZ+9aRjp09RzI012jguypmsdUjPNgl+GU
S4HDgSBRoarNEC+oX1GArCZz05hIP7SpTXk8NLROmJy7MeO4Tc3fCswbDvtu
BQoKPqQLJQRL07Vk1s8ekUbnLOQqq1wQK4GwT237DrTqd1ycbw0Y6yi+VwOc
AGYCcB5uR0XHwtllGBgtecLLc8+Z61HRzDkcAi4k70Hekm8Kqezv3G0HJHYy
2jWM856Nrv8ukxUmkeXa+EfSO6RJf7ROMylsLRApO0FJ3ZEDCGJijctbFzRS
qyEmo1vmfcmAtu/pMedtZX3q3r6UxIIqfeQUZxxTJtjlynzA4jmHTFyJa+Cg
HfxwNIRqc4ByLRlwkJjuOa28m7qRUcx2zUbrMDIOS+Pi4dUHeGqR8XG99LqG
Zs3rhis9eb5fCCNcSq1kpGqDjCO8vV10IfIjjnlvigVaYwo0t/daUaUV9seY
nH6rZqCFBXvF2S8ENHfaVw8A3RBwNZ5JameW54E7aoTeFcuyKzIVIKBQJLZn
IjU5VUrYDyZwgWdIaBb2jmPG6iYmCCGX+Zi4KHPIEwOkaxRWidnM1Ye+u8dH
3s3fNaZxg6vDrPodIM1nn95TrH9wii7nm/ufAI3Onj/p1iNooJ3gaBtafgQ7
bPomHp77pNorOjwDRmpeQZiR12MPvmfabxCd4R87iDcBVbl9NBY7nGRP+9i1
egONg+Kqc6foTiiREkGuoIeBnigwN3SzC+f49vUOX2obM1dpnp4sMO7uZC0m
0yahikT+r1TpLHXVEcdFst7QPx2A4LQM3LYLldX65+GUJ5ybwpGDbYdGs63O
bhu0G/L7DMaekFxYWWm8zdT7NROhWrxA4X3IEXFXBZXzeVE27X8HVpN/9mzf
S2LyM8mcSEp6vGPLgHf5qsh8vWKg5pANNW7dAL/B4RtwlCXzYqmscJCK8AF6
ZoSIjKW4yPrS6KC5I9KqIhOpAM/tLrE+4+wxa5n807tM7XUmcDaMgX9qwaHt
ypSrlBrlSzhSCrCYDOa05yT736wfeum8E2BBhCojwIGPlHl7zKid2OYkyDro
5QiZTTC2nrG54GXaABcElT8Gy9DEUbLPTrjd2xXIQPmCotO8kcvUg446x3ja
SSZ8EJc2RU5p6jZ8gr/IpC4ge8XHyQY2uC7tNCuwaVnn7exHgTJkspTbTiCX
F9gKlWRf9E4XU5tjha2nyPa7b/5PMalZZ+EvDZHzYsuo/YObSGi7/1SZOHm/
xeDL1PEmpKQyQe25O/UHveydkeU9RWvt3uoghci2idznXf7cfwKT0R8P1KDB
jM1gGPAVvYznWrphxg2bJoSA9ENsGOh3ZBogYQdqV1updFqYvAT3xsrLKk9f
zoSP580SUXOxJ4s0sOhffdBHe4KGLBQrHYVouRJrB/Nhm++1N+xhggEQUpsr
V1uFBDHuODr/WCszUp8tOkP1v/AGDhnIPZYaooIX2ryc9CpXj8pZ5DFG6kXE
9q1it0BwVAmEiVm5f63p6w3VxfRJpZTmnnL8YT09ry+bQA9X81pbwpVXX7ye
o3iR86JWdrXs0fIWhQS//CNZUngdjyhaGWARq1GT79cDzsFurvYn9sOdc5yR
7LP1TUMqdRAd/qP90nz7Tdf2aArM8px94L9TNn979PgjjakKZN1/7+d35xkR
O6DsM/ZoLBaRsJfcBedkROW3+3mKxgEyPT5vYqC3QSdtBM5gIL6F83a5x0sV
OXnvDCGZikAgCfbQCyYhwlN8XO2P2iilqKU4i9/wfeb9+DzPXTNywkpoCUO1
cdpcRz3GkVifa75JYuqkdWlEC9A5rf/2Bmn4IPulqdHnweXzO7x1mBzoGEZ/
SSPnzQ6uPaXqwiDKICpFj4TD4mdDhPAHC1D1CGri4vZJuu0G9g5i8j+PIecA
syJ4j/MgY1QEc0RsR7Ense/EWhNVAWLUUQWDk3A+DIDvLTKaxEnclIiJzm/9
fuC50ABiQ2uU6ptZz2i89l7YxO50FU1VRWsT+KBjofvhG68IQX7YQGcvhKxK
i0yAjURmrMiRMfTieNNzdT7PNFCjYYNgzPPIf9F6lX268W9VKRBN4682b6xf
UivtrDoYRTewl3Vgzm6DAsQX7EqsTJ2LLHfsrhBpsOC3B8xcbRmqL3kYFKCO
i2FOawI3MBK8YE46PItg4M46PbHC/CaxBjRkBTYHQaMFhxbUWG+VWWzx7evB
ote4CSfBwmkveqAN3KYn5j0JTLCnl6PkVAfGFgHG1ww0qFkgLoLlXW6sEv1p
RNpQ/IFZ+6Ij2v8THVON/AJid0omO37MpP6+3luZ0q3gEsxhoRCPS3R6JqXs
jktcpvGLhcxc8ugcGUiC6qgoPdif1rD8PUil25cGGgLRVBj8WE2r483kMFhW
1m4XeGSerFe9A5/x45fGppNWsBzQVxJ2gh2puZLNhozwPCdmTEa/UfBpDYiY
caHJT4xEzVzu/gdDodh0iIuImSnxGg0AUty4ubI83A9ukTX6M6Nvzbc1RLZ9
VY3aMhjjJ4bqRn3u8BF+QhLKXGpKMtBIMo6Qj5cRraT2qbm603h6N8ViXQGl
M3Nj4NNqOYHvi41rTWyR2RCDh9AtgxMeh6V1spm+k4p7sFXRVK0uqHXZYrO0
XwW7UKBCfXYISw/JEJJtkOoWY4cTpxsFdp6awuJ9SJ7RLuFGfGV9IlFjRmpb
zS8KHOMu3VP2VlQygU1oQ4ivUwf4oukVzSA60hWlXgIceSXW7hkTxr2QODJC
xUK10HkEhrSESx80WbWDHuSe1lCA1FvngeZSrpl0maFDL1VvbG7oJvD8IG0c
W+SF/UGYXxwhu1JGI0CAGxipk56hr8KMxs9BbJ7bVTzidXfxweXWH8j3jTU/
z5pHsF84hInWekZcpg3xvmVcjK1g4JKu91Di8mweWkgHhtNB3GSqGbanYVOL
+h9g8wN/TnVPgj2NOSs/SUFlUSv99nO+HUYVvNnCdp7HzpmLBkpVrM/Up8d1
JM1KBY3TRn7VUcH4rn+xS7ssQ57cfMlNwNwxxVvjQNegxYuE+jnQrQvbmn7w
Vup+Rt+wq0W+JVOjUvl0/5v9mjtK+iLUktr3JlRD2WR/NVuWH6mSsm3Xy5w4
nF4RGFOlI+W5EM/zBzvHlb5K6aoLBQAbsUGBkf9gXAvCUg+CccewM92YXJVk
6mKYqxR/RQFVwFIMrOZrpZX171OTfexPa51QRDUzt7yj5tU1FPk+FI0kxnKy
DBkVukuySZ4KLtBjt95CzcuCsuQx7T7vyYo1ZXuOF14J8jJ0S9Es0rljvce0
JI3QgiWSL1MYlrHPHfPXj1Hgm60E6X5ECmhumGCGLPSnididBhFNMHHWMLDX
kUN5foUF/38jmUOf+aUuM/BRTpW4HcXqFIGyNKxOVUk8o2STme1h0fo8F+db
oUbvbCpftvvdIHeGJXJnD5RpHHTt1V9a98S2pTBDOKvEf2EqQadH7Wzgnq5c
kA97Z53jp5Blmn2lmD1HXbwX1r0jfQy7YCGd/ahNi+U/lPIEbd+hTRwadOz/
W6yqg1VywYTV5dtmcyZ6tMLj2BGCciTdi0behM/YTXjJh1KL7HAIgdIj65lf
PEMT4iXs4mj32WX9LJ/aNIscpfoAlQ1a9kXMguLTfzgeD/Cy5LyHxQCu8sFC
2sf9xvPns0rlnz7lwBQWysEtZnOKjS5qKuDpOWehXTsT7Jr/iVdIj8FKr3x+
j190wnAIUsNCaNde3l4RUgkkI1+nCCSOLTiKtHYGIXxNj0bSjxr1yHq5wbn7
L7G50ECjc5ca9gtBilH0gipVMCK/TsPcuU/nmwQqM9jHALVKccuONGvBuIVF
Vv8fUv1crEKkT6BKnQtk413SJ2127qqzQBk0MCVreJcYo8zf5Me3mjF8PmF7
uKZd5KiGgA4MZRtB4EnqKDGTuyIpAQoS1e6dgfQADfFuSJMNa1wqBLdrtCv9
YFQBA0f60yFtJF+/jH0+AhG2bJuxqcZ202oSeRwhWOlqnv3T0acBdkAGgO+e
FFo4uBIPvcETAlLvD1nv6v8sPcrgwEjWXmNF5CzzetrHVV7j8MMpCu8pDRPC
dOh0N23OfEL5InEglZyZXmSTwKrhLXsKCVjErEHVq3SehO7Cu5Se1SRLTnBE
1X8MTj+gVOmDINBhqfv5i3/R5Q/kYpgdBPtkXcUAJ/DvbyFmMgBxXHMY0H0W
TPFA0oZUj7ErOqwWP4s5gribQhYiCzHJNFElQDFD0yfoVZIDZBL7NXix/8li
PYcta0jTkHy/WX6fBAEhK8Skjx2ZMkuYIz3rSp5XuklgPo5ABu/2gxo/00ZX
bHqcG4BfoK09X5HmqXrHUtzMfgGDy3QCNMjzqKQ7H0y21CVYvJDoukTu51Jf
NuVYFOby+bsktfz23fmotiUDR0oIsT0wj8etQ4DCtl05QeOjSkeCcYhRtL4M
1UZrasTz9kyUyJ8qIrMfgmxohR+aJaswP+yOBycaLR5KXrFlTuacyeCW2LYY
lO2IFCH3p3tyQxScFjGuYEmJRirZ/EFunCuIJPk5quc4DiCdW7gD3pkA+xQd
aZi4bFWzk99AecvoYqijd/qphz5gnXK6yQYNhPYm7W1uvYUXtfxZT55uMauz
6DOaUKgBlSx7LFE2A5wxuVWRWKgnLEw+k4y2e3OqBgfAcXiyhmM3aqE1FZg5
vIC6SN1PI9XBCcMJxvgXZPdmziFFGxQyRd2kUnLSamm/WImT0rV8OOyM/KKX
cXYWb9NMu0QO/C5wR2FqkOtNMDNxeIpQBOZD2/1FHhbghxz/B+ljtSRwVQkM
3vFDTm3UjBFnTDZW6T9cYBxAV4bnpTq2HMPRo9YqxI4mBLwUCax4WE8qpnFg
LQ9KHxgKXr1MJxXA45nnt9AWbY8fQbFMinH5piaN+x5VWHhabkknX2LaReoT
L+LoQnfgoZelQAy5fedeH/yjxvmvaB/VlmWPazOpRzEQn5Em6P5UlNe2VuW2
S3JnqwwJr43A3lieN1kzDjaZRaJ7QG7Ob/w+hOzIklpDosHm/danTgfKa9cB
IE2aOKxyIN7eJe99MDcYmR7LC0iRTVOr2Fz7EyYr3tElMVOPNifqA5jrxBQA
SHW+0ydP/m/7zoQyOQiuc7gYO3dBJygJpvjnEQRWgHbsPln1mni6cU39SjTg
X5feOS1sdAOeVSyOScNT0Wop31VS9KELuP8FXeel63zZy4TD3HbN3XqIfxjk
WAFY1IMQPJ7ETwMHsG2/Um5tzSwRiYdzbW66kiFelq6zk5696IJO3m2sIE9R
pwgogH9lULatnVemSxprti+9nwdesXaPpSI266syP7hs5livxHwU02OlaHhZ
DG1O90LVMIA91F0gZkd1LSLThtHHopnBa7QtmPuupP27wgDv2RLFSysloAew
hABifhx2FK/bSzW2F47d9Rp5bKf6gkgaCC+jjP6PKVCibftuXx+LfC7wB3m0
6HwP/I1JE2PvvqZt36A5ZhPWSbEwOmkwAnixnvKA0spzwhaQ+ddQO9qy9diO
dBLdhT+V7D+ejdtHyMNUS1tByo/E1loDXdb0dPPRrWlWmWVUv7DetmR5J0e3
zO0br+A7kt0P1w820EOhmYPmB+Hz0x0eeMvm4jyW2J3fbz4MoDAbZHQ1je1n
/GCMLn7wq2fGMFe3mav9SnejTJPA3W1M5jN2Qz0DOz05HSDDK2GlWTiOQm/l
oRjWgb7ZGAaoevyGsnngTT2dmj4Pg8IcDH56tDkDmoj81WHKrxfCXhbl4EkC
NQdxnNoREghHX2jNxPV2I8U44QVaPzopjb39CuRgDvJdN2yOcOvC4wGIlO9J
08RLpSaM6faisBDqCtZpE65OINpAS+/ih7ONz0+MOC2kR9mZsYu/iHcy7xDo
03Zcr3AJnIuXq8nvHxEwjdcf03QRpAg+GZQVer+PEH8z5XOUGflS+TNsMAA2
nLCXRJ6AISgOZTv3bw/0KmJrXhhMcsK765+MS0Cp56RlYXDokgsbiWENUc4o
q9mHVcHeHyJg9/lZNzCGf+/EwekWfdYJL98Ueh5eU+nbpxkwrtsctRIwTbMg
Iif+E6uldgwH+HIT2mobMwlGzcNHxUHKYbYBKPvM6FlvT5uPWMC+Bsqzle8u
izwlz3jUk+EcoYdGf/kF6NJcy3KmU6NbKV4gRfnk2tPu7EbFmFTPLu2O5PtM
99ww/vPg85g874xO9vDYAZpHlWmibh2bqP8FF+wvBuT3Dze+EMHiEB0IXlsm
yoemI1+gWrhILedv1oLxRXxFs61/VQm8BSGdlJqhyXP6viqzeRgLQ9ZS0fPj
KekrJETjrPpyKXQLPFTw0ppIeaZDleF7zN89EmlubvcZVVMdrhrDx8cNbgn0
BbIvO1XpUG87KZk0DtGk8C9QbiztBXr+JcWlFE0BdyKWkLbk6CLRUO7awBjv
uKF8ApV2VzKF/ELt2qoaVfdldoMjxmmgLr1DyjDCypnHEPWYpWRc0ccmC7vp
qelbCKg22aSOHK68PCQzphUj3615lwF5PljinCnfZTi+0wMI4W2+ya8w/Emd
IX3QYha85Hu1AoSxHqgXVudck7StH2N98l9AH+KMm7X3BJuaJfQswYlJ9Ais
s/89xaewWbaZXOB1tqW0xQy+gsiZ0rcs/oQop/sMOOzVOhXPlc/votBFypsw
xle2vDRV5Jwu7nWMyaZDJD56Rlj4FR0OWlJ6vih6GL/qQmp/AdI/HMv2livt
D+o195tE/66a8QA1jCLUtudGzDBy5bVC1uJJBO/rpdvfOJvdkG29nDPqEnzh
enmrXLizxQTMUDx340PqtmkLsu0X2ShLYhySWkOQXIN8nC6IfgQCOS66BYlX
qYe16tiwLENMmz2SZeV4SZPLJqtHgDrt3Z0N+dAg8h6+s6PGCN9RQ5z5/q6T
GCKjxmNIrvdZ91BguTdgnLr9tDVzvY1Io+emVmj/fQbalC4vlt6gLawQCJY/
L/VBS0lXlM7lLC48lTUTDIDViixnGD4tRsDV0ayf+fyT98asmXUFR5W0iz7g
v8r8uLtj960XJFLN71r7jJRaoZOdH2fXWXo38fGvfi8cJ/V0ibqXv04DRj8t
J3btF8tpssZGNfaYM6r9HAH+GDEIohMY9MvwVGiOh1cQ+qCpThEJx7aOhng5
M1fGJzW66vtdb/oMbAV8W1Z/g3XanY6Ne7dol3yrcRaP4gyJ8dkLg1+PwAl6
C5hpGOuWaOz7y76d6wKr7NxnSb2fC3YQ+p4AuiSo4hFTKrwzOol68fwlrzwZ
G8FwAXnp/j17iejf7FCvSsWWPC/ZEF1LaZk0eQ6lbMHpJJMm4Anb637B974S
vKQZUlXL1ozzjK1uDlHixT/xnMnTEMwQGgeCgUdOe+pwJWyIPyVz061OJpy/
WLDP4erMUO4VHZnvTzzdT9uJ1FRjPgj51DzNju7UG+6iRFHmH5BX8fvlgF4E
CUAlrDDxV9IEisqwFbQKfJDhVyqpXl8HX1VDzcRbM8kTI2tQwd/vnnSf+DHX
uKAfnZKl7qqjduhJVgMnVo/0kCBi8wbUQ8X7LnD0SNQBPQOA87Ji6fJjTWch
ub9wAf0q8QrSvXSOD/Wtf/CmsxJjeD2D25CsnlW11Xo7BqX+U/r/+PdDQJxj
KKBxSmfujMEx0ulLXpdkVmbW02EoQT2M9OSCO+B+ibvC09Sqgm17tHrFa1p9
dEpIzI3WFVYOXhh/xzWwtd7xdE4x5GV5rycB8JOy2gm8JlZUGQLFIKYMUlFY
/AFdpIRo23fRRfCKLMMj5ycaYKivZbV/cJtZulTYhDgueX9Q3vIv4E19Xsfx
LMawOfHk7RI0k/vwtLOXkym+iddlZFDVFECI+gjgSQqMW+H6B0qeWw0w5fUJ
f6QBnYJAWbsSBoHkIIRGoa6vYqCuf2Kc4gHS51UU5S+t1Rv+W5Y7aJY7NCms
ZQakkIm8x0mDh26wfrlWtku2cufMUZb+RbP1Z7lrgzSEUGllttlEZt346t0j
1k627BkjGyUXX825A5e12PvOexRo5O7fu0AL2Jm7B4saGWqT3C7rrSl9c8yU
MgQpC3kqsyM/R4dVqHoN7VP+c3k7b9kSYl1Bvzovfc6RafwYjYzur1j84NEj
0drr4dQVbb0bW1VZAX23xqVUwUQ6E7BzSDzA4D5lQtrI7NEyvhS5b9CPwLXe
lcCq+jVe6AM+d4UmXXLmTnXm+EX2vPHrJPVdGanTCwy2ZOY+iQ+0M5kBLzeC
khaNS78vHmklu9DrGP08YtfjJkwBmR/KpHEB75/N9W/D5E49UJ1fwlQaB8xs
PxyGDOJaead4N3BgIMgw+8xpM6yDB8VcbAKnguUMkJzFlzvt3jkQrVfS1Hrk
Jl6B4UigMVR4JN9wx49uwlksRN7jsz4k1PjDt8AZn8UsDswoo/GI2Hpwhecx
bnshsXlHvgF2qBq5EMoa2fdKvHGvq5nPh1/05VVayP0p78d+jdLak20rHvik
vKa1YKXVdd7TreBv95Ohjo7eKO2/AbgYb9R8+gtDsODJ5Pe12P8apkSWWm2q
HIZk924jzj1Co+yXbWwjxl/93Bu6g4+9DWz01XZqP1BXCzyivxfMvoRd9ABL
N/7XT9YucZnFt0KRfVGMYVd/Hsj4wywLzuT+ppZf5V8Tw2eTjmqv0dOezqjB
05hudPnqVVRgb3UMDNbchz3STe8Lbokdz3H7RcfhRujQeZZt2iTuup+g8iIy
5rXgV62nShfNiN+SeCzGHHscsQEiQc7oIJTBoMwpid3Fs2gPChWOQIQD4b1V
rSYFDpx6eNQOVSVk7F6LbT6yFu3CZBcWzhT0sv6wejT7cp+zR0a+yAkQBc1B
Aa9YW65xoE+9/b7u030e1Nh/CTqlSAz/jeMYD8XgiTdJLTu8lQEKc+KsO/z0
5r2jahbMfiTw+S5UHm+dSSk718D35juGnLxsZp4h+AyoIzytZV1tjEJDdjVM
UvtKbc5uNVUWxAEh0bwlCWOs23HeSXKcekjEYyXosTVqI5QUtmjcTvv5p0+A
R/I5Zkb7Du6tfgJuIHZA7u3kU1wc6lcC+oZMUXAyyE5UPA9fWhfo6Nhj8NcQ
mjfSPJkC0IxFKAvWXdCKHGbgFUHaX+1QfAjQ25kBarDPW2jp/AAUJnJ1YwHH
C0Bp4MpJ+RcEH3nPp+vZqXoojtC3aUKJ3Tb4Q2uU87IKE1L8gKvGUs/0c3XV
OL/hZ+K8wYFhoKp2bCwIpQ4SYNfio87Z1hkLKlW1UN4I48zZe3121yYoIfTY
lMq8iji6ydm2rhtgutpK2xG6OPbvIwNGVU05MCKZAlRSvmByReWNmsjNR9ff
c80PtaxI5DUO3uhXP8o5TJ3h4xJOQz8wc9ubt5h8Ao4ia54KtTeVQvR7O3gB
JxhBOOFCxXMDXBcnzME6GrdLKQUCxQfCv12QKstvSFMmwU7ka5WSEZPWQilk
aHb7SQzLH4D6IfXLG07NfXywGMoyOrI0aDpDWf6v70zg+1xcT/ep3EdUZNaL
B3cCZnEESk1ZwOCLiMS3mH7APO1yXdg5F7e37jAx5UTxzv95JIjUbQUPLd7T
vMrJ0QwgCHaWYay6QWZXLHVq8Gu6ZkX4dbAFbvzEcfkBXCxSep7I+TDy9mTL
puiYvjHO4j2RcSl0a/FBPgO6VLebd7XRlxuWXIC6IutvtBOvmp8dGhGiQ6/y
YJ/eT7uk1T0yoG5x+yZLaUNRPZvq+/ZOiIwxnwrUyH/yhw0vooMGCKMoY+45
GJLJ9Hy6mYktKl/PXbL1sHDqwjDh1K5A8CfeWY+IOY25Ufn8gajsY1ZMf9nM
i9YoFOCLYqW7ZkfprjkbtoHQxASiF1yRcT8GridH//t96SvOt/ZRSfvbPVet
QOch7x0zKTnuqQ6nKxwqRXiOFhO/bAV3K9csw16EIvlmshVk3Zd5ks9iSgCi
s0E4yLSREy82J1FczUlHrvMuXnuNL7qP1Nmr60gN/1lrk5w9dXdezxcJzwAe
nyJw3S1HGfOlaEUNy+JkZIrjXgCTvJfmadRgnG7O//Bkdms88pzvVs1oP6D8
sdjTKY118W2nCR1ReAbudJUflY9Ur+qy2ah68MzDVeaOu/R7x3YtEEWOWT3/
qFf1CQ0uo7pOY+LPXaOe8pLWjY3v1rtZ7Hi2CuKhPKRSXJoDX8uqQqOwg0pX
xhHOUJBZRlrdwYFU9QALbKStXaQ8D3OgQBLQztlXxfsMLh0G9/efeTVzijmJ
Qhk0AI0/5Mel0DPgWHdN2qtKjd09LSi1Zwsvq3CsxutNjCOjqInpt2nSbyJg
MezQ1F3SCPxcFntyUtvH5KCMwaVSbZAFAKrCzU/vlv1RfAPLn6WGdvQTrefM
oDAxjECWuIII1hK1m3kKF81L1om6fDwVPx4j/oNlUXPMroAOBrmm5K9/XDL5
COKVTx6kepKbbphS7L0gam3blMRNGub6VMzhfzUR1YtyCme6VB436EhJQHCH
CIRQSPccDp/5G92wyqF4stsa9VDc6kyK+ywPH+ESY8j5sNZWJe3meorisZCg
cI3j6b45MgWUxqV6ls60PNXlA0Yr0ZhdGC5/z6riivqBcvNf1Wz6gb/dfeiP
l/oRYdpWs3NvlPlqU3nxQ2wzXMI94yJx7+VK3bJetGJ8vmcwm8lcnrYHFmMA
BOCErcLbUwC/G1/gmsGRM5N4loNnpOW0qwRVjF4E/JKiADmbPFrL9BKOw8mt
8YV5qSpRFnPmps3hMekzoTK8kKrhm2vigCue0H+5rZJhPkaI4sbqUr5RK0FL
XvPa48nOZLWm7xxDRDtumgwHlKWajedY/EpSj228cgOvUR318FmP8Qlq0u7A
fSy/hILrJeknZJn/BfK2DW+kdBiFg2YgYATLTqvfu54ykwx+YrIiRzaDxRYr
lMAJ/a6bMX2bjcEHbSIWtBT/CgP9sF8XGzumXRNMnp71QRaYcYobV/yYB5ks
eEnXs8aaJqmEHAMucqYdY+gCgNRrepzRo9TL79e6s4oycmMTTuLACKnHHmnr
ZUZZsvdVyEeO3QM44JGPZ6ONGFTgxuDrj7mLlk84Np3Ukw/b8wXhvdw8V9m0
qQ9pyb7UddOdLmWfK+H2W1KlSAZjHmAIn9QKncnAAcIrMC+w3V8K9D96ApP3
DW5L/MOEXPuJ/QPrStVV3FPYy1rPgZHXJKYneE1aSJjz04B8uvobfQhQxese
UX5fDm53k/u0DV1aqjhe5Wv5qmTd49npVc3/AMD9Mj5TyNLNi2XJE76ftQwo
w601+t+fIuiU2lx7pCkntPG7cTIr8c6tRbXPGuaURDuKHdiNoDK3k8vE5FOQ
Ldf81Q1uLljnY9aw0QhkJ2eaNIhoohxLH5132FIx8dDK/ZNpipkFvH0KyieX
RD+AVwWuwPI//T3u01WK8jbokEmthoKh8o9y7bh02TQXKbhp3o9xo0enLlOh
nlK8HY6gxVDbepqe72+Pp++h+P2vt5W13j9zecJvHj0F3DaAKztTuSPyapl7
r5SEJyEeGMe/s2QuIHBmrxn/MW57vc4ISEq6DUuNclJ/L7u6oGPc2pRI3T8d
L6HdMVf/wKwGJxMwILsnd+C+8dQfiym/Zw9aUnjOLvBKj76UTIxBjIlGg8BK
CT5q1yjd9wqUjoHWlTmavnMOt9NQhWlcdBHnhsrCjy4jPskrzptkzVcwd1m7
I7yw6XhI2KQZa5m72guXAYZR/r3o5F6QJibKswigwPi89VMedtqtTn1p7IVh
5PbDhlHdACoVhjQqTfvKospfzWeGM21rIVglLsgVy0Zr0weAQ7r675NYhOJL
OM5q25ESBZYhXSvCvoMi9mJLdG3kgGZDna5QaThg9HM3WWqPZeMojaHCvDxe
mR0nTdi8GZt2XHJ1OaeGBadq/kLbxU5N2JNL9DvGMTXrViOl4thm67OoRJYN
rFehElcbDTAfqJ8FN6KNj9/g9OCBiP++7YwgMbRcqp/cspZzt33WsOiME0PT
YpeHVIahy2XjAK965YglFbudRFR0L7QRc9s2P9D1ODJBodZAmeG5i1XIdpSD
GmayMnQsOTyaIFhID0XIBdBY5okll+mSrS1TF126TqmxhkeVE1L0rBWWdovx
X+XDg7Fs5yyHGeiFJe1BWC/w4aXRgO1nMNW/lZFBfhIeZdphTL+7ALW2cQL6
LDV7hKdn5+MDIq1hXPEvWrOAA3QcWIQPKjnTtZEyOXi6Zb5ai3QhdIzkkarL
C9XhqUo/MiXNb8VfStimsr/lKDp89D934aMEUe0hlibfwDUT/5Y4eN9u1mNV
alDZSCUtuEfhv3OFwI5HJSHH3d4ArOVeNR3w0YAFjTxBHJkP4Tn3ZhmUi6vk
+JB4HC1ZTPeSHIRT62hG6b7xWiDarA2NQEOBFv07Br3rPkkM1MDdx77aYdqA
g7yXtY1wpXflKvCRFm8Qns0KEshaFP/tgBGigEArlHuAYlciXNjX61Tmnu+V
pdM5XXZEtQ9x9zOm3O3zmacQ6PMcXYmvZ9J23At3G6IlyCOl1GR/lERjRbht
/LPYhJ2OpvZ9jUvzydVVgNPma1E/ubX8SMPgsNdieZvst9MTZ/LNOnOtiMRL
ASH5lcM7RYMdCEuaCqNGzKDvRj351LTcFU6rU0XJHrB5pnDdEORsj+x2XVW0
CSLfhHgGkGspmw1iUjIEc1mLLzJwWcoI+0zViBMNpoVw+s3wmoPvo0tGIQrR
Q7xA4UpXhWM5qvfI/ncZKF72cDgWlqeqFLebA880fgMO9dZDPmsXMbUf26Td
HmDShVz/iMhLycbyypNONL6j1CSaYXjxQv7WsMq8G5+tNngpHFLD5QB/euyA
j0m4FTvqGvR+TbZoUf782oJhJUrNmUsbAjtKfeK5xa8CKITGn5B7GyVuIlDg
R592oZ/vZSPeqpqlQzliIxiEnCs92N2IN14FykrFjVfEnY3y2nU8ETyWFBpP
FgVws9ziIi8w006InBOVTxix/gDZUxeMMx/JxCdtkcU9qW041sXdX4n3EKfC
kbMTr5dk/1AR+k2R3ZxQHm/8Ol+cwUtGj9HEKbKVFu1C808wvzx+nHxDVBwe
tzS8dWnGH0YrnLaOctU+j/Jm1JEXn9FTBb5wfuIq7knWkaQ8cVbAPSb8mZ+n
B7yEwX0kTwVEClE7K86nTIxrqP3fEfWyCrFr8Gcmza6xA9Q+MscEdfL6QxkY
oG28HKp7qcg5HJdOji4TkPE4sqDNNcMn5RtQ0W3ruL7yWYUxIea0Jia8AitQ
9Qr+lTj9zmz3hBXib6PguocIZUbmU8mgqhtVXDkwNkH0BOrxomsSNjxscJTA
9tBq2N1JGgzVJVCnpBosT8S9rbOqBdZ43QGqkZvPEXKWUjvY/RLHnGSomtP9
qt9wxNrUzS1Fi1B4zkztfh8MJqAnR06MxyIQNbUakLwWnNUJTbs/FXuX0woY
+4UMRrggKOrKui0N3bCtpTzdP8MYbzCKS8ncxqfD69P/0VXTnCDp3CoExRkH
fTk4dNI2dUW50M2ssHqvdofCv20E84ssRS/Xpl5UWx1GUzAREobX/UZSHW2t
WbB73a8L4oQ2IWpFE2MdQ/FdLtGBJNXoPNW9cv4AVqt8Sxy/p6BCcsbYDvYC
lCJlAJEnRmVGK0yGDXlAwdZoWdN3EeA4FtKA6T0vrMknu15vP3LzAmmmjmwF
z0b24mE9Kg4kQ0V7Djx9JfcYaBzF+RwK+guDmcxnu/OwqKGGdz7PPXYOW5JT
RN7h9GKeTX5giy1h5xbvecS7nLB/WW2dQbikJOVOzlF+Ydv3yIRUbGO+LVSr
JUb4z1CgVzsH34kiBh7obx0Vh7VnYf6mVR4ac4BcnyOa3vLdxjHMAyD7/0B9
owlx6AofQEM76459z7/Eb1A8r0fRaomd1g5S87L47C4Z94Azyl63VZZQu1AG
v1A3UukFakVdW2kCHY5Pz8TzT1AbVo2+6FaEpzxc1H55dIbmOeiT5NjOVagb
FH9kZMkJIw/PayruorIjMKr2ImdEFuyqAFFaFVjhrGKTHxg/sjw3PDdpqD1K
kmoNcpJzY9YhSJvGwIEKlXr1pTdoBMT12cCQDhPiwImx89trZQ4BrxQFUo0a
MgsDTPCPihUb6DAIM/g9Vf1Wl6NNQ3igtk1l728lzxWw9iKKHrOS2yHohMbT
S5hGW+ol2rdpJJArlce+z+r7yyKtyPO7sivFm/koNsRDzFAv03wLp7fhU1kk
3i1rytrvAwlcTSo9oWlR8mN0iLpm/Ui7D3nIhctR5uPvkvTJjrMD2lesQq5G
b4rFjYnbW67mrpzPJox7+MbBgCeSvf58Wxlb5b+g3Ngwh6uYa5nG+If+J4k/
K5gI1HAZ0U2AjAc3Zj5Ki78RyO0Hd4R5DJRJ88DcVC2y7t5SgCMm/yD9Yv+9
YKA9+OcK8KGK0STtJrFQKDeqskAx1V6/6qQ+SV9qXShT929d39ZDvm+nZ/Xy
SOTniAusDLITfWifK1+XdH2LJuAtNNsUmdNXQawlwEuyNt0OZ5GY/anl8v6S
vZQaumBWAMzre23Wkkj8wFWZ2Erqogy6A/mPsIAn6zLHGOgnEZ3PnvSqL8/R
etpG10TGnzPY1GQi6ghJVyQMplbZI18TtHNxzbY2wFfPe7rzKpvr/g12i8Lv
QMG/E7wRaWhWbcq0j/u2UczK6fdV69ZF8n7+aRI8RqGQAWGz4tCVPD2TQSFx
PCFETGb8V6kDGkcxYdy7YnrOX/5SZBZbh5XxxGF8x3cSvCeafzMEnj46HwOa
uwIStwaKP/oqVG5yr/XIrdSMBYhjSu5KduczTbP+ShMeKlysMBvii15KxLM0
IOebXk2SFQj6Tiss6mFv6ZnL5zftw4Za+y9QA9CMZRBDcUWztRBUZTm0YJb/
ZZagbIwdUDi1R1hna3yO+TBgPBzbIaj96lmcMxQXkK42ZOR8SLynN5MHwIIb
g25wGCySQYNISZL+iFm8M13wXI4HYlUcNs9h/l8F6ysdt0qOvffeueQOvPA1
ioYV8gOQNmi8j89MIBPSq3j2ok39CIw51xmOoQNIebkEaQov51db0mJvnb0D
NzqRiz8YyVVx5hBybWIQaRyf/Cs0nek2pcMwKIHA2hREN9jTPXOPR+8HjgmZ
vuLfs6eUDRkORId0XFBR+lFdzfnEYAv20YSmAPjYHqHSp2D/AixQPJ9odSly
LXNjP9d7r7E157/vpNYllgap10FBaRvNYx5WkmXcm07vUtNEhviFHdc0Wg8F
omWIFVqOpvxo4ZDixteFIXHmsyLO7LS05EXrtZIWJM1aw6W5H3KyALqmEbnY
y9dAoHHCb3QCnhbsOG3vKJ+6FMhlOWNkCUjKPzmEkeSw7+4tux8dO2LuTolD
8VlUzEGBWTLB7yWkdMPNI7FZwmKdvFhgzSJjr66wl/ZK6KMo7AD/BZnaCu0Q
XRbSwYF9tDwY+YcanNzH/leCl6Fn2xGupYFPvN8wHygKd3GXD6DVqCrBL+wX
axDZwzNRxQ6cuIW46IjQCZYPVz6I7zUhSuHPxGjmFhpOT9ISojk0x70A3i7s
unS6VPORY7gMgh6NR8qreMPYMEOvjaLKtTkc0WqX0enioq42064Y3OWxWeDL
8rZ6VgQeHCYHJO3SuSNLq6LXFF7wimlIaGUYqLl3ZjmgjweBhK9cDPicwA+X
LIRNqdUnCIBdo/meYOk1tXGHejt2zw6aTFrgJwwbuItfMMO7T0PU/BddpHFF
nczE75jQTVzYuL5xTuWlMJA1VU7oYbQj/AgkD3eet+EUikm+JWuflR/NWFvN
GioMzb2hgKgRASoWitl5AR3CY1AbYgXHpABeS3Uedo2QWqlVLCrAcgWnk7pr
i2fi/cZl3h2IUWskTqPPWKss9lMQ3GToFrAtzJmq7Jrpd/HchTXEC2/PYVKb
6NkT2ryjqaA8D5Njsypa0Y62zoqzdhSnHYn0MP9TIx0svI+WENanKdIa0T1Z
NGl+KQZqPklF0UFezWpIcerZm0CKpMlmVu/9EsozTadfCGAQ727Se/BrLNpq
/OTMC5p/oygn07iuZM7SD4G6zsAAc5PVPGELm0U0bVePCxkMj0tzhOSPSmGM
C2l+S6YXahN28jGydhHpn6P9qGwt9skdtA4+/rsP71+ubzpen6dWIXsPsvqD
rCOYxz3rkDEvgX35TnRJ/GjlhqZlWSs6Ui23ZiamHhXUCEZ/9zPR+iMt3zM/
xIDpsISVAaaMl1sSXERnxdvj3gllhY3OL9n091uXBf3XGlH+86utYCdo3XJU
oEgQS4ZPpFsqvq7od3vxVOVJGrRF5zvAfEEkbs5QBYzYsldzDhOUl3PBGeVp
e6QE5l7AflIpkQpdKm4FnA2QDYZZWfG+3QkNr+FoYqFX2K3rSbWER6kcbev6
dPU1URQjL/BtWUpvALcUeVSutxbwnZx+3tICNv30JTvsJWtxhcXlJqrPQugs
OaJQiTFg5jMaQTsVPQtPhFZ1kdz64xC/iA/mNnkhh99SP9WHP0yQqcgX0YNq
d38NosdBEiEATNumlwQxGWL+ih7+MMDGjoxv3Kv0Ao+oD1JQQAhumz123ZzV
na6OzzSwOGwowg+XM7ypySg5yQXleSLDsSLX0cuHz61wWqohXghMnYPhsK2W
q3aUwrLiHM2JnRVtlMt660284R1lZpktTIVIj5/k/8YS73fF+9Py49JOm+ps
4GaWW2HFuXBdLrnbRQGjZp9LBhIg2zk8XtC7DYHz5pOo3HQkIcvBskIiKahl
+0Yj48XXwaMbcFN3gkrtagwBnWvr9y9eJgpVp8UcZflq2eXrho5mTsI+2gHo
rzRfIn/0cuyOSQjoGQTM3k2BVf/U7+4VPfgVvZ9oZctybCrKPj1fu/mHnxnV
ygkViGLQZ4S8+RY454yWaYwIpA8YaDIaVHSY2y3RBMCLSnou8XhZItrKTeBJ
o+xLSTY4a3BNI0NPiFofVYwGyiWtDUoO2F5+MyxIehidksY1HG4fCaPLcoXX
6iKR+89fHdNItDDnaoH8epAjEIo4dWeeca0d0p7MfJHlnPnKNIg/6rUBzuVB
knnZfXNzmcyvISp+kUmgLC7eEMkXYpPauh1emiJkEPjLraSChLCfJ4tBlHzl
roSQXPEe4bcLHmbGxjmw56aOuTSedEKlcwWKx7Ba3c5V7ZGIW+MyIA2/wCIY
cU3ohZlnVsSIIWectpJcgNsiFkBuuKFO233fR9Sunylf6xL5KXOqW1TaYFkj
qmCTlRaOSLLSxYmg09k4wV/3BcbCq71GE4wXtqOakI5SVaw4RLpDyZTMCypV
xh4K6ESDGVBEVPLVaadvUQe0frOu8A3gRA38PpDWLKXfSI5zgg5xW9j8T+6T
qlwIbzd4pQc9eKPXoNYk2jCQ0YlMi52enEMDbkexfXHIHO+3i/2zPcT1iAAW
qfNSleMGQEmK/3IX7CE/uCR9brRbmLmS2J72dkuW8LwZgE1/ufL/A3PpoGcn
+Ce+yOrwfYXf0CRPb++aO2+A7w3tRWnIvDwnufgQz6eCWJpqb5tW0ymzTxjM
7Jdc32clZOU31xySctOgXZkXdjK0azxJfSKEnUxQnSlbxPAWDKPaqTO46MmK
tvK/qdH9JkdHkmKKCYl5k9+BD9aMuIaXX7UUU+QECFUZEcaK4fVZ6T6lJ/ID
vQJ8fUk1LfOJA11z9l8bofnm6bEEEIcj0rir62R2Uu15WsqdFg5UFYC3ufc6
iQgcV2R+leLtT52by8OE5+XaEN94EAclXuJa8562TU7tJD4RN4Rg7btufRa6
ULN33pVYn9QLaMeZlyU7Lhak/1Hw7Bx0efFmkogAB7nnHRmMYx5OwMxvfMZp
PTDKim463X1RtxQCZM03TsIEfD1Wi1oB8yvNOnmmMApweTNtrjEB1Dy+XygQ
ta7jSUJMHTL0QuyZVyW+rAkyAKF64NXtkVrTtcJlqxLfi+MuPbtApkMmDHlG
stCQbaQ9uuivTOhCzHeXczV4bJW+RPg2ToTZAIXgYUosNBIpat8LM/cad93d
2YV1Yv8R2XCdlWINOWYVZG1rYxiOF2xUiCJ/vo39OjJC5nLYCd2CHQ74o3Y8
WdQtfqFPIwP0QIujSXw5lSvipXpmby+9RmutVtIm6pcgdUy3q+InMaYHeo/B
Z+4Ob/ALdYByDu3uh0jhLR7Sg19kofOkvR+c9ZiAD43qhm9HmR4jfWtp8WTc
/IWziEJwV3TgxMyRUCDSkL0MFX4D+slbvhuDy/LL6GezV/GkhKFs2rW9Gz1o
zTRadfBU7b/zxB95vxRsscBtS3vHhYyVWduyNl8Is1adpXavfMis9arFmuLz
ZvigaKUAbmR9xP15BOFHv92YX/VFfQoUuE/aswxczVyHKFLg4mz1wb4C/AHM
fZCXF/TNOQ3pl/OTsbKka5Az7rUHW+NsEKf2Nq9MFvxlG+sKsS445pNNNxkg
NMQe0MUQBcbrUU6EtT1ziHH/mn0OWnud2QPQ586uxJFUalzZirlRgVB9PM3k
r5YXZUPcuhuYgrIWjWSrqxQg6eFzeZOx77RFy2ag0adh8ldOCblicl6FXnQr
FcNDUjBholXrjxuZfCsTrW1JWi71TyCTy2jIjYsGXYFj1d3Ho7lXkxPcc13Q
FDdKL4ML4GUbBAx5O9F5qU8gShZQ8SGx84eTuMsdoKGrGVaRykAxetayy/ce
ZhDPWws33qE5d/VxvYViDix17tuzCdami4ecTeU9pXCV2ZIQYTaVK67mKY8y
hM/VtHS/61boYNxviYve7d32ZBc8JQSQGjfkxsI3LBEuYn0aCW11UCTKERv2
/vRSb468xXDP43/81bmoF5FVV26TmZArGYa6dO2q3VCc0HKjm+6qbKs8b115
mbjMh5K+iGEnpCuDn6LdXKVvPqvqOiQt4Axen0U+MVLONhV4Is9GSndUtvWC
f02dBn1+Eye4xz8NYjE83gLsTSTA7AZRMVNRUbHj5ruqZoqn0McDinqHUHmP
c+HnThdARFzEFh/LWsoot3bFlHWddynWCu+U0A2jRN5lFQQ966V0rq3UjnCI
/wt71n+W2oLltT0UaFPhHWa8x55U7lpcQZ2ClvwsV4toPwEhPr4WhZO2dheV
7LG99mbUiJaH/1y8wGyS/wg5casgOc4VX9F8ffSy0ngRZ1hY7PuwUtgFXh+Y
zUZ1nbteDtJoQHasK4+7fLcF9zAzCv8BLRiClA7dLPV2tw+TkrTFQRT7Y/c0
ArNknbfecywN+v6KWRmu2QSFc+O+DanoeiQK4jjkSXtUckZ2RDC6N0pf2/Cw
L5msSKcWSGY0sFsrRY3Wji0GlQunRRyLDIOsfqcnvND01wKpeDr0hqoMgnuT
R9ICHaa0/i51kTWw0IU8veBeNoVZD8/JgtYh1AiKBI4Vb8clBF+xb72XiTfR
D0WkaB8G5eCb2NuD82CBIaeii41Q57vcWnc3QedX4fCQMdTBuRKAJ8vE+4o0
95zRLzWZDDEG05UpVyhsftoFtJhlTYq+INYcDgibSHy+kIic1pc6c3ia9UnF
tTRjwi6BjsZ7d0PPec3N7GLmNyRHYY5d24IPjFKkBA/dg03SlUSeqIhsDKQe
hJ8vtXxE8rPS9OFyt0SFAGyuapiqSZSbkAP+LjieB+bfbfBDT6ank2npGJ95
+GGa485ASTfPMmADsJjRxhaGtfEyVCJySztJ1j2V1dEHmhSk5dt4UIj40p/D
SHlJ/Up5l9HCGZZbPeIRC6RcCRizWHO5UkWjNBI5N0sBCOkjmtL7i2V1fd3i
5YOYMNH3KAfUmwscXBM0gnBzpO1lvsU2MX7VST9pm7vAHAY5Vf1f1hi6YTAz
K9j/NaLzs38bA3adQJOHkm1rvfRVCwIFyu24sgpL2PMjoxI49C1E0gdP5xUl
zsoIYr21RsAae8FeHRUfML4xlLutpWIa5PwpADVFRYpiI08n4wRzElvQ8QKJ
mKUx85eGxClCvcXgxG7cpiKMbgY03pPE8vAfU2OVKzFxpEPCQ9CUUJnnll5S
u+gtP+HG1c+b4HMg6cfUiaEM9gw6PfFjRSzclxppFuofjFZSBgP9xfIvsSco
iol+OTmkTAI6vWVkWiYP9kHztLLXqogze7lFyslHBCL4xCe5KFDOTzwD0Fvi
E6IUzMN5dciO5jxZZQdQZ6VinJdCUGuJsZdBvKYFvEoyIBSxZGgacqx5B2U2
17/Fp1DBZo8FqsrBIOqwkksZrvoN/jQVlxvBCzEzM4BKJFRrhQrYKatz3JI8
tRx3cYeDDvj89mBiH4RToIrEIzbn2fI2xaoPAvprSSrhYCQ7TB17JZ8lt16O
ji0eGTwT+SKUwb2/hPK+5wtkfIodyISAxf9dp4OqcaIZLI23q2TcLVOZ9mCM
LOXwimfHnquLvVBunltyga1UPFBjE3Jzl612I/3tMUtJMfDAp4z4HNpZHFJ6
P0GreUXcED00Tlm9nBhHhzoYr2Evlg0wQxc83po02QlOXTrciA0OJXaK1LVY
MD6dH1yjM4OqWLh1YeYYB5Q+MyrJHPWGs6ZJrvcEyk8oBtA5Y/+2bLomAp8i
hC9YO405I4DUT4RAAq5La/kPmsg6lYJTy9r4n8FgT4Ccmq7lwDRCnfLjYRGs
cjJqrs5K7dyuNIjebHJI+AwsAEpQCUV0Awi7uKUzKsko1OXJc9CMvzQ6lgxH
VyRMYpLc7e1PRn4ne6+eHTfpCR2x1ZFGT3Ac3bo1QSw2Dd0K7dHNf2VYn83+
YyMZHhoVPRQrnZ59u7ZmF8Bsp5lVkEn6eiNlfktdz3+iPB+ILACgsoPz8OqN
wEiC5NoHoqQ3wiO3vRwVc6umZ8aA3ZnznX2IrhDtKMFZ5pJfvqlauVvwtNJF
xJ1bp++L2sWf309/0CQFX4mjFjv0mXm8eWnT40R1XA7eKcC7xwZDATDFCg6i
y5qUuvU/OxS3b8VQpRs6wifyhJ7tQBS++BOFR6ul/pB4+RPCKvBi2ncbSM7W
T9noweP4o9SmD6NcbEtdU8n7hYlNKkXd9dVC4EGPaGEYyxqEPCIp7rrczkkh
xAwGy2Ziw9BcTb8OhJMznIZputNlGTLoGG4gKZUeVAtQAhGLA5l7ZCHRtHT2
lFSU9g0fIVvEVDGloAQ61PVjmFvaBgRwlMiSBNJC0n89hCP57EdsixBpGMZV
dGOetwfLheng0JU+sw4T/uuGTWvVuGQI2s//kklGH7xObK7eag2jwibNoDmk
ztsoBYnvU9miCT69Vkt0peinTLF1Wh1KB66oI+5bbdOpq2pc9RPErPfKNWto
cFGRAYjhOVBKLClmMN2OkIR3VoDnWnojLdArO3KeVOazfEgkif5lAQTCjJnv
LcpQ7aLNRPO9GUeFoXiRyBYTD0sW746Pd+O3vu4zgeunEl29WqqQndp8gdo7
YXEp+hd3Uw5hNB3ZS9n5E71TZrvtsY0kme/Ujdv6cuIsq38vhoYdtdazH2y5
A0ANp8leMloLylBVU+1StwFOsDGWVnlgB8xLYWLgMSQo0uCvhUNIEES8RB7q
N3QClfJOMcPFok4eLEBWoUSG1eboZOhni89XneRm4Y2s51XhnGnEznpf3pxA
kRzm0zDnuGbJMb4ydEybGp0LBryqSj8O3yfivxSDohWawpcxDTYrd5Z6uXeD
zi0IrLAmGQNfTITqLXPPHT4M1QkAyorVteEpOY4vsZ+u81VQlUuKOkm3SgUT
Mk0WrZGO6RV3TuuDB+BRqZwNUSfEcpCH7ea37ZyY/365Xc4yfOs3+UXgH+rs
wKmqycZXbtVgFCX/npXriL5CAKR8Bv2PCIz9gVN9Qi+mhRzeg6k1fIm35rI/
npb5P6Ew5R1n2GjCUJbGS8YQAQkt0GX5iiZMdVWE1EmQBxiEX2H9/I62fKWb
M3BKH0aSUL4Uy00oVD6RyD+6eMppZ92vDjpjOruBPhjb2U6zDYk/Bb4d1LlV
6DzSO/Zu4zPZm+WhyYpnWU0TrUvr31AYBj3NjEJM8v5eqqpJsoKyChGzt0m2
DJeTeMahhLL7cO1vGp4B6tqMQoAadyzLj0QkGUqaXmhgEDqYUvPzoLKEFxee
1Ng44xmwq4CQbXYiXh4Bx/V5pF4dnYPHMMpl5jfn2uRIPnI31lIH5RJFhg35
axNhQILRWQfKmyhvekeV5cxNQf8lqd7IfHF71tmjTb1u71m3nN4RMdgDwVa0
xUy+7D5/qh52IWn+oMSckqIQPdIJ7rR0lDSsIIRwVqbOPRCPW73AZr3hcKO0
Gw5kJJTNhu0vfX8nH5nVHGTMU7VPz6UergVwrLxc0aa0ixsT5WJ/fgCovaqa
SaVq6DdEdHQSBr9hMf30wQl+Pjb7BfQmSNr//kCXQw8Ne/+Hdb7uX59iWqxR
oZLBZd7HqvVfOCeg9fryw64FUn328p7OmgPFW/6Ue/uDQUwV+lR6VO85FF/2
gaoJAjQ1NAAFtZGYXh9kjMKZV6DTPFMcQXvD7IlfdNcGMt91R2o90gz9aTVs
kZBYsfTLhcgZuIWMeVVQ0ArbExhdgAgiBOdr6fcAuJohJEjZwvYaMh9I0MiV
MW5Tp/n6RXf/+YLgkcguNiBV+YAtn4isywx3IRBpeMTOs++CupQZ+pS6PBZF
NDLjJ0C+FG+Bh8Mz9oi8ondBxmjVjIGSGIjVU3NRblm4vEQP/+gFjdQZmNGf
S/ajHtdfN7ugLoZO2tRDt366oG4XSS6KNs7xB2aB12pNMeD9x2o4aAxSCCZV
CKOm3WDrtdpYb1sp+ocyZ4DyfvTLro7u/eVc+xdql6aTSzTgS4t/zG63jTQl
Ybq8UqTRmQaoXe3+R0tjzwBZHnRwht50MUtPgMJFPbCtf6mAcOpbEoBPCTGL
8FSkR17HGiiMoPwGzL+IEd8CWbRiRXaRoC/UbrN9JNr2Lla0YI1w0PFNn/4v
wP/YgoC74UVu6j1/wFpFRmzMReLMX0G4hYiGhoY7kg9xtZNMy6BRZTR48REk
8ZeoiUvbkSc49S/X9+cOc+/Mt1I0FrWnftWjJuchRM0oAJinlXKZKe77nDIs
uW7q3hU2Sr8BFwYu3W/7RYu0wP5yzg8xd+rej/jIt/JInQjYVLqV+FemPmF1
OW/55pIjzGnQrRO3TH2lBEgLRqbMeRzASMgN8eQctQ44zZGpKceCusGO718v
jyesvhci+SmHAgCpp7H/+DpTnGJR2zFSSFt1P9Jy2LXIEboZl4URjg54o0ZD
iXrJmt9iVqboT6OKj7ximzfgsc46jIB7Ha3gK2kKemvfmQCE4EsXHrToWViq
fne6qt8AtJKHTMZXwV9VKx0Kw9kzu5uDpdJPCi0uzCgvJ/ZyTfe/iG0h06cz
0rVvApLdz2KuGYHwDvUe0Eg+8h0L3/q08p8QyUve/Z8yT35PUExP7cnOW2RD
ds/Sg/68Ak78XU6KusR9SUKbi6acFhtAaRSuZ6ECXz9c6n3U6alEbNLqc25K
BeJmxRQ9+bTUH4g+5Vp/7wZJAo8QqxIfGvqlcK9NMNg2OAub77CE8iPJfP5S
gWldUbl6xpzp4gP0NA+yPjrG1RKMfqNtJsK4OABt495p0WHQ+OufWFJiJmyc
ZfhQ8fx/ftx8nFJ9r3QSFjrBY6KfhQGFzumREldcm1X3OE60gftWsiPK4KbU
Y+ZVKkrcXM87nrn55Vgbi2hgVLSD2J/tEmGEAuC8XPocCOlXR6VMekUwLEqC
Z6LBfLj27VSynYUk3WG3ihsDW6Aw9qsz4vl00MalkaeGK8GrkaI6La1OdxBH
PzNDoYwOINOaogVLpCvO87NR1mkjP+Z1L5wPr1DWoyLxUuvPiAU+zOwif6NQ
gmwSvMykymFXRA0RkmLVOx7VqmnITtPEtxR0y5B9PSTfVSRtTuShLyPuJ2sc
vqPRJHgVkQIpd4WaICeUMpFBV0u7AaWWtddg+eIUj6iaU2lMwmQ2p1AOuvfy
qbhCLHvq+qEf2FzyfFGBe9qe5pOdC2AN+i2mv/9WaZkX+BJnmyAB4lD9ieYl
7RCS2eEk7Nr07zjj5y4UlQzMos1E0ViNtf07GeI535VgemO5xlkO1IemsU2y
JiG3i8cpiBokT3ZCQLuqZBJMMPYJL/NBsKAx+ri2kF10hLen8Bu/kR+ndrs+
c0JzHe7/AO52XJpeIeYOXxGJXt/56rtEZmSPvwoljlVKYfKo2qsxlzAdt/xU
/ZO3hb36XAqEWaa6bcs5wVa5wzuOcNyH9holv5If0qv8MCCKhBPGwxvMDpml
tgNiVeppKXAgQsoJteTMpQwYp+HGZXPYeR93lZppYAKYLVtZMzbnpHlG/dbx
+GEwclDBv/LzFeYSlvHLJy60Al38vU1HuGsWs7yUyBzLNSOSxQwDT+UZLUgm
xbiZk+ZeRD/Ng6wec78rkchzYzQeUVZNyoadPnGKdVDpeYM/cHZGFVwRJwMg
ZzcRNKohWyp42fFKNjM0VfA8Im/b/fiOXA/7ofugeYQXN3tfTPcTkr1kehM8
v3GEuEVAVZO2bqx1ApqlPWdWhcADkp4YtTauB6mTYyILPUl64kpGSMsBtn7n
Vl80ha9ZmIMtKHakV7CpZAfJZp59tYkm5ysOcLBabxmoG1/ZJ25ffi/5uBYw
nGZVcSYUOqP25xwXJbPi3eSyH+oEN9lqSNSM8LYS2zi9XckBupnkzYeGl3j8
W0oLoJESlx3U+7JhPt23bYbwIFCHIcQGHS/OazHLjg14RLIaKJYI2XAuV1xj
X73UAPEI0rGkzVy2tFPv+kR+ibHrcCRxElT3SXTJO7mM7wAtNUPahx8onOEo
41ZwGhFofrhza7Iii4uHFxHcri+i49XtYOt/ZwEdX2VC7qC9gTumeussSt9k
ttqikLDud3kLQLdWtU6g51IborSfItZ6LOCQ4xNBgsQ0fl8fjJvdlNSZ15U3
/h3zyIcsEybHxng8d4c9a01rmgRj+F9XfP9VY3KJnvKAvXaDtnFktjTUMFjC
LzNzq2yYydWM+VBlXKDUnUXdARK8/0tUcU2IQDVgq0nHmdv/QacqZlCDwvYW
gr+fyqmAep9wYxBoaoAHq6MCBKOyWS7qlbGk4nCRhfLTRz1CH+lu9/LgyEQx
swFI4T1Wh7B8vgTL4R740K+es7JtxvIQKeuBEB0P+geyHyPfLmZKLBmm3cIC
AxluO7zdKahpoYq4skSLJGl9HU8qJS9hfsqUl2D+KiGrDS+08hxlMPEwymg7
MSaXbLYGYbrnKCid7xr5KcX0YjwuScjHaW6ErmIrUzrLLkI2+SF4+fyY2wSk
1utrfkUaRLRtv4IHSIbXXj03uTrkKmfiHyolISDXU+h4GHogXQ4CciXqzGOa
YIirKf1aFbiy0N6BVg0D0C9FXPmmjVjNR6gXWdccyEi7FzriIUmxldwN4jt0
ElKL2Ym9rHxVS2DcMkXSyzTn+lvVd6hBHxEIE/fwYct8XuToPXxkj+NWOJrJ
f4cFYI77hsXn9JQalOq0ZK+jaYt5MqgvURSEgLVp3Ll5iOV4jMPNggECib8o
JoxTrxrRT75WUiL9Kz6ss3PbqNZcpzW9krJRXn//He8cdWlcijQI2vmVH7b4
iq1kCtlEBtv/21YLmpuqJ8j1NUSu2FQ9YHzCJhC4DOBEN/MD9Gqxq3fbDPcp
5qRBhs0LjNmNwfFbnAW+h887oLyLIn9aCxHRENDeKtckln/Kt+tzl5nMPyN1
H+2LIzWxJ2FZ4KOgC+HsHuepmyuYhXs2EE1O6jtU617CCEzn9IKwQFOWRDCz
tlDPRiMXnksQ4oBVuWcKlV5PutUlbdNRSdgT01Auq3/3sxl3jGEGqv3mrCAK
QZ1ml4mKx6WLFfExuTE9yvdWYmqIC4BacgnCS5Fewgp0hURwEvJVPKWu3Aof
zJeOrOH9vRJPqnASUF9QTZl2xk3Is0lBxNLLUhRIrCMGndFwZoVwVhlUrYP1
0ECRMWEzHpwGsDvJGwvc7xqeCow5i+rl4uyQtDZUw8VuyB2X4emDPPgVFdZp
DIsqzFf3S6t0lR7pqCRMrVS6kSIpKYht3eaaBU7J3x3n3bcPs2WXdv8zAb1m
s2vo5OaALA9EXyRxfNS9cfYf3CKB1w0U38CTq6WXWG8y2BAtsEIojosNJ02d
0w/GAtlmuWKTw/LbBQjaxeg7CpkUxpXNcJfUJpZr+MiWm35hwDAABF88hMhw
kackHAuAlkEFN+UXuJgprVY9DyG3Q3TJeLbz94bOAiukNrQL6B3ojQ6y1R83
WB8rNgJwWg9np74cmQiaOg7vwJVYsQQjxBjshTR6FF0g1q51w05FVJwDuP3L
YBclVeVe1YHp8P+HLz2qnUqk88OWB+Gx21I9/BnWlQGE660CEyCVI2YNJDo8
WvSv0p9k1wPivUesb+LOaH4JY4YdRGREDXA6hIUInLTz0x7twn4UDNv/eEOT
5XHj0bcEPmIVGTCksJDhwtTMY15EeULlpxWnthRzfD9s04o7ynGt0usnpKZN
+OOG9Yrwed3ti2ZNewqNYHlAtSpmmdmProMFQG0MMCNmqFrIZi03cyZmIqmA
Xszu69WCxv/HA7blirmVjH71R9/oHL93NyWfV2FTl39e58DQwLcfPddA84G6
K34gB8N65r7cqPQ8lCPbMGwHDMUHjmC5Y6hzTVm377wN1yHMXWXu3iA9rhvR
avyw6qr0RR3f5wH0XNq/KHikf40pen+RvdvJ1rSJres8ecojao4lE6yiRi8+
tjS8iI1reyMr7gBIi2LLCgbaEooz67xdT2B773y8+5AGvf0uBrT9fMNzS7V8
soMXab6ucTpaU2DP4g+q6mWCkq8Ir8EWfN1IlWk7+IfVg0+U7AdFvhE5vyZB
sZ/YkvVsZ7RTnDTvT7USGb09c8W4v/qr9LgmgXkm7Y52bifRHqeukVBPniPM
SdB0bMyG5ZFgi0fRnPUDTYpP6ISJFL4zrAwoca8GAvA5p0i7twNGDmuNoKnA
FKzHlGLrMzS+avspY7caSNAP6qgzsB5M8wDekqjH7N3DHub7Ah5sQ54pZiVs
niUqbYmgk6bWk4FEf37CDKz7n1eB/alc6A9GSDotDvhD9+eQYvLjZ8UsOTLa
xAlZRm1LmK96fORmWoc3EXyiwS7GGAu0m8O0wJwLal/8+AFseD/EpeHOVdDf
41qN0/iPeFkEyoEWqHlT/q+51fVGe6wcDLgbYsto/WQQUqF2wAu2dSeFTpcQ
CjpRqkRiROK56nm1wHMYnElPdqvv3FssQqqxU1ABzo/GRd6lPnTJywfL+fIo
8BO4ha99DDckDdKeUnL2cQy0cPORC5EFP7fk6sVbfrunxe4EIK/gvsdahm/f
LY0eVsp2oLqSWQFeuL8Vtvc7+UPuDFw/s8K7FuGGsXqqRfVGpyDDSnz5d6J9
c/SqDu5eVa+GD+jEctgW90BzFF2akv/NlRQ5SSZyxVlHfMIKL05kHtnl9phC
lQ4RaAK92kbd3whgEUDq6XJ4j7vD2U86HXNcjtchKrNTkVkvcNP8Z1IAgM+/
8bbZ+pbqeHVI+LDy83idhKViC1VdDoG0gCU6Ik+HKy2yunhHYWUTXuIL5HzH
XPGVnPtZZN96fK3qtTGYC82lXPdNUGnG9CYnYuo04HphLYpBd4pATwvZfu9V
/80Iip9APOGKn9k6FvhcWrhNA7qK+0bnLhFg4aZoPXx+RVVJLLfyzP09X9+u
4kDvVX538LJm6Ykv0lslhmOBw5s6Y4Cs8zR7aDwTAlO6ilJH/v2oI4/Zvswy
eLy+R6Cqk1JeXcfMUI3aNZhMyoQZEH1Ya4S4s5+i2iYhopDi7EvVhCEK1LH9
yVYgsRRFiA3J4VlE43PxZ32qOdHGlkxDDc67s8oQQlWmMera22oYWM2YzoNV
j7JP3S/NtayOzANMT5jHIwCnzKY0+y/40m19DT5hLVBcH2hwwoicXHcpmpi9
YfDU4DrrIyUXAEImQeQQ4aVTPWcYYTRdhefljzWXRhwjFHgeetHy+RCTya8a
XZJ6cW4SMDJAZoe5TD5K1QSBNVAXvGmEfp3RHAoykXS7NJ+Z0QQJ14LS+/1C
dScZOnm+Zt4tTEZgL0GFxgx95OiVfZyOk0ov/hBZsr68Vb6FbnaR9Ceyspm+
H1OSJyyeBl7k+4+fIUS0PanZQLIi76A6zNPagjC0AFdclm24d220aJuUFvrN
BqyZ9SbsrQ0tevEvE7Wx/7QDg+ROicGM9ZYw9FP/nBY1UKCzaR5J3GYFGLuE
VDJY+ievYdkmEkyc+9T5Q/vgJNlBHCBnq19Fv1q9REKEfBikTCYcRk3dI7e1
Lmtj2B6V1ekQKodNXzt2AV9p9jFdZVttmfrtbQqg5xwgywy7+9/MGB7YQIP3
GX5DO0XjiBqZLgaQx8JztIf4wblfnsM1dG+K4m6GxZTvM/I9xdncaZJOPlza
8ZQm0W/TuLFVin0J8ajVxRnCGgBF25aLLt3igvYgkZqg+OADAlCwEgLkZ2w2
IFCvZT/4UjCJiMhYc05yDHWhTJBDuFfgu966GsSWW7ZWqFiiJvSroJDiqnPM
eAOJLTpeEry/Zyp/h65+CJ2SFwqO8p+0hW/sF1Q49VopfkzyLcDo6LzfwV0g
FqIVuIqPsiyzjbCwGtYA5491Ox7u3Ba1VShi4AMb/PFOUYYkJAbtQe5uMp3P
Bn0ylsOYQLKwcnej8zdM2GmnP2gJ0weiWHxkr0ckfH6U3t11tCEbmvAcwf0p
xlKjlTmwe5/8DeWWLlXlrxrDefxNy+vTW3+atYb0PPTzwYWIiPPbHUtDvYsx
cexURm2/3dVn9r2oTR5WOmBA9NoO4f8chvRF2WQBQy0j4sh4g+eHsIjanYPY
hnl6Bo4DPe8evJsF7cNPUspr5nIGsbnpps/HmG2izSdh5qkCJQFXY/RPOavt
xmU7xF6mJIqxzlAEF0szMXAQsr5vQNAUWKTby+rRkO4ikHtd63N1x9jJilx6
ZnXznpniANQIV0N58J1M6ZUFEtK+ZNnx8aFimIOJtejWgxIYA0pXUZFN8c/f
4rjTFn5gE9V7s5c/Kw5pjO4+rCc6Kav10ivh6sBpJxxbNKqfGjCeD73sV2iI
EGF6Y/cmH68RxAQZNXeftpK5wpXzXL5M8g8OiyNx81Z9VSYk5jR/B/ThGBD5
Ktcat/NFjffcNdwbYoMdtO3GUPfAi2BSYi/0shSS8DxIQpdRV1C0NAeJOr52
xP6duK8nyDWEh4ryAFmPR3IesoA0TgTxUVqSl/rpk4zJWH366rZMwHlr7Y5A
WBHjj8jU5Z2hqGJFUXTxHyH5gngk/S9hf+jgtEmoekCscuGte3J0cEA0kxBo
g1ZGm6fc+0Xhd0Qq+M55mBFZdBpYNiEabd0XzSc1XYPwwwPd6Mb0JLBX9CYd
PtAqFI5+Amr2OfjQGrlHJeIdIOQHgky1a0feukQL9yBa/3YwxNW49v7heaRe
oyITpL/Vw9GYte8BGGPsT48TOUh+db+fTyCxEF+KXlpvVW8bEf9r9NpQMFyA
S61ODEvvM/qUJBORdbhbjrpB9VbXYLm4ywFkRhymNZAkPSztDufYL4QSJQ0i
2txFlh+/P4TWK1GrWsSW3NC5pmZt78CpRry91fVCTnGfvk9AFudtsEcNGfuC
kiECVtXn9vtPZZTnj8V+FBdzN42a2cZxCUp5pvTjm4gDzRgcZXA7pAf4kx0b
EumcrPjHqFpHdpUtQAYEqTPW6fb3lfqE2itdM7Eiv+p9XMOlav4gbkUHOq2h
y3h1sqPzdOAjY7MbYjc8RCNi2dHGkt/57NfI+4AIXyEKzCfxwAkRYkxCN3UV
8g5hAYLqLuLbX9nkywWDIHgGLyEgF2LjUaU7e+ZzF6nW0vD48oOzKVfKEFH9
jmCa1e4qT1TS4DxoSqPQR80QtnizYK9TpfKIvsre5DQ4L7TMSNsAtaUNDTc6
i2rLLdXsOdBNrY+TPZDzdJ/URZ7I7scD8rvM1SAciQitsaDZFOWSTkx92H2H
gjQ8Wsohojo3ht2ZSyZTijVfyoqxkL8DuXtg/FCnEZMu7jxoOMWGW3gGILiv
q5ZDGU9RNsPn4VfdDFR1Evg1qoT+lSErQAusGvbS14GiayQ9EnedVCg0Ravx
QB+uBTdTbquz+zDHDHGmg/BDgigm28Kx0H47+ZSEeTxcTqGZXDBAKXj2yogZ
5dsaeCecm+IXFzLkUja0aPQcHtcFypCa4DT5a5ZbnYxs+1fH1lpiB3NCp1Pk
vSKvgZsSKf1WnYmzVhtSRWRnZJLlwsftBCRSBDrqs0NfyoJggUUM15H0YfAb
wVxy7Ix9lffrOtq2g+CgnBaaxKwNiIjqcZGyjShW84TmCvOrnfbtD3608Bse
mo8R8h+E+UKm/m9pWGhhkev//4if1wfjdYjbbpMj9A7HOKcsmAHnPALV3r5U
3NYnKady0gMHup26Bw+BXgmGAidHJ4ttZfn3eDQCXhFGnDRTg4tFhiHDfS45
fIPiLRycM2AXp45aOppGOjeDEBagrsif49IN3+q8eK07BhwwZRvc4l7IFBOH
7W3hfJ9HPoLaTHN7HLo+Cx85D/Wup7wg/K5WC4XqI2fH59lzu3rUOiMx3ZjW
OCKknza/Iu7dmuN5b0cm+91DkstZYaHEOfgK1jQUvEg6XjzzI44oKhiYvTDF
3icDTJZvc5V7wdEK3wVxq0NcvZKaUitwHCIBWBAUoKy2hOnim+Tpfgylzb4z
fN/ARc7hLWuHdjkt4JvEIu5yiAFGIyfRzdIb3XcL9gfTjoUfBqj+pqbcZLur
SBpZWsA79aDGbZepE8bmSXo3+tlkah3LyndIH3zEKDqyMUZr00azeR270vIV
q8Emao2tkUzQPv2UQtbUwyE9dFQLKcybJAYupXhzL4VyH3dI/m+aJ4K/+Agp
KuJpEx3UnnyIWw4LeeeLYsKl34FMWvLiDRcOIYLngQS1v06oxlM7Q3CB/43B
bZbhumIvs/XR/Bj0KyMDgAPTbpxvb3wiPQfJ5dGM/A9edinb7283jBAbOMYW
+5Y3x2UOZL9MXtJ2kEGQ5XI2eufnPqdVdVNqBlQYg/JbMUGhO07af7YQQ0/f
4nSBJbTi6CgoCDhwfwI+NVe0Y9EdaHYUAvyq04OFzXOJZGxyKaaaSg+UE8RC
7156Ko5kXO7klCiI9w0Ox/nUzj+828MPvuka6Itkj8tiPPYLFAuJyyJQIlrJ
JmFTcOOSBqL0RIiKtgT73yST4xZw8H+vU3jUNRnpYVrcxHqs8pK7235bpi0r
2/h1/2zacfWVUaf6sfgez23FUv7RnAKPPKcghPIhtb9PcMEwkTScs4Bq2Xfc
C82NyVNybtG6HrIMnCkvWbmO3bfxGiHfjZ1x+nB/OZ5CVMCQ7ZYjhUs3EKj3
Gz3wWH9KWZugEMtqiNpZ+QtqzpU8mLAwkWDHAdElvDRitxQLPIR9Ph6KD/mF
bVLCR52k+FPkoWGhL8WRq8bJ8ZkHWX1FLfwrGVP5c71ycxrgdbCAPNZR173X
e9W3gZvD3FjQ7KzSDANl8AG6FG8MWJOspDSXu4KZGUGyjz0RcfxYVe7+qLZp
GkiKibVHB0a8Y1RIzLlbz1/2f5KADPlFxaPXJEMMc+H/vTgX2VqURiofs4Pi
lyClQ8NJGXDKSF6bTfu1J4OaceqGWeOQFTgFtaamHMXY9rmR38R2MlJwBSzC
8bs+9h4h8soiNHVVsVetDJE42AK0xXzwmq3W9SMprvzMN+F5rj18qyVXUfd8
RnsdPO+YijOccx/nsExeoqI5fQKGabxN2eHUuGCr81t+FLHywGuEFcvBzy1U
QSCGhtbP0BzlaywFS0BbEgO/XUjJudkC48Z+y5xDdKuvGNoj4ryEjS21myVI
mTA3+mmZ6uDSC/jte+/aFNJms6xbDdyqMCORU2kqwcUpkSUqYIWHG+hWFxCL
Eqdp0Up62oDwCpzaANa3ZrWoAFIhGEyLxhlJsdsGrXgkODJWZEPaKWc/vgoC
/z1xExg6XOb8LndYtyeXezznePWRD2//RJhD9gKscau1HUG7otD3U0hQNS1/
pT1L7wqWC7GEhGRHfdU/aUXDBX9hKm37jQUU73xWFiFkwGZpBaVg/fQU0PYv
WcjAGss2Isv43J8+oF/4hOOdMi28oLJpksrlNBqLGcijH7DBpQ7xFwyxe0z8
OOxCrOqFX0hBKStF7PUADlCThDNHfHq+NKxwmnf4PqbQGjIHbYu5V/Ezuz5q
VXMyCj1nbK507oUuI0Ulai7nMaEGJ35gAPLoTPPw4N+vd2FBYVEHh2N0rzWt
bpx8ZO+yADNHE9n83VmdJXgiEJ31fwjzyYtWoJ02Kws2M6STExfxhKltodDf
qbtGZIpnVtRIiB+B8ReUS+yXmgz31SGBlxmH3EbhXX6O5au3mfE344ULLp/e
srYMDhx8TEMjMdMQSkKWaKwjodg607WY+q3Sf/Ed1jfwtzqZXenTpyiqbF7v
McIV4YsXOJkcLA6l2aKCXadFxxdJTT4l2A1VueRGclrc5uwyT0aulRKi2yFc
Yegi/hA1SlbQNxJ94Yzf2J2WMN6NHTmQLmJpvpawaelxZMooR6Bi1FtqPR2N
uQeN14E/P5l3FjZfXIalbq0Y1y1j0WdcFPE02LILl2OaNNUT3m5R4D0ILXRO
VTGLFqjFJFzBV+WUR8OaptHQZoisYjttWB5eXmA2M8sY+rT2050JNEcruW+O
mJ9bC4Tb61POjTM2P3NhSw0LJnbi0ow/4zRoY06neQ5D3Uk5upeMMBlR86aG
6ILfhESDdXLOcMwcRt/ODEYwLx8ncy+/hp5zBpPVLZkDF8sOYPmSRC37oF72
4axVIbZYT2TlrZa9U9uvx9ctjU2HfFTLj5V89g9qAg1eGeqsWRZhtwRW/h/S
IkFxAef/0WmXz74BrK1giiFpWiqq+f6sCHaUBMHhSi2cI2Kk1+mSLaOrV/RG
2TPd1oqRv2Q9YnHDgDywHVNaShdJQOEfhFf4b9dzDMHO8hXc0oAE9gRbKIDY
R0V2GR/fuT+TYfdEd3RkP38msmgRINyXs2yZunYMnqB544i4XqsW0LNqlgjY
cdd5Sjsd+T6wqIHRwU84hUFtFzHQX1ERv50iPPGzmt7c/GivjbQhC93n9fL7
LLs0V6J4xmslcpo4gBeuQprwI/qWRwstuaRMHssJD+sODiuTCGNadkGSkQxt
5H0qsNr940Idd7SjAtkoZrPVgA+AAqk0ZYA5SOFUVNth5jrOW2yTSE1LY3i5
BZFaSrrTSxL5LMBaDPBh5THQqJ7z+W86/QdcQeWOy/4SGJgoOUie5URv9sUJ
dBgfD4Gh7m34KXbwvijIv2616tUNoUXBjZ3EItS++FIcfM9TsG3JcL5MZzMU
z6U8vSsYf2IhXvYQQc7NqGIIoAumXAYfWPd7AsAt/cpdMxVrDROKZv9mTH+V
HDekUDUM5+AO5ch8Z+mra1jDEMRFbDkMkRthJsl3OVufi/lV9R5b5HdNOW5Z
l34uLQvdojBo0WTGYD5a6NiY/5TtY1J0cyJVAz1btdFHZoNvjiEINBZLs4uj
pp3Xi9tOULEQGLwNKxcEwI61w+UFa7yNmRP60QhL/1DC7F1hNju7m7lhkQYl
i2oEbpwQT9+46WfCESgf7dcf5TaF48zylgWS54+gSN8yibTHCxiQIlA2H31Y
5SSnQia4NuUzVN2Zt/6nIeOHgETvLk3YgeD6BTCitKrTA3W7paa/mkZCOZmR
/PGLhneyDNPS3DdREYpQZEZFw9Lz8XYJfsXo0Fbrxfv7rQBJNBrfrdo1miwZ
FL4aUGS3BD+5IEGUX6E2WGsS6gUfLUPnBpy5KlIR3UnzBPyadMRV2Wh+Vv+i
qmVnyfW87WD1gfU9c3++P7J2hZsDWS5C3bHbSro7uvCpSvg16H+9n4J+E/zc
5W/sPP0WBleFKu3YowwV/qTn3jtiB3ggHL8noFD7C6jCaUiopSNM+rk54GMv
ketD2tShMDJ5FDxoL5Qbqiyq3n2zFX/4KVJQInAHeehAt47NRwoIXN1X76Mc
7t3cIo+/yWAzCeT7gFf0bTPTyHNiK/5G0TpvGsmNILgruWuSbyepXG/BcN5D
HJVssooUXrK/pfEQl6c0764XWlUUkdZbh4hSE+ezZnsmWbljobMobxdYf0DC
ZqV6KCaCxZsp2mPXF/azWQNNhsHgVFPUwLwYA5etY78NbR3PbMPXcwGKImb8
zxitwKFQqUBo2z44NAsQsCJbRHSssOU69G/yq0vMOmsIT1UaCJ5N18PwTEFP
yZ9kdUL8girZH1eb2BYfe9HHlw5jGE0MaO8emHM5lri3WtWAAF1n5kMMCioD
kkmE7hvvlBtUQf5+nJy9tg7uCXsik2WXT8yWrpLhsT0e9pFsYeHOTsL82PVr
0w16JeDmab3/SEDt+QwbaOZOYSCFCYNmD1UVu2jnIffds/zV+HyupzlYaa7y
vjZVX8/lpBK/lvN3B2QpFwa+usXDgww4mtvLHgFIn7OG/qYN2f88pPQVn9DP
x4N+leC4ZG2WTlnCa0xmQyDY5M0438BMMuprpeHNR/1p5A6FgkpE1lXzPRn9
7uL3H7vFK4qx5xhpwq+kCm1iX0bH4/70j3D9FCp2E4HKExTFpn6XWZH2EakW
SOz/At+LuS7JQ8EUlJDPAeHtB6obH+PoA72XpPq9DgFu4yF3SR+5diGWevt8
EAO3+TY+HNr8FXl8omdU5S4qhuNoQkvifBBFxEVxJmMSJyi3HmZ8brN3wjZl
H+15GE84AYYvxLGlGAicjXuv5BCD1v+mA1UM9kF1RqOO2uCLq1slzJzs5Rcw
bRadFjEvM17a5HInKnprr5YfRKfeQtS9cn6eA5iqGAU2XepG7gMTx5pZIq98
Mk4TrHyjIh9kO+5BWh8OpvzV0rxIXJnz58H4kFOiqGHoyv1VA+bxTByzMJkM
PGE1e7dYWuzq7pb+5snsQGjtcyFffIjJwXlC7FpFRjXtwmCWh8KMReXbAh5x
iaJAiiwGrwm/mlS7vJE1oxvhx9suPK0d7bEBQZYD7zLUI03FPny23zLP57s/
Q0vQqfA/Gd5Lh2IqP/Axz0Es8hcl8xr/fRDBI6VmqekaJxSbEoYztEIVEa8i
jnmiPiWrfw5ycqLyOn6wX0WQpUNN8dBKbts6F21tI7a/wfZrFyuU39LnnNOL
Jlq+1C+cBupCVWBOxa0W0KgJ0lRk5FjtmLB96f+RWKv9/RiLcbglvNCj1muX
ekZN8/SzF07gBfY8FfgTYeL98nwZ0l+Ot9hR0/DO8jfA/veelF/rdLgvGyoM
cBDCI+4dRst4oIM56BKaKBsHvx3g8R+eVsCZboTGmM+1JaR/9nkfxPHwkGDm
OtOaJAoE5loe+DW+5lhu+p9jVQ8MuLPgzIlQDUv4Cl8h3dN7Od6NecBXHxQk
TGHRP9H7uHnjevglV+PTqx3ku/S6Dpdz6f9WnskOSgDOJmUzajkjO6FBpO4K
Kv1l+93omxpo9DLBqdZU6PvduLQYHLh5Q5q3ASS6adJG2mqiUVEjeuUYr+iw
JXTgjiSaeZBKELIyAvy/EYKNIo0dsgWWb0RY+wKm+5pNriqqygk29P/Webum
/5v19SADDmnBt9Qw+i8M3ysKT7tfui1hTy3XZ871hyMSChtDKa4Yu0TUc9J4
eoL8hRudhuorDqDcDDEIXx9AaNPLhzSyqj2y6jhW97w6XK/Wm4tDZvNj29Sd
aC6IZ0BFpekTkneyFbBnzdgmf8xTuy3M58uwdwHuad5IbmZbwDq1P2DtGAe0
vciqmuOX/S2cWvT4ej5DsFTAiQtQWWvf7iXPyjBDvmMD1xOAC/GmysNWsUjr
CKoiK4GE3eE1l0I2WnBsBPR+8DndFbBfEGXnDQ7Z8ImCR/uVxB/TxIh4udd0
LHz+xooluI0KRTYQWmbAyQQHqbgPEHSiDxwNgPQOs5e1KQ6B0VqCkiOC1UyJ
BGvjDkPokCX8xCDLdp5udDKRi5dCxuq0SS7USQYzbLsebu6pJar1ubQI+KJ4
O9y5waeQDEIn4eeC2/dw6UEfbjh0fJaiaoF3sU6Mb/1lm/F5xJUM72zIb/Om
3PP63hbwXKC0d2/S2ie+6QcA8d9yLa9LtNCie2FL9IHD4qUFqleUhIVpBdwD
PTeEmbs9nMPLpcPAqCre0TvZelOkFmV5ZoXBP1X4gyvgZhSN1cxz5Yq8Yoog
EY3pYqEC+RSqp5EC9c7SK2s8m6bO+T7n8E+w9acHPx3SDkKJuhpBkDl78pJ3
xMMQ+t1/zEaLUzq1BWV4yt8txzEM8jQZRrpyj73RFX2Ka1pNoJS/wAQPUeAw
Atps7S3Qea6BzXdx7YusaHv0aE3YbqcxRcgiqgghS2fqPpqgznTY6RSuP+xS
kO354WNKWEiF1rhM1XDLWbh0nJsf+xHbjuR8MCQLLDlSM9D0ndZER7j7Kr67
v+FxVCeeriyW7/cz/6wcbvXq3A3Gc2cgwFkZbXJfSSEmMnLWy73a6yE2NJ7j
zUug6eTbsuCrmsOQJ0UJD5wvpuu6Jb+XMUSrxkY/RmJVNWO/M5Cr3JE6uaQ4
UWkbdgfXtjJ4HmsYn8yazBboZW/Cnc5SNL48AwX1TKy2OS1x2bt17DBZiFIV
UkbRixBRDZtR1bKJnX5aX8ERS2KiHZ7nc7cjcGo1mu2Xxr8TnO9wiI8Isk5e
Gh7Y8/r8eyN5xy9NHT1QMOd0Zy1WLIUVolExsDRTvzpMgYodcra+VUgvfnVx
gJwDzmwb3YpcM3TxloHMerlcQLh2vUI9Jfh3mAbluVNOiyhlMCTa0K4Jf5Dd
+8ibSzcwEg/hMhdKODs1T98qgzMjNwOxD8vjQkzedtk6vUoKQqR/xisIDP7G
s17oZDYpMsji84QS293jMPfJmyuEfcA2+XDAR0II6qpvACn4ECbLsSNUXDDH
DIQqyy76wVz4aI++xAu8uHsY8odv6wcV8WRHssOsNNRyYYZE7nwoXFlaDeAH
pnZ4idsWA+FzHPuynzqpMU2ghjiEV+/xI8BtZdzHlFsotEODyCudmX9/JrtK
5/vAnCmTyA5iZYmuWzoAxWt3z2Ntt43v3auszju13KCVcuDJrKLFX6HcBb+u
iL5oRauxrHa7jwktS/IcBy/eucKlACDwKaMjVUhoarOo8itHaOacKafk5ILg
BruQbBxL85NRB1CHHYMel129A9OrEgiNG/X5wb8GDHLaJJ96LJFxUiNnaLIp
TW6GdPShw4KGD9wedMD0QsaEm4gugcdDrgSgYkxMl2oUS3nw+IOgiTZlbaHW
aq/vmNHSZW7MU4wUlkYJnIQnV/vyhpqLLV6/GKcOb4KH2u0mgtSm4HGSs2KP
9MFSDcfXQqgNFPeyD1wkMIbsb5wzCqVhO5wEUvqg1yt0FfRFx3KSJXVvM9/Q
0Xu+MbndMMJRwxIy9eSQCC+vME5b+MLG1nRF/iogAw4eFmWjtPDcYqtmcx9b
aHyXhDOZ06HKujQSvmreq1LB2yBKb67ZIX/bHWMv4+mtH7c9B/VxZI7AfEUs
8lPfQr+mrposKGG2Dpk7w2Lfaya7pvjeoMJz7Q2+1ZyJ337BI3XU71i79bNw
mmdd9V4JlI/FOQoBPj8gmayX5DAFk5nMbYMBUeZ/yC7hS//BDAtc9OWMnntO
tbqqqQylzXeXz4UIVnSHWF4ulQPsUpdtuBSKWb40GOQMiSTOGq344umeW8X0
Vdm1apDz++C8Y6kDWxAnnvn20Z2RWcqx+FxxsPsnZhwTlIjtapAnsduTAHV7
hciULFyhMXOXGcaRELB5tkx5SNrzqaiW0VsI4KEpF7TcReSIvVHZs7KnONcX
zgGbe3ej7vS5W3YzGNfsPfUDanO+TghHr7jbuK8Gr1cClBugz1KCMCACxYOW
Eshp7WumlkR5xbZaXCrNQ+eArUCnnrWjJZSTGU7QhuMenuGz5p24rxjRfMQI
r/bnxDHTwSSxwrq4TSg09nw5rPTwVoxVmZiYw0keUKm5dzUFhc5YgFvSblpm
63Ix/gBQ/aywuv4ifsEkzj4fWI9+5ICH4SVJudQ9sQP19wdSm35WoWG8bsLw
L8eeQA9UjNHNcxrRvg30Bu/AKncw7Pw0z5+gk5Zz7nmGBm/9AolN3ht2S+Ku
71Ep5nkW68pAbvt0rpxLH76QFnaokVFXdic3+2HUG8sBhgEqZEjmKuEgCj85
ksFZjLowzbUdva9nq+OZItmth1Jry4SIYpKsf/Hmuc44yRTAk3HlVljz5rsJ
hkoy+Qz/W4RYC6Sxm9/PtGzuirTRumnHZg3Tt80pfXbFBTfYDBlsDZtTdZKB
g4EadH+pIGRYeURntfKE/Z3lgpjzcYoqCenMaEQfEqXuiRXG0Hoxm2aAu3XH
k9SANHnU846KbOMDlAaFwNj2Qtrdgt+0FeqOjHhIcc3KtkAzEMQUAGemNlO/
Etk1yhFV3178XSBLWDKXVrUrNqhKXJ3CVf0VmIzC7gG6xgGyXL7gT/BC5vL2
Og5QwrJhQTdLxhOSwY8+euV7yro2zc7rtKGP4eNAHFUVcHEL+Nv3815pl9Jr
SNOiQmaSKWq8orUtOPV9MUr8B5oyw1A2E5jjGV0uWCJaNn7LHkr9dkfXiS4q
TZGSYNHva47iS+jb9FYtP1vkYQGe0hykU1Zoe9pUf21ER35Ga4nF7CCwqKNz
GvwXqTGV+9UC+cFU58ir67S3oZfmzXKLsK9QT+wSNiCEIRb1OzDRRDVeYaIV
4naKoP+r2tWJPNt5pVaGBUlaLSb9mCk0d4OiFZBtalGCdjSDa4PBzZvzT03X
nGEw7TmXdvQv79Gyd8M3Sl9lou854ertaVDpZcYnXGfB5VN534MGMr/maQ8N
Bv1gGOR1f5HSQOKLpbcRI/WyQQ0w+P3N/kfqd29P+mHiTnX54HO5iHQbrtmG
MVLAlMI6Mt0eHM/E9PQvUle68K97vGllDH4Bs/oqYB6Qlos6b/Av1SS7//z2
BL7Zco1dpX+HsPSVeoB+h4wVH/k/+N0l3LRkPm60ETOrLQr+jTT8KJCk+n+z
9EEUYobHYj+XhyOCHgS7+NRnLNrUOOWT7aPhSkyHzqOtyNhp4KSe8HcioGdQ
I8+WJrB3hP6tR9SXdP9VplZFXg9vx4Ma5gzqzx+9HASse/Tkk2r2hOrcgqM+
WeJ28xj/lhfoj4jOEOm8aaLs0hbqzYIuGk25t+RL7r0k0p9ona2CtvZ/mbSq
X+sOqrE1ga7OewgH6NnYqTUpmPVpCVIEb/EYKkRUX+yNtOV66cUG94Ka/Fg1
d86H7ThoBHoHYD7x9yYf+Wsp2T1JjwbaEDEkLYv1N2S6srVY/bJCJYiy8JLY
3J9XSEzlDC8UVBi4DJi+qBrFPqPSpzROdsu7dp/M+J7usXshtFqULUoe6rsK
suuZq3l6Gii8X+E+A7EoHuaQ2UwqwDRfb/AH604IGjHfC7BQWFE+B3tEiZLO
aTHAKh+Tp/PsdtwRoKeeDgdpjrGF8TB6GwH4uvoERYOISFyAda8e3OgTNVHi
J6uUGt1evELCA+5+ZUoHIt5udFATuomb9O3i+hEcaUQeu5+g8/Sc44nU48pq
2bAE1ET4wZEs1/GPiaDv/Nhpstd/O4cJfXeyN3DIgls7AYOZGA+z9nbLUuVT
zXj5Th2HA2T/u9LPb520k19TZl4LxvVyWXopn5XoM7xFbXGBzeQnI7iyRIAd
kSDCtM1cqj2C5WxY331wOIBRCWLGV8U747F8Ijf/cBUDbqBDZpe2kILSRVRL
ccLuf6MeSXfeH0SSQQyAjps1KOW5waojhu1PcCoShuJjY16mrlxfzKYH+AWB
ldDU4Ye/PKvhBx2wSMTh8pWSIMguBTvvu7qPVv4RVOJuTtwJEi8X7LtUZV5z
tLePJ/UQUhvAcwGqTbGaQ8+9oUikjyTzmejDPwz74srfJSssrRRzOorpz8s7
fa0R9dZ/Okjep884+islqCuv+qwluNtPkqXACn4hjuSOfO4UV1parR/o1JrP
wC0+KfTWLQsWxz7WdWupat2LcXRHeZLxG4v+9tEUK186BbNB5pM8ah7j9ELZ
8HQMULA4+rvhtzazl4hGEC6KwdVvDi9y1Cdz8pssDws7LtuSLiLPbUiKBNUP
pTzwa3V28uhINB6mC9gqFZLGZOH7i2jiHCqzX5NzTBmJ63CGz3KD9oBqFLYd
9YH81598ASeY7qUlcEq5hOo/kfA8ixOi81y4dm7cj3XWAbT0t+MnE+wbtksE
eANfGoWlKsr3Y85X5XCLOXU1Wut4Eln/7EWbQrMmP7Rvt4iFkK/GKgbniugy
dPuGnPU7vr6tuoA7rtaBrldc2rhdx96M/XYM2hbShUaaNf8ixwQSeZO2I4Yn
2kIDBw9f9GSMnl1jg0NHFtx6ZcPUtutH3oIK8I4cJOWedo4hrlzRjiTcp199
CTcvNt56bo2w8O7gxeySIRZUJNyBf1Yzn8WmK7vnlfmAte53B8Yy+hrpkwdF
mlQmi5Jw+XnDTS4Ab5SiEytcmSc2a6Rsr97cq+kf4I4rr4Exv8eeEGZ4dPBp
ZK+mAFS6+kgyJqyy2BVKG035r0XqlAVznYUms6fDd7Xe9zrkxcCPkkKbzJh6
akEXZRDeE4wy6Oj1f7Mo2v+wdOkBgMCWf0H6WlY2TLCW2FDJFwKL/D8cucOS
zQpTJBfvKBn45cpXfqViRfTm80r4JpiHex8IE9VoOA7VKXFP1wk2+UME2T4z
FWp/LnqQPSpx0Qo2kpebF8+x18RVQYNLYZn7HuL/JQlYY/L9M+MKMVHfZDaF
q9tcpeufNMwn/J6q5cYZDY1xGq4nNJGAMghmd2tM0mmN48z8aNTe18JAhCvc
OowUYQQ9peM+bGSruBXKxudIltF63LAb5mZ9u4vTbJSHk81NN5poxOUae8Q5
ojKzr3NHwHwDf3fH/XQOczKLLW++sT7/5MbgFrSzyXRt1tq52E8iFvIsLAb0
txfcBvbx5XV4cYQSfB0l/GgP8loAowFuWTatEJU2sKJt9kELX0BTAFtaFTu2
Stk41nShekWvWCkBnS67TS6uDkFzsVpkSE/d/Yj5TMHpAMIZGwFSQRdvMVOj
K1ZteiomOtl4BxOFXzyfw+2qCKhyIX+JQIa6D0Ia8WMyAntYKfC/hdBvQMS1
bidQHWHjGyE7iuF+0lYsfaCJr1p7T8U+DsAB8yIgYVfKP/i39Xylfekym9iE
0IdSi20xfwhIhRFMB0Q84utBTbpTBWAwyU7y/1MF9piTwbO0LcWO+spKnN+N
7jHuohAtY4lPdD0yBY5kQzMGIR6/h6sMgMmzKBj2qvdz+SAGrQkuCiCUkUqA
f870hleqxcau3dtJzBJ1VOq9M6Jbydd+716hQ3SmpiVRFJ2qrpsFiOOa8RzJ
dxzn9dYPcjT9HvMMO6pVVYdnhwkswWsahA5zL/+ia8lMzpr8EVUTDmMItqNR
PYPL6/7PQePkEARdL62oK5O3hrE8CjtA/MMFJHCr+NrCYGZhMoWIE6QZmJLZ
kX3EAHMhXvElkzXoIRXJC6oMR3S3TjYrjm5LMkKoyxUa1z5l5MZ9AKSmZeGj
/gRcOMVznY5xBxvEmz6t7H9T2LlvtaWf51C3GXkWz3H+lze8QMD5zxwFxqGI
EebpzKzEzhkwqBG8ll+Ep5zLXr6+myU49UNTTAihZiPRye2AbYmukgjyqkCX
xbw09es+mH69nfoq/uUuDR8eCh2cyrn/V85ogJViOaI0UadE1FbliUNlt+1Q
caPJdYKVExBlliwHyThFaexfrJFyHeROYZrth7QgqZWeBN7E7RgpT3gg2LvQ
jVPgwFKV2eFAx1Q5cLjekbz4QUPdgxxBnl7a6W6XchGMIniLKpUqG2HoHYc5
DHq7IhQiOH68f/OOL70Uhl80g2U/GtXJ5sO3jCLzB+VwqRfKTluWuwoRhL3k
govv2Rzmo7fo7OwzaT1Qo9bAKeUVC2YCRcU+FqxVmzdebpoFZowvm1EHhAGP
0EjtmdWsG1UN8V0GV8IXg3KWQ7Weq0C1ZPKHK8o3/f8ip4iMiTOsDG6S3JB9
JlaN3nzqYDX15kyKrjZJ9dxpI/MxqOwnZuIAA7Y3Uu8ZSfdTFzdpgikiYXOk
gxz6H5kXvTugmKsrYyJdEkXcTFvX3Kwf4fNAKwO3o94gOJ53ouMVK4Vx67el
4IKprgIV2I0TJVAkZ1//Og0RCRouNHrlnmccsxZy8zP0n/xYmDF/U+rjRyh1
u5i3CHrViT+gx6UM+LSHEcYbnFP9JKGlEMRR0zRmLqSqEY4Ow77U1ncHfW/g
BT+HS80BAAcJwQg/JhdMzSJhV8DfkVyB911t4lBzBh7s4eOcPR4hkUqOe43Q
CNGTgYg8kMN5aKdSQ2D8MuP7pGktPtFGZrNmmOILAmEMlj0AsXFrhAM6GHEa
yJlKn4nWN/IShje1Ls3+hO4BbbjQgyCtTsgFHut5z8besmUazU8LXNku/G3g
dhH1XJJRIHZrueYYwsd+j2fDbXM2Pc1azA3KrB+NLQo3drxWQOqAwmIaH9nX
ILE6biIajRux9XybCgPLHk7HCc0qc6U020UiX0vQWIyD9iWBwsO70PgcNu4Z
8K4Q4BS4rg+l2Ro46zqreJ89p0nHPORIZkJpFm1NbLkbQCb2X+0XAuP8CseX
u/szdX4irF/ARwamwulLGuhTK/8NQj1ZA0nk3TkOr+0zUBG/ZakT7i59NUVb
I4Gga2tdHqXWXiHhRQYcp5B2/jSLHSmMOWh/nuOeFbqoDTc4oRD8zup9yTnB
8SdDeRWO/HHtPL5qgHBSabj9tXXhELWTGbyoAA6nDBQDXKHfQ9wn0pW8M2Nz
yshIveyf0I72EwkurePQv+wvAXF9rwS+RxObzJVphFUbSwr2ar5ZOrnPMnsX
nL5w7dWlrQGJfYAB+lPYsKVCKhVXlwVqoifgcRax4MQ1RyBrUFY14X7uGVh7
OIMSFDzFJbYsN/wUh6+PnwshXTBEVL/zoADnhznIG5Yg9p4hR6B535FAz2Ad
ZVMV4pRaJnSfm2AbUtZMg1/BhVuhUTw69sJPdESmOSkfry8hxGWymjpgzvjD
KEl3v2lSpM2wFOBhYRB/6T1HmtHaNzV59nvECU4Nb0gxJfDTEjUCsuUZA/68
GGF7mqeVYDWtc4pH99qF0sKAQaBsx18mr9yr3CY6ey+YP6cHhq6ky9Si2ZMl
90zGCt1gY+9oZ2NY7vyTHrayXOSgMzJaIFYSscIxn69Cf4a+SK3svnMWsLWD
TS3rDTPPqzvIvozlpg/OSNRoUY+tkbZadpAngy+AJ0l4UkWC+PzL3ZEI/O9p
yBvcHMJXwLaxeEH9TgwffdNzcp3KlSnQyP1AKkjER+Jgx6FmYu5mlQwlc0t7
9zU80yzjYq/5lUFtrV7nlCUa8h7s3lYx8FUs1HUPcbAiBZZPgOjuHFPJKWo6
SmvqThXWqctPUdMWahCcL8SRRVwWB78nqOFhvPtHUCUeYNoGm+Fz4bZySz/a
yoKueq3ABWwoJ0Y9bomfDvP92JiSY997rZpaCHmu/TJRjKfrU4QU+IIIGI04
3NnWYisjZ3VIYAysyqLpuAG7xf42rA/N4hn0CRMh+5HHem79DRe+ocuug81x
Jl3lomeC/3AuyrwMGDJoJ78jeLwteyW8ZubJPeS3RXo4K0ykEqb9ACfdJT54
v7n4vbmaXjYrj704PWf9kSyJnVM2OiNS4YQAxZKII/hrms1MjwvR0CIMgGrB
jQIK1ThgQbGfsqW9N1kgnQOXlCkrqaxADTc3Ibd8JqQLDbCsJif3HWvsftv2
WgBpJeSXGe8P354CkG+Vgk5orWpe+Iv0lGljenczdQHdRCgZ2S228C/HkIGy
vxfiYFVYRtxrQumxgVlLv8IBOnuf882zR13lKtqnYx68Ry7vWUaspCMMqmZm
90moPWVV7OjF+4DNMcxOpHOs0YicNCU9ux950h3dXdJlzzfZcc6elp0h6G/d
hKskAdGfpcl0eT3kbEgiIxxrdeCZzN1PDCEaU7vkWzP6JRhhuRrFCkCVE8Q8
UE5N+ld5sCQ9RDLnxsOuJsubQP7wE1v+7mOsXg3zNT3mJqGSPwHtZ+pRWTqK
g446OAj6cNBziJdgnXesJD0H4tIDMMvstPZkd8ga7i3Evxi9NgXTUfqpH55Z
aW0O9XB2z29m7zFmbAXanzSqMMYHHkd0mMTxyeIL51ZNyBaxMd3D6bZfSsB4
uPzbxaH8vDa8/b2SAu1LRWzGVd77g4tqao29LePsTpezXpnvgzYdSflu2j9O
2i3Qj5h0RHew6V3CEC516nSG5zwuGdUNQEfz6j0Y61IV3nSO64LZdWtLvrqG
X053+e5eMgZ+K2O/SUEyV1UXqHcUQ0gcsy1hg0FUuZuDjIcj5qmxU076+htl
+TL5OLbsqoPqxzdB+g2l9TjZttpezyeyHp2G9x/DDJRQhPyWct93n7VIpmKD
HLV+wQ4UexhfMYg3EiKuV0Jtca2RZf9CyTOABfxxo04AROcnPWBB4azPr//8
jnRTeOAhQRBTIY4t2feYpv/l7vH3NwCY2iNKegbfZEaFDFx+AFesvUefonEL
BT2HUP6kWFBNnFVkmepKidYrQSOkhL1fHH5lztK6+tb5u8+Vp/bqKw6n6IVO
gVZ0jE8QMaRUTREAmX1dpIHqRubbL//UeXVhAN5+YQr1d+9Px0QLo/HAuRlZ
Ig1vtQ1Faie6JEsoyQCDUgXkU+MlyKVK2YW2gYUFOL4YX6rc3zfJUUtGp0BE
BAwxBfGb3Qycs9Rb/2MpeNb26jz4aU8cNqAs/H67aHPMdxE19Ii01a7ITHCq
iKIBJbxMT/UjczhbMv708YSmFgnjsbt61MGAwp/I5E2UDnoklGR++eod0XQj
uE/XHF+dlKhRhXF585eAkBwL7Uu+/mw1ytPtbHbKdbq8TIP1/W/KBjeqkaKe
H9dPchffhr7YrqR+LcxeSOTOGuCMutC45w+5dof1E4PRHvaA+qTt7DBdVkgi
rTLRBXsEUWLZr0fBqp7JX+E3ZQkz1ZoF53D/TLaTe96VbaMkbi7V9rte/AfJ
ibwCyJUQDWh71x74KcsNpHRI7o5whsYpkBeWldSpJ9Q2+zI7r1g0rLzhQc8d
mijaAQDuvmdAGBBHSZ0YZ/cTOLbd1SbUOjIQ6Rf/YL4ZOv0hSG8PLmrO5tN/
6uL4a1SxlaSEAMw2/OZ3QEaVMA+OJgHdKdmCiNLZe8wnO7fgPpKPJfRTCLwe
EagoL/ovrTnthNNSINjuKC8amGaAcEu3T+Qu4NvBWrO9NjXZxN3vszB5T3zz
lvNLNcXhZnbvf25ATHzC6b1Rk30WERfs/7tO9dwhoAGTgadNO7y6JvXhpVNb
msCTzzUlgBrQ9tE/lmONl2IzN98/wf5V3YVBby4yf02EbvlWyzUVmFDK0xtR
yJX9KFUtrFVHy/DBfzdSM5Qdc/Lc0MIMs8PsNyz4/UxxoQzlqoXH7ppFglpb
4BHZ1hoxYsC8OEoQcMxi2T1aiXScIgXMPHDxQILH8nGy/EYRHLhUgHuk88df
rcTbm01N8h1ERhaCNnRAmpu151WrxhnLwSK7WOTwWaODEK4atFgqAUm9eZfz
96BA/fBvuI5ducT2Cb4nYLHwXPybQJ5gjjLHB/gACmSxepZIclop/PgLvAPa
f5lESbv29e7Ud2MXMXSO6niTX2vtnDIXO4vAlRFjV6vd8mmxEBmNvV42ly7d
b7fHSN6TvhFs86jwbYIkLdMPm+oGJKL5iKxsVZm9ELKXW9ChSt/A4PiFmJU9
OIWZUIDdBDkCdIMqdBbB+WXfYkbwwQl9XiXp0LrvI/XLdW74br3TA8s2YtN7
QrWxXzZRV+c=

`pragma protect end_protected
