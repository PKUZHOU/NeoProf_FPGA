// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
Evnpo/N0p5FzbEBVwBLDe9tNB4PCNeJUMsF3LFjm59wKB/AhFn22IDWTCpmQIhj08mDlHgKmq28u
pCbrL2kfAP8S0e2Gw+SFAxywZnRf+ncrS9JjT3OrAeBjn+7h9UGJDqNg1A0B1OusSRQGRkob7X7g
3UYigaHH0z/LyzxAlQdpMfCVknDfEB34ANNZCXqGLE2Hp2E7s7I9wpVD3knVOmiDMjNYjKprMU/b
JYQ9LV9V0ZAN+fMEQNqKcP4ldgOPFv6H5Tcn73lMPmQjmiBUibFVTRZ5/6XY6c86JKVbqscoFbdo
kYUxccUoD8DEspPUuBjsl6gpTogWXEM0rcoCtw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 91088)
PNBUqIujl70oKtstykwLeaCkmUgfi008A01w/DJCfI5zJSvLftQPhWDXPaxfFkJgupqUMpOjDkDf
btFzAvr8cm+8n8iR1M4+qW+1HA93VYEp5G4HaNAOBy8U6EeLog/9wS8yt02JX4OgsloTpdVseK2D
ua+N7WhOZmjQq84ofvqR4y+6nplOA5owYBbYvI5iC04L/K1KBTo6hep/FVYH6tJbY1GHJ5gg7l5o
lLzvvTSragruQ7NGPHLy/v8Gc4Og6wo9kG2NTKQ2OM8DnO8KTGeVGSAxgH1jBwpGYQ1ELsrQcePD
YH865TEwA/pTpJBkPXEfJbTORQifo5AQv6IVSt6Jn15lZFFOpQFI1tqvMKnWnMej+SRpMDqBGV1e
LlsbSL065ota5b64P6fRRqQf9iVjKONP9VClAtm/BgVW85vE9fZAU3BF7+MzneztM7gLR88ei7d9
YaZNUJRKN7DcjzIAjGxzsoQlwBLdBOMvCz6eCpxlUB/mdSbc/WFDgAaof3tUULFKmUFdNpj7NPqM
BeIKF5Ouqa5v9+7kAZl3e0rau2nrYNV47ZeUIsdPrIaJpfDn5NstHbu16WayHx3S35675CFd1HXk
3sLY5aZDK981uTFGAWVNX4mtsOxYlkUEQIIZl8aJ6RyAbUUQURGGAWMClJmAeFvnZY9OaKuArjXU
0RNmvCewdbLsV/lG27JcER32KpInIbLfR5cUHNU2sJGmeglVVIG0Iza3EPuGlpYt5aI4jwAQbPAs
cxFA229BGSGulD++5K978fkZYLyIgpxwoogcyB4JfdMZsK38RiDONTDGrCPxwgD5lZW/mYEdM8iX
jODcGkZiPTRnLhNG0rFWaqjSCJcgjTz8qWBGWA0HyQeAsrpME2Ze0KQSUToC9ymQNZ8lTJLUDE7y
Xu5kXjFtCLrt2+Hu6cyvv5OttR8ajp1qk+PJCzfBAj9MuzsslMJlYYQ+bNFupbhG3/ZIqVLRC+g6
lYw07Yp8NESOgUqGCy5RoGAQqHvyumFIfLcP8xO+lUq+GdJJqeynNiA4pAnuz5W1UEm0S17Y0tUD
tmxvRBrf38PkZvNzV/AcUcHyVELbmEV/2UY7kXpSDrKSQTXTSyTxkilLmgHdcXVDupT6Iy7X0GDa
Ea+lM0Jj4T23t9md7XOIEIrEX9KiJjKfMB14vvNgzl8xccDMS1De9x0EuYY5n48AlvsRlHS4vxE6
KxgFoHv0pLHju3AzF/uTP0eu9D1pa0TUswmMV1RnpA8tUOcIra2+seOLXiZbgYnTOO23eIaUY9qr
fWLPAZayps+Avucj+uQupcsjuOCN7/4GuSmoTkusosQtPm5dKyewhR1dsxc0d2/WNqH/xceA13Ni
Wq8v7fr3F3XeK8z5snu4IyKczWQ38Ns+ZUU1RWvpFfDeRFu2Q7AY8d8gaEqZAPyFcxEm6zjdDMTa
q6zKRxkhUpBQXTIg2nG1lA3qKws5CE5WDzDbntmNNhm9yHz/yweyRHf3qJPlMjysYAVKU9pxhtvm
lSqyL7TKz7BdBF7rRukd+SHp+HiL8CCvi2zRIA0qdXA3pSVxufZKcZRPlJ5T4eWeKUh+ISgOTS7m
Ii6OxT+7Z+6Ri+SRvFbvzp0PCyikFxsPlRZSEakeHrVIDGgm/tT/yyucrwmN/ABRQlheUe7fz5HN
XIoK7lql0YtHHgv4OMQqzZsPRnAEcwzC5e31zINamIcK7ekrq8TSJHTJChqS0nJztHH6IAAo2U+G
LKWH1NhzQMBuDtNk5R5epeYsdyBTImzAtdvnCq9bbWHfR4pNHULl5HhcPaLwhEtErefUBjs9AoTR
ViKTatF0kQbnjYbWXAFRhiPBraAyJ06z7kmBv3U7W84RJr2IY5Iqir4yoMKi6hvLOUx0IC82jKaF
pgCmZ1bAn7a5eME2QLGna8SVUX3E4OpzT6PagP1NvXry/FgQG34CWPpIeANvgiL21UESRPSE8Ahj
qiWTR+FwpwGXVGjCHiEEpAtcivf1UeiTRT/G0C9Ph1qRJrYZB6OkwRwpn3THPd3b49+SbT1v39rN
xVHzhkn7G46AyvszL0V4DDgnGHxHy2ST8wc96mnBCzhfeiH4v0ciem8R7cVlzsdU6vWNo/3iIzgq
RwcX1B/jasXegW97NRkvHaE1Om3nCclOta33t2vt2OiRzPuPG17w44AifPeOml5FtGO/R7kRKcws
ss1RhOmYrTnOy2I4kPtfUYPYB6wVeeCxRX5ohTKpSclT4iYIsDto9aPTyc4Ur2L1AIwpfZ5dSHmz
/mwAHtZHjLlV1nt5SbLwl/tsMHgArOrYuEEoLwzy8HWgBGh9WsoaAy0xOKJBd+UGPJ91aZUOxugW
UJRVeq8IIx1K45Ufczik9WxanRG+82FFDEXKqADzvqNiayG6+Lq0ZVe0U+da9hVaBpoF8Q7e+SW8
W1OmZZt9f2sRPOanXAy8bIstEhPuMVQIEkSgS9otEjNWkJEO6FA7Ace1VryYnJ1dwvWuLwrRe97l
tzbjmNuSWKzfZtyRsHw10XMLg4awr3mlpuPTzQF/jccHys/EERrJvaga9eiTFolXoH20KqvU7gfF
xiud3h5+XVYvV4jHI2gTYo6w2i0U/7JzKI2Ys5Ea/fD5Ec2Ky+gVYSPDdA7EHsHc430wKXi+LO2q
GnYrJrjnXBhZeXClToo3v/Wb0n0Ukh71mPaHBWk+Eng5G1kkFEodOuoZ/uLT2wO/0tXa04ZG44wq
QDKKvFIRv/o11bxV4UfVpZDulQSTmdvvzj1Q8Hs4Tfi20JRzlbuX1LrG76p3sMGFS0gm4Jak46UQ
6wkRt2dA2q/f5dUvAHgHwHQtTvRSrJmsqG4qtS0KwrLwY6X4yWbO3k6NUp6DCywIdVR77PsAYO3V
CkZ9FFoEFmy+8HPQVzs09IKRtb7BcyGdo0R6fhng08RUVmRHt6tqKF2kk9eoXtWpNoCbS3EwsNLw
GGegB1Jo1oIbfHBw6cCIukl40Wa6FbAvdOA8nn4Kh0aFkZvcLRdh620edPmNOxKtnqjPkCmIkZIx
67tgBsvHMi32oZL4D2UPwYZfk88Lf4PQfu1BMnSKJslVGbQ8LhPYZ1ph3kXle/AHPuu+XbBfQDNH
xVMq+EXOtFGXW3KGEIcuiHzoFhQxDeLY1/SdHBIDO+qJCFy1Q8FSivMyvIPihmMNpcg9YJ0/to+v
5tnZtigceXVk0+0JAUjQ87mLOrOFlC1VqpD8/s9IM96qsLdHRDYHikHYVmI6HX0maYeN07PJ5ZW8
OVDtac0vtEj7eCVrKXHJtRgI4G1vP8pWvyWj4ifReUQwozWIDfQcvsx36vRzgfZ3FVyAFewnmtq/
kC1oklftnA0Wz5+6HrgCjtOzjs5dJyrTYMEA11MbXcKZTq1N5ybn1oZs8XcTPAZe5lkyZuaX8Lmk
VzmBeL3IZAjK0Ky/OuYlbMsglA36DGe0SFZd5dsfh593zGLyfXXL+yrkFP0cjCmzxfjH7lBSFdgw
Ujc/l3FI1x4Yxi8z8LuHoqrFJL3N18qZkRDnKelmVsDYaQg81dIB/YOt0JqV/ZlnUMArIMiQPPHq
h15YPN+o7VF7AOAC9e9bItJn3GY1z/f0Kb9cSSl/iTtEYV3TxuZgbYowgxbj5YyzC9CtG1/kRFUh
oDNNFVkBzJmTjX4+jwQNqjCRKRwRWv12mfu8zEpsnZevnraU4xJRZwm2V/hf9hMHET3u0VQXQSbV
wWXRcPaXrU3TpoEeR2Tj8+t1K03NNiJQCOjwkOwQs7a7pv5lD8y66NvncIW4ed3zjiTEx0cyjKzp
y724eI0P5cQem4CtLzXa5EAdXMS5KinXC2MBHD/2YnLaVBZvB+JIWNEIXQAS+Dc5URD5bbe5TR1A
cQO38p0RoLOS48nKv7gkXf0zpKBawbvf6ip6yJeIgdZWvH2gRaN2LmcuID9Fh1gSgqKdghFZoceZ
fM47mC8fi0yT/A+w7JSlkXFIJucidkc05pIH8i0lIx0MCDzXFk3SryJtp+hFVeQisyAtAmyDjH6i
6rmW5OJXb333leY+6msCC5HM3hcMbKHKslw5XbkW/Mo+sVZnTG/+e0s3tJatjrIdGdxzQpUD4FXo
rDpfGDfxx6JCxGubZZyhauh3DEL65ZnktpGI9NN1D8Nxj3CnZcXiERVfz5k+G5S1jkkmfREoWcri
z/SKxF31mm7i1/RALHI/IagXWSAhP0TiFsns8nrZZ7vI2ROdmGXgCD16IlQqYiMtKTp5buYtBm0u
FCcVNYq5B6UzHuxrj3sUZg1qgaxW6cCWpDmdWF0C1jtKNjGv0xjSUUjOz/wN1IO43XObjaeKBkqI
OJK+aA9SUCeEPqIHOEZV4V39Y2/92FzKR9Bivyr1mLvc4IUxnKRi40sw7jvtpAz7gUBpBsHsjHTA
STvVgyQ8DS9xAaCnRqdoIj0Cy1zY+9hVW73fjn1Sp1Uuf/TEoaur80KfpIKy3fDT/C4y/zWT3Zqm
rUHx0h9O+07y271YZ2nDz4+d3hL3R12tBmDsKrKveq8QQNQlaGqoG8vFWVMNNa4XN1Ir3lhpoT34
aZtKdidpL78CVw6aKGTTqpiV7zmfFZbK5DtNan+QzAjL3KUTueo5734lBFurebmNFYApFnOrj+i9
yCJre2beu3rtzQHl8cBCuyf9rAERrHZNh/T0wBXhLrvC6h3GZdn6hrD4NDB2DabNrHiiUppMTa0p
PpfdHwfDmumTjvRrLSg/qlZ+vtdhHQFwVAeXytvDqsMTGcnFo0Veo63agFwwEW27MV5Ba/dySiwc
i15Huyn21f8O3JRVlyhuu/wLIp5Meaj12j93MelFG95sJXNYzMX9o/f/BKVeY7M9NS58TmpDAi74
7sgB/0+tvMZ0NjLEU6Uq9SZSyVO9Fqhl8TGcS+jhzwZbusP0qiG13md62KNhliXy6rf6tdll2vGx
Rx9A8irhLG3J6moq5XDlQoZx35AH22PC/HFMvtVLpR1Iy7Q7D7S62pqu3JNit5LhbyTDqwhhELuC
gVnUyAx/3q/ppxA93ndqUt5YP4Bk6WNLGbyHYSHt662Nok88BylGX2TzV7dx0ks+DQe01Zc9DDYa
Rhf+mLm38E0hCm8PLSnRxY7J5JOLFD/ZAiEq6UQ+S8zQyuYuk7fq0YGmtHV3c6eXa1ihKl/S8DBP
wN8goh68/6J3MSX5m2cBuTirZZPgBanijleJ3TwjJiUmKysferdUXitvsn63r9medO9LQNFfl0MT
OJucwhFj6QQwBd5J8Bk7bNbOW/at1YPIoBgm8cQUJ/1bmhR7ZKlWFQmcE7Ved5IupYjiOXFM+oia
KAQ1FJx9fi86g0HOP1QuYqdA7WYrzuj//8/BPQoQzrK0Gl2MKOnHywcT3btGY0ZXzbzqycQdA6hH
KIZ2YiwvtQvQeAXSrjhaxv+J9QD5zT05YYkb+1uIvUyqUY71QDyD2RREUy+5StwsfZHbGcRwM/k+
nsjZHK8BLHj1vmKZqMd002w4BEhPeHr1k9IQfifAAB9XZ3ELSwl1YsTlgh/wJ7i7ZNla4A4JuJ9m
zYuUEN1ai95cxTSg6ekailqQh6jliDIn5r+jm4FPnhYd+JNa9dV9gtALEXQpwm2vcCYp64hV22oB
7auMHXBmPRwgtOcClh0g8w+IUAqHjFR4Brp26KPp/af+Dpvg+0EDuGG63Or814+JgGSoGY26VwoB
xG5nB0rheHJGSKLBwdBxuhJ0pyyoKx1yKvIX6C1ixCC9VbG/YhbFCVJYLAcOOVMF3guI99bOJZ5h
HEBLAHnffdh/A4M19i0E1QZQhASsnLaChOEdAWH+UtaXqXEEcWvTyzAM/mvKYTueBGVSOwZ6bI3c
43taxiCRsBLPoPqu+sB9Uf3nd+YdHMCZSrhQmLS04uprqOspNqvmk0PBwDWvu5Mz2Z42Zn/jDARJ
u7+KUTlyrUq1jKWxvChLKd7CS1RZMErxXWfsWF6/+h/t+KtHj3OxpOl5+28l3XoV/6PPSugt8thz
lhkDMdX3r/u4/J3XPrSjH3BbXz+beC2r59EXJtp+FuC6tdC/J+FzYmMkIds5fVuYcsMrWXrSXDqh
xtZAaMqXUROahNiYNbRlmi7YAgVwIeut18k58d5K7qbVabjkqaaKzcjmHOEEPt3r+jGtuqnbGsvb
YhnwQWsSFqgopT97QZqb0QKfO39j7R8N/hoNevQliqaWtDpK+TdkIH5OcA6Ikkk5JgQKkcMsGVZ1
AtCodlyq8CYmZ5sqH3OIxUhS0Xn2eOE1k8BRXqTJAO83+WqPqRLZf+iRsdYHjJyK7ytqwNbmzE7D
kKvSTWdM4+C01hhdILBQDDVTpKdmLiO2276fPq6hcFYQE6dJTmJ6PxIQNowtAOH1CTaYsnqqN0g9
d4g4dkPEfyfp78vpeBSrbcsPptTz+5IeISYzBMKjumS73UMUVZ4DdJ9IU/K64OCPnzn8Xp9A72M8
ix5F3abLFLX4Te70yrIoO8ky8pB1BtMQbjpLbUZaz0FHQHWuGdA6koxdaLm0YC/q8P66dHbgH0eL
b+CspiuuaxyIqezGFJkqNy2Ym9uRoR3I6EF/e31eETHXMlAmVxyZW0uj5iewW08aBPf/G9GhIieP
CHbtTcHHTCXGC3Cm+njT/RHvENniaFP41wqiEZk8FQ67ryHMiG+L/wnzfTtb9fjmYEfILMq4h8NK
iOEPa6XW3h4cg+HLFpHmh9rNE09I2qx2X0hHpY8rbiet6TRWQPgCZt1zp8bcUpJdFA1l+YrvPSiV
Wo185VtsSMT1TQ60mxf2Pytf+ainoT3J0tvQ8nMdx/T8doAzw/Y8NOQcXDV40lUy642yV+I4mGrn
Cvo9ahB6ZgmyDZXr/lqp4A6/wp6/BYf84gETdXtddK78+12jTZAdqUy3tcbxjD1NknOlSK9CJ7cr
cMLNwguRUR46mvQgtFpc3mmQMLD09SKVJbc110FAP7dyKjXcJ8tw/PXbRNHEVAHGiAyQ9NXKdXNn
mh1E3PiDBjodThFfdD9+Eeg6EA4X9qVXGrZoVYGAU/tgl019n3/Hzt1ZmwC25HL1O4b67FU+8JpT
Rmui4yqt4sI6+qtJ59VwWyKszFWrh6H80PLpCtg+iWcQ2YoHwaMJ6vVHIWpL84kLcC1cCCvJ7hT0
cLtNhjYZLNbTmuNFp0+O/dyllirLWaSzVWZxYSE6AjmSIRWtosk47cD2AOvhncgeaCcupnfVz5j1
aClxwbzWqG3+K+RSh3VkCLfos6bbUqA4E4YgweCYj+EZHjKngS94Lo2jgJqcG552RHKuGgPApsL9
Hhy5+Z5WDkMh179QW3vdP9lhMtY/TxvBOQvSD/CgaGvfcD5DYlHAC8dlCnN5ILcbUqCq7HvKYRF4
kXH+q7TymZBuzsTTurkHbxdjBpeUAgffEHTC9TmDCdN+2vqXIwjsP9FTRtoR4R6Lb6BiMznW/bPn
ZA1CgmKgMQlA8shAngVKwz9ObmzFd1jzYBI027cy2Lu/VrWKZrV6yvEgp4SNfhkEIvpsDkF8/tiW
sngt+giMVoy47Vw1wacdyEnguVi96PS7jmqDV7jIKxrmE/b25Zgh3kd9D4dccXa8Du3pKmKZicHE
pewhPSELIZ6CAkrzz1L3pu5h0TORv8cRAPMbHV0IT7iTGxG+S8ROoRI2hq7ffDD5yjfkvemZEezN
iCJ7cS16t6sDNsz9QJ+srzfa8KLgKGbUQ8lPYknThKeSS1slEQvQwFe9vthqqllz6CC9Yf8LTJw7
6j0i7gt6xFH2tTHBmJNsgYSTIRJ4wuuZW0cfhB1MuFHcG3oPjdgXq5WinwPUsuic3vO0jjCPy4Bo
NCQzu7CSIc7qp0jiVlvMJTRoiPjCnUri/cb94SP8i38srFWI7K1NAXl8jPRD9s+8TSL725ZUYlRn
kz+kL31gl0bas9aBO7evIbeIiA5qd3yhaBpJlfoaE1g4zdU1PjYGz84rxEUK+tprcBBzgop99DzU
BAcNd9lP3jglx4Ea/LJdu3v+/jkacJPdBFSBoUmLGUYw5LOg/+8hy5epm3gR5BtLIbE1F+QjdeiO
OhLcbdBXV07Yf4nqUPfkafOWQl7hpvADFO7h1BC3hirfsj9WccH+SyYdmps5xt0GWd4Z7ssASipU
ws1+Hw0Jk04Fl20k7qdy0oYoBDtEuz+3dnx0VJhdXfYfZMvWp/D9lOzYLq9FAKSSyIaCkIK0Gt0M
V0OJL/l0In0ks9VsMwSjHl2bviY0IHOxC349VMy6NUrz5AOy0W3r8AS4CpOQeG4NVahpujk3m29g
zNw8uglxWit/oZuY30CAPyQx/FdkrjHUV97/nb2l3APvBS48zKFZAKMg91kVYyYJXTQGNu6fH3aR
o60A8vy88JxzV+4vFL8BYPUZ+ZQQ0lUbfVtcnCPCsUfDlp87FCDAcF+nCdlH/TZtlzf1m5ZxTzNn
2Mf6fJdNAaXUNrhMyuSddC1MJtGdTm9v2/HdvnSUo2k4Y1+0gt3G59ubZ2VxNycj4BT708ND/T9S
dvq05hmBunskiv9oiC+9zJLyRKFfQLGlbwxeLUsZipYb/MGgeLT43uOK7PNYeTFl2s3FXCbow8XG
QQAPOlZSNHke8hshDB46E5h8Ba0WRpqjEqSnYQex3927dgYhBCH5/2XomogUcOW/YbpwDImjbEar
MPGOEvPiqexIcB/mLaZJUsAvC+U8lQsZfim3cygD2rNjcsaY9q6luFHW7NU8vt6a3J9BULycb+0l
RxAOFstsPLoWXyLrm42Bg7HeV3u1jc5IMjuvfG1gNO68LoCexnwPurmbi8WtgCizhifu3TsHkV6T
bScgAa9R/mr0UWx1Vd45X5IMUlgQkQbS2gZHYvUE57YPZxIglk4MwbrY45v+3RLfNQF7WqdIsdBV
1fZuuyr8BrouSYKgNryM6gW653OGUpHPBsB3dtB5Hp6/9KuIq5X6jXEbT+kMkdSm+goHC8MWYwba
vcSNqt7g3wtBFWkMwAQo2xK9qrNrk9Zv5gpvy4zWpLctBBmxjFg/C44JxEsA271ths54Rp0TZLFN
jNXVzd8zKjhqHeGIsNetGNxe6xz49kBD9J0sUnkOP1yj5wrxfQuHTocaBEdkDfT/3ekqUFoibJMx
HOVODrW0UyksaHk1Ish9islLX7h0SqAX0Gjw8PawQAcQ+Gl8mZBQzyLVnjloRrHt4O+TrZb8xhiD
wawBirjzTH3zUmFlV3GnteABtmxhZF2oJt6DyBHJLSouyb3Ym0RKfg2S3nnXVb2/m1V2xKy31KYC
gZwy+u+942yWLRF4wycQcqqjtt5QwpvjAIxspuqavrmRGxx26+MLU26Kil69q6IgbuUIF3d7UEg+
5VKH+CzgGWsq7qfwlVEILHbgeR8GxW0SsZ9srrHvb/mHTOCUYEt2//VU89Ioqphyh/XAQIjxG9mM
XfrayWyZCTmxJ5UbbwWEG4gyc2nRs47B99MsvTXrVRowdTqMbPzM5IP4nVorESj8WVbvOWmqls51
9E9Fc8jZIJR8h9/ioeVV5wY6E47ihawehkD5wSJdy60YRz+KqCmu9KSvi2C+PTPMVRVs+p2c2yOg
DUjMgICN+gEku5DpqEVyASIke1lKWs60hZq6WzcwvRhGS7gjIQc8Oxl75gfc+zxMa/Mw5x88KS5/
5pDPN/9kTJjuhMLH/MhYFTnORWUC8weni4isxjuwpR2trTAJECWJzvseJJkly2ioq6nutMCfojEK
UNX1mS551zbsdp9Sv4hKGHfpNJl4C6rxr5MDkN1mCNr2Plo/yMvvMOOTy9TjMDGVzFYGkBjBs/qp
vVqQgH8Bpidpm6YC0jspiAo5d4RaPEfICvM+XWlipgQQQZhm1O1pf5Cp0W3FIH95dCpqlYX1Z6Ui
yICO8j5uib0XphMvd87ePuXIF1D2fU7SkpdkYftTWz6b4txV0BfhUP8TpU4F3kXFGXd+1O1D0YEF
PC18CBTaREXKmgPZVY+khGp8Z2qN/YaRtKiNsTPs19HaT06AgL5Kj5bXKJ+zU9ibdsmeOWg5Gppf
a80nmUe0y/m+eP/hIGyscn7Uwykox41bzIwkbX4UkdgMGnD0wiTzcUoL2st7WNdHQT9K+h6+fR2B
ME5fw4G0/kJDSQ0eBfQHPSX/qYZUeFtuCIQNcFAtFR3vMWk8V/qIs4OklGCMSPWuPxUVW9AIfHwH
sdE84Se+JHA9PXGRCEi3Tk2IgdNrfa3XdZwlsziO3t8A1avmJauLduP+EGz7OwXsUc+4SHy4dV5m
X/tUKgkXlpFl7zA/TttTgZ8WZEuVFuhwreBza5OO9hITMjIqQcMHhPMlitYfrVR+PqKBpJLNStjf
jEBHlkpjfuYGK11hDbuGKTVZpK73//9Ogfo69jMFJswEpSx7lRUQh/F0oWbV7jvQXW964o2gWaaG
pJxfCJ5wCOu0Hl+pWqf0QO9zUI/G2RJ9lBdoGszNtxQojxp0A/z7MofZ+l0GiCcs1SN+QOJV/nC/
kkcdkVXrabl7xGDnMAPPfQY7LuFjAsRvzNxKaRH35pV8TSM+jwTp32uYbF9HubEvXqfCgG4ggtJs
uRbUMdCBVHHfhwieWitNjItWe/Xo9Uvm6fvbvShupMUg5lMCQ/TAZ4pn0Q6j2CJfYJdFQY/Dvrqa
exXEGNW0K9Q2mWjbDbxGvpj/jt8ASrnQKsTVN4PrXASWOLafMvNoMK/0BABKAOwsLJeWNCB3kxaJ
+7W9a0sgRXM9OMZs2NA167msBYLXrij/sWwBaUlonjwbvTNyrR9Bp4pmyBmEcQtydo6lfuDST6Ji
Y+Oortp/jJcCny4awxxbNZVYRyE9oVctGzCqNJ/CfEihIwaccyk3Fgq+TpM3ByC7kJP+d8HYyw8k
Rq6LcQ1I1FKEu+th3bc0jxpLgR67DbRyaa0sOaQDs5p5adVZvffOx/nbCR2AijIX0dn4BzJLwfTd
1dPyu5P4cxnxGli0SF0V+O7tx8n9nDd4GC8C+WYDgz82iaWoZ9AKEOjR6cZ7dlzdZDlGaBniYjCv
PGeKa1y8x5zRLW+Ls0+fEexOzqbIeWoOxGXXNI21pg9yks1awQ5H3ReRG8TyXOuAqS8KhCWBF+7P
fIbqYyflT3EPvWpPe+Lxk8v+PHNVZR5BmXwk2IdArFG3dFX5VzwOYziKqR5G92tZmogjDxg6GBQ8
qbKmlB/TtmQ/tlnBLHdrasEItrPrMqbdEM3+aWm86CzslrOH4gXNBHkdG5HxzpBt1e3ujiiBZ5ta
5vM4KG/sbbgufxr3Y1Ag805tpXyl6/IUtNlBpsnCcxl2yHdWveYPIJiIWr78jBYbL+c2nVDK4oBd
YCIZXBo1aB/uU2/9+TveF3j9lEnlFlhk1k4hzTjPn1Jy890CgIiFdwUWpZZirkMH1Kezx5FWQEEv
z++AvBUAPCbXvgPnfkLQAFtFk101/qN1t57NHBAS6wXk3t7r9QzxeWsmhs5scE7gFVYkHsjJRBTP
G+E1UyOSiHIVRdpOK3v5iVLCZ+8ZW3mlmcketJjOiiWW4BpEcgQbK0iLkpgt71oOUQBpmzYctOdj
HU17TGeq5CAwKS8mEB3ufxDzhA85s/zUFDrBlX0eXx6GgsEkaSSRjdL75UExMutt4jonMEduyihy
g+8LMB671UM01NyYJEsheYEMLIEUf9W5zlLMyWTOqA0t34BJIi9IUtElHYWci9jsVHBP2cG8PnDy
RLGm/ANe1QUjCpbpAx/7mJQDtKtc2V9WPQL2oOHAvkA/u906K7Aw6UmyDTgpKqOJQlLPGE9882yr
5xQp09ZWTS5K/jWUD1lkcuyA0IFFDqHqOZo4aa8hFPLuz3szn8140u4x5e7FICAh+3mZMAoVX9/r
M64tdhO8vcoVKMnlS+0H1/E8agAvZU9emgtKb84ThEI/ZrV/i9BIw2RyZO3Y+o2zVR6bTcIgCHgG
pyq/s9vc7XT2De+pUBXrACiVU/ak7MgsiUGfZKDkbvqTow9kcfUMZP+/lJeIYQxRvZcw6tttsDpt
RRKSDQyj89lCAZBF0qgmr7ZmMSezsfJ9BJ6iMLXYBJbYzV34aSaFQ+Uk8c4g+U0qxW4YFURbvNMi
LqMowenx22ErFyjbBfZJGEmIjtwYIZStNvxgRF3Ij295/TUNKpBzHfjCFlDUgoWwc4TwUSY/h7qf
CDv9srca6ZFjIWfPGz+SNZFfSaPjuZcSj17Whlwlv7Us8tr3mlPhrQ8DM3xsrGH9DsZE0GPHqg/0
vrCy932PYKt+zfQ5L5Rvpy0CY1d99NruJaPhkJ4qj+EJR6XxzznXMYasNJ9CgArRPvijet1mN+mV
F/azBrZ4Mp4re5KCG/VQSanUYJVZ3v2P0f2VN6zrbAnIDjkeRK7mHZIO0RuA5YS5sJt0mxgsBGTb
nRQcd9+gudVOZ4k1ghipbSGTjf2rNFYo3XiwKNzPOsV0D/e8qWi71SyAnu/3EPeVh0TY5XXhJ3eo
pF+/bDSAW4jPaKs4KFdJWxPoNErpv9UUnDMi54HGWfbhz7bhbbURsatpxEGslxro6VhoAdWQMs0w
0HgO51Uy1vAD8HDivChpD0BluKJyeMDfxphoFxElS20RZziFx8A0lSwmMxNogmFOlBaqc6rW8Jin
Si5ZLvX1LzpPjcT7bklrA+qChHe+4OSEsRKQ047yJzrg9YTsDcj5gwKr/u2tde/7Vg5WJFrm5iG2
Wo6Bbkwbfu2AAII7+uOzl/jPrIK/5YmxfM9NaLMmrR250e+6PODZAw6VjB0f1COQjmDvMuO7/2KV
0iZymxzyVB8YAtBlT9vz6Xapeb81Q4x5TCmY391Ip2xPzuHr4+5+OPZ1GQdB5KLjLnVyfngIhMbM
yAiVvj0M61PiKTy/rMZb9CUWFocUhJnfmgyyNbwxISh9GXCqSCFssHhA3vb3hraquFYahXUtMCXD
iYCrMCcXkEckyxntyHUg6WDBQm8qrYsbV5PN4Q5cJyTm/vHgaV1KmPqxyigczx3bpQBJd5i+KMD5
H1Uu6l4HThrOrMRkkBEA1f7KJhzNhpZ+wpr76LLgTAFc+cv2euInbp0XU84um/xj2d4ZxBHDMdyT
pIpyM88al6sMSQf9AZC0JSs4yGkj5wj71IE8wlrIaOMW+VscnZXfOVRUQM/Km4diat54Tuh/pA3e
bdRY7rS6XhzdAHBGZ4vQCCMeZTW5AbulmMeyqSHxoJzkVT1DZ4vAHAkQ9aQ71IWUn7qVWotp1UeJ
N9GYrAFmICCshh4gASqNmS1PWtJznWTCL7j3DmI6T6zn1BkntWuydL0BrwZUKdHH0acOEnywmlVJ
PHg12iWBOVIH5+S4hFHEPN9WtKSt/XDK+a9iH7ZoSG8IIT68Xu35UmSv4KwOwTXJPBgAoT+QgXtz
itmrAAF6nFdDG5qGHZeTFZSxtX5IDk5UKxbtHBfH44JXU6IRdXF3lVQGRh/IvDeZlWdGIi67WscG
Xl92UWCwYXJWf+m3+o3EFxCsqTrNzLebKcx0VN5IGccfTgl7/mPeKUA6kCSHGG6nKwds0djnuYh2
N+K7+sWlCRsTkpPyO6fUQyKBF1tnLxhZtzq3tmWOxXO0rAQpaCO0qavoxUMpXJwbaxE1g3xZJy8O
3iKTJ+am2Q7sfWuioSh4SDpQ1PTNin45YOYT+vYeFGNivuUWpJiaxGY2QDcctTFkorTgqvkQ/R7v
w6eB0EcCabks5OaNV4g437ILTIIXGHPPPAUHQcn6itzt93C6Ul3stMqUx1A3V6Z73b5JjnK4IEA3
PHJRJ+Vfdzk5gnokEtag5Vu20TWZhK6u1Jm2jT5/lt+a2h33lIVJNSP2DksD9ZfjIuXMWyCUk1g7
dBE+8ayP2oCA2mJVQ7UZqcJz8fs32sDvoJ5sGT8mTtEKTGVl8Q56+eIkVcvl7PvwvNHQo/F7zGUM
PvajGB/dTv7UcLi4MBELyiwYhpNOZG/9KRC3ZZ63jQJPJdgYKRqahQ93BoAACWwcCraFdSlwhhi5
FSxOQvR1jT1C1ALO1tnExD3w0BTEX20XhUGouL4TUyOEvfY0tqnO9Sq+4KiVGKsiryj+QGs/EqyJ
7wI5NMvNoQ8YF8tBQEBszTCeWMJT0uCBudTNAMU36qTyvo9o6+7oww95v5gIZ95VwmX3QSQ61mcM
8o+LhFjI+DfI+C/g6J4lVAssk/slu5q9x/VYCDBoDPlLo9H21hif/YvHg6jpeVrr9M8i6SvMQCRK
oJJn3ck1eTtYjlWpwP8PCgr2KWjAsqTidZOq5HMzSpmYQXJM+7V9CtEAz5BM1VHvB817TO7yBK/O
EuNR2/Vbu7q283ZIHF02eu3dp7HFPZ3wAzUYUN6Ep07EX3SMx79eRniFgzcWRbW9Cf2N0ZjNbzyu
/dWPMwi1Wvx7zrlzND2mT2/PHyTroOh6fbCTFfSGc/ccEWgQwCP3jX1mWvB6w4lGTlfly7DGToUE
sJWkzV83oZiSsczRrNG679ESeXrB4H4YLox4nfWphYNmGiZD2IzpcfponqM+3DkCL3GSW2UyHAel
zXN0Qb+7p5iohnXD1gHw95p32gzb59gNoKBKUVpGlSebrpLouHTm+edih7rZfTAFtX8C5kG0PfGk
0MArlNmQQ8caPb3wddcFDUotSexp2gSswi/uUhcP5HI2pr563OZx1Kz4kft9TRQxTTITXuGFKBcw
cOqUSfleimH5Hnf1PSL3QTTa10+5JHEa8Wddpk5S40AYE40warTTyPJHmQM6krJUAE0LP6IQPo6k
OLtuSzJETtW6RJ+E92c7ByCUHuIYMcka2NCC+tIV8I28A96NRHIbf3ap/wofmeHwIYzVY2fOQHFU
EyZ05z0RiqBTFo/tVpkNYrayoikH8whW9SXW96ZZC4C7Dl0CDJXF6xCrwBt71UcSersa46H2D8Mi
RSaCGCysWeRuGehOfy/ltPOdevCFUUUHqGcEJPxMgzROpQydMFJkgipZaK9yuHDa8N758mKEoqjL
eznxeg+Bre5AnqlvLZdTQ1Pa9JOMqgwKWaaV4Z5asipgr6xRfDzUIC8knKnU6v26/g3SdBBtdMdF
lbdrkSHMNMMpVLWMHxi1dqmEAL9ghWrvVxcs2uXCD5mLQTVjmYGnBg5aMDAfqGzqpIPHjgBkzD0B
FVzYG64NDg/GAU/NMnMaJDvyGXBNu385VTrAYGy1nHi+GDoOMeqfdlt+tECyMlkr1B1tHXyzCenw
PS0M48jC1qhn026CBORCIBk2gMfiUs0YVPNEOenFO6nCV4GP0RcdJju/4nQY3wyDxoXy26y7qXmI
7aWGDN4Ns67vqcAgS/AOxeOjiQeHcF2LBBLnnOY3zBXtzFEKfJpYrXMj1l327lL0X4PwBEk3j9YP
5DDZ8usii0f+KePAOzxi+3dzLajg6z7xYRQa5ml7qzLi4y4crCf8Y6+G73erVt5wP0NkuQo6hQU6
YBL90s2weZ4eEenSTB6vPNNASjy/Azjz+0F6IU/YpUQrZVt9cBT5MBDTU0pqtEomnLj8dHpK5OJe
zOU7ZA0JwAAw+9Yf+yz7w9gMTfOHkPD22gI2Cy5oLL6NbWL07MZxq+nWlJjhBeSjosXiA+IKlvpH
PqoLu1w8AWY9pyLG1JZRigDPPfWwVdgIZyGhi+vtpija1B/8vBjfJzx9wpcLZcCJ/9LvrRhFUHZE
UkoGZHFhBEhFSnaGjVeNYb1WUrTBdafSx0kj+8XEf1lBQgoCsfmTri4465M8P3i22vSiPojMpaSt
REsDtwmfZQZ2lLTIcxMuym5Xfaj+KK0PEbkEdKEGOJ31eroW0kUgtCHhEJyhhu0CgJcn8BUOLgEc
prLax6D0D5zen9JBy+oCeAnz1VMGkDAZq3dusougOcwQiDKsnNL8t1KjMkuV/g8SUwJFLAslLhGl
UxVX1TfYLDRSIqY9c4CjfmbvxiJE4QLj2o/kts0I0pJLtE34BzMa4QvjF/lOmuKlfbd1+A4m98hb
fl7tAqZw02tqszvT7mkpcdKt3SJBCrblfi5KBcz6yI36AmiCcZorQcbBdt555e5yJZFxX2BcA6G0
nIvx+SEKDS9Cae3CUcWxluHmJ+WR0KB3I5LDdRdTwnbjaBck25jP6qa4bJDoOdXe9mIs8llyUso/
XCXWr7gFyxE2yWzoL9vGSXgbw2Jnfc+EyX74JLEKgvicZ6fPxn0DN53/6DJBMGOFVAz/gamYTaUu
Pz2bVNkgFdo0LBtSbaiCml3WekCZ1qDQ5u5NTr837SO/oaYhXxs2sYqG925FHoPYnr4qrwRwO+AU
0By98BzZ/90SDecw84wELbIjC9p6zXh7tJ37/4V541PZi6G0WgQNj8WJQ3lC+qXCamc+aWtT4Kzs
e7OG3feiHDOapj6idGJxux6ZIPrBcDuyFu9Gz7RUQ7ZM9RdfGrmYim+NljrknwvY4LQM11y4Cva4
hMTiepEKXq511XeR3CWOhIWOwN7/wOodKRGDPgyeg7D70IyFwS61IK8R2ODieWxZaJc/K26T90sg
odbZ5aql3jw5yodLr9xz+58O9Y1goMf4dNwWvO5f0iHt8N5J8P0eEt9ZfK+lnUY5Ud8AV42cwN64
SKYTWmi1ompy2AmbVGfdb5DKL/tyiBnMuDk1nganbsWUwuOwO9qBp0aU2V0ATGy++FgstlYR/U9p
7LF+KCGsD+KE4Up/HLnRRnYzDMwHkF2W7lBQesyBi9qE+LhYLbOjotn0Ah7S1pkrENW4OfMxPZqG
MckqJsEm2lH4OIGXvZBu4ja2VKGl9j7LPQECYwW6gWoZBt3JnGhmTAFZne53ehjRubkADFGUARcH
o2iGN1TLWJvp+94N1zMmEaiyisKewluEAofK5MfDt+H/As26PudFs6agtN7WDlbgRFhZiI6jwakv
yYbQyK4Uy/hZtDLfrE6FKjHHG/pPSev54G4I8nDGfZgiQZgThTOSFCMBRN+1iiH/94tjlI2/3WHH
W6HDJgdKNP7JKqiM2Mbw5Vr7BdTwgwu46qoJabQwRDltynAj2PDAHdldAhdYVDfxU6WRf6hXnZVH
DJHspNsFsorm31Y/H0rfdZdwNDkmPKSsETy8SJjk+JWPcKNOrw3+eIK2DBbonGsRqLr47nK17Grv
aD7zLro3a7jIVMzm70kg8CnJMytqAMEPazy/DFxDvrHlfq1+nTdFlJw6F4rk0ApKcYWAngaLlNlU
0KqGlWxCfLy9FA7CRZteLvczCqhMyQHBIQVhRHIpd4vr8n/U5y5U5K4iq7udX1+DXGfL95TbPYb5
6lZNhivtzNQe8Td4f6vVy5AUp/3fKVRRxi1bNMPv99cHtOMhzbGIFI25zJQXNCL5pugT5LmnVVzz
CYAo84AhMzSMQiw+RM/EN6pi3b+izYORSAFM47Grr7QAWO3o88vaCHYCq1RTi1qn2TuQQ348Ld1r
3xewNLdA93RgRo4Ev9gTcSQ80YB/iaXq/bBZTjMe/N5g6JAt+UUzQNqZnKcTWcwizTDL/TglxoXH
aJw9E31GfOvny64M+j7s6VgT2vxCAlC+i1/XZ0qVlP0RlDL/gRTxj+FkISlWLM+0p7sgrDmZIgqe
pdXP2dmht/M1TWXIeR11C0AOXayATHTJ0Vyd59TpoJ7V/BUEnmiuZUFXUUYLqGpFcOH+1GZWKIwl
umSaQa5Tbex9DkiiZfk6evXSZ8nGXtBY0lSsqtABh9z4+n89N6KNwFy9MLA/7sj/9bhNoXXA3GeT
zQ8YN7nvNVFFFm0G5Z0Jx+oXNlpUelT4utpLoJk/Lq6DEp3ZWTUCZFBtuR21cFWm5XpydSDn0NIj
SknDwtpd7oZ+mHHgjM6kpNYWV+UVrZWeiWIs0YTLCiOGV7bgiyGlOAFG7cyERK8mkIpcopA3Vn91
hn+PV2y02nUunJbOb/4mQIBaX3sovGPFwzwknOzn5nMbVbMF+0fUoHH07WZjhXetHMPxn71KEtdv
tdN5kJugBYyMYcBkYkYnp+IN1/SwvgdRO7SgFXBKuS6OFvvFRM4KIlpoRYsXvcnQ3c8i5IRsxG9F
egrZfdMrGIBZ2QFIxduME7WwKyZ4lE3hdk7h/8Yk81cvr63d1EStik6AIN7CITWZOGhYpmoVEEZp
VVQrLeLheUB9rHzafID1Gx2rh8tM4dW6Zha787Ip5WYAxfDfpvoptuSBbunqNQGVwFxzoNlX8v0b
b//RiLgg1MzWLZRYKdV44Q5AfWzR6WdRnXd2mpK7yECwjqFjskj+IisgKpJr8BoSh4uqdrmJfYUa
yGqvd3L4PLdoA6UUgcoVPbC2EYKQKqbxDOT5O6m7pgO/eK4g1B64rJUfzUmBpMRSDmnY0wNPEs1d
Kd5G7oQPnUYW+nc5S/AUTz4Pv3WAyyXdyxtrhaqWzraP9n/8L8znp9DvMGxCRiDdHL2AaL2UoUix
hdYoBW/Z2L8peNbdRzHcoiTgpyf4RnkBAcsZdEOhnz5jjKG2u6bsXLX+rh57Hjm+0FESQutg4ObK
xw8JJI0uZrGpyTGuco+hc0eHLd9Gyd5uRX7KnM4mtkGkD8inqw9ZXjtK1WonnyUBSZycLM57clYj
+YvHOieD6tN0m/U6ZEQztrnPSU441gbDKtW0faVsugXGd2nwt7nlOmu4BTYIdaF7H3TZX9mahx9W
f11raPo7XZ79IizKNq/NJAJXBYZJYj5CpZJVDUeIEBXWut33GbqgshIF6Nq85CozQ8U1qdimW3Jl
X4d/n3cszDcUB3l+XT6phOZ1xxJvlw25F8HTK6Zbi77HdHbQkmM6xjzf88agDgizdn+LkdorrO4Y
Q0tSyHb6ndtmtuZTV4KazKlmF2GZ4fcRkoMdDHdmyR00BP3QZhJh9ikdD+sj8bmE4voLaAO3enOD
GinGK6YPZ8o9quZS5+D1ZxgKJWCNZWasWNxKYSrsTXYYsaptp3gjD6bfl1VtNk/TzqkWAtaMOt0D
181le2IX1c60Z2jc3KJSNdSFSgAE3YvAXuRuaRATonXIKjWafn4Wqp3L5V0TNypvQmRIXR2Ae9HN
HlQHXMHHM6uHvtYAiaMj0TXUP/K7L4JLuOVuMX2l0/RAon2UH0WD2L/EfpZQjBiBegu2hCLbLHcm
yOi/x/jEmaBmDdl5+oUGv9AV9d6TGie+SsWrl+7q8KgNBrtQUpleAcpA/rbbQvhLjUlWPbPiIMr6
vrfPTonl6dDWJIvO6zesMZAj9R1PsPmCSsWEDTCgdL94GyDsfiUbveODdi+HjtSlRxLAvuVcMVD6
hvgDe06UA7VbHdMcNXVYYVl3u1yaFVdCJK7DOg91XlloifuN3V+h+vZYXL5Hpw2/gw9TjqBAPX+d
yPpr+mWTmuaWBnKpbBk6UWdZD/EDX2a5ynymEo+NeUaE740cMSIjiEQWUb9UqSOlWOdwmMprjrHX
ClqMTpNxb/6nyn85c+gTUOtYbsQIabGEn9Ke582q4AFfqLm0gCwwFwXSYA9n0xbugxz95P50D+zp
bPymsiLrBwHT74F/jPFYKFTxs7Jh2Y7jBdlcIAp8YsFi5SSp3H34Oa7IE4F1QQvSR64UV10G7Fx9
z7fRsDY8yxdDQ+duW67JNPNhiNbPs/2GOU1+LvGYV9zeJCXYjdd7kLZVGPan5tjVjQEEsHvfyUxP
S4MfJBrqsJrMZgDGbzWbk1hqM0n1iMhHW+V6RHf6WqbGW6gMRpRSK/Dkajy24PNV1Xbq0LAOlSAT
H+87f1zLlaSShaQOS52Y2hmznF82i9W0cwFB3pSLkC6v3DtvdPZhClLf9wIaZLED7rmdC13ND3jc
OpM9fgG2IQeU8AVDBYHm90lk5ui7fRuTav62cc92LsisJ/aYrZxDOoituY55EFKh4MoUhwgUgdri
GX2zdHPfkC4E0u8F3xxgH+Srq5zRKg4lVZ1CQZ291+Uh69WJtD4WIoDkYMfBeVOhZ7O9rUcBCbOD
hvAUd9jN7q1L4msO3d84eQhMk36WLoa/ADBDRTBvK8VgKMSnFpuI4bSB0y52vH9YLzcaCd5g1Jqc
FTnjruMMKQdcYUAsrU6XG6E+6b1sBzAvpY6jv6lSdnjdw3oao7OVmwIcdYGVn/VPc8cGXFIThdEL
5QDTrFOgIhAJURxB2xKUFlrCj89Sj0iKdMwJOWSYkHl0h2VjT7b0MVpj5ucFsuM+oaXXy1Uxo3SG
tT/PZa2wJTDVfPQtbHZkUt32iyy7mSS31SQoJ59tozmL8pmlAktVHAK60JwyFm/TagLijMAxhBhw
AYSNHKAdLcFYM8tibRo/xJrBP+oq/d/JAHl3N+yOl3nlpHMCrAsftKt6N/+X4l+WAjf7MRwxOs0g
9oIeRY7EXkqTe1kUrosPqXsIPCw1fDkgVcg79qMGEUP4motaIMM2buIfXQZwN2SjcfFYTa0P1vU+
6V4olH4RVmq7ObBca6AGvu/bH02waWMrZi+Ga/Qkga6JMLYyfoBEbmajdQ0GK6HAY8jsMeU7Kuu3
neS10YQtHFoDzkAq6cxPn2gVMz/AEJb/FhDzn0NDAzaM8N9ipBsOTQvKmRCrXqjZPW+1lRcPEWu0
JzpVYBn/xInuvbER6jd22OdAHVEferWSUxDrnUUSNORBt63jE+xpiVCvacB2hNbVgBrN2fjWCrEd
PxqOoY+fs0aqsujwKRgAH+KuDPTLzFq94G7f2ohU92LgNJOlHbsXS792mKUgrJAyPiEW8lWr7cZL
d0w+2CJbMaxhswSL7cFOn6norzA5lRIjSvcxTUApNlPklrMwm15CX6ZMeNtPezVrq87ANCjnFPHa
TxETbjaOIkyAwlo9C/TOllzl6fTpRNddlVmKE0Uu5s67zjH1tmqzBONW7VwKTtFe3A9Wpr8H/JxO
FPKEOaJWSz+8H2z3J7lhMiiflSLlSwSfi6amjnYvcJUt1VL7YQkqJ2w3UjO1i8eZl+W58flOQ/EA
nBjFl4Kx5I2oWZI+Q7HZhr53pSwbdpJTt+BuG3ufjjAHREU7NPgC79Er/cIYCH/dpOOzglBBRZZ/
vVRW/SXXtslV53x0/Oeld6QxnYHc965HSBY6wZK3ggyN9GsPj9iL6j2fLitMBZzD/413r4WYD7mh
YMW70wPWWEu+s0BXHK5FLacSnt+WHCfOuUjDfygecgD8llbHLzrbVMJvUYFdIxy3Ji7BE0aHu7Lb
8vy0AkvOplIMssOuDsGmgNBOAfrYOqCSF3wi/gux+cSjU5YafdzIHWbRuEA5Uq6D+3/CsNeBGLaE
3ow4dQAUIH+c3lCoYpqsv4k+Pa2aMMrhfl/XRGMyxO3HFfxyznB3iDjnd+1jj8/JcesakqKnQD2V
Eu0jdk+jkt64S6EM/Ix+13+NS0EgXAOYCGW/h/z0ZxAzIEsnEH/oMsJCsJqr3zVNepOSaa/aPOuV
4iN+msRVAor3XlJIcV2wmrE05RvD5o+3Jk9QbFk/OUHD+pEvo+C1zVf7pcYypozIZL8EOpUoMjkz
4qzCEW7T5DnZcuAE+/YyGHEd+QkGyyvGtHnPLadILaBvfauQhztXgK6XSqmLbIc7wfWVdWL3h02q
ffjyvDyzpIYyyGQ9GhfFc78DXAHg0wp3rbwXygJ/cNERKMJXnpBU4IFquKlJBgfjRg5boHnkmkCx
jElvZGMWm7PZ1EngdGiN3pzpwCJLPKulh+Jgnr+6Fpngf+Y2j0Jv1a4CB4lHNqQDYJcHh7hWLSH0
uXexu4DkspLB+Ar3+6pd2nv1zejT8iUgqDwFDhnn9L4gSPpRERomnIfy577muz0CzEKcNEpBj2Z6
bGHD4P+0J3E7eCFfpFGkq0VC3GHwLg+bo69TzvycpuCu9FDpOevQdFt3Ly4Ye8EP7Of3s/Rv7U3l
OTmQzv7tcV3GQeB0b01KKVpJY4aeMh2x+7LJGedKz1mw2KRG7fP9wws27bfBECfaeBETL6STo5VQ
F6TEyV49w1UMAZuVNJ2IuHXN7T2E3POGRXAn/x1Fdg7j355Nrna29ssSfqA2EFqu48PZr5MphSsi
xU/vmuBmUUgi6LHIpfwQ7HEcj6TRiDznSYb2BS44YRvnLc41zic0HRaMh/+cWIDJkdkdAEG89b8O
XiKge49l+trDZHWKVnpCeiZsbzTgFGBQKGPEadXjAT4zKeon7Dp2XbyXKGrmpkNL8LwKQlpCJpVT
K4klk9QsIkijmWS+xFVmUA6XGGRFnL1dWqV54mnwmSRgS3IIpy3ApbUYqc4cAcyecIiG0BqB0t53
HUEyjEl/7qk7rtMDSiQn5L4zfwNhTn2OPpwyP8fMja8NcboMRphpaMt/jMqNWfkQihR0RPuof7f5
yThX94ZsaS1CjALp3mLHg2rlHVOEbbh4hRHo01Bktl0A1i+NLUWYKReVfHltHuf6IhFGH7n+kzvg
1u1HvEt+yY4GDROQe2EIgD5Fxdvw1zu1de9rR8tY4/Xz6kjs5k4cqS6VzZw2nLDXwfzasnot463P
5brzAcbAiQa8OjKPyJLo1eTeBfAttqtpQisr9ns75gQSU0v3rz4bAFadQ7/8TlhfhipB6HmZF2Tp
A4EkFxEbJVI/uB3ZUxeCTqBoU08H82wulU5wbyPlxk3gaoBi6rwE68LZx3f6T5kSv5ZhWEIYeJOA
PzAQMB9kZ6NFhp/xEkHOhWuoq4wiYCydyLS5OZ3QrKNq0i2+5kcFsZ9v3kOjz9QzTIQMIXEVvjdi
TlsoUC5UaGSuo8C8FgubZulkKUZWIArLzZCYrkz4q8HsT4HTL2AiIbxjFaZcV29pgbhY7ohxOySt
8g+0SZR9oPHelap53EL3uh8RoEvDwQPpZy7CD15OvFJ7RSCe8W2v4/+SWL1Q915P3T2UWmqS3zS/
aPNvfzBLRKv8URl/5aHB/O/XTusl5qTlennfAvsspU6/BiTNdUiUPup3RA2QZeA6gEPmcQzu1/9y
fbBZ0sK90r6fq8MR1YL6XgC3TBvFGCdYzdyNEiIs/4qwT2La5WUYtjgDQcLHZl7GzbAErSC5FnIx
hY5CVLBv6v9MH8z3fhw6PEMN34Pus0RDYHw/xzydWSRCEBJMkjOa6CxBKhVUCG+jdRpjZ6OW9lBT
PjqDA0AlNPozKJaUcMAQbQrmJ230zqIfuryLPGHcYJ9Bjg7DVJkhuFjyt8iSYipMyMsbla2PzN7h
nkGtgNp6P3/3v3cz9Uw2Uw7LBO2sxJkB/8tZW9bx23k1QOtITgGqfypcdh9lvbix35gNc9SXOspy
9JwBBx9TqUSsDvcIggmD2VBtaObJeChaBDBLDsaikFmgwgcZ4/yRMe8Su4YaBkt3TJo3F6konnH+
qeRCPqwZ6m4eSdbVjr+VONHBT6s5RsRvw+n1WFhwGrJim1at2fm8hviMAZdFJ63km8mcv0IzE9ZU
ItKU1GxVnLbvOC6d8kkPF4SCCdoA1kNRYcnA+bZPcGplo3lpRUjKaSeej9iUw16MwsItYQHuUtoB
EzjsItpJrVtckSrBniYd+QO9zyzL/tylDGARFJJ6qv75sIceGWKayiKc2eyNEn6tHAbGwSp6eIy7
fvBRZhJh6OuG6hhrVAooMtW+MPdBC55ncnbah77K32/qnvWMIUn+5FQQj3kpAq821coXD+HCbu2k
rY0WTA4xVDv/97L9Mv5/+/wsJVQ8bCl0V96Qs4ByorUs2egRDuMVav/L/hqBggcTaNMLYsfaGi2G
dNX9cop91V4lmCOmM04ta2D2bSBB9mKyIJcD4bablg1tOGoySdCm9b5u5zdR3BkoQK2F0Nm+FscH
rEyfEm8si2P8C/YvynF/3mUeBGVeF+PHCnvfA/fLMIvkZuoo5OYES+XtVdHPWf2KFvvhYi6TKIAm
Cki1Ex39LeWG5aTsaUgwqEBFblAnXlhWLjvvIyr0G19USJjXqT2mvJW/oZSpb1GxB3ZXjSaT6jLN
f5VCZLhCwyk0ASOVmI2dfO5zs14cTDcG+xMK9f+Zuj7WcjgzY71VdMcPyeshQtwK7ZCfCVoROMYY
lQj/YsqKXmZ/78MxNPB6GiIKpWVefGVS4o0LFKK6hqjg++TG2eNf8MTBAEV7fBhny9U1h3eP1XNU
7NkbM5SrSXekwVi9UC6ufsuYSSg2VxXf+OQUgU8kIk1qXoTaX+6IwFKNhD0Z85vhBBbBMubo3u7E
waAf+SP5f8Lwb/VcYPHB4X93u+kxmI+XSDfYArs/PX0cwL4Pqjh1WsemG04/KmJsyWF8d9Uyn//6
qAgmUlwnQBwr+Vog3BxcuTlTWTb0+togzQDymMomCmxNX/0FtUdkMxFlT8Gz0IrHwUYjyAdTWELG
N40ySN+0v4aPnXaydynKIuk9wMiMOVxti4E8giwnIcDkb1Iyt59uqKNzOU39bBLZUWnv0OiiYln9
P+X7HOU3DkFIe+0YQHZdOPydAIrBgNDQFa7HDRAUUcF1wQUKtnR0OB2zzkHT3zhyMKccAC69zrQI
P13CQJcnD1WM4QscsOl/k+cLCd+sara0dLkOtl6AiePNIQyGYRTWsWtMOjxOql3O84r4A9iH56tC
0Q3GLZiIj+fnKC90JHxU8A8zlYqsVY9wxoUxeTgHN9tKp+djs2iEAkMY+h2OyzNStLADG6HdolW2
MPv+fw4KQ+fOTJp10aZaLDCkwo1icQNU8LIK8PNjAyqdhvKskUzMtw5hu5aX4v6mSzWbNMbDn7mn
GsNTWaVH8N8NoD/kbneZWEAQBPY9YLd2vNgKkkHpHomvRwmVVkI5y1r/JVVwIqiinkLsCbV+PKVE
a+Z9IhAyFmRWiTw8uoDeMerUCc0Zj5W8OKEm4IkRWpiDoPwh9b6WHUwQu7CGeCyuu/dBoRsib5RJ
XQreFtGv2pVV5GKPwCd94JstU9tGfjR+yC1Oi5wM+3o+tpyzHunbAkWbisoqCCXGMJtrxM8Ih6Ak
kzC0z4jUTlpiOYR3eDNQFj9P6ofoPH8o2mfumRKdgBREhTUjkKAHXzZ70RYtRCzdWj6SK9BzF3m7
YuZYjLymLphUSfZL1XXqUgPKFeNEZA/LjDJ9dFJEJUY3d8FDTqtEFBLooCNwH+fTVXVzwXBS6m+x
3mGWwxJ6qzXivzyaE0IlccMzr5n5ca2AXzO0VH30o8q1DN+nUB/s2i/RVIcVi0+RF5yXef0aX+UM
VRL9D/yk+lEqajRmtFr+V8UbQqoPLSrpmVex85lIe9oV4yKB5o4MH150pQMfS1tjRqydBkGH7NT3
bbxU/xj66FIykKS5ms09rJNkJWdq1Ygoa2C2YDgbXWGRYJ29JwPrqsaOKEQfvLl92oXMJquBL0cB
soHkwln/CfETTpOyAxpoCBVBltf13Vuk5+T7XkK4uO6YCLWOiovKN3EgWEHOcLBnkD6eghUqc78x
/D4FKCQv9oHeQtBH4lAi/0ci6H603x18WpYqccmxNFDyvMdCkAN5GsVoDmHdhxJFAfjmY8QGt/08
Wc8Y05IAO6tQUXS52+5MrT/70lhtPdkZyRcZeOryLENNIlttGDxgIaF+vqaXnUNcZSMrnXcRqhbM
MOV9XpbdYaqDv7YhvBCo7RKdws0zmgYiM7YAZiH5Q0y5ttceGa9/yMTvGMCcu5aNhjipGhm2C+Ao
tjfy8xShOaK+sI0JPxUafQTrD8Aie4Pc5c+N6nSNYl4qGHij8wasjZtTPP2b8D1wkZ622+HsGZ9K
1U1Ot01U3HLqwSBELpY91DLeVgmNpSroiQOMS5r3RwS1xPARqFfvklidxNFKGsicFblShP+ud8ZG
rW5liKAtVUKRWp1sqbHMvZlTVNoDDQxx8lQVphynEhuWznyTMXmyd309DR9LA1AH1zaPyQO7jyhm
MnOM4s/Y3uI3h0lZgRD4k7/kuVFUS1OG+MZ4YpBxm4DcnA8KpYy/KRPISqw6znNR3qVUsR/GudpV
hK5S8IYXU9Fmo+8u66sTQZFcaMrCDj1bvtbr+kPVoQl3dkPf2kRmTgLesfcYUw9UBp2lMcUnCaSr
2Il+7wPiGL8MXed4ZrmQN+hZNl/RDie7twdH6fefNQqQ0aaU1myfpf82SzWCbzkAhstwSHXgK9tP
Y92cl9bBgILS2p3jXRreVZLRsb9Dz1VhBwB5CdoYjreB/SBip7WkGA529hQ25JFMZ6SkhaQcxlj1
odkB8tm8AryOOAQ38hSSMQ46b/VTFgAqMJeWr32oq95JyBYPCCG0BI/mgFP+fLvyRuHDpBnyti6C
aOYzI86DOc2al+70Y6HWx93aUqYMYHPrNF/zc3MLqqStIzuT3yBiEuFPiT/y9V4JrK90WjhgmJjN
qSNpNpVjwGvbpO0ZgLrc2EtL05CIDJf9iN+/zt9do86SJgfy4IEhg/vdXl3l+8XxuIz+wiyl/GP2
gSH0YkKfZU7epQHrxm7doSYe+fivG8A6BlNRJsuDsOeAC0lmVh/ch0ac5Lca6NrtEH7zZgncuU+z
u70gOp02tweS7LDevNyKaW9MhpzcMXZxiR3gBYdh42BzF3PaKprLsnfy2Wi23twvFvOj+846+CKr
nanvQ6Cf2Qk41AGIkKd8/0vz2J4qPlrXk18ZaWOkMUEUrGm2kENjT0BJ0MXbnyqgTWLWLh9URRtM
QRcBxwYOpAJ+aDVr15Cw+LZNIROK69noNqRnu8ZnY0KJrxiLh7Uc8mPl6IrbYIff59eAs6rEW6SP
7dFIbdt3xnCLlUTO7ojYoI1F9mR9HyGvi3SnASLqAQOi67msbX2NbPN0FfklAPbIUDeCUhA7zMdM
Gd6/tbqPGGto2MMeOwr2FXJ2FfVYdrSrYve1KsTlYD8bCzJPzvXCoU6DiJ9cwVrK94J/bhNwIxMm
TobwFbRJAREjxwGnrgjRm4nUvfkw7sBmfQVTNKX5+XLGUee34doKrL/zoZkFKFHea2ujpZ7vO2Ku
r1uVL8Svpj/9IDscOLK0qFr8SpGJCl8DxBrfcgyUpubH8LfRK1PdcDPVbL8pmOfQmGfD9A5K9Gs9
W01kQq7zpovhQ3hN4awOz/0OmPmFZ+ESWBDnw8kWxKrHQo7hYhWgvmiujpCgK3SXThD7+E+iPqpY
cjFIFxhbQ4Y1TVqiaNStPMN9JVqLhyprjgW/bQ/msiNVkNZTWMlyxn28ZsxPYRLJ+Qn26lWIDUUU
Xi1VipCy0lvKwPfMScLrmviYEyvL91ItYxrqGmqgrS5KomxQh4dASu+clAcvVml3T01AcbTflq1m
y+w8MYWtQNLiaaxUxkJ/GlOMCib+OXTwyT8uWIQTA9vYzQ5ulfoz/pHbO7ksKSyFRZ6WUlKTg1Us
1XhOl8PWo8ofTOKauEQTbgDIQ8v+S/sVMho5wSKt1jpYJQ560UZiYHi4RFHMUs/XCee3p3kJLVzq
kQMeJ5Kj+wubyVg61KH2mApWPUjqutCofQ7zaIUkIDzj2+lahsiyiB1Tna3YvKx+dbSpaZC16bMJ
c+kJhqdvwETPB8BB7EbzKuTf0mC+hpVD8XxGsIUOuycaPYQKc8HRhrpmQaBYrWwiPsZC9PduFaza
A4xf5ON1JxGCh3Fo3BgJnhyv0QoUm0kgrwvETktSeIuQ5yiF475Kj85heZT+GsLSzXl1ppZUfRC2
xp+cB4a5W52u90ImAJ/N1FzFcrWXxwgCdHCtFL4RT9F9T6gWVcIJZhdnaumA9DipViSDqHOm3Ovo
phxdKHoUi1nlmzWkMKp0xAETGAdbkOA9Z5JX4uFoGZICVIQfjQU2HRnrmWiqiYUTkcIJ169/4li9
RW5k5nkSyEL7Es/syHu40Yui/b7NdclSmM6tJxfVEKHoSFa+xEaRk3G4EFiDFqYjo5x1iSCn8xLa
jvFKhGoy85iNMsWs10KSD5L7GTeVvLLcHOttvj7ogNGFO/4D0MFS91/W9YFsqiYLejQJjx77i1dP
yPGuGS0gG3FMv0gerA6w0gy9Jt+qBZyVBVpFNhvWHF5aYkSJvetbLIrUhnUxI3iDQOiSF4RltqAT
NL5Vzvg3TEkOGnKSbV6oiZ7rbdTP+GdA9y7RIbhqjuSZgNZGgB2tNq4x3XMJiHzTUVRGftwbIAP4
XWlhK+KHFXDzmMRG7rX211jsxkPOzi0X7RxBVYKMt4BxwK8uEtay6yTUlDRZkKpBlQayCFV0VEUY
sBZlJ2kHK0lQrn8SintOcVRomKYAAR/VYgw3suZp6Xr6Uo38+lPmg+bMMKTFECSO7TonnVX5F/ff
+U9H5POzdByDb6xlYmOBMA2pOacyI9bZoKkm7SYeWBt60QNJ9jRDrn9evlNMlJFv6CvDym7e7+Bm
2fUvQrXJXdO/oWPmmFfWOBHd+y3Wemi/5SoCp3A4r2KSo9YjDG4Sp5GQNrmxmz1uyfd6td+7OXIx
xZshszbkmddofEjmAR7Bou0upvI0ePkamDhrqCrGagA7oU0izXKd3UbFwEQ8XjPTPfx3iEtYwU85
G6lB+MK40UT7by+cq4ZWNTzDsOfiEV1AgwnO56vmBhKm9Chy5T6eKLE6x/xMJi3vl+jtIQM2/Ef4
CCzo0YGtLKyDOiWXBq+Om715LKwxSs8Y0bG1CuPdZIoQMs6oZEfWqT6VAoYOlkZQzRgTt1s0uCuY
F+OHn7xoX3NyueK+jwSyA7kg65a6q/oepQkmh8mJIiQhx+YkGPfOaguvlq/uTg2mHlMyJOgHC3w1
F2NrUfPbp3eoz7Fzfy8FEZfYTM8JRPUFrn+M8HQFoI1D6D2sjbucaJQ9LJ6MjY6ag3zSFHNCPiax
8dglx3rgBHSKVqmNIGf9yr3e0piZ3l78iU446rxCsbrk973IYYXE2pVAEN4wVAV92NPHPGb4m0x1
CMTycMCQnE9X3yEx+xni8TxAD0mb9kQCF5QTugn5w+Ll+Mj6MJJ86SvaDXQ/eyxG+j/xx1HaHEf1
A+Vasj3jvr11vrbaZvctZKRWX9GhHbj+DlOrRCtmN4lszUlS8c4G9wYFteMjFOMpusf6UKZr0Xls
vMHvrc6w77qctbng8bINZ07/RKubIRK6tb9ErpinIcH8Rp7PPbWIxF2jjYpEgH3kkaTp25dl2PRq
LJA1M5MaeO1Q3kCYufCCtGIHk5ATLtPf7wihliQFvFjNlgg7PziRmCwfPINZZqLE+zAtVL+YTmXN
9ailK6wRw4xAEycaCDGH059TnNBWyxe4i9M2PIU4Wgz1rI1TSPcv9D+CzkRmjsIgG/pVXocjGXGV
yc2pCupV8nvGiuh/WQo7ZRs6Oc6VvsYMm6DvO8yrnyd3aDLNgI6ZV0HZ8z2pRRYPsxWKjHP3CU3K
fg8OtbwypyYRPUDhMzzqWiQEmQ9AParsKucOMLqTRSwfUjVfMSalLkmTUEtTw+M62TvLl+ylljLN
7MDKCZMKJKwDOWK2IOS0QkpQHv8qw71o08XHjqJt8mpULyJQ/r00zTlOdYzDN+qcMrUCoO2FK0Wb
0VfW+UhTApFmVrwH2Xi/ek7w43emwyybWU0k9LYfkq8iPFb94nrsRQ9lbeCJt+HNN8PxjDV/Jg4Y
Jvoo2tSOdFRKZnA72wfizyCRt4JIPvD/X91HjRl4HCKHlwrH4aC6ZTEnbJHYFdnWRxpAQfb0cZvU
KfXNvZS+YBCeUTjHSBMoQl4p6c8fhdJa/IXgixie/v/yMHPrWdMTlcAdPkLokUWakZbp7Rxhp9D2
0TjqpQQWxaKaxG648CqzCXXp0Z8KhZQjsBtArN1KkkM/2jFJdML2z7QbZSPRlBP9f7nEVMteQQFs
urZYEGvjh3dncEI8L3CqmsWOIEReslw1W/h359yHwinDjwk+Ec7T3g3a5UjdEJ7PC2uwvVT/RNBi
aGEEF6FvkVUETxhoK/PkNZk3uPAh49bP5nmjPIxfHaOnyvAjNehfO32TNQiIqUSTbuqbdWoVjZ2Q
Jj4M2NreW7CyQ5mxK7i28T7OBfxibriXCDueDuMzqzRvyee1+jE8seJlf6qkyolIyimN8ntvwUQ7
r/YsrVluxvJr6GQKvupFZA1AG7v2xZ58peRUtuJI88UIESaIoMY2iWBwSpX8gRIcldjVT9u1TT4e
I9O6XeOpREXo0R09Eg+A+2u4bRe3hYl0K3WKptZ8ckhLX0W/UvLU2wEKnLc2YQaCoqpdkCt9twFf
Q4U3vUIzJh8PAJutHNJ4bOdWJW/MY0Ln9N7hXsgdKwsVCHbknjENFBDYvqag5RwVVv5efxKDvcm8
XXYhvoTNLTybtHo0581n/TpN6WAVwyOZUqUozjYKo6dAHrCFpLXwEdqWrqDjUXrwF8ov5BTflqj4
q+AZu7X4k3TDgm8ylDRbTkxeXyykhUUE9rIAcyF/UkF3cqGNRzG26MkJdTLXsZhrLMDk1WdtAdld
/JFAX/aI7G60EeP+u2Dli0eNQ8QbIbfcU+ICZIBPA1JTW3CimQb7uCPN+i86M9CpvP98SpPQ4FSC
YlgSPu4CSL36xBPynv6NmQ2VnIMwCdzSd1iY6sZZUMHsk701gdDa7g+CKR3gGkk6GUfjfM5wEp/V
pn4onoOzz8Qsi/8yNu8bdqatDwklDwyZkkRMj8oZBhiUwFCeNKfbsxYesQlDgqwcg9I8NJbKbA/W
5WRs7K/d9pXTqJACZcLNKOeY9utimzGWk4ZenBA1ncUMcWNkH2rpwn/f/DFVfSIjQ/GX/1Okr1mv
QcN/Bs/5B9PvnK3lj3VeUSoYRgM41hY4BhKsyhgN6ueVFc1fcd/EMQOoTwrTHWybmS8746T0hxDY
/SpnHD0oFvXZKcv2fSPzi+GjnPgwiKvUmTjiP3c5hO6ylfk/ip8A0SJa+laVmagOhHSPlbNv4G93
ml6C8a5IQwp9Tn2Ng01WVryoKqxSlD2WhpwssBRPEqAi92ife2wsp23sOlE3e/PxRhpoJPoBqS5v
tagVV4wtndBbnkToXj9S6I84wtmKhtJlmhg/HHfDovVU+oy3zWxnGdf5xhM4r8IWrmU5xAZMxb3U
P/6XRbcYXidRHl2eaIjagBNx+9+/ijp418c7cYg8xKmUtVbTp6DG5zXyfm4v7hCfS+QsqiltAbXH
Xac6S7K+de9qXJC11jnvOB+U+m/7mUZPeRupLBVv1WlEabIMykRqdnop8HXkkUKE71sil7lXcWSH
JoznFsgGO25Hyz6RmGX18GEd/by/kn9ODu4JZ7BohXKAoP95BJJ/sa+rEixw8EmatwUgzBrr3oQz
9yfY+MJ/87AxxDRNgHrUmJpfgr6aMA0D0C4oLnEb+ZjVg3xuyEUZUXOusALlu8l1RY9KFDSnr2Gg
YnGIsqFEZblA/6Cj6V7JpR76n3Zi8cDdCZMKfiGDKIAUcIiB7sfo03ohYh+KB9uwdPyHMUNp7pbX
o/1TzI9F9fv7bqhw/5vzM8DuwRgTDdUd4kk4LprVKDA7vaFMG2gSVU7gwwE0RoDJltK+V4Mq79da
evRKpLu/gzJP59hHtuJXzlG5ZzSPMOW9MIXLDTJH7EV2XKAJl5z9qCiM69+Pki0LmW5nnz+iKnPa
bKAfido+N5MQ+yNn/U0eW8oP9t2dqs4F+GG5g/KqG7lc83YkffOsXKAMLOs+H4jmrPXvVxjM4/Ad
wIBywGGTD52Qs86q5Cozai3VeHj4a71SU1oaoLUeWGUaDnRHuZA0RYZocrQHolqykxB2XjeHAtLk
Wx2c2PYCPc1jk5WV6douhKPHFuRJToH/Lhp8Hlw7b8U6Lhi7agki2pBwxwBIDekzYw8ZjmP5Qadi
dOD+9EKXSvygXCVtoVVAVd1LneT+DJR47CbMKFkd+IIw9ihcKXXACaAJl5l1LEHg2h5u3WVYCndQ
zcaL1E5D0cZCU1Dxn85nQB6EPrGBaJ77nKl7Eh8uZb78YfYzqu33z70jz4bOjHOOllUx9YHGzLma
53y1pg3ClghBcXHuEq7wzSV2myo33bd/SEskGaanduK14YwPCe7bjCxqy3B/gtNKSRNjRHPCb4V3
yquz/dgTDMgZ532x+gc1B47O+aMCMkAP76ZcsLEUSBZe+js3mqE1VJpZ4tFtkC2FE8vSaJ+DG2P3
i+EdW3NaoMYLeNDDQ7AkCT4ml/BY3BoAaex11PKDXISX/O2r41JW9pwWzNJonEL4Bvs7jjZ68Yut
jGuzBrOcA6Hwc3zQZ3v9oO2j7SOt8UsuCEOKe1qPKfqK2XFFeScS2ArByaQ3KcTymwhMHrKEripX
+aHRQOabO2wzX/hUt7fg0Er5cPU7OU/ocaf17SUUYEDC1SSWrrkn81/FoXsQF14Hnwm+gbqxbwha
TkRM5AROXyocYNCUEQ2JMlU3sXwCYPg/mvYxTBJKzekhcypeYlKh3cJg7gVpFOo7whcUSpjloz5m
OXnSukR5cYPt+elIXRzo7DaxIEoJE5/ByKWcZmKi/gaa+5+yKxcbJpyaDwUAv1Wd7Gs+STfGMapV
Wd/u9+7UvlmM9JOv/2dxw8THXoWpb/dFmyW+KxtxxoGkoHWsCpPZIXxpO40uF6lemlCPgdEEH4c1
9wQoYdbIdULI95+lD6pguixvaRlrKqh6SYxDDiLMShpIMII15GKyEhL5hqAZbRkjawF2o5u4Zxds
hZxKzujTh/GBpJOpNZpXs+eEGSUHzU9Orb6I6/ePZZOhPiZ+aQ0cO4AUjjsIi8Psf2S0g02I90pQ
tpHEgqxtzpp0uEfoUQa3Qg5benHwjGwswr2SNP92OX6wB8d2FA74YlYswwWTYEFz5knhWRsPhwfE
s57KbWsYbfkic2JDE+4jwRTyoAQ+abA19ArKzz6N6ICJMRm0FV8FbZt7YKONI43LLljvDguBPCRq
iRhsJ89qoATocLRbcyypwWEcxCA4/ovjl9PEY01R0VUeGHcoQSIqKy0LgaNkCxVxdBw5dWSIevZ+
Gwv2XlLNU6HI2iH4NY8eueGFAe6BgSwQ99aB/6xjXVm8v96kTmZkVrHPe/0RGBE7QCEeh2yeZgzN
J+dMfw4MVPP5Zfgz1ix/kfpL7pEN0mCfrsabK3v9lV75BJtH4LOCnAvSdlPsm9Lgs9VvRiu7Mdk0
Kg1KYpWAqEeRKXfCraaVNAkuI7w9ch9/t+nHlfvw3gM0e00S3QQdV8WwDwvEDNe93Rf/bbzPfXrT
/YQ8jipz1b65lqaKNgUpDAi5CG85lg0FBJxR1Kx+ELH+KFIwpq8CxHTTqh+jLyI0OVKESIqt039n
MiXIapOmdZfvUIFZXMlAra/qALPWIC/6p3IyK/zRUzTbUt9sQ9YLNCpHE1bAvBUb0xoSMChALJf6
0tD18ltK8xTBKuT89Vfg8O7+qI3wTgyrKS1SyIo06oDP/+FhAoSl1AGjHoiKGZlqmHWyqztiHCZA
mrtAfUxMJBJZI6YXmdbUYtKpw69cnpFXZtYMJRNxQKJV/a/+wrhecbJQxBIrHgYxgui9eQapLaLE
g56N2M4gcEt/WM04nNTpWLTURQZOExDrx3gjZyXHD/+slOM6fAxHJa+vBX9w7SWB2DR2ReD2Q2kM
FC6Vc2Ls44m2mzb9hurFN7WVaLfstpzCd5RQ9JRmo/tZhp5Z/6F3pFFqs2YDXbDUfZGRGQ2mIJUo
wsnSCVDZo93Zkd+iMamSxmVYVEGmDMPrWlONQK01abQg1TcqIGz1tXIhSGuo8VHv2B3am1Qzmkvk
VyvwPX2d0a6KSYhe+H/qSgT0ynxxhdeJTHnDWdN7MSQb6HPQwUnCFl0LFfIbpiYop4dWoYPLRAj0
ZXSuy04uP46Ut59yS6yWHdDyem/ZMjQs4bVh7xqLNO+L9tOq22799URVyAF/DXtJX4bvrD2Sbd+D
79q7r28o87xSz02IpI24f7sUS4vciyiieuXrFvswsBifCcLGpphqiwG90Kgm6E+Ex2nUoQyPis1p
T+usFWKD2no5csLyJEBv6fCVRPgUA87A5RJ8ZKWzWdurXvibQEUM8RpNtSuu8G43+4ginuGBVavm
d/EDu8rDJZ/R7oWx6S1T4rXLeI8ZfXn/oCnyrtF6SHK1+G4aUp6Co2cg5mmdnuSnw1NahKGQEYKN
VF+sM5ExaTeF2Hen15bcfXUV1tzVcMfRY6XaMoSBPaufxQZMah91RWFMhAdMaSRSHoppqcUYzjNB
tN4HcaDs4KqbQqLJtGWWYhgrVT2GqW/Tt756FShnI9zjNf1oQ0XafTqqvf8vci3moUIXpASLIHGz
f8XVTQHNzxQoK8yIq0pPiCQerum93ZxlRz+wnQN3rKwj4N9UADLZpQjkv9gs6p+FmsbEVAu+9UZW
2lkrFoh5TmBtguMIz7rUOWqDcPSJNK0hfnF7s6F4ipT5mPDRH0/SZ/fZzyc+txb22Us4oe0/I0S0
v+J2+sQLAOk0X65DGjxJHh1SSuY9j8HPzgwEyy7acm5WXNOu/WoSaRnG9Pa6/OtrxV7THWm9guen
xtsrnugkzb6Q8vkQwo7u8QJjqrHMymc8SdhraG6XU07J7hJ/bnUpkjWy65AgDxALhXXay51L7Pna
A2bWjuWmEabzIWiuXNjALoM1cXmoLyHuk8waBwp4g8lkiOhS6vW7oOFn5eHw4MAmj89zaOmS1mSk
0+Vzrrj/ODVbnCXqqxOssu0LVvYckdkBeRuLyqZqHo3rKeGvjcRzheS4538ra+iO4R+mMqnR17GN
hSke/sANnno/C2HjMs9c0tJ/odTHsweCFhyK+0Hnyhafgunr1QK0hy1tbkQLp7k3bfXo7qf8dxbQ
SrN1TWbT6Gwj0A6WvMaA5KQz1DTnXA+/+b7kjUKdj7ZiVbIvugLjolPu6qbzXzPaH/xzsN0VRw0y
gwlZZTxnfvHlZxZqZhaqB0+eiq3hG+TcPzfuoW7VkGDSHOuVf7S8hh1moHn4OjNHr1DFKOURf62i
lk68g8ym1bGQWf9/9jtDhPi9nkVEaHg/ZJsb531fFKksB0kzu2ftAa4CzVTIyBmTGnymsVtPLQ8r
4Wqpj3DLtt8v8l+umtJJ7PVtkAikn3yDv9ZHmSdEj3RJWPFZvsHF5GnVgET4u3WpuLd//QBtywJ8
xEBTHPcYDt5RBlF1dQw2yIKbtcaA/N5TQ7616g0OW0gGejg0wUujLwje4XWFiQeZ102e4uPtiQYS
p64BuV2+Xx9in7WG+rXjBOm4vMQPA2kh47iBeQxuM1jTj/TW4iXacRvfpUKPqhlDVGC6EXWRz+C5
RQBzrlWvSs59A1kxFmtwZ0FB7dntSQI8dz3QamzLTZ0KHZB87Vn02UHEiQCF5fulyAYYP+OQmBMi
4+rlG7o+RUuBKF7bz6QGUg/I/nLg7MdC8d449BGdvZDvRTeWMgJrWCcZjmPrDfUNn9HOxH3Ju8/f
yPxbchY18z8RLWF9jdqQ6EPii52sKvYcGaU9J6yKlhXsTs2dtsbJK3sqMD9MzdE1u9APIGDiupWM
ACiHfkyAKh/YhxQ5Hp/sbjnZLwdQQnRHjHAXRQ6MTQOVDAYnnrdYlTJ12263uC6/0j73yX6KxMXS
J6agtmAxG7kEsc+TWVdrKv03YHKkNI86KCL55J4eK2ebc+/zMy1492WQRoF4WwLsqFByN9snMir4
QoC7jAW/VIzH14YxUdh5a0hwc+ZrFWAat00dFq0V2RKkm0j/zsnXbhHNiqrwWDiMw6m3N4STy9fW
7hoPgyV6zA/jo6s6EhZdAcZfhysDc6xlfwarxZe74DQWLRtj8hHga+lndCf+sBw/JGNRYLc9QtC0
X3gkPv5Y3yOtLWhzb2PtatwFD/hRCDTGzdDiVW/V4UKmHRdg952HanUqP0UPP2ETtLj+vH0x1S2Y
H3iXckUKLEiXU5kPARUU79aebWSsf7y1d6SX6W2w5WVHPoUXMMfyjqspMawR/iH0onx1OE2zn0qb
6ewAY8qo+kfrZjXoiFq3qL5PMajl8CZri/Ok3z/etNaO0d0hCE5YtAXF3NUTAbXB0OWbFdmdHLuF
5QreMzuyyCTZeIwzsR8IaD70ZCLzq7FGAZWLhh/aIJPuNuwiMdQiT6W4tW3Hhx34AkfqYQqGavxg
xHOFClptByksadg795eAxwKfTjMPkjiD4a4g6EXbxZyqBC3VctzNQH4V0SfqeH/uhSTBXIpM1a7F
nBinz79Xp6ueYIYx7bYo1dLknpHcJ5+wzTiVpdoG4X/dZ+qV8b3IQGwnEfoboAD7LvX5z6++CGvF
2LyuapFV64AGugPr05SfL150ubOOfVZh4D5zCjU6QRs/UTztPjsggqJJF1KEPMKqEOLsTFhb+n+/
rbcjUPgVZARjcVsWywcoeYEWmfLmesddSBeXNBa5igFdhGim4RxYSVfcDKYcVP7I6s7WWADEEkS2
O6doithzOGG7Lb9ODHSmyGGR6RJnETi++GazQyXVliJQwuuiH7UAEVBiq+CHPSB2OHCcB3rBPhmR
suUQuFThqGCncR5KEYJpB5SW4c7su61JfoPzDWWclmbvrS3U9ep5Xyv2xXaHQkcvFIiKayfmv8eV
dYWt6otlkNlvVNenFeoIRMTcP/7l8ANsFF5ys9WHZuFb/Vw0RO5I+ah0sIoSpT39lCKiNbHCw+AQ
PheeJYakU3rl+8JuD2IwDlQvjb4eQlhASVkEVFNLw97ncvacD644P96RlmS0CQDkeDvshuaBCfZU
dXIJv/U9uf/ZmwgWqBfRQM1WVIZnqDTSSWAQnm3B+DT4AUWQuYEIbKpdhCzL+XuDdWbFNWpjDcPo
2PP0AL1P2FE2iY87UVjqP45acLX3Nnn0sV2kzRB3cLWTmwrwue08MHtb5qjJn8Usy+/BHfnhXmC0
iynj+DOr8R5lUCQIJTSfKunJoOHbFS5b28U2JQpC365oEkJ6HKeOwiJYrGMNhWjXFGJ6AStZu+Ut
n5NNc5jMeJwRwpFkYyMEzyBSgLk4PQWQUUq7hH7oz3g0RfyoARJ3UxaOqBybqHsLKSvTBI7wS6ak
myjNFqc85qW1PqsT4+6bFJYevGiEbADnAhkHsqu32d8+Go8AQLJTTFyZhjnU0LKBAltfQV4JKpzq
aE//1o+O+R1mSHHGHs+c1fWQwpZhvw35oG2i3GixbBfHGd7CmoT+SHONgAbQgWX0Xt+r6gScQOwW
qNsX8A4Svod3FCbnLU7IjfdQL2pUaomd4xBlE4VcKjzh+4O2rGnKBjlrRyHDrJ7kr9dUHoMhG52F
6+aqTfiwCFBMRgEEMl/in5ETXJPxp1ap+IC7cSF4JO+HkW8r7/NI0JW+10OqGtM1Pw10+EfUzJVY
ezb7zI36oHRxg6rm7zUPMtmP+4C5Wl6tF7m2BR9FPqTV5ZaIYSHB4kyL7KYTUi+JxRQu+1sxqRoo
zk+39VVyYgM6uWYKJKZZbYTFiqrY/hSS/3IY4MMu9EAm+pdVLhPa4A5dE6l6NxuqfdkCmLjiegRz
Z0nYjsAYfnAjAMFT/G/zlXaL8G07727055wEVtU3hUuy+bIRUeDcg+f2oCHRpkjwkb0snk8FtwLG
ATf8abSVPn/dODBIlX83MijrPrYorNlXWzcGlNWovd3Vrt1qEA7OJ+vBRkj0oVSIb0ZU+EAUvG2I
7X+QWUX7x4mLy0W7RvLb9T9z5CWns+Ya8xmM/QRTFnDCmck3Rkpnu+Qz1zrnr1RgxR+kSS0c0/7z
UcIOKuGV7+zgf0CCXwsVk/CldVOiaXN/KuTU8Saq2rQWKzY/KkZXxH39JmNiFZFpcraP19SdPvik
d2l12aZT1hZ5B5F8bsJ1YhLphoskpcEA8KFhzTVT/x+ZDIPV0ku+/EZo1uSqjFgOUGN1IHUHeUAl
o7Ibxr8enbdZLqmnOKMcSIuFQYZzlSgvWw8j8mACElHWgaEfVZtSqV0ky68xkYSBrC+hm4nsNpSQ
TbFGPPX05tC5k9m5TyfRfuarH1dDhgmkHJJQe45X5M9si4MLt7s26zHyz4gnYddGVW9nzfDavMPm
iE2BvSutNyNJizQ2PAEbSrfyerEwvkmbUBYlDZiN6I302r8TSLgLf5Q8tDqT00OamrD0VQXM/XMe
pA0eNBiBhTar9vGDtQU8sYV6JWmbR700Rebkw4Jl3bXb+SMLjIlvSBuEGfMjNyPjJlQkW42ykABe
1ejYtl9t5ohTmT4oZrZc0Ri5kZtNlveVoEQkBAj6Ka/WzxfR9OsZips2lduUT41idvxaHBpALoxH
La1SR8GcqymTYad5W2IIe9HoCWtRkHvEDYZPZJiGsl4OT0JOx90c5HJUkDqZ/lj+1ps3Vg3cBKbt
LneIdlBgPpCyy+pOiSqg+uZQyvlXAGVGJm4ahOPwfLkVJKJFx9z7Ub/7BQo3hRZ69HdW/5sglOEH
n3LxGB6GQ0mHRAHd3QPdiul2O/7L6rDALhMSzYwPFLdUNW1mqzlVROkX3psS6w4UTZjuE/Nm+tth
a91wxD7PpZnLRWpQ+NLvmDdhrkuNnHe2kmHhngIDn2/uRbcKESpfrNbfa5Edv2x2lLQqC6MDYNB+
dkR6C74uvmQTS3F3qzQ6jHHKXufhC77AdxLsFWAEDsW9W9egxpGS4Mq9+Upf0O7Rm6oSl+MEoxKs
inIiSBZW3RwtL9BOeutx0hRcLOzVQMF6KeieYpzg2mZlRSBINVB556TmpjmaBM6VdZmlNFOd7s4H
bUf2S00/Wroc+361KTvPxlGAgsqJRzMeGZbWajn+MHB5nf3fOLmBLNuipsZwiBCGVycJZUjJs+Ds
weh+alJKglKZvtnTpI0uRG6KvNlp7DvTdtEa/MfEw5vOr0WmbVXSUaCL3NdaznLxdFlricN2bNrA
kqJ2XJ3IJfTOaYeZwtElqbGcTN39SLJXSZgoDosZLIlFy4lh5Y99IUIcKPVMOUNOrKkaz8rd/3Q6
ECkWKaat9AfWvfMAuEyO3scLCpcZ4KJHtbvjmFZSEv74vCW2FkJHqjSyPvtJ4c7VWo1Ut/UjWStS
XE6luFg4vxBoZajhCpwbZ0bqkbo1qaD8WLDTx2wBgH/W25rqRBzNaqfgMHOU5mxsMUNqtyfzuUYw
W9NWGYx4984E7KZbfVUldiZP6mOOMhi8+dWXGVSOG6j9Cbn4ImgAW5b+g0EmUTiOcH4sCcNEq1TQ
iiF6iExclz+WhvMjyK6+7NnDorJAAL85uarI32DCNKm/v39SwQNfRV9SuAR/C9d8DbG2JV6zaXFL
63QMe3dTxiFGRQ1gK1c29562i2NdCr7OcBMyGlYiuqUhNbYCfxR8rt6bcz8Tbc3CfjWLffP28sj6
Q3N0MghyM7INiIVi4R3LmcqZbbBYN6T4tGAYdsT0rrHyDm583fgoDngelR8eKn/d0YLtQG6MWCP6
WZwm6HXNwQhBS9caI7GCXD7RrM2dPNkZNQfw7KT5ef72oEQfT1/CoPPq98M8T48ZA+U9o/iRSFYU
/J2kT7OaGc+XhHACrD2Jx6Xyb/zQnA7dbEtBSufmEDLHaQEedKy22t32we4zH1Ony3L/hhonk06r
lYvoSGDPesuuObBKPDuogLgoR/t7lp85xbp1DlsRG8IdP9miC1tpya5/okt1W9zOm8gXyxqREGpi
ct8YdHwB35Vq51Svw9ot5DWxEAtFj7k2+2IAfsPefjLVeR5R8L+Efoxs741jSzWxNgWC4wqJ+qdx
MzF4MhR2B652J5Jlxyhv4QluO1qaJ+SOXD0Rkd4r00CHtxAZ9G9UDvGilXPyKWxR6dYMWKaqgEFq
cLS5MQkkWjclxaB6Jjf0j9ssA60vnfOnDaYPfRzV2JnZXcbF0q5ucPv/nYAyFneKpUEyFDZ7QLYf
q4bhANddwwfG8+sDceTZiMZ0Sv5D6OrLMfWZSkDEeBSVKP52r9oPY8URik62vxJPcmKqaLmTqNqh
EQ1MTgIIm4JNxv4BoFvx2hvK8GXCVafIj2lSKLzt6LJmQZ8Nlo+LqbwAirpw+nMMvX2hz/SIhZm0
STIJqLc3Bdt0gv51Ew3RS1cc6aWALBtV4b3/4aK64EFOHb1ny3/WMj5qlWr1DaCzyBtTm+E4h3Ok
qIow7aTsnsjFnBZO1huWuWqJJsKmDAVyRaTUiVQDXRf48TNAZ1LZFbwyY++8vggoN862FbormhSQ
ARuIZMWoJz7/KRLfQMkEXGZdvmqK8KgnyWXslmzfe7WiQ7bbaB4wxF9EUUv4hA0Gzw4nMiPuFq9a
2hNAjDyY5R4aj+57AgLcMdhFR8ZNLyTDDgxeaWZOrIYdWZW6iPSO9S1EL3bEbU+wC4jeXIGBd9kS
zKlwciObeLdbV4v9m1J5wi9W9u0y/93jsh4N0GdirGFF11J+yiocOmbccgxsy9APUxS3wLA86kAA
R+HBpmyX5UpgMXuwR8t//ZLbRU/J9z5dWau8I3G4leBI3DzTIVyweXIFYwH5c5RiP2ZZE5rPdc7d
NxG+YI88IQB9fZWDrzt2KP+FCsaeTv0/YCwB0UIyLzyVItphAUKvJ23ycvPqt6RfUGAomd4PGbcy
1gjlj48cwRSn+y25p/+3IZmpoDpV6T0Ai/2uP5xOoX07/y2qRt2THeWarRdUJUCfJnlsGhZN9VOO
9a+KsrIXe0JnkjQVjqq03yHjjYHGXKYF2HpFceA9y0rDWoKbm6hiK2EroFNqDbPG0kBxuZnjygU+
9ccPBCfNPWBixJ3qUoUY9FngR4o3j/PGqjkSjuCwhzJe3elAN2buPae2PaAWOpsloxrJGus2QePy
78UNvbuDyNEJA1zSNCuXz8O+wBHJbK2rU4WB2tisLDZP1A4rzE8wekL8V/lxpJj9+jQlEHfVmp85
1iPLwEBJ6Y9CEHJbhVERYQV4RmnECJ8o7eN7mELCKTFFGzSRSRFDf6pbhR2pnsTd3/kIuArOOHej
Xb/wbX7EUa5KphrIU/MSRQjXsld1JxfUHLWQnEyrJSfOKTh+ceCZnzE6mf5wQKe96IQeOED6PTON
RH98ggdbYGTikxUEGWgcrAeG6MQM5TObfHVxyIIV28IIHtU0x8nkz7/T1q2lWI3KAAw7IlGmeEee
oK0XMfeXGqNy7dwaOpvqOzu5tbAupn6s7uC6WEqNbenpGHO1xRgFLKN/T8px9gpfagWjpJkOU3PH
iGenxxb+/rj/u4xtpvO1W3OPlBBaxilo5zYuyJa4NX4dPzh+i8Hlh5d7qlvXMDE3WH7xx8/fJ/ni
YagDjT/cfqSxgfE7LGG2/BqEqxQKoAxBxG79OwXOU1e4AcWqZqm/M5gifOFNSS28E/xUNgHqlHuN
E8aDJ3fNhJPlaGA9/1GJNA64YPJTj/3POZthDBiHEQIXraGlHVDPGHmG7OPxmasvZaNVlo5v/I/Q
ZguCkRiBlbkXE3CbE18h2aR6mYcSpRI/EvXU5WVvHSADebzj6EvWDHFq/oQTSRmEBDAvtgUjL/sy
CfqB3K1SlYhU/51Pb72QTy+PlIscQxddzgS3EItc4lc8N7TI3dS4rXncRjedXwMG8dX1MWiM85bP
rQHm2I/mTujPvSlESLMrYK2w07FZCn2RKEKF0ggA0RPMV0Z9rHAEmHy5o5sQwP/TRyhxpLult9Dq
Dd0G+Ik2kvx7Gy0grEW2Z7zUHDHgTaLiGeSn8327ZfQBlmGsvNWlgQV42npXUAecYDYNbRy5qOzj
nZbajTQ5w64gaWZdlgB/X7Pm4k8ABIIqK5UC/uEIlk3Rhjv3nEA9Wqq137GGM0ainu2iZ3bF9k1G
4bLsln9klv6CsZVHwEOLM23eZ/s0UqcuKWlpjn4FNkR9ovKCS369X9NZE+xQpqhcbM/YWv5o68Da
KcrE+EMlsg8KS2p4Q6TL/iB1A/v/A0OBH5gVWN3c3lL1oE5NPUjnCE88QcYou1t+wrkT+mAdamAV
VoCWxHFuCYfki7kIQPJxwKcJOEXNAOHbte08teVJBOR72u4hZqbwW97CS3P0lO/6dmZW1YHAzumI
sxTTsCrVpLPlErQPmO6KLbZmSx9VApU/B2xEyj9jgd2McJnsZNxnwkVoYHMUP5Hwjga1cNi67Ku2
ce83WV0mrpzfL+BfaiWlU04g6xgZk3MoN/0+GiICl5VHZ2OTbH5B0tJ/1xtW9u1gjTA0B2r9T+Fd
qiOCpqYP61Cqm5qFX9mph8nLjia5/WuBt4bEdppe9Kaxm/KHynz4ykJSCDZ1Kc0Fc6KkJHOlVUy9
jn5kjqRlJw3xWmPVqj44I3Wgm3il3feRdW9dh4HvVzcXCQQf0p3YZP2hYruvyLxWWGV26yWP2DXo
juqljkqCnUpgQZ4LB2BdBVeV42y7/DrkBIMjGWSfAWM/I+orFaGc9lTwFDpIs600nsdkMi4Kecho
mxccQGIPMEszLrmh2xYvcwgBOvOMJlyapcyI/b9i8N6tgWin5GIo5vmeyhjTISLWFXnBUJoKZgsC
YEpYm0aCV71x4+29rMU54IpHkDMutu+nSY9z2k6wFvTRbqoNdZ6LNdYLqTuwIlCDAXL9OT25Zzsp
Yp8alAm8NHghcVdHsYLonto3qDaKN5zwyfmKWkFJzKN7tb1pd9r120oHxYB2bym42HLvT8WIqm9u
EJnH5d2t5UGTlx4mNPwZqwGP/BJXY/hDmcOiUatsrXWc35JAYbsw3Keoy3COpDLdE+usceX176RU
xUE1kBYT3h3iwa7qBH856FgYpVcq6GuqrM+ZvQR1CnvKdBoIKlM1rYCcQX2pCpRVOE7oguFeJAGC
Xf3FT+/s8Xzc3gtC2/yqLiUbh/MqcB+itTjij0JAZptTZannmz0Wjc2bLtV7vyhwOFGB9OEhPAgb
yocgeDNlA6N1/V8NXcYPfxu+E72vZHVZ9HeVPQ7dQ0peOMGrdv22y4qcSntUSs/S6qgzjhL/TOmB
E6jdJI+s5+EFeKevmZPyfciEAoN8P6TlN425J+5CBB4Z6TrXD6NrowW7/RZasJg3vDHd8z/iEdCq
HCiebBbyiipeOYpci31e/0QlPHtUrISSvpUN+OHmFfllq+pQdmgR8DZ6IFleJYGUeyztw6oN369s
rcp9jRcTz1CHeRAdwqd2IDOqFIh5qX6cVSW1HiTYfOfYyPdIkvWaeNv93T2TOuC560qRjyscDPmz
0cz5ADzBowd4uEZl0s7OxAHdpkQoG8kOy01MsOcX0CDrBBtfpiOcBot9+EsrDL7zEiTUt2XHNupE
ensFUfPOCxjt7w91n6AoK3AYSlUnr/MPs00f3Fu7NQmljuaYn7NIIHtgkrcKd5z2DjjYYLvZ1HPH
VJFR2lJ95ZNIxj3Ihi5Kk4m0CENu0C1jyCkrSbBnni8PgC5CT7dTtvkl1P7ss4h9Lar1VMf1oLrb
/gfMHvxOHM+/YEtqArX1wTgnwyknbAiCHU1LCbkQscw21iOtTWh2BR09iXd/PdNUM4ghcVnZnga+
pQWq0Axf1+Ho03uPVPXzc3Cw4G8uZsdQXLTT7sQbvFMDP2vbnQEMp5o32ZSCEJ/M+osZ/3Dlcdph
fpUacgnNGGDs87vPqFC0RMxqqW0vxhy+Ehw7S/v0vWElDcjHD4XMJuct+scoYBop1CpV/iwcPdgc
7iAzl8rXarbvVQPLxbc/xemzCiNZjAA+3Gug203W43SBu/wyntFItnGkGZMtWKxY2pJwxTWgaGLe
0U9cRfjQHMg8qRRXFaDGIdoz1066DxmLFUcy5K8e+ykVU1Cxg33HZv98IuaV8CehiSy76hDYzjif
u5hAn1eajU7nJCMYZi5qwfclnGHY6NStDcaE+C+6vwhfeRZITvNTDGD8IsmsjfpF1JbX9oARuZ9+
Zxkr0K40lkOtaU62M5UReM7wxOxAgcnmD/schVL0ESPN+zRK3Ogn/0jCxCv3vDmySah9Cl63InSO
QLlmbYO6EnoOgu8jdffr0JzekHQxiO1MxzuhLav7lNpuBhUn0qNnYFLrR3SSSyfNtt3TunSAUbws
mltn7ZbUlumwOq/D99LQhbvjSwQ4nxug+MbO2pX7z2lefaQPx7xlu7IRzY99UcquJB5uKxMlR/q7
F/W+8ZZZ3VpGFOXvymCx7h4AGtk1Eymnij2/3SmajT9tNjfFvZyIOrqzh+KWmebcZoi9qtSRMh3d
QHVSQ5YTMA5HH8AWetN7Q/RjQwIYHFvqv0T4pcVAftF4ct0TufosomJ268v9cnJ/zdhaA6L+gHmB
KQooWNu4pie+88HIx6btXLjNqb8bu3AOiSS1IYXk4BDiQA8/TYUVHJS/tCXiSVAiSQE3c8unj0Zh
bOOAkeiUxXECPKFLW6+b/bWxIre8SZ7nCIbq/GaZnsbfXXHCW45yPYN7tEIol0+8/7BfFODboV5A
yg+aYOKOzE/WAjBcwc9QdmBep3w8UYyVrCSgSIQUt288XF/OEP9VGhF3SgPHwg0ioKNd5spmLoD9
dUuEbEVjjLfM4BolEad5zSlhpMmStAvNbfFxVrc3Qiqi5nEP4LDyjIv7mooEpeQ8gfaKcvsHsbEv
H8CFk/N1bL6jjaMWLtrwB/+6f3Do/5AHK9guLu+5zdoayGalPTGJ7G/nSMR+JTun5uJDwYDKnNl9
YM0dW9fGuMFlMtcUWDOKfjYp1FlAtYJC4FP4WdKB43xn6RVbhtStF6spqbs6EN5LQpGPu7xCVQWN
fo6OjABonbb6DDCvCjdKrDK86egXKOSgb+sbFWdH2Yqp+p5M8WYdEePwo1VVK+JMLmCrJEy7IZgI
I1wU8vev2XqayeG3U3gRPY7vwOLIrjbQyZRtd7M6H0MiSgs7BM8vaKFZWqmxgPnYbMPzOXRG6s5n
L5jRtEea58gNX/lItv8+MvrbIWfmh6gSh2scOgQft6R7sQkxL1uWCQSm0D3y1jpjhrDOZqUF9aK1
x/Nb3YsRXeXAjcWHtMYPhhexXTMvFBxZinRKZuQmZOp02/KxLO7cWaN/WLdiwca55KNN3ATER5S8
y+9w/PRW32cAUAlkZoVDr5cmAe0ObavVw9u3jBxis9txCDEBMAnJe1gQ6EOjo4k+ErauaaKeT3pr
gjKNDqeZz9ZZ5vSiNcj7h8XHVPQI8/IBH1Or6N3SDDiYqYkd0ErpVYuhR9g594Ynvp5mj/wQeWzF
4JKgZqU7CagfUU3ixENxwYNbgVywqFt2+vi7qKkxgSSLSjx3N8Iv65ExX4lNYB2Lm+x6Q7A5Cxxg
qXedh1xoN9rmWgZXVzf6MaK4oowO1GuSFhBcZNosTloZjgzWS2kEqEpL5O/XsT9N+fZGWSX8ugdJ
zyUDyZqoitukmMzNunCddWmKzbB7g81IKketzV1iMk56eEESDr0bVNjM69vBj3KdssszQvAOfK8d
8YFDPjaxqk25BIHvGyDJVpg4qGCv6crvWH0sWLkplZg7LytITsURoE74sl298MSCKOHeyL9dqg5z
g11b0omvGWoGanRwOkoPy1/2MTFewUQAR3ItM3hhLM64hqPWjHz6iptlZy95mlaHvAMHPqb8ML2c
QrYkxw8lQFrmCLnp1rV2V+al4viBqu79uhSgFETQE2m6q6b7qyL3OTH2jgPvqpkKuLa2C8V+jdfk
1y+sbNHb6mWIUAdm79lpw6FwC7LZuhShRNoP+HwOBZaZi34Ji/Fk22hmGqSMSQBvzekgv3oRp9xv
9gqkv+S8lU78kyVfi3y6dKlTJElbjvEjLz6ndFprl8+g+NhCgBViPsy5bXHITAfXvphiAkV9dYbD
tTcfOZ1T6A+JgwXG7nKfu7cZONVr2i4d6G68mEsoVkFvUI9tjcf5IkOyejEMRe6WwRqXXaXxZ41K
cSxso/8dPWjBD7U41n4DaxMFxDoU2ZkxO207sCrP01blD1KVuoOKAckGh6adj2ND7w3zk54e7tSo
jU53JKxkMs/H/UrpCjVcdbULSoEalTjqU2NU9cdA7UdpAakPUTx1vWFXzl/0T9yelGI5Idvsemta
MfBsOoTQgn6G/2nSYe2wlW/uldYFgUuhfFLnKzKQiMKmMT2+tDPqmZ9Zl+6mvtssve32B6o610qv
9Q3FzVQVkquADrdAAPkUxOmFq6nqIrw8f+GFAdn9456WMy9RY2nqAYXmfuSBIQRScUw+DXWtfJCz
pLNN0gG7ecW0nw4tjShlYTcsuG8+S6OoMQX/1DE5hdr+qLk8WLACDdWMdLdiCV7qLZ1I8SaK8Wtx
BfBsCpUYJR4DjWYax9OpDR9Fiv0j94TF7CnDYQcEmEXKx5pog1OHyFBm85MhKo61Dy16AYg2kusX
75wIT2ptsIB/Dd16i0hCIotMZHNWTLL6lt7a/JdKrAfK+kejlVVmbhIgQShHAJ0aENr36L0/UYdY
oJ0zQtRtYM1St8iRfhGzgWYXfoJL6xVUuc/5UuM5U8fNo2EmTThkhYY42U9iT0mAcKvC3RwfSwjO
2xKwSEt7nQ9QSmVRfGzqbwvgHcqGYRnNWvwnIwf9Fp40Cs8lTsFoYAN612gyMTVe/1S23EJLFz5u
L5yAg0lkLblXOYXM071hrgn9jd8qy64Qhnz4LtOJP7kJkGBj/Fpe/MvuLCafZnLuSV1LOykai/4+
aanFCFvk70GUQyECsOURwVYvmzbBF8ahztLwh/z4lWfKB/xpucEvmnpTcs7W2DrNhOMHg0ckas+J
a1dptG+KGZq85IghyucZXeqqKrAeRs4U5AXhexBB5jEb1RGi2muRT4XPEVAFSAepmjhs6SucOtci
x9TtfxXcqaC+3rd+UgC2eOUwqGQ91RPt/XgsFtxXVatag92dnFilyQQcIpqg8FYhFgWaRS2wObXB
p2mBbAo4aS9fQ7opvdUowRNkgRc8Yk1m333WRzXKKohBcKHpp1Pw3Ii92Ds2/zDCWDPOOjUPYt+m
H5iz+0eLWyWPrdhhyZTH70MLLzWxZahK6QGCERXRcA8kGC35109TvAn7RRnFiQKy1Kb1p/QpCvEd
biT+DQPHFSjbagAyYlLG5bA4aT1MllbEWkb1gcpDlWggVp3Og5rKouQdLjhXMx4tQkVX3WBx7PT/
kLUKIjvnAk2a3aHTeAMC0cPRPj6gD9G9D0NtBGXPzcI8wtDRxHByX/mPf+Ur99qBMqnLJeSanEc5
LvD9YEfPfpzHYOxGEnpz1tMKwBbQs655vHBP52b+QzouLgl9Qs3hVURx0T8nFSpl1trR7kK8uCI6
3NrIohNBbNa/QRUog1F8dwxugLiU6e4mqnJeckw2TcIv1iCJ40IWlLAdITfviAcgXfi8JU/uHof+
XNmMK9JV4vs0d+LDhGiMtTHpVTr4TRQm8FXrzYT0OsxDu5bDPpvrc6o7lBR0WHGoLrVYkDSmlL4k
11RXPMHYHFfG4R3HxNBYyWW4DP7mhuzGQHnPTv8Jm9X7SGYYbO0/yDRt6ej+QgJBOdymdNVaocbD
XpjmHbOhiUdHp3cAlgxRp1ARklP0DKmlaVUpbbTxntVWgZVnlAGHzyV8smN4GBfMh2bKleIlIRki
5WxZMRdcJ2WPHXrR2uHN9UMN83abQWGxOreYq7sH5hhmfmlUsobncr59KoSmjW8L3aLPeqW+Q86T
Xb9L+GO0WEBbkY6PqSn3RMV+v2D4pisA+nijScM7jWPReiZT8Wn+TYspfHIUS6BPoQsNDEUTIqV9
FAWlWF3PCz8f5Jg41fyFtRw9Qs20KaAfQXag9EaU26fGYefTHWR2582e9YQdbL1lf5I/tcuB/A+G
R85nKyPZMswON+QZPS8O0HjVzJge1zbLXApaV7uPapa38LhWR3lU4RDgxlfdHedR+cFg7S4D7qLV
6Qhh0hKf2qyufqjEXhjPZCQFpYdBmXxOVX1obLdTvD1W4Johc/JDn2nXMv+CtWxbURAYIPaiZXs1
Db7QyYKdy0XH5P1nSvb+6jTwdOoOW/dy91/Ii3VwstiinVVzlp0HbJdmcSEHKitiUx/IDhwFop7k
zaY4h7QaluxzpwFIiYW6ghVMaAQ5B26v/pO3oTSMC3KKm5d3OiMwhsHENpazH7esNQi+p/zFRajw
k73axOMrbSgM0FkHnVCgIITL6QWQ29nzWsrV5zjnx3tX7E/zN+aTW+wZXhi3uSZfI+K4Wlfiys6f
eevZay0MvZeOG+OHjhje4sk//INFUnJ5/E8pTXSJjRcUEOilffhCdXT/MjFZgXxYa6FV6DrcrMhe
xehXhidXhaF6pxgBzAJYWsT04cVGid/0OdfpYIvv4n6wXNG77GiBdnsxp+uXfQ3WG8yKVVJswxPi
MbnFm487qbfBipsLcUwTzhFnK6N9tblKPa6pGpIV+hWW6lZGs44O5eAsHjlg4U0Q+Oy0wof5yak/
ZCt4gnTrHXsLlv/0wghULYCAYkRGvRKB8QgS+BGHjn98/oRJcuzXB+fy0Z9LeZBbelOQpTL/1VcE
Gj2dKgsjmIghK5a6wAmSHTcV6/Ejs7c+07uoLc/YSWXv2ar+AkfAll+GLT7/+n/BtFsNBvWWYcXy
sXFF28UJFyiLlJDGploZSqL038Ar2kT/aPdCobBRiJUR2zVnIPOicU7zoDOxTB4Kud2x97P7btYt
FxP5qEOWcoeT/wkxY+yD9aDSzL4Giyiijou+Efmblr4LV4WicD+6iVeUVfc5AiTYxjpej48nBlag
arDkQhtbDQBzAEq764Orzq1trGnecOG6I6VLem3II9nSoxr5ULWH77DWDFjk7t5blt9RUS277gDy
8/k06vCIE7kdHYUnCE7HSQWlUh4nTk5E0z7HOSfrDn70jbJ7WmP4e8kNgT6VpiIpLdzbrL1uUN9Z
aCMPV+FRIH0fo/pj/3uqyumn2qAolobo38H0s4BSNZHVmlteMNTZq6CJwqGAJPIMVikImp07CRRS
dUq2+Wx2M2LxanRxLEqZI+O/EAjFp6bHaDH72jvqE0rEk5k+xx0SUu2YNVck+n+/HHiy2yyr+lKe
gDRFID/YWvwdGxrZov3TcwZdfP/deDgmniyBx6UsoRZUnrjUH1/WWBXr9+anDEwEjz1nR5m3zZIl
raUr1waISGZs+TwWCOW/VzGvKJ7JnzGB9sSXdq22yPaf42UiOVHZEX9MVe64iBLWNfikEVENMujN
tUXHCct4tOGdfuRWrxBeWGH+IpDfhYuVZuLYiVoUVM3wdldoeL2g3qjE5Sn2j7VagKH4As+1+V69
xrQoa35NH2kKQXNikYqclhKxJGOh5b6aRmlGxwO4mFhe6GG9BJjbVccSHYyM1LfsR8EPHzsAdAJD
zRk7awuRNa/j1YtdslIBbaT0IHGAcWtlQe092CZ3qJm/5oKChk88JWfBGpjmCQfFeaqVdC/PMaGo
LQbw7lV9AjlkS8Fyf7bvtsbBayYe2It5XSxvNgi4drVInyS1aHSCt1PXFus0yYhv9OY/cGCvxIFy
tEKLsohbu2DrM/kfgX3BDyq5Um3BpXBSWDQDPHxhFJwzolAcLGMrnkKCYi9fbrg/ThmOypUL+pXQ
os5MdgltlKVgm0xk2uYNUlzNCVA6KvcqfJNNdUuBxUG0ZNfnI4muKv8tDUQIkph8wj+3isFdRqzW
FdfUu9c44ObeE4NlefJ1zUiDelcC3n0wliLJilH/SVtuOAWAAUA5jpMeEfSf24r/AYs7h3K/Lm4i
o8E54684nAMAj0aMoLMMMEY1zGnn1JeKSYjD420xpI8DYQ18ROE6+JlcDq1fwYUsmEH/SkUb2IAD
HLdfAlmttUXQB7yIfrTYY4HBrjbbGpcRvouyCXcqXJHbeVSW0Ihe/Ri0jPRYD+0cYa8Tq7i7Cr4F
LXn7FdBJGiFkyQ964k0NSMyUj/dmYTedxdwZ4liLH8FoIdFMU27kEPnSA0sMhiSFOYsaupucjjD8
CuM7CyLEzJ6N59jMWLRsgrvWnxltFA+BZrAu52jvqu2Xy+SgLNDM5Yft100ENxyqD+AsTrJ8TMGg
Q/b4HumoKh0yMFb5e5fewY51119YQlmYox+M8zRTWfmAOhWwMBm4BHQRM4tipkVkvAdCgU8AFeb1
2pxsxi/VlwNF7J+T1u//VVYuqvYalJdm+swwIVsIC3LxS4jcOazVV+hxP5Qjs0TukaM95VgfRSMl
+WKlR9YDPRpPNEl9aCpiS1924S+C/CC2PBbtuf8Ifrr7sxOGRHYXZ2FZeCzFCKfiZTrcfJCwQOMX
puPvDeyYYt31FqAckL8NmEdUnwEbkvXuHD31lU0p2E0hW3H3MNlg5aMEcFHn4qqxsSLFPmjqrAoY
pSGEbb0q5q9OFMtXMgLCATdJjQPlFoy2CcrpRW5H6mJakwgJBsZNDg/r8HjZPyFvK5lvotjMOH1K
ubw8n9gXO9YWzs/EKJFvnGRNFVxmc5b34rQVlTKh9bt9Vgcw3Cmj/EpgkE1ewrHD7tVZ2RyLekUv
PbpCFthQT4Ln+g+zu2v2YjaqJ7CE9U6BePxIFCi/4HxgT9vMgHC1T8tk1LZkqXUkedc3Ll14ZJEi
8LBG3cvrG4FoNiqTlUJQd6va4OzgKtgSfw/+KWZAq+esIWZx4pitCvJhQKBbpnHDbBDi/djlBv0R
7DdTywdjzM+rCiueJ5GLuJmh7bZGGrVSpIFGmMqvIGX4vmYCqbL4V/2bTgfZmWb4XUzSYIK4xS3T
AgCe02Ys9v2SkilqVDqzFwQmy5hIhCSMcEi5gxjY2nTdt+lR14feAMgCClz2/FmV3bJ8pLoOxfks
8Nic431RCipBLeK5Wz2Dx7wcu1UC8y7XN3hyQ5XoBz1RCcKGH9d4K6Iwd0NNqt5K4TNDgC3tlaOY
HySNKFzA7RwxRUDcs5tCvw+Z9485PGxlMb50XxiqTQEh4b8GSujeVJUhcRbsPM82RTwtyyxLDNr/
Mqqc/8X0jYbQ2HnEPLb9vjPHnk0+jD9tYzrw1NlAJoc20dw/Im7rt07SdxSO1lDP3M/eg3qDdNPO
+Q1TdTdz0eyGe9j0A3DytjOhZyrFV03t5DJsVAjQq3mJ3EePN1tblNT8HIYT1j93Rya09/pZtuvu
mRoKLj7K1anGu2cHClxqh3/BXdSbUscL2QDQ4ox3hMP1np03kUG0Tx9zLsumw+EdlA/GC25CuaO8
Vc0gNDDMu28EOiOsdZIV8QfC2Yq/czjJTdI/ez+fYafhCIba/ScbYxivbMby3h8wIYvvTbZqFAme
HEnk4cwXfhQ9c9GU0/qm3ci2goSDz6QSQw7W5jgoPqnTh7/OfAXezfm04zzGH//GqosU9umfDOa5
FfQ0ovYUgAleMOcYRiNS0PSZ+FdmT24UP7XPLKOX2XhQvSNwGGe7CRqw/7/fYkX8qBZypOuyqps0
VT7hz0AxPLkAsYCRv8RotHhDCraYL14ZUTdwb8lwM+UCcnMiyhR7Ns+D/qHmY5oJ1qbluNsK8x/k
eYBb3ztFuC9CKPdzuERuvK9qPZWbVxeAIIgRunOAdsK4xpsC617Pz1k4tzB9+nHtIyiSqmMSHyAV
5DO6pIpsPUPgruSKp07uLMHFNCmy9jFE6ohvWcr8zD+HSeEoySrsHgq83+RdUqCRzf18PeEmAmzw
yryWF6Szaw+Er8KqWpM6xhcZC7/9vshwdxqRJRTKp4mPTtdbt7Nh+NDaQYSAx8wukSXpWGy7bBBr
+Et+CvmnjoFIoBpZ5u4glDENCLrRweOm5yrvjPlDb2k6gO08x7xTSajD60usK5CEaDKcFnPCqr9t
SjTRcCgvNqvKjORwobcfTK0WTsFJVZVF5UXof+fa+0E76hp2rgkMeRX6gWMHtS6N7hly58V30IGr
QJvsvKXzIFizuo0lir2o9BgsoDYI48sZUOg1lYyHJTLXJZo798+iCnPrxfamjlOZd86h9s+gwMJX
/C6KXi09RwjgVnN556FrgNHqu0aSGKpdzpUYY9ioZiHwKDDt+Vv3Rs3vqvdX4GiCjfTp4XYaGq6J
gOa+ikOHMHSuiBcRLa0RdppSOh9QeXgrNg1fXcjLshJclxhLTG73RlEh4YnAsMEBYowRsHfK1IJA
nh7DuqbJjlbavBzxQ40g1L0kWOcH9ZKIKFE5su+Bh8czE8ylubstmcyA6ZpbmHfNFFnNOaAeipN6
8WFUrQlXMxWa6bNtnKzyw1gU5TobQI+pWg7otLAnAjVxjk3Q/T56S4jJDUN0enziL64REaXzENLf
zbrGqA6FNHw+1BtqLrssRbAUBlNmNlmGV80AvggNwUaIWqC8AaOs8X508qyhB0ChWnd9lRJHNXsb
b4k8Gh3FvhPJoIWekDfnV0LNOuDYAasZO8JO3J/RqopkEs8uzqSKOVnyRB8P/rUdWM6u/0P1KuUL
APQggUkYAzSDwq8eU8lApx6sFcaG0fnqXHgIDLqp3uG4jcxPKVBiU+Bo3HToPm1T86NcIhqlU3kH
2ypXlx1RVGMWN5uhRLTmprb5I/z88NrI1vaqyDQSBnL2/1cRO+aNFvP9BxiHfS8gYj6tF4mCA/We
VJ11aq0tdDtpEPPkmGM6m91owqiyisjbAdKsAfWPgLaqaRJJZh6popJDeqG+NxpkeXGOIDEA1bzH
Q1CfxQfhv2Xa/jBYEi7kbSdDx11ir2mAaQVjjlq5zGiJ84/9cl4GSOo1FpieYwIzeLO1nrS1CoMK
2f43BNdIRXf6TmJkHbc1rs33KAugkYFqHz61ci+iZKOrAjPMMZPUyj1mwTNIj4Sa/K/WyMyfRfNn
MVup2XbK563ql2ByPA8PjKkt9PUOxUPW/3h6psWXNdd96bszzkv/gncbi4hJJ6RRNsSCV2R/zj/r
UpkmXi9wD/KmfqFAKazidYZElm5m4bJQNpl4WdpZKlE0woJdZ2jYLBrGGnwV2Guaq3xUK3lCjFRD
/BO1/Ip2IGw4ARJveEAqTbeIT/waxzeRPz4efC4JP4EbaxtFQtExERtTQU/Xpz/E7dMS3aYS8XLV
DlvIZsfHGAwd7r3JjUSr7tJGbgkAkRrfOg7IH/lUgXdJ3kseViV3wr9BE9NqMh5owxbYPPByvs5h
Istwl9BF69+9kDt29hP13XKhyvO8dRzUfdhVUfq8QN5X5Bm9GR9QMgKIUuUcKYkbYjjZObwmhtOq
qjEaxqnW4Jn/Sk2FshIlhKMZOL06nm/0iLpKT/sFeNZAWJl6SvUVs5/r4U9nw6JR6AiRM+El+tmX
gLfX36JB/2MM9fHcq6TcjjZtvbxYFvERUeg8rtFmMoWttyVReuH4MXOkdQrVEVZUZNHvBrZxitIC
3onCvQgHr3RTSgtUsL6BnHkBXnRsMqUdfyYOEQaNe5HhNZpvkilXmQLnMvc4Hj5EBcJTIhrhLX7J
DgSRirBVnxJ5AAnfmsYq1GhgLUXLFZdNbht4JWeGhiCGdS/1Sy3uLEhXdJQIvifnQspVw2Wjr63y
Wf4Mlt4wkHyjqHi6k+b441Q8LPi0jeyF9EK3uqtZrq/lPKbO3rjCTF3hkOU1ibHpx+vtNV/dMhRL
5Og861r2IvTDute0E7GEfeojjVOr4FxCrrkAXuy8FG6FOXRVIAhMNC3vXZL1QgcqiYQx2bylt00x
q/zVcBML6JO5Xmqpdx1KSvphoalTvNMNfI0nSgtEp0U0AQBq03lKt2uOsRMJDCtasvoi+/TKnSoq
JgilpugUENJ12Xdv6CTA9AWKJ+FuGsEvds0xO1Cjub/M7m5Cm9ev2RxHX3ZDaIXbFnaE3y4xWb2a
FQ80RN84xg384NjLNdkiWXH+uRUMIvQ9r93Wxs2nyAlclBg6ZZpulDie42EmTEGFXlDpHY0mnHRY
rQSqEECgeFh98StO2VnN9PUrbydST+J68DUWhcoivIEDPvADa99YMEYxzIL3BI9VBPDIz9Yea4/1
3SG24IlNEbUVtJewxbANbH+hRYriVZeJsgL2yU0zouE1TAFjKUFfR/jtJ8d1rfqbo8NrvsSQWsCG
YCiIWcUAtODhlDiyj1PVoBYrA0hLdyacn4ZqXnpdznojwURkBazBBI9eLwMaP2Zri8yBPvdDpw7O
nSKKGMj8Uzf82UFl7wX4H/oDLq/OG5y6peDr1Hjum3rPngQIYZ/JXl0Jl+X/0zkyOp6hRLXBkq9g
UA/Mzte/b3dcfK5vj8yDDr1tQCeBVETG1hVnFMrdF665bIifgM7Zesi3gBE7rNlx1hq4OhkojppC
W/UlxvPD8lAvH7eMhGhJrhUlc+ZaTwq8BqydZoogGPhR7xYICd2Qau3NQcbepyR8wTnmNkwcebe3
J89cUz7eM68PLkoC+znw1oZJ/8YPre8ijhzjINyXjSTNJh9StEYf3jl/WygZyy/1Nc1Wor2KPzfO
AS/S9SMrCXjZliVZZzCGq2V1arVg5MS+WRypJ+s/yarmKiy4cZC1z5JYY/cYT6TK9khj6BwXS2lw
2Kj9AaoHSfn95yfAZetxQ+xNtL48aCjsTPO/rhZrcmLHI3W2GL1a4nGZbG32+m0XYRZ94YWj+isc
v8MEaidy3TLacRIeha8nlXqorDqphCa246bX8HunT9866oikYAT9t6J+kF8Euub02X6yobu5r/2z
vhumYKuMXTo3/NdunDoMukXMtT2HU/8bBemk50bxgZW+up+Evvbg6a4z1knOWERGZ6HEZkkDnhuw
WYAHOnZvTp4S4MDjPx1QrlLPT4mopvWiWbt5pZgqo49OTGq9Q2SpKqyoei7Ms42j4o9ZZbsxwToo
PxagOdy6O7LV/CDA6VK95yn4155LALJ4IMn+S/CJt9rX6X3AIMB/rnHsG2NSsAw9edk+X4u84aay
a8/TYBmmmNpzwMAIv+ZBvxPnjhWkrHSebUreAU8Z5iA34aeyEid8+4a5M7nzBLyEvCNTunH9w2aF
9vFsW6eZVPEvfHkslpquIS09HXmJsy+OEs0ZASgTn78GJJUSUXpeElRA3pVVx/kRydUrEC3vU1f2
88FWIw8c3rOj3QNnJIEx3SFZ5tvD8718R4tEwdS8cPTfuuyA0w1jq7qQUgRBpABNpafM69VXD+Rq
zyM7cfEX+ak6V9VE2V5JzMYCcKutGtvAMaCS2LaBlsNfxShYVYfCM+3iCEfa58aHgoKbaJc/pfpX
x+xZWWpdi1suDxkQpojyNSnmIcl3+U1/ylrGSOadX6RCfhU1GN81IHt8bedgr/3litJSwR5BAx0d
ADtFcHPXhIZF6e4AwByyJ8ZSvBbY52/4vWaUbiyEgvirfp1wrbJl1It2+38yv3JuawWH+gS5tj1U
i8b+ANkmG+aBTkPBE/UGQjE4jj2vyQqrjyROITs4hLUd4ECnfbOXEsfLxP2FSCxtYThqpnh2G+eb
i4Qax8bJ4YM56REJemQ4UcC5My7/N3LEIyxSeq90wnFOyOkiTTf6m4hI60ciiElGMC/AmPNUIqqF
qkJmy5VJQh9npus85WlSZk0jSIggunjtpj9Olrq11mlK8Ys95hjrs0svXWLHX0Lg4dk/klaMrUpD
xN9xtkRpcReCqMFnHfmfxc0/TXkYdtGCwr3phfyqTS3kQ8d0p+dxomHYjovXtepSbtTPecGkX5uM
IuxsgPuh0BtfSBqIchd7BmLOwjEVkRigtNXXI+dKWr0WuO3l5xOlIe4mxbBZAawVlhKAHMQdtEWA
Ct0soN4DmDMH1+AZfOPqgYzaribmBTgpqyE89vyasaNCcaYt9JNjKRM8HeAvK4SZUhwk9pRrF6C5
onMCmSSTwEc630j3H3h8RjFGoUd3FsTfa0Q2CZdtZ8+ZduMv0loHDZlq32copJwG6TIRPS2//njS
yr6c+etI1CcECmyC4V2lMdoE+01p4AkeI5yYbXMjJBIqeiOZ/GcHpE3dZxndXGuSftmzbsHi8NN8
75COTl+kTcZmmRztwUnTQl/QsuKfl4N7+yEmAs5ntaeBCjo+mLovc4lPN2+EcJ54lsK3aPHCu0xf
+u7q89/7kqlhz8YaC4eBuMi0Ag/w5ZfqD4yGnlw5EjAhT6VJuJlG7QmFP/uLVGaE8HERLuIaETia
/V7eFsDuc9IktSGkftnHZYAhUyWlh2npI7HqAsuZuyP5mORlW8wJkCLZ5MXzeeJLpG6cncRiNPx4
WiKN3jxgCgtLgV4sipPy0jkC0H1Qog457ZuSlwkLEbldOWYc8OnuuWhv+HAWryncnMl44WDu8Nwv
ke6Nc4XVn59ljk5BwELcJmp8XvESIPtnU/hEdNgb9snc0SOV/dWmDqfIlansXlh3u275fX55osIb
jdALKLhazAEKZ1c01AkzofrU4TsU2uSobcEQxq0tnG8gTfiUU0J4OaEwngrBDl1Fm3OY5Srj+p/t
MAOJTCzDeEeS/gLfpuOfG3hWPHf91wf0hdMfimd+vOyA6NvaunkA+DvMjMVn9L4cSxa2GbNUZxum
MAnvd8X/BaozzmYOYTJLK4dklduWlJXkaEQOyfboLb5qDy/zPcerMYOgyBSLSehNLfZOEiA/0Nke
SbP+2O3kSgWAMyhYEYPihCDWFylgtUqs3piR6VJofY4+pVg8hLv5g+IY7JweEjf45w3FFQQA499d
qwd6n3hc/O41TNAaLdluTY6ZROb7D940WZJOoQTkSjmBvzNGLNSMgYx2O9qpezSlJ2aRxVfUt0E7
J0q3nurKSbXh4NEN1iKS1eHLWyuxtYPGNuBYkoT9lijyRCgNHtZV1S0GUI3H99rO8RfQ44cpTGtp
nLVw4DA0Xc6cG1+Jfx5wyeqJDsXVqUBUbJGLse0Y+lPd0rnKonhh0r6c6a6XlFbhzeAORx2XF8h4
Z46kexyko92h/A1CYecAUCDqdGOmyVecMeLk5YP8bNjsZaed+UUdgS8c0gQNH8sSXBKy9KdyHDeE
JdKQ+s3d02BpYnkWzVRE0HrePclwxK6bSQnrck1Etc6rIljje5Lx8Ls01hwL0sg7ZJAbQ393v2ko
cgbagA2ZhG5V+ESKcfAK4hg7dZCZfZB9hj1JXOZXFgQJTTkW/1dH1+ibivZD/C0RsnDl5hZD5b/5
ViHSNWisogtM4HlTss2m0twleT6N0sueMJOic0VeqHu7FznzZatAwWcupDyoAOXKOrNMg+g4Qjtq
dGFJJcwjNEg8hQH3OpGO2+zYrZK1w7dC4+vObQX6XueKKpuab+ACMFeTotseVhsbO/c69SeV9ewN
3IO8a2AKsfeMTWNVefH68PChhXopL0GBFee+fHnEIT2z5tO2kEVbh5fhXb+na7Q9jVMqWao93+OB
7pyJBFGWKoGuyJXFLp6Ua0nEgxiMIeKd1oqDXvGwwDUpZF9x8bnyJnzGvfR3hq+vehIyko2FA6cz
BBWUydWEMwyVN99K3IXIPgUsQHi9W60xx9rGoSNsbz9mokPSKOBDDOEv3Xj8EiRgoScowBZ+mDG3
kDTBb1L8d8rgmrkfNVlRcU+Mr70UzK3pZVbyHOAk2Y1oOFGop6q1N9hMkYzxhuzUAppdnpZ372WD
UGsfnl9KZDzUCANbHukZeVtJqUs/Mk2PsCgzeBMnqjkBEl4GGZajoLMC9D/Qo5QNzW7ixzNWTHvf
uXCFTADzbqRO531r7jf1K8r/4lDcEjljDmFu1qxhs+8FlzM9fuAAiKHW1lldmi6y5aGT9ZsAuXHe
9Qz3DGHZ+VgL/pEn9DSRla8FmrMDnHZavzldEgxqm5XKVItOoxrekq90HyLRyaRI6OmZfxKeGjcM
IvXB6shzy7aDF5rxw0zgmZZrG9HKaJ0borcYpZ3LR6xsG7jkg0amvSCSTMG5NqVIjcBrrPAaGDXI
x3CCiChw+cR1ZfJsgWETqkupTQCL/aIJfEX8Q3CINGuxSzA+8b0aEfFEqkTht613DmF+a6sJqfNg
SoOFmyOXrC4RyQ1Phe8B3UCpIw5EsF3UdoPtoQzZzJeN09S0VV+UAqQlceoDf6V25CNBqrW0A13J
Vy0QuR2Q9FqFqLqmiUku+kgMqrcAnYsGn3W3yLhjIXfUNAxOfrDQ+ZTmE3f5kybM/7AJOqOgfEER
nga5aHp4kYYwmZmy4niCJMD5oGXzRwxJ5LJsP4/gzSmM2H60+LCjI/yr4s2EUJqwE0Y0xb7sOwEZ
Ld1xvlBWv7J5fHRWm8tXYgcJbJ5BsxjRDkw0/YR0YFsiLwVxqw3PBEBC3Yz7Tlr/WHJDXnw1Ytg6
dvdrY48nKIPqlZy0ZrRLQ+VnpwrnjC3X3qHasngk/gR59db/SSPsrmwAbLbpWl6RW50wK3JV1USi
UeKb7xD7cjR7nNkI90Ug52ITm1HKs5SedB8kwMv66KR0O5B8i7fGUc5ltcJUusLd8I+k+HpDAx9X
YeGBCE+PyzNFSVKuiL39Towc8uetWzK+URpqj79Fomx68L0YuIMi6ceq+M0U9G9ZsfOoNI/Onw/U
VAG/STsUB3xprDZf7cohPUSUtGbQbQ+btcIxhD/pYJslSXLMnKvL9nlGfrKM+b5TqkezYqcXjkOS
cZLcj4ZmCCszQrn8LEQuqmkukbKIMlX+FDScoM5UVP5txnLPl7tHbOv1SQa7SUjfNw2uABfkRdzx
sTYDpkyzjwYLqTNnFDOd+OkzWfKyIG1iaQ4RlVPTzhoq8e0pYjoduLu6uQh1ouEMq7XjsMZgrN1n
vcSx7Wb+lMSomFTw7DcUimcq9mjICjYv6xzeFljR5kmlupeRMiBCYROClZc+C4GNrpMszosOXETf
EhIaKVwNb7GrKb37N45kQe/xjKypJeiGBRtoCAnKkEK4syTabXlo9exnC+n2CeVGLEY60k8Pm1nl
YkIn5r7kb2lWyBTVS5KdYrbDS/s1coU9yD8AbvByZ5HrUCh51tRCEF0jOM18M0Kre32iBk6LZKFC
WET2geuZhLuY5YNMa36JKup5jsdY5DchUpBgX3Kne9VhEmdlLHCsIy5IK7zR8j3j2ig5Ei4eIP7b
BbmPXsIuPh4JZCVL9i5vKzG8NXzE8eAAUc8M+eNfUNMpBKz/Hl+rcJ76g7MNJuT8uresVLKnbkxb
DvI3sQpNbTdNV+yNQHxqxRz3i6c28o1nzx2FSCzZjlzoNUBkL6clSTJyDSw5cHhgTTDbByE8zTVt
zSvEqtcNeuhaSf+25NlvWlJia/yUv6OkOK040bkqbDAOSjcm1ufrvtCP0wqTTABw5rSTXaLDQAF1
qRa1iHqqYLZY/Tf66bjJPaRIkpLoBA+5pJW354xCNfp7sJ32dlCIRg1lmq+1CkIsnGXvF7NR2r7+
2VqvATSZVhmSAo/y2YX3m77IjSUOD0kiY8zDslXUWgXIWFYvkvXBG1bxK4p+ZsQr9SxpVYQvvg1D
TbXEFH84AM5lBWm2WyzLNTR2LPPq9sO8DEz6txaxP0V3Lq6k+s/Bd2BXtnaDvyfkTdGa23h8Bhwc
8lKw31M4E/O0E/Xx1TusVk9SCeO+ZwzFhruStgmGXokgbFzUyJLMh9hAFuQbbSzZo4Qf6iqeUDWG
iUgVzE/oHoe2+EvjyC00FsFeo4p43R09/8HdL2ZI9WrY8Q9EkrmUcHtj2fKRczN0qoWiJC6x0Gje
pboTT+4dj8oYMifjNSzIq46nyTJkgpIO7tZvo8huEYA24VxrAHQ01O3KZedZCjZQp+aPdlVIPTZw
06N/c4eDbcuwHwhierVb34RVH2fTz2o0p0abr37cHM4UEPnkapo2ilZrVv9lFeDSyOgFlA+GY1Lz
loT/E2TAz2U11LaAz9OMBNVpb89huT5wb9yxrPSrk3hevZ03gAlXJVWeKhARhy7gZis4ztxbrCZb
c97b7EAJ7J3V/RuWQ7yDiYY3kos5kgFQjIIItAOI8c+rzl2ehpHRbTKnODPMomJwWIRFRWCUEJFx
cCk3vzAm3RKcfeFnjrXGItgW4dntt7szPPGl30MF3jmotke8dY71GFGWMdpxNl+YSNsAriUlFLbA
9VAptGqZJggjxusZ9YR7M1TEnEx+VJEK6uUbNzvwdpAqiJepZhkzGGFX+slyHU+Yt80durQyrRCL
/RbMgdMAYejQfguS1SpfHL5alVxBJG9Py5otbr65UxRB9kzFTpVulI0BIjgYpi1xOAflwPr5izDW
QZly1fbIaqyNrmPoPgOMbLwYOop58nqD+BT6Uc1lKmuoJRtlIiNr9FhFLWK38Q+Zx/QatwX16fxh
MMfImJ4l1KCDaHp3YBNi25MTxTl6tqB5V74DRk78hzw11Jd05ltdZebt232k29a6jYGTC7TKu6nH
IfBXgiTW8CFXdTqRfdEC23LxPHC8mGapeKjkGTImKwL2XNH9makdbMcwL0Q9FL6EU0j+YSCJbhg2
uzAgftCuYVLAkqdLZ4ZokE/OHO1F/ceqL2f5y+iFF6UhcyWSkHMC3ukVa+kWzHnP+9AfJhiqcz/e
Zukk2m8GRXdtpgWfvUsZBrrqgm6UNX13PRSYGsp8kaNDUw53LiQlw3zGbki/8qkS+51UtMTGg4OP
uDWQpjiLQni+JPejSdCuqM1fzc1CrZwgvhBEdfM0BKjEFQgUypD2HJL9nVM75iM1+w4FfHboRkwz
bczk7q+RsU3rdbqp8zkD/Og6mbEX2eQ0Xu9nK2qdfM2HLL+ZSZodYSuwXO0WnB0U7c7pI5UmewtQ
FYe002wZF6l/UJUI4aJAZWV2BwrGt+T9DsVdB+ua94lSH+GcwlFZWsHJZdmDPZlEjc9qr5EFAAqB
P0Rd1Sjmv1s5KltanGm5EhJVPeat1vMyGqsRLp9ZA25Hqbb8QTpTP4yYxnprzGGqx5zdP9FWbl4s
i7hNzxT1AhdQ4MDsdT5J0xm5PWk5+eQowuYXsRe97iPWwj4uHYDIfRzHXo5lwwxrDGqRCf//zbSV
ZQcuoGuPwUGONv+52E1mqgg21j7Gh6f7l80uJCdkWJ83Zqlp8WAIvplWM3tPIJ83JLk7K6Uljhcf
HINwpP+EyJqea6KTUhY8Fj11SRBk0qLi8JkG+AGxXR3t/oS9QQRdfjuSS5gXYDYR0fYD9MGQoE6e
c1HBqfNsfLccDQaE4zTPFo0tI1HEoXiULDG2qPj3EPCjhb3yoai7GG94fD8jlXzHPkByTMac1hrT
UAk7GKCp1RUgjjLfC71hT9TMVX2PR4gd70r9H3b3BC98JDRkiQ5oay/Kd3foWFrk7aME/YprSwMk
Xhv3zNwqixjCmIhjg7R8HsML/6lKx5VBlVWPnY8ugbtsPQZtLWOzXAwtPz4mWrJBNabMUeeRlWLK
4RupaYt4pFu17JXBT8vxYjfOVng0CRRmMyxt/wYi6Av8QwsKeE64Zs/OZA4qNqIZYY/wWwa8ArZa
CpZMGCSfD9CwcMj9h3sWuIr40pJxuvloCrYLMb5E2DUaPTV4eY6dGoaCXISLPpX+jJEpPQm1640i
ocx6A9wZFtNmL+04ZxMj5iT5oprEDWzSYw5N29U4/XhukaRn87IEVUYpH71YxN9/Bp6fzWibHMCL
XwNJOjTjJpJiOOQETDqJvujSzOABSprb/W05x2NuKHpIdyle29/GBckA9cwtQUd/+IP5wD5icCe/
axsloaWl8ACtNIOg+sm3amAYMBywFi8Y+is76DSK7AikV4d/DDD4wD+ZOGb8mJSgocJKkdttwFCN
+r4OXw3330IQ6RMDvegKCn43ZG2r3i5GHH+JOK1whmg4Wx+yH0gwikjYDUBWfUiGmMULwEEyOtkW
PtE8vn1X3v7ri+MV+0kthJB0opcC+fRjnyBkJ7IiBTN2hxCHt504XJks6ixZ00kgZKPdgdRjkhm/
L/sQWq+ZIm6aOVe1IStoWYYGfKgCyCGmRyEHfWEYOWQXuePptFjvdbFMCEytkW6rxriuczByC5pr
IsojM2ByA370aWvDbDdWr9GZ0RZpxIA2/mWBiSwrNMn0hhgoElonuoKeK4n6boFHSj0/c6oFvXKN
ai8suOiz+jJCes6XtcOXvFE2JIeVA9t7NcaFAoaygbcvZ912Qg8G5hwpX2NrfEFO1NkJJLrL04F+
4PzZAcfec4wgNHrwNMR+tz8NVYJ+NdXpzrBx4JQ2mFKN+PluhwSiXGuMoXGo0y4nznGQdMKJ45YS
pztpvf2F6jiRMGmGjgmK0vzJ4qOm7ngzCgZMTGpoW4n7/IHSldFOy/9VW9bhIn1zy3RCB+8wLiBQ
lwYKFYWjj/krCXufFzd6B3GLD7RwaeiZjMqJyvLoHMyJn/s2zrsx/b2rcZuFUqusINeH9RiWbtBg
KgkgfcBuGT6P1XPgZJhoTW1BTawp+DhdS1vDoOinG46s267zz/opatlNAMf8SUesv7eiqQA2eYfP
Gr4Srtl4khJ6AN6+rafL5OKCZBpYqzyWAVSyQF0sp4wiHVQg3e8ZcnoKAY7naieLi8cD4JnC0c6t
y0rSDuy/RvXtPru4yX7KJG4hti2XD0XA9sbp9yXg+93MpArWzW3cYPI7o+x5aoLnXVgxYItB954+
91ejSTO8qCmygq4w6KWiwKQkGeAgNpjHGhXG322gHLzENsz6B71z3MDtCHc13wErDbi2kyUP2ASU
PMQtqks79L8Ddnv8KlEDo/M5d8uKFOZ03s2x0kre6+VmC4lJrg3erplMHZQT1ztil7Azp7jxW1cS
qJCEfpoyjJCObPyYWZl4dOifq5B5EQQKHnHAIOrBQ5AcTn/odN/KCNay5hgf/rQq2CKqjY9TexH1
nh7FkHBb7V9m5rDohT2YxF0Aeixrcc6YS1WNEhtrx/W1n+sJHSHzz1Djz4K1PO4ZfJtegdiaoXTU
iZDpBCemWXR3ItZlFaxqE9mmh5CqjvVLD73+rlq/WJ2H09w7I8C/aSJxDRqgYr8lcKNt4PGuGIee
YDCgYoPYXqzJIUvh/oYXJA4qzvs5VB3zLKAbis5Dr0wJ0dUXGXSIz0jL3vPslAn+ldMchCIGII7Y
yo9J1Kx5zJGXmnKrXDes+m0YuZ/chhRdQOTHgtx5jkmc52Helom+b2m4yf5d+oUacZ0vHkBuVsCO
lNWvTojK8qLebF1kaNUb28JhyqL7hiJOMuJGQ9ND4r/4sQdfV0PlNhxNlSihxT18RGvjaOamd1Cw
yG8yYhBoTcJ+blJFtJRtLIVSXjwyq0Yn1lxDIrVz3AUFZKvZu/RMIAYdOb2GMHHzouwHP0Mhm/HP
V38Frj8/5P8uTQYvfCrfY704t0Hb2fDXPT1ZIHCg4DMZjkgK+klFezKo2XxibRKtP7rjZaehjjYj
vQGH3wSBR37Fb3q0TkwiPNiJtS+RQ16H+CZemgZo1l1oaw0KfQNCXXkAkWhVlLmwS0bTxHKKPNEv
IfnOGpGzlh/rKuQm2I4OCwN8hHb8I6Evfs8+v12ARV2ODEo9wPUJ+C4q3OviJQfO3bEW6gbdU3p0
zEfwtU5+dXkxbX09KU0d9ZkUl1qSpREswC03Wc7X1pPAYmkThD9qPkglPu6wGWo7j8eD/nWwZSRM
N6rt4zWpJrmWNl/J8tswCeIUU/W2GJ929FkmDB6DyxwTqGgRLIT4WC5erNqMDS7zw6KSJpREUtH+
qCw91mLLVgCOGzm6KgEWemIu4M+WSFJ+uMXU18AKLMxDvnGqyxNkqUjDF0H3GZuMzJ0VfElBk3ar
P/M82opz6OafYKKvO+iGl4PjA+y6UaLuIUkT6+bRwr5v17ixhbjF7oHO6hyWK2SVieAr1/OUHTsw
ehyngfpe8Lpo3POkaUUMrG4sjvQSPqtujo6+nW1J14a7rrCVaxMHISA56ICiz92q4dYH1XFcp7Eo
5ZI8z27fFMs4RRBHuJ7VdpAocRQOgCxqgjkU66HAE8PJAc74o2YEJAPeQdjsbHjhmKrK8IXLGf8D
5HqMtEk2+VJMAZCWCbTSQW1zXmvSZSWbHsAJGX/X0d6h/18wfWG5I8fCbhfNvTjfLsXtk2QVRXlB
lK7lA/O6uXPjRiQJOky3kmZ1FmFN74CoeLeFirJZDzs2hPDDnbemmopmQ29iH0GLwvWb4vCVMS/d
SSWTX+lqdvDiaZgoSzBM74RhRFJf5DjNXmEWsITBi9C5fxKfIcJErnu36eKKILEPE02SV2DOguuL
dDPIQOE30nvWOYXg9HpY0KxCObuv5SnZxVfQjW/L8t+6LvnH04OyEgBvD9CqTq7sPbwgCekjhaPl
LSw4spy/etz1XAbuWVujJozULQd9N5mD9FiluE4EedAHUdI8TIRFupFYSCxBMq3WL0HboPBR0QlP
QpMeJRhMhQuwBZNDkodz8LhjGhjiUCWCoo/2R7j2YaGZD6wQUtVv9eeoSMKVKTo1eznzhO73fvaD
R7/fJmOW5XK2EegEqp/42SRX5RBUdIztONCPKBv+3h/L+qfD1iLh7Q++wAa1d25NjRBrSk449L9C
aVsKC69SKzVqXncBQDHLBIkL03ECDlJL3yqCSXYcVp1Ku+uocUYGThsbM6L53Bo5ORRI49wkVyIh
l7E4mpn2hjOB+UIRY6jaJcwY6U6YRap5EkknU2BtW8jIMjLbkDocX/7vkuqmUwbzdbU72OZIh0p4
z+L4Lg3luMI64UlOH80ZgLRAKS9fmRJ+lUZZcHygDmCkNm4lf3zTHysUSZCcFkIYpJDaxicCHrpC
gNGEcmJzX4qvzla3X3qjNqncAAgR73t5D2T2T3VQjYxGLxmocNZZYPP7AmzhyyszgruCZQ9aT0Kw
b/ZFU+2CrtI+cF34uITczEXiCiVdC9NMgKSRPCDqpNuLkqcS7GMeTDgpsizcSim7tyNPW3D5R9tl
P4VEmczN2wjwz2QbuyM7ID73kSp0GxHj+g091O8me2v7Gp+wvno+egsD0ldBb7mU+Yvvrk9VVUmW
Dc/cz+UTO3M+C9ncNH0UkUoW4GOEBRQTj7R+uGKpj/esBpEjYL/wN+jAJ5bwHtYOo4YfY7fHp/gm
t7XDuD80m7UMtdDVVmapqq5HoKCboXneJ+dtE6I0DW+jf2N7FXpJP3xwcLeGUM9f6Br7v91DkXPZ
BBK1lKPo/XEPHB4rPurtn/Cg+Ztdpi/EVfjEAAMKr0/he5w0Cg11JLFWtSFrPAetMp4bD6Z3ZGXT
O39OilreaRpq8DS1mc+mnlilMMqeeH7PAREk3rnGp9k1syTQ8w3XK3BHbXZApSzjZXBqk+ge5gWx
mk2wW4RBHWHh4iKayisXwqQL3tfRKdISv+M37TNnUrECN1diSSB3ozp8rldxMaya0EBMZDopVfoA
30PDmunmdysqzxY2TKYzkjSGbT7kmK0XUAaA1bv3NbobYn92QZtjwbLmVv1X5b6Q00vSNm5IhtGW
WaT2yMvX1348ZxOGkCDOiyJXvNabrNfQ+SXmtqArHg9d+ybXyh+DmiAU3FjSOkV+C2aYA+l1Uetb
v6w/lh6ac+RG/0ZKtv7CBQIrVi+J8Y1Ct2AF6CdaQVzllwB+53hzCACkdRsxGCkcG8Nb6qOJvIbF
WRvYvlka3h5oB1viG0iN2yMGbqHsqJeFMJKMWUdm2I8E1bBsSdUEYYmx/naKKgVKGQojutsfqNnu
BFXIU1DNTwarOMSi98Zd4ViD2Rv0mEtNO3dNGtwPEK8nzCS0QHiIK8Tco4Ge4IEzXmFqjueLTCnE
Pb70gRwqWCfHwjQgyAz0cDrZGT6hdFGa43wwf2fKtUKGTJzFWlFufK3XUOWUapOlMyuNSU0DqcS9
4XwmHDf+bZCXJI5u8E6SMm7f6sKK7Yu+Jj6DmvS+jYIXVPFGzKkpyfyLX0qi1Q9ThUtMqOvcyA0j
ns0nBPgoq1tnBo33Ok9wFC8tZun9qFrscIeFIJbRnCEPDMdywFz73f0qQGBsyC00srCAOZvVzkBy
IkALS1cJd/3sI1aVIb8MlDWzcaZw50jHDw08HVact9u9NOMwtEIVbXtbF5Wp8VffY61iBNNt6v01
IXtLdXzdBA7HiY4uaPkTONfeDa2tpJsUPQ+NtCNIZ6AweXCW3yUB94Re4t+kxze6N4uJE3HgAziH
tVYpHgF8u3i+7cRCQA/D+xpVAyhgrofhaOi0Kl7dYtwrKh9i85GvrpCBaHHEwsBRww3HxpgUQSdy
NkNUpvTGTdSRcaL0PGC3TC4aFNVuvi65TLJdHcC5GuuaylUNmZCD6JxJXhDdoj4o6VcyoRXIz664
UBU9x9BE1uwsMoR1Mu/HeFH9CwFodR355BzAvzxTG9PnFXPshRwAzhK/EhqH/2cpV7lomgBKqCYo
i/t6aX/ZCtWxJRSk3NottK4T7jfX14bYyYJuUrV61Cl9o77klz8mYlfsrjSngkmXTZexWsMeK/Tw
IBIB66e8TjxVFy7qtji6gw7IT6rLYuzNRLT/TL6oVwYy0EfkVfdBrN3e7uLdiBIfuaDMkU2DLwzC
8JOphg3JL+EWjutQHcpwKE3RizGEgdUlI8MbbbCjDog7UrxCwyaRlz+Joidt18CFlNWb7vmiPrnE
biSxMnDAbU0hRkUHRC3DKmRlIX8Cyw7awz8wz920CmTebBCnEOXce2QxIX12bFafnjYou9yYdALd
vIZ7sE3LJH0o+Lvuqt8A7X4KzLhaClsqKu/3OOltGWPnMEdcuAlf+CGlPFhR5RUtE7nhsMEc78/q
rEieZWJYAAjYDwIUzAls+6N9yiHQbZfEXnEl0Q+NRPxZJGmaYGbVTQSh7TmRSG6JGpsqwGQAc7bA
I8pLDXycQrpjsnFxLmrK2BK4CvijI8Ot2GPsEHyOYpEZNUY7IzfP7GTRG8oZsC5c7Ys3QVkBdboM
HzR56fGr4HwH58BeOxgfzB/Lq9Mc6He4xMJF7idVFfHZh1mod2MAiCTsnwYpl4TJ7TMYOmK0m3NI
fYbsvXuRbpMH96ep0cJFKda3kkVjFeZrpROEvu1ETboBOxvPul1BQ6OAeQIvABBP79hNFETPl/M4
YcRsgB3f9Nxqjvh9XTgaJTn6ThuWjQxoePUs4tuig2mFQ33X6eAZmcSqWj4vUPLYsLgMEFKKln0T
vxc6rWdNXJnNd9KTjw9ctFHAFOXU4D+I296WRsSz6dOEPsNM/Q2g5c70CWuYVT+Yy6cbkMDLn/dR
dho9PTVQC/albZ/XD+QcSobB6LXR4C9KqAFr/BJb/q2qSuUUcPLPR6G64FC1cA9qgtnhgOYrcGFY
E3FwzlijqcqYKx48wZGn3cOFLXvA5GVg5zspsqCRD9UVmLAz5KbdAtB5DXZxodsVMql1OViAQY+X
Ywg0Cv2cdoAkx+h+jmrlwOLxvjWTwkzIzAPAQJLNShx89Afja2N1RIiMXQSQBbjfaxaaXmQRXpNA
u8vmxP8Z/FL3cvFISRZffL+9SQMOV5hxabsE5oaoVsMu22C2vlC5k4BrzosVfSllcSl8ip4SJAOw
aBcbHoNSCoxBBuejuYPTYubrZs8ri1iSqS4KpfaaEjxOXntU2Yj0hH0MlEih0LIwGLw1TOV12x2b
eF/B9qVDQtkvpM3dRdZwiy8gjuU1r/yLBTL9pQYHbaVJ92LIv0lOvJE5ptDNSEvc5k7bmovJa1EL
8J8/oo9d60hi8JbHsaVZ9CuiDXdZFZwq1H/485NQi60k4JlWprIGqXtPmLOAvj84E8AvwEeCfTOU
b3pBlxRRwcovhQGpbKUFKP5/QQkI2pt36yE2JgOpnzdXYAfWIARIEOENrzN7XArRIq4dZWJ3swWs
EGHn34JwzYA0/U+6GKOrl5kJTcN1ThZzs7lEU81O5GarbfQJk3m3Q+qDwQUgg9+pqcFKaN1WOqLe
H4+7WWTFLJ45uOPJ6HbGKZNmeyxQJQD7dECx58kbWxi64k3Zn/610n7NVlMwigC/cUcnN4zxlyr0
3D7f1Yx3cjP4of7cSYI3QLnaZwfBTjFEq02Y9QYInIpT7vDOt5KbBgLK4Q7cR9yNemxIynbH/yR4
fo16VfFvtP1Sgyvyi4JfT39sApuRCnvRPJFigT8ekZUZljXWdSA7p+64DQtAMzpH0kWmmrfTjOvv
G9rQQZdbinC3vJX3HsUK+Z7DeAKTFPwNG98ccl1ei7/XX+aHKQzWaCeQ7T/KA4QwDr9yTxLrTxCK
ViSeE8NYNiRz88zFypdEAQs+KDiTn0V5LBkF14KR/7YXHex0nxn3kv2BsKy1XCMACErSGHh1lk4+
v2+R9d+ytYSv8LpYh7NyzEq14WhMd9svKmF+47O+j1ulo4utW9TohCX3lPPlZcV4iv3DisEhom8j
TjS28LaR1lWTztJSeq1H29R2Rvbz/3T9FPuSAaKBBfHF6TUNTeOishl2j/WN1EWIrzRTLLQ9K2Q5
KjOg9VBWPo2+zWsuQ8dQ/LiaGY7LOMJ7tCAHU0mRqHEwb16jX86mHOBhpFuHG/UMC5RR93xVIgrh
XqdyT5dxf7q8GZTOBICY3FzkYS+UZJUmz1Fv8POO/cG+gE4sG1gWL93AwrgueN5olaugg1nIfZlH
reRPr3dcoiQ8wmGxeDNfF9in6Kp7joq7KS7Oa5y1PGvm+FhVyeWtRgs+xuudYwZ4BcFvba4ZTA2c
sm2IdkzLE23WWQ6pRPs0knjQeBAQi1WYve8Sl2QXjd3EgSzpcAoMpNp0NLQyGxn3r5eOxZAIT3oz
EEzYses2j9PMSvRxErH7FvEj7ncqxRFA2S9gHvJ3j5/J3a/zElzRaJ7nhfrqJrsBamsnxUbz5WgO
K+lH6AOT0gyOvaV66i6L5X+tAWFK/8EnwvGs4hEi+lSWu76q1J1EQC5Szq6aPPUCBQ11BXhX7DZu
7CPHFWVgPFPaxSj+m2wWc2Hs3FtlzGAUXyDKxsPHQBKP5gkfVmiVL/GXMZXN6R51W9jFNbfU+7oY
AOjLcMmvJUZ/4Ggpz0VjkPNXvpaps1M41IrofYo1sQorkSBmGpX4CuatPg3R56K9W67Z2/KQfyyO
52sJaVcpMRSOWZQJnluyRe/XC/a6+Sw92XfVUIEQUJRcQVIdKGonrX22Uvnif7DJ0JTUbgbjE43S
mRFZqnmLkpL2KWLku/hI54UL/+HLXZNuNkLyxUVCO2y9OpsK4iCCm6RZyTRIJcq06csTwV3goojc
ZoNh972ddY1EThU3ZQSHHwe8xpRjw6SjE6D7pnE1GSMFG53nxJweebiL/orsUQ+6aV76rdQcSUPo
ilzv8AiN7G1969bJVlw+B8783I6hqkJXZ3WRV3IC1cn9x7Bmom/BUGokKOs0/LflKQ7kGAU+B+Mb
jx6QaDPo9el+zQDQelCLDJ1Nn3IXXso64778oWSwtdw7rVOYhJwgTVJ4V6nom+ZSGxImQczK+2ol
k2rQodEyRDLEHY2hQI54BA3sZYjEEGObiWfoWkSyiqkH929aO9SZDfcuK+Ff8xTTEv/nxVvqSfPx
eoqXBDbWNpqBG6PI0xZRAdqxOW/hN9tIaEfw0TQK0pZQSGUVqz3tWjaycyIbXdoVagGI0kAlNbG4
C9S4YkhVcJwQZ26c/eTmiecp74lTq+42ykhlKH8LKLdcR0BKMjkSFKqg6Fwoxm8Fx3Zl3SjdXk71
rJpxT1bLeQNjG4fTie49yt8lnkv2uu+LIjvCGkEMdjdygixTErbd9DQ4EwWG1kkEcmplIdQNKQ9E
dDXNy3clyNboJ0tRqLcBZR0aMLIYPzg5vsLSOHyULu0sf/y7jDtv8mMkxoFdxAD6I5TQip1MBcYg
/DpHfT7OcckI5itpdYrwZrMh5Q1IkWZDrwqv5VFIJp9yYeKL74IwYgeeAQ3JmCfJtKE7FS9lgmmb
HHX3ZkfyuXHq6LmJkfgduLBnRHoLt9HJMOTZN9JzLqKe2FNdUdieHAyuEQOwjFfOS47gJu64ILNv
Zlz7VfM58Q370i0dD9a6WdodLGelfdnIxrzzkQcdEEsrqa8b38ocUq8EcLDn92XUV2/7WrHbOFWH
/OXeYmTHuWwH2Sa7zMgucVMQrT+fx1gVcaF4F1vQnHYmLLgnAyHXBsE7FhmYzm9WVW2VSIujAtb9
YP1VH/Pp2Yzr3nbMxo2qLczkaW5i4vrcoLhGS4bvfjB9Y8m/itrI7YfC/XJrrf/eYQaVREYpTCZp
Xh7f39vXek03Llwb/grWTOITB8QMxDQOmgg4fjBFKYiOUWMeEzBdu/ctuhErguOxdtV45mR2ac0D
VJKWXIVilTYLIRpIYbROmmdxiYvU9vpCsNw1uSsveLokKCdNj9UVXa9cq13W+UZqZBdW4oSPJBqF
ojE4toLerh28gck0GFknQGXGrqCAqWhPu1k42tPWlWsiJm5J8glfAHMznxBhH+RnPqi1Kututo3Y
wrRznKPEbMtvf96W1iHZ10YpTckW3YAK80AYKMxhiMp5ZNjbIP115wvab+s4l3JISxdQgGekOTQj
kGvsT8DRjKfODC3Vg5R5wJB7+9A2WqaURDWU1m3kXs52HaW2OJU4b6Y83EkNf+WCMvZt48CyUrAz
SUk44kOzKufXYJtufWANwEWQHu5RATyMIERGRpNyugyfXMkrnPRUXW/hZRHzc6xD6NEqVBaU6e4W
tetTKckeCBcdDC50bs4zNrarmhWXn8B4vwZEjlFSj07fV7OuuWKIeLHQVLKTQ0S33RD0Q9oSgVVJ
1uYMvP5ZJuzhRXN43FLUV8/9bZwRAykSzpqlrJxbblAYtOqB7O6ORMdFYOMD56psh9qfJSAMKqwG
0bImS5bEZMPJW14ux52X6Q0AS+5ioomn51C94+PBDvjnYsfkVRIA9bKkQymqHhbkVnDjldTD7Ufo
AT7ALoP6qEHStbD0eiuXduw0Lc24HfmfOWJNnAeEwThisgPvQlDMzdSnUg9kUvsc+WGojX9WZ9lq
RDC+t9Tnj6wP80MwqPASJSMVzHJeedvYpOipjRHrEJLJMu7SIVSManL7eLjC1F6K6O3vLlcBVwdK
TMgdd6Fmzs5jvQFliLMgXTqL8OVTKGYCI/u12P90HaQJ7pAuQI80JzdcY7LK+SH5qDrXclLRhTY1
hEgBuW9NEmWDNzHbQQmiqFPgJ5HHl1wIZFE1MRTyUuAAiNvNahfh+uwcy9sNAxiqyayYXkFPRXFn
6FATiUFo7t+sfd/Kb+EN8IRtfnmOftiaVlU4ON6N+CJSLYu8Ws1rgjk3IHHmJR6Hz9ACHQmcLU/d
mPbU3L9Z++xY1bOwlSGKsE9DrpHf741v5JvP/iFtD/5G2YYGm3L/FmIw1R8wnY/up70ZEPb1ZWic
avVN+kg+Qg7E68ajRbnz7fPhE/QIooOEkub51lvHN5m6nSEIpMzyqF0+CIyVireIKlrkK/N4cD89
GAnQQ4ndQBjWy8ghQJPezIbstwMSuPov9AHPQtBiK9AJY79i/sJtY8fLu3KhkfoGQ42+0Cm9j65K
D17gjh7/c9sJ9kORchIi4m9aiyaO8DUjSoOYxJ7pBf/P2V8iGhUdS8moA2hMoAWVw0bgZjxxCejC
occnZ2+kBUyGx92ua1VTXXox4PEMTk3I2+aWIZ8IwCc7jxELhN0jxTZ6VMRaQ5SXAPEpxt0XzsZS
zRxZKNmCMobj2yGdOKklftMruy+W68SXQUEM/HVxgiWw0xvn9k7+vSJIRvxiBC5tuHxRdRfXb7YD
aeMYO1kUK5kkknxjdCiYrsT8FLYwDMuKoxy5vwurfd5cc04vYiyyuQwllcKduGFz4WC9OILicgcH
bap4vP993n7+56CVopTSz74tjRQIEC4taeROFrLrSj9p1tK+vu3i1k4uum4cfNAIDRpV7xSKcKYr
gorEg2TAum1gtuuEAuCjyixfultMhqMHQ2iFhWqcx15sdkddvkYC9juzkikkpfXaJVXDVmcq8Wgv
Qr59kAYdQskq3qW8MHxMy7UoXao0f9IkO4MSBWUOOqnOzIz8Ed3Uyy9nl1QRj1fn4Mi+50uXP+as
nQ0SjJtCd2T7sugGFZ4slKpTaqaC2lUFC+MkqZsHSqyxLeo+hTiczh9nc9wxBwZ44ZwPnsAuCwXg
MesQoOPV39vnx6SU1QFw0LhrxJT7Qx0Q6Mnk8XetctC8lDrcCbDG2ZbaHN1Gc/WMFduDEzh97Acx
fjqL5goD3XghWzbVmNWnYC3D/G8BUYkPZ3NjkJJuhigT1sNKumvQTbqtxQ1rPINYa+Ke5FukFZ14
nxNgg0CWY/UiJsqA+n/y+QQVprNmEGI6M7m+wUP27X/+zo+SVhuUqY3hHPFMRd9Ykdg/oauzmziN
v38C/Jbqut0VFm2M2QI46A3W6jFKro/GZXGeeli1d6v6Oz9DzsQj0Jv9UJuIyhb/NkUPr3RbYQXY
YYRr/BNsEkSx9jozJah0izyCOrFqFKXqZm155A1L0cihn1g6BRUopNrzZzxM/268VXLQ11fQIS/s
3BIycAZ6BjZD8iRacIsn08GqXRiOil6YRIMopWqw89IC+1JPjRvnwxqD+CevrFSNT3/9HBv2FM1Z
NmCowIHySAHI4HMTDhbNzry/Dj6jJxD81D1La3CneDMLH9wf94dbIk3FI85R0rMidpj0RDcPUaLs
K8hSPgt9YNz0YQIWzLehRUxdDgW43/0Y5CyWDmhlZkVSrDg8WRcjNpsAwZEjLX6Hh6cuQAN9Fw57
f6FNlZ+MLN81j5YeHTVF2pSnRWxJZbO7fTO9yimbpNbCO+SZedspN9hgglQ4fzjY93RZmNxI8RgP
oA7Ss0Y0iZGuvA+l3mFVAFwTkx7BYJDt/PXtfLELUXSiyL/WNcZoltonVSrLPF1CjDK0+Dw12lbV
gHq0hj3nmFiR5Oa82yXFIKWMJpBsX0bhFxQ0+zY+gICsvIzpq5PubfKIlV1xYcYMufDbL+FdIePu
hXV6ksxREJoIAuyiQRHP54D9GVLeN5SLgq+e3ELGJcTgRHdAhsRBRBG5c+Gqz8qgsVG6fJfVm57o
pvMV6Y35hkK9TCVbPNEk99Bu2RpLLHF98B+jVs+S1AdtrBUFwf1FC8GWZt24F/1XF8phU3yA5d70
CtwLoQE+S5ZmMQ972g/+bR6LredhP7EUU5G0oWP0AXCSJl83LW9SKBV5K+5cS32s0tPBoXT5AuWH
J8uWEX2s/hR8CrMGFxQSj7KudkW0hNzjJazfnlXXrEG/rT0OPyEyaCQU4u8dVvKzRcJnxPm2Hq/R
YF2r3wAnsVuSdPVUP9ukNcxn7RZ6nzN43kpi6IY3pGy29PAr0fU9Pj1z57YPO5QF49MhVKfIiE+E
JQ7FRahAE0qMl6h2oCanqv53HTnTT4VLDGMbd/UriOSbmBRK0XCdsAcyT5WbL5C3CJY57Y6pH7N+
sr8JWcVpgggSBcPVncD/H2of02Yh/nH5Hfh8nMhv+llBpcqLi29ZVABxz/IVHeeTeTjPU+r5jW0S
tUs22lHmGu26JSu93oj69BMCK5upZZS3DPCBYIODQjD7qg4IDtStVOTJ0DJMk7orHZjthvqIKkmN
oxpTIuGwKEDIf4kWTTAwbPXjr2/t0N+Mz/610TXZ+cCefZiJ+4FD0YxcQHAldToBhikcvmmPMp1c
cXl+qO2S+BzAfUMaQpH8JOSTg6q/kyhorKgs8j4oEelf9z8TLLTEaRDU7FyjRhO06S34Eaz8wALE
1QPDRYx5KzZh7M2+ekG1MDyI0GdcGRTdptKj511ciV/LEPSUmbD8gYXEBRKgT3wEWz5f9+XRq/rJ
SZOV1H5KYTQJl1fjxinljor0KGWBIMjhTyz9LCyndrjQj0fX+TSoCmLTiaJzXjYF0OOVAwi3xjF2
L3qkGC3RJLBGlLakovaIEjeDq5OvNB5hEWf3lgpT/NG7ucDNp5wujDdfz/J9ttXU7dBds4ymU/Ek
uDhnHXVMoIr2kmOo5usuJvD9hVbqL9+N7zQ2zUzNBQ7fp/YFusClYAkNCXdtvhfzf3SfO8uEy0VZ
5a6Vp4mMyPVHwLxLWoAZ0n36Nw2Wuinf9A6I8PL1HXLGOVYSeCW1qKqHP9Xl8X/xGeNKOu9iqG8E
3xQwl/dOlw6yRjzYuHm/zhVFxXnlV6d1eUOwaDj+mtRAdsvyZHAE5wv0dL7F/6pVqwdXlqHpNC57
izTzU/vyeWZlzC431CfdyE5zM8spjBXF2mjH72OgHNP1XQQ1/Gim16pA7k0/8WGmrzwykafZaZ1N
6za5fk7BckF0frmTqhzCcQKwRqFob0PniGLVvZcCQMpPLzvnGyT0pbqS1tzyUBhu4qeMuaO7c7nw
WUrTac9VoMqFk/HATUO5n4/ArLnFLZ0G0lnrRV4KnEVW/BMwwDetF5ReLZbTaKEHuqtly89rBxU0
ra+f6+HNsmYHsyukLKEk4kbliWs6SHuhVSY3dRmcqwHkdRiXJ1KGhrpUI4fusRx/czJBHcbNa7k4
Dq9v6VMmtaEX6KEWWsX/QXwJqdOWzwvgAc2A31y4gQUjjVCni7K4qaIJyASqcyDaAt3hfnDTutI0
qhE+WeDY+rmuAVgiqMK6sHZHsbl71qVxPyGj8cfms9ioEbXJaSSYa2TUw6LccQMkYgS1e+k9fNWL
mAERES3bSsIHPq2yYDBr2skIM08VB+2jY58kuanC8j9BJi4yDshbAJV00WCndWY4k792je3olDZU
EnkxWXwlbvXERYYeInji8pvlhbrrU2QESKCbk6QvoAxC3YUrIDCgOKOAPSF1eG5G+vEZbjDXEE1R
DZBTCJLjUt9zOGmuyPomKrgAEwOCqIiSJw7ghYsXEaw+ymdRC/llZOaR8cNyNV7dM0DzNyChcdww
z05DX361XIGDCnHw7Wbj5w43mW2Gblb8gW60TxEJs7flS3FXyIKzDLZ+YbYswfn/aJp+646RWhSb
OoYhenY+iDCtCA4A7Oah3sLwtwgcbrGfFs+7n/G0xY2RIVfu87SYG3wykxZiulSJtO3xAY3htOXI
CQSt5PU759b5yY++WX70qpYCszgdQGoYXhF32xZHTo+kl4596ilbNdeVyOJeUdRhkcO+SFDNUBBb
MHWFnZ/stbFoZA79b0NT98i4z+7EyFloWhdnKn55VZcTDUNxSCuUeVlxfJT4bUPZk1iu3U2GdDij
UVVGOykvyXb2BbuIb/jcaYLGw944K775777urjwRgqyDS66wA3ZtigKpCpBytNW6Wx4etM79F07z
z8i04KmTdLUcAgf4Lo4wrXRIGcP4Wmg2M8eKYpk9QWamn3J8KjjL+1tI6HQ8ilKirrd9xwy/SrYE
gtcFxz90ZuaDrHir5J5KZAJNLxriQvLFwKx1l09KHOiS2wNHuG9SXeyc7QNNYe4XJq2vD47MZK0S
KKcN+r8IVAr+p9LZHxWNJndUG43uPMlRbZyFZQpHxCowN5vr1JAqT7zZ2/Xb4Sbnk/8oFPcloZUk
fKEjvckmxwGQR6mvtfbjPCM3Lw/RCWehkEyZQMIzSZanpstC+kf/qxLjlMW6BMmFsjRm/eFV2pqr
QpqceOKMp7Cgmgt9as1qQH9MsRkJ8ieO4mS7xgGVdVr3vY632cM3+NrmAD8J7PrsesuqF7vd2lC8
iHneIYFt+BTa6xyiydxOux/HQVfB7FEq7Ao7KS2PCNNcpUhNkJdFZHrNrSBbhuuYkoIKAwUKvw7E
fn9ZtyDKE4sF/QNaDzr2qO04wG+n6NbrVIUisVkC2zT6YybOO/k9m7wM8zo4DZXTqoYyjRuH/pFq
0y1GS60pTfI0WkN3j49VlhtByuZADiqTF0I+i/HyklvI7oOM6UJOBXoBGDRfoQWj2W3K9sV3xgk3
1wZZdER8lv8ViJyewHCRMfrOmqddW2E3jhw8V1npuKeMN3WaQv9kVG7FnRttyqMtJdbiezDPLSuM
xgmnsZpPYYmTcop5n09VZRXvpRA+PxWNaSyacqNsXBpn+aRkWeMGyBJhat9XmhKMGiwJzJZt/zKF
7Iv5+NRGotcbandQZEyFCVk+75yUoBgmEyS/wEIdtPw+7M+Lm7VZmh9J9DZ9PIHFzVEr+2StME9R
0cBCKcFgr3kkRihnvQwITI56XA8UxMZ8BIPHxEn68EXliMLWgv1u36gxfbRs2D19yXhPLcCh20th
PJMIRpAncKiqBU6dzQyV7lx3jb2XvmQVJQ6pmuL4tsiJdcn7+nNZr370RNjeCp4r+ta9W4BnG1Iq
j7f8O7WNYKambn69Iag48ZitTYSOrF0wWMpzTl4sseuG+JrW6sOCCXlj40kCKnAsS+qPwymxJApC
KEIkUF3q7WRWwVqcR3o0YcB993GqrAJ1eCmj4OGhQ1NEufcZdoh6nYZPviF0AptF4PPrP8XpmJP6
3zteMr4fSk6vDV70MQUJ45BdChHZ7XJQjDoWRoTpzcwcSk2qQQkgStGyeqmN22BYfXcl2jUXhJh6
7w0QEzqbd+CnlfSLng26geC/iZ34Eo8D4/o+CrdFkp4bR9CGY24dmgQIh7FEHE/mMLhjNfKm0U1a
mma7bJD0oZ79IfAcT1s3DqV9AafQ980HG3+VJkYU8WTSrEmbyg5JuAjjdEqmFh+OjzFsSle/W9HD
aXtzkiMXHzxc7a4D6O77OxGjR3/qUV0NOX3kGLb20IAaqRQ9yHL/S5QEjO3RNGC1AHS25jAVJD1E
BaRXjLUclVZP1YmpBcL5GTjBg/t3LzIwXvX5bJ10ij587UUrxjtlJ9F5VBVeplaJNBW58EoszO1i
ZTYPjcZqEuA/UXJuP1W8mZRJ5vYbUmKcsg7zb/RAsAxy8EAqM/+jBZlzytWQuCm8Cv+gn/yJlJp1
23ZHbz834YhD0I6ADERVGQxW7UnAkwVYClzZw/QvuGfcwo3ITXApfTRsC5BgQn7EzCFNhJRxkUtc
PtP5yxtrjoIYcdk67qiXorSg6cVaTuOhYCdC6AFHbVJlT6cmAHhkQpiXIm2dzZyOtolaTUk5XDuv
bSyzwgC18haBqPrgmNBcN+n8bsFyXgU3AIUEwrQjpuHA4BxrpaUslyzZ/441XV/WXLo8vP292Rfh
2Bbl2kkEIpYZRV1lecdszXi9Z9fx9HiHEW8o5KpHu8nDWDV88KECAK+T9w4T+10DCnQkcWJjwhTh
4iYk9FBEw5VPSW3cHjTg9qtM64UTL/0Ux9lhVl3KQsLWSnSLP6uAYhWQivANDBSJS3Jep6CDUOzj
P6oyoWKlFsV4iwReQRdCwPfMak2q1hTZof0P7B5p5XHtLPs3X5RHl/Wg8ERg6wu9ZHPG8C5P0Rbd
vPjpQsRswBHOudn/sA0Jp0gtu8pJeVnVM8qBi4MbG3rkWlop1dB57bmuSFEBSrI4XUp/FOnqu6sC
AOzmII2OSBJc+uG5MpyaCgkZ5Sy1Vmh0+rn3SxHoLVZ3z7M4MyX8cxfXUMCgCXeJ/658UxCDK/Az
WEW3afxT2aFMhYfx6tISWPUUIOdlGp5wQAGZf3rJ18DagVpz4x77o9J8u6cqDw6OqoZV8l0T1blF
rrcYRJjaW4bJmyY9P3npaKTF+eO3UvvR224xhkkpwJ0/AkSwwVd5FIpYvm0t6vYCsXrJx5p0mAGg
Pb6Rq3sEauy9HMguk/4c5ZkScFKOmyQFjUS5fagda+I97ZjJqoHcKHuHR2OzrCWHaikqUVLCLhDa
arWKwKAZFUhL23+ZC8YmsnXunmVB16bSxuriUHYdnrIrZ0RFZddbwZ8mhD39vULXlA3a6eHF0yZh
KZMXO52/AiRi7ZRZ+ry2LbongsxbBrTrXZKVdrmOh0M+b0QjkT5NcgVa3GNO6vfJoHO8mhO0RON5
LMxFcz4vIRMm13Xi5KjjH5LCuuk2Ifq6S8ORxkOnKBf5WKCYsEVczJAAdWJJJmZzbx+cJP0zMT08
WmXgSBJUJGgrnQkM3rBNkq+QA8AmEUdIeZDi7lVz3Bnzg3iSVa3ekkvKi9sPmKB7hOttjdGZgiI2
YLoN4whnVv5kG7VXb8MLvjwxr0jiHPEli2cWx/QgUCpv3xg2bRvoFCq6VzMOpNIYaq394H5DA3pA
r0Sdk0TVgo2R0z0D9KQ3EU0nUyL7psDXbm/qR0oYFaDm6VDvtMV9sO5GFzBLVtya+onwANq27VLg
1PagQzJ5tNhVHKWgdRWz9ucVdpki0KlPKxHSLRVIZNpFJsNeAI8Zy3aMwkYRGiH/M9DxB/zU65e0
jPMHI5c4474M6jeThPkbz9lnQwEwGevR8Srn+ttnRX3328FPT8NUT0X2h79xioSW2szFlcKrt292
s9XjWt4DjLGFMkayMsWbUTAPkxJiZ2tu34NEqbScyHw7aa04NTP3Kb1bTddaA4WqNfzoLNU2NUJt
hWtZlPt9QGyPnGxjp6Xnv0zdGKezRwutGc1pV5w9PRLlbXbfB+tNajc8HFRj0AojqciCmu/CfraE
ILj5QGUlFjERVFae6N4vb1QKTupJxeoqQv11a8SIfEXsxMsiY78ZEAiVMnCjEDiXT8RGlXW62WQg
eKwhauQ4dJ77y+DfnFfjL3WUn/QkfKzUKYFh64wI2enNRaVzllwrADj6jYjxCax/AufTvLdlKBrO
n8doB+FR3fdQGSCgIFjO0M/2tpULQXnkLLHYMwoGt5yL3lyOPckZna651or6HAGHCo27YVUaTlzt
aa+vHa3ncaso4reJMw6qa1lge9Z/ECTzYWq1w2DRGuaVdiP+UFxWz4OcVVM++kxvmATTSvng9uVR
SKSVOOVoS5tNx5qaoCXkqmjECnSYszF5U8AMVs6Vg9otQEG1DNGpGJbtKxoDivOK3Q0paVjmJU1W
qih0YlrwE8FmruHsQDTLcYsh34jF5sbIP6DwqhVL+oJ4w59NxQJCd+2w0BMRT4L8U+6rUn6CN9L/
ox+s9tmPW8ivEaYqJuWclLgwQsnIvdvqxHZA8Jzu9IR66yGRpA/Wj/39KRt3NetFIm3Qvq2gbA8v
3A64iywfxlXbnSrs0ffzWOjcJ9Wq8bgPR4D7BT8abRFE9w9P6ZOuMQHvXjpraR70HCYggxfuQ9+o
Z2n/ngQSNHrarFcGdKNeOx2vfBCugX6luhqknY1aGnRSpoBxP5mYFdFS0iZdNUXA93LL+wIxjJ3p
dw3AwVHf9sim5DDO0lERDFKvFQWivTknCOKmuWokPuzpbEiDiqWPws+zb+kBC5lF71ysOR4nRa88
7FZQ8UUFeCKJCM/eso646eHopOgkYW3gPjHTkZYoA98EJLbpM6Qu15URJAcf4voWb6tOT8UUyQRt
doepZ3FVHk2RK217XFMIGaDR5hoJMYi3SMvANxDw78qjChWBp7u0ITMY6xQTbHJ33sEuSfg7Uj9s
JqXvIlv/rOnEYHAnBXEgxz2wzqgkgXsTXObfx6SQh5XLHuwc8xcQ1BCQu6zmXmcVsoC4obswbZ6P
YpEbcJNGLwWIp84gdViv/km98td9qe+Ka/q6RpcKt2UDqlgQGus5mJdoG8KI2/+svIUxTnFoIr0T
x1UOWM7S2K87tmkmw8qc0+3o3gHYqg0r7nCuctaFs+jGH9RYud+hlGFv2Llan1KeMt//xH/cEaGh
Il549nrSzTwOO4qp0l5QsWYzYrqWPmMs7XDCn/z6Fr1gLNkjRZlTLbLUwFCHm77G+7qW2mwS7K3A
HccsRTe0zkj3NNZQqXc5gSHytZGzieJv3GKXIxvBjuIXX0P5NPw8dT8XWgyUUjn9idjECBIvsA+B
ieReviNiC8BLfkSlMDCYOZm3Nj8SqWq0HXmWKmPorp2f5SQ/P25g8fOgw5A+VKWbUCs64KLhkvFA
L9r5eKPAjMqnRunqhI7vjr7jbPfvVHxmmK9MxFq5ll8AlOmrE11R/lQ77iMf9e2tfAiOSCEKDMbv
BPpCdBXhDsT1vjF4CRMF+Y/3x7nxb5kzx5sX6Hix9nJGZBVovkWTqBNS+4co/QyYgN7hRaVgwtmY
CLDlMkEiyY7hTfAk2mKh1CIf2fmRpfWnMthdX/kIyTLuqQqrZTIjhm+dsXHpGRiO9AHAS14CZAPF
UHbi+hM/hPSRE+5iQ4wiomhncrU9OzUf3r5sTAzPAMnNSnYunyiayLwLT1zLB7v/BnfS+sQdyTLw
/vVZJXU1i9Rvurvrad7BCqI9RtISdODRF7CMMCWiSiYccUaoGnDcrhOkrUlasNklm6WviLQAaN+e
u0mXMtCKCZ9uEV/9JCKqUeM/ZztSMq0wos/z1rSNQIG0rltT/LXrwdqmuKIsfzWLesH5wIR3Wj//
B/4ui37LzPmcT5JmGcsqV4/ZK6hPG31jK/9Qlr+76kFL3NjrnI1KbtnaxNyU4dOxxlSmA67p3Qsd
8j533vu3HN8KzSlbSVNRFyKLjJkb55+Y4qiQDzKicK+ANDGz9oLCLnImQg9F8CZxqWmgybeCg7lX
3GdT4QnbyUeh3QihvF851HKBleXVTn+8OkSiJObAiaxwDnSjvw2GL1Ozmp4Dyuhmy53/Dg31iTMm
dQiaTcd2JpqMoPgrrXUDZLJrBs7BaFeQ0KaPx7K+x04mvd0NuyMPbCKeVnvOyWFc4jGXbpNQwqDT
SFpgBwbPWMB/UQGuSs/df60z5v+P4R9PM4xO2gBpfWrv3X7VlQqH75l+ZIrHv3O8DZXamYFGzlnS
nb7au9IcFGShThblv8gSgUwWj2RBw4yg3pKs1ptMNpqz6VgHZZvgJd2UruhOi8MOIHCIBtVykEOI
Jw/Ggd3AfDbqFPLbIORRaVuFjNhxEsrG/1m2zxqY9jb037Ai5rb1w13BU4zic2v96v9i+H/0dfAC
wxXSfj5wG+2UTO8PqnDTHNlt4N/AREvre96GJsZ2Vbnkhv9bvAx4y8n4liI/LZKuRUG+EyvRm/x/
suz8bn6hen7raltb10k9jU+JyLWtI7Dfer5138WFwXZ5m8u+58NboCXziQMDLMOyHW5/TCh78K7I
j8SDsBY/zeixSVn2GubbaszzO/OBTVPeuH7MN0xm/3O6Na33Zf8zmiPZD2WAugHJzt7EzNAc2NKK
5ztVaKyvZdDbpvoGvr+UThFSG7gC+gDaoVXVk0NwRq+BGuGMiGHReiHREHntmHNIiTAjf4ZJ2LOR
+c2Y7s4kg97jFa6kroxW/ded6U9T2xfH0Ig6pLQzMBsDnJMoysx2SrE/l4nXCvxKH+3DxZ6i+/17
I640Uwf+eUy5JHeqBZcAf3g6ytCW8n+F6P4NNyAR9g2OWYiV3ib+4BP/XCgrce3Jm3gnQa18ZIXc
MU8hWNTtXUvt9a3HnxJArMy95dUU6sq4M5ipPJqWtlp1c4baToBVV8vtHN8/HLjGCTArDbFBTqmf
+ewZtOldD6O5s3d9gWy9q9uw3ZoLRFi2z7ov5iggCvO+bUAj9OGg2Pu+u317tBtGugFn/3orFsPB
VrGAxxjPXTKp2OS/RJg16BT0EnSnYptjRf5lykqQ5mw0qi6pGScjYZC7yaTlIgWBk1ssfIcPFr4Q
NrN4BwZDFtF2QgDz7L+rNa8qxdWpBjrVqG/K+EO3PH1hPlOzLeKCWv0no+AHaAx2Tukz21V5hO7I
71MStrnW+9dIqt4GanDY0+PanAG1/W4BKC5eODBuExYYhH2M+qWecUMlp/UGtNfSjJ4kL35GUFgt
Mc27ycBoCf1ppRTCeKqvnx5hT5KjjxGOz43N7EH23kaK2F/h5lR/zaMoe59nONsH6DXNVa5oL/e7
gJILjLdw2hCa3LHL7HpP9t+aOU/QYDdyVrujc1+zxkyn4mgDB8qt0DS6JcCywHhz5Ud2WekWSb9Q
DryiJhK9LSX7cUl2GhcSokolFG5oGuhqUHXjqg3cA8m8h+wY8kCOtuHWIuKh8Fk0QVNaDqNZHPEN
bhPXChHi3ooVtNL/bKLotvAKmB/edaDPEAQKRXn+YV1punfyIp2tBAJs3lAMccrZ/IKZEcJ2QhPt
N5w22jpH/tahnDTkO3rvkT0AupeJs0ZOseKK6b3sQlfF57Xb5ckFeVn/vWq9q9dAGdqymrNlTxne
JrMVHkG9hOKMBR433IoweZKSC3/mchcGbknF3n0aQ0qrRRRPvJVXBsHjF9hDY5CSVJPN8ljCN4UX
MIaGupODSHNrlLGCPo0xord1a18wFZUkC3EoU17Rr0ZWOOLYGTbTWEviEu2SwVSo4DpJgA/M/wqO
z23Lvc4394u6xeobIa6I6YqNTDJmQJbYxDYL3wNz6c8JE9+kplpmTTRPpw9oXoEnMr/PyJaXbLcR
8F91lqKk7silcYW8Zf8z3+LXujJC1Q6bfHWusE8XQlGvT70ltQrLPtsKozakeDl4eGAcqN97XYuP
BxzW2mti9p2pt3oBQPLazsvfDFWDqAMNpzH5a+CmyBRYoO/jLs6Ra14UhvD7Dc/dgZ8NXjGzkXOx
A4juvtQOFikTTXMd4PRTFngv6CTZ/qJcZZ+bfVhSbBbPfEj29pasShzw4iQ6bK/ZOkBfYH3JwF4e
tUc0lfPx3+57Yfhio/03LUPcq9Pi6eCEC9/YcQWcKGBS4YCNgytbeu2acLmdX4IU44QyedvmWj4Q
LLU15BPV/izjwp/mD8RiKMWJjGe+hY1RaA/RUi8ZJ2tvws1VhHNfZ5Ck8jGGDmNqqTuduFBV7+iC
gcHjPESBiFdI9aQAeAignIjKZt1qqUFVSjR7d0Go/ErQm42dIIakIH3EhgK26ijQR8hvy8Zqmdzx
9J6HnyWFKXM6+kH1OGhc6nGwk151Y4uoanaSJloK1GBwaTJziyB+Nk0a1DqxTxri1J8QzbT39HZG
Bg7fRk0K3BCE9U+pDGVSMa7b5DQJElfmy+o3v0ZO7tnCRmMUAZHVIyEoL0nizPBM3ZgBZrtf61EB
RCAhxW7BdNouRFfiRS2/ip0gYgL4QSZncWK9VNoldsSMb8xF0hiYEuN90lezmO4PD1bI0P32TkPc
hbkwlT442afdzRqydJiXycT/EvSa4KolUrCXmTHTe3nr4tjMvyl+NCfVxrjMjlrUaDMVhklEw3JW
X6Af9p/Q/HqkiGsnYp0QRP5xmcTPozID2ClqJdlOEsk+ax7+v43HQT2n+devEkiAH0/WdpyQYlw6
D2dO5rz4kMUyM0N1FGFN3fk/Cmo3bqe5otMxpbdVJOMmWRmPY3F//7jAaAMQBUFqE3ubec+T2f95
5I1RSUsA6KtIJFbZXz3F/to+/GOhvaHT51eJOYRxGlgmJbI6b07QJbBJAw+N24OpGv46R0Q8MFAA
fnnh87lM9lSv+133dOZOwOiyK7wuiFdYv7u7fYTDRSHOJG+LnLgT1Qokam63n/Xzdyh0Ae+AlGMA
DSjBz0OFdQ3NcvjWWp+1H5WBeT+sZ52b2OM0nJxu91Hr3OJPGjprTmrpvkQRacB3Fo0YFQoCzzfZ
J7RobKw9yLfI1B8jKa0kCCoFA1UX1yYz0foDugIeBIRcdufy0RSmBQIBEYwCp+6W8ZCRVCthw8bn
UqRN4YuIlWIQj7SBNzD81CLboxV7kfEy3B8P1VX3wlTFwhbjAn7wbZQAMoQkLN9h6mXBipbKUn9J
WBR+y5wl8b2ADCfzK2UpVEh348SMFD0sylFYiCvOz7vCGxZz/xBB6bYiKpTP9DqQa2QHOC6ixxJq
doFbx1QiV1dggU8o/uxfvzW3hgvzlOYXsi4qyfHqEGS7sW7ZbL8feVu1VxC14MnTuuU76NdFDQ29
5y2F2QyNykcUhVvlnFsydsFIrBSwoF1oxgDnjYGZnppF5fu+njRRS/zU76gwh8Xi7/GjFU8soz0/
je/S1oWnf733bKkB2A03UHjSWUbwFV/DYQkxbX3vrApF8XV4G0jlW50hhpaNvdBfQRR0rJRukcPP
ZZelGnU1VsofBUQi0WOxJW8GAZgVeTiIRgyWN8yxVQAGipsjBynV+UGhFsQEefj4Qw//aOykSuGa
L9bRbulDWC96OeOZ7vBgwCABxvQgoNHVZKG9LHOlVIUde1UolPSOm33sGIxEi5ZIjyHy0yABK+Ge
AZtoBfl9SeE+0ldfgaZMpJclSN0kd54I1YJ8EqzF/oDuECk7rE1ZGko8eDV0X8u7E6AY9G4KZVBb
BqfK/8fQAKqS6SmgH+5/v4tyZ/LTdUYrLWjhKAxPh8w5rhiWd6y4gem6dI5YDxI+6OaLvLGp86mY
d58fcOgaMJNBBPiKkITFnz30v6qQc6pOQWtyKygSlJrvFWQHSlWUeGcgYDPqPViV0WU3aNXj6yp5
xVxdKmvBRmthDTmLIYdd+mjzhV3LqEHjKxdJok4axALLhe6HGEEx7qtmNROfAAhF5qR2wj9bXj9R
2+OmQpG521Ulmly4rqRqC/IuOvtZqhTpZWSBlS1eUIPw/qJF/ey6ZCpYhhETwGxx0JDV+ttoR8MX
QCTMEWlT2KG0h/G3QcSuBl3KS3rxaVS3fJ09vDmGmNmXPrcKPMgGPSoVO5V4IxuKUhdBw1Q8pS49
Vh2og9HvDZOjGcWvIaiTex7IoXdMoY4BXiWtZ6szJIxJclyDgY72fQG9fyp4TpVl7aUH8tcGygN+
dhi5jlKzfUw7U7tlyvfh/fDBaXF02wDaET+oOpyXJNz2Jk3AuKZIds5jkSyrbjx0/jPnU80vQM+t
rngQzE7WTny56/ZdRThhkvPAV3zXgjXjAk8xMJU7YXkJ2UQA3Ej5TFPG8Pnr4tQokEBc2ORM3FqM
dhL4k9nB7UZoFoIhXZiejj+olOhF5EGvCFhBBJ9En6Vmsh9Y/84EdIGVou/hdpFghtkUe6bxCsOU
dSWHNrT9mGxZuGveyhy1S/7xqri1m9KwbNCsGWUzHmjpgzp+U1orgLUxvBgj8grJonaTalZlTLW7
kHhY0SgCmhGLIxkpnlC1eBZ23HjFNUKtQWpPEIXeYEZZCTSIjMc2gPNssOmjcAc/1YpPQSVI5VIc
ka7ExD+IUruuRIVFT0WJpYSDE7+L1aJX+gu/vutdY7L81Z9XTWTp+HnWt4A5Y5sxJA+k+p1X+jen
s00+SbsLxoRhpdYToH/+tsJz0andHfwoiM4a7/FbbByPT8Gsr6cUpOQHASJo+EWzxa0gBFyinMo2
CMDwH2o6NssNbpOLBLfm5A4gRnwQHk/3L+dCwEww8p9uCCcKVj/DrNVaDGyAPprSZx0SEzUEuhGV
RG1dDDPg+Cqd9wfomM7W8DLK7xyShlKNqIlZeuJVyn6pOMfGRwfAedj9e9qGcx02G8CXSQKbpDwL
zmzupDMFbYyqTSdjjZXZwX76uV5tYte8guqm1wTOGuZY10oThE4/4EPjMa6aFNAVGAwQGPwCwtrl
BC2C+GU9CpmHglcWOa47bavegZVe7CmKz3EYFx5zCuDVzRNS1ZZnzP26UD72SwjeqiUkMOafxPcG
enWKdOTZ3btmL7ABKtXs/XYakNPLdigjhfvbrkm1YjIaTp2oxjuOqUXaYRKkp9wA9QY4InmsT/sz
IrAHuJIH6bcCduHe5ZAgn3MTGi3uIU8zx9fj3IuDRz0/RJcrew4NdaZv9GFC68xEtFHqvBbSwohM
4QlaYVDm3P1z8nvftEF6oa8Hs5UCV5U/87rZ9njY8UhOPJnGHYCcxGxL4Idd3PwdMc4eMK84GhJa
D6WrF3KEmo66GitB/EerNqvSnPF35/hZpvfSCVn/07LmBJ8MuYOpfiXasurjhBtUMjPmP+3mQ/Sy
ZxTQTfTuRuLMsvD6HPBQoUm3mGuvR7mrMLTgUF8Kx74VT9HoWjOAWKk35Gx9cn3dVndLFojVsGyR
iMwC1Zy9yFhnG0He/aelqxysPf3Pk0PQ5j/mTe+eJG5Kwb6iiMPgR+RwJe5CXoIbxaN3qANOaXLT
oCVtYwF2FxlXL8s3tG7M7jOjjKnhAyov/u+pS5KUyqOGA3LKeORBSFUlV5JXlnt3tHFefRxdwgZ6
BLizsTcxbLBZluB4sYoYREA6xS7iX3N1jCLShPRDr4E4nhabMX0/QYMKpKiVu6gpKx0mMLysHGWx
q2XoA6dO1lvcZF3zL5RiJnC2qorMVZfzqcVaZ88/jrZA5hf2q2SXHNX6r+4LksVwsV1XTSPehLf9
aTrXm8tzyHbc4OEZDzcgvug+OB7uIlhW7LpGYEvqjZeBQmOD1/BoviZklZjfWnVIURlEtkVGUUSG
36JkJg7OV+iuTDW52Zdb4GsE9Us34dNfN3ssDwOEfNdcTMUqAWU5Mbd0sjgtxHJgFy3UDOmws8jv
f/ozKeCMmnTXECwIL3ZfHz7q626D7zhlQcVr2S0G8r6ndvmatOFq1ifSk2lcG/mqDdKZpjKeQcZS
pDfO+4x0Nqa9s+UNsEDrhZxhRuakI5hjIDIBaCfoTuRVJwYRJWX147l6TqK54zx8Z2XUyfji5b0c
MSHP1GSNgWEdd8aNJuGoZsIvbMv7UvE0md2Ygfomcq069cv3KjHUuh1u8wgnCfVm1hvpMiA+RSGn
8+/6ZTJ0+3+2F3HLnRndcebvl2EXzOoYnZw3wEPPlRcLtzimts2TYRdcQVpDxOMn1GarDD/xOdEa
EoXlvaVI0pyjQozd0A6QCMUEEroKS0Dq8tqs7ZQxgb7g/bkzWA8klNIxC0p5ECSW1jc3KZbq6lUW
FXBBt0rXlYZBtxog7dH95zTFgjRifcHw0geb6WV13N16oW1H+u6lCWJ2wN7NKo/6ERzi8/rip/ON
lHr0R8r8i30e8Rj4ZYDPaCK3j40GYHlgIjHnclTydgtuDUNwZu0AYY+GsNiZYj00FKr9Y4T+jNCM
/d1QioQRoCfYMUoWFJXMm11Ooci2ru7icr3ffwO9dwx2LJ3bb6qcPUOS0f/GPRkfTCGHV7RhtqWh
1l04jWoeN/3T6yEIIrRQleGiYvl5Bw01c9aErNhXfq5ld8pAX99n6wbCScXa8GDesDcZKiOCSO3X
Fx0HrErywDp+kkx12UfhQ473WWsr2FlPts49DgoAskS3c2gSJ7kCQTcnFPv53eZPnkJkpvEOVJJS
S3klADYIkJWIin6NzjYVAxrJkR6Nt+GZbzZpl5/EeOTgD/8jrWmwiwtwWZWYhf8J92u0h84KiSQN
BiMDyEHRFA5VD20Rj9EzC/usctN4FA0gRfGGq7JP5KUmw0L9HuTQyd3tBb9KDCz1O04/PCoVKUB2
96ROlPKrQtO/f1ZgRPUhDU83hRF+NW4vLVfvYR/II+95tnwYN87xAfYFa7+Rdne2fG+gFB4hLIZM
zxYeiqmC9ixBKmWoC5xa3wFdii5FbSj0UWC+qMlI5tor05eOohm/X/defHcnXVB3FfxkBTf2oaa3
PVv4jLkE9JpD1BshUkp50TDCzrT41C6w7yMuXeh1jnymvMkAPEPlQj/DE2/tV1+db9Dw6QY12Sj7
ZfRidt73/onX1Q+nU9tV5FVtTJsu5K6rosm2Z4i3OQ8UkfPir8UEpAvxSUvh7lUT++MQo+XmDUyX
axYE0bIHaB+dsx7otO4Dh4O/zHrSJVgApcrKxGa/CyUznf1HvhmUnzvi8D9ft+jtB009F15/kNFY
JiJZumv22/x5PCbU9PZsO334gHzI2n7rzSJu2A+eYHKiDhJv0F4BoSC/zX/81Z6BOr1tXY8E1H8N
kkMXyEXPM47w9deE8BaSPKEzMIiS9ZGRaCPRGdXLAWITZRofRkzlCVJZ0CXl/W4/4zjkWqfp7a9D
+393CUm/3nj8i7FdGrj5cHHzB9XsYCKNBL1NhdCUBDkRtiu4ySvZsK5+7cDyqmGiHh/xcnIlihQe
FLsNiopsQf7cezLpWctMj1ZYe1xsbeu0iQQYG70/jlSdNPhNSKJkvbrldqHBtgSvBwpB6ow9G9MO
vg6Pev5myHHHtKYZPHWH29BrTqpxpnNxDDwVc5nyFAuzt9Nrj8OmKgbIvvppi+wdbJb6SJgjC4U1
GRw2CEhayQBQytCpQofFJ89XnaEyHsiIuWdtPeIK7OVXlOZKj50lTOnDmFuc1ABR9kOjd9EvAbXQ
UShXfPdYrBrMSSmwenTOpZ0ATHKNF2Oh/e4uCfqe+s7pkeiYp6A1TXjjtAdBFpskKIZvRrocd5yN
R+9A1nKEzJtNhdLDdztLXW14TZq+NpMbV91dlsauUUjo4Qh93Dm3SSuxEA/newsFZYE1LemKTjII
eNce1lWwPzTxVM60PO5Da+d7/aovm+7X6m8D5o8KKW2W42yBLxo0+l+sJdgcaQsCave/GvHXPp32
mgeeYiu04e9LjmdKVFG3SUiouflQRcg2yeF4IhzZPxFrmTEaj768jgWf6FZe0UJ8phdqtnFDp/ac
AY9rerCKjz7kpFzHkNPH6OmiKNDCRWKZK4iIz217wdSJSbzkPG0fX13N+T5hzFbbIGkmcvi2ADg3
C7vEuwdaKt4oJgd/k6FBvH/IafaFlQRaDvrqzzuyNBtg2htEjNg4TsGUKlq/xPhAq5aFlelrUbeW
oL7AdxaqFJMvG68Ohl4oGdZq6xj9rj2bgH97lk93PSgZwb8b11yF5mHFJki3TQBCT3P0sD3XRV3w
ZRMQWhGqC4BMeBuiRdckGzBMEPTQLrzASe2aAxiD6U1YVje9FYBE0jSQJvonYvQ9lFTDEqxJRjO2
f+XxMqov0l5ZongGr/o3jG3gnBldQ4fZ9CiRZuMGmjG3fr1Ip8/jRBzk9RUYKX5MeFqRmIaToCUM
4lLLBikdS4LDBTlSMoFahWAVl8CxfQ6KwTBY4kqHJeghTtwIzTAc1I3VAlwd17hp61HcC2D/nzUD
6fyHGU0Hy6pAUqMQ9b6IzIiBXAT1nqaMi2d4cacNoxbWcARWZXm1mR8dsqIR4qxwPYe8I0jiYaDL
WOkhEi7gdTHLiO8rYITXfl75Ijs9Nrg81akBHzexgZDX+K420Poo1JYkrO65dun/p+GxGaBYEI6v
+kz3cofr6tLcn9cW92Nqz+wTpSu8QXtyM1r4IwstagiYa6km2R1bFIAn0EJBGrcR20LaZjG5mhR2
+FziCm3P3d0xBVmxLNQXKDYRJn8X/GYYg6Pwu2UKwsmQ7/UgJxaxHjRwKZANzfZzdl310HgHvWbM
p5vhNpXkmOBefHi1oSLbnk9nYp6ChMWcqKGkrkWk+xOApCPInMfpgrWasTFZTOGlTfTKAdC6Mdpv
PArJB49lnFlmh2vQYWHQG4v9tPznDl35bPdhvYk7xaHP/yXQE6qmkq+072BCwKaNpxdSjcnQwAwT
eNU5BqLmgpwJwls88JXpGB1iGFnvh8wjxA9t6zkllleRQUIcQ/nS6uXm3JymiJF9qQYhihqJmNFq
o5NYuv8ObWeFYSFftBdEfxUjC5VmHWZ5jHso9MMBv6Yl28ebuXrYIznG2ZtQDbUGQpQNNl7mwPU3
b9qXsqSSI6AC/74j5rZjynsQ5LAGsMOCiSAv80CsNrdEEZeDMfqhxOrcY9EBI64X7u4RBvQzqZd3
7pvfpV+q/nA7Zc+y6fKzQmNqqUGafS9y898M1Os2hYKNKcvDOvtG3iBjNGZVN+1rctJE8Ek19J0a
u4acXORh0RbQumSDANoJq+wCwQUvIjBQ0MSqM53IP0D7pUMXzqw9wQ3zxhaRNVMH/kRF6BUTEGma
RSrwFUT0igthL5mLIUIMWNa3gsfVhgtl0CaOsaybe/CCMhnO/W/4bt91BzaYECzpj8DU9TOKuRca
Ci/wVX0tSieb4/KEhYeYHLxEEBw1cshfDxYCeOQNGoEQ5hdfCb4hj4ysPFT6o84mr3ZKTOlo41Gu
hLmWDvf+5vSL/9q6Gi5ifi8SHSQ60HK1BXoLmRlWy4zDkxCrNtVljQbyB1NFQIVj/vQ1rNsBbngn
b0jYgIUsb80IyeAfIsh2dCRDC49/c4WTNXEi68xRW5BxiA23JfidCCPSmHBv75qodZTGhr+B1mXi
s6qQzg+WINzRDglLt+UkOka+TEGetXOumelJsY2t1sXew/4NNrahWlo5rWGnXPcohtIBgICpM1C9
jVib3vcWiVaeMZn7WxnLXWhE8xOgHLZPSMLlXZfMDdPIEZTID0/xB4GMdeYvrEk/iNqAhXqHp0So
qZfVjX0V2dWO59ddyrZAZY60XJKiMM+5EZCago5qDtyn8wBO2Y4z0Kk2QLPb1k/cF0UbL+BX4sc/
7yKOLYG1KxyU6XmGqqBQzYL5YyL9u4iPwf5cLVnaDulByTESrsvZAxQYgeKxE/6dmMQPi41aSeJj
FXt9VASglMKF9ytkRQL46VBH9PAfmjEqAMyteugCVGp1VsHucYHNq3d3aqKRMdGavQbtv/QWC5ze
SU5O3QdGZly3QEjDJtN2Kt/j7ZEyjE0ROFL7rArd3PBmmkshAhr1xk/tdDbhrUg2wNyjoFbHnE1V
pmi1B9563nI5syfFxEt1cayRp9hNYM6+gLJOmZYvAfM22+bXZR4swcu6DWigSntiEv2ZBu28boJL
t2FpQY+sBfqHn+FEbpEb9vEYhuVokyNRiTABJjcKamwjuP9r3kxBEGBlK/DjwOAYQr3p73RfmRah
H066PHNyVWj/aa+zaWhI6QAIreFhGOJbNAJMWgxPmdTL8CC4l8vEF78a/tsTJ6UFxBrmZIKnvaMc
WKX0SZYPw/5shYUOz2tsoJE4nJIHSThsIXA1L6FAFHPmgkYfKyG3sSJrq5TeaNzSYUrzONKSs2VX
+lNpYsXpUEd2ppXmXb+1Wce1+Io2pZs4sG40TBSalSGyu4VzHS2gVx4qWzq1/FPvQNRScBteW1xY
0/G9Azk6hO73QEtA+EtGwSTUfA0IpMDybuWdsOVWzvrETEqV9HDtq9yrX8AOWABNjsD3zz/mx6R6
lqL245Ow2PVhrTKPr+WSnIMbof87cRXwSUOh+YFclKqESrU4MZEx2mJRD6gXaSNg4WZqqkpu2ybd
rUUOca9pazdbMQSMHVBUamKpPxqBuEumMWNz+UfyTvF6EQTF9HxgVxZcllzMRwf6yv09yb4gHox5
kM7xAx0SPqfGn0YxxM3WYowMWcclzJTIKn5MnScf6byS0/nblKJQ0b+f1dWJc8JwPsyqmBEzYZg0
gEZERKQy8NGEpQVOxjHXx9444Djfmelh9yrFtgvwCU/xLBCRoYKWejl88HICOhbEXthnLnsIXZcM
rCT239g+ATi5vZVaFXQYCQc70DbuVd5IhyNFKTBXgs8TdJ2OQLsziJ3kODG5HmM13zOnZPxVxtEJ
V19mlIhJvi8j/a3OZBt5tz7z20kBXdJuevdSLzcd5LmIgJJ66ix9indfcizbsAjqhQjZpaFsnOJV
AiTs2ew3ZHPYPsPAU/O9ZYSSKXE2td6vv//XSZHAOm9HzaUpSAqPqd8EiEbB676v9ZxtZqczfOXZ
/taGSQUsFG++AS8UvWoNOQhOTinEw6FatOPU66SvLoJ9FnG1Wz53IRydD3B9WfIuFAB9dNGAf23d
MwWqh98lER7DvzS1RK2Ila++ILB6q9kVvfbDVtK2nBzcZ6gVq6g7jO3acIAq62nZzYx31TJgQkGV
7mef/H7HuvgYW0jpDlgib8drP/N793uOxE+hOh/Fak0jVRsGBFABTQ2Ktf1r3iUIypCX3nPKk49B
DZRXvjw6NL30GvYlxgQJZlJc0GUKAIrI6lzNB39fZK+U790prbH1+eoy2heAT28n9LFezyHwWliw
U4FlKUGXVFx9j1txFuEANK/Jxz5i9qsNiiJdWKxRR8YlvhDCPsRslrPBEZI8ZRjADScoPoVABXRF
EBDrZqTZjSK5jVJNPcSN3MvYLc496+pnJFfeixl/mPA3z7M0tcx7ZdSlpriLgTuCFtelYro3hIIH
c7xCxj5k1Hwla1FCQCSIik0t4rVk6tjLfO9vm4bqNGem1fpefpZ5PLSbAtgsWcpIIDOxoy/3Lx01
J6CptC1Epf90H6EvjoNM9EOFHKIkH+YwC7z3caoUmMEWR0x9p6wPIIvk34cVqfFS/XIxhIwlvcbv
THVdq72rEYfoL3bPZGAO9DvxQVx6sHddOPYIXQoT9qUPyVI3OeG+P1Fm70YFkiPecT+vE3OVh5ys
031di4u2YCt7we6Hau+zs817acvzRWtIiGY1B8nqxPkTuSulPpb1l74ayD+LF1fWRLd1sjrazmM5
2czGIqXjcJa5AAuSI6g1eTBxcFC6JdCTqVaV3PjhitVi1BebqfkknwRmvpIzgP9uIFAWg0BxGDRJ
DRmJyiSVqUwdeuGOXgdqqDE0VE28+XMZHHHq80NSJcPt63r1DmmDDv789AmcXKYFAwSwsWVG4O+X
gMzdz7m68DbuLpsc3nOTAlt1tGwV2zoipdAWNZCoY5J+wHtZ/7s00RGkmH0E0HXb5Vs3TaQzypoW
gELM3X1lpwTpi/FZ/ktwV3mucSFC1UcXWBoJI7AI6TSuBHxPDqOv+MYO48ZyEFNXU/MCIPAq0c/q
v0B3Loc4eTeAL/3BIESR0OIGi+9lG6XWWDAivjdIqSSd8mKPtiI1O+PV8waz9kia0nejQrNCDVLo
XVWeNMdwKnhldKWhDYoZy9aiXIMxnL0Ab457OEXXHXITAvm+EkWfHst0Qr3y9ubqIE/B7M4qCt4v
c/PDtVeVgka+TfgA5UYnD3AzDWds8RC6ZHXvMIID6+L8G/7idswPiczYWQxQPunc9TZl7QkjpJb3
yVOskyzY7YoXk7djI67saJSk8q4sSPxpUoFXOJvXNQuH3Xly0w91ZCW9+3OzFcecybmcObbzE5Ea
yQNJwJqzoPlQeJYN6f+14ZSPjGBiELYB7F4bQ0TgLPhnMfhhjxSZ5iDzVOQG3ZrplZJ8o9f0fMJA
hYUJGPfLhIiGWXmMW6lDJhoH+FBTrpOHw4AWJRpxze/1zNMAMHE0tFXRV0rQQCw5QhnY0YSXk8B0
Br5p0t5nMlO33qdjLUWJVAd9Gc+CCsDwZWxYRQk0WIZbs4VejEu+FjOoUNaSRqGeSHX9QWKKpvd5
U+iO6YUQI67WfHZHJBwlJWmiJ8UI0saIm7JSIfrp3GS2p53WJb8nit64McQMiMCvLKwsiP+zN8s3
0fsKzlnelAhUGvVbRFS9hC/TY1/n3a0PuPMxnxwvTsuuBtFf5I0bCKszII/Xq94GOzgPlVbj1ZvH
55uEgydj+aOrMBWI37tc4NdouRSNVbHsxZrZ0A/0h2aInUg6br6rJ9uJOW92xE3vMuadgAxdWqxk
j9P7639Vcz9fHVufjRoeilDFHNfrIIpH/FcL5yd3yQ8nNBtBR5S0RwfYNH6FbT2GN0kBHPqDCrDp
avCMdE8F8HEyqVaQp66g6/zFFSFMa/9W4VfofnT7AeghNPBtDhReGYUY3e20T3w0EJqTqjfrVquw
UIz7+IRetLtM1lXI/OwmyNMIhU15GwxiK/GO0Yx75jMRIkgE09M/hSBLCjsKNlPPkzOAqAdvoRLL
4IRyaEdXTo7HBRWO9TaAhoYxYbmiHH4kFI+1LD0HHjOgK4PDAXmqDBiN+lnzQQsxSmJpXS6ZuPxq
g34LxWRnSbT6jyjHEOVQn0227wqBByTh8LQNbYCGiTPnYszA2DOKs6dpx2pSr136jbBnKCOx7P2b
J0ZrYLNzB7Ptn6lzWrxCMKYEvfqhKmrZidiRFDt+HaAfj4nan3azMIfyd+zLgBuW6k6J2TNWhHdQ
iUtVZwa8EA/TXDIe4AsgqlFkRb4/EvGRlsDq50JJEgGhrA312cTixWPntHPk2pqPGB6neN8aIj9E
UcVx2A6IBk9Sq6Se8nsRHl6qvT/P+8CvUn2xYOnpMUYjK0bYR5RyRhM8ECePn2sqwC2YbjYX9bTp
0leaS6DBO7DDdMRSl09tdl9Slzx+Sek1+bI/+Y/jMoTQQzPAj1xUpCP1biaWa3vuLi0t8AvtE9ed
zEwpAQ5m9HlM7hsHPnABaAoEMFdnoBN68HXFCieyAxus8UNpUuvOrdcdhJUDJ056YRQSKPoadYfB
xwx46R+KP4ZOhYk8uEwjW/0ZnGUE2mRjpd2NrR5gdAGHE6Kh/4Erzxd/nxfGfslJLeaPn66Iizyw
cB+10KOsG3JMuTrp4m+jlNzu3MAZXaUIiCHapT2XxkVj4f7HnLyfhjvNv/2rCC7tyq4isM5ZQ5l+
lJTVLf4Nl74HEb9ePBqOtUCOAx6s3KPSfwyb+vRoNsphyhNuXwpvGIBd1dbmQKraj/Y1WZqAeoqh
8/jGqntxZYgTBz/oOt6ryQUJvJjKJowXqPxOUWOmAcj5XEOp5FNBHNEbRC7o9zk6SFqSnMNzP7Vg
/IYaQn24V2IBZtb3OPETpKukI+F8rRBpGERRGXnw2KnqLhMcBQzuZxzq80ql2HFLmNrKWTbI/G59
tusvEpy+QgueV0qHS9Mskr5IsxHLu9cZ4amxG35qK+FCfOPhfTHYprVDO40uVE7rJQd7H1UOxDz0
YXv+uLctxBKAEpYL+XyRJC0VdJArR7BBXy60jce1fPdBZouXxzvaTLVvvLi4MY3/XS3TwFv0LCnK
H628tilpvlzT9QRmy4K8BmseYjdXdfHssTwjAYvxVKqTvhBH2eittAoqKFUQY07tonYHFEfpqi8s
S3Hmm4EpaKczZ0MBR+L6DQ1/dMDG9O7dYXOwhLEbkBRCuZPDgSoM9nPKL5uVi8NegJSgaMfonTEu
no6HfJlSqbF6d9PT6hpsqOUcO+0MpTG1NJRM9mlAk8kcNqfEQh6B7jWZ32l70nx0+Nv0r6brJBlC
3F/1joWYz5wxC/ggSM1SIv/WWnpAL2gw4LvrXPSl9GZa2tsprnmVXkmn2uELYA9NXOjrfJyF1Gnm
6gNFnpnNu5lF3ctb67QpCYCavFei1xSobgMch8Um451iVkNbLDE/FgD9w3/mCmmtcO5MatstczWG
TiSS3M4RonHAvyJAPhHSzA799ClkhffPT/1MOkpltBULsVxY5aRb2NAyGB3+NizxDEoJgYNYjwyc
x+5/VonKrA4D0FImseRRbvjdN7kR429n0C8iYg/kM8lG0z68jBGWX4OyP32PNsM9/C4a4SD7yPWp
9qxEstpcaWqLP7+UcTPlZ0AdDCQTwGzMDTqyQZ7J2Jbm4cKZSUZ/cAR/I5aJR7rGjdgexyq8PGnX
JCwRNzbOLArvQDvQictyAdFElE1HCfyprPDyghf/I4jc+MolZfyPUGjTWHpJrAHVwUjSyWWHPt1I
vENmhw7U+aSDKpqzSWm4PeeOM5kPclwC6Cv+UNdvJfVdF1Qe0QDO8VL/8Y4ccNMHh6ho+vXQk1Ei
slQ3iZ3dKXfh8FJtpQcqzYRd50wEsndK612rpnxr4LY5iP+qAYc8uvrq9NSzHrNTvvp4Q3ryaPQe
xoYh15Nriih6K6v13lAGlwt6HA91lL44x3YtrwWQUf4hzApSaWbwMWx1jrOERtQW+ZMmvj6f4gui
hrkrLALMxQAfiwy+IhZmldt8myX/n6ej7ctup1kKS7nGdXAYMlbYxSUwzAlgKByw40k7CLAJA0Mv
1TazZSILInH9P5hAdkq8cF8YxsJREbTPBSjkE2fjX5d4glftlE6rSzY8w4fmOD72iyeShqfzo+6k
z6K2L0vyQgy3y6u770wnYu0lyJxgbFT+LafYOIea4SZPwCM8Czd3rwt9NVrnFZU30Y1MCWzFeqiD
zZUccc+dHQi8m/wRhP8f8JWkk073gAwU7lGt3hfAblmW7KKCO46pFBqo3gLFpc/rCkIQvZBZSmKk
nJ34t9LKxT6V692iXuL/p1SSefVKLUzmheLzqVyCm3OfeVWwIPdkqK69NngZqz0LH1BRg2xAntIf
SQMM+ruc+120RQ9h/9plewIgkQYB9A2mp+2lnlYUqXIqtOu5uyJj50AAz4albMZnmBPpyT1Edjoj
k/P8m0Iz/3oFh/iBXS8YqfB6GNvHyHBCpxM+DE837dIfu82ngiDPZYmuEjWsdPvCe/FBbxu9OsJQ
yeEk/VEyvRZ+lcTNyDcTVmR8DzepCSjtg79f+4f2fqVz9N0CDMUYW64Eo15H/M9gkMocXcnc12yn
D0x2PWbK943vJPZV29QfTIH8wgMxJlx0aQEBdVPDgccF3eTVgdDzZtHpoVyjisQeV5HP0XGQeOgI
K0MMPmYcyGq0jY38yten8ZyUbBMwn2t6//CvUmCR3iU09fLaPXXHAWJVyURCqPihzQvPa0xS/BfD
5T7CuLvsGle63XM74Pwd0FruPTp5/LvPF4mObihbGEOuURV0AyURzq8C64wFW+PZ9OT40nhspQ7I
+PAft+j1IvlPwzm1XqS1B2IeN4Y9lkqDlT+mgWfIUl19ut84hL0QGBT8WasE91gUmrw6c27ILbIl
wVEsJa3lKX/IE0SRA9eE7GBYe76VMwVFLTwaXi+8dhaahnUGbDZXdVI74H2xrXqfrqvyfpKWCKEX
AwMj762HaKZ1cQwFZeQwmqgfBDU0XdA7KqZdN+2m4Q9dlPkzCEzvkRj7Q1RcEApvW7u1YR87WpDW
PQ5jiCS4iEJe5NrYWLMIV4g2ih1b/CA7lIDncWh/LISQvrsxV1wa7rpGngZ9CBq6y8WU9OZhlypI
iwAuPFY8tnYT8p3uhVKp55hqBmRFbHrHitb4Oib3Ja3kZtgPwvrTOmazj1Xp61265y+kSirAa5m/
NH4HGkEvEKIst0e9lwMaL8ynmTUw9iv4lG9FtedMIfTpDgAOA8/UPedZBEcJkPwlKslOfpiJxPGH
SQjKv7UvAUrSl4IgLVvrhzyL/n6Dk/dRKZ6nm0SP/Sxl5P6opzodaQCkJAFQTbeYOgUoh+IoJcb3
Ifw7HyxPAoIH9YOOoz/PVcUcqcm3cxyhNN3Wf2nNsRnJ+j2dFMN/zjvbiQWRMvZWxVnVbmjspVpE
nFtX+bClZPgAoWdOvGSz63m4uo6SsMl/L94gvo1suBCDnqeJw+M1Qe7h28NbwNDoHzb1WhqkZtoN
Gfv99owc/yv+sAgFKZzSBmdwrdQc74p5Co10Zjs6JSnye39yi8Doe7qAO11hnaCTAlp0bSaQHKPd
5a6DafBp9uHWmO/zAzITabFydJ7yRJ2Frd0ohrdBK7Bb4V2u/GNZHGXdeY+7HhQwXzV/8FmmqOqj
uT5tWmoncR1MPo+4PGLDmzZ7Ab1FVMeZwXAn9nOIM86w0l9nd/HE4Jz7yR88vuZUjldLmhHKvdml
Ofvb0yC6yNwQtQacx5pHcJEeUWm3FodweIuQ9QRHg0vXLMWO/BhzCYG+Kic43PGe1kdL56MLjeD7
IlB3ent1AuI9qSt5QvRk5Upj5AfVYQ50aWxWD/slTqBueslv3x2XDcvaMKHumbMxW9uSRe921mwK
PDtb2KQrSun1nN4ZMl1F0a4wyjfqbk3hWeVtEatUnlUUGoOqLxUzj952uCeY/XCFJFi+4v+Ucl6J
hHgPqgkYuQKG9ol+VGhZnHzChJX0Zch4gKiOY9AtlmLmGFanq+m/oNFL5Eax3LFC36qgSk7pk8Fa
Oq6B2bU7LX4zv3FJ3+Sc5qkiuDJwTJMge2FCYb/yUwH7cMlsqtmJ6IIxMskzUzcVob9jklXkZxwz
9skytl5uVCUrIigJfTJYyMYCLhgSJ98lPFRLLRH06qDRBQOQr7jbgHRq0elrrxQ1ITccbSCSha3Y
g9A1DcJ69REEEce5hRN3YRRhFMrNfz1hnMAtwfnYJCTiUAltjoB4kABUN0VLp3OnU3/smKhvLAla
OtLqHuMD87aHH/T38fDpvsEbY7/MWEteN5wE2S0w8JzAD6C/OGyXUvbgW17SsrcfeHxqny+dY7qV
S8TR/yfyoV0G3xzuPQJHo6h9M3X8UpPf8edAAKGGUNXuWKRMkKMWNAf0kuyTIJOb1Uy085TzwlzY
83eFL2zdAnpovkYWdPsYKPI21CBpM+R6m/ApLg5+Wj0c6QE0kJ/9E82d8qQQtYzRKYEDmFqj3jFZ
jCpYCyiO9eXXQQfzQXA8JRCLgJ4mqahM84JzVh/C6i2K/UIkZa68LUsWyTAoInMAw/v2Yyr0DOwV
zOJMDeGri9MUYHI4SMJ6vEZ+ltMX223q/ajw/FT7LsFWML00EP8ne7Dgw4Mbdcsset2vi+XbpEmE
srHwd3x6YmevnWClqNebYAT78HnPMUaE+EbbMq9yXMfrJnfK3nKGYH5yJMe4Uaw+RrhmpMp2RHYx
QX6OQDA9M9hoEAJLkWiQNbf4jRsK5k1cMugWVM38cHtYnun1mG67K6g26K/klfKkkYbD+iA5CgH8
TPiv370vo1eZfK/+S9wQpBCQxRm5j0oT5YPeZrBRHz+Lqfr1bBqQ5Wr8q05iLTVZefdRgmygE0Tu
v5iPwQcDugpCalqqPE0gzukFLeui5K5gCCcz33eNfrskmbfTXXSrrAdcBsk/eOJylptIwX1Ew2gJ
RWKBkWumBCJzSNQOe9u2ok8ncRq6/J/TtCjVFzCkUWHBMO/1UHFTVeNXHzdtGg6khqat7slZSF5K
S9KPjVKzL/LSvtEImgWmhrc7YYwtUtcpNREUtkiQ8KZVbyJnCxQ5pqyfZ82AZHnsuf6ez4iFbG0a
BC/1Jawew0+hZ+IdbPLh7p3gMLmcWWPLEwdP2CYfY0f/FWV2q4HlxyBAneotY0UiUmSJ4d7Z4WpT
idD/DarGH2gKJWFJkQMgHugHjW9RSSh9qQoIAUQ43j5+GHJ1OSzCW0AaPUVXS6cigMHzGjUmlGx5
9y0cbz1Ovys4Ut9abSWpRk991jNev0bVe21wLlRTFdaH3awXN8leXCOI/76/oL1Nza774VyTrZ0d
RLWcLvwiZpvShkL7zIPLOcKl/ZMRXVDP416+mz7b7+xDb6EC9kM98BzffHSpg6dsEpDGmJHmu6AU
obgIW8n2O0ddtDGFMo0KcuAI3hA0EB8pssNsyo2hndVsaxBnprBpQvKjZ3Gmbrg5csoCiJvEU5gT
wqOgCtDFzVdohwxqBvgCtH9UCW8bqONzNWiYmsO391UxL5mYZ6Lz4TdyNK4AlRwV2/JVkvGvAbWu
W79Ag0w2HYz+viA1EOfSoNcNI9PAE1bXddKaploB3D6qcR+p3pAu93S5fLtIb2iLc4ELby7ZInFE
PizrLLnVK5gzfQl/ymB+cYNTsLU+kFViYLODTVzErIj4S207rDVOdN3LDDxoPrPYkD1+d47EEGBT
8g6R8fTHoW1p6ZnaAd1bPY/u7v436EyP5OCVE/DyqanLtdniReENDYrEHVTIq/Q7CJ0nxxRaZ8P3
4yjrd/qy/Y6PV0NMJJhocJR+EQqp1dJ0eaMIYbH0bRyN7tUqu1ryp0ENUNcJj7ywPYKpkGfgTCVo
PoN4/VnIaS5jhpQBkF2n81JwALW0Vsp0X/cRSci0EcdYynSaGFnR6wQZAj6ZlIk207/APpRgdY+L
8lwVBvsudpq8tJk+90PA1jHpftCSFhmzN3MrdFo6gSrqZcsCRckTotnf+EHcm6zyHand7JZtHBYO
uBLVAR6fLvuuQ4k102LEWkIz8EuXi8QdY6s6rvH0Ek9JkWaZ16s9i8J3BtGR0v/jAJjRmPlEC8+J
0gi/E5yT2ryhBFVCqXqom60XMj7LafSQDxVkgcc48LN7LDM34dqNi4OTreYt5+lfj0xFWtSmjD9D
sL/PXpZIyyrBS9OHv88LvQJ8qVQCL6zhQiamm+A0a7SmXPgiNt/lZxLEdU6RzSEHUrtScxx2cJmE
2PkhceR28jOjgEcjynIGPMV/r6Gb0wrjTjH4TqQBFfoTUAW/ZUX/IMhj030EfsCcknIL8ljMYwgz
ZvK3888dxcihIKXTfWCbpO/tp9DS8EUs6sng3H4FE0XarWrL18LZUOlxhHh+aGqbTmChjD0TU9Sb
bMRXtSz2dX30ICz8B6seBUwlOu90molWhAZ6jBn4Z8z8Q0p3M8WuQocOlGICXP0o2wWCun6O9hIF
Lq+KgTIZNSJya7TrRstGNSk16/Mjl6UrJP3QoC63HqxzTkBxX252pEYqteZSPXDt727sXMK11f8c
nOUbPfN+c8wY4SbrUkuzMP2eHlpDGa4g7jDl8aS9w68Xj8l5zzi10Ts0wvTa6lOwoZawsQDPiEyR
LEyiU1EnOLgJC0gLj6QIDRjW5tSNdfWZVNechaNiewU0ZcDhznp9iB7quPGy49TliCXBAYfOei8e
plDYV4wOyP8e/tzuGwQDbrPdUixpazDlxkXHhbATHgJRY+3eaFzGaVfLiY1STl6jRVICpOADomXT
PIoJgPYCgafgdVyHKqXObq5mbm0EwvvSK7N46lsK0MQlfJmUnaBmKBSSwuy/Q93pwQunsJ37/e0m
V26BsoH9PGRG7u3bOQjJ10qR+gZIytehy4RzeBHS2bbFLs8wjajB/8P0jdYJuhtWwgaQ3pOJgUMH
viHxvPzS2TNZZ6J3f3ppCwIw2sC3IUWu+6N65q8RhP+g2kEnNqOiYVxE/ljEg+JdBkYA7LHBIj/Y
A1T7kBJSIEPaBa5YgF2BPzBoUOIe83NkzO2U+vixUZJlh2j4uV3Yug2P+NpFEnIU+yPJGIbGCIM7
OoyAl7h69GPay2J1nb2VWKW//rZezsJvQ7Km+s6EfEE1PnTtUaWSMyHIaFgmSe4RccZPD+LBOE5r
szCfaHNc6sHRf9Gh416cQrp2WFjmr1QyQUUV6EmJc1PVVWFQD28hnJ18VXFK23Zlb0rdXldzWgiP
W+Qdij0Um/e3vb2CS9X6aw1xdpZ1m8kpdfy+rRaSDIuua3D6JPq6L3eg8mWpKdcTfRCr916NpuME
TpJMeyptMgCJZZ1/vy8AqLN5IcSlvvEqmSif4ihsZKaYUEK2EYUv3NkdsO5YZVlFe0v/5UIfdwf/
FgG0WREZJNsdlKaK3rwlEp8W/gmyQL+Or/IqdMc1H5egQr+VY7NqyocYoXTObBCTbqLvbEYpsQWo
z7Z8KBtjt+FhQZHWrdktr/txVnpVQ9UKSYymp+rcBRkQpamHdpCvsYlzUtJ1yLZ6dJhkyRTTViwd
ib931+e7TCYZcO4Tf5TYHzYYr+TP1cfxgUJkjP9kFfp+4WH2MqD5A3WjtKV2Y0KpUZ1hyQGv5U9n
nk4i0t1qAZ5HFS9GO1jBMc/o2HMQBi0lccZJ8VZ7KiM6Xd3rYWUkWl5AZakm7GKAl3IozZNCEJn+
CQXyIYdmDe23h3CvDJ07pWFVYY8U5VDaw2C4zGgaQyWHUdGOQ1PONQODAtqrIzsNPx0k3hzdxzWZ
coy2ELmbM95jNcpvsG/U0yEHpOBLUGKu5SWZEWfd/pRvB13vYDRns6hHglo2xp8Ou6HkDwZh5nC4
B0BIN08/2n/E0D9xEQypCTITkr8kjIRWF9dVull4/d1yOp5yjvZg6bBoxvMObT88YoHr3eDtxjGT
6cxnxNjiI1cWDdV4I1a3ZmccvNPXL7Ekhw9LBAn7nTTvIqf3ErDYJl8waW7r1FYIwa5e+6U1B3mH
Li4CJvWoJRaEa5OWMXt/K6mlRoEVASQQVHIipcO1C1Tr/Jtj3y63eiuGzhLTgms35ZEyYNLuxt5O
egwDkO/AHoMvrcUVq9QzoPZzxcwBxNsZDKAjTEaKHoLEIjq0SW8fGNQw1OE9gUb2MAzpqjrR+UAE
o+3PKQUArcqlAwa9FTDCQkgRZMNDxOKTjowfLBrjFtLeABv8XpWtd7W7Pawo8phOSXHjdk9bRs5n
JxVqEC4QAVrDkSlPZYX3q+qP9l6q/0Dd6Vz0FoiiuZVQvx6E4zCB8oRYwt43T1TvIMGsZ6yxn/X6
G55WH0L9X5u+lb/sK5UU7XC7Fabik29Zd4pHZ1mP1quST5JC2qsbMzGu1Xsh/4OhflOyHBbfgvO6
FdZo14h9AWxCf5mY7Ag0mC33rZiozAvcHk/SmwrJqdhzerB/jZr/CGYpp4Btf4Qzc5E1RojOVcK+
4bERCzEPtrOvQkq/ujiyKKTon0Vte5/O2lmPllpemMZCSJsgxLIroodivy8jO8T6YWo6Olgn4Btc
aX2SKXwkYnjTlueUelDH0whhht1i5DGD2a82CZhwpGMxhZH2nsD7GwD34BlxVvK/dTCvQpP64Eza
+j9W2QP/yf9Ro42MkSjZD4Wr8hiEYydULUAulyUbhffKtLHLcnl04VYYIWGybXBy+CUaeYT0/oRY
4AHVPcIsdpkGbFbEMxKnhVFrdA7fsH3hEAi2bnJTqHfUcFjF+83XAlB6OSHmDjC8pIaWaubaUSMA
NNt8qrRrkS1ubAnlsEGX9KdojAlzuJqk0QOt/SqYikPqLbZNx+2dWmbX9xGOyWqDHXJcHSqZtEpN
T4rj/9w6Pf8iYc9YzmvlvGa3CmUjYeX2e2dpZfIfrzmu5jnZEwzX+GP4/JtUXyVvxmx/YX/3R3Hg
Mk4DV0SRprOK5BCqhYYMfcvQ2hnsOoIWdEYExc7m15u50PXAISNDtkaHFXJqhG4lP9/wQoY4YOh/
USIkjArtNeAyWxKhw8D7dY7dGkM1e9LD4akVhX2lPWJzsvaNgPO9D7YwLFA5JQ/phVufOShS06b0
cnTeFdUed5rZ/U0McrrzMwBaquTw4nb+Rp+4C8W/KjTrYQGJaqaernwjopuYIt14gy43ogejbCLI
WrdRDvqZC9gxFOyl17jMEWxOLLgMTlWUlLc0o3ZZOJJJCMFEgU+TWks5kOB2z3krfxNF0Ko9pWap
nS3xr3lNI6Vf/aX+HHmLo5Je6jCWGPuQLenzuI8CqoniKlK2vJ/HIRsXusZkr69UpqJCrVJ/EzaE
qcANIN1ef8EaoAp4fjDiYzYMhi2wZPmWLZj4XNua1TSZpOTb640c6js6OZcSxkg2grsGU+m6vhsm
bFnmOE2OBnfdMvMZLrV5JiL9F7qnNoXxvOiJ629OVdVkydoT+Mw3rIHIOWPFuU7R48q17tIk4PxA
LopYTbv9FrhamjjJhnoo+WeysizRr1E8JAj/IRkKT+INCvAAOU9Y5sABXvKUUDaPFcsZBFb5ZhGN
/gXPzlMdeGgicLiNaZlNAszileoZ/43GsayIjjGdn7AG+kk+ACRmS80Bc9KjzriVWfFPThfXKi79
xflNFFCqVCB5sDg+7Fs6t6mQHHNPSnYDBvCMSGEV6gEx5DNhKYtEDNZaOr8KebgmcjL85Dc9HYZf
UUCacrIQw+gYeu/ohE+J1B89gt97wTRWrqgJ800DnvH2Lzs4HEUkP3mQkT2CW8NVNlqPVhuclmlS
7BbpsyM1FUJ4TskWcT8KcuVzUnZTTr/GpWsOZd+i9vOThoGTww/Spf21K1KZbWjKP2z7Fhk956iP
8+6pFmRkAT7OUVPWfQS8a/3T6l4PXzIK22BBrV2PN33HMhis5b+a1WO6DayL9CiAS61mkiB58muM
ZuRufq6vhmatphxUHnd5siA4BM85TnzBrg6xuWKt4D+Bg7ev7he+pvePsOLwJwr1qhI+vSt0gGBF
mRGIZ5dKLQi0r8Re6CPd95BcuXCrGyDfh6ZpBaKJdoiETvuaMaTXIgD6B90TwOFfp5BW/y636F/+
OZPfKZs49tCdJBSDvYefHQGDzFtTb3I58xcRcpOioabbmnWOfkDoPog+L9OKoa/S2cRn4gxVHyxZ
3VeQqTqlkrYUWGDmuh9G60umyVbujvq/Ezv61CtMIWMQcM5QMmFKhQAtik/l+HQRLVSmCKWZDfje
vAy3vlhKC09wfdFX9u7HxEWwlhn7hWZUNNe/rozeeXspdYep95vkdrVd/gY5L0CRvj1cDCrtHzzj
LFOS6BvViJCGedji3B1QhaMqwYUJc2FbqlUDFfDZJgPvuNpyPqfQ85uD1CqflI0TaetMYUD8PlPL
Fx0+hc6vKYFVH4TJ83PcA5RjuHpwADh3AveNWNK6S8tXPIYeNl364goP0VUHdGzbCyWIL1gRtkmD
UO1ZiZWO/IxkhPFl2iVKQSKSsTif+I/LRBlb7mApmK24TDJ0EwEVketAq0MMQ6vfTzOuz7zFCmZ8
XRUPJO3Rcj0HyVIeDfZrEA8jNwtbx1Fqu/CJdtwYhcACzaG3hfbqp0b6qRkx9cdKLJUeu7a0yKvF
mj9HvJoDsnwzsK0ZcInJ/1VKLeZQkDqkDAL1u1B4ddAzsdBPpZZgL0apxy5UMd9wn6NqNw/pq8Vu
oEv05XEO+GbodvuYgujIPaiS0blJ58vKKn1goDMy5P/gjDAW5ZNrZTEOC0z7P7aGd3QEDNlGVvM7
50DEyYhWlDt/T11SJkrs3zJyTzL2iXhw5/aFXueAHBDHOwDGkCVfb+4Cq3Gw/tBtGBK0d5yRae7s
y+CKEJGaGKnv4DKCnjj9pd4k7ECAXL00p28dGOwt4EiEVQHpYM0QZP3x/Zdh1U94cBQP9FidCbyV
lNLev6a2U3Ey2BF1ZT1FJM+0jdkfRFJAzQjjkTPXQzDbaOZGZDfg6gFKrOU/BFft5M9VyoUZ8rzB
W8L+sN0IhAxiCbyV/dnLmr6CztWaYpJmfHZbWlaBbzlZvEbRnEnZG6jK8IZLU+ni5UxC+Wd1Wjxt
CAYtQNer9QlIgDVuNKMP/5D2K2QODp1hXB8GQkesP2Cq3gRnqjBLW5SnrmHbCGvTejnSOQfsJJQ3
o+M8bEwr7yMuk+/PDD6r31LykvxjhKqEawpN921KGlNiRf5SaUW8cmvcf6nI6vzQIv0lY8F1oLWN
/hVR2JvPqqN5rijDPzmUYYRnwqj9a9iQs/364xLoBCDI5PrurD0Nmw0erCnshnHlS5CnJu+rTnqX
QWko8G4Yd7UGJV8YfPM8zEyvs29B51CN4vT1WekK50v+s+7sVdQtHJsPVUy6LrBv7OCIE0EMJ0Ox
A+U0qBV+kbA185s48sgNlLFX45VsfydkxovrmNvnMyfpti41graMEFVtfvvGqLxCUxOU7IdzFcd3
FQgQCHbpQt9AYH+/+Pg5WtyBI2mx4ZvVdxgLfBYwKO/HfOHqePDZC5Du6peGkVFdQnalPwL5dvQr
iuj0D0prE8imlfRxUq38DkU5pyBIYF/NEMlaibxqQS32ighl6mlI9/YL/1AebdP+VxggvNTMNpxX
QDzGLNVumfp9WTFBmzQ4x/k+wuIZx/0IZVs2tfyOqPzCbSvvi2FY9s5JL94whqu8e/ND21queRU5
p6VIzDJ56kbaPr1RCOcEs2wd+v2ye/DUVMoqH/qxqh5OEn+4Q6zkQrEz+hCdWNwZt/YbIwykGmZG
2xjMrmAX8VjjBt+2mnB/JcrXXggAAnRHu0CVZ4Q6pDfwC9F7M5L5TaJmfhAQpTMRaLJTjdBkRiTy
RSTYEzIN93HnbFy6FUF2XJx61Dtj0Yi5YLFRCrbCusR5JXeZbsisMrpqo2dY2/DIV3qeyikJVtfM
p6V8LrlTZ595s5YAoZfIV6/sgR+iueUBYVZbvDPv3P3GC6DHK/1RlVyYXD7q36aLjHytOqAIZYnT
vNyn1N3w8WYGxJw3HydT0k9gDK/DkiRfyD4cZB5MuddM8H4ahlxe6tivoSVy+QK6EuGoUmhPDEev
gX10Bwdt1vL1jvJVsKQ++NmezGWOEcwvN8kr5goI5JY8U9XGVaVNw4uglpad0SPW/Dn3hK9snyrD
IEdpQjfgfdUGNZQsgP4HJ/QLUQrcAodeZUBqgK4LaGc9RN+D0KB49dnjTaPzY0RKPS2foMpq/lh3
AagYYoT1g/6w8NEXjOijIc4sa82p03L6FnTdRz4KnUvh4SunGqetbk6dovbwRyaa63/krFFM/Nym
/1ogL7lYV6XVF82mjd1DiqD1aD6Fln7bt4q9GNP34D2gqvF1HmVOsuG8YGhhPeKL39BSXwUwJc5B
BkpvMukaMf3dwgvmPkdMr7OEjRyhNMsZiRkVRisVQmpELe0pOyJclKCSHuTacLUmknmSqQvo3P/s
/TUU0Pfcsa4H98FfjTLzYMqFVqhehSGIjsXQgzQ1UEeb/yUTlKY8HskxHemvrvUipQ//J6Qzp5Jh
NX04kmgG7Uoj/Tlpf49pEeMaMBm452pnsZjXKbKWUMQtv0E0z2jA7AgG0d2XQIKfbYI9ozoEbmWH
QWihs/4uL9IWD7pcA+jM8UxXz/HBbJcyhSY4X8neOIpzPWI6PsdxpVzxZ+/gpqYWk90OzCXUMEek
2S4LKWI6dch4ZQOFaMEeMNmL92tKon/WGrD2TsvQyrYDAq1gLqBmpI6sxcU3l4xOHtlkA+DWgiON
wI2W5eRs6gpH1L+w8jzBd4KqMwAZokpm6PpboN1U+G/mpXBWesy8K1u4qxoir7JCaDu7V02nW0tw
Enf5A/XBvctSfYh4C8d53euBU5cJZFyVy6eYG49uINeqR8hBxgJeazCgk7DLs7qf9P3v5zpRtmH8
SkN31Fd30BHQOQ6K4nIm/9kVznEG2sGRANT8xljVWCGXhdLRKO5/OJxfR7OOt26X2Wkg7FGXBwzv
jXtNUNGG5wybIMO9ROT4Unmg6DazhRsRDZ02lLb52fvHRCE7pWyUhbZnl58gyjY63KBLqBcrg9bp
ta5BeicD31/lBBG3IDxmjoKuUi+7TsTe1T1lJMX2g5P8e+Mt4YzT+S4rHcUq9kNLRBj5YhWowW8H
0Uz8Jl916Wrk1yeleKSkYp2DM6dUbceY6knyTMRI7pdPOXiuQKV9QcKCe1W/O7K5SAvdJB93TyYS
xbUozH3bWSjNqt3dmAocYHMNqwVdDKQ+vz415T/Uep8bWoPtG9oGVi32H2kY9/VXwj1imWdXaSex
DKxZu+Zzp+O2a4ejpdYaALf1TbCLq330nrDOSoq/XgrMvIJfrjqwITfEbBOuuCPRafjg6Z8Ws2R6
gMmrQB80M/ajluZVtrGTq70hqutmfh9BPh1eYjeQknass5lhTeDZl7bz/6GvscS7k7LCAbIQM3ue
VX9vsOalkme5bfFo0/r96/r+dcIRR9dKUQPjcAHq/xTWm2pIym5CK1d4Ypx4CT3unS11g4ULp9Jp
ctCICdHdzjW5ZGRSU+6XWAfX9Vq8uBpcyXg+z/wFLf/G2yHwZDfMUwACBugxsvpV++aNEitMLTcU
GI7DGZvthiqq/3Sugy0iKAys/l2ZBAYrX+0XID1XVtqlMntMpqKkssfPuw/NEjE2QCHFyYS7Nqra
iUJ6TA15q7vOcwffTjbyLjkjbT72iyu/0ElSyDhLBO4M9gv7eDYLdnhaB2AKA1jYdUrwpWa/UPlU
KjxoYfE2/xDzbe1z9Z1MjWwcUKlnSwSNm48JblDgcjDybcRK/zZApbNrhMM1wtjactP7HFiwOymc
DzZDhATJ0cBd7Rtze6lf0wydVoU7HKWJ5+atgC8w3gnELV5ETesoCngM3AfqxnZLoDcjioh7GAFI
k1HSlaDqd35gn8kNt8xY4U0+gsioxBdYxbmDUIycoRGGqRJaSuiU/UjAGGyDP4CCe/MuCkOwzWzG
/fNPs/Sx+a5mLch7Sy6k/8KVl8HkMp8/AQBCGt1S3tU6M1mnEYV4mWL4YuQ+UkqhVScNtv9mrJRn
Cu+q8qaSsfdRRZpfwOQTvN7TyCMx5smdCwReQf0+DVuftWgo0wsOwuj54mwEFtKYq71mGVcv7Uqi
MJENCAaJuB+WPLavws74xk235llGr4B3ajnvm1/mKiZDcVFTHf9ZcCN+nA2jpZmhAtUeoASHPE1V
X+Tyxv+U1Pt3VAohYzyMwWOwBgLCo5yJa+XmISnwCmSbKJ4z/UmTUlySyc50EcMOZTS0nII4gdFY
sK6vaIHxr+w7Px1zYaVb2lLPJHP9B/ONunGs3veDefIwM0KXFgD/Rfa91gEB8A2zsLKS5Qa4R42x
g6OZigRdcqHD98atI1Enj+Xi3XxCoFYBzQ5OTiM93SKw3x7WyhqwRiv/WseeaS4G/pWu/YxMSI0d
5/qUTyZ9OnCbfSLKAuoDQGHgzdzNu2/siaKsvjMMc6R3EfQAX3DL1dLDjG7llA9lh+/zXNTXGtuu
cZ4O9S8ErFvb9aTC9K8nhrPhFX7i+qQcfbo063SOZR0WzRnRBcx43B26lliNzd60edhrfYkUMcGo
zOhpVjZd3cxSFWBgg6O085HvcZh6zGKrzQ22iMxCmdVF8uHTExhev6AnOJZkeJD4/yTAzyH9l2rQ
FQdXz0FH2JNv9C11LLUjd8IxVY3FTHvE51bUktLd9EUtMCeMFt4mW/6Tugw//MkwUKv/YZb2lee/
uYkBGicXDoGSr+p9wCGy585/KfJr9baHbA52U8bXSEL6vx9Biv18TtcJp8woJuT9fEWwMnkoVAlj
3ceEVFJi91PokMPZsRTs8ixIGH8BgYROK6XA9hUY8rxvGqr6rAx8CIITTRsTsEM0IqpwDCYgqko+
KPfk37LNkDujaVfGkF6H/GeRiYijhlQEyWOR83uDA35O8T/KUBCtuGQIC+szkYFgll1MkhTqfrKz
efBegflW9PXCdC7ZVV1ReteLV30WU0TSNAfSkOygKQ+DNsX+S3lToLb5AixX8QUabWSwvJlNYvDv
k8NdpArTIvAKdgh2USg7eBk4Toa4N3gwTFBeTcTkFkUheqPAlaVwg0/0EwumBmT93kkBVeX93cm0
k/fCyGnt9JeFwyJLMSRBuGf2D0qcL4BhVgXYuh2z0iG9bBszdRjYYUSVG2is/SqsmimoclIVphMx
w6ddnAK999mwqBkyqIH3ztnpr9vTbzJr3TN1gUY5VnwhlY45BefsIQkNTcnVMGb1FG7EuWjWJlbB
224k8ex3ALU/fr13rUf5AA5oa06DolkUWzEt5/LZwEUBLZRg3Szl9xA9lzYSwgYpcWXtUxyQYTRQ
V9l4V2SBE1PxNpbZGoYUjStp8zaBbOWgqsRbsTiXqFX1gdOop+gaiBqbbLGmGWz5Lg2ijpjIGvKV
awGuZOPlJUTDRB4zThmnGEurs1MLEPF5zJ3oo7d1w33B5nwijd5gEVw6VyJRtg6q7YLEWCSwJf6d
fHnXitQC6moM6+HvqUChAPaTN0pfn6JEff9/CLVDymrF72ayXNYo4HPiQ8ASy+fA6jWkb2Hg6vsl
wGgvK0XEecWIZi1mC8L+CTBbuVrIe0bFbThGsUNp4kZF3abHHhI90kTtSkJHFHQ2y0u6ekPN0D2k
CqLwxFgeITbMt748F3LFICqgR0lEhKjpEyVb6Ib1/jtnx9CM7OJK6p4FgSvQTFQd1Q2r6ddA87yT
nfsVJ00TiDflmhOPZjQF5vuKGpyvc6HoQJ1PLnt1Zs4rqhG2Vi6+s4Q8oHtE+6KYuByRBOYYy3Ma
6mv4pwCVuE6S8Tanm2pS5964FDWdHUi+PZ2bZ4ZmmUyQwBtzRDudRVZlv4cZWY3kIhihrRnulEUq
Mftd+TU3KN8Nf9sjduP7Hxi81dIEagk0nPh9sVlOZ7zOKYqwoJNKTQF6igqOkc96MlIMTF3wqmNl
zT8a9jqdlcNT1o54Yittwk7Yf67dBJBgyMcgAIkVBch1kUMoLf5dsPoXYxPGuuuNNqhVT4NmsLEj
RODfQvXT8I7CZNF8wNx57LqhyIvE7pVg56s8xFM3PK25q7EIN7dQ5ZWeOaXF9+ZO2iwYEh9xfaV4
AeOKSlr3gq0f8HIwajYI0Xo0Ao9qfbjZEwttNma31CnIuCenTg7Jz1sTAc1+uthyw/9Cma2JkFbG
E9MxGKzy/Bg/WBcYpnPrqKwp0ote0T62CFb+h55akupylw/zpFH76b133iVNLl246fP/0tCPBwQB
NitLhH0xAG7AfeuoFgCHafToiIC0IBD4KB6A3WhbfkjtRF1tTsNyIEWqnDLEsgdl+KBxE4rid0Bp
dIeqQFAgU0G0QscSQIQLaRUSHWfgZVBA2ARCTmrxXS2md+9Rgi2l7AnoYR4cvdTl6Emho5+qOWib
I9kE8AoBDBtUD7xa1D+/h1kCKKb/cL+g1rVsppgUsOhSwXFubREd3Nic/nb3zmf5C51mdzU5LbIW
OUe6H/9Vb55aTeqhQhjbJZJZLabw3AlbOxTaGGqUyeJnelIxNwcscBx4OVHfM+O/Q7pp3SPzuifd
AEUm8kWcFOvbo2xoYiYBiD64u+qy26j3y9xdnU52CgDE5AIDOBOlwts1OlJQp+bIpzbMEA506zSQ
0aL2iYtLVcNBnLzm80KrR5aNB542NFpelE6iG2fF7KgZPOAyOdVkr3+YDMpZNYMnMrHhHkNKG57b
KsphiXXMC2NK7cJbmRrnM6k4tZjCxm6vKepOv7ymt3RAtO4WT5422lFdMH0baJahRSgztbH64MY6
TjL4SFQYsE/pfask2vii5kuayEZLVg5uVn9QZTA3lo/pWeR9FYZLszza2+bQ7NJvu5vSuDcLhBp+
KUiCGTWIZVmULfs6WN8sflzBaltabCby8wBM5v6K9sS4nYrmHvTLt62IpLdVo2Swjo+BpYhChVdE
guMm35LeFSLw7ATZ7Vx4zgJGyQgW/R9ClJVDq1rCHED9OxzBSWnHKIrLK+zeNoieiBjMpsasANMQ
SbiQtU3JeXQ+mDBsLcUVnuklbU3H35Cgzett1M4M1Jcu3q6kds2PDGz4nRDVlw1D7SGz1oLZ/UXq
/ZB6iiW6wv/Tza0fitDoL14XQ80e6t8JyEQFuLsARa+ypMq8dFe5giuErR2Q1fC9D+lCq80Xv/dS
odNA1LGVzrz0pOlZrAdrACuRgGjaSH008M64YhC4hbihooqD6T03Y1MbKK1pFV2R9w5bHkP35B6D
qzOdyGb4rojHyhN8+bud3qvjmvU+FxL8zU9RbPcv5CkrDs7REEFHSyQJSGfeXGPaYT5fDn3qKrkQ
sQIMYdM2W6aESUVTrLlJacIG+dElgkBHGBWfvSFfgOUzzPq51kM76cGMmvrk4qNEiFNHdIZJR0fl
+EMOLA7LeWv4L82GB2tyD2UU0bp/mKAaprK58fr8RP2xs1EmWnzDsPWfMWIiLlKiMk1hbZ+cFcEj
wmjO5kboOwwY4pNfUXtAmESfR4cfrdb+ZEmp7nVygqBYFDV5GA2SF/uuWmuvD0N6eKW5xIAHtcaF
DgMCO3I0f2F68WXp3yBD7eMwEw69bgPLTV1rYlJV6HP6GicDM+fbNb1sTX9P8ENiZCRM+HoVwfJs
wcxQNwVmpK9uhRTbABZNG7DnGj0FxPyV6MB+4oMPky38LNoWAz5H/2HPorvmimmHSxppWXd3cGM1
IpDekYpgnqXbvHnavwy0Qgl8oYRDMwiKlNztQe65wf08/3Tj3iRdtE5GRePfkG7ODiC0EviOSpE/
9nL++g+CR8q7sAsOkShfK07pvzqOo15PNQCDOz1ombTjzyL7i6pngHxxC9QkP2vJYikEwhnzXfLm
w3aEiCaWVlwyg7eDVmKxFTf2A4earY1tSEpjSd5JDTnYTv0GWImlOEVzEDb9lMlga1pKesP2Me93
J6RxeNcUEKkXfbGxUD7ByqscBQswW7vEQv+/D3PHI0K04J+R9Wu3ycxMTHbnDSjdZmkPrljwYWCX
IWaPbI9+5tquvjq18uixBdMwHB+Igqt61mI7ZL3ChoK1Szkn4girg44QsaqRTbCILacPt5Oh9LwO
5Q8Jv+RYwLkrTm1d2fXSw9Ja6/5XJYL5nrggtuBwGLW910aNcrEq3RwklFiDszrYi9TouQ/PTnh3
XIQ097h7w4N0XQ14knFO5cABzuchiGKuYyOjUZBdH6tdLt5w9Fwu/LHZ8E846wr2p3P0M+sPvkZa
lMGQ1Ve2FdQqhQuT2CKZFOqgMQ91VlylYgHcEvEvBHPals/5Uy+FyLNXraEgquav+due+XSGsMpD
Jj7PO106jjNIf7S00tEGxMUqJDlhsQ9IcXbw2zTwrhqND9/TqvTtDI7s/+8CaWHAppgRV5xxCERu
mwNUN52S24pOEEIf2Glj/iJIKTWMBbEwe81jnDlLVDLDTL3wMmY6m4mlCeu6YHsfJUz/j617JafR
d9dUlA80GluR4YMGlXHlMASGp82x9mxi1lT3B0erXp8Z1M8IfDcujooCGl9whEbxsP9u7hYmJ1WU
Z8c4TYqQM3qRg+BOhaUgvs7Y2C/s6UQvKk4KBQk+ku/jD9Evb0zrU6cL56J5YjuoW9PLq/dtB8Y6
uGFDVIfqUopozHVUUHX3/naRl4Z930EBPQXYmn9ITSJ//I1HqBt9u5c3CaAUjbVhEj0eiN1otLzf
Q+lwv2lgKqC5imESe4ApHJdy/fhRwAqWzExtoWeFyLI8SsNMTRl6nqW6azFqbJItq0MxAjxy9Z66
oCPvFz3O/ffgoqeFKHfa+Es3jVzdxL7wJnZrz2AVqzimSoF1QHg4UfdB9pHcb9nF9ixyjchgNTxY
RNZg+X+oC08VsG6LQsws0VkIEh4HRqN3dj38QXZoVEsodx1E13fIXCmBrZLySVitRHDfsjk5zwM+
1Hptslga9XFdqtwyMHCtXVOI60zmnQe2h0X197SvV/ujEhCAOXKOixECTV3sg0OynofgFaaywMqM
YdPKL+DRxQ3vWldwGgMUnP2g3IffS/TgUcOPL3t/4LhYohxOIHjIXqIDAnqzkln9qqXfX8CcAVTA
q6a3JdQgslGRM9C7c3M4K6y/R6kICLqFIlphUjkiTp+OdFxLIrNvn7SU9ZQrvhjGev9pGOE85y8B
2mQ5VrhN/ovoRTuPD7l5ptqKG9rern7xkpRxspy+jMKyfGXNwmjv0vufbxSbBdu+QJIhN7Y46SAF
evkLTpi9R/36VsrRuo8wWPM6CN79Qgm0IqqIW/JbD/kQELXR54Q1c+JH+oVOBpkLbY2oCxR4mOeq
7AQpqCk7+RkhYCW8nukQX8vgrY1clOMnxGJu5a9r6+hyKU2PTnXGnIzjfR0qd90oLWHj9GDpyv7K
l4wElF2GhR7OvYQOniKb+bW1Sw4bP0B6Yr5ooDHPP4+r15qf/CKRwM9XN6ylcZHK7RbNbhBjSq2L
uW1fVt6yQQqvQ3KvZyF5UwHssM1j4AVBF4RXdO+cHa0qP2Lgz2w+wB8mIfDtXDB4hNhsvc97CYpi
1SkKHT+bApLGjvEb8pa3JLZRBAuldjUsaY9RKaoVVsU+W+Avm8d0iQk+uJxGY0Zvf7ejVyk6p1yL
VX3Gt9d5okZbTGmvc/cf+qcVu3CNoT1oOBVqwkgymH/nWHR0w2MTDmKMFfMdHih3Bssd8DhdJfCl
pTcPb/ZHLUWC7hlfGVRwVS8yBKjCoi6Pu5258c9YCbtn9GBc9gLP9t/osXtFo3u+8suFqWZ+/tEe
+cI6bZm1CzTt9+IX5YCAunwrT0c1ixBYFrFTZ0xcQCUTPMvIJcm+QaXAeqN9Alp9C5uE2JDo0mvy
XU75D3H8gaoA1Tj2GF1/ZItcMWRkBMfKHwAq49pxMC2pUdVNke5A3gJFEMlOLxdRXEpeWL0mWA2N
prMQyTxIa3JjsGdNF64KwE8o6UF2gBsHcaPI1qJEs3RVloB159ZMaEj2NzwMGd+f8zfmesO57F1y
er3N4C9G3jSCSA0jL+URseTSnTWqoAT6JqQQGDK96NPuhC0kvnsn5bAYyHRrWjIL1fnY2rMHameb
z8bIpJDH0nyCn3h9PbZ857NoegsSxTLHAXwH+OdIdElLd4JyZfqRgkotYLxVSQUxyTnKrvFlFH+C
jaRpT4U9cwBa4P7w4kvgmrCUGfJ80euBqMden73nhKFvmYQab+Iy9pWmNMRPw+ImPG8+GkUEQ54l
pdGV44lbJk/5cK4aqVJMZFKS1uwf3Bzredro7++51qbeAcPHcwovWQ0qMl3E6Sy54UWdVjfTtFuW
s4K+2laS/w/dP4y8P0STnWqA16zA3iktn2nRnDddkDOo0Jy+s4YIv2GLuFgn7cYtBPR8ApXIAL9Q
iZVaCVr0pYa1+3Mqy1wihxfkJI12nxiO7lX1oto7UMq/aUkEb2Dp3jiFcwovQmvHRHNSrK7wUwA/
xHSmk4ViUSD6fK32fTlZ5Vy5O9fdmIkgzSEp2RtJPh+5xmDTkBH+Jj1/Od3ZnUppKkvfcD+oCItw
MAD2od3GN7W4ndvrqC4kXAi7/++DUPXObGz/EHg8LU3C/UjNLe8UjhVZVb08+G/PerflKyjuqZoo
rwI6QBKQ4htQIDMfbO0JvVs9PmDr+nx2Tui6eMuNPhQcaVqohEOJUiJ3caYwght/s0bJBosJ16Aa
1mhwPNcUalQN3naw32O1wqWXX+2zL2kmPzXlb8/+ITCRpoNzKYoHvuKvwa+Eg285QWMz0oVAdMJp
189Tz3g/wMmqdtww9s+BKEfR+mrEprP1hPXzkTYKgL+8JOWlnuNCmf91u3GTswtrf3xTWegl6J+4
swXVKjIci0dMHKam6OUE0NoFw8/pCFtsxyp2M+I1/Qxv+J/NWQ80NInSmZjUG8ViGRS3bQiKXlqK
PA5CrlQUdGvuHy0/LHQukgSlgFH38u2As/edtkhyRgN/TnYRITJJAzgKku9jUpTyMvVjY72AlwM8
YmQ+vioRJm2GBIGK/PxmoqA/gda2zyVpa18Egfj09WkFW7WJKm7OMs9y4RoLJoGdKGtKcP3cDa5X
BABwJtClqusLNVJQyrn05PWM6qeZfK9lCc0tuLqgPrkPdKjPrJXFUDaDf9czd7PRpoy72+mzP2+F
JhE6DPqVm4hi8xp120BXXzd9EWD5WZQEEWAsBJ+Rx/U+7tVqPNa/GM8z8aAEZvv4UNfJoT3odNro
ImPOxkRR0ypO2uAcrIzX4Tr5YYHNoPj+d3S+YiDjcZ/NRgOLCj4abd4b/2bbElIMZId5k7nBZjGR
QaXz0FDK291+YlvoDlXHJHShfBP0F2ZVHwdo1PgSUbiah2OxGXX4WISAFww9vLNenWI5Qv82GXpT
nNz+fqNjcrd/46rc18Y1Xol/wa5FzRiJYpL1l+azDb3dqokg+nHcwj5q/WLpmFkP3Wj7KAmzQrDk
hW/op4BEX8VHbB90f121g9aHFIw69bGDVn2DDPXAd42s+Fj5FPi2hBPmIY7yHjYrn/OcVtFt2DHG
1R6erKjgYgGSBPpAupC2PU9ZqTrluLv6ICXRvcvIeB13J95rA0xQam88xvD4QG/4UhHXVXIaHJuh
KFrn0raSKIPBkjdYMvAyfc2o3eY/YCqv1MgHE/8BW3N/eeM5Rl4m+2Z61mmgvUQaBYAfp54nx3Gm
HJ/P0/CISM6oMMKv83O04/EfhoZ9yHd0KYjnxb8+CRkwSFLh/byPG7+wzkvrrmAF1m+v9k58T92A
rUvbEdNqHK0TctVqMSzXaz7cEHchPTSh21oQRWsBnfx4xBAtJr9qWNvoN9qKt0dZ/1YIYAByNzhC
bWF7Oww2MEfDXc35eyyylq1mfAw+1w8264KFQ5VBKi1riRFjI2yKDDt1NABLDphwAZTtOx0AiIjP
YwZLmKn+BUvX/oOyym7rJW47xn/2TWGUmGWFyMroF736+upYzICzTCFs+NqdSMOJm/0zvPrWNmLF
f6C9yVxQ6qq1QDXEqsxUphaA7mrpYx4dNX0vDm1p2FGIFCVXts37U2OMwjOOEgVrl1d29V/oJ4k7
+EjKhbDlizk0o/GbACbvPOCyfkMhjItl7Pke46ZzLrWQHt2wkhAE2qeEkDXG3MIS6TdZHNTS833V
xF+f8yLn183QCTPtZ2pBwiMjF3ot9hm9FTgJ6vWsXqgjyZlfPE1I6CgY3v1v/alDISt02dqzKfBB
lFg9OQ7PIdfGVg0O9pEr+GW0sHMrPfePlEu9ayN4LX3+9VeLbXAHDKAK+p6iDF4FFZ3T9ONq/cXw
HFk4yGP4mEZ2k4EsvAEC1KbWbDC9cSQ3WZiQ/VPWrs30XASsmzwW1/I0RlGKHbF9ZgzVycCUx4wj
OWeuqPqnChwxhErraJ2K/MglwsO+xLGFB4DxqLRA/g9Mu8LYA8ekTukLBkaq4wcxSV47JLo+uFWx
CNvcglXnpmO1y96D00oG6Bcn2UJliU57w4y311LkA2iW+zzGS7wyIg75T8WWK8OC4Jy/pIjQ/UzI
yIknpFm3GBeBvYJTqXH7UuJUcF7bB3DaMHVGSRqLVQByKDF8jq9uXeV+M36/2eWxdzCz83lLTitx
i78SvJvkkU6iE6uA8bvLoCrKjDxOkskTOncrJWc6pICzzE3bG3BQyZ5NwZ+99FXKxtT7Vz46L2Ma
CQepVU/lcPLj5q45KWO2bwhfFg58HSkrVASHWmgzZqRZ0ig0sM3vvDas6ZveQvjY/LL43y2In5mX
BOYb9ygbRYsTfg8Jyu/+V0M3XrnICDxya9CFIaX6jGpypZYEFzK339+wD0wxeSNNjSNXsCkEySgi
WFSkaOIDXkkg2P5pCmDkhBDaRdi38k8WKTiUOkjMuJlXLumGVe/Ta9jHEUho31pI5wfJ2/EzdO5o
xE71VSTFqUeAuh/otu/pny13cml2bCokKcwb0AZj1HUk8096fHAIaANX9usHARk9/lWCm05VgTsJ
7DnThR7nspCVGC1uFT/dejOI0EkbMI24FsuSq+lMAM0Ym/fzXFTriAeFNQk2pZdrvYhCh1TYIZbv
o1M85mScYzSZvHKOxrdYFWpJkj8xuDEE1MncushTLo2RTWC+BrAWsysJ0/8m+KCUOvo0NFVMajsI
IfzGYVMtBCzyVFE1mCYyuVvM0y6clpnWr/91yihFHTglVfDcl48By5nhCcW9WThAN/m4oH5uBge8
Iqb/GARhDN3UN1qCMEAaisH54wvJF3B0D6DKZdkoGdPjvK2AU88+ZWlXOaBrP6R5oDbeM42aeBZT
UhaJ2qo9330MShz0sLSY0WDqW3rXqlKSJk9dJ8pxJ3yk2tL50EmesxfUUqhGEL/JO+io9x1wnMg6
+4AE4HMFXBgIhkNYYCCa2faz1ypYXahFY4HgyO0WLNsNmRdgtpG2+hNFzOgEthhItvWGhM1ZSIuA
7Uzjk7Zrndbn1B1iePEAW8KTxAL2VkaBHUXZUh1i0CgPbDS5M+djnHfy3fza4C58G1+4e+ITWDBR
tlNLPtSXFnFLLwr2Fuai1IAidYd4utSIdHRveSu4/ISm3W1E0i02gCL3dSbjtNEu2d3HCFDopHjo
sWhV4cEHTv9wjAe8T5llw8X/DuTJA0XB1xcUlroBsiiOGpjQd9neOK38ZaW0tSYJD0aBLRA22erw
F1Dhi/8T+1i8My9S5ZY9uweNGLQwPa8TuNqatOmdtJ9Pw/DCollV8pQ+kGmPjlzYw8ZWe72Lzo96
99m2RlXdiee4fnvPtcTyeF5m3cl2M7uqM4YILq+ESm3c+JfCuUrIjCMt1U5njBcAXSSxPc6f1IoK
Tcf48sBKWzRz9H1WzONQK5E0zANnE+O6w6qbSthHovVbAnOGEWyt9xObUypkkUac/LvMasbmhkoE
7EHGdSkmY5gxthB2Y3tjTMNF8Kk+E0O9bq11YjrxvBDUPjdQLb71MVqsv/TNpPyUxU8zqhZmYJ5J
3EMmWGtgrnRZMXwBUKrkRBS6FWO4UrpPx+r0TzKwn5IBkeeFbNQHjGkIa3kEpdzROqH9Di4hkv+1
biKsvqCcqu/qydLjnldp1jeN2KPV7hT3aztln+0XGx9nbsiJqAEkFPxPLcuMszNBW0l099mVU/OI
bFtIZym08r/ZMYL55AQe4VN/Ub6j9NWjNSs9qEwG/P3AOl5hwxFH8dD/nw7L9b83Lj+s8rMqltDq
38raFhF7/c7Eefd2fhXozuQTpORnpiUKYXmxwleWojBRKLrHSzgBcmY3IDOP4Mo9/+O+/00Nt/JH
Bedii2vS53/Kol7CXi/DAN/soxosEq8b/oIcDEJ6pff+T3YWpAb2yWjra77bDQa3kob/Mwj2U/v7
d026xzcYuOMv6cgwqc6+nbANj3V7VeGW9RFVU/fAwuPVAiFP+6/3AZq+Wzl59td7gmudcWFfQ3nP
ZjjGIUyDdrfEduBl1PDfjPtJU6ODZAF6+50AkxBNB+LfOet2SXSh2Ov5OZ1P/dcm8PL2Q6jdAiO+
qGn1G/43A/bMYvkR+XsWGVVRrKCkRePnV4j0l2y6CxXfi8+o58GODyGoUwTxewAkkoNmsDJQlDHt
urWnmW4vsoxt05Nflpv+ilYAhv61H6j27eopBJ0enYfOpoP7ZhODVaessYsvmKwka8D2XMHLiDbj
6Kq4dTsaBMfmgKnh3mOBIkccB6FbXy0KANz4TOMcXNxqPN1fy+0yHJBORl+Hxcg8S58fmAYZKrBR
7cfjj37LE092/U+8lZKYRmt/yN+SXWLF9LpoIdVe5TskasK74DIeIYEva1GJlD2cvxREc+TKKN0u
12Ppk6il1FIsn5yWVd16zQtMuN2FT2ccBIlZeuFT/zND4WhHblCeym0yb+8E5ONBfL4WiMgEfxBq
g9RWBKjqwjGScg0ZbnrnvJEh8DLbtppoMr5WYZtfDB/9dFc1JCZj0M5hP3ngx8ATMXzRm8krFrB8
f+8Xxw/FnFDBqNJ5ShFklYgnaxJ+I7aDe3nvf2PeTbrRoKLT++JSUGOgWQQALi+SoA0aifk2z8lG
dUHpiINMgE4o63N1GrKq9zZ7j8YdiPOBDta/V2m3mG6Q0f8Q6a6IisjsbG4oJyGz80cxcO/QYaeV
j8LWVYcBsHDv7APrPXcTONwuqRrpax6muaqAvLua27sb4apI9e59yQunXyo4wJh6rXFRs9BFS9Q9
Vmf1D535DI+k8TxqGuTW/ic6wEphnajW6wKyg8z6DId4KmNtrL2LZioa2v/915jmRAOiD6H6gv8q
mwZl4fZdqrPPkRauuVso2e52YGIW8J2Tsc8CFp9p8qESPTeCYtUf8eL1+b3HeC6/F5EjwXKrjrF4
SutIaD62FlOS2/e4/JFLUHSvvGYmjgmEN6n19iUAV4DMJUyN3ayFGhASd4gzHdOwRM5+azlWVsfu
2xCGC8tMPbItdLgpPjsa/bpk9Y1hfXIrNG3Z9Amsi0mpHvaY1S2E9NKyyQMC4tAbQdtKU/uW5voz
LFiR+EBz9k7N43t5qVjbRjawuItd7GbcD58LG7qBKRu+lvhEpRluajede0VS9VaPtW2OzIGaI2gx
5R0/SvTtyP/ozVvwEPIjbj4sOQ0n5ObHMrHJEHP4FpEYmh+bm5IH71YjPGyzd5r6/iv443PPcp5i
E3YyjneMBIV5ItYdnB4fiENgWEpflZ3DrIDS2Bi5eF0HFKXlImai0g5pBEalbUBibBKAECp0saMr
kU+0YHFAfAy7RKF126NFUpSHKlBt8N0LHrz1P2c12clYsiCtlLLy4W/qC8LsmazL5KwzZbtS08OI
4M3yEXvNLWB/V1P9G/I5yUjd1YiOAzAP5bYcVJGoTpzZp5gjMd+kLFdthmCM91GJWlppz2Yyr2gf
OknGHE2guss32OyyhaPKJQTFqN/Sb/5D18tPSjd1OBuVUy3szfCsZ7MAoFE3ULsVKws3wnibPtTD
V/t0If6cngqTQIB5MZWiQIEwNdlep5D0A+jnzyDnHjIjMJOZtzB0TLBO/5v64hTMBSSh/6aAzWmw
zr5nN9dMF7zyXDRp9TGLpg2HOeL8xCB9VlyV3NBWoIapGvqE4R6++wydILpE0nKCihVJt+IhnWyJ
zM76UFsT11g+UgUAqvpyG8VLtNSQcy6yXVHHQ2sEKEEbhPcYIETe1tjY8CWdq+N4jJPdrUHA7I6z
2Lx514/VcX9J/kKSsbIAaYQZhbxR5EVQAZ2/3QUb5SirEUTbN/X+JbqdQovRC65iTxWEaiIcenW0
UYSvYnaw/bxPQtIFCEzvFo54ZVry54G5lYXdKylyU9lJ//dikkd66ve8Qk5AESFqheMQwNRJYhf0
Vdeb7ycAk19GiiYu652bDYRUqx1l5AfGvXPg+J6m7x5O0c3gu3M2l1hv+RtImuD9oo85fpk6Hvo0
kUfkUu66XKpA3YYdOF1+/7MsRBxrrHBJw2cdcFaUzKGommuN4AAz50Rh3+A/w/SBZIjNxYmJvyh3
ktMoXKBdw85Y5DkAogwYb6m/bVL8SYJ4eBI4tVMjc0PNOUwPRxj8XnCU0uU7iknhCB5hAErxPiuZ
nyoTGYhutaj+0KiJVvx9h22EX6iC73Lv5GK7CJry8pwTLEk3vGuPmnCJglN4sGOwEGdtYy5nx+7u
K9OrhpU/kKl4j2brxVPy+Z+aAWQj3zbbs6ExD9a2zdwqlUwCv4BxeI+5Y2dR8Gzyf7cxDVZdh1EP
hJbW+DurEL4+lrZmFEBJ8rlwqMVNPWL53SXC1bpwNm0Ssy4pIk5mQ5RNrKA8n6Gt7L+9w97Et8AJ
pZuFGYpMx8vfcL3NLGTV+O3qlY6XBqR6QzZ3DjQcrVebll+6bdE4tLNKPgMKDzGaI2tgWFtsKLdR
acg2LPuEVwiL3v0tfk8aiDwApjfWHeHKE6WSI9Z2is+j7wb4LJMgUtPYZ2buMp3ektYwa+03AtHh
m9DkWoPg9unhZMLuRD3bBG9lMMfrHu3ZEkt2frJjxt3pXlVfRqXXXGdQaDA/Z0nO9RUL8k8hNxXf
LkK3DyON0WBYXkSq+NTWVFoPIMPlILxrnBMqamSK4gzQmfRj2z1uzWjF/pbR8459YYyJzTgkPnYv
+txfK/T7S2LqCnbtF+kfz4SMJ/OFT6sr4LAWUDOvx9uT0Il4BNcOYDrukFH4knvyZzShJ6a8xSTt
+erZklJC7CmTnR6dz7J/0EFt0X8cbYluQNYQK/zpBoKNIxLE8ehqdQIqb9W+K60I/YYtafFWXxDX
KWV96FeRMK3tnue2hSq3jj76F4rKBi00VpmtRpusUQ2/TX+J+tme37Gb+2QoOYh48F/iyu71M0b9
0BJTS6UQ8UFjr/iyTCsrCj+WBpHZZQ2QsgTmUngFARd58guOKD0r0T0gs0L6kpnvGvf5de8TUnXc
3LTyaPDvgVfv1Ktty09ROFgAUlXXVvoxThuh2Bm88JCKIGelDKnhMnbvqO1Fqcxt1GJuPrC308kp
/ml9BldeIUBDE3bKgGuaUBIGKcZLVLvZPnXfwaKbsks6csfHlGQMdzX5Y528g3Fl5Ko0yOVHRNTt
6FrOHxO5MnCnoQ4ZYn2tGJYSNOf+vG+jFEPGkoo7+TCQnNcwngV7xGGWYF2QhrCT+mAZZGRGCdoR
BEfBengOkkGMsJUfAp0eO+tqoHnjryXdG3lebvD/EfJZjno1FXmK+XryTFq/D3K+RQjGI0A7y7Pg
9FwNnHMPgXB0Jn/8Zvz5bdvBKgQDsC/vBDpS4FJGqMyVeB6FJyHAzucI8waoAYFG4ChEJMSoCKyM
QozcwR2C+cjRnYILlyJpAGvDA8n60WI1CS0Jyjx2HzPJYtv0XjImmpYP7V/bG8ZtuKOqH9h743/v
Pt6mD87oPpk0HUoji8dhTdyQqJ4dUMT22Zpub35IsBHT6rUug3+rll67l0Q/gAiyZ2Kqt18AS1Hd
CiiyC2BFISlwcw+XW+5SOWcW03xxTSNnqkFroIz2xkAp40ztY/W2G36kx8S026LwRWdMdkUmhAKx
EmJMHTlviVfzkWlAp0G8Y+s+PIyn6TQh84qx+Cax1ASXaxANVWxBbdxVXViQdLIb3eKAuoOtAzEk
QW1V3mb544P/9JqDC2Oye3BMdBcE2pjyPs1EKzJuXBgiBYZ5BWiP22wxw+lkMLqSRWd6Q8k9sYzT
HeObHuvGY2KV7Dr9rC6K7ffUAv5C+hZEfn0al0NafgUiAR0ZWks7avr51M+lsB15zXfwYqVT5Z+P
TZpQ8Rct+guPz03VCLX6CFAzRS9r8xiuwPeE/L3a2pP2Zh+VhmBihwap1F5V1RA99Iy5QsUcnhHv
SSd3m76VZuuunSd6TuStSes7gHWFVtwpeYlrbA7kDPyt8rJXGT9TtOi3hNQ1JSuulQWXrvf0Toqn
/CngtKbK77vXUwrmQiTLC97vGFaikXmWX5lGKRy5EDI2LHctqg57YAqzvN6sGI4RFnKQPrOG+WbI
Y3BzCth7xtShi9v6RoL/YSz9C/LFDpOASAmg/w+mI/NDcvDIekDbjSnOi8QSEaYJ5h1dO9S+895g
WECyDmZIqdDQ2uXxcu4jgmH5oHj7Nlqg2JARjxxgDP9bUOD7vRkn5Y4gYKQEW3ryZ+ZC7aq7dAHT
D+5QaF3HCQk4lmPDMNbirQMckKN6Moerlp7hkNJG33nDGioeiqs3NctLXFXKl/vWILTODdGBuljw
a8hHjvdjXmHgoN7E458NFAC54rSWb4Kp82OE7mCQ8MJ9a6qWPfFmIg50M+NszCFCoGLmpOHYeUMh
CE68nXX0ja5uVt3w72jdgbRS9AKKS21B0VFx941btltIa3emWh8oP5VRm0z2BjPc26OSujyhH7ll
PWV0hw21p0HyL2FRfJN6aRnRuqiJ2tQPXl0CDbe5lynbdrdSeq3tv0tEtKaMEnKXOJOHoSPhDATD
ZKY=
`pragma protect end_protected
