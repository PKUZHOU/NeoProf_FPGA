// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
aSIUwlVFpR2c+WKgJ7+U1Opbnh8qbB0Fd35DM0G/MtBoiNt+aDNrCZ6If9Rj
E402ff5LhGADNN1tDzmCJqpxpX9/Xushq2ot0VlJ9ctUDSGKrGg8aqPkw5Zl
/g+g4YprwWcB/80ceZxBJkxuPE2pZkuOvhm4I3iIy5gIwHxdsW6EzOv9xU65
IlyRGZpFY6HQ6qxDRNpLuVwwT2ALVENeEB3lf7DFMofPxlykUTZDmZdagW64
MdpV/YyEPD0EqT3+yFzeDntARzzmobsbF0Qzbt9v96siIdYQQe0COPQFPWcG
5VAabVZw6ZvwReChm/pZt8l8Mf+aCYXWrh7qkkCmUA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Q7w3UCjQCQ0XbTC90kCNs3wApOl9Z9RLI1KWz/GH960Scz1ts6BkhXyM1tPt
cHplMHH+n9lkE9KHd8M+i07NxQW7N9D/vaFWAMF2NNkEsLFzdNZlCto/z4oM
YqBvZSxpAlUtTdE8E95bXeWAQpnn5x+f3aAW5n8Py34zNgMwe0uHcCNrTLPH
1CvpT24687skUvlHQ6F+qJ2s7QIoRSG3nPZb0C4weWkL+rT99e1Bb+0pu0za
P/G3YIlLT/TjP4zbRfWlmrHLjLkHdanoH0kUYLHvmdtU3xMXn92SzUx4SWW4
maA0UZUxp/+F1ySgAQ5InxXXXsJ050xssOW+HsTlrg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
GDEBa8/0N8G3i1EPLCiyT2rA8zkLVpUSs7IOXGQd0lFoveaZ8JylCt2gKixm
OZX0c2bY83uHBpLLTfQlbz5cg7yDxLJ1vTQcCBkwbmpiHTq5YpHxXKV8DodX
VuDkLH2intMEJWjOdMrXKr2akYKcCe1BtrCkhVbqLvvZiHhFRME9fA2WT1g6
CDSjvFIquJhSuQfVg6wfqy1V/pzikKmyXmYWUealh5uAW5dGNi1GqU7a2VTN
ifOK90EPICVNOl7GZDtmr3nwswU4C+zNv1TbLLkxlzmr//rd8gj2WMXdESiO
P2ZB8ZlGpSb7iEgkDCC4xpHxC6YFZH7pnz1rXmYWog==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
K3QLgkDWC70C08eV1lLL/ubFvip4dX8AGAONWrKfN6nJCCZ+W/rdV2HRqfLk
ih2y/8Ye0tutJiZ78rt+4dLvSEWq92Lup3dXPtb0daY0GGDy1KQgUUNwZmuT
PtBPOlAxbYhYYZ3xsnT5exgmK5sUOOf1PmK+dCK0wz7uENn8dUI=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
TNad8KRDgn8e8QJLgg2gCCa6bodhFI3VQgAilpAJmL+VPrHVmLPR8dkYXZKc
hEXjYC4nmKdBNDP7RoyVh2jKppTxsrrtldiQYT7bvauNXjrnVOB39iPIDShG
YiNFoH1xLc8TXy2IKwV+JHTntXJEgnd9+IlbR/w+J4efecqn00zWFAE/cOLi
dUtzhEn1PFvkcARfJdzuVpVV84R5y7DJXCOURDm/YDse5SJlbXHDLVIeydQc
yLZ0dOofd+XIDp2LAuq/OvWEexAtZSaICVQUbs4caImLUWWkvC1gcqk07X7x
BErAOb3IJ7vNX9MnNSOiMCxVRfucr2xlnjM/xcZWE5Ht32ZkMJTiiX8vdCmy
VhXr/55YApaqGDqLs1kCOWYR1h+7siCTFZ3SIwf1j5Eh4eVek70hetN/cq12
n+50AA2uDrYfJ/DKTcebbTNEX5b/Id78FVSVXcDtzX+RIXfwbp7ClN1+15hq
sPHwRGt1WBzha/dfwXEchyu9cljiBKem


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
NV+wSiXOQ61ihX7hQCi9+c97Pz/GPEBY21rQJEyGCtVXJjf/rtfnULJ5r7Y3
SzGrbiUZMRRkCBC/mdaHhni6cck8dvb9JmkN/ajfb+TV9hfjMtflVaeWd9+U
YGtnxC+X6syPEeCoAwOKxBs4i1CPOBRSzNEeLEdOWzZJ3X54Nyw=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
RUsZEQqOO6vQhtRZ6FdAWUMqptjEfDkgc9l8SGSm7hQYYn5zNXlkHiRCRxT7
9oy5DlEZhmgffduaM9rfJhC5tY00e0IKMyllJOZ475zeTLZ5dhBFoF/wxqbH
AyTtUMAZHi5rmuLKxaBeLYy3vv53v6BjbD2WUabj5bsp8P+I4n4=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 6800)
`pragma protect data_block
aWSBZ8dPkgFRfUhBPLkw3rof0RobctlZ1XBpcuWucb4tze83KSKopC+3BuLo
Chx2u/J8aTA21tpt9fnp7AfI9vZa6wSlV9qgyEabJQ0bwwG+a6cH/QkP9hVC
ubiabQn6PM/CejT00B8+9fnean0/tr9DfAFuxd68VoSF+pAPXKGx+XH2FHLV
I5cOzyo3TMa/h29Q2ixj2PkdZSCtHBNPT7p9Ls7MEZ1ZWUwtkURXqOGNyiXY
/65NFvff+XBdSl8M8FasqpmB2AVE1/6Hb4JegfsEGdKyCaCVeSJjYl3Ib8V+
9+MULh83AGfZxaRGp/f+Q8uqFP0bXzTFLB2IDqRaJ6QMb+EFYRDtqrnFeDxM
3ipGOpGpojuqUKROIdp5vr9GRJEkh0q4319o0G3GErbMy7PR2WdNH+uyBbjy
hFzHt8OFER+CYGGcevZIWHBUyc8198Jr/2CEWs5YfxikqoBNQVUkVAznq6xP
uIv+MbmVJp4w1UgG4n1doizeVd228rXHM0DNW8Q7yy9M0h6b8DvulnzzDetq
tgpxfqaPcxMcCDL9dCpAe3uXpZOhuVVVzjsHs5tTPumfJWao+cdPNEdnMT5Y
M6DxU3XQ2uZE7FqEvwdbZCE3SquUrMvYcEILTf5wywVHLwjkRyokaF5PhWwy
y2MFN91K+S17urWXA0Q7mo4EdvJRm81AixuYC/VSQ8dhOQDNft3eAGCAgkHv
/hHWkG0yTuBC+rw0hzZ/a3NpbyL+hTJhtm8BXj/JtphyW7dP6MiP8EWojEPO
ncvFJ99WyYt5qR4yUi/SMknp/yJjLfDVWUZfZLnqfB/xJuNM7KlkZcDtt02K
4pYzDH98HiGgPxlIHd/S2mUpatD2CXqiViS/W91V9hXwQuQF1bd1jUihi57B
tkqtPRdQoWy4UpclgSO4XFlOeTf1wgabyv6g7A63GQU3GpbKB8XId6Q++pcn
YOfVyTwnBo8ubK2MobQzFwW25PsG3rY1vDfw8Jky+BbIy5bzOiytot2UX8WX
cEODMd+fgJ/znooTpY/Mw1taqmJfMyQp2vUteWP18HNhfHka1618hN/X8mX4
CLAEkDtfkmbDjM68hiNwSb32woXqTYYWfhIGwudDmp5cWSvoa08Vt+T/BRcl
aPO8/X65upHwt9Cg7HTAX+w6CV69XfQRiHn5lAhgMDjXSzCJplD/fnY80uvO
3ssHGDgF+0x9qE1iXkXYRbeyxvyE71tCMgTARRj4mtE6FgM//Dc0Bmc+1vZx
Lx6SocS3lsqrjDy1rKUcHbYhg7aqw165V+9HrsfHy979tIgsJStQfvmc9goW
6nhaNEPaTBtrNxWaDrpgoTELJARDTIg9QlhS3ktN90gzGlWt/pqjl5b2NI/W
jf4f3Ssaz3GBZ/6nALEn7DT3IziaL1Qo9jeLhCDWsKFy27EwEVAoN3dJtatR
LTIC7mhynU3oc3RHZ7XyvgtO305E6TDYNLjdMLFrh23UL6j6dZKKDOqhNyhk
Eif8dX2aYtXE9zgmLMK1xn4EZNllXvMJzyJLCBNE+BorwhUKOQDVZ3DHGvcM
pSBbklqYr0PD2HVwBWc3VtOqV5GCSgJTQXg1e4NBXycItae3Vp0DJFTTfWOc
S726qghDk3Hx1Zol0jvv+NIfmXIhcBt/Dk/q9D7amXRfRmTGOpJFtFSPwykk
WCH1pB6Q/PFWJdNE7i9csFshZrqb1bFPMxFcvDyMXI8jtL1FTT2LNt0q7fVS
VZ9l1h5V/A+5J0oU4dnHzDquL2jNkkUfh4znFysZpvSosxOPMZacmu0S41L3
S6yaEAiXV6kSTSZ8I4b/RsTdOHl2QLSZ0pCHrD/2vwgDDBHLgsC7ZAW0brl0
Ic03SH9DBl1meAtos0lcyDVREeh/RVICoqI0BA5Ap7BiiApNSvmA+aVWH5fl
GGKPV1RWzPZJlEMrFPAhLTziYpt9M6X5eRypL3awMFwrGpXvQ+AoSaTAjTjd
avNdPMXYk1fmyojZYYc4WkoUIuNsnd0iaa66kb/xAY8j6+zt73zvb0mmG3ij
tBLndKW1ZU1lYqzr++WWvZk8YumSUN4rxbi7iRVyXb5nlF78Sq19jHvwuNos
qKlDEQk0t++iqC951dRXIcYbaiCjJzSMrMBj7HB3waCdyucY0N+jVv0tqFu7
40vs3R/yKOMo2RltbolVdL/E6smBZ71vSbmP7cxZgfu43ZvKF3f049dJZ6Q3
k7DExr2+WY9yW7lVmSrGpJRfFd6u4ZznMVX870cHH74sktxX+USgIFpZRqUB
VIC/yFMlHYqa3E3xzxaz0KPNDR4NReptyOofz9WgWexQC8dmwwyjHyKL05NQ
gC6yr12PAsuwfQg0kykq6mMvE7S3uig5XrKAEc2loKFvLGc8G9Z2ntOmLHa1
OGGLKyeQ88aqEGEv0oQeErtQZKphIubdOeK17RubbhNAJBdqkllHuAcwvJ2L
L4U9PotoNjLc2cqx1hvv9BTLvJq+MpU6H5fJOCCisYBf6p5eWIj/u6cLbSAm
18EVPY/fm+R3yJCHeMc1cDshUTTL6/cHT+EVGL54m/4AcBf5MNo7cbXHOi1n
WJUeEXvtdGjSNJH+KXfWi2zkfiAdBub9B4lPr4ycL0H60tDP34TqBc+CRocl
/Q1Lsoe3z24HuyjaitsZyCJFSzW35h8kHizx1xQPHAO1kybkRe6f2REf2hMM
uXea/VRW+PZHWqHrF6JA3oZDBt346xr1FKp3205o/KJKIN4Mvsh5SsC++a3E
EAruZjbti5xedcQhlNw3XYC2UWZNMHXGiNWfsQcdUOmbcqeIJtlnMHrGRJEg
PpiF9QGySyuYlCTWbr3f0V2y7nSEka+ERezQJQIW6SSoiqPSbeu9KOO1ZSwx
hHWAhgFpWqz6ZVpgqQFC+lAj7xTnmTGOJ8J5OTz7amJaLKURzDxaS1ihlEL4
X7bBrXHRbI9fug9WSyeBRl+OkhID/KQEbaBLtYriV9O7Pxh86Nl0wCFq2VPz
hptfKtv1duUz1RFMYrJXbSDtcDdRPSx12XeHwkDsdHPW5U55ADVXEPZH6UH0
lUidNK6gxLDb8w3R5a+2Dln2fl6Yo1I1JwQxvApJWlg3EVrmfOLZXmB14jLT
0GwmK+9XKDlQ8eTQehIfSN1ED7UbKXdveCY36PGQ2/1l3ihrD+xbrigulCjM
Uhy03kjwxQ8P/gsuxcWllt8TTxCv46HpVpK4PU+c0hJc+YhFxQtM99IbFnmF
5ECoNbGPICjW2zt/XruzTcG6qnoVFJs0Xe0BE1uBgOxK+2z8ymdvsymyq6t2
STsmQxVMcQtqVcm4qfQ+oCCBMPi3VW19+72EQMOWRj708HGzcjDEADJ9FMhY
8Q/I21bQSUQH4TfuClzTb8ProuphaqNBfnVaF1QpWI+I9Wo8QWg7NiyZtmEn
viGd3ITKybXrm1P2tcFY8OR9pqAKDjrzXniSXDl4bvaEHQFgsbG1GRtAsEDp
ETcmDJ3iftmHwjqNymoOpooChrNsD4KuEr4FjD27JGchIMN5B0dtJhpArbHb
0b0zi9+OW/QrTZPBNtciGyykufPRMvfHH4PG2g7JGaPuYgSLka5Eym+JgwdA
56uwzXvHp71QCULHYhwhrauHckDcu/U1yl8kEa7Ye3uPOv2q47c7VQ/Goy0U
NUDh1wbvslBJgtFUu1uLZRywhVN3GztvrxCna/K+O95cMRbk/awY+LZtI2Qy
Nx6P/IuaqzkYGX5dAaOi5Lm18j7AVWoDRqFc54hq1ysasSj8RbXCXWHaxeiy
Ie9tXsv/KMGaRCoY2Bjf7pkdI0NCsiP221ytm4f1ggZs5Q4CdMRav1EpFiKq
xZ2hiGbIDUjt8K2Zq23wUUBk06nQXVTsNjmSe07d96iX0/gBIk9Ek3rO03g2
m6I4I0bWLoUyeAkjQCZ1cpSc8+CQ8DGRnNtjlIuIYT38kgu8iruQ3y818RAS
1SWCutsga9gcbPe8IJwH/UxL9zgXF9QWgTD/86WKl9NxHPA6+sxnSGsIPyFy
mParBJyJE1UYVj5G25XD1WdhrPWeS4BpVSKVYUrhqgGLLILRAkAkPpM90DBV
eRA0GUymGEf4oNz5rw8YoGLG3sPyh6iyhROdAVHwkOwUE+D8iFzYl8PRnEut
1PMVfinaUwvjI8LhIrSSNjRvpIh1NBBvbYdSaxThvr2NwG5aEm+D3QGs///U
3YMpVHAzezc1dm1I4zJQ8VnyPxKwdSZS26eyDtaupIaoCbi4C+6EwXcOX42h
CHbJ7beV0NW9wYZw9BhmANsPDC1iB8pTpRlIJsE6VPtJOIPkcbsLi1nd8qes
ZO252XniIflrmMN6c+fbNqbsyIcWkWmcoD1CT1qZqrbOuAwGB32ft35bDtrh
s4RYHzVbSjq4vaKAkTMgn3rW4tkzR0/4m/YC3r28okodFAts1M9s12pmXaVz
V/SeFKaiTpOOSMV33QD51L6xzYckOOd8eO4pgLQC6+xF+tL32FB09+8h3rvZ
5G3xlevzH8C6bhHN5DwhXhCYIDuN15GOffE1AuMv8O8y5OluQMSwhwrlLK+q
0S/5o3+gfeCUJKDYZxnaoITApOVIUGIyhLUHM2Lf6AL7ftjgHTO/dZwvmJ15
mMnCU1OXoSoHsKR/rhrzhsothOsIhxmWnc84f8pdkCT/4Kt7XHoMfz+Uz8sW
+kB0rKERKIyfSUO0DKIkvPCPMWkLGFZ3QnEkYCjLCm6JVEiLAYcVzl658wM9
XmTG9zqUmN3l6FsvUUVnLdTMWvUmCcKzXzMZYAgPrCVMBL3nSnNARxoHHNp6
d0nv2TBUn0yvAyeTzhgWYuxcWQ6V2nS//IgIpr+CtOnGxHNvSIvfVo3KdTPU
1E/LVUuEEmmrvIL29zr5IQdh6kOdXctqYKgVkz4AtJghQaL1FMWEgYGv3k8h
ia6XDS1auFafvuA+ib2JDQG4NF6D9J1DrjVbalsggxsolNUOW+B5/IlN2z+f
TZcbvcYYv++9ZoHczu8cZnhE3HqQE0DW6CldKxTGjGKa25vFVd4hdTIq2b6v
cFRYUs+2Q9DLHhSsUSnOPJ5W/6STQr9q33v7/d3lySYPHfA1ZtEhNwyiuTPj
a4xYdCAzwxZxI7Msd2Y7gv4R7IcG0I9FqRxwtm26P8x7STE5bfIcIWT9EjtC
GAufRK6ZRRaLQ2WQIzjTwW7rXtnCt26arO4bMHJtwTFbl6xYD3swhfSH3p+8
URoYLKgkDYkk7ec7Wine8s5/HvXbHSbJUndM6OMKAOtrRQE8z02+akow//Rq
PX00MFvBH50AZgubhrHg6OYvXfAMCgRHh+Fv1XrUX3jzGlYVmdMWTGhsLgWO
ATSFP88hQ2Xl8xbSASe/ar98+AaBdjTDdQqSx0eL/PNAIEEMPE1wMfrGsJ9r
D7JraSQzWxpgwkGDszG7Rh/cU7x+pbB69rATctAHxefwb0y4cq/rGn9vWVbp
hIb7kzFtpChf0HONAGcS/aZztXS83RQUJtU97KfigvrvapPJ3hTPTZ+8JZKm
/YlOtu3gIp+BdW9T3zgx/aNiY6ARG/iID3xHz1jL1GHqCwEo77SanHf1LML/
iLlvUCeaF15lEayS2bA826Zs//2iLC6RiYYNxz03o0jzfoWR7HxOm9oXibcI
LFh/jZwiaGbQk+H5+UovZjAgabltPt23rZMqOW8fRXfnqT6Pt2n+iW5NkKJ/
YsIYgdjLx6U9FSil82Y96HqJA3z1/wVzCrOrkN1L6KdrwVEKTSa+eV0sW776
nLeoSbdH5bMTtbAWUzw0HDiYj8C7b8h5/V5TzqyroT/9njEffRXqDCvWGZbJ
DmozHsWekgBdq3FiNGL3YU9OUpXuwxyvTROjwYWybtFX2c/x5y9MO8s79WPV
nlr8124c/8GlceHxIQwANv62UFJhBKWFYh2Rx2Aq5BsoaEHNqkVetQUXEBSO
x6Ti09RalCYr0Bj7UMFJ+KLSc1rKbOTW3LVzaoIlJU0YbLWOMW50X+zti1My
DFB55ShauYOuaZtrdanWTlbByjD4Vhd2PO52Rukfi1JgG3p+sxbVFKYKCsgx
/yjnIOGWzGhaamjRkA0tpeEYTHx5qkHEBdH26S9VoiOYyCsBA7e8QWecush9
qrRzo2jL7QAYSmtlflHp3qhxqhvtBOUGrkNOl0QHqftRWuIXltxAc3Tm42jn
9wWrBhei2elXMAy8wE5kW4tLD5HiKwVJzPqiQbllQuwGS24AHPc8V/o3eat3
ptrx1nkKB/aH00w+sBLPN56jciTazb0tZL03jIb+dInQM+psaShyGB72wzRb
SfK843ocNxm+H87HKdCkax+uJqdKCdIMZjou0iNOn7jgtT8cUUvSJ2sfWJ5W
BU+wc4o7nC8xe8o6R3OonFxZz/8MpXAPWomsw4tqO+1qrodXYI//hBIc6ajv
nD47tW7e+Mi1Y3eF+74WdAUjaPeGk4CANixK4Lp2/Zo6oDoAcqqxAOCNk6JQ
5WNKIPtemz2nSxKuGC4EFcqdguk28u8QDXqvn/n6whZksuuy4AGZ+nSQMDSC
GRUIAtxr8Rm8AXFZwDsx8jndzE1g28xPKyaK/UiZziZaoyjNHZdPZ5Nsa6bL
HDi9lgQLENNtb0WngLeK1z2SHona/Ok/Oih4jQQYDLLwPomV4diOctawUKmL
HPLyfGFgTzWv4qvI/qnvA2/oenSdNdDtr6WRw2yjEINV/jAAhxW35i0mk8SE
YPszJeyfBklfClpFpPkbGs+nrJnBWuIDks5RMN8Z0PaiEuqZykDM+jy9wC8Q
IG1VyRCeJ2DYb5f/wrSJP/C79QQs53DIwLh2UszTGc/T5CRbFn2nLq9nYEiT
mTkx/nF/dqiUaTiUOyPOuM2YB2KNQMu/d39cWNj2pJ5LVPsYgulrnCUO1o2v
YNcC8BXQ+vASsC+qvpw0c2sS3tFqg7dLW+X9yKtGRJNrm8cBSb8Hy1kJ/SCu
Hqaqij/GgK3nucIZrD/19A+oXEmB+WnAAEPEgsWGj9DtH9mAOcMZ03gAO9UK
lnKCjKx4SWjZsPqbuhfPu6Wi/JQsyqJ2/gt0TvvJccN8FulKXFY0X25uX0ja
/D/hNMn6lT+XLsUUo9cUp+TnoO55TbpI5kutXrTgLFN8g5Da+4jlzCyq7Lf2
19wG8VEATKzNMQDZnLFQ+FxZbjPhDlQUnO3HH0Qng23aOwUf1V4aJgezBinR
53PBWTyqCG4ScWvrrDmGJyrg/+vQ5gpqNfXjsbFGneVxrIES9x95RiR0ORF5
8ai5knBm6fxJqntxvSFECObg+CbVF4/1MaTD04dM6rPtbLErOgnEFCWLXklA
u5KsExR35dlcNoW0asOCZYlujYOO1kLStUhJXElVbdvwXoTCoPb2jO9f7NHa
LDgDKaxpJ35/a85Yh1pmIjkNJk6bVndYP1q60d8MLrxYbEBcv7AhtFmfk1GG
5FiyWX7Gy5u2yubXhgao0rtTMr1nqrad6Yoq+WQzvtZeYe9N7kDmjr8XNYSY
AXvJ1EDtycuYWfKXGO2exbCtrwgdyDdJ4+uveJBz4d17bcB4A58YmV12oBuC
2YUvWb58bubS6L7974IzRMNRL5SECDfHWgyI0yBti9BCfsbOPuLcuIJhi7Vl
TfOaqCwgIBxbEEpZjyRS9PcUPOPDeHUqLWzjoT7fbGUyw3QaJKQVnN7hO+JM
soXoJ+mQ+XxZYGz5zCksu6Pz6oWPozotyu7iYNCFFLnHT8pzZpCXvThP15cu
emGUqpopoqvpZH1r1gObpOAkHg3BMpCfURF9RCUAizXypF1FBV6boWZVaHWI
+UW3KTltujnJe4en518We3HZzH699s5Jz2blzHqq2RcWcLHjRk9m/g0nQHbg
lBOwd6mLwnB0798gOWKtdhCgz6OcMUx+1cHlip6Vyrn4TiB97KexdWP5u3Gs
E9sGw4drh06XU6zcj3iVNc+k6XrpGCvThzuZzioGaejaxnDZwTS9bGfmJIcZ
2Yq8nhTx53neqMJNjgTl98n1QI2Eyu66KY0uhUhALHXnOcMx183IQnmbdWDn
euw+rv3q0CV749pXSmrESXILVeMsQSD9Y/UEBkJ0K4Ad3+47cqsqZ9dUcsuQ
g/p0ZmdNWN3eQjDz+RatRRp8+9WqX8bWMCPS3X8VkLwZCketKxGnpfSmbe8L
4oITN/fcyETKfUg9bB4m5rp4z2wi2LMN8TQoNAVufHWt98SUfdWsOrc8p94z
6rhb9viSEIc+Il/Cg7hUU1F+D6cQNIZsFaEXoMDg8rvn52dDkFAHJcVtO3HR
0Jyd26zamYSUvMIBFq0Ei99w0nFGCrIk9x9j6xECPUxcQXfWEQ8WPc5ro8Zg
eFPEYN3bQGNkjoZXGoCYm+BtHiC9m1ACpyj2SxWba0TCv10/+Or1MWmHOoOT
kSJ1ogsgxVKVu0F6LqjPKagtGsdy3um6SJ2PRiQe4QAtpyb4bO8EtA1+dzCs
Ug4hb4XysaK3P0hE2wywU/M7nR/lro3xpxnuh3AhzVqj9DeKJW08zYK7Bkon
sdaRI35SYwcrWWhK2ccHyIEwYSntQ4rdt7fcV9OqJNfeLV++JsBcN2YKtq3z
YgpqIs1SK5ZAM4NgywS7MHTNBlwkWLRJRLHsA8fntg4JC/+hHepaPa0uDonk
eGhHxYzqBBsm7lYMXguNz1/4Z1Hj1q2bxT9x8AgMxIUXRxIJD+2khzimfqvW
1H8B2OJAoSBwf8ez2gTH9zt5IMqm1NyndsulgKvzcIX5XX1RBiqqur9/TwWc
43ozJ0TCWbVedTpcVzkuT2YK8ZlkTDMzdCt92aikxqxoIHKCu8WVuQZXHnzJ
mDCm8xOxfc129cjldE2yOO+Y8BlldytwJ8NaiNzBJ0GMVAQ4I8udK70u8Rse
Gl/FE7d3MsVm0VBdoDDs7g4+sIIALESomzuitLKJx/UAzWvHDQG1FsYmtN+l
a0N5y+l1KsvuyaJNcdFOOScbtqQtsxTeRj8ct1utv3xxZxyVflCPoGqIbaJt
oTq8+2+aevmKCovw+YDjWha5IRcm8DkFxhdkPKkL2nF7VZD6aRZHzteMFP6j
2Tgfg54=

`pragma protect end_protected
