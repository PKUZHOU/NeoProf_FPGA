// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
kX3e9yEqc8GEJ3+jJkkTxbEO7QD88HmsTQ3cI0HQ02UI5JfKE13gDogcK10a
CUc8mbJu4sf04ALKcuEYehgNkHRMxBNT/RanYfph2uLm+Hs5ZyqnnIXc2lbv
BYCbN7dBozn/ztjCSdD/IPAZoQFY77jze2KKXTZE++8p/oDZZJgfpYUGQz+E
QV4eDUXq0VHhKKBNME10vSUe+sb9IUSkGUC5ZndN3DLp+mKKmRgqh5pbZaNL
gXqve4buIo74+UNXlf/ubqPyMvOJgJCbUERgN/2mHD61gKhVbsCDX3umXGm+
moG0Zr2ucwvjkHr7DcaUrHlL0lJeuZpZOpbhJPm5GQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
JwrEQooICzkIa//8HEnhIFbX8rDAJtKeT35hiErEIUnY1P0y9FP2tZW1I0xo
kO6VHAEpnLJzusux7NTkFYJdalLvCV9ik4z80dZlOC7ohu/aM7m+D5c1ZXC9
JK/8exAIY2rTVsKwcJhKmucpUCmciiFIug4SoWwfDdpNRvWeyVQYVr3v43Hj
chJuQ0VaLvT8jwQeKJM6KP7QBZx0sv4E379C/gP7q9ohHdzm2NMe6bk+/M3E
KHMWvuw9cv4iCBOh8IojdKIuOuweqEmubbaGVOrah/ACDiZpHXWxn7oALk9+
6+36eOKMN6K9c1wWeF3fOFJAAuctr0Ujs2VPu9nbWg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ZRtT4uHTHUmrowiPJJr+jD30eAa+eg4zzgowH9e3m6WZauVbvkzw4Ty6kRJr
OVqkhUDfxwB2Dp3kJDFe2E6iudDj09fLSEWZwia9A7HlBgPDp+VsOspnCxQ+
nnNgW7k4GixlqWvjj2GzJIqJBA8RD375TP78uHXjyIio0b+yJS8GNpP9SK0R
U77wiQ+AS0UDRF5eT8TXQUooYOjUXFBgxxbvSGsPJtDdkJIqTzRUBtMuMPzh
TdlP2z73Iz+AZ1YhmgnYMzooimGkDanu5QSBdpkeYbDu5mPaIQyuhIwUPNE9
LNjUoU0winQ9xHYkhOG+OYpS4r/qwJqjBXE+NKKpDQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Y+OgCsuny7GTFmGrZrrc9PzCdRpV+qcAPtnBsqJyTikyaqaOU7hOmN4zHPz0
0cbmtCQHlduGJKXFBpBp/BTwpxsZSJpJS1mjZfuNl+FacYXct5LDRwy497Wc
r8Sqwb7TEtY6VU3psUunbZCfE/bM2QeptZTEMZqeeW3FioPc/UA=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
ptR7w7aFPLRfGwIrmu6dYtxhfFmMRvKHVWmy+PUeINGZ5+w4hKFAmyLy+NlR
ziHlOzFHltLTk3HS++Eaq9IfLRIs4wIum/eGiBvC0k7AZcbY/OFtxGGHCf+v
gQ//HEXYQZl6Un7vzoM8K4myi+COaI2Iwa4KPPpgZIHav3skHHCK77BJbTU4
JvBje9ffmPTFi8snj+AK4LxaBpPQbd4J/G6T6d+bBwK0c0jjxHWQawzySbtK
0SnRZKEw88y1Gd64utrb5xvJa/+SlwztV2UniGDlKCFspv6oh06lTf3qG+7a
uQNCbPw/e+TfMREi5nd0TIOmFKPrVpzDBLUxxSzjPO+5xKfNM/XyhIysO9Kl
S0W8w8UsteuAjIyAH2T6TiihWZaakP7noFghtzNccmjqx06+WfIt0CDvmcJU
WoppxvRxgLjP6Fm6fbhK6JjTFmCY9b01f1XCL9fCAMrr9z6LbNP/slWaatYo
j3vllbU9b+FQ/6Y9VOS7eAU6LUXBbYI5


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
rhFC1Fm3djDwjs2k1POlbFxa6RpKyeXyNw0TQYRnHthn4fGtaG2hfhIEgOVv
7Y97Z05MAs2PtPYDrfx7x6PNgGtH1ZcfKApAm3xQT6k06ukeikbNmspDZP1g
u8kZZHPzNydWiuFZH+ZRzUqaRXHjmqu+2i6YxDWcZF043f9/Bps=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
VfMd8FgJDkyB0JsduLlUt0EvOULWO0byrnD7prbh009TUfaOxyv/vgqKtGh1
MklGFmNqnqb+L9RAlojNOOSIyxG8Ntcih4RuuyVskQ6+wRX7DIZ0XSmFT9wv
gNsVSxIOIdQ2EQO1BvIA8XHXabiWopHYVU+uGbNeb3e725ujEA8=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 57312)
`pragma protect data_block
JWc5u+z+D9KlkOMftzx9jGbogar/7HHzRCHqBnlGIpzOQN9hYQmaOIWRJDc/
MCjqvmNGrcKRbTW+ZFJzQQPlzYCHXdnQTHvGoxi+RapaBY8l3uls73mUJpWZ
zgz4Oq6V7T2H8y1r3r5d8RT1Mq9OjvmgJB2n17DTYbEb+4qforfOrKm4CoPg
0AnqsoKSvCuUgOeARuVubvvh11VvESDKvAlwx68w2tjXeSnB9rwJ6ziSinhO
piWwWmFHo/WZLU7wEw5tJ5pVLFqXe+Wr82ZNX6Jl5dizfXs7x5eM8PJetTvy
VbptuHhbU4en7NLB/erRw3UykIgkKbg4qBBj7ecsbUhpfByt4yZImaJUDMEy
vnAmcTgEuFmTlHqkaM9g+44+Iz97j2l9GXcJLxX0alaGFOXVALCwxtniEvmN
7/1qaiFKLbm+BaGUlKF3kHkq12/V4rRXz5u5s7DS9p7NpAHb28p8HHC/oyVH
uE7PmXu6lyAW/rPdYm4fh3BI3SH3AuXIWhaOLdV55FKSTlkKI4+OwcDUwe5w
+J73iOBDc0O7+NKxoUpoZQy5WIrm+yRMQ3K43LyGoV5S6ljBcKzahTmoZhj2
mb/ncn738QfOu8PPZ/48i0WrIMZGETis5AnR8QexCdhU3/Zu9EE+BZ6qVjGj
sR+km0SPs/E3qPhRB5IcZxskxW+4UFtp+3eK/P99AO910RiAMZr6PBQ/PI2i
KqWfHZRT3XHLnpwN9VYAKRzV3wI1b0DAkesEMQmNXhs9uizWn9xVq2MDpjo3
ZaY/gF6XKG+a8ZC5s6o9xW+hhSBULSwrz9kRzbUD2ggeMuUckBAlOtBQM8lB
w2jliVgd+by31SnI/12BT++g4AV5mv4Jl3lJxlmSYemK583vG7RYQtzgjuMv
F6A+1qmKzDASTrxsL0QnLc4oIGHPnmTjym/9pRca2XBGbqwMqGLi0GL6XLoD
cCzuSqNfDZsAMXRgS/1U0+GcIH6tOBxMzna1if9Hc/LVTG8rMUhClJXv5ht8
lb8Lpn4IV1X9gM6UDsmkbrLBIr8jCvFX0mprNGn6AtNz+C2O+AJj5cjfURuX
IGEubwHY+RW/cKOHXNNWAtUvWJIzFdYM6s8TOrbbdSkO3TUlQOWpqKuy+mHU
QvB6naxGAxDUGb92iEInE0M6Ax6bTWOAifCsguT7r7w3oE07zOgtcCTfu+nw
3EhPa7UBXske5tznPSFvbC9mFM4CzCB+7km4TMM4lYm24K8Xx4EH0pbHo5aW
rIMg/ukxlPySomwbbMTo64jlJRUwufyx4mHA0VJvEmQe+sIoTebA88tnjVU8
YbF2UrsUyq5ftCalL+K9BabFYiYDycToFatrNXVQYx7acWneg1bfLxb+nUea
4hLxOu9mUuFM32yA4hsPFbI6MekUPl/ikE7oeNDxN7VCVQENDW3so8KXvIWg
znq8TlAneVhtNuRxPH1y6//wDRz9wFTXIDzqiP4vb+UNYCfVlyOScwAdn1JH
sFGHwdrnGy9Ica6EUbtS5ZyNg8aVhzPXNlS+bu23F8GEwgEy/93YkBX50im2
LRNQs3J9WHgT1jDExhQKymjLV4VKqFrnCw8rbnegCewvmKRSNSnrvtPYoSj4
JwpjYxv/0DozwFUeN6qG5r+/samnQTrGz6PkPNVZi46hXUngvOn+tpw2rKnb
wVd4kS1EeQAVTPr0flEvY03DLHC7zbcLKae7ojwXOesV+fqy0z9Gnl4cI3eX
oB5xiAF/XfCz2OJjiw9bw/895U3jtMtFVkEU8BtT4NiIqWAhMWz5t4dcrnjm
AhsgtKfuScAv34RZfNmNaSV08b5cCvYwQRG89VAcDDCBo/WRqD5jNQ/VTd0H
qoiMxMoGqxf/GfC31iOz4ZablzKXeOb3+PH/plXdQBMW921nyuenEsGqGUBQ
DI55e0vqGgCJpX2T56OW7f8gBLuwjnD+RKvJ4XY7xpD1K1/h+h5ZZd7xBqii
RJfyUcgzyNEVpMZ54SSKEuewgnZ33ppviiveW0x5cztGs6N32RfdUYODWGgw
/UYQ+mc/pAdrA4ZQVaxrtmotPO9NWWEyDlue7ANJ78y6cbLsA++O7Sz6zgZd
3XL/MAzfSmd8brqXZ6KNTK7mjAwUjEyuOvhMDCRaFhmcUnCZN/onZ2om0VKs
+wma7a1WFOn1iZyaN6msBD4CgcP8xPGyE2XoUMglWUCtswtyV6Kk+s2tKRuQ
B6VLVusSZqhEbDczBztkt9opEzI+SL7ZvD6uskV7QvW4ZJcMlsfhofrNLtwv
XtSeCcDL6WPem93cC0owTacqy3AHn+qp1ODa+W2ulnTsdqnQWlPXBQmk2w8Y
YfZCejRiTa/g4gkfmLWwDRcog+S46EjqCu3yjwqAMLZF6qLXFqtJj6QabyFE
1WLUJ43nBJW1OPwAX3B70QHV03i7DHCxkyleaVa/5zzmPLQ06NfE4nIyu5T0
/GI+/OkDmc8aoy2B5YWkZhJ6+fLxCNbQk2NFvbBuL9TYmfXhiMreRuyOMkr/
8BtsWqD9+T36DIxjQl+sIOwEtLzkcO9irG2SwXq+LXPCJ6Y0Xiwh9HU1J1yt
kQcfThNlOHwazn+NEIVq8KTTofm3qShCUKQvw+F6yECq4Vlc2xhV5kKwbu9w
OVn5wBiDy9sQCx3l0xFJf/0Co3plqJ/gDAv6ZrqBYnqZecaIPdZTdehpb32n
0kX9RtyjrhVuhyeaUXGWJ+ahIiGLB4B8Ut4T8hT+lqw3B01cqDE7PAav6HWU
2buk3mdq/9JvsAEiLmQ6V5U0b29giHVTXCTKBbmBVQgbBaQJD0OtiOUKbS3h
2zF6HojStY1Pd+AfQq1eAYlHNJdvMheLNe1ehMHR9FtrOARm0rP4DLAyj7Pj
nGNqkjmi/fQnt1ITSoPOUFog0fE+QMEoH0vuwBt7MDKMisIbdBld3+wyvGax
FimHEuQIosG03rLpkqrZwSyegeszn0N1CIEQO8L3SFR/StTCqFzspFfNkB1a
Nh7WmWnclYlOnpPk750MbgHoi/IxbyrxMXP9hIIGLWmDCePDjlb8ucv8ddkK
vcXKzhbEjSIXh3eEL148vb0/Ib29kZIAvOWaZ9+z+sPXm+SZ3MESnVdnMZO7
srlQZlE0PoSG+snf5lxqgg3aSWtW3JAoVzkXnGY9mqx6gaxCLAm1LHA3LrNr
koocgUlY3ct7Fvp/o/bWtPdjMENc4Z/PDpBGeplQXc4aB1kzsbJsSP3nVHNj
0b9JnegrwBrfEwPx4zvSj269NtrglUZviJve6ieT0zoGazPfl6UqnBXc8QAW
tvf3Z8DcQvebIpCLIMWx7ibAJtHpWgwLtbC4U1K8UCmDp0FmzOmWm+rJR7NA
/oslKaYevziyNvH9bjQc1iDnIbIl/ZYof2qcbQ5Q0FyI1+BSjSwr6ro3luUj
FdwHpB7ArjHLqTJbgoCkVrYDAboSelJD9ubHEmOMaHCSXBbvcGDRHA67sQyt
5bq5WT6ZVQ1o6sBCTtkk5xH07EAKrq71RRj7hSBL4IVwM1XApKkfkXShy+mr
n/uA7TlSe35mAIYAGtB5CJVWLsZB45ncZsES5mWgOtWEaeXmDdU/bzacGeN2
5a4hjVxIJVErPdZpVRFo18ddgPSFRCEGxbEkN59mqG+6+XeW/bSMyFdJauuy
UkiQUh1oe6wG7KNlAXCA0Kt3bA0i08TIZVWsqSUmz7jUL0AA8LzZfvj2uzR1
cmw1KHl9YiISoK9AA//QIj5xpNShM07viB8K3yF/dU/Zd7S7onP6J+h7ktU+
0P8UbVH3b4NrRDpThVArCLvtpo1PuSYlOZssx6y4lPqu5rbXrC0t5vTTb3iw
3DB6rGrDt4fPV8pPVVQnEmSu/ArBQn7oNIDUtoDRxSquF5QMknaWa0jiYk7j
vKPFvRk31iAvDpQrKsJ0rDdrch3IQDW3SH870AMK0tP6cI1zaDl8O+4t0xL4
GtGxSp01XHlNkuE1KDSdb5UOk8nL4Kub6hw+k2P3i3L7orYsvKC6jil0sPki
p29fzE2pnD2Xf6IAQ1+oFGZDrc/J3smD/NcWW10W4kUMrpOd04vaegk+M8sm
cQYdqg7snPN4GxtAxAyTxMqcVlCdTd6pJdhMZJodF3ARTDtduT5URYwBcNGX
cv3EXZ9Dp5b9YYj1DQ8xblhIbAc4Vw2xGwnod4PuuNYyOOinVJ6UAsfxKJD4
b+4x6h1cmgbVvrimYTQ8RZ+Yf+2CQ3mJZaiNNKfAEbQ7OQY74VzkB83d3TUM
ohHE1oQqRpodrxSE9iowRrpQV6eYog/H4Np3sVBHTaHS1N4Ojg+X4l2i5eMi
VW2wxXE0WMXvw3GPP0qyhZYdpL18en6YqK56a9+40zvPjwf0HxYPsM6Z2Vpt
HSYJyBfTubnp2F034BrbRwSpQ/dST2ZEJrw4b2yHmliyvtH07LyvOvE3WDCy
+ITL3FlIYUXGmqQB8+tyxAETveUUpxA1pKTv5WI1/xjfGrxJLIej04QxA9np
6sEbdSKzq2Z2DRUlRd5AcBL6Hg5/H2hHr8Hy05Bt2s1n1ivyjfBzXUHbPp4W
UuLZmabVPa6GaTtt/5KUDfG5ixSBh45rxl0IuBf+HpmOHb8cOqkuXPc5IEYn
I171zPHSoFB7pDo/jwxjO16B/7un5wkrrFzpRjorpZViHL4spLpxaQbCqSyJ
xqfubx08ND73ixWSfP7ZcAX6esq1iK+y8hBeCAz8X1iSbRlp+3xIAR7zWcaD
i9O9t/beg0ncH8KZNnVH0TSQaFnZEgbnGajv0sg57f6mWU5z7kMtjnS8pxD8
5jEBNtnjyvrIyeqMOqacbAx2PdnBV+cVyKdD6jqX8ZzPoEK5L//IOmfdu2RY
cJ6R1e8P3oNAN9K4+lNC1rNh1fip5fxQER6mhVobE8HpWYwS4tmujwFD1Ow2
aLxgXzU+h5kqpRDqTV0kptQ6P3/tR7RFYd8OL1mTIs/BgDmyx+KX1Z7kS3c5
TooxOXZk90PFtZI3czMCOBXoW9Vv9ru5jL1BWnmQgB7bF865GVjzgI8RVeWP
IY0lV6P1kwc3Jk6paZMDwhlp1SplI3jqsfPyA+XsIs4tn2IaZPl22T/2Kp88
Ku0sRCPzlkjUtj7VjfGUZ1tpqQRp49zglwMad3XKTrvw24yCsPNnWDJh+ULr
zj89+11AlfTXO5S5pYr6cFFP1xEB27UD/rKxJH8JJ5NNZlsh8/524wp2d3v/
TVYOIaPMJW8hcOfOA9LcJ9AZRX3aeVgv1/ME0uRW0/hbQX3fFCqZjHiTsKm0
oeMO4HxFVkGzRw9IeLl/D0NUSotu6pO9FBr3N6ebnlOfH6xPUuQlsPa+wN1I
8uRsU9mU/ZAfiQi8/LOKvL+RJlQUh03N4WCvznJZk49ia55X0XWj1VGPL+2F
1pkmxomPoh8BqOCbWDqmkXHAiOLoyNrgVkKOUq3p40YgNs7t+Lsvq7phf/3h
KaoZwi8rJ4YVbsEcCnIPPf97uwiG4Jic2mCzo7YVsb9CzpGJqdFBOuepg6Y6
D45r9xlV2s96jOAcaWIBISsgNcQpwM1XSiq5YHCSSIy0iA9cTps9KnJ3RB7A
QlWK96adTXIcmebzDJJiD4VqjzEhEQREVlXR7hfEEy2Pm79KKowag18yWuTA
2T/PBWYPjgalYYCildIu/7xKMbM33hQW/xrwDf4Y1/dCpyRYFwnKLZUVQpmV
3jlJEBF0B5W/D9NHJOsVscbFMpBkMUTxy9PEjccV99CGxIOuW5QviEmH5sNQ
qw7UiODeuAHwy91m2ldv/0ovidFPgt+XHm3ozc/VzcV5Fl3Is/EY4K5jcYa8
1iyRXQPzi13KxBX6WwQdW5eFCnerYSS03eO05jonumSuEXfK9dJazJNqbWl6
FELRBjLeD87oyr4mI6XdB8DCzMA6LDSXkrYGF4Qf0pDiKWrb6LZrSzITodse
t2lzcdxBsg9/tEQvRwGdiydb0bxinTykFN2K5gZ1zBEyY0g7D58yPPSZNOtx
QR6KzdgDOy2TxQhDI5rt5mkICGZ68WcOxMs1rpZvs8sqjVnE/rigFM34dvIX
nbrpoYaTvTMxhFEhX/lHpOJTbMZMzSPpPtlsweHHaJybqtpBivLKq4bhvK++
KhzDKqluG2ODg8+tKTVDspy2F4VTpJFk5y8pML5FeO1wVss8ORos1HAjSeD2
I1iyCdYOExbP7lsUgk5brDDhcvzHei9IxyXGcMeiC60qTn3pTAUJmzevenrO
/uMiZo8aIMru237YHFt5D4P9zvxSwkzE9HYZIgVs5xzqa2TGV8y167AQVh4V
M4ieo5T7BnqY1pWO1pav9aeQ03EAwlEfs74YTgvzTXwMhCoOzG5Bp2JNgRP6
KnSTTeGUeg9RJ+6eKnN7PREt46YiJHvozoeT42VxLiBZv51k3vmvFtSjP/VR
1BXoBHb63fwr0YOd+l9ReJ4XeJ47my1mFEGHaW8dtOJNj8z6/3+FaDn4bU/P
A+9tpN6aBepHtyJHolPXNy21FdFmczs9HKgIRxjx6xZxup386S24o75Pc2WK
PsMqnkCtUFEmE5MISLPRpSskil6r35BudVo8DzaIJooepqcnQCHRVbdMmnA4
PTD2t5QrS7jav4KBILh1sIisXqHdMjbVc3cToKkAHzC2RW2t8mvknDkx1ALW
wgwGz34HL+foC5AN6S4OlrdsITsbJkxYNQbGU68+JDYdYtwbrkxV3KvNCfUT
/3sfukykmXBh7Wq3cEquftWrbYd9/VVdAxDntE5AA7KQaLMc7e65CXDf1pC1
NVFpfhp/+SmZz+UbBLP6yyCiAu8D3ZmQk5E7QA0XOoMv1yZZamO4ejjxedGD
z98pX7fbhU+2hpvPMaa4lSdDlEQnIPr7aqniT0mlULiEaGqJ+eQH7/NGZsn5
f5EmuqOxCXcX+Gqw+rUqOP2Y9bQYAu42APiomUc1TMytr7mL07Vs/LYhmEuU
HHwGmaOjY3K6j+9DSpiH/TqIbtROvdG03vwVbY6+un65FIQxWU223Il5HBVy
Lf7+0ZL3eOgfK4ksCFl46aFuohltVjY8RCB3Iwy3FzkvmmFBQc7IXF4wl0OT
ySPpEWDeYFJrrgQD/E4xqFKuVlUVaMk+WCmm1cMJnwWuw9NEWEvS7oZIhb1I
AC69BPITcwbGHmDyKLBv3TFp9GFegyydo2HmmrpNe2ZQ+ghT9sxZPzDdNmvP
s2iKuXrNUXlEXhgRJc+/0LLZiF35NjbjbYCMivZD4pHB4UF4xaLux/feqa8w
kKC5jQFXeYlNCJtI1Md5+cMKTEu6Ndc4mT7leOclTOF7sfR0/UheDdhVzwcj
rn+UaALd2y53A5z88IPRqdX/wE1PeTnzIIMCt8ScHXxskHtJ5xKspdC+uB7u
GOoih33/nTb+/nDkxnZRGcM8TuSLI2pdlppER+nZ4CNFUFfczh/8G+AoZDnM
f/GxHRz9QeFgKs0gBOZIkwl5MGWvonuVkc1L8Gp/E3p74BDsfIYsfbwwPRIe
1Ii3Ary7J24xMtRXueNjZ1s0fpcscR6+0FtCZ/YmgIzY/iJ6+J3wU6YMhINj
GIkKwwT1DsNVq6ypcaTc7Gizn7D0LRA0XqX/+ujtVzoecL1zAzfufEo9/mtt
7E+VsGQxF/2G4Z3ipQOKc2T38keqk8MjVx9BXc7/6gpr5a3obLJtkuu1XXSk
fLFLITLjHqFFIk6N3O4J0LXacBQVkbmD1aZRi79medmofZvdI3B3F64AMv2U
HKly/tyISgKC69dlL0GpacN8HYi7erPa2wF2oiK6tck5ejO79ZCGjQ4Zw9qC
EBQgyG+w2WgQrAHVCZjKmSIEfoTVZO96YW7tgU3cNSAM01+/QEhyuROfuxd2
pTzKEvzwrFq5HFkldJNbLnakE7zHUdbRfv4rTR1LC0M0PUWYzLpRcyE9aiAv
YxQNIrXkzon4fLayQpksOUTYSev8lzKi1GBBVkUBn4/hT6DBvZ8mTyDAKFdX
l73VaH0WjTbiArH2IkH1ds5CNoWn4IOlAyRadhJQ8d5maz3T2V16V4FODQlf
fwCCOySopVhanoBprEFpJnaIXh6fesuMg+d2gEu3YNYG6DTdeQ3pcqZt5jKW
V+yACAeqDN8s8sBYbIDvPOsKZ5bEJdJz/WikJxieisdIjKPnGqmgMl3WUqoE
nL7vwzqiCPBM+fh5PDR2525Xo3Jhr+fWvs3uKRviepQbn0ux8rBwTrhBgZsZ
Eoha+GZrvl8GqZPCwGFjUOsrpkxzsTO8p9C0MhZq+2Vz3m3nxlYumTSWYsYq
UMcJgkl9Pnog/XxLpTd0e60zRu2DG3XLkXhS00Hia8GsY1bHQSIkabc8dkDj
JzLdgQeX72mz9Fh3+X44xylYbMIEYyvObWno8Ko/DxlfQt/1gy5XV3MlKhfD
rV8lPjZgzT7809Ptkq1tAfdd+nSpIapdAY215oxJnX6oQJfWxH1PT+j6d+Q7
demmejllFQADXADC4w7jGi1MzcyVg1UKR/jp5EOF3eB/3vRnYXB7KgUaZrJS
6whBx+0MD0pDqpundwGhvoKNe+3huawYAXTv+Y3qwBh5MYTZ0g+DldM+ZjlY
bD9F5XhTCC+DgFPJ0yxFbHDCDZgIdfm5b2UC8dwF6WaUKD74i9O4sRWU8bXE
vKIHCY5zCLqQo+fqirMHx8LbFqeVeCHORWYKrCeZbGPRijilIrFwZWPdpbgZ
fXB40P8nD897les9ArPzWUJxy4mueXSp9bY+YryhBYil3DgFv8FIvkfLUDXz
tvm55sIALdhZ7SYrU0IE4O8vUOS3hhK46Me05TQwqi0vSdhZpCsrq4Hre5ej
CTFRgeqrP9zlbXcVryYk0zyiqWAi+pZEdk5TZTjVG6th3XremVVIePjcD54m
RHP4Z2qO95nKuUuuBK6wKxxeikpNDcTGB8NPj49WzrLlrCDQHcFwHzP7BlKN
8McBVnL42vIK/MWuxFzcjMKhW7vVHehA8W5/1/IzgBZAMespM4UfcuEw0ykz
H9lk6tVYmIdGRja0qhBobSauhSIiFHDBpqKMVH66t8jcbZrLe6ImBP7xAaVP
ueTgmjFDj9fXLa8v2zRP2qutGMPDXAgOmgPqdP4zscSWRY28AY2x9lqKjyur
3PcdXDtEFG2IatqCfmrOC6vRj4F3goFdRXQ9Nrv410HmptNUS057GMKuOGzv
GTi8NNV+9rBcfOAnJhQkd3OdMRiO8l4G5HCHroytUOOIOvAUxVS5uC0CVO/R
1P7CZog20OM4ie9Oy0aVQD7rG9Iep3C6YFxMHqmh+JLOmDwwHJ+ci5fY5FsA
octfOkdWo6Bbm9qGOOOHahf2/+KC5kZCluve48isfByyOY+Y0p5U0immII41
FwQamdyLamT6THOZBGbAan7E4ONOpNUhpmOgH6onWb1G5uxeRyDef6I7iN05
S6VNeTDtjFhHDuz/7x+wdg+qdk2xvZeyFCsKIEHfsj/CnONFKbwNZaA8bI82
kPJBzpgpW2mNfObA6k6DYhpWU7iiRCnmn+Q/HB//315Jukj0ozdXrbmsEmdD
I8AM/e7Yy3GhHamG8s3QoI9LMAkq72jOZFjy3kaVKInZCSETlu+YeJ5gYFDN
X0xfWVyh4zcf6XhuxjXtoiq4HlAT5Aw2e8V2tJDbqJ6+YpEt6EiGfHtbpuUJ
F8NHq6K1PhNMhVKBB/bJRZ7L93MadI6ACoIgznsshTgawOKfdc6SZKdkQebS
q00wg3IK9FDMsCZcas0oTwiNd8kwRoxJ52F25nm19hlipAmu3KaplHMj/R0i
ZmRVcwD8o2EQAuqafo588yKnymcm0+Cf5k+zFNZEg8yx5VjBH2/5xsfSH+Rs
m0vrysO6mlrS1atabo8XzBlGy/64BtV60CdZ33cyoYl74BW8ZqzUc/d8Wv3O
qTUAd7QEv1bcp1hHTQCgb7ERYER+ZGyzI0LLNRLtyqbiPxxWniIVsGVmuDHq
QnNza13jGFYbfKa5JpPlILOGeheEnxJec2S4HFOWw8uKKAo1T2ZJDLTiFE8C
JeSwANCEo+L5XPPyE7CGH0aaP0enCkv6BKqapLOKyIv8Sl7jDlyIKYW9MBK3
BTsZBMbpatIa9ZdyhCqlmIThw7zjusUhgORptapGzj7qtYkqsBKVu2bMZCzS
4fZsiiLXzCQw8Lu6Nd3+c0Pf5ljZMIpNazCkfE0b0P9plLTmliFHmDv1N7sF
I8Zfu0UII3qzRRRY6Tq0LtuW6WP8D0rTzYEbItzHw5A3YwX2CZBvreJBZrIa
DIaY8MpVb8PPiitwauN5+dr9MIiMqFTxyDV/dOYcXNg+bCMb/8sBH9dS2xy1
UAqBD54TLTMxfK89x8R17vi8TbNhG4gFdYKoqeaHW/Rz4yK+eT1JQd7Ox/dr
eScutu1DPHQc6G6uPFicE7I+oExBnGgIw3dT/yNiUSVBaSuWFNYOIN9jECax
ILeQ+NVxKKqbshhI5krfijJ8BO/3arFfq6ulxAorsVfNuOS7XzcDwFrzZSYS
nGwR6LkCy3R8HkeKjhcrhCtlP08M98XGYq+W1L8bvbMaDBMvKUAqlNfxTdcs
sm5dIfsYG+QYutXYZSNS6iOab8iDH1Ri/1dGwA9/tRwJ/QN5olIiwd4uwvfn
MBGwZoLiNw8fyrEZvACpaaYkuQYm4z8f27jSxOoDiUUFmjgW5xFOtxWcqwMn
DRQjVzAzhrWMIOzlWHAxDp/Fkxy7y7gHAYHyj9Pb6qrIsTZGBCjX4Igix6fY
7MB6ZKKhPF8UurWonHIL7A7mL0f62QZroPveoFx8tsrsF1Zk0jCOm+ZyiRux
97Lhk4I0ObX0aMfgDVKoDgPG6NQZ+Kq545k0asupcPY0yhhQLbZJbWDxMzJL
LFwcmSYWDCjiDN8EqSUzCAmChhlz3Y5JWQQIQxLxw4/FI90bwBwwfTlCEo8P
P6pH12k0vszXlXvTMqn5le8x78QJKsYUKMzsMTadhY2XTQGZcFgpaw5skQeS
BukvvWUX6KhJfoe1vrg6OO+zOfiLOfZg0F726Gm7O/Ademvi4k+9ZbHARkXD
p7xFcPb7hmprELCkUIaPEBjZZxs10CZZ08hvIcY4S+Zz6viA8CwOFc5gONhr
+aqAtxVBfmQCDVvPqMez0dK5B67btGVuNa02tPCvgCBoTAdSDKBv2VD2ba1X
S0cOAICAR+rQlpe68oKoU1Z8U+0xlksVT0Scpr5Z421EBTTLKnKQ8veubdUT
UTFJvXMbPMS/GHYJObZiwSq3TXdIwvXJxQpLpgPUMvWJ4vpTWnWkP9E+yD/n
UhAF0h8SaC6sh7oRt2N6DYvZdJ/Kf5/XqEqWVIydp2WqzOVuZV7uood60G+J
VmxwTlSi4O0iJ347FjL0DgLwhMW9G2sswxjzIJKtL6qAK0YbZFwGQEwHW6k3
oiGZg68m5UgCq234L9PRet+J4g+kG7w7RXRtuwwq6+Bp5rnkE0imWE/Fhat0
Zh4dtoV8xloFnetUdf9YJ7f3kEjjAzfim87u10n89POqexnD68m9riW+M42L
YC2YqmY+2D2t6V5YMHCx2aJ75xPBSCn4cZHmUuuN9T/tVOaRUUUHNtj4rK50
p67NjtnJrWUmDvApMBa5A1IhsoCYkgRHvert8fgP7wXI5G4uSXVjPS33yWoG
Mt6t/SsWqeXcaek95ACh6CjY22d+7gM8BZKKCBFmjBqFRKD9Gl1auCc3MYoq
JB1AVQmVxpPoOntR6h65wWIfUDbX8RdMHgxnrpbbZUIQOSU7T0LvyY9ncr+R
zbpm9+2Y/FFAr6OappWoeZDrMsE8DN7Zbzf2ErUrX8HvgXBDez8peIdEgq9F
MV/zbrrUvdATvdpH2YCDi4RlwrD7e57SSAqkxwyXX6eZgvjgodW/5HEIqbtv
CY/QGKslSpyDCgTf0YWBKvWOQpwBzkSex2gzuU/6emMoHmKZsetT3XzisUUB
N0ULEHgzZTrUbx8RFYgevatWGEM2oK/qAmKvX4nwGUnfrIgfejndpakjGUjd
A1PV/nlReRJgb9p5LskmCQZiskGmGSy/YGtM6sFrah6iqgq2Xt4EII+k2jGZ
9d7y3r6kVuLd0pky4xXOyh2bTOWGLt4f2vDP5pOBJy+jvj7Xoiz6oU2kIDik
VR19IwHXz0yM1CqCPs61bZ6Y46l+dVv+2o+ocaOKwUKJ7dUckEkzfks/sh1/
Qpm+z1a/fy1HorBPuYvM98qYq7S3Ucnc6GLRdG4Wat+cPj06B/xp2n3vDby4
DOwK7yUfZLiUjUdr0AtiKSeAIXgooYLqAaRWlUooMTfBnhxswPkfMtCT85gN
qTnTiIAxUyCSaVm1dVxggXiSjZuaeiUe1FbXbr4crTW8FYf/+BVs07mqaWMV
UQdDrXSklG0ScXG0unqy0/yuvxRPZSSWVC2EWjp/TuOORYIk3RIu4+EUOwY5
Hw3IkVrqK+edxkay/hZtRoNvM2L4nS/7S9mv5wnJB8QpEHwqpBwD2umVRaHM
n48KavzGieN8yA1brpCYx8Xxy3dRZqYxlDcAidtbA16pSfJPr8G+U7ZLSryO
JXdRWZfaMzmglYxtW3d/ZgzEwTHsBZ/7FgPgWeAyta3LQLaj1PR5piGZjVo3
sUybwA1AK56uM8p5vNpcxxswjCTh2a4TCOoNYeVsw9zoGKcXVBLFchjdZS5u
mDBgrB0V93pBTWgovhdQwAmcItHSh6vQxBYg9S1HUVrJTiSijxVrObKIVIpP
/3iRuLVjoq+L9VVXz2GSY73qpyltlled/9W+KiVRSToYqXg2dsFlzuBKy6l3
Qq0vshxxLKGNRIodkNjJ0Pu56KZXl1nEgPDC181a9xp6M/eRocLRUVoTmxQ0
mFuFOdNtN9DBvgH5QDjvQ7X9y8oBv4NRd3FLtgWpYGBtkfUFQcpPlKk1vNCL
DDbPfEozo7BiemfnzWFx2PX5/j9W13ucmiiyc2851DlrlncHt4pzVTIKSPYJ
4Qq2iFoBP3ehjSkJk095s59fksNR+VICZkOBd0mnXVZCsLF7X4SgCky/kTen
/EUbYdbIKmeJk4iFnw1aJL1ViDZXmOe5A8A4wesWiYH2pS13dxFTmwIHwDd8
FZeKaWTyWOOd8nM9u/+74zE/MNT4Ma5dseOzQ/pQLq/CFr+H048ODh0CekFz
JFrRkwCzEtxOdv25XRQxHtbDZhxQ/qIDDLNrqxoUhUyyvY8/gyS7SnoTUlQz
+EpWWb75fD24eUg+BG3Mvk186ifMlu9DHqNbCXEOtTLVLaXnrIaYUerJSAAR
/qVvJMigVINwrB7YDHSfvROFWOFNom70RbyfNeTyvg9Owf91eFoXmjTZ62PO
lDADk+IcQEHVH9ILSGTrU5QuIDo83GHWRpJQZrbs3dmEjrihtEpAOQ235fqJ
D3r0mU0ZpnGYN0mX3VopfFMfNrs+iQUImvWFhC7O03auMoCATZCFUB6pzQo0
wPCD3pwdIppjmfnLxJ6gcQW2lakiBwtq6yZa2VciKLkVl6qvCcjYhBhrLgz5
nWHR++xdncF0nWx5VqIAHC58L/raH1tAA8tnTnpKudWit8h6e/EcfpJRI9Lg
zKNehjxhWPoxZAGlHAWAHcXaKs5/hzjwdXsYJl089GShBnHmOcKEWQ+OMuWy
dMQ8tSMI0IbqOxWd9Ghj1JtdvfFeWa32L8Cgnsq4BmSiJNOdPdD/M8QMOoxy
mvtUKi3lI33gjgfdkK6WtbbfutVy0pq1FvlR67J8Hj0KIDWXhsM1c7DShTEl
p+UqI4tyxoCFsdfe2Ot07oePAcUokCZ3PIb6IkCADV8jNx9L63MokLCTV0vO
rLGzn+XAAydkDjkPI5+1nngS+BDYnNLPMU+F5roMC7Ur+uQvZdvShawlw6PS
xzlPjoBlMFRj+ygOnyw1Exi6fWyLpMaKvad9tAmVKJiKRYy6gXK4hpaaPTw2
yZGQYY6BrS3bSyTdyCA3s4887F11cPwC4wuZ2Fk1XFm6REJsmQSdgtfpfME7
fBWRSbz3I33lEgXZ94DTv8NVByrtk2L9QCS/YHSXfaAv8cClbhf1lz9iExPH
oZyknwwG2tutld8Cb3n7Sp93jtgP41dRgntdDYUuR+LRsb9R61JuHRtobkgD
JFLuF/ETw1AFVdLXZqg7iACYSrf8QHwRPVd59Gf7koRWsFwukS9+AIN0U6j5
e4fRiYMQfrdiUbWY9PFmFfUGyUnVA+ukD4q3fkdFxz29kTAaHmoeiXEtoFpa
ryXQ8Tbm5m3t8YCygOu/fsd8FbIlYEWdZ3d6CD0ygXDExUboX60VSHUxN0xC
igu3gghXlN+im+uq+oYQdVjEsaex14IVPnO21grOhCCK09KgQBkRiihvKG4D
pJN4TJbLxl/m0aQ7Cgc8mEARpF1UhGPRBoQ1zF/3wejupyUu77gaykgPGr8q
ZUOHCAzg80ZDAg6g/pXvnm5HnfSEg5qtuWqoqu68VzDCtSq0p424+W/UJRZw
2RLrqensiNw/CGWzc9zjbaKThOdudUIcUIw4VW1Qs8UuwlOBUogQYAmnC4Ym
MqEflBn5aS0j9ohGM9XG1VLODGK36MW/bSOWDNJJRLpFxYqtVhOoeiRbpUQA
x7rXPJAfw5xsJe+4OTx74hB1Am4jpFmkiOD412HRg9KHBYuqXbwhIf5s3190
u/udxu17bbosJIMQdvneuC5vtBvbuCr4q0nFHQaceiaFcJmvkD458KLrAmpW
1UAKVFvKQ5jn6YnBoV+fp3TZ1Vs1Q1rhEqiX3OgcN9R3TWCFRI6P12uLXpXC
oG3ycUcEBMOnjvSJvnIZkxUMuZdIzTvero/b+XBhqxCpMf/oXLzVVnqJhTRf
enMdQV1F+IHsc0KkyOkcj1p9oaVpfo4dIXtwEOmdtLXrFBF6T7xIqdWypsb/
OxWKHB1d2WNixLgQutTj9a9zwT6b2VwtshHIwFGRXcRv/xvNGphdAQX27pPA
S0XSBosvkMuDK4DRuxgUkjFsCB8plqY28mhNJbtrpmHt9iXabeZKaDdqxvN7
wHmpiktim86KL4TcJbmMqHkKLwvs10JCUsYpMwwgZDIS+eWnFdIfCjSwU3o7
7OqqRvXDwQyKP14KB1iPuyVrgi4gdLJ4efV3Ca+tOIAUORr0PIXUYzD5rp6K
hDphgcFiNs/TKXZ6rPa6oo+c3zsEmbK4KaI5TEauFzNyjVY9DTmG84Urfvwg
39GD9KyQTMpftRa0gWhSB9nfH8OmYhn3rh2LA1mYrkF7Bg18ydUnS5/2qhxh
rPHSR8LbAUa3wObEYJ9tz9ncAEQisgvL6mGSWrXH9YPZTE8yZnHz3BNB8ZsX
SIuHS2l1lHlHrSdUlVFIDFILN2sLaLURavfofg/RgasKlh89bw6TqIKwxNNW
p7csoIte9VHNh1W+H9brk9PFrpDGRb734as4eSKMhgVcxZuNdhtK+L4jg327
bsACZH9iasD8GkXAEFawKWtYlgkui/r0nOitmoDSpcVF/DgWhZtY7e9/2LR0
f+NZmBI/u+QY0Elm2tQ31mdSDLZvvvlubhLleqgKPz98y4v8N9os2E7C6RyQ
S5PD+O1ImFKM61teSlWw1rQsX5HKoZyPWAKuF0iT5bNwj1Z1pwlgB7jH11Bf
dlWan8fM9lcsnuvRkZ8RzeuRNN8xG3mWix+8KZdnaQPAbLO1IBJvNmvIcMQH
gk2TyS14464vWk39WpqTN/JGZTqIhQvD5UXNw1P+cKsUNg487oIhBr26Hzqk
ej/aeyl1NyLZXbeJvJmXDswpoQuTn1nNJQvee68HSsel2Ja0MyWM6Cpcld88
4drTgHPMYFrbjQK8oiEsmmxOwHtNCtNZ09T3epfsYDrUArLYlcLpHXFgJUwT
PBFPTinf+S0gojsxMKAFHumB+pOPK55OUGzRShD228yptcSpa1mcXDmM5HIS
7vE1EKarBgBNfulEtrQGWyI3+/vOcsBQAhBcoIDBWXkG5pXr06et04LZzHa/
kFkdZH3yUDxjqhzFf8KgLHiNogCMp99jSBVBd/wsbOGUbzB++3HtXmuu7iWN
twFDMfu7mLZ2jhFJq6LG5IDYgsz5sPRMDx7Yj1/2yaGJH/mdUEWMeV2UOBd2
PaulENIDoCp+sT964ZzYQbLANlFZlp56ilQXssuilekA3klSCkbp/DElDbtp
w3Fx6qYubJ1GqL8C5mXfo02lkQi/MaOoXa5R5QojKcKMJS25vlzVgXxCXKVT
dkQAFGdNF/y6M2wQ5+87mj3T3TOQbzydY+HPp9S5TxxMBEN6AYOZ99ii5ys1
L6VbTqSxzfmQumofCAX2zR8J5zgnkOmR/z6eYulgsL/lp8WWsrfU7NAcy/OR
F+otEhPdqyVn4BnbRqZslHUrRezKN4YMll2+i3zsTVy71qOLR0lBhn0xdl2t
2ysdm1lknrRk9UAjOHr+YU8G995qFZfX/SQ+ZqLUJYKLQLTqsSrf++l4XZo4
Mpw2Y1UCyPvdYdSPW260OvbelY57yI1RRrh7GlgKoc9x7RgKIKPWWTzwBcrf
kxgXkyiK901ZBrfYvVz6nflCjLHDi6qurUSfZKw8ZQ1VHaPtcm5SMJwfc32h
RuEpGkh4+uX4tDJK4qWEFlPoKALlDSqXenVPCbxv9D9CqIRJ7Rg8Sf1peRF7
WIKgIdArW59ExvYq+2MAfZrQ2dmJeHR4HOkUJJn3+/Sfa9yIjSvBeR/vKzYF
lMatmZub3jIDU+XMsTAaoemMgjTzctxOqwWk9Kstbd/N5aYigb3oHGRWvjdc
n74D33lGuW0dN4sD//ro38jlHLpPu+MOg2TbMwEJGjBCUjt7Bz8KoYlHsIIn
Lt4lATRtWCEdKF/d8/bf1A2l3kpTDbtlN4YgbMjcakk4jWRRDZha5lv7QpIP
fUKoKnYV/18A9xq+0H6WQCi1A1P2159O8sxMGafTUvFzup5Mp+f6xmTx8+OQ
Fnjf7qXIindWkysCd6m2On6zWdr8c2h+mO+QPZEXzsXFCrcP4OOdPKFpMnPX
XsQpqHTE9cFJhydVry+GrOcKXrk/ywRuPp2DvbQWAujPagb3qLP57Vn9ojCM
56bTQNwpvZoeQuT2A3IgQtpOmmGHOEvUePcE0r7rye5IUjEj8SLp9vCfko7+
m8P1nLg1jqrqpPEtLYYpv3VW7NKRPY72/nNx2Xw6WCDByhsNLYU0Hqao44ez
SXzP35BIhbTUu6tXM5xa7bmtOZbnoA2MfQGFYjQzUWusScnu32FhzQsvtHjD
Y2WMNsze/93GdEenYTJ/7a1wqSQHUdpWt6yp8ld7esJGFiqxVXB70IiPPhUu
T2hy7Kin5MB6npuGaxF3RV4IFCKlk5QMfpLFCoFPRSVbT2vlV/1zb26IXJ+7
XkiOC5xE6pcbh/EeLTbBvQCqEM+QmNUTPmw6RUdaBKV6Tum5xbn0Tu6MpIXc
guxLfxw9rOsVglCHiWRrKZ0nfg08uhuBarEDZXPJ4a/qAfz5ZvjQM5TCPQtI
cCViood3Nle1fTjgqAqAT2p9m3/G00b2rFlBN+GwbnBWmfkchk11j+ihnLYi
98bxtzb4iDXp+f/pLGshQj04hJA6S16Xlq/ddyUIM1grg0fNOPZYyW3QD13i
Q67tASFUwYjBvQW0J4y1RDJq2frkd353PzsEi39zKkcP29X2RNs+wODAcOpL
6ABrdoIlQyFvyJJGEkHGgOHti5KMI1OfPOj/ZRy+bTA09j944fGxVO9nWeyT
46KrmGmO6l3SfpSJJQZ1t20s7sEJ5sENXkYKRhv3AQBEsAUfn3JVNfhILnQq
YW/Nllo3p5Ud4jcCVaVaKc0uVP77I0d+M86GluuNwXaHa8+JFC1YLt7TtaRX
DK8oz7o/S7kk+JlDCtcOf/5ccIXG6eDD5Hl2APU/WSz7o8+n9toB307QSwni
8MLJnhLKgwUWb4fns7okAF3eJuGVasuuM3QzaNPrYoXxyz/pE32yjN8tNCNw
0oNAflZytRV9bdaF3TAOeMg0tB+LQXrO+cQANphb3dAgZkGMAdp8XN/42rr7
Z/eQgexb0QZx1/UnLbBvqrW8jBAvLBHp8dm2zHSA3Vhwi0fcVtnBlJ6sG7Yc
fY+PvwQPr/P9V4kCJ8OC+KjCqpV0kV4a1iSNP8IU1SP46TKXypBpWollSn6H
d+GAktXrrInnwRgrtikRy4EhG7SusXi78oujdMZmdjdkvpG0gxKytd44lwRb
tOhu++RDzTVLau2jmokvMEDmYljudae1D727XcGreaT/YJElfbqicFi4WcIV
OXsHqbbptH43U7h5hTV+oSWFCD10q90+KvCZLy08hBi+jSM8/tKaMlhIvpxp
ZXMnLem68F/8v8OMI1HhMxXiaZL594f74MCUz1EcSfuEFPeDMrwznB33S+i5
ZOI5AFI1Nu1n5CPNL/c3745GPc2KFmIr2aBTz/I1ZblLLfWh4Qp9/hw781Hg
DOwAg4IYD6jbDJGtsJFkEpGyOPSNb/fH9xvyvClZpldZ2vhLrei8ySLBbrUz
nVCQUJ/n4L6L9W0Yo1Gd0oKECgUfzMTc/2xnLsBPEvikVqYJQ/Etn6U3rD3q
iL+1bvwnMv/IT7VO19C2Ygtm8NSLCMN4C6l97nVouB/8HEnwlNF9L9i15LmJ
Ma/DinvIsawgTdqE3cvDj4WD0BdLD2lfYMl5dp0iUYp0vRg40YH2Wiv6j12m
T3EATA14sHU3sJ+L7WvlOQ/te0b1vFeBRM8076exmFsRu7l+/AC6atGH70sp
GkbxECGLb8my2CG7/kfwPX/QM/3YSaRChlASBH3xupqSLp7I3PxH2T7urh/M
REUtmClN8ZBHE0ytd9PqSfcXUC1zmSMVEPZWG13A1atCLTuXf4R7LVuxDDHW
0kKNc0br3237KdA7utUC58ugQ+R+SDFI9f5v31qh67nIbptHSWCkCwmqizem
Ai4dAsJvjDP8oNd0zTwG6fiZ7p5hjMr6YqotGKWJOZ/92tG4NmeE9t/+BSn3
HbFZakMKUluZLyQRJ0k1zVnXH44PGaZHtHB36FIL4p82j97u62wfgC99ii+O
buJtPEIXUrBvqLb8tDT7gtfX6qxtJ78ln3zagCMiBFHuUF1PkqDM4kWCT8cN
N4n+YaAERHH/zCMmqzb2iiAW6mzBNR2JGRe1z3N6gdiUQi4Ume/Alh8mqFEJ
4Z8sqOPNjqC1MeRKbQRjsV/6M3fvx3b+xX2kmLHRlVsBgMk6rUeiee7zpsfq
9mOwfTd3y7DdQOGpcGAR2d/i+wtr/CvVBohysOjIof7s5sUKgBcb3M/cd5Bq
cIeZjYHzwgLkqGXu/jALQIvRKaQ08DRslAAg+tPp67Z5LlvJfqO+6ceVELRB
YCITkfdHOyGkcmHN6ByKTuv32MCTa4gZJq12ZaSdcMtKJ/O2LanBoY5xQpKN
NbvKYR8wErmvC1xqPl2Uhx9KcobG0fRzdUQkY+TSWOXAlLPY4wTkFxehlaU9
Z7rz7lvAc4ASdvFubf1xm5LQZ+FcV909ZurBXQ4JW9u53t5pTXL51r3YjVNq
VLILXnO1jowNUMCixU3UgjmusCu2dXN3l2w1tlPQwZjgUncLKk7cbP7QUMfI
bvNvC7/+jlg9OfSEvuGiAGpwgsrhNWDtI1kRbLcfzBwoM50AI1x9a2jko69W
wq3i5sa6nfdcWcwKnwZYAMz19XohBujycCF5sTgSYwyoF3+adaRt4qjjzPva
mqB36GGQntQRJrJMHVblSevu32m1XnnEVkmOmd5M+yYfpDnyiRRJtB2Ouix3
6FEZHnc1YbZiqZQGVJOI1sKIObGUjcRW0B4DbAR4d9LXBV/fqKSHCQbaZKVK
cBqFCgGaJ95cfR00bIMdIeHSnjrc/dZO/WWcgiO+cL7aJJSHD4ro1kwVqvqP
TPkH1mQDg7RUKKakyuF2WUZCyvf6AmO0TEy4osNmbz4okWSuWnd0qLTtU3Ha
pVXFFkTzMZLOsu//GaGuBGF+cajqEVcLyenHn1zaf/mcDKAjdsWZhxqhDlM6
6/z/a31xtabRNhnJ1/RogU/J0YyK/quSVd5i2sKY2b3NCd6cjogQ0g5WLNnE
g43ZaDsTCYZh55dcTgSMjGtQLrTlB1k8me/cgYyoYOgEJV9BAj4obUxPA5zJ
StOUe0W0NNll58RZvwRqpn6/MBRi5rXVUYJLyXfUIBPS7BRUgVPfcuwA7Nc/
CZy1845tQ5L9nQb/bGQkOnn1TNOdx2OfCeo5sZx/6xxs4KdzATlGJXIbSoCS
bACbj/GKEjtaf9jtS1yhiso6vH2uxggFT6Teuig/K+wKzHPoWlQF/czEKhVM
OSTjHzAOKr+AZ5kH8l1GTpmbRE9cUA5M0dq7S0Bp4cqNVV/3P3wHPbQWbncj
MYchnTL9zvzi0jXcimfQkYqy8C9uE3hF99b5TQLlNH4GnxA0SKyKv4Aj1YG+
XQsF51IU5et6L//v23x2L3rmmPYYhEm3St3ypeWgkxY1M3XZ9ZXWs/xDRL+u
DQp5Ste1RMTHQR2AZXgWXBFLZ9K8iAP3BTfhOkqAvewXdBl3SYJt5CTDCrR9
XTyLERx5aVJgEWYxzA4pWISdCst21RTyny0yLAywmHqSTb2Ov7w26VuoG7v4
hFMb6vEfSdSoqD5zQ1s2HWkeS0JC7UxeAVEw8EQriFEhktZBXcaS3osAGXWs
xcFsj/o/g+WsvesNe3A5m2Rpj6o6HvHMvG7VfN8g0Jn9yKFinAS3yL9EiHdi
O8TiG8gB+Iqe8pteKEILTYZD8DF049NP76SxnIwgXozRmHsvH6eRL1GLhIJw
DwKgjydlBTcfEVVUTkL73u29UqxLbx7ncaM7iGrcT/8R3goaGZlKjol9flYv
xr8J6rlODA66ZCVnhCitJRd9rWIafYv4HjtyPBSTYw1lPpemaO29Q1KMCbkk
iJpxKDtNv0AsGZP4sk2Ai8/vDmirHuh9fX9gr5pHIgF5G+Ms8UCwUJSHy/3T
Sg+EVcwelD1y3TNKYqwgWgwDoFJJlxvQXEZAg3yPli2Sk+Csz+/Zeb23DaFl
NQxNsmYhmvLIFXkosYSa6TCGlDKzlommeFU+EZ5KNVfWTJbD6/aYLAAWX3zz
R8eyatIIK2FrwUydfxsDmTEa0lOuM3hWAsR/xNPQ4pvE6ml0dV01dfJaNDZC
UVpXMlfrkBQwb8+mhnSzjeMUVB/ex8r6e2rPEZXTU356s3FbsEj6Fq7mDa+C
pTBrMoYrJwM9dZBm5psrQc8RZ6ghrYv/s31Q8AcMT/6XAY6hFQDD2FwIxs9g
KTLXmwOyEO1SV+/kKPpKGryuL5deUMtUn+dzltB1o4RmV8nMNSkI00MNx5Ls
f/hkZOy73FvOvKaZ099nEqzwr3zQJNVeIpcs4bwLOLBO1iBOCSl+TZbD7Gcg
mfyiXA0g9rkt51pEFnh4xAM6iIkFOQJX6vIuk9+OnR1+g4NANqNqEn0ucegm
M9BkuKZCFiv0cAF5y/zpS8eP15CT0/hwYoBkHcs+eJClGrU7Gh3kyhceOxIl
iYiGTclx2zRh0ONygOhr7hd6peQwnf//FRicN3YST5OWUMViQ2MyYdOKFTeB
+0YnWOLJmTvs/AUASTKX6uLA30uhXnWi2wzobQOdYxNhXKrqvbek4ldE4TFE
W6U5KDc6LxzI9pt2ESJo+CaOJiNYKYmfCFuiaKUWfDtG+3FQIz9ukzSFcYIR
t5F9EoNUYIlo+GwKoYtRjSGvFoMfxFIsE+L6k1dlGMF36BbQyV5gBCN9tgn4
MoX/ZfOVcTPr8w9eF7FNNSMg5+6F5rWqqULusn+SKleQmp8vzaXKozMMbMSq
T6Oae3RtcqhlRDrW9LDpEYHIiHR0ypUa5Ok0InJEeoAmgAtDZ+VV+86bRVGZ
+1dw5OCfYPMjrWru2eBo1x6IdJOf+jbkaA9JCbQmzQzaVidSP9Prui+CzCKz
TtLIowZVUF4oaQ1VeDPnxf0skUXB2TJflhy/jethc8hDU8F0fnQf3L82bTkv
t5awuAAfSN2Ig43Ll2bKE/NHX9C1jOXjYUZZJWZGWjAmDZn+HCk+SMu3NcWT
JzM3IAX0B0JlTilkEipqE0pb9oNvIy2Jb6D6cF+o6i4yKyH5og+apIOf/JE5
Di1Th9iuaOy/dLlc3kXubc43Hvu41C+M4rIc170TjParkUXKbzazbi35JJqM
54IMnGDJG2Gt8BLAR6F5NSRZPDtZX3QiriFAcw8H4jCUfW18lGNeE6s+Xx/w
SJ13yXtcs42TiwqiIA4hC0nyDgnTD5tumrfIF0C8qWzMwmX5p7msKkvaw6Cm
+tLzeKje7olcUiwayGvOnNcHcdyPWeQW5iN60c3Gto3FZj5hg8w/IaOpE8qM
4b3GMtfa9PSSDcf6B1QP/fQPa580F0+7EMwXNovTR725jgcegiCK73lC2YdG
rrpYiOtvPq4yfzLaAT7e8cJmpwhOof384SXBypw37+0TbWKIbd9yn4D68UQX
gh7BU7ruxwWNx7ztOm+M/bKlA5ku3GiuKZ35rRTrv8yg/Q6l4vyQf2dD0AQH
hdjTUpyQKwolbBdbcaLksZFCuHq8SGhHso2YBOltS/7it3rB6gHqIv4ZcEm4
MTugp7NVISNAc7zUYuiuU/cUs4BnU/6ygtNe2B4XbKzElN76FT7uYGay7VzK
FpNXg5BZkqy5WXCLKtZ8gj+aSyOZzJb+bLaHDHhBIN9zI80diqpFf/qyY+aE
W0dsyFjstxUPBbmsrTgYYYRci9I0LAOUxTS93McZHArJcUkf1LSFaDvwQrA6
3siy0wMxgdBQ4ijF85Hv72NO5aQeeVCKAa+t1u3ynVaExe8LYhTN0uuxf5Yq
TGUVSgD5IZsuaPGTzbkA6+jAVmQO1TWIdMRELnYMr2AeWKvh2LyyoAE2RqEN
5icWzdFJcpVgTM9bxWetRGHWMmV7E4zMr4Fm0qoo2jiNSh/WOYYtk0W3r03V
XZlSO1Ko4lhGN/+Asqaukj98SQJ7gq2+vcuF7LbpDA2lMZx3Kn+ljMb532+4
+i5N+SQ4Bs7LlxyyOUnhTm/PcEY4s7mUddOn4E/m4u+cq0v4rchLavfiDpvD
jaiDaJkNTwYRGkEr1e4bq1xxyQcU8smoQNDQ4bVLmBhuLW8dUAfZrFRsIQ9t
wwjRUl58DOtMhThDFvfznsyueNi7pM0bipg9dlYPqrOHEt35HrOjNROeuYZb
9EBtTgDezDBlJs+dun/SKwwQ7NLoFV1jmizQVF4DU8MELTfG8o2jcckwVFJF
uw0Z5hb/UM9a285HcK9IjuXGG7P/VHsbfL02l9CKs10GlIJ8QmxP2MJ9DXrX
fdm2l6/kq43Ct3SRdP22pTwOLWG7Nyc1M4yU+lP/Y3fIzW++pAS28Jo7k1RI
yYCU7dKL2DnFuiOKLQB1uVw1YkPM2hb8RtsNXVxgo2VCfF/VgVlnbRvaQhg9
XXL2Jfbq/nhKRnwW3GGZSwaV05VG/OaP0Gidgmjin1lV0pjz5YihTcBbTkCL
iI/UfBhYhlSGsn9fx11uyW8kGjiYRcV7XiOW+kXIipOMUQIUGf0IK7PFN2aq
PuNyoc1RvJ80ECfTO97Ty4+zBdM8hi4cBF4x8y/K0Bnt44sE6+R86QZS7B6C
JFR2p3SsTiizOq0Nt9qhB7Jn01sFuF1EkxQ1ybKRjMZWtfIP0uHvTWL9wAt8
/hyg5CnDbz2dJfgGoVnP/3B8R/ATvGzKJylGHcFBRGi6qlz3BChlGgneBy43
0WKArruqTiFj6UmzdFIqc77i1wuDPhcnTj/FVJqCFGL86KfX6TfgKcOFxxRr
Srsp5mXuQUCI2YxK8nYYIuv3TbYvhXZAAFLixRe0JgARSDKQDYNeH6lcMUnd
bxmnYz64uCfB4Peddvp9f7qgr8Gd7g92sGe/QulTYMpfZwy5Hr9GuX5FPfzq
/pgnuD/DOQIlgkrqsUjqDox7V4bg2HcruWYZVz+oIume/asAm7O3L5j0r5W9
C4AH/G0kme7a28ojrKv+XyQBJQDLr9RyegmBz5kTuPtZ+7KSjNbTN3FjJDv2
8HlET3YrQ4tDkTEdi6DbCzxMqkPk2bA3rvDrCqfNluQ2zgFjjQ9vtzDxAFLU
CrHHSCuuaSJszOqkEHk6nwx8UE/jP3TT8AAaJ0BOsYGHkEvvjS3Mvl0a8T7I
w68fX+nhi7BQom2nhMzoPjfpKYwkmUZ0dCd7FqDeIgHm65HKKqvil3KUOD3E
xZ1yWlQDUczAn2E9kSP9mYzbE5i7D8W7sOur2ZOf2hNwpUzxbx0kiWr/fZCF
t98cCFTfXwvAR8h+kkXXyfU2XekM+2keIA3kKR4+3IWijmVytgt19Z8fVjNL
Z8quLJbxqcwl4WJgJnnbUXnbATfLDvOEBzKFM9ivblWe936r9O5s5ay/7nLY
9wWEXqoPTvhJekuuLbZm78Bv8oKGU3opelAJgd+EXjCoG5myn4a/tzevTax/
8/VOKSzzCF8nVypDGNtu8UsnI/x2FYy8XnvMUwyaj8bck+v9KQkHEtTlDNg+
E7SxZbllsdmbb9hkj4YlveHJEcFW1zU47iza+Q8AB/JK2huQvCLlplJirbh8
kDUIzhRxF2omRkX86irYBG3xoMInC2pSPDREn5Ro7zBesV0oxL0722R7WTwL
xmdmFHKaqAj9pSdsXnu297SqIUyJY0wa569lV3flrgh8jtQr8RFtUgTfEPmL
CDdD/0B8xLUZ6dutL/cyIPxBiTX+9HGCAVymcdb45mADbQJaYsL0l5W5a2GC
/9pXdfSoYLBE0dxFq9ro5WerTzcy+bLjEbw74WgaFCC5ANCp1/BNRMrC/x8v
qkUbe3bqo0uIZk0xLxlnxZGkib6jqvdGrDjCsytxdmKSZ2ABx5bGb+weroTP
RBHG7pKDVTuTzd0aSqwH25gaEZnOAF3vCd2WdrK2Yd9DRI05pW13uMLSqf0O
iiuLNFcirQbazK/eqEinU4MP5XmPNH4zKz7CZyv44Ub12qP2RI6RKyhqpUuO
qeNvCAko8HFjidv0nDodMLrBRYX5l2yU/oaT4z0kS7NA1Yo6d/7ZKWilxEUl
ul7ZZf34xRuF4WI14unT+dcWZpI96VCS7SY4d1GjjzYW0EkR+Yk4gOpUe7eh
CURRIRMvwGyb7wAlIn1AOUxNMEZ3gc208alKyPRUKAWJvPbwCF44u4YMbWFi
Gtpo5anno0rGl+XgpOUclpWcknGBm9A3NTKc0vWoT1MIHqCprOAFck1xnXth
nI4ZPA/o+Yle3J8aM05a3Evd+oDK3jWqRJGDN1h7QV15lysHK/F9Y+IU3lkr
mCzLtgo+e4w21BqmG+aH9Z4xCnfqAuZYalIX2Oet3k4XuC2/yUHJuLJYQuiM
caO9bXJ+p97xjKaVHeIYhb/g/yInePQ0jx8iGs9PDsXUmmP74KaqdLJ4zgiW
YymuLFCjGH8GmOuKqPFMbOVkKcqtqCBDLA/FGxYGnKx2jT5GsrD23SeaJjCx
I12TNNcqMgg9Pxe0Abr5TQu1XxAl9qTiC1sjnBrHq4Bcj1GpVXBPDByU2E6L
c0iAvUKiQJiTaolOqD0TkK2DOVn50myqG/Vl14iAbgdi16MWhnpHTY/e7cVU
e3UhaCmEgqgtIIZf3KsHgQVPXa2hDkY97mDkCSanfrXAlhaJ/LqNxNZt7iLe
AFiJrdtlAVOoKOu5yiVnJTLNczLI1AtI3QlhpUJ+YgXEAC0XFw1lI5aQCSd2
wTmiIKgI6ItS/lgcxYAkVMj5INEG5OtFWku9PdR7HdMj4haqvJgjQhvYix0K
0jtUvevDyhyh8qGX9LtZjyC7/dLbO3YgDdyxGBur3Cl3IpihsHF4PjdjeVL/
RMlFai8vYKaDNgwBILhdItalAu87/2m1zEqhfCWCnqAAtUralqiLJzkTfg7E
TInzTEXfxcze8Q6xtPGNKs/lOdp4OfAxQs4BnSGPqSN9xzb+WweYmEYmbFC3
KERsDD/cu3ujf49UkISYNf7XPw3ccXhbLkL0ZcXXJbRRv03u2s0G9mKDD2PA
gr+4RCvgxvdJevQ8TvyJ9RazuWyrwkZXQ9y6uV1YlaTcvJXmdHkcqRJYWtXC
GcWOfjDNFWnX6FN1WOC3Xd67wA80aKg34DRD/16zLoDgYcXt8PtCUZVS1AGk
ny8ZW3nZe+ix1rPDrCu9w7HTdtuInVddd+B24+f4uZTfyoJBm+hxv9UC1K4w
x65RgvugQcT3EDvbAjubP+QqNeC7wNGOUeUHm7UUm0XD+p/zzFoL+Q3I5S3X
qc3p/aHoJRwztnV42cNiwKH0iHuJpaOYVni/xRjVHGGPUUgDj4JvVNCFo5zh
fdMmq0gGv67Yc4/yrnTNYYrP9p/VU4o0Gl//WGG2fLAq6D5nNuvz0X76EGpN
3PxJhLjms6Az8+LQdTxdyukIEWeBqYXuwXP71tENJ4Mcvo0/gQD+qgJARF7+
x15a376pruY3OyzIsMJfdtpkgm2SNEtlsq9HIJ7oIKVqR/42D1T3zouxX5ff
Eua+U20j/2Mr0zpkUDw9zFSWKOuMUlmnf83NmLvtx2+zvbAWRYkrMF8OfVE/
ir4VpQWg0TDs5tmsWOu2OQLU1B7fQjGsC2Cq7sTMJSBBUVdb0weWf6mifBwu
OSTZHB2K5Fv2IoHbW+jGUKhpobr06WBiDNU9gtL8rKuDtsyuEs9cAZRCULra
WKW6VvOsUujzQ69gUXaSC39NbWHDikYNhUiTrKJ3kg/hSy4ZXGA5s0EnbVK5
kJcji4Z0Mfz225g2gH3VEmg1K7pZpngllNA3LrwUAyEYZDpTcHNE38r7bvJc
g13Wvw7OF19UJSxngzuFsqlrCGV6YS0d+N50cTIgTJuwDhDBPbLMaVXORNO9
QYDXif5YW0WoNAXEYIny82CaLpnZkkvCzTnm2GHAP9EY16krUlit4r81GIQc
Ff6N+zvZQ4wr68E3LjZjS6SGYWc0lZeHdn8jgbKh0hwhm/ponmp73DPzsyTy
79UWRFPmdkjW2z4FOrsGL6hYtzXUBDCvgKiWWi73159TCFDOAeMwZI6ZvIrx
QaptArsUa2GyVUtbAVaeoAdBze3VmHbFbXTlFjCwkN804NHNHJRc4t8idyEf
Baii2KtRatkb+bM35XnzByeCvNbhV/XMdRKHzB8fsNYaZZtuEvxxR/tTWbJ1
ksz2sL7w6M/sXZjtxJlvufO7gtYdXZEsPXdG8b6PVjUrzLqlXQkc1m/6T7V5
qbkmCTSouABRlOWVk+WvLTqItS1pOxeuAZ0XuKEn7jUloY01fPUjHqtIDIhV
KM8Be2/gHYQr58kAU73JfUls7ToA/LxpiovH5o+VD6sgidWW2cMKW4JljJzJ
wuuZDIQeMsCniU03FsJjPAqaZfOEjku7sxqxUqJC9psNXn0eB/HomJltk350
kX8HjWJ8qX+cICYQsOnNtT5S1WLL6O2D9khgaQ9P6KbIqmPctCXHe3U2SUjj
yqlr+/fo2+ronvX7EVseKlfeQUEzJf0wDHiTSodCEyE7IUtclJeBrz63k9Rw
JNdMB6Di1An8o12YGx4T7O1xSJbASErCGtya5bLshpOfDC7D7T1iPMmvGZon
Pph0d0zbXmCUGpL18iawUyeJCgXysMC/iXdYOcZbALMuaqfa9evJc1DJu7Ej
ZSnlAzw8b5j2Eko1Omfh+GPXOg/iDN06hfFKwfIYgus5vTPL4D1Lx8qCD+RY
h2vMu5FdFJmPAV3hW7OnyzuF5UmoUjVApm60Eg3n+aNrDue+XfLzPBLJZNnF
HNKyKnENUyuJGv3aOVEqIKdNk4gJHIpey0nA5ELnHGsowAHXuVnmZrg18TCb
C4qnAFQquwnwdkIKydqlfIlRlx83Xoy7JcFvBz7DeXEa0cGRzYeyeb3Niq8Q
gpvKhIYGh88ROtXCo3pmiKEdXk3RKCJKIVF1H455b+m7gnV01GB2BNhVNY1z
XKnATPclXYlUHvRFQQXK6v89pYOSsGxpN61BwhHHM8lwP8+bS31CAS28J++R
w+NvcOpvoSR8nsaEsB/p3o+yAs0PJEnX0Pgl1S4PVL3+lTYhiNgpACn7wd81
gsxG29jvTwx1hoFhr63rTBYLdML3h9PZNNhCa6sCUyvRLzQYw/7qi8Bnfgv/
va7fBkChaG3Q+0zDJJK+vU/kiruAzesXyS+atluoPAf+vlRfZ+TcnZSd2Nhn
q5e6NV8pfmo0jFz6BmEpCWxbFEEJQKHt2toBbVsZiDJnAx0Mxe5XEteo3PqC
TlRE6vrS06IYATVF5zvYeYKCjpxZNSYGUb00erfsbJgU93Rdo1/+poMiQcN7
maRZHLpJZZ+u0wb6GQY5sj5IGIY2IUAzU7Utu1Zhj1Cwps9mTDvBZsfcH+ob
1fEvbhdWqSh8elADjHno0765PnAKDqTexivgq1VdlRzqNUdLsyo4dWOJji9J
B9baq96FkkQc5wFV5GXo0YE7KnAm/x7bBLRFGkew161NVC8LNhw6MKa9omnP
PRat9juQrkEmEyoMbNnMW/yd+4szhPFcrJSs2FIdtWsxvsuBqzPetrEWJbKV
6fffzrqfomEeEZbp/XyRdyEgpBwLxhCkG+BbE9vOSetdvJODQeXlsvP/+PPP
hbPr7+Nr7ZhNQMiFpVv5ON2dZ8VCY2ADFUf3mahScHXpIK+SAAbSFpJ0UesQ
ShB/zmjZnXQU37oS5u9ZgcZUmCMTsjtfypV4ZaCXXS7kD2W4GA7AvmiheeTL
X6PTWiAERhfEg2w5uxrWi0J8+Nk3y3yA80JgCMstJBP5ThDK24Oj1NbE7vzS
Fmobv/Sdz98EJensHaGi0mOF3mOLYxfM97N6HHCduvZZcT3akXrnO5AMcK32
Xt9+BRB4xVLpjycQJ+QSeu9WSUtxLgEgceAST/FGygBk4seRhw4MybuyLaGD
Fm8vvBggv01BXmUzo6DwBEE9PPkBiSt7cdDiKpfMvvp4PvdMahYYxvW0CT2V
/M29UgJ58P19ErAFstZiUjPElUbgK73OdCUfcGOzJixHdaE7fxTM+/YdhH9R
vN0hh6PHT4BcL4DdrmSPaCkblK4HJL6r6g1JrRLzPBp4McuxW2u+if1RBXLK
/xlrcsBv4kkIizjQtG2nMMIx9LXWVfVOBhwIsJDfxF9qY3ilnIyx019YxY+Q
ewsz2Aw0xvPcLt4jrEHMNzyYjMAF8wtJRIBZMw3EQfB+nWTMifFTDMjYxOrt
WwlLDbD96v+DoALhmBhYBq13usJmZ0kq+VHwWUDtwEeLE8fryg7RodFSyep5
Lodrf9eTLzAbMQ4pGv1fHP8JHblnSLa7S43OhIR0oyovaXlqMM73MzJ/Iuvr
KDQ4yffFcqnG0ndMiDaITRy/Y3FWsU4JiY/G5UIGYauNHIZjOtcM3lQfM9wW
lAJewWkyQXtqBrutvUQ0vMRSFbiAbI01LYYFkZXAdT/tAQ1/+OVRAzft2hL4
GC+EhqL+s6B1b6jpo6lskpUcwpBFdgc0pwQ0OyeE2kwcQz7+YwIm7VXyz+8D
n4okdtQuIFyF8+FzoMFSHo+UxcAA+yLAUAjBK986FTGFGu/HLtSWABm9vYBE
zbi0e921C/CP/iUXGvOmZ8y9b7O5IkPsT1IMpsPv2LWlpXLt38+VnmleYEUZ
SyMCmhjmPBJBbNaQPxQK+zXuftl6Elcr8TczVGyUPZW4a0uIEr3/h8o+2nxm
HSCFCGJ7IH/juxansbHwdizKid2cPtwaz5O1LKKmyJ16X4vOZ2VCq1tuzPEW
NZNGBplBL4wv4z0X7TYCLyuaEc7N7izsgSeHfnVAE3JhW8Z6zkB3WUCHzZ3V
JLXlz4uEuvbonfmPpA7VE8s0KarOF1JUyhtvJ/riT837FWhpJowvGtqdNAYc
X9AYEIeZC885ONS99R35+yhvYldKDpofyNCNzqxD7haM3R0chx5h9WPlHzWw
fZzEMBkQbmSLikYnmnyLeRSM4eaCpbPeZ2GywnlXaU1fsCAwZ1WpJmfglp+T
0t+s7SmJ9LrF8aJTSakIlTHIYdf6dDaVup+VTBsLJltRV4SOFIia3Zg5ktbm
d+/e5/KNOuyCiQ4MmaoWKpX2KJonwiIUIkoHa5Bl5sNAPnSvUQTGxngDmQ++
FDjkIl7XX1Sro25S3Fvm3mnIsYdi8+5gcPKvWObeOODf6k44L3kiggWrzblt
o685pSjoja/AC3ncCBb75HrxJv+jpF6Dx9wSPChNIAOD/QB1UoR45zVqjPXv
rioeAEBEZkNLg0+urKS/mCtHz1ZXsF61Vgcm6dfJJmq5vL08BrDdcKrjfOXt
2xUdnAttJOnTxk2qWdwb5bzgs1c29lIwSXpU38vmeMEgswk+nUZz6eaLEiLP
FxCurj/+lsOtNp77aZ8COrmHGav5I9hZwNMreq3sMb7fT8QIyE5RBZgHjAtA
mYs/gXRgitzXWisbuhvgALOh+jhe9wwLMGZnXR0CuLWwn40WYZwSTRvLz5IN
NO8jtulQ4B9r9BKmWGGHl4VQ4/aIUi6bXZ3do8dowFKDQWp2Spqz8PrjSLG/
YRL5OVgvKxG8koS/4u1S53NsU98zVCsgt0WzmQesovSB3W3QXH290qEx5oPc
RlDn0QRuMzixv27Kb/3bxDNlMJCIiSnbkl6PdpLosbibYRTqMOIOGzYbtcGk
Ehj0uscNMdKWAG0YHWIsvtIhgORV3OnAnpazekb8ek/TVdH4A1ITyKh/cT/y
ZokWO4JIMl6jMuLuOn4ypyT7D11/JYfxezKxLBVhtMbTaAJuewQvaVeQ1Lf1
EZtUqBkSRsVzljE/cwxT7KWST5DMyVSPTfVsOYfxN9U986hu7VGlXq+bSARv
h6P8DiKwgubTDfs+UYLyPmbuJemKGQO08wm+HEmerq3cx8K38u3bgxaSHfKN
N0D3Mv/tLk2tnHVhOQe7KM0VYWgQGHddRaPaCxNR8L+Yrrhrog7E3+muUEDT
rIeZyH0ACBDA29vGRBlFIsPFNoz6HxKKzld4JYMQGpiLpdijpeJlSG9wt0oH
/oY5u76pqtxOu7Q+w24hRCjilj08d1A3IJag3Y1Pf947GOrYWiA3qhub0O1C
6HARdCFGWGi2VL5hylk6ChS4diZ2LNsXYjia+NtOEp4/QBOllyRYEM9hjijX
XnEaF9mxuW1DvAIYZal6ZSjlZjfNCozqOFN+3S0omuwxF5A326ytiIr/+Huv
kTN3r/89hzu8r0HC1fftwftPJg4GHGWYt+mqqE9Qh7+ANybAGLbSLob5Z5Dr
f9JI4y3/Pticryw4lgv048N4AzBKs/hDZY46afpA17RVXUYD4EwgxJWDpHkm
3Ya/JsnWZ6fIENSLo71/we5ygLq0qNRp7oUyMjpX4+8b4TtdRERQVMdmrdcH
IDqgxb8b/kUcV96QaUwBugsMkZJr4bZGJfKwaY6rk5Krr97BjYD9WpGVRpDO
CPGcv6Oi0M9NUXQDmj2jSvGxWMjrhro/QzwASs13ilZh8QdAvwJfk/oXSJiM
sThYtbp+HZ8XPPqrEqtCVH4wpkihLa7zvZbptR7US8HOv2Uoh6C6RlMYuDST
a8AycdxtiQQYs1iwkC+D82i9dUIBtSDh9soznuhbxEGMAuYBNhSjDoeqq0Zz
uErVwMxAO0jDcjpmWZQcWCxV2wP8KbPNSToRVCNFYRXCXCBKGnEmj+9q6t+F
hQyRTMYgobAn07/yAenrr37BEfy8f1Zam4zNzCc9r1PSgSLNlV9pdaUZAyJI
jZJtadvyttGuHL8HUppKLSc8fODgeRY1IEPtx9x+ddfZMzS77V4RqiS4jQsX
iUVaW6jsXdqJciAs/pyE8UVon0ScuIaqPXdPNcy784NGRaSi9olBDoyQDJfQ
vw6dKVZD1ygOrtwZla2laaWjse7Bymm14NM1UM9ScRhQyfqh4IwYp6MxllTX
KOdvVlSarVv5Ugl607kB+5YjX44i3mHd84VAft18zcjTU/kUWpDO6BD/WIHn
OQ91A6A++934OKuLvuKAXoNmyM4gGG9rnK4JyQ9Tqd9LgmL/AZJxJQPumNNt
gBzsRRxCljSPvYAd6uF8sq75UdObz+VOj2i07M34vYhgowTwksfUvTbMQSYN
DsRhdhTqazgq92QnTFN/fyx2+9MRBRK/3rrHCeVy1mMInXDSktzMy3WjaUw0
VxpUIL/WY0uyISov7LLLvC8MOTQ2ba76KLfuJkq65klA1yr9fokZqxNggYzH
/T6Sqf8EeQtvB7LiB0i/IvzHB3s7KjyAURPThNUobF3iGOdrNZyV3zh3YrZL
iwlfVOPuzhyCygZ7UuvKCZAnuXSSUVSpvoi+csG+dMO92eTS+pZTz3sgGmMn
mIkPsVgHmXdyjfUjlXuLS7nHzZRfpY+PvfMA0U1SS8G5JFG998/y9/payn8X
pDtP4JAgegng+2qzKoPuGmk899amoEt0jLnSBxKL6MCdSzegbzNX/y9sfCwX
pqlaWew9LiqKvvR+xy0WB76f2dP/hvNeG0RQPWUs3bBXiwkIgpzI8Hs8Eb0e
WZK5Bb2aOuUUjtXqGGka52f42a/WcI/QOeyMW1EUSdE1q2Le/RbmrAiOK1vB
NfXOjTo+EqAkYW7YRIb8rq9Feo4hp+P9nXIjg+/M1dMvK0Cks6wjWtgMG0Le
uo6uUQZ2Ijhgp63SntjS81vP/D4IJ8fduGQNlyHu6iSaL7x2s7XczN/Yv0Fn
2330NVbLfcNHtwGSSUktSF6sMTjcjfQjEkXH1RFXaBZKMIpta9SgrAGeXlat
3kWBsJff+bStC706w33Me49dU77alJWoZrfgKWbmfi13UZOFC1NsuYMgty48
G8N3hZWi8TvWyMyFXJHaYNlMVrLCtFBHdY/GPXisx49RnnEzZ7MrfsIh3xFS
GgWO2JNswPXfAAWvFtpAjVe0U07xLLJK+A1LAdNo5tpYENP8UkzLtyh38v1E
Io637cWfsId2Q+AAgJiTuj8HYzNDtNXh0HH0sIfqdQfVM4JffRAJWZltxEiR
BfpOYRTMG8GCG84AmKvC5cc1OLYoudtuOtoF0MkB05M3QxYp8nkKpY07KETq
21OlScPVk4cXBsFtR0/7Vyqo5GcsKzWHPd0nFjvQw7kJ1nFAj/4/5brdDMwZ
+OnmA35kTB6TggTij3ZUVkAbK8vBPOvUXIvZD9bNIKe+N09TbykRNqAN9Xbe
GHb6QWvALttcC28wleJAGpIIunRGzSDmfromZHCrstOrQi5nonat0S9u54XA
AOlxcH9ScOStFSqYGnEAGBYyo5iJmErmd18pC6FN2CS0xTduATLxrUVc3SIP
9oppPNIWYMIMyOzjXvAw2duHf9CNr0ImYe95xySnr44UDKPM5K+lkjpwLhFm
+RZhy8llC7asAhhRDtoGmQqO5wog15PWLqpz7MWU53dd2ozctu2jAb2NQTHE
N3RhI+Bc3WwdIg9Y1b2a45jOK5+zEj7mWd1Nx83r2LW6IOOpcYxDqd/0lGoK
0yor4oTEcKLo9J1GkW2UskzdgNVbdwenIkonZHTQLG/5h7nNWIkx+1g5MdZ5
HSgMQeOF7afSG6e1URNFI3Jq1IAMPeqxVMDT1FaF2+gZvqVNiJDgXJ+UIaU/
BvkTiLm7UHWxEEWCDFlT8WoChisM+iNbH1WfmoWtj9VQiIEkV6/LV/2oS31e
Nz+rB3TIvJkT8IUacoFMop/i3AODu2+fIv0hj/RFROrQ02mgEwbgwaFtZ4J4
BQHvO8Ax1ErpR37ykj3ZD4IESPRr0FlRssQgwMYcJarFm/75iCeu6Owp1pgI
aqYcDWzdwvySANQu1qk7kKYNExwtBzaqA11lui/OWKYmIFN6zFaCUQDHIAFs
2gT2/FeQEYvEeXnNBzap2Tx63okhuxJesT0oC8eztWtsOTrpQIeHyH8QZpIC
4ax5z9dj0Vdh+iW3d8OdwwcZz3TJ+G3cW5Gd9Ql3vf0fo6k1WgPnbP5kFKWn
EFG9HdiIW8LqiIczACuod/oMxSgv7rhLd+tCuNU8y0bcA0Rn4cMANSUN1fyx
rNeYHxGE5GjDnzqOI3zt5mMo3Cfv4AfVjktoenM9pHhtGtvzhLIVmkcRkPJ4
2e8uyDrfvtSvCjzKBXSN5eg2G4y92lMaE/R82bPHW8wuPzro+vB0sgqDmlUQ
mckdN9HKA8D7ULdnkSA6JHtLl2cYHeR39cRhKBafDGiWDIQ73ZkSd37/81ci
LcAd/XaFEQtqsmAj4aEm9LVSRsmd+n2kiaoGtGjIyixkxwDYgj9YH9UNdQzs
Qrl9PDPJVB4Ba/Umf7rFNu84ZlJMck/1NQvi0AHKkne3LdsqbjzN748CJTz+
be2N67afpS/gjcbPmGcUJV/cZNs0CEs/B2wwtqJbBoEP3M9Wy1m5PySJWPBe
PGvR+xRAEo65tMH+EgF+fJ/x+XqiP1Cl9jp6Tyk0zwf4UjhCHLDWZWZ6eaum
129RzNPOYvNqep3hfGCRNW4B6lpQNn3NW8xwCOCS+d2dTPLDXdr2CgvlQjMa
2o3X+0fg/B8huLEndyzvl7+Lu+QHwHMnfTZItX3bJD5nU9Rte9DMMsadOyVY
+njlWH3h0ZxOd1vIeR0GUfYwLeKH9+YAXdrSx/7i2CkLrskgwtyCUcymOAkn
zi/nnGvY35IcMPW9VyMlPTzYYWtdJVJFD1kLqc9OWEaLED9AQ3s38P7vl6dL
7XLU/fKuGtlfAcmyIqTSasnKND5B8hGl81tc4tovYIDknCFOqh5cR706u9IN
FQyUy7zyBtLeIkeVuwkIUvepmL5+rtQoCjURTPSTjGiTirImOX5N0hCoSrYP
dvbo+VVxbNtJbbypnGJVYP6MeqpZVAX+jNRnR9o+gMc7pcSi4plcPSCahnJ9
258JjShUXwa2YCgXeI7+TNnwZh+gy15ktodILJvGn0wuzbXsvoqWY7ItFpy3
jxwJyu4+NsgQTiOJnUZ0zKv4OflDrcaeoHlxqLGIEd+XfWJIZe7TGKb3EcWT
qjfNXcnT8e/e1A19G8Kzyf/WloU9oyVJT2nCzR+B/qDbwCA32W/vIF3LGAKl
OdYrg4EoGoDbuxOGOd62cPyPr41bWcqlyGCS6fJ4vjwqjQp3LxRmD9DwXmWF
q9YX2WIlM4FooMYzezSkslu4gQk2DKwAf3F3prsnnOwyU2jwNri66RHHmcBB
Rn0Woe9LpCDAQw/SyI71x29oRaUV8s/+T5hhH/KZpv2BR2atAK+5klCrUF/U
AH45IntwaRmYb0gs/gCTJ5utrzPfiqb/kvMW9L+k5chCdIDFBZHCcI2MmPBS
XV9weqbMDxHHftAsOvYWmhfnoaQPlfVy0xa4xPkqTXFRknrV01CX4wsvi4Rv
3UXgr9HJ77/6RQ77UM+HfRSRVq84/NgOkJwTgZ7cR1Q9Sh3Xq2dSD3hWUM5L
DcgWsmFLVyxRa6ZKqbuFovgFK0d+vq9/t1ZLWG3cfZiPb7TDYRHL5rdspLjc
Lj8Jf79T7xBpwXflUm1W8P6THtYbXPHjBXcY0zH+Ldl4Ck42vq7Xx0HZaab+
TzVLjZn+3PoQEiRNBC2Xd7x4OwA4yqP4FFkEMOpzwa+p1IlK8cZ4TbKhAJlH
UbQV37fEjFvu7pSe+DO2VyLMRSqbbkWR5x65UjrqyrZwRKg/QcnkTZGuw9ON
gJcKVnF9qDH1fDG/dX3yBprVYkki9j7ZZAmsjd7pBjATevZ+uGKomSoHtCeg
SQLeukLRwL09OnmJkfxkCG1THZAdGvSPgt2+fOfhyvLd8B4zs8V+NTWJ9uYl
9Y0G20ze/qvgQTsrF7bM/0bEMGHJO5fpW8AhkG5A5lB2YAwmb6Z8MU/xkV5n
xvIPxQHyqZeO2MLz31U04r8D7MeUnexVEXu3B6IW1VkI5BVZosfRE5yHPJ/M
2+cH1aJfACV2Np+f4u05Iiq/9loeJhOFSO8mEqmb3I9wzn0bTrIlWxqiKDLo
TlWjGtGzgl/ggBkCEQ5ezuEFj+570u8MTCK0wzA/SINtAJmxSRDZNY3u6CgK
lY5eWQSUkmSFDW+DzAs1LTazxI0XDZeRraYulet8lI/NlKfUj/3G51dmdj+m
Aiv8R8Ff290+Q4ezzgYAH698nrTQN+t8HzWae1dXqgHPSYEA1+CyFF6bdXUB
IrHLW7lULxfhdArW9v0Gx+6SeKwhGTEdIrMW48RLVzoy+RcvK8YivN6NsHCr
+sPYSq8/zSh6uOg9gwOpxFRge597F8xggJdIEPiwckm0Sl685HUeQr5vz+oN
D0TZiBgXAUSw6E98NzRn2byenGFwcFdxjK/VbsvNIe9hyduKTelm8kMXauUC
Qt8RvhdaPYVgZRgVxTiHfOaS2Sai7rQO9T8XXZIifmNddJsWKmayFhjanYVo
UWkXVbIY8SwbDu/YQkfFEOwwCje1bueufBSkDOVCpjBIoNwAGnaoc2BQku/2
DGSGnh0/aRCEztoPpR2lo/bUo7mSSbGrsZkAUZ0KiAGPQAJkHlUwSJXjXNyU
pbIqGcBRW9uFLwTwejIVeRreNkBkQbadhz9azEvrrGf4JrDSwHrOjWqqxEvJ
dQOhcgotSLH9XAZa+sPkv2k3VlRk7twkF7R34vQowyD/dv3T6vVBKF4HCStB
anppt8pHw2uDxotjs+c8a/gFbpvdxRc7/zjOeDhWiPkUYVHyXtypUVrLwiT8
OTZKYFnkEnpScQftYz1UGlRge+xK+ioAAPr7w1vRCIlCsGREX0iFO2lZrgsb
fN9CRtFIgHh21Rkq/dhxL9bQnnk86ON54qrSPO//447wN5Q2CZjHifYt65Qq
ouiNAAFxts/nqCBoVK3Di23pc97xPdFLX1UHgABBJwAKlSF2OUhmMT7D1y4u
ohWa1WjlGIVVs/QzEkTm3uekdhJCPeNZSvGAMqv/28NF7zWRuR3FBLIW1p20
xT3hjGr1QGRIu8rfxhKJ2qt7I+O+1P0xf4MY9Jn8aV0ENNOYi5mZL8PIo3ZO
LRWHLhlTGrhwKBFK34HVbuzt9lsuU6E9G89rMZpiGCFevhGbfPDb6R5G2LZ2
RaR83HWgNHsudiAiwA4MutCxLBCA3frS16k45+Sx1W3NsBJA1+GaRTVQzrrf
G7i25MTiqryzOzbxeAwni1pNDPkLRnkNQejOVR9yVo8rf7cVAu1fa1CsiC2V
CVZraekG51TYdPgi92e1NUohRdBV+AuUM7w0hbOLqjmSS/uVcZMW1YGcVHKt
+/rMPDcC9z/RJWDFjGLZ/g1Zq08HKTV3iOnVw5qooBimsfYpAQWDupFFFxjl
3Q8S81+XuybAc2LmNvUa6viQxNrwL5fn8NH8OdEXka8Sowaqjoj9186wVjHz
naO6msV1F8Q6aHqqlZ1EtSxnQueGzr0IaaZZ+fmtPNozleshxjXgh41moIU0
VV5zRcBgKklnr16QUjP/fNebaJc3xNWQ1oZLUUaBHmfbrJUZeX5CohBsUmcd
MqCg9MFZhED6Ht0tCUNdCxfBUE8dXP1I2hbaoWnVb9EyWKvl+woSx5jdcjzV
Rcwgflg5bXbkKKAjhM4ECertzbQdUD2UzRATwWpjygAQWMa0pXx58XpR8D64
t0mG6YGAKZNmvTthil1zOoka40ad4dbVjG2gm5iFcROPsm087WnN0QltblVk
dIHdEWZb4ZSlve6mXE5F7SOQlNsCPBf047X0gBzKw7mOqq3UyyOAPTSOHusM
2kQKkkveJov0rMWtxfz9iLDX3M6rcalNVMQT8CQG66odL+jUsGWXJiL7dBV/
M0M0bvMWmHPK3Z3l8ul7vwaL4LWd3yl4FWEO/mHQnb+uR2Bx1/zUxrRPExFf
jFwP4MB3U0hClXnK3kVo1e24OsmbJYsZVTKu2oQp/sixpXM3rgsUNdxf2q7U
KFT/ZciP+Ip7WkY/Jle10/XCOCVKIsKZ+k07FN1t4IAklEpd63IpaflZ6cT5
FZ4aoEc+M/sEulGQcALuUSgNSUsifjCN42xADvWq9sYAGJ2AiVwq2HTV92j7
okG+kjrFkXbgQSS1Q6hpxHqjzq9N77T+ahrF5tpooEoz1WdI5BVshrMkiad/
eivgJkqE1mxMEUry9sCTr6KCx64a+VbAlfr9NqQJfRUrZnUAJuZMPL5f4RfL
+jAbakU6jf4BAPP6KwNbxd34NgCtJ3DxUkYTAToBqfyjsFlS2ml0kJjoGJeb
AFBucfASMT0yLshpPmHv/dcS8lq3LH8iNVMMJyKRMk2nx9HnUg/pGkWMvpm7
S6u5ppjvTncdxfwWZXpAogp2pV2Dl8O0r1bcKodMN1Oes2+58JjWOR4M/a8t
0RQVDSesjVbZRaPsTCuTMmBa3Gipd/JoC9zbdvK0k8Ww4Y9aWF1izRovcXh7
U5f0KPZVBkI5QScUT+eZFX1HBjjKNfyELMYPjImJRA/ShTTya6/QQfU1gFCn
/p1OszqJZ2rNaSFLq2kO4td8h8nQNf+CsW77EoiZQVZRC8EF3uL4J56z/luV
pZp4O/Jvrs2kNl3YXaJDbt7TPRWVVaI6OBhffSQ/e11GJB5mnpxryNBH7TKa
kwm14m2EEVN/dIvVt4AsncszEDUIlMC69Lpdx9gTm6Bz3+cmhBv0qxqn1jS1
0hv2W83QC4QE6UDyyIw109Gl7lqZbfLvVsHDypzLaD00aCcQcHXlrfZZWph4
AdDZ6G7jpfEjFavye7Y64+LWO9Wl+7+OrDUAVLe4x2RgrBx50DGRBDj2pqkZ
Nd7g3/AlEEvIMgNZkuZl5y0aqVSmd3iDSN0NHykehWH+aKrV8CW3AJTIaFCy
ntKfw30mCuc5OFs8sN7J9w8ad3H8w1u2ZsYrIoOlOEWLt1C6us1l27PcdDyY
AXG+addqsSre+qa1whQAFIEeKsFeNGo5uvAiwpnOJrdC9VK7kvDVaA17nYlt
FZJJNl+Us4TsPRI5OTe+jfkzbixn28KPBnM8vMaejfRfW4keif+F92hpEk4P
e/rOCmEWY5msfwIrH5pbxr09W6wDaQawHkLoBZcbu++b17tJMxnOj5Tgf4cj
deO44DrqUfDHoaSxhUWfqxjvwEAtYQlYhDqd7cm0/hc5h1J4O+k1vzmDUOn2
oc7vyxDKYUppfGpqjkrtPFcJbOmmVAwEnWT4ytqWy6M08pwd6Du8z+8kVIJe
qgm3vIH96danDkrxvJ9fXE49Js8j8Qcl0iSt1a29Kh4vkeJjbhGKuD8mWkAf
qhGJ4YLBTctbRRFrkDw/Ic4BKAH7pQKEx1ZWpN1tuVVd3fB68IqP+sR7EgSG
LktkWm+bk38nrmcymofE/tRSiHgiNigtkyzPQ9Y2auX8Yp7eJryRPlo6wtyl
jMOfASFLyviXLp6o/5X6AMUSjKfm5wRYoQS/KzYTlII2Y4OWPKUeUZ7CATLr
BjaC54n2AkzM2SR9FCuMr8dh8FvyFSNPCeRoIK3uVxnDa3azEe5CRj/cE7HQ
Y+WAmzK8OKPVf6sesWPKgpM2MZwo6E479fRcr6bvd/K9ojbptqtEz6pnJpff
qgLAB4l9eJOxZYaPW/Efm8FNG1HNKh7gDS8WzNJQ2NYzyU6YClR5jtDfIaaq
8beSMjPpB5QSl0b2367BEEmrc5xSgmLjlhL9DtTAZA4MWSRr8v6Ees6AlMUO
0Q08rV9j6MqEyvW/hPIy0yHDlpBZf7VpheWcd8VjiKZ3G+O6Qfe1ohsVx/QQ
ZEocg2pdNvgpKbY7Kl2yOkeni+kWvDDHbAkUDPNoZiKmr1M7Xdrf3n2CP1FR
J4J9EZxg3UZMPyUQLLjr0QpJ24FFaL+zG5aD4VYRo6GOZrL9Nk/+gT4oNDOb
eSw7zAKa6zRHOclv2TNy/SW5EMNVZnsvWwnPtFIbYRBntSJl+Ink5TaUeizr
QK9Os7IvtT1ybk1xHZXfxTin37mqiEWFT8xKBwh3gH1lcJuEBprtpZfi5ha8
wRvw2T4kh1ewnIVN20CPIbs7TdKgIkdKFtRk+E91AL1xfH2kJp095WWPo8/x
hw5y9xzX0dQgO9NcnKlc5XsshcA3nygw861ar+i8B8YHckZ30+SmTYXIn5S2
DV+Nk50Juc9DCQARUdBIMgeIVIWHsH0UNV9LLnI+e+KKVurJSrnb6W3mP3X+
t67CwYpGbzYoyZwyEAsLpH/ttI2SBXJJARp1ZS2J3qoKRZMbD/vOPaUbOdVQ
LE4xU6eFd94mfAGDL4YILLF/ZIROnymXzrZ4+pjc2sL624IYDMAC43azWWaX
C6GPm70Fp8hQKGayMq+dsLYXoUDI/MCmKg8Ci852Czsved93HbOhr2R8X3p3
7w9kn9KuudCXHk8Q+0mzPkf+eByE8e15zn+ODNMDSyTBii+el1aFqfy34NPS
y4p2RyyN44PNRsnwOANkAhFxe0AXwSIZP46PQtOnjHKxNapJJGh6ufddx95+
843FkzSihJ998JlFwAMeLt412vB2UAtrxubXtLzE6/QPsR8x+prvg8TztMlm
tig91LUEHV9XsVyAqhS76BW127W2RzrQABHHajBdPgZi6IWdvnJwoOGgrDvA
d0sX8dTKXk/ald5hKplh0xspXVK2J4gortnfIhHVc1WedAuEGStGvvj1J9+7
0eHFhGMYYRiJ2gZaHLo5aTTj6mTgdNQxrVTn/H7IhQ5XSNeuKPsmm/1jqB4T
MMKbGZSf+0YARMVyFXq++xsx5s3QtTZQLK1bddms6Lbx1yTdIe8KSIB15I5x
WHw5BDgCtV3+6gcQsa5bDhPHfD7jNIn8BhUOvn+JS+QfzipCZUTtvL85iFqg
FQy/Pvv3dk8A34ipZoJmBfgjzG0LkLj6HrjedWIkmXTMraUlBZVeHkGLuax2
TAiHM4EwHQNNLw6R1praOh6S096I82/+T60404Tu8z5/EKdMeNFNB8h+YKj0
npZaur5oZRKUFOgxakp8/h0KaBcNmyb8/BLwuWtx/nKGJPeNjuQQ3SZIWhcE
eplNMX62y23NeM7BnPwt5xkqq0n2M2NUpYvPFjXV7Bm++42bLIZTxAW8Pvhx
Mfpb17mLYSsc5Okn9B0KoCAj4w+j9p8NA/uAp9a+b98MKLLH/x5mwhxt0Ix2
TwIRUFZn3fSv593Hg1mNuyvXYkYMQkq725pf/YBWcQbXpPivipevBIU2QrmX
i5B1zQupp5Mv9HPJEO6yblRzLJC9aOxy6rZUZq1BpPMSf63ioabZ5ygX94z7
1a23xt/lEBYcmKwmzJXKMqrgaR7K7Q6nY6Gokcxd8Fj6YBLHUl3yznDJxpYQ
L+Q3MOyEnmIJqH/KLiI9MW5ogYD9fZENuYRz1oMxN37FK7HPP8p4LeOluUe0
SuWMUPwfEQK2EauJJcsSvBLwz7MbENPEkGSmkgA5H4DXrrnNTZxYNBXoA8Jw
54/dw2AmTyB7cJsdJUDUZ+pWP41mi7TUIKMrbhxklwFX/FvD5BOKnKtX38Md
40l61XQGWaQHTlned4pkJo6HHt6d9cgIWfTuM4pa9XSL+NhKL0ZmSnb3URwM
0UKcXzLb9CofzJE9YTizrAUQCSDIIJP6unKYbfqBdhmnrkVPOEIOUnd34xdZ
5OucgdupoZ3LVAP5G6BW3J02KpDtQ5LU6BPCp2NnAdm2YPFazR8+FBcu+6Cu
A7ep8YEMrtAYN0NkhxX+BLOyQHDDP/w41Mzjq9QwZIBhWTZKAm8s8osGU+/r
uBB9T2FXo8na201FmN1zNfRs/9t7iCssXwmgUlxRWvvNtZrdRHinmi57RzaI
9L1EXcx29guaF7DkYXzQQEsFfUJClKgo3gB9aEbBualEhyJBQ+llEUfHzrM/
BkPiVn5l22SAItSlZDcxGCGAG54K11kt3uITQ7fvDKjYT19DKWW0eKPdUfod
JNcM2uaztsCJLGheNmvR+WeWh4xh3kPSQXlBQkNltb0z4lHvMn1skmI5BKz/
BDZeR8wSAjcQ/4KFf9MboBPfGd1QpNpDKMSpB9W97O6p82q9YUYcgyH+PoqF
Yv6hSKnHfFvwtfuoxX0FLbMQ91EN14mxvTonBbhVFvF8U6tO/WxAOHkXejZa
Z6UolDavxzbHUUkFDeW8/2kAZeiwnRwtDm1rSrDQfTvejIXA3uW1aqtpgBNt
TM5lo7kA0Jg2T+PZRXd47uEmGi7dkPyFfZcZWjbgMTqO4fT3eZ9LtNcOFrSe
U9pysqusa3yv0QyBDhbyB06laNDeyWvKEMjBWCr5Vz6Ai6kM3e0iRM5qnSMl
e2gUGDtYiyC0WaUXI0JSoY6hsKF/zU3sDD0DnH0FISC6o65TG1u3cSapOB5W
xOhnkN4049WLkQE+UVMinxWVJJC4TnlwEwXBHIFe+RvA+njEbpZybklHYDg0
EtGQ6a9ykb9NYh7wE87qeAFi5HBZpAlwxfDJ5saWEdlBBFuXw75xX3h35Cai
SgSTn+opAYiJ1YWlAGJ66stdJJ8WgdFa3eY5l4myT7AQkYo6iN03qSVs//y6
i+j/KaDVLzlAGlaQ84X2Btw7npn7a4bPLROywAp/UQVt9FzITcIGq0CYfgxz
xl7PqgJECVAX/Kz1yfmrdfSvBga53KW3pcbD9d5v2aTHEHpu5QFrYgdfpjyQ
Ah9xGKVG6c2NpT/OVWeIMmVtWDLKJfjZQUkSklVRoo4wfsvwNsPSxgmWdmoc
Gp4E/TB00ikZARG58/wIwyTvV4jzSDZeSQxpYC8MsCmUmALduPYUw6RSIH/l
Top9BMcFJGLmzEE8/9vMoHgsT3iaWRQ/EHU6iAbtDw337lFxcUID6UgKeCJJ
6M+h86zXujyvlx9MS+qFuXuKQpgKJ6XYQcskLpx75MAzq6JLQs/pDxU9y+Hh
orz4VysCxkPV5WBJD+y5gtZMvC3INN7Mp9Lfu+v3kaNMkXNqmJ5FthPqMap7
lf2Ee4TTwcT84RdqF57M3nxsohf1KnPhKwkhHEmvu5et/cmgXW60NS0rFkmi
hkxJkfyssM1QgBIbdXPWsk/dXfKC2pZ42ScobE0ug7JDdvb+vQhFepuxz6o9
dlUYb7GzUFlF/G4mx91ovd4WUBOwNJBTVuX9HHDcA8zMbkotExFfNmw/19gU
SU2tCOUMdOtoSQGtwdcziy/JRVU/plSZsThZjsjDLpKPHHXUd0IZ/uVjPHrq
tTCP9WeZ/QQz0nz6zO6b5j5guGWVgRLrqVZ76QYFcFHZM5RKNdO2G7YDdr4S
vyY4ORYScSv/0Hv9g6n5MiUWAg7s0Od8RMQmGeHSbsAMFxTrXPpw+BijCRC0
/Myz2MmKJQj+JLqqh6VEugG+QwmnVzhoufTm9z4ir63chpDZPmXJyb+j1jPE
OGebxsE3jWhHgmWMD4suwJzk0ZbZb+4bW1RcRlWriphy/wAkqZgunWfKKWnz
hRLVfGCQRbw6UWAXu7RmtCw/k9dILy5w6FoUhsKDr0XFEKLJCG3oiOQcqaxB
rqixc6y5s17qaRMeewY940T4G0wW7psA+maBFxRY2lyqhVt7QK+vKpw8LIpN
k/qewkMgobbfmhr/fF/o6w+3ZsBEeXmi3oYimiXQtb79YMIsEsSEBVeo1Ifo
C/KzmdynKn3iWUfz4wV7Zm/2GD4T6s1vHGgv2jEeDEo30kFZW8Of/QJ5BbhL
D2wAY4OfaORb32xsPOJfmiE6CgL8CnR8twbt+8w/zpu9fh4LaiqdzTZeUiJ3
sBea6DOw3qO7hNOoGUjCefeJl0I0Kur2DDvUBRobxvlLxqqBDQKJ3YDZy9Hn
FcTrr3TEroSg7zQwcrDsD38JlfYCqXQHK16RGHKfZZ6xsC4eUAUq6yiw6/Yh
b7JF5Dku7qXMtdnelpuCC10oENurP5iZcpW+5dDj75ny9rqyUiCvO56dvDz8
n2Iep5Myhwlpl58nGoGeoPDamGq/k+LZndOIHF71GyjWXHCfNdBcMSMAbQaC
Tr/RtF6Cf3YGLN9m3WygB/yONBCmXn2fgp+LKANg3IyHn5oPE/qaA7/qMUr9
WrzqDpcKua8HI2rw2EKQ9h81M0SZ1N4JQc7GFJSCH2F4lexW/5mNYETv5v+i
dgx8SMR7JI/FkQC9Y6WA/306avfxkfyz1CViXbPc5WclGzwgle+2vAowpAmK
JQ4LyTYsmcead8DSnGG9mFTHF+nNhSSpci/UWWQ4LDkg05RsfMtPHU8ETFFN
QC/gnFxjfkoqIVMYmj8Drsa+59g/PzODaygjIKH0jgWANuMh1Jcn5FPXxlWr
cNbHXGYr1H40GunSf5H+ioQ7Az8CvmXdz6LcwY6cQhsnM+0kwDH6Xd/rLu1x
MzSve49w+yZikTIXiXPsXbWsKzvrodUDZv3keJ2i5IWTjlAHdt7dg0d7PjU0
m6rkgyLq/6K7SR6lmEmiAn8/5+mmStd5I873kVUixpfrc9QI4LTDarxmRG50
8QXZFCC77/N67RvmPpk2Ob9CY0mhPp2F/pdP+pN3hf2N4z+JmzyB85tPvpaI
kjHYNgXBjA8zCoLDvtBISChIkqCECQAvaP9TNkesywrzgIvOzLB94aWD/kyL
FJNaKsHhmbE9NokU5K/WeVixLQj6Gc+3YUGmyZNkuzDEAT3DLqG+0AKo/xeP
mCo5v8Ys4lq8b0rSnAvPYgJ9GJKUt3yECNRGtaHq1XDbGunuvdeM3IcdH8MW
6L/W73oXMyYkbPBQ3jbLiCojAnAwBiyZ59UrzUVNxcAHIqzNO2G3WErP0kT4
4NR0qciGlPM1jYGoe/WX5vaLmDHvXws4raX5Ovp1Mhm+LHkzhj7bw7boHze8
mN1KIpX0UroXwvfV4UD5Y7vOrKWZJqGLoC5CvbqDVYmSlMo0C66mCjbWSHv7
ogZY7bG5hLyK3f8zWUvNq4RSzrAtUwsjSICzDMyXK3t0vIsDIf+2ZLkwfQqS
V3SzVCzSmm+OBIWG8vT0wEgP34JVG+4jVpPv4ABDwDztcxCdfff+7NDr1WRq
MqR2IFHTD4BFYkoSE2z0+LIIClqZCFCOWqtoJ6hXkM3fy0LmZ0omyF5l95r1
G+Dbs9PcEl72yRrTeAuQaDdylbB7QxOek362r0oKREyT6OVVIh0XOSdEkbVx
27C0RRXOlKl/1M8OfJLR5GTyLu7mjLHXj7Mh5tlnXq01z4bHuklTkrpqUJ4Q
+MIvRg35nNNW+1uKI7hquHdZ6GPszhLPzQ/sVOqt7z9ghJD5seMCFA9BRbnf
YVUQpBVr+LcfQF9iOm7zej6WzgPRqZ6UII8s+ghMeirewF77bNCW2gJit27n
2r86ywj9+y8EQmCHv2i7/jl5lDm8NYdV9a4dSDaEqKsNZObsh0dm4L1Q3rV1
f4XVUuOBTAKwwd4GgnfNzy9oZIz/uCZijA+eOP9PexkYwX2bADS5PLOOTsSX
OZ+6F+65nZAjiQ0mYoQP+ot/jANmfXmUycqkvGMlH6ol92ESsTL9aLz/VwF2
VUBuoowNVyB4NNmuvVdu1bEFoXAgKP6I0MuCvgG9xWkFJXhN4Sa4TuGR52Jf
CDmlt9n9mCxZRyspdDFZJU9SHO6LOOcR+Vqt++Ouft+tM1QvqO2sT4fExsfF
Xhd6mdsjNP7dRBTfn5QTZOzxduMgEVL/UN4msQR9TNx3GtYMG67afeKuCTFR
LqnqkPc2NfkBYh71Udeya0DjybtrlBg7ZZ0aueTjGEmrY/r/mD6z8yQoVg+T
xNXVaZKtFWkZHUwyQ6PfACML6gBGNaQj1DesCK4JJ93dAm5W5cVb5u4RTAqO
YWaNtDWqVOn9+C9lOa6YFLQpsBBsDT0Ac678cz4UZcuve6yBnxwUh7mOPG1k
N+u516gRRzJW+rym5yMq2V3tahiGOlhViomlQIU+dyts5GEqElcTltOlJijL
DK47USWtlQqWfzUiHiNUyT9YUk8CBDTRn0Q5eSeGpJGYLg4CTB2Bfr3krokp
aqjS2757X2h//larXKCv3Uvf9qGm0MYTZeuHVcdmqMxIl2ZSDtcFfwhDbXNA
wpaedKgF6LoaOVwmrn+u67T87h7HrIbFzExvjyT8INE3RPl26aOgwHllrD6a
Fq3heVBIRo3tBZxsifWc6hKKo/LzGTOHTz4Y/dljij5M/1ij1ziYmcGfXR1a
EQ8oDz1HwSMURbcZwg9tmnFw+w/PwJSOcqyfwnDw7zDH6fEjrUUT9TojrQuf
ei1JxDbSObeR0w35Ng89UuGLjrx+HuUFNt5yoN1a0uOWL0tD4Sk9+EgyORGv
sjNXsZHGjaIJKz+T7BCjLF/QKyzZXofUjd8Dr/J+53nvrthj0bGtmUsF4Nom
vdbclmN6Tnhyfwfklj8yADM7hb9PsmEoS81MSni6/pfAlS/ePzipqqbQWPdc
4S8q7LE/na9W9WwQ9ggEot1BF3qN+F41nV4eo5pL+ehOL8f+Mbvp5UqrQGk3
4MEmsXtuRygk5xL8zUMk9GZyLSN9zLwVwnAP5xQ7s6Q2EIDDEsZ7MECQff1P
zQfrLxeylHfwvbZmmzu3UOM4zuV6R29S+4KFyXmGt9QTK8FAMUMgWVWKhsVu
rq/ptlgLcGnPNe5npY7koou71L7BrGThQz6CrcaADu9kA/RV+BRbUGeepoVG
F3BD/cLH4bcQGUvDEDgW7fN+TEx7qNjm7a+ev7xgy/q4uhp5YEOli4hxW1Gj
Xg15cvXYDmxwvCBNcQsXFUjMFYDaorsQMSNEK3DItQ8v8U00MBhjveH3t68V
6CQbcKQAckxrvDSNmkJRVjMocb6NCGaeGkAYjF6kOagybdxD5fqcf6FRiE5o
L6JG5T5DvPiJGMD8BRI1ClskozHj1NBW9DocYSIvUPoC8hsSTJ8e/AsMgOti
M/lllUp5RY6th0sDtRpo7U3gmXKfwIi5cjvlBpC8OI9zxz6xkIpfB9+lfHG8
A7K5agSmOdcnL5Wn6m4kCuPz4nipHNhlUQ749xTFfK1dB34nsb9kwQcwtkgw
L9gX3V/pi/ZPalSBVbt4lH3NG1HDSDM+Vlkr4NUytkdJC2FiUipi4Nfwx6TZ
bUi3VHpXBY0OAyUJYhpug1dViqSu1D7tciy9wXKc6moYlel/afRjuWygp66G
eiDJ+gB96Bq7wRrgHgUkf3DXqYi10r8ccJ+jrPIrZk6Y/oYcjifFiHtSpC86
+udLWOORapNLQehBmEUAHdbRBL8+BM7PeBt1U04CfcsfNnwa3Wkp1Tmag6Tx
a94pCVn/XufpuIsTK0qppkNkqQtzz+Qj5dCV98ilc9YK72gKiXANgST8LGKy
poJKV+3w/4Eh9apEj3LhkW4JXTVcORsGyAiqjVMLMr2DeRhENoa99+uTWEqK
6M46zJg9WUF0LVIm3rBiNXUprcXw0WjbYWz2eGsLJrBp+NuZo9ikOTeNfpgo
lRsvzimhrYT/KCVcC0vqPMxE4sZIE9nVeIEXDNtWvAINPzNODb/6/R+l/I/K
CB0OM5LisP7QW31B9IdOzV7IM3T2oQEGa6iQBHubtAo0jrh6r8+ttTwSjfzb
qT04+tbaiOeD9Mjd14UkiwY+WQ37YiNrNEd7pHqb4L7DVFH0WZhsZwbGpc32
fZY6JW3C1KhaEbloJg23wro/WhO5xzYOB0rvwNjqy7heA4kfzE+AvguxOvCX
lXWT81LiIKnWm5LWyeM8XW6o8IemiAtBx68fdXiQE+ohH2n7gtxlNYcaCLHt
TBHSNqcGVGJl9A99RHQQ5PSyRDt95TgrHxKY7f75SwGAvCICPX6VRXHdgyPl
f83jIp25XXNKtaEDiB1LzqECo/AKsgB63shk/BmgecdDfaVv/WhXsSpnUUZ6
zKKVK/SUsaCHIBTcBw1dhrissXnkgdW8wSvyOf0mGr1CWv5GlAPw1+aPmGIx
WDVisiUGyFEKQEF2tPCkkUb6MRaQjtJxpicrLMUMjk6W4XKAUiQUUFsMP0/1
pzzUYDEu5eWCEfbwOzQGIU3+PF2azlcQehWIVNJk8A7j4nhQ6ohJyID5vwqy
6ryZDAWEPEwur7Oyfkz69VOk5v9kOH9hMrBXQqPnsjWU3ZDZ8/8ZDEUdUr4K
lQ+a+G1qtS7FrxFvBw6+naZC3KD1exZLtK7NzbhrjkqUY8Gkjz/ajSwQ9qwx
5G2qhOCsbrJ/B9fDvlWOUoozX/Kbl0aBq2R1PdvLPu+wIEiue17xv8OAna1a
rY7QmnZYRh0hOmGWAoGDpzS+FDR9gXQms8qIsCP6AmbeI4wq3f56PKJBxlzs
pbCrBUw/ejXABuRNaDGzO552r3W5msiC216N/AbpnTVI1J9YYYB4JsSMeqMZ
OYZGmHJT2gClrj6zBd66lpumHb2t32oGEVWsoORI3tel7XG2fZlw1I+0k7CH
Cf2qnEBjnBSvou5Wzyi8NhPgomNPY2VZGmcpyf7kZHCXDkAqRlFA4cncljPg
yDOUKaRzgOinwdgVZ/gxcIQv20ejODZP9h50tHt5vIgkTl49OIrlZjELCAjx
nMt6sxngeK8TFKLl0MFlype6F2MlldVDGGAdVHypP2QJnpPLvxfiBU+fPt0D
eOWFJ3BAtxMAbi5IU3iqsGVZmvyHrbTsLZq0z+s4TGAg7ISjD8r2/Pg8zAUJ
6aI4vCmM1D34ts44M6sjvURxOyNklBB3Z6GSLq5xeL8+6fHkQcRUBhD0hd9C
Qc/7UYtf9LsB7gVK/yj2qo869W7x8nbIGFu8Dzky011SCLTyyB8nX9n+p7/E
PSDzAssIYIWdae2Igpr/N+oak45riygtdjrOeVRb4lmxcyz3ubggwgkQ3BLb
hx5S1cnX3RHfhKDjz2WpFCKjJUq/nvCVAhmLi6h76pwi53L/Mcjl5D4SxXeh
tk8r6P5wFu2madgTGeyaYjFuRczYi/qFutEUL0jEpx5tW+a50qwtF6gCSBBl
j0hwXvCfz6QeKblx8/8oimxuDOIgVsDIB6DHp1/G/pMAlT+KVw86PxYy2aLT
LU9vhiOyvukKTejULxBipzU1+8qftXsspcg6tbWXewPKzNYoo6hlq51CgbZn
QbTQ8F+W74Mh1NCG0+sAoF7begRLLLD8fahS3JdbhI8qvlMNisg767KulefZ
fivzGjyz2lB9qfoEZfH8vlFRxEcLSwT87zYfAdF6XxA9rAeSG+rvAbVt+XeN
Wgb8oXMbebM2XeOt5gyBNMdSIRx0Oo+5/EtEEFqWpGFZnp3pbnibCSqmau74
XMhT6qHoL6C49wzfi0BRQM1OhPtSPv6TeAVMFXB551e44WS/C/L5md3PhgvG
SYKI10Ffus7dIfreN1NVVEsVxMKDfh12ziJ1JUyRzN4CgPCZ8x4SbQzH8SS9
QFAU9vYBW0jfObbDEJUsU+apRzwkwxn/S+ioq3dR/bnuJ9v3rLQSlRNAFjhz
ZMoQPZGblcjGPuZ223XO9xTVKKhUV6E0L9flXdo4AkppBwWBC7jPiewfi9kV
VVvjlhKBapuGPugrFyPpH+9PBv1jY89ABXqFW6E6hglO4e2tPD+4JpThXcd0
jn+7VFDTRx+GpYqSLz8BKJDr/57unzR4xY+eIT5b96u92FFDyC2rV/1kwG6z
521eDyI9gNKanC1Yqh4VLGj0L5wtAwMk8DnyxiIFe15TxpOy+y8UErLXtpbX
OVsoeLJRheQeudJrwmmvoWFJHlSJgLu6J7x7SHP7EbiazJ5+ZuSYg2eZgFO7
9t1EEaJ+hn63PFcOe1pQa9W+hQzDL/sBwwNY3ktqQ5J5xrwjZUNPyI7QedGP
Oc/S6EVM/fl0hiX2iBQSJ+rk6YiaZSp7lsWQRxPc98O8z4QWkrmhuqPO+IoL
DK9IVipDx+CNH4Ii8jNo6DtGbVJKEsLRTuVvd7/2qROMXJpQuHRuEHU+S1ek
rFpGTe0m3rF4FnQT9Qerip6ieQWxA8nlw82EyYMFKvbHUCOz7beb0bGpy+2N
OEyY+1ofPR6YNth71T7ht8JbmgWd2QD8I/q0itt7aSJstPRqEaN6KrqvsROb
NtO3ZQJxdEfDHTMnrxVcRxKBWGpKjiPpyXjWS75X12iPDMyM96ZRCw4QuIep
rY8qwMHd9WCe3fn+Sz7KBH1AIa2bKxsafo16EJepYYe6ZPZ9D+AU7snIpq8R
UoNGw7OG5MYl2t7nj2XUmCDvpH5RLsCWv0qkSVyht153bzLs0B71KDTkP6+z
iMQjRx5/qyIethTQUXp1RBh8wcLW9Lym9q2mVLW8ib6IEbaRI7olOT+Sx2oz
2dXPJv+4+nCkmdbPtXvbff/8KDT2gwOQpL5CHPNsoirnPTWuh1sNaW7CoFUa
+0VjM4Zg/IizDE5Ee+QbC+x9SPuRKa/qyjAwWs05ZivVyyyawIErFFNWZCp1
zpWCJFfo5MNtTb4Mhhs5SUw1Bxvw4wDuHfmw2pXWliIfyg6UXkmUhlsEfcLt
fPvYRkkDvlU29KjM8XdJFODPcf7YGQ9fDTKHWGtjI9whGV9rKxtJQBMFT1MS
sc7pTiK0v3K1i1BVrN/cCmStxdo34/9z1WlzDImxGxl6QQzwWnbp8ePB+32l
dl7fQIlDaurA7uORJ7PO0cGqLJk0JqEvKH8kOTjjv1B8kpriskwbN+Hizu14
1p0EKecib1wvQK+CYGOyqtbn+8JSfL0yXM25tipOgtad62dQqf2KV6B5ycwB
i6AJPfKPtmsAUrHG9FKkMfcetKL+Num2FppESVppCEyS9Vpq0T1Wh9hD139/
2qsE00OR6xiytLEwnA8u9xi5OXSWBPxrzNao4ydYqyt+VdD5FLxf2o6v8wYt
yp3p0qk0cnbmO0Fgry2QzVCrLGCDDqRPeR9Ky+kNNlvh7gLFuR5folNDED5E
9zjuSt9Is82KFPjzvn3FDTBGXHZF5rS63S3pg2IYF3VcxmDVNvjpYesgzw14
PaEH0yx2LsbvfAfck4tuX0t5tE3Sq+kbCtC2+/EoougpSabFicXHrr/63fwn
EWDgTcp6d/BRK6QTafeCxFrZDJyAYJQd/zwNRvzsZIUsHdp9pu1g5qQ+Y3RN
AU0ok2FnUG92wu6hphz/8bxi424TET2/IceAivbz+9Ynt4soBn3Ky68cr0ir
2TYc8HkRs3/ZYK/f1bcINPEZLY//nDwLIdTbuvhBXV0BrbYoHp4rOjDV0Dw7
FGhK7qz6/8VuPS12swTFo5Dg17ANiqC9ERhsojHyAC3CyIdtuEBiTC9c1LQj
GIlmJUAA/PmdTtEYIlt0L5XmXZxbgQNaAfvAW9nvuLEvOppwsyKUb8khg7hM
zRPg/mtV8cQrfGRst8BkUMplyBRZwYMldKNZErB4iyYaKsgeAOeRVII04ORP
YtqJC3KCR2huCd19+v9ROAFOMmhwgj76kYb/HYdYYQmHMpDoAcVRS6mXMy2u
3hX4tEfSH5NJvMam7QJ7qPm/ziXox9k2tiJVLqoO2WGoorwTelbGYQjbIgxm
IUMJI8MMnjgUDSNEAy5Yl4Pzq5jzobUkPbBxuSVVt4Jd9iehDKFu0EOvnphc
CQU0FqAB50+1wOl6L9vniPFw3CmztsyzY1Ema8narNVYozTTmCNM3DaI92hJ
kkDrlxvMfSrqDKAdc+kkS3jo9epvAHElnjYN9sijaRtkC1xL9kMnswAND2nJ
AiTOzly2Pj8uwV1fYdiHn3vYuO7Uy+NgqLWeLrtVaLRMKZ3Ia0t1x2YqZnWp
z5T9Dfd7xTBLrUterZ81wTNazMLWztIbB1ISZZ1VD3HTySXUJ5FLQsxNRvmZ
WGhGEocY4jM3bqS87KRpKDpZju2Fj7mzlpihcGe2t4tbrSfZE4FZGtac6i6W
l96MycR/KJqtc9p9H3fbywKOy0Yyq83PtACgKUl+NBMNDTtQo2klbcbWVEjv
sMZ8aTj6pyJ9KIlZgHsvLAMdfdueILqTX7ZVr0a/zBcjJxtusaBn4X5jud6D
3hWkYYv2ilLfb4HSaKQfs2WrHiyqz63qKmEcc/vz0swcUgSZkybgjLhmlaqM
Lt/nImnXGUevpXeBmOPr+IuH0CHTIonzns5yH6tB4tgppRcVl/RBRApl4iZx
SaolMiFlizd1cya8Yof8oKHEmngS76MPlPQc2Vie7MB5p76mynKTZatJTpsT
eigZP045a7KTOBIqXvwgr4lKhaM21hiu+3l8L0qoE5n7uHO8AcwsnKYPMIss
6OopDfGkJpDuAcMoN2FCb1u7/UcJYUd9FJtyARxU91wD51A02aKVfOgj7zD1
4Xf3hVXCGR3q6wgfsK7/ik83xwHiJ76rWU+O6MyG8+OzSWCtJpprP2IpmJpa
N+oYhyzUURN7WJfrM0vd/u4iMQ1JiLUUUzjS08UpK3okABXZFP1LvPlaSMGF
wtyl+5eVIgDUd2X+oZvAo25zKePOBYX1ua6Zm58ezflF5yJGqRxYXii+ImMd
xtM49ahIKhx/pF9MNNz9padiNzhvdKMp9JsvXN9jbJmhUpOErOcCYIW2iBY1
za9MdGOxnQorZeA20XzctOiOcB3tYH8RP4+bAlc/Ky75HUHySEgqonu2jVHu
StAWR10rk5M/5rRDwkzQif69qZc1nJl7akfAtqlxq0ZMedpZfRz7diu2/8se
K/d6ICgQkdUK2qsOit2o1wqaGJhjsBpjup9gW/Q3C9m9DpONPNlUzWSfhh9P
svEYQCh2jVXissbA1ZDG1/leJiM8akfWirA6iSQ5xXd3gJrxVv85KF0UnYqL
ul0cpoa8nufmeiE9+/MS3SE1tlULyWvjxfhVL84bIlBjyyWde4np+OeQIFuc
UkqGSzRhqIbczfgt9x/Nwt/zZB8m7KUNgCSrZR69H42XBw8Kgmgc/Ydb3H/o
xYeXHVwUz2BdRjjLaepslGvFvcDXKbkfUMbffm4RhTOQnHkNWNF9tiCuSy96
LEVdBFbmhGMJlW81EAOAp7pBcZLq4FGdsaS9mYPRMMJN9hLAuI3Zuihs5UEU
8x+uaJ/mfnZopsc9qtx+Og6pCs/bcWCpjlbTtTya9aq6iJCr3IbkwxtMWHou
TOFyH7qNFHTc+eItlz60p3PEDKvwOB/qR1AkUA3RGzvZCwLxFcQiV2cW/FyL
U/ZQHHM/Jo7n3komnwG3ZVIS79wvOB8rzFBMeUBlEVJiCkQ75XFftA8ws/jC
gCt6lcU5g90/jBdBI4QeTOpF7JR16+THr8JgeukRwEOFwiyIoI1NxhDoZn3k
ssDGpyOByzSftatnsAATYrI6LeX5DULJF0zwEEvJc25QSxPfpI2GRjz5y60G
o2NXjs/B2z/XcW+DqreyyG6xHxt31Cm7V7/qs/bNnyErqNC0U2fI1w/nIeLp
tzpbg3v3JrQWShUDNgPczx1tZbpL9UGFwPossJjvqc+kUDxOf6GeWPuw9hps
3jkm9Sep9ATHV5kICnzken23OLqI4zTJCzp1UJ4aHsp8qijUN62IcypOQljn
ykYN5zsKpY2lTA7EhuYtMRgwIItE8ZPtxS/rrfv++nZXN87hLYd6x7VORGru
MlJJ2WHhOrdXa10ulx2C+iXqmIp50OrW9AaoQIfCOhmryfKKhHFjdegU7v53
nsUES+UoMUhTTMhOvuo19Clg6ffDpb+QgY0oO+Od9kFdfGfw4t6fcxWZN6cP
z09XXOE0X3i6DSL18aGUx+VS0VgY0ryQ98J1Ymx4CAigskhQFxOjVMPF40uy
MroD4V1LDuXwMWnhmI/nrfy68ZCMXBsVDLbhrUibmx1FOcFiTqiNCkRKMu5i
Ps4kJohqM2YKuxrEv78KBReYf+LXpZla0c2uOHjJ39jgiIAz9HcIAUtTMGlo
3H4PDmBybPj/QFfo9P+TIO4s1QOhxwIRkHUYB5fK21O8mWDuOhhhXUIQdIIT
Kcx9ZXLF4zM7vht0Sw36duApR9oY+MbxJk1fzT1QdwTdb3h7ZZwfQ0bTtlF0
luFDC91CZd9S9Byz/V1NpcgKYT2p/kOmYMCFDgOc1aQ9KULJxzocDNcZvIAz
c8EhWuSP6Hy3Bgg317Db6Y2m6JefLIAQVgXcmRHZOCZnjhBa5Mst1vCvEQp9
+vsJ8oNx7klBuxdhD0DafLd8vgC9EZGP6mXuMmKGisj8QNKmGmLE0+8VZnrM
paWXMdvI9IqvtLgpt5kj/rEz/fV/ztllEXtUIMc7RX0U310JACm++v6QO8T0
fpn0Vq04jhGhg+pn9OHVU3xUd2IOhpvI+anFWmNJ5JiBxB70seATuLef6xYg
LtMkdrJ/4XQsd5tllQ29BjvQsIi6RHOYL6fMCnnZdUGhnjlkKwVGhyismhtV
OGJt02jBPaS7EQ1SzVEVWQ9QlMLixnVU4gnzoKTLWGDeYJ2lgqbCrFbT1mHM
fXAjySywL8eNko2THXnbGQHPDUHBHQblYGT1tFdK9gRxdAdHF+1JH8vLPQGJ
MHQN9ei3RdE9riGJXtNZUqjoqMK7D2EZPEQQSH6LWjHUhqeTjZKlHA6SZW6o
G0w1JdQO1/hQi3Mk/GkwzqVe2H2qgwuzuBZrrI1ol5UpxQ32ysgYQvxHDrfx
+Wrwxsr1jm9/trIL9Zjr8CqTucQvFUV/OyVhSq987nTyAmRmDri8qgcO5w6+
uAVPKYWDTpjtzFgojNAAAODWexc5S3XF/w/0WWx9e/2q3/fO2sMoCx7IdKPm
+nJJoJGth6Slf9vOIFsG05UKVjiXZJ/2oRIEhM3zuyaYkHhkf3yUgYHX1l1T
gyOv0BM2wycmNGS5JvfYd6CgH9BiqlDVKY01K0RRhM0lUb+4mbcqA0pJm5bP
r6nz+J0qp0EIGfwwgIMxFLKszxSxqYclqDkLsfkkIcxT4vCf/6auAdw+pgZM
ES3ZHk0FycUiKTJKkN2wJtjUZ1lwSjfKQXzv4BNUiAzNoxrwXWUyRTVSIMS6
2zsFW12Xq0eM1F+ZvD9PfX8jqTdwUx8VSqJ0D34r1Db9zSOJYO49GRv/EJhv
AbK1mTWS+K29Dm6X5O9H12aOTiuT3xVrJoz35qLmrSFtnlaIo+em3HNA3OZI
4gGMQ6ZEERS9D2ICqckvJY96qk5m/Tgg5P2FvBZqxsGPQWDnRAqdW8A1HVoQ
SfP5L46Eosowovgg+EoXmI6cYEfTYPSB2ZCCf1ggl59cdizXGy/5OcnGpbuH
3aG4fCPhlZ4DU3D8jV7W9OPfcIzzIP8ggDwCICM62qWCfO7lXW13+3aINKmY
PAcN29FlxiVsQP3iWF65v7XWNMJCEw8+hRaCT4rWUAnuxyRs2DL4xs3Gbew+
9f2IcUv7FMTUSO3w9USieDMLWiwP9kpgy+p5JfnCJz0jXy6SrYaQp6LyXcyr
biZsfTWD+E/YZf0ii9S9Ckyj5JIfrxeWkPW+rhXyAdlw5aP/ul8Yr7Adj225
a2OD2YVhvsIws6A2ZHh7rVuuL87kTh+ySfTNz0B+Km47SWzNu81lSikdq6dd
gYmnNgiTmsgJ6y4+wNCr9yWfSXEi963tNfadjpQNYJL0qquvAF2gpbkTApI0
mU7Nk7/dQ0qfLrrfSzLhI34dC3VrzSm9PQPmUZAJn/SvvPHDYuNmGRsYdA8X
uoIAHFM/HcJMc3LTVVToUgBK/6fOjc/dIYoifXUaj/2sNv7Drpi9GYNVHu+L
2kElfT4HeJ1Gc0+jHk3T930mk8AGlNfXj1QSLhgIcjw8tIBT8LQuPLeMXWz8
xYRtN58AHpHmTIN6qSZwWUutww1gb6RH6RmqOAbc464khrfNZno5VzeOfdwm
zzmkelEAFMX6rlwRtf5OehCbxOsn8oUhb9UGull7UMjKP+jmJ/d1L6lxg2Lw
FKWmSEAdnYpw7oytt+zb+CK8BFtkq6aMFZpbkfcDwcroabO067SiUe8McdYx
SkkKmCpMk3boam+isDKzygLTURxtK0gUjvM+aEAGYVnupnypX1fWhkzjUjNj
yQp8/5ZhmEJ+dXXeIHZhvO6YBTXWLpV0ukcGKDpMYV1J7T8hWkzu3vZY79az
TQ8aT1p3eibiule8LnPOq7s60aNp+e1cFH7V1JqKUlukrrOeJ7JqRrc0vmlX
Yx68PpPYd8F2ZKOPDnPeKiYIZTJ23GMLJ1dC0i/31JfdWA4SS0WpUuaHikoB
gq28LAQzqW5rOAuPw2DoFe+N3mwq7dnB3Cp9e8QLUBS8cBvjbKr1Et1cRCjm
gAFxN4u7dm8NHCwU3SVgZ4nA2n4OoLU2SPx6RzrGNpwgyCRZrxk1njlH5CDT
7BIUZbzcZxVPSBfHLiU5jAKozO0WTvKwYoybnl0wTOmLY4nSwjTdOBN9GH8b
HUsotBWE1H8aDKenrdte930/rNRFCLL8F8tDk4TQe3/EaNaHdYguYA55BnN5
COMEVrM2mDxPki2EauAqImLZ2RGjctStLiQyw/8sqtngJojUuUpHiIDT6TVq
o+RTWhdBbi2mafTcLZ9YB0Ov0/LLbRJp8t6V8uQ23YdhAgCQJ68k0RGhBlSS
UEsbAMdzsvdz4Q2cDADR2soHDZcY98haNvDAFARsztjmk/ZV2UQAw5OTQhSW
zkmhEQTE3PKhAUbtGITGXqEoL5EzuWBMJENYBXVxe+XEzoSLvsgHkH7vJU5f
IlbbQJe/GundZ2jp9+2uP1csIWCuF/DBrhRcAw3vFPzytWTJ5ZSSmKWn00hs
0nFfBsb3Gaoe31YpQ6rFXGotG7dMbxbheiNc80hpDdjCSgUftP7aSaQ0LEmb
sZ0tSkaiGcOIUMPlAYk2VY0kCQ8YvTdntMqO5QCnhRY5mFrKmfRkEX7Y5cI6
qrhBYIISVp6n1iekAbWDYMQ72gmBro20zQw4hz2PeEHUjhGYiHcC3e8LNGtS
ZLZ0Q38OMme/uucISWbYPGbUbCzyYOaVgYfWXZEOjyn+f94WQbmfI0S/3Dzb
Fyi7lL08dE24HnRuFUr1HKslf3J988uirSYbgwlZmSAt+w93hcYubbtt5tHN
Hn0cz+WQybfFexnx70LNrxkAS5KknEOwojy1IUtO4qwFM4WRQvMf03bK8uij
Gv/GVYbpGX3SnlJLPmwEChEzaKdxRsnrKncGGQJWGM6GKCxh3s8bBK33fF5T
M9zrnUilzvAXnX0cJ6huQ0RWMOEJU/7G07eu1jn5p82bNbrAk3lmyp3ou12x
TYpjz7Qu2n/pD36gyw1G2qJE5sWiWRLK9l3kEm7MaPlnMj9vKytEVkkaWval
YKR/4gIAerRE/ZhhN+6/qzfNUhvjgsxARIoCaR5xGzOpu3K+6s11b+iPa+gn
nDyWFUgAhJ1QQtyFrUi+8lylcgCoEDcrSgtOyARfZPD6xjNzN/xaV/okagSx
6fH/uVIX9HTt1owOJOT7Gg+GAaRv7gV3OeGop6WnvksnD0TCnu3gAy9VJQsX
h3mtP4Ud5jB/j+nrloM45UtnX9jJn8v5vDfYo92FROkcsIrHJ9aw8hyARPcT
cBZMTwtb/3vWy6YxdfG29bL5bYbk2LNL+XHWqCawxfTjoetA6ksXrt4TxPWZ
11PHh0Kgmc8BlvufE48Z5BRQA+d7QFDGu4aSHhT4223AI7EUnc87OF6mNLol
pXxzsiOCir/VZJCidRNwyYDM7+W9oS/TLh4dI8oggRV5LgLs1cO5WD2p0tPX
rJLwFI4Dso3BkKcTQNzQq8giqzZEj+5x4ypqALMLgxttctHzytJuWoIENiqf
FsNhBv0/+qZ87i163ocdBoNDlV45Pz5mmD2Wds3sylNb8C/Z7TF6YIVjp42P
9zpo7ygwAxbWFSOhn5CrXlje+Sgnp/l/T34wdMCtvX9HvTPPgu9UV/MIlcri
7xFkFh3wr6ArUfIB8MOd8vzhsnAknMlUKnq56X+3xQIBQYXqAZEhmDy1/f8P
Fcqn0gXLdHmPbbdrj6QMGU76GRFVIRjvEkz/CXdFtDHmzN2VgOVdfg2uYCdD
zQRXLRkMwvaTAXzHwftGTXMPhxFNSp8VV6xRHyNBFl4r/Wxv3mmOmB8EbcJe
2s5xDzeN84l4+3QmN2vJ63H0vn5vpISTFLEFe0loeEa6dPRx467+9f1U+mIS
QUNX3bJDC1j15pBavcCpETDb4Ku2yiY1vb7gxdwqmLJ2UkhdMslLQKhtTPLF
BhZVhAOV0k8ZsesJqzZkN8+AM1o5W0YTC8kc6tB1tMuWbQP63nYEea/jQG8z
uAd+wDTo34sZV9qmocX+StZKDsV+wwky/1af8awLlICp+Qs4QtMCSgBwU3YH
UMdl7IQjyTe70eliBG+KUne0W00jRg4cRvlyyGujG5+lmzuWoAhErlRAZx0o
cnnsYJAPoU/0tc2ZIV4habE9E7GhHpcyOSdHPltGQuKrN5uqZ51fX/CYC6Nx
pxqf6bGT1XCzCcXzWViEFielLCK7XbchIkxPzBD68zqWi5TQhGyP2Ec/qoJ8
VTYXAwY4eDGsEvGGOyH57dHgF/eJkXD4e5CNohpIK+GtJAhbj40jeK1Q4KLY
UCbZ/bKvfIJ0FmmOcBAeX1UGa0g+rckooN6o0tOsGUm2kw8pzvA531GxquYi
kBPIfzZVtKYchlKwW6pVStPdQNG8HvZzVCkc9C2PQkpJ7eX0FJljGw3jeMly
7cv7rHfFl+Jj5ZIboWt27J2ioLmb/gZD9AXROg1tKjgIDZFGW7hRTfzKnEah
cqiHo0nSUjTCNMDVGZDQNekwyM6hNxRJeEDjSaW28ntRtdO+g4Ebg6G2hvUp
1UxsiX/uCnvSJpxl5oEtqh0EapOP+vaF42rmS6XDrLR6cPordOz8HNfYZkoI
PCFXpBt/1NFve+XnPb6r+dr23BgC4S9bAkjP/4OT+fF0rBaOzxZOKS+B8s04
nVJfuAIbvTFN7RyNNJ+6ZHyk65kqu7BsIDTnfTpiXxhlJsy5+d8T+z0tXYc5
r3u2M2l6ZPhGKd7AK9SkyrEN/LHbfYQCTw4NgPzcUlgSIcZybFQo9Ve/Pm3Y
brLrjTFS33LrRZ5ghID4J6LpYzRsRWBCX7g2lt2S0hwNAjBLw/K8M1t1sKG1
ATUfECy/bOTT05A60KH8YHfBzE4FKExVVERPhddtrobVmrnU2SK68POZFJmQ
KmTS+GTnvc76ExE3Y9IgkoohQGsztGdUhmScChAVSLs2QEiP/bZz/m50PBBo
nt28BrauEJtg1FzaQLfiiPh7lY4UZRBs8zHjdTDG1BnsAPCo6odCjPqaXyfP
znmlArKxa2eMlTgnTnNHxh3fp/MyHcOUWNImAfVHhdBoohua7Nku9/JvIP2j
cVaxj7gfvA3AxL5PPxSnQVeBeZcmxw6mIuKRQ7MJWaYVoFwuU2GOcGJCGcVw
cji+RQrEsFLCjbEADZa8xb4Bb4q/9dXVIj+W0r/aGWhU+aZKS5e8dAXj/3iF
aHLzLyMFhjoyvHSiL9s21LEr/rCqNsYiUYWloUPjSBi+tBqgnOOHyp8rCLjl
NZ+kYf1GvLMU3I+S0Z8h6Goz23o6uP1GafW/D7xviEEM7nCRPNWdNz1DPDah
gznmWZRr/L7rD0wl+F1Fq71ZaDC49c45BGigAaW6aBvOe3fCeamfj46sGxrd
iFIguBpXttqB0DZmY14/ZxYor3J08O9SWT4ffiP84iQoTW2zVlu/yLRhmxHA
UfzLeCVqR28ZErAAiQmLQYtSlPGHG3XxZiGF2jZNxDIy/Ejj1hw052hBLror
xzalr+ukqsJgIk9m3LQWJtCt9NqrhBWIm65YCdM/4hcfmjLENHJQDmDVdMoa
dLGD+iL28T3Z02LIE0Hl3w+IUDfkHNVXdcrbDQFQVF3OvuIPYCNacolRYNaj
XeT7qJzVgCKuL43+RdBsUxZRRNLVLfMttvLN4vlGuwhEBSW3SkiBuomlx6iJ
alzDF8n/q2Q38tlW/rwfPs1hVfusR8O1Yay1BU6vNOLA3sTgoqDFj5+T+Hgo
J7GIZUP39uBfjJ1GZid6OLnfKSbhqgxJ4GlK3apqmlotw9tptIUOvs57vsXw
BJF+I+4U/Vu3GaKyj0OTyC4GoOCiTlCNbmNTnvCYWKyqya+NXrPxcqQ1Dfcj
8MAUx7yhCj6pJfsICDpB90dsh4QhGMqi/+Bm9NmSGkmhfVRtchVYPk6XweSI
h9PWz5sm74ksUjGmqX3OaZfKVQGXaSMqdxqopKIsDKGJkqGBclO5RIj2l34a
hizZwsWnHM1wWKzfO9BSq67gfkgu5/dOpZP22xQ6BIYS0Fp+MaDfbwDlrJur
Kv8r8QXL07jREX/n3Y6ZCdIw9gli4qxSnOmxc/zPSlLjPy9utFCS55iDE47/
f6wjzl8Vh7j1KzRsjJMZk2qtxnUMTXtG70dwk6/d9sHpzvog0lun9+43lyD0
NhKyOmzJocpuPaLiPqSO0aLSSWSM8lQvmtZOJ5mrnE7bh8+5pwqKtfzEUMSU
9QgYXCvI6X+U8LKmzUycV/jWWhLAIWIrU4GTyXxlmAR0YDXEP0p8DDcHEfm1
bVGaQlMeZetTABVtsnODW9nB7KG9blvMMR29WvJsfBzLkQnOYzYIi4KpXwFM
sxDujWRG31k92PNWmV7CnGwbn5dHAXD6fa4RNwp1rrRJH8vsN6W/+pH663kT
MDdH2rXkVQqRB2l3b8Gj73FK5APUDpz6TU1AlPEpLvSAGF4SAY0H96Q76a6u
uMWygCjvict3IwdGdZ7G7iIICsyKVLApCXfGyozYhnydjYOTAVuoVqMx51LX
WHE1ooR1LqJEGzu6fkOxGqS5SftKIy5y5quIeEowH/N6JHxh6q5UZqpBnLgR
QHQVKa/+taSwJFR4HEzGILRHbWJsP4Q2XYC3RqyM35BWBAJIG1dSI0o+ZvMN
FuCpG6rdvNdMMxjRDyAIhj0VIHMSU6bb35wrkVXMXfpgJHY6DXvUozsGaHL9
8vGuF4NVDUuxRekH7ChkYjKPU7rpywb+m/KzlE9GnajwhSXBQIFjZ+lodcxp
12n+858LrXDBmVxBXU//4V8ryM+AXOVaqEbV/Zr2mt1VTvgCf47yLaq7GlVs
8jxNb+a0dgZrRe3NZ4Ck6XKsW67HB52DZs42OsvEJnjfJ3rKPVZesRu1ZcX+
QMMxadhfFbE7NSzfx5mcEFla0AwEzdDHoIrHj4KMD6bEDwJspwNSlaWMs++E
k3UpWRtJkcX2wWm8V6dtCWbjExNtNw2sYYjo7klg4czdiHnYH16cFdZcSqpX
9s08O6vQeys6TiHqD8yZH/9cK02LOx+a6xNsVyTnSjaDM2+cXXLbrb/aCq5M
UuN3M6ZckyDNkHJ25Gu1AfluRikmNP2HSuFmrZGguctdXqVX+WACzmvMXSYE
y50QcyzkCaUzq4apTvHWYDhfGseEXdfSCcL6WQQR13Nphhk8qunYNzMqPMmU
U0YY2tyvRa+SLsrp38JGhaWVTTlCIYjf0r6mtpeHJ7gVIaE5OFxxSmfgohys
XEDhh5BsFhUigMU7RcTgNUEMRvkjwDYJyYtbm60xtA1vCFIlsAVO2l904S0i
NFBO7comnQnTsML0lj10tGlxVr2XYM1E2NzxA1S9wcn7aBFztT8GZRebNK3t
p1G1ukUYidO2mF3okeTYVdUbDLZrwkeKfBCU8u1vskoTvqDOzvTg6b3tTKhV
0QHDwcJHGBbO0T7z3jnCqt8lk0MpinNUxG7oCXo+/52qyocQnNbotFo5ph7g
WMtLfDVEix2KwGPkq7CQcKRbNDELiC27DRh3ZISPwcsLxMnC0oW0hFrQciTQ
4EjJvqo5RECC3IN3YclgDCbs+iKKvJ6xMGMR1MmkxwODhQ9+9iK5CdR9wUPb
AhABZRl6sMoTA8Qv2d2B1BFiD3XUiZMN/JD31B/1Yv5iyrMcpcCD9fczrZ9Q
1UM0ioHgUjrClPoe3cLH5HhsG9SCIacDscEKdSKjhZYtl4YDTH6cQEQfcCtw
MNM+bBre/zCC7rH1f4tgpKYya3P+Ytt6X+tjWFaM3oWx3cGIIArrztPLKtFf
3uVbJI60g7z7edHXuw/5J3cwjeZtf2H+CdtUHe+D/Q1sGE7j91vaCtaB1MsT
VLOf+ab2Lw9Nw/wspUnrPQ7Q6VY4fJSNzEAUU0nEZVxBPHzZ3Kj5jPgd7qPa
zZW9tPYox+emnAQxZsL+Kx+8zr2VUdgpkxnMFzS1EYg6Y7Bkw2Xok2Syu6Px
FRdSufhKAMTjfiKcKaoz7IZPFivgXOJpjpUseQQW3Ji6dH0qZAurrk8OZkHB
kJCGU0vL93VrC2ZdvYH9n8lT+fZ6DaHGTTb8N8JoADSFZ/wnvRVBq7H7/XDG
wkUkJpjbFm9hb8wZfkBdtfVmy4zwfNy9BDAU2mSPnwIIcd/mZ/Lh4itNIm/P
hdEvfrC2MXnOu9j5m0/BBQoitXHehoHvs3N3HfL7ERNq0CG4oDDnd/KzNSh2
tazXUVzyTr8cLtauu0OOoYknmGW/XdTQJ1zNev9TziQVXdCfoP+F+PCsZRb5
EAGRYUtNpt4TfXjs2oXMS2Dh4Ei9WMeILYeqFimWxW8SH10umRxVQNfU2fTj
Yk/KoOXLXu57GezL2MiilC6eDWjLkDaEQhw6n+J0CFI5BxwvvtvHL4KEH/v3
s543/iBFofSvfqDQUeBp6An7CmV1xY17DRn6aP+IbmvcOwV6WJT/cNtzv4L7
yDpoZy0ZMU7AurHy/TVtVhuUFBc6kFvMEsVcPrpEqzkj+xpEjAHpUWiOFx0p
whVQQoZH6/rxW/q2TNXmY5Gnf5EcHg6k3Qu90lCvmUSNrzCZAfhhhWo7cLu4
LvtX/hE5gcCJekMG3BlSRlpYD7QUYc8pgLByRldCfLEuDDlhvVFd4PCf9ol2
VX1cqlbLaSGoST50G6fG0hLigl7wceE0UO7dKcfDXDVvdx8Nw+wWNTrk7zYh
un/wVjowFe7KjeRdZliOMwxQYgNhI/g17AtJH9XDpSEh9Fb4NLZvbiiEuwXX
XYeavOWN/bH47AiqSjNXjTPwTGBFsLM0mHJdpMX9u1HLS35rlU/QHxp/1QWr
yW2bDXpl5dAFhhPKtc229sZaci7oM5SVeppqBKlO8zWFgv92GK6eDBpMxpwO
f5xNDa8GeDL/k6dzZalGSajyAuQ5ShQjqaDI5NyeAFy9JQwemV8iLnoV8sXb
7FLDfAdRYVOfAGLQ9c2zyit6hJg8b+x2n6w8jPi2qD0bJObuOw0F/wzBuovM
vFkBCe881XJrDQHvOhsq08RXu+iXvHW5ABYyRM3omJjsMJ8nmGlYGBHEe82n
9DPWFyJibhWDCI7ZEeIcpiHlr+dJICi6HZzOXMknHRWxOCY5xVIYCb4OUDIV
1t9hxNFBOa5X7ZIGxYeOyosStkOl4FwhPNlD/IWNCodghH5uL41JEs/w06jl
qMdqtTzaIdcYvUMVpXCN7whZK9wiJd90C3qqrFgaRP9/7rvFNY6xwaMV6613
zlzrfuy7kzWYvEKtMSorW1qzdda11rfx3Q80sBdtlYMBo4cgOPXqlji81fsA
mBBLihrYWW0LWjoWW9by0sf/qZmm5dBGAZXojh3RB3XNr26mwFyRNKmwwqYt
hWzAZknJc8/4HoSeGriszQB6y3JJV5leVRJYo6oU3eOcjwHnwztiwXpilM0h
htPAmnKxvDYTbCD4WDgp0eAnbXi2d/6gMtAb6H2jSHN6KRaHCyBmtElJswWj
1Juvwf/F++IRUcWb6fbTNRmz2jYn7qwQbkrC4VzEqmlgAiCwErcBSOALctZC
l5Oqr4IDLCLN4s/9A0Fq/wJPZrcd+4RiZXGa/cMkcm9Hge02ob5HnUF6bhbW
O3Md4Umb+ZRDdfeSjg/lnKSGJLlB9/EtNLEOTNhUsYQfriWuOGHickJmj2j5
476q6H6nIKnNAHIYlU2QVxjrLNXNla9LRTsax+Qi3czKj2f2XKm8XvvxfQHw
HbzFeoI5cRgdQIVOypsifnrDYGs7sY1x9sJmTlvMZ3VKzOlUbdjlg/sRNJ2M
XDHEPAT+PT8ExKCmHqu/inGPSIR0g0YJynhB2531f9n6K1oq2YaCsx7LrH6Y
BITKd9xmBrQZrjz/9e1F4agB+J9X/IcAZKL8Qc1EwYF5A5gI+80+JbgJN+mu
KNpZzway8IxQ6U1vHLFSrZNotbb6cQuJKk4KAIG66OeTIfNoTQV9c1VYjHvS
F+Cf3Glrfrqm3Q0xVYK5gjdrMvLnUGbtB4aSgFjB0eU6NLzAZdzSXw0u+bY+
dKNDSALaeOdbgeWJ/+aMV+Gh2GcKHn2BM78VNR2x3ED/5mpYUpevRkeM/YH3
B9tggRIXHRiDwrVoQgHbqELLXC1ttpOwDjnz/7zIbSUHLxsWQ66qFeFVZXU+
pOV5TdNugmKxua0RiQ4OEmCT/FeQoVjWLTSO0W1zCe3NOPynyqMZn0Gr3rZi
drEfBPvKMLET1TtRDVR6gErONDMRQQzJeQEIZQQ6+YGNqvRObhYMupOucWoi
xjq3Ag5aE6knRe4PSTPXtmjr1hgjnCNx6i3OAfp7GHh7zo4fQTjOTaeknxNM
m07+LbRPTO7LFTxI/VHaxWpgFUsHufZi//xHcqEaTSOcOCbJ8otvmQk8gJcY
3irhXfZP2E1FqRHOcFdpZ2iZs6TdWZZkjH6vs9lXEo117ojUybQz9EQM6UYJ
FXnTK1sceAj6WyaOudJ47QqT7G7JULqsk/31LTFvGJjGE/6LvNraZs8SEBRu
kX9UCB3wCfulMzQDvQcy6VN6pYuFjalb5TQX4o1UWfMy2IEuJl6opm8W8rfD
UX7sBq346NAzx0kbtUbvPIoMCjSiPAkLJ2uQqGRU1MwUN2S4WJ1LXFW0P6Lp
RjXhPnIHQ4//2FtozlWqFXuiGd63zrYftEku8Yjo9pzvl1Y9ZKP+mfaOMJnB
QCBnXRFomx1orSbImfLGOEpK5g68lApb5euRXpIQBilMh7y+rk/bpFXrRYiG
9H0x1KATuHgROBOW3LPOleyFykjlo4LSHCLhhz9FR2BBC2+LH8GhY/H2ov4T
I+VxdT6Rd7dzmn/oeSpmlsTYcEXCYgAD8J26LgCPi8Yn0S3tO3wNHqmkiUXp
P2AufTAbhhDwVejfEecU4kZeFpLaz4pjFuc6dTu72wIJ9G+qn7nnkYLAGitk
JeFwyZwmzTWpWTmi5rXk/R0SnuQNYmd1Irqka8HHYigobMMrKTwarDvknnJ7
r2gtXIzFoZd21xU1Z9dpieUFHzcHmaMT8DEQKS+LUgWQFzS4Y6jTG6PZVvQp
bsuMQYDHkTy2J4Nh8pWV6ttbm/5Q/luR8PMKn5ratQoACUiFyWcVYsgrQlhc
Yx4795UWTKpTOjJZRwyoEgLm/vXe3tP4awLRV0zaG8SpG67uRH3Zlzk2v/Sv
/JhQviCbqIE6DmmAE9ei/oMVP5BORtXjqenIB+QoIz8ug24eMIdqUYCK7hfU
ZycZTeoDG1RKd7hMOiOtOJL0bLttNPVJBrFDtxoHhOi9IIrwXdSp+afhFDo5
y234KJCEZxxnzUNgoeIoPTKrO1aHM1zc4+i/agiXbkGk13nWesnH3CoyfLdG
wAur8KdVrmQWwV4Xyd33mxzvVAQvxtuAfl+hGX3JPkzebQ8HlzHeYfEqFHx/
fQOQAImwpEmJ6aoJezcHGnBsEHY63k37h72BuWiiijlDdeihAJA1nM4Myzqc
9nuVjNOeq41eqoRwlqfa4yox+g1JBKbdHqSRTqBJU210hT4+jpQV1LmvWXUV
Xy1t6g0+WBl1L07aBheHZ9FGntz7ndp9eT2xXUiID/kKa9p5I1bgRmYtcpJN
el83pRGzVwZ932lK3s0quaagVLfKvUngmgtOuej4NpujdlmOCsaAKncdoiVp
1dbO+k9XiXpMGrO/lCqnImimJAuPyGxMc9rKJTBkNcC5bc3eIWOJzHWT/Ndh
SMPH+/fmJeiXXzEqNEaKGsBZuVzA98E5Pdc8/MtPiTRRzqE1sYnr8ApoehE+
B0RnQ0u/hbxpeWKSp9Br5KJvz4oxU4JqZ9UHrKu+2ItVOKUqYmsHZGXDDQnQ
/kAb5cDDGawaPs2iBJPr4d+Y14DFWAK/hKkts+AggrEp0lzG2sCQVwLZ5XmB
6WDU6HMLUX21qq/HanEcEvmwIOq00mKzkT8Jd2f52fTrEnzRFf+mWAfs0Dsk
lzs4TzfMjAmUhGlxI9tSZ+SPcybFtEjtKEVUcb62Qp+z8L2qjw0ZbRRWGJFy
tmqhMxvLiLU9z1rNh0VpT9CHAh8j741S9VZ5prjVA4WQ/DXU1oTTkvjwjG16
JHqwPLOk3ev0HBIrgEtDC1XcQ6V0YFkXHOL9GUJUVmDstLs7cDwu4uUC1Ssx
eT0SJwmy9r69/11q9JwafOYY1OapaLSLbSQi4moDRt4QLSNUph4dhJB0+jJk
h8e//hGNl3EhLqvn+2DWttBtU3bJ5CxPh2V3xkY1zdIvNk4xSE78r23zDn/f
bU982hhD/xpl38QPfhUuqOHTLAb80bEGnVcKnwgu9EPX/TiMjR8xd6GWHWN3
x5SovXTBrr4Pb3/artqb3yUJT+drkYWIpa8T7CSOWiTX/AbiKtJdiOgEuC2M
zEh1A/duDuwiDRtPAMMHRVdnMt9K82lXUROSyvlNzTYn7o8piLEb0IQKUGRp
od7hcwDLvDox9gj1OZCxWsLN+IoPQ5lmi72N4nM8j44rcU0WsKGNegjtVsl9
u5nQ9Kv9vIna5vgyg9gx5udKDbsHPfVYBVePS1ddjnmg0BrBFetu5F6V431U
B7dG1GcGrFBfmmo1fwc7LBpkhEuGDvJxJiUDE/OUVJ3bDZuWXcX5xz+MD7Z5
LZcCzcnnMqX26khxRd6zXEKpWHWsUj1hN4t/I9m1y0SJvULbguheyl7iSHa1
Gpw0gg2AJQa9msU21d2ItXZgx+MTvNOLvwnalZ2laKLoPLDeRbRQmDKKvxWf
DQ035lhJRd0WJklz6sF5fMqRSoShn3ZCBeSmEsBoCBjXCcPX12N1ZbfOq6Ex
3auAwuD1sBnq2+NxRaO7vYCWExwW2/hmEzDzLbpPvPF4uwctl/6fgQNmRHyU
Gg6GknzosP4BA6S8cb1s7ZY2xe4ww0Q41GRqiULXy+rqAfoXsisuVUkkUef0
Dz93cuqdb+T1aLFxPnBd2KcJI7Z3kYjvNmcpakYJsiTTaUZJstqC6IooApVb
KvoSuO5QDUtQQxG2NxI23j3izWLVxfqvdbWUfSt0jllpH2ffxHS45to0kupG
yhHAznbnlIWinzevXzp+0ztNFyovzfYF0L7jETWaBGvhLbQxDAsX0IkZ7hsg
+9QVlp340sd1kJB4Ka3ofi6A8jFZoZpNCyGpDzOD5j6nMLWR+eEkXoYfJHhY
KsPI8aTh5VELtOQCiFTFtJIA5rs2VbmHDqFQOrjgfIifcMNMS/gluMW/TMdW
+olruBzl09AegbGaDbrWu3td1JyPxM7vlfLWspvD/mRN1THkOu9xwHyyU7de
o7LrzqnyWat2/Iu0fwMb58O23fL81dzSMqsivMExcr6TkUtejGQhFUtrTyM1
oZNrsjJm1VqENsdNZDTO1im7aqnzed9gW5ZQ+6SNokrI16BuzLyH040TPAxb
TRTBzZcTYF4tAA/cZJT2Q6OPa0xCubWevobt3Mfy5biWcGQvPKrucTPQ+o30
/zOd552oqc78FNi/Uu4kkLIhovuvZiPUpiyNseQjFpWTrnAGj6/CEEaB+/4f
bQJOGRmEqxUze8C9IVQFiazLStruQaEodhV3COHKep/r6PZYlUWVFwL7PMg+
bmFWrpEj3CJ6VFWrRChyDs/isctE5miNo04xMOVCaWOLph4EDXT9JOGzGfo/
wMkHNfcf6I64TUTMMAPdiGLM8W1hXANiDn4cvFiJWpXZ/rEt2fxtDgObkP2c
zeqxPluWXmNN9jU1n30sx3C0fJFIu59vBAKWnaVxOwyV/ey5at6yL63AhoLq
mtTsmjAQyz+Y4qcveKcDUUYz00lccJHIZeOJWp+GH0T3vOSqn16Gs7sgzSNL
KvdvaEgRlQutx+V4neh2SXUl1skhht4q4f5Xv2/hBC40CnVYJqPWHY+AdLnP
YvEK6WGYf6D2HzFYsL/Duy48AQqsI4mqNMveJF/6sdX0SONWEqbBGI2F0WeZ
ns2kwZ0X74vmNwoW9v5HGbuhTcbG9pFsFLXdFuXq0p8o+jtJ3l52wSnARVrW
FjcCU9ZIknq21SJfaWzqDa3msufHJL+/G7Sfzb2aV46CQI6vK+I2+pJaaFN1
w8ABbxqi9uD4J0/PfDv2VE+cjPFwBGvWOAKNLwQFfS3Om7ar3x41KGi5p/QW
7IRYRyBHoeNL1vMmetFdAuABespKtqJjUOetTm8vapM4VRVaPn1LmK+DictM
OBhbjQ/U2Z9FHllDUgyalTIUg8SOIeeBosTSz65cnTV0rngtjbJKMcUJHLgx
MTQtliJZOVjvmcB4KpU8hAKdVU3700K66tYK9jIMWk5yherVNF1N2GYTFhRG
dS6ellUggt4TP44iAj4dRgFygueD3sKv3Lh/6npnvqBrMP1LcLLzMwQYBEMB
lsyc/8mCmXzBaLiXxDyRND9KT2alsuRj0P0fuiAku9lGmOemXfn0B7jxtNWc
7t25S8OYM6dsJA0rqlJ4LfbnCVd+oDth2dKGsGeaOPFeYyXMTXOhgc/fErzq
G+9xhPqVMdyuV2MGjvmK2QvDtGCNa0wJfpstWBDUyOE0u9RQytbjq2CYZ5Vd
FvFwXipmBtLaHY9lFIm6JFLEMCBPIfag1rqAiLt1Kpcu00cwaXEFcHo5PVOO
Z7avQ6AvaugoDw97dK89k35wp+PVFSOd36oWZJ5C+FTm4c5mmkV1E8CfY6Pl
CyEQMqj9u61lNv5+TocILbiv0lmF8CmpIzLnfKITLgUxOUzPCBez65ZdaPPQ
UAn0Z5aZLv/fqrLPm7cylFxQNyF1q28eN1P01k+Z4gwQyD3qkN5ZSvS8vRrQ
uEtgUtFOoq1UKIrQiA18VCM1N+9PPI1g5XO5Fdedi60KaEyC1vtqCJz6JRcF
VAblbW9+F9F7M+/Zuu1T6bCxLPrnWjJbZ1zgr8MvTOoccY2/XPXgXIVWTsbC
wCxJSwejO1X0fdluKla4UeJA3Ow5JQgdv9mPzOYJuyck40SXFzHUbPifZj3w
Ku7bGLIGF+xasO2MudW6MtkKyDOcqZoBataud09RDfsw5uiMxUYU/iTrGT+F
lo5tMOehPdWvZAMBXCI/TJuPE32mbc0W2E+tF35gFpLis4DUWS01ODWZzVTG
uSBCDLOoSrpUW6rgYPB1LaagnHOrhs33V/ohK8CWt8/SFmOtY4qyuAdScq6b
ebGXxMRdNXLDwYfmH3ZHYrTAz9v8nIh81kLik0YPn6dWEVw0Rc3O5io60XjP
TR42fpoGfiWjJK1D31PafkWTvFFSFMWb+TNb3HiT3XTT1uh/gWmWXbQ8YT8e
q9w+G7uzzvI1sBz6IFCJG/y0IOYi7nuweCySkkJ5DNIG0YGJ7ex/hC7foskX
FpWWG2btCCtEXO5+7VheZVolXD7tM/hOAafSIN9GOY657ebaKyI3olFsJmqB
mmqKI6i/3zrN4ZFlaYtM8yCx0JJ8pG/ZV4GdDg74l1jr/kPdW+c8tql1mdIQ
U+v78lUN/HUBsg9klgq+qBR5t7R13XGa354iQyXmMjIL/FXolyDO4g6j7Sb1
S6YznNeqPGYWUv/96OaUXClusv/N5oLR/UQXzgOoH/FAavPHy3lK3lT6Uqr4
dewFnw1TlhcpzdYh+DXysWbPwYq5rbK2sy/xIhd41XCgbFG7G5NAMfzT4AFz
xrmn/uuMwcyiMIvvWq5miZ3GhBzSEMzLj0KD8M+rz7dJJOq+4uX+I8i0jYcv
QVWHTJWOYnDxmd9XnPuJAlz/UAh9ccsH5PwrB80APaVKuu7GAfp2O0FdnTJ+
SynSHUzFK38LI+LA6hjKBTvJDElSf2qwlqUxwIX6KksEc593/mT/9bPPmiga
ikbqRcaAF3HiZ4i/W28qTl/zU/KVG1Cu11JyBiVe4wK+SwX0tI+Vx/Wdsd+D
J+oqDQJp85x3ku6y5A6qYHY627YLRmF2IgAKyH19ri22da2XXYR6BA8JfRKm
rjdZxzwetKgKsZ39VD3QNhM3F+GOnASorIF40zY87iXB28ltwkfEMTrQvUTG
r/ybEBRoShwlBQz6oMLu//g0UAXZKzyy4GGwa/G9NuaJzVrrvMJ0lITcMHZp
t1675Ql707+IE44LhvrwO821uoKdfW+G4tBBdHNSpg0jhsti/N2MBXZnMCrY
RE5GU3WpvpWRHNCqUvPB7jlHLBeAGxecDMZs0/7ntuBqh7yP/7CcFT/1T6tA
YJcht2n6bb6VOGbhzB9ntFkHvtuw7rwKlqJXwVnnZef0mZjp2J4GI404coRm
WvaTNKzPuD/uFeNrB4BcMnCbryKYEQfH3tuubSalcMVlU3csIS35jV9nA84H
Hw/Fw+JuhFOjCTGZ8T/q8NC7La6BYyEqoiVQ9UvBcpMB5ZG8rFBaXUDnoAIF
8CVe6gdQykc6QtqDU1WhF1McIqJDSfo7XaVdG/9tfFXclkO4qBFWdZPRwM6n
YCiK0RNHaLRkuOepTo1EzLUmHzkWj/70fB77fwkTbdLwMWK2r5U1s+89oeJR
NOX2jz51lqTiI9K573dHoAOe1Cli9ON6hO/WEjtZE2GvstlJ+lnbH7y4eH42
qUkvEULWcUo/DZnd1H81Qykci5sQGCPEiCZEm163Qs3Akp1vuOYlsX0kN/Gx
fIZZva3xdWtbEwe3WmG0Efc9I+cERrWEKZb6tCfEoyZsukoh3YDfJQAtb8xc
8m9LFTzGD4Jc9UdvdSxL4rmbL8Y3lhelhpvAzFoDU/j7uBhTefInXK4KIrLi
jUwjEzPbgyWafbEH05cYoWvu5FifhA3jmwIB+9RaKV/8sqH0Igf5inLkOb6H
YmAkmeQU8OS+pc/ZZPpFyQjKDnTLd7gvp1MDSjkIbBL9diSYo2q6kosMxx/k
2jD62VR+FQA8Iejflh5dDb77AWr9i2lZQG7r0UZMNU6fohh2WKCz2hn8G6d6
eIckuUjQtKJspEtOhhsvfUO2UqRHXY7uAEqPx0Zopn846bgyhml2JZN7+2I/
gKq4CHP6p5nfQPXUsMMRWQ27nWK2uJIjHiLV+tzVMAn0GK+7NqD3SxmUgsN8
4L3H9VU0HLw2fRSNa6M2RX4DNVv79Tq/VWtVUFX8EBDSXaMHJLO/VHvSfMsu
07kjOBB+kv4wnDncvtGk/5CY27uqyZztzad3NazJEi6RwjMK2VdpuBG7fQ4B
zTSp/ElTC730IWeR9zd1fTBIW1GiyXdbss2gzw6svJgK5q6ArX/mPwABZ6hI
8lKl97K7GwZLWbBQ2YxZPrPF02OPa2gm9WAEZ34hTJjv8900znA7g1lKnKUR
BjQs3VfoKHRZ/KMyjc2QuAKgGqMU1asqSg8phYXfTX8ejOwg9wycalCDBSZ8
x8j3Srm129UIq/k2VuZ7lW/jOA1BwHyalH5duzYzYp0LUla4LK46Gb0Y5HIb
uSdBVR44lfGpEyhGT/cL3GtkKZGRBuNZQ5UwEdNMAfhlaAEOS9iD2o0UD70Y
D17y6Gg67h/HPlG5GSzAXO9egyKqUW/1VTLEm6MGtYB7XPpxuivLYcEstQ/W
NsE9nZ+ZUcg9Pb8Iuj4SFYGt5N4ciA5jZnDpMOlNDUdVnz9I9hsA3EeTAnGY
2Y5836wiFcT319D8hwOgw3YSvkr3VfHU3VLrx1w13ofbJlhE3ne1TPkNmrWF
zIA9A8cAOHih+1SNhDfHJsQbE28YNDxZi+Hikhzo7k4ILrHP3rhXD0deq/hX
6bC9QgltSxBBJCNYZnC1IjyXLpJQOJB+xLUtoy3pGKVJCuq1C9Ee20PbxtQA
ZHK9aFFW60PON0ZzSWFp2WhA9HY901I1R8cM5hbzWfuHvPuOXRdm89S6Nu9J
djakRlYETgrvad/pQSylJim+/vmLMV/3QS412aIBK81v/zVsRKt8aA+vpC9I
1cwBKBH3WS7Sociqy5DgRK3LngyNkPAiOieYWxW7kQTOVwM32qbafQw8InNB
6AHZ+a7VtGy7NNJ9ezq7dTMnFfnx61KkiRuODXsgrVH6ejTTSBEu9Q4PCRq8
K2uO1FPJHsUeBvSnM2XlanSgm8ThaQqVenZ9cyh7Dj8KHVxEiVcn2U93vH8j
2PUfn5OGgnivUMbmDGTvFYA6qrXGCZGjNwJLnqHhg6yXy1GPPSdAP/SLjx4z
yJc1xzYjjUR0a8P66cRXSz0tnE2JS3+VkbklhpcAAgWcgbVO8lpgwTDnaTaQ
vrKPi2e7GocNvk0p9p/IeEQCVY5qsc8hDx8AezkfTXJ+R86mEfpCoHzFphiT
so9sn7/m6ve3zKH3Ma63gQ0mSCGpaqD1n9nzcoqlsD5qAG1kZeuQIQ0pVKuH
8xYJMMhdB8giyo6f2FAG6SHF3esqPpQdH0tmI0OaWa9PBxEAvuAEWHMKtb4w
kG4AF/zsQiyhG4erj9dsVZZq9ik1Fgfl7gUtVuXx1A6aqBg8MHsFRH7xdTqR
F/NuXSr6NBfjDgP3w5qKtSV9qNys3S5tm3gGPzdWrxnIt6kYF2EVEA2Euyhl
8a0R3EdEOeVITLmq57jq2OrqpOZcIKsz0tF3kcHz+zKZ0oad0/4o4641bQz+
XHVaOeQAhhfT2864ZU8nUMKfmggGEvy004aoZmcb4qYLZ7WFQEQGPpSiieR9
coibTa37JxQ8jCE1ZO2dE8QgUjNjjpeUXncsBP9bG1jWQ7VPJu5Qoh/54aPu
We3P+GIKCQ7wKakiLb5w/d9Ty3FcoIhbBnMpGCszFb74YHLXtFOqzEVVhMGC
yM8DdwipNFziYCOCvAb+a0gi+Ipi2Vmsjy2Ee416VSTgUwCQOB7h6sAwpKH8
pCbh0X7mJXIiftztBaPRtrAXbv857V35kSGundw+AzgL1GO0SASowPQOP/1w
G4vdpsO+rmtW5lPV4IBHITpi1HatQRuCTX7rEg0fR+lJf8eif6p9aX8CJXA1
yYJsokzKHzUnfqIZFNAQtLJbMa9bN+j0NxG8x1AqlGhVd53H4dWtJMGZS2Gr
QD82zUAiclyIBFXZQ6Lxsi3aOF98DPfEmTUmdoRnQhQMUCxY3VLda9KIOjZ8
LdYMf68zU0JbS59TYKLbwBJm4i9dbMWJYvMcqbOtitnG23K6qponuw/cwPeJ
DqzZ+S9/mJ1ye+wp/9U4fbfgZh5sxEue15K/4t+7hlJI7Qgyk4dqEp8itwqL
tYUMpKRY9kteBLOPwCIFvNqQ9F76zh9LW4iP6x5THMsCdZ9pryC6RmDzZ8XG
HIiYqOtbvHB7NtkiixLehapDZRbX/BnJKlM3haSCyUjsNoMTfWirZnat+ALk
0dkuPiQsskUuo3HK+lwvp9rH31UodfVTBb1RevBnyPBRrL8VYSiFuXetJBue
JJR9tlDUbet+lBnQAiFSC/TO+je3O3hLmTUb4Zl4Gme3pVJfh4CALbGQ9LDC
6y8bg74PYYJQObCfRPiyt3MCz0yA6qEAQGWi588y7mVhD4u2nwNIdrSVUwqT
x/7wESbqO+O8oBFqUfJw3NKekqamObWYFhxI2eIkfOQtMgiKFGBJvVYcjior
yaDRvahJ2lqSdfz41lACowcTjW2Iqlageb62NRIsB2EA0o+7vQw/xSCvv5xJ
HDeMKR4dKpkc+Jdm0iftxBi4dyxA5bEHppr1+UXTXF4mDS1J1QT2xpBmvf+u
QFEVdqGGZ7yWH5HfZAQ7UHHj6k3t7hNuwQyi4ZQSN5elkUF+iSPMcRi06iAf
zF78+z8fg4NuEMU7SZj29hInZq2idxr3SAps8Z1W9pzv7Y83zOKAsBQdLB2Z
VOS+y4TXxiVo5dasmN0kMPSh7VwcMSYQCBZN1p7tJToyD4kgWsplboE3RGjw
DI8IDQEKc2zmOcP7lJJIiB6ZoAVXI4y2l7mTCP+IKFR3na9cMpHyXN/T9DWO
lIlm+8P0z7G6z7mm120988hGpdXdIfvuvRZxlh0HQZHIkOE6RtYEhpQYpGEE
udTTNDVqqOBf+e7uQdC46UAMnFwmKTPjb8uGa2aUExs1Cm0qH5jlJkillr71
I7ygM+FZ2WKmS4n1lbbp9eC3cSsGRkCVVOcDJ2ECW1348dTRpAVgJz9eWLhi
FdukmtKXhRnZS8IFP8+zdUPSKV2d1TVjlZ47imZbwHkg4mzfeekfQ63RW75f
x3gEwVk53bjOMqRwuxTcDD+ghUSQbnPR/OkTubOCuF+5D7kG+2M0RChSFR25
7iUYw4neQH/vfRQ+D/JJrGihaR5yV8BI5ayHwdTcnDv1fV630fYDcI2FBzxv
3AvItjnYR0ra32yN0l/13rgZptK1y4uLGCcAlpjNTQNeyCxoGA7V6ljIzcOj
GIdn41p9APMnpW2HzMfdjmN9jaHg52Le7SqrSFhlmLm9Kk//u9BpzxHh3J3c
ZLhUWUXz7wzJDLdQVSsleEAkpVmviwhqLRJH1THp9pQ+/xrWcylFRiC3/eWz
nCxtbxO+ZLXxue0DviF2rkowgTvM5zg7V7geJuVMFdUnnoF5Zn740wHr2D0J
CMz+VlDHG73D5c63rDMTF6ZqiLN8iklf7WvQ++wdmqN3FGcPgAWwvPFR5Zy5
IJdGVmkfy4BtCqnevfPCVa4jxGgJ/Tp015zsWlZw2ietDLm4lNJIrA1owTim
2Ma221pEm3yQbIHrACHqN6iufIilgFSxg8sn9b2tJyYiHGDtUusBCz0Frlph
/nMKlnqsqEbL+uOLE3KQLDpfstSndAVF7LUZMG9lfTOK/AI9WXVMpMZzUKFQ
9BUIYAaSrhNjRuZWbNc1luRIeHyTg5c49WdbtOHECWw+n6JNp3p2hVkjek3F
waQANn0288mQCKPkpzzm7vs8HHZCYKzvpk+DqGa5c1bm5w3O/vhyVCqcKVJ6
O+3L2OHd6kSdqxMMMDpz8XBNNtMqxeCKdfHiucbijM+uM5Hr6zIGziZQaWZ6
VonrqikOex2n9Zzo46x/ZCjUD6PRTPZFHsmfjThZfLGZPNo6/O7jDlwSzc/z
ZmGfFlazwiips6ZqO4QF+nl+9bctBsYOuok0FlDWtEwmouCJBPaZSQ2SFxRz
6ESfwIMIzO56uXoYL8av77i9jrPpNvrgQUyGQqlGUH5F+ce0t24lGkQAHf2T
BmLs6Ie0lYKCbw+X2nHWcj1JnY8KhyV0MaJ7X3BQBp/WPgFgbQcPWErum5h7
ZrcYwMOKEqrQuGAZ/48bHjtTyxcQWZ0dLhVOVtquwUwy1H+zBzFNvMuX5+Tc
jZg7YDUlulIBbV6EkNQt59FASeIFvMCJNEiBtl9fW9uQ016zuWI8NvPIhPli
zuneYP3eGe9yOyz3hEEaSk0jgUzqn1UxIbN7scND2mQLNmGMO1FuzZJ8BDEk
llPREyCPHv7tlGmlkCNTYZxsC8F91FjErNN2E/RvnzlZsnhpEgyGJ+xvXuGV
ac5Jwc9gFmalJlJtAk1xPbOymI6bOJjxUlCsJV0eTIjz182+gH+IgEESSCfZ
Cj0MRzQqnTU1TGFkRltjzjYqPTY1/TGrZAEx1pQ22d04b4fB5f8/MO8j7VyR
NgQ0xp7q+6OUsk6VsAwQ1+GHCCc+tRnQyA2DxL9Vr2xldl8lE4p2ELah/ERl
lpWd/EQb9U75f9G1YO8M36f0P5wQRMyaHTe3xYNnC01xzFlz8sY3jq+jm2p8
91jS5gE+wq+ngzFYiUtlHGdvfN8gnP8FEHN0wLJ8z+RzdFrKrerpjI4q6PnN
RBaHuvp/uyKezAcT66SX+Rlhs7X1y3EOls7u31uLTrkBKFBtaydFC/CECsoV
3lvcATu77F6TU9+qz0Zq78eR5wom1TWWk9ozdiMjvjWqWmKlR9APPaUQDFYL
wvsOOMmO4z0SNRGOdjZ7HpQCAiHQmG3BB63BXIccf+zS9vUsRiDRoEwgj0qI
KXe5YTDIS64JjCTWGmPfAFnarwvWytqX8OKsqw4nexm2iD745i8+dXVn5sE/
nwgMvt1KLd3zeokl+G1bO6Ka+ls/nyhGp/xui/u7myqEtme0BWSLaDNQM9JK
Mk9J1HnRwoL5L0wkY99ABkBhbCV/4CNxLsfqEe998iEk2SXhWa2U8OWBWjl2
Q154QYM9wbucrQB3FQbtptqKPUvCMlqRoNBLmFJ4yP0QlsRPc91LGjBjY9NJ
z4+0eLzu9W4tYo384ROnEw3Q+NwUVZf+xOk3qS+lmxsCHYE3RQi2uhngcNZm
+q3yODhpVcgZQidBpT+aA9C0uYAhb0+I+N+Yzb2n19jT74A40wby86ncaXCr
SvgjO9rYHgVXTDVFJfQvQG5fC9GX/pKvjxMUrFE46eUI9cjVPhUrd+4r66EY
nUZ7Ubh3Ld1mJ28fWWWa2c0idOVLYJXBZ986PUJ4YH660VH7AoxJu1XUxDcT
xPesaL1wKDLIvgwff0uQUe/cU6ZYVt+Pv6sMVIEhsbZsc7JA0mFFOjmkMUro
81gQw7+2ZGzNsRWY8K0GLtQKV1Httq5+/1Zn0bWKSUVlDG00J2FTzIVuYWjE
p4/5vZ/PRWZqH7Py4yJPrXXwAc04ZylMNakw/f809ptFJUQKAvtQE3uDDSfW
ZqfhNvzBbMfF39GGhJPU36+TAMZPPowJJAfcWy+l6SvQlVamxhSfSsU/YBVF
rxQR6eoSdjsI6Nkvy5/OO0J18wwiV6jQXkjZ

`pragma protect end_protected
