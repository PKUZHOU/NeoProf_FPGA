// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
UTUgs788GjXW6qi0apobtnJOdrvoJapYdWqSMGy9BQbViuF9C5Cx1SQNUgTErTr1nBMpUHH8yvie
QIwkhAe9lLkQB0qrYBLTVfv1JqB/7y4bJlJaCmpbaVMBmaEddkNcd8vODBXNtEYfXCiwWJf7KM3r
I30p3DFDOByu3jQ50xPkOQlnr7mx5tj0A63zDWSKxPv5cyKA1OS1CR7ToXo+TKiBAK6pKqPLyIve
cM1bgB/PP56JaTkbk30XiKhcmCe259wkLvch0GvwplAkAnjReqCuWjtviLdzMpTZ/IOD7VNPY2rN
QL3oNlenw9+MRox8OtvAs+3oWvNf2Naz7lSnNg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 2160)
I8vCXW4ie0E8LouSqXviBshdFP6KG5QjbaIO3aGZkC0vHtGfKeu0WbUYkTP6soPybGHf0/Bk2MBW
fBS+K8APRRVsMG0nMl6xt/sj9eEXL7w1tEot1Qs03QcRkIKoK1ahOI6ubYP7BswH+0pkNXICM+3O
mI+W5geJUIUQoEFcts6YtW8AnGPn9nU4ZygLLriYVu+GDjZgMdczxrubDmU/foR0hwR2E0B1G+Mw
WgFzI6TSiOpIBn4c/PTg/QQZ0sqAFdakDz6PEecOknN8O1sqX9K+MM5kv29KNP8IWq3TZLWJ4sFt
Ia7lduCmy+3wWr1LZ/evg+DMzoYcyTrGq/zOJOzjE4ZkFS+1y9sHo6GRju36ndS1nE4+ccE+oSR7
rVpHmZTx6ZljjeYL1KyJ1y/KKc3GxxzQyZ0p/iNI4fryTV1BZOWv7ig0ND0wLtKU35+nYDij2Qrd
OeffneOvQhGqB3CN9ZOXPkN9dCNXdhFZVGsw9IQF+4mLcDPOmY4BjNnxVSL4TALlQlRqe/uXj16H
4a//9See1T3Z+T1IafxwP6lJCwzTArstPB3dv+iK/mC4XimYxe3w2QOPD/BiOpoquVB/gKnW5QFA
R3+x53G7+OOtkTYZoSLrt+P95oBRGz5d9txqAgnB7cOMxT6keY+3uyzrV+UQURdpT8cBAr8dEgUd
Qrl70Ga76yUZWfVpqb31gZnsbi4eqsQpeBYS1Io0casXI1lW7TxIPajyydtWSx/giTmvHw4OSw4W
+Sy/PdlpWi8R8uUl7mI32plHi6B1BNqJuWfl6rnwL2PBictXRX7dXxQ4JckGyKOM2Bp11Nsw1Y9W
huffaCgqWhJtLDgdSj94Oj1F0TbX5A+PHZxJDo6WCJgKjyj56iRZX1USCqfp6/Vj1GtpbNL/70UY
+LyWzx/D10zIO6q+FlIp08EiH/geRcgSYj1vyaVurg5m4nKAQ+mLYxl0qYYVthlu8BHRS1+4OAK+
n7Zqr/6qEPFlK02+dxRq5PIByTmbQ/1V1u8HZcW5ALZ7uv7xU3DjsJKFjQCYpgBQ0ZqKznxIrpls
q3pdyqqobWgLQv4eeomuULpyyVBbHtiwAKn2cU+ZEBo0U8AgzC5ZXsh9qVUVGEBGjyYIoA5MAV3o
71DRcIYYjtXjOeeHXPSN8WG4XM5Sko0GaYW7UNtJBC1RVTSx+iGpw4YnHQTbHEmHAT+M5ZP83GeK
LjQ5MCXNaLycmxJtUNYNW5RtD/h1I3AjIdawSic5rzCYf8ansEPxoC+2DjC4lQKNd1A9vicn6RL2
YwewqQfyCgpqgVEk+E0KvtNSqU0yRcXqk7rQX4EZSHiDScMpoD3tEnA1qT88JKqo/5a3YEPvcvYh
cf6uwukRs09hWQa66+D0GZsYvuKrhgT9j1IiK7LzE9noWqmkCYEIkhXhuNm9cNknyN6OkeyPnZjH
LeFlOlZ49rWYb5vXXJpAM1Fk4/Vg/5gzh8yHBQ5X4UXuDZ3I/TsuwTMmG1ZSLEt5JKgRfljP0/5D
MpdO4pX/5/EKUzsHc/xHdekfYJJKQHGaeMxRiWzFPLed7LZKQ8zdIctwKyMBkdM9bTf5OsDII+Vq
xDB3u4Ch7pNbIEqwoNjS+RkGmhRvkeTe7yBvSpXADCHPiECB23gnqGOM4kONTB9zXthr1xW4ytK3
hShFF0n87Oqg5Cntx4uatvKk+sC0mnEoEj/H1QjaGmRoHmP97hQcHMGvvb0TcomjTZIyuihA8p4j
pwyPof6XOqExSY8NX6ghFc4G1cCily5n9wv64pbFB6SM2syM9N+AFGILG1dEzIIvjESyf9rFKPW3
byU5ggszWJyfMTxtkUHYngB6u6kX1I2bElad7L2KgFUTAZd2RtyDhkZA8Nbh1fw2QTiZbOOFN3vZ
uLAdLF6o42XE1YRzakGJ+WidnbGySK/hDkNCy6mZO74vNR5CjVVKBRyLxyuXxNZlhgXqh0XJhQPx
uZiv871t4413AymRV2Schi/7eryFqDFz+H2X1i898GWkTZRU7oegWyB8bnTItuehjrCZy1Eybrwl
xaHFXgzQlPHHJ9PWrjuDbvPo3ueRa6oRY8mbCuGRvvj5afpzRninvJh207bl1b/PdlQKkVBxjSEy
vzZCq2MTv+9guxY5YK49++3s58IRknVNPuU6/R+/VkjHyMGLgiNVuiBS1jtOvhbdsIBdlEDAQE0O
bWuQYxGSXfAICyoxCt/BKsKMJNFXR+lV2hQTRGrZfrD1YDZp6bGXfJ1e+ZmJPcKjYmu/08yVCPeI
PzX2/gnjUyF5DyoCoHk5yStsKVXQnm9ysVPdiHbPrFu6hfIQ9T+h94cnoELexJuLox2FpGpwIo6+
N8eB5eCoBAkDcZGEtJvsHCrCQ+H3CgdQS7L7Ai1LbL2i8+CIwD5nqDyP302ojQ4Vo7z4ukNR6b4z
/xN8L+cy0C/MVEcFw+4eGQAmt5cJUlGiRmrvWLjFzg46u5FZOzyI7RLAtuwHsGlwdolWa4iQhyYM
Z1fE1w6uuhTj5dkzKZj6GD+bm5rHT2BfzwtCXqoxRfhL/wV0AnTMcLlLIyAWAdQoNCLWHBLISRyc
S9lKhv7w9Q33NJithVRDhJ80sJiy6kEQfdwzAHx6dttwGGFcg8ybC7BzXRkJyeqtiuIbCHwXw5vE
RE/ipfYn29xsnCZ9rQ6zPMw4B1eJFOyPahuBHQdIkONxkID265U4oOfcFXs34H+CslsgwnNii296
mK9cM1YdACXGXHGZIPS+NRgg1LBeJNcCKyP7me/+dbrepCmujvRC9aSct5LhfFm9UODQfeFDAOBC
wU4fwsgBodtG5xogmzN2jc+9wljjXBhOlw/VCM39o1QitudpCqEXyDDu8hGF1nWSe9fT
`pragma protect end_protected
