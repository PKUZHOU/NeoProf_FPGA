// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
exfycD8COq4pcteM7HZ0FSFlwx5N2sH3OGTigueccZj/rkVB7zE5E9nbkInlT0jO
v7izzmpzaHe/dVMp08t3Zfwtts0lsMZTnCUjaji49YoibzZyTEFDgV/VgnImpbB/
iBkFLAwAHKMKhJtRGfOY7OVcNZbd2SisLo1PzkZjmqXjhup5rCFVBg==
//pragma protect end_key_block
//pragma protect digest_block
sB+b2daELRJ0iKJuCLdeGxnM7mc=
//pragma protect end_digest_block
//pragma protect data_block
Lf34TiCPcYFlw1J0meWV83Nm5a7/RDDgBIX1glJzjLsePf9bAqeDoE+7hj/GxtPJ
obOlCUOH8MTe/tlEqX4CDrtoUSXAVxFVEf1S8bCTRT7eAwkrWwfMh3WVfxY0+7hq
NrEZyOs0n2XvBPip4T9uv41RD99RnFhXNYEijGytkvM2N5JA0nsAgiFxFUw5gLIy
5ReVBKY+e/FIo2/G5Pd0PuUiJFLwZUWcGkzYIOPhv+R4AuBn6WDI2FgHYFa620o6
r7mKGZ2fcI9Ou1h9epM7DpWZT0mlMTXIquxd2jEfGOZQKRPDPTsVOdoor/jrRXX0
NVl/lOdDZrsHbkEcsLSoc8LPsSH4z3dSVdFu7K74wrfP6gpENVZRtYf8A7/zk7OI
sKSjYLOcpu600v/oc1K75fEIxQ0wHY26TzXIolShn0ocPv3CP/2yG0xy9NSmirzh
MGkCM1J7RXSgNTV61pBcLamWNcrfSRkGL3ZqCfJ/Ajfin+Zi8ZrXdNhYQNmfxkRA
TbTZpRNd4UVS0EZlixCjxvFAra15GGU4LMKT0CcRfHSG8MUHVz5ZGsmXhU4HunAA
zV4ZoLTYFiS0tfUwxAXpAxkkV1y22aqqY2TJv85ctVxBWG4kLTiEh+6Tze+gHWNn
8PGk7pxvzVNSHdk/XL8ttxNvenoZKbsnXsxLCJedLbOiNHOi9LlHVAUNpx3/Qxyf
avP0dG9NEQLDJAFXRXsjTCAPF43gWyS79AKaAYsG27If0AsO7ensDFE5UGHXlt9e
bEaEsZ56ChRvRjSHa1eKIO+hi93ItQ4oysYtpn7X6gdS6X0enfMtOqszjpoB6KYB
eheL1ab+3GxHid0oTds6XPlktpEvqc3qGOAbvdMujODi5eg+VgeQtKgLsF7ny8Om
w9c/1JEx4bMhybycXn4mgW2kcVb1Itzq90sBocR/5iTIq+/qI5OPfI1HhCE2bbgq
puIspuYwFLcuWMDF31JnFgEtvUYprpqW7L9rNnHTjr0FTGgBuTAq4rZSPN7hK32V
o+rw1CigtSj4ICi3Ut/JDkCnDxlXZHPcmRZ3ke8VuT6uavbvYFv5SnXEXqSoGIgR
6g2Uz1Eu35Ha2itqo7vneDmiJQ64z3OYVGlGQl/rMVzRPYEGUkFzXnonhPvTJIUG
EubR5xqfFKYLeTqJ4y7x1aNkzDqt9cZyKz7xbLL0B5gIsgPImzoqvchh2rvv5Vws
6Mj71Y5VTm6C16ZhhBwr+ekVYe8rkKeF6SSl6vJhtB2KFeuQZzoZZq5y2vBAfXDF
ikftubu4vIeGHQCXD1HVy+zznN3SKgH4L4+quvtknTHA2/3zjKrp7S4qjpbG9lok
AsgsnAOT/9K1XKVxoQpTLluyLrrIJGxplnxfwFcIK0131BlUdBhJbngNbaQAKMP4
hWZ58heIo0BZ3mDanLNi2reXcQgqPXXSh87Gdb/2MR20wjiLwygokBTYa9py4N0r
sMGRI8NAsjgjZHMLxWry+BiEh75JFxGpncpOJ3X7KJActW8YuFkphGEaWAnCx63S
OuFXeNdiHdm0V2VI+vsD/4BokSmZd2gQAptvxUni8u+1H4gGxAqrgVOSDPbiAJwf
EqybfY+FIog07lDDzx59gzjOGqA0/FSYw44ONQK6KUnSPMmAOQN+yjgNa/ou1+OT
0tMG0b0rfEIlvH9BWL6YnuZ2PEoIYhMxCRbP9Q1TFUsKzutb1j/MVFjUZwSQcIPb
a6CtZTY/AK1Mmsvbw2mAdFUWCHRXTSsbSoUiyCWh/bkkr+lJW6o2XQd3bURze4yB
BkVHP2WLXb4ZBv+I+NbtTwvLecgWEaFE6TSXIUdilcL4+y0AI7PLk0EYobKAmGxv
Mb5b+fOOPfmU2/FQZCWpBRD3DpX5YRzD8Wplwm7nlK7gC5wibJwLQ9msGOaRFWsJ
KSbAx6n/tzGgM5xKS6KNnSwzVicG9VN6xuZcxxuVlosvWH+MueZ9qpFJgl/yFy3v
qcVEYpMtXL53W3b4szJQQy2eSQWP8UObWAMzsRGhb2GmdpV+qM6to557eoao6T2n
TUjNlOFp7SchGAMGeitnksVydSoXx9yhUoE+KTg04M2R15258CeMxthqhr6D5thh
5bXNaZX+Kczu7iuQoXiQ9bY89v0fZECOlF/0GIUrF3fA/roTExDi75QALaJ2Wpb8
7wOIvUx/y6mK3ZCqwiJ+sUAKZ5YIgaucCA200mgccc73oPKLsFWA8HI3d2vSV8ej
i1N7mzXU8elPH4WPpl+h4IPAYa5sI4kNvUvGRiabyFCLTRoXep+gHHf6bLDVLqcU
zMBTWW5l17EAX9LFB2/5Bwu3XpZ3h6ET1jFhNQz6FUmDDT1gGAjj4AbkiJK4SJZV
sj+B2IIUsR9xEYAjc1cXBxeAPzLiyBw2jlk9ztGJnTlNKKxcL7uoUFGexEN51gVE
lUSl4wfF25RGEaOqLsXrX/l5Nj6Iznkb9Wkh0q0uk+zODKadPWyS40L7WLPR0HqW
I8jtcxQNWFdplqjRi/PmZcTzk3MLc84WT7O9EXDjzBjPUwal73lKktJAWDFuwsBa
fOtNJpecleGhGXsPrPNj3MzEdb2Z51UIfsvRxJ4qgTW31MK3883+eXrP+O8FmaXk
tVdmxFiVDkrPl4ZeR+V4VPGBrtfTpcmwyTpK5lxA6DR7Tc5Rd7LdCFD1CgZJ1dTF
22OpVzyXImPx9zP3BQ2Rx/oU2BuANl+vsfLfGNDeC36pzHidt49CxnqPfNGQ/jsa
1dyxRongxguty1nCNR5loGs9xg2VfssNkcxoSeO6DgXSEHkl7ZWP9MgkKjXpWiU8
5vonZe8rCJZpz/y+22/DmQsPapa741u3WlT9vjxuvLVXXfWNPw2t0SSugvtkBRN3
hzJPj+oAHC0tbBOmrUux6C0ZtOa8KZ+gBTnO+UNrsKYm6rhPRE+gL9CkXslurM73
NXrD/Br2SEgjbukw2a7E8BMaNTduy/7qiJ15fyaJfMllSlRpXYdv3LWn/0+CmPnk
bqLydl47i1zeb0Nq+Yo8weQra4R1wwRmfd1HALt/T78Z8qmRoIViw1gcgqTo+J+n
W7fgimWODocDDOKCYoDQJQ88QWfm870Wl1AhGD8k3ZGFg+J+GsKecOshVUjtKQnc
xUfn4O4gs+ohWXnjpwnvOZs+ql/dTbZklRfE7PFCcwlYYV3jB76wYL2yp6vJfewL
5lxquDu08YsgpWiR/0fs5wsW/kTkVsp2nFJMKpGfb5Ci3QSXeiLOfqzYkw2vC2Az
7WNg+zXhSzNxQi99WNeMHiIeW8TSFJTC5gEdbLdnK1OMWB/T9hlvGZTVbn1PFtQK
UKF5heYdzS3XSVRxiQ6gszUmmHP6Tgcoc3bEGis5S/61HqQoQMqyEmzILCI+Q10d
yRBvUGghLsrHpkwUcuh8TAF2cChJcXIopcIYjrStwSSlG/y/OzAXHU+E+IXqwM5k
IurKooW3KQc5gLHlLq5SCn4LHN7an2OBaWqAw5K1JGBRTdUGOlFXksjacXIe5DuW
z+EK/nmpC25uGQjsAurFaCplQ7jFf28wdjSA6yEUTx0dQ+eomp1Ix8/i2c+oBu9S
jcwyL0nhueWRXKx9Rs74kHQRPZhX3itSaas+Fz8DXyuw7xszEM7PjFGcqRogcv0v
S9AjV3aHrzy+yS5s6RynPzwdPZi+cKTGM8onWJ/qXVozHQnMxBbrCu6Cb28AACpX
Ntb8//clVMbahYUa0eQK0ATfRcASLju1UG5uEQm0WZ4bqfPlZ5DGc4Fo1YXHKMW1
KiwkKbF0EOk7tGuapMnbXO6V4RHJTSVYzel5XzzIBBp1a06KD4Bhc/kb81SM3QJH
nAY1JJKAfnAeLMBi2TEbgMb3ZlZXhFg7Rmiwi5Roxj0De3p5DBLaVNz0FOiz5Wtz
ri081ZDv2qxW5pjIJTTpaWwoOZl/gr4QJc8+AcA2tkaYwyF8AAcVPPgHHNQ2iIxX
Bb3xM8AF4+kLjNEnyntZpIOxbciNLzrHWmFCHDOQ1VF6uz+Q5idZ1m1c/cfDeJq5
VIqgaK34gxpsC2vHL6jKndLwXZz70EI6vBQccjrNVeTHruWvGPVDUCWSRu5cuzMu
CiaI4JNgutq9LS6uQ+HReQ9lPpxD1atWX/b+daNid5/NVi6oDPp+2j4+nnij0ELL
dVBJNVPCuzSdj7cC/rOhjccS8qazQ4PrCDNBVfxo4Qlt99jN364K/8lG/6lSAmNx
uEkw5ZYnfVcu2oYQsXskDYph3QL3ebGh5RgFEPeCrHfeifazlYkUWrERKsqr00Nr
J8KSi2pdKvABT6ihi1cSK3A7BxEFgxtMmHCBm8B/2RxwvTZvmAw6cbwPPIzaYpW1
+LVkMu4ls/117T/imiJVhgtYByjmsCZRRGkbMtzRsEeNY+oDeW+Wc/eGxnKNrhg6
76txnkIAmwsB4itISHFca84Ppoy9pIXUJ0zYb+nf0nOzaV5m14cdHo+mIoCc+4wZ
FTZrMjOVcivGTiK8WN3qVXhSDdpV1asVItQZ3ftbyHPd+lTmrWffaX7KzCMeLTXO
D6UPBEFkMDPQ4IGp013N+5KyV0jel0apwqXj+7NmkDm8pJYYP03VkmzbyAUubR73
hlS8Pz1Y6g8TMmTqvUYD8zcDDMh2ioMQTErTKWwblyXOC83BSvLoF1KJG54wohUJ
g/ghd9yf96AgNRmyalRw6CXauNFSgDjNdLRQ/uOL5Ddx14U+DwFAfBKGfKbAJfJi
ZikULYSGdK139fvQEKEkXHkbG94yb46IVn4AO2r4hav+OM0yKpGOk48I3EPPxbwV
824r+/Q53zzf0GyfzpT8HEuBMZwe6Cs84fJOVbYNd3pkCn2Z6+R+9VJGEtZcmcBO
Tb6AXbVBRQrxYFDz5YAj5jZ1zHr9otUmdHnZxjN9pl+ay6OeBmMUyUG3XDVsrmJi
A7WXBtR/ZFOqE9cKV/ETcSLjgFYdTLIdhleBn3AnOQL354++Vd6qEBmwZMs2CB5v
jORB/qTQQkHCokJuAuZrgr7DhvhR6ra2GQdRkoqkrK/FOsKqSjJLNVza6tCYTM1b
LDfFkbb0OKOEhpYgwjB3Ju+Sb6jSZf2RLMgJ43AZlB4j+TsyvChmZ56cwrhu0Bsz
Th+zWnC9mJJUsV5BXA7MDzfo53VFQ5lfLrgJFkC7Ad4gVU/RYDR7PA6YDT0jwQGU
B9WdS5lTXexBzoAPJKFHfstnKzSpqszL2loRVqbjwaE3nGj5PAPK7n97KbE+x+Hg
FSUIW+LMbFwE/Lc+iyqKHQUTUJBWIBdqUXlPttuQtMMf1a+m7p5f1KBp8C2o5jjh
OXEvPt8DcbtQd4/cy1zbEL1MV76cvendL7Snnobj8A4NAv5DEDfxeERAu8Tcoq7k
l/SNXpt4RBq2ixq/f922dS40PoKjBQ8igCHez6mP0e9ceI7Jy94yY15c71wdl966
FaGgwFm7tQEnCuPdJpOakyvoyu/Db+mONnL3eSgyv9oEM6ado4JH0m7cIQRZigFZ
vaZv4rrpkNskGMI/lpqJat9PtgJq2yZ0FlHe54dGnutVAALafsGk++Jal3BNDTW9
UDCRZl50Teyl9WLdMotrKA4V/O8EjV4tQw93HFUxKR/BBN9eKJkwsHSO0QcFDkpO
+qrczxYnnRfgJb8CqvG9gVNKOuE8h+0xaIcgDohVI7ycah0ak4GXqBsjAoz2oIQF
2KO6llV5X/zb/489vQm5CKiunX0kv6G3hcd9gQFr4ISjJ10x3niUigXC2EZPDVzB
sRcxkhoD9b+q6Ln7VQPf000sI3b0Mzd2HOboRA2aj7DQVgmKNrUzDu8ie6VLoqSc
qOhxzXCshoeWoh+qZOHxeNrBJ/teUgh0XTHfA1tRL/5EnXJZAalZkL8ltk8SvtgC
fSnoNw2LDWs7mWFukLdfTdCICjbxS32tl5QPCystx6Mi1yuFkkq2snslu0XadLOw
UJtxi9y6hmFpgX6GNQZabPFfF5bve1jBvjcw4v4um7ywMnVLE6pl+ZuIAWycO6RB
GdjzQOPWluagCnt49vRWAzj57E4/eRICkDTff6goYpO50xznvY3lYZMPFKrRsf3g
d+zrsZTG+PSRAH6DVvHwEzQ5auvydeHBI9ep+6Dn+DjKxjV6Zhduw86t4Jni7XTy
b4VBTvme0NUr6X8sQoZSaRCbBnOhc0CJHQqYnchwZXDXxb0cJ9w9i1SoirV7lyZy
bQlnSftlQADEsM4D0krAlm1kEPlf/7g+G2R5XtwQxMOFp2M7cNuIa/6XK2DEoPRA
yT6f4ohXnGDaaSoqyFrdMQgs8DXsJ1RL/N+/4ayNZASaNnZV2JzfkCTwRKvxSSes
/cyq7yAwH92qk9lrnZ7ZXEl0stTT3zN5TNIHCBsR/lZc3iR2XL0L7B2iNFxPevZq
Dvm8QH+6Yj04Ldx+SVR5i3pIHklz0413ZHfTQc2I76FwwY7WC4pBSpGGRR08+jgs
zCQL5T5z67OriUEylVPo5OyYmltfNwFpD5jJ89O9rcB1eXNH/LlVc1V41n3jZqh0
DN1Df6WIMgbvlno1/r7HamVuG1gnMc7DZXMtHw2C4eXPDhHJqvacUhyYnFhsp5eh
wmN4CECQnv+UDqju4NcImMNmxE/0zd2p7vQbGkytRnwjpNSVFCe1cvY18eZgHG/p
KKrmWjeKYiVVAOzgxc7IbKwbjskudENcwKFMVL6PcaimM42zRLnMiwFSnOjAm9bi
htI/MNYa6r/ifmGFfVr+i9BKwbAhHHuzjDhZP9ZZvMBMm+qmIP6XQIbI/gpWLBTW
fVbhTrmwk5oRi7sO5i9r9LKJAYilbCQv6/76F2bgTDb6utimk0aauILNHydlR6yJ
c+Msmc7I4TlBSQzg+DQLPV/jTi7KOVRori5FufellRyuw0NXna5+PCjMRW+ahmi/
Ec5cC1Wvka9E2UtayiyIjoGJbSLqg3fMlZYq0+4r4ZacTBgTEpxEqEn6d96lYbKs
MhKSTzbdRIhKezm04xjR2sorDFX8RWas2+o6EjbooSqWzboqNg6HhaKyFnQD6Hfz
VZZ9h1WX5BLpFo44NSatG2Z7UmsnZCILBpJ0+4HBJc4iWYRxgucuiQ65KBq7Uvfr
XrTrpDEJwvgKl2CE6qiBwPVJaQYyalPdDLnga7zUezHVvRH7u7mIxCC+MOhLotc2
VtpBFdmFWKhjN4z/OkSh/B6hcB7KgQ3trBQuev2azkHf7ffTh5NOGloISpYY/nQf
ox1VAHyWdENUBJzSHSV/xYOCR/hjxwpxU/88mydFVrGEGXOesP7J0AmU/vLYuoIA
lknAwmPJA8dxUfMUvZUGztrnhzO5Z0apxOkWRq7ox3Vzb01g52+Q33m5s9/p9S/k
teV5yh+EcbYGqRgXeppgzk4T4Y6FTqM9j5IX5FcTa1FQXgmHyuJzq2ODy9MTsUXR
NMmHMvNMARyKyOI3abm9hUwnIRPmjTnvDtSe60Ucz61wjAiEWZRBcez/E+VCjc0w
b0JbUtyb4NXcNJOXHCi2o63s4h2Bhu8O9obrMz641Mepeet77+GBv1YFoJjnx10+
DlPfEY0tP8t9MA/vqzr3wQfFu84spEuxnnZE+hIFZGM2H747HCZ0ZQXJpiz3Q+EG
PUq4epRwXiOd0/19rQmsppE5foeX6IEXUZwfMxIWPLpw6+PlM4T8J/BEtcD3zgG1
FBvg0akiZ86ibv5QF760YebFLPQI292ynIC2AK0Szl7oNGMoGqtKzie/LygmgQgL
vguaLMyoHOk3AxlvwNWq/kQZXUl8iRAqW0xyOf7sSMBd+LRa27PA//HmIfzflq1M
oORdqkZyHmvDZSFxwwqFrHu8X1Ce8H7yDkbOI2ghj1ZNTgAQLbv4PC4K3fwjo02j
jDTfQp0NwqSOeQ50zrKKIm5cGe6WYyc76xsWz+PZQxP0qY24ZJwF+pWetR/UgqBJ
9u1rW7VHxyV+5uikd2YChdPJZ+fm1CcziyV2wpM65HqZ13TQKjBVDiSZ3lcR5I4t
T3iCaOD8LPjx9oqswi0CFZHC143BV0vdU8BcNe3dF2lIhQngWE9bPS1cxOQmxS1v
ajr3sZ4TwwM6iKl4bk/w3/KcYy2LcGgT3Jb0s6w3Iy+x7VkD6gzUaTzUv9LWdFFk
HykHj/Ok9hNDEE3kQx1CVHV8zgfNNiFxjjkoFFf5GZyMXnEjOHkcT0D5Pw2A6hNW
4R2gu3/VZE8hpv5A1MAXuyvk67PsEkcX8UrxRQNG65FzQzl+kwwsPYD7wEKl21cA
xPrZVaGSPvKjgczE80JsdmjjngybROp/dL10N1hVY1zkykmIL2C0DRRXM2oSPZdO
Fow6r8bD5PmXj+BnowZ3WAFsl7WYiCud2bdVGkyK73BB17I/V+/NiWGRqkLoROWv
QYljQbDeuX1h1f78rYLVZP1H/hESlIoYk32n2migSiprjKgRzRtQuTgehLZ5aTIF
M+bjx7lzPB7vI1VcYiSYVn4ryYJ7QJvXRT6PYcDY4+EsZpNvTt3AqHePmCpwHrkE
UVyHccMb+6Vp/NEUU/zypCtZmkYXwvNnicfth+t3pSAa1MqYGSJfHZBLI+3wO7El
NA/zF+DU9MS8sfNa0gnY28vXoWSic+ZcRSRTIDAo6ffeGBdbwE84+3QH6HcJDAqw
Nl6FIQE11wI4mfikf2+aBNydTowrFcRwHwzqNM6h2+/1b55797kOk74hpAOWT8I/
yPoQWRgHitDVZE2rpdE3ok7Xzv/oyOzo9SB4OhKnzFVNoA0ag+E01ka9JOqXqfNr
RELlp6FUnHiFkymxzQaK6uonZeHjFdAm2ViP6J1o7ROVUUqC9aSOF8CPZVS4MyGM
nYKaLE8jSjQ2hBSyLy2A6ZbOCp+Vwfv9ARMWOsSEIG+bHUmMe9YrNfItTyoJJ4NF
fuxhf5pFgou0gdukPTDcFXOJovDy+gGtH/gwHOjLjytehgwrIkbVFcw1Z3VaO55k
a9BZ/DNAFaf0rLwoytgDxtc/hBDAqwSA/sAVN/W7OtCDbNMsgrlT+gqugwMu9umE
qYXuDhsxGNshQtS9z0Aix03TrwIAsu8di9+3lKedIGVrLA+e+xLXLuY16q8Sd2k8
QnPin+yHWuU4k1f6eHjmZ3wHpVZVFy4wPJXwjouZPCyltmVmzS2rZxYY22Z33fiy
BmBAmQs4LZE9irQhdBNIQEAT6evr52w4cNdvbUukcrHGN9idD0mbZ8B7Kqh3tS/V
RtFNUIC2kVUCNXdeeDue1lJw5un5XTSOdONcO3KG9PzZMTH7IMkelshrhyxLbTxj
7Tvj7xHGWNptsgi8CZaIU+mYel46HuGXLg1B/OoknZ3JthjehXzTcb1Jj/uRZ+Bg
cLM//bwLFmnQyfe2PuDlkh2UxLwdTT3C1tBO9jLmxX3UtKE3j7JI3ZXWbFrfvChS
UhrfY7Fgic1l4eGk1TADKe6vG5zr7upc7r+NrVXt5xaMh+ZmRu/lYD6ziuHAp3cb
+bsB91xizWeFuGzz5bOzbsxUSQcbylex/BTiuhsjoI1wxflPJUG8a8zqzNNRcdgB
1PR7o84LwfdSPH9/ZYpjFRb7d4K+O+HFpCfCP2AWK5zbioqNPw3Yg5FgeT0luHHC
1fIlYJd6jHeDqv37xx8jw7b5DZQwcVsWG7B/OFermtG/bkEC902a6wYkW7gql3Z0
l/dFmx+qZV9Z3lGmmOJjFWOfMK0cuXQnvQLn9jGpWNIgolC7U8LfXK/T1DoiI1kH
/9X1D6wpt8lPYXomMFC5fAMxLo3y7vPJ2ShYP/RTZ/7FCtI9lGQlXX8RZFBbn03f
+C81jgkuRQMFajrvHVDpxOzAmGZeOnb/dZ6O5U7x0VQNJuq+eJMJLQNLV+gQ9s8i
kp8ZNKzlvQyoInoT1Dod+aQDqcapPoenOwDO9dwtZrGRdfNv3xgITzn91sed94y+
d99727hgVZxA0mRIKS7gpAXEFD1F+BaYhJ/rUTMhrsq4k9UlYOS6nimGDqTEzZYK
SNTYCAUtdBozegkp11vp4/fne8beoI4VcH0w9iSzSIZYbHfVSU9z32KXvWsaBFU0
vWtDqqFMusKPgtDGTQ/pBQMXw3xorEq66oGeX03kR+hqvNps0PTzcnpP4GcuEXOe
PqPXgcHXJrYpEY5Gy4zmGJ77nJ9FQbJi/35VEydiL7YO0OM9nBSqEzq+pyHBlSob
T2Hk+ag9Gcqeit1Z5WKdh8Eb3RfWhSXcP6eL5elNe1pl1VpO3lLFGioSxMKD1Yyd
0FCK97QQS3cHoFA3QCxU4HVHqesb3RThqBBk34EN5R1nj8eGtn5QZm7DOrlORqNl
DXXZGpcxzp3Gvq4dh9PS1Ytnppvi2dNJNuA3NmygpbzS8pxzH+upYXnj/mrmtZSl
lqTPtu3qTvWqK0GdUPu4fNDE8r/FcKl0Qp9kcnUurZPO7IwdDxbFrqJf0BWomHOo
A1tZtBmjwx4FIHFo3WWJ7MQ1Z16TzPL9YHCU4+VdG6RmQUG5wo6Hj0IOslgApm1k
Q1h0lsJVuZzrrxztY54R1e0kVYnNmZvE3Q2jCaj7TBJV6vMmRUiGbEw9Aj4TH6B3
sowFgQe3HVZZdJRq+naXb0XBn3NhG38tZUQ6F0C3ia4TT6gsJ27ifeHQmQYJKckK
FSPOyWGFlN1w1En755nU2EWLXcMnZDu/yIXgcJsf9tpDYu2h8Tnx7mQT7kS3q6Tx
B4cxtooSVs7s5QCu3exVHPcJkeoAjcYRenmnIJGHNMVYwqI/YxBhAJJ2ejijU43t
rku/uifuoVqUAZhXvnUNlAS+SNnk7cJxVS3TXnlR4cF5A9QlrLURxu91YaKvXHYV
T/dCmNr42I8LYxdgu7sty9ETaMJb0LY5IczkkHSxFga1tfHo+nW2C/5+oGga/f6I
mP+LRuFkcSIu/FJniPv8CI0JzUZpmQB1nFHsRd3zlx9Bpyq6s3rJrm4Cf1EtxiU4
bZ1navEzSzwQY+GYNUqAnE/rNmLGZr8PKlLB73+8IYPJORKGRJAzE9Ps6G6JNr+f
aiqCGuBrwN0D08KAPKGvaBnK95jEbuU0LZpZ3+G5gQBoOb6l2G/kodnSPsu9vgAI
dl0XsIW16KjIB+MH4VcYDRUnkHufhNZ2KPF4xJslUoaTJjDoOt1/4aQXzLUHdmGU
cK3Y/5qMXWZ7E5QzmdWD3/PSrhD5pcQ4iw0INoh3+ohwsBcwfk8C6BAEOMqrdCOl
0kP2jxzo3u/kxKhIZJgB2ibX3ygbxpUXtlJ69OSgZTMOOWEYsf4KYsNjYu9I9cDr
na7GthM4r3/WCtXwFStjqLqp9VkZPAFWo3KrBn+OZ+hnUo6IKKvp5MeYDYSY+omz
nMwGezw87p7lT3IEVpCu3hMMLrRGd+Cvu3UU1iAxcOCsiJEYULyrZ11w+LiYemHk
yypKBoiOMg/LGOAjOSsCuFEAv+7rSlijMSBbxwM571kT6P8CECQT5brReHmD85SL
MYNZEG45WOHWNTEytvaLxgyRvw8R+/NwIgj0QzIPiGkbahx88doDeifuC6HqTS4V
gwZYi12um0eF5T4F3twh7Oo9HLeKom2hxrS64LrMCLI5bp/cZN4btO8gWip3+2Tu
So351pf7gMq9JbJ5PTauNmdkcgeBWN7pgaex8iDQIpS1Vc41nNjmrr0YJYQVb6qb
4nUqtblqoHTqnbDVHw02bObK+wPJZYQqHz78Agi8JETY/enKLgSyQyl3W0L9SmIK
Lv/RVlp8tV+SF3UO9wPn6mGl4iO6RtV0yBxr13wuyuTnWGmzfdDKAJ5meJqYASni
cFQfopEP8g7b2s+/2RxlL0NF4cESNssTL8CwU7ZIpSCc5LELg2cpqr84iUHlzsCS
2aj0sd4Q/f82YT4niwJSAzi1s+zV3yI90k5vs9TEs6cvxWN302h4gnsnE+4Cks38
k2qogTH2leJEhIYXrLbMgV+MlSTAIdHphqKw6XEpfRE8r8rf3fwnzL5v/29Meo2E
GRAmmkSxVFKpguTqOl2QWiiM6FPxBiDzw20hhT2nTg/ivcK7XqD0VnX0tDsKHJQY
Qtif/8KS4UkmUCxKU+mRyO40mm21wahfJIs+qxQJaQuNub3yNxg7O93IS9boLjwC
2MbTpN/sIX1HTx3KZugbsNZQHkAm7ePJXmBIsWdSSNsjud4cW5qLtE2PKSX7qE5P
g/4ESN2IwvQ23YpoozYWTyb1A5OA8UDf2ocNQNpUpTpi2A8DmFQnTx6ZbNma7cii
Fmo6vfMI/7pVJ1EVQqHx7Jja8LWVZ29sLC2OdTNDh/g7g+2l1H/gBYKKsNd7poXD
FmI5tLxjTb9PD5WM4Jmm7wb3JL3ZApltydOJztEWf8pd7NhVHtkXUyQ5/ImLwNdS
/p/v9icmM4SKJ+8miIfTTu2Pcs9/gm6fpPvePh5Dxjm5hDqwZH/PkbHjh8wV/uq8
pE9zRZCJc11UhJeNnvG2cuG4lbA1ovwhTUI6kXY/RclR0hEP1dEHEHorNRnQqm+x
H5zSWaMB2bcsTvbHJOhCdQxCF/utK31x8pvMgrBYrMB3j6L/F2Of9viw1tBM9gKe
UK1yVk8AtlV0txkl8DIFPV14eAHlXrJG0KPCSXyRoGb721VPxV43cyQ5os/W+KLZ
DLNL48eCwUFS4HH0E4ZvoZWSXfw5N7Ox+CwWPyjVBR0cD9etE6VngDSH9213b4rY
Rkx9f65kep5I/km4Gnxe5u2NfobJFqxilqQyXge/zpBsXIdCSEXCHntCKitCs8wa
e48nFF1Mo2Nq679bk4CS1UKxYiHZfc9YfzYEAuz71xuZknYPHvfuuJA1+UTHvLt0
nCbZiZjxicZHskznXaRhHOQPPpVHcj7/LlL3t6EBiVcVHdc/xRGrRT4wbU4Xc+RF
Gd9DcJZC4DZxH9LLO2sHCa6lLCOxbnPiZn6WNWRYErl1bmOaBx6J40YCCYA6VLZr
LuHVBgEVz080ERinSNt/IdSrIlQEZXJfmhzkRbvSbH/kET0P+3N/fuVltbLl+vhQ
OgwfJumJ+kvjxLUPQfl98y9hXlj1HcB2KTpjMjteei399BRYc14tCg9OrGw8ryhU
QivHZfSN8E6mTQXxobHUhzNN0j7SqehAlnwCXESmcWsEplwcS7E1XKliL+00tSiq
IXho/afno+CzCD3TSOi4ilStG5Q3OR69aTVzWM6O83OWkiUaMHNOTXrJKETKLyXQ
xfHXdhSHkZBshd4ZeR4IoExLhrnSXKx8cdzruW++BbU+HEC6qfY7jiShcfZLgyxu
5oVRLVX7Y4xrgOYuR7H3nKmL8OIkAtLiClHWHx3q0JQGT2Rm850fXkTzHyperSz0
rSkEQiWPQZn63Vby5QWkh/qcHURXWCIQON50I9e335/jd9n9dtQjdgQrxL/CAQ/c
CCYr9Nzp4e/odltYAu3LlK40myWIdzrv73uUpCdMI8LvvxSItm38G7U+LGogRyLu
X2KPrgfZehj8vG8zSdQ8uPeCdi0Zi1h7uXbBnhiWoIqmTZZl4TBuZGzKvr6SVwSc
anXGSSSf257n8XypEsoWY8YSAlw0J1f70AM3WY2lnOyquZtHJmPB0juXN0TCNb5i
WQWwxNfxkJznDzT3xA8ZrOHMAi/D49Ix754/ycHwxxix2fMadYyP3Si+fTzEFFzR
N++9IKhgLQ2A9Xn2YAPdmz1PNfKupxpJDpBQS+DAkxBGpqAdlpCnKEvAtTHHXWBj
moT43XpL3ACaeJxaZryjE6PKVxQazBRaB9ykOMYzRuUgYARhhrc//APzNCxnlzn/
v6tS6RXv7FFLNou+86x+i2uQtSpJcBn4K8hJdQPVvFJ2deeQRDCQ1g0vppftaQZB
eTA21Y6KXI9+7HA+YSc/1R8RXfqt408kifPXVNYOvOaU+clw8K7ytJOpiOOxwoe2
/LyfXFRftw5/044kbeEAajRGEi8P/w8JEGC+3HaYcTTEnOhktcqp+tLCJlWQ21ur
8us2lSiqAkFD+ma4XShHheQpuqbcRQwUTZ23rQOCrYXyMn5EeUbCkgrnB2Yqrnve
0dR9XWZlS239aHlpmY31Ksa1tK4IUukZuV4kcIJ3evD4nvA6qa7uar4QgzaC3Ndm
kEuMLNvYIZOmgrFSosLMxJ+bzrxyblXkVwypTkrxisFJbFyS5lYtZECxdlSVcXcJ
W0OR901qK3rmhlSMJLqUXXELdDFH/bPHXuo2kylL0KrI+ku1HZ0fViQROo02B//I
wV6aVx13XsxEWjvrRyRDN3Pk3QTRjl2ciLgapDVr8whw5GPIespMgFvYJIVzTvKC
87UKR6brL6aLBPc/ivjB+ySrcYTfUtP7MwBxfpmWjUZpEyBhS0VEOT2NoBJTDDVj
BtFO3utrwq1pP1sjV4BMg6TUeddX8jszO8O31Xp278H1QKYNgxy57G6OzauGANbb
lEav93f9XGaDOqiEzBLbLtrUmkWcFiDJiNct52eOxRg1WqlT61y3vaj7nTYZp2cU
BAlcxP1+WPrC3GIaVUxLoI87zT+I4z6rv0LzMHRuBWY=
//pragma protect end_data_block
//pragma protect digest_block
FSJs0xBeAnowLanRDFW92DnsnLk=
//pragma protect end_digest_block
//pragma protect end_protected
