// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
cDTQLUh9xyLm5KZdZVJDypdaqBxLRgxJ9nEKptFqzjPQxI3CC68zs5zRr9RpcOHUOiAKGC0si22C
9pnlaiTAtmn1xNpvbh7mpZ7Vog3zhhijEGOnmifgkXZz/BFvmvlzHcglmyW11CgdT25UFG6jLHkW
zcSBxGyDrGDHRwz76AMFgdms0gWCo5phGqOh65TouH40i0FaYtCqYuYefWQhmPpV3VgmDO8XaD1l
UTOTWALNo8sGt6hSW+/Tf3J4+KNWdEHE5aZZrPYZG3gXVj6SA0EMglZ7CnEnAVYoxRcy5czMB0ZB
8EwwKrqLRrrRE0qbah1yQ5/KccMhSgMS/O3iuw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 8496)
/ckeMXIqkEiMGu26+IH5KPCmob4WMdlnp1lxu/A1CsbwLuhHKiRMhMSiSn80QgG5jxAwId7Odtat
yUNE/j5CeUSsdWy8bWGil9izg0TvD7+9mCvG2PZV8FHstv6E6YGhPohyHtuH10P0UcikYKq8oNWV
HB3xRheH0mOFXdDQYrFuk73EfoQDxZKrKSAVp/dHjwE3PK4mRpFu5bv/mGOpTckHVDnyJ5b6EhJ+
WnVE+lNJKzK6X5ZDBlcdE3cNlznXuM6WDoSGGvDfVkYkcYg7+63WQAd+reX2INcOkgXSlA4dQaex
iGz5USHb9DIuLA3/5+XOh6ucVFEovo7Aw/2cjT5TtX0yFGNcjwCzTrh6HCTM6snsFjETL9HmOr4Q
zT1RhkTC5f0FyhwgDR829jzhyjFmPn2+h/m9c2gG0PImf1eFJvM2sizjUn/WnBvd4IOTJSKA0yYO
CUVdorUaqxOYLM9w0PRO7+I7JBNSejpuBvQdLZP4CowTnTlD7BcMLo/vimReAxcNFSXhADPNJA8p
mBBJ9uVPrt1WbiWc3Kc+V6iGz0w9MHe7aYFgig0D3/w2BCJukbh73CXKmEKanle4OTBrTKuQS/Jn
0ytldVTTIcwQf9usa8YDxMcVninG/maFBU2mDcdcky9hbckV6n136SXuHs0X8O4kqx7Rbt+ri4bj
zFAFYJmOJiF/7lEoqbaBwA7rClSknRvPRy9388/GV10EQ+9f2uJP3fPotkkK3YQ4M3bDPAydXiVi
dQLt/r1D6AMo8KvWQ2yciCXUv6qeqYtJHmyzJQ2FQm3Ke7NWuoHOJOmD7v88+GhtRyvrx3/qHLSm
4y6D+C9qwBu5YMnzVgZ6X0CaZVpay+d9SQ8J1yUyqvd5KKFK6mxqyerdsYPZRuywZafBouRfO5rb
ielf93roxk/BxgitovlOxOz4mPeS/4dzMc8rPJmMR+0YsOE/1hL6fcPkSFjm25HXCaAOPAdwNzjl
30I/RmifytbYgLjnbtJuB8FGgZfm8krdzQDEzvwt2w4YdPprGxq7+bbojd36HI4uPvHlP1kOHZ0S
aoFYiXOkPW3YVT9bKvk+02YlGSVXcM1m5Gl98RmasZBPHaSi+Wft1lnCzvXgyEbkDWQrtOWixTA7
QZ9SGbU1YAQ40qultxSYdjXqqFZ3PIMJ+9gBmV0+g5n0m+mJOJjybuLRovzyCv+zUs8iHATJgWdi
yPFzrWwW/XVxqYKTJMJRNGxkJ3avlDF6LAWIVYCk3PWVFYyiLCxAm2EN5wS82B60UQTHJNGszWjO
8DGta4qisdzGIHsrlvMMOZLn+OVMsF9RUaTd5aumyZtsYWX5HzSWOCXDmQ2AUY6aUhhoS4t9+4fG
zixQobFXRDavb143jN+UMUA15LjibjmcN2s2BFLHEfF1CRwfNxnnbVlUOy9nzUP+HzjKHZ/REzfZ
tEe98kArMQLZqaW95g80ARufgRsayr0YYCb2zHmZ2uLPcLTaut9E38Vff8WUCOvGf8CGgIrfgpUU
eLXwGxeT4bpEw8jljHSThiJaYGJQNdforIFaJ0p+qs+BHHC4Fvlz6O8R/W4vcVO3OsAUb7z7AP8E
rPC4ju8U6NX1pLf0xfVE5dK1cwnHNibSgbNGVGJveFDM7SjTLeO/AEXK5i7ppXs/fvWceyA0OeCy
1i7+Eu3P11ugSnpWudQTMu015n84ckXP93nVl3Y1v82x2PCl1l4hvnCQ8oxiivwnx67pKp9fruXI
SHnzx/dnVLgfVFlXguhJ8xHodSd4c5VnbjgFEuEKUMotr/uQ0JEOEOOuRfP6MHKuZtb49mzfzyC+
p8wXOGfilWxdJu+OQqy3ISRIu8VvQcbRnodzkSIJHKe6XER7oca5HmFkl37HT3tpjeXvp1Yb115J
hilQWmOMevxuojvTPbDsXjmMcfuUgW/TD5gLOiIJHT5wN/DJqX1/xU4/UcUsu3vqJBei5dsVoXmV
oREiBTW3NuyGiqfhZV6Qo0oNaI3Rt3FL5uTLwmIYGPdYPdsFAoc9soajr4+u2zuZKcotj2CwHiBk
d9m9HJLaxPcQ8p5GHj9FWIaPZYkSVyNvL59rcwqdOCDxSg3+bqualgNJT48m58gsIy5xAzfsVa+n
7t9P07ob14VCqt1MRHQX72VntO2ePV0AaGABnnoY+tnoRFoi/azpS0Ld0Kpg8L62QGM6EBxh/KeC
OEsOkVaGm40+tJJ5tFimDNZg31c7JcuXPr2kVtHHIiWCQ94r41wvZgz7b4cbAPi0+xEpFFRBVFUj
C5BJg7Qx5AMr2hDRwd/OCTJJj0WOO8tBXzWvYJZ0Qd+0GTEwRHBOv7hjGm5/gZCXV278zTRrQLua
6gyWKRy8YyaGv/gncLBKydKosM/sxyEEs+xHea7rCU9zUv23r/5EBIDQIM14688HdRv74S9YlyVy
lCLKHBgZJf8b32zPR53wq15eWuDUqJne2356OkObx1WzgMhOun2Gasz/dZkqGGSfYRXWGhFi5FsZ
2P4OfvndaQVeBjrP+K+VPwRyAT7WWOFy5gPCIqm7xVljYTffGPE60ZqAjneWHZ4ZLZoJ67GW5odf
25A+ZY31EbMtY3+wpeMc4k+oFyBgKq0ZFXLZw4UFe34kLdiau9og3MCFPBetZtoD2Z+qse0BmELo
y6M85xGwOtbgnrozwlV+Ke8UjMvy9itVSOVhEf1bF0SvJAVMcGAZoAk2ddfZpB7HsdQjZvgk+QLj
I6REKc/vr/2Fxt8hm3gZvliUzTZZR3Zg3Mgm9qEcHAeo9dAI17WoPk/U8ByhaxoTjj/l4n9Tt9+c
CafHDBURlbKrxnW0/1MqqNA94/n+xojKh97zIisx/9flTkM7eI6Oj6x1ja7gaK8ZQf6upFYYpdU6
M8njz/EWcll9mYPzuGihw+mHBfcU3F0hqkjl8q11brwD8UafKnQW8dooDa8Ff50B7MExfjaQImhd
XUDvtJVBOMLlspgJgwxYCruqKJa9OgcIJC6LQWNeSB068EE/Bl8L0X0U4VykBOe9r5YF/oo3fkdc
oCiescbIuSo71dGUHGEj8PLS3xzBHYT7WyJ1j726lR1cUjvifY/1f0Lb5/VHRmsWpCRzqnakEU9V
fNcJj9EGYQZb0P26s6GxOeNSpWTa8X6NMkMLhogBB9+2kCzPQM387KVxNAcqkn1jPcgU3VlBTGsf
d2kHT7Ccy2u4+T2lVjg8P8rUB69Ar9Z3V3sR1YCNb8Jsn97Q1LEgZzfTFHt2KkDVSBrTUmggRNed
/0OL6edwjcVpr7hD/xKvRbzK2rZTbkkP2Gpm92Ku3eu4cr4t+tUcmsvC8lFt/1RMAmo1lfQQGVke
ITKmaqtqiKAIAByo+09SjMggb5a5b40fdQtvph0oomALJn0xUpGqheTneV+rj3w3wTokFW+0Gw9h
CTqsBOjvULygQgBL2TCbKswMGODPLp/UsHd9GmpT1AAnR/JLTEtfSqTJfgZJhw/K7ZPwB7AJqWs6
3ITlR+I6qXo23LY6VdxSdCZafJ8muRs+LwqKhMkePY1M1QO6LqyCmFdOXxzTr2Olv9EqwxA73BFD
TrsWi23vrOPahYfzxXnl6B6rwzf0hYORE86fL/++PWoD6HlObjEQXDKknpFwlgEcrmU2cw7Co7Fu
yb31L5fEVQgkzyd8aiAkaztD7QWxsP5QPdb6j+tPrB+MfpUnSTFYbdGcOE6/uXyn9BmKkgtodnB6
o6qgEIl0sU0byp6uNvVqBUv31WPOg+ImLdCwrYqvVSea+8dnb2K7J/twKe3g9vXzZSqxty8oi41g
HnQqXtaufTuXCSmwwdnHNyWKbAIyf/ZefcNOIghOtW2B9/COCAo2rk2c92f2BZ90YHnZTFSAOtu1
chPWS00arGDq4KgLr0BYRwJDgzduyzLciDmYPM+do7+6DSFJjcMpU6ll3+mMiilO5rCN5rOVVS79
2QkCOeVwtSSDBM1D5lCugGqZadSKCQcdWFowL+ly5SJlSt5Qek8QnZdPmVgs87omiAq8qPMvx3HT
Ibf6mx9H2VL3j6gQoPEpRb1N+l2ebhBgwc18GgITx0iawn5H12sDh3fXM2sjkwgD6mz98hz/nBqr
Ne8plmBUZ/XkvCLUJq/iCkmAzqFIf0psSci6Vo59HVmQJ3GVZnvtDwSSh/O9BRfS/w3v/E8m3TI2
g+McsE3trEsg1KWP/F1L4HFcJUq2baC82RZDfBGL7QIEyau4drXIWGHtgakh9WqUVC+jUMqfJzAB
gBqZ8uuMk//Cox8dalumkgDUpHZ/gfB6wV6PJtY9ohf3tbZ5+N9Ib8DAzJ1TYGvLEhSV9dsJN8gU
baQph+nH/3TntY9wKSlzGJ+z27NCwRz4syDstVKFVLzOsccWhHE4s+RLk7HMjyjn7vr9xj90vb86
6SZgyGR+excogCqTs9vRxg7/TEsakM0IfngNb1Id4N5tL8G87BD7FOQpL4iwPCezbGCcdxf1a6Eo
L1kM+K0p2Fsf2rsh2qUzCBWbZSg5QufaCPNWOjIkLcCASYA01+9w4ehrFUDa8AcVkHjktPwvjwBn
PSf5AdpbI5ag45g6dOP6LNRw5gI/XsIko/sBAPNbCGQjXw28zpu16p5bAjkuAd3RtwW/peuTKEc1
+4B1P0hu59dhr2V3LrCQPsxDyNxFMsI8X/n+q3sbA0jdO8xy/y0BvvWDpfVtNuNcFUPwzCkLXsf6
zsKgZx/j+nV/FUPT4c0HjD+Qs2vmRbCV4ZayG4OrGbulrYPKFCKajk2qRpnfAeFgez6HO/jLHzQS
P/yRWvsUBtzczlktOcqu4bHgJrKMMY0I5q2AQDDHaYj7hoUtHFWh/L6Kxu0mmSWZuwhmvoFo0enn
imFnNz5yaQUbG6XHX8qdGyX02YwN6cKOy8u679XJndEOTHTVtRk4JAgnAEZVB9/jpHNog41S1xJS
SR5hBXGTXFG/DWJcsqWvdHdA3LP6OUtUnjn4bU/uWgH231TGUPzoa3WX3cMbFlmOKoSMKHtAJUiI
UzLA1OGTOumZA+/zf0SHENZtI2HFITP5mqzA39J/Ke+XkKRhrZDadSaGHcUDBmuOJ8sw3K2eIEb4
MpGCLJbFzO5hpeg9JjQnPrqRIMypebkSIJjyIEfLAlfzLBcd4APNrN6fpRIVAUY+LWUDz+Ml0jDg
7zefFoamcro2Ew0cilT/1AxBPHV0TzqblL6DQr2T5Ct1sSwiSm5l+95HcTGBnOHdRBVT+AIFaQrG
WMhudn8KkynArkpIfQJf/p3CAp6OgkgiNvU/uZnfK6oSD6ycR8CaHY2u1faTzVrevY/DanAQEppn
vLouEEUNMbJRhTOxTbQK75ThWRtQ5/CWBo4ueuBUGK3Xt6Z9sSmOWeFAbCUxKVqbDapcREVty7to
38qGO5WGrAb9+zJ5piFrCN+WnfhrCi1xnOynPY9ln+3ku+oa2nUegxRUtLgXyvz+kgDkPV8mFY5+
n7keISLKcM7rT0xnR5O+xDHPC6I6MZWMLxM64cF7/S2bqBm9AQ1RcIF40vd5ez0ufUFLN9ltykk5
u79knSnZtdqEii/mq+8E8nZztxLUEhEEQvY8pn1keUpbPjvI3a5TkOb7/82356ujMlpOwjbqZeGx
gSvGG+WaSF6SX1bGiIM59AN9a9hCZwa/xUnhG5X+xZg9QGC3SZC8+fqslTJzA5UsfTwt3F46dijc
+MJxhR40rfoBYUaKhfisaJ+HGvMR3rL2VYmZ4cPNPZh2KQaaE5X+pnCEsCvKIUxyBfK4ztcrAFu8
wacaoXpaCoIHV/oaMwiB+QHIaCFDA/9vgr0qFxkwGN1MDFcsXKPYQdPmE8tg155AeXmS+qUU1EF+
oaSoEJ3TH6JqfCzKLuyErEeCPRFvjapkTYgFPDP5PI5EbyIpZL/OCqGrX+VxkBE4tgwE57E50Y8j
ZcwXBF2Tsy5GszuaqOCgw+oG1mF6wgI3sJUCamCM403+YHpxDFfANthBEdEHcotUxXNBK/4Nzpj1
Qt8MJ0DIyp3O1YAFP0d53weljwXprG9HnmvL351G2jTgA8yV54Ul2T5DkY/1dY9zrlC+hmhgLpGY
nN2yAI7ieefiYb6t39Q/FhULKNbj961F2IRvWR6UG49hDpEV2KQGOyq+bzo+2iMKVDqDFQdydL4y
BX3asdz9BopSv9/cEIQNhttHvSZqi1w5hNEamyC+SF9dmYZ+nrLQS1h3+peBBum9bCalTjgraet1
q6ddxeKLAH/9G79ASWuO8ZcNZelp4o6CohCyV33NAeSnWccDw/p0wIlnObXZDNXjK5Is6A5vtQsH
vqGpi1W2U7HS+Jh9Gxvd1nr5vza8F2WJ0IAYo0kYr2aDwXg1eKYTea/zfTO3VPi4+YoVEWveX21z
9PaR+hMzkLj6LZY/KXWZ4UDBiWj74RSLjheJGEv9eoChqTlHMmW+E7lhC39FGqarmvij3w0reBXF
y+RQswlpY34XxeSdshtvEK3M0IM9rRLcONHsgrIQ3sAbPJzp9bber/aqb2pEVI19sZ9hoExjS8f3
8izsiqvFvjNgjc3DlzX+oFljoY/6cPnP632UFys2yb1uxSkKajgrghoY3KpoO5Nv2GVvddWq8JLS
qW9RcXCe9uoE3bKIUz4fJpjZrfteLAG/aut20fVwDxPwGVzU5C2E3n29Q/DdAbqdCCTR7WFXepaj
y6QggTwk+8RnmvHus6Cn1Z6AbWAjQoL1//UU1UHYaHDggYK4ngWoC1uweLu/7+P7BmST/ZMavy50
yMotJp+PT5M5Swhjr9AO7vKykueZ7nfvp40nr+PstQfv2twFP8Dwox17+qJ2dNqMo2c2A7+5nSdl
FWD338Lmaz9tuaiLNHVp4KlcxXuQ+xNkNangbrQgibGgfGn1t9cRuLNQff9i8yKk58A4+UjxiI/1
ikLD6BCubyauhwUxQgktjLJRrv61xb7iq+L9/WvmSAe7OvTuWBy4gedw5Atgqf7zGfqhQf9rkboi
KfvgiGq+3g/BbPBf7LDuyCHnHMXOsWMisfVD/s5UypNAssBTfGoOi2b/6pJNfX6bsjXX5fdboYv3
StBqYnT4W4YWIpAKPbPTOIyRH/EilRWWpdacVhW1v2tSMscQAeO19eqLJHfTBu75DM/TbLKJ/SNO
E/btoK9gfUhEwC9dfYwVKWcZPNob/c3ldjQ1a5HKQaeY+6CRJyLzrfpOf8R/78Da8zelYmCo4LLj
PI74Vx7bf9/BMO5mzkrYsaCc9vW4/cgnRoMvhWtNMIesxGhkFcg/m3WihsmcD0A7hd9c1hBrIKjP
0CfOA7vTFwlGYIseYp9zTh8flA088M3edHupwGOTv7d1r7Usa91q5Id/9JPanF+xIlVG96FWvpRr
NkJ0qjG7RxDEG1I62LKd1mPMIwGfSTeYq6g/4dVY+dEBrVphZv5r6Sd7Jrf+sCM0s1nrTST7u6TF
R3CQDJyw+gmuK7Mb4vjvGF1eCcZoU0GZosPSlb/mVVFzIuNNUB1UVcuJ9ft2G/oPsuRUmMtEKa86
sgPQLolOiZXlsSrPYAuxjgrl5d6WdJJXvC+DsHgDwyYKSzdVVPh8P6cTa36+jJYNkunCa/j+eAE1
KikTEZpNg23cWhJUq7tNyzNPXI4P/vNnJiB9iBZlUmPTgMvUSiBaXKMx165LChcRKkA0NChG0DA8
z06hEgEv18XxwLwMUK1uioIccEJnTSvmiPINKV8ulmvDYQ1nEoZvzNGWVBWqWl/ZXVCFIOIaXS5B
h5xkjzZ8mG8WfHe0lWEcxm4GW4xzPtgeejp0dwczwtVP19W1xm2NcE/Bh7U8NYQHxv8APy5IDfuj
hA1bVNAxMlrFeW2zTcqwSA8rztyO04DwRuWx2B/O6g/vu8JL2A3szbjI79AhftoDYJz7T6Kd2uAl
lrKP9b14PyNEeH9WNAraM+ADXaw9eAf2dwGy7H0AMGRrFqvBOwIkHvQSKmIHwRiV59aqwG7rLV78
XB0rRF+k6QeHTUnFaJNIE1DMiJkYM7xI4h9mRdT51KgJ7dznFo9yirXjFH7rAnCRNZkCoVah5nbB
mXNkVNTaSmfuWtXw0hQswXQLwDqiPcTC/sRDNeiUuT8qfYgqWVjErqwyJQSxrDUFqh1AX7S3qFoH
nnbHBGnVeDI43KQ7qzbWiFB1nLOAmcGJfyi3QS51/5w/PkK4hY7w1AFGUoVSyt4ZO/4LfNNJd8Y5
sKwEPqy9UertnHJkRqax63Csd0eLbNrAgRewN91NlZqpnal9oDrKhbzjC8zDqVuikBxod7Dw2/En
kTppy/XGw43dheMYtyntoDsvX7EAEZrc5sWGi7KP1u1Ic3k7lyVJx33I1+/6iVgwFqo6PmNNVZMG
XWBPAxlano/77/ybQuJ4iNFiX1MKmwDO71R7EMSklFUaR6+ER1MLx1iAQNpNIa1XCeAUK5gRhnxU
2CiwYBBjhccycSbAAkChxZYi5fqPCGo0GOduwpB6XgsM/IgiyNyCVreVb58YWN40Av4sCndqQW27
w/QFN37fd4nf/rzmoCpwZKOjCRXRS38cC5IKNZsZXtSTIgExZo0bY3Qt6t/k1MV3H27M9Ycd254l
tPn/Pp7yO5pJOPUwNdfiXEBxykQfvXYJ3W3Hbjn0HfhmFJbIjLMlJH8Uct4Jp96eOLRQbd6DF4sT
hMmOMQUbFGALtOdc+XZRzN7xXep9BRVQsk2O1I46dFziLQfQF94NtG8dyDXcq5mV0MKvVH4Gl/3x
IUtnzbl1bOog6Zhr8jiS9LWf+SMSJDUkzj2SaWkB+2kkzKyiD/UK4XKwillQxRpRDOuApTXj4DN8
mjSE1JkGzeunQoC2nWt/SPkEpBg5dNytrEianc6CyP4+A9n2+8n3ddNOxiJdbxebGMSx7o/zsP5d
ScBWSu6rqXcjQRWGmpW8WA0WaiNGiG+U8+J3HBDxMdkbOy89zHZlUQ0yav+GDvVd//dUAgy/boXt
1iKQRLLA3R66lvgAr+4Kho6BipwXEEXR9yTnzi2Hkv+tWbinpWIFWHyvsBvvwuLlMQeA/2JQrakO
l3c/qVqwoBNhtXuL/Ibh11cH2/zmqEBLcIzFi3iMQgwBOJVwlj+MdQD3d6RfHa7f82iFGKDDdhpb
7FIinDrwklhWCVX3V9xzQOt7972/HYbZ0pmNODnOalWQP7XmIljheOP0JFwb1faE1bL5g2FTQaR/
MrOwu2qQJK23gMs65Mj2qR+uUEi9RsxkH0ui9NF3QUJZhxVBPYbPONaO8dMVreQg8rxj+C31nIf7
fPFY4N+fMpt4I1kI/qcHji3eriTSGyNd1RKaBVZg/m12w7NLIg6zB62nR+XMaH4zPZuCxoCTi/l9
dAYMmYSwFOiWBHzV7sxS5bzH4TUraXEyjg5xmfW69JNEkDnKHyQJgcxwIeCKKuW2Cxecze+ccouN
VTZLe5vrhfgDogxrw3iVNTIEyLgdNbzlUr58MpttJNOxeM5E5RVRqrnhNSr66Bw76PNNeM7tw9uj
a0bjWzqpYw4+Nei2Qzgqc69F7XPnfGtcHMMA0g3vXQg7YNd2ydi3OiI7QU7gPJwj4pcGpYQ/OmKF
CA6vNUDB0N1/wbWNlbQH+OKGS3A0Vg3ijFgyM9vIdqe34Gs//IY840oilixTf2ujUubx9T0uBx8g
ddG2usZ9mdSVNm0h7sKr8toY3nNNVhRyc/h/LQmeckRIWFMCUkspobN+1gzUUqyOKyCKrgrP7zjc
yj1/gvpFnRDtPNWbP6ckbG3Dzm7RYL/gQ8ydyvRr71S7t380DqIrhnXJUbBb6WG/CUpI8gDXHF31
jiinedIc0GN7uVE2qoinvze2b60SbRWlhNbqxYACYRAm1wIuov9rxnr/TNURBh0suj7pxv4uNkwC
vxHPhQEC0TB5IJW0hi3LKFYAqrcsgNXYXDkk1Q79ok0LK7JLTUGwSC/QDha5PGZHqC3asz24m5zi
//IT+OC7KEd2fhAnqAMvHknXDl5TveJJHzJ1InpPbCDjHfEo8PfK7XKwgoJA3tVtDF+W21oYt9H1
QBYuPsPgLf7vabszo4B7+QpK3woSXcfQJiKObVHDuuIIz1SlSSclZbz4l1YQIhrZzpECi0kDS2s3
MBngS2QdKcx50345BsaGYnlxlbbXIFPlY6JDWco/bbxluCXfzLPiJDARbgHVEC1apM+RO6p5symL
M+nuHhchKxC6ntSExvGB1q2WrAYWwMwpDfhKH+k8dfEIKaPmp8dVlrf0S4iUisvJnfAxgfG0jj5L
ZOcZLdOjybfQxADe8KE1X5tne61LJyGsVFaQCBpX6uBNbqcfXabquA1TC9jjIT6lgzjZhpzn7xkH
KxWZpFDJgsfAYUzh7H7wYPY4MoSruuLqGYHvnzqhkdc84DkVzj/AysnJS7jpFMDFJP/H5HxmDZnz
yUpmyImVGKSU6yF+aMiXpvGgmg9pNwphMenwRGOLYOvUwrzpGE2Nf0XEcFmTV3/SlctSIX/UGSd4
aURG8DM1L6+702QHGmIZd6pjIggs7OoO8HdxuQegvLPg862iFi9HOnymOlevmJNccdUQ51IUg69O
BO9H8sNoPi0fNZ5nOn9VSJ7/7FNc4Ib9XyizRId+f701z/qiKVymyDeNBA+WpNC+BtNtvPU4XYb9
n5fKoIgOjny3dDDW5jkmmU8y9TAwgpxvt36mylaVN/OjbJp88nS/EdSVXqWIAH7Ws5F00oJCQ1sB
+SsFbqBATk84zLeSOPvd2BMXiKz55A/A0s/13OQFwYb4TFH5tZAi6yte8F4zwKoAIz3NTTMZNjml
ZupXvbTdotMbnBp8nkr6SBAXZCxnn1FvyYSt15OZxbfXR9wyWCjw7inRigSmDIerJSc3SYkxCaOI
HmP9M912/Xt8nXK/qVjAWzcujooUKY/t5iaYnjpAJDQTHBeipnnk6pV81+CbAGuc128OsZPzEk6g
hztJ3R+ynBEFS6fivT/CxesSybAoCl+6wp00pcV0bi3rKD3clHkM0HZ2gyfKbDnG2T3tVCobHh3O
cAB6EbHSgMXZGZAI4Uf0aOM7F1WbZaC3PKH7delehVjZo9zBn0wzubrQVF/kSgEgCj3ul95HuM3g
jWClUJ/o/h5TufboMmGqYzaIRayBX+8BYIVfZaOaMODE51O4qlm7K5gzGcftQ+Lc4QPcdb40gz+L
LenBt3tnoA6A/DqEB3lmCfh6IvJr3CF7EDpIACNSspT/d9L7TrFWrIQhLVGWQQeBzG2mw0xAgLn1
WoPUR0S0peYWZ85wBn2Hnabrou9bMzcFumoZiKAF4sGqBlMw4XD0ZuMxXZuJR4yB1o0bwVRjHzIb
DDvM
`pragma protect end_protected
