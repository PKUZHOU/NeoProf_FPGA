// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
L3DMCkWskHnBX2Kov/bLeANpkySs93wRCbzZG0OEiCdi/BZbpwm7HISG/D143iR7
m98axVjEJobw/mJ4HHvaHxGBCnG7QIS2fWnm8NTe1Lecg6WxqW0KSmLfMX4UfMaX
Bi9jJpVrrXLf3fMpUKKxGxuCs7qqVkVBu2RI8TgAFRvOcKPS1Og5dg==
//pragma protect end_key_block
//pragma protect digest_block
rOir2tNS6n9FzlztmAIs1D/1DNQ=
//pragma protect end_digest_block
//pragma protect data_block
qm/o+X+J+jwh/yjVWCk7Yf6lOQQxHDMy/I9FaDAIBV5XLuf460MTvTB7K/g3GQLx
VHxuaPadsWBarS8QGGVTKDfCVN7TDXfbmrAfRoVrYyDgerN9b9dXNFyBmbSJKk4X
Vi20ouopXWgRwU9nsPec576KBKZGqDPNJL0qdjSWqhj783gka4RIIWtSEH47xSOF
9Y/8ZN5fFwXSUYdX1k6l3CzymOJhnh2w6CkvR+n2gywFu7WOuUm2SkyEiRGCUKEB
4OZxthAKmpHOU0pF/53LhY5vpZ+466/sOYBAZHo4ik/Gs3ZdXC7LsR8xeG56BDNc
IOJMaB/QU/5lTjVpIUp+dearan/DdL16L7rUhl6NbH6HpDDl8szIEL7kqGzc6BCF
Hh3GYTBRun2gBszfWQLKhlFJKP7uH7myOAJqkz0vpCoQ+Gr3CoQylMaOqniSybpp
xAYh6tmVYxuseT/c2ODQcZeiUIMc+SSx2+gH0UXxdOkcfUBrpXk6hO03J/1HDXFW
CM3rtYPzdimc2kJ6FrOBeKlIrVzMcTq+2qeyAq0ZFo+WaSjnMW1t2GEHmBXQpMIJ
EMYb69ptP4YmsA9sIGZf03pcq1Pdo9Q0jWVEiiDQtCTh7p7ANr323JyAC9eNY0q9
WxD4mUExL1dUJ7TZzu3hpl57O8n943a58lNZe7LQYRkV9pCXSq1fX37bNPzBn16Z
vTmXMg9dE0anIBn9YAFbIHXoGaNhQwLeYPTtkFtquYNPrtxZQnYl6UdyRmLbaPIq
ANNNLEfwFzEHtYDEOsHgkOSwFvBG1IL1N0q7VulbjaeA0aOJ9aIqHNLtVabsVyx8
4t7RhzmWbSTwofIr7syAtdtsw4fFq77notYaCXY6eh9+UfNEI4fAHtfXDhFTIF0b
pKMBJX5qtiK9v4BGKSBoa0A0ohOg8KK5ij5NZgJgAauMM7c1kZim+Zv1/cI9Odzh
9wLl7PsXTCnYTQD4Sz/7SGk3z1y1VnC2UNdH36lozKI2j8PBo3f6IV8q27NnoZch
AbmgPXfLorINn4W4uKkmGGa1YavwjpAa9izvTXni1CJjjuto1C6/ozJE6940S4vO
xq3X2fCWa+caGnxkGkza9qE5OJ7hx1vvkyDphGFQ3icGOtc0M8Z35nMfgyNIhh2b
zddiW5F6tYAIW8l+Pl+amMt3cVOFb4+zdZbo0c9i+dVmWRrcy62GQggCCoNzsGa8
WWnXzScGzgpdSQqOiewUuVfeL5cbgzmVq5fVogdIqnFMGbpoTeid4hG6sMif6JkK
aKKXPwWQo9EUMkKx4GngAtLhyoSvpy2050O9QieahQfzU+K07bofemTXhMcx7Gpw
e1bwDy/GoASvMQHL9BqyvF5ig2o60+WqM0Tcvc2TaQ8seiyjjgOKKTcCY13o6v0O
5ME2WNtuho8YCrnMHspQ8zUslApz9kJTO19qYBiqIUNDZ4uqjLllmovN8WGfdolp
FpTDcNTXrdi2+EJU4e1ww2y0go6lxi+dT60YWaY+P5RNq3poCjmq3hBWbu5zO8Im
07cwbMMQg1qaq7eHaMeTxc2YT4HMQEWMfSnPmqfrgoVRq49rFj2fwuZdamhnj+Hm
g5g1+hXcVrUDOXZvY3HG8cW211mvDzB+4q8InPE4HN1dvKMwNtLir2UwQk0mnFXl
+fILrf7F3zESAgoJCMZVjrUDpxaZEbL94RC1rXVdqUDdIRj/I5iFvxPO8AGfvLdT
HhC9yY5bSxOXVaLadVi8X4j+rgZsd7ciFtfsgtw4+0uoL0W6IuMLjcWYRoIAUXv8
QRJcxHk7RTDmY63hzMKXrya4GQT2qS82GuT3YB84S7WPwIJbhUS6fzr0Yy734Mdd
G/TJDgi3PbR4ArgLBRaBd+MR53ulVW7iKopme2d713rUldw35WyTED+xD058KOEF
qLNMTUL0z70APF/IHLezdTXU6JFmHGZ9O3IKn6B5jy5m0n9f9WvI0DsGT4yTULjs
dIfTqTf6CjwpKfSqZG/lKTMJO9FNtocBad7FoZe/LxkBq/WDHOQbnGh4U7tYvT7t
cmzE5cu7rTsbx55gI715ChHzt7WthIRkQEEsdLRYyGg/+EuyePJS1SuRlOMMEf4Y
dPp44bQubNabJyg3z0WZNmscmLJxPSK+jypdJ5vYNxHdFPwbuNI6jRvwuwlnDMsM
pNdhLfbxPOdc/OrYhsJNHaiZetWilWZqD6LMTx6eKDhRGpFrIe8Owtl9h9n6NY1i
CXnaYG2x6gp39d7P8gVLpsQ8D910CMKgsN0B+hypCpzgY09j9S6UJLL0xrQXLErC
QQ1Ds6LYM9kpVZcltJnVKALJGVdCBSflSoJPG9AuDsmS4ndOcFCZze53pQxYR8Mz
1cXfjfSO8TmK8XVjtQocuOAElcqmknxfrwv3TRDRBNbc296TNZ5qto66oOTeZ8d+
zy9LucMSyFYQZaJeGHXZ3/xkThgetx0qp4xjcagUksEoMXfgaB9kiKspq6+QQbvP
vEaodH8KjtFRABYSun0ZeId4+WUjuzFey3gENvvXHlU+yk0yaxImQp/ekFPEBfat
uRxUqsCkCr1Qr6iKqzHtCMmTTtv/ZyUeDKuDW1pJbnBOuLzYi05ZgZ+aEZtbUKyN
AhqiMWk8MfVpprl2D/+L1lb36O0s1EdDblMrpOyElens0r3wZOdt6Jah/TWze7qm
T7mQOEFD+rJ1rRur3CqlE/qz47UjcpmAKLmEEgPitAL92pSiRKhyuJcTnfvJWqhx
Yok9ju3VS1DwQ9DzNXPFr0BAfaIXbp1vCaiZYs2ncaUKJ5FXpmK1/0DyBzl02DT6
lGdieCa2YtbLMsygZzajw/csVuWW6dCMiG0tCXdaPpvmevI82bSlflUIVWfxfjQX
fIgChGA5ySNXqCJgQCN8kMfWM/dzoRF8CUcqW5YURvkuFVlfI3e5VsLNEMXMOyCo
E8hx/4K5XoDh/sFfc4vP2I0B9gosv7Zae9IN4ica9VTvfGiG1cOSzDnRK0ENhiHp
zHl/ha5iINXMIg9m73ltQ2um7WRysiSXnKFGBI8qLLysgddeITzFgk3Km9+3TIAr
30EK/zcYO+rzzL6f781cocn+4vVm03Eiq330oljjImonPDS7mEG8U5W8pwVA8Xza
AZcy4sbbl+vNR0wOsHraxZYNTLrmQ91syXpCQEy4u2mITarGrkeY6YSn3PFuFOgR
h6uaF/AD6MiK4X4T4ajIiOuIPMClq+9gEYKyVpEUtGuZIAeMvG+Xisi2fkCo9MKH
LGVJkONnujIG/lOWXhcaEU85mf9xyhi4k16Kh2Jd0fxLAsBZoJgGHjV18E3Ausjo
ogo5Qpv7GO+6PYUFD7w89AqHGs/1IqEvRIorskqhF5N13AJ//aQRxIVJ1DWXYgPQ
l5YGRQNeXABUW10rzdj4IcWPLt+1Puw0dyumVYLFPNYkC7Ep6ui+L5DZj2m3X5tE
J59cOHwhBEVy0eDK/Hhxi0jAiPeabJceJ6jIdXLAhpnhsCJQi3ie5YGf1JuvSU+n
shORVjioGlNUxwtj/GLe6QirmqinNOyRp4jTOBwRFOpINj8Df5s5R0pINOQr3cMS
s5ZvhuTB5c1v06uzdjv9vy75pT18D64Wt7PTnjMAW7fn7pzbTpwLDyLbbOpHq8Dq
2rgV+hQEU0HxaxOKHFgzqNnWEVqExRR6wNjHg8jtipHq4ALgVmoCtMZ10Bj0Ax0V
jnwFzq0Xw3Wr9DkLjcieK4vUhV67SnzPIWmivPLLa/6NesWqDxUHGb0S7vbWZedD
WlvVy9SPNs8uEUXIGApEFzqS/4OS4P0q/ogObRZIGq+CkW5eQvbDy8ZXvnvQXN/0
dWVGt4ArNDeLo9buoNXdHo7avEkFt+daGM4slfq6mSFtB+2Z4ASnJoVU5zvOvGIE
5cbVXh3GGildG5KgUMbVAI62/3vmry//ELsTlm2QsxxzHARvAOVo+EsEOmrOvVP0
MrU75lJQxh1+yYwCblqy7tgll+HMMRcNwjv5S55l/cIs7Eko8drKsuvlO7SJRJca
ZfgpTSuJ0VHigHQHPwFiiHtMKT7TpUb9+60akLiMxW8UdGiyglrRzVKPBRCFccY4
zR9G7wzbogz2C0S+fM26lc2bemsUqmvg0BYWnZke3VQvA4cxIXwLZt/akICyniIx
edyifE57XnlmQwYlDUanwaars5VVD2KOyNzzVthNmlA3ajqU6A7iLB2ztjVxV9lS
LOWA6RUQfFHhZq4QHHOV5+b+OAzfoVlVnZ7jGw+E5aHQE7k29b5jRgg9usRNrlCo
wa6aIdqn+CPjYfQMng32K1FGHC7pKoQ8PyT8Pw47lyp4aLsQgcAvWxP0R4yI9tb6
bURN2OKPsTq8rKkxCz0op6k3RT1EPVTw94XLy/4Gk2tioUpbKjHOYJudPTMRdul0
xd3QeElRNoxPEqVsA99pE9W5/4qioc3yLeUgsYgFSGjmSReIVtSq2ErklYZqI+aq
JFiwlAl3I/XQkFB/aNa34bLZIpz2lAcV2hj19edvERA5FDBcf2vQdzUIgnueCO86
A2ThXrLxibCJOQ6k4e54axX1jR2a/h3aRJEaRudaAjImQoV4276QXIbP0PKesB9z
151LxShWRGhYCXgCQp+UamANYbU8+yCU2FqF3efyYUQZhWVbUBmFhskrh46qYdzZ
Nr6Hsw+xkgYN3PZs2F3tRSXn6NQaaAac/g9YtfeQzR1vymQQ85pP5ttWvRbf6OAb
kvwu9gBUyyrXPzV0gNTPODanqNdyBuEy13Jm7alqUSZUPTt5Sy6Svd2PeP1eqVuS
5kZV1G6yhFAu86f3dS65dsmVj+6JhkOxDqGrocI2Kpuswj42pyxTd93463rYmDOQ
Zqa/3Fcw4GV/jKL2ml13ULYcdBqN8n39EGlGk727g+NbtLI0t5DhGOrt4TTQBB5D
3Z+tweJjQLPbvk+shMkeUiLare415Mz7l5RNKM5aCUrNiSREy4KyuXwcf4CN5aZD
P4fuQ/e655AkiRl8qEni2CZKqWVZ9qXA5qgUVElI5E8aAg51n9Z3luqPySDdqQ+c
Vdcg/uvRQhOSfVGwahiiU7l5iUVZccEdzaEzrbrnQOOzNt0d05zYlaaCX4oGgczP
EUE7KZQ9IhIwL41kjdIQgsAYc9Aeboa3phNNf4JPYj7+WtlgucWvQyALwV+ffp7K
S6kOT1+GSb9T+dZw/hhh2OUJ6HeR4+1NXT0s9olkM50aIQyq2+9n02BU/HAn/TuP
Yj5MKMMAM9jDjpNDTpGPEwfZ0183bkWkMlNqB/ht8+xNo0D+5EuBkjoVuHqPpCyS
5ueN0KqOMKnOk8td3AEtFKlP56+m2Xucpn5J5lo8S5XoPieJNUcHwqxJhqJTtN5V
2u/XZUQzBx7P4ixA3VS6/Ji9Q8GBuJTGUpH+1uS+mfGFjNnG+YaF+LcjfmhuWS+7
ro3cAzFPRRxF1eJJOhaoc1GVV/hYgZWb4Oa5GrRHLOuZpcSIi8SHzHidAKZFRJga
EGx81Un7/iBhxH2OiSQoxtvDqNxsHCKDZ5dhxQN0ovCtnkyjX+xdMuRG4GnNGajZ
rwqAxToWOizovwO7DpkXyYxY0/vGntjFpcfQnBmociOlw2PRz0jiRZ0QxrRo629y
JMm7R95IUXP+AXuT4Cg+VPZSagDMEOVEfwxIJ6x71TE4DeNU5obewFrakshn+b6Q
9scOLsVC4oNzfj7WeFXX+X0aZMp9GNUyMjTqsZr9q3y9mySTOL2IhRVP5EoVtWL8
vmVMdlgdt0qQUsbepJtuvLBgtG7rBzxMioM8nhitQsLOrnrNK4c/QoHgZNofZ7wx
Z/AiZxOTWGovUWkBpYO9ixboucDrWVq92BMjcyLNb51ZGxsOuxKLjW7H15MxRoGz
8rRVXy1NynEu0KjK3VLHHkr5/YkUE1Iaw6FBXLpFIkXBKDyPBZmlykiHa5YCMl5H
Ms6WCZbTv0tgIrNTs9+5AkeXlKeI20wdXMNGyrjhAiNfT3+qLdXWlC1LnWXR4X0/
ZKeiOybKu0tuNtQCKyhM2BDdpL/Nk4P151Bs+bBbI5RpC0mquGaonc0MaQMoDG8f
kiJGL2L91KciFnKyj2FWlx8+puvw9+dvTf9xdrTc+otqF34XZUjftVhqdK/hLMBL
X665XxqMv2pNOaxy5O9qreA9kbp7SvxcUJUeINb5chslGnpsY7M5BtSR1zBp1Cqz
I9P46gdQogKIr7kXKAUr/W813UgJJQ6eJvQ8238qr3YdRcRecbys2W7r9W13S0UQ
XXtwb2gR2+I2sfZcSxvZJ64GSQf34d6NYDS+QxaHi+JOTBvPaki9wbEz5ewSEBoN
ewsMnm+lfiQ6qmgAdfJAo9d/M7+/toPLAsxxn1PzX9mhfwigvR+UJdLXRJm84a/p
8pBlF8O8nE+t/4CCuoHc8yhOvuLelAuILrjESWbiBgGLgZ3pO+RXglm9zGPtGkEG
hwwnmjd+gbREpVdB8mFhEV2g451mQvl1fEXzayObg0a4mSboVMMInKeZOULBlcTo
BweSrDWslKgbPfp6sHgUQ9K2HuvFj8kMt7xa3j7ZHW5HlYM6fisrDFu6TQqacUVT
PLvJDg7SKbP+pUsDZSD96TH6Fyk0W1u5qjcVGIHFO6T8KiWwg8pUcee2dQV3fVJ7
kVH4xpypwyaDFukalDp5LlRQ/4Rp+4JToExzh+gSIyiEoBzv8dGeFEW/Z7WAZJu/
n0qf3Gs6BewIeDpv/SynYhRwwy3qOU9vdZQgJSvA0QAG8mNadpF1pkyA9y4QRTTT
2PjV3zZJRKLbZwTgHQ6mX4PMnC5gEwt3U4bTMJch7dk4cJapqIfFGHA4NrBXrt0e
PBQQ66sEnSyNkModGEKdp7i22kqv0wpQ73ikSObW2JLC2U5l7eegRBggy7DBXST7
iGN9YbqcEFbO465n3qMGHBsf+UqvinR/WdmEM8HyYjjoTmnmCsXl2NID7S8jLaB4
YTcqOF6cVbNQ4oYQfgWGX6aiiKp+31hm3dHZjRUpqkmr25AuMhXnFr70E3ojuqfb
6mzRjyHnBS7p5yntZSdB7wyzMaMFT3TxHq/hDz4nY1yyv4piJfEZTpC0pucgnZBi
bjrDc2fNBeFb/m6ahgwBBY9sdHfbd3c4/QMLb7VzPQspKN0C/1ErYaCMJQ1vDm44
BQJIZQpYJWMu11XOuO1ZqffvWnnz4SyvibtGQJ286R+GDTzz7Ks/XPuV/etnm+r7
fB455fss4z5uqyL45vPkbApC78v6i0zrmehEv9GTrvj3M3qQSewoPyr/974cpmvq
tMtD6IODq9fkQqKWEw/8STTCMDkFQItnz3LAKAySYofjvm8Y8kU6bOVZB8lX9P3h
y1YcTkiXnJFIxFMeaqJb+6hfKr+s40nbkprSKj1RqY+knzAvo3IVi/TiOCEvCgze
tPXfJB/tADg80n1ZsSW+swAQEULUdCagw1Ind4sB5ybe6PeLmGlLV4pBNTsYKLb6
8fs65/ghX32JniuSvI8P7MV7UN7slpu4B4ypTE40Kvtpn1efj5G4FVAmopEhZd3K
BgNvIuC2ZM3cyAHHCUspc3rgnOORJYN9cP8uwm3usoaPyneIB5zOjN8HY005bY7r
D0HWDvqpu86dXmVWQzVFG08z4iryhftZkFfwTGNnEj+kcckPAM6LcI6a+ST5HfkS
tPAqiRDgE/jm4CUCWLZhU6rRHneTF0tNjovWTchJy+sDWvfsTHM6RoAuaUeyxUgY
7LmsTJ+jwo0VzmKWD7E4J3AcbL8tDeMPRcVVuJWW0uO9TuPwCDgjGsVRG3k08SOi
7Ej/yEXDdFSekYphrNnpBCTACBXdIcw2PJTbazP9XkYLE3oQoPjqGoJ95lo/c3h5
gvIkKNJNtR3q15FA/31pccHyjeKXMRlrbkAdORAKYBpaqrRxyFdS4pNnbQyEy5Mi
zC31OflbH2+yOrnVjZ2RLubYjoPWlyBJ0owT7KTuO3AJCTB/0qSEFkYaj8z1KkB/
ERJ08fNjb4/mDxKIYoRZP4tu7X+zlrd7r+Bds5v28QCnbLUXBCcce5L1qYC6p2RV
QRRWnjeuP9uhUAy2P58QAZgvBY7cRuLv1KVca20ZZk43CdGfoDxCthZfWUfEanXF
Tlnij++xXhShjpvXYgTXlsjH2Js19bVSC4fE7TOzWDoWH4/uzAGmRGSv+4h6iIln
+rxmOoatjxQWo9QWXxYhhFb+pTmAbcgvNGLMGGuaAL7VAVlbcqABeUGWLi6QmXgg
o2T9iOHO2C85aqOXD/K0g6XUr0tT1p3snMKtkzAzG7MTohUxKEXq8F0oFUYm8QaS
6oltJUT3mjSQmjG02cKsfFDLQ2ENZy6Q9POVc0QbDZrowhCL3bu1s03Y34TUm/Fy
DMMcyZ3tm6SSAuRpax/5U7riXlhALEMjrGPjkvUx8b7ZiOyGn0LVjTxt/oSWMyZL
UGD6A42TCPXiT7o0h87RB110pbUQT/HIpmzal+DlpRkkB3nfNbjLLW8hQKbSfnM5
GqZ+N4kJWZuu87NL22l8Hc8Ka9b984hEyQsqfzLqJtJ7ojagBj7vhVo76rkO5wwF
LTeu3cBm/dRd7hrVzxS55F1uuvNvVwEE7IRTw+IEPTTyeq1mBt63sPXfj4xGvY4f
8C8nuSQVMWEp/lz4K03JQjTOrARWs/6Uf6DDGnL4wTWNkbQmoslWugeGus4477W4
DI1qKR2nA8PEWx39vT5VjFkb9ZUZVjERTNu66omCHlrvDyfnGch38856v46/vRD0
hsVTs+Vz/DrxU03h2eUHmJ1B6bfRURhEZCewXTs31RShXaRnQrCFn1eY5XjFksbR
gwZqyMbnFspCicy7e5MfquZm93MwSZ5m1lFWEV+SpF3Y+blxsHIEdAIug18on7RZ
3aIUt51OPhnL29JgoGmxtDSnj7xybCeSWs3jIjYchW19op0mpPlQOT1UBPr7otAj
/1VPwgEpFEzv3cAQPbfe7FNPk71Y6wFSvi/Tx3Zmz6fZUPTN+3avvsKehZ81YpJR
xQVWiMdlS9KPCbxend3m587ZLJIjSnJlUo9OeYgMXPb0nKd2RdXkMPcxuCf4SJ45
wCvi9hniD2MdI8GAjBwEGJnorAteqO42CC4BV4V5UToB8rmAgBcY6lRRDWn3vEzE
jOUHdfI1rIo2bz4wxKF7yiKfkKp90az+BPaDI8HBr6kPvRcutUZ4eJJZaVn0Y52y
MEgBomcgINNF8eRjUUWZKAXs0ctsZzeBahfFzte2AdaEuTgc8JWK96KFVsyarKyR
xEA1HJQzRHl8YIJ2Fm7lbuqnNwuXS14i1nM/zLQaCrcfNGJuUGXUnBfe7IHflWWG
A37s/wMAU3zygAX4QYotzWDKIPM0CDFD7vO0c50yplUjhYZcC7QIC4bELz1XUzNH
kptCfRz/zpCYAkF9scRMlKHR5xMp+nq42/8yLiBZOHZLWE+xqP/hi9LccT8P1wRP
B3rTWL63OaXZuwYjg/g5lswmwUUh2kfkO6/kdC3w3ll6kBJNDXrzIhaQV0eX4fFV
SA8L9Ury0JrEL/unMr498pMZQ1ygxBlLJ4gZ4lXJP1RXk094HDBHb6kc4IiwAf/G
/NhIqa7xCHOE0ljmY8QSJk4gB1YE2uvE+nQRP13URHxv0H1KPG4fhBz4yFaAjY1h
fMFeIUURaWi97HgbfGff6P9/ZJMUSEZlBf6hyRzEDFwMi52xWMj5yPXJsu5JKBvi
9gRh5OSMQt9/MxG5numoeepzmEXRNaUnzBEyF+qIGF39qnjMDS4hmeInQWLmz8ss
nQbrlNqIm+xGxoe2hwtyJF7daGLFq40g+xWque/zJu7WLRDJqW+7z/Q5S2KwS9We
iPtH1uMaDJ+c5jvV1iy2T/zoSUEa1Br8ArgdNF/AeL9zcxZjOb5WxNOaUfumQl39
+ETHtRBpLskSHDlrTJ3IxW6qyZWJ1aPyUWnvMKLjGFEpvVux3tans9U8vg7HxD6K
adG0cQAWG2MoyIOeXhTE3C1xjMNlqUeawUMm2Upg0Grf2i791Hjc6jzGLPf9V+gD
629mopPQQl6QvuWYKyqVfnlRfrMvqJ9ckFN9jK4MmB4xEbGcuMnL9mb6417cIAKW
Z79rpopheu6Bw2B8Uf+V3qxCYCL1kTXg9FDnfQrptloeLDYAOV4Y0XvOnBiQYSc7
zJE6vH/IBpgjOQV0NM/rdzK64C+sTu6QYMlWA2POry2a2RMq75xqObPZXQIVKCFb
TUih2uews30GZCpr6Lwx4zUT8FRr2RcLYIW4xS1YbR4tPNR11Qn/IwkWdNTCgx21
UNkO5m3x3le8Do00aoyvuGrypvp34lwzW5aaAbttqsYXXmzaSM8xzGJUIDFeWoua
CVytE1OivCu4pVgYwQeK+9WpW770FKUSs8BaCrycXFooQGlAMpWxtpON+xr7xoHH
chfo5va7tP/FMmhqrv5WGdxhsaxfGWFSAfcUVxy99cY4G6Ge21rKhm4fA/8EWdN/
vSor496/Lz26CsCPcA4FzN/O3vk6sh0k0rS3oPQBKBEyO/MDCCeGEW+0qcvDt8d6
m1iipKAjEOAVGiM/oztiR8t2GL3SHv4W+uF7JJARzFoVuQx9p8y4KJltHPWt3g89
xjrjvJ6fwlWjDebdWiNNT3BKF7Xoi++0P4YfSL7wqBUdOqv5gFgQihWNAqPlq22+
RwaQyb/Lkga+x68xXUxnBwK9Z1vOKGII2hf9mfWnd+9J1jACrtB/ulDnfiKX0YBx
YjyrZiB+XW15KF5K7OzPUAsQqF78VGP5zal/UxvWsCQfbnEwUYhfmG/KAFC2MfMN
UiJH1a2dI3O8jGJVitvUk28cPhr/Fv8TY4NFvpCnIhuW+mQi5m/qOH+hH6FHwfyE
4BZo1XI0CD/q+e5LMWKmMn0KmzyzK8mTrjDhRVfCnIezvhc5ja3uaM4sS6U5S9QQ
P4aNdptQ7UudeXbdQmhkQGBSLwzdh2Qtqm4W5oWanWkgR1cDG8gk9/RMXM115nQ2
IqZxtaNCW1RktdQIBeeVlvg8MnIHauH3xfi7i1gODY+RbfcwRjAhijsS42JApS2B
+4aqGzX6jVap6F11au9RkFKquS3tWAuuoXT/NQ2uODAnuYhMLmkeS+xDNdVGFZSH
deiZibPRWThR/MyhaGHPmRTifZC5kK0sbJHkj3s1LH1V38kFaXFjrOut2s/nhT1k
5rOBZ3+7KZJQS62QhJTcr/8/HJmGsx3IerxL4y9ohk+p2rgkjsx4OcYEU/AQMBMC
xSYS/OJRsrdMQLuJy0YZRIy5PrcjJ+M+nTlmH8CEilkGCNOjRXch+EsG7RjdN8to
z4E6qo2XmAg9NByip81J/qWApYanTk/OkmTOQqhX/PHSXNNlweNR294bpXzR4QqH
MMHYr/2Wc5GAUiJ3XpH7ZJqZdD1+Nw/qB0RSfkIf6d3GIN2boQKzrKknt7rZQs1v
FWWbeO8r+9pKxbXez/YFDnFk92t7BnUAfH18VNeDQNoCsg2u6nyByJcQdIqbI/Ye
x1ugInk8ZopBklI1WjnlzsnPPEXgxevB9685G00uysZ71XDhwWmrwwX04MLp6Mfh
qIf1Hnsak4sDQhZEjK5Be4j3h2CkLherFmJuqSaDMJ1Bdyqmhq4bMdFZr+INDltg
b9II+mzcvQIKm/8XG8dksINSQGXt67xEqqre4qF1Jkst2jPrpr36qWwfO0mPswrd
/JmM5bDEJSJEuZ5AnFbfw1vhmCJrlYnUCRB9F+0SULSmUlXblbjGFh3iMdFeT0P5
ZN6qwroxsuI35IYcNXM3/MrJmNKa459/e5epQN7Z9A5kHKmwRXmwsZ3KOPG3KyXI
VVda63xih7LloKsi5BWL8tB5yCaC8I9zHOs/JP/TOWK2wC1+Ah6jBWRkKGXr4Vjs
poQnobDu6D7hOdfsTFx6c7tA+CY3Ja3pI+BglssPBEHT2uqw0bYgiIkK4dZ8yjAa
7VotWyjTs5+K59oHuLgnrUlHOJyu8rZ2Eo/GSyr1t+BbyFmINkMbtLlhf56SESnv
GhYEzxO5kSgHqwPgoMor2w7YaWfZp3rYCgCWa5zDfLaKLp2LP7s+xJpTyUGg+3Nn
Vz8prPCaadBHtF7hvFPLp1hsmbWZecWM/8ybGzVPzSN3aE9KMqiOFPESUXG5rtXI
8FRBtKxTBASi30ojMALMxvPNBjUoIS0zKYLsA2dVfKo87PM6nSeJ9IIBtxZN5dU+
Gvws1iKGOiq3Q7NUGvYy3+PtU9jr8J9zckYjqv7XDsl7iPNLN/bvMOQoSFsB7/hY
rln7Y9Ymn1pqR9Z7ccstHxHtU1gYAuLYvUK25IJC2CiZEL+ezLzdHBpVi3a3PpZI
6lYR3Cqrz3GAiiZ3gNsLyoZl/1fsxF+KuFmy1tm8OKHgXDcf1MXGo+8CNmUBdDBe
tYXkRsfEz699RYqw9Bp96OcP1LZRiVPJLAVskJt9JBQoJYtBavkjaqyHf13vdxT8
09gOrV/yEOGtpudSszbl3yZGLb72WkKq1xzHHlHGj6C8UyICUKJpSr8TdKRKAefp
grIFuqsnhDRmCqUw4pM93RSc+V+4/uVoTqUcpM8KvdD9tTUPV6hnRsqwXVPYcL/B
Bras+EYFElTjhs1AWR5XyVSvdSfGRDfNeDmz3MbgmNcaSDupdUntw7znePjLABFy
3K4ouURieGsBlW9ZvcGhqLvgZBqZ7OS+df7htXKYrGXef9MqraT9uvL3kabp1wbA
PgjLj3irngfjiHvT1vyZR+NV8uViaphqlVHbXtvxJSZh2zt49b1HBxLp9XqEApNh
mZw63J0H9CSGHr6fjk2wRl21msblW6evdbr+oBJDyxAKNsgn4XmFpkpRJ3zSiunh
x8IC3t8iMyjTOKwhtoWF35/qQcFVd132FWCw+XG1q1CdJpBxcvt8paThWOrKRLh7
AqjicZn4/tTvRjQAnxzuX2WF9tLxO6Nvujl+GG0tI57BhZAxDXmHgSIdIwKh+Yvw
DkggvCU4XZ19QEPM36+CudFvEHai3x+CQ2wBrZC72AvHw0Pcoy+1rBo0c7ww4VTy
+UPwET5KJs2bqk1Tt68HXnCcP7r3jEyiigEgP8vmY173526PA9zdbMaB6bP00wFR
GtS+enXNwK+bhwscViOtK9ILBN7CBvsdVL+VPBJPftNlZUdfueS4IukQNBXNib/z
QfODy4ZhPQl5O1bqUVDXK73K0BCMQY/jM5UmwEpgFz+Am9zK/tyilnehafrN2JnV
c37ePqREj2Lf30W4TgyAeQz17MOlrJuGvX9nxQCWxrUzyY4KdSX/bsmhajezpDIp
gH13nnIe5Gmo/67P57NO0eR9n9bjKT52xuUEV+dURxeq258Uvf7iLXF2+SjJ/gQD
V10BMz7tAk/lemtaBm+zmLo3gJPFv6Aam4huVnQPNxeJrWbEt/nnA80F0xKUW+Y8
RAAA8re2GNXTPaxxjilSad0qitAZihgDE1PyxA7EyTiDdFsourV8OI1mTuoJ+4dz
eB+vxblwL2lF6vdiBhj4u4HwQdgtq3l1m7YuSzUy4pKr+rautsZhW+Ra5cWiU+oY
MwhQH2MuoLgnPDtSi2MrI++Vcuh6f88J/C65AgG85Vofm88KXb4XIaLMZjWpva0y
IkaQ2S6tgzqIvrFCNjoFFOJnxmdEOIsl+Kpnc95Mk49yP555/8l5ZHdFUbSF7dx4
/EOP4YShKSr+d8WVNDS/SVSBiMh4zL21gVI0khxbqsGBzovfn2TJNS7/ydCGK3ou
QPaRrxZkA9BjaLWYHMcgIGHdOCPn+iLEcItHFMhswPp1npW9EatG4/KzocAgW+P0
K8Dhro/dL8Kj7ZqOjAVBT5534eCfUhNCQXSXnN2EabIGr0cqdAOjQiw5PspaMgG2
L234FLjnynhS0cEsajDaATUbY3ulls2T2ygPjXXd8xI98PB+GQ8p5XqjjkYDYvhP
54MK2ggajn5TzH3oA14n98nvO1YWhaJ17fxl6gnhU88C8PaMdQQYqB3eFh0js5Ou
bIy+0v47ndx5fLPHUzb+0NCkS4Zd6o58eswbpQy7g/guWf0qJh99ul1HnWy8QYVH
FhAltUfNOTARcHjOWiaBcgVDH2OCCghcJppWw68YutyO94jfD1aA0xX2Ar/+nuC5
s+Hugw6Pzit8fz8p0G+PNXZVCHBIh8kcwHiDF7Qwdpxsq+v5op9G/v9aXm/XTEPd
vjXb698Nq8n5kDcpPV8TpnwusNd6bYJijnIz9UjPnXsc2un2P07qAagDwNIEusaw
LvDZf4lFKnGsyVnlXenCiXxYv+M142tgITAZS49AqTMo8DUiOy9JgNOBwHw2lukq
gD3bMZBF7vic1tZM9cfnkz++3hiNsYm42ZlXsEp3/JbgToq+KQebdMP9ZCW7/J2d
As654KdFZBvrkHhnm2zyk/my3lI18+1vbmvUoS4E5Ee4SVWGtMrLP9S4xlD3r+iF
miZioGIntKl0b/Wu/VV1TVzrLGR4+FewuccDt6//Kz91k5NmfXumh3i6Oe3KtYII
8kt+1QMpG+KMG5nykdz9F48iGRjE3HdE7EHrmEwJ8eQtQUMbtdE3o1BWs0oRWBES
YT3Pm3i9aIrmmwNQPUy+y8SUDBlZGIfwaazW/H+v6Icb/ai+oM2iEDJy6ybVKuw8
dRziKQ7eDJQ/hoAtYYaKlLSA+V07wGp4/ihHkxC8vzWuUj5mfOdPgOZ4gtQ+Mm6q
OGUEu36f7R5XDaoArQWC0ZJk8vdIxyGYtC8uruLvo//EUzmWlEh4crOdPJ0GsDwe
q4O8Uv5/yQaKQ4l9lNCXNasoPUF0d/JZNO65u947JwEBeLPoBiVECNYG2Nr1UxBT
IBfxurr8BE+4mLIx2oSBSjoDK7Nwj8vmEMdL3H/bCItuLX7yOIV0Ky5+R3Zw2AN7
1TYqQyeiJtjnYVSH1gPjDCJVme+OKXSeGdzVLjjUo8k2S5iJLUGdjBCo0dG/v5e4
WCO+vo3T1SLvjgLpQJvItSzcY/N5MsmOXxCRqoJ5qYLlE3FQ/jXr8g39oy1R6XJO
69HSJC63MrVeVL417a9Jjawe24voAlNA67YsnbgpvvrHgvEO+r250+ma0mMtC1BB
6mYygIrKx9TO5bfeqiRtu1whHjBKw/0oMTbuZS+q0zt+xeemf+jRHibM5B1YOkAq
9ddR+uwo/asT9AK4Ri7ai6ftpuVTxAI/WekMUZlsjbyVWxpvpNOhwHsHKeWik8f5
mO3mfHBCf9M69/zfIkrtGKgpmLFpCN7fh2n2y6DFAKnGrHn/vf990qqry3NoOOHa
XjgL9QdsAOXui8qLTFkEUw3nshAxUTV2aY/30UQR6PlGbD0S56vzcX1nChZVgmPW
yMCQcwvbkJ4eICA/rAoI/3yJWZHc1AnRHYlQqGlBIlVV4Uc3Y9SNjK6w2pA4lRyJ
HZClkA9Wi7Nr/gAC2wh2ylBgtepMjCSVCeuk7KyU1NmE7u9RkI3p+8EsxhbAWhGv
xW1+HIjevq2dbmO7TkzsT+ErJOWJOVeW6PYad+UAppjZfH3UPyoNY8pHK5yaLkEV
bbmo6ZWRD+fhSSmeknWSZmt+zbqo2AEl7hvIMdWiEXRu2U/PM+EhAzRdHTn9djOK
xOoO5fJO1yosZOS76edaUx4Bi/LQZt19SC6gqUXHwukC+fUXoeBGQQeYFlUvCTqz
GfOYqtOPUkLLWgZRJXUMfr71Wj7I9VCfXRMRKExRM5nEQzzOrGihzD5UaQpa7eRf
rIAiTFdSz6pcP9jsfUL0p+jcPQ56aibiJCsstsP7KaQfCjnf4XazihiDGqkbMniS
0NcWTUR07Bb8P1XjFQBP++5reTZo2SAJySy+xJkbbVJ8u49Es9Rjfs+lxwxn8h0i
ey21hlMiv3YzU77fAFXXQO42/WSU5HnMnZI9LBn7/qCXv7IzKphb7jJDVo1KvvIL
xdYCS2OhB2cXAbbGKblxYaCfJd8LPBuh2YA6yjzlbMsgs0dKJR7SSiVUT4GMlX1Q
IAcwRpOmBUDcarBTIxaK9IT6ANbmnQhrxRRr6lyUJuMYFBZipprveSCUsDiztfIO
2BQi5W29cTmbAwzoc/PI3VJV0CZ2px3379cC9RTql9bOhQTmGNN9tOyZDkjyfDFq
Cs8EJl3q1PhKrV4XlYSD8pL7MZ8ZE+Q8ovROjTe7YOTU7ILSsWYSko/RBu9+yqIe
ZZ23WebIaeGTpsyoY99obFDyhvQDIU50rgpHxMXGhhi04T+KpyY+v7KTzksbb3h7
K0MgE6YYUiVlWJsyEz+5w3ZaVxP3a+3LQoqoBHQrknLZmbRvxKJXN2QKpMSUkBgv
e3q+9lR2I2A+L7eFCkjaQfzyOOd1BnkwFcjH+itOXSsM5MGqmvd7gnMeaBGeshc/
/htY2+DpwJMERQbUnuJE195E8e2XtmvVXYHHrCUslVc0XWfHfMVjsNzfduNvrcS1
5I66RqaOis29SXwB5o/MS+5/kVCPTPG/E1CFmyEDSSb4dcZ2i6LOHRQ/i4bgeMk9
ZjxYgwRal9AcEolUvS/HfHoS6Ji2/4+aXpb5CqENkoGDrum5hf2WiYxhRqQZvIsP
Tcv8y6Qpe8w6/qCrLtUOPAz/7998JU3ck65DLII3FFg4LeX8NDY4duJD+GeDopxL
T18PN6y8aZ6RBYfqhEOyLNI4i7ypChieI22fqac/JXJQHK8F+/YryaxmdqEtH1u1
fZI+cZ+JfLaoLY06hcVBnDZFFGqI0jETmqsEd96cNBVydWJ3zi8BjwQEUTveSRBb
0vCAvzZQIMKG5PhyFqNxqiJsOgf02zHR42G2Ro3jiaib6dA/QPEcQCCBhrIz44gy
RQrL6bS3T4jveM70uaVyqCwzbLYvXlti6+lmTNJmyowTMcJR0oLWqzq4cVAL6zDf
mP8Km/Kl2nJW50I4WzRgiCg/lWBYpaIFbPlBi2I6jbAn6hsx0Bhpr8FBO9pWHRTr
7+zHrYmSG5fdD5CctGVJtCbXVyXYfBPnEjS43gUJup3Tw1q4NGS+SsS7CZMxaD3g
0XB0HyQ6DSEbu2sIYGXTzmeRtoP6UOCeWcH9HF/2KjuPVdTlSrq7d5qNGnOI5zCJ
fWuXjudKMhXuPYE7lATe17VTBiXMY1+fsQaSydI0R9+OWA50pEKduPppGiEoVllv
9hkOZkD2usNkkvrI0F2ClLbveE/tkMpQLh3Y3N8rS5maC52JWiWdGIAHxzYOc8P8
Nnqwf/ov89lq8uT+PMvepHNwFbwlIXKaWQWyISWIjxul8s1tIONv301MaM2aKLCn
is0VX2mayc42Jyhh1heXA/xHQRmPQCj63SBih2e3M1DmQiaKG9x3qSqZdtWRBZlu
hp/luSd4klW8Fmqx8b7cLDnjqOVaIjARh/JUwlH18EFyZ18PRxbcggy8gM484PtS
oO2ojF41p4+auoBdyu18IvSkbFAWxvSlEn01pjewmH9UJj73Uogdn2ONpZgnMHMC
tx3p951asxFgwzp42OxtVZCw4FZMx0nlZASh71Ry88ftJ/H5wrWdgrjOO8ZpbagG
uY6vgXv27sUQCwUTj+uJWCk056yIXsKjxLqPdwBSSjRJDZUqhrLZknp1YSiiEWw2
bXg/DBxYJAxPY1K99gZv+xgI6pRSGnvvVK8fHFrEMn0lnL+WCl3XTpslX+PLAZ2u
p1ZEpq0wndkgRPko/7EOeN2aq6wcQfONpeRXz+lw4sbJ/oxx52YigGmsqjyJ6yv5
EAzJwv9hRWElvLXkNIF+5EvMon7gz8jEwM5PWgTTKgSwykitBSTnXHNkfeotnyfT
SqcwkVHLbCVgQa2S/qtOw93o8DL2S7/PU/cJbvPtqBB4K6xGWoTzBnv6zNitL8o8
wQVa7WzH3F7wjHPc/ApybpEP5HjKC48LbmZgaDqwZbIGMfB5Qctu0EUNb29nyYN+
3563OcD9ncGm87I2MY/5gsxz6jGLVUyNKWMA8KKx6MNXFaGbp1yljtPPygjQh+3l
4ST3J06d+oTuRfPd6yA5Aiv6BMb5OnkZK1laAwHHKqtoKvU8WBF+gSFJsf2U2jiF
r+7sV9mceJFXPx7sAxF+Col6+4cziC57YLT714j7sGt1rWpPvvWulqINPlmYcNS3
qg8gVrf5MIoOL784AjQ2sdYcIY2S8h2QKFprMjzUm7K2vs4JzFHIbN1hZh/VkYMU
k0vXx742JsMDZV8pshaxM+9j7HjsJwhx/NCmrPwgVJsxN8ZuVX0LcF75I/j9cHR5
BIHXy+6Z2Wz8pvFCk7neFzjDu7xt1x4tTSEAVnfQ9MNlSCnSDPvVFH08TyBzTwVl
2lVILNJZj9gxtXKT1eUTHnYW7Qypu4jXzwdMDM0/WiG0/TzCOn1H/d7ihNf4t780
x2wDvxjmqg6Jm/5UpK/GTF+MnlDCVmyVSfWWmKqAT+zzf8yzeM9WLVwssR2oa8BI
j1bg2nprDSqhQIXxpripuC88eQucF0ABoUgwWZrp/EG8CQ6UQjT5nhSDDEEv2POW
SRI/0H/2Vzx2Y3FS/FieuhhTWGNjcpSwlYVMUgYJ7TsW+KOAWFxPsmbUQIaLawRE
ITzdOMPTZ8yEyHMaHciLt1OS2BF7Y3zHT22xBeTyvSZDSyM8CobHZVWeYwAOt870
mm9KuRo+Pf+yVH/pDdGb0/1Q48krz8+cdQEcgj7jmRQoRbi4lZ2u/sUMw5Fqs8MM
Kax20BeC8JWRVI0YLZdqEEOSS9pdo+xS9zvT7Ki531KJwn5GZF9udY3taxZmvNaz
AFL/EuYp3JMBeWWLDPB6eyA5Q9UxSweZvxFLiHm/PJyMAtAbTR/TXQPxN6cLZdYZ
iy8ch1uXg/b6LxPWB0muYlSA9Y4NfHDCJcOjPWB4YVuoVfXDm1ATw1cWDaiUoaIk
0q4qau+juMK6GBu7UO8clWCn6d8DPs4MRDjN8cbVtl0rYLt1d4UVosCbfo/f1xd7
Q/Hzeo3Y9SyiTc6VvkoC2NYJU3kkgpjLoF9uooH8EOeC6uuH9YhXk81eV/QU9p5Z
LAqR6PH3Cm8E/H5ohfVyAAu6g1jaK0TdJR3r838NDWP2G9Ytb6zrfsl/AAgEBwu0
BlwmqmbPSY+0pb2fwQ4NgP26LWq0vVesmPpvE4N+3rjMq3M3LJhiFyERE3bqdEIY
8ebzWGHOSvL56RXG1tzyyTCSIhDHDjtcVTTjebRv9VPz7vYzoqMyo+u3jtiFEITz
1mktn+B+91p+L4b6mxdwMR0tm4ObNGGHSyq99eXOdCgtNH9MjmZPFaSk3Hy5kuQ6
JZH42SYYepFgzkdoHuEcXJLYJDu7MqzZOtltkJLIo0JFY4rcqG9ouWZbRHmm6pMP
jjXfzxrvc865MkdeyC9aNje7pv5yU8BzeW1nRgdp4k9BoV8c29R+sM5aDSFQgFAx
nk7ak4GN3lYhtcmIjvWPEdg6TfYrj5MKLW+ltiYWF890XsKXSJGuQFsGg+PGul8e
zLh+WAaBYsjcTo6LF+4AlzgmHUf0iHruFKiNt+kobVJW5dnom8p6qlmoh0WhI5sQ
jAJlfvxmZG3IUaBSnpnPvvlUYbGkTzBOoaxtvczD9AGCrLJ65u7dnDqI4AC8T6wH
9jKQOK7BjKXm0dLZv4YkdvtjfncHbXYHEmUxyjs3m1+F94Kvcr12qq6FQx19BCOV
VAhdsybP3hXFdy3k9N3zpZXE1usQXSvSyFpYQc1kccnAbceq7VWKx9n6ezX5JB2E
UTFKVu3Jl6P8OvUbQ39NyLgZKf5bktcjy8UH9uOe8dEqbSb7lDjbc4OSHl0rN0Cw
T149tKfsPm1xLnNVZoSHxYHtyloLGklCeNobrpd/0qkf1EVWl+HWokiY+VmB2oOk
213zmPeLx7JHjgZTSa7Kv2pnKK9VZmBqzybQnW5b30sLHjezYzlfB8ou3wIEVqMc
jsxn6XQuOG77BHYA6UAcZqn2xfpkJua23biHAMRxK1sLnEK5MFPYfr3OBN+ZqzBb
bLquyOddoueyJhFAbEb3MW2JMJXddBLZRoo8LVPlgQXWVu/M3r/BhjWssH1pfLXH
WWcr4r0U0tDnza1r0qbNexYUg4j3VrJ8vGQsNX9LH7h0rggawXZfE2c2XNPpdTHX
iojczCQKZntfGLhELQtS+FgjUtsg3+SrLC9sDofghNm8MgDdeX8+CRql1twqVILs
pfILjv9eqxOJbEouBWE17ojz3JleTMoC7yM6kNsjMjuNYGdCD+UHV98YKOtGp7D2
RPTV0ANBKNtV56Sxn1AAmtd8whG2/itRPj6xmWsCiEBhV/6Ja4SFdezVf4wON9C2
NuzlYg7bpMyDu/wZB+REunbqVKYxy+Bk+hyzTgLmAtAD3iQHQMqEAFW9+4UrM4C+
6TfOJxvqTAp6urgnyStXCB1AihQjbRw9NdL4usMyA/gC8Xg35ffjGf6yUPjox5Bq
jh/rtbOjkcNlV5WPdIypxm4RYJgP2RZDiCgcKyrMlrU0XHi5W7OoskrCVY3Xpve2
j3dKGSeUPQAUGNMbxWrKCnQfiCc/5CZS4TUVHzcvQzK9yzKHlSj5Wdao+MkiyHXO
H7TNo3d6kfpmT4QIff2LZZyRdOF5i/vstiWnD0MJjnXeNpwVUdkOT0/bs1RTg50f
mmkbMEbSqsQj7rQPn63jfOpe/ZsOeTYmnhzg9l+P90HV1xYAgkd6kkkTnULMSrFQ
hGEPpKwtYZt+nOpD5TR3q0MWfUH/klp1DvH9MbYjPNgJlrDyr3VAxqgB+eEYnE/7
eB0HGBHCOCAmwx2FoFFJ2k3fyGRH/sTACzOcKPNCeNH46ay0OMZ7RLAxvHK+Fufy
4FlEAgXGjOUEqQYp85IzUDsuQOGTHwweHAJf4c1BR3FA93UZunal3qXGjmpvI70K
5tIE6/9fBxFip6D5r9tWp2Au/9nM6gf0DtHbbjdtQHclPWMCHQPrWXcOPe+0Tw6o
BYUunTKAkrWNDmopMNjijWVRUoarn8+DyfOsqbopYsLZKEBFmc8fzXAWopp9rsZx
8bSNNdtA/mL3ixhp9nn+QY8aZqAkGtGBzu2X4KCUOZunKBt2AldfvqonD8CZaEDM
FmeW+Su9K+wN9+aUDj8hXwqsPsdp4D2IKfYMuWX8YZJzhRy3QDpdNXO01Ze2foY5
Gi1hcLp4f95sKP2SbZ81kM2rkj0sNp6bIE+K49wO5Eo5TX23DgBPqF6i5H0HeDhk
1+FkQuEyTEtBIc0B8pvo25l3Gfkk4egRJ6OrRq0GbAGwMsjO/LOPbe1PDwYqAqQR
hpVfKfDD58jJIFMS1KXeZzhmYAcajvEOQkLAf4SpSRd0GntOPUzrFmgydDI/7awg
DFLc7YsjNw/zAwDAnEX/YqGK+ut2C/IsFy2aNKs9ZXmrWAptG9RS5OJpLpJSE9Ir
ifBfJPSUKi0jptSXrEBA29ZU1s4mfUTErX/DMixds6OJQSgpokcq5nQc7tzfwFXZ
aU2smYqCSUhZJ5erCuPODmz7p3XXs4hTnpwukal45ezHeCC9RLFPPtw3XDvLAgVp
PDxdr/nlBqCaJN6TUE7atICgIkg+Z+2nxsSLJ9bWOQLMpI/sCfrIHb3qmYMvYZVY
rQimQnQCMxShPrk6zF7016NgyEzS9EMQCHDoMi+9CWAWONGw9Xn1NFdtHBesn/4v
iW//4Uh2EgLBh/S7qGz7YLAJV3ZwprzCqKdBBwJHrov86jlXfQJJeUj0Xbss7PHx
v+YZWkuJY6UM6YTFVQCMsy6yt5AzqS5M64Q69gtzlyuGt2/ec9nOfM9h/esStNmd
C4cmMxjgoSPJmLBdWNlplLC3JWGp4E0ErOz+Oad2hvFGIOS08tWEflpvfgalXun+
JDgZqiVOrnzc42h7TmqvQfAzpO1tp/iWz6hiA5WyqILbFwD90iiOVQstI4XFlPLB
+thEUmu9Gc1YwEtpCXCJOQ2NAYp2wVbQNj6CuS2FzaHd828oEo15XkOrm6t6Ih+U
806emxEnpOHnVb3ya+rm6NWA3uyi0Zorg2KfyWE0S4v48uD3hUX+/xUBOQrzGIUX
ho55B/gkZDSjf06iGWG64g7CN5TBhKQALNJ5aywFFnz0svXrZPy4nFaqEdN5l/H0
oYJptRBlO4u1c94TLSVo6AlIquZaiF15Z27zKHeC8RIv4U7dwY1/9n879hdG3cih
opfDQY5YvjePM9duIUVuArfmKzAvOgT98hRJXppIJc7H7E5dC1uk0fuFEZBhF02M
XK/CW88kVQGeoHVTA1dom/odfmZC7iiIwNbSWDp3VOKW0inSKJaq+LRZYXk2xUxb
M5ShqO+KGZorHW/BkjzxyXz0st+24XlbxAB1iE3WteYR+b7ckmcaquc14lKn4XY0
rFJ/xE/nNIGdMzrnIjHK0oIG4BIIvOZfTuAOKVVUcx8uGbO9se0FETdTluDleYs4
IGSaYOhKULFn8ugw40kLPtl9ouuy00BXiROvr2+QfswvUMXH7n8gZ81dI/efuaLq
VB2p/fbZ0mpSEkAJwkKzlH6DXRTsmYLx2eLpBAwyts7PoEMlz3hYz23DNdGivQ9k
/lvDICurLbr0I0yXOiYeniKivJMPy67nww57ZL+yuT+Cwbq7ipcPNJN3x6ZmEtcA
qTR0MyE5FMFow4Hx7TfdXFO708Z8eHFbaho53tvgwBRxEzDKcdPHR/Yh7R6zNwzv
RFz8HIqaYmcMKSsSstpvzCx/Dz+YFZcx0DSVIHUVplgVu0Ed4UDiFzAxT93sIhzu
JWwIWB/apahYPgjfhgFk5NNhQmYIG9+SMqDKqxEMWlzj7XyzrdnelqnEgwkiMEfg
YlKFUNgRufH4/35C68IhYnLi+xR8D7sZ5hg14tDVshvXRSXMoWsua1KyxfZkBFqR
/v0A8HAvlo8bPk9ts2pSVrK0oqxUg2IzAV4ekqJeVFGZPuH8D75kMhup8/wZ94CP
NoF3kBfUpHcPBXiI+fw5xNXAg3vFTghUirKM7BqCA8dYQK6lLpeb4/h7VCsYwASz
VpEUD7lmI+92u94y8mwWAcOEmjlQxsQiQxzs/ifSgmcpz4077ylpC8TMcbtGer22
s7P2yybOOgRrvwNLYUOcXEPlxUHf3+Z3qut1fGgTM1OBzCtSs7UlulB4qO0fa1JA
0V75c4T58C3tQ48m0pUKWT2uzBtNlh4ha3MgAJgILw6aXupIQwqK1pR2NW/GE3C7
M1NRjbYuj27Yz2FLCr7g028Mn61QDbuXBiigrTCLIv4fW5p7iQJ9cmc30r3Zt4RR
9Lsjry5AC+Vs22y7D25TXBb6UcqjPapaEXtm0NXHIU1/BnSR56tCpHGTetFHHvxU
vC4G+vt0Y2FDiuK7EfbHulSFaXFb7Z7HFZ/ZOOlOxMXT6l/X8oehleDJSWw4ejKQ
yliEwwnu6rm+xChLt4Ivpw4TzT1UF0Q7g6Z/10vuQ36kq5BdPqrp234sTnAq+l5V
wUzn48dYk40Fkhb9AkDpumwDFSt5JHh04Rmqw4MErZJ8lPCu8djUVj1UMm5MSUha
ytFDeBwkaLItxWEo1bZDm7tQbuV2vZjrtVMCQO8oVXXmG54MloX4k3dt0Dd2dSRj
ru/cQjMUhzuFmeIVpRd8y8uLOklAivXKK11v5GQ9WamJjnmYqKlYG+YFmnMwVxZG
vS0g8WZk7B/jkYKylyehm0ZH2cFLqNnVBMFSOzG6+ouBDLWgITPcT4F1S8KEKEz6
Fr/PFtxXVk8VdBe0RhcoJ73nITkTNPzJFs7Y1YnG1HSSJ87cruWIiLsineq7/ED4
QPW+GdgqT2qR0bHXTv5ARaLElQSaUCwQZ+XTm6MGHGHnLh8n7bi7NVngjdCfeWoP
1ytwEUK450qigaRisuoYdhjmKSj2jgn8AsA2Bdxp+/QKKUevshUZl1nwJljvyG9n
HIcPzZURC1/NJx00N8umUukVJb0N25N9oLyUoC8kjjWNnO5f/7CtL/nq9mxwcJUV
oiYWQ6+Rdyc02OKZVkt5yGUrw/1XGmJPjniTINcqHRkmJeqC5k7Wcjciz32DPmPT
Ehpcxxf+QEWqXP12v4zxDMlrnS3hYcOp0kBBQ9lFIXocm6cqByZEpTLbL4JXxC8s
VOrECpMGDCewRsuMBJ3zoKBDXHX2ELV2DZZZbgn0L8jb7lqzxzsPlu/BSvpW4onR
PBosPk2WyycHfSgQEfOhEeu0VB1z87DxGBnWltgzPG/j0LUyqVVEID/sub1JQImn
0cLPHk+ZuKmTFn7XAl+wGaSDY6DuGUy4jNk6QHvAas7yZP6yRvyXqjLDZEkX4axf
/lMmi4V920WjgMRfUdbctSr//0vQNku4QTiH19zHQaPnry4IcNxygsAHFOE+DcCh
oYCA637RX+HIgQHCGNX3sDEBjo17EUoFK9/mbKtwedH1uYOYL6B6JXQMN3wxreYP
NuTQ1v8nwduQM0kI+FrY2lsNMDK/5DD0BEdxti3RuUc1GYyeD42PELyZO1yad49H
Xh/fy4hjC4+jjGHSp+meipGh2WbMIFOGaGTE7kilX3PGX5LpqSf/K0UYU3FMxKdW
9Uxs2WpbItMEujuvaQAZBxAhB2jSg3MlRFi70xeFNMC9Nmyg0NEynKPxmR9qtqaZ
VT40hLamk4pAL3NUt4IQNmXhaU86Dk8rkAZpu9t03WNF7ynXdcdV/WJJqH/zseRl
ugrRUkP9FcDvsim2halXzD2p/xmT4NI7+DPOGBANuR8Xh4ohBDVSY6axSCazA921
7yHRo3O3WjDQE1y+BdusYdnplmJRv1qG0nm6+5XgIplkQqENAqQCrh1QKxX40Aps
mCoK8C2gUTxnEdATC6kuQb+Tipa+ldVPaF73uIsLtatD919PHe2W97SPzyhJlQQ1
j5V4UxtGIWLfJlZ3+LC5kkeRIz6/RCmuHffk1dq00G98YtjMO6dwWllGnGHN91WL
ALfyQNNLhAbpvZ/tfuN4hDwhz5avHHsGZjXewR/1RGFHdfAeGJLR9eZZSnGAaUsv
zFx3nyJWFR3tK9JHg15VJHSR+USaH/qv/tx76zK9TOgeO02PR5HntGbTihCyEW2f
uiSQ28FTmy+HcRaWC8ve7RsKT187oJjfT9vuxkJDAHsF/2zuomDCHKLXEGCGS3l9
94b2vhqbrFm5hzS81o6m2LSvVxJxPK/8E+uNToZHAmQ41Np4/P9SEfCnqeEQmiiW
83uzYUG4kCdAUwOfiwsPnKopl5qMyumpMgLPiouvFzMck0CxqgP+6ov7l8/EGO9d
hltn/35zXQRkzaVpdDYj6RxAqyOAT7+zHa2+yH8g2/5URrbwcm39XjYRAzhO74+P
Zz+WUavJ/379RnpC6B4Ozb3lICiGPJ7V6CHBLh6uhv5C64jlUwXQyB/aotb3J4TC
9yW+EG1IEepLpn6Q8qdhqMGatpAZ2LSdBIDsHy+ilZTcdE1MvaaIArFvzwEsZoHh
IaxFOsJXA1jxmmxsrMenaDe3fEj3UY3K4jy55o96ipf9iq5dcIEuuVa3Z5PbS70D
c9ZxKdlZrNdbicxIlWHFM6LAdyYvv9ZjIGc4gJUW13Nt+bb4e16nrrjSkDVFHF9c
CGPXUnc8YiylmnGBWoMUpzN3KCvPs/YUrCISOUyEBDxQowzeus+mCznAkBIemOL2
YfAzTS3O1vLHIYsZaTLttRFtRlbgSstrsjQ0Po51oJYTiQIzbZhJ45VmzoxC6Omt
SN39u4Ru45qEb0KHSVgfx3VzdORwoA47hFYnXo5wMpvfURA9KqxnKnpHT0YUXcha
d7GIXPONeayNHAMRd6pjjXXAeieYvi6KBopeEzjg0hT6Lj/T5Gtm8dfylg5L2cD1
Fvap38IEtE5Ad/H+WXSeZjGNbZDOZyYHsEoXGV1eAftK/mbJzR5/9VO/G3G/tuV7
vmlSA75ZfCsg9Ob3H7OYf84eYQtrsdX9jnTPT8p9IM7a8S734euQcc0ajdBrCta6
GY/ubKDGLg5jHwkh2+kJL1v/MEvflv1WNgzjgslbnWCOK0hVWrjrCf3Jph9kd53r
rMbvXlBrCAolB/cIw9J984Pw5BgK4rqAijWejqVzRFsBN8dwxijAO0jRZYkOyJE9
HEco5HN16uTC2eGXK5PtspOrF5DoUC5qxmXbWGQUL12hwQYPl3YA9jizof3AlNSY
l8rPrSeoSoKXTJVe4ZqeK3ghUtzlr0YMxaN8vWIKsTOcGnR/eT66D3zAWs4m7VDu
vtgtyIHpSRdzmwa/EChduLsaLyqlr70cK8InY1Rm6I75c9yd0PzI95DVZgvYyynQ
cn5gXgeyQmq33J+BLcrjPidZyRlhuIoB7Tn3NMUtlLLwL4dhIZuwY+MAdDZgpEms
ApNs0uqAPSJd9FZ3iVT8toZEN5YRrkoWtt5b88wnbCDnGkYMiJAVoEpe8iXUJR6d
idXn80bKBx2R4YeBJifRjeO43w3w3Tn8hR/iDG/+SeU1f67ww4X9a5yeyPo3u+cS
Sn2SAGQhxqd1R3xDs7BzovaLbeyi/xBo+O6WEygj2IKNjzoe+zMOYwwfFNn3NX/y
FfDx7FbXxaNI9LR4W1LplSggTK+IcaIJFpBsbntagNlvAEAipa9QOYQo2U3PnhH0
wVQyoIh8PIZzXrXjAKBiCzBo8HSOF+uO3An3xdNWj799087Tpp9J9C95N+G95RGy
Vz93HZcLTWmL7Dbny+mVfmAtxa7rzKPxdhxnJ71aIZUimed0OevucTT9ThhhG2b2
kJz4zGikcm+GXfR3pZrfAZVAf6ylzs0vNCWhyKee0T85uct495VfLtLWFRJOXBuI
+M5M3C2YyoPBP5zYgmOj17w4ZW79cIMerwDqJhPbtqq47f0KNkRlonGjaEQFWWT7
dIU5Ypt2ZnC6iaOcw2tZe6zDVDQ8DLBbRydQ32vPnD6y/C/FmSTSSBH1g4lJEv3n
LI1IPULF5NHTuAmtY3fD6paxzkllnmtVOPYjNqaaCkCNoeVKAb1WdptkaKrs7vR0
XYijyMA1PwBnKKXyyHzatDpcKOQLu1FfWlqQl+A/n04T1685MPSj8sxb9qWIw7qL
KLz3rR7qamA1vv2A3xK3cRyT0n14LsFq0fheCAiLLn3PS6pr3ZZedB6Yo3+w+D2t
GbwwH2dUDBQGb9HAYdsLWwbybEL7plyuKFin3yUd28jSHRjGGGSPJwgJzWzSWDq4
TGna2RPq6pSgIVjdUf3AmBHgzxl2t3a5458oLhqGmFBUyUcr3MOwrXului+/PTx+
MmCfaTXGlpzt6yr4JWYwbHmZs02JiuPTi++bEw4gKI3XA7Nh7O7g9AZxVSE3g1ze
pJPkSsa9FWQCUIyjieHb51EH+WPqQUobGcRkm5Sh+hJuFQDGZOBeUhMTnBlFlApq
7rB1JXP08PQH6QS2N4WhVLeWVet5ZxmFTj7KizJ8XLl1+q2pGfJ2dJpwPqiv/aTY
rb/cDGMenCZp41/Sv70RLGhyXp2j4HXOw7FjXu4piiqvvBNkfXHeO2B31/SRBMqU
dwASQkuB2K1suRcEnf966XdiONkW+kPCZDcDvsGPuSpMc5KI8Epa1Dy48rmnB8yd
7V5ymHvBcYJjYzXmkUkaZdt6j/laOpAR8J4H8d6jly+uE7Fb6/bb+WT1JORSjVOf
ZHXbEqs8OWa6ni6Uql19O2ALnYotRR3sXhcXdJoEN+wYT7r47TditY04aDgBV3Hx
jlEyNAdxop+MG/fR/T7TCYEY8JI8fabeV7ugvAQglJZZIUvvhkSTnMhfz7WlHL6C
w3AiMYpOGVNbSaD2T/g9LBZ7mFJd5wJY+/HzBw4o39zUy888q6fnanRlYYr0jGJN
tPULtSDd2uRJcna+s6JAERpkmbExPrOA6VUddPPrIOQqIkjJ8rV1s7xa2hseldth
oW4YveIlYE2mZF2SCA+aic/GIHdxk6lkca44sNlDm0v1W+FvCdExUr13UM17NDSr
CkWE2iGs023QV48lS8mcGx3/fuKjAhmkhLXsoH9BssXSK7TiLkHSetA+amxorzzc
TrCZhfsqrN7LElf9JMqRG1KSZj5euJpNyvFPEilR6AwWOuemSq0Tv91HcYU+lNCl
yclBq9pOOvShEdjd+OI4kiUtS2AfR50eH4KSh2mr2s0fkGcnO6HJXP5TW+ci6Lcg
4SBCI+SG67myCw07IBXSDcesch3ngk3nhnLdbqDP8CQpAEGr7hd7TaNw2U3I9lQ3
Zfbp8UVNoyDUFTgC4zxWTPKUmyuIUnu/9MhA3itLOPkjYdxsu+b8D6DQKktQO6xx
EPtV9gVdveKTQIL78pqMxwwEDwddC3v9JDOt3+sAJpzUcEW+KsKgnCDtvk+WIFHy
GiJvqcMpWTZAgbGN9RaI6Z71W2/h5ZKjf2OzRIWaOxZU1lkoZJnZDYWOnzdayvRb
DWXcFroGI6U2PR1JJZV8yeNrvePmTcOyUSeO78veBN4Dd6hHOH9Xmfz9WuQ0xK8j
9c9mNb6phXSiuzwJ+Q18+E74dZ6S5Ka9Nf04wmok2ig9jQFEC7vVyt9PBukCNeyH
V8Cs2EbsR5Wr/oGgKHSBi3t+Q4yfblt/wuucryN53Iae9anwPLVHpsyFeVKFptIF
GC4P1k845BmUHmLiTrV2sachX6nVM4QDTTA5EmWOnS/MIV2d5DdpFUl0XLkyLvPP
509Gwdvz6bv2O/MVo+83wT51V7LZUcXB/IqZ0J5GkNmZI4CVFFs98aTpmcpRBna2
sm2GuY4t4cC9nV64LwVEhvjaQCPn7y0iDQ5hTSwyhkhQ+9nv829goECpWKCPGMca
JLxHFKWAziXo3rIqf1c7/mXfEJ3cXbxRwkJ6mUO7qL/Lc6RE1fxqKVwiA+gvKBxN
IzRLpyu4I5DNu51gtDuA1aa1YO3zE8/ev16bnkBJjAhA1vJkCvlOUu5mnRfH6x/r
WMgqkt3M8TL6bO9OXe0MFmXyf/Q6a658HJpBKBKmJo2xFy29+T3JjexsTZ+zkg95
ERKuOLV1YFqKY6Ald+mxWz1SkE2+Cu8sO2I/52sPXHqO2De/pfqzXMjwFV3dIjbO
W3x41RsbDqDnmCEwJj1zWmfqm6XcUw6pZn/ngxx50N7CWCK+LYIGcF3nezQdtIeq
9PfOiCHrHB3Fwcj+TrTca2JKqBzBH9Zs6ZAEs5IQG8oli6t3mjGyO0PkTa00aZeH
2xsA/wqyD+pe7nrOivGe7PrVhKJz0f+wM/u6p56u6USp5/Q65RnMT3fWWD2AB6ee
VVShmwPpAxdz0esZ97aJ9rhxeLpdG+Jp6PdSj0IjspfQSrSmGJ1cqMx92eEowzjh
biGB3ohEAL+FSGgRKIiVtldpWDr8gqAXV6qHeMTr5zxmqjXcZNeX4B4ZoQKMhQXn
7d2o4VX+8VZq9walBIDJO7y9oq6J07d7J4/sTjTamCZRCt3N1GJbX8YD4WCX6u9o
42Pnn2OfojaQjKYOQzW79frbM0ixTlxOR0yXMeRd4l4J+fNrKqKXQyOgOiV5dMMO
5zBtCOQnqS786d7+7E9Q2rsu8p8mOWXDsIPP2tVoZL1p4HUyX1YlqAOwFaH/2p4O
H6qX2/DBWY+FxCyS+AAz7+obF49E+ZiPnDQeb/URoMmqskf/P33Q1iRweRxuCs6w
ojJYxgR/BTUMuWfVsDGj43qiNacjlEgRNl50oL4/FjklP96+XAdAoK9sM0F3f2Qa
Z22+06SoDbv3hvVbN8ObVi6Tt1wop4uVWWagSvgwIBarj7C+QhAw0nFCHeOkjgZR
U+nkmg95XfPWQXikuuTix79SD39eWSG6CLkHYAl5Nvmh6qi7Rbzdx6PAZL5sFInv
1F31ujUsdbZU6mdvHITf6s5toIFdd1K2hnABE8Ll2tHo2IlhuEbVjTzPabQFnjV5
HNTXnv8+T3IQUbCk6W7AEcLSQhy5MvMqcxZq4Wx8t2iSW4icfjuOZMN/L7ZVXFzo
Uv77t8FoAXPCrAP2M+wfY8eUnDqzotG4Jx6vahBlf4v3UgL6yr7c3+KzGGXNU0UA
l0wWjsXnWoHdzBHnRVwrlxqn8C/RvnFp2h+oiqMh7pY91U3o10bV98BdUbQ2Nn4/
L0SIclXm4b6NJl1w5kswi/SDhlp0nbN/EfzKQBa7JWBkaeFSblIx72OZn4f3qvxj
Pw9xMeXHBcmbQKksGKFRftScbdiz56sXjWJWPNUp6beQe0pLSqJiSDTSSKj3yc8W
F5nScuR6jyZUI1sBKLr8xhZ9FDlQwHEgya2usZ6Ph/K2xiW2bxkESdvLh+tFVr46
3vJRijb8h3P4mDowa+khx4rIEQE5HYBDysfECGGupGsOVTLPQxne8EgBOG/AzK03
eDKLL69p0ZsvR3WppZsZhFaA7VXtACihvboD6hpwIQChWViOerg3vvR93V3xHETn
BKPSyIRgn03XCKtXqg8NSLxoU/+P7a8P8F1FnFenn2Lvqs0fbqUchVwgjrzQ3EVx
guPqdy48WuhcF4QVffv6c3kMKNp8m+TMGRe1O1Ez8gqCalANH+uy17wI4XapMRsA
pbiqj1YH0WWJn+UUJuGDxvXegpOMlFIGtlE/eIiu3BJwKDxyL5Z0wxdxaO5lgeJy
gOhrdc8paX2n5kmyVuBoZxji7YQ9D+dVm4rAeQtmPwMhe0yYcTy+mIkx92tAokCs
deBqLqQneVITI24gyrlXnOpfQUdUMMMEtPpcISU47DwOoQLltFfCWOVrtbbmaMkW
is2I5/fAnlt8WGA9lOb7o/bRYWNXnwZ1IUxlj2qna+5jd3RBKFGkZUR+1twfQwc9
heH+7izf/BVCaKg9ZBQdFCuWGK8c8bVjkWVLpudYXD8uy5v8V76oLAx0GiZVeFFG
/fViXuxa4uAaBD69VY27jBQY30a3pkVlKeZBrjDJAmHpIeNimxuD0XsxfKdkOOx4
UQeuLeGunDi7hI8gDnH86NRhb3XXwZtopbALtW42CqPQY9ZfeMzlpcI1k0XHqCHr
xQTgoL2OP6lAKklg+NzPjNhKKT/XMbMB+VLjqCeO777rVdGiYrb5Y289gdviDAWW
yg9b05wJL6jOkJOdwO10bm8H/DrRnEvLFk00A4yy6y5ozuiNl0fKpvszzANuARD5
ObfirM732MhlEyyJmQhB+BhPbyg2MPFYMWEcV13ww/BjIMsZGWCFUb9BtBBYyYoB
kXK9ClO7fB+EGBfMSqE1EBbZXSIJVkoAe2V17Do13RRbeIihZxs7HXFVV+Qj1USN
3501gf9Rv860ddzslZu4Q/1o++h9oeEutvzTvlYuqKAurJIAewsUiVlaitLqtaWi
rwVgQk7JOoLNMvom+x8im1Ua3375bBEphqxsnpNuOJzaxZWLAztxg5rG15vardYp
LKG+SdgurDaWfKJIbf1HCghz8GM9boARWuva/32S/rCaKG4cN8Ch508EhnQFqJbn
eZxwvq/X1hNau/Cdv6VwKJEwmW/hrx7bO9L4F7Q84YRVo0qjEa8h1uCVVjLjLVxG
WG61z8vt5zZTgZA5oA1qB/kX9QrY3KZE39mKl9tt/dROmyEOjhUMb/THTFh6nu8x
NZYN5tXNrIDb85Msf1fiubYwMEwJ47RbMn6H4oE7mC7evNO7+jbtyxRChblHCQa6
wQzjFDLC7WyCKSc9gYEchsQl7V9krqXiPPWPhNRJuvJKLUwX59DeQmbulPGJPIFR
ZIr8oOawyumriZ0JAim5nEmEBeiSwe5RxSQdVoY3fpB8aW79Mo9VgtVmc7KCpL4L
PYxjbzDQv2Z/ze1adPSZBiZQL1n1RO/yWlAsr8mqXwWm+nlk6ucMNfr70RXv8EGn
UgYn7DuF1byPul4vduV/W7Cc0b5Jr1GcDuBAhp6Fm7JKlBJ1ydc4L+42Z0/siHUo
JJD2ZlreHR8i46Sc1dipthm7SZVfZXLmsMY3QXco5wWSyYthnHTZ4OcKZLMumw0+
UxrcqAOoA86OcgXsq7ySnL9J+2SKDBOECPSZurdzEvdvNq8BS74Frr/US2QxaPqZ
VzxBQ7kkRZ3h3py6kLbUtfYqKjbr7HjH+uktdxW3bqSxVW8e2RS+UCCoXaeGN/RG
kmUXALLtxz3yo1jYnVjHTlh+2MZMCgdUexF1nhsa6wnw8sBgqpQgyngfyzV/p86u
/030dEua3FqYMObgcJCAA0rTpSykDlebK9tR2mo6dlIHEReraXGsbD8mLnAO4H0p
7Ki6w8E/f34DklcpM2gveYYWjywEGQBVlbb6ji1648ewFiYujxdyahgzF1c9oE6W
yEkSeMzhkR8DY0PM014J/HdTST7CHYuVVKuzNH6US6BYjYqF0Efd5Z1t89V/gepc
GO26r0dEtGkTfZ/OTumFTRzLBjrOFtntCy5lHTwjCmi1gFQrAolF8m8ZkR9OLoBe
V9hPZ4LkUnr22vs2RXFb1LqzH9/UcNizRKCTWQ6H6Nbnqqd8zetm5cegWNRj59Nc
2l6RISxXZIS/EEIfsQZWl62HKEadE4jp6jM+rA0qHXfevzMEikroKsZxuQriWPCN
4+5PYgVGveRbh2Az3NPWMvvJPmLBjgSif3YUgHPDu54pBpgZbndVnkE4kZRpjcUV
3xkGIKC6r3Ju1r3GDg0xKQuqgL8kXGs+x/bGCrK9o0vDcw06w4EWMiZhrxCZgN3y
wtzIF9DDoRQbgtjemzcq1l2nmxsqgSLUKPTZt2+1QCfOMh/RZoiD//tpVMS5iG7o
0IrUhS03Rz7O8VAp4TUnEB6SgeAYbfUPsOoQu/nL7DnE1qymUpSrq+tMFEW7saM1
zlk9fR6bwxhLHbPRxJ8epEZohakOGhLjWQBUId7lL9wYljEoU6XNL7HSrHeoNzyo
Nfq7lRZrB7j1LKpuGWFzYuorFZnJHJE2oPlohMeDP3TqvOdVsKN6Rby0KalFWUcR
r4uiKcuH22aBoeg4WmfwEbga6AzTIrRp3E3cXovSK79Vw6/NJht0tnTaBGUNVjOE
K2r4ZwGCLUHPlfxOTAR7hkzj9dnsoKy0bA9JuhggFRo8QoFzy2pQsBnvKvnI2ef6
01b0n9OMkIZPPKeU3gY644/GOVV11Sexv6lOX0nO0BdmE7wxuyB+edBKTMyRnNxx
TurDsME4Ec3Jz4DL3kNlbo4dxoN6mAKLDSRjQdHlgKk6vaQX59SLf1mOoGfmi5Zp
eSCbsh11h3HZOrJSnmTVgeDFG5X2UaEtwtHqqtQW+f3dV9KHtc0LQpvWdX7BwtS3
x0KDqKAr4VXegqEGkfUGIToNX/+VJBBP46zirKFpTxMFd54ftEMy5Eg1LtYcWKTJ
wSKOYSKYFlyPZnUoFiXLxFWHZVU7QYqSu9KSLfzHEl2sqtdYk9B/PGR2rpsuehu3
7QApjiK34/nhrtbQs800XiEZ3YhnMoKIVfNv4Fj4r1R89SbuDCpD9hHWdZVxDCTS
xfCgvoUtxe1xmtZ6cQAqwPj2m5PJwKwtzhdhLRYBAFbjLDyqd7YvhtEFwTaXbzI3
bmtojtTDOJewpbjTxmYnF9WLz5q1fbohssCG7P3paoBnMt/5RvvAvzU1/xrm5Dx0
wpPMOIHSZSe8N51hUYHkrlLsGfHLR7jZ6eVOEfYhQimZetYDVZOynquv0WsSbr++
azxzInmQUh5HjfojsseM8G+wZk9D993vyTxfQXsnvnoXEjT7zIuZp2XsYEa1ORxG
R/qcieqy3rGDuOqPhsyItD6EoZEaqKh9i353s5qsgkyXV35Fk6ZuPqCAFjaovpWp
2Jl6TwbTqqiVVoxwjVktOjJhWHDxJ+dN50NXkJwawKSVIjyW7/tDuB+ITUQSw+4d
ASAtXejDIZyTKFIzQMbfe1b8uipIoE0cI+z8oWWtYgd9AXlj3h5H663WFCtNjWVI
yySTBP/sfpSGqw7Sjy4KAHr9+LZeuKrz9X7H5LJtGIr11cwRdSZS83hC6NMpKh67
nLxmab0XHTFWtLE7X5w4aQ1SDc0FjhQN0FDwUWMS/i/3SI98WdHZHXsPcr+yVCip
NEOWzYveQ+8z/htnC1qKhcLbCkHw1wXGo6FkjiutDWZeok7tX+7ytYHthQ2LXJq2
YDX5tk414NusuICHj9jMVPlsRLDthG+IAwVtX6M7PodeJZZDv+vpy8kgLMACdApc
DEuLuc3w1zqUOw51XQ/jckuST68IHc5vB6Rr+483cTJQB1dFKM+ETLAsxgMyXeaU
l/uf4ZvT67iFa+DU5M4/zDv+AiasbCE2QWgWxOYGMg14aoGW4C3O8a01nqCk0joX
ILX1mRqhkwrTe2XrJ4O8Wc4CkxMhUgh5ICn/C9D9nv3FxvKDB+47uAzlQbNnDqGM
KE65lqsNJaiEZCa+c2hTMKUBZkpmugd1clWU5zi6fSHyhpY3AITncSjIHgzxgXhG
YaPk3KeP9hjIhUHPmn4FVunsyZWK6fMo+ex03Fo9lCb0TuydEQJWnqXXLYeRTXF4
z/rdn7vx+NHMYusd9/q5eml39NcsHeWQX7GC4A3CB2ONAAHXvmHlgViO9ty2BP0G
TmuK8pMcDU7rHmBk1L4h15N9JcuBb8t0vjoRh14+gqBatVy9KZYtmJZOqYE7oy4H
hIvg0KngsXT62UAjXoTvgm9G1rREPZ013U7YNF5MZs4iNuQyK6cqLi05Kyc4wsHl
LK4ENeesUPWiWMAxRsI8RSEcFS3Yrs1b/UfEmHii0q7TWrFnnIVupCGE6MXsV1Yk
qfnl9rrPm78NltyaogjApAG19Ti/6EGN/aEBqHjh9lVF9WbTBl3Uj0QShHJvzUGn
Mc9PNwnNmpi3oP/pa/IKwr+J9um6XzBbnE7PeYqIWWCmavY+JxcyMKF0/5Z0l8Bh
xwx8FV2/D7LhdteIpeY9sMJs2g4KDQas/39Tny4vM7m00F4kO8a2jj1yP83/prPM
M7wUSbuexKnzWG/fSAUV+x2Kx86euBPm39ByxYFCwGYUi1uBqBr/ORO7HNWuDv6b
qzEtJpe7U8Mq6erSR+3nAhl81V6gH3vScXuPmBDVzl3MgCZ8fmcrInXaJ/gu7aI7
RskAkI5C+XiHSQIpcxfqFuLZqudFmqMZcLDG/Yux3N48goMbU+OXjO4bmMRI5w3N
J3XyL2kDkRLUudK5JfjgTcv7PxhDP9uv4tvwavzhBvPjE47xlgXsfcz+tEiA5kmp
QmzlzHbfEUngCYQqx13GLY6xHxIu/EzxldFzBaqyaejwImnQP/Sa1MJ8/+uqdymH
8pjoLCcB7b52Wl8dpvgnSDtqRDDhmhhR9cOp3tPRXZYwbQ9WsbybquqGX3Rq0gK6
2EGmFjtxxlPqwxKWvZQPVxUupg/P5iX6XY43Xw198gedVcNQLrMzAPa+C2O1ghfM
eIecUFi/+Rk1MY0MV8A8HPGt47LPyNYCjz1f+pV9TnTsXCBva2KYptxdHUzfMSnZ
ks3YqowG3uwE4PxNT9FUjuPYFj/XYHFYN58U/zvNBo08qO21oF1imHUFiEw680/N
7mnQ6iCs9Hhlgax8M+BSmWAtCCmNijO2lf2SmcIAWNs0vV0W2whTwvHCcAzL38rQ
qAToPOE07XO8d61i9Ionyfc1kfR+ar3ulxu+TcEhoOnl/wAMDWd/t/8B5jNBLAvY
WHar7xD/9TCArRibaCwRa56k77ZoQNj++OMHMKj81arktWPmtG75SYHBaGFV/j2x
nl3pjziJGE4+cl8A4pENS+nZOChqhzy9HzppJP4O7523b7b8nHKQ4wklgkd6EL/b
JIsrWdME5/Q7i9o3gZpJ1aF+/7ZbBQBkPkHhMctmFGORuTsASAx+F/U20bhaHZAr
ZwfQwGGSiNS6bPO9+bMc2QHfJNRwnVcTz+wksy6Q+fBRaGI4Lt2lFuxgYTtX3Ib7
ojUegqP/sFesEtLly6tHF4YIxD0Ar9MNjjtbbhxM8+rzqxKjIY5TYeFgXXTDsL9Y
zr+HXo7UUiixS2i5Jjx3xfQqGAV6BbBg42NoqUsIcRqZpEwRv3QyLfdkUUYHQMK8
idcLujcv/PY8Xh68SZxcnk6hmL7/LR/uFO+bK96hr9WHA9Y05SoTzvSLhzhQLqjW
Qn5XPkI0uM9+2WHv62M4YNX0ggkIjGV4a/aPMnlFUeRYBKYxrSGEHqBlZoOGH1XR
+K4z8S37R0qndFdDpb2Qepo3VfIZm3wm31o4OEE5FsiMCaM3jjoczBqcz0QacYcU
PvFep1EzeLsZpPNz/Io8qGtAgMZ4V9JwpG5Rb1wo1BViy2ORTWDzBnKKuT6BTNsa
y296u1JrHCcfmxy6JgH499EVQXfNhYPepvTdFr9gum6mJRXu4zLKBL2Tfuw7IfGg
6mUk614coq7zypbRZQ0AYzS7a1EhqWQT3W0zY4fblgPSEUFoJ/ps/7jxMfbP7bOE
ykQ6X8ms2ebuXvRAc07XvX8hN1CfOszdz7Y/r00P5T018qJ0gvayUApVuqhjF0RV
C0s6DnItMi8EWuYZfqjoRxrQEtWDNMKll2m4I5wCMMcba1AxCHMSgce1KOEyTEDX
6vxfZsBivwBnao/j0bcM2Q66OFx2Z41FmlvRBtc8bJz9GBZb2T0p2Ld3S8cgRvih
p7JgwFEkhtEZM/xywznNcbSOY8597dBSNGP3dL2lQD+NcSgSAQq1orDyluOQ0xmX
JUjT12EiZhjELde8Nbr422ZZ/M4PQckm2OgGpAptJCT6q4fofqphYy9nzAAx1Rq8
KexJhq4xopKKxDFyWaqQNpw4asU6pvFZUx8D7RSpyT9MYS1cYIx5yPcaiCj2kwxj
U04+f4udo8xT4Ih4yIJUEPdaFZSGn8Zvi4iWCvKLrn0iWaq02iy5GaJCEuwpz2b4
hKK2bAZhQmPln/aGktN3efqPONpIp1g/ZiYAV03+WUFWQkDjC/cB/KiIxWa2sgTy
JCkwzEz2j66X7EsNF6CSDa83mplQftYEZ+8DveadvzyferYTh1fM0z7nsIbHU01H
OmEzQkGLE3UYn0jZOCMZ3tywOsFWuRtGEUX6D2TAkXwO/NOXeVkXZUwsgVXz2D6O
U/kdp0TJHYyGm2ozxqkeNpaSkR02gF9yRjIy0LSo8E7OCQbaWGm26AUWKmcIHiRe
PpEpvwIb3aWerFqqxeKyVsL+ndbqS8vKW19Zip/RSr6xc/GGPDZNdfKI0XfzNNGK
fRY6Sn36BSsec64xKBnNMemx+nkcjBl5MgrSxB8pBB9KZY160jGc+bFS5bTTVglK
PKILsOrdY4NpHHvLoXXelb2Rb6ueZBd5QAurGgJm57jU3GwUiE8p1jgxFkyk379N
JskW2Vcv3GGw83db2oo0xfT+QY8ttzgTr6GbkOUXOUzmUHerit3vKUHXUGSas9iu
1ARBzTH6RhSpzjyV5fNsCLZOZ0HVJx3RUb/ziwtRPx8HLvQ17Lz/0xumjf3lGKve
et6urB9OI6EgONSTj4S6p5EtAu20+6MkOXtVk67fToI9QaTfSdA0LMxMkOGeR2Ln
J1tYbXseY28jUbwdLnO3/eV4xkvyLFUrDNQCqQezuenC1ku3jPq6WiE1XumTv8Z2
VxhfNZ05uOyyrwZSTkmgLzysqvsRZATxUp1HUhAxu2xjmH8nAhDYfBScKBcgGF/n
cYLIG+Vm5APllHdQMdNwOZZrTeVT7WujJEj+uGhgpcJb1dnFdHwQPYTQ/9cUYc0N
CgkllYE4c/tVgv7s+s7bT1uO7F6Pafco5qfT4t2mOf0aBucfDMp9Lb8BiBH2Z6k0
bNoI5u7UvjPiXXV5J8iYCRcG7Fa2nYrh5Uq5wh+V6OG1F5XaAhl8PEErF31Av4FE
u1eGU1DT4PZ70/csi4bLIk8CzxSS9CkLd4u1BxQyiJRGyte81gWvcqJHfsjgVzxG
CSgcaaEcwS7B7J4KnHjh4EeA1JniUI48f0l0tlYg1VRhRKFfVuSwmUSLwr9g6mXW
64NkzwBtepv8BJLe9A2vRAI4/Lkn0QuW2vQTdx8npSU1pvTQtHEWyB5p+6eI2CN/
0OZG0WMxdcEQJ6uV0bS1+YA5dM3RnMoxyTOWvhvRlfcutLNHcaqAvsq45qJkrGJT
cz0POq/lsHMCG3QxgNzaP7RXxcM5BrFxqw758+Qi9zoRoa4Xx8UB1KpNd/MmiRLu
FRgNIT4dJVIlfJqo8h3q3oRsCYD3neQfcjVZ2xpiMd2pSMrOY93AfGSHjJtTl5gj
fBJvq/h9orC2mN+BMjCzllBPgpDRxfbKfMWtqnx3p1OD1gjMruvsAHeeWvosD0fI
tnNu2DQHbIy0qnzgH2/hUMkEobqKkaV3IZktpFDB5tCrvjwP5145pYyacIImjA+N
p3itWtRz6wQTq+CSNoHHbSohWGkUyjYO8Q7og37xIP2HjYrfzAE/IRgZ3Pxfa8oY
x+ysQJwnnq1IKUWsXjNglO/0EHLfinci/9hm2izw+L5eBJmajMXEDIfWhRuLoIRq
TxbEw8wFW1JawY7DC6YHhVoqw4lGPyiDiFDWLEuXQFIczm1Rmb/YaBXc6v442Hzo
yKQ/8xkOlWZkKPXeuo2yCEFSo+aNR/+YAriWkFTq4bRvVq03g1qPI0Axi/jJLXZX
PgPn+eGurZIkyBLrEciDLI1ynvWgyaplMgzUdHD/kakBEw0B4aGXCTSFtZE+znOE
iR9Tr4h3TwehJhqltspkI5WPY3sVf/NzcHNuQY/pdCkq1sCYfnm4NP1y+d876khH
iEN64xXldRLu344I2SK9QaPNXRLXaWMZFCFeKoxKXKzxfpLNrG10IBX1amwnahoF
c9bEBcJzUWU3qOS4p7UpvDPypPlS8YDkZJ0MQsZoNG7qZy8k/FWPSI+FmuJ/iFrf
OLJjdClXSYuOdndRcZ7vMlFr6NC2D2Joc8sWy6HxhcjBmFEv6ud4LYEdNknbrnz1
njEoxnHddQmbQKx3d0lR2AJiNH4WeLKsQe9O4cY2Bbh6vjcVFE4JWpQc316ts6T8
JGG66hB+X9jpyZXvvHCuBxHjD4+QTSjvLcWT7j55sOFvuqUjIPQUsAPdMSA6znBs
ANOkmFoildOMJpNb4axvCUvFxt2Rk9r/Xq7LlPmujvf7R0V5gNE+DedmHhjIXT4b
dxkw2vZ2/ejOZbyEtyXxDZDle959hs3pFihaN4vKVoS8EMyW6K2DNeNgDBFA9Vv5
+t3p2q/zTAao6KKwIArT/QfJaAwzTnelA8VTla9I2ha7AeTigS2iayKFzaRdvIt1
pzLjq9DYyu5qlw8U7Jgxr6w2lFmbnv+qGIFnoZd/8nz6oXaOtPC9ZfogkuQTWkbg
3lXOh6b7eQM+6Phk0rTGYPgEtgVRsb6m43JlUgQtPHpQsJYd6pnLenVZSnB819n7
NLmzu8fjvA4MHGyltFf++SBjlWb0JImHYH8LqiX1wVdkFCZ3cKw7xgW3OfRAYiYA
8fkFusCYyYuGJHvIL5LMwFJ53WZiwn8jIRQ8F44dDS/KlY46f7g/FdcncPwJVHFq
wgv/fO5EjyIsO7vgkIRGco6s+b5Q328OXLYYU35l2+N3js31erGVohszK7N0DHhB
PJqHbxDWX51fUf2nuK7FuFhRtgi7gZgFhH1FnCt4v6KRAode2iVWZ+QTxS0+EZeE
I5vop9L0DCiIF3q6SvMrJzQ4vYJKSxZ9VoELc+G0QvPuwfZE56CCvwVGicgdX3Bw
YLzsirg/6AsDt9aLRV2W9AVDy/o2lSd5A2VW3jff2B8U39wu38Z/W07eEJc6MfQK
n7Xg7siV1RjFa+mm5RAE/TcpU18B7p01e9vOCYj0grLZr3DHyi8dPS1IA4vFxJ82
DaxMAYlp7kyzbGW+47jtlhWtkhnrLY6x7uZ9WAEqotC4Jxp04ShpzTclSz95xXR5
iueSEe04KQwt1Liyh2yVj8ImzlcqkmviPpPwYpaIK6TzXyosEQ5HzQNOsnhWeiLo
XqxzhdSCwHqRQwYC4VqvlIVPARGCL6DfzWZUi2+sR7YAoPXq3t8R335FCy04gWGu
gX91ABcjVkg5OsyzSQ+1S4u2fGiE+2cOf9EfknboHlvwFyfRB9jpWnIWG97pgyse
a8p849Ll+PcQx21cJI/gz9ZbpeH+XApdNmFfxVjsPdLoNFXUMaTZjWos1FK3I2c9
5ogsW39iUfZsXiiIcSQYy13kgG+ZMi+pIloF8YZPDV724e689UqKEp1oJr3Js1Gk
LVcJpWO/Ht2A4HBFSrFAwC+CPR1Brkk3mh0gDP8oAQgQDPeXjxwFD4b1buz8V3oB
TLM0esSh8pQAfGw3N9j/melY58VxbFQVtMlF3FOmN4hWDaDeRMec1NGA0DNGfrXw
KHWRPWjAl4VEKD8ymghLpw4VKvyqPzFWk85KoCsLpnn+ZicSQKuWOv8TK0XyOsV3
+Lx979C+/XOWgOqruyDhrM4bmLjFlnaW3D9lGKdWFI8yLR+oouNhrxwCXq+2Oj4k
9ifPN2YvLOgn2I4ubCUKayaJ/5mBWbidNROgOoAxq68OROm5sQunjwvunLOCDSZ+
xcIR13zHw4TEdUqY2bedL1p5hrKFDY2icqdCSvpdL/fwekes4xOhjKhaLVw78c+u
gx3Pk4Y0uENE63R2qyF5mQMJGPDF5DBEQnu5Ls0QRxDZo7kAyE0Phmt9xIeGIO9q
BgOvdLz+SHSkqK1HSiBNSM3BGJr9vuqWZhH97XU0a9EYteel5eDLTLTLxazGjaQ/
rm40YXiGSSmldMqfReuCESN+SAaWyR5sZvXCYdC1f0K9dfKHNfjYhpnJJQ52ojhS
IsvDrQUsffU4xspUgrhAYGUmCo3N4/GoJH9PubtPMW9K00zz/Tz94SZNSwnKetAN
Vuj7nijDFBCCArEjTyU2EsUnfgTuLahq1zm6jw0GoFjckLHg+Rlailnp3GaGlgcO
OwByw9Mw8VrKR69MqGzgJUr4nkUdPm5L9WfDDetMHJfGX50Wspl+PJVfAOD4XpO+
evbgyMXaRqOpD/SgFSWxbAA0FBjrUOqsRooQURRS4PZMo+J3jK1WXH87EYIlXNXg
86iF261ssD5hSABS8rlFbu2GqXzPR0ME1eu9eW7t8s/+H4l4j9eselahRrIoOvvl
3OKbvNT9GB2p6wwdhBPGzPV22X6smCfNsYIzOXL335R6En0rF35fT1okmWONCpUh
R0jO/eRPL3i997p/rK4bDoFV3iwIaSrqOd+6qJS89NGbHYyW1ICwjK9vQLQ0kxhk
LKo5Cvup15K2rrSOnt9/5+4RbNzTG74UA+GKelaJTJSc2V/jdOqsz23kYhTN4nl/
nVgLH698QevXBxh1z7GdzYw5znemDpwafldC1wZ5XbWiDszq0yLrZrNAvOmjg7tA
4O7dG3Sc06QKUbAltozyTTB/u5m1JEJFCYHwJ6UKty6KMdA9dbJSzbmhAxYASArW
9x6+NODlanoyOibTm8AttuZcEgioLpwVzBXcGzIWTWTD/r213Dy5KtmfD3mq1eNi
qzZeTrGK+V5RHyzvwRv1ixo2IKO8GLqQhxZxxlQ3P+f+vkcaSAvYa843ly1DFVtQ
SDvIdhaG68VwVvMU7kZva1KwCg31WxnWWQ9Vb7AApQW8GJAGdiyZdxFp01sgeTrs
3RatQBWg5EgSXTxRGv3LHgVCdJ+kMYGwl7F9YwQLf/4LNPjfIm9VVey4qQhsE+4s
5Kfd1u0Vqpja4OXNfCs4+Fr9ul7FpWLOOzrvl8NRkOUsrgcFumlQvmHbCTKYW4rk
mCsB8RZDhCgrYpjjcUB2un2rGfZLH/3qHfdGw3261+xGGFX9K9NQi5ZT66ODU/yF
/SUI9VuLG/jD6r4kWAHeihWfFbNPqDr3qvEtOrj0nTijBQU4lC/ERZIMkK2Uq3pS
295lOZLMx0Fok9x0XtdtvnzS9pp18FNbD2wChLGe594fZUld94XR842Zp+he3hIR
GT+/CTMubd+/FOAlSLPB2J4EI0nQbeDUydr0GwgrOsGbh9QK41EFkZzV3S56C5zK
8SN9Y3U5KR2UEb0SWDJIuE+OyxRXqMRhjfgu+f3pblaeICdZEiblIt6ONo10bJo4
D1LUDZZl8ziMNcBeytkGKvmgKKP0DSBTDjEQc3fATDEm0Y2zNZ5rRDHipTURaOVk
qxLEMp/2NXJWA5S/udedb5EEQBxk51RoSgck+L03U7xBoIUzcePMc+uYiZE/BnWu
p/irSUCcJbVbUwqkBjkoH89a/o1/VeUGvCkQM319qGDicWnN30NIkEvHM+R0afw9
F0QzNW7WTA6YeTlDCuBPj9uFVkC3/AFTXiR/hA16tM56YLtQ3OzCZqL9/AjXcVlZ
Czupb1Na0Dj8plSCM4ReiwjsYfOv1HCQuxTrAGHiWx9knXaYd190tIHM+jN2sq/b
riJE2iFpODrdRf4K5xjWEi7sfT5uvDx4sNk7Q3jNCaCvcFClY7wdn2fmml431HJ1
B1x1A8SYKFaKpZCiCfqmNX8stjiezqMTRgIyKxBcE3mLF0PWKEfaSLNYGUuTC5f0
IuasNbbTGXZLLfGCnqK03lR5kqfMpeaLLmPg4bvvdWNjOtNeXhmvvPP7lkK3a1t4
O/fJmDVUbK6+uxImjnH8JdzzxARhTRVDybq/LAI40g4c1q5nIosQYn0l8N5Yz4Ms
btyxxkwJz6oAo6oEJCCxA5dAKPthQ1nVaN1PmxEUOJG0AjtWaL5CNSOrQFvIqPX7
dk3GDpRpe80YDRcvh+4ngi3ag1VrDCcz929r/j72ACWDGtOwmzEhyms2qL6xdnKI
rHogAqLNyBosBV2fKpU0InDM1PWHfHzegvvticwC1lsm9zQKZ8kJy2wiblbTBeO+
HINQWa5bYTjO4xMVPx7TCVBxcM20lEFBB/ZLISjIiXOozZ3iJ8ACSBHutSvT25bw
vqicY01SqVe/lmrhJU4XkhzHynWvZSLWBnvmsywgaXLfXuvSIa7jG+kGv4cy2Lwv
YkH8f088tiTx9AtkD7vVwqPzCQrjrolQfIJgIMvtOlc0NlaO2JeMSDQ4Z6WpOANG
EF0B7WJP1vNm6ztI2QAqBds1BvSRY3QQvm8pEoJwRpRNrttT4d551CiS8ndRCmAr
Bccc5Uc8YxRu1okQbPCldVC3/BrUiZIqOnfFLiWOhqoR7GDzyUqHrhx1aQ3KpYtx
gGWr8sS+XRhtTsbiHt3Rdz+LZoz6GSiRdqnbwKBBiODKDCq9WeknoH4kRSLe0auB
tjm6s88Ss3HM+qHiHxRxzhnGtSlsqJ80LUhFGJUZTUhRg3E65iGjH2q7tMVdyN8D
pHIrX9nuTmLEutZYXjcu5p4AanTwLh6Vjb2tlOk7KM41lJ3zggAfFTRh3H+s5Q74
L96GTG1BvtizF/yjFjtVr5Qkc8rejg8XmLTlrl83z8/1LqFtW5RfPbTrGyjcDM8w
/k2vulMNsqBWKeCKHBb6NKyRlyxt4duCTg2fz9IXtl9TIBNtQzhUjYv222+gEgZq
4znHfJuyDExHQ6AZSm+YWWKBXp0Aw+MYir5fcXUi66Q77Gt9mhaojs05f/SlmXx3
pbbO89AWS55/+lnc9K2hPd7WSuzkTkdqZLgslVdStFEM/A81jg/g6y0NJj34Wgsz
Ygy0MI4XmlVbfui2RcrW+rAF5VKJh1DxpgGXGkzsKKkWflIwJ1ehNgyZ2xYr6n9/
78qzuZGYJjaRDNpO54irbe0XkDf6yqRW9uVvqN5AJoeUw7NuJKeghTNZKNwG+iK+
m771u4Aoq8ldgr7cKWp5SmcNkkT24gDskvZBXpjr/nX0zUfmr03+y3rhmajDkblA
7XhYe4XLDgc9R+W3/DRWvsZv5szhVxol78uWf3mH3SKFwMgU8bCalf7esOwVkcDt
FlNwEwrESjDwxeo5MC/89xolVUq36+J6Tacf4J100CbDwhZ+PPDgA54JTivlWz0u
SIDekYkmF0scm32KlkCoWHoPBt/UCOm8X6p3DpeY3NcPfv0qPWsYu8XBwiYm4tGR
yPg9sp3btp1OsCDL3739E8cJvOPT+UOtZtBirNbtoQSQbSFdBK7Syok34e0ciYE6
mdYJcnUHitv6+DoEDgX/f4cnOiXstH4rBDWmk4k+yDZdSHzCMvliQDKetfgujEvX
+3VeNL/ArixRvSjTCUPn1Xh4nOA8cVHzotg9OS4PYvYLfbyRn3oxRBRjBh204JiU
9MCk4qhheZkee0REP95U1SoQJW3NjEGBeUfVI7xCWNPekFfe0N7xPQj5fwx4HJfl
WI8fD2aYPkD3xnm3AmN6CnxhvdoHd++xbsVLZgHHR17GYu/XqPQ8Fpl6/vo/4/Hc
Idf/5qOaX6IvhHbeEsZCTJUpuRHNJotBgh3+V8SBZ8V8aPoHEAQuCrxPhuhTLTp+
0hpjRyPaOSCdbrgAJsB8rUsbEk1AppAMQUpfy9MR7lsdnHpzRAHRdbQSwcc3vtti
pCuoUEIuzjpGTPlHEd63IL3GU4aGaTvezqNbtiJXEH49q/Khm6lwZY4no3aP50/7
63Frllu10suJjNdk82Qx7ZJT2WhJul4Cqk8o/PWL/o/43zqwNgzgMTRO+SDY9mOh
c8WTlslt1/TQ3eW4kYUL91bdsbmJKQ2y11veE5xRNn4Gl/8FLG0g0z0VWWcYZmsS
6XkJWiCfnY+CTW88dDN8uyHGoYtOsBZ9i32lJgXimTLi6F1gfxG07XM6YEZu6icu
ARNPWaKiOoX9edhzsfzQoky9fIPjB6Uh1ZYrYfA2UV0sRFNyGWifjJ0CjtftDcgM
PogI2j7IkYgbpux9OJkvoP/CYj/s1CrzzfHlMrpGGuDk2zmXlfI2Kwm22mLaMUJV
dtyUkjoYFlAl5Y1RnnAqVyaJmuYTUHIz53q3zSRaKM3FXaUsJEmBxxTFmT1+w7BY
JgQQC5Y/zSq9Kcv/qwZgah/CJtRDiRhdHY1ED4Xq6TkPsZNFcrT5HdusXecgb70j
W/9b/guzcik3lhxyBYgvB1xKftVSYvkmpYqiSzCk4ALkk0EynH6J/us6V0QsD5Ak
EmuVcQGO6IbhAUDvZebFLGUO9a+vlt8zcVen08fOgj5D7scV4pp7ToZarX48fs1H
qn/hryXcEGS6eDo45oBA5SZsDpacQwzXNDzkAd+7LEYjkKU++gKpzpO2CnudobW1
lag+7sq++ZglfBlTpx0Y0q4mpMZoGvFNy+l25VbkvGiQcE6mclp9cTlAR/477o71
Qagb0Vu3CpRSw3upxtotSvnucjMdXl/yJeSfic1MpnedaxTF5QFRPXDn+IIrWWjq
bCc/IeAaZFVkjBIHdZ7B0oPaNIK49A08Ld8IG4/l3N7B/eG3wTTB11eFjPu+L3jn
8tKnEW6sn4HuR/I15YmmlsjHKqSQprVUHAe4EpH76JzReNX3vhkb+ILa4hzZ8ifk
4vDgu8NQ+Bhj+dcH18aoLCRlWaksm8svUW3G1FAs55lF9QlaOSs+amWSMRfe0ozV
QJ87oIPM2dbBi5EU7y0qdn2aYsjBfbYF1i+Rj6z+6jsxotLMoGCrFIwNWK7I0cqz
4Brbzv2z8NtG5vw0oKGkChLb7LnLNsaTyjV7y4619YXz56fU6Y/VuL2n56Wf9hLp
RWkaezWaje3G7edLoqkFMqUx4SqBmPxQhJINHq6IEbHcpsm3KcAHVp+pkS5e1JGG
sFebJ09k5BcvEGVUEhdteUfwMJ2qS22H7fF8f1DpVcT+mF73aHs95FVHzrwmpntY
7YDH/Sagkmt3EJc4+on4USH1lmAYNEOXKiFib2nLYzy58zS6HymzxJkLTeNlONZr
/XFT/NMcak5Rqyqkhvgr+sfA7LMLIy8EFChuDSdzF0LOE8NAvfyAcC6hgODqYTRs
yr+nX9ghfbciIWmxhkKr1jkzgxg+DXm3HvXGfmbdBu+1YEZl43dU4+oWbCznelCr
3RdsmmEiZG7SWO4AjmlKjvA7YAFMQda+XPwS5aZVhtZaFnFeksHynfF8++oOwA7t
Y8LMYhfMgkXAWWIhsBKKtB/TuEWjIOO44h+dVgGrKqN1v8dp9srTDDoS5XDaVgYh
5Mg/2I6ajrRFbPkBoXRVxXHblfU64GwgaiyYwG3U4NWw7UKOiPY/F1RfLPhOAkal
IfZW2e9KC9L65l5IEwwSDfyRvitnQa64vRXutExNhNCEE/h4a4XjnaR22bUmKxd4
GRJvFLz+msr0mjCBd2e9XvYpPPRwB2EpvFj+SW//+hume8m38Bv7HZzvFI2oRNUj
45pM6rCAd7ZcARWOjm3O+7Wv6qS4feJV8BJkIW326008Hqltu+pOged504XJwftv
CLxqtz2nIE/26+ebJ9MnKxpDddV9EyeBsBvezBXkA4FtnpEO/sRZMNjgzNTrwKCg
0vjXE/RSX+Zhmylk8yhHNPW9xdljoVba+ILSqPRTEFGlWKhiYJx7mpp4VdwsQAUO
WhUrd1/EmB1rfEucIGmaVUDwZJyyo3JrtwNNfNgKRicyL/6/7ALDia2TRF7AqJqJ
/oiXqx9V5S4FScDx6SV9J576XZIxX3Em1LTaUa9JcoSwSJJhPVCRXKZXOr9AuZfr
zrrAkZFrCV/GSv+I/rckBG5d6qBHHC7tTnDIIcjwK74EyQ9hOSpsT6lT33zoNzNb
ahVIXhP2P8GbSd9DeEPwZEua2aESXXimfSjLxE87DNsRh8nqggw668t32NoI1SJr
gEVmeheri/ZoMe8N+WuRZFuEFk5kem3014RZXDqGC8VlqY/aU7ZLszK9CA0eWrr9
w3YRajAxuhGFffwblV+EVfGskWwutqBUsrwxvMuCmxrwzhxNZt4oGuZcmUfh7kRA
bTFoR3bdaZImdZ8KNDticnNNkQyipoesVLuFKSqGpGPoJIJHeXB9oIw1Ia3RyaPm
/0NqnbLpITueoddr+qU04Tmv+p6PjmDEu2HDOqi65V5NFAJxGCXKXSojkK/OxuQ+
beqSKJdenC0axcVUZ4QdGXoYNaUIGKKf01GYSLKQ0j58Rg+nR/qAO7sOEnH6oeY6
rbKiaO0albjzlZeaaHQMKUmGQmB8baBnFKyizd9IoBF355m6XgYNPNttAwuD03P9
AKD5w7W4wierEfvioI47ijztYB6ARvXrKYohUT0zaooGWrHBCVz0ZwkZ+fLxHiNf
4+rG2iV+yLepM6zoBrD1oF9Yklhe+ncdWVSN/ZGKUkW9eoXM5czBf5QyuB/UKH3W
E3y7jY3l8csz0IBLBfyXIpTG8T+Hds1ZV3y9/9fRlxQSphdkgZKda+4NWjvKpJ0v
cVwjNl49pgcLoBVsALQFZy3jsIeZrkKPJXWNX1ioAPPFAdBmqGCyZtRcg5n5KBxc
0P1huhUunNRKFBZt62bDzB2pgnNjfewwc1tZ/H0XcJrZwr8dq1tcPHleSSJIEjvF
5KdT2Uf/gqODZnSSdGO8x14+WPfA0ahHoi4EWCfFKWabeRvVy1dDsVkEcn4/eUsQ
AlUNJmRj4ANAdBO8RUnsFasY+gpsqGc4YqodCBQX17y4GYseDvIXeOPtJbWYFt88
XTWqTjoueuIG1dP7Yiu0WO55VJZDiumeXKbZU5cRlWmICurfGcsBCqYz0tr8bkbQ
N6Dbbsuj6NJar6RMZ4pLcS6CztZIccPeK7aTxLvEyrCb9LnkDEVuScExc/7MPpe1
u5+8AIHi5xvP5zffe0WJIC8GlaVgwUG4b/XzrUj8Irvz+ZrqIQp4UqKlyDM31LNW
KcvBvyJ2Kw/olhoPq4V6wjCfeQa4MuJRlF2+GY/4VGITaHcv1i+el3xOXqosxFXt
c2EZ1QRWLKNyzXrTG46+U3npgF80PnYzCu23vF1x6n2KwL8EffunL14PSF4FxISG
z99X6TGCIOvHD02DCHsiRZL2+W6ItbZUK+NL39OtfhycrG+5ts7PS1JMolPnInJS
N/4+cjzjGYYrTeGmZe/+FaM9ppG6e29H0LU+2irRv/jORWDw3Q9aVp7vPeRQGyry
+fdTMHhYkAfSQhRGjJM05uG6co+mQp3cIrSw4+p5YxAdRl7dWB4/EKL0rYe2n3IH
Imza2yNnM4/IvJbhYjzb9KVl9MV2eNdeZ7maXgN/3QfKOUM49q8Oo30EQ6HcylFe
Qo/zJAY5Cs2oz1x5aalMDO3StBiW+0srCC0vniBMi0KPMPxhK9bQQJ/195MSedzF
tfnsHsT0mCWHnGB0fOqbcEnujGLwk9R1iTs8+zdgQULheIFSxsTd74LyV+JVXulW
9WtpA9gdDXNGA+LjGAZq3UwA9bMSjoSF0Y+92aFw8C+WmFbGs49s46jJBuJG8sN5
XOw0QSV7iF2P1dgAgjONK7o2zmhdKQ4Fvc4g6aux78xebgGjP6OTEKE5LSZES53i
ubqTekAjL0BRsd5ROxTgDlaSHLyzLLrWzKUdf/u+x4tH5YNOajrM75tXuwWLWN2C
Sp+H2dL/pOqzmo3qU9K23acLU63CjzrtH+v61YTiIRXBbH6qc5Uc8BOrY79Ppr9+
u09RHPu0tg2dLVwUr19x9Ca0A2OCnmSVaqafOk7xSTCekPIVHXJvJQK51LYYERqE
9Yoey/j53yjQ/izNCHfeky7g8XnOYw/Z60jN7+cTGJNmvVbKcxWPDvNfU8aXUD/o
uNaRIThnSqWQh6dA2niconpFA4Ia/f9gU9XIuXMQUvNXKKvcTZ8Wpn3AopRyZLaU
xwKTFgXjK8t01fQ3WafDd4Pn+ScLtwLQYJKhB6/u8AZ1pk3MFMlp5ZCLrz98dY/p
r8Fb510FQ340d5La8ArXUoIXIL7AgcOdZXT0g0IlnFk99tOjnVDEnMBjzO0vJUgN
+2KYEw2tCrSLOqF9iYm0kIevUUuk1xHKHllzi9JxH9nrdzLmDbc7w3gQfv5Fs9yu
vT8NyBKfBj3mogkf2rMNHPiYNNekLn+dlx1rRUvabxZj9GPbrvVFS2y83F+idEjY
9hOdPB1dWqeAfld8pTexfWYZcKEakUiCUQ3qF9XxkbCEI1DP93Qa2kFIQ094hbTk
x/C+72mP7/kefSC9H3S93pWqc75w9XN6CO8deY4MIoLEp9AYHutyc9txdpERHsoI
30Q7JgdWmU0lWsjLKV3dQuhufR73dw81ha71VeEwQJcx6F/y5y3xJ1Acbkm6uNKO
eekXQI1IYrxd7UZ8bbFPUiYCrJ8+G6hcrEx6F8DmZDCib4DyCMZ8/T4qwh0z8qmW
UHelV4fh1uHlDquvMAYmhJPJlpF7plgHzwRJ9Foyvu6qrWwyyMun9VsWRq/DPmTY
9WtYjrZQq5V3SHmvPZNQi3Sml1qdgxBhQgOZafIpzE7hvk9C9BCPMwIksXTkZHAG
B+eiAR1Q5xNxZI2XXN+yH4vLZxeLJPm2AShIfExk/PP+Hrq/47EzRKQam28sh8cN
NfbQKPkPPJT0MUguzlR0nRgTvXypUDQ4feaMvaCYMDfFlwdlOYjX+59S0jQ2l7io
FRNYdpb7fZetD0iWidyYRAwJQnodXENxq+WnPxYrsC72+gmNoBqjCMd4fSJMltC0
RA6YfuomkSBMsKQaURVCwMstC1nwE6/1CxLIxMegvsa8zdw1TXbbVU6pTNDn2AI0
hdPyiU1EfcBmliedUdtpaXT+2NeQWckVOhwY/ccYstK6etytHbb/l6QKyWS7TeOR
5jnp1+ESiuzE5U3NICKWeAY+Ds1a8vPpjYUoriZTwtcp8gOw9owXbNXSVnbTPBDK
GVuDIdeq8leCGyrg9m9EqIUuQEqdro0mapY5GhIkCX4DQAhMgAHiCDM+sr4GdA0W
cPi//RUlPxRSF21N7kpuuSOVnuPD/akFD7jrDs0m2BV0RS+Nvt7NxMkP8dJ8qHgS
5qdYj/0rmW1d6lY2WQV62UzFEav4+8A6Ue6j+RHBpx7VEeiXc2F8WDkIDjDFeEOb
YfYyPP/rnCVynUiDv659TwvfXJwh/VXRfBfluCfdGA9l9xFutwBM12APvhKqWgMa
Bbx8lYJAHIK87ax0OI9B0Cn22hdT1LwuhrVIMcj+55y5gUAcptRCRtZtD5Ft1S4W
VWNkkfrR8gzA/uC6yx0vc31k9Mz3hVjdjKCg/tKCLav/nlSJW71xgASrwsarkqUV
QK7Rl/tbrIqEOUZd9RyqeKTOWMfJEAThIiZPcVqNoB9rsIUAZYEGM4jkHrxQZKoh
XVtOCBwoXSwyVNobn7Sh5is/hGEzClfRPH1jsYlZiZ/ENWo+WTffI/6l2NfONNsI
Ps0jYUjzTsbASOkXKQDwA9XZrv5TTpP9PI8ZfVEL4i/pZi6J7eMqRiwIPUWdshdD
7+f6iQVzH/CWwR3PGhdsux6PkNcPixQZUNuDeMukpay+ywXEZie3KXxOkyI/CaQx
8uDoiAkJtOrvnOgXQGDfItq9tkMeheLacCpuZloF1wHLeRIO0K3nyecPxnsUtSy1
I0xLMt1Xm5ZzDUWji4J3UJO2usF+d3sYncfjsCRANM3nGVMuyA8Mwuns69jzSQ7K
UZUMQpKBafxbnimY1vaYXGlpqYyfaALBaOh4VSrPKQtc8V/PIfpqBZpjkc644Jmf
pzM4yroKCJj/BtgJvOhVoWsC4mFhuoe2GBzYD1glR9V2BMze/cPTp8cCao2oDa5O
0IQIDsnZt9egoGxUTzQdFcv31dJqMWdtx05yb0/hdEBVeoPtqL4VglV65XJeaTde
NKwedZjeaOHcKtukm6kp6W7Snv7gZOHFkcq1gIsJ94ZHac4vngoza0ip62Pj+hkk
4uNZtZ2gC/XmPV+5RuLbS0IqZfinoqw1hx+1Kf3Nj3zOW/zn4+YFfcIG3exrfXS1
Vuy09RUZglqdDjt8zu0AkmSJ9Y2xHvQ+zR/LE4qfMc0Ofh4FcCE7FETyqVa7U2R7
viWi9OlAhcZqcsTe8NQsUGGOMb96TikOxcKCjxcGr6EteYGNlkpXD602PQ3MCcT1
rGa4I587YfkrvDJ1NfUKjYatrTayWIcWZNulofMk6Aj7T6dWTZ4pJALPZFfQjAVL
Vhqizy0tGD1XPi3foGMiE+5VhWtFJu5UWLMxIhju9m4m7edNi8jFslZsgLQwORWH
48tiHp1HcRmEocP/grxWoHBNq4IfMM10ONETgpeKO4g8W03Wr08cYQfV0xrNXo7M
OB49/cWiW+kGfVH6G6pzn/SdXAtjUw3OaXe33tDSFoSHyCC7dndUSv7nSxPZnHmX
QEY5pprX5SaTj4WLHveASjvWGhESwC3ygfo0hk2iGjdVt7lyqc/omtlejZ3keQaI
b3W2pOxR3loxsPf/Ni2/MfAHZmePnGjzmX07HUhHsFSZ86kLLPjk6OSPsjTvAV7q
vmNeMfoRXn8NDYE5OCRLg+rBm72cf53KQAmMrHvd6cMXSDoouIe9VzzhfSB4BAxz
fO1QIc5TEwxdLb5cHDfDCxubkWrwmJb7YZ0aK/e9k2gh0ZI9RZXxH0dciqiIym4d
SOujgKtD0ZNzUAjz0G3cnRHVKMHsFnJsmL+reM0QVCjCXJKHC8atgTz+QdpOPTPK
4OjNheFDEq+NuJd3JpZYlCi8eJEvYsnqSI97gtgnp/BEK+N6jdypsxPfVrrFxS5a
Vgd2gl0NpwK7t+ioiCQFpjvUh1NHfGCeyS1YAH52nt+dizXLSC1KNYCACPp8hXmj
Hg1xqkd/wArN0X31hyZ1kv1FEmhEJ0kTiicBdF0fxDuNhsFIXxDCxwaguIp2yBnt
0y8fy5frClAo9weE+ynZgYMeZvbnmRfJ5q6I0nlhxi3DazvLj+Sfe8MQqE5OsNcq
YFHzsjEFIg02bmvWGks92TYXBTjJqihHRXdmRlehloF/rgk9tywRlliqpwtMRlWS
nF8cNkhHVCTnA9p6qd1U/or+D2wWzOFtwSQM/U5AAPDc08e3Em3J94advkHfEPy9
r6LpxbH5cjA8s4F+bhdamrV+HMnz8w5MgfaWtKvyz+1I7QznCZqUDApEomLbs1Dv
e9SNhnCGn0JmoTqN8OZ42ANmpNvxwil/TgY9lugaymdlzVrjg0lAKRyoVc20aubJ
sAwMxzfG4XAGeBLVz7o8RpXgBWzR4yGb9kLK8bqKu+5eHHYWV+oTsjWUGVDAvB/G
U2b5xwin+ZguB9kgL3BI2zMjrfFo0Mybj9YFo1pwCe9BQaX6DSWjbdiDSr1abkSn
2J08n87AuQ1YJFsTYKB68/t1ZTXdJ0WmNdW6I10msk+brCMa9QYbwd1oKEzr6m+h
YY2fAK0kDBtgYAa4s9gaVifIvGawDceUCx1wQiS5zsZJPKEVaVDUAU8oSLj5UWp4
3AfJoP0UYZkDB6gFiWmyxs2Tt+yR85J2NjlFuZGzIoz59Qw6H3fb/W/1rWTep1N0
LzTsoJHCkDq9gGryCoM1Uy6HILYRiDC3nC0InsYSVtSzdBKQgPulwXoH49RZcxPK
3eP/VzcJNldnXlfXHCvFo7rFXgJ9hWytZ0Uzk1B0f+mF5w++So2JwBSDixxedKm8
PhLCNpZ7cjSwLvBDkRI0WTuEalukj9uJWNMfKiV/gSp0zweCsjvr6C6JMEDtOBxv
e1xklkZtXMLJH85viKGyAlbMeQFxG5ZuwBzFxgyj9F6ZFXQt3EzcQTEXS+r9q0oE
fjD3+GIzwFYF9JV8f74UpnYqdq4u5T+L0IM1+OW9gy8iQH2DmStRX3NdOtejDyrf
ronTf5e2d/YzX0loJz1OdFfzbtkotEDeSBH5+I/f8yww/kFOJ1bsr41lPanvrM49
+/+WptGdYHKkVJQIPd6HSaoVaT2bUy74j20uQffV8Kw+wDoQAOnSb2FOQKTGlzux
MQ3EmeGIqZ9Ku1ue7KjPth/IrCkTefZNKvG9GrVLeznHYjxXBkDdsZ8d+9Nt+f5E
N8iw/ivxCOgvksBBkMej9CwSkOr1j2zDs/ZRBVZoTF0tYpeNtwrEfPSSEjDbGAzg
08QtemCK2blbnF1ztxTl+vCbgZtlTlPQsem/Rt8lhcNJNcX5S+LW5F4S5ahllc+Z
dBB4bB8eBAr5sfrmps54aK2PNXv6SG8kVSorTq8/uERcPniDrGyuL0RNUN8Uzj0Y
YpCLeSIltfr8wYxITs/K0/cJTp/uvn9UzG6vIjxTIYybK+H86oMzzBc+1OHGRHSr
EwVbgZfuHIGh43hENtZFJ2tGINRZxm/HTJPgNYuHd4y5HJZEWzNuncydykxEFmok
JwjE78n+u0x+d2+ZdvvHQQi0JkRjoQXfQzGn6tPeIajt2VRciNNgJDZkETmKi7Dr
gPUXxdXUr62ztLcvfqU3VzkbXgCJKubKWtq/4c9eynCeYmXuo1pI5KtAMPymqIK6
GDOUrm3n1f212h+KV8METQCJNQ4iIH9MfLeQP6ixef0kXs6i+HynFjHDM3eqwR4V
vxEzwMZI17Sky7i7fWIMDT8LOjYDuejzPKTE5DRRmlTfRZ1kE1/AEbfV3hMkblb4
VB9MmJ4Dj0z8AZtXB267r/71/68eJAG/ut5WRQe1Fo7wgdPlKmnt3FSvvD7ivvu8
sSf6GkmSZVR9H/RKR6ebYr+2uMD5RUXefDSPpPCesWDGj1vryOPVUPzAgbt6HWqT
KQ7oYVOl0fnVQcUtvv2oQgNZTNgH39xboKUWp8xhFyW+f+a6ezgHChYAK3RrF4Rh
rFqso6AWV8+2qz3Z+vEONRgrrahByDat5PSnT/JR1pcHpgI9k4XeXR7PEeE0cYEb
XrCnQAURHapouF9weAEQ8R0kNQHJ7M+VFIJUvgXisY2e/OVOWneRInkZhkYjoNFB
jzLAwt1HqFDDO6xiHcJ3fQK3BmgU7LEmne+w+2Cjo/Pmd2V2agbubYtuZMhsB3te
QbH7PmRQROiLtg5lggLbBnxDw/iKWEMLMGniyAdR5yCoXQ1ldXKPUZU7EwmiPOW3
FuqkrervcdXnelBMLbe06+kL8uwYzKGC0b9b+gGlhNGTBM/0Hxy3j14aaK4ZBxY0
g5LymXzUJPZvTCG22Y88WHc7zzps5nS5kQCFx6/XrSPg2Ge0frLUjLxlI04Bo//l
VujYqaPqMgRh4W5qP+pjkmnIqjx1O//ZkdJs0M5lkJ0KpVlditBAXBejuxvjdQDl
6RKi24bDavcX8CZbfxUR9pIrjJ7QMMc0imVXnj6sK5wGdHmWpq12j6sbBm7Sx7Kk
hIxq1uFHBVHt+wCy5cEGgna388NtilUauhOPYEyo/0MqaA6Q7o8SP4TSgpNWkjFt
17m9e47M4PXSlFfRFkNO10rwYDFOlo9Cwp1PaHrCHsnVoWpbvyfw1xATELdYNm09
vgLIGMo+Jqf+a89p2NGXySPK3p8zvovCQ9WYkoXWtApApKGIDFjJ3S0MtRlFJR+G
n7LKsHp1YUCK2EGLRLRPhSffAsY0iP5S6q3utHl/1vJD/Hrhqbrl2fU2Aky1uPwp
4y9CT75p02Y9hRxUvjuV13zYe1lYUBEW7LHf7StZQcmUCUJ82Z7F7G3GzWxjvCTu
GeQ+Ag4g9CSDDB/q4lbUcoldr7Niso+pZ+1oTb3g30QIoc0u4AtOsSUXLGhQhYxN
rqSz1341a9jFcMbinBSK3pgtbguQnzkIMbAhLlFXiSMV5FxVtFo8E3i+1/QXG7gJ
ZtvSxEbcaunOwBNvg4UsJcZ8MPaoDeoC68lvL4vjj+XuzcR89Y7jsVd3eyHgrC/O
eoxbASNf/K1yA1R9zeDjrNZ06iversq6hGJXjiMRw1D9sjtnijd9yobUkHiPaRsO
9MGHUq4WQ/51OcC2TFQFOo1AG9hFnY0RjDbO9sroqGz3BLerrAl+dVmDtRdiON8e
/2VwUYAnOOnmQtt+su47XyqKi3PDbSbJsmcXMuuvLU2W2bko0LQ3CNZc3uFkksKe
WZpqIP0+y/evpBgS0tmSx3HlRBS1p9O9qq+7wsMj2zvLALzKrK5yvUuS8Vz/5O2P
j5AuboRsMCj3xa5+9JUP/NiwSZo6Cfh29ftsuIKFGmEt8EnBK7ldG7SsU+GzJHJl
WIacxeZe/yVUVKMMFGutklt7/DeKitHZ4wgMWdoIsYm2s3H6nfwGBmbarUBKei5S
/PMG2XKtuK1p0+RKsUkWSLvMCs7wPo3yWMNM4FWXDfsHKu5IREiRGPHuNJrNYN/+
naNZkanbxATVnKOGaSgWTJV6Po0z5GbqvDtq6Kv6bTgnRcw1Kva+VhtaczyA1qTG
REbvY7JFcz4Ze3J2eW1jbVzmv7fPSdO+NOTuNJzBDuingePfgeDiYjS9MvnfFIyd
vuyAiFguPR691CXegC2YNZfPfj9sR5akzg8ur+EYfXqoU0wWSnEDGNiRUgw6qoDw
loCn5BJbbY7oSoKMOc5Sn2EEaN73QEVUJfw8IyE8xXfi1DOBuMXEWLLntbomh/TX
d6mGAapQvlbJfdgxl+5v2lfIPMM0LrIn7rDQZLGp+wxvG83v3rkc4eLgAYMALZqK
juHN4V+s6Dlgtsv5ZsY0BMOHGo+zoFK17+ycSKP3OeY2iCAHULFwFELvo4QgUW3d
pqLPx8XXAIdBkBmzViVugrQYIz7q9aTd1h22MVmvsDm4YrhXzAG4ptlnCGBH2ZL0
tJ4WgbyOeL38+Fx5iVAPAB+LxOKeHDovfhqStdXT3zM8MW8CsRgpW4t3CHGEsuFk
e5W/a570rQJPmXeNge13xeKIeZ106KXskgk+j20p66O54xevCx3V6uaFZtbyeqdR
6q3Cxz8OttfVHF4xJCV9J13tcAsjAsGVjPSP29yeVb0dVM0qSh2fFSB3pOC3spuJ
UIYaGDwA3vF9Pu/w8p4iy9wnqJgwIDeP3+Iou/u4unhs1e+G69CcIDoI7bpLbMyx
66kXoZuAlQZTX4JfSOX33THvjO5B7a/UxZTIjgHUXlYLxTVXNgBhBSdnnn9UKBjv
m5rShXTFyy4DimFndyS1CGI71HDJXTgZipAZJ8y3gDfY75GmP60TcP6Ho79GwRBU
NfFnnH1cdMqWl1UwzNqcEq+N4uVxefCWn5SLaUIyiIlgZVy/M7ltd/F5A6k5R3kB
HyZmcZbLTPCzi7KryHmG+djY86OfnXN0mIdQ0eu6B6O+kdSXFh+jR2zGfxN64DDG
/xOWMzRfLzS2bVo2OuwdjKbqQxzzLhP5jEzR52AkixPYFpmH/joTaObBQwgDq+kt
ezVYlCFsrNJgFE/9PmWzvhctvpONtsaD9lbHkjsJmoetGqn3a5eONKK2WELetIJ+
0AcV5OLzFaMWjmXe2mw0V86qZF3jRtjhd7T622kPkHQ0KsWQrw0Q6Ushz9r39Sah
1cwZEF2+dOPWmwOIYx5AkLFmTVTSvUFRtFDA6ltWbPrEVoWp1Na1DjINGN/rFNNa
I3xU7qukGU6CQUjK9CmK6tOJvHmnJjqIPmiVFGEyzG0Wbw9KTno/7Vgj77VfxGgB
VQTnOA65qCQYfkJVsas6XRWfCUYyNFwMqIkPtZY6azXzmaCCgS11KwBPWS9IsB18
/b8YOxWIN7Xz2tp2emyDKgM0DJMpFfocenBNTF225JhEr0vutIBcS03KPYNbJ6sG
3qlPFH6h9/2NdGzE1NeT7MDH9zTpgvJlfXqbWXRUsL/5BwncLAMBr4K6FYqeY218
qElB7mSpIr+x1fQr39rAuKVZoWm5YpNPVXujetwcCqClqxSwi+I6PQBP4oqc3ePZ
Hn9xRo3clLY5KDTnrIY8lJfTCA7F3liXTJ3zjU5d2IOF0I8MCVmX9QlDfgmlodmO
68xi++IPKS/V02WA6PHtbzBhH7QN52Mz4jNKH6qKRDvZojMy5dQXvMEwqVYkGGLn
2ZydlOheK60lbJd90c0SHAsXhy00UPxDhkBdLZW3Ki/DQa++ttJDO4FchsmNcoGX
qrBeTkIxnn9SeWSvU5tHe2V/daOCUbFHWOivRok1jQ8SqSsQ+9Tdtcz+cR5AoDsT
69kYqJbjfWqhAH6F7IsJARfDKXL+mlcS7l/ZI9oN7+sdXAZ+9jgAKox3/d1eOkus
sFDltQjV9VB4CvftSH7kbc3sY88jP0WHt0y0B2anicZWuyN65XFzXG7TMMhN8ut0
3B9lLJWOEkQPwlI32Rlu95nZJyr3GkUNNrwypzXignHBAuj0r/pAqCyog/KRZcCU
F2t23cuPGSP9MG1SkDEiQJBcs/YNHw2jqer+DnzJaYzUZmYTzsKGMfxgDx/cQJsX
AEUI3Jw5R5dlCk2H8hDUUAOvwRAMVEiZUxk0OMAJZyo8m5ry7xufS36NLSjqqMLd
dBcRL+b1YIbHVpUNz35nZcLSofE38Cl18Qm9BLPphrWmNKLbYfFRS1OMseuEaG2q
bNlDyyNIN0FxBgzkBWfHBHwqoI6caTha2UkCfGJ5ItYm00k7BCRCq7LMVW2Nfba0
lsoAQVs5OPWY8L6DrtEURFuHzxyFGaCpvgUEZO/y1zDW4sC3rkdDH7yvGn3jNStM
7OtqNgHCRzBkQ1Af54ha54ms4qmdcafG2l9yavxg2NHEeNIxOmkyViBJwEXFCafe
SWGJd42rQDyTkXZVURGW48Er0Cuxv0rLikQBHRZU+5MAJOsWtO4qXozo0BL3qUjP
Pj4H92XOb73FsNBi6T8oh5i5sKP87ZHl6mrefFrqIcAVC9kTGZoPS+5aKbCzAhwc
dr3WGbeAVaCXlFsbPlcJ4MkIn1yUSdPvvbmHSLbSlp98UrTaKZ/udvwpZe89zFe5
6vKwMj6V3cNTZVKKqs0aoBjpdQYZ/vouC4jQjfatFFIGvw8iqUBbkE17vGjM2XfN
Do/XSR80dKm1ZL0lB9+f2C98IL/kN+j8c/3rGLJ0zTvD0CuSOUvu44EFy1FmTAaX
ACi/nRV6vrpjkHHsRdLYmYAz2/VyVAk7UbbREAyboF9CedCJD5ccDFL0OuG3FilA
wBqQeER2z0PJN/VuGpYyJeKDiMUlQwN0Hi3V1gWISRXxJ4iWreHr1YQeivlgSXlt
MSryb4X8cxtr0JXKseM9Vw2lR7YNZhm50J1cBULD5+vBypneJHLEDu/RDUPZ7SF5
p4vLq6uFASjA2n4k15fkRpT7HstABfNmz2VLHZd9meJrHS9E9hxWq0rIA3dA/7Bo
0MIDSaMtT8CVBTzYLNFJ4jx3RbbdaRqzJioBcRvsmrQa2ew9RRBfVahWGLY/Y9mR
VINyS5E5Oy+a5R0y5Sip5TSGWNzCnaTFcY7OYWAVNG0QSic0Oj3lXvv2M1K1ebWk
i2OnnWFU0sXHHqFMTAh5xFYa9qqvjpnyEAIDL4ReveKzox1jS5PgOKqbp0RuqAmD
OEh1yFL7lMfqUpTvB/I1O28Dn8NDI71NHp4bUu5Fx/DONv7PahSLb0d0NHren6lP
RI4A23R/FiWWzsA4SS7L/qLF2vzwzWD6NRjPIl/SqS0vAn4utkB0cd3VeLiGNvl/
4357eTxGJk04HMbF/kPyKrN1vEWq8tu4qnTK/O8scMAw3jMQNTDgSCfKkTE5YVAL
28pBcBFyWcK/NvJqLrfrArZnN6MOLKkBV8shMxR6lzh/epOZB8Vv1+tvfmfSjIeg
q0xLoiIee60USH02S5qbq1h/dyo33YU4A6qEvNUYdaoV+WLq8a636QkjQRULhUCc
1ZpKQ82cXo8q8byIlOX7on5ymGDJi/d79ExjkfNH4M+TDmVFF9y0WfGCfCLScZ6l
iwKY5KIQ11vPbNgYBLHs/8K4+eaDrsA6csOgWp9GrUjMxnkglDd7ckQjB0XjOyeS
07tIZS/2G1aTsnwH3SYIJ35ymbwX+IzaL7OpNih1zgn/dYEBxe1jjONNFbp11LlI
2gjBP59R7sKTpNO+/oYWiq3n6x+nmoSGAmtGVm+MndCdlkm4tVhbKMZ5vyXlECnU
l4OZwNzYPsdXSCnJtljBsMS5Qg66rIugJ2KpUyYfsJhlrk4/yJzfqL/1bFLi4YGU
rHGxDa8CIecOo3N+5n0Lw30Xo3GNI0dresns6C+58NKoESM6WH9aYx63mSLkzqSj
7/K0dbwIKo17fz6bxRni/pRzbCDsDC+V2QFcvK8sJOXvLm3KDtZ1l3bWU0bYV4qQ
OUD7XLhb9F8LEB5ugcvwHGhyD5RjCumz/SmpvaPoBYj2crs5xI0lyMxHEoH4SMTS
QdpLwUDUThibCV9nZv+eSJ43DIdj/XQ4hMO59eGOrIhk2VZ0m3o2Oikja03x1AZo
sB0Pj0/bqbCJ06pNqIcXHNZlljnPifzO2y+OpTITYZOg3uV12N7Qw729FurozcJe
WHm64vyj7cLhKSb04A7eqrRwAej5S4544Z9VovfTZhTcj4UnN2oSYLV6AjksoFTP
QbQc+aHem9aNCVvSHBrglGH/iOgZrlEOQu8LiI18zNJYEQeLGQae1j7g29EJXtMg
qY48j3kqTR7N59JaKDkYxDh08a2YPCtk1T4mb3vgHMXlRP5bdckHnwQ/9TF2mWAT
CpA+QCuRy5hYjLgJEX4EB/wFc++HfPE83pkwJUy5lo8BCVaBNi+Tl+/N5xSiSYIb
8bNpMQAFm4dOFurWw8/QuAQQtJHNP5gRKrBWrACOZDkoW8iwuUMlrIgKrjtBlOKT
YWAu/d0aiPCoxAmGCI5DzSvac+7mnZ5l361n75C+mbf+pEJNNi0FygSPHdkhNd8f
MXWsgZCpsa12s/kz7fDAocvEdXKyBuZDpCZepY1aDviCKIGYMeRj9Ir2+L6ADlSJ
qqbWwqaHVdQ2jPgocz1G17GHoRBgOPrPEYjtDQMuTX9M8QRxUkIVUwEjSnjhDA/G
ufl4WA/eSb/qUYwSi2KIrhD1kTEBkreHH0otnPK+2x2qDCR6PEbQnJgCfUGJ4Q1p
fDwH/bWkLwiJdYswnihL8V2RY42fRogIudxRx83b4rewqjBDzIJvz3Ct36e4GW5X
/sOfbLy8Z+z84BKZABZRBLHjaRvYgGZqKlRAIorIXsMjvvngyTRTIIO3su//wx26
zIu4jFalDy9OY7DU/J2w64I0eP+rA12Z7cFemu7fu9J+ezY1HJn8TC9N2WMXDWK6
9nPqIuVTIRCwMtY4JHfYFaaWcT+SwJj1qf0kLLoe7dJcbh5gX2VaV1WAKCetdH4p
Eiarct0pWse4XLX+5BGq6n6qozcFVN/2to0UOG0NVt1M2Jl8tJ98zfGNRjPcK8UD
SpvYaHAQbtp4Ixt1EbjYAEDGQ9v82Scjx8nfxdpOXdgM7trRq+3PTOCfTdMve0At
hXoD3Oa0wxxO1yCwEjm8rS3f4el2HpFLFfaDdvCzMchCiQUCfJScEz4RWaUuAmsc
TnYYmkejb7Y7UsiXfGkUVaBfW8fbVjKQA2jGy/H0TGvAFatIddi5INgEHPCt4QwF
opV8d44KEnubWvx+tn+M3Y2xqXbakdxgdpeYj0Jdo10BSLvSE2qJUsIYkkgNHzeP
2erLlTTQSnuYCSJrWaul01FAc8LfSkeNq6/1x2iL0Dc9x+lvPTbgAFG3up/rrGZA
W2W265jLW4dD5iXtn0zrjNvju/nzeMIM+D7dDQ1ufe0SYGdx3rdlpuaydXbMbPdt
7/9yYoADOY8AWThON8rzEg7zvLVyEp6u3bOjBCFSlYSHYP7ytZI+dXCpT0rE4u+H
jix1xKodDzvguzGjFWDlVnczeaZ/m750imITr6twVPhBHqnJoXlJRbJkDt2IOiBu
jjPAP2pI2Na2EPEVdq4+2xzvauIr/uCcv8vxnHV04W/+Q4ia/dWVJBPknVC73Pqe
wWbL9G/xGGZSAYsuH+MjQ/fhDJTWIRjOThj9CSxiecsM6FXW8ku7j5JE3pZGOh4l
LhITKto7crlX4j7robZXQW4FmufM3lBQdpp4JCYCwGs7g3BZUpc7uq8VZoK3yiue
zVJNpC32StidP7qJ7ZOHb2JJZfh6NLung5hJPr+Km1U0BmWUOpYPslwJp61WWdLP
a8uL7NH9L755ofe0bLSz2LmoldhOsOJAScg0X3M0qW/M+HQ/ivRA/Ge+3pP0yKSw
Wo8mJxMgsb0Per3Wc7tMiLc8QYMZU7iFFg7Z+X4KsvLPKR/bCtKDhqnGXDbimAwe
sCyRM19dSMHjXfVmo8kGjFBoZ3kX2SvmNiGIzvK12v1P48zL3I/FlwHD3lC6fDeO
ujgLhIJ6vZ1zEgg6nWFjCgfi3GvR8z4NiiGexDUqdyf8JkQ0Y9aQ3Bv5V/qvoORN
d6USs0Ax+57o1P5mYgk4HI5TjlFDvQfZPzXvg9pspCT/7BgJTWxmr8oCEKvu+AUI
F2YsB6LJcZ9ycOwqzkYd7kPGY2DwfRbr14bmmGxc+6g5GRTYipW2llfrV8p8nA+2
78Y98c/RgOeQm8y4f17Adhqj5SUCyWjBrJcQxGPeg/UKK93ZQA3GA40m58u9qJwl
SFuEJoLgpVG8wgFFkLhCKIZWU8xnBLZr9TbzswNGH5Mij11R0VYb5O2oXkf/GeYi
CFjogjyC6SfB6hbaxxG1SYV68DClQdNAYX8XRtbTwyu2zhfipicn8UBzXCuu9lQ0
G2AV85XLrj0ZkCTQzfKKcZ86k/i8Y0YNIATL7frvYc161cc7okDJgAFPPzh5ethv
uFv5lK/uYQXANzmOj4M3Kmgj5/EdSOnaiDOM1+rPk7KZOFOOSeT2Y2vhEsaWjZHr
C9cZZ8tIv9q9cgQt5qKxQ5EPu9F6JmPoWlsM/A5LcRCWahCVucccp3OSE2MnzXqU
K5Ic0mQb8Mi0DDSAbDEPr1aNYMxpJVorHfwSgXcqwFiTuYPLTrJQBnKZH/vPu1ip
o4s+WXIyZVWzofGq9SsYQ5nqIi1dKJGMgxnx8vzMtJmgICwkgRDMmJXQIeBXTHrV
PCxXTbSvtY0wSi07fkdg6so5gpd1xK0tenpcYTVcHqR96qqo3H7To4ziCDYcUC7p
jGHjYmMtcVWs6OE9PxuuClaZq0XVLB5iGvGVg1N2kAjSLQSK2YUiN33d1FRC0NOJ
0z16i40Ay4sz3ETwMSPqQqgyx1+sY3l5CaX6xvzSWRgZGEmbI6jkzEN548CR38dD
96g+h8LbNMH/GjiK0kObOyqRmN5BVwlebwV2Byg32iu00OGFIOHTGogxvyHgW+eV
AwhlAxI73aJl8Bkd6IkGZkBVkgu41cPbMfBNCx1UcABf9YebzKW+tuREVJduJsWR
P/q9w0RbBv6NEjpk9KAnAkCS2iR3kwhl7effOX9X+JemzsV0DjilG49Agb90xOfK
a0WHm7GmXadu1A4oRfpEqC2frE9Ai7Lhhg5eBNGwj1DkvU8nZqchbl2J5qzc6z/i
2p9mcSz/f57yNBpA//DL4PHoqeTeYVOOdmHfd9tA4JJ16TwG0gNqSRi36zTkp12N
NHaU+ymymUh9LVSZm6ioOI6dLCE7a6+dyBvjjOOOpSkEFmIOaQhMiyzsi5TkKjRV
n9s9X6Z2u4S5clxbjILUUyQqHFL0WT5N+e1gL3nOfh8xUlj2MtPxQSLNwYbCm/RN
3DG+D9Hpx+Es/qmZrkl/RKOKYBBQBFI055Z5SbXhhg+MiFLFEnkmmeAaUoBxa8xI
A922IOQ7/QMjCqciGdogHORTVNnXSBG6tdrDZxBeNcQhQwBgPIdrueH9Ft17BEap
O7R7SaLJ3BEuQXjnLkRRPgcEI9fp8M7+45j3HI2/XOW99QAU8RURIjbPRtHztlb3
dNxX4aWfssKgnI+1lpC7+rh0xm93wYTIEI6KEfTlbw3ygzrUPRPSEM8jk+5hzkmd
zBf19vhUal83YTpCvPnvUbn/ZB8YMUXv2LWE3VRJtjc1MrDzD/0E6Rzzx7UcqkSD
GZ/PQ+bF+tOElFMWtX+dW8esP+dRVerpibmm1ky5sagvQ0+6SImv2uktKsxGuEsI
4RV5VPB5PV68DLMky2FtIIfrkPjeZf2dK8elLphxFzh7Gdheldz8d8zJK6DKXUMM
7HFiwfzc+NzvygQh4jHNNb/0ZtCRxladP+RLffqXIfvsjY7W/m05vO2xl2V13SCe
t2HnktU7bXwbN34w8wdliuPKM3aJbDFHVi1AZ0TPq5FnMX3mtofxJjHKTO2cZKN1
1b6WthT7uzhURSQdBj53M3OHYcT5v1dClq75VQtWJGm7I9iapE0Co270fDx8i1mk
00dA+d7FvCUWhjT20ybHfT2l4ZKGyekxnbnQkWIZFvqiQUhKikMuKXHWWsMdow1+
YvwSzVu38neS7POMFd45F1BkLzJ3e+jYWlye5jV/yNy7HqXGNXfpRSOYHb+LRDLH
S4IPgJG3WFLhwhxz0H5yInSnEkk/ZAWbTADYHv7FKkzBg4nhCyYhFrE79o11UnMB
IWYCL3extz9TPm6jrQGIka1TvbEMrUrrez6YTIqVL7LokC81Q5BLdVXATV41QkIX
2qCZEYEzVQeud75kQEy+BM1MCpmqEuUMnLVUKTQC3lciQSrgF9QCKE6QlNBcTXs+
GVMp8dqxIBa/zXrfgyzBIaPxFpUPTx9llx6N5Ip+Q4DQJc43sNN4OIQ/irsAJWVV
8BDhda580clvsmGbCW8/fCrMK8AzG8c5Fvd6YmV39pJASZlEcQ2YAaN3PhjODaIU
D3taLZztTRglF22ivbgwxtFWna9G+jxtG9EjHmQ8JDvEWXPX1mYa5QU47rzfVKbL
y3RZtFLOo26vy241jHTLTltgSUPpvfqpyG2d3CGbxcYOWCdHwZRCuCcqrD8taU2B
qjVc7BsS2OGV8OWQIBlX/biURgridPjqvH1yUKIYyzfCbye+vD9nroZAL2Li1qX8
fN3YiLUl2jeLpiwMmgvvjKlEctPjKhZnfBDCfXit2lv2puPW0YkSVwmCH/KH62Hk
joCzN8tE/Ubrr+g96R1pPdDhClPzM7wkPfAn6XOIGPwJ9nuzshi62ayVuRYipsDT
x0MVhHypFNjfLPhxCp+zZpEb1R0IxJdjVyiM2nqr5Ps8BmAOCg/CCvlHjWkG5O3O
DeT/GNajSoTGjpMqLK2rSwWIiL++MtIL8zm2TGxGKFzuyLDzkVZbPTtuwRVStH7n
YqkWXGp3x53QZ5Udjsqg1LOQ0FFd9omQIyU0pNrbj5EmacDQvJ6BBGFcsyQ5j5ER
jElx2gdYCARa7CHKYqGnQtrZGdlGQLBFkkRQ7/fvAjwiqMYvAlo9af/+QJ5uClUC
Xs+Ao197UqcPg9WicPnrazcJhVBxU4rn+br3l2O8F7xkV2L3WXbMdlSXrwSxsN9C
hCOOKB0vQjUArUfVOghtHD+9bmtASe7W6mRrZdcDYDPw4Ts+a1ciBT2edtho0Wu3
q5GbjVeb3KRwA29GnvnLqJm5LILBtbPOWsYvjR8A1wjFeZJ3FMZ+En0AdLEL24lo
dFOp/8R9Jkaj5Vqsg0ErxYA62C/iXfW1mmLXRhZTfy9TJax0ypUBY2Msrdil3Mea
fKho0mK/7qr0UpEybYM7QwXNlEPpSCWmyFyFBMfUPwMDcs7rgmQPoISIWwXrMQrQ
mAXdfjGDTvzDD+tac6UD+HI0SaR3EbyD65yO7We063yORG4J6YLgEmjTeWedu9ff
SlmR5yC7YobdXNBEBOdv8F33CwZmxKdMkGB15i1A3YfBMk2b7PpLXfhP2iMYpJUW
FUV4YHPPZjO7ooESQnae1cTubIIMc7fZ4F0So3/pxqq1eEgl7X5IHy9Emf8TiY7F
SKqITxnzAxY2HtbI9zjNYn+/rPVlo118swBs3V992/o/bv2qwo4zv0mWjje1Y88B
qRvuJpPG9XYQFqtZxo6MmwCPYxSCBi6r68a4LRNJ+rDs2jobhBdcQ52o4YT5ZhDF
4VKrxFf2Xhpgg7Xf1U1oFhQP6W+COTrLgLZIWV3Y+M7qYbY6s+K/vzqQs4eEltus
UThH+IOio5LeOPDSUony8qYWG7ZY9mWdmCu3x7cQ3Z0WxpYCUBVK6ldfvPUT9OQW
CcJXMgrJ4NLJrzAf0BU78OPGu3lFDcSydOMpwPG/fTU10Lesyfl8D2qhHqy2BbfN
1CWs2ziTrTG3Ku3WG+vBWvGFj4HYNwu980j7pOrd0cM/FLqRkio9id89zg0bVK2q
fZgNXjPEBLWG6tKfnzdydfCUdPBVbhHd0C81B4KAY00wrdWhsoodAVOsbZnVWJwz
BLMHh8Xx/TjAzLTS4As5O7UgEFHYK+4A1Wlnav9YhrxxGU3vCmfnkY4M1Rdnkek1
pTq5SCD86MRDlRc3hbiLghzDHtXwGJjDa6sWzNgImPAyjN8D/sJCvuP6Bzp06wSx
9k6XzcKnZZuZlpoWIH6RjKSEFERjSjQkaAyB7gT5L9wxd9/Y7smf8RVNn8WHEp9G
1r/CAotY+MuA84DdhPOsU9yKfmzqeHjmxvRJb6MK9FSsR9IdrNubjFEBHngFoiON
OArO7lj/1wLBe9Yii2UYftIL0neALuvddPEfLpWwRMswEgN2tsCuJDby+W5LSrwW
EfraN2bQfDXHK+pcJ71Hnnwr0o3r7tQdRoO3u+Zgj4vluOZ8BcNt+rEAZPk6+E4y
DN2akASshtaa5PI0ZIJ/T52hWSriGK90nsJrWabudRzYqt6nYljDn45fN4zW/c4X
IB6BOURdFJ0aEKKbffwymEpervVGiWo5swMUoua5JkNwgOML9M7TbxC8dwUQeyk2
FPV+O+SSF7yqPwooBWs1Q/ocJ2h+N0Q/+FQYLj6hHw/apxEEHMGiTtdQhDftbYl2
GUhloH+BTXSSkYKOzbBDS63eRjFVh0EUVCnbCXWx0ILkDQ1pzPMYYgVOjBBrUX86
WV5KmMwA+gk9YgB5ntCzftnAeu2oGEvotuNJjs4KK03B3JUKI4rALO1Sj6+3oJO7
+xzvRVrDs4Ibk1QxSDWYtkAjkrK08N30gOY/lnSI9sv6Ag69wzHLiOYpKjIkesRR
LFUx9X69qeogSLAejtzVqjNz/K+D2epoWcNlOwrB8VxjJC1lqdBZ4kZT9aNUenh6
UK2MUg4WjErQtWrJXTSAUSpKU7caEGpAQou8YpCQWlZA//0NYkuk6llzheEH8Ypl
i/e/s2TyA+Wn+3tVDoOxgF0jj+AYoOFipKkm3xLCzG72NPTcQ00xpz4a0c9a9Aqn
5BQAF0EGn19ATpu3SO2JrIfe/twoWNwFkZ4FLPxvvff6sVat6DjQ/qBSOx8j2bX2
B0L4ParkNzmQzsQduaCXroCM7ix8MziRTpB/GFHCggNZCDmV3htNfYJf7+QL21xw
R+v9OhV0rbD5M7nDJzy3jlWIQji648OA59auIBJh5Z069BYvtH3tTlCLghYbrUeW
brezM1gXr4td+WwRsbPd2dKFmj1YEYSOLQ34DvLpyEele9ePjowXFIJM7xIUX77B
zEHz1I002pX8LrcktPFX5k464a7qTyGS5242P2bVXqRk3+q5kaV5asKCDmCUF32H
Zb691lgucyV/yU2mbSOw91lKUYgv/jPjtaWbKVl73BNhVqEZJQq+gMTYkffx9u+N
WiAGYoGH1EYKPkxDy/jiZdNrvkuZj1zn8hsf8oonew28ohBcWyvGqMObj24K0nmg
bqYpjxNpDC1EM2EqmvjTnUW83P2muVEioAyvt+ZbFQkSszyQEj0uBsRzcdHpgkkI
kvviGdhC8in4rqyPuc0kjlHAJMntEnZPRdy/r/svsYZYctwrOfbXFj2oPkSdQMln
Xw4TFbTR7GgGRsCq7jbu6KOCdLs1Cui+7sE5NbGH8D80slQtAy0DYqFUpwo9ltSs
mdFkDzeUEijnVf8pkGGz+0T5aPczRyvyQozUNJbqZUxTCmXSjrJp0lAR5AqlJZly
Qc+lTGkT6pJFgbiS3mD/FTUfqxVsqrKg3GvXC8+MkrRHseEvGRAC5pKgWshQvBrJ
K6KneSdNwo+6cqFM8gTVYkM/Gx0wWvjQeXbHBN+IJVRrN41+xGoRoXwAjieXRWAk
An89t4d1EzgMB+WCuAVMGUMevWT4I7gr/7KVEKS3LXegJn0R+G4mfgBCFxV6CBZJ
J7pidz8PhR8hcog7AMDniTMPv1pqmoDaNtOw7rsCCgs8fiGmp2fK574f0FKbGcuc
VVv1DmAjrfpakS0kNdV4xk+DJgB5Rt2P3W8Au1M/B2arGzdAjp313SsXUeGpQx57
zrMSEcnG0iQ4CeAlTpl3iyQRWsDICHHaLn7TkjuGSpsNLej4oDsv8I3ZffjTWKBs
9SLPpGGaWnyANj8QXhXrJ+1G5KfdjCRtifqynYQ7w9JHtVHQo09Ny7MscpD62gZR
rOuEw1b2aO7KJZWtDrDtez+umtFGL719izDmsx/aWkY+WRjpMBVGHYr1uc/LMssd
rLpv3rta/KQbBCRCA/XHXgeNhAwuGEcTmzXWhzyPvo6HmHm4aYme+tJ2lrOdTXnh
g08/yPMK0nUqTBO3WhFE4PkBnsTZ9bkqwn48SfUJ+IVYMJKLZniOqIyAbpttl6c7
l5+YB1X2AsSYLJn2FGxen72mqLwsolfS/i02ZDenn6RxcVl2wrERhP0GB61Y/XCo
qkv4McH8CnBbLi6NSIoDh20oSBeVhlVLSWHMlq8emna/0G5OsrebK1RRbrA5iUej
Pmvf4FPKxKXAfCubu6p3VWMqce85NwryeA6OdKp+vkzC3Fd+d9xRPMpV+8KplQ8f
lD+Ap/dvSaOnb9fK8r35GBu/vXW2yUeKsYSS7RGb8mkngcpJkrTTLXiOzULdXapz
m3mMODHGxhlpM/57q20iJvipFSzPggvWElHfOIU/M32X1ZiQVQ/hCvysMxACdb3t
v6UDjJxI8xSHsre5lbRdKgPg/JaKek0/K9NR6jIHoYLX6u8Bwgi6XRlooMKydbdy
SXO/tNTqdWSDZm6TLrtAskralWNGpV51iC1bNG0R4kDqrGAlIq7jvuG+xKm0HZjQ
AmqRZPj1o/YwYmrPAhfrR1fhd6FYMEElOrkXZ/YXPueG9rKjKCnfuon/TzFrhict
2+8MlFFksPJaau7qaJCbwz8ml0b+wDE8Z1MXyhfXKxeuzjrBAKXUJkmQAmzbqpCg
morf/PO4rP2vewY0lbMc6WNWppIUpQoevhk4/gLVIeTThTyRNBKTI2NHZq3TPNBr
lMUg8bGKjxWpPx0Grcxa9R4vbIEPJ1LSN0lvfWnkGJrjGaW3gEze2qvV4S88KBvA
2CtnCn+VvfQiYG+lL0Fy53fWrvron/OTC7VvuXD/4knUzWVTXUfeSJXINSJgHk1m
NlbE9c/zbRGVKptDg3p/c9kQEX8dhx4QLRcr/WjkoG1ZBQ9vQnxVaiUvj74878ud
6xwNlsMmZ73bYFcUeDrHntWsTbbFJizmjSpJ63T8JOWxrm75SV0SpiE4g3fjkERv
HY1EX0o7cYr7djnzBq+iNMQt+rFDGsJvr/H3m21qD96eZ71RggDRQg0G3FV4KgMU
KBGLB2MKmspzSqSN2gEw9W0crRI3iXVClDpXwX2eKbvYVfLijWDpQNOrqiL7+jgS
ZHPr+3Tdjibn9u8qd30vTmys/vMj+9JZQqdHHfHOUbYAWjwYlL5ynC1QkdROAUMJ
7MxiXjd1JUvy8WynzBRzXOfM9BwlI5VSH3QY0QnyHhigRdaJo2V8NaQ/ROsNigss
g/WvEe2gZzv1gDTa/Dio650Ally9Xrzg7VQTHpFqAnfVj14S9m4L4VYv12SSEjSm
qUkcGIrqqr5WhVdeffsEI1zMef7prDIFd8/0y4wzic2gPdX8DOPvWEnMOaKaHzpX
mlR7s1t6LaoJc1Q+ux3uWn051rYzR5fQuU+0jUaHUgbkKL5/uI+GilQrdLivJEY5
/hEwv+4yHMBk9179j4nJo4op9iPDMADojankwMIefEKpaZQquveoxmXQnsR5KG7s
bm/lb/Mx1lY3jDbaVKXP63PhB6v+13+KgajI9nLY9aX9Wk7xpUGWBUCEs8YrSI0G
DDXpLsJwVs4hqY+H5clOBhkly8Ity5SICF1+qKqgv50Tw7Pb0Qk6+Fq5oX8k+uPl
PzlOQR/mEJhhte2Za4SgwJWdsI1DU74TcwtihMcN8sOFJqMTdvqmhQ7wQossdnok
jXtL9ciHFs9Wf+WaQHd8BMpi6pY31qRvxq9gxyfEUKlZPlmyFwc5W7cwHFRraS3L
oxvoD/0nFmlYSza/QPCGXv4PG3Z/WirFCSinyDG+H67fmyn+TNHY+/wJr3XQYOB8
Jl3O3TY0p/ce4teS9Wl1EjDrXJAzKrpCeREM3FfxK6H8MHTzSu9Pskm2/VV7Vnjm
xWyB4RxpwSCqSoeINak0L9zygm6aBBA5XS3YCRo9Kv5UffAPpSG7KP23KCN2/9MF
jlQnJCBvQePFz4MV4s4ceB+PdGv1V7TbTFj/tWwCjVoRU1VBrpIpagR73R1ixC/H
1M0HADHoNj2g+0qJBoSmVyj5DdStmbGlVSrRmTvt0tMRMjfm3KAwqj6pobWy8N8T
/8mtKwgKu0zEEt26C++EfjNQI2rPpeX8XAVB/NCUlAIYojd1NRw6ynV3rBXkibq9
lPcQB7NUViIuGcFMNGWnFHv66sdzJCEgA77pLGrjsqjkAJ9SGRHL0G6skovXStql
74TVbQhVmwV8GghJ6kE+Nn88Me3yJvYDZX2a66XIVkCus+2ezlTayM8he8J3xmZl
qJ+p9PB1Y3gXgimoS2mTGDovELydRBrVb92E1pG5K8IuOTLn5Mhrs/iGSSk4Y2sd
B0uKMAOUZ5zRPty16Kyk5q5AcgrkH+ZwbPgwyn1xv7Gles+1xEIj0GJF2+F9z+y9
DmI0LLxy+vIfGadwY2Ijf8YOBNyDSAIOLjdCDY7CXeIAzXL739am/07DgKQMGkKq
TtxzBewy0dfQNbgDor6/vFJ5GlV08sl8MF2JAbfY5D65tC3dsGTIyPjR4FoiC1V5
DDlkgbHC8t85jRZuGRJWs5qijKnh/+mOcoZM7IfrDB+bAQDakDdMaQqQ1pjiG9DV
ldUmpKBd23+AHYbLkApOVlAqz/SVCrN8L8mDTSkpSdTdofkqSNrr2x4KRWuIvuVD
qjYDJMgAzSd6J5hvfFjSRJGFrr6YcMbIQBIuoppbLatYd3Ak2gmEyJB/BlBp0PsC
HM/UdrQ26NTEh+rDEMMl8V+FubcgSTv7mAk2YvYeHO9nGJlp8xEQB5qp6eYOEFyo
tHwrR3cpvUIKmz8qQWsVFdQNKBZE/FqanjxJ6W5v2g4gKnBVnWO6EXRzIOgKneTh
ptmBcIRpfLyLIGP1CAc6PKZrTH38lPmHRgeT13ALtcw+L7SZcm3INvhC/7jk1Qyh
HUiv6cKA81wTO4h+8k0in/+9f+wiuvZQsf4hq4vTyEv+FPWnYLc8OKkA9PyDU+aH
+6cZ2zkKSj3HZXSfbxeWKxpzASnGMBo+DbA1J+qorUMgeRd1OlxXo0yLBK5fSqo2
YhFMXghQgM1e/zNQRE83OMbFyGuQKDlhLuaMDHxGiw+Zrfco6QwysVp9nZZHO/r/
AIlnpO0bFAvopW73YmTCzTeh5vsWaBKdSgADBJTMdlDVLNO1AG+mFg6h9GWBe1m2
4n9UXEHjM0Dmku368OHIQvZOYBs96ugF2gckRhDaMUTsaYGjvt1Ocg0//A48on9j
YhvQnvP3LU06DfKJROgaAdmV2cSgDwJ9QFMo5WADEQ8hImIq2H7JjecXCWzVYvKe
kOxEL2aUvvwI/0u254PlyCrlEhmvnIAaNc5VrlsvdkpmIvWXGs/xMkP4U8wTVqD2
KfD39NC9tS2JA3z51Quc1TU88ChVAN36+ypXVsGHWQ2jkEi0tHSMtOc75R5O2lc/
AFuDBGt5wikJpAUd7dCi7JvG/xVEJ5iPV7jLVs+N5uIOILtyZ8MkB+pEN1empVI6
WzJOFFfuGch0+l3TlwdDEgjwJiIj7iW3DEVTPiKN45zutLpDy1pizjkCdCpzIazn
PvYKj/LtMX/6MT2hZe6LdIJ1tGGgFd7nx8996IDkXsKtSpg9TUske5QJaWp0Pjv1
uOd+7ik5BEfKMTxxmuKl0c74J5Gr/D79bxI9AmYiWkMW/OUBEYARASWMcxymLH9G
BWdeBVRBq5gVRipG5LN5M6npqoq22J4AH8GlLfudluuBusHTl3RPQ312rv7/rimh
2hiqNi/PK7Y5GuNUuA40+bBEWOcgfiHHHra6bAa+Bk1S3YpDQq4T2V5OjsqiYLkd
ziNiBtIuKmQ0HeOOcje1yNxtTijyC6GcVxGJaEKtPv6InICHAWQLACQILJzra0D5
xDR4xduAs0pU2qAj0JuFvRHGAVG5yCo1fNP/qwbD8haktPGM7OivEGBIO7ijDrl2
CME7HlpuMSkO5dH+oY5CdCXLg6ngyDmWuFUWeTpjMkIH0ajPZc9WnacBfqH5SW6s
lKJgfMPwPct2UuM+mJB1j+gYj4GdBhMFY1PInXve4QCrCTy817EZ8Bx/QoaYYpuR
+pWkZr8dDE3J4BvUb1+tC5mwr1PzRcA6VSn8YFqk54n+Oy9SiOaumEYd2sk479f7
cFgVmLwo98EkXnSdH2R9J6KzoVPj9mDl5YKDT5ZhTsUgZmvG3jlRnFzrpyDjw2Xq
CgTpQow2ehMYVL7KBXGUy1m5aho6lCIZe+4wZbgF0O/0GkW4YdQnf4gvQCDCy3Nd
Ip7VVWTLNVscvesJ8BqM4UWuKBjRLX36gLX7HQf73whwKvc9MI7pB5fpvw2HHZfP
org9Ejxf4ThPt/MaG/arrRdvsALpb12vB6Up+LimYMMqGFnV3eHwGB1zstJfNOqx
k963DLwg6SAUcJj/MAAIqXdkta09gpbONBKLYmb8HPBjeGgkxrAgIgtscpQpRtDC
P1YUMIUPnoisLCSPz+XnKYiKGXzRCeiiTQwPMyN2yAbupTwLqlrmZGDS6EUJAnxj
6zodJmbk6ML5UbgKNiHXX7xJ9IaXRmyPCT7aaac2gVJyezqn8EiARhVlBzqI4URn
57OzmeCsx5Et9RqezGwmiQq0mP2S0PZpsC/kNQLlHS0JhEJsNktHTC7YmLIzF4RU
4T6Ye/jh04UX+et0W3YF43e/KYgryZeDAz6c01TqyhbEf7sNP3+7zRVwsYGi1bvr
0nCTDbFptHzroD7rRtgCG2UXPkfAi4iVY1yeayyqlDwLzmNTj0+3ehtTB9JMgV4Z
RnkN/ocijr1hrT81lUhfWR3Sf3IjogfLO4b1HPLblmwnkvqWzDyKI1fMLL1GyBNu
Mda41V1EhqblipMHSFnGUWjJcdKf6Gp7JX1VV7au86uJfNqd6FB6KYloA7C78mVC
KRLUH06jd6LCHR4NwQcswTODxd7CoYaMEvrOtHSMJQOqoE3dVoe1YvEaQa/Af46f
0CMc4jMjuNvTtKPmF/jXsnJsS/MLmxZwOvV+QA8gAjw9pdmKRf3sxnjAgFENQB1g
AqKHaMW35hOCryhhebTjcpmVfBc5pifjaFF1fn/VdLCt3ACfNHX7XNTlR7/9ZBa/
eqEZgM9b/qYyOezC7wlBpIiOc79IQ2zYazyk7r4/QLkGhfxXJN0Ni2rgmz/hQM4h
LRLGdgryULg4mXecwLUBGhBIRghmRe6qULBId6duJ2/4evnoRnPw5ZosejaHcnvH
poLnVaxN0IFi2TkwxqImfV2yjUcz7e8g3Ed7QM/tNTpI4BkwzCC+Hvoz8E+3YEIc
pr+t+0FWhqLK/RjbGdMWBL6yFnNm0PxIRtToAY80OC/+KQhyr2jPQP+Y7b6lERCu
RkBERqgdiPEPVFCQ/V0ucg9kL48A3iym9k51S70xAMgZw8UBuZzWL8Efw2cZuxYf
Ei7GPvgcyaa2QK3cf/39xg9BMUWNmsRG7ykqyabVGljiyCnB4pCjrZa296kXAuLS
c0rzQKBfvLN77W4Wv1gqUq9VRS5N8D+hmGT+2o0RDovO1/kxChg+HybL3BOzVs/R
YUiFEKzmnE8i6UBDtXIdUbyh6zICToAqBK5UpeAPM9hvVI1TU2J2N+Ou1DXtNK8P
CQr68jHkorNGWmi0I93EDFKX7BrUDRYbXatIEK+JKG4V4lvf2zC+ANLBkrKctaIw
b95EtmIwhF9k/V/dYd9QYg7xl7e6YRdKD5r+JONvFWV7OBVDJCtm2/7gsKAyO5uo
iQozF/JdOWprzLnRBya/oLoLnfkp8Hge2X/0pE/phdy0hOQjE06MD2jwsVpUOLDi
JamNMoifOPsAZkMWp9PCTaOQNF96hJwiPIB8UYliJMWVWCGJwR2+r/BFv0twtbao
G0E/jei0nCVB8W+KCwuQmCO9KsmYYyVLhITZ33qFJeYpkeWSykd8i4xyJ4nd/1V8
9lftanT5t4uq87VlkVr15SEZUmrEuVXrPJ9agFE3hrPGErAKiXz+oHkk/iN4KQCe
DhPe95cycqfMTDYLZa+E0ZyA0uIEAUMUaF0oqkoVEv6Ll62w17wzR84ShNO7mxZO
qC51DbYSS/KjhFSByJql33w0S7y3EBbozFfVZ1kRweE9/TZV6KdR/MrPlP4oM25/
G8PaEc1vz8yjjsgX8FgG4JJA/6WKfOEmB5/0r7yRxwfolKsEkBjLM9+yGzYr1kcX
5/8un6urG7e413I0NLL9PA4Jzq7Qg3ZQz+AoDCu5VL2Zw/QArkgh+HedxheD8Bhx
qxJgDS2xZPdOEtCbyvgheDBLaEBC3fLFCg0G0ANbChVFU0UHrfdKi3vWL2v8VoPy
HWw+z2JSmC2di/4bqKF1gnLAn7EXXV1KAnzype2CZZJRlNCikeREVDm7vYGqCpT3
eLFCGv3vwBaT7TS2BA7xUnESF6/QaJHYSTmTVoVmleYDA8BXddE9hH24uct5QNM7
XSi9RclYK9y38+Djgioovv9h0klrxwyHjnLSvy7A/gq8bzYEjvcEUIzAVazD30P4
oAWSs+NZ8RQO82nyx4Y4SXS7POZoyk+qH3ZC26ijpO5f4LhpKaiRXITuJZfeVwJu
ZAL6Ebp9ubIoE40KpgMw++9pKSt+ICIrFNF0njeZ9eMfeXcYcHIRRGj9CaIFXEcq
4iEOsOH65Pp6YyiTDpL02cC3+MvN8IL0ccdUc2/cs4xUhqGJk8oL0nMBEKtMSimj
PM9JrBMJgUvBmqn67gRmVkisjMMOJDM1NHPZRS/X9vnbk7yat/fI++PDUbeF+G55
CovU64MmLmy8mg7P+qyEMYSfcRgTxHAZz3UarFKIQF+RmfFaDqqc/qZ/i81yP1ee
J0tfOE7o0pJTx7n30QJegoJBShUL0eEDbOcxcSCF6eL1Hq0VPdhkaQffSqTL53Ia
X78SDg/7oIbpimg5FqKuQithN1PstjZcYdzXQBRZtC6jdoxcBs2MfsbkcOMUagmb
WvoOyORf5qj/hXPLs2QkK4JziZD7R8lvoJSIHWNmQrKjO7XQl9MFEiLdyuOQL7iK
sRpGVV9HqBQAiWGQ5ipT0Hclmfu/rY9efdJZmfTtXaPJMNHoYlUwD3V1XDBGYKJx
+rEnqdlf1pXqYncNKeL2eUuz6BpSTQC7tXU1W20b6Od4omVtPZ52Q2F5fPpl8vkr
Y6BThiQj5Hucs9+4fX4PUr641iRilJOIZ95vB/qBUBQiP+rsEH9Mu8zG9RG/+XHY
8LHZBeBTLIHVwyu65kjcRSLT90pLnVNUTm9o54QtaMCm3gmPEbshl3M6FlWSPhD0
XRZC/40x7TE05ipdqrlI7uGDpUjn29JsupZhDp5TKMjnYR5yBUzedrb/Dv3XST1E
B2N4W1/iFKczbZyRjMNlksLzRTu3yAjx0jPkyCBJrM53byVGrG9pVWxUMJw2e2k+
zMD0bbCOJcLGvQ3NAOLvVEQeWa9fwVXkhqILvIGoR6O0PkNWUs22dnhjdNL3ig3K
QiD2fgltXeh4gumO5sWyGzfECMs4iYcrX33Hcw6HLHqN+rsbP33+N/O1G4p1pCfE
1th096mCxzSoWwHoHWkYZp0UU91DAHsJVyAGu3+O90v8McroXzBUc1pkzgFPERfI
+6vvuEQwUAfekztsg/e1HR5TaUqCEk82jL1gL2lJinU0RhqSjk2MyGNPLuvVzeZD
nDSKZWN2Htk0W6oghRd14WcoUiaB+wMTBgy8VSzl7MKc3sFHRSAqXEGIK4La0On9
A8vHKZZDeq2vqe9MTMlTcaSbreeIGNmtli8Z/idXqyRXp8GN6AWSIIxWLwmR0tcM
X+Szro82uFv1owi81wyLhV49AjI2V9uNjXk4DIcKIHp/u9JOAUaWQlo05QkXFMaa
sBYB5JMSqyDbdreDSry33FkLJak0Zv1C7p/XYlD1D5s7DKGkbTKBqO9xpVoHk5sP
PrZnasS2FqjHLf47wATNTqEAuLyB0SLvoZiE2nBZ/mfDXxL60Xuta4H7EzBChMLS
9da+pVeGrhmNwgciY2VTpcmOqmGGVHMKfO9Z9e1Ka8wc3XBGH2+/jSpNfAtZ0CG5
016jFkJ6C/8/gUvXQLbzKUsugAlgofCovyNRpefDPh/0xt6uy4vkblDFRHvUrXyF
//9ijBB/PI8W25hB+oA23ML1sbx9d5gMDhuO6ow4uod00G+nex2axmGj1FLiFHGi
kynjhHv5YrPdDDn3amtN/Uj6iwHC/DZczSeA4C/Fda29BpP9c145QM9Oh5mn21FP
kVZO+ejQgUCqagAW5X4Z2BZOrzX4MQgGRusW/8pneyFasqDV+aC5HkDnsJVIpg+B
Z9xGUHRzXa2Lku8O7B7hZsBn0yz/NnOdqR/Hd6+gZwDo2dhaaCMgYm/RNqDOUEbK
SkbhCbOcF6zAW9wgL9DJ5v0x3y8WmyjZazGv6w1LyaX7PP696CJEJeBn2xdsGCp5
vxdvqmgmPdiZ8j5XRMzA8R9eNCaTjcCuZ6TtxI+/QP7fBrB4HAe6l7zq1lLI69Ov
BNB0WfRe91RvxoWCvtm3Z9C3yLk/rN/E5F2QXM1iiEQNNZ+HJud5D2trWKMSHylI
Rh+2jQ8DPzMOf8OWypbzD2wtNAwdk9UrKDP2ipHfbMFueCtTXTBtjW8p1BGy0bSH
8CJ5BbnEo2DJkMN/a1kbTo+fzKwfoXYBHLUUBKMu9WrHLGKYjQG/QOxrdQ8p4u/V
IGyrXTjNx9LZb2c8l1qBDnZkmJpubG1/j08DBggp6BxJNF0COczBaFvmXONCFzSV
9WFlCzgXc40T+OGr2qnui1U+DakbLEPB2xqyg1DD5T8KFbYfSZEzcDFQ84Dmxvf6
DcEc/ap4oW24N6UikAnBySuktstv+OUZMqCp8qgQJbhT/jVXbozPAj3zLaH0sj2n
CLZtvwbBp6JcfKFi6U46A1NOesN6VL8kmv7fFYGMCKDyzoeW58Liwyk6qEOP4abd
B5DCD3KO7tdQiQpXzbXCWZExOHx/TPSDEkNaAzScD3Pzsj8hndOFauZThbMi/WBq
+QpcDtrJ4I0UUHhYqZnQ2MglpKhpqaZoMYcU0VBwxeEuT2ojEkmCE3v2j2z/ne0i
qrL2KZ8+/ebiHMLLHKneYKRebUqEywV8NqcA56GWpzU5G+mNuI+6w3cnV0DMCv+K
0/dL8iqX0SnzCcB7ckChk/nQE2Pp3nuLjHsdzYuYGeXl+9QFdqvpWGBFLdJ2Rqdg
7UwwaizUG4qDIdYNMkI6TjYF5xbYACq/KJwV7Y+zC6f01iH/j7AEyLYUmyBosOU7
sooLqwb6K8TNAXVXuM8CkESBLDJe5IDFZ91krCmkDNhslqCysJipILTwt7PBLChz
f16DVDLoAwjaZI4q4wj9AbvZ5XrfD7LRSvaXeK+6/sdzhNwDaCPfNZLBSvxJQIap
z7e9xwzt+AhM7MExpt1+vLrwUhRbZ+KUyKn9SBTslj4I+NA0P6wUcy2fGHGvKhTk
HKxcS9bsxhXYtKqwN3OyN1SsfejrN3gGV4ZNMZ3DcYv5dHR0XubbR0e1rZu2Qb9S
LbR+x1WcjzfVdxFJCppMvurloJ1hAxlI5ZOAjh9R4GcK+BouiGT2gJvcMivZJpQU
HYKeyg6J8f5J+WnObtj5cSRKD/nrgeyOJ/gTM5a2ODpManb4ZqWSDGpRKxeG6liI
Swo+j4TXOoK5RVH9KNRmDJb7qiqD73gYGfPNCTMpS4fthEA4SQfT3Ycsu+F3sWtg
sQ5DsYFXCwqcE1311h5Ul88C97yEZ3mucvRHyJisFExC0uR8hJsSp5T7fHChrMPu
U86cxP7ZCticEUGQOF8WcyF4fH9zmzDxswvhl6vF9x/6FjhRWjpSRJsMc/EFl3N9
PO87levRsYFt6XkIvpmwB/cbBkf/QcmFJMQGvzJXsdZ6FIYffFYdmTQrbU2834Jk
mYHeiKAGc4vEI81IPeFIfS9hYmLhKcMCIjLPiRYjp0vdhuQlOiPby3SFuI732gUA
wzsT6K6B494BZO1sJPhZ7xBxiMRuFXQk2ovWbIdfpTg/VS5lylCjN6O3yX3RJJy3
IBCYOz1gK53ypvsqnqCUCqniTZ27zcG1q1QbKoQ4K6TPH4ZYw5Txce44tJ2tXgP8
yMNwavk6UsQzngYOjgAXN+BEltZ1n2k8kWlMMWv+gOQGRu/WVVUwUnVoQQrn97YP

//pragma protect end_data_block
//pragma protect digest_block
XFQf6916lLMGVUsdZR4S87b3QxE=
//pragma protect end_digest_block
//pragma protect end_protected
